��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���ጨ��KN�`��[��h����z\�RG�K��Mb��1�X��d2�t��_s+h�za��1�J�u�䁣�!����ef�������j�Uڧ�f�l
��������yY�w�|���puvHJ
Mg����/c��^9�����Gi����ՀEw��MXYO�rr���=5"���Z0w��.%�-B��Q��r�g�
�o\M׀c`�y85�9�gX聋6�e"�Z ]IWA��O��3C�5E�IL��!�$�\0��|��r
�Г�L��{3&�8zp�p_s�O���*IY�t���k�P��_�ӫ�����Кr�k��4L(�#�BV���o�m��s&"n���!���K���nv��'hP���L�:ZH ��X��˃MH*�=��T)?0	W��H��]�	mɳƤi�\F.��\N_�ņ��S��
�R��Y��mv-]~C:��*y�W�hP��oS�{9(�/�e��ꈭ܏�pX籚����X����"�~ԅ�qC	'�]{ʔ��oB��ŊR�� ��2�>Z�tb�Sߑ��Fgr'AНa@�n���o���r�0֏��Cޝ�d�+	�H����h։ayK���Is�G�B��b�R�Q;S�J�P!���oɈ�n�z;��B�11,���L�^���ߕL&���m�$Ԝ����(Y�C�p��@�E��y�+�-uS"��v[���{I\fPg�>�$ (��$���Pc�A
9B?�{l��ы��l\�����d$�ʓbV^#l���#k4�2/�W~�H�/a����F؇.6r]
��+����f��{I�MLF���K����d�Q��a��D`��K��1\�͂��O �4�zAL�	 �>�R��ݜ1�uJo��cy**z��\M��7���/rNDq�6�<^Ҷ��+
  ��E��4e�'�����Ō����b���9�,��b&|�j(Z���␒�ݾ�,aȰ�D�P��~��+�:AȽ��f�?Ӷ�(O-�H��:�� �C�@@v�g�3�p/�e�� #N�·W���3�%���(����V,�|��Ǝ����y�ɵf����,�z����i����nX�"�T@.�PgH}M�궔?�zk��y`8��);����9�ӆB�c�����Z�WIM���ݜ!�nY�-Y�tm�l���m�]� ��T�W��o�Y�$Z�X�g�[�6�k�k�f+���6�����eõ������)e�=�k�z�����\V�K�Ӝ|)���Ƕ>��Y(�R��,����շ�2cC?���?�:1�7&�f�^��<D߂=/n����	!�O�����:?7�jxN�4�w��Y$���an�)����ݭ����x1oKMx#8� kxl̼X�z���]CB��:��>+СXО�`L�J[��}I�Z=�7�tT��8�WS�ՊO5{��`.��\I��h��aZF]���9��4��Ð��i�$R�p�#J��Bֿl4�X:NY���D��F7��ǎ���"���N��.H5�c��=Jg��WI�!�$�"�v�NP�j�����U��Џ�W"�KE"mM!��ss���2�A�H��.]�ï��ر��8�;}�}j�kp�
 ���a;��ܗ".��(�-d:}��ʰ)4��M��� .^�%����O�c��a���m��30�Y��D7ED����j��B�_��8h�^����/���s�\4��㽓[��	�Ú��{�>����X�J ͹�x��ӥ/3���B��@dWʞ-M�B��ɶ/7\3��Zz(v��^�2�uЇ�`
�F��3�^�¾�qu�,B9۠1!���N�8�����ǐ��
TB�|����[��|���g`v@�.���
�PM5lK���<�|<��W�����%X,z�1��|Vb���6�̧�a���$��LNiy�8|�	�iDR���D	AǤ��+��R�t�GP`�]��2��MVxK��h���)�~�Y��+r>�jC������"���<@*������ۮ�D(I���s�G�a���S�8�\;�B2`�Ek��.��8�t��췓Nm��玻9���]/�sG$��l:�7��w �0���b��?S�R����quK���M�]g�o�=��!$H%��l8n���C	}��A:�~��7�NT��1�S��?	]J���2u��[4��[��A�+Qv3zA�\�~�0�e��ؐ���u�שmn�=���ϼ��g��B�5�<���ɕ����X��T��K=��՚
[b�����X�)r�=W��s� �����2w����Ok	��By��$}��LB�� ��o
i�ExD���~� �
�%��� >M���EQ���n��
�m��^?l��q�7~��P��X���
3�����ݪ���%r�La�l��)�M`���;���P��Zｭcψ��DEh��<���2q�Q�Y���$)3.�3��@�c���M ���������H�vm��%�:t�c,pcp��@@��.3���ߓ3 �F�sq�������M�e�p�e���x�����Z^����J	{u��tK^�Mq|?����/2����g0�r���:O�\��s>��/�`3�O4r��b�O.j[���R�p_�X��&nq�>3�_�<ّoG�Di}����zb{e���"D/�X�۞s]kă�7p��
��K�OCp.���I���-�h��g'�I�q��'��ek'��R���4�~�D�����1��f�������	jc-��g��P�x�p��Sa�cD��IYvv@�4�-D�H�Y��� ����'f�#t��Q�J۲f}���>l��8��W�/ΌT2[�;V8��ǘv�=�y.�ɳJŬ�5��]�/���[F�;^me
X$��:O�+iR�~y)�&~d�j �]+$�F'<wD���m�J(ߦD�i+E��m r�w��h�_�At���Q��&�kַ6���	�4�zE�q��>8(r���9Pϴ8��>vvBr�����"A3;Bi#�h�k?��Yէ(�"�x�����Ö-��w��T;M�jp�YP}�^�0Z�\��jC��,N�kYb0j2q)�7��I?����x��_��Gy_�ߏ|��ۗ��75����N�!�zi(-LZҦ����P@���^��N�q?Q�F�X���x+w��B\�h�^�t:�Hqv�޻C�Zd�s�� ;�;�p�����' p2Q���NA��[T+��r)�FrNe�-�+`������2vZ��KX�A��i�,s�"���\�dJ�7R�N�'�j�M��]�4��{�ѡ�5�yp�=��������5?��M�F�/�&�l�eZ���ħh�Ȭ�.Y�w)�R6�G����N�j���̾l���&3|y^�X�"o7KJ�P���t"�Q�-�5�ͳFd�^߫��\�5..哪碮�W笉��%���2��D(HS��3m^'}OV�lN���g���G�'ur˙��ֵ���nL�n�+��T)�3!hf�TEN��bS�ͬ��7�5��Q��	è[��=��� � ݾ�g�)��V��A<�t<:Y�Je�4���y� t�KC�ura�s}MǪWd�X�wPu'd�g�S�
��"�U�Ki)5k$R���ޖ��e�<��u~JJ�
��~��?�Vc��<x�Dtxf����a���E�10� ��O���ZShi��];ҫ6H�f�i7���ߠ88�P��v��C�����{hp�`0�m������D�`