��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�y�Sy�;��>��&�MA�)Cʌtg���e�8~�����=H�9����.k������U��U�Xe���M�b�(	
'�m��_�S,(
>ɢ&T^5�[Kم~�WA��Mb�c#�<˃#:}��6͕��F��O�j�7���'AF�9��'�ƹrq�9�p�
o�'�w=��v��("�|��ӏ�I�\.�V�����)���cB�չ6�t3sꀚ u?�({��_x�W������!�`�e�H�H���|�-�YY�
ꆞ �Ӟ냨��e���S�kFd�v�e����y�*D���G�>����+�ᩜu�f�x�I���*��/1\1����r�2�*M_�4j�t�'{)ȳ:�A��!���ש��6�D`��Js�[�a�O[�G�O.�����}�9�����E���;I҄0"}̙�������@pi?%D;�4=�6��`w�:���{����)T�y��ҕ�B��F"z/.��.�%�g}�|HW���c_QEխ7u�s�}?�ه��F|�����čg��ډ�+�!�aC���w�ŧ��A�M�ξ%�37m���x� ���3:9�@[fU\�Fz��Xh�����h�*Cy�i/�[J��H���Z�i�	���#�*�G.��և ��ֲ0��Q�s��9k�7MJ`���%k"��o�Y���Uu�}�G�2+f.�DU�Oī����I�
ٜr�1"Š`F)Wd_�? �Qi�]װ�'c�R���lƨ� a�� �ɯ�4����iҎ�E� do\5��3J��[�:VӦ������E$x�f@J��V|M�G�ql�:}��e��	k�Q����`� ^�Ea#��5&R� o��i�rY��C�n֮R��QM�'aq;8YfC���BR�Q<�?ēU�Z���f�c��7&#�Y��.����_�MX�H|���	�E�̹q]�	QR=�ßBPM�ҡ�+��+73 ��B�h��cP��D��qu�h���
zY�56	h3s�ތ"Š�ɗ� �x��^o�t�w�7F�91S��ɠ �0d��5bR��~���k�W}��ӫ�yx�����#�l?�,�}r�o�8{�B��Z�{���t�-��=}������jNܤ�ƹA���(͆�-9��jr���4�Ơ�^��\��>���/K�`U�x��~�9�ذ2�Zj,�d��,�<d���s���ꅾ�$�2m�������<:��n�ׇ6I� ����� \��)��j�9�%(k�� �6�F(�)�ƶ��d�^�a��ŻϮ�ɩ�ï���+kBU�/�Bl�!uxB_,�4� �4��ߐ9���r�K�	!��a}[&���ɬ<%��6�|[��"��ɖD��fp�<Q�	7ާc�*]ilMw"�&��S�D[���{/\�p�X3����]�~x�����f�(�8y�q ��z]�G��;�?f;����;�	:��
2R��a�ߕȳ�8��4n�?s.C$a<U�:�����P�ZUcl���GF����0QA���x'�3�
6���]��4��|�WT��ˠ�#�[I-�@.]�f��mc��}�vcW�<�-2&�:� x����{C�j+K�T���Fw���]�Z�&����/ҝ�x�>9B���%Γp�ety�G� ��~'+�4$�Y��Ux|:Ky��p�X���t�!`��~F�/UƧ+�3"�`��}�|jpz�!ؐ��4)�o�'5�%��PR-�{����H�v��E-K�М*�b#�~'�#��#v�(�b/����A�b�A��~:�É�~�)��+o3���h�v�3����,��Kh`t���E���KG�ϰ�X�Ƨ�&`$�@�Z��ٶ/��{q�G�xFO�K-4;�8o��� *�򂣗x}\P6�����K��^�$�o�R,X���k���-�k&��n�%t�J6�9�݀��ޭ�)Bpɰf�ۣb��|Q�ɐHCC��$}x��
$��R�Y��Gi�7�s��5�J���vES��--���7��M�!N�nX�h�W��(�ھ�&܆�`�P�Dm�<ѓ"?37��6W�Qj��$���Tl���g���^i �2�������^�ɫ�5�4@Pf4,Ǘ��g�-1:�Q�g
ߨu����<�T��l�l
�����L �$V��վ"���'E�S
�vĝZæ�B>�ȹz�%�?*�(�Y1�.V�d C���淪��?y�_\*���N��Q5U=`��+&MOg�3 èi����߈��7�@����XQ-�FY+�c�~rOS����a���F�X���A���g�2�P�ӆ���'P��y��
���3�ll��n�B���,yΥ�RFb`Ֆ�d�����b`�E�c�����<Ǘ������r��b�I+{�'"{����#9q�vUS�>��&�[kLT(������S�Ju��i�4<��$3�sdC�צ��}Q�Ǳ�g�<
I����a�6��kBp����(��6ăxx�ǧ���]�����f��q.ٌ���9��b��Q/&ҧ��0Ӎ\t�����#�MՃ�C�
6�E�� �{N I 3?~��I	�nl��y�"�����:�J�z� >���̑c�����V�s��$����;�&^`N
���=	J^�Kd%�{���s�~:s#�L)��-E�mF�/������x��^�xB˙��2�6Hr��x0+f�ڪ
ƀ�۝n.��:_^鰤����签�"��Yo����z�/�$ז2k��p(BF�)Q"�XW�~F<3~'33��0��GQi��I��G1� ���W���d�7������"��ƈ0�N��̌�<�v���#$7Й��p��#˾�nF�ߕ�I�+�D��i�G!l�D/���t�h�c��mQ� 
 Q�7�~�����l9O�
�Ĕ;lM���k��-i7�=�M��L������hH�����V�	U���l�|���v����A��$�Zz	4��o�0ԙ�팑�y�;:3���;.O��K�@�e�0��,?�A��)j��<�|D���4ゲu2�PTm�\m���h*x�H�E����ۡpR��-�,�1�E�C�N��.g��X��P?��KB)�����l��r��г�U��|~<�:��P+!��p�NY Nz�.�+���y`o�y�������F��{�|���`o:���`����;�%�\��MH�T}`��3�����yf2.��5|��i��R�)Gn#�P���#5.�r�0��!_,�~=��e4L��Dٺ��VBI�ו���c��"v���f���y2��8d��'�`Qu�_��K��Kҍ�������w��X�¹g��̢���p���{))u��?��0N1�a�.�����էE4�IX�)Y�Cnb��W��쟞7�!�(~;W�rI��e�+�����Fr�f΅j�z{�']{�%!a��k1�ԟ<��<5�x�#[��,�i�+��E�Y�C�=��iUlT��Vn6V���!��H���{���.<��i�� ��$MO*��
��W��a{�N:zGG���z�eI�)ｉ��6φGs�A	�,mW�`���N�IKdӴ��g0��J��Jk�%׭V�������ƴ�����
6��t�R�<a瞑n�bA�nneI��z�O�Ф�k�����u�::_�x�d�~�z_1�a��M�Q�Ϯ�*��M�(�w����MG��C�m�IŌ��@�5n�\��\Ҋ{�����[k��8�E�{���~/�~�'���\���Ɉ�p �?9|�
�^6��A��F�y�v��2ߘ��BU�|��8u'fڔ��0U�U���=� ���+�隞��vK�� oԙ|���w#z�F��t�˗?�2Ï[�$����g='�1�g��Yr���&!���tJ�mdح&��okdP��H���=��'>����m?�͝j�f�r��2���&�y�R8Q���S�����LpTٜ f�e�]Sx��9�'H�zt� �~��i�p��Ơs~R� ��Y�(ɔ��a��s5ԟ����7��S�P\�f�p2�Q��2���ڰ����uYQ�T�b2o)�-f�\�Z{$�b|�g���!����&���E�f��o�?�v�Lj�hI��j�[�O?�R;�� ����3���͉�4Q�^ϯ�]�稚�������> �IrT�3��jb�1R�Ѣ�P��ɾ~�`�u�Gu��*p"�d)sa3pa곋��� e4�VJ&���_�+����%�<M E1����Ֆ>�!�Z�]�wX��D�I:_�{�"Q��nHG���HȧO��ح�BTJ�j𜂐NَiO��@�0�%Rg�UC$��+'-bd�PT�`(���:y��<�w�2�����O*g6�t<6r�5�~����jyN��{_�G���0ra�d&�5��)�/n�᭟ =�VϢ":pBs�o�.1ۢ����-c���Π����u`���H���&|<p�S���"��݌��ɸ^V�I����h7��R���H�.�i��� {$�QT��;d��Ձ��6�GZ�����!+���;�+�s���5�'z`{�}?��s����O��H�E^��Ʉ~y����'f���W a��m��'�Z��[�y����"�0�N �=�܄��4  ��صz��tShk7�.�d	20o��_������+�m��]��{��D�8ٮ��^H�
�!�Q�I�*]6>(o��
fX���2F��j����BOۿ�Wvd
�A�T���������l�E��;�r>���q�8����a��@�8�os*�۪�P�w���7�,��c�tuff4~9����%�J�=�\�?<ܘ3gZ��<7R\�&���ڒ�v'{/�3m�sinWk���00���΅j�9Ժ��w�>�h{$�)L��ĹSܯ��	T�_ď��Yt��B�����6��%�a�r���Ri���.A�/�»����Ci{�������;��Ya��o����,�T�VG� S�B'y\��_O�Q�6���^o\��6�s�I	��%��]8�s4ʼ�%G���u&��vJ8���{�h�z������7�t��n J����Z+�h��?Dce7Xo?�@�k��+�,��r�ή�UC��IC�������� L�#ۼ�����}ƶE6���#�{=c�C�y_���mX�g�	��M&��ao�����G�%�J츌ʔ��l�Ь,�P5H��A�Z��n��\/9m��DyӎМN#�~v�%\���WU�e�[F b����hrڰ�����7�q��5�wGW^mr�D'̶X����IJj����i)t�t8���Ś^�w�{E�,`6ʰ��)�C�蝫`�G�-���=���k���go� c�Ȉ�0��dvd�8:0�n�("�@�o�f�T�GGA+`�r�y� �%6�M�_!}7��c"��M6ʘFX( 4Qc��u`r�5k֭,p	D*�y������L��O��t�QD=�_�V����b���s��t�sE+�����)�1���X0�q�׌��q����-*��|�6�P���*�Da�:�0���Wqitsq��v��=���/�K%���@i��ޝjF�uAjf�����'�=rp��T���_6���\�����;�E���:��l�)dr�H�7$+Gn�8`k@J��A�E����\�Y%[~��?xp�&mw��u�gII_�ldV��i��Y���K���{?��O��i�G��"��0d3�X9�#j˲ �щԵ�2ۨ�f;P�P�5j�f��fD���eK
q��eWd������bc1w��1�#rC9d�kC��aT�� O�-�Tz��;yd��7�NN3�"f&��3��N;6=����dږ/��0Sӧc������GX�x�Qh�ҵT�<�A�@��qЌ�B���Gd����3E���\��)�X�b�׶�l�y[��
|�6��.e���`m� '��������\U��W{o�W{X�6K&�eY	,��l59�4�����ǰ���ԣ�5�Z����d[}��-��8@�n�3;/BN5=���_�w���l�|��o��1���d�%�����׍Oh�r�6��;���u~q9�hw?�H;c9���	k�!��&b���M�֏*� ���I��(�J�|�ĺ<�7����`�hJA��I�ʨ�V�?��"8-0���G�zZ�"ŤB�Q�䷆lUz�f�} �{�~@[��G���������XK�ԋi�%Ɵ�}ݟ�j���H�"[���9���a�a;��ȰC�]�u��?�,��ݯ :�#���������e�E��TD��/�|B����u@��񁰑G9}����Y@����oF���p��&�S=���������{�_���/��	>��\��z&OO�����=������	-��H�A���{`J���)a�1�Cq�e���o8+��7���kԾ��1���b���g�Di���T�ݹ�S��w��4^����Nh
������*�-��[�L��RgW�i��Y=���˧�C2�HL�&����+ð�c��>���|�޸B܃ 5��*�d97JKb=��u��<�g��h̍r8s�pX��T����Y1������޲����g���w���&��!G܂}�6��|uW^��K���{��9$_*���H'��tKѬ����Uxd�Km�C�:Z,�=a�������|0��i	]������}��D��tT�����(	lo' �W�����{{�]��Pou�yx(mo.�t�1��']F�BğA��j�O4�z����`�� K��Ƒ�J����}n+g��L�5�?�7Hڂ����;�\^3�o{��셪��|rD����Ʌ>j�f�J�jJ���q�T@���@��|��|!3n��hҒR�*JE P����;�l�쑪��s��1���괻Q�=b(�=�j0���vi�Eb.dd�l�f�o}s�m�k��@I���J�AR�ڗ�0;�3���xS���A>"8||A��:����L(���Xk�T�j��Jia JLڠxe�NM8�wmB7=�?դ�T�k�Gn��� ��;�
g��w4"�8g�>6riV��S���'�8���r��b"�0��&V�y�!��T�d�W��a��8��@�J�K�[!�v,c�(���~"c˭6�
J[����r��=�"��x{u�
G��)��z�o�x� �����l�&�RO��y?�Dc��2�j��ѫf�c)��ܝz橧���xԿQ��lg>��QEݴU�Fn���~�q��KԀ�u�(��|XR���(����z̄���o9����C���pd�-���&φ~�m3zf���v"���%(�kI�F�6�9@��P�@�lvЯ͚`���JmIin /yq6]��@D�ѥw�XM,�=Ƥ�0�� ��x�϶����C�����SQ�QUsl$ �E$�[�+J,�TvN@C"�Ë�4�
d��#?��:���Øk�_��=��z��|t��Q3ɋO��G}�no*�ο��8 J�Q��ތГO��/:f%�/���-���X�q�Y�K��dYlt$m_�u�qdk.\������R�� �Ff�q^��b��4rvbs] ���؍k�H��w `ķ\��s{1�/g�|���h,$�54�e�GK�B��e���M������^E�eꐇ�[Ƒ���%<����{gޫb+}�h2�$	��y&��y�0 A1H�V� n���Z&M�2��ꁦ�q�K�1���̵�����Ň/	�67����K�a4٭Tځv61Y�	@�����5ݱ;�S�f6��ؤ����7`��w�d��PKxK�b�d�%缥�{HA`}L7���b���˜��r��J٘�9�㬡b��r�P�)�����l��If�b�