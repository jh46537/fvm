��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E��Ӫ�-N���=��_�@Q�:�7�����n�KyJPq��QIVC|w#�18������c
�X�e�n��8��Vgdz`*}��LW���$�s6�j�E�r�bǙ�����.A:�U<����Y���:�*��^#t�2�U��0��d�	�Y���W`�A�<���������(>s\�#W��Z���XgG�����p?��"#6E�Y�!��_��2���m�C�Ҭ�b��QD�;WG�ت�����8{U��x����b n�GX�E8,R�x��Q�ͼr�խ�y��9\���Th6�f��f&Pi/��:T͙m���^��,�+'Ծ�û���DO�����c�a8�A��G����/'%��5�����*A.X�s�y{E7n��qn��X0���� |����5���.���t:��y3ak�t���&���6��G=�g&o����	"4@�Y�^�{�:�ɡ�HM<���%u�}⨤�v���o�V$~BެWw��y��L��|�2#>�]�Zc�&3R��g��6�f#��uO��,��D��!IN\�Rީ�7�xf�^���{r;Q��sظ��X�t��fZ)�pjbL�3�>��?�7�ˣ��Df�ɴ�vyT�}*��Xك;�t���Y{����#����p����f��z9�����L���:ӤZ�����+q�t�e�)C�B"L�K~t�my�O���T ������.T��X"�_�7�P�V���l�	�A�I�Op�
k�L��{�	�n�N������[����G�FQ-��̕���}���"qN�1a"Px�N�n�{z��O��H>�3V��>�����WJm;2$x�AȱHE�u@v��!j��֬�4'm�S^OV��l���Gx��=��gH�[Rs륙&���|oG.�&ۉs,'fMR*�/���S���zO�eP��İ�l��|N�W��/�s�>n'��e��Խz�oӐK�����Q���1��c�r�5�c��*���7aRE�FZ�H�k-#�����d��(.EkP���_{�����F+</l�j
+aN4�a�]B(cAr� �|�a�~I�i>x<��w�r�[)%����+�n�n7�v�dy�3�l����0�'z.yy�Ң.�ʲ�菽�X9�-�Ba_��^�v���禍jW^Au���u�?�{��'�&с�Ó@�g"�F�W��HEO�
PM�!&>����m���� |��,��h9%�m*�O~�淔 #O��o�Y�m:�O�s������P̃�b�_�䱮�VS������=zOD���`��\_����8N��!�D���u�w���~0�Mm�>j�ݿD���{��INEAo�$��f�=�6'a�i��������:�bfE�9c����E��r9�?U�B�ܑ��[�痘:�~�+
�5}8n�"]9�Z���l�k��3��eDU�{{�y��J���M��\ 3�":��u���Nr[�EZ$[��L3�O�������o�/k���"-�g��'2?/VE_,�e
$�SUA� Dhy���[U����W�b�5�0F���5��g"��j@�z[�����eP