��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#���gXݤ����R�Z�.�7bY�C-R��1S?=��sO�w��p)��2N���Jz{�6"yU��wY�YwP���C1K��MH�}2�����*y�{�i����naC�Md��H���t�eJ����t�����Q*�^�~���W���QRSR@bG��>F3cj���E^:�{�<Z:S���-F��
Q�T�X`�3��p>0&T�#QLK����g�8����"��#%��dQ�!��_��X���ը��{��[��Z�߶CXXUg*��x�.��ɕ@��Fb�F(��o���*Y���^����/3��W�j�ˈ��漐���]�g�dg�\f��þi��kro�Y ��$�n�]QG�
ƯWΆ�����,�Q2��^?3n��2A?G]b����/���ΛOH/I+Z�4C8��7�рCN7E9�ڼn�!�%�wv���ݸ2g��y��i��_Ǚ,�+~8[P9E�@��D\� �D�t�u�|u�C�����Б�]����S���)3�>uZΧ:È�Z����LC��
Rb�s/�yfi�a	���N��Ŕ�>�; $�2e:�m1Z��0�U�����M�����ʇ����z�=?-ڀ[*n�$,O���d�z^��'M���U��� �NK����0�gf Vn�\�ڳD�����BOP1�X5����y��Ɨ�gT��Hс�nK$<�OUB�0����X?�����F���~ˡ�Z���(�A�
TS/Š@'���u���2�F�:�'����1��J�	T�|~�N�"B��� ��S�&cVR�+��6F'�}�r����ئ�\�oڼ�Qq�2���]��E>s�E_R���4��-��ۊ��ѥ;O|���1��� �i�������?,���|��X��H���x�2�^yF���߀�f�4�L��IuHK��`	�����s~�c��}�'-"Լ���� ��Ƴ<rwG31��mE����[�T+����e�\3�~0�->�`m��K��_L/�DBQ�����@�]!����� ��^����Q8Y�ԃ:���d��bp�/��ճB��}bA���2��*��N��r��,>��S�!3��<�����?VM+c�F�&�	�J���������Ĵ��H�Q{�1�*(�V��2YU��C$�D
�-|8[��"y
��6ɻ��hC�3��-AR� �33�^�Cb�xq������� �~Z���f8P���!Y�傦Zw�*q��M���&Rı����!(��"<�3��ߚe�ü?��X\�U}M�9��`���8�ϋa���!�.��1����B��.��ܤ+NKW�m^�U��:��['!x�[�ޔ�zy����`|��Ⱦ@[_5��|K���{$j=w���˚W%�>6�֩Yu���䍃Wf�� �O�^�Xs��՝���%��r��0Q��d�[���&rMZ��紫G'�.�*�_l��?��#����fIy���#��'b�&�ҡ~�S�P�S��Vc�p����
gk�4�ۀ�8��N����p�򸗖5Ytӣ�8&{lmU��8�����W�'a.�C��*H��)��]�Χ*C;�z<�;Ef������;���m�G"͢��3@*N�rw�{(�$��m��In�Y?�MDdkK�ߤ�hw**D�)P�9�CZ�zd�E���q.&�/�΀��(s���2҃I�#�>�@=�k=v|�Z�괯rκC��$���r���c����Y`��l��T�5U"ÐS��4{�LMo|��++��:��*H��+��3�����Xr�k����$���<�}�_b�[7z��ܔ&�t�`��NKn��5WQ<$M�\�p��]���ՖLR�M�C�Z܆B9�Ò�z�|3
��UU0)'*���+��̏��`������2⏊x}�m��+h����
?[
mvwM�7���Qx{y{��m�e�Ru/�]�}�0��OS�N`�H��(�@�Y�?��5:�kX��+~[�+������ۀ^R�f��M�zM�����{Z-��*� ��2&��6}�W�Z��5X׸�~~8h��p�e�	�Eiɗ0P6�*j���n�$N�l���nd�͛Q펓�ؽ˃�:}�L#�h�j��&�t���~5<������������z�hX���`%"Znه��6��n����h~ޮЌ{�8Ӱ��C��7�C�lw�=��K�n���G�7�$l����C�^= J~o���.��}����h��v�D�W���!U�y�)�V���v�kl�nD�ddW�^��-s��R~C�}Ӏ�Ɉ'���yi�!ş��X3���K���F�,*Eu�Q]����ЏUja��A��K��J${(]?շ�c]ݿ�6�劙sg��6�" ƽZ�]�k���&���L�\߱��fܮ�p�Pb^���v���"J���Gtx�y<=����L9U���l3�tV��7K�������3Ӧ�TAok�j�]��ސHZ^�ҦY)!��椘��fzOږ~������>[r���K������y���T_��`����l?���y��js��
:��JD؏���Q]>�_IY{�ʧ=�IdY���B�YY���h��^Y_.�&0s����_��$�s�n�}��N���5b��S+��pv�D�U��*i���s<��,�ԛMn@T�IF���EwK8��^T��8���k�z�Ve�����C�L�b1ˁC�1/���-�D��"(�9�_�n,K���u���!��q��ѳ��2�@]C����9��ŗ��9Y�'j�"㯈	�AA�=��W�qrT���S�y�.)א�=-�*uk-t&q�,�B	<&b�3���^0�6~�g�[mJ�����y/�(I�:��ݭ��Lj�ICZ���flA�����S{�k�F������Y ɺ-R|k]��^��Ϧn
�-�K�(��/��#W�!p�=��kʜv��Xq�����e�w!��O��u��ZՐ}Jj^�v��9���o��@0_!c:��$��~��-�j�M�A�x�0i���| 2t��2�.kޮ��X�3���ج�7�R��v��#�ޡE]�=e{a�v�r[e�r�m�y�T���
a�V��|�#~��״�ns�+C�:jB�؄r��)~�9��S{��8�)�,DTFu`�f �	J��9������\��E�	<��OZ`�U?���LU�+����n�����)��R�G�h�L�Y� ;���`��_S�T��N;�q>�a��q �Ȥ=�,��_�r�����+���_� �x����K�=�/~&��L�T[͸�/�4wEr�)=��M�ͬU���ͻT���1�24˸5��Dh�M������5b7i�� ��o�0��v�����jT���UhB�P��/�T��&ފ|�X��]	�Gk���xG�!�����b�w��FW�Э��8S:������L���0�g)�H�P7��ҢGf�v�+��X,������(�T���픾yO�-βj�Z�tC���.��HЋ�|�-J��3��HɚmZc��3)�,�űā�G�L`y�-�e��樬)�ِ3���G,g�k�>�=�.��s|2�D4,�a����B"�[�W�)�4����舘�`u�˜��<K\�u�*M-���2�5?	"*��n,X����f5t8�j�C��	㳜��.Ľ�<�jm^F���� �4�yvS�V)b`�{�.eP�g�Vn������K@p����ϼ�~ܛs����~LEk��!���^��6�H7
�{@qE��aԝ�yr����=K�
�p�:]&~�G�b8��'��5�$������au"�)�	@ЊVTJ	_�2�ʣ��0�З	�+ܔ)�.�V�so?���XI���`��p@z��>ڲ�	��cQ��߃C�y��*���{�¯�f<���\wR�E���I順A�A
,:�l��P ��xX��a�����MA�aw�^��ژ8P�b�� )~���9a�}f��Bl��V2��ǹ�Ntb�f�ȍ�_�sB�-�J�F�%�\�fL�F������U�?d��2�������r�z��,P��]fT�pmL$FP��͟�o�@��u�����yI�^���+c��k���_�J(�Q�4�|��1$bh�{x�b����j<vQ����l��@�<9!6��Uq�k���J<��[�|v�����di�h#)��k0{�(��D �Y����{o�e�q�q|Fa�4%��}���j���R�X#6:8_����$+G:��!��[��X��5}gD�lbqLy`t�|��%Ͽ�����ľ�a��#�CoN�\%��c0�]ƿ-����h�<F]�K�K��?eC� �n�����Tك��5̄RVl幰�a��`4��}����p(����s���:	���iK�e?2Rka������<�xCڏj5#!�9���X(4
�n>�u�X�x{xFA�,D����l �.��|?�&�{��M#�6i1�U��Vv��W��MW̶
7����[#��q?Ҿ˰q�z�"�9�=g'IQO�v��b8eP�j\O�q+P�c�WyJ`'��#��&EVMw����a������ꄯL9���Z��ghB��B�������V��� �9��o��6����O����O)J���0�����"O��\Qܔ����fP�|�ӫJ���z�ʆ��gi�{��/�!K��!	���Hy��bG'�g�H v�<�+y�p;�l� �)�u)���Gp�e<T�?�#�Z9h����h�q���W1|�.�{k�L�8cO!k2�
ѩ]������a���Gc*�{կ�(��w����d��X�]wTYDK
v�x4�_t6�t���v�<�N�q��x���X�E>����M1����0`F��sk��n�d����4���i��@3rE9c�I�I�&����ͯy{eX�y%��&�o ��%��k�nD�lп/~"IՎ��ڊЃ����*��%V/�hr��k�=q�p�L��p3]�M>@��ڊ�.���E��Qr0x���98���Ǐ�$�5_+B�*�;�1p{�l��k�����E*�Д���c�V�Qe.��]Q_�#����C�HY�`4=�n:���-��*�3$�n�Hh���~�·q�p�|�u}��0�t�ʳ��wS	_����3%�A҃랖��Z9��2��t��n��y�v"�]���h�����1Ϸ�:��	��nL#�?.D�s�Pg��;M����ś��vHG��
��z�բZW�U��C�|y�=\
8'�L�1�^kv[�H��%��U(�u�qM�~�J�W��HfvF*�S	��1��Tw��K���`�q3�6Bp�V���۹f�� r߉T8�M��^'��e�/����|vP�n_7�UΥ�^�k8��z(��8U��7l�,!�4�ap�l^�Zt��q�]#��s�����P��Q�5�A'�F5@MF �Dh�8�$/�y�f[3��5R�;d�hT�}|j��Zz����}�O�\��dsp�[E�-ݼ��O�^����|�=�n��C�����L�%��+
��ڟ�Y��Yp`�%F&���O�S�o��	W������~�l������Z���%f���N������)
�4g%9�\��O�ˁj:�,�0}����XW<|}tV��m��MHi@XN�����$��ϥ���G&`]��!�����l�k0�J���c(���p�����}�oR�qB�3�/�N��X�� �{�O����S\Uɘ���#\t�V(TB6�r�g
HT������S.�%j�%����:�&-(C��XL�W=�w�nU����cW���A���r_����eu*�C�m?K"d�g$�j�G�k�t�pA�������=�w+B�jq��WSGH���f7��$��|>(֏��w�|�����V��х_�&������J$�\4�L�\�]�A�T�̄2(߿��H�7��'.d��w���|X6�oG��K��,�ֲ�l�)d���Q���`�b.۾dE����N�XvXR�{�b��t+�������M���$@�pL���ɏ�A�O� �Jѝ-N4��(4Y�@����ű���1�
��d��N���|aӨ���ӄ�mճhQ�)�T@�v���ESGb�7M~�e�};'���k0њ��I�C'�Ac�d0&Ne�xo���I#Pq� �}4����(���+-rx�*E���+����PO��(ҝ �L�Pt�.}�aklg@mL�Q_����@�����WZ'G?�>-XIዉDw����`��V��� ��#�f�+�~`����[Ι�-�>s4F4�H	]�V��'�aD����:1��^�T�����z�.�|�`}�����C�m�K���i�F���{��@���s�_��!6lRS��q�� �j���7�{��CF�~e��ʶv���/IZ��5$!�ޭ?_�#��J�9��~{��)�� ٚl��wbށ�����S��Kb����@5!�;����F:�!���"u����S��M���6GF�/�H3�;�і1>�X��2d�4�܆�T4h�V�H�7�ǿ�ӟi���CZ���v��
ٚ��/.J�c"J�L�}���J�� d�}�h�S[��3!#��8i�%��z6����t$�W���}��_��.-��=4��4�}��c�����+���u&��wvc<e����Τ�������w��t���%hY�>a�_W%�k�)jʹ�e�Tk"����T=�k�<0Iql�s��东~�zM�lZ�j8Yhj�p����A��N-���W�j٥t~��)���U�|��6�����%yW�ę�߂~��Ro
�Q���">�Q�d�$s��8O��B)����P
�s�VQSD**�6�#��!�ao�P���f�G�0�ι�T�i�,\&ߘTA���#,��(%n�q���g�5�j���4f>�3g���u#Ca뙖3Q(�-o�U8|�Lo�����&�{��Q�.8�����v]p�'׸ȱtD=��zo�ӭ���/��m��"J0����ejgt֫�������L���I��_<���}��[[Ί�l��fT�8��w�G-��C��p�}���u;���V���kF�#}�;j���D�]�2l�߀�nw2e]t�x[�O�uUj��q{�ǩ����F�7d9�5�E�+ђv}�`�@풝�(I��%���Ǆ�-�U��'�urp��o ���Pa��ԗ�ҿ����Hh���Jv�<�i�)4�h�+�"'B��p�g��?����L:~q7Q��j�:��i�מ���j����szx���=��[�|��)ep�;����b�:�4-(���.iȌ�{���D��y���߷8x8����u�6�!P'��ҡ��x
�i�z�K�yz��!"�Tj�Z�4��>K�e$��U�3�X0�~��U����Z K��vykV!�9��t�[kֹz�=�
:j��ԒBl뢉4*)h����4QNl���7��yA�l|����}�Vte�u�f H�g�p�M��P�o�_�4; �%��5N����y:���T�䭌?u�z8>����
8=	�0.��8R�����(�4)3�#(����B&oE�Cc��h���������Z~A��i����-���@�<��;���	#�_ɒlkj��O�!���3�qcp�EF���X��~�lAU���d�hZ���s6�cL�Y�Q����@iR����cWA���˨����g�T���J^��9߉e.@/��6P�(��|��y�[�/������qp�+u"��o�f��I�$�G`��g�tB?�&zTP �sZz�zi-t�燎��# /q$�Dm��ޅ��q�i���^�3����W��EȒ���FKn�:X��$��C��A�����Oۇ��qTwN��5۵�?�'�(Õe�':R�f�qOf[.XDX�����Q�\�V���o��TH��1!�L�8�nqc�!w���Z�9�\�&D%|�&��-�/召�S�F5�GL�4�]�����)0"J���j�Xg���������U3q��0I�����I�Re�C�G"7��Vqv�>��0��3%;������S�L����,��T���ӝ"�GSy��w1c����y�z�]7-=�I�(�'<�=ְ�9|#й���Y�z����8M�sJ�C�k� ��T@h�X+�q��~����msqz����g��wTr��iu�L�nY��FDֽa��9ճ'G���y��Ch�=�ϝS�v�Tÿ�1+B �33K5qhۇSp�P����S=Z�G��ku��5͟��G�t����vZ��-��D�w��f��]��U�ι�$q�9W�q���?�N ���.)����b]��t�9��E�pY�.�<����I��4�K�a�MH/���dO� �#�QT$s��2��e�P���׼U���T�L�I�AB���{���.d�-�����8����e�-�X8%�p��/��9{߬L<�M����)�p6Ek�fcg
)دH�x��p�2�l+�Rա/��� �ˬW(�\�2�|�ΰ��V�g���b��Aߢ��ş���\y1��$�9->m��g~�5>�P���&V�' d*>�r��P��~��'�w-["&ܤ�Yb<z��f<�g�Ez)���Y��A.�S�� ���ќ9��k����ճ��p�!>b������c5׮Ґ�X�A7Q�Wu(�^YW��e� (v�@���oh/�D������ܽ�Y��!�̙c�h��⦣(��6Y�|?��	�#[���8>~\U�#�w��+��.Ʃ��Qj�(mm�1�5}�.��`ő&mI�p��B�Vh�c8�*��ils��+�׊�Xکt���ې�Z2���d{��=B]���[�Ѕ�&�+-���	��ݎ�~��Ys<��$@"���4$�U��Aĕ� .AJ(B,[� l�5��*'�xv[��ߏ1m:�R8�ƼP�m�״iY���S�3`�iʍ��jJ
B|��5�n�Ax�AI	�lA���_���3Ž^�3��DR�T�v�������LV
�G]�th�tj��3��NX�%F�S}kc���c��1�"�=��nife�)ڐ��X��R�]M	��4�"�-HzM�uT<,)T��_A�}�t���}���sB��=�*|�P�>�t[���O�\����$���;�"�����h�OMv�vMI���/���;����'�0�AZCvC��F[,y!Gw����(To!�w�@�+�SLct1�=f������n���L �34���g��#��'"#p�y��cϋ��vH���nӃx?GGPO%n)	�O�<�L��$�X��	]�/s��x��h��;/a�Z>;Zs�7֍�!�_�3�m���x_%Y�G3>%}�H��S2�G+6�x��t���н�PE�͕�e���h��ֶ �!�b�-����T�I}��U٣[�f�������{	��RS�O�Ll?S���&QM!o���r��7��S��OX"�UBIS�'�����=���h'~�G���:�� ��jg��=�b��lKB��L�G���T\qqF�f{�%�����ה�ް	${v�5��K���.��xɇ+�o��K��N"�yo�pΔ��Z�@�/;����T�
ڮW��1�PF�S;�d�$ �}-E9���P8C�a�w�=������T�bS$���	Q��ɚ��.; Ss��Yi��qcu��\��6��&g�d�|�W��ja(�,X��"Q\�S!���<Jx�	��
o��r�Ȥʊ�!����@������U���0�t���C^BR�����U�Ig�!�˽�[�kBuyE�t*@�܄�[��Ј��	���](Y�3���{w\Ny��H^�t�}��B5sF��Q���g��x�q�Iu Q����~)ξ�Z�PU�4���P���V�W�n�5*?���A.�3w�E)���[QȀEx3rK�'�hX�߆��qK�8�1���, �]��|�4��w�%����F����_���p�m�1E�_�~O��Zz�}��v�\�F�?�9�e8*�{hf�����B�8�͜ ie!���ӮyJp+q`^�7"��[�����#�F�R���2�Y�X�HZ(�!�~���T����Dy�l)�;˝��@���m:5�vk�1�[v� ���x8#��i^�p�$�� �p�b���Wl!xB������Qt���^�E���z7�㩩���9������X�\�� �S�m#���tz{�"�`��q�� ���-���a�����2�Ab��0�0����f�O�|9c�f�~B�4`:D�(H�>+��u!hU�~;�~����z8K��}��V>��U�8��@�1�Q}Ie���p�懷�|�Xj�;���1�Q\��̬?r�o���/D�{������t�8��{���Gy� ����'��d��UD�Y��6<e��]�W�O�]�z����[�@��#��T��Z��o瑗G��-�����ŠK�E��؃"fFg�k��?yۥwפ5�+T�xw��
Z��`f�p�v�nn�?'a����9nc�4!q��!f<l}k��L���|�W����m�p�bL�2�2�����΍��͝�e�������7����(�VK��W��n�L��@I�g��OϿ{� �<O�.tb�ʽ(8��$�=����	�!+�k^1ϣF�~�}����S-�������6�`�:�����.P��[�r��|�8@N�=�)�Q��#,â҃�K�93�I����"Iqqa����T���fwMm`�J��$a�D�*����o��_;�[&ˏ}U���E#���~���,�>������RE"�ø��M��\�@V�|_�#�&����q�
݈F�I�$8%$�K�/��ᴕ�y���B�D|�N:������`D�)�-kzjD��=�H�Dʼz$�BZ���/7�i��ڞ�X�D��ms�|8�=|kت��:��4��R�,V.��/nHb�`U%�Z�w1�O�zBcdx�3\��~���j��uŜ�|�o7�[+���I��u��F�� ]���1� ���^#�YnA��I^����b�YcA�7�^�)|�����`7n����2���0� ��z�C|9S,�Ń�n:zxp�������2��\�~�E#��_e�TIY�i���t��H�܊�i�V�m��p�����)8ux_riL}]���V�t�8���J� ){�y.$>W\�|�Yf��O���??�Ԁ���TԔA���z����X�;����,�!�}��z�)��BɘA'B�� ��~�����1�	�����d�0�����hwT��j+]��9 �}p|-�-�M��ڙH3�Te+Lg�S�ېR����pЖW�0�y���_�^_l j��R�A>,n�y���YaS�|~ Cȅ-7z��`m���>�*��N�/&%��I����)2�L��1�����TY2M9t�OՂ�C1y��/�T)��qM3�\T��ya��
���I����'�rœ�H	�9�N �*�
�l{�-�M�5�Xj�m�����5+�+�O�����(�"l�h���d]����YT�����K���9�R�{����R�ʚ�hNc�c�Ӧ���&B4�JT�J��4�� ��єS��5��m�,y/dQ�����R��xvH�Eg�V�Z�f��!R�uv=}��P�tnYI����A�#���6rD��++��F<��G��&`Yϡ�A��uT�Ї�=���	%0Q6��؈�6?�
�� �t����Ք�'��#W��Jd�],Cw�Y�l�ZU����;Ţ�<bD�P�
5��oys���-.���y8���%�����o��_�\u*,	�N5���k�����'ǘ��f�E3�\����.W�~c=џˎ�	�us �J��E�f���=��О�A��	s�v�����0z�a���=P��+<����``,m��=,����Ĥ满�5��3/O�����q�:O;oeoE@#ܝ3�9��56X	n��v�2�@�j���t*u�3�z�z�P�*��̈C�$�Ǻ}������O��EV��@�T��%��d�2��%M��Ƙk����!�-[�EK�/{]��W+�붟n�F�
�W����{�l��4>���C���櫘��$Aa�~a���X���hB^`��V
{�3����M$[洩m_Q��w`�ͬےtS��M"ç�9�Rk.+
P��W����}�W����nuI�jkT�!�h�+�����W�#e9�x�d���L���Z��)�GǴ+���cdե]��H��V�\�qֈ��y悥f��j�z����VG��_��r�*��F��p�Ǆ\ջ%��&�>�"K["�0K���L(T3��=�a��� c�V`V%�q�3�E��&d���$�,�$-��T0'j%��E:�>�W��s�'-W$�ϸ.�w��1_g?�K��9n���6�y_'1�\h�3���{(��K׹��&��mt5�B����������
/ ��*7���e�����_��E��a�J}�@�J�f�