��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbT�L�!�4��~u!�:��0�� T�^d�V�0��Z��������7n�+�qB�$�)-����f��p��p���'��?�������������g��
CZ�·����;��7�eRp���ɘ������'������1s�1��[mR}��3E��rP�l+*���K�� �зM�9�4���!Y&���u��85�7iG��C��q0'UƴE�+۫�v�԰�O� !�,�n��	���+�(o~�q�� ��cR	F�A�cD��Z�*��p[_��-NF���V������o���	�>+��Ѯ��i#�'�|���8}���L�xV�)rl��>�Ѫ��$� �de09�D8H����
��f(gd_�\`"�
Y��H�t�L*���vE�	>z#A�BU���V4��KV��Y�;�V��A�j$�/:P�7k�����Y���ҥ�>�H	���̨�����Y.��b�N�]7��˻���o�u-�d�1�1���忳�'
v2C7�R�l��VQɼ�=BQ��&|q��B࢈��E���<r��f�'\w��B���'���t5�^n��ac��v� ��*T_FE�NIY��9��.}yǽ�_B��i�U�u~�Ӓ=`�yZ!d��yߚ��2;����O��i}P7L�����R�}k���i��m0=<�G�|�����g��
��$�Pڏ`g ��u�<�ƴ�� �~t��i~��{D�����6EB��2��Ԓ0X�
�1Zl�֥������6�b":�h�Cs5��`��M����CRk$�'B�fU\�(�	G���i<�۩>rAm�J�K}����֝\�n�/����aA�w���3(Hd�g��{`kL"�� Ȃ7��-:nJ=�<A��� ���Gcq�3s	 :�������e7�T�kQ=���O��z����[}zUVG8?���&p���eQT|<�#.c!~�����Kճ����1m�rW�}��^ֺ��.���^T��|������녘Z3 �@h>
�9��ex�(/7t�\�t2'(E"�ɵ����>��9 �qЀ�X@���]1D^�V˱)X�đت�\��D�����ʳ��э'�2��A��W���H�S��ӟ���7��Vَp�;�)pP��Ƕ �[q��"��#8	a�+�Y����[�>�N��WY>�,�[T�/��|�q�nM�z�l�#u}2�� *{�u 2ϒiCά~����r��r�q�R�c]���EO��D`Aw(���^1��:�W�%"m!�w�[
3M|Kys���-�7�wf���|��{�Ú͡# ���}����-kG���!\sb2����>�^y�eIĲK	���%kN�3�x��l�Q��a��Z���ൾ���B��)k����)�=e�˅�.��Ei�_�9�n�/�(�r�^UX�zlz��ܢb���ez�#1��L�;��?��B��j�w��`.���Y��8�eL����F:��`K������8�g�!|�J }|�DU/TI��$3�K0���ɒ;����_�丰~<u>���^y���W��K
z�&P��L�t�:�NUb^�KX���z��ܰ0���";g,�����*݈�W�y<��J��_LTF~<K�" ��azV}C����c*!4���:x���<&!��Jm{�$�,ҝK�3?�$�;����f���[�l4-'M*%�?���c p�w��EdNI�Jz�s�vh0�Q���͉?D�'��#=�.@���bq�؋af� �#˒�1e�I�"�|{r�q�|���7���5�R<��$�>��c�U:�u���U�[E�W�ʳ~��X5��U�	3
�vs�zf�taX�"1q�ʙ;+�P�/��d�3MNJ�!�����Ub>#��t2G.tݳLA��4K	�s�f~u�Dy�����K�ؠ�4J�^�'�u]��}�>,Csڥ���g�Ȑ nΡ8	�nH�Wi{��)�_�(�C�@��R��wO!+q�^	h0�N�����@�H� �p�����z��(itZz�w�D���r�g�=~js�`�@��M�Ǐ[X+<l�Q*n?w���`����:��B	��6����["d�u�>���Ew����=��3��x|?܎��7B{�Ts�s�iN:��O���E�t2bŏGdAL!ʱZ���S�X���#v ��vo5�����mq���݄�J�����F��Z� l:ր�D|�'iw�I���du�X��	��*��2���e�l�����4Ȍ��eF��p�U�0���i-�磝����F^ ���oz����/��qo� �b���o�;��SlQY/�y��(�@)���,��3��6�����dH��K5"��8�2VZ�g;Lw�&^�[��+�Q~�t��:��:37j;�h ^X]$�L���.R�HG�Gf%W��S;�.�WK�]����C:��d�1]��[�`���vn�PP�� �'9�+k��|�L�3��>�����W��	÷��d���5s|����2���IrC�Y�����,U,��o�5om����8Q���՘�g�f�,�tN�Q6C�N�w��`��,�7V��iw�QR��2�k�r�4�t6ӵ��w^ڋ`4.H�5�^B����ޡ
ZA��E�1}q����s�xfH�;��W��v<�����vgǼ���#�B�.����B�󵇼^�x¹k��9R����OJ4B�Uj����4R���+��5\\�:��u2��j�Qh�<�^�K�=yn�H�����ܥ�^~fr؎�std�󚵚�hH��%D� �ks���:�Ok�X�]��%_�/X�2�ɲ��O�;yc���mK&��$��1D�Q���Y��*F��������/�!�]����eôYs���E������y�\��� �R�c�� P�V�9��5��}���C4t���_�S�R��j\LFeNE��(��%D �qQx�C�S�W����Fbl��j^O~��r|`������&+L �O9�'�d�o�w�{j�Y�{�w�!����u���O�t�����!��DI�פ{xi�tm��Ua2:�.N-c2�ih��֗�A�i���J��p��Ć��{�`�6K�l[�.�c��ee��
��蒹E${?�
Kr�����{5~�,yP����K/rt�d���ydqS?X[h�	��2���_N�E�?�ȃ!�EDy�*1	�\{��7#��w�G����ڞ�;�`�!t�Ϩ���Z���$�V�=��Z�y7(�m�ɞ�V]$SH�4���M�m�W�|7�|6�Ǚ�,��rw�)~�!�.���g�s0�*o擄��[�����A�7���o�W���CH&����B�N{���\ά��PN�\`P��#�rk�:�hp�}��%���ߒ�u�; p'��Tv���Ȭ10�8W�I3g�!e�~l��ԃ��U^��S��m�@�f(7C�c��2�o?%sV����o�)@I�X�QէiUc}l7��-���ި$����tT���G��
Z�@S�<�P��'K+����ʭ-��c��|�hs�hk�p>'���Kd�������Nc:<����W�p�Y��XŎ�,���&�:Sԣ.s	㎊mW�U��+�\	)4�=d�����I�w�c�~�k>-u��H|Ju��z ga�ပ�N�V�G�z��@)�T(]4���䨌���x7� ^Z��x b-h�Y���4Ʌ'��K������1z����Ю:viQSqPm�7�s�_]�ူ
����d.��{sO!�{�@�޳t��Ʉ�/׆�����8�omPܾ����{�!"WC�$w�#�\���t�|��鮃~�2WR������צ���׌�,��N�;U�W�.У�E� j�)%��s��D��ȳ~�����H+��X�QG9<��}QR���!��/�p�����iq���>(�+�29['������w�C�It.)�~�?�aN[�d�K�-��
��m�;����[��V�JD$;��g�����F	���s�~����ˣ�@a�, ��4L���[�Ѫ��d��QB�-tKP�#�)��<�9;q	/z�(�S7�}5JYC3�|h�g��/�f2���"KeF�AMn�!<����"*%ȳS�-Ka�r��S!hfǄ������ǚ�-�� ���=��.Ш��y]cb���3�/�,��%��WQ��m�=�k���z:W&a���y��0������?fJ�j0����PT��mؒ�d �9t�G�<ư_q ���ɖ�W���< ��$��:�p�DC�&�Eߟd��H/�����O�[�4��"ڤ�K�_VD��D�7�|?��c�A[S?��p�+�t+ߵ�*^�b���U
��A���{+T�#���9rI�eP9,��~UUv�E���7����z�x��U.�eqA��M2O'��x�F�r@u���T��c��.K�_��_�/�|�4�T�X��)�T����%���uYy��0`ԏ�Tѫ�T��Z=\���Kz+]ɮ-��n4�M�ۗ�j�-����)�D�Xb�t[5�{nі]�
�:����������^o1/"�wU�2����K��0��m/FSS(/��Q��[D�Z�t����*�����>�d㯬�T"P�LZ��:Φ�z���\۪@I�
�Xf�RU��늤-��G�����
.�1�"�@�TA�	�Jz��g���G��&)���-���S�t�y�Xj2��|�a�;:0�����h�CM�_���W��$��S �d3��U-��TUb��'g����(p�o�1��ح���Cb�"^������\�
\��m]d��g��X���~� a56)~��O�:q�����0��g���-�o��i��<�98�#ֽ)�z7Ή �by���gsi��&�&� +�N�,t����qـ�����O׌����`r{Ga	����1���"�#���#.e��lo�N1�N
�lD�Ea�J7�$[/���p�H�PD��wt�+�Z��G�d�qR�\3��Y>��\�j�L}T�fRߚ6����`�)�KK[�HG��j�	�>Ɨi�Da�-^3�^��r8�|AA��> �qѪ�h7T�D:Fb�}�Ad��&"Ϩ> ���qC�S�p��A��_�xG:�M����Iן�?Q����z�c5�A�Wœ��fS�s`���;<��a�����4N�?��������gv�,�[��٢�p>�sWᯤ
l~"�+t���%W~$4<S_���W{�Xq'��}kM�n�ε9uZ�O0���:�O	ߌ3�`�V����ʚ���ߕ��9����X���.��p����1 k��4\��x�/��ԄepuZΘ4�0��{�es������+5�*��	�)�� �_�Z�JY2��(�]0��k�We\�@RC�rQ`ú(	:�Xn���Y
Y�G�cZa5��v�:���������G���-�(^���� l�?WFuwf���N�|j+�C�={��Ϛ�<$'p��x�b@���5[�b�K�Z��-����Y�M�d+��y��D>�4�� %l.���.�6���oҫmM�x:H0ss�R�d���XWvC���X�V�W�2!����=��i��&,�N+����3-O��^z�j�Ȁ|�j�	dQ&K��A�f���4Oc��*�)X0�Pܒ<����i'�l�g/�=��p��:б-	�k'۹ใP[�h��&5x��<3�����j��N�����>�洑�o�z�~���V��:SJ��Q�,�}+�kU��c6�
AY�ŭ0m�<��0K�t����k!�䰱��H��ɚ��'S�}�h��)� �0����T�^���5�>� 6y��K��v5K��)N���q����S�T�6����?"�5#bB�>�JMW���tӳ$�P �5�� y�}���{J�H?��cY!|]��e�0*b*
�g֠��[��FF[&w�f��I��� ��V�;����.�B�U�
��A�W���$�r��+l
iNΖ�Ǎ�G�f�Q674�j��1
�!���{U�S�	w_�OW�hp�/~�T�)������Sو����iV��"��V��W]`xS�!:5�f;tuX
�cɋ|�&DC����l.��N��	����|hc���#Z�"̣�6���Z��X��v7�`��@��7��H�e�>�^��$'D��P��h���;{U�m�A���,A�����\�5�&�x���f�6�)����ϰ&g�Ò��K����G��ׅ*	,�(���J@%خӿR�(.�\�UӨ5�0��[ОZ<�uVO��+�r$�e�9�D��ˠ���BV5(�����߸��L�����ò�h�U� %�" "�z��F6b�A�dSp
䬝��l�P����P�#�oհ]G�Z@�b^��c?.ӒN2��?YhsG^�D�x����u���JND���6�_��ȅg;�'$�RQ�*n�+��q@��4����������oO��d�3
�����w��/��#wI'=����+����q�HH��� ܛ�����]2�M��w��2zWI���7�����5��[)&�֜U�O��!+�q���	���0T�����K]H-���K��w0�5�<A���m0	px?N= ��P�M\�J%��hg�����^�'s�e��Y��2�{�����p�d�܁�'��� p}�y���f)�0 &2e�dġ΄+�c��W�b�ǣ	�d>��Pv�l��^����{+��ʚ-��]51�x4��޸,Q t�|��6�A��
��Ai��|�(Hf�(E"��0Q�������|~�(����l;�2�Z,���F '��Ǟ˒ԬwP��}�������ɲ�<�(6 �v��Fq���:�/�=)beJ����n���:=+k�*��=�ӂ����0Tu�k`)/�`?@��s'#]�����2-Z�5���e�==�㱟B��E̄4�x^��� vX_���o(���A��q �9!��]V	�\m�ն\kZ|��9���Y.�R�C�~���,My��$-�K�w
�h1���O������1�?ꗠ�:���0����:Bp��aw�����H��T�$ߠ�R"���G�&L?�6\���u�YpD�*3�x�C�]�R�lU8�5�W�nB��wa
�t�з+�������1�B��o�;X���f0q.�(_�<O�IV=�ps���K�@�ft[N2�J��[����D�I)�����=��q�۔Dtv��0�8���Q�%���%�����t���O%}�ï� T���К�Ȋp�������#��i���7����ю�?� �`�]��)=1�����z�q�F!<\s����,���2-K�
y�� ��܂�b��D���0�t.�Y��.*�%��7��k���m�0����9l�C{�q�3��:ky��$�X��z��ay^�+��'P�������r��Y?�x�f8[-KoZ< ʊ7z�v!��S�5j����2 o���7���:�=��N��Bt�n�6a{7�=a5�A�-5rШ�����2{�-AM���Z��1�ʅo�w���7��럗gs��+6"�o�9��:�#)��Z��(�}��5��MBC`������v�u-��7�������MQ��9����k޲�0	 ��G�&6�48���_����lo��n0Y�I�lT@�`���[.�5#���0��1���c���,|�<{��	]�S�*%�_��
�A��{Q't�}��v&��:G*�kP���ZM�3
Ч�5t·����ț�C[�M�>�H1���D��黽���g��"R�'%���REJ�������S�:|��tz�59���:���\76/7��+�:��óG��|�<�8H�[������'���˗�3G�}����I�ٜ�R����n䀶�i�em�2��G�x�*O���[�T�(���8�������}R�*����p��zQ�o��BZ��9�mF5���~L����#�d�F;�~8��c�+K�����7�����9Z(U�eT�{Q�}�q�zc`�65��)��g�j7�	�ѹ#Vɟ�� �Ta��7�q�G��بƉ��bJ� 7{�v�*�{p�!��h�O�|W��5�Z���c [a�v
�9���=h��[��ٷx����	`nΌ\G���0�,�TI?Ip�Uf����&ӓ���t\�q�[��%��̘�h�n1;\��!�L�����!O�#�e��@{(p�mG/GMrlk�{�,���PC2{O����x�#�j��Q_C���O���ۏ)X7�ϸZR���[�fѺ8��mp��=��'�h[�f@�A��WtF(@пt��Ll�L��J<,X*��Wѡ�Rd�Q�BR���R4�Q�R/N����No~�H�����9L�UF��80�+p��"�d�m`��:H�ǽ&�Y
2����ڧ$�"P *�yW�P���>��Q�[SZ�z��+J��Nхv�I��v�<
� 7�\�e$ǻ�Z>mQ$�V2?� �;�����
��.�`8ˆp�F�	'2q��:4Xn/�L����}w�/�E��IB��np����iY�?�k�-(�9�R!ӯ\�s����z�>)3�v������nk�0[C���B�n�Rúpf^B-��q��ź�7:�N�\�̹��N�[��ҲˬEfiR{��(�_���"Lxɩb�W)c�/�=x��S��Y�x�h�;�>��p̿��0kE�L�z+�!�fW6��Ut}��~4ի�T�ߩ�j"Z�M٥�tө�Y��uA�zc���[�����H����9!�<_ViBA�p}r;�_��eוF��AE/3'M��%~ϋ@�7��0�pϥ����p�f=�dd .^���s|�Zȅ}����f�=>^�oj)��}�]�.B��snG䋷n��p�"���HU}bbF����Z�Z��CŐe�A�*y�e��TR�&�.l�*n��e�S�A"5�#�eL�z{���X�������7�D(��{uҔ+��\�?�g3�;}Q6n�ߘ����P��;�jG�T���Dn�Tbȫd���b�ܨp����{a�B�X�d�S�ڪ-��)V����F�b1�O� >�F-<�pه��@ȕ"�љ���5ޅ@����	̖x� 7(#�_�W�!��K4p�-w��n�'�󥠁�3��O����g���MH�J���4�x��f������2��5;I�.q�9��[W�
�S��W���R�=�n*�M� �]�2��=�Ћ��t��0+*�s��1�\����X��kHʳ�Y#1;<�?^/��m�Ċ}�%tg|4���a���Ƒ���s_�%�QR����:���6�G�	�>R �W0.�JS�L�RNwD��P��iS}(Q���1v��f_�3�v�����G�s���W4�5'�!���O��E�=B�(�P	��v�#F���n�aK{�b�]�z[eO�s��i�+*��:����p�L�x�C���_.j�j�3����Е}��"�d�ޱ�>jo��[��>������qx���>�{����-���O�@�v�z8[,=���S�{�@��=W�rN\
��voő��]�	p��[p�V�j7�g�w���0�(��G�-�f�6��-�~�^���8�x��K/� ��El�4Wg���?�JeZ��v������5���$��̋�p���k- �
�Q��P��Y"�ԫ��OZd��ڦ�VĘ��w���ˈҁ
�NW�/Ӯ��r�cK�#��L	#m�@թ}���,�o��(��O"� I��S1�.r.!�c8��~u�խ5������@��V��|-��:��1c�˒���xS��B|���\p��_��w+	����{ b<Ъï1<��i��l��鐲LG������_J����v�E6`Q��s}ߊA�{0��փ��KR��*J�aA�n�=[���֩�����MFW�a�/�tGl���̱�����2[<�w���\��bEA��Jx���}V�<���'x&�7q�I/�7xXP�q��{����>j�#�A5��[�N;wߊ@�1й_��w��lՁ��uv/;���|[��Z���q�k�Ћ^4QH�2�
�R�3���q�ޏ�bWy��͒Q8N�?�\�0�7�Pew�l?�A�`��|&��9.F��[m��  l��.r��b��\C��C��=���}Ά��2f����4�Z��y���[�E����L��i�d�C��C����d��zBʚ����Ƚ�QIe%N���? ��e��,r)olo@���x�ǭ�z�ݫ��N�W[[S˴q�1G2��	6F�=%*�σ���l���mJ4s�S|'y񮀦*�0�c�f��ky{ZŸX
���dB�0�M���i�&$Vdhx	l�R��&I;�P��)�>�/*�e��� ���o��2��	��)ն�H���1�cf�������'�3��\oǅ=7�W�ӀLt��D�99�`�h�u�:����˔M��t��y*4�ξ�󄰯R���rd�`�S�R-���xZ���	z�D���W�k���w?�5����p�����20�g��M;NQ�8�~eK��h	���0�O��{�o���fO>Q��b��dj��������]Gu�ڌn�>�p�$2C����I ;���B)���<I~K�P�7I>����f��������3�R��e�YtthR��wU�}�y�Z>��yօ.�~_�6{�_f�h��<��f��`�4�D��QƩ���nښ���0#"i��=[^�j��%�tY+0�˻خ-v6A"0��4����
�%R{�F�bW���7��Z�0�����������ri��*���V���d��o�ͤJ�S~�&������iL]x\깫�W;7�U�g(i�1'cq���G�[]���Ī���K����{���vS�DB�\0u/�*_><���+�/Y���7�^}^��C�߮h����J6��ë��d�������dF=�@�"Jv��P��P�f��|��ey��.���n׊5(n��V��iG��Qq�B����oN�G:f���2~@��8����ьZ�f/e>�-UO�dm�^�P��`%�_j�T�E��Bid|�l��H<�kF	� Ԭ:+�uI��dv��A��6�P���xN�9��D�I@��P�u����xe�>Ay&���~�*�v;�T+�65�dw�z��s���`�ML�P�7���*��w;����nP�~J�Q�Y��ߝD�_��c������H�02�sK
Л���-/�X����<\��sw��|T��I�g�ߒ���g��8�)f(�rq(z���>i�G8@��6����1r�������6f/y�BFԭaP�4M#h$T�������w��f�9n��[��ٺ)%Ëۏ 3�����F�W���×K��OD'�<qm{^(�����ĄZ �ߘ�wP�v$��[H���4��  &$@`��'����I	�^��`g�~�z	Y�ƤejF\|��F�S�(���W����ʨ��}��o��,�s��g}��)�M,�oԁ?����SH@.�T�ݺǣ�Bܶ���G����E9�#��|8ʒ��8xz%�&����E�i} O�\��6z�W��c_�����ҹ9���ㅰ�w�T��f�8ɟ��>/=�d[8@�������[mT�`��ԥ�}�c���77���&���M��eؙ�ٜ/QYI�c}ҍ��X��0<�_3t*���������g�5^`�K�|R�����u1*Vi8P��S�5�:�^��~�Ev�O'���uNuV����e�+��p-���n������@��MQۣ���1�q�F�zikIz<�p>�Q $/�OIi���4^<Eހ��qM�0Q�B$�A����IS" ���]�����,l���ީ��]W�qE�I(e��ڞ���6c������2��T@���hʚ��y�~��hBX���Aڳ/W�z�'�	�Bu^GMn�]J���ז��Lo���10���ǱDr�rg�3>ҟan�l7�LB��K#��tp	6^9Yτ�?�{�[x�qG���S.9��3#,�I�N��Y��IT  `<�>�S�U�g����΃�s��X/���W&��e|-�Ws�u���]���P}Ô��K���Dc�i�퉤�#�y�������M\�T4��#et�����Ge��B'�y�����=b���0�PC��.��'W�<WUa؁��	cK���Ç\��i�dQƜ����@�r�xl�Y��
jma5xы[�'d���{ٔ�7�#���B�9?a&�E��y{>k�E��59m��|]~F��BBhc�����o�����f�]r����������[e+�}u�K�\�\���HM'`�Vo�E���"P�������Ѱ��w�/0ŢT>������ŝJ����������ŸC7�,� ��y֙�.��z}�ߢ=��q��-�W�E��EL��=�#ay�8(|�7ٙ��J'��g*�B�H)�X,�PjPk	H~j<z�;�ǆ��~O��o�QϹq����|F�n��%��3���Y�Z���a�N���E���а�)��`($�_��jjLla+ֈ� [��!GA�W�%�Ϻ�C(�H�MF�A�9t���#'p*H�h�hLʜ���5G�����r�+�;O���u��.���X�)~&�<����7�ummI|���ゖz��o�Rt�/��<�U���?���r-�z�;�]Ԑ���]U:.G"G(�<��~�7�[Pr�X�U��E�"vb=�сi ��X �������LaN��_w��d�"1�y=�	����.uʛWj��a���ib��¤)����y��m�ijF��$vr�+DYitD������ ���+��Q�&�0�N�QE���7i�T�u��
�!+J+ι�m�wk��$=w׻wI���`AŌi�nw�z����5�:��ۀ��y��ڳk�5		���โ�ƙ���a$B��\�A�Ew��� >�}>��p�a!�L�����j�e��?�Z��)kT՞���R����O�w�r�]��B�m��"��V�ع_��1�Q�5�'UD���?��������zI��o�������#�N1C#��U4UU�K�dԗ��g0�,��g>�B'�rk�H���fw��kGǫ�<_>W��Q����"��Q�d�S�o`����E��j������4���G|�6&$����jA�Ozy��d@�WQ$��L�5����8e3���S���.�؂^V�t�+�k b����M8���f�5Eq�;�g�����Y��S�hjI��v������F�';�L����=M6vSus�ޓ�D�)e��e�x�~i(dl3����"���8C�9t[��^�?J��)��t]ߝ�!���a�(�8@�5��kL��rJ+�{���9� <
��,��Z����sK�"�.�����"��h�~����w6h�R�����z
r��41�#UxG��T:�tñl�$��lO�6r�a��s����$�s~����[�W�#���>�An�y�������T����J
�4���5ػ��~p�j��T[1>���Q���h`�G�@�y�c��� ���|��`fe��9�R�W*�K��;� ��R��pǘ6�vdѪ3�pI^�'a/�cӴi~y�°�{l����רp���K�`��*{�C%|��k3-��A��Yn�Q\�?���#k��:>����}�`�+�`�kF^��$�~�I�?��D�x?�˨ʻ��V,�$��c�$�U��� �LToV�o�.f j��N��!��*��i��SʅD��S!0w� Q�D���6��{Zˡ1	�ͺ�3������Uv"CD�C�ZSv��\:��B�اA����c��S�Yn���9 ������!�>nO��?�<_h�	�y�87i��Ma�Y��"l�Y�kS�DcD���	��隆)���ƿz#T��D�1_"�[��x3c�O].\�岛���W'�H}I)|2������k�;��Hq!�yw�]����� ZQ����dV���y8��> d;��鸍�%��.T�e�WN�@�BJ��a6���2F_��=�Q[�n�~8
���)SCi�C��4
��#�d���
W�d=�ҽA�����y�2;xg�{���C!�5E����w2S�@�e�I�* J����*y!WK�Xu{��5c�::3*lR�������ƾ�+��4��m�a̚�9E2Nm�et�
��"L�[�K�;ß��*�J!�S���FrƟ�C>�0��},�!�<u�\�-�ԯliB��TJ�&��ݲZ�3��%�yx&[�{���tH��|����3��-�.�a��НQξ\���g�J��������㬵<�q����Qٴ�ѩg���uu�'+��ː�PF�4(I�A,Qqt�@�����:�L~�v��D��<�*hj-ʫY�ݽ�*�Ց'V��ٻ+� Gԏ[�奟���W�c�	����JK
�_�c6y�M	M_�smC)�������7}�����ѥT�����+��h����Œ\b�^�,�!������o�̠ǡ���6L^���Lx!H�)2\��|��Ѣ`�a]�z�M�,� ��X��Vڗ0R�,Et�GHh,��>p�VQ�.�p�=C=S���i�J��8 �V�e��UR�+�UJ����c����(�)�J�_$�������1�8�H6�NS`�ԺT�_��I���-��}m�g�nAL*l�\V	���W�.�����A6�챂Y�
���Y5,�c��S,�n�MR�>r��]_	�43d� %;���=9́��u�	�+Q�Y���X�-�c]ݨ��f������0�Ȁ��hx8bGF�ŗEǢ+w
�츄�����U�$�O���*�W�	N2#���bf���[��S����N����.� ��r�U�um�D�[��'K�Z������mi���t6��-��B#.�&��9�3J��2������J��*�O-��H%Z%bZ�H�i�+YbPU���tm��Z$�ޥ�s�(���}�4d�圓-�aҺLo��M姝���\�ʰ�!	{?72j�놺+k$X����`���u�f)ʠ�I��z��F0����2�u&�����dU�/C�l&
�jn;��t��q^��Z������ r3Vob�#�Ea��E9hݰ��