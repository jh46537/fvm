��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C��_�+��+��^���vZ�r�Ln��5��[�nj����R�fء�`��vW����慵e�d�s"�2.,�'�={���I�s�O�*W�Mt�`�X�n%��mUe
k^Ubۦ�D���
�<��ŕzї>>�"J�����_Y�3�S���dG������QKh�% !@xj;�c���2`2�t�\���ĸ/��=�C�(���T�#����p.HT�
"v.�ȍ�������Obu�i����~�1�{��G�,��1��#����y�k+�1���z Me�T�߀�1^���%_�K�/#�5}$�N��)@��ó	\����P�t?�N�b��z�ԓt��ms _�΁�g���kƆ�3C4;U?05Q��hKY���ۛ'Wg������@=U2���v�B@��'�1�XC!;�`(*&Lc�8��l�;��o��)? �x��	1��7p��]�V�A���c�)��׷�D�4��F����D�m�<@=�<�|>�_��|F�4��0Ø�4��d���}���O�&]*ɹo^������/�lB�f������)D��?�	��Z�����f�|�J���7�칌
�L�2�9#�{|F?���������i���|�A1�&O�
)��pݤ�{��j�ݙ���?r�_���p��i�Sf�V�����)�XΎ#��k_�06��2T�B����-f�!`~�\^t;�W@�DC������Li/$22�PoiXEO���1ZT��*�ut���ʯ]aЂ�A�#�Q�Gj�Z��|)	~�E�aВu�ߓ��ꋭr���ӉkK!���whI���@p���P�)�<9?�o@�^�7���S�	X6bQuZ��>w�|�~}f�ْ��I�T���^��&ytO��Ve��nC���7��`�vp�9\�.:�r�'�7������ok_��̅KK¥˫��͢HD3B�z�5�K��i �i�9,��/�,�)�?�g{{�5�J5U���'i�Zئ�����d�|G0>AA�<��j�E������V�� �	>�'3D�r!�x��ھ�!@,�Dq�g�{3c����5U{���q�o���w�h��>�2^Ks\ֶ�#�N8� �d�J�#b"r�\����h���i�ޟ�,�%'M����+���#�aϏ^UC���*����<$�jӻf#/���6Q�b�E��� �h�|�Z0OR.^.J�o/U�
&�������h��`��?Zo�e�^��{��K��>�P�!���T�H��e��`������^� .�3�.`��Y%UK�g���k��F��G��%j�K����}�$F��R��7�����kdh��A0�5Yh):�d�~0\���R�\g�pN�����|��_���/���U?ES����n��޲�g��W&U�Iݙ�����l�v��H>�ߵ��f0w��G\:�k��2vh
Gjk���P�ۈ�p녀�T�2���<�7�w�X'��Vш��#>̋�}��`��O���1E�[�����\ؗ�C�m��~E��#4o@�	H��:��k����"h�|J�0� صp��e���Y8]l�J��D���N�Ս�� �����L�)��ѳB�*]�ɉ'Tf�&�t�KlFw��ǜ����/i� �lI�D����U
�q��S��K�|��Qb�-C<�ƞtq�D{u�Ѐ���x�D�饴�mg��j���j��1P���!O���?%��=y�v!�Nb:NK�6J�'
�![@c�\7���$݋��=m���@_y��y7I=��j��}�WwBl�8�R{d*o|�{�?K�0a(��-�P��鶃(%rr��9�C���W�M�4Y�#��E(+}�Qr�*��6rrK���tV�EL�#o
Eo�xz3�g�&x�G�"���]Zi!��o��X��BnY����h�i`bB��I��N�F�:�UPHo����Q�t�q�뵈$1䮚��rtm{�"��U���#��򿛥�0_����]�<}�<;q�*=S+	%h�wM���D��s�z���b�O�-IRᕒ(fޯ�MId,�%	c͗Ұ�͠,}	5�y�_��=�d�zV�Ŷ7hZ݀DRUy9�����V�n���1���oa707�.о'�uN��n�Ȼ�6���a��_`��Y����<�O!�-|3;i-aX�ǚ �����/�lBE�ss�k�X�[V;x�s��B���KI��{��3�Ø��H�	�Y�'n|�x2X ��i�h޽^Go˷NM�kK����N�K���UY���bþ���=��qq7ˡ��tu��-i��w�M�{�%!����<�6W^ө�q]!� q�*p���������ӻh5����*��x��ሃg|ςs>:Jӡ�R�)A�:FM1�3G�y��L��ӌ���σ��	h��L�f-���|*u3h��v���@�ϫu�zz�� �p�	��e�[�f�%&P"˧v�" \X��~?â��5����SQ&���9�%�-�
��o�\Nvq�o9�^l��yi%���[�ON�t���Pj��NʛJ8�Z![���<���������x�c�c���"�,	n��\�-��l]�u�t�o�
oo�H���"�'�m��pMK����Ӣ]2pU.
��8�r���2+�*�L�,<�U\�D���"J+���!���}^��(E:?�ngz�V�g��w�ZB�D#�����$����W�_~�V�_L^�P
o�����sÄxp��+�C)<(X=P�
/�ۤ ҘrH~��k�����l^.8B/�+�z?\��E�FA� �a1�a��#�d�H��~�&=Q[�<���ڟ��1yG	�I���8�5;�Q�Wx_L������k�`�ݴ���U��ƾ�d��~��˟�댏�KL�-�,�b�WV���~|E(�O�K�!J�G� x-G9���q�ݘi�������������[/��S�u�<f�z�v�u�(��D��Iv*����'������`M����HT8<"�3������PY���4V%�X����їCĂ�I/�'u��%BX���Y'�PD� {���P�#8�¯?��P�j堌���d��/M��쁼�`�/�A��m���XU i�,����0��TI�σ=���9z�ы����Dbd��9�rj��o�I��ڹ�l��tj֬J��7/%%��0�J3�^yh�F������A�s���5�_�k�m/.��u�]���q>2k��Օ��A�"�%saV�>��@ŭ.m�&La :;r�Uuh�7�3����/�aۋ0^��^�h'�,K��wJyFz��.���V�K�����O�C�Oݳ2W���[����J�0�6:��j.�W�m�7��}#�\X
TRt�0A?���C��S/di+��0팪�v��P�?B�G�վQ�35v�,-#�,T�f,gS�=����r)�� H�qw(֎n:#G���p�RAŬ��RukP�fr��Z�?�c!���K&=�	4����j����&uO�~[%��.I!_�l_��<{6r�4"���@�ߣ��v��K(E����.�M�����:�%�6:n�	F�7�݂��k�o>h�x�@j��n���@;���W
A]��)��
�GrVӴ������ed�A?tHQ��*ܜv�{��o������V�	��S�jIÙ��N㧭&�CH��D:Lw�,��*�?P�� X0������w�)��3���.H6����^J�[�������
J�"�q+6��щ+�-���p7�yku��1���`EC �M��(8���+�.2���}wrLvm�kP���<��H��9�bZ�c����D����{e�����D�q��yM[�û��R6Im#��<)�����G��\����GаS�e���yc��[� �c��0������d`��f� ���h4/|�ӑk��S�*4iۏ�Ѫ0��5��>��ډu0Kr��*��1�A7BǾ`����F���R�rC	ø�i�}n`��!3yK�*׻���K��p�o�qH�B�w����cq:YVY�@+�Bi��� pgr�j�C.�}c`Y~J~�	W��`�)�ݘw�O���nj�� H��:��[�&�/�M�U��Ћ`�2�|5|�vGY?����@q4�ꏱYյ����&h	�a�aq;�\`��&���Xf-Bo)�z�G�V�$���OVl����j ��u��hDr
tD�Nk�s"̬���zkҜU#�ڪ����� ��Z��z�T2EB�n3�Ӡ�)��;�,/ot���#?[T�,�J��nJz����1j�a�7�"8M���n�N�9�U&T��s��]�U�+�?�ׂ�s�F�5�}�,
�
uq������z �u�`f� (�������g&~F��~��Yބ��������#�]-���a=�]�.#�Z`8��Ftc���6ƞñe�	k����y����V��~�̻Zܱ{�D��ב�`�^b;W�"$B�������N�jf=�j��e�dq�KY�G���[B6�͞>�����@��ښH{W����Qm���uh0��,����%k�]#`�̇�Gf2�Id��"�e1:��Ζ���ko��ŉP= Ol�d�"rN��(L[̝�)��U ~}�?�͂��S��b/]إ�2���{c&s�~�G�<��1����]Ň��F�@��N�N>��s��wAM���x�F�#��D��ǿ��hCQ�9�H��#�(��{��ރ�a3�y�ړ�F]߄���6e흼(X��J �YVX"[�8ٙHs����s�%5�̌�\a5����7��������(v��H�+jL�YԐ~u4��U���:��vWϔ�֗���:&���#��0V�2�	+ɧ{�?��	��a����ъ7ƈ�A;��E/`B$��]|9�����Jc�Sx�B���1m�y�o��\ń	q3Y���Q�3��2��o�V'�@A�k-T��a˃��@���<�0q�L=?�.T5������4=�v��B��˃��{�}׏��ř��P�ώ�#?>�/{��� �C�:�= �(�RK޿���c}����$���3F0�]�.��h�]��P"uj͇�.�Հ����lt����eե�s9��L]�7���DL�{b�t��;��|7�Y,Tcm���iӵq�����Xr*'��j>=m,ZF|oTHցs[^�:�/`��Ϣ)�j wP�I�S=�8�x���F��M$�J&t�2)�><�i8.�Y�H:��q���7���Pm���җ��}B&_�FD���3�jQx�(3������x��L��p�c��
=NJ�S0J��m,������w}>PQʠ���� �T���!�upB$��D�����P(5�d�`�� ��S�^����\�B��ER-�=��~�[��E��i�pb��#�U��7�F���}]P������<K�O9d�#��j��NX�@	��K����y�rKl��@�8&j�J!]x6��<Q^q*6���q�.H@�(7�@{�۸5�E��J�̫�|ć=*@��YLXԼ��i�Խ$�,�+�L_m����ŗ�?��kR�=� 9�Ҙ���L�b?�6��)�����+C�kƱw���\rj>�K�'s�F<H �O��C9h��Ѹ�n�g�� %������ ����B�D�w�z�����K�4��T�}ti��H�&��})6�"9zB	�"B�H����OX��h��  O�t��m�@�?�[�b���g᥾��d�QE)��)�$��Sy@:���c>�5�}r��&�9���2�g ��"م�.k���pLE�� bw+[��w�� ��DZ��	�Wr�'����<?�q�Gu����������x�p��dM[D�6�Μ�qɃ�5���fB�ßoY�6z�V�3�7���z��h���_s�[c���?ʎ��Ly^��9���S�'a�ASV���[�#��;m��Aҕ�5:֬����2��������yx�@|_˔�&��4z�袇�]
G��)DgG3�l��D�_��r��������f��鋔h�X�ӾFc}9\̘
�*�^��Q�$����|%U���` �ꡏpx�lF3HXa��[�ճ����G�ϧ�r��1��z7�.S��C�eR��c�At��Ao��g�3C?�c��'� �8����,�6I�����ߌ}"m~ڇ�zPu����&B}�>:��κ��0d[��b�����Ri=�(��"�㉅ɒI�1]��T�#�v(�m_�F-�|��ĒҬ��8��^i~�O���fF��6�u3����4ǇZ.�
2�"O)��l%?��xQj�	s�o*��iz1B���I�:�-�ϖ�K��+s��]?9�־GYrKL�-G4�
�h�J��E�UI�1p�zM9�� D��%���A�a�P��@(�lhZ�4꒞�ֽ�OZ�U���(�Y�{�o�t���t�����w��V5���DTBF�ba�Ei�Q�W���g�jcL��ӭ���9��j�EQB0R3%՗��yf�zv0h��p8�Iy�� X�~6y4�v�p��8P���_��f�m��gv�B��T�N�e�@p��QjF�:^�Ԛ&�#���:p$��:{%K-��n���͝����y�BU�h2 ��-2�i���V^2��=S\y���݆p	_��R��BN:4����q2uNZ`k8Ix��DS�˪WY��r��Z�M��?G�a���jD�ΰ����nu_E��
�r��5���Q�]*{�77Z�#��N�CÛ�M��RU~r��q` �1��ϒ�=����ٝ��LLw�Ad0k�1|<��N�>��Ei3ޤz��{�sst�=�J�!)]]�QR�إY���RK�_fK�r3{*�-��ھ��1]��p�kYl�R1�D�WVW`�:��7V�V���jj���	�.C,]��{=�Ϝ �9��5����g�;���'u�8����K���C�e-=� �k ��&H�t�&�:l�(�����%�;��l�Y�X�S#٦T]0������3E6��ux�>���,c$�BlcT2Z�:}<��d�D$k�Kf��>�K��C�9������5]��Ky9���MZ���n(�!pl�W`9�.��'�}�|�a�@��@ټ}U�_M���@E�x�t��gj(���
��b�6zw�L ��ˌ,fa���p�x�h�y8O�S<��*(��]��<�Vۋ�+/��y�G۞�KH���Xm6(Y17-���c�2��)Up_�pL(�y�3c�5�f݌ԏ�йƈg�f�W&7]ӡvRi0�6r7��%؃n"�pV���G���*	T�Z.&Xo|Ә���M�S����8�,&=���3e~&o��G1z��Z�=٫o8x4b �D����J��W�hRL!���)�|)��Y��<|4o9%yx�SE�Ñ��51��_X���Ef	b�@�Q.�
6{���1�{#RNL̈́>����\oĒ�5��
; t:�ZF��IࡪVe�<b#/����QY:�d�]�Iy�6ݧ�w�f����Z
;l
n��):R�� ���G��Y٣�?�S�$�zT�Q��rD�#�T�����C�Px"�����:�2͠=���~_��̹N)����ة�F;}�Yi��!���������}�Hf[^&�pM�M��A�����'y'8"Q�ޖ�6Q2��?X�ނ Px�J%~.xF(�hO���D�����n�n��ɞ:@�y�c�[!ڃU��>���g�@�����N�J�c�I˗�
����ZJ��*�TC��u��n��/84'���S�Q8%�鬼f�Ѥ��:a�\�H���ʽ��3�`�w��#���_���Og�n�{�&~��d�\H����,u9�\����#�+��������[����]"�T]=����;�-ƾPodw$a<o�C7�O)!���3����4���f/,.M���T�W�BZLG;WO{5���s0J��Ko/�����}9�;QW&�L�:\
����;�_�����p��u׿�?��B���:�>9�k��vջ��R��f'�Ĕ~�Cu��Я�bY�����ɪE����h�=ONԅ������ꬅҰ�~j�̱��Y7I-?�t~���|.:)�p=�fo�|������~�#�A���r��իW�f� 'U}�s��$Q8/��4G���<\ �j2���(�C��h&a�	�����~3�h�8j<��>C����:>�O<<�+u�Q� ��$K�#��r�j]�P��6��*TBˎT
8��,k���٘q�+=���m�����`Œ��&H�%Y7�;G�����]oJ��n����OF�k��?�=�VD�����&D�X���ၤ,�i�i�)>e�&��<;�V��ġ�h~���هWEn4a�΍�Ds��^QWA�j�/
~[{ܪ�)vޝB
�(�笔l���K�V	L� 6�rũ�8��F����=@хΉ���L�� ��;6�����y��o��sN&f��0\�����8�zPEɱ)�O������KH)����*��-i�!�� �[��yp��>���v�\�̃��Mv�Яw؏A�3R��~�c���Av����6a#$Q9���x���/,��t�
��ә]ј3�,��|��.��l���@v�/q5�;�ZV����:�%�|ʻc�1͟i��rq4�B8��Җ#�.��sJ=	�"�$�d0���KA��	��G�5�j�M+�z�C��V�;^����B-h
���5!>�����x}�5
��CBQ��`q����ǻIE�����A���DE���-A]�m�X<����C;{KG�@��'���l`&�d[�7���%f��+�A;/YU$h�RI��J�M��Ȇ߄���#��-����%m~0����驅�Vs��L���t�`W�ڏ�8@��S�3�.E�r{T�pQ��ΒbR����^����W���)�;C�o�̃�c�d���"n~>^K�EN0�����S]bV}H��/g�V��*�	��%Ck�[9��-4aIE���4tA?Qɩ�)��7�q_:W"�D�C��c ��}�g��é�Qg��}���� ��y<楘=���`T�4T|�Q��Cޗ�y#��m2�^r�U�Dy+�h|��5
�E`W[�˵��zP(K�K{2�n���G�%G�͜��|.�_�j����p�Gw����8B<_�J�Ӊb0-Df3�1� 諯�za8bC���d�\�L����dUo_�PF��×���?���UG| ����M;A�����䂅�\�Y��"�/�V۱L@��89�@�Y:�*C�D��0O��"�2<���$3����멖�]��.4ڱV.���8?�~��܇�Ft�=L�Z�x�<�)�P4���!���:**8_zM�q�4����_�]����m|}A��5� �Y�Uq�w���Aj9.��n.��28l�;8��B�tƶ})#�^�Os�x��?��q�`L�b�J�����e��4$�F�X�~�"W�Q����oy����a�	���	���l���B�N�щ��EN[����VX�ѹ��c�n<���N��ԂYL��Y�J�?�ػ��F�0�ңqS�;��n'�.u�D1,���8n� Du�f@��䵔:��>���]V<�gr�+�m\�u�J��@Fq�g3~����F��g.,I�ɞ��5�¤�GI��'���Gnr�]���Yi�H<y�/W�O��;�A]-R37����[|�~�B��3gU�kB��i8�����9!Ho+�WQ�h{
�P����*�%+.��3OA�1�8˸�&�$���
���M)���:A~��<�E>�Ew"Օ�����x��Qcݺ���)I}[F�����h�o7�T�k[0����`O�8w��\��}�K2Н'P�VO|h � R�O�D(?z��r��B�zy�e*�/L��k� �����YbXb;}BO�S�l
���Lʛzz��z�*��%3�+�����lL�kn����M���X��EP�5RT��e��fx�R��8�~V|�����y���g��`[�V�Q��l���ƌs���D�I�f��E��N�݂mR;x;")�2//����^Iu��.@�/�&τR9�*1���}�z�8x�m"�J���B���iO�b�{��w�t+$���v��1��,��A���xK��-FX�
G�0gn�Ǻ�~�)��1�!�؎�V�``2�뙏#t�pN��]��B;�أ��4�^�=o_���b �W���T'�3�~ ��hg!	8��jb�`<\���P�4Ӭ4��ȯ	r��8�_��,�F�&�$�5�sH%�$��x�G�Zs