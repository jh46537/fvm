��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{9v#ɋ*�j���-=���2sȣzx��M?H��חsY�]�Ļ�}ȦؠIwٯ7��+���9�O.����!ąQ���:�隼V�}���"�>�N�����x8o����Q�(u����aQ�ݪ�HR7�����g��Mڣ�jE�+���B�<����o��%?�?��x?���.����5ФȍDo���y���܎�%R4�������w1)I�D�3��5��[�B�	��;��˙�49!�&w��=
���wDK\���4�K�)M�@%�)F9�%񏁹�8YL�v�껁�+���%'��:�S����/�ЀpRs�ɴ��+Z���$�>���k���2�51�4ؕ6�/��o�5������w�Y2�h�5�W��\�BHrI�_74Bt�-R�?sGLig Vl� t唨��'RT�A�ףu}�Q�ܪBy�Z�;!�ݍ>�,�pٛ��G����h�����J���h��=�7�e��I4#�5��$�OX�FM�z��IP:K�UD�X�l �K�_-� ,�H�8��VC��3�� �쾮��u8Vu�8|����t)�ݳ�8Ҝ�����\۩T���xHZ�]l�i,>�X�3�򿳒�����nρjžw�"��pj�\�Z}T�H�k��C� t&��Ĵ�N�!��=�M 炄�� �/��6��5���m�`���8b����E�D�a�����P�k�U�:s�)�����%�aM�vK=Y�xd͐6/���זA�	bN���k����<c��o9#|���������2Yܴ.�DAĜ+~�ה�9)U��C�Gv���_4�#�F3�<���e�L.[�ń�r��!�<����{>�(�m9b[Yɖ����&�ޘ� ]ݨ	��ks� ��^�ì�I/G9,�ND G�YϷ7{c�<��5�1��\z7�>�Z��0}]D�`=���H�ߟ��˜���T�˖����`�?=�FvżC��h\E�zټ*,�G�\C�)z��ړ'y�cP2H��Ȇ"j��=���R������&����l(�I�3�RC&Rf���A��R�{_��������	�y��C�gۍ�a�����֥���7}��D�F"L�2�?/n�%�#�*���L��Nf�tfn�N�!zb��z](��Ko7>����gH��3N�j������\n�=k�O�h�:}Z�ݧ|��c����G �����oF���K��?�Ap�xﺼ*��J�d�,��P'�GI���@/oz����s��o��H��ґ=�|��j!�I�WUE��T���p9-am�?�+�#\]���I�G�\�d���O9$�V���r���q�!%PC�Fӗ��웍S�Ű�����褌�~Q\j�%�q����֪�k��_��P��M��։��=]Qi��7��	!�Ĳ���9M A��������<_�^L>hY��u���!�ub;۱Vz�TY�<�����>Oz�u]�Pr����0�wr٫.VN
IoU��J��?�KFǛO��t�T���g������op�լc��B����de~�(��b�]��.{V߀�����ą��/p��r_�ɥ���E4Z�H:�`#z��G�HF�~���\�>�%�#�нA�Cp7��t0�P��Ŵ�n�]����1O:�C��rWor۶ƨ21�#J��j�c[^N���{�4z�wБ�;3���|>���%��N��'�]��VU*1�w��ԭ���o�f�QJ3�yz��[eԊ3���Z���rpB�"~�r�YX��}^�TM�e.nv��G�'��'���h�|�V릶�a\��	`� 19�ۤ�?n���W��Th�w%+4�!K�C�}8>�uBRU��ד�ع���q��CZ>\~�l��	ȣK�M�]����'Ds`�ŷ�@S{c�p�<�  �H֕��pU�n�U,��?
����}f���5�I�c��!��,���ׂ$c�/@����L��1�t����YE������O�XІ�l���{6��a�:��Z��8�+CD�y�Vo_�P�bF�iC ^c�B@�n��h��V|�밚2.\�
��xk�PNC���u�f"E���@T�����:�5�Y2uk���4���]��?�2�3�(/9d��ts��𠳎�	}�_�w�u���Xbi��E��,��j��N%�R �\��s�aH�	���:�n��A��vz�{d8^�d��C*���ݮ�8� R�zWg��������H#x�3�H?�^�P,B*���mb
�D���>&��Vʤ�T�7rE8i��6(���f����d���#L��v��ɇ� -��t���ĵ��I�4�V��D=�Ҟ����jl!�Zg+�f���y�]�%h�0���;����5J�,!��Ű�=���!(?��T|��� ��.�HT9����]F�\Z��,xD�q�4�,'�%��b���:�}z���Ar}XUi6���R�eܮx:9�ˡ���G�划̵��5�Q	�)�#��7t[ƌ���S�F>��.��b�������k����* ����K�8�N���9^!��"a9,�V���a�D�:֙Uq(Ae�-�YĄ�5����TB8Dg/U�D:�v[��i��U�eʾeq�9R:��v)��0����P�M��m[�Z�N���<LV�z͓Ȕ�6uU�0��<��-��>���	#.��K�hW(.����(_��j�%��ɗp3��)�}�b��۫�@zb�0��z��EV��P�f\W �� ��m�4�F�
��2��?�@
�M>�,SO��>X����wa��U�υ����d�H�e���.��jq��M��Yӗ��3cXq�c�R����Y|U?�L-�M���b딽��a+�����H ^�f�ML�K�{+�����O���3a��vw|\��S�J㟮lnxx7�d��W�A��)�k�B,��=x���W����?eAt��{<yڤ~��0�,�A�A�T��
�5�t&{���p~��^c���؁�O^�ж���|�-ߟ�(�Y�m�J;���Ƹ��:�̚n��?��P��W�_��[�P�3�׌���G�~���D>e]���]�eЃ�z�lc0N�f�#�*��He�����iju�� �5�?Ѫ'k3�h��*%��?�;���f�ҡ#p�����?}|��SE�E���\dy�6��۬��W����b��	6,���k������8��q�I� �G�A�E�p^���I�[�p��x��N�����ѷ/ W!K�*��V�N��!}7xɩ��3�p>ݾIg��/�Ƞ�X!��	��̈�WAe^"�},ӆ��| 暯b�d/�X�rPD���zԥE,�s��P	h��շ�~����\�G�$)��~�O+(nG�� eq�E⅒�׸b}��覂q�e&�����,S*u�`���uR �c �R
�; ��*��P�qW��T��-��A�z�P��iF*>c{ݤ?�h��¢�=ѣ��PT&��������բ���Y�jr/RЋ���;� _k,�w���ړ��1|�i"wGےB�%�U�Wa�C�K�%��R�>�z���3+u�E����o����3x3ӌ�a�ְ��o��&��6�#��P�,<�n��bC����9�t ��r�%���ʢ�luR�I#��3��IA����ٸ-o'T�ރ#o��PKE���k�('Ǣ%E���/.z�Y�6�c�`�p��m�`����9��~3����O<|]�j� ��
��f����]_�8�~�e����>���F!�}�B��N��o��T�Hۧ��<�h��T���OE��=�l �����k�oR�@���j�C �g��s�<�a��k�η��Dg�XX���d�EmT�mA\w�}���;��g�ٰZVi�s���C�y��*�C�u\����|�-"n���μf�=T�d@�Q�`��]�l��
�q��Z�n���(m���X��f)�n�|�WL�N(�/ߚ��Lg4N6�*�W�*�IM�܅��i�@��
.h�+��x�+�ƍ��F�s|e��=���F����2;�~I7�m4��Șژ�f�kB����E���T3wZ���d@nr-Օܒ�� z�漸'�.�$���:4&EY�'���s���g����RA�3��qT���X��"B��ʢr�Kb��rΓ�$��YO�^.z6^(T��
/�.�O��-UdZ���k͛ug`Ǿ���lk��j��fm�>�-�}Σ�<m�z.mX���blNط�������'m��w�'݅�h��h�	2]�K�F	����S��K���g�r���t;��1t�x7��-w�$�Bl���[���e��<�:�͕Θsg�"�Y��� ٪h�:5�kъ����C�dLq�6�^�8�����j�R��Ƞ�����~j���x��ܬfh]�̌2�1��D�(�eW��V7��0$]�*a��m�[Ⱦ�C'���1�rT�{Ț���	�O�}��9m8��|2�=�Ub-���=�{�S�Ј]�^�n`�/����&�Rt��d6�t��͛(����7�Ͷx�4�]EP��8z�Q^��Rs����jӖm\U��4�M?M���)��n���(����)��[�BTс������C۰e�:x��!�b��7����e��M$P��6{ӝ4��'&�^����v��v��!���5J����8|m�)�-4<;������'t��W6W#���H������
�z��g;����1�o���&��2"6bg�'�~�
��N���;��s�������9o;�XmdD��v���)k�I5?�kx�Ê�A�#�ve"����+��a�R������/�\���B�᥹<#4ƣ��iH��D�e#��Z J��:Q�i*�U�N�Rp=��!�� �-B�,�T���
	��YSg��܀P�J�I��~��,Y�����>ħxq|���e��$�ēj�8?��W�����y=UZ�'4�W�Ϻ+~����z4�̘`C����Iӫ%�D~����y-B����҆3�G�Pߖ�!�j��E�K7�ˤ�8�?P�6᠙[�V�7j�Z��(��y�=����"xR�ֽ>��4�����!P�F�R��"Du��p��	`��in�`&�`��xAͦ7����r�g����7?6���:�ӷ�]YF~�MQ�Z�!���3��?�><���Rm�6Zƾ�jr����r�3����K�D>ddS,ߐ�>K�:�bAi�|�$avʑL��gժI#xGz�\��@�X�-�Ly����Q�(��@�k�l3�9���$Ʉ���=����F�O��[�o������iH��ֻ���3Qv�u��q���Q�6�kȵ�Hr&+b�����]ς*��=�����<@`*P��ֲ���T0�]�H����IJ�HV]��𯶧�H���|��t*�pU��j�z0
�b�|�-���V_[6��S�/�Q�`��AV�z̯d5��-q�W���W6�.	�`��(G�a�ФZ�I�U�|�����`n� �lv��`?�=/�� k��ۡf&��N�@TE*<[TRb�������oy\Ў�L 傆q{�;HKt 4���A:W�n�i�����j���2������gÿ��t��p�� �P\\Z#v}��߱a�23_��d��}��ar��m('�%��b9�)�mg��r�/�Hd�ĿBT��� �o*�+�T��H&��h�a'
��.xb�%l�`��qW�K8D�z)��������㥻}�2KIK��pˍ�`��Co�	����E�z��N/YYQF��>�%���0@��ݡk�[�kʬ#� g���;*�1���F���%7slYs�����ND�Ӄ�ݟB&6d���X�I�M�bn�9��6qn�'���qݔ�����z<��*Ob[���Z��9&iB�I�`�ќ�ԟ]0L����?�Wc��RTo�e�\K�|��kr��3أ`1F�������ݚb���:[��* ���R�$�閂u��I
�&߬� �!���k��<���Z ���(�t!�oNr����]����3��?���dJ0M�5]�*�(�oxH����8�Z%��h ����6/$�4B:�h7])J�j��"��6�X���C.���p�b�(��
Hf��g��q]vᐂ �����Y�kF�8�T�
m� a)T��@����Ek��˱�TYձ�=��Sk�/�������J8�o��0vӃ�b��/N<�W7�H�r���o�%����e����MxěF��9yn����&�(?�q�J9>q����Gɟ$e������0v�
or�hp J�J���Z�7:-�x|#l��q}dM�Z+���]�?�Y{���ݽͣ�%}8d�^�Elh�K���Z��z]P���"M�D�?h�0��a^�҂`�;���ϧ[((|��������)��,}�Q�M���Zx��_I��V����s:y$�|���������6�.�|I&e��9T�h���ؖ��x���z�/�;���2��n�xP���� �#+����TI���2K���(�y�:
��D�u�`���������5sh���2�ׄ3�Fͼ]�2dE��
�ٷ�X���*1Y�KE�Ld�sA���"cL��W<Z7Jq�����.�=���EHJP�o���=����Y�F&�l�����O���`H|���,:U����O���]��і��!̕�Q=<��Z���u
�1}�.�ߏ��T�K�X���K%��b"w��lM��$;i�bm<����Z̓7&u)$��Ȁ�� ������_�O�Lc}&�5
�Gm�8[�A3�;�	T��o�7z�K%����������=��d̫�=��ޅ0 ���sz�D���(� ��X)|f{���rW�I��g=�x̄����C�)`E�?g���H�ߙ]D���%�f�s����b��qN;×��� �?���F��ԙ��9j��Y�+;�L�O��Y�����SЍG���wtF�<̕���Α����cW��9N��`���"A�Y1_��w]+��>	�����}�g�`�"���t�����s�e��j'f�� %����N�V�h���YY?)���+%9vd���5���41%�0��3���� _Y���h��;�#Ci}+���i��]/E+z>��N�5��C�է�Kiv��|o�[�7(��f��Å����D�)(�=݌
�A�wiqG��t%{�jb�!b�\Τ���t���Z�g*���@�����F�b�~��\��S�B=�ڙ
�|h,�XqXj:ᐐ����7#�(���th�v�fGh��ȐYn�wT��@���t,�^.=��	N�16䧞xr^�MqW�r�:�޹�
��(3Q��&㈑oJ��`�����,~��ZH�ç�]��ќ�"�#���y+#���E-(=���wd�3#�k*g;,tN���S��|���Y�Ux[1ᦄ�!�:���9@_��˃�}���(�ќAAri7K����rH���`L�I9�o����h8^�eJ>���ė2�FPL�t�������z�=����Q�N!s�ZO�zsY�^�����_ry4�UeSs�'S������4Gu/�3�>B��7���t�.� x��׽��#np2ivv���zvyQ�Z4�pAf|�/�i�>>�i�@��Ý-V�~G�w��;~�X�h-7e"Ԉ��� [���%��(��m�{�S}x�!�M��P����}D�\�}h�`e���X��NȜ��I�6�h��b��LT�%����>j������x�x���2�@|�ج.��4=:��q�*�5n�A��.L�?E] ��7M�x�4�-��ww4��>��E�ghu�6���d#���[��!��/h���\h��:mP�S�ǧD#<U.c>�~�蝤ڡ<T����!*�h�a�4� 0_7��6r?y�YֱͿ��灺���M��%H�}�k�����n�����`u?lw��F9��Xw�������%�S�_���es3[Lũ#}.�/#O���;^b韤�f�D�9]��G�
p��]!�ϻQ���^3Yt
^oF5'0!�L8����O�m���]�gf�E+�����ْ�ŵ�6��]:t�'�}J̵�3gP�c�(1�(���v��5��þN����}�<X6��7�mS�3>�`3�-e�R�}�7݃+��H��,�w�����zFP<��c��@��>�DJ����L{�p��+��r�,�el��j��t��j�3@��$�$�����4z	`���IE�Z����j;�M�#,%Q�SW�fpyw���èq/pd�����˪��+�z����������`�K�GֶI�S�Sc{8��u���>��X���8����ꥣ|Io�~b��5*ǭ�2,T�G�	�_D)��Ru�vj�sP$�n<7�M������2�<��_xwM�nҏr+g����Q9&[y�x(�^KLvX���^-nŮe�J��Sy��;�m=�p�����y-B��6�J� p����vR~`�|�}缙oql��9�s8��Mwf����(��n� G�M2��F�c���R�PZOBs�fz�|x�T���s��KaJ��Y�_�W�����ԕ�,��l43������kÏq�}nw�Kh�!=��F���y�����K�zi����
�	�<�C�W�+&�e�����IL��w�tn���h)��WKٟ�g��C�[&Xe��d{o���	v81丮�Ekn�L|�5!u���L��Pc�����U��KZ�!�f��-�&M �����g���8U1i�T��e���� �&��;����
��c�U6�:��h��g·��B:�@��y�>�f�ڹsY�a��f�,;�=�p���]Ё�C�
�GA/�Tn�Ы~��e��dg%hm@Ѩ?/}���kZɷ�-cY!ŷ��P��7u�W��+��wk��w��@������7�W�J�հ�dR>��;G� ����P��9U���k�_�<�6n��E�n �>u[XL~RI�c��ԨoV��l��I����?������y�	�>&��k���2������^��ו����C� ����h4����(3��rD�m�~ꕮ�94�?A�6�a�v}y�D�nLIHO�C���fR��ԙ{��G�f^�!�  ��Dsb*�)�O��eH��ˣ�2߻wa��PL�3������ϔ�-��`���H�u��xy�N5��]��HI�R�R�O��3���N ���os-Fcc*7�ݲ��|K�4K+��җ�S.�*KN4w�@���h����S��܇��2A`�QUT�i��"S}i��a��+މ���3�kT�TV�P��tV��މ�SZ�n7;��W�;����,1G�L�X�HJ0L+,�/
"��?�d$�3��.ię�`�΁T"��jW���56���[v�~���v�#�i�~�@8��`�R9�˧��]�?,6�)`����(O�������9��4�=\!���y�@�tr�˙�^���im^�О��㽳�$L�8"w-��A@��Y�g����+��h+5�&!gJHq�u���1��J�cc0t�G8�އn����/&{�^��{O�^�� 3?��iR�hEM��pթC�~kw`X!����E7:��G�z�� �yV1OX�!X�yy��:'g�ג�l*�0��->Lٺ0����g�kl�:�9���Q�l`&����\ W+1��wz�#�jb^)�Lq�[�{�u��B�� >�yl��Nφ�ef;B��{�*�,$���WX����vatuv%~&���bC>������e�?|6�c�q�ڎ���{~�s�~+ö8���q��9�R���}��>N�:r"ֵ������N�+j��TjU'�)5aoґh|�qvb,��$�N����Fp���,��P�)z�R�5,Ah��Ñ��g�^+����`�_�Q�F/ =��eoƗ�D4���;����MX<t��9k�J�����,�)�S=VO7�j��K	����]�c�gxvǂHd?7�&"���P���؋�I�cd{Ĺ��³��=�(��S��{����������;u5��3dǠW�!|,	՜rv�Y�N�+�3�,2ba_�w�M3u��z�`�mP�r�Z�.EW�u�J����Pp&��cʩ�u�-vt���k�LUd�^�I��h�`�
�|���輄Fc��|+(�9���Y)E��ј�O}�������3a�����.{ zjx7����nxC�؝���~���]B�!
xp�)�)_]Nq%���� OsH�{�O������N~�$��k��9���f8��x��Tj�U�)�K�)+[n�^�'I�3�\�曤����.�Ѱ�@�������Idn��>0�B��725%��G�$l�t�I�!}Y��vGc@+G�O���[���>o��/�|)�#�X�Ҋ�������G��e���iF7��77/J�����/2�{<������m�U熲6>�i�&w��E��Y>��~����y���V*jD6B�~��&i�=J\��B�N�l G�Qw��䆤nd���:�p_5�w:�A�m<~럘S/'�I5���W�nx�JU�V�؈�fq��m��g�(d	�j	 �n?��y��y��ʵ�1�݂{W������;��~��E�N�T	� hd/f@�R�iFH� ��B�H^8W�Y�"�N]oN[LkFY`?��Ί)xp�BiX��7�+�?J����]>��=��}����M�ҋ�yd��2p٠�s(^�����}O䎾�X����A�t���I�IL����Ά�Pِ��M����4�T)��>��p��p�
BG�P������P�a:I�~��N�e�.V�����{m���[�`��Ǘ,�iǙ�^��h�N���D��A�Y��R3zjD�}���x��=�	]˴�>N�6�`|T1�"�%v�9�|�,�{-'ٜ^1�Uo.��������:k`�μ�yv�f.�1��'}S-WJ�Bx=��-��'�c�Y{��wR�F7Kn����v���я_T�J����b�z�-�	,e.+����@��$����)�t��-�ff����1�4�j!�VҖ>�M��Ο��i�/�7ZbX"|�Q4���|E���$8��2D��LP>�HCa�	�Y~�@����iD�L��=Ѥe��s=@�������D=y\=�B�����	�e�5v+�_�m��>S	N9�O��kI��U�z:~����#�u=��% ��l�L3�i&��B$�<�?wt�#0��d�w�h�"���B�9\A�D�m����I�*��k��/|��ea'J���v�&�`a^6U_��v�Wԏ4��Ŭiub�8�5�\@�!3��?�g����䚀s�0�jzуd�.&��*�j_�;�b�����'aDV��	�n�W����ON�9pL����x��Қ��EW��o�v%�H�UVD��y�=���	�
�0{9�ҋ��Rd<��Q�ķABjs&A}|�SLz���T_:GR/	�#�Zl�y6�[)\�rF�L���'�K{RS��N�W?�&�Pue�	=��[������\�}���(NF5��
n=4����H��8�|��@(l�� �������?�ڕY�U�{�(�l�&��X~��)J�uٍ���s�ږlmn����ڮ�;}6d�,����~tkW�-l�=s�{z"�V�q�H#�JgaӢM��-Y�Z1U�6�y�|	S�qV֒�'����O�C���h�X�(bZU����$a{���P c���x(NuXA�gV��9��[���V='}�O��<�Ɂ3`,��V5E2���Z:���r�5k�n�_t�ST��1Yl"֛\IJ���L-��>�y��eb!��\T��9xlw`��ETe�0�<���=&�*s�J�Ht��ܮ�,�4�k�H�vb�~y��T��c�?,��
;�5�"��߬�h�)#�쌰P�;)�k+Af�mk��{&�'g�1ҕ�E�|��)rJ���3�S���#L��s�VՉ˷TW�;��u�0J�KϜj��O�������?��lNB��\5��ٛ\^#Q�<��Y�ϝj����j��4��	_D}V������~O�)=� �����}�jd&��,ùQL���Y�-g�"�����]�����Դ���5���PC�!�{Nli��7�)��޽bHp; ��ȟ���/��&$k�Ap7w)�\��\P���L")E2��OA��:���?�7\�x4��ز�+ǢY��U��%N��3a�14��Z����A��X�� l2��4�;��p7cb%`�= ����׉��c��u���ҭ�`/M���չ����l�J��V>�Sq�Ĕ�U,��3���"95�ܟv˺�#���*��{� t[�Љ�O�f�i5�7�6�>����/�������@���,B-��%�9���L�soP�O�K�ĳ�+�J�ES�k<�@]q8�>[Y���Vy�o�^��CAo�wJ{	tY�� ;��@�Z!���j|�3�
��?�h�%��TɈ��iA�=W�è����S�đg�o����n��1�;�'�xq�Ü�2�=%�V!�K������j��f�j)*��A��@\�-�Ns���[Hj���Q�,�A��km���
<x�����s