��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E����pbT6o4���_R�&�l37��17u�]pO��*�+:��gvʑ)QH	�.ΏkP�	�.�O���zϠ>�a�6�����Y�{$�-���%�A��/|�Ԙy���!2������P���m��\.^yK6�p�����$��n�ӧS���:����v�[�A�,+YÊ��Ȟ��V8Ϙx�K���V�O�L��� 11o�dKY�^�$���Z�f92�;�v��.�t�෣{��k��C(�E��ҷ|���V�}@�i�9AEE��ZL�$����tI8� �!�@;�*8��!Q~�C��LKr=��� ڜ���Vi�6�	�C���	+��gA{�h�2��Z"�5���eZ�w�0�$w*���C�$�Ч>n�5�������I%1%s�d�|lGL��uԉ���1t�P�op��A�E������⓴Y<Ι,j8����R�RR�5 &u~��Ȍ���HDl�Gɤ�z��{�?;��8��	C��9����P��Wu8����j<�N���'�8b�RuK�t06�y�x�"��!:E�(�������B��ddm��ɀː/J��ax+�u[b��q�ʹW����/h9N�g�/�B@2�nPu��{:��+WM�x���0�dՇ��OҖ�ń�~��oA�R�!	.�Ә+ۋB`����2?m5�P������?
9h��L�6�}WOlV�
v\|�S�2d���4������)��K(!��Շ��ݑs�BH�o��.]�я�=/�H�@B-9��G�˕�ˤ�F�(�3���=8Rz\kӚޟ&m���qd���DX�M�[��Jw#w�[�3
�j��聪
O�Vj5&�&��'�KP�U�����(��F��c��Y.�mE�~�! dاZ7=�	������uUWM**��nt��Ar�RV dw;x�D48�u�)�+M@��!�S�/��IR�+ݢ�m9��bܭ�O��4üA����K#��*�y��`�>l1�"f)� ���� �t��+��~<go����8��ʷe�[��3Q5�z~��G��W��x�#P��TjZ�;ex�h�!F�5�&��`L<�S��AX�b�� u�F7nf-��#m��N�X������|Kg�g&�ۡO��Z����o�~��ܖf~,[K�<�\C��;�bV����hY�jr3��]V]�7�l�Y�݊�:5gLNz�p��ǫ�䮓��ie�W<5����X�]ۻi��jo���v�C����}w�P�k��8T6���(�m��4b�d��ɴ���j���_,W�!^�����dϡ����;��o��}����u�6�[��B���>�32L��0%J��[�B�o$i���ٞ�j͠�_��z��&o�����v�1��v�5�᠂��9;$���/�K͟48%�&UP6���al��K�~���R��CNN�m��Q-�s�@eq�'F���� &��\]�fa���j
��KuVwЪ��4�%N���Ѵ�1tF|XN�c �u#{�'MnQ��{s��ku�\��&f;�����>�,դm����3玵�Vd�y˂ 8Jk�T�g�t˜�u@��Xa�J*��R����knr�屹��_�����S�����#b�qb��xc�Î���+�r��/Q����0�X���K�Qh[�hа,�s|jCH��
�xF�2���:�\]�O'�$����2YЦ�� ��|h�M�H��Md�c���6ަ�/���2\Sh �;T#��v��}p�ϔ�.��d�΢��ԧ��6\c�����ƈM*�A�7�����pm	�đ :������M�E�"��J#��D��L�xS��Yߌ
s�rr�A)��-^���i��$�'�w���]u#"p�{��-H/DwVv����v5n��ͅ�^���������SE�y���K�/�����PÒ�����%�g�j������jT(�p�©O�q��}�� �����R��]�J���}����Qi��3�7���rT(۪2��g־g��O��r����F��;��eb�^ rL�L<��|0o��,B��i�$������:6��������cG���I��g���/�bԁ��6��e��zբ!ifU�����ִ4�$01���e��H|´ ������I��6�_`�u��Gx��oF�jnۧ�$�8�(��� }Ͼ�R����$3���%ǕR���*��?~sD���Dgrp���A�&��$b<}o"@�O���}���A�wE%7��� ��zn~�6/pĶ4jw�����Y��Ar(�>%��s#���k�S��E^���V:�i����E�(�PrɉXr�r��c�r�����cv�G��|*��`E�.��U�mP�#;R���,�bqO��zm��Qf�3��3�ǚ,H�X=��wWN�2)>��<�����sz)G~֋rǊ�.��oqF��csbW��&IFu3����R�c��v��!y��r$� �.��i�L�n{�UfM��t���@�����&�QWv��D�n�M*�X(��A��=�l��݅���k�I7�1 8r��3��ȝH�uu�d�{�~����:4��@ D���u}r27e���t8"ϥ��I�Kl0�4qt_���5.q�V`/�uڑ�XJ-���gL����#�p��*?��
l���կ�e��pE�/���)�/?%~p�w�O��j7G����6��W�OTqDݑ�9g�<���Y�z�q�4���O#�g�SlhśT��Řo���Tm\)ۡ����,�zLꗅBZ�P�o'~q��yo�J�{l�z����11�f�M)GҼE1|<J騟��B.�4J�7q������;HO*U�W�;�吻v2�%�ƍ�"`3A��y'�;�3h'�����˩l� ��6M��.���>�[6v�}���A���$]2i�������s�U��Q\�P2��gR~�^Ʌ��[�G����f2�i���8�kXBM����[��G�����m�f��M#�5C��|�^��\�I0�M� /J�G��"����^�=�]�i	�I��t�"��Τ�B{����	-�x|��|{	�X`�}m�Њu��;|�c9��� ��
2 ��e#Rc(�j8�[F�}�x0L�-!ǉ6<W�M��\����`N���H|�	����]�ܮ3��1>+�/�Q�!���i]]�Ltw�[��t�&B���G�459 �%O��)Y�T�z��5��u&�^J]����O�=6
��w?6�r��34f 2�7����Y&�l��_��.1�`D����e~�u:}ȍ�4tC�9]�숌��ɟ4X/� xS;v˒�i5��_�-����o-�.��iĄ:��j��ӊ������I��Rn����8EXБ��]�iϲI����UI!W�{�8J]k�;��}*D�9�6��i�H�oS�<�5�͘���^;,��f)�'�I�AS0�C�N��B�T��1�s�LMI$2b�*]���f��#����(��8?}���M!�T��^�~P8~Y?�/��!��z@]*}���1����":�i\ ��!a�h���^	����S�Ľ)P�!`y{��/���>�#2�����eRk�v	�u5
V�=�����C�9G��%�vԳ9��\ !�����a�,/���A:c�M�?�<�����j�Ϳ)Y�S�d
,�i���O��f�f׽�Us���<[���k��{ s�$٦��+�y��12?R���xlJ�˦�n+\� I��T�%��|��V��-d��=(,o9��덱	>��/���\6��&�p]r��t�LH]��ƴ/��Q�8K#�r5{
�ɳ�;�,�(��u�����ۮ�WlH�Q	_�ǯh���&�n�pVy�F�St[2���&8��v}��J#i�NNdѾ;}���Qfn*';�Ûd�Qw�Dz�|֝�FA�%�	Z@O��S%�,�$?e��,�0�uL����Ap�@:�jw����>x�]f��Μ�Σ�;OX�kfF�}���$��������2<	�Y�*��$,gEL����aL.�n�R�E�+�A_-'��[��O	�5[�Bs�[��.��7W4�VQ���ꡊ�K#��[x%E��Al,�1b|�mϱq�=`����-3⫊�L���s���{����+�>R��"��W��Y>��3�5FN������ aA0R�\� +���b���Nb�ð�)�E+(%���u�r���n��f��tQ6�A 4L>�1v��"��\��������ΰ�������$��k|o�mܴ��^��l�^o���3��QjY��|*L�c�@w��V�����@dw������c����]����3%���W8�uj�Ǝm�0C�b���i�fcM�p.zVK��ܯf`
{��n�(|���f�\O�pʅ� �'tr�~���9�W�z�o��iA~���~گ�N������(�}+��wk���-y�_Ӗ��	�Hf�/\���5����5��<�)�tǀ��,)ސ�aҊ5����kr�λ����1p�BP��g��+"�6g�
��
�	/,zϦMўD�t	A'1T�
�~����k1�u8v���"9��˔