��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&n!��0��>�h9�N-Fo���Ĳ:��������&z*ON^N�+ͷ,:�:�8�w��������hP����9�֍���eF,م�����}�65 v&ˉD*N�t��ޚ��x����Vn�����;"g�iNq�h6�VA��Μvі�g,$���S[J��-�~�n������Rj�B���E��M�<5��W �2!fk�9�:݂z�<IY�۴YC&@�_�9>�¹+�\�a�g�O`����)�qҞ��8��=o�؆�X�`8)��xu��
�`�D��(N]�{��I����I�6��]���l��T������tr��u>�/�8m�����j�l����Z��姂%Oa��vF�9�O.� Pt�y@5C�=��P<
c�f�|�����ӊ"P��-�U�NUS��:�n1ao�������&��,X��5��H���(	����qK�Q@4K����h�a��)Z/ҞEī��;�]�7t��X��]Y��w�#�W}Nw� ��u�"��0��o�s9�aSWr��WR�F�#lY�ۈ+z��܇$���׹ ��U$�-n؃*/m�خH>����f�M�� s�W�D�(;[���-�K6���;�M�OLVy �z���a��٫{�mV������$x�rE�F�,�٩(�<���<��Co�Τ,�(������p�E��=�Ä��8�҂��R���I�g+%?p���,���0�r�%�9IȂr�����m����
99p/�Lq���6� �c/:�w������|�Uԁ�,��u΋��S��e��4��x����6��À���"o+�8���B�qGbi���*Eo�u�SRS�P���V��j��zH6���_�3�1�֮q;Ľ��S��3�����Dn��H^A������W������`��un�����)T�r\��d�pN�Th=�����(W��\��+V#Q���v���F�q8r'��D;
j6fn�eo<���8l�,g��U��ȓ5_�L��>YC#��65���v(�u�w�;%~·l��ϺN"��R��ʬ�%,h��ar��CN���e2� �H[V�����Bws�+�q0=�6�>W \P�ި��?���L9K��R��[�gz�ɦ���N
��!s>K���*��P%�kH��=���[�X�Q�m>(�^ƭBo�l�H��ݞ�B6�Y�~C��YH4�+?Т�ᴷ��@�-Cye�\b�����[_w�OZDƧ؄>\����^�7��HM'^I1^��ؕ�Ug���ϾR��	��(^���p�1U��.�L��t޻wœ�B����2�6��QGY�mc��7��x�h�!���v������' �Ɗn+��Q�֮U� ��WwT٭n�:b9���0��L ��������|�U���5p�ΐ���+�jz��4R�Y5�_Σ��'��mS���>C.�C��U��u�0g�������C����A��y2�
�t~1R�`%��ͩ��S\w����eX��=�7d���2:m��+*r~�N�/t���凪ͣ����	��a <V��F�wo������G(x���������@@/;������Z|���K�v� W(�9W���$��ddC�:XS;��D=�?�E��L���+�����L�o���ЎC�aܞ�
��z
2
�`A��	<a�+Z�@��l�viŅQ+��z�9 �P�i�l`�+��-����\�T�E��#����ymE�A���K�U� ��x���ueyKWN�]�fv��#�m����Ί�i`��wlNV~lǧeC�0��y�O]���36�p�"�s
��R�EQ.��t�� �g@���ddo����l�{5�(�ѬD�H�sHw���E���#�z���?.�E�,����̲��xW���ֿX�4:�_vl�5��`E��8��@
��V��=M7]�)<$� �m�P�xvlJ�1�N�e��c������ӋᚷV3��昜#IR�S�{U�+U(���6P?!4����?v��8�.��<����NT77�p��o��yb����8 ���Gs�
�80u���me+~�-�_�d�A�����To�	ɩ���<���r=�q�^MR��/�e	<�)��������S�s�hV�ݷ-���M��zlU����|�":�
��N+Mڰ�f�ƥ�_ۅ+|A:U�fȿ���5��T�;��(iD,fH��ػ�lbf��������t�|�̞��g,=:�`���A��R[�0Q�8�,��K'�]� ��� ��3TٚW�e�+ᾦ$�M�q*pX?0��Ԟz�|��I�i���̱s��$3�Ik2������0����"����Z�5]pך�f�h�~�X���u�:G��7���z|z��ָ����-��B<�+r��`���ƙ;ӛ����MN�ﺺ@���I�W��N�B%J��6y�&���Tm�fyz6�7	a����K�j.?��Ր��	�-�\C��4#���f�E�v@�|n��P��~ev]��H����Y؁^1�R}tR��z����p��	�����x�~GvY�g��I�����c�!$
䆚10��|/�� 9s��g�f3+t�e��0!V�O�x��Q�+8��-���U�V	� �/>CqPSV�u~���?�gQf��
r �D8$���m��GR��n�vV���%�3�2�/@ǝ�D�2ӈ�5�C������@�묝�\�t0:��K�vNOT,��u��fm��8�Ԓc���F�!ᕳ���m���o�f~}�afy��>��nx7�Uƒ���Wp����sm%CnesI'ԗ�&�	ˊ�k������	^��d���Q2,!{�iQ�Y�N����0��y�)�w��4�i���O~�5MR��E˸�Vu���P���2��Ew}�j#7�:):��2�	7Gu�Wg�|[�57���i]��rWM/9SH]�, JӤ�"N���Ѥb��z[����/{��XF����7�>�u	�z"�'P�������1�D>�^���kV+<�2�N:e�*�+��TPx��"��!�M4p��w���BvUP0=�f!��2r�����Q�4�U��:J�79>^���)��FH���7r�j���C@	�%�ٛs))]p�����faޜ�Y8rL��7=[2�`3���VfE��/���'Ȭ���m�?�H5������ʶ9�ަ���/l> [kmn�C�{!�*���-�_m�@J��ʏ����k��u�UĿUk�70q�N��J.쒞��ev0��'�{ϊa������(�~����e=�<d��]��3�V�ĩɫ1�ˈ{6(.�Y}/�m�T&��P�ލ�ʹ����4dc�6�ap�P�N}N�D����eu$�5I�Έ���<�t��%�ng,�a�x�����#���r�;D(�{&>A�I{���� -ܥ&ƈk!QXn�1��#��y�"�"<wD��[�::ŭ<SU5�:whÓ"����S&#�D�hus/(�S/��x��[\�U�i�2�UWwO�CΔ���=.�4�5,�G�q`ᒝ"���&�jn�PK��*����?��1���4=X�#�xҔ��v�*���(h�pEz�3H��p�lm��W��c]�(�cۗTRk���8LJ)V9x^�����4"��I#�W��q��a�;�䫤�cc��J��L�\���_���s�� h�su�
K��X��[���6��,�p�h��{'k���_�D��W�2# �n �����55�ѫ?�>Xְ�^��҈쏳x���r�����>"�c�ޗ�𕋹����4��|3~��kՓh�	Vx�`s�mSI�r�pY��U%Q��f_i���d����m6��e?��NQ!�3bJ�r��\>���:yJc9��Ҝ��j):Z�y����nX	�2r=w�u���U�Q�t]��ž�;
�xMʭb0I��@�|A]7�ɭpO�kS���l�q�k���!���aO�嚏̱9�衂L�z�Ax�����T��'��U3�zC�-#�n7�X�(��h��M4���O�X�C�2r��+�)'�O�a����ݤ+�#�w�`�oɍ����7�i��i#D)s��P���}��D�B�������5W X"w� F���C�U�"���qP|�s#��nz/+�:e�%;�%��G$���I�af���4k�-'�wE��1\>������h-�bT^t�Jw�a6�p���Vk=�.T<�虍Ý=�5t��Fq@���4���'����sʕ��V�8�ko<���
���X(7�}�|�f���(���gͫօ�ѾF��f����Q=O��d��$K�1�a�m�u<�SDv��Rݲ]�@C���E�!����@.ә琻uލ�f�#��B��;�`2A��*�m/�]elb�����dVO/����;�5_k����\{h_|�iPW�Dm��G$t����it��ҕ2����ZE�x
��A
=2�ޖD���}�Q�C�s�-hZ�;1�ݾS$���I�� D�QG�!T����/��� ���.&��_��[�-:�Z���]����:C�;W�(���iH:@����x��#`Y4K9#:�s�L���(غ��!���%5�mV��4��n`�$���8�%����#3\\7k���.Q���I��e�A{)�)�����S��k���<'1�er�sa���%Yw������<�-����=��g�c�ڋ��.,{�&Ld=7Hq9�R�N$�B}F�R��zi�pZ�|���e�F�I!��1���K��P%`�
m.qN�����l�L,L�ӆd��c�{�#U:�]()�!���Ye��(S.Vbt�EAu�t�׶�����5wƙ"
*&]6��P�Ҿ�p\L�t��1m͙R8aR�-��-!��&4��f�[���j�H��}Ĺ�S��Zٻ	��t1[���3z|`�V�ݚ�},a����ϲS�hp�*1�C����&��\��NLq%�W~�ׄPi�R?�ϛ4�5�o��]� �2�����V9lGX<��)���l2WKۉ�!2�ٟ���@Wj#Zq ��VP
���:���J�Jm�n�����&b[�cC �ڛL�9���i��@Q�:$F����4޾��!)$\X��'Г���c ���xy���BI����S��.(�^#��wND�P���c��j�I���4��d����p��7\��4�#����hð�s�v���\҂�S����p&���s��|�[ ��32��	�O