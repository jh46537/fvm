��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a�
�Ys����'Gc�$��@	[��%�ײ�Q�tZ g��xK��J�H	E��J݂��}ݗ��e<8N<���cա��b W�t�f�f�(COE=�(D��sU��G��+Z�D#�ڠ�U�Ӌ�q����X�5r����^��'�M�}?i�:���)Z,?<f���?�y�Ҥ������,�c�	�r�EV�$e�j�U��_壬�R8V��
����Bᐊ�jkӷ|��Ť��Z��mcsZ�a��9@��)LM��������B_��TG%`�q7����AT���;�
����Jr"��@�a eI3@�&[d����Yؠ5l���-O����m�܄���&9I��P"�������|�g!f*G��6h�,�Bl���h@Lyr��(M`x�%��ٿ۰O�VՆ_S��a^�+Y7���lw�	��iL�O���w��eA��x�0��^ah/N����RKIL�V�#XpT�}^��Uq[����7��bu0c�C�A'm����Z��(Djx8�k{�ӟ�"�]V��N��]�}L�1�M�͋M�p�~�q^���V�4�P?w�+.C���P)��@�}L+)�z!3�t��n"���=�DF��B/�H�Ϛ3�:I����(�u/�ސ+֋Z�>bW`:ZDF'����2_&����V��R\�e��D�TcK/&f���$Ys��|,w�����vCGMm����9��>�Y+��ӈ���u!w��z�X��:�[Ky$Re�ۿp?*�kj�<����ӣX�WXk�\�짲ᛧg߹y@��';��%�����[{�VfL�ay��n,̈~�.y-)�t(�����H�������(����2[�o��5ŀ�$'�	bFrk�&����P��?/Mr`�X0�з!���)�2*��К��٭	���E��^�|��!]& ��U'�������7�� ��~2b��I�m<,'Z�D&ЁO�����b�?�"K(`[��N���l�-���f'ߚ[��#x�7�f�9{$��f^���DD����%0��F�yz�a-G��^�w������z���%��9hNBojr�l����b���d	l%vT�@�#m������%;}DO��47s���i���
�e�(�)x��:K�.[]��
�#�0s���l+Gr=Q�X㽒�'%ΛJ�
U��>�Lo��"��.JǴ]���l(��4Jj����J�Bp3��>���T���9�)�Y���S�@Ȃ�3���Ϧ&�
썱�ۚl� S�nG��]8�^0�W{R�c�����н�@Ɠ�M����5���@U�gY2z\^ܩ�{����]xI�����3��0�r���X�4�=?%����B|���Z�&M��Ն�~1���8"��9,H��G��n�d���jXQ���r�ڲ�w����{��|He�%ޔ���#��'�1�Kx�D���:$$�MzOa�n�2�d1�y�;	�dw�z�=����U��գ8�����Im1��&r�8�K%Xs9�1�P�[�X��m+�jx�j#���d��%�w�@��,��A�M\R��R\h��\�3U�����vHQ^?�0:��s��_ V�\U��j8�!گz6#a��o�j��g��[��}�-��M�]�t�U�L�2�̃�X "a)��N�-�e�whH�Ե��aY,��,au�{_0XX5-��A�o+mE��-��q����R��CBޭ� ���^��Z=�do���^��Xg�3ݖ����U�V��_����d@��Mtu�H�|,	�հ�W�5����̈́�~C�ww���b͐��_���j"����pѓ��̀D�c-�>�`6bh]}V}��1�b���W�k�	�fӦ�:��u�������M�Kw�*��0�g`��$���	4A��& F|�E2m���wz�0n����}�;slX���}�^s�	?�������m��PsU��9 ��D�w(̄��c�	��-�`��_A�o��`�v��K��Z�P�n�}�Օ��*T�*����v���b�g׵�K/�),�d�I�M>Y��Jp���|��I?��)�ܔ����������=�HmnP����i?o�ROn�dL�N�FV4u��a2���&�S,6��C�	[2]�r�����uyX���c"��*)3��1֏�%,8�))�SN)��^�G�X �1��Fڜ3�|��!�)+6n���;��]3=�iNP�����狤gg�Q��@ru��R�����pTw��XgG�Űɒ��È���d�n�;�����>u�l�CrDj�QA�У�Ӏ ��4����IC�7\��)U��R4��%����YΫ��5�G_�X�L�=+B���|��0-ݏ���W����Jr���G��w�ƚfh��A�g+��BGe�E��%����Z� �r�u�{��"����Z&�rmp~�ݐǽM�^G�X�R
`m�[�ot=���i��飜������{喧hP[]��Ʌ�}�#+����(#g���Z3��z-��Ԙ�3� Gá6a��	���7R�{W$�� ���y�e-j�.1��0]K����3�ؔ�R���zjKQ�<Id�_����bwR�+m�O���d��TQa��t�;!W�?fǁ-��"�$����ˆ�?���E�~��ID�ͣotRP-�!k~��?�cEH�}<'���4�v*����h/���X����pѭ8�5�>����Ǘ\/���.�J�5��r�z��g�
�0���,�G�m@�w���G�Z�c;�E4%�`�p�����p�.�r�菋{�5�tq�t��u�I�+��\�;�e�KӤS-B�I�7݅#� �_߱zN��u��t����AJZ0rl��~�9_�n-��.�C�#��=IP�:�s
�%��^���s�
/B.�0���9�^\��e�(A�lp�Q�5���㙬��Q��������BY���R��~������董�g��3|�d� ]TsE.��ٙ1Ϭ����:�e�@ s,T���1A�U��r��Io�i��&�+"D+h��X�� 5n��k>��$�=��¤Eh�M2��[�<�r���mg�����-���/݉��rKE	���W]p�T�\t.���^	��yl��8��r�������$QyL.�2�L܄���3�p�U�K�fZJ.sv���F.$���b��F.�ǋ�sW�6�6<�{��El�����.w�dU��bC��:T|� .�����98��f[6�L������(�ۇu�.���,!V3Ml�߉�i�fjҭ���d�@̈́UZ����4��a�.t�!�n����q;!6e��F&T'�B4�Hnj��o��Es��k�-}�3~-�����00%�k��H�V�[�RD���!��>�ģ�brLD�.���%	���J�?��w'��W�yL��������YWKk����`��Z��@�I�S����-�@�N���j��5�ch��޿���.����;��pz��> 'r\�mrx�C�����}^��TIF���9�!��z���9�ழ�^�����4�'~�l�`�����l`rW��[j(8E!���-�j�+	O�VI�J�#��	j���mT΄nǟTίdN�`�[�=�y��Z�L\H�o<�dc��1w7>��7�Y��g��]q�łi{��0`)��[�'kk�䑘��3X������l'D��}�~13x`4?dwdܵMj���}�����`���*ZQ�$5���M}ȭ�*L8-O�c{}�֊gͥ�n�k��C돜1�f6���4b:~�}D.8(��I�'������[�&�\Lf�{��o`��k��[\:�Ǡ4�=�#������KH�g������E�����E�F�t�ǔ��4O�W-�fbC���o}�]2�x�-�y�������������t��!�Ć �����9h�,"�˯ "�Ǽ.�q�M�G�5'�N�A��>wQ=�볡��	����s��c���|�C-�/~+����k��Tr{�
i��*�c&q�$O��#�4t������pa)''��(4��d�Qg�ZRz�p�������I'��h��U�5���r�3�o��.,aM��k�ܲ�}Ν k<t��K@��ۺ��5�@)b�jG��^�︽@Ի-Jmn�R���վ�G���b�gd���i�������(��Y�1���|�ٖ��7@��P���cڪBU�����l%%V
6��ظXi6�b����b��]θ�hi��O���H&Y��D-��)MI��4o^s�9t�bn��P���l�I�[zhJ�⡮e�?�d�Xr�\�+�c5�48OA7�_��N՘v��~8�=PZ���+��`�2/̒���Zu����,��U~^�⽱�������VMI�7V�p��y��c�;�eև��(Bў���΄T���GѶ���dYU�V=pPPZ�N�a���gQC��ߩ�m�`k$�8�m�f�㓗)�FN�ŵ32=x�>C�3�ȵ�Ŵ��N�F% D[�Ts�R�cO�:��ҡ���P�@����EQG�z	RI�툭��Ŵ�TF�s|H��َ:2!|]Ǎa1 0�u��c`�s7hG�)�]����Jp�f����b�a�Pm��b��7f�:�C;�4mq$S�GO9�K�~����e�IFO� j����ql�j�'�!Q��J��}�]L��FY�"\�I6�π_z�,|�܁�m�=��T��
�i���>y����r:< ���"�d���)�f�!#[�e��_�+�b�و+�W9.�a�/:ge�^�����(pN[�����;H��b*5�3��rTϪ#+�-��y�*�U�:��*�⶜1�35��1�C��u��qr�WZ�d�H�p�TQ%��u�U:�1r�B(]3㚙�
�֘6���~�m���"��d�FnX���`�";6�8��s��i����b(�l)��-
�N�D�����<������e(�s�.k��:�y���摷�������L�&J�?�闚8�pn��}�Xկ$Z̩�=� �>^��a�{�1 �+l�#�'��b�G~�BW�Q�A �⛏�ɽ���Se^<b{�N[ԉ6��LI,/!I7,�v�W0,�� ���[+��*)'.ՖkA��/�9A���f^fc�:ae]�P�P(��b�-�4(�%C�{����@�����=��^Q3�2 <�f�)��Ά`�2.,��_P���p��8��V9"���)���d���8���m��+I��x��d�t���e�3ocn ���rV@q�5���K��+��;g��r ���� ��5��Oșc�'F=0�F̻H��P�eoSC��8�*e�0Gw����nZ)�*eܥ/qRF�1b͏ ��$�J��-ƫ��<iHI-���TcuX4�\�UZ�㹤<����+�a�J�j9����K��~kӾtJQ�0�z<��2P9M��C�[�����,v41�
M~���[a#��u��g�d�=�ݸUD��<$�J$��
&{����U��z�G\2f?E!�&.K��{����}Ƹ?�䠞��R	���yk.���Uf�JJbٸ�WNض�z�Y!M����XA���D���e�r�T�q�1 �O�#��L�L�R$�f��TH�6�ә5)A�[�l�a2��e��������	������VL5�o:o���إ;S�lV�,�Ͽ�wJO	�>�1��ys&<���g����X*���%Y�v�yv�AY�NU�0_53�@,g��h����	&�]���*����F������1%�V5�&N�T��%��~�w1��<Q�-�7�W�d�A(��۟�S��a��WBZ��ԵO�m�}m���w�qR��#a[����w�j߮�Fc�OA��L��I&=��`ꜷ6�.[at���`|���q�t��q�>C���6��ź]Z3.��nԾ��d�4�[`f{�^�̡��>���P` �a=H>`sy��\R�A�|Te񳕕e�� ��G�À���JX0�NN5��!��	���(����~�z��/ M��ٝG\RK���p��$�$�љm7��d�d�N���7.��vλͥ|7�1=J؁�C�F_���Y3ǈ,'�3��IgN�6��$�����p��R�Z+�
˲|zc �xZ�/(Ү3����� ���9��Ʊ8Z�1�r8�W��Ue*r~m�,���w[ Ƙ���e!c��U��̢�!9X�겫D�����S��T��i���zp?��o���^�D.�07��iu"��TO0,�4@@�d��Kq��e	��P}HT�K�AoY���m0��*�Ġ5x���</+Vή��.v��c��^����S#>�{���D��@+��y��X�Ԑc������yo�.��9���Q�wj��kU��@ҝ6�Ҷ�W���;3/
���_Jc"�WJ��q'
������ALk �ϱ k�5!.�犵�Z�X�%n�5�I�'���(�_����G�З�f)E �����@�D�jw�VM�����r�)��|ZeȞ?.���\�F��s��=3� ���v�ޱ��~wm_�u~d�+�n��MQ�bݓ9F���bI��2%�Ս"Ֆ��K��9�eXBu݆E�t�ɒ����