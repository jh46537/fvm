// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GysNz7X4RZJby7H3iwVDyGkgiv7nVWGCS9e2Q3pDtZ/2ggtsIesGQ/MBLAuSZX6o
aJC3b+UrnuV0nLgI3UYbM016nCgpjQJ+ZPUYjxZvt0kuC+rNzHVzg2gkZDsEaA3n
pmzDjDa0LZcFCyxwoa+VATTH2OXNEBmoiafYhmJnSYg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29216)
t8S4xz/lf7zvVkl/i0Wfw9WqbPo/t6trqYE0R/m34FqGmUDJWLLWgdDAe3G5hwjx
ZvRqBn6Bqd8z2hoBW4M7qL8RF7u3HFs4WeJSAHhq1CHmM/siHfu8WgFvJr23J072
CWpgPJ4ythy9ky5jjlV8kWMqep53PCi3mw682vEbHarqJRf6O+Sz0LpWeiDW00M6
+bLtrKfvIS37fm5c1p2rGX1FfRqQS5pPQ54HkWiNhnimj3u0hFRZbHPzTbbQWN9f
62icOcYjqF2VmpM4LZ1HOYwwFHVqM8FlZ95E48HlUkmoeb1opoFbMmoe2kmQ2sI7
KzuCyE353XqeirbQyMMDm703fyuu4skgmwsNQPHjVzIgzJGecbtKgwU9VCPkkSg/
IsdkPSaX7x8AZJ9WKz+E0b2GGE+YcBoD01aXV6oCMUHSqU97CJ7B3FQjORGMXY/N
74AFR7meR3Gb9H1G8g8McGfyCqPzRLVo3pH4Vg8sEOBggbgV/qSlmDPOW/YAXh1I
sgkBeH+qH+Rv56ryikmvOCFa1TAWJIBQM0e8v4tJhMNfk9bGe7ZPmPxSrDC26ZQN
MHsE/WmR71Pmh/TCfvkguvx1UQ/LIDM/EplpSHLp/dB3DPCSCmTz5+q5WR4JFnn2
USpthtb6OsAWiZf6WVTVnNOmkAcLUrS4TGHQlx3URKBW1jONSJwNy3vthhMhheqF
/D+EkrP7Ota3VrwPJCl7sxy3ZLFVc7t1drwWQp7QgYhdDVg2hDheXf/4UdSdNDFJ
eroT10aKqw7VgOI9H+aTuaJHGYDUbBNk8LLYyOC1DQLoH6eevRiGKoFhm6m0RYwQ
8X/RvMD2AbvNMBBxBJg+uyNoVxfz/Clq3lsM9O0xPr94ctIZyDRZzj9UednhX6D0
RK7BR+F6/y0JpKqzk9+DwVnStlBueDghbo769+g1nTRkpPN/DIMX5kDhDqOCyV4j
TMahY4E7ZqBDCSgV2+I2F8rW8gwWRmVLt2iMVWpYf9HtnkfsImc4CM6AaLq2N8G0
wwQ+6h41BeQVnGSB2rQNur874Mm5HNOqFomcWJ+SLBCRkMmaaQhVhW/WxnSpd6ni
8OKhxKasafqvj1jbukXaLZSJhTBPF1gmon5fp1NCDTpyI0aTZvfJIJhJBWu2bYKE
66kFrEUprRx7rd36CYl4W2lXdxjDz2L3MNZpFfYRXnLxDyFNb2UD5IwuoCRjUwXx
Afi3IwsSU/NMpoHPNb6nvW8IIcDZ1oBiPARovTI8jHXeRQMPQ6yA7qJhM8D3DFBQ
aZ8t7EELlGmLei3UAQMQOGlY+vzAlbfUrRC+oxgwpdRqbQAxoivlKlHMxpO/YK5Y
bJuNgu/i3jFv/YiKCAgxof7uLb/XRIOqKv2AgoVHhjHW9HRExjhUX2YHee6p3jYW
/ouwbJVyVN58TKwg65O3xCe9nEd+nSjwU2h9kNQymIEvw8aGA2IKTD1epx8q3uM0
l8uoO8F+UFn/stY6dAxIGVK6DKKCJZ/ZlfDpAzSdDRhjKBalnBqbox9+n1DVLXuY
cGeQYB8tbTW8yoSJBrWNakAGfjFCiYXTDPI1r6yRTFNVWzkHGycIIDsqi9bqpE3w
IjC3FIlZjz4qv91TZTRS3XwPrDZPeSpKHbTDwz230/7KxK6He3TagD8fwrjXgFTu
MX6ln7+NJitV7tnyQ3AbwduTcxlASI2k474MNnbSCz2b4XnnEUZS8HQP4L1gOVF5
p7qn+xwVyAHCue/u31PdNnjdEm4pWR06doOlZDHMhXmPbLR4e4h/dIGhk5ZI4ZfL
coFrh0xTakYgkqeXX8r7XspVtvwCTFgTT6R6+lSEJxU5pu37ftB7gsEm7NXibtkN
pDw6v3P+9V0cNKh4trbjpa3AWNSYtCuvIQyhdWrrNzRdqzhWbFTX7d9zdFdRklct
tK8CFLR+r3bpef0OFSwwI5nkYXrUEqXe8xJJf2eakf3SvjkIa8LIoKlrc+0yR2mg
urdMeQcRHiwiou55Y3jPEEh7iuI23yYQvzh+hoF7pURbwKF0O7HE1dB8W5op8FuE
K+0W6BD7HSqF4x21v5M1/PF5J62kritC3/QfLvPx6z0751B3CjC6xLyqOemYb/fz
KLTQVRt0z6NMYomvoZ+RrC8E8heLZtFyNAKccLnuxMxNOILJa7JARKHZ9XyKHeB2
2puooAXPw6CZTJT7enZ6LEnXYRhCTptBSvdYE6GA1J6wr1KM7oVuw4rsnaR4DT3Y
O5s7EKjkAi0OzBTZ9agrrhVfEEsH55S8FKEKkdtBZBmdpOmODZApKdy77uBWBtRS
NCxCJgvPIo7uOsor/PnRZk7KE+lN6X6WT8gs1pQcl+WL/vIJh3zfsaUYOPYzwQWU
dQcnbqZ9F9OE0a8pub8ljSI1DHVyXmLhaaqaspkoctlF3jXKqXZk9jchK+5Hk0W6
CP0NjMmKG20zXGvn0i+PePzKG2VBkwr4t7KAVJua9imiRpeeg593UKtfmjDo98vY
PPvepcv/fN7J6grmz7v0XLRj/huv1icmtzFET65AFqVcrdXyILqF6+RSQZJTks1D
7IoNrY4kapIu3NvULU9AYZP74cbfDReVAIn67I71g3pum7kyVhH0QVUKVa1gcWnD
Fp7fZEV2N1R/mPqdhdjXc5jeS8hT0Zg0FvsH3NihQOZ3UukaP+WaJ+TbhfiN6tri
0y0DJ55FTj8IOdetvxe9h8XxWY+Z1vfyHsIZdli6don4QYCnHPus4iWwq9/nocw7
eZD1BP57mh0KOMzsruS4HUQcYqmalVBeY75XKbaY6b2itRGaxfEvaS6YtWTQB0u5
qmLQp3EqfHpjM8RAFsAdS/NFYwCAc7HEbLcYwxGRJgd0dpRqWY8HOzjeag8fhsR0
O/2GqSR87152uym2FwJ80RPktstfsu37KglfUvDt3CX3+vU2l+UwHwHEvdfgunne
mP1BG6zsjsQznoMaiQsZaC1oDuSOEMG0izvDUtvbQQ2flVFSntRIUfvpDsuULECL
lMtpGgS3uNnbKu9Mn7BjmNBNZCHuzyFp4jdOF5Kd6z5cuNH6YygHIwciO+OCxPFh
NIzyTc69q0r8R6VGwGIQrvk2l4PgD0O5pstlBlWozabzjAveeLRD2lVWFKcoIUwb
+CwpTFgn8tY7EvS5yH7TwRghTBohsmmhaFzvoxBO1JyLlxgKHcyL/oViI1woms7D
2DAnLSoI8Nxt6KhsfPgXKnsVbN6TI5BTVJT5hTyjFU4s/iEyU5VRiQVq6+sp4GLc
+VMIM9o+B7AzmZhvMsR8VSyrS1zRl4zYnFY98E6JMairxYiFH2x+YnQIeGi9ijXU
DkBWhhzXBv7fWjKFCLD6luSUx/c0P63b72KdZ2xNh6O72vazEKS233rhy6iikNw7
o4DCVSw7hUKAEXwLjzPxmK2u86o2sVll47hwKLnFs3mialV+oh7msylMtcp+zz9C
yK+i9qsn4zZ7JQWjMsqyyZiHQbmV3UgihIFl3UwTM0iYa8/U6bP0s3IJ9g0dc+Cm
SLfjfBaPJjgb+/LzxKu9ChgPKc1YRwwgvnIO2bMP9TFdPEXFDTgPXNRqbjAc1Jtv
AHuEtfuq1LsrHW34bhh1rJxRb6E+0nMQT4paKjClzbqtYkABX5uyxq2DQRNYrqMG
Um5n57UqZ/rahp7LAqcrygCjMEcZHjnwpC+4/hw393nCzF4JNZxRCyFtnOO7RAY1
ijbZWDSWK3kHEj58DTk7apMBJ8yJTGiAXU+4ubxrKelAOdopwGA72JUM93Dm31jt
mepPdki8WwLy/bBagul0u7bS4X84Rt+E7BH51snWdoODL8OLB5nudSnfCN036Zu4
PGvB2En7lflLjZf7l5xxkvI8A1uAfVakelNabZd6Md8kkKpe9VULxqGJNnkcYTZj
qDT9OxtWDgi1gKxJrcN4BOpW5J7nJE5lAyjjxUAgX4sUVUb//NLaiHuoylH8UU+Z
gUgqM4ifI0sQvmeCFZX6OdLUx2yCrBomi2f0e5iGJIbhL8G0GeQLHxNIaSdxT3O0
rqF3DYCJegeUTKVOft+AtIywHRhJp4meNkIBo15HaaN8EW36geV++VWA8T5lw7Oq
amjWAxQePVTCahqS/4GkFoKCWDYdw6hIiCLN7XLXFDGv8g2ZcYxm1Ru6ImQgmqtJ
o6VDJFhaI0vHkW7hOeRez5P/zSrR3rwseb19hr9LjWSsxT4xkb2ajKcWYbs/qGih
IOOybYlfkUgve2/WFfYOQFOR6scC29GmmoqIAG2CnTt1xmLLj8SN5Ir1oRVGL5DA
D9SGh0Hsp6znwlKLG8UsTtr1geRAfX+hieSqALXQkIsyMakd4SQBWceMZb23cf5I
emwKhk7VubR7/Q4Sg5y1yCd5MToD3896qE7Kw/dB9KNDxHcfTKeEpGrF9ycsoK9D
nLGHhsniRM9bJQN/jf0id8uMJWpdyK1Oo7IPF5Jm9SCWQtNHTVTP2AhJ758fpmvr
kCZDEfjxIDnjJB7YAgEFZ0mow0lFQN9t4zerXnW1Jvk+Jm9XDxCgmf3KnfxcxZDs
mOJtrRfsrsrURzaUrTz7p9++vcVaVyqaslQtfU9JCcnl+a17yXCINkFy+bqjxkwq
VkdleUHWXx8HoZcSLqK7bZ5UxVMk5xyuPkiEGfCFpb1rrwfbsTaIdtncSbx+MiA6
HOxzNYIu33Q9unhQ1gAB3GoSm/3aSD0eGbd4ykLwFCU27LWu5ND07Jd+oaoJOL5S
Qnb6uea7xR/UVuF6X+ILPh/62TC1ggE938jgjvcAvSzYcL9Oh/3RDzJsJOq7OCF2
zvJFkJ45d8zDqrkfOzAXslXH4PqGVuquxPSnp7J0gSd8Tr90JVC9lXkdByGWifiB
l/JyvlEVmS4KvLy5OUOnLx3VDUREtEXCqte8IKqCIxYk2qHOU1u7oz5KOfMsBp3T
Ie//vipZy4Dg/y4iB+skPsUp4s9tnxMhg5pe6tFRcWG7UWHP2cKKyU6FsFUshLmU
KyYeN9TdfSzBKw8h/5ltyQATKaUQBNEgnK5SFQcTZ1tTix3NE3f4scUdssdXZnWl
O9sYUFS0uMS+7VUqxtqlQ4xMGtgfl+fXlhJya563Vh7jI2E3jjQWkFe4meqLCMi7
N5hbnyDBVy0lQrCcvZzqxEaOZnzupMjMXQPQTIlXYCxFtNl2mn8cachiqaUhv++U
xNOYyXSD0m3MUNrc7fJRkmCmeDGMNtdusQ/4BpQ1Zpcnw6VRGNZtxcmI8jtpaTbt
bHz4sH/A/yg/hhaRkioMqabzIRcGWwS1gDZuU+UeJ8d4xzgjVEz/LEZD7M/y3yua
QJjGbFG0Zd4S/FwTq6OOdWW1Rz44TAdguh1m0yGnxAXsxLnNmy8FMrx8hY1i+jQw
ImGsGSBj0TcW1Z4upCoM8lFBb8PTXrYf96yInmgoP2xt74lOSVMgB/ohfnfq5Lpu
C5d7LGW3ju+T+l7LVClk63h5iPtW8QNazsxlE0+vWHJMYCwZM2lqjzXzjp6rV/mM
Zmy5YEHBa3m2t/wMMWIO52eKoOGjiMlx907Zzr1iXu8aDoGj0Sl7ziPRzF4IBNG+
q+NRb+lX03V/APXKKl0uq/SCFIMFP3BzeRc8+FuKuWixBS/T2SNTquoDm3GsmrKH
ZSYnU28+l/ECqiRfxc936bm8vMCeucZcV0jtOHLaTQkDVCUPpL805cfdjRWxCBhd
NXSqPNv0VxQqZaFAFbSIV366pcoa4IoOztQH1KbuqUsIpZeFMNPTjBQ/DFhrlYPu
t5WGUaxfSrXT8gAxVEAAXkYZEJ1k98X9z3C6+16pPT+Jv1twQowo6t2ePebzJAa1
r4KHBWVqK5ezr3SLv66H9oPW1agkOHMspzCmup8chVO4QbgCtprO667W9RignH2k
AI8GCL3rPklmRS7OB7vCSZ0roalP+w5gdAN2oyEkIZ0gB2ePSZ14caITL6fsn9KX
puHm9fmNQ6dh3HbbzabILiIp5CjlMFTMYoR3jfNzyAFe2ZbUNFusWhdqhkJmlgQG
WMtlk+jg3QU9Qw2//xGG2MuzPZ3wZ90WTtrrsgu7Wt3xIpEloyxCAu5FNpr/nJ/l
Ks0sgvFxzCJ8yLcsSbyIUF9wamXuf1DYmpUZUT4HwfoeGS54ffSeuoaNhT+2DQst
KpIB5aW2PdS5G1bFo/oJGJsl1JQzhHovatpELRrzUSP6YElkvRsZ+nvXNxXyp8Q1
ui9ouOdzgWDQXu0GPuloo2pCs4BPqy6HbEVuz+MXnFXpc+7VNOdabH1K6wgA13ym
93W5hYrGBnPUhq7SGMsNHanklobyYPubkKrYOD9H769zh/LJ62s+7rC7EVqnYBFK
kdyYI/1R5gv+fW41qtFj2tRwAlYHrohImQBN5S0htPk594OmzryEDJV43zi6L4xo
K9yEBKVuXqiBYoGje7IdIfqmYKZ9yWmFUa2KesrCyQdYjLW7sKjy3KXeWi1o59lQ
KERbBNKto8WN8TzyxzE6zYmTNS22QbkMFujxopAQ0NOJ/bzQwzgbM24veE8kVLwX
UIBo0SjkemNjBOD0sNjx74YjvLXFeGYEjeVjMGotO2lEqijTQhV3nXXCB+Owjua+
YUHhx086biSjkIE1Vbz7A18ZJz8fZyI9hkzN4zlAGBIMnxiurkKcG3foRiPu1z7Y
i/U6dplk0yWRO01m59iTQZOxCvjkp1laS3Xiltqtwp2sZir7Dde6vOMlKkfxhakw
52v+hlY3HcCGdZkdOrhZEx8Aja8p1o8kMvypah6AwFrtlA9DK4Dk+ivaFOh80zIE
O5te+BfdmWn2e/gRHpKhmni+xMNZjqMA6SC3bkzE4hzNO9F4qJzfzLgbRnDGsgr1
hbLzwaRxZLzZ0TuXXR2oeT22M0VzwSqU0xnbjck2Za/W++9JYjBYzpwTqX9hiUpi
9bQE0anqDLKYntz8IZzy+n2cIG6CXrtevg3Rf8aNFzBewa7fHT/xIVMCAHJI6zyT
aPCr/SRduMVsP0sfr8+8skrSaMx3pa+djMqXCo+DJMJXVmYgp/ECTKzfMmaCeg29
852dx80ZUnqCSFMf4vJh+3b5HXHuGKfS8iXfYvGG4gNiq0G1A87UjF9L6EZRMNJW
KbSTzpg4moVvHtmTeCcleDuxBfVv2qzdezKH0wPb/0gYdvhCXq/SICPwYD61+tPc
C3ji5obaalA8vlmPfl0HRSZ+CfApTfdFmVwlo275a29Z/rWcLhxDOpD/Tjj+Uf2H
iapMUGyY7eApqPBFFeW+VeCVTq38k959tUjjzbp7zXGyAIE+WysgIYEJQBEhLO6i
Q4T4nQPIjF3lVP5q4ehyBOdpbicT5bTowXpVYlNry7zcPNb5dDgdaCzY9N899kh1
WDaHUM5lJ9YQJnaygDBB06YSXXK7+ywDxVZ8OlPtaQADyyeCnTYgKtBiag1/2IDm
5dPslshWzJNBwN1dJWcVG2k8LcgEviAWU/WzALYWrAfYhyBwEzqDgtUcCvUqplM2
1k2z+FMNBjf0tfCrv6MkZcEbywRwl6/5FhPSmbo7AvI8HqQJVHhLSjLNpFW3DTdZ
tt+KeWLkXzeStZrT3TB0pPezjbuOUbEUC0dhzYI2Ib6QzSkAvEFskic2jsY4ZSq9
q7HGkJdJkmk4CrAk6u8e6gSG/XRF8zI6A3fnDylOO+Is5EEf72i2V5EfuBvP8nZY
j5vgKqelb7RzRfoOJhTwguv2Dheiv01NwBMFp3oMS/hs0H12TMFLVEfVLiSIjfZd
9yH933cw5B8i/mFe9IC1mAJ6WBA5d6cxa8UQ68hNg2RaKrv80rC/WEMedf9AK8xr
hKEh/gdwLGqgwZGAhmJX9S8CV3qRy/5vjjh0uszeTxh5g8Iw+8g1cavDdIXdAkIl
71lppiLTH6/ZB00FYfSKgJuV9l4RzGUJqnldLEu4IyHTuBb2G5StutJlubAXoVIT
EeaIVDUuyzmiF5fIwROu5IrNpmtElQsomOwlxXYJ6knXERgtyEGNtHkAP53MDt6m
eaxDCGDV1iyh4sHmml6528EoJJ/heBtcoXVtzrdgD1Eh4kwhqV2GblC7O9XIEgwY
+JNv2EaQm5a8dY4mYgtkw3CSnVzMH0KZYsK/cvDsak3SUVSm49EZo4f491SQj6Oz
LpnGCfLYc7eVNqF90ND0xVBafQ2Ll/kNiK/367Ft0VESDPj0RiMsPWeYR7FW1Fh6
UYlJb/FTJDWiIwg0mVK5pu/rVouUnfgiwGNHlsAMIy2m6MgT7Uz+7G98owmq+esY
dnJg+krsskKsNk6CcsyaqpPrtZImlZJB0Sr72GGsFSQikFd4YkyHJhidQF4zr29L
WEThogiHgJCwq2dcZUyjh7hKVvrP7eeqrypZ2TYQUT4LiSKxhudRETsC0hSHvg1G
HdI0JsMnYqDt3iZc9SGA2JNRYuMPK87VaWy/Q4hOopIiJcOdQKWB9dz6TdcAHoAn
WUqVLD/zpk870n/OcfrcEAKEQFtjMO51P8UCgji5R8zvExy1GLde9j2/UCW0Bh47
KVdF43n2wm+JQcSjrP09GiddiC27U+aCnsHuJjhzbAcTDpkLyj1lT4t6BjDv8FMg
rqTnO7G8JRpmxrAKyklpH47FNrkQkhI7KsXFztY11NBjidOaWn4HHJJZ5X8inQOc
u1yFTksZfFKrv+H/EeVjIdL0BuZfYmFQWrkzQYOLCn9PkKrkoNkBDwIk8Y5msgzf
o5UrhPUWMT92+NSG+skHGUT733pV0x/m9dbcUkRJc+FkrbN8CVA9c2Q2ygYGrmv6
6mf9Rw7PGktR164mtDianj/d3TLU2YQ5KC92yvAw3yLvVjmLHnK4IHSPnBtqUitN
ZY8HV3FByw3IBIjk+BTGlVZQA0MxSNySs/h15H1tVrMgC6HEM616EbTS0XeI0IQl
F3IAlpbWMVzQ4Ne6S4aYKres+nG1dBHvqnCsMbZupIMdVL5QwywRkwTFNVAgkN7r
v2Ic8YQFz78JIlWLkXtV19bOQ+RxEhxT7MIFK9/e4EYuqRJpJFmtrdvthrlmmGBG
Gg6IuPQoqEA//lXA5SPFl1uiStJFSEZVw3kfAf/YsJMNPWSM7AxpSA78ckUBlubf
u4qfQcfOJSGzn8vSduivy1uCY8gLJq5TBhgCuWFjmEb6/7g4ijX4audY+zqWCN5z
kpi8/t3HzW5u9ip9kxTomlp01PC8qX7Qtc8CrAsmqGa7q0nFSFKxrURZBbifPwTV
jLAxybgbQkGDp7BYzjL7twS5kJHXDBr2+mv6OFuoKxm0cY/59rgjdIGPa27809cY
tU3pXj7hJXMLGS4zSFFAEqnjYDGIDpQipgxP3Iwq2IaZ/sCSi8h/zU5ammy3LkQp
FZVN+jXZQbjTQJnJJS+Hsarx7ww86dVAXPuj3uToGMRh0lLBT7iQgDnc4VErIUcx
Q78xvIoaiR2oRN+g9Qktsnn8fvWvahlVP7bNBRWdX1rqe80GOgfApmVTZdHwLQhZ
U/JZnAv+p9qUXxuReDxQ2BRRtiMXVwz9IgsSpMK/1wg3ZVzgEVO2rFUg2+wrsG/9
ugAn84UyN5PfZw1hVPkhpXqfPe8U4HrJUxySzPSEI7VnfPr/KRObpj6db/yk45HP
dYnn6UnrdqArWnkVzRD5wBvqjKW9mkvKwF0wD9mSxZfQ/vxQ11GBmGIdOuYyi+fN
kjjv6duoyTmwI7jcVYQyTFbk8HyfJ3DjzXNT0lalTT3Qa+HO7T+dAWjJc4Ovatt5
XA7FVeWYDXKBRj2bOq34iUkcfrLZJTqKKc0FvPrqvzM37yOMSNdDcUkVLi8dBluD
H+XFJmSqEEKVytZ59sJas8b4Hs3fQMBMNduvbf3edQZTErhgDERHj8jjuHrotXy0
FuKCV1VA1T64AzeuI3i/gcynVp5hBbqXmw97BiDvkFt+KoEIA9SeLBBOLYJGB9rw
208HTM3iy9qN12F4g51iVCd/PoUD8a4pM5iEOU9TldDI59UJqKqEQS73sOSGr6pI
Rh9AjJJhJuOltLiU4/4DnkNz6/fNb+2O26vC/ZMewfZr5t87/PL5zk0AT77TPuCm
Dyxlu3A+eGJJ4mvE+k7meAZV1kHFRYg0xN5dpoJ7lczGkiG/kVVYgg1cIQp0UW1f
hfqbjixJ+uNyV3sKqDE/a0Ccjkptc9HRh1EcwVHa0oCgATJIaHeHScNiz3N62VsC
Tma9BnFyoKZmHmJ6pm6hhzF0Ad0mcMAodI/U6OVWw9gzUkRb/BjlichPXXQkdbtm
IA5Zx01moqjjjPsMyKnJgtNpjMm8EcEqvkBXBdNlyZUGj6gh6oyJpKkBk6yH7TVA
jYJ9lwgH/6D8TIzHzn3vcJwSC7JnBlgzPLemSFKWsLTk9900qAezktHlJvGCF7f+
PeGAWJHk1IEqw86yt0FPG7qUwYpk6EOLfrAahIvhzVdpQqKznRY7JRhSw42VJnLS
Rl1eoyEUnQAk4tBOPfgMRoyAIXorcjABnvWDNrPl34wlcjcpWHLLZ63fcDUv8YYE
AEFlVLCHAK3U0fux6E7kIfy7QOMKJxqP5Y0hsqYatSopEMv/CqXDdSKCEtXPAAUF
1+Bk/96RZM1MJMtfEje5Xo6GOB919CH65DI2BE081fG2kdXlVtGkCs5I1puXbvfq
H+ewBr9KMNQWlEfZ+cI0mM+Tv9uC4bvUvaYOQwVc4g5V6/7Yt/OreO8xPvuYzK+c
CxnKdVx6EfFY5h3UdmdD4+4AZXku4LIemYSmO+l0O/s0h+55T7J3c8NjKa1myNBk
aaPAT849wXeYcCa/CBvyGKkype5bXWlVBfsLnwVbZJ+JLA8ouf0iw9mtxFOOjn+b
BbD4R+r7vZppezBoikMWXfXpdBBmqCq9YzQDQ6zHfv0NWs4Ea3NWgD2rt8QmOpPk
XKUNrpbzyW706A8dAR8B0m5MhSba0+RdFtVegkW0WnHjzWoJAKiakuPniXtBu13+
z7sEBNYXoUlauaoEgQ341N7DSCyjPKsXTIn+SJXQinzGDMhmtRSW3/MIlmtFgQeT
7ayjOHHILfeuwad4G7dhAkKxAxY6FkIQn/GiWvAg42tjebfi156W+FFXB6+/+KKb
1RMrE/n7X7SyzIN23LQ4TbjhNg9o2e6OYGLdyGZBfTWFNvzK99SHyvkziXaUV65g
RyPm8TF1HNKnseXQ/hTpXKLAeh/Xlcjt73TRih5KWhjzAa39AdUnGZe476DT15FD
fL/UjxNwR3D3fpm3uFdnzHtAh9Rn2Fc0gUHuX+BbVWz1aZz725NbuakhNfU3MDOe
QiP5guHrIbQqnKoOONFHrHg/M/tv3vrhWLlfwRXVduSggnHglbBH4eqb8HISgbdR
NsE7VvrW1pHWp1K9K+P4NxtDYkgwgiKR06VjiQOjkkNdmwFJGrluefIn+GInVI1P
v0ALYkpyd9geoQA0oyBwDCBS+KWsWTCcuXY+VzK9WM2tvi1qtuzVuPqujo0l/E6S
HRJlPr2+7r7Wm+55Q1WEfHkyIsEoWzEXeDEZnWJWIk5Gg1tGKyhQrMoMlQBLpu+W
JJO7f63mF9ri2Cdu9MRSiQiuQIH8oeJQOzRSl26G+gosvT+euffyapHWDdAaSHzd
kUpZje56vbBYHfAbZBDjlKDb3DwZmugN+Wp7aiPMcAdvGrga7w0NRZ0cCa1VqUYc
o7JoYrfGoV2vgbjWbVEMBYJBCX6YY3Vd9bvDQvHx1GVNTnwbexVyrx/ZDux5UW7E
gobMBprHeuRK5DbqmfsYT8OYnVhvA3UeZUeecFRVz+uQldJBWS/4xaaKFGWkkMHG
GGqMp5ZpNnqVgru4j+M4x26KdGe/lh6n8XWLIghd+JnGpak8luNJnlL3IZqbX9JU
+iChGyswj+EZqEqbU0qasixXQ0lQocwyjR2R4WKsbMS8HOiJJScp5o1A5ajX/154
ZaoQaSV4sQXlcUH61Thztx9qFa3BwqqyB4DDiA/qS6TgpUmTo6Aa8uBy+uim+oR0
yKM+eNz4C5eQNa2R/1+uGvb+6ghFcWN3l+C/EvcbWBY5OhctJHFoE/MVlLqNHa61
vkuh/tRvwMN6w1DmAxAHl2cFvjmW/Ta0IL8sFYR8qhkqxP/P30MXA334GCmyZ4Dc
gTOaluouTBWnZFhovHaXFNlvfKMZWO5hBkvLBHPNHd5w854arkgB4RBoYW/aC5Mn
P6c3ogp3DoRTPQzYD5C556CJyxNB/z2S1+G664RfvpcitXoJaLaU47cgnt/J5frs
TsinE47dVhwP95Pko8FK2E26KarWSxaybJQNe+0ReOWfIVHLEP0d/okMCfnQmr4k
sEn2MlY3ZIC0RmQ1Uhfs/6JFOr8rLsNeWIz5U478Tm4+lvhSLIPl/RDbe1FGEF0b
jqUzYRN6zKT1l2gFBNuYpnma/bme5JQSJMXHsE2oKdm8b077UfE4zjzvH12Cn5F0
+r42iPNdWfOUKRArgOZ0EFFBpUnIiS4pHsMoxWudPcLmL9E/fM2G7Ccgrg/MMfVF
+8AiTZTsKq3z6ds0KL542KO/RCQ7I4GTQPOyUEnILTJ4lVmIXKc24NRQ/MS5UPRN
sUGpZ5e41XKMrTfGh/b/JxewBt3/ogIIOwQPRXbKMv6xHk1Q+9lZreUsCodqwAZ5
1YMts3h5m3coyZLxxSBbzEGuPdBIrWrPFsDa6PZB1SP3jeRJpsI08eQZms6QIElu
t0ZsbywN0wtQZ94od4rwyGixNsyRJOhM8ONhdQSeiA50ex4OcCcnheg2PDogN5Y4
lv2uBr15M/DR03sDWI95icqv1lY+d7O07WJlssDnbkO2pQC0LZp2koQv3GGecZWY
bmK7+SIP0pHthKEyTm9CGDgY91lt1kdV+QJ4PWJUyWAUj4n6jS0RjEqR0nBwpHDR
nnfPc/soh2m54tYPrMM8Qu8tLKs613vm0S8e0L7sylerO71C5w71A8ogBgqMTA/q
npT0eSUJidhXhc4Wf26hSIXbR9X7XCxrN/I5c9dqxhE3VUnZPWN1N8fueXnbXyKJ
rNd9muHkY1aGEyWdXxlpPtZU5aMFiSY1GFtursVdMcIXAgxgXuZTVnK7kUdM3zru
pRd5U2QHlhLBdsH2/majxluJjwx3T6MRAP5vJKeeb0vA06gnjdp6rLMfrazH1mgx
3+YvS5Vg120UQ7XIkiW1TzTvBej+3ZNg0BuLM6IU/Y7q1CNXVrnw65/crViVqcfh
EcSmp79LGyGt/vGLn6T7tkkw3gSa0ZX+LMDJ7RedB9+kp8zR+xEYcuREtMBArWJF
ETi1BGIgTZB2iClupocTn+UiR4eR71rBOz6CTBZkM0CXGX72zgBRCqa+hZe4NqCC
Zs2TxzrbDhQch9Gf0L/lub30Obh8L2jj4NFEH6MJ/IyzUxi6G0v1N7ozvQp8Tss2
gdcROWPUA13/5AYoUQ6MBTOjnW0FsFMqbxx5T9mmuQ/84fpkt4ttjzLY5vHHaZmd
kUyA53WCLshFIqLt1VFFCulLYqXPJVvnG0o2VyYY92cQJddEYMj+AbjRQku0o4w/
L4eovYXdKd++5bhs6UfVRlLP59pE6ctsECJO0OyFyP3MipZUJAO2SHk7nSXzCWqO
/IM3ANe/WEZysEdhgN56aGvtGsCZtJhRRFDcVlD16liABoBTSvo+3/9BTSR79qKK
v6IDrTgp6Di6QcJsD8ZUb49imF/GxoCBJyMv5Z/8ouOnZZi6GaXVtjSvzufxSXJO
l7YMQ6AJjqgpgZxNRtgOK11RgSzQiQRJe70MZPqiq1oyEhVHzqZxhs84IxlhDYN6
V0FREYWwFiS+Hf6uv6hlqJFVQmLpYpfN66ptQxVArBoHGp+tcMjI73aa7sVETEgh
vYIUhYmoQoyxE6PupHlmw8WsDN/N0BWG/aPpcfGlZLMYNrYy08FY8nHGImU4vc1f
iTLsdzDvbCV3rB3iSTVtFB7xSeDuigIeKoREUHcWdmlOUn4x6uukw5SdsgUbeIVq
yqOnACb9iEnAdz65ly6FFUguMHo2G0/SECMAwhG50fAWBBKmzJJvuzuu0FsNlLjV
eApyvJoYvVS3Qk0upwKfG7otNr4r37ZcYcPghxcouFejgMJA3gyd9QQi3EFFSn48
+mGa4VPf3whRRqKPR1VRxabXcF5Y4AgLDuE5PAoddZYYW/r4Jyc18IpypmCQYEyv
tADkGm2+e7qvhjrPgnBZA7XpxCOE+UM+TOVb24mBFMLozC4EpIo1sbw+o8esN7Ll
rTKc5KKg22ffvdC1xT6qzygISJkPFepGVUEZsp94eSOcAu/4wT6TE/3Su7glIjYI
KwB3ERxJzjF5QwY/Uff470EKyFKTdKsqtg6aOIAY7qM5B4Q0jtC/uPH187jmq/F1
he+a7mrY8S6V8QlL1wsZy0wQTF5qk8lgmW2EE9LVDwMIZfc9SHaox/Z0w5HSj6zE
2O/sULfWqxmpE0ePE5e2V1jDG7dRb9H+z70cF7+k1LiCWd0JVZTfNzfyWFSSi48V
hrsTIubKIHOwmuL0ycEH/VxaVaK5muGxbAYr8h8iKOByGG+FSqh3As5bx4SHlCaS
ZIYx/WFkoCR5Klrr3anCy1qg7gwmVkKraLFzPezOX57IX80HJTwElDVm0HyNT7LS
UxlWOTvA0F/Kkkq1iOYFwwrj4SKL9RXL3dWX0whamwZZMYUv9q/DuQ2TpAbqxGz7
NoaY1DWfirVoXWRX9LkM2Ax75o3rgcKYY65tMTv5pddgkRf/pGudUgSpCIY+jtoS
CsQHo9umYFP+10EzNHVikY2Py5J+JgFlxU7Y0iNHg3r1xJlC6VyVoE/GKZfOcImJ
apgTqL48L3BMOQ6CdJWw++lVufNjpiQz+bRW8xgY0kXkpVgrD4NNkcyAlUecn/E6
JMO64BnZmFvIRVqFSDjhRvBM9wMVkU3PrGpgTr86lglMd3Li6W0LeETJ8vUZ97FA
vy7u5mqrXe83Udy5KRpc20TkKGsH+XgvUmpppfq7H0thrTyQCXfx4ZAKLcl8y/th
cx0jhobsvIOT/pNH5e5Xffcf0Kp+SPHyDhKnizF7Hn7RxLmR96hHUqDZNxdjIizW
fv2+g8Cr/jNvJcsjBaFH3435cQcraTwA67wIwYryTYJ33oDifpeWO5lTzontNjLN
65+7+fNiMN1mkT0sxJmzhPOVmCwadh8lhG6tJ2KvEauOFC4yIFwH1M9jWJVLATpx
JlBZQorRrn4r2e0ZMN/2iDX2TuE3ldo9rQXbHLEud4u0wtzWG4qm0bIAn9xOB4+8
3x8EPrkuzoCCIJoayyAPpIeIH55w1uiJ+uKRoiBgsOBrM/gbjudcNCFm7xWx1XZd
eqegx90J/vEX6am+iqfkPGV4oCEFdb2Gc8Ltke42t3ZuL4OORbmZUfFNeo8XKeoJ
GImntRfVJwRp22r6JQ1wmSGrMF4vhbaY2qe2ERIpwwdEJAjcYVVnlntV0W7a6u68
9p5jn+/F7txp8erNi9rz6XSJ5XuJhn0C+xDG/ZFqScfbzohsv09lpPGL0eQQ/4y9
pSWVqQeEFKIAbr+9PErwRjnkPz1Vt5GikNb4/h1V8aIU7FqBPUuoWNKdX+GNR/5R
7R2CfrBNYB+C25M0mjzTkeELnAA6Jhqt3fdA/zonoSkTIBH6O6abU/KUZz1k2EC4
PJKyc9dlO9C/xyDHB9ylpOtva7io95OAlMMVIk1w7vxldl+FJbob7Kfs1/S0ILLP
ZtEGR4vd35NUsMQcocfdF5yN4yKwdKLCgreGt5uP0dfOopeVOCoUtNYOvJY1NBcS
ZZY/Vh8KZJo1Rfu46GAjb8UxSTVJwU5CdVkyB9S9diZI3/FNG54i83hb3BLIqeuf
+7qRyBepG1VzFhKqziVfxfA1VzxntK5d45Zh829fPtgKc9/or6ipTYFQaXi0Y35q
0yiSUgllt9KoBCKrcd0/MfbWulDBHLSwHhsN10qDx/TGKDhrD+w0L3mqLBsOeYoX
rEAeztRwhf/W/RUKsPfP6JitbSP8IszrVSA6OYx18lkJ9Y8/6TUUCAa9xxB10+aQ
A71Vh60KUHTRv/m3PMF1xNIfFF7k3glE+LSWbn5MH0zEorTt6svmvvP3corhMA1r
2MuZ00b9lmHqhX4+bBDJK99rdOQuoTObnpnkjKOjEKMs8MpHQeWY1mZ5i2P9peZA
sjIe9EmGmQg0DVrJZrIKAn9rAr8jPZ80YPcLBQSyaAVR9oYzwrnZb1L65r80L2Bj
WG74i0jQh5CblM3LG8SODf5gZuCumYWRa1mpyh7Mv3mlzrGDu6HfEV2w4x4uKfOZ
5PmnSyl15KISeECZeCT4qY6/Uu/WdhtY0gi7jtY/g6TuABfE9GLC8guH7s/oK6Ow
FXXYGU/K264fSJig546f6U9skYA5/SstdY9oUJtN16MFfMHi6qn+kmINwxrQ7V7x
YA7Zrrd/hD0vMyBs62fLpl8mjElfp7qyKaREZ3WAnn4oW92RnMmGCLFfiLysyFmt
X7pavt01rwwL8H7B6rhl7t2SkZ/krX+wIibNBCpY+Wutwp/PRFXfUaf9dyGIy+c5
6rIPoO4aHdP0OvIfpMy6hCN3jSS2Ee4FAYnPyPvE+ctWTb2UPWPr6CK9uGtmejNH
FRHC2O+5rkvIJaLA8bJb1F1df7lfy7SFCc1Z7YK1lVqBPBzgBRjeoJ9GniLvI28U
U+/agfOPSN6kQxvMKaFVO+8avc9NIJ9ZaWMOO6+eSHnZj+lIRxOkukKjZJdeTYMU
M21iBLw6g7FVAhp80k1/Ca15aTa5v3AKPM9jFIQGM/ESd/JVpmy7yjHV0E+JmXt5
O6njOIPnZ7ftBQv2Fs3SvErg7rwBtkH+zpRLOZsni3oBaEqrj0Maqie4+89p/bGg
5xJeT4taz7rHZKGinhCcwIR+HRWFTx5S6E3QuGZsUatl86qrdaqzdgV9zHTOGZpM
hIiqUsE84wP0HC8PfYG4O8cBUEifkqTEyGYFABsSi0SMCGqCivqlrK11MWvh6pa0
grvBUZ7nhsWaHzLxVECk8vQPJyYASQixacF+FlGyAeRwIE0MAJDB55ndRRFbgigP
2ZWcSdLoMOHNFN1It2EBLkeExUjff/Z/2k2KHy71lDBshwXCEmJk80lSrLGHOMMT
1YnQ+U4YU6q6Aidhp2ZiuQNYfx4VfVR4W1t2gGXJjYI6Ekgy8QKpkh1IqF8Cw0ax
HmQsdsZYCnpu89LoTgUwBdQCiT/UfxbPMtbWYkkmRRFWds1Un+WJSnNSCaG8dqoq
V4G1lyLPes0uIdmfJ2cLdi9Q8+baYdN9XsEWGdaWcPbOlBdDtLq3rjojRUq/MnvF
h+ueRAWgrjJCvWA1XUKnN9rWTWvrAIpXpDamttLJhrTvKHvYUIZ/qRjSpiMTtGXl
qN6U6IJmd3jqLc3MPqFA5QZiGNNsWs62EphwHAUVSoIRh3SSCK1iWqcgZaiNDMuR
SKTNFJr6BEg7Q9Nw9DHhGyq15KxtXACyOvc9Y8R0qUsdwP4KLAt9DYz22y5mdYYV
2sGQs+Idgj7k7jb85sDwNgB6JgA2kaIiJJadBfG5XUvxCBn5+0GZ72IVW2wOjlNg
lE2b5v0rWosYGY2Fyg6LQWXvZ2XPBImV82R/jFAcFTlgdXFlmZn8SvrVoQKXJNZ5
563UWTLvK7MK2GfrVFZLSffE78P9a5waNVEE5UyRfjZFVcvtk8ewgNLUsCueaFPm
bRne0ZkktxGCYf19BemMTUEbm0O4RgoIQJ3nlQUf8qEuSqW5gNuyGKNBTFNU+5Y1
xdBFF4LREbJzak9WBrrKlezjz5U9i59FvRRAqRrQG7oVygjdLlvs5XYafwFbnb7W
VYWc+YrSF1sOf/KMvd8ZS8Rgy45Cgg6bUzpuotodkQaNKVa+GXHMA35tNvSrYevb
q8thnzg7NQmf2AB6yaSYcTcaohOIOSZg/65oIoM6nFpQUa2ETYhPjh+EPhnBKJNJ
A81o6sE7BAV9Ji+cLgVOg0q9p9eXvoi3vLl+r9DBPYqX5btSmkLi0gi1oZopTjBn
EE7sUGaEDIgI6fEU/lTFnDPhBgMWNxMKYBAZfIfYaI0DqQ0LUKxqRwHGQYYSA+HR
/V2PUhbllbHki+ckzzZERwO09B1FoBv/Fkta8x82fhusVI0Ne+t9zsQ7qWm3frNH
wW3+RPpkrzvN0NOcsCURpMzyMqPcUXQG9bjZwwRIENOwGr42joZP4ekgOEj0X81x
WPxD2rfhGCIlRN/zG1NjoPgMlw5LWygtLFkZiBG3uFrn9a0BDcVlVGzfplMgrGzY
L0CUC/O65+jpgwkcSniTzH5qSxBq2+NULj8VVTSwg7C/f8qp5m08crCWgd/HEEdb
orVSqUp7Cz81diD0MxUcL+kzZzSB7dw21TTYq+t6GUPtAVs9Z9OzPvJSg6fYIkMa
xOZwz4t9wjLls/hsxCOqICTvUqv/pBYLlU65a6Fc4IfKGN4uR13Cfs3vdxKAISmc
TqCHYQ7PqHuVlH+TQZTjskddiYelAx1n+LH4T8i5sxUZc7ku58WLQycKmkhv+fj9
slLkQIBVeb3TTN5S7ukoV7O6UU82Yrt6DWEri6HYbf+rKNcluMNDJZlVjXk4cPUX
depEYhUBnly6DxMtcrkMl+dVJicEcBjRrXk81Is3y69toFgLxqf89seikkugaVoA
sC0I6/OjWNJIoepIOCcSmtYYe9+fR+dIWxMuwcUAJT8Q1f/P5ifw0vVufZqIleEA
R/Tf7h/GnQB0Bu2p9L5ERPTj2GVVvGNBuHBd8GVwGz3VzhZjQCdbpasMwIA4W619
cy438Kud7VX2KTKXlHmjY4CY0qv3fsLsGzhZ4JtfHNj4nE+oo2ORGUStwW/kTA4J
bVLHSlNHKAALnkmqtKMuBOVjkHvDuq1spl4dVpNa548G98TCl0zN3u7/YwvA7SkJ
HxpR/zJ/h/VdTorBhmkYd/4Tl44kHTemYpg7DOm1uUUohzODaSA5dnzZDF4CyuO4
rHektzXbdwq9L+RFGI6Z76yeRBi79I/JnWP+HOpDOtJRjFeS9p2AMEPR1Vp/ZAGi
k9LQe4aulNW4fs4SDcERXAL6iTiEvNt/4NqP0x1fcg1QjLDJoUlTWZHWvb13HEwi
xDBImYosgMkX8aXwmYolgOgmXhWYVAp0j5m3H2Z1qeE7QlE3R7hIRPsTtA/l5wFC
B/2Ii7K0/Qmc57yEqhm0MpnPWATHrdYWgg+TYZZdGDE+S228BzHGnoe1is+Fc8ol
iAaMfyDJlSiWrMOcIqRop3aGnIvI4w0xu4ro9u/lXSrw0nk69gGAQFjt27sXpxc0
smOW5UmPCbArqGFeiZHreiXLzrNlHRoMXzz/Jognp632/DOclI0pV5ZWthhhn439
DmMwyHVnwLN+TmNlDm3YAdeZ5JRkR0oicFUkuFlQq2rE7JPUD56OuP6PSZcsY0dZ
S0i3qyOVrMU96l9U8RRIDoaqDjslwAPyLVOSZp74Wcd7VyobyYEqvOqMr/xM8XiJ
G0sH04JMawxgxU5a/7N5pIJ8lTFoz0yZ+oDBDKKmHDCDI4EER+1SAHVbT2ex/8u4
HVXfDUPvn36l+l66Jl8cgZQgrjm35/J7ROCrUbzcB1civ+fdxNUPZeingTDKDSaE
RS41RQzsXxF5uT3DabevuW7nCWsZP7wRpJUWc2242Wpb7A3QVmjVT5RyPYhHCAOn
Ci2qOXB50Jw8K3LVjQhKf3jA9nw4BL4HPAF5OShATYxPUdKsZcMujSFuQmsKSliE
A74R8DJzuvthzZULzA58vYwUYTyU0YXnBHItaQ8MvUz3l4TK1b7InxTtRq7XZCii
kxUbP7MC+XhhI46CG2kRgjGDwUj1KS7P4bNX0hTeqa57Wgkhb2CAvIRo0K2JjlDq
KIy49x1DMfskDEEi7htSJJpqIPe4EgA4gDO6SctnHIm2+plVkSLHqoItxFCNz8yz
IuipW0YuHKVdCw8EibmrpQ+3RwC/D2JnIKMsR5PbDNcY5tzEj5o2WV7mC6Sqptza
aH8XHXhiDinZBJejONgjqI14DqkHQQB1Nwi+Pf+MNd9PRP4ohXSs0YuPuNewt5Ty
2WHczcSy8dKhvXx/tKh4GsGRwPWYRaa/nh4f+5u/Pl1/w/7OUzWw3TEx63IKTfQ2
oFI1oNVkjV6vKXICKKAt4Y6pXMQJwSds7oPkqi9Ap+MzUeBvZ+B7vfB2YG8ZWE2D
f9fjaP/0jqIp9LRT8kVSrSkB05bVN7xU9yBZKUf77sWXfBI7O5L2Qj4rU/lE+nW9
A3SwNOeDqndYZx/aKAFyYrzXpXFFsrMEUR2Wp6uFUNNuzJzkCswMzAKN1Aajwd9v
1wQPy/kNnpmVk3KElu3yWsrRyl1VKZoJlunGtxTpYwRkgl5eSfjp2yDqRcsvjxfj
9IKzDNvHwG+yzWUbr6/LYAdtUC7OcMvEgK2+mW10WfbuMcIhaVzEXvT9c5Uagopw
6WYW/nD8YHjZ48KMdtnEpoSCVWGI7tpgz3PuThfKP0D8I6/PdTMxyshOacqH03Es
haHv46OsD1M9YdN5Nw1j8CokYL5uoEc3h/Da7J6xYs1s+OV5CHQDxcBxCfge0EVk
QjwrN2YQCISMaYh1VclFWDTH/fqFwMHK2wS7hqnwAjBnyS7yTb/xteyvw2D1tLQw
tr+wWyRDRLPdjRCAiRZ/kzL42nIXYHubAca9rKhtYCQKvajQ1c2vYf27sAcjCWRW
x+hXnQNqY8PmTurhcnoziGkHP1GirXozbTnbUcnqqmlbeTXWESOQtTGfRnu46IBC
ExYna+H0pKawif4DFx7gnxQ2buan9C/c6h1+08dlqNtRF4c43WwhB/qShii+vOU2
m1TIOGeltc4kl99jskQOAAFSiesT8PeqexRFW56HJfVOWhT6ewP/Jr8fEB9AuOH3
Xm/lif9E7nOQZXGjF6JFqwNCY7199rNEBLOaiuGY9pUcW5+cmJt9Jz+P55da4UP9
zgtTRd0wUFXfiyWW42sYzfxpgBUeovleKnQgxcHMmwp6f02tBEQLWbmjF0Fg/XkR
dlakUL28WmL+Dd1ssJFUoFJH6LUsOoRVTZapjvigswWIvwM+tovooetOEZKN8LQ1
d0Syb/iRps7tuTys+j6o+hUp/wnwxfQ0ONefcAcufejOJgyrb88FDdL5PMs9xYcQ
YARdP6Bx7k8ncRHCRzGgmvUnfJHC6LGw6FUFqEOpjIWgIITMqfY+jA+shcgIEpGL
AaFfLpfutLKqmqbSIM396ezk2UnmYhOuPOHOFEmjQIFUFLkE9OfWMqkJVs9Bud71
ghuKxkP3Bm7sVVFrW5laHS8iHy8S6kdrUuAElwPd4R1lnlw+kUEvutq7VPSteO5D
6XL8TG2EqtvQCSTUX9Xy1rqw9iPfOHTdPETrJwRxcvzHabVn0Cud9nnuLLJhjEhy
brTQxz3xdNnC4J5Yk5RaDxDIJfIkPCL7/xAZkch/vytFRVWZry382gGYKnLieDLo
QrEN3jPuJPwh9QtDQvLASDfJ95Km71ZFN1zrgz1Q8DcJ1SXtLJ1pmwoTBSJX4++7
E+ivwbOxVtjdiLRwi1vOiLmak08xgALt+L9+Dq+RqjiDjuSgF2xUZQmTEnwrfXmH
XGVQv68sCI6YT3X9FA1agp21T+x7Fp10aNz6EKTeDGWCxJfhJ4nTXLqfAYqWCNdp
r03XKCWAvl6kUgNx3vsYrhxTBBUNYU11bx3CSwtcVf/lIm7yTl10K7zhm5dSbfdn
OPNoERWAxGRjeL/LMW6S8TGh6ORpxGnK/ca2O8+nQCgZJ448D1ul979psjBNcJC8
7CBjCOgwueMOXPUNWy4MGR9uzXAekedQ6dSsHw8Nod1AQmjLRNM+QB9/qG0g0xqX
rgTAynE6zfgm3xjLqOR/HlfqwB6UkwziNzIplstg2lnjp12Jt0tPQk405utbXCbz
JDN/q92BAquSZHssmvlNvYKn2WnlRrR52nccJCql0UW7URQ30zXBSoZCGcrWHNgh
+1RlvffObXMHcJmHS8sekQvDg35EEiVTNmwffgC8I4bSkFXMOIF1R2UT/9GZ5Tat
Cr4JaRylZo5j7DfaQxDOzLRndExaUBRBOxq/MSz0FIrRgZIKd/EfkBX2QIu75bzZ
WKIJn4qTJwMdm+3P6j8iE4W83DfEF6ItwmEyzgBfzHN54wWooLjxZgERv5DSNWRy
ofXgg6Poc8WsdziCtNnWhwKdtQk0pk7UAVlbMNsJg7rOIpNT0324zB8nLf6nhSkJ
rMCmWUXAemeyRjc5o21RnjzFayHIn6o1Vout4F8xKzMr76saM+77aYWOGbodtyuc
b5ODhuKWFADXKzOe8sx2KdWHe/ugBjT6slNcnaF0e1TyTIAynH9T3/Ed12kNmW64
2xjePGxjbygsqwqtV0hRpdVAZCmKWtuighs4YZK+3dWRucSmPO1kw8WI31o/lD3P
61dzhztXw7oNNrCWLCN07fs6II7i+BE3ihfSSxu2As1n7jrOTpLtMC5S+1OeiyoT
5H3BBmy5lOESitbHcXLWRXyArRE9Ryuz5WWIF6TXLl6rHFlZ3Q8ltu3/Wlei+97k
6Pifu5oHbPYmWbn3w3Vu6VoRWd9kla8hhc74dhEkI3brnk8dOhbSDJ0zr8fELCqJ
F/dAwPq627HNKqJrSxnvPBNzVCZKyOdm6KKTF1zAW3WhR9XLLMKq8O19ccN2D2e9
xYd2juoZ7XUdvxBrSc6cOk3oSFdFuP+o3xR5kiQ4aqmLrbbBRnMik8oNuvqmUHzS
CyEBW0huXW31u4IsWTQYir8S4a0cSIPvqkXSRxtl7fHasWBzDt4M2by1C+LAYez9
WcMqcXBIN0slp3KohywBA5ZpXuWMaWfm+YuZj3MS4yhC9ZgBh4Nq0yqVkRftLOxd
bEn6eeRTxT/FhIQy0lFuVS3iud9IRT6bxTylkksZhlNS24hPgYmQRfWxBQ4K/TWV
nf0AwCz6VHxUAyi8Yh0KjceaR0lTWImq/IMaPriz74d/AffdSWtzXFtD7FcfNQFS
hpvyUde1StvwYpxXcBfTlLSbAD+rKoA6gZTQFfLdP5RHpurhq3IFcIufgKhSTESW
C/K6FzESfGwRwxgvZMzNSO4pTuliPwt9rbXbC3onivylQgJACgsxbKhnyZ4A/zE0
2y1g69jd2GcJcRdTZ5N/+jMZjih3kZtGsC04yIgpj6blpWDwD2pQikaaOwIIiPKd
mFHYqrEyqM637Eidb+97R2oVhejlEZB+OeI8FFLwBmMVoPnxqxod+Itsz/KhnzJw
HJS4KDD02fzysvIOlzRrIbyl7Pof3vrxauL6A2rUPXJ27METWFZzIzAzkr1Vp6Ti
+sBYuU+vCIUwr3HMEyrQr4ncsaOWIjEltvyEfy0Sy79aUtNMt60OonZOdPmSf51C
NTzOfH5yvTZBuLCoakkx6B6oeuPdYRV98aRkxc4fFgdcPXNdu6GSKe9kh3iOaL2E
6NW9Vjdazp2clP1ujna/JGQolc50CmnxgMLfSPB1t7FeoW/iFxOpjKPFzizl581N
ueSA2A9GMm05OYDht/0MWvh4sV5T79JwMPyltkH9fwSb/PpClXp7Jx77lkStgCVq
j/BzcCm3ulzzZEYucnio8oz8y3VIB5uXWo2rbPPxQKhT4eKPVckVKItS3kPUVRsh
vaH0K7B41pXNJJyb9sLZ0wsOQUnB8IlmLWgWdvQG9n9BuDB3UsglTgdnT7eSfL4v
U3QO6k2tf5mo+90D93UE1rclQbYtI7sHDO3qtDhlfMcjxpFU8fFH82CHlHOoD6ND
Ty1HOFw1WE79uq73wyY2kdAPw4A7u00J1S1xMXG2GV9ToFXyouSs0+ANAdqFywv0
Np4pqtXbgy1nWrh3aDPliqXSVyJKWT5qOJVkMPYKqT2RHxHNsVG3xgyQjZWPJYrW
kPoqyLEoXSWcTKwtD6JhMVjVoRsjK7aQ3sRCO19jZjQeXe3KY2l5hCklNNF0o/eE
81FvMhCmbHwc9m5lu7PAjd7bhL9yOSl5YRiq9/gT1IHIN6sgByuRqX0l6Y/NHWcv
c11jHPtUQ0y4L7AiS6K0DmD+8M1G2yogxyASS2CsIq5L/ixBt2bfZDGfyHa0c36r
PFI0DRgiHYHlptENGcUYg8LANCXsqR+cOM1hH10syye1HcUjSzuQLzQT8mEpuLET
mMcYkkKrDfps+UapUzfjTO13ZutmvKBa0TktmTiytuOvxZzMQp9YQvogmg29z8SO
vvgBSU/Tof8jVin3ovEFGxO2e94I+vonNzF4VsUgqdnEbPLNkuyPc0GyaCHpKyPv
pxwpPXL3mW78lXorSz/CcFqp1ZOmHExIJXlkKEPV6CyqVr/7Wb0QmHvdBa/TV/Pg
5tdrVT6+1YGlQvldCBw8zdfzExKMX/a02B8FOSS7CsXjTHP8ERd4NBxNMDJncSmS
jx8lMnfxIoc4d798fO05Uk8Q+Wu/zh+xS3pVOA7UNuLMjpJB5ecui3wUDeyiAyYY
nf/ctBpaLbjkEp7rVLdkbB/f6H6E3hkpcEEyLzUTfGxbLM7cYKRViFbK9Vi/Fxhr
qRzfjEsI0YivbA96PluejdSOAf8058gTcomYfxlQHkVHf6ta7x++xwfK+5cmkAOA
WPg5tfnCNtetN4vO1UQnwQWuV8uAY9/l7svoGo3wInQL27OUPZ1C71Dxbd6QUu1j
COTLoksnbKq9FT7+LzbPlZSQj+K0kl237XZmesIPv1Sd/wgOrSt/Ub+DXEogX5rt
NOlIrFCLWPzk/Kk1XXIBKtA60+JGKoComgbOBr/7TAD6WUs7uTx0pu0NpsI3pN+G
cpifMrlBB5pc4oxZUDPeGJFoEoRu4Z2pxHGhy1KzEjmiew/jPbOkT3OPzxItcw2B
WdQMHQQJwm/yFSwSStMFqcVGk5huzjJN7ZoXLa9J2QUdLjdp+Uli7VsdeN3g7T6m
5qN2yEOb+CDvQmJU+PjjcPkt4MWl0Pw3P75RcglbOdZ5B48CLaHRREl7zukzwNP1
LwK4Gv60gIM9xPMG7d+ENEkP1CAOae/w9jMpwUzB0jzzyM7CE2isgUPBGIpSHjaU
awep7VfZ/Fo06Juu1WY5NQvJ0ateogHAEMLe4NHW7Z4FyP6T5YBmLmbD6sFS8YIU
VL/e4fVGut8UNotzxsoTzMFFuYKvp0cMi3W82h0g6OHXcpem2sXx/fCyuF9nHUJJ
cSjKTzFenV6arS/QbQuy9OfCjQ1DYOgEgQzJdzxyNP8Wb8yihztShlIHGadwicFR
zqTYkPUEGi9Kaa3ivDlCgDE0vZ7zhXI4D8or8VQAMxIyx3Z3si0AjeDuh7B7Er1F
RfbglTKGMyDXbyLKulEG4pGhsx9Z1zHM5se3QrYyegp4R69UOT/AoFWMKuWZt0Pz
dwHUu9XoT+FfVLZQeMzBs5BK5fLqeLVyS01e7OCbVP4GfBNmRx9aczTx7TCfBbvT
fPKFIV8m2LFkDH97Kxe2UTauqv/BIaxoU9Afcj0FJiw6qzJiMMN8tIcBVoYD3dD/
We8QiVmKgvEkBwXZbFzcZzX9Ojhs0Tu4obxSmItkvDYhONTHcNxOYbM4y9OLb5XV
78C/6m2nVshrFIRK6k3EG/g7sz/flWPSFJnUNlPwsZXzkGSptWXRN6MMdlhheQCK
QD6JsjsmEKXXWM5xCrq48OwOcH+hlJxcFD0rvYV/jrTmeaxjYgXK+IPY8+7qpKyd
2DQOPVIQIs9r1typ6tFOoCmnL1aFk0Vo1cGfbuyZr5hH0pKvfgqG7A6DtCbQyLSO
kjJpc9zB/7/r5DqDPg+96E5MoocG2beMXC7hHsaN5QoXEWIIoC2BW4Bec+54A1BC
7D2rQJjwDV+T7M0jPZIZsm4ChI3gYt1Kj5prl9fFk6ezhWMDXMxSsKp3Q8iqoGFi
QNHIw5Yv1l2xWli9oj7aYWkvf+2ntEFp0RHvvyTfMAKos9fCGY4JN0yAgBYfCVO/
x13BuDhfSjdvkGPUROtP2mlX5PrzK5v6hk1oyaVswPCeXLHMVBz6QQcvJqRllMlN
pl4SxbPWINLmEYtaWu/PhNCA+Z5OCfIhnH7SXsOB80rS1bAh4Bhr1+P3EkBJleTy
rnqPFb8kcmIuW9I6bLjxkFT3mDo2WW9pB3/krDIU1Rzh48YV0q66CIA0G/j//KMB
LsMOYay3idDez14weJGcQH/Wevv74EproVLmbvMYWc5gwo45GNlmMQFUPWvRNCod
Z6qrIkSzZ3n3qR6Qi/8bSz7cJX1Sj8jjmKVeCq80NNL22dLpj34TRfxggwrQWGmC
o1xDN+ya48SKuCMA6dgoxzd1BnfZtsxICotyMnmj/XO6K3Mqum9EkiYbfa7Zcv/c
mwb5OUMNJMUO2ZCr1XNJ0w+c0pd0/QNWJC+OFhp319qVMxqL+cBh2+Irzehb3MLa
ziz1eF6jvR91SLH4DYnQGEmxXm8a3lAbQQHZpR7jo1g1bCYkSRDAwIORPEKsR8+p
pVd9dvBHdeGvaS/I3/Vl5RvjPlj6il8Dne1brXBHdvZLU7l/OsrI43IlRDgPUR3I
V4PyuS4W9s0mfal0EKezgUqwQ6E9egT1yKMsK4tr8HPuA0DMy9oWUh3itVz1YV+t
Azc5rxZ/rEu67L2qwnQ8mJ3BgoqugqDOfbPFP+Sb6fJvYIoVzY1uv0kzPUbfeLsI
H7DjD8icYcBAh8HgBz25EoMQluEgvi/MWtdJsOyaqcwgydYXukDv/RRwdwAfoCHz
RXQqfiubY3oqh5ZCxN6NN4Y8S73qMd8AuC7X2Xdnrzof+3v8ABw23KMWLjz4Sr1B
F8evqqw3uOLQ6asYrK7SvqyVMV/8eQiQzCpeq1Rxd0lF5MUdC9BqfrYTTBeIbr+3
mE06tEWS4Pi62FytbaWHNbu6FBH9gUjjbGpjmRpB+LMi+UciO5AlJhyuRpadffZC
Gv7c6ZcTv5AKv4TP8aK3az9/ZgcvtcXBkew0cD+q9AZMDH9WTTbFMy/2ldz50KSn
87KAR71AfPGmima2Cg8Hj2aspA3lpx4D7zO/r2AbnFEBNlJgSMy4fPh79E43RDMC
FHPSdTICY7kZVn3nTOmJh+PJCSK5pQB5rM5QizNnRr4kEvBevaG5jch5HjJZOF3/
s6j3NdQpDsQb4V45FnxN9A+vBMSGIHhukIz1Po+FhcfSh1gZZ4m9t58aIL60nBe6
RMYYpNhL8ljrgArBmOT5dGRg3YAlV03sBHlOl05iT1R4Qf7kriLtXZqoxUsnqwFo
Pl1mDcmXSxh9uyS2+ac37Y3iL6t7KRgSZ3BpnIWxxkioJleyBDxY5uzn5+X4fU2L
gQ2bxqYRklxmMjfn4gLK3CBWhzTQGUytNDZzUEZ/JZEZjyQ7+Bcnpon3YSzN36Qd
CqQm2DwGf4nDtouxw7eydMGsYiGuqz0n4CY2n2mMKuKAhYdmz99JgRweRhZQNoX7
IjMcdAIGFpxHyEqmfjOvmH+cc155qxSZjcJDK9vC8gSsp+RFF/S2PgTjDFGCvyfm
1RtKSYW2gb06oGU0BtM1/LzYAJiU7gu/avLAGBd8Ogg7CXDKAvJFzqBReuwSxyi+
T4QJYPX+KG4khayplbrH3CTNHK7YFwVCPQ746nyYFZ9QNYcwOhCc6Ig7PfU7PU8W
gyFfd5bYvgJsoQZDGqT4yU+CIk66QmWvr/FuMP6enygkefDb9+RpPoDchuXmnpxS
py9JTyBYYKdPKgA1Iu1UZVZrbl4XgGvckU+umCzfeVsbIcVl+ucbwva4OphOs+mQ
RupXJz2TeWSvQQeLAnztv0AAknN+Vl9hMqSI9f8BqpXka5zb5VaJMggRF3pF+m5M
uZTDbENmsR8PImenIRdxkMX62Skhh7h0RJTmr1hhU3fw0lBuY/mk9CyirzF/SNg5
ZIj8QX8noT9fKG7ssy2pSRCx38NPHw6fcNDXVc1nZJHueWs3zJ7dnwJJvoLf2uKB
/RklzGDgrSUmKGdfIfco7Be25QtQRmmX9CjKVmR1ksr2ErgXmmG7e7YuJSgea1N7
P7GUEJyaQO7tUVLQa3aD6XIKAri81tSMqKcBGsi9Mbs/v7UrZ4AQshBOuPo0QMCD
hi/VACVxKiUtX+jYC7MFu4lgCSbE3Xhmbakmu16PZKP0Dju9iDaxMOZhsVkR3SyD
7SXhK0iW88OCEQAjaJN5fDEE4XjUlyOgHRbQWp//jbR3KD6ng8G9SWezWl3SaVz9
iZe5WbyVCBVtqwJfXRuAF9pdHhyI5KvTUSycTdGH9ev3yHCpErzvuzeSvbXvHbI8
I1eEdTmXVX8WnBFcHREnv7TWumwQfQ8xG4z2pNPyGwZUoqDQGAOLU8nFYM38fYib
Aw1cjTV0U+qnrqOnnuitUTlVPYn30RhyS7D4/J0LqVcbxDHCmwzIyonI684EN5f2
d+QWq1JOAvY/kx9/N9m73ROJLN7H6GWyro61YyuEwQ0/lrJRLQJUJCwAeC6E3MQ8
I32OM5QrYGw0SMCqzE2oAXPR/JPc6HW1YNipxa+Z46rVQ80/rAzuALvRROCXFd2R
1E9rB+m04uHdBesF709Fydk1fsPGfoeKomEjZcj2523T4CxoFx/dfRUgiTf4uBWw
JkYATuShS0AoelEqxv0kp46yd52FqAbphKVwArSrDzjWA3F/LYekwUKoNw5VZS/U
VQsVg4DTdeIXip1s0Bv8dLDr3XzScaOafAJ4kLFH6PBrhIgT1bN/9iwyjC70ykAJ
Bz4+eipPHw+H5hp42ZZh9T6cdQTp97gTa18p52wilEqaNEn1mBUESKiXYnHWN6RL
+pvgNNoDL2yXN77C/6U426AC9qfB1bwY4RuxSHtMptMVuQHGtKsUTCKO/DKzts51
2qUsaJDRRAxM/rT5FoW/4Vu4jovjHl/prIddq2eBKaC/MwdpTPMnzDmuZnKSzmWk
HpQgkBy6kxfYqlnp28CqZvxBMnTotisWp0+qn+LQMmA7IHDFIE+nznaYnUuUF84v
6pBObJCau1Fu/wzM1h93TJDvC+pNqbDdLGtgAlg6fcRGarfp3rD5SITl0hHAJIP2
eTKWYEld5Q1xp2BAYststJc477Jz06bTE5K7QDLfZrz2Jswm6DCXYdVOaZF1rdxB
F2BphkVFwDoQ9uMYaP3eSKti77hJoJ79zdFSY2ffs25C+L3vF993O5nj9yK0Trqi
j93nmzTUyV0IJdQKQ5zeD3TlqXMMGyZvVwydOIEac/GlMxt9B1YOWrKAgJLhJo64
OmIoFygBIpXShHUMaPj3ehA/Zg7zujUsH64EVMDFijKyKZ9NxJgEZaaFg3jWY8wB
T5Mk9a6cK8kq9HwE9xRiQNOTlevy+OtmV4NKyT/qzu6gIgn5pbuQPYJi1VowKbKr
WfuRcmGmYOIM4FRRa/1BLhxT93DJXSbyuYnUMAEC4e1gCa14qSshND9xeZEPwphd
tYuKSpl91XfgX3Hx1OIIRcRQLGUbOGDz4BPqE7R4FvpBSBD15ueSAFzfLLQ66yYH
nhmUIjWwYbAGta9zBCHqrRXnx5I97iODKMd3Vzv5Kc8BzZW8GFPOwQ1MhtfyuSi3
zaqoUox0+znw/2Kks33ktZC36gI6tkfCCjtUr/DHW7BdfITEImSYFZDxaId9lR4w
yXUi7n3p7Ea/s6ZjxyW6/uFfVK1fD6lt8QBzZUGoUtuzO04edBEmth8W1tstc7A2
OJJQCmpzA6Ot6NAE/SkJL7QjV9s9b9iEeX0anM8SWPYdhXDkWd8G+tu7nPc1C1cM
8u/sdqGgqrAp/0U7obLIQCjIiuv9Rr+hjtHaTf8/bo4KxZwTLUem62kxC0xMiN6q
mgR/B8xDJ1tYu/WLQYPe9KeMDhoMrTQLSe1880WeGuuQjM5dkq0+piokRCLj1D2G
s4NzR8YCp3L3AAb3iJ5UYS+uslKdpLqMFhboouWN53cdkOCgpSzrV9fInjhsux58
bCWgZzW3unSyl/BFlW1DP/iQsnEuJ9j4wsfUVc+cMDkdQj9fnKu4zwc5dkQRGquq
2wXDrQCTGIACwdcdtD6bk5snBZcsOwdmzbJvpzzMJvShzOwrxqEf1itRAMZRqETT
AADGjbKVRpoJ2t0BMLe7V5XKA9DP1G1N4Upy4OCfTdadELqqE16vukx4TwNrCXF1
d91TDvpNTqxXXGiGt5mDQ79sEjwebqHoiQYoIAFRAlEvpX7JCne5lVwhgkozStNU
IrODUMwdlZHRoHK8ry3zJmyH2oCJXAYKf4NeJNHBu/Qo59Eu+e9fX4D9o7iu4A2e
pfvlDSLREaq01af5R54FsD3OS/K1H6bnhoiJioZ3wsmFuPdpWaIyefkoxx4BdQRd
TkdS/maRZtJc790PA7bxWzAY0eP0jVR7WX2xM4tbATXg/2bxns+YV2X5zG2wamwz
BrwLk9IMDkyNartUE9lY+UI9YbEKSFNOwQa87hSlyegh27yEAgN4/fmFR6/c7bk0
74B7is5oNat94E/lwBxgRdbLe5HGYKYkSq8k8ovWOjMulqS13VYk1N99FyLYJ3QN
K9SfdZMVP0xMer/0Nd5mQfxSE8k63OUv/bzavgIiDadYNjEp+bKJl/jIKbR74hFu
J73A9mGlXuioXxmZgbTHsX5tLXUCiPcWgvUV4GuQ34WR1doWi1N700JWCRkxEbtT
CwO3rCR74OdPxP+wU1JcybKdp0+7EbtLuq6mikvkAOmlrS4mJX3y1+7BLHRBJLbm
hn0RrBGnIRgNLr/7b3AJJkwGn9EEXeud3KRsheX4V0xGda6mRrM/VHkI80t1W97P
/HFMXhyfTxqI0A3bAtyjbMqeYpppOzFzTRu0s8+8y+S5N43rMS8SxwnB+5KyolbZ
MAugKhbp/7feqF7QKgQicWcxsKi8NRnavvsxU9g8oSvq04Sn2QeIv4b+N6vdbcK8
+VRY7Ards4BK3vOXcPFnxACoG8FRjfCr8UBN4Uje2xExNGKYFiJ7CthajwqFZQeq
DUkHcXsKLcno7YGyBHQKfBJGeFbP4DIps9kFJmPt3fKBSXhq8/NQXJKgMM1Aaw9W
B6URDLPnQ7BVc6Wg0kgU/OtWHI7jfBcLEu5WHx65TFDn6F3jRfUgRoS202OAczv0
pmfwz5a821NptEkSq0yb7ZF205SA+5pb2AkzQ3pQ0wetcmAtIPTACSfHW5eaXqs2
AcKg+2mnD9ka0GdnjMeMnnIgXWJunb6072Ox3m+wmaELe+aKfAs2q2yZFZFy0wUt
/+JXauuSixU8zFdUXle4YJ4VOYHax1LvR/4pIiVcZcVvOhAAs/ieybGVDutAhV+F
ZckqXoIO9roIPSlKIFm2Q69z8ZyplB6ONVw8W6jqYIk01srCABvwDLFaAONd9MtI
LX/i5tdH8TnRN1PW1q1qZ/kGbpa+8wWpLJUv3FTO1fXWwL3zQnjk1yDVaor4hT23
RE4/Y3TaoGsrLqCTJ+cl72a7aOvVK0Q/4PHUnmRmibAt3GxknsymSThkFgGW6S9O
m3igR2JWjeA9aKYJGY8ffUpai+t3DU/pYBpU6QBQxPvK/b50H/D3mJASETeVNjYZ
9mE4YqjpoJ3m/BOUXqL6VUARYOU+Up+N7itqzvgZV/3+hSYFvkYyYdOHsTuOkiE7
Leo1iuIBY+UnEK9aaH/5x1SOF80wLUAPV3XS2mWwS5SGSHv3kvXHarrnWu2ivDaY
n3WTa/X+2XpnsPP7p94NsMsa08zQ977UuWaDZ7hFFL7F+r2KqFD3ai9hKH4Z0y6S
iAxGExPQ9vbnBFOOZp9KnBy6qgu1Eo1UseqtnXJiK76y7fcjJ4+JOUEKyrsjT2Tk
x+ZUvLAhCjkHZkbD8O5Ka8zT62CpXtvFw9UzOWPS+bC9evZUKPJKnVMUYE7Ks/Qd
CyX34nVZ6PFy51eU32czVIctA5pxdi0/FOHEMVsShkGtcrDBihQzpvSyLqAJ8iY3
Jd+fmZ0mPG+k6cvQYEGEvERtnbzs81avdcU/57/Ile3iiPwwkpxOtste+qkm/2Dt
3rSm9hHi1WgHFhF6JosJjchVoaHvVMi9iJAk5hUXSRYv4R2BgK5w/cGSUGclf/Mw
B4a2nCaAL8l8KS+1JVlSkhLKusvKAie9JRVNQ88Z5NACe5utTlrlENcSTjbmXve8
y2hcOUQBuXTiE3tOvydqaH6IDJ4SjSf/w2v4TN4vKM4IpDwNqXMSAYFDZghCg4xn
YWkyPAr+3THTZW2Fli3uc6BH6P3hhyE4ywuaTANqHCgpAYc/KEuEjfU3Ia137qP9
CrqGoJAitmL0/M1SPJfeox/Bg6ZXvU0Nr/FzaeRM7TJg6LkEAkMXkX1ONGOJuRuV
h3VMZYj7tcEg/gBMTDzEVsT7pQeCB1YKHJycQ5P3cRB49vdAHLa84Yt6zU14VnCa
rMAmK6cZ7WuLohUAz1VB+IrT8jtgfseBIw1e66aZ9EONInx5Psp983n26ysGi8jg
ANnGy973SLDxtUltXceaM0CrQ8fuivddAsyQ9QqVaqH/BjqZ7SqC6zdblB+3aUcW
h0p6IborFmCJbu467pzE2ZIMZ7YTChwQvg8cVxMdI/GyCkTYuepvDCxzN1LTgK2e
p2VjyefnConBoGht9THebdIkZMChl/44bgogjUo+koq0lhN0URLW6ri4hdlP/PxE
x+tBmoc/7Uml6e4WlmenjTFAX+yc9mkkj9Z7v88/7+FsjB3fnt4Pcykhgma5QLV7
uxXIzg64nTBDjqQM7OaGY85oh01PRIGj1otodU8C+5v5Npy2DrgYUAStLZtEXK6R
BHxiuOxVfm+jw/zEXdQYqVZf4yZ71MV9vzvM29XUIs07I+L/1Cud/m/Eo+e9gqKM
SH3z7y6jwTKuxv72HrsQW0fJfaXdJx+Nqzc5HsMf4INTr9aV65kuW8LX72+RxvbP
VLg5F7nXILWoSCJwjq0C8KRVPLHk2S9QZJylzEALUHZn1JA5fcu85OR3ZP0GidPs
I5E7Ksu/HMbybqAh+mVK8maq2SKzNhVgn5pIF+ZYkFSeVet7TwYR8so5lhexLVFv
SNxUqyARHBc2MllFNTC54wIychghwVODG4be2w9MUByaykD+FiKxfOM+k4P03nHP
X7/qEGNp9e7/0Yq0qtPxYb9dTPj8YYLfdoABWzZeIUMCOWgM3WnyObLQ+a4BcKkW
t5m3bslx1zV62CePnZCSXZ78IghU1hiiPOYqqItKY2yIKIlQFyDbTnfLg6lHIxjX
bdOwJup0yT2kp0tKax/2QxQatRW5f7iWxH5vo2uFcMhAKXtuAyRBne2uq1QVDV/O
NHvNFuJI5PZkiFTs7ciKFBC1GmwKasAOBKgqinhditPRRlUVIFkyJG9tmSxdyzH6
C7AC7PFju/jpueQUw7VgAHaNot3Bb+EySoxwy7U+WCZUVd2BiFUACjQ2K1njxKr+
+dTW8XpA+MZxh0LoghIqApfQZ1PO7zIBV/XRwCKIwGfln3doANny6l9T3phvd2QD
fCNwcaLzDAuAYhA7V1jLaCJpDvYcriYtZXu+BiregGqfqEm/ScA0tputLaMkwfuc
wCw8HY9rHO/GeTpVMHsFTfl8oycP3oYWnTzSf7kbxrJpWWo5QwdzmeigbOZO5S7+
AgTAqgUIzg2uDsh6fj2/umlqlCr1RTuhN6ypvN8+fc1BGtWzpt4w15tpm0DrndUb
O6wmBI4cUXicx8Wbmso1nMnpxrPhVITVQESOcNZkIKjt6jK6Bxk0sPxlAolnZD2g
lTVPeSXXvXL18WpGvY1h/um17VIWpklFhnPez1m3QkOyaezYyj6gnyDZQKtZFm3d
A9Lo5BY5pEygsHM3h+K+yyrSCNw8tH1iVCkMNHZ0CNywXhAdzFClgdhqNTtcEyJ/
zzBNvlaGjFwdY9SBxGGh02O/T5cpnRilI8qZvZ12ltbl8xF8euKlG2oT+oUrXCte
WrIIHfUtRVu4VKp3RJ33F5/LjZCEbpxvDyG81Yy2nzSO3cd9Oxpbbd7sm2W/cz1O
o1iY8RsEvsM3CCLo982negRwvhsUUK3WZEq0BLa1w+b0iJOvK4A8HxfY4uE/np1K
lJJGJuZ1KhUEPlIWqpUZkvIRqEgvEn5gSU4E4CfB9kSIDy/+6UhZFlZHnraaxtSp
fM9DgfKXNnBPbAvjA0kWp9wu6OW0h9l/WSFZwnczmoUi2LSvxR3JOG7ABCHd+gnC
F6brIZ6OB0r5CGZ3akfqmQlFVTR0J6KtT7j2KVupHMtG2bpme7u5gpbCxZ89yrnd
pPnXd8dUPwX8xDObmuYo5d2wlk5L0jLEu3pEZA1xdGV+IR8/jD/r4kB/+YzLCLuS
gP9B/xvdnWnhtZBTRT1YEIhV+/Z4KYExTxDEApihRySJLKeQxuUVHYzTVu1fSPRk
GLIJ9m8DBjm0TOf/hQ3BGZKp+xoKRskcUPtkiGpxCJ3uMJY1C2QsYjlKmFntbdQC
WtznPSSAXL1arO18UYnqTND8MDYNW1wXgSBbnA/OeNfBXDOtY6vhzu95ULuDoK50
SLXZIyGDSNHNQFLEYaYTUD7AOxmMmerfnwIVzzsuYHbfxUNDeseIUmh49UI8ELyp
zzWftrkjdmde5xbFPYochqdf0hqaycTvUES5WI6rNuPvqlj5AxneKu3Iru9L0iit
1rOmt0poeVd+MagxbjupSUEzuFM3ZgEAGec1grJR/xeSZz/YuOLu3nl4cfqvikrk
rCRt86dDo8XRbUsYSscSUnTVQ/65qRwIPGvr6jGsCtboMI8tfN84C6HSwahCGshL
Ry2CNP9rV9VCtyN37DEtC7ssmHZf44zy7FeWhg3EOyaPbsJN5dIfLHRzHj7HBRXv
JpPb05SwG639RWjpQGyNqRuYb/e5zghDDfydzOhcJmKYwTp+NL2Pqe67UcgaWLsk
SPnNp75JpJMBS9bTww09SbVMn9OQjPXr1O4BtYXjIgokCbZ3bKo8WcJ0uGHA/MR1
J2WYouXdMiNuKOpg2CEM3TZy4sYFkcCvvyk1JI7FBHvkEBEmQJp4eFfPpAZSxFut
DW1Zv+TZRiXpxqwctDb66qY8fVvL7EvOVopmKAf2+55xhJFVI7L2QpvwBdzCJOVn
j90Rsh8zN0DEkMkRnLMJKm7fOcjSviMdV5S8InCz6ZwekPPMxcfXbuo1BYyir7jG
0Kaivm939qC3cTPqhjZDs3tSHIj3Ofh/X+0kfo9GDrvYnQ9NFaN/COsTPBRHKul+
lIaiZXyOxnB+MnjqVa2neolhtDn8FVZJSyPAu9CC8jq/hP3UiumEOY4ka6LzWb5e
MFarExvTORUhYVh/PST13M2dr/ROL7UAEHmX/1tnKkrw1QzG8ar0Y6/ueK4j4X4p
pIHXGBufBGuH1QRwESvmq0iW3lE0caHl1aAKhE8/jJW3JThFP0Fh8HfM6Ksl4V1a
rl4JHQ/439Aqv7k4QKrfJZ5rEZ3w8WuRXn01kK27n+nJF6BGR4CfyxLAJnTHmvIM
GITVnagfliuj46oSitotp5Uf1Vmengel6PhYiJJsoFl53GisZPCJX+p1imtxxx1l
FSUYMAQnMkPjKzXFft/99iA2IYHoruBEGH9pdPgpt1JQSvokj74Dja4Bq6Vw2i21
J4PABnD4UT3r0rgzkZB72LwPKmB/faHTXWujyFMAPTtVjtfBf9j5FblJYMSjA089
127NfxiXM5dYveQxQZEor3TvjTPXV6uwjOUwj/7aSIIjtHhPDhReyjdbx7E2HzDh
Gc/cSingGjY537PfD/x8ffZw4bThNR45j8N+Yy7nec86WiyUfGBiOHgOwI52C3fe
BJfbFjemnyzIMrAi+KcYZjvpdUTrN6w7IWwOOFOUYtOHWqEhQsWr2iZQgtgt1+6j
KkaRb8Ionk8asZym5zfdosfjjpLNnmKVDbP3F67v6hg9A/R7cOmuxMN5iuYtXfV0
6JhaRjs4B77NkRbaSpkkCNfATwnD9vXHNqZCaDWKeGdNQjyeNVxBkJjtLzo9Qmhb
nLCSzWMnlXFURnlkOyfA0+JvJ/HPgiQ6ysdYBQOUlJDFW/wgA4NS1D38GcpXyjd9
VezOBfBaIv2bvcRVR5/j3cNotBuQJVHg1rsFMn9R0hUNGPjq+mfa/510uCZZxFI9
17h7L0YMo58L8+PwikiQI9rKyre63M1U9Z4KNPkqJv5OJsWzJ0sSaK5Gi5hrtvEc
2P/LJ+HeRk5QrRveqKrN0JvPUdqMZbz40SB8GITh5mGv9yBaKRxXW18jmNWAd7om
zaYwf4irsM0jAX7nKQTjwnw4nvnSjq6V8FVzRLxbgVuEQkIm7i/kiub5z7t9g59Y
yiEpEOoyOf070j2a6VgKZtPP3LFVnR/s1gKdzmcNVI9h39I+Kc5ygdYEGClIqIkV
jT3MTJsAQncnEyCAjpikRXrC4TmltbKps6RnqSkNEZZmPA73QTU49acDYyZWtKVp
fkwQMJHarKV1NA4M4oO+zJhgg7p+GRkIti/khCzVSOEzYzXty761U4kSUhfKIHsM
dDTxqYLDE+pqGdQc4uWddTRIJk+uBzd2l8L/zL98yl7OQbYCp3uHC52luy4cxTkH
sa826Lff2w1loFlrrAyaXf2niYvqTWy0LPDYY5wRKeCSF6VYeyebBOm1NIzrh2Vj
Jj/QzR1oPylAdcGYXT3D8veHuFV/fF7eLQwyBfR/H8sBpd6ok41ZadfOlr4eogn7
QFKoyYQbW7eunpmdH243yCZBnG8hRwKA9nHfchf8RcpN1bM+DBAeCE0ujuVwMojc
qLkYSRR3VNiTwoPjD41X6R7/t8olLAXLgsaHPGcGxbcj9tYmRSxOfNwvmvHhv08z
dpguNZz+OdBRDDhbkdKybcEPRGFvA9C9QCbZyRZ2wwuvIc2eCwIsldh76xUF5GrL
RJf6EERCevCarJa4dXh1Cb1fF4ZshJa6/OrPI8f592+n7bi3iNPjluxcWjKWarNn
Vx5vJyEJ6q3BjS0MNGbX2vAH+qb81fVCG4GD19KAoOhIzqh5Torfd3P3rxfxh6HF
EZqTt6GDSBmUqEEqy+fCIqiEoRDZBHbV2D1n45V+zZcQC/h6DGGkX3TsHbnjQId2
F/OPkTUqvD1XiEXtjtWlGNDRGJlT1+WR4PGdyzA7tawpDRe5f7VUEJ6jrr4cigHu
9bvGeEqyL5y1YUeTHnI8yX6mYWNCgDUYyeDO+zXFJfVuxcvz8/EJVCanXY2g0rTk
WnjAfazeDqSkC0MUMIN5XKvtresWWyRUiFzR1VGbOmkfAbHlC0IkroYIZRsfQ+Io
5I3fJwHCCOiHpmCs4mHuxZwxf1aaw4nsJk8Oe2EhhMA0ypb8uNTj6mXA7U3+xLfu
4vNLeiXCw/AJN/Rf11FAl5ZJhPcb7mzl3Rv0JfPiFFQlB5RN4JPR2yHt1kBAdJ71
ESFNOSCvnnXjDZ3+U9E7XKle7AEuh/xzlVtte1w9BWnwroMF9HGUGQhLHW9WvLQb
krY6yMcKhXedBy6WUATui7gXC9I87skpFr7P3fYmqK/29RNsABCIx4yUaOPFKVkn
SdV1oQbkswxe5SZ5o8lXM+Pul+lnERGLtPnFO2QTtq16xoxUW5GJRGW1RUoCnDuc
dlV4vHgs6L5uI5kBUz+OtEyDqjeWoQo9srnbcJGPPTl+ganq1EP0XtRRzzFofF07
XxGoCgNMKv2scyzRAkxCW8ccbzMzN0Q7eQgUEc8G+ZjvZ+tmRaCF/BmKlLJs2Z87
B4hX9y4+U7IQefDuEzpaNIGVR2dTuEmexYIW7tfOndULO6QX90MJ8YbyhKARqavB
mFk6IsMcfLn8U8EyPwtFtuEC5GrrolNZLpsxRl6nIdyLfnBhU+zJPkVDe7NR7063
UFFwMuoGgH+Ipfhvc1cRDXo1Bmfos1zhCPi+DrGhwXqBhKvwBgS+rqRBAbQ+i3pA
AoZDdB8fM5Xz2BZJSJr/ek1GRR2tNl+FbGQ6nbe+wosdxQbotwue2bNbvbaFSJoZ
ueavVMs7nLcKQI+bskZfi3f7MAPSJ7Sow1pav1Jk4r52vujxzm/IwRiwh8DdZQve
GeOUVOnrvYBaVXCIVM/kltynQbjY2ee3meTyVT7pnIEoghcZCy42cm3zvgJ/BeZ8
U2f3TE7Jl9MWCInKsMG6hPy6EyRbCPtRMvEhgYppH3opxCzemdPv4uV1dZfSwVcm
g+wfhJSc60y3LFAB8wicVIgDO3NOID6jcWrS4d4Dk2IkjZQlKFnAMKZBQwn1+C9d
1vyKqww52BFN+4Qkf8FrxP78uXQXQVvPoK6v11TR2oogUkQWW15q/ZsJOtNjstM3
VylUia+pzLPXD9rO9qx163QD3Qehv97S17e84Qwt0vGB+O2gKnSUAypbiirKkLTv
T6lgBYwHGHetpIlrTcaVB5MPe/ye1PAVPG/4VuZsaa8rlgDptjXb3bUuadd2Rbxm
B05YmyKBr/kuxxwnGBl/OYS+vCnxALjoLvYwAv6Kl5ZGQq0FMr+72xkZjzn+8FOj
z9wX/O/3u7a6TLBR5DMEsQprMnjIlwyr01VmWUwjbMHxINOLikTNt66vREaNpG1B
XxyxJ69j85cRrf05ZsylLw6ln9MaUA6kCK8qFQ4hdsO1J+v9XL2KMDM8Rsk/Jckw
irClc0o0vjmvRh6CFAMvRVOtmZWhWuVU6SFpBLVigV6UmlhgJVOep+SxdweNZsCj
sbt5O3weqpbK8FQoJNQeAQ+TBrprLPTfh9rT/QSRczSgfrVMJU3sZwiumnvSJ3/n
2eABLXYLx+VM434EgWOc6Ey97SmcLjfiJopb5xaGqYw1JPFK/WmYqlMrDnWc5aqL
Ujif+pqlMIMStAc4L/5dAJqkaOVEazZzzUMsf1qnT3slPZGoD4F1oXM/bDrHe4fq
ukWlqbM2OihBpW3XLqITvYNk/pTZ2M6hqSsblH4gQb1VYuAbuOLt8fYAQTi0MZoQ
hBqxJ3uHakhNroCC9+OlVZSZI4D8cTNOqjBqqkOZe88dIce7fJ2gUwKCKGt2DhVk
dP3UYfQ+eL5hCeGg31m0ZQ33CHtwLQk49xB472eji8o=
`pragma protect end_protected
