��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�Gf�`x��S�.Ao�vZ5��]f��;=O~\��3�I���Y~�l*�/��:��By��af@O��6�J���Co�58�׃�x������1��DcC���mJ���Y��Dg?��YV���X�
Lzig/G�,AT�[G]�
(1с��-��� $^��n��7@�6(���D��v'���0-l�o�މ0ޔ������D�SF,U3�>���	uY�i)�֥������'+T�t���3tk5���3��9'+"�1tkg��p�[��:���_ֱo�����:�V�sd^qP��~²bd'���X�����U��=)�%�"3H�W�������z��ܷ5:�U��G����s3��YKV���9-)��6j̕�tP�?�1lql���;5-��q��	���s��v۶J��`�S�h�c�	8)&�����qTV�뇗�~����¾ǰ�5Z��L0��4��;�
"�B�q>��${�[��� J��7\�� )���&���w��I��t66����a�=>��2k�/�u�\��ijԬ��={�Ԓ�c�D�	5��-��
7�䔏���Qw��՞����@p�bywI�l �ɮ������[�MaLOg(D4������kC��r�=��p<Dߴ2t��5�S���D���IzOA �u�;b����|�Zu���Z���D��ZiR4�E,�E�Y�����;J��Slt�R��b���ì*�c��Rw��&�F�Gu��^�1ߖN�/e� ׃1�(�I�K]�"Z�-��p�����v�[2�?�9e�t{���>��*���]|#�,��v��%���b�����q���\��l��?�Ќt����5� MI�Z��6��>�y�����PA�:ם	�b�G�7E_V�(�ٴ�.=���S��8w8�q�/{jч��|��_|#V��3��'�ù6d��*�EG��z�r�Q٠�=���Uw~�ߨ���mDT�+�GM�\]��@y��U�Oh3�u<V�0�N�<6A�k���̍�%jZT����sxs]VDMt(��K��CN���?�ԙ{�n 飕B�\�\~�@�L�Gd ���ͽ��&mcɸ�g>��[��Q��b�AC�·�!F��h �ӷrG�>��r���J.T;�~��Y���M���YK��n�5$3��b4��
�&^��1n���h􃉑Fh��0��4�V��>k�]��3�N��Uo$���ph#::&��Ef�]����+e1c	e�IdY�!�p���gD��>4q�uގI��cOP3㫧Z"��LMG ��o��2f�v%n��Y��ErK�0C�v�}ǾD���Zfҳt}������W��u�Rǃ����j��%��2$�r4�-��2�x����iX��~-�P��r�E�>���^�]��@?�i�5$[W���O��O�	�NRm��#�����r<��yCu��D�[���+��<�rA i�ʲ���PdɆE�z��r7_�;�nUҊB�4��H�Lg;û�T�'����LS_!�LH���ŏ�Q��`d��6w�������oZ�i�1�P��ˀR�q�U[����ҢT)�̕ʕ5.WrC�h�;���k5�Oy�h���+V�� �1���Qp�D�p�-�м'�'�A���&}q�.��T���ڌ�����&�F�j풆a�����H��0@P����"��%%�T������~��i������O���[�G��PTLL��1^~(�^���]���,��vu���~���e�굢�tڻ
f�Kfm��{ۯ���( ����A�ѕ��xM�nbO�h��(��_��x��U o�<.�y�0W�|^���f-�~&�4��� ��\w�K�ټ���5�����\	C��WҲ���^��'���+ώ�MF��"�JfU�����5��+�FO���������1���3G�}�?���z���['������"+ 6)S��� ><�u���Q��s,�C�5����놱s��Z��[Ћ�Ɖ����Or���'�e����i�!�yk�,+���$2�w����N�<9�O�+��
���-����3�m���O&��,�L/r���v*
��'^FV���t�LQ�{6�a"]4 ���s�Y��l���셴rT,R�$��cM�'� $�ϓ�b�+���f���[E���!�妱�c���NH�ޚD�C�3b�6����SqS�7_Ф��`]�Uf�,ǰz$����H��f�`��H����oCg�0���9G�*X�}s+��<��D���9ࡒ7a�wG�$p�3U���jk���P*.Qk�G}�x�����s��"������!����
m�H�^$�Zv����u��Ɔ�Z4���4|e� +�M�5�'��\�x}�l��o�ݔ�X�4�>���L��0~�.�t_�,��7�(t'����ۂwW�C{�q¨�k������Q�D�o���ҿ�'X���̮�&��@yå��ζ5NS�fM���f�%��o.r�^5�o��HZ�N�Oh��`{�ԣf%W���{,�>ᴔ�&ѥ�Y��(A~��TPl/ �,�h3h!�7|\Y�6�W�_��pCy]W�;5v$[��Uj�ٿ��ujt��%3:da	�s�SAl4��R
�.����/>��d^d�{m�?���������y.R�7���1��<���+��F��_�%;r��N`J�V�Ǻ\t�jiheu����t:�F-DonG���<X�����r�P���>�mX��+/c�آ�X@�,�^E�(N0^�JBA�>-�-�|�6��RQ�&�q����jǃ{�Í�b��Dk>�3����й�n}BѦ~42t�/�3).&��$�͆2<�,��HHʥ}�j��n8pJ)�*ňK��b���с�K�<��%`WHHø�>��U5@vn'�{V�uC��}�uC�j��L�=#@L�OF?���D}`�>�:�WN ����\�;��OB����r��>�.dB0�Z/{���NBS]�̥��7�J����{��(S|��o5�c�R%� K����,�r�&���"j��=%�����!b2%k�O9��I<s*|)ѱi���TY|R�G`J�����׎�*�y�+��u�%�����<�UfT�"�Z���hvwΑ�og{0��X�
��֤1γ��S�1�f#ϫ)Y�|��Fׄw�<��L��J�� �J�u�U/�)	$�	r��\p��~R�)��1L-I#&6Nj,L'�.e��v���Ʒ={ҿp�.�فU�*#��:���'�7���3��X�mX8�|�����X�&?����0Wރl4�QKC^�Nf	�C�~�ώ�&[(����H��/��Onk?�J��� �
�% ��*fަ�r�Q�j̴}SKo}g<�g+���Ϻ���k	���<��>�(��:B$���Ԃ��I��9�X�e��/sW�����c��Z�x&���.���\��NO{R�<Ï��l�C�x0z�NҦoos�#3�5�*R�y_�&�0�;ۊ�֎x��gg&�?��t��Y� ET�3�"x���`��>�l$%x�V������U^ޮ�٥"��`�Nz>jO�;�o9F������İmtGSykP�GH$�M!�F�C�j7�$����Q�2C�4�m������b�G����p;��}<9jݻLz�g=r	�n��hh�m_���i�<�����1��D2�T3(�a�Q%�pst�l9�D�-����>U�z����T�`]wX�Is�l�a`Ce��.�t,�3�a�%�)�Q̾���U��ݡ���|J ���~��p7<	��UP
K0��'~t�M���r^$��~�&4t�z� �p������[�V$��0kI�a��
���5�L�B48��T�K�;���έ�n����.��mhI�?���@�޺�`R��쮳��Z�ٻ��C���95�Cm�H�t��A��1d�}�t�ŭ��Є�S�a��=(�Ѥ�Ѱ Z��&��Y�)g��qԗ�BpZ��ׯ��)#���t����Qkj�o9|O2w���$w(Z��� AN��g����ReBD�y�:RMƋb�)��/w���mhڟ
	��a𦣺->�m��-Ӱ�>ȇ�����Zi��)� ��\/�g��^�%��f�/�}Y��p[Z���:�1��&	��Gs������B�W�� x�T��۟�8�W+>Ď����HXRߺ����0��v���[ &ٓ/�Ơ͘�̲��G��F�z
�c�P����.��즌Q*����y
��T��h�~��kAN��1�l��"��Se�X�H>�x���&`�f)%#�)�&->�C"�(߈.
4�[4k���	���5��VUꫂ�x�8�Q��<o<�֓�T�U�m���� ��"�p����1�����'�@*�,Zy0��9o�\](�7�o���s�P�0=���l*0y�q��V���t;4o��ܥ2��� ���/[^KPj�B1V10��jΉ��++7�kCM��4\�G����U�L�[*G+@Xj/�;�Z�n�{�[��ݙ3)�y{���?���0��p^�$ ��a?N��|(���;x)��3��AL�=�[`���m���AZ��܈2��(�[k�}ƌ���TC��-��	&���q��$����|��Ii����P¿��a�d؁��1�*w��W��*2�Sb��1�>",�悵i˙y��_-�v��q@x��#�~V�ˠl\%-:Ȟ$�#g��k>5�(`����^R$iʟ���g^GX�q�[�h����
�Ȟ�h|��js�c5˭�y���g����&��/V�C[���+6�R1�C�71$Y<��fb��G2/�E�}tN��а�J�"�&�0Ґ��'ߞ�",U�O�8жL�r�W���;~�+�ܤ?&&5c����Ǐq��Ab��h?oK��*"�~��K@ɾ(u\"�bD/���h!�����&BW&\_�-��FiJ>��T*�]X&# :��-�$켗N�����	�DM�t�`Q�����7�X����?���2����z��_Aa�a����&h�؞��ˎ��/�_�y(��TZ�_!$�oS��mb_mo�lt�B��=�-�܀�_�H��ZDizM�=��f�'�P���_�5���=�:=�qrY'gd�}#b��Tqq�4c1���3���h[�{G1}�kׯ��ä
p����E�x�}dP�f���fY0�WVd�ێ�\>�'�ѐx�B��b`|"2%�HQ��&����A��)�3d��
�t���q��
ł1��z��QnG�	���2��s뢑�o���=�8	���0�jjjp?�!�m�F�=Nl��tH�FM�O'��/0.VL��@l���K�n
�aG�UGф	M�ŝK�����s&;e-�N	���\��r�H�|�TF�[��Ze<���2NrM=��a�1N�{���&�ӥ�S��D-�2�`��Y�-�����^:q�ڬ��)�h���wW�]K��ag��5�:�2��fIOf�Lބ_�ZV��XwAW �5��w\�Sƾ�M�s�{/a;�$�ɵM'��:!�Q�6K��%�N	�6��_����9�h���da��?);�v��W������`]�Ƥ��F;�)\�^&���˯){/�V�����PJz�����dzG6��@#r��3��)B+z�gm� ��X�<�U"o���Q]�$���ע@��Zr��������;�x3�lt�u>�4�]��lo\A��T���B�����V��%0����]R�/����ަO���T�Y�s���2�j�B�ó(��l*L��A0L=aS�z���LW��i���Z�	���Gw�g=N�n��'F@="ykq��v�r	��KX��j�@��{��4o�G����6�#�(WƬuJ���
�n7vi/UC��ѿ� iH�, �V�Ll�������s�������A�R�`{����2�����:x-u��������u�@N˵��F�4P��'����[
G$Ӄ���L�pw�h��T�R�������b ۜ�����)C��[}��nx�N��¢��x��ӽ��g�5*��Rs���0������8w�����N,Y�F�2�I�^M*s�NU���wU6�Kǽz	ۉ�a������Vp�'� � J��NBX�U6.%��(�	=B�\}h��G�}M[`��|(LA��{&u;z��ڃ��OaMƞ�j�ϝ��E�����?�Mi�*�#� �7_�u1h�!3�$.p�ᦰ�b}~n��D�~R�toH�ٴ��~��l!�G�	֡����v�F|6%� �N�Y���mI���`�\�ƣM��(uJ2�O���,��s��H�D��:��zo�����$/��0�����I�*�h?0���̣ipf*>�ږ����PҶLP{�U�Z��B�t�Nϡ��r� x��	,:}Z���Nx����%Z\�| ǆ����"��\YT������q4u~;	��A���*$�:�2�`�}�>*c�W<^���j��;*|�|-�u�݋U"��S��ETe�%i+���Nb����0:�TM��V�c��N��I�����Z(��7��]�G6�A��+��uN�����dIm�CWC5����3"X�4[hZ"��7,���U��.96 0ڭO�p��X��	��ӎP�[�]��Gq	��xr,���0�Z��HRϢ_�k�F�he�nv_�tVD�^���dq��xe�\\�L��P������j�'#1F݄w�EIKXXq�mA%40%B����sۧ�@�G�!F7H����]��-��ϳ��͗C�n�����z���6�'�h�U ��{ͪO�;�j�{��<0ԇ��\w01h��h�d�b��ѹ/[��$1���0Pj� ����X�`r����n)X>_0/��;�l��ysЬ��X��R@�Do�M)ar�7���o��	1>E�������<f���S�
�,	T�,
"�3� p:mr6΁���~ҿo�1�zj~ùv��ɧRj�������[�ҮI�=���%�l'z�Q��*Ì�mz�z��0x#��;����V�f�Ƒ�m�(X&�P�p�~.�*��g�,�|�� �����,;��g��P�pT���#	�mke��jL��?�����h��?����=�)�ǈ�Z���LH��8�����'��&@
a���Ib��h	K� �I� ��^�9+�:�F@Y�2;8>�J�blH��¡(�c�[�n!%U�T�+���`��t�)$Ր� ����>�WS�< BKZ�㋪z;z-�9��#����9�8A3@.�_�n9��������>��j�1�e:9�)<�I�w�*�}��.��?���c�2QP6!����I�#��y3����_�rِ�]%����]Н���+�YEB��f8���)彀�d��0~}�3y�ظ��`Jۨ��s��A�y�f#]�ûgճ��ϵtv=�WM(Zi~Ѹ�3���sIxg�	��v�׾x\�<nU��A����K�}4����C�'�	A�5���>�pQ���Y"��)�5.�s�OϚ��vO�.�g����T�ل0S<��jx�����|�_HWv�6��,ǴJsi���հV�Kx�X@˱�p��StIA����iE�3c$����]��J��^b_�&z(Y�13\ V��F�D3ph�b��ۧI �A�������/ʌ�	��4w�U�C!]��@�R&If�r��ׇ����@ZgF�<	V��Tސ�~;�I�,>��e&�PC���v�1`�ZT`N��u�o��y]�A��rl95uDˊ�6=���I ]9�T�|��]P$I?f��n�-�-Oi�[�ڋp>Þ�j����;���Mr��7�b��6�ȃI�&b���3$��� �����E4FU"`�"}��0�t����^����E+����n�eO�%�ܔ|��\��a��N�;�2�o�'���h5Ǩ{��d�h���)�Tu�хW%����#)���O� Պ3��?�#�!w�BIUs�G��s\��գ�0���V�.]�32G�$b�Xu��e�%;A6���x	X+[�xg�������A�ʙ�����Ʋ�L���Tef��=AI=�����8����L�[6H�)MSm�wX� ��Ut�S����V���Ф�$�P���C�BNw�;��4hH�ܿ��c����Q�?e�ٳ��l�A���P��&���`kB�����8��c�����38x���G|��]�Eʇ�S"���b�f��'���`�z���*�'+$��8:w�*�ذ,J��P�]5D���������)�"\�m"��^�KD��O�~�/i-�{��q��#���A��NI���)8�����Li�d1Y���bz�-��\�V=�Z�4GbEZ���V+��G��S�^��=���S� |f�ѽ-*���,s���$ԇ�#�qpU���Ar��o��oT[���x�l��7�gP�Y*�م��1	h@�*Q�����엠ۓ_���d�g5�/8B��/�6�ލ��[}Ln�m'z`v���1�S�y�j3v�h�<�xB;��<'|b���:Q�q�o�`��6�|���Yυ����+b�j�9fF1w�3��]{��<s������*2� ��� ��gqن�BY����`}���%�pr{g��`u�a:39��~��C����FNѴ��i�׻	1o5l��RB����!��ӣ]g�E&����?��V�DD㛊s<�p���@�����1�(�ܔ�H�_w:=�	�u;�2�B�H���1hع��!�����+3����2W��9j���Q����7J��P���d�
�\�.�����R�y�l�&c���*F×�����H��<�"��� �=�Y)!�*�`�W�e���Gi��E-�s9�.27��<]R����|�T)��a#G_c%��~��tbܱ=4ln��,:$ȋ���Z.�G�H�km:'��/�䍣�����|`;��$ ?�+?�.�5�m�����"��ש�N��&�j�A��.�=t��Zr=<�I,(�j/@T�������,�����m�O�����P�Q���
M�WN�=�.�,/c�0A��'�X�q��+�(L�W�i�C\}P����h�)Zg���:��^�>i�Hр<���d���(_�p��P��x����m���{��L0΁JW얾�.��e�y��cK��n.�v�gśh��y��1�U}+�B���J���5��[���)�Q�\�Cob�Q���06D�O|C�=J�\kC���I�l�{������4�N�q��X�����Qjx�`�������{2�AOr畳��q�(F�7�omRf[o��cu�R��'�%�J5�y�������/F�<K0��O��y�B:v�S�!z (�n#�1A��aSShfp�ړ���ɎB�,Q���IϏ9��cP���� ��o�ׯ�
@�@�#�?�R!���C�cb[��s�l�PG+{�M���([I1��L>���֭+V\����ˍj�SU��=�ie����:`\-yG�AW���x�1���N�߱/��p�G�3��f������.1X'q�,���$g�K��l>ٶ�)�DH����$�@���w��Ub����M��<˸�;�`�o�k��$Kf����9���eY��(���p�8�9g9�"��Y%����8�,��ʐ�%�p�e��%�Zw9��7j��l��,�8�}��\~�J�e����Y�(�y�^�T~���;K���'6�+|������8�r��X�����-3�}=�B��/i����g׿K���ݡ�y�C��_�0!�j$=(�r���]i~'X������N��-_�<�Uw�6�峘���}�+����v����VB5�k>��yD�-'oǷi�*@�H)�j� BQF�XD���5�1��K6,�kQn�����A��ۙ""ܔR�/�C�:���j�^�W% �į׼��\b�gK2���Z1�L�(T�UU���ڠ����A��l��X�h��a�4s�.����Q0�*	�f���!�����]�8�2�d��]�,q"�]��G�/�BdD2��$��.0(O��jl����(H�	p��J�U��
/�1�cXҞ冨�h����g����M��SJ�N毹��8����W,��%��ps��c�bq�YT�{�<�(q���R�*@���4�S.9#h9�߼㵨�o�̠���d�U�3}-z[�!����M��26v'���\���Jh"a<"Mt�E�f��^}L��H��G�z���KA���k�����>�$��/��*�����7"5�Ȅ�OQ���x��$��#�	�����W#�+�C~�$]���-x»��b7��'1o�Kc�?w~�i�b@W���%�A�7G��F�OB�`j�di|�$��D��Gx��gɮ,e$!����m���b?�J4m���F��H�8T=�f ��������`qCΪx��-�����q���O��恍�+�	�V9P�������b��W�����i̴EЭ	zԞ���95����2�/!�z���Zh�WCX�>�'�g��lU��,�â���2�
p�C$�6��3(|���e+;Z����O�Wm�/�a:;���PgOU���B�Dy��$;N�@�6������.���p�/��O)�K����~�>%l r=_3E[��V���ιʠ/8��2�+\��V*р�K���&qR7'�U�NNu�X��굇<H�>E�����yd�t1�dX��Ҋ�A�lϐ0z�|�TJ��r9<]͵�c���I�ѽ��i"�p��F!���,s4�O��m���W���R�Ի���m)��.�23r"�	��E��]ݸ����`9�O�z�Y��Nj�����t����`�cb�Cֿ�5I>�5�[�Ԓ�a(���`1Ex#p�r�|^�Ľs�ԫ�}�#}�p�%,K3^�O�ys|��h؎	�h5'%H+�����X�~z����Î�3��L2e�@��j��h��q��}����/c��v��Z�����$7q�@FU���+��bəH��8v�1t�+�-����Y����܃���,*�(~���Tu��i+�` k"�\|�[��f����	