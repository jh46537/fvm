��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���q��՛������@�oa�R��Iz1A�#`�ԀP��Iqh�3��F�`�ҥ����c�
K4#����ge��T5��G�z�4��R��\3jU�;Ѫ.Xq��d���D��nmac��V�ܕ�;�)=�(?0�י+�k�襮=�%�YO������鏷w��>�s]��6�t�u�;]��4���!����q��
1�xF!b������.����\�2�X���`���~���4�k2Y�a�w�7=�E�u��#��_f�g�:�S|.�� �֞/^���J���,\*��p�#�0k�|
]c(��7��ȩ�'�Q�	�kR-`~���Zk8�$'��x��A1����Ko�� _'-l_���\��
+*�q�k�����V�LZ\?rŮ5�xwpP�V�22m��w�j�{!��;�Fs����]U�ӂt0������M|��L�{U�o\H8D\���í���&3C�#B�x��h���G����g'�M5���P+�@�K���Z�T1��	�ϕ>����N}t��l�tCfSݮ�U�+2T�S`�DV��#�y=�����/xn1%s{>S}|�R
Fл��YA�VCr�q�5`$֋�\QB'��oq���>��y�H�mS�>�}!G%�B*!7�W���ۋ���{QJge������!L�>o���I�Zs|�͸|��vW���rY�}�A�yPL�Uݕ87�]�D
�v#��)�S��}i�vZ1.�ai9l>f�0���mFX�0^�J,Q���O~]���o�[�r�{�?�o]R��� :k�8C";���RF��re���`n��0T����O|S,S>W��c�yf�VrvC<��Z@�z�84�3Tn�HN(5ǅ]iz_�}teνh���+7�!Rٞ�n��cz�M�P3�p�$Eu~KgNܾ��ۨ��\fz��,٬���'5�cN���f�VNw7ߍڿ/�A��o�����x�@�T���ѣR��	H��M��R�#��>.w��7�vR����O�}�Y~Q�mF'�&�}�7th�+LB�M�D&7	��Ec���?��B�6�b�9J�=t�{l�M����B�����9��Y�"EQ��k�:'��wHa;s��>����16��	߇!o&/�;G���yubc[�𔈹|���Q&Y���X���N�G��H�x4R�[�����nh�;� ���w���<yA��JDk�<�N���jB�������;�5�9wץ��l"sc�]U�
�XVP�ןn�;�w(�J����������H��s�����c�6�$'�ݾ^lS"�\6��=�[�8+h9z�3<�$�l��k 6��G��@��!~M�nFCu[�a��h����fr��[G�U٣�7�K���&��F��)��+�B�m��\G��`���]ѕ� ���=���
Z�C��7���=���䏻-:�K��v$(���=��k�#��<�lg���D�6�G�P�v�^�C��R�v/����ӗ�PڑĢ��E	d�D�?�%�f�D�!�����-� ly��!d�N���.`�x�'4 �"�ף���~��9ݥ�hnJ&���H/#=���Z24%~��$��n�� 
� �e����|,�V{��T��@n`�[}�j�*���c`?y8λ��iD��v��MRh��E4�&��nih@���}��ӂ�~i%��Y�H�@��N'|��)�ĩK�KD���1~�޸�L܏HW:�? ������};��'Rx0����
�,W.���K��H���%<�%e���w�HW�gPsN5!��΃��_�O)V���v[Y�}��͒o�g�/��G�Lë' Q�ZP�+��'����+����tF�"����������㑆Q� b���E�.64�ʼ�M&�r��8C��o��E{�ph���D�%,"���y�2�Ok�Q�n:��/Z"��na�X,m�AAq��=>ػl�����~��-���τ����6�E�["��Ƹ�^S�_��dIPݞ�-�0�"�+�e����l�l�t�d���*����V��?�XMD(Ĕ���R�<r3l6?�t�H��ԁ �N�UF#�8tLF�8���bBڀ�͵�!k�ǇgA�w�����F�^��9^_@�Zҕ�"���1�P�lVʠ�+^65�{��]R��>�ʇ.�"C6p(�n��D�s׎�`�6|kk\N���raRJ�T�#RE�4�A#�4*$�c�ѱ쌓�*�~�c�ws9k���g�'�p~��c��hG�ӕ�Xzs2?U��h�cd΂]+A��ydYV.�l�U(0~��C)'�:�!�u8 =τ���\!9�uN��E:3���ҽa�>�bg�0� ��������NW_'X�L� �\qD0�q��0�r�;T�JY�2L,#I��M�Olr8 �����������t�~#�eѾ�����bLYF_���Z��!�\���_��@;�s��3'������e����ǩ:�?_�9�ÚP�kM;���	 �m+\��Î���|��jy��bG^q��:5�����B���|n�>XZ4Bވ�x�*>T�󲳤�Iz�I���ޱ�+Y�gE��8P��v[0斟]�����[i�|���eP���A/�~�`�K\�*�0�J&U���Y���y�fUx0p܆�������kY�||\[7�Al�1����-�x��Be��@�a#t�|�b�U�&Z8���Q���B����\O��
�������[��e�6�?���	9�������|����WI
���	}��2�e�T˥�j�0��a��->������!�IL��4��F��ؾf�x����W9��Y�w�� �C�G���h���O�]�8�R^����!!��K���5%����a�6d>��GqZО�?�Y�00����D���n��@=��rE��?�ޑQ*�>���Y���x�+��Sv4��Ց~�j�-�M�rا��G�F>�j5;nV��sH]�ٿl��tI~}�?	W:�l���Ծ�#&�-��Rx>�^��<� +�p&++���G<�4y���Y�Y�S�K˅�`�(={!�m�Z� ~M��IV=#TNܽ�����;m���qg�w��9��X�!��6�DW^��<F�`���8��J�Ձ5c᪔�щ��Y�ž?�9
��b��+bt�SN�;���Y&0�^qK �ܦ�h<�)#{���/�N$���88�f���Il���w���=��Ҋ�K��f[�����3嘘�I�(;�KH�e#!DCt���o��w��mw�\$'�P�c�u�²�P�
�'���؟o�I+�Z�pz�D7�j�9<p��1v5+o5g�e�$A��Ȩ��F;�<$�=G5�<TD8��G��3�e��yV�v��z��+,!%Zp�+���]�4*�,��:Lc��b��w�2gO7�Y_V�G�X��<���G@��WSo�Q3��A��ӿ����f�v{�lg�jB
X(��ʊX�V�p/)l� �1�v^>���	$�fv�̎�h�tw&���'�[�ZҪ9��<k�J��5ˎ�����>����ܵyb�R_ �|cn���6�b	�����i]�NY~}8(z�BP�1��,���Z#� �7����#m��A}jC�g��= �V�	�ј��G�弋�L<m���/	XR>巍��>�'zdtՂީ�~���x9��:e+,�	7�'����*��P�Cy���X�F�[��[.�LE-	����ތ�%B�$c�γ�56W:P}UC11D����}�79�E���:X�Oqw����fG�q�&���T����ؔ��N��Rւ"��F���Ys�$CQ��eX�S����!�M)�=��G��==��¬+�Ȯ��0Uy�d*Q ��\�:��[�P�RLH�f�����h-�{�q�)�A֓7�]� (���R�M2e�"��#�*yh%}��~T�]��XD뮶@T������-��ɪ���xٿǳn�gSny�4u^�����%���8�O�^� ���&T-�Me-)��6o����'�����҂=���h5b���^򭼅]_B��O4�ߝ�#�����b_v���6�����FV���bZ*����h�����$�Ф ����&���\(g�G `X-���	�AE?@t��'���5��ɥ�\��O?M��'�I�O�W]���9>�����RT����
�	���}������ q�)hX��5��qs�7E&{��P���e�H��g�r!L]��R�S�n���� l�8�o���d�=��F+��#�-;�[�60|�	u��"k��J2�>/o/��+W��J@�|�Nϧ�1�+�L��l#�ol�0�I�`�+��[�Y��,��ځ�c�t����E}��#/[gzk$�d�H[��:q����oR�l̠�]���q��ѳ��-ب�z������~��nk��}��W�ȅ�<��bZzR�1�"�0sBi� ����`�g���_�z�����1�UfkǑ��
W;7��{=�hX+�=5�2��G�d��z73o�
 �Y� ��s2�����z���ɅUOƸT�l�@|�;R��/�i�9��niOcr�4"�Ks�ZWv�.�\U^H���ph|?�J��'r����7���A��g:�SW�_�����֢y�nQ*_}�i���?�6N��*�&�o�%��a|DCS��z್B��k�ʘQ�W�C�l��m��j�� ԛj"�K
&���H�g��R��K�5xA�Qy,C��)W��@L%����LY9EoȀ��<�WN�f�&	 �C�B�����?;nvA�Q.����8Y��Ez�u�-R�����x�Mm� �&;[�G�k�����ܬ�^����g�#�=ݹ힆�b�s��9
�tI���L�m��n�ӄ���N���j�}������d|�nV0/���(���w�81܎҂T>��=>�9�-��ɴ�7	���U�X"�����r��a�}�
FCd�[	~�Y�\
-�'�jc.44,Jl�+���fy�#��	����{�Ý�C��Q
#jz�<�C�V�pmi�,tvTi�5&W��T|�Ez�!1@�ەrG'��B���s}Ҳ�'��Z��:��e���?/k�o�ʂ�`1��}�M1J�QmTgp
r������E�'��5�w�'�!9t$����(.?DlH���"cBT�KIY��!yx�,dY�{��)�|��y�#(����X������5��-��Q���S���s7��BD�1kG�P�G')˛��gȝ��C�Z�ՍCI����A&x�)6&���W��z���
gg�jn�9��5�Y�F>�F
��ӛ}����$��|
͞���I;UL��EHۻ�)ueTO��
�Z�VsϽ���;+��Ynލ�8%��y�Vt}�}����â��=/���պhQn"*�+������g����$ܶ�yVf�(�<����`�-��_��fR��;��jΦĒ� �_F����ES6��Y�EI����Ċ�G���>��
*��^+TxɽQ	�ق�Ϲ�2��͖���v�-�4Ka����3Ry�G�V�-M�"�x9(a`k���`=��A��l�ȩ�n���:�8�#�u�y����T!����S��o��C�'V/J5U�������N.�J��R��><��"n@�*ɧ�й��sa������Z�1}���qw��M�jD�hI &7}!Q��/jЈ�w���H�8�X��� ڜT���ҕX�@�B��)bMD�҅�����Rɝ#d����1d=']����uڪ��R�f�Y�VKP
�|�l��,v���Er�ea�D �}�X�&,p��&��E
��%��������D�
�{{�9���o�.Q�l'�z< @��!�*b%j8*[B�I������5�_��g��	t�����bz|�v��CU��?�F&�Q����7���0A�˱��0���Fq�򲽈�E�kakS�QJ�&����օ���5�%ޒ~}���x���3�a��\,|D/��������6�^$���^��t��$��^CY���VM�ƃ~��F�
�%,��ﭯM�j���̂Ƞ�z�Vr��F�#��/�r�B���(��k�e��V���ZI��{��r�ϔmʴF<ු�Fs��ǋN��l��$�
���(nm\�!wjDaeGѻ(�����P�������V*?i2謚�;�#I���t�̠�F�j�0ҟ]���=_�f#:BXZo�B F#�³��G�����4n}0w3����G\ds9ɋ;�<hI����p<!x)��{�z�e]z5����$,�)w�K��#���v�t2�{�݈0t v��1�"9�E�����P�ݘ: S��,��c/�v�W��B�<!��@	���\j��	�VM �����_Z�1 S:X[�[�����.��<wiG�ܹ#�o��܊�uŰݏ}�_�<������)�1�I�5$Տ�m��3�;�ź�.o\�����<q�����:�-}��������me�� a����kt�{uI0�P�J�p�d�L�z��rLo�â��ub�o-�va�mD�F�*���9�Ĭ�h�=pfw^u��	ۼx��U4,'�l;5��1�:�����hC���ݠzt���'�y�w}:����%C��<T�m�U g^�.�X����2���R����UrW��~�|���#&���(���J<Q���sD��p�§���O�9��Ȩr�{_#"TB�sӟ��q
��c���Y}�/��&u�]~g�[, V�%l/�
�᭚�i�V�=��ٜ�q��H�Dͭ
,o�~k�����Ď�q�-"�ܦ�����t��B��N��'�Y H^#g:^i��ń^-Y.�F�h����{�XXRKK�`�� �P��q��M�	�`��6M����W/Y�B;| ֙�S�V��Gax ��f�DC��[����ެ]�����sX�H��v�N�o~S�u1#�2q���ng)��+Q<wH����7V&i[�g��c��I�u�$��<��˼���⑎ɔ���L�A�)�]���(^p����f\�Xd�*걪�3�s�H=��>����GA�b���OCEvy\�N̸�"�B�� ǐ���;F�4M���`��2XZb��D�-�W��K��3�2��ֺChJ�Y~��B�\���TJ�x�ǄPF��L��U�vā�Y��bl���	������]��x�\0�Nl1�e.ڿ��w<Q���`�ag���ȸF5p9����2�ф�}bB���1*D�G{r/��x-Oes��W#�~_���B�V�1m�����K->��rӓڡt,C?���)6����k�"�&�����W̐o�� +c���)�������/��ڣﵚ�����+~f:U���r�J��TC���qs���'��fLe��������-+<߸�BI����:�H��.uҳ��������ZX���`�]����Y�su� ��/b$ ���g�;F��%:�gv�}Ԅ�g��K Uv9~��z^�շ����-��>R�f-4�v���5��<=�%{Γ%^Y*9+bb�747/��|�$Բ�������*��_��?c4��ۦ��>:�?��q.El4���v�3�k�Z(£��tD�q�d��7�>V^;�ډʘ��4��7yC�g7ĉl�הz����g��x
��}��h&�S_��)�SA���@	�,:��Uλ
�������d�|b_KO��B
ۅI+vQ��Hɮ"ȟ�:�2�O�q���2H-���q�)�z�d���6'�O{�S�$���^���D�X�����O�i9�1"ߞ��~*��.E;�����)3��|�V}hlb�f�	޶�Ȏ�`�@�N�&M��n@W���f�FЖjc~� �G#�\q@3��ޫNI鉊f���c�C��!,��کa�M(V����/6-����R�uL��RW��&������#�ݛ�և'\���%�ė��Ck�(`g𐿶��+�}�YH��&���m�-���zA&pj����҃�Wp��I��k�.ƻLI����������M?%Nw!s03�F1k���9P���ԗPJ�5�H�32b�$n�+e�[�Ր�
��U��"�؈��/k�( ��݂��g��F �F��D�T�Q?��H��Ћ��֬��~v���b�؉Ne�&0%�^���p�-�j���~�(����/���2��0�WgnJ��Ey}9���w>Kx����t,'��9X����[.H61�ŷ�5G����x�yܿdr�<æ��(�"u�-��o��u��`�-�XK�]ñܤ���B㬷~)Y���~G�ĽeٽD��%��|֢5ݗ�;3T�	�.�hU���Y���H�z�[��h4�7��ʅ�7NN7tⴾҝqh��&QX���-�/g�8[ar��z<���p�E��`��#q�"Db$��Ig��>��e�@�����[,�$x��R�#��֨j������q��umژ��,��c����2%�QS�{�z�ھm7��o�y�7ԙF⫟�Lt�63��R�@��;�p���.`��Z��%���$L
u�rS�NmhF%��x�F��1���������֌���ˈ�Vq���F!��6U4�]W�<�} [<#:�O W�̮��Ȕ�!*���b�\\��߈)hu�����>g{�f5�"�=�ɽq�(����3�� �_&�%����ȴ�����=��:�%�-N�f��On|�o�J.�hzPEP&ꒁ��i����0L�A7=������F��[[��\6#c�6��6T?q�+��p�@��MǥVY���T;kǀ��ݞZd� Ww%���t�iJ�\�}y�/�$�`���ŷ�#5_]�����yg��)�E��&%ca=�:�o��jD7"�NEL��o;�����d�QDUh��.1[K.�(R\
��k�# �>�4ߡ8��T,��3�l�#���X��m��:�!�Ʊ�X�`@`�B����{��zگ��:�T�j<aJ���'�؞x��?�Z}R!���:P�t�/�LB�3w&C�犨+h��:��r\;����_3�����H-�N�1;f� JdC��v-D�QԬT����|��SXrVN��L��K"��`ڤe�Ͽ@���a�$[SO^p@�W�A �l�ӥ�
ßt�va+b�!:����9l�G���B�m���M��/�1O������(H��/U����J��72�j�5��0x�a�5m�0}9� �A�+�Gٹ��@~Xf&������D��@-˫���]�Yݩ��Ɨ�v^�ғ��$�pR���쎯��R�թ!T����Zg�IM%�^��AW�D0��}ɼ�ZpW��
S�
g�aE�Hkem����zӳ䖹[���*�]&?8�����a>?{hߕ��ED�F�zѺ����v�
4�c.��b��	m��N7��Z�4Q� �QdY���L�`1������]��l�w�,<H���W�b��ߨcY�^�������$��TP����^@�JC�|���O��<��MlU�K��Аl��l���-�v����j���S#�S�n�h0`L�R��T������'3	��8:@:����[��\9����6d �NXMØ�AW�)t-�������H��*Ð�e�)���	B߉�:x��N©8vI�'��0?�aD�6E��qm�F͐��))�Tw��Y^����6P@��%	��W�� 3��i�����3��P>�jc��)�V��٠n�M�ٜ���a{�<[ÏͮF���/��������|�a��-�)i����Ѱ� ���:�����M�ӯ�Hq\v�Nn���N�qC��r�-	�d;N�"����F����mL_�>�q�k��}a9+Wx kQ�$UY�n�\��$��I��xp[)x�����X'P�M޼�pc�+�6[2\Yh7�ej�����}]�+V�D�K3ޮ%��֟%��[:_���΀$jNw���N�6.��Rejj��Bu~���O�ܮb[���9F�aۿM���@���_�4'���� �6�6\8k�s:Zc�&�'��`��R7x.��3�P$��h��Y�D��7.��Ob={w*��z�)A{s�������d��:���$�Ô�"������ݰ�� ����g"3�`�!�����w$��:�nԒ��Nj�������4i��~��R���Tڔc �C'כ�qL���� �~���sΒ����Nʻ^yAIR�d��ټ��b�A1�x����M�-5�'�:�$��R�&+v7&�,M�(ה0j[�]S�W[P��uW�9{�~��ܬ'flL�	�bP�#ڰ��A�PɈ��Kg���X�L��0D��t�e
&J
���y���v�ћ�[ Ǉ�~@��JuZ��]��P ����a1DȆě�'p��%�(:W����y�)D�SBi[�|�[K��%��!�x����*��G)u��N�_��`��~�`!�0��+���[���!��Z'I��h�P��Xĕs �U����*����B�gR��c�E�ЏQ`o�����0�!�����aލ�ؾh0R;���J�ǅ��e9�E��C�Q����YI���p�y��K��r�h���՞'�����v��Ύ2/�>n��3\�5�ӄ���Y��c1Q5fp�"�~l�Ղ�l��<Q����&_�\�i���:�|ڶ&69F��Fd�ɟ��A-J\%m�^�[�Vx��)�����D`a�e��8�K�x��9� �[��k���K����"�Q��\&��Sqʀh��7>�_�` ��7���R��6c��$�0>Y����Y��31�+�t�kp��X&��]�����*�4tyP�B�k����⫣�Kt��3��X"�΍}MT�����z��l*�_�-V�"t~����Qb��'�a����o��H���3o
��&�sv�t�$&�n��e���"��F�=D��]b�#��sb�_0h"�P��6���������WJ@_W^aC����R}w$�B�:8���ނ��gpX�aF�I�����L��H6��9E��N˦n��[�8J�����0������������	. ������x��M�5�.pP��|��N��1���pF�C���������M�Z��ˎs�T���MB�,��<�/Rq��Q(�ʀpL� j��V^�$P�9u���O����g�)d��@tSG����|l�ć���s���'j.�q�z
��#�[gj�x�4�]Ko�a)��(�08��z}�E� �����~��[͒�t�cweG(�]���2	�j~ű���pXmg� �[�)���	��n���
 .�0���rٳX������=���_���q{!�lI�@���_�0�6U!<Ǒ� ��`m�獥,�rQ��V�0�
�
�y������0Ϣ�{���a������.׀���?�������q8��Dì�������s��� �z9�����h���NyM�z��A���%
̆ ��RZ�������釿�d;���jv7�)]���dB��j�b�6��h�/�t�2���&]���ѡ�2�փ�`��F��S]]���ra{�1���mTގ���=�0�ߔq*�tk�?���E4�N%ә�H2�>͑cbN���xw���s�a�qy�֖,��DU{���q?X�hVJ�#G����<5�/�"�Xd�5�mІ�bb;���?V��V`KoB"����_PчZ�V�M��,	iz
:���R�ß����U�:Nh���@�Y���g���@%C���(3��[�­h��vb�2L����[�-��`� +�% LP���?>Rb�� �m�����#�Ch�萉��:{���4��	6��+���~@n
W�8D ��1e�3�Fn&���uv-�W��!N`�MgHB@K��l(�[e�j�(d���U\�318h��d}=��cO�P�����<�m���9\9�6UDm�Kd��#����Zwv��_�hY���^�62ɤ�m��q�x�/�a�t��Rs&!���4_-�x�����)F��0c�*���!I6�������(�E��E���\�b�:�z��I7/�@�p�߬N[�婤+I�W��#�q�)O� %^rG��U5Ա�ښ:�Z=�B�|��d����{>�.�ۙ����/�c�6$�|�P�k2sC7���d��ĔW��	&�v���nC�F�F�J1Q~�����׉�E��6y� ��|�ehC��V��X�-#m7:ߺ0��-"F_U@]m��C��z�&�'�����D���_!�ܝ��-��T��D��eN�'���
�4�f���ϢI�U^������&�q(o�?I�{i�����Qu��r͙0�V�jJ��Lo���"�h��,ii��47�( ;�'ٰU���Z��L��Qӧ��;|U!
�+D!�c��0E�˃V0/}�� �5��Ue�˕����:� �x�Q؅3�������$*/�<��3ٕ���C�#�U�7Ѷ���f\�Q����2�]Z�i�_��,�Ҹ��vK��̝�Q4���^8�~)�fj�o�)6��6\&tM�5�/���!ר��?�{/�R'���<�`_����C�(��qeA����|�o�����l�����>�iA����B~��kT+W{ܧ	X��+�PN��0�'Fsm�62��(�I���%�d�.�`��"'ˮ�x?B�����[��u�bF�Fr}�.�0Q�	H2@s�l���^7��u��}��<HD|('-(���dM��Eᣩ��\����wYK�rݓ�SB*�#�y�6�P�@�ƀTs��b+j+A�NW���3�Z��JEk�����X��y��niԸȐ�O��a��E��4ލ��4��J*�I*��ه�s:�Y����Fs
��v.��iGyřB��%g�����{r@q�R+��A$�T�sU��X<T>Z$^�C�A/�Ɏʿ�Å's�<��Q&}�R�6W���e|�
���bQ�Wvx��mą�����k ^�<����s�͉NtW��T�1�B4�-�J���*7l q�P�2i;�9_����^Qv�ʭ@v�*�N�n�ܻ(��>D�7MfE��xe�@�nBZ�I2F�!3���}[ �GS��k�{���eb�Z�#O�[���*+�,�իw�����("j��ӻ�b6J.�Qs��P�[�⒐�����E�wI�V��R��/���yUT&��G���O�+&�}�_ƈ�����_{�j+ ObC��������f:{��(�Џ�[�o��HӸeA�TK^ԛㅃC��@k���;�,b�?8s2�N��'�i]��"��O=?Ǫ�WZ`���	\�xh��	�IL�J����d��Jr#��oli�"���_'��V�mҜ���2��4�&y�{T��������&ݪ6��Аv-ŕÔ��H㛡�8x�b�ca�q�$
��1m���Z�m�L���x�ܶ�w���ɪ��g� N�F��[�,;ml�� C���d�|���Z� �'rQ�EஎJ�7�w��d�bLs������±d� �:���j	�܋���4�XB����գ�ϡ���j�k<�����E3���!!�յm<ý}"`���o��ß��ی�5�Vpȋ�B-�;����] �A��H����L�����l=8�P&A=�=;�O�?����s�W�p��`�9X_�x9�Q�"�B�˓�:;ӭ?��t钪�h�r;w�������oB�
�iN���QǶiU���|���|�n�b_��W�^o���,�o�2���L`;]�Y�����h&  =ÖB����B���=�+$;��Z�O�6i��~����I|�޴��$�!|��ue���,�z�3	~LR��ϵ��Xs~�&�,s�އ"~S�0����������jBl�b[*�?+6�UrMT�Ø`��«!����l�9��g���#$b�c·Biy��B�9h8�n�`aן�k��x!E�w�@@!�h�W9���;np'����7�ʹ��*��S�"WVD���������h~�N�"���_l����Y�N	K>i��dy�S�k�_����I���9k>�̟5,��@�t"�M�h�����S���#ku�A�"2w���2j�z �/�Įi`�S�Hx��T��6>�mD�2b/��� ��n
�,��g�I�������=�:�|w����j`����:�لx������I	�|�x�
G�h���滼��	$s������H��\2��ȈD��q���N���̴�7� q������	i�E��%~���`ߋ������GʞA�k����Ћ�c�T$?�c���������f��;^��LW'�.t�գm"HP�.��0�m8��d�kk������*�:w�{�?�%�G&�^��L'3�r�M!��M��I�vg����_ƥ:�Wo���e���y�\Y�@��`X�|A�*m]B����Q�<u�>����Nm����WЎ��aNdD�1�~����lK�Zp�"��7�I$W=�JpB�d8ƶ�E%h�r)�k�O�pQ���mYI�d�b�P�q�yQ��^W&�����A`���c���{n�W4���u�>A��5�\\ �6r��݅�@�_��MJ-�so9��)�\�ʷ����}�G�k�ʘS�X�v#�a�������p^�e���`��o}�R0𞫹����
�͜/���=�;0�V$��#�+��B-�z��+u���!,�%A�y���vɅw�߭�O�Ɛ�����y�`�f`�\K���S�R�IQ�Э��J���8Grh~t�1~�{�!����)��K�.���+ʗt�������jJ�YZ푢��6���"�UaH��A��{W�"�9��ݫKd${�Q{˃9��W�ʠ|io�}\W�i�F;w�UZ׵����9"���/�y4,[�м?�^<m���.j�|��IL���;;�,K⊬F����.	� 腸��d:�ü
u]#�2i�=D�r���sΌv��1b��^�����Ooׂ��'m��=Iw����z1e�h�FTj��w�v�xn_�i�jT�X�9ǎ���9b&�#��
	�=5��>5</:�
#�9I8c�W�Gxݖw�ݛB���E��a�RY;�7�/$!�:Ec����Z���A�e?9�bJ�/4���Փwa�K��9JE�ՉcpwT�б������_����1�Ò#�x";��#�C<k�h%]�ySʱ��ףT3svS�p��OJB�Rs�M�6fCvߜ�z}^�c�EǛ��=�d�s��( c]<C>J��4���K�+�|hZ,3�����Vq�|�!l�]]�]*��G��Y�CC�$+�E��-l۟�r��;��n�0���LP�y�j��	�8��)�ٗU��J��jȄaf��ע(���+M��z���5�&��;�����Q51��l�U���v�>�(4�a��Fz�+��)Ʈ��!i�Ś#�[�Taj!���/�(�gL�ڿ�O�ζ����$�@�%��͐/�� �O{C�'	+�w�M�"9.9-����@i&!��ԫ�Z�Z�|^X�����D?��Z�-�,y,�_��&ЃrP,E閈���7-���ƃ����WD�C�B�C/���^�K�D�`�!��:�j���[��;�|��p����罈�G�jqI�]@OAr�,�U�,��_�!��tڠuN�~�!�$��gd��K'��C�<���� U�Y�m�����l���d��L�Q��\�s��.P����"��i��7�=���5��z�hYO'��D�1��%rz~BP�Q$/��@�e��cl�N��ď͖M��Aa���2�Gh!.8-w�z��Z���C���'��^����9o�bp~H�W`��S��Ğ�q�� ��n֖#���pP�RC���?������[̛�l��7���
��"�[qc�?D�f�������Z��,�mV�t� �fth��e�Tn��WB���5G���S���^���"lm�j�g{Sn��1�_J_�,'Ⓨ1� m_�B��V�C@o6����ţ㵘\��f���ʘ�?*�"�v�V^���{��}tn�	���~�|��d�\�Ύ@�I��!�cNO��N�����TW��59ЈO��Ȥ����-�����H�s��O+��L�b_��c���|�q���;���_��"�O�Hk�z�:��qO�-��^]��ʗ~�7�������;E�e�AwTG�"�� ����5���&嵽�u�$�4K�;# w�Ñ�7ss�z0�>��Wh�����\>�,�����-<͘��N��3��V!v60/��9U�ؑ��r'�Z,s�����ޓiM�ø�,��X�\7�V�~m��H�G�!�J�A� ��.a�q��a��a���o�"_���Aʛ-�����h�rO1��>���U��	[*0���Zh5R=�3�
��+����y������:��M2�q�`�+k��)�$a�jj1�$X"j�[�Q��G�Ҵ��t��q���J�Y�&�Ay��PƼ>��r >�r��%�2+~�<���yMrV�E�9��,�{���}�QS�]s�$�슶�������P��ayщ� ���P]��I\�����f���49k�����'���|���V��g:Ϳ!H�(�Qk��+����ב^�|ch����4
e/u@.�Mm9��>�����G:�g����.+������yB�mJ�m��� ��<����Z�d�	�T�i�d���?�~1��!����R9\��װ�QQ�����}j� �n�%�l]�q��7;P�u���|}C�;���:��"� H��z̞�0|�n�9R���=kn~7�q{��2ɚG`&<z�c���]�Ϩ���&Ǽ���$);04.�t�t��(ihI#'�������t�y0w������џy$�n��Ο�������
&�����cy�wk��6䩫�ahD 8{ĺ��"���i��JE|1�t�\��ճhjH�������yH����8��g��-�T�6׈r:�|�(�y�A/;z%�lg"c����l8mg B���YV��ɱ�h9�r	� +;�n���EG�B������3�>���N��+*�vdɔ��P�dGy���&[��rˤ����+fl�i: �5����c��a���Ϙj�6���n\�O��"��!�0���GÑ`��E��*$�ݨ(�Sc	t�q�(ƛ����pjj�w�����0��LBA��7��T�HCuB��"�y'T.ű+&��VF�MZ���G�B|*�ڡ?��Q�s��}���n�L1m�b��R3�(fgE#�eɂ��۳N%�;/6Hsz�SLz&#SOVAaYo�����܌ނ��( \�KŪ���Ow����t�0�sv�+S`XE.4[� ����8����#^�,�L�@]p=�qܨ@���v�& gSO%8�4��_�9��6Q��xS��z����;Wq��u�)���Q���$~�+���W�Q�۫�p��T2�k4�e�3��Άˇ�.�p��D�.^(0��,;�֬��SҐ0��x�C��oW��VA³vWϳ�`�,�ڤ8��{���K�����������b�'o���vn �85W��Z��N����9���jf � �T�fR~@��
�����Nz5������)��H�Mˌ2�_�=�M��i���IG�sy*"m��_,$�,\��7�m���e��V�&"�>��;�	�+�5�y�*#蹝*����;�Oyw"n��O=�i���e�	�FF���TD���j�9 ���1�ӻ�aU�m�x�b̏�hC���aL��gU�Į���X�}���ʵZ~*oQ��^4S!(3~�;Ur -#<@��0#~A�������������D9��&d�n�a(|�-��Lٕ�����i'�/P=՟ ኪxm�@Nj�-��e�J$`��q�"���������kB�+DT��O��>�<2�:D�[��;�Ώ���;R�)'7rќC�$�#rE#��@�_���K��l�	>�w쯣���i=^��`4A�P9���u��q�OG� I������$n�!k�T��⌳91�o�*���YW�Ɲz>=�(�w��f�B�S{$��P��|���Ō1��V�/؏>w��x���򸾻�8Q#��.N`|�[�u�F�����	��KE8 �]�`Q��nXd���؟^�E�٧�Y~���M�1�,��{Q?G-�����fIP8*[���U"�x���.�s�~.����.���_�ze�a�K���dV�AuǏj�wh<t�t��8ꔍkA�N�V�*��O�}�+�?.O$��Ai��1q�Z�9_�8IՃ�t�3��a�߸sIZ�+���`'���PF�zHqU�^����t1jS��	t]A��L��#O�bAS�n��{��uT$���z(Ih5u�r`C��,rhֻ�v-'q�je��,s�<�H��z�ܤ� ��۲Hu��}�**���ǲSv�J�
R�.�^�X�sHb�,䩮�;DdAp����j��+�����)d�|}+@�������[%�&��0�]+V9w'Y�=%��1;;�xBJ>��/��'�����(��4�a�4��7�u�s��i�,[��7 �wm�IK����7����£&�1��6��{Cî��g�LI�
y�	ו��%`<�R2��X�r�^�e����5��I��V&�h~�iVv�Ih�-zQ`	�LÆ�Xm����I2��:!�� z/��q����'���~�߀+�c$[��=g�`�<1��X~���9D�Y}7�5�)��S��fj�T�D���葉_��Vs`R�;��֪t%��jn�TI�"����B79��4��M*��l�ZU��2sj���kN����5�C ��p�ρ�ahԃs(�M�Ov����?nP���׿j�VP��(!�
�z��J����6yG��ʺG���X�?�q'�xѯn� �7Q���#��ڥ�������/t/Q~�T�W�?9��!_��c��kIp��'�pM|?��}-�_�]A����JPg;+c"E��&������!"-���w�S�_���~�H�A*�Pa��4
�\�$x�5+��[���R5��W�0�t[�����<�5٥� ����k�i��D4�����#����
6�Xszd�K���������jFW�̽��|O���*������q�io�E�¼��;�͈l%���~)�c���>�pK��K�à�R��HK45�/���]z콣�G�P�������{�p=JH�9M�N�E-��X�!fՊ��O�.Y�`q������(v��.%�ƍ��F,�~�������f���}6vgz��@���28𜝆���O'j9�A
!&FF��� Mx��홚�>N7��z;*�wA0�o\�
��W�EN;�Q���TX�����Ր�L ����w��mo�Շ��k��{�E7'��pc3Ed^���QBL��{�U����sT_�/X5�\��>�������(%�Ogr���LI<�6�E��E��8u�1G���?$:.�@^\v/�p�(r3>��F���*�&��ʩz\9�ٹ;��{*�^���qR���4��/�%��Q��2
7��5��|D�X�wYgI�c07��Jbc��a-���<�P����2��,@�2���ķ?q�;/�Q ��@�P��YX��N��|�q�r�^���Du/y��%E[�����W)��&����%���\���4 �L�p�������+��֤z�&n�UU��`��I�1��`R�>��-���	I,W�������< >��E���B��[#;�)��5z�5��"T'D��ڈڀub1�Sw���A��[W�Hݷ#	�c���I��9�-M3�xH_����I�U��_�H��Cnzg:{�fWa�;/�pb�B�V=�C45��jӀ��r�ۮ�Rhu\7��B������F�f"�yv-�Ɣm�Q���G�9�?$i�ڰ?6��{k�U�PO���3~YѺ"��t�.�m���(kqg"a^��6�j6{Z�k �"0\��:Tn�Uhv�qn����l����:���VLv�o�� �C��bt��i��@��($�DY���}��u����ҹ¹�����9��#�U''�.=m%u��Lq�!�Qv�bd\,�7<�~�B�)
3X������+!��B.�7�\b�)��\�Ҏ=�����aD�^$FQ��]j�љ۝���{�Ax�.�f$�c��r̗�$X�sf=�ʿw�#���E((�1"u_gk]����;�oS�>ʞ:R7���+�����<:4ڦMs^{3'�q�^Ry�v!���dz��u�9��^�f�M3�e���ck�����H{�ˋ�#,c�DAy�=:m(w:�Vq~��a�CP�q'L���@ǈ��M�)���x�Q��P���ڥ��Hp��FB�ڶK�/�Q�[)A���1��9ԥ�ɱ�zC�1��v�e|���J��v0�F����s��\�r��d�_�wË}a���ɒM9������1��%i��� Ĺ�{��Ӏ\�"�6��:o &N�����E��gD��E���*����9����N��8|��Mc3��ظE�m7ꑢ���Yfg�Oq �=��k\���J�a䍜�Ҍo�30����-�`��@iTI�r�!����:���`Ӡ�2;�{Ԟ3`�Ѻ*O։��~x���mp�熿)1��[C�����r|`�t�&9������.~f)���^XNMV�	x?�H %��N ��C��{�V�dz't��DshA߉�,��X�i��f�s���Ȁ>IN��iC�B9ê�l�:�6+����^G˸�׼�/(���E	�}L��9s����&V|�M���6�S���5}����0=�V�dLb=��������O���ÿp#R��퀕瀊S扰���GJ��Aȥ3zs�iA�ur��֦LvѰ�"�M�@���{x��GӓQ���,�kz넃�&�%�Ǭ��Z5���h~����.�r7�	�x]�����<d0�t�f�I�iò�K_�p�YF}��m�D�;�l�Xe��~��V��d+������^O���D���:�Mk���w�*	(���RY[�a�K��T(�7/G�=�>eN]�[#�Ua=���̄!˂�j���3v&��4���9o������7���O�3r���Y����YP \oV]���;T�F��Y<ӈ�8�o_%ޱ���
�H���a�P�!u�K~��NЬ+����cq,|�Tǲ����7�b����aک�����C-��?����TBq�B�{��� 8"�w�D���p�:��b�����F+���/��[���C��@����ja�c4"��U����W�h���O���,Z�,�ʅ.k��'}M�H���3={U��y+�8��7W�]96�J�xw��Ȯ𦞀D��jL�$!J��G��~د&sXD�M~?,�lN�>��r�gP��J]��N�8~�q��n@�r�i�"˱�Ј�������WiB��t��}�1�3>� J�Q����zۈ$�w��a�^m,�O��s1�w����6c�o�琵M�.�>):Oz����k�x���c�!U�km��l�A�Lq�کvQ���C�s}ԥ�B����|�䃕�>`gu:�G2A�,æx�Ό��$��W�bp�$��#(��Q��{��<٩}��5�0`�I�G�����rq1X�*�/����.��n�>_�����F� �G(q���5*)
����T�[��,�}�,G��!��0xt�ꬅt)� C�|j-�g�34���~h"�Q=Z�j ��d���KEJ��=l&�=(����ݬ��'�1�ˎ�8FP�O��Bb��d����}��o����͑7�H�z���q��B���ӻ7״��}��~�N�eH���|g��D��b���0��r�*�S(�06�C�h�ЭV�e�޻ ːA�n��$C���<�a���̤��-�P�1W��AW^��xSe<�Մ�K��C+�
@��U�A�j>�"�US<s��N4h��ߎ�0�R���M�b�o�2K�������T�����1�<��?�.�:M��)�(�Z)
�u('�B'�D��a��ۯV(�'���=go�S����Q�1]^kJ�*�����4����=H����3�dxa�i�X`~�G#�=c,~��N-���nL��\1��@�M��;�Z����[mB:��#�o�1�X˨5L}B��F������_)������@#fp����lK�y�\���N���(h��������]��z�{�����-�9��X0�W�a�`"�k
�R[��5����B�s�C��Pp�B�1�S� 5~'z�����|�x_k�P5"��@}�*v�%�|U����%ώi��e��:��������8ߐ�8f�4��͙�c�?��Q-R��'VSѵѷ�!I��M����M����_|��� ��$��%̃��9�90#���٤���Z{�,��J��z�)�i
F�J�����O|�V�o�FM[p���]���(pC�Y;�4"_�i3tg�+@+�b�����P):*���}B/T<��dK%K �N?u.��<��N8��<�z
�4�'j�T9������^_W�H�a��a���c'z�w7�V��zp֋N�<Tj�(A��"�d]�x'y����d�+F�5��ct�1{B��~:H����pSH��`$���f{���>�H"F��!�W/z��ؿ�����@Y��6��V�����J�	��޹�B�T#N^��Ģ!��+N'QP�5�v�ô�V��7|2�u�\�u�VߍK�Nyd�P�.��Ҋe�\��:;��\u�#�ۥ;ƙ`��ʬ�rO0��/���yMW=�����_nxB��w�߃�U-�J�BƟ �w�78���!�=�࿔�h�����ח�1iȲ�`K����WHk�ћp��u�)å��o~Q�2.N�/���V�@_�ğ�A�R�8���1��fn����d�H!����?�,݁��B���!�(`����ج\d�we�s���Ϭ�5�V��ġ썢_��V��Vr�Ъ��A"�[=W/�~�����R�z������J�`�S,Fh>v����H�cn!#5ᴘ���P�le�	o:��"�آ7'D�9����Ө�;��RJUT��}=,��u ��xT���Ǩ5�H%��t���y7ML�p��y�Rd7�_(��_O������2�� �H��\�5�t��-O�qC4O[ջ{����E��P\����J��/ʯ��"u�� �����Z������ �X����0d�L]wQ8�{�y�,<��?����p�m�z���1V�
uJ�|��D���������\�`�r��i����&P.͉�Q�O0��0����Q�W,�A�
�0��:�.7e�H�?iv5O�guԉS�Hm��km�Cq��y���D�o��@�=��$�en��Qomr�l! �%��NO����:��}�O�E�s�?k��֠K��H�]w%�(&
�B6s��B�C�|���m\�˽~��m�\��]i�0�4�B3�bT��<_V�n(�C������κ��.� �M�����Շw�R��I���T�����\o�Tm�ד�
�yR�L���<�z���;�����v@�p���o�Buz;dy�)eQ:g ;�3�j�l�me��2�g�*�nL�i$qM�� Z��;��]~��*�k��e!���a��;��H���.�L�$�޺��l��(�d��`'�:��>9�����{��bʨxt��t��"h9~�-��p�C@ΛF���ֲ�la*�ŉ�ܕ��.~l�/_&�bI''�Ճ)s�%�j�]�Y� QQ9ZY��ٟ�ȹ����k�DNf&� ��� ��R�)K�1s'H��÷��Ԩ�q/0��|�d�e?�
6W��e�ڊ����I�#W��ќ�)<�"���|8�f*G("�! w�k��<ۖ���u��%G��ߋvǷ�/?V����o_{6$�hm
�A�ܕ-����i���R;����0A��7� ��o�����R���+��x<tv ���ql�A>���m0~@�{��Ւ<���D-,�xy���l+E��6��X/��Z��+��ā9}�ku
�'�/�����V�7*s�3��=O*ю��Sdӣ08w�c��-�%0.5~�G���~0�c��%8�ɴ�u���כ�~�@7�����gJ9�D_��C���"�i����˪�Y{eԒ$I�?M��Ѡ�B|����ƛK!��)#��v_����y�X�=��J�n�dJ!�)[�Jj]<���il���e�Gʜ�;̾x;�3��)<W"�ʵ\�	�V<�𷑗�����ݨV�ۡ����h�7�9���c��I���I���₇O�����b�V�:g���I2��v��閚=So�o��g+B=�t�6����Ν���I�r�g�YC�p�89K��/�x�6!/��:W��y|ڹ�Al"|�ĔvK-y%��0-j%��W
����j���?s�*y�$�Cgq�L׭8�	T<=p������C���%_#K�҉?����~��ZM�wX�{U@��8���G/���>*�ȫ-8�Ů!T�a�׍h�e�� �� M����)�ʫ�슨J!�Bl�X0gj攜�V#�^<^��S'b"�?����V���0������n$7���E�+<�u��R.o܁�d#����S�¹�-�<����k��;���W��0�W������{)LP����=�9�����#	�"�E�R�Xk�*�ϻ �T�������u�U��%����oe�5%�Q�G*�F���H*Ȯ	�t��G[�Q%r�=�b+C�5��_�/�U&���Ռ��HJf��L���6IB�b��`�il	����� �=`�P,䌋�҆��-�i�{���ԷNsX�v���	A��3��C��s+����'�V��:��e��2��_�f�������&�j�j����y��y�CB�h���~RO+��c����e4	T��N���܌�(����!�W贑��{��H?5?��;��מ�T�3$���I�������t.6�Nk��t�E���FJ�4�-��t`5]:����s������-`I���Y<Ĳ�������"r�A��u2
��&%��X��a?�LV%�c�1)��`�GK���9�Mc���o���:��,M�1R�_)($�}��_M���D-��;QT�Α��O��y����L��"W#����&�`�u�`�6k� Y���AP��IIC�,�4h��4,t)Z0��0��(%�V���Wo�q;�,�\��͇jْ�� �4��0U�����5Ty�:tqYk����҆��l!�� �b�0<��AU&l��!�_D��!����qP�V��[�9Q�Y���Wm��Od���I5l�U��}]�i�V��m�DQI��{݀�^��c��Q���{�Nw����E�B��o1Va�I�#��}�j�d��B����	�p�{�7l�~:��=j����2l��������tH	{����3aRtڼ۸(v$����Wd�x��.���0N�<G���T��g[a��*	�[����$(o1y�5�H���O%o�	��_Q�~���>ҵ`ܰ�GKR6J�$�F�������xT�F�]v*��`ԣt3�WӔ0� <~iT:��0T�g��U���).����]%�LTA�2��z�VVb�8p
>�yW��M�F-M�ӽ�x�T��P�\񅒂J��4v��G�N3.M3k5��6dp�H��R��	�����N��x��i?�S��0�#g�sx���Yo��+��ű�ݳ^X���G��'���.��ƚ���eX��t�Y޷X��z�,��Dk�����<���@U�	!ehQ�\<��n��~��	���.!�Va��-C��<��s8��*e���l�!����:z��1AN��"cfO^m�i�fLz�/����^���4"ڴ�Su���n+��wt�3�F�Ǭ���4��u�V��J��1���A�~ic��z���a/�9�G����j�ܸt�@A��ѝ��A�Q�F =��z���US�r=փ���˜�M"�7�j`g��{��^[��1��c��B~	m2�YS�ՍM��f�b��a���aK��Y0^�RZd\tU�)>\�����%��̋Z�J3�Y}���}e��u�����o&��kD� dxk�kL+���ˆ�� �g�?[vު�� ��*3�ԚC�wO>
w�@f^/�	���>hN�������#尶�q.��,4͍4���`�׋��q-��?�NL,���cj����p��㰧2\5Հ�X���l�|�X9�A�2�i1��Q|�f�-Gٵ��|"�L� 9���"b����NN�Us�NW��Vn�RQs�WX�HU�iA�+x9�2ע�m)��!֛n:�f����������A�L}��~K�R��uP	�X2C��mק��mk��Zd��2�9P��s�lTe�6�+�&kX�!��x�	(����q���[�X�_,��F8�j.̣�įi�	Y&H���A�T�q��CZD�V-�h��粃�{��EF#]<5U���{�蹹e]�Ŀ�ЍWt���+h��1ʻTv�4
JD�y9����[(��!@���v%1J`^)ּ+"Wc�2�(�z�T��k�*���I 6շ9��y�#B�s�wl&3�d�;�(��ak�&p�UX��O��y�ʅvi��9i��%�-������^�;�y�d/�h:� �����KY#ի^j8���+B@p�!ԃ��!(�?��.9{����&shyBv�J@t�bn���i^�m
B���f���"π�&l�`j��%AW��[W.�hC�R�Z��>��괒g�a�'4���c��,��;�ȷ�ҋ��9ڬ�k���&8����J$Q�?�ĕ���CH���6ng�BE�2B>�����kI|�rG����5!m��k:)���׷��/F\2'��q�Ƕ¥�Ci-䷤�	oofAv9bώ5w��e�y�94qꬢ�2Fƣ��MC��Q���s0v�ś[o_85��sK�ȴ���O����F3�z���[b�K��ԙ�c�ֈ�/�dA�m�RY>ל���UX�-6��o�[61���� ��W]� �h�V�'�t���:] �b�1Q0"0"
2꟏�8�J8afm�d�Qx!��ןU�t ����_�(�f���A[6������!�w��έ��F�H
�W�
S4JS"���O�Wؽ50�K�K���D!i���VC�<���o0&K\J} Z�q���p��	j�!�ˋm�lp�#^	Twhi��dc-h�2
\�,���Aq+dX�ʫ`*D�x	.|X~ˏ���k>�55���<?�[hv�Iq�{���mcWE������
d�仜rr*�A�z�."�3����P�}�n]���I[lv�vJ"�55?��6f_l
0��v����4��Y�2s"&ؚr,\���)k�)<��\�u��&S(U�3lK�#B�&O[�d��9:>ο1.0�������!b�4�-�����@��10s�1�e�5�m���PJ��b���Suy�3��_�Q�X��$M*�f��Zax�UQ=0BG�s4*E�j�4�R��� ���"��\؋�p<�$��S3B�w �P�<>?�x��X0qڐH�qF;rC�Tߒ�n��l!!�T@x��Æ���e^�б�}$9'��ΌXLrPa� ��Qk��&	����;΢rh=�hz./��T]:���r����J�hg[Ҵf���⡥��:�[-k��+eX�*t�U��#�;���U��e��F(0]��k�X��ީ��m�b&��@��_��>��4=����<��d9��m$R��O��R���U����f��s�d��&��<ŝ`C6�=G�n�V���S���.F�-X����ӻ��?].�{<��;�V�D����>�D�,A҉��i���>5>\tK���(�_5m�ʲ�[�������@��R�F��PL
�m5�J�9�J�1�r�P�O>I��l�O�F-{f���Ktve����Ĺ���,%SxQ�Ю�)u[Z_aXv���IE&҇Fs5�BP�\r'��/����`?H�k9�:ib�҉�.�N㩉o7�Ί���MR�+�F�[U�O[���?�	�̌�t���񓜴��=vv����R450n�rۏhh�-�� ������0雚�Ճ�Y`� �0x�&���傷�K�.�!�M#����Bo)�M�y��k_�o�3��5��b�l(%c��#z�HUD����GJ��^{�gC�N� �QLB��e�9�� �LCk&9}�\�������
,,�	,E�{=�9�C΀� ���{��*`�'��|�X��g���C�m�2������W�ֻ�$_�#+��&!}\>F2�u_A��~23,-'��S����M<�hj�L��.�
Ǘ�z'�`����*խ���+���?)��{L���B����S\'�L�m'+wy$Ʉث�AU�eh0Cq9�ܝt�'ER�e� �v�}Ӄ	@�����L��:���m2�7ˇһ���b���?��Tt-jm3������*3A������s�CX��	[��3B�(&U����ZF�� /�#�W�<0N����B�ҜE�����чr������%[����q(�`�x+h_?�]�=̓7S������\��s���W�AJ
�~=ʩ��N�u����.lh�>�� )�kz�������a���[Ù�cࠒ���TGL�������?��OzY7W�⿤�TC��D��<7},&�57l��k>
������+��P ��l�fX�!��C�
VAV�]]����c%d��t��K���jN������K�C�	�e�z�x��NF��]V۠Z�\�ԗ��&�x�TY�3��5�����B����c/�l���� ~� aqA-�m�A�#3��d C����YMg���?���sl�E��:iu[�^v'�O��X�Es�Rt��ą�a����ɧ�s��D�� :l�V��լ޾%]7F�l���?��_:g(�Qإ�B>m�~g���8�Wn�6�2��E��"����>��DG�,�μ#���F*Ov�W��D�:�7�!ܭX*"�ge���e�L�'�mlʒǕ����KO�$���Հ癹�.�.��C��U����P܍2m�����F�o|��
�[��@��Twp�5�O��mЛ��W����M�H>� ���LE�/�g� �YC<N�y���]ߣۖa���˨�*J��܄�s��J����(�f ���K:f�v�P�%��Z+����["=;E�QU�y~���%�u�87�.�t�uU�!�ت0VQ�j�g�U�c�����u�G?�q�3�#�����kl�-�F/�_o�v3Ųdh4C�.��g�����&��H��U���*?�-�����|y�K��^�c��l�aL��b�?�pv�Φp���,:�^��ɧ9���s�����0�!�7K8ap�L�g�WD�u�(p�Ԍ���>Il���e��䴲)L=�Tf���9��5���q3�u!X���T��q�lA�W�������G�X!�W����ӱ8ƅe�ӻ���r�h�#�U���`��{e'L�p�6M������ӊ*�q�2�W��ZSX�̵s���^p�pF�a�.�w����5I�.�2�~�K�
��j�&�nܛ���M7�b�x�7x��|�
"�����g> ��ι:���D�U�_��ģ��;�����ѥ����>��f�tQA�)�j$�x�D��)U�M�8����|&����Ћ���rA�/{�/L2��}}Sˊ嶥ĭ����O�ɈT�w���i�.�O��Y�����𦃃1��#��z@ֲv�%�^ �[:���'�H�m&��,642�	 �ȁ�RMv�~\g�l�3�4C��`��xi� �ɚ�����;�9�R�5YOO��}9��k�0��A�\[Т����Y���9gb8�Q�K03�y��hiI)wi
��B�/_ iy�Є,��.izmY����@�x�9�*�$y���lH�wasi�'���)�����2��&����L���iv#EK슾zW�ಏ��ȽnwC#���Y�>���Y7 ��uظ(��
�����c�6PW������:�MA_aq��pܛi�j���������kM���W�[�M�m���(�W�Ba��a�;�H�0R{i��jn�ĠQ�a ��H�+�ڮ[Lanh?�b�%�����p��M�y �$]p|�0d�l5�����h�%*��+�'��[?�1�#�a��!N���zg)N����3ϲ��F�}lY��_iBs�v�7	�Vk*W�\U�Pwl�ת���}�F�� e�4���y�I���¢c�&nz�Uz����E����)>����y����*����[�9��:�A{#��������5�!Q��:�$��_
7����XML!�1���^�F.�����X~�.;�ti4NЀ��F
��H{&��e��f��p��f�u��cK�����Z.��ѫC:��2�fhi$��:��I�9@\����ORSog��\͘�ԓ���Tv䖑�/�/15�QaԴ���C2�D�+JD[�fgZ���c������I_��w��R��:�O��Oݕ��W��~�STu��	�Q��a�5dQn���kb~$�z�]%��x��A�ɖ؏2A@�Ŋ�Q}R:A��U�'m���R:K�����ٍcCu������BDٚ�6̬2���^7T���]���M�]:�>�0efT94H֔ԏ�����GPo��[9���1�|�F���Hn۫��̝6ж�m��-�~<]1�
#V�Z��|#��jؐO��d|�xB��ay�)�W%��4g�|��_�S�Y�o�(=�"��ֺw��|ᵫ�5�L �,���p�w*$��̈�3��=T�  �
���N�k$��-g�k#ބ�9��ʻ -p;MZ�R���bH�[gb�D�����N�*���"?4��k���3���Y��Ga�Ru}=��BG�9�̕/~h!��Mf�o��%Z�KN�QZ�u�gX�:�C֊
�֕��EU6�Q '�T�{s�3V�T;�*�ڑ����n\�m�����h��I��|��>~Σ�}%t*��u=�Cl�E=�\���Q^��2w������BҔ��D�k�+�R�U�fLKW��Ki��������T�J�<*t���Rb��V:��#�S+ո����jlumWN�; '�b��75C0իB�r�� (����&�>՝h��|���H�[D�u������l�9`�*7���h};�V%��X�\�L�����eZp�a79�G�"�gS�L~2��vV���8�)������ݖ�D���"������Ø��Uj��u"T�#WVj���g�$ko���ѽ�z�P(?e��(�j�b�T&Zڐu.��4���/�5҈J�j&K"
TU"U�)��b_�����a|+�۶�.��b�d�����)�r���GSP/������t��MS�aD2 k(�1C!~�7#��d�"�>_p�S��7|ͭ�1g@ �\d-�c@f��]3a� /�P�ϸ����۱5��h�� _�>{�+�au�h#i����a�7�#�#�� )(��<Of����@��%��%KQ�j�-ڸ��Me��<����LJ�7��a}�J��`Wx�����~�`8�g�R%pn����oy;	 [GB��M���U���v-pyF�4��Y�R�s�e+(�-�aȽ��)�W� ����^ã����OK�&���� &~.{�hYG)T����t��L(�引Ș��ڨ���a?��c���	Qɯ5��ϕx`��9���%�e�u2��_$�A�������S@KB��2[1�B�&{�rCX�n��5���!��q����y���VC_4ᐆ�a&7EJ�s�'�։�6��|�}^12��%8�n<�]�yb��pv.�g��	�΁Ѱw�e�Ǩ��B��w��cv�Q����&�4�Ǜ�����d{㯀T��M朖�B�6B���4m����)Nܟl���_tg�5�H�5��?W4i.0TԜ؉�ݧ#�ڷV���,�~)Q%]��L+^�RN���?98��A��e�(�t3Y��ؒ�_N��9�<%���o�m��к�N��K�h�П.D_ڷ��u1!�S��^��T���z�{_�-9�8[��:�\?��y϶�N�1�ĕ�SC��*��y#!��S��MS��@y��7�@:v��s�j���+��N)<lSp� �V�<��aɎ[������A�f�$ F&Bc�����J�W���2�I�N"~�28S"��B��}'���mȪ��*�hiQ���DKO���]��M�B�Ï�a��g'Q=~Vh("BŦV1����X7��,$�iݽqa5�R�t.?�
s�w�7�E�����G�o�Y����
�0��i�*��=��n�
-x(���d����yf
�L��[x�����yw\�#�/�zz4��߃��S��?Ey��@� s�A�Amw�(��97����q�\}�UӖC[~�P9�뭍2�Xc.,���r��-i��)Գ�ԅ��W���r4C�P���)BO�uJ���?���Q�	ZH��N�Ar�>,ʤa�|�6IzC��ķ���FW�"�I���ע:PW���E��`(;�d���ӵ�4�J�h���X]�KY#zl��'δ��u�CP�Zu׋�0g��(Ɇ通D�}2��6��2h�L���T1��#��ml�(�d�qK�,��� ר%��0��*p�8J�˼�~��Єc��ϳJ��Ư�+u�~�]5�y�łR�~M��0Lcd����} +F�@�zFE��(�r�OpA8D�k�QQH�'��[1�i��h�@��n��ãb��;���P�=Iy�s�����h�KשB�~���H��Hzٜ���\�K�sj�K_�Ag�USzwӛ�Ģk��⵪��{7^�K�x���h��Ok���㕙����9v���G����nH�S�-�D���X���Gv�zC�� �;{���6����)y��l�����w��DN��<��7�|�~e{ ��mٯ]��YP{��ݝH��6+���1�����`�atHV�@ֹx!�Ʀ]�n͠0����Z�� �t�K�]�����0EҜ±���@f��7D;
4+ՁX�)��Q��l�h��?�Մ'��:.[X�&<�������_j��tdg���q�8�:��.j1$�=�jMuZ��(��Ӌ��T�yV$"�X�H�F�I�/ %�Z�n��9т-D��X��ɱ:R�Џ�t����tK�D�!מ��_�mքv���h��Z��8��-xc\�r�]S����^6� �Y����?��h��r ��N���:��7�㾍�1�镼���x��[��g����$�~�Ę��	p3�س�t�&�pR����oʜ�r��v�1�WQ�^�zBF?c z��yJ�r��V�#��őU�S1C��$5=h=�����^�̗=E{Hp
fa�Z�:_����'�g���R�dt���ՋH"4I!�M��GU ���k0߲7���k���� sE�ױ��b�<��w�,5��^Y����[��*���O/�3Z�	��L�jD�N�,�O��~fD���}�2Pv���v.����ܯ@���)�oI�D��C�ߵw���w�Tu�蒼O�.��h��<#0�4qs��o@HI�`C��T�����e������n�ǵ���m(�7Ռ�J{(k[��.�{rȖ@�]ކ8|��|��N�|��a��{�!Y`0/����sr�����7����F%P8(��8����%��Ź=�F-�pmG��2�Vf�;��1��g�-��$�2��sc����ɇ]YP�ת�N�*#�)�����5E�)]�zi����`��((��ѵ�pe�h<���g�k9�q���S��X����	s�$�Jڙ	,b;�
��B	�&�}�&�r�\���$G�2��,�1��~x�}��kjڶ��H�jil��#��^�鯷������C/o#�kR!3���0'��)��.3��:g��^f�/,�NVm�js����`b9�L��P���-�)�>'��_���þe-�_�[���3�p�k��]]�n2,ڸC��zp��M��AP�R�bZ�;v�[hw�'��HPIaA'�	��!���K(fS�3|���g��ʇ��E��9u�&�3$�`�Ȱ-u}����㰲�����p��æ�6i���o:���S����/����m
���r���3��t0
��g�����/�:B=�M` �3֜>�+6z���,�_eXOQ���v�9p���(x�*&����ƣQ/�Y�tcƚB�KI��_Ǹ����;ޙ�(Ԍ�&�q�]�%���R�yk,�*�6j}��y�Ǖ������%	;ڰ����ʷ�u�8�a.�
�}Դ\	u�P����G�d���8
u^�|�Gr�YF��a��]%�d�S���\B����k`&E�`F���X翭�Jag�l�[�#?��.x%)L�ˍq�G�O[咕�i�)���@�I ���o�Hm�aZ��^g6^����"G���!S\1������C��o������ķ~lp�to9�/\$Z���:�������3xA��'�*�*�U�UBTċ�G9#[s\����Y3�
o��Q���c�1{�A��X��*u.9�0����3_��%��F���옗�\�|j�y�y��=�D�JX��5���|�����ސ�!mF�N��V� Q�`e�7���������'>�{x�nvݭ�n�K5�TOw���H�g������SP��'��A1����f�..��
`H��dA����}4H��� ���'6�����-�Ҕ�9�Đ�o�+��D]2��*l#�]g!V��KSZd��!n���p�E��0?d��������u׃�~&��Ѡ`�S�e�	���	���+����|����G�pE�kW2wq��PF�E gѲ+Y6�K!��&��?���Y�)uW˚-���T�n`D�����f�D�1��u���;\Y��@���a�4��"���8�����o�`1"��WZ����JՅl�k�Ҧ��3�{K�~���0�~Xr�='��h��7a@��?I
2�	S�I���0���cEg�j]�V����Qg�Ԁ�d�ˤ6��Vւ��,�]u5a|izH��c2����cǳ��~�B�F��C�6�M�D6��H�;�G�uLwy��ŗ{�)+��CӖ��5�~�Wh/L�%��GFN<
������B���?�74��L�Rԉ}<�O��j�&�]��`\i����~\�¿�"�Yw?����Đ!Kʰj��8f����C7�����g�=
�*}J(;0r&�� ,�M1�R�E����*윢_���E�\,�$��J�R�Y}�LF����^J��$��ͳw�����r��+2S�68`{(��Pg9CmW4EកI�;���L� �K�2k/~k�q�E[Z�(�5���Zqc[,|-8��`�]�fq
����8���FӢvRg} H�g��|V#@�����kX�M�B���kN6Jh���&�!9��I�\�׋`i�Q-b�PD��s���"x�z����.��g/p���R�5�����"�	��$cYid��:͍�#Q7U�c+4]�f_mFcr�r�!�f�ٛC���E�sd�U�Wb�^���
:aE���!���W;T�"so���,Y��]N.�g>y���3�x<�����aM�D���Nʼ������1;�P�J�Z"^D�F��"�j�+�����2��"J�>�L�g��X*��K�����;�W��8�5��F�{���	����]�	}��s�C-�GH	[@��d~}����-S�\Ԕ�դ�D����8�:��L���m�Q0�A.��.��=ך �$��8X�3�S5��I/����X,S;�>�ft�����W����s�Ʊ^}R��:onN�ا��:b��-r�m2����}�8��yc>�bAk)
�G���#��p��v1�	�3A^'�����w<T��|��&P�Xz��`��6���*�����oGD綏��1r�8��f�G��V�fu^&��Q?�����`�����]�j�����vvk��� g�q�rY�u�$e/������wd]@�K!^<�U#���QM7p�w����pw���Ym��"�/ػ���K@����w���iI���|�ā��Y��͔��Xb.O��Y��hG�1��t|��8�[�~��6/����=�,�f�-o8�����2Z��.־v���˶��85�#�N���/�Q�-F�s��"��Μ�j�,q ��v1u�ש������:i) -G��V����A�a�|9 BX)/��M����c�Y3��D�U��1��������YN�K4��9 ���jĕ��Au���lK�IM�����ڪΑ��;����A�}�{���-��:			�@T{�F#��:��G~����hà5_���A��	\\�#6�Μz|j- ��߀K��6��^9é�7�,�u8Hcw?9�1�M������QOɏKs[V4Fٓ1z�qI���s��	KBRرJ���-�)ܝЮ��P���9f��A��M%�'!2����b���ݵ@���7�iR\��z�,ѣ���p>���`�!��^�ehǇ��)�[7�d㘇رE�{g9+R��ƷB!��lх*��[�~�ĝ�e���F��$�hܲ�%��ûs���p�p�r���ys��6��~��K�-9�a��P�<[��=�2�-��}�hki�חJ?�l�y+^u�����R������	([� �~��tQ>i~�a��%9�w��A��O�|a�S����n@�1�bz(c2�KH���q{�We�H�=�X%�Ԥ�����.̽L����:?(a��7�|>%\>I�'��r I���}������m���G��?���O����b����2�.ESbk:�m��Qj�#�H��Nb�y��(��+�5sϳ&S��(����l�c�hp�GB>��@d��Cz��6��NJE4;��h���b~+��t\��a��;�
�uJ"��y{Fz��L�Y����ɆBg#�#��PQ�G-�q��6:k��*��c�]*
��=���M���Gc]3:�1~����O׳mRP2�p��3�����2vP.pڈ�ҧ̐�� �KT��3��ݎ���8�A���<��w�1�h��[�˖K�^�Yhd�860˙�+�ީ�Z1�@���^!�]��C!D`5��\��|N�aUe��C�M��F �YQPBt�
a%��P#��ԗ4B�E4iL��8��n�.Y���TH����J�+v����ze:��k\����M\Dg�F��y$�tEӏ(A͠�% �w��� Xq�t��A��|s>L�|jj��=��p�Z,�wz �*w?��D�bը�&�k�V#�'D��S/���k�V���Ǳ0M��������`�F8#��(#��>����	��T�ev��t1�g]���.fN����:��f;e�:Jk�o�ʓ��{�)z�Mj;"�/lC� t+��8�l~km;�v"3���B��f�q���a*w�0�����4�+��8Q�仒kQ�:�
/�C��eH�k�yP1�Ǝ��V��TY�^fγ��-d�H�%FL��!��o׶ ?�Om��ղ���Л�γ�e�d6)�a�c���M@;[�٣���9T�)�u��em�ݗ���lK�w!)l1��[;d��g<\?w�����C3��U|��h� ���V�	kx�!˫c���
��\�ai���µ��i��$g"�$��u�9��.��D�&�.)rx�?R
��ܽ���E���aq�:���@�kn��樔�)�2|���48To<
8�}x� p�E��b�A&g ��l$�Nn�+�8��*�������k )b�(#�Uk��RM�vX�Z�|����r�w��rM�&3D�Y��B2�[�+[ �+vET,���2��X�	i�~����1ѿ���g��'&G��o����,����]����* �V QS��y��z<��)@U�+7����p̬�(��:�"<R�V�Z��:�Y�Oe�B��8*�7�6���|vn��ǔ3�Ƭ��`H뼖�L��kBYR5/�`l��p�ޒM����6�kp��-/
$��zE��5>�9;hb��n2�z?>ΧtǊ�`/'i� :,S"m�^�'��+h��yb�>�H>bl�s&+~��ک�M�s{gdx��G��Yn�0z��'��H#�q����h�)��*�e"����+�h�ώ��|�{[|�n *�B���]�jI���P�S�)V�y�*��W�k�R�P)�" ��x;=�SGZI��_R����k'�i�`�RYL!&6,�e��lȵYo�D��5�\���F%f��`���&��ԬTO��F
�WŨ��U$n�q�% ���x$38��s��QDę�hZ|t��T�׻s���G��"NC7�N;��L��$�V�N�y���	|�$��o�)���%�-��|	ݭobe���Q�'WԠ4�N)�/f�v�a%"5|?�l��%��||�.�O�%��!Bw�����lNs��7��mu�����d`������%�