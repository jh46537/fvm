��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0�����(�_?V~��
�r�-�ǥ�bߣ��\Hj�1 u��>j�f��o唌�����b(@4b�P���/t�Ħ�<�#�gQ�b	�o�;.�'_��`�@eA�QT�<�F�_�P'�?��ug&`3z�:Jz��"��l��ʡ5e�7�؄Mg�_��h�����'��<��n/�'���˝bm's�9Kz���������,���/FK�=���߆}���6���鷼��(*�õ�[o�
��M�܃QMߚ$��9�t�B�z�q9�xl_9BG,@���ϭMŬ�CݞVq{�m�9�E��1�s&��s�:2���~�Z�pD9��z\C���N`��?D�1ٰEB�4��ϔ!��픣��#�9b}��"d�)򜶞����2]]ISꃅ47|EM�N�6�R�em���ی��GS#YŞ犇d_�����d�Q*�a���z���1���f���o�D7^>@$�V�� ��U�
��O���RD��g�U��N�UY�w%����K.�C�t�ވ�J;S!M؁�A�{���������>��Vo�q�c�"� W���?���� ��ŬZ^�ri2��Ⱥ�i�a��{��RJ����+,�+-d:A������T���C4ѧ)������'�Џ�uh�䬭��'D���.��?����r)��V斕�߁4y�� @�����C�8o\�K@��PY.���D���{=�7���4�м�d[9@����)\�x����s"h��Z��2e�F�u��#���$7T�\��02y~١����W�]�3[y��Z(SH��Oc�n7>�9� `$�`��9o�b��R�q/zzΆ��R!q|aeq�h,Ffh�0 �8��W�I'7M��#}�\cġ;iw���0UЯ�4,��J�=x�_��~d0�@[���t^{�����u�Q����qG�J�r�k���Y�����)`Rn�O&��8�f8C�g��K�Q���)���Bƛ���3�ֿ�;�>]e%��).1w����� �7u��!
�����o�S,�K�F�c�K��tˋ�n�6�"44�R�)�R'�����pm��#��H���Zh:�����u"_�p���k������dM7�G�-�¹�[�:]-5F	����(�����U�#��'r�*H:��_7B����#��
t;��Fg�Bk�ilU�2Bp0�	5~ݥ�l��g@���5e�_��&�-P�ګ�$����kS/�'V4�b�\�\��8����f��Q~3f�:�+V��B��H[�~����w5klp����,;�̙P��g��� �]��8��_�N@�f`?�L�U��ʩ��qB<2�����8Ϯ1(H*@G���RB����1}Nl��۫�6���+�×/ٶT�rr�!Pn���Z�ĸv#B����S��f�4{�Ӽ�Tlt��Z��̬s���E<1����"g?Y��i�fm��es�P	����Ûs9�
P����G^؈,I��<�֮W��{ ������q�嘙�+�M��GA��-v@t�5'��`$ޛ�3'��u��*Oci 
�H'?F�ʼ��N�-��������!nA�����_��H��C�oLn*�ޯ�|��HBw���)έ�w�d��s�b�!�$sQ�=��l��AP4c�I�Go^�ky�P�$���4�Fn��ڠ�kPM�FÇ�9���r��G	j�4O�!?皱7ӷx���U�����Ώ6�_,hі�o!�g4o��w ɸ�R.7���9π,{��VMЀ�.%㔪SfW�?N�:T���r��C��r�[9���F��/T��-��t���cHS���;���J�!P���Ӛ����chq�'��%��'o�I��|�FF�E.Y��Rth$#���g5�O�*Tx. .&c��jꮧ�͜d��Hڴ�X�/���wdDP/]N��>�j6fs�	l7.���s�'1�p8#9�Ҥl�}�滗�`c�١A���2�X�<�1]�u #�/a�/��N��(U�Ik���Փ�m��4��+��2��9�=�|˵�qAɭ�/d��E?s +�K)F�}i���^J��A�@9MkM��Kj��{UH��m��JbCBh-����d2�5�R#']���Q�?:zWJ�Aā��V'f����n8���֡H������?3����C��C��J��~6�=K"!%h"�SV���]6���\��ה��O�<��罫�Y��Հ)�PI�V�>�v�Hs����V���D�l@�=�p���C�M�x2�{���.��������0�����xw�.ԧ?R����2�=ĔD}±:Gޗ'1Y�G�;O�U�����Ȟ�̀;{
� �~��JZ�x�"N'���b,/�mǵC������k����]Y'��V8O�C 	0��LeA��=�M�[R
��l{ut�qdJ�S6h	������E�c��I�>�?O��	�J�͇dC(h.��h���Oo"[	a�T��=x�@�g����6t-���[79�*#�E�K��~�b2���	{�@k�"��/����������x�ͭ}�K� �{���E���_�!a�oL�s�Lm���~��S��-vW��w���"
�:�r �:�>�1�����\a�ϔȬ�d��=H~�v�X��a���v�9@Ʈ8��.D��e�,�76�$�.S�����y�ј��K��p�i��i�B��|�_��?K%H0��Zݜh��	La���>�Y)��^Laai��*�G���W�5��ηY���T7��ﭩ�ӏ�BPH#o�ы��=}����Hj���c�bg��fߤMߴ#γ~
3�|#o�U��=��EcpW���E��$�F>���X���vD<ԃ��Y�d�l��O�*7�ʮ��*���Ģf��^j	�	A��2�ǥO!�O���n���I�`Зcz�!Sڥ�x�UD��zo	�YS�=�!;��������{���X(,�{���x6�-��F�3vu&�n>7ax���W}Z�OR�u4<��w��{�C��;&AD�]��^��8�X�э%-*m����D��ݘ���E'0|d���$�;�:cW2�M���H�o�f5a���z��5i	XJ(`�ڑ�]��_�.t`��5��'��1�
M��P�`��n5/24Z��s�h~�%rʫ.x���JL��}ö)˘�Oke��1��||�P'm�ZSOT/��`��&�q��F-ƲkMӸH���H�{I}�J�zy���!s_�B���:�g��or�4S,vp/o�P��)�P-sk�b�ݸh{
�UW,VZ��N��E