��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��ߨ�=�]	7�N�)3�M�Ρ� ��B
�i�k<֐�1(�/h�"�+r��ҏ�X�fИ`��6.[���L����Sg�$|����x���
����v�95|b�fUw��e#���`r�|�QZ3E�*��e$㩥�֢H.���a9��[��}h��P����{7DI�y*��f`�K�>BW�{�����z��<�	&u2��<��q-F�zB��0�t�c\��L��U�Z���T�u�o|^��G�)�=�d�so,�yr���o�L1/�%�o ��)X�A��f�H9=<~�/�f�ԑb��ޝ��X����3�5�_�O��AX��ˡr*`�}�1	��83pPR]�B~ƫ�ug�D����2�9� �����/E=4�pzD�<QCY^��}h[
KV �����{��g$_�_@�6��F��7c��m^�<E��.r����@���E�X����K�)���ʶl��q����^���3&:j���C�/����\����\��f��y
0m�K!�oHg�h���{�/�l-��s�.�{w�)�����`��-�O�p5.�v���74��c�h��P̿з$�����K4��{��&Ӷ��*z�Е��S=a��IDJ�����:Ļ��)b��ݘ1k�u.s�p��DZ�t���t�X�r#":'�7��i���^��%G�N���+�!�ꬕt�7+��F�6���5�nUTw����͆�Vo��145�����Z	h�S���O�\P9cE���9mz�=[h����O�e��p�k��t��_�7b����T�vij�0{!��	.�YM[_��*
����ǽӋ��G�hv3A��L+i�)iF�;�i��Q���ό�Y躰��"^�2��B�d<��8��i�����D�^��Qa�]�x�rl��X&m�Ђ����k�>h�^��(o}*�Ո��6{l>2�.`N7��<3~|�����c��僞(�ʌ�"�)�r��]�OB�_��2gm�>���(*�i[��Ϲ�ݾ�]�u���*��J�W��skƟ}���`<M?Q�I�u���]	�G&xa�=4�⡴v�,dR�$6��<�b��C1��nb�����G�2�T��Cs=�W$-�e�J��b[C�Sv�.�n��8��_�Uˮ�&e]�$>J��\�3�͒:�p��h$�<�5:2�:���e�Ȣ�S$4g�[��(_{�_}����H#�Go��|c6h3�,�s7vV.�yѵ9wQ3PL�ZM��ݬ�O�L=�\G��#S�� �J�&�F��Ի&u�+�Y���r���$y�X u}�i��Ű�����t��ȸ�%�j���G?�$f�����6ƦZ �c�@H�����N�
)�9_�:�\p��=��o�v>%��w�984�r֓���
0��.������gbͷ���Oˤ :G��k���D^���U��[��Pt�[��Xa#W���R���3�+�?L���4�Z�����j�/8�=`��XKj�~ �Q}~
��gZ����AX�w0�*��;r�EڲE&J�y�P(f�����;�ա�������c&�{��AFc�������k� t�߶@d�M���/F���������#��D.��&]���a�Pݖ�OK6�Zl7�����0� �q)�3�ȣ�-�Jܬ'ęaňJ������Yq$1n$���=zZ/w�iSx�O�6��kďޅ���?Z�8'�x"��0�C��Y%NOӌq ��8j��E�h���mh��S� 6�u�S,;Z�|��$dn��}���m��h4�����$�S����h��؉M�gl��2C~h�2v^)�~����L�r3�lS����pҴ,=fD��?>[F���c��v�VK�HO�G�@��_�t�3w6َ��wV�) -_���!�W� �~��h��+�OA�NǵHh�>�:w�k�n3����R�
\n�e���!���"�7rF��$����km��1LOm^:�Xm�H^w&v 5Ms�ȿ��V�K�F�;��2�d=̂vÃ儴��� ����M5���ט�O=x������8�C��%�w9� ��[G�I�w޵�Q�u��_ׇ�}Q����B��f�� �����B�d��,�9[���	��A��"��qlKt�� ɰ��o��k5Bٰ�c�#�#����O�QKhs���0�ʄ1[{�&x@� �7��b�?�a^�J����צ�d���^�@���W��i�lz��[� 1y��F#h_�1����y(t�踻W?~|�F�G5T/I�m��x:<Y���<���@���]��� %#W�B�6��3�h�a<�ʲ�ŧe��'Q�^�u��k��\bq�@�o��WF&!!�2Ǩ���V�< .�6��{���J6n�t{Q���Ӽ�%����jI����i�}�Kʇ*��)u����<�=
vC�4�	�H%Uڢ(�1���:�(S�f��ʫ&��i�O~�f��S&)B:��F^�֢���^M_����f
����t�l� ۓ�+
Sw�B��Ş_�J���/�H
8�N!��"�y�f�>�Yٰ	����{�['��J����5��.���%�lw�IM3ݠk#O��E�){X#"����s7�~Y�·������k�Ę�쁈�jVy���@��T�i�"r���@����`K.��gQ���3��0���G�8T{b���2a�P��\�)+���D�=$�+S�׮Jñ?ϕ\!D�t������?���І����fW�8��/�ͥM-���9n�'�B7��p�=P�/���ɡ�8�!߁����`P���Eѕ�1ɐz,T�9j�����:�Ɏ�z?Q����:h�l���f|Z�3NpZ��h{vJs�b�I�k[�_��\/�9�#Hϝ0Ab�&��/�pV�O>Xx�����A|$����N�&���9�V�lt��k9�� qi�Y<OBW����@�Sg�7�2�Z{#�	0���:�դ�ɝ*�]ܵ/�U���l�<�-�V�Z3X�J�x�{���Ph2�,L���.R"��3���-����c�Tv�i?`I����&8a	)��l�[i��`ߗ��c��AI�$ޝ�wD\�Z���ygG{�ܡ&1�α?kI�5�n������:<�YQ>{�-����wd4&��<g���&�An��đ,%%��.#���f|b��0�N�L�p�T�a��@ӂ������,D�e��ZMH�u��׿�������`����PH�"Z�yRʲ8�}����Eyʗ��d�ߙ��&=�$7�GvLF4�t{�|��	0�@Rw:�zO坩�8%�����?�0\���!��(��(#r1> �Yk�0�?��"��)˶ϯ7絠��h��-;���ĥ�;���s��"���j؇5��}����)SZ�����(bM�s0��'�q��0к?���LQ<���ꔪ^�\�gR��S=�h2��~.�祳�EZ��$p���L�M��j��r�ӻ, ��}���}
���n�����(�(QR)d3A.��ńˡ
O�>��*p�|ޢA����Z�o�1s��%]��ky��^�I_���N�Kk������PK�YZĩ@����"(# hDg`�]�G��#)1�����\\�G�!`�f