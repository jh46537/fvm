��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c\�esR&{������o�T�e�Z�/��`%�����1�2��g\D"[ޏ�F�
܌�)�u�lg�h���T�Rfc��h��H��H�q���,�+��f؞F�La���q���Y�ޓ�J*u/(H�u��^�򧵖=�L�A%���o�a��o����?|t(Y����:$�31��Ax��cR�t��cXun�	�<��{j�L`_�m!\��X�/�����~�u�`\����?y�?��T���h2Bf���F�=/	p��^�󙁚�H��'��b*�f��_����?K�D16,����1t�&���kĔ�u�#� hY�^e�Rl�np/|��k(U��-��Y{�d�˧v|G�/ڏ�{ZHQ�T�go�T=);�Z��ϙ;�h6��������e�#w�j?��5kp�J����h�?�YD���.�?ڝ�� �E���ؽ���\ dWw{�e��?�vM�Of�{L��i?�`��m�= H�Q�S	�� ��Ե�Xl4���
C������лq��`�P�=�fH��N��w��7$7�gPS@�N[��~� J�t�Sd���)	r�`���-)���>y�@޿�oէ	��"�	ˍ�m�T��u�=ѮSٔ0�?If7�8AS��=!΍y�h��c��h��ER��10<�:{w#��圮�H��tx��H�J�9�$�z����ǎ����@Rp�#�5��a
��V�IN���c�)%�~՞=p��6�������E~IG��8�P��Z�a�x�e��&,n-*��>.r���?�A��*���P@���Q��Hw��coeY�XMii-�7r�[2������	��g��y�ɢt��nхR��;��������L'O^e�����p�D����[��[���_��	�<����M^庅xڧ?�q{o^,:�j/_���8��
,�֎�DN
T�!\��!�80��B4-ܯ�	^�9p���u���cU$��K�����<,���3�A^3C9J��\O�M��Ӂ�}+����-�&2�K�}�]f6��[�=r��٭����-��Jjl��'�Y0P��q%�ˎ�{A�\����d����=���-��T�)�C�#'�6T��E����kDr3.�����}���+f�fйA5��O��my�bU�Vf�N����K(H�����6 ;:�5@n���~Ӭ��n�-�ṃ�*�ט��F?k���'��e,F��\�R��G�����v�[EYd��PG��Q(�&�⼖f7�v�T%�O��r)B*��/w��Sati�$хn��H�qf�}t���h�=T��zc�7<�%�����9�(Ƥ��H�'Rdm�Z�zp(ԝ�h����m�����gu
�k��8Hi��n��H`�L9H�̧:F�h7�4W�ؑ�b��^�&�;�dTm(�/M{����N����ޯ���[��A`qʚ(�2��c:���{�{��q��4�	W�i��)RZ}�����2�,��=���h�[�?�Ɏ3{�#S��m�+�U�pt*j*
O�M[(�O�W��ϛx�;֯��$?�~ynP4����q&�i�C��ye|��$jf�N<6W�l�q����(������ihJ��UH������I�d��ؑ�n�m}-�M���H1�v��3�c�����,�1(�޻U�޸oL�N�L#y���c������9K1<�ey��jL��&�(��<n�u�h��@�W	����=X���](SV~x}����lwVXm� ߱L�05���:|�,�}Ӝ���l�\�]6�i�_BbU���r-D��	4��l�~��O�5���#@E�p���g�~!��u���@�����0Q6n������G�TB�'�Fӏ^����#�Ce�Ť���.�W�/A;�ZϮbo���&�Q� �zr�a/Ē���%�;0�XG�65%	�n�bE�J+z_���&����G������7�  Pg'�6ʅ)�C����H@j�a��"��w���T�eѵ�e�ˢOMm/�X���C'թ@�!eά�֦5���3�}��,��\M��(�_e��7�B��5ak����g���Hܟ���'IܛA�J���;��;�6N�27�/0
��/ۉ�ʆA�E?�R���K�,g%_k�ŷ�4�l�9�(�s3�3�d���}��u}dU��߀�;�x�#�led�.|i�6�N�w��8���
������i���w����.2�!�?��U�sf�D��m���1�E�~iE��0�� j���i)3�]��i	��Il�\�I�h������Gy����<$��g9<��#�����Uesy�?�f�1��ԈtFr��+�C���k�"=.��c�������U��������.�Sd��>�o5UT���c\G��'�_�䲑���4),J2_��썁��e�K��߸���<��?-d|z�b����7�y���XU���V>���'b:�MD�G�ݗ��!��0�dрJчȚ�w*/~�,���)´�A>Բ���t�9IH�V��l��\�)����@?�	<MX���F�|0�ZטѺ:���H�p+�����a��T�懻���i�ǌx��!���cCB�ޝ~!q}M�4܉�kޢ�FN^ ���"9�u�MD��F�+;�.�����S]\�yv�J�=+=[����$�$E�Y�l�6gbԅ�����Z�7�2���vF%�.�!�h���v>���=��Ƀ�~wf	��v�8lo'`X"`my5,"ۆ<-�֥���[���M^�@)��V�B<��2U�/�L���qh1Ya�s("��me��*�㠊"4��f����Q�����>~�B�7���u>�����LW3@�ldT�b_��q��,�N����>�%m��)�<8RC&�N+�~?��}o�FA7X��R�l4��=;��&d�D>�B��,��ƙ���wS�m5a-���wu��U����o3�g�!Iϊ��`��fƣ>��gc>�0F�o���	%�7�'�U	:o�ִ�w9')��Q��J �+�� �g9C��t��N$��-穽c!4���5] �V1:]6l� ���P!���[q�t{��%\W�m�h�%�e��T	h��{+�����w"��d��$�n=�%�Ư0�fyۋ��cO殮n����WH�{&�fc�8G��ZJ�P��Gd���f�U�uլ���)�C|ɽ{��@��t��7Q�"B 
�-�ۣ�vm��pů��� �����I�-���1�p�6��$�P��%��z%��&3��-0�N�z�ow�$-���N�E����=����]##�>Y��ء��kT�o?��PZv��ێ��ꨁ��N��MzL;�$X-�dF^t鹧2������'��܄=L�
�9F7�F�ϗ7��u��@ �J�a=o��1|�wx�&�B%���lqt;G��
J,�X��D{+�2v}�5��9�M=I�6W�]ҫA���� S�3�T�{�p��.�W6D 	U k��.��8A����R�K��_�s]4ü����9x���y�zy��+�JBy^��l]�!�a]������N}�-�z�	~�ZY[�5>�')$�pq���"f��_��F
4:|H.�����n̖�Xͬ]擋ٸ�&
E���'1��2���{mt�?�A�q0_`�0a��]��i��TaC"	���so���%Bndiq��6p��*�0�F�(T
�-s�Ӊ�Rʬ�K�0�"��k�%������=*f>;��CSl�t�J�b�>���F��Ay���[Ïp����wue47!�>�Ҽˌ��u�ti���`����U��n�`3'Nk`�,�"���p���]]��P�)> �R�IЋ�OS�h���*�<�o^]n�-�<'$�6s�cS� |K9��&����E���&�>>B!-%)݅wV�hs
�3|F���]+�f6cѹ
<9�͌;(����>�^�_�˖.{u���?��mxv�5s��i���qc��0���3N>���Oï� 'y�҉�mA#ip�c�t�L�w5G�ͯu,�O��JuR	}3���I��k��A.]]���6>��|��v��R?���`�����ДGXz`c��HjQψ�����簟���7�=f��T�*'o4mI���P�x�(>v�Kh��09O+ڳaOX�a-	S�Jn�}��B��Y�
��r�>v��}ݚ5	�`iO�٥)`�;�������
�wF+�Ѽ|�%ݛϞF������_�a U�7T��չw��������y.2�Z�E�2����)B�CF��{��?3���ԏ�dϛ�	�v�3��@�[~1P�쐩^.l ��*!�TvAz�ogy�S���U$���xz<�)k~:����pn����vJ
?��b>��7 '�(�2��c��W�9�Z:r���[�NM��Z6I�3�%�'?-��XZj�QJdCFh��0 ޥ��p�sYhuqϡÈ�`�1��t�Y���x������ͮū�j	��֮����(}�}:D����������j�m
�R�m��J�P�Mm�w��e�Mպ�C\���R	9�͓��QW/lh)��Q�W��c���:��L�sT
�![�Q��݊���N__�����o�J*-��m.�t$��ۂ�
�~6E\�o�P2R4in�,i��"d�W��k��w*0�reC�=��C�ZW�ʖ��78mYf���|�ت�����.�m9d?�=�*��錽���*�ڮ��?�q��g�X���F������U=ޙ�:�<�|��@�G#S|�t8�N�w�կH����Y�������6��OD_%��O�;f�l��ak=&KiAޘ��0�4�k��_\�7��s�dw�J�b��l�i�9����Ų�K��(�7#LPo>�Q���y?z��p�d��g��O ���p6�J�{Q�l��F���W_�=�?c+�]�G~
�@iR�ؖ�Y����M�7V���M�1cet��#��(�[efW�7RpH~�Ku�#�[��x�Ū�g`-��NP"�ݜ�3�(�%΁I��?k����Mq�� 1�)	�����{�5?�4Ѐ��=��0��?�0��G��G^��j5W)�Օ��..�_�����C���N��|w�.�i��	xĉX�V�A)+h~��)�zu8�Y�7�T��!��"9�%�%�7{n;�j���Ql5H�EB�� ��"�--@eCĐ�����	��p,2�Sۖ��ȿL��jh�u�w�Ws��� X�[��B�������Kw�4���� �s�׫�{��D��O=TҳW�me��'�;��p�����t�T
f�aXa�H�A�J�H~Z���&W��:�WJH�6`�ԣ�$��"��y+�b�O�(��S>�*��r����N5���2�V}hr��"���F���W��ڧ����~`6�S4d(�(|i�UW}n9٪���4�k�{@ /*��ҧǶ��աG�M�z��e��bԆ&��i7���=g]C�?"��|0"���!�H��A���.~��߭< y��H��ù[jF�A�������e>��bY(���p���A����jZ���1�?�~�0	�"`��8C�eǦ�� 4K>�>֟���w1_��b�5�}I��7�Vw虜��@��N瞼�Hɧ.Gm)�C]��� �H�1�c���*�+�<�Ճm��yO���P������^��.Vx�("ad7���?/��v�'h�:��c̹_�N+M��NN���bА�!��Ue��1^G��v��L����\�!	"Q�-T~����.\��4����%p_b����p�����_�^h4�|�I�c( �]�%k.����Y�J�����y����"L�^ik��b�u1*�6��X��`ւ$l������a�u���);JW�QFn*�
�6�z�A�b)�3q�*T
hn�6*�S&E�0�M]��6�q^8������o��'W{�c�)0z��k8�h��m<�*wv+_�j�}���0�!>�ʪL���.����N�+���/�q�d����a��"y�а��%/]���y58Q�cAzŬ�u
�D�j�7<�n������*�O�X�=�a�ٕP!u���z/��O�z�R�$�Mn���֞û����ɥo+,��f����i>��vd6)����:	�?]/%�ԁ�s���D3��CK_X\�x�˿�ŹJ�硅,
lU_���T#��_�~"A�+<M�k�b��D䈍��jP^5l>zr9�R��Ae�n�r	�7�4�f	�ۿ��҆Y�2��Es]]��3:�� ��y$�s0����V|��V���^��+G5�>�r�3��$�(&j�<(5U�%�����UO5mJ��b�D���X5NE�u0���>�4�!1��P��iP��e�Fe���_	�}qh��Rt�Wu�}�LL�����G�{6��nT�������WL�
�[��Ԛ����a;�ju��ɗ���EB�0tUg�S5�~J�W# ��hv�Iг�V}�7�A���R�ďw�����q��G����p����"E�CCK�����[������(�N�ȶ��=Ԍ�$S�?��G)\o��2-�l�o�i���M#�b��E���Y�C�"T����ar�!�<�����c��4�V�uw}U��%�i��N�Iq�Т��;�����t�T]x>ERf�g��7��
`�nm�� �H�7]�O���}�.�ۜ��t��/"8�J�G�W+#"VE���� �����]����^^�P��ǟ�:;y�ݏ�t��l�d5�mZ�9�S�0. �cƈ���b�w�q	r��Bu�Lѻ��$k]JgU���F@BB'\dS�C� ���JR��Sii%I�}q2�\~$f�1&���I����p�t5�K�#i�=��)���/&��$o���yߦ ~������V[�+J��=�u�B�)���6;��%�_�t�|A!��l���V��qwU���xmғ`YN�ظOG_L=?^��u�w$}�u�(�Ch��6�y>�$�j,*#G�s�o��|�c~����sL_�_�b`�	4q��b�h��NA��^fpOǈ�$����������^�e1���8�;1L���L� ����V��yI;�ơ�[�f��q���"�����.%���>���s�5���㤞�nj�}H���Sǟ�`C�Ђ���OC��5����c�Ӎk(c�3\�=��u���rf����)�W4�䛌�&��y5���bǴ����R�̔\�D���M��t����4���ʆ�=�_WU��Y����*�
k�`��il1�k� �XJx������曋w���Q���`ٚ���-p�_i�nt:3a�ݷC�^����κj��t=�Ş��eP��M�1*��=������x��	�?*�u �+�`�@F�yEO�_��yUj����ä�"M9#��W��k�.�����>�<IF�������X,��R���S-v���^��m�=U֚s��R�ҩ�P j�d�Q��r�����B(!�
�Qd���jgE
N8��e�RM�����x�T�Ɯ����#1�`�5D��״v72�ݏܘ}���6�$A�,r�U8'������ʾ�W�ȠC���V8��K�T�ҽ�3F2��>�����j�����I�hj!H��V�D��g�""í��å@�ܫ��(�ד|[�N�M^���MS�mw��\�0�i��^7:��M+'M �ʏPˉw�(��]�U�dU�"b�u? �*o���U�&��bO���W𭸮��l �Ym�����O�Rۚ�I ~�����B9s2��$rw{A&:L���Q���R�l1ʞ0��gŦ��f��d>�b�۽�
�BvRc�އ5$�M�k������fyl��e~�H���/��Q��v`+���I�m����&(�T�Cw�!��\]Ň?���⍇�Ƌ�K�=��6��B�V�
CYeL�oW�u-G}۫bS]��n������Mƀ�mpH��rp]���5-0{�?�-rXaG
(�ا�\�A"r�z7��z������·���w�3�/!�?��n}2�g	%2Y������B���29C!�"��G��R��T��j'SJOސ�%"��;�b
�R���/S����asU{�������wթu�w�Uc�
���d�k;�W�t�z/�+C�u������N��Tce	���;(�*���3n���.���q�3��\מтyK���B�0>3��*-��sgeoc4^��^E6�>:DȊ�ȼ���?���ؘm��ۢ0g��i�ν�8�h.��{��x����)`���](��/�9�&�X��&]nQZ� !V���Ȫ�~�&D�hq�O$�Е�%˝�� �XS@m:���Z��}G����JB9�����YL���Q����N���e���`R�����f�*��v�1!M%GA��bҨ;j�¹]r��9��<��U�\y���GN2:0�L���������>�cҁ��#����D/H{!(�$�X�`��"3��'��7�ڞ��@2t��ۭ	��S�}�N�Qx�.w1�N�1,��#�������O�t��.��1�DK�28ߒ�1	Qj	���|m�m籱eB��1=~�{� �$����L]�
�$H�
Ց��u�S�s@���ߑy�,�9>8��'0v7������.zC�� �ɒ�ص�P@�1a��V��4�K�2�1V4��c�Æ��9�p ��3�+5kcUNn���2;������>T,��=�-܂r�D���0ς���JZ�?�h�+� Y�@�!Ó����J~����aM���"����s������+S�gJ�R�}h]�����c^*��2-�5����]h���b�08�7�`��QKE��7��[o����R'm5����`橭|�^�$���T�Խ�ϬM˦ �oK���o5�[m�4L�C���C��5\4�h[��o�kih>�� %�*O��r�=�TN�7��D*m�/�7��AYnFA&%�9_�->���b㸊3�K_ ���/����ha����O�o2VK����Y�]��9dc���[�=B���"�C��RvO�L &8q�d�K��~�%����(|W|o�?�#=?�5a�am��
�g�?�a��x_z,��t$��Zo��S8�J�2b� o]�nO��żj��H������r�5	�0fj%3�rK\���	�ܦ+�,�rf�0{��k�đ떕!o/����-i�]�
\�� P��۵[�$��$m��
�h�>���kl[g ��&�l�b�h���RLH�}W{��yU���ES���l�
��B,l7ʘ/��4
��,R��ya0}�>	�+P���T��lRh�8� �rTq��q�7�	����O��)�=#d�zK.�)��q�ݑ��m��Ǭv�)�7�����Ưc*+�wK���ŀW����4_��ıD:]g�́s祟��/.���,*-4M(���c_&
Ѻ	&8:�|�d��L6����RzS��N	�c���S��X����nM�� r7_�< ���_�8*]�4����.�*��Ud@��h�v\��&D:ާ	�1���{u�&/�(��Gx�ZZ����'R�%����ú�Oӽ�����p�A�n)���<��q��vm��0�X�??� ��,�|�-֭�ڑU-�k�p,�˹M�d�7(��F�$� 7.~R(�XI�"��v@Wy w$�ʭ��2�U���I��<�:`�,���-�;7�jd�k�-A���Kq.L�Y��7M6��{��+