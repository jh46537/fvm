// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EdZOsJR/M84nPlFpABi0kEFEDHIeXTZDKdSJqlkY13WDiGHeVz6abOEc26mne2Y8
dnGfJkC/kflnpGae6h5JXETT5rdJmuGbIQ6UUkm6Uzu4p+clLvsXyx+k+tz/Lp3z
F9WN7hj4GIn1zuv8rQMI5Z4WDMJtiRjcZjAGmgsS4iE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21664)
vTdaHVl99w/4nuHjvZXuItCKWPwf1KdfBfcSf1qJtYx6tpkikuF7osUB1buZ9Aed
vK3RLrGGajc8dGNMdGIrOEcyzL8hTwKSBE3W+CEgHmAQDXom9IPlb9qAo+kzhSGW
bINhvorhxJURmlB/F02EovnUqoyZPFOb9PNGt31ffB3S1vW1MYR9wx+krMxUi7QQ
Y95cg8qQb5X9OOjOQ58peDiV8BgcR8CV2+g5CpwiQ4bm99gAchgj++UrBY8okzd/
UTRsMTxt4xSI/Y1s/w7urG1N+3aCXEtgYh5qmGgkPxZ8Osnsw9n6XtWQa/9ZA7w5
N7UutyySqUuxMdkU/SNkcncDPtdXfBzq3A0XHt3Yx+k+wV8DeeWPBFRdQnRBYZeL
sbjDhM1cU80QG/9FHexdstIhIim0mj83zDrN8sExbsCuMjN+r343l7yjZ8yDvNAw
F98UqeI8h7peLkfWwp0dNI2+5aAnW6b4bo6HrqsKFY6nZB92dhkcP9sEdJexDQbp
eVMVqX9ixhD+oUzASdmqQIVSfTkMPS9vqpo+/N0xYynZWJ1n7YE1oVnmg6R0KUAI
+u5wvQfh0Z5FeLuH0qHTrSj4JaSBe4yTLSPGNMV5gVnkFeR1IYlP7q432xQ7uTig
C3JBZXnPoCIFfnZKmtj6UuKfjcR2akignh1WtzfFiYEEIijsAOPT7rmS6C+HKmxO
rZt7L/jPUhbT0xJX+0VaqGwkMQE/28TKMuLv5ocyc45mKnRZGhawL+LNaPxeuwUj
fbPWrqlQpdEm0pE2/tj1q6xPFzX+vLtvFmZSrXGovI7Thc3lY0rRM+DRH6S3+lfq
i+TXSpFK3yAMkx18REgsbzcoIMVUfLV1Ln3n1plwdJdosZnMwpd2YN4U9bM0B/pi
qK89zfpJXYGo6ciNm7/o11L0Uzhh4z8pfnkS1/NPgnuLSSGsmycIlfVV0iYMQyiT
3EMQz88twl+W4ao6K4uDewc2aPbDz0EBOJ8iVvb/G2ktzsBRyNgGkrvQ0WlqFail
pUuPuqpqMLMqQuXJHr7NOaaOi6HU13rjaCFsTc+DuL4XfUqE0L8BRx3jrMYzzX0Y
4c1ZvIxxY5qLfXlTzvwD5hxu18cXBIpf0L9TRW1tz0kfsxHvW7opf8U6yv8Hhbk7
iG0QHA0ZUgYh3FD3UcGYrsGVzVoEQTIr5MGNTue8gfpNiOsD8J2rzumszu0996VP
Xh3nLEDjQ+avhYUtU8rNK70oWMFOEgP6SgNme9NcwadpgNfHTajCo8L5I8xDayNl
padkMnB7zLn0zuSpV4XzxI2aTbosGm64IK7AQcJOCOpSrP20TWlm38gd/3E5Q/7i
X+R0zRZm+KH1a0uLsuhEzF3BRKCfkh0Hbtm3XsNHzuvRU48JN0UWv6xcbfiGEw5o
JlOBQY+yttpGVXeFDAwMRA78GN20c1BcMhIK1teAebi+Cu68B6ryEyJwFJnPUWG7
EnbCJ4LKDHRPn0pe7MGrmCmfRNf2TNvux9HuKWQ0SkoKxHpUik44u00PAAtUwb1z
55oPnK/eATizCM+bM2+j5mx70xlCDpHTp1bwIt2LEeiN+qSUIopoT0O4KAx1XcsX
O/sNKx758C04ZTt19o+XfVtFIwsjgGcwdcmfPCH0JsP2kVl98XshIjEs7+1vWnPO
DMHjnmtGHVcNIoEsbwouCbhFRa2iwvXh92hOQni4lplTghsvDrqNP35Nc1GnAV9B
sR4zOE5hVdFhBNtKHbp9IxFju4Ymh5A+/pe2n5IB+gMEvg7UItL7lYHUAQ+d/ZEj
bKoFu6ZSc9aKnkSw0z9Jd2t1HdMl3xUVz9Q0neO2egYffGZBxe43FFbLjqVNC9xv
Li8nd2pODPCU1PZZkVKpYxXduHqmS4Ga+eWbkElLQ0J8fxWEtQaRDj55EISGqCBA
F3ZwACctxbIITUBzRUF17ciOmWrFYby2p23mZUnyKRS1mL4QHiD8jUJJBoc7Y1Ed
k7L0ygjUxCILJtd8KUvINryV6GfYSzNSZvfPUeyBN4GGFzNvUW8M1vELTmpM/bqW
Bf5LEFvP90ybUxVBi0XCsMD96Jm7poXotjBwvE4nepk1F5DNuS/01dpE57McSHAz
IwRXBSqubUR5lbRF0XMc/y/3bvMDEJZHYzI9iV0xZILgRKM8K+ZvnH5PFZQcd1op
fwnLptOZ2zj/4q9PTwnLnjk6Da0CAtmkRTOigTCFbMc5Zqwg1BGFePvkH2Pmdidg
0q0jhIQt23ZNDoSloGC9zkynq2xsy9htHX1yYnn4BViLWpMcQxMweYovm/MnPInH
BzVQfJRp5Yfkqf/MhmloYpM7OX9oyYefxAPVfgho9OoPoPQbumHC7UrwxnoGTeV4
WtgWT01csbWqDU7gtLaX8JgYxhbw/zUgt4tX9tZ9bOxywH57paXgnXlzynnd5aJp
l+1/SPjGA9RSDZcLpT8kOIrGXlu+c8MNM2Vo667HXpKsvBbagUAYVMqRfEteJdqR
uMIa5/yCN7YDmMC1w3RdqsylAoVXbJ12AYNY7suOnzUEM9cptInEvkdHryAy67p6
yQ6k7xbJijEemNSrJyzJmgC0PpxErWSXpJt/cSXZbzdkdoDR0PRJN55r3yb4yCIk
OSAlcsqe3vYeaRupGG5cOF37VCHLDfjSFGUbnKpSwMA/AA6Clnu/vZG0tiR3rFcC
9DxGN3KZRn7tIAnMlQ0SQmso6ly3Dp8oGmaJyJHhrxR0a5NLxV4ka7KkkqCBCD0b
GubsixIY9BeuclXORxH4B72cc8a3pBz05dk91k031VxjTDkwHdyCXw296+A3JceP
J1G8ciwMj87CisBHVqIyaHl61whx1a6j8YuWSPUTq5DwSh54kYxVl6YCFY8SmOb/
L8yuCLtJID/GZrvirm0Q9yME1x1PobtAe9FeyDu/iXkt2po5fndvaWKyAVfWYKzW
gCXVfr0EzEP7xY5bf4vdTTGMOKwMDpb9fqSXqC1WpiCOKpaV39GndFgMxaa3iYvG
rt3i28TE/xwYeuyIQa0teKaDrUiuFxrM8DqWTOsbPzJLL51fgLQ0HAQMO0AgncAJ
EPmKmR2gsaC/wwlYgy84NPgk0bJsTZbEn6kH/F7rw7mi8qu8eY8s8YwYsOZKedFe
ZIcpis2y9iaLS2v4KLwbCmkUsLhTaPRmX5tDHxi1EPPYUvb81MHzUFXy9rItQLid
EI85o0PFtW2LFK29d9vrEztF+w4auL6YyFjcjKojCc+FJKlJjk15xMgJGr8qdSY1
TPHl9Q/RzzfOJdfYfNoQvwby+dmmFVRyfW1EAOZAwuczPVjSULXjfon2/6UtcX9A
utgHB0RVbx7ZsS1PikIxjbIhUhDXm/yKFQ2E41Av6IRjX47myDy55AcVVeNOP3WE
DsD8FYQNnFn4wfngu1Q0JJz/tJuxWP0dtErXhtsSUTECI2fZH40qBbg+LOhk0NHf
jcoS+r4gmERHN+SyvrBjaA0q0mtMi7+unhyaCwogmq7MnDckvfW3bamWiBQ9EB9u
3sS3+VrUByUVbSgYVfzJu1YFSZHqw/24wp98ta9Ap1PgJ1mJLLiTT0koz6yPCUVU
kaFz+IihXgmqBv586IYDqeNOodPwzPdx1D1QHTPyM6yhvPq7AV0q/q+GHhJMa+Ya
kNXogoNqdFIQEsSk5MHEXj+pAzBfzUWtB1HiHKr5oEeVZEMk3u9vLIn07JxWM0cc
7aP1QiLk3wrxzVxdKti+5ksKGRf3GSmXCm2X+vFodflySBlae0icQ8C/qyeZvmck
iOFb5OBhPApJhtKjPpyM9ivFQ5QFSChXilsp/ew+XNcCGZxO2bdrowyxlLz1tS3O
PTedKz8itUQcLyqZiqDCMxFMvXZ0IcqYpwVFhIJtTCF2QNqmsCji6Ge0yOhXJvul
cakCT/3D2SMsSLdqok2h1cpRX7nISmHv1fFM7Cd1Jmuk/BRTJj7Sri01AHtzMIIS
3Vm7cqfK0DVRLooHIM8p0Pm7PgJRr1nvWN3NUsA1liBHCRUkwWSpppKExPe4GY4l
s1i+gJv6NS+8jjUxwzOMJAmyB9wL5xwP/i0cmc6Q9h7NGE8VXSPMw14qAD8vaEdM
kiMQQNxjV8DHQSWeWm8HR4fU0eZWIsWFTp+Jp59QHXQeacLHoQJ8CgA/ZHLYORQ9
Mvtat9XMn3uh0E7KGceOaqZ+4tgrG5nb3vTUaCtEwJrrw9+o1293i+U3rA/ndTN5
1R2FZtRQgqMQxnNxCvkvlNumSec2H45murx5FvPx3mNOcwO3gBtSxK3RTCULjknK
KtlZ1xSzYjkCifMtxb0/wyqtAUDxZeHIydQRXxt5EjtduZgNdkItKkNYj3wDpG6Y
HE0w0ogk56FmilSkgDrua1+44VS9ur+9M2PzezGqYPxdjwMm6H0265HL4HqudRz0
AtYHLJM0H1y6ZBNJ0aCh6BxUfhidMy2SHSQJqrUVAH1Dki2ci2lPEIhhYc6gOtrx
zjCGgyCHbVm5JfXrS+I3pw5ppCeUhnaJMFDQ0yPjA572eJmsunaHvLCG/CvFuemA
zmyJ0rjOisKWZbZgcq2J8v7+SgbnZ+7IY2JPPXokLZ4LpYTsL22wGp/DM6w2Bf8O
CJtgl+dmsWHhxVaDtDHQc4tio/YPgw8qKAC77xDLtJkzTf8x1+igZfE174KOgf/B
Kzaggc1SU0GgykiuFaEbpUAeAsZ4YFh2q0rSaFhIwc832iKTTxyeTRIOic+4yNFa
ywYEUYiOh3qtykpv3TA4IIKr9e/IeRu25cliiTMtSkYwdzW2MfsvYWjdAfwPczcw
9675/objYloRF5Hn94TmbSSIH8W4daI3iOl97ZxPJBSlxLEX3TlRkqicOeX8VAXe
O2jn+w9xVdQwcAmwBThUu7jIfSRK12j1FJyqIA1Jm1pNstxIigmUwK9Z6z7XGQHe
4FWxPZzKzQfvWgqP9Y95ip/rcxkBqQ4GvkaHEjLUlvwVFnbTzDxMFt4AcheTRRaO
00Qyq7wSrwskaf4r5nEq3GuvtFdDuTaojnGjhH6WZN2dx2xOdgyHYwilkiDQhWxA
iUX3tvkciRv7yNIk6CYyjkMShKHAyLkyB5UD2tRekgi+Ov4hOR/5E9jVzBtICdxl
fwtgMCQVUad3nn0H8eqD2HrC7FIrx5ZnCYM1x6Z92XDdLwDwr/lMdTQ9XqrwwgJy
VkJLAzkzvyHD8FP8vf51UvfWX8WKuPFmsOl2oKZjZ7xAjxaWnOFeQAQoaEuwTUWt
f9k5bvY2qM88Q+x+N0+ViOcXXXKqG80gqQzNjQvPmoVXc4TRRpaBWkrJgSZUvlI7
p2iczYmABAv4WWlZJsrUP+YCnwweanGdTRlWWR3YLICCJ8S8eXnv5Kx/iC8BSVZ1
Vum0XcVBnbYvk602bKZlxLMI9DfoiQUlejqe/KYLd84klJHbWVtHyn7WzlTf4aO+
mkqOnMuGdu/m90LYJxXeIiyCJe46Nh62ClZUOckT9eVNq8pNCQAOJ2OHPzdq+7RC
4VsqzTiBJRpi2kigL0LXk3CXipwHeTQhSuWKoG4qFaSqvYmmETYap73ulc+SsOXH
URwbGTj7lNmM6iCPbKhwtgFj0870k7qn6l2qzvUY3KJ+zmwKbiNjtyXzEqVQAzui
oJJP7jIgLWQDW7XXHi9NTrTbXiI48o1oGSXMkq2IQvTiXe5nfxXKc/bAv8s03uBY
ImVrdubLmpY6oj6HBCGHntlZpXDPH9leXrGi2TAL/GqIdxoeF9/urKFSrPkf4GU6
En4tDuwiIRgeIUZouo4SxxLA9ouSo8/eycIjc8lj5NqyedmFg/8KvpeYR6BIdEIg
JLlsmSUAkso4lu4w/9YyGy3g7KkyfE+UFaLP/imK/opMymgHjDdjCNEm2O42DCzH
6hPRpxnTap/33MmE8bewQryiJwPPglbt21VKb7qaU+BCNpYNGh8fKnoiyA4Z7Exx
4T9jvSjVmfVXkYshOwpWK8K6JQVuC1jTVmgd3PKWANzQ9Kg4MU+EOozSjYZPrvlV
xxEYO0mShdHOZJ7/csb8nQjtrR6PvcMbpHsR9GiUhcle1kEPIe1zpS34j+X6gQbe
sP2U5KRGGQ+kLNL8fLQnkI8u2fd3u/HefyZf9BWOmz2mp4t4VSkWjnSGRcv/UY91
iddKiy/3O4HCjnoKLwn8Xw8LtgDXpQaIEx6kF/Ns6bK1lviq9BAmfhDC6iNnv+Hq
joRPvCmWuY4+aRayXkW5vUwpqe597bsTCa4R5Oe6cnId/zWoOR+gBU4ksPMDAHIX
doLqp5GkYWW8//2TmDe/5C9ei1Spa6Gpp5BzTh+m3OdzmhkpM0fS6KMQd+UErSUi
ksRBkNJw17vYIXfencg6NUB92BteV9o20WmE8hjjlzSUe7q0P6+emdtiWilNUbPF
V3Ks58jWuIzt+l9Z/VFtDEiU/2NmdMHOo9dlGJ/BtQScDx4qe56Ua5AcN/7dDmuD
R8K/MMXrsjaOparJbRl5wz7ot2vIKgi/7jIDH0qGFqIidBtBRSsgQB9NpWjnYrTr
gyLmLCujt8+e8jW+Iabar7zLDGA4s+e7DvGteI+4T8rNk9U3utS4Z5PBU1nXbPxA
avfdzILVpnp5GxMRQeqaqZGNLY5lPVW6eE2vO6awE2qdvruYiNWF7BvTTA9XHPMH
tcII4kQxZsyZBsBUITcoSUvDMvAdDNdEpyBGN0R7vPnm8/bcxReVV8G1fjOzC+Pm
EXwIxjZscTu8dmxSERWoWc8FT0Tqas7MtHV2VrxcoxWUxvAMaGDTVQskNYUZt9e2
Roif84Mdhp9XX2axO0EV9YKsKvwYFdRJbWoV7Uto/px6n+qLm/AfZF8RuD1hYiIY
ces7nLQUqlr4e6A+1Xf4cTk02qH+ytbd6PAMCQ0wle5nyydUE3c7cBapBxM2SdBH
G6NT8z8qELPaVeXPxuA1oEkfgiuJVIzbJ/9Z9IFLhsfaVZSZImDkA6nJAvxEgfuc
rLZ18dlfGUu39bW41Ki1i8CtrJWndX5aE8tRnkOHfMEwSHTfVd37S4ekmE50pBh6
xMIjK2KUpoQ+xAyM2hvQtWmsy6hj+sf8RnPlUt6KbQ/nw8/Vl0aBlXmsCUKYcCIN
NJ+pJ2jeC5edV2Ag0YT956023e/TN1ip/i1RgX0HW9OA3D/sk0jSNKk3uSeoxok2
v6VA4aRx6WlNUkV9jhiGbHprgBJdkG3R2N0zA+rU/pdivDLfanY9Hg3oeaD8eNmL
VYZRVH5buHs4FiHfVBMIW6moSg+2wvctY/Tf0H/pRhafPIgqOm22rpXjSR4Slqpi
YY1d8vbrOvQXLS36g48irIsSw24XHJPuwegXUY5aYYBqzlReORpOTPvw+InEH1Nj
peNdLS2F5ekkbNAm5AzID580wDZSX3mDKGYkuY9q/Vi322OWXY+QcIu9eYc+ST00
vEB6woonSBo8P/+cTzHAgTfqfP+fPTejfzSLupyVHP0ezcttA2u15by1Tdsy4Oo0
B0wpS/NGC726n4Bg8yRwWFJun5cYH+iG7/Zs/p3yhA1RGXTv1AruRtoMoL1ylSrL
gVt28vzCXt2y0jxNjMuhivabPrXS+z1b6F8IJW2UBPzDVmW7++uJeZ49gKUDHklO
VjmwkA7DeEdCyn0OcPMvL1PGVn/E1gfoOdH671S4yGYaqSP545nECJf39K4UqUOA
0DvWoWZVVqGnaFwd5LgJurhFhvzlNMHuXPL0+ZqbjHDBkl3dSkEdxN7auSpAc56D
vmPwRWdOEIykkzBw9k34DRFpVH8+3vC7gN18QQgHdOlDVUxAfHSZNdIGIPOPS/xD
mmnAP9DUxnd4KFewm1t32HTh65mX81uLnmEHdR37TGmeXrbQP/npxYzRMpKeN4Iz
xliAUhpuIuVkM7NricVJCKXii4lHmPCI0Pz/QGH1WXShWR2JdPBbowmqcpF2kzua
k7qHachoojypQ6H01m87j5LHeb17eqb9dZR+A6ZeTu4wbcldRzdi1Rb5GziP0H/I
+B6xmXhzpqvjW672Hd9e2bIn8XAsXeogsITAd0rkre1EPePnBcCBfa0txd3LGLVy
8qhKPS2/YNjf+pSuB7ckaCVPdJSy7TXv/4oIKWc6fmhVRl/sGNdwrbgRP8E5EIvS
YxPfW1a0f+LBTRAj97AN/BGeeAPFt9B5ttEBIMRlmGitZirPjzqaGQAAyCvupmzc
LirU1O9UaTNI7VmluhGhWQ3WctNFeIcUTPY7K/nMwK/m1ZKYBPbp1Zw2kHTUoFuH
ZeObGcUzYt/7ziVAhRSFivtfCFwiNXNg6fGNFC56+MZHspGLRAgY0w3DYvAjtKu4
hgEOTBIEUjRveTadKty4kPB9YSj5++qllbSn9Nya7C2GHc8d/euJO6TbqZOB1gbc
Ucs8OyX1c59nYyCtOZpEkHWHb02BwSwL/GY/C0SNbD36o3H5Pt69nph8HPhB0rBM
KyqyBMpuDb8RTgTbbs20lW4l/zqW+H7yf2GUyczSv89GR4eubvxUHQnVmz8l1lEO
N6cQpUBFZ8V+9BOD9Rtf+IME8iL7GTeKH2SRMUH0lsZgyxofqg8o4sOat7T5a5Ca
cfNrGVqZhTA3kbbEEwCnJFTtpnPpcqj41O0mf71IzbqpHj4QtKWJKMTU3xhIC+lB
helUaClOvlFAfjAwOKvJ9VhGwOXl+1wdhT7JVomUnqN2u3aknze5RuXK+rvJspuY
QaQ2WN07ynZ0BCjeelSNp5Zxj/uth63cKAi0bXmPYm4IKc0Mo85yvCwWKAeCf0wc
eZi2gyff2AFSkoQtn7b1DSeOybTILnHFnbwDzMI4Eo+xvUv/Qn5FYfS9af521FQG
e38Jp+soHeLJVCM0JdRJF151jSGS+tzHfuCD6U8HrWe3c+QDTnBiUEzl04Or33Mv
Gc41B3WuDEo9jTWjUwFn978dHMf2BArMPm5ZvJujYjJ3uMcNXVGxS4/Q509YbWEf
w0I0Bm8IMuEsk6ZNxN32WaYtmYDjt7Qp39kx1SiN3S+SLZkscLVU8NeACyP0LGdh
PFSDc+a59lTPAPo0sMeeY9kUPZvRWlNcbu8r6SqpeBScPRGmDrv2daV3FCrUM0SB
/b1nUUgu/vfBIaKyW6NBcPT3e5R0j12HZQ+eUQinExcUr0tzVPSWL18ArV0vuB4K
qbtUjp/HKbBxKhnEvtD//cMhJXA7VIUTxMIU3nm9jPS66+4kUtgXiQmziur9CmYH
bHfWAvR0D0fucRHNnuHbu2laqqAQ1NFJU5nx6rPYX5dknTC0wVD7tcMSsGpEnA50
kMBOVKhbH0jpOUx40RPV3nkZYyrErq4UeA734ezinbj7eQXMbPu/bS4iujFPe3BC
PG+GL9eLEdPZMRORXvWv2AEflKc+ee90/DkdYYLUUU8jWLgD2XGtEKwGyEFZc3v8
SMFgT+hYfVp5wUE0iuLwOw6RJeOYcId3T6iGZrMkVTUtAS7VUajLu43St8lS7BPd
J0P5tBrUdjPjKx4y9wWlCodC4lv9lcW7YujODMURg6znMyvZD7uw725Hmax4l7G/
eYSwbemdYlMg1upKC9JQ1xlHwvKWzuAyE+/Wv7m4unF0tEtnd56PA9AZjrWQeKpW
msu6N83OUk+Bp3KtVgJaEntED2OoKiFR217AD2tHoy/lhW1N4MfuJ9w8TSuGXYt9
NV7fsroEsPIdkyyR3aMseUpSSz0Qn9I+xXp49jbLIqlXm6VH9XI2PiyviAxvCaU8
WaLrg9uhY64y20PFWrxN41iw3XVg2t9DYkvTe2lbt2o9ixZuDsRotfrOaoiI7O+9
xu/vlmFebe5TbWD3kuJzItSN9LYJGmYuIo5K/bomqpEy4ppWMcCDeEKMcgnzbP/9
OWoA4DCnWvLbiXiNFmFkywFb3NN6keOT34EVAQ0aCQ0ROHo5QeGJpVBrEWxI54/W
3iW4K35ytv4DtLMxeoaI/V8Viye571s+Aj9UIJbCt/fHnIUzcEGQUh+hSudddR/v
TvAY9BAV+OkBrJvw+c9rKYzw/F+EhRCSc0ybilWTSXw5w4Qig9vQHkn4KTeg2C4U
5VMFQTD0gSq4ZeZIOsigI7xQrzEnNrIQ44anVp7gsaQ9wn/hVe3T2fbxTWMS7UA+
NqD2QTvWYQVfcbuGgxMxp4yHzddN7wxJswnJP4J3dY6RGu1DZRqkLmUXWDEs9EJR
KnakHRj9o9HI6nYk5IVxgQtePHeugNyayd0NHeBIyLf1SNNsCxF4pQx5ogaGSf6n
QLmGw4Tc3ruwsimxZekzyY+Fdyyzk5zFTNJfYG/3OOb8miUYSkh8OrjB6usNGiNG
Ahk/DXnlH0tEQdji64BPvtk7UwnJeC0G0PBumdXwtZYU0ggpOGfkCvQzjeLfCyZk
J4aYINKHm8X1JYu/4AneQSZOFSEEGrY/hoNHqLg8WsO+jAUASWMTQjzsR5UpsIHY
/JVOckS1B5nhec4A/F9JVDfg9bNqd4NhKd67cD4EXaABMrkks29XEwT9xPHb9ICj
mH696IbTrSp7Mjz3q/N5tS6O9etzVZD8wSXwVxy/HrC6ObQaIsig3pMz+22YsPCU
VbhrifVPWD12HyQoA6zaiDAmVFzL2hSDNJ8MTMGhEKmO8zT+NLM4b02LcqwmVIRw
F2oBbH7JpJH98X4koZrJVilPBLPgG5VzLtdoJhaTbwGr8bFt+dgD+fMcYK3Yyl3/
2XyPeE1QHH2zlXWjK5HxihDN2A9aXHN4lsMwfT0ww50BmcyCqJw4861Dbri7YwkR
LIpDaj802f/IcnEqZrRCzWTwgVr/Q4xL/RcJPNsGvq3sZmtVlgRCyvYxnga0/5QL
NGER8KUFwlp8jVqetJXoZkKkkmPF9R/lXZhWXdg799Aub+d2ajxhr9lGVlty6TW0
b4OEiKb2mKCmzbpmUzPF3oVFcRJBi4YyGMMhBiSnvBzvjfgaU/+8o+px2ZMaPgHo
7hqPiNY/J3+4t94oQ7uEqOmzVviNzemqU2pW+DrPmq4osYccUwkcisAuKZV8bMbT
xCBLKZlvrwjfIB4oH4b2tq5//pJvCfJlSxot8Cz7tdqgFUhH0eycYMfFZ5Fl656Z
Qw7j4A4fuhd2LWCk564SaH6TI4+Vs//9vkSXK2sf4AiR9ivhGUEriyJc5Q/X8BhA
wdkbYuARYssexxPFlzqvrnTTwASk55TxypJ0H6AVgSIEqvB6sJqAbDf2MvXBhPmZ
h0dXlnq0f36bxoqFHeC3P7IPgGgIyiGFWvLPoHMfvjHXXDMCZ3H8FSLUTkGMzy3g
IUWt2XCWK09dATIy2kkrhqQ4xbtgCtsLCERZmEFwoOkRQCAXpmmBJzzXYnkRio1R
EriiLXV1mElm4pR7osAV10PEkq+7SVMTjvI8fhYOs9GepNfxLat7egHBMCbroV50
PLNL6FjCIYSyXcLCfkDf2FJjF82SvAQuCca5BK37Da2Vl/NUY1wB5wUGUPZkWgrX
+uRvv0xhRuZ7zRVNNDRRRjgmqx9GIxr0IV2gxaaj6i2hKVwFS0CAWPFOdbJ0i2ln
BnkPO0A7gZOX1bs7sRXF2nAx3171/2GJSMtqtbAZ0Ta3B2RYi+TNZXbhyPUyxHPs
COn6v5JR0xqglzEErRYzHGtSdz8258OJzlsqpdaErjsE1BKDRb34Bcs/7rq1i3/Q
gIvAmfUqhGXisiLQnMKcpZODl5eW3y/0TCyBA853K3JjMcJGz/pL8p00sLXCXOdf
yuh2vfgCVTxbFHgoDBx5dYBe0tgHW8skyjFbjMEVmFc/DuZTqLdCnh8pSbK6AWXL
S/R8Lczp74pQw7zUVGJxHG2atbO3MAhR3uuAEN6LgtxxrmLYPnmmJxnJ8Xx3vMIH
Lp9/+qzsONh5rOHBulNfKB6pQqoz3DAFwug1daZMgFGirYfhN8vQOxJuikIJwJqK
+yLM0YN5ZRXRQMlUCUKq68MkRgLvETPohWhVtO4i+Yyq2MYyZagxCKK+8onv6p2s
zS7sjcF0x95pmAv7JlVeTdt6M0+RtDc7uvACoPjqOitVoixP5dbkWeTQNPRMOFbz
VSS+hUsLVVzmSmhUO2z6NEPX6EqPhUfmv8yFRiLx+jgvA4Zbp2n916Ems6zmCyqt
KtMA4bRD/mRldxxQCBf1kLVYLkLGLikfrYHUYjBnWNdgHdSGQqDDHvSTVkxmzGX3
udW6oTttJw3tUYpY5OEeju1n6y4T/XELdwFWrRT4ryhRhlJYM+2swrnmxQCUJTI5
LlAa4ir9vwJKOI6Fp2ZCEHgE5UIAHg8Lib9XS+fM73T4EGcr7WkLP5ZH4ZL+iewp
Wt/j8TZf/YIVxgNxlTzGreSWtslB0xsvRXSR4USUjaR6Qkv/FVqux+9EYYFPJtQs
FkT+VWpuo5dZK/8KKp30ThVzqxneHEsH4gCZ3bT+QT/BfotMELQA2Qv3Mk9Or4k3
4gVHc+wyvSZmJ5DjLTB0X43YFmEOiPXoDObSsXJOU6H8fmO4s1+/Kkb0ubG9x6lS
P3BklUPa3t4qL2X4JBOR1HwEWLPQp60s3dvObrs34rfqMWxx5we0KRk9HAk8hayu
GmuSQAPJEqw95zloC9q0L0l5iUT06ob/in5Or0iUnzkYk9q7ZbwSfKfYgpY/UMGG
7t40/XvLKdWW+v7EEWSAetb0EB2/SKZiqFYK8ZdakRENftH0EWhdPh6r5RulRT+d
GIs/xBW7QbpLVvuMumiSPlC7pqU9BwWv2hxfBrW0KuGIQC0N9OytTGVaSaLhDQw+
GO8KxX98AqU9waZN7vbmXhhkGllM31oFuUBDanQ56+WaMv8VpM91AUZyn5KZpbzn
wzvUmDF9VoOvmRKAYl0xhTPNWuTVgtyITcZz8fJMOKxLSTadZrqdHBeOkhMx1Pak
wthBBYA3rakrA1bGs/7rkJXCgUCzEDCbLqkOvpM3cv1axLPy5f5zHx3nHCXDWT3K
w+bKATYNe0gwObPPSI6yx3CwMW8lESBeeYMlpA97EoIJQFltDEl5JHDiHvh/1+dz
vqUSTx1HVeh6S1UNt7Dqwzyo5BbkYvSZGXODWyyAZRqi/9NghGnPMn4ETH6QOfmp
G+FXGlXzRFEnDfAeaQklEBVUDFAowM1NHt4YDEuTNnRoeerNUL62mDRmT0jpBp7i
zGeLe87XlszGdjK+DokD+ldPwRS+xgTehYAmP71Ly8RWec7p4y/geJWbsBKbXnMX
QLiYNBiObkXyU2dwyVadqmhI42HEauPEk5AoaRYqN1Sde5jos8oR+WYgAfsfmvQZ
7g2pyhaNZiGJ54HW8ObAgN583i/fxodMxbyV0VjQSqGQxpGn/rC7xtMyhsxC7XAB
AtdIIiJjmKDRgPMBILjUYed3I9Wy7rxhgZn+8YDuxHIoCjCCM4Yc9rgOHUXeYyWB
lBdcteM94a9JovxRSNMhotivZUkoSQN8L8Q1YH9+TlRt7okb08xsY+pvy+Rcg9lm
9uW3taFc/lSk02Ook5+8T6bYZWnb/oPT/6Y2UZQO+lIOG3ufKoNd14Q0B/iCG+um
nkbQxB9bzx9iUxhGw5kyg9qoGhdtNFlRb0mHk/oBu6cGLVQDx8mRZAKt4SGw+LyS
qkQu+G4NuG+8jfOP7wo5w1bBltzdVLcqenQEyxeqPoVRDOq/jSq2THzfsigzVnt2
lMosMUvIdNhNPF1jM5cTaWEGDUq05SKFJtPSXR+49rVIRwQ7NGlFmGGMrYTzwBhk
SqW7gPXNbXEW4EjaijxTrS6fKm4IN9VBeCISXD1bhG+NI4DrqCabQ3y1D4M1miLC
jGt49slwRrTOQraUdVcloTgWEy7RxUm2yOe7Vfdy+vHHgHGr6i1JEYgQlFjELjAd
wVQs/de+Tdvw/yxMx9h7Fs3wGWCIaZYWLUba86SCw8vzlRnEJ7NzTEPlz72JbKcL
5uWWl+gP43Hg63gfKqJ6KI8ZkBARXI3GkQcoNvYymYLrG2VVnCpw1S+Q1CqkN/4Q
9Gvg72uVhSGair0G0rSSKY65ULXxxTZi0Mjm2kz82a90HgnnmzdIvOCLWkiKwNek
6YRjEastvpTO99ExLQKLwvRQUdMX5Y4uhjymO9rapL6WnkOtLCmNlrOcmpui7uoa
tReuylr5QvYeV1ZE+lOVarJsD36PUPxUiPxmdGWFj4qUDDSZujJi1DigRPZgn3l4
Z4lyMT2xrR/agXfok+nbLubphyMx6v1DXqpBZWJwHFJ1xmPjz1Ci5huC3nIdslZ+
6OYJgb3ZX8oEMkDrrL9JSlFWqdfnj4Ik3yLO/oPD6G91Uf2OOvVQoXVVp09nKPdp
be/DDhyISG6+FjkQoaWvfE0b2qh1K2eQKI/LsSFE2N6+aYS4AWxRJ+Tz8QLZnCF3
K6MUXgDy0OQDoc/Q69UdVj1HE09INBVBQoeh2RgN73sbVjvZpBLIi0GS5gGkcZEF
z8K1mMLAe/X47lggRs4so7xgparhMEs9UjjDOCQM+FJFRMLGbsRzYT2j2RCh9vhR
/GxMLfJnzC2/ak/fiU6I0OZNrjT/+S0zXCN1EaQYDnS9nxyxTeeQk6s3mkoOzQ2c
CSEcV9y2GaVwLHFyMmKyuakgICRbrqizRmrXs4WwKTrxFi0ZhSVdeTtt3BZtLEc6
cdWe78cAXJ/Nxh7lRxy9U7p1o1Y5pA5DNGtVhKHJdpu7vD3wHcUCX9bDQ5ig4sTG
RVV2VmB9H2jgnZ4+vBHoDldNYjSpTFuWffVgiHBwIw3a2q0EzQJxlp+6SjTu+sbz
NcZFzmh23Ywr5Ld26+9CFOVUBxiszGWv6m+PMTieuSEZPPRd5mOZ/z4NDRJrCqp7
cnQILfqG9FnXKvXYZoNsyiK43e1quKiLzEuMVxeSkfizrpjcvgkOCTmr1kRtA3Ei
FW6Z3snaET1/LoEKvwpYTf7JdbCMKkm8YW5aP/aTFkSb9WoPFft2izxx5UKNYTyV
glA65CbnUmavMSVBQtlNmnuuttUkM1TR461XoY9/NgKnnCp1eRvD9RVUJi43ZjA3
29VB8byhvLphzbNn1k9rm9H35Z4u28C5ZQCO1KFmXWOAwWlN5YUjVkBegMcqqTyx
dSRCS7E/bB4FgY138iigFqSOGRzAYcxCuiyQqdLeijzkf25xpgO4Zu0Pseq5B4Ed
RytvKBIXEziJmwTUKlRyIhk6XOw6l1tHnUfJLUOfwlP1DY4sYGFlY12o4NZ4d+aX
iUKzqm9sBjNsmovBcC/pFVLKZEu1tQAp13ghCBge0ZnmbfgV8kYo8mBdspCPUVUB
QM6O/ukaDPQLh8rf/mEn7FEueiO6vdMsLiQmFQy4X82VLCa7DtWtpkT+d7spuZsa
oqa1rJuninyKqZuY7EoFvz8yR8U0MS+v1E1McN3U69U6mlIRd4S883L8k72UHEI7
kLXbjGsYaa6q6PCboz8gyZnI+6VQmpdr4MWMOxnfY2L1lxR0RczBVLKWlkJxlvk7
7G+n6TSKUmzud8D0xV+k4hzS/OpAw2Q1GKWTQ385BGkNXBif9VU592sot9tVdKX6
gbOCYhHKdXWVsNdosloGkMe+fDsjRGUf4DSRVJgwJEjNZKhwmoxBr94M5taqAgjW
ULk+dIy5gGig8iKnFZYMPJzXDU2YJv0aIum95TquDEeQ6fOVSu6IylU1yIuP8yUU
K0CmBrUFPgQfRdr8Pe+qLWtp2lCZONYz7/L85qGwnKkWssusuo1EIK4IK4B6oPpL
+ls1Nr9v4VM07f4UXpF/4/A6CBM/FbBk/dt34QfJfMxmQJdZr1K+mWxP5ozrwX4P
4rtVEIabuDcyepApqc5uyC+Ag5a7jMYzHkNNmRcP4rtt3dtWnhLKfKUq9gyoTFI+
2j3E+VeDGP+BXPrkquNKtLoD/hlA6afPnwXor4AfkRTgZwPdMvicvHqTNr/lUoHX
eLppXtBzH7eKDfNjfHZcFcp0575xWIq0Ir7BCVjrLve76v/vNikuD1v27Fhb/N9c
vEJdsdmjU+1qdDb7HTBMLhPxPrUao9yp19A8sgBmF/Ss+NUrP017P9u4vNnXhoJ5
m+cobZnRp/1JH4evwwtpDtkYh/ZoMarAd2UleSUotUXglEm419Vb0Sofp0/oJRvF
E2D3J1Gv01hgX/A0lu6G6d43Z63CxDQG1GRcrSJrsN2SoDkWAdrS1LsF3hK/Nz2y
W7n0kHxyy94H/fdmfScDDvjqEHNOjbeFrRc8ZLFY9oi9FeGQmv2mmzSlIdhlKilk
4EpLN2ZN6l3n/7IZMltRu36t3udWh4BIeJXefrMkfHwfqe1e3vzQQx3YtjsSmDkX
70dqfqOkMEY/awQWIPncJ7mGdPNG9Kzmz9+tzj6XnobL5YlegJYvAqoLcxqiOcte
/BPijAW7c1MmVdwL4MU1+wlNEFa8m/nkKsArwTKP5Z0NpxGqzbscqiRw+huo6qAL
ea4DaHyMZYwA4aza1xg8VSFTIuPnr7Gksm8IazgaGh/snKRmYFZ6qVFAlE/AUYYw
U3ncX6gRAKxxs5XSO9ivFkrCRSMtB3sf6zbdcYldk2xFX3d13YLw2tKHeBwQRVPv
yvB4mWy/HlRpgaCrNWEzbgnnLRZGOGwDjIJTSYHqIJuQu47icl65jsqf75BfYJfh
iILO6znZ9sSTvwBVDSCN1w0aTx4DorxTLwoTqvdt53xLbbzmktYmJ5fIWcu0ljyW
pxmvXlowyFEpoehompZ5iM1e5paDC6/qcKqLKViu9MzuHN731J/MVO2u1j7U9bZx
KaV+O7/Io6Iu+QTTrm1RjEc2W8Lnz67IymkvYbTTEUqHiVqc8I2c3kCUy8ypY8AO
SP7foaSwS3EuygX67/59ziHEreEBFUQJC2r4GlQ0pR1tcyCLcy1WFlmnf5enqetx
33W/69+a/64UGae8NyTDBJCCWbbu+7I/zo4Pme9MRdUKkf0ohPMliTBe4uBnDzjo
Gdpj5xf6mnAQUXka5ZRr91OzID8zuu13B3/zjMO663XskQyB3qeK/TsuBOMlSy9b
U1h5gHFIRdBXw8LJJ4hvpi2cn4NVLl/ecn5kR2qhieuM7rCrM+3GfWWSbrMiPChi
CpGFrF6dZM0nWiWi77UDvo7J0WhLMisJ77Mf6ttrVUmXa6ZpD9oy9zTftABppX5z
9MS5ZVnfadyNTJxhYSiHaE+SneAOT7lqIBN4Kv1Af2r3id+Hu6y/4Sb41DOblDlc
uTi8LFuEvdw+TYWmk88HYkQVFd9nrTQ0UR183pBCQqlItUPVtN7+TIBYt8JTiOwK
VD11GhS4YV46zm4K1PF5wIQ9aD/zzjWSe1dsBzthyLfCumr6ggEmTnhRA3UUt05x
IHkj9uCUcmiuS/GYAw5+QJt3GuCPqIUBiqgkghwcQFOwbEaKmlEkq/vKdHvDrizp
gbX9rU7Fudpk4CM/OqVQRlpr3nmQenChz6WYHOatuwfat276aU37DcalADfUPBxM
Es7liqhcPOr6lTb522jP3z4uN+mDx5mvbckslqycJJJnmGsCXAdfoxvXKNL2AAau
38twwS3tLEMLZdE4gItgSbtQkjUSjUaRqXHjgXAJLk/mdAKyouNA4M6jRdGQU82H
tRqUu7XNR3HHn6PlJW0QdlWAIZxPQRSxkmK5l3z1tsyoZhY/rwq9hlM0peZDVtVS
mdWJorH/GT7ubbgGxEhB+zFsGCYwHOr8BqjCwbPXIJmCTaNxd/4MtV0o03MsCRez
XsWK2OFZC1szxFmDjoaQm/0pUcdU2zVVzY7eI1Sk/w0qyTLrhHM4lTW7SQNYMNEy
ji4iPWprMD9paYXmTWvgb3r/yYIZ1OIv9gwkUVj+u9xtvFstviFEdyonajfMNeB/
b+oyNtPDRJ5eyzRKPxNfyB6xmU3aTNdjgEiBilHXQYWeNitv0jzH50MuSHy8oUr9
zLUCHXTJc2V2CKI701givcCcPAD6F6ugcqgypx6vnicH/s6vJ8K69BTgJD+HIY/4
OaiegyojYaNwiDdNFbDegi3wKp3XsmjIuCfWq24HVZ/To8DLUIwkoNPeqMeBoCDi
a0kq4p9BB79GGO0NLyWkrTDWZBzLR2T+j3FmiQOdVTWB1AbBBV0DS1SMITMwVF+/
5AUjjyamNVRI9DSKWx7lsSmHEvO/4QYQc9eVdJ7+o/J0slvzcEPhQ8vZ+3KqTl/+
nmyANbTkuWczyUTh3qWbaObUNM9B+uyWEAWWJHdjy9Ft5KxLBoWD4buPFq140RFD
KH+oIDoiamBcEjBVZM38OlcIgOcZJCee6PDYEEPwbZw+ctlyS+lnAp5PZFTjMomZ
xM7ZWAazerP2Qj8dGsUH6rruIJ6kgjc7WpeF3lViOgfJJfaF4HSax8J6LPvVYine
yBB2njygg+iKhqFKEH6qkT02B7n3+Haco2m6DcobgcCXAobgKGFZfLSvxyfmWxoj
pDR0Mk7z62AYxHoGSLUQJoHnAcb3hhPJHXDXqJG2GBt7TDvIL/nJeWrgKu2oQakq
DL4C6mB7VZHy4BvyxZ8RXsLUbQJDgDAX0fKMN7ipSqv1/ugCuNhdHDuvT+4iDJjL
f4BNBb19FRvmrnX5jeYDJqWiMEtkq0Dp4QrusU7+SXuRVynlaAiaLT2XnjyfINBM
6qF1lD2DxLL1Iu966ve0N1Lcq3UWo34x7b8FKZcxdsQJrmF/9B7mUM4Cb+1LrBgC
wj+zXC/HQpv/4obP0d0HFpFUtxmIN8KqBpTsclgWwdOAxo5rom/0EHiXqLOlCbf1
3lMhd5LoFS+UqjNl3w7FmIW5XU58z2DdVdTsDKz+T8FK3REZVu2oexe7+dLlGFEL
dIvsOKDu1/2myIEU5TKzb5GXs3aKxgnfvJuJFMngxl9+RfJAmnGsqQt3aAQuR6iW
9txpbSFk9qNNhc0rTMm8uu1M6hA+1birbz4ktRKaub1ZFuSaMmVzzkl1dYxQ3a3f
9UhkpQU/aTaLYHo2ABRRZs8R/pqLPxMafUpyVnyXfZgBmg4bqJIx/PW76+FwZH/d
OV4nH3hoLnCkAnrhmUOxbBH0zncNF+qBXKdw56Tz1WB20vZTHniD0ndTFl/l4jz8
F5Jbi6V2HvGDN0kvxWNey+lC5zjy32wbxHr9o7R/BS7qLtW5bmtgRu5ueTomPHn2
BwSxqdg08tp4gWi0o60mjYd/YELsgjhVM7Jqg1KszDK4RUuYhQ/NLyUTjc3sLH6B
ZFe4XvcuYPkBQSlD8zAzN4AtmF0T0tqUUzLNbztQgWVENjx4M5rCQIFs2e5F0P50
DTdYUhT7pkgI0Oge74kxuN8fJKSG73fp13/3S9mNH0E/Iq8MhddM6Nnoseuba2hF
YhTGWGqp4KuAo2U3CGrtkYaMqCdF15bxPcMgaI1oVK3BrSRthxHldxkORT+jVS7y
CCENYbwQht3douRr3X+XErW1XMtdE1ci1fo8xF9m0IQuxN7xZny5R1mI83WI0uRS
kR6iQ2rOKau1IJTyUQjRQbbQOuxRoM4Er5/hNmbcGhe/HitqgdgGvAEciom4Xkvb
PoyPnKrL7u+zSokWUCHVj8Q2LL+phIVThWoHEIpD13Bt/BxPUFSKd7SihRYA2P2Z
VuwzzFWm3cfSgDTK23vWe2sSBDHFu0cx8crWxqM5W6ItiZay444ro3jgXQ9Gyq3R
rTFBS3VsjCmMfIBefeAgcMnVeX4BHoej7fwuSYk0OTX3/kVHqFMlNtdBQqjYjhru
2Yyi8bH3zpCkcqPsj6iGnAesg+n9W86K8krBkryJALqNBsEkjBYwhPPIIHDywFU0
2egw4lyFeIeS9r9fguL1WxCIb4ou5Ke7W9qbC3i1TnfzN2LvqnMUBeOzSr9RZaHL
Xc4XRxH8jby7nC3oTCbE8YaRPF/chWwuASVRRZ89ZDPZ3xvi9jAoV/iPMcH/TMTw
7t9Zx4EBH4YmAgVaCEH5bNppqHT1LVq9Lff9VXPvIIcvH9zwOYP2Ywi388byjY1e
/6P4x5lrmg6J+pmR0DsyX9Jha4CtOl1pqzQj/IAVoAkzpz+vfUHMydNqNy7u7hme
8mjSvlSKbjyYJSJi5rb+g9PLgiT2B37eaIqQKSy+asXfA9Mtt17pqKZwRpMeEZLm
S0jkqsuewaP90lt9Xu7icxsUocGZlVb/M6HPa6yIojvY6JHKbITR/u8BTEjVOf8v
7H8uTYmVZyinuArqkkvEDFDxDnO7Svi/thxa0Ahp42tXEQFUbw+e89gPKH1EaU6+
Ka4U863ZG3TuBHQ3MoME6URm6rkWFNdN1TVOYwo9XbQRgAB1zgiP2gT5yprPUbiN
TwJvcaVp+1KXj7/4IQVRqBeScOOH5sbM2AlIk0WfuPhbMF1KecP1ZSudtaCttSV+
beBXvYANK1AhbsETnHTCyWvu4svOZSOedTYAVldVp6KueNG1OxRJF82L0gSmW2zi
DeU7UVlf1jfTCVqAVEP8BOcjxM3m9D5loHEBsic/lL9z2FkDUkUL2s676i3fJ6wJ
1Y+qKlkUwGv55BdaOYXPNXmIrwvahXZCdEoSjj/oLcEeHC2qD1Hh/I+vWxq129Ld
rOkzRp30bpoM691A6wPPb2SMLWYzF0dJv+uJgHqEAFozCS2fSYegRsZVofn0DCkS
Asx8l/F5t9jB/rs0m1SpCerXqrGq3hg/E8QppAVxt5MOGdBuZSBYRzrfK8APlp6b
aTVSi8K4+iTXyUlDXNRxGvAmfIbpXtvAUm6w+d+bOur4Re9SidRNx6O+V8c3LIJs
Tiksp7ubD0QsGUw7WBZ2qqMewipswXesh32ZjUKUWht6ckRF+pqJvXcKccqKJT4i
1NqGhkExzxZ869qsIN10HbORTGLBKOax8hKv1Pgxha+bEB0VgATLgSs7WeNznv0r
KrbtRPfHDVG/d++bjUEFXPs5R1a/bjiXfxJwqQehB1+EmKHRmf1Ca9L5SepPTaNI
JXCmLJiILQ65uvvW255Bmcp1RI+8PMrkq1V8QtbHjJhM8uFdBLYgEWCixjhRk31B
4h9lqehQLSW+zLPdBADw5PNwUfVqwG5Rbx/mGa53WAeOefCg1rIN4+ZpoavSvFn1
2xsBbOYnAZ8fLIViFskN6lUEFP+9JO0ZszxEe1YtioMe18CP3/kAmFiJHURB3CPw
be7NWA35fwdUsINqCD3m8AH6mDZlKbwgvmjqHN01dwLel90XEsHbsRyTuqZ4CASC
1gc0Fnosxs64NQp24t8XbnLJ8a4PGIKwKw+Bo3mAmkwYci599k43HJ3g+amxfeAd
DqXtqNlaRzhc7AwfJUIqyPVDk8DyK9yuiXK2zoxYVREbgQrjnEZyM/SYpEY/jPxE
EbjxzpseYN7D5vHt4lEQ+tYUtu/tvf/5ExIfvU3EzQpUYYrY/kb30jzzkr9wbT4i
EZXzfMXKQ1CDWamdeB8nDIbqfyQrIYveX4z8R0MWF9Zu4I9fuWmDanFS7bf/d8AH
t263WyUBJ7E2vZhB04gX/Jc92CNO0kgBDigex2aITJOzmQ5IApckfyJ3MEqpMM4q
Jfp0yuVS2xhiYwU075YV1GndcJkUsPHJ1VEmX9AT+fWQblxs6zuCkvWmDvH1M1Q0
Ah5udSiiq99XZUZPshG4GO2B1j+X2TKc5Trabbt81rzKWmuOkk4Rk5hU66q2ggHF
jI2FzuGpRz7asPFrXLIK0lTEqUwHXmw+x61tX5xx1BQsAivMq7sOT6jVLjHcMC/t
rx9YLNKQA4bDTY/2lSOAJAMILhyCBZBUJgcQQHudBQxL0ATTxof0jDxpNuSBtqfM
0dmz7MukGFSAMOQYbMtGULOtivlKCMB9s3d0jg2kCMnDiT4qTmdx+f1zhiV5yHoH
pambVdYDPbVYJ7xHGP6nnMqAAubQobABzc+jNjp/aSmn/gUKfgdMcbKax5YlkHlO
KQp9ZiZJESyiX9u60p/yGIRM/drLYizWiHDXEHbHwo9HMWyrRiorf0FthIH5eAgE
1mvmpGwzAJmpC+lxEsKgQBV+5HL2+++sozrhDeWWCSWngS9GoFhGE6+/exjuiH+I
LAWqzpjIe20lrgFJ+oWjXMo59xAzqnK0JC/fNTdQ2WClLQABS4pGQXffc7occ3f/
EgZHYqnoBnrCCqX8yI6mUqZsjoNXCast7pPWo46mrPyTKgyd93r5yTwAO+mmOje6
VXYcGIVNb2cEK7/ZJroBLylnXXM8Nj5i9mr6TMkEBXeMzLmS7ZuMFo2oZqFrH+RR
pK4iT3hEjUL0zfmqpoU95LBTmsbU8khMqKKEuP0mdsO1z56iNxUv3WzM0wKQE6je
t5K/9no45HYBUT7r0qQxg6hLRYBMyety5AP59g9pRy80gwph1R5fVK4F6REgE3fT
LBJ8R87VjiYx87buwtLNxVHJX86niRFIU1KiaeMbfRO4J5yPwp1yPDEw6FbtTgL0
1JaXlg0KJSRqYj/I8x18ch33tFwP7iE8KqzCNQW172v9G4KqCsdA0kKFZH0H2OY2
1zg7oB5hN/Mpa5H+NjOqo5p1evyELomJb1mobJ+o7+GXn7I4+DfG6c4Od6h4RM5V
EZ0dNFBKvyOx4BYXYhJrhfLHCraUXInwJhb0naxv6L6pXv34fa31GpDWsGKYZ99L
bcqyWRsmQ5+N094L5lOlm/7xbcBKn516xYd28Bjc+ThDdQi1G1oOaC5CZ3Z/6HGj
T/9XoZ58wzWADWJP/id6UhGI3EEtfPsgz4fLUFvELDEIlpqiaJn5lYcURm2f8yoH
CS+CuINu+EHBrk49yY7Ha8gt4TzoPgJp2pgDtH0sdMDYIz35x6wmioyMQdyLLIm2
tDUVAW3To/VdlO1H8FzqclydX5bN8OWTCjoeRKYSahgCcMfETV/UsOP4LtMgad32
dZbWqIIF0f7zmmiEXi+5yHGViGLPhclMAQuUTBcfDk5NubUwPwLKZp39KTag4DFr
BnsT2eAJw6JW+KSJoAgPovc0SfeVuI/jTE3f7s1PK+npwejJuZlbOJLV3aUx0YKR
lJMffrnqbgxxIZ93xLRJqU/EzN11OlM3KhCdhXMsQuOsG4z06QkNWWulg/0nKz3n
WfEDpU+D0L0el9ArpqsxcxVQIfNzW8Q1wMQeB6gD4CW/jnUTOsZfYpuWfUp3plHb
CH+S8n46VkCa07PpLUMEcwN7osfY9awpf6eQjWZI1bOrMVnYFwqUXcOvBhS0E6xL
+/YZsS7tM8s9sTJv7qf6V2HSm2WhfBrvwfdmZvcUmWqhMZUeMcskmMjrTtVgYbHf
un2jAmYsUD5YXw7Vd8Qb3ceD/aaOv0QPwz91o8XPIymEsfOwCow1ju22BS9dwZO7
2SV0uyxA+g8h5UBi379fDFkUqCaw8c9BMhiTyqgrsWvwCoX08J98U96bB5/K3MYX
k4DXs7RoZdOUPZ+x8Qsy4rIui8GXNTK/bj1TFx2VUeFM4YfzkiuEDbY98SG/fnfg
7kXfMSZkC1FmiyZM9+DyLdOPLTcKl17uHa0RdcH85YcrlP9jdjduRc0+a3/3lCRF
fKVr/kaWA4pDgKy51xbqCYda0P3rz7RTWFhA7oLuDkmO6cRifvm9MRmcxX93SiQg
7TE0kV5Tw0ILacD3paEZ0Zfj01AWcH4NKZj2J/iQ3qPFGNNFJNu1QBYhD04RFaZf
7yq9U+7i31Ledf0NPPBYK3okbryyWdLUyMqk404EBz/cHgBxHswvt2082WwFNgjz
VAJH+Ft22KYELfA4JoHR5oip1FY0j3luRr+WxwpvIhr9Tiofgk7tHI2VxG3rncdr
M+3jICPim2cisbrj17islCV9Zy3bLacb2dHSflYrjp8AzzgTh7+EP+SoTzmpPc0K
tgoec210k2YT5NBaQMfu7Sg6ZBdc/1rVdXgjTYxITZKQAtierU9BvCM9ee1MO03l
D2b/s14lFTIhmZPVlc2pp3Hh72V5I+ozUoOYbeikrAMwM8P6QMV6pjan7nxGcnxh
wRTkdDvv1XrER7bo+BOAkUWVs6WER8iRuZXrhk1PwnDVm2TgDuFJHwOgah35+a7F
8qwUwfVxJoTH+Qv2SwT2UKPCJOLgaPfpHyD814LHgFKopijXqx5IzyQPnS6B1YTY
LBbHiQY9rYWLBVUXSCQUvyloHbrnoVii9nGdSjYjKxWW1uQ03iUcqYi7spgRHjCS
MJv5Hs8e2LdVYpDM9y4xWSy4SQSg/U71akdNEgzBzG1M1DMp4Jz86XlmZnac/wgs
97L0h+0G3boMpXqrJ4Kb0y0h2oR6dvTDXF8z2sxkjCpvmgsd30Pfb/F1Eoc0F2e+
94/zKVRvcTBSfoNDCN3B+ws2kQ3BjOtEBnPnOrqByTB3OYu5kOwBBCWT8RV7VXdP
B4aMc3od5DBOdJMGVvhh+8o7DLbM4cXZRbiMlSpcXOzuk2f0Zuo4i/9t4M1Br55M
6QfGkck4+A7yDyW81h2vH+BwOW6iWth+YhR5nuM/MCM4t7Rkp0OLNtSmk2Mw4vI0
GLdtb2J1VTlqQlsR75k9Qn3fhrwcTN/6fUu7QW8CH1Fl6cmBkR5xzV7Rp4t923mu
RQHtGIr7Ki7h26pP5zf7DIdUzWHd8JwZOV7T2TAd/4X8KIsv80lw9p9un3lpkolQ
O+QV2d8jzQNhp9M+TfVoAp87ufUDlqx+l8GkK9H0NpP91xfC1kweRnUIHJrnIGEF
pv07MTxdBmUrbUUm1WQjA0qZup/Kzrwmti/kEIz70SD+N7gemq1L6Ybiqs6oPstm
BUt4eLAmkHZAbGPTM/Bs7cosIbYTHZ6K6GKMfG4nv1X0E2sHntmQqRKq+QeluD9m
xcaG8Priy/hUVAXFCRYdIncRvbY2epv9l2ItORChRxAp/I34L6SoLKULxy7HIevy
nwRztgE55rdqwbZEcG930tBVkex6TwV6IaVvKfFytqxLF8Zb9+4nkihZDnW/ouO7
dVF7Uo7IBEw2PkqpUMLpXsa2tuKy+ZbF6ideJNQZcoO6uy6FeCp+VXAEEu7oYZx5
ZXuut0dIPKjUQUNxNo0R4jaL/MvKUVnPG6vNiaVcW/s5PvxSBYyVrarKhD3eMh1t
jg1J9XtrBrndHXmaXAse0l2klZV1f8s1M8iY6gViX7WBhpVsV+TCCqMNlpifBvr9
1Ou2V9PzTo51dbAf7gXut1oacV+EM0vVhCNMm5kWFkSLyZrYmZRVaQ7bvAevXT1q
0jJ9yCS1k8xBT3hZziyQaEWDa/kmemU6KbnWQR8Uq/5Q27y/u+lrOwQJXZSN1b7+
3IrH05+5OYXqdWEpFimJc8AsOZuUfZ3iB+uJf3iljmpD0RzgDLOOk9hvH4E2lUrp
YHHVd3vpnTdLV5btvPtVdpX4BNtCXbxpeaduRwv/ahR1EBRZzDa7cG+zPHiWKvMv
s2+vimcYRv3wEdJ7w2nKWh/2fVoqSrVlIjS+RV7e8v3epBiySxvHyvMpcGzYBSSX
i9/MDD4U+A/17wJdAfqtu11gmtTTi/K6UBkv202V2VIz2h6+E3dtDftzI4VAZbsM
u6OebDvETrIHGodeRryOW7Dztoa4129KyuK+odKXLtp4MUDvLlChRI1mDBzxP8VK
guMSmqQLL3XS0mynkEJvRyy9vAQdK2RzRweU3mPgF0gTg1a+4R3I8ZmIsJB16k9I
Bfd9TahcumAwlsype0D1ppCkTyAEh9jYtp7aO82uTH+LVlx33aPj/Sg+WeAxJSb6
VPBPZzVvBs50uAchV4hTviiAKbBDyyvw0JYgnszSjJDf8smtcUuwkJF92c44aQHS
SNgCvoNgfPsJEqDDA/9FpmZUWVIFqbqR33xQt2jeyNg/EKXaps93z/8TEKmXhmQh
jP3VOBnIrM4zyJ11trUnObybaiYgoUJvh+mIlUWokzXxCvl3qpj1JrllH5h+xF8Z
7PnZSYQNx3yLisN0DK3b1RFmm1OTqPWJ1RaM85LSZ3jdmr9BFXW4Q/EBvvT7SA9k
N17Oob6AYhRNrGi47JQbS77VgI6o/7ehkKm1Y+lQfJIuYY3ikVdYgsbnhaQYdVA7
ouQHaAuMClUeI1IABWlhgvIaZHytuSM+sUkBHOFNf8mwOVUC9yli6sfibBxDHKt9
2GqFVA8HM0Lnr+EFtDudWwWJyNXskOSfkeFdHZ8piWxgi+rG9FiT/aR/CWRDmAHc
LXsUSSldiBmjXi7EYLSPgxjaVCrLmG562en9VcLPcwjBJe7cna7qHsp7hiO9SQEH
eq6hmNa8MrWtkdRJzrzuhlQlkndM9YUMwcilakdqOSkUqFS8PtZu0APy3t1+d54b
/9VcLrTkYGPJ1HCCIZ1RUYmDq7hqfLf2du/jz8oR6KToJoA38PHIozmNxY7L+zvc
Oi02kkF7Fri7d4NevOo/N5zOWXwxg781cID9224Z/p7XFtpiW1KeDFqJI2wfPx+e
6TegQxuas2LwCXN6Hp7IhzcDfiD/iD5/5eSFNlYNJq9QLZmQ+BTxVPyg5eu6D9An
BkOWFpPouUzep5hyd73B2zfTOP+HKXgAI1Hh95NVNY+daZ3a8Hd3SzV8Lyxvy6lz
QPog0+RsN8ScFWiGaowWICa6ClidzkKiDA7JQLT5h0ODKSJwNWRouvGrDSB7nMMd
F8faTW8Ps/g7cLa7I/9dO8efcfv2+VAEtJRp2+g12RRTDoMUhzbKikrAKRnQTGv8
ePBtwTudM1cBq52380XiQDBHkDji3RWIxCyqDR6iAZAhuqpLk7TAHTTae2885k1+
eL1jo6YSnEDjcrcfItJZaPrUcoyiRm5uFzDxeZJv2QX8S79tVP/RyQOiR3WreeJm
J1mTI3JvD64Ga3vibOtykPr434NDNI2u0W/k0LMr/WsxT5YU6REVLBZHmbsVKmpl
6fiik35mkCXJZcNj0TtY+8PqmkDNFUDfVV0hVGkOB0dm31p74BpEwXDoJljebJOd
eQutQhIknMlSrwQo65aKiGRi7evV38Yj0xVsZ+2WpHf8J/2I04xAB9wXROnp2A1r
flIdfcUNLHpgwPEJPHTRZbn9JhJIv3GJURKlwe2u09sHdeC+b6tIDwmq0YgsvWPP
H2YU8HS8/Q5I+6n5u7Ak+0D6KCAsqWH/nc8/XDjMpZy3X/ZWmD2LzI2hmvhzgckC
+WHBVL0F4HzBCmBtncy3mILZsKscVJm1iG51Qst0iI7HgUB405OobJsDosLHsJvN
Fw363wnpmGoQuVeWLB5qXXTEf27Bq/nhb79vF7XPtzzLLdeiU/Dg+GkF7JJ83G45
jgeYUXHOPE2uQpXFsRbp/uzjYcnb5wf+PrSVO6S/98mQxsqNzbhFgxHMStwMOGil
awU7ZgdJfNBrK0u4YcHCBLVXoXZXJ5oh0iHO806/tfRqBsMkLPgeRRqjnQNLxQoT
9shJiOVDV6MQcuJNS4Dz+IDPdrss1dlGoLdpTDKJILzXJQnwwTSc/nDSmSeM34Ra
EUiNvut/OKC0FYjkuPj1WPdz1a1SAeSbYzVvHRRf5nnXmrzHg0VCjHXXouHp3LWc
QTCkKi/MzBZCRCz8W3QsCkOhbZMFRel5zI546cp8rvIUBqxN1WPuoe1cpouvraJZ
UBssyFVIzXCtj6UtiF+6g3+biKaIobLRytIXKoKh50yx2gc130jtiYc81LDGEm9O
HDD8B7cFFBYK/i5jTQsun4JNuy3acKk7IlzXs3dGV/YRMJz1GKInrgi2TXDOnGwm
YUpPZ6FTbpP2jPTuh8g8cE7hI5nh/Y1W24RbZQphGV+QvVZQryzkkGHeoMTk2oZ8
2/kqffJyeQy0HMvkOgVcG7BD+z6jD+UHCVn8Sv3j9DGgakS2b+x2FKNI9nyaLNM4
mMnJtcNgLez21xm6QtDrr/0tW/PeXBpjL+8W9Jg0s0x8B15QTjxLVpYeiBoNs0IH
WteVfKO2Ym5UlNGOakAgr5AvLus8MRy/GE6ReTOhSeogJLwQBfzud+1f97Eeq3Ws
YYNAlcVRRv6SEtWE+7Dz9jESycYu/k1Ds1ROLcie7dmZY6YS2X4fXkIQe0+Mje/w
WOfuXRytz7ggMouKMby+uWu+Le92sGCUmXMHrUSV4osytK0GMTCyVBBPdPT9owx+
GHMBFbimDHncdCd/hAhE8j6Wq1/bXgpI5cuzLwcuTt3LoXJ/znTwnzTVipfViyy8
Ic8MnkD2x+ULYpg9WSl/wYmfxDjm0qLwWpR9iTBpgo9zlGxp7/c+vMjz92R4RJDU
dksDEJ1iVR/t17oTXdrrVRjEBgbqZHasAWvQnrMeszK1Wj9bCb8EcNF8oaEsKVKK
+AjAnSSt8qvrhbaTye58OYZaejKoaRuGjEGnhuwVoM99NaNttyh90ENK53agXhv3
R8RLA7gf6xXYZbTIhUtg+uEH/CfO+l/5aWFoLlfNtiB72gpCANO0YrhFTxXOooxe
CQgIQEdJT4OiLpDEHQyTWYEa0fViSuHgmZu0S2W1vBSr44irQ5hyOP+AjticOxIN
vBCDvllZb0oke8aUApZbVkTxKPoUm5SBDWnOZYQx4frQW0ZyQXMD+67aTfQrYuTO
rfJp7+phEcwkRJoEB+Fa66mh6imyLC0ZK69NWgJEj+8r3xdoJS6ALq8RD1L2QggE
2dL5ps6zYcFVmjVbjBoLyQIKD/U+7KpmKbVP+6ih9na0F5YdfVr71EAlvKKw9jJQ
Hi8BsORFs5Rl9bXeTQFWgu9+roAbB66X7O/GiC+hBDbqUsIhdTrB3aiWRQjwI5kI
03h2BA8HIKq/jPA38Yd8VkZuSn3h92pOZtP1rQH4mc7S7LTrL6YDpdnL73tdA/rK
S4NVWLWOTU3jExF4zG5H5KKRS5uQ1lkJR2xSG3slyYfOJeFdYk9nwBWqjALbeVjz
D52bccdqXVppRr/OKp1F5CNCNy8xnU9gpaUzANDsFo4IAWMSd+gJ/UogSoczaqA7
JVe1WJSIU9gJqP6lla+TtplOY5UKb7EUPte6Nh5dTESYN+8PweWPOnY7V5GZGHoH
M1xjCq2uo8nRGh68etHIrw==
`pragma protect end_protected
