// megafunction wizard: %Stratix V Hard IP for PCI Express v14.0%
// GENERATION: XML
// pcie3.v

// Generated using ACDS version 14.0 205 at 2014.09.25.03:51:45

`timescale 1 ps / 1 ps
module pcie3 
#(
        parameter FORCE_GEN2,
        parameter VENDOR_ID,
        parameter DEVICE_ID,
        parameter INCREASE_DRIVE_STRENGTH,
        parameter DEBUG_WIDTH
)
(
		input  wire         npor,               //               npor.npor
		input  wire         pin_perst,          //                   .pin_perst
		input  wire [11:0]  lmi_addr,           //                lmi.lmi_addr
		input  wire [31:0]  lmi_din,            //                   .lmi_din
		input  wire         lmi_rden,           //                   .lmi_rden
		input  wire         lmi_wren,           //                   .lmi_wren
		output wire         lmi_ack,            //                   .lmi_ack
		output wire [31:0]  lmi_dout,           //                   .lmi_dout
		input  wire [4:0]   hpg_ctrler,         //          config_tl.hpg_ctrler
		output wire [3:0]   tl_cfg_add,         //                   .tl_cfg_add
		output wire [31:0]  tl_cfg_ctl,         //                   .tl_cfg_ctl
		output wire [52:0]  tl_cfg_sts,         //                   .tl_cfg_sts
		input  wire [6:0]   cpl_err,            //                   .cpl_err
		input  wire         cpl_pending,        //                   .cpl_pending
		input  wire         pm_auxpwr,          //         power_mngt.pm_auxpwr
		input  wire [9:0]   pm_data,            //                   .pm_data
		input  wire         pme_to_cr,          //                   .pme_to_cr
		input  wire         pm_event,           //                   .pm_event
		output wire         pme_to_sr,          //                   .pme_to_sr
		output wire [0:0]   rx_st_sop,          //              rx_st.startofpacket
		output wire [0:0]   rx_st_eop,          //                   .endofpacket
		output wire [0:0]   rx_st_err,          //                   .error
		output wire [0:0]   rx_st_valid,        //                   .valid
		output wire [1:0]   rx_st_empty,        //                   .empty
		input  wire         rx_st_ready,        //                   .ready
		output wire [255:0] rx_st_data,         //                   .data
		output wire [7:0]   rx_st_bar,          //          rx_bar_be.rx_st_bar
		input  wire         rx_st_mask,         //                   .rx_st_mask
		input  wire [0:0]   tx_st_sop,          //              tx_st.startofpacket
		input  wire [0:0]   tx_st_eop,          //                   .endofpacket
		input  wire [0:0]   tx_st_err,          //                   .error
		input  wire [0:0]   tx_st_valid,        //                   .valid
		input  wire [1:0]   tx_st_empty,        //                   .empty
		output wire         tx_st_ready,        //                   .ready
		input  wire [255:0] tx_st_data,         //                   .data
		output wire [11:0]  tx_cred_datafccp,   //            tx_cred.tx_cred_datafccp
		output wire [11:0]  tx_cred_datafcnp,   //                   .tx_cred_datafcnp
		output wire [11:0]  tx_cred_datafcp,    //                   .tx_cred_datafcp
		output wire [5:0]   tx_cred_fchipcons,  //                   .tx_cred_fchipcons
		output wire [5:0]   tx_cred_fcinfinite, //                   .tx_cred_fcinfinite
		output wire [7:0]   tx_cred_hdrfccp,    //                   .tx_cred_hdrfccp
		output wire [7:0]   tx_cred_hdrfcnp,    //                   .tx_cred_hdrfcnp
		output wire [7:0]   tx_cred_hdrfcp,     //                   .tx_cred_hdrfcp
		input  wire         pld_clk,            //            pld_clk.clk
		output wire         coreclkout_hip,     //     coreclkout_hip.clk
		input  wire         refclk,             //             refclk.clk
		output wire         reset_status,       //            hip_rst.reset_status
		output wire         serdes_pll_locked,  //                   .serdes_pll_locked
		output wire         pld_clk_inuse,      //                   .pld_clk_inuse
		input  wire         pld_core_ready,     //                   .pld_core_ready
		output wire         testin_zero,        //                   .testin_zero
		input  wire [769:0] reconfig_to_xcvr,   //   reconfig_to_xcvr.reconfig_to_xcvr
		output wire [505:0] reconfig_from_xcvr, // reconfig_from_xcvr.reconfig_from_xcvr
		input  wire         rx_in0,             //         hip_serial.rx_in0
		input  wire         rx_in1,             //                   .rx_in1
		input  wire         rx_in2,             //                   .rx_in2
		input  wire         rx_in3,             //                   .rx_in3
		input  wire         rx_in4,             //                   .rx_in4
		input  wire         rx_in5,             //                   .rx_in5
		input  wire         rx_in6,             //                   .rx_in6
		input  wire         rx_in7,             //                   .rx_in7
		output wire         tx_out0,            //                   .tx_out0
		output wire         tx_out1,            //                   .tx_out1
		output wire         tx_out2,            //                   .tx_out2
		output wire         tx_out3,            //                   .tx_out3
		output wire         tx_out4,            //                   .tx_out4
		output wire         tx_out5,            //                   .tx_out5
		output wire         tx_out6,            //                   .tx_out6
		output wire         tx_out7,            //                   .tx_out7
		input  wire         sim_pipe_pclk_in,   //           hip_pipe.sim_pipe_pclk_in
		output wire [1:0]   sim_pipe_rate,      //                   .sim_pipe_rate
		output wire [4:0]   sim_ltssmstate,     //                   .sim_ltssmstate
		output wire [2:0]   eidleinfersel0,     //                   .eidleinfersel0
		output wire [2:0]   eidleinfersel1,     //                   .eidleinfersel1
		output wire [2:0]   eidleinfersel2,     //                   .eidleinfersel2
		output wire [2:0]   eidleinfersel3,     //                   .eidleinfersel3
		output wire [2:0]   eidleinfersel4,     //                   .eidleinfersel4
		output wire [2:0]   eidleinfersel5,     //                   .eidleinfersel5
		output wire [2:0]   eidleinfersel6,     //                   .eidleinfersel6
		output wire [2:0]   eidleinfersel7,     //                   .eidleinfersel7
		output wire [1:0]   powerdown0,         //                   .powerdown0
		output wire [1:0]   powerdown1,         //                   .powerdown1
		output wire [1:0]   powerdown2,         //                   .powerdown2
		output wire [1:0]   powerdown3,         //                   .powerdown3
		output wire [1:0]   powerdown4,         //                   .powerdown4
		output wire [1:0]   powerdown5,         //                   .powerdown5
		output wire [1:0]   powerdown6,         //                   .powerdown6
		output wire [1:0]   powerdown7,         //                   .powerdown7
		output wire         rxpolarity0,        //                   .rxpolarity0
		output wire         rxpolarity1,        //                   .rxpolarity1
		output wire         rxpolarity2,        //                   .rxpolarity2
		output wire         rxpolarity3,        //                   .rxpolarity3
		output wire         rxpolarity4,        //                   .rxpolarity4
		output wire         rxpolarity5,        //                   .rxpolarity5
		output wire         rxpolarity6,        //                   .rxpolarity6
		output wire         rxpolarity7,        //                   .rxpolarity7
		output wire         txcompl0,           //                   .txcompl0
		output wire         txcompl1,           //                   .txcompl1
		output wire         txcompl2,           //                   .txcompl2
		output wire         txcompl3,           //                   .txcompl3
		output wire         txcompl4,           //                   .txcompl4
		output wire         txcompl5,           //                   .txcompl5
		output wire         txcompl6,           //                   .txcompl6
		output wire         txcompl7,           //                   .txcompl7
		output wire [7:0]   txdata0,            //                   .txdata0
		output wire [7:0]   txdata1,            //                   .txdata1
		output wire [7:0]   txdata2,            //                   .txdata2
		output wire [7:0]   txdata3,            //                   .txdata3
		output wire [7:0]   txdata4,            //                   .txdata4
		output wire [7:0]   txdata5,            //                   .txdata5
		output wire [7:0]   txdata6,            //                   .txdata6
		output wire [7:0]   txdata7,            //                   .txdata7
		output wire         txdatak0,           //                   .txdatak0
		output wire         txdatak1,           //                   .txdatak1
		output wire         txdatak2,           //                   .txdatak2
		output wire         txdatak3,           //                   .txdatak3
		output wire         txdatak4,           //                   .txdatak4
		output wire         txdatak5,           //                   .txdatak5
		output wire         txdatak6,           //                   .txdatak6
		output wire         txdatak7,           //                   .txdatak7
		output wire         txdetectrx0,        //                   .txdetectrx0
		output wire         txdetectrx1,        //                   .txdetectrx1
		output wire         txdetectrx2,        //                   .txdetectrx2
		output wire         txdetectrx3,        //                   .txdetectrx3
		output wire         txdetectrx4,        //                   .txdetectrx4
		output wire         txdetectrx5,        //                   .txdetectrx5
		output wire         txdetectrx6,        //                   .txdetectrx6
		output wire         txdetectrx7,        //                   .txdetectrx7
		output wire         txelecidle0,        //                   .txelecidle0
		output wire         txelecidle1,        //                   .txelecidle1
		output wire         txelecidle2,        //                   .txelecidle2
		output wire         txelecidle3,        //                   .txelecidle3
		output wire         txelecidle4,        //                   .txelecidle4
		output wire         txelecidle5,        //                   .txelecidle5
		output wire         txelecidle6,        //                   .txelecidle6
		output wire         txelecidle7,        //                   .txelecidle7
		output wire         txdeemph0,          //                   .txdeemph0
		output wire         txdeemph1,          //                   .txdeemph1
		output wire         txdeemph2,          //                   .txdeemph2
		output wire         txdeemph3,          //                   .txdeemph3
		output wire         txdeemph4,          //                   .txdeemph4
		output wire         txdeemph5,          //                   .txdeemph5
		output wire         txdeemph6,          //                   .txdeemph6
		output wire         txdeemph7,          //                   .txdeemph7
		output wire [2:0]   txmargin0,          //                   .txmargin0
		output wire [2:0]   txmargin1,          //                   .txmargin1
		output wire [2:0]   txmargin2,          //                   .txmargin2
		output wire [2:0]   txmargin3,          //                   .txmargin3
		output wire [2:0]   txmargin4,          //                   .txmargin4
		output wire [2:0]   txmargin5,          //                   .txmargin5
		output wire [2:0]   txmargin6,          //                   .txmargin6
		output wire [2:0]   txmargin7,          //                   .txmargin7
		output wire         txswing0,           //                   .txswing0
		output wire         txswing1,           //                   .txswing1
		output wire         txswing2,           //                   .txswing2
		output wire         txswing3,           //                   .txswing3
		output wire         txswing4,           //                   .txswing4
		output wire         txswing5,           //                   .txswing5
		output wire         txswing6,           //                   .txswing6
		output wire         txswing7,           //                   .txswing7
		input  wire         phystatus0,         //                   .phystatus0
		input  wire         phystatus1,         //                   .phystatus1
		input  wire         phystatus2,         //                   .phystatus2
		input  wire         phystatus3,         //                   .phystatus3
		input  wire         phystatus4,         //                   .phystatus4
		input  wire         phystatus5,         //                   .phystatus5
		input  wire         phystatus6,         //                   .phystatus6
		input  wire         phystatus7,         //                   .phystatus7
		input  wire [7:0]   rxdata0,            //                   .rxdata0
		input  wire [7:0]   rxdata1,            //                   .rxdata1
		input  wire [7:0]   rxdata2,            //                   .rxdata2
		input  wire [7:0]   rxdata3,            //                   .rxdata3
		input  wire [7:0]   rxdata4,            //                   .rxdata4
		input  wire [7:0]   rxdata5,            //                   .rxdata5
		input  wire [7:0]   rxdata6,            //                   .rxdata6
		input  wire [7:0]   rxdata7,            //                   .rxdata7
		input  wire         rxdatak0,           //                   .rxdatak0
		input  wire         rxdatak1,           //                   .rxdatak1
		input  wire         rxdatak2,           //                   .rxdatak2
		input  wire         rxdatak3,           //                   .rxdatak3
		input  wire         rxdatak4,           //                   .rxdatak4
		input  wire         rxdatak5,           //                   .rxdatak5
		input  wire         rxdatak6,           //                   .rxdatak6
		input  wire         rxdatak7,           //                   .rxdatak7
		input  wire         rxelecidle0,        //                   .rxelecidle0
		input  wire         rxelecidle1,        //                   .rxelecidle1
		input  wire         rxelecidle2,        //                   .rxelecidle2
		input  wire         rxelecidle3,        //                   .rxelecidle3
		input  wire         rxelecidle4,        //                   .rxelecidle4
		input  wire         rxelecidle5,        //                   .rxelecidle5
		input  wire         rxelecidle6,        //                   .rxelecidle6
		input  wire         rxelecidle7,        //                   .rxelecidle7
		input  wire [2:0]   rxstatus0,          //                   .rxstatus0
		input  wire [2:0]   rxstatus1,          //                   .rxstatus1
		input  wire [2:0]   rxstatus2,          //                   .rxstatus2
		input  wire [2:0]   rxstatus3,          //                   .rxstatus3
		input  wire [2:0]   rxstatus4,          //                   .rxstatus4
		input  wire [2:0]   rxstatus5,          //                   .rxstatus5
		input  wire [2:0]   rxstatus6,          //                   .rxstatus6
		input  wire [2:0]   rxstatus7,          //                   .rxstatus7
		input  wire         rxvalid0,           //                   .rxvalid0
		input  wire         rxvalid1,           //                   .rxvalid1
		input  wire         rxvalid2,           //                   .rxvalid2
		input  wire         rxvalid3,           //                   .rxvalid3
		input  wire         rxvalid4,           //                   .rxvalid4
		input  wire         rxvalid5,           //                   .rxvalid5
		input  wire         rxvalid6,           //                   .rxvalid6
		input  wire         rxvalid7,           //                   .rxvalid7
		input  wire         app_int_sts,        //            int_msi.app_int_sts
		input  wire [4:0]   app_msi_num,        //                   .app_msi_num
		input  wire         app_msi_req,        //                   .app_msi_req
		input  wire [2:0]   app_msi_tc,         //                   .app_msi_tc
		output wire         app_int_ack,        //                   .app_int_ack
		output wire         app_msi_ack,        //                   .app_msi_ack
		input  wire [31:0]  test_in,            //           hip_ctrl.test_in
		input  wire         simu_mode_pipe,     //                   .simu_mode_pipe
		output wire         derr_cor_ext_rcv,   //         hip_status.derr_cor_ext_rcv
		output wire         derr_cor_ext_rpl,   //                   .derr_cor_ext_rpl
		output wire         derr_rpl,           //                   .derr_rpl
		output wire         dlup,               //                   .dlup
		output wire         dlup_exit,          //                   .dlup_exit
		output wire         ev128ns,            //                   .ev128ns
		output wire         ev1us,              //                   .ev1us
		output wire         hotrst_exit,        //                   .hotrst_exit
		output wire [3:0]   int_status,         //                   .int_status
		output wire         l2_exit,            //                   .l2_exit
		output wire [3:0]   lane_act,           //                   .lane_act
		output wire [4:0]   ltssmstate,         //                   .ltssmstate
		output wire         rx_par_err,         //                   .rx_par_err
		output wire [1:0]   tx_par_err,         //                   .tx_par_err
		output wire         cfg_par_err,        //                   .cfg_par_err
		output wire [7:0]   ko_cpl_spc_header,  //                   .ko_cpl_spc_header
		output wire [11:0]  ko_cpl_spc_data,    //                   .ko_cpl_spc_data
		output wire [1:0]   currentspeed,       //   hip_currentspeed.currentspeed
		output wire [DEBUG_WIDTH-1:0]   debug
	);

	altpcie_sv_hip_ast_hwtcl #(
        .DEBUG_WIDTH                              (DEBUG_WIDTH),
		.ACDS_VERSION_HWTCL                       ("14.0"),
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              (FORCE_GEN2 == 1 ? "Gen2 (5.0 Gbps)" : "Gen3 (8.0 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("3.0"),
		.ast_width_hwtcl                          ("Avalon-ST 256-bit"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.use_ast_parity                           (0),
		.multiple_packets_per_cycle_hwtcl         (0),
		.in_cvp_mode_hwtcl                        (0),
		.use_pci_ext_hwtcl                        (0),
		.use_pcie_ext_hwtcl                       (0),
		.use_config_bypass_hwtcl                  (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.hip_reconfig_hwtcl                       (0),
		.hip_tag_checking_hwtcl                   (1),
		.enable_power_on_rst_pulse_hwtcl          (1),
		.enable_pcisigtest_hwtcl                  (0),
		.bar0_size_mask_hwtcl                     (24),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Disabled"),
		.bar0_prefetchable_hwtcl                  ("Disabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (0),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.expansion_base_address_register_hwtcl    (0),
		.io_window_addr_width_hwtcl               (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.vendor_id_hwtcl                          (VENDOR_ID), //(4466),  // Microsoft
		.device_id_hwtcl                          (DEVICE_ID), //(57345), // HIP 0
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (16711680),
		.subsystem_vendor_id_hwtcl                (0),
		.subsystem_device_id_hwtcl                (0),
		.max_payload_size_hwtcl                   (256),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (1),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (40960),
		.user_id_hwtcl                            (0),
		.vsec_rev_hwtcl                           (0),
		.pcie_toolkit_enable_hwtcl                ("false"),
		.millisecond_cycle_count_hwtcl            (248500),
		.port_width_be_hwtcl                      (32),
		.port_width_data_hwtcl                    (256),
		.gen3_dcbal_en_hwtcl                      (1),
		.enable_pipe32_sim_hwtcl                  (0),
		.fixed_preset_on                          (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("true"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (770),
		.reconfig_from_xcvr_width                 (506),
		.single_rx_detect_hwtcl                   (0),
		.hip_hard_reset_hwtcl                     (0),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15),
		.hwtcl_override_g3rxcoef                  (0),   // Don't override because not all params here aren't the correct defaults
		.gen3_coeff_1_hwtcl                       ( (INCREASE_DRIVE_STRENGTH == 1) ? 9 : 7 ),   // 7 -- default, 9 -- increased drive
		.gen3_coeff_1_sel_hwtcl                   ("preset_1"),
		.gen3_coeff_1_preset_hint_hwtcl           (0),
		.gen3_coeff_1_nxtber_more_ptr_hwtcl       ( (INCREASE_DRIVE_STRENGTH == 1) ? 2 : 1 ),   // 1 -- default, 2 -- Selecting P4 regardless of BER 
		.gen3_coeff_1_nxtber_more_hwtcl           ("g3_coeff_1_nxtber_more"),
		.gen3_coeff_1_nxtber_less_ptr_hwtcl       (1),
		.gen3_coeff_1_nxtber_less_hwtcl           ("g3_coeff_1_nxtber_less"),
		.gen3_coeff_1_reqber_hwtcl                (0),
		.gen3_coeff_1_ber_meas_hwtcl              (2),
		.gen3_coeff_2_hwtcl                       (0),
		.gen3_coeff_2_sel_hwtcl                   ("preset_2"),
		.gen3_coeff_2_preset_hint_hwtcl           (0),
		.gen3_coeff_2_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_2_nxtber_more_hwtcl           ("g3_coeff_2_nxtber_more"),
		.gen3_coeff_2_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_2_nxtber_less_hwtcl           ("g3_coeff_2_nxtber_less"),
		.gen3_coeff_2_reqber_hwtcl                (0),
		.gen3_coeff_2_ber_meas_hwtcl              (0),
		.gen3_coeff_3_hwtcl                       ((INCREASE_DRIVE_STRENGTH == 1) ? 9 : 7), // 7 -- default, 9 -- AEQ Waiting state for 1st selected preset
		.gen3_coeff_3_sel_hwtcl                   ("preset_3"),
		.gen3_coeff_3_preset_hint_hwtcl           (0),
		.gen3_coeff_3_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_3_nxtber_more_hwtcl           ("g3_coeff_3_nxtber_more"),
		.gen3_coeff_3_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_3_nxtber_less_hwtcl           ("g3_coeff_3_nxtber_less"),
		.gen3_coeff_3_reqber_hwtcl                (0),
		.gen3_coeff_3_ber_meas_hwtcl              (0),
		.gen3_coeff_4_hwtcl                       (0),
		.gen3_coeff_4_sel_hwtcl                   ("preset_4"),
		.gen3_coeff_4_preset_hint_hwtcl           (0),
		.gen3_coeff_4_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_4_nxtber_more_hwtcl           ("g3_coeff_4_nxtber_more"),
		.gen3_coeff_4_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_4_nxtber_less_hwtcl           ("g3_coeff_4_nxtber_less"),
		.gen3_coeff_4_reqber_hwtcl                (0),
		.gen3_coeff_4_ber_meas_hwtcl              (0),
		.gen3_coeff_5_hwtcl                       (0),
		.gen3_coeff_5_sel_hwtcl                   ("preset_5"),
		.gen3_coeff_5_preset_hint_hwtcl           (0),
		.gen3_coeff_5_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_5_nxtber_more_hwtcl           ("g3_coeff_5_nxtber_more"),
		.gen3_coeff_5_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_5_nxtber_less_hwtcl           ("g3_coeff_5_nxtber_less"),
		.gen3_coeff_5_reqber_hwtcl                (0),
		.gen3_coeff_5_ber_meas_hwtcl              (0),
		.gen3_coeff_6_hwtcl                       (0),
		.gen3_coeff_6_sel_hwtcl                   ("preset_6"),
		.gen3_coeff_6_preset_hint_hwtcl           (0),
		.gen3_coeff_6_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_6_nxtber_more_hwtcl           ("g3_coeff_6_nxtber_more"),
		.gen3_coeff_6_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_6_nxtber_less_hwtcl           ("g3_coeff_6_nxtber_less"),
		.gen3_coeff_6_reqber_hwtcl                (0),
		.gen3_coeff_6_ber_meas_hwtcl              (0),
		.gen3_coeff_7_hwtcl                       (0),
		.gen3_coeff_7_sel_hwtcl                   ("preset_7"),
		.gen3_coeff_7_preset_hint_hwtcl           (0),
		.gen3_coeff_7_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_7_nxtber_more_hwtcl           ("g3_coeff_7_nxtber_more"),
		.gen3_coeff_7_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_7_nxtber_less_hwtcl           ("g3_coeff_7_nxtber_less"),
		.gen3_coeff_7_reqber_hwtcl                (0),
		.gen3_coeff_7_ber_meas_hwtcl              (0),
		.gen3_coeff_8_hwtcl                       (0),
		.gen3_coeff_8_sel_hwtcl                   ("preset_8"),
		.gen3_coeff_8_preset_hint_hwtcl           (0),
		.gen3_coeff_8_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_8_nxtber_more_hwtcl           ("g3_coeff_8_nxtber_more"),
		.gen3_coeff_8_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_8_nxtber_less_hwtcl           ("g3_coeff_8_nxtber_less"),
		.gen3_coeff_8_reqber_hwtcl                (0),
		.gen3_coeff_8_ber_meas_hwtcl              (0),
		.gen3_coeff_9_hwtcl                       (0),
		.gen3_coeff_9_sel_hwtcl                   ("preset_9"),
		.gen3_coeff_9_preset_hint_hwtcl           (0),
		.gen3_coeff_9_nxtber_more_ptr_hwtcl       (0),
		.gen3_coeff_9_nxtber_more_hwtcl           ("g3_coeff_9_nxtber_more"),
		.gen3_coeff_9_nxtber_less_ptr_hwtcl       (0),
		.gen3_coeff_9_nxtber_less_hwtcl           ("g3_coeff_9_nxtber_less"),
		.gen3_coeff_9_reqber_hwtcl                (0),
		.gen3_coeff_9_ber_meas_hwtcl              (0),
		.gen3_coeff_10_hwtcl                      (0),
		.gen3_coeff_10_sel_hwtcl                  ("preset_10"),
		.gen3_coeff_10_preset_hint_hwtcl          (0),
		.gen3_coeff_10_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_10_nxtber_more_hwtcl          ("g3_coeff_10_nxtber_more"),
		.gen3_coeff_10_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_10_nxtber_less_hwtcl          ("g3_coeff_10_nxtber_less"),
		.gen3_coeff_10_reqber_hwtcl               (0),
		.gen3_coeff_10_ber_meas_hwtcl             (0),
		.gen3_coeff_11_hwtcl                      (0),
		.gen3_coeff_11_sel_hwtcl                  ("preset_11"),
		.gen3_coeff_11_preset_hint_hwtcl          (0),
		.gen3_coeff_11_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_11_nxtber_more_hwtcl          ("g3_coeff_11_nxtber_more"),
		.gen3_coeff_11_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_11_nxtber_less_hwtcl          ("g3_coeff_11_nxtber_less"),
		.gen3_coeff_11_reqber_hwtcl               (0),
		.gen3_coeff_11_ber_meas_hwtcl             (0),
		.gen3_coeff_12_hwtcl                      (0),
		.gen3_coeff_12_sel_hwtcl                  ("preset_12"),
		.gen3_coeff_12_preset_hint_hwtcl          (0),
		.gen3_coeff_12_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_12_nxtber_more_hwtcl          ("g3_coeff_12_nxtber_more"),
		.gen3_coeff_12_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_12_nxtber_less_hwtcl          ("g3_coeff_12_nxtber_less"),
		.gen3_coeff_12_reqber_hwtcl               (0),
		.gen3_coeff_12_ber_meas_hwtcl             (0),
		.gen3_coeff_13_hwtcl                      (0),
		.gen3_coeff_13_sel_hwtcl                  ("preset_13"),
		.gen3_coeff_13_preset_hint_hwtcl          (0),
		.gen3_coeff_13_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_13_nxtber_more_hwtcl          ("g3_coeff_13_nxtber_more"),
		.gen3_coeff_13_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_13_nxtber_less_hwtcl          ("g3_coeff_13_nxtber_less"),
		.gen3_coeff_13_reqber_hwtcl               (0),
		.gen3_coeff_13_ber_meas_hwtcl             (0),
		.gen3_coeff_14_hwtcl                      (0),
		.gen3_coeff_14_sel_hwtcl                  ("preset_14"),
		.gen3_coeff_14_preset_hint_hwtcl          (0),
		.gen3_coeff_14_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_14_nxtber_more_hwtcl          ("g3_coeff_14_nxtber_more"),
		.gen3_coeff_14_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_14_nxtber_less_hwtcl          ("g3_coeff_14_nxtber_less"),
		.gen3_coeff_14_reqber_hwtcl               (0),
		.gen3_coeff_14_ber_meas_hwtcl             (0),
		.gen3_coeff_15_hwtcl                      (0),
		.gen3_coeff_15_sel_hwtcl                  ("preset_15"),
		.gen3_coeff_15_preset_hint_hwtcl          (0),
		.gen3_coeff_15_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_15_nxtber_more_hwtcl          ("g3_coeff_15_nxtber_more"),
		.gen3_coeff_15_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_15_nxtber_less_hwtcl          ("g3_coeff_15_nxtber_less"),
		.gen3_coeff_15_reqber_hwtcl               (0),
		.gen3_coeff_15_ber_meas_hwtcl             (0),
		.gen3_coeff_16_hwtcl                      (0),
		.gen3_coeff_16_sel_hwtcl                  ("preset_16"),
		.gen3_coeff_16_preset_hint_hwtcl          (0),
		.gen3_coeff_16_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_16_nxtber_more_hwtcl          ("g3_coeff_16_nxtber_more"),
		.gen3_coeff_16_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_16_nxtber_less_hwtcl          ("g3_coeff_16_nxtber_less"),
		.gen3_coeff_16_reqber_hwtcl               (0),
		.gen3_coeff_16_ber_meas_hwtcl             (0),
		.gen3_coeff_17_hwtcl                      (0),
		.gen3_coeff_17_sel_hwtcl                  ("preset_17"),
		.gen3_coeff_17_preset_hint_hwtcl          (0),
		.gen3_coeff_17_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_17_nxtber_more_hwtcl          ("g3_coeff_17_nxtber_more"),
		.gen3_coeff_17_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_17_nxtber_less_hwtcl          ("g3_coeff_17_nxtber_less"),
		.gen3_coeff_17_reqber_hwtcl               (0),
		.gen3_coeff_17_ber_meas_hwtcl             (0),
		.gen3_coeff_18_hwtcl                      (0),
		.gen3_coeff_18_sel_hwtcl                  ("preset_18"),
		.gen3_coeff_18_preset_hint_hwtcl          (0),
		.gen3_coeff_18_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_18_nxtber_more_hwtcl          ("g3_coeff_18_nxtber_more"),
		.gen3_coeff_18_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_18_nxtber_less_hwtcl          ("g3_coeff_18_nxtber_less"),
		.gen3_coeff_18_reqber_hwtcl               (0),
		.gen3_coeff_18_ber_meas_hwtcl             (0),
		.gen3_coeff_19_hwtcl                      (0),
		.gen3_coeff_19_sel_hwtcl                  ("preset_19"),
		.gen3_coeff_19_preset_hint_hwtcl          (0),
		.gen3_coeff_19_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_19_nxtber_more_hwtcl          ("g3_coeff_19_nxtber_more"),
		.gen3_coeff_19_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_19_nxtber_less_hwtcl          ("g3_coeff_19_nxtber_less"),
		.gen3_coeff_19_reqber_hwtcl               (0),
		.gen3_coeff_19_ber_meas_hwtcl             (0),
		.gen3_coeff_20_hwtcl                      (0),
		.gen3_coeff_20_sel_hwtcl                  ("preset_20"),
		.gen3_coeff_20_preset_hint_hwtcl          (0),
		.gen3_coeff_20_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_20_nxtber_more_hwtcl          ("g3_coeff_20_nxtber_more"),
		.gen3_coeff_20_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_20_nxtber_less_hwtcl          ("g3_coeff_20_nxtber_less"),
		.gen3_coeff_20_reqber_hwtcl               (0),
		.gen3_coeff_20_ber_meas_hwtcl             (0),
		.gen3_coeff_21_hwtcl                      (0),
		.gen3_coeff_21_sel_hwtcl                  ("preset_21"),
		.gen3_coeff_21_preset_hint_hwtcl          (0),
		.gen3_coeff_21_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_21_nxtber_more_hwtcl          ("g3_coeff_21_nxtber_more"),
		.gen3_coeff_21_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_21_nxtber_less_hwtcl          ("g3_coeff_21_nxtber_less"),
		.gen3_coeff_21_reqber_hwtcl               (0),
		.gen3_coeff_21_ber_meas_hwtcl             (0),
		.gen3_coeff_22_hwtcl                      (0),
		.gen3_coeff_22_sel_hwtcl                  ("preset_22"),
		.gen3_coeff_22_preset_hint_hwtcl          (0),
		.gen3_coeff_22_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_22_nxtber_more_hwtcl          ("g3_coeff_22_nxtber_more"),
		.gen3_coeff_22_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_22_nxtber_less_hwtcl          ("g3_coeff_22_nxtber_less"),
		.gen3_coeff_22_reqber_hwtcl               (0),
		.gen3_coeff_22_ber_meas_hwtcl             (0),
		.gen3_coeff_23_hwtcl                      (0),
		.gen3_coeff_23_sel_hwtcl                  ("preset_23"),
		.gen3_coeff_23_preset_hint_hwtcl          (0),
		.gen3_coeff_23_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_23_nxtber_more_hwtcl          ("g3_coeff_23_nxtber_more"),
		.gen3_coeff_23_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_23_nxtber_less_hwtcl          ("g3_coeff_23_nxtber_less"),
		.gen3_coeff_23_reqber_hwtcl               (0),
		.gen3_coeff_23_ber_meas_hwtcl             (0),
		.gen3_coeff_24_hwtcl                      (0),
		.gen3_coeff_24_sel_hwtcl                  ("preset_24"),
		.gen3_coeff_24_preset_hint_hwtcl          (0),
		.gen3_coeff_24_nxtber_more_ptr_hwtcl      (0),
		.gen3_coeff_24_nxtber_more_hwtcl          ("g3_coeff_24_nxtber_more"),
		.gen3_coeff_24_nxtber_less_ptr_hwtcl      (0),
		.gen3_coeff_24_nxtber_less_hwtcl          ("g3_coeff_24_nxtber_less"),
		.gen3_coeff_24_reqber_hwtcl               (0),
		.gen3_coeff_24_ber_meas_hwtcl             (0),
		.hwtcl_override_g3txcoef                  (0),
		.gen3_preset_coeff_1_hwtcl                (0),
		.gen3_preset_coeff_2_hwtcl                (0),
		.gen3_preset_coeff_3_hwtcl                (0),
		.gen3_preset_coeff_4_hwtcl                (0),
		.gen3_preset_coeff_5_hwtcl                (0),
		.gen3_preset_coeff_6_hwtcl                (0),
		.gen3_preset_coeff_7_hwtcl                (0),
		.gen3_preset_coeff_8_hwtcl                (0),
		.gen3_preset_coeff_9_hwtcl                (0),
		.gen3_preset_coeff_10_hwtcl               (0),
		.gen3_preset_coeff_11_hwtcl               (0),
		.gen3_low_freq_hwtcl                      (0),
		.full_swing_hwtcl                         (35),
		.gen3_full_swing_hwtcl                    (35),
		.use_atx_pll_hwtcl                        (0),
		.low_latency_mode_hwtcl                   (1)
	) pcie3_inst (
		.npor                   (npor),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //               npor.npor
		.pin_perst              (pin_perst),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .pin_perst
		.lmi_addr               (lmi_addr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                lmi.lmi_addr
		.lmi_din                (lmi_din),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .lmi_din
		.lmi_rden               (lmi_rden),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .lmi_rden
		.lmi_wren               (lmi_wren),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .lmi_wren
		.lmi_ack                (lmi_ack),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .lmi_ack
		.lmi_dout               (lmi_dout),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .lmi_dout
		.hpg_ctrler             (hpg_ctrler),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //          config_tl.hpg_ctrler
		.tl_cfg_add             (tl_cfg_add),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .tl_cfg_add
		.tl_cfg_ctl             (tl_cfg_ctl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .tl_cfg_ctl
		.tl_cfg_sts             (tl_cfg_sts),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .tl_cfg_sts
		.cpl_err                (cpl_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .cpl_err
		.cpl_pending            (cpl_pending),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .cpl_pending
		.pm_auxpwr              (pm_auxpwr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //         power_mngt.pm_auxpwr
		.pm_data                (pm_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .pm_data
		.pme_to_cr              (pme_to_cr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .pme_to_cr
		.pm_event               (pm_event),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .pm_event
		.pme_to_sr              (pme_to_sr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .pme_to_sr
		.rx_st_sop              (rx_st_sop),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //              rx_st.startofpacket
		.rx_st_eop              (rx_st_eop),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .endofpacket
		.rx_st_err              (rx_st_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .error
		.rx_st_valid            (rx_st_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .valid
		.rx_st_empty            (rx_st_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .empty
		.rx_st_ready            (rx_st_ready),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .ready
		.rx_st_data             (rx_st_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .data
		.rx_st_bar              (rx_st_bar),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //          rx_bar_be.rx_st_bar
		.rx_st_mask             (rx_st_mask),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .rx_st_mask
		.tx_st_sop              (tx_st_sop),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //              tx_st.startofpacket
		.tx_st_eop              (tx_st_eop),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .endofpacket
		.tx_st_err              (tx_st_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .error
		.tx_st_valid            (tx_st_valid),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .valid
		.tx_st_empty            (tx_st_empty),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .empty
		.tx_st_ready            (tx_st_ready),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .ready
		.tx_st_data             (tx_st_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .data
		.tx_cred_datafccp       (tx_cred_datafccp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //            tx_cred.tx_cred_datafccp
		.tx_cred_datafcnp       (tx_cred_datafcnp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .tx_cred_datafcnp
		.tx_cred_datafcp        (tx_cred_datafcp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .tx_cred_datafcp
		.tx_cred_fchipcons      (tx_cred_fchipcons),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .tx_cred_fchipcons
		.tx_cred_fcinfinite     (tx_cred_fcinfinite),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              //                   .tx_cred_fcinfinite
		.tx_cred_hdrfccp        (tx_cred_hdrfccp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .tx_cred_hdrfccp
		.tx_cred_hdrfcnp        (tx_cred_hdrfcnp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .tx_cred_hdrfcnp
		.tx_cred_hdrfcp         (tx_cred_hdrfcp),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .tx_cred_hdrfcp
		.pld_clk                (pld_clk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //            pld_clk.clk
		.coreclkout_hip         (coreclkout_hip),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //     coreclkout_hip.clk
		.refclk                 (refclk),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //             refclk.clk
		.reset_status           (reset_status),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //            hip_rst.reset_status
		.serdes_pll_locked      (serdes_pll_locked),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .serdes_pll_locked
		.pld_clk_inuse          (pld_clk_inuse),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .pld_clk_inuse
		.pld_core_ready         (pld_core_ready),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .pld_core_ready
		.testin_zero            (testin_zero),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .testin_zero
		.reconfig_to_xcvr       (reconfig_to_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr     (reconfig_from_xcvr),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              // reconfig_from_xcvr.reconfig_from_xcvr
		.rx_in0                 (rx_in0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //         hip_serial.rx_in0
		.rx_in1                 (rx_in1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_in1
		.rx_in2                 (rx_in2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_in2
		.rx_in3                 (rx_in3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_in3
		.rx_in4                 (rx_in4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_in4
		.rx_in5                 (rx_in5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_in5
		.rx_in6                 (rx_in6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_in6
		.rx_in7                 (rx_in7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //                   .rx_in7
		.tx_out0                (tx_out0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out0
		.tx_out1                (tx_out1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out1
		.tx_out2                (tx_out2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out2
		.tx_out3                (tx_out3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out3
		.tx_out4                (tx_out4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out4
		.tx_out5                (tx_out5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out5
		.tx_out6                (tx_out6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out6
		.tx_out7                (tx_out7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .tx_out7
		.sim_pipe_pclk_in       (sim_pipe_pclk_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //           hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate          (sim_pipe_rate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   //                   .sim_pipe_rate
		.sim_ltssmstate         (sim_ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .sim_ltssmstate
		.eidleinfersel0         (eidleinfersel0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel0
		.eidleinfersel1         (eidleinfersel1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel1
		.eidleinfersel2         (eidleinfersel2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel2
		.eidleinfersel3         (eidleinfersel3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel3
		.eidleinfersel4         (eidleinfersel4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel4
		.eidleinfersel5         (eidleinfersel5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel5
		.eidleinfersel6         (eidleinfersel6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel6
		.eidleinfersel7         (eidleinfersel7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .eidleinfersel7
		.powerdown0             (powerdown0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown0
		.powerdown1             (powerdown1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown1
		.powerdown2             (powerdown2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown2
		.powerdown3             (powerdown3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown3
		.powerdown4             (powerdown4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown4
		.powerdown5             (powerdown5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown5
		.powerdown6             (powerdown6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown6
		.powerdown7             (powerdown7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .powerdown7
		.rxpolarity0            (rxpolarity0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity0
		.rxpolarity1            (rxpolarity1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity1
		.rxpolarity2            (rxpolarity2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity2
		.rxpolarity3            (rxpolarity3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity3
		.rxpolarity4            (rxpolarity4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity4
		.rxpolarity5            (rxpolarity5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity5
		.rxpolarity6            (rxpolarity6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity6
		.rxpolarity7            (rxpolarity7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxpolarity7
		.txcompl0               (txcompl0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl0
		.txcompl1               (txcompl1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl1
		.txcompl2               (txcompl2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl2
		.txcompl3               (txcompl3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl3
		.txcompl4               (txcompl4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl4
		.txcompl5               (txcompl5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl5
		.txcompl6               (txcompl6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl6
		.txcompl7               (txcompl7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txcompl7
		.txdata0                (txdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata0
		.txdata1                (txdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata1
		.txdata2                (txdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata2
		.txdata3                (txdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata3
		.txdata4                (txdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata4
		.txdata5                (txdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata5
		.txdata6                (txdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata6
		.txdata7                (txdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .txdata7
		.txdatak0               (txdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak0
		.txdatak1               (txdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak1
		.txdatak2               (txdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak2
		.txdatak3               (txdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak3
		.txdatak4               (txdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak4
		.txdatak5               (txdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak5
		.txdatak6               (txdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak6
		.txdatak7               (txdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txdatak7
		.txdetectrx0            (txdetectrx0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx0
		.txdetectrx1            (txdetectrx1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx1
		.txdetectrx2            (txdetectrx2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx2
		.txdetectrx3            (txdetectrx3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx3
		.txdetectrx4            (txdetectrx4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx4
		.txdetectrx5            (txdetectrx5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx5
		.txdetectrx6            (txdetectrx6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx6
		.txdetectrx7            (txdetectrx7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txdetectrx7
		.txelecidle0            (txelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle0
		.txelecidle1            (txelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle1
		.txelecidle2            (txelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle2
		.txelecidle3            (txelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle3
		.txelecidle4            (txelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle4
		.txelecidle5            (txelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle5
		.txelecidle6            (txelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle6
		.txelecidle7            (txelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .txelecidle7
		.txdeemph0              (txdeemph0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph0
		.txdeemph1              (txdeemph1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph1
		.txdeemph2              (txdeemph2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph2
		.txdeemph3              (txdeemph3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph3
		.txdeemph4              (txdeemph4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph4
		.txdeemph5              (txdeemph5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph5
		.txdeemph6              (txdeemph6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph6
		.txdeemph7              (txdeemph7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txdeemph7
		.txmargin0              (txmargin0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin0
		.txmargin1              (txmargin1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin1
		.txmargin2              (txmargin2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin2
		.txmargin3              (txmargin3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin3
		.txmargin4              (txmargin4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin4
		.txmargin5              (txmargin5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin5
		.txmargin6              (txmargin6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin6
		.txmargin7              (txmargin7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .txmargin7
		.txswing0               (txswing0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing0
		.txswing1               (txswing1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing1
		.txswing2               (txswing2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing2
		.txswing3               (txswing3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing3
		.txswing4               (txswing4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing4
		.txswing5               (txswing5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing5
		.txswing6               (txswing6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing6
		.txswing7               (txswing7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .txswing7
		.phystatus0             (phystatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus0
		.phystatus1             (phystatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus1
		.phystatus2             (phystatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus2
		.phystatus3             (phystatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus3
		.phystatus4             (phystatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus4
		.phystatus5             (phystatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus5
		.phystatus6             (phystatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus6
		.phystatus7             (phystatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .phystatus7
		.rxdata0                (rxdata0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata0
		.rxdata1                (rxdata1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata1
		.rxdata2                (rxdata2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata2
		.rxdata3                (rxdata3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata3
		.rxdata4                (rxdata4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata4
		.rxdata5                (rxdata5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata5
		.rxdata6                (rxdata6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata6
		.rxdata7                (rxdata7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .rxdata7
		.rxdatak0               (rxdatak0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak0
		.rxdatak1               (rxdatak1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak1
		.rxdatak2               (rxdatak2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak2
		.rxdatak3               (rxdatak3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak3
		.rxdatak4               (rxdatak4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak4
		.rxdatak5               (rxdatak5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak5
		.rxdatak6               (rxdatak6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak6
		.rxdatak7               (rxdatak7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxdatak7
		.rxelecidle0            (rxelecidle0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle0
		.rxelecidle1            (rxelecidle1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle1
		.rxelecidle2            (rxelecidle2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle2
		.rxelecidle3            (rxelecidle3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle3
		.rxelecidle4            (rxelecidle4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle4
		.rxelecidle5            (rxelecidle5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle5
		.rxelecidle6            (rxelecidle6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle6
		.rxelecidle7            (rxelecidle7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .rxelecidle7
		.rxstatus0              (rxstatus0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus0
		.rxstatus1              (rxstatus1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus1
		.rxstatus2              (rxstatus2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus2
		.rxstatus3              (rxstatus3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus3
		.rxstatus4              (rxstatus4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus4
		.rxstatus5              (rxstatus5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus5
		.rxstatus6              (rxstatus6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus6
		.rxstatus7              (rxstatus7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .rxstatus7
		.rxvalid0               (rxvalid0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid0
		.rxvalid1               (rxvalid1),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid1
		.rxvalid2               (rxvalid2),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid2
		.rxvalid3               (rxvalid3),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid3
		.rxvalid4               (rxvalid4),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid4
		.rxvalid5               (rxvalid5),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid5
		.rxvalid6               (rxvalid6),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid6
		.rxvalid7               (rxvalid7),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .rxvalid7
		.app_int_sts            (app_int_sts),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //            int_msi.app_int_sts
		.app_msi_num            (app_msi_num),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .app_msi_num
		.app_msi_req            (app_msi_req),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .app_msi_req
		.app_msi_tc             (app_msi_tc),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .app_msi_tc
		.app_int_ack            (app_int_ack),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .app_int_ack
		.app_msi_ack            (app_msi_ack),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .app_msi_ack
		.test_in                (test_in),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //           hip_ctrl.test_in
		.simu_mode_pipe         (simu_mode_pipe),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //                   .simu_mode_pipe
		.derr_cor_ext_rcv       (derr_cor_ext_rcv),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //         hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl       (derr_cor_ext_rpl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //                   .derr_cor_ext_rpl
		.derr_rpl               (derr_rpl),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .derr_rpl
		.dlup                   (dlup),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //                   .dlup
		.dlup_exit              (dlup_exit),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       //                   .dlup_exit
		.ev128ns                (ev128ns),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .ev128ns
		.ev1us                  (ev1us),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //                   .ev1us
		.hotrst_exit            (hotrst_exit),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .hotrst_exit
		.int_status             (int_status),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .int_status
		.l2_exit                (l2_exit),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //                   .l2_exit
		.lane_act               (lane_act),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //                   .lane_act
		.ltssmstate             (ltssmstate),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .ltssmstate
		.rx_par_err             (rx_par_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .rx_par_err
		.tx_par_err             (tx_par_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //                   .tx_par_err
		.cfg_par_err            (cfg_par_err),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //                   .cfg_par_err
		.ko_cpl_spc_header      (ko_cpl_spc_header),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //                   .ko_cpl_spc_header
		.ko_cpl_spc_data        (ko_cpl_spc_data),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 //                   .ko_cpl_spc_data
		.currentspeed           (currentspeed),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    //   hip_currentspeed.currentspeed
		.rx_st_parity           (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.rx_st_be               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.tx_st_parity           (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.tx_cons_cred_sel       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.sim_pipe_pclk_out      (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.rxdataskip0            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip1            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip2            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip3            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip4            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip5            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip6            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxdataskip7            (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst0               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst1               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst2               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst3               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst4               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst5               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst6               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxblkst7               (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxsynchd0              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd1              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd2              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd3              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd4              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd5              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd6              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxsynchd7              (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.rxfreqlocked0          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked1          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked2          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked3          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked4          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked5          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked6          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.rxfreqlocked7          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.currentcoeff0          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff1          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff2          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff3          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff4          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff5          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff6          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentcoeff7          (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset0       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset1       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset2       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset3       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset4       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset5       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset6       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.currentrxpreset7       (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd0              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd1              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd2              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd3              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd4              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd5              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd6              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txsynchd7              (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst0               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst1               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst2               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst3               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst4               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst5               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst6               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.txblkst7               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.aer_msi_num            (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.pex_msi_num            (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.serr_out               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.hip_reconfig_clk       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_rst_n     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_address   (10'b0000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  //        (terminated)
		.hip_reconfig_read      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_write     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_writedata (16'b0000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.hip_reconfig_byte_en   (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.ser_shift_load         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.interface_sel          (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_link2csr         (13'b0000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               //        (terminated)
		.cfgbp_comclk_reg       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_extsy_reg        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_max_pload        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
		.cfgbp_tx_ecrcgen       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_rx_ecrchk        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_secbus           (8'b00000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     //        (terminated)
		.cfgbp_linkcsr_bit0     (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_tx_req_pm        (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_tx_typ_pm        (3'b000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          //        (terminated)
		.cfgbp_req_phypm        (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
		.cfgbp_req_phycfg       (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
		.cfgbp_vc0_tcmap_pld    (7'b0000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      //        (terminated)
		.cfgbp_inh_dllp         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_inh_tx_tlp       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_req_wake         (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cfgbp_link3_ctl        (2'b00),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           //        (terminated)
		.cseb_rddata            (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cseb_rdresponse        (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.cseb_waitrequest       (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cseb_wrresponse        (5'b00000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        //        (terminated)
		.cseb_wrresp_valid      (1'b0),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.cseb_rddata_parity     (4'b0000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         //        (terminated)
		.reservedin             (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            //        (terminated)
		.tlbfm_in               (),                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                //        (terminated)
		.tlbfm_out              (1001'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.rxfc_cplbuf_ovf        (),
		.debug                  (debug)
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2014 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_pcie_sv_hip_ast" version="14.0" >
// Retrieval info: 	<generic name="design_environment_hwtcl" value="NATIVE" />
// Retrieval info: 	<generic name="ACDS_VERSION_HWTCL" value="14.0" />
// Retrieval info: 	<generic name="INTENDED_DEVICE_FAMILY" value="Stratix V" />
// Retrieval info: 	<generic name="pcie_qsys" value="1" />
// Retrieval info: 	<generic name="lane_mask_hwtcl" value="x8" />
// Retrieval info: 	<generic name="gen123_lane_rate_mode_hwtcl" value="Gen3 (8.0 Gbps)" />
// Retrieval info: 	<generic name="port_type_hwtcl" value="Native endpoint" />
// Retrieval info: 	<generic name="pcie_spec_version_hwtcl" value="3.0" />
// Retrieval info: 	<generic name="ast_width_hwtcl" value="Avalon-ST 256-bit" />
// Retrieval info: 	<generic name="rxbuffer_rxreq_hwtcl" value="Low" />
// Retrieval info: 	<generic name="pll_refclk_freq_hwtcl" value="100 MHz" />
// Retrieval info: 	<generic name="set_pld_clk_x1_625MHz_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_rx_st_be_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_ast_parity" value="0" />
// Retrieval info: 	<generic name="multiple_packets_per_cycle_hwtcl" value="0" />
// Retrieval info: 	<generic name="in_cvp_mode_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_tx_cons_cred_sel_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_pci_ext_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_pcie_ext_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_config_bypass_hwtcl" value="0" />
// Retrieval info: 	<generic name="enable_tl_only_sim_hwtcl" value="0" />
// Retrieval info: 	<generic name="hip_reconfig_hwtcl" value="0" />
// Retrieval info: 	<generic name="hip_tag_checking_hwtcl" value="1" />
// Retrieval info: 	<generic name="enable_power_on_rst_pulse_hwtcl" value="0" />
// Retrieval info: 	<generic name="enable_pcisigtest_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar0_type_hwtcl" value="2" />
// Retrieval info: 	<generic name="bar0_size_mask_hwtcl" value="24" />
// Retrieval info: 	<generic name="bar1_type_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar1_size_mask_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar2_type_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar2_size_mask_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar3_type_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar3_size_mask_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar4_type_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar4_size_mask_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar5_type_hwtcl" value="0" />
// Retrieval info: 	<generic name="bar5_size_mask_hwtcl" value="0" />
// Retrieval info: 	<generic name="expansion_base_address_register_hwtcl" value="0" />
// Retrieval info: 	<generic name="io_window_addr_width_hwtcl" value="0" />
// Retrieval info: 	<generic name="prefetchable_mem_window_addr_width_hwtcl" value="0" />
// Retrieval info: 	<generic name="vendor_id_hwtcl" value="4466" />
// Retrieval info: 	<generic name="device_id_hwtcl" value="57345" />
// Retrieval info: 	<generic name="revision_id_hwtcl" value="1" />
// Retrieval info: 	<generic name="class_code_hwtcl" value="16711680" />
// Retrieval info: 	<generic name="subsystem_vendor_id_hwtcl" value="0" />
// Retrieval info: 	<generic name="subsystem_device_id_hwtcl" value="0" />
// Retrieval info: 	<generic name="max_payload_size_hwtcl" value="256" />
// Retrieval info: 	<generic name="extend_tag_field_hwtcl" value="32" />
// Retrieval info: 	<generic name="completion_timeout_hwtcl" value="ABCD" />
// Retrieval info: 	<generic name="enable_completion_timeout_disable_hwtcl" value="1" />
// Retrieval info: 	<generic name="use_aer_hwtcl" value="1" />
// Retrieval info: 	<generic name="ecrc_check_capable_hwtcl" value="0" />
// Retrieval info: 	<generic name="ecrc_gen_capable_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_crc_forwarding_hwtcl" value="0" />
// Retrieval info: 	<generic name="track_rxfc_cplbuf_ovf_hwtcl" value="0" />
// Retrieval info: 	<generic name="port_link_number_hwtcl" value="1" />
// Retrieval info: 	<generic name="dll_active_report_support_hwtcl" value="0" />
// Retrieval info: 	<generic name="surprise_down_error_support_hwtcl" value="0" />
// Retrieval info: 	<generic name="slotclkcfg_hwtcl" value="1" />
// Retrieval info: 	<generic name="msi_multi_message_capable_hwtcl" value="4" />
// Retrieval info: 	<generic name="msi_64bit_addressing_capable_hwtcl" value="true" />
// Retrieval info: 	<generic name="msi_masking_capable_hwtcl" value="false" />
// Retrieval info: 	<generic name="msi_support_hwtcl" value="true" />
// Retrieval info: 	<generic name="enable_function_msix_support_hwtcl" value="0" />
// Retrieval info: 	<generic name="msix_table_size_hwtcl" value="0" />
// Retrieval info: 	<generic name="msix_table_offset_hwtcl" value="0" />
// Retrieval info: 	<generic name="msix_table_bir_hwtcl" value="0" />
// Retrieval info: 	<generic name="msix_pba_offset_hwtcl" value="0" />
// Retrieval info: 	<generic name="msix_pba_bir_hwtcl" value="0" />
// Retrieval info: 	<generic name="enable_slot_register_hwtcl" value="0" />
// Retrieval info: 	<generic name="slot_power_scale_hwtcl" value="0" />
// Retrieval info: 	<generic name="slot_power_limit_hwtcl" value="0" />
// Retrieval info: 	<generic name="slot_number_hwtcl" value="0" />
// Retrieval info: 	<generic name="endpoint_l0_latency_hwtcl" value="0" />
// Retrieval info: 	<generic name="endpoint_l1_latency_hwtcl" value="0" />
// Retrieval info: 	<generic name="vsec_id_hwtcl" value="40960" />
// Retrieval info: 	<generic name="user_id_hwtcl" value="0" />
// Retrieval info: 	<generic name="vsec_rev_hwtcl" value="0" />
// Retrieval info: 	<generic name="pcie_toolkit_enable_hwtcl" value="false" />
// Retrieval info: 	<generic name="enable_pipe32_sim_hwtcl" value="0" />
// Retrieval info: 	<generic name="enable_pipe32_phyip_ser_driver_hwtcl" value="0" />
// Retrieval info: 	<generic name="fixed_preset_on" value="0" />
// Retrieval info: 	<generic name="advanced_default_parameter_override" value="0" />
// Retrieval info: 	<generic name="override_tbpartner_driver_setting_hwtcl" value="0" />
// Retrieval info: 	<generic name="override_rxbuffer_cred_preset" value="0" />
// Retrieval info: 	<generic name="gen3_rxfreqlock_counter_hwtcl" value="0" />
// Retrieval info: 	<generic name="force_hrc" value="0" />
// Retrieval info: 	<generic name="force_src" value="0" />
// Retrieval info: 	<generic name="serial_sim_hwtcl" value="1" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_bypass_cdc" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_enable_rx_buffer_checking" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_disable_link_x2_support" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_wrong_device_id" value="disable" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_data_pack_rx" value="disable" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_ltssm_1ms_timeout" value="disable" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_ltssm_freqlocked_check" value="disable" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_deskew_comma" value="com_deskw" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_device_number" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_pipex1_debug_sel" value="disable" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_pclk_out_sel" value="pclk" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_no_soft_reset" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_maximum_current" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_d1_support" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_d2_support" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_d0_pme" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_d1_pme" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_d2_pme" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_d3_hot_pme" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_d3_cold_pme" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_low_priority_vc" value="single_vc" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_disable_snoop_packet" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_enable_l1_aspm" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_set_l0s" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_l1_exit_latency_sameclock" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_l1_exit_latency_diffclock" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_hot_plug_support" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_extended_tag_reset" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_no_command_completed" value="true" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_interrupt_pin" value="inta" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_bridge_port_vga_enable" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_bridge_port_ssid_support" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_ssvid" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_ssid" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_eie_before_nfts_count" value="4" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_gen2_diffclock_nfts_count" value="255" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_gen2_sameclock_nfts_count" value="255" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_l0_exit_latency_sameclock" value="6" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_l0_exit_latency_diffclock" value="6" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_op_routing" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_op_completer_32bit" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_op_completer_64bit" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_cas_completer_128bit" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_ltr_mechanism" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_tph_completer" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_extended_format_field" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_atomic_malformed" value="true" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_flr_capability" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_enable_adapter_half_rate_mode" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_vc0_clk_enable" value="true" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_register_pipe_signals" value="false" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_skp_os_gen3_count" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_tx_cdc_almost_empty" value="5" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_rx_l0s_count_idl" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_cdc_dummy_insert_limit" value="11" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_ei_delay_powerdown_count" value="10" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_skp_os_schedule_count" value="0" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_fc_init_timer" value="1024" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_l01_entry_latency" value="31" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_flow_control_update_count" value="30" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_flow_control_timeout_count" value="200" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_retry_buffer_last_active_address" value="2047" />
// Retrieval info: 	<generic name="advanced_default_hwtcl_reserved_debug" value="0" />
// Retrieval info: 	<generic name="hwtcl_override_g2_txvod" value="1" />
// Retrieval info: 	<generic name="rpre_emph_a_val_hwtcl" value="9" />
// Retrieval info: 	<generic name="rpre_emph_b_val_hwtcl" value="0" />
// Retrieval info: 	<generic name="rpre_emph_c_val_hwtcl" value="16" />
// Retrieval info: 	<generic name="rpre_emph_d_val_hwtcl" value="13" />
// Retrieval info: 	<generic name="rpre_emph_e_val_hwtcl" value="5" />
// Retrieval info: 	<generic name="rvod_sel_a_val_hwtcl" value="42" />
// Retrieval info: 	<generic name="rvod_sel_b_val_hwtcl" value="38" />
// Retrieval info: 	<generic name="rvod_sel_c_val_hwtcl" value="38" />
// Retrieval info: 	<generic name="rvod_sel_d_val_hwtcl" value="43" />
// Retrieval info: 	<generic name="rvod_sel_e_val_hwtcl" value="15" />
// Retrieval info: 	<generic name="hwtcl_override_g3rxcoef" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_1_hwtcl" value="7" />
// Retrieval info: 	<generic name="gen3_coeff_1_sel_hwtcl" value="preset_1" />
// Retrieval info: 	<generic name="gen3_coeff_1_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_1_nxtber_more_ptr_hwtcl" value="1" />
// Retrieval info: 	<generic name="gen3_coeff_1_nxtber_more_hwtcl" value="g3_coeff_1_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_1_nxtber_less_ptr_hwtcl" value="1" />
// Retrieval info: 	<generic name="gen3_coeff_1_nxtber_less_hwtcl" value="g3_coeff_1_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_1_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_1_ber_meas_hwtcl" value="2" />
// Retrieval info: 	<generic name="gen3_coeff_2_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_2_sel_hwtcl" value="preset_2" />
// Retrieval info: 	<generic name="gen3_coeff_2_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_2_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_2_nxtber_more_hwtcl" value="g3_coeff_2_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_2_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_2_nxtber_less_hwtcl" value="g3_coeff_2_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_2_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_2_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_3_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_3_sel_hwtcl" value="preset_3" />
// Retrieval info: 	<generic name="gen3_coeff_3_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_3_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_3_nxtber_more_hwtcl" value="g3_coeff_3_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_3_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_3_nxtber_less_hwtcl" value="g3_coeff_3_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_3_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_3_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_4_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_4_sel_hwtcl" value="preset_4" />
// Retrieval info: 	<generic name="gen3_coeff_4_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_4_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_4_nxtber_more_hwtcl" value="g3_coeff_4_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_4_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_4_nxtber_less_hwtcl" value="g3_coeff_4_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_4_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_4_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_5_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_5_sel_hwtcl" value="preset_5" />
// Retrieval info: 	<generic name="gen3_coeff_5_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_5_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_5_nxtber_more_hwtcl" value="g3_coeff_5_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_5_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_5_nxtber_less_hwtcl" value="g3_coeff_5_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_5_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_5_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_6_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_6_sel_hwtcl" value="preset_6" />
// Retrieval info: 	<generic name="gen3_coeff_6_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_6_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_6_nxtber_more_hwtcl" value="g3_coeff_6_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_6_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_6_nxtber_less_hwtcl" value="g3_coeff_6_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_6_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_6_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_7_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_7_sel_hwtcl" value="preset_7" />
// Retrieval info: 	<generic name="gen3_coeff_7_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_7_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_7_nxtber_more_hwtcl" value="g3_coeff_7_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_7_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_7_nxtber_less_hwtcl" value="g3_coeff_7_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_7_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_7_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_8_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_8_sel_hwtcl" value="preset_8" />
// Retrieval info: 	<generic name="gen3_coeff_8_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_8_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_8_nxtber_more_hwtcl" value="g3_coeff_8_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_8_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_8_nxtber_less_hwtcl" value="g3_coeff_8_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_8_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_8_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_9_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_9_sel_hwtcl" value="preset_9" />
// Retrieval info: 	<generic name="gen3_coeff_9_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_9_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_9_nxtber_more_hwtcl" value="g3_coeff_9_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_9_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_9_nxtber_less_hwtcl" value="g3_coeff_9_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_9_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_9_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_10_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_10_sel_hwtcl" value="preset_10" />
// Retrieval info: 	<generic name="gen3_coeff_10_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_10_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_10_nxtber_more_hwtcl" value="g3_coeff_10_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_10_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_10_nxtber_less_hwtcl" value="g3_coeff_10_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_10_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_10_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_11_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_11_sel_hwtcl" value="preset_11" />
// Retrieval info: 	<generic name="gen3_coeff_11_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_11_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_11_nxtber_more_hwtcl" value="g3_coeff_11_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_11_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_11_nxtber_less_hwtcl" value="g3_coeff_11_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_11_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_11_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_12_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_12_sel_hwtcl" value="preset_12" />
// Retrieval info: 	<generic name="gen3_coeff_12_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_12_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_12_nxtber_more_hwtcl" value="g3_coeff_12_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_12_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_12_nxtber_less_hwtcl" value="g3_coeff_12_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_12_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_12_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_13_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_13_sel_hwtcl" value="preset_13" />
// Retrieval info: 	<generic name="gen3_coeff_13_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_13_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_13_nxtber_more_hwtcl" value="g3_coeff_13_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_13_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_13_nxtber_less_hwtcl" value="g3_coeff_13_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_13_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_13_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_14_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_14_sel_hwtcl" value="preset_14" />
// Retrieval info: 	<generic name="gen3_coeff_14_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_14_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_14_nxtber_more_hwtcl" value="g3_coeff_14_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_14_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_14_nxtber_less_hwtcl" value="g3_coeff_14_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_14_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_14_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_15_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_15_sel_hwtcl" value="preset_15" />
// Retrieval info: 	<generic name="gen3_coeff_15_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_15_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_15_nxtber_more_hwtcl" value="g3_coeff_15_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_15_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_15_nxtber_less_hwtcl" value="g3_coeff_15_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_15_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_15_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_16_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_16_sel_hwtcl" value="preset_16" />
// Retrieval info: 	<generic name="gen3_coeff_16_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_16_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_16_nxtber_more_hwtcl" value="g3_coeff_16_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_16_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_16_nxtber_less_hwtcl" value="g3_coeff_16_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_16_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_16_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_17_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_17_sel_hwtcl" value="preset_17" />
// Retrieval info: 	<generic name="gen3_coeff_17_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_17_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_17_nxtber_more_hwtcl" value="g3_coeff_17_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_17_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_17_nxtber_less_hwtcl" value="g3_coeff_17_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_17_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_17_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_18_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_18_sel_hwtcl" value="preset_18" />
// Retrieval info: 	<generic name="gen3_coeff_18_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_18_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_18_nxtber_more_hwtcl" value="g3_coeff_18_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_18_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_18_nxtber_less_hwtcl" value="g3_coeff_18_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_18_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_18_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_19_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_19_sel_hwtcl" value="preset_19" />
// Retrieval info: 	<generic name="gen3_coeff_19_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_19_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_19_nxtber_more_hwtcl" value="g3_coeff_19_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_19_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_19_nxtber_less_hwtcl" value="g3_coeff_19_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_19_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_19_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_20_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_20_sel_hwtcl" value="preset_20" />
// Retrieval info: 	<generic name="gen3_coeff_20_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_20_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_20_nxtber_more_hwtcl" value="g3_coeff_20_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_20_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_20_nxtber_less_hwtcl" value="g3_coeff_20_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_20_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_20_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_21_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_21_sel_hwtcl" value="preset_21" />
// Retrieval info: 	<generic name="gen3_coeff_21_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_21_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_21_nxtber_more_hwtcl" value="g3_coeff_21_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_21_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_21_nxtber_less_hwtcl" value="g3_coeff_21_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_21_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_21_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_22_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_22_sel_hwtcl" value="preset_22" />
// Retrieval info: 	<generic name="gen3_coeff_22_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_22_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_22_nxtber_more_hwtcl" value="g3_coeff_22_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_22_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_22_nxtber_less_hwtcl" value="g3_coeff_22_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_22_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_22_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_23_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_23_sel_hwtcl" value="preset_23" />
// Retrieval info: 	<generic name="gen3_coeff_23_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_23_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_23_nxtber_more_hwtcl" value="g3_coeff_23_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_23_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_23_nxtber_less_hwtcl" value="g3_coeff_23_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_23_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_23_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_24_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_24_sel_hwtcl" value="preset_24" />
// Retrieval info: 	<generic name="gen3_coeff_24_preset_hint_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_24_nxtber_more_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_24_nxtber_more_hwtcl" value="g3_coeff_24_nxtber_more" />
// Retrieval info: 	<generic name="gen3_coeff_24_nxtber_less_ptr_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_24_nxtber_less_hwtcl" value="g3_coeff_24_nxtber_less" />
// Retrieval info: 	<generic name="gen3_coeff_24_reqber_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_coeff_24_ber_meas_hwtcl" value="0" />
// Retrieval info: 	<generic name="hwtcl_override_g3txcoef" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_1_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_2_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_3_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_4_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_5_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_6_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_7_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_8_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_9_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_10_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_preset_coeff_11_hwtcl" value="0" />
// Retrieval info: 	<generic name="gen3_low_freq_hwtcl" value="0" />
// Retrieval info: 	<generic name="full_swing_hwtcl" value="35" />
// Retrieval info: 	<generic name="gen3_full_swing_hwtcl" value="35" />
// Retrieval info: 	<generic name="change_deemphasis_hwtcl" value="0" />
// Retrieval info: 	<generic name="use_atx_pll_hwtcl" value="0" />
// Retrieval info: 	<generic name="low_latency_mode_hwtcl" value="1" />
// Retrieval info: </instance>
// IPFS_FILES : pcie3.vo
// RELATED_FILES: pcie3.v, altpcie_sv_hip_ast_hwtcl.v, altpcie_hip_256_pipen1b.v, altpcie_rs_serdes.v, altpcie_rs_hip.v, altpcie_ptk.sv, altera_xcvr_functions.sv, sv_pcs.sv, sv_pcs_ch.sv, sv_pma.sv, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, sv_rx_pma.sv, sv_tx_pma.sv, sv_tx_pma_ch.sv, sv_xcvr_h.sv, sv_xcvr_avmm_csr.sv, sv_xcvr_avmm_dcd.sv, sv_xcvr_avmm.sv, sv_xcvr_data_adapter.sv, sv_xcvr_native.sv, sv_xcvr_plls.sv, alt_xcvr_resync.sv, sv_hssi_10g_rx_pcs_rbc.sv, sv_hssi_10g_tx_pcs_rbc.sv, sv_hssi_8g_rx_pcs_rbc.sv, sv_hssi_8g_tx_pcs_rbc.sv, sv_hssi_8g_pcs_aggregate_rbc.sv, sv_hssi_common_pcs_pma_interface_rbc.sv, sv_hssi_common_pld_pcs_interface_rbc.sv, sv_hssi_pipe_gen1_2_rbc.sv, sv_hssi_pipe_gen3_rbc.sv, sv_hssi_rx_pcs_pma_interface_rbc.sv, sv_hssi_rx_pld_pcs_interface_rbc.sv, sv_hssi_tx_pcs_pma_interface_rbc.sv, sv_hssi_tx_pld_pcs_interface_rbc.sv, sv_xcvr_emsip_adapter.sv, sv_xcvr_pipe_native.sv, alt_xcvr_reconfig_h.sv, altpcie_reconfig_driver.sv
