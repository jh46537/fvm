��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�c���]�uJ]�u����`�/�_.�~���8�l3V	n����H�|U�ݬ�h"�����~��ܓ �ňPZ%�ԄQ��muZ`{ܡ6�є����w�,��f�/�͑�g�؀Q���3�%��"�uVY����)��XSHq&�~�KK�a�pΊ��54X���m�ڬ��x�$\�i���#��,tL�)e� �;�ּ4�W���&�j�����O���2��1֖Eo�G�Kw��WW��{��+���;|�F)�)Bƻ�Sl�%��i�������:/?E(�k
�E���2Q�����C_���/J��Yq,4I4B��+��&����'N����k���UT����͍ԗ�D�c�Ă������FT�of�f��L�{�bU�����̖'�u�m+��5�D ��k��2f��wxR[ Beƃ��$���%�O.̃�49��ڳ\ �
�P8�mm*���_b� �����G��D�`ae�eV�;,�z�7��!���O�'����d�8͂c��KT a֮Y*���[5��f��£h>��|��~FF�hA���u��~oIT59��f�U���	���lz��m��W�}��㶺�%������J>�V��6�	Ch�u��}�o�d
l����s�*P"���z-Į��M��<�A� �d��QYc=jfp �gx����1��d�8��у8���s�d��JO�����ju{�$�� �� ��9V."�X�hE_��,#��v66}�	��u�+�th�����X��GC�s,S�F12�+�s�k3����~����ʒ�z��"�����{U|đ<���#��G�׃G�����dYM���7Z%����)�A�j�k�G�>�v�Fg*��"�Ն��c�p�3���M�|:ѿ]�ty��y�U�:R!G+��s)�<;���,K}�n���Xي����"�#I�a80:+�Y�G�[_e)H�4s��y��Q��!��N���l�Y	������o=��N;�F4e�4�TG!f�o�ho׌\��"��O�9kђ�0hN�������XX	�l�<&u�K7�I�ﰒ?��7��U�yHϷ������B9z�k�Cjż�Q�`'�CR����#і��񒢦�b#~�Ls|�̟�8������U�v�}�����	�
�D��7)������|��}L�ǲ��[m�.hs�7엑m�a��e�t�.$F�O/:/�\Ic���H煋`G^�;q���f��W2mP9�!v=�����9j)�B<��p?+���L�/��������wR��~f��2�c��>�W�EǦ���3ߦ�t~�����&_��G�;����9��,��H ` l!���wg��0�pN;���d�W�J�`��P��Sz�>{%Q%��a���^#l��Э��~}@&����J����G%4�9L]�fl���6yi���r���	9��N�����E7&\�HH줘����9�!W��-�����*�Riԟ��`��f#�m���;pi��S��>̮ �u �����k9u͍�sN	�1����/�w��@����IƔ����b,�ɑ���[y�	{N�[Y��fʉx�;{�'����rC���H~@��q��M��Hkw�P���0�b���E�T���m
GC&j�N�u��ÅVU�Ӌ�=Ǆ/����oUw��:nۨ��t�[:�F���	З�H�P�B��xʓh韵�����y>��/JL�l����f+"rg����������ci��7����4�9$m����O�4���'�9�)?����� R�2/L��sZ��72$&yH��\���و�Y)�@l����@f��i���db]�q*t��wC�s�M$a�7`��^�`� �����Q�����Zv�x\���I�h�gA��gR6�J�O卜���Ͷ�BfyL��;a�喣I�p�م���<�����\��j�P�9l�%UV�����`���t����S���CjEӯ>��+��[�Qt�YU�	���[?��nh�  ���PDd/l���� B�QԘ�yK[�
p���L<��=W`|LQ��#�T���+���\���h��	��s�y�ў`�6<o2�6L#�YJXi@�P�Yϩ��r��Y9�Qe�`�	���R�Z��x���Am�����M�&�zZ�]-��wH���7�'ʇ�[�y������Ħ)z9�%���l�!��xE�I���;�>�k_�U�55�G����+�F��,�gd�}�+�%�s�qH�Q-��Yq�ʈ,���o�&��r��#�c'? r�M�/&G%ܵ��;P�-�l��H����@��g������6䱅2�y�. �3�E�|�+����J-`�)�N��]��Q;����b���iR����;����r���4k+��#C��Z0�Sy��:�ECFZ�O)(O��x����ϵ,�R>l����)%+��C|h���Ro���w�+��!6d��LOцC�L�^���r��-m5{��B�R�\�Q��G�r���!����x���8��"o��W|��̝���e
�F�J��~ �SLǚ��2�EoHbp�߰d�:,��d�L^p�K�����M3�����jy�g�ݰ��մ�(�G�u�}��2Mu�3}2(��ǫ���z���m̫�
�rRe�+�W^<`(T
��C)Y.8A-^�/9Z(��|�=7�Z���,ȿD��o+�Gђ�QDy�s�������������(�,�<��p~�Z�+��X{e&���s�������C)��솛8ؠZ8�IY� �Y��"r=D�p�-c�1�"�E���`s��ӎ�NoU]�2�9��o��6�k�FK�ŋ1媱�yGf��0]%��qu���A.e_|�y�˕�3gT`���Bz����ms|��/�rY�W{xC���D�+�:��4ji}�`ڐ��2�l�؝�ؕ�����o��]�gc�h�#HF�/*�&�����ƸK�#�������o'�R�P@�S��I���]3�1l�n�K�T�k�w�NS�r��u!��*�f$=�3��Jv�����mg}ߏ����AZ�Y!B�T�(DA��2��\�T�	�J�l���j���w��H"�v+����[?��6�GrDºB=�+ a�gY����J1Ԛ}�*7C��M`ҍ�-puz$PYE�!�d6�u�V<ZL�D����A۰���Y��31�ַ��{�I��/��#[�H�@�� ��G(�^�X��C���۞
�l�_��>�拳=*V���m�Y،��)y��z��!Gڴ
�f.�3�5£ZJ�����0�߻BŻ�T�e���̐E�,3�؉�kv=w5x?5J	F�