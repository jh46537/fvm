��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�n�~Q��x�vHB>���8�'`m���v䪇��rBR�r�u@U�l�{�����߼.$8d�8y������kp���?g6�����o��_�H��J٠�O��d�,��l�f�%�Ч������L{ 	���,#����v��*�� f^��n	��j��Հ�*�uZ�ز��z�V�/Q�8�3CJf���}�0��G���g+��<��1�Gv��I��8�L���(\�+F�:�w�7~�?���ݵ
~�������G{I]H4���h!Z�f�(1�vO�{�$�m�~\�vYep9.�[wwHQ����-��\�nTF��A��q��&p��u�I��Y�	�Φn���فԮB��A���H�$��A$�{���۴$	p}�M���'d0����:�A�D�:W��̧���tvB��D[��Ѯ5�����i���W�K��}����gMS �#�w!����̮�=C�6���S4纕��'-m�y�;��-N�J�3-6��.�y�������8�Z=�GaV^��p5l7,�-���k6�$Ŀ�ؓb4icʙ�i�C��&فX���f0�ض�)����o7��p�w!��B-,�C&*���az��� #���ːi>ElrN+5��mF�_�57y���h�s�џ�,�.�ӹ�5ج$C�H9^��r��o��,--�^����pM`B�P���?�c���_�����@�u?Bt�,0'�7yM>�~_��6;� d���^�i�0�P�I��MDU�G|�L�����l�Cq� ��!���u�u�o���8!�-^
-G�Ac�'������wY�#�Á��C���JGWR+�g�ɀ����{4��&CI�1����RSѴ������&KW�+G>�i�@y{9=�iε�gn�*�ʈ�v�s�T�b5� ���ǒ�������BP�dʾ\l;�0x�Z	�2 k�%�&_c�Z8��;��t���r?J��½�B���5z�`�F�|��c�`���~����?��v�;����X��D+]���f�
�n �����ѫ<6�ZF� 
x��G�6M-��5��X
�`�Uд��8��!��ri���"��:=[~���S�?ޟT�e�`��)��!Ί��
�u
 r*���.�柤M'��$��6����x'� �v���-(��U��MK��̐3��X��՚�om���J��/Dł#���\.� ���n8����+;¹6��}�U��Q6L`�lnz�E�1�f� �D�39([x�X�M�j���F1�{�$�p�Oa����������j���h����)�>}��q��3����O=l��r�!b�9�U�zB�q/Fث���.�{j�n�7� ����K��@QF��'>�TM����aq����ك��a�\��KI���gz�,��_~��o���{���{�솸�ұ�Lr����.�FE(kz��.�Ր����5��M�_������V'��"﹑�aS].�Ki��8z�M��A5kKi��������z̼����ow+hF�YO���q���y���
{���t��IK��N��]�!Z��f�.c��$a����t+Gt����[Ta�_����]/n�y4�wm.�nRs�K��AbH�a�(�פ��w~U�&.��o��] � i�q�������ì t��Gw~ۛ�(8������^0�F�2���O�1	�D�t.��x�!+@�%���zI��R��"��qɰr�^	��5j�Z��c�jt�&��ȶ�Nb^�W9��+��Fک�X{0�� �Ӆ#�:���Q$���8ɨVVvG�=
	q4�%�P�ZVE@�w���w������� u�<�IC�2P�����o����N��ּ[�̧���.����h��kg�\�}��[�*�����_�7��1lϤ�U�ODr{ࡇQx%��fQx�uF>͇=�ޔ��._wLң9(��j<�� �Y/ �v�O�=�e�|xU�O��@�@�Z�dl�q"JK���C�գJR{�!�r!��<�"17�Ӟ�=����q1Q'nk��"�b���7Z��Y�c�ߧXf&:��%e	�?D��ax~1���kXd�>��2s�@�_8m-�3���F�a�C�S������Vi� ZZ?%j���@о�-1�g�%q���HC^)DeO�P��tF~�:�#Af]��2~������g賬0��t�Y,���*Θ9GGr���n�UaC*���Ġ�u�g��]Q��"n6�N��Un�(�ǹ7�84���FM�r�l�F�H���,gޫ��| 1���>h�b��b.��"آ]��]AG�8������(�yMz�Η���\��?Ԅ,��c����e�[���\thNg*MıM��o.��+-�)��͔jX��`61�Ir��p�2Y1)��,;ĺ�a����q���M&�YuP>�]j�a�,�E'���y����a�S5C����dZ��a�YI���:e!+��z�2�&�&rh�RC�B���=��)CLn޵\�V�g2x�zx�(�+�:�4��%u�#�Z��F�����V��N&�C��(E6G��֦�f^�����;�I뿒y��a���<��`!L (��ٙ:��|7t��=]*�.�D��4�b,��DqȾ��̄(3�$��`a#wb@�o����~��q����#;��A�(�&��d����q�`�r�ɕRPb:�N���<q������^�k�l�~����~��s��0��aO��`���1�l��n�3���!ѹ�������!��pt���r���p�+���w�8�nP�e���ě:�ԙ~WM��µ�1�}8�����F|��.Y�5��ȴ�]n�-U#�-z:j��/\	�]Jv3��*��U�J)�91����S&��'��+���b�@��22�C�N<�-�b�ā�ڃ��\sg�9�'�w�Uo��k+sE�,�R8���>Ğ"��Q�������M��zچc�3�06�כ�/P��b��rWCjd��q<��!!�SfH(!.��"Z�%փ5�j]ӗAn�p�0���s��N�u2^Yj�D1�0Iql�������^n+�a�<��o��d�#�i�b��*X� :O Ji��8��!���_@M=W�n���N߭���d�C%��Ox5��:JH'��x�J�5�1�1��ChX�����gr��`�DX5��08��a�<��'k��9�0"��k�h,kdf�>;\�,o�o���d$�6'�,�L�!����-E�����]������[����C� �LĐ��h(�.ɘ��<a%�JtFFc/G�F�&��g/W�=>�մf�KsA"� �]�C\��;�����ƧoLO�Q'ي��$ǲ�4:��lO$�\�F$��Ӗ��]	�#��Ɇ�'Mz <�N�4�+V�ؽ�S���0 m"���Ł�e.[t�(�˹��
V�Ee��Zz�'�q�Si!]��8��y�N�$rn��!Y��{+���<�ƌF���C]$B�a�t�͸HPB�у��,�y#H�!�O!O��m-��	��T�G1��m�T5����^�M��LV0y+h38��~�Q)'Ăλc�������f��a߈�t�^zZ)����J�F.����o ����JC`Hzw���~�jiy%<��~��t[f͟U�x��'����n�@���aJ5��s�8K�;���%jF@����pvҗ{v#���L�a�����H�"�+&$�^8��Y�<��N�)�,�S��0�R��:��A��(rQ��u:�w]�#Q�|NŶ��k6�1���������f9�����H���L7�}������m�OVwB�|)P�������_	��w�.��	<9Bq��ґtl�Rs�곎�(=@GԾ�9��Q�b�Y��OMdX}��C��S���Tk���;y�95�ǂ���/Ky�a�ϝ��Z�y3=�������2~�3�.�|�3'K4uز״�f��CX��"6�jͧ9Ʊp�Qd,YA�=TtT��n�������6�2�ħr�)	��}<O��e}3�x��7��n��Jy?�����a~˟��b��#�GG��*�<�Ƽ��=��J�5�?.~VL5s���,�8� �Ҽ�v�f3���c��N�K����G7?��J4v����v����_����QK��
����Aw��id�Ķ3��b��Y�^-��slǉYT��8}i>@K�ѭ�~D�L��i�LTt���2���B����ˍT���`l�$��z�a&�aQ��9�&V.%���s��q�g-+3�!��h�a��T�|�)�����,t��!�v��{}H�k���񚱟=y�#Go�=���W���3�����ռHNCl�zp|�3x�z�p��x��B� ���ߒ��K����M���8�e�QhF�(t��e�%������NoƂ ��o�m*��i�Fyo�R�����]���;m��h�j(�}=���ю��ݦ��A��=cı�e٥！�94F����+���fW(�_�ի�O����>*�zsЭ�T���Sk�o@�L|���od8)^�'`��܏z�+������0�F7�rvvϖO��(ͻ�4�8�1�/`y���`o#(�ZuˊS�V=�����=��TƑM��KXf�|8pՍ����ߘ�|��Wdp��d����&Bd}�x�����z��y�D:�Dt�KE�B^M\��+#zbo,�S���
ڂE�OGZ���f$}V!^�:�`B>�q�8�,׾EK�]z87����<zƒ�~D�w��+L?�pp���L�P2H�V�L�ӧM�z/~3I��ȥ��z6C1�;��ZrQ��O/~+ϥ�9x]1
�o�	`�0IX'��k��ҕ�(J*	�~T�WLCb�'�O�v�rU�gX�,���tC?�sƛ8���'7�i�z~ӛ�J���$B^�p�$�~��(�PI�2R��W1.�^�~�`��M�4��R��Q�qw2R�͊&p�G�J:7��w�-(�j�9,/���S�40�޸�҉#��IA
���Z֝��V���`�uE@H��zj4e���|ՇN|>#:I0(5��ɨ�����4�?�Yi/�kу+�Ih�؏V��N��Vi��G�<�'��"�I8�g�忉�0�WE����<P[����;�h�\4�G)�K^(2���۵ΨVu�d���[���6vgɡe����<Y���0S���*X�L)�}\��fM'o�2��O���g��9B�[f�ѩW�&�OK�&�"Ð���m��TW���\/a%V'E�%�u�ċ#���D�~1�nf�a����c���zD�F}_�KQ�-�q��2"�)z,��\��*���Ay��+F!9��;���u9s�����:�xJ���t��0G�d�r����