��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�-No�?�j:C�]�;�%Q7�j&N�fV� �&��o},�<ӈ2�����MI�(4�E�@mm 2I�.Ǽ�j����}L��Mx���RS�xu��e�n{?8y��นm�(��)*����2����5Au����;��jl2���ܮ���[��{h�pSb��l�g+�-O6�`��F���\��N �a��%,����zA!I��JLBICU��J��g�,�0�fRf�a�K�m}�}b�P���.Y��tt�5:MC�Xj&|L����9�w�X�eA��[8��?H�_��Z��/"��� � -Bo�/ύ�(�3p"�=z�jd�t٧0�g�n�y�b�N�B�C�4�#��:@ Hgͤ�5�eO�C�r�A:�Zs�%�g�z�l"����4t�����7H�j��E"�|F'o���Ͱl9iG����l�?�X�h�V�ApY¼o[�&��ǡ���tj�9�@�Z��3c���Ff�A�j(>\nP��{��S��aL��<�xc]P���U!���:G�`��j�W>W�4���-��PT*~��5#ǓLD;h�10��߀�lg��B��.ܭ��2�*l%��?!W�L�ۤ�a�X��EcO$+^��O�i/�XTR4��������GiX��q�y^�z����Y�F�e����i�t��v?���DTpܤ�|o�l-�NW¹��B������U.̄S#y	����ZR	�ߓ��hF
�=�.#��`���t�v*&|�U�瞶�xT��Q"�����G�h�N�C��+��/��~,[$�fz�61k�[Uh2�JKi�ڀ�T5T\(G��h��QT�ěu���1ޠa)��}�b��0���;L��;���Q!�D��*/����W(w����BF*�^iE'�ͱÃ�=-� ߹2�9����������F�g�>=�BsCq��#�;�foiZᶒ��ZȰ#�%.Y�z_R�?ԣH=q��� q\�rd<��`�l#��C��x�Bq���g�C�%�:��Y>A�]-=Z�a:�A�V,�k�fu�W�]�?�#��5l�n�O��4�n���q�u�"K/5`@�Lp��\����W�o��r}���Ri�x;��H�8}��+��)��J��xH������[K���!y�wy?8�:����UuU,���ث���:���=��V)XY�"��R��{����aTO)	^��ϝ�`%�����tC����h��5Po����'�8b(uC��*c��'���7"6������yiZ)f`���9����GWi?��<=�T�,�|C�5��(�n*/�#�0"��}�;�.�x6[�i�$![D�H�k�Z~먥d]F\�k���JW������\��	�aa^�v�hթ&�E
�}�hX�Z;4ô�doPAmuXt����"�ϋ�Nq���?2�vy�&�jq��c0p�Ȭ}:!���^���a� ���(聸E$�Å\'	����\t�B��ڛ�XC(~���9.,�?>��^#9̟�B,�5\G��s���$�=����o��)D��K�����8���tWPG��7h�^ٵ�Kxޙ�A����w$Q�T+�\?�r���E߼��˕���=ʯ7!'+���{�����V��i��ϫ�����F�І�Xuk@�\�@l~��W��z�҅�Q��D۳o)��b,��S����</��6½~��_�Q����am����QIfʛ'�����s�E5.i�c��#M
tr�Ny�y��.?�iڦ�����h�o_3�Ȁ(P�oE^b!�K7�='L)�-1Yko{���R��%�8�U���%M'8�+E`|��K�G���L����n<.�S	�A� ^+4���\�B���%֜~3��,�es�t��1 V��靨H���^��CNc��G��O8e�a֕I�5�;����'.D�h�[*��O�z�z�L�d���lT����G�����P���I��ޟS~F�q�c$1�����V�P�{k�Uz3I��|����0�x`���I\j�N3�lk/�l�"%�.f蹒����7�(
 �4��I,���r�2�-�N���_�����ׂ��ܒ\�Z^�O{ѕS����e������-�!��ؾT���pX(}�����4�\4������@n�V�ti�m+���,>Y��jtJ���B�bϡ��>}���A5ت�(Bg�^��z�Is.v��|� G� ���Z�*ַ!KZ9o���d���;����F)�w]�Hr������ �6��/4?+<����r�~�gL	�򘢕�`x i_�C��65
E�VFB8���B?>�X��i������8�pG�J��{rI��ĳ��2�]�;B��V��x�;!2sc/ ��#��d��Ԕ�T���ǁEL�ܰ"���C�-���zA�ã��aU�n���A�O`��1i�+6�����������A�A�߄__8�����ҝ�ӯ��o��A�R�0�Xj�!d{N�R�3LONg1,$Y��v3b0F�m��������c�3EZ��QM2�b?��:��2��pO.�^���cy\����ٙ.W�O�1��Ź�w���/�
#TD���� 4��xݮ�����靫�����b���~�L|)�C�^au���}'�t\n��M�PA�$�ɉlSl�p�v^�a�u�kV�w�K7�b����C8�K}��5`�nV����O�8R~c+yֻe�)�U\X�P؈�݌`�i<^c`7
	���I�F�f���NA��=�����.P����R�i��zۿ��e%t��0\N�g�0
��5�p��L�'ȿC]��s羏+񩈕�@|?Ϝ8�t���e�PM��!��U���1\�6�s��Q�"[�(��P�:!��)��Y#���jy�^��JLP�w�����g����ua5��{�j�YMx�le.�O�k��B��
*�C��}�E��UՑ3�'�!�>��30�<Iz�Κo▕�5�G�b�l�&c�"��J"�]̏��AIblwz�_�P��Vf��������}/_<�&�^�l1|�M����]�y6�zZt�J[���.t$���m���&���i� s�ҿ�c�,^���m����D��Ƒ�rz�����k���ʆB����z��f��,{H�Qpf��K��JQ;��  YQV����0=�;!58�f��m���
��GC���-�4@z��g��T�,,�5�n�+O?P-�a��6��`X��<�f/8s�_�Kj��%����I�Pmh ����c,0����I"4r��y>��(;Ps�~̞6%���R�v2�T���cX��