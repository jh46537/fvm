��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�y�Sy�;��>��&�MA�)Cʌtg���e�8~�����=H�9����.k������U��U�Xe���M�b�(	
'�m��_�S,(
>ɢ&T^5�[Kم~�WA��Mb�c#�<˃#:}��6͕��F��O�j�7���'AF�9��'�ƹrq�9�p�
o�'�w=��v��("�|��ӏ�I�\.�V�����)���cB�չ6�t3sꀚ u?�({��_x�W������!�`�e�H�H���|�-�YY�
ꆞ �Ӟ냨��e���S�kFd�v�e����y�*D���G�>����+�ᩜu�f�x�I���*��/1\1����r�2�*M_�4j�t�'{)ȳ:�A��!���ש��6�D`��Js�[�a�O[�G�O.�����}�9�����E���;I҄0"}̙�������@pi?%D;�4�Q��L�<Cat��jB%Ra��68:�*�w=�M;�mӠ �1"9��2P�}����2�S���%*�G�;#�-\�-4:�nI�`�>3)��2�'ɇg������'�a�h���_�Ӳ8V}*S������O��.����8����O�v��$lc�^��4hf�2qw��SA����)���'l���<�� �/r����-�t'c�������._��l�ө�R1*���\�ɜz_�&c[�Hk���I�䵧0��nBzB��h�!�h��>��W�c�/�,����L�Х){K7��(~���1�^:DmA��ק�B?�d��
�)(���_��u�ۍ.!Ȣ�ZE9��ꥵ����A���%��A�8�l�����W3ۉ���D��j������3��hqz�U������"<C3��
��[-D�,�r3�]ˉ�28��D�L�$�����ʹ�ʬ��v�"a��ܩi2��/�rHh��Z�p�g�Ce/.J�������F�[��N�hh��!�NV�`hS�>�И�*Ou@@���,dDvc�x'I�B۾���\)��G���?x�]��t)���Tu�Ġg���tґ�Y�����Tt�͢�բЍ�=k�P`�<?��:�w�o- ���iEk�c���gH�#������z��/�"�^��Ȯ:�� @֙�����eP���\�Y��q'b6��el<� ���ȼ��ҏq�x�pThtR��6�$@���=�l84`��z$��Y��N�D�=X�'}h�Y5*��mBלm�	+Ҧ5��"�4'�:��#�ҝr�h�4�(L�Guh�� �[�۳~��J��QV!�
<3�NZz���1e�z3�+?�<J��R�;Ѝ8A#��?�`�S�w�^��jp������#��٨O�Xe.�iJ;_c�U�3�*�9���5L�:�ܑ� �X�OO����An&U��VO*ֆ��&����C��L�#�6{�-ݪ�������׏�����.�F*n��C��'�`�{N���P7���"PT&�L���}������)��BiϹ!`UV&����B*���Q�H�x>��c㠺KF�R�~��Q���j�˔
��ɉA����e_B�v�׽h�2�/Z��Fϊ�a����#~�Z�$"�x�|ϴ��^�b��1g@l8+RE�꾒5�c|@���ӥd�7��4y�Մr���y�́9�L�G�^W9��рI�pz	��=K�r�a	������E�U�j�Qm����r�%/��u�F.���]���ף��~Kļ{p��m9���sWD_�σ���IR�^@��UL��	`�T�u����@^V͗S����f.FF\M*ýЏ�=#�:���h�`n��HzI�ᖿ	�U����'�-��v���=Ee��C�����sS�������sm�u���q�$�%"��bi$d(N������L��X[�	��ˆ|�G�d�@��k��c��.ޅO��%��7h���j���a���c�GJ�ݛT�A�ir!x.�;��dNh~�>�c�4�$��DߺM8\��W����e�os�6C'RƠ�φy��p}��rh��ۊ�����LDk�e�=m�A6������J1{I��Ya�V�R����]�id&K^`um�@�'�����26��ڲLk�(r�����ڰ���p$9�1p.ό){�T��LTa�US�7����>�'��b���F�m��-��ųũ�U�R#4�:�"ˑXΒm�UO����Q�c�UO�B]Mt@^�j�5���^2u�3iw��sͥG����8"���T� ����?�qr����3�<l�r��D��diѝf�L>Ѯ*-Q(�~b�=��hB5<�p/��;�0�3r��Q��<� |�O[�:L���Nm��:�K�IQU ��3�T�*r�K�W���F�_�l?.q�7m'������|)}�ߡ�[��cիW�Z��R�	�z��tz�'�9-���!�N3f^�K������V���eV�}��nĉCV>���˿��w�uK'~��<I}���QҭG��5'�jD�;u|����B��0V��&pzl��h�su����s��.�A��ч�����s@'L�|hހ�ܧ)�,��b���y1�tnH�Lߍ�<��b�� ̨FuFTbE��/O�g��Ra @ۭ�bd��>��lA���F�=X��@��#���:�&)��p��FiA�2ڧL�lDKn��>���u����*�f�"�v�ېŵ^VމK>NA�X1��~�P����rV���*~�Ҿew��[�'mt1�o�f���f�0u��\��U��*^>c�ڸ�_�R�Z�5,�ߤ�~�B�:�G����ӗ�>r;���� <��ld�/-�WƎ��d�>)s\L,��Q!{T h�ӻ�*R���=eD|�G�qt�$���k�糙���ߦ�#�8�W�\5	qk�j=>�L�5�nv��!�C�*�S�w��q��/'P���M��8̲o���x��I���i��%����i���/]����V!�)��]j>3F�T!�K�������x6��ͧ<g�
^����L��&]��s��(�("�e����}O
ر+c8¬�L�{��1��:Zr<�H�k`�r�l�x��~\YIG�BX�{uࢋ�eN�rh��v.?�B:@_���.��`�=���%PO(��j5�D-���ܘU+�>Qȹ����:F+�@�mWd$l`m����)���Q��3��n�C�?}������r�H��qlDd�2G{�����e�w���kS49�S�d��*ʉ�ZoW� �K?��*YM�\w)!U�da�q��g�r2��FKca��-z-W%����9u�tʲt8�e	Ee_^ ���`���+��2�?��e��ˍ�SVz>�艀�@�kY��99�'n��A$mW����6s��%e�H��� '}��	w)�tR��w����3���c������X�3PGy��A��_�_�����l�b���vH]��	�e/o*�|]e��z�����H����{��\���c���!g]I����ٽXSL����|3%/@�BK5c������J�F�@&��xbZ��A������4���N\�:��.ĲWs,���{9��u�Nɾ�azeIw�}_腒= �>�ߘ�%>v�p:�<&�Y�ƴ��&����st��^��L��=T�������VS��3H-f%N��ŴD��5�nөh���,��#Rp�L6��Q��¨���"]^%��t���.�|�F�)���*.:̓/}b�u}n$�����!6O�����3�9YRJ���a[m-����M?;͊�WU�@S��h�R�+�+�ݦ���[�dB��K��e@������6[2ˉ��  �dL�-�ofE����Y?�����
S'��J�:�A�]}�	_�ф- �v�wm�Y2�X�w��	���m{��cޞDc 0�"�o�qX]��O���h��P���[�S�p�z��c~�%)��?���S�qv�&IcH��@v'�W������CТ���;������
O�z����߼s��H��We�|1�w��Ro��-�ٱ�e�G{
#�K�"Q%��&"fѐ3�I�O}]�4$ s�c]6�؁�u�C�/d���.��j	¸�<~���.N���Q�e�G�B�v۫��e������P>zy���.s�m8��E������>����$^�(��g��ˊ��9��!ۂ�	������%����a�g����%�1U�V��=X�& v�H
���Bڲ:L��+�t�I�Ahޚ�t�\	T�B�clEN����Ά�[�2�R6[��f�8�冷�B����c�%v9�&C�`����yo%kN��CU脸`EX��0������nϴ���B7}]�1�$�o��\0X%*���9����=���"���T�/�Y`#��z^�^0��.���=f�F7PR�!�A|2�����_+ŏ���i�F �"\������R9*F|j��;4����M�!��[�i,
��prx�	o[83`�SȰN�$h��K'��r���%Jh<�۷�K����=��.�J5 ��/�w׈�M�)E�8��W(���UZyTo�o��@gbA��3CL.�Mi��:um���.�	K_y��8l�&�M��b}��-Me��Yh�Xn�������[%��P܄g��,�����d<�V�K�z�S������VYo�ȶޛ<�
<5�X�u$i�е�'KWۧ{���<f��g褾�u u�:''JۋU��)�R� |�;�w5�4��>Z��E"t�+���J{(�3�:�vjxX�mqtSu(-�	���h�(�?u�u��.E�7�]���Y�̶��N}ߚ��b
��W�$��el��;�+����vpS�.P���Y�h�gDL&y&�9��V��6~�j��"x�N��#i{�{b`�	^��ۯ�T���B�+��EnH��3h��N�[�A)��߅��~c%�� Ȗ��J7�jɴ�6�a���@��ϩ����o�R �����v��
��4��@����45��<�k�L>V&�Vqd��T����h��FC��(�:�&�u��cI���mE̌}M(V�������כ�a��>3�(��pp�_҄p��'��5���rlTEqZW9�Y�\�_0��i�넎��!�:���I��V�P�ȯ�<w:r{T^���V��)�i��-�;C~�`� >�&dK��:KbM���Z5Is�mNɏ��g�'�B�pG�j�
�|��8Pg�Ğ7��na�O�n�hk-̺^���y��ıJ�m�dÈ6���0h]���L��xT�c�W�>� ��`O�yF�8ǋZo�k�9�L�D3ʓ�ΞF�2 Ȳ�N��6��ў��%^�$ZS7�$bZ	k�5G�r�M���<�ɺ_�lrL�;!Ӥ~��#}�P�.=��e2��܄c��)���H����UK��B���W_�5�v�Z=��Kj�~�}Ď�򶹶�$z�Ik$5.�Q�\���9m�[�1�yMc'�$`�#x�bwc/����o�iB���2�t�Ӑ����K6[CHrf-g���K���E��R#��h��`H�H���
� P��d'b���ʀi���qAų�Qr�w�չ�1,i�
Ұ�s����0��ʑ {nЎu66>�m��.��5��k|p�	p-k��m3W. ��x����w6�Bg�w��^?n�8l��5��K_h�2�*6�ZB�.�VT[f�'`?���u�Q������qy�b#��#���o�u��렰v�1�������B}��=��6���˘�!�Y8��V#+M��f�Dˁ�^"r�@�25���v��*����\�03�,K�S��T�a�%z��/]֯�:�����!�������Bp�7�]� L^Ho�fx�����;�_v�r$������e���o��qy���!63]�T�_��x�^�^�	�]4��ؚ_C���rpIE����ç�G�[^������zp�O�	:	�?A���if�K�R"h�O��t/�wl�T603�\Q,p�w�=��T��Ifg�W%��u
�(L`Jl���L���