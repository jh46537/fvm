��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~�HA�W���~�Z�T�K����"�1z���.XӜ[>�iq�)�R���D{���*�ۍ�;�*�Yɝ�,nS5��z���.�? ���H��&��:U�Ԯ�`Y�բ��$� ���>8ՉU_M6��B��˲i���	7��� �a���6̷v%%1��c��#��\�<�p�-������=6����a��ڍ
����E�$�]<G��SbS�v�KJ�P��@q0������9���P�0FzdY��(&!~@ɵ> hRU�Í�z�4�	y�v�ޭ��'TbA�Q�g��-�i�Ӟ���\�2�s�slʿ#��ԇ�ķ� �hnZ|Gzu-�6qG�C*��+B��.�o���s������q�`���|���M�7O�/�'���'.��uq�3�x.�f�	���N|��"L��i�Q.�Z���ްtl{���p�{mc�(�	 �?����v[�r⸷�?�W��i%�,���T&��T�=���8:]�NM���-�պyf<ٟ�zX�V]��C"��oft&�g48�mv��vE�?���1�S�!1W�=�v��|e�{ޅMH���ġ������k#>�l��
������Ԛ�M�D�C���Vò�E�$�2RW���Ib/�_��~����&�RP'�ȱ�.��r�������i%I��b3R��pJz�i}3�͐�H �h0GR:}-m�1䫄����cg�-�H8L��G2�c�Ko�;u����9�&�e���D���Eh���plfq������8�K�E����K1�Z��^J�@�����x��L���s-��i�^�xLi`�D#��^f�jjO����g�VN#	� N��Z� �ܙh^�c?W=�S��~\�v�8A��؏㤙�`J���nv���C�_��/��)�5������aA�^[��<�-KO-��
��,a/��uG�$�@��v�2i翌�b^$l�|3X���9�\P�jyN�B��:>�:$�kY{]�kv�t5Yw��8�aې���CmkBĬ��G��p�n�ҿ�`@�Ds�U�� �.� ��>`��/��>��y���8�1�<��kҠГLpO���K(E� K�2/Ɋ�� �&�yi�Fjj��xvzg�9F_��/���0q�Ӧe�o�#K�U�L@��w3�	>�ʲO^$� �P^�=
wm�;Fnݤ2�?��Bl6~�I���GCp�ݒI��eQ6E�']�L�%Arr�R5P!~��V���>'5h�58�R�gm%�;q���_���ݷZ_\H�v��5ǝ�z�^~_����#��0�Bv�!����TGQ�?��hDЬ�E�����m�|�@��Q�Z����6�����R�:��E!�+���Q�hSٯ\���x�an�0@q���;x��m�!�ǩv(`�>�L�[/PB������V�/�۲�aA���[��d���e��I�>%G)��h�oS���}_Y9Yl���L�Cr��V�0ވ.���f��ɃN27΁�7y�m��c0x0wmHd�*����PfH��϶�!�3���y�� Ďu5��G�2'�V/�$!��������&�m*m�y��a	�e0�"9���@��m�x�`��1�ˢc7����7N��9%��4L�k�i�'d
isђL}�<N��v�9���E��P�"}������))�Y�s�{.�
�'��d.�Eߡ������{׿x�l=�u/��q>@f�uX�/B�
ZؒOM�}�7��+C h��~�|RQs�x8 ѕ�V ����#����Ŕ�h�� ��țb�%'�b�/[L��Y���ȗ+=��[��D���c2Ǵ�6W�G.ū��d�SIߣ����%����b�F��Q�m�6\
���m��I�������KF��9*8�!��MA}�F��?Cy���s��U�c���0oa��i��a�����4�R8Ҋ��c�WGij��V0�@��A���S�>�-�� �t}.��n{O�x@�l���2� �8u����4Ql�䕒r���ŸI`���U��a�zx�@�V3E
qIz���ig5K��qb�E��1�>��_�V{ h�	։q��99�_e��9-'��Sh�i�u[Ͱ��))6P��������&�8#��>~�� �J*.<t���q#o�O�{��8׊}�(Ւ���0c��R�/�p�\�i��P��U��ds/Ŧ�]�227lm�	���:I�e�B09�]�;h��m�z���C���tRn\)TW���W�+�<f ��ْ���b�uW�� �t#)A��O+6pi!�d������@�kZ:�(y���y�.��R���Kn�
�T.P����!�8fT_��լ!���2��"��3�YE[�myӉ<l�k�P}8$i��N>��Jv�$�lXͽu*��}��|�s��{��  ����E8���"�%`��{��N-��'��!�3�Q�F�u�������Р����]6A�a�!b�:���֒��;�c�ό����}4(���S���OZ�x/����;��xK�9kBD��dE��y�t�-��d�F������I2Ge+,���[���W�C#�ϩ�ZR���4���c ��s��DFZ�&9|��u;Ap,ߑ`�l�
�5B���T��7#�f����!0Y�#�c���3��q�����	'"��S�Ç82�U�d�[���_��S���:�Ed�I��|ѧ�GU=�7Қp�BUA��x�@��^s\d�Gp���%_\�R�W��J��L���������գ��R(u�D�����Pۡ�@�J@G����jE���S�b��q�}�����P�AC�7�:qOk�t���Mh��(Z#���˩�+�w=,�ay�Z��~��\K;hJ����J\.x��r��šTU�anl��o)a\nId/��s��`	�z;$��3��u��΀X^��<�!�LH��d�Z?G�+���o��F���w��%o/� �L�	�n�R��m�a������F�<�F�n��1�v\�9�Wj�q�{�c�����ʶ��m���Ly���?�t3�vv��n���*�����G>�3p�[�(�N���9=}~6̅S7E{������7Ȏ����!re���_gm�B1-���<׆�xN 6�[wSj��9JL�CN��G�����|�)wj�&���v�%�v*AidO�.B=��(@�K�`O;�Yȗ�,W����%ZGomG�:I�����c̆��@�H��Ux�ys)̔I���*W�WI�hj�Zo� �fR�uwyJ����CS6��LQ8�y���\/�5-ꩅ$ugkI#���.X������ζ��/���}���
��%�^�<xk��+Bm�XۑK/��A��מW-ČV���BϮY���f_�MZhL?Z���27�
��4h�w�����U���Y�%_���L �Cr�r9�N��Y΋K"T�,9��Y�6>̩�����"�O��!{���4�8QW�$�գ�5��2L����
�ޣ�l���W3�*i�BX�w�k~iEyj�3?����y�'j��(�[Α5�2s�<��GL�$~�k�����n��,9�YTf�l2A���CU���H��/<�"AYŐ��q㙵��*����oK�Gk����L,)�;���US��. ��:�� I~|�`�W0*�/7��h՘��sP��5
%��|�,�}�RtU����ކ��|�nN��s�1�u�f�RtP�3&�.c��<ܵC�2���7��%�7�݋|n@eH7_�pV�ٙ��i3���Q\�YŐs���������tS<T8�c����:���PD�(	���^�R�Mc[�TE-1j5q���{YT3}�+�Q��� ?MR#��'J����!��v���2B�EҴl��2�Q���
^�wj��gD�y�c�+�F�sk���`P`�4���o׈��c}�m%5m�T�a<&Q������|�f���*�W����R�c!��1]Qe�^�p��հ�!��ZdR���~�lOd�Rgx:�x��y$}z��l��z���Q9~QO0،Q�lu%~d7���I��|���h4�I�+���G�L����H����{��`��7:�3�A��6�.��W�P��(3b����ɿ2�W⍣M�R��:��(l�1�ɧ�T3~�`\�feGN<����X�B�ꌥ� ���9!4G;�y悝��i�xɝ�J�Z������5�;��T��z���"n�()4v-�j��d�S�����:ރR���g��?q#�Z��c���5�6&�(��*V�"�1��3�yY���2�kHq!�r6�ّ{�Pz-���k'����?�QK��.:�-e�:�