��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzG&jI�#�aW������r�zj�P��)�'�S�s�D��m�PG�d��?��PJ_d��BTD͞��2�I��#�)�X�an�!`��sc�ɵ��P;����OP����-��C �q��y�!N����J�Q5��Mpz�_��xջ�6�y|D��uDG9聱*��Va8�~���#�*t����h����!düF����
��S�~]cDD��yDq��+�p�YA��χ'"Y��"�!�	���l+h�ϐ�gk@T-�߱t	��J��:��m?���/�<�
����O����\��ԈL�1k�S�+L;w���J��;�WA�������Z��q���)rl��R%)����X�՜��J�+n�C[�am �Z�45�n!M�̷5�('� ����ٿع[���μH/X@�\��w��M5�S'�{�Npe<&B���0q�Bʬ�T�N��us�	.���Cߪ��>G���|�4�Os0�!?��~�"���Ӥ�d��Ig�"+�`���z�ӹ��OudLv��$�S@��>�x[��~L�@�l����I�*
K)����s̳�<*|����gb���f��v|!|`]���~�A��o"��?~�[3[4
h`rF��+�B]��s����,�	<E�] [t�eL
���9���j���Ί\�L0Q�d��eS'��k�.`?l�b�{c��Y����j�jެ�n9q�|�(<�d�D	u�-'��~���mw��sçB#ԟh��Pvs�J��V�ɻ�u��/���V)��S�����fq���ϟ[��P�lZ%�0����~�r�"�	�m�Y�Y��FKџ���d��1l2�9Қ[��D$O�����5f
�|*x�p��¶�ix��}�&��ݖ�x!Uɤ�-�S�ǿ�2�����L��+oZ��Zq�*3��Y.�3����/=��U�z���ѣ]�����^�+a�(jWQ��^zj���J*��7�y4���/�(�/�C�|��rI���)ܡ9���gEޏ^d�N��o7?���������KJ^�b�-�5�B���,�\�p�V�;�p�W\c���<�Y��OZ�N��/�z]����є�~��&���ӹ`9V�o���� p�g�D�j�$,"㗊.��_(�)��c�1�J5;��cg��ZY��З0���A&�.��=�����ʕ����>rl9�J�I�umI��	 B��;�ӬA�=��F��kJ�w���$�?�g�j4�D�C�c����Q-���YC��I��6u>�� ��<�Q#���O8��)�؄s�£�Eb��9ȡn�H64g� �	��'��̐r/#�qa��{uOAǲ��/i�ϖG��G�r7>�Bġ?}H�n{4���W�z �5��}8�CgIJ��1[W�����'Y�>跘OYy!����T��qZ� �/J2S�V��IR�̂�7�>�T~fb�F���GBm:�2�+��5��߽�8@^���/M�Cz��������\��u�l���I���7#��.D��]��FgT��ی��C_sδ�X�h\���:�dŋY.FW��v/:r����|�V}�"����+�ѣw�`���3{"ww�����z�o_J��L0�Ć����\o���r��vF�)�)3�)�HI�Fs����^��_�`g������:�s%�w�:�|�E�^�:R�WU�{.����l�>�Pަ	uxCˈӸ��׾�UO�H��?hG���=c���_K��{XM����6��<[>0�)�1$�r���YG������/�<&3�&̧�L4٨<�3�ᙳ�\imۋIK���̏w�*�'��k��%�eN�Vz��;��-ld:�>/��
�T��FG�*�|$��R�����#���;1�$��c(ɉ��_Kw�3sRV#����UK�q������b�r:#�S��é��è��r։Ӽp0X&����6f���
�*�:&.�f=���# ���Q��"�9���n�>�:]�3�%H@��1(��*�e�~�����v5�٘|#E�e�4�>�L��^&��q��%��џ�_`k\��f�+�??nppd�[fP�:�(Կj%��;�\��V� �Ay�;e a���^z���X���q&�V��[:`Z�]�*>#�-ۨ�k�sC,�~&�3�mSD��ɵ����\