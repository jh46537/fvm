��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���Ox���0��?T�}�D�yBl98�锛�l	`�ġ	d}�:��PƸ����~��R��o�K�jV�,R����vy���3����O���Z�����g�̼A��v�{�7
��5�¾����B�C����������r}�:ش)qqa���·����BW�4����"V�CL�zhXo�e��6kT]xl(���%lT'�W���'�N�V#�L�`�`�Xy�6$���:��9I��ì=P��uS�I�w��������F��<��s��y�i�u�����ml�G")�O�4����}�,r��𯴢}�鑪 _@�y�Tkt}��8!�JŜ�>9��C �gl���-����{���Z�*� 9�[�B���c�M�͠�+�G�Yy"TGz_'l��2/;��	^F�/	b2�ܕ�Z���./k7iǶ�>��R nS�}O�i|�y��|N��yJ\
�U#xi��|爫m^��I��6 �!�Qڔ"	�Yj���+��!�k}4�q5�0�:O�1�.M�ϹW>e+.���/�	M�;�P�R�K~Ea� }�]B+ �� !E�N:�x>�@[�s��4 .���>4��G�ڒ�b��9�����o�H�6�5�ާL�,B�
��ϴ�sL�/�Q?+���eƗ�:W�ML��0bc��R�Z�%��#�?g0tndٵoQ� ��U�z��`�T=�[�z�J����������\I�ZB)Lh�Cۘ�_v~J�_��}�����^c��cSb-��ae���U���29��l��U:���舛1��6���S6�����3��q(���Z��a}�ί����H��
Ա3.XV�(L���~/xG<�3���n���bԠ��Sl.�����^��F��ʢ\j^��N�8|DX"��'㏽��T��/9�ysӴ
�%�Ev��oI����G���J�!i�d�P�lZ�ޔv[�����-~�Ub������g�m\E���i��E�׈@�8m��T৽��8W������%�)
�![�:���%YD�UV&��Ա�����;v%}E�h�(���!�S�#��4�g�\WD6�Z�]��ɎZ��jsFnqF�tvHE}n:1�����b�P;M4�:�У��r;7��ک��|�<��:RM��������`�k�Ƀ�ܸT꾴X�-1���an�L�_�#/if"[$��]��ʆ[iT�[.��ԭiTٔ٠Κl���X��Z};�]�}4TSƉ�,>/~�i[���yL,��c��2"�
�h&��f� x�yJ��f�!)Y5�s�S6������F���UO�U���
a��16\;��3�O����C�٧%��\�>��H�,���܁kׅ7C9
�i;��ctq�i�I�'��'�R�]��N�����Ǖ���a{$NQ۠"����w�9Xtn4a��#z�d|C@����CѕM����M�?� �\�3h}�a��/�x����(��j�bfJ]�B<�s��_��ԁܭNўK+h��䪭0�/p�`���I�G��b��
G�͒����Yf-"��"T�9�l�h�����>��;���䤾�� �,����Fc~����;��.��� ��7=��ր�pz^�GU"����	�;a'?�֎p���ߒ�¼*��x���vwn�^�k�U��uJC�I`�����R&x�..ۙ2�#V��t��Ni�����n�(mg|��1y�=��:��@�/4�k�$v��y��NpmxR��2z�.�Z�,���>䥀�	�\\�u��v�{\*��:+K�*]�����v��~H�^���GɁ}k"����W�c�X�Vv�ע��_duR�K��8�Ϝ�+�=O�eR�^�Y��h��L�iP���<^��<B �������{��'g�<�|;Q�3ܺ�N7Z�X� }7�p��jl��N��|����ϕ� %jz�^��^��=1�KkL�~�--C��0[3jO�`l'����q3�HQNz���a8SD8�}����X_\��*>�ʸϩV'�,e@�[\���UE�~]wވ��t=�!�o��O����b/`q5�>��Ci��P�����H��j�G2��h�r��lQ��MHe�[o:�ſ-�~~��Lh�1Ǚ~-��KX���w�s�.���E�KF��Ԉމ
�'��<(�����/Bi��M3��z��{t��������O�ș  �����!�����$��}��z�Fi�P��J���Y%�(�9�����B��wr'��L�N�x�7�Z�-S��S��%�2^&م��.�0�%�����5Ǒ�^�� �����c�6P��2dPƠ=��c3��"/eu�ťl����<H[��`7#r.����w��"���'���(o���R#'ܱ���@)�S��l`Q��P�)ڭpR�����\>i���3i�!�U�{���ŝ�Q��Ï�-�D�
�MP����ͅ*�!���$�aJ�j�P�& 8ʼ.��2#()��١��3֩vE2ʄeݤE,3?b��w�pi�8�߾�Gσ<����9l�GccۘTS�J�H>��[��g�Z�ۘ�f?��n��A�����zO�nr�5����²1��7�[�"��$��e�������l'oMϪz�T���J�g��"(��X�������JB�]`+L�As��%���T���k<�ZC�gK���`)�b��K;84��-x%�������[�{�W�:�v�C�����Z����B��+��)攰 �ARZ�e�=씐A����Vg�_�A��>xy�%���q��R�*G�.i��d��i26�N~Yaf%�ԕĩ�5��f�~�`w��i��,-$ȾВ�ZM&>L��0$������\=��*���A�`H����ԫ����e�1���l��y:[ѕT1m��ߵ2�i��x�Z_��,m������oT(_����!�̿[��l�^"{bN/n�j�����~l�k��>�&�l�;l��"�c{C�`��c����-������f	���G��4.�ch�[G+Ю;`���&�̂
��I$x����)��H�g:^�G�B`��'g �aaj����D���nV��|Z���90��۪=ԚJ��j�.�^�a�/�⇹�@�X��Yq�,8�ͮ%-�نt�fwͬ����ŝ�ى���8�to���Eɹ�����R!��Gx������l�%��ga���á�}k_��C���Ǎ���v�+'r	���}�;�~|��f�qfuGz[ ����,R����޴��ܲ�1F��AQ�/��2l�Xú��R�F�&�n��X�\wҍض�Eq�^{Bv�:��9.iuqw֎�q*%	�ad�$�,ST��k����=1��/���U�'Z��@b�v��A9�����Ij(��WE�>�mȰ.�����֥Qw&���V�����j�%1V�=o%E쒘E��6�$��1�̰�ڀ��k�|��8C���jI6'�x�&HlP2��ԗ��>��;}���دM�nnAZzN�F�1S��΃��~��m7(c�V�xY��T�E�	��nU2Ã3��ٓ��G�K=88���6<��H�.u�a���l��A�F�-�J�`�m=c��O�0�/��PVQ�e��(���l����Y܏�u��7�3Z�4N���2N`�f�Q�dh���e��pұ�fE�)���@a�R�����%�Uj�v<���
��DM��Mu��t]�r��~��#GpL����t��Y5���׫��>���a�6WIO]P4�}3�ДI��ItO��8W��<��UuV�#ShE�0hȱj�jq+0����q��e��qan�3�1A�j�]�ѕc��f�� 7�鐿��ZI��]Ln>m�UHq �K�����Q]�\߉�\�(ɋ@��<}3�jJ�^�=�j3�2��c���dT��[GM�.&���n�V�Z<��{�-2)Nk�v���@����1G�1B&<��=L*��7����l���0^`�h?9�Y�4��%���Z��W�S��Y�I��a��Yu�d �:�^�BeK-��t�jG��+���#�sl�:6���~y�°�qơ�S5FK�o�u�tͶp���N�$���I
 �v?9��F�o�����p�d��QO �S���YK����\�Us����/ԣ���)��V����~tZ�[��MUP@�v𮐘�>$�9$5
�tiv��,_�U��'��p�89�&�0�c�L7Ѿ�����<f��ϼ�"���Ӥ�XlǴ�!��I�k�_��*�$�]��c���qK�����3-|wB���" ��0P�y��@h��Bucy�Sw�ku�����8����c��݄���Tk6�%�Ď0:ŏ�%��n�,n�������8�ǹ�TH��i^�bi���9ꨛ)u�m���Mj�.h{ �l$ߢ~�>�:%l���J�?���@����:�^ec�?|�չY�v�����f�@�˻
�QT4�և?�+;����Yء���h�?E-M�o�)�-ڢhP��gy��e�v�*���O�d؎M!�+hw��)��C�/���>�pF]�D:4����r�o��&܏%e�֏IM'Zhv@-�vy���1+ƽ0�f�2�R[c�.EX�g� r�!��2�_	:�a��L��q�k����l�iS:��m~��B���JSkZ�Oˊq�}�wx�S��K��Yi�����L C\����~Y���f��NB�ʛ��#��m�d�8Q���(��L��h� ����Q���4ؾ,�W�.�k�F�B�u�eH����d(S�?��%qL�q��処��dģdeƉ+�RiL~�$pL	6�T�x~��Й1f���t΢�-`^����c�Vͪ�v�� �D	<3�y��w����x�#a�;�W�|R �L�+�((�P�s�4����[���ұ��r�cof�]��'�CS%�l�[@5'����Gj�����AQ��b�{���c�w�t�ֱW�#�K3?A�Ӟw*<jCu�жrqY?I/ID���ל2�QU�CE���_N�MŊm4�Ʒz��'n�k�IA� ��pd$�0a�[jڵڸ�xIE�Ɂ�l}�̡���`�"�X�]���G��Dչ��E��	R4���'K�[��X����M�؉7ˈ
]�pǨ}�-�N�A\��Fp}��O��E�ڨ�+�0,|�%�Y��
�r�зr������ tI����9:�Q��
H�p�=����iAY�����엸�ji�2@!p�)QH���hE��&u��&��m�A�y\��L�#룗;Fø$i+�,q��;��`�ŅXc��rI̦5/�w������$��֊�=�B��rY& �Oy���b�va�z�#Y�䳱Yv`"���R�!!I/Q�2�$.��w��~F�Sa���� ����
3��0:+�n.�ߦ.r?������3��}���3cMTb�h���OA����'��՝�x�������;���Mo�F����L���{7�vg9����hd�?�&鴸�K�{��-!1"�*������yAQӔ��[E��:EXCx=�F�5�t�}Ҳ�ЩK�Mv/1^��O�������qv�jgG��7�W��;Dk�vG���8@K�_^���*t||�~}�@��Zrd��R�}T�/��r�C��ɛ�W+a��z����y`#��)xfD�!/�̳*+������\��J�0K�1Jʓ֣򗝮���{L�����8^���K-�P��䒻3�|	7���ԃ�LU�D�RŞ���22w.�P2�KP� ����ް�,JZ��	�V{͛�������9+����Xߩ��-��g�_�g�~%���jl�3?b��F;V���(�,/�f�2}�^��d�T��:�aW�7�l2r�AzӅ�cZn~��Y�j�gE����	j��M��Z���BQi@/�=3�����ɖE�/���	2�(@|����
QrH5�u����ґM�d��Z(�q4��C��x��>��չ�`� �[����Kޱ�_�4 �T;���g�}H�ʲE�}�:�/H�8��l���P�
�S�ˆN�� ���5k){.+��O��l��Qq)0�2�k_]PP��ӵ�b�v
$Y�����xe����hF+��WR4��Oít���x�W��呟V~{q�Y�|���d��^���v��8�+�')�`1��~2x;���7��x}��@��x��͚��|��׽���D}����~�0��=��kG��E�43�6;G!��9���Y���,�:Z*}���Mf�l�
��b�]��n�BA��J�t��-Z����6�#�q臅[���ʜg���Q|�/�_����4�e}��	���r�!����V�Y��O��]d���������^1�;���G�%�6���>^؉�T]�E'D��txu��s�S�֣ڮ��Odp�Zi�	6�ɒ&�����hX�1��P�9�F�d�֯9L�J�_��1���ڔ��")�����x�t�����؁K5:���I��#^`I�v����9
�g]��A��5Z��C~dIћ,��9|8Ơ�4��H��(���=*c�`M�KW.�3���I��m��,{M���7�������1�l��p�� ˷�1�d����k�+2V(���"f�<#DK�����eO
Vʅ{6$��i7��E�ñ(��vH���f	����Ml�4�1L/!N�\ۚ��+�3��<��,��%�������S�1Hkd�+8�џ��=�>�ƀj ��h�a`��È���I��;1ds���8>�QQ�Fi�}���4��ۅ4D��ʩe�;w�F�J��V�5�#��@�;�ϲ�#�e�d�	��_�U��ޗOyV �Z�x��ſ�����-�t�/�!��{�p���X�1ݱw�j	F�֧�9`$gh_�d3��	i��~�cM%f����$]���c����|�L�8՜�e�^�,Y��}nϸ	�as@}�_MP���M�-�����q��hK̳�X��H�c�+Q��B�b0���
��x<�͠��Ѫ����¼P�i:H-Q�<⬗��u�Koqp۝���6�qt|T���~�!:���ZT�m~�������u���V�%U�|i3jkq���)mP���áט��1�~Wc^�q�EL3RuL�������+�;�{8��������B5tv}A&i��ʒ��������"��9��e@]Z�̤�?�K$�1����W��E8@��K���!�2B��K�%��wNឧ��i%�b����s]G#������cun浠���S�L}q��rT5h���aV_��.�}�۹�Ԡ�nPM}���L�����VӚ��x�#�D��|�#=��=lhR)P���X�E��]ö�c�o[�l��+A�n��U?W�׉v-�S�؊ߘDN�l�Or��Z��z�zl�����Y��1M:^�;�r���K�sM����1���{���d@��|T�)��@�áu�4�B�bB���(�F&��.��@E}cI%%�� ��}��+���7���k	��B�;yy�֊�2�� ��i�dƧ� ���=(i�/�{�������`S�����߄�ٍY޳v�M����]��{e6N#8Q�u+���B"+h�Ϳ��	�j�>��.@X_�M��Y�=��w�6s|�/*v��}co��'8(����p���