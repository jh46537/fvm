��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��At�JD��>�dtW����.��E�?8~ƣ�8������k 8SE��O��������9�����џ��W����oUdf��ߣ,E���M���F z2�ѩK�	����b<��Qy"V8�2*X{5�MG^v���^�2ON��[Wg�ow����q���?�\�P�����s�N	}��������0w_�ٝ�L��S"�ri�6r�ħ��!�|�0�S���p6�c�p� ;�I~�6(B��6��� D���\��ue�\��� ����_Mp�HӧE�`ǫ��#E��o qa�$������`��VIS}q=kr��ɢ������e���T��#�"� ���5志�ͅ�
簄�]"��DZ�8�ݺ�jh^c&��Gֽ'D>�� �`��@~#:��D�8>f&mCi{֥+��'�$5������`���'��L$N��"���)d�r�!�=N���N<����9:Qt��*c\�h�$��\�D�(YX�~�7.#<\�S�_o<�Æ_��R�v҄.5���m:P��W��X�ɾ��.#���b=	��hq����xK-k��x��)�j�&������To�$���t�U��~�{�=y�
�반j�
�|�4[��`���)Q����RK��F�����.�M%,9�qU�y�,Z�(p���=W�G�B$q�i|}γ׉A���Է/w7����lm�'����!��8�<�A�ܪ9PЮMjf_=g�R��o�6��Wu������Wd&KȔ�ܹ}�64�#�H����	�c�N��TaG@l5�ʬ��������ޑ�����\��5 �~�=%W{j�p#���2Y�93;���C)����6>7��/3��xp	�b�ی����M3\�IK���Dt���ڝ�c$���Oh�U��8m&$q�����:�(�������+,���Qx�b�)k���
M+R�8'<ď��_'����NrX�fYn��7�u~HqqV�\&�����:�C�S�N�49	b���q��c��z�$�g�s�
�
nf����p�3���ae����w������q窵wtÑٙ����T�[W]P'��Y��5F�l!8��`���j�'���Q�w��wV.t!� lZ�~��lr��x4
����"^3(+v��c���m إ�T���줰#\�J0�%.�	v���5���$����� �`�~v�[��#��wO78��v�za��E�ٹ�����{���-(�V"*�`q�'�����/f#�C~%�L�G��%�;E�@۽�Cu����}����0J��7�$�=R�̹�jƀ�
os5��ᯪ�Op�r�tg��X�UBZ�&	b���&*�s��o�*h�5r����s(㍕k;J��7d�x�>R��3C܉�Bv�#����]�!y�Ͻ�BjΗ:ﮓ��s�]�#���A���fKY*E�c��[B�E�Vr�-� E����1ɏ�o�o��Ř{͝t��9�Ƞa�,��s5�D)u���[f��WV�":�1�����Z��� ^@_���fq5�!	�I��
�J���S�6�	q ���u/�ljQ�O�\!���g�*oM�)72?p��WΥ�@*6�����Ʌb�/&��,���W�d�g��)o;����4�l���Z�#Bp�ŝ�Z�[�]����s�!�ळ4�@��k6�{B��VӲk�a��͇#F����ˎ0+�#�.���=,.�O�M���[��*������-8b�gy�P����a��+N���R�}��z��D �y�M���S���\��IH�x&��Xq���5����SX�ݎ��ASd[uY�<����o�\R����~s���<k��j|�m�������d��2C�<BZ
L#-�B�_17���Tθ�3T����*���ْ���[>�@,ߟ �Mt-񯜄��f5){�e���4�}�8ǲ?��] ���w"��m
�����v��m� ��������I�"Z�	����1`��D�z�94-7�o�iE^I]g�i�m9J�Y����-���x.d���-*e){�<�|��I�#�G-�����i�7Ĕz��!A�~��Cǘ�/���<��r�C^�S��R�K�:2Q-�Qm��S9FK�.侞��	��RW����a#)��N������45Ӡ�X�;����/��2p��?}����8@O���0�#��zؓG`zD	x�a~ړhEȃ^�pn�9s���n(��V�>7�A��u�A/��7l����[��u�f]
�(́�Ʒ�?R�ݜ	|��S�GR��Ҭ�E}x��b�'��_
��Jb&��}�r�
�g(����	,Ӯ����Xu�Pm0nQu��#����yBR~�3f�t׫�5������s��qj�,@'��WU�J���mU�8&�̘@ ���,B֤Bwo��` �C#�e�P(-%v�P�o�b��E� ]�dǵ���M$Ze8Ke:�oՁ�}���� �QR���g�e��a�K�4B�ld�&��:M�Pr��u��q��V-G���s�Wc]�ᴆ� ]��欏Ӈ�l!�>�Fї+�H: ��. ����\Ө�)aK�P�����_�2:"�*������4��b�t
4O�b4�����pf�I<�b��E?���CYC��J�Ʀ��0QsT���}�e�Zqi_��U��ORڈ�^ C�ɣ��	q�_�^7ٍ_�ּ;W��JGK��e�P|{'3�$�,E{5�[�ʛiW}\�Gٔϟ������9ǖɯ(�y���`�g2�Y����C�w�t
i�ͰB��a�6�.:]Ot�pj]ڝ�R�u-����yQ*�}�"�%?E+72r3�AX�$� �?�+gj��'K��u������,�P��ε�SKW�;<�L!zb}1�+Я`���j��2�fF�Y��ʁ��@V��yT9�p����!���<4�S{k �[E{�#�B�2��%Q�۝����h�~S%	{	�e���5���~��4_�Ъ���
 s�����E��vʻ�@E��6���}QXA��z��3�L3�LB��gjv��أPi�si�ף�&u���ZX�%0x����� ����%pr+��쥥W�u�1(q_����~Y����u��e�������/>\]�*̈9F�o�7wk�H�J	��˳���n���#ڑ� *о���&�v���7��v�d�^q���K_z�����g߹�.�pJ'l�5�� H ���j@n�,ݕ�űOq`��ٗ�@Z��e�?��@ZB���Z1�?�bu�}ɜ/��'�EzLK�_�7ju@�Ǆ���"�y-߾��nq�Bݹ��7d�f)�a�R���OOi*����g��0��Z)K�Gs32���L�6:�*�B&���}�R3��}G�'x��iY��<��M'a?9��_���,ME�j���������A��#B�A#���`��֗�桖q���C�N��ݵRN���t�G��� ��V^%Xξ��c�Dsf�-V樬���qnJ�+�S����G��O��)Hu|� `��.H,%��3!&ӿp��f����u1����CLXQq#�
�(��BG���L8� ��H�V��Xe�[D/�����]�{��
E8<�����M�w�a�u�����g7f����g�Zt�a��
	.��U�e��z\հ�|?ꞎ����5��}�2�YA�3×?��a�������/��r�{������ �e9�	[��O+��j�� Qeb��AM����fM��g��;l�����4�\�~���تjA{�̣�5P�`]�z� �'���5��F��QG%n�uz � [Q�Kz=q6` #6�N�6��v�'Կ��Kk�(ׯș(;Ԯ���uBUv��]�ɰف�X~������z��CO��F��Dt�4Yz�B���ŷi�{爗��������e�[��3����G��o��{�Z䝾���}��pkS餃Ӻ�77�p�@F�=����Ykz������8�G 8�N�|Z�q���`���Z!yH�D���a�&�C�Nu���Y"��; �b���z/� �J��_v���r�E�ׅ߫w����b篏�[%c���׏���xg�a����nKp���j������mM�����񦊾8	=�*"~}��#��e�Uc��ǘ�4m_��^��ʧ�P�EQr�U�旣#���5AB��X�H�w��xm2�'�F���s�3�L��S=]T��9La�(N��ѓqNs�x_�U]�K*[����M���B)�ݐ�Gh���2X��qI�y»�)�$
k������
(��͊-��C��nz��^q}]n���@���##�ח4>�/+������u<RP��f������ɫ�C�
ʲ� �[�j�����}+�G٭�ꯣ��Ҵ�Jz�TkM*���)4�*7��5>wv��zG��t��jbPO� ���f�?~�~T{��J��.�W���
;9 �I��߆A;�����Bi�E�&���|�V����|�3��<+ݴM׼J��2q�.���+��p�wE���|t�
�v���Wr����z�j��9�P���QQ���ig y�j���.�!�/r�