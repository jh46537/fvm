��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����G��l��"�Fe]=�/>�"�3Nع}EJ0���U4�q��q��i��[�3W9^�LU�3k<�ҋ�͙.$w{�d#?ŧ�.�&���\�FaAG��Ƚ6�o�� ~[Z���~s��c!��ء���]N;k����h ���ZAcd�q�4S3�*S���k�!�[�>�Gf����tZf�ث���Ta�z;TcP�.�Dz�Wt�'�KC���h�����D�����5G�j~7���w�q]M�����u��ɲ�9�#���ƈBt�L�Q1.q4���v{��і��гX��"K��8Z!żD T/�P��x^�அ�#�U8Kr�%��;�:�o*ΧքF�K���.�cۇD������,Ih�w�qf���}f�iq��N�AΕ�H�����[_&�Xa�!^䆎����VV$��e=ۈ�4s���&	Ψ����QI�_�ZO{�a#K��<�2#�큚u�E:�y�n�%t��I_J�h�T�m��.�34Gږ�:'unZOЫJ���*�z	�:S�'��[=�����󷽠��B�a/T>Cs}�����b&��9u@'e�6 �,>ݧI�aA�S[��\����[��6�JZ)Ӓ��ɒ�=5O� ��w+*�8��-�o�! �l�n(.gnX����G�$����(�I�_9�{�iL��tV<�0�.�8��\6�L~�;�8��;�6#�J�[bY�y�;�r���Hd#����x4 ������aޛa�?;��3�\�]�����Gu@|�vj��,<W:�:o��pT�L�����ùy���� n��6�`�<Ȕ�>'ˊ(��P�?cuL��r��I ��F
0�T�:�{`�9���{3�˵���[�Oۿ�h�7�fth������*���ǌʀ"pr�WB>�'����j'vE.玧���!Ƙޠ�AΟ�>r�gEo/���;6���u0́�&w�n	��\�uK���ה�9x��� s���;eJdAW�Zz<�����x�z��2cn���"|�����E�;���~P�0�1ZGI@���aŵ�LϢ�@�j�n�!��.n'��.+"q�o���rf��R\*�՛