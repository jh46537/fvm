��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��V-�@m��Yx�W����A�.�ƋB8/dq�4z
�2z���,�k�������^�	���/��O�pf��$���:�!� h����-�
+�pe�$"���𝘹�qT1��)�*�8���|��&�U��.(vJ���?�2E_d�S�S��g�m�6����J�]�G�6<���{�rNř@��A��)�Z=?>��fV-}�
�T2����?���.�����ٷ��u������|�
]���b�V̎& �Af�v���ĕ����UHU�w̲���
�<	[{ssxa�Y.:�r��54c��0)�t�z�u�XL�JK��_�z]�X�
���J�ZaG�,�|ię��Ѿ@�N,������e�"�2}&4p�8]NՏR��e�F��/��+�_�)=��U2})7�=�`�vr��T��(	�\X��p�p��1�7�*��hv;}���(o��ۄ��o�|�+�a,�%�.$�
�U �L��6X��ݷ���n�k[�=\�e�F�/U V1߃�Z�
9�Pç�JEG9�{��MJvX���&�cݷ�\��X;K����<�P"�Αgw���i��J��~��0v���5#*f�����s��Rk�vOP���ø�j1b`�T�C���IZܼ�%�)6Y��h)��, �W��)�0�=`+V㎗���(��T��>�*-�d< �ݴ�<�A�Ek�,��L�(VGnAc�Lʲ԰ƅ��
9�ȉ2���No�̵v��"�~�~ނ����c������G������Ht5���:����T�j���7EdEi��6�;>��0�*��O:��MG�hu0'��x���`}���f ��gЌ�/|�dV0�N??Ͷ�"�=P�\�{Qh �����|#��������Os⦅��ne�:<�9��8*��:A������ �f^�nQ�QK#��O/V�׷����q���m��2��f��i�6����'2�.���ݎ�=S��?֠S9g�e��j��!xf��t������Φ�*�9)�oqɴc�HZn�v�,>�J��`]��ǒ�.f-�0�5��7#�Y�3@��L^����"+0Vk@c��/� ��g���l��qgMWpsqQ'��k��dٹ�����*V Ѷz:��F'��q�����1��Ń���~R�1�q�f���c)cG���A�y��w��,�!��[C�9�����'Kug���
���sN=�A�N�a�U���is�.h^W�*y�ج���%��� �v�:U%/�4��I�A�,�@�~7˃�q�j�4M�D	��Q������+��E6�W��n���.����j$4�:S��xʻ�/'��S�@�=�� ��.+m3�����@ �rvUr#�G�)]l\'��O�ѻR�;��wj&��IN��q/��WV�D���b��`�Zl��`�O/��5�s..�9��P��~�+m�~�
lT)P��N�TW�`Qs�����Ӯ�!㱲̊W-�2�(`,��ӳ�$K�/Y�!(Ydۘz� E�u6j��I3L�s��0esNl��N����:ZЩ+9�j�s��ۓ��ew����>�;��}�w�i��x0�
���-ë$���`E2��k�V�����]v��mTq��j��$a6!�ቋT\d��1:h*T���_��}���A@&�\Nք9��L��� ��v����Y�t��C�����H�v�l���D�$���Tu�%Z�o,�����<9��碎#FS�Z'�;̓�*]m��V-�#Y��+v{�ێ'��'�U'Q�c�/0=�r��ߟ܋]��~l'-�n�L�#�F=���Ut>�����є]��]	C�D�����&�g��}��b���#^�I����Pps�	�t� (������7���"b��\��cr9�2ȩ%@Y�JN�8���Ѻ�r��������Rt�V�I�e�F@�e����
8Z��z=z��r(����V��$���⒣\�M�������N��XѫԄZ�$�g���bn���ԧ��,r2`����n�T��3��P�6C$��}jϘ@�'�τP�ܚr�Q����C�F��qX�5D	�Q��N�%���`E}śԦ1;
8���� +i=��_֭�ޜf���&
I|����!@��4��L ����R�����>�D@AK��ъ�n�����g؀�Ի-1�tnc�:�����5!�	�����i_��Ђ�c�z�w��ӈ-	�� �[���TR<�"ȉ/R�k�)~�gf�� �
]�䢌����XS��=U��i�zрw�G����	l�]�@��;�8�?�k=�ŷ3;f�qZ�b��U�񉋊w)�V0-a%XAYf[�η�L�0���)�B˴�w)��䲪#R�H�0��v.Ss����nŢ����O����רu@;�x��:�䎰~ܕ�ƽ+|9�32��&��"ׂi���mHo=I����c�c�b���R��p�b�Fu���`�p�
1g>�����ͽ�c`�9�� {��bǧM�8�&�(��^�"oVm@Wg��
�ro�h�`�S'k�� j�Y��]�����8�-��o�ͳ�Z�hƥ� �Y5��X��%�M�hrػ��	|a�U
XZaO[�"���u������S�L�T�����B�vݻĨ�d�߮�n3b)�Q�\#BG%�Q�=p;��ۆ3�/��
�s���de�rm���D�^�^�?�# 
�^Z���&nFr��0>��j�k0v�*ٲ�>�����2?Gݽ)�4�'"b�b
î¿���tB���yCx�k��٩��,eex?C��o�z���xX�JH`�8/�7[4-�o-X�u��l��sR<s��!��r�9��b�`4�aͮc�LW�T΂^���8�|_P�:| ��d�E9 ����?��6�tQ�T����N����o�{������E��U�*�eQeh�5�G$Bx&B���*�� ?�Q���g0<2�Y��W��#cD��U��"W�h��ؖu�(���)Ԇ���y��Y��K��=�^�׀�Ś[�\�K���X�:�7IU�v�C���?�o�.?QW m�-��BN���fĘ^�����4;�����@0O�u�Z�svdm6儢/�@�$��`)1��]r/�?s�B9}�"M�_~Hʃ��|HaF3��b�M��ȽGYV9���q��G�r%n�7��ƌ��Ztxu�8�O�op�%�T�˾�_�\�g'AZW�����������c�_���3�-Q@ "��Ib�ߧ���q��nR�Γ���{V�y��x���쯅�_G˓T[�����l��C�2����&1�y0�c� e(�Txg6��J6�A��l�b_�,�K��4[�����r�4����Ƀ�
�7ꞥ������BPpdBXm���vԪNt��^���gG9�d�����I&[����l��� �u�M����خ�I1��h����ZU����_<�$�h{j�����	�M���s��-�1�EE�I
v�ZlBkp��$.Z��Lw$��J�J���-&ĭ=��2�K8�y�K$�T\���w�c��������Q.�.��L�:��;[�s�"���DC���<�)���������c�XJ���;s���Km������L�G�b]�������&0ѩ8�u	��S���K�[��=s��G��a�K9.��z�&v���MRA�YNuFV<G��	�F�\�i��J8ƶ���V����y"7�po�Kd��#mu@�C׹&<�F9>t�p)�[)�2H��S*R�.7�7e���w�@o�� :������/d?(�#Q�	��m���C�$`�(-a޼SC9fu����&�Z<��$Р�	p`C�}u�r6\L������|̩�̏C}�%H�Ex!H�|������-4�J-Y?EСA\6"��o��aO�������~�Zs�����Sn� �.���J ��֎Ʈ��cC�m4�l����V��&!;Z��aJ�F偧:��2��~ :j�)�L��mTS��w����A����W��[�=��$�R!P��w�B�W.��]<��&	�9��.�&�Ƹ.�׫^�3`���
��?>���r�w����/�S(ɣ�Y��r�����o:��A@��㓯FL&�:�ڌ��ԭ�D��8���1��d9k����)!��v�Ky���"-��nZ?� ݤ���YV����"�W�PB��D���2�D��%ra�� �K���, �����G����ܘ��o#8��킬��ƭ��DK����ն�5d��}�r���1'H&�.�,$l����ن���%G2�wc�	]~?��17����$wQ�y���\P2��mН�Q�Wt�'ʮ�ׅy��v��.U������`�0��R�Ik���pN83u\Z���Ύ5��8��y��(v��l{g�Zr�Ɩq\��y����Z �ohk�2tD��R�h�fqg(��]\S~�T:.������P��ч��B�Q�ͅ[s�srQ�����mʘ=�� 8b�:+�C��b0D�ɑ����y����0�W|q�3��n�@�U��W[A����9:���w����P`��^s$�$R���*��ʸft����\��:0K�GQ �(_��P��f�{E`�g� `]���~�cl�-h�M ��%!��?�42O���QN��}�}�bOHӷP9x�Um��T��u��e��?��0핋;�Ji�D۫���3�=�S���d�'�Z�֗�p��V��Xǰ�w��.܊|�Xn�\�"���)��G��*<�}w%��n&	���vXӨ����*���
�Z��^�xJ�mA��U�(��g]�h��r'��7��N���lhG�Tzn��J��p{�������'A�(��W���P����"�ԘK�u��krݙV��������Q��v1R2�Y�[㉽�&�� J��.L���ɘ���/hj�àu7�Ͼ��}׎�y���и7E�M����Y�cdQ˽��=�u��p��G"�p!��Sa��1��������Q�����w�?J��i��c�9�&F~�Y�o�}����u���ly..V�Ce`}b�UX�`��9a�+�?�f�T�c�u/ߕ�����{�����D+��87n��GpJ��~b�H$�-�����)��}1c=u�\6-�L�dW"���T��J��������y��4��ޑ;I�n�h��xr�ѷ�rL��T>��g��Q:K�:���Ia��I	�v���:p2^Z����.�� �?Q�_{���1�D�-��/s1�굯�R��YQ�+٥��w��:�]�4.�A��W�ξo󭖟>]w�L�r����ҒR���<B��N R��p_ߊ4A���fv?�2R�~f�W�w/be�<��KG6
�p�� ���i���^E��/�3�%��[!,���(����v�VA�7$LG�F8u�}�OZZBfTkh��(���S�A7���ǬW����t�[���({1}�|�<��\���1�7R��_���mEWM���D����%i#z�3��xУ
)tc-6ړ�f^��:��<�gsH�6�ӭ�6�t����<����fPM������'������vR˩���E{(���`wu{�v��2m���-�=�W^���1����J'
M���0�՝�⇠5���j'ɭ����OЄ�@X1��r6~�"������+Pi���+�>ZN,*SW�`=��IUj�7�ڤ�NjR��ŨqD�6V�&)(S�C$>��e�5�9��vѐ��-Po�7F�\�w�ߖL�Uc�{!5\��9�""U��#4��E^�z^���vQ-���&e$Q0�v�|γ�Mc,Hߗ�w+u+I�ٷ&9�2��#O������8�^L����/	�
��w����s<֣�����H��X����t�Z��:�Z����O�%K^F�V,���$x��V+�-�I2N�/�\����|X�A�|�G��ש��¬�1�~oE�����٪��K�l��t���3KQf�1E4�
��_�ȣ��E`pd��ڏi*��q���!�t&U�"�zH�M�:��%�\`�UC���/���e��P�Wrj�\���65�%��;ny~g�7?Q!�\��0�|&�W����̴O��K>)qo��z��)�[C3i�=��LY�A�, ��8�����&�ѥW�my�$�z]�r�籠a����#`9Mh���2�SkA̟z�4*�Rz��~�O��A;�7��߯'a�E��~�"q�[9+�w��Ӟ,��"|h��j�2+�C4�������o�}+M�B�v'n"�@#�b/,#������̬����o���ޓ�5i)�/�>*?W�}�L,����?�����i*UA�Ѽ��2
�as
�c�*/~�z�����&��^���?��lj���;�6�y�R�Ѝ���%b��P��u'3�)�7t�� �D�m�}*��M,A�fZ�t��0��_�Z�dͼ[�ur������l�@���޾����6�9/�&�!�5��Mo�l������(��{5���,�+c㗭�"�w�0q�� ����h���k25�՞T�zm
+�H4�q�F�x�L����u�N���r�\��q"{��,[�|O��b���h)��PN1�yD_~��o�7f�����ik�K��n��Ķ��	��ST]܈>�sw��_���;���d_��d!$q���8̑G�$�ham(S��(O1jk8aZ�@cWy�M���[eX�<��%�;;,<�e
�Q�>?)�b��֎=nAe*]}O��T:,e��`�;�m����w�Xo��"���;}��DQܸ� ���7�x��N�A����{@���O��J ��	�ca8i֐"���r�QQ1�r���H�?g嬒��A�J���j�:�M1�Rłr�7�h��2|��$�s��{á2�	���vVG)��~�&���L�%C�ٔ�������#�,����^�Memݼ��Mc׏z��y�1|wTO�b��S�7�}�ۯU���	씕vI�����r���Ƒ��&�Z�l��"ϲ_9����c�+��G�#;·�n