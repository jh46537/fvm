// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sdYOwon60A8kM55GhzhTIv0MMCh3LWAsvKHYgrptC9jwBGOSKWepPn0XSO+COpn/
uFCm/EsTCjaYJg8lyCquEyUIXkTduceiipMfUTTsQailLMqY0q641NdBTzCgK7rP
9cC2OfbnPXdFe4avPQfZXE43tKhth3I+Sm+1sPZbm6M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11712)
JFmQuhpwx2eGk/3w8QUhTPtm6yCKv1DyYFL2nPlqusZNPpW5644REmSiIBw+xFFW
mrOV75emFvUGAMj75i2wQvG3MUtRuPqsqjUrPES2c5iPQxatn07xsS+TfAndasYW
44cmgwwONXLTeoBy2x9dRzpMMpOnzVeccN3/zLtchvH7Bu50zYaWQKH5dOU3xzOD
PL/fTYVsFAfLQ7oGAIV409VxDSYXX3Eog65xHswSGnwjI3Z392GwrrP4puFzVa1F
6IcgNpSyK+RyfuPuQTeH1gZ/+82Txzp/KVmuYQlfro3uKQ5oQ97XiPQr3BQ0Pgc6
nrB1BvVE653X0/KsneK1/Lguw7tgX7QXwTqzatecxIH9pgl2MrhGM7FRUO0C1v/V
2hy/tDfquq33cFdAWA2TFsMyTiyAu4Mmmv5dZXPTFGQ8/jzOApJZ+x4Nzoms7u8C
syfSsJZMcl3N8d7E0apOsSNj1mv8DiDspvh/2agS7ZEm0wDsFYgOiz6djbprk6ge
cQtCDZh63/QQjcCHsOG8ILatUOTOcdXgGEdX0//mcSiFokWeXONTxvws+1v7l4Tl
rngwB3di6UcFDoBsPq5QdoJAQma6PR12BWYwPjKWyMYtPVHKDCdQjT3jo1WTIHro
09nfb3uCZVu1zhcaVa0946JWWzfqtpLTdioc9gzlhcKdyH1f+IHn0geQILmbph13
LKzDfpz2G+zlkTzdGNAFsTxk+briAi03V2VrOExbhi8ciuOZIzyElwM6u0Rmmqkh
17xvptOQ9pE0bqwyy8gfzcQXfB9kIpjQ2H72zQjgD6LHJaQJVMu1oFv0VNY83j5S
bXk4Vpm9agqw99WM+0SiveMOBv1k/jayTrRtyQ6E0lNy3fUitwFFSKd1ycLJ7PP7
mXuCTeJXSbSv+X2f77XAet1n12z33n/L+KTGeNCPR5+BYMK2W9ilz7UN17MVKeYU
sHZyAYBTGBOecu6lkVAUopAsdxK5KPSpjKqmoh6+5uFrEHfuY61p/AoQ1IMAoDfw
/29OF/ByXnwoiHtZyp04zsNkmZ83pOL8pQp5hB8oyYMVqvA+nagRGJN+kjyFvrce
/Tmlddu0xVM7NcjN+naEjsIjh5rDjdjAo+S818U1+DU0OYFzhfUUFMrJvykTAZ8X
zKfG0Mspt01c9yLCernVn9N+WAwIRxBjVKv6LKOHe4CSp2aKbRiTZBmHGcEvveDQ
8qAn2STh+44htsVZPf/Su8SV2wyewCr+U5gPbll7Qbo58UyiY9CyW9SjmRNMaKIB
9Fz7F87y64AkVKr61g8NjANtF8+Dh0ZaU79x89xPZ9yLbBI33NN7wBviwUSplUm6
vV7jNp+rSAw7lRuzT7Lx3uOJAwPqOox5snaujlgPGIXx0nJlL3rLdfUkWT1bHFTq
b+K/zME+23wlDrBqWOTUPglxPN/zrQ5RyF+ITAVzqSAv8k7nzSsxt+zhNFy9xZU4
nKjis9HnSGZeT0AiEmqPYVCGNHeIwQ0O8339+sdZKdSeURFUmzptdWtdc00+c7fS
1+zTq2D49L2oS64ZfVYLbikkcJYOYG8yzqr+cWL6+GJsMjKmgOJznRF34KjbLrfo
hSFt0StGsCgCOS9p/yYX9UGnFQWi/1FSq1ETDdlWd6geDkMyDhmW+2nOtg7Rw6gl
WXJ35umkb/dAM31QpL/2r8pXzvC5+6x3LGS6//gCB3huzYppzAsP99mf0/PgnUHe
plXgFTwr9IT2Pnm+EAXbhJtj06vmm5DEfyQ4DXCDcGaP7dpyriAYUmtEVP40AuIz
mnZzH6zI293QpuNncf6X9XfrtLwB5byUg+LiQUEQG7BxsHRVNgMKQBV5AwSFHoNT
h7p02KrMHuFj/IPAjkDyvN9wIXKnZDZ7eUfIHSl5ZFe8bgWCDrBCYZfd5YZkxGx4
Q04avnW18ECUrgrq6CjYW3w4btJrc42dyZ8WCPb5i6FKhg9zXqXLBqYukOMposIu
RdM876T1kyNvBSHM7alMx++jLyDd90a4OgFpyXRJv1JtZXbxPDOGY2sy7bC0nGTH
I4yaiOqj/gn8dibm/nQkwQZa5JtXSkQf2ZD/bXJxP3iElAkuooPrF0T5v/zq0qet
V1AxkYq1hPotlcwcqqDeKN8UjgBL5jH5u4+/TVeM66w8vUuLE61GDmY/9dMi6T3C
3A6mgNbyIrMmY3MELe/99n8jakA6Cr4rYhSDHPVrendudKaJeBV62OXaR+ciOJFS
pIkUck9Ge9ldJHaAXC6LdRl+N8wxDZgNfGcjkVzoEZuWiF71SFOEdoOmrexlfbie
XyE5lBB6ca/heJmiLR12x4YeHLCZfDlhrz313DAMX7bgRyL1yQvAeih4b/cgbRSB
kRomFE2PPGJ6ddgfaE48a3GZHEH5Q+wRA7c4gd3cs9vbJ7lnYUJ1ZjCaPTjdEMOm
VWvd83fmYDX5Wby1SiM7awjdD9fB1K9BuNKRd9/cAhEk/8XJYcbTbDkpbLZuJC+G
0Q8PQRWen2XCQN+WXuL9sLCjSrw1Gnc7dgzKmJUrKgGqhmANGBrhkleR2f4XaS/3
Ee+nyU/iKCDB6XcjVAXNDBWnt47Pj6Vor34kGRZomYRT57WtftTqEKJKviDmEkai
EDjWU8IDgBafDbSrMt2mRPyWBEaLcgGC++s0JEwm+PyNMtUcsYLUL1mHoJDZWPfZ
acEBbt7tgwl4HszC66MRNbi84Mo1KZSvFfRbvIb5tCv4a/NTBIIuTt4LyLmG1//7
tArTzxncrmGW+vsyoP4lPow3baTu3f/eW3mLIQvWvEFcY/w+La/S0Fw1HOvtw4Xg
cCobX6gjRyEV/HH8yhdfmYMFZKeu7NghYw+BqpsSD+yc+6NvP+wnzaKGXj7dtazE
s/5girRy/deUc+4vzisP/tGGi4TkVjpgPpcK/ZtQVdqyBYNlCEKElRiqpkz8S8Mn
XSc4r0wK2Ty9hEX3opcA0suQrFZ6LaVuVArtfWBAF/OWvEpuPttKGOmxJ7AGW6de
9iZJWknil+aN9RSCJcMN+mGQAT8FeDsfDzqjiOWwaHJ9KyZMV4NrjMfjLxqKMeYm
rfA0+9TM9jHMCMXroylmMAoMz5Ui2Fw6psTdcsLj/Ovbsqiyezf2NLuvdA7+Hhvr
JqMsMg6hlJMwoOO339ZnnGyBHS1hZUuFhzhobpDcIbua0uXzwM05qZh9izMvNedk
Rr5JF0apMTx1gVKot/n08yzTTaMmeExwl7ybudzGEd4kNAMJM7/ikAT+BzDxDBkG
l9j2RpBG7+hmZoWm2HhlhYQ4EVLjgYvis9tWw6kaa3ght76JZcWzL4aLDR9vBkuF
6iamrYi7WyVKYELSIvSmW5mUhLAbx+yEGv5eVPT3In+GC3xnmgp2yGHw49lKVbyU
yYcRIuTMcppnp3SbOM5MNffEy1pA7bWknUbATjjlzqu9N9ZHSp/ssqyFKBXkxXlc
iJAjBe0+N9XE0gEo1tm5e2ioTedqiUaZDi40MH7qRxrJDSicHUQPSc6qISlf4NBl
R+mpDUGB31UX1aD70wdLt+xEgWZLS83ecxq51lDf1eii//gdgsknlYdEZlBFfNWN
p8E1YOebVFbGAzw3N1bXwmSvrPEP2o5Nf26gt6NgoqDge/pV8rKEO1zDVT049RVa
PP3oJD07OZNJxpRsiQPu+2TBQkVGMrt0J2msFf8OuMdjZZxUH7aE3h6vduC4zELs
myWGcziN3nimc6ccSKekSrivrgcYaA5IRzxrrCVd2eEHbQdK9x0zYabxGB3vdK6E
dvQb/WI2b5ngf/LFR+jRFtN0xzigXi5TrUM210r+1v0CRMRo5bNgTSE9PxeO04OI
tYspYfmAp6zdHWYaya+VTgKlQgGPfE2DV6mLqIKIMhiem8GA1zHWeg6I+9j8iK6Y
gskWvqyB4/Qs7xalmpsIMwx/u5ZaHsNfsM6THKvGunBb1uwCWelp7vcrsT2jMsdi
kJZXlkTXoLFONG1MF5S8e9K0f8Q6m1GvI5jfrk/v7zSzQOz5Ej5hp6qHb3gE5hDB
bOrfLBwZ/KlC2yKc9YGK1GUzBFjFEN1+EewyjPUDA5PBeLgwB1G+NoRVfLaXErjj
HuWiFb0q+DhKAI5bNYrIl75skoKGJuYbsV73N4aaTaA11AqT2ruHdL5qWaajBKE0
d/tw+0/vLqHetaIUniiZ4HNvO+StbplTkozjE1VhOuE0/B7e21WMN5Wr47klqqCa
2A2mSwyjqcvpdyHT11ff2Jd0Dsz3ca0UDOE80bfaVxdG95S7qA188cxHMcBLtDUF
YkP8FcKxMa72x8bXgSNNftfwlNjQgJ/s+BL9ywNKtx0dcw6vWFvLet1Az0lO+w7X
GZbsJiytVg97+FDukiUwrwJvUjiwj2sYu7aATIIlCPoRcM5EAZ3hkZtruwxqloBr
3+pCWRTXLsmCIBsW0U1OYPHj/RIGlYcKhCF6URoK8B7MqwYy3k0MuaT9pjkZ7w2h
ZeSATKKT/CQko2tgQ3daUukhqcPIgVp+G3ZDSs9/V7prVZ+hd6lkKEwiNy1nNWpD
kOgANhDSYI3yFE1EFlannG7/eFjMzOS+0xSdYzQXFxn8kDQSAfxwouv50Uc6Xv7R
a+/35hylbprZWJ1+zkUuD53bZIpNIS1oP4ibot7MIa5WS3zzBkqkSBN4hKDcglIL
nZzGLLvebYV3ms4BL5oWYK1mEhy3xxn/GlQdCTwbngDiLYWAPwOUqryw/PB7AXD0
XIRXR3CixZBOkRqAiy7MdtE6wMX73/EbTASuVmQKPUnNm3K2b3RynGwjTh57ZEiL
U58WpO2C/vdgCnJwtfCpjKpZXYtfrh48lqBzr+BI6w9LSo9uh0bi/mRbUg0mv16x
Xyhjn66tNVZ33j8Xs7bWaIzllqPAfX3eiosyztEtRc3K2dUzTlai00++JszM4c+E
O9sMze45O9JJaiVM0HBNGzXsrIUTtXzkdrIF0iIJu1wHBADgvGyqF18PYlGdNJ+u
nyqqE07Nzqkz/DpvZie3y1EYDq2Cvtssa4ixvL7teFp+sJpvsERwT7xYvyW2mNUb
AQYmffWySey+u1H/KHR+j1bUJmt+mFUmdeAJmSvIFgncN0T4dUloRHOqAZjXQKtW
3bvhhh881IywHfC02YPb9IzX+Yw7s4779MqN78Jcb2JXfSLZKZffmFvwlKiI3Tj+
HN3Fl6lEf4X9DZ+k0xOQLnGhsLbgxN1hT+ZG5YU5kFhPS/sNSfQ5nc8IzOGvXT8e
cOz+Y4wbXV2dqdrafNAWs0IErkSh9cyiTuEJgQCglBim4jU3IqIahKo1qSh+9bTK
7in1lY+qp0ZIJNodgSKrn6XVtQv8T5/SAwFpevRV9i6btoO00U8hN8tP1DIc2ZVN
LS2i1RX5dFQ0/fG5gwZRF35y3n2h0d8bNzPq61VgnOaXGbKLb8wAVM0NZLL1bV+O
DnCRFfQ9XqRy8u/DjuDN+J6CalS2oEXcWAQ26NrL1nQNuQ13OosolfSXF76yQb8+
LBod5d2BjBpIUUmHTmUiyqWruKehGutXY+xlulAfZSdVLe03LrQGpk1uu1NeOMqC
U+LTmPCFUYSx7k1YenSP0EJYOJtd50gvkYkE6SY64+wStXHGqGpFXHbkR+4cPlLP
sWHJjNJ5NyX89pnDRnSR0p08gpd5+0hAZDUMpGJD+nIAc252p/OaY6hArtd8ltkI
MQ0rCdZ+l0OOM9NMduiuUMlS9OtDmD2EFKL6a3pnGmq14BBVKME364a7c/6HpAWq
dFWIdAWBNy3A5UyrWRAv5FUBjQQkHIhgEKVGh7WIpSrdru344KgTCqsOdwKq4rTM
QDLFjKPj6hbpQ2Gy+xYJTvNM2nbFk4cz41pVz+8sZjCFAd021dZt+LwO9Fu1rMEt
6Skfv3PbTa7nkdOKenzvP4BnZafwFCaNybZMpBknF6VO2jsfCwS4/LaJOx6OWV7x
jSXOp6RhRwbXvUWWccXfpRHiFr98xvozHxdicAkvGLK3Ya0fcM/Va0ckeZO3VlWt
R0YMOCJCxHwXlp1NXDNbfpBUviwnMmNZSu2QsYi/ReEpQU3xcQXeMpZH4ec+o8Ln
Ien1aXTisGuyKObwbgpDMHzpHSbcn9/0BG5dP8Gf+ucYcA/DPLNN+mUiBu4A29Fe
42y/S/+MvtfhXHk+iG5SnaNg1fmu6AgKBT+aXqKE0hsDoy/SeGDRzlR2ePWD1CQX
pDEptxstiv6amu5KSZ7VuqzyTgNecSBBjcugMkxrki7vgHi0+dppfiPwacvh38GA
erzZ/wXEMj0NKQD1KQgMDkjhzysNdVXG6+TR78gRj5Kt4whWoWiAZJ5H4B4wX4ZQ
/Ke2R9a4ptkMQnVeAILxbCbhtnd/DPbi9GsFPa09CL8WEHtc9ksB6xMIiwTULGFF
R3YsweCRAVf+iyG0w7iY5+XngqAS4Ye1bPUOWiOWQn5s/6dTjQH8HVC02JXOGrbF
TiW2BBazgU3QZpskSoa2/4AU7Z8GFR4uHpLV2JM2wK43gt03CbdJq3zMawFEDVbk
j944DihZcxvAFpD8Zr2SS8CWe9W1Ew1SXvaQPAZrUrthAHfB+buxxYhUGTiRiP4+
sgkcFZOs0PpbgvM9s5LxNH9w3DDqAhQOTKrbV7Rr/fzwVeDkF+6+XQgFvY/6V38m
0PFyy2AI8zcYnXca0qkHEkwoheRIjR+7yRtH4p/7/JBMMrh6uV35DJ6pzswf3GiO
gfQ2tq9aXh8B2KE43kL3H85DZ/h0X0Scnv/jF/bS9QkgED79u8fcDjGGr5tRsuFq
Cr1cKmNKyKtdcqw0rMFvMafughjwFu0K3dadEt2+3p69vNqiuMh8vY2rCJ4I9gL7
6Zp7BgnC179YcqhpjskZTg7+vvQOAIucfhK582zc1SlWtb+NPhTyTEcCzH8evk44
uN+vuivP0WCZG3Af1d2/wy91tI68ECTgsM3hfmbA2hER6g7XKvkAwe3BmJcQFGaU
UQY+pe8CEsJ1nPd/wWsA+BKDz4hmEamt9C8CivZHlC4GR0+qbPX8gL+IQW7EhYAs
QUQK5GWhrh5mRMmXEwhaSuI/hZNfZccssr4lhpIvil7EdnfvHiongE0oTmA16Aex
kehPwFx1gNdKbUk0Ne7MLrUuWCUTvMTM+bb1pCvTiFXljsH2USDJ4xcDbZydCiSX
Ig1xlxS5RdhCR0TU12zGWFHDAIIi3KtH1VmanVBLMSM2RXKHiACbt2WI2xqip8I2
N3UsanpmlaqbplGqKu+u0T7xDLIK39rN1Or/ElTefSVOrGQydkexP84nKzM7dJRl
1e8x+2+r2vbzKXwc5rmD0YIJXIB/Cm2wP4A7Hc8diatBrvYdv4Gjt7QJMdwz3iDQ
/SQQNGieI9RXsl0fMhVIpmj9EHrO7ljxANlXSk2mnZs74Llr6EMxf2fcJ+7o5Xsb
akDhkT7hQZdkFdrDGdMNCV2P9s6agunsrejjb8MuiCcKajaEXz+3YUsOsw+gHz1Q
oZCZIXL44VpQ7J7+1C1Zngag5Qm3Vyx6KDIoAkGS+CkVkQVeojA+3srj664fzwD/
jrR4dG34eCaXBouMUeBKQPjPwPpvQpYgaB8TfzsM0LjM/2zdlivrKKjaV8cWBmHI
zo87bzl+WUg4roas+yydoBH+AKBXDaAsHCLODDtqwO/6tIFNj3m+Ng1GnLsStPzm
CgEJAGpFJD1rDNAj9RRenzYcp5C5kLWLsXg4VlpFcOJdZGuRSAWDc/8GDcv/y2+I
q/ubdQWMeBvI5/QySq3wBqRS0J7XGqc+/we1XEmYd1ztj6ESNosAOtt2czN0OYzl
D8/bJDMmKrx+TQpLpV/Cy9fu2RkhSYhEpw7JPkYUszToLMPcP9u6vSSTS9Fylx5R
lLVJNJLF1BcMwrcNKTbH3tr7Xm017cGq/uhyInFJn37pXDOFbDKymND3zY+Pjmnv
SCUInppnmhEO+X/jnAVXa76qEQ9kiAruWgHHs8xjY6AtUATeTfHU38sS0ab/XJCb
9hqirpoMesCeewX4eRDOMB5VLjYfGP3XpgLk6fDcQGe9ELzgiFPDXMT6mX3AdAll
/rfSxNK4ItRtXOlMXTXDAqDAY7/QUFo/Zdf9BYwsJoI4LEHPp8/UGIlN0Ro6laSS
65UDBL22u+SEWyjGvugN8mZV2N9PxfnDwQHbN0WWVoFhY3URkGuOvQcIXM7D/P2k
EbMwVLHWiAIN/Tdl1p7p1rMn4cY/SRfWLkRKWy5q7UPKV0hv30POWsSbhJRTuJfF
aAguar/XGhRzr6Nr1eZAYWsyT1GVeU+R1XEsGzwlclcPGwBPIdDdppNI/Zpxzn+n
FmPlCY3YPzW3SR+OIO4jbwHUuJ14sye99mRKPd7qAisQtkhsOfEDSnD+9gljXUbI
BztMTkU7L3gJLrw4gafqKmGYVrL8fBV3buwIKaYZiE9sceLpYPmFQbZ6hYp6Dtnr
TzhmRgS99v3HdDPU5aG4CWoL2WNUD0Gxq6HKrDIyqITA3cos/cNVPry7SbjGklPK
nq2/Z/qMz9Rh0DmGif0JTfBWKz6Paog9STX59DRvWZi4rOpT6+yvQu5esnhvURL/
THwo1JXSB6rY77Jhle89Ub6ENSFc4bpk+RSXlZee2gPqgaS+FkGKsb6Wx1JkVDsT
PhQZ62J/eyY8wPrN5/5Wzllrb8KLxFG/91m+VQpbz5CAGUut0FrHVsMsS5aLDtkZ
yF6VqjSCzYz2q7u2RpL46OZElfSOIPB4aiBDNZ92d/c/pGJuxHXbsZQYJW34mhJL
Dd77ap5tN0omEn7B7SAwKtoQkHEUocM+3pL82mIzqNH5p7JCergdo29nziSvSCf2
L/UHx3AAfzMJCisJ9PBIAzu1jAU6kpx5C+x7JFqgCLvMlaupHzuofKvbZCOKvh87
4pXwXYOXKwJPYQAu5aOVzEGgCLp8F2qE9XNjtbEGVH+hEmB+of1EMiPXZ8Vs3lEI
223U6jXSxehNv/O3IGNPfOEaZWpfjZhmNfeNiSZhda55jeBTrN5g4lQ5Jev0jU3T
k4z6A61XWBtIRxzMPW5TttBYHsGY4V++vUhPuY30m8G/DCk9RawjhO1uoy178psK
m9SwjW7gg5uRUlhC80TTaV94ZMNgRLftDlbiEuCoo5l22tryYXRnIR5JpgyY2Cn/
MrapGdHZHL8TlmG47BcdUpn7GIvCM1ZyRxR3R9YRtOGf6gyb3MHDsH90tBkqIcId
4oZs9wjJ/aFnBXI3OW9ES9BMF+AC2PE4ODypOeSZsiiAktET/02vUT0GVckITMDE
phESfhdUvnzEAIMJ/eiv7nbLWdvRh0Uv+iJgzDfRIZ+YkTIZHlDIAuqvIRDV4eP/
X8aB5EoPsBHgsMntOvZiFHlrk3bwlwIwcmc1JAVb1PY76A+kHfn69Pruqyb6Afdt
mCP4n0RsBr9c6/q8uaPEeu/7vaAswzFMvrIqmapySvdjAMJq3/2P+Z+WV3gDyhpl
UuJ4PR/aK+hMII5j5UcxbDUd5DQIDbG55eWPt3/ufIwedQNfIoJtkxzC3qZrLQZa
eJtTldlPMlAPpLDRbrOUKf4I7gY9PdqrE2w3ZvslCEpJOGGBkw9R+RyxoXixacMs
cdpbGA2PpRI/aTEjDiVP0dPDT1xMTy4CTJtQjVJJXjHmATQVZkk2RzqdzIGUXxUt
T4EZMQtGqjQKSW/xZcZH6Bmnkd9Jq26a5sDF122k+xxB9Xo6mbKY2DLMf3mDgv7r
C9PDDABDCVRPJf7PJq7MYF5SLp9/GAtHGfWaYKqVqcABo6DnYlFDGfu4k1j9xUg1
Y9wLkD+hUhomee6gQPi1UWOCS3eT66AbdypHGucLlU9lw+6Mpn2q7k8Fla5HmoKF
BQD22OWJgJ0sN4ovTQDfC/h96kx6x5jfuPbWMnhiIeGlpJ5MGW4PgG0UijB/FKbL
lVZOmT74DLU44+sTlos/0mOx+DzodUDYHUq4wGlAfTsvzVeBlJdb14pSqqBf6EPD
lwKROxxpALfMvkL/aGu+BlyJ8MEWIaJkPisICqUwQ3/nd6XwS/rKbIZ04Tkw0+5V
57lMosn7B5CkR0J3E/QTAbRZJLcHeWWkPLYBecEfZGB2RQ9jvB8YM5d8Y+vzkr/M
0cEoEzZWGh7VSgXFwcXhTplfh+hkGZKZATQKOujGNNSo9YVQCiCkQV29SP9F6DGr
Y+5wYLUYlWGmu/9fXHcodl86LyLWpyo+965qaaoV7Rr2lBzi/fXkx5ruJKulxXx0
HqY1DTHoV5/PqCXEST1Rqia+m9rMW0CIH+B6RySKwlLnDaPhGwh4O8KEapUDr2cr
+IWsFFuUYUcPIt69ZdolvP5xgoB53zmR/3uIDdHul3rx7P6DtF9L9J67UgiLHzHw
VxWA8c0AluJcFFV+4z6zaM7WgG8XnQBn1O4wpg8QF6DgcK07ZrdZMd6LqX2hCx1/
wfynJiE3RpKXJg1pKOA+4rA01mlE2QI+q1kZhQiZ1/j6aPBm5OAueUA56AWftodL
K0lglCk9ks3vSC0qaT6/oI7G2R4OIvdJa4E2NVNqRyY/ZvifTwgwdBnig0gg2Np3
ASduNwxX/JuxNR8j8qx7EhBvXoGuM0OC36mnGLuOTqVPA9LCt0YeqNpGAaiUBWVe
03PPXjzjH1Ja4vNez0ZuQAqPUnFORYly9SaAVAceJuOJln3GFv0SErkdMvCqsqi4
Kn19Rj2Qv8BP2vk+TMjGkjsdrvFMHGABO+6At3dkiZtSmCQwAd3OtiZ4mWim/8Vu
tCblWbntnHO7OasWRmCcM+KZ6fC8HKnDs4YsRCvkKOZB6T2gsptudOxBOmKoAHB2
nnyDp865bT//reJIegp+G+saGa+jS0xb5c2A+F+yty5aGoyhS7DabQAWvrPA35FD
vBYBEBGMOsc8MQCAxTB285tE8SOg+JKquR/I8t/xYwPw9hqEkclv1+1FGcIEarQ8
hZyOvHy6nD00GBJiZlCJCKKGw0r49Gb9G2F6WuDEZGeuKyKBwv8YE17TjJp4OcTF
lzHB10xBmEW+XGUYRDBuNWA3mmnYC/LaVN8/sJvVwk61v48HR0+d0+ilgiRzMgJC
qK9vGfSsYlXQWdNwMlt29KZWPwTmAEsP+QaXC94EAz4gdoaHVCM4agY1zDNMcNjq
eGGXdQ/Z+NnBq649s1KPjXgLXG6cGTETbZdGiRhIHXEMTKakt953rVXquYBXcMr4
LelR5eSOww6yhmTbBl1JoH4N9m1F6cA7NB2PVat4ZYB8B3wzWLI+GYpzQu7YPgJm
32ur1NBAL46ZJQ7HkaKaXjJ+0TGhVl7SRXsgvtRaf9cjQcKWAyKksx7g6mRW68Jj
cYU2xfY35degVv7B1QoWWaGXeW7KpEvCL3aTkTBzChC5bYIEpPIAAI1+eYB6lHSZ
seLeIufWwiG5LZcMrTwTW1vQgI1Dil2XaWzYMaRupNcVow/U7PSqT/jvv8uyayiV
POtY+H6USfbvSlSD23CyxgDGB+7EPUbArwS7TqK37NdH7VFn1KFDGYW1Bt80N/Qj
zHHqklDewj2d8XcnKp0oAgUB7V2PyL10oszcUWArJmdG+dy1yEvEZ9b8je1c1Xnw
CZZ8B6I8P1UUK/DQItaCo8MB6e1bQ5xetcJ70IsE+UFUpKhOBXNkE0wAL0GSpdFq
SLqqOHhWNb6DYK9XlWYiusAiswdRVoEvddxERRxJld9q7Bzdi5VRX5ypJEndup0n
RQp+VcPYfRZr6u+84QwBu4A7Yk5aLkHEgRvBEDhgmkYAZ3firEFihkfifqCwAss5
829G8H15UBJkIbRZZMXibOQV97am99NAqxeWYFEOqBPM9WAugyYclmejJzpDJ5RM
5qXngSFzYKf3HzND5KHnnvtRCSGVyfoVcU5rwRkGtaJ8NwYA8wcOq5hPznNANaIW
6ImZaQAJwBHOvOUH+4Y9qzudpvYlitVuHeg1Vn/0a6fUnA2aefsrUvnnynvRtsmq
/v8zAS0+dx3BDMPtXUD4Z7b3RmBU9ArJjukL+11pU94JCXW7Awmvq7CDVHjSUIhZ
Rr2G/g222pWBDsfFQp3Ru+Zh6cJ/2+y+2aj/PrxxOeD5rETiYlG9sCCEL8ITAHth
ze6THs2022Qypf/Va0bXX/nzIvZ1bt+7LJN+CzmNpfcEF/uDfxzEhOwq4CiJQwNW
XZzHK4loQTzV9oWavzyaHeDt+537wyPT+zMLdCcvpqIzyi6w8RB6epvuKvTdSsqA
xNTOgVcNW++Akb97lQrTlLpRaYm7y+UzX6HiQRaF1RZhkre9JT9G3EmdWr5VtCwC
8JKFX7hJkJya/jlbZpCIZmUg5wLZqOCrtCnF+AJv6845n2O3q1VlXEGhXyQ5YaMY
tqGmepX9jkyPhbcGNcDq4Mei++VJuCWq+YSw/Gqjih7vMSCOf5v4O52BOFosxr7w
r0tttWoIcXB1JBOG8CX4oWatZq7kfww2KL4zf+Q9vs1lcWLdUO20Rn8ZrFPBJ8ld
PLL8MPBi9wMb1FuWTgx0TuYxYzvzKbCdNv07IawBj5acONs1h433/uxdnchx2PRO
RH5281CisozR4tmgpj4phvx3qB90AlPR7qgAoSi7lSy1uxLiJWOU+gQxG6a3IVDn
aLz0CZEcJrUf3zX5XPU1xp5lrjLcBOktjpN28LR05TTtKjoYFuQ9Zopx5iz3lIs4
28ei2dF+WB5wXyX+dPiKfmOx3hYhVzj3K4yFHXhn4iAiyOrN4Rdq+87qOV4nq45F
Ah0jUt8jfdidhRhtWpIOmAWxgxZ9Ksq6qgqqsEkUfZXH3rmCBSW0Cw2aOtc3BHBf
/+wrNVaNJETilo8SpIpxmiq/fPuyWhMtGGNhpl1siCHe4RaLIbt3w+T0k+9z4ueb
8Wfbeeujg6YKicyNO993JDv1jCbterwVW/Rj6vrEmSkWwej2v6wDhbFzFcF9pwz3
dKeo9K+fhbDtYsIQlZT40tx4+gnuq4xW5ZpmoPpjWzF4/Ggz/JnANB5RNMSWsuJ7
MRgtz7AZWKmJmc7oMpArpXSt+6HwACZF3eNErH8pzh/tNsKR7G+XjVPG7YdSCvFe
isVS0OzaN8Ennve4Ry/Yjf4zeAVwO6frNTp5KJtH/smFF5gtlk+v+Pzc45GQ8g8X
QHv/32LWlWwr8QhRgojJXzmSsOLVQGnWpJXv4fAeslzFzYMbS/LL3BC04byBQ2s4
lI6JvSztZ+bH4O7RORgI0uRIgzBy/v4m/kt4W4BqRxlev11PxU0ja863P2EmpUIN
EB0eILkQCOwHZtQ37G79FlZ9FlaU7Q4TicwiWm3l072qhTucTqSRonZjc4R5n+1+
2y9ijNmN7tIvgdNTEg2ncplYoXkyMHC5ecOqk2dQs0NvRdLHljd3aFWh7qppkkJP
ICH66Rx8Bl0QBHHR72n+3Z1o42NCBxdDQryRQen2BIKo1mDIi8DyHX3nYZClTu+E
Fv1UA5A4KzJTC35a+tv/sAGKQxWdA1lhW9+eLksj7yu7SmUC5d3u5yH8MiEXnVoa
+GeUA7XPlxmMHbCGRc4XWfnaJaCF8G5aPkxp1kOMcDapwNRSKqroL+4pI+9CFYqQ
LA1kohdrqGoGkD1nny7r7hcHzUjeZTon5dWBGpMX8B/iwPBReb2JulVNnkyrL9fe
uX4bCc98bAxa3ZdWw7IA+lhUQOQMZhls/Y4ezbijB+sZWiXmF/i+56i71dhUzpi4
wR5dI6dg32t2l7S6QrW1XjA80Jo0R0bkbZYtGWfhH+HmwzfW5O+ivdQA7SEZnqgP
Zu+PFYJKfo2npFmY7XhDJVBRLYalU2BGaPEU9C7hkEE6V2DwzYjowOzboqYZJ2Gb
j2u1Yf6Xefk86uhLQ68qCfFvXi2ddUF/Efqi8V95Uv7dqzexQ3JtCJvG/FwjfqEy
FzWhdW9acWq5I8YjZarNjPIRoMQBq1RQ//Cxo75+C5Mg0UvBykNdzL6T31vMnd/+
NB7m6FdRMhjCGBtDCOGZr4vPe+Iocqnk3L0yjwIO5x/Avq1oj46lRO0LMkYLE/vd
O5/0SB4Fb5/2SrLkvWBILI8GyQf8Asu/IWW6GEsujsHmSiRq4NzyEcScWRbNfQ7c
zSRshT5ijfgbRgOUK6Q4WKeWVIK1SYndxLGu4FotUsgR7WQH6FAWNsb/PH8pBvHU
jBUyS8/xhRF6Ys/Wv7gidBEiK6Sbm3Tg2rgN9UoU9qBkh/XpkiXe1VySGkKkH5wZ
+VnrS2UgACElMYF0fJB8+PsYr+0CcQK8cV+IqxFv4VxRuGy33hR6KBaxkz4+9yDC
5SFlI8dOkQ3PFcc4xQM5nWKlii/jAOnrLXnfSF0wh3DAcTSpJh/1F6h/y/zeyDbw
kJAO6moCxP5G5xUBClnSRCjSkXuz2Wq4gwqCMevEvYYnYOfoGmM+cnvfq0ZyQuxe
oxevOjPcW1rbil3cZqTiw+gqOz6eaOInaYvZacTT3+G66rvTbtjMQO39L/Imaf/b
rGvaxLHCOoxwY5wMqbfuJUUV4E576d65+8w1bydEi6EUFA/h0BsAqBblfH24naF1
Aj5LjznJvlyZ0BlnnmGcfwvba3ki1oXdFnYtn1BqU0o6rTV64C4NxCAGZvPmUFb+
gqazSCZlXuoiDC1cq9FFTG9AmbePHwCKdSkZEDQ2x+e/8j+uYh8Wq5uYlGuYh6Eh
p7CMLF527EPomPhvnxxEXAMnZPylZwNj86JAKpAPB52r5VcrL8BbnH0bC0j2eSk7
hwZtozi0y/hCRorG2DxUOPEMCxDfb/PnMHzZafUMQMOA3RPvJYayewV8bt+E/qDj
9cyQlY4eNyaW5r4P4IC7DoLLJEdQymE5KsPi1246XEaVMmqVZadKqT1UVxS74Guh
MgEaw5Z2rWr0v4V5MOvbkYm01BFq2Es9oDJPXcXXwfnxWqPrpbFHpVVL9VglR4fz
xXvdl0JUEFSTqfnwj/jXLwJHa317cTe2BLR2Zz5DDKe92SRDKdOQ8365C6ASdSZY
yiuBlfxLPSdl5pU6Q4zPaerr163GyQVi/O/Hfi5X8SQUj5zPtWY9OK/erW0fHKOI
yr7DMzPun5WD+yZhADhbc1R1c++UVls6nriy0ogJbvqt746zHjvGMURkgIVEdYCE
j+7Qo6ZZLvdN98xuiVYAbKBxDBPFOhwXtGYAwVhkvGPQlSnCwirX8e+8XUmME/0p
MQ0CeSg4BfoJ5WaGPlXtNKzkr7TD1amRlmUH05x1T5M00qcrcGjrswPZ6i6KUOTO
29x70Y6Bu4GlvUoMTi3OLY7R8ORdAFB2s4D0X9uCVuxTUZekphHuQvJRvaCpck4n
KEcf8NCNrrh609WbvxzqlF0QLTVw4Lcx73N/fA4vufpUJc56zbAKaovgTvzGMb0F
n7zdB+6hYTFapCg7w15MUWxsabqfnQts6r2NmIyoE8XEgOkJ13RyH98f8odkLwRz
pA2Wp/dawUSsu4cCgGqUMl2W4UWCCqa0G3Qe2Huiscn3C8C1dsle1ouI3YVClBvO
OqVia4x2Yx/Hpu7238j4qCHO4yo/cF16RUbvq1XYN5MI0LOyAH9/9vVeBXrav3bK
jVN/Wk7vVdQ1npSiyZ/8C+Rfc0OONcyrpOMPctcAu3wHCIoKm1P9RrHd3urJv78Y
`pragma protect end_protected
