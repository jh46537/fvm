��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����p�0�F���)�ã~d�:����f=�n����l�@>O�Њ�۸"�#~����f����S��UT���������בJ���\/��2����r�X����`Ir�K_�x6YV����(�/�~�k�q}����;)���3~�=�FgBBKO.��}�@��z���̥x�6;���X<�����~2�M�2��$)�sFaa��4����9Q@���e:TWrt���z6c)�<�~q\M6�'����/ q	-��# � � ?!3�m���{�D@� �+P>�e�<>��]zF0�P}��N�в\� �Jy�Ǚ�j�qAw�IX�Q�2�6�o7�O�7w<S��H���y7
W��w�Ӯ�T��Qg�"D��^�U�L��u~I=�5U�$��n5p�V����B�E"i��z�MPBo�,{�օ9����Ka��s\�^�d�h�z$U�/�C��Z��B��Qs]I>^���-J�Q�4֢=��~Oq~
V���qIͨiu�$֤2�|���g�J=���w��Ob�o-�a�����,?���ғ�۔�Ov��`=�w\�j�T�x3����rz��GM�,�����Kђ�^�ɎZ�r��R5y]��37�/m���ǫ��/6'Wl7a,
��1HL�C����%�����m*���S�B��%3���7��8[Фd�H�f���6��0 � ��޼QY6�vm=m�붪���+�~�P�\��ơ81�v�b�!@ �x_d����|��n4e�V��pAw5E9)mDr:�4�\�q��7�;��>���4d���iW�b�][��=�!ӎk!�+��b�݈Nܢ7y�T�}�X2�r�u��B�;�5Ta���N���A�:l����U݀Q٤�ld¾�/��*�a �P��2
X�+ �=�,�;��Ǘ��(�5�I�� �Y�΀~|��U`%>�����ZT�]��g�0^��nw���q���jӜ�r=����K!}��u3*�>G^J�X�l�����ZB#HP1t*�#Ҝ�����g=�����Q�G�\E�l-�A��c1�l�b�:n�9Cc�{y�>�	ݞ��/��2R�C;�����^�;�Vl���T�M�iJ�
7�&̩8�I�dCH��,Q��L\]���ףb�c��]�Y�sx���_�6�"K/DM��4p�Q��YD�D=�G�P�u�~p�N@�u�O�2�6�Wt�q�i�[���t�X	�� �F<����8�\q���~����{^������z�,��)�|�4�V��{�M���� j��!<LBsZ���AJ`A(륐'�8'0�Ǣ�P��{�����B�3�s�r|)r�QÝ�,{Hԓ:LH����rKw-:2St��Ie�P[�_����^�8f=w��jc�Q ���"��T�i�n�Vӿ�m��Y��}f������m�j٠R�	6ZL�l��s�Y�*+\�m٭���&>-V�ǈB���[���<��k$ǔ*�3g/b�5�m&���}% �����rW}`����)禉��#�xE��}�LD����S�&ud\[r�4��,�7���"�ept+]&�	�*�Ur]�lg��6`:�,�%N.nޝO�c�}��hhXM)k��꣸�M:�v3S��vW��`� ����1�r,����9XH?���ƺ�ج^������wP۩^G�&8ljɦ|���|P���V�.���D.4��c���O f�q�&Q�4s]&���@�� ���7�O����He0�����C��l]�HlѳA}�Rto����.Yaq]�MY�����%���x�S�%��&�&�o\fQH��\3E,n�LM��|?8�kf���!s��\1�A��4�D�m+�B��)�MB5��3hmovX����Nk����r���HGA�Z��D�g�Y3��Ͻ�w* �?ՅV��5�J=��ƌ����>�V����#7��;��Q��5�p�"}�s9[�B9Y<�S�ӥ=[k#���y�	*)��z��Qb5�:�-"B�]��'��ki��B!I��?�#�yhtIW�H�w���c"q%�¤��� 
�JU��$!�/�/���ɧ1���^��#P�s��)"���6]�W��_�p�i��F{)I�I&�zVi�(u�(4ԓ�WGA����C|*p�o)#�(o�nn� q�&�
�U�zP4*���&d*_��j���eTc����p�:��ݧ^��&�I�e�q�-S6I��׻0C���������i�K\���?��{�!��mC$�}u]u!ig�E��xZ���C�Js��"~�`���ic���軰BM!cv+"��U��r���AΧuF?���J1"��m�\�z�K��=U<��Ɉ\p�a�>Cܹ�vS���;�1<�!`�.�ɀ��7�K�б5��N��5�p; L����K?�_Z�[>�M),���B�����G����JV90��?%�	���I7�g�}.�ʌ���.Ӕ���BS$Q�K�2խn���S/����2"��I��4&C��8��w�B��dϽ����&�C��{�?h�-,>0���h<��Q�ր�:�^���%���.�����>;�/R��r�N[D�9��+����V�6B�K�kNk�^>�Q��?������)��he��\���Fb�r��'�߯��>��G�'�����y�d��8�=��ZO��Lv�|�afW	��Î���N�M��nC�	�Ox'��<�X�x���*g@�X��y��(�����A��$ܿ��o���|�����Ş�����l}�yi����x]�r���T�'?��(f���[����ū��֨ɮ@3R��ݣ_�Z�fS���g�w�e�f�6��.Tt�(���Y�ݼ{@9�a8wUZ� ��q^��\n �u��d�@CU��"ʮE���%�s>��x���	�:'&�պW�k:�m�>�=�n�۰:��W�]X������6A�sTu?��Wk�W9Z�V/
U?�&��� �J��Y���o��?��N�Ƥ}�1h���b�E��Ė��C^[z��g��&��9�R��p�����2l���Ҭ>�^=���Z�����S�wg!��R��nԐp��yM ��[FU?�54�!�e�=�QƓ*g�L�kFT��z�y�k�0�q�̲a���Q��N�����a�E�������`�Ѓ�2�V�{۵f@u)J@�*��bO���W�y�TH�C�U= �0�|`3X���ͦM�S�����C=�g�$OR�2�U�ϧ���y�}g��RD9.��z�]�1˗�S\��N�0�����
^�9�#�g,Td*�ƤW����2s�hZx�RS�FF���l*�=����ZJԕ�4�����#�Y���^�?r�º��ڒ�N/�N�����9�i֥�+3���������D���<��� \&�����_>��TR��~b���_nz�[�R�9��	D�:����z�Vge�Є���|���90�Z��)q�彩�ҋ� �³��R���k�v���<��%���22�"�@��$�'����z�s��;��3@�+���_�>׏�F�K��{O_��\�#�E��:a1�/�8B�E/i1.��@�Pg{��	�0{ SbTp#A��=�7�0�X6�Gw8[�Sg�m�k���L|)�:�߯�W��$D�Eϵ���d�\��YS/)a���v�r�~´�=�q�G�۰�Pr�W��^�����r+p�"�M��_����K�.by�7�Rz4��?�{_�0��^ >�:��|H�ǈ�V^"�#hC��s�4W�#�z+Hp����܇o]>���dYrG�O�,4�q��o�������7�Y�&4�#����ܖ?p��*]47 IS�^��(�+U�c@�~�춁qv|QO|�\������^\���Z�h�A�0t���=��mK!��S��##�'Ϲkl�s�C��VѥpP��dg����)�����PKnO�����1L�<iI�ϛTy�DG�C����P���t�06���Д�{��e���8H�W�~�w��j ��=�IDm��P�j��C5=�Q��20_�^W�@�A�,:C�6����v�:獉l�����n�Sh�^A�g�������)m�t�m�����9Em�e~G� �ؤ��z��*EW�<��O�Ͼ�E�gT���8�B~�@��S�86.I^ݥXyyA#�vz{@ρ��V�-Q�b者�}?|����u�(?�$"t�����O�wV.���df\�|y���*i��"�C	��|qW�'SJŽ��i}i$k�g��gd��9��>����;�����n�0���0
�UJ�(dF��R���Z�I�\��\+�X���
yhq3�@|L�|�W�C�Y>8=d��!�h@ݶ�զnj$�u�f8�?T������ܵ�N�' � 5�J��d��aL7$(����jH.d�-N�F�)��%$r��˯�⍜3�~�bݴ��hL��ǀ��;�_x�q�ۖ���i��[�Q�;TQ�f)?8��a��8NF���,�E��pU�h�f�yU`��X��T�!���=W&��VI">�u�Ny5G�-��[�?+�1�ppҋ����}� ;y�F�C��ξM��X��9z��w�Ѹ�Z6AF��4}�B{�K��=K7���xժ�>�o�o���4��i��tT��+��gh� �_�*�^J���5�(8�krԓ���$1�xf�HĄ�+�;�=%�U���8��2��s�_,�"���՜�p�ךn�U�ۦ�c�}��2vT����p�MT�#zJ劀
;��0Y���$����i�iO�,.,�p�%B~��u?T�;R�h*��ç�8�����h��z����@�x�|��3�c��<�U[Tb�'@��NƷ�/)��d�:�Nw�3ov��>w�F��$� �QD���>l�/!�є%h��_@&�T4�����8��iu��`���2��S��[�u���[��������ûk��&B;�����E���Q{��v�$D[�e>W]ޯ��tQe�� �!��@V] ���,��#����S�^dsal�����ͻ0���<k繳� 9V��0����*�FI��kQ?�/������_�NB���95���/'������Ťdrw�Y�h�i���N��\�^�Ff?��ö�Xj0{�h�kN�>[����=�[��ۙٸhS8�d>v�S?܎����$�����
?���l"q��ge�A����J?X?��r?b��\���񂴅�����A|����a��dm"�/��O-;!��H%�|ܠ�.N�@�ۓ�	��e�S��٩,�>p�ד`��T'�����݂v6�;��ɠ[:�\���O}&�:�cF�%/#Tj���%����81���d�����^�}̾�xaܬq�zM$n�M.��M��*"!������&�[��/���v���ES���p��7��֝k<��a�6�M`�\	#� D��~�rG�Wf��,;�c^��3�'�XΞ�ƍ�N��GRmh�(���g�q-x�"��x-U%l�
7����%XK�G]�X�F���>jH��S[�lV�	$_�����y%��L+�&V��[�{�c{şhG��޶ު���&�x2u�E�fVP��i�!笩
�U�d�OF�Z�s6j�,_פּ��)�=3�?�����?��5}��?G�<I�ޛ���?"h#���Խ�}��2��"��T���i:�����ȸTD6sy��][ʠ�ep�����M�����"�ݎ4�
.#���y�^X+l�<8�MJx,z�k�(실<a����\�v� R�d�U�$��5��h��cN͆�r@;']��S�/I�2#�y��&���6��Y�d�Г���F�u
�`Q8���˝H�����ҌK,�?�H/��QZ���;72}���� ���֧t)��D������TX����P��n�Fe����r��z�D\�����*�5�0���W���-��tҫb�'�e&��ӂ�!�Ǖ�W�T�5��C�3`�D<��D��� [�~*.�?@&����zV%�Z��T�����4�[�^-M�x��#f�^�&�N�׉ȥ�G�+��4�h�|(�[	��4�u {x��z{`k����~��i^>�����]��M�Y�R|��;^�Dϫ���/�d]�N�/1���5{�:q �Շ]������Kl���B��c�Ig�8ld�@'p���w�n�:6�f����S������oi����<���"��l����{~q�sz����5�c��@,wb�)�6Iɧ ����j�_�M��Ѭu��|��Kaj�g�O��E�\Ʈ��Y[j�Ɖ`�hEx����t+}֘k��sr��H��gP�
�������c.��z\� ��g�؄@z^����X��d�o���3�d\<�=D�&���Rx���c��"��㭅9F!�A+Ő����Qn]?{#ħo��i!�/��/�\�sRi�b�WG���郑3��oJ��ZRCe+�/  j��M��Hk>���+���B�S�bywP=D(�-C]U����g�+�S~j���G%F�uH�E�U՗�]��$kS �o>��ی�V�'$�[�9���F���E���t�XIȯ?���=�{��F7�c<�\=��l,���� �P��W�Ā\�P����~Q�[ޝ�ixp�i`��%G-���A��&p��	�v��E�^L��An�����m��.Ϋ���p� 548aQa���`9h��	���12i9ł����A����V_"D�.���;��v�� k�	8�.���%��
y����V�Zܻ�/��f�Yf���g�/V���<�D��ZLD�w[�8ʰsKB�����?"�q� �޺�r��	�Nld�T�AnYɧR�DS�s@��^�%Q����]iW����Y _�
[vUl�)6�r}1��x$������Cp*X���TC�f�Pw��%1X^����'b4�h>��8p�aʏʷf���Y����ښW�N�x0��ij'%�z�:_��քI@���oL1x��8o8	�-L"�S>1����#m
l��T]�K�dG��-{��<Z���b.�fCƿ���C�ȴD.Tg��T�I���!�n��Ȭpk(䊵�� }n���Գ E���9��C��hL���a������(go�`4TKa Y?�*Wve3����\)�A��1h�h��g�=���Ir�^hv�@>��+��}��]��t��k�E��p�5�	7	��ie��l?��L�}�6���&qg6���n�k/5,ca�%ʰ��
�	������!$B�qWی�<%$���ߨ���N:�?csp�g��r�J㧔Q��P[��ˋ��i�o���1�؎�C{l�XQ�V��eb�����MO����ݗӚ�:�)^	,b�z�-����z)@����0�82~��ޥ��#2�����5`F��/��e���	9A;E�ݶ
�����C�f<T#���s�V@�.
����~���� ��țk@�%�jw��Q�|�� �G�x�A�S�{F�e�y�1�A�ﳆ�4ֳ~��B�����P={��q2}ʁ ���i��{��E�&�п��\��v|%��<����W�2+M'x�S�W��	c�AT+RfL���!?A���(,k���σz�a��I� w��u�����S�o���|�G�� ��vGXY�$o�s��09�|��^��Wg���	AG^A��d���C��䓦x��0}���[B: !�=��Դ�"�̒���I:xX䳬[ti�Y�DM>E�0�f3��`$sk�W:�}HmQ��n��J�2��Z����H�b`5) ӹ�"}���v��nM�[!W�����8§��S�aʩ*?��Y&�0�3�^n���*��(���7������ն�>�?��o�ը��9�����wE�IP�f���;���F_%YdB��l2g"�y��U�Q�`�(�@�B
X��T��6���M��g�
�`e�&[\c�����s�x0���E�kҠ6�`�G��YQ���U��e[]�Sp2�W
75�� ܠΓV|:�|_����Z�;���z�C����U��fdNY�\6� mM�YA�ƌ�n��1,��%f ����8������P��b�;M�-o_BT�Ě��`�"��_َɝ��q���WX�#E������m����?�<8O�]>����K��j��%�Ly�,�����y�/����r�y�$�
	�C��d|(�B��/ڌ�l�\;&��Vf�"�y,�닏թ4Rn�*Š	�ᾤKc���Pcƫ.�Z���L�W^Vs���w왈Ɣ�z�T�NO
)j�n�;MXd׼«��rN�LX�ϵCp�t: .�tj�6;()��+���&�J�t��-��?�B��W�:��
�U������R�y��f썣������Sᩇ�󔖻����W����<�_X�V߿��69�E��{_Ȉ�-Ԙt0\�L*BVb^]�i���|b���
g@��[�W	�[�ӕ�IIj!�8"��J1�A�A�QK���=+�&� ��.mye�n!��-D��FxH��	�o��X���&Z�y<����������u�s�g�%ȧ�R�x�����Y�[����XJ؀3��anO� a�H,��$XN�I>�D��}8K�cj|bc,��M�}R��Ԟ�&������~��8	&��NØ�j���ԠF�"Uk��Z�p�@]�����k�M�
g,.����Lzqcz�6��Wײ�9���M�]��8�bs�[�H@Ej��4�hو�K&���X���*R�DQ|����|�:p$ �"��	[��r/��VSK�}{���z��NL`r�����/X_P�-R���=��LI4�Yq�^�am�9�+6��t5B�[�T��:��������8����/o1t)�T5�gv�%�eC�S��PHJ��5�C�l�4�%p�=]k=�:$?)p:P��:?Ԫ�v@�����(EC��j�O#�ގ�VT��s%��͂�)`��*�5�r�MG���׾A�b\Ό��N݀`�d��4�:Ш��г
B�ۭ����b)T������B!SP�H���4Ĕ�,����Ȁ_�����qp=�ǳh�	ȹY�|��K����	�#�7���������+
��b��,H�r����UE4�rG��Kɀ��\��ᶧ�	�!7����D[P���1����¹�k���`��1.��=��lo�khA}1��x[a�-飕㒕����,����%HyKt$����\���s��0h�� �;�
*V�'�Ѷ�C7����;��{���xu�O����L��:b��j~���԰6a�J��N�а��6N#Y�\�9�]��ȆL����6LO�<��p�!�J��?P/�P7�++{b*���)P`���-q=/<