��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*�����W51R����\�Բ���I:hިHm�{#1��`,]�F����=���8M*�ҧ5 ��O;$ʢ�#ӵm����za�0R�DkYΫ��;\��ҿ���J0��^=��)T6a���za�ѯ���ׄs��b\�*��&�jT�3��t�x̬�����o�����T�#�� "�dB|��ꣀ"_�,.Rw &���C�}޲����Fg;:!-o�2�+JsB�&�v/��4�ڦiJ�.��xe���RE�/(��o�]������a=]�,l2l�CA�@��u�:�Սv��D��r6�Uy�R��m��()`m�[�B�M��X���2��4E��9gZ���I��{��U9���5�q9�U�] �,������uއ7��+eI7�U?&i�F�<L_fv�1B �� #\�H�6o��~j���p��*�>��t�vn0 ��VC��z�ǨՄHP^�u��ZEا��������bb�o�����Μ�>����C.�@��9C%�Y����A��r�xU���'���z����{$]�����8�j��s �L`� (���O����&Ų!&E�n��W2۞�w�1�s�ѷ�H�yWJ�e���+�P����`����t2�2A��/�]��@ED�a�@g1�������o�5t��YI-��,$M�QD���c�AJ$�xO��C����T���ka�U��\����)=������z�Ƅ׻��h��a?"�\��8Š&Ijz{D<��c�����a�M��o}�	'7Y@k�G�N��м��h莑}���Do��`?y9�Fg�EO-�D��=F�<j֖.�(���7�1��i�=z�+z�%N�H����Q��1X@��9?�a��
bT������ �+�<`i7!��w7dc���i������ʠs��B���@��\�n=<Uz���������ˮ��ђ���2o4v�a�����-�����Q�|\���\���R m���� ^&��
��ၳgQ@K=��lA���j�!C��y0Z���<#l�O���.ˤ��ؾM⚂_F0<.�����ͺC}�U|�(��cz���Im�rq���5\��M�C8S�%Nvheo��aeP��&�Pk�TCd�.C��ϵbQ�02�>��@iʃr�V`1:Z��;�����,��������Cr.ԼW���=�Ϥ���l�=����k� )�*"vkH╗]�,�۱�	U.Ƙ.t�8C��\�L5��EC@Aq�wJf�t9�3�8�CUDjTvyK��ͨ�0�=]�J��k���'6�bG���1�����;��s¥�숟W����������$Ĕxs=SO����Ǡ�+��/1����Fv쓽1;:A�(�se����w��$� lD��y�{^���֌ڨ�2�a¥����:zb�)&.q�\�ߝ5|�F=�ȀV�m�p ���2�o"h�����H7�2�� ̷����1�kPa����6��Aܩ��v~*�47�2,�3/R���@�i��`��U �&��s�����{Wq~�Tu%�Pba#⓴Qא�v���7,�un�m����@i��m(���6��b�(t�q��y�X[�ܡr8j�U�`�OU�n|�9��|��d�� �g�|��)�����~a���)Z`�P�����w�a�}=�s"'�X�a��i�qI=���׮���x�j�V�*2�s�V�@b	DM�~,~�}�5��|ر�,)�ρ{#ߡ�%��w����?���j�h}�	ʉ�"���(�$wX���۬�P�o�Y�Sf9�k{��r^�C ���w(����c)�³,���r�$��g!!�t��[>\�u�޲ք8Q�V�-l��ڥ�mB���CE"c�d#?i�ݨ*"��l���vr��S���?�#`C����5��㲕곐㙓+�Vh����M���Bᖕ�e�'3��\��B�]>���-��g�4(B݈8��/�Mc����g�̔X���e�I �%��$<�X4���U��q�tY{���#p3�>�ת�C�\���x�1�
���LL��N��齬V��6��A����/��x��Q3�MB��k�[T������wvan������� ~ܱ�P�!n�-	��lRU�c���(�ǒ�m�XǗ�1
�͋��cI��p��"7�;���UH.�U,��.XkÜT��17���h@~�w�0��U����C�	l�Tj� �l���9�����߉��pFv��~�3�u�y�`K�R*]0Ox��SƖ.�ː�(��m���"/_��}4��d����d���Zo1��?����Mb!~��K�0̹�%�(�82�'Y�>mͅ��!��!x�&%z�߲��a�4���L����w_��'�c�H��6R��d��'׌+�%~�j��<�+����k~�9k���\��WZ�V ee?����\�K�|K�Ka���4~�cY,;0J��ro��C���Uc���R��Ջ�C7J3��k�i/?��,"�Ԥ&G��[�R�
��	[�Y��N�$�U��REu���,`�O7�z�F���7g��`�]OQ�JxID�,ϬJ��B������袄�����j7�ո��i�Ų�c����QX��Ц�Z�>g����;��Y<�����,ذۋ���3�E�vH+�D���q0�r������^�;*���7mR�8X
:�%E��B��1r��/o�n6K\7e�R�Kǒ�8������~f�~|�;28����D�A���/F�->qPdyO;J�7�O���R�T�(�`�?�D4!:(��;k�����J��Ir[��yv��S������JzǪ *O?�*0�L:�7�4�O�.�O`}:F���)����(�]>�Y��:H�Nƺ$�@��\��A��Z4��1�m��{�Dk״<"���B8�˲�R�@��4}x�Y}��f��Ǿ�������_���Y���T0^I�'�B�V�,Q)�7p�<:�N��
�xHг���)_��~D�N�2��ycn��|g� �FL�O=[�Lw6V*"BB����V���뿯������ty���@��6�(�e��(�{��*���h�� �A�!&�g7�6`{#�"├(����v�s����[���7���M��l���`��u'I
�-��%+����o:9a�����!jCD�=����
�[
���i�`dΥ$����Zx�jn�.�q՟��E`fZz������r�&�cm#�?���(gRTd[X���B��~d��^�������ìz>g�I�`j�N�w�	\�*��8�GW��|[�Y��|_�ܵ���F����m0}G����ж@�����g_������1�N�r�0 bk���C8
�Y1,�ś�U����ɨ�7�����!��I'Κ�v���L�=g�U�_Q�w�^�����!�c��nI;�j���-9�nH��3��ݗz�q�[h-P�7��b?���A��]�@P1�|���G6W�sPw6����h��#=�RM8���/i���iy�����OHOe|P`��L��{ȱ��k�����}���QUL-�c=�7<���U��.�e��̨2�T�U<3	��^���FI�؝+���T��f�e;/�0���8.q��]��T�B�'O���^�$Y%��)'G�~����_�]��+��BF��T�Ve��+��#�ۄ�����wH�m��;!Kט���O����w2���x(i���@����������i�� �ʍ�]m5;v�T��,`���@��fa@A��ۈ��Ճ��Y�K��0r0����m�ˠk5�zq(�c0}}��|�q<�Jj{�WSU�Y#�&�X�����%�Q�T��FʼC)v��'{�/k��PNe�Ǥ��JZnb�}��QA�;��#@�c��E�}�?��D���h�_��@�`E�bu�X) �@�����V=�p����kk$�w��;���� Lc��M���QT�P���f���]?�ŭv��Gx�%z3�DѺ�/e��4}~v4��)p�-u5�=�.7PQ����E�RKOA��v���7?=۝��f�O�gZiZ�%a% $��%�aսĎj��z�$��ӑ������;����`o�QX�w;	)ڲ���,�<2\'��>��@.�X�����@���z��=ȱmzư�^nI1x3��N:��?�{��.n`�=Co��@DH�{j�T��m�&0Hɾ�ȅ�#���4��ɑ�.\I��E�i��GqPU�y�Y,d��erۡ��A�͹a��iᓝ)aP|�+�|�/c��a��d2A4��ߝҖ,o�ωힷ��ԅ�����&#M�����
W��$P�&����}�|�,����m$����!����ls�#�׫/�D�N��c�Za���J�LC��l1W"bᳶ��0=WA-�����)h��	ld\��I嘈R�0˜��O�L C꺶[�}i�Q֬c��5�!���!S�1�k��P���ɔ�ӆ��w:J��S�'�<� (���!�]LF �5q(7�4�y��%�:{�����4s����h�@ B'�	d����k�����.����0Xr���Y�Vq�C�}�RC���_
|�|���V��<`;�d�I�Q���\��Ѣ O<��wJ��3ͧ}�pj(l(\��ZT}3~�YKS:"G��";/t�z�~)�9��(1�&+H�� �d	� N95�b�)*�2`�8T��Od��ʅ]�s3�E2���H
0��Q�g�~�(L\�T�k���׻\��JGS�p�F�`�M�P�	���l@XF�H�R����G2q���H;�:�} �}6���+?��qS=n�P��M�$1�%mȾ,w6Q	�BĘ#�I��8`�88��O^�gCz��	�q�U:4�v �+��籓ӗ�U�Z`�<����_^=�@"�-
�e���G�1����:���
��Ts