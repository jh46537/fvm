// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cii/H9KrVUSRoNv8fZ0vLfWabF0S1f0QKPszlV/Z/CNfTaZ6NSgfH8PRKG+B3VJ+
nYWFgHmRZLrPhtQRPfcn8liaUCncYqdsij5dCnDGqq1Y+zDjUW3Ph6hhJkUn8QJY
gi3ZdHOaS8Xzz1jB3W/tm/dYiYRIK3FyfnjF6bo8/YQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8992)
ZbEir7tHSSf6ZPShYD09vjXsJXB9ejjRC+p39pm3c69tMe9QDQ/U7NEKAYaLK0/4
Xqx2VJRhWsdOvWuPW8T6xxSK5XDCwtgkpO39MCDN1128dqlysAer72aFR9bn1QeI
LAC+JBmS13k6WkEAhuZwN5kI93hI9qWvhTN0XAiQ6U0rBseQlI1m/CnSSQiKYAst
Lse/As2q2uC/OEOS4ntP49gZ2Ry4WrqeR8pqnV4JQ8A5mc7RCqTaxO4oPJg1jT2Y
TQnvjYk/od/J+JdjCvJjfCVaqlvGiP3fziMAAz9oybSiRULz2vADQ++x8gGwOOVv
1+hHdMtRxqghhdOrv+ccXy4VLtaeChzn7u77/6VP9ooM8YvagZ2RM/446tVT7ktf
JU/hwPMwBbIWtykZ4dpS0bKr0HCgudLaL5rt2N0QcvgV64HlJrINf5l0d7tdUaZB
B+jigoMaXzoN48Rmaeq/zKr/W5jq1Bdig+cR9LLxNH4ZlbS/uXO0VEIeYS3QLuOI
uXanZ0MVwkCdhel2FDzqsPfnS2fq7JnjjC9f5aDW7Wj/pGEsGi5IoplsPzxY59KE
lRFw3eI84eiP5fA1I3lWzqBSFr+ioAtPh/5pxvsX1NJ0OP16iLkO5+/Ecvy747vE
JxKnX0IoeUeoyDOzX+2bN57thPg4IjHT2lAd32MaY0r4SssrjBwQ1UdeTYha2QzP
IA4aPat+F0PvgU3CmIWhCG7ExeW65mAUwKpd8DB9/7PbiQMgS2YYOXavye3PZ0hl
UDLoudjMHNIfpuZA+Ldb4pVBWdsPITcbdNhlKtn2ant0kgt2zrWAij+WzPizaAFn
BwaMWpdMdQTFb5aRjvrQiHowaLpZ9RJ4SrgiNBLCW4YN/iI8X6D19msNIbHasSk3
yxyx4wGUeSNJrxUhrTWjzE5yL3LQlgEbW6Ik1eC/Xy8EGf2pxHJggFd54KSmThTe
C7j42gSQs41RIlAv1yTfa0UGhphhVcGQJMwwIdlN77jPk1H3/yhU+ADhTePaZrqD
TKbNS2Q4r/jVNhOe+RrsRaSwcjO2rXs1VvBcH3VUArGS4YPdks+ZnX6Uusq6rXOi
3y9SPyAvfQo7vy+7POIGfTNSTV9En14Gl7ejEt4u+zQHPLMWiJ9VR645Ot8hawEf
gsoAbE2cGya+UMUuQfUsVnLxjc4au//daitVjDUBNTmA8o3bH4ZYNSRaXtdZ815z
Ka1VtiQpFgzbfyVXh/lvsheGldvyTH7oTWFLDEia4PDYwpr/9Ujjd8+NHBqqlQsR
c3IPMxGAeSZPlCQyKddpmEiWKaAsUUN2w/6SsTl/yJaw1GEdRawMCp++WLVDum2r
w0A+JGkSb63dth85kxlmwEaWjJIKpm90iIp2cIEUczmnzDkp5HjJOJv40lPOS+KS
xw1Y62rRFZHC05pLuC8vMVAiRoOvGrWkZ5vHXHkNExmMLDUE3fhzRA6mv/odvBp+
+kHY+VTDz70CFEXxHqPAIrm0PwWqrCIkIIoJ9JBZoBEYQlk2xQigMkTzNE4q+0NG
BRfzUYC+ma3icfs8kKi7eP5kaOVAW9Yr7P7Bc64GsKPPCAYjXbvtth2qKPYfix93
gxiCaZU41gE0NsGj/1mzyuvgMGzK8jG0L3MlgzFbu187G0RE2b8i6302iNm4fAct
1dnmPqrQ6bdl7SqhbBcyUG7Gv8nkyB//ZVWqx1Gjz2jpqEijN5cRLBu+J0B7Kl3E
HldCJJPaEokiNhGS6Am2g/g1ammQYpc/irLSvmSwkSbAguBF9sEz2b/ZssISBUCE
+8Pan864oKAxEkqXNTk1qCLBDoEhg0oCreBIwjkTVXnHMLhFaCSoVxQKTqjhG7Xq
AsImy9pXAjmryj4bWPG5aFCUcHshZp8KNUkEIMsYZYp5zbGvyBKVYf9zDJeJq+9E
aJj2367OzQnwDUTCasIFzTx8aPugkfZ0JhZ7OJLbqvxwXJS9UPG1lTdLKqQI+SoN
gHRYGBS8r4SvAdHmjmelDT+kntTKj0hWhMdHFgMH9ZbZDJNBkIoE4ovk7G+C3EEr
mCUWFyq2uiQq1mTd1vv4E/4bdPFzp9ir1dOV4V1X1iiXHUvFPqu9FsJ+3Bl09v/C
QYw5AiH4jPhrVYqU0+To7ejYfC6FMFDrqh4oZzs+NTIpwePKtOza6c5nhTMJY9mR
Is846exooXADyH9OleKWGjvSvBtD72UJ74N83TmyidGzHluf2J0AcU20UACfyvY7
bcysKY8ov1eqj1EsGcVN3ZHnjayvl1zl9+H+kQthqducyOYqFpXuedfoef/cFnDW
FWzrupxpbvafywe+w5NWQMIXZZaGxy9OuHctWjj+FO1cGXV/5mNCN9tWxIIOdhWT
gHGRljHp67exHtKiTGY0nfbtpTusS2mjzLKCsYJEl0b29wXW4hP4cSbTlGgnz7z5
vEA+0AtBPr0nJfo0tmWRKhQShMBkpBPK3LAadIhT5n6hlOd2ug+N2BkY2QRLHp6Q
V3PO65UubblstMhN9NuooOk3HJhli60hsRFGAqGSVRumVTTCLMaHlKlZVyILQj4T
BJb+0l7hn8nTBts2SXJChF++MTs3CmH/OElenkDtY6BENNC0XKOyP9qlHmp66JQo
hBcjEV+wtQxUKRgHwXKeJI7BVC/3etWJB6BskUWfUJ8Bz+yG3yy9qoSY79OFo0LP
sRc8w/PsCMVq2G49FlDCZE73UpojqExTFCeD3dA/v5SFpefMAOklIiXfaBUq32Gd
Q+Y/vD58uAwBWD1ISyp35ekMsI4Nr48PLI/RkvwnY4xBeEh/YZvnGpYNdGqxxrRz
l7vd4XuyZowDC5fABDo3Q8pal4Z/JEZ9DMHAcSvMmiz7tCT5K+zBxmxKwqIHKdcB
qF9ZEToBc6S3IJvQaK2nyxQaTLfSWDnz8V24cKWgWl9hq4EkJ3YbnFRZph5I0HzP
/I7ePX1dq4FkVpa14hYEPFtEuWYtykCpQb9qCbPOTXtNEy9ZkOgeLHZNSW1ru8Sl
ODopOtS5Plbcp+EzXPzxnPBJfnXnozZPw9A6FXmL53fbFolsaNwDViThMKUzZQwm
SluABaifXLovHno+zxXTaP3aqsNI19YhBtHzpKsN7ClKs4bp/8ePx7APzhO48vJw
nYOiJqsV50Nos40Wbmy6FDqW1IARJPML5ksAF6Jmk35jfWo10NgQJUHiFUOaRlLY
H+SZxHD4XA62srlk3eM3RuR/qX9kvAeX3yyULLgF3AwYaiwMudW0XkDOaQNC8bRo
quCtx01rSxvZMGeVEzQBJ8I+xuLUZBTB0iAgnHDV0fDgeUF5pzQ24lmFdcgvbLcq
96+e5cfVCojNXbs1kho1gNZdqT7d0YNVBavIAzfVLSITCRuxk2JQgoFMJfmB1U6G
BTkf2hhOYJh5tNvxrrGtZdsoHE4ceYoMv3ZbXg5zOy1P8gVNp+jHK4c5rq+ry2fi
ulbWZYQuVw2lWSTXlwjBBskjumkVdlVrDS73xxfzwCcxmv8BUzujsCUAmIi/eOtM
T5GciBd86KPhvG0XunHmuh9s59HG4BKtmPbZ4co+28y/xE1kXU5NyeQRhRAptuNZ
wowuxXtubM5aUZLpZZ0vpJAzRkPqdlJ487F9pteYmULb80WhQHLW+bUZJtbf6v65
8BOJGpfBloYnGXUOBGl4ucFM47gJl7R6gsuP3tyaYqC/wpmzKjiMjm0oaowUj5Ou
71cnqELPDp4x4vmhDu2+CLIaWjeS9I2KW6MrwVLDlFCUlMThMZ2X4zWLBJx2O03K
Ag5S/LOuiCXj8hDtdDNnOZIg1lnXloiHVnGRodFFpGpRQD49Aqjmtrovhh5R+Oqw
0Jf/v9Htla+KJJRyJvAP3WbQ4Reh2f7iD293SkI+SK898YCXuw49e2AzA/n8fPtv
ycm7po0Cs7rcgBRhxvRVj8b7p9/G0CYxfTMCzm+c3kub72AAOw7S0SimtKf77+yS
MwANGv6C2juzV3z5BGm+SX98nTthI/Yp1/O24Mf0pr+W6VipFjtnD6Q2dBil9pEp
HH20uA4Dr7r5mc/yc2uTd7JCztl80lBuKAa8RhgHaejED1/3XnB9d43dJqOwz/w7
RQES/722++BehwshrmSltaIHc7lY6JjJASmZslzxscTSFHfW3nUMW9YPx2XXvK3w
pYx3/t29MEiNnR+FXQbEmW+zz+IFp4JaVjxMmIA3oV0HPEWkmTbBYE0qdjXra0pm
by28MEY/oCJB6BvTXg/HtXD3csfkq9XdpHPP4eWEP9c+jiCBkuwAxftpmLR+wU5P
2h7+Bpad8ZO0vUXCGXhNWay2exuCQSW0GwExr8uMrY8ASTMioQsVmKZ3lEnF/v7T
aP1lnhnKBiiqa/s+Y6wLucN76DnIPeuquTl+XLK/okBt1aqVkyEyZRPYTZ0M1I+T
D3YnSi1fnPVNB23VdEMdn+zLi0G7eMcn6wKwWNbt/kGgAoA5G7IQn4a6IcgyF9b9
9H8EfxVySWmVeKUZKTMJH7O1mJRPRas9Uxd63bgTUbAYc9gkRRj+b/BE8BuGosgu
O8rew5ViX1GrFZbp50BVtgsaue4oHTI2EczInHeDcPZYm6lExqSVNKq/IXBJYDIU
3jbISFKLOIquIEqT5I8PIZv2SWATecKeH+dET+FwQIyYHsmhTYOGtXkioiyebjj1
Sw9YAyFkd8UxVSs15+SjdmhZP3h7Vv7nVhElPnRks9/ygOGbmF5wBapX4T/fm7dt
KraV6CJHs3zxbkI95l0TH1DuXoyYmUtUe0b26SurGw9PSYn+s3UdH7rgaEHWc5WC
dTF5MkANE3DO6JlJvVZTM7FH7RYt2CeZcy4mp4GKyEa7jyR/wFq68t2haoBZipfH
/HBOcwTlewofS9bwPnfu0zfljNs7VzN0MIG2Vr3GU5j+inXGIB+fAqGsoKWhweer
73vy3ArKha0q5Svz/SyRdkL/Yi3knEAtSUZGv1RmqLlD4AvskgsDexEWas3x0VPf
Bf+5LNr9OK1y0WxtyFjWRbdbz5bxHnqb3nKs2E5z0ESWalNrB2IYi6PZJO2OnvK7
C6JpW7cHlMZxQblbiEumIgHDEKfRkQLx6oBJD8YQZH/6LFP0RqNDmAUkxZUhA3fO
PUvHmNO+A8RYpq094fbNhie4/XdAsT3dkt1Led/xWojA1jEXOhAiw0gV9B5PYll6
UY2Z+MbqkOl9a1bRdZdfM8Fv4Ejs/t4A5RoMUOhRR/sHl3K1AHuj88w1g/UQFGr9
4e2UdBV+bjjeL6ab+cErtPd2pvQF35+p5nfdO0foe9QqfBY2Gd5PF+c3/YQcV1nQ
Neel3zkDj4wcrfD49Z+4NzRoRB2KlA+f2MdmRAjbbNrXtT2jovJ/nO5pHPOKRxvU
QWLqJ7//xLaEHEkJ1h4BXKx3FtOe6aq4Sl9/YTe/7K74yew+e73IqAaIIYT8gJN0
GWlhx9/70NT+zoV0qnD3gNmvwutNubjS3tgeveciZyUxvvLwdC2ySd99WOLBAhTP
Hep0CBVzydGsZQWO2xfbOf16rRa7qjAEXrkFMoCl2NO0dQkVoeJQBl/csTt18nm1
ySOLLTb8AmZymrrS/GabZ1basYrUYR520DwFRNwWpLyzRs53aGoASxLmaU5hKY++
/IJ6R6FmOKosm/0mUgWUqOOgRbWHSncyX26UdR0xTXbAt1QaS5msbh4sHbyRYy/s
/WrJIX3HvQ+m6eH42cTGZOSdwxwCsuZ00NeUvSIvGjp7BwxPyd3R2e+nr9AHbi62
IbewDb8AxWMbFfwWKD6wi3VFtH28qLIHKdEo8skUCIEytrujtIuTZEMU3cSl7E/w
b6BtQEmvxG7vW4cXmnpeYLUq37C/tTeJENjUvWiKHNjz2CuTfkV6nQ1hsFcG6WVQ
qNL/V7FkX0RGAxcYLPLP3HZVkKsh2jkYuTeM+qrADl0gEPOpiaBtXLT3m9znBoXn
x9vOHJoobsOy/6BTrx8dejzWSmB/hQLpzbl4sJwD+yBsfKZdwZJ6bmsmg7Tl/jyR
4T75h8g4fhbMigyJbM53OxO1dcgbB08UmFTGoZpTk4kRfBk52EHRrTUtPEmkuyE7
1nokDoDhaa83MbFkyaKRq4uULq9xgIcppNBsXf3ifKKAPg7+IMFedJO3/ouXV96P
8BNnPLZFeANg4M8SGJRxcZyw7eON6TUVE+MQJ8c1dCnKVjmpQswz1f02SDEPRhmt
MLireP8IlbyIFlOiz477mf71Zg2AJJHxZTe9BXGNewZyAPlWCx42Y+RAIVPW2xRx
TJFcXKnZ1Y5b9aUAi6emlluP1bEdgnPPW7eWBqRp9UwpbusqG0CVZG5HAq8esB7w
L7Lpv+Mta2NmRQgxU0TNgy51LscPBU11Y3VZtMI3FkRqpVfY0wXeniKqFMQQHh1X
HYItErXuBaPToqVDOuh2v+LTslZceQ0d9bdjWJZ8QO1MIkMlRDNKoDPNjAl3Cia3
3HOO5JIACif/vS2I/M+5RfAOPhhSDWaiSSwB/Z3LhQsODBxUCDdvCVSzumux7JIV
WodDf3EPUsAsU6J4s8GhnvihbXQQ4ohh+5nLynb/LFmVY8dOO95LJFHPN+GhA21u
XEJEk+Ht+Xf9P+f7+W1PZJNjvqcE8CV71mfhb5q7OoWGS3SiswEf7ZSaVGyJQyLn
yMlWrHpzeow28wo91jGI1d/BPStM803wU15NS7LLByU0ei6A/PwjOougsAR6qcv2
ORSJmy+90IasGIGfSZARtziL9pzO5oshROuQ3uCa7b4fzSVR+NbUPKcyZhOWZa1G
IGGR5tGocUJFjgPq6OeEuZiKAN+UaIE8XNEb1bqzTmby/cWOYIn6v9GVZ0qWsZNw
ayOfeiwhWDkGJcFzgZj6Tko6Dn8rlh5NOJfitJipG9c5VPHYZVKXPED++SfrS9sA
oUohQUrS7LeW4oRULsHgIeZUQ5zEN6bu1TbRognvobS+R+wHvmFyCNTLd5Br6Wpx
r7GGyp3dAbONk+gMkuGMhisqVcc+fF0s2Izlklz9xVsZRjA6Eil6IR7PjCnx8W66
4Zt2dqcFt9wnNaR4ZYVesV4Q0+VID5PL0B8bfV+R4rn9FBibYovfY0sRHcsd65Iu
XLTvBwsxbhAWPzawGSNKRwjh+ZYUgPeykT5+VlgCB16aC8GdAvkGAXBs9f0R6x2I
hUwKgxed9+uV81XQKe4W5qvsMbZUxDCv9MpOeUOuEdlEMoTTGRdoOLXPlpMOnbE9
V1tuP2zjbwuD4Ew5Y+A8h0jC+EG15RgRZeg2H6r7seq8vc/7EnX7ExWtAk0hoJ1V
wpYFlG+ApZ1c+pbDlb+3pWynVjb7VKyPtfSoTTa0Rdkom7PAPHL1aTy1rBNdFuyM
CdP+7oD3TMp/dwW7j2cUOSqjSvNqysLXW6G96pT77hvmWv6IaQB/IGE4F4qST0EM
yX36KeaKK1aTo6xDzX2TueEyi8iEGixq8XQmlDgwJhA4V/2XBhZzvsMpGTaIaayt
wRaNhFw+C0kDdB+YXrGksUjibdnguDqiA+YeMdATe63YaL0s+BFXi4HWsNY6EWWl
GcQV8O/ud7rlpsJjvNVGGY40SrcTNIM6QX3pJgElFvyOLBMz+rA7s0JjKx2jtVd6
7bo2IfWMUugxEx5OBudllJMAJYcLYMZHdz3194DfRFGcvTAwaEZK+ptTJXXZB4A2
6jWF3ftYhBnlwrByyHTt2ZyZhhldGEWK4q3qJ5futVZqlAENQEoP0mfoKn2aBDVX
AK0Dj8ujky0dVnISlqRz1UbWn4zIUQqMq7+WOUza/V7VbeCIfcPESeVKXuOC+yaN
hyAxb3rjz06H0xdcBVHYE6Fm9fbQJ86ArwpCdXrUsCnN4b5nOA4HJ717KygoRTG8
UUs4rOuqUhTdlkXSJjvaTbqLyx9jBCsdrz69Z+0ZNXGu/ybGiujXMZmhHP3kY8m0
SOc7EH64j2gEobEY03ja7eBR9hifM6+caTfDQwArzX/1MIHs/bwkTWbgyDqAfYAd
Qrtfwo+wnmN9fLALSJt+I5LaMCVJYXRFPSwL1kLnTeJoLIbgO1ueN9Kev1ec23FA
Y806nhnQfM+4FjUk1HOYDAjsnjH1DUk9L3c8tm+4O8vDA2O4Q5UD8getCp0AzSRS
Ls6hX0B44ZovcYPBOS83fVmmqB0NEWrsfLxI96TdhE7NsKbqhHE1Hl/JONbjC2Gw
0JMWpBLv4Aky5GlUrZkxmIqZUA1zmAITs9Dnwrr1zSODOMn9+x8e9uAr015VHRtz
Ew98qZ7ZRmrVW4kFbOsm6ALuToU4C6777WYRrmu4nqXY+Z9mc9rPu4LF2g7XP8PK
H0WVozxFCGrflmjkwOIc2JpsL+YGt601E1puvXUvixwqROPSAduCzn3Xkapq+zLI
Coqq9s5j+sG2SLLej+we9tXVpailjv3GodO9EWn+uD2Cu13ect6k4Y/6xZNogoXl
TID7GPdWmUAOD/r+JOxEns0ikmyC/QOhFMEReSgfEB7BYUoVZaIVVGcR+JNrNyWp
fFlA+X3T9k40akj2FKO7voXYv85cuTLRSE9fp5XB7ibZB7gOUFxQhr86U3fpnpdi
Vjz60mvMaHkzQXyhEaG5vVcWq/dtSNiamQhKqN9welFR5Wr1SIdj65vbuXiPXFuQ
vAIQzXb29mvtPcTtS6eM5aSlqb9Imgw/wKrjmZ4N7vAq1ZTKiOOiihXfLa3AJo6N
D6zIHRHN1MUe/7gcBy7zGitagRbN1eWTqLvg6y/7e1S7zZ3sMmKY+B4vv/YE4/KN
wq6Wkg07xX7+Ys0usBSrLq9vtf5iuU5kY8JouFKGB2IAYmvMkR9Jxl3DcEbj9Nsj
J8mgM6pA0cx4JK4EozFfiizrQlx51uT6P5pZA9Yda9+5ANFOy5B8Y0/TMZChPWRm
rWnBx0cLnS5a+Oo6vlXSwqAA7l0Zw9nQVfCsEB1lpetoWGqMiaUeD6yZmxFy+JyS
gOfAcpnWbrJQyzPPSvcumbax8ydf40NyeIj0lfcerprZvbe23lZcNr+LO7z130DH
49UbHamMUzAUPKUOqnDDfE7XxMPPEotfuD0wkSBNEXDtQ6iLGjOoweY4NGaUame9
PldNvQ5WJT9AfFxMbwP9AMzbrQ02QwrzHjcYcFHCDlAM0UU4ZHwL1uceEDnTVWu5
EMnTfwZNT8O4s9aFZ0CjBlIXK7QnXzovyhJLydQMKJl2pxY60S2hla09TE4lqLKz
ZGjtPv2gyBKxJZkb40m+GLtrOcJoFxSBVPT+cGU7gf0aikDOqJe8JptVdoHRjCkj
89YFkQfuXux5S0+daihWTq1GTt8l6QlUJN4zOa54ETG6mhY9G5xe/nmK9zBq7l6X
rX3VTULJwQGa+VGHqytR8lA++Zp5XzW8I/LuP7OvxtBCkQDqirQhFJBL2oFZHEDR
K6meqyHI2CxqxfhoqIm4AUpQwWH40YMxbHOqiJHgfcazaChqBT0vtk2eH3lA5G/V
b5WkWvPUCLQE3XuN41Yfkd0ECeYwWhdPe1UCU4wNyyp+Z5RtNBHtnmHAlzzHCTP0
eJbva5DiO/jmy2Tcvu41+Ghag1Cs6dmkg3/dBY/bNpTRhR2geF6RfTtToHBCoIpy
7CAY/B9V4JRbt3tdEbia4IB+G5Ki7bxe6omANZNkmrusU/SEXKnFmWBiPBErtBa2
z9YKFyxwdiCS6ek6eROdAePl4NRgEF5RZ6Vh4HfzWWxjMbb/b+a3qZj5Wo75umWC
AIZoJwnXlfqIDE5GXqHv1/wkxKoHqJ3oHl/asaRMD2/9zozkomsBjT5ojFXUDRqK
tu3FrGLK/Hpjv0We3pzO13dyyiFVOZOpUwBKYGQColdPzwnD6qwqnPrQOVfRBaN9
gzuZtU4Q13tdv66dph6RLHfq3I0JRHEJ0WD0zE0AZ/jkspuWIhTPqoObaWcFsi5+
KJHx3X5+FtEqMIjz8WdG6TCpYTYBOTPXhyVpxKbbPUhBazgSjRBgbC+mVxdQOEd/
4/yKWp5XK6kgNEGl37xVzIk39nIYiflcGJ3MemEFcSOIeSJfV5w+95g6uq+Fk5c4
wdAo3Dy2ROq9lDROANjMNutHjijh2Dim9gSSgAxROCGPBHS8UzcDGU/cRChhJwwW
CvJRg+Y2TTkvYamd7kBG920yqXqyoFH51QmPwoJAUWPWUyL5FNn8IEnR+PQlW69h
EgJOuyxzKh32Tv9iH5ySt7z6gXMNug1OafhO8MxOOjYzvMG0EI+/aOo97jSgjD2a
HPPlKwlFYPOowSCxFq6o4Q8aWa5Fm1WvtZnPj/O4dO93/MiyjVnfVelv1BS9Hv96
fNEnUE0SbPxesMzOynYMUoqaS58JPQTHgP+rNvdW9wijt53ADtY6Rb2gquDnxsOj
gnCJ2FcZ+nUynUa/+zVIMYn8pKsLeqrwwJfOs3epKmrzeZ111A6uORq149ea604N
UzTWhaoI+hE1+vjEyXWsDW76x/rDp8ZCHGpV4Yk3K40Bpm83JKZdb9WhRDm4rfJ2
Ej0GUoh7CuIiOIoDGwLxDmhSUi6yAiRdb9k7qVM7QbI4+W8CWeKzDCj/4OBbM+Te
n3fAAI8apZhYYmXTyTTqVtRnq3CG/+KTWnpEmsW/b/UwtTVMsB9zgcPbVnApqGiA
/kaSToI6Otd1ixCM5MIeYwMDtKev5URbET/TOnnnRUxnDXS7d3pohWA9aZvNKlo4
teEWogz9Xb7QGeKPT98RMxyQFo0DT9/ROiUjrcXJoPLFjRY1dmKLNCt2VU6sDRmO
u2zD1qCJk9PSIQfY3XqbeN2fiaZYXJbC95AZBA/a+LsadZFeLVREgSpBr3n24TUg
7Nht6EJ1D8L+TutSG6CHreeE7sG1Oh1UJf3oE0FMjBDTsCdGUas47lS0YHW7lgbN
UxCjadN1s7OM+ZyB8Crooqo+AslqX02k32rzlLi+eJVvdtl2/5aFVu9IUO0Xq7gQ
JiMu5wAHDAU5djJpSNLQ4UDA9R8K1dDDkT6dVFaRcORIjG2sVerFEl7wzX4zhPXy
SwcxrK3nK3/jG1D7qgrRsuvw6y39+zurGmzjra8nTwXz41RxO85f5glWMZYwCIGR
EuPxdx/mAg+c5Uo1OvkwzFs3zv1AnOf7XBFcY4JpyS6cFu/YSfMdItLQhvaWqSuD
wsSmiio5SoCjH9GBcktSkfe0qePucG6tZhPJsVcSu3N4nBTveed1DQfGr5YswRxl
uzuov58P7xtUTQNMKJ0JEfqNYh//IRI3CVCfs54jwVkuZFRNZ7/EuVv+kbrIHrca
Z/1PHDOKPWPl535fMHdKJBgOTL3K7FnAfd7wj4AUz8O14tDdQiiZBNnm05IDhJkj
YNb0ZOnpTNfGOaC3Rc+yn9VPO4SpQpiFav2QgkCMLE5L470wttmfihWR3ma3skzY
2Fm5IlCCNSd3cbQFihkWWWMC5HKEI8IEhCzcFcF6u6FUP7xG4mKg3G1Ax4hY6Ktm
5v3EH2JEVm6WxvAJtfP43Ia11QuqLSz07DNHbniHtiy8TWhZ/Y4mMZhruJjRJiIU
V4bVTUXwo2Kh5FKJ/mPIfhVLoxbucaS3qNnROO7+NgYSMb4XBplopXABBIWrYbSD
b4ce1w5riA5W6abmakOW8bIifq9suqtzVI2yGllGSIvyZApCdhSo1l/22cSyQiVo
uh8DJyYfqafo13zdkt5H2sNbCoDolSp7mnmz9a4/3Ba34bL+ApeIoqCJw67+cIKr
eeZ/f5iLBmm/DNUdn4j+mACHWk96ONqrEojMc7ceRGjdDPwRCHzgf8+S1RtodYVQ
7IFAnd0zsREFONE4nFvmXDmIHpS7baOCvnPCaM/webVeabr7r2lf/W9KKXxeul4i
9RwTyd0wHdyZNMkJias3CmzL04JSAsdMEl9CKuWXw//8z9k9poTvsr1GNPYd2a4g
0g4oYhFcdInKOf3BzjnTMrhSyHvDuRMryMFa/UaSpXFnFJ7iA6HGAMPOM8YblQWQ
CQOJrCX1XeoPBrtjjece/g==
`pragma protect end_protected
