��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]ǂ��O��˰�	JL\=����"pI�: `�r��+i���B�Cp���,��1��o��(V�M�`SqkH㵊Kp9�=�3�1`OE�'`A���MV�������AO�I�\;��1(R�9z�)2ژ�w�)!,�:x��A�����o����;q�����g�ļ����O"�jb{���U�m ,zt���Q�������yAR)7-�#�vGCUÚ���,��˗��u�r�zE�ρ��i�g	�E��e��jk�#Q�\�W�}Ul�G���CG#�`����7���D�!�=�l�\��\����-8u�2_r�M\u9��Y�[�A��{If�ؗ��&X�����^uw���o���\�\Nm2��=���n�&\��b4�mN_+�`��D�>��t��.CA�}� ��oퟸ2���?غjz8'WD��Kީ�I0�H�0��H%*��4���