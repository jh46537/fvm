��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
��䂍F3�`�Em��IL�t}�4WVn�r$��Ӓ��dk�U��U|�����{ ��s�z�~b�À�b�L}�,^xt�y탄�9�0k`۞\
���'�lO{�P��f�g7쿜.���,�r���H>���W��+�;�S(��}��V����$(�xkO��ÙbR���B����qJȬm�\KB�5f��-8�x�@$�ߗ��h���LZ&U�/�����6�U(��/՟e�]D(O-Eܫ��[�e+I>�OY�ᖧ�<�)p�?(�{����õF��7[��
��N�Ñ�B�l�]j＆z��[%H�� X�,�O�� ���V�D0���{|���Geݿ��������om��)}�ŭ(�HJl�[�NJ�7x��b�;��u8@�="Qf46�8kĄ}����e���8-z�Xb~y��� ���QW�+&�z��Z�u�)A �1�\;[JGq"<8%�$&�O~��+d��:a��r�ގ�<Hw�3�Z%��py�܎[j�P�6F��e��)V
��y�xq?iK�7��&�iߗ���5��A��Ll:ki�E�ř�	Q�����k<���3�3��ݦ�;l�Wrl]x�o��#�V�q�]��UI�
j/�?�j�wL�}�j�����X˿�85����\/�p ��YƋ?A��u
~u�J�u�_�1�[;R��g�~������Ux��t�[S:�D���5�{�?�
c��k:�G���Z������Ԧ��K0�?��3`��W��&Ѳۻ	���b���vpz�J��Q�rX9m���Q!{�UCˑ'��$��2�9M���V��٤":O�5�W[��;�%Z>���k���펷�X)��4~��U�u$r���r�V	~j�3��+h��t�1aPռr0��~sQ@���K�90��t�w�0)S���%L��Q��+��C���=�D��dE����*����=HXB{�y��� �S.ұ�h���Ev���^��|�^N"8E�(�V*r����Dp�"%�ə3����{9�����4��I�;��)�`���3[C��6��#�-"����6cwi�a�QM��ę���S�l�g��$q<o���#�+�P.<�� �Bա���}��ȿa�;o�a_��#���k�h�,�9��P�5M<_\�B?W��3�1�Ԕ�}䑚}�=Ft��J8j�#�t�'�U	X���]r7+�r�t���ے�-���Y'7%\�}h~.'0<>]���M����TO��+";���cYK�z%�W���k�7t��u��/�y��@�R`��D=A%��qoĪ3f�$�b:>�'b8�#)��(\;*N�L�f]g#-�3B7����tjU�KC��֟�e����6N��d8r� ((mk��Q��w��=����ף�n����Є;��*��ت��q��p�}�˹�e�f�5 ��&��Pd�J����x��U��#A�Z��D }s��2.�ɷ䆜��WW��0�Ͼ��o���<w'�U]T�D�ah&9�@�A���$��%Eg�]�P�M��Rk:�>�t��Ԗ_S����mF�; 8�h	ʷ%y ��4�t��t�!8��	i�+P�ʿ���<cv��`�3~N	����i�6ALT�nI���q4(U�������[Sw��xN�ػd��3" �^g�/�E�.T]4<�΢�*Yf�O�����"�NQ�����[�-��K�t�S����Cr�����w�`BP,ͽyb��\?[��}��jys�\|���0�v�ɗ�i��vAVa��D$ʝ�^�dܮ�7�7��T4@�P�����Z���{
ш�/����y3�8��00v���wYGd��cN�~؆��0����M��'-�I�^�D�Ϩ��tA����.�J�џ�_R�0MѸ��3f�<����X�� ����WB��KrƮޗ�	��(w��%|���KZ��
��
��8�t����uкp,��M�jIUPX�u�O�1分���ٜJn���A�N)M���)�S�x f��D�&u;�h:�hY֊ =J��E��<�R�_�h�r���tN7|?�z/c�`bKx����%�k������1���v��� M�a�~1����8b*/7�\�[�����p�j�Q��1i�S�%-������Wk��n�`��t�] r���TiM�t�h]#�+ضUzm��"�2��'w̶B2�Q���k�Q�A&��N���̐��~��_�q=��}�.�aI�]�$7z"��<T���Ej��H�\/�w芏F��{�]�?XPl�2���S�ڬ�(0���O����Q��\�hD���ޏ�9`E ��f�G���nu{@�����#Ʊ����Y�(w�;���^Î������`n���� ]���s#�zXU+�by��!*��ɘ
C�:N��OfU�����rD���^}qQ8R��$�,u�d��������m��ɩ�ҿ��U,��j���A���x<G-��zc�����w-���~cq����	��s�wI@�D*��<���{�5�w<��7� ��?�V��YG\�}���m��́T�k/�N�D�+6��]�mOq��I$9l6A .~�5{��1
8{6Mc�#�t�;(���x�@I�k��m ����ԧ�*^�B�u�{0; K��/1�kZ۝��y]��2���K��U$�.��(e�Ԥ'r��=���a�� ����3��޴�7+��[�l2���K-�޽���:V20�hA-�0�H�CɆr8Z���b�"��W��õ�ɔy���\<3!4���[N=�ua��s\��-�(ѝ��;y��86G��K&a��6?�����gn����o��������T��Y�-;����\6)�y���xTF �Q$~����웑@o�'e�Wq-|ܺF),���0γ���:��
�k0�4�Gao`��X2��ŝX�2�MbL'���[����2`�h��>Љ����2M���cifEN���?N�G�����^�(��2+�,�R�i���2�m33�K��Bѥ�cQ6t/�n���tH�r�`�0��������/��*���:gP{�+��@Cm �B��[�iY-Ee'$#���T<�7��8J�8��x,��dF���QD��.F=Y�׍��w�R�%3&2�}��/��^�����n���?�M�Y�f���z��r�h �{�:z�%5�U�y<'5���T\��/�UO�O�#D��ȋ:޻%�9���a:#���
J� U�n��׮g[0x_�x�Z���w#C��ʑ�껹|dS@IS�&�@�����@{���e��S!7���{Mf�����l�2�=�1{�-G폎V>��v)�on��� �a�mx�"�զ�P�߮˰�q�w{|�ϱãG�lhc�yǦ2Z��s�J�'u�i#0/`�����}W�؝�Uu�pO���3|R#�~���ꕲ�8����w$O�CRJ؉l����@���ؽ`��6��b�a�qzS�_�����-9sM�}�	c�K =鍇�v����O|7��l&�5~�,�q�x@U?P�p x�r��5}a57����d 2G'SR0d�j��1뺶$Z�,��B��=����zq��mҨ����{͓u�x�>wcԑ�([X������,���6�1�(y���f|:��g��G�{\-B���3�V��斝>�j�`|���%4(7�-�eA@�)�͝p�&��(Ee��BU�Z $5n(��N�l�Y����H9r9~5H9��wMp��q�o�Q#G�gz'��� �/�ur/>�l�+?��	�����U���a�(h�pb�<&!��^#!_�/��B��G�麨�ԫ$�+S8ջʋzz
�rf�=a�9R<���}�E �� 2�1i��h������:����������se[ɒZ���۷�Gw��q�i���Seڲ��X��:���S��QY7*�vZ+{N�5
��aJc�h���Qލٖ��U��8s��F����4]����8�乕k���c��)?1U�˿��m!����C��48�%/xª��ĒF����Kٿ	�?a�e�tӚ3$vɯ�����mLgV�(�W� ����P�5�7�W�<	��T�S�K�m�#�"��`� V��\�П�V���j19�e%��qO�5���$����f�f@�u$�s��X8;�K:�u���G�p6RA_Ƕ�1�"��5��?w��FݫV�S��^cʅ� "�-�"(y�u�J�ސ���8�|�)�vtv���I�L�c�1�9|��Y��e��D��a�p��y����>^M4�|;OC�v`ݛ�o��WJec�M�F��C�Vn�{K�HTwP�Z%Ik�8�P0�ޗEKX�0)*���T�o�[���F��J������WKzQ-tlJXc���*�}g�洵�sp�3���5�K����u��A8"RJ7��`��}�&�~�[�!�zB\�%�6�\�&ʙ����q��s]�C�^�%�V6�����pZ�-����K_XjL���ueQ#�y�9S�c�MZ���\��n��z1�g��
,���d��x�k��$[n��<1$�z�B��̾��#�&�5�)�JY=�g�	&�+l��]���~U��C���n*%����B{���Lƥuvs�P�E���A��)m�pʁ�'�=Z�(K E����=A̲-�B`����~d(��ZI�K~������)��xXk�X�2��eI֩Zs���lo��tPc)9�}�.�qa��g~�r��gwZ鉿0M�\�7I�ݚ3��������=
��b�����{��3\�lo���9������b��zs&����<%.i����K���[�Z�Oekx��x��f��Y��q��΋^\\W����0�ćtc(�����t�8�R�(�c��ӑ/��dΰ��F�Mf.�&�'a�̅b�m�����U0+|mw�`qt��{��؎���D���k�b>�[Vt�N�x���CN-'�b7�0Rn��ڞ���P���j:���@D��nq*V�ט���@�_Y*�Xal�6�`[L�[��\u�V蜺A9�����)	ez̕xL�)e���fv�|.��j�9��6$FkD���Z8��T7pJ|���#�$�F�ܠB hl�8����C7�֌>����A���?��7��������a�� 0�����U��L;kpJ_?Y����Y�4��8����+��F�L�|N�r&D@}��Ŵ�vwЫ
F��d����QM?��F��	��Q���s��bH�Hn���TO��%���"\��K�&Gd��3 �R��z8BU�%�V��ĕ�%�+)[�(G��h�V:qG�Eo��!yQ�K�Bx.:��*BAo�|�Nl�D��<��c��>̩��/3��>�}�(���]h��������ۨo����	�	�Ur��( �,/�$޷ �$��*b���LJܲ����� R�-��JA<sL����%s�������n� �v�z���_�����i</ �������E�Pr��C��¨ˣ�k��� A�0�W>|��g<:,R���N�s�
�|A�АE��m��`�*�ʪ3�k�l�n)|�Hۛˎ�mj7RU�{J��ͥq���m
 �[0fb�l��B�#Ȋ{��ۏ47�������ь���	p�e�#ܚ広�JH>�u����#u0<n���DJ�AH+��`";�6�����C�_���;�S	V� j�),������X�LkY�%��9\�R�z����0�JV�&��������^�eeZ��%?ڃ)/��h��*�W�������gFD:E���q�܏7FU}�' v%�`�2��ֳ'��B��̏@я�����(�����0�0�[nU=@k`hNq�5���O���ѿ�&��G�>�Z� 6����gZ�%�М6�O��U��<DեX�;G�~
*7�j{c��P���d�`3�F�3B5���_����_$ǚ��#�w�:s�����A~*~��Q�h+/<������
�3ST�>�N4��N�Y8V�,�
�0�t+	Z���_�]��P	����ӟ�,�R��{�S|���̙#zRe�����xo�>����m6���9�y���_�2�3<��tiR+�^	S��� H9�"MP���u>����چL�z��*M�����F���ȁu���'ڢ�����tk�^��@����E���me�4SMX��fHD�
7N���m2�ɻ��/6��:�SyZ������t�b�}E���-�;��-�3x��1�@Ȱm�w���V[�Ѯ���[&��o[Xgv5�M�|�_X��)���˰�~~s�ؗ{u�KT�=�++e@�C4�b��&�� jO#T�Fő�C'���Ȅ�M�^���U7?�<c81���� u&&ß�h��x^�ݎ$���g���W
 �g͵*6�X�*�4�.RM>����s
�YO}#����xE�r��﮻�!�$CF�:|�TN�$~G �.@���`����GA�.@_�+Ɉ1(�U� ��}�����٘��u8>�W6������&�E�S���J=J9?x���X\�+]�NL�x�7|�b�3��/ś��[7GeS���ѱ37^�צ�fA^�L�$R}	�49��Ks��V���uw�$g��a�k�0w#<�{���Eq]�1!��s�.��	$E�NW(�j�D��e΅�.*��㾂�}�)A�vq�d�f,;/����=� �n��
����F�� a3<�C��*h�3�N0���'�����4P�<܍��h)�8
�����>�g�[]��?�ɩh��pue��6��Eu#��յ����:^W0N��2���Fo��-����Dn�ئ�S�]�y��.����]��*�L�<�Iߗ��YI�,a���LĲ3N�$<�u��3��w��ޥ����4\x��7.�>�ZM�-��[=�ʥ�|�(�o���o2P��1��n��Kн���Y7JI��AS�I_����-��?��i��SZ-i�����|NL�k��=|�(����An&����`^���
hM�S8h�Z��j�A)����*6&�N)��\n��L\G@�a�g�	pͲ��88������|y<T0�k�bzO�A�UYƤ���,�[�2�"�"�9#~g�7�K�M�!����G�KN��<��V;�o���18Bsՙ�esJ�n�R�-7�:�����R���TM�nE�vu����;�Ǐ�W����g�&hr~��_�l3�͑5+��!O��h�HzMww�*��kD�b��WA;�g��j~��G)�-���v�&�<�c�EM�z�.��u�pa�����5U�/���po�<h���G���v�=�6r(HHz�`�x�r�Xz������J
خ��#�D+ޅ�dZL��iPi�����Vı�zR:�i�8=K6���e=�5�=H��<_ZLx�̔t�f�xD���izOuk�I�5 ��{;��w7��� &��/X�KK�Q�9�0���W���r>H�� K^��p��
l�?���ĕD��4�V�?3B��E�Њ��믐"���;U�Rp�(�Y�9����`2�53f:�,U�>�����F���9 ��5(��o�T�]�d��N~�aJtkZ}���հ������K�w��k8wڤ�d�� ��A8ǖ�z2_�F�B��? ��,��a�z�P�[�u�Þ
���E�i,h�c|��N�@�Y��dL~cC��n��:�3r^f����V���ND���Y�H��H܁�5dѮ��]eSHq*p5{Cq'�Q4�ě[]v�ӧ�{��$W?RS���� <��C�[e��vt����eG#���X��;�A����'�32�k�6�XЇ��e6��&������7��͞<��	)^���e�!z֊W�����\��L�U՞�a�#��#y����S��7e���j�������ʱi>��|�� �T	N��kc�(h���I��h�h\襘BQ�z4��b4ե�9'��ߪ��v$ &>��¹�Fp����?�	w�:��:K�px�Ba!�(��	 �K(��`�`�5�?G@@���!�|���Q���W�q�I�4%���E�xw�Cv��s�
>?/X �K��2���\�[��(�lj�`�'�u>ˏ��P=䇂F�x����S��,tYµX��z��q!j�����n(��
2�e�ƜU��MjD��A���YI燊i��-/� ������`��q�wO�[	(٣��@��D#f�=�"�\���$��'&q�k8�[�X�"F�e����8.G���	�U!6Vq)5p7��̊�����B�8�`��_#l������ͼ�,iݜ��~&�(�����]X�f?����OYtC ��0��!Yb���&��=P@�=J���tmF���0�1x�V7̬�c��0��0�Vk,�~�����I(�3c;s+�\3��L���^E�J��XT�^R<�v;����&��:�lh����1�g}�%>��@�R*Gp��"��,5�4��dyh3u�ΣOkŚ�{�2b�_���I���H/�[�f�x�Q���{��X4��i�y�>�S^Ab�S�U�^�*������1�k������r��H����g�H.�lf��?�����:����RGr*��V`�u�aP�G���qJ�٬:p��^%�hK
̻�(V+`�8����L��ۣ�&#��X����3s�`�"h�^�y�������A�]2����;�d�	����)������5�}W�Ic�l�=щ+;ҦkU�W����sjjƸ�eqa�$чU�K�U�Y�"�d
)���U6(��!�rM%򞖿��yz"�������c͹A���r�= *�o�#�r�B?[>�W#�)�)��,H�D�Io�Kɽ0e�N��k�`x����;��5�%)CP�b����-3�o-Q+�)�[6~�P:�r�"��1�v����J���N��Х�����ʒ������E&���TE��~�����" A�J�o4H��$��B�d�m�"�E�+,*��Tֺi��q�� ���w�p���F�V�Q1�����x�\��t��=k͟) uէ��\wj���[s �&����"�=�m��v�C}�o��Б�/j�}כ�ڥ��g�O�R����v����C�*������H���lm�M�9�e�M���O�'<��޳UE��>�qJY�bh�_j��pX���ؔ�ǰ��lM	>+)k��� +}�C#��c<2��ϔ�C�s�h���c�L�.]27��%��z��l�ar��_N����o�0|��vEpl�p��,#=:+qO��:�
���-�Z:s_�g+٘�����,#vq�di���ؙ(��xl�WK�tp_��Ѐ�!�@.\<��l������	�pU�+��W�TB��E^x7�=�JS-���U�Z �1S�c�ױ�@^:������
m��K�Ή����}�s�r����@D�ʟ��/���1��c\����]租׃{Gv�:�*��m{5�w�S	}e���.y�w��hb�%�Q��.Q���E��>�;�?h���X(�rz2��PL�����N`$$����-$�^��0�P���ws����^л��v��Nl��+��M)���N���������k�h�/�f�:�c��҂5o��=�4�2�	�ƙT5J�e�V5�v�&��q{~���:Di�2w�ir�����~�JЯg������7�M�;��L1U�=TLY�΅���b��Y��*�� �(��J0�1�Wzp��"9 �|]���F�Uėd��A�BDՙG����\N��%��(Z$@Mo�j�#v����\��|\�o�[����$��$�������4��Q�Ϸ��*y����� �[�A�3\qB���� f"�5v�p��3��<S(�]��~KE�V�T��O���Q�f���B=�����AϮ�sDʷs�Q��+�h���0�U�_�ϭ�B�$_�E�bS@����@ĺ�P�r���B�6�ev?�˯l�-�n���ۋ�.����a�묵CV�]i�(���*=�����W��!��tnR�&+¡���:�ۄM�#Ǟ�sՅ}�Be��O�ijɊ�F^2[�_��R�틪�<�P��u�R�0�3��pZ�N����T��rS�(��_��L�nw>�qe�l�C[�P;1]�Ñ������rvѢ� <��Ӏ�ȉsv�\m��� ����w�ʂ�+��Q
<=�y�r|��R�μ o:��'�o��B�Dk�S<u#Z��0���H{)�W�X�ܣ�1L��[<�"�}m�����M�`>���)��euۑ|ޚ���7�m���Kw��9S	�N�0�E{l��2|���]1^2'�[��`��<�q�����t��ϕ��`��΢)����E���������aĸP�%+�L��|B܀I��t'����-���Df�EF�-�wcWg�p��b�P�>K�8�t+�-�dڅ��#J�>�U32u���Jƍ������u���2p������;���m9Vx��\3c��E�l%��z�E��d^�oB���.�ˢŋ��3�	�ĩ�R���a}�]��;�>,	��V��ݩ���z�v��j�3I����b4i*hu�wp���*:�kN�����-#�a̙�Y=��0�9�+ƍ��K�^�LE�q�}��鎯��Gzz��Z�L����$�!�[��� '�A��#�e���}�LCd�jH�W���������Se���< ����ܸ��o�xk�l��D|e�|C[hl�N���4(F�T����xd�'7S^չ��bĭ�/ܳ|r]��\��;����N{���`a�2#M��YN�
�MZC��J�ā�BiM9g%i�^[5��,�g���@�b�v�D:��$�57K]M�yh+#�VA�Թ�K%i�T�>W�~o��I��2�p�	'�ʶ�D�q
0(��u�7�k=�%�Հ%�s�nkdX�X�x��
9�]�����6��7+['�Tq ��R�����Ҍ�r�Ktt�jۭ0�t��5�fM|�N�c�͋��8�S�:Hs��N	gT��Bf����u�����R�kZ�~H���\_��#�!`�U[�w}6��L4����>0F$t�)�YI��%�����uS����[�N�u#(G 2�L�/A�M.��!v�@k�	�"u��d���p׏�yw�!I��շ��N��ɶ�Z��۔�u��m>6���F恨m*�!�4$)��c�8-:����Ey@��wm8�4��*GO��$�H���2��Sx�vz�w�=M�:\L|�0C3Նf�:����,
��ך,�V�Mv:n��V��n�yfl��wE����>RV��9Y�4(Y���h�b紗���&Kՙ�w��0 kj9����C�l_Jv�E�9&3�hIfi-EYH�����_<n�hR�-p$��?�u3!�	��0��U��-~�57F���0�Ǡ�c�ת����}��&�����b���BHo��o7Bq(�^m����qf��Bp(�T2�t,�q�7奺}���~�g1n�4oY֪k��kH1�^���*���є�/��@���FnX<��?��1��������4/�d�a��ow�ȕ���~=��O�u��o�OĶ7pњ�)FU�������M�U�U�2(L�L8�����C(���a�kf�v����r�&�1IR}w(9�� !��s%��r?���is~Q��-��}T�NL#>���Ӷz�}�͠봯-�����F�۱` �gHr4]�%+c��GXt�*��#�j��X�,���ݰoN�< :�ѣ�H(#;�}����9c��F�4�V�m�(GZ�ѓ��>&m�c��7�l���=�bFr���t�f.C?k0��_�x����)��϶�y8�L�V{��-������+i���+w���K�wϵ:PK�/�m�'�?�4�މ�w1<��d=�D�E�}�0~Yr�Ш),�z�CrbH|�]G�<�iM��	��n_���u��5���v�-��%�؉m�bq�4Z�!|?�#���غ��lp}���yx&!P%�"d�Ӊݯj̀�
4ݕ���i�������i�F`�^�0�xM���qʈW&�� ܀����T�0����_Ss����{�wi�όN+�����`��O2m�y�u�9 �s�cU�� ����V�<�҈x��2@a�F�1������:�k����_+ز�dB���ɀ|�U0Fwi�Si���F+�0ǈ	�!�'&4�wX�Y朂
:ɚ�vC���~����S���J�n	�Z*�i=��g�d�j�I�@��Ph_�h�v�\�I�{��s���`k�-B���#�J_��������I�|6ゕl֋���tuj���Ȅ���q��x�����gP�z�"��F:C�}�[h��}�����5뵄-1e I$&�|��I��q�k�?��Q��D��=��]̢/q��;�O�W��_zY.���/�l2B�����!_gS�.N��Tx<j�韨^���[�\���F	gpF�m�Κ^�F�ɣ0��d�f!�w�S�m9e�º;�D��y7����=��|�9mV0�mJ��"�?%��ҐA�9 �42Y�����Y-¼���s���ZM�xr���AD�D�%E�P�Z^���AHTX�H���t���T2)N&k�
<xdR�¡M,���n���ݘ�8P�05�D��Q����2�'�B[���=@���τ�#�-3���Q\.\ 
���L;I�L
�Aj̘�%�9�:3''^�$�Tl��_�	��tY�a�>x���;\��)��c�T �:ϡ|A���i�$�)�A�*S K*dR�M�[�h�-��<FyL�t��ˣ�ku+�?c��Lex�x���K��q��R<�(�� ���������"�w���{-�ITC.���u�AЃ]i���@E��@��j]Tϲ�(s��s)Fy�D������z�N��0�Wl��@�	�&:-�A)���,!6�D)cח&�ـ:]%�H�3P⧯����T;�ʶ,4æ(�x1SC�V�0���� ��4(`B!�R�Ub���P�B��4l�o�T���7E�AIu26�0� �ኘ��t�Ӡ�����
�f��s'�^PIg=���a��ƽ��/��?\�Χp&;A!���+�e�v�J6d�[�HT��bo�(X��h�'��NÄaeh�����:3�07���T���b.�A!�e����l%Lp�Q_�FM�[�y	�������̤�>���]AX4�J�53��i�=-TΞ?��oKS�b25q$�mԁ����&!�����eM�k;tӭ�s�Q¸�V$��0���^�w�i&iΘ)�Tt��8��e��i�x�"��+��4��3�@�Y¼G^����GQ����P��5���|�w�ßm��=a�/D>���7{+*A
RM�dյ⛯r��_4�{S�	m8��ð^�M����)���<Ψ Ʒ����n��`�b}T�8�����&�V�.�<2Z:���@��v'�0�$�͚�=�Ʈ��H�LW<�m8�P��'��B�!!gSK�AME3�*���s)'���q~qgb~j5����&GK�`Lu����?�=���$$/�&��0��:���˙WR�Sy��g���xj|�P/����?vL�c�h!�^5���(����T錗�g�GS�_q^���|�����N�C�ˢ�̨��� g��8���oh�n4�$m*�7�%��� a��Jb��y�,�Q��
b�E��ʲ��湃[��ƅH��Rނ0��$�.���8��g�[X��ȋ���E �:���wƶ�͑[]P&��d9��o�g�J�\�����?��\/1��=�\����	����+7�K�b���d�m'�*��a��R��PB�8yrq3U�GH�P���,4f�J��3��B��R���ާԥ�᝚܈+keA���x�\�v�n�$�\\�W�{'��|V8�|�L�v�M��_�L�Y����n�hʷؙ����1�e�J�kP�m8�R���j,
�T�y�&��>�ե��&3?{Hn��-�8������^������$-�r��)�Z`L��
��P,Ɨ<��VNj2�}�i7�������v��g�SL;�
tk#����.���94��S��U;.-$�������ԂV��q�*@[�n/�T���&e�Px��tT~Yv��'<��HW�D��q�ܬdK���5��b����^Z5v�e/�����nM��!��/ё3�4p4��g��Wj�H?.Q�P`���<�s�rnmK0�̠뛹��g��P;؊w2^(B�,� �A�Q\D5r���\wZƐM%����S�q*��c ���!���۠(�Q���Ei����M�s��cL�5�1b�%A�'1hI\����i��(Ҿ�|���I��7F�6vO����*�9AVR���+U�����0����e;�M��
�^#���%B��c9<�2��!�`ak����
ǳ����1l��Г��/n�\1Y"���)_�B��nX�\>��͙5*-��]��ϥ�����-���op�15���b�G�$���zvU��܏mͧh���{Z�F�`�j����7$�j�TG@��@Ƀ�e^n�z��1V��sTw�����MtS�d���ui��������v v����`�Y}U ���al�*@����sUB9�>X;=۲f��!�&����]#z�ȧ{q2�D�S=ݝ	W���L�r2�T�_/�}R]I�L��C�Α�͔��n`)�R�I7�F8�;sj��RP>�a3&�O��=�_<�j5A��:����0��9�w����of���1PՆ=<D���a %[j{��-�p��~�5
I��Ƙ����$�D��H�'�����@�U,F�lD���o�O*>��� A�b|-��;9�vh`跒��]�/�T:��l����1�.����]��0X���1}P1�R��([_��@��ݟ ��th�����B��vī0���pw~�\���8�v�t9��e��5r����j�@4�@�.�-[��NG�@���E�Vi�v�P"��ԥ�������Ԫ��~/��e
�R����G����>ۤm�h?e�@|:D.��\�:W�֏za�p������m��P���)n"_
E+��5bb�r��b&Ls�I��PE�W O{%�"�$X^c`��F�ޡ��/�6���[�gQ���ƿ�篌�B�k�����#����+�<����-�	����l��\I����'2_����=�1e������{��|��18;~L_�0�ƇS�s���_��gˡ��X$�m�؎Z���/��= ��hc�)��s�-�FZU�MK��h�y��{�o�J�����V���U<5�/��,8�I[I�찱�"�K�|fsq��hG9ǜ �E�`e�� f.����K���	�iU-���6Tu>�h<-"�"d�`�,]��΂��} Q�����;�#���i��N�	�)Ϗ�Q�`2���.�j��N(�;��B��̂ nP��*5B�>�Ʃ#y�A���[���~�+��b��,����a�����-�H��A���H�@�!�.�#� xWfX
&f�Iƥ�#�Y�Ĺ4����^����`����4�〷�2��bR}$�b˸l��c�dS%w��ch�r�z$������� ��)q���#���)�49#� ���Gs^�k��$��g�{��0qG��"ទ̀VleO=8�½BH��U����&��Qxs1ߋ5%�}�0����xs�IW�=�r�qL��b�@L�y��&��0��aL���Ё�s���_K(���;��xv���w�1�YaѐY@�KN�%Jd�Y��/Ӵ~�3`l�V�/1��(=�&����{��� �n$��w�mJ�1�f,\�;�S�C��#��̯\�=ցn���{��H����Y�@��A+��c@8QV���,�������x(�!����Ͻ��7I��-޳��T鞓��ⰰζ�*��SD�-=��E�N\�F���l�Ƽ���d9��u���BۑC�NO�a�����9����Ժ(�Q7~^z7�����nM�]�r�I��5��Ng�dkC�V�J�8GQ�2�Ɔ�j��ѧ��(#-�
����*q��eP�WعA���ؚ��)׶ /H2�)�����=�57B �m���v8��A���N� �N;=� �N~Qէ�U!�4�����${U7G` �;����ϲ?纻�8ި�}f�����z�/\_պ+rq�:ӳ&]�G��DL�6jg�V����iPo���i���5�2��� j�'K���-�W�6�-fWSw��p�P�a�AjC;��Ff>v煡�A�$��~3�����_�z-���5&YG�� �kV��S�8���F�{N-��Q[�{j���� i�k6���r��K���7�� �z����޳X�.ho4���5b`�X�ï��ԕ�����EF̎K��2�D�}<�rU���F=I�pt���CC�\ck|x��=^Vu��%h�OD	{��Z���|�2}Is��W�5�]����w'A%�V=P_�
H��vg��D.B��9_CIa|��P`�-���LR�Q�y���yi�4,+,/H�e[�	�zi�S��xa���,ݵħ�"���Oy�Tm=D���w�Ϥ��Z@\�mB�[Ɲ�OS���"��C�T��/ϓ}8�^|>m,��4��(/�qb�E�y��R뗣��*dj����g~֫Q��`cq�.�s#��D*�1�<�tzM���s< g�yqL�3.�������8m�~75���Ars^���m�����x�%��EEݧ�_��=yx��+��\����M��ti����X�a������,��~ C7�V��D���S��٩(�u�`�.�A�e���'
�kL8ylgwo������p��j���{�](�9�]6t��"^�	����I�|���z�"h���~AH�:�/�M�?�b�u���Q��wtR�V�{�	�Bc�A��$����s���@]�p|F�0�#�-0�<�v�SPV��s�x��ܩ�x�F{0�|�Fv�����J8ˠ����6�ݮ +7�������c24����4�BDw���MC�_:t���^��Ԯ�&�4]9���h4U=L�t��P? �U���J�2wꇫ�Rr%�|ۄ�~b�AcOABjK+�����������f�Wt��_DD��;���u`O�ˢ.JNHy{����Q�M��X>���4�綝�sR���
��>A��Z�����?!�����QП�Hⅹ{J�9�C�\�p1Y�k�]�!^z�R}8I��{���dW0{?q���g{��j�2����s���X��`�$}�oc�i����.�hF]�JU�������x*T5s_j+���mœ�8Co9�-��4*�2+�{�>M�fM��j�쿠	�Z'k]��%���S���
�u:x�;(F��%�!Ӗ��F�+�{Ѝ<����	X,�-���2 Ck���A�,I;��W8;Iѡ	ޏH�G�P��*���gx�Mf8&�҇�Anb��H� �Fgw��/n�if���gsT��mE��/�I[���'?��b�_��>J��:�j3@|�T����i' ���L�a���s}Ԍ~a�$�5CLOͻ^u� �����وӭ�̬8W���~h�5�f�j�,V�ar���@�d�
v���8����R��Mb�s��2Z���*��~Ͷ3&lq�M%.��7(��9A��~�`�^K%�@�w��ۤ},�y�G���l�*_��� ��`	��O�_p �J�n���nt�vgW���%z�F-v=F�w��/w�����c��� �P?����f�>��.�� ��S��5�;�4���c,bp�ɻ�ԓ�����#4['����c]m�zJ� �3'��s�%����=���wf������'��(�k����zd=�=���	ȍ�kY����Uؤ��3�Y����Sy?��i?3�?�]����c��{i��jr��	t&�a��Q��	�^$�\�h�^����f��$������$s�3�(�!�)��e�7W��1W�H8��Iav)?�͔��L��=S�J��XfQ>ϐ��#=�ʦ�5�/���t��l�D�. �u�d잮q��#b�S-�%%�����Iq��rF��I�m
�*�����(2~�e����]Jd�K��`�)�7J޻/�2���1r+k�9����Ƭ���d{�p���a_*�\��v��W)c���b}x��ixr�����.�8��+����HP��>7���� >��?:i���g����H�A3�F��
L�����>�h�ɕ5��������&b��@�K1�.����vFT�6��d�Q���t�@���uu,}T���4���^�Ηi�kQ�o
���o����ݪ�2�ܵ�����o+��