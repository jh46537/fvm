��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�z吴�)b���ΡrϷ���	�J�|56=�#�#�Pf꾍�F���Z���j�eG<�hЪ�r/w�O�M4Q�B�dB)��ʁ)�����ҨP���#|O[5��'{d뎪��l��C"3��~��R�p�"܈�������ag��?_a��fX���d��smۓU}���>�O�iwƛ�=��ˑ��d�i��F	FO��{�i�����UB�O�I�]j����x�%��1���lC���?�Y�����Z�[���륙��RQ�x���1~lі�F�T�<��7��ض�K(��B�PN�C��)e���d�bU4@_뜽�����f�QR�R��b�:��G�34���A�q7�}�A"�/�@���p��`�`��p�p�FaH��<Z2?C�{,ɗ\R�ڻSZ
�>��j�q��Y����m�k�*a?�Pl_����%�ۢ�SJjhĪguO��/d�&?�7ү�o�u�N��Vp=�&�(U˴n _z�yU�>���!�Ch�
ywA�ꬠ�.��W�%�913�:"h_���Z����5�'S"�>%o�B����=��	��F��<��됰'�8�"h�D^F�ꦱ��o�,*0WIx�:��|�O�ŕnD~GV��ZY���~���F��4���Yc\�`��X#�th���v��3���H�Ce�h���x@�I+Qoa�KEE��t7���i�;,����t�p�3 �[�~�����`Uf.�r�Λśz�m4t�l���[n��f{�X(?E9X��՜fk�����C�~eQ��lF�>~�������@�Qd���Y4pK����視��\�Q�t�(�{x��ZB�U0��{��1�����-G>9��������[��Y��&J.�V&9���ɼA���dV�v/kY�l��ֵ�P��q&
����\��?��H��g�M��F�NL�<
����ֲ�鹻��.������>z\�r�z�~���$/׷������hO��(e�U*����X��\���(���]���Lu���[��֓��F�"�(n7Ç+C]O�_��	�31̈́j�G���K�s�O��Tk��z/٭������[w�U�5X�z���K�-�I}Kj/�����h#`��g��sz�=������*l�$��]>�Pq�\�dK���U�8E���Y[mdS6sO��L2��{�q�$ǚo�"M��n�wy�h=ʸ[�ǥ��O08,z"�EK"J���΅��ξ07,U'u�P����cΩ������41?���C���|�P�������*��c����1��@��� j����yj��l0��&\�@l��ǟ�vel�ޱ���J����.�F�_QZ\A��jJ�i� 7kp�y�S��MJ_�{�)k_���$��f�xN�T (9!`ٌ��eo�A�S��%^�#�L�&-N��Y�{<��7dz���@��L�$5"�&K̘�{���6��^���7+$np�PU��Z��{e�{H���d6'q�;��,�h�o�f�d��h�+Z�tF�v�b�層�z�N�o��O|zٹI��X'�l�]C��"�:r��,!o��v�h��:��3n��5<���w�瑯��"Y�4��tj�޸O0���9�A�Ҩ�I;���s]_��8᢬��u�/�%�aw�n\
����z�G|�N�g���g)vMi�f=�xBv��hC�A���a��b��C���>��>I��z�$쉇(��J�ʬ����쮋����t�Pa�x���?N^W�����p�-��� m�Ve7����z��a�A���<��4�SG��a"��C�C��{�ug{h��1!=	��q��y���{�Vj�^1ِʼ��Ic��'O�ocU�7&�;(�/}7�}l����G\v�,��1-�%^,�YZf�U+�_e���\���ɨ�}����=���',h��5w����-��x�vkv=G� ci?oiK�q4�[�K��U��I���m����㙏l�C�O��Ǫ2��� [wF&�Uv���LAI�p�����~@�a;����k�:�2��C�3NO(]� �?1�Ձ
��"�1�}��f����0�HW�[�}�A{(���`�6G��%�<��\�s��3��鲀�������惚Ln�\2�r_O��̎�o��̼&�ԑ� 8�G�`�#�KY�_��|�R�U�
%�f�r"�q8�1	�q!{@l�NP����$��j��1����A��-��.C�������&�zi����K�� FM�O�(4�y�`Qc� }� �d��ϛ��O�:�W&pw�6�����pE���r���GX���$�#�U�TbAݽ�&m�5�ӿ�R�n�\c�u*�'�qj�Re�M�¿c9���9:��18T0R��6��K�ї#�ޖ����P��wƶ���1F���q뀮g[����"�U,��ƅc��F��d��"�N���M�<P�:y4���Wxkؖ�Ŋa�d�6�n���A	�A�}�?�[C帅v��Q�O�F/�I	B	��Ut��I�-b'��W�B&��dR�7aJ�S�t�b�6k��Ζ�2��uU"�
ct�2!�p�|S���2G�l�E}���kz�fb�rў9�����e�-��q�[��y�����4_��z���Jh����<����t��࢒�k�	�����JGk������Q50m���t<�M9��Nڡ���*�B�����B�!u:�܅	��V�aӢ�J��s����l�@Nl�������|�n����wAHK9q�2�bj<��o񮈧���L�oXB�V�O�����ׁ!�K&n|��'o�If��2���˞x���go����w��ֻ�7��Q����$->��+�P)§�jY>�#,�doR�~%%�Y�ll6.��*L�7�B�[G�m�ip���
�f�n��'�4��T8a�5f:�kn��)��T�7�EjbS�Ʃ�h�]8�_�h�c���l��tS���o|�9���*V`Q�����Σ�v+6O達b�~�I����^Z��y�� �5 �"����]Ϙ��5����5? �;�@B����}W}:X`��K��	vk���"̸[>"͞)B!���v��zd�5��M���vn�wtU7���ڣ����O�k�N�k5M�������.m��P�U�_� �LHM��I�ʈ�5�����سf�do|#eG%N�b���N�����;�K r·m�����gap�C�0%ku�1�2�0u���m��z����W�M��b]��.��f1v�nEx3n�������>yU�Y�)��'|��O��p���� 9��J�%@ff*ʩ�e�ֿ�<k����l_�Yw�F��h)a}^�Oim��f���F�ѕFP��'P��Z�ӽ{	@�{X�I�(@捎��w��f��L�QV�OId�FW�,lѲ�Iz��-�Ǜg� ۚ!IyH��P��D�=hG	_ ٜ�b�9��۠hB�t�GU��f"P��ԁ�ЕdB��B�f&��`�ql �
�W���UOL�fA�9LM����V���%�j��>�����Wd����E�v���x0��xR!��$/���w�.���LDΒM����d���B�� T��k n���Y�V88�ZZ���W��ZK���`���l�k揸�`x_+�����T�14��*��,5�|@���]��Q� x���
��]E�<[�x!k"U��\���l�G'8��z%H�y�˱%Q|���_�=E�$�;1�ԓw��=���*	��4�0��$m�;����G5����ym�)a���O�aY����8��j���c�Q���07�)��zf��;ݰ.���)�J�8jC49Ʉd�d�~(��D�"�-�_�l�Q��$a��C�q9��Icb��6����6e�[L5�YXjQ��L��0Mr"5�eM� ��RA���Y��4JRB���g�+�`^���;��T�~�eP�ιu�)��詤�!����nH����޵��\�0Hk��a��
�(�6ωK�=��^�% n�0���3�7���懻��7~X}��n��G���r�H��4�Ϫ�/����$��v	�Eъ�{��ȁʲl9_1.��6M��;ˌ�4�����30E|\PF�W|"�8/K�^�[7YyǨ��"�bk#�=7����?�`$KT���a�%��r>�Ɉwz�U��{i|Dy�5�L�B+�WxT��r^%�D→�� �ܘ��Z�=ڮ0� ��T������0�K�p���
z\>��y[��FQ�˚k�{N�5	'�J��;L�9��[nW}R��l�x��5��)���~��\d�_�MY��4��C_���ێ�-��}��d6t�C�/{��(a��eH���qP��d�R�`E �So
�V�2eMM��K�)˕%�i�'���S8!c"�?��X�76Nf-΅��vhs3/����f�4���$q��s���}�r�/&�+��Ҝ7l5���y������b7mW%&Ew�2�a�eq�w��T�@$QF�cpf%G�7��9�[LJı"������ ���/���Km�`3�:j�����Z���~��$˿�-�w�1��ӗ����uΠ�lT���� u�k>c��p�y��=���Ɛ��v¼`6<�K2�	��y���xyi�5J����:5��Jӱ�9�=kw�K d@'�ۗ��ET̷�v��S_񢱚#״�H+"��C���L�6�  )Xa���%luy�*[��
�
���#����
(#⋁.Q;��r����d,	�N����pw���;����沃z�(�J��{� �-5���w{`3�Ҽf5�����3��ĝ݃��R|Ƭ|�jcY��K "e�Cw�DKQ�����+��)����J���m	靸�q�c�؇!-��Y*�mW�������a��H'�$C�2����	�(>�h�%�a�
%��,�R'9L�OLu�����2����)�4&N�p��EGeʹ3�I[LM�)�X� R��惭h���(�>e_ñvc)���G��xJۑ���|f��sOįFߘ�5,�b�#Px�87����B�!��$M)dh�uɕX�TV�)�1��#���Ad�*e��*��>Ȇd�MC03��UM38K�8��*�%�7��"������"�"x�eF(<Q�Y�CIx8�ppL�=R= ��}EB���|f�5�z��� z�(��.~�}9�O�sǑȑf��$�Qĺ�~nzzZpnp��s���k8�ṕ�_g:uel`�LÚ'�����ʹU�_!�,ء����rFu�S소%L66�!v⩱���1{� ��������d0������� ����	�w�j<,�5-:���7���P~�>M�"����#�瓕��7���T��!^s:͹<9ʑ�5�x���ob�0�$1�l������e�����Oj�p!dE�RY�=�)��9gh�����Y��֍Շ�61Q���<O���ۃA�鸨Z+@�c�;4�Ϋ �wn���S����n�O��rHTd�+�E-�G�Dx�Q��n��?��Z	�Gys(���M'8�c�F��d7�����ĝPA8�&mh쫕�t�y�~9 A�,�g��A�#L��Π�M*�~ #���alaOz�W�3�'�*ƍ�ė��<��^��L�e��果�~��J����?�)+�v�?4�É�QQ�Nb�1g]ag�H�#U��r����٩�)��}�c�!�������tj�7P��Ńu�F��S�>�C��܃�:��S၌(��)a|���T��{�-xI���<�y3J�D���,=�_�`���;e�X��Ur��)�`S��aNY��߱�Rh`��E�瑔t�m�������������Ȼ�V{<ܴ����c�.��v�iK�<��d��J:���,��I�N�L~�H���M&.&���-�:r����Q����������%=г��,���?԰/X�����
(2�M8%�=i��� r)��n��P'&�z� ҁ�c
 ��N0'lpr&�.���+��Q�:��h���wO+<��'�� %:��{��g׃v�x%��%�xU���"/ט4ں�@�x�y���H[�9��VhT�$R�4���9I*փ�͂
��%�+l��,$�V�Y�"�d�6�Q2�g?����n(��Yශ ��Ļ��QݯJt��vm
4ZD%Ir�������i̬Kl&��P���+Q<w��+o�9��[�᭯XO��J��샕 ����fS�n���T�D�v5���.{��<���K/���l#�U-��]����6��46˥g`b�pY(u��Q�˪%C!�[c?��OFAJ�3i)��<!3ԶEƱ��0f4�c���7���<^(Ո�Y�G;�b�m�5.��&��>�"����.	�K��4'�j�\���=[�D��o$Ur��W`���q8#�q�����s�C�yZ��kУ��C%/7>������=FFСʏho��]�;�z��
SfŞp�.�=I\�ቮ�!���n���tE�dD'Y��_N2��nq��'� µ�	'���Z�DbQ]]W���r��� ��GOv������L����m�r�K3�X�A�Nn�8s8>o��j�ۺ�� ��
�k쩂ֳ�h��cׇ��thALK��^�o���&�n�y��;�{����r��)�H�%�}iPx�݋�����J������JS�e[t��y��GI]~+�(wܢ��}�B#�A`&����B��ц]�c�;/���q {<�Y�������vI�Z 3D}lw ��6`q��6�,�&�;�DJ�>�jN�qQa]g#�sZ�6�%�оT���#Umr�gZ'�F���=n�s�%�M�9&m#�>�3�~��7{鏀A^�+�D۫�ٔ�����Prj����!ԣ�Ԧ����)\ w��1�9
a΋���8)ԟ�6�o�r�)��!�ۨ7J��)A{��H�/�Wflspg+�j���W��!؞�N��1=�HZ�� y�0*�֍��Nt���I8f����]�}�<��%󥶡jf� �6�K:k
��-�3.l���G6a�Hˑ���(��_�������'X�f�M�d�$��q3��lj�(�_`��D�A�(І`�2u4���WEjϟ�n��m[89�-�����7'*��أQ��啫�%��o	����_����߶U[���Gx)�<�����E�f2@m�IT5Ǥ���ep:�Wm�еX��:f�$��Z��>�:���v�h��QQ-�E�p���
,f=u6�d%�"���$����y�g#H�&T��&����,��(r�DlNB�}��m�GOro� fp�{9W���	����'7n�'�;�ku�yk����鐽��zs��d��g�����0Xhl�C��P�K��'���	�r��wMJ*@n;^�lu��4)���ut��_�uߺ����5���k�$�xPJ��P���[���?��;���J$8��ˋ���'՛�׼���ٞ,��_0�v���nZ�{������#�*&���7|���}�pF=~.��w�B;�YǷ���4�C$�E�LJ�{��P�ӵԦŇ�Z�20�������a�J�H�COO���Ïn޴�״�s�KK5��V'^�~f��mȅ#䙘��ܽ�
4��A@mhWf��K韷:h������"��fI�3���m1_�J�ߖT_i"l�n�U������Ŕ0vV�ΰ?#�ѦOl}i6_t:�r"���"*I�o�Փ;��� *QR{����Z9д	m2�v��C
�6�pmg����z�����S�=`�2 �M���ZH<�L7�>x]u5QP��B޴��-i/̸��%���J�q������R���5Z��M���A-#I-�s�I8:"�kRB��a��=ϵ�S~@�K��r���9����[R�,�Y!z�P{�[x*=H�/���ӄS�,��?����H�tE$г���n6�0�so�M�i�c��"���k�p��{�� Mv�E�$Q�c,�1P��!�i^�����;8���L�����1e⯯��~�@�릐�z�hRJ�U<��C�Aw�a���鶔Z�t4M)��M��fӧN�a�23�%��W��g�仫�﵊[Kgc]�Z��sRà1�Uq���E�s�zW�R�g�P���`� %������+q�r4��=ɬ�P?b��q��{�D�;��Ψ^��`�Y����u�1��ۤ ;�7r)���R�� �s�Z��<�ɏ_����<]���n�m�"���}�Z%��8Ϙ>\��g�=�L�:t!(����H\���F"��H�dI0&��Y��ے}�_����8KY��"����a��e�U�Zvxkr싡?q�o*�+��HaF���E�����-@=�Ru�`�gW:����x����������%�TX��Pg�`c�N����^��X�Z�ˀ>͟�LÙ�N���>dň�yRu`��S���6fW�U2.�F���GT���̀���Dō>`��o6�B�>�.�U#�s�e�_��{z��n�dZ~������М�6��BIsJ�G)�׵���\Z�0pa�-�����x�9FWE�p�����>�Q�}�'�{��j���]8m��r�gG�.�%�eS�_����V6�[��V�c�|#�����՚�7Ҋ�vI��� �	�tŔ[J'1��'��r@N,ż�		�y嵲W����;�~��;�����	=��!1���妏�c�r���9����'G=�[���� ��O^�ܕ#����4��Bb�0I6.��0�8��$��^�b`�eI��tG�M��-|!a�C�n�	.�d�h�1f�2��j����?L�=M��
�m����<)����Њ|p�H-E���독*���}��9$�V�p��ݜ��E*Rũ(`�o�9%�S�熞�o����J6�������	-}���S7X�5�y�d%�lJ$�i��?��Oc��yaw֨R�4�M��R� ����7�`�Ą�d,��U�ix�B,��464��]�Q(����!�`��C?�����m2:��b(ZAMr4� 5oF��i�����i��VYT�[͝A^-	}�`�<��Y*�o���z�l~Z}R��h����c�]����I�����y0sY���ͨ�@�FP<o��g�_PE��ѓO�����=D�1k{*C��Y$�D1�ވ��m]�b�R���fѠ%�N���<u�F��P�v�ߊA߹#�X��32\���/�\�'������KQ�|<rR�#}�F��`��|c���5�o���쿄���>��
�'�x�RM�G�j0��kcd.=f� ��#�jĒh ��Q������{�lF�C.��Tx� |<���J�+���9V�&�;ި"��q�Xଥv齡���?�򺰉�stI��S�H���`��gc0on:�g�V���qv�p%ܡ˞�Z�tᬄ�г�K(2�����B�+�1��:��AnkK���� ��XM1��n�-�w�Z�Y�۠�F���[˸���N�o�!sΩ�e�P-�L��ڰ>Q<�� q�k��4U`h�2�m�ޓc�^���������?�X�2E|�[8Õ�2�0Ԕ���34�]��9� )ݤ߇P`�#,���#�j[ca��4���^w�X��ـ);�~7��I�3�