��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z��W	x(�}��>�W�h���z�ģ�l�%����F&����=;����|�� k�'b_��P�X�H�[8�bNw��a5N[F���?T(���N!)𣞱.jqg=G RN^�£�@����sE��΋�R,�Ӎq�9�q��փ�'K��	�$@s�&>�U;���Q�Kvb��_�s �GKE�  �+�H���.c��(;��ծΕ6įO�\��-��X!��Q����oQAdt"-FT�G�dA��پ�2#�r`�i��%����Н5�-50+73-�o���V<��x|A�Ѹ�AE�����\�H

��Q��vXn���: �'ʥjP�t�b�j�Ogz��ټ�$��u��?/Ƿ �!�������j�τ�Y�^6!�ل5@�s�H��N���׬ƈ���r����+.�?�΄m�ԟX�<��>pV���]p��L�i	���`{Xy9��|�QK)��*���=J7-�8�9�Y}J�w�F=E�;���X�<}��_OM�_�%Ha@[7���7��g�ޢ*8�l$��b���v��@�k��0K�U�'�f��g��0�6't��c��M-w��ԣ�C�k����t�&Y���D���s�XI<D���7�n�j$�0D)?�.[���	BߗZ;��JO{�>����i��es�COx.�m�V?����оr_�ɞ�\n	r�>x��w4~�Y�J�G*0@�j��貌6� �w��Jخ��qN���,��wI;�b��-i��M�M@.��0�}8��g�M��7dL��^I5���hыu%V?+�]i=Ʒ�W���N����Ȼ�������ڐ�:.�����/BG7���)�]�ML������ژ�%UpS��_~�-���R�Pi��/p��ɞ�R����B�2
��u�k�|���T�됵�//���W�Y=)�k��L<����I<��B	�`9��-��ɓ����E��ю��%t�Gm���餓�Lr��ee+m�w�jbuǕ�$��%�[L�+3��DVL',\ja�\�d*�E���37l�U>�A�<3�5� �]�$`���,!�D�d^D+�?6Q+��(=�hf�K�(r?]�ؠX�R'��ZQb�-�Q����k�����Z�켜7�/�U�Agڑ�az�(��DvoG{3��m4BU���t��F���T������	����
��Zw�z��}�C�n��KWO{��74���>f�[�s��u��}�-f:6�
�����޵�VZ���A�U%}t�Oۃ���|V����l|m��{Pl���:���3��%v�i�Q,���S������� B �;�v�&� WG�	8�w+�g8m��@H�����<��&Z���^3�O���1j�}�z�B�S�ˍ���U&�k8�"�W��8Q�
����h�dF|��	�V���+�8QzS���Nx}���N�X�-6%�d��>^��,��Ax�h��Z�,��sy��}W�}J~H�I�/�į[K����a8J>BJvh���j)��y5k�=��<���,���@��X�*?etyX8�Y�GC[h���ER���]�'H2 }zre/ל�V�q.��#չշ����%6�Ț�����!"X�G0�s�u\X	�]��V
��b�{=�w��A�HUV1ڹ�e��澒�cɰ���#���Y@Z��tꌳ�z�\�咵9C�G�k������+ԉZ=�>�qo~V���c3���W)AE�<k>��X �(,6�����4�iD�,�dxM��@A4���3_ޕ���^�>{�J;�X�� ְ��m�<Ϟ'�(JM@t �,���Ц&�����k�(f��[rv��		����`��+5TyP���z.�J���6����/[{,�T�����KZ��d�d���^���-<��b�R�
��|ĄW~jˁb{@wQ�Pc4���Fz�q��B,��g��ӫe\����`��a��6�R$J�ߒ�YS��7͎�`�9�Ra_Ƚb����b_���D�0=蛴`���HmqL��yxyM�,��	���FM���7�Zpɿs(���C��fu��G��y�t^��bC��]��i�[E¡�����eM��Q�aM���o.`�橤�M����&z'�N/���zܢD?2�v�'�0]�Eq&�n^A��Z�J���CR�!U��u�]GA���-zpV��K�٤$wT<��T�(�ZA1n�~��c�e��r~��/����R�C�'ϭhPB��kb�/*����5S����l�2¹*K��y0ؑ�2�3g�$G �A�Lͼd=|�Ā�A��s�=v���Z�bJ�g�q;��<-�L�������	�h�jFj�A}�^m#�GW����y��v�����\�ȃ�2�.uV��ʞ9�.kJ.��m�f2�������v�T�����ɒ(�M21��Y	�}�oB��4�PIV<,s�o�NC��n��R�3}5O�T,5��ɹօ����H�!E�{Ii��}����-L�Q|��̣z�Mp���6��Z�͕��Ѥ��X���&�+Q"z�s`�(��Vv�xYv��=[ĒX��R��,"�n�_`q1e2Ytȫ��;�T�y%�o��/��/^ڪ���9`H���&��`���T��=7�eX_�	��M��P�]3��٪1s���� d���q����xgĒ��Wt<%B�������B��<��	B%�y�!�����<=_�:i65د�o���Ƴ�$xY�� ������G�E=vuQ0#���W��ԹVL�
Q��:p}��t�8P6�J,�;�*CNA�N�cMUy�n�W#�� "�C}ݍ��
���e[i1�����^R0V�O1I?��c�t��i��x��ޙ���eا���˩�N��}������D�v��Fv�@n�:��fʒ��.�'��ď���]za�~/�}(�ր�z��nhzF��	-�jJ�͘�A�;s���(���YW��s|����{�l/��|u��,��9 ٟ�p@�д�=��no-�O�p릥8�Z��[�z�Ш��T�JG��̀j��D��,�����<���So������@�KMӿ��û=L���-5��R����QsM�����L,����;ؖ�����J���5�����^�=�����@%���%�1�������3e��C��D��Z��G��&��-~�����8��Z�q*��������p�W���1&̿�[�)�'�Q榱� ӹ�2���b��>RZ�q%w�9`����߮ȳ������;�u4~9��_k!�z�%���J���B�D�\�Q�_e��L�4���:��p$�N�T��#��ջ�:�k�+�,֋��Ж��J�EB(v3�^ ��K���Dn�Cđ��E;kVp ׃]������Rl�G\��`��|�f��?�P���xCh�h |[H	ٕ����f{n&Z��(�� 4��\z�S�\|`Ce{kT�C��������J���nѡ6r�09%�2��]O\Xf�ųFjFSJ�d 3��^hr��i`�D�+�-m���CEz�h����i�C_N/>
e�RĠ;���p�������1'����ʀ�Ed�t����D1Q��f�h�Ԧ+�3K$(Lh|����r\�����K
Rv����f�aKb�d�����C��U����(��Ĵ���x@z@x�p�J�U�ԇe2`�-���s��[sr����$���uǙ&��GU¤4>�`+6�n3���_��r��7�[]HU\���W��@�9)�"m�dt�V��k�bx�).oek��IYe����m����Dm�m�C����N��b�%_Բ����]��G�OȔ�$���W�k.��~�9�1&�Ht3���ʐ�Ȑ�U�{�E�z��xw����Բ"~���iFɿX��>Sv�����4<��^�����7VA~Ú
E��;d0�0Y��X������j� ����Ё+O㗦�AҖ e�5�o�����,Q��Cp����9r��%7�R�fr�15���B<"��|�{�ĊTm\�������7���ѧZXpW;x��f�|�3R�-�K�%#��Ċ�Xթ���]����S����3���^n=Z M�g��k������m7A�?	cuP`�7L�'^x������HhI丠m�=@^nt�U�A_��d�G[D
�(��AE}>B��p@�j�t�Tj���4���לG�UU��Jw �xG���Ç�zX��3?ɭ��B�$Ta�ZPF��fs�8&�zY���;"���N��l�E|KB��Ip���Pۓ�|��li�Y�B=�ي��e�E��2>�'��d��mI"v_�\w �B�&[:�xGT��;���1q�Ķ� �M�0�{���(/%0�E�$�>s�\�����BPMG|P�r��.`�U��C�ޭ�����Q>�k�ސ��=XY!t�!����+����'�H�3�ȣǁ��v$�bG�{�	�t8�?>�\�г�=���)�U����Q(�g�ILI*����{,B�	S��u���Y�]�6,M�U�ެ���j�F���R�he>	e�s.C�;#:�����W��]Z�X�*?c)�b����L��<����~a���e�?0y�Z�<��+gж��a��t��(J�d��f�+�y�b$��}��&O"���o �T"��hx���ɘ��qgLt�(�d��u;1k^L�`��0��J���d�$�(�m�W�j��	J�h�l�?�l����0}m	�4���G�H�ٺ�F���\!�RT��D#�`�W+��>9�dƈT���r�Ԏ)r(YWlp]��1��l�v�� ��-���&���X����q<�ڐ��x�\�?C��!dN�K���tz�u	�yF*�{�������l�v�������v<�6��H�F�.��mq+�BE���&����4�|���S�s�(�(A���ӪZE�[��d~�]����k�`us�EsM���٪��j���x����-�,��7���Ew4��G�&���9s�"��{b�"�N̦�l����5woﺱ��&����xV��R���d��	��K�ޘ�}�y��Sq2yYQ�sVBf�O�
'=��ñ^ȕû��;�|����,\�Y�
ԛ;(yxt�F+Cs�id3�vY1����b��9m����j@$��|s��9���&o�:tP��I���������p=~�%O[�o>��shZ����yu�~yu��[���B��b3ߔܨ���l��@Qp�3����s�,�W�V4�lLPh�2��^��p��0
�#�η����Ax_}��;8�0�=��co�NM06���f�3ڸ��)ü�i�ӗϏ��h[en]�����r����ni1�ir	 �W��� OU,V �����a܆�|
���ه�c�z�g�m�!7�v�l���V7�Q�� kZc�{N�����:��\O��v�X
��g-K^rCpI�!*��1���X���l�:���'^sq��V���9r,#�_���*nl��=�����)��y�f`�v�{��aH+>I����;�f�T�<��'�\x3%"ڍ�c�#���	F�%���5�I����V(�Փ�}�_Ht����ןT\W��������X�S���L_�D;����HXXm؎��ɗ�����:���|)�jw�����W�7��l��*�gfo�C¼�\N�%�;���~�+�qDheZ����~rdX�d������_'/������A�?8U}�z��������ז�Vv�\�-?1��\��XX�=��_����`1X�u�&̻"���F��b�����4S�NO�����ǵ�%7������S�jeuMd}�����=�O������Z��1�	U���ʫ���t�+���[�$CJ
�2�k3�a��ѱGf��ԏ��*�
���P��cI����qa�.�z��Շ	�.�r�*C��%�ZL�я��cz��ٵ�1����Mc"���T��re�+�8�['։��Ur k�)���"k����}	��nZ�I�)����)�]������}У�a&E\~�a�B��xw�e�K�d��5����b��N'��l���s��IP�'��
�f�`��m��w��*5@N�]G��d��5v��E��[(I�L|z�t�"�f�J�4�Ǐ�Qi�{��كl9D5 ���F���(��~��e�%d%��
x�IiuOp�6su;\d��s>��5E��쥚+�Ư+�J8j�1R��������y��p}��o9�f܃SQ�[뙒r͙9�5$����tl�q��������
	�򃗏Bz��h��7_�̮�̷�Z��d��N r[K	R�,�*���,�VH_�AQ�X!�?�(��~���J��Syc+J���8u��DDnﲂ ���jÕЧ⪡��\z���t쎶&v��j�Jn�X�,�U�CUh⁣9EIT�t>�פ�� ���2����8{9�Z`b��m3�B�坹��A�F����Ȥ����<z��6iJ5��DAG݌��F�9�6�=.[g?�0�W�E����h�=h�9J+ǟY������(*>�[�R`��pə
���%sֱeI����1�(li�y�ש�n[6�5aP�~W+���W("�޶D^~�*�` %��c;��rK.��+TY�C~����Q�!�������(��[�w���������'H����}vE{mP�*�3�'/p���2!�c�5�ey�;�Rl|���>k1 ^�QW{2��������j��KY�����(�NN��y%,���U���I�r��C=�3V�� 8<����2�m~:�°bX��g��Yx��b�Y���\�p���oQ��uFv�v/�r��3R��\��y�^V4�����5^���X�9l����>�ko�*��yH&��'8���:���Za�̢lS]�4�3^}�͗�:q���7}�������م�����o�\r�Nh� ;Nq�ʍD��r���K�-x�
X��>
f�d;0 ~u%7�ޡ��%`���%�{dJ��ZM{��>i5���&#�c�.�j��A� K=��zĤt'�7-sv�'YW��V����؍Z�Cċ���I��*�n��۴��J?��i�e7�t�A�dx��23�YMZn��'��ݲy��$���H�p	�Vt�<"�p_�2n��v��3�O�r%&
��3 1�)�����G%�@1�(x��}u��W܂��R�H��S�0�q`1xJ&�4tRL/_7
���%0���u4�c��H�$��NW	75|t�g�&F�bKZQ�V�;���/#������>�B��9�Gv�ٍ����^"8���Kk8:T*�i0z���E�ȏ1D̃�2=���[QU���>E(��BN�;4ID�!B��!vn�����#!�sCК|j�0�ÇT4�>���E��.Cuƨ�|nq6㄂���8����FEWM��i����$iTj��K�AS��^�G�Q�B�M�^�Ѝ�ACo�qΜ����,� ����󗝳PY��E�jژ��ѫ3�b�ߚ~��w�sH����7��,V��� k�7s��������t�er��l�'8�q��"<f�~Àq�T��ϩ�D��FP�k��r�;\u�]�U�X������*�<�L�$��>�&-���^�㙢4w�փ:<Vg�[��vz	�Le�U6�0X1�@'?��4� �*wʲs柞��H��<Y�̃�_!P���E^�ܛq��C�td�|���s�6���������R��gV SO�#�W��v���e�Bj�������h@}���@�h\��iR�0V���~Ĺo6a~+Lx*}U�9�đ	Ȥ�T7e��ȱ�푥h���D�w��Z�N�&yw _D�!�ϊ"�N��-֏��0�I��˼ѽ�b��
q����\�ά���T>`ԯ4�?Cȣ���#��C���B�-�A!"`bd��߮#�:gI������i̓�Ű���ug�tPcz�}�4Ϡb�f��2Gv� 8�
]�F:��n7�qI��x�,:��a8������b��k��ޥ���M�����f.rZ��y�/�\8`��WT�q������o�'3��nvu�,�*�������#����Ry�'��0va|w2�)b�N�[t���i|��}��T��bf������]���{�k�VA�BN�����d���<��~���PY4�/����t�e~B��|����{��_��9̈;���R7�3~�q�DV\�4~��=�x��S� ��Æ&�niW���	�|�S+��!��2���c �="K�;��]��������9V0\���)�ޏo�r.�'��/�h]��r����?����#�i��~��<֨��m�h�!�/6 Z�k���Kn�A�M�(B�`�(���ʩm%��ib����Zǁ/�'��u���MN̆c�dQ���SV�8����u��z���<�w�0�2�a��Ǝ7��$�~~ִ��g�ڻ�:�1��G�I�����V8�U5�_J�I��T�4Ar�_3�suOF�u9��),uo�.ȈЊ���*D.�l��׷�J���!^j���� a�eGb2�v���JyJ? �bX6��"�ǌ�7	{c/n@á�UIl��R���c��1*���&�Pm��.�z���C^��pj�}�G7�}/�*=��HL���[�v��,k|'�#�k���C)t`3�2F�Xn��B1sK��r�[��D(����nfޗ�:�� �
ٴ-������S�%�̞tq���o�g"����,���n7�+jI�E 8B����wHKx�=�����d�:~���{Z�2�M��z�F6תgs���Vou�xޟFE\I�9P���ߌ,a@�q-��3cMI(��XD�0� #����*�y�/vFlR�^2���)I���d���T�U��]G ��r�R���jFW�#=�"n�sM���TB���gd!wx�v�޶4P��oX �Ձ�sg��}�rDBk�e+���Nt�!,���h<Eа+g�y�ͦ(�M�IA\Go�T�H��uSƽ��J�\��;��W_k!T�vbő���8�^	Oe'�R�IU����s�$چ(�<O��X��J���\���,s��q�����^�e9;m��{�"��9�P�o��]�BD�'�S�G��
�3*G����2�ݶ`4c��&Y��ԧ������Y����?��}�r)������� P(�6tz�O̤���Y��[���&΀�� ��<O*�[�9����i���5U��o��g���y �w`|h*\JxȽ�"�F(�u^��7(��8��`�Uϒ��Or����Mv����t��ͳ4���l_MŖ�� �Y���Z&�U9�EUd^iV���[�t��ZSW`�̒���y��̻���qR�-���G�&�~dP�Z�����z�ӫ���Ƕ�$x��'3�8��~��e`�li �
���ɂ�lhZw|��& 7�{�;�ۣ�t@M�����;���=��B	��Mh�As����լ�eu�Q!���D�������:��(s~9F^j��YJq�ޝ��d>؞b�ώ����﮼3�g�5�n�'��6�r�����B�����!>�_xO�Si����.��-�3y��v�I�X��uv[�m�`�R��DD
S��}�޳�2��ȇZ��n�m�8���Ly���.�*�r)ڏE�8
]�6E��<�K6��F�>B�QыЩa.;�^U���7��M��5��[�n�~"��њԡ?��6\�э x�'Q�ZEY�s���jI�^Z�]y���Sh��ǯ%N��j�R���'�0ʱ�"`�E�c0��/r"�.�F/jW���X��=����s8=��͏⤩2���M��1��W�I J�l��v�:�uՎaE��`�φ?��*�Nn˾��K�I�娱s�}Uh�Us�C	+��w���h��Ko��H�W���/̃�4l��*H����ڔ�'B�!�<S�2�S$)M�`��p�6\C�EI,+Ȝm�/v�~g&��wt�Ǿ��s�*5�ղ��ķ���WOl2
P(�
�ၵ"�`��\OSM�D�Y}�/Ʉ�}��� ����(��'�[��b�0�{m�SU��UаE�F�ʲ�⟷q1���=;���?oN�;w��Ů׍w��`I��ݠ�o(�*��F���J�'�����h�}G,�l�nn4����P���D�+v0C:^�8��ly�%�4�Y`H�\*Lqw���󅂢��^K�q�e��Rd,BEs^g�TT�b���ͳWi��Z��I3�>��}RV`�m�f�fS�z� ��39�7�v�v�c.tX/����JG��4��@m��w�b�e��ܛ0a��b��L8uE'�^j�Rq:��a0�m���A�����(���	[o���}��ˉ�q��Re�?h{���?����.pZ���^�����=���*��x���r_4��N������5/�Q�/C��9��M�]��{��B��k�9� T�	��	��-�2$
�L���f�P�Z�&��x�~�<�#>�ߢ��h��R���,��vHh�P���v��>�1|v>@��K`/'\ce����0�|;)�0(�k��1;�����_$f�)�L�Z�s�I�c��o��Z=-r���X�uO��5%�ǰ�sn9H�9��pcjC�b7z(����,i�{<��]�߸��ӕ\�:��©ڐ�D�?Z��`��4���Y�����/��? Bl/̋G�x���|Go�^�:*�Mx�^�)����6.�����*0�g&�z�gq=�1�����Է�����Tq ����C)��	<HM�Wش�Gǚ���a�"��,F��
�����Yx15Ԣ�ó|�+�X�2���G+m�G�pA�e�	��P����|��7���"Y���z �;-�p��t���v?�bj��W�c�{���b�P����,��#|�폒��7����lnM�X�%�X+���s���b�Y�cO�iͿ#�D���g�J���߀��'�=G�kF0rj-b�%ұ��r"��ڊ�����&a0�L��(Cl2D�fbE�$4��.�[�b�)����Ҭ�Te�M�A�J�_`����S5�n���-K<�q�� ���)�F����Y#E�H9�r}�!;�_Y�c�Ƅ�U�*�����3�i�BV��p��W�Ƙ;���?�Y�'7�N�؏���٤��h]-�$��A�c6�i
���Jz��(/D�F���t�dm�%���_�t܅�Tf�vn������{	�5:�}�Bן��:��#E	���m��]���Q���#�#D��8��Q��^��a�Aq��} �L|L�x��iz&����y�q88-�V�&�Ƨ\�)��[�����.�\+P +�U45���y�"�KJ���T�C��v��{�9q�7Vb���8�1ʲK'��𦷤�%On��.�%r��z�!�������UJ��!6V�V"�|�`�I D��o�d-5}d�J�ϣ�ф(SP���D��h�x��򾴝n�
2�H�7���aN�\����,3ŗƔ˻�P���|���{� PɲA��̝aPڏ��I�$e��)M�;(v���!�����.p�K��"<���HSR�ی�ݚF����NӪ��GXB�h��|��eF�����V%d��fj�R@��e[��t�Y�&q�9�N�hҬ��=7J+���B |���К�qw����y��d�k�C�xw��Z�	�5������:ޖ�3����o�' C�/N��J��+S�JX���F��=�z)s��ߏ���͑���5%ݏZ���G��&:����z���C�E���^�����*qX�r����bTBh&z�f��`
8�[J"�	S�3FO���ʩ	����ݗk�Ta�J 8�Q\ҺIh��qnv�W����=#g��R���z)Ыg8�r��0���p�"�U��L��Ґ��^��VHh�0*������M�ĥiu����h�x�
�^m��Xn{ �pc��fѬ����'{UW
_-}�~���	[pq0T2����y.o�^�
q�uڊ��n��(�������L����u�{�̜����r�$�R{lDsP5���j�Z�0l�H%���W����
�{X�*j��̥1�P�#2-�#����hUi62=)uʼ����b(�i�-q��ޏ$qM������k���˗�!����I������W��t�o$G�iʇ�%��+��p��p�g؟���g�s�UMyy�����@&��I�VX)78�*�\V�d.^BTq��R�m��T$��oq���z��DU�<-(��t*t>+��ڲ0`5�t���\��s���'�RN���_�������{ʰ����=���d��fl9�O��ԉ��EuB�|ݏ��-�ɹe�e�(=0XYj������5{���ŭV�=(pH2ʾ�pDr"��5zC��]9��ߺ����0�V5y�>���s��J���w"VΘ�g��p����M�u�;+�Ep�=Z���C*��a��R���<����h����G}r(�T�}��y�a��l��ӻBvs��_�� -5Z�c���O��} �OA��0@cg9gfP�ڰS��Z6ƮP���1өAEF�wG���0�H��&tJ��̴�§��IN}�l��v�MV�8' �Е"et�IT՞n"� �U�5KCC뼟��o����:�P|2Q����n�5�}b R�Ľj1 ��"�+N<��#p��9�f��{�!�O���"�'�y��P$Z���Ƣ��+��x0�Sg+Ƶ\q��%�|��N#XH>C{׫eX�����Z	�uo.�mE���O�)�k]w����>��Ng �(e�M_������}Q�]�"=1������x�Mʭ�^�z\?�Mr��W���@��\�5q��k	iK�it���Ȳ󬚕�_�M>�R��QЇ�#�����S��'[�7�ް}�}3f��������F>Q��g��������1����B�RW�q���q��2��|���`\�T?P�zQ��$U���M`���~?rfýW���5���'ſ%������Pvr?S9��oZ*�����8�C1���������Z���#
��E���J��4G�F�u��gm''�3K��x�s?*��t[��E�X+�$��5R!S�q]�x��KҲhD�J��	g$�0���=5��Z��
lQ�J�Ɩ-�0�6����P4�aq3��-�4��ф;5K�Ϯ=q\�`.�k'�
.ǂ_ �OE�&+�Dʝf�}4;i&�;2�����憷`D�b��
Ź剈�:�z�`�Bk�4�/�Hؚ<�8�ڜ7�9����+�TK|�
��Dm �������q
�:|��")+M��|�9��Dj�*�d/���;����p�$�Es��B?y�4�,<��&��hj��)rz�:Ӷ���������oL'�E	 _?D����J	�a��>P	?��5kvt?}�$���!�+J�;-!��ke˴�9�f>h9������E]�V���,��4ˌ�����yПƼ,;���tw�p��_���⧁D�p�+]o���N��q�4ف�V�p��IL 	jK�l
h�vs���ON^+����緪��h/����3`:@��z��!W<�ح]ԭԊ�w�Uw��N慀���WN�^�(Cÿ���ʭ��C��X"O{���8zYZ�nS�2]���S|�	1Jd�~��ӇC�hw��w`�å�kܐc��|�Z�z�k!~I+a�"f���;����<��eL[h�ҙ�M�_!�礏��7�%��z�W��xI�Q�ND<�.��"[��fZ����}�)4�6��;'�I���A��@����֡���{>��m:��<��$GV.c/�l�U�a��}ӆO�Z�0т�Z|b��n��ao�.H�`���#��Ơ��?̬�`�b�ͬu�z1��;%���N�4���pd@�
��S�Q%+���h�;��wΑ:lq�#�e��1�ѐ`�99M.*�n3�����J�� ��.�x)<��Ɂ�{�^�SK$�z<\���J,C<X���5ڃQ�)��@�B�Xϰ����@��u����Z��|��M�"9!3�Z����r�b�����F8����D@~��V��zƖ�)^X��`���J]'�q@�;��D��c=�:��y�GGԠ�I6��zM��1���l�ի��f��M��?^�F��!�@pCj�����
U�T��/��0�\^S�Qt��W��(�蟉x��G������Xh���?e�����J���Y�N2{@��|��+kl�����7ݴt���N(��<����z�)x��/b�l���'�XY��@�����*3b%$s�Nvx�����U��P�\
M6�f+�4�(�l��q�!ˑ8mbV�����Vn��B��Yf��O���($�?����%�����Yu%r
˼08��ud�Q����;��%	��4:�L%�d	 �1�{j��֞	�� �`h�����甝q�I�S:߸iy�i��䥷��ב��<~׭4T8����'+CX:)J<�fo^d��.���#.��Cr*�/A'u]`�y��/�"�MX�Z�H��t)rM�;�����?���{:Z��z֫�0z���p��r�/s�r����r��B�mcF����M;mp�w�Q��1:ўHc�	]'�/*e�D�EjÇs�D��15=�t�BjhR��a�O�r��wod�X�ל�4X��������t%�6���ߌ=�˰�~���O�����6,(��.d<9<��!�0o�^��������K�U�;q��.�1f��b���Z"�*l�"fXeX:3)�ܡ����ݘ�E��?y�lq��PB�A�`��@H�#��l��&����ζ6ߜ�y	�Eqxy�/xF�K����
K�1``�5�`m������:{�LbA07�S���Ui�Q+w��:��E�,W��R���:u?�QQ��j�A�|�+d��e����v�N:Ճ2Xŋ�f�+Ɩ��# ��;��f���s��3q!�q6����	��ˮ��N��=�h>l�t"�6m?���+x`��U�1�y���Olt	���h� �*h9!�#V�u�%���Xf됿Ӆo�e��Q��8���U�i�7�0��Noy2�������RN߬��N�Ǣ��˪C�b�8�!�Y�t��\��@������n�	�Jo}��fn"r̈;���d��z���8>	T�*���7���	0��@��M�Q��ɋ�e��������:���Q��Y�>B�6�b�	��:pj���E���1��Ύ������a��lB{�4SE�'f���x:�آns'�&�-�z���a�@�_��C�X�́�H�ـ*�F<�ab?=ʣt���`��[!A �g�3T�W��!e�e"t�*$�p
��]Ȃ;�݂;lh`�A?曶x=@E�߳���	T����wQ�&\p�+>٬W��\
s�� �Qq�63Fw��h��)_�_�-�f�AP	������FϤ"�:�v��]�Nl}�8�	q��z�6�#	�&UE�z�W ~��5\n�^�_r�n[t�ji�R�~��R��wA�����)	�o�0\\���хw�ݫE�c=�`+`��
q+o�����-|P"��i�駺qNb�d[X_�Z+=�ˎ�J'�;	��0�����u�f�WCF� CEMї����dϣ4i�������Hc�t�Uš�� ��eе�4��\N#nJfy9&�#U���CX�E$7��f��݃z}}��
����c<3uO�:.z���lHt!`��0b�>MW��m��.�۠{��d��,��Ҝ�[:[��L­%%m�ҫc
mU�fгQ��˰��魷�̀��#�P/D_vC1�n ґ�?� k�Z@WnS�6�ݜ^Q��x��?
xnz�M@��LEw`8_�쫘!SI-�V��D��+�� vg̔5�|��+�0�ņ^�DdU��T����q��2����صT�'�js9�|�eP;^�7�,�_���iW[��\�;^1Z=��}�u��ɨ��&�l�F�1��&�0"z��2pB�j��y[�=ȈĈ`��]�
��jٶ4ˍq΁��J�kɥ�g�x�cE| ��m��4W�ECL��BW���ď���ԉ�9�(�dg�o��~�D8��񓛜��b���G�υ��o���.	��r(���K�}��C	*�A㺟/t4��>�v8�XUi����2a���+	=u9�r�?W+�*�7�mg�gZ�phyݱ�N���x��fF��<��C*VM��a�q ���V�&b���6-�4��A+���0��?*4��#��b �����_����n�D����l�ff)���xoBm=��.g0b�ޢw�T�ҧ6��� ��5̏�o-�XTf�C6W�?Ң��N��VL1������3�\�O�����UxE 2�
<��R��+.yC 3���z��>V<��ؼ��7�����aC_�7gwX���?��h%$�mF���g�f��[Ķ��*��Np+"��ƴ1sZ$j�| �zwr��7�~T��R�>����ac+D�P�&�ڙ,���5צBl��9��q+�5%rM�8�X�6׫d~���Wn4]�Y���+����r����yb�x�"ј7
�[��e8���U&U4�f˰�ƀ18�����+m��u��!�L����j]��Rz�f�ޘ_VPp��!�icԸ�cr�2�|w�Q�2���M�6^��O�-:��"���S��t6.� �M�Tf�doaH��-k9N��6��VE������r2�d�Ϟ�<t;v���"��ô����ϖ[�tf|} ���nS#,��u, pcܵw����R"�z�n��К�O:�~��`,gjvX�.jn��lB��q��\?˷����]��h���ݪ��(��/����(<a�1�;��r�jM�;e��DZ�ZBl�jM��?C�"����\��H�[4�B��oS!�qץ�A��l��afw����U�Hi�����Ψ�݂�F��/u� ��aa�$.ƕ|<~K�_qLǯ�f̪r a��&}�9�H!!��`����n*���2��q8f1>����k= ٘��}���VU\�����*�[�h�d���+)^�J��Hl�=d�ǿ�F��!��}��Ӧ��	U��}N�M߰�a��%�}�����i��S���Fz�~�_%��
�F���-����A]hX�
�M=%vΓ�.������rq����r�Ҿ���g��v9F$ 6�Xe5��:�6��h��H�}�L3C�����R�7$���q�+��pZ#��=#r(�rX��9�xɰI,改ly�$�3��ƱU�4 ��d��ϛ��'���`[%������S$9w�kXY�:c�����8�Y���A��M��@�RT`�ێK �U���~}�Ɨt��(/�T[����qWX��rv����8�����	�`&k�Ff�O���#Xʗ�6��ӈ2�c����j��|�+�8�9̄S���'Y1x06|ysln"l�'3��#@#�$����G"U��^�j����U�OF ?��p(%$p���s$Rh��y?������2�:�t�jo�H��Jn@��ʻ��!pG�G)|��`o���O�����n��!7����[����������'��#I�͝�>`3������c�V�X�ۉ������&H���k�W,fZh����<j��������{5�ٛ�r����`���7��BG�={c���R��ݩެ����K�	�s�]��I	����S$�l�V)]}�1��#@A��R�5���eH�E��#���7���HT�\'Y�쬮�̘+�)�/MRHt$P�o����B��Sӥ/�� %o.x����=����ׇ x&�]���s:v*�|r�G	��?BS�����J�M�4�uE�k�@��F��4��O�5¤2ի��p*��֨�*Ա,*�E�J�������)}�p��;��e�v��X�+��5<��L���3���U,e7IUڝ�G��l�6	]�^��E^��j2�����G�.9�(M됕F��KߔfP�l�C�g��5�+�{�<�%.v�m,?u�w=�T���@���.�H�>9�s�\t6�����3
n$p���a�m.�Vj��v��溶�@���<h��l 3���Df�cSZ��	o�ڻ�%��"@8����#q7�r�M����UJ����͛�a.)��V��P�leP�tR,(m?|�s_?������o���{P�^m揷��`Fj������s�p���)IP��!~�뼘��ܮk=�óp�g�n�Ӽ;QK�>s&u�A.�J���yr磆�0"ܩu��k^�FuUVzY�B0�0P�1�;<��t1r/��r`���b����'[�4�3^},Q���@�s+�T ��������aSG����^A&��n�
�x����7�wҋ�4f���e�TAm?vN1h�j�럳�t�o72�-!'�X���mc���$a�wl��)�o]�7����6h	�5�@���ܺ�b���N�"�J)��2M���i����+�� ���wB� �����G_^���W�ܺ����y�6H���(_7�.��Y��-v�h�@V��KW���tt��/q�"�{:��"F�'=��]O#�:������<{��R�H�f� o��Ld3A�ͫee�s���|L���G�őkO�J��Pk]J��U�7����������l�-SzF� �����G��j���� D��luO�W��Ivn��`ST_�E��զ�1ݾ�3ۍ~5֎�Z>/�0�>�H7�"��KÁ>��@(���4�j�w�l?�D��tB����w@��F��"��$��@z�K:����9�,1�1�x��5��nRL�ׇ�R.KwЍ� i<�7 �"���v�w�"Z��������}�H�X!���L��&����P�������g�f����r�A����'M<
��:၈�M�a<`�[�b?ڔ���*�ʤh���^�mf^H�
 V�t���r%R!&�q�<��=�],٘X�f�]S��'m<�Gkɑ�;�Hm��W5+=�pC��� ����G�E���Z�l���QW�w�X�x�aEn��v�}�5�IB�����7|����@����s����Ac��L�G�F>X=o�v��<����㊟��vÅOS�6���Zf�b��wi�P�&K���[˝[��1Ɇ3��@ʇ�[}ߦ?�(��B�ht][���!l�%r��j;��>�0ـ[�&o�q����s�<j=J�8�>[΅��\��Fˡ��L�s�B�Dd^)��v�y#F�p����R[]\��/:&��3T��ʖ.�(��S�FNO�0�"�Z����mܤ�����Sk�ۘf�����������,���a�ʠ�kq(�}a�_\3�?X%~Wm_Y!@7�rSt��1�=ϋ���=��"󉰙�dz�3�6>g����%����k���e��)=}N�;��R�L��f�˻��6�Ŝ��}�]�
|?�lC��l�� ;RlϐCɰC��6�3�x�����w^�k��\tͥ���!y��r�%�I���(��Y�m�8��>=��@	������QBH%A#�(�R� �4�˔�	@	�/�����?Ά��R0���mW��Е���N�u93=vǸd{7e����bi3��0����F��I!�NϷ���9�DuVq~oE(����m�dX�2�"	�U�	��=}�C��^��_��Ϋx�rȀOZ�	|ѽ�wVL.��������چ�A=/�a�)J�TEpS����e5��S۫���y�[��P��qdb��7 �v�[`�0"J��ػU�m�&�`�R�RA�2%��D���R����1W�~!a�j�aAI�����8��`��,�@!���%S�C.���3Pkγ�בq�$PΡ��Z�C���B���-	���nyQ;�W�7�1��ꭹdD����N
|wv�__�>���c�_��(�J�YNH@��]�CU���u�Y�o��v']X�7Ԝ�\R	������Gw>E���z��>�ٜgf��tZ��eCd39e_� ���A�2�V�	�=�I���A�K��E����o]��2�L�����s|�C��}�*�U��?,��S��Y�p&�m��#{#��F�z+F�l�<��g6؀�SB�iZu2&��M�	��IB�HC	����mO��t���r������X3��U���m�v{c�����ƔmG�B-]� �P=A� Nd �f�8N��R-	Xy���sO� =��UpO:$�n,�2�kԘ�M��*�5��;à�݇�*��p6ъv�
�S�<[�M̕mл~8�|��7ȥnI��K�&&��!X�e[���h�z���C���>�9q�É�q��s�}�w�X�Z�����h5�)P�]u�����&⢻�����4i�2q�$jd��I�#��/�t�/��#�Ri�+x�,�@*�/�[r����ljO����~#�4p�=��C��W��31��d��gs�`1�J���0N.mQk�gGa��r�]Fj3�;��my����e��+�<��-WL��ˈ��hۂ��$����J��?��#a����L򻃱������=��NĂc���ܹ,� >|l�	�H��2P��l�K���e8ʳ2@�I�2`���y&�k�O�1o��T������#����Z�B(�&�)�Y
�]Y��Ù�E�fo,2u�-
�^mY����e�(P����-E'H��!�D�Lmd�cs
43(��ׯ�}�i�	vx'g6܋N���\����?k�{6���U��ZA�̮��m�*9P��$!��'�*�`3�ݭ�}0�,����B0Zs�H���į�������6���vư��π=BC��qa�Iܫ�M�q�e8\���o�w9&6
l?�C�D2خ���L5�g�����)+T_z��*hfsڙ;����t�)v��jMsV��l�A��a��YK+`!\�^�~*�@F�������c�IU�r���N!�P
���yϬ���V�#"+�s
6�S-g��g��Ë�H-|���iGI���Ι|Jy��ʳ� FF�d��LZk�u2H������ա���hr]����E�1�}y���Q���I0�1��%Ep�S���e��@46l���iD6Ȩ9�\�%&dʠ���e�=�������r�U�x}�:���zw2�H�}�Nl�tP��4WwMN�&����`eKEc��&����|�4dMC�ǝMw�S��	������x��W�[�qp
�c���z��?*����$�nR����M4Av� {��+���O�/�,f�w fJ����m����i�r#���~@Fn�����1�[�N������Ƥi�W,�P�G��0*��;Q�<��uS�f�&'�h����tS�<�Ì� ����IT�;6�D%�Ϡ��C�9�hb��V�R:7�*��; �Ѳ=d��LVB�7��滶Ejt��&����*�7�Cf���4<���j;(�Xt��z�o�E]�Eb�Z�Y[(-�>O�?�ڐ��1ڿa�3��I��c~Կ���������y��vD�t����!p5�%���	߯��*�D�.3�]=(�}v���<�`���T�w2SLs��t�b��)N���>��J�lQ��}>�0��Ǖ"me��_�0��فmO�{{&�KF%�)\�� �M�$�@�V��W�}��Jd|�O�O��xD�1�r�K{=�=���gt��h@���\u�?�"�b��կ�9�+QG����F�?�g[<����ϐ�C�"[���sBS�C��(��L�XiL)-a�BT��R��Y4�|�5�V��C���Y����,Ԃ�V^x;�m�]���`+@}'�� ���չZ{�hWש���誃�"W���<��9<���\������)�]B���1�j�ϓ�t	ax��Y|�]��k�c9]n䎺��+�+Tzyf_j�� ���Ƅ����"�TU��W����n�(�H�;��"ۤ�T�n$"���b��TK�i��	�IO�$�/��L�=�h�E�0��%1�*rg8��?uD�:`����ޘ!�uK�i��{�!�	��<ʝ�����AA1C�=1�#���-d�6g����{T07<09U�8�ԳQ�&�m�����,��c� �ϳ-���\F0��bR�F�vI�-r�$|	��hZ0��KEKZ�Q�_�R��N�:��44ˣӓ���j-|$�5��g�M2H�`�h���l7dx4��jە��m� JEܝx��8��;�Zoy�)��ל���DP�gq��ؕ5����z+�
лr�­;ޞp�v���4-�Un�c�baF_/��5 �GP3g��B}z���V��n	�7ns�����$�c��`��-���(bZ�ͬ�z2��P{b���ԩ�.�~��7�z�H5�l�ʶΦ7�����{k� �V����+K�n[�˄j{��ƖS�����F6�)�tS��!�e5�u�<�܆1T:C��z}&���fR���������1ip������񿽀����R���جV�^�����m��P�O�(��H8Q0��W-PW�.���̕����݆��t+o�g6m�ㅅ����`h)� �9m��iЯ��v`���rs�ZJ�Gp���Δ*gR�F�z�;۔���7��寍�;m:G�[�^�g^�*�7�xBL��!���)�[Ȋ?�bm���O�w�pm��0$٣T[i1��z�%�3�Fഝ�wn���� u��F�օ?	�̼1v�����@=֍�Xࠌ�!�t�B��W�^���R���8�T�9-��Cǁ��H��v����:!�n�j6W������8Q���R��Q\��J�I�K�C�f�#[h�ʼ�P`��Z�޸oU�i�n��^��)����;�)CB��r���㣋�`�7p}��	~y�dpޘ��4(k�Kf7��Ɣ�Ƀ���E���9Qs
�t�`qYi��N�C��g���H����!1�-v�B�"����0Q)W�91Wk�#P)F�#���q���2(�8�-e�"�L��qga�<� ����No�-.���B%{�`��O��6h�	��cz�l�uc2{3�a(^	���E��|=����·?Ӝ��Uzb��X����@�ŝ�~�ǡ���Ã�P�=�) �����o�s �����ԍ�� ��&�f�|0���>#����l�Ȫn�@ݖBE9��:L��N @�惡�pWAɳ����2"�� F[���䱹ݮ~u����l�_AY�d�P���{q�+��l>9��#!t"��a^s��U�&A܃a�B�Y<�|ψ�F6J��/���I{�7�':�Z�֕K�u������=h_�7���A��"���f�w�<���V�xh�<�y ��[�T�@@�*݇�����¸�")��M꿅�cv�x��Y��ś�O���9���!���%�F���μ(����{��{�r�!�`=�����5�����LԶѮF�o�N���p�VM�g���զmf�����J�T��o�Nf"Y�J��Xchm��B։�*W�k�R�V{�V�}��v�p�����P��7ֽ�m��p�8,���U>����'j5�-.���"����+jK�%$�n��_yhf�E�.�;&��\5*8p��Zq�OI��Z��3��6���m�s���T�j��g� ��F�b��k�>Y�M�����ύ�&��a�����.7��*���lf���q��w�V��96+��cp{��^Ě˕t+��\��
}c�ŤM3?��nGXz�w�/��x���W��\cX4l<�2���V��)�#n��--��%�8�`Tlo�����q}�I�m�^E���n���Vk�۳;���(ɭ`Q�t@:��W`W��Wŀ�h �W����1Zݣ� �o8�Y��-�������\�^p����4�U��x�{
[�0�{j���nڋ���a���MO�|q.��=��Aݟ�8���f������ #���3H������p{$T�~�fu���������>���:ox����o�eTu|"�
|�A�8|H�!:�������opY44�H�R1cJ��{�Nr^@�!�gLrY��y:�ꪢPk��$�ח�yv��/{��O��=?���J��%��[�F�	TY��c��~R:#q��ikt�7;]PZ�xx�Y��`{����]�5�$���qun-��-D��x�y�u��Jw6���py���)\K%Xh�sD�����̆\���п�G'���X�
o���9i}���\ ��V�K�[9nϾn�Ƽ!N>`�h���7��"�S(�8�(g����������z���N���'
(7y���2�<h�X�'N&\��	j�e2F�n�%ٲ� �X�w����*&gg0���o��>%/���U4����)��0;U�G�i��J����x��r��>f�E�����z	oo�B��f�X�z9�q|�eC�V�f�X��דQK�fi�P<�?R{��D�d������:M2O�7��`�wp{�Z����ꎋq��x��y�e���<(!+���1�M<wQ,)(�1�S�qiҾo�8@�p��ź�.��g�!��c�+�[��RM�%'�E���3�	/��g�EG}Kq�g]�`��*!V��W�[8�++�+�*�>i�A��$�_j�v�NC-��i�_j�J�i���<��+����:���7@dq��fC�ykյ6,����J0 ���5@"Z��43��B�tTj�������j��ah��g�8�-fJўH�X׳�	����r]�Z�A�R	���(��Ήy�i,��&|�= ����0�~X���1��Eq<�4�Ƴ,��o�f/Lj�=���Fǘe~D���W��)�l,^�D�m1�5-A��j���Q���jG( p���gɟ�V���k���h��cTsʗc���Xp�v�W����Zn.��s�p���.n� ��g��I�z�.�P��5w���@��[46�R2S�2�]��YJ�c��PK{�(��?�J���K�c�/�澭ŗj��z�儃S�C��jc�$�?�e���h}Ta8�de~�|,�LQ/�iuM��#��N{C��KQa੾k R��Eҩ�T��:AGé���N��J]���V�+�,����b�!'su��f%PsM:�0m����m��hTD㷿�6��w5ʋ槴��b�c��ȯI/�r�?��"z?�6�]v�
9U��Ɗ ��-��������t�U��
����DtaX[��n��ӽ�Ax-����d��a��3�.���X�)��㕴ʢ�h����8^UOTE�K���b���Z��_L�6��n�J��ŁΟ�{�;��8�>L	m������;��Ks�Uף�|�m�f�"Y�)���7����iL�|��`ضt}X�"Z�@�?F��e��+L8P����q�n���s�a��8�[�=k�d��U1����PeO15Ce#�i��:�%��
Fn�kK��]7��󓆁�E�Q>�[�������+A@�ڻZ��4á�]�����6��o���TqR�m��>��۝�Ui(!e�4�`7�@@��!Yga������'�Y�5��k�T��~]�H(sv����=�;ά���md��9�G^H@2��g\4\y��R+�J5˳���B����2CP��p�(�`��:ބU����K����_����6�ߌ�,���ս�����2�����ѓ��C��s���<��m���'�����g:�-Y���n8l�N3�?~��̟�ucx�U��WԆS*����{��S�s�e'r�8�߳������TɏÙ�^]05���x�����M/
q�Q��+a��zrT��w�{��`2�����!�Ji� ��U�]���O��}Z�#E���yHS$�T��� ;"j���yR:��ZQ�7�k�w�gl��機j�59@����!f����D�#�z$hL-��$W�`���CES\F�S��'P���)�H��At
���#�a�s��ò��+y�d?y���=�.j��*�o����\���.\��V�pGEN|�8���5q�N���QN�x"����o��?���g�du��i񼓠i������&��&4������.��o⽂�H�� �,qq���3����X�r���J�� QJ	�(�Z:>�������A1����j-��.����_�d�h��s��D�r$ȼ9�~Y"07f���{�*O9��\��T�	��tG�;�"��0���!L��l���l��ʙ��y�]@_��l5}���ԋ�.*�6,����Ѹ���%�Y�^�p�GϹ>K꾥
ś���o�δ9�E�dIc��e���m��I��Ju�����G�,6� !��l���\�'>�4�Exz�!�k�m?���Sa�u�)W�1v�>��������� ��HՋ9��(;�׹�o&ѹ�90��=@�A@&A�%7B,���7?n���*�]��4G�f���}�Zg��U|A<Bq�j���L����%u�d�c+\� s]ZI�'���L��Gi4�
��#;�E���H�*�L#"RɘEd[���i�P�������;"-Q���, 𢟕��b�s��?g����K�h��ymV��/T�o�!4[~�'>]+�E	36�[t"ƫ���Q�	�L�pr�81m^�Mݔ^���,���%����H���:r����������d�C�����T��Tl���']�7A#p�������\�EKG����,� ��^�kq	ȋ�V_(� l�-k�Z�m'��d>��N\�Yh"��� r �`��2�6�ʷ���lM2�u���;P����'���CU_(�I5\��S�-P��RTz���K��A0q�K9܃�*X��,�8�ɳ��n���iYY�I�4`��T٪=���q���uu��yV=+�Yq�)�D{���趶TbkC�O~ք����֏�����0t��z�~Y��"�����:�S�0Z��r�b�������ȉ��t�R�x�+	R�|i��~ٹ�[{u�״0O$��i�b�h�;�����d\�l@:ɤf�����c�|;QX��^��?ӉD��a"����ZN��T���Y�p+}�H����ܹa3Ƴ�Ɲ&�v+w_:���w�E�<���� ��W˸�<6J馤�\��O�i��'��r�Y��0<�!d+[���2�M3�7LTo��a�`�9W�*Tǌ�	1��#�Ęj$ȁJ�n:*�=Uj=�R�=�F�mCJ���U�뮳���:}�]Ȭ[���R��yJ]��+o7�>��Di�������*ߜ�}�.�:`
���i���]��|w�b*R���������6�9�,_�v�1m#6j��a^X�sV�� !2��`��X/����~� Շ~��Ho���X�-5�F,3�ݓ]q��z5�&�~4_z�S���@1��b�uw�4�(�E���v�� 4���,�Q���@����1>P=|�!�t�Ƈ��`�5��{-��k�n�si��ݴ7}��0d%?�0�Pz�]멲^�&�|`X�Y	Y�"����V��mF�K'�fc�P&�@�$%Q��&��݅!5!i)����d`i%��|4,�l��p獨��㤺C
��8����G�P�ҽ�,4�/�}l��'���	OD�d��<)�aJw�`��<�{.�dc��y�\gAH�z�k��H	��?��%�IE �bp�R�Q��ƃM��bF�m��Qáp����q3�)_��[ CQ'EVp��;.X�Y)�� �:i����X�as�W���P���F2\�]Fz�y!�Y%�H;¼:�O��ݰ8tւ-�5��k�j ����\�z�r�����5/�ɿ��ISǇ~�uǴA����K2��м��x� �ȼv��iژ[ͧ9?C�k"U�����������͟9RӶ���jq_,9xy}ᆁ�@gu(*p�
�[�!y�_~���P�o�^�U.��.��c���+�O�U���	61��w0Q����&w!��<�(������i����!��z���C�"cU)��X����(f��{�a�. �Y�_��EB��+ڍOl����y�T�yU�q�p�қ������aÙt{�\�1J���(F��nX$��y� <������J�F���ebM �g]=w����݌L�0+`��`p�ȏ=z��mڦ����Y'�s�M�~�����J|�4���Bt�en8�^�u�f1G��5����$=���!Mܰ���T4SK��kI�����S;"�\�`2�ڔC��||�Hu�2������A�h�=���f�@o�3Tm��{h���c��V񣌭o�����HS�\i�Si#����K �ZgR�d_D��U��.^�s&�o�О���o��"|�#�K���o��#:�h�����<C�k��ABZ�)PX���O,�����	ya�zs�T؊o�	�#���7%�ͤՒa^'���*c�k�>	z����MշN8b�J�Բ~FF�f0~����w�7��2�Me@�~``�����7P�2�NH��؁���aif~]���~���__�r�&Y��ZKV�)�.�{;;�J��Ψ���xh������&������hex$�]+�q:3^&	�_i@W�AT��o�U��Ovդ|�5����jv�(�Wm�@2��3z�r�����E�9�-�v"��S��>h�^�Qt@��I��I_w�M�/$e����EB�E�`����֬D��p����ע�V������B7
�>y~��u��y����!��F�����m���]X�(��0h%�˟��o��h$����^�G�<�d����+����\����Kٜ��9��
͊�6����+����(/-�PHw�"���\�&5�Xe�Z(�I_�;S��tZ��^#b�ds�l�<m(���\ ���u��;��V��;*��F|�k|�,��NhwL%d���k��|i����aYu���Pb�4=� z!
4EY�s�Z���PQ�y���j��;����w�����O.��xA������ �0o�j'r�Ĺ���h�m���y�q���0�('o\ɡ��{��rޞ��  �G���8�wV�,fX�PJ���t"C1��Eo.No���_�������(YU�&��R[n�����E�~C!��r?W2>�Y">Y�Ac{��tjVyIA+_uWf$�R��+�'>'�''J�/]m�^�T2x\�w��V�|0S@͑��Q,�z���t.����_�3[~�A��	��"��%�
��7�v�W�_��:8�)���i�X�����%�
�����Ⱥ\wʆ+<��/aڐ������6�ĉ���iH�),ӑ�ڙ�LI�ԛ���ڲ�_܇>A�fD`ʧ�׊���3��w�Y$ܟ�L�2�)��� ��
�d7���.הc�c椡O���>����/����i��]�;���J��GƱ�t߄���C�m�<���L�O۸Y<~F�゠y(_�H�˛����	o|䨜�P^u�:�譞دԹ�&��QP���:����m7�UIw���끣G���1~O:����'[]eƴ<�س~�}�4"�i��X�s�t?�B�5�ð������3�r�:P����k)�D�m)�1n�^�ֽE��'�\G��K��m_C���+^e����=V�g��z&��Ħi��:���y��p�`�=\� �31�	�$cI��"���7��j&{���|LE*��cqƈ5�2)�_��n��Y��r�ɜ�O�,�nD*��x4���W��j"W��T?p�����6%��a��
�~�!����p�44q&�	�L���'���sW!� *즷�0�t?'�T:��{ij4P���Ԙ�t?�]G|�3�F��.5��d��3X>�7S���7�FΧo�H�&ж��`u���3{��#� 8���G?��i�:����Ad�q�mʠ�/wW?:�-,�9o<��Ow���۽!Jw�W�o��ʊI}���o�!�C������� ����\{��4������r3n��c,�U�P��*��c�˩���.O�ۮL\��W�s-��Z
D�xr����Q��3G3��%�����ֶ�z@K�݅Km2Ƚ�jk�ޞ+�tf��j�FhЌ���i5�@p\n0�_���!'m��A���>y����#��� �Τ](Ұ'2�}�հqKp�`)c���sl��#�3�)6_O|E��tX�|0�m���e�DZˤ��}�^�Y*�Ŋ�J������Ю�-3�����_����(P��s,����ou+,�LI�*M�j������1Q��q���!BH��0��A/Gn������V��)/��ó�ڂ��Kb}Z5ɷj�>&��z1�H݆��80�?
�4��+�^\@#y�i��^	�0S�
7��9�y�P�-�F�ͳ��OzHpã(��I�:�����Ԛmi�D8�ŝ��9l�	�$U6d��|+q}�|pJկ����2�|�=Y��ϛI��؀�|VDj��������y3��W���(`�3T�m&��n��M�T�Jj���&���
��b\Ε���܀qf��"���k_?۞�*�F`�!�DY���4��i%&U��n���2j
�@��J+yG���i
��i�wS�Ѵ�9�a�Qf� �,1�( �74z���	ˬw.���d���i�]�[�b���L��і^Bk����b�$���,�7�$4TF���]���
iX���$�E?;P;eu8j��%Y��.�W2���jNA��BM\u�L�j�^�]�2��XL�Z|6�+w��B�������-��M�[�K�C����K%
�-���pO�������/�5ѷ����a�Ʋ%�o�"U��3�ݴ�-
RDk�F��ߜiqF��3�kg�$ލ�1A��7o��Q1��\$�]k���'�	f���,q�邩�GؓE�
��u�`O ��/nX�I���F*��[��^�*�?�i���O�ê�1@:*�V����Mv�0H�>|�i�w��zx
�{�GW$Yu�����I��/?��E����#-���&g��:�	�6�%�F���'�\h(t�]�$|�������_�'���F+��7��_�/�J���X�k�b,+��zKw;����*���8P��%W�6�T>R9�8�w����d���x$��^S^;Yi�\s"�T8�{�(��#����zH��P�E�?����̐,L�*���8v���1r����nҸ�ە(N���xі��f���N�j��M�y�SW�"Q7|�Њ�g�V� �l���-?���Е 2�V�۞'�Ѿ{��[�`^�ё�.:�D��a�읻V�]g�T�U	,{/����ǻ�VB����S0��N�3g���5�t�Y�����(�H3P��^w�������Oz3��+j��e����}Q�(^)��ת�9���:�t�WCRI����N|�v��Upb�� _C�+�H�>ޡȳ>p�ԑ�v��A��g�4�L�ڲ�]rpmU�O�X@�JL�"|�E{|��ͨ�7���&�A:Q@A�{3Uy����e��)A��
M׷�pxȌ��Y�Tqnv��x�eԗ�W�b�@�WX�7"�i���2�2c:�횊dm�i��0 ��7e�p.�t�B_��K
�m�������%�Ek�J�x`+e�󕰊��zJ����t\��M拚(��z�|}����E���aC����SE���-np	��%+��<�G7^��1A1��l�U�ЙcZIeER��f��x�in���ʛ��֯	��I��?,aI�W��Mb�U~2�&Ux�*|"��F���B�]G�G�*��A��y�ǽ1�T��M����4Ƶ �I�*Ar₱s�s���ՂV0A���RصlF9E�?�8�������属��0�
If��_|��)�9&�����n�1��l�U�=9�1)�f��
��HGĎ��z[�@L����cO���)�aG�W��Ƭ��~���?$D��QF]&`ϰ|"�<+�:�&yߑg9mka���YI[�#�R�K�`��hv�XAӇ	��=M|������eҎ��_?@�B�Y�a�v����p��N��u��sC�Ç��������=e\\h1��-���|�cv��]��S-�!����AT?	r96��xd)F����q-h{/<��V�8��`�쵟���ht%��n9ADھ��u��}���"�P��Q^����RԑPi��m��6DV�V�����}6[�*ϱp'��b�R�!~|�E��]�L���ï�N`�s�����_a�_��7�m��c"���)m����/C;Zxkx�h:�<C��1�g*/�
�	�6tD#ޑd3/ϝ�OL�˄���}��ϗi�Ҟ��t
�(��L����9}��|�Ox���
�Rl�E=�F��J��W[�U�4儊?�9�G�n^�r�e�d��`ژEf����T�>Q �i*��Oٗ�묬آ���ߥ�!��:��>�\x3��]�iOX�o	<C#��;��5T����a�����U٘��vrQzʛ�]����pu=�}��82;l�69XIQ�vނ�s\��1�hݻ/w��Ot����̜�!��֪w�z�~�:X��2�Ww��{~S��0�(o<���)F���C���k�(��Ϙ�����s������G��Q�B?A)2�>C���ʖ��|�s_��a������ş
��c��ת��+-��_�a���,��"�J���=�L�i<�ӕ�ٺ��B��ē�虖Cgu��0sQ �ѕ4�������Aj�2B����c��?K��|���Z��6��m�QpE�9&�{�����=��L���w��I6&�zR�gq�rW��<ܩ���wħ��JZL����߭���e9e���<DTd-s��?�1Ah
��B��"�΄-�S����P���!���r��/�"��hdԮ�(��{�r��^6���c�[OX�w�l��)�)�q�x�_$?܂=G=K	%���Ro/7+�8m�,��}=�1g�Ζ,�ʞ3����.
{^��J�4��n��3���iӌIaH��!���ފϊ�7+�Ę����T��N+!�ha�I�!v�K_�Z �i������^��)�?2�q�����
�)��	��A�K��N0��&2�<�@�B������]{�#(7��w&��kE�Q�ӟp��Uɪz�Ղ�1��`��Y�5H9���Ur�ļ	J�q��9[����.�\B����p�����u.!6��` ��2@
� *��0�&��f��u0�ݒ��KT�#�`��T������YD}<�-��9�p���qjIJ	N�$/_c��Rv־av-�l�J�0��"���ViqD$���-�"[z�F��z�������j���V��U�N�ȎBx�2����d+�њ4��a�R0W��w ���^,#l��X���+��SB3������j�hy�̷FEO�,\��#���`�qga@��MRh�8t��\"�B^����/�t��G@�C���:�4�L�R�-�GP�������Gi��h1����r�.���{Z��Ѫ��C�������E��B�oM����)(p|���)�����H�]\�b�z���2Y����l L��2�o=Hc�9��w�BK�G��7%����W�}Jy��3 ��ȹ�<Ev���׽�d��,�^�13"L��m��=`"��eM-(k�x��= 	�BS܎wr��e�e���:��^��;�<��.��y ���Y<l���F�2a�zVJ�����Ş�6�1��,C`YvRM�
vXKk��u$�PG�Y5��m�"�o(�fq,�I�a�K�g��{�|�k.v�䌉.�������"ojX;��
�~�x���|W�~���SPI��[���p+-$l������Ӻ��>͊Ee-�;�g�y)N�?���#��_�WD��O�Y�Ś\Y�����7���S=��Y�4� ����Ȏ����j&�"b�|��F�_����pI����S
��D���y�,�� *VH2)�{��n�0j�ȸ]qO db��)��3�H�._�,�����'6�8�}�'�ƌ�W*6��w��J������L�\�R]K�[�p�Ƶ�m(]rUf�5ޣ��em���^{ߠ`�挐�� �9�DS����xdx�)|��M���8��>{M�wnXS�H�ۂ5G��[�(���T��Z���=��41؃�R-�Cv�R�4�+�J2�#�%��a��R��^�`6�K��R �2r���᫑������r�� U��i﨩d�ru��Wde� ��,2�DO)"�ܑfgh���oDDH�܅�U�5�G��/%F�dɑ����r+���E7���Q�v�Đ��_�ǯ�Z�)�P���gR"��Ј��2ԕk8�`�٨[�G��Q�.9�,��HD�H2�"�0% '���! ��~6�rf�~�����[�$��ɮG��6g����#�Gb��̑��2x7�BCVd��������"��K�D�AfN��D���j	����z1�K���.;��m�5!e|^�;��3�h�=�ӿ(N!��� ٵ6�p�D`�aёd�y��,���ZG��/@ʱ�Jm@�2.r�R.�<& ���'��z�t���}�rߥ@)�*;i��9����>ƷP�Y)���r|��8)ME�GPOb(�υ
c�DӲ=�$� {ѣh�1`Kxw�/9�g�.$U���vB�*�r�0� E(���K����,8Me	Vy�/�Z�H�e�ro�׫є\QI���_x6�H��`B91����w����˾�'c�������Ȕ��
)�,�6,��K�qd� �n�M�1l�q��t�A5�J_���� U�u�>M����(��"���%f���}�s�YM�0���iI�^~��P}�A�Zp�p�mUL|}�/_68�fR�c���y�h�J��:Pk��TN蝟FL���Zh��L
��MM���{�{�]����� �q��jE��ח?��7Сv�}�l5'��{m�,�~x.P<�3�G�~Wb��_���[�Gj�,�)8��i&۩�q���k9�s}�(�� ��g��J��{�_;�5O�l�T6�B]�C�>�;�k��g�N�D>��~�I�l��"��ĈS��P>�p�����ej,��<ҙ��ڥS_IGP�Q�?�b����d}�i�Sa�Ӛ��=���!��:[�'�*C�W�duUبK��5VD�F�3^��B�<���2 c�5*��ezR}h+r�� C�UNB���Mk�w�3���I�bn���!N��YC��=>~]���s+w���|�0*z���O*�Vh���bF}CUٜ!iPS[/��Z�Ѝ�.sʝ��ͨN�
�1�ZQ��;����,7v�/��S�8��Kx�vZ)e��4&[��V!�gba2S6(�r�x���-���n.��RG��Y}�i�N����F�YM(!Y89���j�߆�4-�o����N��MZܶ
�������Τ��+�l�����ñ¨�n�y�M��zu�/�ƨѡ.��)}����8��5&����P*�x���a�;J����P9Q�\a�`p���U��I2��xJ�~I�&R>�29�$\���ů
vr�c���2���$����}�P7Jk���˜a��-�\���#�I�u�-��%#ۥ�u[�!Ru��<�ْH�ev����]����������`L)0� CD��N}*���ݫ@Rh.F�!�%�]8ּ+O��W��R���'����s�}��cF�Y@r��bT�Q�R�QFd�'m�5����I=�|��ⴾ;���&���|_w�4�)��1�TX{����#l��g*�a�㩉G�@�P�u���4q�g���[�G8�x8�P�m0��n���v�±3�h1��=�iVw�t��!�`��>^k�f��h�:��+�vMI���o��)�y �����Q�9���(7�w�@>[�����k�w��s f(����˖�7���G��2Lz�0D���qAS
�vnij4,��h��D�j�^_HO�N��i����`�A%�Hi\ �.�ʘz>��tW����q�q/24h��ݭ6m���py	���zc^����N��Ow�wH#�����xv�y�d���$�J�~���&L�R�M _�r�����.��A��F�
[�P+�!���3�ѻ�][�c��/X���=��r�O7彈�ˠӟ=�w�K��;��;�>�����Fd,�c�smIe��'N�2�$��E��$�%ٷ���vPƈ�I����j���Zi��7�3��A�}�H�dnN�O4{�n$�O*��˷7�r��Uڼ�<�됭\d^Rt����8�����Κ�-V�ͬ����	'>#�(����j��VZ��#(gP�y1�e-5�ZLV�x��O2�a1=��i���4���ۮm �CUT�p�'��,���1G���w�a��gfwl�0��$����"����bL������?=���|�a��G�G�����.��~��>Y���5���3����b-m�g�� b7��M����&��gS�W�+��ꖎ�!b���QU1.�7׼�8�:�D�dx��'�q��kP2!X@���!��oGUtT�s���P:Or뙔>DŪ�$Q��P��9w��,u��_��޾�q�@7L�֢Е#�<�#���V\	���H4���޿!�@M�5��_C�w��G����*�?� P� �'eD�����W4�E0��7|�0�����F�k*rHJ��^�S&�>���1}�Rmx%���$��������0Je财7g ���1�/�sz��J��4�I
YZ�G�K��(q����Wk�1�������<���hM��l:��>�U��������0�0��V�;�-��1w]�[gw\��G��t��R�pu�%ᜟ�@�)5S�ُ-��C�`|k�h�}�>�T܇qG���^�CC���2r#&�F�W,��0r���a�P*�r���*!�	���j� E�1�ݐ�n���ǅ*j�	oFY�3�Q6���s�Q^(6h�-&,�������u�[��#E�L�_Q�ʘ7���\��ȼ��K�@��jn<_?��H�ϫ��#�S���+pX#X+�M�/�/ꜳ�/�s:�ݽ|%-Y-�N��g�T3�^��K$[�V ��^�D��,��ִ"�>�v_�%��6���Ŝ��ɹ��n3�(��O\�rt�I����|Sٷ�to|�8�)�_��Jjƃ�z]P��8��j�������eД��lt����P��Q-?L�=󤳫��mՉާ);����-l$��U���Ս��S"�v�R"p�t4ʮ{
l��7_ǵ"߲A��2\=�-�6K�tF�[�OO��"ȸ��>������@\���˚�J��,u�0s[���01���a�b$@QA����&�t�'	����Er�a֏��A����S�7!�Pd�����9=y6JX��=ŉBd1�wS����C�{���k�r,�J�I�h}C�ohdpM@aPWS�|�����[�����E���*3R�h�Q���t�2�ȏ�D����d�w[4��KI̦��`�y��9�i�9m�X�
>+���.[���'�)�wb+?$b�Bl��]=$�Q�*B8����o��zu%|mL���K�h"����)����&A�pT\��ҏFZp(ju�|�p&v;jrj�����>b����5|�Z������L���f:4:|}��@?L�t�d��B�& e���oF�<!տ ��/�$1��f�u ���5D�rD�p�@����Z�*ɤ_��yUeǢȯN����#K좻Ί�\N�/ו��ږ1�5�n�`�o���2t^K}9�gx���W�#��<���BȎ�F�eȒ�CE�8�b��[���U�м�ZY�8W�3	tZ��V�,f+�'�k�6�d$G����B��/�2�9
�L��ieCc�S��ޥ�b�3�R$p���X�u/��V�#Vћ��YݒAy�M��E��MI����p�z�Hp[p&�?�yp���A%��.W%\u�\U+�S��))�'�2������L�� �9H��Q�\�>��سʭ����ѿ�˶�M ��ey7+�:M�����j|7�z����r]�JrH~��WJ^H��,�|jɽv;�K��@$���ɾ=�U���U��`��o��R9��ҎI��o�/d4�w��e�0��Ď����2SFr��:N�#�YUW7�Ҟl���g�A��O�U�>���#\8�,ZB6���-�Z�r{��j���g���\$G���D�ړɆUqX�\
l��b�Vli���� ��.�,cP%�^����s���D�P+~к&N��>Of�s�*�dŧ>Xbsx�����+�!ݘ�R��� ��
u�Y+* �/򘰖F`y ���o�,놰=�T^Xs+�ڞ�]1LI6Qq���ڔjG�Y#CT<u�+��z+p'�I���I:�~l�m2Q�z0�p#1ő_�#2��Q��N/����1�9�뙟�2<�]��"yH�0����2��Q�����F}�ɦط��8%5�l|���r�΁�.QZ��zô�q�mp���4v@�h���q�7���C.LApɣ�,�4�仾<|���EB��/�Q�B�Y֩��?c��P��=T���@6c����5��zhc� $��b)��W@��&o^Љ����m���O%��Γ���U+��Ǧ�yiԠ��W$"j��De�Ȼ�W�d�>������&��6<�A�%=�&�f�i����$ce�Q�gS$ټQ�͏0#�p#ޤ�#����v[D��ַ~=���8�_�i��rX�DG��'��(�v$� �?{]�V0�M�{��$�l���Q�'4�2+t߶��.Y2���C�x ��lE����Ȍ�؁��I����p&l���e�=⊠��5:��9I�N9&NúRt݄$(i�qme�9Vc͉K�����00���d흔���2�%6WP%k��x���i���,
РaHC+r�s��jg�4�v,�B��A��"��4��5A���3�'1b$�d�����x"��-�v0zf��-������fFi�eE�ԝtA<*�e��U  �L��D
;qh#sܟ�)Ǣ/J��^q?3%wV�.4�@��a�1��}����	�Q��K�q�XS���u�{^��� i������5�{�匯o�c� �a��b�#�e�#��ή�k����b����4�&;�H|\k,EUΝ@�Jǅ���;`��dH{�N���cB'�D�}-�w9�m��x:@I��;"�`iB'�++*��O��GX��#���1�*/�cI�d% ��Ҙ�',�n��8nE�[;h�`����@��xk��0I�T�*��P��hW�ͪV�J+=,�^k}���Z'(�K�^u�V=����ʢ��U�KګȺ����vBO��8���̸����0�T�?WH/�]m�nURb���K�b)���{E.�Lh�=ͿR�	��8�������������+f��/���+���#y�F���f�k����V{A�b�H�JY~Q"��Q�\�h��z�$����a%�n�YZ�jR{�z�o�V"�S���퓪��|S��:K(�f�r��C�����cm��ХhNu������0L��qOoK,t�\נ{��l`����-��ő����&��x���+R�� ���鐾�����z9�T���.n�fÈ�,�_��kI�K��9�z��]ͬ��.B�z+9��0�]����"a�]�v	SB��T�2�r��P6��^�F5r0[m�݁w�d�i�!����_��p����6�	��|�	�� ;�s�$CC� tV╒�f���w��Z@�k_��"�^	Y�!x̨��K%���o�n֩��z虇
p��쀳��1�5�+���p��]:U�c��^�ј

)�Fl������f��yu��]QHi�j�;�<s&'�k���e�	VI(Z_�����i��x��W�N����~9|�)�a'���O��Bs��kBq������lx �[�~$�HjD��OH&o兎V	ՠc�k��CA[ƌ#7e�k��mn�����<]�=D\U�/���)uwh�G(�~��~�EB\�E��023�l@�kd1$j�/+F��~쎕̓�x�>�{�:,��) K�����h�b��A����ӿ�eL��+�LrN����,��#X�
�r_9@{��?ʛ *i˚��%��C(��R��sϟqн��r�,��{�U�9w����?�-�껞
T�޽LYz
�8H��Wq�k� ��kI�ϸXk����-��P�"���l�`�	پo����:�����W��zpȞ��P9*�An����X�F��I4���.оTp#M�.���qv�u�����4�3�1�ɧZQ�59J�SŒ	,�LG������wHN�~0��fc��:	j�E�G zP�;d�>&�BU #}g|	X�j��@���e�������$ B�2(�d��� �7�BC14�Y��}z6��cZ�K��Zt�u.��g|�ɡ9�
)�(=bXzlg�0�P_����qE��ԏ��_DƇl�h���Za��Ő/�O��sC�.6���`�nA��wL�T�y�C����%���Ji��n�`��Çgi�i	G���`\}ٹ������V���q�	��.�D��i"C��w�[?����
�w
t��G�b��B�5����vB�8G���:�OW���f��/<u�z (^n_	!�&��u����w�vC�B��4�^�j�Tj��s���X��A��A!n���*����^k;<�uL�N�n0��,0�J�v#�Z�	��%��}m�?Xr�3�$���r�Y�dy����f��������A����g9j�G+�8������j'���b�=�F������~��<;�.���ǐE�Gδ�?1�����2��\N㝵�.�|�h�3�-��+U��ai�(��Wr����D&�yE�§: n�<��~����h����)�!%ݫG{O�h�C�c��5�4��0�L�cӖs�Zͅ+,��C[Y��ᵮ���Uz��a��u7ڳ��]sU7���|���%�0�e�r�2�_�|��'f�P_X&����-3rMY�z���(�B��z&fp���mN��%X�b%��J���6^w�h��S4�+
l�,�H��%`��NL�x\}!g���IR��g�ǯ��09��j��c	�u�e��1l��b:�k_qK��2�|�󀤚��o&����}�Z�Q��:��
����^�Q��FZG��OAg�����8lWʤ�<�ܾ����ܬ���k8��2 �ѱ��j�Ԃ�0{�Fc��rV����P�y��l�fOV���h�t�0�G/!��W����%(��XnN�)����}�v]|/��\j�zxɈ��
7r1.��_zEczh�y7(�1�w@�n��r<��2Z�'���O��n�Q
2-�0$�w$��7�;sO�o��ʹ�9\J���HQ�W��tY^Z�a� y��5��p
����S���z<�����r���C�drĴ�������պ�g
T��w`�VQhG���:�f�ϖ�׿^f,6��$���h�l˴�Ɲ|������E<��%cU�z�Zԯ�T.Öa^6i�I���o:7�N��|B!z>O� �Ԓ���a�lO?KZ�)�%��`�UN�h/��Á��>�:Y�*"EY�B�����K�ϭ��K��Eh?��Æ���s�0D:��s�vm�wV���u[.�a��43~�M$Wz'[��Y�u���n�IHy�&��`3q��7�,&�m�2�2�����)�-t���޾ez�9
|H3sg![+JCX��t3�H"�o��8!�gD8��,�=�KYc�}�ʄKQF�@A�����f� �	�>g���ʃt��Y�6�Ax"���<�v�G�����]q��=h�(��2ֿ���}������m�p�@:�]�{�
��ɲڈq�3��N��tŉ��Y�3z�X���������ذe2�]��Na��˽PH�	dZ����A��\4g���L�`l��K�:��j���t-��l:�Q�� ^���z[��C;���1�?�CYsO�0-�P�&�䕶��̡�&�P�L�ZFGfcf^�2k���;I���H�	6b��>����;�`�[��\.{j�y?������e���r�t}�~5!��%�_�s@�1���G�T{�%�
�:.�Zm����Ûݨ�F
��7 ׀����X�Ә������ƳdDJ�o.��$���A|���

I��Mv�����i YV@�oࣃ-���A-�g�1#1B ga�0�k5<_�3�j�����%�;I��"��g�o�3���l���@#z��r�t�؂N���?Շ[*���D���5�,6�����S�$ m�YU-k{H���
5ب�d��8ƶ�E�˚+��$�5��
���fRW�ʲ�{��h��'H
]uC�9�l��iD������x��1���o��k������&7в��޾I\ڂ���-|���՞��k�@h����kY�dM����6���
r=�MH6�\�!\��
�'�{�/ɵ���aa5[[�Cbo���- ��Le�\ԟ��_��<
]��Q�nY�����(���s�A��d�_^Q�7ʠ&�vV���\y]�M
aH.j
��#+��pG�����A���46x�[�X�"@�W�mE/1WL8=Q�Xc㍼r2j!=k�r�Lp*����l^�n�+���B �K]C3AF��6�- X��oӏ��6���u�\^�K���;u+q� �8��DQ9%�X�o��pr@��@$ځ�,[`����d���+�^��(2�GW1f�L�,��MMT�/���� ��Ϣ ��:����T�I�
�3�Ս���h�E�~�O�|�u&<^���Y`'� B����:2�s "=ې�jm�|^2�?��8;����Jܨ�����r�� �g0�5����2�����<���i,�\p	��l�=�頷���	3ipj^�DC����9�o���ʯ��vAU��y�[�>�i�L�w�P��
���V�b U5)vg"���r�WS�Z��*�\��f�o	He�7���\��P���C3_�{��9�w�[�Ց���˜� 
���Oz����q{"ɰ��ܕe���Jh�+K��pn��-E�m�G�����Dn��|4�t�81��D.1}�����N����/M6��Î0�P���Qr�,@����8j�I\�����U�;\�*��)qd*HY�7�̻pӺ;H���'5[P����{M�v����RxȔ7����#�#�/��+�'1�!�������@Yڣ:	;��P�K�+k�N� ��S�P<Q�مJ�R��nn�����WM��m(�R��J�C �;�z�ܝ�e��Y�ገ�qPPo�����أBC}�nf�L�_�����݉R����Iw&{LA_Ԫ�Y�Fdi��
�y�Z��S�[7�0�.�T�&�k����}�M�A$���)m9s���2<U����?��n*��<����Pxאq��E�
�_c �KU ���������i�5��Q<t�!�-���V,�p�)�X_�\��k�����\���b�D&Bߐ����t�� �6��tK0�,�!I�N<V��H��J��$b7NH��P���g�tX�kl��8��[5N�ݢ�"2�TY�B쁌�7����#�b���^O���8�P"��c��*��;ht2a�ѬW�%�4�U��T4}��-x����K5s�jiơ�r
2�����g�T����Ţ�49K�4u��_�*ϗ�Yp��@��a�6�8�P1H>bX��B�����=�U<���^/�ڭ�K!��++��_���ʾp���@gC��z�q^�4���c�D*� *wyYY��A�Kp瑁 O̿pU�H$>�K�c1B=B�����.	t�Gz`ng�VZ[�6���c_�n\�Yο[��{П������T.����3�QI���k�0�)��R��R�գ����G��ӫ���c��k'ҷ���T��c!䑠5cB�U�#k���q<�4��ڨC#�8��\8A]w���7�M̒�a�#6��A��h'$1���4���Y��?�@�����f�3���q��	=��^F������7h=j|û�C���Csk� &�j�/P{�9�����ҹ7�p+0h���8Ρ����Q(�EN���X}=��(�a��NU�wI}X����y���XŎ�']��ԅ��s��8$�Sa��22Ɯ���l����9�&�*EDed�g�t|�1ԑS�=���ʢ��ĝl�
�n=Nw� �tT�2�=�Bϩ��mc{�Ju0KN�f��������%>Ŷ�33�nv��Ri��4���_##v[�i�R�(��Yļf�"L|��.�n�:�j�u��5NU#�@v{)�"�ɎN�|1�a�g����o��*IJf#����޶5�K����n!��c�<u�Gso)ݗ��n��jd�����tj/]��4=;#ކ��nFH��`c�5��p�cw���1�z�{St 4%rP�)�}:�W�rH7��'֙-q���R�˭� ��uGCM�2�C2���������N�W߅�+o��D��~�۬U���`���B.���:DPD�,��g��Xs
��f_	�m�I��9��N�DWR�xA+v�V5!��#yP�i�{h��3HZ�W�]u5�y��"C��ɛZm���W�V�u����V�_�! 1��(����k�=5\12t����A�9xm/�g�YL��bV�a�Tr�tȾV݋���)��9Q�?�`�ø#Z2�HV0&F�
��Ne��0�����ѣa�����w�7~�`Z<�f0����8�F��|�gl/���g��d��^bqc{�z ��d�P:�r�ҩ��f����?*:�r�W �����_����eL�]� ��V$���5-AV��>ZQ�=��O�N�uS���0�����ā�Kz�?�o�&���>�Qr����,>�
&�v�dXo�a�a��8��%�cd��� ;l��%�� d'�JU�-⌄3�a��H�-G|���x�����;�	���*]�1�\���
�>ݒ�J�K8Ɉ?���B���g.I(JŨ����>ta2l�'y��o���x�6:�ꪏN��hp��.���d�CcK��5��j��BDT�X"�(��z`*K�/�Ϫ52�:D��<�_1A���:ɠ]c���}pDπ����,8r�
�7`�p�[uH5��9�<*<'�yw^xR��^���\�+���rwr����t�~2��W)�u��]�����áZ�q���]-Iv�+|�&��(����_s�O��,���ߌ5-v���RdX��2M��k��e�j��y��j��̎8���K�����Ō�S��m�.8e��ޓvރF+�9LS���X��Q�� l�x��Xx_�ڥ�S�B�%L2��Y3�H�E����f���#SA���{2MC"-�ۿ�64����7����d�4�x�	��	���Y�������8��?�A�'�z�&��XQ��Q�3�"����a��
�9�����ȾIx��t��ƈ�
n�A������g�3�ȽOjas�Wg�wh�#�\˕�R��̓�O�8ʲ��O4otE楉Z�(H�}��μ�p�1> �r	�تYәp�Q΋�y�Ez�'AyR�T�gɭ�Ķo��]t�`΀|S��fy0�&��ݤY4t2�@p5�5Y�:U1�����	''�r�(�&!�����%��4�cv��o�`ӈ���(�:��F�����k�1Wi{��2�����~�$\�����h&E)���#����uI��f��^B6�����P�q}����i��%��g�6$��(Y�m`U �-6:� ��
�H����wgI��L�i�l��QW���H��f�@t`�z���Hl���ȿ�����&1�
�Or'�;�rv�
�a����(�NQ ��'�h p� �0Տ���{�`nA���]������5/Z�^ �uHԇ�6��^Q�����'� '�bQ.�N�e	�!j�כ�,wћ���>ً�����8vxЦ���3p�t�;IcU8�ry�W鯷}�0���ڄvT �3�����LO�Q@�&���]�UN:����G���i����D���Y+{�0v��6���O�-��v�=Y�b9�[���l^q�Y�*	l��$�̀�s��8�3��&Ԗ�ܝ�;z�ct�֫��MPo��Q����-������{��&�+��5�C����w�%�V�lP�h�,��d��qnF��&�o>����GN��F]�]��p�I�T0��˘��vݦh
��d�t
����뾃*5���Q�^�6�=Z��gtm�]ybJ˻~A��qrg�����������ϧ}ދ%���e��yV	�E$��f�Q�6�� w��.���'�i^Q������#����N'K-c&�aj���3;\�����{�%<��E�C��|5�S(A���,58�Q8�������%ш&U�]l���v���l䄉kݞl��\��Ms�:�R<��`1�l�k�N<|�-c���#�b�OH���r@_i��Ԁ�-�9�������p6s�D�n��$e��\�;p}O�U�%�,���W�$ٜg�����=4�wB��/CnR0�����.�v_Kd��S��E��^��+�&��j�Ӑ�+��F4�b���3 �(O/50���.%{4TYb~+��7��ȥl�!��;���F���(����a��ܽ�U��Z�x����i��5��w��gՔ">��j��i9a���"�6>~->Un�U�P��R�!�ذO�0e"҂���&��K ��(�a��9�e;����C�c{	�Y�!����
�혿aںyڴ�>oy�<�ۍ���"��F^��g���z��M���#Ԏ'�F�|�˜�2v�w�����q0T��۸X���X���KU�P���*d=�fa���0�o�g�i�2��G�Uh���2�l�9h��Sy�fR�6=���4����B�U�`J�K�{+/��/�D�E9ɼ?���r�ۛy?s��)e)��V�G�^��R��`U�\�L"D?�Cp��!;�U�d�3���S����r�R� �M}P<H�>�vHD�![R#0�5<֚Q�閳j׈�f��kFG2+�Hٲ~�5?�==[H�L�5��[�e�v��'Be}����a.�Gч���q���g�
+�>�@r��̰��i�b�K� ��s~�7�
����7�5�N�?@�Nʕ�ٹ~I������f͒�9�uy�(�`�c�}m��b�7J��f-��7Ȕ�Ch�(���-0a�C!|!��8�����&���:���.u�N1jiI���3��9-�{�d��vG3�	ڞ ��W��T�,��<��b8[+>� ���Rv)|PC+S�u*�Y���o?�7!D�C\���l�m٩�$�Z`�!݅����~��,p��h0�]�d	Wy'���:-�8�\6B����o��	7YQu�,����"VaK���=��e�U'`��͵[�9����V���� {f�����/�]S���^�˴C����O?&�/_���K�.X;5�A�,4��
����;! F����J�d�������֨Q�w�����8* ����X�8 ׳�;b�M�8����ğr(���BܻJϊ]�bt�]��qa�H��j��]�/Ԥ.�r��X5u�˻p"�U��6�Wr@�S噹n�A��mv�{��.9��7�����!%��Z2���AIQ��6�ޫd����<H(�ۯQ�'�C�!���_f����ڟ:�����@�u!X�ơ��nn�!7���ȳD�m�PDNw�5�;f6�l:�X٩A��$9.h�B����A
�\?E�������t�9&	�P�&���*�.�6V<H_���D��P�^Y�s�&��|�B!9ՂA4�Б\#�G�G:��D��C��r�ؐv��M��f3��U�L�Y�2�����y��ࣸt6�,a@�<Q�Qs<������JC�ʡœ����~�ê ��΀��ܺ15]~}�e�f���-A�L����7�����t���-�P�"�C�_1�	e���Թ�F��b��N�W�B��g��bϠ7F=�r蠋�'޽���O�bi�H�����^ gU9On��W��B�w?�Л�W��# �lb;o�t����l��g�SW���8$	�B��>#�.�7;�M:�@�6C��uҶ�����@Y�l�<$�����zzW�%���N���1Zn��>�VPϬp@�4V����Lx �/e�J�����|9���������n(O���!�k�Ye��%�+oe�\���mh�Hvpᓡ���VQ��zG*\�;����#je�� �@��4�^$��t�&��> ��BuAie��c��9��Oӯ�-�ȁGPQ_�ܕ�V.����wJ�)^	U�d�[4�I��f�K�$֚Y��M�1�$O��P;#Y��uQ���Ȓ,k���g4��l((M¥��ZkFWl��G�D����:�Q,�u��/$_΃���0f%d��_����vtϨ#��O��fb��^�p��0��JﾔG��l5#���dI|�+!����&H��~>l����@��:$x����5�6t�׆W~ �?���*�ͮBG�t� ��x�N/3�#��@g	K|������^���#<��O.�A�mf�)��D��5;q�<��f� ���{�w��@SsU]�k����e�3.��C�v��f���enB���s��,�5#��\oĺ�3�Y�*��&K�x�������f
M��H��D1Qbo�;���OPGg��{=�e�S�;��h"KK#�@��L���L40���%��l�4_#+X�3�����Oy�����Ql�b���������ש�<m���z�����քM��m�Oo�x�-�DU�2�g�cD�b諞�@Q9��
�e�yE�L-��~"*&�RQ����~�Y�֚a��?Jy�Áay�Q�ΐJ7(���^i�k�z/�r~�O?���}��b&V�7$�����ȹL��ǦȮ������S�-8�O�}��΃��+�w��/�X�of��m��nl�����v�%��$Xx]VF�.�C�9���-v'E������Fs�~�W�<e�g���	2Z�5>�jĬ*	�j�&A��+<���1�H�ɘ!����W��T5����3[��/Ҍ'Pu��[�(��_��ceP� 7SJ������=��l�&J��@P� "�s��Y�St�"��c\���R�����m�-n�u��j��j+��0Y�B�<CL��l=v�P�˷�땶�%�!��7<*�p���t=.�̌�;�Ϝ&�K���'�9D���*�	8\��dWrr1���P 6��8E�aW[՜�����(�L�=���E�
�*?�f�������0r�xu�eHQ��Z)�T��D�:qT���@d)Q���g�0�Q;��ۮtZ(πk���We�S�Z�F3y(K�b7V�/}ː����d{J�-��m��s�}w��t�Qw|�@��]W��:Q�Xޭ|m%���怓��ДX�G}(��lloY��ҺW��4�Y"1~T(�+E�з��T��gw��N:�;�W�=��@3B�W؛����ˮ�(E�	?(^Q�ߏ�x�}�G���4ڭ�� �j'm����d�0��^X&Bz�O�& )t�a�Ϟ^(�9��~.w�-�"���w�?��9���Hx���2uSU��k�5���GO̡�N.E����l�[jW����h���"��VҼ��3d~�V����u����f�����{F9��:����ӀH��� �GrƢ�oV�^@� �~.�#���j*�y?��C��ÿOi�<�W��^wH8��F�{�����e��tO񨕰�(2Oد��u���{×�LH,ʺ�D����h��[rܸ���O����L�T/�8Sa����JЄF�,��}��PR���{�M��p̣�������S3�n��0�������h`ϸ4V�U���� ��2۷Xj��� o�ʆ�{�ȁ\˫�}wĉekG�XB���������v�]m���qcIss=(��f��ȳ]�UK���#5V�1n!���k�1_pk*���#���c��Gm�jK�MV$�����KԬD+M�����Z�9�������K�n47��g��;��{���H)<��@0r����i��rt����${L�c���?q�O���N�|�|��H���[%w2�;�U��R��oq�����_��&Ʈk.A�S��k� xr�('3���a���S��~ ǇB�9��0�A8�w��y"�(G%�n�u�U@T��~�	U͸��U���W�Z�wW����E���Z�ԟJ�s�2��{��G*W>��Ya�BW��ӝ�Q��t{��RO)f$��e�L��[���-F��uY��4��7CJ�aΤ�)gE���oE����r"�����y� �Me����O싒r�K?-p\n���&��+���	�kJ�0��2��Û�I��'b2��vDμ�\�vP�%E���\0/��2KE����ʳ&�k�j�X�a��	5�>�<�P���9R�� ʷw�O/6N������s�q�����&A7�ӟ���3`s�PL�'���������Jr��U�j��;����y��M:����W�fl�++u�/j|���W"UzQ��L�[@���>���^_�4	>��y)�@e�A�B�H�X@C��Z%�9a�������9{!�}[<�^4�+M��?�� p=H��S�ܠ�q��JeY�	�����z�G(�#8f�DR��<���{�]Ï���Z˱�>�dg�X��|�+���mL���q����+�%�~�U�2
|q����{���f�"�p�Y&��Z�0�����"'���^[���&:6�e��U�2�%��J�S��}��Sj� /k�r�K��e��B�z�lU�I�����vve�&p.���Ǹ��ǅzոTj�I5�v��v��貨q~e����l����г=3r�t��s4*�]����t�!J�U��c�r�k����Tc���4��o��=����C�x�@�j�`i(�I5j�4�<�J���ؐ��#;L�{��X��m��䬁^TU��C6g5g����ٿ�]�n�(�$���DD��f7��ai�D�r�X$��3P�Qs�[�p�bh�@*����"	�sxv������H�� (lBڨ\�Q
����FN��K�b�t���?�|{"h!���T#�j�F�+��zʐ�������͸E�Lib���ᨰ�;���;!�@��>W$���*�ap�������nR��/�5��.�RM�p��z�Z�z~}���M:��/q��P%�@�<�R���&(�S�u��s�27d�7h�IB��M�6r��� ��������ϸ:x��R:n$�G9�z��<�-{>�D_M�H��q�>�V�Q��t%�gb�V�ټc�A�����p��	�k������1�P$��j��3�fa�H�Ȥ����m�g�,ؑ�_�>�M�=dK��#pdU�mSZ����ʅ4X�P��}�?P.%��Z��*����@������I5�e�e	��
Q v�\nWh/4�J>���_:�E���e�jY7�5��a ���������^/�~v�s��$ؽ|��0&��hT�tF��lp�M��S/kKt��~M)��П�B�u(��Іf\+���Vt��16����:Q�V�()-c*	?,떱�%�O�j%a�D���O�Lni�?}��T�7�ܹ�*k�����~\��v)������2M�u��;�B���954A#��Rw7�a��`mH �b�:��烾wp*o��p1`��fE
����@[H��.=s���s+c<vm�F�L�rC�,eM-���=G����#I�XK������k1sn|��Rx�ԥ*��6�P4�krnz9�&?#� ���iz�|�A9�(^��a7;��}v��%w#���3��S��R/#�H��Mp���pt�XmiٝO{i
����d���ג�_G�@O�=�G���=�w���0D<��s�lv�Bk��� 
泶,��2��řd�����owW�1����Y�j���	�Z�ŝү/u?�bF��an�Vиh�z҉�M����ۊ�:i� +h��E�Q�u�k��O��eM��O��_ְ�
���;�'�M�(�#�X�.�_�㴡�7��Y���{�c�N��.��ΙmiI�)�E\����h���D��M�zn�r?�e���9���{�q��V�p>yʒmܲ ���*�b�꠪�Jd�7���ǐ����ZgQg��[&g1=���Dr���7�ksA nNO���Np������	O	�k�BW|�Q@k[���h%�V{Tift-����_�#�:Ϫ~t2���Ҕ�mm��O;v�]@ۥE膄���4"W�Ӟ����\����2&`����W���w��DA���M�!�j���F�_O��rgZ�au���[l��T	��F>��9��V*|d�6�\��Q�O����,��p��1�fB���]i(�/}J��G��ԧ�~��htF�aKw���]�gҧVP���P�B��`=���Ռ뽈���Fr�0��X����{��TƬ�V"0d��0}�I���"9ן�`Ϫ���Np�0�YP,�z�T��5z¸a(%l�C��M<������	3cN�=�M�^���]Y`�&�=ΖO��k��dbһq���f��l\�������Q�ڒa)��g��������q�&��z/���["h�ͣ��g��4fYJ+����q-9#w�£�^N�kL�}�"��g�6\ė�'��ا�Mm��)�CҒ�L��,�JI��2U�K	 V�Τ��D��BC�'�l�3)^���HJykX�.�gI�[�7��3�L�L�4��fR�P����B���5x+��������t^ �'�1hs��*���a{l�eܛb��P`�D�p�B�WM&����FXl��;�}����@(/S/�Z�7�9�F/�x4l甛\��N��*��8�><�${d��}~���X��64�Hi x}�g%�l����ά�S�=�+��1��D��a��;��Z�G�����Vv��G��_h'��X��-�Ǝ�p��X��_�eً]`9Aӌ*��)��������Č�����J� ��Ӈ֖�9����n��:6���G/Aƪ�Pwv��]���M�li?G�y\W�l&��#�լ1"!a��`2��	�g���%���q�+��MO��RR;�,��|����yf��S�ٕ��3!,�V����cm��[|�������}ՠ���z�[Ѝp�oɎ}D�֩v2 A���<�|⯯��_���C_�M޲N!nð~`��1�z�w��E7��b�ܱ��1�������˨*A�K�70�j���Ft�]�#�p}eXH�x�l��&��1k��4G>�3��|�Y}��l�P�s�(�����׊f�`AҚTlCD»��4m0���>�n�^� �1w%w��U��z�qq ��x�I�u�6����]����#���_�,"+�:dW2M�{5�|�Jd�а:�I2�Sj�1��|I��� 2b"�s*iS�u�v�j'�^I�G�<�A����yA���Ax8������7Vۀ�~3�it)��҄�U�5�8Q�Hp�r��.�+��jS�C���GvT��B�$;��T�۰�<� ���^b��-Z��MUm�^���w�
��Se�b�����o/���b�� �?�X��*�ڨ���Ư�Y����l���]���;��c�XL�5�k�醥ɕ������/PmX�\�&w|��JD^�9��FA�E�!=�z�Q��[��
̙�\��(|T�� ��v��\#��Bh�k~�ST�sOԡ�8"v��4Š1#lmkdRs�Nl�&�:n��p��K��}�c1�d���*�O��k�n�Mƙ�z�|y�m��"�x IIη����q5��r>C��o�������z��-y��;�+�Z�0�my�jjd}[tS4"�P�h�x�p<�}b��}߽0�A�L�����i��k/�j6l3@�}'�D�2Y�L_� ʬ*�n�j��o�6��T<C����q�W=����	򚽤�T�9i���@�k�@O]E��y�l��5�
nUd����(�(f��&$z�ds�}p�s�
�RUR[���=,���:�x�~��Z��X��^�#ŨLt��:��BB��ג�]dl
cB�_A׻�g�~r���J �(Wa82��h~��e�)�`LC�z�3�@!LZ�#gv���N\�����yT���MA 	����Up|�V	��M���-�����I]|���ӡS_�����4��$Y��R�{��S�?S'`�s��9��g��50��a�W��a����4��k)$q�K��t�y��`I�Wa(Zʾ��~��؟k9&��|�&�
������O���� ���'f=x���SR0���g 6��\"B�Rt\�2'��a̠(%�}�`\]��T/ZR 4�k�BR�4B'D+7Q�5������'��m�`A؜���=H�q�E���g�Щ��-�&';��_���l�y��'�>m��d���t�Ljց�4N�q:w�X5�C|���'m�p
6^\�)7�X� �J3���un���K���S���@;�6~�^u���&	���W
&Ϣ
�J@����[��o8�r���2x��h���{ UMq�����c���)�zww(�I���@�R�6�q!ʜĺ���nO)��y��i8)��؆	�����]�i����[
!�[��%� 1�˹R��'0�	έ��_5`�9둮���)2��ؼع�'�y^Ǆ��s�fj���H��r�dֱ�f;��"�%�:*�>͟��7� u�H�U�y蒖&PS��h����p�����YHa�	�^U౏EF��fH��O�~3��ڊ@5�GZo�}�Ȭ����5���^�ka.Q]z��6�^��4�+���}��v��0I�!�$"k��@Qyx�lbM�
�3��0E\�,oD�2��7�Lr���A�jbG�-�\j���n@̬$��L����zҾW��[��Z&ȯ�D����\<�x"?�+��N_g� V[¢�+��/�����(`h�oX(�u� �> >V�F�aHb́C���<�Q��-7IնR��ZWI=���\{a%i��Z-b��3��!��ͫf�⹮�X� ��R�7f�{|�|�1-�S	�K�&�z�	�0�� �Dt��^E�
�ױ�r���-?����n��l#�H�8�f���1P�?���]��C}�D��t�TO�9���`Sq��Ø7��R8a��]>���-s���@pi_�Ė�a@��6��!���I��d�:娣�u���Gͫ�;N攉{��r�CV����q^���IhC^x���7�.���c~�֛lN��w����?;!�<��(�p_��W���j"G��S)+������6�'� ���) ]@ݙNU��E�=���I���ރ<8G;�>�g�z ��YM�.[�[J�"(v�F���x͙����7�0~��B�� �C�/ؿ���8R7_L�(f�v�ġΒ�&9+$)l�|F�Ed��Xd%��۽��6e8��*���l�W�18"o�oZWA�¼¬�"V���*,Э.e^I�;$���⒦��Үv���S����
ɹ�ҥ�q�tf�d(�^��t�!:�t�0Ĵ*|!���99�ӓ����]Q�Rx:�Wz[��D����kA��t�?�	�k�i���:>�O�k��6�J�Ϝ�!�SKݤt*M,Z<�h� J�^���ym������y��x���s��ı��a�eb@O�-1+�%�dd����h���?����	=��\����0Dԉ��YL(ԱL�|��ٔ�^<b9��<B��H�|L�r#����q1�i���!�+^���:���*��I}��?�)M�U	a��ݢ���(L%�\H�r����J�Ut��2n��jH���W��ȥ$�4�I�"�6P ��>1̐��Ү�Y^S�೹@�(�k�'�� i�h`�m���MJ�%f�2��%�+~�Rz��P�R�˘!�T������0��[�c�ڿa���* �]O�39�B�zΔ��9Ϥ��(a�pfz�/�,[�	�T�
����~¢̂y��k����?C������!�ݚJ�.K��Z��AH��_
[�fƮ-�k��}4WW�}w�F\��G���1O��M�����om�L���U��0ޑ�/���������M�p�����<**Ǘn��Ü�~��֫A�x�օj�U�L)�(�]�IOe��֎N����\~«����2U�a�g9��Oa���\��O�OCI��u��+����D@�ǻ���3=�X�8�
�u�A^����*�Ah�-�8�AW^�W��w%FQ�Z���A�'1T#{��'���#�qyo����6��_-�tՕ�DC�*K�4Q��`�;��~�[Oe<�6b���~�m�B
m�*���x��߂墥�����S�D"��dO�����4��Qr/���<|9����;{�8���p�~��Pb3k[��S���W� ?�t\S�Dv�x��M����Jͽ][�L荻����5���U�_��z��G��%*�w��XZ�}Z٤D�1��Lw��z2���Y�lx��3%�'�J��m5�P�سQW�8�/Z%g�O4	���-�e�U��P�̐	�(���L}���k�u�K�$�di�����t.4ǻ�/�&��	M�r%�[H="w���+��1L.�s.�!�1:׿���Il1� �E�އ� �Sd�$$� ��M���X� 	Q������9q�F�_Fj��� T���up���P��`~]d5�M;��U�TN�"�sb.N�b�&Z�(L��S# ˭s8�`��dT� �-��ւ>C�E�mhQoѳ^�|ài[�?�/%
�i�]�H|9#�/�#� b�L�w�(��l:l=�m��Md��.9+���c']y�L��[]�;�`�ڹ�S��ϕ:�i�����=xR9�N�QY
}Ô��r�RV�]���'87wb��]����mk0)��.w�/���˩�i١5BZ߲��Ǌ��+���4i��ʱTw����m��B�+;x���Ʊ�h�l��ˇ���QO/�����W�y@������GU!����@V�I^����n�3u�,�w�+DL�`!j1��6*ئ���5�51L��	"�L:�������3�n?XcW4փ��H-�8�-N�h?P���y0�v����iћ�:b�Տw�|��t;̹�3;�T�8西|�{A�t��m���'c�e3��;�|�� �N�ʍ>b���Gf'rU�����]X4���ʫ� ����8mr��2�'�B��@t�$s�Q[E=�]:sˍ�m� �+��F��
�T�q�q��o����iD6�SI�*�R(!A�/0ՠ� ��}������b@�Q<�\^5�}�����eoY� 'sS��!>pO4Q�S�?6@�-Q�Kڴ;�MvBd>h�<�0w��Y�=�> �
���WhyU�/4��X�K�{o�7�zG�z�������|v�r��cr��7�f�wS�����C��WVe$m��w�n��
E	�9*NKS=FƯ ���@Y��oٲ7�ka�i�+ʓ��4�g��
w��q^��L�n<~�6�����J?)�b��]�y�_�{��A��":�{7���C����VG�A��0�Ya����Q�}*� :_f s�,��g�O����]CA�5x��j�.��j�y�o)�i'�f�h��ӌ�Kx�G��i;..� ����v'x���qב�~��a���Ά*��~�&i�tā>�P��=�$��z� y ��hPBa�$�1d7i��@�2<����u�[��Cy-���mg�O�����5��t=}X���$�$�x��K~1�>C;%�d�uǣٰ� ��8�e$Bt�15���M�"]�Qs�7�o1�����-��G���gk 1� a��#Sٷ�F�M:O7$� ��A�Fyt�K1�x}؝����p�Or�8!9�)
S�t�}O���ؤ����>a� ���AWJ>��u�2�����4T?���x�54�{���yWZч�&��"'n�W����)*��Vn�)�ahE�ǅC��b��פ:���m��5�&��0c�p�:8�����	��W #�"�p��q�H�y�h�-�(~�G8�Y�@��n$�����0�d�Pٯ���|��	�ȡ�Tފ햖�=�\@�(i4�>w_��f�g�� ��>���f�߮�\bՕa'��G1�}
O��Yo�(J ��j`�z�ƌ	��S:��
�w���5���;���S����C9�A��f�n�yd���?��29Z����S.V��ϼ>�$,j���11��X���Q���s�6kE?Ԩ�'c��{��M����
'n�a/�_{�p�;.r5����[!��_�	Y�)z2K~�K��dU�s�_ �p�H5Ii�����ʭMR<�[����^�5�Knˏ)%,a~��Z�u}]����Q��I]M��Y��K�-�,b!�l,s�� u��^f�e*	�F??�ˆ�G˛��ȗ�؇@��b�������<����2��M�i	i�_�0�1�]����*T�����Ҋ�
Sh��Ke���Ac�\~I�շ�t��-W��哃E|��ӃԺ��Ԝ0�-z)�Z\��2:�S�~;}�o6K����qC#��s�fڈx�ߥ�*W��Qd�����<��o��^e�5���p�����T��a#e��v����Xl�Զ�LC��S��pq�C>�ъ�T��`��Ip��$��wZ|c�2���c�%y�A�R��I�{%ߧu��.���O0��/��zS"�_%#�c�P쒭!��j��>ɗm��k�n��擞��uI�Ė�8�#���t%=����e���@܈�s�8�zi��h}$W�.��:/Hx�2��_��:ô��O=2G;w���k�C��9c�H�.�5lpfJx	_w��+fqD�*��Y|ٱ���W����a3U�+?%㌎�$��?�p��_k:}��}O�hQ�V"��8��i%�UK���z�|����Ծ�ь$�d�����ӷD�4�s�DG
�[�#������X�W���4�n9�z�,���_�����_G;������������$�6����^����=�P0�A�>���%��"�{�6;����kD�ಅ�I��8]�����S���m�O��cTAm���M������ �_�_�-Z��./q�Uuɿ�_*ѡ�Dfi���I��Շ�9IY r��eI��(GZ	�T;|d2��r=�o�*C��o��/���i|Q��JǑ��Ou-�K�x�~ۈ-;�?�QҧCb�Z�0D0�~���ǂ� �?2c��ٲ-�v�5��ljn�V#�ոXd8`��+�1n� *�Wv�Dȩb������8m�l8�e�5eq�S��W�4̸H�6zj	��p!��<�O3�E\�|/lùmU��N��_�"Ӻ��)�z�ݟ���b�MDf+��v��J�?hu�YT�I��oj`��@�ѿ���>�Q�s��݅5M�"	��>T�(}��ar��a���Y'x���7�L�Zu��1�u��] 1�5#P�#/Y�3�F�Z�2���j�o�^�ڷo^ADE�:!	���*�*,�vmk(\�=tn���`��
VV��/����_�"0osv��Z
�b�s<��-P� ɘ����*��U
�8@�����ӕ�@�Ƶ�{�s%�nԅj~zC��A�*�c]��C�v�?C���e��ř�jG�d|�~Q�Z�y;#�+7��A��ֽ�h�FQ�	5�m�uN�Z7Vo3;`������v)�[�C��E��{@G���A0��B#��n>`5L��Y�_,�h$Y���D�ҬL-��%w�տj%4sESg������,��%��T�"��Cd��G5��H�!�W�������7oƂ؜s刕��j�q�+�	s��ys�ǆ�w�:���O��jB��>��4��/�]�Ղs�7��fdk!�}�C�6.{�4}f�r5�L�}�#@^�렜����T�fr1�͵�,�a��o5�$� �-�$�煔K�S�ʆz#�W���Js4�ѠT2�hT8Z`|U��4��Ģ��u�j��F�}T� ��i�
��ϟ�(kj�v?�ND�l�&�vl�3�S]wl�H�x���>Nb:�~��3�rn��i� ЉE6���2�{�+�=O�Y`ǂ����}"�� o��@��`Қ$��`hL36��J������/:ǽ�_�=&O�)=�P����ag�� F�j��}$'[o��۞������A(��^��j��������)6�C�^v���������%�����l�MQ�ސ��3��2e�����.�ix5��!=�� |ы]^��Q}�a��qW_��İ��0�Q�����sL��9;
fF�9Bv3�)Lw�ӿ������%A���.�+��`�K��e�=b@ 8��+����'��'"�1���3�}b���dU6�����m�~�X�}7�b�۪RB��K+�j��[Pم��`��h&}YK�������'���\��0�J�6ΞwWY>�� s���ks�F��w(I8�7�oKiV/=�Kh6:FNYs���z�
T�z���捛Ko���S�'q��"�w��co9�-)+�W��8�DX�~S+Tf�n�Y^1���z�՝�m:�p�y������23En�X���5V=�d�- }�N$Y^L�p�D���m����i<G�{��	�Ђ$0���e:��1�F���5�k��]�O��{0�k+'���$��2P��� � 3�Q�1�1&7EܤS_��Xk�S�`�i���W���ne��5��#�b#k?�_J�7Y���B���tը�SQ�0�7dc/E�vtM�̗����Y�A�t��ORMӨjV��7��+��ضji.N�1���2�}Z�z&�&��'����B�Pb�p�&�ՀlƯ=I�0V��8���짺�	�(#���+wd���X�>�׌}tv��,�٘����5�j�?N��@!�(���k�������< '��~��i���C�(��{Y�x>��椔Xm,�,XkB�XȓȂ��ɛ-]��2��I����Sa�����*7|��
m m�'A.F]��LR���EF5�v�/* �++#l���˄��+>GhJglz?9��6Ϭ�����$${�D�t�W1æn�S����4��!.7�ՀA�=�m�����Bm�U�8B
��.�qڱ��/m;�Je�g1����-�'
8� Sۥ�f���o�6Em��跢��rϊ� �:e6Y1�5����
� �6�X��,q��Et1(�L�a�����M��<��4=�%���T�"Ff"w�������#�JP�B���\.�!f���>5�m��(>�R���vxP��H��zȅ�����}@���{�*|˂����.�k��SH`d-�&po�
1��X0a5�^��hE)}f�e�'q��չcs[G�K���Q��A(��dV7�ړF5"]�~b�{�"_�>0��:��Q|�H������H�iV�|���l\~�=��GS,l ��"��I���?�طx��q�
ș�k�b��V>����J*r��,�`g�p�gӍ�;��~k[XY��M?c�b��Ҏ�����.�"�	܇���w"�L~�i������\}���i.[7~d,�;u�p�!i�ojP(F���v�"1Ɏ�y�h�A�{L%']��2�^��0e�ߥ���z�P~�N��~$i��ǵ͂T �,�=sAoT��ٴ�7e��ǔ�u�42D�X�zoB�0G	�q��U�+�ty9��Qb9u_�6�;��;{�h�CRE�N�Eb�J�5Ftz���%�#��^V$�������ψ4&x�]��xeb��0����������U<r᪳"���*���̧{<�����R�G���F�-�.%��J�0���SN\rF�p ��uIeOղ����{x��6���Z�ui_�	H�/5�"J�?ョa�7-�dM#���G�!/�1��PB|��Q�)���
���c��`�7|۳ӄ��V�>��2�R�^z�Qo�������?{i4�UN��cI�(ff�Il!���H�!�L~�ԩ�JC[�E�Z��H�z�<D�}���
�}h�Ty<��7���]����~[eAV�0/�X��O�~P�~"����ήF!8�'q8Z|���Vu��9>@��|u 8�dWk������m�Lq���M@V�IJ��B��M۝�'p��H	�54�%i�!��;��M~����N�9��8ҙ�[�7)����������A��&�i饲e�gr��"_�f|f���5�s��)�w�c���58�
��HB�&��K��O��	c��`)���e�?��I?<i3'9/yF:o#�gQ��� {9erc��w�J ALЊ�����{�A,��a��,�8��yK�?z�OC"�|+����e�ĩw�4c3�o"�����k��.��Fj�,ٙ5�	eF�$��SkB�M~�2mlZ9�A�0�;�[e�{h��M��L�s�����A,./��2�"�*�4��Q���,��*ӏ�[�- �����"ف縖�S���cQ7	��x�h_�zcLYS3��Cm #&�Cg��/5M^���hE��?�.���A�	�|gM*���Ȓ���sbY���iQ
����i��i
�^�er���Z���v��v-Ǥ��2�n|f��ׯ���ԏ���n��@&D�<��D��1�wmApQ$8��G`.@�E;�K��c��q����J�b,?��s�~;6��ݥK�a���ԳٗcAh),��V�Q�>B`�[��q=����bL@B�]�u��������(`��Cx���o5�����n3�i�	���y΀�gjh9��pO�Qk�
	����-qB0�}����z'��+;Zх_N��	��H�wJ��U��[�"�f$��A�O�x�)�k����l%=S�\��/��1��^/?���$!7�������6�/�͢,f6"�ЕdDg�GP��tp왌��Õ��3�������tڐ�|�˥�!/А<�5D��� W�!�I��(y7,��,�N�;W��U�%�_��z�����%-Fn�p,��"��=[I�Wtt��a�.r��[0��x�f�"�˜����iW1G-�
�_m��p2Yd�*���іT�3��<`������������9s��2�� INA��5�����I��3����N ڀ�G���������ڑ�S�M�=�s�y��MĬ��[��G����������f	cʲ�j�r_�Vz�M�C�����th���b؃���`��쏥�;��,wײ��� �Ћ�
���p�$���`xav���W&=Gw@�짔���/�l�V�>�2�3��Q�׫iQh��dy^<�4!6"��/�6��w���Ǭ��V/���nRfR��\4��;�;�={/��Bb@Z�nHk���*!�(�H����
��8���Z��D������b�}P��� ��$:�i���5�6����r�4@�|�C��Tk�k���R��"�����:��E^�.�\�?J�C��caYk�h��L�˹��0��R�B�\�r�4�B���O�X�l���D������ٷj<H�/9~�� 8h9|Bּk�i���AlJ�f�v�h`Ba�Q���*��YI���Y%�D3�}X���^i���=��WL�x_�KTcMP4����(��#���[
�|�(z�� ��1 i9���ex��`�q���>u% q�<r�e*��*����Pև�S�P?�ڸ�2/چ���l�\ȗ�c��t�qoڇ�s�얡[�H�����4�"=tWt	Wm'�B+ I�Yi�@��� ,��A�Hr�]�(�8�;0�n4���h�l��b��b\��L^�L��mh4y���(���d'�X�"W֛G5�$^�k�gZ��V0�k��>?*䲳x����	�r��%�U�M���iJ(��II�� @Gw$RzG(�;Ek��������f�t� CT'ZZ��1g��e$x��7������>J � S?���c��F����Z#��N���[f���4�71�j��?wo������/��k��V3C���;B7Tr�w�F��p�B=��;���QU�_���D���C�	%_�oo'��a\�e��7��!�^Uf.c��E�7X��CW��ʂ3����H%�	J��~��n�~�9��ىmw�goȢ��
sW�� ���4��B�#!4��F.f�r3�
[�_}��*�n�4Ș�wثxǷ�lHʟ��#Ak��y��^HcF����;FG � r� ���V�e��:�񬫣�6�}�z�B�W{Q	C٪l������}�ʎ���9� ��*Z�/ ����R��m�mr��A���Ss�	�rQw}�qY>���6�w�uf��[�a+U*o�n�U���I�:9���Y�8a�w�Q�s������ i'=�W�Dw}8M�L>s[+(5у�K�H��-��=��8����T���Q��Ve�L�A�e�hDW�Woψ&����Һ�Tṥ��v�s�� I�W�(�Լ7")
�8j|"��Y��+��۪>�;�SL�:K��ҷC���hq��v>P��� u N%F3���r��aE��9'��;�g�@���nVRhɐ�g�:��?�	��f���;���F��M��La�O����6^z��PK����g�pCe���[��I�ʽ�%���F,�`.eL-I��W~7>��D;#��U�!���g�d���\��;>^������!��4�D��ÁD�p�O.`|W��MGO�ʈY�wj����<�V��Z"�� d�=�U�iq���/�TNz���"AH^�+@h�������+�>7Z�O	 �gt|�M;�Âr�ǥt���e�D<���s�6�AQ�p8��j?���c6F���p���k�׫:-c�|�9�a��re+�X����������Іv6 M�VsY��쯭�����ak�y�Cl`�J�U��j�e,�(-�wWj6;���D�	0�J�@Yڄb���=�I������A�?���#D�r&�o�:[�42Oyg*�4�rgCW�9�-Q�Yw�2��������U��;c��a��0*���T�IL�X�j��-è����%qM ��<#U��62y��U3O�an��'^�ђ������1s	^
*�/�e2ag>������q�k3�<|���^K|f������Ђ�E�!��ɯӰ�f�_���S��α��i����7�=m+̖p���'Pb���	z�Tq|�{z=�rE�ɱ���J�hL��ct������0?�gH_t�^�n�:'�M��^%������i���y1�.e{���e��>�I3a�S
̭qoV.[���ƠN�����NS ���y8�&�,���y�*�������9$O_��q^�t(�{Ag{ď��^1q�I�X��H�!���t��-�����_�ލt�oi�Sk�� ����	���
5�yM���w�\�Ѥzo_��=��M��+i��8}:=Z?Z>��#�D��nxI�X#����C~n�أ�v�յ�JZ�N5�P���Wj '9W��]�[��0-����q�q\�
[Ӭ��\��p�M�ۥ�k8H���w(�$C�X;�&b���$��9y-N���ye� �3���Hd)�J��rW�_�K҄F�4%��l�*N�����*���n��������c�� os���_Lɛ`�\��W�����?��j�h����\4�����զLK�c�Z���E�[.�)7up�ż�,��=45q��?^BA"�����E6�j�������̉��|l)�Y?��<ZuF�Jp4�R�4�P{�,���~���^�"�KG�MD�* @�����삠'g9e"{��՘��*�����ᛢ�\�r�i�_-@���a�xS�5���6R�#���lTʡ��(Z���d:k��f���+lE�Z2�&�|�\p1=I쓱����3��G���
�-��=��DU����I�%��sA(*����Ã$��j�IJ�a�/�cU�x�9�p�o|��e�޻X��+1�B����D�T��lK�4�]w���F]r	@��n7���/&yH
R��t�YY�<�Om(t�_�DF+NO�X��� "��t@�ǟm�:?���]9teLt#vU>֒E��qaQ�O�.�KC@�/'�����K㭟|%t���:[���a�B1z�y�o�_Lƨ�����TE6����C�m?���f3�Qp�+RQ�XshT̈6�+��B@���j��D������Ζ a�RZPУ=gz�!��eX�6N]�����!���X���cqW݄֙7��]8!�ژ���>��ئ�M��:?oL�3BL#�7����D~Z�;�J���$]�=:��N��$�َQGЩ��9"'ӷK�<�܄����X�+O�s�87T�������y_��S2<3C��!�{z�x٢�7h-/C�2�q+��ҫ8W�}�!K�s=:�좸� m��ݒ(�!6�5c�HM`p��5��u�F�2�FJ
�e�F�?�+�[�)�O��R���9[f�e� ���!u�G|���Ց��ӌ�\�{n��A�����tk���lcG����"z^�gh/���xC+b�*��VG��ƈ�qJpf��vh `����A1�{�Ѵ$boԤ���^��͒[Ύ���4�0��k95ӅSCٌJ�X𕼽w��r�*�bm���2>[��=N��p�j��&�pPN�g� "��s����޾����+�b����`>1���V����#����(tS�s��y�%;�y��@_D��B���&v��ճӑN6���'L�p{���yG,��mJt\�KF٧�R�OV-�R�d��M�okl�cE��,žO|����?x�eq06����Is�ǆ)���fM�v^M)��2�)?c�^z�*��7."gB���K����tRa����~�Km��D[w���M�t��kB��)�R��D�߬�ܯ�@�J?<���l��sU�
#+�GL�?�jd?��I�M���CL�\�����Ӿv�*�^����^���xw罃~͉���X��H���vj�/S�Mvi4x���E���ҙ0S�&��� W��DޏS��J<���\�
Y��!W2h�U�W`��[0]�l���U��Q}�&]$���v����f�D�1��c��F�ىh��x�4�I�������c�%Ӄ!���UN�5�(Ό*���eC�PS�t��O�Zn��U`��r.�L��@�P���? ����j����~��l^�8�O�F=�S�_�&��R�h1.�J�>M�/ٟ�*����F�ib�����E~?A�����w���-T	��e3��gg�
/�&!�%�^���?ᅍa��k˘���U=L�����vB���I��E�1�����ܤwE�<�r��m����AH�ť[���I�����N���p�r�oĎ/g��(v9��:���uM)wV���.Ԑ��?&-���k)  ��:��Y�!�	K��J3��4�y����뵏1����~d啯ޭ�
;�AaMfmJn1�ߏ���}��$����Z��b	$��%�R��Ǖ]Mk��`�o f�tQ���T�+��B5&8t��Q�jn��}A���m���s_	�j�(j%�>M��jH~R�T�-�E*�wt���r�t��j��n�����u�憰�e@^�U^������|t|v�Q�^��QS���XVo���W�;��׻ے��6N4̀�{�#P�X`��f!r�U0��	[���2F��;�|N�P#A����%��8���W�[,�8��.S�e���'=&#9�i�a}~�\�0���H3�@������.cj#�������'�b�R�B�#SR��9�M��?�7. Ѩ�ەRvf�S��3
7Q��Z�v���K�wAw����Rd7�v�!�Ä1��&^8`���qqq�r�mQis ��D��67�*T� (��ڒ�D0�@���P[�	�F�2f�,����N�]V	[>���!(�2�Z\�]����͕@;�{r-��(��i��]��J!%��.ML�+C���vN|�_j����l���i5�0��&2|@r��&3�zRs]������h�F�<Z� 4�J'��Rw�ѳӭ���/޴�K������տ�����:�i&h�"�ֲ={�}(�J����U���>��(�^w��K�(�-\��vQ��V�������	8��נJ�w����΀os�*l_1�u�[��$�q�� ��7�o��N��rl3�7�B�!G0ke�O�:3{n��}��O%��W� ,&&b�Rn%m�rtd�OA7����ArGm����x\� ���o��b���k��Z0�^'ֈR�2�- ������V��+����pP]ai�HKg7���=zNU�o��Q�P2l�S��y�ҹpJ3
�U=�	�0� ItM/Up��39�Rw���y���G���,���`��ʖ�K�[�{ZMN��h�`��H3�)�.�h�@�2%�!'���Ά~>	<G=�W]L%D��<C@T�E9�aö-��6���^yv���8FBbN�8���`�ˬAX��J�^��!�#�s;�x�a0d�ِl]3��$�uO���F���6���eRZ��~�-2�Ź~�j ��_x �d�>T����B�2S�][��D46�c;+��K�@��ip�IgR|�&b�k7$�s�V���`�q��C��Kk1�cz��C����"��d�G`T7�h��OtXtr��,�*�WNx.���}7
��z /4��x�흏c�b�`�ҝ�Q웫��ѻLMl_�J����ZU�jj�E����=�֯� G���U���{��m:��zT���lE�1�h�*��%�κ�<�J�>�"�1$_��
X��ӎ��!���3�^�xpD�M!��y�D���� �BU!`�25�����Ԑ"d�`J	� h����� �� +�fޯ��~�ו���D\`zS��&#�!���X��d?�|���;P%���d��`�ĔLMwN *H�bw��o.6����<T��ŗ,p���Ɗ1�u������&�5V�$� O��񸃯��v|�N�s��}39/�иB@�+�:r��kRL��Ԡ38dT�:0tI� C�"v8G�C�U�XF?t����H]�fs^ZEU��̠7/��Za�_˯��񊺠%\W%�����ơ>�(���"�F2��4�GT�sm�����F���_���4�P�甠=}	�E�Z�I�;�:�v���,N��s࿧���0`�}��$�n�%��!֣��&r��z��� �c5�"�W���U0H$��m�X{��b��4��x��E`�$cn����B�k
t��CWy@��	��-���I�n�s�(}��oX��.��,���
�7f��� sB,�{Nu���xf�7��eېd"PF`�i.�����?
�Ѯݑ!Y��8���E��wn�o��r�ny�~N;��@-�j��l�"���3�F� �`;�G����&�&����Ҩ0�O�q�Rm%�dp�D	�G&g%�`�'����]��J!*�vc���FAoa�E�6B��[V� 2����{^) ~�8�m�
���i:Sxm�� O�2���@|!u��NK�k�(ONy_A��y-��/��>���k�E���}��7����n괉��sK��e�!�W	�*���d���6�;��3Ѿ��#wS���(�ʷ�P6~�J�A':k~AϠ�-Cr �=�~h�	�e�1���u�/ydqh�h�(V��i;��ɞ(���G.�o�}Sa3��\�szg_�wB���P~��xN�G��)n�(�)�A6Є�~z�lf�n� Y�e⺍��}YE�'SOy�5GI��-P���)���\���
K���2����(�:�8$
Я�"����-��z{��uעE46�(3��I6z7�����[�D�3&㢊~{љ�i�B��7�gaZ�^�y�E �;O�����]_�p`MC0��2��=S�\����3�������&�`�0N:׽�mL|�c+�4.;��"IW&[�������qo�x�t�s`��� +X�>Kr�̑h������c[Yd���2T�.9�B4�Eܣ�ʁ���������aA�I*���!��-{(`3��<k���]���n�o��2�����g��4��h�@���Z��ظ��&�TU_��L�(7�0݇���\I��fd=@8���z�hJd<ڠ�d����A_fťF"�
\/���2�%�|s[ږf7Z	<G8曟��B��x����'W�����'\?DgM��t.���]/Xg�c��l�f�GV��~ぱ�s�[���C'�4�λ'X���ElB������cV���k�O_�H�$7��@�L�Q� �ܒ�c:������(R�m�4Yc��ԟ���6
�L����,�Y.��/z�l¨
|Y~)���\%�ZbFJrfBZ%_a4w�)���q��Mw/K�ך��~%�)�v�P�<52U�nO��;Q]�/DWBї��<U���\v�i�O���>c��h�#�i�֪X�8
���b�\�Tz�����!Y���G�fB�0[�a����C�ֈ����[r�j�i@�����ƛE�Z/��=��?�P֝H�n����>��]���l�M��E6� g�rUY�z:�cbJA�1������wC|/H>z���G��� Ѫ^�����wщZ:!o�Hl8pL�����<��'��c�H"����~���6G���L�/�n4ym|v|��@�O���[B�4���ud�\^mJ^�b��1j^��L%�w�C�9���L�h�\��0}f~VTE���@�M7�U��
����Լ�HN=�&����O�Ǐ��l�U9U�]&�vm�t����_\��R�}���Q��F}���z�p�@��K��/n�#^��²�,���K��r�5�VY'`�#7��KF���#�xKw��ۋ�����f�6'� ����ڞ�8-_�U{��F��2EFZ���0���t�?�cݤ3��?A�ƙ�H�y��]P#!z�Ҥ!ӳ��@�LG�"�GT��'�����=2]
�[a@�����vKk3I��U�\����l�S�5�Z���H�޶����~��[�����K}!İ�k� ������d���)D��"W�QR��޶����,�\Ȉ{��h�̦����:�;�v�&i��8�����T~�����[��?��P'n��я�%�w�/:�xYp*j�.(����</��B�L�t���ޟ.��=�^E� z3k��c�����P������eK�K��0폃�ƌ`���n�S	�Ϧ[�z	%宅~�Sf�F�$H�6,���\M�x��������Lc/�*"�룖��9n��COl:���j[�=R\Q��Aq��*� |�?�\{f)0<+\�j\�}�C"�R���z���X3+�"Q9�B$j[�Q}~>,uH} ���؄�7QL#� :e׺�(��>�4Ȕ��7U��Ε�	���;��i�?���D�n���Q�%����T|�;DǨ�T��ԇ�fX�n��p�ބ�(���^�JO�8��H�k`4:u8�R9���>i�ޢ��ڞ9?n�8������[��X�{�)zx��GvC%��O%y����EF�U� �8��xJ��a�l�E�?E�i��G��Z�|o�(�+�@�ۤO��̮��f���u�vB	�9������4OF��I���@<xZ�N3ZY�]7AY�����?@8���MBq}7{\�j�WL¾%�����3��H�?j�{(j��&_8^h��w��#`_�g$��l4
��8ӜP�%Ѭg�sB��mEO���$\��1��f��~(�C�d���w��JMv�<�a��e�p9��y������3	�H�b��WN
�L.{�EYB\���B�pb�.��o]��a�ʤ�����|���Q�&ݪx�������Y���6�����W՟_���뀩�?���'hL�>!��K�D��bs����1�5�>m_%�9���>�'���3;���]�8��Y��i������\0����`wg���,RF�UT�����O^��DW��e*��WO�1�����0QRt8O5��ũP��7`�;aE���,�,�?Hj��gʸņ�tR�<�[��y�(�㋞����W�avj���I�d��}��S?,�qC�\?5�m
P��ؾ�����0|+o�'�^��?�h"�y^�{���������MN������+l����Mv���Tl��6Ŏ��,�,�= '��j+P�ژ�a>'�̧�s�:4_�oG38�mR�#�T��+����uQ���5�w��֯e@���6.`��T����A�{�\�Pʙ� 4���G��\|�H"5�Sǩ��6�\�:��Z�m`�k�'kT*��W�r�dʱ@Q �vw�F���޽���5Sۖ>�Sw��]7�&�����T�E���˃z�����F�6"�Ʈ�җ�	�Gub�?
d��v�ﰍW�]-�{wS�W���5�Tw0��?�& uZ?���P�����=�+�r�6�z�"v���������m��bu%ů��tj�'�(�I{ѳ�V_L�K������<��-�=���9����x��8�l��'���	�DH���Ȼƞ����:a����&�+v+nh�4��kT\��ڷRhX�_�!*�D����(���W��
�ڣ�:K��דzO�e��qm'��
Js�k�$�0�f�Lv��̓ę4-Z@m�s�M��꽷�wҚ�Y��I����ڹtlL3��
|�WG;K�j�w�-�]%$8�[UyT>ɹ�|<:����5�~���%���ʏ�)u��d�_�GJ5���i�$�ŤSLe|.ώZ��v�S*�F��e����E���1���>[z���[�qf*3��:Բ�yA��l^�%���	\���'tɐ>W ��������ȯ* {Bٟ@�7�b|Q�C��La7f �;�����sL�	ߓW�f;��uّ�Ċ��X6��ܰ��%`�\sB�g�X��T��EsA8ҥ�~�?z_�N$��w�Hvj߀	���DF�&�D� -.��CÓ@�Wdy,
�1�����N^%,���:(6�r��H�ݳ=dLo��oё�fUR��3��!]��Z��C�����{PGb��5<�ϾY��&�4]�nm��2�=Ӳ�ZZ�׀dڼ�nItѬ�y�]v�k�H����i������DG�� ]dL�p9�ϵ��N������u�"� L/j�#��c�ѪY���B<���IG�#S���<h8,�Q�l�l�1��i[<���Ra�'�ue��.�Y�Q$�B2�_�ۚ�i� f��A=^�N�Si���C��`��%�{������B�S�<P%N]���,�n�-� ������=t�YUNK��f�db܃����%�[E�:8��l}#Jߗ��'������R���ݵ���%�
��61XG�yz��b�O�7[�� 5!�`u�#����y�Sxd���(���tR��j�WB^)jh�Vv�/Fg��6õ�y3=�>�u�ktt�s�[��e���Tb����'�B�!�*\̂ă��?�׺� ㄗ��Ǉ�H���9���)�Z�`#��7ɴ=���9��W(��Wj՞�|�eb���O�G���oZ}�[�]���V�+jC�B����Ҥ!��)"唦β�9&�q��zU�c�<�����bW�$p�K�Pog�ic�?���;��g�B��mt��K���NL��L'�5Ϥ�Ym''Ț��<7���K��V���C7�����)��`��%^�h�Yj/K�:s��k0�vS��T�l;�*�Z�y��IAmi���3�J&���τ�ݡ�c��o#�Q��_Er��C���7yA���O�O� @LĻ;������*+�}�V�x)�<���e䦔M���{�0��{������ܘ�O�!.K�6&�IS� +�A��~��p+�lA�t�
���k��iث,�z��M&��~�)k�)�~� ќ
t��-��ޅ�MD��A< .MmՐUH}�BzB�v���@�$-[_�=fe2�@#_D����e�(�{�D���@ͮ��A��2:����9FV��TO&/T��X"������k�&r�梺ߣ�uӕ�~�����wI�9��0�;-�&p����B��)��Ó�{�"� ��,=�k,��҈��� �7^��X$%nu�JMcS�e�#p��~ �	Ip� �9���2w{5o���P5���ȫ�J�$t��}u	4�Yg%����9T�ҏA����3�߃��m������?���N$U����3�.�E������6��6B��|G���ô<N�>z�>�4$]Q�P�������@�y�J�5�]��
7���Jә�#���lS��;?&��Vk����8�."a�r��:W�ܬ�*��+s��	�J�ӂ��X���z�@�C�-�e⻰�eN��@����}96����'��8c��j��[1�$JG���7Di�!��tlJ��mR��:`26��A����Q��m]세�Y���*�Lb��̥�	�(|�a���33�C�	k�M=�N��h�[oG1l�A�d���}MV�A\8��G�_������C� ��>f�*^�����xѷj��ä�8�c�txPy�գ����J0t�&܀���������4҉ת;4�|��Zp��a��S�M"��"�4�v�oRl�����?LR¯��Ux+�ѥ�k�����HQS ��!�`��C}�/@������n��A���}����l�a�Aa��Ɩa��	��ݪ&eZ���AZ�TH��������GV��Q�ȼ�=�r��O�9/0Oe3r�t�I&��>�]VX��v����ґ4����;u׼�ɷ0\�t��$�4�PA�D[���hH�By�, �w��H�Ć�&�����0\=�a�*�ZP�T��-�����)�l��%�N�b��h�뢐���PQld����q�p�
&�.L錡��f���PM�Wf@X�pV�i�x��w�rbhMDDXv<;*����R}�$�����(��:���^e]#f�3�|,ޡ��p�h��������Y'�������/�{ȿv�I��'o��?�:�%��Mj����N�EH�v�+`�����El=L��ҬT�2E��UH��fE�Հ��;�٧B��>X�si�������'-�Ur����C����3]�U"�����<����V	��$�Kͭ1�Y��R%-b#�� ��{o��]�_��6�v*̯S�iU}��.�n��I����'b=X����o�D{��]N2��������&]�v�ӛ�z$�F�c��Zs�5%��e.}ܵ~"��'jf1��p]+���a9��5�ߌ�H��`�p��WRJ��ߚP'f�>Ws�A�xF�w����b��tF#9@�a#�+^0�s,�>-���a�#��A!�:�#{�������;����̘.9%й��-48e��T}�_]��h��B���L�NO3�z#�n�uY�C�W��;s�ߴ��V��Fٜ��OKO��S|s��(�x������D��g����5�c	F̀�2_�R��e%:]\L����)�>7�E�%��>���n� 쇱��RZ�u������D�p�I�\L�X"fv��>�F/I���P�T��)�FR4�ʯ�j ^��:�k$oRY��x�_0)�ل`�#Ôݜ�z�>�Xq�q\��z�N�=�kK���d��;�F�ɒ�Ʉ����c�[T����x'��Od��RM���j󆍵�u&���I�
��&(�ʂ����>����/��c%zs^PK�#�6��26{q26�:2�'���>þ3Ͻg���ve9U�تo�L$�M
���I��r�)��\���K7�&4��l�"-}����s����Gu�-�0�췱Ti.�U?��@9���%~��9p~s��`�J����.O�Ո(r�ٹQC���d�w@���������~��)&�u�5��f�y?i�k��Ϙ�SAcG<��:y�Vө &��&~
E��{��̖�􄉨��6�����!R[��ژp����m>�����ܨQ����t���Ӯ�	���Q�Ad�5X� �h��8U6h��=�)0�e��Bz Vw�xbxu��M���0�� Ny���f�{��Q���͊2�FͅICC�}(ٓ�8vjk��w�3}GA�ڱ�������ݚ��xqLo+zs:~�VS1�(�zը�(����jF3�>_V�%�U[b(���S)� f55V���U?@��[��P�mC���C����LǦ���E�����JU9N`޴^��p�5���	����c�������2��g��>.ֲֺd(R�p��㮨�� R�g#�fc�u��RF����vA�x�Y�A��d��>L�2��浥`�7�e>_H�#��1�3�4����7��l�*tk�Ky.慙�����	r�;�J� h�����-� ��
�h�B����7�D�l|����M-�Ak]��h�h�N��bB�����BҸ����c��J�(]�XD-oL������@`	�`=1P�L��&����K��<��� ��o�ޔ�㽖F
B�p%KebI�jy`?�N?��ϴ"�����Ԕ �\,��%�
>�H.oxp�|������&�#ߪ�����p��4�[P��S9�U:�1��� �并��Aj�Z��C�aWP�����7�
0}��/�=��=�h��8��k�u�n��8��C��V��X9Ex�E��=pZ�},\k�-�1r��U�������gHE]f�2�d7
��Ͳkc�AKܻ��Y���czL��	ro�7+3������HS����a����"t��>#���D������GӘ ���lp���f����3��,���C��_�qd�/�=o'(�̣��C��d���itR4R��0v�ԇ � T��J,������l�Լ:�敊�P\(٥�z��G�15E{�u��|�����$����QzF��܊��6V�v�3�BJ0��+A�G~{��<�̀���rC�8�b��J����� ��W쨛7"c��Y�K����]�;O3� ިG[�<��a3r�ð]r���c��Fr�]ʛ�(���	t��O苋 Si�7"Ï`��PrM���Fa�o�u�,�����ô1h�?��l/�k0������ҶvF� q���a��(b���(|��Cł*9lk����88��g`�A�н��g��|�h.7�6g$ӱZpN�)������!�7���?5��OKR�B{�a6g֌�c&2����Ru=*E�3�,E"M6�=㬸��`RA�ǁi��"~��zM�8*��%|I��uy�hԃN��u;��J>|�w�i�u�k�lJ�'�b?�ɿPR�v�x'�f�
����{OU��ǏC��8�yҌ��s�b	�W���r��eEW4G��<Q����.Cu��i�cv��K3���"���M�^���C�`n�K��� ��(�|4�q�.p#��bcZ��7#�P��{������a�&�*.VP�øF�c$����@�t��T�V��i],�6HuW�S)rʪ��y��3�e��@{j?� ފ����j��<W�@B�-;~X4^�e�F.��s�y|E�m:&�n��^٣r��<\����瀭�Jo{%��21�4�N/�M�*Mh!���܆�u��`/�=��O�f�?�eV���)�am~7������J��_��i0k�W��/n�/>~���'��␣�W7�u�"��7�X/�g���<�����8WHG:!���U�0�����pF�݊64��d,b��&���3�iuSM�%�:K`k�% ��-�t�1��$�I�z����;��$�4;?F\L��+��f�ZRp���"�=�qc-{Q�a�JL�M�~����y$.	�9U�$L�Zl=��e���R����!9��y_�Ն�d�}d����̻wv�j����	���Ⰸ��9�M���N�_�3?��s�G�06��b��}�O����ƀ�0��9�et�X��YD�W=(���4@<���G#�����K� 8/E :/�YV�5��Y�.�@������`vº�{�<&��{3�c�ld�؄�Fv�$b���z���v�Y�V�~�ny]�������ժ��_|t�ܿ�c�����Fh��}��0tG��qO]���%¸���b7<����L��O�	Ҍ ��OsH��|jK�b>E��˙<v���b��/q.�O�9ſ��C���2Cg�8��#KvY	%H��~�;n�b�����Ȧ�˸�y�FD%�#l�Ftw�k�m����J���(�p�\}G G�W��X?�>�/��ZY8rL��&�q�E9�t���#L����n�`0܉FJ�n��*��M{W+qSK/����+G��z�]�
y-�)X�Bm4+�z~*����L��C���P���B0�u���
u�(����)����V�z;߲ O	���	䒚����[-����&�쨪yb���XsU%����k��C$����
�j�H����hHʏ��;p�:K*o$~���]^j��W��M\����dr:������o���d
*'Rj��Y�$ob�oբ�)|�Ymo�H���&=6�`n塲Ȇ:�2M�h��ձaV��������M����Ω��v�s����f���Uj�⿅�l�(H�]���v/���h%	���h���M;��똈S���k��)�^�#���=G�-h��y۔ b�zJ;���%�q[R~���I�_��x*w��^
�N+�S�R~V8B9��;�%���_��I3ģ箁��&�A�Tr���َ1/��8+���yujp)=w�w��A���!�J��9�e7�ٳ�W3'�f~@q�#�:�v�?��!�Ţ��
)F8\�NM(��f�)������o���b����I�8��U�er��Yog�è�3��_b�&la��gK&���4��-��8�*�ȩ�)����x�p���cf{d���3��۪_I@��'��[sO�%M�z�ȀB�H��K�0'��W"��k~��^��@]�S�$H*k���n���`��׶����/�����v��+�f#���<��=.�T���K��t��g��:��� 	�/�ڧ�$����-�ƧL.�,2KeU\��|βn�bL�U墭���0�Y��M���Z�K-�>� �H���A��V�!�{㈡� y�7�s�vm!&��b����TsQ���1�U�X^��(笔��>������l�S���a��y����������U'e2(ܽ��Y�Һr��oI&0�E�г�K�YIs�xu�w�yW3	3����	48���̴�b>��3��6���L� �w��B�w���%FJqV�\�!>®J���R<�J�$��g�]�m�Ie�ewttv'����`�O����:���i��4]w1�GId�{ͣ���Q���F��Ϥ�*���l��'�7�:�ߤ1�
5{xјs�OLH��s����l�]��/�]�ԅ^���,9][�|2-[����,H�F�C]U��l�B��L��I1����E��>���wi5c����a����q�� �Rߓ��2�N�v<�D��1�UvOF���`OANU#*�ҽA���?:[�'��Ai<��mx�̾��𸹼��g!=�F�OW�{�\V�v��Ӭ��A����`���Z�7,6�t�=G��Rt����/[�)�r�a�L�D\�E���5�2<�Yʁ�ysn�Ӓ��p�l����Cu�K��!^�݃��:w46�2����=cݵ�zQ+�4mn]E��2z݋�r�p�}��,�h��ڦg���;��;n"����u�[ǨW��G��&M��Q��;c��U���c��[z��Lڲo8_E�|eRJi)�!rW��%]��v���\� �)0�ξ?�����#�vD�%��M�Z]^؎+�^s�E"�֑�J��@%��6[�b����ط���J�T|8�ı0��A;��zhX�+�N��=|��]G-�Rˇυ�V3��&glr�r�d|��s#�u��)
B��g��U �X�z9b�2oB+������y��͕��i�0���>�I�۽���⍁b�I�`G�6c`�0�����C�q����k�w(k��`Q沿S�EBC=�ql~˧�����ލ�ç]`�{��
n�m�6��/Y�V�Ou��c���re�f�1d����w�EI)å�h�J�J�1ZtJ��G7��"�)7i��S�dh^�E�O�~�,��M�	��nȔ3�`�*Rw�%�Y���� ��U��ʌ;GM��]�����=dش��2�����/�Q'z�m8�g���ۢЪ�m��^�$��#Թ� �r���C�=J�'�ÎNp�2$]��3<��I��_�3&�#�>��#�i2�]�a�ZN����-���,֓ s�n�g]s8w����X�(�aU=�Gj�0�C�U̬q�˰|j��z��>É�G��{�x��O��-?T�CL-���Ɏ����I���~�HBҽ�BJAcf��3���t�m~��u�]�#��IJ``o�HB�,��Jgutr`G�mp<�@��� �V�@H�
s�MB�+y�f�ا�ٱ�%H��N��Ϸ��S��y�	��n�����O
�s��L���u�4�����|?n��x��6 ���z��r3�o��E��uE���5�@�ś	��@�,�EX����ɮ��kds�9�M\�� �n���A�N�������N!�� �1A�������K���^܋��A�8 =�-V��JX9 7mKBjw w�ۢ�f|wA3�Nm�D吏�b���Y��/���ѕ��a�(SG�y�g�y�.%�08rw,�y�{��o��0�sŻ����b�~V����h�n�j6���o�0�N8<��W[��S-�3��&2�?(fA�C�������>�g6�J㩏J��5�Q��{W< B�O� G8@R���uKF7E�߳�l�(�`�Kuǩ6 ��X`�*���4���3�ߔ�I���^�?�����8(]��Ě��m�mzB�Σ�u�Z�4�kʈ�@���b�p�V�ܠ�_�Vb[,���b�`q�ؘ��Ћ*���;�9���i9�����
	� ��j��pp����tp\�udu�T4u% �9�8�	�j�W5۠i�Dy�Φ�d��4�aM"�ո)3�躎�(�@��y</6������g����<Ba�s� ���U|��F�ϙ���ҭ��'8.�a��XSS�9���������	�Ym��"r�g�p{��tq_�W���Lȷ�JR]�+��R�8W�~~���#��x��p��B��%����c�[j�o
��	�ui ��Db@_�[B�l���rh��{LH�"�F�]L9��Q�ƌx����:��Gt�m�9&-��+0�Z񻌉A�U���l� ��F��q���b����ڄ�(��!��.�1�u�����o��e���`�� ��˚ J�.��Z�mҭS�����p̚9��D1�0���ފ́џ-�@3n�oG���7bK�Q��y8��I;�]�����k]%F�g�g�`�BGpX� ����r�	|~�j�7n�XlO�����nP�*
�U�DD��GpQ�X �+Zk�ɨu�4%uT�D;���2� ����<DW���JT2���E�e��,����8.��J-�o��o[f��_K�"� /�� �+��T;�KU8>CY�G||q��h9 V��@��T�e�ٝ��1�>Ģ�N�� ��sҦ�;��uA�2^-]�����Ь4��<B̌�~)j~�ߊ5-��%h�<�x?s�W�`��8
z�@����؍��`d������k�VK;࣫�׻�_��,`s��mRl��giX�E��e.&A�ڈ�`~�*���� ��~�p�W���A��`�\�F�t:Z~��-*H�$����{�}`8%J�&�-]��9�ӻE�
�P#�93�Ape�%��.F\`�X���C/ak�rF>я�^��IM�_�v���ϡ�fs�`������FD���#BΠֲ w�a�@�VM��s�G�*_M��DT��'�B[�|<�q|����ce7�{���Ko���ʺ��C+s����̼o�����Y���m��?谺˟ԋ_>3��h܁�78�O�#1��%�q5�,�g�'�M���JQ��=������9���;Kq<���-f"ε-sef)��^rf�B77\���3H�:p��3k�ʔ���4�f~Z�Ǻ�Y�,xx7�-���+cc�䥶�7:h�K��|��e�aQZ�ۘ�R/���nY3�����ا�����9�+��nZޮ�n�q_�E����	;'���;n_I �R9�S��=OGr�����F�R���>� CMA�!�h�����ZJV�%&���%�����5��	h��p>����@'P�T1���B�W�.�c�8��9������Ng�?��`�	��*�\=���O��R^+�?�is9�488�9G*������c�sk�d��G��Nv@R�'½���^�OU��H��i�����$�/��~����c'j�le�6�Ќ٥�_Ǡ�XK�s���"TD=Z0�z!�yCH1���r��h�g�y>3}.�rx�y
��L1~����@�ˠ��Q�	��nՔc8g+3o u��+V���?��E���X���Q���WF9ڇdnx �e楏���Y���4e{��	�2��ƪ�p�kI�ȳc6�y��s����Qh�|��㲫����^���f3dԚO;ͅ�v%�H�8�?,�v�k���ҷ�N���Mf�:�O)Q�_�R�Իz�G�Mc�C������4�ۥ.4PH�\͊Ʉh�yU�~�R�0�2�\���
&�H�N~d�H.�{v��X�.آ���pd��,pb��'{cO��bTv�@�r\�y������/�B:7{���6�p�����D�O����m^U�)���l E?�_C}*޾p ������,�ɕ������Ș�r�z�ڛ�E|62R.�u�$?�2.�%y�M��_���-���� PC^�Q��Y7O����wڎ\�z`e�_=X�~+��A��\jZ6?$�?��j-�!��2��Y�Otͫ<�q��/�bE��,&`��2����ہ�����)zc�V����	qf_k�~P%F�--_��EA1�V����������G�̲�r���ةV�=]��o�j�;�E`�\�nT�i��������PZ��eO�+�Ԋ�@��wo�b�
-�^��;�+��Os(9�$�	A$�0��tTA6�?rF��n\������r�=��s_�����t�����~�cC�c�oN�q	�\��?���D�����4�Ml��
w�?��("�Y�;L�y:���Y����H��[�9{Ŧs�*��e�0�%�h?p��<MYgD#�(CD��Ƙ�<��'���<��8��t\�4
�Y��ZMU�C�z�x�U�� �w<zI��{�$���F�6ʏ�P�/\�=�"�l&j�^�4��/-U���Գu�i��!{�_}H���+��C����WR(�M�e�*Ɵ�x��d��L���60O�h�gbq����p����d `H�5ކ��� 8v�n�-�����ڞ��醂Q���ϝ�;�LN�
0���<⣽4��{@���<����Vd��M���נ.v�B�������E'� ��v���t������'`|2u���ٔE9i}юa���!*�D@;�t��(PS�yؠP�kԉ$���R�aC�~�.ia�r0z+�Kw7� �6kSNp�
��V��5������gE�,�ޱ���3L���@�R��o?�S�)����#fߛG{$Y�E������;ÃI��l�V��%��1#�/���#���(�<c�o�\�k�:��6��&h�yjr�}N׽��WW�VF�V��LƖ7��>��6�W�ߨ�kK�ޭ(����`3u.u`6I�^�97ܔ����n��}=�8I�i�k�S�yV>����{��3:�	�Ym�ѵ�I�4Ǎ��r�X l�E��¡�:W��Pv���}2����3��e�J�@@�6�U���	�@8`N�.��u�����Z���Q�"3�c�8To�E%_��;[-�Sf7�T�G��v��@�/qrQ��1��>��=ܶ\b@8%Rα��镼�{�M(�b���Z F�����ĤA�����PX${+hə)*�%�����n���^�E'^�#�MGC9�F��ge�򛏴�`� 7���j �w���/��z0�:d�u��i.(n�C�?9�Y�"�B�V1���F��� ��,��Gh�E�����#���P0�Y+���E�����j��X ��*�LWu�b��NuG�65�5l��S^q��X[J��*����v��:K�d�9��(�	��fM�&�,I.��iw+�0"Oӗ��وӬ�¹�~t{ךx���r;�r�w�F�G��a�@��,�Zɋ�9�2�B��w)7��H�c �Zél\k#��=�c�/�U�pљ��yl�/Sća&��U��z ��$I�	�>����WnWM#�~`���A���|!�_�v���%�6	�B�Wq6�F��Lt{�~٠$uk�X�@��?ߥ�t�����:��dUGJ��Dg�jD����L>?5�"]
ał��������'��F]+���	г�4;7�}���Q �3L����f2xۃ�C@J/�T8�ob�-u^d���>y��m>��&J4����yj�#�Ԅ8�ζ�V{�0��X����G2��@�:�<�>^�ZYͬ�
�]�w��T�6�9���"x-�"��i�n�*�B��?6��,n���6��;���̧��[��(��.�q�d�~y�?$0q!:6@%r>;>w�$tr�Y1��A�L���i�:Ǎ�Y�SkB.��Q��s7PQiT�g@�/��	?��h��V�ۅnE Ai�	Y�����.OE˚G�i��D��W�� 7�J�Y:�]��o^N�s~K��fPA'e���D-�����w�b<�[�۰����M^"�M�:�=�Q�����C͓�6I��(.7����׋B%���|>�cα]=��)�I��(��Sh"��c����'[���GT��?=�RE���q��1�g�e�l�wBjQj��� o�FX ����v��P>���ֺ�/[H���?��������Ⱦ�z��윌�ۢ�P�Hrz���Æ�I�j�H��%MO1�`Iȟ7�=�:`����|���ջ�jf�������V�A��U<�	mo��qMؓ"i$�|�@�Ҫ��,�Uf,?��˃�^�6�+�!NQ�"0w�$��4�F~X�����V!솹_��}/7�����l����ŭ`���Z�Ǩ�{�5G�Ι9�@a��0;V�Y<��j$A3�LX���h���C$�kV���>BZ� �ͼ��T�t 8�F�DD��<�_�Ϝ�۩�T�ë�A3�*��t�]���C�kَG��%��>�I0(�*�o��E�㒝�����1C��]�w�ߖG�+�ӱj����רiymh]�;cq�^k�B*jK���{B��"�m鎧�{�"���
�S�ٙ �!$�,�A�^��[]T���`f@N����M�"Yc3�o�`~@�B��#��TXs#�X(O5雨����R>~�S1'=<yV홋�.u�$�0���?�s�`�^��l��"��5�h�3SOh��%��E*��Q��r�r�A��ݕH�r`��O��p�e!�&�a�D�� 1��t�&c�k�%#�S�V���kkd��n��AH�u�9�����_�D�u�p�ﵵ�폕����&B}>]qs�Ũ��n6�=�a�J�����j���� ;�#����餬洹���<e|#rI�?lLY�3����K���U�
1ȍ4��b`��ÈҋH��vu�w�C1/�|�����%�WC/hL����i�"P$R3,`8E����HoU��C�N�������̥(oͯ�r�\	������rpW6���׏������J Nu�\�����d��LIDʴbT�	�˝p
>J�P�c�����<����4ɘ��|�֤v�#�'������kah�	�����S��r����FS�vָ~���|�����T2�����~�ޖ�qaG���e��d��l>��Q�%��{N}e��q��l_N�S��	Fu@-?Iv(Bֳ��VJ�ju����U_�-r| �6\����#-՗ͭ��R��R��wCg�����ժ\���L'g����'��������s�	5����ɂe��sv��T��8jҩ�i��8�K6���� �d���v<"�p\�}�Cr���8�
@S�.��ɕ��ޏ�$w]���q���}2��t�o�Q<?fG���.{�1c�d#Hp��! ~����1���f�{�)Q�Gx(0�O�!h�����j�[�/K��h!�B�N�K�(v0x��y�> ����͞*Ѡ͈���`���þe��)����n.<РW��1�%#� G�����C	b���"	V�MS�%���#/T���++�ߊ�G�����k���w=[�Ւמ��6/C�ST�R<�����O~�ݏ��Ab͘�+@����� UW�e�Yxا����ElA�L<V`��ڠ9�(�"���D;��Ȫ��:�|�m��(�f%�p>�'\~O)K�Y(	����Y
�X!C�Zn�22�^JY�*h]{%�|�=5&��qdB�'�Qy	z���a��.��9H�@p�������xj���4.��<i��`�O�<�,7�L��I�"H�)��E��/ڦ���ti�/t�Z�J�t�T3���J$A�|j1��d�!��5�m%�nj/�j]��IOq�!66�vb[��ΐ�����3vI@P����M�ȓ����q��Fm�c,ؗ(��'_� <�nhŰ�lH�+r�N�0����#��G��5��p��<B�G���YO�y߂�~��x��0�|���^r�Ή��i$#S�x�
���P�(�K*�]1�.	���3��c<�D��B�N Ԧ�W7��A[�"�#,}_ˁa�U�}��n�CJ���@��/-妶�T�!�/�&�Ea�9�v�Úe���i"�I�B�S�Ӓt9��n��N,?���.a�tF���mn�K@X��z��z	�p�@�+{����!�H�@fG��y���
B����Dx�u��	^�m���(f^��y=���4.����l�oq$0��5�W9�&� �DY��H�;�#�f��K�v�#�'Y>��K��P*��9����Z���^�� П�a-{�����rh}d�C�lO�߿�сW3~k}��3ܭ !M�%j�L_΅���C�{�4�ÔQ-��-�vuu83�)�)�^�#�$��I@��z<�Y7�Y���F�P�ha�Pr�
���m5�.Br[�46�y�������D��y|���+>�gRӜt;����/�~ j�'��ȧ��1��%���&����D��hN��Ѩ_i"���.�a��B�(��4���&��v��w�d�װ 䶀�~��AQ�F��NDc�v��R�q�d�z�cAX�2~@�/���{oF�l_�ؠ�rN�U>�;ˋ1[յ�AOZ��o��#�½��,��_5�D�[."V�qeȤ�t��I�@��G��S�g�'��:������ ��UC&��<�hk$!	�s�'b>dT�����LG�@������t��Br$���W� �H:e��{�SU�wV`LNt�>7�	�J�U"F��箧H|#Y�����,]��x��~��esUuM�w'('�Ƞ���5R��3#��$s��
dEV9� Q�jӝהE*�-�F��U�U��4��ή�9O��|ާnv���	��ko�9����ُJN)�̊(�Q4C���~�5�|��5)��1̉���Ɇ�Hf�mNq8vS�������@���_Qh/`M���!�8���>Wփ+ÿ酌{W�n��c�Eo�ӂÓ��S���R�S��j	��[e�,!w��3�e�r[t]��L������ޭ�=^/SPӮi�mh��@{�HL� �Ze���r!�(�Ud�0G�i9����5r��ȰR&H�,�$�,��߃���k�lܓr_e��<�m�STH�Jđ�)b"�~m����A5j��/dȺo$�[/a�	7���`�KT-�Pc�ǐQ��s?�p�P��sݯkC<`/�4)jN`�	n���*�緪Od�L�EW\[����pL$����}��
Y��'7)��)U��ǫ�O�؏����	P6r k���T�?U���ky�+���:�@��[�eJ�������!tW?k�%>P��K��,`-E"S%`�u
:rՇ�q<��h:�chZ�/+H�먮1��1��E�P#6;�x[kS���|����mN�Py��>|=�bE����X	��bb����a`���}��M	��k�E7���,�%�֡��b�V�PA�|����K��D�K{@��ݽ������.Q\���L������rtf@C� t��N͑�j�܆��p�	L��cƂG�S"��9 ����O����)�E���U����Ы�+ғ����ڣ�8Y�\����Q��卓�x�H-��]`㢾��LcsQ^�ᰮ>cL�@�n(--=_;a6�R3A|��`��R3�!�l�����jeE`��C
11��4(q��T�bgw�O��8��d��eI%�si45S�X�f�M� )f���]�Rq�}p*�p;�c)�Ģ:���w�݃1�����с�DX�Sn= <��.�ft�f��΅�plw(�t'�����\p�׉�[�>.�Ԭ�m��cW�����ښ�2Cx�'��V&tH�C	4�a�2�?��@��@띢�3t�a;z�D-]!��*�d�|�H��Y�u(UG�HΏ���@�器[��Y�8=��B�$p �s8�(�sE�&=Ҥ���Bn�6��<4�9�nX��Epu�B��	�!~�=���JM�Y�r`Dla�FV�Nd�c	��q��(�뫯�ι�A$�
Ϥ��g�:�~���	$��	����e�%� 2�Δ�Φ�c�N��N1�v���zw �^�����=��w����܆��4��v�i�b��Y�β�~���T���_N �y�'V��QG��Ķ0��_�sz���`*A���)-�@�v�;�/*ONX���~z;��U��y9h�t��K|��bzu���?Z�֙8���Y'�m�����?��3'���콆��kA[n,k�fr�ú�2�!��WI����<�+�#wA�gwS�v�X�psՒ�5X�Z��&H��������<O�hcB���2�T��+ �<!�f�4[ �#a�$D���PB���n��Q�upώ�`�Yl��)�9�)�I��2��b�?�M�n:@j��߀w�W1�~�m63κJ&oj��v�Q�4s�N��V���mu�&�5h���8�6O�W�2�����DSd\<b���/�����Qt�T�<%�]�Y���!��t��W@͠y�Y��YѾ�J���pF7�P�On��}L�Z�Q�&�g�h�(�_~�-���w�d���X��x�8�cL�2�.�d&u�<�2������ ߽�z����!��|B��`j�+��mו6�MXg�`���|Q��R�7�t�oh��(���S�I���	�X��w7�*���o���0F^��^�"15�$BZHՉ��,�I]��g�&mF����z-�Z��/Ua�,�t#�Y��w�v�7�Nokջx���8��{��	r9Ts�n�Z���A�	�Y��6zVXH�z0���Gl����E�K~�hQj�����5�9ǿTt��HA�C��ѰS�Ez-c(5
�+L��&��u�S�g���"Rw�}p0%��8܍~�4$:�!�#�	��%�0y�6?���m���L���"��%6�`�u���@�������%:��:fm��@��=�)�`_�`�Ĩ���'���h;l�EpT>��C0 ����y��ʳme��ę�OR�sNR��Ս����
��c��A�G�:��9#�t}�Z�^�-Ϗ��d���a��%]D祇�6�Ŧ\��$��@���
N`�N�����ןwN�7�^��t��!n�ʥPb'HUO%�}*A�QD�i�9�r���p�L�V��/���`��@��`������>�����1Hf���S4���4�4�HwF�Cyy��v�������K5J�u%�����_�(j��ei�	���^�6���Zh?-���A`p����'�&u=�>�0�����L��a��8���x��w���Dk�x�ԩ�]�3�7����%B���w��c��Z�����T�p 6��v�>���9�f�T=NO�0�~���4����'b��Y����,�Os�R�����$����r<��'��ťts���p�~N���Y��B�y��*���ݡ{F�m���V�@r:��$8� A��U;(�(��t�c/���_�����S�����mI�V!���e����r*mq��5�S!�����R��۟G"\M�'1�[�Ρ�e΀TUN�zak�s�sӽ�-w]NtĞ"˺��{>#i��.�W4�D���¼J�;��������:y4?vz�幩'�hE�Q%L�B>���*o�3�!S��ׂ�U��}�O���,�B��Ù[���T2�W�ㅹ����!!\(=?G~>g(>Ft>���%d�����=\��rF)$=]H����3�"3�fӄ���[O��\E���]I���.Y��U��֜����-c05$�Z��.u��+��/��,��nS��-�4������엝���M�0g�sj��w�*`�F�(f�j�T�_ݳS��=J��Q!��+k�_����3n �� ���a�y�D�	�Wq���w7�j�d�r�S��x���(�u"��y��Gi�Qi����pt˳�^q*/�W��J��1{��>D�HS�6�F,�N���N�!Z���,�P��g�"�˗� O17�"�C�O��c�9�o���7�a�V�Jj���N��-m��ڞ�!Bo�q�B�Dn�:1ޝ!M������7�IIReb�ʊ�5ף��^̱Sf�0�QO��^TN�t���������\��2�
jΏ?; /Ռ ½�x�:�Hy ����y��Kh�5�g��nI�l�C�9M~E��_爨l�bebd[2���ŗ{���X������y��)U�W�����݃�����CC�e�zк��)M�<�l�M�5�V�!>L"!Y�'-��5oqs��^im�W��l�=B�p�6QD�`竔��[<C���{�[�ƥv�?$X��O��Cgfa!e.(?����#�$���fv�t�3�-����녨r�Zq�!�BY3��7����H��1U]<&�L*2���Z ��.��<���J�3>�F�d ��z>��U���m(�E��{�Ge�!�#l�w�g9�M�N�U5kt��yQ� ĠP�$XȘ���A�E��K�-��<G��J�Ӧ�U�.
Q:{&� �wfH�%�N�Vt��{�J�|�&�n]��'g�b���W�*��gҼO�K�)�!9m��������Ɏ��i�����}q����h�`�ّp]4��K#iV�3�Ө.
��hYK��Gw.�՜ ��CҤ�O|�G��!���p�F<�Z
��!������ݶA��(	P,U�p��H�i��4���Ѡ�7��b�u@e?�^��ܓ,�Ge(RO\�7�	~��P���g'3C�ǚX����M:����� � �a�ta��x�M<�k�8�g��ok���Z��|��y=?� �\y^.uG�G0C��*wZ%4�rk��A?vz+]��y�xv�dk�Z�C[�+�?�*��7�hW:#K��z���|t՞�^a��ŰƜV>��Vs�	䤡>Z�KF*W��xjC���4ݏ�@��,(7`�Z��Q�������G���'����.��V���I�F�&��/?�^.T�קxl���B����*Ez��"����`���6F��s�N�{��j~$�>ϋRh�سD���i׌�V�05F1��b+�3E�Fp,E���J�SIX?ý��� �~�3j3�����:E�a�ͽLT/�桀���Tb�`���&z��f�bO�&/m����bv���8��O��-�u��5��+b��VQ.��V4�5hy~|�c&�!�������3%�cl��+O%Bc4�H�h,׏|�����}Ю����7Y�!$�Xpp���m��MIN;����#{Z�a�j�LŇ�s���f���p��ٶH���dy��^;S��AN��i*�W���U�2n�zUVP�d�&���j�(;���k�
2|h�8�S�m�h�|k��D���])0�u���wN`��
%R�g��{zސ_�����KR������� �)����2/	
B��|�"0��p[6�7�j�^���5�(.}�J�U�B�~�����E��9L������D�f�Th$�榸�F����T�R%T[@��/"��X�u�۪k.(��gF��>!]e�ّ(\�B��b�c��E��̸��N0�����y�P~��e�Z��{�l*��o�^4~����T�3����k�wL�������gLi�/�\���	E��1��R,i���iFP}�uP�
;H����q��7���I��3���7NMe���B�%��4��$��j��J�b��FO�o90*O�9���`��ƈ�
�W~3����k��	r,'��L]��X��k�J�_	���.��Y�~�P��G�e�7#r�E|�s���޶׳?��V_�#s����s"�|��1�S�'�w��I�ҫ��R�*b�=k�V�͑L�!̖�����e��.�
�=����T����:�y�Q���Nly喎C���ͥچ��9x� ��m����搿��c F�!����E)�g��Ҭ��À�xE�r�g_�/$���0!m2��j�o���m�	v�>�u�͡ %���;�Ů
�]!���"�a�$G�N"�=�	��-����{:��2��@_[��#A��i�'_2	�P�m�`�����tG�[��4�B�阇�}�PO?ƍ՝�<ްD�	:%��rq"Q@����\��̟w�f�6˂6�$���W�N�vy��|� rX�#�ϟ�1~V�G�C�ǳѨ�4U�ԓ�?������T�æRA�����I.����ʩ���yX�=��,|��]V�6/H���?y	��R�!@V�*0�u�dH�f�{g:w�����Z�����v�VGb��X%�b�(v�5x�_��� (�x(?�Լ�t�������'Qo�D���Q�xG@���X�
P�� 3��_u/�P:ř<�b�%tQ��
��Oɔ���:(��CɐZM��&)�"6(ۑ�l�SlN���n����|-�FYEvӟ�|N�V���[�1|�:��MZ��!S�3h����п���%[lK��xF��v���8R,���`:��4�$]k�í`��C+�rV)Lޙi�
��g��-@D����������	��$�\������ȷ�O_����,]縃��I""3�%�u=���}$;�OHK�JA�|�!R����V�/R�e6��� ��ug�=��}��%��R�*�X��7�bZ�ҁ�T�6��2�Kw��m+������A�&�'Y*�:�ۓ?���^�6S�6�&궳n�+�_�+�sғV����;��ߎ̿�#o�*�(�м�LC�O�k0nl*��vՇG@H�區&�bul|�χ��}�d�s	����Z ��Jx�O(Q�KD�"~�E�܍zH�Q+ [���;FOōy�4E\������QNJ�#"�e�B+ql�rԲ
RgĠ�MAH�C��s�p����+���'�L�{1�+tZ�$��"(W�9"u�^�6�z~��綋�G�GF���}�v�9.��8n#�Lb	����%Hi�ݲ�S�� zc�`g��@��߅t������%�]��[���5v�����:�r5������ע%��= �J�h��w��m"�y&�]$ї�����m8��@���6���Ԡ��|��5�=��`�y����7=��tn���QN�&��k+���-��T!_F�Rjd�d�'��A(Xo��ƈ�ۗ�BxD�(0�Ĉ��4�p��%Q�G�.�9*ŁI���'j�P!UU�hX� &tQ��CP��������u>4�����@\�hmL��j��m���N�a&���_��ʹӐ{�]~�B�ЬEڥ�e L6e�Ր�ո?���-�>|)4%gD'+�<�6^1�4�3���5�׵ջXs|'Q ���z�
��
�>�GJ�QL���H�4��U5�??)NĻ��ی��Z�g�H�ԝ���iڰ�*��_r�>�O�@+"�(��e1���	�cW]��Pg��$2"�[�m�a�K)�I��.��4&�ݵ�ѱ���6�""�J���}:�g��q�_�g?��u�~M2��	��o8���=��쐷k���yB��2��X`�lƂ`��wS����V٤عi�@�Y e�a'��oN�U�V7.Ϥ��Rf�;,�gܯ3� g=�_9i㳄��ZT�/v���?º�7�
YI^����3�}xj[��p�*�f��e.<] +�ⱦ�|��)���61i��r���&<@���(���oXO�=uR��/�G��{-�l[x���eJ]3�P�}��ƽb�Y@1>�W��v�歭)PH��ƲWഒ,|y+0D���8I��q`���$e�IC���ٖ'g� ��3����S���
���'d��w>&�<�ꝡ���7���k�?�,7	����E߽L�=��{F!���x� V>�{k:L G�S�\3���	��4��]�!$�4	R��?�%*��ɡۇ�����?-W�(�������[U��+,KjG#Ѱ�΢b�'kc~��T��Vd.I���T��M7h�^��Qm����A�:��a���ܐ���bDM����(�;��	�2ݖxcc��.����C2�m)�}�����K�<\$�V�9�H+3�:����c^Z+��π)q�S��ǃ������f�0��~l]�7p��#�2�*��Ix��:ot���|�M.8p��o�X���/��~l&[R���X&*K�#��Y���S����T&tp���vh�5l$wDm�:m��s����0�{Um]��!�$ТSƙ����8��ɣM��=�e�?��ݔ( ��z�3�g7���O2C_�:�ϙ/�B+t��ډ��qB�eP�,��N}Z���.���%�	/�(�U�U�L1$�k�u}�y��dn3G�I�㧴%������u�5"�����u��R!�?�u�4Bl/����:Q;�j"-c1���!�����*�;�d�o�q4e���<ٱY�y�Z���&����D�ݼ6=W'GJ5v�ꨈ✰�FfnN��Ҁ���B�s���W-`C�֓F�~XO��YZeO ��&���6o��l7!� ����銟�P�Y����:M���t����2��mL��^@N)���#����+�b���#�T��ct?�~A��` ���m*|�Ǆ�&cdNիQ�Q�Q���{��t�SЊ��\��!bw=�k\4k���s�v�߂Jr$�?\|CnW��y�u�4���2젛�H�i�B\�"ia�h���2�z������	]\I6�"��j`=+��k+����(��5����F��O������R�1� �(
�'ӧ(��^�?K-i'�Ä��	��Uz�����{x�둒��T���ogJ�&�^�Hɮ�گ>��0o���_8���C ��BW�-�0���8����^��7=Q=��sk0�~x7�h�2K�$��)h	g鱲[���>
�af�
`�C���:����������q# �3 Z�@G�Bd�������6�O;��}�(#|�W\���^�s��U3�mL�8�f�<K�lE�h6�2�2��Z�ks�s({C�:d�3�ď���m��,n���r;h�R����)���˶��M��ŠAic�p��h΁R;߈��y =�-o$�k�g�$����*ƴ?��}���n��'����� >3Q��X�[Й,2%�-�����fK��K6�@>��4[�2D��28����?;�K�c�*��{������M8��e��S�j�(K�y۔��r�?��O\NS���[��՞E2N��'�"q%n���5+�12CF�x�4b@u��y�aV颎U*\�!KP2Bk"���a��s��~�<>Ұ����~�_%�q����.ߞ_��8�~|ʎ~�ݔ�x���&�欞�/�O�$��ƋDN� �H��+I}�(��a��ŠzY�-��S�!�w��(4|���vaa�4(����$�2�������C\-|�h3�\���E��(i�֙��mq=zPּ�*��_gS�d�P�4�H����������X:-K���{v�,1L}4��66k���ɹ�{�Rc���WNn�z�XZP�&%�.38�xV�}}���rL���ی���-�g�j�c^���m��1q49�mv�O�w�k�u7�M��c��Z�W�@�)p�^!��������) w�U5|/�7����ijRq�v#p?Q,���9����W7���M.20�����1<Z�XB ?ά"*�%V���1	� ���s;�`��M�o)82�pG�oNYk{��kv6<աZ��:��|���O��Nڴ�u�V���ʀG=G���U���2}u�&�e�v��#H�X�UGt�3�S.K���HR�(j�Q&,� O$L�8sҀ{:.&hx���A-�L�{�<3QpI�
�T��N"��v���D��{�w���.*���'�g����iFht0����T�6��@��W��@�NP��'k�ߧ�,��uW'.D�a�:�鹖H�s�I{��̦��5�gEȇ���2�B`Z|6!�T�g��{�z���~K1���҇;}x��'�lJF��HB�oA����� ���YW�W��(�>� �E��j��~|� �0�\���<%��+<�t���kX��>�w9ɦ�y;,wX:@9�L=�'I�q�\=eM$ ��͵��[��0).+�%�x���ʊ>u����I扯� Q(	�ş�c��hhM���B0+Y����%?��Z���lZ=�1* s��g F6����ڃ>a��]�?�����G����U��lNe!�������p�����"y\V:{����
r=����8x2A��;yQ[1���k�+�梶�\�f�+�a�}�M~͗=�O������l�u��ߘ��:����Fr&�0�b8>Ȑ.k���:���c����o=�3�q�oF �?832tpS�)7����$4����/���+�f�Z@�����I��t/r�Z1慢��ӹIvM����}���c�N��F'N��7�T(Ux^m�4m,\��&�*N���U���:��,�:0�	L�6��p������b�u�~ϭ�:���&9�����b�'���+Jd��jy��<�$I��`�8Ɍ��/"O��w"�S8����p2��?��Bp-�")s�Ok�3�~o�U]BS���ړ1��8�R�a��L�$^b��F�r.�f
Gb�P�7��7;��}��yqf�4�Ȟ�_:Q9]L�1�&P�`�nŪ��[n�S��Q���Ѯl� z��}��]���[��v+˪`b���'L32Ǳ��As8Cڀ�M�Q�J��`Ԙ�e'R³ F�b����׬;J�~��_��g����1�����?��
v3_�\A�SH҃�D���P��6��fA��_b��3ZXxZ�h���F�QJ�"����$�+���Ń2�)���/"�O�}#g�nr�;��H�߱�sF ~�����lo�
��t'���aO�k��;�|��r콯����~���j�S�!������c�vҢX�ߠ��x�#�Lo��*�(<m�CA�dj���`{����a����TQ��r�fO�1Roq+z�Y:g�Z�����7ؽ<#˻X.E��Yևqa��<��{Qו�<έ;��_��*��h��Ό$$��yF.p(��6���V;q��ϥ��Q[�P�\�_|N0?�s��-Iʳ"F�(��c�]˴���#��=��{�(rZ�=���uk�S΍N���96dݨ1{"؄�"��d�����؄�Yg`�C���-�!7<l�Y��C����E��4kJ��८����#$����=e>�����,3���y�̮}�kg[�q}Zy@J0=Ix����[J�Kt�-�P���4}�S�(U�&̏A��7��T���A�u���(*=2�b:��+w��f�Y���S �IYr""}��,i�o%����?�(��
ҧ�e�7���Su�se7[g�/��&�v��޵����t ��5Q �YKu*����Ř�����H���듮lb�򘟕�"�MN�M��y�"�o��{�~�U���/
���;z_@�?��&�!�G�P+[�W�RS%v�����֚�B��ֻ�T.��; ��Yz�':Y�j�49Gl�5�Y���pCh�����g��ɴ��|�� eG�C$G~�`B�S$|��.��`�[���U��U�;�k_�~ֿgg��:$���-H��
D?y�$�C�JV3��f��ç�� ���k�����u2��#�(*M����Y��������Db�a�_����%��1���3�/<Mԁ�~1c��fg$�4az]�o���Y&j��8A��Ab��_ዱ-F�!UBL��D�wF]ǫ�?�EZ)z4Ǹ�&|�X����1
�7w�[Cuo��5O�LO5�^���K̗Xo�!(-� S�ՠs��U�J�	��y�[0�݄��z��y�as{W��.Ǒ�ty��֊����M�Ԉ�|5t���Ơq����o���s���f[Y�K��`+6t{����|�/'��j}iY���bŁJƷj�/H22����/�I�2��=�����k!�Y�?(q�v�V�d��g� |���(6��;���8�x�;����u��~)0�+*�_]d�ޱLg*v���n���הC�L�WT��)��������)K;�*e눣����7Y�{�`��+�]O.���#ZF��a�ud��^���Uǥ�� ��2�2x}Fj�w�N�C�8v̓:>	�[�!���B��&'����Mܐ��5O���W���Fd5��'�p/��S��H�/7%��݆*;RY�W9;���J�����Âg�)�-�0�/�3�	��ngO�K�_5[����:md�T��
�\���@�G�m Y����Q��}G�:o��4��G�n��מt���]���� ���ȫ�]���)%V�/�J�o���u���}��1��}@05Q�=
�@	� W=2`X��P�p�"�~�ux�u�k��a)1fd������%#��a_G Aq�*���fp<�K/�V�Ds�-WC��+P ��. k�rp�aH�K~s4F����+ug����$^���6H�a�'�bK]G8��b1C8Jͧs��e!�,�t�!��kVF�E�f�Lɘ��?,�$��OA��k/_/A�m�W�8�KW&R~r&�ƓI(q�6�h��|'��;Ig�6朎�����Gè�H<@��N�U�tq

o}g�h4ه0V��S�L�h<�qH����<É���Q-YS?�,q���V��a�m�� o1�C���Q���S�m�dO�4�`i����/2.�9"��0�?d�%qw�6-�����m֔�?L�,\+�aC��=��Z0���o�n�Ez��q���{��]˔ٺ�e��eB�(⼢��f������] |��eia��!��7_.��|]M�j��w��(�h�=�IҮ�z�e�TsR7��d8i3wo1��'�!B� Q�+:8�x��<�"��4$�B����$ݜk^a�Ì^�}��?n`\�C�Ϋ��m�q�M���K0?��x�>R�1I_��>م���P*�d�e���0V+��@&�6r�ಲ�p_ay����wU4��
�
�V���8�p�V��V��V��S8�O���\Gr�������������y�液_����9��s�ƿ��������X��*9�HH",&%�͞�e�b=�S�z��qSVa�㜐�u@��1��%Ʒ���+3.�0e��'��v��/$�:-ώaJs.�x$v��y�rx`��� ��u�$�b�5�|���Aڗqg�����1:���"d�zT�d���o]a���x>�l��>7f��d�:��*Du�b��ǌ@�k��8���ߗұA�}t]��ދ���qd�9�*���� �|��1N��+j�c��m�u�����a����;؏�z���I�v�[�k���7}���gM��'�X=�ƽ�[��@��f������`gF�t�5�vrU��h�p�M���ٮ�9��+�z��'��U�ơр�:˞�O#��A����3'_�^<�.�[#f��U_�9r�MĂO6${���̭��Vk��T��W����1���J+Ք�eƛ:��j���^�e�o�/��pHAoyH�[��^jJ:��ڷ�QFmc��)x
H��I�\��yoN�M�&�1���j9w�)�[��41�í@`��T��4rH�I"����^�J�����M� I��4��?���![0I����v��1wfRO���:4��d���?�Ø�������Q{K�!{Rď�`dȈj��i7$�K�/W����҃27Y	h���C��������8���[��Zo]x�t�-{H��rM�X�p��y8���1]v8�?�!2�Q0;.��Yv�����).�)@������*l���k�r�����F&��<��%�^�o��!�!3��F3��\���aF�ȅ���]XP �δo31%�g��tPs|a�7ƨ���`�@��U,�ӿ�8@�>��y���t��وMޮ{Ԯp�o�ce���8��Y0<$�7/���Ĕ��ibP�7a2�o�� ;���[�*�������H�zR���O��_�(��h��|���,�N��N�Gh��zޚ�I�M��(D-`�Nq�a_{5��(z<�k/��4���C�v���&���F\"�o~`�\�:��~"��y�<鏯\)9���<�����X:_��n�ѧ��%���Q��=�?{�:�#㷎Y���ri��l����W���ǇU�`�>�=�S�QI�ˍ.i��w� M��v��������&���O�Q�Pg��9c�9H�R����᯽0N`k�V��Py�a���<6�OPB��ޕ9����/�(4+ ��!�~^�iBԋ��y��8�P�#�l"����W�t�?a��֟��toY����%�̒�q�E3ǡ�O(H�~�aU�M 9X���,G���]40ٲ6@��!���aȘ6v���U.{�/qK�����&�@k���0��`�5��O#p^�3d)��H�f����3�Z�J�\��`�M\i���a�C4D��Hk�g&�p�=Q^�1�&=?��?|������B�����%��R�3k-VK���5J����(2�ը᱗扊����b�%C��9U�%L�x�M���
���)��+b�����dv,����r��a�̲c�:R~�$��g�v��B�Pj�#M��M����x���l\�W�I`����|RGa��pUu
��{����'�=1�aX4ܪ�g�����#`�V�h�+��)�j�w]q�R=���\v\��CcEI�e��%�48 B�G��Y�l�a�u�ٽ�5����#�׺;���k1p�RSC�N|�hι��ѡLs�SCL�'��7�J�J�a,���^��ul�/���6���6N�Qw��m�|z�X�qDB�KkbѾ�ϵ�H�E=VBb*�aI��-���3�� ����^���@Z��j�����/��B7a���7ܔ	���bJd�s��׽+ob>�hk��RG\$�x�o�� �x�"p����n)Q77� _��:~�l�Iy,~��i�ّ�]e%���Bi?(��7�IihXֺ;��uy�{x��$hH���mFR�ʞ�լIKԊ��&���T��i� ��C?睯*�$�!����\�+&^�7��v*:9��)1�R6 %<��h_�1��0k�!�8�,cVz������hU��s�G���Bq��)���
K�Ctg���N�;�o;���${� �p+�R��>����0��޻VCy*r����qZjǲ*�����ҥ���k`������	v��'mD�=U��Q�� ��Yr��eL#�t�;��S�\Cō��Fd�VZ��y>�!y&�� ��<��q�䫦�l�48��|8��5����h�j�s�ְ�:������C�}u����;_����g9M�Kr��nM��6J��&O�B&�e�?�Zʼ�e8����0y�	'�����}����h�������襢Z�=�>V} .S�@� 7�2�g/@0���|0��!Z�i��m�X�Gx2v�!��O��n���hyeڴ,3u�`��	�mL(�$R��G��dx^�W��HT��C�e�Gf��1(�HΫ�/(��K�'��c��5�[wj��!����C&/�Gz]v������W�������n��<��-��"��c��=t���%l�P>�g�U7��<S9J�K11$�Cx�l�V�х]���2"yCi��"��yYf�A��k3�)VN�Q�40���Kh�Y'fleي�v��c[���hs���B'U�V�[����D�+�^�{��}>���e�[���$�(V.d�)�z���m�Py>Kq�4���8�{|�|&N�ص%��[<Օ�a�H��wBاrp�e'�椐��>��bŠ����̬��Ƶ2�㦁�,f�}�Ϸ�������\S�=n"i��hk�8�EJ۫)����f*V"?7𭡛��Z�؁H��]Y
��օ�X�9w*k#カ��������}��A��ђ�����md�<�����Gt���:j�B�ST����!���B�¼9�ܤ����Je[��)�澫s�F��iN$Gt��� �s�En���.�fQ!��dG�K��9'�nS�7�j���=�/�L����{E.f�f;�(����^h=IФ�(�u��
�q&Z�[ts�q���&�p�M�;��Ȃ���Enl���8Z���?>�ۏ�[&d������yֹ�d��;Y�	r�H��je�Pg��Z�k+z���E��ҧ�v
�����ѰuDS�O_�v���	)VM�	��L��	�()*N����Ih]G�����tK�8̶�ևh�<�h��5w�!{�λ�t���[`9�kN���ǣpy����A	ŋ3ɜi�p�L������~��}�K|-Qjk���O��N����^l� ���#L
����!(���z5�^dR~�ƿ^hz�$Q����LB
��1���t�;�/�a�̗L�pT�Ƨ?{����x��~m�;⌭^j6��{l�eO	�kj�X��DΚ�� ����$#��|T1Q��V�lc�������Jė�Y�iP�*�ۅ��f�N�/~�S�;'��`��M�T��k��9��e#�(
�>-��A�[|�5"�:�Y� �gp�J#&�@1�����L����+��TD�	��Pќ/��&�Ý�J��Z��}���
RQ�{�.w�:&u���~-!*\�9ȧ$���_��5�@���)�e�KoZs/$v����}	�H�&����H\����_���D��Qѽ������:���)��/�z	zm�s�>zHm���'����$ϲX�y�Rמ2�d"�X�\Vo��R�|��ľ><0��$�@LB%�,���	YO�p�c�N���a�����	��8p�ۧ-��N�$:�B�(��s�ւQ��@uJ~��ܞ���u����yo��ިvI
�"��"��{/v��39ӑ)��u�ʴ�b��B���X����W��w�P>\�"����	&�V�l���Ш����[����; =�n\�e �;w��>��&p����@7�3�+�k/� X_�|��6	S'+��#hd_��ӎH���}H����<���uC�i�����6��&��0S�!H�4�~�o�`�<:�&^��8dq}�o�o�Pt��_:�Mq�̦ѧ�&�0
%��E��tS�i�\��x�c�p䌪�p/��d�Z~�1ⱋwQ2]��.�n+�-�IQ�;�WXP���4Δ�����i�H�����F_:&p��-A�K+��cm��s��M8�,�j���=�B���`�����YB
�����)�FX�Z�,�m�nuD9J9x
5��dF_�-�Hn��r��a�di�d�DXz�Ā3���>��8����A�Ղu3S��oh)�j�v��m���JK��f�����\�,���@�F1��O)~�ɼ[󭺖��V,B�":s�����[Gz&9���~����iG��3��������f��i(��*���ޓ��}�},�/'���S{o�"�^ɑ�_�:���g�Ӕ�G�jˈC���౜O������)�Θ*���	[G�=�}/�m��{ �wG��ؐ^�l:9yl��5G�A��:�\�$I�v\��e�8�Y|*�I��}� ����tR� ��wOO���5봛�b���1E'��X� {nݓa�C��S"s�~{
BM�M�q��N��͹�����m���ܡ�.���OWԂ�s�js �����^�l5If�m`,mYR(�rP�WbMG)��	�
���ZVk�XI(r]�raAa�*�^g����q$ ��OäR����O/Y�qĊ��Z$���̬�N��$����M���/�g�������%;Q���}�	�D�t�
��'��i��Gwq~ϛ����A�f0��~嫮Ce}�G�x
�C~�RD�����05�ȮHF���'$�~#�����y~��WR����|�/IfV�0V�|1�1����7�������-j��`2�7� I�HCA��4�^Q��������ؿOP=&�Vi>�,�Hٙ���/�&�f�V��K�o=-�ϫ,������H� 9��4j�8.��£��!W�yWi��"��&����(T���j�?5��4�(��CS%
����{��栜�=E1��U-��f�Ӹ��&�C�y(�F�½�~���^����,���̣|̖�U�&2��ڒb<�aZ�������b�ۨ$϶��7��5�TE���r&:F�0A���o��e~47@�
�3��g޽R�0�+�.�����������<�"6��w���z�Z����W/ǋ�5��n�����S}��E'^D�|�k��^��\C���\�Me����ݿ��0bFJ�֬�
s�_�KK��z�)ɬ	�,~UuH�K����*���A� ��?��v��:$I.����q�!�q퉃B�9�?�2�GI:v�{���9�(�5O(����Xt�\��J,H������B�m���X�ٻR[QͲ`7����jG�'쀺}N��p�k�dC�^ika˾�!�B�<�dw��
�o�YȫT����s.I��]�����q\F��N�
z.�m�J��9r�yZ�r AJ�	YgE3u���|T�<��U�=��н�7{�+Xh!�-��N�>[�x\,e�^pD�,?����O��T�zي��������,&�R%`�(�VO٥Y��W:ά����#dJ^3�f�m/�(�9���gd�9ޤ9]�)'��*1�O��3`��Y������4  �"	�����^ ��$� Y��Yovʞ|8���_R�N�?�4(��[�uk�؜J�>��;/���&�9�u�-b�l	~��$�v8� EԿY0�Y��v[������n��-�Νc��3dʸ ��Y�Wf�K򌼟s�e���$��Z&���h��{��R�|��}�޾�MA֟`�s��#d�w ��=��گ[J�@��?e+���,h9��l�MC�4�F�A�7_5��+��q��<GF�l���wΕp�R�>x_HHk?������$2��94�@�``���+�{���<�5.�*�U�
�B�U>x7��u��p�����`��>k��s�>�� �m��G�$��EV�1?�6zJr�w�z4��;;Z7Q�@U��`���C�_J�f@�n]#tau6��>�
xr�է�?g���꟧z&\��e��qW{�@)LY����tf����L�öx�n�W*'.|����\z/f�5�-�4� Srh�G�¼��$u����{��ȧ�@���9��n�d�}���~�<�����8���c�q{
1q��v��Ӧ��ιC����2�`g���������/��X衳E����""Ur��0M0���k@��>p�1�Z���I���F�ﲘ��]q���
��}��e{���2� ��KcjY/]R�^Ç�!��X(�|t�b�V�K�Dk/�;��J�M�|ʠv4�SG	rˣk�}~��i��Hէ��`��pW� $���G��t-��T�e���#�U�K�RI��^���G�^���s_�q1N����>��T���$�����>]E8��q�������gs#R�(�bd�@��A���I��ͺ9:0�>�E�P%c'���o�N�>tT#N>z��Do=������M���%
W�=�E�N���m�"���x�J��<`��5@lus�_TX�{���ǉ��_�t-�܌ǜ �"��"&�l_N1�O&8T������`*�Y�>����7�\�>�)ylC �r�IgËQ��>��]���R���'-zK��kU%�B�$�C�F.x݁,9S� uWu�O�K�^�\mD�k�Z�1]1QUб��e�U�ƍ�V�\��o�P�TT�E4+���u{�A��I�����5��lL��.�Z0GZq��1�9��R�q�'��]/.�ka����xI�d���W�x<h?�?��kv X��5�S��<�ŵQ	0<���I���Ɋ�!!dB�el9Ӑ�#��B��W��l���/��Ia�)
�*��'�ަ�
V�bF�~L�0_�v��"���w����l�@[6*,�_���V���L��s�C�lh�Q�>�h2�K��	�YB�6�9-��w$D��$!���aL�{3��>n��l�v@ض<!q������Fԁ��RB)ϓ��5+��n��e�)������/��egM�:nQwv�=�wd�Vk���4�Ô6
��e����(4�[X��mUo�?��<\Y�V��z�z��vYZ���oR��Kj-�W@c�0�����0��o��f�����j!%�g,O�Q�1g5`+���A�0;��:kl�pn���u���e�bA�l%�Kd��5�0�H�b� q������~�ݘ�[� ��x*t���y�N7�E�w�hH���f�*+�Ϗ�R��k����)� ��� ߂ k+/͌����[��$��"�,%�K��/����>�ex��k��5�sl�1��hg��I�mL��O��loTr$R�'���	�������.�i�W#X*J���ռ�Y�?���ҞD���R�
S�ي��Hܙ���:����{�.j�D�W�.��OyL��u�>J�S�B�M��b��'���pV��ɭ���RJ�-��l Փ�H�����Q��q�FD�RS����Y򭃩�����J��Ϻ��QT���JQ.Add�^��/�'�� IM� ��b��� ^���<�uh��|F[j�\E=My��nw���]V�BH�IQ>�M���؛L^���8����A�V�t�N�y�gQ1ƦL���8z�8���ط�җ{��.�����𽌪ޱ'�"U���b�zI
?}�/�1I��;�p�q�ug	[v��5�	d�ֹ4��#J��*�L=@$}�bx ��Pt�N�)�'���`ɼ���=ӷ{іukv?���v~���=���*{ �^��z��x/�д���retq��w3u�k=l��(*�ul�g���r/z�
tl�й�J�۷��U��U7t|��P�|!?���Q�/������%i8��f����Ɵ�O�aٶ���GK��6_#T��A�z�^*����ϕ��%�1FG�Zb�F\�9�a�ͣ�*I�:~������[Z:�6��3�|�,�X�E�����W)�y�W��.���m���3�T�\�#���0c�^��&D�N�4�k�N�/`N��>}�7��P:�<M���Ї=��&��M"�f���n�̳�ۅU���r��F^�F��X��^[�Oe�:d%Ai��R���
��"r�1��M��@�^Do+Z��F�R�W�P�������WG	��w���cߗ�u֋P=���9Fh��85�\4��k�&Bܟ����GUh#��-v���Wc����gu����RJ�q��o���pk�h�8P�,<�ͺ�m�^."'��m��i7�Jk���;w�s頚��]��5l/����a��r������Z^�uc�O�7P�,���ζE���}oXc{i?��#����͂�1^M�k��������v�7β��5	�/���@����\;���ށ��c�r2����Ŏ?fZ��� ,��$��eݮ3Ӫ��t�ҋ���ݔʲk��٨9[���(# [���W�@�A��o=9��v��6����'p2/�[d'3q�[fHʼ����dߋv�(2r�|v��᥻wi �dV�i���j�~�;�\���� r����<��c) Z8����"�� 0o��\M�ą�Lia�b��G�&�J=:��y������z��0&/��;��fʟ6��)@Me�q���,Y������kB�C�b<���b�o<����m��h�4pU֊�\�tm�Z��]�ꌯ�/����a3#�,t��;q[��]Op9p����F���Y���-튔һ�tf�P��%��X�s��&��k�,^�K�G��g��`j�f"�L}�=�X���y_�U�a��Y��;_��*Ҡ�U�o~�븀��m��1�t�1�2aU�1V�[E[���Po(�W"�Y�fķԱ�}�.g|8ߜ�:���K��{�L#�8� ���+�:$�DT�n�"���|�J��-�����x�~��K]�(h����5��5�$q~9�b�/O�F%�¾��W��H�o:|��37�jJ^���g83~���z��Ef�;" ѥ����s_p�h_�����@��B�/`���,���b�7/$q^O�-��bC�N�~@��߸a*�?>!v}��y�j��'PV+���P��U2�l�q��w�KY�t\��<h�Ϋ�"���	OV���ם�x2 U�JP.�o��vepc�|��6� �:G�WJ	�m{��R�O3�H&]��0$d�&���~�3�BP��0'���3���^��L��BA��ѵT>�S�? �� /���g$[�L�����r�d'�1�j����!�?��[ +��RI�[
�%�P8��*P껭�L�<�v�>lrvys���&ع�L���l��I����GN�u
�0����� (��O�p���jB(�/��\�5�����(q���Yƅcc񗬑@��^DK����ouܱ" ����q�-����e׼�[b�z���Z���$�R��DA��'"3$j#�v�z��c�1,ʃ?�^���l
(�R�σz�F���~7��Z�߈��i�;�=��4o����y�ŎK�7��H��	�c��g3.�h�Y��eY��E���6�k�(���uQ�Rf��u��A$
��>jZqh�xil :)�x٫.�qMW�2���GF
�*=�Z|@3v�@~lP�G�|���R���w�wU�s��r.Z%S�hh� '���v��	��z�̸���D�7)?�p��Y�������ti+&��`8E�5|k8��Kvp)������_����8�3Wg��s���Wޟ�*3~ib�S�}��F���F	���6���#���ǌ�3�4c����nɈe%��ͬV`�pפ��9��Ը62*��A�p?�mnf�� ��Ak>T�;�<���O�#�I vÐy-�yiTrq�ev��>8�l���+3Q_w���	�r:i(��n�L�A�vY@�z�Ssv5�9ǀ�LV���5s��j �S��� T%���Y�/�f�\�i�� �]�	�H
 ~1	��ʺH��]�ݣ���s�ϭ{�\��p�6�������OF�'� P�肹�7��Cś3�^P�i���lq��9�n����<o���DXN��w��I�tzL��B=T�X��L�)C���GI-;�yuN���� ���1鶮�i��^�)�T���\lߤ3�S�����i���[ձ��8AE��ER=d�#r6����/Zg�`q2�tC����j�<֗hx����������( 2�!�������x��h3f]df(�h*�?���'��|��7��;��^~���1��.���gC����c��"�^�����Q��"��|"�c'Q�K2��;��F�W*q#X�z}t��nƨ�Dqg��s6mSG},RL��¬�����~�{\׺��i�"w�~d�o�ƅ��I^���z��ä��"Pqd}�Q�`e�:�!��S<�j�r�A�H��ھ?G/8�	�����._yy���C��4�����sS�K�_�z�>2J��k����[�?RŴ˼�g[)I9�
$%$�ܰ�a�K�NQ5���,��l�RNw�JإyQqc��0-��@
�>t%�v1�P�YB��>
e�����},��D�9��3�'�\�G|�����īh�m�J
p+OZ7$�� Ų���1�$�����Lr���̛Ǜ�V��*9��J�?bA�A���"��l� A�h��6����mO,���rc%�ȹ]�y�D&�{_MIº�a�a�$��V4���ֶ�DG/�L���4R�E�������y�7d�Й}r܁�3X� ���q�`yh������ץ1^�;}��V�`�gW}^�P���IN�Kd� ��nt8&��V��d����F�?����}�\5ac�~u��k�,m5G}�kE|���7�� �pV���f��cm	�:t�,��qyh2�B*�9ִ�@{.^�j�/�&�fU����&�;�N�1��cIR}yp���Q��6��a�zX1�B@IA#g�^��0x�U�UJ�t&���|��l%Ma��>�"V����_k�X�I9s�t��xɒp�Nu��CHe�ș�0�/�T�Z/_�XH���|D��R6�}'��,�}��)�:�^5��Z�"$p�vږΰ��wPpa���kU/$-s�ҽB��kaTW��n	b?�5y!Q8>>v�j�ѝ�Q��jn��,D.g1�4�'�Z�\7Z�cw��@|��>��x�+^�˜+nm�9T��g?���Ö����rGHobA$o�M�0�HNɆ"���Z��hT9��T����|�"�a7Ȩ�6ȯ����YTn�2�a��=>����R+pQE��������ZE]����7C]��/'<����K��]�'�#�����ͨ�{�Q^�U�<:����!7O5��+{�'z��JM�a�^�X6�/J���{l��}:��fޔ�S��W�!�J"Q��P��<Ɓu��9a�H7�o׎�*uD�p��i���m�^ ��9���VT��V�Xc#�����oT��p�*r��:6g�{iB��Ep�O�
q;��m�Jb��g��ίG��ys�uI��L�d%���l6~��5z���x��U��&s��8~UC�׌��)n �vx�?�{��A�4h�hȠ�7���@XjX��?z�|cH>�,Gt�[��16Z�E�0,�JA"N��[TծiJ�4�h��1<Z�L?QQ���;�_�\��<��}I �l�oq�\�U/׬�;z��ԭ%�(D�R��̈�:��ÿ6��u��k��j��k�űG����@�b=OJ0'�r=@vrf�䤻k�n�=��8�<����y��S��z�~�|�X����oC2V�0EWxu��5X}q{�*G��f�AE(huT���G�)�{4����Ԥ�Y#�F}qzp����s���ٷ֬c��8QM��˥ zL�vA�\��e��l�����  A��!t5���/�8�څ��d�w��7�{�ܐ)���h}�m�M�ҭG��k�['��d��S��q�*YT�uB�'�
�X�����gO��}DL:���`��.���U��a�l9�U���W3�~�x��̻G��{i�<���E��
�S�Qys2���x�G��{mɕj�&*����Јi(�g2t���Sj�63��m�Z�'`~�Zg?u����NWUf�3$$wD��a-7��w�a��T�+��R��܇$�[��i����oK����-tᯱ�?i<a2J����u]��EwY;�L�r��H��%*#�<(S����X��[G���ަ��@�\N��|�2���OS���j'�S
_�7�oϋ���Ͳ��P�O��֮oD&����F )�K
��'�d<MK��Ǜ)zE'F�����̾��C9���!l	���k�^�z��J1����	�* �+�I�=��,���ڊ�§�u�O���^5���V�;2�^�,ʇC��#��6���S3c�O�E3�h|s�*V�����l"�̣MO(3xO�0v<��?������-�\\���X�	���E�}+� �h��έ���l�/ͬ����#�<��¦��w+��ȩ�°�2I���m08�3��L�Q�O����N�sM��#`:�p�h���w�� ��8�rz�_�0��L�@	Ȉ�E�Muە��i�#�A�/�V���t�K���L5ΓSa�c�pv	�D����y�VOfU-�}�M�,�
��-qe�U�	���v�
$3�Ɖ����AQa�'��O��wO	a>g�c���R�^����u�!��IY�SI�}b�1�/�zE�QQB�|M7@n�B�lD 6@��Q����r�k�8��Ƴn^E}���#\퓊k$��O�jގc�O��F1"�p���Ӱo'���i��
M�w��	�2�A=Qk{b/��>(w�گ��c{ސXI�Q�3���*���؜����e����t�0jw6�9�T����b�#��<���h�J��<#���|Z0�G����7�7�azLbhc��Z��7&/
�ƀr�Vo�==YՌz���!X9��`����˕d��%w�j֬��o\I��cM�kՁ��� ����]/ϱ=:U.�R�jn�GJ�l�p9O����k��l\�s�;�5��������n{���Q �Ye "��Z\Un`	񮤴�pZ�Ɠ4'E��_�b�"b��C�jo����c�u����j ��}apڶ��A�i�ə�7��8�v�}nM?t�##�o+n�d3\qBu�fdW��均˗�t���E(+��(^�1�3,t;l ���g+���o�E\���sz��J�]��ʕ?wH��)�Y���q���2�nD}�����=*;O(�TqV�� n�#6��0�:0~"�@��q�&E ��w�C�eh�sm�m����Pd�Y-�t�)s��X��z���9�Q�O
������(���H�7)�3]�D����S0IFk��������>b3T�|���0[��������?�]$�F,!��\�Bc0����՞ʏF�(�^B��?�b�#�K%3��ҁVٺ���$�!B�^���Z�2!��!��f{7����%A*���J��ĭ�f�K����M���D�� ��b�nq�_u�=G���l�A�\�n0�DD����`Z� ��i�a�����M����9��6�oo��pm���&�IX��E�f��5�F�����oY��_~p���}��O�Ol0��[�|��'��p?_�2�`��
�g&�/.T��r���+]����"� �S�©U]¥<Y�z�ȫ� ��d�f��:JkN �H@LufG�~g���\X+�I�Fg��8X`��}�ȎlA�T��U6�eÃ%����GQC;�ղ>�Xd���x�n�6��e >.���;G,��}�  s��ł���x]M�=ڐͨM���0�(VÌbn�̄����i��J�t�'#�\�=�O�#TVd�N$?��m�AJ��>Qe9����Z��W� �3�������\����/�X1h�9'�jy�5R���W$_-Sa��&ܥq�����v� |؏����U(��t���:�x���M )W�
B���Ic��֒�� �"�,��N���C	m�����Z=W_������A��;۽Ү�d�4$Ƀ�zr=�8(7ހ����3�7��xi�/y���8�82�8]~�`K^k�}R�I����s�vb6�5�n�U����"P� [��v��r��J�� ͧ�Nm�)��7���rH�Ͽ�����N[�g��K�RR���So,���W_	D��lZE�-%G��ґ9]�|��&�'d��Zf��/��_��@W��G�G�hPI ���]��[�s-�'	��)�ԕ�^���ۇ�R��������60덿��m�K��"�
}�E�6�t;sҢH�"�=��
���2+������j/Ր�jGyY��U�^>�N;^ A+Þ\����*;�پ�P%%
̛��^+�9�"P⏼+Zv���Y:����o�]cr�(!���=�w��n���;�-IJ���C��[CW�VPhx�ͭ��"
M�zo�V��;]K��I�+�^�7����Ff0��ch�)��i`9�ro;y�f�ӀI�� e�G1>�M�S׫�u��쩾�D���Ǫ˨;��_�Z���oR|�hf!:����ѹ��h��0���&m��sθ/�1�^�z���i^�En�I�T� Ӌ>����BU�/�s>Qqj?K_����[��t
�ÓqUx�:<���?Z!I �����g�q^��#�i�K�jN�E���밆�H���,2��w��M?^/�B���]���c`?��`���&I�����[@0�x)�}��E��̥�E$R޷��U��$Q�V����]���l,��&�C7�aEW�o0:�#��8������.`�+������Ε<�Z�;���i�����P�����%��h�L5߮��f� p��10,� �,W�g�3l5���4�u�>�ȇ���RzpT/�lV��6O�v�������'
5�@������X*�
��vu�>≖h�g
N�BU�2�T����`�eB��4r��s��G�r���k���|����w��&��u!�p� ����Z;x��s��,���q)�S���P�c�%;ԄVG�fxh:LY��&�Q��"��(�F	 7�F�����sP��R�z\sv<$��U�vϑ/��������?6��U�Dws�R����ˁ��q&0~f����	^C~��YL���L0YH�|��F=���o��Ѥ��6�Penbl@�AK�P��� j�%5���$�ӈA��V����N���3]��e�S�%}�H]�Ȧ��3^cmD^�f4B����g���Yh�f�B~G"\B"j��폥3�4�f:�rt.�s2�O�j��<��ytڜ���0*�� ��i�~<^��t��_��?��yđ٫�!���p���$��*-�'p����M׻�����2���ƹ&�]�v�7�މ#r�F����s��j�<��@Q@R$��UY�=-mUÐbk_`i�RGOI��dN��3����m��o�Vנ�p����	��`U[��N&�� X���9��I%��AU��iZ<Z��LIl����H�s`y���g�|bLf�D�i��R�k���y&{ov�����ا[{�޲���#�ZH��/�A��m ���_��ɹ�B�s�^i��x�%C����dt���(~	�'���ا�k���vW3�4���gv6�l�!��Oy�*q={��O�g�D���X�'��%V�cO�� ��g��c�!�?mz����sr]�����J�8��anM���D�Y1��Ŝ��L���4D�/]�
�E|t��A�YD�ŗ$���1�LG�q*�"��+ܹ��2�[�(Tʥg�$�ŏr�?��9@5�=q��UC��i׎Lh�^�I_ۇy�G�WO�1X���%����7jF_��pW��̙e����}�@C���kj��}�B-q��7��"�a^�㏄��h\6j�p"j��񎞸��{��w�\Jv�W}� /A}�	�?)�t��K��Z�z������{�#�h�f�i w6?BL`+�J̡/)n�fo�}\��м�����m��zR��5���O�^��t�Z�ì�yi���?���Q��U@���"]s2o(v|LyF4Y��]�[����,c�lx�$\��&*��q��î�Z�Io�^G{q�\&d��?(��okiA�/�4�eC�a��N8b;�~�����v�̶�����i��I�7ӂ�|>R���(�$o������[w��$������}hmAӓ�֥�L2y�k�ѷ�d�O�p䜍��i�o��3j˛.m��0��\_�7����M����*]�Y*�A����>;��+�Ȓt9��9T+1qx24��z;��t�? $iI�B�SUu�Y�����i"hHC~�:��{�<I�FL��W2����+���"_�ji{�J �w�0�G'��P}g�'�j��+�}sc�\P��{r���"S��@ns
A�	W{�ˋ[Uk`7�}�R�N/rb���1�e���88P�3i� ����G��D�	m�Ӎ�qtlqtt�Kɾ�����j�����"*�B���K���@��α:�<�%���n��慦�1<Q�&jd�Dgo���Ueb�S��hH���]���!P5q8�ͅ�L"������@�K�7��grn��7�}4������ Ǘou�Zvǝ�P�A ��B4�w]�6�B��Z|�T���`��UmёT͇%'����Y	��n)�̑޻z!ÓbZ<���3q"�5��+i���PS�7��+�8!�����{R����J��6�ڲ�����jcmY�7�3�rFæ�/ �����݉p��C��+���z�L͘B3ob�"�pPD��b�2W�g2ʞ�1Џ2q'�G���R]zF:?��Q�lEfH�1X輞X���a~�.~���Xz3A�[
r�$P"������6�sO��%'!Y�+���$���jSd]�A;5J��R����ΖY͘dCWf,Ͼ�C&��<�f"%�qa�h-}�޹k}|�ɿ��l��W5�W@��4��h��^�"���W=S{(I,��Z��FWZb�� �d��е�Y@z+M^b������*ng$�6�ݼ����]��\?�?ف{���l�*��2p�Z�F�Φ#��}���D����+T���,
�ޥ��P�g�βJγ�����T~�yD� ��a�R�z��+i;bȉ�B�~�M2h�T*b�AȝY�o�/m����NM�
�
��.J�������Y�J��|����Hku��EE̸�����\Vzs��	����nOi_�+���.���EH��bvb�����?L��k(;�Я(����(
E�hA����]��w`����o�)�G5ȧ��{yw��	d�8[>���l���O�*<�$�z��fT����]��:Y .�T���~R�n�g�m�1]GD��L BnM	Y��^�+�`^�d�Y���s0¤�m׻r\ibU,��d�I?.U�ۤ0L�类�E�Q���}���Q2����3� �K��]��B�N�	@����Z!����V���IƝ�I��L*z%V/��YKG��Z�Y����lk)=��;Ր?.lp��A���%z�F,���PۀR䄘�?!i����!l9� ��/�&��ݜ�o�t bl��0�.�Ĕ��M�)�_e�RjA�4�\��.�ɀ��čy����&����{��a]���&�zy�|^�fT@�=N�U�N�igT�5�O��9� 5�O�K��Y}�ELW����n�Pl�
X6q� C��*8��c��Egp��&CF_2"nYxL�g*O�)�a2���@s����b�Z@��	��㵆���s�/Q��v�;�!)F�o~F;*W����h`��ܛ5&*�#|�U�[�5�����uDW��_��J�+��JK�P�KKT��u��5�j�A�/�Xa�ړ�S��F�uj�M���U� _T����bG6LQ3�r�oP��2���-�5f&H٢�	L��ʑ��uǀ�(@\����9��c�U�R��p�|e*ܶ�s���������em�.((�t��� i��Ɛ��~`�������X�}��7cQv����K�(���zAC�*���T��� ��!��H��7���|`<M�`�{c�6�΋�)b'Ѿ��{�^Z3;B��*B�בc���.iڟ��
eC�j�k�d�fǣ���aj�-���'����$��a�b^4�F]��tL�f�;{��Q<9hl`H��@��3�$r!���ŉs��ZE�ߺ!��Vs�|e���fҫ0�"p�z~=H>ٯ[�li������@.7��l��ܱ�j��Ii�o�<��]e���p���;�dz}T��?!5����&g���d?��x�E^��������ǈh3\��vφb#Ȇb����}�ħQ�~��𺶌���z��[l������m\|���3�Z�V��|����j�V|;����T�>�b�>���^=e�^�s!8Z?��&D�����,��n���\���a𲴀�4�,IK����1��I��^#�Xb��ԅ��lX�e��=����ںhQ���,�l�>��j��b�ӬX��W�J�g�y׿bFX�nN�lO��������4�,��dj��l�"&vn�&~���WSUkj���gL$���Ӡ���/��y���%!-8`�3l9��m;�@)��?3A/'�p�cV�q�k$�b̟e|o�h�Ƒ�Q�w�/���iR�U[�i��GE�4U`c��k�t��-��]�z�_��J��ϫ�g�����>v���	H(jBr!qd�y�ݻk���
�l@�
� 0>�m#�]r�m\���b��m��p�~G�@��o����oj� f�3�
�֏ ��Me����(O��f�шx��9O��뽢�� S`�Q-�7"��-�ʐ�0�ֲr@K�T�x_�d�kL�m�M�@ �uQ���NњD��v��S�-�%����wK��'�~j�KY���GYa][���.����EY����!��G
��0dV�1�F堗%��\d�wm�հ�^�{	[���;���ul�ў!��%�J��_
�D�:�����l1D�}�"r�=V���ִ��A�#y�d�?�Ϝ�'g��1�c�2������{;S�&ȇ꼮�%�vL��Jǆ	DH�?����~}�_��'\^��'�ZL>̎��2'����zB� 7y-�DA�V��[�.y+�5�W`j���p;(��Iw'39�̑��-���5�B3��?� I�~�k�c�����:�?��6P]!6I������^���X�~kh ��kng���{���k��^�񙓩���L�[�	w����`E�IC���^����H1�����g7��(eE؍?��AK~�!�vЃ��`euL�;�x.�0cfA=��lV4�@n��P��&�D� �G��#:�Q�{��-;ފsG�s�\�J3�y�Z��5B7]K�y�;��/�������"�А6~�vk�?�I$1��dx���p[~����w�X�%���o-�P&��
ID�o:�|q���=�U.8�YP4�.g����2������!����"�*>�l�0��V_)�{�?g������(�ݱ� ��_��NҤIc4g !�t�ULa�!J=
Q�%<��H
�T�8�=�)i�N�u畳���R����˂6���0C
}3d�f(���m	�l��(-�X�Gc��O���S����O��Y��s�J!7�Jٱ�<2�R�XڲLK�$���9�cz��g?��,v:S�I���姃u_����;o�^��86oxD�KB~a����+R-��*K� a?G,l�3�b�<l x�C�x� ���~}��i4�k�Q�Ǉ����Ǯ|b��������)��-�o��8���K�tT��E�R��X�GQR iƢӖ1�<�>pWR�y��d�<��{�4o����Q�!��>1�:7x�3"�x|O���n��T�UTR譞��2����z9^6.�0�LƋ��ES��H�x�-�?ª�볈Zk��L���^�*��䌵5@=wv�ʛLN)qlv����q%X�oGd�ѥ������~�Y�LP��Rq5�]O9��`���&�*�-k��"+��8�4>@A��gצ$�qM064������)W���S���dͶ��:�q�g������TA�Ll���7��XI�<C��м�F�8@����:��#�\�꒕u�����=�np�~��t�0]}cڗ��� G��6�*����%����ą���1d8����uV�Ҷ;9�(��)��r�-�Ś3Y`��E��jf~�yeME>`�Sz�X4o�Kl�	�4�r<������������LP���~�	(��R�zn�L���],bB��l��ggH�W]��$	ʱ�.6רz,4�Iv\{H�Mx��t�9���H#Q|�&f�Vm󀒕k���R���;J��T
>xCH������������F�Ai�G�ro���nW��{#w�Ld(Z>�p�W)'���:�ѧ���M�4�u|�����*��jRg�'�S��X��y���}��4�C@�J��f�Ž� #���۳�.�2U��<q�W�+��eO'�r`=q��\7���Y5�"Ó��H!�j0}ң˒��v�����O��_������|��D�|R~R$��8V����;'��nc���p��o�7���� $��:�G��*�܎8j��=��]_�=�YB)�i��5T�H`֘�!��4���ty�~���*1 ���1h�
~0�D촨dz:��YƑ��~Ǌ�^�~�E���6�����i��O�ߣ����]��ԥi?��U#��у+����Q$~���h	Lt��f�7�^�G:�_I�:��\L��wg�@���G�����.q?t�� ���fjw[�1�ډܢ��<U��2�~~�����q,i_r��*:��9����hM�yq��?�w���7��O\x:\�Reˑ��C��zd�yݺ�my�`|���|{�V��/����A�	P�F��Y� �,C��	�=�"<�
n�oA��#ߣ([j��Ȏ�v������ἂx�(�x)�T&;�d��?~�p�R}F�L�[���)(1���w�HG�G���+�!*�A�^?h��QR�/���Ƨ�ɣR�y�2 B_��"���I�!�^����JH8�yJ*)v0��.�!k���l^��~��%���ν~fZǨY�_[:t�A,��>�*��^sj��72����?c�ND��֖�zd$��C��>D{�Mω^]G�� �S�a�T{L^�c��'�Et8�"͖uF�ڋZ
s��4�&H����CX�%��L9L�q�d���?�;IZ'٥����0�M}�vsĩXw�- ߦs�`�|�̀�LmzߐU�>S)��QU�s�����,���{F&=�~���l��](7���V�>�~��;e����x�XoI�c�%��C��X�OH  ��09�:�Po2�AɮG9iKS}Qx{8��܋c=V9��h�/���DJ)���5��'/��lo���B�$�Uf؆�X�J��K}[+�AU��`%���#Py�g���r{\֞?8�V�Q�=�؟�����"��h������ W#�Ӑ�(Z�sCdt齱�4�@ڕ�F>��\��`�����#�Kh�(t����;R�Rȱx��#�h�X!����>�����qrUlX�t���c�����~dh![xɘ�<3�����';�j'1��zɟ��;�R�X����5��Y+D]It��G���LO��0����ס�F�j�2�a.�7��[��=�/?�+�N=2o\�1�� �v�8�?]���_�#鞋B�ƴQǣn,�ō���З�������,©��*_��+��<K�9Zo��j�tR��(]ʑ�9y}�o�z��{Y��45��k��X����>BI�	ԇ
�Ϩ����k#��A�gf��?�Y�Q<�G��<1<aU��SZMM�Yb{��Ā�M�g��+������sA[r���~�Lf-4Vh��"�xNe�����N7�i
��8:w�Q�P�q��w�[i�0����q�������_�T����Fp'�Ů�E���̩�T���� �ܔ�	]�ߧ���T	��hON�"�j*��8E��n�+'С����F����{=��%t$���~q1+�eƧ�r�����.��)��QSc����o�d!����:�����ض�
k�4�g?ϼ�4�����w��"�g8�LNdrE�¶�1m����ss�)�(��	Ȼᔢ�<��oga'�Y�����(��Ggh�_�hp8���A�(S��L�f����Q*�w�Am��К�P�$���WD]���@譽�9��֬#*5a ]m��F^_N��?۳���,w\�T��Gnw.��F���
=l�8�x-S!>e�Fh�3K:����{8@S�Q<Cmf���$<p�b==�2��"�
��<t0c��2�l�c
����އ:�-Qz�+�}�^��<-c�zq)���v.��m�]�r"�B���r7e�vX�v��~@"S�yްe���vE�b�'��z�x��,��/-w��w6�D/x�y�gK�n���1��m�I�� V'�Z�r�Y�3����Ǿ�z������Ć�x���Ԕๅ�<�>wW�ԭ�,^�/�"���[M�.���%�6Rhp��K"� 
�1(��U#&��^�1>O��:�L�X���F�k@�&0q�����tI�Ug�nP5_�.�Ic!�R��t���E���1�\�̜v��v�!{���T�CH��o��W�ejz�i�#��Us�eN�\��"A!�bK��w�����-��H�J���������7>�WUh�x[����d�Z�Oe����$���#{��5Lu���>(0�{	hj�Bs�~R���xY��)�>b����o.d7���M���� �ن��9��|Uˑ\݁����Wl������Dh����B3��A9��$�=�&w�����!�[�<�����l6�y���������wcy�w��P�go:1O��s\��<���;��,:NZMؒ�<���/��'?���N���'bJ�a��j��ԋ(K�i��F�2����I��9X���{�2&�B0�O��O���2d�I؏i��M<�t}�&B��o���K�|��/*k���G�g�:�؎(�q�ؐ��Q����fŊ8��!^��ɿǙ`�(۴y�,2q�Y�Q����:KiW�Z�p9�ᾷa=��J ��p�X����\?!�\� �X�A��������e-�j�������!����t*߆�aA�޴A2�M��ڟ�2��:���^�K:���`-��kFi�ň覡���U�|����U�[�<�ڣ���o~oԩ�r~%��-m
��1�s����Z2|���<c*+�?�-��hx�#b��O]$ry'�n�^�y݈Mf�-�������l$ �	+�������������LH�N\B(�k7В\���w�}|"���'q@pK�"�XV�d�!"&Z�~��ހM�2�hK���޾�ޡ[v��5
����.����F4���Ev�p�����9��(���9$�k�~��e}�M�"����$�h�`v>���`���l��1\�Nս	
�_�ݐ@�����G�,��WGxh���������l�cLil����<���A�R�)�;�eh��a�ƨ	�0�m���&��-��/B�ʯ_����w�h�)kIp��Wյ��|�C"ǕlM~�ȩh13�p]O�Y�z��-e� t�}q��A�����e�:�9[ �v(�͛�>�`׍�nrC�>�LWw��rB{!�n�NV�����-����>R5���wS�|m�y	vv�Q��`̄�,�F׮���o��Ⱦ�[��+�	��g?Z1�b��-^e�
q�î��b�͍-�<zW�������$�8$K���i�1�I[��ׅ�.r������~m��POi�/*�=�1L[g�!��.���%�����V��w��`���;'H��W.���P��	�&>���s�_�o������(�����PBC-�Ӊ���)�W�/�jz��0x�vf��c�৏����������!k�I�x��H����������%�Γ�wH���?��-8`1����a��E{�&#f��]:�w�y���D��r/�������� ���Nl�:ȍ=r����h?����L���s����@�K��P���`
;I
L�f�Bm@@�v(�<��5R�� ��� �#��7�-zq����h��HIM0GƶK��p6�5�ʣ���_�`��.J���Tݮ��:{L�fyo�*Cd��\��PX8�[O�c�L�A��(�]�m.S��+9}�
d��t�+��H�=������W�Us`��,=��%���;q�"L���WM{�h���e+�5�E��$�#h���Q=5UJ�.��0�&'C���FEt��쐹�i
�9��2�!�GV��5����c�!�����v���h��=�~/��Iuݲw��c�$q�3/�p���}��XL��WG;:P����B	/7�Hcޟ���D��9�cl�+*AH�|_\}��e�G�i���������{S�=�ƣ����G���M�Z���*~�neE�>
���A�0Ւ<����~�ռ�[����⸧��n�­�qHZ3~�t5��`���V
b}#�J<{^ǩ1�����>j�&m怶b�X6��J������ E��$tѯ_��.�7$�˘?j7S5(4��W&����Ly �]���ωڹ��(!�)��:ʭkL�<I���ƠaO���PD��^o��~o��	4a|��Ar���z��"/����j��>�}Ҝ�t����[},��|���L)�J�]\i�̱�g����5�����%��P&�?dSI�#i�'�}���Yx$�u%�ڑ�.!ѽ�i@������ͱ�E��+����}Vi�*f�J�"6\�+��H��s`/E����C��\yAx�0���"�n������,C[����Br����R��<���( �U_��Uhs�|-��щ�(�g�x#��*M�� �I�AzI��g60�:��$ʐ-~M0���j�gN�rb>��9Y�잆aS�����0���*���c�r��ND�O;F�b�=�M��xVHU�+�:~�d�z�o5�2��AW��"cFzq��K��n���~Z�H�"�c��ʮ�t�����Ȼ��2�����)���s�I�e�,	1����S/�gG��
�����z�$�a���v���C&t����y�5.p'v[G7�#S�l9	���?p%3/O�X��&��5����0��El[�'X
ߪ��4#C�=<Q6�gg{V8qB����+,������u�}s
-��J3�ΪÅ�����3�p��u�"o�>��߬��R�>���]l�`nX�M���~�s�'@ f\;@��P�61�i�˝��y�_E�G3nK�F��H��65u�~�ث)[/�xSȂxܐ�b�$�m���nW�~oƅV�N!�XK�qoר _�iil݈+�������' ~��3>�D3g���k⪤�%m��`������1x���D�x��[�,�=b�lO(ak����lu�TX��z�K��O"jf��eY��+��Hu��߿ �U�f��7`M
 pb:u��Qwa'8��{�q�?��?�;�D!�kyٿ���i�w��NŐ�f�?��2(�Yq��=��׫{��T�x|�.Ӌ�g'�m�9}9��P�f&9T��!�����3e��'���i��!E��ɦI�[i���+���Uwf��e�^me���U���L���
���JW^�:Z�q�~¯�4�('K�㡓���`��m�P	�}5��gpGƟ%V/6�G��G^)*���E�
R�?")�1���:�c����rl��<1v7�ܕ{�4=���1�7IQK�����N�3�YL]�%�\��#ͷ���=��Tg�����ϡ���|�uSy&���]IʊS����xl��ac�P܌�78Ӓ]��ރ���Im֐ۻ*P�|���(u�kfU�����J|�#���n���w-�wG�0�
�S���Y���¼Np��K_���Ѭy�	�h�.�E�Y�����?+/ys��fG$�X��TdEa��Zg���0T����$0�����iOc�>�JÐ1�$J���\����n����Gة3�P�V�-�a{?
�U?1�xҶ�9�&/��\sS�c�������A43�RkWqF����F8t�A�]B>��yҼ��))���ǃ�k=k����/姛�E���C3������;'���-բ�U�#df�y��+`�%"�:熎�>|�Y�\�W�%�P�y&�c��92��sٖ�ۜ�����CƙT��ԓke�%7���}�r�D�l)�kD�RZ��9?�Y�wsR���k5F�m����@,P<妞���v�?�Lz�Q
��v�\xm_��]�J�Be��[<\��m"ޠ!�I�-��ã�/�Gˀ�cR	�����].�(�� nb������u2��ia"]L.v��߼d���t���+���!�HO�/����+n���G�cٟ��V��aU��OWoU%�5��S��7���P� m97R�����:���(�X/n�� �T>5�,���M00k񧢁ҩ��*�v5"~���'�Iþ�<��W��+*��3۽�����fwE!x�qQ�PR�P�͋cU�x«��kfC���ϸ݊k�����޹Ƣ�įp'0�"�gU0����Æ�T���c����s����&��m
cãJR(��ӫ�����N��W�5a���1��/�i�;���{��'!��=���<t��HɞX��ɿ}��a��a? ��[Ԋ.��}N,.�h��7,O��+ -�h��:>�=K#����eS�B���
eu�v�i�G�PָUZ�Sf�4�-���H2�"G{Gat�V�9UU(�%y_���v_T-P�Lj&����A�!\���b��8~�|�X$�P搀��f^0�n� b��5��F0�^�֛�7�Iy�]5��Z�dM#L!�;�6���F���^���[�M�#C�P2=-�Ĭ���_ ��΁��.����p�rG]�����1�so��٧\���S޴�.V�C����˟ָj��C
���QŏmB�lm�{���M��-z6� ����9�j�ޣ�F:.`vd}�|_�]:F�T}*G�����y�	���;A�q�Q����^8k�����{^[�Az"\����ě���!�����vO$���kyog��\uv>j�G�L��,B�W_�z���A��o_Yo�.�
�@�;o|Fs�!��ۿ�@<����s���^+�h�h�I�"��9�^�R���iS��̦,1"Lݿůr��\S�OP�;F̓G��9\?���Z�:��WA1�w���z�dj�\:GyF_��^0��S9^�6����O|�9@+=��m�|o%悹{t�A����͕N�)��!�ke��TP 
.>��@�k�Y���w!�����G�a�����9�G�
j��ԩٰ͚9BF���_�ŻF�O��#6�K�X(<>�YCmY�<�H���T'�r�B���GUr�W\I�/˲R_"�:�"��_ �4T�T:߆�d�4GG�y�?��R��*�{���m刿J�h�k��׋_��E[��|'�B�!�+�-�}DW�l�՘�;*R�q�Mb�_�2��M#� ����R�k?j=�z�hvTL,�Y�""FP���j�]������u&ϟ�ȘYL�4�z����-���Κ����&h�m�{�b[^7�+����`ٽ�5-��bcDU�n���}�!�I�U?ҥ�D\޸�V�P�Ȓja�<�c���ў�H�J��c��v���t�3f:���o��:G�Ap��t e�Pe��ׇA��@WJ�R)� ޢOn��o�nsnu�{�L݄Z\����H��5#i��Ǎ�=̂�gu��d�!�Q[j����U���$�
��DƔn
T�R�5�"�F��3�d;��Z;��f����NQ�i+o�����_�hU��w�_d��'#� ɝo��.c�{GwR��Ք�؋N���[:�|U#&M�Q��?�CW^�C�EX��yu��<�q:��b�t���K`��I��e��/�ͩ��a0ČB����F��
��n)u�?�V#�U�Ɨd��&L�vŖ�@��.�>j�8��x��'\G����U�nI�jj�1�C���d�7���yF�\�H�3���4��Di�=3e�h0�����ؠ�3k���p�{����+77�&J՜����w&���I�)��G!����0�a�� d�玅�	}������s�,z��2(�]v�T?L���|�`��_)��(�㦾�ѳM����V�
F]�\G��A�u��Z��"zEB��c6�s�Dqo��!%V%�Rn���s8?8|��ҫ�� G:�^��Uv5�#q�~	f m�\�i����o�4tc�l�q�Kce�i(������<(}Z�/フ���Z��ʅ;�
�Ճ����%[���C�o>Z$������-�͕P�A�~�O����w���DcX���qw��t�?Ƚ�O�_���R�LL��/U_j*�:#m��r�I����[�!SH(+Ch��-+p>f�h6L�z�2�N~9���o������ņXA��E����O�@՞�.�a�B�]�HTobh
�Q�.��q'G���&���޺ӳ�<�� �by��U�!=�6���l�-Ly}�_%&MKL�M�1Lo:V���l�u�DR�j�p��J�
��|�'��o�ōH��֢����7pҤ���-0z���a�%1��.kn
�Z�8sh�֍���{FWk�vL�nb7����U�a�Y�o��	n�}p�	C���A�΁��>�	�٤�F�͍򿣥^�����%D.��M��ly��tgsƛt+�d�!�qt���ϑ��{�P��,��״�̮hϯ�I�0�P�.�.ǐ�uw
 $~4'�9��&t��H����u���p@��F����C�UotO��<1�z�*��2�_mG�S��c��9��C�mM���<ѴF�0�U��3�[��jݴ����`��v�
=O o�h���ρ8؅��ax�Ohu��^�;��sD%g�ۤ�>�����\ܰi��f=��N�3�pj����:�N�4�q���VS��a�	��1�e_6g����+�-��H'N�$p���l�����X'��]�uV��;#nH^�b�H���nmMG��jm����P�PFl;2]v��(R~C�Eh�ȑq�EE��(�?�x˧���;	�l�.яM��0�t���7��0>��e�+�lV��r�,SyW�� ֢�`�[�I!��߆�^�o�����J9-������о��h�3[�(��rTh�d��.��P�!,(�F����f]%�\,="Hqd�l����I�(�'=m~Yh��Gax/t���8`T综|�Lc|�C8�9��ڮ�`�b'��!���792�h���Atn���q�����j���.�湡"����/���>iQ���������rLOW��=
�~[�dB�_�e����n��g��j���:Pg���8�����<{����b�m��
�e�����w���o~E��N�~��D�H�ڼ��A���≵��W�sD;���s�M��'ߚ�M2��d0�:��~{]/?W��(p���03��2U>��+D�GH+0+$$�ߖD���c��;��h��?���`�K�-	�����t�~t�~R�8�7�l��}Dm�z@����L1/e��`��s��yt�aɜ�~N 0�o��k!���9�J4��Md\@�m���S�%�7����Es�0�Hd���R�p+'{���h
nw@P�]L������C[�me��l\ݻ��_�b����~| ��iE��*��a��Lֶf�gtõ��q/�P�g����e���Ǎ�Z�7�gWa���f)ɻP@~��~�*2
X����)�j�g2�T�s�_%M�1	�t�a�˳��x�7`�V���d����¢�4��xK!?kݚ�s��V<t�����瞥7�C�ݭ����w~ls���h o,dU�����܉��e�+h�r�~��Y	zIA���KU��)��8����f���z��\�,���U��T�� ��V�:�I�6T�!�1��e9Ƀ<hS�L�~�I肠c���FZ�9X�+�}�ݎe�aH��2	0�k���E%`M #1L�R����D!#�4�J�����`;n�I-�=�n�&�~�oE�0���m��Om�,�;���6��L��>'�CD��w��-q�Ih%e�H1�K�[��;�U�W�.~E���r�2�������w �.�ԎY�P�W�\o�4�2���s9�S��u2��"��O��Юa�7혬R�gW4��o7˻�Gq.�J����,�E�]�xg�H�]Ut������*]��R�e�Y���ņ7�p�ceiہ�����nV2����&���)����y�F��K�S�%Z���llSp+gcIB�;��I���,�R��\�ASf+g�]E��n�H�M_��!��7��pm-�.	�����M��g�,�G"�KMP���܀sL�.]VL��B]��e�����^��3R-�F9��xix�p��,��T3��0�^�
͖�d'&+O;��$���>�كL���[�
謾V��i���0A�N�x������>Y5�pj���3������$e�pr�ݹ��=��O���O��'F+zo�X'J_��Q*�N��o�lߺy�H�p��� ��]�e4!�!-a7��ݬ+��t''>gI�*vXq��^�a����	��-�3�b�#<�w��*�Â�I���	��Hb��,�fX\�1�G����9��kd!���@H��/�v������k���Nh����|��}DV?Ns�RWכۆK��3��YN�3������k.W|��G���J�:�G#U,�!��S6�̾���'PG���<8�O9�����k�m��lww1<R���'4�-���>`W���,'1 !j��}� ���B\\JKB�R맯�����cS!��V��"����d=�_Wԇ�K�C���Am�8� �� Ë#-}ˑ	 c�2�t���r�����8�~w��Y �b[�8K ��R�\��{�Qzh�<�����q��Ln��=Os�0��f��W���u<,�~S��F5���D��J����D_�V�����o�/7o=yM��\�5�}�T�S�@�ϊ0en'T'��l� Ύop�H���Uҡ��x�&��@%Z�*,����֮���L���O˃��HH�p�e�rBcy(�3מ���5!zl�JLǰ�P���Ĝ���:��:��]�A����;��nM)j�O4"��X#�K�-k�r�$U��`�3��Xt|�A~�i�r|���F�����`N1�5}4ǘ�ҺqK +���fz(�I&�+W�#�rm@���`:�x���h"���J����V���2Ȑ��CC(��Vb4P�� k�����ʇ����p-�G5�j��X�\��I9M��wE'2�� �Ce�cS��ig�b�1�ݬ��n�@S�,?^��n�m�*�	/3���J�-&pk��ۜ�1��q��Be[�m:��ה��;�$y'bE;�J�uz�*���ـ��h�4f^E��՗�O4�G��a����u�o��ʗ�*����C�4=ډ[�k$�Ӥ�Ρ-��c��B��Lb�+�-3%� !,�Z�y��5���R$O� �D*�O��2{�GȘ�޾�OQ����]?���p��_"%��5�����w�Ty��w�������O����Rz~�$�7s}��Ȳ�-_����t�XfFT� 5�T��բ�+`�S_�Pd>:���d�2.56�e�;����D�������aȔ>�k0�f"�c��A��:��n���a��ߗZ��i룳�U��+sE ��O�>�"����A��P�u*I,9$�@��q��f�H��?&��c*L}Ⱦ�nΐr�,����\I�9-R[�}��	L������aj����E �E-=��.8�Д��_F�`�-��[�(b	�,��=�+#�� ��x�f;�S��,ڟq֊�6!��	��*JO+����0��I?^�9�\(�G=k-Kp_�S"u�몳�w}��ZO+����K���o��8�i 
�Y�HH�ѷiP�Ռ���z����5R0C�{������͢�zx�]���*��8��U�ާ(
	�)��
Ȍd��$��O.T��u��9j����v���	�~�j�*nuI�c�J ��d�m-&X7Ⱦ��	�U�����(��Q,*8`���|�n[�{���а��fu~	�T��L����g���7�h�E��MY+e�����T���֥�`,�˅~ڋr��S���1�{���)/�[��r"[�~��¶��,*�ii��;4��^�ڦ ⼾��=�ڠ�E��j�I�_vxt8۝.��+ʏ�F�<�!���M�0�q`#+�΅G�V)Ə��(�\(��X�/��'9z0X�:|�g�m�#�Y�ٙ�ђ���+�r���m󭟢a�~�&���Z�{��z�##�&
W��qt�9��W���3�y�C�l�����h�B�Vy��}\r����'振5����u���tB���*��ID<���d�ǉ�8Gm.���e�9rt�E>��\���o���}xZ� h<����|����9q5����~g��6'@y���CRB�D?�p���Y��JE�7~-���������G%��!����k!�u��P8n��/孩-�T����ΪG�q
��g1�4�W�3��^b���Ι�������e%�&>�\�0~��i��}u�/٭����d�Y��%�9q��?b��8�u'���f|��N���y�{�(�_�ŵA�� 
��4q��ւ�:�5��Fj{
���>SF>������^��(��6��ㅛ�&����r Tֺ��~l��\)M�}��짆lʿ��ޢt�r,��\���k�oh=$�=�������Y^E���5k������hw���'�ȱS�`6�Хã���T�*N�aΦ���Lڙ��+*����m8_��2d��cNn>t���>gz�\n�4��ᓧ�l��0n,c�k���O���j�m|�N�ԜJ���[�yN���wfN��R��\�v���W�茴f�����*���=d/K��ψ*֬���F|��CV���j)з4��Ѓ��rײ30?@N���k\�`��A6�":Xu��`��e��Mް���2#K@$iBT�\����o�A�۞ k3D�H	��8pG���vM4��K���J�d�YD��1�"{����	���<g�tc/w�ȡ�㻣y\�,�E�c��cƨl�(^�61EQVbAQ��y��Na�i���);��@Ũ$���YM�"$�]@i	��0D�@*�'Ն�.�^w��?�v��	#�F�z8�[�"�c�!
���O\3�?5J��l|���Ĕ$VS�
�]s�ĴdZ؂`&�8���{��"X�����B	�gB�tZ�x�`����	Z�N)������)4b�Z�A�i��1a��e��n�r����j��7Bԋ�����a3��Ed��岊�k�I��]֔>�V�]���7�ߋ��i_j�~>R-����J�!I/�\�H _�My�r�-�W���ZQ�E�:zi�
1����H��DDX�f���!B��B�"���s�f&t/R�h~�~����WA������p�`G��Awi�SW��}��<Ґs�JL;H�t�eebΓWks��Y1qЅ��<q����(�i��ɢ�|K��NL���, ?�m�	%uZ?�d
�E����+�-2YΒ�F�e�M��y3ǔ]�'Ni�U/�E�dA��Y��yD~i^��P��N�D���,]=�����(�W�~�$��vz6>$�|���b�E���b1�����-����p��g�?��'m/㼣�-��z	2=��8 4�4����T~f����HTj\�m )_Аa�eL?~��e��x�B2�n?�clN���Ƀ

ƕ�	��U�ڑm��!�¿�:��P^�Zxg���(��Is:�K��
�m� ڱ�J~��	K�Y.�1���.i���U�Ű�)73dq���\NuJJS���>��H�WJ8�����7���.Ç���jJ�YJn�Z��I��f���.$�qj�FP�Z88��3'��>����K��^r�].Ȱ���Z?j�5�~[�~5P�ω��^�{�E�HŸd*m�Ag4�6=B�7�ŧ^�e�
1(#�pa�u��xi((h���,JqA���I��?o��Չz�-��p�AH�%�
��S��d�)Q�;��n貒u*U�]��Xh�� �����Wz�Dૉ0PqrF(ROq��"�s����`�1�&�������z
�}r�qؙw`������֋� Y!�#{|���l�o��Ld1�����`yq�z�6W��[
�s���ǣ��Q�]�r���H6�U��	l������}M~ڤA��c�>��A�p��V�Hu;�Ě�bDy?A��	�;��E�ғ���b�[��`e\voy~C19K� �3�'�P����� �'%������S�FרC��D��O��a�kS��:&�3�X��C=}@�#Q��`����^~����)L���t2��D�m��$�b/�0M�B�Wh_��w�9��8�!�}H��!�|{�"���[h>~Oc�x��TGK��\,�D[���вYp:�$��[w7X�!n�~����<J��K�n�M'�����vJ�~�锥(�duAf)4{\	/�G��[��讀Ȳ�E�?�8+_�p��_Kk&���n3JA���4�ʕ�>��cB<*Jw,<Dhk�C�4�e���.ި-mށ�WR�����'�pP�)}��T���8�~���8��pj����V���ꒀ�>��'\����8-B�fo1�=�{S�G��8"���z���W����0�S$>�%f�[+7���ɳ'8�ʤE���h��V��F4�IC��J�i��"����T�+6�\��]u���s����]*��@>?(�#�n>��sF�F	u��k�@8xۼ8�E�NVW�l�(��qk�[�����a�y�*p�cfP��.��y�z�DE�~K��0��,��?&��Z���Ą�c2vPϛ�l6�Kz�D����[��U飑WIB\:����p:UP<��5���Ԟ��mՍ���`f�e����m����^T�Ut�~��Y��;T��Th��Xj^�������|9�-�̍�9�^0�f��Q�i��'�$D����*5mѳ��+T:�r��o�S��P�A�4S����Ӊ�����&Je�	� �I^�bӛ_���w�1�5aL��9����V]�@�����I����.\C$&��r���3&m��,A�og-�቟.����E������>PW��Q�%���6�=Ȟ��� 3���9$2���ɻᓉ��+�&j>@UP�چℊ���y�'(�KJJQѣ_��Id�"��( �@�(��k�	�D�_N[&"����N��8*��l�l�Ϲ̥=^�6@�T1�ϩf���w�uP,C꣨�)GՏ��>:��j1/�tp��L�|�bf��A%��gQ�=e�0J��ѡ4�k}c,cNu��W.��Ϭ`���������z�;ʆ�&�{��-++�o���D��ͳ���pH�X��{���%�1�l��VY�%I/��K'��-�8��3�!M>�!f9[�ڹެ&��Ƒ���5미C�G־^{��6PO���˥Dv~�;�a��\K@�8u���d��h61�q��(@�������x���Z� R��b4(4���[sԉ�Ì��Y�a���,k��0��!VZh{MVb���\7�!(m�(~�`��/��N+]��+x�������V9
�Д�����z����/!ql���0ǖh����n�Ui��غ���o�r@� 
T+���%��t�����M��	0�d$�_V�Wx����������o(�R����S�<U鐠L��	U�yj��=2YC�@�u��i
�H{�Ptu���c��׎���x(�H���� �)eE��L���|% =G3%U���vŃ@�Q���.�(�c�V�O���!ӛ0s���h��Z� �ρ�y��)
�D��k����f0�y�нy#Z2pg;v��{�qb�&�C�]Pq�<���%�6 �����;�?�Wa��z�m;��(~)�=t0��d��z���>�"�7�Q�|Ţ��hW��ԇ�;)v�,�#��������p�x��������ө7�p��Sx	�1r�Y��y��y�ƺ8F�`��?�ߋ=�oy��1H��#[�kT�"����n�Zʁg���&|�r�֤Xu����-$�q���U��0���q�يP�����E�x�Z6�&{x�`ݩ���0{+����@B��P��m��bb;HD�0�I��b���*LAT��A[jy8������2�w��$[*�J�^C�T�k�[!�S2h���D}���B�m�r�Y�ǽ��D�m�z���nl����~[�����F�!���;�1���?4�Ė���!@-:=	
�(ˇ3���\-�n%��"�^8�H���|(�����F�2Y�?q�%��0Qэ��aՏ�����b2C��G���}��T'���~�y��Qs%&:�/����A7�_CǧMvd|ʯ��h#���2Y}{&�%��[�6j�Ds�Cd4�Ә��A�0�����p�����,�v{g �5���}�e�l�����o${�m���@u*П7�O�����z��<�~ȴ��I��F	�Oʘ�(	�KX6�D'u���1�5��6������{Ћ��`{|�����#�įW�#��W�n�V�Wǁ���;c-�zdN�CHkcg���cr5�56YdC�X���_�m`ѽ�;���U���;��S�zs'|�w�����OfiG����U�~i�:�oӅ<�����6��p^���w�/Q��Dw�C��Î~8�U
�g�^nÿ�+n@@�q�����嘠5�=�>~���I�������
���P9��o�
�ޝ]�`/�}���,�>�ү��7T�Lg�잍��ґ�ܕ�-d���H|�9{'ڑ�0W-�~�"��v:"��V��;:�1?YK�M�0�t^�����t�d����@�ݽi�ߩ��#���=�"������ɒ	^�]�^o�j���T�I�v2�;��&;�p�w�(�n�U���)NU9�(�����;R*� `�H��t�D��K��t$�1����j�7��x�:M�qn���ft�H'5��b<D2h;�
B�1�L������{m�&D<Z^��n͝s��e+4�#�S I�	��M+	9T��x8ŝ�ͺ��_��d>�prr����h�B�Q�p�����%��VD�:���*�#��
�DؾZ����j�ĉ��ܿ�
Ձ����f�g�Ɇ����o�Cy�L_j�O3�.�}"�WE�����������,��� c%�ϏtYcͬ�C�cm�>�K�쭥*���C�ʱR���i� � �%�|�z��NH���@���g�p�t���7��^��+'o2��љ���t���%W'B�.�� �_9k=��������
aU�"�ͣ|�yё���n�xw�Gv!��vrM��B�#m��IO�+�ӎ�1s�c�!bs:f�Dbe��(����3[��SvE��/(��yH���ֱ�?�_�1A>D�v���CU����{)�,N��L%Sszn~�K`��B	o{i%�HqM��
��`9�ERqY�MyQ��)t/I!z�Uj�y�VEO��*k�?��5�$י=�<����B����#ɼrH8,�d�x\S&��<�R��O�{{	DcVu��@�/t���!8��T�+��|��~���aI`��|cS,�4���]�0�&J6���*M�j���|Y��ϲ����k�4g0��`tU�����x���@�;'�8����1�v���A��ܲ}�c4�Eb�/;C�J���GeR��"����R�T�x���j�i�P5*�c{ƣ���EQH��I�'sW`��Tx�B%%�t��;�!�l�}��6�M��Ҳ����L�І"Û}�zZa�v\��[��}�ş>���4=Y0��k�D�˚`
<&�����ҭ�S��K&��@I��Bd���P�?��.S����t�|��R�Ez2K����(a�������|'�gwm���94(&��*	�ndV���}��T�Bo�h>�Z��I4F%�	glw&�Zy�D����	Z�sV�)�����m4��-=B��lN��j��8����T�-Eҵh��H�'9l�}8(�gnkYf�h�`��Q~ut'�ɻK���
���_�8g��M��Q$�N��玄q�v(��v5,/�m��*z���o`�3�V���a>J�cM<�"��hyzOa���}���Q�>�Qlu>��*�{�ZM���J"��Tcd�C�HӏY�����QJp{������m{Ŗ[�z��pҳ�<i�k�:f]��Jq�]k��xuP��Cr� 5˾��-�Y�	;揈*��'�?���`����+�Q��E��~�� �'�~�w�_����e� �f��s
��ݐ9=�R!2l?@�J��ٙ��(����s�0��V����.ܥ�7?�1���������3���^���G�V,�x��([;� � �ٓe�
:�I��at	�ȓ�x�a�,{��iV�b<�����:wAZ;V]C��elglZo�{�� ���ӧC�Y^qA��"
�~�G<'�����<�}�@.7Z�C��S�U�K�)ݩq=�_�)s6��8�M�Q]o���.��b�g��E��ʆ��S#���IdĦ���KJXw�����)'�W�����*�4d�ZB������Pa6u�|�.>1��u�e��
7M(��1�85��1c}��/�n:���q�,ɴI3�=o�3anT^ ��mٽ?|#P�V��|�g=K���~���`����ʛXZ/Kqp9�i�{A3�!H���v9f7�(WԀ�u8����w��T��w�^��Uz�δ��&_��?�	gQ���Jݴ�ƣʆ�L��B+Yn�?�ݜ��q_{�i�w>(�-����S7�%U},c%n~�#=,��_)�x�;F�sN�/-��	�|5Nq�ԧ�P��P��n���t͍�`HB�F�ܿ�����sŻ�=�MSy�ky�G�X>t 1��޶I߈���m�Z"m�tbW�@�>xM�����u��u/w8IR+�A{季�Р�*|���>�;oM;	�;�ڲ�N~��PE�����R][+KԽ�"�9(=P+	�U��S`q[�x�.V�L���cI�L�[r�����|%�#	�A�A��yp��E[��/�ʹH˫\���\�-��sv��|U]�|`����2O��<B�8���2�W���_���E����$�#�d[��o�l�!��4���`\U�GԔ�Q>>�(�^��WZt!�<�n���ي��E�lK%ڭ�8|t�(60����L������9�}Q�I�c"�*�PZ����b�T�D�y�RN��d��2�SN� �9 �r�to�hG�I���/)�bp"{@`�f�ǂJ�#��ﰪ$2���(�
g�B�'g�j`cb�$w/XA��dF��ЭD��g�&߿fo��a�M�&G I��C�.��n�^(}�q7i>7���m�C��Խ �.�&�(��֭+��U��Ӣ���2b�;ia!F~�Q�0�<
��`�^1�^k��V�E@7�&�0 ���FdʏW��7|��7�fjt��_�� ��G�����"��ԒRO�����G���^��D�(ͦ�
�!�>�zG<x@	z�V^9j>d0�f(`fyo��7]M�>����q����~��N��9�*k���TD�n�T)b[KEO�$����S�h��c'� �C7]�§��e��ȧ{�} �j6�t(�s�C�|�̒t	=V���=Ҵ���<}7���q��\D5��ы��xFՂ �nr��*���b$/��3�9&o����_�
l Y��F8�ꛮ�~��Y�~�~Ltؿ�x��ŀ��Aݸ幅��Z��\�B
)�4!D����O��X���K[�)��J����ֶ�}v�'�C̣�z�)@��[鎅�mP
���`�<�}�)�G�~px�Q����E�>j��L�Z��|<O�3$���kKTL�%�G�\�F��.;Z�����/>.{���ȑ�4Mn�oz�q�{�P�m�8E��$����
� Y��#-2�g�X�^��q�k�L�o�GZ"��x3�h،�o)����l	��v��ǯ�p��-`MFx@�5��8䂢,��ɹ~����D��_�����w?mv��T�W*�Q���Ps�ٶaq߁h��0��������{�6U08���
�D+ΰݨ�Eim;�"�rRXxPe��34��e�wr��`��1L����7����N�鬔$�)�~��i_Z�#)vY��ܰI]K��pϣ����5�:��`�j;��d�Fpz��n2җ��Z��6�da�DB�rZRˋ2���e��T��e�f���SE:AwRV+A�t��[&��&���0%@Z�����J���5����j.!����cn&�Lk��{���}r-����N����xk�� ����\�k�ɷ��e�&�[�=���M�&����!��������f��������=�1	3-��Z���E{��:4eE ��	����ʮ'���Ӧ/��ٍ��J5]�!��Zp+{󮇇`��hl_�χoz͛��D�2�+<?�ھE�s�>j�_�6-��A���z?�H�T�y�YH�N����؜l�@:�z�nз&ꙹ�$��G�v �Z�2���X��=�jw���;'�z�G�k�l�/��)�~�{r��>�.Y�!JX�JT�dK�<�E"��<�����k��mR���%�e�B���-�h��z�������݋ѩ����{LFW��11�}�<�*h
����ߙ�%q/�k���ٲn����|�C�kGXBW���Ē���V���Z�@SG,�ݔU_����X�f<#K}������*(Z�F: Cؕ�b5?iȦ�K&`�x�x�l"E����zť�����k��ZBv�R[,U d[���	�=�؉��7�-������2��?��j�n5��'ɓ�ѹ~�M�1�7��VPw�E������	� ��~����uPc��QJg��4���k�E/Z�u����DW�jJ���'�qn[����O@���=��igXT��a��睆�����qIj�WH��	������9d7+ZA����R�ǃ*B�pH��=9���U_y1pӨ�������~'�"K���_�x�ڊ4!��$<_��V��-W���RhJ!�������1g6-e��0�r'��<)�X�N�;`o��ߕH��^��k����?�9Ya���uK�"�-qDP�r��t���u^�K����^v���ކ��{�< �ly{�t���\9�����G�+1�*>�(����A����S�qm���������V��d'���2O:W"���`7���l�*�֠�x�	�29*>'r���p��:St�,Z�>n��X��� ؄15����!VY�]�̼M���-����P�;�(m�[vh��M��^wq����rݾ��D�C,�$�����Ua�F~� �:�{���JYX�R�f(v�(\J����5�?2�6�Te-��`�~C������"H�Řl~n=�z��E�0�ڭ�HݸT�\�e&�{��n��m�-y��9���w������2�y�C5𷩶T�����}]aUgn9� ����Hq��9���0#��^£A���N�J ��	���,����L�Й	�ab����V�n<󅼸r��7�=�%A���{l��l2��ʂ�=��ݢ���<H��N�N�0�E+�t�q{�~�Y���Ȁo�t�U��s�Rh��4��ć�.(��Sɾbݭ����)�B�.��Cc��sX��G�y���3��qx�A�xyuU���ʅ;3>�����Yt�3��dcVK�5H�׺B�s�'"�24�r���| ���*:]t̅��	���;Y�o�=YVȀ�� {U�B�,WvT�̼��.*���l��e֕q+J+Z��ڇ/8�ɡ&�h���75�w��ɚ��u'^�Ʋ������� b4����fM���D��[�O=wp�������#�<��`�L  0���7'kވ�V�?�#[i:�/�`�>���������X1�M���;����K�>��ZJ��X\\m��E�/��Re%�f�V�.9e��Kc�툹�ƦC滕tz*N72���V��a��xI�=�GˎY��^9�0���7�4�cI���;Ml�u2K'��P4��d�
��7����p,)$��b�������*�EzII�X�|v����EA\���'����v`���/Y�N2.��3��޸>R�,��oQ��x5h����	�3{N���73����}">ꤐS��O���[���n�!L6��y47�m[������h2`����,*B*u@4Z%v"���z2������q����q��$Vaȵ�&���Ս�������r�̷lpU�m�h>�@����K#'Z$xz���^���5��!��+��#�%���������F!^*��	��GS�1��$N��W ��P$:���"��b4 c�8˘>�d!󶡁�UD�	/���2 ��_
�lbi	�'}��鉼��Wl7�hT����_���[����UpA��!���~<�}��-�]��׺(g5u,e:U.2�g��e��=�]5�[��.��U��/K&UZFr|U<}QG��*5a�XV��Q���޵�x��Ȳ�g�N"@��W��Ni�Os?��j��U�nk��	w	E|fQ4Y�l�L�A[C�w�?Pf�. K�}��C��O���KabU���OF�Gs$ھE4�/$E�^=� 0' ���1�`�֬��e����Bz�(���gB"��j�ԯZ��]����eñ׊�����:x�����jxvN�_��I3�nv���/]�};K��P�ͩ*�e�G�tyl�#:�y���"u�N������
�삄�m+Pwl��$j~Ɋ	�#W�u�H*}'�9�#��%B#�u)*!Sg/�B�JcAw	o!�����~)q����I�sщ��>��,�����"XC!��7��X�_�C��
Te��,�6E�r�S����TiA�][pjk��)FC4�D�����Ꮐ���0x��P�!5�%C2�f�U���L�f�)�u�:<oK�M3|;�&��v��pv =��U�Y�<݀&�N%V�%���-l�J"��H�d��<��[��[{6�M����%k�|FdsG�4r���T���2�xJ�;�����^cq��[����I��ȃ�Xc�1��Ԙ�b;�<O������|��wt�M��{:�V������%��2G�z��~�;�p/%�K.��&����ƧY "g���-=�o|79�6���
���kg��o,%G�2�y�#��m��<M�G��p��5)�Ԥ�͛����G���^�d,y�o����G��ZjR�^�s��;��ˤ�ٱ��b��7i�=����5���rd��)h �f�P}��%���l�3�NT=9��Y�?��oL���� :Z�b�����{�C����j��4����6j�l���7`ﹽ��H�R-����n�ٞT�E�C�дAC�r&I��r�;�oTQ�˟�0x�B���p���"�G��5��C��b�/�lr��"��F��<�|�T8DM�J�R0��T)�p����qQ��,x��I�dӒ��׃��w`	k�L{���-c�\X<���s���a�<��H_�JU���[�/�"���<[>�� ��
8� ��lD��.UB� <�Z���j��Z�Q��1�� ݤ�rB� ҄�8Z7�X����qXhgh��7��]N�)  �3�VA�&�����"�qҮ��Z�BN��LPu���K��;R�&��m����O�}�s�ehC$��F�nL���d�l&�>�Z9'̕W��n���n?�`���<U�x�W�<���4���<&AsF:{�%���K���/仓X�
�UC�n���4%O�cr�$*DL���A��zz�U0�{�4�1T���JC��b_����6+$�6P!)�����f��C-�x�ၹk�F���Ǐ� ���҄�1��<�j�,w���i��)&-�7�J���N���f.�Ω���8Q����;���$�6���l�HR)2���׮EV����.x��!u�en%H"�RQ��&9��T΢��X�j]�4��l��F�����^6�Z}P��}�	��AO��.��\z�-i�@���14��%�X�H����ꔪ	�$�$'�+с�� P�9�]�+8&��Tz��+.R>�6����	���nz���g^x�eD��	<����0�B��c��2�~�ǒ?��U�`2#軤Ǚ帒jD��;<w`��)��D��O��i�3�^$Wt�q8��'������#8�בҘ>|�<P�FK��U�O���"}���E���e�_�+5�iF��2u�<�;(�����>���|�L�1��j�֬]�\m$�'�"��w���rH&�{���A��ǹ����&P �#�]pLK�n�� $s[ �o�߷�Z����;n_�1Eo�������F�ղUK�����>���]>�����PA��\�$����~�*��u���Ȑ��zl#�V��eD�:�q�8��$��)ZX��>kkpKi�����X�p�ey����J`(!K���5cބ�� �E���b�O����O���S�"���
�E"��#����6����P@ܤ�d�@�@M�eo.>�O #�E_
=�Ԕ�^q'EM8��)�^��NW�,�_�X��62Z���l��	�kL����&�_K$��p�xLc��:(L!Z�a���w��m�X�
�7���[jk�tѢ{`^"f'Y�X�]�I&q�l3������bi�qW���	�~��w;Q}-=%�:�Q(5H���me+�W#��
w���������Z}M4/ȃG�9V�m?<K��Wq�a5�^�x~�^7C�������(*� I�yY���.e��`+Q���}f��f{͏��v&��K�r���|@gFK�98�G��+"�ꪘ�61ݒ�5���@��l�JXs��E���A��H�8D$�A���;�ȣ�/��1赻`99ǆ������C�ɔ
���T������fm&��-��J��3�y�gH1��>5t�W1��fb�Xأ#�צ����-60���;c~��u�*�)bk�8�r����]� �E��.O�~��t��C�8�QbT׼p�m�ڪ��K׃�L=�ŏ��n�u��X�A0`���`/�iM��m8%�΋K�͋F�t�w�v8�����¤��Pk �l���)p�a�b��¸1c���n
E�
�hU���O������9Y�g2�La�C:�!(pq����n2.`6��<M�0�#�]�`�%�qVB}Mc`�$T��w��f�Z��ߧa�	�u�6|C�d�����y�c�3����ʅ���|q��D�t>�ɈՏK�`<�xV\��Cx\/�&�KV���ńҶ�=2`Mw4�ea󙚑oc��c��Uӊ?P3t16�I}�&g�$��h8i�5j@J���mU��1�҃��_x<���D�9���i�ߔ����6��� �6�t�^�����W�?*���Ԡ��֏%�c����!U3�j��%���S�Qj!T���vd���<�� WB�M���-e��{J�9�0�8(�_ć�;��`�H�R0R��^���Wj�V1�7����"�&?�&�"�?w�P���f�0x�~�*.|lo�� ����7����u�50�9�k�V��e/��܃Ĳps�Qߺ��1��P��d�3]M-Ix����uϿ7.��x���sG���Q�J"S��DY�|Z� c�A`E�a|,B�[FJg����R�jnn�{&\֋1��w������mܰPknT�v��q��~�%�T�E�R�� ���F�}`�|�0�0�]s�kDM �*- Z،�Nw�ɔ�3g�dX������x-�٩s���$������.��ו�r�=3��c��d{l))���<@-�]Α4���%|A�
@�
I�3:=�O& �yO�w7�)_�Ng���ID�}k�������#X%"E�v�7�ߢ!�Wl��v�$�wحk�K߬��ۛ�Ua�5��� 5���N��7��yR$��K-O��d+�q��7�3䆄���ba��D3q;E�Q�Y��*���i�	��L�G��[��.;�����U<�	3+s9n����E��󘓭d̨}�)$���g��.�:�ݽF��Pm&RCZTq�o7?�ц���X&�%X�͛1��M`Y�>4g�(4<�~��pB���T�_Y�9��m�fl�� � V�BS��{���Ĳ3n(`\�(�C��� �T���Jw�F�%=hӛ���6R���B-[٘1mMA0�&�}�bh����(w�vg� n­�7��C�>�0�v|�?Z�R%��[d��$�~����ÿPL��8˰���E|��9��&Ti�o�TIA6-���P"�%1���u2��.6�8�޿hP0AN�R-�����ǯl$6h�S7��;���V�,W�+:oϪƷ'?F���di]kk�S-!}^B9=H�wI*_B��5
��G��Ar���3�\��9�ڽ���N؜�h#��/|Ƃ��i+�ߟ�z	o�BJ�L�r�OM�3雥�I2��U�tD��35�k8�87��Ձ���0%Fc�+�3α�Q�>)Rq�T.��؜_	2_��]�;C/���jFq��	�,��8X$�������(.ɫ�/%l������:Cݼ5��)G2��8_�m�X ��N(O,5�_�E´�����KQq�l�=����-Llw�Jʓ�� e��]_8=�R��OY?&����Ԩ��wZ�g�sD�����T<�BaHj��p
@�Z���ռ��)�B����, u�.³z�������z��곅����I�y=��)=]����^	�w!��f~��h�S��{��(������9��"�����Pv�U��e�LJ�zrը�q6*9��u&�u���6��ص�q�P��+��~HXl��ݜ�Fܹ$r �ެh1g?~��1�$'�XS Z߻�<�����{<G>(�y�)�AD���(_;���l����\���e�?�bS�#|�S	(��LKp���&��{�C
��p�V��&+�Rl�R�iS�
�W��+!O��9�BWDɞ%���+�`A� Jy�A��+��m�B������ZH��"E����Ȥ[�	 �r�7�����&m������4h��z��#�P��Wg�r(�~7-�ԁ"ijE��(�L��[NV7��j�'���DĭђZy�*0"��Y}y���&4���u��))�[��pu�)	I�C�uS�,���G��b�� g4�B��R�A�
p�0H��X
	�]�
��$�$é=�����['����
�����N���{�X��c��� ȀoB���mY~xp.�P�C�jpgZ�Jv=�G״!�/�D��D��c��N"=E=��*��� �KjU�a��B�����A���tڶE˪�,���T*�`���<�r ��뇌�;G6�^��ݓ�R���U�|��L>�(��8G錽�(���s'��ѷ����;�J��H���� �Z@��˔	���L9���Z �����wY�Sw��uo"\#7ƜoR!�(ñ�_~��O��9��Ň�/-.ME���A'��U�$���-�˦� ���?t����.�.�57��i�U�{=�I:W�����?<hu�.;\�~�X�د�:��F؉i�2xC�*��_#�*&m��~@�~��*��n�i���v�Jҳ���%����?���y���IT�SKz�Va(��"��T��J+3D�I3'�l�$�����!��vJj��޾���I;�Y%k�$�~��z:��h*q�����
_�q��^�[�d/I/_8�/�0��~� �a/�2˶QWd�-Lt�@���<e���\��?�:�5(�J�I�QZ4D��| �
/¥Y�����ͤ]ʫ�o�k��慵w�K4Y_v:e��w�����1'�e�@z0�c�����ش�6y��O�����mH��c�5u��f��  A���T�Q�y�P�D^��B���S~�����B���ٵ�#lny�JL����Ýi*�%���F@���kB��yӟ�����f��	�,�)�v��l��)��Cv�`lt[�)��Y)O�u��]��a�������8�W�;��Y����$�����&��	͠}�$�|f�aX��n�1��+�A��4T&��O���h[������a��.�u�rϸ����1��T�NΪ��V��>�Zf�[Y���ټy-���Z�vI�~������0k`#�KE�c^���T�"���;�TE�b3CߺC�a)� ���q����J,{]X�O̏?wE�VS�T�0��j8�����mQ#r����kXX�d�t�'�U�~Q�d֕�� �ٶ�;SQ������1��v�{��}K6���ю5������;�s�����)�����N�	�|�yb�NBV�J�o;����أ� ��`S��r��@�D�~����cP�w�_LL�^����p� �΃���5�B�Gx'NjݜoU�^�������=�>�z*G�^�{�$O���ξ��VU���MWZB�V�.ݺї��� �#��r�܈<H��`%n�-E����+.�~3(v9EZ�G�E*�1���~R����ߞ��EiӨQ�'\s@��l�LQ�k	<Yo�wTy�Z��/�̀��J�8�)l~����*.@����������ܔ�x���O玷�7eL&^C��R��3n�-gp�U�8?�xpY
���W]�%^Y�+�Z�w�R�B}�>�� ���nl�b~�1#�ڹS�G�ejbNtqA3۽���I��VdHuhMWX��Y��!��T���-64���|,�H���校�|�����A�m,�q�k^�@��$+�pB��TG� �1ƥ⼢�_Z����-u^P��N_�S���a�
j�
�ey�\\(^}��D �j��C:�X�4���\�K����V�&Q<@��"���9rVE�(�{�aVU�R�aTH	Zq�9f��ok�����m4\��r��k B�k|*�[y��vi���dT!�F���G��ڗ|��;��KZ���*Ӳ��yDd(2ԩq���Dҏ��VV=k�RqjH����QR\�iǽ��� ��GE�`D#g�R�D ���H���]]�u/�rEl�v_��vH)^�o�6���ZH�;69��cb:���H�EeT���JJ��9��1S@(ڍO��Ra^1������%Ξ	g����e�d -�U�%�p(D��o�Zd(�����ў���^���ٸ\�ot*��1��g���er�G7MMV l��^tAՍ��x��Vuޒi��`�| ����vc�V����շ�1Xe�$7؉5⢒H�/9��i�F϶�g����>��dL�����3�õ����0���&���Ԉd���J*�w^
�S�$�i�I5�F��Y�'+�J��a�?J�l_�d~<��c�6b�-�c�ǯļ��f0))��c5�쨄�}�7��ֵ��;�YBY� ���X��W����3�E{$Uݖ19����o���[?��;�e�B����l\�H��ӹD=LKn̓OB�&ץ����x���Y)�ҝ�W�$�ۄv)�� �[�	p�v���ʿ"�!��m�$��n�7$�?�W���OH�������j�#X�,~�C��e9��QjE]O�e1�'{�&A�Ԓv�I��X`���p�S��?:8��^by0���-���7~�3.�N�F�g�Yk�z��~�<E�m_��������T��q<j�z��0B�gy4�?؁�e���뉑>�����=�a�-X�h�������������&����w�w����n[�ʧ�L�ğVD]�W�ܙk&�����{)K�Sp=n<5p����7_%��CW�����G'#��p�(������������9�:t��l������U���J�Vԡ��tY���/��i;�S�B:9�PCug��	������I��k�A�_+�W,�<�lĢ�T�?� 'R�.�d�Iu_��/�=ԭ�1l� �t]���&�6í�^���l���3�7�SG�j���?��W�r<�HT�?I7Ev��J�< 
5`�{���=��Q�@��%����%�������D��hx��y��vK�a�φ�-����`Z���n�����I��"e)%�bLU��U�(�R�f��F��0�Cn����PL�((c���!7D���i�1ߧK	�M>l���� (R���YL���r7�:�5�� 7�Ab3p�A���+;R����b1�tE�����`�`M�p�:7 ��j�EXF���c2��y�[|)��3Dq/������\P�&��ȥ8t�����%-�^�^Sb!���R���5�D	�{~��w�
|�7� N�!䣁g�#���Q��<�D/��F��	��F��"-5�=�4
��l� ��l�6�h�S�h�t��ʜ�Ǉ�q���58*Pv���U^�':�7������\��8�q���ߟ��T΁싲o �u5 ,�>w����cZڻ'xc�`�E�n���c����%�l��Y�֣-��k�5��}~wAB
�&��Mpm��<��^����N}�(��T�~f�/O)ܛ�G��MM%�G�H�v֏�(�%c��;�urT ~	W��dS�� �Y%	xv�e�k�����
�hp��[�Q1:����Y�3M�ty����=Q��$�I��Z�>���=�W������ j�����YXm�M\D�^h^�'b�COLW1�r�;�k{;T
��)���=U�Cx��I����m�&�^�	Cˑ=���h�*[=T�g�����7q�hc�o��=$t^�H�l�KP�2b|B(Ռ�G���x5ً�c�`17��Z��r7t�2Yl��+0��۪��INO$��� ����|,��9�+�[C \.`Sϱ���(|VF�T#,4I*�]����
Vg9}I6r�S�\AF�VS2h�l�.MW�`;�V}"K���ղ�U�����D�G-�ҏ��H�yFqrY*�4ߕ��S�D��A��#Β�A�j��Q��v) �U��]����e��@2ʒ^,���~���v8IV4!葾:Om��!F��P��d(եm+�� /�q �^��ۤ1n�������>�֦�cj{z�N�	�wE_y�	Z�8�������?�y��$Q�tv�<9O�h��S��gb�q�=��Ul��y�K��N$�y�s��[�v*Z�<��(�E]�
��6d��3�f����e���U����p=�Pԑ�M�
�9�S@ĉ�Zr���7]U �����_��w�S6�\8�,÷�עM:;29��!��-�w�]U[�g���rH��윀��B���c-�OS��Z�p��N��H�gaK��c�"��{ )B�����S����̲Q/}>)�L�s��R*?�Fr��>�~�"�b݄���
m�uM��)k�;Y'�:��ڇ7l^��@1� ݔ���^�Q�`���3��*VEU��̗��lH�|+�N-Hӕ�E��Y�D6gv����G>�{�c�	:������.^��1�A����V?�zdШ=Z����:ǹ�4]�%X�w�� ���ڮ���D#�OԫK�w|:h�δ;4ze]�5V4l�I�r�o]b�G�>dwA������T�|*�7&]7",��(��	�#�G�&{z΍ ��&"�nq���騽1�,�r+�x�
O�p@�1��ɵ��ULM�f��M86�F[w��-�G�6&�A��A~z����#���Y�c}��Ոس��_Q^n��u+���#��8�PU�Dl451p\	�A��|��S���m�8J?$��)΀	Q�Z:zA��]w4:21����MC��)�7��$���ҏ��~���P!_����G#�_ϐ���!e���;G�8�e�9��
���1#(<��L�Ђ�ہ�*�`z�����(-��ǝq)�$�f�'}�<���p���_:��X�����sX��� \�_3��Ț��a�_��w�8�{GG2/}�*o_�6>���j	��4/R�O��v<4 �O�a2��+�UԖ|���;�%T�k���V�_�bvd:}�o��c�k���	��ϛɩa/�3�/�HI�l�M�^���e��Q�C�"��f�b�Y�o��(�2g�E���Naq���8`h+"�&����{F{A�]�F�"H(\P�yZ\l���+t�v�^{����[*O@����q���u��V!k]g���j����0Qˍ/B�ʐ�H�.�*抋��+Gڔ�n�[X��\������Z)�k�U�yp_�[�	Ȕ;:�N���(�6xe����Ci�ϕ0��Z����j�`����@&!�E��W�̶�'i$fZ�Q�Z�+#�:�e�'���5}���l���>�FG_�
�l�:q	F��c���S� .
���KD" +�h�X�VV_������Z�lA�KY)cJ_i�͋n(>��\+$��jC�+d�iɊ�ݍ'/M^���"��G;�M?��!JJ?}�Ѱ85�w�P>��	#Zf8+�ywq���=ħګ� �$��$�1�3I"?aKVЁ�^P����R�i�@kI��~�D���L�\�M�Na�NL��-���_�V�@Y������WcR�e��3�mqSϞ�-E ] ÞL�4ϼ���}�A�tQ
��Y�	�W�20��[��Գ-��Rc=>U�{?�WɠN�s^ ��b���(���A.��[��S�qD�f(�{Rr=8�IL9yCxY���<|Yj���ll�H��S�Y�*R@�W���d�����Ji�1�xkƬ��X/�Iɡm�<#�hu���8�kl������~�nb�G�&����z��3LKN�P�`�B�w|�9)�w���Ū�4	��x#K.3hqi�����l�&���h��o�}�i2�9�l�8��k��=Ka¹K��Ej�d��1�x��4�hR�vT@wz�R{Y�k��S�˘�4ŉ��8�=E�4aXn^ 'Fa�S	���p;%�'$�f<�h�%������Ԯ�5L�*B1)�,_��`l�Q��w3�*%�p�B��A6��CM�r�@ԙ�1�-��U�gG+�n�+�үs+\G�y��wI��.��ԌHv ��s8�����+K�8�k9>&QP�r���qP.!�1P���-�v!�2E�4�ٔ<������_�6���0113�_[�7q*|�OB��A4�rj��vo÷g�)H�t�<(��=�K7)r�����l�T���ϕ�=k[4@RU��9w�Qg�V���W<����m�����""��Ō1�ZJ%r�Hu�~&��£���'�½R��ʌ���J!0 ���|��.%Ġ)�����jn)���,�Zs���u��m�6F]l��>�F5j��ɔe����'�8��6����@��R��R���ϛG�s���z8 �0��q谣�/f�c���� ��JX^�- 0��q���FN����c���kȐ���}Ű��b���8��1��C��K�����J'_o��u����?/�Dm�l���U6���/��NZ��o��0Yk�� >��Bp�e_����\��3��3h�O�>�i�{%VV�D�������j�>�h����4Zg���$;�	��'	�y���l�,�躗�X4�v2{��{��I׿��~jb�0>�l۠x�ճ�Q�B*&����;�h�<�'����TK-X�%B_����>�k��ub�'�ZJ��
]�����F��}�07��������5�W�hWvM����_�?�%�Gz�#p:dk��wEW=��rT�ⴰ�Y=�n�fcKֈ*9���m\�;-�ӊ�����eec)mǈ�h��dɿR�2�_���s�J5y�'>CF��QfF]zԶ[�� #_x}�gW��5���a�W1B���8��bώASA��vj��o8���㛗U���Ԣ�����xFU�:�'}M;��^PN�~+k^h��&�~�
D»t絒�@���P=ދ����
� �~�&��~��E�ay��XnA�ɐR�����̏��&�_�&�6��OR��%`Cӱ4���pO)�����|Eq�������"6����C.�$KR>��@�+�+�,1~��5;^�����Y�_�����ߵ��0����7l�w�)��*�EH^/'�|_Ϡ:�|��{���t�ѧ�)g�U���|�gğ�{�]���c����/@�r����E�{0�x3���dg�h1}RKr��d1c��� ����ev��iޓ�G/ tY���S��+��	t��Ӏ&d��"]'=r��k�~���ﳒ�25����䱊�0h��a#�h��Pr6��������6	��k�*&���[]���`����Jk3'�,��Y�T�/�G ��q�և�g�u�h��ٹ���<��(��=��'#��RE}\��\8`ԜS�t��L���j�f���;�q�LE��&7�����Y�LB�Y�����B@���t�>��I��;��1mƗ��zug��L҇�@q	��ٖE8��X�K�GO{�2�z|]���<��r�`�W�t�zϤȻ�^�z�U�Q� +8$ÓZ��^[�1e���Ya�H!N�н�3+�@:tj��a��8��1[ȩ���bz��B�`��-�mҘ�^�f��T��&s�����-Q'�Å�* ���2�/{�����	��?�;u�?s�G���)a�z�!��2#0à�,V�H%��ERf�����`�mk4(v.J�O�m���}es�yßN�>q�.�g�4�gu�o�!�y�h�p1{�Dw�;�n �m�Q^����y�6�c��}3?I�|���g��������u<�������pTz��,��8���S��+h�e����з�E{�:h�ZNI.D�F�D�n%o�@uM���e����%���4ex��	"���?n
2�臨{;��o4#x�쇈KC��'��&�RA64�Y=X�u���:;1	@ �����IgUj��I�z�\�p6lb����'���B�����-�j�{�����N���A����#�kz��"��Eȁ�ĥ��vg�T�9���0!�7�K�.M���o���(���ʞ}%��y�����'�Z�VO�6H�$X��1k��Ȅ�jJW^�븫>o1�Y��ޮ�v.�a6x!��RyI�:9�# �
�Rc1��}�KY�)���R��0�H9��A�����|@j�7`�u���b���Q'�g�7^���;%G�ē����Vt<T�vEK��v9��T�m��斒!�ď���b�8༡�{��4���g)Q�M��4@Fd"�@\A�M? �Q�Nݰ�Â.0ֆ�~nW�Ey�[򮕀m�R�{�'+w]ue6W�Iɒ�_v����;��a��曗���y�П6��ױ��E���;_p��:�^��H�\�1��޷���cr\Akhʭ�s�uk򙵃�)�V
G�Ї?k�z��	��/���o�_*��:t��$�V:��I3[:O�z�������g�������%����Jos�E��Ƒ��NQEV��P��=3�c�e��k�N��	�l�W&~p���E&
�hs]�#gjS<&�5�Q�xt6֠M�y�u�@m�K\{8��Vq!�%�=�Dy՛β�	�F���/]B����2����}�G@�Jh��+v����랠JLa1u��q ,t�G�,=S�#�6�U�5�{��N��Q�٭a�wݏ1�y6�E��y���ȳy!�n�	��_v'2'%X�R�汶��M�~��ĉ�r)h��W�R�&�#N��ѹBF9"�� �'�1����<��w��M�� ���hV��M����J�+�d�!�c�`<o�#%.���u��q��ݷ^�%ʸ�\A鮻�_�4���Mee'0��������pR@���"�?����8�Z`\R
b�����BFB#����\@�� �nW��_��L�՚�.�Xf:��ϭ���b%���I
���0m7��ӶV$�Mk�'3�Wn>炶��7�����(>q������L�6IS���{�����x:]�ྠq$���x��`};GF���!	SI�{}�_W�!�R�6]��C9��a�602Gӗ�6��P+��x��.O�Ř�>����j0�k"�`QT�U���uH�N�-;���`rH���jyv��:  cރ���=%����p�k�i�3�����*|�5Vf����|Gx�]9�4s�ˣ�M��O0��=V�L�r��)=�e����n����Bø���=�=���a�� �2lݵw�ǀ�+f����}Ү��?�M���o�4f�	˿1�9l�z�"����C֌j���*�{���6ƞ3�Ѥ%�	CQ�h��id�8:c��>5`zDc��&��2�$h�39э9�Y]�,2ì T4�l@�N['V���o\)��QJq�j���'����1�?2y�=8��]s�#���#�Rp���=$|VԎ��d�K����،�����8���q�5��<�������$��R9�/��(I�t;���
���Ȼ���w��]W Y���_w��b*O��-�eަA��E ��:�u��G&��s��s\�QX"�doPL?�����1ڦ1�Hե��Qy�ܰ^��Є�0F2���~v�%mc͔4�j�
~d*I���^���dY]���� ��y�Os5�X�3��Mgd�: S?�-��ʿ)E'�S$������*ݻ�Q��ߞ?R7LR�i33*V�,��<�־ZN��`:�KU�a�B�*H~Vi%�6~���Gm����z�Wb��+���F��ZjE�( �G�Zma��R_�0��T���"�m����~��%���Yn���� � l�cye9>��<pf=CՄ�*g�X��H0�t$3�,T���|cv��;���.K���V���Ճ�YjĢdJ��4����/����l5jFpx��T�q��q��7�4k1�K��Nt� 
 z��d��ps�ָ�΢ ��@�W��C�z7R�9U�J��Q���ں�l|���Kp4�+ˊ��>T��kRuYC�'0�H�,��(L:Z-��x�����{�jh�yҜx�Y%7���2�J�U�A�Y��8�x
���U�֓�V��������d�c3�d��ˠ� ��Y��
9u�?n������8��4yT�V]NFk��įa`1�ylP͔
�{��L�,E	K�[T�/H�N�菬l9n�CT�W(u���d�ő�(�Dy�G �ݳ��Z�(qnA�P�!�w �������������|FBAJL��pc��;��=@����%ٟPo��YO[��%��˅��Q�)��s����U�Y�V�S�>a8h��{����
v
��w0as�OhO��������۪n?k�9�h�|�c�M>���h�!$�O�@Ot�����1�!�	���:�Lg��wI;�Y<q�9�;����[_�h�*��&go�୰$\~
�4��xb/0��8�T����}g�TZff|E�	#�D�\��`Q0��k�A��/0ߓ����B���-B\$�(}&!��/C��ސpYs���~��L�2tW�;����=+���\�˼�%
A���1���)�ʅ��-&57��X�u���>Wr�%�MBw���H+�����/��5���Z�O�A*�|ra[�Yh'��]M&��O)��7���=~�X�B�;������ti�Ս�����BJ�S���1� ��TUah���7K7����p�t�2ߛ�LU�z�k�\��$i�=���YSy���W(.WI�0�]I�Ϯ{A�h��tēH�M���I��	�Pd�Z��3����n���s��$u�$#��_������X�`A�u� ��wtD���%�ֳߛp��b��A��p�L���`$dg���g�]f�1�A��_�G�C�@IՑ;���6u �
��[��Y�h���`]m�2�\p����� ���u�&v%��Y�'�y�����v�"�O����/�"����8ފ��ҳ��W?��h̟�M��ρ��w���()WK��@5��kCc�xwa@*��?�����8��r��ɘ���$��n��-�kz�n��:�i�U���$?^k�ˏ����eY9|B��%���թ2<���I�%#�{��6u.b�d�#�];Ӑ���d��H������z:շ6�� ��~�u!�P�Y���@�F7���V1~�3�-(6J��ZR-c �m�R�=3/OFWR����3�]������j���疘�]/�&G��"M���g�L%�>_T^��͔t]˲���n��u� �U�[�^�J�������_�j��Ź���q��!����`tII���{��V�����FrE�h�G7�$48���d�0d�+ac)٢��W���YpiN���'b���z]���]<^斤�(�{/��`W;��?H�͍$�q��E|�fIŀ|�A��gj8u����� 0�]�����V���khOq����"�ܭ�5�T�9�NuX�Md�A�E��9��_+(������M�pl��ip�m�d5�3*��r2+�R�[h��!��|���E$�2�@�A�e��J:��`���83�y&(~�������<�x)\O������������Yй��G�Y�4�)��D|2��z�Y�`��Yѽ(�@�p�������� ��ad;.��q�m�,�%~W�s��3�s�2�M2�P�p�2p��Y�2`< y�E��KO��i�J^f���m�z���% Ёr�G���Q�Ρ6ٿ����}Չ���Y�_c��7��O��6[r0����;������=�T�s����zQ�*
�"�J���E^�2oy��j�P��([QK]���f%�Z��fF�W�|���PA#k����B�mpYr3V�s�U`����LP��y�*�[��Ǚ��N�m��R�AX�cg; �����wTVSv`Z���׵?�7*��c���#<����0�7 ��^.�);Y��g���8�'n�Ł\!^�2�5��P����"�L���Ye�#'��o�6��6guZ��������%�b>��c�I�E��
�� %M�LY���4�*�	�Խ����y^/���:���u딤�.�V�է�q���BIеF>��2}F0��mR��ȝXcd�(s)��SM�� �OB��rP�҆�Uڸ�os=f�h�IPyD���Z�D�:~t8�2���Hᠼް�/�-�Z��^dS���6'���P%bN��7��.ъ��*.���_#@˯gΣ�e� �P�4J0M���*�iA+I�z߭�?/Q`8�Y��ii\1��ų}̷C���N�&�����u�B	⍤�Fh��F�Sk'4�~�Ѭ�����kg3�?~ͼ�h�BN��bV������~vϯ�Ѕـ9�hן~���׼`ES��=�y�̤ꫮT:ف��x�[�Ɉj�.ǔ���l"�I����c:��B�MK�e�jʂ�)Qo(�r+ץ��=���64��9j��d>C��g��M����Y�yV]+��}f	������n����.�郿7"���.��w��]�򘯰��H�P�p�gq���+@!G�ۂԲCҸt�&�`fȦ��{��
�z����0q?�жs%2l #������:H{+*�Sߊ��_���D��6QZ���y�do�����3�N�_�6�A9p�5p�	γX�í��P��2C?���S��w�\O��G"��nv-���2|Ç9kFԶM�%Y�td���	����Z���LV���*�G�ǋ9����P����F9]�W�0����\l�T���}Â�����Z+`���AD�A&)�s�ɴ�����:N�������=^���ͭ���K8�?��=�-�U峉��%2[r�� @���-O��؝.7B��>T��(3B�;؋�ľ9*�[���M��4���x!�@]8\�T/�F~��� �\R��6����������(�k�!�řo��u/��ߋ�p��KI�M����L=x���D����^�\�"��;�ڛ� }�w�<óq�ƫ]��<us��.݁в�ɷOЭ��"]��=cW�~�(��1��rDĚ�����W���)*i�um�I�$*���j�?��,�i�5)�Ôt�a#2�3 �Bjv�����7{}"���D2������1������Ano͌x��1%�,�` N"��U$h�{�5�(�}��~��B�q��AH�1e\$��$��ln�x����;b���}�.�) H�ڗ$y]JD[�����K(K��DW~dG��n+\_�K=�鈳��,�F�xk|Ar緍�E� �Ⱦ`���
M쇓��i��Yw���FT}�"�y����y�%����z�QLRVt��'�Ryj�G���l8�H��"�}H���g%�5Ql��{Ͳ�]���0��O"Č9���r��8ѽ�T��tf���ґ����%��Ծ�@h��χ/A5	���p��e�����qfR�I��'eƙ�q�k��h�����+���",ԪU���a,R�q�����T�KI�l͜|4�'��,%v�W�Ѝ$?\_yoKص�!�uNZY��T���p$[d��"�|��>7��������G���ư��x��}������w>O��Η�^6!��O�ET�M�Z�2{4�2�%��$h���H�?Ik�`���c�/��RL4�X� 1��1t�@U�m%P��65��ɑI�!¼�O�0P��E6���ՙ�H2��Gˑ�	���@6�i��	�F�l�v6�NBԹ�[�(�s�l����'�8��G����Ѫ��Lɦ���� �P^�t�����J���B��[�
Dظ�z$����Ƞ�cE�d5Bq��tB����Wo�x4]�d�'�n��tS^&����@�|$��=.T�3�`]�ߙ���-s~���g�)S�T��g,"Ŧ�mع��'��>�{����Zt<���8�@L���Zc5���{��d��Fd�v�&�_�*�a��3�aC:uA.@�l�=!;pu����lSg'a�{/�E�g\�=ӁMC�ɺ�=m��w?s�-��=~�y��3e�9�g��gz��OSL��8��~[�nţ L;g��omU7���#�9a�.vT��]MN��A�9��z4�G����V�{5�cT���[d?T����|���1<E���Ȅ�w̞BT!�� �ʎ��_�E?۹���7��g���tokYvgޮ�!��t@�0�������4��$�F³{��)���g�{`�$����;��
�P/��a��A�'�1Wr�s��p$�T��c�&/Ƴ���:�gh�7��-j�o��a2rl�-�V��<�.}�R�(,f�[�b��e�/��;��#S:��2Ü��t�dׇ�8[Rk��?�~�N�M8k�#Y��6  Яcdh0��s���Tk��뙉��Cb1�=9s���A�O6���5W���搖E~c�61�_[elU�"�'
G�� 5�,8��+��v�(���"<j2Pl
��u�A����a;��#n���sT��<IM�GP��;�*UD�O���v�ыGw�:a�0:��'1q�K��Yz3d_�eև��F;T�`$x��R�B�f2b�?ot�Ci�`��bnFV�d��2<v=�U!�2�ynRM� f9�'���ˢ������P�7����I�g�q(��ë�ҿ�w�IWGg���Lu���:ƺ�p�E3��{� �B� ��Rc�A��u�틿�7IZA8�uW�K+DŌ�K���z����ق��ms5@�5�74:�#:so,:��74_�#4��p�&}�p�q�s
a]U�7r�fft�ߋ1�6���v10��+fv_�j��0�Qk�����'�c���*a/h�;�����o0�	��&���p���t"M���o3Γ�������("x�1Ji>0Gң-����Ч�g����	�-�x��m�v'����"ã���j��-�\D��6�d�e���z�rؿ��Pʂ���d�oj�+<�R��D��m��記γ�a�;_�`C���)X,H���f`g���;ᆕ�H�C���ЏM�
���-��7�y�i:$��XR����"���sX��Q�V#z�v���������Q+<��Vg�;�+_唢���|[s�����(M,	��ؽK��n�9��E���eFkYb�`1��UK���gnv"Hv�QzHi��}O�U�H@��ƽu+t��Jf�)�Y/�j�:����-���1���6ʿ>O��뮫�b�<@~A�4e�,;mK�)����m�(�pˌ2J@.]A��S���J Y�)�[h�y���ع��O���������a�|���rA�``�T3uS��Nd�!jl(�5��)����������,L�M�l3I>������L���H�Ⱦ���hDFd��|i|�U�F�� �ǀK��tQ��8jF׉G���aG�:0�4ڿ*\y��?vp�ʵn��\ �z% ����I��o�REh�,��u��w	ve=�l�q� b�~|՗�Ṵr\��,9�W�o_��,<�i���B�@��R!�H��	 ��D��朏�����Ը1WP}�.<.q�;P�(�R��J�T�7Ī������<�"Τ}q��Z̶�]�ղ7:s.�n����c���9�n<
��a��l�#�[9�c`jr\bo����0R:���B�Q ���-���ۖ>ܰ�-��?m���%ȸ�z%#�X[�4<D�'�}����FJ�zU�E��]�N8hc�e�Y��I�9/�1iZ.�����.��hp�Ǌ�i(���	��d̗��蘋�eH��'�s��}$�%$	Q�
�14���p�ߤ���SJ� �2�ʊG=Eݯ�!ԣ�Ӌ�(��1���(���LV�-:��~���;��MˬٞN���i�A�s
w��&���R��' g�`�)9�����x��O8a�U@�]+�aɼ��x?��P8��D��}��pí^��z@6�d���E8�$w�G��������X�ZnQ?�*�_���j�,C���
����y���dfQ*����_/�54�B�%J�i����r=�G��m��Љ~kȕ��� ^��_�fOuOV�⣀�����-��=<�ad���k�E�O9���sL@AH�W��������K�-2!L^?����x����H}���DAզ�%k<�(�tB�d�7h��%d���'�g�>/v��%�E�lZ�Ƈ��U8��Id�����Lь���o������ַJ�ܪ�a�BP���	^�c�T}-�n�f��߄�t5>���
�!�:8Fg��r�<��F�/k��Sx>�DÔp��0e��x��R���e�J�G@<_Q���3�1Yvx���,�$kD�e&���K�@�5�g���0b�C�?8�{G�9�E�p��f�\UM7���t/�Q�s�ޜ�-���2Td�/�'(Y����w�ഴ+�^�[��T��<iM�5�ʧ�Oׄ4Ӈ`z-T�?���O�)�t=��칒�8]�ĥ��Cc��Eb,����g��*��W�T�j�5��[�W��� ���/�wR�q9�8}͊�>_���@��]�g�,�Ja�>�����P�B#���pp_tX5=�+`6��T9!�v�+G7��z$E�!��[�rKy���:D�]a��ЗM5���
��\�h��F���n��<�^��,_ކ Ѻ9��5�Q��ڐ�����Q�j� Y]�A���0/Ĩ�ӏ�b��4�>E���8���=inȮ��`��������z�<��[��#X��&��3��6�m?\�i��B�6�!�rbT����.��4<�9�ǎ���3�?�������ZZ(�8�"��h���.BN�iL.�zD&�-jo�Atv߶��:?�x&:U8f�����x�'�$��حB�R�����j�ի/�Z��łj?p*G|��������0�,-~�A�g)ZI<�f?N8fNaTE�Er����4	v5��Ue�R2m���mY��ˣ��k㲝��D��7R�k'��(�h�fP}a�.(����~�5�����F	�eJp)ۯ���hO��
Rܤ�>������bިo�_�p�ny��C��,��us2�eWP/6���1�\�����Ɯ���.|� �S۟Z�}Y�b�ѝ��L:)��1��l(��T���n�B�gJ��a�{��4�[#���A�A��ҹ���1b��T��M#c��P�-[��aLvcp����������j��|���I-���
]�� �\�Nhv��)��z76v_�tx��Q%Ϸ����8*�5�$�=���zٌa��I�nBΑ��7��᫈��V���]�4���B��|y�2� >���ʲ���6��LL�޲�J��,��:��  �)�S�Ro4�%�iy�g�q���~�)q!\�Z�a�*�SjGV�\[MU�ցP7B��8�ط0���{�Ǚ�S�|�VW��!�=��st�QHQ1:~"�]�kV�p��� �`��X%�#-I�+�h-�d�x�ve��iZ��q(���I{��Cqq2�^�Z��D"K힓�T��� �.��ܦ�!@�?Ls��Ρ&|��"K��N��y�hD�*x��D�2\d�\�.C����x�,��ݷ��:���B�v0\b�h��ym��%�s@)���G|<��������;B�p~{�T�b�ju���vI ����)�9bfB8�Uh�v=��z����ĐE��a���j��z�������T16��'�7���^�QN����gaB����>�C��Xu��0H����*�VU�ڡ>����o����-PC0�|Z���9�Lq�ES�l�Q([�H���
����@��s@ܘNU�i1��qy�l|���er�#�i�c��*���63`'eV�+���t�0Y�_����r���܁�[�͕(��� �i�YI=q4���ޭ���T�%̸r�m��:�1EM��&�+�ē%s����+�#���l��*:���2�\gP���:�Z�F4����OW���do�`��W�-����U����]Yޒ��౭E�/q2���(Bi��DtZ`���ALf+Ʈ��ipY.��_�D�r'�J��|T�&D ?���!�$��ԎŪ��I!��w'��!<zO��F��&S���E�|;c�JO���8
}M�u�]J<Uia�/o�%{����A!�J;�r�bJ5�F:,�H��;�n!!��63���}�8��`3�_77v�{�6u{�)�st�ƒe]�0P�n �@��k�/,$ZW��z��*lu��T�?N�m�fT�en�����uܔ�8I�N�ɳ�C��,�<�v�?r��'}�����WI�nQsf�	
�3�m,�,{D%��w����\-�|��m�
��m��E,,ӟp�`�s��"T8���%p'�n��F���(ɜZ&�`Ky�j�ug�3�g�.0�A��K�cca��}+è�� =��S7��H����=����j������E ���)�����g&�����L�V�1��E_'��&M.���A�v�ErF���8x��yU� k7C�ɢ���'�=6��Y��+ ����H��������dǰwiH���F�Z�V��{Dۦ�,�}	m\��2JҶ�m'E�\��l�X�4��5�B�o!0����s���̡���uZ\s%�� ���YZ��f`T�.����] N�_�Ů��&K��ĺ���nK%U��X>\��+�DY~{�囲ʧ�yQHt���=��5W�H�3ڔ�v��|FP�t1�=�G�b�Z-��{+;`m�1��#��Yl�,�dUTĝ3A5b��*��ހ����,ѵ#w�q�\��[c���8H�h�Hv�tU��~���*/�=�a�6Q(ꌙ����Wmzb:*�1�����K!��,��c���$,�7>T�E���8�a�[��%����C˷�ҁ���+�4A����!O  ��@���;Pf�b�o)����)���Cb�K��u�X�l�Y�n�c3�|����Qu���r���eV�
M
��b���g���������Eؙ2G��M7���͂��+�o8d[b;�����ò=zF�K��Ϗ>;������u.������� Q��k_�Y��������U� MȖ(!T݌�����>;��9t�����;�"QRZ1��W�*Q��p�v�JU��޴���\��J)�?�^8$8X:5��i�&�Tg�0B�	) 0`YҌ�WGN�8:���f�7�Ӳ�*agZ�B�V !���.;g��7�:�T5�~�6��?��1f��3�>��А�	_��.��Oxz�eD��h���)#���'���F�zήn��V���f����D >���.�h2A�0���;|J�-��b3n�!�B=RxC�k��-t�I������j\�\R�˷�O7W�Ӷ�M��tg�ۅ��4�x�F�h!U#�&��[��^s.�/�\�ѐX���SUZ�{O�&Q��,L��*��;���z̪Y@G�a�N�(�U� ���}rXp|�kSk�ͮ��CI=��K�wQ 3�3�������Cl��9 �������*���HG#��*!��&�3�g��oj*L����S�\n��#��B�b'��9�C���p�T�w�pܐc����@}�Ҿ2�������P�ɗT[¡(�\��|���H:�=��)�)I��Ե�q8z|f�I��>zd�ܝ�*��*�1Q��4l��^c�^M��JB�&;V?��)g���`�  ��f=�2G�Y��t�<N���Ew����ozM��; >1v/AR��0��j���(E�xæy�*�b���ٍ$V�	WZ׎0�[C�,؂�:����6�!=&�-]�}ӕ��N���/D��~�%���nmu�0�~3�sw�tȪ�O��+�س��6��-���in�*q|8���i�%�@����ȸSEXm~SM�7�>�y���rGk��*>�ț���_)կ���6�Z$�y�T�*�� ���6�K�B%N�f�%�øk�YO��}��{���}{;oA���+St�����,�r�dr�n=�"2��+�Q`�6�M^�@��cX�G���N\�L[1�%� <��A�R��Q�k��3؆�rC�O��S�%1^d��$@��pjȈ�*��Նm����U�B��Y+:cA�U/ǝ)ݗY���¨��}U�-0 &�(�AF���N@d
��E�C\�X���������e��.G����:\f��9w�^�)[o�E�_��WӁ+��h�w]/0Zyq_.�#W*b��2XAsٗ>u���۵�;L���9	��R�dpđ+�Я�찚n_>a���m��é@�ߩ*����En�>k���y	����.dݠ�!t/���R8�9� �E��.�{����>�I�bʰa�7�6�W��<��4�ь�0���M��m]<�Fs��'�I��ѣ���ӹ��cP.��W���P�]	O�;SIt�p�..��P�A Ȍ�¼	���U���<���kת�~+�CKȁ��7�c��\8�ݏ$�؉!ā(�PE��H%/�����"�����] +=b<TAghat��ы+�X�oX��/����=M U�y�ͨ�svt�A�Rŗ��ޤύ�<r,AtV��}��Fh��1$yr�l�H��E-]�KkMODa���y���^�Ф?_͏?-������o���	������P~	�z
��qmO�M�*�p�e�1@�,mO)��t�<?���ca��d��Q%D����y`�)0����8�H��&	eqU�Ӓ��!>hv�*��Ƽc��Gb ��5��>Yl#/��|�����-l(]��2O�b����	��Z:��?�R��llz��3 /�q�:+],���$��1_�6��<�Z}43ѰRn֮,ڀ&�!�r�)���(��^��f� )�xɀ�&Ap�D�Ѐ�Fr>�V��������>gXO���h�sy�̞31N���qL�LV0�)��:��YI���Y��4�鍳ǈ��N#�ǹ�x/-�����$ڍ$�]N�ta���x�K�a7��V��p㊱���
�۱�q@2RJ>����O��췸�1f;�P���GE��XgE�������`��:.�m��MY�7��3A��p���w��ܙ	����V$K	d�1�x{s�K��	��G]Xk�#����s�q9RH��oer���~'�����]��JJ�W��G���
�e�[69"~Κ�m���'�aYDAK���O���Ke���2X��{��rw�����y�f�t�Y`�S�l��e!�G}��]8�,�oE�!����[�P'`F���cM�uHd�v����5���X��4�5����G	0��i&OC�(g��|��}EB�5n��'w*W�9�5~��'�]ۡ"���$FƋ=�Dߍ����8���|#�H�g�Ȧh�%Ԟ@����<��a�W�2�&cD�砫'�1X�:=S
(��ё��s��=�������e0�
15}2�D��z�o�A�OFɺ;Mɚ�����ҿ��'H��TE��:�a�n����ǫP��u@�@�&�qZ���f<W�ˋ�'N�(Gl>��d��F���񂪖>_w/@�mF���T�����MC1�'y��Jӵ�t�R�~�\gw�imʵ�P%3�A(5dG�͌�����9�$M�3SR����.��4����Vִ�c�R��I��x�a�+�9�m�%R�RY��4��� V�:�zW�fR|Sh%��!��)��I6h��5�%҃��q�`��^�GA��Ub͡ڏ 4�i��]�p���RфMCf�C��M�bE�M�iH^���çx�
��Du����^Δ8���O�m��o^�B�+b�9Ǽ���ɬ-��2�ZI�&�/�)����2��:;M�h��,�\�Z��tw�=$-'�ej�&�M�$OdW�m����i�܂0[ZX���vg�)Wن��A��UGy(=�C�*4}H�
Wks	����;APۨC�g��Q��J�Y(��g�{m4W�]���)�����<�,�y��KR#'��4pfa}�����94+M��Rn��ۣ(+������~ncTq���� �X��B�`��l}P6��b��44�ߺ��G��;(R,u!O��n�:��G/�߫�떚uCQ��2[�K�y ��J��M���}�l��Ɣ��6NX�x�4*�N�Pnr��lck�rձܩF;���nu���&ᠢ�&I��\rSM{*q릙{��-�g�ٶ�F�¹ �F��T��$�����G>�qP���rl$1���lQ��l/�0�7���R���wb?eV+䧈D[(nJ���c.U�$����o{ϑ8�'Z���W@T!���o1��N�z��W�'�,&_c!��o_�"I�(~������M�pIX�� �;��f���1�ҳ�<}Z����ztq�d 4B�|N��\����Wz!��V;aɄ2:��p�MtXs>�����6N&�7n:Z�X_����"����3>(\�Y#w.�L
�O�'�g8i��uC��|�?Q�*5�<q��m�A���K#�LNF���z��LX5��s0?*4i�E��S7���G"���6`���(\��(�����V'�V�3�W	;��Ӎ7�>^�������3ob�M 1Ɍq�d7;Pb �Ξ[a n�z���,0}谿^Z�}��*��˅_�(�7B��AJb����S<�� P��� ��5�Տ�X�G�R���Ƶ.ifp؛K�,��6v \l��Y�
��B��W]Y���M)�@#91��PiX��̗Z�dC��RPf���*�[�p�U߅GN����;kk"o�&{Az�!eT=���	�U!�Eݶ��w�/��j8@8��/(��p�*ec���{7S�K��\���r���}�\�8���O?�g�gLg�^�^�l�=���R-��R�5lࢻ7,��/�YobNZ]%�npCnȯ�Wˁ�n����Ӑy`Z��뿕�!�����wuR��
��b�2JG�&��%�7���d�Z���ܕ�y�̵U��]���FQ}��jό�!�Sx�>�lU��o6��~آ�;�X��@��W�qy<�k�L�K��_{$�+V��ZN�A�Z�����d	w�8�5x�3�\���L���a2�y��/��b/īe���&���ҿ]ܒ Zn�,0#�>����@"��!��׋�3OEw.��T����I��j^2Ԋ��ʾrs�ࠍ��d�1�G"�ռ�k�A$u�L����U&x�]m�gyf������S 2�s��#�R�׋gx��Ȼ/����0,[�w�Wv�i���Ie褭��Z)g��C�N
��YXN��XU��#U�����[|��bǈ"��8���'�2.����+W�F�F��2�hh�Y�Lv\c���|��
��%����q��+�(w�Z	�BI������C�]<�{�7?*��h((Ɏ�ud.����,}����}s��T�O�Q\�[�f�g90��J=[���ZU��[z����M%8b�+w2%(��v�E�yK�ũ�Z����� ��f��2bf����S�Ϡ�>�y�
cX`���R�l����N=v�s�R�"MD�n{����95��Żm�g^�F,����
Q�z��z`7J�eSy�bY��x�������o��r�k+梷//�>�C���7,���{tp��UvA,�7%t�_H����*���Y����[�ec�K繑@#RyEz,I�㕊�e2����d��W��AU\0��,N�l�8�ͣTe9�N?1@(�������\�es*��Р3�+׿��' c���������Djwn&���r�\���Tv"���-����oTXC�<�eW9L��1�Z�O��ђ3.c��OAH���3C�) �6�~�Rs�3�1��y�P��"m(�.�-["��,�ꆂRF �~�jbb[2��Ȑ��L:.�_)��cW����,��Lf�^��T�Bq��ޭM��KFڻ�q
��pA�����s� Lxz�#
�jZ�8iC��,R ��$^M�q��⢻�J�;�q"��x�b��͚B���j��x?q'��?Kǡ�VS�հ&u���nQm��w3��i��9���[�Ob H$�� �1��ϡ7�&K�=�N�$��J��EM�����t��k��0���v�k1�u=���@�@��\BGT�:݋Me���ڡS�w."�|�3�=�*���TE�otA����+fM����kz 6j�2��1NL�JK.fۅ:(h��`��7�?�S�������a&~ؒ�sy�����s�+�������V��K�!A%f�V%�%�hu]��/�
�h�"��:�ԕA�
�F)��b��R�o��f�������S�ʪB�;�]�����(�Ҁb=Z��q�4��e��d핡j��F����MW�Z�6w���C���'C�b�f����{�h�A'`U#�?��m���{���6!c��ǱN� u6	sjV0�Ku�������qb�Zʶ2[q�i眬�[��b�mǘ��q�b�Ҝ��E(íl%�o�L��ڪ7H�xn��:�X�Q���Oi�����y���߉/J�-@f
���o�t�f+`x�^�'�4s�\{����ܼ/!�E��[�����W\)Q��(��	[r���X����7ж(�ߪ���)	�cy_ȳ4i��g��H�����o����P�~\�+^*�/��~���e�o�����x�Q�f�?��}_�)V$-��h7�d��<z^=?$ì.�/�1!f��o��˞�Ύ�I���[�q1������že�w��\�[�/!X	�_�R17_ͦ�1� �·1x�o\�B7��5<@����3R��ٓ\X�UC{}\�b��ǗJ%A�@��w5���� jd|];�t'PJ"s~��gg!��X����[��5��Ñ���O���`ݴ��BxF���c���D���X<�U� �l��J��v��m �����)R�ɝ03�k�i����-�L��!:�_[_gbr��uRu�)���#�*M�>~P?�)��z�A�6r{�۸na�ڏ.���:����s7�:zڎI��G�9�ۛ���?��� �.I��7�7�+9M`ľ!�Z�)���6		A�RrI�ڟFr��Y��e3URؒ�T穊.F::���v_��B�g8�T�Q���
r!?L.�p�+_��vc����"��#�&E�� lJe{6��[L���Y./~��֒�?��>��lW��n՟�lU�͂
��)�3�O�&�q��+Urp1{�6��U��C W�=��n:��c�����;��H~�"?���W�y���y�x�y���AL�K��L�y� �=�>'�ouh��L��͟"��4ǈ��!	P��t����c)��/p�L�3���f���.�OJp�܂ܤ4���=�!TU]��'�h���e
�y�?c�;���>�����h��ϏD��
4�g�t�G�oZX% �>�_��TW����lY��]�V8�1U�h%�{�3�܅��ΩflB�wWF�N���0N�C�ԫ�tP��)o^�L�vY�����f���V@���QI!p��ӳCD�n��S���>�t�)f�y��{#��<Nz��N�9S�VdSՄ�Nl�|;�gv�͊��=-�x{㿖���!8�.;���J�!h�UB�m�C|�΢�(S&iU�/��Ҷ����4آsʄ�r�3B��"��v������M�@�E�QA�}T���!��*��x��-�p�f;8�=;��{!�6˾���b�H/c�<���E�RCp?ɩ��C�Ώ�
&�XQm#뀣�� ��Z&�蜽"�����d���n_P����6x�*~���a�X��$� w����C��m�,�]�
B5oU��p��=>���<������M%V�c�Bwbq���r.��mihjh�b��s���D��o�{����޵�
�ހEO�aB��p�n׹�<���)*y�K��ý���U�"_�5"�0���2�(�?����hj�����c��_�B��Z��:�0��#�x��J�&U��*�ąv?$�^��,1� ����];�C�p��#��X���Lk���@����M`���_��=v� �}��}�̏6E�-���S�-y> �$�%�a���3�l]F�x����^p@XE��| �<�w�̅ф.H�o6lHH��[͏���a.�*����f�"i���b���U�ᾔ
�y�mQ9�4y�������*|�'���N����(��xk�Q-��^`��XT-�Տ++�[H�ē�X��J������5Fod�C�H��q�A�yR#B)�����^����Y��<�]5rU~+\�"�HY4�u1�v'�(�Qѡ>T�k��nm��bgwoo��v����,���2gP��}K��tZkM�Y�oo��L����<b1yC����Q[��4�����8<�Sױ�y��'
���bW�O2鼽6�_��˻��{O��ABL���y�*L��;	��d�r�2|A9x[ѳ�P�6"N�-�|�"2�e�<�0����IUO�H����>r|-��$�i�+EټV��J<ل�6Z��诊����4�u䓧�5�jw����� ����fX��A���y�ӖE��r�����$�� ����6�3s,�6?�9���C�;�&��ћ�1�T�y|C�"���au-/s��`�"�v~��{��Iͩh ��q��X��=8�I�;v���?�VP���B�u��,ȁ���H풋�q��l>������s��M� �XO��&�t~��y���2���Ӆ�kv���y�t]	�M@���x���	'��<6�蟽����<<����٫��˖�2[��+j\9��+<�LOO��U�ˑ�z?:�����9CN2;��ʛ��Q�5a����ݺd�Pp����?!,�_�]���F�a���Z��͖�%�/�bg9��2{�a��D�[~',̖� u�l��!�D�RL�zE�N��rM�����C���İ�̅�3j��}��N�cz�:�Mដ��["�	�s�w.~=
= R�c��̬���M~�#��{�u*:R�/9�46�!��W�҄�M
!����Uٜ{j뀅wM5��}鸩7)�n�0��TH��G��9���$!%�Z�Z�[h�∞�
���?��o�2��E�4>���NQ�3E3.�?ZS'�!�>a����-�!�3d7�����I�h�H��b�V�F�Y���Gեo����"k����iH���
��?,)f�u/d˳�k�AM�>���̧� �@Q\<��/t��?�]/#�|�P��|���Z:�������I��l'��[��^��v������