��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}�������B�`ה��u��&Z��d���d�~��h�a�h�f��%��+�E?L���ɫR�P�>�Of��fV�U#ʴ�I{f�0�H�ԕ����%p@O�P�k�k\=ۦ�}1�����D"�������6��3�<�ev���Z:���r��V'��y�Ti%_U�Yb~ޛ�����2�&�Bď��4������9>�&����?��y<������Σ�*ZtO����~��I��h7~-��,4�Ή���� �ט�0<�(U~}r,�	k��2G�w���?�K�s��R��_6>R�"A�Z=�9�C��>������u|��ق �I���Z�l��羿B9����7���V�7��=����D7NM�����b�9u*��aIJ�c#��ɷ�T��Ǌ���0��e�!�9�Cz|�[���y�-T4��;��h�c�P��$�?0G����+W�e�(Јc�Td+}yx��@(�Q�8X'�gXH�});�r�Bo�4}jv%�}�TT��-y%��[�]�|$�1��`G�k�MQF�g�����9H��[��1�|�H⌂n��,��\?���%O��� y�v���F8�����'9��|���槈>��#����kԽ��*AIZ���E�Y���Bk���1,W������o��^OZ�S��55�#�<��95�.Y$O`�N��ǎb<�b��s��g@jh����љ"Gk�Dc��p���@9��p��0$:�ztB9jX��t,� :,s�����L�`�4�֌j�5���Ɗ�ꪵ$-�x�3?|��~P?��ҽm:N���U�+�)�0,j��_��bL���s�ƭOdn4��ŕ��95�ĭ.�G���gg��l�r4���8q�[�6����4�×?J�PI�MR%�e~m8� �ނ�'��I��J�� ���D�EZC��?+�pO����V�!���GéV2v"vRG$�Km2�ڻ㞥��wg@Ѧ�͞q;�>���{��
���[.S����ޣ~�eT b�L˻��U=����y���Ƚ���$��!{�	�-+.=�8�x �v�pei1e�����nx�5vL�9~T���
<��+(��-�/�u�z�(����!cn"1�lL��SZ	)
�+�]����FPov�|���-УO䭄/�b?m�f]ӟ�|�	�E?:Q�҇�!�vx�K���|å䲟����Un��u1���6W��7��0�h3�߸89،0�0���Ur����c�[�2���B�y-P=:-{�`�q�1"��r�eܵ���c ��>��!�"dY~����J�PR[.U��������d�\��[���ݼc}OT���(L'WŽ�w����ڳ9ZkpU�2��@9ھL�W�Js�Nj�m'�vG˳.�QTv9�"�"ڣ�9@=�i�o'Mw�0��־IJ�H�"zs3:���z� H[�J�����f�V+�i���&`�R.*j��8�w��;�ְ�w��9=*0�)rx�~�6�f#S�w���@u��@^��"���ɫ'��d���X�}硥��f`����:حb�K�^��n�Ոk���rq_�$�������*T�J��8K�ܣ)o���lӃ���ݍ��F�yc��B����W��E2�n��<m5؜������em���^��[D�d�J�f���T�4�cJS��*h��{�	 ��ko��������!�����s���xu��#]���"�b.ů�iW{A��Vw%:�"���碵��H� ��&�X�������� ���
��Rs����1ݥ���_��h����Q��o_�]����!i/
f�4I�,!��57�%�y�k��~�&8K�~��x9(h�w������6���b?�W�X��[T��#�u{��2O�u"@�7��J�ɐU��N����eg�4�z�JƼ��{��_�c8�D�W��r�����Jn��!�������Iӷ�W��G-�xS�̩NY���K�U�5����oG��Yy|��R|�5���r 7(�7'l����J@\�f�ݛŜF��Q2N���Q��y�e��#�%�*�^���h�`&��rv��i��1^��}����4&/}����,[6o���n8�;��e(>�z)_�č)m	�=�#V*�u~��`z�#w�H�@�nv�7�W�5/v��G��Ö�� ��He��ƐMe,U&2�?p� �PK�)tJzԏ�2dUG?�55�ǇGf4�:�D�R/�}J|�o.���?	� %H+�H�+F�X�]w��Fy�y�\V;�BN]�4\��AO+r�����^��<c|,��A�&����d�3b����ը$�D�k��ͥ\�+��j�_]F]Yў�''���G������ز�WW�*1�'$����i������D��|�^;w�1Q��A�
�>\����GC���Ls?H��zܝ�1��p!����[�U�D�h����<�x~���`� ���p4q�nlQ��eJ� 4��W�m��DԎ�
WC6�}N�1�3KdNd�]_+�F '��s�z����9)��n���l�hdr �9�:��<�F�W����A�����iBm�-Ұk�j��~�^��QVw�������J�4T���s���u����d��N�h���#ǯaҚW�8(�ݲy��� ������bF�a9��~)z��[Ǭ	/!�B�;X�
�װ��{��������Fy�ڰ��+1+�"�a .�IBr������E�^\�h�P+����4.�f�|O���xKZvx����%�\m��dWD}F�Ʌ+�w@I��d�;�he�T�׈VcB�9G���Y��)�ׅ��ji�t*ciq�	<������I��E��1R8�=J�i@���_�.�/�J�@J�)�a�R��~J����3'/��4���֩9|^�G�@�wS�m�������亹����������SSI��*��R�Ŵ�bR�,�%�*������P^��v s�~a�n�-kV`�k�,��Ú�[��41ۖ8#�`�ϜчR`c������!����J�]k<0�V8t�.��-HlS�Q-�nS�������F�n�pd�"t"��	���q��&-�9A)a	I�P��Jl�ɽ/[u9O}���!$��3!�z�{(am���_�.di,� 5CɁa�A�]�}�9��i�s�����&q��0��'��(��~-.'�F��xb^�峫�|A<ˠb�o�8����켛>��5��Ur�6��s��$-O��W^��V��J��8�y�ԡ��ǚ
�D_v��Q�W��0y-?&��h'Q2�&��ф�G)� ���������(%!#NT4��-ߖ_�զ�&5<���v*�#IL��D��{wA&C��ڑr8|,B�KNDf�On�E���цl��uֻ	~K&~�$ܕ���F�H�QoP���}Kj�WgX8"�������p�E�#<RQ37]���ʾʝ����kjT����G�V�Ê��rX�g�����NV,������{�~x2T��=i���y!uC��0�|�m�$���M5�g')g��l._-�f3=V�M<��V�-�9�49�B�c>?�ޫ�����5y���;���CuJ��&l�i��td���Ya A5~�P�5nE�jX���@�.�]w�z��[�4�(>�쳕�w	�ă��`�X8��R|��h}d>'��~=��݆��j�8�rB�o	�D�V��M�Pt��XG��7���5���a�-G�7�*g�.�I�B`Ȼ�����B6vXַ�jI�Op16h�k�?TBL�H@n�n+J�O���B�=	����h�Л%C_D�;�W|&��2�ʤ fb�B�����l�@E��8z�to;ʃM�l��I�z.���+�lph�=.����V,f�Z���|7j!a�T��Z����� ~?�i$so+VT��&�i���S�
w�H���n�o�g�GC������}���h-��ů�݇㑠!������v�3񩾍�1jQ`9 s5�2�:�K�"����x�B�H��ۉ�Og�wg=eu�(g��M�NG�BYj���@�U,i(����A{;�k��'%�����xC����)�E7G?}�A�`ŉ��×1**g��n��&��������ʲ�]�լnӁ��U``-
��{R�xX?�n,p���^�c�K�|���2�Nљ��������-}���p�B�5"��I1�V9�U��7����`H��8�Q��!:���R}7�49����O���%+1A�$3j^�����t#��麶�)µ|��ũԐ�6?��$*>J�XZ���@V�pּ�mO0h����).��]�J�ꉕ�o5q�-F +,��������Z�� ����c2L�aO���T6���è �~߿�/qa�?(/6uc^Rѵ��E>ph�|ApM��&+�n?:i�̼���"���X�ү<�׃�ׁ�d��L.K������r�N^���%��n��e�b���T�./U�����ʷ��:4?�m>�ցdfO����QS��7&�.@�s���>ڶ�َ4 ���_����V;�����z	.�L�#�g�H.��G���QE�se���@�5q�@����\7�1e_��*�b!|FE��&�zu�72k��Jy����^�U-%P��	�=�����T3*��&%��2_�ڳ��BWȫu~�d�B
y��i�~+�2<P
Y�D��\<�x���