��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�P�UL	�s���U�P��� 9B4�(*��kC>S��k	:����4���pqo�.o�zI��rjFF�/���j ����tp�|���!*S:ԣ��4�7�L��J�s�{+:` �,N`A�DX.�sJ���*�B�-�:��K"9~}$�"7Q䦮��}��mH5[e���'T?�;�]��-~y[9������k_�2�V�{[c	���=���-X���<�)o�G����]σ��dy�v']�;���<Ir��J��1���$���8ă�T�;8)m�T�qh�>��LJn�ݐ���U����j�NPk��f�/��h��Ow��c"��_\��%ř��s��l��KW�a�L��+�ţ [���I|/�siu0�̰��F�
�:�U�b�4��M$��.�n�ْ����mي=�^¿��ݩ�`��_엔$9Urzfl����4�s��ϯ�բ�.�DHL��%�i�v��+���[�	�?أ��!�U���x���*(��!H������oYV��J
�:�@�;y��w
~�w�`b��1ZY�l�E��9#w�_��@8�����e I/i�ȿX��z�M7��5vm`�OZ�2¼�ep�,sw馗+�s���}����0�
�$xlU�@�����u���G4�7T���6�c���|��lw�k�}�����Nk�IbR^�K�~��$�c���0�IC���x�?���w�����y�Z�Q�ΐp+r51���oBbkJ�8�� 	���)�~��v�qL�8G�r2�d<�7�C��ҙ#�/x�J�֖]�A����L��*^��������P�y�l��s4L�(�!Ҏ���a!���<#��_����2y�z���*�s���O�ʒ�.azTdzJW�LJ�f;k�d̈́]h�e=�h�s����VQ#;���[bt�Â�B�m��>���iL- .��� O���	��e����	"��ni��A: �O n���RmO���A��N�-����tZӿ�:o��Ϡ�{������[� �x���K�F
;�N�̷|��S�D)�J�&�����#R�N��i_W4{P�!�4��|����*�H�g���g=�l��O��e�)�n���� ͞�Q�yV�^���R]��K}���4���:&���Mw:�#�R��)�2V��.T1R���H�j�ޣ\IP��x�I�:î�"����M�D�4��������<��AȌ$�J�L���YX�d��.��F	��r%�
���7�N E�Ճ�2��ލ��Bzr�m�ӌ-�)\�}4��W�
�xl9�0�t���d
�ԛ�-��5�q�z��ℎ5h0��x��ǣ>i������%P}�\���Yמ�l�.��?�	<Y٤{�? ��ݾ�6L�^w2��o~�\RT;�6������U-|U	-��t�X"��PC}׀�j��9%|<�v(v���/�j�j��4�;���i��`�pb�%�(��ud�mc�gX���J�
|��<���d���L#�S(SpS��^��q��
��<����n�X>`nPȴ�QLc%:(����]�u����1�ipXo}(�,�XX;۱~��C^a���U�� h�M8`R&ƨV^�.{VZ�y����bFK��O�W�:��w�����=�7�r����a����&�T��;���`.(��l��1��?7�L0�RB`oMD*]ͺV�-_3���{G2P��Q1�yN
���6��w�Z�E
.:G(�yv�Cm{��HK`]����?>�h���3�4���c#P����CɱpA�H�׬�}~"5���;@aY�>����]��w�D�^���w��~ˀ������U/VV��S�@-|�HպAwfI�Q,1�����8[�b�IJA7�D^a�xc��ĨӘ�tU��?U�5��`/�(<�2��	�Ӳ��*	��|�/�%�y��}���*�0�Y���nS۪����;�ST���,F՛pm���7���8
N��6��#Z���g�ߞ�Ӡ�Y���7�L��3�o���r�ibJ|k)����4۶(p�w��zcY�����N�F�#p���-��8�#�����X^$�y̖ ʀ�UI��2[�M�xY[o��a�w�U�d4m!s*�t��W�Ld^U7��3��ԗZ��t`�Y��� ��ݶ�$$�I��;	t6���r6ɚ]�ֲ�eP.G&$��Zp%.�o����Ӵ_����+��WJ�l��,��I��Aؘl��i�G���>W�gK��TZ���`��Q��� 9�������T��$����<��?v�'��g�D\�/���&��;nxP���'=��U����6
I��VSb�
�(������F:�/m��Y"��S�����R�lN�0���l�R>�?6�̎���|swn�_��!�>!9��m'�~s���<�7[�o[�o���ψ�2�V���֤
v�6����\����&���X��Ӥ*]cz���=���9�o�P���M#�^p>â�CU����!z�L�s��`ЦL��X?g�����hϗKjЮ�E��@���D6� %�oK*g�*e߮L�����DW��:%\��snp'(���������}���t�mj�F����-$���x��Q�i�
 uqwP+9?�������e+��u^����TyK$�����t�WGo�����.ə:tL7gm��0��9۽�5X"Ɲ[\i�N�6|����\7���(��ş!�gn�O+���z����=R�߸�|.R��l�S�.{���3ʬ&��mP�sf��
P�<�SmA�����΋=wf��@_�X4�ZB;���5b�tVM���L&֮qJ)�wT�9V����R��zk��q����:� Ԟ���ɽ�	��,5o��k|cݙ��mf�b'G�f6M~���jM'�=�m���r�Ymn�x_��t������SY�n�])"r�"�.���jL�	�]��I���N2Ab�(]����"�)������ ��;��ˇ���"[���8�nڈm755��d��)�������K
|N��`�<p��IѾ��Yt�MV�?���mf⯓��q�е��sXuYcu��/���I��^������F��l͑��	���K}�x�>L��%;��f����JaO[�[�[�|@���]����X�~��O�G�>�����Ұ�D�)�*9���Ղ�|BViz;�pKFi?���4�F����S�Ŋ���4b�ӌp癩���J�GEC����D����K� �Iv��3�0�T�ƂȢ��&�,����5ts�Y��k�װ�H{��;z���I*�������!���7V����ֱ�m�"Rmħ��8��(h���C�n;W��C_�jz�t����4�a7ؤ�Y�4n
ݤ�e��4
l�[���H���j2�	���؞�6�8d�0�Z.#����.q	��t�3A�X
��{�&��2% ~�6� ��%RJ[62n@��CS�$�L�N�D+��W�	��(
T�b�H/乖�����ѳ�+Hfz"?��eFU4��(�K,���5Uy�8��(*�<k[^"�g�3
W-�������Q�&���{��ǧ� ������a�bS��	��k>�US�D��&~q>�ǈ��u��Md˵Y�k$"j ��u�n+)f+C����G�v��FwD~Ų��K��!���Qe$
\Q^8K�)0s�<�E��1[f�BT̋V�kd�5#�|][8˳��[YѶG������bD����ED^Kv���q�G�e~���	 Np�PH�$Ѯ&��p��/?�����Xo8�ߠ+Uv�x�#&I�C�ۧs�����E��{[�Eɠ��S���(6����rh���}u#(����ƳNVa=�uv,H�K�2 \ٟ��J�2���:��p�%��� _՘�y����>`�����T]��飌���\�
$�
A����ת�m�s�F<�����2�8���E���Ӈ\��@2�-)��Q�胥(�ȠT�b�k����`�<��r�"A\w)�D�u*R��Cʑ��hR�>Ǣ�L� �^v�5�n������H�Ԙ<3% 3M�՛�oc<j��D���� ��=�vm�h�.�o��}(�9	k�7�� �UL�dD���2o�ߏ[al�� �D.;w��0\i�[ٟ����lh�"��@`�������ߒ�Ŝ#"g����>���I��`��rp񺎀Sq�X��U���8�ލ1�2�?��}ӂ�4P�!�IE��ח�I��k,��Fy~QK��L��zD�����w�?������Ve�`��`��k��j�Ҳ�C���]x$A����{Әg K�@�b�B�VT\����R��G�%��A�S��)r=�~_�����W����BD�|�"�X��t�.*��t�,��fR&��#%�#.��1]W��+�z��i9�|�=������_��{EtDƶ"H56��_M#P��ʅ��P��A_Ԛ�8G��s�ܞK�҈�������am_��+MM�:�Ѝ���ǭO.���b퀉�ޓ��3|��dWt��c����܌O��_����iÈg���n}̬ȑ�@z8��Ȧ�R��D{o�d��坩a^���û*��$����z�QK7UXvO��`I6.MS�`�C�w���o�A�R��&M���Ĉ�c��..1O��)����I����{�����~�=��r�&�h����5v�f�k�j�9�熏H��<����t2HG\9�k���e��〨����Tz�T��S�j�n���V� #tr���d��2&��l�J���j�/�����-'4l�s�O��1KĞ���|NfR!�-|�^��&?�������:���:&5ך�7!	����T��xw�#V�޵�.��S�V�us��
!c5c�!R���e~��Q#��89a5U�Ӧ���j˭)�?f|�s�E���C�`�I�X��AgL&ܴ54�I/��������Q���Z��J4��),jbS���N"i�v�u�ؓz�|O�?�%����A�蘴~��h�ex�Ky�Kq�K��s9�����/t�$�v@&F޵�����-���|~[���g4��^<{l	ɐ���.�؆�h��j��ŝBw�Q