��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�ףe��	�A`������I���;���a���^�]���O��oҎ�t�~��N0�=+�Xs��=3B�@�cT'���Ǖ,ç	�9��%�ْ�o�q��9�ˉJD���{��y���N�N.�qC�@Hv����7hk�ү�VpK�ξ�W+��6X�D���a����r��1�NBcV��sj�^}�%/�-u��s��D����&���-E �b�q�P�>��K��}���F����m=/1C�t�d�^��)�}����l�Cn�Ҵ]ţ�݁�'wR��ۤ@���7L^�G�G{��<���+&#�8��Zf�:ћ�'�C):8���Q�a����c~X���v�Ip��`���Md*.�m,HR�r�jw�an ����������_������7����g����yN2>��&�r�W����F��7O��ALc��k�b7�0�)���� e��b>��9�,Npys��Da)�ٚ�˛�����Y1��v@��{f+���1Ȕ�tI�1��SԼ�>}4���֨���9�T���ȴ��e�Z�Yw0�������Q�n�:�n_���Fg�{K�#���Ϋ�-;\T���?�cA��>H�@0��A~淂4Vl�]Q��*���@���*�]�h9!"�k:a�tC�Դ�$�v]���Px  �5Y[~ܟ�5-��{�-��F�iv�&�#%T�(�Qg��9Ӫ����nb�=���׬�I�"���)V�1 v�b� +k�%Xn���Dŉ��~ PNYT�YN�0-ۆ��#^��yb?��v�r�/�U|\����9R�0�s9�+0t�-��+G��]�=��<��yZ��9X�}go�W��/�j���'�h���(��.�4�/��z����w�W3_��!��i��ulRKD �2��n��WXU~J���F�vj�Ld�fG[}�'�h��,����ΜLf���35���批���ﲯw���I�f5������&��(9����Z{|��}�7���}<�ܟ
��n���0�!�o��y��F�$�f���L��N�������lz��8��L� ^j�'�)#�KskԿw��g֭��j��|�%�kc�N����ǹR��ɟH�eo�|^C�.j���/��~�:G�	�s�vW�¥j��uZ��.����bW���a�l�N�)��*����fî��2>Y�i��L�Q���Zd\++<�o��\��)H0�z�2��v��~��-h-�Z��0=��	
<Eٶ���(6(�Φ����T��R<v �Z�:t��QQ�n|����6Ϟ9���p�.��.u�-��}�����C��z8��f��Bs
p�9}�)����Ƌ�Z�����v��9�n�h���.!��ݫ�
\���<?��@�#=�X�ʿ߰���3�<?	����*�Y������-�Qe���s$Rn<w�It���+�7��j��V�՝];~b9f���JK�4���"��< ғ%��&�@�=����i$�]��x���bb�E��eD&wo����k�qb�̈́,/�	�|�܊o�{���/r�D��CA�ޫ�@0}�\kF����A8p26.&y�mn y5��M���`���5J;���w�V��̑���9k��q'n ��L�A���o�����+�#1n��	���^nz�_�qxI��)������G'/�o_�$��j�����h�D�Go�@�h��X���_�����[�oB��-Ґ)�S� �vT/��%�Q	���l���D��	�-P�����7AD2��
���͉����V�,��A�?Fǻa�j��5a����B��B�<<�e��������d�{��F�c�o6�l-�e6]�'ݫ.��K]�q/��͊9sx���Ș@8V3>D�bMhh+�ہ�6����K�;u�:ERzlbf�=���wo�Vp0&DW�M�Yn����&!�<<鳲�����V��r�)ݠ7�vjz���3�~C~}w�����D� ~��`�k��	�U���!u�B����$*������,mtl�G�t���S9�"�3H[��V�P���ɺ
��$���m|�AQ��Vۿ_ta-H�G��a $K�}?��,���)�b�m��b����/+٣(���0�(��ޠD�i�굊