��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a��S]/�k�q�&�S;�YX���L� �L0�4sI�1]���B^��}���N��P�k���]3�C�)�4�9�CJ�JS֐x����q˫��w��d�lQ��>^���RTZI֊N���@�3�����y�B�ǀˉE�{n�`5݂/�*� �W� z)�R����9Ƚ�����C�,<M���M_�B�<�Zju���F�?����+�hj�g@^(3pb�n��Z-�@�wm8w!n�����֔�;�Nw�/�������wU��!�)s�|m�2o��Q�-�VۘӀ��dM���k��#�b���g;m�`d7J�@5uر�� �т�a�	\}'�HT��:���!���L�t��<ӣ�mZ�Ԏ=S=���5D�"6�]t��p&� �Р�䴙�f5u�T��E[u˝�r��z4@����=��K﷋�aD���խ")c�B�x1�E�7v�-�h3��JҮ2�^�)@�����k9��c��˚����@�����/�2��̀rz,6,D-^�Ӗ�@$q3&,��虄/�N��$d�3�� ��t���K�j���݁�:`��ұ@�{�Dt���j%�@����6�8ζ����wT.��UT� ���ÁJDM����m}��ϡ_v�o�O���)*<��TW�]H�t���J���1J0�}�
��pu2�}�>�C�tGm*�����9X%�u�3}����W6�Џ�7L(��|���f(��T%�!�����捭?���X�G<ܵ$1�y�4��J�DIRsh�!��1;�K� " �Й}DL�:ѥk�S���V?�Ӌ�v<�\W1������ZLq9�N�h����ͥ��admO{
����DM��t�f��?^�|��ښ��Z���桇x�B����JET�c��=�P���"�3dm�2�wD`�H�������3��@�M����4�lYcz�)s��k��j�e"�e�
�|��N�s�6b�)>%�A�C)����~�#�˷����묌n�%U�q�2i��S#�JG�7���κ�zK�M������8��<`�����<�S8]�"�Pݷ��ͱ%��ɼ��JǓ���y�Q����>w��l�p�S����&���r��d7�����L�D����K.� ���CҪ�V��R�^��R��M�%Ӷx�����4�y���v֔"�$}�=�u .���G���(�X���TUWx�,TJ��/>E�u��I��Ñ�墘��< �;Y�B���O��6��bmC����o�l���a�JD����Ч$�"O��d,��(�Y���.w�m�8�:s(p���&�o�ީQQ%�=�����b=����mRI}�q�t�n�!P''��M��	����$��ORO�`"��ќDJ|CT�]if�j_��y��I���JJ�(oas�h�\P�ni�@�a	��A�fS�H��H+��" 𴆀�^�B�K�QZ���"�{&j�%X��P ��~D/�*������i~����m��wM�1�Ҵgt�C��gm�H�H���N�ƅ�H���I�;�}Ut�(>?����9N�#en�r�=���\��ȩ=�@�(���$Hֵ�Zt�S릻���.���a/�P���������Z,[��Ʌg)B�.we��5�-���w����=�<G�3�	gt�̂�:�����{0��\ڠ�w���6�U��6����PoZ,!��C�8����+���� @�Kz�G�0�̄Uס���e|����*lQ��-k<��z~��F6��S�7��uh%@�AX�fh���H�}����q_"�MZ�f�x����_�`��в���06��C�\�PS�J���K���SV�	�t1���jI�r�Ƕ�8)W L����3�w}�m:��+S�z�H��眈S{� ��t=� v��Z�HNַ�?�-�I=���W%�#�Q�s଒�!d�����$H��Suu�� !�OD��H}<�j��I��\A��g5���#����LQZ�*U�$7����4
��h��=A��	3����ۊ��O���N�T$��m
bW�goN|�=�7e��훐*+r�/:���\����+�B�p��%����d.���ቤ��"���+��:7r)l%�� ���4�a―�<�㺟��Z6S��v�"�Z�/r�w7�O��F���"ލ̰ޞPU�
�^j��}���>;fP�]����'hy+j�n�;o�6S:1��G��@C�ھ=�g��!�^�OW͟\�Jx@Rbv�@��p�<���W4?�����`=�In������*�^#[fx��!���(����a��FG��t�۶��kX�}*��8���V�lތ����1��@�@�T~�<����;̛4��Jr;>o�A$��D���U�0"1�5h�Ciny
���Up�nY�ͧ�)P�� �ݓ�� r.R���3^�'�%���`��h���be��a�(�/}�%����-�[��}�[��]e�t��q.W����TЊ�Ad3zRSA���
d�j�D9�ոvz�Y�1�5��W�fQq>��!#m�7����?U���J� Ǚ��t���prm1}�u5)�6���<U��,
�E�i�K�K&':�W����<7<۷
��T�,0���1kmk@�Yּ�h���\7�e4[7��RWf3y����ܿdų^�݂�Ox���ң�G�p��ԫRj^��&&�K=Ã3ڨ�W�A��`w ��\5��o� W��1.�o��}�gd�f��_h�
�o���<��Ϛ+�_��	�Do\�	�����,7�lx�X� T��+��q2�!4;���:-|�퉐*i���JM�~���@�}�8Ղ�j�H��NL��|�%���A1G�ny�r�*������B�����kl*V �'�������ۄ�U��hj$̱k~ి]9ւHѮ=T0����0<�u��%fݥ#�����@O
��Z����U��'j�p���4�����$�a#��W������	�l����e��bd�֭��a7F~��jvm�	Z�i8�J��Ξ��c�fH���o�zN<���E��b�4��V�	e�e�m���{BC���t*��@��ɣy��.����7���lM4�h�k�ia(}�C�n���q��|�\XiP�:�v��/�k
J�5�*�ˏI�׮�-�weє���C��-����~#��ʸDlb���I��n��]����������E-�D t�f���A��?H�]���/X���e}���̡& 	}-g�Q�Un�=�֩[�<b�mw|��J���*?ܠ�Ĩ�ݜQ��kwެ9����M@">�
B=�q�>����GG�v���?�E�X�s�&��Xd=#aaJ�H��K9x�'�NA�v�� �6R�Jrl�>r�~s����.dR�q�L��c3s�t��!�ɬ���������}�X���n����;O�
ny��}$N;��z��O���O��n��>���)�FE-�(�G��F>y�H���M��L�-ߵ|g�	/`�x�[��k�)u��vm������P�/��ug�=�}�^����?g��q���׼0$�(fI?Ew�q��rK��s�r�O�|���\G�D��,�H�A�
��G&��� ��B�ӫ�#��W�w�����f�ޏI�z�����~��7�P�q���ر�)V����Q�ʬL�x�So�M4]�4{��JM������?�� OexP�
�.��cA/�\�J�5�M:!�\�~�"f�_�J A���ZG�_O���{GX���
�[�,%���v;A}<�⵭g��Si�ߢ-2�B�_N�`sd�a˘�ր�1��N���Ք(�a�&�P�"�t:O�GZ�	�	n0	�� �i|����A�b��3Q
=�11���o�s)g���Y��J|7�Ko�PQڳ��w|�-ת*�;��8��|kQ�4��*�T�֐@�u����P�i&c���y�u��`�?7��`��/�D�Pi���f���#α��9+5�r�B��c��T��k�K2��V'$qDֵQ(F��:l�QV�����.dt�eɏ�"��#b/+�u�t����p�]/%��}��o^���vr�%ðH {�6ڔ��L@:��wP6��c2ee�r�^�HU��:鮰�%�%��y륱�t��&�t�w����´����5Ü~ꘫՀ��u`�f���3��
��UES�<�z<�S�/�L�*HVmz����ш�Ջ������0�)��m�^�?��N)P�z��¾y��te�1f�(��yF�F�(J��g��F��|��������EI/m/k��\�u�#q���v���73��yx�u�T��{HCwZfCCLb�����0D�g۳z�xb�0�����G�������j��/O�'Q|,n��|�]�Z���0A+���w6҅����D0�o���\A���f�g��I��۬���1��v���(��R��8	�y�T3���X�,X�
�؅&�5r~Θ���|  �@��>��\��R�9]���\�Z��G��) Q��hl��8�F���X ��q�;d���t!����g�h2�}OV�,�RU��S|_�nL0���^�GY�JY20@�^_��{S�S�
nj��0�b�e2���\�aE��w90â��o㢌
`�ޯ�Φ�[�P��\m�:�=�M���[��+��*>C,w�T���
��$Oo�4���x�'��7j�f���Ew�EθiU��Z_��{��;(��[Mh�N��C;`&(�?w��RP�s��p��?��pr����g!���s�n�q\�?���{����a6h&�/�e����HҜ*N%E��?g<��Xm�Gj׊UH�m��˧����%0�����y�����P����G�G��0cJ�s1]/���R3�:�z�*��n@�������zd��0�%���N���![Ř��_9��%U��P��TS�Z1d���D�7	gs�|%$S��������fc�s��]ـz����
gt ���v�؛*�c��>'��4ǚ�zLTq����dV	���$NN�� ֿj�r�Գ��71�#֬-",|3Q�Z��'s�B6aE�^VT���Qn�~C�৥W�gZ_6�� ʒ�m4?$�֘�&l�W����_��ʜ>(���Y�I>e����)��?�+���|DW���Y�K��R���;�gtI�����=�q��N�X�Ips���(�e�Oc�(���"�o㑀�|R�j�^N/�İp�:x�-�Z�N��9��h鲖i��TN��"vH]�o�^���a1�
hQ�n�X]�{����%*l:�T�nK���W�I��A�V�6ӿ��w�W�Od�	)�%t0c-�:m<���"J���3!��IR��Q'�����<�Is`���V)�G�>��B�s�x��*W�C��˃���U�ҝ����E�A?�g�Y�,
0g.��~�a�{m"����'��قدK&c$�{n�����Hs���7r�lΐ&/�^ �N�U�z�E��t��1�iD���7`�x�{��Ь"�����ąsl�9��|�����\�47��K]��