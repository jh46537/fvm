��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��eڴ��XD/=���~U=����.eKUl )�xE�>uE�}�:�"�J=t-���=:Xw2��u!v_�Ģj��wr_N*�HGa��� H�Ak����_�R�}[e�n�W-i|H�)vśǍ��'C�~aq(�{��3�۔?Ut�vs��AsHzI>t$�'XWs	>�2�R�t��e=4�N�P w�C#��Z��A�0:ϻ��{D����X�b��FAiF�k�"饀�����o�Y�e���|"���y�ϑ]��X�V>o�b�'��Q��'Z��xa����_�X�E-{�R&	s�����E�)�`��
�4������L�f�A>6_6�8i'���|�D�$q5���E�8ӷ4	B@�&.e�]ѱh�I�C�.g��x�Ew,��Zno�
 ٹ`�[�!����8�.��3�C������L�-I_D f�t�#36{iv��Ķ��W���A�Y�����D#ƿ�S���]��S�13����H���u&����bbJ⠛R�)�WQe�¡�wy�{���0M(�@�dl�C�^��o�ٺ;��
�,���15�e+>鎴����Y+fi���6�R��B�{��_p�XT�n�΃T�%�d���u�"�J�3����O�
^%�.�_���v^
�.)��_[��G �H����1�,���1mBb�0�d��i�1�U���
����Gє���
s�M�j"�Y��N)0�]�*�]]�P�+>0��2�]I
`�����G?�����;��{�@ס�/d���t�=P�����e�NJ����4o��M⽏�)�� � �sHTr2��Ju^ˆ��G.� f���6��A�Â{�mٜU��k�C��8��/�Q����5b�B��Q�0Cᢌ~���ӍQ̧�Ԁ���o&r��*�bU�X��~�`��o�ֽ���܃2���m���[Qi��tgט�{���.�u� ��Y��|�W�Fd����
ؤ��N��u�W��r�{�O؃QWH1X���c@S��aRðw�ri�E�������|�����Gl������a4,��^wc#��X9�Dt'#?U="�G��z ����o��qG�B�	CP�gB���Aj&�5~��h!���r��է�Z�Z�LM����9�6�=���mV�S��]v���b�_t��F� �I^���H�M��/E����Y���:�EuvW4�5�qh�sx��+U��v�Nhw��~&�'+ڜrk��%2Q���x/N�RY�\.B��|=��p�v�Z��}�H����r�[g��vb�Ō#;T֍�����嘯Z��gFON��R��P�_��|��bN*8�Iv:<ܼ������<Jڲtp�X�����X7���aZ|q���#@�
׹Ӑ�A���Pbk���>Pf����yo+,gc��o;Nm	T��G���q/�]� ä�B*�E�xSul�/�J�GNb�p}4�C0E�q����,׍+x�\/;XR;����hڿa�>7�P-E�$�E|o<*��.��4����*1ZI�-��*�nq��rАh��n>f��q����G�l��t!�K%�[AÀPa��mFc�b��)��~�+�fL���g�mݩ�+��8�d@�r��:����x���v�%�P���{�,�9���U"S��٧�0���>��M�cC��oؾ�nI�)��	�7K����b7�K�O��b��wRI��GQ21�o��H�k��n��j��y�upD��0_��V��#�B���ayߢ����j��n5O�/O�����&�h�<ؖ���W����ȞC!�]C�g>��0�Cm�V:�*��Q�ѲѮz���)�㗭�x$�@K�*	/�w�o��_�4�sӇ�7uJWF뜇��:�;z�b3��Z�K���zq�(�N� ������~������<J���/XMF��~������2z`*y"$�6�ȱ�x��p���<.E%#L�g���3�GS/�IF�q)v
žC�~�*(T
=o���I���	��8���T����"���Pc}�+!�I a� L(3x��'ZP�Y]>�>Kb^��Ц�1���H-
<�v�G���ʔ�V���;�k}�k�:ҫ �"y�Y������G��>�m)w��V��A �^�}�v�|f�$�V���q`�4��S��FO,��#]?]����gk2OՎB]'����I�D`��}��7�O'%�͆ND���_�]���?��"���L��K1xPpl�m���< Q���$v:z�D�^�$��I�sU�^���(Kf	2���OYn�Q����͖�އ���yfo4*X��ś\��o�"�&LZ���A�(l'X�u{[��5Ű���c�F|�N�yBV\!����߿���Z#6�Ո	�����m�2�ݻ���3����و�J�/����*�$��Q�'2�Y�E�s�'��0�S�3����?����4��C�\��P���h�(�c�v\� �S�w���`c��}�ҷ�{S3(7����3~���x�'N��nҡ��ZH�ٮ��*� ���dG�Z6�F⅖�eD4ě\�+e�p6[���@L�_����ЍQ� ���ݑ*|��E����ɲ%b������Ͳh�����v�<��湄�k�Uʰ�z���5��b�7j�we��Q�n��KT��ˏ?��뇥��}]�95S���*Z7�"�֍Ho6���k��Z0��$E�g��M����r�Rn���i��Y���+vL��dkD�����H��$��ŸeY���~W�$(�K�ɍ�<P���~Vے#���g�^h�2��x�JW/�_����H���M~��ߨP�0��pC�첤ʞL�*�7XpxV{��s�ӹ:���U�x���rB�vGIO�p�iNQ�J#�T��2E�� ���Q+�l�C�n9�	jzy�8�_>ӌ��h��<��n��"߲�v��@�vS�Y1�s�}��l�oK�y�<Z$�W~,���L�9�1cng��~9�/����	~�m�:I��sf�F��}�������j�C�Z�^2�$TXYVn���<��}8�Z�`��.���\bJ����Di�`���N�i?+�xJ�Hv��&��֔�ga`5��n��#��n�7��[��xt��|���cH���
W�q;9���;DȔ��S��w��� ��߱�2�G%�[[���@��)}f"����;�Z(��\�F�"����q+�nF�~'�b��5��i�:�l��a"����^d!Bʪ׶q_��Y[V�i�S�}��t(��CH��N鴰��9�؝�H4Y����Z���w��n��Ѝ~����yr�à�Җ%���1��#Fvw������
�D�Mo=f,��3���O�p�G��5{]*��ųےI�3�����#ԙ��ɗ �Lae8I�Lj��>��������ˎ�;~^�� ����Nio����zJZc����[�j)O��qg��1��8�"waN\�LE�Q|�H�W<�_�Y}5��/���y1$�J��h�l�v�S�2�;���.�g�c{��8�Og��{��~��pcX_�� �ꐕ,�Z�n[7�����Z�a�/���ri;�4�R�	쁋��2�08r	�8��k�Tʝ4�B���v�0��E�)�D��RG�����Se����I���6{ ����"��8��C�<CM2�f&�a�j�fѡ�8fM�W�j|FAWe^����1���o�r�'>P�Æ�M'��>�M[�Y��@x���4U����0����V�L�_�Yh�ĳ"Y���kP�G�(%���E�Ya�*u|!CO��s��%
�φi�G�w}�q�x�B%�N۳Y�]�B�8a��^����1�+�ƫG���Oc�V�d�?�$5&��1���Q"mƫ���>Hs�t�ޜ���%����ےge��A*{И9�CF]AԜ�0PHw��t�ͪ�X�<�h[�07���O?�����M���,�������ei�%u㯢��owh�#qK9Z~��FM��f���ԡ��]30'�e8H��6c�F}�d�5�k�G�s�:8P�����i;��+�7�sj^�~��l��Nyk��/w^T�&g2�>���A�;���Q&W9'\YI]�ݩ�Rp䲫Scꀻ�P�
�5,oU�hT��z��bډ��]�pE�ْd��h ���I���򔠋,��v�Bv~+�jg����~�,J�_��^k���П���%�RTu~�����=@�,