��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VHՉ�bs!���v���%�G;ҊK�|sjF�M\���]���<��	/�[�����>���J�>j�f�R��Q�m�Y��-���&5����c��>mfM�~���Ŵ��M
��ݎ�Q�J��9q`n뤬Oտ)U�Dv��T�Fr~<�����������f\��a��R��_5M������t��T�I�t�|��Z��@�j�0"Zب �¹m���m
F-[��h
{B��D�3l��+������9�י��LP�ܷ��Ep�]P�.�7�?�9B���A���)�W=8s���|ꍎ��	�~_Y�q�~��A5#i\�;����/M��IT�������,}��#j�mJ���PJ_�%��Q_"E�B�jI��ϐ^���,�d8��!荦���a+�Z�B�gIW�6&e]_�5�����'� ;r��	-�����N8`��a��
�$1z� B��xNs�+P\��R��G��	F�aD0}�g��OP sTQ/g�`b��?`�I�ۘ��Ur�<I��v�aN�"�F�p �$��Z�a��D���"!�f%j�,��'3a���ߡ^g\{cڠ9f��:�r�n<��P���>�8,�x�AZД�k�į��O����zK:!>���:�)�彨Ð}_L��ky[ny��X����p	ka�~v�v�b�g�/Ǳ[+���������j�_�y��<2js��=a�7/��I�xA�$�L�kEє�dɋA�Nb7ȹiLt����3Wo�{w!_!j�������U_p[g$��X��C��s��ɩ�(�������[(�a?�c�+q5��/F\��m_�Se�H���F8�cC�T]q�ڂ)W�P�C���k�������9Z՟��>Mn��`6�E�E{�cp����Q�t��	�A�t���f�B9x���Ȼ�<V
�����&1cEˢ@�� 4�gm�sJ����#lY�Q���W"�{ԍo����5~�� �h)p�*�VT������*:��W��"S�9Gʘ^}�䗗�k.vw��I��e�X�@��l�� ��O\������dl�0Xt2u�����:Y��h�e��X��בֿ�ͱ՞+��6��Ѱ�r���<~n��z]b+&6����s�����:e�*�{����q��)'5�}�����PWÑ:��?yF�����wl��V�p@����ϱQic�+Q2�L��Z� �R�xu5�e�6��l>^U)N#s���?]�!<k��%|��f9�\(l��	 )���DD�M��T�[C)D
��&gRѠ
�����@��	w�2�︌��va��Iմ���� �䳝���A�2K'�nM���d4�mC��􋾲#Q��>x8�n*+#.
q�&�{�LC��8�}b	x 71�}9�6t��� ��N�������O�������uH����V�uVh@��/��L\�#眇p6��wͬG���t
�6���Њ�:\�N~jpD@���F���m>�x\��c�UH�<J.�����):yyG�b�B=91��1Qඌ���K9��+��D��S��0\��TSʣB�:��\]����F7z�~�O5h�&�"���rL`#���ZI�!�)�����ax#�->;=��ꪒ�҉�P��Rݤ<Bm���!A�U�Sv]{�h��}��0"�2R�a�X����� {$�K�MQ�M��d��h�?�)ƼZK�����wH�"�.��of���.�It�W`�Uɧ��K�mC` �O�MY���G���\�z�V�[KhIA�y}2��3��nx�_�%;9���nK���
+ ���_x\�"�8������&�H�8[g"��.ڊ�e��=	*LC� }/����ZW�̀�%v���i��ɓ�p藄��^`��ҦpI���ij����(��u��%ĵiF����&�0�4>`9��ǭ��t��6-�=>'9 p�S��j��	͛�T.�/�Ӭ�$fvT|Fz31q����HhԼ)9q��ʕ����x����{�g#FD����'g�n-za����F�^O-(���4M�m�9�o�{"=�%шO*�нU�~&2E��p|�$@���~F���XJ��l�e�A���kɅd �'�$��%F�}2y����@�A��]/J�ڨ:ۙ49�X�I,F,�}Γ-���$���!0��f�F�b�����*Cn���Jԕ�ta�&o���Q�W�=g�`���x��B��U��B�Z��0�9樠�>1�uҒ��z�A�[`9��1v�m~A|�Ą̤�MbE�TE��>8b��S�ei����˘���;����}��K��r5Ed"�dh��/LCdW
�]6�s3M� �C�E���i�X�»�Tȸ�+X��\=���vă�žqU$�o�g�ashܾ��kt�;�����!^�Wm,�a|\�����k��ӹ�Ce�zc�=�$�&����ŏn�@3��B���?�;�g�\D
*���#66�1�<L61[��"٩�Q�
��C�<5�(j��<���U?=#&W�PIk�03r�Zje^c�� `euV�$���Z�`V^9uMA�1I��}Oy�]>t_����e���b?m��*d�� �T���]床ᒒ���z(�X[RY���>r��B.ʹ$�̬���S��Gy/ZR�#*�D��,phcM��g����4�Mwو��j/at%|&j���͂�'ߥ%y�8D�D��cc\�K���Xj��.k'���Cdf<��n���_�rY���e�4���MgR��w[��;�6�M�?`"��f�[=v�V|��4��7�Oۖ�A�?N��
[� e��-G�s����uE��h�2��ڷ�]��UN咇���tN��r7;� �ɏ��-��"[0�,�P��O�����.��
@@�jn�kkmc�&�"s�䯰�h���'ɣ���tS�d��`ts���`E��s<��sI0�kG��?%���F*v�#��qC{ b�"Q�"_�z�l�e�趢l�ǐ��t��� �4dX��o���=�q����{W�W�4B	���jʪ�P��`�j=�npY�̎���1F�*4�A�
�Tas�����kE�$N����{�x����c�t�#~�瓧�l��m �w��U����9TZ������Z���E��\&��G��kq[k�H.��
�����&8t<�O��N���t;�g�]�<��,rm��D	����1���k�Bk�1�Tc�q�4p��(|��#$���\�����[���f�h��UI����l7�Ä[9}v�"�Ѝ���=ݎIN%���힕֣�.�g�UT&�x�.�}$�����񍻅��ʿ]�!�Q( ��_�_��ǣ�^Gw�c9<?,���Ѓ�� ��WD��ϡ�nl#Q�ɖ$�:�`%��Sg��_�E@xq8�z���7r o�Ia�H�,�[k�h����CN	��nkk.�v(��G15��U�i�}Z�M<��}�A*"�����gd^�����Gx��Ą.�w��R�X73$
���⸜��v������f��PNyǃS�����:l+��m9jz핯U2���2���BaT��oRڪ�كd��1\��������=���+���S�C�1�������'n>�Ln���I�}���;a�f�hk��X������"p�G9U�����+���?�7y�)}Y��5�7,�w�L���5K1{d9�ח�� \�q����U��5w.^'	
�k9�^��zB�<�a��������<��G�X���z��oT�t�ݍ��)���(������vIF2��Ǽ���h��P�'�*�Øӏ�Z{�х���lgY]��%:"�;H��D����N������Qъ*��]
y#���Ⱉ�)̞�kx���3PMj���^z��V_������`�:�?y	�A>�K��Ց��}�QrL8�r�NT]po"wp,G����8��팘E`c�d�˫I�)�|�׺� �!���x0���* ��KxŻc��-���!�]��;���Y/r������z�@�YD����U��|0֖�|���s
ؔ��*8
nK�G�(������%YA�$z�.��{|?���j{���wYe��,�͝��9;��PĶ&���͋���w@V�d��,�~W[6�X�����\��*�'�_|���R�0�D�UX>���43=��3�Fj�Vi�s�L g�������;y�(��3� NV����	�(7�Ǧ2va4s%��x�|������·X:�R �ތ�ެ�T4Qs*^�$��]�
8}l?:�F�P@=��¡��Ą�We46��~y��ܭ���WT�$	J����Ʒ�Cr�<�Q�n���s0�S�DvŴ�����f?�§��ò�[cg~���Js �7���X��s�ar	f�Rp�	My�NA�0�9��b����i����1R�å���3����1b���nbl�9<t����1&��j�쮥�S�ѓ:����˘{T�`��v�3�9�!���#h/
�1.E���?�W��bp�R0cy���R��K0���e����u��w��
����?��t����Y�ԃvP����H�zi�K��L�19���t9��|�-������X�{��y[#2��%�W��ri���-��tJ�qv'�@��A%�59�t��[������5�P	oon�L�_�$��#�fr�T���1��@M�]�N6�š6�|���2 �>)H����8[_/1j1��v���/f�1$pV�p�\�&����spD��8����V��s��|�P�o�H���&��T�[bΕ+D3˟Wl@��-4v��zŽ�t�ǲ�@fN
Й޺-p+f��۟�� ^	�sޚ�q1����eG���!Z^<�G��b輓��3��������b/'�dA j��SY�n8B���!]����.��%@�uJ���)�r�,�o���\�W��"0��o�^�k4�z�1�m_��ȯg�z�Ƹ�/$���emb��r���
��f��4��w�1�Mu��[���<�w 
���J@��/m@�����cd{-�?(o��s?Ap�;��*�IɈ�+��x|Z]�pQ�� ���~��u���m��tP�ul��y��_r%���\ ��p.C5�hy�i <{��Ot�������X��];Y�7V}�1����X���
�?l�(,�(/��:��l��`����_���e�v�upy��t��0"�����k����v>���2�.+ܙ����z򵔀i�����'�A�Mdɫ/ON܆�G^��O�/QQT�W]=0�ŗ���?T��]�1��Yp8����n�tΰ�n��ln����NY�Ahɜ�Rc��	����}�vپ�?��r��-v�%�����8+�k����X�=���ޝ�H��Y�N%��Tv�,o!̺\;{ ��& �_�?_�wXOw����F���F��#K{�u��ж����f��關��j���>��\w�sD5E�b��[Q�j�Ka����/:�������ҼmS���Q�+Fg��i#I�x����i,��vL��B(��I�H����B���Ο�G��v�=m\��g?�a�·l2���Ս6���V��� �|Օ)&q`1BZ=�Bh�>����0�����)xR��ӫ�M��/3�~�P���I�9���<2�����U�Ҍ��d��
��,��0�dG���7eV���+�`��� *c0H�3��6�����M�b7J���p$�~�ЪñKDbs�#y��v]f��~1��w-��6�%����c�'o��W��z�i@`��F�����a+p��(Z�D��r�jm��u��V�F�{-ж,X�N��	��c�Hpe��#��Dz���U{'�q���Ӣ�:ʅ�5ᜠu��,�|RߝMT ��&wF�?u�gZ��R�>�i]���
���T<B�a�{��v �����x�&\0��� Cssp���|��n��Nه�7>L���DF�VuTI��sbbBI+ۀ���08�~��4bjOz	N��}t{����L�Ca �H�Nۙ�Z�@> ��~3�e� �Y[�g�~��z�c�X����ʯ�:�BS���m��zy�ڄd:Z3.^Љ&>�$7Yǉof�R2����K��@G~�߻�N �	5�X��m�11-3߱��� ĳ���qB���Ŭ�{si��~
كjZˉ�X׉��� ��ť׌��e
w�d�ܥGi�`.z��X)���6z4�e��Q~����T"�I��(;�h�o��G��x�-V4K�J����P�K��j�+9����E�O�H���A�#�+����Z��Q�RPvfP�F��	Y�r$�ȗ�?�;�șs����}�}rf�?��O�
r>�~�����^[��õb��񌑬��w�Dս��x)��$�]7��?�ڹ(��G�=\�NS����H��X���#�u�(&�R�7u2Ԡ�Ѹ��d�K��N]t?�9^-m����sn�g=����8�W���.����S�]�&M��@�&�g�d��/��6����i�`��~k��x�|��:���M2��Q�b����{~\pQ���u�]AEq���t2����Xi��E�0����|�]�?�xb�l gN�B����ʣE�۵C]�9�K%nJ� ����`+F9�o�Mvrx��߻�,�Ý`ݙ�!Wdp�?�ϝpdHAՑmfu��#���o�z�茩����V4�\��,Vshp���rW��O��3r�b`���:�8�*u��rw��T�)�����0�ƚ��d*�7c|ɋYA��:(y�4A*�B���j��/�����(�ú�0������)�]��IQ>E����c�t�k
?���M�f�o�*6�n?ص2��w�M�'b׋#`9�!0� ��d��������7-g���_�`�.e��&��}��}R��Z��hL�j}_`ʿ@N��:�{��y�Zn�^_���v�����>WB�)�zx�܂�BLJ�3��&O���w�0���c����e�����(��h[�o�7Ԥ��xxgm����
Y��O��~^�;r3Ļ�Vx+.S>���Q�'$;X�A5@�2},w��4�#1a��}��6Q�k��E�:�h_��@�]�d^���R1��Nt�مJegm�M#��ML�G�҂fXXxX?�>�������U5�'G�_,+cL