��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9��͇��<��R�v7��ASEoV�6�l��%S�,V� pD�hh�Z�A�2J�}���,m�-�Ki��F�U�Q���>�H.Ydr�/�Q^û�-H�<26z���uU]3m�p�wQ��m���g�3����Y�X�^*���Y��?M�x[�fN`�A�� $!��Q-���y�k[��A �	�=�S$�E��@���MC��'"=��e��������~��d�,є�#�^�dާ��LF��?s��?��F���9�Z�q��db��f�\�0ӵ����
H�V�S���gL���I�g�e+E��y�����]���Vr�͝�[Fް+�����:Qwa�yI��ckW4�3f2{�<�o1�?�mN/6�s�G�#�#�c�@��T1B������s��6�O6D�{u�x�F_�jֶ���@�4Q=���u�4�;�
D`�x'�
C�ȱ�9H�"��2�5��-U�s.�j�1-�u�m�<O�PR��5ȉ�H�P�n�d�v����A#��7�T�_z����Ů#��b��M�O�NS!�&Jia䅾|���*jΐ u�*;X��&Y;
�w,dӗZ�2�L�^EX�L��a�j�� >�o��Bv�:�:K���?ԍe�\(����2-����^B�D^�nN��	�\���J��� �_X`�!�gr�z�֧��Q����{4}Ha�������E
��*$@z�����O0%�ŵWTK*��8$^*�f��Ζn��<�����-��'o>�;���������aeV�6�~�����rdzK0B�LAs8xb��$��>�V08�ТP��F;����)xM8�p�)������tꟑ�C��.8q߻�q�����q��m۴�p��V�������?%��N��캭N3�)�%M2�^�����;:��8ze0�����>9CU�H_�Xh�cesg�X���H�z��[؈.\�����U�&�rҔ;��ƎE4�/����韀T�jn�p���Ǧ-��x�{�
��7t0�YSx����5��v�{��l@��♙���7��]b��~D��h��ӻ�۵�⢬K�ү_rQ@VLA�+�u�_h9 ����M��B1�s����H-ˤd�F�+2@S��c�y��㝷�¦VN���(ӦP����]뱵�#�[^�X`UZn/c�o����y�+�.Ņ� ������>���`|O;\�Ns�� �fN����d�?��џU��: ���Q���9�±�:�<���9|1D��L��L��`�����O	1��i�Dܧ� b�Ǧx-X������*��qv���ߖ�#U�8x����73{�;�����]2<C����q����݅�˙��l����>a0��8*�N	JO8��w�N�W�ŉ�65f��Պe2��P�A3������W_���V�J�|io���3��Qn��Y9Z�V=OF�n��d���	��t kO��S�F���I����aq�|��,�[zͥ�?cl{@$uL�c�9��_���ǥ���C$���B2­�wo�1�~a�`$�f��ՁSK+gMc
w<Ic)��O��X�b;��K��8�< ���BU�t��ʕj(��HJ#����|~�����8^$�TOm�*�g�j� ƅ�x|�O/ĭLA��4�̅��n�ƮJ��0�{G��s�]�%Y>Q�^muJ\�۟lC��K3��#�v��ύ�|�Q�ےl~/h�O��~���n-�
Iq��r��IF�y(~�:��zߧA��\�t=��1˴u�W��U���Pt����N�-����ĳ>�2�=_���݇`��p��͡�2d�Εe��|Ⓞr��L�	rg�5����f	�Q��g���鯟�j�$�W,l~@f�]|�z���`��@�Q�0D��w�~�X{M�C ��z�R-4x���93�g��7$YS �Ľ��>���~U"r螺�k}�@W��L�ȾPўh��>TݱJ5䢸vܶ��Έ��?��~-�I�%51�E�ߠu%�;��4A�
۪Ƙ����,�byj�i:=g�$�7'�?H�b��@	�.�7n�ڳ
`�д??qg
Z�:��ǀ�摋�b�]�.���rk�~�˪�S�ll�II&\��.����nCx��zX�Rֻ����{�hkd,���~*v���1�e�6���t�=�[H�h~�m\�m^�q��#G���3Ϗ�w���s�U���)��CTS[Y^WC��0�Ł �|�[��\�> �m������i�U}�puZ�E�WZ�����4V��^��\ ?o�OҋvhG���.�C"�v��`��m6�A�a��A~��ʻو<?v�Uݴ�Vp�B�	,�} �S9�>Gn�B����OU7&w4�2�I�����2�BYp�3V�A
8��4�c����y�4�c{X�Iݎ&O��u�����#����s��2�&��X�K��R��A���_N�L�6ʏ�DIU����� �5&�#���fb =(�Wp�%?6q��& ��Ed��h�6V`��Ɓ� �>	�#=��FF��j�+�E�%Ή_^��62 _�j�K�e)g�B-	�g8{>��|��Q�2hu��A8�Աa���,t�L ٕ$�V �wҌA��`=v�u��I��l{�E�
s��®�˫�o��\���D[^�,�K)�厌q���(A��T��\�Ƈ��-l0�;���C��?��-m	
���n�B��	��7��dzpyEl�J���A
�>���Z,B���g��.�,C�!3���z{�VqH~��g������9OW�ʘ��3U������ڤ����8�8�TZ*`�/���15�K؄	���Ԭv�i<�M }�[@�-{�Μ�}^�^VBgn���	�]��U�c��S�nz`RӺ�����r��#�Fw�E�j����
iL�\h�(o)��9ՈI׭�թ��%�SL�;��Jn��y�q�NE�Qw"��a!�������}+���y��*�ԘH�ёZ�n���hw�6�ZA$��XOm�N��5�O�)"4�4�t�'R%�^��@A:��H���m>;���Ԥ]f�����C�x��(�L�] qb*�(��)�����0���#���(�i���n�6il0�p3�%�����=���Q���>���S�Iun1Y���enN7�7k�6�b�G�3R�'j��F��{���՜�25i7�.P�T�F0��ဟ����F��3-�M�dO)�R����cp&�z������_�_)����*6��$A�-`��S�e����( ֲ�%�~�����q��VF��R�k1��}Z��D���]\��.���a��8�h�s=��(�2(2P'aBD;�uJ������������&\# ���)o=Vmo�C5�[�@G���-f�(�w�!f�e�
������,�{���2�mw�&j�V���b!����`��dt¥�lz�Nt���ĉG�&�d�3��S�����t.֒�[<mj�Ed//��d��PP�SW�1өn�r�+tU�
��k�F۾�u���y�����_�	��0d9
��M����2��7��oB���b�hx@���[M�m�jiP ��R���%Rm�u�"�du�wJ���֔�Tx��'xZ�6�%���	�CY �<,S�B�����;�~^��=B�R� 4S�2/E�g��F�F����}�V
vm���i6���Ahk��A.Cd3a!�G߇��_��?B�c���yI���w<�aAο�haJ�hE�2Ѷ��p�`� 7N{)8��Ԏ�_�����~�W�"�ƆD�u�QcB
g�|Y��Es�E���NR�葴C��Q�ۃ�x�H�4��p�:�&Ut��W�5��:�1b@ckbOKL6�ܭ��D�� 4�o۞d;9�e��� ��������{Iȸ=Ƥ�+��56��j_�����0eWuZi���.N�[�����"���>VS���N?���d��o�d��
8��k���a;����7C?f�S@��L����.�
v�^�۞�Z�G�_�	��JC�7|x�7ݐo�,.z\�r��LYi�/|�����2T۹��o� '�$�`Hg	V6��'܀�E���z��ۣ2�9~G	���|hsT�MU����V�~6�p���_�wӚ�o ��s�6J�,�[�õ�m��O�t�z����=J�W@�i��՝1[�v�S�At�#�#���ye�s�Yaװ�ܚF"�2�`��O"�dj[�b�l�F~�)�0��j�PʉL��.0�r8}�Mj)�+{���s
KG|��i)��W�l�(�|��1�ǿ��@�.(�>�����.�I�=����3u�[\���ID��4/�.�_o����q=�'3D)+��Y���fȖA�9�����'^��2hV���xNyl:l�'����?0q�Z�k���`4~U�%���M����`8��WًE�po���ԥw '
gjf��c���(�[.|����Tl�8��W�V�oP�@���*��ؘ��zG��b�L��ٍ�cy����_j(?9�&^/50�Yu�l\�nR�Ck{[�7��}a��c���D��O�^-t�ױ�Jwt������Ԙa��f��q�)�S����/<_V������h�N����G_y� �y(��lzt;���h��wGb�O���^��_��T�W�����ޚK�4v�'a�#�]I�As]����0�����tvm��q0K:
�����!�=���:[%�ȝ,o6� 9~㡋�؂�2��HY�d�
��O���gI�H7��; 7oFI�x�ԛy�O\MN�܅W��,o�	>��42�߲7g���n�� ���{�K�tM�Z��y%'H+3��X|;h��%��������o��΁�Pm/@���,5��}`�U��37HK���@gG�.(u��|����Kr���7p�smc���9`]����1E�ZgS%�+a�TI8��ᐰ��j'��-���d�hӂ�
:E�7��Q�Ep��67�ZFŪm_b�n||�\g{.R�ñ��t$xm�bk�K6�6&����O�1��3�VWܩ%�
�&�LB���H5+X-s�I^y�*��
���fyz�X�l��B�����