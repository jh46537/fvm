��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��&��e�uDb���JG�����*�<�oBr����a�%��X�H�\�d�ʷqDb�Da{���M�a����+��zVrX�{��Tg�bG��[�<&i���|���F�sb���w)�Q �#�,��Z7e�����c�؄	���A���Os���?�
�0�'�ݗ���B�M,��ڭ𝽏q�3�P,*��{Dz���M������6��M��aM[AtsT�(0�9�\9��(E�ڊ�0\+��n�<���?Q��H4��= �pv�n�qo���Q�㕡.��6�*�u/Uצ�pt9(��(��L�{��.<x����q�]I0o�]Fd���ƉS?U���QǗY� l.@��!4�.���
�H�gr�Vm�,O�(w����6�c��� ^�êH�\8^:��94�\���rf�̯qR'����|������$�{�������Z"r��V�|��H�[3n�K0��4�9���T�d�k]ZH�Lr���ҽ���:t2L̹��Ǳ�%j���"���Bu��%N�՟!���%c[����l��)N���#l�yA/Uy61��:Ka�|=���IB} +��-M�#�ܬ�+*/ ��[q)(��zݟ{օ�t�ܾ꺉�Y��Ћ���?��_���n�Gb���up�l��D"R�3_�-p�p$5�>����yQ_"�[��p�%�"_Cw�S*���X��%��0�Rx��HP�c82�)�: Y�õ�FIK�vBv�C��ÿ�N�f��ӎ�}�� �i�b8���*2���H���6.GXjkQn�&gv�@wY}����{W� up�)��|bl�{`�o��+�0��w����qH+�-I�,�����#K����}\���sÿ�J����i9U����`���
�A��hج�Y=�,������k���Aɞ�0A�+L_�!z�5�*��S��t�����y�!���!;���_$���M+�BJ:1��g(JHmz�<�R������6<�c���dDf�&�[J���t�}ĉ�<&�����ĸl�>J�fk�*���@���=p+ʊ �����2gIj���Yq�P��;tJ�g��Np�PhB]0ߣ�ɏE�Ocz�'$_�[�
�p�=H�S\*3�l�\&a	�T� &��lZG�|Ws�*��r���9[���K�0���իG����Ip.���.TI�"ؠ<���)�fé�w��n����*	��9C0���ӳ�(c�|�X|��*t&��!��&1�^*�1%\E.|��?h�+��N�S1��K�Tޅ\8n�k1�+wsSV�;� �_�9�8N�yTH��	�)�B_N�X�Q�0
�3:�g�k�F*L2��Eǡ������s���n�)�����Ѵ���Ծ<HL>F��Cǟ�yQ܉+iUP���V'=��F�ᭋ��Ԧiu�9�i�g�R�*��7(+�^�h�����{=,2� �0֘xC�@��ñB����xI�
܋�ʨ�p%�V3S�Z�Ĥ&�J�H�g�mA�0A��w���䙘N��굛�����),�?�o.$�:��&�*~h�Q-�;�!��DNƭ�qH�	 �fҁ>�`)��`�}��>��G)��/J�f�MK�K�r�ug�F����P���j@@�L]3���#I��7����W�h���<%;u���?z߿�3-�Lc����.
�Y��=��	�z�ל�����2���v����-��G��i�7�@���bm��N��|��K��4�FB�Ԝ�Q��o�Cwt}�8wG0"c�A�[�/���n]!ԐO��s �U��E��G0~��z%:n?oHRE񖀎*ʨb�a�pJ��9ߧ�7�/kl�[*��g9T�n����;��j�R�؝��$J�@���be��7xr��m��N+��S�&Res�����T�N�<�韗�ˋ��sC�G6�
V�Es���%�_����Aq{PL@�8p�9�ݴ�[r�,B�&��sae Uf�7%�^O3
�����;���$9�`�9%�r�@�j5W{�Kܺ����UE��`�~i�wݪ/Y����H��ŧ��R=�!�wR�F<�T���50U���[۲l�8�+��e���lhbڍ���M8
��9�$h�nV�9'!���DN^.� ��3���3o��c�}��~�5�{�<�a����9�����\^H�h�(ƨΎ���yX�qA��g��Q��v9n#�z���lܸZ#�lr���hEl�l���thHl��s�Q����+$��R�z��"ȏ��C^�{���{�����~>�t��"$ltn�@���Ob�����F���[�ς�Ͷ9F��^��nQ,�r݀o���	q^۟��*�~���h��:Y�S�\A���Ik�*��ڥ�!��w���q�T���z�,JMk�ٜ��Uҳ�\%��dsţgO^t[d�_^���G�~X''���E����(�,	g����-pב����&���߳��2��u��r��?����`�@�.��^z���{�7���E��c�R�Mwjd��(�� 8h:<�� *�7R�ťI�c�@�����@�bZB��w�G*�KH���`�~A�H����0֨�1�_l�+ ����~�_u���`�t���6\�n�,*�����o����G߭!�-�"~��{���:?j�����v*��0��2	���Wy�s���W�w��]�V�oa@΅�@l��[{��=��Bnq�lxce@F?�~Gk�F����]J�<�!;֍�EE��gC�B��S'����o4R��L~@W���,걨<+��l����i�¶>�x%rZ� ���-���f|̳�/�h��n�q��?͛U��;�.G�⤓���Qq�W��� ���%�!�J��L'����si�k�ؿ��^cOk��W�`�%7Z�E��%�H�J�@ك�B<)-�vS0&0su��$����KO�u5�_�]$��"L�`��X@�H\�.�\�,�Ƃ�e5e-�Cu�z���[�_���*[���o_��?|*�W���Hʏ[�>��{d���g�������ǌWc����u���HG��o�v�7�����ɞfSݥ�1<$Om���׋�4j'��V�Xۈ�3���´��e�OT�
���?�Aw�r�z>ۼʟ�D7(,{ :Q�k�˽ڢ��fZu9Eh�Y��Ng��ӳڊ��Ƽ0N��U1̆�Dt?�Ə�B��u0�h'�C�K��v�w��{��ۤ,߮�����@(E�-��c�=vYXh�ʀLV���2a��65�Q?�����{z�<ImB�li##���^���0���6�"�)�bT�7��mǺLҊ�{1C2����#�1��F�B!!9�5 �z�4!DK�T~�#J��7i=Ix�4n5��=�-������s¦�P�KԎ/Fֹ��5�휷�Z���N���(�_L����p�Y�D����w$7s�Ԉ�}13���$
<������o4��#8�ڣ:���~գ��iV�,1��ܼ�p���40NT)�%�_��?�Ŗq�u����1�a�V����YK���㠝p����>T(��6�檶D�IP���+��
��S��3v8�t�f�\"��}�#��AUs1��I F��@c�X�` �O+�0>.��'a����F��K7_���VK���6�ֶ�Ґx�H�q�u��1 �Lr3�^�>�zG����c��@բ�.p������~gb��%�!Lj�F8a~7�ކJ�8��A����ʁ$�T	��&q����ص�u٣�N&Ÿ��Z�e"� W�f6�K��}�4?_#��>;���+�`�w}1�H�M�P\NI����KF|�C<o�t�u��c:��+.�W~V��/�М��c�e|�-G>�k_���?���c�.;Ƹ��������:V$�	��|��l�idp�=�9����vE=y��kיТ�?�`������3�����3�l���>�NSc�SOY���(l;(fش�V�xV4�ʻU��UV���"[X8S1�J�fE�5f�আ�����_�i�x���������9JZ!��M�nɋ���* !�j��o��}�9HԬo���ݧ������N׉���Gyh$ �"�d��1��ae�C��^{k�>t\�]��3ܶ���h�΅%����c٭p�8R��|Xk5��ACt��*9�u�K��(&u�����ɉV'y��E���&�U�=w�*�t< I���{��ầ Ju�����(�Y�Zg�Qc���O�����0<�K, ��}������R��NI���ɬ<��Y@�����Pf�\��f &&z���mB�ۡ��W`�|���_���Q�o�8��ٙ>l��DGې/P��\��r 7����Wv�(����,=�&z�n~;S*�n�ܲ���b�n���RP�~�ߊ�r�ݔ,#�Ju�<϶*=)��9�=:����H��$'�R�Gn��Oܼ_��a�ԧ4��\O���a�"/G$��V�\I���4k��>{r����ak��V">9�W�8�&]:��^|����D�+���[�vm��yS��`�hx�2��d2\e0�5������Q���%���>��>B��yAO�;�H�?G���$��{+:e>���*����	"�
�����1�(}�WT��-ȫ�H��s���6lL�^(���#�����(�[|�lQO�� �z"a�ZA���ڵZ��w�$���K��X��R=�.��[�$v
�������m��
��Z�Im�22����YYSO�h���/����(�Vz�<2GG�/LB��y�1˴:�E�q)�9ꁥ�_�)���r��lG ���{�.�g��ѿJ� ���Qk-����������z�K��������U���������0,4�^�7��e�Mu��X�	�FSuuo+�L�����[��O1) �3�K�L��%����(����Jk0��o,�'ݓ[cl�7C&`o	W�����9�߅�2|!O���R&�kگ�: j���0���.��!����C�b��M��/>�l��6\m_L��#	�6h��z�ǆ-��Fm���O���b�R�R���bV�Q��u�E��A�a���zd�0y�X��hPk&h �L�XS%?��>���J@(�x�r�h��W��Vs�Jd@[�i��9�����k�<�
�o[�B���,���3V
�ʄ���C⯖�6Ct�	����)��M�b�# ���>�"�,�ݡP�?��#ͩB	��(��*���}O���J�:X�݀��`�סNNt梄��{�ќ$���ȁ��K�Q9� Kr��1�m��i��opڅ�B���q����l�>�Z�k�:�_���F�m'%�_��9[��S�cZ�ųJ��C>��HΞ9��[�-cS}:ܮ-�R�SF��a�1l����i��zu�G�u*�kx�lhu�M��Jx�� V�p&�j=��l��b0އs����~l��y���k�W��Vո�`G]d���ډׯ��5������u�3��K�^���Kk���G�5̖]w�$MR��n�?��u����zP�͙�a�g�^Y�n7	��0����1)*�SNR?s/��$�ǲ-+�Cjb��w��Q��*�:�<ge]�x�eU23u����Xn��ķi0�/�S�q��MÃ.��d�uy�|gE���{z>�� �[@N�vTOu�24>���l���$��LG�f
�7������KJx����^��Q� ��Z�{A!j�C��As}Mbk{�mqcA�'�J��l��y6]��5[��)�wU���FD$v���7�45*���B�c�|
�XD��Ҁ)�s��<�Yjڀ��d�Zr��H� �X42zP���!�
 �L^���@I_#�?ۺ]�_��K�����$���tb_�x��G�E�ۗ�w-��H1�M�˅rY�1u�B����"Qӈ��%$�Hӌ�+(DcG�/�D&!�Jѝ>ef�K?�_���B;�kz��^��v-!C��$@g7#+�^�����5}3�$9�A	��"��vc�t��$�y8��Bu�R:���,�M[�����ց~s��N��W"�o������<+h u�&	{5	�[�*�c��^6�t��'��Ԏ����$$Lb^b&�.�����+��P2E���k�UxKF7��l��Yݶ\J�(q)E�"�D��B%��rF޸�no�i�����ɦE� @��++��@7�i�y=c��u��E��@��������<����\�܁��熦'/��
FyC�4Bϥ��E<��o~�R��tJ��琕�Y�L/')Y�p�OA<;/����6��+�g��ͨ|�Kn����r��o �c�kD HU����S�z�u�8f"l8����Ta�{����3,B.��Iٵ%�(S4���<�Vg�t���v��3�/���Z=������Ud&F�m��n��[��z��%���e5n��k{_f�d��rQ�9;K�����Y��=����R�zo�����X	K��x�,��`���u�5)��Pi���8�@�p���=X��r��q,����Su1���m?�ܝ劅�����Y|߭�6��q����&�����c��7'��!���`�K�YL��n.qq�Ш�o�Hs��D�J�O� 2|����U%D �����m_g��&�� ���'SflQ<��n�,^k�
�����&����I�b�7�<�|� �-���'�D��>����Sڰ��{�m[_KQ�����˹����Ï^����n�}� ��>��k-c*�=s�	#U��K�����}�;zx�k������ce��gQ�J0��0%ٖ��_�s��%ӚH����k~�~nvf�z6�4�Ԥ�4%+o��tU�*��(�1��m.�%!͞Jӛq�����&��̛d��J�%��r��y��!-L�$��Z�+�O#fS�sY ?��am�[3]
;4�뜋�$;�89_�8�*{�@_����!���nE&�H������6��z���٨�ȭOJ�ʍ��E�� �w�a��REz����@��g����Q!���<͘�[�hA�H�P<���L:"K���#D�_�(��q���yK�|�|o����9hio��u�3 �xب���k�T�_�)~˪�H9hNϴ�Q�O��0��e�����F6���VE���oǂL�s��]y�G}��be�^�@��2�Aow�V<LBb�qw�D�Bt�(�x��֩�Ʋ�P@bp���K�#�1^8W��R��]���Ǝ[��ṓ���EB�g��K��Z��r�K�H�#Zo���<]�L�FV�o6�i�YS0��tJ��Sc��J ���|Ub��`S��҃�9Ւ���Mb�q��9ļ�Fy�f��ގ�U��h	���BK��T�:GΙG�,��`�o�V�m��=����O��l�Fa�qBw��x�Q\��l�(QD�Hu�*��z�]KUa} EƠ=��I�uV�w����Jj��:,Q6�q�K��`��c������q>�,k�{5���lC��\$R�R��o�*��x9g����Ѻh#r�/��J��O9�C]M/�eg��P,7�t\je��MʣXi�&��o{U�O=рgfY�=�Ok�^-T���|�%��.�� h��`��n�8p\8�]���w�`��G;����=��(�8��A��$�'јr*+f;}!����"���s�H
x��0"�H��_ �%!��>�fF�$uh��J�e��J�g\ ��\J��?9�N��Pb?Z���=�
�nK�>�Z|�?5/���`� d���)�y���Y�}�>�:��$��s�pحr�%��s'�u��%����3խ�U��v��T��pq��6�%bwpRQvSHG��<��"�Dk�:Doo�뉗Q˳<�J�f��"�g����[=#>M=,�I�z '����c��U��!jVL�����ȑ"�)*�ĺ��*�_(��!�cο�$�*�S�ҽb�$���{��=t��[���?���.��>��OO��/�c�dJ�p�vѫ
v!��Ė[��x��]H�`:HZt�ɮ�}B����b��D�tv�W�=��d��!I9�z�vȸS�@�zR��wW*3��-PB<Za�W�ڋl�	
��ǂ��T�KO��h���a����& 6r@sg��N]"[g�a�����'D>�-��'�-� !�|����X��D�R�
�,���#kA�=a#`U�6�O���S׬ٮ{��t��Wt'D�6��~����U9��j�L��9{���x�wźV�ؙ�T��ݛ�vέ}�Xȁ����ӹ5+|��B��י<f�,�'ay����0���B5�!B1'/UV��ņ��߁ɏ���v:��1�����/�s�yQ\\u���Г�(�l_r�>�6���`�hp����c�P��9�q��v(=
a7.�,�?�@d-e�K��b���&��`hj�2�5����s"ל��	�<hnJ��P�I#�ro�l�:�4���+�3]��8K��5m�X(��6��8�����lW�9��|װIXpjĭ<NK����/ۼ�!���R�[�[���.�o�~�����P��%��5}ط~���T�EY�X1��T��ȿ��i\ �K��næd����/�ۗ`!=QⳒT�7���Y�)F����/w`�x�L�~w1O]&v�&�R�.Mb�%��t��T���'W�qj�����-�����l�R�a��]�>�����s��@23	�1
f+?dذJZ�8Q<�79�s�X.�����3�=L���8�k[+����1��K�`��!�M[R����� B�⣙CxzDr~w?�A�t/~����2��p�4[s� �w��B�I����m���鞈f����y�Q�T��ݾ��Y��MtŔ���W9���l@s��_,�k7�����^���^��P�@:�fS�1���7+d�^˕��y���|�2>_��Ҏ���nY.Dړ-oJ|ʗE������}y��?���:�N�r����j��������+k��ܘ6	H�-x�{�.'�o�5�2�'��Ud��E���-kY�/��
��t�vK�N�2d [��]��{ި�V�x@��%o��i��83T��<�����s�8vt xY��-�q�,j�Ac͂��u���dc��x�)��A���F\��cKn�%],'U"��Z:9#�����m)�Ý��R���[��:���(I���bq��� �}Y�3��;b��Չ�t;�ܞ5� 1���|���[_c|C}+�����JB₼��A���`4oem��kE��\m��E)n�/��Li�1�Ţ�R�ݘ~ŋ"�T�����芲�0����2
��+~9���^ �A��LU0��|�,w�1�͉�J]>�X|D�2��e���_�	�nS'Č ��j��m=%�$𘦒C�	����d{�FV�K��Ô�q��4asН'��Q��Ӻ�u�z�<��!;t�[2k�{��6����n{����e�j����8N�e��U�ur�L��3��q�^�s6�����m�����
���DF5,���|��Le��C~�R�V+@E3�W~vM,-��6*0rC��"q��gL����6>:�إ��'/0�qVOZ*�T�7D�t��@X�O��~�#��"���He}�`�Q�P�s�����$a��%�t m���}7RPT�_�V
p�P�� m	�'M�#�O���l��o���	C �*i3en���O]e�$ɖ���O�zy��x�M���O����o��c��b�t>g@�v>��'o����X�g�n-�VA#w�K�
��D���7�"�H+>�a��$������ui��+ �X�n?N0��#7=*F����4&TG"���';^)���ha��X.` o����x���d#H�ԏ�-y�z���|�>\������"Z����^_`c�,74AȒ�����u#ƪ���]���<}�lLi�	/M>�)Z&�5=���cv�^),�_;U��?-�k����밬'�S̷{�h� �=9����c�)1$�0�9d7�pY�qBL���}������{f�N�0>2|�e�KO���i:b���b�O) ߺ/� ��]^�u��@Y[Y"�K8�R �P��B+}h��`н*�#d��)$)e\%��/�:���=���k����aY�){�xޭkkٶT�~7\?�?���A�%���2㏨ :&HS����D��t1��s��G�f[%�hAv�&��c$v��n�GUOJޖw
·Ng�+`EYQ�T�P�������o��V197`L?<��lF�Y�s�C��ͫ�1��E_ JNC����%3��2m��B"��vL���!q�1���� a�g��[u��L�r��[8
�/���8��K��pme	�;`�C��Y�����T�}��~LSU�0=^gI�Z���3-dN5���{�:9d�4�2��>��Njb��tB�G��7��W���WsZ�3�Mg��2�C�I����Td���랉��n)�v��ADe��� ՠ	�X #����;�H״m|���k~
���G���L���J<�Ԩ�E�;��{un�78��XN?�˾A�]q�i$�|��8�0���3��
�"1����@|��#Dtj^
�Zޯ�Grt=�êm&�Da���!�j��Ii��F�_D��
$�5Qݮ$��!�E��pef�0�}k˰>^L��~������,x�Ww��5�~;n+��1�4l��;R/� I{�'���0#b9��p����~h�̝�dR� ���z��n�%�Z��E���t&�����$ѹ�b���8�]����VLBN���K�z��A����@
IDF�q��9�4i5JL+���c9�:��0���7�=w���o�cg�<��a�&΍n�� ����$֦�/�${��,�?O_�'S�x�������Y���|~�D�����oM���j�E��,�m�)>~ᾉ~U	���N8z����Bl��e>ac('�@���+���ba�eG�o�k=��ҧA]N��XTy9��	υL��B�WO`�T�<L�X&+��id���_��Q�3-��aF�z:�D�����Z��&� ���$����S�2A�����1ڽ5��P���kW+fql� R���߃ "!�!�\]^�1脬��F%�tzR��?"��{�w�]�s7YK㑸�ƙ����� *@���UC`XSyF�B j;n+{b����bl,r����S?���U#-����#�ZwR8��Vg����U��14k<���^>4B|fSlWj�묬(�f`!cYA�grK��?I޿ vZ���l�6+ ��RoTo����
1C)>���K����	+Qn�ͻ:1�'6�4F
{(�@CF=�=��t�����M�&��ȕyGjq!!J�ÑX���[�$�ΩH���+C$S��?E�y@�D�c\��N�����D�x�����)˲s.��&��X�����s�r]!��f�|<��)  ��C|����\�~��fV�:wQi��݃p8�}+/v��D�6	o����v��V�u�a>nƌl'��XМo��j���ʘ�	?@4�F,M�BH��i_�N���k�T��8`�VKpu�`��Uԓq��;���i��V�R���V�^<�Pe�M�vA�vX�xQ��r=}8�H|ֶ\p~�*P|��gk���7���^�s4�P	��k�,��(3�[+X����<�8��?6�d3�(��3��/�E3z������uҥC9��o��^L.,�Z,B;����#=Q�X��`�CZdR��3��)�0��<��^{+b�>?ٽ������W��;t���zx�(<W���-Jޝ*۸��If7���n
ɔp�D�<jkKi�XªT�X��g^��3x`�L���EC̒�bR��C��v4���_p��n��2r�n���ҹZ�߽�9�<0�(g�+=�G��\>H=	�4y"1��$*�A09����
�޹ބ�����^z�K1/�*�Y���#�WBupK2]�-.�D	�t�!~�I�R�Y̯�Pv�@�86T�>J�P�r�=�����P�!� -R�GWd܆rVf �	>S�ab�DU�`(��d��z��H$9&ߗ�!\�TS�3���9�y:c}��A�[:��XL�u����?_�N�&|��I���z���9�$|�J�����J)�AC�«��I �y)qZ�1,�-�y�j#���Wd��O�D�LM?���w�2�~+�\ox��?hGr����C|�܃�<F��,���w��f\i_�����(�k@$�?�.�˃��`�pH���MU`�Q�ni_�#�Mz�������ӯ���;��`$���P����,�Ga�5_S���,|_D5,������"xB��*x�1q��ٔW*�@�1u��������@�)�v�Xvg�b���L�Ğ��d��Wf��o�j:< ��|��8��K�զ>��}���w=(DHz�}�@-\�)L͘8��-5�X����%�"|��þ��d+#~���,qm���ީ!����&����K6���#ǐ�P\{pǁ)��������90�Ld�6����;.��Az"�#�2h���R����D��`O)dD,�kix!iu.��|�� �h���+�w�g�V�r��74�`e�/U˫��q(��-RM��A,~�ˎ���d`N��R��䬗�� C<y��/2���B��&iDnn7���-�q�����^��E��kc:/Ŕt=d��BO���r��cTQf�y�".�&�� ��7��L���/8�M��L ��W��|��?�4�e9~6��Ȥv�ݕ�Y����K�#z��X' ;�P�W'q ��e�4�]Q�{W��W{"vi�Ð� ���V�`0ԃ��C�/��m��g�3tc�N�3
�o&{�_��i� WDәvߏ=j��Ch�y�D��砱����fVt��t^B�m�a�R��UsC7xK�r��77�� ��Mٝ��7�')b��'**R(�������M�81�M?�M������|n�a��>D���&�0&vp����!p����/���e�Y�mV��I��˜c���������7�d���9��/��s�_�j�T]}?S�z)��*T�ʃO��x3!�Drih�o<�U�7���Jtö�|i��f�q�i�ڭ��Mm��H?�<�/�j���$�4��N;k�bb+��U�z2�6/��
-SYƘ�z�Iz�ӳ+J�xrnp�{d<�+a��T�\��G��oSk����W��x����+����C�XL��m7���v[��b������ڪ�u�V�u��\�nt6ѫ;�cA�s��P��y{äIe�2=�N-�c�H�H�&�^N"q����ت]@��u� ��C���v˸��	�:�`[����K�8_j:��kX�a�{�5��[ 0��F��;�U	�yE�0���K�'����c�.��܄��@�	�ڱl�cB9Y���6D�&z�簽)�D�S�e߮.1@�7T|[��}u3���:q:��,������Y�2֡a����B�%?_1�Uu���>�j�S�g��!ƹb|�GF�w�pz(�н�I��]��+��$�*�x���(/q��S�튐Kɞ�t��nP��������y�3����V���p��H����%_�������}��V�@;b6*΢d�&������.(�ӡ��^A���k��8|��T7�����_�|�S�����4]\Tn�Hfm��e7!��#Tq�K�xzY(&�S�����-����9#��}n���mLAڷ��K�	+���k6�����`J�d�N��Cωp`]�`1l����'h���AX�����ڪh��l#Wz��	�����9i^�tX�ƣO�oI>nU�Pʐ}1���SFs`?*O��A�wqukD�<niE+�ά&i�	�s�Ł�@��S�wz�$
r"1%pͥ1�����$�B'Q��r	�5QG+�(����*��v%�(�VF�h���WѦ��Tl$���2���f���N��Pnc�W�/��O4I�q�����Of�(���/l��W.��������r�p�Gr�z��zu�.n��y�_�TW�9宬�5��ql+$�94f��������ކj�%�.Fd���CB=x_op�����g���A�GE(�m�p8~���n��#ݼ��&&�m�S���,w�I�W̾'��绰m�L��(����9���	�I���?ސ�T�(�%~5��x�7����?A�&6z���){M?.ؐ@aɍ��U�P�
CZ���N�Uk�&�*�ӡȕ���T	S�����q1y���4�'�9��P�4��u&�%K��i�]U��+�}�Pz���N��߰B�\a���0nu�).��bM��� և�h"��D�6T�'��dx�w!����[KS_����(�ȴ�v�C��W����jZMP�MV�%�_�Ӳ��<�c�	u��{�����������k�c<�	��]�������O*��~T�=�m�Lvg�n�"�xo���Hcv�����g��d��m�SԈ�5.��"�8Y�]att��E��{�mq��%L2�`.'}��[R'덨����i�' �
��4jF����@�Y��S��$b�n��h��>�Go�'�ͰB�w0�Ż8EY	kc�[|6�+-���#�<>���e~~7�"��9X3�b�iݱ���y��	��L2��e��|�ܤʦ��`P����Kk|NA`�wL���S���a��5G��۫���t�����!gv��jF�+vC�_@o��/�UR�"��b�Y'Yb2a��e)�-�=(g'xi���9�L�3σ��=L���@������S Y���1I0�D�{�&ݕ7���aw�T�:�PH�Z�+�v�����x�^�O�S�h��w�t8'���>��N�m,�yq��A| �!t�'T�m�8��Y�>8��Zl7t_8B��^�e'�{#�9t��;f��q��KŸإ�����-��C����D��bz�������a����{ۈ���0��#��ej���w���I������m�r2T2����l<�m�:a)��R�)M��۵���N&4a����\��I[4	�~��omn��u�I�Wkٷ��l�C={jlg����5��pG[��J�O��G8�����aN&/c��s��5}B�l01�CX>P[Vza��4lk(�G�ɡ~`�pD���}	��"�e� ����Ö��T.�^�dMb��%�ޅ���~�^g8a���0����Wxܛ�A���qŬ��?�)}
� i�3�|kda�.��ҹ�)QD��ȝ^\�X�k
m�_��`�k�Fb4z���zF���5q)�R�AY��fPe����&*�j9D�w|��2���>(ɇ	I&B�K`����P|��U�C*�f#E�A=3��V͕4���3bѬ5���*M�ٞX��l��L8d���sz�l�L���rَ���gr
i�g�o�j��x��V�k���7�]	,��8x)�645P����t�`\=���h^�N� &��{&Q�����]���E�Fr�zv��H/^*ө�D �@�v�V��E���@/�o�;!�͛���K%S��S�N�'0"�����b0]#��<Y�/�ס� �j��(c�},٠���C�P]!�qR�����B젼<��/ҬϵL���3���2�Ww@�B�P��U��2���b���c�6ׅ×dQE��^�D.�_&H���7�w%68d�j��Ln�	�V��L$ ��#�'�/����}�R��P�y��-'� 2����>m��@��B.�}e�2F�I�1�0��T�Te
[n��Wx�^�6�DE��!:su8����r��rê�-�8�P��+J�F�;3�P;��.}n���od~w�iS_�Q�b���{�}f��^O�n.�#v�ž�h�e��.E���o����3�a�c�F8�E+��5�98R�6��u��XX�H¥kś|���שsf����!�	de�~i�ี�7=��t��1Ι����/�w��(|�t�,�|��gZp%�&
�k^�?���i]>�.�p�P���[�����֫³��}5��4��Ѵ.�	�L�%s�2-��2/���KӒ&shJ��5��5���sz�!���j���{#	/E�����k��S;��`���<C��2MN3���9qy|�-1q]�:�� A�>���1l�����9�6�#�}*��%��.4kc�1J�@���f����>��5��jMz�L?otE�9�t�d%�YߞZc(���o��5]��`���}�ġ�7��$��g�`P��.����^W"5��{�:�P�}Q�U��fg3�+����2
��.D�7_i���B�#6�����]��J,�xMs�x!D?�u3l֫y�z�S�@'�㜿��z��U��ː�4�ȣ�-|��~`�LA%��#f��L,Ჽ� >�¯rN��ͬWM�OJf���$�}Z/�솜�n�P�������EY���>�M>��ܿ�K9��ׯf�ZG�/	IA�^Z��"TO^	1����ʦ��T��8;�k׾���^ɜ���޹��|0\���d����aC'�y�zl�Bͱ������iڸ�{�/�ҸQ4bx�H�)�8��6��8V��/�@��-�*�ZJ�O1$0F;'u�G�D�pU�����HS�!S�3؝|97��=N�ԗ�Z�S�%`
��w��Â���X��T~��5-�������m��@���_i�ƛ�Z�q��~���nD�%����4I�Χb��?1�V���r��j��1�6�{NgYwW��If��vV+��v�Ӄ���V�e����Kۦ��~mn��z������"ё��ܝ�E8���)5s	ͦ�.ӭ���+���2�0� �#��d�ȿ����\��T��l�u<
�,�7-�N|�{S��z�b|�����(�a��?�nXߤo�������Uz�Jr`嫳������m^����Z�iI>����T��P0e��D�{� s�Q�jx�[N�u��,�h ΀�|m��g�DAU{᷊������{�}���ӊ����Q��[�!�D5:t��6�Gl0=\C[�����B#��`�:Ŷ1|��au���Y�_�Y6K$�S�A~�6�K�<!�&���=(��x{���7z� �&՛zd+���S��E���`�Pqv��~b�X�~��9J�8��8"^�giIпח������?��J[F��d+�lx�R�Ed`��F��9n�vvl=էߒUT�^��P~�
�`12�����wn#N �f��FtA �j��K� ��uLp��]����9�Y�������?�0�᝘c�!�<=����{5��U���ZF︷l⭑z�I������u�`]w��Ǩ\%{� ��;;�N�ob8���C��?j['7�ʬ1��tb�qD�:Q��pY���y:X���9��J�H�e�?_��FF�`��仇�o�	��|4��TT]!��=�����|�c��*�d*��$���4:q8���b+kD�|��{�P��U��`�2I_�0�]OQ�0x��mV��X���(	0S��C\��R:���GtC
���T'r9�E52���V����ּ}t׹��|�[4�=p{)\�d�TγH����4��_@���!Y�9�3b����Hw4��H�xI=A%�Vi�SM$u����ۻ�J���T�f�v��e��W�<��'I��;�<"�):�AN&�D����ӥ-8���]3����n$k�-f���g	�XG\�C���ZV'��Rp�ml\'�r��-��0[�<B�Q��yks��G�nb=p2!KJ���~��+s�I�whu�k���K�� }.�N"U�:-�+I<��i�܆���cv*��������u�ےVz�b6��o���i������,�̣���P�q�0�T���{�u�ֵ��yOz�����1���w?��:�;1D,��[8�ӂ[��;����D-y�@��/`�[�bctN�f���|�+Dyߠ��YpÛ���U�V����h}��}���U�������#P��D��6ł2��-}�m�	"~�j!WI��Y��y�.5]Qþ.
�\jpg�H�
�v�<Y���mcV���K��/2�������A!{�7�λp�V�`���J��.���}�������,1�N�c�����n�
|��+�)-��L�س����5Uw$2�$�d ��df��5��m���^������[}�}nEIL`��q1�'+"h["eD��n?�-P�{]�	I�o�4j�Ғ��Y�V��UD��S	���֑�H%Ӛ��h�G믬5�T�e$4C��6k��׎n8XȒv�=�RY:C�Lc�j�o�Z�]ʹ�?���j-�uP���$��n뺇zW���-�i���݋��^F�Q��aN�x�M//K"l����?��*w,�!���
�˳_�3�9BDK�	�iNbn�m;Z�>���;�[�_�k����r� 
�q�����������}�Y�N�N�������{�6�l':���#��ćv_QL�R������bd��Q�%0,����׎���)�F��cb0U���i��_�[x~,�+�;��$o0���*Rͪ��Rsݾϗ9*��F�З�[��j�2���f떀Z�u��_f����xynv@�%ӄ�j�By��i��r$�c�Ș��ZzJ�eԸ 2�Sз�`z*���׋m�#=o�)���N��|�[PL+���Q�����i8���l���ne=k������p'5>�E�m��Q�	5����\$�;��x�
�ځ�Akx4ԣF��|J{�����������w���P�-r-z:�*C�o���-���#Jf�]��e�b.��?a�1(�N�q��l,����T�@��#�]�R�N������|!�+�'������϶"h�X���պ�p�JSQcj���L�@��ᙠ�����3ղ�*��+0��1	�Ϛz���k��W�����헧��j�n5��Z�)0!N �R ㉃X�l�χ�R	�%c��{�\����X�6�&��̪*�՜{B���G�_�3?Z7y�����F�)�mŗ��m��\7CWH�o�ݢ?8W�o��L��[����waǮ��G�N���	�#�}i6'�+ ��O_n~���ȼ|�Ħ������7��bq�t���V�n�*Z�L
����a�������
�B^
�&6�!6��]43��խN���|��Y��Y��ِ3J��0���Y�%�]/h�h�|���:s�u����1��tx���cidĸ�aF����W�z`�O�ՠ�e��Bc��\�(4�rH��~6+��.H���5�˅�*�T`K�m�n}��g�唼�q��t�n>'Y,�Lp�p��}`�CB���\��s���ժn��O���+�D ��#]��+`�_N�n_+���7#�<.&;$C��
���8Ž�,�Ų�$�Y��A��Aw��Ȝ��+��Ԅ�hE3�+�B�3N_�塲���ħ����p��{�6'�"��S�����T&i�1����˰�w�Ē�Be��c�N[�o;�/[�����h]�*�q���'d`�>��R!2`=��}�:���ӟ�O�c_l��i��9�?��4�\�)�{\���5e��"d��$���$�k���f�Y�\Y��zh�-�mZr䰺���{9�1N�'H�q���q%U�u���۔�v.���N��I��c���Γ�ˈ/A��M�G�b���gM��c5�8�����"��J����Cr �"�_�Z=m�pn;�E�X�lp��m�ȈCvᣋ>4O���ha#��]�˄~�(hϋ�yaZxR@������Y�IIb�B�@��D �}�U���)��m�ʟj��߃��Wx4b���+��y�I<�����2nL�XI��b��F�٥k�0�J)W6�Cl�場]�hL>!G���͘<��
�(v{�UA�n�B�&���d �*�%�� �.���4�OS)��|pI���|=_k=��������vQ�HK=5=�b��^t{��j)��ț���U��)֮,�*�!���h] �j�җ�~o�$�;N\�=��Ϥ"���֔Móa�ƿdָ��'��nŝ]��a41���s������/�:����A��p��q���H����wE��)�y��Wy����Fz�j�<����Dj;���ڽ�-��X��b�%EN@��D=�%a���=K.�v�-�`�[�`7��[�I�4�k������Rg���~q��i��M�[yuF��ICmY3��W%�SMW�z�$���D����\ ��mb�42�vD�3�ۻ�Mvq���o���ʉ�-����\<�c�<��k�w����S��9��Z)M�<��3�f�I�{�n]�K��A�Ѳ��p�rZ��z���i�
�?�g,�ۡ�}���̬�lZ{E)��5��(�h�-��\�8ǐؔ���3��w�	F`1���K��y�)iU	�>2��\.�&H�Um̖�\D|r�*2_Bfg>�-&�T"��k��]wf�A��u��"!��?�Lj&�f�D��=��۞�g�ũޅ�i�QL4{�c��NG���>�%#�r�m��u�8/h�I&Kͨ��"#!��u|1qYS5�祒�NrG�.��Ԉ�
�\���)�n�~��S3iɤ�K���v�<!/��F6�r�W�����
}�+o��&����Bc6 �0
�m>�0�FB���넘o{��K���w�W��Dׯ��~F��{K��=�]���:.[Q5gƬ��+��-۶�lk��g	g�\�+N�]v'�)}���V�[�Ȁ��~8>7�cC�ì[�4D;�Hy�o���%�E�fG��?�&�
����$���Ux�nD��̂���~�6^[S���0L��;��yS����.����/&�^���t��r�:�|U���H�TQU�e
L,U�L�9�-�(��-��d4m/N��8=އ����"8&A���)���}�(޴�j�,��2A",I����NŖ��ew����4��*�,���9���%}��W�9�{c7�O�����wGw���/�a5�q4�-�?�(��C�����깘�/�;:�.U_=�W��;�A��>�B	!G��ܯ�\�J�cn̩�S�Q��dv%��J��`19��+�N<��#�˚�DG:u�}e�z�)fy�=M��a�ķt��<HЉΎ��дE�)�r��PhWK�}T��Uj?��p@/6m5{��E�h��9m`\�]s~��=[��׼�ӊ�>,���L�X�[=?�&������"Z[���f�nÔ"�L�%�s�q���R${L��QΎ�֎J
�n�xzO;�D���b+'q�d���^���K��a�!��^C���?3�m�9��z�����֣�k{��r��W+�iG:Β��hm�ּ�� �,*��ߩ6F�i����m#3��a�Z"����mkZ=��3�x�uժ��|`��'�w�օ$,PJq�y����Z��L�<�Y�!ު�2F�=����I{j(�Gʽ���ݬяi>�TR�~ӊ���U5��C��dT�I������i���6�w�ڒ��$�s��|G�g��1.B�����2�鯎���ZI��|�����x�w	���7�!5؏c%��(޿���v�D�C����#��yq����t�r6�@�9$���g{/I��
�W�
���U���q��Ƣuݼ"���v@l��O(��e|��N�2~4`�~eW��2�s[����7�[z3"�߈ܲ: %��G��M�������^��k�kf�o�ýA�J�<�ļN�sY��Ӝ���1�`|'�-�lBSU0j�>�21xq)
G0��nQY�j���w�� ��j�J���+�f��Sa{��)#�i�@yy���n)RUX��	���¡L�n��{6.�u>e�r�Ȁ��{���β����45  �~�5>v{���o���kۣ��G�_I�m����5�}5߇'�=UNcQ��F5�Ih8xŏL��EGм��Z�+�pxpav{�7:s��
�°R�5�PN���'�����w�J��:�p�G4T銕N&��j�[Ђ$$�*����F	���hM��џ��v��������!��){ ٠K��B�_�Oq���6}�5ϓ"���L��31�*�_�F&�����l��}D%:���1�X�ṿgN{�EL>�}���9T�8�N�[��;�T�V�J��>���jWz���9����J���ʄ,�(�=�7��8�+���wg��B����X���}���k�.�f&pm���`
�qo���a1��i�`���5�(ѭi��e��3�Ҟb��k?|���E��#ؓ؏�	6	
�Q>�1��2 %'��G�a�H[)`�K�����:�2۽ȧJ�1�Њd��q�϶0T1Rp+Ɇ�:�'̘9�����CJi'NiSyM��N�����B�F�tɾ��$ڐ��)�m��`ua+�I�^R5����������gVb�A;�R�= �&ρ�[ʙ�Y�e��cg��'?��s�Z�6�S��IL%y�8��n*3sm�;E��)5C�v$JSY|�Hv)�[!3�!,G"�1V�B�<�{���y����	�F��dzr�$��!��6��y[�<ц펜=�D����9f֑+���
�f�ͳ=x��Ʋ�ₜ�t���Pv3oZ�U����$���[��I�r�gy��������̎���z³�����S-��*��Q�f߇>v�EI������h�(��|jvg9�nn��]�����(}�&e��;�E�����r�l;��ā�cqr������ۿ7q����� m2��4�����)��P'<?�F����4���a����Y��q�J��WK+�W�6ed�M���K~��¤� S&�~� ��Ƹv���c�\�7�;g����7�g��Tym�}���#���~�__A�}��A �#@]�!�s8g������;S����8N7Ⱦ�N��
��{�j1����ߤv1@���}>o��R�p�gy1��4�	T͊���sAk�����qz��5��[ˈ76͜�n�2h��M�D)���A�!$_���y̶�pc�pM���,W����3��S�o9e�����⇢�Be���c�Bj�~ͬf[?����b�CW���c+?Q^����a���Յ�?�3"SA����Nk0xٸ�b+�Bu�1�[�f������t�v��&J�y$'��"Q|P��3�y3�� �f�f(�����w�:º%�:�Wҹ�U>|�H���N�{=�t�� iy{����`�Xr����E�օx����r�q�:?f1
��/.���#r0a�A��kߌw4�9��3��+���x:!��]7�4d3��e�*�ɬӏ�V��Gh9JRV���5�fg���Ԝ�0�;p��X������[�݃YC��qɛP?���?���a���@ߨ�u��k�YM0�=��K����b���p簎�����H�n�o�ƅ[#++�IF;�؃�O�[f��I��n�w�+��9C�؈I<G��u#�.��Zx@�Q�42������[F&��4}�����t	�u�鋲_Hk�ḻƕ.�Ŏ���������?B�J�W3A��?;��a@��B�#?�L�Lo�Y0�r��7�3��p�"�<�[+z��&j[��N�Q�ȇE~�� �O�ԝ��е�z`��B+mWQ� �PT��z<��Ƚ�i�����8�rB5M����r���_
�
2�����WIQ��w���)̼W�������Ȍ���^���#@��n��.@��)��Hi��z`�z苴�)ih0��@�-=�\Nl��2xqGfƖ�K�՞UL?`no�*��"M(�P��FL%wہ��)B ��{���.���חa���W=�kzxi��!�D���8Q5 O�~V^�X.}�gK������Ţ�mӔ���Y��s��C=m�� 1?��S�0�㷡PON���R|�N��B(�7��j_ڣ�����(�v��xVTC1F�v	E1�'һP� ]��:3����$�Մ��� +��{������1Ժ�����W��؛��z�%H$��c|d��cM����|V <��6�댻!U�;,��9o{��Ė(�C�� �l-c���C�E�Rv���Y/
�H��_�OA��D�3�	)y �ي��]w��[-���E�[�4�ZZn�pcKެ臁�F|N����b̉���� XU,�!�Y�b��a(�?\���I���E�j=�頧q�1;mB�G�
;.���v��{�&���΁y�����Km2���-�Ol7�b^4�k�<2���r!|E�e�7�)�	�� w}��H��.@_��]�g~sw樆�@��z�T"iLp�����c��O�*r":jif���g>�7��5�(��CC�9q�L�xkq�![7��%��-��{�Lm�<X��M����ьf�u��0-�������:3�LP�����|�{u��g}�^�}xO�&1%��~���U)�Q]W��I��I$���%��L�7��4�`��N��s��-ʨ���� �=a���뤯��P����נ̒�P)<�{�orp rf��}�䕴QX1���MO����h�6n�W�9����h�$mX���\�S��]rR˾�J!8���x�J�I��,>
 ^�f�pc��p/ =/"�b���'�/o"d
���r���y�#��Ŏ�>��{��h[fq�;�O��f��&�Ju�<��� ���Ƅ.�7� �mrC�]��GL���24�=��H	�����+�����v�6A-��)%���tm�B��X
�뻦P�L��` ��঴��sӲ�'`��SE��e�k�1�&4�l�����wߋǑ�C6t	���A� N��\䷇�$���y�U�(���=��+5��〫h  \4�,�'�� �:e���IA�E��{�����<"�0,���ml��+�1-�6��L���z�rcCM����QR��Cq��F��������)*��=��V����e���:D#@����'��/#��֥	���X'g��S>��Ԇ��kj1 ,�]�nXܠT̄�I�>�b[�%d���è��p7�T~��\��j@����!I��E�t�}��l�k�ً���%뼤�iŬ!��%XpJ�D£m(���4�r3�%u5���mϻ��M*ݐ����U� ܺȰ�J.��p �3T��U,�R犃�#��+,$g�GN(�3	�O�v�5��{p��iS+T������yخ��sq�M��^�MTe�U��y��t��'	z�&7P( {����6�虬��|L]�#x̷6���L�|��e흏���P]��v�����3���DW� �w�7DJ�\��C�ĵ���q���]����˕ܐ���U� 5�5��ֿc��/	zЃg�}�ҷ~�x9�Í�AϿIǋI+�nL�&�6�
A�V��`  fJ^�[ć��jR#��y�`"s���`�+���w���N���*�Ǣ0.O1\v���&�Vʢ�t��}R�D`& �L��	�� PUG��PZ���uq	D��/z�^�ʉzd�CL�����I���}9�O��.o_�b9��{�f�� ��3����V�*ͻ����B����M;��jgY}�g��A���`��Lv	��Թ�y$q���Rѻ�#�����X��n	�r�fd�k�/�/,
5�{��pDvV��Bu�fc��1��!����j���
4A{O"��i���1X���E��精�g�k��2��胪��[���:K���+� !)�����Ȇ@��
�T�����K4���%�w�uw�/F��ٳ�>N!�t1�4�#,,���72��:���H>7� ?ć���"��sWU%�A�***�4qg��Lȕn����f�R��AUv���A4�X	B�-�ui�B�ܜ�m�o�G�x|��No&fc5{��9��h๐�Z��_y��Jn zyi�+>&�o'J>�ו}��7d�_��x\BI�7ԙ���B�7�ݐ�I����B�g���eOh�~����ڗ�d!�9�R��u���h�\rݻ3ƭ��E$���>�g�I,w$	na\׺Y\�� �>A]����n��\6��P��mk�}���^3��̎��l��?�p��#��{)�G{ |��n��I?	O��OԐ �A���:�萲�H���-�c��3���-��#�_]�BbG���B����L�ƈ�������챌b]%����]�*���צ2�YU
���k?��`f�Ϥ�iW�����4�?;����R�&���f����m[�!���nL���9�mT��s"��5��+�2�瓛n���~�A�^��y=9n��ey/<���F�!� �Q�x*�嘢YS��f��*��)7��T]/4~ό1�Ȕ���҆oe#�5�ǋ�Y�Ȋ5�D�(􍟘�X��}�Բ����z��Z2("��V���.��"�������v��T�翑[�rC&��v1ڻ�h�H��