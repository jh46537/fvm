��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#�~�,o#��uIk�˥W��.��-Y�S~d~rIi�2~�������ǡlS�,BA���z�a"��Pj��j@�l�hv�7گC��H���(�m0���]4A����_s?2tb�߅z��U;���ʯ�d�T�?�\4�?��Ub����J�'LƊ-Ú�gV�]�`�����T�rP���9K�ި
]1@#]����J>�[*�e��	���}�u�H��/(��7�u��{@<ɔ���e6?]���fC�Q
,��ɠAEp;��䵉]���]\6�����Y��,��*u=�fմ��Ű)þ��-3?:�bZ��E�i��uJ�4=%9�<�[��>�X9��<���)_ֳew���q��(����E�GbC������- ���[��\[X��	G�6X�=mG1.�-��/� �~L.у*��~��)yg`t��&���(�=Z�&�d�Ӹ��W�y/i��K��Z_��Dh��u����z�D�S=�"�y	����N>��P��!���t��	��:|+����>�N��D���;q���J��C=�%��<�d9���(X�_�P|6�����}m'6b��GG֞�1�J�p�,��x2�z��®;Ů��I�*y�<"Qŵ�hȵ]�\��}8�M��E���+ÒBw�ۡ�M>��i����o��{k2��]Ԇm�y�ތ� #�N=���H��}�wPe8;�.T��:�WP�&��3iQK?�S~b�i��.�"BZ�Mr�hG�F��8?�%�� :>�({���O^�=��{Y�I2�%q!�=�w:$��;�<�J��OA���t�kL܊��1����v<9��!���rH�%a����N)�Q�6������B6�E����МP�.A $ӶȎ��[n5Ȳy1t�V,
��������k�1��iv78�E��$�c����W�$mb�)��wR��tI�G��o?���#�+C���3�iv:�úY���}�`�L�##�X�jL'��j4��M�!b���w��pw=~'�<5Xܹμ٭�Vkr����1��F+j���V>��nk�W���WJ�{�����qM �~�Zk�Ym? 5��ئ=�Ot���{q4���{�7�d>�޲b{�l���z==���Z����"�����aL-��-P�:�OE
����#�A��!	���}�z��~|�_���s�0��G��#�O]���/�����i�v=���e��~b�-���g;vu:C�"=�����W�Z�əi�گ�?� \��N�*D9F��y�b*�_a�jDI��♔�"2h)��1�6+b讀�Xݹ��m��:��\m�d�%�lK�L�P�:jU@�O9���u���O��mdq�P��'K,��ؙ,$���՗!}Xf���9����������Yɺ���bQ���ʘD�;��;�@Z$�<;�ci��r��uC�Jwq�-'��I�X�)l�<��|l�ǩ��
�P�<�91�:�FhYù��6:��*��m�bTf.�}ub��yϺ2�vD]�Y	v�5DmΙ���J:�&��2;6���N8E4n�-�{8"O���-(k�|���i��!�
��ψ��q��|��qόl��9����҅t==����pL�Tfލ�D��Y1�`�A��Q�Ƚޏ ��q��  $(�]�?��dE��R�<
ZҚh���X�}9��s�vjoQ����y�k��J6�������2�����WOd۷�@*m_�8&I�很!K,%N��[?��]�|�@7p��m��>��\�AZN�H�n�*}�\
3r�'��l�JW��
芠���ǌĜ@�᤽cj��4E���F{LKͻ���b�h��!����}�Y�r��GPD����tQ�[r�s��'|&�����2�H�m� f�t��9��C°�E�>��2����j�:��:��5���+� e;���I�f'U���J|?jZG���!!��x�_�\��"L%�w�Y��7`����b\�Nܴ�;Qq�i�lSM������&$:=�R9����*]ݗ�
ϣ:��B�����.+5Hp��k4�`�g�ѧ6����&�Jc]�ť5���!6�D�J�ζ��JAԀ>��ڬ���CSn|�Y�RmA���'j�o��q������D+{�7
(&W��GLz��;���9�H���8�����*9�Qi�ˣ!W���_�I�~qg?X��;�����[��;�.Vme{�P!	��]��@��زN�