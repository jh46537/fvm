��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�/�CZ�0 �^r��s��<��v���~�"<����IblQ=�Q �qc��=��/d��,2Q��R�~�����tz����g�������$%g�*�B�WC%�)�,]������$�s�qhz-i�9f�i�HݠL�6��᜝>M��O�OT����墛�!d:��+�e��; �}z�L
<��.� q;m�.��ܟPA^Wg�QJ%�\!�w�շ�o#S�h�{(��]�K&b��!��e1j����o�&f_	�UI������26���k�c�뜑�+�I�����lZ���gw�`1��n�{����RA�G7�Eԟ\�O��|�š��ڕ{}G�����j:��$&��cX�<!�+�~��j�C�&m  ����I�c=��	�㒛�j(�2|-ร�BR�z$���>s�	�L���=q6�� >-�^��s��:�����A�g��ᶶ������D%I1|,A���l�|E	�}�ۋ�h����"sh��L���r��~@��|���>�ޥ�R��,`����Bv�61���ݥM�w����ס�tI�����Q��o�`�F�)?=y&�[xw�iU�;>�j*RH	3k�ϗ���
��i�{�Լ_�G������[2�c1�+���TL��Wiԅi�����j]�/<��Qֹ
ի�SM��7I����^������:�D���U͵��Kf0��7��GhL/��	����������&���L�	�^��{5B��t lN����|G��SS�l8����&�s���s�R΀�⛮���a����[�+},���Ŕ6X �O)���ܕ P֜�� �Œ�t��pQ'����Z ��	f�h�z�w_��H�y�T��������DNK�N�� lq=h�B��/^�!m|��jTJ.�|ȠW���M)�т-�%�SDkm�k�����c�7``��\0r�@I����DM�Et�Dc���t5��ZT~?8F~�%<�.��0���у�~��Z�m�j�.����1*�K�$��84��AM\����IM.��-�똣�n�X������ T�`Q��抠^��R�Y�U�D͚����
��v�,8i��FOTo���k�a��'®M�]=�g�&BzέQ���f��v�A��;GN�!q-e~�����Q���{��ϋ*�7�ɉ��"	\|A�LS�uo���u��Wc�=/0��"T����>�>���#����>�Ӿv'*��/��uB\�F�%noӃ��̍�E������E!�	�{���*��8�̈N0+6iOFb��pc�+-bji�����v��ov��H:Hægkdk�]��Ɂ�8E�m]�+Y	�i-3�w�;�U��1A�����8�U{�w����V~�hf}��P�#�db6>t$�*M�-GF��Sd֩��_R`.��W�A��B���R��l�bR"���Mo��c7�p�,pb��h1���b!�{�+yx��-�V�k��9�h	u0��&jn��*yi�\qĔ�ڪ�g�CO?8M�͹<E�CSĿ��Q~"@�Kq�Qsȃ��W��c$�twW�*rPo�P�G��̫n����`�#���,�26��HbE�OE������/g	�V}�Gz⊢�9�����X�Z�R^�����
���˚����R6�ek�Σ.>h#�%��Ş蔀��.R����y��s^�^_$���>��0'�y��Q�
��,���=_:�� &*N��2�ۦ;���3���;s&�M��XȾ�����b�x�ʫ��v���n����C�B���p%��מ	�^�9䈼)�C����C)���c�(���"�3�ĦpaN�Y����+�1�x[MW�q�(�{<T$l�Ҙ�pWb���D�ld���&�*Z�co�?x^ڵ����0��ض��TS�]܌#	{���)����!��G�p� �%FG�<Z8�u<Y���5��N���W�� ���z��u��6o��i�����-���S|졞�Nߞ���2f6�����"�|X���(�.BO"ﷰ�C�(Y��+Ī�q�E����g��L���g2QB�Zħ��p��R����1Q`�|��0�&�!R���Z����pW̋櫮S�?�5`-&�e��U���#���U�x
Fd��x�<�� ����|>��v�y&��l&=��<@R�����M9
-$�M�@��7�U`����V���.Mk��3�t�\> }Y�_)gŊcȪ�����>�$���G�����ƣcA�S%_��(V���F�cc�z�,L�I�m!���:y�ע�V��^0�6|�TE�61D$��qG���s=͌y�S gD�]:->G<�Z?���XE����Id��f��*,Z{�Q��5̀6�}P0��aG��B�s7��c8o����HϝA���L�A�ref��*�:]��8�ɓ�b��L����u�(��R1�$���j����l 멃��n�{���=�5�)����D�@0 zV[ t�#�h�Oi�Z��+5^�fG��d���M���h�����z�2vz=�*^���-ױhp*u��W5#��ҏ ��(�)~E�{���B�l�m'�bY���(�yO��w��ۏR�	5׽�_�:��9ca��b.�����O=7Ҍ�~U�9|��^
J���AL`i\X�&�J�u�Vl7�Ld.���k$#��$��<�pµ4�Q���Ƞ�{�
�0��5S�B�L�	�����;iv@��h�f�)�ʌ�zǺ#