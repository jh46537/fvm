// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tnkDck7ii+PKkCouxROPQCiE9vlaMaDLjDrYNTlMvcw4j+1D8EFyLA1rCVjNQNk3
1qZr0gE4on22PdqWYK7YwwTTWotY2WZLbElYXV7UZPgaxamj+pDseXyD9pmh5vJn
2VIA9FYImOnlSxNkBlaQLiNSii5h9WNcIcA1JBvAHbA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20768)
+WtgVlqyKk6cmXEcI910RvtQ4nLP4ZvqPJ4134momng5YraH/9DrHPr/hRmU1WeO
3waP9BaQzia+WxmSL4cCgemgT6XgbtZ0Pkg7uhnYMH9vXwggyA3cWJiJhGq7D8rF
HuXwii/hcikTeBLi2A2EOaNXASl1RSXlut/UFNnNr+ZYEFanMt+JRjVa3sOQAAsg
MICmZFUWZ9wj83i5l5ZfyyLcp/4HT1AmYmpSHAeZcNA2c4+OR3dscR1MXDEAC77n
oOtTXq2Z/Ubsr7Rxhf4tiSgF8WbpFTxM8Nl3g7FfU9Ylg2Kvovm9qRs5KZazE4xE
F6BZ6EzyBxOazWcJVegsYQifdiFK8SRgjBDK39lryvEtDH5qEDh3eGg7EOvrNAQ1
PdhqlSWYFR+4RrR57avwjxH+VeT+Q67kZVUCTQxfz22N6iysXODkPbf2Yi4yDSt/
x/4gIx0wunNFnDqZ/nxleaStrzBoFivT9kagMa2T/+iS6h8yU10VYkaHa95Y7eN2
JTHPMnRwhUWeFl4FL8ff4/oMeFBNLzKsZsmNxwvtDLSkDYniUF92jeLwYibtPewo
A61KVDBN1ZH5HPNaTVvRKqFX0CPTD7KmQ4bfXG0FORC92WjAqbDE4Izu8esSnWMG
FnUECKskYovDdOFdpTJX/obbHyM2/AJ9TDlxisKulmPVFwK/OvYK/oBh9/OfqZSr
zQ+5fe7ZWaizDP0VlfITkmhlYhAYeCv7/1lpkiNcPYmK7zRpX7x++fhBuqeCoorw
kKEAU8LfQ6bdgE8IuwTh1nbxR81dy2sDmdWeh5oQ1uOPuPTeMpL27cTsgahISAN+
J3+6xYBN5FPB+8J4Y2BKSzd0nks2xbUDhz2LgrslN/11k8BdAi+5TnXRml7GEbGN
If15eeosIIJ02M0Dk8Rw9OEGzQ1QDQewzaLAoJEdt8UL5eaae6hMHIXRTEe3ITiP
oEhw1i0PiRkczs8xJIWKDLhe6UiovIZH98qBrDwm82qC/5MGh2SBa7qlA3q+nnet
Hfovond+WZR/lXqJhm4gZN4tCtRQnZC8LOtWMONnt/oKeh5T8A3LntJuJJtCUig2
WIYNRWMfEjST3r8Je9Y9QBQ8Udba9NkZOVgo7XzZcNuOzja5O5NL/Dev7aPqpcM+
fZvO2DH+coKhndKGXY37uhtrN47UxGZJx8VJ2+PkTICLwbO562Qqjh+G1w+4Icqx
OT451xO+cmS9R/ATS/Ay+iV2FakzzqSVE4dY/o1RtnXiv1N+TjC4XMyH2k8wEFX+
lZDRqqj5/kwvPiblJDTv9nIhjXoeH6OwmlMXV6Vu0SuVbLsclcP2VpUzjItY6uy6
5/rd4SAs4cDToP0cn/rsrPuurMMsWGIOdJXC6tDZpEwqFdaA1bRVaJvAq/qvzpcR
NIk6D83gJkXgVnisoq01a6JWzodvplm4gh+x2J8maUdSjRxAH6IEr6IqGa/6Yr5h
zLl43uROgIjLz0SUQJTYRojTJT48iTV/OGlam3AfdR5jVvdVbYqS05fku4bxgpyc
Iw0E3zmOvSnbN8r4z7BIklbG0ipAvPkQ3K5/F8Kd4eWDS0Ys+YKedrLMYzicF64B
nekZt7hv5F28McEZEkNnUiY+/xUdltD2DFtAPgHdo8S2vKATexePfiXWXq7NKUOB
TxTWU9a4Fxd1NOdsURuCDNeO2qxXfJ3/bTDLatZKsuZg+ylqzC0zKbKd5AGTiL9u
vulbLl+uSMtXbJNlj16kxS4A4aV/iTiEPhuMNcQJN7gZE/UMnCtIa4U4ogl2m8+F
uz96ZcN2s1uumVUeN+jHqnOwh5VuBIimdWCHXCHxTozKXDaYXGmo2NGkdNqsOH6P
hdR939slAAK2i+IZfHgHI6WB275iv4nP4BrXUv8HxgG+17H+YAtCIGY4+hAZCRfp
1Qr5NL3TrhDlKS/5INe6LtQrzLmTxSFiXOy4LvRldI93BNCYQtDCsanW099WrXC1
8+l4qv9qkS9EZHmsuyQWDqmjHtTzuWTZssEVI6P4yFONWflojHWMeGRrUQVEjoOY
ojq9IjXO+RgoYBclRAOUEx/5iylfinZNCuV3EtUk3+k8uGdzJokcaCXVEkaVYpp/
fXbzmBPiSN5azIwe4wdDfPgQqUlap51oOui9QyNlLH3vXhxnjy4kfPNZNhR16n4I
CXsDa7Rfql/vOgOGS+GosmJ82Dv4ZGnb7Y9Ctp6WPxpxYs7rPWxhZ+Y3A2pnYsjY
YbAE7RFX8lNllHJhgVSG42muorMqXoNjt0T0O05WaHOCdHoVQnFwpUDOUAGyihHz
v25epsRmRB8RVhpCmwIQq4z9s7BL7z8dYhOEQLGt5swBWKt8+JHGUCIY1lfy+kan
jVR5udz54PYGGniKqCqhSqgqzI3Ri/c3gjqVAGaS+GTtgN0yYUncOqb2ryVyed5C
OyiTRoEgnTfKw5z0psVxfJf+7KTc18GQLWX7rX9uNAkkcVZjoPQzyAMphpe4BkoU
vA/fFML4F59EaydBH4fbwtmbWmVrLQ8FafX1jKVbKpE4Vk5D548uDhA++3ekoNio
MZOQZp3ojyAktucP+CnDOa4gbFzbBSm35JAPiZ6pNRdT3kQfbe+MjfVnpLIeurcx
2EcC1P/klIlUKoe39fQ9nhgDa9Cf3QswBJty31JOWZtBW9xW/rmPNZxD4eBxX4X2
0odcg8tMqcmUQRgt9n0zzQY0dNwMq9Jp0vLzSZif8aMKeVg190OXlJxp2Uhrb8+A
7QqN7QWhhD1jgtbmecNcS4sOkwZeVWRkR1lZsT1OkERICEjDpTnDYOkJ+PkgNh/s
WXIRmL1SaHcMNknKqqydygGxBpprhMMU73SpXd0IyFLGj7nOaGbFZcOBM0zNPoh0
LEbVrmH9O6wsaYx1+kVxaI65i/CQmToeOFiram19I3jAt7GRoAK+b70r1gRBaxIt
n6DOTbK2WXlR4msa8OrFz0KRyRn4Bym+MPec3TPdLg3unAzIpacLso/xioX2Op31
D/Y0j2k5CA27O0snNBV/g6erQ+UPonpHphGOj5pLIKJLgx51LNfaCv4Cdij2KX52
QbcIR58CO0UeTHoUODwDMSHXx87wJWr3xSI241Aa4ciIQItgMb35rlnSm3rOP3rc
huQpUsbyPG+Y4VtqdHmh0As7XDSMLEnrQ1MgICsjnETca5yW3Dg6+Iw1C076WB4t
b6LdPDyH++DPJN1XMMdCChvS3WLfRBXuwFyfZir+p41u1zU/SrMHpQTzUZALU3hv
JcnTMi9ya4ZxFqwugvuJcbyc66/WuRg03/8PauT8UvHs+kBuUb83U50xOWLsHqPN
0JO5ret0qp21EU0ILeH6p6gInvhq0RCE6NEd4UTLh8+O6vg4ywGs0OU+IpjmJrsw
629vPjbRBtYKpFWHoLnnUBFyHSlY9eaY09yjif6Uio1gBpeg4vwW1usvVDLk9H24
namNtBCrqXJddoE+XYbJX69RRDxH9W2M39Omj4Ss75fPKeYiXHtqFGhtie9qxTD0
q5Qlr4YmuOrVMniFNpI3HGkCmsXr5qTlmRttiqQXOCSmJ3SZSTslpPsehjvc4x9Y
kI8Dk7r722LAsGgwND/5Bq5vE7jcrc+m8JXOWCY5y7+9XZ9QM18XFVZGHQOGZYxN
3bqQwGnRM+kPhaTGiuqYa3hVozMBr4EQLR4lpJpmshi98Sr5s6sJHXXaSr9wYvBe
6KCKZK4khYbccYB+UcmG7hm/7n8BfeahdOokKl5xPEUyx7UIL2ebLkWrxecnV3rR
/9PxWkS4p2Pblj8BKzEN6JgDzW38QFkcVn9wD7B0EcQNDWOrEXk9vL0OrgR1ZTPg
z8MB3PIla7BA99w9cTbfdeOW4Q2I3AXi9mKTZPj9BSZiKya11MrpzKNTwhgIPxio
QSQvWYUbJgRNIBkCv6zUmiNZT269OX+PZmUS2u/DI7g9fCD74ACRyJgZ2EOlGA+z
rC6uGV9ZjAElcDCkuSbWGHkfZCxJ5xn0OqesUcmIW4ABPgry7TryWYR0g2pgUv4M
KRm0O2hfbLJzS0hLExl9vG2sQo50kZaa/1xjJSwZetb2z5Yt1xEq5zEI19N2hoDd
ksD5Z7mP9d/Wi7gVtssW+I79wu3LeaS81jfNZsm5GlIWuwwqCd8uZ50FHHabXhDM
61HyOo4YNYOZGxtKy4bHMfOpidGsBTX1Jhy1eqytw/2L35HXc6njbsCvUoGx+bgF
dMwBp41BGnjwRBOeoChtwl336VUvxTr6xoAvj25OtsWakoa3MRR1at+gr+RdEiJ5
aMihX8vRo+7PJ2XEOW1aPlo4J33idtS0TtiIAX/r8TI7Lu7sy72Q4jjDuAJKwLKd
uqGI/xymDr0WtciE8z+8pC4tTlHHTRiZLRfBQm7f220eyE5tBk+S5do4nE8nDYeg
C+JRzAofVA+w8/tlu34IseLC2ozfKssP9m2NT5bpYXWlx/D7hyWcI95lgvfqnwQM
NYXldpoarX/+SsXC/0PXeJThW2eJL4iP8KLQz7ruPYEfXmCNP3ypZIu1ZDpESpGY
6oS/qm9FiZAXnyKi5hviCX5sCLVMpDfxKiPNWrjYiHPnLFeygCNGiPzo2qj7pCd7
+vCJynNhekCRS7BiVj5AhJ++6Bprms4KtLtZhGdUMQgm/2JUNGkDk/3V+JAFRSOm
cMOS7+7w7j+mgk28MGsIW2Gr2eFiIGfAzvDMN7fIJcNuRLZR7nSit+CyHMT0o1EI
m5vMdZN9ZlKWjO7Zo617C5IhD15ku15AR9PJtfg7xe2uNlhujGDI9bhzI/TrN0J/
VXHokZ6F4fzW+JrZEQjHgv/hOS2KiaNrWVFld0O2fcH4c4sq5Im20bAfXTblJgXC
1Al6G4E2QG1eldy2gd6mkD7NoTb67QPq0Ylh8CEDAppkLh2xK0D2rPJ7JkvoMOG5
EnpgnbLkjYT5tFjfxO3nfgTDHZIpD9ELhE2KcXxPbt6mxmu13LTnXilO8Kb0aziI
p7Fn+8a0suYTei1AhHAJCab1fo7fFAXOogkkvQOSlaUc4I1+ttfyq1HLZPCM3JNX
7rjr1a8e5E2CAhGZvRWjBWE4RbqAlu+vcWODLz8QRZsPdX7gs3ImnOtFmtmUL1dU
ZOQLVuxUll1jZHMOf3tcBr+ak52PEgzHjLhUEX0yPyq8QCsUdFxIwx2ddufn0Dac
HnpdvhGhlyIJ8EQujeWEmIaFSbUapF9s4Zp7Q9qRIABsg+FQNE+poYVs8H4lssp7
cadFBlYfuWbiRHpBF+CUrYUiXNqlL87zvWtbeJAnRzLbayPaHdJax1Z+jlizmQE/
sA5B4zMocV79+2JqeBr9VYF1E8DEOvWOWygLRsE1Jm7vrrycmSJYApv3KpVG8nRj
Luus6u0PI+oVpp6ilfPSn4Si1SLzB7oGPtK9j/Fu+b71BDYSRXQ0p/IW7ckZOrtm
sz0C5zPejXhGzOnTYIq/iwyVGERRoH8x4p0W6FAIy/z6QDDRZR0Uhp4TM3/Yy7gC
rof7tpFOd6aRo4q3gryaD2UFizm18wrAgdad4UQWIo7RgSkI8GgctSb8twIQVRxt
ACbWQ5jbmymZu8thXBuOw2QHsQ61jE0tFbOLaX3Krzxjmjy4o0Ax/CMB68AFESDj
KABOOuUrJSGQcoF17AObRNbPkzwXZrONubnI1kcNQvYQuQOZCFn2L5JCZlQd9er5
tXcDskE27lx9lOCjhXWI3icNRzeQmGLJkJSsAVDKe+p3XDoHv/g8LldZsFWjNuY9
z2x11ksNJJvyCYqwokqVzE3fk43cMG2FloUZwkbJ5oPqyLAn6MzMGhxfaVG77IlZ
+qpZIe1/1+NMFmTRIkRz6ASuXwxtOYCRuMYicxMHTsk+kR7UspXbrvYGWwtkZLi6
oh3GjhXNku1yBPwKSVed7nx1bJbEo9dqHCi2TjnypMVpKa0oEi1h+d/FmGUpEhGr
krVMhBLBs2RmEir+Nuc/WZhSX7eFkxFUWbfQJbDFReKsC9UjiNdoGXy4cLieVZfO
IxIVOqaj2f+kPFu5eia9ArCjuJt/alXKB+JoS100dpn1czYMc6K4wMJj9wRZ5vf8
dlPLEe4OhpJ3N02oR4XjQZKv2HtHYvvf46/iNSNDf4ueazhd4qwrX2f8HKYH9wQR
3A9MW8bdkqzgPjnOay0EDI4G4gi1Nkg0Eq7qWt7KppezWKTafFv7+KI7BLY5AGlE
cnN4+0bpGF9EvXvzOrhmFOOW47YUN7S+qMFDOyxwjtT3+UWsVQRrrOh4zt0lUIEH
YRsW8VRTk77Q0ifQIyVpqu5OCFfz2JONqwz7vV47sC3YEr+danVfhJrdwzqGXOhZ
1OaK1TdrAkbRnNFWyPuMjQJBAtgvd6WvSIs0Wq5JFAmwsSxKGClklSZflLem+2/9
irVI2yGrA4tknJMsoVG2JFmpd33nNZAf/71GZ09jXXK2eLJlUnVRS5XPdgx5tCC5
49G5qn43I3Gz71MWyHUcARAr3P2aB0cbpppvvqLyawoCQhfQZRSCHL3nHBpTEFBw
2cMAn9epMHFjy9diConUl1HaAcEZh35I0PPBgQm3QsI/ZQo/DFAdGcVz9IgkZNTC
mmHZyU+/XDvaVZiSNSAFSgaCiUb8FtOBEhWigfL/ej7S/4T/fiVm0upOctgXQ7wt
oa4c+gGywI4EupZGe6NaunvtU1b4qJ4Y9a2hNpnu/w5OvWmaPAZ80NzPmy97fON5
cv+DU0XE8qtX8i/kWJ4/6k6DH/pKnUIvAGmTeCcdMLsQCw27PdBOQDdi15Ea81cA
NCtIOek1s9l4KdXwAaRRVVOZQUr8Fev72UXa+5xM8xbFzcVYlw+R5ce+ahINFSzM
qURi23o/ct0UJHI/kyoTsiDZNV5Zz9NcEJSgZTCZD4s5AxWGeiVBj+B/GLxZLGWr
35jP+YDY6XZdYuyF3QFrDIVIhIhDyLry2D8VfMfbHchGj8AjF1RKsvS9Q+cEMrup
HWzKq1zvVTklz7iT2Kng8bApYpoMIzjDRkh5U3NrN4kvx1nnpBPZ6//GM1zGGPIZ
9x3fRgLouaIzDGXfpLAPy5Trz6wsA6S6JMxdPYYi1e3FskdMQZWUxHS23amRhx8F
bzsk0MZMJBkAZNrwNQQWEK+K+GEGZq/Gx1ZLkd/xTmoRtQgKiEX+ylDsHDpg5OJW
W/EWAvlH2wCjbwvH8A9ofco3wir2rJjYohf1I8aN5OkhojAbqFmknoDeCexKQnGG
3fd8kvHu69u2VQ4tJM6tkNZagxCjqDeGmrVi7hflmN0dTgHAakxwwxNhWKvUbUh3
IqASiwm8kJmwmUaYDlH7sJcZsj9vsoKiA+kIlhaxx1UDD+SNJix1WOtrd66xCJd4
kmAJM84kt2+SXFpGX+NwUG1FBdM0YX6PgB0ylonqHiQzFYgmW1Vww9uCSA8og8KP
LospnlEYWMYdAQPPUGLKkjAAusiGoqiiUOXCr5Z40BO/vDsmArQ9wuSf5M39U3Jc
nZl6I2p2ZkgqffBp8sOopXSw7bQ87claMX7aAUyYRqmNi7KNgg30RquMUTo2DOd2
AsSIZ+3mVpdUInewOg+3lQMDdfnrXrNSQxV0uuh6BEFmQ3gXqqNAAY2867MbAqXO
Ug2/5iWSqxny6LmzuoSG0L+BcmLCYu432qVad4q72elIdtdO6QsxzLo4c7r9qA1O
XgL8cuIgjTf6noNdTm19acmgYzxIxQT5A5xjsZ4m5lJ13OJ/FSBY3zGXENwBqqHi
M2dCAathvJyZQ4HIDjdcg5onyvY0zLOlw04stQeGJmd45mpH3pC6cQuwBStgZaXK
gAyGl7lxDjHCF1Ja4oJlajoHvlvx2Y2aoTOHYUO8pitN1WO7GjYlyyO+sJy/qWMl
9tmWw3lSJYBKy2VR9gHwFw/oPTHLH260cVTbFp0AVCPjKV4opWtftSYdoGip4er3
0OKs1mpSbXi1rMhzNuo4W1wWjLAJQDGLqs3fhirikEoC/9/4HltQqIeeMEYMg8Et
cmjMkkNUpT5FYUxMTegbIU/GPwWxh+3igqKbOkgsJNSdOtrWc63OfdxXnzgtoIeS
fz5bedE2VANqG8LB3aZmRaxDcz9/Xc0R+pOTE76lslxTXbLhDrBCYmmh91s0kjTh
lFXDhv9EBlxcOY/jW2cFCjZ9XxMAyVuxY8hKrLa/NNDchkZnNS69HwKX6zilMPTX
PrC0AJVzOhH17GskPlufzt/fuMkjC4/RKyxQqnepfg+HKSu2SqVPZ6H4mfnXvpVi
lFS7wISkfPA2oNpwTdwHggl/HEKdjbrSZPUQdwj/59TQIK7KSjmSDwb/MDwYixxy
4i0Uy+wnWs2ii+DRzPUguhKXUP7TPo1Orpcyop59PZn9xsYSAPNPQuDIc2LsjdT2
qcN5acqGHV2V4zVxhKbsG/rwQaYWKKPii54F0DKvE74W27yskh8efc5c36ukgqZW
m7alSs4fHdMM7n82AIVXEWYwsjaBvFsz4bnmgVq1RVeR3vmZyujGN9esPBSt/KJ8
Lx+QRRr1z3HnTVaswKpC1YqEC/spO3GnB+h7ptcM/AOzAadozB9fIYHCDG9UUfIm
3QaFPL3jpxZiwj6KeNJYxF5WsIz2VvCcy4ZWOhPt+5CYuJZbNuYdwvzWdkUVCkI1
rKaABTgXN9K2/M5Onqs3A4SmAN9cQMRhOwxCM/tqcYcjO1Xx9+23PM3AC+MikmnU
ogBMZkb2bZDVJhdABo1sw7FnFLGLAjXCPIc01SO+ZmpnhNw499K8uRE0RQ2pU6Mr
+XOsv8FF/eVIBygnjBHgCzPeWES5kYbtjKskelcikt8n/HiOgY7R91noMu+jvV9m
kHCz3joZHBlzP4M/NPPb/WjhKA8+b2hANUmAACtJ7kH2353oVx+/JiStHECmQeHg
tT7ZVpBelenwsgQna6ZAdor7Vw4uhmEqb8EVZtG2rG/4QRslJ2LNtVOk8MqxitIi
JGplK7DurDyNeFsM8GeaxmyanoeV4+mQ8X5ZYjVGpnbUYVbW1EPzNW9Jtwhqn99S
9bwZ2OL/CUZ9230NLyUSCDijHQsvDO5sLnqguAg7+T2XCTvUIUFBttyZt335SW1S
WTFAuK6stcxtsmagU42nFZGcqMCbcDy18S5mIx5dlOSFdmagGWDK4m2plJmjJEky
av3Oo0z1XuJ0WdlAgYujqlOsOiHenTqYxGZUAqDCsYyt+hcs0UitzQ0VXk32Owbz
ATu6E1OWJZzMj/0LAiBsU87st7jmBH7488BfFXY0WOtNEQ1zvKHyafFzWRR/oh6q
yiU8NuPiq8Utiq7DMtEPQqs1uos/DmcZ+alX/keQWyjDEKG5JgR8fpfJhhlDjvBX
vmv26bMaESHwCJACo4HMfE/nYi9IMSpgT/qHdT5JsedgcmfLZf3ufF4Fdqgore+Z
r5axMyGHjXp8wF0+x0/wI3It1hYZMpSgnjE4/q5OZlLn80Ytgb9/em9c9CXyLsS4
Tjgwi6/ytNywMzyPgxpWEVzkF/fSoL5IUjQmUUwFfz+oTKNYax80QU6AW7c4M/XW
tgmaZp2XHGk0NTg7KfNAa4+kfxp4C3NVEhG+gT/RUyv7hThZewpnOKwIGf27mNqd
sgFAcheqnIyclMYwiRqIs3wKruXFwBbZmuKgPLkWLZ5zGHTx+PW5Afkfde7iGu5X
FroUB+fjYBbQJcnBJHPsfU/4T1bhtR/7cGe/z94stD4mkkItBtb9l9cNnpwnrAI8
zCD/2ztmHqn+obwAC3dLOPYLeBWSgvVsZPezgOSYHqWIXYIOKQDFrRcmPxJxFYWz
TMgvISHPyrKoNqkHVr06/bBeJZoU20vdH2uNbUQRitYdHoffH3THqfw0AQmVqW/9
GhS2OFUioLJ9f8wzOn09IVqzWfwQHSltj3XGYpYm4SE3GfK2MF1R9scBCdwU7PIf
3DG6LX9pudyB9ktZH2uBDJvm8X6OzRWmWrR0eOTl/GskkCzBNT9kmKUuqfZjj3E4
iiy4vGjHCNli8s6wTE1Fe0AU/IzEhI0Ls40bqG+991JWaYq74jt9sDtmkbfsIuja
jPqBEb8sqLw5B7j7H2VzBXQtKnzrnEK15PR5buua0G2k1/P8cGt6/OFGRzWDQO79
fvrt8QzWhG2Pu0JwhhPmeG4AzCxuvFpzxyIZUIhVEGIDRtEyZXVKodvz5+Lw5n3d
LB0HQdDtHSXzir9MHVLsLbFWGF2gkTH6UxG4p3ZkaVAamBvXe9N0vUzS2QCjaHuV
09C3YRe6X4QPujK3LcUESU460CRZ3ikdmbkowaZvTH/x0dr2LZ78pFcamzJTZHWT
gLcw7jsNXFo37fiOCvFNFtKjsGL5G8Z40QSf2F/DNzoXrOS3yu+fi9P98yqygjdH
2kiWTnMMBXo7DXCo99DNq0Tixhbxr1rSBhfMdwvCL8UbiELGCyxB8wmaNHkLba3l
aOfVbvq7VMXwOfeEpDqzuK6PstPVZefsq4uk8oJwXWnHJxBVRs47QtHV7mgH6OnN
x4kVyPrL1+l0dlVZopDxfWkKvy/7dI7yqLtCFlhXgX4Zf/YipjchabSjKMpGra4B
YdrYLAxTal1Z1TQGtR6ff1TmAPHPvvUijOqPuwIOB/Wchn4i0ikLNacwpCL3iPlq
za/tpqXa3cUEV3Xev7MERJjjmz9/CRdaDXRFZbD2tuja4FafLN6YQOsc9i+FqiAT
UXdayhHMaK3pKSM2ch2puYiQAusGVNmAP9PNokRtShUHTA5XzYCyMUVUlntXFdZh
EFxDjjrii3u2L2yNUFE6EM8U1zM+DCCBu9zVm/iddJGq4TwAh+kdFqERZLwvsveN
h7/p3AOb6DXOBVRbFzyK+YdosSVR2JKk/i+TYnE37IHx2R9xx8OLI2RozGu2idoW
169LKIwAyTVIcehFtTAO8/XM4G7Lgvkm7l5hhOe1LXT9IQggbQpvQk+72X5ez30z
NH0NCusFDPGX4gCbTyHPnBkGESMiE5sfgCz/qZ5XDvsllUEKR9eBe5XUMJqBo4TB
nIKN3oIv+boaln9GdGW5BHu8R6Yp4AkJJy7RW8rD5+RVWqUZUANz2dOt98gyjP2u
x2XC8Qj0UvRyEDTY30vGxaiTWt3fCj46fR/mqWgdrbfMFxNzGgoo+YN/yzb5Mj2L
pBMZLYzk+XnfLzF1Ti2HfRcta3LbaKGOd9VWwa/ADVkYlS/BtGgRIVvc/htRZm1n
AWgqLxxa6FR+jK6j2CMgzISt0GuqJahcGUYI+P/JC0kyTLZbUe/B9kV/wqjKVdVM
G4RZYUf/SEGy0W6xhrg98EHS7xBASfvwhDT+3CIhQ0JIDLwGsdH9QkbSB5lx2Yv5
cBwPwDIFM6wme9mH08OZ/rbPcK1qPdiy7aNR13984KKCGpdljhMs25b4FG2MC6DL
iTl3AGZVMyvJTInh25NnJR6YsxdkOhBKlXOAuCe79rFiZJQZ2YM1+g6psK2j1gau
t/7mcpHIMxvrW7sfenMHDiYgvdiKBXvfGC9q8xl7+7GMiOYuxVr+k9ICLzC6U1Vv
3xSREMA8AU18OkAQiahlhWc7CL+rNga6sHnsezoPCOVWW6bu4zBmdbrLQk59W1Dv
y1r44Ka8uIJjQ7+64e7ZnhS0fY+yayW1AcERek3kRKGS6dSbMN0gsTc8QFA1pWRk
hGOmxpUTFh4IIBP/jVbcr89TfNH69BT3/nXDqWTTKLMMYzFTPWyIc918U9Iuc0jZ
gFR/6tzAhZT8uPOAQ5h+GqodvEu7b4uOyeFsEiNyWUeCaQD4nOV4d98fbaNcFlVW
1n0WczK2mszLeygKRE+9u47OPQC4KnAEaGWJHp1FkSIOTPgtEIMEXcTx6RAgNURT
t+rITn095RW6wJeUYxubXOk2c5/LECVEgxyattxMJjbPOfCJ3zIMwfZwC8TdfNAm
1npjpoCx34nzAnOOR5KflI0fhgzetLbBaywztswF6M4b+SgK7C+bj1bB4yEt4vbK
HMtdO/zTA8L10L8N7T1SSM5H3JgnOvfboz7FTYe+69bl6u9hU1VGo+k99bCF8gCM
zuRf3Vlvwap7ICqDW0zuLOwFdurT3Ph/3K2Kw5K5ZCadBzRQfQt31RKNeYyejk84
5GuOOxzvrngmUqnMZ0l5gaIaO8Uj78YGK2m4yrSlZlO/mM0GxYJfNgI9x819k1/X
3/BVEsD7pLOi151acTPWXtslX8hHFhjZsYe/MtiSdalLNBoXEd9bSoiJN7TWq7tv
5O2Gl6UVedWHz+hvtQS1jlYS49Q5rKmhWnAX1yvJbM7mA76CbG0BNf7H/apxrV/R
qBQQWNt7teOd6IVy0W8Xd8WzzGPQctPCYbExRbzyV7h1aQK1mg7xApOxF9X/AQKm
wx5TgIa9nT77Z/LMBWUPbdbiV1euBFAqdxqW1VBa2QScRqxkf+KQsHXSiYp/tDrb
XvSK7CYTLOXdXZboyhWcvNg4CTK9Xj7PoZS3bW3pqB5I5jiByVJLAW3QZeNFgLlY
DKyQYl2l2bi8KkfupNhVKEfI9JboARyZ00O/cx9T9YJEk2xKYuB59+ZvUnv3dXX8
EaZmonmcGJ3qbXRjm0lWA9TpsT9pUgzf+/XP52ZJoHphyz8Mrx5rr3uQWEbiMkAj
+UqI0xB3o+Q1SgKs//JCagqtTfNJv/6Dptml2LOoYDURGRHqFOE/DYxN/iXNfYIB
LIy8lXG6BMndyOr/6s81XE9MyjrsD5wbtr0q+oZX+xeWVwTWyhyyCkXJ87t2aPVg
wLbBFh9Yn3uuGOSMlsPSpptTg1DoY4nBAN0dSrEiIINsOV9/06IQUW3X6MhJwroa
Y6lGynOC7xYbMOUgCCftFQ49CyMkX9m+iQ3z6VVrJec9dYNEDF9nq+TGT/gavsc8
B538bmxgA56I+MitBstCXu4fYgCWbvl6Y9yIqGfr9USqSmuWhW66Mzj8HcpYUoxm
idEZSI0f84pU/XKT2qlobuKYXZo+zkUYa8jCUouKUPE6sw008p9xfzZcy1IVMCHe
ZlI1FUdtfkMI2GW38Gc3RxYAhzp6yItBa12IkM2UXlfXYHICXLBvdLQZZefGEuva
u6lRpHXkaBlq11RFMR6Gd5eVbXt3IKUeznP7pJbSDgknpjB5VJ6N0rhf6Db4oOUx
m5pMR/P3WeAmbRybSK7n5Dt7RjMF0y58BbLGcoFbEHavQgp9rSydZUPj+Ap7F50J
53OX1EwEE8yg3rT1SsX1wzN68LltwJ9/xjQdRX2Ko+DegnXjnma/Sor/4Z6F4CUI
Eeve2L5hEuV3wBb93oLjIPHqxWmFbQ/ZBRh+NBO0Tqf5hdY/kiSmt+LxjmzwekU4
Pv4fb6G07Jus/wG9ZwOvzrwanZXppjX5/Qq5pMGYxXx1gtG/SH5ih5PBd4uZi8ln
I7x9715it8zkEWbVt4ZlH5E2ZkU82iUabQeU62+eGj/3c8lc5qXn2V5S4RIKRRgK
aiMKwKZDiecYTZjLa1dRRUI9niKO6pKvjdDjhXbsxI5UZA4cANYckXR1NdLz81sl
AR/vztPHu3z3WChL4+wM+GvojxTEPpkDZEG5kfZJvTheDIOdT5/NMzSp674/XHkL
mQ1Cz0+LxXFKDbyhGO5eGtpmiZJRLX1wzwPb4eg1I35dtt9Y2U6Z7wyfliInvejZ
ZmjP5JDe//qqa/4dMxBeynCkT12pa+JL/to6fzqWELM90sQ4LrG9LzDy6G3MwQAB
uo0kla6xlrdJxo/hZYRrL6E1rSAAwjad1UE/V2slNlZTzOAL5hJrtDaqrNgdCE87
3Vt2qUUVD280dwvjohcl78vMF6RS23GTAeHUkRB6nMgb+5eB9I8KT07843GvH3Rd
UC78rrJDVFC5VJVurGLjdOniHOQyIa4ZaHvv8uF285GBu7wcEg+ig0/VCuduUIaA
TArtuNIhh9t8NcA6DtQILOr5qrQyw709jEVoNT0AmQ4cZzX4MivUueTkufwO5OU+
Vb+t08rw9Ki02B2dehLyTWt3owih+Z1Bri8+uQ+PHY2ScFoLba5H+xgwV2d8/BFM
qfvEO2Y/ufwAQTaA6bUZIXB93Ze2/sCroQdEEQj+eoE76te2t+AsesrXpBoR8cYL
rtK69TCxK7CH7Pk4GVlCDCAl4PbynRXJDMOiyyHGf43i9oM1Ug4QO6H+LRQKpxDR
mhkBflgYHi4otNcXECHt0cf68MinkF0nQkoFfLvrJRGSmy1Qdipji6aLjcSevAmd
jtAKBUePs/kZq46Az/ziK1HroSf/ytByLj7SavLlMzcqjJ4U+I+45RX6lc21aVAv
ZgW4/VudLQ4e9uqT83JkUb1uyOf2itfdXh/zq+ZlM7EH++NmOgd1xo0XsXrtfFc5
Ylx5vYmyRs6SI5EF9oq9YYkz251cUkzK0ghmuG0Kq8ysv77j/f6cusPNf7hx2FQE
okzlDTiwAByq6jouUqYUeVeBY/LlNDuBV2iPpfT6iD08IG6lQ7rOEHtnv7hE+aV7
D3qdFVAlTffGugGXg4vKWt5alGrqnwTUV6wGn8qjlmusey7HZnYQz9ZTCFBq2p1E
6hm7KYHExwdffKwdb18wxxDEZPsTbz2+ebrMDEw/jRKqZGDFYHip7I7aC6Jz+v9i
La7VEnKzJ9cBAUfkNYg6uIC+x33x4Miqio1Km/idM0seCcqqsseoz+D6lTFnGI2h
M2qNx2QSl1YfwRh5iQp3Zadi8sb6u+GTmRuOwqotF+jl2ymo469J3uKQZ2u7Cvk/
7HOCawtg6OIpFawqqTS474zNwPWGQhlqySHiICicuR3P3chHrr85UWs/OArPhx1g
jdatTEgfqKzEjK0Pu3fOy2CLpoHKHAB3ij/ikdbSroMzNoLCXV/pVltUu49Fjp3I
nRvXvPNypI/JkiKqfKDrw4c8rWl0SAM1vfhpxG7g1HNWgxwj4V8pBGa8nhAQP+SQ
/sNsstesVZPv8gswizynjQG2jTNGZiP7/xHIvdyRVMvyXx/1UorV/7xzxFEM6y3Q
fdoT1oYV89qQHRZl7OJIzzcG6ZcGym4Rs87gKi+s/JloU5MF8yZzBRVrzUx5/xKF
bAQ+zGhZSJ8WI0aWnuAxyibIA+g32cMbvtfWd2NvUkM3drVfD6AujTj8/YDiM013
pANFQvX95muzWf770nbdwSmj4jYQhYPWdlDbBZK9cT8G/vv+pfMjVNIG2XA7jlF+
LBRZimXbfXKh+QipZt4AoXdjNS93snoAPT4bjGG+R8KtuSoQZpnGACnYv68tV3Sg
AMtdvLvZXqrUYlyZXkeI4GoNV/GZr2dZLnECRxEPBTJCjF+SAcT3inQaAGZFuNTi
vOymoDwg1tVFWFe5Gyg/gfrxx1eKyRtntTgbeR4YFFsiTaCC7scSrYAo+LA71FHh
NAHQgFO7CW/EK1O9a3KAsoWzy5K9H5Fez+zdqvV1OL+fiI/00KNGWyjVkxSsAWpa
jBWBBfpML+yOA0vqIC/WsK1brKekZdE+qEJZnU3bqx3He21ou8uSL+uvx265UznI
tpzAlkf8Hb9DqfbqHAhteIBZibplw35zMZuZGcDWmALssEZA834C72Qb3TaV65CP
l3ne1Ju8smalwSUuoJKN0S+NOhdwnQKq+UM6cE8aYP1rhgpibLYVrWs65f5Tyx+/
FytMVfhTyMlrkPCnu6CLookrid7MMoO3zWbp2hRq2d8z4rb20ZgvMx/xKAyY2Cq+
qtkyivz0Ey8LzDvvmztm2ot6u+ZpkDHQ7E+uheDiJwkdLxsa2OMl3M7PCNVJ0ov/
4hkSy7OQLHq4aFspWFol79YXBjFEO3C21YYsnYpiTXeyv7OC487E7Eyp7+Ef3iTf
i4AaDSEj8UF8xKf/5tr1NKO07ieaaksmvzOxIJdQnwBQIET1OxorcgESTUj2NHKw
EBWvvAthj0gKwZ04R5McehDwVsxFySceXRvgXuZOLJdPiZtcS4X4b2M7XaUnFR6L
9rubHl9dsMLGGyhzRZ5cCA5CBLi3n8eeto9SIQ6MD7Hji3MfyMybT7n4dxj1jpkl
yF65FX8pFtWEMAuLS3NU8Yla3Debsh+Xl0eEsSAFyYuW6kHUL5NyIVcAW8VX9GlN
qVz3Jq/1ED9M6Iq+ao2ZSc/fg1B6zRQwHgXndIB8FzLsSbMMOTnVWmptfzKzFj4a
Sg4tCpEBSluoP3lNAh92jIzBGP/6ZpfhFeaknme9UuqA+r5VsxHBaTHbFwYjQV60
Ui2r+XrowbxLX7H7H9X6UmP0W3BkIa+lPWCvVWc4uUfUVdnnH3GsKZLvVL5iupF4
yDb9VYTICF1JnnnU/VhNL6MGwspOQoSm82PA9TKBg47ZFBnKxQVTp27P6C2Xsrx/
4Tuh6ciQ70wQxnxKA5aZxOlY9UJeKOKwfFKIVFtOpDwpyXtJyFdrHgO9IOBLI6Sz
0b9kNXrfnbPV0xS9NRy8z3Fve2eSv5gq46tE2INDTDhJo1rBeSdXEYV1aLYuIg4A
VWYEDzRAhR8g4vbKYdzhcXZ0b85F5fZUMHRxs+ILUPc3i/mmPNKyTIa/2OpyamaA
dtOFj3oYuK/913C9dyJ/qV6hh8fRwwBUuDyQa8jBUUyW+P/hEVXx7Z/jBpueuyeF
0lyug+/VSyfqWujvzpHMKpKr3sXKwIZElWSu0gThxSbCKrde0T+W11YJlLGJAQ9C
KT8LL26I4V4nnyb2RsLGMhduJaodo8wt7hf+8aU7gbYEDunmbV1K73iL6FGjv5bG
NlySSGLTz4uPYKLTqFQrWzzbc+KvslE2usu2eFNN4sAN5kxUmxMWJAyjG0Ip1pCt
AS/p1PQIKY+ALi3j68tswzIIoBse6KXXpWUSYlP1FiKn1Wq3ynR+71ZWoKQR882Y
wJLcP+//baJ6kueTJX5fD4EVE64zEwdrr+NLMB36fMIpJPvg10YyGag55ntcWDE5
5W3yeF1BKfS/mN3V1VNqEVQi//kRXizdJYfrLbM8f5Np9fB+k+UESMDP6Fhby8io
JB0UJSv/SWTlRCqWh8T1/GAkTGQ2BIA1wlQxWrDqTINroz9dydoRFFMI3o18Qxk9
JnMEZrq9D98M5bpMAA1tNEcDMLPTi8gKwjf3gvdtaOdRvWlEfkTV+R8Zi93RVJXd
c69exVDQoNeGVACnw0MNwJao9uB6o0y/9yqOoYf0HGGGGQSrS3PVyGhLdfbqvijG
WG2BQVF99aejhJN1+Dfroc6yk3Re6oJLYfYzDs1SQDQBjkdUWJrTwbA3g1KrHyvi
LHNMa4wujTZO4UNGwtWp6vs8FAY2S8lBKnLIiqEQUF7Khwq0YwDT29y+X3NqQ9sC
JGCn0of7imMPLX7wCVvPc825hSdtIO/e1Ls6B2sKDPHNNS4U2Z8NRjDR62ZWdABY
fiWEKtnPaUpGbh67vsSTUk1wzzh+dmgJ3P0A2wdBY/J7Fic8lVRJf6/HdZ8AvUxw
AfkP7pSMSG50JQYEpw1FM1fdXxmwL+2cG1SWXPIbT2A1XPzmTGqfMsSaEtUNIcxW
5di3DIC9VybHT9TGLj4i5ZwV3jOb96xsIi4Keml+4wiHCyf2qar37NL0tLI/T6z7
1hkVy5But4Z0VX5Ef0OugpT0cGHUJLYR+n3WXyBN6sv9wcVV2TEesosKKft/i5Du
Fx4lwL/qZRLtDqHCxPUtEnsLF7fytTYXXw2jYyVUZqB9zlu9tbqqzGAtPd5L3kxw
dlD1NJ8aGfN+o1ryIwFDAG8vEUxqOK6Zb1J4E+FDGYYIQE6UaWp03yZqtK4jwpkc
/U3+OC4Ibe+/QnYj1D5slCUmTnJG6cRSnKkKHz5BLXO4HNhU60R47cP0VBmv3l/i
KrT9ZjSnDHSKFiDeCbFw6tjhZH8D716Dw5jh/3YTdMkKzufZT48mXtJtIIelqKi4
lNKxqkoSf1/96SVJaW0BmpSmsn31bcI7ASFUDSJlr8hVmUwH7O252fAjC2cuVt4r
U48MHVkhGyjh6cco46kQlOFZl0F8zQ8e5S5q8o1mprojR2Yj9xbH2j2hacsXJTtO
TvBL1uV3RtUWg3zakRhV+6V8iyIyUHvf5Dp8QmuE/G7YQoS+NcYSPyngm8l2yXcG
P38H9gvnI6nD47UYGYR7aUM9VISd7pkjogvfxLmrCuhVj2FvN1oRsfA3iPjlw43Z
/cjHs87xQQ+I9K6ZGfGpXD38dzwLyVIyT4G6DPcrW1mL497XULk+u6n7GlYVX74Z
KodNzsZ4FovaXO5JPQHJO/Y6wLzHZpNqwLz64CLJ+yHAeZM5+/YKgyc1PTvypBQZ
Ge7N3mva6j6sohG5rcSSPGAHREp11BA+awCamQKgHxFwMmEz8f4jjz+zkgwbVuP2
I0yomfHYm50K1uZ6N9ihTslfeQll453v8H2R5iUxxxzLDww6QX69bsScMfOY4KBZ
xAbcqMJSqsbLq+Fzy+bqIJ85zVwtdHMSzCtlQscIipdu4kGZb+DRTYNoph2QeRv4
bx9o/Sud46WV/6CkpnY07nGP4zwboTOfZU/emPnaQpECztx067ICTfrFelKlELRx
Y14PaVMWatj01GvTaqRF90JVePz/c9faQIQaMjUb+c3Wr3WkrzmJF+8mvyUo/yVT
UVu4L9t/+LwacuBtbPAVRA/v+0KL/OFmECdiyySjzEA3Uk5UYJrGl1d7YU9nWhWd
K1Md+AxXwj2HReQGuKMRhgyBfzVqb+SumBYRLYvTKzbmNOzHOXOWPYX/4A8AqCsp
1DV1seDi5GO4cmptsk6uRh5g63SsjLSe1LQzYYpg21bLfDmoZONFLTpYdLuy3TnC
1w6iWSfaO5s47zo6TehVe17Xd/Zgzv/oOG9Rsr+KiR/ycjfFY/EDYjK6A8vZfWoP
OW76+MGuZvFiHf4HYdO2Q4LrweQq/bB5tcApHtCWM0Zr+UVLwruMckyd2YNfX9sl
WO72jGhb1RKl0rug69GjHp4gj/3qO+Sp4ReSaVv0KSRAdlhwKh0S4Rsa1XrevIG4
gYi10A+R3b7fkwLnH90LPqwA+0WMm7FHXZYx3FNW+NP1vg0YRC34TH6RAQeuxn6r
eSijpiP4efYOu0ZqUYfIxU6qMpCzYW5rePrhfZsmiAURX93UjJxXBKSeNVN0NQw0
n9EhsryEMcjHsKbhRfmOVxQPEUyFJZxBJp7/224lddikhNjECQc7SvZBtowuH3Kx
IdIZq8KxSOegxN0HF185yHL0sAJVnLkc6okIGv6vhrVaEXPkTFZBTtKiM2VQU3l5
WjHblnwstOKVs2m2RQ92oPQbk8dpZqtgrW6bQCuxCRnjp7qXGi5gpQmTxccWHluu
AC+/cFVbEXuPxtED1m25Frt0Rljs7KoiGJDh72+WUo82Z8/ouQ6/cWS1eV+pin9g
yOfmn810hfuYdzVC2OZ7o1XBnPpssL4/JLDEujnVwkY5skvnpBLkxWIzkb5ff5Yf
xuxeD/qDpkiWcijPkONouv6BCp1ppq44L3p63H4GAU0OmTh6/ZvFX4bmpkowOJ9Y
DJHUdeV5Lmo1tNgmdPYEp4CK78y0OWBk5if1nm/ISfRN6ggcK1I1QqJo8qA0A04P
MQV+94rCFkKeAylCCVJA6Tes7eZy+w9Ywo74/PUOgqWrfM1Kh5P2JiraA7FCCh3l
luHmzlonelAEn2NMRKzqagM7lSoPsogsNvGBEgDEKMPOIyO6bQD/lm+8g+z/YdyB
XhMQAZjIbBJuRYpD8ngDiahmCA06KgRNPqvzI6uXsakPOjLH6V5JD6m0AS0eP/xA
9CI+IcjFnO5IBVyo4cLcZzL9kBylXHzcBEmoX+yR019i522HCULhI3TekjGQAnaB
cX1WQXCEy6WMuBSYRWY+aajZKnAIU5YnWhCLi4BCTgeLiS4RUSuXdtR86HTy88lI
TnwR//5DZ9PMHOj2MBRQ98AiNDPpVy3jM+vW/4oTa4JVypHXq395pUGnt4o4Tvh0
XZRstgA5As3OzuNYmwzJ+MPI97CXrLz5eQrL5RStEf/AaPI2g0E2sjfQxWW89yQK
cWkkw084LMa98up132yyFwcbQT46/+Fagu/imkWkMHPsXI7Wf5qZ5IfKYHzN/RAu
pfZFmylen57nZY5sXhxhMokhws0DO/HKWF2ArD7X321wUAcUhkzPUIdcOF6Jfrfv
PzJDVMVl7Nsv/75jMXVy4dNEIZpr8DLx7yIeAIAEujk4WPdRGReq+MVFmMndS/2K
h4T+1irh4Vl/wQnbukEpcRW5bNauxu+Bm0KBfE5vPWKAomkYvoY3QAZQ9t+TBVGx
71WUJlO2B3azoPpo01S0rCdy2eZnNInaD+JkJe9okBxP+wCm6crk+Ppd6Trf+l4w
32MsjWrMZStQOmxeF4hBsuFR1rH9v90Bfgg+pfV3+Sg+OuoZWyMI/KHlRnExdmss
2WxV3MMJsnlq3Z7/wweHWFXy6lblrEYwvRx3vcOBzgo8mCbKvPAIrBK8ZIvb8SsC
bmEdc2hb8esthaOq4370Gd/CxizjhedoShSO8V/s1TCBNPglBS34yQWmDgaDhzG5
0hr9kEUBuV2qG5xZS0/M2sa6qPpS8phOQR5CwNgRwsXpbKaikzscP338ulZSSral
7dyJ2zMnb5a1C2L4Eoj0vMX/sXJGnnm0OA+0N9+YAFigAyva2RqkMggrFOu0mvdJ
IX8iMmA1k3ltPHUFVMSJe2f4+SRobeYDnhrGfJbVvmfDgmZGriucEXZ5O67sAZAM
YyhgVotHj491ukHLSKixSj1Rmgxm7Z/YN+KypUc/damLAgxIy11yVg6sxaU9DU75
0XSnMRXxPElnyKp9V18xUYKBjk8h26OC2Zgcy880f+LQ1SuiTavIabqKeeJxHg0y
QK3HKZEkJDzjLm8ORyZOfdgXxsR8zEUtkRhvOvY6z4+CXuMs4GX/W4+IhG0XbQWq
Fh9eu9u7EWyyO+CsPwYZzc9YSHpDxrkFdeQFOtOybrugRbzBYSX+/1CpzqXuBRMU
6OLQGyYkPhIOQ/vCzXzBOBCCBFCi9LYl9ZfMOjYFzVgROhT/ce7+c2/U4EEh6WVt
NnCqksC/gKAd2VA6vAv3xyyj2r1D/eaXivo/26sNwd9y6KNrXEh+vVVitG4vfNO6
DetnAfbBmpfFn5yBmsUYjXZFTpsAGTPhhHZ5CEHhDx3nUxmPp7cwof7aMCv2Av0g
jE1MswQW+20SZhOZZ9oDRv9d+ijwunP7sziY9dUvNRle0tEkJ57rSAcwEWLQGprk
uwdPdVTUL/nllGzqT0ePRss54TVpEZLrNhe1COfWryHmkSBnnRlzwTkqH+NHa6Rs
thxYYmmYmdyPgLw7HtqC5WML5MuiRfPKBZPcggN+tVGNleqLAHVFZUhVmL345s3E
ItA8jSH7kQBei/3+pk0U+L4h4vL2D337Ox8Ogc0BQ5+rGSn/BfmY1ghKpE7Q0Lej
LnWkD3MqjRLiCFsvjBSg/g0qSxFud52M3uTAvSjG2pHQWpv2KvdlGJXaIyUDV709
V0E1DuzrMHOXxWILz0xfxGGRjuE3NNIagL6z2iw5dWAuv6/nmGmC6zp91JRXesbB
u0laWlTmXYNqkh7J2Qy/3j82957rYmj4e9gZ47Uu5Vv25Qz0wk3swhFfhp3dsmas
RhZiihv2gIeMGwqHPe6n9/cOXxW660oYqHm1yjYZ6HNmQoHG4gzC0B/55Rne2GPB
akrpvzFSJtdi5DZHTrNTCeyhGkB7Avkq8qW2qALH6qHVFabuRDy8p73P0xjvMKKz
/K7lubu0+i0n7HCzAGxfMGFe+asrH7hKrfFLXkrck1k0kHNS6Vb92kvRSrg2tVLG
PS3V5AipaXhytf4I9JwqVS0F4xKwuhUgqKP6bjO/4sqBxO99ut43JDangT4S2OFm
rLD40923hjFCZnJylJ9N+a0Y6a5gwBgJbV8fU66jiKrZKt+/ELXol1BJlwjen/24
EeHvYlxJGp/B6Q4RWmFpZ2l+m/Je5E4htKS0ppVjsDJ3QmS4xiqkmGaCfOl+TAZZ
Q4Dpqi7Jm7fyChJhU4zzVL60o5FEGQvrgp2arQLV2M017WNbjUisrDKj5I+drrmz
gCWbOf1qe9S1EwvY2pP7dNLHK3iuRM0iT5r9j4ochix8SYiKApl/GmVhpFhWBDWd
dEmwYC97g9M7UWUeBnLW6ymETs/kJLxazJHWk9GRxJMUKST2BCNJJlKdG2OCA46r
opYfB+Pr0RD48AcmK7tG7t5mDlHg6kXWxnRCjoUMcywDX5IIh+L1ChgiJLgOhsRj
tHKltUq+qxAbJ30mBm1QiwJbEQVm6aaqtRG8DiLN3PmAuRh9B5dzdQ3R9iggGPMY
drjqnkLVNGO7D5896LcbtGxjOSqqoMJonAr+gpRJO8W71o+dDSeh+1Is4dZb/xzR
KinQaPd/mLg8oX0QgTPGE1HZomOnGBF3Zo5KKzFT+YlkWrasywpLdmVg9WgqvaW8
HDuNSHnnuHs8jF8viDWL0yK29gOVxhT6ATTQcGK+XlL7P6uDw75sr8tYCzjOlUkr
yvi81MFmiwlZ2ayVp0vAHWxArqwTa/YPZrJNi7TvKlK8R0u32xmnAzcPPINupgGX
4N4lM5+5eRmkYf9IWMs0YmGamO+52uFToiiiV870IA5NY+MScqRtmUT5P3+zekrS
TUWd8uFg8TWCveSj3/SvLXH0mG/VfC/rqYEoshxHONCkd9NnDup6gOx+nbYhAJo1
ZLe9SOa3N6jVUmDhrQNBYLoiJ0CDOiFOBUgZXYS+fKKeszvC3wo2qirSzPyqJjBY
nir5oth5LObiajrWCHEmHVTeAc6IGgQ7fj9CUGyaNn9MphVmkVPTQGfzRKAbxwkk
4tl4Szb0bjR3VfeKbAWjkQYQfT+BkE6nRtYUw3KWGUuGNjo6lEAERT3TWCdqcdkj
3TLBNy1SkMFBEhG6+/Z7xa+QWA3ogW23Nv31AAfHMVYPKpDB9DOxubtOb59HoveH
Qdd+mNZgw8bhfMj3LlUP+P6qGjMoiqegSuAn0UgFZgt37WHMaJtNuuFV1wLDooxX
uNOYliMvEvYAmQ269vZ+HR4v6Gccm6cwX6U0rmCJzKG5KO6Vd12zzNX+pLUD9+2H
EGql7oRf3aXM57Cn2uU8KtgH3/dYQp9j9aYpwUYt1YUtbHF5n9fzNP/5Eh9Sfl2P
hAbmFLgTre1Gxa54wQ447/VgdUEeadqyt22Ya/UDyN4mO65ALW3dO3r27WoeHqr/
aekImxzi4xwartmKGyR/XRsvpZ0LZ8SAk45QJvHx43IFdd+sLlx/PhzLcKtIWMN1
lFFmo1w2C7pO8rKpugnzNJQunz6t+R0AasaLpA2Fq7K+KxSCcmZXdHxMk/GRpE4k
zxukJ6cqr7VPBtahkZjbeIMoLyomkYSL08BO+oxdwho3DWc4F5JBuWvLJxYq2G0C
0Z6nF1o1KuUTed8d7jdI6RaS4QeKmJNj597+gBDStEB51kIhFfMN8o+JpmdS4mBB
NnM2zy+UPZAR3BfiCkpCBvrEYDRqScA0QWsN+gpEJNy1UJ4lXmafp6ClADHax0AN
mA2VENJqwuFYj1mJTNfRAMHwteLnqVf9RTghTxM1dDErjKCrGrvf50yg/xb2U6iM
S1xAgfDjNO7teX1GvBOIdE72flebtAtUeUPXlZXsMVeAj0eeLa29MpCkyvGYzaV2
GetLGkQ4EaFq1rLYG/jw6n2azbB2WgBcJI6jps3y3NJv+78w/FeA7jDgyL1NZSAP
OjmZSVQ61RSmDkUZrXsYyN28/9wEOPzUEtlA/gc467Bg/D5wDrgT/Pyin/DVkZct
EVjFUTGQIS55v22+BYOueYNu0GqVu3Jpks+yVi5ffirs/eJPi1FEBU0rJYqEqMmj
7poYr2ZWfuRp3U2aSiy4G+fTHRNf1aaRrf4NW11xBuV+EBcIcDgVqJvWw7XWx9qE
MlxqB2Wid/kgWI6tiPAH68a8ZjuApY9i2t4/yixNcltZ5Q4/5vY6ixMSY3+OLLHG
lSvmZ51vksiKPaJo/G29JzQcuMws6dcgdYw69UCWnps8ajLGN8+u3RkgkpSJ0IGA
TBorFIMUmj01cM59P2N+3MlSz956JjegzsckN2YAXNmP1Kqe919Md7VNQLXQ/ehI
wKKiLic6hU9Ca7lZuq4V6xQgmtC4F81bm0Bx71oVaS4gaD1DJmReGXKMjbjnHthw
z1Mz7aoNPCTcI6Fwn7NGxIqj05VkTkiuVf5UEzUvU2SeU+1Jh8FQ+4T51EuA/bSB
EOUjERxdH6KoLCLgphuFJM4KkERi16/hyXVop7D8g37tIBtr4Bd32taWfX9+/5/X
G8yoG0Bwsq18KN8idLgrZGMymeubAvmPggSLo8ktcaOvGTGQYdWqz7YFzUplmPIk
wWv0yEkuG8x04+jk+/X7Wh2R8lcuAIhOZPEij7+moe2Y6KgLYx2Gv3a36xvCgSqX
8K0/jJDKYPQWyPybYBEFyqvEXLQhqNyloSDZtcmAJt3WcMi1aU1NHFw/D3FW//DD
sDbwlIqtnqwd3XvXhi+0Da8JJ6JJJ+MW4WiNra8keUai8MBaAoyyvjsj9H1MrsMg
PeapTWYUvacVFKKkueNwGXKKUe2uihkX/zWYMlI1t9UI32VPYIoOFe0e15fulmjA
xwlur1pcU2jQthSTiW9VnjWSB9DkyRKpFHR5DBM7NoMngXhiQjJcHcxDKW7ffdAG
62UyywsfpP8O4eJGXb1Fe7esGa6Q/TTi8aWjH9joWEmUq2nNTszXYzkpzctH5/ep
0jKw6K3PLNdOLQuEq6NMOMHBe+1zTG/m2yZT1wcr86xuVMBep1e3C9eGLcaw4vAt
5gYyI1dbuPaMPG+b7f9GHbFMhw9DW4N7sBMaWDgy5ZNx8CIiZjVkI3Q8kLAtQ7ja
wMay76qHonhrgI9h/HeMky9fm9iGQkbx6NbhreFUNf9IBI/+Dvjnc57W+Hf8YN9N
Up2M/8NdtQyKY2vnr2TH5sNpFrUk+38h7yduXp6sibwfe+qtEqJtSgdpl3I1yVek
NkRHMObZ2gqfForyWmvMz/AVmDAW3vwk0q2M0OnDimH560w8dF+hMqD8x5zlPSnC
oOwzr1J0I0bPrMSa+UNrpfXvWW13VOoSxjo9emUX5+BaExTglkR7sK+O3W5r7lWU
i/pMjd/JurjPLFBjHj3JgG7DQ5pPLOYoy9D04lpNLxHE9iwDByBx6HuUwNpIB0GZ
xKeJrd+Z4aoxrEFibeO/8pGNr90XbR89HlYKAcHa96IttfFKaVqNwoHPzrAFl+QV
wzh/I1ZPUgkewc4vA928oOYGbPJmNdByvA9BwlJkjEwaoSO2HiPngozo1QL1vmMt
H8CiNvLOn7NEFgL45ZrfxB7inwOoDS4dcD+KLESBYi0VLSvxXiTIu1M0p/jby9zl
86UKsr8z8Re9Tqo2mkepNUpFL6dXD+VJyT6uOzZ2b5BPfE/W8kBMu8VWEfOf0eeD
CZj7Hx46cTz5HD5c6XX9jCO/iA5Ijr0xJGPK41IMQV3D0No7kytq2xiQZx1jpJvK
34JGepxjfuQiLXlT1Hp8BA4aFIabVEPnwVs7JRtlhnc70ard8hITLvYoa9gpEVJi
6T9lqbiQ3aYYdceD9jmUr4OrH2EdNW8WeexM6C9O5bW3Pv04d81m5yrxPSJeerSL
6/WhtjHm7V/zUqFzCTJkmOQJ5SQG5MgTEH1CvpZVbwFEZ16yOlfDfTnFs9iHN5UJ
/AQTnODVKEa6SZafvc6lZZY7MC1EZE7n/uOfpKpY+HMFZvqBPf3ZjIKhK1sCLDme
Fb3VLRD4JJB8DLoODZd4hbBsekVvhmBVeVV0KuOA+zf6u95P+mdpbMFVMe+2g7FM
QL7XVLAvPgnsLiNT1n6C+DImYJFRI7bTLvw4ZXas1AdFxUKgqDYw0CdbjuvOOSAE
pjmzBnQjRcSjMh5tpourMurlWdkDq17Mr6aQ4J9QT76ME4rcdChWc65fc6OV/tPt
rNyQPX6nmW1RR0Kj8F0ZFtthot9J85njCWDMcO8kR9NTB0dYh3acOHKb08oeM4aM
xzS5jl9ZYmMEXBEunp6QCs2Bo2qPyCcoNXNYCKSdfnpRyVd38b+ZzILZnvrA8RlG
m9KA22MjPdRFZBcjpnfdDnFUerbrpKRyCkoOTyQNeoGrlr0pambhkRRHPtYnA3Om
qM/SSo0jyMeMi97zkbJkEFKiE1CtoooX0cLN+iM6phCZfR4bhqrEb2ZLxuaqRrm5
i2xVFmwM+bXeBlE3nrm478bYGj4GJ27HrfdqqtucEc3nqw2DKVDUe8LxSCMqgBQB
9zzYOgrlwSg4mKsCdCRt0DXZSSKZplzRvgB/jOq45o7AdbHYnkz6kcgUookg20wG
k4UlDETQUN47BJpF+9pm4T7FIGAeN2H++LS62+A3Jxcm4NAeT5quhsc0GesWbLQ3
9SJi6gZJcVpw6AefO6TlwokFG1qyT9QYZWM7iXjVP2AMKHejO6OL3cX0bVnu8c1L
Lnq+m8/rJ7edtZTOmwybOEQZBYzo25MdAAy7NFu175sNm//MNXcPOXcj5Ap6xrtO
TV0lti9LiVP4jNXCW+Z381ifbmY/aZeQtci8nzMee3jDbd0qd2WoMrZXeoVxIbTs
/1N4DkdSuXVk+ndNeBIdpBjiuY1MGka58/RNlE/Y7lAivq2fP1tUxsl2jiyt1wfo
inAauCVk7dBcIWf1ghaVHZXKBrgSbk3MW7DOqjnVyUNY9GXCtLj8QPM+Bz0icvl6
3lXmnR5U3iUfawf6yLVFYJDjcIi0aW8pE3mcePOqmZBIDRqaXZR0Cm6w+0x9tcLW
Glfd5HxAbsGa22QWM8wbSEtYqyIr7co3xm4nrWs6XNg3mFH9Yz1TXwJP4r6m/iFg
sfuHQQEndmC9B/mIqeXCgcibKdN1349P6E41oPP8W6r+LphXJIfoRnOPa1Tqq1ud
WDkrH4uq4ghRKJ45GZxz8w0wry9nY28fpMY0kZH7H7+aY9KkHp+OP0jfNFOQyf1m
mLPTOUADqzImK0YzSgsLNbGKFGmHY1slYKzjQxYlxAOGcu/11KmR3gHEvGGr0cDm
JChUfqxPeO40+65LQ0pWByruFY4mwXMXYJoVeTIdAJB+pf2edqPX+4FQMnfrFRnI
syCfoPsBhyOEbTcNyBa4EdeyNtMQkUCKnywDCDQ/F1kMR3HWNBVTwFNCiBsQNbfw
PtBaqO/y5836m8P6A2NY+7apIkqCO0F7WVD0GAB2hfz0ixkX2WLCsTZ6zf0qKNWD
fwYxWohglGP98OCw/NFUvGp+k9dEUpucq7pXXZOuw/chK3/8GFdQPg9KSiFiI/W6
hTTLnw9zkWm4ZX4pf6NR1fii6lcDy6nbfilfjXURWQRsl2ZZF4ojE9uVQXQUXbNd
zy+zhZ1GnOXsTgjiKAtxenoL/VX2b9NOCaykJWQOwspIN7mL0/2fV1lVdUainjN9
MKqjrsxcVQHjYqbzQYtrdK6THFcM3XVg3hWyML3UgRWyFRSouC4xEZbkeQlgctQw
ibUmqzqnWjuE87wUuq3KZ5KHYs044Z95/JCKIVlBnTzCutHVKO76Fp2Bg6NEsSxv
WikLEEt/qwprh1JhGpzEpFfBHKxeHQFbSy59noiWU9HJ1QjOKuZ3wXxdaZKabTaH
y4SNxIBHH8tMOmjEfpr7K6dav3vOpf+W4ZkxAbz+pxdKaZtMHLTwWdLncmBGclJZ
IOC5t3tGDlpfaLQgjLe8NyV3aP55z3d9NmhYClfvhOY=
`pragma protect end_protected
