��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�q�E��	YjpA������2o&����ޛ@��	�&��O!�Q�p����B�]*#����Q�9��]�I�Ȧ���S���볲X���q�𧺯9G$�$��5��#ě�Av�<lŬ76s�_
�*���p/=�S$�;�1�$ƺ1l�`�d��c8��h���J���r�P��<X3�O�6�C��i��֦C���wш�yj�3ϻ��UJp�t� !qٯ��p���&��O�n�:����MO�x��}ٴ�曆K�0���T����L&����f���%��l1��G:��)�[�i_��p�Wc���W�쪉��������c"n9�9�.D��� �	�#��N���]��ӬZo[�`�np�� ��@5�� �S��`�k"�FdIoa7s�>.��5S��)�"�P�A��:�������V�MY{���X��]a7<���f���N�J����ꌽ�A�ܳ����j��y����Y�ܦ�5�� ����	��[V�:� Y�Jm�L�Aq�1��e���T�^>d�����ꈼX�u�^�Ӵ:^q�0�� �/DG�8|;ᤸgV����G�mM�����A}�|漑
3��xY5\�B���I&x�]�ϭ�	�_�jM����ȵ�BW���nl�d<��g�L��<v:�>�Jg�L;�B�>0}m$v�C0W�	3���i�Vx�L1,�ln�O�+w"K��~\���h�dt�K?U}ݎ�]5
mԇUǯ�V�%�u�h�����I�"��LE����(��Dz�[_�+sW��uU[�f�*a؁�W3�d�����,��h/�0j��K�"�p�@j��h�%&�za��yv�h�P
j @���.1�j?;��W�d�hf�YPl�F��vF~�b�_&�23Y*>�0��Pj���O�0h��\���g��M3}^��(�LȀ��p��b��Ơ!���W��P�������} ɵqUG`0ˋ/�!yS>$�5���'m��>A�\�L�2dߜ�pb�5g�±`��S=���r�B������L������D���IA.6�u&����E�\��_`O�h�9��c������p_��"?����P�It�q+:1��j��_�ã���x���WYh�.�=M��,Cnh9R�'�ml/\����?�Uo�%�]�|�H��{�N�R���t���&�Q�j7�]B�dq�W�Y�T�w����XDۛ%ŲK'!q_(q���J�!$�zC��˸e�����1	x�2n�T���2�t��Ѷ��0O3,�2Ӂ�}�r��+w��3���ԝ�ۂ@j7�V�b5���ݯ �F���B�P��������;�����|�U�����~Ok>�Ԃ!��W�7����~,/��)�Bp ��7��g�N��v�(mT�K���֣F���M�o$�44*?��sLI�w�~į��Ŝ�$�Bh�#�
��0��s�B)0>?�._�7~�B�7�V�y أ���O�,#dǒ���Y�����g]W
�:��6C[M�̎Q�~����z��S�Q��ܝ�H���m���u?��I�V6�>5�O��z��U�MX~_��!����&~�h }_t�u>в�c&�[���&�c�b$ŕ{���2�Z�Z2]���nI״z��R$J����F��p/<a$��qǠ ����sر�l�1�0)i��+^h��$�P��3۾L!��G
��Q������evG���v!;W<77��D�-h��ɖ��m��=c�}��Q[�}�������vf�,��P�d+�~�m��Fl�2��aXZ*�
�<�� 3k�$5��	�[�w+
�:Lf�"�,�ԇ�d�ve�%�H�.��V�"�t>=p������6�\k�酻�RK�χydO��'Rd��>��|v����I�g��U� �5�8)f����y��׼��]H�`g9G�<&W��G�>v9[���Ͼb	�:Sq��YfTy��Hg/�ne����i�� �)ZP.1���=F}70}��mHl�y�p饧�w�'0���I���/Ԣ��$dQ�(x�u|�	�1�^���k�j�S���e��+�#�F�D��lg�i�S����}��..34j���0�����E"p����ʹ�/q�q`!�9�qZ����<1��aĬ��z P�`�2�d�������$�K�0�\�>Yè:7+� �&�o�]cι��Wm�^Y}�kh�ֈ���[��i��Җ:,�tٻX ]�th',�'B��i����#J�mtǣ�S��Z����߂`j 4�w��7��ʱ�Q�S�# �w���$-]��=APD���3N�|���u��&��#��ի��l�k����
�Y����Lh�n��%������I�ʺf�Eg��w>"�O����YS��g����p(����fH�6���`C�P��t{�l>ɽ��kb�8�i�Y2tl  ����ݭ�}bc�W�΍{�>�5./�T$���S7a��d����`�Ұ�:$	��l�]wdp]�j��B�<�)�|I9(�(u�5Νj�C>�{Ś}��p�?��:�u��Gk�(D��"L�0�!
����c_\skn:��wX��;��\*"[�^�����;鉊 �w��h��t3�Ⱦ�~� �.Wo�P2;لtWw�;�-�zm��x\�������L���:����BTs[�'�j0N�k���.&��[�X�o�h���C@�ÿf��X�/�G0��=�o$7�\�c*������S2�'4����̄�E�AA'�@��j2ؓr��������Yp�$v"t(n��]����]������|�����Z o�K�Gq�O��!�ATԬ�3��Bz[,1Խ����ssyi�0Y;԰S5b�p�Y�[*�o�s��#T�Yf	P�y�Y�F�x=��[���d �Ǹ
G��e�����ߊA QE�� U�9��C�D]������IP$��F�j��8�a����]+��"Z�	��6���Q���p8{���Q0V���@��a\!iJ/����O	�m�Q��'F�S�N���������4%F��/q�0�a6Rh�Qdۛ6��~���#�����$�<g�7OKW���s�ĴpETy����۱�e�]�̂w.C*�Bް�r�~K�o�W�t0�IAN�1�����=>��W�;ɁM�p���b��kXhpE?�;p�:C%��-����~�^�C��&$��hQrEH���!s.��S�4u��h����z@8��
p�� XS^��tw	I�*���A'Ҿ[�A�pa��U�Hv8r�j���a��_DGf���'nv�SJJ����;�*��\K��wWp�Ԉ����R+�ū��=X�YC2��mu>U����%��D���
��amLс��,�x��>Z��"��;n�ޒ}�ܴ	���q4�u%JП�K�xϞX���'�eb�C`�]ȭ��9�����0ҝ%Q!��ybXŘ����k���cN�P��⇨�M��7w�Lj�����R0Ԡ�1��7d���[#�$!��w�x*$|zaD7��5;>��yC���B�&}�o_�7�u,��T��6�O�(?�9��p#t�q�<\�E_���Cog��#�e�}G�>ƕyc=�K�#6aH�o�)���̔��{z�}���Ѩ�m8eG(��4t�T5:s} �D#�<�:磄���V�H����Z*�:}���r��Q��N#��Ąe؛!'4��=D�)[��Q�Nj ���+b�5[��e�Mq��ز�݋+QY�3���b�`�\֛i��/�C�BP�����#�z"q���h�����]�E��q�Sh���j��O=�O�0�0~C�k8��Xr�6`����<�(C&V�k =�+t�O��H8�?�.���t���o��܈we��AnP���;��y&C�󚚪X�(۬�C�]S*g�'A��s��	�Q>��wϕ4�;6)��S��l�.�-���4-����S���4�
7{~nL��뒲��:�6���#ރ2��E���=������?ۓ�!c��2Im�� �g�}D!��p�ׁ}�i�N�m��Ͱ���*�����j���.?.qO�3��V��K��L�9�1^ϗZ>g�|�ł}�F�wJ�>��֙���� ���Y�{q�R�����J�+jwƧ͜n#
��j����i+��ņ��L"��>{��Ju��6��-*Jh����t2�Cy֫�*��AK�r
�C\�ܳE��5j�_
�HOu�u07k��LF��T2�e�%0UTs k�M'����пSZ�'�Y�r�I���0�C���6����		EJ����&)q�k�Vu�m�.G�U܁);�����5 Q��v?�P�V7 :R� { 9]�.��{U�:��V��	4�]m�|3]B�Z.>G�F��(?��=e������.�P�����Jf�-!C�]܆��Do��3�c/}���gK��%�@�n��f�RI�<N_drj��xS�������Q���W���_7�� �߶���)�.�fv�%�{�}�"�8#[�1��\�R�\#?�!}�9��yj�~f���9�c��[bI�`p�e��a�j���#�9�\������l �����L'6ѷ�[�CI���!�~�7�4�jm��h���aL�o����e�]2���GR�_TK/��>K/}i�Z����$e�h�J�0da6F����CL,��>P4��q� Kx '��X�/v߉E��3�ZE���&CFՐ2�b��`qS�����c�����Br��T�A��a�kB$�l���֖��t�Bs~Ues�ܪ�4��5yw���R�Cr�v[��'>s\U߆ �k�/�Z�}"�	Sy��H���j̟�A��UnB<��d�D&b���0�M�������)>�q� �Ty2U"�)HtK˘�Σ`�����K!�emͣ��V^��k�q�0Y\�}���q�9���� ��L|�6�"S�>��`C,z<��O�dU|��vg�L�k��x�e��;�����t���p}��{qW(׍+�HΦ_�q��æ�J	��Ph�=,���*+ �
�\�ꇾ\���M�Jy*a�}.�w��l�����T�0~ׇ�oyP~�|��˳s���||Cpp޷"�i$1K!1��`����|���H��q�$ �M��"�'�邯Pw�f4`�i�*Љ�Go��OAB�]�*��R�lk~Yd����ܡ��0y̦���ID�Ћ���3+y� �10A���Kp�:��ǭM�Æ���+�=���,>���Z'E�]�������%�xT�Q����Pa��jͥ�A�;�jzN�G��8|`���GO�Z�"/�(u^�:x:s��ͅR_����e�{-�>?�4d�À���!'�q�d2B�z�[f�|��z�ְ�n�_L�c�j�"{��,�,UU�yVks�k������kң7�@�sT�s*���?2���U��4�	 4�笽��[>ߐ��FIM
�_�f#X�{�A�kX;�@-RX��������R{)Z�0�iS7@����)>XP�����������hm����X�uP��"ڴegR�6>'�@�iZ�:p|�D�3ǡp�Ak~z�V��Ev��~7I�{BH�K�_�E]������W9);�'v���;��n�c�s�Om�e��G��`��mS���~�8��w�b�.=Bی���ڒ-{���-�߫t��^�ʅ�LK�����ad4�l�4-: {��p<+pT��(�4X
v��#�������n�-�6�Y�Y|�c�?E&?eAv�0������{���b^q���D�>D%r|<��BC ~��Og���-x%�mQ<UN���'�#�&��~��8u��W~Ծ$�ᶟ��ONZ������J.m��~�ʺy�cd[N���I]��p��	��[H�wtE��8�8�遘+��0�˜��$.��U��x���q��ו����=��u4��	���r ������1%��������7A�	�A9
'Po�`"�";t��4�Kn��4��CU��Bh���B�K�ӟh�C��:�xw���[�Ŋ���]L�<���׆�������}�9>Z�ݮ�c��/z��g2��_BS����"�!��%�c���+�]��陿EŔ���ä8e<d�v���}]q��H�P0�M8�2ђwy�N��>.-�>�g�$���Z<���`z|�~/���ՑvG=T~F)W��C�?��-���ϛ��\��p�*1���B���Ϭ��P�Id�rx"IҾ'�'�$�b�N���z�iaV��U\%<i=x�Φ��ߊY�s��s���.�eTG�R�A֛4bL���{�Hڲ�
�)u�+gU��J�{ZV9��ѹ�]��TˎK���\��J�b��!�RG���0�o�l��%C@�{s��G>��I/��F�O[��)K�:7]DX�Э,����I�k��g�$i�5wi:�o��b�n?V��.3r����Y����)h�hܱm����[W�8��V�ͨ��T�ܥ�6����=D�w+~� P�ڔ�A��;���=x�93[�+�7�H�7�����)�էf�w�0��|��q�`�𣽿�N�eܛ��f-��4o���v`d[�s����^��10����<����_�p#)���n�QeR����qR��r`��ԅp,R�]�"�䠌TX�SM�M)Z��$��% '�[�1��_t2 7#po{���t�uͲPL=�鉶-�PA�����[͢�ù�q]-��:��*Ϫan@~�ZOf����� +o����*K�����~�l�r��F�y�A^�{�M�)L����zo��"�pkH2�TYҫOñ�e�J�3m�H��uH�T��M��G�H�m�X*���%v�^	NUA@���n�(���k�1�4�]0�@��s<BI@��ơ���^�H=ٔ仆d/����9��bz���D�,"%�:A�yŲ��d��in�-B��w6Xm�W�8t;�H����g�kMr��w��jI����mj�7�h�a;�b_��<��Ji��I�HTy�	�4Y�F$�X��'
x�[$�Ύ~����֛�iB�.�`a'폋1���.�b��a�������2Կ_�G��9V=G�X�����m:�B?�JF�z�K0��������A�X[��	/G��~-hru{����w����)!Eu��Q��7@�&z�k�=gV(�ͷ�A�|��5<1�e����?%���$���<vK��:�06'x�h�4~䉬7�3�E\�G^R#�
� l�S��b�~��@?�)��׬YW��YSN���[��=ᣖH<����T%��Q�8�R�q#h��r6z��q�rM�U}�����8�m.�a	-#q}���&�_Rt�Q�G�Fr ����1D�����$4��O��QS��<;��w�r�c�`�N�������9`5��\䘲+�P��둎�Xަ�y45���Ū��l��I�������8C~����I�Qy��^���9K��9�l�̶�+�l�H��O�
n���o���ݖℒ&G��1 �/�w��Y��C���U�P��������^����m&쯶�J_J�3��b��'��y��<����=Z�{ F��4�*ѫ�rȝ|(.͖`���]!U��NuYi�%���7�ox��Xí/J��[�U���ˑ�����UE;�xm8�ܣ 3��=,�I��H Dz��%0Q��%LPt��S!,L�v�6�9.Ͻ�t����3�y�ZؙV���&��Wl��ؽ�u��hK_5>4��,մ0)-�-8�n��D��"=�<���#��A�E,���@���}���մ�6�W��"g�x��E���#P�e3�%l.��z�vUHK�}���KeQ[�+̄R}�6��V���bk:�.�y+\P�"[kZ	�}��V�s	ws�~���>as����~���I��H��?֠1,�㒦V����X�[�]�X�׽�Ee���	�]�� ��:�\d|�Ս�P.��d,���M�=Լ� /c�����&�
�����߸���]ƥ��o�ܭj9� ��gS6�4���WD��l��#Zer��X�PR�>ñ��K����M8���u�ѩ!����f�]s��]�����L��I=�� g4��L���`۫�vĠ�Lm�-� k��QF�%Wh�qX�8�_�F���!���=�JSO$��]לa�|ۆ��h��`�Kʋ��p���)(V�
��c��F̡���W�Ȼ�� 1�4^� Z��j�
T-6��(�������5�>�$wWx��I|�h�=<O&��Ug��p-U���.��O�cnUtQ:�ؠ�-)���AW���� h�k��g1�����
��*�)���^.�H1��|�W̻�cJۇ�vz������O;ݻЦ-��+}�	�x���ޑm!�^(4-�5""I���I���s�Zo��`%=f�A˄P&:�����S� �i����b�pcP��+�����Sxj=F�	x��BM���^E�����HVHĦ���˲$��7�:�sW�Q����3�M���<�}�"��F�?*=|�<>:p�&��^"|��
�y�"�,��}y���Z���8JOI�xC��g�۴�u�Ĭ�c6���E�� ��9��p9���c��*I#&U+��I����+��R���g�ⶎ&,��H��TAߺ�"y��B���W'���5���;�������	���j�^ܠ�:��2�}���s�Z95�O��u�@;��O��f-Z�R��'ӎ#���7�޶�-�!N�΢���r��LN�u�n�P<{R$h���<P�0�Ďd�|��7D�顣툶S��V)��ŧ�B(k��H���P1f�L�2�O1�
��������P����<}�+�I�;���]��f������}!nE�,�V��2/$v�ݜ�����%�G�����Z^^O�V���"���S��:��h̾_��$�IۼA�A��*�qu7��ղu-f��e(�Nt7�o�7_^�X�a���/��i΂4�韅�>�O2�������V1��T�e�ɠ���=�߰�4��b}�z��11sž��9��h�3����~��eŞ�+o��0k +j����ن���w1N��`o�촫�� ����o�[W|8���%9B }��e�R�^}a���y�[ڽ��]X��;����r�~5����ή92�9��L���Z�2V�.��Ҁn����bIں�a37n|���)f�p�̫��E�S3������D�=���>���ƣJ�܃��L�i-�� ��q��Y�?Zʲ.� .��ɴ���?�@� +�\�8��bQ��ܛ�l���j=��.�t��?p����ue����q�q?��lh���\'IK�j� �f�.��S�M;�$�8�	cɼ��ȵ�ya_�OB	»��u������S���z%L��>��ͣ}]�`H�N�je8ʔ��:8৺AH��� NH��e�8&��<�uq��R��&�~DzI:B?pRf���)}"]�Sk�,⥧Z��&����M�;B��(B+3�/����,Go��mFV��&u�Sj���V�aaB������ҔePO]@c�]dhz��F'�����n����x[�|қ8����y	�y��h��V}_Y2��Y涁��Fʃ��A+Qϳr�Z��:�]6v�s:"V�M3���9`�Ƈ���%�p/�e$tP��{�Y!���A�G��N���*��e�7<��V�d_���=Ll�ީq;tv���$�.@�+Ϥm
�D��MKF �q�X���������U��I�ǈ�V�� L����;p����aW�0u���"rt= ;+W�a��f[-�U�c��T�w�+�"��q�/	�e�PŇ���j��zs:H[,��@���T԰��v�X��
-M��.�Lo�a����#yy���1����ȕ0
P4�ފ����s�
�A$�[����q��˿����Z� ��4�o�J֏ǽ |��f��LҐ������4T�Q�u~�1X�$��e��Dz)�'�<�b}88&�&ǳR�ȌF�e�n��LB�%VW&��0i�_2�:H�&���=��d�s�26� kc��a��������s`tZِ�q��3O�l����~���p��A��`#ZJNޕCE��W.��1萢��އ������4��Y%�>��_�v��4'���U���*��6����[a�p2"\��>t�/����렡��󳡽�'���Ќ�P���r�޹�5�.�F����n����i�:-��?^c�du�Ն�@'c��u%Ʊ�שZ�cӊ���#���6T�@��<:`]��$4�O�(� }�&�J��G0>�m�S�]}=k+�0s�}�'�p�UeiJ��r���j��<Eϴ�����g�������0��b��͢��K�>P�}f�Z�9��y)�?�v"AB$mt{�r��d�0��3pI4+pt�r�d8H�����+��aigŒJK%K�J��g�aG;M��K"��v1?��}��H�sy��նHD�� ���nTA��:ܓT��z���� E\��U�q� �/~L���M���
����٧�@�����o�l��.�6�L��2,��������-��jz�a]��
"������?�iz{[E��O#@�d�4|� �a��5�}�b�A˔ѯ �")M�4��D2XQ.Z�61�pvܢ�@c��~�*�5��rL^p�Ǻq��# ƿv7�%�i+Cc�+x�Z�B�B���L�Q������ZH�T�h
bL��^f����[�9:��{�q�y�$Z���U��~8�Ԑ;�[9���Ҏ X~�Іd8�� D���lp��s�=t�f�1^Q }߄��N�>�s��,|�<�k p�B���&�P�5k���uپ<M������	��г�� ���v�[�@�\5�v��	�ξd���5c^2�%�^Še�L�7v0�q��Q�~�,Fv�Y�8�(�_��m�Pﱮf�x1�o��b Vg�~-q���ť���p�ء��#"/��ap_}�$~FΟb�o�qO�Np����)�x���d�\]������}η!�wj�)8���<Ώ�(�ۀ[�do�A�7�`ɣ�b�X^���A-:X�C4�ܯ�hW��[G<(�Eޜ/F"��#��љ��?sfsg�O˚^:{�=���/2��7=�u������1�ߥO{_ui�C��h���iu�= ��8��$� K�hb�b�Q��>�a����W�6�)@�dMW�[�#K���: ��魜���	��bq�造N����B �-�j�����K0���� ��|y �OZ1`�E�"�t;��\� ��;GU?2�5,���6�v�0������` ����6��F���#j��U��,H���Kk�� �1)="p)��`O�P�A))��"����5[vJ�� ���������<�5�:��훀�~���Q�z,k�,Fx� C�3�o���d�mI Aw>�7\H�[
k��f)Sq7I��,&����6(��S�c�8�3�B�ܝ�E�E3.���`��mά��7�xK_�m�+����}���]n=\��n�sJ|0T�&f;�e=��>C��̖�(Ɖ$�'�۝4�%�IO�� eC�}��柦K�Zi�i_�sYYWZܬ7QN��5C�<��O��ى�L`a�����?ܑ��D��_!�5��7����&�~-�w�<ܟK�%����倚hir�z-h����g	�Z�3�4F�܇�~p��w҈p3
#\O������Nm�&HF� ~HÖR��q$sp�o��BD$��@��S=���h��cwH��//��9��[�|_���e����=<Q��Nu���q�?����}�]�t�I�G�5��E6M]j�{���0B���%b~��|���JUt�z،
"i3<�Sk$�ݏ��DSg���UT��2Z�]���9i�v�#��V���_Ff��U�����s�#C�j#���mx�<ڀ�7�(�)��o�ĭO*ri.����Ttv��W���07�~ye΅ �f�`�٪������
��Q�:�dv�F4�i�%�0{A6�Z,���iV������m�����c��.��d���0�&��>(��}���6$�͂� G�����)��h����Mo$Kɬ1n��
��4�29�[�� h,5�/T��Do2�?0�슃J��=Pv��b9��?���k;T
'�c���ɠ��E���L~%�r^lk��#vC���H9+%1���y,<��`�E��><���Z)B���II��U����L���;$���3T�j�|f�3�og\�!�kdD
�\���I��.ғ��%�o���e�*(rZ��[;t| ڴ�cuLy��:8��P��L~L��V?>�iE�����g.��AI�K����e]��r�|R8��ma�y�~�W��������`�dX��t���UeI��\^���xF?HWٓ�A��Kr-cK�w���FΦئ���hea�n>-���lC04u���%�	r�{�sXۓp�H��d�tѴg�uetX����(ml�^�mbPW�����(�f��)��?Uem߻(}���M�Z���L�S���a4���<��</�A�������E��8�Y~Pַf�?�"�#4�p1=|*Y_��鄱���_q6������d��w�)_�I���Ar_;Ķ6�^��$1:0�KjX W3-�I�}��wB{>a���DNk�C4>�'"v�H��`:_X��F����g%�rYИ���Pjf&�I�4�������0Њ��b0�2�=��EK��,8 ����:#�+;���r�e=�_[��j+j,��������0���0���1���ѹw)�VQ��{��D����/V���e��Q,�-���ЋG���ʎ�.�8����m�i��������l���s0n��R5����{��H�`dE������@tr?1n�>�M7��,Vu�m�L:MB��9ف��mM;;Q1�7I�C�?#���@.�%�$��?�q� S��R�1B�5؏>��K�-�;t)��t\j(p�iz�,޸���p*(l�0��5��!Qa{x��8Պ/G��d��	֦*h�tw]�@H��;�8��X��o�U��$m�Xu�eP-���N�X(F ����FV�@�]
C�t`b|@IY�uQ�Z%�,zsS��A,~���}�%�B��r�4��\�2�+'U*7��y�:s��cW�7i���i�СK�|}�T����S��}R�q~Nb|LT2XFג9��RE����{|�Thۯ�#о͌����B���$�5'E���x�ufz�򳺝Ά�}��H��Qc�2�[�t6|Pz���`f�M�-H�����{�x�?�۳l�{��=N�xU��YՈ����'�2�+��V}�Cs[Y���{t_S�I$�I0յ��hZH�� |K�`]�������ԩ�~̢��8lCu������kڍ�^�tΟ+���R��NDN�7��ƹ{�)kƫ" �V6�sܻ�ٝ�Xֆ6�����MF�k�fH�_7�X,�y)+��`�&��t�TZ���3�R����Yg���6������*fn�K#�FZP�F;O �x�[�6�'��+�0'`���������g}�	�gsOM�TɏQ�Id8fv�ܣg�7X�� �O����f�x�����o2����%�>#��C͒08IK��'N�=w��k�5�+��&��<�.0}<LMr�1�QZқ,����j��A����2�#g3��gِ����eҜ�i�z��_����M���hx:ڋ1[�G�
+^�|{)���4y�:�0;;̼v���W�aK8��������Ӧ"Y��jC�EM2���@��!f���^ߺ��ʾPl�d,����5�9=�hJ���ր	 toIn�	�\#�}�ԟD��B0�؁��Jhn/�4H�|�W	u)��J��3�Bڐ�nM@Ak���6CҌ� (H~[:Jō��0]�w�Aҽ]EWq=EG�x����۸g�>2��M6��N�'��!��w+R������)�)��0����m��fA�|�"r7`�5�&�N���r�hbH�c��H�O���O�u(�<"Y����*�L���j+dq��d�Y�=�[�s�$i�k�����|��᥇<�����0��)2D7)]�I}�W�U����#�0�t�)������t^HG��^g�s��GJ;�l.1������!��r���3�r��mvy�����n.WNa�%��#I���1#y�s�{�# ����٘Q��V��-Ooé}r9b�T��f|s~)��gĴ����
��}r{��� ��5r���iȥ�z,�U3h�.Kc�Žss��/ojF.������m\�Rm`������}�QY4�Q���I��`V!q��'��w��!{�jf�./�����M�����KH[vTO}��Mv��6�
oSzt]ׄO�~p�����J��_�ZH�a���7X�U��u��@;���="�l������PΤ�<�?�t}��Iw�5�!
�RJ����;�w�d�l��N8&���'��>(S�(����⯩����9܈� ��_�T:>9	�6��%L�{:X6�N�ɏ��AL�s��]���`��1n�R&a��Cr�U}�DK&�w-kz�Y�5D����{�.��Ȑlt�JpB7�p$(2��ud��a�k�>>�����B{J��έ��."�'JDu�ͦЫ@� Hs� ���*8oDb�J�6�{~ϱ_�ÈSnJ+�ԃ���*K*G�i%f��d�����$�s��::ղ��JOr�����Rϣ���"�@A?��+�>�����g�J.FIW�XU��ݽb�D�n�Y����1mP��}E�/�E@���Ѐ7�'X������VY��n4
���u�{�֮'ҙ�G������k��>�ȓ�9����	���� v#������WFKn�%�4�b�3�Wk#Q�6,H�3��HSD\0枀���E1<b�M*�^&�Br�⍝kӌ8�D1�v2?��H�n�z��r��
W��H}N����_�EԜK��Y��Hk��=�9�&)9q�`�)��m-d�i��N5��ّ�L�
�P� � �Ծd��ǣ����5��;!f�i�@����g)�b�Y��&�D�)|�
Ռh���f���ߞw���,�ܬ��`8K�!�"L<�=��+�
��_{����؄2�A-��n�4`*X��b�w�tQ�
O1O36��&*�X��!1\ry����rg�;??
U0�tcX�d\�n<U��i��P�p�����,E�fZG>3[qz���G�زW��@�U$��N��I[��%�t�gV���`���5U>j�e_��E�f���x�f�3=wO�����Z�!2#hX��.q%�8`�΀N�QnmÉh$��P[��$�4�P��a��hx�mC��1H��3-��Ӌ�2����hv+fK�[hu�+Os7�ێJ2��U�-��7�M��7�0�+�3�'ƅԡ?�T�C5� ���n0	�H�2��M��[��A���+y5�qF&��U쩋�#��e3LN�4�� (��N 9b��@�X��&Q��78���v��:�.������ԃ�O\(7�#4��t���I�>�V��iל{Z.��tR �惟��,ܻ�$G��������p�#�f?�e�"Ex�x��?��'�^��g�X�}wFݐ�}��a�F�nt�V���Ku�ʰ]��qZ����.�"�%Z�߲�U0m��9�ؘ� ^p�X)9��h{
�6���"W��k�w�ط@y�!7e-E�loA^�ރ�� +�S�Ã	��}{E��6v�HW&�mh��X�.���J������BdW������{YOlE��-�p�C���*Cb��"�<��?�_���>��W'>�{�/ �� 9�n�*xs���'h����0��q�:f������++>��0������,� �=F��	�/^{{8��Z?�R)�[�KZ�/�w1L'�R��Ԏ���..�H����\4��n-��zF��U�J��9i�Z9� ��U҉{���o�ۊ��pͩ��V�k众/n����l=��${�����s�P�T\���t2}�����i�)��%˜�,7 �=�Hk�=
�ޙ��
��0�Jk;b�"���#�=��wg��b�F��p��VW��@�
Z����ԭq�b��=g���: <�����}(�����`��	ߦ��p
��ޙJp�Kf;�u����{����<����P���k�f����%w�-l�Ϋ�`�Ŋ�ڛ��l�	�J�
[��z�dd�N���&����G�������k����ܲJ������t������m�R��-�G����}u����e��N������T�^��/eNo�S���1��u��N�%�g�'���)G~�yk7������v�/��:vY^�1�fB��.FM<���0�_�?�;3��VI���	�M!9#$.�V-����ѯ#J&���δ�:7�#tJ��j�^�x��9��  NI	W�5���7�4�Rّ*SN���1�Kى6�fӷb	W"k��t�C�(��4�`F_y�)(���`b��T��7�Ӏ��˾F���o߁I(���;Z�r�E��T��U��d����5d�,a���Q=�8��Hۘ��Z)nU���MĠ���]��$�C,�Ë�pk�<���J�>��9b�I���>�?�7���|��W�jW�N�)+t�
�*lV�9���o��kw쾟,�G����ʻ������M��7� UOC�o�_�聭�Z.����Z!ي�8���5z��yT!��g�=�����P,�w�ѿwl�Y*[� ��'�G���V����P���JR{��� ���q5�\�Ұ37#��o����^�c�9�%���)`��Q��҉������1`�p/��e�tɡ�&ִ�e�����mUи�p�O���8��p(B�|qF6����E���i.`�G_��y^cNѣ�bW&�+�Ш�$�Ì�rʳ}��I�=�@��D�d�+��W2�[�?<Fp]��Oأ��z̯�\�iJ�[����+</�q�]��/菃�;҃b>��KmY�^����(=���$�L�-�p�"�bSA�b�i���fK�{e�=���(�]�A��CE᙭&��	�yA��G��?�y:���p�,rw��!�B��+/��'�b�� �]�'��E�@3�M�C��sE���?NC �$��g�j(j�ŷB��LM[r�����箚*f�����-��M3���������Ĵ�#;��Է�G�lm�9��b�v�H..d�6'����Xm�+�^�ƒR�!�V����01 �Ţ�mwD�a��&T'��U���w빵�Q�׸�!��<晴�{��͂+Z@�!�@��0�ˈ�TI_�5ڥSˑ�6�]�Z���u����U6�@��˥���^ұv�/��G��R+?ٰ���i��"�
猌�e�Z�ߺi9'\�IZ��㹄���bzR  =���2Ϫ�w�a�n���_�D+2*ThQ�['��J�h'�Q�� ~@[�sRh*�
)�y�N��~�r���C�[v�	�u�{ �b'/���	N�BMd�>�M�u�(+F(��@��[����r��TШD����+�웬�[Y���Է�a����HJ�VYb'Z���a�r&�y�S���W������D��[*�A�ζ�<yV�����~n�3��OF�ZΝ������,ט���n��3P>x����=��@b@h�s�Z8��Xr��ŲG/L���Դ B�4�N(���F;�ZysbfYҌ���=�I�x�Z%"X 2�3�Ճ��b�d�<&�&Y�-�qѾIAt�����E���Ņ�tV�?fn�NW�>y���B��3��]hJ�䨽�k$�� Л��*�k<lS�L�Ek�j�oﬁ���^�.��t �P?P`4��7T����kD�� �~��A�n�o�������&��x�����ZX�zJGow�Y���0[b�m�TU����lkt;���6W>cq�p�p�sߘ��=��s�}&If��y�����_�Qr����c��mŐm��zL��Z#�c�|B{�c�w%�Ц8Q3%|ϑ�kž���.̛�+�l�S���&�%^����9�F2��O4�%(d05 .j�����_>P�|�&�KJ�+�	�8;q�Dd�m�QG{�{g��o�2�yUg`:��N��K)1h��#�.�k7���~�{��(�M����LO��c�Z��j�0��s��<"?��`W�Ш��� ����8 w� >�$3��
�ц�=��V�w+��xFnߨ)atz��)R��0QY��D��O�-��n��[�7��6��5�-�{���Xm;U�p��1I��e�����[f��8W�	d��ܩs��/�2�倯�J�6�#e}�h��ErDH��R�����\oN�A�&�8��h��bF�K'&�i�����ra�����*�L��zƬ�G�ZB�����i����7ywK��f��nC�,���=���WX�{�A��|Y�t�l���b���+�2.]�2�+�&ui/�.��"#��u0��]��go5����ϊ�
�e✘�����/"g ol�o�OLW���-)��;5�-`�$c�Nn�Jm*�����X^7��l��dN���5cx<\��G�	��-�w!?��,1�,�.���o>�UQO�����8�+т+�Qv�����|2S��O����}��@��4��������UP��'҅��� �J;?�Ъ7�s|����!��F>F����V���f�y�c�F
9��# ����˛u�%n@s�%˭<�pr�������J�f
�?�h���M��!���O��VCd0��� �^?$޺/Lpӣt)�)��+�eb���\ғ�.)*B�<~��8oϬ�t��AI�A��V�O�U-��9Y�ͼ�����f��M�o8����vC�̑�Y�5-�῵�V�����3kT��bk$n��ndP�����z��V7X/���c���oc�u�L\����]�rZ�9r8Օp����kd֌2w��.��>�RXi"��e�K��hXm�t��coqŔs1�f"lJﮛ��W�T!@΃�B՗4����/�[�̭ɢ:s���_��9	���b��p���QB��}�ڛO3��lԥ�m�Z��I��HH-��o��*�nv�8w;�V�B�Vd���zgP�(��h}�E �{+�
d�P5�{�c��*x��S�
�B Ի|�,�%�rh_�p�ĉ�ʢ2U��H�+��߆�����<��;���0����A�dGe�$��}������Gga���l@+�C��&�����+�Y�2_R����"�;Q\��2籤[6�pH�랫�낼���pU��mn�[��tX����[��_HuX�c��xӠ�?:�SjP`���g�m��Ѝ��JX!jWÌ�.�ۉ]i��X�
�d���d�D�<5���P����k����wʱ�a�#iũ���E-�Z Y_^+���99;�Tu�7~i����'.�%�:9����ݜr�a�� ���z��qz���5�:��T�3Jh��|W��@��r��ݙ��y��4�qm�a`�|5�s����0��e�dv3\;R�99Ëʢ�:�a���	A�K���g�[���R���E��l��Eg�L���ٵ>zn�Shǝ��\�X�M�3�bc�vT�8@4�U��=- B��?�N��a�
L�� ��g[of�F�Xb�l{�U�]�kX���K��̣�����c԰uZ�v��?ꂾ��>p���S����VX�,|�Q΂�Z��� �k�u��-�KM�c�o1��7��#ᎈ9$g���o�Ʌ���#1�.�8��uƦ�UT��5t�P-�A��[S�/�'f0�!��HT0�����"�K��䘰#�VąW��fҵ�����kNac�~�`�|CiZ��;�1�U�6O�$���a�b*/s�+���4ps��</�)��\& r̩��'�T�)k+���V�LX�<'M�%S���N}A��LΆ ۰�'K�_l]0E�1<��f��[�e��%�&]5��NUC0�>�G5z�b�<�; ��$�a�
-�_��rxne�|�v���r?X��'��\՟ �4b��S\7a������K�S�T�f8�'D;%^���/�ud؞'�_��>��D�tt��m�b�MW�ש��Ѻ�G��(�i4Ɠ�qp1�2�Dh�W��-��c<�8V)��kӾǨ}�~�vĎ>��0^̢�1�u��������e&J�6�Ng!g��N�����Y�"؍�-�v5���!*�V{v��c%�r$��))�h��9#�i�i�P��mci#���:gN4S+MG��͍N�$� �ϩ�&}d�lA����b�¹��b`�e����g��V
=A���^�<���T��W�Ǉ$�ͰA�"�&$�v�دt�ɽj0�I��Z���  �i�D�����6�u��3�k=n3pSk5�ґ_�x[=?v����������b�Z�ͬaza=�!	�j����\�"�B����o�p38^�)�Q��PX+<bj>]H���͍{��x�m���A�*����W@�d�D�T��4����/.Rj��^���)�|��<�*|ݒF��lɍ����d�C����x�RB���UU��:���O�.K#�W������}>]<���m?\~��