��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���� 6�:$���mQ�$��z��˙Y��ˍΣq�(jh��Pܬr��eۖ�����\ΈNt5��.�[�c�	o���kZ���H�Jl�F{���2�������[�u=�;���n�x��i�J��A.��>#v�c`�H�Y+��P�	~�����"��@�&7�����.��C���G�����`�4F&�[]*^� ��,�1�89"l�P�F�M�#)��*3ú2/~��Ƅ��j�;'�"����,����������l`��� �B���t�+t �����	�� ���k � ܙ�&���"�&�R��D�1߄k5��\X��y�d���=�Rt"�����ts�ܡ#�;@��?l��r��a��-j�I�%>�2u�W?x?�3B���G�Mp����?�����[�8���U���ݰ88��-ef)�;O�^�{�И���-�ݥ>Q�Y��4X���&���̆6����"�,,�b�uxL��#���*�m,��@�1��.-B�T�
44�8Bi7&��إE�w孁���I2Q�X(����*���%C�.@�"}�k�Հ?�v�M�1��h��	�$`t�u����#e�/�MhH;��C���<�ڀ��
��5�����pN�Z4d�����zw^���{)��W�c#�hG��n�y��6���M��a;�u�f>��sh!�9br �w|/~�o>=�'d(��Kc��e�3�,�6{�@����T�f07W�@����Ol��#ԉ�sŋ
��	����C���i�[��+��_yD�
�ی����E;68��y�bHg��r@k���2�'�_r���[���$���z>U��j ��ъ�@J�ۺ��l\SմM��C���l���1
���b��_����G�Q�ì(V�3�G-E%4�� ~��U�PƢĜ����R�%�9���B!� �a-���8ҫG{G#��B%�H�i��� �5�%h?�9ʥo�����c"K�����j;7�M[�kO�� ����VK7^(�D:�� �
L�,���]r߱�����`�����]���#,ʗ���4������[1�ñ/���&�`q�����_?��V+q���%c,�� �P��'���S�+�.׼�S˿ (;��St��ڕ�����y�gD.�ޘ�=����f�ƨB��濹��hb�o'��|.�����]�V���vδ�����O�\?��vK�E�r���?��.� �O�AE�.�~a"���խL��`�LB��݆��5�6�p�h��G��-�!�Z��bY�ncۻ�\��v�ą��p�\Z�b��PR��/f<���*֑q�̯�J������@�K�YW�G��1�u$`_.�(���� ���z	<>�кTc-I�Y8��Ng����x"@yN  ����'���6�m�w��'��she:J��\�V�t?x�N�a��<�mu���ӝ!%§�j,�L��Th��w5j/r�wH��t#N}[�����w�k{�-�� �Mn��E�IQCO�$Z��xY}�5���>s�����������e�2H���BjYg�z��dd-u/teЈx6��!��&�MjGW��c|���7���G����e�,M����fZ�}�o#Z�n_�yJ�i��:��^��F��|��~G;O9�K8O74��C<KQ�g����Ar���1_5;��^xm�b���f��3����Z��E^c.�7Ǌc��D�����`�)�,�.�
ԋ��ݙ���3/��a+N�Ghu#���yFʑn���f@���̗Ժq_xS���)�n���7�!����'N�zDn �5`�K��(f�G�L�<��I'����-m&��U0���&ۮ�]&��A��?23%�%kj�rU�������s���r�ۿ��<�b���L���H�d^-T����HiJ��u�|4V�TʪE���R W��p�UB����?�S��N��%�~K��=Nd�d \S7��Gb�LXl�L��V�s�V�֧V�X�]���$'9e���n�`���LzR����E<:e_H�h�R�\t�#@ԳNrb��bt8h%��y	���a��n��y�	�ϐꄳH(�ۆ�!'��gh����N|N�NG��]xDbj�Y�q"h
��,�ɦ�Y.�
-�D���v� �T;�#�Huɍ�i!�J����wD�ώ/�+N��O$gg�Kj��ҕBjY�(M�������Oş1_�@s��%x0;cz��W��r9W~h�&qP?�Zi��ؔT�S��F�ǖ#3-ց��Xvi�ĭ�{'�b�?���x:�J ��v )Z�?��v.�e_�� UNW�R���;�*�S�g&bk�em��4X���h3l�Ɔ���g��^�ظ���
*uK������! �܀#�m��ǔ�ضʂ��(*�#��W�/!�N�e	VwZ7��"�����غ���ŋ���������f@�J���'�[�%�I&<�Q웚��@������ڄBATU�MwcZ��2��6���N:3?\��O�}+}̲�C6��u� ; Љ�aG�����g��QʥE��	�t����7�M#)
9����'w�E�OW��)ɋ��5�� 0�?���n\�ύ�c��Rx����re,P�?��E���v�3�W-���q�^���~�jY�<<����
�s{4[��D@9;�w��|�-
Pr�ۼ	WSQ� i�=��m�mg#qp�RS0��"B��"��;0���߲��nYg�D/Ƌrp��;2h�Ī�f!���a�������b���5S�<�c��(�P�Qu���Z�/D akӜ���ɵ2/��
�/�9��0X���p��ڱ� Q}K����I�[@�cZ���܌0�a��i��mR�3�Å��|��zm�C�s���IJķح�M�N�*a0en#�2��[�2P���^��ˀ�,?Vʉ\�������\��Y�+����NuF��A���|���!��5��S��KP�Z|�JC����M��s�+J��D��(II���NKús&���Ōݑ�H����8ѐ[p��-?�HS�����v�+�YTe��v�~�}P�����ޕ̇��ʛgT��F��Q�7z�B#]o������h��C�·�>�i�Yv���Yv��ab��O�5�$���i ^��C��m��!zŔ��,�s���R�j��i.+��V���:GhZ���R��)�	�;h���(����ƹ���@���D��ݜ�2����&C,�:��V�{��ƒQj,`����&k�d����mK�؁º
��Y�A{�y��I��d_"K�5��\������_�X:J����Q;<͟].P�����E^`hE���H �ʘ���R���J�g�\�˅v�r��sN�D��_r�j��������Z8��|��hvHB�S��P��4���i&��r���t�3J��p��eU�����ć$Z�s����Z\X��Nac ]'�����_,[�i����}i���CX���\���p싘-9��3���B��Ҳ^|�����KJX��-"�l)\e�;Z�v֔&3��'���Z��;5Ӯ蟢�S���Ӵz�1���"�gGS>k搖m��w���)Yq����%ZuT0�`���,_j�cu4Ⱉ�C�ܹA��S���2�Lz������ .�;A��/YN��rg�g�ԏ��׏Sa �Xa5����Qռj�a ���y&3$�a�����TTπ�TC�Q�=�"����6r�SZK
��� �1��J�"h�jP,�JI�[����,��=|I�4��0�����x

�+ZK�l��ػZ���/��u�xIuGz�@MK4�`�o�!m\u,	��\s�Z�;���z�z��2��a�k��/� rd�p�<��q���)̀FB�{9�
��G�t�����rOU�@\k��1#ny��
�L��#P��ML��*{��O<Q�J� Z�38P=���핰�ea�[�ڇ�=ΊT�&��)g	D\��1RE�f���|�A֪�
2H��pR�	�<i�K�U����чŻJ�F�[즛.���>-ޓ2�)m��x��߲7����f�Y���!����5���^N+h�B	�`��ϗg=�H�7	D���c*Ix����W�Ç<��"eXQ�˅q{�XXc�]�?v�F`PdOA-5����h�����e�p�E��Ez�U&�>��9���U�����C�B`�+]��Mi0)���dG���:�zgb 3��A�@_Z4��t�gB=J{�Ϛj�؈� ����[��
�I������=�Ɩ����o�fg�M�&�ә���z��HHcj#ﻉVݶ/f{�Q��[��p�79����6�J�J���3NO��H���S���r�f����d�DZ�`��K��������ۇ�Z��Cۅ�J�^죜��T�x4G�&ى�yF�����Z���0I����Mro[8d���3���`H�4N��r��u\a�+�/��4;.��o�	O���x��f�1�X�����$O��t�������7�Ӳl��c����r9�W�ϙ��m���P��O�aR6 /�����@I�� �o,��,&�]PT�����ĩ/e�~ �apc�ы0j���'��;$�6�%����a�X�9�x�π���HF��������u.�I^@�� ���9��?���o��FJ�?�n��B������'<�F"�V��NҴ֜��J����ftsW�������@� �4�Cy�!
���=��\���鐱�u4�G%��$A���q��I ̫�� �Ab���m�ۘY䥝r"*����6B���*bo<�,f�4�!���4A�Lc8��x�7��f�\l$����5�J�ޟ[SZ�"m6�i��s<�-���rP���d����f3>AAP��ֲ��d���*X��j���mK�u���<��Uq�"Q�D��� �#�+5���u���f-g쉉��l�o�߫��?��á(��G8~�
u��ޜ�0�7���#)w��IZ�攼��RHY����jR�Vp��p~V�������>�9����~��h:B�)�nm	�:�!�?Suz��"b|�E�/�\��I������ Ҁ")������܅�A: �3�)��C~�w�e:0�Jm