��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�~��"yAfEi�)�����B
��۩C4JA?ϋ���n����g�ҕ8[���!�܅r(�=����UG�O((�K�`�0�t�s��hP�D)�w�xJ�[K_
�ԈYJ���LݷV�2�콷iF���}Kq�I�q��h���H�i���m�����-�bH1�)��Z�ٍ�jӰtr˥V�ڥ��L���|��qѷ�&GDq��ʻ<�����n �Ꝿ��d�T�\j.+�wH^E����C�]��b��`g���[~?Ӷ/�}3�oN��ѭc�2!	�PC������B�+q�z��*����� ��z^˥���ER�J��d �-+T��o�9��h�:V�%|�]�i�E�GJ��4�G�xn�XV�Gü�g�4�a�K����ѥZ5j#��T$3�"��!��K�jt�%�8��2�Rk�h�ﾃ�!�����B��y�����W���&��&0��ɜ�ࣼmZ"�O��S���O{o��6�c._�M�TĜj��[�nń��񡗆��d�
�N{f�Z�ú��e������=M��K���������<��/:�T� �H��c�d�a��[�ӧ��7A�����D�;���Ŋ4�>��gґq��xʱS����Ogt�r��j�q}��߽n�M��@)�L�q%Qe=�&g��� ����d �:�d���^=7�O^��K4�DW�PX�����h��~8��a2PƼs�Ky�����G_�����I)��C����[�A�j�!����dm�$�AGL#Z��$�e��
��W^Q�q������b��bL`y�Z�,��p���ǹ��_�#�I���\�b釭M�� ��=�V��Z�5�Y��D"����2����-�̜�9tKw��s؆
4�gi�[���;e���*�N�a�,Q���Q]e7���yZE�%����f�z[%aZ����=���,Օ�RHޟ��V:��K�^[��`�'���`��/����t�)U��#t�����zS8�Ɣ�T|rl-ᥲzGr������ͭ^����Ϝ{@<�/�E�2�%2�I��<����(�c���j�B����C�b���g2ʜ�-xLo�W�ܠd-|���_k]��H�i:+��������2��u��\�*�k��|Nu%�fo?p�;��^�{���y��\���0�v��#xʔ��lۋ��\p������\�����q���K�I�԰��|�k{̱�����Biū��L�v}_�d{�<��a^)�f�I�u�Y����^F���+d��!v��Xy=�6�&��L�/�[-ǫ�kF	o>��"|��R!*fX��Ez��������nEs8�G)f�2*&@+�s+]�@=��2��ؽ1�)�������$��7@��Pde������=���jŃ�?�H��TYf���L������¾�������6j�Mg�������CL�l���ֈ�E���7�ڃ�CG��m7A��-G�5;*6�7��m-�ZJ�ܕՊ�dhǷ�Z��&jS�lts˺U	&pu=���_�(��r��ƞ}"������M]��q PGtj��� k�����vD�,0K��ؓφ�/��tl���/9��	$�S<�!�A��QF�e��-G�d̓��P�btz!�o ҊFi��)�C�1�����sL�����?����k�E�8���z�:�g"��u%���PO�@�C� ԛ�r�9���#������$
��11��jp�z�0	`��f&�A��E������aP��H޹5��ߕ�CW�,&/��l�M��a�(��ww&4J��7g�4x-�K9_f?�f1��Y����E��UGȠY^�?�5?������5��I�'_�2J�����\�#���fqȘ��:����GY���E��ΓN}s�Q�g\TS��Y����o��4�pN|d��x�]7P3MN�(�"�I��?�=��v�M���H�0A�2q����P	��
�����%]K	��Χ�]C����&�d�,��Q������܈~]�[6)������u�1($u����5����߳T�&򾂮����Ȗ$�7�q��P��2��o�),���H��ÿ"Պ�A��j�{.����J\�{y��1޸�[��jq���F3ȼ��=�O@^uK�45������O�	�3���m���V�����z�$�Q�UB�Yn��4�˱��tQ�N�dQW|��ӥ�|4���=`Gc6��\Z�J��½�fó�DG(x#���h��j{I�ǧG?�L��'�F�@��ו"�W�O�6�*3�p&.C����ND�"����o�b��7�'�[ ] g�H�����^%r�
�G�mcU9�c����́rez��"�*�?E�U�`y�]��g��ǋBAڰ��OsnMP7���$j#_��*}���&�ܪ*��ۧ�U��(6R	g��iq����Q���x���\c��:~��hw���O�72�u�ޥ-� �36�����LV�b�^����l�n��z\v�W�NMya��@�lt�{4גҀ��]��[ĸ�3){�	yM������!;@ci� )\IɳC�/�'v�ڊw��K����o�xgz���Yk��H^�A9哺���sw5��XVp��8���F�g���Kq!�ge�̩J&�C�5G��>�*
VɭȚ����_���/.Z��p�1�.��E�A����2�s/r=�Фѵ7,f�������oP�lb�T!	"����om6����|n�2��D�I�mLchd7��[p9O�C�yխ�E$T�T�	�с�XF�G�q\��T6;���ce;����<7'�V� �$�Ӑ�a-ӷI�D�D���ݫa<:]d������� �|����-86%=>�%.��3����Y-�_F��zA�dH��k�Ơ�5��ތ�BKB"�M9^RII�$��X_��� 5ʖ8�ēţ�l� f����kK4���*�o�5�1G\�p�e���I���:-�~���-����oY�M��d|)�a2�s�~�x�V�~?�V�CW�1H��6��Ģ*/�3�+A��������5������<R���R���(V}J*�w@(���k�o�3�#D�t8v�]9��8Tع����.�a�Jeh
���E�ҏ"�,��&���\��ڕrA���q
n��� �	P�ȵ��X�.�K�-]�n����1���v#[s����-h.g�����N��i�5c!X�$qEإ{˞����E�y��p��:a�'9���TX$�a~��D\~y�x�m�f4�f��hk���@�L9υe��9�����Io9�$�^� �F٣�Z���<f����+��EC�[�n��\�܆i$��]t���5��B����?�d�į���|��Dr��0���>s�'��_�Z�pr$�bA&!��0��w6�8��n/��mo 5^�N�.�g2e���8��3=�}Na0F�F|�i�l<��
҃��{�� ��R �C}�?+­c�8�.<����\��xD����bb�q���\��8���0R��2�c��b�ĭS�w��9�d��������)e<�/e#	NR���⧅hc4�D<ع6��mȒ�:�T0~��Ůx��8�3/�x!zL�XG(0�%��eq,�i���$r��8̀����ȩ��/�X��$���}�yf����&M��K�s�g�[���n�9;�m{���i
Z�騉��\,��l���Q⥌@��l��̩�#�A^�o������C��A��
�Y`'�~s�
�w��`��:ى:�Y��N�;3VIA�g0�I\5-���bNS�s���ۡ�`rJb�h*�C�?f�,�~�0��3�~�UNJ�vdev�3!�	��C�"�����Ҫ~�C@�[�d�|�F���j�=���
&͞�*�71�>H��e�5f�Y1�s�ZqY��3i{K�ͺ���cL?g���{��� 1��[O����8�B�˽D�� ���x��d�������6v�l�z_��7��~yi-��6�_V��~�:�o�Ub�<I+�ヵ�1Y¾�hC�<�k�L��P��{�c�)lA���]�7�s� ^�����������6���/p�F���k�X�҇�X4m�P��)D�.L��ki��q���&��3�q�e Q{Y-L���-؃t/}��\�����c;R@�E)k��V�ºk�/P�u��)C�YU�&w1?Ҹ��!���1W�+�xO��=,JȧdK	���J�Ϊ�?�ۙÈ��������g�K�a%V � bQ�c2��!��Ț����>��煕�s�P�|O�4^�_1w�����}]�w�2�K��4�{ڱ.�»��n��������x�Be �v+����n�:�����em�>��qGڋe�A]>�54QJ'�8���s�%�	°��1f�>��Tc�8��|N�����~���N�z��õ�a����\�������'�ei�ީ�γ�\/`sA �j�M"x��9�u�D�" 'IS��m��NN�u� +$Nji+�<�Ě�l��o(3�-��gቲ|�Ĝ� ��ѵw���<L��ݽk�O
�G]��t`>y�+-I�bKD�Th�.�
+5Cݳг�$�]��/��C�t���ena��elW�PU��oH����jH�f�.��z��t�wy����D�������;;<�z�M}�N����C~�10^0gי�N�m�b��� B9��V�<�)�R!MCKc�TG�͓�"���T�,/@]�}��׶Y�'��:�	�#��d#l(-�SB@��\���t�򪙲k��e}��������J��TDV*�N��C�y�4��*��TQ��Ě�U��#�h� �J{.��%�:���c.����u�h�����o�U�Q:�m
��!���lt��JXo��?��8W1������Y&S{GTZ�%G @Q>-NB�|��Y�g��x�U��ɇm�j�o��<̥/g��-C]ӯ��c�"�j��ܷ��j��ឺ��N=B�-�l�����M�R���Ф$cڭø��K-����AQN�=T��A*��0QK�n����?���N���[�mnY(�8��A��#e\<9��}@y Do�#�C�#(��oKxKP�^{�94���V�&&�f��H�wW���B�b��:��X���}P=��G��Ξ��s�%(C����i��;F�?3�Rg��n�״� /��L�E{+�UppN��E���n����z�Z�J9���;#U2�"�g�%E2w*LC��}�����ܘ��S��2ӎt�J�&�iJ��٤'�KZsQ SI�1� zQv�R� �v�ө�.ݨ�?o$I]Z���M�9i�Cf�'���݀`K���Y	x0���U�	BO<�N�A�z +g��j��'��9$Q(�p�;�;�Ҷ�*M��ɂ��S���g�yО�@��������]��|w� +p;|B
�R�Q��M�7HK��,0�J'o	�&�,�6�R3������:/Yy܂��X)T�b�-�|���cy�}���| �:�f4�ÍЊ��<��;�����H$2}�+�n��h��c�3���sa��YL�mz�71��&�+�E�}��j#��U���@���
����� 8�IQ��g��I���HFqY�Û��`pw������T�E��L���P�E*rM�����w��eft+B�:�KΨ����1d���5�Ѝ��%2��$+��?�nOv��mMX����y�j���w���*�����/G��ّ���w��5��Q�qp�q��<��A��GP�{�a)��Rj�v��eO����xwmd����'�j�^����7劝�t��<N�"NI��=,���{tx.�;��c�_��mL� �nX�p9FyP���,�{P�>/�����Q�s�,{�V��`[{���pK��[�`ьm�T�名��5�+\.�  G�ٚR9��j�wg.�{om�5�D:����@����� ���N���h�y\[�_+�L�Z��Yt\�R�Yƍ�5��v�})u�U�ĵ�r�ٕ�N m�!8WG��o�-�@/W�{qv:��ܹ���?s�0�cxB���k�����lh�w�	x����ǭ�?W1��AYytr�f8�Q�~z�[_G�OÁ��.Q�F�6{��vje�$���2� �r\�Ъ�jg�!���;�g΍G8Ҹ.��7����@t;}�!c \|����<�\�o5z(Ӭ2{4�� �N}�]@�E_ފxW��@�(T��<^�����@'a/���R�<\��X�C���|�-j Q�KW�7�����s�A=o�}��
�@��S�+*p�{���:��p�2�BaD�6��'�D��p���[5����J�b'��������,��]��7����_Z70F��t}�ӔA+J��a��|����2�7�v^�\to����:���;gf�R���q�K��qN��Ȇ��z�A��6=�b��j��_�U�]���_(ZTS Ui�ݺ���:@��j��fr*y�3���x��h���̽���?A��$�g������-�B�)M�[��l�{����W�.� Y����[��I�Dq'sw��{2^26�a����\�*.WL�YT�(�2S3�'%��//������@�=��y���n�� {�:?6K�z*��ڏ޶gR�P��]���1�JǷ�Dn��e�/�������9 ��R��đ�q���d��uWvѼ����Y�O{��-mO�:N�C�� c|�a�L�4IqS���=�]�F�E|՛t���	2�N�'���悘a0]i�T��<q %#m�dK|\��<�ޘ��E�;�>i���RK��`�����~ta�AiD���8Ɓ�^2���@��sv!�n!P_�SZ�ǉq���ꯞ�"�IdέVC�%�5(��ѵeL7sG��7�3Q@v�3JY�s����I���4�>sӃT��{=U����g���L�z����)��(����9I̗��&n �޵���Ha�6��I� F��O�񳑴k�l�]���N�Opi��`4eʽ�t�nBv>L��0�W�E���/�&�}Z;�&�bA�X��xj �V�~�y��An\�(��%Y

�I@L$�Y�t�]�w����S@p��;R��~�w]r����$ɳ��Xkf,�. ��;7��޾���M��ҴO�ҦP�a�$\ú���Z�ɔI���2��]���!�}�~��]=�u�T��b�1,0P��f�̮�̗���d��g�Z�(\��mH�X+��7C��%D�R?��7��7;뛬U��Հkl�k�Ät\������j�w���B�������kcг��I���9�T��%������ʊ��zj�-��d�3!�4���ەxW��e�C�JϏB�� %Cnmn~�Bx�h�M��Z�p|E2�g�\K�jh8>L�rv
��.�{E6:����*�?��䐟��&�f<�q3��I^òx��˷�D�kv�e��6S3K)��O4O��/�/�(<ǟj���<I��7Qj  �����_WJ*.��>C4���wK��ǧ�K7�d�.VM�w�`�s�,O���
��*�
�a1�`ަKMT�w�\6���/�rӈ�:<'�����A�9a��	�έQ,����-�f"��qf��ٮ� �K���[V�~�Q?s��o��fƄ"k�@��u�l9.61��(o��S��*��������"8��BP2�y�3�|�>=aΰ�Nt��D2H���$<��=��s��l���:JJ�݊�K���m����h�S�?v�8�E�c*��M`�a����-f�O�u/�4���&�t�X�C�ME3�I�o�p��m:���%�̴pnC^�mw�r@�LT/�S$S�kk|�C�<@����O`�5������s����� ��Hf���)G��n��B4( BͱX��? ���� @~�S�*�v0�|4��/g����r6S;!�� �t�$9�(Ŷf�V1:R#w��ݣ|*aw��y�=��q���G���Q��>�J��_��R�2�#��0�����'��|SG'B��^�����e��T�������2���e����Q�#f��h
K-P��Ҕ�B�D7���mP�����.$��� !	�̨������PV8"Y�HU���A���d3,�n��^�@���nTi�J���|�e}]f�n���$��&[�,Wb��$G�����/rQ��T>%Ը� �^�lC�����AɏC	�=���C�7�Fw�`��X��_��ûv�5��q\���vA�S����Y}�UU�*e+xh3q�.� ���mXB��+0a,���ĥ)����l^�y���;��j�9~����M��7�.�s�2i�["�>W����e@y[p�H}?�ǭ90 ŏv/��;Ԝ��#4�P&7e��LC5�	gE($>�����k�A�ķ���Jܖc�Ǘ�Mξ�+Z��E�CƱ�آd�M{#Ł����E�&�( �'��8FY4;��3��\���]��p��Q̽w�������-d��Inڤ��`�?RD�(�u��V�&���($"�)�;Y�r,s�(�M!�f��9����c�.C�kr��1�hq�ɠ�`�u.X���w�`��v�MP<����=:��|r�����T�)��d��4� g-@d��_>'�'�'��&G�p��2�]�I:ai��!땳��W8?��/У�8��Ǳq��,��3�O�7 ���������L�`�́�X�H��='nm���"!�vE���":����0r4�q���d7�yz�	�����H��v��R�Q?����_kJ�2�)��@���\	�!~�)�"ξ����>�J)|hk��u��?s4�
ڸ�4�H�u	L�)n��Q��`���\�b+�Q&���N��7kE���Ùj�y՛"�ךI({��ϰ�c*������#|�0v�zD	X@ڗ���X�#�<�,� �6��j)�NM��{(.�ĨJ�#���a�1��6{<�8og�ex�AIX�1��GΑ�+Azh��L��]?;�ag^I�`���]�Kjb���BSU�������^ʾ)�_+��\��Ym��Fn��j���������_e���i}͛!Aw�k�����n��V�U�~����<$�V��ՙN�9�ZȵR��IWh�9��iJ�(�e�͘{���jt��Ӫ�b;77K��v�!���L���k؉:J'����
OR)����{m,Q"%�Y"@�Qʫ�	wF�B��;�lX��'i�?��uf�2���V�
svV�� �E�m9K�c�� Io�sȜ�D]�S[pK\U��%�P���w��4�� �c�4�[c¼�0��9 ���2�f����xH/Rn��P��2�k��p ����w�S���e�L@����c�!QX��G C���C
�b:D�2f��>�X�2��P��)EcOt gdȞ7�7����é)H�e5������[Eq�N�N~�N^V�����]E4DB\ʥ�2�:rr�J�}��1 C01�,�d��.��Oǘ������@�=q��~��j�m/�g������9Dw���bż�q
@&�����v�Sq�����W�n ��6�iÙ���F��%����Ү�3���>��L��W�2�%����w���,rB�4��.U��&���Vy��'�f��!."ѕX2
�؎�K܇�_X�]�7��'�0���v\�t�Z�
����x�7���tG[���Ef�!Q��=�BƌN��9?�1_);��2�1Z�S�2x�����l�|1��n�������T��9�<�mc�g�m�ol���Mk��xO�ċ}E��N�e"��+��
��1E�~�y��p��FJ4l�]���f@�O��oW�%&Q�AY)_�ݛ A�c�e־D�e�B༞���7s&&,:a���B{�ve��!g�r��K���$�t�"��أ�yc�_�tcg0'l�j�7:��Q.��J��Nh���|�v�R#�FK)F{�)�J��?x�D;(�ȥ9��8{UG�ZHٯ!1�Ĥһ�_�n ��'H�~��Mj�r���N�/0�U���"����S�7�(_�k ޠ��um��IA�٧�6'�hgo�}����
me�G���H�:��c��n�w��<�yK�ˎD ��9�c�%W�6-�@���鄩J)���c6Ȼփm#�Q�T�%م��Y�+h�࠱�E�<5r��H��B�J5��x<Z��{�1�:/�7�)|L���5R<@·כ�zy��eG�8�9o̹(+��+M1�����-g�d��:�[�i$mm@2��0�ƣ?2ɻ���:u� =	?���� ������ؑ=�����d�%�v�Cbh�y�V(<������4��gG����*��T��F�<r��}W����e4�?eG��/7��x
��#
�Cy{-���tP2d�?g��{�SΠ\�`���XK˽���?>_f��W	E��A"j%�[{�1έ&�x���W:+O'뮾炌㴝�m��4�y�,��v���/�ǴP%s)e3�CA�[�}��)vnB��qz��_����.��i�1Q����;�Ͷ�A�NҐ`�Ls�5���=�����
9�#�V�6vg:�"�׻[�R3��?eP�����"�Hf��@�`oQ��˳7�o!z�x��D����g��R�S����5�?��{��y��@��玖�.ɭ'��Pa�k�F�R��oa/�� )4�v$���� ����]#Q��J�C�P��#q�Ж��J�d��UD��㟅�	%��?ӈ�� �(	nQv�C�,�ہ�<���f{Vk�ג)I��(��L� �өH���MUf����_�͹��ܠi�Ř��U@�\^��QAap����t��wx;� �h���ޯ."��i�x���g�i!�.�	�#��ʎ����(����i�Z+�t`�2�:lT�{/o�k�W
F�>����UP\aܐ`�;%�����)��~a�&���{�20����n���U>�x5�%��|o�ڌ�E���%t�E�Ϣ�����	ɪq��ܰ%�>A��G���ZҟZw'!��)�B�2.�j�n.�eV\�l��4��K��Fu�z-��4Ї�z����՘�0�Q/�^���w�(BU�(ǄyW3�T*���W0���n�&oy���?b�
���3"Ag|x�*�e����^jn�W�VC\	��r���}M�ow`�ɾF[w���iP��a+�D���ŐIk��AK�w��w�.&r�Iw�M�ÅB(����ޝ7�x���hr�\�!|�3��sOH�����jD%-`y���NȆگn�s������ �#�K}�}(65VC������c����\O��[�ڴ<-݅�&&���c��]��dG�䋟�;,`"y����\���o$R� �2��p��lGH0(�H���
�Y���?���BXv���4�O���� �=(?|ͅ iSKZ��L�׶���V��O�1c��S,��Y����H�Kqx�a��{�i�~���w�/n����� ?4춟��{]#��R�q[���8>_"a�N�O;�R��{����6�渄�8�R=��p�)� �ڪt�6��:Ӯ�k!;�:�*�%�g�`���UB��~Z��>^�Y2��4]N�)���Nւ��\�D�~���	����Cw��)��qS=3�[r�Tb2X�B�����j�ϊgA4��]��,�,Ծ�,��\G�A9$��XW�pCKû����5�9̯��u ��5��@ת*�"J��'�`��t�,P���(�&� �)*=B��W-BP��xp�Ң(c�E�����n�P���G�&