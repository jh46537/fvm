��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ� g�I��Jw=���c#hN�j(r��Ҹ�@���{ zM���T�wY�Z1�����I:/Ҥ�����	WMЍ4�
{�٢(��:(7�p� �[4	�D�}�*��z��'�*;J\�������y�Y�!9�;��S��H�4ͱ=iT�����r�Tfg|���*A�*zA���] H��H�7��m���I��:�.���?���j=�N��;J�<<��㌱<_^�1c8�����?@�"3LG���L^S�S��qQk��akM��ݶ�� ��@O�`�i�\��9�l�6�{핹�r��)�k5v��^hQg�@�S�)����Bc-Y��I.I�d����z@�pR�e��Y}�sf�!�SΆ�����\���.�xH��U�P�پ�V�+�J�Xk�i+�>�vM+���޺�$�.�sl�ʯ�<��]�7T�.� �]���+��.$��鳮�wSd�([����.��-T�(�z�1�-������5���y�o���{�؛��?����'k%l*�
`K�"z�i�"�;IQ��'"�hpɞ�ȭ~$��Z��T���F�(�O��u���mܼ��3_ŋ`ȦX��"�A���	���$��!|\aQw���OHK5��V��$�<��q�d�7�M��%|��hǭ��١�Qu���EU���\��m��J��&���s;��o���%��{��r>��_Ѫ�$�����K�5�Ii�f~>�����"Y�6�o�t��ok.�~����Z7����&�m�ik|�p�T�DS\�-��LӮx;i��Y�n�" 	�ߘW�w��k��t����(�	k_, �-��J8��fQY�I�g�z�t[�F�\~� ��Lt*,�H������;g�Z���p�_��G��}�ED^���7`6���X�R~��2Ur�%�$SL�*��{�S+=���p���[��� �Iӌ&����W&��9��ˇ�ь�ܔ����a�����bF���%�3C;p��)N)�E��,�ʗ_�)Qm)`�J��Rɔ�dHj��f"�y+)^�:����$-��]���E^��3/B�i(���0j��F�������Ӯ-��e+�>U��'	�Q����'>������`�>GRbDkfj�7f���;�Ʊɪ�����V�G�=\YĔ��n����Lra�G���meb�M��j���W�9�����-��������#�p�ݗ��3�_�z�f�g���y�@�1�"�SB���oƭ�я�Sܳ�,���������e�M�x��	5���'k����d~}5I�qf���/��k*���hG9*��\�f�ti܍{X0��ƫ�����W����f��H1��ɽIĨ�+��+Ϡ� ��?t���#&�jE�F#Ƣ�C��۔���=�`��5v�uX�8�B�4MdE�{Ӯ��!i��\Ŕ�]w6h�5��Ԟ��p98P؛���Tϻ�=�1�z}7��� ��0i�%��{:&Ұ�V��m�q`ߕ�vtv]�gY�3�<�:!mŵ�[�Ȕ�x��J2���a��RXw���6�޽u�AsL@Z�w;�YTjk�g�ni��7�-��ޘ��A6!=�#���z�_Guz��u{s3� ��Z����D�Z��C�c