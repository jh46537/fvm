// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:17 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c7oHIDY14YmFCEW7SrC5O9kAFzU+E4QEe/O20AJiOcRmwW0OFuPfeL44qTZHkEmh
h7fJhU6aEtiTIQ2OkdiIuoVuwhQNL8i4EbMohPEqvlGKQfDwvlqkipwRO9TdWCd1
fFhmGxAwnE/OtaXA+O6Y+ZdwgvMziPe+bH3NakN69uU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5792)
152lqvB/wkxRUS+GUb0nu6NOKAybFvEwLg4l0xxnDhB44IjQrQvGZO1F6vb+9LkR
6O+YVDvVOEYOB7Czs6rQlU5NBMx3O4zFdGgObRg+0X2hzuopHP8IpgGK7XtJTHde
KqISrLTt9jWBiCqDYsJ9XPWRrLsI73mw3oPorxKhmbnaux7+NecdeYNFPylZJRwd
B+jxQqSIbra/70q1SK/6aGYTtQycdFutC5EQsDwTbL2ttoPPnbXrVAm8Jkb+IQ/4
19dH1kEFDj1vIFY7f7FXpvxTZPQO4Fi58D5ST2qnWgV190KdsV6Vad1/N81vfTFO
xm/7TngczghZjdri9jZkb6Iveikh4MtM151EsYdr1ra4LctS30n7vyBPVcFtBRXn
tmgcBM4/ySW45adQbte4GFbPERK3lCDHJBDxa/XhFs4fiutIihTij4vrRNtHAhWM
Ryc568S0TJJEIY3rdTAr4Cufh/J0PSUsA8nJ9Ob+6MLrYBy1jLCvgOM/8AwiFKaR
A3LpmE7D5fectE4jdMVBQ86giszwZ86L83c4FMwC7YmJ7171yxSDduIJPXFa4T7O
e4z6j/QALjYuEYMyN7Uwmnb4mdu71iCyL2Bql5eDreUdDaNUXhGQ4cGPD92GtR0A
RxIJSj1nZ9gg744YW3XeCnolnF9OkHfRH2T6n6oKzoiR/36nrvYsOgDTwz149hn/
u+FS8qNt7CM5dRx5Y5CzGpfqZbx4/NoHvKz+EhMlYP8FS2iP8/PJqdzu/kgK53W+
i2XKvrYCZ+l/LBhrmyjLBzObOqegH/tUR04IvlQ8wONLbASj0pSJ7gVIJYBHcYcE
SmXSwm5pr4NqB0znfB070kzIGjHgFkIDG4+FNDrcz5I9NZ+yMOSMm6yC52BRvbXA
TRwK9XW5NQQZcnC47WEV1Kcx7gI0turTVnBZjp/2I7sxCgZb1KUC4Ed1INvCHCZ9
7AB4E07s9dKyBDSXfRS3+Ed4Cf/PhPN/egpuFNoZgjRsx86vfgjkaDFOBJBPtq4s
T+nEzZTOrPGZpdGq4ukIjwZ184nfmlsEhewHtJqb4bl0BtohALgl9ENeMY8mwuLV
yclTWsFMaH3hEqTCuYFFteNuy3h44805OsCUdUikB71ZkchKGfPpI4RSVhC3a0po
j4Ii56P86duFLc2y0n3N/3QqE/ig/mGkJh1M7SKnG8o8obQ0p8XCz0bb/C9uu1JX
Dcplo07ZLF8QivgwFjUwP01Uo98dILd+RaAW2H87h1Wwsi1dhidrUk2E9uFdqc92
2WiLV7jnMsm5IQADRXTeu5veJGQi82XF0szkOJyrFW5rUiRJIZ4AdRKBMBIa44Mu
iD1MPKPOGK5fOn0SkcmQSSToUNWDAZ/rcGGbL+66G7b+VpkEAgieofk6Ikg3D2Jh
eoMKMredH6uOqfCQA8WuQzUe6Q4oANTzOdRZvVRLahBmpUIgshg2PNGnemOEhCvY
ZZLiEo2zzcxKyDbg7oiIl0tfUtj4GASWTa3LYydG9ILkJ8kf+WsGjE1PdjrOcyjS
ndLiKP6Z9B+O1PdnX5R6syw4tsGSPAaXTQ97ds9nl2kyB1UdtyNx50fe0g1pyRDb
5j7uuI19izWo7b0zvgUS6LOagBfSQP1/wNOSvENYmTmhJqvu8rFL0yuEHZ7s3Nyc
N1u7yiyyHJI+y6Zw0XYQIuZwX1fF221qyOYjLCq3+wc9dwalFyCifYzDXbzStq8P
adzEddzh2n+cJSppvzmI01tFpaDTPY7EMHVSozd93BwAJhPPNytS2fDUHcNRPLRx
7Tnj0jOiosM+hSw1KIwyBiCzG/UFDBn40A7BXLL9BJeMe3c8eQrnOKbqHxxy7uMw
BOIfq1Jwd1Q+qrdrG0s0O58DpH6pTeINqx346vudt3kuk4tlYdORq8lCxpWJb6dY
yForhAJupjDLyqa9ymcrBMn4q2fltBAFWXxsJVA9kRdvsCqcXrwu+RxIdsy2T8JS
68+56WMViNvMMDTVQ15e+kWteJ2egRK4bd7yH0NwGpBYHpNQARjCFJCmzVbI0udM
Bz+lXl/BHwpkBw/J82LoerDUJjlYWidrCzGFIQtzL21mTL4Y5+LJ27m34efEvMgN
fSQgpwhygWt1WVe2fSPWQzoU67IUcWJUc/9BOUQsL3mb3/ZMEn13yMOHfhdTmR8v
SPE2XwO3sDzh78HsU4zw3asNONU3/G/X9TyxwIILnW9niggMg1yBX+F42Miv6HZE
UIqWRwxbcRpm9l+oQMutqlN/dAl+1l6CxKRQgIdhIAkI5qqtGjBvtaPxZuEh4ads
jFyffHSiTPpFbUST2FEuCQq1F92EdeFO9wXntb9fVgbkzKy8f6bO8fwIrLNBMiUQ
GysMdUKP/wF3N+X0jZDuyOkyfYgC0A7XxiCCdpXz7UcFJT2HCq7sv20PkcjKy/P+
VR+gg5CeIUUxMJq88HwgyfBe+EaSa7wTc4hx2jbE9AMLTBdNQdkf04p/6GSZoZMl
cMybH6Jxewi9l11+KjTScRj+rRCq4yMdm7weA2wsIFS+WCRjFZzUss7cdNBtAt54
NEJuO+G/0ecWGfVC0W4Q1TMZUNHiObfNoB37nwCroJ2+C4pDcIuBPFbyFFzSq9Lp
Z/WqgCIt6bTGM53tp9+8X5w2Wu71NAfMwBvRHuCynLc/NSTg01vBDSYfayJT08FH
c8GlzBEw/h4oQAh+Mk9j3VqP7Qa2UaEVEuraegtRJj2OTjqQueO/E8NPD+LLnqpA
2oVtPByPOm24sOd0TQmxXuGduxFjrTMWM1rmKErRSDwf09OfV4aMtwImm90Oyl43
++RM9v84lU/WDkYgktkQFNvz68oButJ39Fv2OdijfHaBqRJzj1YuB3KrSgb7fWv5
qkjX+up3zj/Fl+gcZ8WttDWie27K1ur2lgWniCToA5bx+0KoV1ureNQBGCrxkHRP
VlycUOJm79k3APf017bGMWFJr9dcseS0Yeh9I1T8Q+CSZz6T5SxWPWxfrxPppf3p
FlEtgouwUEI/x4jgBmLEi2HP8qhdTOsSOeY2V2LTZrDk333DrdLw9R9LD+AtKwdD
VgFhUIRxe1Ul9IEclHyBVRr7KZcf3+q2IxJL0nadtfHEJnsEVwHTmBiZ9J7zvhit
IzRBT4LZ9UYxN34MtVYvx4VnCvDq/UrhocsmrVzLf20K+OadNrmoZt5WsNQhjcii
oArC9ThbDiPysgGWWEtpL6mAjhXLEZl6AYmjkH7w2hUhNQJ2apNNxoYIuLcGFhpu
+0nOw1ElL8FsB8d03HHdnqE2HqLo00reEKDT5zQtq8exwY5uIP+Oj3CxPtbO9u8U
qTUvqqDlOttplWVcz6XLkYmfA34Dm4fOcCWUKoCNMr+BVMWPueMTZFRhWp97k0Cz
9eo+2Zt7BlnZrRKm8LI/FU8EWtEU8xbH3NZcOTAr91lwB6KTRXhNaklimU687nEx
nctHl4vBtuLciNrKoFbxW8SY0/5+8rluZa9mdDkW3dLGtClcX4UkT3GSwO1RKJWV
KXVNPJQvR1h1MBr1CYK79MogHZyTchuF3u4zJYdRgWuyU0cQ9RIv0M+XxuQ6dUsK
Opk+ITCHy68r84Gd9E2LnVOyWz78a/VPGG+qSWg4hSurm5VQc0zGvbk6LkEKJ8ru
YX0FNal8oat7hw5uKCGW+tyB527z6y2oBLGWqm7YbEA4kgwaQWmrIgmGJBRvYE2o
YoJpFBvgo21/NNLwx+9HlsdYr3QEB2cuKnT5bmgeXWN2LUd/yuIPbY2NMH26Ay7d
8yjGJCBv2C/av9h+60yU/TidoCPRLcWFCNrVs3zm7o2dKITDIP4QHwVsNem10LlP
4dL3BtKqI551mkP63uIVC0eGCkH02yJhLVzCmJqFJ2XfFRtkomI6xaKkQPF1tkkS
lnhR1k/IF05+uwDz6lHTy4D7FGYWiq6tT/6p35OpDys4OUL1SWFFtPHZkeaXBMhZ
KN6IKmPaedVViEphlWmIulaC1REqvuPYyMJSUQ//KzBEmNC9GhOCd+hJ5mQM7qui
ZwZCIKIf+wkmhVg1bkSjGOvB3F29URHeSKbOmxanDS/eIoFgapM5JuK4yP/WKNpO
bnIS4/62LP4OCJrb9tfAvhcYjJFTHzyz84AGJCUbB+U9VqhLsDMEqSxeQb80SmDi
jiBQbWc8J8QZH5w5B8ES80pvPKdeyuezCkOVZk1PJkkP3ei0nMLHecX8DQGjiUMi
wl69jOYGjyzUWFz3qkd4EbYBSPuRXY+pn3HXfll0iqDx5ysNT45ZZ7CmfBD+LbfN
PJ3zodS8Lckv8kE4MVAzAHn10XiI92y1MsjrP70w4INRanarOgZC3WNF/T14ndiH
mVTtAdXVBGwK9UyEMCYFNFoj5/5fk0ixhtZTX/a2YKu/lqwxsluiYTsi+EAa4Iy7
5Q2eUmIIEil+hJFMufUNThLAGKH/gP+w5WD0hnC/c9E1FGZCMJjprUFjkJK4FxlL
xrCcIotiB/x8DQOhFt4Xx0FbI6tyW9EQoEcJVdGNOMJhl5TtCUgAdvfCpyKz+aYy
TBFyy6Ca7UTtg5n63FNy4XaO+D8Bruw8rO8QRSL8tzUSTE1Ts+RsOUNhXEoK3NHX
cH4MzG0vbHDul8iBReIZWT2NyL7/DmPCHsLDhUdY6O3B8axwGWPn6fmyanxouEl+
U+DBLRQvjZuys5HGROUZy5Q/K3fBr22E1iOwtRaGuTUkBZCq3r6BoO+sgBC1Cj3S
9QUGto7GiO5BZvs538gTCZKwQj48Smds1+t0ewuHH+bkCDoEYttMnSenx9dC0gIx
ZR2bPCkO5NYxsmTMxGtSYWdl777AppyJARr1TMz+YlnrO2FW0vegVEHEW9p4jAOi
yHIv2eSJ84wXxTCAaheAQ29xSnrjyD0cfg8e+po1dmT2fDYcuCQtEzqe27x9aLVH
cRF+RgjR+ax85bn2tVVa+tLNeXrdzE5gwtu9X8N1Sey4l9lrAto9WNLjBuiSo8DV
OuQc0VIPaiTOB34QmHq1EF1TngVQ7phDELVsyvRjrn7afoOHVgPXY0l5GcG8c5xB
AH+7ST9Zvn+G09XN0L4/UYodYUxDXnjK8bwC6EOOFhjQSsh2JrWc/gx06sIR9cx4
AAAZsjGNXnbrJX6mlX/b8cqZYvp7Mj9IfvmjLass0U9GOe7kKsY08DcsLAkZcGhJ
a3BXP3FfpcWerrNdLuc/P+PWjfCPFCPgEDNu/00ua+sIRIQHZXbSHA58mdljK/gI
hGFfvxJ7PiIGKCoLDZRUzdualMYS41jEWhlH1S5FFcjzcE6pyM5wYf88RkcQ8qjF
GGEhDbjT+nBii7teitde/EdagPiCvqrcHCNy8IUeFeHKPkY+Re8xF1y2FoPlBU7L
mQaKAyaYMe3VfQZPsKuinzCUwDRFR2NEHSC5d1XZOXGm4AEd3epnR3qEIThV/CB1
b9Dq35z+lJWqvAS0ow0qUs6WVXooD3BkhoHizf90MGRagylQ+rynF2xBFAlu8nUy
yjkfiHv2YvQ+9aD8l7xn5IuXKAU4IaheHTq3SE5O0ltNF1/MYyNijXeL68ZweLBj
yPaAvvA3M4iLrMoRwaBW4/uUe2MM30ElRO9LPwam9rPjxi7HQncgyxmOMBdCC1/2
JMdLMMFLlJkqVMQdFrfy+BgwT49DJU03eeBDUrByDV449royn3P1k6zwQQ1e5rsR
WK+ir/6EBAi/tOwsQwnIZ6jFS8LAkk2GaoFz2pQhTPHcMulRPHNv6b4Uy6XSGFTX
06BmCpCJfQxT8UI67mUKGnFbv0L+mbEDrUEGFmmCFQ2GnvLnzOj/IvC87v0S+CKm
CP0cUHjG/DRTpQcxj8ayHgIgCEXyKFCLWBeipo5iMhg2pQJax/Bo/gvwEYyVc9ir
wDwGj1Ty2NyB46roR8Fe7tVGDr5XKMtgZUk8rxeZy4Y7AlQ/A9/yp2lZnryWX7K6
eR6S7iuAxwcJsKYwjt/8lufND+OCW26lj0AKWpSDVr+3XrBhfYIWDmp4Jak/bno6
IO0xYEFkr9PVbvNMc9BoAgsiwQ2fxJoxsjr1KMJ8JRvJzD53Gzf799CU6RslOc/9
A16XES0WBZa+EO/9foyorS6YR+Rt/tMdN9dDP1bx1hhyCUct0tIt2CP9NvVBiAGf
J8kOrjJzy8apv4qCpUoYVL/j6bMDd2GtOo7Kxycf2TlXp16LLdrLA9X8j/rBxH9D
Sfi48NOCgVrs1fR4lMZcT6PoTXwT1pnVgoo+iUbZxVeeIwStRmxY79jmUQLikEbP
quPdczyg6h8fDe3vmYIY21OfrM8mtic/KaGxGPakydQQy5JsoDK6PGrm59aSGN5a
GCM3Gv3TtX4OYm7F9MnvK0fKjzjmO+E48+NrWQ2uJW7jrzCwdN1Cv+wn4pF3O4X+
cUVmiWAu8hhH0ZCx8t7y4AUZArBLJPA87NqRqG6GvR2CE1eD520zP4Vm7u7oLD2Z
Xcbn6vhR1yUnDg87cuM766KLwDNKRWcyZSNmwy9mO5W6y9TxFGCo+TW4iemsh3xc
eQM6tQHjg88d+eXupgUUPborCl5wKNtGSG8k6pgfQ2o0gaRRZsTfV785yDpQLedU
QRQYoRirjL/DaCmouqxbP6l5KfkWB8nN30WL2+AJzIM4wP1omLn5ZswBx+fofSHz
1+9HA8OIF0kExktr1ztkPW0EwNlTc6HzQagTm237wtR4cXK/aui/30mG+hjq+696
Cx9tpnAU3pdWdWTXj1zPW0tw+pILyc0ChuifO7e/sjfl79RoUJkDtIuNF+8Apn3K
AZA/6eYUUxhsZBG+Dfsrv0GsbZcAgfxuFnkqqSSAjWMe/AUTvYpHTB4avXOp9ti1
vGFA3uyUd3roWIJKiBn3kZxhqYLsJNo6JH2lOIJynS9ukSfYO08vYtsi5UliURfq
8OxgWyy0n0xBpOdIp84e3eWSxDty7kkfVnJIXluZQiQo5smTamHMSMSU+SrdXxKd
q0DVQ0lqa9clYW5r5QmUk6EpWIMoU5IK+n4HKyb7fa6hSSOeVkbWO0d4+zvGnSlx
LM7vhiFsAlCfAslAzTi97Kv9cNfjtsRVpvLQRMFLrniNOrj2qN3grZjLVFr6Q/nk
Kv5gPrurzvg1VWWB+MQFWoVMNvPV4GntKxpvDmgod/xus9tQLFTRP/nfvmgy5QBR
uaXaO+nP6CrGia4bXcmCDPvZDoxArmyaKYEWH5cpjbDIpAc4MhwnPjD2XCDp8d+h
s8xvnWRuO8a3FwhyjtDV9/gWukesQXEGZL6lFYWlC2kleeMFm3eGoQDDDPyaOU3b
Ox6mIrIgCQGY1dQfKUimaRRc5QzPFF3xP5jpH4m2Dr7g+yS2yrtdmCGq01Jf4VLn
3hZmGTKu2/R7n2h4v2jNUySr9Gjua1OotJ6vy5S0mhmL2N+/bm1806yhLi98Fi2L
X/3ygRp/qn1sDf+QX6qSUSOa3aRpp9u5eyLZt2kchm6s9M7RyecbKugMHuqGVwNq
oqxnwqUj3Qjo2gbjt8stwe/TXNz/EV6dDLNSJhEtbrSnp+hQtgDCB8uqYtaA+7K8
sHGlJzQzQdrN+IwoLLDzn1j8+MP5jkCRUsd2D8YWB9MFvDIGoMEQw2/Z3Dtn5/aP
0CS4St9VwQoT0I0kQNCfMVzkHB+toQzcIUU44r9ktEgNunI/q3wTlmkoRCBfRE8C
tWnvrHtqNmjiCxOh3qqsUcqTikewuc4OIxPJIXvlXFA=
`pragma protect end_protected
