��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��eڴ��XD/=���~U=����.eKUl )�xE�>uE�}�:�"�J=t-���=:X0?%r�H���3��x5@|���	�HF��L<�l�17&��-��d�g�GD|u��V]���j68�[l�	����z��Mj=��O�� �^�.`���=�B ���뢹�mM��?�vAFu�5�l�S\(]���P�+~����Ѹ��r�J'���d��Ӆ�I�ԁ"[���6B�}\��y%�]^D��.��i����x�x�V1'����˕�tJ_���)>���g߻
ItO�F�RE����?�6+Zx��(�O�+))ʎ�e����F}�����̊���a��2��`f�r�@��nT�@F���'��d%�)�`q��q���W����!���֮�PP5<���%�V���&Q4��M������<u�� Zyg��?n��u�n9K8�ԅ[x�K�� $��k��\�䲧���Q�,5�(iW��&��9�rv�#�u����Cn���ts�!u|I��΋�0,�r�*nڕ�e�X0�|��,�]�bw�_(�{Z�P����0*rpi�EBY,#����
4��nB)@l�ۓ���{ٟ�Y灂��7���TB,Y��wɠ_C4�leO��3�Zp�_0��4<D��z}l��u㸒��M0��A�z}w,����ך�t!��#��m��i�cz�v� 6ӕ	�'R�=���p���Bx��6�%Z�idT�eÊŧ�F@���Iep|<�E<��ؼ����m��͇]����+]-O���m���td���]�� �t��
��L\��2�냈v�v�{.oD:��n�2�O�q�T�8'~���a��%Y�+���.,H�Wc#C�b$7 z��3J�,��A�Q[������2���b��Dm�;tT|����,\p���~??����"��!w�V?lP�)
�1T�0�Y��؄��7Uxk�c`U�iO�����H
���N���� �<�������J�|��� δ@K줊ʑ�SNr1���yc�1[��zE�4�7q"����T�~*������@���)v���v�yaA9�L�F�TYMˆ�׏DǤW/����\�(�� ]5����kۧ�j0�GV��֞�)�ɇ��߳%L��������$H�N��Ě+��?'��a\$R��<��Y��]�-"���W_�7��Å����V����J������w�H/�Ef�caƔ���'Bn,����6�S����Ӑy>y=��{���MMr0��r�e�ut^y}��j��P��u���U*Hu�C����O(b�+M�Y\)�k�]�9h}�/���G
o�?�A��C�1�R�!+Ƹ�IB�ȹ�F��)����
�[/��1��|\7����Y�l?�w��]ъvY_�"�+�rg��P�f�i��M�3Eky ��`j�ߛb ��G�x��t2�!��EBu<��9�{�������Ql����L?UE?[��,x��V���5n�7mQ�
��l�7G�,�75�>Qd��*G ���w�A���� ��e{��N�l0�Ò��������$MPǓ*lA�v�d�v9�*˜G�6N{�F���$}p�8WP�~��z�s����M��DY�9KxS}�`�p��p�Lf��.�m�{
C�/$gP�E�¤1�Y����"b��/I#��b�y9ScN��+c|٭'#i���)s!�f��dOt�P�a��ᇈ����X�fRe0��*���i?�$ ����7���3jX�hp
)�և�*l���ָ�����:G/9�pu�=�o}� �ؐ���L����-���HX����Fqd~��y�{���m�2j�������\s��@��4��e���m�����1�?�V�ܣTQ0aKfe�� �u�Aq��y�d8r&8��љ�Na�s��]���LFuZ��r�r�1bh�ѽL_�^t�Gp�,Dh�V���X*�ŗ��Rʹ�l>��
 �,��M�n������q�#�C���w0!�6j��T�o��2i
dR=m�H|t�,,��L�809g�#��Ed�e�E�NH�-�CY}�犬_0����;�E��3^��E˂��C.�I�Ȯ�@=����IH���}����F��M�SA+k�]v��[e;꺅���F�����8�4��-Sb'h������V�d�iU�աR)�8uĆ�E�'�O"7kM��F�H�s�|��Gq��I��gj��tNv;�<f��y--�LN�inf0;���>m������fUvV �@qGוֹQ#���(@ �H[�TEغ��v����N��|�����9	��*L���N���^���5DCE�`��ݨ�(+/�}�:�n]�?��5�S�=�Vc����n6�Z���� e� ��0_��O�
2eX�d��=x���L�I��Νu�������[�5M��M�PyVy�{p�����&z=�܉���`mHI˨�$n�W.78�`�ࢺ�ONVx�4¹���!�G�����c�D��o���7�X��F��:�xE��<Zu��ˑ�l��V�g��s�
/.�l<+�	�֎����yL��4=����TD�S�{ƒ����dY���rP�#�] ��es慄��^\�������SSs�A�����淘���K��s{�#j�TZC	#��tonϬ[��$|<�m�|*���4�G��D̆��Qk�*t�`-�P��q+A��
�믯��{'fM�����d �*]��|��#���O!��w�C�c�rL�Xm�ܷV7����3����`�5c�=E߂�4�R�G&~��DC��K���
U�{�p'C?��������L<�S��ig?;�;�c-xgH����t��ll���Oe7X�i�O\�]��r �R���nKt�i��L�y
�b:���G�	p�Ԇ@��Y�����&��U�SGrLǵj�i0�E�oG�����@����w�ONh��h#-f�����=��y���_GHE!~7��d��$���E���-%�WL���j3�4o\TlE�/g��k���vh�`;�'���X�od�M�0	��!$�Ա� �]�i)�:&9��#}�:���=L�X�-���Lq,�E�z;�=�;����Wߧ�9���f�!l;���t��F��v�p�m�����?7�
\HoˋtM�P*��
�3���xZ�|���!PeR��ssK����u���6fd�"���|���̻<������;��?M��o�������R[���s��:?ʓ��;�w|_���(E�9���w n�+��!t��`/��5/A?=�<i���}��:�k�W�#p���!��_�� ����r|�=P$\�����R5w˄�Qҽ��ElO���l]�a�¡���6��8��͖$��؅g¦4�vn$��@y�O�/4�0��)��;��-�t�M����R6����hl=N��k��]�ʄ��*���)�T�Vk��B����1G��r]������	u�ฏ�H�H<��U�]�\�Zy�X�������-������:7�7�e�P�����,�0�gX�<�I�����~<א�TH�w��B��e>�hN��6B��)��3�����QRޏ�w�4�e1{�Κ�!a�m��������Q"V�����gJb�$���^��W�H��U�3ZO($$,A���n��J�"eRX���ɹ�_T�K���f��	W
j#�n�9�+{ �.����}�����k1���7��P�i�1y%�*�����/[��BW���ɯ� �;P�'	�RӞ�x3'�C��̲�S>�]���b\ƑQ�-9J�P&>��+�����.��ރ�D��^���ă�R�e�$7�^�������#������Y1~(_T+J�w^4�hG���Ҷ9x��)��kbyK��j�b�Q�:�%�*%��(��EV&v�������=���>��#p#HЫ���I�]fu,���	z�4g�?f����J�$]\$J�P�L��3l�\�)d�w�#ï'�5��7��}Y�t[��|�M�������X]|s�3����Y	������)����/��}��ϱ����P<e���'Y�Ҷ	�Y�����hlw�y��t��Bju=�^�K�z�Ņo�=t%�L
8�:y坵�p��=Y���x���'[H��H����Q�hM����uK~w��9ٴ���/�J��f����C8�� �O�Ac5��ET0=v�^�� D`vM͢�k
v���u�8�o[�_���ċEl��RSE�s�흄���]3x-ԙ�(HY��O�5\��6_��)V�Vh���&"���U�@�lr�d^%�SQ�e�Xi<^�ɸ��f}���j�pF5XyB74k�f DoϏ�)�s������^�3)N��c�e�����m����ZȌʺ�nL��I�n�[�SE��M��<�ǐ3��.kֺG���\��M˙�0,�Ue��M���r�j�x*FϨ��~uk��G��4�b乮�=��L���ۅٚ��
���pCʲ����__pX̒�l*���5B췯r=W�HP�Ҽ��m�0B/
��Uؾ=�}z�CC\ﻶ�0I�u�)0��T��'Ň�OI�!.:L������.bkO�)��sW��\�+НOMb�x%���+n�/Q���˩��a�e=���s�oZ����'=���lR+Ff.eW2��<f'�=�V�/�t0f��d�0z�Z>+�m>�3GǠw�ј�� x�x����߁(ʵ)k!x�6��5��`�I�{���/�S(y�~'���@ͤ7_Pa�DJf3���v�0���nX�!;m��;	*w�BKj���C��W�Q~̟��H-��G�y��)�%ɖ	�GB�����Y�}y|�uN6{'���ZrT�I�O���>��.i�Ptc-����� �"vfaIO���l�����!��T}����~�Aia5Fde�Atػʇ��uw�4�k�1�L��nT�a��lK�<�d^h�*��B��ũ+��ո�|���'��.q�%'t�ang��
\�OX^8���,����o��?֟v��|�$iO=>y"̰"l$)�+y��9��׺�=FO&�+�4@V	7L�t�.ѳ�����m�Z�Kvm�
(�Ntlu~�!G��C3�!٭��hH��Kb?� KlB_Q�4�ud,�?�B&]������,,UPTۑ��rov즴�G.fMr_J!���9����D��X��K�ɰ�)־���Zܮ
�FF{�������T:�ް�r�bwq}5M��@��>C�'!�F=���6���M��x��*�Yy%/7]X�vC
ܻ'�I.��Q{C�&��]�F��=N�S��(`�U+z	�Ԥ[m�ma�&�f�o'�pK���6<�H'E�:&'���dlńd�K�z�0(��N�3��:�R�YN"�w�*ɑ�t��3y8A"Ix��-���y'��$Gm`J�r�)t��-v���vC�&P#_n����� ��óKO&f��_@r�=7|d�iI�����aԒ(&�m��/�{a��!��x?&Ҳ��Hqi��ר��#�2�U���x|D���Bzp�"���54w���#�N�η~^���b�E����{sI[U�N����w��p�S6���׆��鏻+�t��?<���IߵzG|�P�=p�oB�K�H�e�j�����(�Ni��8'.�M��Z}0���X���?M���@��3�t�4�'xS�K������ѳ��KZ&z)OU��N��_bV�ϰ�H
 �fѿ��{\�;�i�(��1]��&���V�A�n�ƢJ��z�Ɓ������������n��\;k�ϡ��\�Z	>ݺ��#tꍵY�'�
SG�	!`�}����ZE�q��p�t�\Um�[������Y�176v����l���� ����L�ֳ��z�/�*�^�݂(����i�nY9�@���cgu��.֧&����HS̝�F�V��wYV���O4E]hN�A���E�8�i����R��3u�\ٌK�p"�J�&�=��A��,� .T�L��4= �7H��q6� �˨�/���r/���X�3��&0`�k!h� ���{"O�����y�_�V9n4\�}�r;&��2�)Y�e��!����Q��ֽ�]���q���$	+c�'�Kҋ�$�m����]ii!��'�5�^wnP�㼍ȼ蟾5_��hQ=����/�ؕ0�d�\����E�u�m�[Ɛ��0`*�G�2]�uɈ&�|�yT��,4Ӊf �LU���W2t��ׂ���<�=��F��?��|V�@?L��֟��(L5C�7�zm�8X���Le|��$?R�D:��VK�,7o��ں���?t��s����Z8��v~���4 H���<-��2�>ҵ�~�j��������rPw� ���Ҁ[��ss�3�I�������v����(��h��b.��9�+���ls"��>9R�t}�uF�?V�U$I�+�cFB�I�zڊ�� �9�e���*��cp�ԇ��,pV�]��@7�8:�m�C?v���j�[#R���n�����i������E��UvMߢ�M�2
��\b�� �Rwġ��[��8�A�)���K��.�:�(4�y`�#H&���Jz��h��u��*��]�>�1���D߶�QC�0�8(TS_��2L��W�R�U�N�����#�Fڳ x0�5���gu[�2[�wa����*�F@r����roG�U^BT,*kn�P�����G��ຠ�����8��ů�9�e�K�����жB��R�#S��,�cw�篱ߣm�Ot�ש���={�Z�q$�q�Г!;�6�W��v�bÆ���8�
�]�c��|��=*��$F��dq�·�R� ���8�I�?��)��!&Z�͙#!ǁi�+ӧ_}Ay~Y�f�dw�l��%�&�!sҝR�K���GȺ��S7\��'/ �M������{ �xK#�P��V��7�0J��2��c��2m�]iF��^2�b_GT�@����)�=0Ӡ����J�9������ NM�k�0eਛ��1I�ޕT���q�
/^�Q~r��B�\���iߠ���O���pTB<>��� ��R^Gg����� �W냣����7�����;}M6,����� M�8�� nA����N�Q�vf��F$2�'�菧�\ND$-ioj8�n#�� �t��k�����Ԙ~Ԁm����8(�L +HQ8+�����}�<��:-�#+C{�E��=\��z�M3Y�XN��Zڸ�&Jo�,W�����:����%Ol��2�ӣ�u�Oڽ�>�$$FC^~�ɇ�郒%���������=q2��:`KQ����kH�<���(6	Ŵ�ML��D�l����zLN�{E���+�8flQ� �3�7&~LX��;פM���̦�2���}yn2[z��@�I�t]E�8o�+'z{w�cD�]&2�9���-��;Q SOW?! xIǵɯ��n#��9:H�NJ�=�� �����F�:[!@ݥ{R���umW���g��pCA��ym�%/��E�#��	�1�<�+��= ��U
@4H3���$0�cX �^�2����>2�Qe?7����?�	�Q���&AVw�2�Y�4L�����������br$U�m��a��5?bE�>D�2���,��0������S� �w�(�dZ�d���d�������|�Xc�����*��K��3۱\�"��s\zB+.�����ڴ�`+K��y����
�SVh�g�i�~BZ�a����4��� nIM��e��-�~P�y҅B)�� F!���Z�ʾM���[6��6�-~��HbhW�2�;����rR8�+9,~��ӌ,��1j���]���~a��<s��p�����2��bЍ�m�z����.�ݻ�/I?�q��V����H	XƉg�u(��p�}�G�:vr�9���U,4E�Ah��;[�ZGnoi+x>a�i���TԵ��yV߁�q1�7���q{>�'zƘ���D�pO���!�6�g�$ۅs�P�����\Q���$&�ڷ ��7�k��^�1,*��9&?���!�L��?sZ�-�q��wd�b�=�����cM���1e��]j>����+Jo��<��(������?�+���!c��'�0b��9k@���l��_XRn��gr�C�A�1������^���j�{5��ڞm�;������$*�i/�Q�w��f+����.�+�������P�vqxofX�b��Nc�U^�'�R.R�&��ZwP������q��afFS���9o��?^&c�Yp�;4T+g��d�EL�0�J�5L�Fd%��^N�>^ ��t�{+��v�Oa�ԞZ�i�7or��x�\��ovƻ����X�|4�է�������D+3w΃����y������`܏v�o��4w)Gl�2Ք�>��A���-ۀ��� mM�6�Ůh }}���T��C-Y��g#�W{��,��c,r8���.)z�>r"��O��E������i�����̰��uv��U�N'
<ڡ�PX��ˏi4C�|3��V�2D_��B�����b�쥽�D҃��_��A��wG�O�ۼAk�㊒����#7�W���t� g[�6L9�# pL�U�Ucaw�K+̫tA�zƜ�oɱK
f����O�fC�v���оA����|8ĵ+yo=ี8��S���n��g��	
��N�V�	l��VH�	d� �>���-,�~��e�Z�g;�T���`�,Z5*>e���h5��V}����]pȠ��ZW�xę�,E��w��є�c��ղ��"��l̈wu�X-��9�V���/`d�${K����.�naC�.5BL�S�/�\�3����f�j}b���0�;��S)uEA:P�[[_1�;'��~iQǭ�@�U���H�3ڏ�n�`k��窒�LB����!>!�rG �jP�W*��&���`S�EfSQ� ?�5�;���r���;W��؇|e��<vA恇���Z�	����+]ń�CCv�sU8����jc����gMR�g`Y�����E�N���T@��𤞁���r��)���)�{��������.b3����6̞�8�;��&�/v�I�#��m9�z���hv#�Q֙: M@���ˊ�x����H�8سc�h��߰BZ��A�ggr�_^8uv5%�tL��(�<c��e���e�Ƴ�F/^梓��t��/,�������i�Ғ�����%>�\�`yH_�S�u��;�Q��z��MJ��ap��%") �Ld���a�m���`���vN������'����?0�.6��?���+��)�{��p=�l<|5b�w(�zD�#u�	�kW����P���_��R]jINe1n��rG�B?����Lnja����������~Ɣ\���8�b���0&��[�p��5*h�F���f���/z֕c\�J%O�DKX�7��[s�ӹ��+K��H���}-U�ƺ���y��8��䂯��Ai>�!]C~��9��}�G�+�1��2B�e6z�X��8���E�X��ʆ�?��h��_��b����mU�T���k��c���т�pPr�p»B��)˲�Cs�iw� �����JZu乙K���;ј���-)#!�Q�0�a�j�^Ԋ���g�q�i���pr,���(�E8r���j%8QЏ+�0�ɦ��=�r��r����ɤZ���ݺ����#���)$�ƙ�$irZHF�m� �	J�a)�@���#�;3��@����2�H�m54�!�ju|QsNV�L��D3?�b@0��aL�nL�PF�-x�eҠc%�[D���R�����x\@Q�p�:-�¡���;� �)n��$/�P��c&��p,�9(��Q��m��V�G�!Hh��R�ͮ��rSí)�2��Θ�v6>��s��Z����Cq[_-[i��f]�Y�i<�S�:L9���|�s�>Xn�0��#�q�~���B��nQ90}�����hV�c��ر�,��ٖ0lV�5�_N턫��P՘1j_����O��}�-�V��#<�e���3����G��v(5���{Upy�&}�[qj
B@_}�9ޟ��8�z
��F$'-�M��-���l�^h�7w��n���ЉC�K����l��7�ɺ��۫S0۲����#*l������੩uuk��#>�%P����*�"��]��C\�ӭ��R] ;�t��˖�{ ���m�T�����L���eh �,32g��E�V����&����g�°��(n����M(Yz�T������Ɓ~l_�����н�Z�!	*C�� ]!wL]�z�,��_�c��]G�����XV ��`}��9X��en���#4?H/.sc����^���a�B��D1K�_��,F��c�ܦgێ������������>ud�����6�G��㶖�>��6=���Ͳ�mk�MD`�Q}���A ���9:+@ᾄk�\%����1��0��s�b%� ��GTu�!�D�c܋/2%zVDMu$E[�
-�M�:�_^w���<�p����q��y�=Ⱦ��޵��-a�ѳo����ޤ���;?y�&0��P�^�pk�5*�t�\a�i�3N�� p�A`�H^��7g: I��Z�[c������\�TD�LK��B����VeҠ��.�d�/�������D0I���`�e���&��>�"�\[܈�s-���h���g�Q=.m�����P�������1��dI��F��T�)���2�u>�sa�Ey���eo73�b�6�� 5'��7�]�HlE��Ԧ/4E���ğ�:;�n׬{����&��=��%6,�4H��5�Ftx���Oh�� �p�G�Da����[�u������&���$��+�_��^�J�g�Q�q�]mY�]�	�(��rexwg��2 `,�V����<�Tg ���C�굺Ԍ��A�; K(�ҴKC�.OӢܠ�W�*�?����a�pƧe�ؒT� �:6`�K0�{4g�.����	l��B
XH�k�z�n�֥�G;�6���H����6���P���V�X��������B�F ��&u��b^.3��������v\g�f��q�6ar	<���B��<T� Er��S��_��P�j
zX���"B��J�C��Sp��̃⥍հ2�1i2����ujm�ŋ<�2�s̗M�:-ȁ!��mq��D�ݑ�ѿ��@����抽�bx��?��i�EeW�\β�Q�;3�X�D�ܐ��/gDJ������J9f�65[���eL�9FU`7T
 %���֊��0�I�oҧ��wV���7ö�ÖN�3�%�LR&�M�Nh1F�nP�|�i;�?��u4�����@�F�y_���`aw6 &�*C5���,��oכd����o�t;�'��x$?tUŸ���<z#,=86fK��(L��ߓ �!q^q�<�a1��������n�8�p�.�b�s�5n����#O�
_fp_�'Ջ>�pTU���p��󛪘�ц��1xd��.v��������*f�Q������^gY�F�X�}5��C'W$�z4��w������,���f�~�ʒ�3Q'��;���@M;ԁx���7���7�86��#���a]X�����P��2UM���:/R��g��?��r��z�$�9��q	q9P`��(�}A�X�*�lI��*��z{j��sNlO�L.͵P��Zr�2��3N��[Xs/c,>-釗��g6���G�RAiĎ�PK�P{�iG�Y�k�O�E�8���DSk��%�:b���s'=����J�����������[&��k��wsj%wt+����W1�&���LB&�"$0B�:�K�����B	!�\�҉��`9����M�o�V�YJ��`㪍�yi���V==1L���&G��@��� ͬ�}0I-�{�"C�_F�е`hBv� -%D{��vF���RY��ت�zFU���|G+�i�u�ۿ��0q��@������1q� �].�QR�l#2�������v�#�5]pfrw�o���+j�&1-�6�kDdgv ��b{�&�tp��`�7E���9��xr5�f-�G�zL��'n� �Y���zV�<���s㥸7����5��rN����� sV��yϱl7�$ZB�t�~�UM����T��>�楄.�š�{�hV���� �6�BH+ᬦD���n�G����CHl����3�r��ia��<����񛿳�g������;6/<�~�)a~d!�٨�p*v�ޱF;��*g�F�/��i%���Ď}��qQ>����i�ùR���zg���6�}��s��3�4fZZ`�2�eaBe-��M$̓���G��~~:�w�PN)���I�������'8�:?�p4#_K�F�]*61f\m�y�`)��lS�Yv;S*m�b��~m��� �EZT�ͭ������	$[��W[4}v慛��O�lڞ�RW��>����V�����"��n_��c�t�K=3�f�D�U5���/�N���ո��)����*��ɜ;ܚ6*F����˘��)����0�S�Kљ.h�1%��/<<lf�w+��_hĞ�0Y�}�	���Y�X���<�,�� ��o"N��~�{�i�l��b�DqdX��:�l���Gf`�s�!�8�n�����+����ޜ�C�xZ9��C��Ԡ�!���K�*-t{����ӥ
UA�]^�w�(33j�1qP/����=�uV�ъ P�h2�T��Aے���k�d��k�m�P\�ܔ�ȱ�^��3����n���$�?��Q����.����2����x�t9��O��m:��H?dO���s�[#~T�M��"E�-#��"ͭ�4�,��Ǵ8x�1eXA/i�(��d^ ��n'_�D�2?&�C�%�{�c96�����sȄ<5���/"f��_��
^�N�H%��.m���0b���9vn'��,UA�4ȃ�ɻ�^����&���=��ĳ�SZ%{�Iڻ�$U��&aF���I��8��͙d�ПX�q��âR�͔?R��s4%G@��|#��G�;p�������Y��*٣��=p0:�\���&I������������!���9ZM ��v���e.a~cJ�
.�B(fJI1苚B�ϕw�̍����4����q���?v�*�S�����L�G����I]����<U�4�Hu�d�n�!Z�LC �#%�d6B�)����Wt�xS��M��c. �?�F@h��xɦ�iq�t�l�,?��h�I��^K�5)f]����{�Ff�S7�����C��R���uf��C����m#.����_Vx�߽Vt����`�#�Q(�^ uZ��د��]ȁ��S���U�@�k���9РCl1v�B��[�F�+�ӡ��Ų;RD.�S��	ãe�	6PJ�S��A%(5d2O(Z"~	���k�~�P^�g�SN���"���.��Y��5�����׳�Ӌo+h$�vD����i��'��`��p%0>�3y�E裮��?\��׳qT��l��{�Q5z��c� �3������3!����c:�w��c<��5��^�ED�L�*��k �*簤���������L$X\�
���j��1�~����𡄳�EG��S�~��":_�H�a5!=y���A'8� z����ts���N$3��VU�Ī�]��F�KqV��cuۓ��]�PDb��h�U3����)?��4:�pqFB6�H	_;��/��r�c'�Χ�fۗ����K�j�h���!�m��p$M3� 	�@%fz������w�w��"�T�{w�4����D�4�n��}�`���ׁA�T%&��ߌCme�Mȫp������c��b-f�s��bCe��,�][��S<�R��]��Es�E7�ck|����l̢j*#���u�z�s8��\}�A�mC"T�nȪ�"d�q>�����'�[��>]4k�nqa��O�;j�����̐S�a�~'ћ�X�2��r
=�]��-+���=D�X�f�u �q���1�9BWg�4�e�/!%�>]?���+a@� �b�����l�M~����%���~��>�C�u���.W�jK�} ���F�U��-l��g&�L�P�#�35��9�\vx���h�6�]/Ƌ��H9�e_�%$���|UG���Ƒs�G�����>�<�!���*-��T�n��U�ߓ���m����"%���sMv�~��U���6�\Q��#��'5�l,�ܖa�����3H���3��
�����6jwR[{�w?ZbYH-QU�eX�n3_�䓍`��.��=���T��U�FR�}_��E�E�Fz�fi�׵\�[P�Yp�I9��YH�~N�!G��;���;��E7�g��ӗ3�G����������w���Lq�P���YJ�׼̞{�B�V��=��]�4~�R$�m$Oj Q��MK