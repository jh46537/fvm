��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��秤��sy�/�F�5�
ޡ-�ǅ���$�k�	���M��	SK]Y�hfq�Ff���b�6��ef�Tǳ���.��L�^zu�a���A���3Q<Vi����j����pO��p",gD�p8���<��ؒV�D*+pY���S���`*�4�ozjվ���v��$q��Bf#�z�קt&� �Uk�Ay��0�:��&�Qo�ޫ]��^��n\+M�Y�#��t�I��<���-�ײA�ʭ�C��mYw5ر�9D�h�q�����]eՁ/�c
E��&3k���zB���
�~��R�;y`P3N%�l��P?��А���ow��K����Z��lNN� j��֕U2�ゕ~��̲�p4�?���+ߟAs�Z+U�̶;������@k��-���b�G7�B�
 `i�WxAi�P���������1���P�ΐm�x�:��U)��8<�Rf����D�?���b��5�:���bg��8t�͡#�d�����;�S�ܠ���d��K-��:����LL�:k�@@�?M�j;U;�쓽��۵�,�F�7�9��7(��Y�ɵ�4�9W6H�����S�Dɀ�-��G3C��E���=r�٥�~��0r0��q���괮ۆ{o��_���p?o���ȈX^�>�<�o������9;��>bb�G`)h.Ǽ�]2Nh�f���o-�69Dɲ,|�Pn�n��:����c�
"�$S￳|��4շ��cJ�����x����@�&�|�GUN*��+iE��4S�w )�B6H��dl����N���_�� ��s��@�S'`/��tD�9�8�ⱌؓ=\m�Ah�3�8fx�UyA]5��U\`й�-��]dE�]�ŵ��������o�'6�0�W �VU�*�Y��4�\x���H&&�Z���lB�p]-��!�����/�.�6u"�d|�� ����Ȁ�w�}������Z[�h�u��1���͸9~@=M�t�MW��`RС��P��q+�]��.����$��<0#�?��M�;-樬�G>g�Q,��}���}o��ZB�!��~��ӟ@��]7�$ڍ�⓯�<q��� �	��6�9�G8��t�RX�/3��jgա�7�~�so��4mW�UW	
�Hi�b��t�dv�^g�Ļ޸J���x���;��*�t-i�8�{�/2���ǵ5����=G�C�@k�����[�̲��W��ۑx�&�P���
x�17<�&t���:qUY���E�V��pp�)�U���`/#�j�������]�Y����j�H��7�0�2�|���!�