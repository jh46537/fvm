��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���C1��
��4��$�6vW��a��9a�#E���}�k��?�|_(W]�?���D���޷��!�h.�:�p@�A�ҹ��mJ���=��jf���Y�\k�
=��of��.�>���ݞ���χh�s��W?׼t��=��ѥ� +}�B�}�M�.3�y�]��2��@�0p�o��H���p7X)���.���t��!s3\.�H��w�U��>�c��CK��^Z���OXW5�!XU,�K���/���;���[��ɗ�t$/���4�#�|��0�P�� ��5�n�E7x���)A���o��/#���?	p$��YOe�	�B�́Խ�0���H(�P0U�����wkT�N�$��(��jU�M)1	����g�*����ݻ�U!1��{�&0�^�|��"��ݠ��Y͝=��`��U�޾l$h��=Ӊ�l&�/�0����L�;����=�j4lC\n�WJҎذ�QH��Y7O8��}A�k�~;hĢo\��!��3��=�D�lC$��8��5��1L��#�Y�4G�i��;8���J[�W[��.q�Qz2�nʼE�"|���dg�"��%���KDxΘ��q��H�N�׊3Gj#�9� >��|�ś�s
�@ĳ��w� q��l�:%(����k.u���6�|�Y%���3S��hz��bqO��nV�����*�z�>�|"���_o�6s��w\��&W2�I�oKR��?�G_T�?:������ߏ\`7
���8�n��	,���r�_�.�Pi*q
߇��mh��8`�0L����IO�־DST�P�2��~L��E�p���£?Q����iX9�{}/����zi�>��?���Y���~��ƌ�A��a�����Q�s�6я���j~�K�O�����E���P
�|H�چJȃ��}($/�b"˕����\�����6xj^�#mv�bKYx7�'	���7�0hz=�����ע ��/����Mĳ��!�:X������?8�b�ox��6��m�C��#�Dn��� #t��F��C-� (
���v���E�3���]Z�N��>����PdU������\~@f4!=�?p���e
=9�l���-%Y������O�1�B��b| �S��B��gLw��=�G�-�#Z�B.��p�
f���?/r���Q�um��s�^Bk��y�	�o��e�xmR�gl����xJ�����>xGVڻOD�r��
LG:��>���v��s���1��_�A�#��	N��OuCP�����|���_r���V��R���)qn9
v�9�`Ʌb��L��^�*�s�_|�p�\���w��#��S�[ƕ4֨�h
��ON�r�ҩW��\�7ޝ��d2�3�,����&O���+��s���zĎ� M=�fr,r���ló4�	#n�H�F���4lMds���(�K��B7MZ��-��C9����w��R�BH�� dc�~�1�oJ�L<g|c�x�/�;�Yl?�����ƙI?��E�5�cڳy��&1X����4��*����w�|9@t�ћ����Jܱ�U҉I�����@�<���L��������qb��*�=LJ�z�1y�/���:OF��ZS6Kih������Xd6#`X�wg ��Ӆߦ|�˩�k��<V�?�&�O�� �,��O'��X��{kn.<�qY���FB��:�m�̈́��?o�/���@�#[[�������&hB x�������1�*;VK�B�Ed���9<���3(��u�k�𻊡x��\�M��}�nu�q����m�����H���	�����T+]�n�Cn���-�0'�p_z��+��k�D��[���<B>����A���@8دw�m��=�qN��5��~�c9����p��Lk����E_^d�$�iq\þ�e$��\6�� ��Q�M�!����gmʖ��i�0�ٴ���/�-��1�Y@e+�OM��z
�(��B�O8���y��+�����2bJ'��[�v���&y>�Yʘ���Xџ�9��;@4�������öq(3б���(q;�G��h<OS��N�~#����Zub��-!��1��9B�͜'�׮�V�����8_q�➍��Ѓ�'�̫��J�{��!���Ϟa/-Pʖ�S$� dm"5a�͞�m7Ob��w���^���
�����6<����&���#0�M3�(=��%�C:�]��?|4DZ�P�ޜf��;)��~<�%{8W/0�{&�cf� {��UK�V�w�mҷ�
���ts5��j3ؒ�D�n7L���&Ȏ��G/��X.�r冓��i�{�����Ğ�h{��8id�@��j�tb�~z!W�;���#�}7I�,W�&_�,Ti��@:���K}�Ԕ��h}{1�_\8u��񨎳�IT�m�#��ͨ�6�ж ��7?-Ǆ7�<	[���$�D��/f���ރ�pv�$æ�2M�3?����J�Ԗm�&��Rc�`�B�Ox��:��%�+µR�CF���^�����_���w�oʶЩ�(����s\G[�1 'dl�؝�x2�"��T����o�2ރ���)��q�ۦ���8o��0��ϝt����^���~���`)��E�qFOY��:���m ��d>�'�����D�J�K�r�7̋��(��"U�gm-�0��|J/�]h�r�w-�컆�@Cx�(1d<٥.ѥ�����h�D-��jR��#�g�+�/�#l�.�?����@�THol�aPZ���@�ի�p�#5�,:3ݤmK����
��������r��=���°6P�ܱg^ȍ%^����Xx�ߤesw7g�k���:�Q�eK�� ���T%�`4H�カ�L-��
"�Iٷo2!q�?C�ٷ
y?[u︟����Z&���v9�!�mejr7C|�
5т�:<�����nF�F��j-��(�0����ʾ���,����i�A��L`���9I����w�������o�����#�y|� Q�ܽJ�U�:����7¶Ց�/��$���ڧCe��u����RݷE*��� ���k;T�W^��;�#��s��yuC�M�|���3|Z����[/��R��N��d�x�ek���Xҋ<�x�_����Y�15=��?�RP�4���P9�&� �A8j�%7�I�]�wo&��b�\�L��t��(�p#�7')���P\�5�[߰����}�htB��$mS6�Ӵ�p�QxM�顨��(���#0p�\֘$��~ �5��,������uKGuH��uԣ��~��g-��Wɚ���ғ����������j��OJ6�Xjݑy�S�	�oE7��NQ^9Ň��RPf� �~T�iZs�cM�&M�D:�[z4�n��mr|��Z	��)'4ڧ��b�,I̠��R?���0Et�����8<76b�������[� �z�VA���\b���q��\65o	��_(��8�2����kz�m�F���"X�ƽc�k�9��~������ȵ����"�&S��wppsxR�<�>�&��ET����F�?GjoT'|<(��/����j�mSC��?�6O�'����f盧b���no}�I�K�:G�$#��8I\a.�\Qsȟ:z mA��vWr���ZǕ1%����	��F[+��_��eSud7��: ;�=�2�ROL+y�R��Ƭ�id���Z(+�\>�f[�Iݔ �ڃ��ⵄZ7�;�&<6W
!�8���]�DNz@vUί���4��c|]o�r���֜�"���U'v~���N��8�lh��@
j�/���l�~�$䜮:)3�|ǹ��Q�d�.��b[�a�P&T連lD�����agdϝ=��|Ss�MN��~�n�MܲW�L�~�Η�f�U�i���x�1vy\�L�sG��1�'�b�v�I����B��<�2����������jл����H�{�Wx�� 	�_�_��e�:����}y�/չ��aL��0VR����4��7�0׾ ����A��ȗ�٪E�_/Ti�X�ɤ�$,C����#��'>���-��H�׺ÍH����:.*`��r��0g�o!r�2�W�� vT�A����qF�it��;_o�����S�s9��l�V.9��r0˔�����<ꮤʵ��/���ɟ�Z����׃N8����
O00������[��!c�k�2�o�#��g!�ۃ|E���a�3��ߢ�G�c�K��-@!5P&)��3��	�sO2���p)+��2�E�Lp],�W8�iT�OY���'�M�'�#�9��1�=���^y��2
�>b�>E� �.�/���;f����('�(���kO`ʻzQ�px��ū�!%���@'4����A�}t[L؞=|��&���U,&'e��%�*��1v�m���H_/��ͬv��^��x�Rui�7QYv��%U���/67��C#���!����S�X9E!?���2U���6�"<��1VY�H�Gd߬6<�p
{���J��14{ER��DK^��<�!}���<5�A;�%~?|j���/�,j5�q͡v���Z�A$Л5�A`"״L2�)7����
�[C<������u�L�3��6����R�\k{I d���V���z�dOFT>����Ad{G��qaі^����P��Pu�[�S��Ǟ�X��y��s`�	���;�$��ߐ� <��{ot��q��\���`y���9��Y���a�Tr�i?��ot D6�����)K?�n���+�?�C��;Oe��C��ER�;�`�Z�6�������h�U�1��6�������e��S#�MCt���M�X[6���N�_�>n/Rx;~o��^X�q�C���4W���m?p�B|�P:��祝���Y\�n���6f�T���?��#�l,�iE����溸v$g��]'�N*��"l���{۵hi�
������H,{��**��L-�Idh쫯������-%;�4,�ouK��?CFƃ�M{�U�^ٻ���?c���S<93~�
�-�����7���;���;�>xy�B+�ň-+m��<m/��
���A��b�
Y����sP�{�!6�O
�\�b�.�X��d��1}9�:NôȺV�w��'R��D��ʶ6�16?�ԭ�f/�z�ޢ3ڮ]k����݂����J��H�C�����vN6��ȭF������w	��h����[͠d�_+�{�_Vh�W��=k�I��'"�;7S}O�w�A�U�p��AT.�ٸ�Mm�l�ܛsDR;<�S?O���;W���ɶ���2�� ��{���T0^w�DX�2\�^VD�j��6c�kI�3��j�4��|�D��d�i�͚^������)�B�ٷS[��i�#�b�����9��s&�3sme�����m���&�(qU���W�?��s�S�������ZRjo������VI���ck[�@S�(6B�R��`��Q(P��_���ߡ�:8w���q#�e�7�#�D�8�zק2�>���_�v�ş�wuJ��`M�E�M9��O0�*��[g+*���L�XyL�	{K��*�:�Q�Ч��B���%��U��
�K-�*ws!�B}��6�����14�G�w�2�i���ٞ�;�f5)�}C���Ǵo�a�����Վ���b����@�ʧ��v��6� ���B�>y9,�=���T�xW1UӨ-'�fL�����
�]{B.�����ŹH��0�ݚ>�4+�
�e�)�R�|�
EaU�U���|S$���+!F����K�=ڢz�r�l�6B�}o���zr)H���v���:�݃c�O���̘�/�%0���C_����UK:��` bf�;]�'2(γ��'�"K;U �i�X5�����:��Uފ��w���ŭ���qHkIyќ��S1)�xJ+��w�w���/R.�̟�XA6�æ>����>��
zސV!E�	��Z�f.�x�*�W��r�BF'�q�֖Ѩ���U.R6Tx�( l#ag���������s\!F�Y�K�,y��;U�q��"��>��^\�ڶ�V�ϕ��t�Gz8M}�D7���Q"�jhU^����tv��t��U
;*9��w��}�ڑI�y�M<U�.2x#^~���ޯ�X5�tGP��#$ʴre1�oH;�3=+t��SмY��J��4����5W-x��X#Ś�#�
����n#s�o���q��>A���;���Klf�
���q3j6�N�/��S��O[��'����^�%#4&%X0�����ؗ�*�p(��Ə?kF��Y���#	�F粁G���:�����稡�J7�fM���Ǽ,��N�^�\YxO�K�K��T20�>(.6�cAd�%���w{����
$��[ע�W��4��@�/�Al���8-���;� qj�6h[����5��[��Z"Z-3u`2�L�N
�Q�,�Б��)�������.a�,�BC���5=�MH��LӰwŰx�	��]'����c������\T�3b3V��xr�\�w�</�d<< �Cj�p�w�,09����Y-�p�Db>�"y4�\O�tqWH���*�L<�f�2�
��0IMa�`����׀Y'j�X�&;����#UN]sz����@�!�<�vz5+Ɯ�'y}%�FH?���G��ے�N�A�e� �4Z�c���qm6���`$�_@��Q'Hs��f>U���I�{Y��v�<�\i���!:���])BC�����z���Qψ~�l��G����3=�Q�k��{�v�e/w�>CŘ����"�vTZ��DWMr�K������0�̫��v�~y�FU�U�]�e\�9eVx�J������9��� �S?^����($���b6�1��~�
d��@OTP���S$� �2��)}��?���d�@Wh�S۶8߬�	.a�3��%|�o��[�r��~�0�K��<&�}p�w��Pa��������9Yt;a���X� <��O�C�޵�A�gh�C�0��т�w��^�ܘ(��\Q.W�9�>K>��x�I�<Լ�ݙ����`q����4	�L��؆�d�����1�\X0@�'�޸�D$^c�� �=ߐw/i|�w!�����fx�w�)Q�V��L�!{@1�O�9e~������x����9�	L�lÇA�<��ל?�Ԏ"�2�⊩}��V'��`й��E�?{�r�g�%98(��E�\ґ#g��d���H�<n�S% �&�
�%���*ֈn�}�}A��n�S`�X�	�M����B��&Ho�ꮯt\��L�n+�=�	��$�;�� ��aƀg�P����ɘ��E'��r��r+��|c5�P�OB���
l
A����a���?�U!z�d��-W��,[����Th��L���/�ю��0;>�n�A �ȇ
rgg��?w�?��b�� 2�	j8�!ݻ"�qK�[Z�Pav��cv0`��V��!�)�e�U͕��@~~��Fj�q'F#G����c�����9��o{V2��-(⨴�Dw�|����
���ԷH�j��|�>�b�Yl�1��b��L�
�x�@��M�z�5����TL2w �k�'��-�2B��=�Y��r���(�rd�4��kĮb>t~�ЩeN�����>6�������ޣO�M�f��/G�$B�{Q}�'$��6�Sx�&8��7��*T��BO;�3��Y[%k�'�epy���-$�P!�I<����W��i���&���$�_X�%���	� �jP�"%�.��yI�Ts8]e�&P���<�E�c$jމ�E$�9[���JD�L��6|�]h��!���;K�������:5��U�n�������������@��)�6�Oi�{9�����l�j�t�:4�Р�R3�l|Bn!���W��bHvY9
lGd�c~�a�A�Q�̾�^[L��=�6���Ǻ�Wc0�k�>n�Z`՚�V>zl�� �d�Zi�gb�0�a�x&׭h���G�D,�G�g���VL̛{$i->�F����Ɣ�k�Ϡl�EK�ϫَ�c��I��yʌ���U�]�3	׸�;����xR�-�`��������JNP�_6,�U�)%}y�m6i&k2%�m�6K�p���q|���Q#�����U��F2U®���w�n��Ƒ쟥-�r��P �@�`ն�Zf��(����?@8�"�QR��?�E��ȥ�]ÀW���ౝ��<���Ž�b�]t�q�����((tz�u�	Ѷ��aD��܋a-u�>.�� �RLHR=xj��4gգ��D�6S����� ��U @P|�x
� +9�ހ}������6�������x%z�����c��v��W#������H6o�w(:�e�Ga����S�Ǐ�n��+�[����Lem8/��.' ���N*HWP�����r�"����c�H�D0�l/��P�G���Ҡ�qp�	�OW��c/:�l�J�C�Muު�[2�/}�� �aEj�'o��� 