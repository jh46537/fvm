��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���ymc����#��בsb]b�k������p��<�xÚ^Z��ߖr�S��7���X��[hEa�fv�"%�%�Z(m��3�����xq��k[�,H7Y�C���=_���d��;��ˈ�ɥPSJ0���r�ȽD�"æ�Jҡq3L��|�|b��+�Ē���p�-������x6�l�E~,�*OQ?q����g�CW��P�ЛYA �3ex�{ޒ(pj|et([1_�c�5֗Xp���d[%�r�޻zU�(i�m�hZ�˔��R���S|B4��T��	x�[�N�*�������pB����a�]^b~������:ї�5ҩ8d	W �)��Mm�ԜP�Hζ��z�o��'�"@+Y���ug'��e����y�R���a���E���q��SO �K:��y�5!kTF��[�NHC1~��'��l2n�o.��^���t�3�*�UK �}�1i=c��#8v-b���~R��*��X��>��J^����v9:�^A��L��ļ�1�A��C�3��I���P ���
A�܄qz�{�x��N����b��LAdUF�:���wHN}t�e�$������fb�c�m�:���Oz�QY�΋���"V\"��1w������#� �R�L�F�`�F�7�W��B�*0�6��S.#F���"��]7�BB�B���)ӫG�ʦ��*0�qy:���l�ꖁ�V�َͺYD�.����d��pLkWFk1�LMT[ez�1������ /3�Q,��ݡY,m�igA�T-n���/�ҷ�w#fT��2O��
g8#�B'��_)�T��u���@�|@tE�T�-m��;j�L�@���Poau�s*f�(�<�]V͉ڑ�'��M��q��}S���O����؆k�/s�pB�{�_�_�m�F؛)Ų�筒L�4H�����f�j�I�I#	�Y.��TaԔ�Q�#C��#�x9 �����Q� ��>��af�Ozw!@������<\C�^b��?��.(�y�zL�]�ތ�a���Ȥt�*
��扗�m���7am�e5��!Y)L�#f֤��=K��W��� �k�4�8���;�s�8]�p����%�&�ϒ��d���Pv\gγ7E��4a�st�-�Q�'�5�6��c�����/J�������s�����Q-���@� �^��"���@�Gn��Zsɖ/ڑ!�n$C�o���n��!D�/���V����<�|x���}��ǃ�(x.h= Ե��Q;t?1o z�l�GԒDU7�şi8)��� ����[��+�_d ?Vb��q
�t��z�ۤ��[7�ݰm��4��L��g��� ��1nO|:ۨ$���hZ;te�u�f��jQ�-���.P��zV}��ce�ny�p��|����#X�St��"Ͻ�;�.�j��L����I%�r综en��N���EXK:	9�ϗHq���#s�=�t%8F	a���~��T5�
�@h���ۡ��tё����܍AKQ6���ʰ�@pP�y)�|����@�gܾ<�s���t���$Zxf����=� ����8��f��^��c$}~��FPL�m>k Mb�M�h�����CW2�O*q�J��[����gh{՘����a�^}���
�:��IJ-���Od�VW	���{�>:i؈ut��B5;��� �T8�