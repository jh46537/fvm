��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�q�E��	YjpA������2o&�0���c�LڄX?�i��+�#��7J�n北�����J��kƧ�6���+{E�b��pڢ v�U��4��WL`d%�Zx�Һ�|�N2L�\����-�1s����#�+��l��"����1,h�'� ��a��I�k����^	w��G�Z��k(\H�9���# \����5AA�f��~o�ItMi������)Mn���e�4eӜ�^�����[)�F�0�?��~��w(-�f�sS��c��7����3��/��ֲm=o@=0�*QR��$�Ym*2�ծ>"�j��MZ�)є���8���'.��]����Ai��b$'�c�]7�a&���S���,�'1�O�U2�"�7�;@�医�.G��C^K�F]���_�3ϸsN���ј��`a3mWQ����UJ��|���9�~�4�<�>R����t�����wt޲�MV��D���z5}�)�����F��º�q�9_��bX�����}�d�ڨ+5�8�j�3�b2��\�]Q�G�d���OWQ]�1�	�>O�Kb��#�<�����n=�3v��ޅ�b�zs��g�۝�����x�w�hAlz������S�K��P��I��-p��OĴe�j���O����ќ�\芷���#3�'R����*Zr��\0�{�N&�����g�x!��X�[�`Zp#��RW\��.��C���ƹ�B���uMs�V��	�\��7bL=�H��&	p��h�8"�X�V�1F���:�S�-0gD�/��-���^���ݥH\R:
�:7軒r΃8�kVq�W����ܘ�^$�F�C�v���RO��@���bī�
bY�3�8D�G�l�Q��+dE��*̵I�GR[��,m ^	%�L��!sf��f�Ъ�E�q�tC�ym�4<����^R��nOrnm
&�<7L�9�[�2�ax2�Q'��d��dC����'�*I�z��5�߻ay]4�j�P�/�րv{�ɬ��Q���y`���pL>�� fX^�:�*���]<pP���J�3r�K���F��8[�4�#�����1�ÅH#[5`�|wn6�@�{/a�O����N����
�X�|�haE��܄l�F��\_C�w�3��Y"{�	.�ND0�HBVF���g~3�O'a�#�`��(���٩�Y����r�#!�����#�~�ǭ������4&�0��#I��^��G(N�ly�kT{Dy6�ƨ���B뚸od6\�(F��J������F/�U�k!u� |������E�?Y3�-0�5��Y�X{�29ip�mo���y��B*ZPF'��#bEw`�z:n�r�0�G!:�G��R 12X�a�"T6�w1��u�-
�͌8(�]xم-1L��u�cB�2L�7e��W�2Kr `���7�����b��h3����Z��HZ OI�����c����)77ˊ#�$�z,��ag �?_�?�"�#V�T����A�|��0��	��R����z%�_Ȕ:�<��]!k����jZ\0d�:r$���;�6�O�ʓ�P�YS���aoH(�]�x�xy�VMS-��A(���`�_�F>VX���ZL_���=%r�HI��S���C�j3N�
��}*�/7�u�J�Kq���V�m���ޯ`�zk[�7��<�[�&���j@�)�|ى�p��|@a)�H�o�B�Eé�]��	�0SA��Sm�
loYEpJ'�.�]m==T�,?P׼�~,Wgߔld1]w�j*��
�9>[�0T+<��$�^-`TI6*�`Ɖ]Ņ�Nd���]��X奝p�O�t�Z �◖��1��x���ع2�B*��u;i{j���AB�K��p��w?�-)�[�6�T_�B�# ��X}�O+�+&��P�'d_A��CX�#)��I��a���ڢ�7���4!D�e�=��JZ��(v#2豘�����k���)0i^��ԉ8;�A�Y�&1CS��XF6?Z{�T��Kj,���$��O5�)Q_�q%ݎ�.R�8Ly�F����to��!�]�� ��Ɉ+�d1��UJ m�p���k(D3��׍���r~cc�]�\�ױXC~|��g�_�v!�Є�k�^a�ă�e��]���d2����<@]e	��Ѷ��" 0<�Lw��9�1�	��M�p�|K~T�����,jk�W�Q�#�K̭Ln�ZO,0�R�Egq[���F�:��;Θ���f
�:�
�º���z��W }hͫ}��^e�<��o:�%;YHWCX~����%�`m�(���)g�s�z��w�����S���Q��W�'�Z��ָ���=Ja�AR�GQ���>川��G�jm���*$�V�,����-gTg�Tl̊B]�O�4�Ьf0_M��U��6����[����Z�!(pG�d�|�qM�n\�+,�Sf��Z�q��i~�KS�99۪��b%������~��^0���o���Np����{��ߚ|�&H�=�j��I������x��ٟ�-�|v� k�]wL�+�Q4�f�PP��Ng��ذ2r��F|*b�X1P �9��