��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]X@PQ-� O� ��G����G/�����!kY!�w�cZ�5�iϭD�M�W� ��-ݲ,c����t3���b�!�ȋUB�l����́g��)����6���%�!RF/ ��Dr~kvxK���xp�Uޢ%�V�d�z�����9;-m��;o,bY�c�΢&L	�
\lDo�}@�����VNWD#�!+���Y�vs�1	z�%-<�F�4�Z��%��Ү�?��Uܡ#ʓ_�ۮ2�O�PR'�)��;�(a}��t���F7�ւ�[̒�����۸��#4ͤBJCMT��8:./WHI�� ������u�(����fեe}�r���!��ם��٩$Ox��/Ȉ�&g+ z�Y�W,û67f�w���P��I���i�=%G���O\#�f�R&c���:	��9H�}�t	�_�r�͖ <�Ȑ;%� `k;[ݷ�I�c�F�a��It��H�QIV�-�&���x0�DCq�4���UVe��x�<�{ִ.\P�����	�C�k}ƄT#�������>�Vŧ0Z�Q�눮�9�Y(>k%L��v�grJ�Q�c`�@���Ҿ��)���kH3y:I@k@0$��Ҿ�$����{3���xR����RQ\��pTh~�N5\�ǭ�Ͼ�;�)�۸���"
^�ML��3PBQ8�m��c�#�í�D$m��8�榄�8r��(E_�p�N��ve5.�b�mNG?W�����\�����'1AW�F)���p��6��(�{��&��6��CN�Ҳ�~���դ^/;}���Vs$y.}�5�E�$�v��hi��A���H��.$��n&��؝���X3Q��n����$9+r�ȹB�x=���W>&ŷ{E��3L����Vy�k^T��ۦi���R:�`���aF\�����2�ހ���EkxG�}�q�4�p7��%;r��{yf��Em|��W+��2�.6�G�7pZk+"��������u���V�a�W����+��>	���mI����L�z�Y~S�c�����ao(cp����G�1��G����]1�l����d@7��ί���H񋛡v�ǣF�_�@�L0���zkY��Un�ϼS������U�;��3Nm�s��s�v<r�m�̷��^E�ww�l#̈��b�D(�}�L;�8i�B-
4�Q;�cm�i�]�x��xS	C�d7��VN�E�|m�ƾ�G)8�6^�t_&�wpt�	�퉁k)�iC�9b"c}������Y�ʁd�:0}���D�>L�ö�ם�_�x=�Oz]Q|nm����!���Gr��c�9 @ܢ�����V�|dF!����U�=u�P<��Fj��4ގV�Jɛ <�t�]rD��ڶ��!m�Ͱ�P���k6���u S@����::��CS���V���3��#qP�y>E�1����R]�[;����RC͇{K�"����ʧ�X9�����h�Z�U�c�S���v49V+x�Ϟ�������{�[�9,0���)����!�2J�����f��!Mጄtz�gZbwT�DR���.]f�Z��"n�f�-���4n���[�N�=�k2�ˈS�I1)8��w6w��ӫ��v�����:{æ��!m-C.��v�h
�~��P�;�p��[�0�c���VmC�8�w�`��M�x4��u�ɐU[2�,���qJ�HT�+�8�2!�0k#�n��H�N�b���,�E\�`�̧��F�9��\S��D ���
Y�/�. �e�V�3n~�k5))Q)-6�]9bQw����b5-�6 �KIQ�{7tpÕ_e�4�X;!h�$�á�P��q	�:}�Ur@	 ��;�W5���V/�Z�q,l��Yے��&<c���JdX�Pq�����l���8�aa��\���tg)����B�^9� �У�$�O�'糎"ߏ�bt�VJ�3��YM��NK{�ːoڽ�*(xsH�s�|�oF����tLn�i�.n���b����t�8)��1J�)��m���O�A���?�(�Ľ��_^�{�lF�?y%��K��[�uuȘ����h��t@�L�m�ga�CBr�8M�Ϗ�m3X�nd^ϱю�#��d2�4y!sס�+`	���U*��l`��"���9y��:~�=��g��B���~z��6��"K)FL%�v��%H���R䟎Av�zb-������nИ�[gb2��rO��l�>펫j�h\�x��ú��A��Xp�h�*�2��d��V��
���ɼ_N ]��m�FΟ*��+��8ؕ�I=^����a��)<�C���cE�@�ރ�s�׌��$�~�&�v$��y*;j#OM7�$8�e�F���=�Mi��EZ�@��G�d��|O����
�^Ux�����mո���$Fqб!e���(�X���J��%�o^����P�?�k^��7ohA=G�*��,��I���"s�dU=�ﻛ���T�ϊ���A�<�M��� eC��b?�,�⃜��17t��A��+Ք3�`�"һv7�Ƅʦ�
����I�JYv�usx�O/��D{�ēD�U�H�\r�`�������Wt�}����ܱǕv�})���'/��VdI��%�2��m�d9��ɶ������<�y��JKI5��oB��H� k��kQ��7��m��΅��JM�(���@�)��A���Ƃ���wIIx O\��Q�բ�t���XO/R��
�J�v�uo��g'�*De��S��S�ػ�=�%��F���2����K�'cFϛ2�����$��j��{�sS_�&FaѸBa/,���L���7�X�b7���r乭�c��� [s�]�}��rֳqU�/Tw�b9�d�1��.�
 ]�pM�/L�#Ϸ�����K̊�����yٓ)n*��^A�6�9`P�����r/�r�z�sԲ��oW�@�p�1��@��5Ə:t����v���=G����w�[��{��/㐊�e�6X��y�m�����o����<A~P�l�������=W/��lh\�С�sP�'�6�S����T6<��{1���Y���q��=T��$dCi���!��H�qG����1/��;�#O�UD�o�LcQ���»[�PK* �?�R)�T�W��FH�j��p��,�	tv�,u<�ޙ&W�:	�g��A�t���>����Q?��o�i��m���r�0����a�9��Ȋ�Wh�@^lA�o���e�� ���&.ESW�һ3�Hc'���Ǖ�7!:�2S��d~�-�f�������`�%�b�'��(h��,L��s��꬀�Q����GhB�H%�*T��[3���͈4=�Ǉ�?��ײ��\���g�D���/�Ύ���aK��?��ڶn�*�+�ˆ��*��hm�Em���<U�*٫9��>g�I�]��^r��q�|�H���DMW�h��ETl�Էk�"�ɂ�4`�&���״��g���O,euU$#�]��LRNƝ"8�7�E|h���q�u;({KW��%�Pt�diS�} �_l�� 
	b�t	4gi�Fd���}*�Ak��G��T�o��Zd?���]
C�����>_֭z(-Ff��\) N��q����}|���5t��C�����|����닁��-��X���Rٺ�C ��G�<t�#{;��:�X�P/�J��kI}Z�\�@QNk�>`d� _t|	�c�J_���é?������m�z�g�����D��#T���]���"��US�d�N�x����gT!�������t��-'f!K�"�CV6�IߍۋO�~p�z�n����$8:	���6a���6���ҋ0��� M΂������K����lhNP��XX��edz�1Y]B���sgpY�����%織V���نL��P�5]3����i1�1c��k�@^6�Ǽ����Ę\db]��jS����H�҈��}	g>���:��)���{�zAt�Δ�U$�� l���f����R��E���� �����/ܝ�iC�xVy"
YAfb�lG�L�U��9M�lh��?SR�,����j?��NO���v��X��ctJ����t�F8`��bq#O+�d�[u����AJZ���v��K来��
e6v�c�-�V�g�+n��G.��s�ME��=V�2|&(q"S��e$Va8�ΰe r�j�o�ʖ�bM�n��Z�<��̣����������-p�|�Ǘqq��}��~���d��3� 2��Zk�b!����K������Ȟi�&�-��;7��9A��{4<�?��NA�MBz��/��}@g���/Lk�w��Ԛ���;��#k�N�^P����7��5�ԌLc���:CA��]���m�H8��K�BJGz��;AF����G2���5.~}�f�'���b�/�ޤ:�6�s믙2�<�J��-u�L�m^��'*��_�ʛ��͹N�E�z����g�`NT�r� �Hw�D%|*�^�hI_�����z���P�v!�*`��d�n絼>ᓝ�2a��]�Cϔn�!��w��_�o!�DX�x]�Cr/�E9E��RF�R��;���,�Z_�@F�C�H�9����� �*� O�F�Mrk/;U,E|�����y�� �i�vCE�VL2R�r��W���l�}}��nU��v�S�b�8�l_t5�w�����g����M����7�dj׉��L��r)h�f�H~���h0��~4Rɡ��~�笟^�ƪ��a�
����N�|_8���?��$U��oZ�/K:#���\��0�?��F�$+��fe�ޅ�e��+}���.��r�Ү�d�D����*�1�op���|Ww�Ǜ4ke�D�?~xg�0:KQ<��o[Fp�.a���Ye��%�����p`�G%o�$����Ȼ`��|�h�K�8]L�8XJ�W{4�I�pC~םL�~�o��>~�����X��<�!jч+�����0�&�i��$�پxzi�]>n��y�����8<�7A�tR�X�n�;�;�E؜�?����N�gB*�S!�uv�N o:?��g�k@FB��	hEު�٥��b4KH?7�з�7%�sM��g`8$�^jO�����F'��*P_ȍs�._&�x���*L�]�"���9�f(X�&1������|������^:A�g׷{+��J/c� ��N�����bb5�x}|S���$3� W��h%<��@��:-�V�>���=;jKJ�� ��ހQ�{;�bXy�,�%�G���V���b�ѕrs�"�b����y	��~Q��j��!
E�&O츫F��,{��na��"�`�9���,�ѣ�T�
4?d�{6�!�O=�b�����n�+��-?�m<<4۳k��SP�!W0���D� B7�;��߮kO����d#�P	O���e�QD�*���6�%����nAE�eO���� �J�۾�4r���){\�瀮�@�K����B<K<���P����Bt����#Wr2x�ȁL����31ԱN� �h���܁awU<c*�Q7���G��w���`�:���RP�����n8�l�*~,Qt�yC�Ԩv&W���C����S&<��yO���.�̽�~�����u��%>S�e���� �i�z_��:�P� Zu=n$E��zXp쭅��K�Cլ����ȅ��)�~L��@r�	�M@�������|=c�&��.�0!T�<\�Í軡����[��3:=��׋�3�Z$0g?Rx
bհ2��p2D��!mn*�y^������f��I 1�����Q	j�=��E'"���@ݗ$k6Ǵ-���ΥQ�Y �A�˦�����_�Quyo����E5���_d0�"�)gx��"b�aeE�������f����)�$ppɰ7�q�rm��&�6�:�������`��ߧ�6��g���o�K�K~��(��b�
��p%К�ں��Ώػ�I�\��vp�؂Ý�<a���&����ez���� 9ԡP���؈8G��]8�����C0��m�Y�+թ��n$H�qB����@Nf�RI��
�5���rR���*IbQ�~��o���mA�����R�m�r\�Mf��iJ�qг=7�ǔ="�����m�ܬ�����>r�n��ˡd����]��
�֥��7��~����R���b�\g����X>TdK��.���>a��"��M;�E`� ��{pJg�C�z�?��$����{X��8g�g�W�]4�y��߻�fFR��ly"��چw{�Gޫ�ٲw��%(�9Q���3���aޯz�����B���Ҳ[Q�B���$�9�O��5�z��1�W��OI,Wќ1��K]�0�s�[>��P�#���u .������yhJN�pLeő#'�1I�b� �����+����y3���XM(]`�4:fw�Q��l�.�z�9�+���A�˦&�^�!�=�����M�*Z.�@�B%.C�����I�Ck}�H�QxU؁.�j�<r����Y���4���������ൄ4�Y������7Y�$M����J��&av�Q�Mrrh'.����_� WN�H�I��k!Tג���x��g8��qgP*_�%�hZ�b�u��R����5�E��1�'݃��_EK-=���Ǖ G�4J��rO������@�H�:i�Үʂ�L]ċB�λ22.�񆍩<a�g0�W���t0�V�7=�Xᜀ̜�c@:��\|V��w3u���mDEѕb�+	�Y�������}��elҐ�=��=t�`n�_�#�����K�H���%J9H������T�u���b`��;�{۰;ř+B����>!�F��������I��?=$�����q�c�rg�0�ؒϘ�����Q�owoyBKҼ�͘��Bj��J���';��v�$O�3͡2�Z@Gss��Gʯ�a��!���`]�R�{��<N��ʧ[I\�/�`��f�)2ʹ��*�9��)�^UR��ٷ<֊�� G�~[�Fc{g�XT��)�ܝS}����t�i4����g��R��B�D=�{�=��ba�:k��~j�=B
��A�猭�(ՙ�)� 2
y�ӕ�9'�����@�ԗJ�|/v�1�]��x�N��]�aU,�z ��5F_��������9�hk�K�*$�V˂�
�<V1�;q�:+�֨5ǂs��y��B�:\���3]�����א�_;��?S�����]l��y���0U�o�N�uTA	�1���['�2nI�om����I�L;�`׼ŀsO,��|����۠�w�>����e �$�M�C:�ۥ� ߣ�g�E���[UW@T|H^�J8 w��<��پ���t;uyp�\��m�����h�f�"��i�F�B��6�XN	�����n��@L�aE}��ݡ}�C4V^���J�����)��*��x�,$0�	N9�mG�O��I"Э(�o�3]��$�q��D��@����[�]\
�GJ���Mra�J���T�yP��UQ-�|�7'�+�`x�xx�ԡ֛u�6��&�J��C�����o7{�"ds�h���i���q�����bQ�J�8��Bѣ&�$�r⹗�p����kp��r�1���
{�箿����72�[h[ǃ��nc6�m ��7ѦJX����V@n7͟����L�&5�ț	^��7��
��Yo��3S$�k�稨N��0������Y"�%���f�0ľHy�ȍ��w�8�I�9�+�\;���h(b��ۧVO��A�<D$8z�SO��>��'Ut`��=�Il��V���*�k��*���X�v{�����V���ػin�m�S;kNǝl��wx]��tc����@�R4�=�B���RY)�����G^W��=͜ ��X	����`��ч����")���9��p���W�p�)܆a�4/��b�E�1r$C�Lm�V�;�}�hh�)��2lM܅lN(�Gg1�l�H�T�d��b~XOrl b���Hvg�r	v��y$����i@VgS���$.!r�R4Y���ow�3u!�A��U��C,�yޘ�hZ`���mn�X)�1���ϛ��ɧx�c��ӄlH\J���G����k��pw����I�г!+�֩�z���R�j/I��#�£r���tF6F=1e#�;tOc-��ț�� L� [��I ��;{�9>f���S����tx�g�G�{��f�)w�@]_;�Fb�'N����Ei\t�}���♳�����h��I��8{$~S��N��Ф�-��*�3����D�Ɔ	6UnJ�4|�S7T*t���dLL�L0r�a���ړ�b���7���4�'d��U`�i��W�Tʉ��:�y=����/��[�ѓá��K��M�ż���#��2�TE�(^�}��m��ox7`�����5'W{�1�,\��߿[R�H��̾ޚ�)��=�����O����^H��Z�3��n��e]�t��4��=��˹/��d��h�q����jxh7�P����尹��5LYt]�߿TmB�M��^��i&x�m�o�I�����˽t�|ɞA׳��I���٠JC�u��	�)���̌��͐=t���x3Χ�
�?v�kr&���}g�Vc(7z����_�3���<ƻ����_%ݷ�����A���J���݆ M߆��2�]�O� ڑ֮ƀKL�a{�ҽ���ϸ~Db�ܶ�E>pb��Ċ�R�J�s�s�Ύ:��w�s���^}V����
ĺ%�ZN5@���L������y)_!���SP[�"PL���?:���u�[ֈ3Q�m� �_����M���B_LV�C-71��A�;��>���\O�o��9 ��-����
���g(�H�UB����p_�-u��}��NyS}<�
̀��&<��#_c��̿��]#��(P�G��p���Y~}���`�(��A~��|g�t}�=k QE~�d-v��G�.�����r�~ǉG?���LF2+��ͧ�����(�y�g0�H(���� h�y�f��ٽl)F$��*f�ٛ������u���u�x��Z��}���.$@/R����h��P��]i�����Ez,b�$W�#�R�K�������?�w�GLI6���&�XA�(�`�!�4�u�F��&p�1�O�d�?�#�gX�HP��Q���J�7,pZ�����?֟�见�}S�9���3:�7�6��V��*d�V2�5�r��8{��
�����f����_�)��I�����]�,��[�Q/�x[��J���h��Z�5/�f�l����([�)e��$��ͷ���gB�Z:��@��?V^����~0ֵؼc�L�H>��"}��rL���s{�u��9gR��T�t�#�)��.f>���w35�02V	�0]�g�X�O]{S��)���V�[ÛǛ=�s��]B����E�*�;&�D�N�����G�Ƣ��@�]P��֊!s?�-��x�d1�C}��@�z
����=��3��9"
�3��`Y��3���Dm��Sg��,	'�񃏒�D���=[��Th�	���w�����P��q��P���G�Y�c�j���[$�yRL��z�8�BS�Cn�:��-%��H7���~T�H;0���:��o��
��uZ�w(DT �7"��&
]�@������XIs!{��Ȭ�ˇ,���
���F��%T��h4�uX�����*���f
-�g��A:κ�t��c��`�$#J�ɉ�e�i�_'Uz���Yz5W#�W��Ņ_J�q� V5C�$DxΞ����B�ML�'���+�>����g�6R���A1��wW�������L�u�Տ�������Q��7.��D/��	!k�C�0���,O � �:�d��h�ȅJ��`]�a�ީ�c+�C>��ʒx�2/�<�$Xo1�H|�+d��|j�Aa�;/=+	b�-���M�Y�(���x��{��.�'��).k�&��|3)��ka�
�6�U�t�3G��Oǧ�B�:2���Q��'<@�$Ѥ�]k�I�� {]����)�6j�gFy�d<�q�Ӎ`yD�G�Rϭ�"Fȥ�cV�b>��xj�b*V�L�+��6��.T����[�L[�G#�;sV`H5������P�!~G���*株8���o�5�k��ﻹ�q�R"�A�f��돖�㮆��k:e�Ȍ�������g����SImo���隼$J��<����w����g�!%S����B�����32�HOE�9��y�s�V��)4�׎��F� �z/��*�4�}ٖK�����d�O�"��D�-[���6/v������=�g\
��-�
���&6�h����gؾp8%�\r�}�o�r�B��7�3�pI�Q�1�Duŋ��������i���z���ع���Z����0��XlE�bW�Զ8�`%�bN`�Wv�;@����5�3#ŕM�k���\���������z}�)^BV���b+~D*!5�s�Y�N�%􋊑�w���m�Բ�B)�>���AI��^^S�������0�u;.�RTHpZs�m�DPA=��P����{�6ո0Z4<�bt@n>�u�n�y6��W�v��+��[�A c���l�Ƴ�}�n���Q��Z����3���K����x$f���(�O�=���8u�$;�~��:�]��K�`��K��	�C��cި)�̉3�ׯ��Ɇaxv��Y��ށsǯ��!��6��q�6��F!�2�`���X���2獂r��e
y2M�4��i�e�-���[9 �h���4}�E�uஶ���	��t����D�/�Y���D��F��ݠW.���R����ੑ���h֕��^ ��M(�c�"Eǋ��4y���pC�8l�s�uǝ�3��|���HP�uPD��N2E��'6�]CW�sG�;�/�[^��V)�n�}N�q}���w�p^_ʙxu�d��j|'�O���	���X��,AIDO~ï
��.eI��B7��A�-�ǈ��|h</��r��4�$`�f�e&Ҍ�~�B4������"�v���[��b�r�J��86�^|j�ޣ���D��$w��%BG�Dmá�-
d)g���@ks `,����)E��̪Mu���X\���:e]9#�f���2G��������2"@xH���e�]Ä��� ަ����sǲ��$�� ��Fb�5.;���r0�������=���G�{�u�� �ψء�-�T��a@_��#����Y�%2�ٜ����K�����C.��j�G7��XV+z�՚Ȱ�񈄭�-�REx�C�Ff����(ʼ6�62}+FJ�b���5��*��*�/3��kѸW��]?��k�V쓁�;��YO��EKE�	���I��+�GN+��R>t>yO�̲r��rZ�gSш.��\�*G�˹L`�"��������6-���E��%��_��Aӈ���PNVcg�Bp��%�3:��2�����N���T�q�h}D�����"�$+�o�^ݿW�_��]7�4%P�j���c��0HS�!Ryh�p���������7Џq�u���I+�������hs&�>�]G��As7��M�5��2����?.��k�!A��G�C��e�qI�וW��=#8�f_?��f��u,}��S9/=H^G�-C�U��
q|�ɍ��BCB3�~��ۊ��W��}@���E�T�/G����H���E�>�f�\m<mBT���^�Y�I��1�.��/0�ے�ΊHHf�e^�t'q�l�bp�T��:�c�/h(����C� 8{�f#>x��������(]?����Qɺa��I�J���#��z���)fW�
�%�la;��D�r=���e������I~v�AJ�����_��P�B�Y�K����	d�.�y�!|��A9踔��c��R�`V��,k�S�����RTR:X��3.-����l?�Ԑ�y0���ׂ!�ۭ�:��f����R''�y^���K* d��@.�0�3�2ns��L�}��r�]c5XZ�U6��1��\�I����!��dZ����-�_
w�s���V����\u�ʮ�������*;�F�6F�AJ��#�`�"��A�����6�m�J�id�J��&cϾ��gs� g̬�b͟�����L:v�C	�{!%3�\Z���;�/�����Yz�����J�����nS�J�(��ש����eK���#��Q��#�n��l����ȡ�1M�/l*A@�.F����2���}
��c��v���wSb���2�I��⇒z,��~�j����.A�O��!�@&?�&l�P\m��P�"*�F��&=���V�j&j{t���N��N�m����o��<�_���\�T�f���z�M�`A+ ����K1�fׯBZ����+��$3/�'0LQd���q�27|�0Ԟ5���D�-��������3�/�9��VP�;5�%�?���s��lgݎ,9:��q�ƶE��|�?{���P2pn��y9G=�P�ǟ����?��Z�O��j(>;x��O%�%��k8Y
dzj���e���d���9=ޭ��^�-���~^`u�w2�R*t}�
 ~+�Uw8�TKv-̕qx	�t<跗��O�v��L����cͱuSAT�+����R���b��O�?��x���'CF�ڢ�f�-;��/���Ch�����\jꝂ����UW=Z�Cv�9��J�<Y0�y1��&�,�0������~���p��m�����P�#&���i�p�J�.�N�gwA��L<GR�K��+CWd�-ZUjE�3&�G��҈���5�Az��1g��B�=��8�Ý�W��,�ơ�?�xҒ����j6��<����K��o����nvH������j�k����lJD(ͽ�[�|�� �ɨ��߭i-�j�*xCo	:}C�$�Δ����&7��I��û��U��*��k�`���Vb����ݒl��E$�Xw���%+	�&��b��*��nIa_B�l���"!*D��Y��rY��;'�7��&Qْ_n�'�-&q���f�ۉ#���uXs-��Z�̚$�?k��h3�\::?+�ێCƣCk�
+��$�}'��=MU��G�z�S*�����+q��{�"Ѫ����AL�e�}�A�
^�	{w��1-'�䳍ʜ>CBc�ۉ�:`�p|���8/`�M�J�uQ9�5	��{�}��	�r\�z��N���!DpZ�ߏ\#̩���9U��<��a�PH��Q'"m� �A�����8G�${�,�O���1Yж�(&Mc���@�Z��\�� ��W9[�h��Q�+��<����hϏ��m���ߋPG�ϑ��p��F��ʵ���t6j��j�r�۝��R���^�9~��t�E
�80�:Z*O|�^�:�Gh��%�B/�Խb}Q�ě	_½ěm��y��9{�+��qv��e��f��0/�M)���E�)u���_F� Ң�0��	�AX"��#%k�^��&w��W�$_R7鷃܆� 1��0[3Z��AV��r��<%e��il�4~`� �-a�[~y0(h���2Ѕy�"��^H ��C~`l�k"$&�+��[��29:%�GH��m$u��p9�@筼l8�D$�Nd�r������չ�u��iآƲ��6:m�'��T��m���QKn�n���IX�n*�t����5��3̼`��������#:�`��45�y��E�8"���0D���'z�?��>7��X�SOF��Z��Ƣ�oJ�{���2Y�(�#��A�����Ȥ���P���P�:�+ܚ�X�ew������ee�Ay<�9����C�An�Jn�%$���I'!���Y��tI��G���y�����Le@+^�����"�HF��*�Q������Ξ��'9�d�p[�ﳭ��&>�N�Q�Jw�Γ!�!���w��t;' �AtB�{o���ʵ/����E补t���	�#c,Y^)\7�,q�H
�_"�������^x&8���(U�\��Z��|n���T�1�ʭ�8��� x��>������=/1;Q�:!��(�p��X ӏ��0��2~�_�o&G`��4P�UJ{������4��4��(�Td��)Y֔u��|�0y׾2f����:O9ݰ��5�s�ղ�ꇮ��z�&�#�OU�t�-��L� 19l3f��m�<��o�}�;��{x<��k������rI����oA.���"�t��U�Oթ4�=�g�)#{��;�Frĉ�VŨV�}OWz��}�[�÷��\'�i	6&*�ܐ�pZ}��|�j��h���Y?&Y�);�(.۠E�Z�T��2��VY��|�ʥ��9̵���Ø�>!z�O�G��0+�bTF��VAD�)R�����u�*�z�/�_�ʬ�I��ӧYv��0��\W`�G]L��uǡs�O�t��)�O�/�m��i�t\.XX�������(7ڂx����D�{j�Hܰ� �]�h��>��������E#3�ek;69N�Xx��Y��S�.�٠yj� #��D\Z'��MA�w�A��׮��I��<��jn�w��S������7�\#�loLN3�vU�G��X���N�W�"r���Q}qjg*ՔrB���WCe���V^a���P6�$�iOqeE�݆��ڣ�������m�<nB�uR���V�\�3X���1�=8�Ǚ��+�]ѧTa���)K���G�vO֯�<�ُCy�$\�E�x�}>i��;PoWE�s��Ix�*& ����P�C��B�:�uԵ�c+�qΧ��}QD���N����B�Jv�����,���:_�@F��r����a���`4��o)�\���)�C6��)<� .�F�7�򅍷z��&�ҸBEN��=�(�#�b�}�l�ɔd�Q��)���#���= ���uX0m_%k3bQ���O8�� 	���Ѯ������YVh��G!��V���w�퐿D����,�j��G0ll؁�k����T�4Q'��eWO���WU'���h�<a� ��O��ӉexP��G�?`������*O�|���	������(:XA}�Y� z�l�T�o5����'�`��*|�8H� ��UmPt:̼���%�΢`�#э�s�S��J�C#;7 ���r%���ƙg�j ���AG�'s��^�?�� r��k�d���y0l��
ZBCĒ���Ѣ��ֆǜl���ZϹ�^[�����Y1�4i(�MKi[�Rj�{�[mo|�)g�s̰��kx�v�ߩ�����3�v���z�h�J��4i�(�Jm�v����j?'�z\9>�\L_���~����>�2�r,� �n���D8��|U��Zѻ�,�k�#�b(\3�R�eb��H��?���5�t����
�p�$�&�����4@v�6-��Z��p�[?<&�O��G��Z2�ȋ��,���PB��2T�Dae�0�t�k2�e���
��X�Ű�, ˠI�>�t��<acQj���^��)�	U�[����ߋ��T�!�<d��J���V=�"������wҿMT���7%�%+�Nhj��M�l��?��j��Ń=�WA	VkH�TР_jL�
��3��`{�.rvOg���.H���v�p������[�߀\86���4�O�ϭ�	DySPl��Ҷy~�`�~6��}��c]L��GWs�v��aW�A�
���M��2j-��V�*�~;"R�k)'�l�Q \����D �8i�����b��,_����!s�2c4��2LI,���C��!�@�_j�D�I,��jf)p!���:��8'#�E���R���*����a�ȧ-���8tD-��S�T
�dr���>J�]j���q���dCGٚ�0~�{�_Ť,&�Ks�?;7+�ͱ����è#���4H�1X�q�M��z�,[v8�+Q�Ҁ�����pm���e�k�w�"���Ҙ�W��T�`l4K�Ƽ�O�GT����W/�_*p; ��1�eNbM�Ń���$4���(M/��^~n�VH��b�?��&/3ύ����p	�D�b���h.:�r�U����3��w�X����� �����FV���t����%]�*��w�@4�S�8��!��P����-!J]-���QW���XZL��������t���k��'���1�Եc�O`�,B�S�u3���r�A�+�h:���ٴb��N��������S���c�)��T�P�7�kvdw���#�!��#�%��\�?�=����?g�<Vy�:����
�E���$�6RkN���:d9�5鐺.�W*��}B�;._jH��]�b6cK��N��u�3�&�\�
7��Y�!y��1��f� A�'�=H��ly�r�Q�қ��.��S����QP�R@\v�Gs�;��a\~[6mVԅ��&(k���Q3�0R2�K�mm�������77�8��&�($J>�F�����t��:���V�D� ;��L���  _h�W̷����k����L	��Q�(/M{�挿��7L�a�!B��4*%��C��4w�/t�ҳ�4�� ��X�/c5��k�tOr�5MF���"�9���G�P���V�'�ȓ�&���k�zp��z�?r�`I;���[@��}�%���qת)xs�N]��9�A���H3�IͩC��poľ}�.Z�c�p�����^lnb$h���6��Hf���ǘ�t�Y� 㸶b8.��ఃڪp;6b��6׃ ͒m�gaX��!�p�Z�d�����C4y�:���;�Vf�v)��#r��U�O�ԉ�y ���8՝#�fug_`)e\���N�ވ�Id|���V�<A���N+ Ad*��[s�~�'2����bB��7~D�OLQȝ�x���!DF����n1@냏
��� _S��t�!�l=���nx��G�
-����o~��k@r��3�2k7l-Vޱ�O���Ζ}�$�
�_Vt�,�I�#�?W�I�j2c����y�҈h6N��IbT�@;��Q95Tq�(�%P�k������HԐ��i�ViT�奈޹��2�b$���V/���|q{u�z�8%���KP�^�k�P0=[ے�X%�u�V+���:��������L�y�:wݥE�փۡ�!��L�V���,�ۘ��}�7�_q{R�R�_6�]'�уh��1�>�~���i6�T��U�d�Z��CW@)�P2ߨ���o�����U% K5�e�l����i��T��{��ͥ���D��NnaL"l殬�23WTVC��o
��[yL���@��r�뱞'�I�^L��k5�,�sF�^�LA��M�4���W��ӡ�q|�^�@��u [�O�a�"����7��.�(&y�Y�
k���j������p��=yϘ�/���U'
�-D�>N�<z�^��-���y����`�R���"�|n,�n��n.�����Q�9k	�������hp���b�a�b��&mc��x�`k#�j#ɰN���4��WQX65!��-�*G��6*!��C#�߅����%T�I����8�r����3�7`�n�h��}���"�5uW�_T��S�gW�DEL�79m�h*�5��x�c��N���=�	��w�z+��Ƃo�o���rʟ���M��9����n'L�Oq��U���B;/���A���z��f�.�)#6��X)�zDto�[?�Bt����0��15~ t� �25�-���[�hh�����b����&�U���ؕ�3<�J�O��{�XIZ���ד7�����b��c����L�^��*22<\5���Φ�	��i9`�)��� �,� j��tt��o[��?���u�wc�ݭQɧ-8�Mƫ��'�y�{0XP��߁����'
�Q;'vUt�1�Ϟ8�NT*�Iw�B�<�6[��i�-���;�q$iX�U�}R�.����H<u���a��jvq��{-V��Q���gߙ���j�g����-�8 ��\��P ۋ+�
c���U���d�O�#@��nˊrk�OE�r$c�N�&z���7q�ljq���R�m����6�j���i3�<�iw��l����ӥCG��ER
*߇�q�h�7ͣj�kS��6U�6��� �j9��6j��L���w�6���^Ŝ*���5ZWyL�Dn��
��9�z֝RT���I`�T���(�;���c�46��'��t�/G�����4�+��E���kx�`�O$�	�u2�Z�D�u�2���uow�Mh�GB��5�䈌<1���&^Eȧj?E3{ma窇���-�<[`i��)�`u�D�
����?mp��kT��X��U��^)�qL�i.
�7�ߗ�K۱�n�y��V"_���C��m���*xɅ�}'������Ƥ-�����U?���9�!֕��"a��鈘鬹��?�\��������q�<6E�����.x�]B���P�&�\A����42�g�1����uik6�l��(n��T�s�Q��_*#5��.L�Ph�u8�Oh��(:�`qz���i�J󓘧L����*����k㚻���ZSz�^|8�c��Z-3N&ku����
y�[
&Kg`��ե	���*g��xH"%/���XC[�*��3�KOEY�&��U �N�s�!7����p�C�t����h)����ouF�x^�F��O�aʑ	Q� (���ΉM��=��a*�1j���chڪ4��R^C��ynf(�~������N��5[�muˠ����4�+����w�ͼ�}�-k0�'���*5-�P���i��Wk�9sP���?�6��C�]/ �Q�(9�^�	����Z��U0_�`>K�XXd���%�.@S�i�����lJڻ���rytȜ��&$�"�ti�IT�v���c������UD��I.�)���>��"d��+�jcw���]�����U2@�/��Ķ!���L� �$�֝U�`&��o�`Rv)-_A0N�O\7hcY�?L{�']��^��Z�AIM�B�5l�e�r��(�����W���'�qi>)�H�r�9[�ſ�����ۀ})=�(f��Чy�K��<O���5 ��3g�*qG��Ýj���0��oIGKv�}�g=@]�ݰ�@b�-������>�< ���l���G8�U��1'�6v�i�����2�:͙)T��â���B�c�˴
 O\0�ĉK\�j6�/;5I�Cb��]�`vd+l�^��FU�wg�\�CLؘ����
�b�_j���yc���s�yXW�M��ݛd��zf����
�"��9'in�V�����zs�����kൣY3��Ӗ4�^�{-�j:��	�>gc<�c�]��<����������3���"RJ�o������'�K�5�E�0C$�❥�I�{�T��W�,zqE��Ee�yl��V���кُ��*�Y�p���652�	.��a�p22��<l?�c����\|f7����������
$g���^��nR�����7s�?����W�.�7���#�~a�x��G�]��7����Z+v�i�y�>𵭹�!FV��k�T9�K�&7ӫX;��~,Ⱦ��8�h�O��N��k�q��U��/������wE,�J���ڳ#&�#-Ո�:ڻ�f{d~;l�}5���[�_����V�ʥ�n����m� ����4W�hƓ����s�,��~��J�5?�i#O��&���_6ʘ�[lF',�&�!YxÃp}���EK�:z�G�^�+90����P0uƜK9#�T��3��S(����thI���w�gFs)9l�V{�K[�P��K�)p�CX�����+Ï?�4h j;&8 ����8��"&�'�+o�9f\�>O�-GV}.C'kc%	�}Z�Q��Щ�P�����'�Ηq��������2#�ce�F�L����A�O�	e�>$:�_��6KLye�N����;������S��|�~e ���9\�ƒ��D'�5��79�`�gq�h����s=�W⛋�y'ތ{��'�8�@
�ߖ�B1�'��e�M�Y�@܇���׶j4����K���q �Z��#��xƠf?���N��bm�ZJ�n�Y^T�����P]�O�H8B������$q*	w�#8��B��5��bL�YU�.LYki��	�P�<�ߧy[�V)�����i{Tp��?�~Z���B��Wl��JC�n�P`��HH��.,R3Y*�	m���.�����2�_�v
����(R�{�!�T`�.�*p��װ�dVͅ��d�̍4R���e�u>}��I~bo0�������g�eh�(��`&��`��Dp'�Ȃ9Z��m����>3;�v�͛��Dy�5�x@��󻂶>����O���'p�/P�jr���ږ��\������.z�����
 ,�X���F���j��g'��-ܮ�Ρ����򤌦 <ki~f�V"XD�Z0�uA<i�X#�����z�3�����#L�$��!L��sZ�&�4IW+d!w�/aW�Ĩ�𵘇�]`���{�Q:rh�O.��bT�K��ڭ�Ϸ��7��v=�ׄ7�'8¸=ң勮``��b�*_���:!Aّ)y�H��d���-jB�؈���%x�{�p��㔿�?�f?8�K5�1%�".�@���$��[��/յC/a	��BpͿ�������9�FF���_O��mc�wH�FdI9�u���}�͡M�Z���"�(�byo�Iy~VjEGiE�=�7ݧ�P��{ B9���>��۰Sҡ'��,�.�>�c,У>dz�3�GQOtF��Д:p�6w.�5����C.:���cWg�� ~#�)P	\ŷ(��;W��Y]�;����
��0�tQM�j���H�����F��D���R�#�pӛ-����̩ZU�<�|���6�ǩ�kCFz�����!~/�B�r)[�j!���e���$�x�Z�٣��O��*�/;����Vf�V`�,<�t��O��R���k��;}�'-��)�ą�ڣo,�|Ȥ��(S���qUtN1�a6�r��ƺ�n4�O�����!bv�`q��"���&�=|��bHá����{�&/ܓ��ϝ$Cу��&i�W�ހ�����A�B1:�Ju-41S��"��\�svh=zc�g2cH�o�ENP���'Ȟ+�֟�W�'eMG�;��So�N�1a'��H��~Ro-vw]E>J�����1���ê�2krw"8�U��H�h� �ڮ��U�C}�%�Tɭ�I� ,9����$�0�#�T�����,E��!!�R�_g16/�� �|�+W�un��!�(DE��O�f��o�r%�)�+rfߨ���"\&ک�*`�����Q�_d��Z	�{B�|=�v|g��FO�C���4w`7����ҫ��N�N��u�z�D�KV�pU��M"�����:�#eUV\��3g3%��	-"�#/�U����/���ڜ�2!~���\�?uP���E%&WK5M��no�}ݎItR�6Y�q�ħ{���?���ݘ~�p�O�ћrV�{�lp������+(?��F΀�ZQ׹�۲"��^�폛�R��O��]�引=��^-X�)nI����߄B��j/�Ц8e~&'HF��"��F�bVi�wx�b�%����*ñ¾A[���#�GLh�/��@�to@�`�h�U��,p�Z-��R�]��GiL�@W�8�N
��]%տ0���P3�>=NG[���*��h��z���a���/�sBE�ĥ[&$����NJ�I��컗�䫍B�Ѓ��;��X���EG�ɻ]_����֔8Nx�H�U��ZV`��e�K���%HA��?��),�������g�c�T2(��G�y��_Xu���U �Ͽ	��ē_B�{#�3�N&1B����ouN]OMe�5��>���Dm��߃����5�/�4�'���P2���GHZ7ފlf�P�|7b�;0N|���5<�<�E���$�oU�^,l�� ��z�&��(�ϳ0�q�en8�����Ch	�&$������9"s��{���f%o��趨f�(+X{�!�*��T���t�uz�bzy,(��;U�U���PO��H_�,��T�2��'M�F�M�k����Y�Od�Bv3��<��Ke�a�$;o.K��aH���Khe*a���^����y~���ѻ"��\��X�G�	��ب��EZ���"���Gd-2L�j9��Gn�~�A����F�n��P�pa2]��F�Ȕ2/�al�~W����EfE��Ἅ��!�����$I�쓖9���sRrd����bG,:)�Lˣ�J{��lYC	�R�p�O;���i~Ɣk�<c�HKzl_�"b�>�w��Zt#�<뷺�{t ��r�.���uR���L�&�f�A[iSQ���m�a�4o�~��Kk�zy�,��+.��$gE�����r�Ph��n=^(�M�ʶ� �[�I��t!��W�w��tVѽ��K�l�	���]����)E��0������H-zʞ��˥�P�2��"~�O�c���P�~���賱2�)�2�\8i�<�9怅��vE	��ؙٜ�f�D��_y���Joˁ�f�v�:��q�6*8���?�;��U�<�VMs���Ҡss��A��a)TUwMl,b��/o��Ы�ٜI�&1��Q𭖦������u�C������|�̖7PB*')�)�]j/��/N�u���h�Q*�7Tq��U�)k��u}���4o�
#[RIb���
���p��2����{I�-S�i~%k��ܖh��<d%S>å�-*�"�d����DN�GK\�`Z�Y�^��/v���U���O�G��nP��|]m��8�v�C�Pٝ:^�{�q�z8�C��\���R�7�� H�-����dHo���s����1��Y8��=��$�p\xG}sC���6�