��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c\�esR&{������o�T�e�Z�/��`%�����1�2��g\D"[ޏ�F�
܌�)�u�lg�h���T�Rfz��9�x��+�E���6�e]��@��<�9�Kb�[JYh��<�"{��Xw~�ti��ZS��{�(1�|T��]F��R����x�f���w���%,n�uG=�@m������+g�#�4�n����n�z-���:bp���%Zx]�_�rqi�Qh�M��jIS���%�(���4�҆E����Ù��p��8�^���Nۿv�_�𭟥Y����A��zxN%Uc�Iԫ౐����.f0]4>�d��!����<�9,�H�8���oe�Q/4�[Z�����g2y��� ��'�S��3�>kڻ��\��h4XeR�uGVCRZ�|��ƒe��F�lEH%2�m^��Pbڻ�N=5��F�����In:�Tƥ��65��c�f�N�u�z�%�`�]��ُJc�xi��?k�����(E͍gHcH��]����0
�"$N��u2
����6d(����<�Þ�E7~t�e��A|~PXV`���[�}g����P�my�BpP�Ē��г\J|�0}xi_5C��L��M�a4�ס�|�QlFzD�2��*[����x�O^L�m+�3$y=��P8�Ւ~����Aj<��l���K}�%N����L\.7~6�!bn�<�5��V�Xհ�����9���_��h�Ŗͷ(��.V`���L�ļ�.�Cb�X �RE�޷�	�7�:���YV�]�d¡���n7���ˈq��!1L	S�ܧ35k>Q�wV�_KW��I�,��CZ�)~#�'��s/��L��^��c49-��F(�ԗ|���A��fx����Zݗ��f�Ktv��̂ea��i�(t���<:����T�X�z�F�1|
�l,h���5�<�lv��Ն�� Z)�Iq�>[Y��7-$��7PD��?��M��ǉ���n__��E�^��G�'�r�W\��t�G���Ӳ"`�\��8߷h�����G�+�6�=э��]��y&F��ehiJ���P^�~�z�l=)ޞh�a�1��qF�����i����"�l����Ac$ў�O��[B�d8�3_ ��&K4;u�ҋ&5� �
��A^š/����S�m�xd�o�v�`�$����9���y�7�g�-s�/F�#��z֩Y�
�W��Ȯ�~'���~�ߒ��B\<l��/M�fhe4�69�S5���p����@E�(��|���8U��������8��a��A۶��C>fw49��_��c�:ؓQ'�˩�ܡI���ܨu/�}��-�+%�i\�BİސY&�)��e�9��dz�m��b�jXeJB8���Vv�~8]#U�&�h�-+����t�qye��K�h����@�;K�޸�5'�.)��;�p�y]��
�퓦��i�Ǹ�[���-�S����|p���;+�3nE��ۣ�~�^����`c.A˔Qs� �;yW�s��q>*�Z6��	5�Fɠ�����v ��K'�CB�����̄F[u��Ð.�*���� �s����d]��D6

��-�~o�g�:�Kё˂�L2�t,hl��7'�������^�@ڄ�
���n)CeM5ihZ��(���c��Qg�GI��Vi�6�FP�BU�jZbPѷ�]ډ���l{�z{��&�JQ��XS[Cac��\��+��!���.ʝo-�yS�(�8�j��ߚ��Q����n߼���(j��͹�nå�(Zh���idWoE�*��{^�	�K�����c�i�$F�>��cJ˯��Y�"��3)��W�c)��f
ۈ����]�S �����_70K~m� [��6� �nh��gb+�#:\��d�ϔ���[�-��u�A�E6����w�<��-�%��n����@���J���mtW�zxVy�@�YP'�(e���}��?ޟ�o@���y�R��-�ˡ��_k� �M��r��eq'�0�O�}���Tir�߅�Z���KVg��KRp�"���F��Y-�5"�Dd��̵:[ 5P�[^В�dh��'���C�~�D��ևmmc#h�������`�^?�T��Af����5c��q��Mb��D"�] ;/ו��l n:�w��b�ϐO6�9��#��/��xת��Hդ�Q�ʲ���6�,,H�_7��t`��h<��N�4��T�6�V���~�u��y�=��y�g�R�Kc�����fb�f7}��I}.����kˊY���
��d��OW�A��rt��k��]uN����i��^ֳ(����|H����6���|�ݪy���h���GSw2�ԟ��}����P�!�O��M����5E��Sw���X�B(hnbƋ΀��6��
/���SP-w�A�1��v�]q�C�����7?�Mȵ��b�j���&]�dBh4��x=�؆.����x@FR�أ~2�A�V���'�L-D5�-RK�x�H�2EΣ�o&T_&|[�2��O�����>2ك���Or#��:lh@5p{Cf8�D��\��}��6z�R�����`�C�P�,?�f4+�t�O�|B�*���K�m-1�mBmW��pj�z*��01�k�
�>ب~F��ي\�P^sE�D3N��X[O2�B�r�a��/0H�OB�X+u#!��rͥ�N���@�W%� fGil�O<�yzda9��Cpn������;)4����G�Z ���V�] ��@h⬋8!�O�'�	���-�mtu}0o���"�m��px�ҵ�TS?���(Qd�����q�)/Q\?-����"��՛�dM.Z�Oْ�����OvJ$�9(�'_73T2*�&��^]��v�&`V}DHa�e]}f"��	5�ڬ͗����XDB|i:��|��(2}!�j���J2� ��Nܓ�<��R����Z�g^���m��	�x��[��[�L��Xp#$��b�R���&D����>s/�D�LZ_U��f���,�
]⦞�ι����vW.u�R!P8�Ġ:فYFH�S^� .�ݧ�O���+q0����j�	�;>z���K�-��0+�=�mྒྷ�w���=~�Si?n���.=��ͽA�Y6Gn9�/��t�6<cX��|)8�ql��;�~R���{��"�]*}�"�s݃(�+>|G���ǵ��4�Bٺt1y��U��{S-�4H�d�Q&���WO���F?`roy����"�	gH�s�LCG������zO
��*����k������03�דR؊3��Q����W�m����[�D[�w�����Y�`e�c^�i4����E{8ut���  ʹ�VL|�y��չ7p:�a�Ƙ����Ϸ�&�JyM�B~ȤRZ����o�}g��f�ΘkԼ,��#������@��3{�8"��a����i�Z���%v펍�L���u�
Q3�t����2e*��)K�E�W6gT�ۨԓ�eOI�p�!��J�ĕ��L��Rw�O9՜]�g�k�O�7:�Ax�:C ��!�^\P��'�Uy�b��s%�z#�h!s���jq-$+PM�]�q{Mo~ItY.ص���ˁa�O?M��Ҕ��p�v퍩x��g��1U�Y����KV�ؖ�S�<N*�7!k W;Fb"K�^j��f�nH�wߠ;�Q����>�C��ۡ�0,�?ɉKz^#��/J$�/�pm���a���x�1@!S�� ��|#qY��+��N6(���5��� ���vF��4���7��4���9�ae-�`GqFHDژ��(ه&pÈ*�!>.v쨗�#AJup���o�4�:��~ �mKP�RQ��W~�B3��@P����|V+��&�N�L���Y�o�p��_�u����#�(��D�;""��7 @<�����90�ýi���wB�k]JVC�a;�_��j��(��3\:ʮs����.r��ϙ��m��me��Z�M���:U��0>7$�E��9!s�B�a�,4�W'�bY��o�a7q���̓�*����t���t�*GQB�YRr ��]S߮b�\a�8"����ckq��w�p�=�;����1�p
�8ZC͏7�g3f׼������0� �sFi�(~�t1Eϙ^-*\KH�ʠ�#�.\2z�������	K� \ӟ"0��-��H��:4]c~%�
���[|$h�����-?�!+F! N3/�~�fG��lW���Ğ^R��:<\%��\\���Lο;/o�g����v�d���obn��c)E�Y����肹���'D�
U��R3x%Ra�m��/?7���������d�*��L��na�S��.<���mf�g���Mk�M���M�of��[�t`��	��ex4C�����p��q�V���jO���ٹr{,)��R�����!:!�SaN��x�<�T�A�b����("���,��چZ�m[���xV�[�8�a���#m�(�0��eq��nQܧ��/�c��	G�,�v���:���-xM�5ת(��!����
�7_s��(z��5���)�ھg��Z�|�W�ہ��>��N0�F5ɁJ�(VJ���M-/_}�E����vbI�����n���������x-�pi���R�[���|U� zҀ��3;!y���eG��ຜ~�Mu�U��@_`A�t�N�@�O� �s@f�juuD��v�������)��45����c(mA��������v�6q�X��8G6cQ<9	jv� �|�!B�-�������;j�����"��o^*a�$�mn� nWk,j�gB۟���p|�^�$�@�K����]���J(�cj��F8���P�Z�����PB��?�q�_��	m��:��q@M@��c�������N?����)�[�5�|l�T�I���;������9���战A�ut�+1xʳ�z�8�Ӯ@�?��5`���Kك)SV���`��c��@�1;	\�|��j`҄�����iB.����� ���!��tZ�UBq���9B �n�J4��8	�<�t�K�q%�]g��p�e��Sf��g�0��7����c���e���;ޙOV��e�é��<�1�!�!✤�E��&��q��Wh��A3[Nk��.�]3�pX�Z�0����hRF�8?����HUv>���ѵ��2aA��ͳu��	�(�}MJ2�n��¢�GH)���6��c�[;�Ͼ��D����u��|�^��D�!�� y����6����ԣ���+�#�I�<��~�����U ����iv���:�*�s��s�&�B<y�2bc4*��7���Y��Xe�@�=�[薡�x56�j�h�i���W��I�A�IZ�xO&��ų�5���:Uuk�	�rXB&6� x�G'JḾC���E}Г����w���Y���d1?=S��:�r)ź���"���WY��$��e?��Ԫ��S����yF,��7P	�*�;r
� �cOV;��B�^��7?
��{( �Gc��s�s)���Q���E��#�K/k���F4[��b�'���U9,U�_�a�s�ªo��0�f���Dj\Su�8�?� �F���tr;���s�iR�=f]V�{W�x[�09��p����j��uނ�&��Yt�۵� g��O��<Ĭ���Sqw�O9Dg�N	�e;m�p�t�e���J�g��Y��wˢ�7O�B�rR�0��L#;�����a'�?X�F��a~k&X{�[�㊞�0^:	������k9H�b|"���S�R����;ɬ��G�r�L.������q8^w@���W6����T�o�-�t�c����Q�A����~P<<����K��k�'���Mw�0?��Cj�X�&շ�9�,��⣬4a:=����vS�j�s.��b;�4�hҏ�m�j��m�"��(��Ʀ?ı�T��E���$û��jƌzO4��{�m�ջ�O툅�"m͑�JE<6����s�R�ȼ]�'p�!��>��L�M�!p��������+*Zv��Ԙ<�	
�����2��9��t�l{щR��l��y,�iJ����q|�H���O�5����0.7�	g:��x[\��֌�>k�Ne���[�����ZT��\ʘ�D�I���%o䶧�ڴ<@����w��J���I�������<ur�U��b&t:�ymz����s�N,KV�/
��XRU�@���5m �yoWyzN�O�^���/0�ؙ�e�,٫]8V� =�5�[C8�G�Zo4�2�@��R��PďV����Lj�9�{
���)�
�pE�RE{��ޱ��{/�I���m8&���i�N�H�;\�`��Jq͌�e���9�[�5���z�`=�������q=�����6�~9��T�0K������� @���e�!'9�7�+�G��ӛ����\9L}���*���+��^�<�ӌcy�Į�wT��W���EW`�Ş
tח㢍Jߟ�g�R�t��E*�2����	�I$�#`�������e��z멮�*3��`����Qf� /B�rbö[�ߓST�h�)������SR�;�hs%�Pv�e:Ltg�\��p�e� >��\�=�_Tn)�	�L�Ѵ6)��7���P|�9�'�����.w9�������ܗ_B?�Yg/yס��|G��L/���zr+q�W�0㺷�+�$���4�xD���؛�φ.mU�)����Ws�{y��b[RW��̛m0z2?�8N���74Of�j*::�.�*z0h�d��m&��]�9�D}C�O:�0��[��
w+	zւG8����9���g�,(������������|�iK��c=��3<�U������h:�q�w1\m$�٢�1E����f�����u~���> WUPsEi~�!�.��5�	���)u�XuW��;%s�8��aH�������Q��׍CN~��ByFXM�2<;�|��t�Jk,�y��٧1v(�#B#���5�����\�eK���*1���Ӟ�$���ݷ��F��*3�Y�����M�Cz[p�ӧ�NA��ԏp��M�"�#f��}��+��T瘪9��y�u��
���X��X�38E#Y�4mI�����4��6ns�c��%�.z���Hg25c0��$ĥ�/?��i)�N��_t#���ps��|Z��D� T�ʈD�<t�_>Ch�	�EWm+���j䯨���o9�4���XK����Χ�=��1�����z�ڈ�����Z�7�5F_��Sf����sk���R�G�A{��<Je��l����I/ ��$�M����ER	�1�QƁf�X�Y�7�6�<��gEJ�D������_��aikz+�E��pj�&��hk�	��F�l�~%+�����&��G0�m������a`��3k�O�v`���y[@�4��{� ��==��^�@1���.I��a�ƹ�#��<��=*��դ��o�=��^[Q'i��&����7uJZSC��1`�Ku��6y�	H�:~�tS�;��ұ������������&�&U�5�,�a��1��I�ݙ� C���B�%�R�Y�ءB{�aժ�|���9V�O8��$V��a��3�V!r`��^�������0e����i�Q�2݄C�c�{]�{p9�`M�^)+oNcl����c���c{��/�U ���$�~��s�֦p�6b t1x�4	�)�Z�7�x�qzx5�������v�T���j��ZM�c2���U�N;��[����(��b:c$�����;�EN&.�j�?����Xh���g��^�a{g@�F^�@� �41|U)��W��x�.x^%�\�,k��a&|t��Sڿ�B�s��SvP�þ���
h�QMȮ���)1�����=��c���r!�*��W)Z2�05���L	嗘� �r��E�k�mT��A�"�!+L��͢���{eZa���[L��%�� ��׀Q1#�(�2�:Czg0�5�r��{*������b�ʄh Δ��ϝl4��7�,�6���^���V���߰�6]���I����Ư�<�[V�9B/���0Z7�'/�	.k�u�����a����;�?M�q���ɔ���1�x�ܙ
[l�C��yͷ-�Lљ���4���J�\c���箮�wO�I{K�`����K��lc�D�� n��vtC��-�y~����`��~�"�3t:i:��v���������3����ƚd��v3{�OG�o�-d���+N^��>���&~\HV'͜�?�53�Ƕ�z��Q��s>�-���K�BdkEL~��g�__X3��P��RV�z��Q��zPڦn� =��l8{�S�u`.=�(o��Б���~Q2�C�_C���T�����{���=@�ƾ��'��b2\\�^0Ό�IJ�a�eb�5�@WG*�������0�S}�����[��Ȁ���J����Vl�a#���Sx5�K�^���Q��ZB����{��Y�`͍xf���j��>��B��"
�m��c����f���~��HJ�������	����I�=�F��s�2��KVD�q�S��/#��� e������p�氪�lPLCy@3x�C�L��QD	ʝO,t����:K ÝQ~�Wz9������C*��cCSzVh<ir�?�� ܦ�)2ކ�F�N3_���̟fܽ0��>�9A�V��P�:ш�9�V��_�Kq�WV�P�H���`S�$S�*�*��/�� �,&�f���b�%bL���ڸ��ae�]M4T��H��=wĨ�󚑧}Za��H�p��qQ����Z^�E�a>ٯ�e���>��s��FF!Wq���7F�����[���>�x��Lb��ƕ���i��>�&��-m�_�5J\T,�ZVP�M�_p�@`_"��ֻ)j�{\���� �âM��E��� �s� ���M��Lf�,C�&�ޠ/�
	
��*c���6�_��/�+�S�tL�C^ru�d��sb�^���]:��A���+�9XP�^ޔ��k��'�6�j���BN�(���m�d�W#�>�W����ߌt [U$��<��rƝ~�a�L�2��V��`���vضy�{M�Q{�^�_����TƤ�����I�lky#�"�y��x�b$Y�G�Nu^DpɆ��h�s:��?�k�uh!�ONNڬ;a���I�8{�i�7��F�7f��'_lE+C������Uz��9:�0�A2��dc�ozb�q�̕T�>p덣�cw+���X|�QT�'�q�@�Q���3e-�_�h���|[>!V���@��t������c�C��$�P��.�l�ca��lrS�{�ţ!�A@���I���~_gܥ�z��}kٌ�z�\�a�]���E�Y����t҇f��$ۣ�����
����؅����ie�3t>?���� ��~M:��6����	��\U���}��Q2���R�D�����V�#iBY�K�k�Q���5 �e&I��b��k-wУDuGmB��~ 5%U7���U1��d��^IES�W=�J�R��9z0�=�7u~��|BK9�TwjB��yV?�M=FdA���¢Oae[� �� ��%8�����%�0�9@܊j�
=݊��*C�J�9��@�X(�7'��}~4�E�ȡ*-�&��yt����EƍsĤ�i���+��k��Ü0,E�dzv�@X����}�;-�.�t��~o[9˂����.�R�H׿�A�;�����B
c�_�$d�!�=z��5$t���#Ѻu�H)�5:���ѭC4c���-@�����(�Ԇx�mI���k��h#G�6%Q��w�����~�L��NZ���!M����S�%�_��w�CQ��7��Y�j�2b&P�yr��6a�	UB��Ԁ�`���@*~�OA��(o�.b���p*�><���+�`�Fu"��#pۻ\c$�=��p��7@o�Aѩ��^ F�:��ml�+7���ƜH�}���PL��u_ÌsLQE��� @{8*�n��<�6D���"NH��5x>����[7Y���l<�4����!��ս�~�O�G�*�伶�z�n n��⅘J,�������>��o�}Ȓ��4�g�{/5�]i���z}��e��g�L��'��]��'�
��� ��zj%bӪ37��=�tq	m���a�
�ʓK�;꘱1/�Ӧ7��'�|AFE��p�౼O}�?�>�A�8�;����9C�ɊD��e��y upcM��%V����|�n��USt�A���ј���n�i��(��#��汹́�o����+`��=��8'��KC���2�(��v�(��O��U�RXic�~���xx��� �
i���
���=.�0tK��@�J��PZ�h,��$9z�R�[b	z`��t�&�x��4P��QS�ܳ�ȳ�ΘÆ���`R%���W��l��É�q�xɄ{�����-�g���K��b��u4�I5^��}��T�@��[�qK�c������
�h��		_	��xޓ��H���?bQ��v��]�x]��	WqV��3�q�7LU�/��WnPsn/q�d�
	�Y�r���VerNYY�m�(]o����J�e�@-+�[�Da�ԫ)���BK�j8B��On�< |����Z'��=G)p�f�e֘�����z�	�G#�X�����)���g�ۍ-���2�e�.�i�ƅ�G�h��E)�)��w���4�~���d>;.#�2��@2�&�C~���A�q��ǆ�6h���p?�
��v�+J˔�g1�k~嚟�7�C
�ؙp�5SC 5���z��\Y�e� =�(�����\�i�����ơ^BU_��Y���>JNR�f�Xe�̎V����]
��R>.�߾gn&}�*��q�k�
�r���*x�NQݎ��\��R������=a'�@Y�'U�����S�r�߻�	�oC�w�[������`Xb���=q?(ݰ���^PB��\p+����ܹS	��ψI5�q�=>�[��%��6y!-%
�]Ӻ�[a~�ݸWI#�:KG-���P=�ޟ�!�t���k���G-�Fi�M����f��y��y�*t��<Clc ��n&�n�բ�pƌ�`��b��r:����-��(r{j�R�Ͻ��ɀE�S
PK�o)�.80-��@��CŞX�d�:�_5jB�x���Š��%�us'��aPQ���X$��f��n��Υ��R�Z�c���sUb��nrr<?R'�%1"���Q��Y��罷�*>�-$?^p�Ƅ�v�ʁ׻�U�
�Ѳ#��?�-��7�8��u��+"r�V�L�_�roI��f�)$Єqb�2I��"�i6Y���5.�U�٦0^�S�6y�*p+�����&r�g,n���C/?�?�z,�t���Y�F�U�����E0����4�Xѷ���IhN��]��C�2��֘�V��9@Ī*/�����GC}�xT���m��{�T7���5K{]$��񽳀�����PS�cq��.�CY�[��y��ko������5&Y��zi-�v(��ֽt3�ƒU�&���}��ych�I���&�'�f�E&%�'!�2�m�h�JHִ����M�BGP�̡����z.1j=c�Z۪)���!H;g�������1v _��-^�ʟ�w�������c�d�մ_&�l��uʥ7�j{��O�j������޿��&b��kTP�f)Z��K�	�r���s�)��|��Ȝ�ߜ�0"*�ܭ��<�<$�L��ɰ5˫����p��)4y�CW�ʇ�l�pNE9��n� $�)o��=���B+�t�H�Bґ� ��21^Vg�;g�Ĵ�[#y$ؼ�#�B���P͚�^��MۍT�], �"K���N�A�r�2���7�Mo��HK����0�]>Wֆ8چn y�-y;�3���x�|��K���"�!M��Ϋ�ВS�!
fWMF`E��H�[�Z�e���UJʻ6GB$>���g�j�Eqs�IP@=�w6:ֶ��k�*J��u�ǺoCɈHJM	����Y� %)_+j�e�$�Ic�z)���osG��Y9�:4Ma���6�?R��xÊ�׍b��~`'����SJR>;�1��D�a����l�'#�����f�b)U6�tH��5����H1B�'M%����
����ҩ��vC�8]x�dL"X������ŊӫV�P��E�4�͖[z�
'�.�NE��f���k�"$(�TAG�S�P�$��@�Ε��Z�JԲ}�5D�2M�J��5�%�{@:Fd�tG}��i XX2�������41��������ʇ�?��b�l��_)���+�@�zw�f"�X�yW��j��$��۶ŮA�*G��Y�Y�({�|M�7��k�=�-N-�,�t���{ZM�r��í�H��K+���
x��3�	,7���s�;�E���"�fI�IɄZ�R�T��g��ehu��y
��0��S�D�ي�?�+�۔���#zq��|.�� p�Z)f�R����KK�א7��-P��cߙ���r^����m�� �f�n�%(X!�YR�}���t�@�	K���3E�<���EI"��ˑb�L^h+���K��K��ek�kE�m\��f:��ώN�K 1̠-�/�p�`O��vK|]�E1�r��.��ޓI5��"#Z�.�T����z)qN�9a/(]�Hp8���9A;���)qQ�5�Ŭ��K�,�t���W�@��t�R7��[�T�KBuH��Wd�Co�*H�t��)��H��b@8p{��d�\�i�3��s21��4/uAw�Ɛ���я`2���y�����WR~��M+`*��aӤi#B�F)in�[W�/?\J	����QY�&fA������B��0����ꗱ�KW8��!�p��7�s�"�;�=o����}b��,���tn74�!���Q�i��q��DIB#�0���¥���'T�S<�/����>��Jܰ����<o��p��[0ʟ]WP*�m �e��[Ό4�MX�:#��;�"T��Z<l.;����
�.�ݬ����:+�p���rJ:r9�r��!P�|C7AA���.�d�oM{La\��u�]Nkq����A��8Ep��n`����B����
m
Z���O��&��'oeal�Y���&?D�?X��#�Mmt�\�&���lꆁ�I`��gi��,���
��ϫwG�\m@��"�W�Sh����a:*C��ˡ�Uu��]�T.�5H΁[�"BWn��z��W��|�D���MI�K�Ig���;N���7H�cY�o�J�ʅ�qY�`k���~�p��s҂��C�n/�̀\��0"�,���M��E咬:I?b��[(e�n�����;��I��⋃J������Gw���~���I�11�^�0H��������&���X�/��6���GuAL�f�n@���o��w�6���|h
�w_�!�qI��%ܺ�m�����AiU� <&�:hr���r��P/{��h��k�P�ˮ9�}'����dnZ��_�^�ݐ����$��E��m�&����}�
"~�hdG�ԏd%�����FK;�XrU��6Vq7��]��le�\�	�=r��48�w 5����e_=�aL�pC���G���b>�^���Xܩ7!�� Z�i��c��Vm��I�ރ��%Q���.���	?�ש�{M�����nV�4,`NW�4Y���%Ea���)=��&p*�s��*������F��-)�/hF�q��1���n�r�X/_��Q�UF����F��2��K��n:�.�ݑ�
�c�v��a��@<�� ꊥ�Y0	9�Y*�*ӂ�����"fZ1"�~m�]'8a k��ST/F�+)�S>`ل焣G��Z��E��+M;��A��u\[�sE�-0�t])�y,	�t1��b7�Cs������1�Ud��8��w�ԛ��B���$TWFA���X0�VaI�r��)�I��� �g�>A���k�C���)EQ�(��H��J���!»e��"_�Z?��v8ǡR0�SbC�Mue��P�=�GeT0곸f�Ֆw�Ҥ��r��n�`:]Kғ�n�pqg}\���H�~<��Q���\�b5��TWҢ��vMo��G6�Xz���E�<��.6י)v��K�/~*��7� "mY�7K�sO��zQ"��#�?�nv�~@������4�+v����Z~�>&T��	s��P���J%I��>*ߗ�"�?{��1+E/�^$+ق��5���[��ҵ�J���W��C���l�2O�
�/M�ɕ�}��;��y��2F5�u�:|B2�\y�M
�,�ɦ���P�[�]y��@�-�����* 7���tdPN7kӭ5/�����{�p��[V�a9��WmQ�}��A����-��|�zL���P��TO��N�_��e��C,
����otVv�3f�z�x�٦=�A��BP����p$�X���
e6�bl�u"t�*�\�g�CT�
�w�M��TL�à����m?�.i�i���~���s�*�q�_�k�뇃3���/'��]D0ƴ��A�Ew.���4Qʣ��*ncGQ�9��.��t�H' :S9�W.i��C���"(0�y�� �(W��3P��aɗ�"��b�pA��� �z/�A1�:O���-)�k��B�}ʛP\AZ�c�j�».?�ۗ'���o�.�ҝ3J�$#��a?��B��	q�~��g��Q{{��V��}!�'��F�$�a�a� z3A�R>}������d�˟�y�"�$���.����3R��*��MG+b��EF��7Ը"u
8��ߤ^� ���_�`y�qY
6��'ϭQ)��� �'�˕�#�+]P�8"��1��󌻅��i8�?�Av���s��K�#� p{�������hM����O�e��8g7V�KLB #�K�o����`����d��q�ȑZ����V�8a�NȀc��|�)H#𘆵]\G�����@x�9W��RU��آl�f#0���Q���#��yk��G�'���W��NY�q�inP�,u<�%�o��ѩwq��QKh��&��p{$O=n�ܐB�4�/��!����tA��;G���+?(P���G�p� ��X��匍��o/��`"���L^�O%�EX!