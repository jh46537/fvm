// ntv_serdes_2ln.v

// Generated using ACDS version 13.0 153 at 2013.05.02.12:00:12

`timescale 1 ps / 1 ps
module ntv_serdes_2ln (
		input  wire [1:0]   pll_powerdown,      //      pll_powerdown.pll_powerdown
		input  wire [1:0]   tx_analogreset,     //     tx_analogreset.tx_analogreset
		input  wire [1:0]   tx_digitalreset,    //    tx_digitalreset.tx_digitalreset
		input  wire [0:0]   tx_pll_refclk,      //      tx_pll_refclk.tx_pll_refclk
		output wire [1:0]   tx_serial_data,     //     tx_serial_data.tx_serial_data
		output wire [1:0]   pll_locked,         //         pll_locked.pll_locked
		input  wire [1:0]   rx_analogreset,     //     rx_analogreset.rx_analogreset
		input  wire [1:0]   rx_digitalreset,    //    rx_digitalreset.rx_digitalreset
		input  wire [0:0]   rx_cdr_refclk,      //      rx_cdr_refclk.rx_cdr_refclk
		output wire [1:0]   rx_pma_clkout,      //      rx_pma_clkout.rx_pma_clkout
		input  wire [1:0]   rx_serial_data,     //     rx_serial_data.rx_serial_data
		input  wire [1:0]   rx_clkslip,         //         rx_clkslip.rx_clkslip
		input  wire [1:0]   rx_set_locktodata,  //  rx_set_locktodata.rx_set_locktodata
		input  wire [1:0]   rx_set_locktoref,   //   rx_set_locktoref.rx_set_locktoref
		output wire [1:0]   rx_is_lockedtoref,  //  rx_is_lockedtoref.rx_is_lockedtoref
		output wire [1:0]   rx_is_lockedtodata, // rx_is_lockedtodata.rx_is_lockedtodata
		input  wire [1:0]   rx_seriallpbken,    //    rx_seriallpbken.rx_seriallpbken
		input  wire [127:0] tx_parallel_data,   //   tx_parallel_data.tx_parallel_data
		output wire [127:0] rx_parallel_data,   //   rx_parallel_data.rx_parallel_data
		input  wire [1:0]   tx_10g_coreclkin,   //   tx_10g_coreclkin.tx_10g_coreclkin
		input  wire [1:0]   rx_10g_coreclkin,   //   rx_10g_coreclkin.rx_10g_coreclkin
		output wire [1:0]   tx_10g_clkout,      //      tx_10g_clkout.tx_10g_clkout
		output wire [1:0]   rx_10g_clkout,      //      rx_10g_clkout.rx_10g_clkout
		input  wire [17:0]  tx_10g_control,     //     tx_10g_control.tx_10g_control
		output wire [19:0]  rx_10g_control,     //     rx_10g_control.rx_10g_control
		input  wire [1:0]   tx_10g_data_valid,  //  tx_10g_data_valid.tx_10g_data_valid
		output wire [1:0]   tx_10g_fifo_full,   //   tx_10g_fifo_full.tx_10g_fifo_full
		output wire [1:0]   tx_10g_fifo_pfull,  //  tx_10g_fifo_pfull.tx_10g_fifo_pfull
		output wire [1:0]   tx_10g_fifo_empty,  //  tx_10g_fifo_empty.tx_10g_fifo_empty
		output wire [1:0]   tx_10g_fifo_pempty, // tx_10g_fifo_pempty.tx_10g_fifo_pempty
		input  wire [1:0]   rx_10g_fifo_rd_en,  //  rx_10g_fifo_rd_en.rx_10g_fifo_rd_en
		output wire [1:0]   rx_10g_data_valid,  //  rx_10g_data_valid.rx_10g_data_valid
		output wire [1:0]   rx_10g_fifo_full,   //   rx_10g_fifo_full.rx_10g_fifo_full
		output wire [1:0]   rx_10g_fifo_pfull,  //  rx_10g_fifo_pfull.rx_10g_fifo_pfull
		output wire [1:0]   rx_10g_fifo_empty,  //  rx_10g_fifo_empty.rx_10g_fifo_empty
		output wire [1:0]   rx_10g_fifo_pempty, // rx_10g_fifo_pempty.rx_10g_fifo_pempty
		input  wire [1:0]   rx_10g_bitslip,     //     rx_10g_bitslip.rx_10g_bitslip
		output wire [1:0]   tx_cal_busy,        //        tx_cal_busy.tx_cal_busy
		output wire [1:0]   rx_cal_busy,        //        rx_cal_busy.rx_cal_busy
		input  wire [279:0] reconfig_to_xcvr,   //   reconfig_to_xcvr.reconfig_to_xcvr
		output wire [183:0] reconfig_from_xcvr  // reconfig_from_xcvr.reconfig_from_xcvr
	);

	altera_xcvr_native_sv #(
		.tx_enable                       (1),
		.rx_enable                       (1),
		.enable_std                      (0),
		.enable_teng                     (1),
		.data_path_select                ("10G"),
		.channels                        (2),
		.bonded_mode                     ("non_bonded"),
		.data_rate                       ("2500 Mbps"),
		.pma_width                       (40),
		.tx_pma_clk_div                  (1),
		.tx_pma_txdetectrx_ctrl          (0),
		.pll_reconfig_enable             (0),
		.pll_external_enable             (0),
		.pll_data_rate                   ("2500 Mbps"),
		.pll_type                        ("ATX"),
		.pll_network_select              ("x1"),
		.plls                            (1),
		.pll_select                      (0),
		.pll_refclk_cnt                  (1),
		.pll_refclk_select               ("0"),
		.pll_refclk_freq                 ("625.0 MHz"),
		.pll_feedback_path               ("internal"),
		.cdr_reconfig_enable             (0),
		.cdr_refclk_cnt                  (1),
		.cdr_refclk_select               (0),
		.cdr_refclk_freq                 ("625.0 MHz"),
		.rx_ppm_detect_threshold         ("1000"),
		.rx_clkslip_enable               (1),
		.std_protocol_hint               ("basic"),
		.std_pcs_pma_width               (10),
		.std_low_latency_bypass_enable   (0),
		.std_tx_pcfifo_mode              ("low_latency"),
		.std_rx_pcfifo_mode              ("low_latency"),
		.std_rx_byte_order_enable        (0),
		.std_rx_byte_order_mode          ("manual"),
		.std_rx_byte_order_width         (10),
		.std_rx_byte_order_symbol_count  (1),
		.std_rx_byte_order_pattern       ("0"),
		.std_rx_byte_order_pad           ("0"),
		.std_tx_byte_ser_enable          (0),
		.std_rx_byte_deser_enable        (0),
		.std_tx_8b10b_enable             (0),
		.std_tx_8b10b_disp_ctrl_enable   (0),
		.std_rx_8b10b_enable             (0),
		.std_rx_rmfifo_enable            (0),
		.std_rx_rmfifo_pattern_p         ("00000"),
		.std_rx_rmfifo_pattern_n         ("00000"),
		.std_tx_bitslip_enable           (0),
		.std_rx_word_aligner_mode        ("bit_slip"),
		.std_rx_word_aligner_pattern_len (7),
		.std_rx_word_aligner_pattern     ("0000000000"),
		.std_rx_word_aligner_rknumber    (3),
		.std_rx_word_aligner_renumber    (3),
		.std_rx_word_aligner_rgnumber    (3),
		.std_rx_run_length_val           (31),
		.std_tx_bitrev_enable            (0),
		.std_rx_bitrev_enable            (0),
		.std_rx_byterev_enable           (0),
		.std_tx_polinv_enable            (0),
		.std_rx_polinv_enable            (0),
		.teng_protocol_hint              ("basic"),
		.teng_pcs_pma_width              (40),
		.teng_pld_pcs_width              (66),
		.teng_txfifo_mode                ("phase_comp"),
		.teng_txfifo_full                (31),
		.teng_txfifo_empty               (0),
		.teng_txfifo_pfull               (23),
		.teng_txfifo_pempty              (2),
		.teng_rxfifo_mode                ("phase_comp"),
		.teng_rxfifo_full                (31),
		.teng_rxfifo_empty               (0),
		.teng_rxfifo_pfull               (23),
		.teng_rxfifo_pempty              (2),
		.teng_rxfifo_align_del           (0),
		.teng_rxfifo_control_del         (0),
		.teng_tx_frmgen_enable           (0),
		.teng_tx_frmgen_user_length      (2048),
		.teng_tx_frmgen_burst_enable     (0),
		.teng_rx_frmsync_enable          (0),
		.teng_rx_frmsync_user_length     (2048),
		.teng_frmgensync_diag_word       ("6400000000000000"),
		.teng_frmgensync_scrm_word       ("2800000000000000"),
		.teng_frmgensync_skip_word       ("1e1e1e1e1e1e1e1e"),
		.teng_frmgensync_sync_word       ("78f678f678f678f6"),
		.teng_tx_sh_err                  (0),
		.teng_tx_crcgen_enable           (0),
		.teng_rx_crcchk_enable           (0),
		.teng_tx_64b66b_enable           (0),
		.teng_rx_64b66b_enable           (0),
		.teng_tx_scram_enable            (0),
		.teng_tx_scram_user_seed         ("000000000000000"),
		.teng_rx_descram_enable          (0),
		.teng_tx_dispgen_enable          (0),
		.teng_rx_dispchk_enable          (0),
		.teng_rx_blksync_enable          (0),
		.teng_tx_polinv_enable           (0),
		.teng_tx_bitslip_enable          (0),
		.teng_rx_polinv_enable           (0),
		.teng_rx_bitslip_enable          (0)
	) ntv_serdes_2ln_inst (
		.pll_powerdown             (pll_powerdown),                                                                                                                                                         //      pll_powerdown.pll_powerdown
		.tx_analogreset            (tx_analogreset),                                                                                                                                                        //     tx_analogreset.tx_analogreset
		.tx_digitalreset           (tx_digitalreset),                                                                                                                                                       //    tx_digitalreset.tx_digitalreset
		.tx_pll_refclk             (tx_pll_refclk),                                                                                                                                                         //      tx_pll_refclk.tx_pll_refclk
		.tx_serial_data            (tx_serial_data),                                                                                                                                                        //     tx_serial_data.tx_serial_data
		.pll_locked                (pll_locked),                                                                                                                                                            //         pll_locked.pll_locked
		.rx_analogreset            (rx_analogreset),                                                                                                                                                        //     rx_analogreset.rx_analogreset
		.rx_digitalreset           (rx_digitalreset),                                                                                                                                                       //    rx_digitalreset.rx_digitalreset
		.rx_cdr_refclk             (rx_cdr_refclk),                                                                                                                                                         //      rx_cdr_refclk.rx_cdr_refclk
		.rx_pma_clkout             (rx_pma_clkout),                                                                                                                                                         //      rx_pma_clkout.rx_pma_clkout
		.rx_serial_data            (rx_serial_data),                                                                                                                                                        //     rx_serial_data.rx_serial_data
		.rx_clkslip                (rx_clkslip),                                                                                                                                                            //         rx_clkslip.rx_clkslip
		.rx_set_locktodata         (rx_set_locktodata),                                                                                                                                                     //  rx_set_locktodata.rx_set_locktodata
		.rx_set_locktoref          (rx_set_locktoref),                                                                                                                                                      //   rx_set_locktoref.rx_set_locktoref
		.rx_is_lockedtoref         (rx_is_lockedtoref),                                                                                                                                                     //  rx_is_lockedtoref.rx_is_lockedtoref
		.rx_is_lockedtodata        (rx_is_lockedtodata),                                                                                                                                                    // rx_is_lockedtodata.rx_is_lockedtodata
		.rx_seriallpbken           (rx_seriallpbken),                                                                                                                                                       //    rx_seriallpbken.rx_seriallpbken
		.tx_parallel_data          (tx_parallel_data),                                                                                                                                                      //   tx_parallel_data.tx_parallel_data
		.rx_parallel_data          (rx_parallel_data),                                                                                                                                                      //   rx_parallel_data.rx_parallel_data
		.tx_10g_coreclkin          (tx_10g_coreclkin),                                                                                                                                                      //   tx_10g_coreclkin.tx_10g_coreclkin
		.rx_10g_coreclkin          (rx_10g_coreclkin),                                                                                                                                                      //   rx_10g_coreclkin.rx_10g_coreclkin
		.tx_10g_clkout             (tx_10g_clkout),                                                                                                                                                         //      tx_10g_clkout.tx_10g_clkout
		.rx_10g_clkout             (rx_10g_clkout),                                                                                                                                                         //      rx_10g_clkout.rx_10g_clkout
		.tx_10g_control            (tx_10g_control),                                                                                                                                                        //     tx_10g_control.tx_10g_control
		.rx_10g_control            (rx_10g_control),                                                                                                                                                        //     rx_10g_control.rx_10g_control
		.tx_10g_data_valid         (tx_10g_data_valid),                                                                                                                                                     //  tx_10g_data_valid.tx_10g_data_valid
		.tx_10g_fifo_full          (tx_10g_fifo_full),                                                                                                                                                      //   tx_10g_fifo_full.tx_10g_fifo_full
		.tx_10g_fifo_pfull         (tx_10g_fifo_pfull),                                                                                                                                                     //  tx_10g_fifo_pfull.tx_10g_fifo_pfull
		.tx_10g_fifo_empty         (tx_10g_fifo_empty),                                                                                                                                                     //  tx_10g_fifo_empty.tx_10g_fifo_empty
		.tx_10g_fifo_pempty        (tx_10g_fifo_pempty),                                                                                                                                                    // tx_10g_fifo_pempty.tx_10g_fifo_pempty
		.rx_10g_fifo_rd_en         (rx_10g_fifo_rd_en),                                                                                                                                                     //  rx_10g_fifo_rd_en.rx_10g_fifo_rd_en
		.rx_10g_data_valid         (rx_10g_data_valid),                                                                                                                                                     //  rx_10g_data_valid.rx_10g_data_valid
		.rx_10g_fifo_full          (rx_10g_fifo_full),                                                                                                                                                      //   rx_10g_fifo_full.rx_10g_fifo_full
		.rx_10g_fifo_pfull         (rx_10g_fifo_pfull),                                                                                                                                                     //  rx_10g_fifo_pfull.rx_10g_fifo_pfull
		.rx_10g_fifo_empty         (rx_10g_fifo_empty),                                                                                                                                                     //  rx_10g_fifo_empty.rx_10g_fifo_empty
		.rx_10g_fifo_pempty        (rx_10g_fifo_pempty),                                                                                                                                                    // rx_10g_fifo_pempty.rx_10g_fifo_pempty
		.rx_10g_bitslip            (rx_10g_bitslip),                                                                                                                                                        //     rx_10g_bitslip.rx_10g_bitslip
		.tx_cal_busy               (tx_cal_busy),                                                                                                                                                           //        tx_cal_busy.tx_cal_busy
		.rx_cal_busy               (rx_cal_busy),                                                                                                                                                           //        rx_cal_busy.rx_cal_busy
		.reconfig_to_xcvr          (reconfig_to_xcvr),                                                                                                                                                      //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (reconfig_from_xcvr),                                                                                                                                                    // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_pma_clkout             (),                                                                                                                                                                      //        (terminated)
		.tx_pma_parallel_data      (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.ext_pll_clk               (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_pma_parallel_data      (),                                                                                                                                                                      //        (terminated)
		.rx_clklow                 (),                                                                                                                                                                      //        (terminated)
		.rx_fref                   (),                                                                                                                                                                      //        (terminated)
		.rx_signaldetect           (),                                                                                                                                                                      //        (terminated)
		.rx_pma_qpipulldn          (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_pma_qpipullup          (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_pma_qpipulldn          (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_pma_txdetectrx         (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_pma_rxfound            (),                                                                                                                                                                      //        (terminated)
		.tx_std_coreclkin          (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_std_coreclkin          (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_std_clkout             (),                                                                                                                                                                      //        (terminated)
		.rx_std_clkout             (),                                                                                                                                                                      //        (terminated)
		.rx_std_prbs_done          (),                                                                                                                                                                      //        (terminated)
		.rx_std_prbs_err           (),                                                                                                                                                                      //        (terminated)
		.tx_std_pcfifo_full        (),                                                                                                                                                                      //        (terminated)
		.tx_std_pcfifo_empty       (),                                                                                                                                                                      //        (terminated)
		.rx_std_pcfifo_full        (),                                                                                                                                                                      //        (terminated)
		.rx_std_pcfifo_empty       (),                                                                                                                                                                      //        (terminated)
		.rx_std_byteorder_ena      (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_std_byteorder_flag     (),                                                                                                                                                                      //        (terminated)
		.rx_std_rmfifo_full        (),                                                                                                                                                                      //        (terminated)
		.rx_std_rmfifo_empty       (),                                                                                                                                                                      //        (terminated)
		.rx_std_wa_patternalign    (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_std_wa_a1a2size        (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_std_bitslipboundarysel (10'b0000000000),                                                                                                                                                        //        (terminated)
		.rx_std_bitslipboundarysel (),                                                                                                                                                                      //        (terminated)
		.rx_std_bitslip            (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_std_runlength_err      (),                                                                                                                                                                      //        (terminated)
		.rx_std_bitrev_ena         (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_std_byterev_ena        (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_std_polinv             (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_std_polinv             (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_std_elecidle           (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_std_signaldetect       (),                                                                                                                                                                      //        (terminated)
		.rx_10g_clk33out           (),                                                                                                                                                                      //        (terminated)
		.rx_10g_prbs_err_clr       (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_10g_prbs_done          (),                                                                                                                                                                      //        (terminated)
		.rx_10g_prbs_err           (),                                                                                                                                                                      //        (terminated)
		.tx_10g_fifo_del           (),                                                                                                                                                                      //        (terminated)
		.tx_10g_fifo_insert        (),                                                                                                                                                                      //        (terminated)
		.rx_10g_fifo_del           (),                                                                                                                                                                      //        (terminated)
		.rx_10g_fifo_insert        (),                                                                                                                                                                      //        (terminated)
		.rx_10g_fifo_align_val     (),                                                                                                                                                                      //        (terminated)
		.rx_10g_fifo_align_clr     (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_10g_fifo_align_en      (2'b00),                                                                                                                                                                 //        (terminated)
		.tx_10g_frame              (),                                                                                                                                                                      //        (terminated)
		.tx_10g_frame_diag_status  (4'b0000),                                                                                                                                                               //        (terminated)
		.tx_10g_frame_burst_en     (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_10g_frame              (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_lock         (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_mfrm_err     (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_sync_err     (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_skip_ins     (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_pyld_ins     (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_skip_err     (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_diag_err     (),                                                                                                                                                                      //        (terminated)
		.rx_10g_frame_diag_status  (),                                                                                                                                                                      //        (terminated)
		.rx_10g_crc32_err          (),                                                                                                                                                                      //        (terminated)
		.rx_10g_descram_err        (),                                                                                                                                                                      //        (terminated)
		.rx_10g_blk_lock           (),                                                                                                                                                                      //        (terminated)
		.rx_10g_blk_sh_err         (),                                                                                                                                                                      //        (terminated)
		.tx_10g_bitslip            (14'b00000000000000),                                                                                                                                                    //        (terminated)
		.rx_10g_highber            (),                                                                                                                                                                      //        (terminated)
		.rx_10g_highber_clr_cnt    (2'b00),                                                                                                                                                                 //        (terminated)
		.rx_10g_clr_errblk_count   (2'b00)                                                                                                                                                                  //        (terminated)
	);

endmodule
