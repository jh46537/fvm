��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)������ɷ$neU�f�_�`@��8�����Y�c?����ؑ�#���W۪�v��5��3f���D~a����5-�i^� ��Ȃ�kt)xA9wѴ�4擃��k���n�.KG��9o\�D�UJ<���N��rgئ�,�)~���P40�xv�툒o��'K����9%|iU`��kA���M�!��:l��ak
���8��'  g�ߋ<�{��O�fHi��'Gh/�h>�1���g�.8�C�>r�]�R.�Rp�eP
1����e%�~/�,�7��_/0�I������n���YD��O|K���P��۟��
D	�u����R�;����1\cfR�b���%�#'��b����?��,#���؂ѿ@��L�,�_�YAe{?h������~y��sIo�$1��?(BY���X ��V��0�P�r='��w�5O��"���Wht��"[���v�unq�;���TLu�@��%���Z,�M�Ym��ђ��Y����l��8#-Tn=�3�a����C��ۑߜc/����+!R��j�`5��X$ĒƩ"�e�;��������ݖ郞ᨵfa7&O�^ݭ2y+$�3�c!佮zL�̼O�Ԉu�xU�Bۗ4	�@=�v��|.����.M& �Q�H�`�8ɪ܎쿿! N%I<�\�ɜ'�� ~���#~1�>�~|a;�q��f��*C�ӡ	��kv��]�)!���WT�����Xs���f	~M'��">n6��#�Ǒ�MZ
��b�́3 �8����l\:�u�:�5���[[���t�0��x�����7�O��B���ߊ��ǘ����P잖��NF>�Ab�0T�c5f�ޔa8]��5Y�C{��+�ܠ�$��g*B>Cӭ�56Do;ILڗ�	
$��5=L)��G���!�>�o*��隞+:�z���T��9�?T_ː0��J�ʵW�@�P���|���'�>�����kP{�Ѻ'���#D1��5ٕ���}�~n+��)ۂ�P���?yp�^�3P!{�9��U�]�Cc��5�3�4�-ʵ�����_y���'�7���W�+ ���so�m�1����/[��ul+gq=�5��C�cE�0)�-����l�MJ���ddP��%qc��߀�>LQc
{-w��oF }�ϵ���~*������FU���1�W{ ��/2�8��i�r�)31S�uvI�E~�m�,�Pj)�X��m4�r3ݸ��i����c� ��΢\���-�h�\qt�K,�.K��<T�R����N#W�!3�����7������y�������F�ߕ-��:�.��b�l9��/O3�\RF��5�1o�F�vO�9q�
*�Q"�^?e׵qp����eM�UI��C�Ct|��7<�< `�Z�X��*W�lJ�n�o�tԀ����S��%D�{�}W��? �8Xb�*3&^�}-sZ8�]ȍ5�K�����o����!���&j���r���_-��1�hg�m��Q�����YT�x�'%�Ӫ�^�!��3�������$�X(�W�-�V��ȴ�^�K�������6{Ş���w$":jc�p�jUI�����+9�����}x7�D{D�«*�[ha�	~�{g��0��@�`ǈ��h�_������Ց�5�:B8]��ڇƪ�w�|�LA��K'���ӱxY{%�/<��|�m�D��,�~���-�����CHv%,�m�)�����;�7'�}EC}�DP�$�%�y��g��5t؏��ӡR���{�G�-�@տ��I"��a�LrދD�~���V��ıb�R!��:N���Y��9r�c�������9��Qh_�2<���cFm�ӯ�l�1{���|���<�|���B����5~�C"Yx7Z
wf�U�A��p|!�Q�X-�^���p�{�IyԝA$C� y��7�-��4h���������Z{\6e>aR�?K�d������	a�%/Y��	xC�2�P�����9��w��h��j�����34~R�w�)���~!��u�h��1�z�͊<u�n��P^C�pq�RJEE��d@�	)J�nn���Qr5����J;��X����]��v��Ʈ"X�b�u(��S�T�T{ܱ��nRCm)[B��{�� �$��1�`G�C|=��5ޡQ��#j��y�;��Q��S�y�yת��.# ���4�^!
�ǃ�p�֨��.�KM�'�F�n;�����҅x5{	j�$Y~�1+Χ�O�q|�)�~!�p���h�9}2��:i�|ܔP���f��$|�"m8Yz {(M�Ǩ�#����+;�B^ش���qPj�<�	��oJsi%N�+Q������|�1�꯷�%o���:��u�.��iL���ImR)��J����DFwhM)eJoY̥ǄUΞM������-+��j̥���^�lW窸a��\p��͡��N��5�tk���L���5FZ�]+z9���*� ���$�d������u�D�Vݥ��{�_|���4Zle��u�9`J��� 	�;[��7�RW�̲C�\�5YH��gpkw�����$�t�N�;�A� ���f�ω$�c�d3�>
�R�[�A�M**�;y&�4w��y��Nw���\s
7�MG��4�0G�P�@c�k��מ���/�.�|KߘM�1�=���bc��1J��7%�罧����X泦�#�*@��A�A8.tq�q��{�Kg�v�]����J�?�m�p�N.oK�B*�\�=~����fě^/�Xn�~s��2p,�y��e�D{����B��������&F�8�jY<G!�±]X��B_R�އ�q��ϴ��I!��Bx�H-�C3��s���p(�J��{�R���`мy#Ѥ���X	��/�޼mxK�5��Ŗ49���e��1�5�=�ʽC�ϦT
��#�a�1��nH{&��X������u�ܴ1��\T��ɞP�3�Ä>�N{"ԛ�^Տ3��Z
�*?�({_5s��T�?I-� tnq9�j��=Y��0_�O2-ê(b�$֗�&<�wK?�?e��발�P�d�:4,��;vD,E�F��-LM�m*��/	�+�$!mqם���.?E�g};S�<X�?�,�����z��/�\�?���&$�#T�%2=��
"�	L-=��p��&����v���F�_Y���Ner����se~�� 7�ޓ�t��ކH�G܎=���#��[�Q̢��~+?�2��[p@n�uv��������X�[fy&��EՁv娕VZ2'n7,�,�(����U��[g����'3����[��8�̪��XV|w3��Mv+�������0NZG�,�Cz�Gf��!�gg�	KP_?�J#�R�a��(�G�YK 2q���������]c��*�;�6����A�Ǡl�Ĥp��`���5@�p�V最B�YP�J�?t�^1��%��
�n7t�r͢�oW@�Y����S��h�ښC�gn��C+��pJ� �z��y6e:��=��?Ä{���t[���SMey�_ʻ����k��-��:��v/�pTI
@vk�Bs�хH"{Orh)$�ʫ݃���$�ax���m�PZp:�:��Z{:h)F���
U���^��D�K�8��\�l?��Z<��VoD��MB�f�*��c��[%��=���{0=�P�]�����w`hhR!�/��/X���K��9I���N!���W���ߴ��\��r]�X3�$��-��'�DH��I�J�w2[�\7BW'��x�����q����*�
K ė��hrl,q�x�O�$7f!
�E�'��0͐Jk��W�OZ���ۅ�T��qţ���,�nu�;���&"L�P��D�q���j��R�<+�i�>����4.N���i�1����[�za��~���p�$n���2xs�:P|q��)�>���(���N��{d��z�C	��&%�Z帪�S������W�~�.H~���S������if�����t(�<NS���?�~����^���_~��ϳ�C�(5=�n�HZ��o���Hc�o��b*���,�=L� _�{�u�S��-[H�P^���"s�4��O�r&М�I��|��m-3�l5�����Zڤ;���ȹ:G٢+�������{��{0F½����I���(�� �}�	M�ͧ��