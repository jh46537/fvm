��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7�-�W����9���?tUo�2y�h�j�Nx�"��u��yQΎ��v3���Q٬���/o��5 �}Ღ�Q<&�'��':���uڀ�줏�|i�5m�]Z���h���z���lY����(Z���{/����k׌~5/��Ϋ�x��1���I�>u����ա��� ���#�V�&!U$�.�z����,�JAa�X�}�g�&�JrX-V�(��G�?�0�������B�fn�X�{`f>�/a����K���O���\�a�()>AK�x4�r^�<M� ny6J�H�jr|�ɡ��!�bX����	w[Źc_-�ˋ���,8�dJ���^@��i 81O;ee��պ��fe�'���aʪ#Ӛ� 6��+���D	GRu� ����1)ۍ?`�Ӿ��V�C�N՝U��6C�}����m�D҉e�o��[��w������l8���\Ԛ�c�	��'���}T�f��ߔ(��8eb�"9����B߂�Z5G�#�����ƍ���WչɛJ	��k[��`v�pA4[g���Z��ĭFW��E=�T&	����6�&�ô r�d�=���Vߌ�pH�Fc��B�,O]���~?�nf�Q(I�9YѲ~�>�y%��қ$��DQ�����p;����R�~�Dc����f�p`ջ�mr��[m���H�B�+�ߜW��.�ܤ�:��É�>>�>M}��;��@ʼvԹg̀�����Ly���1���4�?�e��T� �nЄ��A]ip3>���4���������q��Z��gqs{�&�/���E��b�D��-��Z.l��%`&��U��z�׮&}�����C�/����Q+B��T���i����Caz���j����uD�7�?f���[��9�=�˦��1�C^J/�sni���&2��^�n��������
}��ᩏ7���ޙ|�2>�9�	�#�pp�sd����`F�J@z9�k��l���8m�bo}�
�Ё6���J��Rv���A�J�"���o�t��#�-b+�O!��_EZ���Y�~�~|h�:�Q��V�3������-~����>���]��{'��w^|�nn�ĉ� #>� JIÍZ�
��$i(nN�a!<n����eݛ5Ȗ�~�K�Y�V����}Gh;�[?ʒ��p�+���9(�N�C���Qs�]���"4ftI'4�x6�n�}w}%DP�
vZ�:�el�4j\t�B���:�B�S�0Ȭ����lM�1����߭��pkb y���#SG/��}5t��yhT{���m?�)��1�j3�����r�5^��7Pea��j]ca���2��Jtڒid+dYN��g-q�(͑�rtu�/����ң9�#�'��U��9�Ë�a��ῥ�ڑ-�m�r�i�dsOɳn���L��7����<f�8^�XQ�ze�6�|�Ր�0	����*�����
L�Z���f�`{'5�	���X�	�9��aFЗ���7��M��'�0���U�}nO��wA	񗴰kBl@3܆�-c����VA��*�����Ϩ|�)�rQ�)���ИT�b�,p��Gɩ��e^F}��v��Z�Z<a��6���Qa���'EL�l��(W͓+V{^O	A͝I��ӫ��<z8��������@�)�Ւ���iM��y?.�h� �8Oߩ� kՠ���Ot����#�z�"0d*r��6eV��m2�?�B~�G?bv�{�[DMz�$�գ+f�.���J� A��B^i�3���ʑ��K�b��"�C��T��/�D�}a!F�8a|�h�v��D�.|F߯q�X�@���SW�o}���tUU�H��Fn�~ET&�A�Ã+Z>��9��-9��������>
�?�ɞ�,����-c�m�U�s���&�X��/uo%��;�)���L`L�P�n�����C��]��~�p>ljz�ғj������	mG��aZ	2]�Q����� ���@X4|b3j	3-|�4wXޗ���Ƈ�L3Y
�8�]'��	��B�i���#��*Fh��y.����%0}���]�ֲ��?8�Y�w�w��+(�X�`Y�)�@�ﭥI�	r�O����)쁗A[&�!������'�ěJ��r���EHY�ns��L8��1{��z\�Aq5~@��B�6��Rƽⳓ5-��(�L��J|cԇ|�
����Mh�."+����|� 63d幧�!���D������lOX�v��e�澹6��B�R"W�+�N7�/���	�_״\-io���	x����wI�	��	;?.�@�ة�؉!���[�6f�����/����v�6�5���j'U�|����y�Ty+�{���Ɠ�ۋ!�	�1��!OĢ(�A�7x��J���BTqdk�]y��o���)��~.��G�R'��R����x~� uW�����o{C˚4L5�W�EB��8�0������*LK����&ɔ�lI�ô�FH
��y�o�3�P4�z��Ɇ�_g&�%�D�*�PZ�ۧ��~l9��Q����eP
�A�l���3xp��}kG��Y����?�RmkCw��Vg��R4�u��=�	���hcò�����0ȤI&��m}�R��pכ������I��*�d�Dst��^�f�Ʃ��׍h�xd���Q�8�?Ä�P1Y �!�#57DԂ���њ!�`L5��9Ս�?����+��P��{�-�:�5��p���&b����J3Kr�qm$1קx.3�>A��ٳ^�a���@�fɋ6�䎳 3�q;G����Au3��$�ע�a}����1U���@�U�����Q�2C�?NC�Ma�W4w-џ�j����Cn�G���oV�j�;gV�'��˕�┅�ޛ���x�w�
��׆{7��Vv� ��|(\�2K�ة��R\~-��'�Ҝ��/�|�|��=K��L�SwX?v�J֯*b|E����F�*-O�����Ei�q����B��U�������P:�P�J�g��eAp�u��_�ɬ��>�t���y�6�r��ʋ�z#p���OK�̎�-6`��`7i�͊V5cej��r�}��D��0dH/2��i>���dd��l�i���¾4
����-�B?���^~*]�x��ܴ��>�ȍ����_��#XJؐXp��Wb.C~҉���by˯���Y8?�~j�ރ��+�"��.�՚��:�[��}O�..�����1>y��q>B�}p=41��s*�.��N���P��c�|苊QҀ����ʑ\����Fv=��5���f���I�>�[Y=2�G��=���Nj�4{c���|�~�IuJ2ߙ�Tq`��69��V��J��E�y��-��6Y�I}�zlŤ⥎�d�C��y^أ�AP��Y?n��T�sg��9Xli�`�k.xX�Z����Mh�o�YS%��6�_�a��Y�&<����d��|Y^�,=*�~AZ�J&"C��@���c�ݣeɷ����Z�vvA��ޤꩊ�ꛭ��)���Eȝk���w
�߶%�\�q�<R�U�n�H}46������T>< ��Sx�,����=1�����5�4�*�|��.��q;a>�H<�&��w��Ƃ��J���e"�TSBl{:gnF1aE/X���*�Q�Ʀ�\B)���e�j�v5�O�GB>ή+�n���k:�a3�<_��F&��)��(�9/����
�6t4X��l蕣\ʎ��D��G�D)�d�鮩@ ;X���;,T�5�4�s?�O}OEn,��6�W$2�'"�8� ��熡�b��[:G���������m�g����/3��~l���)s=�_��J��:�ь��&)|ȹ�h{�k�xDգ� �j�y���5��n8��c�M�Is�/m_~DXk���|�W1<��Uډ�Ȭa��2\��|P>�_���R�ؓ(QEw��D�>�K�̴��{�y"��yd�&�G����te��R��4����w���0.��"�l먒
�Z�ӱ�'k�zU=\w����WϳT�i�e�M�9&f�B�-�4d%��]G����)?��z�K�^�M��'k�H��2��GW�}ݍ��;�l���F��D���)\I��^���?���F�k��5��!���}6��QE�-�ֵ�n*)D�$��U~ܼ��..�>X�}H���/8h?��,��xf�,��=��>N���2��_^x� ��b����`I�p`�r��0y8J#�����ӧ�@��B�~U�#?��K&��y�ƪ���^zժ5��9�ٝ�ҡ��T#skU;���f�D���� Xs�t�-Ga@��������L�9��)�i�}N4�!���|)��翽��ç�_	�Y$%r={�V��'�2���W��x���E�I�[�����M`Dv\�J��� z��N����.y0�p��{Dm/�A�rfns�Bw�c<�%k���N0zuq���'���V�|�2ѹ�3���^��,�Ʃ*��U��|��b	�E���]5�z�J��#�j[�.
��;��Ǔ���((7pD�Z�������\�y�~nA�+�x=�nT��o�+�l�eW�蹿��J����׈s�v��)��;s�����HT�a�k@4��E���<I�f�4�[��G	��%�Mgǫ|]���x�\ �<�fW���3������''��u��>�,�:��t��
�% ���0�[����8��ЕO�iVϑ����pO.h��8�d�*��aKdI���g+�]�9ؒL�O8w��|7Pt=�m�*��_IR��	��X�Xl9��j �a�dŵ�t�:��񫑸P>\��M��Z�g1?7�uIj�)%�����^�o�=r����J����Hx��:V{=\�'$�$�2aڒr�hָ�f�Cu
F�V%�/0G[F�S&ng�FYnS�]��n4����}n�*�_�ڊ�RDjR��8CR�u�>�u1"���&,("H�I���˽�Q��r���>xQ�t*�Sݭ��o��!�˜\H�F��E|<��ߛ?�1#jd�����?+�6p��{�D<�v]S��QS\s.Q�P���q�+��`�>R!�G�/��6�y����x��	W�9�q��ʰ>e�ݹr�3V��M$V�W_�hhl�M^�S�+%ge'�}�e�v(PU���U��k��3���u�C�H���:s
G:Q��%-��+�����^CT%L�|�����%.��ls�O�y�jǖ��3Y{g	�!%/�%e%�s���0�n�4D��1�/U�n^��5�Ou�D�>�FEJ��̖����my&����R�H���B���@Feo:P�gG���Q�8^�"T��[�U��H_5��N��_,�<�mMT
����'~v~v�=w5��o�p$ C�]Ez:ؑ)�i���X�gĕ��|k:��O<��e,��2x�@`� k�D)��SiĆ� D���]�A��������˖_�q���a`����fEp�a��@m��m�R�/H�Y���h���1��1#�@�T��`���z�%�y�@/����bd�m�۝��ć�\:}bhDm�'��>�Ԭ鸡�&Rm�w�ܿQE�[e"�.��a��;p�=�T�
 �!'��e�n�
u�	qQUS%�	�Ot��F=b�>T����L�6� o�D'V�A��A���S�<e�B��7��&�_y���_x���ֶ!���o!�b!V��sޠ��^�B�[\*ԚZj����-�� y��A������j���ho��o��5C�}�D�{��!�â7{Q�*Ye�"�m�k�Mg��?�m����G6�	��aa��S��(Chi�Q�90��;����7AR� !�'�X( ��do9��w�,�`��VR�e&����~L�� /�#o.����{^
��	A�ݮ`ǹnO��ܿ�ۡK}&��
��v��'�o�<��٫5�_|{�p
��K�+!�v%k���S��N�`OFs��+t��Ȯ�=>O�M�]���0� j��"ط�L�y㎺�b�Z���� P"5�hݘ��aCS�¨��-��B_�_�����"�"����jls�#W�'4�?p���2�pl*k���{g���V8&X�	���]z6F�'S8?��H�bmÂ�η�l���y$Ͽ7Wa4�:;<��i=s������0PL�?����no�0\�3�x���q��Nm����-~@i�-6Ww�@ґ*�s)q�f��3����g�O�H(���x�Y�s�jɅ�Q����_� ����%E��T�!(�V�`g�����yN-1�n	�*֟/���C�^�����xt]��-˾3���s�S3����ܩ����dԮ��,�)�S>�{�_��IA����!#���:O"�QZ�ٵ��N�U�Xa�qn���Y�Vܯ����U)PVX�����pL�=_���?RW�̾�H
x���'W���?ʁ�PrH㳔���AylJF����w�o$oV�;��f�aJB��٦�����I�'=�:8MS�#��a�J@��=d
�m�+_�̙M� ���F;]TEn�t�N�q<�%�
�x�z͕%�A��v㉾�My>9҂y e3��dH�4��I͠E�|��L,:d\w�J�ÖP��h�,��r��ʪ�Sl7}�I�f�d)b,T�7���Y�;R�-��m{�����3�����M��%�E9Sywo�O?��^��� ��@^T�x5	�j�cM�+������f�|���R�Ӯ<:R(b�Sp�t(�K�'���M2J�A�B���2[۸�Z�IV����$�0��G����zPLX!�+�ĝ,�q5�@
|��(������?�vP�7�mO��V�آ��bBg��\	�5koA��^D-�{��!^����~G�-uv���A�y�:@>Y��A����:���S�����"c�}l=��͖_)k���AG�@�����l��]dүR�p~�)�f[	8���/��81C�������>��e���᳐1Qi��~
г���{HIL�a$�]�uR�p��C����܇�W�����������:�ɬō���8+(�X�}�W��ީ�tr|��~a��wB���]l�Cr��C���ʴU��"�)�B8K�K����9�e�>���RٜI{��+t��b_� z�ؖ�a�d=�%�͚�;�G���֫G��4�H���u .ua��޸([x�[*O�.+v/%�ґlA��i�2!o.�v��n.����[�[�ͼ�+��o������[[̙U�;�5��C����D��v�o�Y�{�T,��&5,�&&�&x��=E��!v9I�Ur�:s1+����0?v![��*Q7qQ�/?qŞ*^���ٚ���c-'C�@�az.Z�(o����-�(ϰ[�uNk�A®�A(M��r��$j�Z9����t�ˣ�rIY�\[��OH���熉c�Y���i��~�;_���E��K�1��P ZP$"�u��7����^_�Ӌ{�o]�Z��YFN�.�U0Ý]s���Im��j[���_t����*��&�y�'�+������i�	�]:�4�z�_��㏳a�p>�>�[���LvrL������N���ƈ/!r��3��HH�༞�D�� ����0��w��7s�$�yo���g��e$����4d6*�̿:�e���k%K�\1�D?��<&uޛ�q�-���ϫ�Y���Y��H�]�]r��� �
A�[T�-h�% �yҳl�������8_�ԕ��-��tNB)�K)f