// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lKDXjPAtnXhUouy1xRQSSs+bMaJhrLcfDICnOoireSLz3VBuh5HOeN2JiGFDlGPz
rG4N5G2LoX4DaYUIEdsUSI63/M+hQfWOoQci+eubhX/GMBC70x2WAInvkwHIwEAS
d+Y5HiBu+GzaM25kT0UlKm0WzZTLqN4XhfefYCh5+NM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8928)
ZhLV8/CCdlnYroSkWIeM+NLEv27eeqU3IpPfoGqtx4Ii+LmbvWovQbXhEpvvOimz
6wx87dix9kQ2kv25WGUZ85/s+Q+vkb0vwPreMVY7E+rMXpInq/LKAd5tm3Q0+hiD
Fi3yhE8I63myYApOp2dSnpX8ThbWDXA/QqGEUiMxIhXEySvZwJ1M3iY+5VVpG5lG
QybSCuX5szvFEn+ctnm0qqADDqADVmzGl9cP2GJIl3rIt5n71fxZmNLpcFMF4/yL
DZd0aMzZhaQU/G9EanJSXbh2cGsJYIf9MCMkSCiSWQxD8i/clpfkpQ8YE1+t24O9
txdY9hzlJo37IACfIR2V5s7bLRUwzfXvcuOM8pphOJICpJVUfj6f1snajBHX5CVr
NckYGXM/HqumufbjZsPZFKigJezDgZ4JR0VALnh/PI9j4ND1E2k8Ar164UnkGzLK
VcKBh46jdkgBd4FgRMf4x+erXHY6ppBBHs1jV2jtDkzeFAfkcqEH82jU//+H6uQd
acjp9M7aFM5enEE2SbB0LKJ7bxbHrbtp95sKbPbn13EfCqki3V1KaDAH7BvIZDPL
ZY0baez+5ioFLYhZl9yOuFdM9832VzQBvnxo83R0e3cdi46goZu3Sba/EAiTM+sz
lXBUumsk8wnEL6qmuwfwOykjYPhWYLx3+LQ8ABM3/ur71PX5Q5dWaFMWG5DrPwjS
cvQCJxwCcwEHzuTBtaA3BSGzTVxegTcntGROlJ6WaYyMZ7EfJo4chJybspVsPE1Q
vnM7i/1QrSTw2Ny+/XOZCzRZB71vm1bv/YUrX1+WJdMkJpQzdBPYmE5p5nZqzzdB
bjtIggBfohiEx1ZPjtL3KFRKQBe+1oIHOUFViwtV/Un0OQ3VsBGTps3CH4K5BQ0g
5EMMEVkARfVFvtn1zWx32VxOCMemS3tEvtkZud+ImdZXFADbZVK/NvnDEv+eOzCW
sU4flu8PXLsctDR3BY1ArafTDwAPyBojWeezhLOgEl44FyCPBWqpWuyTE6djNuxA
xuY/gfWZzG1YPUITmBRCkqtib/MrOqnka9xROtZAN5bXGwkYDCEPYYVYTuB5u2rF
q47pWgH5nI6gl2jtWl43IcSL0YQK1/1a79jnDvwjYbTTyT3bzle5U3a8Xwd81HOm
Dr786/urH0MDXtFejPBp/hFccXm4CVh9jAGuVwxuHVDRo6MARzHTohWHkX2N3Tvt
EPw+lAmO2LrF6Gte97UL7wyNndXi2Jww5x9bVkYfbWLxXYYjYKHTvqDuazZPN1IO
2Z1cQNgf97/AJc9EN+A458KNa5rCWK2qAwz9MSFYJUmjmXSdRSV4YgeC0xDSsl4T
jAVBDlpmPANLKMKhYb7WjxYQweQD4u7TibWHZTGfJ15RWLouIRYXMsR89plr6MeY
Zm/UGQkNPeFcDlHdGk35H7QjgcaOiH8T0B/ERlubFbdfyusSH+px3r3Do9wJKkzG
TY3guRMB+PSNUBn/eWfW22GrSreCXXd72AwQgb5odzn7zz0YvBqKafaRHkUIZDx7
qiRr88/jYSPfRm0xhFLI3jS38L7LSzxhfTBgfRGNMYNxmrj07e5MNDlFyieq9ks/
Pssn4yX0llbr4URhmMd81eGpFa0dBiOZUEn6BH5MalSUS/dWDRky8Yx5oyi8wB66
rR/TzB7XeF0N9ybnvsrYSVHnjV6+jsNcUB2l0dpAbTQTSYBG4NZ1VDCBD3cgpK/I
wzQ0PNiAa227MaPWgZjetIRQrizTLyW/Y2tDLicTaLXvNfhdltwyr9wJRtoSsLPw
Eq0D5KWzW+bkUhlPU7FSF1TB5eZEceboMh2yHmMrzWjs5+EVy25G3VfstCOe15C5
QTCATMQppw3zv3Ik8lDK45+5z8T1NzsUrEJ+Rb3gXbZCwp7KbMTjAf1L+fYXZ4Ou
eQXHZBuzvo8W+8u1lAxF1/NAsR7rQknYYMFIKiaf+21cRaHhBoTO5FAUPyqKKfD7
zbb7bFRjRV1Q8Z2MwbKOYzSplyWg79/Kuk4N3Yy/mQ/zvIHQDT6Awb5xrB7UXEV9
qeIxL9ADnnq1IfUe+eNAv6Keng6AbqebRIqE0Gs9BKA4HcfRH1ASAVyylihrvXl6
w/jcrXz6/BR4UTb2RZ218JhZXib7rSRbojkH9UL41sSQCqjXStVjSVCRMdO1lXFB
fVj5KLNd82tqqOqEgpZDg2wpjx3zHZ0nKeAwaiTXq37Nt/nvOJNeKl3Cwy/n8XOO
OLZ7tSKlvJN/6i15xaX87Z1ZhQQvtCSZAaoJNe7Kg3gRacYIjDxEP5CPlZL3rAv8
CJYldP0OjRpWKSiZOagWpjvuEUpYOrkjtWRg2QxmCasU+L/LYcL7G9aNOYAAQKXc
cQ2B682CuhvCPxEKQitB3rE+R10nbuoORxs4lpV3LzRxG8oGiBx5YT5panLCgzTM
9K43WMv+uQ3J2KCbKya0fXnxP/2lyfhGoL7z+QTuFbfI6XOurZDHwRFFSj0xmNgW
x+b6Srz0y+mPZsNlXJGXx5rTc2VnuUHHieXzuqRIIzGHUGd2kg8ya1rONQZnRpfq
cGZh7Z7Ak2H2Zgd9R3momrL7CQJDb4YItvUu/+/Qy3RRUVBnWTUNWnm6fTEricbc
+cMMncSCp8mH0pQ/F9tpBxuwJ8GhfAwKWbDXXi5v5CSRS/rVaqyeVRIoHb8i9bXT
jmlN07tCQV8B6sUl2x8ijOUDh3r1Osq7aybSL+1Q9YwCc8Z+8ZVOG1gSgGOt6DKb
Frb+Y6ES5hVdeBYaUQ/ftD+WqnPd9gRTa6c1xW+3vek+toChN2qThamRXRuD+hPe
fEHfZGO5fz2dRQSZrYSx6WGor0QHnicemwnNN7ycWQnh8lg1zf5CDa6dgt8QSFx4
tcriKWquVHDXzPr1Havdha12fJ12BseZjYCVZwCNx6zBaJbW9l6dchc2cT53WW5Q
+Xrn24BUZwjPQS+1QmzAr6eu+kJeIABUCKUMbnKgLe0A/RoExlpeJObAbPOfxKss
ohxr3MrYhTR+QQNaF4YOGrUwYSF3Mxyy2EpNQ8upl4KZyWWSfFIZm6B+XBIsf7cB
DYGh64Qcq9QDJcwk6gEpGoyFaPXdhSXV95x6P/P81Xrq3jnF9Hp/LeRMvexzJFJt
SL4G1W464BBdfK+0eBpiq4jpT6NpehO09hmV9CD0y3FteH3HSqNY2MGqX4H2zjFW
Ir1oSvDI2kbyWN1l9lTWQc3PcN6Xva50oz0Z1lwIOqhUiK90pq338FkwtZJZbD8b
Gsg2MqVzDT3Vs8uq0adq8lXrSIww5+hDyegt/IzRbV9jQI1HD8H7Via8iSZc6QvT
U1h2EbYA0MSdtVajFqhKLH/1U2IJk6djDsb5ERBeAEv76pyiXbPUyUeTlHrc6nKC
n14uQ7yb9pmvRUty60Sa4w958vYj+j9qgITSm+noNPLARyJrR+YgjvaKXQnmiWHK
nJe2tLLaUIfWX4GiyFHz67SeX8NdVaxSSepRFp85bOmnKP1JVJdO20fgXXvapzaS
R7YqoFkTLlTT8nTQvRaXwOuG3amu1w/8Q4ujP24zetfeNSUQDfFLulY3bt3plir8
U9486gFQAVoA8YciuTTkngjZeDqudFQ4tIDwNNNjjmSwed+Cixj5qVAc/dHlTkmp
UB/I23/NAkCeM6r3w63NIte5WwX3m+Al3Ri+MVzTit3hGZDGRGSDcvqfHZZPLaG6
mN6ZL4Vy/lMXQlP/DV8ei9KuCw1fIPhpwsy51zLkApyUfmQYqIwH0s2bO93ZBW73
O1YpEkxk4dtoooovWh5l66jp7m7T1v/eNMkK3UkEwIJ+JadaPCYTkHeFjkFsinYs
doBcRRZqN0MAY/OPE5L0+1Og+ffA/SwFTkHkH4gC5hiSG2c65c2E6FJoyQ4UBGQy
eD9715R1rsitH+pFmMS3TBa8NMy4+qk7dQ/DxDW45nS+msNGtBRsyN1A8Fnhy9u9
N7yciwJALHM0NP9ZVlJ6qZXh9JQt9LCri3euFUVXNXOyT/+vpgpQ2UPqGK45QZB9
PJQe5fwWpWlX8xS5i+kzkBKg/7emrt4OngK1Ul1LH5iQPr3+RUPbF1xtA9dU6mhf
mLfZWNUAzmtZESuIPiEIxlArLvn+tJgJde+MSQpaGwFl52HzQx9NBYo7f6wHyliO
eo8KOBZpMpc1uu+MQPTJRxyKLdfJ6HhUuR0G9cTXah/GtK37bbDBRhV3NjhxDauV
Ts8Eq+Wi9i7NqgowmwWmCfCc2f7bn/z/swWNVYPjOzoNXwtgt/iHcRLAQyGxJQ5p
w7WjwBWdo8eAzpdzwQa9cLzgAMtYCsDrCWJt4EN+zt7mu6JHpfxIoN9zp4a/mAU/
QAXuE0Qe6w/1rxSzQOEq/acemjCCtfdvDdYZ8NGIkxgwbH4D34S6lfftAHWDdRDD
gzsdizLSW/HwyJJUkYbim50+205SMtvD3RVisFYB4++kU+B4WCsoUT3dRzU47qGm
T8bRmMeQdHWzMTXRgS2FVw8a7BZedKxXPyycALBnj3IQns9bp2T9Fng64zjeb5tv
UM52y8QN8Euz6J+GJL5SjlVtvU0nA1vOy+2r5DnHEbOVRgQ72kOUwMVjlbsffNO+
bIWcYV/QgS5uC9kRaZD5gNFmWshgPPGq22rdyOH+bA+d7nai4LFWVKNXzCvf9smJ
apo6FgJoqzQf6c72vXyD/Wzlz73m1+bzyPbZISEEs9JXuKc+rLf69fdtdrVMHI/X
DMtIJFpiojni+f6PBmei49FDTN4iAVgliRgQwNMGbcZclX++WhfQe6DgPgXKwUxl
BIiu86eibjkIZguAq2DPeT9SMKoWRAqY+vp5kS9zvwVzn699zsGl+MGYKyTBIWqY
tXV/Tp6nJ+y8vz1FIwUDSVtMpevO9TUw2vRvjiAyn4urxn6kXg/Y7FY8ANKEvbbS
zWP/lBWGFwRa2TxgimNYVjkHoO2uJKcNcmXL4YFewpl81/vKOObXVcei3/PcqywW
aEFZmozEXGPRoh7CY381G1ZX9ykGVSEHjAwFMKOrz/IaJi4+JjXl55eyhMy7QB4D
81UMP85fQh47N3iho8Yx/fQtRzdubfUECQ51Gm1DeLMXGlxHwTU6QnnknVBWuq24
JN+7MRI1qYcFHd3kPH+RSI2k4fdt/2nwlgs7dL6K7WHhfIZPewbM1WcEUIM4rIIm
rsIoio+dldUc/gzFnDXm6byo9PHlcA4dR/Pg/tz89660CJ1HlQkKUHq4iq/NiXgb
t6Lv2vNFBdHZLX3YXFrMNSSQs1QqLSwwTpNh9bOryXPhOBdi9d4ip+NJIE4p5OD7
kxlDo9qcyu/EWEZSQTSzbI4x0lpDQpoBad8Mwtiq8mN/dcHnv/2LtwitUNy5ZD5F
zWP2IE07Yj03q4scZtSONaIQ4Nr+6hvWkDCoNcBZ0f55UhlF718ZSj2vnoVzpKLf
jFh8gLJG2VGDS4TgeqgnhLwSCiUj1pDV/4o399DD+z0yhkyK0YMSqyWghEYs0xzk
VTI31lfXDOmNrfQOzUvcUGEqV1BRACE5HMjlzGwDgFdAwkq1zb0Q44Q9prT2Pg8I
xsqtHa75R/6eMKvtfG1d/LaayhI8h3JWdDgO9tfZ00YzuRBpUXPnMY7/niVF7/n9
AeNBogJX5/VRsV3NYOA2bWD+bu7Pomz5V0iaUdri5oedP46sIltyCOngr1MV65Lt
NanxrytL/oMttcGXENap5azqYKzJdl3tMJtrh/dqvTEJLZbIofhsYITwqxtONkxm
RbgiL8+qPYRaHlKuxPmcvx8HES3e0hSZoxSqMDO68YMmdyIPekLaXt9ValeP/Zqo
nDaXamYRkMayljUHwBGBmDZ/8SF3DeFAO8TP2ibhGbMz1y6YXePf7J6E4ZsOjGKe
nngr4BkDavkBplEcaayD3iDN3Fo5Y15fruMt2t8yE1UdivzzGay+5NeCxee5mJRR
8i7yI7R60SDcAljA7We18tRshPevoe1QiKcUTrH3qd6f3SFcKMDcSws5/j3sVUDB
jP5hiszocI1zjp17PTzupMNZ5cUHuuDjwCGK1HtebyFLvveRBB4Hw5ENzo/xIco0
KO5qpalR75hx43sEyLGm0kPL1muei+fIKhOr39vwPoLk23uwi6xsfHN4zJTi83J6
HAqurax3XmlpiToNGEfKNsnJVH7VbizBMHofUh/OkdTpEQJ51bjLrN2V8sHKOMkP
e0E5y9SS5lc0R7uZnnl6VU9XWBV6cBdaxuPBKpQOX9uLqpDOoeOFJDisNnmJzK4e
ZF+ztGsh3BhoxXmoHhSa2S0zD10GV4ADLSp96IPBGgqZzCwSdm6jtejtJuduBFWh
6cxc4C2bA3ro3mfy+usVsr7OG6aa010RF5Io+2hY+PUgcVrTkI6dURX6U/2Es3Cf
d3r5edIboTDFEAKZB8pm41G3Zmhc2wFmltdXMyhy8FIMGdmr2rKYZsxZ60tHc8xo
scIbhA5WZkc5ma/fkpbYj3GXCONGxqzLHTH/crEpgDvopFwLxJyrpstt07IYFkGX
Rb6KMS7ZHF7dvNjt0eH4pHgFOxrkn5VdpPQjuy830EQ1L94Nm7GdYyuQPrIWpiqk
gakrh3Fm/mLxGDnmdKfbeeu4d8hJAU9fiml0mKCSgtGbzY32UtFQPc1c1tXvg8iD
RDguy8sAbklQ88Wl+CLRgaYobef+G4NJoUyeIQ88WTcK5ya8Kz+ak7NKL1xdLdww
4lqI0uswG5WGgMvHXFMsANPRzcq8Vb6AGi1jz6PHyhRap0h+avHp8wKSDkublFXY
BUbOlFbMh09U0YPMx1iVete1qETkr4aiIRoADzVpQMAvMe6V0glvD2KTgicHw59x
G6LAX81wVemG1pbA/+adS0hFUDOkfl/NEPQpP0uRPcyKMPLKDNb0LeVlJpCcw/Dp
33ESEzMMfWU4MO8zV2DFuZgcNWo8cVEsCbtvuK8/3e/It5h4E7MsPB3yf6bnhkQE
AGdyeXT6xUyrQtznwVu6re666GWiPLXL7/UwmpYK47mOYafNLZgFBqzdedyMk+yn
z68PniLeF1Z2bJwjuFKBiqeYPfUWpoa6fGLs+yZq4cZxwn3p1u1Y1ecW5DEgDISb
gmhLYqnkfZ87Cjj2IO6sGDExB4HqzMynW58xbf5wChdgtkDpVbGi4rblovmfJ70a
8oj5cAWFil9d0Kow6MqlXkYEZYNQlV3kJyw2o1F5NP3igZwRt2C4ciOir/YeY0o9
YNF/xZdTH3SPP2hVGOIBxPHNUAlkwqiTDLnSvZ9i6rKceDJ3YvXTOi+KnTdQP0fB
zGkfNHH4czp2NZrGuctZlzGgogBN2lnAaEIyxouDHXwfI3c7kItKJk9rSL7EYmcf
qkXxWwWEflfmnnv0DrNn1uu1jfW8+CjkzaIm7MkwVrLJTJ3FWKAvCtdytoO+M0Px
KkKCt9yBebBfg6Rha8R+dkKWknGlIc+hEK0k1o1QEDecbmllRoMo9lBpnTwdzHuU
jLXm4PzGNUOIHkg8PeJfDXj3FqMbXLOlpo3NEGzn1aB2q/PoND2E0YL/ofOWflLr
pm5p4MGMLKzCxrtZdM8yvyIecDWvMe5zoz3o/ewdhRwlywt/1QnIXT68Pr3hjVV4
j0ePyAdNNZQmaYT2E1HiHyikUTHzIgInjsOn18cfHsxI1YCjLDIbLxNa/wydtDu2
jjjB8ySbQFEffbO4zku08f3CCMVzznRxxmYxwVDu7R4o4NkcVtP8IqSAnAQpvagm
/C/dH7okcUmfLITz+fIr/e/59aJSjw6di4nb2JYQmddSDRVo1Z1u5y14Olr/Oq1Z
1pvYMYzWvab7homwXoL51AFwSoUAjBdEFPUvpguEPE3R4GNG2oRyahgkaLTUQD9i
0k1SIbxA4jCPZreMmKpLk18SVg1yC0clBobgEQX4ub7L0UiQ/pPAlMbS5FluCK5V
S3AOCSLiCesl/R9pF2Dk0mN+EOlA3wcFmyycLC1MQaBp4xz3W5Q/pvA4bJlrqROA
u0uDcDgF/EEiB01uyurFeLsXjLQepgEP/1QW8FbUejSrek305vcBIBioy4qSEYhC
cH6hGz4AABeNvSbQeMPCTKUc3vTqAmXpJziHBJRAcpO2pxqPjPMEmR1s+R8Anrua
s3LF5gxS96j37ZhhJxaOw7DR+wTrHdQzL09aqDFM6BkBkacZlluulPYk3TuWEcTr
4ReFssX/x6jFaLPgrDLl/fTANWBPhXrT+McvpdWlxIBcW5Weedo/w6nW9JHodEP/
V6nhi3PtxF9UmMFwX/p7ekmyqZa/4d1bHX0J+x3WerCLjwTaQUYGP37TMUCJ28uv
3eWkL3NlN5Q6dN3bbYP2XwKA9vYU7mCigRuxDvo8/EvMRYA7/EhZTWKD/u341cGP
pENXjL6oVSTtPSbWOIY/Z41K8XNPXPEPJZc7Hdr0xLESt4icue5brBxQrVcj4fqA
35X895fgLtyW1N5pCkD1YFzHGSjyF2cn3kLM2wtnli61FWGuKSnDZQtTm5+JMgwe
MDQia0VJh7FA+IVuwimwde0GObcT8kpcUBp0edhjczytuFT9h1kglQeJ2YaJJ7mJ
sgeFiTrOzkL2OIXhWZtMEdEdD9am1NYxpmZFN6Pywbzv444isOX0ykaPAmG+JBZm
dsgUbVTiD4bun0BwXWJghoKGD5I9vvEbPzJaGU41ClZoXsWvxaQ/NjfsOk2h2tgV
IzMFuCl3QwCHzFxhxdDRPVJGNrAT5qdB6eUJ4QS6g3ME4V9hSzQgfa6HA0TIq6Wf
+x1nPT1Nb0Zd+/kdYkjHCLVKu/q0nLkDIMe5ZwUH11SZ81BDkxcj9nePorwTcP2X
HAQp9q34ovmk3UvrkpP/kmimKxVrf6kSzcVf2qEO+lPqZqZkBxp8WrEkRHZhLRnL
HmfJPZbyv5UZApgOwnToe1eBi09edtzzDnkvX4z0GJiiYKfSY22w0gUZNj7E/Mq5
eKhhpA7mPfP/Vfw6HOVRmSlDRwXldKzvXDdewInT+uBmFhwXheLZry7pRAWYGMdp
jONqZnuH5SWbvRa6+W2AcI37jxA9rT2oRK9w1RebC9lD2rUrM6wkrvGg+u1+MEgy
QYZYoY20lhh6f8U4S657LX4qXDZizDvbzgZhl23wBA9/b23LfPYJuQXNYOasXGKN
PhUT8p6d35qRh5qD5MRY+Gjlwx1e5OUM8peDeLcckuiBnho4lQzFvoty4kqn9YaP
9S7aPQsUW4vw4uOZeaWJjmTbL0rqwtdhyUJT0AH0qdq048zNpMvPC4zbZIFVW1tE
yEVTJtFHv9JY4R+xZjf8MpTHTgsR7RHqvyzi1Q6/pzQuHH9mkL5TM/QcRQtU/Up9
jr6e8y1rTdv40CBwKz7XWIcsL2TtbV9OX8WuCcb+OKpDNjl0/5qg2wS/+lKLZqc1
XYMQaymsWkX/98RmRJgADfe2hbXJJnleU+p1bv2IWxty9o0v3JlB0ClXkcHLsXER
Veo/uGSKHg2lk7pzIOUjvzGv+3xrzSyvFqzl2G04NxyOKyUZ3X+66gs65B8SNaHx
H/NcV0oRem6X8mVEDK34TMH/wXX9qBjUsbxTpE/HqXmU8oXR7lLSiTAG+vc6KsyY
V44rFrraXLN0ZjTqNBizQcOipcechAzLEKYr2Gi13557AebIFL4iUEvQ+Y3mjgeu
ueHeojJjU3132I8OzMCCgSV3m5ey+KC8JubJ975yEkjoq9cgzCXtpEQjqW2yCkDk
v3/GEzPYCkBys0rvL4y3BlbDS3H4/ZrL94umaveHMpopiWdPUGP0AeBVtZ1elWph
2ZSIYYQX/3jaIjsO29ekK4KmmCjOVOemIdErZXCK2IJ5wEcPcTqx1c1P6mDc+SIr
QnZgBlL3JkN6q3B+eRf5BADhLiSpB7TpIFP05gSXP48NMLwLDtRNPr90/grXga2x
YqKAKsVycsNHA9UW1Gsx7GuCZkv8OSFbWghf50tMbEgWGu4OU+acRB8sAMCHYPJ1
ZVZ2csPI6gey0n5sgU1yILK80UX5jzX0Hn959wFMFnk0n4YikpbcuN3F9eNSHh98
DI2GKNwy3ad1oABpO2B3jpVMu7dMe2MSCJ3hamLhHSUN998NmT9vcl7a3wUfSWAI
tStYkpZgDMUggLinDU+59Y+VrqL6JEQUoGkehet1/J/K2g8Cu0wD+L6M1XnmNjJR
61vidGrsgonUZBTJxTKB7KETOBqdokh9+nUs14PItjvsNWb/qq0aTinI2FvNTPU8
VpqzbO1ZYXb3VTJL8e5Df/gjtaRJcF0kOp+K+SMsOOCXQj4w8Aatffz7xdn7VRCd
DltxNjKoTYmd7anUacdK4fbP5wBZI/AgvznDGYCwo0QElrOVNspFy+HKdphBo96/
rjHQl/Py6nlFCIrgRWu0ZBcQdaXPiedL578Y2yIHb4vbaAoX+S/8YgfDuJsAGDOe
4uCi7iqgB126mPh0QoepAW2h6RI/hFWHWGiVQf186VFnEFfdA89R0pMBc19qV6wW
+0Mk6fRIG1fxq/rEjA9r3krzY1xxcG84kXC+iJ1mFJlABWhUnmMqOrAGzxeSZnnr
ceeJ6MueaZ1gBpA02EYpukZjKgzu7CiuKI2kGDsXxNw9sFNP1pftfo1syr8VfFb+
mucx9ojd3XQwFNaYCkpxQCbfQx5PXLfFZmGSkAg825LEk2jlkCeywl+lMwlA+A8P
p5CLnraryAaYFSDvK4vnk5i9UtSBlUznRBZMzLbnvYjSmj/hF0EjPPgKE6cnZEvM
uRNYHqjVAWPbkkqWH2fYFeRHhKdZ9lS45WTaykoIYYUKOKrRPnr4Mw4xDxucwifo
kMnLQD06B366TXXlq8L3zXTxf6ND2LyGN31rT8F91e2ZiHCeffP7dmpQgdfMmxvT
2ghABK/qZQ/eX220rQ+OxGs2sKJJdM4sF1pP6Um0Xc+52aBEauLXpU4lctx+9QVT
KlDVxXnI0HGPO01OS0QFE4THb9CkVO1Was3OtxPKWilaL34Xbazzkzh1VBFqvEhd
ZPLbNIPToDP4A+qesFe/a3nBh6azFN06tEXjiaGLeHcoNL3p2l8J0w5R4hkvD/8t
gSnKBcYIuvrBwA0CPbxlpf3YuQx1Z0UcXYyNWagB9brPh/8PrC3tOyVOjTwSvKv6
Xvcl2bsaiXpcHo4j8iALp0zsHDBzOozVCuVx2Nrnc3sQMAfKByO5AwxFbt/Hu/Ea
Dw4ogAokowRBaCqXLiIwaeoXJyrh2MCfLR0xGVGrfihpcT8GV7ywXO9Dl4NuNUBP
jp62txnQXGo6Z5zfsI3EmM0kU47+sIV3o18V670w9I0hC7gxiEOH2yf/rhAgB0tr
WIdB8nylc95Pi2Qn4FgbAc4vVY0kxJwTBOmfA1ECAyeq2beRlVD7Y9C65Av6iesH
1DN/4XeVmtBB04yI4bagFOkVam29TA4daHCxYFZTb1IXQJKNDgX0VuS5E79CuF/N
7OGX03/nXD8N+sHQV9+YuMGMz+cmjDHMOqjLQvqtzTXTUfFXfpOXc4buLYryEFf1
gZ5Icy9JhTDTRoCwRkF3in7oLARv1yhSKgwRGGuF7Dz/DC7/mC8IzaHr/fHy2vUw
GVfa5CsvNorbfy69qTKKV6WzjF9lY3UjdpwyAkNu9nIgnSSgwjbKyj6qZv/Ip3PN
VZZYZFHlyLW2xjxN6+ZryM19P9Xpci6pXQmbRDoEsDl6HoOYn8BGefb9MHUhrp/R
xTYMljD217ynYVtLGN23g6SfBC3dMMBZsy/jUBdw+/lIoHuRKgFQIRPdVGlnvMYP
rfaqM0wxx+3nW0z9GXdNnstDNQA0mr/t0MFhwqWP4wjIY9MvcYihBItkM0O0T7qZ
Zg5UdweX3bHtoqMT1ETrM+ab1MJvF27AbFnnpurzUHzpcHFZroLEz+zrB3f8fV/9
`pragma protect end_protected
