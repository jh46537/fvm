// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PSQawq2/lUBhqKlBml/uyXXAbKrncm4HEw/upoNomb0pbl3DSkzkCs5+wDViVCM0
MJESx6y4y5WLquDzZ/fCdgTpyqIf4/3VmECOLBcIjMJxR9K4Qa5XLx3dKIqRNzCD
lCtaHsMFl+LNa3GOOiz3zZIlCmi1tNXv80Fk3xxzTtE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16304)
8P9az2SV2RPRCUOC+wy+u1jl64exjImvF35k3Kw6GhlZUpEpyT7i8XQQbWezUhvj
Zo8Nlxf0IS56HjYBtjjnd7QxsMp/ehtkBorwk7bHxrfv4w5MYswhhwBTKBPeErU3
A3AG6qggs7tggAGitkKY1qNdzdIC6mq02Z0GYvkH9pYRUV7CqDUgZwR9Lzwr+Joy
VT7+q3AsorKyEaPT4tDoWPkSyx1ygHKLG8I7nKZ+MyfKh0tGe6pqvACDZpuU1J3X
oOLQQJ3jNLp51KNmNjcWXozf678LPKWcaaVX9xUxKdaB1sl6hH2Zk1J625PFTrPv
3rZq5Zl9dfGnFVfrMEtCjX9eLJG+U9/3wLqdrquYIIBgpXoVlnpoC5/wMfjNqJzi
HVtDjKy7vfsDho7xtmNrMgtcYeUPuZsCbeN7IXWplkwsTBpnhep9FxBvVDsGgUre
bAPFozk2CtBhGLpwrWcdxz0/vL2oRr2PGjdSb3XumKEdhYPz3dW7gLj3rPVGGB9A
HiAAIQRIYNYWXNFrzTJAPZ87klYwvtH5G4ACiQD+a8gpAcnWCHZwd9IE9eIQIbMm
JIoTvwg1TWzGl8Mivu7xBMAeg3lR72Z2xPg/UOWRml5h2HyqhAHFz65qydkvUrAY
M1UN3KU2cUXZ6jhom2RWKa8T8oM4F5vRAYFU1gQmO9XyZ17FxU2LvWVrbYSz1eOb
QOHrHObb7lgUPbEzNRQP9ZrGwshJfL5aOWsI4zBWStl4O8GBxg9taWUi2RkueKbY
S1jdL0lDP7DqCKehqefyeMpUjAp3yOrm4GSLKzuqrOAplbXhMNDUzBJC3VmBunHf
vGDs53RzJwn+E5WUzLzXUEppgUIGWVCW20/iR8gotFFZ7wdcKW2emUkCODGXlv9W
9p/HXyunv7rq0qcQ4f5j8ykuZIu+pszxkRiI5oDcDyti46hbX+6kCEiXigmYuCGm
3Lh83IMER2Ec09MYMoiz4SsWZwX9gSzBc+mx3L7LsxRbLwGUAefboKvHx+bcGG5+
EiAblMtbNXSyBTw35jkm1bBYtztkPzWMKn1R0euNEwTJl+R391aJEu3uAY8QEl0P
ia+R9y1P4KBLsxog8IeNWSmhqqVpX8/aozOfHMQE7spOHEemMeIoLU0ztEY2NS6P
3uYzsSA67ZCbU/4/P6QYoLUFKk6dI9NIf6PbWrQ6IVNWuE5Lcu9kqvEqKg3KsLvY
+H9/a4kgMs5+CR8pSx/5IkmOvV6ehTNR4dxOolfJyFVbmMgpxDNEq8T7AumCnlFH
AEF7omB8ImMVESKdBZJBu7tVhDeAQZbpDZLZiOG/1NqD+GjtYcTCyYz/t2BfcNbs
Mf/Nm7UCGsbxaQdaZ99ba3glWeUsshK5OR0WuApWle73/OcM7FgboglcKlChZEjx
mc77mtgnbUKIb0YrKyDljyxPWUbaKhkwaqt8Xi+isiwZaHMk3g5PWmYhEtTd6qRd
BkxeJ7VAC36WzenNV3Cn4OM0869/s3RZUmAe0a8Q0s+ji+1bsrFvVps74acZsYc7
n93TOGwgD5W8oT4JwDh0LPFsmgiL6ehVcOrHPk+LjmKfJnB0QdFPs6mm0mpUbHFz
pyoMl55yf9z0JAaCj3KaPVskROCwPLGHd0DjbKaHRlnH+4z2Mdsv65e9GJBHcqvK
+iWiFLUIcWTmHwsLGsvPdMDY8vUQUUiuyWFGERwxBb3OeGkm8vZrOpoomvqnkDDL
pRsPmZ8L4JIKzOQuSTJOwwLWcc8jPA6Yu7TqK73iWL4FxGdV+H5XdyXcklp+/NFE
X1uZRwT/ehClpJ3v4l1W3j2KyaGNVNy1xkBSYfo5NUO4QCKRzVQvgcuqsqq9Y5W4
fZAR4nLcb52CoP+hD4Z7hHMJcoa3CJmb9b9Zybdxi5eUNRT6Fq5nIvAB0i0EBPWH
3RT/bloNcSFZtHp1l4zpGFKCKzUvdnFL+vLXOumVNQ96damwPq2Tvq6RNpnzUWxX
0Khl4BuR8uF0tJ8xl/wFfGArFA09MLq3/iJ4FK0VETU7Wu970JQrqMVvMKA6CLGT
cdnPeIMX3OEtCM+Ae/LKzTND7ad69tTrr79ifv7eY+l1+fik/x8yNcXib4DQR+C2
Wqs/rUONUYDKWTZ+CN2tTgAVqixdJLBdT7lENenVlW17fOZO88Sn7vn06UatmIx+
bj9DFXJJze+e7Hiht3lrmBIDTRVwmeBJ0Vpn6kz2UFJRDqRGiDAzi4epGaiLe9X+
RMbq6AZvOFgYOBZopkBmFnHx5SSBlFswDOfTOaKukjkdmsTlI2Tc/KQpnu/Wsa+g
8H4/2/p+lDmGXr29R8yNnRWkPFMlLb6PpmwF2wpIoZZCD2n/90crjFyiRzwSXxDu
5PRWtsxFG1WpP9PLFADzYhtO1WvGx6OtVkwe0B6SGckWc8xX6d3BshVpZdon7z4Z
hnkEC7mCdK7hc7Bt6HCvx1v9mlVVga/ZH/h3x9DVcOhjyz7ew3iR452yzpUXa8lu
zzyn86Ter5KhXWaeU2UKdX6dSLGOzub1FoRsISgg1iLtOBFKF1Xf9PxU9j6nS0+Z
zCMDtW5aPIxiL051YX+7oJIn9WFwwMyuHPSGg9rS0lOYGVfy5rAglLv05pQY9tCs
tpbST35k9F3toCwmH8ZV2me9fkg6mCpIc0iahgXMtkrakWwduyrFGeAH7HtPT9OM
aPFVSon8Bjt0O1orZgLfmkcqqE2VAUqZee96jUrJO7n6OoYpKNSlO7XLlHy2RqEe
0yt7capgi4x0Jn7x7j3AXviZxpzvsUEAN+ZHVdi2/KsPeWr//3pXHCC0aCNY+3cw
927TMXO+78GyU6vI2vXufSovIAfI1j4yxqcMfxsmBS74aKwBpv91H++hKnIIg64O
QAi55qj+7jCsazz8/d60c9xUN9Py/P3BDnJKSQln0Xuq/iHLeujl7d4ysJcpIUi6
OPNH4X7ngb9D9sDk2hQ3gslRphKVE1mYwiM1v87cUGNmer5M+8P0ND9HO2089hJe
b5/dgYNRc8PX3D4xnOkN6w2U/hD3p8ZrJx6LcGHU/RyquIaCeL77UzIR1iIWoHEQ
ann9oKPmFViW+87iBpdUrCC3bw2WtQog89Lo739ZtbRRRsCoLndU/EUIfR1xW+zc
Vb3u1Ueu/vz5TOy5J6CTUzAgPoY0xr7ORsbIWEpcWFjyGY4RIhgjv789cOEStzjI
drHD5nbQ4NWG7KYDE7x5aL1rT3yHqvXKPwrCnWDLbBzn8vQ6VNTRLRI6FEBCwr4E
qUfZrzaX7NHxyMIE2hCg64EXcfrGkVbE8+0tkx19AVHXls8kOVgGaK3/BCD+vo/q
g+s8XHbiZ63X2nIR/IwAV8imZkND2OFDbKy4YK0sm9v7HwUCeOT6mmUW3YyHYG39
DvMgOVHbaQYSSp2pLa20W/OMFUDJ4Zau2BtEdPRhM3d5ZLx3FZeDN28R+/HewVfM
alm3aucNCYndwT7zWAb6pUHd93LJTYY0tsRD/5s0EPQCMpKmch6OCmvAMw0nana7
+gGde2lNrp9cr+deX+kO4dgmET9oQWPUgBMjBmNs19f0zTfel3TlEHPU48mgXWAQ
/tSQrzrbTkcs0+3d/1DQrR6NIo+9lrYGZx0yv6k7w5I9sNog+4XJnTW6z1ua3zX+
vE1VsnIhqwMb9pA8BjcI+EACejOVX/1RrxAAXiHab1k/tLjl5w1HMlVIlLbyvjgr
fwKFnIlYs3Ef4dE84RTkTrInGXJjAgd/tmvrbjjT8k90vJ1CstBrSj/B2lp5k3eQ
iUEG70GZC+s7syZHOx4dlMicDN2nixRExQYOeRCahLJN4f0Pu1HuMZ7mmlJBIroQ
sqQy0lZzWCNxG68FMC2TIssptZd72/hsKIrtlXoUIxT+qeMUMwT+3xHRyoPcPCgi
t24fJF7GYA1gyC79qCyCnjg1sU2ClHi7cw0LvvP26tgnwxCKH8mVMzoxVfTA446O
jFZQVWAzAhjlMRRlMBphc6DJQrOH72fmMbg0EICUx036YpiBQ9AxgM3McykuBRRY
pJ9HhoufnfrOviQhf3o1XbRyTqqfzU5T/B4WwN89wbjEwB3V84s3LIROqj8ObFwE
4yWk5ard7ncFnac7Tsa813r8UiJoVt7vbtQWQGocR+oYcU0tbY9X5KjE0Xf3H/Bm
r/Ho5QR54ydE6IQKhqwkXIVW19dhaNZeSS0fmHEq/AsYndmf26B73bO0pleTEnTj
MJg3bpNiMNX1e6rF019ewoMUN/x0gTcwgQ9Iezo7gjetNWzjEWMRlgQU4OgFMWUq
FM5tDGVtdm2e0qDj/YesarRzQhZWHNrNuf1IM9qsxlKspngpemwJ9CbeoS1y3i0m
kfvTTfZlcqgJ8uBJRqsVj+ZSj5qV7+p1pWwL8780A5HC/ysdSLOPbsRQfH4iNdK4
gAJHeZdxoQNmr2XtRiG5XhWhzw5XtPVmnezHGd47322/+hGhbs5clCS0Vd0YdIkC
pa58eOL9w349CR8jdPmjsoGcXbKHWN6FCY8oXxEwh0o3eoE6xhuCr96Kcm3ULBfG
iVupzUShhNJ3Z0mtlrm5dkaHtndOlZE435whiV841hkbNN+G9o6twtQEsoCRpaZI
maoT5SB1Kmxa48pYivbBROdELpdmks/hDKAo+iQGwHprxtc+q7EZT8xiEAkqWuO+
NHGc3w+UcldSbUISUpMLYaczamQIZ1TfmjpcEX3NmtgF7yce6+fxfYPUUUnzVmAA
Yx8LD3F8t+9kZ2OQojfvkwmjLxJgSy2jCraYoPGTPJGtV2BRqKOREPNGotm9USwc
kP5wmK7kkpUcm99emQBcaGdVHVRrX2yxYqggUirBNeDK53rKpBkNrZgZ2L8t9Eor
/uppD5fJRuB+O69c0IqMAuUeasn78grphCsdzVTbuBNszWL24KARtTbQWYRy0G9T
q/qzv5dm+KnLiavvoc2rbf81h13aQxDKb+H5LHjGUKFlT8k5yQg1VRjtMWHaJK7+
MHegcUoIWRPWsUNwlVG7Hx72QZJapoZsWU+VRRlIJkoXxqHPk/nUGn9/n6vx9H+N
JAnKBzxZDYgVUF1Mx8JJ7pPRdduKfqhRqqjvhTXpmH6zQbCBan4d2Iv2CKJz8uet
WoTT7WZ2epdLBcvxofJDZgjtT5nswsPBi+InIkEtEDYl4WYI4m7YAWdPLSGGKJLH
wWEloKr2nLj6Uv1b4PXWM39OCatiQKHbezhok0BeyABAc8OI3SriIgMpBZgP/FM5
biXQxWAaIgpzx9TaE3espJ3aJR3yGlKC+SYsau4m5k6yzYlcqp8mfcas+0QUo7ef
zimyxS1V6bDi8FV4F3V8aMm21SE9aeflsCFpB9xKTa6OlXS4K6afW85e2kO5XUbe
8G5OFNlJdjfbr2sOEcKSdW+L/H+HfT93dK+u/ASTN93kRI2P1D5QdssFke9epHfw
pxptd34oRabGCY1ucNBtyRYgfkjq9OwYM3CyoXIZj4+/Zl2NTia7/m7yc+HvNmZ5
ht3nEkvc9LibTluYl96NBd+QJV0ARk33qHnRu+nPPaxKTM/iaIBYPeJxHpndNdeu
h/l2d6EoP2ESVDrVDkW8Mv8jJQI6mduodLJkxT3FEpXt28rJWxjJNeWzk1ql6Yak
dLo5c1AV9/nHaP5dF8pca1ZiVtPzBJGxYGm//DgbaHjaE5gJdFJ+tcKiXiM8ey69
p66ngIefmPGiBAg046Sg4CMDGrtPBn2X9A15IDyKPAl6ZAfaTi6ItZF115GotevV
/k/Y62SOhlvOyCPu20TqdPsjIQfsVHZ6YnLMEq0UddI0NYDJS4e0usO1JB103i7X
JlDNQRZ88DZ+gkhNBUAWrRnZBnVA7pocc+mDoRe34dAOYfkHr/F3CTMvmqgvoj9d
3aJOBfirYOeH4lvUbyfFad0pGkBaUHmXbtD0DjmBot4xCQ8zH27w+ia8ghptSVQo
VOrwBsaiujT+bfM0TUZY4KLVHqPsJ4PQ61mEYHhbfzQhE+AWuP3Nnc+md9VsR/S5
NzNGbfpW+h44cmvdRQYwBdmtVuTYQyYND09gWMjGpOle0glCLRsD5yBlMYDRUXx5
DZdMCBPSTXvtg0p7BlOwjJbo4quk5WLaQUVlXK3UY2rOcn/zLDW2mOgnKj6GQbZY
Og7xW0VaW3pw7EXx/U0hleZ/6Kewac+cQR/C8rMKTXYnQbP8IhcgwZcO+KiegthW
kaVHY0P+Ym83ebYXesPZPk8r+rmLZ2SOimUQL1Rw8AlP6fgPEby7ZqVALJqg75aL
s62JWtRHH1hmNAdbQBZE3kNJF4yc2jrI/rtXsF8ZDoTxx3lgxY89587gx9Vs9xWN
dlSGh1U6HRFZimTl1yrJUP8xD+oQIZzyEH0irqkcoQK7MzSceh6SCox/FCVnDdJE
sHbILoGKBBgMAT3xQFYKNJirujbL8XUvVtBAvpJbOQ107JyoAHHr9d7eilGCs8us
WdVSKzOdiOi5fLyjgxIeMtsgEEM5ALzsxnLcYXrrV/kqRyPAjNA/7MMxKAp+S3CN
4h1WiWSVnPsXQoaX1ZvXII7acn5YuhYKhG7pQec987rqNLmeyj4dj3zJlhD5g4CS
ReoywbmKTh+JrbjWUP086if9d66LGxoMI2BieSEWuqy0wY0dlhVjobfvAgjwr2XE
OHyaamHtHbTvCFK8eJUnsvzs6VYWPPe1Kiz2g/kgjau+IukRmJc25jKAP4Yy7bPm
8LqA1CLaFcoG1hIrTdxfJyFsB8yAmneRau5tsdGtaXXdpEyZ0tI9KHrIoOQ88DK7
eQ6RPFoworWXVABMqpX080pVY8Svmm7HENJ33G9CpUaQnl5UIZbJel0pzEHxdw1T
Aw2avEFrEqxZVx+1LanFCbKaP5HGtLa0dvW7eI2V8El5s6zQuMveKTqyhQz52LeT
YVT4NWttFIMXGYDZo1TbUhVJqlm6V9RMGXj4RbPjGrz4CIvJGMrR1tseqsIEmxAz
f6YNW3jRZ+8aIn6ZuNPOZSQ7pF4aWBDwsKR+wnx5IXwDje8X8bHnEdBbNvD7yMvi
dik8e1/sDaIZAsaujAOtf3k0PkEtvk6mpVfBVtu+qEqjO5WDEnnhwyoBBLpMC096
n8QX6qz29QodcNUnC6XxittG0ScMw674xTagrGmoMJHsG3wLBta++8gWGmH9BShU
Tt7Qzio5z1PcAnldCp5BYFbWqWYkY/vHoV0AQWL3RXy6szF16149ElkZCD+qkUqW
SIAvX/OOABgpPMs2sUPMP1lfZLMCWgsJM/IDuv8JcYQGfLpExfyhlKI5yUOtkOAc
tOGEjKXh8nGIU8SbG/a/tCRVYC+KxHmLRLkZP0D0olph57R3nWSP9jKU0cpaR9TW
vgEhgjnokXlZE6+7z2QxcMtfVgptJ9tVvBooRMF9SnSyzNPlENe7SMV8MUJxpAQv
mr+9jG0/NGUOC7V8w1hFg8GzCis3ZSDrKZmovwuB1H3OyOk7apfyb4ifTJK+/Lrz
PeaSKlAX6Xd3RKqMhNgWGG+5AQiHko9Oo+RQ6f8gL5oOO0XODinHP1yjW1aSqSDk
m1lWi0hQj7Le9BluTU7rzV6T4ZHDC6pAo6GMiSZt3QOieHE20ElypZz9sLXn8iJi
85AkmIfySgLtDyh+qDrdpwFluDsnHkC56Gn61Lu7pYNR1DkKC6FKgyj6Dn0h8IvH
F5TJnkMXzUJI0lNbp8s9LROKjHUu2j8jIgJpD+KvIZrO0GOrX9BwiSaY+T8P3mFi
UTXUJ9vjgB2Z+Gof2ycbypspUa+hYvhINNHMKGpBawF6KIzJygatMk23/1csALcv
BHIg7ZoI23gOZ+EghK4H7KxFOWBBNkLlp7TQeQb3bm+VHjhUnq1U5sFN+7rZoSku
5Wg2SJ67S3swvMF8ZWOQsVG10/jhOVqO3uc3GEXM/L+K4+W32bvUReU6ENpm4Lht
KDZxntwNJcwHJ+Sm6dvkkg2yr5GKWgah80O/2NeMGLTLL1I4vnaCsnZsCkXP33M/
dQP4ZsWRacXrfTq5Dqxqyyx/1RbkhHgI8yb2vU4RXKw0WZtrR4L/TTm6XaZwiP8h
HC5y4AqofgKK4I4y77/fsquGzh5z6stu804JAubbriSYBi2SYFleT/83i3KsKI3s
dgje7HoY7N3UpTls9EPGZAO6HNWbHOW6pbsdC/fg41rwfxtIra3MDxZv2+AAbRrW
CXq2QTCHSbLN4RcAGcr7cZNREWhSKmkWmmeuNOyE7AlqjyKd9lSsKkAu5SoQXaqB
GhWeZeNUQjoXxYa5SrMSDmyMWOJGBH0jObIJRqP30M0kpMd16aGDc9FyV9ZEAefF
FwxHKI+wutalLjxiuT1irkP+sAlf9AhXSzHHZ3R8yCFlWDN166lOTTavyACt3SRE
GWAx7tc/r6vNNkwpLAe0oDPy8WlotoGSqEGyYxjjQprqOIbX1RG4XkF3KrT2oK3s
9/tN7VLQD+Jn5UJ/0dgFY0IGLw7T8UwVXA0cxh1AZgOd53TRA2LI5E/r1iXDQb3y
snVDtUJWnGcW7LebsKQRyO2/BEQqJneGyyJL9JTjdeNZGh/SHHcHxXiuL3+ZBvAX
VdM1Kl7kWwov1lZvVJrH8RMEOZWPUEDGQXHarndv1VmE7XSaC1WclzpcK2JbDeZQ
pQTE7ii010i+IRs3OPzsYx1TZ5/oRZ2hHyyjRIP3Ke8gmXV6G82ZOvHLabmEa50+
IpYfoy7F1/auoOiJSn/oj5xpbspW879yQmHFEmGSXeXzHN9vP13W9m40n+7fUkEw
tsh40M1qtu57nq0piOPyHx3Sn+3WtBM2SdUbTh/JnDPkvgqUtbl551O1yJPx5NbG
W9gNjnzHh76oBy/zMHx8/VS07c2I2KRrM7jLG/8BkYPnKMkddizPv6Zm1Uh6pAeJ
e6BZUx/P7GDojSwaZPpwSc+IfkkiHwQ4b3eU3ZNHNPdImMmmZHUdHZqsZIy5irHa
hruz1lR0uiu0EZ6OI9UysAfYrYEC16MZKccCxg6Xin0irx8S1vUM0FmclgdQMI6Q
rI/DDDmDu5BqbzaoSU4IuVP10fU94yjD34MpsCWkjpCu8ct13s8t5hinLGcz1kSj
gfOg0f7szFhqNBv3Jjrpdi/+Ghhk237Z668hwI6QLHBZjwQLKe6PCjQKNN2gSXsI
5DGLZtHGYUAzbfg7mZZ/6kVtvecD3fBsNaq5GHS2LPaWhStcrxT9JWCKLokBW2nH
45/ZC3eh8H3nsfTAupAcZYJYI7B9UzBPEw5oWc+oK20FbqFjJHQy22q/W0ZKfBzy
CEsVED4EB76vnAa8RirSugNA4S2ZOJClYK4+yTcafuPokoGPnQoDENddMTfyhOwT
TYFJqidcVxQxbzyW6OVmhlUMhOfpC+JGAwLymau8oP//QGJciOa9gcYepU4Z33Zn
GI1x6luC4/JyymIcOydhoG0OgsHuILhNhDteIgPEvQCO7ntpu7oCY9GftNGJ2IIt
94AE1ngzHuztbLBbYG3m4ypom3h8gkvBuMYYBQVK4soHTPnL+9yO1vHKrYqCt9pD
I4P0XB2+nzwY5sYGuJ3zEKHOy0sAgVsYVjnRlhRDF6gvSf2OlFZ8+WgkoIJABuPg
BsYAN3r6FtLmTnqt0DuS7nn3K44r8M9TrKgaJmqNRfxNT7NK7DW8OCnEikMUf8kO
gih3yCWq8V9t932tmJdCG3+lC9+gv5dJfodVvCZlMe6tHGKHH//uTE34A7f6wFRz
PF2lA367NoZsA1gnM6muHXIZRFP3XBayDmKjatgwQzc69IcMnupres/58h0mDH91
V4BQiu+1lFg8LcT6kKhdLxOC7rn1zIoY+lL3XuqWNM2kM76iZUWGE2nh3Pzylqua
T7U7zalHDj4DH/YfF3MGLZ7rPHB9DekZ+Iyp0i9TILIqMuUYqNMrXCZYC56Vc9ER
wn3UGGDp+xoc+LfUaGAOLcCOUiJU6QyBtY+b89izcNWZTQuIivaZK7QbFi3vCm44
2yH4CTm8Be3Hh1y8EhX36UWnEc3dR/qPTUltA5wJ/X71Bgk5iVMkAaqiclcgfVSE
Y0gYWaOlg2HsHIkqG5CmciW51bcGFWbzdn2CPFERJd1tIGY2XtQb2c0DjrrCF8QI
xNOFY1UGHvx27xYa/wjy+jldevvxdJalhJdHbNyqe+YSN3u3W1KPLFzEhBQbmuzb
zb1/s6XbKF1jSUnqcTs9c9TWqiQ95w/YFjM6CuwyUqKbyRkTkEcl+MZCoAJgxRlp
oAM43MoGroMvvEEJGAadqT0NR66SkTdiuR4gR1E03QX5qwvauk007J1xCruBO+mP
V07Mwg/Iyk4weZjptcjqmvbvZuItudp22dN4h6S2NRgwkc/zz5wn+ooLIqDQ5mGM
1fY+JEX/5Peo40N83ab7DtObP6uK4NZlyY5xTvD2JXdYSZEKGxLgKxGLHEFGHoZ2
4HukF0jawp1AFkbZ70pIQPNMmIBUiR7KAdbcNfKZ5tZFnUMCrsXtabwgBoI2zmAO
RB6HL+btfHBujo09UmSGWwoBqTrpHLHpcfowN3R+VojwJZgNHJDP8dQY20yW4Hpf
C3iODK5z5/YEvz8Njw14RSZ04htBJXzMdYxb4YJRKrxEq2MC2woipTUAbCKmFY6z
+9Q72s9DgBMMmWPNXrhuTLb5eW/as9thcyS2ZTVnc/Poq2R4GU9LuSWo8NmdRXa9
rEWd7mDHqYG+xPU9D1wOg2XerjAIUb/qx8XiuEOa5GJiqhLg71FA627deh571Ejk
RSS1dIdjboh8qThCvrTEem0ekPM8Zs9vrkHKJSkjdBriMBi24v+5kaLEUhg0+cT1
3G3Tb9V7CqC/vKvMBIyMVFOrYkE5Qp5qQehK2sHObS4hI3C9MfSFHCDwXVknYev6
C/1v06iMFwwmMmvbbdriMpQCLViciAZZk29k89IPb/Mp+GAdmdoBul/aaqf2MVuV
Fb4PotPVsq1Htup+vSNSp7AX+OWl4AJ2Fo4JzEVTptHuYgxW94BmeK3pQ+JthQZm
dzaTl1bB3/udaSCVtNay/lqEdazwNK8i6ef/gsOuThsXdQ2wm1BFF3UZTra+mmCr
6f3J754cL54viqwFQKeOC/IenGKqV/HRcg4nISAaErGsQdQ7aBMWWP67vo0lb8ir
vsFlU9aBOaHSbNxIBduWRqmv6ckd0uVVou1Od+kAnWiaYCi/78xsLFfptUvJ7W2r
l5UGKFKplK14AwpcGtzifcjFf1EbGDQvqG5W3zYDsPFeYLptjwRi+UFnHToOo9H5
Ld2j2maeT8iNpqe0VBw+NpifVLGNSxD4PxaJBNr00IUWCqOraLPqe4zcXVYB4AEj
FA1oiFwZQ/VgzQn4sxWD2RQaOPMx1DjRse9FdjYwfk1ZCmMIf7Xey3G03Ln5038S
Bww66l2gss4F2wm4ISFlI/zmMTYfK5cSsVLDZhOJxSYXpZHHqIlYYt09FWXcPycy
RTd3wB+3zE4EffrM/edmrYzF9bdipW45f1NCd4zrWo82vSgEdx0zeJPchr2nGjV7
JKdN6APIBk1k0h3AtDWNupXao7NeVL/r50H/WE3KLkdqao4ycpCooebpP6UZ51Tj
O1BGs2T3H+18gGgTefUUN0SwqIWj/y6FQ5f+B+L4npGsPxummWJ6Thjmt/nhZoaM
zeJi8WmziUqlSBhnhIgPL/LCt1Jvf/9UxAjJHRoryBgXBgkma0nmNpxZTUlHliYo
hLbzoGj4aVWD8VAB6AI9UGmfS9YI+elxvAc7/+fis605IPiVSey9m6+BqIFqB2u0
lcMbc0Eja/AOgmIJWn/hBPtJ25cEjCp2ZnsEBOA9f+/xiTJtI3bkU9aHS1O7KQhD
SvIhyB5w9d2tVzTSVjt4ZNt5LDNR1cuiipu9+X/Cuh2+YTezGSyyimi6pHpv2jP+
/5ju4FHdQBSIoZbELsEdDxfizOWsrN0breM8mAK2080hHUu9ePVrjpkbfmleYuj+
sJoTz/ElDA4S/QTIGJnW0BAQM8mPxuATdQse8nkAq777U6WEk9h11TKUrkjSCHhf
iyVHYOaFGmUdQNg20mGdY77AT/atPxz4PZT4/S8EVGezhzhy2f6KPXKq3KrN+c9N
AFuPAbT+LKsiMZU4jFmVQEBANTXQ7dFjP7bnTvMj1DcmchOPmLFFKew4MlsweAya
ANVzjKKb2IoVLmudPG7lX28LuKIcY3nRfpei0VhdnI0ZtB3KQsUrXXH97iIUcr6J
NPUQF1KH61rQ9K6lwHC2D1LTVJjd4/X04JNzXLOoStfvDNpc0kOULUokSH3sdSv2
htxFVZX5ZAZAQiFJxgreq1LqkZj+uQrLKEn0wysWg7/CrDoydvw4o2M/Vg8lboGz
JjPgwFj88YzHpQziEttnGkUN5dB5NuopjCA5/CKhNxJmFCBDMUucZwFx5xUffZLU
EpzZVuZfR+XxIuQhv6cA/z9FgST/v7t0zG9AwgzrZ5RWkVMMvbdsdDfZ0UCJWucU
7iqwwFXiTLJZkdqeizLMaE3bQwp/m4zM2v2kLHaiuwqMiJumlN8d8xGylrOniZ/7
4hzmFkLwjVDoMZPg97PSq7lWS808pdZuqJlBlYibMm0QuTLcUuYtkGSUdermBgat
vna1cTzbCJRxXEqfBxxDlJ4O0CrXWumlFdqFn7zMPC3wX7qJelomeLgcBPcCP41d
7M6RDbYHHkmP5u3A9Jx2/n2a56FM+vsU84j0qtDqQGb5Bs2CL3aYwV3M4Mf3I6k7
txS0w48mHu/M7pN2RvNhVKuxSzFDXgFzhNUCbjJAhiswDscsh+cen8psz7GJFGrb
0s4DajEtWmtM6jOP1qBVpduew4qiTHNcbT6JgxA9QgZZnTzqqEgddlioLjzNd/Eo
893zl/4P6lFGgMe7uAWuFwQ9Ej6KHxVE2XFgg0ebyfgPc7Rk+gEz945ImgL+20nj
eA5I00+T8jfNhH8T+Tapkl6kWfwyLP6qMqnAc0EBADK028K6h5HPXpLmLWDPjhQA
K5cafziRSkTjah2/UJSvV0ju28YxC0yQxnkKwQCYNZz3U+61t8/BlCeDtv3RyL1/
4hKoMtTF/L9EFKwxFUBcc2wuTr4MveIDNCzmcLx76ejEtPxx98h3BkJIYu99ShjC
IA9L3VnQJMW6i7NEeVoIWWNBtdmeqdNMKIc5ijJtHspb8Ukj+qubcHP4kNwu3P8X
A9AM4g/XYJT7ys2Pa+/phXzKk3v4AlZ/wPKhQtPkWEpc2Chb4r7qPjAgWN1AkeHM
5OYqdAZfj6jkdP8Qtrjk+G+QCYX9Yozkyaz2j55lCm+dUvyzvcy+H3xFBhcYsykg
EXatvcHAfPQIXQ0rVQsg5lDdcM9ziXnoTNcv2vYxvN6wvvpNF6zxjV2knEZ0NWu1
/NDkL7PpuZlv35Bhi2Dlzmmm/lbAQhit13xZ5+yuhccxTI6ZuhKBgJWllhbIvTHj
daHbqFtezDxKMQLpOHDRECwpJ4CIdVrKX7/SU0sCxfz/y4Px+H9R1IDFHGIEc+3u
u8LP8otCNi4FNZ2aWCnUHeS7hSIn+wcFMtw6BmDNlFt6wwTrlkbnYX84YfRx+6ke
Wq7l6afyggDNi3kzEhOawVaKeZoexQ+D0VPAt/v2PqJtTTdKqrS6biovqalslFrQ
ol1CkPCKV/Uq7iO10wRX7OonQxMImq/mYl5RpcbTQBWSQJMjnudPLQ6bDMxTYcGm
USvn4u9FH9CqxFI2XzV6JhRf3cvcG6jp9uZ4BqpJ4u5NXeSGxXTFk2W3BrHa/N1/
rs+Qeb9Qo4jaBzr52dzvpUj6Orhh/vyPT9dVO3QaMu9AopkF01Eb3OuxWQKCkI+N
j6v9MQ7iGQs0CmT2aJAFIuYAOdGuzwkQvxOZ7pf1MLKPo0PyN2pd/TRb3WTKRQFR
TEJyyhWHD67G0JdenUi80ff1G0mNRAD3v311xTdSu/Hd2Avn6EMGIpKWorsrPAts
1lq53Y9G8nW2+R6GdqV/2I7wPOW3yOSwjQnEplOjES/aHZhMpVQqLUuwbPwl2YWc
X8toLfBVh+g6YhBc4eIDjyYadaY7FmuEJ5IxfoKc7HtQN00Gs+/a4MjvYkOdYXtk
ip6xHd7qLRHr2U29ciP2W4DkZp2zQLgbhi2mQBSHr0m7Dodd8L9hCbgdebiGAPOd
cK+sp7MoA45xh+d29rprfukeIwCcKNk9fT3kuhLj20ZDAkvEXURkWZ2+0jeZk0ZZ
iXIF33KeermMqY0osZH5+1eJAe0w0bl/u01hGhStd8oG0kBOpOPX3y61UbaD1LRd
AlZRumX8i2Du2D7rxI/LObFcHbmOOJLw2CB1qRXRkUR4xk34amxTGU65YOFOIgwa
fRJB/E+g+RywKw5KO5yCEpvSHoLv6EE8c5vZLEzmH1k/EvCvltGdd6HwR4ji/QzH
QC6m4PMlsV8qD/5wFd2ALJ3o3VteJ3fWPQBjkLYyTpT2QXNTGKjY868oWF/R1a4V
nPnR+wwnxDQ8EBywGN3PXkMVdx2OCJNzknOSxqzqdE6gPBs/7RxYrf6BvVXPgp7P
6kakg/Lo1WgnjUvTfJHL1dxzgHX9nHRI2U7J2zf5jFZKej9mfg6iWOf8+Tw0Xo0Z
CSCgLy6q4lGymY1pe/MhroPour2txYpJ7++kdSM+6JDcq0aaBz5ULZPv7Ad1NKjM
CQHsqShqkM7m0Xju7I9J3GqlK2qp+0sL8CmA8WkPPzeG68unQr72J/iQmji+iQfB
FVLABneGaTNAW72Q5AmgERQ6QNmje8sMAqPG0PopB56BrI3bU4+ZfM6iSiVz4QQ2
Hj0H+/Yc2przYTlBtuA03sqwRZHEtXqqLkInlIcI8W/TJbKWzJHyaDs214WfsGKB
WzP60aGmy4KgDUx1bUCIQ+6zD+oDhPtd5gPuiyw+RwBHQqhB22KhqY4JDSulrDsc
oOW1xGf2mD4IfVyjqaeeL4l2hKpWRM1dQhYyp9dc6EnVV5p6zc9FaS7HepCPYZRu
MEmQAqe5l/gP2xBTzw7V2ShQ5Ml7wWfhft5wVS1FzvFd1PLpNkpa+2tX2GhtvOBz
I6NymZe2S8uuZUg1dGeAP405K7RmWMgEZxQne96u2dUf6JtsavnjNYJzmjYnIffi
6K8Ey2HKPReu/i97MpE4n1Gn/AvVw3rT0sdfGeC32iNj5ZviW7QlxWgrLdKzpdGL
PUESeu0jsRa7UwnwA/CaQaHTdEwD/VXy2rMEfQ/CqbMcTwLt3cNfxcByEMjWIiUJ
43vZwJE6FH8LcBJ8+qVpHxZF8Zb9OUwbrXqJaHjGrwjLL6oZ+R0aFvoOfcMNRiA/
mjh7IbC4I6Z15G4Tz72ENkxUeBAAT/30hSHLRb+pnJRuspVs0q8vet8clu3B47uK
8OJHCw8St4ZY/Mw6s4ItTq6Uo5//fJE4mrmF8DWxyMtc4fNsyFDwGba2w66LIE/0
Adw+umvF5m8F0D4Q+uEYFWS1TEdTORKDZp+oRyJypDom0Xy65yyaaeGpBIksK5Ei
/U7TiungQ6phPlV4DRY5cjDdsU9SSf/l0WJ0k1bQnBNhxSNPAg4ctW+oOwP++HHE
tmnv4Z0JjN8z6heF6HwrLCkV9qwMksfP8+JSQ87ix/QVzA6h6MKkpjl0FtxQ6yak
lJ+rO3pBTmhqiGQpVzklET6oxSqEd/4tfaZsRIPFxksVZ6TH4uj6m4pYuYbv/Kej
V8f6rCKjxknFLZfwG6lAiL2behgWyylGuXcgEuQJL93akDKh5nuFmpZvYOle0NBW
DkFfhhswcE4O+Mi8Zpufd3Trli5LPgvwZwBHrA0OK5Sg5tu5ur5HKmS8djob2c/r
k9yRxSXVBvTWp3OhyUSDU/ucNNm6hhUB9ISIn/uMS+yTO5xjPMj2XG+H5znrVzri
4t+IANXwKkBk/gNKSqivTIEzO5W2NabkgYgEnnFhNjGFL7UZnXUQexWG5rstEthG
U4qthpTGQhniShg4M5R/Wgjrj6Ho2ESIhtXi0vkcRbCSM2bctF5ZYkvJ5KnWC+uY
dxLFKka2a8jycXNxKbX/lEZIYnwnNH6RIyhB3VF8OOeRhMOzpNG7JDxQAa/UFWM0
zW2WuloV6UCvu3j0yUTV0LmqQOFlLBfMtvbvMp2BiMXVFdylxMZtcBw9qflEFLMa
7y8MzVhaH/wwogm3NnR2ZClQQ3ogBfTHBDNNqwZGxvod2XBw4NnOdH+2A/SVjUWM
mEn9lfcMT+R37BnHlsOXFF/W1FzANoh45ND3kwSB47VuHbc0Rnx0p92qCwxtanXd
Pc38tEb0I0fOMW0gb2QFq9c6o2nZzUjT5BSJOxyAXxkgE+3B4W1ApkvQ7W78w/sc
28ElBOMzRlqUg7kjRQG5JhLs9/jLxQbqbcisD5bVjftN+VoM9tttgqeMObQRq/qE
/+VS9U5JADSiM/io+7Rby0LTkx2QRYy3/eNFZ53cITDzVBNvaQExM7JvQ0BehlP6
+gxFAauBcsVn8pm3iTZGyrvrjU94eiCay69bpEx9/SDtBtyyl4e/ET8zFfdA/0ec
BTNxlSS/+Ta+9x3g3D5BYS2evxrZSPGi5SVnQKa6cO6NqIb8WrqLUP2baUzG4HRf
5S+2ftTvMK8/oBHFmWkY9etnUenjgmwWThdsmWIGN7bkXUlO3JtHeOXtbygYbltk
RDFWw0wmhpOZmA9mj4ei0AlynTPYYZUE04FkT7HKvLlMkQxhuettQcmy03XnFXdx
jMIEqt0v9FwFs9eE+/gI0cmE4I9aXKyj68e/NsGKTyD3xAxlXeORnbuyYgRZbXjd
UM4sNNyubkb/EEbtNS5v8l7n76/xqNjgPctsLlAwOEnyPHebXPRNQxzF2fRU1r8X
0nKvQQE+psNuaoGq/IDCX5pR5DFAnLkGbcRdUUJ2RRmzbFuKWYOjHLoSkYAr2+vo
0zvbChMRin+jh+m6i9iDjBSe6uRdwOXtVFrMkhjQX/vRUrsGvwZYHdR4jLk6gTT0
YCIoYRuiFCNmHRWWsburtiJz1rE9LywUpbbIXqQrgtGtOH+BjUM373PcUUjwo5Xm
Dd55GP6VFoZCYG5CPV2kqyNJCl3nsLxTIyG0oZ4BaJ/sl2u31hMRbW+iNO0j5I1y
PgPaYuXufsPODnC9mphxwvwM7vyVpha5W1gGkgYcuEuLf8gtF6EP+vytcY2lf+yC
c62uGfSf0qQHz9euhSLGrvpXLrGSu09w+4wwF10rfEJTsfUFhJSpLzbHkvQXICzQ
aP8krOkVAsWDMMtj106rPBQIUAOUD2EDrnHsD/bpdseb9/zVZwNGU4Juqozy8Dof
2h5jiqTldTs7mv6EMw/qQf/HZAG26xLwxjFIQgFngEbPWLOZvzAw9QhkuBR8YkQw
s7e/sy3f/TbMz+A+7Pa5FIzX14YoaLq1UlWU9BGb4+SAhveVOYnMuG38vXW8hXrc
TZVAZmdD31TQdfRtg7aOj+IWEUjXgvn/mdZP/RjDg/q/vvB0hhF86H97DuQhzr1I
Zhwk47z8cK5zaDJnyn5kA2PsWSdkjtoxd7qBMYkf+Ts8YOYEfgxcHsUAElH1ySY9
ccomhBnojsD0mcATbWw+QNB27UoPCNFgEETQipcTFfNV8Z0Rn8S2JxPc2d/wuAsF
xDxEHjyEQf5Hnl4ZoqFdeLavFzsD8QEIrzG5t5Mf+NKzs3LKe4HODu1jE8RvK2OQ
Wj0Ud2QNj8jn2xMMpTEu/kHe0QLLPP8ybS5/sHyq6UCZ2Zrqx5wuCVTyzQ1RlX2l
ljZYEzaxEtXx2HF0Y/CPBw1dIg3okOHkjdeVMt4gSb9lWPE7Ao0WDg+d/DhWJ0Kt
GX/MZVW/CJKhtI9B5P6mBayfXrQPhFPMZuCfBcFBcbUyqUMbVcxCaZ7yykH5F5Mi
6YX/IbXSyHQhUdKPzDALV2nIHECUZg2Ltrq3IP8ZjB9UXZ359wj9zPKOoRruvNQi
1lJTavJpl9h3T7zC0nvC+zrrRmVSB9F4FfePKUhNdDufHyzNlHjgNKHGvtQoqhM5
nW6qc6o2j4xiE9YXNgkEa/Yu0bBg9rXyyNG2ahpxp2HzZ+aEW/Y5YLbSU5oo1i0a
PHxPiSHjSrQ9rVhbdfb17kuckY7ee/CEZT0ZiOlnjcnsxtL1B4hfctDq/aCOT+bf
/aKarUEcId1ws64sDJqhX9ThgxgFXboEt6GAdM1asyOFH7J3N9u5z++7ZUxcQZg5
NeDxGwrCmrmFAra9KEuMqZ9kcQmrhysMUxgU9+9bv82t8Gw0xAvyr1dqD5jK5xyd
nG+sNW+0CKznfDA7/iljx2ZCErngvfZal1bHftXELgJe5in9XXp9rhQqvMtZg+K1
TxPED5djK9wt5mfYTBzYAQ274tSIt3jIKsi7kBPy6y5BGol5zme5R/fxMl7fPR1b
ZGVTqtysVCVpioe/b2O7QQIa7s4U9M4J48oSIvvfuwah+cRut82CWZW50KuczJfO
LcMLw72mRL10zHXmLl7YyJZDXKrgnTbuhQVGEqEg5s5jdVSq4kwYSKUFONsfoKXW
IXPbTsmx3Bi5kr1hb4PaS1XDQgyqklbaffi5uLOk3pSCWHP0+L9xzMrjnR9NsIfj
lv+V2oRmpXZkW/5+bYqXotCpPUhKqcVSIt0C50b0QLoWyVLc89cOQ47jlbK9t2BS
8W/XJDoNMFRJb5ypO4y1QUGOQkVomn9l/UfK+9BBpx637K8pUTQbSN/f8OZGnwB8
htynIfEUhwlbvTmESsaO9QP0VuYEZtSkETbtsXVOrRbIUUP89R9QZED/KBs0XSjE
Rx/bXDeWImREYOnCRHDvimQzi4BJg/nCnidhZb9+baWGsgejYSsEP0yIvZHu624v
KVynmzuHkZrNYr3hvtcq2HkzU53jdHVz/mXlys5HVMIF1JkS4Ji6UUs+llHPnkd8
HpgV1TOvHScP38Sr66IZBNpv6t9Uzv+aH8YxxSJWZKiasZd/zJV5Uezd4Ty2ytvP
sw4AG6ItdEwS2pf+k1qORA3pTEjo/T+hiLpvgzUI+hbYqLKRQCqECu/fBIJn/5er
aT1HhdWoM5yah9iif2WUA48X4CRJZKmJ1vmD0lObhNVN6OmRxGYa1P9Rb7+h7AI5
NOSSTZbqWsRYZlZTliGLU10gW87B/zZb/zyA43niDfLyUpwlA9DFJ6Es7o9Lkl3w
oTWUhTnltsRFfpiAJINJgtn/R0IDAxxasm4amd+eyyUlL5TgpaByXb9ZAV3dcMxv
fux2RjYIyO7cvPjUZj7uxvFZtbootNs2wKE4cn31KO1W5LOwnz597TE+yHZZ1IXT
2OBd4A0ylSNxK48b86Nt2flLy7h/A/N4pXwcNzEsaUqv5nPm9Agp+Xhux+3kjwIL
5qOKBASH5b7wo5tkMng5ZBCjFBNiOm47wNOsq0LAukkL9jaqByxNVniVt1Rrax5R
F6ceA8P+jtOGY5U3YA/YiUHz6/lrvn9p1rg6gpZPKQd/LdiFwTbkwGpEhfnlz2/u
tipL8F2OMXn6xx9+E57A+4SDiRh05osOiZCcZuoRRPnG/qwbYZUomKZ5nsw6Nzhq
wlmg1Ycxh2Yhfg/pRZIBn7bhu3ILvzmGd7hxD5Zx1d2FnhA+/R6KGhk7AEc7Z55q
4qjXxPARHaifA13pB8CWMA9hc9OZzNWRhBJu5RT9I8KztggFZ10VlbuyCNT9eX/g
0EF1fY+pArCZyLns4QAOBD8KQBoA1xlj1dL85/R9c8opfmF7Riv7WgGkfSBKC1pU
UgK1G9lsqhynDWIQRI+megBB8K0VKhJZulXUNytYetcyVoq+WAWYsnNzOn3jc2fv
LuHlrrflPsEsBhxelm5OSNXs5ISnRsnhDiyM5f0o56wDwDYo71C0N0ibM+4fJHi9
/MmCRjetRIeLTREfCJKXY9f95abXaBYtdJBPQRnIRvgqxdfgS8kxXxwyI4Rczaaw
NJmsWG4ILNmCNdd88KQf+oXE9XybeVMjArea4hDY0lHGVBxtHJUR+Y1sjqn68Dsh
mO5RZOuagYDrOIp7hOa2Fj0OSf01B6s09aKjK8fiKTUqxrrO+lgiWi648hFob1Yo
vBPEsGQ0p2dbUq010tPEDnMTihwPM/37LKlRSNAX7r29Mylj7zQbq8Gn/7ynqk9x
90zo6+VfeUBPoPFJ64yxZmKY8llk7vxdzbeggkHfjlgxbXT5iMBw7rvSjCKrln+N
a+tzJMPyI0FffGfd0AISWuW2SvbaZgIjeXDDejwIV6XNXx9qhvjmXzUrbUAOjpki
fCf+g5G6dOoRcfUcB9ZsA0DE0c0VYoneMK1Zjy1g42R2SJtN8YNX8XrNXrspYnyY
jB8nHv3w+j0K6hVfG2bLnu7UHu9xpYC7MueLCLzkbPvsWJ9ZngCa6xfGWBYOE1+O
Ho9E7yMi2q4rFenIKvjKbAyN5umgPeIUi9tsn5PkgG1hWLRtQdeeUVhAicFh9qWN
S8FtLbYWtPcP/rXJIEV5iORH50JYaiB8qT1Ck5Xxomd+lD4BIugHPPfVsRgbA8SK
PV2yrUOy+K0dzcwJDgdBaHlgox4VatLbsc4DTZOGRQO/BPzvIHbinERjqO53WmXg
05qqIMyjbgFZhsT0SVWobuKVWFzk2+AfENUyxneITUqj9ewTehrXnIBcvjszPc8c
8WAadSiz5kSVGCSSG48LykAmJOkdU+UDSto/xjADF5cUZv/svCD8P9wIq5xgW4zt
7HQL6wvhc14HJVuygC178EKWfHlVhJWgRm+wMYgPfDTkQK8ldnhjzIxwjgC6MOeF
WjTNzWLWkbIx9q7GBlGU4/V7KXr3feVzJR/PT26Y3Qrf7PBOryNVYQ3HgluaKwgS
0KZeGwF0Cw0tHI0fuS32mrbrpvXcc0qDCenXdgR9ncQyzvJzW9rTWp2qckcMt4dP
Wznu0RKuN4M2G2VwREXO7QI3kkzGU98Tzdj8QVCc8BusybzP/3XNWFgPGlbfuDWu
AA8r97mlxnTJHOXgFKOS5zEyaQvhrll4WlaGrNNk1ZgTmjbzc0IeF7lNibcAMGvL
S6GhZrIu/mvrEF/oPnxB3PlZCQZk0zExqNRJ0Iv0vOThZa/Dkzd6B+fa76tYaHTh
IVoRwzCzzlBDIwWvzchrlz1JyGExej7Nwl2kuqtzwUJXdO0lPPYsGxcOA4BXSfHS
+1ArYQA0E9dFNhDuaEoxwHf2VaVqmtj/2q8CU488JipCJRBPP28Hl4W4RnGvb+X9
UfVN4x5wS4FkGn7j7dwawpU+yfCz2mce1El21ws2IAbp3mW3mQpU7wVOBpOKI5S4
f2fxjUCfTszoBu3AVWB0BiohVAzfQq7yN4afN9RdQFH32pH5McKXgw2UlomA9TOo
2pgFjPPwvce3ls0o/FIvaxiF6JpnOnKeTQTPtxDJj6akAt6dL0A2vahKBQX8z+4J
N1zMRJbiJS9sA1OOicfDH6N7Axi06ufAj8D/vN9c/bIXjw/3K+HQOY8mHo/xtyi1
fXlyghbh3eHlCaxcknnFRzdQFI21sh6ZbLqKuf2VogQiFjqsZkBDhqPb9bB4UJLj
068ax//pXs759bwbHsd5DHr2PLD6PNXw1zW/78HqT6jJOkx0t5eLP1CtRE3A/H5f
KwnDiZweT2FRhUXzSSFBNQ5gvMR7XJA+ipZAJC30OjyVreHWHPt0gRUPZmQC7pLm
03vSIy692Ox/dRQ8pm/xo6ckw11F4cq+XbNs5aW0vINaJypAWpzcKVjobbhExhs/
tiQBpbr+zZ/pt9oMK30hWbVaUQpKWWk9zSqvzFx+OnQ=
`pragma protect end_protected
