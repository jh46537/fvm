��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&-\X�ǅ�2�.*(VuM_J���U$�`�ß]���Vn�A�1�����)�}��
RZ��)!�vc�x�\/7���mi{�l�Oj��υ�ª�W߄�JA�;��'E5;�%7?G����Ǡ���%!���ݑ����f���K-�c��	�����w�MF(�bW�.��'s2_>���ǀ�cu=�J��<FRY����M�f���:���y�ƅd�sL�e��m{��C�c#��؟q���)���R��7��aq��̕#�h?UԗCT簈;��_pNb�lR�Dx��SO�����G�Îq��4$[��0�33]�1���.U3z���T��[<�����f�C�5�\���"|l�t=JAd�xL�i����
2dsߵ ����C�'sZ�ʚ8����rr&ۘM��ث5H��
����q�X��p�V�������(�~��BS�z��%u�%��7;����}���Y�l"m��?��|�TS��>�$�E��̘�FG��mЗ�[���dŷ�o�hu���V��'A^��u9鸄<�/�n��.��"�P�e��NBc������-ҷc��G�u*3˓Yu�V����3 �\w;��/Jۃ��d/�#��zxK(X�n_]��`0*�`<���#*��e.�/���<Q��\�HeF|���K�+[��En��;�R���JT�ˌ�&�l���q�+B�]�p�n`r:���Eyi	���
���lE�{�դlx��!�پ`ϙ�iդ��l�G'��R�/��}& �P�[�ӥ�@H�(
�{M� �3uc�{K�#Q}*�u�"�$'���3a�s`���$�7��T;#�H1C;lƿ;m��4٘@t&6Y�zgmq�?*��g@S���;fzn�Ǎ�^����-�HiHQ
-}�?mK���%�:����pM�L����Mٮ�<� ����ѫ���w�A���#���e���0ϣ� (c�e7�dz���By>�c)W��K�5Y�!��z-,�Ԝ����̞���$�_:����\:������Djd\�+1�g����6iE;���7�=�Y�ԥ����]�:�3@C0Y�[�)�&��n`���y��!��H���@z�%�\K��<���z�L�҄b��X������]�-�5_%{������8���}��0�����IvB�?Op-�"��P�*��癢�X�^K���i��e�-e-�h�����M�#�1o@VqIR��jr��� z�B���J}^�`�)���
�D�lJE�zzjb�\0��n{�fh�eM�2(:ȉ�������{�UT�[O�g���V������r�S��49���P�p9NB���h��C�ۡ+�C�u%_�.�7�@����z���K�+X��iX"\!O5���	�6B��+��&<z�DzR�(�\�<����A��Hwq�\m������H�y��Tp���B��Rӯacj�C��+C��M�p�� ��Ky�����ʌs��{�����ԉ?)k7ݒ鱪�PAlB7-7��k00��k�LI��,t��"}y^��}�)rLƚS���Q#G�0����ПЗR�~F?CD?*Q�T����S�*�dcdp�̊���Z_H�\3�+�
鑝��7�� ���^�,�&8~���C��S_�t�i����d䞧clb���.|�w�#>��Y�'�(��E?�V`xZ��M]�EsntC9�Q$�;Z�6ˣ_�K�3�D�zx_p)�X��7k���H���yu*�MyNSΚ�X������:�<F{u62?��}E���k]b����ן��.ťl��UKYC�P����)�	0D��ġ?���F��-��·SD�R��&\���<���� ��;��²����~��$ڪ��4V᯺�㵬���ER~Z�C��&�*�)߄����z�pۛ�V��Z�9%R�^1��ߑ�,j�@�GFɒ��3�,�o�4z���kZ}��p���*�^���EV�V6EB���;����`,�����j����
a��C5|d�O�=�SY�[���юԀ+�Q��7�t�}O�搡%�I%�g���Y�� ����=��HRc��Q#�(!��*"�=d�8	w�y-�uj��'�N�?RhE����<�0��f�1���Y��]��m�vMv�y\��� ��1�oO�X�5���%��PkB ��E�6_Q��=�_� oq
��Q�Ǉ����qz�lC0/��?�	�x��z��x{m�EU	�^�51�n�4$�!�'(\Jd'��9��a��Z�E%\]\���ܟdq6|�PZ��k6���}f�ۏt��e-������ͪW?t�ӯ���4����3y̿�P/����Yy}u���y�mA1��yCN	��Q���ً�hG���f�	�N�+{��Pt�q`O#K����e��1>��ڱ�[Z��d���"~��y�s'�8.��R'��3������=.MNV�w|"cC����;�?q������k�1Sy=���UA09\x�|	��>ݫp��0�EQ���xʃ�F�	�|��Xi̻_�ͪ�B� _�n.C���Fv�h�c��>E��{��A���&1��Q\?��^:<}Th�V��M��yQJ�b�� 	y��������5�o��Pd��ۇ�9�^̄�E�F^)�E��)d9�RY�Z�`o�U�j�����g�(w��f��hw�钚�[�u꧃Ba�M�ԍ <C)>vF�Pe�ל������[��4w���{L��jŵg���}��?��ˁ��εX��s���-=�I1��t����)��w�YGf��˹ i��ET����^kB7����_��8�-n_u����v�#�*�m'@���E@%�[���2)��!���^���Y������A"5�y_S���(�1{n�!������z����&8>�ܭ<a1&5��r�
P�z�-��2F_4�V�E��$�u2A1<�	t�lb����-9�-AY�0Wg3��e:�T�AǏ�$��N9��m����&	��Xm��RGvO��,z����+�V+3�A	��_��5g�{'�@|[�u-<�5\0��KW�%�N����>���ٳrv�T�ʟ�QoI�4a�EP$n�B�K��`�J򞞽S��0fn�ښK�v�G�����q��ST甾N<���U��{k����\R&�B��$g�"u��2M�]��-,�� �}���I�6���%	�/`��#��ֲw����×�6a��m����*5E�q��'k�O��!�o&FDD&��^�syB�?� ��c�	�V,�fZ�er8�w;I��m�#�����0�tXJL�������$�1�+;�Dp��@ �:H��ѧV�"4��@L�l���T\�J�žU��g�̗�KX-`j1J,�_�GJ'���ɂ��K�Q���,��VX��0S-9;�b�i�3)���J��� m�����T$ j��SC�=�����ο|u��	�;�)LJw�9i�\�XDI��Ѕ~��Ƙx�}�f47��=�����;�-t�R� V�̘`R���a���~���`5I�:�t\�p�}�Ӟ�|r&��a�����D�\�]�!2���HC^n�y�ۿ	�=V@x�Q��7����k���;�'�u5[�hL�YS����iP�(�P&������>?и��N�^1,�`U�c]A_�y��z���y
:-��WEVi�����C��
v���y�'S~&t����h1ޝBܨ�D~��Fq�+���HG�c����4�i3U��ɉ6�R���F9QI"���2{M*MݱS���?���N8�0���rj���|���op�,�G���`���*֕�ݙ�J�T�Xs�:-�Qu�PM��9���6d���q4u� s8m�K\��$�f�fVd-�;��� �#���?n�����yR�.S=$x��ͧ/V�,g?��#���6�Uc�*;�6�7En������t���%�����N��x���(.�w_�溍���.ឥ%�V�O�Ն ���_�!�`l�R4�Z�tv/��a�Ź�O�W��<͖���CH�/o������IN��1�����+>T�Ч���J�J	pl�j��|�8;��gU�3���Ǳ�	���U\�"f� ��t[.o=�/Ul�;?�8[Ķ(wP[��㉥� �ה�c��{���u��s�0��y���+>ym��5N�d���q*�悺U��^.����P���6w��C��iS��J31͢�j�"Zyؕ S$>���}u)0F�?���}�75z@�ݴ�y��� \�.i��iPl[ssP����
RP�~����QQ�)�O9�#oq9�sHf�?$�{}SjB
a~}��>��RgS(H���	��m#�|c}j�o����%���M/��q�m^��T�~�x#KI1�cFYb��Ѡ���!�f��&Ny���e�8��m@Y|mJaQ�р�T�D�C�4c�(p�=���<���¦<�lh�T�Ҙ��1Dcѻo����GЋVpCYC8HX�i�Q��2"��Ne	��u9�04��JR��U����
�b�y��$u����?�����y;;m�1�z�%�K8�� ��� f��I��?����Zr6����[�z-��|��~+
��YA�0��	*��,X[HG}4���0�&�	U��!��&y��@��U��b���ťkɂwJnk��p���鴘�K9��}��&R�n�n͙�H����$��/< YEx���c��.\:?_�U��&����0�����󠥬-���2���Џ�K�d��/�ϔ�)������b i�*�;�	��?<8t/^Ri8��]�lg�w��U��lh%��c%�E�ΛrI�إ'�����h]�N�!��Jj6�#���}r>X�sngS0O��;��P~������圴�U�[�x+� *F��C�F�ve�7W'�
�:�z@#kˡ�x3�`�Nq��r�&��Ο�����
5����'U����]L��R6�8��� 'h/�S��h3����n&�k�u��s��W:����;ڴ��ab�䢍u@���ȞVIz���9YL![$�Ow�1�a��}]�}��238�A�_=1�o`zH'*���=��~ba6�?>P(�K��l#��U����]���pI��T�w	�KK[�ϓ{������O6]�Dx�)t��b4%�x��=j�Ŷ��{���G��և݃�����Uy�h��F'��y�%��UFE�q��!�����<?r�%���H��<,8���K�i���Bo��Gv�m%V�,���mv�k޴]J��OP����E�����*�dT��{�N�U�}�t-�in����m��k��*	Q}�;�ThB`�u�9B�a��ɿ�<<l(�C%�c�D�_~)$ ��L���}�2�{hƈ���d���7�f��G�))�E��b��?��Dp��{$���$�4Qa����x#�y�b5�L�׀�|���vq���n�G��nċ�8~g��E��{鸪
��?<-..�QB�?���e�U�N�	ˢQ��m%�!a�U��زy�����.�Q��u����u�װR�'��Y���ě#X��7�))�U��J3j��q&S%��H�|���`��,��fx��
_�w"Yٞ�	��W������6��r�Q�&��$H���0�u8Xӿ�V٧J۳�Zz|{W�UZ�!�7���v����){������U(&<�vC���x�8�Ȩ�wR�ɨfY�=61y�k��NX���$��~��~��80�a����E��O�I���A���D�n�k���l���
���_x�DG����?��k�P8�Af�zI'/�xm�v�:�<��qZ�俻��ڂ>'r���6�_�w�&՝Z�f9�fn�.�z�)Tś
���m�.�����ia��O|��f{�S����(�^4H�@�+[1�'�Ё��Gb?�gկ���Kf�yPN�������r'"?N��͢��G��^�K迪�#n.UOR���T"�U�;";2�u�|;M�͈:'J_b���  ��T�*/��[�k��\�zDFͅ��n֍���X[Q�ϫ#����ä6�b`/"���k��Rwu�L�\ͥ��FKjt��¨u��$$k=��҇DI���M�K6B�:���i��F�z:��4�ݯ����������D�fd+��K�ś�4X�����<Y��$.ր#QM�n��k�md�>�?�|�`w�Q)4�p�o�}�	�mU��L����b{�߄�tL��=(IQp���@��Yg�K�2�I��f"
�bɬ� ����;�HAX�(�,��M$��?;�k RC,w��@E*�zR
G�O���q�xA4w�lg��hצ�8�4z�6����z_��C5����Mq��ٹL�G�g�*��&��9�e�DU$�"Șw��k7��m{Y;MS�?&�+�,N�<�S��vn������y��1S�t�7�f��,:��^:"U^0�{�쿞h*�Y��	��Y��ZV�f������,x�p%`-��Y�8r��?���]�����1!�}�UR@1��=�р淚�ʠ�FC��닙-E��-N����аےI��h�����9�āTәA�`9�}$��ܪ����f`���b����4�<:�!:�����OCʂ�?Ӆ>a�>zqo�>,�V��;S���!�T�pA�D4��I�h�:��w}麓ӓ扢$�2b��;!�G��T-:VW��@[�=@��PX�׀7	TS׍��uo�`}Hk
��`o��p������[���l^��f�I)^1ە�m�dN���`��2��x��VbdRp����$���zmpy�lء�Q�� �o��5�Xԙ_��D�|��D*�:�z�Ξ�
-������,e�I�?�紈����K�f�S
hm�rN�\_����#B�2����Q����W�,*�M?�t�<'ܤ��q부Q�+���e6��V�5{��	2[v�bXƔ��<��`V�j��~<�������2�xn�~M�*:{?���ݢ�Q�H�u
����04�ϜH!�#?�'��K):gL�L��[�h)eA�bv���HN��*��{>��U�	�o�f���?��/�4r6���il�Z�f�N�"�r����G'�ӫ��/ʣ��Dh*/�4���d <<N������0�@����7��׃C0�j�N���H�$.�:��!��GE@�PGҰ��=��X�`��)�����T�s},����{�ak��0�,�l`����0((�~f*�6�P�m��|�M���Q��A��%�PP��z `��؆��+k��:�,G���iP�Gd@u7L(j�Tz?@ߛ�TwV�i���*X���0����A��C3�ܡ�����D!���m���3��_Tm�ͣ[�\ȃ)�YX/���?�z��1��!LV�[�t�r����b��$gN�Qe��FEc�)i��T���n����+�Q���*Aa>�F�J�Qx������lib<ŷ����%1ZC�4�l�:-~�Կp�1݇8�ӂ�Ξ/ٌ���. S�֔��=��e�e�/?6lP�nw���k��1�	��}���:�@�~*=HD#��aY�j�~�����p�h�i�)\�G��V;m/��+�� �����{�h]�ɟoj����f�Y*����﷪9!��%σQ�S��Á8om��E���v