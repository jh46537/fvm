��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[��]�,�����X���H�ѷXF(v t�V;�]lvTH�sF-�zt��:��I	D�Q�+����L ����P�K�V��4�w����8zk� A^
�]P�8��r��*��-|Y�7�� 
a	U֒�n�!�ӽf ��p$ҕT1�"X{M��h+��#���nM�^l-�K���J�;�S�p<�&V���f�l	�ƿ�������z���y⩖݈�AR��+�YV�:�>�mKH�5ч�����ឋ����Ǽf��ʳ以.}�P��l��7O[8�xPp"<zU��\��F����7T-��y��.zFoZ��i�n�ˉ1���CY¿'[ϩ��Mt|�F�M����B�mp�C'�N�`b�%���>�ml�7�:�(%��}���N�KG���/oz���W�C�A�5��b�pZ/a� �N� F���])	u
�YԐ`#�m�(��ɹ�x:�����A���%M �~�Nd�0�s!:��|^w�����i�+2K2�|uء�0���bk�[Q
���p���%��{HG��6x&�����?��Q�]WՒ�^���ز$aϙL�˛f'I�n�uW��]��?�v���`�����E� �(�v�	��Iv��*��*���
b�Q*�gǱ��F�#��U�˯z�V}���ÿ���������l�Hfl���|�}PW\1]�S�S�+VM)o'�s;�#n�@ώ�vI_ �A[\�#��)����ذ�=�|{D��|j}��_��JHR���ድC�N��+P�m5�`~��O6*Y�
.��&�}�8u��fۂׇqb��缣f�rRT�?���r߅�cEY1CE��7e�����z%�,l�E�E�9�ə�������I?�|�!~��'!XK�����+kpq�b�˜^(�^~in��P�EUfβ8��6A�q��	�$X$W��1f���"��������?��H7G��Z��3�#R�d�5�׼Ϊ3ev�^9]!%����N��r<?�l�k����8��vy8#dB�F���YD�M���50Ɣ��:b�*��i��Wӳ��4������m�Ɲ(I��akf���7e��d^����r5�_�=ycqbAn�]��jlX��׃�ߦ2ԓ��+��^w�Ǳ��5�ja�U�%z���DȨ��ci��O��޻�6 .����^b�#?��+�k}O�T�&�xzy��%������v���h�w�q�!jһ�����z%��(m.��J^L���nxD��'���?�Ʌs�2`E1k������?����~R�k�?�,p�=U���ӽ�RO�Մd91̪�5f�/x���� ]<H�-9��u�����|�����Z�{�"��=i�oH�� b���3N�Q���s�l�Cg�c�\$�@�֯SA�@g�jcv�ڔI���E�*���RI�w���CLE��{��BZ��r,�ͥۈ���?w�b^צ2`c�0�EB�����3���ڽ�����qJU����Q&ڤ^����C��)Z��$<� lQ�A��٧�B"P����#Ӏ�6�%������V�Â.tO�ZW}���-gr�Q�y�[��N+8�Nea�6�JR�+��FJ-/q~��U���B��n��{�N�٤I����t����CüT�{�3c���ܣAN�,Ի�
w�r.U�z2��Xn��3�g�of%�<t�p��ޣ�s'0���M�����:�����T��&��x+��v��ի�vמ�����Fl+Iy��ec5ß c��۔-'�� ���
T��U��趢*Q<�$�Ѩ^W�p��+M�z��S"i���-G\�K���+�CO@ٽF�%���"�U����ڴbbS�rϏ��� �-�x�]gX�4�rւm���H��N������
,&�/y:�����fSa#|�Ǒ�h��7�"�����=c�#�b���{U�����t���s��>�o��K���h�4�PZ�@Pk�L��ţ�<°ӎ�o��l.O�)@��-Y%�Ӻ�鉩�*�O~�`�LCw__n{�-:E�=h	����Ɂr�Eu\]QtW��
���R�г_$�� rz9����涥�V�]�6��E�>7��� 4���W=�^
[!����*�TA����y{���s-����Aa�K��{����-	IN^��1��:�x*��e\�`x;��Z(��j0�#��>����DPqL�oOK����/�G챆���?0ش_�Ґ,���^jI ����H�^~%�Z���tV�U�����U>ٷc�*|s8oگ؍ǣ��*yj\���M��x�ĢS�s�Ӫ�XQ��f���v@(o@#�p��ũ��Sho�SČ˾�@�(G��R�T�v�4(nw7>g����� N�����J��B��7D�*��dX7�����:R��	6�a~Ÿ�<1�ޱx�����ƴ*��g�%�s��.J6M�ނ����d%��;��%4�I�%�en����� ln���9�w����� �s�Ğf�����q� #pT�^���'���?����Q�t��a����i��.~+�y�&���+�� �sm�y�p8��s�<w%��<AR֚�t�� ��|����I��mb\P]Ι�iu����iG�h�A��h!���Z��2�3����t%���l��	Y,�o���g��Wƛ�Q�Vw�� �.m˥,�a����(RI7�I�jm��[vny�y��q����hv�f;�N+�|4<$J6�����'����#�Z�B�s�Y�gYH�f	�tǑ4RCQ�w4gbt3�JM��zd�岌|�h���/���ǦO{���^�p�(Q��k<�������9�5��|0q��������6%�J�9J�涹=VnǛ��}��
(Ι���#��P
;�H߰�'h�w�煼�,�a��[Q��ܥWT�v�[���xHYBD���o����m_d�8��lSu����~�}A���~�ch:�z��;�ug�Amȍv"�-17R_�10��2I�τ�4��L���7lL)�]1��}���w՟��|%�,!�쇡j.����j/��y�m�to��9Tj`?�3m�A�<%�l�_Z?���7��D�Eq;s��g��z{��WW����H?W�N�3��-���f��!��~q������.��A��V�B�'D������{y�w����\"ʋ�@�^�y&>E��@'�*z�^5U���o�OS� T���H� �9�ǟ� ���@\����g�GXZ
�qs�sڇ�n�݃g�*�2t=\f
V���V��,-H���J�4�b��>gÆf��LC�g�]�	�zɋm���D����(� �ҜXUʸ�Ԓy����B�[gH��])P4�fP� ٩��`
�ӑ��q���x �ߨ�/^n�]��'u��U�J��Wr�[E�4� :���u��˱�>/�E����j\�M8�QF���v�v����Z1���T���!��.R��M�P�m�rD}�t#��;��y=���*��z���7�Ybm��|dgR*�?I�!$��H�h�b4&_�E���dBo'4ר��p/|!=h�1� B?{����y������~���8�����5CI'Z�;�o4�f�|!�\Z��s|j�@���d�/�O�	�\(���U���t��UsQ�%"Vh(�' ��+rӗ�e���b)���P|�)�<��������	�+�a�����c@ٰF���ja��e|޴�4���R7��d�+���esB�����b��g��rO��t�@K�Ofk��9����,lV�� r�F��[��$��O�c��.k>��mT�a���1��s+�9MDkH�`�}�8;���ףV�,��f"�I@���pD�@����)l�؝;�E��i&X[S����Lh[�D\a�u�����ju�h�АR.�����w���p������MӀ�8*4G|ye#l���9.�Fm`�p��1fHi�ۮm���-0��Ķ��h<��[ŕ�1 u�2���MZH���'X����9���9dxt�,k ;�������F��d.��c8^��	t���#�L��,�rܚ�>�!C.�2��V��z����~흞qF�����96�� �&Xj��}�9�oA>��!ٴd�<��6�woCb�Y�U_��쯆|����EF؉��'�D���-C�.��9�OP.j�-�c��� �y��A;��&ztm+�Bz�kN�J�J����� �H�&��)D���]&2	�`n�3��2
1��Y<#�y��ׄ{�yL�v�,åW���n�l:v?��L>4�\� ?����E����Wj��G�3X���F��D�;�����&�G�\	���/wo�����S�˯��?m{�HȴNS���kC$%N��@�ݭk�P��Yz9��U7���rY��.PY�@���<JC��H.�+�B.t�wG)�e�s\�c���gV qIX���#�څߍO^{��B��o��;�v��ڦ�P�ů�I4�%hB5A,.e. c!RL��{u)9*��.N%w�*n�u��D���4�mjp�����8������A�uB9lq'����l������9�T.���j�_�CW#0)�i�w������v��i4�a���$�q������v5#�:���k�<�ؼwC�˱,�U��
�w�(���|�w��eԝ��0DP.��@��\'~��e� +o" S�޽4g�^,Y���ވT��;S�F�����I��?�`سf�ZX��T=n�R&�j���Kܤ���������s+�����
}��jf`c�:&S��g�%H��7-!,U36�D�ޫ!]�Ʋ�S����Yh�0��.t�;)ny\gj�r�,I���T�9�Н�K9��U��g�u��N/����U�^߈�P e__��䩇P�}��mR�b��{�i�ݎ�&V�MմYԁ�,pǈy].���}�As}��9
j�9i�� U�6�FnX�U��@
-�U���+�Հm28��[!��F,O��m���`��~��4�=�T���P�B�����%�)���t���Z�Ǹ.qˉ�1��
�E�h���-7����X���U�f�
@KA��d�G�׃g^`V �hn��*�֯K�TZZ��wt�Wμ���;��z���bo �ݨ�xW5QA%NXk0L�?x{�ă�5U49��WS��0n��-���q	j��fo~�Z��1"��d�j^��͔����i��4�LU�q>���T����pl�,�ST�<}6"l����]$�m��iź��d�`]YKQO�O��P����E 8���̆B�?�Z�N�pl�8�y�=��x�V��=��vf��p���;�3�/YF��He�o4 �%�`ag͙�YK���7x� ����.�{bO��( ���w�E9�9Khߐ�w. AM�dTq?�o��� ܑ7���7�J�B�K�	ʅ��Ȉ�m�[ٙ����2㻩,�owm�D�i���۶k%��� �H�bl�.-��:�RJ^&Tq.x�(�-$@�bU���A�͠a��T���}�J�|���^�K+��0Y��v��&�A!��A��ɐ�X?�=$�(�YkBz'�`Ţ�K��*ed)��h�>�)dv1 egQ;]�g��GL���ޔ�}�:���PLG��s�R�3�j����Ho�d�u��5A��/�"�J��Ϝ(S'8���R��pa�WP�4}�x��褝���ȸ�wYG5-�.PI�I��+o5?�g�����7���5�k^A��`?�R�O(� ��W��m1�����a�Vϣ�>?���I	<-t᫷t_# �Ǘ�m�H淳 ��x��J�� �d"s���W^*�f�N���0�C��`�H��(s�P�<��_����h�j�xA�:(�x���άZnX�����x����������iy��in�6���H����v�[k6�T����Ȥ��{ޛhT��io�o�����>��;ie�`����W�	�N��Ձ���O�7�[�M!�g�ڗ�H_\ޑ"0䕼�	4�y��|p��HdT%�̀�'�t�U󚩲�����Y�aiH_��"����^��-�����靕��N�IG��;�:>�$�����}���"Xy����f�:����&�s
'9N�k���fsg��ʬ����̌a���(l��xVN���\�˥�_w��z���I�c�ݏ+y��>�ᐖ�Ŏ���(�4P��r���s @�+���pw~�G頹�v�n��,�[ab�zLo�*Y!T�����|p1�c�y��lBi�)��X�����c;о�� RJIja�45�mE� ���y�5��Kt+z#�Z��Z�����jxF_�}n�}*����5��GM�(Zd�v(�{X��?b�#eO���1D�I=EZ�_ƪ�<�㻥���j� �(A����O	+x ��"���cz�"�m��ɛ�E�����(�!s�1�D7ᅳ���pe���ۥ���t�C��u�z�Ϳ�˹ۧORAK  �N��aJf�t��'R�KN��!�4T���"��~&t�d�:N(-+AXl3��?I�T��],[a�&��$�N�
P*I�@y����p�u�Ś��>T�Z-�{�͸Q�ɜ/�����9a�#��.�c��d-���s� ���¼M1�{���#hT���D��!b8I�tA���##ՙ�Lۤ
�e���Ҍ����Ƙp��)��@)�����BwP��4y>�\���?ٰ�p��!D5�����E0Kcƶ�K��7$���C���Uxc}2�����'k�,̾q��VefXۿ Eg���f�^�H�}�Y=`���q.��U��-�6�z����hڇe�7%A/��qZ�"7�[פ;��T�z��y�|6 �b�����퉒�p�;M�.^��=ꅮ7+9j��Z�+p�Җ�~�<�Vz�0�c��V��Wr
����Y��D����+���h��(5b�@�3�iSw)���"e�V+~���B*ZdVQ�z�3A}�oO��yD��+Ĭ0�gϖ��f�m�Ϣ�e��(=�O�rZ��>!}5Ip���V��c�����2�h�ZI��r�
� ւ��B7��cG,ߟ�L����������*�o�x�����I��ڜ�~�k�/14�)	:�v�1ؚ+5�%<1�9��3��k5�Rp��H���0^��uo�G�7�~Q�.x0n!� w�q"g����K��7��� �=�����2p��EQ��>�s��3�)��Xw_�-���K�|e�(Ȭ�vn���VS�� �\��l	�H!��f�R��PM⌉�(�wJ�:�����K���ǆ8�̤��Ժ��?��aر��l o�]��DY���w���h�>����������<;j� &�'R�Yg�#��h�c~r\a8�g������«�`3`s{:�&�@DC��c}áw�zFQֽ6��r�
�F��pb_�)a�}a����7��x�OHx�r���މj��-O^��Z��C�X==�ط�q�и_�.M%�(-&����\��lLȂ��	���]�Z	`*3x�?�����Z�T���h��&:�쌾��"Ɔ��z2��2�r7��\��)�Na�/��l����I5�bV�3��Q\1^�@�hbUu��$�),�0�5LF���{1�(%-��/�2�CiI>  \��4�"u{	8��6���{�$rc�O���qz�����3Z3ŀ��5,s&��%;#�ŭ���ɩ�]�u1�2@H�~e ��2���������'�G��s\<M�S@�����_�"�9�$0�u#8�b�M���$nx�3}����p�Rk^9���o͸�}�.(�ޛ*�o�|j��i����eYB�)^E��jqUGicqu��_��vrM�]�>=�f�a�A��"��[��|�c���Q����c�{�J��S�q5z]x���N�/kةX��xe|�����dPӑ�'7�������i{ɇ�{�ϧkψs3#����,��5Hl����뀊aC8�z�3���H&+g
�7�<
���@pزx*t�a�I+�Fb�)��儰n'�z�ԯ��{�C}Ϥ^��1��C�";"� �t��@�t��c�Z_��;�����X�ӓb,ߌ����\�K�n#["��Cyڬ�ުu�W&�U�_��d�ީ��C�^���>%�	��{]�>�W����D;c��f��t�sjR�Gp�shi}}�i�C頋z��i��b��@�{�M��=