��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��b*]���I��̞m��w^o;�2qblFȔ����C�e�sU0X�81q��bE<�?Z-�h$K����w0J�(}�iz�C%x*�S�&�<x��Q�K2�oXKun:���o��ɶ� ���WÌ\�_`��~l��sh�֐�@��Q로�)�U!���w5�Vh�9���g$���/R��SB3�1��g�T��a�� � ~f��y����P"r�4��1+�������}���{Apv ��|�_О\N��N!�t���82�r��Ư���wB�揝�#�(�E�V�"�[}�'�~}���]ڮ0��jɀ�R�rf�o��HW!��]��&j����!��r�۔�� �������0�B��]���5n*2I�m���9�e9L@��Gv)�жr^L#�>T���=Q	�tQڤJ,H����t�p|�J���}[�O���ǶL���l�X��&�%�[9�k^��,zt=%ȫ������1E�����G�h�� �	�}���me\v �������K��\���raL���ʹ馈M>kx5vH�M:���U6��4�07;J�I��A�+#p7���J�8�(����e�0Q��^����]�Y��*�[Uw�N9�2)��ܫlJ/��pY�R	��p�.?���X����y�K+��WZ���;�ڛ!��X�6S�r~G�"�/�ӻ�ص-o.ffZ��d栟�8�y]��9���vY�t�]_\�&��+R���<D���B�X��jl0yk�5�@���Q�r������K�\�l��5v��@�I��7��K��w*\6=s}��C�t4z�Q6Ud��E=�=��7��p%���1�k��{l�?i閞X��qb�_��?�m�|�v�Я_�_h��@mS��c0τ�I�;b���dj�ͧ��-	��֚.���,)����%�$Z�퉒��C@���4I� ȃ�od������S>��AMő���]�Mej��X�P��8��)�&�-�,������7�ſ�@�{�X�ٷ�c��n�w��@�f�uҖr����-�R�����~��e���;�(U�Tce�+�ww��7�&��jQ�*�X�����Y�1[5��`�����&u/�E7��	�e:�\�M����UC��>�r�iV��bm(+�sgF�������g��-�r�̼�0:��`&����x����z���ĭrd�&m��M^GE���R�L�q�� ,��#�׌R�a�nF��AE�-��	$W��v-x�&�v��UR���՝�IB"���4�B��>�]��2��F��p�2+�`(���ѹ�k"���4�(y���n��U�|Ag� �a5�{s�~O0-wrR 2ynC�K~���=D7J��G�}��c���G�����+hY�P+.f�ZC��%�+&n'�a)�*��֟�2�"���ܩ�k��q܌�D0��R�n�u��M��&���y�=�f���y�'2A����yM�My'n7��h<pJ䋓�����{(�y<&��ݴr�u���,!�ɕ7���Q�_@@�{��iT���%+{m����5���.җ�.s���϶]74t�{�\=�wv�%O���{OB��v���%�mlH�s�&�j��x�$c'�j��^���M`}Q��%X��!���� a��EW�d>A[Y��g�8��)�VD�w����H����$:	J����>1<8LJd��=�e/)�d�ҫwxղ�H�+~��w��o
t��.�����[��o��k<����E\���_]��y����,ax�e���~�[l'�!`��e�zw����+#i%��48{@�^�u��nȸ8�gzBq`�n��Cx���+�q���0)D�&�A�!7�m�e6���r�z6$��#�q�3 V+�?2�6ώZZN�C��?c���N��G�wMX֔}�@��ď�r���g<θU�+��mQHa�c��ab��`�7I���>��P����;\m��n�3�3�k�7�@?F%�$��h�ۺ��9��h�R�H�p|Ћ̦�׈������2^�;XA D2N��1X��/�)`n|{E���v��Zv4h��6S�Β��
 g�&S�>P�@�d����^�+S�����r�
��J_�\�J��ݮ��ߎ�fs��%������
.�=?�`�@�P7g
6��`6t�(f8�{���U8w��v0����cg�>�z�q�_x.�w�(?8�9��<�a
�E�@����y HچqB>&��R&n5���p���s�3n�AD;���v�2�%(��ԉ� �|s�����4z���v��ʾ�ø
,ڵ��ΐ��X�B�&s�?_���k�L���������R(��t��\lj���t���e��$f6#��&b���͚4�x�~��3WUl=ʀ���cF�3@���b2��{�jk�߈&OD�Q_hŪ��P����#� �����u�C����Ofu#���^�5\�=Eɕ��pX�t��F�U��f���J�JԴ9�F/~?~�B*"��D�����c�BN�������������,6�90����(<��Fn& �o������(h�T���Ϫ֊EX8;ĥX�\�'��!�_�	��:����j�l$A�h1k��&�2c
���ч��Te[��d�#�
�R��i�ӛC�H_k6�Q���@��Ueo��G�@p���4��5iG�~��e����C��f�w��M��>�~�M�ӋL�ݶ�b�]4j��p���I;X�龌�Ԃ��$���g9�\\'*�km���93���Z)�$?k[�|Ì��"^�-/�?*�r$���HC8���/�7�"e$���P@��:�(7�HO#�`���	�t��*�s��4��I�o��H�K�dpe�߂=�$l�i��\�A$��dp b6>��^A������f�B�O^�C�"Qw~��O�@���s���w��Mm� ���ڗ��=f�����̌��sL���r<}���O�B����wF,���
}\_��(�Ai)��\5�JS��B80]9���,��*�@����D!_�]$9ם���$�o��H�}Iߥ�Bl�H��F��9���=p_ �։�͍B��#�m�]��޴4@���"�I�I5!y��lF+�ĐC[g.�p�0�
zY�MV7C-w
�A
x\�\�����&9��M���>��_��bap6���Y����^�7�J�%�˅� �b����r	����n�4��"$2}N�6��_u2�οz���j��v �׆���*���C��՗����I2��!M�^&-u���18f��nd8��K��Y�R�0���FFX�?!ֲ���x���rG�HX�m�H��
A�u�T��S�����8e��>���Np��勡��*��*D�sO1O��
{?��I���g�)={�n�7R;���x
{����'ݐ���MQ��(P4�s�W����u�#k��ن��pGŕf�6���\��zm�0	=�u�����X��v�X�X�)��j�Z��TL�Jq"" e��Y�B��Q����t=P�n��~X:�Rł.t�R��{�J(3i}�!�_�>#��L��c�ČW��&]���
=TG����0�J�tuS�p)�]�	���	^eVK��a�s67)u�!�E���Q�n��jc�c
le��x"A���RQqaLVU'����m���%°8E�n��"�)m�����`4PI-Hc����n9g�ʥ��a&.�lM$
+a�13Χ�>G�@^�د��<�B7�0N����6:��x	a��P�X�#���c4}�i@� �Ɔ|C�ܱV��Cv�BK��Qd����2)}�ow�j��q�#���iTo���{t���@ W�}��r6�r���?��t<�݉��ЈӦ.�u�)<�}A��`��zM�P:J��9A۠��Y ���;UT˺鲹O0����8�AL't��2	�����s
������+���.�:��<�� ^���Q��R�sRЕ��v@2��	�?�%A2K������K��\N��ps&\/	d]K`e�k�lj��C_�sɝW��O'�MO�&x��3"7U36����E#����KŇl����s���Y<K�yw1L�.V|̘��K��k8�Adm�zƃ�۴�m�A%U%5�4�S��R��e���_�����x��AB��		��*�,�u�iK�I�\KQ�iϰYi��B�'NvP��E�� p��� \��!���	�>"�;��>�x&<L9i������)���m7�µ�&�WMBGkr~δ��b��톁K9([�F�jĮ�m��Y^dO7�z�q@�謟����l\a�N�^�3F�%%���A��9I���:YAZ/K���������ͷ󺵽��eR������O�!����|�3&k~xe)|�������-��YϾ��|�d@,�N�M�)��>/7g�QC��oW��#��i���99� }���Հ�qϲ�f�>#�M��_�;[�5�$�9Km������o�Ӄ���F�"=sF��&����v;��
uTРCe������������i}ϧͦ� 1m쉘�4VI9��3Uy�J��[�)E	d�)(T�h4bL���a��l�ǫ���Ӝ�\}BŹyV�t�_�<N7 �p\�,,^�׵öBB�gYd��!tx��i�tͼdڤ����&>e�FL�@�����7�c����M�^gjv ���3��Ąb-��o4��D9{X���Ӂ yD�ی��J�ό��co@ͱ�NdG�"Ċt�' }[��W���
�~0h�0:�������J��zè��ޚK`�')�HDp`c�(E���>;�&o�#�7���,�5K/��Dp81����
{k_��7�)�fLս����~�2�*0|�:�$[F!�!�b8�N�G���;3�c�/����@Xʤ_9
Y���"Ww�!~jǌF-K�#:�c+�rj�)�CF�\��H�1��`?�/����jl#M�$��^�3Xg���/MT��y��|��o}6J�D�U���%toϏ�}�ꔐ®}���Oy��� }!C�=���x|�`(�n[׵KW�>��6�����/�,��mHG�:[���Y��W�o� _��WzX��K�<t�Jf������