��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�]���{��)���o��8"OON��Q?�@z�W1p�e~K�T��ojA<^�<r����=?�Z3=�������ҥ��'��l26�af��K�3���!K!�����i����>���	��m Ƨ>��!��Ą2]��m(���0![K�e��g�}�}����,é�mb���o=s���
�QT5&��s[?�N	˵m�p���A�H]�?��s�ߙ,=���
Ԡ��,���E�}��c�m�ln�D �6�U7\��${5��u��^�vve�(/��7�5+ryv�|=X)�������V��TW߰T)���,yC����c������}6�P��"�If�QG/g�|-�2��Lݲ3m��q$ॿKRd��n��0fv�c���=\Xc�I��^��Dr%�Π��j����b8��%=�p܃DL��w�ި�K�d����[��/R����)=�-�v��p���_�����*r�.�.������c�o��(���
w��������;�������.$xf!"ݠ�������d]�GX�[&�p9���!_���0���\V��Dn���Q�����*�w�ݍ�2)��J����+�L�B�PI�����B����V�^;Հ�:���`�3`O��&٠�m*��~�s=�Ĉ|{Bjz�7̙�4O��]#զ��r�a����i�9 �¿�)�
6	`̉kl:����_�D �$S�C��*�X�.-����uao�����^8����*�U7�mQ�>�}�z�P6�GB,5�kRг#b�F�7�ߡް���rY*>a���?k�gN��~��,��^@�l{N��nx_������ßg�K��h����K�L9c�`����1A�',�d������«��s؄��s�U�㜇�Uɶ8�H�-f��mkd	d�?!هM/�R31[��{�������P%����A�}RwSl�$��BïD��V�(@[�,�����&�"�ûz�,w*��!��&�f�O<�^m�֚�����6���t��9�Uj�|��i��Y8$m�4HĊD��\]?�����SBޡN�vG\3°Ͼt�O2g�r��)"�!m��z��B�{��zXM>;�ks��y�k{0������s��[��qu�� ��4q�MFػ�?��q��Ew�o� ��xz�A�?U�Ii橋���� T(��LL���/�\뉁�\3h���-@f2�求�+!P������D�8Z���0����.()���Su���z����Z�#�q��,�Y�e�K���$���`���;<p�>���t��O�	��H4��9�gd��z��+�S]�W�#�g)S�0~�x�W'�J=Y!�3cj�QR:�a�,��}��N;��'���s��)�$3�j�m�8M�ǹ���ƽ���`&}@�nZn �`��sV�\r�Ǳ<)�޼� I��5���r:9ja�;�D6ׁ�f8hQGt���uA3�n���h͵����vi�u�t6���|����sd��x���S��y����p�'N�����f�q5�
^�'���L�>rҔ}*���{��e��AJ�8�c��i|�BrQ,sZ�������~1�f]j����R~)z�Y�H�"���Κy�
�0��A�6C_��d2���/�@�Ab���c�nI�}g�~D�q��ţ׼����n�h�a�?��*�)����&�բ����)� ڏ�1�z��w��B�?`!�$��*�:����V�f]fj",��+�c���T�r�1C��:7<�4B�
������U�1+k��J-��S0>a�+J�j��_�Vt|r���\��?a�T��3�:q9k�1�t���_R���c��(�H�@��i7!�q�jź�Y5nS�ڐ��J��t�����$`����HF�D����0���P���lRE
H����;���v,�:D.LB&�.v*kb� ��$%�ZfN&��n���P,@8��tQo�q1m��ws"�۲ҏ�[�Uy��!�\V��g&&c ��G������̓��M�p[��o-1g���$���0qMQ�B�
����X�����޴{�,=��X'+E�����C�,��5\}��h������K�"9���"�&7uTՐ��m�NR+���p��B��qV�6y��1��q�@7~t��5D�\��'+�L���ݵ��[�A��H+K�o�v��}�D����b�}j��3��k�W t��2+�y�ථ�,t�$�b�dojr�v�E;k��A;�P i���w�<�{>N��5�ʯpd�苯�^�t��q�ۿ����g"r'x�o�d��������S��bIlFQK��N���x���r&֌�R��j���t_��DI��KsB�э ��㇗�[ �_h�� r��"a5��TE���Zm��d	��K��}*zS!LY.X6����*H���	��2�o�a}�bn��[��n������R���C��(��k��k��c��|m��N&�,���n�6A`Q�S�uk�]|�.��%�Ep>���ؙo,N&���;��5�G�g���N���q��=�H�D�x�J@�{\��ZF��h�F���)��d�UZ8Ѭ�Nh�Y]�R�l�H��B�U\<g�q�����QI�+�s�`��2A�h,������M�uYO� ��&�e���y�您�f�=����s���$�$A��� -SB����T��R:l[�U,�.kB�ؘk����:�v�О�d7�oJ�f-��VHS_�גV�l�M�j�ɱԕ��o��u'�x%��yip-�����>U������_��*6;b���t�Ȕ�Y��Jܙ�ifWA���]��|�:+��`�vc����.��T�Ƚ��Q�UB+�G�(��o�I�w������(��P2�7�mN�R��� ��eqv�����|Q\D�ݾT��>a�$��Ú��Qi���5")%�%��r!J=�7�ʵwZ�r&��mTk�U���'v�e���=�?�˫X�[\.���k�D�g�i6_� ���O�)OݗГ@�Y���:3��n���}��T<�pA)��2��
b �;ȹߢ��)�u��q��z�rV;�Ǖ���DfY���I�m:��G���X�.��?���Q���;�HOOMd�[-��R��5��0 ��?e1�4�9c��vɓRn�Q��Fʧ�.���]Mk\�y��c�Ĳ��|�pq�hU���7#�Ã�6�#xF�Z*�װ���Yb���x/,�*���sSSL�"�	��	�O��
��*>���v38!cB�8�����º^-�LƁ4�-�z"־kz��CD���~O��^TE��;�خȬ���2a���"��*��� ;�jF~�Ӓ�5�924��^�6��C(��o6$�h$���3"�Q�+�l�����8�̷W)sF�K�2ڍ��i���zƷ>,
�Æwl�yq�Ϥ�M�wM"U�H
��2�pa�>��@}�>�KoeEL�h��ZP|WH��dP؝fU�҇�\M3r���~C:�����0[
�l0�l�/���Xi�s\d��׫�ћ�	�.�}y��<��2(�<T ������-���.���ҳTz`���E�[�Z��JƖ9Nƞ'Э���Jƾr��^0�ʍH���]rܔQ����Oy�9^)��;"��4WO>=5��s}��f�mN!�c�s���B�	��޼V�50P���,��[���S��?��r�)�lF����Jty=*G��a�4��x��g;�t� �K?���Or-�9�ͦ�O�V��x���C���p9�#�́�8�l��yj>PKT4>�V*+���=/U]�>�T�5X���0��-���DDA~��:+��Gv�qah!��p��S߅�gۉ�f��< ��R��	���1)~=o"Y�O�
}��p����|̠�E{�lmɖ�U-,.�gQ���W��ƚ�E�� �Ġ�z�U�~�5'�"Z��ؑ�9�R�E��g�y��1���*L�7ҹ�﨔0xf�V�R֒??�?��s؍�n8b��h��8����H��{l�t6)xB�A0��<K����}�wF(|��V&ag܋����hu��a� ��P��۔�*���Z���4,�C��(���.��C���\���?	Ȁ��q�#���6l�j��\�P1�N��f��O�mR��0s'ؑS�Љ�(�.K��0@/H]h�@J�3\�g�Oͳ�u÷�v"B�D���p .}L�v�r�m�ˬ~�83X�[��$�7IL�rw�vU�{���g3 `-�`�}�V2|�X�ɇ!����9��{������St&"B�jpO<-�:�87b^�dH��S"����/\JzC
k�?Ț���Z`(,rMc�3y�mYmƇbܝ��c�`�A�q�I�E�^����@�ϯ�;�wJ���z�}��	�m��NE���BQk�(�3�H���\���է�Kt�A������>_,���Ar12��.��R��`�؋F_�Ȥn�*b��̅&bD"�ڨ�a<`�hD�e=k��8�V1t�����V��P���>����U?��i��6���X����`�wRy��~싯�E��u���+���93Ж��Hӡ���K��s���L����d����QW;����	�����g;���G(�����\ņq��� (��Rn�ٞ��J����	Zom�S��S��7D�)E�=�/T��_�r��Q��&ᩬ'���T˰��1���lk�����ǫ���0J��G輭�M����;,�71�(��l��j�Ҿ�P@@��G=C�ǻ����Sրh�QU�)� �xA{�]C� ���ki�b&O��B9Ӑ�Q5���%�B�K�dJ�]�L�� �ȳG��E�U懙\��[��
�kTj�yx�@���q��jB�"͍}�P@U��O|-�EJ�$�<��dשp��.u'�i�w��#!M��jX]� �C]���$("�g�Eƾ�U�{=�>��h�t�_�i,u$;!D��;5o6M�߸��-~�D�J�G�=���xe�ך~��v;gSG_ϩ����B��Y�|Z�{�k�JI��R�ixw�Ӝ�ڞ
��|�ng^l������?���$���u��o>n��nheV��)�^��>��&ځ��nN� �(���w7(GRJ�1��b��$�X�&�A+�A°��'��>�v �����+�S5�AD�����v�Ý�y�#��I䥐>S&��z�K&�e�-�b� ��ME�q> �<(�B@�W��gQ�,u���IL�]�10j��UA	�#6S:0M��!�\�R&~�2��Q�Ξ*{a�S���Z�cL�dّ͆W�Alɝ���߾`���=n���5&�-{2ӌmUNY)�曮Z��ʖ�����5�0�cv^.���j}��u�vB)�V���GNӿ�V�@�]��� ��E1�]��2;*�S)r�<,������Ȁ�}�
�P�d�&�`�*���	���J�;
*jA�k �^��2��X�rX�\lA�zǿ��f�n"���-�&�������V���\C~�I�g�~�8���K���h`bF������J�z��5���Ճ���%���_��'$����2�Ou��є5�IQ-dˬk�b2��PL��;O�7&ʶ��Dw���]J�`C��mL��wc-�.4��`_���g����fH���߆$�/����9��.�<��^������0	<]��7�wD���e4;�=M9�Q�N����
��]4������� �#��~�ID�d⽡n0����H�_ײ�ׄ����"�/�M�vN�ӓ���!
���?��uй�i�/}�W3�<�"����&)kP�H��r���u���\v)�i�Ϙ��������l��&�	d#�sg�b��w	Q�%�q'z�ݿ��|�_ �gߜ�</���OmZ���tu� �h�BK�q�N^I��Xg�"��ot<��`����﬈���5�*o �NKz����g��َ��ݍ�30A׬�����:���Gh��c���<ϼI�MÝ��&X��$&ꭩd�d��{�wv7M�q�G����n���U|﯌M;���3��-��rt1��0�S� u�3�[�� ��fPh�VP_�	�g�$�;�H�	���#�p_j�0'ũ�n��U��cq@���1�Z{��t �~��^�������4��$<�5B��!�1 I��ٖ��]��'N�5�$���!}ɭw%)%֒�^�2�
O�l5���XY���e�o���3�G.@���(c1��ǹ��5�X�(�_N{�@�V3�xT�U���"�@�rv�~�o�����p0�0T5�N�.�"U@�]���p~A'ů���y>bwsHT�d�)�S ݟs�щGU�Q�{Yf��8��8����շ�8x�D~�1p��l�=EM��.ns����/o�h��hJ�r�U3�o�����r�5�"<kv��4!��x�Δ@����ɪ� �7��w�..���w6��B�p�V�'������E��=�|��㈃r\C�3np�Qs��㶶���=8oh��F�}V5Z���3�6�F�L'��7ux�cme�`c.���g�5���^}�[,i�on��Ǵdh�u/�b��1�"=�V��L0����1��G����(�/���������O�"4�����):�`Z{��[�T��4x�P��NR�<_��ou%&��ls��1`�T�Ǻ����~J'�t/���G��_P]���K�&������Uz9Ơ+��2n`�'��Ym@�St�mV��&�,SK��E�����?G8��#(J����v�cGy�sǉ�?B�5,qS�%�-%&uN�ʴS�3 �Uن]9
g���L>C�����M���#�	��=y	K鰯�~��?�#0�2�n׬i���.�F�H���wٮ5�q�q�k"[�j]��F�<$�mZ�1Y��!O�{�,'�XI�ÖFmg���J��c0&)��p`V� ��	����<k�Ua�`��O�� YOQ��\��+���W�-(o
��p�s�a��i43+�?�eJP��$��b�Y����k�U2t�����~�@���t��3�� U����s�mN�Oe^��ͳ9'�o���r�ᬌ1�{7� �s��*۔E��M.�C]T�*�^ܑ�9�Լb'�yyx��x��v"�W>@�H�Գ�Î��k»l�0t�U�i�=�P��Mh15�wMGsR��ͤ&B��廠��|�)�Y�jh�,1���v�=Z4�ڏ�c�1-ӆ0��+� �E~��{�kv�1c:��oV�3�� F~�+���g��X�����"/�Ư�dY&��M+��	(+5�NuWo;�,�����׃$k�@�����g�Dd�Z�l"���>��}/���F?Ï�ws�a��?�� ��n9	�D�8�5�p}b����ZpU�7��e�"}05�pC����{�z�(`]2��$�ίw���Qw�8��/����t���y�p/b�KKɟ@����F/f\����o�$sô��+���A/��Ճ�c_���o��П?L�8�D�6�h�,��Bߜ!)�7cn9>7ka����7<cs{��ⴰ"�hZ���6j?l;4I���}��s��[��ER��P�+k���������6���yxh�&�	�?(g:t��9 �&�$�=���(fy���Qi�H��z�F�aX�,R|����������HZUֺ����G�>z��
��5�Vt�~��=�.L�l1�Q���V���.%j�����>��j?�M�a�T��r$����JX�G����C^�.��͟&�,���o!�O ��%� �B �\�e��;,T�SRuqcRK��C���	xW9�vn����f[3G=�[�em���J���5
��h8�ψ����h�xeO3�M�,�ȫf|����{�����W
D�6�r��"-�
Y"(6C����)�H�o�x���w�j��8�&T�+�~}_Ō�U��H��9|��5��V������]2��������c��RY�O���T�V��su��K�X{ld�3Q����N���MH㡱5 �5�O�f��	9��3����d��\5d+;�{-9:Ab��H��!S���R�Q\��@�	n�n:��[�ܞ Y.��v�m�����I�)BQM�,AMu�W^�5�ؑ1H�*C��S���2Çq��}f��#�L��o��5���&?=w��ssuX*�ؕ��S�j�����B��
,J�.'�Dx�:3�ʭ�m�$�l���^����ߕ�c̊�7��9�t��e�'b�!	V$���ƃ����d�X�_����Gr�{�U���1n���d��q���a؍�u�8\�M��j�~{|�	Cv�X��O[\�uz�ᛇ Z�ْ⦁�m���q٤�W�-���Z��������"�0^VZ��N��C*�q�����;���~�O��}�EM�OP)xy�S"��<8	j>������p`����ϰg`[�R9 �"r�+̿K�2������4-o=e�^�$$����S/@��B�g{["�´?C@A�!i��H2��c�,�iP���y��Ԑͫg���%u�/�������R��w�u\�±#��Q7��{Qs�4�� �1�HL!�H^�ː{\��o��SH�^8�F�s�d�~0����=�zÏ�5�,5�|z<��l��l���X��1C�?aZSu�Qv�~L�$$���v�Ai�N��[�W;�s�"j��'�s��fGB�okT��$R��Ԝ�??=F�	�:�^+�g��l�n�j�&ҿ��%��-��H9l�	L�Wgn_�"�Z���Q��E"�BۭN'슠�na!x��Kp��a})�	-o��ꆩ|Ċ����;��Ȟ<~1qb�h#��ǬX�ޙyKn�ϲndb� ��9g�n�/�u�Q��!Ù�j��CC�����P3ێ"H.��0���@iF6����e��Ӥ����M���X��=�gxƺ�θR�F~-b�B���1h>��m��h:Q�����m"
z2(w 2�
k�L?1�0��\hKp2�ꢙ���
{co��V��ԃ,��n��}�[W�Z[�&�P��M����<�J�um�eQ�g�M2�*պر��-�JU��߱��kj��`���,�ԢO��h�
3�0�͹;f�5�e�O�����:���5�}ӯ!���blj��X�fr0����F�ݪX�c�W4F��Rm Xvw��d=��ks��|��!>O��q��2v��ܧ�`�8�}��E0�Rq,�)�Vq��u���DB����S8?36)I�0-u{:8�c��\�$�lo��1,P1dki���1P��)���x�<�⻌�˔��~m�RM$�eBwP,��:}�s]�$�=���7s�U�m:��8G�ԕ� �^C�:���`ڛs�u�r�"�?��s:� �c�"(�zV�M'�3��]����������3*lqe2��yw��=��MXS��5L�X������7Q�Y�1��m��R���f�W9���fbh�`^�Ep���w12��L�H5m��w���gsRjɵ�����]�Xv�R�kN^du����w��GV߬�E�hC<t�f<�^����H�d�}�l��z����S���o���4��QtRY
a�;����FE+�U�c?n82/c��Nd�mw�kɿ��2�AC�}���QgK?��� �Ԉ=�IN�K�-����Ǹ���(��D����(���m�P1A*w�|5j�1�By��t%��P�8�CT�8+D���P�:�����Ipq����1���$�9&��D�%��.Ӌ�C�c�`exЏ���]�U�x&y�s��f��_<�'�\��#"�wzBc5i�,9\t�.�Ws�����e�p�d� ��\��G��y�|�� �>h�9E��t�v?���T}^��*�����^�����R���9�JkJ,��G����Z��ץ��|��'��ii�b�g_��;�d�7o�[�ʿ��x�c�m�ym� �����[�o�����}��*2w�� ���x� O��'�,�6���W}�%4�7�p�
�M1�{R�G�K>�0�z0'�󤱷��o	]�~n��  5���>��.���X���>�\�L�4P��P*f��H9��-d��� ,r�V�){���50_��):����0R��1����6W���z�3�wSF���K:���rA|��b����B?	2�;�#�شg���ʥ�����z����h������S�����9�t��~�o�Ó}1�1R���H9f9����>U�M�yS�~�D{?�r�I>)[��cz��.L���W��|���Cċ��r��!TK�	u^�l ;����
)���>���b9����2'���Ɨ ��[�+�28�D����~D=�2�p�$	ɗlq����6+���xU��d��	x����3W�?t�zY���N�D��|޴��0��$?!$�i�ڌ,\���*P4�2f\<ޤ�\�iI.W_o�g�����9�w��^��w�tƇ,i���k�l�e2f�`!��2oD���0H0����0��v����xd?��l
ak �7'1
��sQ.	M)�5�GduR���?k���6%�{<rt�8RB�'����f�
tg����w��@��^�mFd�0��c�}�W'<Pb�6L�3��6����]��=v�W�p ?'Y�	�k�gR����,ச���V��?��6������)0��J�e���^?����>`����[��+�}M��^Ɇ��2��7��y{8l`����*�5H�L��K[�[�S� ���I��w����\���l�ި�5�N���͑$٢ʹ������uj��KN�����N/X��,��w��ڳ�y���wo���4s�MV�7�)W�:�j��B��pY1�g	���

����#%.�4� !(��Za�RD���Q|J�j���!�z[s���(�O��s�1v��̆yc�~�;��d����6X���N���1Zo%�.���5噥�i��ޏ�ee�?!��s₷��6*5M�_שջ�R���,P�E_����(7ȃ��@4�3�b��3h1�Z{���j��a�V��2´���;}|N�Kט��gF����+���p��#����5���R�K|���eu��+G��+�����1E*��e�����"pz��$6���S�u���7=Fs�$9V���#�aP�ǫf�`TU��r�Uty	���_)�C�M{�� ՟�^\�[b�Uc1
ҁ�
P��&�V)�o��N�!
�y!W#�XwȓV"P�
kx�1�%�ޤаA0m�/�P�9��8�]!�� ^��2j'��hl�=��̶SQyt�}�qc�J�ŝ��/�~�;_f�A���f��xd��0�~dL`��$5��	Qh��W�H:���g-)�hbW�>U��?��hG�f��C"V���}I�h�b�$����'F;(TD��8��$��������K=\HĹL�D�����d\S7b�T��W��l����l���-����y��}�m�/�f_�����*�W��	K�̊����.p�]�	�7����ԕ�%�2�r^ح�%�%%�{�M� �K�7ޯ�¶�|�&�����z���Բ���,SM�1�8�{|{�������;smc��8.��,���e��=B�ޡ/2����y?,��&YN�ל=���*W{Z�?�F0�=�5Ԡ"'(�ʾ����r
�i˘Fg��ԎG�
�
�dzm�05ˁ�Uc�|���*�)0�[��7!��b@�7HI�CQ69^�7T� ��:���{D��CX��O����:�3A������L$�{[D,��u���=w��*�v�W����r� ���4��ԛ�!�ٗ>8�<:��'�E�W=;�5A���2+�u;2���������ݹ����C�\zq�]��td|?u�F�����m�I�2�+=Y�6�� �Ǭ�+��!2i	�Y�F��>���kǑ��T���$�]qL�Wu�D���+�~Ptc��AI��9V�B��佧�.�^_�x#����d�����C��������B�ǰ7��W���1�1p��@l���{���-�0�n7 E�T*���ýt���n8z�lQ[�8B�u��U���Z$5<K/(�7n0�x*���ۻLf̤�(�C���50��lֿC�&�6ˎ�],�{T�1/�?5eD�<՚wۀ,-�݌���+u��GiFi�l#X ����`Z&\y)�"���U�ت}[�Ŵvժ�c�R�&x�ϑ�7Yv0W�e�N�,"|��s�_�s��#����!*/4�:��Wp�:��*��R�˯:��h&|˧��7��V�w`|�����5G�����o1��3&;`�f�=��~�JkOO0�w�+�p8�9r���\�8\^k��/ݓ�rF�Mp9pQ)O�}�!���6�6{^_�[��������K��q��?+�ahur�̲~PYG�BvN���FC͟��Y��sɮ��Ի^��V�{)���ż"3]Qi� �_,�[)�t�,ktVFܢ�@LK�`����CӨBt��NX�;%�):�rF\�����i�0�H�è�U�&�eJ�j�?��� ��j��(*M��Oq�)`$�
���m��Ǚv�n����(!{�v�O8�5����a#���ݢ����zn�"�UFlm��[�F<h�]�����6V&s:�{��o�£��G�Y�(}�#MVʿ�d��[�I;Z�*J��7���c����a��0g�M�9�^}$��!� w���Ǉe��Ҟ������|v��R4'��"P$zJ�91�F$f��T���'� �?q��x�a*kH����6��f�_��,��P����i[���tl)n7���E��1�J�|���u���4��w)n����G>k{-l�P���r��ڹ��P���V)>�``���[�d�m��bv�<dk�L,�Ɉ)�
��r�y�Bߧ�/�X�OX�,j�Ϝwe�Q<��y��Dh����