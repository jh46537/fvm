��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�`��L�o��<�T��u_T2�MA��Rɸ��~�u�Қ��r���=���]� �� ���H�+�LQB���=��V��پu�~!5�Im��`bw�U�㛬�\���_�R��Ԟ�&��p��qm���K���������H,e9��]�vCj�l��2�V�n��˺1Y�	f��׬��D�ڙԱ�Z>�-�����/�Zw�g1���U�ZCK���b���ud;Q,�8H��Gk�����{#��`k�/"�0խK��Щ��'F��s�Q�ٍ5D16Db�(���Ue�;"k��Y5�%�5�N�]]��Ugx`��׳[�(�,9H��ʭ��3:Z��b�+$ϧ~ԨI���#t���H�|OUh�<�3,�^�ɛ'?ܯ�6<����p�b�M^�� J��pr}�=F�\��(:�z�w=��?�2@,~���\�&PC��AW4���,z#d���N���C�_"`���\:��թv����̉�T7u)�)�H	���00~������������^k�F�ǩ��\�%vt���Ϫ��q,Y��\/�n��n�������ME���W�d{���H�!�
>��Uω��D�n�#�z�'�R��{+� V���@��f�$�R�̌�Vqu@�����ҭ��#��|ߜ������2���2*�r�_J�ܝ�OMM<S��|$S�Jh�{Xl�m�}k��6��z�n#�P`��n�K ԕ� �xD+�hY�*��ܓ��������r�uB��'\�tCH��ۡQӣn��?$|���
r��`Y�0f��%�!B$�Q��2b�� ���ۆsL
w����PV�{ZV�Ԣ�q�n3��?�l#��S����
���N�3�±{H�Â���������@3ƾ�����z��xH��lgn1����1�6��i-�E������㠃�[*�F��_$i�g&�@�{/���,m�J���FLkk'b�Ѵ�G���P`��zP�Q|!�w��>A�j���O�P�Fk!߳�X�۸���R_�,F=b��u�{9a����}�K�5L8�<����3��Z���,��a�_RaTP( E	}S&��2�F�B�!�5FZfQ�0�O��?���7��ܹ1����MB����.j����g�o`��N�7��q��y$��&�)xGb�嬽#�0"^�Y8�h� �*BQ�V�m�c�?ϣ걖c%�$k�	T{��"�1�8~L
�Y�D��D�������e�M>9������<��da�uT���v��:j)-�]U�>=@h��['���2�7�p2J������QD�U$��I��h�#k8]U��`�+_��} 2x�� @��W,VЃkT3��ܣ��Z���=������n�6�M��ʋQ��I�z�q�� �A]�rz��p)E�1���o�9��P��H=�K�KF��/.�Y��-��7�4�\��O�߇���yĀ���+�H�!q*z6�7����US�b�@
���,����j\�p"DC!$���\��쫡������QsA�����Ñ��ZK�P!5T�q9L�0�, &�b�R��5�Ѝ�i�=E��aeA�}�ml¸���%ι>pkyq�Dg��"R�l��i�~?������(�F	�ɨ�	mFr䱵��#����kR5!e���qM���"A2���9_����.�&Po���cL����:��!��Z��E}�X`��l���^��0BQ$Xq��]~��%x)j0-�\5�^�K"��zk	L�,��Np��U���I�~o��B
i�?�B�Q��+O?Cm���ڬB�+܍�C�<�n�Ғ�|� B�����<�Y���.�ا�kCv|6�'F+�-/�!Ů��y�t�g���Z�_5+�Ĳ�1-N�7��C�dTax����\�+	�Y���2hF�l`W;R�H�%%��.��h/C��$X��t��ЌL<ߊ�u�U�����:+�
�DW.�+ �])CV��"����P���%�Y8(��8��"�Nz��Q�[��z<:��X�8���)I���B�޶�l�=�Oj�BOߎ����x�:N�!��k*����$&LȎ�\]�2<��~�,^뀱��e�mZ��[�Lxc�|k�)�^(�2���L�i?QG��$H���� �AP]�y�-AT�]$����3�)���9<�wh��|��Wv;[��Fv���O\m��Vu�}�ʜq�T����"���z2�؈��9�)�)�Z_k��f��c��x�HXa�|o�J14:h�^x�%])��A�aM�A.L�QF*� �}n��(�:��unOŘ�mV�D��e>��(����JߙK�/PM�A�c����6�LY�Y��[����Z�+��C^��#Ji��{�9&h�*��Sw��GYRO�N�8KQ�4[)�W�ZV+�r�9�[94���Ê2̮!�,�_BƑ�����u�h��-n�Vn�5*��4�Rи3M4����a^d)cWajXz�A,3G[��,��L;��F��q��j^x MB���Q�b޵R�]ۜX[�X���A�]�v��eD����ZQ=g*|=��=�'�[��2bY���bd)��N���୕����PB���������Y;e�x�˴�5����V��l�ޚS�umFH�Q�+�a9�`1�J�Ye�!X���%G��uv �����l��?G�M�������:Ę��
})����aCn ��!T�Mca�9��'�yQ��3�1�0�?\��c��v�QMe�+�����v�Nd�l)[��a\���W�v1���X�"���1c%ڀ�)�s��4	���S$�=�?/����ؗm���$�X.���n��]��DD���`txO�wXv�k�I�[~L��	qCR=/��-�s>���0�}	�V �����&�����k3��F��񫨧UΘ�C�Z,򕲀p�tI�&P�,@A7| V����D�A����l�7�x����Ԃg�:����Ĺ/i�|���<�UJ��e8f:���Jb�H&�������r6�=�T�n��y..��ә�/5��݉P[�߂L��㚽QGc��U��w�V����.?�Tl�_#-�j�I��8���^'��?�������Զh���ߝ�N�Dt(޻�)��7@1�p{�+ڡFţ$��d%�f�@͵_-�
�F%ѫeH�@�P�W�.�+%��jPzx���,f����*!{ҫ�܌�U\�*@�|Q��z53F����S�ڝ�.ۧ@аW��&��`Z�v�"�G�1V`�= ���C��L��5GX#>�M�D8�kk��F<�g:v�:ƣp�ц��In���7���a[�g��$x��}Kr�y�h��X��J��-��)�,�3�eFRK��y+~������e)�6NI2�����-*��WY�u�����Z�&�^�M��nU�<W��_H±8�Ik�[_W����&4�}��}�M�C �7���Ү'����kt�Ap�����tP�:�>_�@c=�S@�����:�4�ޘ:�,^[�t�X�--�i�σ�'�TI(ε��"&@�YP�`�D��`TJ����=PX@��c�ö~'�b#F>�u I�E4�)oy	���D]c0��9�
���8�c�686vu5��D�f��^ҋ�-�L�bl���#y1�DfH��ַ	����'
1��rﳋ����T�<�\a�R��%���ǲ$u�5I=�6�HǄM4t�P66!#
�Snh�������b߱U��BNlY�h%o������m��c�~��zw6�q�'	R@�����LĘ��:�
	B�[��j�@��xu��8 �&�j5�' $�p�� 7�H�;1O�/\���蹍������ B��C��w��eW��� (
�F@���Qk��B�A�N�b](��n��J��������'(\�4��g�(m܍��	�*��7�jJg)
���������`��XHz1���f�~�#3��cl�׾ݣej��������6�y1�JTJ�>��"��(��훈�Rw�����a�t����'d
H�&_x8�i\�+N�Lr��g{��F��dbuY�'�2�g��b��Z����%�Ս��p�S�7�i�J�fW3���N�i���K��O~KXʶ0�X$�\Ba�̶k��M�9q�p{�>�.�"�ȅ���Av-�M�r92M�qt/���Dg����'�7�xY�烦/�#U{�9dK2Ap��,��&N�*�
�,@�Ԝ8c�k�B������=E61|�S�d5�Ԡ��)~���
h�~�T�g�=D���g3��q�[���SsC+�˝����b��	=����D�^��C^���QK��$&	p�¼��3���d*��s�V��}�����8Ɓ��[�d?����۷:ܖ�Z{���B��)�%dq:y�i=X�:V��ų�Hj���*U�ckc�wQ��%xv��g>x��M���'�汁w��c��J��l�[N��k�ҧ륂���ے̅�>]!#Jᴾp�:E���Ϸ�?�0��+�z�.k/�;u�vp��̈́h�ZPWXh�����'?H��{/��ҍd��0����z5��y��9�&�l��E/Lw��V@� ��bX�ø��sC�l�U�/s�j6v��z�N�%F�����P9�]�Pܳv���Q̜پޥہf��g[�^�Z���\�'��X����5�tE��^.i�R�ęB�UL1�0ꆩ��� �-�E��R�ÜO}�����r2H�R?�j����q��DI�a8?5��F�Ơt�D��D�~J��iU��RK��������=!�8�h� 0$�����r3����>���m!���ӆƾ�#���,,�3�ɖz��| �j�n�od�U!O;7����@7���r���Q�˳����-�S~��$\���;��<j���X�Ɔ*��x"O��tg�Hܖ�D����c?!��^�pl*�.`1	��^��/u�l��?�:�}׺iPl��'��A����<�w����"@0���-�l���}����Pj��������� �M8�cITCh��q��w;�V$�z8�DvO�<[@I2��2�;z��C��1K���̬�~�c�,��