��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�=WM�Q؅T޺HݱCV.�!ͭbs�.�8�y�U't���V��ăb��%F�#4*�O�ЈSxK4���mlZH��C�>��\���u2�c��́<q�~	�(�$�����G���F�O����6wU<�,�-��O*��G���	Z�/�쮣b^"*T����'|��c'�%���\�֧ʈ��O�_bl6�_c�!����V�e \Iϫ�=�d��h�#�)�(�cA�7��yq���R�^��o��m�/��9_�u��yՍ;1�%1?�Y�IP��3��^�\V��W�,��37Hc��L��T/sq���J�'� �1�x�;�hP����e��7=�]-�l+wĽ�־ؙ�[e�̊�V��L,�,�3�;��w�c�Eg
�C}���`��P�]�bZ�Tk:bco��ڙ�K��"T�@������9���'V5=��V3T�&|]�m��)=F����ye�PʹpK-�ej]�䅼��A��ڒ%Ʒ�@6B��!H/'�6i�
�m�aSς���QwQ\@���a�%ӌ�>��
=1^+��-eLP�V��花�ڣt���&�k� a�r�l����{�ܓ]v����Z�uv��由��&mlZ�G������r���OFjt��1 ts^s
Z0�!��=2������;��;�]o�!�Xry�x��]zc�=�<��'��&�rE�����٧Xz��^��5f�>Z�f���o�����7S�r���Lv(6�k�VPWTjD���,	��~�7�9"�d�4�ƪ�C�O�սAX�s^KoB���.����� Vg�W:����8���6���W����ٞ!G�m�,�"#������m�|�ڀo��2���O���{���\��I˒o� 4Za�o�5}˫$�r{�!.������^w�x�O1�/�t����W�g,�iF�畟�޾#~yG��n�8;�jB����ʔVpvq�WC��gD^��2�a����O�~X�w�ߔ�h�X�z6G���;V���qg����\w�+�H�$�R?�^%��/� H&󝯪G �xkD�k}��zD����~,��{Gs��7���q�F�+hCL�$��#�z����ꃠ{��s�U�o�/�"H��6/5kCd��<W���
w}ݝ]��`e�RO�92v	ϼ�	e�*ַ�.�*ĺ��<�wu���"��pw���(�Q�
`�ۢ��l�~+������m���]	�J[|]�u5��)����}������Q[>��)��XϬ�w��� A׌�y�1���ŝ<?'w[�}�>�!���i�PV�5�t����
^���5����P��L�5<2A�:
xl����
��5İ�W�BR��5wm�������w��iUI�wp *�S��4�u�7���W���`#oT& 9�?��4_'Q��; G���Y�*�\��fd�ʏ����)���4p��[L/��]���%`�6��������Ks| y@ ���Ѣ��l�|���<�����m���(%�{����C/��iR���}Ң��h6�����{�:�DDr�_�֫�\����54?�k�"=�C��شO��G�=Xm�!s��4 �d)s� ����fqM�c�r�}\x�ՙr�V@�J|����Z>��a��Մ�K��7��U]��%V��6��?��aUZ��\?&�#s�r�DL�sQ���>W�Ջ�]m����W=ao����g�����i�#W/��ϡ땢�J���!��׀��8�;�Z�H��G����`���2�����q�����P�+��c�#&�2)�V�ި�COllk?�� �\h;�v��.Z6� �Rg;Pz�;�l�s+� ��=U�7�t��?��7ɨ���Y�T<��$�YJd����Τa����H�+�O����0[~#&@�
dW����o5v�Џ���gb��A���_L�U�O��a~6$�Nq��N�}B��}H��>=�}�C�G���@��*� & �'�_�#��0Vș� ����J�`/���6g�����E)�S��o�ۉ?p�S/�7"p�P��^�/s ���K�k|+�8L׈��@�=�5���mwԉ�kQp[�S�=�`��E^�(]h�