// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:43:32 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
O6Qnq+TvUJ5RZaPb8cmSXnLXrInM0l/huTI5V3bByENkgzXqgaVG3Gw64z/WprKf
wTz3Q5YOmdBrUyVobG/yOb0SqktL7QxQirRNOMvmWVTi0ED1C4xKV5e0dy6ZypTu
Zfai5eEA9u1DdfvmHZ45mik0dmNBpfJO/8lAry+vPus=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4336)
7BOQv2L6dplaoQmx13n2h8IPmzqC6Z3jbVsMPjXHJY0fmbhyxN7ByrK+cEo6Upkx
xcz2uDLgaeWgglA5kv88G666BCRUVWOLL7y6O+uHZucWsrBT1PFRdNvglWcCCimw
yR3jSqOoyMeyQUKoVde0cE2c/du63ftre9JC7Yp0/HOS+TUPbzzgQ5M39Fbd0Kqw
H20O2eqoSRwANFdI5iTH+akv2yVKzEFSHjmv+WB7k4VEpxCIPcpSSWhD61phh5GI
jt5B66+/8Ys1SzIsb3GQymSozAJ5OVxUfKUau4Um+pvNxntCvIPsngkWC/mHJuNa
gwTDW5aznLVkfkq6NMDAhX0g3SY5Ca/ALKXkbzRHjDBf6/+2CsrybyOYN0wKWFZg
rsJrhUiOXQXosH7T+scHoO8Bc30sJ2n52oG5IfKb5yV4ieom6YKiB3+tqF3PM3Bc
BxJiaF7eNijH16GQWVIN57HBnwfzicxGwtpBzmFDM+1e1UGRyairxDCHCdOxkOGP
rRF3kSqD4x5KjPiyWbLRaLNqg7vZN+RnoE64lYNtEo6cqL/tQ0HvRuapTbBZckH5
pMSlmRfbqJ4dl90RVz2RqQUlluo9jj2m9QoV50kYkgaGYsjD5LOi1IAhmUaM3yPU
19ZyFNVxBd2kPrw73pMC9C++ZkdZOBPPwe3d6auLaOO6YzGYAB/D3LGlORYJSu//
bL8he9BaQJKxjF5cA2gAlz8qu0NciBtp9OK5tmy38ySWg8zcKqmzs5i629SxRhyF
KNzmw929dIOkEJ6tSHZwL/J8uMuDRhi0/NCFPn7alc3uN8Q4WfUxbzYJMD5Au5v7
r+gxflV2W3Br+MCwVof5IBJv+XgOs9AzqulPp/M9uhWliWRNvwXnHvbjPPLdDCtO
iCmGhbyv0q8oarkmMM4hN5I5hqgyIikq1rcM8moIUqn9S7Fud5JU/UoSvxKYIFQH
fyKgm1juC9jbjvAiy8d+IRzo5jSQsRhE7K+a1FFFXpfnuYeXeLMpVUjW5xLg7bkI
++TARlEjHz9lFcwZYbXdJbQq3TZSBzSaq5OVIelW+zA5GpM7DyMbkJpMf8YjztHv
HSMoPIzYkElIK7ruNdfofsdqI5nJ2rBHzuNrShvb4xPvI8bwPqqmDOrNZBuGBD03
SJ1bCt4H8lsAX5c0EaFAQ/BID7RA+6STrR6yob4RFNIawN0AKCxduwBctS2yr31/
4D1Ch9H8w3Vk/XjGx/zXXlVBrSSISUN6dXfsbBYQWgurrNpycsOSzn/S5dd9PSfm
ewMpW594EoK769lgrSMfNMaNUDDIqpguLDZMBgrknvBwjvFwfzEGCThV9MqeW3oI
rla5XkbQfUkYYDoSjRJ7Q+7/+fMqZhrchTrPWGjZnQ6me+fRrpb1s6x+mgwJfkhY
wv4+R0a/PcY/nlfsc7kRFRDm+G5GUbaTkwuFMzlJwu95mDWMm+KqL8vHzxqtxSUR
rnOek9KLbVOCthK5QlYvPOR7H01+afUM+snrFLFenWY6CJOu73mUZasDNvHywi27
cFkPRUcUXL++rLeekDeeX/qLOn+AdIvovnfL1xqDKR5LxYA/I61GKscIWnfILfud
+lIsob+QpeOc67v45L8Xr+T+InVUMvuhbdX7ZHr/OEt0VW5PNllfgXFyRhWStUra
F4zSISg2eqrWmKRrfv1P4091gccaPLHHYv6pPtWq1eF8Kw8b7oNENmm+j0mZDUA6
S37ERHLeEV3cZo60hl/WLkjF4OmYDpiNDrX4AgT1LQyfTRgBpRMIPv4mp5XpL7m8
1ft6AFm8U7VIK0XK8NvGpc+k8WQAiH0KZy639GYTpDNybJ/wLHDD9WRWeAFhWYZ+
uz6eM43qzryWYB3f4Z7bsqbMYi87XJk3w4nafJeescFqCx+MBqWHTzM50dv1bc8s
gfzPvXpHdqVjQ//OkQvazgsWzCqj4xjXKbnKM6eMSNbvmcKdA06+FEvdmOHLkcxC
yAbJfsUFCfUBVCFZXfAg8FMtTN/SpN0ymrMhdXJAaVz8veFHkFrTTOz/I9SNnaLW
SnWiXmnH2Asn1nVwM/XaKFbKC3+cBHFh/atLfDx8EgtUGE4xRi40zm2HKqMfI51q
++uG4ENCEAskIgpO3Wc5h4wQPy6N/yH8YuSk1nIPb3BnL43r59fjws8oNEOZGbZn
MpbTEjw2ecOuuwszaWy3bQwdyzPGTp7TEx7ECc5/HukQCpAW4VsnjoHOMZuw9TVQ
VG5/yNWtgKVy7pBbrJX550tRYILMk6GCDaBIzS0/yJjFYaUmvo0/RIDCG8+ClBfj
93KlmV7e4b4kE9YjJI7gkqPgjZijWhy8fBdRb5nkSRt8SvFR9aaoCD9sBhuWecwq
KQuiyY90yWATmT97GROeWkzBdjxQIUezonP4k3jqqRcjmsgYt8p/7TqokUJv/CQa
OdHxrNx92C9+oduMxrsBywDZvGTXi+v+noJKDP0wwX4EXSC22Co1EF+neLpyOmOq
mHLNys3dyfqWYJD8ZGOJrh+WEWGHovOy6H6nZe33u1Ikvwj/sIR4rXEe7ue4WFdH
6L9QVEcAGg0gXp+N06iIpWpt21KoLiGsccchYf8byZDoTx42nABesDkYLz2cJ6yd
SYlwcbDUS3b88+pwcozeWv59MLwzfZhMLBRGguyBuWcw9RBHoy7s/zw/CMOeBGxN
gUX94lczqqCSdmkeJgBvWZ8YKCtBvrNyxIve9FKJkrogMdFM0cL6d15LCiRC5gSJ
S+moqa3S/9Q2kgS0E7asoo74naBXYAPfLhFqzrOMTkc6HYldUeleiu+TXwMTzWcd
9ywEacMkLJ3SkxVSbq7+g9E4L4oyqIlTisO8LCMbVYpWcyoc4K+DZwdLgOd18Osz
O52c9t9QkfRGp51zIZxwwFD2aWJDMUXkJGnfN6ib8BPkAQpn1l5DVI3riUeXtWTy
llZYjh7KzbYNQEdVV6hCocBaIg36o5yh1aHJGdvs0dVgv+XZ2FCn4JwMFefWSJ6D
7UW1M1TCVdeWLzTAcJuIPvyucX4DneLymjyZKg2I0VjjY+OrXtZOosLBWO06/L2T
06xW05sA7Y7RoBDRkNO677hM6lxley3SxseWpE/EK3Ejp+NoVI/YZId4zWyEUnA5
aB1wpQHOdxTeoQny7KIk642CnNA4ksIcVfYMJHeF4jrzGJlmO8Miu6wt5/6xr0VT
dfYlmxu8lKiOZmGV/8jZ61ckp03XO20mkfl/D1SC2WrFehtkOEhZc3XYCUYNN5dm
xgQpNO0DcS1esQoywyfTDUr1WlDqxUiEznVxBTF3FBJVnpWGaOOIqJHV2YV493ff
kgCaUsazAWB4ZI2yvM2dQ9STzkSb/XPuxvBaMAeEGbHgXInj5QSGAkl1Lr4YMfiW
14JU8+q+uxfSjRo0yOxOy4NgIzh0Xcht9LlGt/bZmXvbC604o0M5NKxtPgnlp3wK
iEigqpLcetkZBUWRu32EGJ60Ym+m4ZZq6Z3SZ5bvr2QveLxwDKVDUjZL+Yp3yB5a
ilQG09VfcGowWK3sg7CbmGFo4Knm/vrfPakA6Oa6+286maggmbD7AKid6jdYljCy
fjyyYyect6Ggtd7PuiM4gUNq5GhEiknOllHkyBzNsh2Ew4NVFKC3ah6FUm7ddq2U
5AqZyI55vbLm7fAOuU5SJsVc7qzUt2OzGG6wZWiEvQEi4vZMrYEHi8wAp9f1NzHZ
dx1kg3WnxwHsrJEGfuyAgohELzN8tEsKtAUBvkjja9OCyQPPCil3LOzFwewKMfjB
jzvhejcq9F5JF/ZtNxS5hSpczVgjqfQTuHqICaF8OQ2GfxsmHwGYHJUbGjNj8/ZY
eN+vrMU5vDhoBrH7UZVRH8c2/+dBBc1vgkX1JIaoo5suQnwtSAfnJ8UgUfvN5FVt
/+swfZCSK8qCOvncRHW/WuSTdpmWaNpGKUfIr8ZI+Cb9JZzKnjvGSYkwKq8h20rj
akXCCLbbN8xTidEzt6ufpi9fGQA7FApkbGMrwV4XrvtEiE+6U9sdu6U0gazVtHLt
s1J46dc+NESi15bwEViS5BRV06qH5+4Zj7lUNwIVVj9UKSmCy2Is5rztFVcsrCLn
jflgnytfRi2RYhGJ8Bzo8KRqscurijnDjrzCimMc37tnxlKIPrSmw/2NmMhbaY7U
bysDBQvZ2JZqmevHsM2JJaVt7266vqSbdJn1NLCdPTIQh2+o1cbYmzmzWIItgomZ
6Dv80A1NLjPnuISHX76bpNOPozG7m+eb96aDGsX3omccq7ygCj2BqL/aFSmUEvru
m/5zwWcD6pi5HmjerpDNM5mlnwHTUnL2PjQYuxYDpwQVR/ITJJqcK43LlYZijqGR
2wD04vqGJwSf2Ku2NoLjt1PJViCJkl5JEPPO2T4mF5hQAs9b914Hck5wgV4CoGE1
g6rD3NMHQAouGIKDGJCMRzm0IjEZSc0dCbT/XPTxa/O4x4z5uVe4R7iliYYuN3ve
/JU+bH1KolOb3BkYRaCEQOKkAEiEpBX/+lcV+NhSB1OA29OSOWoxr4D+JWnvBJS0
gs4Q0YP6s55oCRvVbRg2YxnpPJqWoJMk+giM4cLWoOwOYryKJPBkJU019+LgWd+X
fmCH3j/AsBL4rlc5nbYGiI4XWjKmR8E6A/WuNkB6Xxxlr/l65ALiiGNjsEIgydmU
4zqicOxsbJSk1PEKKyvJUidzVCOMSwdcBBP8P/g2CgX125AE4psOdJObS3Ty/GgK
+rpHDvWd2i5lpowio0nhNK5ZAy5AnYWD6IAJZ4+wMjl8LG17XMHuht+GYXjF3Usw
lT3EC0DduOyvbdw+ala4PbnZS5vCMQOVNDNo6XMeBmPVmCuw+tJo4C4nnIKE+RVI
A5o6fM+ky78NIQR/yJXlwnTP96XnXtacjYVz30o5eD13GomNH7N5GTP7NYGZIClE
5ZRnIkMzW1qs2ciJJu+Fu8uto6xHFZvcspwc4VXrDfJnNaQa2VcT45bJsNSiiSoi
b/b3yVzpdnf8XM89mi1VfoHbwZSkmwqJPhNUEzM4oAan/00ufddfyc2ZQEGffrZd
vOEcbT+dfh+tO2RqC9WWiK7iZAyTfBpK4ohzwmBL5xFGKbSs7jImSOnPkgwgWFLL
nGDk2eWay2jUuIbLhDyAjSW2zl3f8x57z4eoGVUImCq793PqysrY9PAZiPbfXHOG
FEt8EgKUU84AiIl5m1DSFansuxkfcwhKtYK+Pb0N1nF/SpIctnZAvHeYzCdiGPeb
97pc6LcOa5pcnnCA+TIsALdPGXIdC0QzlQo+lw3wx1Qgi8K5zPT9TOlmI77goZok
R8CVP3errhdNylQ/fxioZAQxASD/rzJF5wnl+gVHAu6GPfjwphsbA1tEQw7q1evC
MFFDjdv+qfNrKKZ5czbRdjy4hAWn+58TcbLEQsO3RmiP+HgFdk8b7oTDW/TbVkjx
T3o1hYPPPblh9nKHhRjMlgX2Z0HD8WNfE3jSZyh8aKkv0DCW/SHnTGsoyuQXepzt
w70m+ljVZD57SP1zfimxu8yTsrrAoiyzMw8C+IBm2J6ejPxLKI2hdi9Y6bMpm1f2
ikZXKM5EjYWVWFklDgkvNwtEf3Pm3Nqu/WL0twLlEHm7oP/bboOK4kN57kwZVFyw
gUjiTgFPmJTKHyWHKkZnYipFerTvo+JYjk8YQHQfS7J6RHB/HtYGZsp0Z1Uh//RV
RaZ4oFsHNIhk3iH/hq//K1Z0lb6waDH0yX5lmva23avua5R99wfqRTga9EsUEQUY
FkX8j2f210SlccWdYboVzQ==
`pragma protect end_protected
