��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW˰���b8Ԓ��.���걜�IO��G7?TnKq��U��?0 ̣���;[�tr��F}�S���B0��%>���t�@�\խN/�\��n�Q�`��bO�6G�5�BD��'y!�ho�o��켚7��y�p�p�^f�>3/��u=y���Ƹ61t����d��ҹ�vT��;�hn`/}��C����Rs)��ajnN/)c	@� W�h8��0LxHE4���pOK�Мƚ��
�&��k�!�W�W��ws@���5�l�h8��'j���*�䞗�/���c%�G$�B��"�=���3Z�2����P���"~�)+��P�%�}�������4�D�J��)N����F�>�C��#"� �LT`�����&ƒ1�[��"��UE�߯�@äh �#��9�ږ2��ܷ3�kf��4�b��1S�
	YU�;%W��G��mFh�h��h���_1Ա\��d= j����I�%�!
��� b�Mtu��Q�{ �$��m����^9�F`R���@	��/�l� ���l�6��(����o��I(��)�]	 ������͑��R/^�貵fr���]���)��j����3��ebT�~s�6��t/�$3�H&��m9;ֺ���|���
�Բ��H>#�S�(�r	��|F��Đ��c;2�Zs,���[S%���9ZSj�����v��C�U
m{��3���꜄;	������0�NK��v�����W�+�]HN�6V�	)���殭�3Ղa�����ԑ>vA���\u3�|^FdX��e�Y���!`XU'�a����i��v+�8�c�L���k �Ә��=`�x�.h�?�E0Ҡ\xuHW} �;�]vP�&�Ѓ��S�?�)el���������0ߪ���V3LIbɎ�9�;��n[�h�:�pj�H1��=R���I)�|����=� �|;:��O��BC�����Z�Q�3����f6���ql��c�	��2�"���6]��@�Я�|��닟�(W�{�y�4��C�;t
 V-��!�ņ��p.��)ɘT�1 ,�2	�Ty]T48�f3��`{X�L�Y�xm�&��.>��$�8u��8̔Zyz{����]ï�'j��^=����2�`���0È�|-\��C�$��;`MP������h�uDP>	�m��R�F�]���M�����/D��Ʋ�R�FZ�|�y!x�Z�����4q�0ϓ�P���x�Ӕ#���F��m]�1~L'��֦�# ��xOg�5G-G�l����z��6Y2�z3*��S�	oj��TM�K���T[���[�)�R�b��F���>ʤ���.�H�i�{#·�X���  ,�r��g"G!�Ot̘�J�J ��yz����U&�_���6u#�B�R�L�y)$�و[s��he+Q!�d�y�3dO���ԙayr�'8��D��v4`���Ϝ��(�c}ƫSv��k�)7�����%�K?UZF	���
j�v��ȋ�ɇ�#��ك���4���rG��$�f���`����:4*2wX�ܮ��۫��&�����.찌as��=�vS�c���Q���x�t��A�tȮ��1�2~hD3f��~�/�%��o����*׀�E�̑�ۅ���*�ּ Z�d��������yt��ypf��x�K����L��Q�֋� &$�ϐ������ 䪵p��?T��"m�/q{������<�e4��Ş���`���L�c��B�?U�ZT�D̪�i;D��U3U*l^��G�6�ͅt�)�J_���	��l�* �Z�O���<�L��߼͉�,h�s�y�$�drZ�xd�!7)L�	-��Q�/��,s��6<�f���2�G�!�T�ȸ�)Pr����rfZ[@h{�VK��%~I%���x@�l�^�I����\5*'�Ꞹp >g��0I,�K1wo�Xml}Z��j��'K�H3�����غѤ;�w���ex�v����GZF��L\R���.�Q ���y��E��_[Õ���Lo����!q>�E��aC��<�;��<d]"{�,喬�>�=��a#�Wtʯ+�-I�� @�jU)R�t���� ��_�����K��OȂ�:M��	�5"�\��IgcB@~ّ��@R|]Cv ��Ew����B��WeZ��]���/��Ju��>��5Rr�M�f��G7�+���F,�А�i�E�5Է�/-K��h�v����V�t�n&
��~������*�*��.��̑Y��	�K��b9�B]K4S�s��6 ����4�I"�(�uZ@�AP���s�/����j���LrH�$�jŹ��7l*R�7��w��Ԕ�_�K��m��I�~j��(�5�(�@��<Š�En��oo��q~Y'���?���j!/IM
�M!ߞ�����.�҅8b2�j (�J��U�Q�jROi�k*����&^%��G��X�R�б����zHS���e�R�5���O�gw�&����41��?�<�O�Ą��>ޖ����7ib��˱�)�����G�{W >�,税k�S�8�a2:��>D^�+0�:�����zԩ�C�ޞ�{��~�/n5��$�f@�=t�+x���������J�s�%�>����B�{$����
#��MB���$J̷�?
���bV	��m�U���ED�C��iOY̴"m&���1h�/荁3�5��]˧]�k ��rT��zm뉟Xg�v!$%<R9r�%8ux��Y���D�+ߘ�MI���;��d������mkֽ-Aa~Z_7�	���Ax\f@9i�p<L.�6le�I륇�_{ (�8�ܤr~���\���;z�Y������p���(s������h����
U�]P��l����8+��Bum�Eʰ��>`ʒ(�ԛ	����kX�l��!����
ߋ�/�sg��^FL{��I��qJzu�z,b�?%�vu��+�^�[4<D���̅2sg�'�u�N;��ZiU; �s^��+F񏽕��tj�l\�����s�(���X�AԟF ��։��G���K�(�U����)G�9,EgRU)�j���������R����F�c7\�n�S�k%�U�y�5�N�.x���	u|и�Wh1�O��SM�@c��3D\ �	4� �5���2�G�QDT2�+$�@���I� y�-rs��zc�
k �Q !ǲ̕�"8*����fJ�ð*�H>R1:��տ�?��&	C�a�:�Ϫ�����r -�n��$�fo�@�J���΋����`��>���:��m >sV�l��cT��AE��t=�߱�tI���2��z_�n�K;����(�A[��'��s+���$���uE�����R��1*^;&K�g�8Fᒡ;�'��;V�5�����p��c�)V�{5��NQ�C��1$�����x�z�0�j#bQ12ig�m�~�ƒ9�J&k�GG՟��x�~t�m�ܴR��:t;�����R���D��/z\͋u	F�VH�1�\l�=3�u���PD${��Us=Q�=<�F,66�� �&y�)$ӼsT����c#��6ʥf�ڝ	�oj�������,Ы7ӝt�ɭ�}�5T�,����:�U�] �.*_`�J�v�^��Ś��.�������4@M ���j�� >��v����� OmV�E�zٴ��'Sцh[�.��?D1l�a8f�t3��46]���G�����g�W�\�g�����ّ	�zzSnGY�gy��zGb�/D��b3��ݦKR5�(>ާ���q@o%��g��W��?��_W���<�N:��7�e��\1��ʸh<�"])i�G�������	Z���u��EFk	�a�SoF�;Q��p�L�w�׍�BM�?Dk5T��(�usE��H]�y�4ܘ��ut�(6��YF�ֶղ�{�q��T �h�����t9W[A���0��kU���r��7��RR�����ەw��:\]��鱻U\͖���6F���H�u�چ/Ӑ�H;���e�u"�p�j~��N�<��c�<b��u;���#�gu2���;L�4��2P��TϘ�@�W�S�giG��2�5�3���r�ơ�8	=ܖ �w����:�6tJKPgh2��M��v�R���&��'��wK����Y�J���!�e�r۹� �Z��a �V9�m���D#�u�6�N| �n��&D8X��n�|�*�>�U-�H�{m"���|���'�9��<{g�4 )���]$�D��J-��	}��ǅ�*vNu}F�eLi��o����ќ]������=�7)���&�@|kh�����v�j!�"F�JaH�vg���=��g��(]���n�w��WN�f@�]B�_�v@	c�U%��j���ޒPx���R�F�t�c��"?�'NW�m���,"�`��o
6oA����WZ�p�|���x�xs( �\���P�G{����C�B"��޴O��X=��7Yo}��%&ukfB�~]��R/Ԃ�����'.Ic�ey�0���|ȷ;��V	8��7�U����]�Gf=�!��+��K���Tp�X��Er=q�wV,��|�ddz*s`��M���%�@�9���� ��[�Sw�|������u�I����z��~���g� �сע�LR(T��,p���C`�齕��o�����d��X��J�H�"nl��	�����(M�/]5����t�F2�؉�R6S��]+!�D��o�����:LYu�g�1�ϫĵg�L��C�2&7���������Kt?gP���u`[�oj ���CbdV|Ω�=�Bo;���3o�y츰��w8V(�&��T`hC#M�U�~e �?�(ȮvÅ{���Z�40���Eɑ9��'`�I-ǪO�6M�9Z�M��w(׼&`N�h�e���rNh9-B���E^�PL�<�
�������K5����/�
:���.eޭ���q�<{�#��C6o���O�'�*R8�F�>=�Sl�n�V�d�ϲ�s�e���~C�9q�wz+C�򏂙c�V�n�ם����|�� �E��Ӱ��:L�Hr��E`|���0��ر2�ī|:l� ��l���v��̟��EB�5��*�w��b	v�jc�=�?x"���=����G�lm�4�9i��7@?�@�A�2������D�����QF��F���#Q��@iT�b �Ґ��2�8b��&O�Aj�"Bޮ�Z�+a��.�fK#��G�k~i.E�)Q*���D-��,�H*�y����z/�����p0���6`����j���D��0�A:�����$�U7��VՐ�k��S\�`���XB���A��̟��@����?��d��؜{����QY6�Iy�+�(�{R'�����q.����9�6�'[�@�{]9�������"J���w���gX��y��ͻo��({�M�.vC�l�|_xx�q>�WN	��e��R��#�.8����r%\_9'����j$|#���'�|��վW6�*�[�����q笡�r�ν=��U{�:��R�Nur��h߆�����C�����ST/D=������E�?�L���悞�ؽ�{W\�
��Ɇ���UO�lS-�0@OT�#�պ�WDq45>d'��℀5����!��FrI���j���5�c�E���|m'���
L����]���J%H�M\��r�MQS��QR����k�J��Zx:T�y�x����F$+/i17,ݵ��!���TI�?�2����F�{V��ҿ����b��Ϫ\��49dy�B�!���j|�i~;Y5D�+Y:��3%��q�fi;�׻�Xҝf��uA���<��n_�� R��
1;��)�r��b����e�]�� GLJaҋX.JȌ�dw���L���:c �
�* ��tQ4j�sq�h	�.����0�dۀ�)U������4}l�G��.��d� *B�}����Xo��oX!�h���4������p��9���jk�*�7~���-�9Ӌ�\`i.+Scw-hI�-����dh��F汛+��}�� �n-�"ݝ����#7���:��ϕLV�/���A�mMP��R�����-��v��	�^���.x�@�>��ެ(��B�.�t]��)#��-R�eC�x�&���5�H��u7�H��"U�]�+����o�6�-<7�c|L���  H-�����!�Vj���/W��^o��< �Q�qE���	�¤�I��]�ą^1�[g�zw�<�W;���u�Xt*�"��,�"�L�����Y8t.!�f�a�<��.o
���{�1P�5:�����G�=��Ъ�"����\�kEɩ�1��H��ң��+�4O�H:l��єb� ��Z!���Xj �m���K-�f,G��~�zY"R�s��/�x�(�J�bC����]E��w.�ei;:���Zy1�^ܨ�\a:�^���G��C_q[��_�^�}3�nf�*�zx�_P�����n*��%���% y�5��h�z����_}q22�1������T��������Ap$�c�K��dt#���Y�N(��V�}���h�ܖ�m�8�{�Ǳ�&�mӼҪ���b>���:n�~�o��!A���%B�%
����s�>��L/ة�P�-e�+{_7F���ՈHW�HsJ<��]�p�a���)Ě��I�l����vK��[�3O/�֖��
���d*�QN�1Y;�0�/C�ƺ��cI��e#�Ї��O��\�m���V6$� �1���*��Wi�B��oP�p�����Uy��a:U�4_����?eq��������h&4��з�m6{��ԆF��;�x���l�(�;�S(���e7J���8	�y�
�*4���Ȃ(B}��i�tɼ����Z�� ��3�i�vTq@�]��U�<'�S�T��| ��K������b�6�|zo�OoW�ʱ����0_q-&`�r��n�F���
�N'��y.�V����ڢ���r�0/�����?�Dx:_'*�jǪ[��g���X��p��p,��~��z��3Ctfb|l���cC
.͢
�4��n��F7z �ޑ�C�$%1�C[��Չ#Qv���b}�d��@?za/�
k��W�J���[��*)_S��*L��lfc���8�x�/��8��>v��������2DB�oXH�$������e����&PP�)�k��y��W�7��G��q~�*T���&��T���4�>z�I�+f���U�G�����v�S��"k����B��l�o���)�7����7���&�b�׃	��^�C�DW1k��')o1�?SĻ��j�=�
(�a�ۺ���+����х#!zB�>��8r��œh�y��t`R��1M(=���f�U��$��&��=vX�ʾhҕ;"�g�C}>���?�v��hс�>X't6��pW�v<(1wo�WO���j�#n��&u�h���81��'%)\f�̷w��j$���
2���8��Ќ���
5o��GH�d};���L�J��;���"�:*4<[�Q�������������rtb7�{� _Z,R�6J'��dg�Ӄ±�:�v�V_���?���Q��'��=��@�P���!�=����+���0EǱ��� �9�5��]O�c�}M�Tv��4��#�w�Tm]Pހ�w9V�<����dq��Z�FF��c4��?�*���m����y�L:�pysr�N�t#�4D\�Ϝ����W�.�:�<�я�[ ��CB��qr�IB�	2g=G���9=��F����Ј�]� ?�8ar?���vx�����/�¢M$c�0ٿ�܃�lg5m���S�\����������mٽ��"�l�nv?���$�� �#��z��U���'�g���'�l����S)01���S7}cJ\�c��Y�گ���1�P*�5�RZ��F�}p
��9�;�f 9��<5S�}�n��z�JU��$�ޗ�&��qI��f0G,��$8RW>�0��Y���]U����{I]0��;Ը���'!� ���~�{]+�Ƨ̆�?�� �\���j8*��5�A�0��Oۓ,��yS0���{z�0�ؗ��
1:@5�F���X
Y�Ԁ�Vہ������g06;܀��9O���{Kz-���'�����8Llb�ڜ�4ε�oa$�C�XjW+qe���Q����R�r���OOT}@?��x��=��+����T�D���V�\8��QO	%3��&sV�OJ���<�R�V��J�1�(��((�����[��&Ϊk�D#n��eU�9�hv�.�X˛4t*��Q��;+��t�T%͉@E�xD����[,J�Yх���B�gNs�^����v�����`��_�w�r�S�0 �1_*#ܐJ�����vz�Z:���P)W���I}1N�F}e��-���-O�A��DCx= Qe�A;�$w�������~�J�����F˷Ef����$&EF�J9��}��9�Ӭ�[��'��IÐ�����6��S�U��$Haq�m���s���#i�����'��X�)��`�s��N���`2'���B�L��#HC#r��4�*��.D#�h���������,)��ʣ��%�F�K_%�E�y��zҸ����܅�+�X ���@�(�!_��s�ĺ����7�5�U~/y�������V���J؟��������aN�T��(Q#{��vмޔT�20O��6o\�q��<�<MN�Gk�[IIӑvDa*G=�����sx��$o����D�²����TOp8"Cq9�rqÍ<�82�N��P3 �b��P�_T�h�ku��D��DRjj��YH�Zd�hf��̯.	�t�?��syT��02�nڶH3���f7��e���[�\��:BLt�C�~C�`凣���-��H���i���{������w�����`t��U�B���%�ӡ-�o�s�K;xm!zt����J�s����<4�w�덅��adb��>� Ci������k-T�x&�sm]��o�S��@ઢ8K#���16�P��؈s��y���R|͊�1'�8,
�/����zm�o�| �WʚV�Xd:�Zo��rJ��ul�fiK��GJ֋h-pD7�^��?o/f�
ֳ#m:Pb7D�lW�8�qF�]�B���Wɇ�E��Z[%��2���h��H^�4t���fGjA�HD�[;hS�3 Ш�j��c�[Yc.^q��MCG�C~"{�lEȻJ��hP�kOGrMR1q�����k������y�#j2�VJ�K���Q@��j�8���E�&����%�DP؟�W�A��$f/"�*��X�c?�aS��L�υIe ˡ'I�f�B{�d�]�,נ$���Eb�+�@8c�ɉ�/\��`b��Q����+�&{�+�E�PU`�%w	^��}���S�[u&���}�J1W`z[�e��猙�˫Tb��T���0��|8���_<cH�����_�ϋ!��'�>4
9[r3߆�d*��P���Y !�x�1I|`�ӌ�/ia��S��ˣ�q�t	��֕��G]�q�I��a��w��ґ��� az|��CX�q�l��f��u�"�_n�2h����Y���nC`	;��'tPh7��ؽ�<���R#@؀�I�g��7ܕ��>Hd@��w��ݜ�@;��æ$v�\N�%�e�
�~����7��{�I.�YcIt<o�DZ�ƨ}F/� WeÙ	7Vh��8�*Ro�</e���e��	��� �.` ���Զ�P�+�-��ae�#~t1P���8�1JE��U��(�^Zp��^o�sR�>qW�5��
;~����p��hR�@P׏Z �V�ώǐ`o*����HY�����b
��Q��� �֬	������ES����I�r��o���;�& �1F��6�JoaS�3��~�LH�F��˃0�@�9E�̳�Dv��x��e���2Z�����Rl4��Ɇ�+ZO�j���#X�Y�b�sik�ʯ+OR��J�P�i���F_�����&f�q������<��뺬0��Z�:5�Ë?L�A������Yl{I�ss��'��P��eҭp���gU7��v2~�Γ�����������sԹX�h�d\֌�8@"�+�*<YgMНza6�Q���^�����yl;8g�,��O�ҚU-�������j��3��>.��J
�1�� ��H�����vJ��� ��7����B!3,�_�Q@^N�lٶ\�4fu�w13����a�����rs�Æ�*K��S�����$�,ݛ�L/:�܏	ħUy~�xNܽ��g�Đ��;�;	L��D�VPT.���ql��{�f�Q��G�@�R���E5P([}l�h�}H��
c@�������T��S�(k`5�;	mD��
��T�m�&	!�����+�����/g����E�G��BʘG�H"�R9R׌4qh̿5MB��&���!|��gm����)*B�5f�������U������y�п�A��CQ,��iV������FE��ɿZ����Y�щ��u%�ګwU�M�D�A./	��X�]K�u���Wj��\Mlg�d
�EE=��	E`��F#�Se'�%�� �|���#
�S�Dj�����\C�vNha��ْ&�v��~��(�cf�o�W�n��F���W&'xaSD�zy�,zN����,z?���H���Zm���w>Ί!�VF �v�Zu��]�}���>ь���C[<]W[�<�m�8_Ƀ_C��S�C�͗�62���ߛƷ�[?������u T"n5$�`M|f҉��Χ�QL*�	�Ħs�=�mc�L	��S��;���,	k/�fDX
Ĩy�}#+&���[Pb�la�Y��|�������c���
J2b������j�\������Mve�U���Q���&?4��]�enj�(2�)C��_�U??��~D���/ex�~VNq>8.c����m7�4�{��J!+���y�:N Ed�5��lҽ��p�j��j>����x�Rv$��R�10�44��d���3QCL�Ѹ��i^?���F$�D=?Y޲��zMO���|O&�v?�>��J�7�uQ�D��Gcc�Wh%�$�5�(���}c��w�IB��Ux�J���U�i.��}f�J��:�z��F�����o;:��Qh�O%���,̍V�M�O���w��qgm^��1�z�*��Y%}�]ϻ;{��A��*�������� Vjc�L�쑸h�y�߷����܏.�����y�Ykv
/��*���^�f�Y>�m`ǠmԶu�k��[�e�����Tg�_\����{;��P�����&aoAsP~ _�'��tt�.،��d���H.�Ft^- ,���eb��_��CB�P��S1[)�`�wD�*�L>��0<oS�u5[~�Z�W`,آᓷY"�lni����=o�"T|ܼ�� �rp�#̪���",�>Vȏ2�L&�1[`-@0�"��VQT��V��#[$Z�� �"�c ��!���1I�$G��|��_��,�P�Ag����`���4���#_50΍�%�y�戀sϩ��@?tj!��u,bo�����v�%:3��)��_�E�YP$���Ccί�H���w_�e�:��F"��d�L�&2&a�wH*�3n*d��B�X���6+��v&68�gg[����\xJ@d]#d��F�)�!�fu�ݰ3
����ܮ,	#��lw4Δ��b�Q������G�\c�a �z~8Yv�Q�κct@�m;=�PS��������`G��
����-���5<�h���8i���(�))���W�MN�|�-��n�,���ǅ#G��@|�jV�����A�!ӈ���^٠R�Eg�����t١їl��vYb�~����!Ϯq90y9��u�Ƅ?�>K���'%��$<�R�Q������CC�-*|���ܯ�gU3�.h�d�To�Qn�"�^�[}���	�����!1F��3�[�;VP�V�����l��uӢp���T�V4d�9�D�$f�/��>�YJ��"�&�@j/+�p�X��y`!�&20���$�0��k|S�(Ӻ��O��,!p<u�k�A��S�%�cJ�[��Vi|c�.�P���p\��I<�Bi��C(�?�Ers�	�$���%��!�w�� ����w^��X�/;
��7�Xcyh痸�s����S+cl��jFz�٦�!�X&�����x �l�?o�I=6��j���p�#��`phk��tH+sQ.]�3(؀)N��l��P��2��݄x�����3=;۴�5�GVw�bZ�F���O[�֜K�}B^���,jF��[���W�}��Nd���4q�jgn�C@�b"Q(��ot�[��z'=}�P��`U����#7j�^b����������xP�ę{����~�%z�S�Pa%�-P�d�����є��˄Q�5nk�=Y5��oW��/�
&L̥F���Rd�I�-��!'J��$=q�Z������=u o����Q��J3�o�N��I5jEDtn��E4+fG�����d�M纝v�u��%�Fsó���PCIӟn��l�6o��ĺN8&�IJx/�����q��|9Y�Hx���`�(����a����z u�ԗ�(jtmb B�+�f�3{�}��b��T	�Ǻ��
�,iJEʉ�@��d��"Q5�{(�H����~��i9
:dEQ���'8�ǄR�*QLt�Z3�5it�������fBDz� EK	�m��^������!¿�'qMN�H�(U��n��&ԧ-��:Շbq�J���%���i�9�C��t�!"m�0?�>�5�FJcj�Լ���B�٦i.�Iy�#�:������Wx�c���R8���AH�c%lb�o߻�-�����Z��@vM� grs����6�w+V^-���yپJ�{���Z��Sj�XV���D��"�iI<�ִ��x5E

�A�~,��Ӡ��o�"�Y���Ӑ�}~VY��*;g�YOњ��=��\K^?��_��*�����q�5�Cå��([��x�lu��� �D�\z9s��1L��&����3S�I�X�+,����G� ڱ���Y.'w�&�D䳅��I���+����M�Mr��Z��%n3L����, ��TȮ�>6-�ou|a�� zlX:q��vH������I�/�m'H^��-���V�gTx���6��g�ɠn��ٿKj	}�i��P����l|߁�$y:�u@�5%�^s�)M�+�M{j�Ӟ9E�����q��Y�)��u��w�9��aL�~���n&�z>��>\E���kl²��oH%ԏ�w���o"H����V�A�~�R�2Ԧ��U��w�+���f���U ���V?��*# c��;��|��g{����s���D�͈Z��g�q�ѕ��P+�gT#��[�n���7B�Ҽ�%�i,���b-Qڏ����*��\�S��]���q;�r���,��X~�
ջ)9cPN�3�뢬���S6�U����&ՉTV�k���j[����HJ��_�-����hv�@��f�r�a�9������y��4Z���,;�����\��=��]{���Q����"7����5����3$Ғ䷖}��n��wׅ�R��q��Dx{�ج��cE���`j�\	K�/�񀗡\�K��p�`у��煣5��$���י�P-��{/H�9���ķ0` x��ΆR�Gndv�G;ʎ1/��dg_t�ż�+�˷��亐��Q���|�(�6�zU��Ř�ӞJ�g�����҇/�e����ȏ<R�<^¨3!� ����#n!^I�tg)ME'Z�S�x�G@R��@=��7z��昵�⻲7��JD�a@Q�{%����DM�Ի5? ����U�ޚ��h0�	 �Յ��.?F�Ccg���H��+���3�m�س-0�ň�/�R�B��e��)<̞hS�2ZF�ޝio͇~���m@�G�Ex�c�qX͛�#�!.�� �_c;�v�#��R����<��g�� ��'ֳ��w��\�-ʳ�!z�k�F��Ѹ~����$�<
���q���'��eKh�G�n+3��Q�IIȲf����aي�a�D��
i҇��'�PųN��R�4��D"B���+[��s1�K�m�[��oW�v7J�ϷP%�v��RN_�rzL� �Լ���єQ/�>tD3i:^1|�"���Jm$�� �mf^���q�F��?]7�Q�Ѽ�1ec��̗�i��J.�y�4�f�4Q�5��N@
��А/��5Wsd�Á�\�ޛ0 ���(�L�+m�0��ۙ�
h�\T�k�@<<8�����q�4q�_��A�|��� ���#Y;q͆�V�K⶘�Cj	̉#�;LӼpڣ����w�$��',5M��ys.z~�[2��G`f7~���j�?�g��%��x�Xs$�N�'�o���l�
��� {pST����>�=�5`ۃ[��9I�m����?!�D]�L9z\������Ő[۵d�n���D�ΌH*���t!͇MW{)ޚ.:���m��r6�?J�`P�� )ӄM��
��fy�#Lg�M�9}�Y�"���FђUf����zz�p��S�w�̣:�Q��p�6 LEMIhG��Rk��f8z,l��R�@�%�N.�Oŭ�?��ɬ�BJ��> \8�{���}�샍���|#����Y�Ve�<?;0eGo�keg��?e �9�X��V>.�>�u���M�t�e/�Ls�ۃ�$
jH�G���0��"�J�ԼtB�!��H�Ⱦ���-
;���i=��_3�t�i�$�g��Tj�|�mR�LEՄ���o���R~��7�D��s'�ر��j�C�Eo�߸�cS�ag�qU�>����)Ӷ&0is?��q�f1p�����v%���j�^c�Cm̍�c&f�ש��C�:��6�ue�k�6ϣO�f���B���J("���e�ɹ[g~���֩���#\!H&�g7�;*sp
=�����@GW|o�� Q�7΂n^���I�O�/���{�i$�K0ݶ��O��i^|Ne�@�ˮ���{+���,��i6�OkA:ӷ��3��,��)؇ �KTx��ڊ��	�;����P$|�U/f��"��y�Og�������䄩rI�D�}`�eD���v��4,��4�)�F�X�$����\�%Y{����}��$�`�n��3�/�3����j��e�r�hu/xm�%ˈ���H�ă #�o�#�Oo#x܅$����9^�՛:��:Q@ns��k�Z\u��+��~�b�<�^��y���m�ͼ���qa�{ʘh�b����:��Q���&
@���]@hiiy*#v�QȲsv���gѼ��7C[`f�_�q�J��1�y�i�e�!r�2:$�<(���7l�im΢t���fj��Y�Sk{�G�v�F���m'�����V�3ǆ)ُ����X�^�ލ��5��I� �ը0�}c0���������Q��T�J���'�W/�MH�J���u�4 ���$��d?.���1�:��V
��XVD /֏����8�0R�h����r�^Z@Ã<k�.rvEƋP��}c�����'��9%8�D~Wڒ�R��+$�PCnsDE�H�)�~=�2Y����IZEP�+�e��RF�(�xAW}�$�-�U�/��}�{�ӊ|ul�l��$\Nz �O��6�O.����)�4�kK�`h�b�c�G�7�p5{�a9(����Uȕ��R앇)�D_���� L���{���TЉ�$*�[���fX�hgĒ��)2��J����K�����| 71�/A���
<�%l�,3��n�f`��x��\�9��e�����U����Q�w:F	'����H<˺"u|�����^?8üΘ�,*z�خ�+���:c�����}���4�H ����'.3._�FN��훇*U��9���kQݤ�tq�R�K�-�09��o4��:�aPl��ԗ&G�=h`06���#��g��*-2*���S�CM�8����ߏ O5���<n�Pbϱ���asR���2��JͷN�?ek�,/�г�$��-��N��ր��TDM���֔,+�P��Uyآ�*�2��~k�	|��Ww�Yͼ�6�]�BO����/a��(��}D��[~]�*@;F�U�e�����풄����2m�M��`{~��=�O�U���`�rf{�V�1,]%��Z�y먨�pl>,��EK��4�z�
ȣIQ���M�L��l�il&�	~�YSN� ��u�Q�#+Bx<�v^�0.Hy�n�jx��!����3�����L+�x�сO��%�P2��C��DVV^�f��� t��Wd�ϸ��k��#�p�pd�A�l�{��5���v	˱�H�t�*b��]`w����aa�1�3-�K���ٱ����ifK�A�\��y�<$��[K:b,(	��J%7+�J�(pǦ��ݵ��w���Y��l.�դ�D�HV��K�,��U_5
�O@&2���H7g�߷Z۟�S�EFB��쓼�z,"�����ar��Q�ثɉ/�m�xs�v����aR�݄k9jvhx<�7%-=~kc9�����bb��90�?4鑝f5c9lgC^�_5N�(���q VO��"v�q���\�&����ıޢ�:�����*]��J��ٓK?=�.�,�Õ���f(�L�R&wJ�ݱ�~v�n��9��8pw�Q��7�;�)��AS����Ժ�ͤ�mi�8���\#�EF�U�2�'#x �����g�RE���$z�
����ch���` 6���99ݴ���_�(�"�ir�2���Se�[��<2��`�BAT�pT���>�@�_���^Y!u]HWT�=�9b�gfp����Rx6Q6�@��\�@�"ٓ7��J�\�����r�)�f��� ��ݷעG�N�C;/#z�mݼTc���=̳��~k��L5xݻ7��9�JV��ER��SDE��.�q��>$��tX�<�E��:�<$=X���\��f�+���5/ЂT-c�խ���7��lEA3U7v� L��4l*`ƽ����e���K��w��(W[�����%����n�C�H�W�Iö��)��)&ېD ߨO���� ����w���tE�jIm@3�p�%��c36^L[�ܳ��v���ߟ%ƌ�l�A���(�՘�'��j7"j���n�s�����f�S�ϔ8^�8�J��~0R���;3� 镓�P���55���O�9O)W��~p��х|�՟Q�f����G�\p��P���b	��NI���IZ�OY����Ek&=(,"*&xv�L8�����T�$T�{�5#�2
jm�b�� �a�x7�6HO�=-�Q<>߲3�MF�Q�;!Lt����V^�5��M�3��7SITDK+h>��/b&��ާq:��5Q:�[`f�"%Ԝq�q��)��"z堐����x��Ż����ȝ�+b/b�Tj��*n1 AE��Ӯ��e`��v[�ÌХn�_n�'͹��5���%�_	Z�h�ħZug�-�Ia�Mo���L�D6�b�����e�m&��=�&�T�u���x8`}_����x����I�������i�