��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9M!@eW:�Po��+?A�1X���T
���� �o����D������Iyz��� ���H����t�CeCX_�]�C��W�7�U	6�҆!��K�*)�� IĆQQ��b�P�AI����	�h�2�ޡ�}2��?8�6���H]1@���Z݊쓎�Z��|���6?�7��yX|P.�3��Ě���Ŕ���a�*��� +�ѡ�
-0C���^�4� �®X��x5�J'�����#�( n�`l#ۦ=/���TG�h�5��U���6r2�nqf&��k�&�$�aBA�ȱ�0[�3�5P�v�����<Da�v�ŔSc�44SFu34�fr�aK�/�M���6���vv-�<����Z�S�a�&������67*,.�鼕"FP����(�1ع��1qԣ��Bے��;�����xZ��X��,��"A�^4�( C^#�N&�/ǚ�O�a����S<��,��v߮-��^c�>��Cm5�'�bd��0z����!�w�Q1j�0r�&o����Sܚ[�s�F���w�^l���lp�?�l��u�o:��WT%�G����Kvz/S;`�]E���x{�F�j�C�e�v�9�U�a[R�����5�������/�a�lck�t��;�*�]������R�%o����U�T�D����@�I�p���~d��.5A����yD`Aϼ׮S�l�L�	��QG������2T*�IS� �]��9�R�f�7���Fj"��h�EXeW�D���]� \ʰ�%��~�=�� B���L����6��s^,���إsKJ����	�i%�Rm}D���(�k��(⿞!�=PW ��[�9����5;_���E��_�Ϯ�ׇ�,�<���}�$
�*F���4�Cņܝ�FmHe��
Q����)��`jQBf��@p`r@���O�k�t��) Z���U�Eg����{�i�3EZ߱�o����o����1�UzIn
��{63�`mN�7�3�#��*G?�2!�Q5��y���F�U�_��ED�0)�Kka�I�f3��˞�q�+�Z���<��9������?uE�Ki��-	G8>�s>*��w�~W�hs�Y�c_1d�T�C�%����{FtmS`�m����@w � ���t+x��md���9��<�Z�0��[2����9��m��p$,~BD���攢⟽#56��٤������o�1c���=L�\��GN�9^1=X椧��L�[Sxd�9��sO�i.��g��&1������m �����[Q�x�lE�Lz�rXU�^G-�
��,jb�U��nZ�J��6]���\���T�e��^���ɒ�$�1^$ڥL�H\uBϢ��/�
��`T�3�����N�����X�D�H���"<oO��3=�j+�����'���5�i�M֧�v(ă����Po���<� W�߲b����h���0V�X*� �_��}cS���Oц7��c��A�#�p��U�gj�j�{�mE�w�W�ɟI`�/��:�1/R���`<ć���F�_�*b�x�6㭼,wB҆��\κ���1]Wg���p�B{��F[���wƧ�����d�=�
T����>@�@��?t�����/g�ꮮ�'f-��ڧ�w����a�I��P9@�J>ܯ��5�a~@���..vU�����D��A�A�3.�����`bj�匜��
�q���agݦ���ل؀Laƅ�ָ\鷡�����h�2��Ng�qM� Aq�mK�0W��xكAֺ�����X�� ��)��]e�_u>��/ _łQAr�ZF3�k��c����Z\ʹ��m�&����E	�N���3H�u���$t�]��R+RA�v4�n[�8�Z��z�9Z50�1���g�1�
�	�K�� ���u�o:�G����&<���=�?T��%C��Q�͞/e��$������ۇ��#+|�ѵ�ѩ�A'��_tk�U�g5r����Y;�.|x��;�����p�W��h��Y\,������ ��+Ŧ��E ���&�d}�T�D��Z�[��(�"ܯ^�?��X�e�r)l:�dms�Q'qb�G���x߁��Կ�U$%T��#|�"����+��\|��U3<���R
���1��RF�/�$^�D^-^��Qad�8���Gt)0C���#�܀h�K���fp>�O(��{��i�V��kz6Q�s�8�M���xq`���ׅ��)�I��Oin�'��l�|P4M$֣�qKF2x`j�æ���QWN��~�z���^�uSl�J�˸�����:|���	���jt����ݝޖ�t��"�0;��\Q}��z��/�1���@�*�T��lB����>s_�%P�m�g7���*L\�pv�*_p�f!]_��\��s��X��Xz�`Ώ)~:�QGoR��etȍ��|X�*I�����>&;6Յa�w戚�e��/�R5�"a�.�՟�4+)Jb�� Zx'�fC��x��ɬ��18��jmw�`g���-f���7���m3d�[�fna�
1��J�=���q�B��tLĢ�ϚFXv��F$�a�L��Gj�f�Wd܂C����� ܈nj�|ȿ�Ƣ��Ϣ�5q\%�<�;0���K����!�6/����ҥ�A����<й�Ծ�ҢO��vGNe��}3dIڛȟGL����r��ڿYe�/F_҉7HO�G�H���t������!(�7�3��*� Z�$�� ���تqj�K]�D�e~�E�/$�Y���g�3Zc��i��(8`�1�/�9�W<@B��t'��g4����^���.�-4ec��>�onJ�sI�������ʸ4��S����ъIԵ�e`F��3c���!����DC�4rz�2�!U�se�����<爴�V蟂���/=L�H[��FH�,C~Z��0�\
�R���6X�z��t �vKM+����,Nb�y$�����0�`���&D�*�Qz��΢�(����X�@O뚄HG���g�3�{pK7uɤN��^I�����tc.O+�#1�?G{���d�������h7 ��k���1�_y�����v����,�#��7���}�6MĶ�Wg�E�mq����O�^�E[�+��m�h���ݾ�զ�t��)��^n����g�u !@T��͛<�R�ε>��!��[-���WT��#|F��j�s�Up���f|%ێE�����bIr�x{Su�<x�:xs�Xk^`�Q�X
�Ο��=�����k��.���E���#ӯ��X��:��t�t�����В���i�֠]|���{��Gަs�h��~.�&�y���W�83���O�������Bۗʜ�D�#�"��#���\Ub�w���q�Y�8��NrA�xL��L���;�kB�M�	��=ʢl_������*w,"X�Շ7�閐G7\��vaG����9�gl��|�]�46DK���Ok�]gT߉��Zb�%-���H��O}�������,@�6��3�+�Z���j����5Sm�������D�6M������Y*j"o6}��m×^��j&�p*����jT�ֺ�F�d����vI��/E��L��ԡ�/��#��R��l��N����A��&��������=[$w�hk�i�(GgTi�p���xI�$v��,)&��`I��j��vI�x'�Pg�t�e�L@���ǫqpz�R7g_%�jX���x&^�gd�S�kϧ�k=�����.���EC���x��/՗D�f,ͼr`ii'�i lTΌ
��Ȕ|b�y���\Qh�5��FĒN����f�	^��#U����I�!�l��l����	���8�S|�)*�8Lo�u��7��(�O|A�o�R\��]�����a}-o(k�"�y��eD͜�&��xOxЕ��O�pN�t�rv_L�z��c[c_	UL���ݯ�2�
�<ZR��n��s�-���Q���J�Q:�]7A���8�S��c�
�d)�s(�d�6���}m[��_^��
fO�BA�K�����L����~u����3��
Jd�.����҆�0�V�n�B��=* �ʀJ����j!*�H ��0�<�19��#C�ujT���n��νNAu��_�V�vZօ\���uj#�r kN�Y[_(I|�&�̢�b_��5*e����/�VS�<�I�p+�{[4�!{��rbA�� �y��Ӈ5��Ӳ���Dn�eU��]��~~px!������[@��� ;�{5Mh�c�i��c�.�\ȖVg�E��tc����I����E�u�`�A�}E�����$��Fqs����$^��ψ�a�	=�ْ&'F��K�Nt�������;���r�T��Uq����>�@���A�ld֤����֝B��"����)n��՝̠!��^}������HH�G�m	-	
ԬX�BK�� �8�~�m�J�jÄ5{[�j��ɪ�u%a��
�7��Q~3�,��<;��5Q$a(Y�0J�P�k�V�څd�3ɰ�wtѪ����-D���N6�^i�un��y�/f#�|�b��yo*g��,���5���T('��r��B �����OD<���Xȫ��g8�<�$���
��0/Y�z��V�Ls[	u`�]�H0�8)�ʟ�' �
�qM��Qj�6�
zt�Ý��4q�����E�du�l��],z/�#B�;`�����j�v�l��p[��<�\4���{��.���o��ʚ��6\ҙ߆ç�w�f4x߽%y��q�u�29u盜˿�y@N�#v�%�X�lm�q�&�������e�?�=�F�_~�z��`�߯��b�`�Y���qA���t�X���޷ ��E��P����A��S�5�9��A��ֺ�]vP��餝U.�fYVh��zmk�L��Q��MJ��@�K��!'mf�ͮCi�W{�ԝ�����C��%��sCiv���#�-Q�r��<�󂟣��r��"U˾j|f�zֺ"�p�������f�pd�DP
��Xw��'�:m��,g*�_Ն���8?���q3Cj�˧����d'@;;;2