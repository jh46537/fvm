��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{��P��f��Oz��Q�O̱�� ��D�м�rT��AGpR'�?�j\�d���7`q�h�K���`�k�b�r�MA*t��E��ɘF����K����̀t�i'�)š|�b@�j8|�^\зE@�Z$c �ה.��y_2���K�ڕ����T�^o�'"��/� �m-�}�+sLú~}f���Q�q��q_ r����^�ɰf��&�R5��B�
_�� �w
kMZԟ:"1�C.d-ˣ����x?�q�<Njkc9l�N��n�ڞʛl%q����j�����i�a�#)<pOj/1�L�}���b���E%���_�"B�����Ȣ��Wd����w֖�k X�6�I�Д���a�|�A�+��~<��4v`�J��mF'�u����׶���%14��,
P���\=�F,�|�;$QZ�f�8�Z-�B�sB7�_zh�X�9���Uf��T��Cr?�/�m��	�G(�5�f+�����y&Qo3BOOXq����˹V(d���F�
˂��(��K�O��I%�Fd�N3{����t��`��!��U�Ŵ�(�~i��<.d�;��ҙp�2��V����t���/�X�*�����*�q���H�aѻ�-_u��]ƅ^�����.3�C�a�>n�!}�#�xGA�R�C��N�l��.�	�(�m���Z^+�.V�cj�?�
�A��$�y����#
��^�o}���:��K*o��n���A����6W�;�R��]�0�K���o��%���KeY�ב���4P����b��`7���{'��Ǳ�eC%$��M�x�����g�}P`^�7;�61�Z��E��=-0���W�,�����V�Ǳ�J���ʹ��!C+3��zHX��.�{����}G-�ݫ#�R�EO���/�<K��
<K��J5��Ē����FI]9S� �
ȸfa���#x�fr��]J�G�P�t1\g��/FJ�d�]s�#�RǓ�����5J�	�BǥS%ރA��B���L���&wZ�J0\��r촲J�/Ƌ�����X�[2SQb�H��d�����y��y��.b'�Ɋ��l�K�L�ۤΧA�3x�d��� ���n9����FZ�m`A2�5�=k�i����z���-�F�%�ϼ�<?�/���^G��7}���cﻣ�U�7��(b�BH+!�%S�=PO�-�2%��)��n�O_�e�ꯚy1�����l�	��4�&8&J)w)\�7k��9����I���W���6I"�`p�R
��k`��1C�Cʐ�<��B�UX�y<X��g�l"_����&���� 3BL�엻Zj���m;u�1N6�EM�q��@�3Gлvg:N��H{�k0���AAd��?
a�0T�-�6<߅�p��DF#.i�u��INj<M�Y2��N�x��z�ЊȞ���V�|xn-
U]�7�u}�us3��E=��s���KW@}�24F�D /=�5�[�^�rl#���#�9�.[s�@c�"��.�k�$��r4@�qB+Z����V�!�� ss�{�p�#׏��n�'\�>
�L�<(uV�����sAb2���n+&<MF��q>#������ҳ���J��������,V����s��}�R��kb r�-�QveR���ſ��+�Is��f� 8W�?�y4���� |GF���j�h�zY,5��E�z�qT��g��0W�*�_��i�}W�޹���)�QA�r��ן�?�6	t�1T>�[߻E��kuU���_7w��4����2X���6�2=�q�< l%!r� ��N`j΍���/
�;�t|kSb
�&p\f��(a���iD>�A����.���V�Flpq�:܃Om�<G�49��&蔹����?��|Sݲ��]l공Q�>\Lm����~a�+>���\%����h2$R�d�Pg=��� mEٝ����i&㊃G��������<��K�����a�s��Q7�-g�Њ j�=nb�z�쫎����ѻK������H%��G���׼6���'�smc��A�`^�Yz�67���Mj�"�}��L�Thr[[�B�	C�=��Q������1������B��^��	ڂ�	�6R���G����Ӌ���$��s�{��U�[��$� �Pc�ldu����r�t����M��;���yq��m���)D6�W�|İ4Qv7. @��
�eo�K]�n��b�(\���|R'��	���x�Z~/P�ż�9�����p��"�=3JO�Թ:� �Q�o�6=|D����nx�Q���J�~޻�f23��_q�퉴�eoY�u8�=c0d���+#��4��I�83
��ϏT�o��C���ӓ���
R�m�ܱ��X׌q� �p.F�0�ۼd��~1*Y�ՍR�A��k�#�:��`޶Cz��S�`�-乓x�Cu�N�۞K��q!�,ն@�[���z���O���ae�]�'��5��&�}�Y����Lwf#QG��{���HB�a����3�G��A��a� ZoM�Q�=��m��{��i+�IkIܮL�I���Ѐ�w�cחk��$H��
a�h
	���DB��Z���q"m�����(�1�+���.�I�-�G�� wa�_TYrX��Gǚ�8À�<����y�JϷS�X'��5����0�6�;s!�@��]�kh&yP'o�.�Vx����;�/Yz���;��^�ᤖ�H�簙�UT���Ds��5��nE_ˑo�^W!$�(2�Q,�7�4�x�Z� ���}�ֶ���9����H�1;���`�bST������[�%��'\��,�=is�!�Vq:��!N�)y����o\S������ȓ�@p�[:ć;���^X�0��`�a�22V� [N��w�~B!%7���B�e,|��`3�dA����B7�0��� �G�H�<[_*����L��B�Ro�FZ�"bW��!��]He-��`~�_D��G
9�ك�_&�""P���)J��zH�X|���?t!��Z�)['4��F�-^=�D&cl�ꅴ�&FU�N0�摎�HLF�eF���6�澏��"�ph�3����0�ܾѡ�+�ƹ�-B�f�~��xU-���m���4���i��tX/K��B��Q�R�]1���x�@9`I���֣t�T��ة0"�a^�%���{�W:�5.���mh(��,b����d壅3���ܿA.�~�I��m6j襷4�ϏwI��'��L?\E�n�k��H��w]h��%���+���{u��}E[펵���L_�����'�l�܀5o�ў� �}�?w��Ķr]��6<��X�7�^YIu,8I�&|���D��:.��k:��E/�N�q���o6�x�<Vu��L�-K�b/ƞ�������쇆"�������M�v��B�Z�f@\$BVA�(o<� ��`�B��Zr�E�3�|z{�jľV�M:��b��J,��Qec�͝�V�_�0���;�v�IĜ�	��%Ѿ�#��g�yW�:��^`$��Hn�J$�a�)�3\ok��m�<
��_W	��m�`;:���s֐��}i4�!�A'��!����En�z�J�)Rr�����v�WDSղ�b|,:6��Q�!7�[����Ƴ܂8Z{�m�m2rS�1�NL�Y��s�W ���;))��mS�/�%������ށ�q��>��Sm��� j�t��n�T z	4��b?^}��}w����̪��ɖ�h籴�7�Ի�4{*�KR>��1��	W{NB��@g��˗�	��Cq׸�$��4��WBo�k��o`�
ȥ�H,x?��T����%�5	���Ͱ"��B���Ư͏�����]���j<�g4ǇJ"�����u�� �>�߬U/̠��Ů�q1Ѕ�`(�-��:>�z�:�e&
d�I������"I&��L�A	E���ϑ�6X��FC�~�U ��?����Ņ0����B���}�6.�Oi���T��_�:y���z_r��DB�40E$}~�d U0��c�'�&�īy)M~�� c�xw5O=7���b�ǘ����'�"�:���a���ل�[۰�؜�yCU+)�	�,�J?�V)�P��VY���u��TA�Nd`YQ�*�LRlc���?^+хy�5���9ǲ����֧��`�sz���9̈9jnԍme��[U���D@;��{��ܖ(�X	��!��mYh�l���S?�a#��p�
E�hQ0.� �M}�w�j�Q�."ܻ�~������-܁Di;�A��GyTv�{�	�@Ѥ	]�;��i�(I%�v���/��ڑt�g�tS���4R?�����f4�i�m�>X/�8��{2ߌ����P�^�D���n�O��3�7�2b������v�s������o�za��7��"�ľ���I�W_�(h.E/��2�9��a�r�r?���v�[���V0�/�+{7���-ZE�^;��s�v܆7�8}Z�9����L��E����`M�ul�{j^�����RB�|c�ΰʁ���:��k}�X��AQc[�uhL8��SVJ���b3��e�hT�eN��46 �\
X6=�騐[����3�w�H,	��;�Nt5䞩��^VmLX�v��`Jۧ�@{��<�<j��� 3N4����:�P����a��!W�a�)��X����e��B3(N,�������a�ń*e_��/aEӘ,2]�|Oc�O��k� ��Ͱ�͋$y��vn���������K��R�Ȃ�]Ǩk2
�o�N���.h�VP�*�a��r�6��@l�;<��.���
jp�h��;�z ���#�Q��{�2L%8����G��|{g�캮��C��W�@Į��Р*���;�̑t�[�*�6${���[Nn�����Q�X�)
�`��!W��6�?���T����PD��?��[y.�E� �4����3��������+sѽ#7�-$�M⊙�������ҟ�""����ą��0���,]S��/��5�3)h�0<����I��Bk�o��e3a�M����	���U<�&9�/��g��O��MJh�0��{�U �6�Q&�U,�=B�N�i6��w��_2��0+nи�=:����)X�^hgٽ&�����E��o�D��l�֏X^���� 7 ][�%�<����/�.�'�e<�9k��mò~�',�F�`�3���6�<��ОqA��.h����M��>����P+o�7+L��i��'T���m������e��,40`��8l�; .l4���&��0��,)e�ݷ�=s�n
���g�O�kN�͸�@H�:�Y#��+ٮ�^Ȩ������o�-jy�շ�!Eo5ƾ�E�\�)��᷌�%+�?B��,t?Sz0y�G�I'��w[/F���:��H�5����J��yZ�Ҍ���|���͠FW��@94���^A^��n�CZ�HB
q���M�.+�5��1���qf��Gv���r�'�>	�>P}t�	0�?-�����}��z��:�nb(V'!4e�@]�X������7��zi��H�݂*d#s
�j������Ue��qm��%tC�~�I�䷰���]�β^C&9�7z�!�߾���K��$`4��fr#|#V�i�������E�\�강����tz�u���BvK�nr5����*�H�C����K��ࣝn5�(>�۳��q�{�;���^rcXN) ��}dx�'�px8�#�
�ȃ6��e`�O�E!=:j5���p��fW|$�9���ڤ]x@ł��kGˮ%ʖG=��`�`���x���.�9jZm�]��L|�j_�;x���Xo/�H����襭�=+��	e��N0.:h��/;���V��П����2���j�ѫ�k/v	�ݾ�EB(K1� �QϟZ&�7�<��I7�819��a(3���&xA�?m��bpyf��� x�B׆�ј��g�����1�Z�?���^�����7_��C_�'$#�]�o��mD)R�Zɘ���T��[=��)7T>EQ�C͓���v
�%��=$�Š4�]�����,4����G��[��:�*U��K��:S�ۿ<���?�X����\�О��s���j�	���%�M��íh��cGK�!���+`�Е�@'`c-5�-���UE掴c��#~�fu�!�샬�fOM�L�1���i����d��f`�X�T�j��]�$k��u>��u���J��T�� �y�'�3U���bL�C��Ix���Ǹ���僰C�lƫ`�OBu����� |��̔+�l��թ2oF��¢[w��_l�B=j��z�dm���7;D<5�����a2o>v�U:7��{�Ot��n�y�/iG�vo/�r�GI�ަ0d���`��F�^�4����r��?{KٟK��T�d����#�˟���6��M	#�2[���0��.L�"T������WN�,�e������ܖ;Go�2��G7�4��}���hes�Ã���F�y��,5��0��H"��J�l;o�Ղ���(/���)���"*�Ŗ��]?m�N�ɓoz�>u�-~B�������a�5�[%���+,Y�T�\� ��RtM������b�q�5u��C}��b��~���p�Q�>/	��G�e���Ta�B#�V�tc

��@|<�5��(X�4���$Aܔ>_�@:�]O��B>�Q�վ>uF������=���;b]�^\X:{�l*4$K�@ͬ(�pr��q�AJ5��������	bb2�J��RՈ�&������aMI��up7�<��]' u��\��r�.��:�6Ѷ3ZI��j�O�h���Nj��r[YH O����-(y�~�����AvTΰ|7�����۔���+\�o0� 0��K<��t��� "K�t�P�]-TQ��쨼� D��ɾ,`5S}�k��J��x�_�0�1q�Js��������g����8}R�95�u_X\B|.#V����͢�C%��i<��q����� 'ZW�Xv_}x�p�Ջ�@��]��/i8����Y�ieF�����h�?��3��Uz�{:M��P��c�R;bD��3�C�]���ո1ݞ�d�$\���dBF��uaK��e�(��
kfBͽeD�Τ'�Ha���d��1`>"���r���v;�x	'�����B<�^!�{�K+�b����WS�Qâ
�ݯ�@�����~i�o�R�~[�ޡzx�hD��S��V�>x�3]�ڐt��' ��}���J�Aؖ6Ȗ�$� �q{8��%,ņ�2��~@l����%/Ix�`���a���~u�/ނz�p�&Y�Gn��Ӧ���O���8!"��E��[��V/��Ar(깖�z�c�a �G��8����-��'㌄"�����p�*I_�'��_9�����l\���2&���ᙽZ�xW�M���y�?�WM0@x���+^$ j}Ɠ���ħ*�-I��h����QP���n�#O�D��c���"ք�BY6i������)=�i斁O>�|�癫؜���ԣ(v�,�	���#�%�õ�����P�P�e�9��/ �0AhzT˓\q�VR��j?2��@q3�)C��l�p<�DE۫8P�V��Џ!�Gbs
�+��/�j�Xa��W��*��X.��s�J	��>�΁J��r)�I���+O��y��-��=@�Ě�����;�z`%�3U�_c�տ�w���b�V<v�7<A�Nع�sG��'�~�6���/� 4�$5m�/[Bf9Q�"�SUBK�4�"�u�d�mT�$q��2�Q��=��3�=�}ٴ�u/B�6^���^b�У6��O���!�`?�5,���D�5����xZ���A���u�.y�D�=$���7o`"��
0���U"_��*bxY��]>���.H�\&��P�'X�P9��U�D=����{��gۅ�@��IFTw���2�v��I��d�K��!I���·�Ĥbǀs�Y�O��d���l9��3oh���2&�(�%����PJ�����D�P�g����%����ij��P���]#^5JC�ݠ,aO�����/L�%�.<���m/dm�R$  ��W)+���*3����Q���Q�^�o�^,�fQ����O��oy���V�$��J�sl����Z"�y��]P��^�Cnp:�V�]k@q��!�B4� ��E������c�Z���'Ư�1� ԛ����"$���24���0�b����s�����6i,3x�L��[l�A�hev٢5��^P���o��W'*ЗbӲ9rʑ��;DE���y2���V���K.r!cwZ���?��$5	A��&�7Z�޼61W�u�p��쾽�[	��yK�xO�ĸ�hZ�D[Sw�_�,�����
�_���&�$�j]�័�aڈ�c����d�Z��|ß�â�*��Y�C���eHIr�k�u0�>x8�8L��<[��냧~����b`�:�yG��w�x5E6N%�q�e�E�7(Q�s[��"�4�\hw�=s�!o2�3�N2�l�DzH�HF�U�7��`�L�F@��ȶ��}D�o��E��������0��/ͭD��T�@0�7�`d��/���H����)5��{%�IX��4�������F�e'*T�6��{�%A���X�@L��Ϳ�(��d�ҫ8�3S�6�;�u�����+��<'S�l�2F��j'��i��Ǝ�9�m�k� ob�����].���Xt�ìOM��푷��3�㩆3@&����td��!j�Wjw^	�-��ij�Rm�/�h���<����
�|�v����C�gѮ�5�`�]GvQ��S�
�,n		��ٛ��v����2G;q���29x�����;֋��ۣ� �4� ����y%��
�Hb��=bD�+�(�gBh��ﺌ�;�|<�������&e��2�'�2�� ��.6O3	��[I��a�Oa�Bh
^�����͎�_k�E����S���4�/QDQ���<<f�Qg��N��{c�fA���.!V�
��?���_�fl [�Y���,�1"�@���>��r:/��a�9��#�)b
�������4ڼ}KZ�Z���(�,o��Uz��9M�{��lS�7�P��@�<�9g;a������]RS��$R�%Iz	����/���a���ĕrT{$�ҟ��@AL��g����&��0��xX��Uk��9"~�H�)��� ��iJi��� �@����q��vO+L���f�V>�u�Ա1��ݢ��)���5��[(��6n����4�}�P��j$�& �Wr�ǻ��T����-`wU+�� 5��P `��3�ۜ*�v�h��19o��	R��6��h�6۟և7a�ۜ�'�a���!��ie5RG�T�X��fn��:�����ٻ��z?u�� �ܕo��A����2J���C�����}M5䚉�*|x�aɣ��B�����)�ӊ��2^r�5CJhf����{��rm5Z�b���	�dt)�ν�� ���FX:�([v��}�qX�����tC��J/ǥ�`�vK� y0B/v�V'p}U�e$nw���Q�$R���K�Ú�65�5кe�	���Y��	ҷb�����%Jv���	��+�틣4���7�,f^7�Cd�]����M�NZ��N}��҅<�#�g��",#k��83����n|7�u�:�oFW�3`�k�lf,�l ����7���˜�� �^SQ9R��*=5�%�6%�2�WB�N	n�hp9s�����T�d|�x��X9Vz&������.Q4(��<q4��b;$�A��tfbLؒ|���wZ�s)w�}f�{�t����j.6��%�=��MBOv�Y���'<����I�yE�14@u�ҡ�{�@MѸJ$}��~���)���68j+K�Dj꙲W����ѝ� gJ\*t���l�U1/`�$�#�t5AIq�2Ç�
�sH�s�b�����-jY=|s��]�"u3���)��84�c�[�t���ax*G��L��oAb���[�^�xL��@��jr�U~Gy�s{��[�T]l�xL*R�����t �3�7��\o󘾄�IerQ���y]�0Xn8�����\���6�d��9%s&����./,^�9�D,r��!�_y��t�w���.{9���1px�F�һ�@!��q`��_�~�*�w	0JA���̘��C�*)M�k����	��M�/w8�4�e����"�]��9әeXB�S������f,�z�W�{h������9����^����.�L���0��y���^�o�H�$@����7Ӆ�I����!	 �����$�=��N�r@������z�]Js��h�b����ۦ�BC�I����t@%L�b»�*s�$_�@���+�f�F����suX6�Uw՛�u��2(D�Bo���~�?��2���BEܻ��m1���(�a��xy�csاTtq?�;n��l��s�)�9����˿^�}���*�3�|��m���r\S�"E3Ҕb+�X�U�	�.ğSz;
>�ɭ�[B������]i���� }��a�#)<�M�u�����&�ݖ�M��(X$�i !i9>6���~��NlI �
W����3�.ڃ�!AV��%T�s����w��u��E<�Ryf������p���K�?7�����"�>z
^Lt��ar<Ԕ��
�����2\��F�4P@�P�告@�����҈N7��sZ��w�f�+A�x�g�^�����N�x�S�`��$U����E/YQX����BQ0K�D�P�����)��M���-Y���M����Im��_7�jE/�H���Q�J�������]�c�����/j������P�ЂDq��#��M�.�8Q��$����9�͂93#Vlx�h"�z:�1�ğ�p�T�'�z�wB;<�g+ Қz�G���H�L���D��H�^cՙ�#h��E�`a�מ�"�������i7��&�>�͢mU���{��ڡILÞ��|H�4N��o����?�{F��`P��[p����$W(� g�T�?+ee�&� ���7�,�%��;0�P��`ID���$R2�x@����P��