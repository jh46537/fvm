��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ� g�I��Jw=���c#hN�j(r��Ҹ�@���us���pDl�h#D�����|HB]�l?7v�]F!̔�E��#K�$��yW��K=��j�M��bv�H�b:q�	y��|��L�VaqC�`��H?L��\F��m|P�3�C��k'm�69��w���+���~��:�ȇ��Ki�s�|E+6�/�T;�#P��n���QS��<W2�)�4��UN8μ�럡ݰ<����㸛� $�r|/��Av˽���:��+V�tz&�0�!�"~z���6���e�w�+F���G�v�l��O�C�P������<����7YmGB"M�S�_��b�b��ɀ��ɴ��2�U�J�#D�Q�Sq��?ιS���*��nI���Xn��n��X��3��A��o	=��{���e��g������-I��>۱j(��LL:_��ڲ	
4o���������ܜ�h�n	��T'-O*6ք��8 s$	� �JB���	��u�V����q���9����cP"��~2���V3�nt#�n�Y[��!g~�R�ےE^���ޞS�\#��lq���[��p��r���$�E�׷�s��YD:��t�� ���1�����:f���mO�
�eJ�.l����	}s\c�v�c��EE,�S i� �yBE4ڞ[p�aChHT��vH��0B{i�.���_�s�;xw���h"����K�Y�m[0�/����*4�Z��Q:ʁP� p�J���Q��)��PϘ��R�cC US�gH����c�8<n:G�:�E� $�^4�-�"�at�P<)�:S+�Y��{s��I�sbx��N	~�%�4|����Xt��� -̊����C�}I�׉�� �~ŕw��˽9'־��R�6�;r���\����;��`s�X�Y��H�R��/��j4��^>���QL�1����|�]f�U��1L&�Ȕ����7�HC�6�6$�R�s�����;�k�*��Z��0�Jݖȧ|S:�C��QD�a�$��k�=������_��ވ��?���(zl�N�@���A����� }���m�Z�R������̈́�Ќ�ȭ��sD����>����",��Lp�[��􇎄��a���F#��У�Jhl�8FU���a��I
bJ��L�Mt�9V��m�	:u���`P6pz�d�^D�ȫ���M����R Bix�O~�m�LJ4/��t�u	t��鶷F�Lfk�TM#  J�蘠Kz� �KA���D$�k���M�veG�V��V��Ai_���:�^�٘U�r���Qa�hO��՗6^o�����p�K^5R�,����t�s��� ���p1/����a�0���I�!>.Jy��SY]�e��/65������>_H�Q��Q���dZ�ғ�X,~V�/�|����
]��L� !��~��%�W$�?� L:��0?_����qK�>#�W�{HF'C�Jh�=*U�]�!�+��|�4@�v�E��2��Sp�'"��Z��I=Q��ϟ���̇Ձ�?ȅ��*����fO�v�FNf���>�ν���ݑj����ބ�J����Ҁ�Gzv�KQ��8=�5���~&�%9u��2���ӟ�@�(37���64�@���y�G�s��O��H�Bw'�� ��������Mwm>����%u��L!�6B��؃g�b�ަ�0�#�/%�����BaB�=3�^64�Xc�g�P {^�-J�;��z�&�F�)�`�|�,h㴘ZskU֔1�i{��g6�/
bF �F��K�+�F��P���N�>%�@��;gq�7�(�q������A2��^ �u�٩��%���/�-�[x����b���\ʦ��M��\P{�]�{�|�՜��F)�)}96�9uB�݋ꝅ�3LT
�J/�?�alk��AT'�=M��w�/6Qc�|��4$K�L�9��`����N�16���.�rw���W�d�t����ga-��c�x6~ 7<���<$}A��k	n��_e��9�*���n&^h���1ڴ	�
�\�R"��� Y��qt�M���e�\D�z.(а4����B҆��✧�ԕsў�دty�b�����.b�|�X#�J�֜g'e�����)[��;6���^R���`��=��%૦�h�6�>��J�,)����qc��4�XZ�{
�8{�̯�������Tx�x���T��1�<b��<�^o�/���X��f�[7�Y���M��6�+d�B-[��V�}3�+{�����̫�ݯ��p[�`�>��>����NRۧ쟋����YXG�1]7.sr��)7���Č�A~r�˔Q18K'�0��S���O<���7S�ԙ�p�T���ZXz���4��aLxy�S��-~-u��5��(+��,#yM7t>����X֞.�����B���65xWh�w�)c�3��e��̒X�M`^�b��E"j}�������w�����9��+���s���T��c����Js����Ʊp0�ʒ��u �ny,���7��>U�x���QZ��Ą{�CHFx���� ��g�� �2��(6��2V-5�VT,<�f���a1�0����o΁Z	���n���/��3�4IYM����(D�d+�	�u����&���\�X�m���ǔH4�."��3��)����@v��B�̡��w��	躳�F�^G�΋ߑ��ۢk��<��"��&�ʏ��1��@[��6����'8�e,�r�};����B����}�(��lJ������Clm��� �!P[�3�Pf����<!���%qf��w�fP	�ݜ�"�6�]5�4)��]��cJG�̦�ʈ/�aݍ�j�JF�c�o��Dx@H�{v-rŐ�WN��j�?��ԏ��g�A8���֡r��6[��\��L2(�g�R#�07b�IE,��9Ȣ����T�c��w���\F���V�~E���J8���5@��-��3.5t��PGV]������J��3��)�|q��?0# �4��"�=����k�������шᖯ��E�h��uQe�b���ʥay����?�
4����%��[1�f
��)++u�mk�(�(�L����&k����k%��n�Iy-�J��J$�8����?� v�(>��~\���nI��)X����)���3�}\`݂��\|���m!�����O��v}ըP%��b6L�wm�C9�
R�ey�XGHt�?z�)��OY�%(�,^�^�EQ�-�L��B��~��Lt�n�Eoz���C͗p\(�>�:%r�]�C,�_>d�u�h{R��7Hl3?�W+����}��M�M���� }�^�B	w��ܡ�k����l�C�/�m�hoB.Tϥv�(��^��M�s\�� <�pj�F�pl�ii��$@p��	 =��	�nJ%���5� 3�Dʷ�%�C��w���-Gµ}ӰlV���껽�0�;n˄>�9�N\��uVW�_c�m�nv��?��,'�m�W6��5ĶeAGx�,V��vP$��d]��3N�ʭ`"���I>Њ=��(܃g��.T[��V��AU�����3�]�j�mV�L�*|�7R���/d>�'��8�!2��@�-B<�4>[�  	�e�����7Í����a��)p�4!ח���#�ͻ��i�,*9��I��xA���o�Wd�B��w6/eR�D�����PD�R� }fK��m�oܿ>_@�����Y	��{�(CK��2�������|�Z�^K,{��� �s�U�]_+'_��~	4)����)��@:�E����i�_��(>��)"�a`]2���u��h~��(M��đM�>�uW����"*+���	�R��hM�		3ć�8A�АtoD�9���l�vb$����N�mZ�2�����hȠQ�.~��� �p�\���*\���>�R��m8�%G����� �gnĦ�Nia�q�+����1����� 3ex�[
��Ro���
'�;�%O�����桁���R4 � �{��y�rVg�������=���N�c}�g�� ����������WHX̳I@e��H�E���a��l��]�< �6�<�%�͑Ll��i�V������fʁ���~,}��{��+�zŨ(ي�}f���>J8-К?��ݑ��"�K#�Vzp�3��k	!�$z6LM�j�y.�@BM��Q�
	Lw�,�5�����N�<h@k�� �=4P�-:?��n6���Y�xt�a��ZX(���_J�a���L���QK�r�*6��`6�@��$����j8��g�_�{�s��x`g�RZ�N��ˌ��|�.�N��K����_YCy}��Gr�I%OԔ8�ͩ=»ڑ}R{�X>6���d��(�������C��bg�kK��d߫7`�W=�H��ȗ%b�GZЁ����j���(��kĉ���l�4�&�~}�b�|�s.��2�%5]�nҚ��;Ī��Z�}�]�Z�Ӑ�N�a�/�l�}pIX���^�h�j�a�JO����[L�����is�?�WM��{.&��R���]�q�El��@9�JCx�H^	vL]�.{����u�U޴P~����qW��4ÜT.���:ζ��oL-h>�6��a���<R�ъ�����g�^�0c��� ��#�]�[ދ��BV���]���TmCb-n�|�Qc?���A����� tcuںH&J.��!���R�<�eq����r����)z�;9M��h��AL�G������񵵕ڈ�� ��ᡦ� D���4�{�GB6�r]�ۺΟ���<�O!=�����`p2i/�g���~� v�+���������w]#�Q�'�,����"��k�n����N���%f�1R���� aO �~� �o/�yL��r�,hb�7����k��� �\yz5߫Ч��ԣ�Oh44j�SG�vE��}��'����S��L;r�N�Ŋ���Eu��}��<���8��(ۭ�2�C���t�n)#�ӇCj��;W|���č�⩒b)�C�N��F��!��eڣ����ʶ�E���# ��7I�!���ZeßB��7���:Ny�H�5��[Z��E�p�?��,�2��>ɍ��?C7L�x��@a*k=Qe,�|t�����Ѐ�I�Iè?��5 @#D�N(�w�Ir����~�j�Pf�*>J�\��ݣ
f�`�����Ǝ���}?��3;������K,V��1Պ��$N�/.�K|� I�X�Vh�;c��M��LE�聯���5c� `(��a��ȉ�r�͋�$+�3���V���q�l�y%�b�3�d�.��@H�����{e�1v^F�F��^�wq�R]�f�����{Na�q��M�T��J]-����|�
{��p��Ş9���3��c&8,������c0@ѽש�&��q+��x涝����W=��~u��}cX�[8��@x���}h�Ѝ�� T����Bm,��2�K��PE���x� j��ZsE�MTv��YȦ%S�#��"�ǫU��b�H��H  �����G���Ճbk��S���,v�@�u���"����o5�/��q>Gז���QAHXo�p]*��,���Y�#���\��sv���%�+������[�$DϊlvW��@��6A�^�ʊR��ĀB�}�C�ܩ�Qky_����~��	�	�2��˾-U��|Nu�9aj8�-|�g�	:3��n��E����ϸSQ�����B9�XI�5�58�����8e�?+���s����3Mb��=\�i�{Q�8^˹��%4ơ@�t��e��31��	��y˴��MQ����J�EN��C����雐.Q?_�V��52�������h>d�}q�-W��Q���.��t���p:5X��r���c��h���^JK�������x�=
 *��.��Z��8-t�=w��J��B>��U��&��Y�f�l� K5{S�QH��'�-��Pw�#����X��:�s��O�}��0��;�*�/��9ڭlq9_|�)�,�n��wd�cGP�,����%"q6�z�<0��� #a�o/u����>���\%����c���ҹ�L=<����Ql�)�´�2*��&,K�u��0�Y���"3�;%��x}���Z��B��Z�L����Ty�iߓ"*7�v?��6�<q¢_#ć"b�2\��󮺲����;}6�2�kt��E.�Sv�M�E`��1�e5��bT�,]�C��n	�_���1��Y��:����O��2���qs;i���_)�>Q��C��I�����:�G�Ԩ������l�c
,��Mm��pp[�<�K^�`��K�:(Op�ړ�E{�Z��w�5
�cwB^�a�4�������ꠘdI",>b(zb��3��6`��3�GXI��IWϛ*�a��?�q�-���;K�0���ž��;�:��8��l��M�#H���v�p$Ù����R��������]{���-��e�s1���������&�V{i�k�����d��8M�[�T�@3�4B�]ޕ���:U�i�
	��,� 
���z#�M� ���R�K�|@�³$�.���vE(�\�������}.}xe�4�eN�#��C泶&Nxa��B�KڹrE>�7������>c�k�OW�j�]������r��K-�Ù�C���i����MZW�[X�M��+��5�;܇D �e���-�f+�/�c�:���Q�{���b+�)H�g0��ۀ&�������?~�~�OŸ����~0/�ͲqF8�.	$#�z�KXg!$]\^YV�Ť�K~���ח�jO9�/�\�4N�|�J���<K�e���Jj�־�^Vdb�̵�9A������w:�X�ݘ��L�焹Qۙ�����u+�V�ewU�8�(k*k���>�
y��~��X�u���x/F��>��I�{�E����%�+��<9b^��zh�u�x���㵱m$�ļO���dp�T�>O��0ç��[��J���m��G(�Į,�p�!vXe`u��}��or��*+��`M��s�GEW��I}e�g�+s��G.�J��M5�*�����S;7��Ͽ�;�q��
�}#��k�+(t�T��t��O�+�F�P��I�ϓ��R]a�e�;����?��G��V+X��a|̉怴��-������]; �M�\�z�vn��^�4��>��N��(EK+vd@-@�$�`k�3��tetoda�b0!�{����NdE���m�s ��U.$w���:�/�{ ���Y�ӻ{�q@P(- ف��vޚj�J���[Z���c������+G]�x�Ìy��;�E������b�N^ԺG�=�C)�T�Z�>�O�����D�z��pl�j�v=���p��) ���g��9@L_�-���>���c!��(`�C�)�_2�-��n]����kr���Z��/'�s�!���1~��w��J��.�CAp��i�	/���@�ږUg��
��;m�q�� �Q.�q]|�~�B[����i����2�F�Ns�7:��6(J�}�V{W�L��gm���N��6�T�u��f낱$��P����2˘�P��nI�� �G;"h����[˥���.��6��ď�$P0�T0ݫa��AݪP��Ӕ~�L��<`�h)�z�yO���ɭ�a?F�a7	a'�l��`�^�^~��L~��c$�oT��$�J���G��?�� ��8�)�)�VU�A}��s�#���0��Mɼ
(t���X���������\�BA�O�"f�{�)�Ho}m��s/t��[WQ���9�lb���DY3���:���NW7�.�^�C2�Qt�2�$���|ZC��YI��뭹�"������B�V\�գ6�4�@�|�� �7,K�L��~���<�����ض�-C��j�n��V|�����J���K�ƽ*�.�l��2���&t�C��$�ZV�AbiW��yJoP�)��U'Q��.m䇦R��ډ�w�q=�V�	"�0��O���Bt)�m�ׄo�wo�@O�����eX�(.�T���e�]P ��>�SM��!�3.l��p���+�Z!��#x�;���l�?�K�N�q��M�4P)����s�����L��1��ץjLg �P��ҙ׻%hif,w���&y[	�xv�A�����Uwf�U��ፒr�1�&60ܠ}Ѐv\��?�� �����ק	MI}$�gªe��.E�u��2��nY�|*U�����-:��R7�%������cӽѡ�g)�Rt��6~x/Fɪ��!�@���e3h�#�K��Nx(d� ӕT���.���2�Mve&�������D�^�,CҰ��(�ys�_��[��� tKc�D�g_�H��s��s�z��;��$����LJ�7rK�,�Xg��@Z�L� ��JV��/Gr*��:(@%;���(9s�)�uIJNў��b��?��V3��.�-������9�O�Z�|U����!=�yC+�����黎�7E2BOF�[��'@�v�,����^��]hk���y�_�`OgZ+g:\���s��#�R4�L;��91�f�L����)=��j�+Z�|�#�{��B�h��)�|w�aX�6F� ��j�"�4���M6��d��/��5���"[��1WV��R�f�������c[i-=e D��^eg��/������ʽ�=��u���w!1 pIcB��ڍ��84����������A#��2(���`@�Ϋ�F�zB1�+�'f���w9K1c�N)?^=a��������4��B�����H&B�	n��C7�ʌjGu|��=/���U�������(q������J�iZ��ᑮ��7ȭ�uth�_��|�1�+���5��V,fw�� �L,t�w�6AI�y��4.�v����o\���q��/��(=���ȟ�;��|-��x�Ja��1B�s���v��͵����hL����Mr��.l�v
%%Y`���C>=���D�l��L'���RҘ�NZ~�����H����u�j����~|ϗWP����V�$Q�}ם@M�4��hN\���dr�Ľы�1���l����z^�����&�m��F���1��)�Ox����1���u"�4U����b��R�n�a*��I���]}�|��qH�������s6�M>kv�������)�~���P�`�1����Խ)���(���4�����*Ns�9	%�2<UDR����+l=�HTߦ�:u�?�C���M&�_3�V+��q([���@�U&���r(0!?xY�aI-�a�?�q}���5��昖�`DF4j4R����G�X��w��
#�z�D8��6%�9�&�πW�ȚE�9�a�>�L�6s��G(���=�Z=������-��[�՛��Ck��c���i�}"�%$������I���q��Z�>��cÊ$��s�������� \iw�r6L��B����o�!�|�n��&#�^�9�d��,V�D3�ޘ���6�Ђ�Q߾zB��a'�kg�}R�tyF�w�˅ƙCk�̥I��B���ך}�C恵,�A���@|�!I�p:Qڶ�F,P�r�<�h�uKŗm< /�ޞ�֪�IS��<�^��yz�&[���_p/��,�%3tq�����{��[�۸K��~������G���<;xΦ��c�ϻ�u���5'<��d$���ǰ�m({����&�f$��Ax���Y���`.s1��o�.����9�X���j�uw����<�5>%�m||Z
Es��
��Pf�Pp>����̟?σc�)�;��Uezz��ڻ+�W��ɝ
�=d|cw���\��W�	m���6ٝn�L�K�j�������Z����#�l5��59{�����q�28t�ǥ^s�����f�[>*��:�T�L=������ԉY!�Jd�M��U��ӣ�R�9x���z�A�����\_���	�+'!z��~��!.i��3v
�-����İO�V����^T8�Ȝ��O
�Ud�A��%�e�p-H�Ra�iԫd���)�zk���ZCK{&o���;��[�D��}[ ����B���I���IS�$��м�O�����K��/�����X��XC�=�_�����$k��v��,�	s��i8��Ǵ+da\Cx���]��^��JfA�%�l'��Ny3g.���`K��.ZuC{-NKtÊ)L�����p��7�ҟ�#� ���V��,Rjh��Hr�����Ka�}Soo�I�����+�z�8"@O� �:�����\��*�4! ,���2�kw�q(�gH�[j�y�Ւ�UGY�Q<�d��i���� ���&���� �.��i2@�w/�\�B�W�b����[�>��19�L>7��p���b]�-j�Q>��l��*��/lqA$��Q��M�a�&�`�
Tht������/X&�8���	S�jA���Vu��M7i��(��5�lj�!�O$U��	��v�Y��1|�ʜ���R����U$����Ê�9�^@'ɲ�Z��ǳ0��U	m$�ھtF
�jcO������xX"���x�le^����)N7�}ذ����"�Q�_�RP��� d��!�b0�g�K-��b6�
�F���r��K!s�^pjPt6�|�I��}�TJ�n�b1�&�IK%�Cn�H����/1$��fͷ�����|y�p�����z����[Ԯm;�)�( ��q4M����%��^h�Z��:�T~Z�!�0��r<��p�~�X�)�$��D� yQg/|�X��d��,+U���${��6}�~����G���n�~9u�<HZ5�����{��=���:�$v�;֬v.~��6���Z�=U�:ڮe%'�(��^�,�湩X�?t�IEA�C����7�*T�`!}so�sBr�;�����)\�Sc	#6�-��?*����9��hST.y��!��*;�ƀ�g���V �e˛���Z,W�Dúj@�w�]���8����qPs�n��}�Ԫ��q�������������[	��� �0��Y4��_!tq63�#��r1czc�n