��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B����R����l�JxM%�$$���E`�����o)lh
6[#V&L�.2�%���1��(|6����"o���F�Q�,���-eQZ��m4�`�b(�I���w2�Λn�J�~������%@��~��� `aG<l~�tG&9��!���Щ� �;գc]���6`�AO鞱����r���D_?���0�����a/��3oE�p�:>�]������+��M�Q�'̌�����{	%�92�L�,ԋvm]�"3�F��Lr򱗼ݣ�65�R�?�}5Jj�%0Š������'�P$f~Ad
ң<Be�7Z��4U`oHj��3���܅K@��6��	����u��//���Z��ŉY�3�[37jV葝��;�[�˟h�ą�x-5��aDX�:�/�)���@F��+W�Z42a����G�>�mr��ʢ	k@C��j���Ww��v6��r��4����*�G7��� ��ap��eu���)�]MKw��� X�;�w��m=�7���;8R�2��� �a�T�:��x�1��Vk>�e�(9By��O�b�G����?�;-/$j���#�z	���:&��N'&�|�5X��Y����@ܛ�9�ޔ��{�^��#Z�&��ٲ|ow�lZY��%0o6w�@�u�ݡ6^ao�w5C�u.�K%����U)8VhZ���Q��K��C'`������(6Y?P@��|8��\B�����B9Q��d��Fy1���vi�*�|��Y��lH�VM�"J>]�ٚ����0PC>x�mJ�o ���8�XT�N����W�)V�g��R�-|�j�Qf��c�\7�j�{!����վ����AW�^��D�D��W�~=0�O��gg�˖q�p� ��#���!�Z�I�h�DvP�M�G�M����@��ǮV�� y���L�>g}��i]�7Zv�.A��d��]ŻV�.7���Zx��ܞaH%��=�Jy���M��HW44?�|��;w�8����9a���	�z��1H�(�'����a˶G��S��2n[ ��:�\���%��_ )&�������K�u�X{<f`���t-���T�tA�9�j����a}� ��/����r! �4�����_��Ͽk3;^0Y���HE� l�������e�$:�[}O妡<���d����0�4�ӯ�T��R�t�PD�| }�����[���6����
��i[^�3hjũӢ�uO�`϶��ȓZT8�&_��6%�#L��N��7H��M��ؾ ��sٯG�J��9g(8v��?����#�M����F,3�.g��bg���0���h��J	Z���K_#'�1���s��"d�t9������+�P�1a�I�+@�C���퍀�K���$H'��Ld�.�fl��Uw/�B�?#��G+�	�b��H��%�\�Ͻ�J����KRR������vrd��K^!$`ޟ��2��Nx���'}ޙ��6�b���;;�Bײ���)���Unm7\���	�M0(c�ف!�<��L3�wa+!ǀF���0�ϙV|�x��:7*u�5���/$7*C�@w-]�2p�n��Ʌ>�=�Kuܷ����U�'o6/6��mOȅ��ҩogd^j�*���>\�W��iN.;±�X�g�`���D&z��b��e"l}Y#Ɍ�a�{�t�g�[����հx�X¶�� ����:�	�ư��D@�Ii	Kls���bb��u5�e��AȔ˛�f2��&3K%'Z��t��˞,Ĭ����(׬�;���Q�s�m��A�s�ϽI����r[s6\�8Pm2��:p����D4:8�3^�=��ӣye�<�Îa"N�"�!�Ƨ���]��V@���ґ�:�7�9"�Q�Zh��(,o��Q�$��!��+ķ�P^�y垱�ՠ���	�b�(��y�]���q�;�{��EI�H��jpvP>}Z��*9�Θz�0�k�M�{����X�1t}�X7���̐���,*{�\D� /�������`!�K�c[�][�3>Z����T ��5glp�����ִ�C?��
�W?�o�b_r{��ƪw~%���d��UgK��a�W���	�p7Nb�ٝC:�(˝lˤ�u�`bŘ��
1�r�AU�nUD�r�eH�ą�Y���6�jqO�����[�����
���J�[;�@?2��������͞m���D/�0~4۬}�>��1�jT��ʰ,fna4�%^��"��%_ie�~?��S���бN�*R/��wL��Iቢ��6�.	����ہ0�����ù(�&��8��!nn��0fGjU����o4�p��"�4�&�7Y�E�ϸӓ{�V�'y �ڜ>sۀa3B��l���0h�J�Do�׊Yz����%���m��t����B�ksX@��r���N�A����'�=?\�T4���|���yc�s��{�P��{�_���GoSg����A�j�i��w�y�<������kx����ėʖ�YH���֊8¨�J�f� lG_6�e����W
��*0��6�*�}!v&���tߡ��� }� �ET��hx*��Y;�\���dY6;$��i�����&�~D+Nah4�a���7»j>ʱ����Hc?A�#��,H+�&�Eś�#th����8��ӬB5���IN�Xu�5�4�/{Yx�6��>zs�J�^�A_��>ʚ$ń��(GR����d�sk���8������'��î�Q�d�'d�5������i���˓��YdSs"-Ч`�K���J���]�G�C3�;�d�I�y�Bj/ah�m�Cp�18��ۚ�)W�%�1����(�"�ߺ���yp>��
�>C�-n�o�v��|x*d���`��g1�?��/�I�� B�h��f@tŜ:\���8�*�E�j��F�:IlH��D*v� \�g�5�B�=�'�����Bh(hA�+���|�|Xϯ�m��^����Oa�_طy&�ݓ�쩪���Y��n��O�<��L���% |4|W��B�b!;������ˊ΋P{�]@Mռ���*+�����
�R]/��WzA�7��6{����m�`��g�V��[I��u�᰺R��8�%y�k��ۧ�TR��Hb�.|c&�l�z6̾�����ua�{U��RO�(r�Ǚ�I�)�ߖFF�2�v��SzP\6�L����I���a�E������}�4�3%]B�qt�?�bA%SJ�yۥ�,F��dR�pO{�'%a!1U[��R�䟓���:���y����x�#R4�hFŻ(.�8#��{�`�����(���-����n�GH��ڙo57�"���e�=*�$'K�U�ʐa�d���C�2�Cn�r�gD���WռC��6�&�1�ճ��U�� ����c>��B�6�=r�C���e����|<�ܢ�8b�N���*���D�AMo��c����0r��b D��.�j�TϺ�?���~'(`�zް���bע* 5�ǂ��R���N�K߇��4��!8ʘ&�{?^��&@�]���wd]{6w5�ű软ՉA����'����W��y��5�z�B��$t��m�P�ۊ�8����/h���}���XK�u�P����7e�����g�6��c�k��LP
ii )�.a3ԉ�Rs�{����m�&����1��[4~�v�����`�W6��00���������y�������k,�K��V��5�irs���C3r��k�bg\϶3&(�H��֣y'1���s�K{��;&ה�'[�"E"�f
˟��6U��i.�p(�H�Y �²�/tK�\�k|ղ��������q�\;΅~�����/r�8,���}��վ��ɹO���������Q����]2$�H�{����Fⶮ	P彻�;���^��#��^���_��Bӆi��u��F��$��"��F�WlhƊ�,Z��#��n[��w�X����:ğ�Q5q��g��0���~u0G��b��N�f���.�*%���hO�03��ԙ��؆:���G�B�:�#ɸ�4� F̕`��
���7�q�XN���+�L�np�0"yf��b�U��)�waT �����	?M�n��FY:�('�@�]�j������pJLBm���ޜV�A�l��)V5� (��_�3� �0������e�V)I��6��3� �ڮ�����	F� �@�K�K�{�Lr�b%�7/�)���,�f�������\���.\�gE�<���]-����!�o���J���z�d]Ivu7����3��I�_���o�b�\�=����t0��/uR��-2u�X�,�����!����~B��K5��<6L�=y��Y&z8"�!�c��ˤ����!N#lVY���[���
����f�L7����7sԔd� \�6=���>��M/�5>������m��7
�\o�p]�~]�d��5@��,KJ��:�]�kl����^��e���"V!���}p�32��`��������CV�$�����o��`���������{���5�� ]��Z�#u�t6l�r�CQ� k��lx�co��$E͞��X ����pd ���ܺ��Ve��^?mv+�H�����%1i����/�r�(w���>���Ȅ� _��6O������	',炨���0ɮ���%�ww� =P��i�\y�[ag�N�dQ�3�x?�h�f��Ⱦ�̖/��?+*�i_�pl�Sێ��X�V#3B&���{�	�Z�v�є��3��U��Z'%z"���VMW����E�Sѐ�or�lr�4��WDZ䈢08�p-3����H�[����;��t�榶���+C]��٩��>��.����-��C|)�L+��j�/Ju���P������p���ߊ�O���,�FJۋ���1:��aS�H$���ED�L[sõ�û�W2�2/	Ȁ}^V1�{��k݉�� ������(9���`w�}��tq~yڅ�Šn�SG�#��J
�w�]�(�%�&Kp�?��ix7�D�w�~��w'9V.�;E#���W����l�	�^�x���I�Pt/Ll3`����b�J���M.d.S#�!��펐��0�T��Mt���q�u�I��4�n��qc�;#Ǐ@�K1�%U��Ѷ�ϵ����0w8�!a����;P,*"Մ�߻^G��rC�U�NO�`�U�-�R����D|?��޴*��߼;r�>�Q�V��_���XK�5�%0���>�nNtB'�v�I�
��i�5�%�wr�٥H���tvz�Q��;#����u�m+�ژB��+�N�M�p�f�d�=4y|��kĜ���P} ,hH0°"��A�q���)�	���ĺp9��%����.]����M����!��]|���q�^;r��w$ Z�� (2�w�2�O��Jh9QN���)�8�-S`u�Ҥe�=K�9�$�@���:&f`\I{g�1u�H���`C�p �t5|kJ�խJ;y�hO��pc�q%=�$=
�����Y����5l-�
!1�F,��(��󝽉p�����;����u�UG#@�+��Q��$�z&7#�O��ȆoK�/�NT�w�9�S�((�[a<�Aݗ^�!zE`�UD�q�2�Ȥ�e:���ۄ�^C�na]���E�g�&4+O*t���Ώ�rG����)�����W�&էt�Α���k�����'��ec�����]�_K��������̟	'l􏾁�]h�qD�@�j>)�2\��:��	�pN�`g�[Y�:|��;��e�^�U7����HOQP.�FWCLJ��#�K[{�Ͽ\���zas�8��bVٸe�p�}���	I��b>��u���/�̗�����زf�t��&v���E�%S�zfyNW�ezB�:A}���.�ETqW��tO��OB=y�����j������>�����D�ʬ�(c�*����!���%.���(Q�\)�{^� ���y�{=��F*]�ք�m��E
�!��2�I�^v�`�)��>�c�~����ᅾKL��<8����Iׯ�!��g��Kؿ����o���8��P��Gr�M*�|�� enB
�s\��13S$E.ĺ:��>������<q0%���|VV/j��եma�rh�%k<Y��=7�-�Fa�a�~=�����&�m!Է��H.��7=1b� ~�h;����V��nx�&�i'�	�ٲ���wUM�:Ը��9Q�;���������m��l5-���a*.�U��(�X�܊�W�,n>�w"�<��@_�b����]#ͬO�g�ޢE�'2��WW�c��|��6�~@ZPc�U��_��dJ-B�PP��ƳA�>~H<Nzb!sy �4>�e�PVvݛ������H�H���Y!C�y�x�Ȅ�:�n4�����eU�D%�hY�Ã[���>���6[{�����1�|�ձ<>Z��Մ����`��ݙ���axh�E����H��s�;���?ڜ}#��p����OEZ!e�Ʀ1.�����y�������T@[�� �߱��U�`ݽ�7� ����
����O���!x���
�4ʀ��9�<[(U��z\(�m�n�V�Mi�c����B⶞���`v3��D�	o瓚'�qd�º��-Aݞ)%'�1]�~wآ�G���4J����F��T��1]�Z�9]۵q����J����s:��d�8�j8�����,n=|H�W��J�GycTb8d���k˖�KG�s�cY�u��%=����U�j�	7����	D2�?#Fs�bFB���qo���=�\q�JB��Y'�2j�;��4���R�Mb~Y�4���-�˝�;n�RX@_�f���s7ׂ�
���^J���I`�n�"m�3��H7��?�9�Àn��2̘0AǾ�,��~6�}3Q<W?j�/���Ci�y���݄`��+
�]�i��!�]��_�������>*rzH6�A8�m���(#+��L���-O�6LZ��6�� �T8�N G�����<���m���n�%8���K��){ ��o�uw��Ш�t^����	�
v��ޓ\��n"�d �����]�?�~7���b]Vo�Pe]|�>�6	� �W�m��CR���']쨺�	Z|+G�tf��$}-��"���DH�<���1�h4(k+������d��j�Z��r8���<�b�j쩉ڑ ���g�9
b)� P�U�w+�g|&�{;_�D;ڕ�7mTyU����Xu��X�U���MF����rG��|HQ=��������G�;����E<v
��a^�J��_��`dO1``����������{h��Z$p	~ҭK�ʏ�����0�js�������&�=���J1�)("���7�fj�ϟ�S�!�+�4�7�>��������]qs o1���n3�ξ@�q����� �|��9�,IT�O~�;�׺i��k��i���
ز���T��b��r��!U_�N�`(��DʣWܮ�<c�շ��*ca>$Ey��*�Cf�tO�2�N6\F�q.b@�N���=��3G��(��l�����