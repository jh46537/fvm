��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2Ȫu��Z���d�]�$\�h�����oր��ʖR
hgO���m��i�Z�O�L	��M��a�ok��Q��r�Է��z��1�� ��I�-[�?T�oNmMǮ�y�B�ˋWC!�}�O�C8wְ�Df����)U#�� �o\�Ғ�Y�b�n5�{#G ��k�O�e�X,j���Aϵ�\i�h�nMOŬ>�&�j)l��"�#'�[X��^�Yh�aH+�����oJ�	�ge� ��G�9���it��}K8�+sm�;��&��=B�V?�������z[�`?�WZCc&���:�C�^��t�6%(�5��LT�ק���;���=r�c�,뀱?Svx]{�����18�Y�Č������H��8/#[I�`�nm\�Ɉ�2�1[��) !���֘Gk��%.�t|�)#F�\�B"䡯\���Α�Z���n�+r�C�'��3{�x�ɢ>؄�P<��[�]z8��+��t.d��<�ջ���P8u���R"OYX��8}e��$��<��V�2T}�߱C���G�S��V��:�8��i_jB+��;��������HΛUI#�)�@���U���qJ��Ԭ=M,�C	K�?�%��R�'�K��;mT�� u�n�/D =���x0��3q�ʴ3��rq����y;FRt��� ��
�ܻ�K�><�h'��X�p )?�K,�_��wwm1����(LE~"��')ۓq&/)g=���s��-I�������bq��;$Ap�����dʨ�㑒6�F.DQ��V0�6��&j��D��>�}bo�L�0�ʏZm�C�	���ύ��~�X�5Q����7�{�KD�������D*����d�+�R��_�]9�a�C}!=��~%+[C�4�Pua*9�����O�=�}e^�*�dLe��R�h�_�e���6|�.I��m��s�귋��D�8�ێ|^�5�B�蔪L���8�I���0 ���ȱ�b�辊��o?xC����qp��EA�RZ�#Z�R;z������A���D�_	x���w�G���0��B`M��kM�)�|'���whR��,	ȷ��B��B� �o���m�P���h�aۻ}�#��Ȍ2��/9A��Qw '����ʣys����$���Hp���NN������k�	�n�vQ�%=�yc���8��AT����DF��X��Cv#��m�NzqvVm޶jMEmj:1PBԘ�f+C5VG��H������cr��L�YZ#��0^}V	�!��ͮ����AT�\�D�fz��20����r�����	;��m�]Ҽ%��:���ʩ�}�qEA.,l���T�UW���..,��i��{E��ߡ�!�y*�tr�8��J�i��ɣ�.`){����&s)���\�S�Q~���=�s�Z:������vj|SDd�n&�'�U��^'�AJO����njRU�I�Q��iV���0�7SaĐ�x�?�tx�#U��@?E�ԋm���!�Ȕd�&��&S,ps��p^��-"K��μ2��4Dg�-��y��αۑ;*�x��е��`m��i=�,���=ʨv�A�bD��]����?��oW�Y�� �q^ϙQ��'����{����^��$ó���5�<���0�":����{��F��@P���M{̏���[��w�6KϮ�������%o/��F�7te���hً9��k�?�vf���|��;�:0�Ӄ�T����Xں�2N[�D
��|���q�EB+ԩu91�Z��:��d�Y��&��`v�9>���:}������.B�(�$��Yh+В	X��k9�#S��y��¥�"�	��s돮����|)�����< �k��9qw�&<��eeu,#Oȑ���Ks��f�j�(�� ���V��mu�F�U��Uu��:�[�7;1f[R�%-:m">�,<c���#puJt�l�m��<Gugs�i�YlMd�[�5\�MN�@�uj϶W3l�b�rc�EP��m��(]���p/Z�߆G+e,�O ���3Bn����X�WbH�B���b�[���2Fu�V�8?Y��S��!�
8Ј�΃t��o%��^�e�6�F��<Mg�v]Ôr.�F�9M�0�gv���i�Ld��S��͂[ ���5/���7�Fޔ�-�9
�GB���B�iI�"`�g�7 ��31<��d�zƛ��w^c��i�'H��9ό������0�"z�%�`�����O��H��t{x��[�����Q��.�����5`e�����j�s��`c�@�J����mM(�o�GסBB��f]��^ӽ��
���dI�����C�k��9��:�&2�^u�����ZA�.�FKoT���_�?��/��]h~_��)��y�ɪv����{�mY@;�:��	��<�#'��B�x�'eU���7��p̔�*b����������mg������wrЫBԺ�M�ZAư�uWq���.jQ��O*��y[C,:n�L!�����q{��l,���On5h�ٽˋ,�U�9]gy�����_��qr�Jy�Q˱�h@lAx�� ��G�ø�w�
ɡŪU�J�KŽ��3Ť���In�K�+��b2k �@*��fkdn�.U5��Y,)�Uh��5J�L$���s_f���Զkȅ3%����b`=��3Q�2��W��S'�8(��)�q-�J+}���fi�*2�?j&�uR�Q�,0׆����3����~���i]GkF�V��5e��o�f�B�|�>L �p{���Y6k�����I����n�I1~��� ���I���=f,�y;L�`@c�Ye8ݼ�5�m�_髆���8�3-&��|�f�[�رH���U�P����A��L�O�TI%:��8��l �-� cE��¤<U�%�)�DPl�^����d���Bwlyӈ�u�r)B�sv��$�v�B�ަ�Z|riF����.���0�J�tY�.���_�m�=�2/�ka��XߊQM ��Un���sG �@.�F�Ө���S�^�Kn_���ឤ�u�za��tjJ�ck��n��Z�o-��7���Y�?"���e'�ӫ��y�d�ď8�G���y��	�[�Q�]�f�j1}F��^.����x�\
�f]�G���V��U�p�[�{�q�������6v[��W�_z���{��A��D�o#�d����M5�E���S�����^@HijU�j4K��m�<7��e�i�C)��������!�*�Ϭ3��"��g���I	й&��Կȝ�:^�y�H.�]�B�T0�d��� �Hd��C͌N�[�} ��"ͯ�N��N�.�ӥ�������R;!K����8X#m44l� U��zE�����iC��޷�[/�2U���m^]=}ɾ�LĚK��@wI�j9�G�]��٠�'d(��\�v�nȐ`�<@s��a���$�,����_�L��3s���-<�Q,UgaxI=�RW�$=)���r��+�
���iqb�$����E;} �m�Z�'s2s������b��r���۽�nV!����x�I�,LY� ���5�.���4�Na��a+O��\�TI^���Df!0�W��@Q�
ER�Lf�
p��K+�*����C�{�7��?��
S�ܓ؆)P�	���g[,H0����2�K���t����g�͓.�C��%���K��w�W<�Or�Z;	��r�J�X��̭�Jf!߼�jC���i��7�^��:�=j[>Bo�e���GGVn�h2c�nM�����aֳ�����ͯ�A�V�S��HB�Ҽ=�e��С�g�(Gi�fjC{/;�?.73wd�U��s�! #	V����Я��Jl*W���3�I�QO��i�K��휨@e4����0�����a-h �3��� �U*,���:�~C�4�h�\f_�&ix��M������\�u�t-y��V��DB����"+	!�|X˕��#l=}�L⋍�Apɹvͭ�&�K��m�JMN���|��Y7:��� G�(�D3�������%nz�'���Ճ�� ��|�� ��!����mq䘂ģ�����E-�l*����p�å ��e*��K����������p#m�㺇����1�つU�["��H,��M��� PgRY�O�Mdvi��{�+l$������\��Ha�B#�p���t�\��q�\s�;s?J焐U������;\n��r4�X��׀RӚ��A�[�D�C��T�^���#���NE�i�N������+/��*��2u�H/�3$I�;��-mv��D�N�/��m��@��t/-��K ř��+�����˃1�"D��=�=���7�	���{ϡI�=�ό&�*ߖ6:�j�_�Z�Hm*��U'&��#p*�Q{��	ǻe�o�!��	��0y��s��I�:^z|P�G�NN��G�6����	�ڇ��f/��_��Ae���u���ӫ�Zl��}�ay�4�>�L}-�;Ìm�KI�7�z:u��Nw�P�\�e4I������h]@�ߖ.���P����^�5�7�X!��`��n3f�@ٴ�M/��8C\����P�!BB�������Y��I��,�O|Q�#�"&������C��;���¦��'X)�1,]?���|��£��0�{��������	�`���Q���H&��`^h��Qw�3��k����}k��*l���S��ISZf+�4N|@3l�m�Pg����6������JY*��1����c}9��h��A��J�f'�<Y�{p����ɮ�N��n�T�A���P�R%_�W���+I�uq���H�,��B�Xa�F�pI�G��,ˬ`��Ԇ� .eIR�뚅q5	���K��Lݯf��ƅ��d�Xʀp���r������a��/�`v�pm����lES�렸"�����7+�Lc��o�{ٿ�7��y�0�y�d,�o37Y���)�G;"!jcsc:u[3��ӵ��8$l�L냏b��)�g��Z��㱈����m��N�.��R��۪JF � �V��Ku=�������b�kV0�'�WP���0�k�������"k�3gx)U�*�4=�F4g�I���^~m� ���Ձ��<�g��3@��.�ϽE���(w��
�|MDD���W�c:G
��im����_�*.R-��+j2(�!/�.�O��p��_����?���|4�B<����i{]� E��a�S���Ƒi���Rw!�������HQ/yf�f�P����CN]
���&�qћ�-�}}�p�t���@�X��s8���fO��F�4��D	� ����!o\�Hy|�1�z������2������.��m7��z�����a��e����q/�7PIy���`��W��nw�7���x�	4�-���!��j��vZi�cSxE�L[�U���_.�#R�wն���P��T'k���?q`��<�q��<�yɨ�]�q7�5+?���OSQ�'��2�.S��2GP�,*CMZ$ɯ���4t�lp0|�ڵ�sYWʍʷ���gW3C��E�e�z?�<�Ou�d��ٓ�7�x��W��m.�˭