��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B�6ƨ��J���t�&��a0��8�ڪ�!r�FEX���K�������rs/��/��E	��"6����z(qN���;1�q��M��<�S��{ �8L�F�˞ ܦ,��h7G�C��i�nܒ�ġQAɡ|@���L\\�E�T��z�:�BD�W�t��O�㋸�����NS�2�x�!s���� ���a�.���A��R�E��w䢀h��z97�2�'�S1���C��a��G��Qu,����#ѕ��_�Ol�w�+�_,-]�A�_U8�'��$%�2����?А�ʿ��$#�5�X۴���b�"�d�l�{�������Ĺ��Q*�R;.�qKvZM^���b4����Pd�~�jF)N�WxeK�Rp*E/ވzȺ֒��TW�%�
� �k���˜ef���H f��n=ɳbW�W�4���7��N<�^h��[�j��=���3�A-Ӝ�L	�/�{�	3�ë��n�[�F�#B�~)2w#z�ћ3����	z�������K7���#��X�t��D9[��X������B���*{��E�oK�L�ZT�t�<�߹)���7�?�QJCa�a�q����a��IWb��c	+�UwRꮭ@b?n-��5\UC��J*�,����OFQr�R`�	���"�!�*RA"n	?8Z$8ws�8#X�:������r֙�[CMap�r�>��.}�N�氖����UY�؝��#�8��Υ"�&�Adl;?"`6��y�7N)?���:%g�ֹ���L�w�ch;]]���u:�C��G��R��B�l�K^mM)\t�in�e$�0>RW���g�N9ya�w$d�e�əqdt?�W��S(�`�����B����BGi�c��
��FzR��1'X��G����-��4�s\���&Ye�Z���N|� l��Q���������bp�A+]�z[�:� 2EAܥ�?��	�-w
�#Y��=�P�с��5�)�ᓒҧ��Ϊs(ƄO{���*@fXso�k]���ϧ�U쨽����:��ω���g܌5Z�Up7��<(�ޞM������I4�`�`�ɩ#Li6�3��'iH�,p����@o��[���-�h��;5���)U��V�8�c���f�'���>��3��t���䪠�e)�B�/�؄����r<�g��o�`�����4B���om+G��}g�����z��(�I˙�|-�����#S $�`K�,s�W����Q���<&_�����:��~J��f�c��Vv�9C�X����寅35�n��P�����̜�yJ���|�h#���Ӝ�CT&�a1~�B:?�گ�L��Z� �~]��4+m���;�hl��{�8D�Z���g�J��~�z��r���y}Qg$T��hq���"�3��n�&{"�.�'
3E�c��n�x =i��3NX;}�t���� �7����P�e>��}����g~6�!p�7��|�	�Z�a��0!e!�s�Am�9�K~��	��?m����yC ��wI��\�S�9�C�w����v�F��*�g����#�+9�v��s7�X{�CYg��x�]��ǬM?^-������� ��N��2T�����;p���,yy�I���L.Q���0k�{��#��2$\2�kcm3��H���uŗ -g^�Gno����'��Iz̻�ǵmH|���b����7���T�lf�~���g�F:C��d��R��ҭ�S|��?�)ٿ"��Ӱݒ�5H����o�93�?G��Jk���� �W���6�xx��,&��޼U��Y�P�n}L��o;����.L�M�	*D���z]���Q5# ?A�3 *臥�~lY@��r����/�w��c.�����Â=��g���+@0׻}�ߦ�Kv���gdzq�pW�t i�?���7�9��z.H���Qb�k���g=���{|�&��Yr����R����|�w%M��U�|��B	Cs�.����?�厈�z�r�h;��c�3i��묍������*�f��m�bO��@�\��ݵ31�H?E�L�Yw��H*%�F��1�jju�*���X\�\#�ge~�;����-{ߔ6u�/��xM��xV*��^�Fg��i��q�(��v��4y��^%L~�uƱ����A0���T�Ϻ2�r1�H-��<�1�>-�3G�);>>7�ar��QN�H>�5̞��ݥ
� ���k�p�r>�M�fP��`�ӷC�˸Iv�}M�������W���:�_�d�8�Хaa����1���A�>�-����*�D*�N|�_��[���`k�w��6;Pi˝�����c��Qg�]�,Q&ăO��v->A��PJ�?48���?�[~��2^!��v�	ش��� 1��>V��u[�+��3���A��z�+�`Y��\o�/�2�-[؃=?����JQ��<3�H����1K�ny�@_�݊����F4��G"p���ˉ���Z��h�${3�Y2������S��]��-�	/t��y���n���Tث��U��a���^HqP��.�RȌ�8�`��d���ٱ��j3��HUFjI�5#��,�����5g���BW2I*:��j�)�'wB��f���r�J��b��\/�[d���y�h���T�ǇhMŲf4,OI#*�7�7�w�jC�<ʺ� v�C��pX�(q�B��ҥ�+���H��l����7+@ 7^6�T�q�[HU��ݼ�����ޝ��j�����)y��x�����W���0�U�/�s"f�	&yK%9K�Q�RS+7
/�%a�k�ٮ�%H�A��O��δ,.aI;�7��Z�7�:Q���VOa���X��?��J�J� �p�P�ki|�8����ƗZ��p[[x筩Jt���g�(3����Ꮰ�a�w�F�Z�w�݇-CT;.~���>u`S�H�vr����A��f�51�6���o�s���"�B'Oz�%k�l�'��5���&�5i �N#Q^�����' ��~fr<��K�.:I�t�(�.	��]ѽ��+�oɐ�)�&�]� ��y�9����ef=u��O��|���/ R��'�Q��GK�5�hs�-�f�Rt���kA.7Bs;&�=�u��_G�]<��T�T/�\���_�� ����՝G�]��'�d:d��zs�L���x�����E~����t���p�Vd:�i�}����x�d�kz�b.1�D}�HB0�y%_o�B5w%HW7jh��][z%r�)H��H%���T΋�p77�l�M�>��2�����L\(�I$	����U(�C�C'Ǟ���[�_���i6���؞ݵPa.4|�|��K�Z,l�2������@��H�B��Ə��Ty�j͘+��ȣ�(����+�p?��~'���*�x�[Q�������*����!�-|N���V�(�8��E����v�f�4�@/���wEz/�_��	a�QC��M�o��������/�N�e�c����냌�F� A�����J$$d��Y�h���1�����ДU�?�;Y��f��m��!n5;G[��X�V��	X�i��wͅ�N��:0DՌ�	{����U��f˳	a���hv���9V�I/�P�5I����\E�yM��%J=���m���&�i��)Mx��<\V(�����"fiv�!y�����h����^uC5I�߹<q�W�|��W�䴥Oncdݑ�Q����H���g��YG�9�X`�0�]5Pk�
[�<�L5�蠂�Ɔ���C:﵏D>v�,���h�j6=O0:�dq�]h�|�y����2&t翏���D!4lM �lVJ ^� �
lf-����.��U���ֲ$Lb�J�����x95h��T=�7���*�|2;�ǥ��1�͛ҵ�k\1�ݮ_��߶\���1pgfd����¬^����ӶlAk�,���ߚ�2B�S��BGAB�[N(5O�G��z��}󑠭934��Y}�j&�@�wm9�EzEy�2B�r���v���s��(�j�O2w�L�t+��$Ma�hf9�7���U�L�O���^�)��L��ȣR�0����g,7��zr9&�_�odt�8;�Mf�cc}�g38�`�'�h�B�'P+r,�me���h��zZ3����Y�8�Fi�2!�/6�̨�|	�2f=�+T��>
<&�1o�f֣�Ց��D4-��u:�H%'#�]�
�Zv��?wXEf���ͥ��G�Ffz��1�Jyh�o��O�#����(ˣ��^�@��hd�?�fu���Ԡ�q�v�䯡�:� �C:&N�a���	vʄ���؟�Ͷ��T0�0�1J�TVK�	���E�T ӣC����2E��;`�A�Ҷ�����qw;ɽ����d�T�:�%��ɤ�G�Ѧ�g�:G�j�
�C��*<ʭ3�T��$p�#���"K?�^���">}
�;�[���5�p+��s�:����(%�t�n�T��=�}��ɮ�Ӥ�- !o�5�����Կ*���H?���I��b�z|��+
�0�EvW��&����LƱ匈L��?����{1���/H
ad^do�q�H��Z)�
 Z�b��44'��5�Nkj��b��h:A����6J�赶@]��m��~4j���S�ì�F�A+�J��$�|�����,xq�����x�4#)؆lv�W��3Wae`[T^v*F�qD��`���@j�Q��PzDcA1��= u���	Oi=Z(�&�;��Ba_u3G�Oq���vs79�cfH5�oǅ���_ћ�˰0U �9S�& �GS�����fR�p��y�==!>��֍dGٿˆ�6i|��	r���
��$,;��i�-q�V {�߻�M}f7D�_�*��h̟ӛ�bSJ9%��ptx.:�>���7iη�X�}��?#DQ�1ϫ�K:)5A���ާs �ު?�\Z��׷�h��_A_�}!h�#>IM��e�N8MF���V����k����_ *��������Av�䗉�6�\�'7
 �ʕ�X#�K�L�,N'r��ٯ?����b�1X�_�
��r_y_E\������+�	x����=��p�Hs����˱��u��7����]�],�D�O�\ֲ�?~ǵ�'��Vb�͞
���7XB�\������7\��QA�7b�'�O|���K;�:{t�S�S���=#~p�į/���11Q���l9j
-��H&X�-���o�L��xR3���x���Lx�r1�Լ�����	  B�? ��[ݍ��/Q=��i���ȅmd�o5����T���^*���ǐ����K�˰y�NU�pԔf�����jz���Tݬ�ߝ~Va�a�b*�;ʯ]N��L��e���ח;�C*?� 5���&"���eܹa���?\��ҶS�F���'P�u#�E��
� ��0��bݍ�*�*�O(��K�e@����U>>s�aY�Ʀ�u^�'�}��7&ܕ���ݖ�L17�P8���혢��D��~�ْ�cx�̻���*�������.c�A:�F�c��a�z�𞩓�����*��{�L����=������9��d���f1�˱�W� ;+-t�� X��ت�p�y/�QC5�2��;N1B����ItB��V�����l{�0[jDh�6űl�H��dyq*7A|$�is;=�~|�*�vE
T�=ǡ���O���'OY�E\ȁ���Q\B��d�g���o�@��Դ&�7�ѿ�(-|��{��7
"L���/G���<�oݰ:��ֲ��۴܇�{~\H;Y���܈42|u<E�Ag�)ȶ|�餣���O�ޝZ]6�t�+��yL���M*�	0�tȖ���
H|�s&�bn.�9C�7���ʕ_�!_�s�2ud�ϫJG�������}����O��.������@#��&@��ָ���6�3��F�,D;W��t�|�1w������B�k�8݆�y���y��H���X%�^��x��!§T�C��[ ���3�P�^h�BDl��`|�.�#@�θ.��:jk{��,��K�L�3D�c��δ����m\�ë{�yБ<Տ�<�2