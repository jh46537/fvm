��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���a�%�sK��h���/a�y���v��=��w�����:�y$f�*,�RA\��S����ћW;�U���T�Ǔ�q�0`�eѓ^����8YU?to�Pb�I�����9���������:����l	�~�Y���)���L8�|m[P��Z�ј�79Ӄ���e<���_�����^�2�����
v��;�{a�<Vx3�-�����ٍ��/�[�mg������o2����@�m�e�?ኂ��l:g(Ozl8S
�-�CW�gF�5�դ����>��'K�:���ϵA��8�l��X�0S����b&�7�%)����!�h/Sq�㾴.��"��w[�Xe2�.ƿm�?�g0ۉ.�*9D��>[ˬ�?]#��m�g+��;��Lb�W%��"�����n�F�`��VW��th��Y*�1 ��a�|�!D�+�iN��	��O�!��x-�'b��Xt�+�t2��&���Q�Sn'aP��������p���5v#�Gf�\O��7�3��}���_�!��5v�����$���Os��8���+�o���7MJ� �&A�H>{w~��H�?�N�Qȑ-e�U�&u'|��9o�j�
s�/��>�`�5��5p����IG#���Ę��d���ܺ���k��g-�Tn���\��w:�oB�g&� ;d��/^;�/�9�_�S�a��u�fĖ_V-
������:���r6�01J�s[�n���p�����y��&�� O��ы��y8�hT	UfȆ'�T����v�5��!!�&�F&�Q���y��ZM:�f��m�]��d�4IVx|�q��Q�Ғ��N4ɦ��d���	�VW��O���P/#i�hJ>�����)FN@�ҡ��.�!�u�L�z�eSF�!��b!�`5H
`1듐�=^�d[�z���)���.e�0���U̯��y��M�b����6��v��C%����#2J�s�Q̿�A_������r�o����X�ĭl:��!����a��� ��1��O~�iM���� kbb�E}���s���c����[l�b�yw�v&�s�L��g`�Zbmy��e�~J��> b��<�žx���Z��>5��'��k	ӖN�z�<S�$�+%B4����yR���{oY���D$E�x�:#/ ��mV����]Hw�Y6�|�V����"��b�̀��D�vv��Ϩ�e��og�2�f�ue�av]LTJGJs�ȱ�n��v�����}���.?��=Z,�!JK�����։��v�2�&:�m&��+�4�I��~;��ڕ8n���]�m3��v
4����:��b,��W݆/�ި?��u�Z����e	�@2w^�+�d�`�_g�@���I���X���D�����mP��c!	F��5���B��Ho\n�pȀ�%Dۊ&��U?F�9p�>�<s#�EB��/�������1��޽+��i<���[��A�u�y~PdʫȈ'K]b�:ι��j���	���,0s7���a_� ��X�n�&8z�g�Z��Jϋs��j�g
��^�y�H2osܵE:ryg����|�w�?��6i&̼q��	��<�;�Sw_wa����B�B�,���Z��y�-����PޮS�,N!J&�Q�x���Bc"،�����tE>�_����Ք.ȿ�o������I�Y$ ����{��+s��g���%$/u"�G�Eq�cY���a�/���&$�A�/��J�&�q�8^NuDμeV�=�i
�6}u+���!:U{m���*~�L:tNr_�v	QW9H�2��@sF��TQ�W��$��-+� �-�F=p�x<mľ��RLt�})�x<'e�Yh;����|��^�����~�F�u.������^����tRn�J��$��ʎ�{Mp����"������_40���t��#�5����A��@��h4$�F�����MI诲��ŉ��Y�En��G���\�,kc��$�--�Ո��t�#�軝��2l3�on�a l0cE��U���%�}�\��� ��D���̵B[��_+��P�E�n�r�n#DXa\�o�7]�:�WE%�C�
���� �F�,U��w=�`�	g<� �^��0|Yh��_ѯC	���a=��n�8C)t�^a}��P�"�躜�2�<J�����x����}���J��)�twlk��.��M����4�n)��:�~�&���&c�@]�[���i�Ys��6�1��/T���I�zZ$8&���凎��a�RtWY��UQ�-�"�ߴ�H��B���f�����ݏNp�8����G4P�2�df����2}�B�'�s���VUIC���b�f �O}��X�W �ʗ�ɅmC$TQ���2�T��{f�+�/��Ѐ-X�R�i�_�v��m�@�
�ۤ���hY:w�3���tX'�� zђ۳�dI�Y��9Xř;����avQ&�[�nv��V9Rծs��/<��|@랰��'g$��ST0��z����s�f:ēe�M�M�-=�`�»������VO$�O�!.%L��((��Ho�{���2�#�q;+ϯ��vo s����2Zi�2fk ,���[+h����zڳXj���vg�ݢ�l�z��N{�v�q�<03���P]ŮK&+�P�1��1�i��ȸi"<Lڮ7��*p� �Am.{��% !j-������W��	��=��Ε�4���	a��itХi��'cB��3ǨīH�ޑ�nw�t�=�]�Z/%יw���٪�[��pI�(���(�SV���7$�.6C��ރ=4j؛#^��By�9p��q��!�#EK�F�ͬ��9D��Wz��~jl�Q��v��Мgf�^�Q���H̄�n"�3{o4Hl䬘��$X˟��i_��R��;�[��h��:(�̼\�$�@�/=�#��kbE�BC���|p�7e�4��� s�v� Mz+�k��x=ػ
G�����l�@�tE^��+�-4kds�
�h���9�m'�Ѯš@ЉN4��M퉼8n0��Bê*���i�|펌M�ǝ�j��(�ł�m�5F��d����%�aĒ;��v�d�������/M�y���Eub�l�m�<�)_���)8�I)<8)H����z�6=UQŢ՛Dt�L/����>8�i����.)c�Ҥ�	9��c�kvŚk��z��?r%Z���ڀ��jA�Gf׎θ'[�e�_���QqI���kY��K$������l��B�z3�/��H&	��1̅*��ƴA�r�n50g��v�����i�ȇn�ठ���m�I_^������?LOɼP+�W2�z��O�4+��U̜TK����)bic�krQ֢���n�[07c;+�4�!m��;��MF�ٚaClO,��7b$����Ńh2�k>����y$��'b�e⭼iժ�[R�vvdO1��)k�X�O��eB�sĞz�n��$��,��\^4}^lΈzw�?埸�5Qf)|�ڲ���ٌ�^
'�����v|�0�j���*6fҍ�lՅL���Q^�O����C�+�����B�%̧�±F����:���G��&jU\�C�P�L\u�]��Ӳ'x�	&��l�Mm�؀h2�FaF��� ��y���@�o�Yk�h�0\��t^����0�5����z���IbE�q�i�)+�Ǒ\7 �"M���O���=�	�6��p{�����0�N	�QƱ漤^��~�5+83���Y�yzW�~n�J�I�<߸Q![�h�F�8�*�i��a�>�ne��c�)�ױ�i�[��<A�3��7v�H2V�l�ڼ�>Q���4��*�/�c����p��\���t����}�C�>cX�wtK����W�Y3�n݌y]�L�C�\����0	�ʧ����]f��zQ�~� ��
�"a�*n�e�6����~!bts����A��T,l�=us?��j�O�#��Z��M.��������<�ta+w+�ѵ�ϖF�=��-Y\�PQ�)��+�rA������=}4���M�Bs`���UU�)[_��x���s̿�Ep
�c��%m�OJ�|��!G��zͳ���3���&��^*��F�lI��u&�*Ʌvݨ�0#�����Հ.���nt�}�&� ��(Vy!a����](�粢���R�!�5P��M�\�iӦ�����y]֜?2�8qC��[w�{�����;h�������d\��9��Ji͉3Ԕ[�����t-�.G�O�Z��5}��j  �׳d�ئ��w<����Ji�.8t�ҟפYeb3�d�ހ�]P{��4;�h�
�VO+�#R��9�!� �wK�>ׁ����>/�9t�@jL(�����`��82A�|�/��Ӌu���O�����Tof,W���q�@�����
PxL,��`�7;�w�(r9vMs[�`y���Ԯ2�3��5����߰������l��p9��T�[Zj9�/���G��Q�%��*RV�Fl3p�"�)�L��;i���1YV*�����ZU��,MU+��$�+�����J���6�l��]W	OO�љ��m��X;�eѴ�/��?�k$���PA�z�?s�[K�v�j`h�z��@�����h��	�Rn{�M��2��٣��]�GYqG�*�vns*��~��Td.{�F� �RQ8r���K�K�t���:c���}1l�ckA���T��O��9Qkn�����w�s�寞(���<��5�!ڶY)���J��(�:������^^��_�V_G�����}��$<�h'�teis�Z�sb-JyqAg=h<�2��.�$���
��&Z�4:�����ͶWz�GT��En��&�FM�͂_9���sDK��<i��#:��U��B���.~ (^�09cv\����-�'��&���3%�% b��]����Y���t7%�ut��X:
��g��{��D��T
y$�B�L7�7_�^�~�V:�w� ���/�ګ�?��Gʦ�+���A}_/��a,jH)W�\�CqiB�)��WUR GF�������,�Ǌ� ����#�H���Ǖ1��u�ѫ7������+�+�{��Q��Α��Uj�/y��X�[����3r�a�>:���?�~#|C��~f�tm�R���iY4�������_��)�v��Ŗ��4�r�v��o�	 ��.����ӟX��q��f��89g��?Lѳfq�ۂ�N����c�t����Ni�$\��p��H�N|)岆��h>�OWӭ�oC?f�>=�8K*˨P�ElksnG�;V�c]�W֫�7�$����s����_����1��{rp�S������I���Ĵ�y��& r��[�n'�_XN��6*��͋j�*��e� .����)��w��D�H���Uu�~������P�M�_��(4��G�{%^~�L]�i�,-��]lV۸'4�A�h���'Net,��IZ�x�#�=�p��⠂�B�����T��2wh�w�V&~,	�K����ՌZR�2��(h{���R~Np�W��T�( os��5IRYvc���LⒷݳ}`_e�ԙ��E�k����\͠H�*�w�%�%h�h�g��s >x����O�}�J������ڼ-�)/��]�� �V"���Q�$�(�#6\?��tU\,�M�Sr�����N����ko`�i�S5F=KD#-=�]Ŭ�x�M�@%���ت�ֹ�{�~zsgT&��~��� x���`3D;_z7��Y�㆒$&�b�|�[ރ��4�T7H������PO����D7�B֜�v�6��vg�wU�ê��v@��2��8�*��-H��	�*C���y�(�Z��m��D)mA��ݩ���e;�&#`�0��CLb>��+&�ל�,�^K�02��$Ԏ͘(KY-A+���HWV�x�*��h7��@�@~�"qt�&�Y��u���b0a8���`ACr�k��(n4z��G�Z�iJل�T��]������t�87���K�s��͑��+o;�P=�/�c��x��N�2iyxʍ�U4y�i��?[1�ND`"N)�����9#�t�{��q���jHO�%��;Z�������-F��%�fo���x�^�ˍ?�S������Ȭ�|��L]��w�}�2���!Y/�fQ��솣)MAڊ$V�_��g�)&]�`�[=4[�w�3�ӵ�b^����B�_��B����\H� �M���8��Vg`���1�!����ۦg;���N��"~R�.�8d�8�%羁oL�ڼ�Yy�6��6g�SJV�Z�*�� ����*��.m)�:_�%R��5͆Ӎ����.h
�>5F��b��a}���<������(�]?�V>�J�va`OMhi���}�iN��zл�-�zcI�cĈ�7�b��E�A��j�3|VZ^���_�����_���׈lK��,���0�vI�[5�d�P{��8�@VP3�����(_7k�Y*����� i�A�(�A<�ٶ�T����^��ۨ��'|0�t_�o���K��l�����ô�;b��B��C�1�Y,�%T��ʃ�{�h�wz��+��b�5�9�V��̄����T��'��.Q�#�:m,	�ۺ1O�m})�O@l��%��e,#�sn�sLz�W箏a�0#��mj�*�5�ѯ�V�?�2K��,�?8T%�:����E���MN�lZ|6Z�������Xo%RkF�{{�V���CQ�i�����S���>$%�w�q�x�X��������j�ȶȱ�.42�n慅�L/U�(z�WQ�ڴ���e�3ݵG���L���_�ms�)Z�d:�P�W_���$����MK��p��D���U�B����D޲������-a���%�|�f��r�Gh�D.3�FK���A���v�P�3'-�O\����ϚE�����_���[tA��*�CdmI`��z��f�A�tNt<1V����79�u�ulE{{���}e@p�Jz%�Ln.ܜH�{�j,h���m�ߣ�^�����"x��]�a��)����h�!�¹�YЈ$�_�+9h5�U��{5�D�
��R���3��y�@�}��X�1����p1-���Y��s<�}1��L��8G4�����ŕ�=؋5�x�vİ1�	λ�,*�f�mp�.��Gk7�kkDt���l��q8'�����њ3U�@K�JQ�O$�I�V|˾
�A�g:�+��5��?������o�fh��g��T��-��G��+��b�o%K�n�9��a�<o&�_�us��sdF+��H0Tʋ��ܘw��)���KY�m�7"� �|17ϕX�J	��kE\��'\�Q�}�x�>vlB������;�WMu��y�2�^��ce/Ih��4�#�gCk�:U����l1
<��P��<3G��F��''XQ��j�B 1~��?\�QUجI�Dm��#L91E
v&�f�IY��qcH��ق��A�s/������$��0gJuX����ߪ��6/����@0�j��v�M��c�j^��]5Xv7P4�0[�&�vG�췮���pp������<�~�;�m�l\����-1�f��=�3uϟ�b���KA�Ae՘�6z�V�ݳ\$i��dс�I��D�,�j�d�&�!� ��n��������MD1�q� ��/MGvж�ڵ�K����Ķ6��ok��24Ynh�"V@��������
���tNL��ڌ�ŵ�-t/�'��U��/��:�t���f;��o_��$"��gHd������7��1���e��Kֳq%�^����mr�KQ�����'�_;��$䇆��)�]JUd'�q�#� �g&V��:��8ya��&�n3àcc;��@}�
����M�<V\�%:h��D$*�v|?�M�B�CV*@Fz�&���,`�e�����������$��5�����
i���Mn�?�	U�I���{�7�V�@�+1S��.�{P㪁xt�]��������V�Na��c�QW΀uVӃ���	�]V�s1��t-:�j�0�lX-'e�F ,^��f�����p�;x�8���[)�Une�2�`w����:R$&��5������1�'�~�J"qѫ��-��,8(���^(F��������ٛ��YȊ{��� ��B/��<*�����Ow{$^�/l>�+��	 .h�"����.毾�郱�@�:^%�j�r@�-;X���%��K�"�y��'���fo��-z$$��9�kcď5e!�d ���X6�C�7ϕ0��V(;����~�� e�@2��ݜA�g'��{���b�uP���.�76	R��d���:�F@�\"'*s3,M�B1`���^����-��Q��e��'���_��n��!��~��PU�X˸R���뽣����h��O�T�����C�!��vC�@s�����k ���c��<���v���YΈ�?o|�<.��3r��n�R�*[��Cr�1���B<.@�r0��X��>UK��rw���BI��.�ٞ`7,9�6�wt�;�n�Ux�|��4���I|!����0[�c�&M�#/���	t��c���?Agþ�#�R�G�rk�Tv-��_4�����{U>-�&��yw�7����{9��JY���δ��"�A����Y߃����GN:��Zկ��;���M)M��9�?�o�VϠ2{䩸����%�f�YE��R���G������g� ��I{;NG�8��O&��Qg�����2������?͜�Kz�$���`´ΐC���Ā�W��e��h��3�gpY�[`����d���S�XM�<����|7Fs��ܧ��(�%2*�(>9�!�]K�7�U�Qi��W�)ʤm�A��w^��kz����z;�15G9�b�kXq��G���8�Zq����ZOEЙ�o$4S6Ȭ3�5����S6�	�_J��ǆ~M������	�����Uvgy0���������U�ZS�����g�����$��!Һ��l��A9��(ٿ*��;�N�3�$|J�֯h���:��̜�r�����,�Fl*�0�,a��0��~Z��,�,{�(n��R �4�^��r��6K�|�I����w�TJ�FJ�E��\�2���#&#�~���<C�����S ��+,:��m��z����h.!,%v���)�)G�:�׆�́��t�m�7@,n�2N5�����O$!�Sۭ��^�qWpzi�#�-"q~����p�����)&���C#�L���5�*; �sz����k�4e˻�?�j/Y�ŧ�m�\Ϥ��a�6�/�S��R7��#�Q:�뎼r'��0�HR�u:.U�~~�W|��Hj]��L�Z��7f~������y�>ûj~�Nj3���W��`yD�,�5���[��B^g�}��b���;W9L�_�J����4ʩIdI��e��f?�g��LɫF�ֶ�bY��~y�q\YH�'\Nq�5���e���Kt�uX[�tW+u�5S�V\���`��bP5����:��w���KJ����`UJFlg�P�%�:g`�
�sw���<�l�;�'w1,x,K�kb�
[zUc�6"�us�^�j�e�@c�s�='2n��������P�f�B���v�Ð�&����mE�
d��~BH\��;��{�>���7$�s���9������ ��CtR	P�h�b�F;|�Y�`�&H���ƣ-+TJT�1��Ʒ�g=p��4P�f�]��&c�>9��v�v�6�F�e��������g��������S(�"�@�Z��3��AwW�|�qGt�}-�],�san�ȧ�F�R���w)1I�Z�,ª	B�4��Ry��e���H��KE�i@Ԫ奖I4
Vz�s!�2ؤ-S�;���g�"�o7��ܚr��&(��p�xӘ�6sK^�:�~S�7��5����-�!�-�$�}9~]+���n��7|`����"sJ�l.�ļ��
�͑T ܠo�	�0�NoT���n��  #�A�� ��{��cZȷo��a*��(%8����>B*yw>�pC�л?���l��v���@���j�`��.��P�TI*���Z�8Q%JX\�<:��̡<�o�tH����YW�h�Ǫ�0'd?z�����\��-�mrcC����qa��1��M̊�v�G��L�<�r�:��l�&E�6���Z�%�`-a�z��ܪ�"�ZQ�P��i?�}�s��Ө��<	��|G!�L'�>�����+c����u��2%����/ �D�f�<M"