��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xMMh0n��f���X�h�ʨ���H�P�e�Iܷ �>Z{�&���|�@�X�wF�R�s�H����'Ʋn�4�ûD�&8��q���TD9*g?V#E��@f��l�������GEXT#?
�5��RZ�F�P�ޣZ�e�g��)���O����*L;9���
_���qci?6�g���}��c��0o�av�UM�Gb@��#�+m�m2��5�?���w�`�VSi��\_�}m0�];��qf��Y�*1s�
G�n��g��sir����,v��P.�ݛ�ލ�S��L>�%6@yuP�3T���$�� ��4H�ws�_)��m��U�h9��؉�`��z	���ir,9�
��6&����F8J��19,��X�2�:F?t�B���jP�r3��<vige��-��^;w��؊���� txK�N]nr�!�
0iPg���Al����J�����KF��� �^\��j,�Z�^"��-8M5�s?����c$��4��s(g��3x�����:Y��KlX�%�.5)r�M�d�w}���i=R�Tm}�|�2�:�W�F�AF��k:r�[Q'8�`�#�ZҬ6d��2��tAF-H�k5����3���X���11�* �{#{m�u|�ۆ)��ncK���S~��Oo��J ��7h�e���-��3m�$2�&��Q�4���̕�B{���-t�NqoXe6����Ԉ����֯<Vf���<�8ٓ��sD��ͩ��/h"%e�����G07�Pt�S"O^3�8�1�ǈAt�t�9QU`�SNk��εa܌����[&2��lXt:fi�r(��x�K�>��6G1*8w+_�o���.�ۡQُ>�Im'��I/q������]��mF���lu�����_ �/�yLѾ�\��o^��ʵ,��*�T�~1*2�����]:��+8y+iX[�hY)?y�����`�������i���ԂTp��xi�mw\���٭pۊN�ʽ�x�6'�N�	�	�ڪZ\EBf;ī�����!
̯�)�+��?�������w�,%,C�i+��"�fj-�YΎɸ`V�7>'������6� ?��K	=��`e��r��9�����T�zr���/�PM����A����)�2�00N�{7� lbP)zQD���_K� �=F6{��և2�U�z��D���Ie�6?���L�K:���b����4�]�'�_����=��r���h�'abES�首_rWZ�z<X�"w%�7�tr~Z�Ǎ)�6Ҙw1���L�Ko~�^4��X2��u�b�Bx���ޱg.���:h� S��̊�~<^�p0�>�C������j8W[=rqx�[d�-��:S�5���I��ǅ�R���X� #�����hO��T�p��ݞ�W��)ia��L�ƃ��ܹ����0����zI�:�U�A:�1yp+��H=}��ܙ��$���c���G�/P�m��n�V��v;���`w+��0l9LUN;����>�B
(�{H#D�f̚)�3$��d��~x���n�n��Q�,�"���$���%�w�#�	�
����mJ� -����U����*�D0TZа��ẘj��̗�*�D5>2)u���]w��\g8�?��Q��Vv��� եi����5/`�`�ߕF��C�3�;�� �.��l�Ӏ[ƞ-�3!�*��,�}D�۹f�z�D˪��?����J В���}$�c�A:Ԥ��@�)Z��bė5�hߞ�����9p�����E,�"��x�Tiuo8��H�!]�{�i�s�#��Y��Vʡ�}G72�&2Rڝ�XR�����8�J(�n�g�[���l��z" Ufq51M�Jo�L�P�^M��V�]���r!��1Qj}��h�����>ڭ=�<�\M�?����SB��ed�Qs�i����*�i���o�l</� f��üz��g�F���T�;4s�[*��'($��[�'M����D��9�썙�P����-S
cCC΋GPM�hm��.��@P��]١��@V&��/Da�mc:ŷ���iy&��z�}#��D���̨�'��z�v�	�V$Dt���>�}3��^	����?֌OR}F�ͅ�/	�����ba>�/t��0S.;� ^�
�'4M��r��⇗	?�AL��vF�D�Z�y��@	�Ty?��v�-����3�N���~��f~j8��ҁ	`�:M�\]�8Fp���Q5eG\�c�O��l���ף�eX��7����{4�S]�-+����j�
�D�R$��">2�L�sco/���uW�d �}~�6�n��0��Y�-^*�pF�[K�fQ�-���EdR��P��<�SݖB%Ͼ��p\u�0��m	�nKAV�p��Mi,g���O����t��3RR��r��j��G������&��0A�:�ch`)�� �
Fj��J	�z��:���p�ǽ�ߓ�������4��~��d���F��:8;���]�H
`m��r�~/�.m�Q)������h��+�����6�"lP�L�j�K���o��2K��wа�T�~���o���X�B�"H���6����!~`���٠�;�p�A��PXg���G�!´ػ��ֲ℁L^���ǟ�0
ɾس����2����c���Λi��.=z]'A����%�����[�jc���1P��Z�ݰ�;�q��7��`D��Z������ʶ�m>�=�a�8�8N�'L�a�|����I��3n�1��^*Cw��^:�ԤaE0-<H
��hB�U��L� �	�Jȍ�e�. u|���v��5����Et0�.��%�#���{3�Qn�x&%C[���/@�� ����eY� �y<w���E�*�i^����i��\�:k�"���?4���e�� �O�|�3�yP���q��TѲ� h�/_P��̛^��~l�aS�pp�w NN����j��n�8��ʻ�Xt	Ӟ��p�������V��f臚�IRE=w�n�j�U'q�xch�s�Hs$uղ���+p##��[OzM;��U�ah���ey���U�Iy���}D��tp�ޜ��gƂ�����7Ƅ}rI�5d���)�$l�9_�4B`��KY��spF��ҩ2���j�EF�`��>xm-�|���	�ҫ_ky��)����E<9>����du7�4yC
[I=�ٓ�=�!����/��g��7������W�d��<�D�?��	��ꇠ�.��;�{���S8*��	�� ��[�z�̯ݬ6�Ӹ�%�:�[�$��:��#���`9䜨�ua�3!��+d"o�p�������{�PK�̃N��pi�s��M����z��_g�b���������=Xs�(/X3U$�1��A
��(7�
�C��N̯O|���%T�s�)��w�'��f1N$�n����'�D2k�u͗�S�Z�jѲZ�X�I٪�g��~�<�;*��ec�:��}��2?��sB�&O���0M\�oԉų�ǖ���:�|rQ���okœGv;�!M�a�$]u�}}
�ފuk'hb��!��v%}�-�$�
�ֆ<!n!�<C&��|�V?0oM�zQ_P�G��>"���XЎloC��Bt4��;��.yv��͖���=�����$��#�ey��l�4�,�
Oߓ��	E��P]���Ii�-��_�-6؟�$Wvh�}S�?�% &�+���dq�J��g~�AޭD��������#�I��F31Y� �Qz\�D�v��z��!�dJ6$��g�����=�t$�����t��Ʃo9P*�1���[��0������(�� Ns���Qm٦���̓��n]eZ����k�����]��mq3�/b"����Y?e �Lo��"\�u�Js��>�@ݯ�\�A}�O�5D�1ķ��º_�ϭ�yQV��0:�?���w������$l�.qSK���Тq B6�u*/H�V�\?Q��MA�cbd��/���<���x5>X�2�a���BA�i���/xCj����XzaEG��x�����܆ފ��ܤFN���#�$�{>T��+_���.$�a8��.H�P5�s�oucKG�?�^o�k묬OC �����o��[�����T�mq�G�v|�m閜�'0'#��A��� ��1�^[���m���>�9>��Ŷ�F��}�n�G7��=�D�#��}mF����P&Z��Թ�M��EG�k�T��YQ� 3?q�����3�r%���X\���=�?�Z�g2�9�+j5�W1��s����wSˌ���V���QG5ur}T+����������+��]��\D��m�/@�߂�݈�CeWE<y��"J�J�����]�f�H�W$O�1���������D�@Z��R���>�E�`= $�ڲ����i/���U�U���$wS3�A���Y�oZ72��t1�z#b�Hɝ8������8���l���'"ǯ� ��������vS��~�T�9"�Y$KhW(�$6�	�v��Ӭ� �J�۠��o5��wL�iϱ�JЈp~,�}�����*?!��}b~6��\�q�X�3F�ƞ��9H��W�  �$��e._��|.��}��g2�	c��݄ｵ�c�y�/�j�,��R�u��TIa7���o-��5�H��.��!RP $�x��������/��K��C�P���R��ɤ�l�^���}�G/����ZZ a�;N]T�b�d#��YAJ�E
<�S���8�
�h�ͩ�	�G�7ǩn>�u����8=qJ��~4 Ft]�Ύ*�7���A�r���S�F�[W{����{圁NY>}�P��P���L^Ƒ�>V��S�ۄ��+��4�1�w~.{+�8�_��/�3�ҙ�e��\���t�H����s�vgA��k����*���
+ j�!�i�E�l����`��C#��n�0��v���J��kv�K6r��,e��	�҆�(��ݿb��B7P� ��A$D�Ƒ|a�x��D�� �KA>A\��X��CA�wui nP�Py�)�SiK���u�)�"-�s���b]����(yn��"�(�=>%�Q��Q$� �D��6��p՚�=��(ޤ�<���\�"������#ˢ9�z������x�!_��#Wh��ᨹ޼�������V:��+��P@C ����=�q� 	x���['���l�9�H���M�`e�8�ڏVd���� m}��F�����f��+Xfn%�&��&z$>����Z-7,������vAϝ�&}@�^GS�{�W�$N�w8PR��_6.3^���E�]���ʧ��T�D& �E���3�.�	\^C�o�C�[v�7ey�M�p��Ć@,�p��';W����k�!Z�EfUR�u}��G���}�Kx�3�Ԫi��dkV6��L���S�x#"#�d)�dQAbD��1,邬�u�\�j�A�n�}0)OU'��H6 ߸5Ge�L��
�`J�'t�ndH��ᴌ��p	����ɡ��d�2�"�f�����O>����������:=���@e.����6�S����� f�Y��P�Q����W��5��^	����$�DS�h�����5ܤ�k�xo���� ��l�^)$�������}(��17W�T��qX���F`8����P�R���`o���$�������tsu���u�9$W���l�%�C��J��>�b����'d��1��	ƒG����Ø�y=1&��a�#ږ���+�d_N���p�<y�]0�>�.!��2��D�����A!�"�9�:��Ԭ#3��
�q�A��dGH�[��ʌ�z-���j��w
,��@�1�,�=�o)0�p��8�����>A��?��P�R�Ʊ�} CۭjM�*�2$�6r��'�O���P����y������ԍ���T�8ھ�-9o~w=��$��4Qt0��a��7+�PA��6��#xr�ۑ�ހ�)F��jg��	����xLa0�G�I3Na�@3���
�����P�!U	��B�`>��? �h�:�y$5����L�X]�Y�F\�ƃj�i��JS{�����d���ޫ��	:_���Ba�^��uG�:��ǚN�qd-yM�vM�(!%��4q��d�xI�V����N}��%��E�4]۽#�`8����qOi��FI�$�H���B�����^��R���a*�:!�d�-����� _�Fv����4�c����[eb��Xۏwr��8U\�1�4��q.z�55��o�����Vd��Ҝ���K�iZZ~�����˝]�䒵I⠊I�n����}9o=މp�(���n��ivsw	�_�no2�%������Xk�J�|T 	QkLx0�Ӝ"�x�X�bp�JT���w^�H�	�{k���^ �d�w�Y��qBϴB��}����qP�`^��1�'�`�'��,9�ic t��p�4��C+c EAs�ۄ�������ﯘ��؟�>݌���x���;�|���k�9&O��J�ET��_�Fw̅����4��2�Ow�#Y]���Hp S��A�����b��t1��ƈ��;�;ġy�y
�':�y�!��7њl�x70��ؖ��h
d�d+���q�23	��G��{-��kӎ�<�tGZ��qjoׇ=0��9-��E>����}<|�j��}q|?��&:���6�l�.�)�ƃ�%�(��������}�~����؂���\�_�Y���HlT�� �5��Q`��Q�Z��Ͳ��ElɿF2�b;�����1�&S[�_�+嬃VԮMK��j�N�(��	����;Y�F�9�Y""I@�[��؞���0��VdD�w�FB��eNϡ���|��,��ԇ���'��y�ܝTW+��*��0=�6���/��Ǩ^	T.0Z�����%CV�k�1��y��q�����Tk�~����^�V�a����i3��B
��=�ˁUF���\O�y�Ab9u�ӑ�$x�N`O�S�md�Po-�G������>�ʹ�q�d\.�^b�YM�cUCΛ�5}��1q�N�|��U��+��ՙ?����9n���w̔|V1�(2����4�H>]{庂��iR�(��CwBS�M��'�EQ�����,e��\����>�� J��R+�"��U_��̖29d
]�^k(�M����Ig~�f��țI)x>���u�s��g1)wc�2�T��U�|n`m7��s���zGEq�����։����l���L��S�#m5\!���3�<XRfQ��|�Et1+�+��nU�c*`Qj%F[Ȯ���ܸ�:�Y�[l啂�{s}�B�Udϭc����T�0qk��G�k��|i�3L���5)a�k��
����G��~�)��E�4�%�x�TW����k����@{k���	�C�4�zT�hJD;0 !������:�6M�V�46�+?R�h��o�ӑv�R(�W�3|l2��M]=�CfYL����^4��l�5�h�K��RD )6��1���$�T
��Z7ں�r=�ѯ�O�7�U~41��,ps���!�����8Wd^V��ru�匑�q�h	�P4��,��Q��������aȓ���6��{�� ��V�oU-	����U��"��S���}TU
��?_)ž�ˤ�2�x-!z�D5�!�Bm���-�\)�q��U��%�rǮ�� TO��ш����)|�dr��% �nt���B"H�����Q����l ��R���z�!��I��sI�Ev�I�<w�����/?�����e���q_5���p�+뚺�k��'|���j��J;�.���%���C���!^2u,�������A��46=('T-�{���oD�ߡ��]��(�*�Ut�
�ޢV��������Bw���;�P�X�lAu����@��rA��9X%�=V#i~	/[��A��ѱ��"##��ΣO�N�:U�^��}b�ļ+�. �&��p�Oވ�G�7�l�����a�X�ʛB�R���ۏ���[�Uq�U�ǧJ��ܒ�K�a�HD����?|��YJs'lZ9k?)��>�M
�7��QP�uQ>F:s�2n���V��@��\�U%�}�����"^�+������v�?`�J�9a��o����y����uxA�,�|�����Ü�幟~�w�;�-��	W�~�!�v-мO_��� L�tw�O|�ፋP=��Q5�*�O�A�m���Q���7��mtO�_3}�C���z6�Ql&��ـU��b�V��� }"&d_tj�v@���Pg��[��[�������Z�D�r��Hnn�)X��I��{n�^.����o����˜u(�Ib���^�.K���JCZ�;��eiZ���O��v�Nz�W�7�<)7W��ʁï���͒׏��-�n�.ɺ҉�5���^�Ρ��q)�{E`�=�[����ë��g�fD����a�7_��� �|�
�r��*�_9oUqΪ��Ky�2���+�G?4+*#�3�J��e ����Y4;덆p)��P<�J�Ƣ�.\:�����@/C7r��(��-g���e�1�1%���;u"F��L/O\=L�	3w,�)}�������:�� sI�uH�*�b�bK�=�C�dI��
���N��V��"�5h�1�H���E+�,��}w�p�45��y��g�4W��4�	�R/ _т��M��	؋x�ϣJ+5�P�d]��ߧ)��oa#d��*�@���N� �����^�Pr}i�m��@p4�d�f1睓��WV���
���4R�,�C l�ag:�
U�4gF){ʤo�ӂ�E�y���O}i��Jϫ�̯�+{����J�4�|i�L���u��@e��6;��?w]���?��Q���%�ˢ|1҉����w���YOn� �aF�w�BX~U��3ɸOat�m)�L�x+ۍp��ĭ�N��Cf7����c��F��7ɯ��`ZspP��[en�-[�xt�v�S���+��^|ΆX�3aNyP���Ez��F-Q�O�2�:`n�������F��,��s�7y*`�0�Ȑj����8�R�I�}7�_�W!��O&�p��C�Z@^�� �8�&&�������#��3]y ��x;Jw�n�@X�s9��C�iom��)_�S�����QVXp�F��}��.}:�b_j;M�cm W%-GD�`U�,:��Q���I{>]ú��B{�� ���"�|{�F� i�gk��C�\+����n����m�.O]H���� ���c^�/���Ĕ_���G�&�a/v�X�hV��JY��Oo���G�}���!t����4�����?c519��>�R���a^�^{�����H�5B= o�����5"ET"A1���2s(����X�`�Z�:e��m����R ��/��-�B�x��E���E�	%��H��n�i-�B'#-��h���ޑ� �Wjg!)����4'�e��A�s��u�"ׯ��]d_�8̑[�e��$��JV>
��L�Re����<wi�<l���[d#K�Af�h9Ԡ����[�B�༇Ǖ���߾1����������B}tz���mܲdyzRbXKK����[�b-�Y{�k����)X�c���9>������_��-�\b=]y[����`�T�@Pg���>�����6E�����!Z���ܒ���ﮣ��kq�'�bDB���,�NׯX=��[�*x�h�q�2�X._�+