��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG��%�}~���~�<cZN�X���Ĳ��Y��$_V�(MT��Ĩܠ2��l�9-S������d�����\������ U�̉���E���A�{n�g��r��*�q�@���_�q��X�5��YP k�١�u��|I�Zi&+��c���tʱ�e�R��On���u�pu?RM��2�Xd�P��1\k�R]�8h���~��!7�����U����b��n�z�>[��DIK��WN2�yz� _�0�\�x$���uw~Ozʰ(���ռc s_��һ �n[�\��z
��QC�)��B(����SJ�f�Dv�&�����y��W�}�0�,Tݗ���'U�jcҬ��Ǥע4�n��|sK!��m�`�-��������^%�]h6����e�.�E��~:�z׿o�_[�c5�6Q�M*�J���(���n���L~|E����MZa�m/b4�!y� ����E�_1�����N��@S��y�����J+ �<��
m�=�ϳ%|���m3�<�v��5nT���
A�<5^|z��V��\��I��A�@�akjd��9��%�g��k��Z��g�e^��@�>��!. ����գ�2�F<����"08���A����GQ�x��Ԅ&m���{y��sɶ¾
;�Ӆ�78Ì����	����YF�g��q�����X�?[N�V�u�?�5�Zn�����U��z�N�2O~�x�
�����Y'n@ Pl|�t��Z�\?�ڦ�)���M�Õ��7�O�=ݾ��x0L��7pـē�����ej>z�S��O(%)$�5�5�vUg������Y¿Q杻f������S�A��4t	-F xdϺvި�0�ܮ[�)&���.��	Z4�"]􂈣0r��)�܇��C�Bz=*��O���Ņ�J�b��oP��3��>W�p7h�y)}�/0U�L}l(�єEC5�w�Ζd�R#A��i�Y8�<7��*� ���h��J�
�9�s߄���ݟL�1h�r��pyx����)�7e\�v�B�;�"�(3�ӛS���j	s���FH0����6���#o�l�ys��y�*MP��ܨ
ۺ���X�bF}���.c|`���2�ў�{X,�;u��sp��lrhcf��mdl!sV�츦j�Q�BH{ֽ%F����m�{mjO�.1�)F$�!��`3|J�-Um�"=�\�,��[�ZAF2O�pLȤ�s]��X�K���N�:�m��ۈ9��W��s�lSÚ^����CI����L35�cdP|3�����[��ʃ��{���dE$��;W�
.õr.�1q/.�� ���s�-Ī�S_,��G`�qa��A-0�xQ��d�٧��F�B���%���ʹ�u���d,3� '&��\�U����������,��FH���D �A4.��2~�U����<o1��X2y�Y�u���7��'NOg��8=t�Dt���I#I����x�U�N�z���R�l6��(���?#��?�,���|؂��q��5��8*�:-�oIUB<38	���|W�5�>���G�� қ�׵��wY�����h���-_� ZɇJ����Wȿ�|�F�pT��z���������t�M�LRH��%W�];S�2�h�VmcU7��m���>9�c{a�)"�+��Z����JV���t }!�tG>�ϢwY���p\)Cj0�d��tN��[���@��g���U���9Řj���^�%��y��0Q���,[ �@7@͈>�j7����p��#c���S�c������
�.7��.��:bu�׼;筃�Ļ��z�T�s�.�fCٻ�b'j&�����A�=�c��@j2˸����V�tIɄ&�(��)1��Q�]7��^t 9���ʁ���6�I��
?�'?�#y>��P�����vk���g5����	p��`�~��9pz(ҷ��Vt�d�ǽ�I��Wa�ui.�*�~�#��"�'+*���c܊�vu ��ت/�K���@�* b�53Ȕ�O�u�Xw
� �mZQ�mR���;��b����O�/3�9������-�AYP�&a�[}Ab�#��bz~����� ?}�h�`�
����	q�`��Pk�x�s=X��f*Y�2�M&�q	�]i&j[�Z]:?��# ie5���&a���{ǭ���3T]����T��Y�Ӊ\��\j�j��oq�	Qơ'm n�v`ԟM�FF�_WO\F�J�{p���5�]�L��m���-sa�y�_�UQ����:��`7�Ì�h�k��% C(��W!1{9�O����Q/���:Ο����%yp��웇���0����?b7��a��狥H�3'���{4(�o��N�L+�2���Ji�G1[F�6���I��� @��]7 "�,<�_���Q`�����-���_���e����ױnQ8�A,omAzU.��5J��I,TX����UެcZ�3v�9�Pc������-���ՉX���sM�������л!ikd�r�C��9_�ْ	�dp+����V[�nu���Q'��^��M�C�m�[?0|���T&��L����� `%��@��)����׶k��w���j�ɶN!�J[c��)m�nUC�!ĮU�,!UV�휶1��-^��rk#���_��No[W�3e!
]πvK���o<ջ�p� �`�����7V��ރ����"¥"��i�^2U�������;�,�)t��.I���U� ;����r���긹�� ���Oq'Y�)�2X~��}����"(�ͬ��լ�	vw ���\q%�U��vqRĠ���v|Y��<��2�������=.�.��5='�:�g�dv��>5��C���3�_��;���*�ϼ�)0�����*�y1�߮"NտK��|�ǽF�U���y�e�Fٸ�e\�}.���8}Nιx:��;�K�A'wd8���%�wpH����f�l0�uA6=�fN���z�T�ot����m�ɢ]B��������;n]�gY���ҍ0�9o��wA\KDs����}�\�G���Qo����	oe�=���Gzu��6��<r�Ai���'D�T�q�V��&�@$ �'���/7��*��A�/����6]��b|?��˱d(�R�N�φ�6��0��ia��W���<�uG�e�� ��]�ӧe��*@��z��y�M�E�vX�88y�_�thU3%�P>�p�;^A�Ō�l��t��eH��[���Qp�=�ۧ2�� ��D�9�9�L��k��?�Zץ<�r�~9�.�N�'A�N��A�� յ�tD�ኹ������3+4����$s�ͨ��~����,�R�T�?�6�r z�G3h�w�n���u�{�e�O�na�j�R�}뺕aŸS�d�o��Q�D�[+�%�s�\S��=|`�0B�3xǌ�\eGu��n�wq�}ka�.6~H;�.���,�8>�Yۃ��%?}i�qh7@OV=��X�@-N�����Nu�)�Ť�ÌG S�}X�ބ`�s�Fm��s�1\�h۔��V��zm�tƎ�?N�]\��]�zD_�8]h�hY�g(_��$����j�k�-{:X�-)XҐs�Z��2.���u�D0�.���N�ԧ�<��sDO�-�|CGo�K|H���.����`zkP'<׬�Y>��n$�a;9�=�Ǔe��$6;ΕPG�ΤH4�5a���(��"ġ���Pf4<9��+��)\h�JLBr]F58�24�-z��g~.
�|�v��zW��um~4)iv}m�3U)r�����=�H�n��}�֏�H���6oxv5�ݭI��U"G<thg��+���^MM�	>/|w��U�F���D�8�-Z�9F��|�fyB���WP�Q�z�ۍ�����1W��r�V�Ai�q�8o�#�qf3�N�>�p5�r�n�P��16 [5��'z���$��{,Ԥ���-�xD�~d������N���㹕��̹	3�n�A��s�z����JR�7�W)?I� ��N���]q�FZ^�G�6�Yhs3M˘$ږ�ևE�u�C������l��R&-z��Y�O��jX��г4�M�{h���d��rAzVl=;���0��fD�c��
���&Ԃ�)����`�q֘�#I×��s�]�r��	�u��C]	����0���Ӹ;�mʆZх�e@������t�j�T��^%��z��h�X��N���xz�������ο�����Yr�R�d9�7���i,��*�LV��"����	ʾ ��I�ǀO?�������<&}N��
�!%��<e��vȘǁH�U@� ��iR�[��%�Էt\����3Ye3>�	)V:Te0&��0��5�*����x���B#E�jb������2���_"�p��OMA;���|Q�d ���GJ�d_c�}������u��H:3�@����p����kF]�cpe��E���� �>v'2�T\B��TW0./�Ю��4(}���:o��aN��U��zMx8͠��\�Q��6���j#}+tu���G��QM��ZI�����z��^��r�)�7|�;���0��ҧR��6��C=1G��D�s��P����g�x��?��
z��{ȨW>�>pT^�'_2���v$�g������x�v`F�g�\�2h���/��F�vC���{!ꃲ(��l�}S�2C��&���H�� #�����Hu	D9^�a9�#����/"��ߖY��n��Iׇ$��
��O��{�I�Y�c�M$�{X�;�*�dH�ӳ���f;(H[C�Q�S�F�wh�K
�Ӝ�-�W��d'��Jn 0t�I�_��0��i�bsh�o|X،2���0�v39=(�4��9�����Kk�P�7 ޹���ȰO���ð�W�Ow�9ּd�a�/R#=HK耡u&��A!�;���Z��~����H8K�@3��VAҫ9�mf�!�}���f£�� �rC<:�)쿾Bo��OnV��q�|�y2������GyQ}_����I����ލ�NW��6m��貍����>��4�n���3���TH�C��zb�z�:�[���	aU�;]����1�tz4~Jh�Q�j�#��r��d�e.B,���?r