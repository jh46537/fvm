��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�c���]�uJ]�u����`����#������`��`��yu��;^n�A����b��G����I��+�L�Z���������B]]�
���a��5@0,�@����W���U���Y���p��1�f��?�ɗ,����j����n�{.��Ƞ�$'=Yr7�~k��$� �q�;Q���'
n;M+����JH�����B��Eh��ݻx��$�m�R^`컔@I�f�|�9Tz?��H�s����b����F2<�n?߄.c֤�v��c-^�]j����oza��Ɋ_߶�Y�n:p�D}��?��Q���질�"Lr��A+���s�BK���,}��ݺa���dg>�`o��NZ��H3��������'WD�7g+�UZd��t%T�l'��g�0�L�0[�
O~T��{�B+D�3s� ?Úǟ�u�W�68�{�Z4�|Oۓ��&SL��� �����|s�
{z�v]*���t���F���RYr�B�d���\���LC:f�����o���Y��� ����{��Pj�����*����l���QcqL�ZC&h����Ιl�m���#8�d�~=<���P�ؚ8J�h�P��nק����Qv�.���ʃ��ɇ�͞���}�f@�0��c�HWHD���y�⯛t�Cv7%�M���l>�H노Z���rƢ��v����WZfd3Ʃp�֭�I��`l�ٻ�dR��� ԷT��o��I8h�y��G9�^iƄq�_��?�-�A�
ط�j��r���)�
��������K/��%.��;:6qe퇢�mZ���h�,;O��/JV�w�ܷ>Q�;E��o���|E�;�,�8��;�\��(��8��uNM)��;��ս8_��W��%-��}k���+��ݕ�=��:y�h׺��a�2���{���m/=��	^�`��ʁx��*��)5/�ѓQ&%�S��W���T�"���?E���&�U�t�g�T��⤼r��鰛�M��,��8������a(������S���a�J+k��Ҷ����5���gV6A�lj��5��=e��0����7J��U�ۓ{�$x��E�I���;
���Ts�6M��f�J��jR[�M����O�<���H��3��q�;�}�8�'��+���}X�)���<2[��P#��'.艬L�5<xJ��ŝ��X���"C9�����;P��7���pp%�*��ԟpt�j҄�)pB0u��q��߭L��os`p�f�n��P����z��8S��?t7"������S��ڷ�7Vnb����z�:���%�5�R��@�׌1�Y�y<񾤪Ҏ1��ãR��~)�[�kp���잘e�gp}I����$�E���M������ɳ����-�ƽ-�g��U�U�O�C�k�[�fj�嚢���]tV�$�ͳe�t7��e���x���V��2EK;��d��++�#_�E���Wm1P�o��޽ug#F��j~$���c�p��C\��O�dI#i�{���kw5����������pZ�wϛa�v�8�M�V-ω�H�yPĭ��"�;��vi�9��Pk�3<7�K�\�RM�܁cg�I>����C�
���P#N���7�i�?=���{o.�������1<��Wsa� ��(�;��IiJ��5�R,ajF���g�}� �[j��~�8ᷣQ��k�� ��[�O�1�H�h��!RZG���A[���/Mcu���2�v�֌��P�㹼M��?��?�b�_�B~��,Y���	fx	g�&�Sou�+V����tه���Uc�tX����qP̖ݲ�C�ԁ.�\=�'�~,/��VM��g�M��x�R�r���1��e��ff�|��F�b*���^�<���F�Y٤�#f���P�Itܺ�ͤ���,���59Ǯ˂V���{L�]6���t���!*���K�'���wD���V����91�ǫo�( �r��E_��s`����YT�4��?�u�HH����Ç���w�
�o��1g��@s�ʦ/�*���Z�w�1�E���o�PRa�����Sm�=Ց�!�t��ӭ��T8�bYh�u������|e�e�3o¡����L�! ��o$���:��kXt�j{�Ϥ�j��;I>L��<���-x�#h �ih��t*_�TRI׫~�^�*P��[�i��ud�� ���ub=i �x:fD�}P�턻-G5}�X0�Y(8������ɭ�d!��R�2;%����� ��t *�t�Z2�4��%���j�$�%mQ{�]�Dʣ��{bԲ_۶�(U�&0<�K��à�n�������^���ʬS�T��)�<�n�=�����>N�r'���(D���%�u�dCZ�1zg��A/�ڰ�&�}sns��k yJ���e?������6	i�)	�t'�/"Xa@��d�|w3 7�3���>*z��e��}�k��_A���|)x*�z2��:U/���<�q���Y<w'T=kG�M"`��ҤO8����2��H� y�؜������րwK��i�J:َ�ŧ�c�`=�n�P��~ @�F^�7���&r�Vc���j�##�*?⽁:	��5��O41v�� ��>���%�*X-��.K���p�
e�3ω�9���*S==0C�G\�Z#Bث����M�O>	�$�1���S��/��5��nūڿR"±����#~@�=�w����	��B��\����.ǌ�.M�1BW�i	.#x�j���[�����
T�