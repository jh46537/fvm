��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9��m������G|S7���X� bU��5V*dFi�0����X���c�j8w)h�m����Aַ5����z�t�T�W\�hdY[C�ģ�u���V�E֦V.j�])y�p�`m�u�O���(��YU�C"�)�δ�3��*�@[��7p�ɠ��͞�!�J#�#ڇ�����ϧR����!�>cƌhb�%z��	1'N/Pz'��`@�A8���=���s>�d�?.	!�+|y�r���Bc1�7��"I]�`K4u�4�����]�,�E������a������iD���D�M�0��
I�h��y��i��#z:&f��I"��z�����~<UnE�����ҁ�<5��C��5w�aD�b������wS��o4��L;5�(���,0,ކ0�dM\�\�T{�?�nkN0	
�ju�Y�������2<o�����܄�+�j��r�~-�a��'q~3~�&��-.E�/$�{�?I@���E����;ͣ�o����Sy�#߿,��x��H8p9�K"�J!µ�+��W��y<�z�+,���"-GA7���p�
O��=5`� f�������'�J�׫x������B�Y�
W�� �����oХ��L%�\���O&�ʊ��`ԛ���[t� ff� �J�0���H����T�
d	Y�}R�?�6�DG�ƈ���X����>	dg���;O�*	���>A�������CL��X=}�&l����ˠ��BW	���$�c%���M#.�{��PMW>���y�Yp�:e�7���Q�}+�w736��=j�w����Q=�1���G~-T�6�o�K�f�s��O�� ��&_���8�����6��ix/���T��BhB�$���(s���YF�����ę �܍ �����~Nd?J�*i���BP��֛b �6����c4
�����jo�=��	Y1RJ�f�n�7�Ўu�����U�_�$�(���Dϐ�����tq�)4o���iH����R�Y�\��J4t߫���F�jJm0�0_rs%�@�:h��~���gCj���R�`��yE#��!藅���N�K.kor6ṵC{�v�Bm){�Q�ɔcފ��c����s5��«[iʞ���*oI�9H���hCfWu1wn�E�$yR`ڹ�̲G�_��Sh��{K����2%��0��زD#g���q�����3��.C_*..�BÍ۳$���)܌�3E�� &༢������8����-Cf���aQiև���e�N7���$��ה�[��F��gH4��&��2����kk��1k��aބ�_��n	������Ħ�⵱cQZ�иŁ��E�bV����u���I��%�0�:l�Q��5���F��ҝ,�J%~xm`QF��W0wi�)pǊ�L�bH���:�����s"_�>r���>IZ�Ev��o��{�<�CGXL�H���3�l��`,]G1=���އ�����J�.�-۰����W�6176�s�9p\��p9x��Hϓ�b�!�V�[;���B"�O�~j�Ѷ���h�ϵ�q�d���	��O�_�\GX����Yr3y��6��t�2/kɹ����ިS�F
����S{�\��aݭ.������u�j�V�K��X1nQ���`�k�q_���?�fV�����O��h�@��Ч�q�_���7���qC��,5qC�C���X}�������"�Az���/d�H�V�D�P�D��u���l���-���VH��x^��F<	"L+�?ΐ�E�Bs����o^�A5���S����
w/�8,�kh���"���=,c&���Fr���4�h��x��T7�G���YF�c>o�m)�G�I�u��T�6��g흇��+���>Y�B�k���U���Q��HO�}�7Q��a�A�������L��I��h��P]�KM�45��:e?����׃,<-�Cy�a\{�a/+��DU��٬L{�)F[��%�/��e�vv��B��n]3��=bs�|�`Q����{G�G�Wqt$@�@P��>����	�RqA�V����P�v�޻�.����-����$�B�zD�ćN���Kʕ����~�1�1Jw��Ri��H3-�)hJ.�"[|mE�?L맂�dMͳ �|�P��r�=�Z0�_Ք;}�9�#B�<�~�ʞ������j+���i̦�y��W%_C:F&)���r'(0�����$c�����ѥ_�́}/��҃����xHm[F�>@���Fzm�>�o�ݿe��q�ᮇ<�T)+�&Y�F�K�1BD f��'Z�$P>���s�=��;tR�}�>�|i&��Tf�����?�^��J�;�k�y�y�sAu�w�9��bw�@��'��YI�X+��@q�������g_��0�H�]���Pk2�d�T54������s!K���i	��i�����1�iq�
qLi�`.`�YO���J4ɫ����'(��FW�=ט�f?�xf�.����\��];bYղ:4�Z7"��J�h�r(�r�e}�u��rdRU����� �j���qx:��"��IQE���S��SK'k�A����_�7e����a�=b������f���WRm���G'ȸմOEM����NC>��c%A+c��c���8an5f���OB�~"3�6� FЪ��� �!w���T�?h�LAV
��'|k�/-n��eZ��F���Z|Lm\͟�Kޖw�>��ǭ#V��