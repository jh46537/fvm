// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TavtoRUH5Rl1SxPhv/SDuuJP/urJ4vBaohwU1ziMlIyX64fZzjT6c0rrATXgno7A
TqrxIIZvGuVqMYkadGcKh1QFK31HkrH+2AKcYsgntWb15ejN5GXAaRZin0FJiybT
CK2GKU/FrplsE1/ZdSnr3XWJHR3Vg5x4roMKfQnlxQk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32816)
dsHrNGqSui6rAoHRqSw2WqivShfRhG803JsomZtzYEZokgEihnxjAa08pAHLVu15
N4zhHiilZ3eZNI+UyvcKRER1q45yF3kMUnha5bjzxS+1Zs2WhMyHlX4C9f7ehPCn
cbYrd46mI8D4/8+HX+e3uxjTFGOULACu7A6P4LaQyKGhwwXM0/TIPVmOD2a0gc07
EMcM4CQbdUdZeVsGT7mEEFxdT0IRWlNaTRM4L0yb5p8U4sVzOhoM43ZTNldflBAI
X+JikZAyOsLSvxoOdVyrGQWMZ35VFO6r7a11I12Nc56VZcHUIDT74A0kuGsLg8W1
9fdAIWRjAygs5dyMQgrYK3M1VgN20ziLUgl9n0VgkxciNUqxdSbni1fgdLXn43R3
tPsdUFlJCWLWdfEuikvc5J01gchHas8lx5c4RF928Z/2YxAyw2Jnd1EBRA/V68y0
Ed2oyj+dx/WTiLiFbmSIjrFzBsSEtKPNeqGT/8jKIJ31JXOCGI6q5l5dGkRWeQMv
B6WI0Tbp+VBxkHHT4rhoIqdL3CMGCqyXMlmLsq6sMD0gXB/tM6PyMtDmdAJ6irDO
u2HEz18CbvmQ2Jyl7uKci/JMUQpvQMYNmRm75kOVKglbU1jd9Y+x8Saa9/WGgs1V
6tTa888a8YOas/oPWGgGzzxKieC3lJj0M/dR3cTy9IXZkkO0jsKVecc9T2SuZVyC
K7B3K7LGSGt33ZOHd32VF83C+GxoYLBg8uJMC547dulFDxLyz3Iu9CFsOsSZHg05
iW76gCcyRcOU37IzACOU7EN6veBDQiB85OlT097+FG8ZUB2X1W8xqo8U3EIQfgdU
FJMoAlCvh21pPsdH1rqTtlprWGYUxbUUpCNiDqvVSiQTi7KxMcKG6x2ZbZ0mSXlI
qOn+DIgnoMf28D4fhFDZhtGluAgdkdIHJUAZQr7Qodd49PLtNAIQwUqeD1EAixwO
2iEQtPNV6cugJvGTg4cuG6SJPau0EKpRSQIJiDxAPCWBn0VNc4cd0nMHs/GsTgNe
5DU0hp3fOp2t1H7j1kogsUQVt2tTOXJAd/ro2i2s+6pj13cEZ3ou9ZqXI19FxJ7E
uSx5UBElJkY31B66Ox0W7xtmphOh9KS8TAr2mOMNxKl2bzILRDSA5n8KE/VNK0LC
tGgBBUkKlShN8+6UqAsEn55xWQPdrhdttUVgZ4cg85WNWJeCbsoafO/UQlGnK46X
Y86Xl8QmQsWFFHb3ymAyX9VQP3BXDlukfAf1ddQ+R206l+4pXJZHeOGmwFbaslA9
ja6CbtnaPbYQlKQZPgnjkFR9KEFa2wMGfcxe1FyZo+j53Aqj+TIhLBqN3sYXKUgo
JAPJm2No7Q8IFcxTXWjd8MwHsO//5uhpmMy+zeqgYIfkhPsYvrWpOTLx8WiYlmae
AOLqGIVtjPMn/x87L4PApXCnJe9GOza+F0UppD8SsIisZLMdRpADMMyJ1KuPVcSB
kpn2Ra10vRq+rVbkF7dv3kYHbOmPq891aPmklvotfkykxobKSDBZdIW7K3eD3K4s
k+8caXBnIraCxVSbk1CUWrux5vEzhPiayNVpv5KmmWsZ5UT2jNuSfKhJG65VmDS0
Jgq+jQh8TUGA7+lspa7FDgpyMXQCWSx3Ag00giAfSakuD7awAJ3liGnCsAhRiehH
5K4XJyrAAV0XeXDfHhUQTLrBfjPm1PbipoJOAJklKRCEhVgQmBfI9Trw04yxspUb
uIC+3Mb9xu/OHhFa4n7t0aqAHFx4ar5CeK6LzsyyTInizWo/aRpavUxJGyPCKVmU
0sdaP3zYHQhLM96SSa7nw1/hHJFOHpXR4Bn5Ohy/R5ZKThUzvewQgBNCmhiVGZtf
I0X9D0ua5EsQoh17oe75fOMTzGcyCrvx3Gg8LYNbpCfdRhYXcTiQyaGmno1T924H
o1yUwnZo6lWmmx3isp3mKTTUUZI/2W5i0ikHjNWnxvVzhxuo33byrO4Uu/tsAGPL
T0ol9GeQ6tuW7hcCXj8f6UOUVihCDswSHFpim/SC9VyTSww5pBm6FAhWjFtxv6jN
GykuoukGxQmLwnIFBq6AVmxJxD49Lo/xEokgXQxzsYTkUBc0/zuhI/Rn/DkWMRD1
8XK6b/OfDduWKx36ZVYxRZlIlQV2rSS3MUDmLd+ETUqV09b9/iYWysu7jjEJmPVr
a4x+eVEUGc/43hkcTTE0qapJP4XW3K58acTjieQMaMyVG9mzqcFOsG3Eu7QfrsgF
uX3Vw8y/DwHnvPCnc7rUiTMDkN7SWcUtiChxB5y9DllezMxeeA8PofGQmWAqI8o9
WFHpu2smA44KJUVr4HYeCPShCTmzmqPMb6eV64I16Hjwzpqq0VIoEKRha1JaICql
5t8EngMquSc5dhNY/gjBUDy3KBlA8LvH04ksptjM1fbZfnEAmdxGsEW9f9PabgDG
mcBYHewmZBlrQmz461XmP7mVY3TSkGdFCDs60XRLrM/gjn9N93vI1ExwKsBYKEjm
Omi6ZMDc+MR4OwvrWk3EkZoruw4NBK46ewe9il2n2I30+VxgIsA9YbPtyLItqLLD
uXNH2jfR+B6WWRnDJNmlSNzMN7su3RHleU8v/E+IjvFxBO2vrxLeJ+SDX3jegqVp
c4AyCwm1vcXb+co77Sofq+Pp8/PSvbd6hUzoR5STipGIj/KkV4SiIv1KCAMP3gsT
2t3eBIEzfM3/eFtK0ko6+x0O+2ogRSUFnvORehyklNq5Zeb5VHWRz2pxVuc4r5DD
SKUhrIklI6LmqIrU2JsHGVj5zQObfQYhT8Ts7OaT4Z1R/uaNXcO/z0NLatsRkLcP
zBXjvcny1dBxTRqQjeMVnnJCeFZcHi6XWbAfItbhL/RLFO9UH9oFlqhtZU32EARN
ZG5xBqt1gpfzV6q8ettVNFrNFbJcDFNWggAsz16GmpXrt8GYfGn/P9atLJ68LbuR
QPnOkzVgZomhzHP1X8rqHJpCJr7S2UYwBwK43uCLRPaABa9x7aXIYwW2C42eUjSW
d9jyirbAowx+HJ0QQzCkTncVo4/22opjR2AK5CYTEoJPSk4CKdXl8Iv9zNeqBU0A
SX2J/81NXPUP6Ep5GVwOUFnsOFd1hbu/J02bBd3R1hxkIfYAYnfrAQ4nCCaA4vP4
fEutbdo/mI32PCa50vKmLVvNQAEwwo3xIhYne6AGFsCimmunseWfelFjzei0B2z9
pZFbHZIVX5e8YseDuWa3S9j43FO7Ej7/3Vfr9bOZDywN6IFjcfAXpYU3c4dYkT22
D1gl4L5jAUuHSYJAptUzJGtFOjwuDvD7juQBEcz1AM9fTTAEjKHt3DV+6qqdzgp4
ZYRmqK43c8/bK5AIDGVzXYJ8CP/SSX/63fK8vKGCsyyuramWG3EdWkJgsXbbkKfx
9UySDI5AVqiocfNJnvz7wqM5pKEhvWJJFepZrKCZ98zQTnvG1dOFTzr2576d2uz8
RTaQID1rcxMGM7nFDkJNABkXenEjH1WRFKuz7XTLfSy0jT9N8eICjYRxJl7sNTDP
l0MnU+Tye8dnmzbd4xlH20bvZ9DSwdPpQ3blhMFtigKR/Tl8+XHuN+4XdKoehOP6
aCbvbKJ1QEcSxJ5GnPycp91qDsBQEQ39c+q6m8IA9opjculDrZW2hTXKf2kCCqrs
WEWBtkCnpqAZVCfYlBcRjpG3JkpOhDGoULQeWDtzR1UAZ6OR2WQneJdn7yVR9eRy
N96PL+/7UL6s/Ek+IODF41g1jNGBe27fjCjGvUudA+U7ErDGjwtHSViRAgt+VSdU
+DKqwLFiPRrJfndBDEq415mrmdH8H5casiugiRV4Bh7DZ3njp4+9LbpT63vmoAKe
z4tKF4iGqr3OiQNzd97dxihPs4yqjhtNlZXvqVlrMnekoRT6EkBN8XV7OKhNrhjk
Jc0e7Mr8ayEeu9mYyrBSVew0eWLaVV/RiEPxJRIDUeAbSaMomlulV96gfbrdPy45
L0Gq5Gwn2c0b2+WB1MY7kIERnJhAEdM3fUmrs3rPLk5pY9DmcEGCaUoKS+Q/G/0R
C32TdZ18xInH5AkReBvDfLuCizEmx7w5vh249nZuj6eHtx2RcCOkrshGqK5ClV/Y
UBowFPypb1FQ2aOgKWFXAIhOdyJTInPE2wE/ghb4ocb1igT2+Yd/vdDGdDCdXE63
aspNkntXwsARR1S/6cliwn6CToRxWGsuAzvZaJTSj9gXCIg8mkb/8CeqmgEUiwZD
ECQoV2Qh6SLLixs+sUpfltRUIDxSnj2DzdNfZbES/Klc9IPK4UAh03P4puDnidh6
sok3urzthqXcKYrCj52VNmdGCbHKqg14Y3w5iXDlzqrLOYB7mhTUTWSFKjTC5cn/
qkQWe2GIMRyRPSFJ2IMGM8rDaBEbk5/sFi68wZIMGyGHZoAPSi5Twarhn4kF7Zl4
ISXMT5gp6VqqKW33fy9G28jwl4hwKfCm9+2AiT56ZwnmdcfH0ZCnVX9NuaI06MKZ
0CdaHCDdktK6SHznpjJWoi0dsjQU7UbwexTZeWSic47Sqq5/NS8G4XWfUdF1KXfl
AD/wRXYuaQ0L8Huj9WciM6Xs7GyWgjzLuOq9KXlW2CbXHfVgmYAIJ55W2642PVij
P5vqFLaoRpH69gZzV1Jo7H3D6M1i2rdJrzZXBrS0GI5YldNimEE0KhLa0v5NwMha
lUWO6xRThBqLe8xtuUOQy9tzQYiUDT9bx8wK5RpI0hlYwSjDuFLREiLMl+kBv6M3
n/pnbJMA6oa0hEWUrNOkm3vUzYkr8lr++QBPYX0uXIskjN5rAKS59BBOEvOuR288
r/ME6FXXPspmBlagUREK2ez8P3aWjrl0IROtkf36zZZ890tEpBtY4FNuc7sBcAnp
8Y4mp1bruCnha4TsWSYZSNACFVbng+FVge7b+o8JUTxz/z31Sj6KwYQSc80WJbUq
3tliVzwyGOu8GUH1x77GrdLyB5SlVMiJdTNtjls/E0Me7eaF/XeVJXbi8aFz/30g
ZY2nFfjhAd6UCfIffbUJu6OZNqfw4O8t9kvWqtgD1uCowOIAte9v1C87bqMWczwT
Y4QnrU3114Z/rYeff9/TEKoZMAs5gZA1vhhDjya1iXE4zfLNeobNig1PuvWxMQEN
Ox50Sif3PNmO14+kKSN/8zxMYpAgiN/cpL0FZzBsX9yqdOg3CO/4j+BaZKKHbP/+
l52GdskEsOnUCSGeT9Kw3zCL6prTxDpdT9g+AB4q6+s45KMD5FQ2+LrO4xJPaaR7
7Ykwle273ktCO/v2R8qTh7Xy5AHG9Y5wVGL2TzENxI1Pvd5AZJYDMzbVGt+oZ2Ta
qmwmR2qskusZQfvxi0fSLI+ekYLSdW/ew0oB5til3Pzb2p2uYokDm12RS8DzV8of
ChJZtl+4wN4dK6T57vXAc/jeGr3Pfyrxd+yTpAx2efO7+dXfuRL/Sh6flaLziBCb
zCvuKi1XSy/gp/sZjI0Mh1llXQli33IMpAbVuaQonVC6nYpFAZMh+LCMHJnQot/I
ZWISno3KtZwgaH480EQaGg7E+7yFP8AI+h2WALCjr9Z+TRlbEmg0yIQ1zF6mQv9I
wG/YPphW8j510FURYXJBa723o+Stv/gCb585Bvp+fYfKY5vGlpajkyPtgVLKvcpA
bNHrAFbdqo9OE2r6YERSkzqXMjGUXhNjOqSYbhZtcpbhbaTc+AOg7NpaXX4A4gXK
3Y3bi3a+V4dS/5eqfFN0KFRDx3vJqNBnVBjlGg5glYPWNtWcsHxC4mwT+JgrK3Ur
jZspil459zW7g0/2zxNfADC+cooz4wjGxWOwYbgVyhDE7Z3iRYW1ssPfrAsn7KMc
p7DUTHph5wbwnX/6UyJUB+/iX7JFs4m/Dz3qPBLt+RIgDcYcRuYIQCubdTgOhgrb
46f7NarI8p00ZO2jYCo0hXKE+ElZu0VhuiMSYNNy+Lqk+g7CRRpgKvKqULqXF6Ce
FZfEoD+a0wm3cUsn/aTfWkLb0Bh5vHh6aIl71KZ6DXulgWQx31m5xNR1z2wYh5l8
jNJZN4PLjVjrntcAmxBOTCGfbckaJoCK+TPqDDNu7DtHQ/5V5N+g4qWHXaoUNVPH
w7TbY7Rd8yGI9RzmTfhDPtEEOrY8wkXPVtx9jjfw5U57M3faYBu2APymQd8KKDqv
Zd7TG7Vc8eqsFk7q6WJlrzQ4oiiAaHKVgtYwZB8d21A3T2RaVPaFZcMk/XWjuwAQ
ep0xY6OjH/LJvfJRHyXJoaXVt/9B449Dz9qBiItTIvfBkVw3fLsGNU1Et+hyNTZ9
OedPGD53x/B2u/AejrQg6KvlCxbguPtPMKXU9d5ExPdv2B9rVCdHtXND4VBzNSB3
Fxik2jXeK80yH4Tkv5wM1fdEmKMyKfBGLfEvp0Ffu6w8qIDpNYlLojGb2Wj+Ac/v
B+DzBh0DpciHceqRAgVKJyid20DxfVx/Y7FtPZ5sISy+OI8B4NbxGoO51j/uKe2s
uf4gHWlzWzIZN+CHBZecszHEBzfIRlHYqF57clNXQv5n737bWf2wLzh0c2Yd9Wv1
m2J62jQ8PjRBHo/hANL5C9BKDgVSMfOkFT8ZUf7yUNKmUfpqfp4+ZC+FJHFL6qeW
VM4u9glf9H4KgHb18vhqIhq/R624XXzSuwX/MNUFUx3DTT35KsZKudfE1M/TizHn
es8UqR7vWS/d1dCxXcD3KQJcEkBKkPHm4aOgrni0yVt7775ae3D3gzTuddAps1bx
whlt3GduByRTQSr/fUkFjujHTUNwZEAhGx1pCToer5cDnIBUS/9ZRbMwvcTN8HxS
YnYRDrYQr3yQmYN2sJUghBsqorvowzPPW9X+gsAIBozg3IQ466mUr6vOTn+ljLHH
P2zlghiDRQaKxxSKtU89BDBbMPx4Rcq+fstBGfnlxoQv8PiQBFPRazfI3IODcm+L
Ql026Z5cdE0UI3iuc73j6NiPORjqQ0/iaJk6wrRcBZCGu3WAD2/fnUi02mB/Y+X4
AYJiU7cgOsFiTuKubGrxSWLi4Ncft5CYhN8rcWiL8MKGPcim4wQRFYF0MwPiACvu
fCbtCLGdTqCTBsBaocbwFove1hefz38fBvjWzXzJZJiNmWo4bXSXPbsweKZ64exK
+KoQjTZwb6z+XKM1j19n8AqBu9AwcWk4KQCWzjk5nAq9ObzAJrsTQgR2nqmOw2lk
ShRcb/4J4cF5mVY4AAPd6V4aj+xw4enG9H6GQOsH2YGBqilyIV34kG2l1fbX/SAm
Lj721SZXLEbeBUt32RLCOrN8zKKWJjxpcOFHgzxc2yoVduKrLgsKd+fiwc6Ha9kC
ahirTFplOGqxIo2/1drX21brKXNq9xG26xQfnmpzg7messZ0NhBwFMoCF2s5o2Ch
4ekzttE6cNBzP8k60586VmGkTHFIjP9ktELD5i4yKCSWm+QQGTq3Nb+FXz23bas1
MEm5cZUxS81JBMlaVmErPHWenRsXTVj+4M0fd9T4cWHi1HcysTFdwnbhfku0MEEF
C0qSuenBiMDxHDyoL2bciXKL3JHzmweExDn4KotfaF65QFF8knUDci1zCIVjYYDS
o09RQsMtDnl70bzEg1K8S6rPUW/3b1itFA0dw+s3dyMJOf590H16NyTpdcdyBsyW
RR83Z9IrH4sOZV6EFqmQr9UUVJlaTLg78j9+daiHZDiJdWBc+/1SbXPxqZC4Aced
p9TiYPk2gsG2uhEE2aTvu9oT4aZAKi8KZjsLOKe1ys1V4VX8V8cPF3eYyE7JQR57
ohSMDubraRuc3khaCJ6tu+D6tjAcGhTwCP0webmRAZrDmxU8PU5dCJGAhA4zMeh/
6JwNcpPZkM7YXLWVNXV2sVFFRi6iiNthE5Das68BukrpvfKAPF2k/ri9Xxtch/Cg
RJnQjJsA26Pyr9A14JAxFMTq9UfSc4n+yske+VuN5gBMVJKSYL5LihxesSgLRPSd
jvS8XK/moOlYXIdtguFyDaX1LKgviHxW11v8ybsOwxoZq/rKddt09JMdBvAHx2gI
aLLlf01BETirGlwogA90oGNxNo5keS0PxmUwxryJaZhXQcqU31gDwtKaDkw+f+ko
65ZDwwLhCMYi8NfKjDg35iG0qPhZL/7gK08HKd1nP2pBTdhs9J9giQC4eVNh8RdW
ZN720ZHxwh6mbhHussAQtkCAVedHMqIrp7WAplXpB4y6vMPhzggbzpi2tC5xpqa3
xZe85TufkRBl7jNDb7eGZhSrm71Xy5a+wJWi8tvNEAzAkkicbzvkau2JAAv3UJle
+SHLCGx18B8WYrGgZkoH2lVsBeuRl9pbcNC7F0qr3xn36nw+abEYIH6Mo0tSGpK/
c7+8fOq8VjSOH3gqR3d30UbjsTrI6aBh0nd12si6b6GYvt/wGXismrQpH6IMD3uE
Pagtmutf7mY3wNZ1mLPz/dXVgh+j0yX9nNBfp8LSfeZJND9di3pr4rXz05C5gQZG
xlHg2oxt/Wn4Bdn9n4GPawLaoXVfOLzhkFayuxNuYP6hEhKtjRoeFpmAG9Mnl/+l
UmDNGZ4EDbjOc+H3fXmlhmQk6O/vj7qakoN1hNC+OsXRlrj3dYF1w7cJRV5Egw9o
6xu2p+4VU+GRk1hcL7EQZrgNpyJiRaizE7kPTv/3F8x7AoJOsZ7X7NVDYcvh0Pl5
2xY4KE2aleorXrSGgao+NzNJQsUuit1FmAgchsXUEMEQyv1nn7ElzClyW36N/wnS
1ygY0lDfVVyOiNA8Ss6Ezd23oWgg4BhB/nZaTwFemWTndXl9dWGtkqyghDQyJ0hk
GyEfcD2WrVRgJdLVz6bobWoSaxigzoF10GjLxqCiag63qvxxR+tIZgy9jVRjFWcW
dsEFtceQfk4zHFa5k4RUy4m8Z3uVbdCt2vNMkavu1mS8j0APN5RLHWqlZ52s0Rx3
/+0NjIwJgTFxsA4DDXwdSAgEW6BZ+aCWPAbpec3dXQCgw3itctkduac0qdoUeYVm
RwsOAFiY3CQSQkGob4yRbxQz57vc9dthCqWEH8YQ/46zFzt+17z2XuXzd4y54CUQ
aDVOIClB3bY7/qEVIBupaIL5sDfD3+2lOFmJUZAE4q+w8Qq2KLFJ7UBFKltW+OKm
aK2AnlDJ43HlSd5ynlQDB41ctqZ5laNxWtXF5QcgRQYefhy/AbAikffQDAaUPqf0
Xj+me9Kf5/NsZ+c79z5/+MTAYj1z7spHJNJ4E8IKIJ7CKX7wyJ15qPKw420OUMDT
IwJwZ2zp4I+WDZYdJwAGABL/uXoH9IIgjhVQh8UnxM3sCSjnJDDEyckq+BKoPCTt
0HXPT2fvlnB3z6Fp8qnRtvsZtOwYQueCmWoghxPhAxgDSDH1SE3Vf7N5yQgRLoJ/
CzVfBw9U/5IvdMWagwgNvKvvXuCYquEAwu6jP7OEm0auaiIOaQLB285yQ7D7HXEt
GpjLmA8AEt4StSRL49/w5lhI9/ntZ336GhJT+EipN1JEkkt3+XAHFxIo3YZawMyT
809y4t97nYR2cN7ck5YnnpvXx6zPVvvbahf/QLxM6hljhBiDczelFqEy1sE+0ym9
9X8JB5nsLI6jcio0NWyWUUJkvoIN7w3MJbwtjldl0FkJG6S4tGsEede1zO8LxedH
BhiOkt+aLBy9qOBxNe8SlPH7vUeFUE5qL8xBCwdh7MAckuOHJtjqQi4t/nhvxzQK
7yN4ZyoH1rxn2zSt0lIuGpDXzvQcTzkCZqoudLFAC7RWL8mDjX3n8cqUCEbdPrC2
cR+Cd+7Idegd78nhZiqJxKtkU/R+pR+XpW6HEh3mKh0194gYVg/N5MdJMP8HuGSb
i4CwaBnZvSSnDpDOFm6RvmI3HsYIbQjFvPQHHzd9wW0/mAA4+BH1UvTJHUIwmWxL
6iCoYA/04sFv9PUqCwwcZTb5Ik+le7TW1RMcHoOra4HTC5Lr7nTnYKl/EqfSFuai
HjdDCxB1CW7uFMSWJ4PUwaqdWx7AWFpfIB2gNznFw1jpMq2O1GFX3tf2aOFSC0iC
tf8GXql97TKSyDLKBifkVpk+MXvo9xF5GwVGSj01p4UoKbbzH6ckpfUp8OgzZ4lb
o0NC2uORmRMgRjioQwdT09zBE4eT9Sv9BwVWaEGQJ8I3cGqIVWG8KEfStOgMFCst
Waom7VClIIYyGfN6U+ygTY2alNJ8pj9vAlLBAra7c4lSSQ+N6d99ZjNJk4iecc3E
dy/kDvM/nybT3K4Ymar0g4YnvlORcqITw3KFzy38MJaUFej90WnwcGnjlBYs9Zen
Yktt5WPe0pYI+NEJFYZKTHPR8WiRI3SqgUCwTED7NA1T5kIX1hTOosFrY+HCARMM
xiT/Ng0MQLhhcVkzMjGB8AXujdiFpJpTOBmvAczIwiH0KiG4OTqPPrv8Y9GQiinW
BLxKLlRnuebw/bW3CuWtCMJQTx7sYt4Woad+Sv7iwPsTOZMdgdF8+RFc+VB/ksZ2
Qd4kHdCYuFLbinpHRpamuGqIvw8jYhZvkIzDlfm8PqrCP966kDbxVdiqh7dN+6Yy
blf7uVpshw8neYI4rWZw6VLQLqk7cbwI+AeBDsg59Ag4jAqmdah0bORZFNP2Q/WZ
JASccfYlxhY+prG5RYl8gn+NzcYhOpabLPp+Co8EkwmOIgF6cWE/LCYTJl8HhhZ9
Gufmga++lg3AQvHjGhU8sld6BMV9Mdot5pN7+fDT+uJgqRhpe8A5PpVB4bA6Unza
+0lWQ3OEUaDB71AlqXEQ34xTXVBZB3oASIILzo5ns4KCA9zxXV6wkR2btZIwCwMw
aWC0X9A79OyzNxJGqbUYBfgeYvTPws3FuGk1MnWriT7RH2sHBWfValxPDjn7O0Kf
aH3uy9t0BloFR6L3W31uPIY7doG7iGtoKG62aeHEJIKzWhi6MvJGwdQOoR6q2Rcb
rgryA0uOpeIen8FTWj6Yf0Y5dZcKlZ7BG96NqWzgdxlvSpdJw1Mn3IEdsS5kOrkC
BfjqUNuZRlDi+5L/BZOzocVC5cuJcWzVqQvrXPMxe08duOAoBvGI5IEWLaK6FPCp
I4Mjb6uKpO14smrQ12gOaoPpt5jukIZWwvfaeRdflxD/4LDkobJ0TVbxCLfVblsc
spD870wRilxUBFfwvdBQ/GjCxFpbKzFM3823ZFE6KIsh8O0QL4kEWcLoZjMTw3DG
oBXvoYGESLNN/8TxL5m+TiXkt2ab+kiTgt/pdzBIwf+VmVhymVAs0asoMtEjLMVO
FbnBrOiIaASGI/NFRQdTPAKhXnJzwDATX/NKo1Dag4vmXjXQ+k8sUFTSizUnvwIG
xMp1ko8wAmuDbuo9lmSk+Px4K4/nWxta3DfRmCyRbHys1BqCaMcIEZ7QI3pTlm9d
XyhNNybev70jIBCfE1PeWZI+I5R6x9+sucpninDd2Zf7FWA41ybkRNImsErmYfm0
jR3WjjPbavM21BZzlhf97VrKY3rSGiiwNcglBb71k+crQq/yf+PHclqY1ZZWG6Dv
x70NLMjOmFGNy5uW+U4YcdgYuqukOVb9vldHuRY4YyZQa+GX2GBcnIPC8IrzztZB
ZglNcSRJHhdBcp5yvb2VR6/QcfgaEurlSgFWW1Zdv9x/9h1ljexbn1AQofWUFjME
dfDzdawIACRFUUJ9NfpFOmtwSRrcTJZWNpl2aM85xIJgsjsIopHQwAY+DwquOnOf
K/O34Hih6yPu9WE6VtBidfKWOC+q4ZZU8KgMiUD1xzPBgsZpbUevwpYpkpUJj4oM
96oUm7SaYpGTOLcasABeneQsTVfT/UbxO2tIHRQVyicezMT1Tnr9uoKHmkDoyG/Q
ycU/ZP2sgr1Q8gPg9d8TWQXqw0yksPL1UCt8/4Kiy+gxQ1nVfg3UJbuHFJfbMFCv
fxKdm9KoQmoYol4Ci4EFGox9TG3XY8PWzkAEk82NzzIvKTsiabAE4DyxBr0aNTMn
VKULLxu8qSspws4rvC/EiJ0QNpkVCAB7BQ1DOUvMSYz6sEg434UiXUCXvYm877vi
nB0q4/S6Nxz4HuI+uKemzAcChYpy1RPkNfKNofIxYEiv7PZR2iEXgviZsHTB9b1v
c76Cf2bZhAPxOsgEGbepEsewJfZNIlCKfC2rMOdYt7K7oAat4g+e/sslOV4kF5+o
rsz/KZ19DwK3vZOzSZrAtUhxcxJAiSsOWs0R7mHSGrtOa5M/Y947YL09PsuwKZiL
eyhjKbeSDX9oay3j3yePLcIXrkb0vbk6tm0BasIY3inlI3fLmwjNXssVdsj2td/3
L8BNhl9jT7VYHga8dVFHHfSMA209BrOsUk/r7KEtPpUUJyGfEhS0NYgdpFqtJ6F1
7rP9Ia+n/wYcz7dsP5dP9VoHqCbjioCxx7i/E69+g16/Q7PgQ4naGdBZujb/7Kqp
K5yLPJJm3z1Ht9Iejpb/1rx0RL5k/A8PCPkzbNClFw+6o2Yn+Yyq1of1dZAGNVVS
HgoFSdmFpc4wqhWAPR3wCiUENDc2uXEXqv0J42mlAofhR5ftQt3Z1aNXXJVZ/8Bq
DQClwoFwMpjLOs9u3HIy9fjpFC/VV9IRLFu7ek+Ux7mBXk2WMsE9pf/yLsrSGnns
FD22aiqmq1x34Qf9rr2YhXbAzYGFsP3rfE8EywvoKZBj2PPs5HZrCtqfp36vZynq
uF1Q5LsOt45fGgKAITWthq3/nsdJT/2qRC4NDvpWKoQvXYui9gescwV29ZuC1y09
G4sBvodxXj2oNkwRFQbvSppj2g26cgcq3qMUV2m0H97QDmoWIGf4P4sVPg4oLag6
7ID/fO/FvN8NKhXWoaosfDjyNWgmvNbwD0nLl5PJXweaJS65JzbDyTN1FkO+HMOO
12RH6UfSrV+Tpbe9ca2bONhPKxJ4phvGQSnMoDkJWXY7A/af0xpHyGHK5Vx3Ua9y
hYoGNHSmOu/OdaUkAkTawL36RzTFTTL/Rc28/Vq/bbe6UYad578b4ieycEoRXpWG
U7rEfvNgBdWLkVLlwuqB+vHeMBFZIAapC0NjcRkvVL7WR3Z6Y9IbgvqK7JiWW2z1
fyDj8aGenOWWbyARPS6jzpTTkzO5aWG2t/Qz+vAXNQRqCeWYmTLejXb2OMY9UWDu
Y4aaHwVzCSFtlbcCD2C7XKUwOIeWMJ040By+bustZbci0dsUxEDi0U87QEL2nFA1
kPoObLT1e7QQ7DGEwpJNt/l78DpY7iqr2pFstva1yDKLnfBBHev0G4pMtT3dzjo5
+Jy3SOCBHn9hHqNg0a5ocpW7RyxqW40IGh7FEImdE1SCTS4BOxgaU9kkdB0jaDBL
Z7XiYqujVDEo0tFb2UlDzxKvHSw7clBMUv57TcaPz5Xkqgy91SAGvwtJV5aRfLvV
uHeoBkl775HpVCkKUzS1aEdA/B8nxJJvh9jK5E77VJUvP95cNXpYbxgVvIyIw6h4
svujcKQUGtWT5rXB0aC7dWzV7XKI0TA0Vr9sTEp2K4ptwcHap7uCBZIP2IVNVkQx
cZcAgbSL4ymi/jYMa5RO7Is9Besgz3t1CStaH4YkuEhW/L8c0OGUllM5khWhm+cf
brB6HuZ4MHiAfdDJp/GSDVAE9fZVeeZ4LPNazSioxhHoTlhIW0PGOcn9V51/rOiA
U2VGyQfc6B81QmCanHOC2fMPecgNRH1nI8eDNHPqiiEoYnrbZJPz2gE1Pq5x7fyr
WKrIUBi4tN95eBCKX4miNBb2k0XtAfQuE3R5BjXM4qOTWTPB87XSTHgwt7xjnH8T
r7hyCtZdsp/4p7maI0F6kva6T5zlHmRy59A5S5NNcAD8ldF1ZU4zQ3G5F95xZjMV
ZBS/gxCnjeY7cdR2+RYdB+5IALNlIzQ7m8c3K2sPYbLDibPO/M8h+LhuA8KC3cMu
jMOk9csMI8eXCrVjx/Iri3SgneCTK5jxcyVhKBIT/PKKqenV+lqnSCY8rce41ZET
J+TomB1aWdQPv0iaI+7E19qgoIEPqaBJfio8Q6E+5RLTRJTl3XmooQPdMGfkwIh0
KqAkH32AafBDcKMrtc6V6I6ZY+yyq2sGylZE2Vkywd4xRAX/cP58y2GwO+QS0ta4
ZqrPgo6pnN+Gt9MoQhLK4BZvoOVYyqy6iIf/MYwEFrBVmtiafNz2dZT7jsElePpH
mqbWlpuP+V8FNbWO9NxURMdsAXJ2x/1Hz37+22tMEpt8cR3zOCNQR2DprKzLwSYs
LoIxfBOK+JB14jpZAuXWeko12JEet7QfWxPHPSK26sjxTVGoYq7/E/cjf/2+dkyc
CUgZbv20yaRpGDr/bpOQy725zEriBaQo3ysgkUDiad7tR1VSt/rii9D0pFXRmmZi
nC5a8b4mtgXRV9lxT4jProwJv5r32YbbRNSZWFfh7PGIaXukQC6xuM8AOm/IBbg1
zfUwvdSE8CoqHF1HXGJV7YHIeIqHFFltE40CVZPHVeZyrCP0jKiI1TMgO4vdNMbu
/wOl3cFjVDERezLBxqnQ6+svUjzmPfRlI9hkmoRnR+hEAJfc3YTKS4W20tEmwiSE
nFFfDpIi+R99MVgJ/Zm1RLskJ9tNY8gZPV7obgZeFYalqmoVuUJaVTfQMH4/SsAA
Iv6VfVc1xzasOA/ZjvuPmY8sh3j5PbnlISf/TS3dbuha5l6lSPbY0WMhrD8wSpI9
jrMGDKJ/KjcDPpDczZVVxlEsrBFp2U6AgkLN+v1egezpFH4ZBQ9qHwg86BZF3l8z
4HtaOGFnzF+gqcLW0JJqm7eiJ4WVZ3LTbbeX0IEY5x4rOnlbCQW+X4yxcqdrwdBQ
+KQbYItacqYhuaTC7llqCmFqk+PoeXq9ean2+Ta/RGmFVw8SQT0AeKY9fyxnB5aQ
RgfqaUPlOFYm6iwRvp7wst7ouJjVRDttTUZukTczecnxDMAZ7K37qtS312pyJAyp
AlGB6Z+lSGyNBKcRpQMFJ3C+lr85yT6IfYmreMYS9aZf2iaxtU8ucWeW8T4BpImr
2dIetB4ov+ZKMVj7PLqdcYmg4vYeIixd+jdzpotp5akpyu3PrxcV/gZG0lxaQBNk
x4L/Bj8OwufgAFD85W0G3zfonSYH8wv4BhkW5bRvpgzTU80ZDpql81YUgzWo9eC0
jnUZ/RJWW6bJkyq5G+zGZqjXtTnxJwQh2yHRbcXYutnNgkbEh6kzfViuj7/y1l7P
ViSYw6xecvzyaxelQrv3MM9fPySN237KTbRamx3Dc7MRxxsWBqqTM1GN04TodYvA
aehEpHojo0EYyO/YF0QmVSsMZ9aePsgkgZlu85lMjMr4d9lyFDb++qZVIhIiSr1P
a+pS4trrM/iuEBtLBiO/OHt+RHyyufZ3z1dwOubDF1dF3hz2/42zrj4DbOAbiKK7
2z4IWthtxRpYsBeA0jkJPGkzafVytsaOxMx73g2wMQZ8DUAgW0PWSiA2ff+LZD+V
CWuupEs7vUEZ8yledLVLLIKwcIsN7u+VEkIvKN9k5DE/1aB13CGT3uQ5EPcS8pPF
AUzW4wUlLqttaFnxyiuj1NtG/6l0LrsnJolW0A0rPTCjhbyS8dDX7eYAqDhrBMHF
pP+iQ0e6O/jGvKoUJcqNREVkA2vS1IS1GxTGYwvpRqhlgD6wmxN7dZDxEEqZ+2gr
2pKQkBgbnqEn+Rqn6ab98faSHHfk/EqwlxFVLWaCcRWg5h/tx96xLAi7XFDNoMhy
G/G8qfQqEertgiTDqpiUlvOgkGwzrhe+QENw4zMYZDi/S0K2wdKpGwIG029Mn6qw
KGPJe7Q5e/8mPW0SbUUfsiZp+hgRf7c7QJeto4vjob+kNDw9DgX95+BSeg0kSPj4
OhcCLzb6Lkpbsr19jsZ8Ly8qAqNY9cOTm/esVU+YyJpf+7pfYRA7Kociqa1bzXY0
a/nE99hx/Gv81diCM4at+t1dMfc+lG9G2TLOJRBPG3zl2li6RHU3vJqZx15dPIyF
LB86YpGnHEM6cgPudO5M3lC11FBXMJOD/Rk7l3zbWiSRZ/a7vxOHivSXJrSO+gDT
totCPdfmrb74IDKvSePGA4VBQlIao4aHiMD+TQzdJECveX1le8WYeXd+x7eotT/J
cGK6CHueRuRlF3ML5QNYscr+KBLnaozSNx4Hxb6Z0vAJJxnnR/OVwQaX/433gTfa
MyWUXNwWOFH02+AoQ1LSL/Tanw/KLCK4A0szKRlOpBffUS2vjx76Y9a1ewGO/iPR
k28Xd6lrG6LUTNuCpK9Uynf3t/M7K4JSaaUjhqH13iE92BebdatzmyDtRT3KiRBE
q6maUFDZ/USXvofJ/M4Q8E0iH34EdJcyYPyBDyMl0t8SMFpPYSXTC84O9KpoZKg+
0cbH8kkoFa2SLOgomXeThASkf00WjFOibOeHKyZyRTHMV8+HoUccpc3O6Lt9+y7k
1y0pb3XF4UrqCHzkB9glHqRHkq8hehcprEhgQUmfPjBpHvBy+lbe99CgGlzMG6HT
+WLbJqstfXe4gVtAWfOsA5rttO06YYmOXhuq6PaBTOvJK2kW6z3Bs4Y4DjZlKO4L
oUpWm8ucfySW6PKx2KWdfq5IWECjQ6oSpWdpWXyCrSdfVeyvYFcpb+03j4HQxO4w
M66pRfTqyElgl+C8/mX49PApwVV87sWBQVy2SVdvsqJzgPhKvwz7wVJsoWxHMcpI
WLV6K81cz5SN6ZLelkXZnxuPTBbYme4GaIkW1jYgxPCTbGbGhV7nHVHffSrtbg4l
PuwintpQcL8c5CQfBh8WRWR77HDwiFhOmK1Q66/Hf0QkH/6rJy9bjCcR5YsEolLU
RlZKyDoX4aciDoQcLkvx+uKxXfzCu9fc45iKvisrfXNcOspyXwPEa9oRuKcRFgsS
Ah7c10YRSOrBnEmDxNlUMN+lXqBBVOmj4JKjK7n9XH3JVgc8lhoK66OA1Ru5AsQC
XcgJSmSgFUsviU04NTUgvbB3bUteeoM2Dz5QtArA0PY9C5P6yvUBwCk7Jsd3lgSD
448qEXI/ORLqCn0/+vKnm6V54IrbNImVGyZ08LnI4eobo2ZRxztMoQ44Lgz39hJH
H4pqR0Cv4s140CibycZ3Qocwm2qHyJO3ijmyUrIOPsGr677/Qae+UXD3IOBoF67D
Jr8cmbyakjOp+2Rbmn7j9CDhqlh14vVT7Xs0Aav1EgA9tTkiNp3RFJrTxwle7TQc
iJKzkvZghWn2NQ9JVTpAF+Cmza8g7u6zEBGc8T9bybyyujOUSisQhDgkpOhd4Gui
Vaw6gLCClspuxqq69yvM0ORT0YGh9WBcD2+dYjnVmjagJO/rcNnarMfCDLBtk75U
/SJZYvm+YtlMIHJyP6QQxF8B8ibbx8YVJCUoxgWi8k1xc6LHtutqoull4PuEWy5z
mjF7e7tzE+sO1yNXl5U6YJOkH7H1uiOViciQNXPHlHTIUf7qtG/CwdaghdToYKD5
FCJ5xqum/fWlsyUO7mXSA8G885jOcK0V8iwDTKJeru0ILlohbKRkA7SA2y6ULGg8
6HMWn86ZWzaWvei+A1W9vA66aLKSQh0ouKA4WWXYWQcz9Qtpe0Ht6KgOD90kLb6r
eTNFORxbFK0K6girj3QXouk5fYyYsjqchq97b/4w3TxXg4nhpQ5Ln2WTegKdw/zC
8r9loliDhnU7Y6R/hSJbdV7ZiXnSmwHQzsIen11N+2JV4JmoDm2Uxq5oTTBW2NrS
xqY4MGwu2NhCtfhzcHofOrV6jhNpOvp/7lNC61TeXPJZb2gpyCVNmQ4p8uwnphCk
55ESG6Ogtw1jqPQ8tw2KUWDN+x0oWd64Czk6A38QI8j23/lXbJUxPIkidiBULXq4
oZoRKORCSCxN1reev31Su4mDYL0dkwowFbQzLsJed3TXXlHaIYvSD7G1xXcpZ2RM
PS+4AYCd9ERruPxyCjKcctzJeAUXDjVxN/7n2JdmhGt99nls8Qmbk0GYYV7l3oNl
4iVLCm/+d1liq7zJC5y8LT4Io9jNeFzOJJUAofNott7VCHHKV0hXehCxO7IHbzGV
Tf+BmS/7TS+Drju5JwLorSJ4u1jaQgDlcC2xgcu6jHjV1w37/kE/1OnSvJw7L5bt
d7rRKQ2iT3Wxa9zzSlClMhKiXTYvjaeCGmJ6i+JoVLH/cCB9d0MPS/cIdkXIGRic
gYIh3Z+oJLhVuXuxl/m0WJvvdeK+a7+1atTb44aKOrVsnGGgBeuBQPvOsmIBv9Bu
idJnVqqo2uh2v/kHvsrvqErfCRwv6go8UytRF6BvVqlbOPVfnFfIM9WHVEKlGIst
AGsoaXTc/YI7Jed9CDPIzyhesv97ncbSMqKdddDzd/03t/inHDJcb8EUjGvidarg
3akVGnMe1eXLlLbbT/nle9Sm3XWIfTrrDeTZPD8EIgJ4ELDwopLcYG96ouIw7RFB
6qJvxuBXYi1UGc1kBUrV9PPO/2W8ACWASC0JrnRYQFnoQ1QqYxzreSP6K1pYxUyk
e1fPA+12EtpF1kxJDk0nTKUSd4J6mvCpy4EeLPPPLFgZsw0Ddwf+71+tdElssVe6
nXyYvduK18ap58qiXYc0siZIjdYfWgqJn/C+DKGoxyAX7QPgAym33TskivSWleyY
azrgj9aavvKJS6V0OmQbhWlI8wZxmVedAx1+SOtQ9s5sWX1d7SWRrg7f/47SEWVL
gqiJ58iqFHpZp92xIhdAdBL3gpzo5QlToRjTH7AO4x42EmIzhNMhUiPX9eZa5uEY
Ca8BZQaHSx7ptazoy9JVZR3B3kEDCdqhw3ot26vh/cq4b+zi1kGl/yaCrTiIcGC2
7jMRSQURUQeRKt8VE44OgRkdYeuT922RYfdeAQZEb31f6r90c61P9qnOFVqq1R8G
cW6EPD9H05dkul+QM6yWqpLh0GWzVpfInalBUZXopQ17WZWAtAQPLgchWg5/MaAC
rHsdeXgex6kjqkfzGbZkOOLvNCWBobGfTjjwKdp2VAMVQH1VlBznEFof7QZ2nBdk
PfDfOaDa5vrkgQ3+Sjg4FZOh2sdi11OLEfHw03oQl7beWMHYd/Gphqm+wq3RRGJv
vQh2eK6JSzSsrJtk4FcxapbAvklJQ08K634+4nFH0U0FoOvBVAJWtl590eKR4Dui
SjUiBpNcwzSyE+BJAB7xXHX/3vodSnvdC3Re4/+khKGGOoX+5pkGnCX3QFTf1n3d
Zidb1or7VnR1AOT7OyvcHXzjxb/MnB1TLYzzBgt/A8o+vC8nS0m8HV7j1NgyzB5H
L9AQwjgpqQMolR2itwguMAF8v4g7LM1DavmnYlUZjRC8xeRwaBDPu502qJtKj9/o
Slf6i1uWuIgng1MD9JxE6/OsUm+t6/wFWPdAGaAh2gykXRHKAWKhy7ZU1sfaHxEu
vVK7/nyBkAVdkd2lxj/b3RCiLOvy7fxQiBdo0BHhqG6YYl9uPenlRwOxDQ8/+feU
7mm7dKd8bmodkDxJdTPWXRPDnY/0D0CzzupL5xbMQRknPBWfi5WZqqI7yFoQW1AO
ZwHMgSrF1H7DRep5AKXWJU/XfJErhFfaBtKG946zU8NyPNSdCMNPg5Tjr/Cs2z6c
AYovzx/GZrNLNuxGcoclHM/DMOJUkEue6ExiwV06vHdZSoDb1VXWhCCePF1N7Mun
YCZxQNjAEmQKCqqr+uqOnAXAV6GERhlrxn7F4Z25zhZI2n0Tv3xYHPmMNsDqVP0R
Ksxeo3tYLZJv8d9tL09z7yAI53YNjR1DKm5Lq+hFafWC1bd5l/4AKhQngiZW7eCf
jHCel4zcKnAmMfQFYBUDfLOSplw8dePauanhCiv6AMPrKg7nZTzsN1hU+cKtht0E
gdN4C2ruLYBcunCF+TWhVGKjIKLjvOG8/XQjw8Whedgj3s7dnMc94SMsVrtoFTn5
o+W/E7+Vkfad3JyQ2Rn71N6feR1VdSmkcBFlMyH7yLrT25CdcOthzhVJvRwAqK+y
ECOr8MqPuoL8Y0UPy43euSHdFUFTVNjZrxywvfJ7ClLbL+cFhV/+XQSZjt78jH7S
N+2fTmW5dhRWF0l0uxYpPTdo+Ii//3cR/DLNucAsu3eNQrkwKPkv5YmY7MuiRa4y
ekrU78/HkukjvS67VL0czJLTe4yUB8gr7VkW9fuc01MpeCNyeTFhgmpo18ciivL4
ufBnxydDjjkRC+xfybRZT6Ffg/bTjjyMwWKQy4O0WSxw9zVczcNCGA31OZVA/IQe
0yl7MD44hCI5SM46ufT0luUcm2kFVLJ5nynr3qdeaCHu7tPm7H9caefA9BV22f40
6IDa3cT/cSwDbFSZGcWUQz/zkF5LvjRLRtk3ARaNKJhfH3OZiUDkbEtxruh26tjT
tfOXJ4hcaMLk6q1nkIkZXNn3AMQ31GrCwkmD+HvDriRE+7jT3gVZA9INAzywEbol
9aZAK1v4GXVG0ncG1dgXL+Aetcu7DTayafDKBuxaw+OlIWWhMGTHxjLNK4wevC8s
0HLZ8x37CkAMRpndC/1zy+JlMHYirrR5dqXqFHzzJ4KvHkh3t79HfaZG4/+3Gb2H
7QWIUBtDWmw/aaHMaCtk9yE/HkYvv8+bVhcWKhXGslhGQP7sEHPYSe4dWvspUUTn
fNUKyqn3HiMFMzHZoo1VgVarrrnpHNWLQ7esfZNEsRWTmLY02cYv+nKerbnIuddq
DymglJ/3DNdaJArGF7Cxz5YEFTEwpeQLlqDb1tKYC3/bBJv3Z6SLVYIrarx+7Up9
XbFC4t0c1EhOWJN3wJefvfIzDczIJ4819tRkyJ20LjhippN2x7wjBGH8xZ2s+ojg
Sct7w/TVkepdb89t5bq8i6KCkiZi1f/M5wS38txJXjpdD3eMHDFoS9E075eXc3DE
fWz1B78J0PYC9twQoOgqA8XKORVkrq/KsdfHULuUZzEkTDoo6vcPkq/zPdKMBQEw
jsBE7wbOUSaemaa8pDGffk8VDPHM3EKkC6BfON88AQKieuoOQU78c6qSCdqUO7ZL
9GCo0vvkSktbb2ul6UdDPM26NB0gjZrC+PBHaA1BxKraPmkVGuDaKiJpAOV+faCv
1CExGLv/NxGQeVKRcLyekFFXg6SgqYKjczkp7y2F0TzsmoeD+yI9R42Yn6cp9aH+
BplGwjXVgjBLmC3mYgF+kFnacRI+FkW/c3vHdrludi81G8W+Fc46HT7UX9sXww/a
TMautEQ/IvD2LM9PA13kv7zgZjfmcEgcQarUUMV0vMfRIwpXzkpsZT7isOGSsVQn
DXzVdw/51IqbxQ7H6yrZimOxEs60lSDhXAw9gey88VL/E9i5a8cff/hkuGPwwnVW
nuFv5i9RBR+ZCxJ9CKoaeace7Exb0mLOezI+UdUAxqjezJfQbKicxW4ZoOyy2n8/
d/EP8UY7b+1sfAsplY3EXXjuKfPPaMFVrqlbOSkZIshEybY5Yszi2VV0WZ2JojpQ
InrSXhYm1yNPlUw4hJv0QFt6yIcSvSmw8sbH07L3hpNBkeFJ88/fpTRNtv/Gkfke
q/WNi+yT1W1mp/1ObQzif+SU+3MoM0EM+JWoa9BXp2HCSgfL/egIQZ9kAaQFogIN
lE3d+/il+1bViXP7tD1I1jhqhxc9G05t09xpZmZ7uPYBykLadh/LUkDYg5/MuBP8
k1AU1xroNG4mp7y5CnJqDsBzvN2UtOaqFjxCtUrGwbNaG/SD9qgQlLUrZKbzOhED
8xhaAiaj3kOUJmxz+CGVskrZFdvaL6E3DDwA7kuUCWdjGJasJ4F6SYjoN/2pXIom
LSG2M0EiLEr1LBX6IAoakrCKQ4FMmO4oRTHdBkXecz2lqBtwMig06MLwJ47Lw+9y
2VkR9A9miI1WhR0A16OZV/twWCQwYBsArIxKbusRakOIu1qTV2juDypKC1p0rlPS
6SODgMfHH/sZJtJ0PfN6qHbesGjzgXeHnGxnzIb9uGPLRVHvUt9qcnZuknnorrsY
kRYkJdtra0apoJn3Om29Y/oF+IUuZelxNDT9PhOmnsREggTwSjZv1o6F9Aq7VEgc
qsIwY6pTz2Dm3dojhjD/gSVR4h3GLBLKozd8RL7KeU9vEpwj3v1bnelGUJqRYzEo
G25ZZ7P+gUU2sjNvMLsTGLg1OVvc1jl++xFjzw5Pqgj/dSovYgah5ssU5/OFFuYn
j9Hc+woBKyaC3nd223K9AuXaeGPHaFaWgmGlgv+dxXdZAvCR0gtVcH2xXtvq7HAv
VWHstp1uBgRGO77eM5AoS5ghmYqV3YIdLuKMibE5E4NY2Oblgo0ZMEBlWuUSwXcA
WX3GDIFdHRtVLnvpHYY1g0U10GB3CS9kKgIcT6XBKdIqO8UOpIUZHEkbrnp/1ivA
w/lTkloc3M9DQeYtaY+dY4mTTvfC5Oc0voblhcjrjMMk0NFHNTNCPUlU5Es+zEal
VapPgjCqH5RKW3B3IG9zqxxQP5LX3AW8+qDUwTZAZfpqBze3FWHbjpac54czSZV/
8w120M02XCT3BRw24+AzNwX5GLh1WE2fCGFo3vu/y/O56XZcoVKw5B+ezF0lxQRB
xVzuckkMhcOsP+D/kkvynyigiVenJoUGbDw8PzQ0ToB4WboZqgK+naZG8iPLjJF+
OkWDsy650tOJ6SkIN3CM/8/QgGext0hYgB09wBG5CI9cm3CAER/gQMtv1QwjS4EY
m7I5zWVju4HNfs4pIE3oWsJuQvIMncrCxp4oXtBxfsWsrPOONbDdyc2soHjc4jkC
uzSO6DGHhCyvakb7qqB3bvNh1J6D/we8oDn/GFhUeLfHIhgdkgdRGKavcHGA/POC
eGJHJNL0ssnk7AoGQRl+ov2sS7jxzgFNER9dMNr9lniE020u0iM4wkR2slsX/ddB
jgVl34AA/odLpafnPmVnwmKq7L8vhhxiOrdLih9M/P0zHGsRQ+DQgCiSDZ9j+Blh
yWAQ4eVo655tta8zdhwIJRXkKwiI0nZZgnj2A2S2vFtQhHFvzUzKxfaRS+harVXz
bR0iPGol8QwSuFz6yuM2qFnaTShpcS7ol63/ZJk9HvwtkjZ0WxX5alcUszAsal6h
e/7U/quy+51jy5UHBLc+zgEZxUCHJTejY3NlLHbnPhaPEO9LhFJGmo7nCfUhsC62
8Qzy0O4+FGqsWnmr31xKk1LjfnyXOqyCjAirmKqvXcOIvzLsBxGo51aFtWCa88ta
Sjsmsp7HCqBy9L8DOcjkMlRibweVDesGyCEjN6equoSgvW/vAx7b3v5dfQe7OYC9
zCGVD75ZEynDjCOJbtFZMI/kcaa2UKSR0V+Rreqkd0ZyBSoZp5oKtKKTy/33yLIo
0Ja18CkpRn/WpusrIICMoVF9Uqo0wbMShRhYDEuk4+wgwrTRpT9KQDy4bkcpnfDv
YqPmsnpIXuZcpFERNd0Yspdhp4hy0oE6DxqFMFDCcBzLzzDpNH/4Rirmb3U8aNPX
jbLRJIhN9yTmcMHKfT06d5dWuA4aaCSF2jbyUDY5FWbkebj23gGo4nwUdznAkBtu
QERQJ9M61xafC7uti7riU86xGxKck1CmunpVw7pQz7O5gj9lRSs0kYT0mPG/QzWv
MLn7oojwx5IvRj5AWls1FkNPulnBwWOm1CeYveMtKgz9PkRzHB3VRGkwFhw4Oz07
Mbg9LjGOu9tsCv6jZ+/VnPNQXlgzqkGclRJTvVpq7JnKdsWmNYaMRaWy4ZYPrs9I
SeGOP38P9r1k7dR+9hnxFpM3uESaBPzeXs2mINR0+irLobcBF1RciNa/GmqTyVAe
CiM2WNZW7Z36A3iI3aVAOLhthNYCPBwNVHxMvhT7KGPA/sPkhA12VP+JO3DLYoj/
c/+vm6etLd5eaSE1544LCClgHE0KxSj2Uw2yYUe9lFBQab9bhiCbOkbWv4w+xmAl
Z4lyi8pRuqoD6JKb7X8qhIhwilUZdv4S1o82YeTdR1QLT2nlXXY2TFLTAdfNG/bD
bwpJltZTyj3h9UMu0PaAMZtlw7TTBHPzoS41y8vPja4lH+Lbz06ysh8mjuwzMUOO
m6yzqLW7btJRneddnxDfsMbqOul+BpVE5kND3C/CUzzd/oJjw2kLg7jtizuYRkNc
9MV7FGITyQn6KysmSdFtGx3bKGgwRR8F2tmrQb9pHyz7OvdlerBrcW7YcHPiFQ6K
ozRNimOmvt2hwoDRRgaFFM2Z+mnjMk63wR6dWboPx7YrWrSIL2BI05UBsKI4Cs5f
24L5Iw/HuguX6qCLpAWukjSjl6IfMVauO+ga5agMyQV+CoMoxm6ubw3chodojIsl
ej3Y5k/rBWB4C/axP5VQBFlEURvLQtxTiBb0ln6a/Dxdm8k7uG+rhhp9VOusIJUu
C5KuIAEXVdF65i2DZijLgaz84wOBTBgtOSIfbWE/zRYhx7qPAxw3+fJdx9yu4cZK
UlTd8KP6WocVOo/9VU6gcoYnynmjyLzXRaJHMCXhHaeKBrZsG4+PB2e+ze1c/6VF
B2WvtMI6lUWzDvQtv09rukBEZxIkvNRFywMElojokIw39DiGyf6LImJZX5x8ikRF
Qbm6bEi5BkvzjhLNz+fET8JOhbbJJ/LRzVIbAOZlDhdEG4tFm2bXhc2hUSt9c3Sv
NbU3q38Doa8LZ0h6Jx090X6m6GDb62Z8BFMMELgHXR0dfJkh5KXeomg83/2DH9cg
4W1+FQBITRlk5J3+/Mfo8cBun/tBoCNf6LyegN2w12bj7eEQgKlVR/lQWuVyVDB3
cEB3sMUsQ1h+vhOl+Yaedyq7fUQemEVena7bj+w5FOWY5Em82XItBb0FbCLwNNP1
1QF5eH+g6X5pNbC7gRtp6OMKKQWQpaWn54hQeuQ6IAzs2UvErDFINezd9OUbtas1
X8mgR9dQR3udpRlAXZmt8EnV4qZscnbIO9BXHYNkrf4xOytaeTtFO0lyzt2nOXin
nmouFiqNUPbHOAXpoTRYPyg/b6VUQAAcKsni4hC/7YddX7jxRK5kfKcGrcSgfhn8
BqPO04mcWMAHv5SkS1TbNjc6vSKUSqR5Z7mul/8lu+ilvIMs0SmUfdPziGBJ370q
b1ewPGQFWQQEdhrM2JY/h5o9uogHXpNgjPHQL2DT38n8FYsNw+AovTOMFx8fUc+h
F7h4DhgDpJZGX3ETE099hmzpPY3l7S/1ZHaU19CvqPBEWiY4rdfnqaA9yqsjqQB3
9eSnHLZe0FsIKcG+sNqn+lQAwYL+toHrfH57Z4ihu+qS34k0JBcKJofIWCIvC/Pl
c2va13aYJAWiDXTmYOuPkBB5adm1AxNDYd1RnOXt0I0e/atxa6umSLxCpujGgaC/
o4y5bX1nMbcdx/Xf1v6nNyqwPWmJSbhM1RuxW6kMWKxOLB9pqdeJHl7WB9xGpyhN
4IDJ/mwKuSuQ3L/YIPzU45vjgf7V+S3E9KFpwe5LxjbbRV0LzKrU6dvXt8lKf556
aJMlMyHkJlD9q2tcX5J1IoI3BNFVz0k84J+n/VrsjpnEo2SOSLw/RZhyHIS3oCvT
qc5TKA0TDswF0g52ld0QvqYQxFQyRzXcum45tomjebU4Jn0xgStX9Y/0iF0bWURm
Kb5Q988OVNxdi7CZFFgd9R466x2w9cVsIiiL/fsW6DigP6xVm06ukRD66F6sbaMR
H43Ff7EE1RImbv75I3IxDmUXU4y5dWaigAuTR3/H9w08/S3uPtApfh15tXPoEn/U
gkgx5pVnFrnr3pYdxL5+RpIF+WmMRLTc+uYqPBhBRNB89PrpoqFzeimoQjndVozT
nXVnQDhjPKWpSjEP7RaXlYmBHqsA0GXO9nYUSxxx3Y+fT2mIbu+ohlB9yJow7KLZ
C0ZxnVzwDZ6bXaWmskzRZBH90PfGo5ObbPrTZybUzWV0ZvXe3pO6hZSmQ52SNLCP
e7dJzO6XbJoYMH2RN/B7KzgfvEOGts5+9VlLCQM/NowA1DGv2/8pbU2UD8I6grr/
epeEgsaxFc9UMjSRpNsBI1d0D1fVHDw/B624UfsjBuwavMKLFXzg5Idth68dGxQW
mmDJZIpd6Rgpor1xrzB/EcCp+Ozs5lyMOTyfgNPteqoM5MAfdxe70ZcSIFD3eidF
fGkyuLSadTNTWvVF99pPt1jWHdu3MO/8G2FJPpd1bl+QTiFncjjyyDQ0Ck8X9qCQ
CCEhDs8A9PhfXoqBjrvug/UsxlolZEvj9dOBjVbbBopMMze35ffPoKUBGllbuWKv
SLhmrAuCrokIlu5OKEulqyhvIMVw4VRbeeGdIWCJmklOLygQWNDJ/Pt38NAvZdzh
DWcVJMbigd/b4qL8LGE3dIPoTEoFhgD6hN/b1WsLgx+yHrQJTbY0O2OjsymZDAmO
nsWdqmgRFdqqmaRhiRZ7zayPdCnFeRpFybQxr/9hxbiK/uicul8dtBomVu+lmY/C
JB9s6MGVGBtQsQQxPN0wrUJt5AIXsdaIO8rIMxOc98PYnTExUXX+Kh1iswK8AVXP
oAnT/4JTEIhmi8Ram29nmj0i6t5KErUrgGdHX8ogS7TGAA+Ak5RK0m17d0p3DdY8
5GuSQGwmcGuZymS50ELdDF2sRGqpASUSGwG9E5gyjxAQrYi9QxqAfQXt6J9iYERm
yqJxVZX12DnZ4sY+Ay6YSbxtUhyG6/lnYQo7wjZyQJ8r5rPj0SCyEg/R+BG8ppnL
oUj67P+GtvTOLw7oDHR6l1j9xRnYA+/HPDIfPqkRYF5UNgpOTRLtXeH1VPoCYJgx
ThQJU2HdTgfHt9G8BTwisRh2bsW4NbPvk8xWgLbpd7W1GyppaX//uhRnSVMaiV8M
/Zw9I96Z2UVO30UZqKJeFvSl7wehbjZmYY4lKdJhbaTStLmpQCsomzQFe2o0SbA9
7gtJ0Y6b8BRxrwkNO+X/PCPVQwnfUGFXSR0lqgQAceZUBTx7QlMSa3uPYVy8HPTr
SinPOgAeDX1mKBDXbbjR9YVsG56BwvCC8Gl3sppFkRV/TuoE7qJGBc4qCSgXy0b6
xyRSwdZ8FXcV8BMIA8H9C4MpQj4ykBKuTdpruRQngP4n3Fabr2W5Nd5m+HpuJvaD
8X6/CCDnnMS066W3Gfm8Mv8ZeGEpgtefYB2BgKX3CH+1uQDVqeCXX6xnkct14GGH
ziYKczE9o5ZGERbz/wCi20dDj9se0CXAVMXIvgaXDSCmqiATn5tpfLvek/Ij8dHw
rbl/c85ohbXo+jltOcu9MIO77yveXJnBjBf22kwvuoUV7VP377MU5+Jf+2Eqn2uf
ZEAN3jvDykUeXe6wQqmsvAeW4u43l8sOX3v2E8lxMIR9BAiu4CWT4oq0AbZ0VHCv
yYkObMgZLmI5I56WxeD3lPn/97tnkVgBKpYuHgZFpJSOqLd+wG8px9pFq/TuCBEy
k6Z2i7RYsM4Kp3HxX++dPsQ7yGUza17DQJ5mAVSNMc82pkdiYDA/biNZEJoASEiI
X3zXQYJSBzLmarfDgiVhjehAF0flgQlJPyTXzed7UeJ3GQuh0/CrdK3ew/f8OcUS
JqrOFR1qyJUv3Dbd1/HYwQ1L3L55PdiYhim0wNyZJsJEEE7MJaUF4cAAtj4kqRX9
hOKWFTSDGmu0hKe1KtIJ7Ch9w6NhBPCOJHVNq4OPVF/w/K46hv+h2FQ0UZowNOze
O9BMqMcS0gBECZQ2b92YwA9Qm+ItCRua/g34xUGLMMn/VWetl14z3YRWeVAQTFQy
LcD7sfwF4ZJwQJPe2Tym0TLM0OzQEcrqAwrIp2t7EuQ27vJ8u5qyR3891TBykO7w
H3fDYt8Owr5Wz9Gw9mVMnnNt+xRxqiKJOXEPdoHTQpQpndJBk7MNAFvNYFz+/8e8
y7bIVhCBi5km+m/moTtwiW3ef8GyW0qk6FSmb/zuLr+eGLUEz5bKXrf+Xzda7NjX
EKGXx9VVNfaHfrqKNoJRYP0qXU3lPi5w9EjIBFkUcbgDEfRPaC3AXeusdXu6rp1Q
z2adXg9SoR1t5Dh1hm5WDEyKLsfQb1YVa4ZMVekAuWI1lDjrOlXPmeQpDoadNEK7
SnvEUYrEJGRDEVweygUdaJ7K0HZiyrwFLjOCDyKAxfmqelS2uZNvNg+fmmoo6LNm
rAT63nq2hmVP/x/bno4k856C6v8tcvz08/qeQJ7bLPUytVBp34LGvSZdiDi8gRo0
smZOyuacFcTp0kh1kwtbLhXIAVHA/WrBRGIbIsoo+K0eQnwXNiMDRQwAE1HbWYYE
zYcqewpuEeRKJYQw1TFtu8chEJSU/D3yqhezz9KHHCEgid9ZIuXuoFwvq2eB03dV
sAVEtesNutm2R6JF6YwVV9VhrJepI2Amj9FWhxJMuOyud9AJgxWAZ3el+9tynZHu
v17Qlp7J6zgeVCzNaas4xtrIq/2Abt6GgvBEC29jw/5QQnWGpx8MV/JJbhyrqopI
SLMGG95u/aXGBQ423GkrwjUObd/lLaaI4yL2lGeGN07Az0J9eKvweo4ESsZZqQ+4
aROaiikaurwVkDu2hjCyu1ahVuLXp15/l5GGd2y5i6Gqegyvg/FJ0oe8vRDnxIFC
O4xaKM90nBcxwsxrDafpVwYj+S9MCATlVMqs8Q695THwSLt80LspkTxEtlQjc/kW
zppBqkIgyOiPn1qpUgx8DB1wDeK1UAnzIACeid0ofoNPhoV+mlwYFVjvmvh7evaT
ohySPHxhGTWXpz6kuObP+L0PQPeiJU2EeMpXVAIcNR9MMgaUfr5bhHeQxzJPAkUx
u+OC1tpspaohJE/FhnNw+rttP7YVN5ctZigfCvWX/efbqV0pZKkMXXQDVyFMowFq
Qz4Kt8gkaCbkqnSuNwDqA2Y6ZIhxAEEKbv1oe7EXKmfTKe4v3pihKqC5t8+d8rat
6KhJzYWHHdC36HalwawmO7w7ckN+WvLG/pilEagbIHeBB0nwSTtiRDNezQempRW+
15DWqnqjlt7bjBlH38kJc9eTtXvIX1HsYCovzHZH5S8mVXitRQZoRiUu99Ojj5fl
yhofeUQxX+sxApAS1YUxVpJsmGtw6CUXpiXax89XDvHGcDHH/Ft3biO/mf/fpNEy
QtGKYtj0/wzIwzsLdeLIOlOIW91fCPIMoZIf2bU2dVdwaEKDPc/NsFW9k7ZgbY+l
40FOAciwtn7F8bM8F++YOUOp5ekF/x/v8+tlPeA9wCZZLQ9epsCeDP7rf0y4nQD/
UmPG0cuy2WZFwH/zXSHkuKemc124kuRMW/hrC/xd0MOT/r4AVyYqGyUDnh5aNdSq
oF5kvpiST0wgptDF7BzrcwAj4YhAKm7lxLLR6y+zyEUejOhWjqUl3TyykQ7VGTi8
A2e+b5WPdqpv9sgncBFhIEQANZ14/oKjuTm/vX4/IftexaFC5OzkAb0poUQ3OVFY
/LKZBL7f88dEIvf2S61+nqXGuVGM5s53XvY+ReuJLQIkE72/+IXJ0f7cWe7AmWV9
1Khg8E9u1Y1zdgKoYiYhto7niHrVc+qxQHwR/ujrcdGSjX4Bp5787AYwdbETsfDH
yKYyah54fAftUAeD0KmH7YahLTGnnbn64djTsxFV0/uq5BGOCrTKXWjTCmLzoz93
x7/emX8c+mpBqDMi63oTOBGSg7+YTUPNsErQ87KYTfdPTX9SE7qWUicFiDz5xr6c
Ef03EKL4xMjHdNjRMEXVXgVx3lvoZEKFqum/ktqbFatXSqU6iZ24deywxvVIM5xp
0pdRQ92H+/9ifYVXvbKFP8chXVh6l9/iJM/bPfuU507RYCQGcT8eSfzX+h+O7nOo
YespGU2EzCI4lN19RaJ95N4NOlXwBzLdBplSKZwnp+CnCcSA4Zsk8G4QPMDKwkMn
/b6TJsyEHmq+5UpdDRTHqD6jY+covwQZaoMzsYx9wp1Nm17GaVgHScOJkaMV64ju
CLrXZDzBXPhe8iAKZzrt/fLF7eHL+PV9W0XLKG7iuZqfZ3T9eAR5R9Gks1GvdJyo
NE96dqHlEmWcRe9oa/zN1vlOt9NZLmOFuV5JvdkyE3LepCF7qsIcuXLiBgP/HpCd
UIfOoiOxMhfQXyGCJQ++MmcrVkGzixU245ZPp8H35DEPJqy1Uv7s6LRnui8pqzam
0eFpGZtFQ/AlhA1mKN0OHl8aqe1jSftl71tESHrhqHG2UdscRkS3dgoqZf/otAsY
GZV5wpLEoDJnHTIB1VdFeBwwW/V8GJ3ndXIBtMjeudsk7zQNUn0WpVkfjNNDYQ0G
r7rIYM4Bky9ArgEbnJNab3n2iLcUmnFYUs6peeMyPrjdz+FR/4EYIcEj8rhtI9ek
63H+v0SNB/D8mb8B9G0WmKzI20a/J3jgopzIPxjaLCSvsUXs+U0p3TeecMMbS30j
s7gWFD0jH9cEg6/zqYp1prBuPqYE+wcWo7XyF94Bg1BOLdIIHciJLe1Jgvz2bZHZ
Xm0d/gOl5SflnCYnworJDWQNFd4rikDddqvdzxb+aH7tLJSlGoKEsZ7tcXkXllCv
X1KWSasGaXzSJl2/D0FvsJ8fd386jLRIuf1tJF1l4nvvzx9II92kvl9ogKNccjeA
e/RP5QDaUcKibrN16lQwC/TFKtcTrTfScnYDUNS8w6kM6Z430rDFV09nIxifKfFX
bmgECEKueLw825ovpphDW1egym/kzodpUNJvt0O8x3NfV5ejGXe9fSm4y77e8N8i
hMOO5cXMAfSYR9bGiUHZd1FLLboQCkzan5JD30FFPAa2i7uvwQxB9lg8Qw78L4mn
sj8HCvzOiTu1+SfiDhxYy//UisH274wRC4W8mHXyOEvRDwbnJz0x0ZiKloQ693kj
U9tTSr5eW0OcKYtg5CXqgM7Vl++4CSOVR7bOz2mNXyDqxfwmwh3JAfTZfAjort0M
Jm+RfPuPMbTi/RJIfXgxAOVc+mGrLEh467GgUl/thE0NiTRuihRHDWlhCYspISrZ
dXlnd4ewHEoTyxxB2l6NHJdk1BVqVGpytQ8DmUhEHMB4bojsDKvxOimYSZbOJSbB
lTs2HfWMrw9RAlUnSMBsqQycY70HRvYPCjtXoKfsi1bIycgE2nbCAXcSdYY+rcxZ
QqB1G058ZXyybuLK2XpPQsZBqiFMWv55Frd5SvvujDWqMQP2JMoZh/fC1jWfAslM
pFvClXuR2uyftYwK7NczR/1xdtmASbCkjXq7JzZptCEKk9oSeafJcNT6NTTi1ef7
FU4kwhZd0AayAbUolk2mFXl65/A3tF/oLgzxlxZCHAr8AQe9S0pwJ2Beo/KjwUzN
1+5rNBKRrAQFRz1fY7xvCfq8z2B9M/phvh4IRhMtqz2HZXdk8ubNy26Z8iCj09gC
bq9QJaGDvv4M1u5+2TLGiWHZc/+QmB8Fy8kRr5wJTp8KvtwUfAcxagcoJWaPNHuM
BHVlYuG4uPitQSoNRnl7Jl7mvJmwsXfnSnMyMQb2QOUD9fydwofrRyQpUJmF25CI
lvEQGWnyZdkLUJDJW0Dnzg3DnZwFr6GMwsO0RKHlAt2alDsuvbwXDPy3G58pVMtz
N1cOm5LjnnW4rJkXymCEpHm83Bhm46GYzrPen+JlODXIWbPrT5g5+xT2rea1mBXk
8TRGW6ePLPVn9joeZjJM0bjPL5Gif+dKFBY3JlzCnbWO96UvhJEy3KLNN14im24t
AEH+YjhLPU5PTR75rBHUCJ7eaNDwZZ1wtLL9o3g7rvnPp/vFk59hpd+0YRZX5XUG
CGAZDjic1LtCKyNuS5YrjaC9VwJ0tmpXeWOBZgP+TzV3YCH+9y6SdocNHXeZHSU8
UedVApFyetaMoqpZzdrA7SIByR2/pesoAyhMmbbrBfuiEZUAHo5R9V+FF2fOvkZe
1YaTty4R7d8h72Ukac0YVnFnRUp1y4mG3KEzN+mHE2SYEQBwA/Er8kuwNOM+12xm
aoItjSVCqHVGBGurrrU1+zJR3DxidG5eAtPCpXRahISwNldOhOIvpiGhZCSDH2yo
pCW2s2N6AN8xY8KJnbidLzmbk5GqYuy/vDQitghxedsDVwJ4pOS190Ti82We2EvZ
7CXFetAV56iN9kVF5bEHSHYG4m4hDgNd6RFa0NeoXVeJOCL8D3Y3GEtscbC5cGbd
wL7Ts3LKhvDmZ0A1Mgy6htZ2K4kv7OyDZPdtnNFm78mW8oPOhOGcqIJhQzuZYdjO
grJvTILGhJk2Ugwmb65esxwWlEseHARwlCDBvD/hL7pTpEeeYR75hK53eIM6iHzH
X39rsOIDNkwL3QjA4zbkfdCerdMFVgLBCOc+x3sC6xFLncX5qG8GEEXCKLhQpcpB
G/hWVvNo5goOB6JGNmLE02XGTQjB3WorUycgG5BbxwJsfrg6p7vwCFojdqkfNYfx
5sd90N/PMOzDG3+XmIGI9CQCNIfEDXOg4gsK+CIQ7gOzGncTCrRRy0J71gMfCCSV
2wMMW1L+nx+Gwn6M0fJ/i0waVCENdgeoWe7lZ7d/64SM/ybBlh0sltbIeMSrKD0h
rzmTAxhJLhUdVZzj4CR0Uq/nljK5814jCCwXwqzf1MHVCWUV4v4IQdV0I1kT43D8
xb1dTC8mGqAiUkCSVvjt5s64Be3pS/D0tpxXxd/yMFSHPkEYvgJyrnkI1GA16jov
KeP3dOEUsCmwIXpzxVpd8EPNKPAnFHcxQ4i5otNPv2EnYTjCY9hXnvr1qVqzRrX0
nDQtfTNcsxqVMIncxMB39hW35TC6AOLk4b78wcB0OM4ThUHPflRhKwpFKwnyQp+J
XHhbrM1f1D85wa2lWAEjCM++1Cp+zqoRBliTSDjfgnyXHcJp1pYBZsHbNtIOdk7c
YZcpZBLqMTZdyJuW7Lfiu9PFbAchVj5IfIowseo8TqBJkHB+J5kp3fIUp/EFKGll
iP2yNP6g0Zq/djdLT/6ms0l01H9n4ONe5q5ZDzaGEfNQX0LniX8ZoGqsIuzzs+mf
CdXTJpUrpPDR2NLiI3Oqe7VvQdG5dX7xsd8fgrhEBOrhQR35s1fONd5Ise/cSuam
Sl6NJzu2qs6HvBnKAeTmi490hmPStHOq2RJIxR6CplZvK4hCLqpl0MLKcPTIl4Im
11niy0ZiWAm5WlrlVfm2XgN2me7ahfi9J+2VxheeP48uP00BsD3cERGzm/lwZgjX
gx9GsJ0gOEmY55GTkQ3I25MloFNZ3bhKr3LAvNMNGczPBPkl9Km/SqUfAWNB5I3e
HCdJugFLrL8j6IwWHV75TV5F/7PcrhaNfrchQmW40fyJi40OlORs33cGKV25ECYm
db/666eQNWL/6TBCc8f5kR07ealICnZoCflfYb2SzuRoJ5mVQu6gjjJwMOBO3LO2
KxWPxmHfZSIp0mncofJNFeAI3gN3Kf9VdXe2JKMMD9rIaCIUOcNPGx9paKJ5pndU
dxduON+xnqEygTge5atOe3unVY4YV0DQSJ1HGtXyz5UFs+sa9gDlLrIsZdzpKhjr
smY1ztYNtHtH+ohBoMqoE4HaBumSYzHeCpoU+0x7YGHl1ZhWltAO8piXKLRVoWGi
/p9MKXvFSbQuic8cnD5N+PsvDXjtbumh8ffE1euzd1niMQAMq9fJ0ryu8etpBeXd
iMEa751Rde4CI0hrDKpHWSog7TuEO7Spjk16MhmzV7K2QsnAEEwASheP73gAvZhb
i+XSzXs1v66UJATBjUn3Dw/yv2uIIT2ULMzuvxEiS6s6qizBjQpIjmqvWxNN3rf0
IhwHuUhSiiNuMLqB4WayLqYQ+etpliWTpojyW88dMZq+G2RJn1RwMYWksh7JrAfI
7ypS55na0NNH2LyaM5XVsXZxrAS8Wq5RStqVzZX/09BQ/Vh+dRRd6Fp9YCzexdIQ
NS4+Mw+Ofv1Z1bzwGCyCQZlSfcfqUaER3eq+xae92Y4pCkvyZERft6OWXqbO9JJV
8dE5ssUMD35HZhX9cehYL/I5jqAPXjPw/dSUDYRLu/8DXjMhZxIZ7QUmK8Lpf4Jd
kW129QYZc9GhHfumwQ5u8OAJopJKP3/fsupi+LQF9EAq9mrfoSlEyH4Kp9uH7cYM
dswbnX3llIkaxjXumhTke9oXIEjNKNX02OsLae8VoL7JXGit5eLiLGd1M5gxQhHt
9GDJNZpgVYbgqFZqDXwKy6BKfNrjr+nx4+8CTD/SQ4g3+oekMbvGDukSib+AhTUx
yl88D+wV5qL80yI+Oyk8JdGflrp9PAdpibs6+6+pHqqACAIumHqxuBvwosilmTej
xmfGni4vaV3sdd3sxcmwFuWJGydUbCPTg63LwRZcUm2wEkxo75ST7YR9feU0zxYZ
zV5TNlO71+Ogc4ZrQzXpOorD97KFiKu5xSwaja/BceV9id5MF0HbaDRZ0GvqKyCN
aNrXXZlGoBBPXZqQd5SxIIHoDg4v9L4om/GP/6c+PzqAiecn4ra775pRmpJ0i0Hl
vqh1ziPasc/ASE6pKeLEYPpOwe5MlAcSW1R3xVoNQz4dUBDrTlCFAmpXM1AQuvKf
ReBYAuDHArmzBWZ7jvdcwGSe/bcOTIiffbG3oflNMa5/6e/ZVZWph2GvX/umaW2/
4C/n3pyC3R8eVTDyEZTiS6GciUzDvROqgg93vKgpMJDTVCySbe5nMGSzqG7Yrqz/
MJXfoiBNJJEeK3pgL0AKZ0h1z8N7G7xt3abnhVKgh6OfZIlIaTYGvpwK8r/H7IwL
luJywEXjlGEJMQjazy11pddHHYikBA67r2USS9rZ0oKo6SfYv6AYbpf/twLJaGY8
S1dXTiPuzVZxvG6OiH8csvP0ntvi+s3Fpn+Ge2o0UyjHoB9iWNzGIpiM3WqPxC6T
3QQidNrGxcI33LEWZlEq2xWk++jFCNAqJdQKbBtow3r919GX8/G59KsAK8fS/wY+
yn4ouy01OmGf/JPcLiwKvzrxymoiSgI8SKmg+pysWHo6BCNorlBWe0UVCVxncspC
UZgiIvL99YYomsnVFDn76WL4HtqeKz3EKluTXq9cjMJfQm/m2RlA1Ew/M1z/6zE3
LDZQ0hlLk4Jw0iBo/CB0rYX9oBvpJKNq8zsfR/Xih24J3e7OZcKiWJSBzh0k1MsC
fFYGsCVvNx4MfDUQIPVKt30P+G8U0O/NyTr+wQzOfoeqstJJjgXiLQ4ULXrhe+2G
z3fczvZsjBtmAKdm6PLv8c3VRbj3wJ05uHFmiXA+2hkrCPal025aHJE0fh/NfZLp
RKKZA7dBI0URZuV/fCU2OYySQcbCguups361fHDmxs3T2NIM+LxQmV2iB8tANO92
23RxFlA2sDn8deXBx3x54C2/b95Zh9ENBqcOPFe8xbCiIqIWyAq3e4kfCCoI5zEP
MwmW6LRGg+7VvO+P91Zm3tKMZANfRCZ6UZfSyYHzGlqjxCjjVCp0EUvBVgseok0P
BZfyY+cI8Iy+iZfrq8DXUckqHBmOAVx9l8d98NDCjGNkyLY2XEZ56jcO5IdzxY/K
AxFdd0yFh+H+LfucXmTAEa5qn6tW66Aob/56g48USjYirt+9Lmah4dMeBEufficR
H0iVScBqMiX7fEilgLW7JZHb1SM71TK/oWqT9dTRExkSAeZpcs84HrR96GhcoN7K
z7NlU8kpjaVKl1eI3xgpkiB4sy10DVw0+9iOnvCk0s7Sbtg9Lj32IMxKEZd8tKX/
cy01xFFaDDcCo70syRYwEYc4i15sbIvUhSVr7cfGKEba3M17vfoJ7Kf2rSNW66vG
z/Bp1BJLfG2o4SKmFX7pd8rOlPPVjM4F3war0VTcwp8rNykpjDvZRuismdsyRgPZ
ESah+1ngNmhhOafEv0PLPE3cJ8fIshNUGnvwTdD8qSPpCxMIt44vRX2ev05o0y6b
MKw6eJpWw96QEaaVIrG4WN3InO6Vc43V7OfL9A4nNYuHlTsurRqS3sCefKfCEwKM
wTBPdfZ3eVLo+wbpYrxqHu2uQfQL3pIJqodk1sJ75IsrAclwK11JeJ9xtwlBj+Cy
fJb5hYq5ZKrcH024SpcGAmsFYSu7Uw/WXOK0EtpdTlFKeCB+YkH07E5MRM8DTnbR
oXJxG3aD01Y1wrE5chGlOvubTWZ2adiiQz+dkvSoqe4GOoDenaV+rfmogBgvvvUg
yJCleFXXNrEqS+p0ZSP5od4upUJn2mKM7yaSXrPqLF/yTEF+ZRYkVHMhbsMdErW/
bhaPhmea4h5tWJJziyZzESVU6FbGp03Y8Y0gNeBD6DUnvVv+ZeCqwCIIpgtIUKCx
3JfuZ5sdO0mLA6KiOhWnXLc+0/9q1o17PDCxAFgH+aG+vYHpNfKQ+75mjBHbL7nK
qPz6hpR3+hmeop1fE1nzSrdfDUN1ITTqHyp4T+uaiHtAA3alaKpzy+2miTq26ts/
TM4dqB0kcrGXRBJfeJ30Fnz14mhEgJGFq0Nx4em3kNqiKNJtvtrqZ0/pcrCEAwOp
eoUAtVF/sMJBpT/57wg8GQOxuBgsdMSZ3/Kndoan74NWD8eOiHYsx/W7H5YkrN87
TDMqG2ylmy/fChPpQzzjKYh0AWP1lCqGIhoaVDYtakwOTsjM/J+WYUqylCA6CbS1
RKJdeTkVtiSMAEHvLDJ0o0MlMdVoQVUnX4xP8ThfbPWRMX448Wa4hMv502gtGv+F
JAjpWsSOIwNqtvaNoNo3c69jksOqUcNo884FSltWn6puQ5aUCZmT6lwq45cG6Fzr
B1fOBe3vqKDvJS25qHwfGkx5y8QrbKmhzkqALT2Q56bQwqr1ptxee8yhaeGe51lQ
3tvvrzPInZVZpnP6dSQMvhv3fQARpnfsH8QBpyHul0NspPePGIwhBzOPyvtA9n09
Zw9QIE2F3B+WjcTh6fVe0Af/vIyqqkLI0h8kMSa33r2TJGEAPSlwfy3aPQgKgvvB
o7ghiGM2EXe9SXat5Z9k9Q3x4mMMfthtq+sAmpk03xMM5kmpDy/IPjdyeNs/xyE1
VNyVGQvBCffba370UUWxBSFAoGxVhUJmktR26y6btP6TKHCRIDyDY6fvgh0la268
39bYy/ijZLSRRb7gflH6hr4eF0luZztA6Is1LbRXTnw4FHEz0p9PZDiqvQ0fz/mF
kT9qBtERDjrh4OLQMMnN+BMWblq8sCTIYk9ZgRovyJGrn0MHFLc8vnxUJZWrl70K
ZCuButeapmabegOg1YPROgU5UbglqTRwvhc3zKiqu6AeoEjA/QxA2VbIcei+3XIC
ZHN45X9ILv+QJ721jPleQwp8EBkYwrHylkuFYPpoayih0IRwFJcDcn8MfUrFQCZB
jh5izgtLyb5F4pdH2Tu8kftfkWe2hqtZHmSGJ8yhDHnoSRgBGU/vld1mxkQFQiIa
Q94Ba1xN1CxJhoo133Wx1Jw/02Yp37EFzgudbeJS99NHCfU1mSy78uBh5RdOBvQ9
MViSWCQB5mdy8pDNR+dgXHok1bFf+d77hQQAS34hyENK/4VocfPSlhe1l4HMI2px
AXHX1a22/2CwO4NDLyF7jFRLceg6UkWynpyRwb8zlqj33+vN3pgYqQvI4yFUWxh/
ERaY8kJlSm1bOii1x2vsNruQQTfCv8kFob+eDgFa9GceJrv05/aY8hI3dmO/mFJc
2OE3n0GZn6rIg01NwmcXSSP/M6e6WymszMKCGOUKVG5urefLdbl5VgDuTE+TEIPw
1zdcAiQSiP9+UzjO+PkrwKZJq210/5KQGdgw7FI0DtVdMY1Lt18DSbB5or+VzuhV
Iw/wnEZ3/flxMUaEsdM3Fma1vJBZ76AlKIPQZRYpRQliqOGuYc+jHvGuo/0/NJqJ
NZ99sEcy8DQrP+ZuqLGR34QSIMdUNlQzi6VJX8N0a7576dUhybCGbLosUSaLlX4d
Lbf0v23KcmyQU9i3+oLnfTlfGWsuLaEI8qdbf5tqmUB8KPSKOfC+dTqL6AotT/Kd
bdkMkglqZ4/n8NBVIFw9Yl8SLYjphNuDU1WcUpF9YwrD0z02+3pkJ43Xitd7gK3p
AnnaaEJDyx1oVMB9poPvwXMvcEZ3LSr5uxsBarKZ5yQ8wcpN65ckTApsI5nbMQkK
qKNspsWAoRTERq0CdsB/m58wLhMHtbWh9t916Ej7YszPxGNGPQp4zi6O46A77D2K
tPIsT4lke0DSKaEdIHiRheTvdKHYMOULjVnRYg9kwYKrDG+jtme0F+I7M07p2dHO
V6cSU09pOTVvZYN9n3MTIoZ/DqMWTz+m9d5BQ6CQBC3oikXUy/0BDreWhRgjnzuj
te39ON3ox9Go1HXAgcEMAD0X+Zj8C6CoJR1LySCx+h1NtDwAZGB0SKuVgL8Vpho/
Pv1vRIb3/1CiAz4nUtWGtfYJu0rFC6t/YqqiPexLbnvg4igal7aqWnU1UDtboYwB
GpSDywLki19eT5OC2FLMr6HALUdmjMTt3ePNFmb8bDiN7pd6gTu/y/GNoDTk4ojn
ZrSbQJ+4rmk9hEAhGP6D+CPbwEDwwn7PN4jD6L3bZTJnCq7er4mxnR+HkMCfOtQC
WRzQ/eJEXswZyMt6A2tGBmOvMacYhndlWrVFeIIFysq2xxmz1jtifREn8RrwLqSs
6u3BybcY5Ci77U7t7j01IYSyERzCdMSki3s0tGkPGFvVEmsSOTQDwY0DTy3fv/1Y
sA25N6mIVzBVs/QhAKWjDJz2TwDXpkAMl2fFd9DHpF93FybUrW8eJsAbycP47/wB
xHeMjRq19xSVuIuYVD2E5G1us/rwvdlIG0dk5HDOwe8q9vYOnyYKeSNlDFypaF97
P83Ad5roCvcHaucE3dsZgo5g0GJJMRwYYT8suLWatZ5t6yN/3NqCO4w9uzMBHKOF
OhasSvg5D2fnCdpBhmxvtTd6HiB0BKV7sBYYWyzerxhhaOsQyJKMOIMUG/6XOCll
FBGy3z6pFAzjsbvgr5HFZGGI+jSxpZFCeLHUZevrZM7HqtyZqDLXb+iV9ESbhFLG
LM1m8nwM3N5CEm3pFOulcRt2gj0dQVRIHYzogUFyTuHvKF8805PEQHYvRTUK5GpE
tRjpNrvbrSszI1fMvmN5LPUpTiWm0swioiV7UVgk3IHvUuZ3HmBUnP/hHvmq9OOC
fxJCZJNA6JKTToJ1UmICZkqq3fTp2SlnpDrGI75WtCrxZkWVj08I+MwqlYnIoWlG
RW26UyBHAA9T8dRAL5HS8iRR/OUCZYgWAKv0rqMNsrwQ5vr/x0KI77L2YR8CAQKU
v5/Xh6QucIHo4GYB6r5JllEY+Qn3LHxx2n0it5OrBGjU7UA8jV4liDlOwy3LBoSz
Gc63mBVLuy5Guim0ivyqA7k4uqmPf38PAbUvKEnoJ/+ieuh199sh5rD6VJWJvmyZ
GALKgMgXar2hATy81qeJSB5DjVoXxq2pvCH9p6/o0IpWoSEsOUe7ydBoOuG/WQUk
5WKFgTWc7QFiLHKa4rlqIfyYtIXO3RaexzfCZXyeQ55TitRukaNK8vSDrLATX7lx
6v1O09XIRZnhBZXjfRjmSvtXaKtIXQyVpFU82w39ie12diQf15COz/IEkJi7j88U
Lo1hFDhpCypa8mvMspt6RzbxjQeg0cPDZTF8Sy/oE5VRMk9BmrJSEKeUClV6kMh6
Bq93tRGSEvsAxRiCGiVsMzQFrkkHLljQBwx5s1VHfoJAod71AsejxEJTeejv7Moc
6YBAQ8E3FNLziKs87srFO8t4Hf+qGEtZ4/ezX2TcAzHsdBf05GaOkKuLkP5Oo4b7
N8mpxirsRkUQXHH936ir+pgwQj4fxsBasDwGug2fQCOw+mSFXUQnB5puBlHNj2Tr
KHTpeMARIPznpU9XJVdk2Cl4A/0H6hOBVdwvPFWHrifpEo5BIVP2pb3KPnhmDUmV
EEZUzlYz6wCm2Ttka00lQUYVniWPdydXm14dk1KwLqWDuQXYv53hOFCSjavKihgb
yTr3X8N+UnAsbnXP5XazXxqC2RVehM4h++yaEx8xWhw3DLj40+1MCyK3lusVzs9k
0/BL95kjhYh9EsC0lhIh65ZXTKVrqaLF/qNrx+ZjPMWzZu6kJraVFW9hBVtlfL4n
JEAeEb9Rbe3q7ajk1zCciQx5X2HEQn98FgsJg0MxpW+nJYw+/xfU1uvrHt0DGDgL
5Q1ANRbfnFehtizG0OTa5Fa3DzCB8aaZCgE0taFRvdDhpuD9Z0C6yzSYlQZTHfnC
9KR7YzcwtM2UU1n7nBC1DlM7aBKsmL68x7s61jpGOSGAw1LF4J28wSiUN77Dmip4
gHtzuy+9QVBSAQn9eoD64hTaCIAmWAmugGyEO4PrwiUshxVaTQi4MsJhxr25BcnA
+7pBxAxtW/EkZPiIMGbEkpZAAaq31tX5U9YFti4npxnp8Oz8ysLkftEe/JNqdbWr
6sZAyVi+XvxGOabWZkbMSyvcQZJZifcUanhGv0d0jFNZKtdWJOeoRPvn6aznRekv
lgQxO6qoE/9ZnhUFlicRR5796/0hk4V/61+rh37kpCCm6VHqYYiTgTnw+Ldn6XGu
ck83oPNt2XTC8512ABVgxb+6K1be6Ns9MUzTfqwdwgg/MsHPgCj7NlUEdbn4Axrt
aMcvCVglXhvoIJ61Py59gnJmAfYloBoG0Ld/3xA4buhvqH+zDRKtQmnpDrNc1RDg
Fdfiojovb6d5d5sCOIIC7nOcAQ7KIG0fsY8UWJQ3tPziHW7XLXDY7ngDw3M4bJMd
SrIlyTHvAaNbtUoOiTp9DuHankUnrdHQAbPlpPjSvKOLyXltWxYck7/ydb/jNUgP
lDS+SiyhaHVF2z+SXGXp7dlNeHuq9fiCcGcHVyRKWNSrQ77nvughCGJIqv/0EHIN
7oRTHdDv6o6CxGT3TS/KrH/vm4EJ8ouO/bhZhKDaIlF5A1CUKILHI8UgwnQzskBM
ngkp0HUrI7QM7Q0cufmhcEyUEKJNHwlydtHKwFQOSkpFcs1BzL7F+YvAP55og6Oo
3ryh9yaNakQhf9w/vpSFzqFxPs+/wcCQ3RUcgBuo7W1ZUPYeOJqsFN9dOCBpS8mF
9tCQ+Idc/e/C9qUtMG6dYUqJuqYKg/Bkg47nQIKATdNRAT4MQ2oTVBGCnv2IHk0c
GwqjLGy0L1puh+3RufyBfZz6+yCaQLbnF1tzSNKgLl4J08mBEV2lPvatxcyXxyJF
FLZF1gUY0YjH2doTkGrAAHhzKDjoetJohKp6lbofLCR3EtMgt3tj1v4VAkNKGWm7
9ZM3lhLjy2JMxbcQHf/7S1qvvHPaO4zlKSI97bxNAYLhEcVHCYGxatjk4wOBNCwl
9cHSVIVqYwS+sQijW1KsnlO11YDGjVYyCrlMja5zK24kOZviCBZl7hf076yFCnsk
RMcy/wSgIHoe13rqXesULqN3vdyHSb0h1FF5kreL7vcFsvm3JtE3HArL28ZlWTVf
ujBeCAWrRJj3IagOSJ0FhEO1X4Ob8lAI8egIEJz8jb5OgOd2biq4v6X/exGkp14i
gY67YQAD9KuDWi3rWyel4SsbgroOTjFQPhE5hxSr0UdF7lHUP3wbcMqJESRqimKU
EALDb14bwG95vncHLbppxC2UynF3RczdIMkF7vadp+8/3EbT4WrADIQqurR3++ov
vwhc+OI4Qn3Lbm4YzlerUo3JB3OxA4bUImsU8VFeA0E+c/vz/aeA3JJM+Whrtail
Ya8uyJ/ZmkdDEVfemh9kVLmLycwEuHCgreAuvAlfXmkrQPuCyzsLZ8p6kGzzLvJH
V37nAB2uk76zYCbQK5wQxzjLntCR2SVWxOG75gc1ui3Th1cDUeOjTDJIVzww3ll3
GJCb1iGYSPtEGlOrYOWE2kchsMc5rI2vt5AMpkIL2jqN16qlCh6snuZOrWVs19cW
pUV9X3WVLjwh32hHVbFYOJiSC4k7qqhxNrznyJUQNvKU9paU/W+iFgawivZcZ3Tv
pPsLWmhm11eLH/Vr4B6yAXUpSib9WGUFKaW44/4Y4HwMu9lYIoLNTYIiMOM9tJ9+
BrxEUu8TMGUiEQx/reyPDpOjNc7gyp/GfUK6T9Z2SZBAV8/pNVSkKN5k8yT8EaM6
V4KzWo92Of0UdfvrLKhbkNsBCDfuoi4/DiM6Y7eXnZh2DJRcGUMnm/G8KBCawj5i
MtyhiDJdU58yW9Nh48DQSo25ZzlgHec3dk3q0jJThJi9rNzOVbtQE8QKj3ARHtS0
GyQFPgV3QBENXxG2VHuO7o3Ihc2Pw72lGjRsCUPmtUOoCb/c5wYt24ukB7w+7KyT
HxakAEHNsC6+9IS+4yqp4Y3wKMRU3Mup5c06f9xcPX44GbhlrCSU0fG6p30Lwqs5
y+759nyvYs1Rc3V1/azml81wXC5cLfvnh0bJ4j3WNJdeW2e9q5gzw3vRsMcBXW9K
LKLFuIaHjoGduZTPOWD5y70mTkDlgG5pmSxKT75rAe9lHVQ3o5MMoZUD7KwtSpjn
nqFKwAxXrinYXIyMsZMj5YnT3hbh4nESmwSlWHlhBEIrMFr6u8I5eM6xsdA2sDJb
jzwzJfgQe3B2QbxpH+4sM89LdkhVm3H3CUKRwLwL4SfZ9PJrYX19dePMoISX5Z9A
4uoNmtrEAWUBqcGZXnkRTBYbbuZkgB45AfFUZdEieiRSp53KWgrig6T52Q2wbA8E
HSB/i46HZAtApFQhHpxV5DeB7riVMc8C/Wpbyt8nfDmYpWj0e9IshIsq/Rg6mUcZ
QPrUusl07NpYdqkCxbgnWtEj2HZvV6QR/bOPIejeWY+ukwWAZSNQz9Sf7HY40Qxu
5wf/GFeeodDmZ4ngqpj7Ht4TZkYhReXT/yRtDCbNmoX0/04Xu6fty2W7KkYJ/8UW
OPofM05olN7OBFPMelksU36tBWauYCHUh8PXZ2W2iy9XL1evu9l+M5btOTV9OjT8
ZpZSWs862PuaG0r6KXU/nNRPwboAEKurbG6cxw1+bhiT8uduENdv1ryXfOlRFm7x
akp079Iy4K4Kip1nJ637aPWbvtQMRIEUBNxZPspJWjwSdvteVUkxpv/4xhtlkhRj
L0zZmkXxqsQlorf3XdGznoUopfzbZg6SyDMl86pQGLmvEOs/eIrby4OQ5qqnJshZ
MiV96s1h/51Wy9Xw7SMnXPw/KlwP1MC1Jh58qD46JVmdNW3l+4B5p1lBV/Dhiv1f
E+B7w9rKFSDnPDo5t1ctUv6IE82VKkt0MbL8f+eDTPe9kpVhoFkbYj01XPVwzP2T
cIkK1QswwmPpmbIBamaF08BkWt56fjnO/dcZdQeJ0+6DLX/YFv4UncWV+uyL0t//
MgFgTkW8L+5xQEvGZnDqps3fTOoSQ/d2mI4S32SA3cfnHGnbynHnkR7/2rf76B5V
ZaWgEojLoJMkC6Vc4PnKpMU/v5VxdVV6LiN3C7FRt6i51nhdqFKwJUCs4uPHqTBY
VYHViRfre9ynKLZGiqK1YM8rTMyFsTbrAf1nmk9/QiPdygwpzEfRlztnSEtWWw7W
gmM6P3rzCFWE+JawVtOF+rDtLY+nZOwlXKWYTjFSc0XEF2vMpfbZUVq7LVhxxqRa
M2FM44ZmmtHoKG27gjV/IyMU3987Nl3+7IS/DEwuSt9ZVi+NiaW+snwzLxePdN7/
8g1PpOjs5FljFMcifMwu5gh+Um9vx7G3YIsMG4xnodSHjwELsoOMhG8W8u6I9yce
xfNnWDra1oLP/SjAhurzSFgLEDlDH/SkMsexlYY4Dg0lCRDx6+58udOmMXN3vVHg
pnHJzxH+2IBbMkIQBQQCufWGmKiSimJwW/wTxaf9mqitswCo6bkupJXitbAF0XEP
O108DYIC6vE/iK1/VfJbXKhjfp9l5loy7vrpY+d9zpWtJPsQL7/zEA4M2hKTBWs0
Oubkfk5DoLCotCI5Dt8Fqg9esb6ZLXxabpZ+2mo2cSs1XNg04KoE2oVG1V+4o0eC
BYzlzeh/jOLPMFBoJjaGM5j0PswpeFPYuDj4bG8H5hboblnV/PvtyFoQExYvg8+q
TUnYiuytNZz79yd02U4Cu1oQcr2Fp/UczpKByX4pSmTNkxycD2nB1Ul2p64hjU0g
W7EqVSo3cI/c4rx5C3YKMtIDpIxTcs/NOUJfUQXmzCM=
`pragma protect end_protected
