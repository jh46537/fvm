��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2Ȫu��Z���d�]�$\�h�����oր��ʖR
hgO���m��i�Z�O�L	��M��a�ok��Q��r�Է��z��1�� ��I�-[�?T�oNmMǮ�y�B�ˋWC!�}�O�C8wְ�Df����)U#�� �o\�Ғ�Y�b�n5�{#G ��k�O�e�X,j���Aϵ�\i�h�nMOŬ>�&�j)l��"�#'�[X��^�Yh�aH+�����oJ�	�ge� ��G�9���it��}K8�+sm�;��&��=B�V?�������z[�`?�WZCc&���:�C�^��t�6%(�5��LT�ק���;���=r�c�,뀱?Svx]{�����18�Y�Č������H��8/#[I�`�nm\�Ɉ�2�1[��) !���֘Gk��%.�t|�)#F�\�B"䡯\���Α�Z���n�+r�C�'��3{�x�ɢ>؄�P<��[�]z8��+��t.d��<�ջ���P8u���R"OYX��8}e��$��<��V�2T}�߱C���G�S��V��:�8��i_jB+��;��������HΛUI#�)�@���U���qJ��Ԭ=M,�C	K�?�%��R�'�K��;mT�� u�n�/D =���x0��3q�ʴ3��rq����y;FRt��� ��
�ܻ�K�><�h'��X�p )?�K,�_��wwm1����(LE~"��')ۓq&/)g=���s��-I�������bq��;$Ap�����dʨ�㑒6�F.DQ��V0�6��&j��D��>�}bo�L�0�ʏZm�C�	���ύ��~�X�5Q����7�{�KD�������D*����d�+�R��_�]9�a�C}!=��~%+[C�4�Pua*9�����O�=�}e^�*�dLe��R�h�_�e���6|�.I��m��s�귋��D�8�ێ|^�5�B�蔪L���8�I���0 ���ȱ�b�辊��o?xC����qp��EA�RZ�#Z�R;z������A���D�_	x���w�G���0��B`M��kM�)�|'���whR��,	ȷ��B��B� �o���m�P���h�aۻ}�#��Ȍ2��/9A��Qw '����ʣys����$���Hp���NN������k�	�n�vQ�%=�yc���8��AT����DF��X��Cv#��m�NzqvVm޶jMEmj:1PBԘ�f+C5VG��H������cr��L�YZ#��0^}V	�!��ͮ����AT�\�D�fz��20����r�����	;��m�]Ҽ%��:���ʩ�}�qEA.,l���T�UW���..,��i��{E��ߡ�!�y*�tr�8��J�i��ɣ�.`){����&s)���\�S�Q~���=�s�Z:������vj|SDd�n&�'�U��^'�AJO����njRU�I�Q��iV���0�7SaĐ�x�?�tx�#U��@?E�ԋm���!�Ȕd�&��&S,ps��p^��-"K��μ2��4Dg�-��y��αۑ;*�x��е��`m��i=�,���=ʨv�A�bD��]����?��oW�Y�� �q^ϙQ��'����{����^��$ó���5�<���0�":����{��F��@P���M{̏���[��w�6KϮ�������%o/��F�7te���hً9��k�?�vf���|��;�:0�Ӄ�T����Xں�2N[�D
��|���q�EB+ԩu91�Z��:��d�Y��&��`v�9>���:}������.B�(�$��Yh+В	X��k9�#S��y��¥�"�	��s돮����|)�����< �k��9qw�&<��eeu,#Oȑ���Ks��f�j�(�� ���V��mu�F�U��Uu��:�[�7;1f[R�%-:m">�,<c���#puJt�l�m��<Gugs�i�YlMd�[�5\�MN�@�uj϶W3l�b�rc�EP��m��(]���p/Z�߆G+e,�O ���3Bn����X�WbH�B���b�[���2Fu�V�8?Y��S��!�
8Ј�΃t��o%��^�e�6�F��<Mg�v]Ôr.�F�9M�0�gv���i�Ld��S��͂[ ���5/���7�Fޔ�-�9
�GB���B�iI�"`�g�7 ��31<��d�zƛ��w^c��i�'H��9ό������0�"z�%�`�����O��H��t{x��[�����Q��.�����5`e�����j�s��`c�@�J����mM(�o�GסBB��f]��^ӽ��
���dI�����C�k��9��:�&2�^u�����ZA�.�FKoT���_�?��/��]h~_��)��y�ɪv����{�mY@;�:��	��<�#'��B�x�'eU���7��p̔�*b����������mg������wrЫBԺ�M�ZAư�uWq���.jQ��O*��y[C,:n�L!�����q{��l,���On5h�ٽˋ,�U�9]gy�����_��qr�Jy�Q˱�h@lAx�� ��G�ø�w�
ɡŪU�J�KŽ��3Ť���In�K�+��b2k �@*��fkdn�.U5��Y,)�Uh��5J�L$���s_f���Զkȅ3%����b`=��3Q�2[�}�t��ղ@��5޳?��ʱ��/���%��6��'%m�������4���>o@m����O�ah�37 �C�p��'-(���q�U�	�炕���O���/6�hV0����z�[��j�A�'�nV��x��u�H��NG�sJ�~'��Ć�Sz�4�4�6���Z�9 ����l�RS���f�ʠ6��L�ߺnfO���x�?@d腅�Ů��
y��6�|�@r���g��Q�QH��+>��rzxg�"�F4��ϯM���U�k{l@Q�D��#��r�~�b3�l=�XliWk���`���5�/0�&�	3T2�tk{�$�F��H�׷,VU��tB�]1J�1%�2��|��Pw�5�����a�X�x�>���U-��Z�c��?qt^ZP���'�E�O��h�Qaqk^�Jr�����&hl�� ����1� }��֥h��oUcJ"lGvj�΀���LH��	P�;��/��s�(�'^^
���o�����g�^��n�.w1���;�Y�K%�T����^�?pf��6Bz1NP;8��k1"[N�W��osVR;=���M���P�q���`q1]���}O2I�¨΅�3���-��1q�(�~qܢa������,�����t ,�Yk�qZ����P�3rx\����>����6���(k��#E o�V��� ��AQ4ܰS���k�}<�R'��xn6�)��g�� ��r&Jz*{������
g�S9�`,)�d@�gf)��1�z�(�ܚ��q�Ӱk��d�ԌL$8�(n[Ǻq����r�?�Ȫ��b?�_�J���7g��~�d��D��<%��cWUtS]fܝ9��]��l�kl�4H��zVR�� �^�%I��T{�9�B-�<=>�Ns�a���V�w�@崗�&J��[�K�����(����h�*��
�k\A �f.}P#iU��ƚlɱ�/d�*���7v�
�u<n�@0�A]���Nj��D���)=i.��$�0�&�/�Z��!-I��Z�Ő���-`rbL;���[���"a��xf�<�C*��+FYe��o9�n�q���"a�=�SU�M��Bxz��O /H�<:\�}�Hr�׽��0�el1�����o�n6��E꤫�0N�a����Ŀcf�x�L��Gv���ZCF���W@�;�k.�T�WnA��5�M���<�k�W�p�K؂b��o�^:���~�5��5s~�|#��j���{��`�['�o'��������t
��g���H�|>�9[xY	�,�j���q�ͼ0ČV�K�@�ٺ���="�2�5r�ZT�Fm��ƈK��;�� �����b=!Tq!Ǩ�R:A�4jVQ���w�ʻ�pZ�9֞�[w?nR ;�����ZqJ;R6
w#��ȶ󄆀ԧ��8B�Iw/�C��El�phX��	)����&>1X��U7I1ޣ�T"Ҍ�����Q(�;(U�0(�����͟�׃�,�1=�d�n�����.�"F�F��=�����~jJ���t�P�"����b����t�ѫ�B�ϷRr��E��3��߹���(�;���n���\�ծ�j�Hc��5*��L��<�t5TA��+�2Bb��xB�d���c��{!�&�弓��9t W� �M4�s�ڤ�C�}8-�����u���A��BS#�|}�0Ǚ��tnV V#qEd�[R��S�Ͷ�,Sg�	>6ݳ���'�2|<�!�~~N���~Ec�y���x)ֽ~��%ש6���'e�'4�^���4ym��ͩU�`�nPJ|\V3%�km����/�"��]i��!�r�����mu��s�=�*W���Ej�K�j�B'	b�ޠ�ʙ��l���۔*���(�A�9�xM��L�'X����~&o��S�ŋC/�¸�2��)�4y�T4ʏ���[>�n��Vz��CD��A}����v=��:� /x���g�
��о1��XTvR�"X�F��5]`>��H�c�G�T�B�N������]yx���rh~�ew�=#���,�g�*O��uS7�@+��]x�H>�	�ث���{XᏨ�8�,��3@鎻�ף*;	�����J�]R�%�1?���Xx��u���_�&A����N`��0H4Wtt��&�5HB��5��-9����F� ����k��{ʎ����C����P&]d�_ÏN��CA�5	.��^�F��.�|�,$����U��XfY+�7���o���j5%�҉��� �.�	
�g+Y�G�=Sw=4��$ϓY^�d�F��&1��m�*nסo�]"~Y-!�hç���������f�6�Nm��%������T����H[D�I �5��C&���B�ԗ	����b�{��n#<G}0rR���wh/F�ڦ^��
�0�9��(W����8�1ĵ�z��O�De- ��~��@E��Zmq�6�p�~n�E��7~zG�uO�3�夓���"�	���`XHiC�������4���͔ԄQ��,N �E}��������J��7$��h]��Λ���4� ^|�g8���͋3b�-���U�=dl>�F��$����
3!ݹ�kº�� 7.UJ��8��cB�N��>�ՑS�L�*����a���^�Ⱦ�Y,
��'}㒸?l�t���5���i�՞�@��(�]��>`E�?T_�k���{(�+�O~5��E��G�k��""��zZ��a0���q�`Ī�,(�K�(p���bʷ����f5�`��-���A�MT��+]]�&C�k$��Mݎ���=�?�M����q��`�%f-	g����g�LEZC�{D/��-��9���6Æ_n'@�	�CH*oR�zt�N������#�j����&���ى�[��F��P27ͬ�����'�3p���$��U��A/��j��x%��J��b