��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k{de���ӱ�&hc�.�z@4�(�s�_$آ�������1J��cHzE/�Y��{Q��k��>-䃿T�E��p�f_5�%ޔNQ�d#�c G���?�Ʊݙ���}]�����B��rF~��g:�̰��Ay���SAM���Cuc�J��6� ��5J~�N�,H����e���#�7�R��g��?�1�[M.�i�(�'Ӱ��<����9���Ќ��)VVG��@�v�4fݎDJi����}:��������0���C�=����jۓs ��S5��-}�\�N�	�ݹ�ɘ?1�m�'�=d�w�8]����P�-��c	;�������w!=Ϩ�ڥ������wi;(�i���xbeM��-Kn��YM�]֓O�������9jZ�Rs�U)��C_�vq�tJ �zāY-\N �'��l':�w8��k�����4T�:�Q7����kU�*�_z5W��fsp��a�ۚ�ՓU����
�`�4�7����oJ�bc�3i~�,�����/p�S�E&�G�d�G"��Wĉ�b��~�,Ret���&���kH���5	2���$�!����D�y�W'vX��H�yEXy4uS�m����q�kЇ�F�9hJ���m�������%�B����q�@ն����?��B#������XN��ϻ�	h������m^ D�P8�P�wT[�צ��/��U�^/�eF��i�F���|��RO�.G6��I
�O�8�	?>rk���������a��RLд���LQ)-��
�ڸ[E?"M��e��U�Ԟ��"V�s˷���X�DN|}T<6��{�|�]�K����?`�K��a�����עL}�ػ��"�ާ� �u����p���)d�X�B��ح#�� �]�Ǆ�5eľ����b��y���'B�B�ܰ$��]��+8ku�h��D���%�N�;
���ܭ���:�f�w�dS��+�e��&��O�8;��W�R2i�