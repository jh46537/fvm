��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�q�E��	YjpA������2o&�0���c�LڄX?�i��+�#��7J�n北�����J��kƧ�6���+{E�b��pڢ v�U��4��WL`d%�Zx�Һ�|�N2L�\����-�1s����#�+��l��"����1,h�'� ��a��I�k����^	w��G�Z��k(\H�9���# \����5AA�f��~o�ItMi������)Mn���e�4eӜ�^�����[)�F�0�?��~��w(-�f�sS��c��7����3��/��ֲm=o@=0�*QR��$�Ym*2�ծ>"�j��MZ�)є���8���'.��]����Ai��b$'�c�]7�a&���S���,�'1�O�U2�"�7�;@�医�.G��C^K�F]���_�3ϸsN���ј��`a3mWQ����UJ��|���9�~�4�3vf�b��aw��_��nm'M������-Z|��0,t�f��06D�x���kv�?�����Jޤ�l��V����8���K%�&>3�������������K[��lh�rꕩ��gl��!vrS�]�`����֝M�/�c*ז��S�Yy�
�.��Q_ۍ1��I�9��a�nX�k"�f_XW�D��5��6������m8�Z�'�%GvG	0L�boK�H��1M\��چ�H��t5���U�Zy��/e/��S�q�[u|����1s��` 遑�d�ʘ���#�O��P�E�\�1��
��>�[%T��S��:���q�	�K�˟t��������_J �%T�c[*�+P�7�s��:�4�і��/���i.-��x�a/d�;�=JJ�͗t�����#c�ۢ�74�k��o���_L%��N��0��AB&ͷ���	j�չ�d]K=]��\X'"n\�:�&��?g<��D��&�p4߻5T�� +��EvA�j�C��A#d`Ѝ�p�T46����~��޵��`D=���X�uZY+0Z���+=:愯�Q�D���&>_9Ѱv!>�ݥQ�����/e�׆�Rގx���d��&V���T����[�� �9��Ɂ��<]Ét"����b`��fW�����]I�9�0���{z�=Sд��J I����!�D;z����2� �7����rF�`�w���1OT/'Z}��e��\7�ƪ+�q����ucw��B�R��f3=��G��c��^́����z�b�������v�Nɑ5�1��T-��G|���C�_DY�������1�޵�����}����.����|"�A���)p�	O�a)G ��$*%1F���0z�1��N2�Pd �KF��fO"�%��u�����m׃�"�J�q����.m���BT3��k���_��K�Fސ�zA	�z�6�T�&���!F�V�� �J�p(��E�]�N M� i"ٖ�������#���y��y��h��8��K�f*A�6�tѮe-q�eôT�p�GW��V׬;�@ �M4�'�o�h�����_?ˇ�~�*X4��RF$3��(Yʀ��˂�|{��٫#G�d�(I��zܽ��"��氵�������F:f�/�|�)3��,�* @�8�_��S�XB��RZQ_�vUU�ʂ��b�l��"�4�˯x����-�Zf��H0���z���CA;�v�� ^
{P�JcV�I~�Yx@��� #;��m�q��^�3(��3�5�7���%��ޤ_�K�g�����7/W���/��(P��Ԛ]r]���pͽH��=4�,]�罥LiZ��[8��Y<�j�fA��T�b6O
t��QmT���{��䑢�vJ�r��qN��'�A\[vO�m�w�kC�x�����#�&+��u[�5�+x<Z�_i������=�@����v�wMۏՇ7(��$u_P�(c�o��m�,���y�yx��?'����xL��3�7�����}nt�QWހ3U�����o�6:Q�L[ Z������O��fCY_���E�L�Ϥ��Jø���5I�_���v�Ê.Tf��C��
en=uz����9�tOsqg���w�i��O�D�C���>��*̱2�Z䷉ϾԔ�c�
я��Jt܏}�����@�>�pb���4�5�~X��c ��hC��w���C}�Ts;������D=���?%��D�"%���$�Q�ȓ��ׅJ��Hχ~[Г��`�%0��@]���y/�,eR���Fu��r��^�����X�Z��J>ܬ(La[��tҦd �o�Vz�4%*~/��& �j����55'�
�œ�0wa�#v/�/��\ۚ���� �uZ	��n�ZB�y�[h��w�ZQ���W�;��CM�;DX_�UF=u�R�ۥ�Kؘ��l�i��r'��5��P�q�9��]�H����}�Vԓ3Rd���V$).�$_�Yr&���@��g��v	�%��x�~^���>�[V�s�vYLa��4PfΪ)^��ΫѾ���U��Ո�k+�5Q�dW���a�rB1�h���(��Y����ל��8'x��=u�4�*���8�h�A��(i�"�ʧ�^U�/�!�i��\Ⱦ�y�~V
�Y���|W�R�*�
�'C�=c��!Z��@�z]sz�<��s%�0:r���p�0��;�}�M�1j�A%�1.�Gī���7�-�n�ѥJ	<��:8�:5iw�:��I�q��S����A����}���l����|�f��J9���q�C�{��<���\�J��hѹ���{[Ծ���9V9B!�ҧa�L����E�~�-Z��5��t/i}5���ʈ5�N �gJ�Z�4i�|���C�ޥ��̐�C�C˪	Ys��5+�<Ln�A
NbꝦ{o����k	�����x����W\�A��S�H����;��}���X n@:��-�Q,U	�M���c�SS-�xqx��l�ܷ��X��쨗�Α��4iCf�M�A)l/ɹ�1�k��7�%w���'}S$u��L�+�<u�,��^�자�ܭ�	�h[�}m�
��oH-��]�|ɷ2�fض�IO)���x,y3B��������%��FCs�Y��B�a�Ʉ3�&4��`�� Dj�81�lv��Z����s�-F��[���3� ���3������1�b����?K�)�݊�n�