��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{���b�e��_�@�*��Ht�'��p�z`��A�s\겸��S���5W��\!{ә�Y�ea��S�~B.Z2�_CPCk4���zmD�D,�Y0 � \s�i�E �1���i(�2�0[j�!���G��A�$�l6�a�St��CJ���@70Bg6f�;��}� 0Ipj���&%n�W��iy�R*��ý$��4wj��`� �G����'ѡ�k�:�}���/���!*]�S�t��ǿ�����@+�sL�����B����Vc*���:Y�ϣ�FO����*�s	]����� '���q��0�����@n@x�:��嵌�;@M��n�yݍ����V ��a��xS�B���a�,�Y�N_&Zll����4|�M��(I�g����Z��࿯�sw�mO�*)O�� �������z��p�5Zil����B��O~	ݪ�{��g�׎���B0؝��0l�
X�Gg�����5��q�b���}Q	�oa�5Ds}��+)�	ޞ�U���~�ЫP?sT���-H�"����4rT���K��lR�n��F)�a�y�|^��+hvHz�+��|~�?��=Ñ���
p4
y�ƋZ��b"qn�:��-z�%đ�	��2�E0?�*��
(��ހ�eb<��]cQ��1IhW��1�ܺ�������{�8�m�?T��д7?�8���>ď���뜒ϐ?ư�婕��ǬiV�+	t{�;�B���
����d��GM�KDu��z^��L>H 0�OdmnN�KB�iq���
��N'���c�j��� ́>�����-���i(x;��v(c�@U]f�����Uq3�}`YH�TQ��K?��l��-��xv�!x<�o�X0k�=nyu�Lq�y����A�!?�|���N�Iq[
F�Ճ�����OW"�a!�I\"��?j���N��8Aa�K�n��r��v��I��H㼆,��0I��$��+�t�n���u��ߵ��P�l{=�NIq �@-}e�K��p&k��	����T�ؔ��������3Ư�f�󇦱��a\�=��H�#�iV˅$MJ�`��ۍ�VJN�AӱT�&����kfn��Au�jx��&�;�U��!���h���5(�(�-Y`p�C̓e�j'�)y��g�tw:g��]�,��2��ww�SS�ɴh��Kr��*�3V/0%��S�V-����i��d P����j/,A�6u�V���Wl��������Z;Q;E 泸0��g�`J��1/�p�~�B�8��Ζ�O���=�A����!�}O-��Hzk�I�Y�A"۝M�{�N^��A E�������k@[��':rT�X���e�O�V-��A��2/Ŏ�;���A�;��8�ލ�T4��'E;�3Ҩ�B�n�͚ �1���
V٨�Rm늮1�W\>-0%�I�I���ic��~��rf�(�K4�z���8r�ߤ�߷�G�����/.��:�aI�+��Cr��0W��kI�.j?>R��0�^�<��
 ���_E��+��,�#86����'-1�[��� �<a�R6���Z�)#���ݏ������ �k�(6E�E[a�@�zf��M |j:�.}��k� �<+�]TX�X�b���O]�Ja�F��=B@�f'����P�g-������=s�,r6���E[���α�]I"�f��*�6������u��Aj��,o_��^����y޳��/�b93�h���`��)����P��d��c:BG�p'b�
�[!��)���wl���r�a[���b���9�����]���o�����`S{�n���i�&��g��\�=�-6y��1C��r����@*1������ 	ӳ��2�F��hf��8�U ����:̈�|H�(��a����a�%��>��Nh�I�ҩq���¯�$�.U�f����iy��Q�l�D�~�l%�iF�:q ϗW��AOѡ�T�G���&	�v��B�+��o�E�V�1揰L�+'?/'a��y�30՝0R�R<; 3���0M׍3��M�cJ
�2��L�C?�1��c'K#��6��(I&ljd����!�����y�ԩ���ճZq�,��=Q����ӧ��]�E�[�g�b���ڑF��WǕ��E�#�b�"3Y�X�A��i2�Y!*�g��EP)�]���|���H�[<�S��팦����\�'\ �~�3��WN�\k����/�v��4~
�����~�-�Jzʛ��/٥�k�	�RZ��Y6�翛{���p7~��7��'��dE�8�#*����e|;���jj��\�����L�u%�ރ��R�������~z����j���b�G=��{r2��d���K�����{Ne�L@�W�	�l Z�h�ixDě�������(r�o޾��A�Dl�=��=����k� �B�Yy�m����Q�
�X��B��=��@�Dp��\8ӈ��P0Y�Qu��,�V�=F˄)��k`��2刺�\`�W�#Eܓ I��f��.��Ǔ@rR]Q��k�N)�_0�Tw�Hx`zD�@���<�2 ���M0��~b���5��&��K"T���&�1�����ba	A�娌�WB����.�ՆW��u+(?6��1d9)��d�����ڼ��E̳���PqF�&"Ջ8��Br[�j��zV�ϴA���0H�-�c���Y�=��,auj6+�1��=WX�i1K1�0>½w
2֩�ɋ�cc	̮��̼Դ�[��G�U��uB���-OK�Hp��٦y���x����M�