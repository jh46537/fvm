��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��b*]���I��̞m����
��6&r.Vm �qx�������
��VQ�����QF���9d�7>V9�<* ��>�����qf��:�_W���6��v��x� 	�ە��A�E��0ړ;�W���e`��a�"/�??��+��.������pK����#=��Άzp�l���Б�M���k��E�ѻ{���k�����)��+OB��w�S&�)K���'s�y�"�ѵ�j�����X��~�x�;���*m�-D�S!u�,��Y��5'.|uJ�a�v��Jyy�n���^�9o!_8�~8R4[O�[��R�J*N�\Ԇ�t6#�&��1���,N��*ng�U&�{����<��$%ݫR��ڐ�dt$�<gJ,��Oj��v	WZ6�g*7�h���Q�	�>ϗ�Ǳ�DT�Ͼ��lE��g��
w�:��KH��8��+G�� ��7,Lb���c�y����q�QŠԥ��l��y�'��B9.�v��KP�t�.b�������6�;^�q�w[�'��A+�����;��$B^/�g�U�T4f��j�R;�J�o0�T4�~����O��Ln Y�9��͌X5��$=�yL�q2����y�@���U��%6Nx����ג?�V,��5j���Z�R�0M�3iv����mO��	�ra���v��F*_��"흜�Z��s���M�o�v񯚱�*�Fh������;P���b���:�Oz2 �D��#�� js��f `��<�z�A�u��BTߞ¢�U%*F+��zb���bQ�<I���/��@��b����z� ��_:$3cݧJ:;�2�,�SmmV%]��'����h+�_:��x?G��]�ҋ�	$J�s ��-)�Ft�%ŤƉ$h|��]�1���80�ی7�b�<�z��y�Ku��&��3�֬��=Ipa�V0HYL�e�B�2��p%"����=���!�����nYY+���X�����J��x�$(�5�(w�Þ���i	�Y?�:�<,:�%l�M�҆U�.!�=�$=ox�5��3<1��Ju��V��A���3�xQ�=ߣ�:�5����惮�����@(�C!B�Ȟ�~�)~n�|��˛���~؞)�	���b:��=�}V?Á�V?p՝���@T�H�Ѵ�q�x�1�%|�l��o�<�����H�'���HBh6g&]K]�Ѥ��"[���C�4�M����ڀ�qDt(�ħ�ـc���N&�1�t�F�s���z���x�|	s,��z5�����V�=rz�&��G��H�8N�V�5�-���#C��5�"� ����A]SX�UT���60� �{�U+8���BM'm�e�At�a2��ِ=eU���@���^��
d�t�E�.�
�2���)HtSfv*k�'�?�l��ب��l�pٙN��Y_@����T'�e�9���ǰ�B4��5eni��z�߁������
��0F��"�J�I�1C�L�Q���bO�Md�V�߭�ߥ��h� _,��3���;t�h�Y�����	�*q��ȳ�4��1�֢it�S��P��P�4�	�<�8B�?�P�7&�g@1�����xy#�i���F�յ�i���`(d��-�bm�_`1��Q$�^@���B���y�`�OǯL��b3=���j�OѬ�@��G�o��!�7�)��Zb�y�%�-iB�qT��Έ��㎽�<�,w���|�|71TCB�/*�tV��6a|�}-k�6ŨnoUO��'���kpY��~٢��G��#�o���F�������$e�0��j	��c�98�� &�s�9RZ]����)>�T��_��ܠ����~�C3f�4V�������������,9��΃Sy-�]�y,S����o��f@5s�ꗙ_�^D���.���0t$7��<!zFQ�=o�2cI���~�^�'���ܱ&0�hDכ�0��״@xL�>c����"�J����]�����vB_q��W
{Z��xl���c]4�x���A����j�@��Ϙc�v���Eoͯ�|B�!���%/I�E�ų3��"�ԫ��N9H�gQ�={p����	��mu��TC�y(Z��?�V�,�:���:���yO�����^i���V�{)�P(�=4����+��''�����Ɏv�pR6~qg�y�1(���+�lsq��BY/�ޑ0C]H�!��qX\1,�s�ˣ�8Y��EN*|J!���}N�\W�h���'��E9^:�-�Q�q3w^B��J1�}�H�#��&�c��*�O���S���2�#\��C��A���T|4%�1�YeT`��ص;$5�o���m�����՘� �ϒ9��S�I<t:�@������mk��2X^�*�j�@֖����|y�N�K*��,�_�	���	�4����Y%�;
�2���X���s7��m�na�I#l��&G����q�ށ81F�H��d�(`'QN�G}��ş��oZX��cC�-s(Р�,�4=_ h�6��^�\G̍'�8v^;�5�>�y����u�` K OX=۠��*��h4��8nYv��L���{����%��^U��N�Ѭ��C��H���j�}~u�WqKb���!g�22�佗f{�V����h�z 
�BK��[i!t\�����J���úq�ļ��G�sب�R���"������ �O�!�r��&%A�U��IW͹.�>��oSf�+vqA���17�n��Z7�@���A�۲3����V�}(���݋�	#�~Ț�P~@��翙��_R��	N�,r�	�fy�dWʘ�J�~���2�Be���Y��(�����L�@_Z��8�֧��ީ���|z���'���᮹Ա�l�B8,K�����i�͊���]�<��%J����������\�j�m��~	�5t煆�3�G��
��w�Q��8MOFm3f�b>��JT���D���WVnh�h �ܯy�@�3�>&�hFT�[��H/�<�h�w}�mj��-���<+H*$X�;���y�X�ㆠ������w�Ӏ#g������Y57�oO���i�i*��(B�� ��M���f��Ӑk����?ͮ�����$-s�^)�u)�����L����l� ���9�޲���5�-��)��\h|b�jm��M��o�-6��2wt����͆SgI;si�����V�_�?�!�	�s[�\/ɂ�����r�_�`7;��׃�4��]��/�t#B
M�I�"��;��1�?7e�M������� G��~Jt�T�%";���=��2x��#�f�Ĭ,�#�蘭W�I�ٿ��;�F��S�Y�3�O���!k}Q��r+�/ýpW��P&'��b�CKz+wz����>4_!C��Qn^4�E4;���>�&o�f¿�qUW,.c��R]F,�&u)�d�-I8�x�3 {5����P���/����qh�I�a4~m�ⶨ� ���.NY�W�k˷�ͭY��:���E�-G��2L����cľ�L��M�f���aHCޣ�6"�< '�uD*������jJS�����0���:����.Luv�bM�p������6;:kH$��m�����U�j���[1m�1��Ka��|�,g	����&m{�˵�`�+������{DX&���e7�D��RS���{MYIe�PT�x�����^��w��'�����v�έ���i�\ka���]/x�=��/���둬Y�oz�=��H�M������������X6�'�b�;l��2�U��b�Scj���y�/�=~�����>���/b
h�+Q�,�m��8�{�f��Ikyn/���w4���M���E���FY��J����J�Xk��"!�F���+�i"�lf���r�&�k�Y��W����p��9�<m��A>pn5f�K�� lV�]�UxO�/����-���i��v��V�v�J�m��%А�Nk���	�(6]#d�����:PF��35P�����8+!/��?�6�?�L=�|�Q���Żz>O�S z�qXޡ��2ǚho�-n���ݓ�Ņ��M��a�DV#���>���t"��?3SB�`[%T
Z��W��/'�τS2M�dD�>��A0�&���P�ُ��l�և���H���& f�A��ر��џEx��j��C��	v���*�2E� ���;f*ܲ�l[��)�	v*:w�l����D��(�ȭ͝7���5���9���Q,K5/z������7��ҵA�R��,w:ZEx���|8�~�}�϶�.�;�8 ��h���C�6�1o��z�qo��a�不X	�Y�
��GSP:��fȊp����!*�� ��ɠ��-W3$��V�2o���	Ra(=�?d1�f�XO�U�%ؚf1�o��1N_����g��#=,c��o���^c�`���:{RôHhRS ׊��m�z+���v�_u�Ǚ�\�i���lCIw���|A*��͚�e�B�����n�w"�<e �p���Su�
)T�M}:�y�����s�h���P�j��\�'��D2��]�q��v�f�4b���{ҭ��n
q��z�K���%:)ȇ��PT��Z�Ĺ�?�!���7ٷ��V�5��E�L����|�]'0`�+�XR�Ug5���خ���.��>�tn�z��</QI���d��8*�~�� ���w��X�}��O��g���D���9� ��Nii4���0~u�t��&6��yZ��vƠ3s�E�F<d�5�m�*U�:\�>U�4W���fR�
�����0{ٶ}������~A������s��xC\��>�㋓H���P t�k�B{#�*6
t�GG�W�wL@;�b����|E�]G9�eN���ǃ*zp�{�g�-H�a@ԖҾ������v���F]ӓ`��!�T�EC�iu7�=p�E��sG4,��+� I�;wP�1NR�*��5R�pI��v�X�K;���ʋ9�e�oя,��F��G����p,�����&,�M=sa%����a:Є2&}5J�{�ql�i��Bʵ�П$;rx$����aYɃ�_�]#�P�0�'�?4nk�,�x��8=��Pw	:0�1�"�o��Y�g�8��މ}�aj'R�XrbR7�
<u����xE�t.H�l�J�p[���poM���8�볙�Ԩ�0G�a�$����$ķ�;��B_�/�[1۶gJix�u|O��v�8��1v�Na��N]N�L����_!����� ����M�ͶXI��٭Og����c|�&,Ȗ��>�<���7�S�8�j��p!*�O�ϰ���0Y��ެ�� cGT�������9x�̴�:A-"��H���9�;�MlK�:�Pf�t �c"�Ħ+nİc�j����a��џ�.�J+���TA������
�~�#
�"�e�6���\�`B���kv�zs&)�KB
��΄�8���ޕ�a�:��e��2�wc��L,z�i�����n��^���m�z��.A�����}�s�Lf��`��I��)G�x{��@�]46���N��t�ܚ ��d �coɉ2;�7�X��$�;���<0��