��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�"Ivf��[��#����-���� �C������lNT�׫D=V�D�S��-5r**sw��b!�,3����QD��4��6*�o� �r>�a�6�Ē���Q�Ϙ �1���m��-\w���[�d�X�i�����7hYt�A�5���2����x�KEd��K3��/�]�C��Ĩ�����`W��o��? ��'��F{��������7F�����愗A_��|'h�جQA����%�8�۸R��aK>�.�W��Gm@}f��z����2�؋���m��\M�B��Y�\F���}��v�0�7ן�w	 i�{��݁�>��< ��Z8k�zhM�eO��o�B�[�3�m� Y�xF�Km���Kȥk�S,U�W�+��W��[��\�����I�N$ED�B��M�Cˁ�_�!��R9�U�l��OM��а4�!�$��D
M��L����#��!��_� �ES�������$	z��
_% ���Ά�?�,����p���p������O
�������}@Sއ< �}W7p@���� �"�1QsXӜ7B]n.�(����Q��p��:[c��>�0��Fn�+��!d���yu=���ep�j���j�q%t��ϯOj��`u��o�a�jp|}�t�K�8�&7�LNs�s�@�����ǹ�7	��t~�my����n�l<PT���x{�0B��7 b<�|�B �4���ْA����Ёѡ�l�Ic��m�*e��:Wі����Ot�)�K$��YI�³K���B�	Ě�S�5�d|D�S�aa���n�("�>�]��8��J�WT�V/����4aY~�ˊ��U����d���CU[��Cڤ������zX����T�2Y�$�z�˱����a�[��~'L��:�}��CK�/�'��)[��i8�@1��N��5%�y�p�I�f&���Z�Vf���Z/�)Q\�v�f� �d��O�g�}F	�$�e&\�L�V �!ȥQt]<F�Ng��ȣf�z�����Gi�kփ��j����w9�Z�3��5K�ѬK��i�fjQ�ڎ���/`O-�<�abS����E�����Ph ���N����
���m=&����Am�C�b�u��]}��J1�Z��o�����q�]�����u_6G{ްv:8-hl��<rF�h��\�O����N.K�Bc��L�r�o�������!zn��Lr@{�i���ژPg�E�K�ğ��ی7��YY� ���5�y4��گx�1�R�c����e�դI��q'U������P�#�Sn�D�G^��
�ۗ��*�}�4��ٽM�(6�&���#Mm���{y�	Sj��� =˴�fW֥ -[���r$�.�W���5+�v9��'sk������,26�����ƞ^��ϑ�-��.XX�s�xЪ?�w��v�7�CB��l�q�@Ȝ*��ܨ�1�8L�����}geN���b�.p��m��BLg���Fg��1�FxD��Fx��0�ʎ��L������ M�$��U��8�Q��Tyˬ�$�2��nϸ�����\1� S�2r�KB�J��n�]�>��Tլl���IS����<�]��C,�Y�YT�ͤ�,;!8��O���A��pF�	��E3OpV����xpF���������������R���w8b2�� ���id�kDU-�uf���z+�k_�g�&]?��u�8�������i%H8��B���3�5v�j"P��Y�̾Ę����+/������0�`\t�V��43�{��=�l=I�,j�\4��@G�T`VzX@��y͡�Y	G<��A����wL�*�,�� �|��G�b,��!o��6\�B�0���j5 �Ե̊k�t��+�սq/8�b!Ir��y�o���l���(q�A<�5V���)_�i��������:}_�y�Id($�r p�S��g��-c�;���^�"B��T�u�p*�"3�<���SG��������*V��eY�C��1���iJF�sO�vo�M��[�٧�2�d�[�Ź�c�Q���5���1&���F����S������|+]�n� Ƶ�G)����܆A!t�9cnY6[ù�X�Mn�*��7���<pl�`��d(��[�(1������}�TM�ۇ��;�)���n�t i�αY�)����N�Ӛ~����l`|���J�mG+��$q!9�$��ϐ4�V�$k4��I�ҶoM�WE=��-���E1e �����&�~.K>hH��ca��gc	�uk��4�=�-����}��D�:��Q��F��Cv0�M4��8��g��Fԍj.�wX-��N�.�^D���Dĩim5 �͚��<M��c��M'���9L=k#�pE��cΜ�#qIr5��@��������-i�s��a�ܩ���72��#ٖ�HS�*8��Pd����؟m���'��kl�%sT���P�d~G��gi��H�b2��lx�1e���Xl���cȆ�<�S)43P���zTnt�X�؜K��d��3V���Aj'�l�z�t�AP��Q��%�	���R���\b!��ʇlz[q ��J�z�rV�ή�l@�)RA������ö���|'�h��.V�����֤������Վ�7lJlm��ݨ�/�7[��޶���w�b#(O�
�(�B�P��mP��w���!��4�}Յ�o�D�(��O�G&�wQ7R)�R�%�m�X�|8��x��
%E������e��b:2��� �9>�����[�G�;��n)t�D4M
�����$/��Ě�/WU�<d���U�\���渍r������25��� �߸7Ͽ�]��P1ZCи^(�'���j��MF�AkE����`C���w/>������n��V�v�f��u�ǭY�l��g�9o��Q��C�!B�ͧ|*���
�d�p�o;@[�qi4�m�r'tE��b� ʓß3��S[�$G�:U�
���ocw�5��e�ށ�;[O�!
�љ�$�1R5�r������6��赧~=��=B�P�po�՘Ɔ�گ+s�.�<K$\0�ry�z��!����ŉ%�M�X�B�ꅌ��c6����"�s�y �*�v���qV������b���aA)��R�n)���`���Uї|MU���H��%m*��&h��Mq�@�D�(�?�j�ȿ�dh��+����[Į����?3F�E��_ m�z=[>��ƨ�~�|Mz�h��(��_Jvrޫ��DQ���d�[%�N��g�Й��ww)R���:�x�)��������}�7��e��q4�DO��SG� ��d�� ?ݎ�饉����科��Y����k�ְ���<�QBg{~؏��L�m ��[1k������Qe��Bcc��y��0