��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�k*b���f^��g�{u;��X�+�wE���:�ִ�J�B��ܿD ��؀-�(�.���2��k�aɸ�Z��p�II�Vp����Ё���^�V���1��W�����6<AI7� Z�QHֶ����Ԟ����h�"�;M��a䐅��ٙ:͕�0�X�iFf)'~~�i�q�;�{��S{6��%�-�U8�� ɻ+6�2N��J�}%J��ه��W�,h�@�w˳~�@��x��5n0%��֬MI�oA�}s�v�E�:��� �y���B�i+����<�DʰA�����Ɏ�2�|o"է����ˣs!�2�Epf'��lm�q�J+���:O8�w�u7%"��[4���Ce�}��Z�0����9g}\i��>��s'�I�v�0-��3�C8���j��+Dn݄竴>#�+�Ul)�B��?��0� Y�\U�e����"`�<@ۂ�Jfv�"Dy��r���Y@:"<���hTf�@0�-�	_Hܣ'�Zl����z3�����7���_Q�z�pQ�V^t*Ύ#f����"����j���
wĂ�Y�7�z�M��F��2}!M��rX7�5�݂!nRnT�����2z��%���'��3��:���w��	�MZ�{ba�@�蘼`Qf,���Ws�JqD��'�8Ae*����KŃߓV���H���*�8r���`��cP�+xN�7����D鷸ZX��W`���A��DU;�	������6�ځ��8e�}��RRP��1���mGNxm�`�T�k�,j1[^˻ �k'x�Ɩ��k9���8��7�s]�/]t���ϸ���NԤ=�V��G�/Gr\]@W�|Ͷ���(���ϯm�TO�G^h���c���nx3$�A��1��$�=�jn��Z���"���uE��#�w����+��
���
>)Z�ńL�2����)���m��C�=Jx���x��r>~GԈ)��"Řj~�E��y���g�,�M��A��CR%���zo���t&�5Hw�v�t��r��hZ�f��^�_����Ɵy��8��MT��a�	�C#�҂es��D1"���g�yU�k�՝E��/��� V��W�ͱ-'�xW5�����L^�8��=���)L�9�`>k"!N�4T��8�}8��;�*JB����l�T��e�;�u�e���:��L���WN�n)�K܃��)z�l&:E�1�n�Jy����X�T~R�`��Kp�����8ԱAe"l�Fo��i�c�<nBpk?�f�w�M��3��Ϯ�{�*�k	7Cm��\�4��XJv:�E�>x��Hikp�xU�������vM'���+< �ZT=��;Y�S2��|	���h�I$g���W�@����a?L��ˊ��Rg�;cR6����Y���e!��Pa���NȒZI6�?�(�t5�Ԩ\�{��t��q�W��-+�M����<�'j�� Ng�w�ў������������_�r,+�$�Ŀ��w���x{� n=l�ݖ�}�iCBBƜo�� d��(J,_��ƚ`o	q�w�����L-^Ηl.��o��zH3QӯYQ�+:�c;���'�+��d�H���G谰Q`�Sg�'E
�G�Ɗ^D���7Y����SW�E�QMi�b1Y�p��5F����6