// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:20 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nZ3r+xmFtVDIdgVhj7Qx/3NYYjqnyk+7EVKT+6zV+tDkF/22a7uSCtCeWkRXboSl
keU8PghLs40NIeMUfPOsHSupmsWEP97xRpdioOz4BNi8SX1bXfveiHupYJwa5HHx
lfMicaRYjudI/6Xqg72wE0xh2S+6OtBilVhkUvoLGPI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4544)
hQu2wjoOhTg3Q8CLROGX7WU+x4ifM62W8f7xKj/KmiQyCAHXBoLHOgAzLze5ypJf
wQm23XYb0q1YQOhF/SlIU1oNgCMapU76NFvmmsMGHa0RORJcD/MYewCZwdKqvJ+R
IJrf1q2vs9ZZJDnEYXCp4ADvE4QKrKTr6zzE9IdS6CpZ/aBd959CUqiHBDB7w37i
9UwL8e5yxlh9qNjLFJm76x2foIN83cWxFK5WNPBDCa/qc61aE+ie0W6JDTPiW8L5
6+GNXp5Mgiv718z4HlQL5YGuFNGw+Af2mnQd5U4u+Wa+sFeVvZWOUmpn2UncBsU5
eMjRcUvVlyQpDLAkp8jMXHpXLKXvqF5CLxXFJ6o+lrUNOMYPWt8o0sF+Uwd6RJ0S
Eoz/0SIDQhQA/d8AmnntndkioUbYkhpPoJXX7R++dlBRlBIvnUna7mAX66jszVIC
FXy6Z2OJanriA16IH77cYOEHH7ni/nHfXcNQyhxBLAkdl0+rpAXpyuk93hDVSpbI
U5l/smYZAr0AvRcHw+11/BEU6uDHP2T396EoxN4iEUlEr57+Btzqt37eEBsTV5q7
W7vx1FhdZGPHcjVfYtooUavtf6JKjetXsxQEqy8Cn+WWSn8xLVjBafRwWwyo/VpJ
C6ci3P4t2Ig0X+wFosde0E3uRIGzqocfy52vA9FWp7TtMOWweb5omFyXoLrKT8XQ
EdnVuQ7KtBI6AHlpz1bmDXdnxDj+tJT4Gu7LwuLyUNsQBOGMe/nRSfvjCcw4LzgW
ufCN3S/FVEKc1V4ENkoLIOolqiKo0ldDD/j+kHtjWMG6g6MXcgQL+hKk9rTKmr+W
H6zgYgLy7CIbKFVYMC9nOARO43qsx10yzC3/bSJ8zfe2iTqC+3xLRqiWDda+ygGx
Vm4YkUW6B7WL+CBXu4m35tWzR/b18pVPbZDqJCDvTN5mgJLd20x1uNAm2ucqyLqg
q+upE+fWGCp91oYSrCUYxzdvdp5X1W6pv1A58x07wcxarcJajxaW2tvt3LfPeqFQ
/RGGH+qsumF9mQzpdqzlu9ryWNh0FPkpzcQx74nUBADz7F+i9a7Dq0k7uNtevNGB
JgfhzHA2SJdrZsUsNqPkD8paisp6Rh1w8uFR+PTB5B0GZoEdM6l6jO7kZeuSn79J
zKlJz+VhpdIf35pA+6mO2OKrc1JOhlFxL1jzM2r0sBh4CRSbxWKJNNFMaqWbJifa
Riq55rJ297zLD8/tV6e8lSXgMwx7bYnUzraI5QPLeSCfad2z1FpxLBSMIgjwj2Bx
G1wldxo69dbDVF/As/CCN9Z1naf/lLTEVj49NbT92gYLVzUfHCL6DzqyTZnJE/o6
rvxgaK1B3SnlgQnDDvYoexODSVuK9I61RONzgu2MuXN1Mt+xIoztbOa/3rHnY0hR
kmeMiToPKFOrqqnoC25230ASqljvLFlWGDkvZdrYmngIBvsJeG4NF4aZ0oX+BDEr
Dz/rG+10cyrtP8FHmkNPZS78Lx5Hqc/YGZSxS/9OKQkC1/j+z2m8GGqslu93Fzu0
e3yNHIJWxP2viNhrl2WFY1FD5G54d5IjWnnEfFRNOkaIVHrNP8ACjl7jjAXL3VIo
IG7uGrm2a/vc7rkBKfS6VwrJ1mLID4EjSPNEagKT58BnoQiZinm8JSAQYdmkofMc
KHREu/94W1OQlmEntOo/46Xd0Mz0VarGXI0WnKs4vVmymLHfP9CMy9bBJ+hStxl2
u7T+Z17s4EzHX7g7WiAXFnqJpJcqxLLahxs/2mL2uqs5KtsxX56PoWKc8jEeXsxN
wRRFZB7d540VEx93OXXiu1ItrcgvVmKC6UAJr9+6Yco6p8536Se8iI5+0Q7FNehR
oVCRjLva2o+ZwsrakAl/f+kIL8Jl/5cbdVVQIOFCuMuDpGuoMJH56ABb0WhyBVyJ
EP27hHxZ2sF3r1G1EXbML79Z9Am89GtEr6vPaD2xGGq+Iovh1o2GglPAvpPEziJL
a3cM7GHw5E6GknHxuB7vNY5aZW2w1fXrlkUdCgNbRoT8/wG7bBtB4CrCaoEkq9Sb
hOwiPF9/+kcJJ4hd40dpMdgM81Pzs+duzYNG/Zz9Hig/rw941NY5zdFitF2itT7E
Phpy82dYj0zNkcTgX6IYERqJqQqWHLwVSx2NdOh3gXKKDExI7pSMnhBQJH2prfFC
YQZZs0UIdOBjZgcYAxdpTxgMuAiN4x6WKtDslBEf2IXkdihvdSuLef3/RWyne2za
dsYV9VnCjwYIwKkxWZoiNjiKBmrVVN0+mudJDQA3n9eoY/iSbO7NGiwOzsioliRy
EJgqXs+tUV6rEXqRyh309vmF/w4HmGByy1T9l/WCrcL4Bj5hzsPEhA4ZjN4S5aJW
0ysga97LLw3kkpQA3G+3arJ65DLHv19y329u9KyCKBXfnkQjxIo+W0r0VMaeCmMj
6q8pZKzPP/k5hDNV5GxlEprApmU4bPwZ7fSHk3GD/e/6Jkl8/Yaa9ls2f2MhvxRw
D4WKpjq8PXeeGfq3GQh92wTA+Vh1O16IIuhDKoEDhJmzggEVghL/E5UA0d54bdsz
tVYSHl0ExoPs7kI7HNfpo05u2TqXWGNGlxStdJ7K+qo8ZQ0lFPEZErp2IbBm57Hq
DyJMVzEY9MLi/vQj2O8TZTyKlNun785WCSbOPjvlh0DtBwEG2yT7patdmD2+JPk4
kV+auw3dlBT5duoHov8eKRN+oeDxf7OGT+v+kykKtWx0WtZDeQHxcvYCnPfWEVe+
1GO+0DOCGOJINRN2aYORPCkUkrFP5QLi8at/qE/9ismLwsustiWBt6suzPzGwNW1
YjYHXN25p8wkBoG2GxDNmU+N0Q3avfHyUHMTJbwKo5lYHfWonkO6jAQpXFuH2vas
01fprd33ofWSHaM2Qi8o8lOLhM/V7ovoFUPfyQB+Tz9279eFjJAc14GBve1zp3yE
G+BGDGTjunQf0Hla1me8ORBX+yb6qVbSnbF1U+GMHFRyzruDcI8zzxBZAizZjR14
h9TWijiwq3Te8FPMlsab4MJ/V4TmEhBOC+5hnmLSKPN6LwBs889Agfb7wkj7QwaP
vOHqXsBu2tBrShZqV65QKnJMH0bSJg8//2dPQujaSOKVfOyFNvpwg53QmUC6XFON
BIVWrQjEU+HCyFbGBZB3r30v4a0p64/tVXGAB7vO7i1oOcA6Xq1UDfWNChKR1qbn
pK1IRbKSGMvvGFd9x+Erb/0gMy/g/f6GK0jDUH6pPu5iV7uXaAHxrEH/2ErhujL/
yvr7q+oRFk3Bso+noohI1dP1YBnbuhl5zdBrLIiMmo8dQzelEJhL5qfbYmyPZD8f
57tga5AjjUBEofQ0DVuDRTPPS1kWYRdQPXF3R2JMOGeFkwrRHXJGZTDWenolWNOa
tRskNkHMTuJgy89fMWKVLq6DxLyuSP7HsBHotu2sjCA7I78cECLrdTknjqfuwTc5
dSLC/6nwLFoHICSQNiYmAv/GRXvcYw5N6cgsoELMjOABUgRNFuv4/UbwPSreZa9m
wuETVvmrdJSRwiE9lOQ8LfNPrwMtrgoutKi3UNAcZL81x2KbiJj9rvDbwtR3oUY8
wiUECWaEXVJy3DBXXZkM5Uz61jdyl+B6mqCRL9iqFEQt3qXS9qgsfojP2WVhJETN
qr3z430KiWyPzmZG+avQLNVjnZCrLbyPgYL9zJXElw28RHbUkp5eE3k04qQjq5uq
2AV3r3PDL6k7Y1JSxvPUu32JlvzoILoQztzcTkPDwK8+MQ8RDnSoJEQOLlNrOrgE
Qr5J01YOy7dRSbjEMt749/Lrbob4gmKsLFSvTCnxCqtP+AS/wNV0djSp1f67t2+u
fh63tbZAKUNwyuOfPIfr04vBCU1BQg+oqnQqmTC1GxTP3PTTZcxWNGcIcEpJN8Gx
JnhlUWeCkpOgoN2Lhpr0kuIPYRUJf4x/7WQDt+miz+dPt92AaarJMafqPv92g6tB
uvoDE6F97opy1jDHPnLItwXXgI3JW79uIY85rtem/p+jFiAZOEXzxXqKU5e/Xazx
J8AX11s1eSJ2+uu/TGggyQRi10p/gU9RGTBQ9jQh0bsnT7QesjL4tVbdbyz4z+6B
tcAPH/0ah4LeJaLcEoCTeQ6I7Gn7tkVyoh83PJZrW8YZD2djcbth86ZP5PybBdT8
Js0IyEmf4EQ28i+kiSJvK75TsOuJfh7IMlll1sOkJetoqKyqBAcFhJqFEKYZJYiy
n39e3H7hZegNCx1tKFDaau3gjkT7BAsMghs2BLZapCd2mXL/pvMFLYg/USjSbez8
wHlj/DDFGnEM2LpvRJxuKa3WPdTnnHGJ8UO2TYmCEFCoeF/asLCA0MKwgnuuMPk5
T5ELc2lf3HGV8q5VqFp26YkpUZ2+q0anuHHQZucHl/2AgKCdia3uyXgbz1OkNBpz
utAgnjVtiDB3GzlYbkQuazdqxfqkACBq88jgTyeasjBK/oUrmC0V614/p69e7MaD
skA6ACJrS6P4+e/Mgwwz40T9v8TsqG/CbPXejvhwwpK0hN8ogPNrfKsVvVuGPd0V
myhASgH6PuaKuzq1JDvywYkp/HkTZscTE7hKA+eVZPL/EcRs9RpymUaulqeQjljl
kiT7Em+KpiXN+kA1mrlnd1dEcMvBoyju+GlenuX5gPJF6IaW+o82l/VN0C4mWlui
/S/5yohqhWY36j2gfNAxfBmqznUrbQBUSokLdFrj+Wdov6gWjYXe40CN2xlMFdFN
8+iwxerXHAEZCHVJaQiJYoKUFQEijN5q1CbF7SOf+E0AdwIYWY5tdGBMk70ZdVGL
G9LwaNVPpgbalyQSHAl8lu7lolfgeV0xx8s+AmIfJxDusp2u8wGw8gbxmcXg0QCa
QnM+rL37Yk271hrvOkGVuN72y320TFUWkgd6Z//RirwzLf9ScwIwJhWqry8AtIFW
ueX+1YIaAQLX1w8mwIQbe06H2DQRHqzEDNbsyAbxctELyprZ/xF9aTpyfF0eytk8
nVCmn5+NM+dq7dgaPnBfaOmXjZ10KItEk+EEGNprZ8Jmcesg6xWPCc3v1tUlvWir
DBsODw7d7vVWrGxz3+uDPFiWbu9M/IyLYm9jyJXxwCcNI0bKGOalpnOPWc2ulE4V
0Yo1UBtdJ8dUM0UW7he5YfdBLqNXvGeweolBBlOqULzpfP9w3pp0MivK6zB5omtv
+NCMWhTjjZNxfhSorOc1Kb1eZ6PI8t8roqHH2LYAph5xjdEnmy7ZK2XrM9CvqCAM
bKq9tq1euJldoETbh5PlkbuHaYg7fazCoTIXV5O0izV98txe+HR5QULmoL3GMTEa
kHcu0jbPFCZbx98N/ruD72Jlaj7BBvP0iq1mVw9pADEZbN+YXkA7mtJFdsnYM+sP
0imx/811DJZjxl0A+CF2Pz5YnvT7Zs/DsRdlix6WXWxZyE/1pwEgZA52Fp7wF3tx
IkryHeNdHcOHG3f9ySD0A2pD1btNZ8Vv8Xw2kXRZbe+NDiC/7UJs9b3kNAozCWbo
r5Cy/h1xKQrAkdKezjw+4W6vRPM1UuOGaCNzFLxGE4ZgQYrgM5SGpgrA1EVNJ+qz
AFwBABkHkJ8txAxZAPYFZ+ARS0ityus8p2b38VJZUIxG22a8TX3vQo51IaSbl5rc
RlqZ/6cYzqTQE7JKbn8VwJhnasrvSiZNZeOtCnq7zmTHr9pvNdkQvIVown49BZVZ
EYsKgIMdiD/9F8j9ck8teJRIRnfwrZ07V6sn+QAWlHFeJAnfnpWg76M0k2M8a2lc
xRFCEiYPnvQrgUAV7hbv83y9vVFtpimMV8Y5oV9+S8+sRKgCQh4fWHHh8Mulz1Ec
1IF4vrhT7ITY2D8sMPIY2q66CVoNZ4i8AaZ34MipsS4K33NXm8y4xYoP7/B4cMTD
oFKmj7KNnrl4pZNMEUY28bPzAx8BKtGCecirDv7umG0/bgT/TuGROQ/kj6kJk10v
Oino6L9GYAsPfF2upyuRv6JmXQ16kzOYM9PYyQvnXpF/32TwYP+0IVFiHSIWGfif
SWT487otqylSIhYdO6dBPmO4+pqL069u+Wre1o0fJGE=
`pragma protect end_protected
