��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�y�Sy�;��>��&�MA�)Cʌtg���e�8~�����=H�9����.k������U��U�Xe���M�b�(	
'�m��_�S,(
>ɢ&T^5�[Kم~�WA��Mb�c#�<˃#:}��6͕��F��O�j�7���'AF�9��'�ƹrq�9�p�
o�'�w=��v��("�|��ӏ�I�\.�V�����)���cB�չ6�t3sꀚ u?�({��_x�W������!�`�e�H�H���|�-�YY�
ꆞ �Ӟ냨��e���S�kFd�v�e����y�*D���G�>����+�ᩜu�f�x�I���*��/1\1����r�2�*M_�4j�t�'{)ȳ:�A��!���ש��6�D`��Js�[�a�O[�G�O.�����}�9�����E���;I҄0"}̙�������@pi?%D;�4�]Aӂ �`
|ܐ�e�p3��D�"����F���O��vm�� �T���>my��N��q9}�m���є����w���Try�	��
25��	y�o��2^3+��s�G�"\�3������-Xof+Z���v����:�S�jXD4=u�A([��
�W��S�Z�j�gߜГl���3���(����U�TLO��~A���L��V�5b
�Y0[V�>�_�u��%4�d�:d�y�|�ڨ���{Ǭ,�0�˄���+	�!(=!^�'���5�(2�>8��z�T�0������Bz�:�4��j�&����v�����p�"k�[����]����h�ɗ��: �,*���<IY�5u{B�{�Dk�b*ퟭt���rZ���ĀU�������f��166=�	I��ҋu��L�5ߘ�,����{�1,/��.r�\A����X�BÑ@�vv��*(Ed�=@%K�r%@�:"�M����-���/��G)�#��5�}m��~��酅t��|YY�U>�#\�o�U����Z����s���A�ȘR��آ� n���Q���M*���ŀZ�>�K�9��ZMDt1.gwb�6����E__v�m8��Y/ԱtQH�vZrfp�|v:�|�Y���	7i����|}o��v4���6�B::)��=�#��ܝ�t��?.�I������!��wP�J��,�Ͻs�E:��I*�ֱ�7��0����ZҹRQ����/�=+{���2�j������R�11B����Ѭ���MyNz��g]9<��9�v츼�-�4�����A�L���YG���LE�cY#1��1�W���?�&�=�(dG0z�$�Y�r ����4�ʡwc@����� �*F`�7y���17K�����⾇��^�hN��4��:P�"Ap:2���:�\��������^���N/�#bP�E��K��~�d�;�9��1�t/ئo�]�7.��PE�!��3|E�	K��:���N��F�+�D BCu�����,���'\Uݐ3�`�W��xc���&߱/��p�^/��6k)��L����1� φ�Ne��@���l%����N���5�Q� F�I�Z�6C1U��6Da�@=u	
����mEG2�0Fk���V�ܭ����;L|� tĠ2�!�uT/�=D�O�nĤ���:R;���q0�w���a�x)��z;d�B��T��/o@�v�@5�����#�փ���9��O&�g��Oҟ��<k����"�����וe�x3fGy���������Ҷ��?���m*���m���$�<'��#�X-��{����W��QYO���&�]����n���P��t�M��0X��"����2Y�%�"I�w�3�:�!�k��m��vݎ9y^��͟ז�����gQX�ѿ��Ȋ@_�w~�?�c<ք�(��8Se�C� �q\Y��� ���k�8hz<D
i�J5�0�U����>+�(F��~qu�L���P9��ᾰ���V(�x(�����m��;YG���y�/t�_��Z��'Y�V��-v��(Q���Q�����wj����.����
�)�
y�,�N�>v��/��1���	/�|t󠈖b���'�e�=/+��G�+6��(=\I� ��0��4�vQ�D"R��a�q	�}	�u��'��m������N�&������ˮ�z��B�����rj1�����tZ]�,m;�cv�~�N�>�S��(�9�{�#�ґ�u�s��V�QVݮ�cś�m4[ ��d�B!���Lӭ�&޻iI}n����j^�=�~�R��b=9�¾W�@*=�)�آ�z���[Kɟ8<�W�&|�|�X���X}�me5�#�v=m�* z"dT���X��L�o�qaζn`���QP3` ~4��ժ\;��W� �C�u�R<�������a�hx���)�uz�z�`����Dq��Q�1��|4]���-�j�?�;�_�,SI�� N!��~J�4F��&�6뚭��d%"�9�g��P�o�j��V���7jl�boVõ��K�Ɛ�]A��9R3�bD��6hH�hO/߮��U��/WBL�},j^��K=)�,�f��Y�=�	��ҡE`�WDg���-pd��d�'���)c=Z�ݝ�<v�)�4^������]3���֏�n����eJR�g�d�I=C1Zk�[��h9��|�b�X�{q�(�h�wsM$��N��