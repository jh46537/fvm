��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽�����Z���i$�?��w�Z�2j|d;�����]��W�>X��'.lg���빒Ņ��(�>�Ss���p��LP�L��&�l�pg� �Qs��G�3�L���f.=ZX��=�*�!ut�g3��U�|�p��q�C�X�\��G��r`��ut�2`�-�@>���k5T"�H�]%T'c>zf�����	gbm�^��8�tb��I�X���t�����ص���zk�s��2�M��h[�k��F�۹�&�̎v�A)�!�����Ǌ�L�=i���X�e��":X�2浂?��'���Scvn�SI�r�G䦄W��ٌ8���|��z����b1J�,�h�#��4s�_x��/v�f�V���0��&HCl�
�:�)0�!�\|����,|0�^�/��c(������Ī2�ӵ�ڿ%:��i����-���������g��9v.�l�ޓ�ވ#ks����D��B���
E\�ǟM�I�'-�Abh��|���� jv���${/�p0��l�zXq��;l�y�W{"F�����_�s ���ٿ�~�N19C�c��AY�~pk�)x�6<�I}ܧ�8'=�V��@��ߕy�hi�U�%_�I�Ԍ��9qn���@�g�0�[F�
*�)��ԭ��7g�J~�.g~���*F�_�c����VI�r�5��K�_�e;T�Unn�5���Z�vrQyc�橃��QvnLl�a�|&�o���-ŀ�I-��wkm�u���.����)��n
��J9Z��T���5\���/��91P�E�h}.m�Z�7����j�����jzƟ>���|q��w�!��g���9����4��a�1����1�����y�L��φA�$�v�����8ԟ�q�=��Ȅy_4V=B��4Ms�`J��;)��s�X��' ��.�Vʸ�F���3�]#�A	�����<s^$ږ{uZ�MM.S�_����U���*��^�S̞��_��V�/��������[��L'<�]+l��0��vw�������~vTb��	M�鰪ڹ��lA��m:�
f�;�4��,Q�܂k��[(�1��H\>"l^oZ�����	����B�|p��9~�3�[��/���(K��m�Ӓm�d�=���>0�ʲ-:���S^4��s	Za���=��[G�6��K�b��\2˖��/l�Bz�z���"OF�ߘ��c_��J��� _G��v��[�pl�8\t���t�����~�`�G e5�Ж��$r��6�b"�эtV������!j��4u������2�����_�t!�g��������-�]�3d��N5Fh�����c��Z=mv51b�����Za�͒m��P��':�t�6���g��ҡ��4�04�d�)��m'n�C�6����x�-U0.�#���9�Rl2�di��\-�l�"/���þ��_��
��.�;ɂ&[i��ʖB�"_44���ޭ�埙P} �>Ԃ�z "yP?�����\���9M0���8��cA�CWWu��{���l�D�-0ݺ�̈́��9�1�k�ğ�)e��Q2�}�W�cP|2]��p�WF��{z}��]�����;�9Sl=�ld?�g/���wn����\z��T�"���[0�4�.?�p�@myp:���~���b'ͼ ~�frґN�^�v0�/�)`����E��Ep�ʤg���Y��������< I\X��˾l�5�G��_1Fâ�����L��E��E$ݘን�c��s7��J� ��7�z�A�jM�d�?������T��dQ���[X\�W�-9S=�x���K>��*ĵ���u�Ǵ�	9���re��ו�-��ǎR}�����և��$βԂ	BS]�8Tib�&�-������?]K�]6����;/�+ұ4����Į��p�v���4�oȲ�OpG@�(�9+UI �[ݾ؋yq-�D:+j��ժ�k���io�~	}��NTX�$W:tO�-;ʆlJLM.�F����|�\����D�+�O�:�U��_�g4��g�0��~j���gw�+�7b���DB�7�<�<�g�Jf#(}�����9_d,��	�|�qrV���@��~,��M������]��5�c�b�����Zq3�'�Z�����3�o&h��M������j�	��A��zϺ�2��d�p��6��J�������	�>�iD�\��N���5d��I_=A�|��.K��UT{��M㹧�z�熳0����b9Ц��.�a��y��{pP���>m�y5z�# ���d;Y�=3�c#Ԍ����G`�M�L�y�]Ka[˴<V� �q>��ϊ���?M%\Vs�`q�E�RF�U�m�g/�T�6��4�B������֙t�\ٴ�|��
�̑_�X:���q�.
6�젖si��ɽ�ˊt���[�Tmˋ;���\�E��2�[�K�
�g�y@l�8<#
�3v��E�q�O�Y��A��XCE�v��f��+m��~��� ���)��Q����z��J�:&�o��|����[?i�#I��Ȥ/��HE���hBr��x�^��<�����{b����W�mH�4���_�����K*Or=sGU������c�y&��<{��g�v-�=#�yŊ�����*k����'�ȫ�hs���v�=����g���8�b>^�j*��)��>�U@6z�TŜ�hV+Y7�=��ϙ�So0[�0h���+�_�?�h`�F�/��2H��K�'{���M���W�-����^ށ�~ľ�sB����6���m�v,XmO�1]�".�1��(.G���La�������GU������$�X�X����J�\m���/Wq/r�jnP �U�*]G)4f�*@�ցW�A�(���$cl��D��ֽd�6�[��x���eN<��J�1�s*�k����vB<�H���y���V��k�q09�SP6 ��F��T=z�^54g��I�o!T����F�#�S�RR�{���� =^��\v�i��*r�L1Zh&_޿�V�~Х~W&X�d��хČ��R�z4I$"m�y2ߢB1���Q�Q�%HǤ������n+�G9r���e��m�t������!;Vw���:��5��hc�؄�{h)��i�3��\�V�$a]=�wpYUžɊ4�Jv1v��/H��(�[~�9��Si��Y���(5��c����G���3W��^���>���ш�Y:�7��H��5aW|��5��4lZ����9�X�Ȃ����qq�� %`�����z��`��?�N�Ĺ���%�[9>e�.���B�ܢ@P	(Fj�;�C��e�ɿ�E��́>�w�87Q~R?=��ot߸"�M2����bF_s6��z"�L� �!�A�3�Pg��B�бM���|6>�
9��kg@��s/���͌�~��l�A>�����5K��P�����g��hi��I;�2~��C�d8$F-a9��
�Yvz�ǂo~&�`��"�}�
yl�y�B}u��2�t_�&:b�<q��|����y<|kz+�S:����6>�U�PZϓ��[F1'K�z��U���<8��4!%�+*7�
H�Y[�
+�|��BGe�����ށů����vu��*��s�]AT��	�J��-*���<49�<�*ϱ�)zϼ����U��M-/����&#"ePǋN|]�п�����2٫_m�M?4�V�4��N�~���˄w��8�\�rs� W�?��^P6���x&RSS��'�xؚ�Ȓ�P��`�s��j�T/0ļ%�ئ<*��?�
�_�iJa=��䪝�r���tq���3v�|���O��s
cr��)��˵�53��.s�,8u�#lm�4�e <A� �RG2\|g�\�<}b��X�>JkX�ʵ>ʒ���������̺��m�<)��6�X��N�!m�Ax._z�����_̱M���:<��}��/9DRg��@��1�Ӆa��M
�=��y�=;�����0/ʛ�q(go��I,�])���\ni�Pxk�Hu���"j���y�3M��� �ɂN����d�����W@ڀG�U��V*%^��Cx�&��^�<*ƢDL�KC@91�Ƚ\)̚��	J�,�2V���XO?0nBZ���A�
��G�����!�닽+$Z��
���� 0裹�r��DU}�$��(�i��+=�@"��)�D��b�Gb��7[n�ZJvԃ�Q�S���i�/ �@%KT���xD��"R̄��#��:��u�l��'b�h�:�����SQϹ���a:�B�J�� �AYr�G�=�|mҊ?����J�p��x֡*�����:��z7>ii6�s�:�`����?>a��rmN�D��@�	ԫ������ΜF�3��5�i=)5K@`Ș�`ه��yIi������v�_*�h�c���'3Ӛ�˅�7�_�h)ɾC�"����qݩ�o̚�'q��+w�n�t�Q�]�0� ��	�YMga���%J��ǁ�/R��A�*#�ԭ���I��m��UD�<,2�Vc����/,�X @%1���(U���}����8(��2�N���Ư:"O:l0��.��OЁ��?��2��yb�j�'��1���TW%�Y�'����u*!�A�fp�Ǒ:y����9;�jHg��|�X'W��P*J��d�^���~�	 ZV��܁	�bİB1��Y�qi��a=� +��ũ�.��sC(=�5�Ƅ�0	s���Tx�Y��j$^Āt2����9m��H��ܖ0;1@7P������);���Pa���j���W�	����jsu]i�iZ߷�d�6�u�5oA6�s��)u�I�%b�K�VA�:Ɓ�yy�֙�o�X�����%��k/ЬfMj��� RZ"�����z���t8�Ώ�0�[���$reU�D�4	TC)���جVn�0�[r�,B7��	�"�=��h��V��������|��\�6ߊT�l�ӧшā�Z50����}�&�*�/�G���S0�θ�x��[P�4��zQ2����e�e$(�����D�J��Q[:I�Ρ��=[��X����!g��^d2�"��D(U��s�<�v�������m�q �ś��2���A,u]S3������-������tx�pt���3c����!�,����c�M�~���~t�G'Y���8<?Xrkhm��[%.�Z��$�>�C�/s�o�-r���d��/�
uꧢ
�z0jYĢ7���<�{ט4�b�Q�-.��>��}��.�D�+��2o��@�Tb�J�jj_�r��2ζũy:�-|š�>0��e���qW��ǋ�rG�R|9|�D��-��u��25�'��s3�I�ޥb��J�%CL���I�kޡc@ͦ���ng�(�_;�Z̭����
T}(J!g	N0ˮm�����ת_C�=K	�@��P���
��6�뚯:'�J��~� �jma1�5�`�{�D�H4�]��/%�h^��r�/��P#��y��Y�����juv?�5�gu�xO��;5��^]���-<�L�N��!uv�4 �ٷ�+�(g8������~���o�!�;M_d��h�:\yRm��3�֒@;u+��%|e��f��Gf�7�W�|�]�_	��g|��D�5�#|��1&����'@�Y[E,mnC�u�"^�j��M��:�n����r����*�$�j�����R�_�i��Jt��n�^v�〨{��yp�u�M���RA��Do<S�{{�)�~�FV��������(����#V�U������&�f��Z�&� cxz�m�2lU���	A���D�jU���a���>�&"^V^V_����ލ�n���W=��?b ����,�6�՝�a��Z��=�R�la��jػ.^#�vq�\�T˱�OT��j�C�-�
���aj���
{�~ڝ���Q�����F��\ΗЉ�3�	�H�j�^�&63��G��N����ʬN��H`�es[:�	��o�1A밒ib�����Ȅ�<^�Q:����G�] e��\E��,,��w�Z�$(a)�Gjڗ�WE(��qpqr��t���h������ɮ��0"f��J��q���}J�M�8�ʴE���|� ,6�Z{��a�5MBK�7$�f"�4tT�#�mKn�/���:���خI���n'4�����c�3]����Y�;p���<{��h���� � Qj�B^7����u�EI�5�;�E���t�����
.!���Aw�PO��f>< ez�cm^6��w�q�N�LW���|յ3����bD�V���x��'��#܉G�WV�˅�Z=�-�A'�f! i<V����os����N�z��C�;mbDKؖ|�Ц[fR@���n�(1F��0�=G��뿚��!���c�I����4���&^���jUi���S��\;��Z��:ǧ�G�U�ҡ��5ܤ��jw�f���f��'����Bd�����&�~�r^����6ก �	0+S7��3�3Wi�A}q";���zW�2d�P��m�ѕ��>;�����BS"p�BO�9�1�<�3�pD�uD�8!9��Zj���������;1��w����~�!\]<GI�R�Q�n��w,Md�\�&��*�.�y��A��^%��v!^���b�$�((���=����[���M���چ*����9�C����)0grV�f�R��&��*��W�C�=�q�L��Y�Q��9��(�h�D�Р����y!0�<a�"ӌ�~��㵽��1�H�A��ͽ{��^w'�]�u��ʥU|$�D��t�b�L�,l����ޯ�]p1^�����%�e�71�S��&H�dy(Ԡj��Ò���+&taM��Ծ��~c���D�*҆	d4������f���[�!S3!��f�{�%�k���6�"��[�i�<���~�`�HssG�H:��B�����G�t���۩r�,(��><��BZ�Hm���H�KW��Z\�8sCI�w�l�k�p@�;z<��eے��_���5)���?�˪��5�GL����8Qbk����|�,�JW.��`4�&a��Y��8����tuX$�ʯ��������m���u�fR�[���\�Xn���]�\k��'�N��XV<�=�XPӓ܂�_*���o-+Rb���le��c��v�B�Q��gP�2$
�l7��@E�켻�L�@W
Vf�!�a��Nm���C�_�8�DId��;��8�~m�Tl�9mmK7��1�� Ɛn����cȬ��[Y�����?���(���,Ktt�[*S�L��b�2�ryyYY��S����Kg'�쐵W�E�q�tυI�t�<��W�f/��5��%U�ezI�!��D,��˿�^��g�"�P�����u�X 5��ߏ6��e�U����HBv\���7���ƺ?��
��b��Wb�(=~�4�^�ʝ5��V:����@p�^��7]V�2@��A[���A]�;<z8v~8�&El"�$ ^�i&s�ܫ� oX��	��.O���T�Rc-�
v��p�R����=��m1�i�X䍎��b�.&�5��&gz9�L��ҋp��+N�V͈Oܟt�d.)#�A�F^�'~���9;]���=�udT�4�&#�zV���U^,�߫~�A3t������%��ƏV/�g��;�����$�Q�!�/���+����F�rF-(c*�f��i��D��]V3�3�Sy��D�*����	͜�Ka�8n�ʀ�9O������[�c�������^Vd���~�L���&����+�?�Y$�2�¢�s���)N�]�\���X]�5��m{�ʽ�G�q�%*#�Pڄ:�:Qo0�G58$��N�N[��N�O��JX=KQ�[5��SM�'�,D��[3,�j���r�x�A�&������BI���J؈�k�H�Z�f��|��Z+��C ��(P�#�h�jO��#�� 8��[��Q^��}~�|Q$��������	Q�Nh�d:~@#N[y��z���@��=*OԾ�[6���k��5�Z}I�\]�ƭvZ���9�Q��UUF�L�w {�8w�lD*S�����N+�*P���60�����ĉF	�DP!�)���m�Og0x�x\�GC��{��f�z�k׻�TE��_QS�0�7����f#�nv���$`�cp'u>�mr���ϔu�Υ�G����z��!��\5�cW�$��}��?U�i0t1��]�0����#�Id,��e�p�)om� x���]'$s'+�]��+����@�ɉ��MJxўot���+��l_)�VQf��kB����Ek��xǙ�M�����Lz%��8;�B�sO�~�ٞ[Y΀I�
-�lx��,)�̜"³��?z���;���z�+��Cd���&��M)�D������P�����v�`Z�z�)T�S�as
^�0�� +�j����Q��0����3#���@�� e��@B֡tS��N�-0^��`�{�[ ��`�ru�I$�(dJ�"�r�Xa"z3�O0-����#'�Gۖ]sl�Qz���霼Q��ӣ�ɓ��;�S��� 
�$Y�qCe"W��{��Q6�iz[�=��>��� ,��1>��r?���e�K�c�T����V�3I������AR�>�|H�y��
�ӧ�#Y�����)�s��. ���s~�3ۤ���E5�%����<�-v~�"�����f�X�F��o:L��Tw{���� �Ac���W�K2�WډY~���zk���,l�^����v�;�O-����,�5!l�_dD��lqI��9)g�{DR��D�/��2��"��_�D�+�w�I�����Ʈ@�� 2%Q8��"ߪ}j��Q<�y�)� Ś��^u�G��������O{�4�oۂ���}�q���S
��d�<�g:�`���a^��v�隭F-,�u�[����Fik�e_���$3H
р�����}�������R��=�����q��Ār�N���n��HC�v[6�.��ߌ$��81⦴l`.L��b��
��L�������Ҧ�������>�W�\|F�/�G7� %���q�|���.�U],��p�Nq�o9�k�`}b�[,��.�h�w����w��~v��2�0Ed�m�h+��Up�vײ:P�G�+����cёfS�-'M�v���lƱ9c�.����(������ٕy��������Bm�_F�����Ċ���r�(!���u1�-���'o���;�	���O���&�ƣ_��^�m��\9��M�� �����>�7
��0�G���&2���P�F��/�"tDN����<礪j��۷d��<�U#�,��y��aT�k���+.��Z�NI���9�r��ٜ6�b��04F���Bª�݁*ړ�<����@��Lv�T8����|;Vz�����v���p�,=<UĤ�}�̷�i;�����
��G �h�pIf[d��%�T�~6$���JU��9:հ
����� ��^��i ����|n�˓�ˊ,�ly��Jwjd���Ə#�e�U���N��Gp��̚��������"7$)U+<s$=�B�{�G�\r]yR����T1�+�3�Zi���",b�A!el��d�F�Nn����'ɱz�ypY��l�ֹ*���{.ݞ�M(q��rK8� ��s�%�ĕ��H�z����Yg�Q�Z�U%]�Bȿ��Υ-/�W��Ü�B�ur�o� K�_�*i���OyU6"�tn��1�J�e�7m�t�v�	�+�s�YW
:�p/顼��uE,4�r����`��G�r�����h��_�m�}�J\,��E�Y�R۞�d.w�M�D$U/�y���ڐ�Hsl�S>R�����ek��\����B�޿Ƶ���"9���>�.�,�2�؄k%���&��spm3*��*ٗ��W��XMY���T��P����qK�T�����9����،�� _���o�DC7<�K�žw�r;Y�_����")���{�^��N�{�q|57�� ������ܲ�L�����.��"���H}���t����䗔�t��̜�+
=>sЕ��^��o#Υ�pg�.�IN*�u;�]�;\�yP��]t�B �Mb���L}���\:��������
FN��S=L�O�bVU��>�-��J�O��5�?�2GŤܙ�
�v~�q�AU��A���V4<3�%R���̗��?�|�d�	�O�F�VN�kmf�Y#�a`P��|��Pfѝ�lE���[�3&��*�5Ŵ�l����S�bܟ����3'���ĳ�L��OI�@өp�rC�D�&��50��+w�2rխ���~���֌xX��̶N�-����0�>�\`k���ydP�>�&�dT;6齠J<,I%�tF�)�a%7��#*x��.l�'7��Տ�� V7�T[��襄5�A>57����_ӷDJB4����ׯ�nכ�����P��(9���-���ؒ� Q<dA҆����k�{b������*z���K&;g�>�ů� ��*Q#�@]X(H������ s8#���r��-.�	�1*a@��`�9]��g>pnY�=�t�V���QȘ�=���H�<�+_���HM-A#l�2�h�^/��M	������}�)
8��՗��(#�3���a���D�"#�%vH<[�P�FR@A�;�0�z�#QKX(^�{�Ϯ�C�8]R�\�Ą7�	-�v��Gsa�$��@�-/�!n�
<������/ci�/��dJ���+O�vN�Ȉ���`S�O1��I���GA���n�.���Ӧ��w-,�#>ϝq$j��̹����r�{��D>����q�I��~�Kܪ3٤|��� �֓�	�\pNJMn̤ ��I`��IF�ꎓ$���<c�xX+�{w��%��̕u���o¬�{إ@gP����4���lΠd|��Ξ��$r�=�4H�ݩBͽKb|�c'GO'\%�á�n)Yh����uZ+xD��0�8*8;�b��I.2�Z��e�g�iǂ=}؏bp�Y'O��aE�="��w	�18�����Q`�ϑ�����)5h�� ;Yv=~�ԩ��>4�|�	q�t$�����;{yḋsG�!w��
�	^+Q��b���9爵}�u��A{ˌ�����5���]�\\�O"�Z�����?�;� �@���nj�g��g��Mڌ�W���V"�An�C�7�J�m�ʐ�X��|�u�Q����gEVhM�4�QR���J0M"�#��J"> Y�('~���7����;6Y�4�[�f�ª��	Z>i\�JCY�b���I}Q��������!AS�S�/��_~n.HëGJ�%d�i���%Ţ�*&*���[���i��x����O�M�Y��I矓��� �^��#�+���Xj5���9��O,*Fk�]�
���]t��sA��D0fi���*�*I�}���̉H�L������S������S믙á}��UΞabh�)���b���� ��d��&�]e�Z.{#��ʁ�5�]�-�� �Ӊ�{��Sc�p�<�p���	q°a?5���y�.�������|9ʹ�އT|��}cz�F�d����>�g<G~�'߷�	�:Z�VO�'q^��s���7����O�t�f_�b)�эd��R$*��0v�Z�['R�����pK��S�_��?��O����tGb:sy����8����>����p�-.��K t|_$��"��(��V��p;�Y�;�����:��Vځ����V2à?��Ƭ�0dG3-��k�����@�+k�'���0!K�Y���'�2����27@
�=��:Yc���c|E&m2��~�r��� �k��b�
Ŷ���}ݩ�	k��Aʦ�>��R����Gj��Z3n�ǀ�N �`�"�8����T�Jg�n�Fٯ���/a�t�A�S2�3m���Kcjަe�@�������x	���,2�l?[�:�PB�d�ZI�q?�"��t�O�@{��WVm�$$��w�X�K�����l�"s�`-	�����I�x�b��%��|ԛ>��c�=L�ne�=�P��GfUUn�?t)��v�Z�X�B#}� W4J�BkRMZ�p�&v�]L�}�Ӫ{u�x��	c���V�1��}��z�%"�Wߋr��0M��Ǯ�����14$�P7�6�e�l�H��0j�f�>�)�$�����2V�d��R���h�GY=N�~�T��8�v;E�7v�g8���X��Q�ICf��EX<a��~=ZTD�����c<��j�{%� �.nv��C@w� ���f���w�!����� M�hJZA�JZ.��^_H��a;6zr���q�m��B8��������3K�x[�G���҆	�Z7�|���� �^�C+��|����`mY�ƢF\:��
2�@`>�Nmz)��q�S<�����A���Ц�F�\�����@k�m�/B�]������X�Ac�\f{q��G�&x>tsb�6]������6���aS��%�,�e�Ȉ���/<M��7$2���[M���ʻp���v}��{��йx�pU�#�A��#����{��,�Y��A�y�S۔Ļ?��Z����=wI��8���Ǎ��j����myQb�r�;:=i����*�/2F-�s�	e������t���$e!|��t�bfo����E��҈D�F����C�����6C7ʏ�37S�g��Jf����X�$#�IBKh�;�0���],���%�,á��iF]͟��n5o�Vۈ�#X: ��l��5�p[h�YNi���R�#^��ل!���(�NئO<�2˜�t��u5&������k���8��e�'<UHG�m�4z�'��x��G����)f:b�C��2i[=�]x��8�	����) ~���/�}p�U���3�A��+O�Peۚt�Q����0�ReB�����a?F��t�2*x�H��8*�_x;���u;�؊���!y�_=����:�ÿ55�B wݎ�q� �9�5���'LF���3��f��u��PU_Q����]L]�T�U��f��Ϻu]�;|e#�ل
�M-51�����܃T�8�{ �jջF>|<M�v��V%`=ׁPp�y�\t��k�����4S��c�O���I���`��g���Qè+���I�P��;���Z��^1��ò8��U�������V�H����ħ���_��Ad�������I�e7�Um�s�z���Ǵ��?w�^��n4mќ�+�H����z��p�����4��k��o�0o`NHi:��>�u�Nnf��~\2�ǰRh�b�+�\f��io[�	���ԕ��!z�a���R� �H�ړZ{�w~�p�sqB�O���4�m��vW܄^�F�7{qj�N�Q ��a Ws�3�%�M>�;�z)�����rCQQ.�kF�
P-y����Y� <S��6Fy����w�<��e�S���	o��[�
�h��o��L���]:W�ι%u{ ?ũ��'��Z�;�|�P#ߟ��wW��r�b@wx��0��՝��ጟ�jQ˾���G��!�oL 1���t�K�.HS��A��M�y}�,1�?T������0��A���D�����7>�\?�-��Ѽ���4�:�����2��<U+Y�J@���l,DbRS�W�6F����9ϰ\\�JX�9��v�
YH�*��b�
�DPz��E�* �iӦC1��)�cG�s$�;�s�e;$zt�wۨ�f�:���X����0ų6-�<�V��`�Hc/}b��BLϳ3��К���/�(��^��&��Ŭ"0G������� �1�jj3@(��&��e���nЁ�ܚp�L�����������-��j��yJ��&��U`bo����R]C�\�m�#ʜ�"���]v��W���%|�����������Q4=���n�V2���3@>����$�֥���iL�'��ēܜ�����m��Zv�h85���T�E�^��G��2�rKb\}�O��J�����}Q�T1v�	I���V�J)�֚�������V���ğ~�+ƈ�vEl���*�f��c�d�3��{ca9��,����WVo��D�=�M�qIm=�b�5�=�߅���O�gOˎ�~{�C2؊���;v���g�l�K6�T�S�hÈ.�RA��k�@��i��P���{7(�݅����T	�����Qg��]	oOg����9ӽ:O�7���-�}��c���8�&"h�{(� �^#��AB-~�Z��:��> ���T��>r���z�$���`�%B���c��Y㭀�^s�78�<Ԙ\�r*7�pY�ß8���e����.��S"��o�E0���':��;x_�'��9;��Qoںh)��{�������|���Iy@�$���~�ϠO-�[6���n���ɮ��H�[,���E�1Z~��f�u7�� ���&�o���*�@1�Y�	�3��ѭ�:�g���M9�,�iz�q n��1%�w�����2�1��V̶��7,��Y��qޙP.Ҿ��4����R�'4F��������k�_�e�;�q�DvU�S]��Pi���z G�_����R����{��4Kaj� ��\�\C��WH����9���񬗇���!6|�|������GE&���>���pܨ�����oo{D�,%��v8���W�N��Jo x7[�H�#',�����wC��=�Y�ҴW���[S���C1�
�L�x
���D#p�^9kg���6����dŧꐯe?��a��*
�"%I���!k	V!R亻[Ѓf���`P*�������A'O�_
M��e���Q��Z]$(CX��"`^�G�˓5C�B��IYH�6��4�����G1�����qO h�f_]�|�mI�������չq����U��%����年z���7�]Y��K�ڄ�!�7#�*��:���Q3z�e�"I�,z,X���O�n��}a^��s31`�ޠ��Ė�_ʨ>����x_zS@[�S����DH&��X���l �)��-R��21�rx�ـ��ӝ;e;#!�Jl����[%ˑ����R�r\v��΃�b��Y̥�k�6�y���<�]��wV��An(��(څ�C5��d�E�,�n�]!��c�ѿ` kxβ���j�+x��sC��O�G��c.� K��S�T�.
��d+��@�6˟i-8/'.�#O=&|"��F=۵�4��[�fZ�nn�� ~����m��R���0�ހ^�yC����Z�l�<S��Dg��; �����$��so��V+�\�f���}�.� \�78��2�T!/ �١�1:�󅠑�}Go1.L��7�!d���n�����GT�}-L����ӗ�C܉����ѴDbBFy�K�������zV(O�L�i�co�+�9WT�3�Y��i����+1pT��*-��#=�	d� Z�;]%iOl�0EB����������JD��%�h�R��P��\�l;�J�cp4����f���7{3|�}�[��n,���L��1�)B��Y@�p�����Dۯ�/�Fe��Չ�/�`�S<�I;�t����[z�]m`9:��5�J��H]NtҾ�����[;"Nrq�Z	�pK��n�5�z׬�X[�f&M:i��W+��-�i� a�.;.gIVi�(��헤:��q�a�n�r���b�CO7�Ϊ?��C$h�'E�0�V)�#{������q�@�R|�ẢZ��OL�c;��{v����{���>��z�.L7f�RP�	�vq*�g��r�EZH&S��F��YN���vNY3\׵;W��Qxݸ	:��E���z���������$D��M3��G���n������:?�rI�8"���=�� ]�TN<(�Y.��B>{��po�����&��o�"L)��&
�=�"
�	���Pg� Bb����k׆����L6�	�������BD�j�3w�P���;�nGA�⽩�Yd��\��?v��Z��̤�0�9��ym�ܲ�b(_��ᘷk��8�n��~�a�w�:`v��H�fI[�Ոϔ�{����jX>f����|�݅fu��W��N�:񕖂��w���PNF�'��7�z��Gߗ��Jغ�G*�:���`�r��yg�����
m����[�(L�~}e�tE�B|2-+Rl�a��=�C�W4Y������Q�˂�Z��v����ߥ��ف��&+8�N�7tj�G�<bx�W8*l؄���01x%�8Nˈ!�K���F�kq�Q��3���-���L�@{+	/.n5e�fG��2� N�����c*Ԡ�o![�/
���|?���k−���&QL��q�_�&!u������. V����	�3�� �
���]�0�t5toD�"��]i�S�����1*�ѽ[h�U�+�����/�Lw��x��
˶tу	|�'ȿ"D@�&A h�T��Z�������n���c ��L�R�ޥa�uل����L)Κ�c�=l�ة>�ڟˌq��ra�ꯑ���*�Y4ry��wT��{[|T�&�5O��q���I�<�h�W@��j����Җ�*�	��>T�7^V*;��?@X+�%�����g���l3�w���tl}�~�@��F��#�+b��{��鶀��mA�A`�(��}���ŢsYp6ҕ.�^�-c�X������}�'`�����TZނso�����S)��t�I��c�\�A�}K�ϯ�u�t��?�^��s��r�f�`����AH"/@nL�y �EU�b��>����lN�h���Ա?��^�n��Ҕ0��5)*�}��d�'����"���?]T��?&Cd��#B��G
0�h�8%�����!���y/5�i�kp%k�t3y�d6�g�l�Y�$������Z��P$ E���G�B(��#���l�Ll@�rݰ��Lb�LE����8�T'�N:w� k�!�z��F)�'I�EI�E�K�m~��\��">,m�����?c��<����#LΧb�@�ey��q4U`4��[}�r`�z-dJG�1	fZ����m[�5{���e2&���Hc̸�DdB'�Ys�U�G�����{"_��&�F����%Q}"��������U�/�rL���Կ~����m�5���MU��r�=��X^��Q�h8Z;U��6i�Z3R;��,�7	�)�	4R��%�S��y���Ǹ?��Fg՘��[�������� ��h�.��_Յ��V:'!��`�;̆r�T+R2Pʛ����~�vXh#=틞�I޴0[����0�ġ��N�s�Xv�傔9mY�]3qL"_	�����~˛��H�=��<��H��e�J�E��R
E#e*�.t�B��o��e�W}z$�� �
w*��G���.]��	4;s{v�<t�}��P �8��PXn4db�EA�����Ҕ��$��k��7��\�8?(�$���ͧ=���qF�H���W(j���A����np%�3�$jS)�Yǔ�Sq5f�Z�I���˽o\�>���3h*h��O�1gb�{G{��[�L�B��J���&������Ԥ��`�\�$�+!��qj>�鱚׺J��ؖ��ދz	.�'cd��he� J�˰D��j�&1OJ�I(�vz�]���hs�fs������FP�n��'.�8���a+�e:O�'H�qP��'Co��9>4����}7g1G�����d���	�홑�@�T��U>%V(�ԁ,i}\���0Xn�h¦�z�s2$aNG���H��D]<����|{��z�ݨ{m-MS8�Q����Hy��f�,��:��0۠#��l6�����?R~��N��l��]!&��������j�șe���K����Qb��L豋�_t��&���?�Hg���#�~�l�J��$F��k�c�Ȋ螀V�!�Z�~�ՒJ��3W6��)mJ
 q?!L��Y��>ƔTv14d�>�
wx�4�>{��s_ ��¦��+�
��%��τ�L���\�Ω)vn������������
�,$K��_�*g�����qH�r�*�{s̐��MaE�!�A\�������4�[�l�d����s�^ �N'
0U�=ւ�0���J��t!����;	p�%�W]�F�?��`��ۅژ���x��!��|ՆCJA���TN��ly�ݡj�ϾnI��"��T����c���j�C�)	e�M���ϩ��`M��(�����|�Œ�NQ�VW�'0d><��������%��_� I�
���V�,�l�di24��'ů���9���g��CK�uA��R�V���E	�����.����r��7:qh��B2)��-�Q �k����[m������CF�	�G'�2��A�c}�ͮ���+� n�6����=
��R/�"#�����)��z��<��f~��l10.&z.��I7%]t@���Q�Սkrgf�83D{��Em��e�͸u��WT������ڪ�*�d�C����L#:�wV[�	���(hB5��lC2��v{��=��to�uۍ%.���Tں�S~xv�C���q�y�m�V�{�sf��Yc�F�Xd���`����ըAU��~fG�i3�gZ_��R�ڲ$>��)�BH6O�����	I�"���(�B^�4����֧i��_NSQ�q��BrΔ�Vk;�1�Q�]q�]H��f�a�,�������(�=#��C�����S�	��1miE&��Pby�A+v�AA�G>����Hg�	Ty�LB�8�3s��[!W�r���fb�I�,ȴ�r�0(�A�72�wQd��.��:.�%
E�"8��U*.����L,L�zA�+��*�y��J*E��z���qM{�&���4�¤���ZO^�:v��y�Ќ m[����;�����H,0ޓH�;줄�R4m/���:qr @�z�`a���g��+��[���A\���<��]�#z<}�#� 
�#���/n�՚lh&L���4�L�W_�jg����7���]�1���$�S1FM�o�Kv�`��E4��n�mi)��gc�I�)Hs��X��piV�b��y����^y׋�y�L/�X��qy�|�@�D���>8�n�E�Tڲ����F .��y��Z�ų����]��g��3o�j�hn�p�!�b�'�:�;���r���'83(��m�F|��%B�b(C��؊�y����
=��^q��-=0��4�G�{UnU{CNvaJ%�i:�KJ��ݷ�����R�`v-Pb2z@�ꟶ��ֹ�5Δ�^j:��hh�C�@I�=D��^��������mI��Fo� p��{���Q׊�M�1lI��y8A}ֲ�"r�Լ������.�N5>��p�0���;Vk��@v^R^�&�9� �!_J\ɱ$+g��q����	�_���7����F�}E����XxP9�OY��5mF1]M�bQ�we'�Sk�+LA���:ơ��9�����5�m��']�J
��O�{��ԯz��>��IøA|�<�y#p��	H�#�%ݙ2�s�=r�nmB}��R�<��}�0x��A(K\W��<�4�(�8��oa~پ���.��~O��sp8<#��ڏ�t�!�WCs�W��O&�9tr�67�D-��M5zz��@��\E�����E���KM~����_9n5��E=?�����l�.E,o�Ɗ[U�d���u�mn�C�*��+ K1K���=��(E̊��%h0QL{��}��1i6�L�}���~Q�$�ɓ�ݮa��r��!�+cD�K|p)������CW��א:8U�Z�Ϻ��R��Z����T���F����'-J�˨��CS���8b�\��e����`'u���R�$�,���\sу���i�o� b��c�Tt/n�vr���E3b���.��������{�?��ĳ��&�Ǭ��`�����2C�/��u�]��Eq~�#aj`�C�l9�>������vt�2L� #vh���8���������}`���e��w�jCky�uy���jq]r�ی6��q������D�=樛��˅�8��yC�aķ����y��v��.K^�q�?�I�;7h(�}_�ן�Y��$�~��n��k�ʏ5ǻ�*4�jE`t��}�R��<s���-�,3���UB�(G���	|�������-��e�z��!N��Ef���nL>>���C1����D��"��iH�J�^��T�I���U������~��Kp��V!���G�,Ĺt�N;�9�l�۷���M�)۫v�"M�)�X���\�fcb�.pt����/Ӊ����cf��~7 J�T���48��]io�od��ޔ�1;�n$��1u/3��mu�+<|#��?��氀`�T�+�n��2P��!o��.	�]Z ������4�}�_q�L{��G|
���~P@ D?Ib?p)C��<�h�5Cx��tC��2� 0}h�h⢻_s[N�x�ˍE {�9b��bɧ]R��H���C��/^��D� [�7+��������*���U�t��L�M8؞�0S��?��٥IP�	�k>��%��/�"��[����Ѵ1�Ԣa@
(1q:��r�q�y�u��d+�׍fPl��Jk�nX;G���E�}~��ӯҤ��+y�DB%VQy���h���p�:�
�d�RzFζ���/�`��^�y\�M-��+u��Q�eF_��Zޗ'*Є0�s�5��/��m�d/]=i"(���?�	ġ�oЀ�_f�59���5/�������m^��_����ծ�s��	�0��e�[��9�1��u`ڮ<�`U�d�����@"WR�ͱK?��������F�S�M��_� ��m*�"a���a�:Y�X}��:"�ϊ�F���%�⮁+A%C�R�=�!�����["L�(!�zM�v�0P��̿'�_-��^Sj���qo��}��`��x��ak�������)=qЧ��e���E�L�i�Q�F�{;��Fޥ�����V/����j�m��ll�G˝�=�e�6�+&��W�66���u�X���Ŗ�V���v�{k��g+���l��P�����T�A�����k�N�D�6%�����W�|LhDo,��&����'"���t�7m�p�av�!�Q�)��X��\9�y��"8�x��Y���},��9��>w�2�pĵ̀vp͌Α|��2�}*�1��y̑~I7C7~��td��RmV25�A�@��NnW��'��Æz+�ZوK�y��a���F�!~A�py͆]�2�%֑����TU�p�d�v5�ڽ���/���bF��<E�Ҧ���G,J�o��ܼ�e����0�kU䳶�97I�@�<��J�A�ٞ�K�}�3;�+ORH/���'���	냈��P��Roeж�0�������v,�������De��[�L�|������+�	�gf�����'�ԗJ�?G3n�b~�-��7��Λ 0��[T�7ɾΝ�T�~�_G,�f�ا=k��`�ydd<�׬\�'s]�������jM��U�5719/�� �J�O�G��,������ó�Whr����A�wf�����#ٟ�Y9ڠ���"��5��1�J� p\w ��'�sc�K��,D�U*����!�ͥ��R ��ͬ_@�D:��E�E;����GsEǨu��eƨƔ��`���֬�`�w���߯���k9:�D�F	J|��ӹ����5􀅨D�є6�ֿc*����Q��=����ߎ�w̺r���P��xg7�٤�h9���b�C�z�a��u�0E�"o��` N�+A;�̫{.<JM]���'�Z�!�d�g������D�nE���M��^��P36����Z�_�!%d;-4��n$��j�� 	ʄ=&�/��L�t5���%��t�i[�Tۗ��<S���5v���W��}�@J%�"�x�	ڍ3X�#�w�J3�ݹ��Urf���7n���{��1�ۚ�gj���_˚�(Z��T�F�9;�*�F��\9t��iP�`��'��U"�����:�e;!K�� ���[LI��ä),|v�J�U�wq�5� ���� 	I�-&�v �t��y�'���N X!WL�Pv	$�4�U�T��D�����L�j���k˘c���4�����XW{��4�ޣeq��$�z��{��R�^j�O:�d� ��3>���q�����}��L���1��vz)��=���K��b6(L(P�Ⱥ�����iՉ��͗�-�w������J�&e-��U�����B���� ���t�:b��DV^j��f�n�Q�FQ�'D�2�Vq�[��*�t���4���Z�a]�(�������#w����M�:A�����ɬ@���G(k]h�0d.�xIL����Y� ��K�>6�?/��w(���i0�fx��W:2_�ӫ9���i?&��wh��T��_�v�/��z�Y���&\(!U}��R)��Ϳ���BzB�/��� �Qm2=�7.�����n���CX}S/ �}��xx`�_D���`A �.Zd.�.EhM����M����cd[���0?+eG�'Pha�4�,���q�6���b��ӕ^0E�-w�����,�7���p�Fr���kh��r1�l�-�je:6k;�;491K?�\��=��[��P��&[�b�"Lж�;l����V��	E�a�����e
Ir(��3V�BbzC?Me��n�+$.޹�^<��&�f>�q+�ߥʡs�-j������&>5�M���� ��Q�`�/Վ��u2F!p�c/��C���$Ih3t�s@ʟ�'|em�lPN����ʢ�6#I����T~����mn@m3��+#�˨U�_=;K�Ȏۘ�>���Ҋ���¡�U��UM�����U�Ba����+��'.�Pq�O��'�M?�2J\�d�n� ��(��O�J������x.dh�z���C�>(�A�bF�Ϥ��鎙�[�q��-�6/�4���W�����>���X��I0`nW�VH�>�G�@�f� ��}ݯ
Q[�g|�>@��	9��b_>��]N~�;������ԗk�|�������F���bJ(���5/�8�WP�כY�>�>䅅~��i�+�{@����7�^\̸� p�����`���o��xUW���Xk$}�wg��Rn]0S1�p8!�)�p����jʃ<�M��
 Ғ` M�O߸���g3d�{�ǝ~�n�pw�7���[Y�K��g���lj{��h�����_r��#���❋��Ծ3�ܧ�pn�b�5iL`�����ȁ2u������v��매�Q�c�´q��v��6�ͳ���"�%�u�W�Fa��G6m=�����O�%���e��x����o�ܸwİB�.`���7�������}z�1��X�(_���#J�/RL1�e!I^Uу�_g߆��\B c���h��/ϫ���6h�!�	v��5M����{G�R�z���C��-���7qʘ��0R���V���O+��Iz����w_��%]qN7��RӒ�eRO��?dڲ�^�t�h��B9����ZAhXܺ(q_�՜R�jW�cq�������c����V����ҳ/�9�w(c�!��ܬ9��m��*�x�0��wdd�=��߽X��6��:wd�h��5w�����ɒ7��-����|k�Ğ�7�a�yJ�f�g���^��G����8��fv���5U�Y���CzC~�kO`�N�2��Xb4�[\B�c�L���|��c���n�vH���l]�՟CkN1r�f�[]�5��7�T��Z���Z��{�V%�jI�T�d�,u�k��}��d˝e^����qȴ5���n��*K{����׉�H$	�F{6J�+	�'�{7P���O���,)��%�I@y��j�J�9���i�P��kp�,���o���@��7���n�6!����X�F�c��e���Pe��]�<g�#ЪN���%��i�90R�Z��dӎu�2vV��Q��2�y�]។��d޿��]ك���RFVuֈS{�d��/�|
��l�<~��C^��7=2�������v���Y��=}'��qe�Z�:����������d�����qʬ�ɁZ����sJ�`�2���4�Wf��͸�E���Rؚ`mٛ����à���*���f�8�B���SO��BJ�FM�G������j�T�4C�?�1�T�|�7E0qZ�\1���w�e}/����@���X^v���*�,����d!w;�����`s9�'"H^Xsř��v�l��dP(���.��c�}�>U5�`_/�]���w$��Y��|Oތ���|n�x�>���4���3b*��d�
����>|,�ML{��0�(Sȟm]O��x�t�M���F-�0դ6N���#���?<Oc�"
�Sh�EGg��AM�A�o���_�j�q
so�7J���A�ۆ��63>�z#�y�	ƘX@䂐��EI���it1<����~6R��?�A�y���l/�qa~��'9V��N�RD�!�~�yʤL(�t����2�W'��1N��ϙy�;-��QB�x.�ǺIқ���m4�D�$N��%Kj�=:8��?aY���2��$/0����<��.�6�u-b]���\�B�fts��d�x�&۹�I�����4d��ᑈ��y]~�*fӋrS`�^sm�"a�+�\�lu����
ju��`�m�P���|3P��3�U���)�\���BS������R�h�N�;�P�d{�[�m��=U�K�Y��\�����M���M��ʝ	��|�Fd�PgK�� ���������=�hASTC��HS�3�3J��F?#�4 �@sĜ�uQjHB��d��HTa�&@-@��Q��$��r���Y`���3�jy�R���U>�"��/��*p$���։�w�$y@&<d'��
?�� ��;��B�_#��ёQv�����E�<�=G�`}��c��
�ݡS�MզYöɶ�6-���e�HKD��rm%�Hمbk`�3�r�[�6�ID�������n��o�8�.d��q��[���ID��V,vd� =
��~������~s����о��U�Tf��eqA<ӻ�B�րx8��jԞ��ʰ����T���� :2[X�;g��{H�w[����w=l\�d������I�M�O�Pz�5�G(y���Q��w)�шt���B���f[��[��G���"��2���b���e�f�9ݎ��
%e5)<���t��6h�6;�r�R���k%�������R�����H�����H�x�wƃ�!�hc�D�"���~*���j�����>*4����/����#JS�1��&��.b��E8e���8�����02��s� [����Bx�q����? ��	��������z��t7z���j �.�����ҳ���78����۴����7�IZ����p�_RX��ێ�(�Q
m����h���*b�d���K���7Q?]�8��5����f����� ��q�N|-�zx\- *߂5�e��'��8�z}��9��9'��;�?����P㎚ʪM)l�5����k��t�~~���4�����Q���q���Z~�M��s��O�8+6b_�0�B�8ĭ�r�Μ���,��-Wd^{�]�Kȧ��ǘRͣ�!�8ߐձ]1�ҾB=U%�]�V��}>�9�.#C��ԆX���ɪZX��R�^_���<T,�߱e�h�]��M��t�B5dc��o�*"!�~n���UzV�d0�<K*���l�t��PQf�\������T����ܔ-˔��91�.����&VX�leG���aB�4{���d(��\��E^��|1Il@����	^_Đ��n���h�)��l�W��W�й)���2f�u�`�}R����B�YA�-݋o��ݒt>��#�0,	<K�.�҃�Q5ʷ���{�̇Uҫ�y�F�0%��D*9}�fq�3-��u�2c �;���~�{����41$�dgh�3��e�f�1�DJ����:�뽋t�$w��8�L�{V������7� ��:~�s;�1��Mí��Z�{$��3�!��Kg��?�YQ��x��{IKQݍu��C���H6PD�ӵ���ʪ��g¯�`.A~�3��� ��FL?;4���z_��i��/�NW���l[έT5}O�S�P��
s�D�T�$hͲts �l�w��̍����1����D�Wp���I6�,u��&��5A����Z�=�+N�ќ�[C+9��b��4Gx�_���:b>�:s��	��0�5I^�tB����C�8�"M��-ϝE�u.\\\:�;��M�>j7]T��������م�u���`��u,������ �;��p��@����P�ꚃ>.�G����6k�sp#�RFb����#_���O����U���~p蹵�Pi:5.Yv'v.��H(2���|��.��z~CX�Z���:�U��Y�[�d�Hy�v����i���2T-c��h�wNF����ө6+��nu��TZ��B�����=�x#���am</�6��� O�c��}O�H�OO�G�C�j�h�*������>�V��D������mآ����3��e��	)�_J�
JW2=p�K�W-�>�Ȕ��3�*����@A%�j��h�z�Z�>�i�@�3�����O�"ȨPi�O,�X�,JڤKЁ��	��E��(y�L�PN,#��[��k���z=
�	|�8E���ɒ�O��ܞO>g"�m3[�0C� 4q�3�	�t���_������t���KIb�-����� ���秱z�g�
�O��[u<un�^�ݧ"��?j��y3��@J�Q�V�g4������&�
�,��6������\�]�粿� ����F;B�p�k}���ҎK�_)���=�2��O�OF�Ba�GF�J߆<G��F���J!q�!��<Ů����5�����֨K� u��骀n��\����p������>�<F{p"�������������L�rxj��x��NQ	A�����n	�g���X�M�Sca󺹵u�3|�>��K˱��-�'Fs4IB���5���9�kD���+���f��Z�L]���y�\���8���%���&ح�}CxJ�2��6���	!+e���'8&��VJ<ެx��x���p8ßI����,���mI"{g��O;q�ϔ��GG;!L-���ྰ���'���D��ف��r��[��,�V�fa7��l�n?sz�WJP���&hRVf�lE%��o�g1�BXǿ4xҨ6�x�tE��}��{� ��S�Y��9�.w(��ڴ����1��Q�Դ˰e���[�a�^�Xp7OI�*�=���!{���5�.#���k�7���gf9ÿDXES~�<��������\�[y'U{��	�ڝ˸�)m�bN�F��<�y-�|m�;���ة�y��.m�s8��%�]�%����M5rk �`�\�m�*h�k]�.�~��+̤&ه���2`��L��h�����������kʱ�v���Z^�"��(���⳾b`�G��������d��̬g�
R��'��؝�_T����� ��j|-/��9��+O����#y��Mh�f�&0�hP��Ǳ���?�7������I��Ŝk,�i�3��1�g
�oPfG�h�X�ۋ�|r�C������T5%�F���kj6�\r����	E�ΎS!��%�-���oߞ�_��B�s��r��ߜ8��S�Ӧ�-Jts~�Z�zi�Es Ć��=W��O�׶�0T�ۻZs��w���zaVx:	/�k<��(m��!X��%@�r6��rkO�=�g�\���X�D^K�abl�	Ϳ�)3��K�n�ٳt�шw�e|�k�c	�D�0��*[i���~A�.��q�5o��/�	/$'�˧�)�9<�qk�ݵ����K�!���a���P�t)� Z��Th���XQ�dh��®]R��o
�ь�ؾ��"W[հZ+[�L��]�dXe�N�����x�
@?Uo���I��4�5�&<3��t8cV'��i���]@ٮ}��=7�l��O�_ SY��>>���ó_�ۉ�wll�rx	������3Hk�t�)�>@�nG��������۵&��*
��Y��h��P�g�PP^���;����5��Uv] ߥNi~���i��*�>nat�Ͱa���K6���\j�鋆c�%:|3����'~\K G�,��//O��]s�KN�L�pi[��7����g�N@�,�(���1���^�$Ռ�ǥ�CZDN4��2K#�:h=�o�,�5'��3�O�a�_R� ����c}[!C�(w��F���j�9غB^GN��{�� �"���=L�AcJ���[����~M�rA��e���������7�o�o[�cd!�����#"Ӈ�Sq���H
f3C(�g�j��k���${(�)@W�A�*���P�G��I㳡'ڿ�"�ʼ�x�2ۍ��ue�y�r����<��ߵF��0:��6P<d�:̪}��D$7��Uj�"���F��tg�(�b+{g�~�"�p�kY�(5���o��ȯ�sU�!�IQ�W�
*AzIh���mH��G������R�����WҡI�U_���%��XW�Dط�Q�F8ý�XÂ	D:��! G�v-M�6�B:7���R�voz���>�`@�5�f�#�^=`0n�0��y)�|���N�U�+ ,�H�D�51')�[ rU���[4/��N��TE,��5h��k�Q��M�L�A��y`UiZ�S���7�F~���i�}��W��4f�0гA�d��ki�y��:�5�������a��A!�)�J�<���Мl7�D��ȼg����Ց�_%~��V"�dh��?s�0�X�>�[�r���>u��0Ԫ�珇���_��K�:�� ��W����[�d����X��C��%G]���rs���n��_�O�0�#X ����K޶ K��19B�x�����U�u��"�S��_9�c;�B��*sQW���ũ�Z. ���o�Ƙ ��N<[e-U؟�KTH��N��5vr��gK��w��䨞���.v�w�McB���}��bɱ/���9 \iײ�>�G�P�%��yl�_^�+<��D����F�aۃ
����jS6m	+	��֞_$gy��:�-T��RfN%^8fM��^�[ܔ
�V~N���y�Ԛb��Ǧ�~g��̇�t�����33����i��g7H8o&�l��%}�(���챢y|��#�H�!\��-�����:	��p��S5�GL�����\s����W��7�=�G4�@>o`������匯��u�sU�q�|LeFK������J�ó�>P>l���q�-�/T��ddDnz�.Q;�hV=1?�X���(A��v"U�BtR�Ȋ)�cƤ�\mY�t�>"~��O�
���U����Le8��#���:,p4w�|�w���{0(���Oڜc���5��q���g��eU���SЪ�X 4"ZU�
��*vl3��xI}�t�Ȱ�ېT��CF�u��RD\ӄ���Vu��V��g�!���Fv Y��D{Z6a�$C4R2:ۊ��!�~���IFD�E9u�tQ���0�%Y�അ2 �(��9ʾ�ݣ�G�PF�bʏ�z��3@��k���8p�^o}���K]*���2��sMs�G�.��O�'�����_P�]T�.��9��������[�c �\��z�#K�[��w�O��{s�^T҆A��2~�F>������x0@"�J����Rڐҡ�w۪���,Y�m-�H�Ԝ�[�I�u����׋�Ԃ���)Ã������\�E)+������k�g�9���6���c��j���x���[m����5�K6��\A����H���S�+v#
wt�MN���*_��~�
F��O� ���Z��G=��$sT�m9����v&h����=l�M](���cH=����IH?.݁���<+���֎������ɗ=sB�c_��I��į1t�+?�\�,PņӀ5G�E�*��Zu��t���=s�+N)�j��-��_��x�@�$���GMT~�j3o��<�-գ�{��N�w�#X��!�8���&�-w���bJ�ƙJ-�:�&
�i
ay��dz��w[B�Q&ݽ���z(�Cj&h�S2ʔ.���k�}4WYs囤�Y�˱ �`�	{�.�6�idF1�,w��T�q�3]������k�
�=��D����U3���@Z�"�˔Tt�Qү{s\�����96��&3�UBgiʸ�K�?�{MgB҂�����M�蹧�����n��iI�-���%�{�=�\��6�z<�v�����h���ZgН��ReF���f����JŇ����|�)[Ɋ�h�^r�ߛL;�'	)=!��c+�08�����R� �dB�e��? 6 �+�D͗�?��$A$�q�N�J�_����0W���=� �b|/��Y����Z�՚��F������{e�򍓕r����.ӆ���Cȫ�6�}��F���im���d*~����	��	'���k����#��m�^D�N����2�K&�I��dp*Kŗ����� {��[�Ldu�x����Lغ
���]�%zR�,̟�3
-����v��Gɮ�����
g���ؚ5�j�	���1p���Ļ�r_4Sڇ\9;��FS&0�'cW���9�K����[J�k���ٗ�O	G�P��� ��PFs����?F]�Ě ��;��*|�D��h�r;n�n�#e:g�#���
2�`!&<d>>֭0�����FR�����>�32O�W/�R_���&7�sYd|P+DWLϘLI�´ne�M��E��6X/'M���@�*ZUp
$2����O?����j[�R�o@���5�
&i�rp�0�a�=����o"��>4˹����1���h/�%D5���������5wPix�Q�@m<���T�Q4.���W=�$FQ5Y�����BR���#�*��f}θ<d�q�qZ)\���z'�����`��R+&ǽ�:�=� ��o��z��F�8|%���ϩHT+����NA:��(L�DA:'3�z��t�j7F�؄b�������C��l(����6�Ր�XS�N!�8<�0H��Ŋg'z�-��$)����tLe�����g��������Z�(z��qS���@[�"c�,g��S:��J|�wOH�A��W�ɋ�ъ�}��v����9��^�Z*�d'8^r?=�#��o�R�!�2�� �˕�Վ�o�9%��;_�d](���娯�=���As�p�Ψ�4D����S"��]>�)�F6C�[&;	�"��rnkd,�6�ӄQ�AE��%Aʹ��������ajo�)]d E��!��,[o���MI�L[i}K���N���y����+i����8��Y�P��ä#n�:�/���P��r�LjqqW͚F��6 ^���6L���&i*C��<�uQ���� �g+�P�ϓ��	�˵�(��qMw%ip�{=Ԓ
C� N��JԪr�����h��	�NT��JF-�{��@"��X����ti�r�����M��~ӱ	1�(�]�Ȫ��w��,VǙ�)>�|�d�f��e,�	��DN#����۬��IlMi��Ŧ{�ڧ���W�<]FB��㣍��M��M\�9 �V]�8��L�XBZm���'�=��Z���"%3�Z����M�i��
�u��hf>�Lص£8%Տ/ �8?�s�bs2�`*B�&�����1Ŕ�I�??Q�1{�K�$*�������[�+�Ϙn��b�c�C���IJ�Ῡ`���3���'u�7�̓?P���_�+
�N鱺��Z�f���P����*@ɡ��'n�L
��Ȑ'�N;�yx��=�Ǯv����a��E�BЁ��R�_G� n^V����7���@
ɚ�I�(?�qQiQ&��`���Q�I��zM�7��k�s�J@/��N %b
<�^
��]��R�S��;�Rs�E���b��*mAb����R�u��`$$�w�6��n��o �<?�0�GM�i�3�;��J��ʆC��=LN���S�y��>��{Q�Xl���K�,d9�ȋ�~$���[�����a-A�nl��v���L�N9����ԟu��.�mz���}�UA�55ښ
ߝ�BF�x��/�Ad���:=F�����m�<��(u��Ϝ�Z��?jbL*�51�? �W.(��I(-<�Q-��]�w������p�	y�khk�7��mQq��n�'<ڍ�Y�Tqf$�R�ޫ�����
�c�v�.Щ�
��������bN���@����JD��$w�*D>��<�ؑ��H�"?�{�.�fO��C��P��0LGV4��E2�v�>槙�~��|vL,-Sj�9URS�7��n�Fd�q	E��	?�� �3���a�-%�5%�Cgs�����.B�@��
5�ݭ㥆�=�[�m��F���{u��DXfJ��EڬʚW��/���G~hx�`a;����dv���T�⺎Z��A�L�v�Viy���P��OrZ/�
x�Q>&䃃���5����Gp d33�i�
����s�D�H�b�ws�<h3<��1����S��P�퍡���|7�-�7g G�&]��Gz����/�:(_���2h�W\g$�S�{0T���Psl��*�|%����E�;�����;|e���a%$x�,����j�==���y@��v�cD�ޯ"?���=~k[�1� �n{�j
��f�C�>xq	�|k��y��}B��a[)xؘ{�ѐ3PA�n��D(��Dc�k���9����+��/�Og��	�P7S��cLу���<��K��U�O�S�֒��:e:�ؤ�ӫY�Ҽ�J���==9��2���D�H
v`�"��x	�O&҇~݆��jg/jθq>tt$S�D���� ��>�]O���z��r��8�"o9$�3���0�݈;�7Bm� ��Ԙ�c�G�ϰX�,�d{O��NQ5 �)�p'H�J�bJ�N�2����Ç-}
qĴK������4iI�&�:�Mkȗ���5j�����D�s���L/wU�e��:?�R�bHe�f�X?x�f_��!r6�hq˴�s��`^����(�W�C�Mtx��b���׵w��r�
�4����+�wh@��p�V�*t:B���b����p�'�7��u#:k>;D�'�Qg�O����5��5���{�My��G.�Z��y���K���ћ�lh)���Ż9"��0����O&��__��	�B��ol?������E���B�����>�G[����IH�o~�}��$F6���v���l��X������vR��XNx��4C��K ǌ����$k.6!^|6����6vN��<���X���h���+��/���*
��X���ǰǌU\�D́ɑ���&N!ӎIeI�O|*C�N�^��z�&�XC,��g�Û����N�b�Dܿ�'�T���Pߩ���T\WNצ�K�o�cHD�ccL��JɅ���i:`�Hr�]�4A�#x��x����dE,�w�l�7�~���-��&�V<����K���n;��m��`��Z8z�xbo��h�/ƇD}�s0ж��ִ�4r�!Hb�C���
��֎��iv׎^�Ƌ�T���2��p�����i���S> RYՔ�ؔH7ꪉ��ֲ2#�Lh\��Wr`�\�y��j"YX� _���V�r��O7?� ���˥w��B�����#n�P����������d'&�2� �1�I�R C�[���z�Z�"@��;Oʄ:��=$��:VA�PGe��Q֣>���&<Q0lO�R�y��1v	�04ٮ�2PDh/����ZY)R�aw�{f�N8ח]ِ��7�V��!t!F�I�b\n���=���ũ���3�[��|��K�6=�X��2'� �ܝ�ѓ" Ő�H�V`�;Aӊ�܃��xdx"�}�3k���DM������\B����A�ϯEP�����i�8�0��Te@ ��:8a)s���?Qm�{�\����5׭��lnN�v�I��s�Lp+�e�]��mT�\j6pK���0�����'����b���/p
�̕�&"��z�C�%Ţ}������F��O�#�e�<�Ƴ�,�A"�:�s��+o�/w�'P#�I�v��z@p��Xw���?�L��݆x��)嘀(M*�+��W�Y�����J��9LҰ��i0�y�ɣ$-/�m�Q�ض�nO�ɐG�)��P@;�4Y|���k�����->��tc%�k��K����$�D+�15�sw�]!%A�;=z�K���r̔N��@0gq��N������
�'��&D��I:���{>gw���-B� %紖L�H*�������������Ԓ��[C5�ԟ��t/I�'w������$�9А�ɷ:�K��v�@t����T�vç폛�i�����\_ct'�~�6�i� ��u������g��4m�Q�cŲYBڕ�F�Fb��J��@���;�G�b9i���H��_�-��t�e[��̡P��b���N�VT|�ԛ�(v�%lKb�m\V@�G!"Exu��pw��r��-U@f3����)�!汢{�Z��:u�S�l��}����J 䑢B��cz6�_�x��wǤ7��&A�*v�����_Q<J���i�r�**].��n�N�q��Չb ri�X�hMřCЛ�H�4��+����v�&����,�V����q�!�{�~s�oW�߽�m��Ƹ9A��B�@����T`�7w<	}����?鑍��~W�A�BZ
��w��7��aBV��`5��vU�M4¼�i>���+���n+�P)7�C��AT<K�~A�J#������Cn�}Z�0t#$��#��	���4�.%Q�v���\��{��{��D������p>��L��~��_��oa��8?&mEt`5_<S�MU�hT�.�|ϫ��/�j�����_�3G)H�Q�}�Vi"�T[ʩ9:V4�n�^��ǁUZ�:������r���LEpd�<o�����&V�O�M�8j+jQG����`�8^l�'î�+��IlA�Z�W��ʝ}2�u����8�����K_|�I�V�20y�'IS \AR��^��lb)~|������������.�h`�+�<�|��3�cPsu����L����`
�g9y�pY-j� ��!�,���V�C@���]�d5;'e	��z�������QZ�,����7��39�)��+L�Q���J8b؈ ?��r��K�x��?7p]M^B5��r���jR]ʫ���zt�5�w�W����QV��.W�ᔕ�i�^NP"ɭ�w��:a[�|�)g��5�?u�3@R[��7��^���{5����pw��Bz���j��tX��݋d��&1["06�Պ�ߧ���qSA>
QNZ�*N7u�����*�O�]� +����� ;6>Y�uuP�9���r��R��w�h�Nב:�a�Ā uM�m������1���v<�4h���vA,���beFF��{���V6Efe����R}�����Ow��	�G5���Z"���\�u��ol�F����Y���)m�h�V���OY�^��\d�AJ�q��2<��g�0��ro'#² %��0*gu_� ���a����%��h�3�b��ٝh�,����C²Շ(�j����~O>Ш"�[o. "l�q)"���#�	D8�]�~y�1m{a8��tX��By��3%���k����� ��&���N�a�kt�%M�:�Dv�mtP��й#î �r�7]aI�JդW��$�;ȶI�ؒ��2��A�؝"���E*y��[^���
�tA�W퍦 [�k1|Y�_8wJ���[I�wJ,����>2�2V��N	����QM��(Ȥ�L7�y�.��K���<�?
��f`9`$�w���MW`���bm�+6�JV�DB��d[bX�o�W!����iW��O�za�%�ǡ���&|I����2��cj2g��l���*�إd�jҹ�F���T��L�ooQjmsԩN�~�)q�~���>�����<*�z���DP,�LYO��o��מ��;l�h�飔��V*�.�o�>�i�P�/8�7�����|��g�?#�������y���ȯ_Z!��3�����q�&j��'�[T�Ϭ�����Aۢ����!IfҼ���u>�iV'kRWZJZ@rP�ٖ�2��#�;�g1šl;:���F������A�_�����Hh�f��@��[н2	b�b�p�-���`g�C�����+������i�n�f��������ʉINl� �UA���v���e��4�H�b��*�����2̯?W��s�)X\��ꦱ�]>�ayz	�a��D�n�S�1�d���f�H��6<F�!R��28j�}h�����O�Rj[s�̜�rΦQ�5|}�H���N�����j��J4!$�4q��U���0�.���*%�2>��a����4�:e"�b�c�O�7�K��v���c�G�����?�t�P,�K��@��C<�mtIб��=��f.�]��O-di�Q�c�_(Gtσ���K����Ae"���8�M4Me���������o8����m���&���H�Q���uB����e�$��E��[���J����&`�C�)���ު�z����1�X����ӡ���<��p���,��ɞ�;�7�`v!q����nuZ�5tғ�͛�`�Q�1�3���=kv!�Q�1�� �?�d��pE�V�t�ִ���.��v0�ѣ�<��D1t0��3�v;���|1�O�����&���Vz��
�&��ƕ)�tYnԇr�~�TzΡA�Ųw��E��Z�(��XR(�i�����ݧa1�΅�6I�ae��f�f8{e�؇)_+Wu�:��*��
���B��ɿ^���	q���	�7N~0Z��^�#�S��ئ��A��ew�gn��G�ȱ]���,������'ډ�}?S��.��T�L)�=��=C,��dc�~w;t󷾌� wb|�&���B�%{�G��H}�'V���U�����c�ʺ*�8�k+"�p���<|<��<_�7�x�L�	%k����Z[ �g}�DV0�3*E��߼�,�{��"��'�����=����b��eF�/�\��.�^�?�ş7T:�0�@�vD��wbU�D����k�c~]�M��?�Ӕ17�SD.1��r��T�	��H`�tYa�
���@��.����i��#��\'��Q?-�h�x���@,{��C���x�Z�����u�v���� 5�.���.��%yZLP,c�ʁiH�yD��m�y����='���r>U�q{\T��I���)���=�L��q���XQm׀KY��N�Zĩ(S�t`�f�����E,31]->��-�[��� �Irń��e�@���׀К��-������~�e�_#�;�έ��_-�!k�6���y��xښ�k���+@�$� ��/���RK|hmaodժ)�!���N�}�C�0�:�&��
>Q�e*�8���<�ѩ�X�V<Z\�
ټBd��L�X�����o��Q��uc!Q�h3}\Z׫��Lr�^�w[�J��}^I�@���6>�r7P���F9yx6�5/3�k�Fў�W���]R/R�z�K��ww+T���7�˘0�����(�7$�mW���bcncWh�C� �e
��/*��f0dM3rD~���k������4�֟�}R��;�f���V�*��.�L���@��w�YȘWf��Q@OdS�\�k-N~���3E�}�����G����,Qb�����s$L��?z�$ad�5��H������ȯ\㞇��Xv�EъKl��0a����(��Ŕ���P���Sf��?���,�1y��N"�ز4�kchs��g�oU��׃�����i�\���z���G{�CLbuk��<�vY��ڔ�('��F_mP/�_���쏳������	�Վ���a�.�5�W�ΐ���8��7[$�<r*K��(���2��e|�^úqb�r��|�?%U���/������E���)q��`�ھ=�h2F�����sD��8ӓ7(ܗ%e���̽�!�Sk޿��P���O�T�M�f�{�$������pj$ r�$�dQ���6�h�%}#8�����]�5��ؕ,���`SН�4��Wp��Մ��	��ٝz���T���$��~��K�ju%s�'�)9b.%v��o^��0ۄ�Y �#_�C�r@��_$>�9V󠽔_�s�G����d�d�T��L�ٽ�s�ᅽ�}涛�R�2b��J��
'�l΄&��OH�0�_���ׇK�t4�nZ�@���ؾ����ծ�/λ���|��O���~�em�?�ݏ�򋢥L�V�������峎v�2�q&��
�����)�D�[b��=ցTYP��+܉m��Q~,��o?�$;��=��DF��Cӷ��/�Ko��»N�ȕ� ^�
��bp���U��W����Tas$6.���,���.Q�y3Eĺ�%��ה����JM"�{Y򸈬��O��=��?Y��U�G�@[���d������(��`^)��OÂp���s���7�j&�l�j����tI������*���6)��	����lY0h�<dd�H��D��*Ap
���YB���N����J90��YEr�vBr�!�$��dL9J��V������6:�K0Z���&w~�Xȍ~G�=�)�����6J�r�<�=�T^����e��'�#�o-��w���i���W��F�zD>��?��徬����e�� ~���`��s���K���SX�vm3^��̣�k�#Q�q���Z*`ݥf4t)�g��b:d>τ�w��2�m(�V_�롧��7�c�����g3ۓl��T�b�P���?�=��k�#)of�9U,��T�*t'��m�1`�FX
Y�@l��ӛjKІL�/�Ǭ��]+�m�� 6�b���6�j��#5��A�����H�+�b<3�fsɱ�R�3T�^����=�[��a�����1eH!n�{������؃u�W�����muYX_1p������m�k� �G�?�,���)���_��޺!�h�z9� v�ĥ}X;I����I�>��U��d��.�p��G��⏜���C�z��	�@O2�����,�k���j�2��*�M5n�63�̋�`�kII������̒zU�]�C1����&���0T�7�����Z����=-?�n�����ӝ�e#�K4%+�'!�Op�F�s\�>�+�ot��,'��#n� ���KC|��JRP;"��a��\�i$3���V�o��-�7�U�C-��|��gwk��dH���\��ЛT��P���>ʟ����{�fF%Y��i�ԮgGy��[�������Ѩ��7�Q�[�>DZ��4����)�0d�i�Z�5�l�p������T\�k�P]��B���-5�o��_%�OG��$U�����P�i��� �F8������+E��G�k�㻻����{ڢd&�x3ۂ�Y�jPZbqd$'����c���M��]ܰ���K�0r���7T�-}����e��b`�#��0��L5����r��(�Yt���<t���>�jIs^cF��l�ׅ}����)��-�1��U�;��gU��s�u�17L�ɇ����I��<qj7귦�j�=h!�K����ﱟ�f��h��Gi�-PU��!G�S�P�dM��w�&�%�~`1Ke�����R��|"9���ܬ�pR�#]}ɾ/棁��%�@&�jz�yBk'������1�HJюŸ��j+�b2����0M�����j��T��	�4��I���Y��uo��@{B�l�Bd�ayW���Odv�yq��
&N�U��.�	�C�q3�#�˷�}��փr"'$\Yxe��K�1�ޕ$I�|��B������� ��ߢ�2�F�`	��u�I`T��n/�5-�{\�H 3��Gά�A�O�X�m����e�#���0�^#�z����7�odaU���1:����go�:	�$o����e�ҿ��z]!K~Z����ytD��-@���	��ٛH���^%��B'n�I�_��(*���_�M�߈e��KBĨⴚ�2��v��[�'׮��Fԍ����4p����0Ok�d��'z��[R4ƵO(6{d�)���q�uO����Ck:1z<U��^��w٘Y�S�|mMnA�5O�O�%�(�CD����?`��eg{l��r���wCT��~�� ��}'�\V`�2mJ�wJ��_z�P���"�1�owAä���V�J�d-�b��)� {$"�}&�)Y���������cN,�ȡ�Y�X��e�r\���_�$P�|V.nї�����ۛ��ҏ@|�*��L���s��%x`"Sl軄�	ܼ�������/�%\������=�_@�~��پ��pC��}4�+s8��0 ���{��q$7�j�����\r���xp���ۉ���hpӽ���:�]u�h6ä�}�2��ز8����5J�!�P���M����
8_�z��z�y[�r;���^�L��Q=�	,�Wie�0Aut	�������w2{s�J��g1��=R�^cs�>���Ӗ 2M悛�xl6��7W�6�;�6]�������� ���Yy���s���Ur]P��"6�Z��Lk_�����yn��yӬ�ӵ'�׷�n%#]�ɾ�.���P�u�0���hB)\���v�Kut���e��l@�/� a\j����S`�XͨY��IY�l�$䓻!�}��K(���2'�������R�0��R�5	\���-���9��}���V7��d�j:0ǥ�TP7���aT�3�A�b���߻�% �8�))g���_y/XW���1�"i32o�5{P��O�1kU"�O[�%�� ��'���3$d��	cj�ޠAv.�,�L%�}8Q���vF��B(�����V;^���=�"����u6���"
�?b�8��� t�%\��[s��׸�c-_��#e����.�K�I���6D}�@���AP ��w�b��{<=�h-����\���{��;���Q�1����`;:�2�x��}���n�[�զR!bT	b���Ծ�К�N����2����^'�)�B�@3�����f��!Z��G@N���3v���r��C�R��UJ����
���Y�E��fP���D��:�C���5.� �N�{���D,}�uݰ�,��U򋾽�fV>�~!�?��;�`l̶��E(�sOm(g8�������6R}
F�{`�v3�WDҚ�x��x�+���
 ��<��du8�ϢZ��r�BE
]j�ݝ�˞�M��Z�Hy��z�oz�����8BM��UL�E��8C�(s�����W��)!��@eF�u�Ԋ�P�b�x!?��vUZ�rj<��5�(M�ێQ���τu��*��Eo��8\����K��a9qz"ue]�J�b��Y�#��	�pN�d����3�*�_I�d]�����݂l�&4���]��S��Pݞ�V�z(a�����ۨj�yɤg�Ȇ�=�ERMdv��+a���,�d�?�#��3A��>���"T�N�g&���o�E��H�_�C�I��9�J�H�2q���ո���)o���o�%����˯0#ۡ©���$zC��p��>`����􉍙�d�&�>�`���bg�K�/%.����,q���$�����X�K�Y��sЫ)�<)Wk$&�������/����v���Q+z(�pW��>^�կF)��tB����E��F>�g��D��{:���Cp�](11�w�AG�)��[�a�R�̞�y���y�l����KV�RU�[6���d��1����,p XY�1�D�&�'P*?rHGR�(H@u��^$5�������V����76yd�G+s�4i�Tqv��'����J�a�pr�yVi	$:�o@�/�(&j�Cq	�wM�p/փ)iS�=��{���?��Vʂ.���'6����+m����q�T����d_v����L2�Y��x�[��IB{u�<9���/t=`�U���KY5��C>`h���|i�4^�&��Q>Kj�E��6s��+�z(�l��-����ji�~��r׋���;-Vj��b"ހ�g��Iؾ?�����x��Ɵ�b_�,'=�g����(�C��,�v�6��-)���T���z%rJ2��MD��\�Ivs֠|N�~K�M�	_ �Mwe��m>�<h�o�u��S�G@��D�[�H�<R�h
���W����\}.���<��*8�O=X������f�g��鷊����I!ZՕg�n�/ĝ*v��^�*��2��Jv���^�b�98L	��iN����T���Ej,�H6�H 5�8FR���Q�V�\�cܪR����m�͵�G�����T�?�+�W�vܙ�[n/�����4���5ѓ�K��H�ǆ�Z�%��誆�'ꪱZ6T�M��w �"���3���
��X~�}�#d�[�zxrE��eb=���P<g�?��䴯�	�4�B�ysx�kQ3��Á3E<3�k�A���RPYډ�z�Bw�b��QG������*�Y�s���d��~l5s#��x��Q���6)�i��G�fN�6� O'�Tg.�4�j�h��8�*����y[D�@�U'�wKW�j^dw�P���hFDUd!aJ�J�ת��kF�V�%\e��ϭ�FH��f2�0���W�cBZ��^��1(Ӈ\q���� ؒ/�)f�|u�^��/,�6� �)͐3��|l������W��a,����f�Gxe�R=G���	���گ�Yb�j 7�N�񉿥�.�D��TuQ7: e:�2lr�T-���a[����E�t���8�5B�^e����?���zAԮ�8��I1����l�9��2f��$�T��7��Ģ��?��Z�4�,,�d�%��d�tc�o�BU���6�������$�G��{tl�ܶ��u��\��u�|�2&-�9ɪ�L�~M7�J��b�?\Lb�U���c0�
R�<p>�����Fh����?��$Z �L9�fѭ���E����Y��nl"�D��Խ��޼8�7�c�$_|�6�vȻ�4�%��|N�z�C%���G2g�+Ie�� N�̳EP&�25����g_���cR��)Č��Z��U6R0��1+��
+[-*=�K)�nC;��W~A��ܪ`",z�Fji�߶W�?X ���5��g|�n�r��$a�o�+]�����^ބ� �(�A~���١.G�C
Kj�M�'{ϔ�M7�9�e4y=�z��E�Z�F���G�
�Q�_��WP���.�|�����~̷��m������?fi��!8�a�L$��,JRtw9�Kg���j(N��:��$��=���TƊ>����BY����N����s�Wo�C���wݺ�!��w��oPw�ͥz'G�+>/�b�̣�h��̓P� X�N���US��UZ}��I��f��BĚ5O��zr�uc��*Zb/\��>zU�X�(�T6�f	�{j�pǜ~+7�*�O��Q,��S?=�̦jV&�������gG�{�y���`7mҳ����Lqp�Y�9%�Kc_-�}���NB�eD_}V��:]���*e���$�Cnvq�ޘ�R�j��l�w������&�����qe����O�or�2���w�6p��ن*�P���aw����ѐICp�|��iw����� ���
�6�~s�|x�8`�	J]��N�"V��/$..nE�
�K���}�����ʛ���4�W���z�|-k}��S���_��������/i#ceDjB�k�>1�)����Z�*�MpD��g�zP���̝N�(&�6o4�L,�l� �FF?t&l7w9�O����ˣeg+e�������J����@wNE�!�J6�.�My�b�J�2p���ǁl�GQ����+��ceq�I��z������i�x�q
����G�ߝ�(�o�
(��$Z����Mm�.�����\���X���2W�Z"q��F��T�����t�t��/k�"�a���:��|�R�����GO�ZpCpи��v~���<�ʖ�YT���YS^��$E�и7Bn�������߼)�:� O���=�yrƈt�D:�K%�,��۟�U��2��7K)R]m��C��$tm�%M;l�E�+���l�*�qߛ��4�� O���Gw�y3�.I}�)��?R��õ��o�о�ߍ����DZ��\<,oGMK�)%�#�,�԰��V��E�7�W�C93��Ϋ�/&o�4�kJ�;R������!�$�X����n�%����	�bM��T]��1%3e#t�$��r�.���j.�N���;?Zu/y�3JïDT�ω���%�)�?�=�@M���Dz�@�0B���
�GŁ$�AX*!���g=� �����&�Rp��U��Ӽ���v���11�@��*���y��2ܙb̹lz���5z	�z�ky��f#C�r����S��K��h�p���H�$��cPƁ&��[})�f�N�jeЈ�M�붱����s.b�a��N�w�ƨ	�aA�	ӣm�ӛ�o+�^�˫Sy���[�e�խg��
�@�+t&&H�i)���܆ ��`�6��>���}!�⵰��W�-�Fx���<lq�%u�]^�E���OGhk��_I���Ƌ����-"OF�����InR6���$#���|����m"�.XP'Ј��Z�]ɾ�M�(�f�i����hޜ�Daq�:i�JM�bB� -�	Q��h�ϑ`n9F�4Q�q��m����<�Nǉ�*tIU�~	�[Ժ2�:8�8n-+�g��/Б��؟�����WN�dA�M� ?j!���`� �((��d�ʘ�-�'�=��ki^ ���6�i��e���sĤ�b�԰�a!�+�A"-A �24=0ׯȪrd��*�o��ܣ͇��!)�yc����u!^�NoLbj��x�-�^��gN��  BT-l�yF��C�����C�@h ����Qÿɼu�'��ƨl�$��U���6�?b׈«b�]
�΅����l���y��f ;��+����pwf�-�~�)Na�e�jÀ�'0�h_ˍ�l��Nq'�>:0B���[�*h�$�Ş�a����|C��QC�`����Eۉ,�8xƍ>���b��H��2����8�5c�Ӎ1.�~f����$ ���Ŭa��f �y�ð�{�J�|^�d�$#�S耣{�/�J��Ȉo5�` Śh9M��r���M_�;�}��L�0��ǁ��y��7{��N���}Z�r"򷑉sC.�Χ��:b�f������,+5C
|�kh����c�jn�6��������P<��!A���&}�.:ZC�;T@�ǟ¤+��mu�> �ؙX���POöQ�_�����ƚ�C`��GqW0��_)�[r!���x �k�.���J���䶦���r=!�+~�'��6�\!"u2ŦF�~/�Sl
k��\���]�襏���J����b-2�7o��EA���s��m)ް@np,�� ����f���1����H�-n��>�g��j���0C?g��n������Y)�)���J\K��,�3�?��0����fO��	�*iJ��s�I��.d+z/�����DBuy�k����v*:g�'�$���$�@�i%m ��<�%L�84�2�ڈ?��i#Y�/��韦�]pm���\S*�oW�U��ͺP�7Y���LJ+�eg���}�k�#��n3+VC��F|��#&	���L��)}\��]�sT��3y.'̀���F6���#\ƃ���Ԛ�c7�	��S��B�>��P}��A�]�����X�0�#��ܾ�d�VZ7�@~/Ǻ�XL'�q��g`-Nv����+��o�"���_5^���ᖎ�N����۹�c�8�S�[�³����[��w]���"[�MBZ��`M�~�����)n���3�M͌������mlD�ݟC��+�U�%�1Q�ۍ�>8���ӿ����m���@�e�lN��P��ut��tF)r��b_�~m���g,�����8ku�������m��55gD(�A��ݢ�A�E9:a�,��У�p���C���z΢Sv��(ĩ�}����V,�	���~�Q�����}�J�@����o���n�S��x�+~��+~��!�Q�ZXU�(c� �n�~��f�8΍3H�~oI&@����p�9����P4v<ʊ*b�pV<a8�g#��"ԓ�Q����qi�I�[�hQ��I]FR넳O�]����ѽ��9�;6v۰.	�#�v���ܛs&���o���Рڣuq�ޤ��J	j��U��)���d��3%*�ɽ
m�B�n�-1�'���z�%{z�<	MRW+y�βVĖȡ{�H�J,S���A9�p絑���f_(v��R0x�dx�r����p�I���"���D�	_ӎĂ�WGy�3E���^o3".�~���GV3�g�����%|��s-)�)��i�4���.�����❔!���,�[�R���5{�o�����Ŀ�|$�[��Eƒ[�>^��-�Nd���]�ɼ���!c���s�Gyسm����/+TN�>�[��t�Q�B�䗀�;�9�l��FR�(i��%�&�9�'��bL�nXX�f\���~����-K��P�+�W����D6=�0-���[�G¦{@Ti缆��ڦi���k��e'�0Cxۨ�!f\|�%�fF��y
N	?��B���Î':�'mn:�J��RR�ue��=o�^V�x`ʨDD�Ki�"W?{ �\p���ɍ"\E�T���Q�/��ζ;����T�nFdD�|u��1���Sy$Vl��5�1	�5Aĵ[+OoG;�~�(��0����A7�>�����)i>���Zb��Ƨq(����Љ��ۄ��d`v/@�"��G訝�'�C��-�<ҙ���~�˛����FQ�?^y�A�6�B��_�b�R.�}����.%&�@�HZ,�P�f�|�H�4���fb֑1Y��Wϳ�4���R;m�Yp	1k���M+wI` ~O��;i� ���T�.�Zv���)%4�/�u4���XT�$��/��������9����z��ޛ?i��7���r\َ�Dg�i�l���%1=��`��X�V�D���)���o;�&�S���~c�.�=���I�����P-�	s��s��>J���_�\F�}us7�:N���Q��[����vW���GQ�e�2��a�yA��T__�W6i�@�V8�z�-��v����I���&�t��a^�o�0�����hϳ#8Ht>����c��b���P4�Ͽ\���\r^��	>�[~wv2�h�()��Z������,��=��Q�vȦpgl�t�V��Kb��{���	GYf��V��#Z@IV���9���۶�"��2�*�YF�i�T|fy)Y����}��*�T�@Ta1�,4i'����.�c �:m4?LHl�,A���Y��p$p��I���uQ�����M�;�RyU� 0�e����/b�0��8�����reJ!�	x���
�qr��m �O�����>���n�}�4a���9]�	��,|����}�c�To��A��l�3��O�Bt��2����r6�I?xO2���A
b���-�H�8���X��Ĝ@�rH��{bp�QPˤ&����T9�|���Yl��eD�,ý{���� �����^\����V�n�v�0;����{��88;X�3����m�?�zt=3������t�+���[������߀�|=�<M��!,�&�����**��� W��:jW�+G�v��!�r�k�a�o6Qv�#��c�x���k:
e�2�ST���T�qh^q��vWK�7���ʅ, �ʢ!D{�q��	<����WB��cs�#��`P��!e���������@H��K�`�˟�ƒF��z�f�^׆z�a|�6�vu�@<�_`*9%�<��<� Y��!��v�4�š=�/��EBA�/��q��8��"�r�>�tx�����88]���@��*���ܽPJz,�;<������U,x�x�nLb���F���>���@�$ߺ�W~��P�7&�� F|�'d���A���D���T�˯�1�;����㚪�^M�,_E;*t�� z<�:����5c�6��S]�_IE\n�r9M�߷���K0I��r#]�?��ia�&����?d��̞�������g��k���ۿf���õ-v8Z�i����Noj-9<�+�1�Af},y�4���Q������L˲�Z*�8 ]��0p��_b��B��Ġ�dr�U�����ف;�U��@d@R`�71��N Tt����D�S�Ev�����ջ��� ����t��:���cO-T)2ߖH巗&��	�Ԥ��b�%<���ı����Bv���"784�^��m}>���F�Rs�%���"���U�r8�
�s�j�&��#��Dǲ27�p�&4K�����Bp�Լg-�\Z��^�1b�F� ��ӱ0�t�u�~B�r$Kλ* (+(�\�?�ݍ٧ge}�l���V�&DZ�lb�[��m���>= Pl�Q�I��S{��w>�k!��(���$l�<V��K�^�1^x��	I&�ċ���X�����&��@?��+֥B����������a9= UHf�@w�[�ݥDKzN*�Ȃp���) [C�.p�#+��EZ���.�C
�'��}�g��-pu���*kd�	]W��&��p���E=�g���hD�������f� �L.��4�X( �:���j�j���M���n:�1JB�՞��}���r��C*h��s�9@Y�yNy�<�h�i��+� �\�Hg���6δJ��wVr���Uޞd��M��#�]��_o}y�V�(1i����y�F��z�?!)<�p��,�) a�����1Z
��;�������_�୍�k�c��ޖ��/
Q3ưGm5,��|���?F
F[o�_��	&*�A�m0���\��w�٥�j7K�ኈ��=ܺ�m5��}9��"6��D�P0]d�ɱ�f�jl���K�i�r '�w���ܛ%��A֦���І,�;������I��b]����@�,q-�UN��Sday��]�R�������_ߍ���� )3�z>$��x������t����Z�ăCp
���xJx���CDJ��V)�9�qVn?A�1E0���3u�x_b�A��n����L��h>m(7���7#'�ѫ`�#WS�k�'͐��\��O���u[���M�6�<��ұ�o=����iυ]Xr�:o&�Q=<�������x��*���-�W�U#��OQ��P*)], 	].U؁��A��n�[Yx�StF=5�v�Ijc!wmڗ�v����Y�t�%���M�����^Ⱦ���"�Ӕ���V����4�ٯ�V����G�h��?���t(1����ن�?�1�B�o�~�J�4B���b��6x,ܖ�h�ԓJ�5eo��񴓊�6H��m@��~,�e���<�@N�f!���(mF<��[ʠ\��F�9��#w��3T1�t�����J�L/�*_
����o����2D�	�5�k���N�/�a���7�ͫ/�h0�Ah��[������K��:jt���N��L ��.G�y�:۟y��xh|X��D���Tȧ��v�2KqC#�/�w87f��i�;�9)b�1Bغ��N�����Ē��h�'�����)������p��o�1�Uԁ�R�����|3�v���S��3k�FR�o�NW��k�}^|�0�b�(.�y+���e3�����cB��ֽ�w���Q�5|m�d	��t)y:|�
zB��/�-O(��G��3��Z�4x�ȨU�H̗GRàq�W2�wu��̏5[��������)� ����g���k�*�c���1Ǫ:M�4h�j��5O(�~�3C
T�'+2	�˶Lg���l�u���X�cD9*5UF
VI�a"�E�S�����T�r�6�j*MC�_���y�`	����k��Υ����F�d�e�WQ�����B�L L��@�+��s3��At�c
�M�=�=�LW��a���%���HN�[��U�q4���|mjTzm-����L������]��a��wܡnY�x��a�c_k0&�?3�"H��D��z����${ ��zs�\�E�����1Dz:�$�)Q�lh 0��ݍ��
�3�����\~H�(�<Y��O*���B;x�����2�/��)����%$�0�D�5��/Œ�i�,=!o?�U��i+�	�k�&Q�¶	�@�4f���7!su�?�T�]	?e�rh��]^©)���aT�j��Q�j���_;3�^���:5xO�ࠐ��r��"X�_��z��w;,sEN�4>�CǶ�hx���T�no���}�)ʐ;ۛ�L.���/��.w�H��|�BR/¦�j�h�����X�2�� xY��I�D�#�N�7e�_�p����yN)��#m��y
K�|'��M�ax,�u%��|_�fѓ�?��1��: ��[_���)X�#�淧FN�(���߲̊�� fP��t�'��๯��#�pS��t�����WVX��8ƃ�8u�h�n��c�,8l�O�Yu 76W¸h!mZ���o����ABy���o(���n���t�[���&�Ƣ��)�ݸ8��K<YѶ�p�s`���B�[׷}��|/)�K��A@�h�<=��)���BppY�Y�+Q�|(U�r��gd���n��L�mb�,m �Kݷ��r�r����
t>J�9�(m�[��s�V�LhBZ59tvýW�,A�=T�u�
G#&�F�H�٣ִ��(�"�֢U�\@'#��m�+a���	��\K��8�T��R�"�PB���"�0�C+|�������{v�OF�
Xgމ�ٝ�6B? _�!�P�I�����;���{�T���/KBD���U1�� f|�������˱�Q���=QG>�ь��^/�i�LڼB��;�?��T8�;���LK����;�愐(H�k�&)��-��<o��@IO#pW=��*'40;�"ޓ�s�0�֍���;��H���G�&N�0���܏a�(�"����[Et"��=����A;��x��e=���'�`��R�U`�������@_�T�
�C7��t�Ƕ�'~$��f���c�U�j6��C���K� �B�ꎵ�/�e��a�/Sa�R�U�&��kۦTq���`�W��)�$�O/�����s��9[�?j���57$��.�G��Z�fh���KXs�m/y'E��Y��2{· �6�ao����j�,E��r�^;�m�x��%oZ��V�>�Ѧ����Ǚv2K ̸v���-�������g��;1)K徕@�����6��\[)���cf����T*�#��A`�&7�7V��!�seG��l*Nb��7Je�?>�uP���A��-�Q!q�9�I�i��&�v�$��g����7���j�o���[���q(�#T����`�98��u0t�tJ!Z��|X�0�*��\^�R	f�~"|�����2c��~���PS.�>�0���Vg�.����|��.J0d?6�;�&�����<�C�d|tSwS�ͼ�X&ޚ�D���kK�1�qs�$���.�w ����fh�)j��d��0�!c#�(:���������K�܃U�E�!���7f���4t6T;J�K���c�Wr�X�S�'75_�j�B%�h��p�b�2��G�ÿ��(��l�ѝ�;��|��fR4��Zي������*@�V�>����E����a�����p%v�a(���j���x�V�V!+�=sk�qsc��%b��n��+ѩr6_���&������rOE�=.��TE�$�bST���ѳ���f�'S}��^��C����U�fˍJ$����;S������W:l��1�DD�B&��ΙC���o;�����l� 4������Cc�r�g'�
���V�j�o��%��V����|����v�簤�i��*�OM?j`�w�4���3;�͙!և�ܽ��O�N��J�o�hI6���@���Y��Z��Y�|In	`E�����Į��J�T�[��*b5���R+����3��s�_�B�L�B�܎����s�{!���-�|r�+��qD��WE.E]���G>YjzH Vy�Q`�iK	��� ��E,���Ɛ}��Xh]���Ui��"�hz/��nF.v+�P+��$bNM$�8"s��dA��61��k�Ü��pT枋�1g)��^�Xt\�u��ܮt�8˙�.��NI�S;��K�E��i�+�;9Qh�	чaGP'���@��J�˽�s�.v������Ŵ��
� �Y>�Q�p�(Jf�+V�%��R/MO0�fbF�rȟ�6�L"_��b`9��
��3�54{��p���&J�1ʠ5�rΩ�Q?:����FIଇD3�^n2D`,<� �v��d�ڕ�]�*�c�qR����s���Iپl0��Ԙn	�^��v7�����/��X�����"V#и ɍ��!��:=r������'y1��l�(�
�.m]���L5�nѾ �L�~O���f�r
܃*�`�!���h�uK�S�me���LY}�8f���'��d�ܥ Efr\���:���D�CY��*� ������i;3��hh1@�K��j���4�f��ou������C�r`]T.���;��E�-��P1�7��<��u�,�ʻ��X�,o��5Q�GH�4`����H�|EVS����m�;8�˄wU0$�5��G����s��t6�K��K8s�
>Y�����9�
㩲���,3��i_c^��z�Q&��~�s�]��k���d�;���/�q3�JLw�x&/ײ�'8!��)û����W+���Лif�]NB�
2���q&Z�XN��R���D�!R�  ���= 9%Mb�p�|�Ɂ�W)J������t*�<����=l�]�*k������e�g�t.�HhC�ࢧ�7�}K��l+ᨅ���\��k�d�Wm�.),a<Z[ɿ�Kd5>�Q���6����9��_Ow�������lʮ�e��t���iY��N���Ⱨ#8̛�2K�����	0���IP0In�j 1<O���2r�h�S�2�X��>>�}�[W�pX��s�c��3Gh{�:�9�v�r�2xw��/y�{ i�q��SLi!�Nˤ�ˤ��?���F�/���p���W$-��ꮦ�E��'��*��2 gOw�"i|��?��gӚ���,�.7���\k'��5�k�g�q`ŕ�����L������aL'e���`s�&"�%���� �zv����?����.QM�9���,/vGyM�v��Xh��`E@c1� �C�	.S���h=w@;����"�[;DF��ųw7�� �V��@e�~�R��Ⱦl�/X�r��n�� �����A�-�Edqx&q&�d�W'S�o����C��k�R�=��|���b+�;!Y��G�t5��,��b�$���,5�����8�Z=nsĭvk�
�*��Hߍ+�X{��B��G�f�ȕ~��3d	��HГ烁�0`�Ќ�$��^ WuTn<�V���a��ɜҜk9�:v(N&����|REI[��a.��5Z��X�K1�܌$��.��Fh��Z��{~cX�5��+����v�S�_Jф=�4�E`a$W�5���o,9Ve��/�8�=�S��^}Х~��L; ����{�������F�\6k�ZfA8oi�������2���:��U�	��g�/SP�D~; 2�l7�]<tQU�dڂe�tH	lW���y6[�.��,�	��1�$_��q�V[�r�"�ֿ��7���T��V'�T3��b�ǖ��as5�Q���w��-�~-d>Y�?�1���K&�/�R��3��
=߬-��hǌ�L�����$`�=/6��$� � 5M��p+��C��]��(��!y�8�5���_����Q��P*�:�9~�#������b��#Ӷ)2���N;��b����"'º/⻚�I�Aڟ��$�v�����W��#��`*f�����KlO(�(o��E-Ʒ�qZ�?%',�e'����r	�Kc�TZ�iV��X�瘾��<~q�T='٣���S�mզj�Ȉ����K� E%j%2�h^}�����`�M)׷��eo~�s׃��|�[�~�,7�$j?9����d�w2jp*Js�3���(�i��?#J�yI��}u��T�Sؘ&�5�������r�-	r�[e��|�I�I���䦁vһb�|�-ժ$���!��':�u��	����)l�|����R�35��M,^���C΀@�R�R�.Z)����cB/��E��"uf�ࢨ��hPU@ѫI������`(וx�oD�:��v&I�"=.-
�a�1*�Tu��zA	0* ��>��yv�C�*�/7�8c�@M��#P%a�_@�������!�U������o;
MF�;���^�QXj�q�ҫP4շ��8
zW�V#�3Ҧ1��|�~��C���ii/u�X������@@��I���{+Q=��������,/�L����O��6���c�,���]��z��7E��?�Or�m����%��sOd����A��O���٨#p��:�"�5å��-��vPj^�Z]w��
d���v��-z#2=����]gn���V]$nb���	2�k\0��IED�U���ps�5�:b6��!��1ȆNR�L�"�hkϢ�%-w��rO�Y�x5��������yo����LQɼ~�S���0�T�3�a.�<�Jg ��,j(��40�[n���C�¸�Ys�捋=rz���e-�׽DE�kF��E ��`�-�X�fB�XEc�E�S�Z:�@�����e�����˟��ϤraQ\�D%�1�I�:t�1u"f�-��!�a���5�*��.��p3&Uj���tl ~"�����B?�)�aK���q��/�F�����P��}~f�UVE�>_M|������;&��3[{�Znh�54!% 	A\F������1���ʚZ%Dir����H�N�j�,��=����iY\ju.L�ڪͼ��.s;����g�8�>���Y�z��BZ2�o��U�̐H���{&�H]D����N��0P���R��WJI^pw�kab3Q1�i��f��T�=[1��"�pFK�4S7���R�aB�݅i����i�j��}V�ߠ�b�Cr�2���M� a�&�:���1 �ˆh��G�S�5VְF;�P�B����7�e���H�>� �=�()lG�έ#�C�TY�/�%�db�+vU��<��M洔�&��\AIoa&]��T賬�-g��� B�9C�߁η\�x9�� ���?3��tL"���E�d����9�[A�:v��K��������-Sj�y�5��Ա	j���5�P��󱛴4)D8f9w��R,��r�<\ײ먑r���K�r1#j��-�T}VQ�"w��{N���-V\��0�dq���&��>u�GW���$Ss(N�����0�h�z�l�U�"����P���l�V��Κ����`M]����1����=-&/L\��$d��7�Ȕ)�+ ��Z��Q����:癒8�WZ&��2��*�v05�O`��<EV���a�)%��O�p�o"�/"�JnO9�TB��>%$6H�y��X�˯R�o5R�BI�t"��U���_n�Z�Hu��_�2Q �
A�tt3=D�i��m�,zE�ppx[����_��{�г�K�⻭* �vF6̯9����/�~ �̅�ݲ��1�s��F�M`r��څ������ ��-��>#��dY��t�inɄZ pq�2�_4�\�䓶����e�!��Bz|K��A����#3("��G��y}�9ڶ.u���d��'�5�q��餳Q�s ��C*�9�6��R7�e�ٻ{��oؤl�HA�k�@���IH�LR6-w�z|��t^�'�fZ����3���G�z��y��
J��K�ˌj�l;�0�Zj#* ��єe�\xVX��
ІU���Z��h�b�Id$d�:���+roʝ�b^��z����AzEx�U��6�M�}�Կ��[p�)��D�Y+���h����G�&f�幵��lИ��rw�њ�#��ز�nh<Q��#^�,P��]�5��'
?�΍�zF� ��'2� �.Evh�j�V�DEфU�gt�3��+&@�׌
���g `_,�A������C(� �y��ښg@E_���4��j���^���%��D�"R��?C �JJ�V)�kԉ` �<�u~:��`?�ܑ ��*�e�('y���$�8놉9U������օ]a��k`X�N�*Q2�?���1��;���iS R�N�r�OlG	����ŜS��o���/*ʷ�M�X�2��X'�G�m+�Wx�1_�x�~���c�6��M>]��o��[�驝��E�b��E^)�⼑1:�ӈ&?�C�Y�Ru���f����|��#g⾨��,��Eʝ���r�u�N݌��O�&���h�	w�j��a�;qO�\������Z\�]EO�q���A^Z�&҄��cEqa*����`Z]L�����
h@�oH!���j�ж ���Ջ2���u���nz䅍Տ2�e��6kC�4K�7�x�60��C��`~N�g�¤�݌����p�ͣD��>�c�_U�DE�`�79���F�-T�;�՚d��sZq��(��1>X�NHs-��Xx��m�xg�H��S�n�r�Aq`[k���V�x�ŵR5�ھ�&24�g�?x9,�JLc�pug7�Gp�2lF�	S�[����)��v%Ak�Ԯ
)����z�,5�u�T-ܫ���M��T]�w�a��B!��S�f)��̮�����F.݀A:�G��t<E��S.h�u�e�G��O�CIE.�w@g��>�4�L�=�M����G<�[0�J�|�8��X[����َ�JhA�& vR� nk|��}��qU�A�B�5��{g0�U�	��%.k����W:�����{ �b��f�:�Mr����"��������w��λ��}���8���Fm��b׆��@�� <��"��iDj�?2:m~$�}|%s�ԫ�a�qY#_@5OFʍ3Dl�m�� ����5b�6
>�y��B�5nl��'6�#Z"�W�� 2:�y���/��teX*����8OkC��������w ���DC����?\�n��]�Y���:�K��aP��H(_�m/�A�v��g��hj���� �^5])�$��@C�wz������U6b�@h �n�3�M�O^�$���.�a2L��6��7��S�AЫ&��<�)�rX��w㰽�*�s���G[�t����1��jg?byaˑ�H?̪�x��b�m���YK-�`���c�z���zb��G3=i�As��(�� ��T����\L�K��n�}�3��h�u�Ĉ;�A<6�S"�v�υ��niҀD�Քx�nG����������P#�WIc��hT]�!�����e�W0�WI�m&7�����^�!��t����V�Z��b��B�KŚ8!g��&G�7!��y�b��[,(������Z+A)g��B]E���������1Э'=(�u�l,9��/�������t���B��v��L���n�� [���cʢ�D�1Q�v&�:T�Z�~��(��(�����{�n����'��L#�h'��-N"�¬�?�}�~_B�A�Ƈ�����LJ�cy�	 �'Q��d�T�F�ҨP�k��VO���<��cD{�r��k���H#\A�r����	Rg���Asܳ`>�8�~�乇�c�5��h��+Ɗ_�S��ll(Q'΍y��	l�:���[(�f�au�Zg,r%��H��靅� ����2���o3E<�o.�t���Z���s\�w�Od��96���J���U� �N#����3��D��t>���vW�W�4,��F�����l�虃��f�F�R_����c��;�Z�.�S��� X\�[RP'z��P)���
��n�3F;����
�PXWi���$���>�ފK�\���s�D���\��wy�{��h��<�2T�l/��S���DS;͓�g����K�uw�q@�h��XII�U�v�ɰx[�7�G�u[��^OT��m���v���b^2����a�/(��3�aF��x���AH�����+^pG�� ���Ρf�GV���N��ER�.c�/P��;�|3��31���n���r^}�[�L�`�T&M�5��c^���Bj��,�b���3D���g�"}R�D�
&6��WD#�<r�Xѩ�oQ�KYpl����YOV�� 9�O�U����;}��+�����V�8�	j ��#�Z���ͦ�Bt����G~RI|7D�$4�:�`$�P�5A���oR�����Ǫ1r٧h�U�.N��7-7�B9�.��� ^�X9�]#�
�K��0&�=V���Hk�3/c���Y�[kL't�7�)��O�.`�E�D�UD��?2f��/8r�p�~�#�V�4p-c]��Nm�����30���)�-8П����}mؤX%LP��s�!Yed�� )�K�9�س����<�Y���[�P�ٲj���q��A�%˻{\�V)I��f�H���`;]O�T�P�g8��-���'�g喐�OmL�"����av*��B37�p����X�-egS�@��8��|J�(~1�y�s�]���V8�=fM�T��a�}�c\ю�M��G���ʤ�1[݌Ix�lX��og�@��
?U�h3����z�5�55_QMi\��n�`�;AFF�d5] Y��p��%.�`腾�������x+�I���^��\3X��1%��{��$=�nf��/~������qs�|�m�]<f�m�EbF
(;H�5��=�w���s���FH��|�j��&h����a/f������|�1���]�%T�� �Ze�̫��7[��Rp�7���j7�0E�_빲��#'6��Lr��A�&�N0����n��Y�a�+������^^�n���:j���c��⋶�����N��W������=�7��/�(\L9s��-��Q��px�>2|���Khv���A��gx��ָM��57�E^�+7b��=��0eOn;��+�1&b��숩��UG����K3+�?+���H���z�Sw�N�����ob� �|���tA�����t���rT�UB���5;lK��h�b�����&�Al8���Y>��XC�7k 	 ����v��J�0KQ��4�H-V �����nVb�r{�"��J*�2ں~'�!sU(Ŀ&{ģV��O��tbo^q��C�5c
�Ԍ�T]��8�c���*Dn��%�ذ[306w���rY����Z��J�?h5������~��!���C�i\�J�M�f�l�7o����'qg�#݇$�-�YM;�
���h����،��W�{ד��H
�~^� �[�����t����p��Ǌ���8�Q�CuǼl�)�ck�/�*־��v���ޕ���h?�է�uǵ�����h���z	ws�/	�]��+��U�����ع�C��@pH�%gT&��]��.�D���1:�Ȁp,(�P���\q�<���_KХ]��{�ڑ��l�(�.>y�ēN�|��gKaC�`�푸�&Y�_���B��Tf+h���I@���{�ۛWZw�`O�r�a!lxӹi-teAgo�=ۑ���^��@{%��BE@H�!�N��D.t�ü�&�8�^~U�u��2�"{�[�*��t��hQ6��쇈��͊2k5	�V���V�I�㻲	�/y@n����Xf����cO^8�L�\�~�3-l�)�~�����q
ڪ�Yp4�e�Fu`���%n$b�r�A���J��!�x�Y���U�P���`p _>r+�2�kA"5_�Z!��V�U-h�.��W�_�����"�T�=���y����i֗nDgk��^�kQ������`s���0������gIQ�^�2Г��bdi��
��E�x����&#�0de�K{V^Ҧ���üC�F*ö��?S�(𝫧q��7�� %��/n������J�B(�q`���W�'[)��~��^�Kg��t�zR�ok+-m$�����9����`���Dj:"�&���]w����`h>��C����&�BT��l��p���lF�;A�:�ۢUHU�Ԟ5�(���G��.�g�Wl%������M9y"�9�X����dal�q'!��H��;���l�!���r�q������.�n�n�����l�e}��μ�&kHa�C��'�{�g$���H1sLǡmr]���WB�I������_!D�̽�5�y^%�z��B��V�dSRE��u���p�b��@B]8_uRș�|U��%aH�C&��Z�`;���`$W�;�mbR����2���R1;�c�e�۹�|���F�)�[.�W�M�j���~N[D3�F�Yz wB�F�|���s- �bw<�r�е�X�����0J�A����O�Ϗvm�]��i؀�]���)��Yދ����Qz�yD�g����.�~X�()�W�C�< Se�g������xa��20���d���3.�l�����FM}cC}��7j���)9�|�
��o0�����rr�T�aC��ygaIxU@�3�����ۻ�,�a%K�e���F*�8B�v1�CTw�������˙ŷg�E��i�bĸ���k����R�E�ᐺs��'H+�n��)�S��R?�Ik���i�[��
\m<|�5|��F��F�����s�����o�%*f�I�4	�k�2P~[�`�%����`#�'k}����[��D�Vo���osSX(��tz�)���<��I�k�'�OT�I��W��!N�$@�ǲ>K�,]�R�"U���V�q�Z��M�kf�&q"A���F�
��n��A�(��S3�%��$��h�*�x��<;m�c?;�'�����p�we	2{E�	�9�H���q�X� ���>�W�|:�0xoy��o�h�[#�O�¡2�@c�g��Ucx� 0� f�$<����A���fCN�
W)�k��σ�x̙�:ۘ^�����:<��������;qqb��q@��;�Lz�7�h�ʔ����m߭�+m���TR����ì�ތH��\U�b��Sob�g�Ty[E����>�^��k��"g��(<�[wj�Ynݥ=[��k��M*Y����hG,�YyĥcOn�@��v	�KÕ�G��w$�.%_�@:I�9h9����h��<����+i��O���iX�7�U,�.��ϴ�bG(_0×�6���	�tԭ�l�%v�<��6���3�0'�de��g�{Ar�{fr�#��#rԸ�c�m`�\�[N�����wߋ���%,��w�ue�w)ڮl����Jt�+�&��RY	nYs"9y����mF�%������]:I&��G䜿G�j����W��t��:Gk�K(sЋ���0��PN<��;:u��B�����n�oo�6���{H������V�k'i��&%�(9O %��U��
ҖHGB]���[�Qm��f7�����z���k�5Q[ I�'�'�$��\ኵw�{S�Z&L�Ȫ�sv�&{\
����,ͺ��	�G���NNn��W�#
�XV��j���� T�q�3�P˛S���-��f*�e�7��Z��M\� ��p��Ĳ^I�=�N���٧�0��I�������0��%a��@��T=?�C=��ya�U,��^���D�z��;2�v�����`~خ�eq���A�xh�I[sg��:��_�a��;E��4]�(ob�+�W6�J��q���+�r�b�ÝH|`c����	�Gc�s��\�U�LX�m8'��l�|��D���P�	� �%c?#��,��U�#RQ���2�� R��O��/��<U��	���^bs�1&fbHȁ�r/�2�B����6���X%~�ܕ��ɵ-��&W���r=#D �v��1C�e=�� Zؕ+�ڈS�p*�3���}���w�_d�&����rO��P�+�����c�1�t�3}�����M�Y� �b��qO@
�P�9��V(%�2Ȧ~a���c	��q�J ������ٝR�'�q���
�.{!�w���'k)��ɋf�_"b'�8�q?WY���z#�$y��UC�V
�c�1==2���A?�s���L�˼�^ ���������0+��\T'Z呻L%�b��޼Rk����vǿ�rV(��ͅ�}i��G�T�/��+ꑫ0��7m��I�GG�Mǂ�w|\4}��q��"9jL8.�c�I�U"is�8�����98 �����ἝFr�(r��tBGn2(LS������Ue3ޑ�Y�!0]2=Y�43Ky��1Xe�l{l�����y�ՂJS�ɕƝ�Ҧ!�n��Fc��w�z"�kRl7�R/g�뺜�TB2g=���~}�jZ��¶_B�r\�Q�ԟ��"r���W�]�V�L5~뀓qѡ{���.)eϮH�iqN���f�vs`��|*�6�;s�QE����֜�D�_A�� ��,~58xf賊b����o��}�j|Yb���2<�(�1x���644Ip�R(�f�C	ʑ���5}�=��D��u�ַ�q�d�k�S7<�as����*�o�$Za"0}�@p:?!��Щ�fR��Gr#���cbn�㖨�5;^�K�si��tz1x�8ɸ*�t8�?o,�,��~P��x�7x�����7�ƅ��ZY�T�r{Nɺ9Ү[C�MǑ|V�v43�&P/�j�`���ߩ��_������4R'��h�#�":s�p�Wp��k<0:f0��B}P@#��B6O+��#�e����	�ێchPd�O����b�>&݈��[T ���^�KɎ.�ywAo*Y;�j���a���R���#Z�2�Gq�m��|�u�r��J�7y���VCna��n��]��]@z�N� 0�#IA�h���"e�v��8$r�-��=B�]"��� �,���I�O��ej$%C��Umʀ�6�f�	�����'}�(�9�=��;ѳ\�:�k�/��3}S�a6<@&�ģ��y���
���!}5��^f�O���\��^�
{��W�&[k��x ���2�2��	��$5�&�r��/�IP��01�"Rհ�nE�W�kp~����OGY^�Y���'�ۃ
��^2�ۨ��bC�çc�|�Y�W΃�QH�w�B�dܕޭ&8RW��ϋ� K,e"3�⣲�[A L��r�˛�DX��a������⊲� I0"��(&��W_���~v�yd�4���J��`��J��g�P�L�r0�kES52����J�Zk�:t@��}vC�v[*m�L�<e��4��zQ��$��M�[�5���C��U�IO�>�����0z�S�����A�����f��P1�)m�2"�%E� �gP�,�!MkzI"�$*5��$�|�����)���>Y�n�F�)�ToɺF�v����s�G����i�q��l������.ڒ�6��`%N3S���s�k"��s��Q�i���I>z_�Ł�>�NTo.;�"����$Ceb�i*\���S� ��`(����FpY����bN	3�`^j�n��/!c���A�^��f�0(��#_r�{}0�q��ZEi���ONmM�N�W䢴�(7	n��W52� +r]�&Q ���W�M��¥��ǿ�"�I�?�9d��0|,�$%"�AKkA;���#+��ЃM�8	@�5-_�pZ�9a����^�D���8C��W8h�K>D���U��P�jޒ�+���������i��	Eu�/�rQ*����
F���){��&�ji�:��
� ;�����7=�ڽ��R�n���0��K�	���&8م�,0��t'�;���ɶ��hɦ�F{��F0�RfG8J��v����+d*��{�#Y��Q��� i�F��N���$"�-��sgXA��˽7ux�	�N,����a'��dVQ�3��,���#�J<Ek�:{E�Ts�8<�ܯ�����R�j�����\��G�J��C7�����"���)���6>U-UO䝵@�5�b�W�<L�E�Ϲ�oL2@��=��W������k����4��|��S62?CaT����}�/�4 bz�b��/H����t!a�^c9�i�BQ��:!�-0�UǊ�`oM�� �)��'Sm�Bz'�D�I<�%R�v]'Q~ϗz͎�c:���@8,���|�Z�ۅ�i�?�!�+�J���
6�l�������ʦ���шt}�~ֱMO�>t��q��{�o�C���K,�m
3�R���KL��
5���w�z��[�B�kp>��e�A���_n�*��MK��l�.O�%)�v���oц�Wn7T$!�h���q���|̣x�̱�cj�)�e��[��#���)��O�CT�h�QxF\-�-a)��ػ��Q�&�Sd����l2�`��)�Wt,��T��|[.u��-�	��>���1l<�.�S�?�7=z,�O"V�7�x\��h{�:da�5V�s��}�J˯�gVl(c=�	�3���ٕa�{����Yh�w�Y�t�<�_��<�k'g���L�n��F"�
�ޣ ���#�%[��&��ۗ�)K�豮)w|��:@W��_F�ڽ��<��ո�'x��� ���s���a��3����=���/���1����0����J��ȷ UvM���ٱ��<�)�o���\���W�G�Xd)�4���X*-�%a�'�����V?�U?��'��%��
߁��X�蜯kݍ���'�HW�GIuE�lĈ�p��^{w��d���}�U��n�Ft�@�$��΃L
b?+�NBIj7r�teEa|d�Y�V��-g��S��h�͑�,��_NC_��d��9���c�$ʀ�<�xj\}ъy���rb�7$�z��ŵ.+m�ʀ�i����Wo8[��	��h%�zS%�]h��Kl+����p��?>����tg�����W-�+bv .�kؖ����JZP�	c�'���]��J4�S�6�8���ܻ)E�B�Du��Bѻ�����8(S�DbO�N3d�כ�w�Q�+�j+�&���rɟ��.d�U�y�UH���/&��cP�x��x��`�`A�_	�Oc�^�(y�~�;��l�)�c�:ŮPiB�$]���|�f���'ݴ��SnQy�,R��s�����^p�a5"�T7hJ�k�4)�p��i��p"��&�s3�����h���6ۺ�!���C����:&1�#;��^�	����u���\��b��j�C�?/S���㡨C��*g~�x��:�oA�=�:b�]|rK7t�+ #>��m��>cM<o3�r1Z�i��%� �Jg�w2EK�[�*ؕ���7ƹ��?�h=�>��_�HG;�p&j1<CNo!32�V?Y�c1��ᩇ��Q�?->9�HJp�_�+1V_v�'D9��ɘ
�1t����'[��H�s��?�A:�7>��v��R��2EVѽ�����Pb�	R�ls)U�6����g�f��m�k°~ss�Q$B��d��D�F,��,��v��p���m&���QW��|'��TX,���~j�bf2>6���t��M--i�:/�!�xnD?����kH�V%tDh*?�g'��G��B�����J3{����U^�"WC�W�9A$���[�>��A�%c�*G;2���Qk�I�s�Ɗ��X�`.׶��pV�u���T��@��@3N�jY��x��B*%'���$D6�<ɪ�[w�9p�N�>ȨX�"�ϐ���W�W�GA̙g����(�f��h|l�S��Aջ)9X�\�\�Ϲ�ud[��V��gnƩо����K���l7F�;��D�Uk�0w��cs(��G�Dr��FB��Wr���P��5>�g�.�� o[�e�a�F>�ǭ��G�D��R��������|7�d��zri����9O�3h����D8��Ood� �D�i��8�F��)�g!��jS��Y�9+I;I�N��j�yp �5�.�ހe�UU�*��?�᪲�΃P3���`9�B�p��k|�Q�b}��j��Y[�T�C{I�Fc��Bp����4< ���L{����H�'�e���k��14��	�{����M1�L�f����z�`#�Y�}�,	>�{`�ۖ�ZP`���r�gܬ��%DӰ��G��
l�� OLs��t�n�vS�C^��+��7��
�	v.+g-T�W�@<�q�	 ����#xw�A>{�,�``��ஃ� f�����o8;ۊI^�8g�*u%�媚RW��tE����r�t�q4���7�?�c�����;�yr&��W�C-M5��?=��ጟ���ԝ���:��ӝJ>���Ls�(����3-ʂ�S ���<�B���"��6<�e�}�'��1�L-�_�/`�R�.�2�[�Y� ����,=��[�O{ʅ�S����t|S8����b�Քt>N��,�N�w��T��.*�P
T��L��FH8;�|�{D�1��~��$�?�|5Xrh�r&O�O_�����%��C�c�}@iː�E�3]��B��Z�_�d���������p|	�A���F��V��P����]:�5qH��n�+�9ƨٽ[�˝�{�.0�9Ad�?����n~+�@�X�,If]�v������S��l��C�H���KA��������%��#5�f�T�����c��|;շ�t�����DVL�Ɖ�`�tS�xa�&i���v^p���g�[�>�få�j;��;Ս�;b��ꤷȣ�K��x�8�%U#NB�	r�X�i��D��L�����1�M��ǡ;�BP=B��F�D�V��	�?v��l�$�C�I����W�~�� 3�=5@p�k�eOͯ"�7R���PM~̏�Z�u�U���"�VP�-��Nu=u�$�[�Sΐ��X�<5
j�Mb��ƶ�r3Fv�I�4fd�kq�#[w�i����L�f2�>\����(XV^)�$̞=�I�����:U��
�p���^��|�B����K֟>��N��lH��aj�	rGY�ǖ�N��h�C?�a�>G�SP�y+�����-p�"YBV���
T�3�lO��y��/(�cKK�C��?!g2�df�g!�;C�T֕�@��G�65���Lnm4�����I�"?��S���_��cJ�1ߙU���Qd�G9@�5ŀ�%�,Yuz獼}(�f�$�sE6?� ����ؔk?���	ɾ�[cd�H�P��<aaL�v���\�z����¾�p�/۳�e�c�2�W�n\0:#��/�Qݩ�R�����}m�;��H����}k�,Ҋ������A����'�h�=2|���K�w���6H���t.+c�ZS��9A�s&#�9/ҍ����ʻ~y%��5 c�M��7��.�G�t�T����HNPh<<��E��@�C�
���W5��A�-ϟyUM�y��nN!���)!�Ya��=vWG9���  3cNoʬ��HT�����I�W��ع}O�=��~��� ��gBg��ǹ�WŚ���'K�r[���~�t�����e�B�
� ����Se k߲��[4��}n4��+.���͉;��n��R���Z� �*�:ޚ���!�u *^�`b��~�F��oR:�9���q3�Њ�D"����]]�_ <����
��t:V�zPE���Ib��@�M9��"gT���nH�״� a�{|�HK��]�}�{�Q2�3�u°h)��@Mǈ�"�M��g�Q{��U>� ���O2[Κz��vX@�t�"
�� ?�����={͠��-|�?拑A�Q��p.��UOuí�a��F�W�������z�f..aĈ% ͹�W&Q�>A�����T��?s��� ��8�������nw������L�k�R)u����͊2���y]����#wSb��s�/.G$�ɭɲB�N� *
&rh�zA�-ᝅ$��.x���?�+��J�� x�gMByˑ欏ˑA�fg�	_K���X/���4ے��nG�y$��y��1�c�.WX���m�y��5ęT������\y���=б˧�xs�qA�	�2kzG�H?�\����W�˸���݌�=�㜆AY�^,�0n-S����[�$��Q�)<�l�4��ޞ�
3_�������g�fO����C6�v�ݔM}�$/��QA��l��Xj#�k�%�$(���ǵ����ـ�9��ʈWdj3�q8C�����З��f`��=P��)���cS�T4`��R���{�c����v'�����b�9=�V\Z�7m��In��(�z�q�/'�V���ɔR�w�d�-0��;s��J�iɅO>�m��'5\f�����$���-��sL� H��pY������!��w^��'����a�þ��)%~��u�R�.��hI��N2���N�s=��!?�c�X��T6`%Ĥ9�c���+�<�p�a��%��=JװE��h��%�,S2���c1r��!������SS�w����L�nSǥ9i��L�m�����y/A���wX�pB�b�Kk;T���s�:G����Q�f��׏	>}�,��o���ֿA�q1�Z����_ܓ�^����]�1Wu.Ƨn��v�����$�o��c<���I$��41f�a�O�O�ݸ�D��BX�:V_����>��}�����B��!��~#�V!�L�x�y��=��JV�|K.�ͽ�+��'"}^�J�*�!�e3�092p*��A�&�T�in(�N���)��v��p-�k��y��G�e�[�_ �1Bz)W�:�\+
�z�Ɥ�t*��8NFF5=,�҇e���o���Md���c7I�s���2���V{8�{�g��)�w�k����fFD&�(MdD�j׫�Y7�����X�js�^n�5oY�F2\D6f�@��wiCͲΰ����R%YS�<��R� ����l�A���e��/K3L ���7��^��	�O��4AW�K����|%	~D��"������P�,`X�^�dE�7�J�1�a_�x�~���}�"��WUbt�^�i�ـ����)�2ѼYy�$�%(x�A�<�C5?i�Y2w��$��/7t[��Pjzԏ����KF>wY���p���a �ţZ�.;yY��-z>אv��KK�GO�:Nr�Y��&fb�j���j��y�^#W���T��]�������U�����Z�F+{;�!w�r��H:�%��kv��4������ڿh�EXr\|OS��$��N�z�>(�e��s��S�뭙Q�M��`\���<P,6���Q^�r����hx��0S�0,=i���.�(٤���!wh��cK`+R\Ho�O��c���h�o�,��<W�"	�T��Ǐ,D~b\�z��6�b���M�v��1�K�
�+�R���H��o ��Lʟ��f��8z�T��3�@d����Ny�7��< )_�%��O7`U���k�N�6+�hc�\eɽ<����)�G|_sw��N˾zB����e�.��!MV��=*z2�%�-�{<GׄI�H�+�e=��U��3�{P��W	`VDE�uD����3Cw�a�[�>RQ�K2���]l6e����mz�;������;��}ksw�ʀ7qF%��3��만R�'�Z	g9�$��� (�7{���d[49`�T�����zJᜒF���;lP��;$�w�����\��2	`��%X�k`�m85v�ըצ��h�����s�YZ68+���p1�z�X-ގ��e�ժ~�&�&TZ]Y�HQ��0=yjqq?l���1OEF35�B��?���(^�;����<�7�yS���K���0� %y�o{�C���@c��ۻ�4��A�=�%Z���E���[�����;�U��j-x��W�*3��p�l�.�4N9Y�Β���7C�ʒh2^[3�����֮�W=�ⷾ_^����C.����-�W�8��*;��@�UʟM �sJϬ�
��3�=���#s|N>�Щ���k|HŠ����#B=A�!ų�����O�3�4���[���G���Z})���[Ҩ\]h�{?�r�s��4�"D�l��J��{��_3��#���� '����:�O�z�0j��˳k2co��*ʔ�<<��O!�n�����{O0�U�\[(awHה@�UO���)��>����Ãcd�
��K^�i�8�,=xÊ��#��cI��a���`U��{��z�'��t2ʂ��(���~B������;�7�+,č�;N7���}�
�)9e���s���n�)9�vֹP����Q�7b�$<8��%�B���Ɗ\�t�X�$$v{� B��^D��j�$�\��>�����'�Z��Oı(&�X>.�c��CҝW��r:z��V�Bu�h����_���Q�0��Rr
��CJ�K��T��H�w����?���W�6yqô���8�6�����b	B�R��5?��������e̥yEfvq�U�LK���䶴@1�����J4�� 򇱴Q�O�B1�3,8�K��,wͬ��
_�>�i�Ӽ�m�O�]��}�%f���w�WeC7\#�����7��7�A+V@��������,{5��6���`���ݻ���hY�|����\t.ډ7��0&��Nu��t�wws�x�-Ay��S���W��ۿ�/p
��!m%0F�J��J~���%%��\'l3o�-�76٠�;FC~O��Ι
�c�ұgZ���a�3�P������w�1K��H�� s$�aS�7p?D��;+ȫ�v��x���� v�}�g՝v���Њ�#o�+f�p���c��a�b�U��00��kOϦ�#4k}����L��W��v�w�����G|���*�6����[;�)B�\�����ж��.i��Bՙt!�.����-c�!��e�N�fL�s�ݮ�@F��T�z��S�מ�L���Ȱ��ݤպ*或m���T��ĕ�g��)�h�QU
�w�:�<�(�	��g��@�RṄ�O�G�p�.̻��3gR)���Q���z��+��Q���u.�(dNu���D�{�-i2�p.��-:#�-~l@����٘=4�����R���X�Wjp�U'��a����H��ݘ"x-u/���W��8����p��
���Râr��LA2e�	iuw��zRN�8^q>�x���ZUh�����^����I��=a6�V���|��-�e�MC�\L����]���2uW�0=�h��5U�U��rΞ�(I�<���m\[#�%~�)�	���{���5Ofxq�a-��l��K)��{�OK��#U_Y#��OUD��[B>m���~*�9�4��O>:���v�ngE��,S-7M�z�9p5�w_e��x^�x��
�abL���%��Jf�F�"r��}e��A�#aH*��7�~�:����@ml���`�Q�5�ĹƉ\����s&{e��g�oky�Z�����C|ن&�h|.��4�X��H����9�۾���$&i7iN��$X/�o���.u��t�v+����N�\�YG*���S��y��g����>8�zAJ��P����	��f��i<uc�����%Ep� L���Ũ #��w�`�@���M��������]�ԡ�V3��N��Ρ&����~�s�۫j*b3,#�Ht�T���y�5���6��R��+`����
���p:K��$���O5��k��J�JFh:��8�:�0`�����((KL�7�ċgF�3yp ,�%�?���Qӱ
���
���ua����%t-����ĥW��jV��ۥ;��>�v#�6Tw0c�^�q���N��q*g�u[�f�5��>}(���v	��ۊ��YF����ҕv8:����z�)�2�ۍ9�������	{�uP�P'��g.�`��Q�L�f�z>��$�������k�v4e�A{ȶ֞�xt�:�V ~C� ~�O鹢��|���=���θ���W�����PE%�aD�����M��wo�ʋ~��������8�fY���Nm� 4l�碙�ܾ�&�1HƳ�.`^ö������Q���	��������o���?ε<i8�=�[�7�/g�FP�Q<s��)<�gz�]
��[bN����U����f]O���+��WEљ�/���1�y������;5e�����fN+��h�RFZ��������#������楼��L��.�N�w�<��?�`0�-�(� ���:k��k�����̝�J5ks� ��<�t3�}q�����_��UX��)?�q%�"�:���'/z�=eg�8�C��;��V�"IR��=i)�����2PQI��N�!����dڢK��wE̺A�������96j�"IK���%ȸP���s�� JD��Vk%? �+��j"�����!̈��
�sP{��F~��Fo8�&q�Z����d$�t�jlލ��bⒼY�!���`8-"#H2�?4>Dyr����q��(>�-�z�v�(�"��Eחph�U�mKY>�D�t������`�6�7��sX=w���M�˽x�7�eK:y=�K�^+��m�z��A����`����	x�Wo�Ը��V0�� �h�'�������d�2ѓ�́��h<�}I[pn�s�ʫ5m�h�_FJ�� <3�A�G4�p�p(6F
��D�Un�����5��Y�������7�.�<wЏ�^lR�=@K%��_��ր�X���r�G�%�ǺČ��B�ؿ���U�����B`'�'+�<��ӎ�]�@�ߛ�+�#S^���t�^\�ݣ^�1U��@�n�MTm����FA<�J[�B�8��"Ns��(), B	��Om���Ѧ��n�b4���������r�%R8������ҥ��k�sT���������E��_�"�Ve�q� Ju~�:1��be{VՏ~�Nkᔧ �AKši�T1������?�?~0Wrl}�E��Ϝ��Ȫp�03�?��0~¶��O'|�h�t�m�^,��<���m?w�3��=[�ĥ���M5�|X Gy��l�J�{�M���ĭ��?A0j�s�o��kFeQa�չ�ȗ�Čk�Do�zU��Z������oPn���~�-AQ�d`�������ݲ&Q�c��W����2=&M签3�k���Ahɥ+@��S7M�h�����*�;J �i��M/��MR
am�J���^�ڑ����W�(d( �'*Z��3D���)e4��^߻&j�\ϋiqT��;W���P��`�bw8.;�5ŝ��$�p?V\�YH,$1[��/��j=1�ʱ�R�Y�b�"_L������Q8r�����C��b��ge�iX�;�Q؋ mv ޛ�cO-����{��ey;�C��.���#���ަ9��%m�$Ղ]z���ݘ��쐃�T ���C�~�"[9_)�F-���S7"
�+���42XlB�j�"��%�S�C�w�94�	��Y�a��bF`�R.�������qD-.9mջ��xF��Q��������+ ��A�0�T5
�?�ye�Π���`G��X0
�JD��IW�ҡ����v��<�G6�����}|���D}z�謙TX"�z��1���K�ykC�m����{�N�A=�2V�oȀ��_"��.�G����sb�:)2`E��[Cg<Ɵ�a�v7y�U3�Q�*g�'5Tw[��OH=�P*�Ӱ ��qq��~:p�Aq�EN0k�ޫ�˸\8y�Fl��.f��Y��U;���ǜ)�3Bs��܄��Mk ���v{��>]�?�n*9Ҭl �s�m�Bд��O~�RJ��r��pG�p����|Uа?�V?��De�	$?�Ւdh_c���F\�h;	_~���e��e���S�ܘa0��I�4$�V?q���G���Z�BBi�Tt2YВ{Qެ)g�\���>������ԑ��U]fp/Pˬ�:�MDUw)�I��y��7_�/,g`��;e�*��0>O�\<�w�s|_���O��@�f��7|5��J�ڨ��A��a�>�s7�xA�D�*��U G^��f��e֤�Qy�4�_� �e��K�_}�DsS�k�����!u�@�U���+o/�@�tG����&���n�!���ܲ�S8$Z3�يY�^�u4��]O$2�(����z �a�!��Y|}����c��Ğ��c<[`M�N�7qsr����E!��>�ҏ$��"�ҟɐ����,M�!�W0�q.�r:	�S�N
������51��\�O�����_���)�HE�vg��T�=_j��i�	 #���NM �	�3	Q�+��6W){ȸ�f��O�}���z�R�dq�J�2¬`?��}�힆p�r-�C�w���U�.mŪm	,�We�n�}��d���S�HCOAC�'TQ��
)�������UJg/f�Ph�v��X�#����8f�rP�\���ў��Ֆ�ܧ���w��%��HVg�[ G���p���f[��/61��d���↽��hut��H�/�6��܉C.��è�}B���#4(�鐕� T����A��c��GtI`~&�j�����$GU��u�bb_(�!�^>I����$�-�����]��7�hM)������d6<�B�G��6D�U��SdX1(�e
�j�PEyLsM�K��4 ;!�����Ȕ������}�ܼ_H�$G�I�kO2%�2���D�Z}J��M�{Y�)�%*��N�x�H�=�d�<Fd�OG��}g�o�3�r��+�N��V	~���jQ��)t��"l�[�b�4��q��&�:&���d��>P�I�˫��U��� غC򰲡7��oD��x�r�[��t�������n�n�x�����Yfa�s���hD֡�\��-p!�~��	ͧe9��W�΁��ʰ2h2���5�
�)'��˒*�s��)���;��1�H-4�����*_5�b.�q�I�9��vE�>�ҹ�(��d̿{���]������6��>~�8����E,_�b����8�S�����ñ Ωo*g��T�2��h���I��ɩ�d5���b#�J�{���q>g!�1`>� ��]g�H+��t"L�/�>�ud��څ�ܶF�w�OiB^!$l�)��� �����/F�}���U��ϝ.H���R��1y�5�[����U,#|���qU���.o̖�ܐ�M�N��M�ti�F`&pn���kʍ��rv���^�)�[�؁���9�v�]̓.D��Y߃%��4c��,�7��v����KWo�������e��U?�>� ��-$�ф���M���x��,ༀ�Fo%xR�د�r�f���Q�w���$�%��];��_p��~�5�)�l�ڷ4gV"w�t��2d��(l	g@������I���܂0�U�N�­�k�/S0���ھڬ��ŬLE-!�5X*DP&�dTD=-e�ɦz�pO��X:�v����2������m`�k������	��K�(�/��o�k�|��if�7��J�FC��"e��V���R$�
"��; $)r1�k���d���/{��	�o�{ڵR��o�G�v����#���N5c�vh��w?l���o�)a&�=�#��x��"H}���J����hܪ���U�M�Y��Q(�9-��`f��{�2t-��V�x��TIoS���4]�f(*���&�[_�3����볪@(��P�-��6���t�x0�>9�5\[�a����P�?��ӰRY��qhL�6���sG�/�`�cf�.�{�y�NssNF�U{G�HY:j�|��&��0٤=W1�x�`�I�,ȫS\,���r)�����B���R�cu+����9y����<q�Wە��4Uh�o��Sl�V������;���8���H\{�"X
� %wx���M�����_=(i�e3%�2���d�/yq^$JS��	RT�I({��(k����,4ȉ{+E7����r�}"<(�:�6Z�.aE�Cȓ@0�޳�oF+pe�D3
\V��d7��v�gG����6f�������1hǗ�Z�a85�P��N�Ӂa��R)���fK#��@��1!<Nh)�`�������A�(5� �K�h<R:�{#.���޽�F"��R�3��(�����kl�������%�Yk����+�{�ev'��?�Bk]|h؛��v���u�,��}�b���Ho.�,���Sz^���(w~a7��B>��@�/O�!`ɉC�C�CV�����;��v$�9�G�h������e�,?Mpl��.��Q6,��z[����8�a� �j�Ƽ<@1�4	��3��؉�2��u;[}����,H9!�@7.
E˲oU˴�(�y�K�"7[9��G
�0f��*���}��e�!XH�vpr��2|�e)�uF}�y+; )���&i�Aua�+�}?�5�%�4&o_b��dCTJ��>���-���/ �Ul�Ps��q���SH1�_d[Ax��5C@���rc�ymq۲Qq��ZGq�@�6PZ緪��9��"9Hz5*���r�L����
�K*Z�-?s��BE�ݍ��M��F�h�TΤ����X�E�z@���N�>f��:nttOA�eT�Ms �9p&pQ� �#���M�ϲ���1�X��K<��3����+PU􇼠��t��u�B0�\�%�!��Vp1"��*��EÇ�V�,� I��9�Y�w������o��0�[	�MHЈY��]!n��e4�g�b���Nn?�c��
>x�y��;�����$4�Z<"?M�=	F �txԛ}Cc���ã^�C�U�3�t�qq��C�[�Q0�y��)H���k'^yv�5)07#�f�!L���g^���2q�ɇ���Կ��8Z_��F�D�m�d����#9d�@ ���Et�!@�Ĝ��<s�>���cL�z?��NROp[��]2DlI	�����۸c�oG�=�j�k9x���;�t|���@�7�ާ�B4�a���5��k*O"VV��N���ʞH@�G2H�x��c����Nڭ��5�\^�i�Wك�ފ��HWW����X�)�= �G��뜼I�.�X��:���t���_=V��%����(7���H匧l!K˸�q���z@Kz��x���Kg�Yb?$"�Z^�f'�56C�=�I+�$��E��f�����G����B�W�҄G���J�ƽ��U��^su��|$�ݰ*&)_��*��L{��"�u���dGa��:N�	7�*���*Ͳr��8RS�w_u��~�*>li<���^�mߌF�T�/:J����x|0Ė����U`<q43�߆��;Pv~�b�=�r�g/Q�ǆD]ͦ3�_��f�z�C�p���s$j%����5��l�l�y��ñ��x/���\bk�8׫j���R3�iZ+3+�����:��!o�:���%s�����˵/w����N�����g�r�-Ҋ��K8E' � �d��Ș�E�Sl��èA���:�㋟�a��&��(����t�����~���V���	x�K���7Σ7U�U��`⫣%�Y.��#��w�g%Z� pS��0�U7�����V�"YE�j��Nk�"f��N���F��ي�O≥Ἒg(J0� &�W�a������8"��������͐��I����o�P0V��2_0{�~(A��v$&Bܑ�s���A��&��Nl�H�����М.���x�fe�#�X��t�����T��<$k�{E�� $������8O�4E����琏�<'H1���c�$s(G��U$`E�y�j9�&2�r����IF�,�\^�f\��n�*��d�x�M|oڋ�1�M�H�����[�'I�X&���n���ȍwҖ���/d'��>-��ev�;h�L)E�I��91���ߪ�c��ُ�Oo�����{����y���֐�Aa�{���3���қ�x3 P��9������n���k}s�˖SK�0��}��_�=ƭ�DCh��O�Շ�
�E�
���������`��S�nI|<�w���Cr[A5��PD���S�d���ï3���a��b��s��.����M��R�oX�,P����ڻy.�8�֍q���~�/�
�̥��-̈́�ڦPi���َ̥z��N�kz|���h������9�W|�n�$���t��ַ΅���,M���m��'xl��+]L�/���㿞�nMA�&IT���i��� %u�$9R���B9�gj��bc^�K[��"��X���x9�(���ķ���fk��"�w�z⧣]�+�B�\�"q�O��ሗg��ߣa����N&�~��Pg\�e7�k���w��8�����-T��U����("�ˁG��<A��v��k��	�J�wNt�9�f�#��f��ۆ9����O�{n��0��m��v�H����dW����g5%�'� ��(i�h�]�F~��R�pDس�L&aZH�z�|P��U�Y��B"�����l��0Ĥٶ�?)��!�,JO}��z	� �id�$/���2؇�/��[m���G����������)�^drڢ�/h��A�r6�vewh��SO[l����tv���Ӗ�l"Q0	�/У&���ԋlt�W\߷b��$�K���A~�z��c��Jy���d����D�f;�\�M��鸫Z�mG٠�c��.Ns&���2�O0o�v�/�ϝ�!��J�(����i��6H|��&�ej��Q|�ރ�م�Dw��Վ�	��atV<p���(��tc2fỦ�)������Rc��,���ٌ�5%#�e݉�Z�%j�-�	��¸�G�I��*_-ZbtrC����Lx�JO"���N'~��G�P��7��>��P��\7���F��>��gD�Z���e0$��o�h��rƑ�M�,�iQ��{��ĥ9�q�D�X���K9�_
9;��P�mbr/�坂1�F��	�Юb�5_�H�6"�؃K��S�~����z �k�� �Aeq.��U|��a����n��W�ރ_�<��"�M[<@�h%1
��W(%�3����]���-+F#�L8�2�����M{��_��q<�I�ރ���������J�Gf!u" 2�����=���nc�Ff�U��[�_��XƕuE{Yqr
�\d�H��� ̿g���l�
{�w�E��!�@`���n�ׅ�L�}�l5�w���Xe&x$'�.�~�P6���{���־�=
����wg�w�/W��=�푃�Lp2|Ki���f2{>��@'�jȰ�B?��*�bv��5`�+]��Ll�T���x�;~�g�B��>c�ݮ�v�S2����E�	����U(�3�:`$��1/7�(A%��pA���P��!�v�j�`�v���mQ�2�@���٘�o"��	�r$�����tn>+J|ޱ���C{���r����m��h���G3s~#��:{5v�%���ܗ)[$�?��:�����;� YK���^9y����K��[z�