��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��秤��sy�/�F�5�
7X9�W�,�e��9�0tgX��M�ᰞlt��e�������$W��̑Ԑ�������xGQ���I���O�i\S�o��"�8�G8Ë��l�ܑ�M�vX|5.�ԇ�s��/���(�&pۗ�Ha���p�{p/��??�\�0�g��/�#� �d�{8;;��2����G�p)�I�Cٗ�6 wb� ��t��{7��)�H�{����4?$�-���g����;�t���]�V�wW���\����A�.K��Q9_9;(X�5�k�hx��U�T��-qP�3\��|y_���`�.=t���lۍ������������(���-���`�@�)��{~Wzfn��&�������SQ�P��#�51�s]iuДKWGw��!���o�RA\K�&�ǽ��͋�tXLc*�7q�Cr������ɢꎍ��\!ж�0������Y�� ���WI���B/JԆmq�)=�t	�k8\Q�I����i@��q�+A��$�m����3Q�i�w�ѩ�o�9��o�����҈��q!�Ha����~2 �}��R��,���,��� w�(��]�/	v�8WN�T�4�F5��7�&�r����oЄSr��4nR<O_n#R��|P�<�i�o/�~�eg�0*N ,��I�Wc���'�w�1BL.��i4Zk��b�84`R�5���f�7՗���p���4�n�dڂ�#�4���dbe蠳w�h(��pk�B�}�Å��7Q��e�e��k˅5�m d����=���,r�������˱�q��ֳ"�Fw.�Gn�2�<-]��k"�I�oys�xTj��h)��{�oE�aaoLg�>��x���i�r���+�!��T�2{Ҝ�.m��#���^:�Y�|H���H���i^�/Mܤ�Y��y���������;��lV��&V^:�̰���\�����i	�Zf�˖�+)ń����A�5WgB�`��L��B�cg��X"�o[O��}Q����[E��T�'�|������̑GCK�֎�@+
�}�Y��pJ��TU͙�he�KJ��NL4K�鸰�@�_��jWYxmΔ�=�h�
�>��.���lȰ1�L�expʚZ���ry?�k�����P8��`Q�`�a��F��K�PC�W��(�H3� �2�e�[�ja�
pB�;c�"A�'}V����*����:s啫���rO#��>y��lXj��n�%>4F�>�T%ߡ���n���
�����qFe�搅����xC�882cM��r����2i='���8�]�w�����C�̐Y=q�	e$�����ڍ�<��32�Η�$��(dJU�".%2�_��SҸ�N�Zz3��H��1�sՈ@�f%�	����W-���9��"�g���Â�d�Uʊ3�~�����o�nU�p/X?%ݞ5�e(�������m��/�^���Ј"�y2��"�9h�3���y�m+�ȯ��-��۝1����{c������ܑ}n>p��.
�����`��-m���!LJ�Vcc�InƁ�c�7ġ����t���L��B��`ՍE;3��s9�L�I��솵~t}-&�֠�X~Y7����F�@�_F2�����o%
���;��v}���cC�4B��߯���R��z��`'�_��u�_���-��_] M��ۋ�YE�w��Ə ?�jd���G�	��wZ��ֺ�ƫ3�E����shTv8ʁ�^�z=B�;���o����m#ur���4�!ۧ�,G�g4X�.5KϺ�M��F} Ƶ��Ͷ�c0�%>RP��?�hGx��2���@�J#zЃ4y�c�as��;�i�8�}���2���%5;2jn�8c!ͣ�Ưn�4
����F)b����?5_6�m`Z����S�ՈA���/�8ڐ|�˽���b�j��V���p�'?zf��6�Z��� �
�`�xaxj)O��F���$�A�Z��1���I�fp���G5���%�B����L�f,�GOu�������I =���1p�Pt@%G��(�`5��*�eg��o3���B��C�&O�Se-�͉���,t�b�?-ȳ�yp�Y\�tt?�>��8��ĸ7��~�5)s/`b���j����JI�/���KO7s�L"U���Vꀼh��7G2��xc�|/U��:
���+tA����~vٖ�Pn�8�K���D������M7�M��d·JO�^�;�{bS�T_.
.��݇h�m1�ֈ5�����.�J��:tV̟�\_yd��+�S��n�׭����V��FW� ��&wzO@��6gdz>f}}ν�Ѻ�,��숡�Ad����b��z!���ܭHJ���K?n���E�
��8��WI몜�&�'�sk��b�/د�8jk�@(�J�u;�k�A(�m���m��E��N]��t]��4�O�lR��(CwD��׿Q�b�����!���7��n9���eW7� �qeO�6�Q���I�����>��6�ph��Zv�;^	�B��H�2�C3-���G�+ȹUZ�
t��|+�9Z���yR��
*��\13�h.N����=D����0f�(��6?Z*��DS��k��=~��`^�언���}�.��uǇ�"�rz��o�B�S�s���0!��p�c�;��Y;y��\%�aq�"�W�Χð���tĜr�ƀRo|&�ֺJ��6j�[���~a��.���� \���n��ٞS�<�Y
��y��8�e�2��	J�C�NM�*\`x�F\�F�� ����ґK��JCBH�2m�\���F�qI��4_��]-�~�;�U�)���_&?���IY��BA��@W�w�1۞�m<f�gU�):&$��?��R
�ڛ,2��I��s��p�oȟ1 �C��b��9IҜt�>�]�S�� Ti�y~f���C���d�*�~P�X����D��,!����]�W��85�5mH�bT�W��Gxr����ɷM����e��^��Ǯ=�������!5a�A�y���f�����P�nv�n��ojᵿ��=ҫ |S3r�:.x7D��=�ϕV?罼�9uo�h����2�ض}LO��=��1��9Hӏ�˽^P��`d9͞%ܹǷ]���|�Щ�Ա�ۈ
�ӕ+�G�F�١ ��|��
�"�2�˖M�#�S�"nE:���vX�~��ef[`��-��y͈�"i��&�����o6�Ġ&r�ҏo,1��!���u ˚+`vASh�n�ڎ�jg�}d��r��X���1��-�}Oh�l������[����+�6�țR{8��#A�6M��GP9���+���O#�%�^d�+�Y[A����� P���D�ܦ� �,!"�W���Շ���Ʌ2Kh���{���y'�q^́�Y3u�}��{)k���%����;혉A���c�7�����Ajv����� 4�;g$��L��k[*�q�A�(��S0p�_�G!� ߱���O8�D'�����{񛪄l
���#=�R	8U�����9��oBzL@ �l�>���#6M��E���R}�Y�B���>΄�z|5
��د�ڼ�io�_��#���aH݄Q8F��y5]�	N�J8r��*nH��SMu�J�G�F�/Qf@�"4���@�Ow��9������3�Zv3k8�Ͻ��Jn(A�^UV�`� t�9Ch��Y�o�K��{N���[
�X��5+`�?'\I ��>](��P��� ���T�3�ޞñʜ��M��d^.�������g�(w�t�(ʎ��Xp�s�S5u�ZL��ځ��&*p�E�N*U>��M�bQ"�A$�f<Qcl~3�� 	������E�7A��x���*EB���䰜B�,�[��l�11twT#w���w�e;��5�TC*�Ő���ϼ6b
��Z�������ԖX�)�*ݪ[�5�&�pά6C��؜_0�T�ӱ��L|[��S:f��������<oeI�u!fiXO,T�-CQ �}���5���f6��������y"S�~�����;����I��ɞw�8�O���(���%2�	���dC���������R�`���
`�뎍�<�?q�k�,��&Ɗ��dؓ�F�e@�$>�����z�ʙs`��X���\���_��۬�B�P�k�s�T�oo̜�K�n�s2��ɬ����ndNr 4�H�D�=��I��8��!~(OnA���~w�U���"ZQ��Wn$[��A�] [���Zʭ���-@��0ΛMch�I��J�<|֤a,�EE��Yvɠ��%G�#U��yk�����|^�/�흆h��}i8��;ߒ�}!�/��^!	��G��|�*��0v��L���1�ܟI�l�:/ú�#P8�N��W���+���%�%��ŨD�LAL�;(�/*f .�W�e�BQ�����L5�G�՚=��Gx�2`�3�J�W5��8����x�l��"�w�O��&�չ�h���;9KJP#�&J��&�	�m�Ko0��ދA�j}GB?	$���!����]�3��X��H�̥އs�����zh9��8�]s�:������s����C�6#��ZM&����M���V��^5	��W�Ռ�Z7SIDt���/m0	9>.����B9����~�� ��+8q�OrDՑ	�GR�@�q:�����/b��i!�;���m+ޫw�aJ_@��T��]Gz��߯P���{�R��x;_���=�`:w��/������
Ib%B
�N�Ġ��D���c_�Z{:�5�u���*\i���@��%�z�S���g�
�o���f���\{�_���|�E���<V�[ͥ@+��`��F+[�!"x��4�I[;��"ĳ�����I��z�~0���	\\۱%���ޯ��}�E��_*�������g��1���%���惴�,�"��^��|4�)=�ڂ[��)�n��@������GɕN�7=ZϽ�R�34�;'�8R���tp�	������J��"��#+��֗�'���9DȢ����E�V�B������6�×Ƨ �8�~�D���F���Ib�W�8����EC�e�X[|i����)桬��z�sRW��w��q�uЛT��"���������]S���$�����-!iD?��]'��ץ�g�#�8�n�[�t�؛)w�C�d3�V=ƼKi��4p{so�n$���q$����6#�Q��U��`��+�@��CFJ  �4-�e�J�܌�}�O��2�as.��n�.�댳N�o�!�~5���6����@B��|�y�-�e݈-�(�j〟��
���ᙆv`�e.���u G����M�	n:��mW��XΌj��rb��k�vD�)-��ъ2�K�~���$Mj�a��PьRF��6Ց�X��S��8���>|�r�	}�������:5�4�H��o��o����.�0����A�`��Id����xV��T}"�cE}�+ˬ2���;s=�\�^�C�e���~-�g���/�c��vC��Y�S�G�;��?�Y���؂�+���]{�:�������EKONBZ���[
�rh�v&vLeE[LҦ�	�b,��,Wf�'ݷ��5�{?
V�Ӷnt����A��t(�e]�Xm�A�sy,zZ�Z*����͔�D�F�\� ��j��7���~V/S���h��R:'�#'�{%E3S��SO)�NTY��E����`��,�	���|�$M+�����a�/��D$j\��ܶ���s���?���>����6|�ʳ~�Q��d�;��?:�8ͥ�I����I���'\���2،�s��AM�(<'
�F8)Y��[�$����xU��'�Q\4�u}_U=z*�� ����9d!�e�RB���
d���pM��_����M�QWˋb³�`�#�y�Hy�����S(M�_gz��uzg�ܗr�߇���$���h��>� d�*g�nPn�R#�X�F�((�k_#�#w�K�;#���tvW����o_�Јʣ��Fy;ڮHΈ9�nY)9A�V.��zJ�K�e��x�B���X���C�Ь0�Ƕ�ǽ3k�(�R
E���7	��E���̈����.��jAđ�ŝ����+�Vb�_OX���o$�?�o�
�$Q��^_1��!�s�%�"cl����IO���/1�p_�q'7^)V�*c;�����J�pL�����KQ���7t�sT��AS]S�Ecq��'˔�B�x8=H�z��U�0/���8#A1��B�D����"xW.�n�wȜvs����s����z^ڲ����j�ʩ��n���pL�d�� x����b9L'�ɵ���湯2��M7����)!���ak��e�r5�J���e�^n7��v? Z�^�+���p L���Q̪�_�8fM2�,����8���{Eng��޹#W����q�TT��8���>soA�/wzL��LB�w7���;:�J���cvQ�u�0$�e�kR���e��Bc�(J8�
5���
�<(�U��v��|�q�����o��,��	q�w�w���q���m/�*�`��#��c��tK�ǡ��]Yc5�ƭ5��G���a�a�<����62<����nƟ�95�1��h8J���l���;��K.��k[A	��k,�������׺���ّ�?څnAŃ	�ue3��UN$;�(:V6iA��� G�]�����;V�J8T�y�I�|��1F��H�n^�T�M��ï�/܃� ��NK?4+zg�J���G�.ڿ�<u q��>p� ��@y��`9e�P�K�)�� "����c˱��j����Aݿ)yEB_+�׍5��<���ˆE�j�.��cc���h"�+��/-tN���݈�{?��I Z�ut��TC��ö���\�����$�1�Մ��-�Z�I��I͋�/�(R� 7j�^W�&�K�F���.�PE����` �.�Ln;T&kv7�:JG2r'!ɵ)L���3��G�T�o�1�8HX�.�K6 ��f�&��iDF�@)ܹ��b�DR��&w��&`��)O�2W�^}�!Kkڒ� ��2+)c�;*�Jv^PC�\��Hʮ��!�ʮ��y	�Z+�_�-��������J�>֛3�4?v;��F�����Iv��0�m�m��6�@�Í�:��ڿܩ#�
�yz���X>.Aޤ�^��O�"���W�{�gO2��Te"l_�dJ5��]��N7Alf-�((s*�kP�����M�gʑ�[����ǩ��G�� �/�k �1K `�tWv狓�{�������.��Ne������j�ms��λ����Nq ����8;G/բ��f�����[^��Ҏ�;�5h����Mqr��AQ�c芞�U���A�����EGӏ�9���YZ�?�5QmJ��[ʄ�{�Ei�{Z���A^w��DSj�/n�7`�]���_D��L@X8�}�Oς:�h�5��Ў��9:�(�Ȉ�{eX@�4ǜ���S��=�<t)���q�l���"��=�&�NQ��Ki�j�#��ۼF�](������s"������ݸ�7�Q��*OZмG�1�a�Wg���G�?3w���i�[S�㏰�Ox,�C+�[8ѯc$c|D.����������Oݲ;�a&�%�jB�Ƹ�"�v��l���v��xIpv�#�w�Y�h���ۦm�N��n�Sp�7�� �)t��z�00|���¹��J�\u�J�Z�b>�n�F綸���t����ʶ�$oe~�ï��O2>wq��(	�	E<�& �I��]"� GZwL��>���qn�p����K92E�\,Vx$�7�*;<'0Pt�Ʊ�۟�?Kxa��:�'�IGNt��ǃ�W��r��޼ C/v���_��5���a�+z�A�+�����(��fsG�/��_ǚ���>)�<�5����q<ǣ�~��G�혭�},�G�Ҡ���e+ �(�:�J6_�8�`)ځ������sl��#҈j0nQ�h3��Ԏ���z��3���f��'�#�"��}{���Θ;ա'\��г��6-��� ���������|�&��̀{�)�T"v��LWۇt1���� y�ÏGCJ�j1���A�!�����c�r���pQ"�����F=��\���i����S�e��P!�� J����İ#R�~���V�p�A�C.�;������+/�4�YZćj{�v�u�3�����툹��'RLҬ�v��8:AL�b+h�@#�Zγc�`��E��j5ݦjv��,d$�Μ*�V�I�}�N�������8)�jH������t=HLX���fўI���F+�E��IT���>���+� �Q$D��ih� �4�� ��������� �`��1J(��90l��ں�Xb�Hl�k/+���z�j� Rm�������.,򞬔�����M0�J��M�����t��G)* ����y'�UA �?n���\~tW�k����KR&<U�=�����V�����5g�͝c�(m"��8�a(i�W�d!L)lƜ{o1�nc��������G��ǌ2�����浪;m����>�V��撂Q�M�m�7��vzd����+�N��TR��vu#rI�d�b7��gHk��Ԉ��$��c3��i��NNj� �XdW��������a�\�J�^� ��k\5��ս��+U&7�� 9�WTC))k�N���6V�I��:mm�X��P���!:q�L�/��y�)G�(�w����ᝒ��
�fRg>O��?*���#��:{����(�7���NW�����a/~�_�|��H�)5z^���G!�H��x������K�a�AZԏE*����6y�=���E��-�Pc�_�n�m@7rHG�T����mt�(
�Q����gk)R%?�.��7�Q�Eʾ~�e�&����t�x4��� �3m��>�I����*Y�������Fc��?!�O(+E�S���*�&&�����`1��C��Zj�sp��_���~g��X��),�G�aGf�����أ���BP�Щ�[�X�&!��g�h�N���DD��s�Y�ϡ_a��W��"�!~W�囹2B���T����7�.��7���$�01��萾x�S�0ٙz�l�LrG�{�=i�τ:�t#ӵs�J��FW�Vf5��4Z#V iS%F^��w��U#�0�[9#���(����;R8�xL�Ǿ���:���۶f�!CC3[��ɏ1�L*��T�qS�Tvz7UM��/k~ƺ�|Hq��4T�p�Y�l�����!���2�)�:	�y#��Ё�������I)i5}&V*(��,_&�l|N_�z?rx���5��3qq2>0��0O��R�-^i$�����x#X�32��&p"V�)"\Z7>�Δ�©�k��մ��_�/���%�� ���0�`p�U�x�n*�ۨ�����fg�xq��Z�sy. *��ؠ��7��uP��/'�Do��K��ф��3l�l0i��KD�����~�o �Y-�����|&�P���Qo�ơc����&����6�GU�iaP� JO?<(J��PZ��8ce�NO�X?�=��Հk=3�(�h>7�LZ�EDh'�$M H�c����pNAC0�Vш������v�IE%w��J���3E���oD�{o�1D�.wcu��W�����0�e��,�i�����`^���S��ӹt@���=~���QK�+�2!C�0V8�{�	ýH,�@���Gf�o��Q��/��	��M�L£��9^����!q���X�
�ϡ��a��:)���b(z�TXZ�k@Z����k5��bz-�i�*_�Q8|�o�yψ:�a�c��(��-�r�rr4�$�VR\�>��|"/IBWFJ�� �7OK����c:���aU���*{�آЦ^�Řs��nth�jV�,�t��*|,��bj�����\����]̠�����A���`޸���=�s�]�x&Y(�.�>eS��6�T��{v������RR�Y�Vj%�6�<73t@�D�I��,ZmR���ςL�r^�Ş��g9�ȿqǖ��ϟ> sFl���7V�<a����+��3��h���0HV,?7C#3���o~����u�pM��]{b�>���N%��aM>����c�M�H����7�l��}%�^��M����50j˼����K�v緀c7�|&��Ҧ��_/�p�}����.�-\)�4#����P���ߩ�-�W��.�m��q�3K%��(��I
�v�v-�18�bWMc퟼�gߧ*r6򨤿JUz��7d��'6�Yݠ�>��Mx~p���E��A[Y:��b��j�/?��~��c�gb�>���*��|��޹�oy#D��@|�Fq�L�r�̫�Gl���%Ȥ�.�hH-U�|c�����A?�#Ҁ���w�(��<�8��Џ�M򾏣�M7B Z䯒1Ǖ�4�����?#%����Æ�Bx���j���!�����ȣSb��R�2�c aa���J9�q�aR����F�+>�r��2O���u}̩̓��9�î�����%��S�p��Ԓ�	k?�������Q�>�o�$�U�ĭ���a��(\��A�'���Q�7|T"s��#��~+�Q���=��bpf_t�� O_Oѵ���++�W�n(�)��	+>S)��w#��e�/�K�w̒�Lsdx� ��I�������2a_#v��U\�{�`G�Sۄ6�'0��kQ����dp���{��->������|��P��Z�m`z��'OF�wq��^��r\�	\�"�ׄ��#\���5���];g1z�HNN�x�� �j񄷤>-,��<���S�� �q>�o�y��������a�X;S`����k����.j9�V���V���F�_�|Ue��΋+P;���#���A��M	��|~�&�ӏA�{�p{�����>L���w���vG�O��O昳�|ĉTJũ���P���d@/��z�A��@pY�v�*��L9c���@�9�)j����q�w��}S��>���,�`\��eҧ��{�K�3���g^��m1����A�7ɬ�Łg�����2)�(t�+L������M��4TV�y�4�K�C�r���?n���2���v�QZ��{+����*�P;9S�:���v����K���Ga�,�k��b'I�}:���1i6z��U��]�T'ߺ�5����5�I/6�1u07CB} :�x%��e��P��몾��_�ulN=�:�:,g��=6xd���>�F�G��;�۶Ɲ�I*��(�&��p&�2����Cy�[���*"�
 �3N�&��tuf*T4�ջ<�_�y�_֜_8l5h�z������<ج�7��F��6%$٨��s-��
�I3�5�:�����~v��թC�|���1;D�EKߘ7Z�n?g��:�uI���d�?�]<kl8F�ϞS�������q%v��x�"�;±&�y�0v|c+z"���A�Ep����f�b�K8���?���L8V�/�G�l���2�Q�&$���]C�Zzހ��x#�������,���-E��#��������'=t��Eپ���<0Ȉ,ya�5$|UWX	�4u3� �_=X�%i�#I2 ��oU5<����Ae]�[�O���UGcz��\%�r��0t�cK�#���u�7�`\��3$1��w��v˯��l��fC���]!��B8�ÓD���/ �WR��_�)Tq�0[���O���\ު�K�� EPևזe���<��s��ݚ~����(��=�^zsFE:�X�R�X��Pr[�yY*Ws����y[�2�]�������#�g	�Z�R�����5��:DB�hI�����^K&WW�0'��d��Tة(�Y��ep�����
�������M��lK{��]����=��X>AO
d-ʴy��ق+�.O�e�%BN�BiS���,�������|Y�����']N��q��l�Q��Rg����A(�t.�<�����Q��� �j��E9`��b�����O�l������h���Ab8�2t���:����Q�l���~Yӿ�u�<QÕ���R����v��w��/u�e.TX��\3h>ǡ��ټ��U֔� bǡ����	T�઄�a�����/\�?j�����TmΣxq,[/�!a���e��h@���š�/S��u2����y�4`,�Ͼ`��vuS!Us ���t�n��
)��
qv�E��ʕP��o�_>��OwԝX��0L�QQ�,?�C�0�%��3���)�?@ǆ��6�SӺڼv���ܷ�����
��{M�p�o��/�p��ev�`u3�������ϥS��0��]�v��㍯b�:�=�WC�R��������Lw8����KlY���I�@\��3����b�L��N�o��"���?D��F��\'䧲�˵��2� ]ƶb=_����T�O���*�w����"�u���_T���}����RC,���dK���[^�,���-(�Ŏ2��c����C�}�����W^��2�Q{�i��٣���3���=�Cw)a�4}1��%&��\�# "m�;�6�ïkT�i�����ʦHb�P=��7��|U�!2�h� JH���P�}�T�%:����� �֖9o`_���+Dw��t�y������ �lA�a����hr�B�R:gF@}s���U��U Qi�s��^�VI�j�d�E�j�G�������#���Ł�����n��S}2�0Y;C��a3�����JNX�������=$�4���d������~d@�tn}$k|](�u���'�����JEl��è<D���M��1��#ڔV\�b��H��"B�̤
Ic>|e~89����+X����ޥ� ��`��_��2 yZ�L�R53EM=NN��?�T[\b@d ~����Q���8Z��H���3s:^y�4��?`����4��QUl��
�ᰣ#��O@�s>��q2:*�9.�;�q!�Q��ݢ����fQ"DTO�,$ ��u�j�T������(^9)M:���p��R;�o����O���%�a���\�Z��FЦ7���.�%�N_,���������R�O�[f��R���
Az�s�����o�.��ݫD<EJ���*"��^g����|F�=qd��i�gb{	^V�ӝ���8�!dZL�e���EV��0<����C-=</6	����i�J��Kw����;h����,�g��ʎDYAֆF@R�.�%�i��y�~&n:˻[���-�̔�Ra=7-����O�!�p��;B&����$ ���U���{37Q�fKI�)��F�&��p��d�᳡�M(�*]��:Wf�ɸ��|hO#U'�$N�'D�� ��P7z��?C ��g�y�c�ϐ;�:keD4
N&�?\S���f�+8X�`�9���ϭ�g��e����ULl�h3ʫ����1C��ؠJ��*[��ɉ��l��8�<�|)jK�}%k/��i�̟���f�eN:�=��H�-;9���*����6,����ǐ�^G/�B��=w��if�y���m��1��?X
E�e��F<��G~)ϓ� �I`@քh���#/��-	�}ғ�.��OG�TC���q���_�D�0��S �[�D�ך�{ݼTu���l���|9s��Y( ��2�g�������߰q%���N�W\��R������O�|]���0\�LLЙ��ͯ���Vנb��
�_8�-ū������V�+=hn��$\�b����	-�Aǽ�n5��4�ӷ?eSgu��/�wG�VYJ�U���(.�=�R�=٧��vd����E��x9h��{9�v�aN6 d��A�^��i�䣧�ܹE3�c���$�R��R�:�mL֞;���0�KJb�(����Z�7M=� ~Z5�P�O��g�1	�U�'5�'/�����
&�sJ>
��ԉ��{�� �Ww)���V�<�#]-u��d�X�ջ
�H��Ԡ���~gQ -��[o��ш�h��}��TAu�C�v\OKg�MG ���\�ۮ*�{ƔO���@#�цsn�a��ih+��eup|�4�$�0vM{��ܠ��f�O=��L�Z�՛�}�F���o��&���E���ZD���5밭��Y*
x�5q��uQU/i~��	vq��`Ex��#(''���Lm��\���R��\z�ts�H����u��A,��#�O���T��!�o� E(w���J��2��$/Mm<?���GRH��� e�x�K���`��8�?-��[,2�CZ��M�����;%���la��W�J.��<틌}�'��/��l��*�+�@��������XG�|2�\�5�~�؉�$���� X��-��H�C��f�G�=3AY<d�CFGf	|[O�u �u
��`S���{�7,Z q V��l�P0V�`$bg�a���n#���Ө����z�Z�:�Dh^ 2�% �8��C7a��"f��vi�T�K� �F�賅��D�>Ww|�4��Lj���W�㕇٫�hJ����j�п����ِ�^��nZ��\��q�c���,ݔse?�i�-Y�k�]���c#��g� Ư!����B)ea5[#�� :�b�,s���R%�(>�����ћ%�;n��
L��8*vH��n��\����g�Ʋ�!�D�oy�ը�d��Crgt�ż��|���F:v�c��������-�4��pΆ%!�|�Y{���8�"�e��`�`��
���QS&]2|����y�sP��o��  ,���TI3�5��#v�S�j��56�"N���sW�X�2>j6J=��A����Y�U@J�1�$���v�߃.=+'�-}D��y6 �I�f�7�LSf4^Ԫ] �?�qkN�����M���]Dp�,��J�����,YW��d����$# ��Q�_&��a���T���45s��j�3-KC\E������H���艊k
>�Th?����д��ּ����VWI>y=b��7�͉���`ez��1���L��/�"�a2a �@��-���u�*�uP�(�����6k�����,��F��c���d������t	����C��7Z��p� ��J��\!bw����
C�\�h�d���o�iI�1}�H4��4�c�A�Ep��U ޱ���L��v=z��[R�!�{^M�م��[k�,_�~���w)/�9�d�\/q�����TA@����?]p���}���«�G8(H�w	��lOS��E�q ��2<��U���f#�E'���C)�U����y4�ļ#%���]���x�84������z:ƭ�c��P!�BO�X���F���^i`J�l�R1a�T�$xchXz����?�8Qr��C{D�ʃsB�t��:���9��~&��@{I�b�g n�,%��e���{�-��_{9����r-�I�}WPU`�f�ҁ���~�&���}*�^��L���?�cJL��#V�������ᇼ�cb�c< m����F�����F�!�*��eL��̾kJ�T�e$ֲ�F�|UR�y�Gj8j��HH�K�3�`y���c��4	=�&�Yzg1+t7(HVڦOX�!�714%^ͭ���X@D�%��
��Ą��!�,CԆ�.����F^����	��;�솳����q.}~w5ʛ��x��$#c��]�o�V�~L���~�[���j|�k\"��3��N9��L+��׫�g6Q���nA-ʣ���;���ڨ7M��(�Ba��#��^�H�-�:<��-6��/��k��<Kc3���O\7w�Z��Y�ƆzfT9oUm�ʸ��_;� Z����F��,�Ϯ�NS���ៗ���������A7�y̜I���0�yg�:��U������V7���E�׭��`M*�h�=.�ʡn�'�{�TUwE9M���C`}\�A�9�����d�:� ���L�����׋5�-	�zE�M4� �w�*V\�v�
vA�5�d=�U��.���� �%H��'���y����C���~��B�oN��E��o�I1o�T�	�C�s����F40\z������-��U-cx:�̖���sy,\�E�B�[V>s�$6A�|'c�S�EH�@��x$��3�e�4e���������Ԏ�F��X���/e�Z_ƿƪs�v{�����q<������(X��I�����2���\3���S�x>�L����GFYQe�&N4x2&#d�Sч�<D~��.x�륷>L���r�dE��b�1�@s�z�÷I�Š���H�(0gZ�z� ���	�zO�+F�F����L�`�X��[+u��b,ݹ^�4Yp�9�άs9!��5�vG���8�{À��6�NbU�
���*����������ݦ_������4�gl�^����]#��9K�=�|~ſ!�b��C�w���u�g��O��r��lo���j#���L	1�5�7?�hΤi��P��^|^��m/�K��i��=�V�m+T�t��U%����c���5�+Ͼ�Q
WHd�4L/\o`��s
����jcA�|�6�f7¸OK��D	�[ ��'@�v}�i�`f���o�f� �2|�(աc'΀J]�� ����}�>33�u�.�?Y)�Uy悅34���0$~;��2�Zh�c^�/�&�%�.��N�'�Y�v=5��/d�y��ꥄ��gw#P�h�]�/�i�iW�a�3b�	0z2yٲ,�(i4�kT�[���N��{=kiwq#�|�_�l�߫��55��Y2/Kb���c#t�U����Ԫ��0�%�����V�ui��$SA:�x�D����쏜%v��|C�[�����(R�����p�V��o5e�{Z��x��w`�N��74!���Q�Z<�|��}ޟ]���������9���ԇ���	1�o��˩���3{M^�Ӕ�+	6g�`Ǒ7�7���{v��х��(�HqWOׯ J��{�J%P#&�����.����V�v��+ȗ��>s�f8wB&p��3�g+߳x�|�S�CW�E�BRr�6����)�A$���^�TB�>���@����.K����>�c�e��_�*���Ʉ���1[�Q����G��l���,���;��G�rg?�u��� �h��e��ZԊ�Tqn����{
���GAt��Z[�`��z@�Ͷ��8�Ǐ&QL�꯽�F�i�wC�$�B��o�g���FG���=C�k��i���٬9�c�f%=�uD�p��́�{l����T8�%�2�@S萩�Շ����@G=��'S2�C��a�A#}�&�U��[�kOR[_�2Sge��/LW��5u۔����,��[F�UJ.�*p��A S/�O�-��^Ԏ0�we���5�J��-�ª6����=ŗ�b_�ֶL�!j�PM%8>�0��a��Ej��,�N�w7�)K�A�'�D.a82g)��nL%3��n.=��"�`��C
y����o�{��z�,�ʂ� ������_��0AҴ�R��E��#dnmm���X%H���.���)���^�mͥ�9��ssA5�Kg�	2R�$�1l?t�+C��)�*&�g[�ms����S}KfM��E�P�TU!�� c�i\�R�M/��e��af3e4���ʊ%���	��e�u����c)R����d��Ɩ���@�('0�5���o��}z�s�H�8��T_�u��Q���"��mU�f��_�Qߺ�:�S2w,H�xv�=����ZT,�yv�dVw?��_�_�����fsk0� iT�[��D��p`�ό]f*?��Y[�W$�g2<����A5��p�ӫ�GP�e|%N���B��u'�U+�)�١��_)�"���I��"j�w�}e�{�f�0~,�:( M�i�8����J>�3B+�dp��OQ���b1�,����ݩ�3G����Q�;��8�
C2R��!�.��V�^�`σ��R�ٞXՌ�Q��h�cZ��Ǜ�	q���K
2f#����'w~��ږV+	�L��^"����tk�uc��� �G��"���T��w�V��s�q��J��[������6ɻ,�__c��~d����X�I�Au�Bs�h瘱RiN�4�ZJw<��2dM�Tި�SsF�j�&�f2jj�f�����i���맷�GS[��a78���xw S�����m{�z�R�����,o_��m}����D�7�aw�=
b�M����Cb�e��Ѷ�0i��;���rn� �u�C�ѽՅL�`�:x�_��
<��	�ʦ���CGS\����{�������/*D�?���~�yiP�56���dC�Ag`���D^δ��"s��I��BX�w�s��U�l�-{#!g*,��R-˲���N��b�QX��T��nZ�#�'�5AO�}�{�h���.����ח��]�8U�V.~@�{��vY���*8�@��P*P����:��'�0sA��Qi�c�#��B�S>p�V�S�A!jR�T�؂N)��+�.m�k����s�n�����T5�.ޖπ�̮�[�z��K�'D�5T!�#�������<GQs�����m[�"Ig����K����
�Q��O���@n?��� 6'�x�Dҕ3p���=E�>U[1Z�m�vs�7AN��~4�s
8�V�A�ɹ�X6CӴ3�u����� w�9��H�J�b=�b*�p�0dF|6�w�a��4VTr�-&����/ס����h�O�0���H��`�{dG�?�!��șg�2��goCg�فcH�{�����B�-f��c��i�ɲ�h>�6���IP��د�=m������ƺ_m;�w�y�m�]�[-!R�F�&��5_�a��CFx��wUN����E�;�fz���ʚ>5��K!{�ʪ�"�	�`2XM��ڔx0ɴe.�I0&�@���y���Z,B��dSG�g����+�?k���}��s{�ͼ�)�84L�[�&�,|r��^����-�mh%Y�K�H�kv']o��a��ǧo�g⸓T��^ɩs�z�$���Z�Ÿ�S���|I=NH��O���O�qZF�����b��i˄1��ڂ@z&!x��>
\�^�|�g��pFU
x�CFT�`���`r��W�\�Ɛ�W�z�e�Ō��ګ}�O��"Q��:�/�R���q|�w�@l��7�MS|gֆ�m����-�����:{8��J9��L�v@Ǉ� �����Z���s'X�m�I>#	�Z�"�5>�f!+{�w����h�,x��1� �����y��P�p6I�fmY(?����\�����	K;��@/�u�aUi�Ž�K�F	'���{�	E�[�K�S����o5<�m�6̫>(����۴��,��Ǘ; wq���8���.�SA���I�t�f��F��h&<-�iY�����RMJ)���^'�_�Ծ�7���U1K2�d�T�α#��*ļv�ᗃ�H��q��3�N���q �٨X
����wb����As4u��JԌ3WU�#'k ,讧�������"+�S����l&�н�h&N�� �;B��Yd��U-��?�D�T�BeO���E,��0
ƕ��s�������Q��lm�f����]�5)�68�v>�.݅`���55�z~�>.?o_�3!���:�w����h'q\�������O[+-�3����!�q��{����
�K�=]_�-�akx����/�i|g.'"���Fp�)%`"�8�Ѷ��U��]�m)(p|�����wo�:,>�5�ݜ�H4Mk�mYɒ�h����cW�b��;[�5G��>�4�'" u�q^h�41���=� hv��g�,���[j�貪�'���m<�)�F@��ƠK�����jBps��S�%堞�s�,dCM�/�3��5#ߐ�m(n!����e�x ϧn,��t�A��\= ���k�F$B[���T��D�>{�k�����H2���|�%��*6(�v5�>������O��F]MRm�H�Ǩ��/l�
nݮDku��Ш$xF�+sǒS�G�X~p&�Htp.�A�]0�YM՚#�*1����;b�����잡�q�YsƼR���<�e]�>~n����p�9w�'��̞G>�И7<n>�9Gދ����+oّ�x�A�`#7�i�E&c�ƷN���d��%��+7!ʧΟ�nFU�뚎���W�D���d��z���K�yWī�}��֋�|��kv���-"+��-IM��R���x�q��Wj�����V��~���|x�w-fa$lU���j_�;M����V����Z������[�ł8@�H���c� ư�Y>��Z-6�In�z���xuo��x #���4K�m��`o��+��@�Z�������D����w��gQ
�⮔I(�0�t�R�C��<����k�2?� �h���7f�f{��ca�ei�,n�vS�	�w�Io7������pT�]&�]����&e�����!4�h�3$�D���Ư*�oTU��-�Q������df<�Ui��u�N�vK�z&w9r:5<P�h�����[�D4�ҭy�����@��<�� ��鐱B�T�C�1�.��@p��Hn��5��b$�q�h�̊_�ި�(Z����CYڦ�YH&�j(��v�XTm�]1�k$!(Y\	"�徽�dո
o)�sP�-7'r}�@��#��46�C4Y?��,�0�$��Ul�^�}�#a
*R����"��ċ�ݳ(�e���t N��p��[����S�3x֏WO�z�
�,�a��{oρ�U��N�s������'����A���$&*��]5�]�ҫ�n>I��aX��"��d���ɢYH������@�8}�/�g�� �(�=e k��[	��n/��T��Oh�Ǭ3�UX�]Ś�Q��i��]3S�iF*<��m�]潚U��%鶹��MiG��L	
�#����@2B�(nv�f���A|k��m�_,�� ���t�c���J^0�@��)/�S����
�h��W�=��4�<h�g�<p��Aa�M�6<�K]�VYd��D�{B�*�X�>:�;�|���j��Y���Wh�%ݝ����j$W�Mv��>}�ڻ��#�(ȶ�Y�Sol� a�7Y� ����
�O3�˾-J�0h��|�B��z��[)l�0-����\��[lF��|L�Z�i��b��9_�=��$�� ��g�eDeM+��Y��q���/(�m�����8�ϥ�URH�Q��I��
竜'L�B>Qu��r,D������N�˲��RK�{4?Dl�k�YN=�o�G߫�dhJe
��1��i��������~�b�������d1'��8�;d��2�EuX`z�1��m�����%��@"՘����NĝX]�{ �򏷩W���Sm��ʋJ0��Hy�cyG.e,E%O�8��; �˖{�˟R�2��X�p�!�=�G���/��Z��s���+ ��=ŵ�a��:$B�EN�X�>�r�ኘ�; XpΜ���ym���+�YĦ�E�J^��bg�@"�>�~֏/�  ԫ/�.������{%k��=�W�Be#+�H��vI���I��/��6�+C�N���8��[�ߒ�]�g+5�3�i�/͕�g��]Q�:�f���L&{�
�����T�z2��aJ�k�w��j �k���D�{�82緌-�IV��)�"D��R��(���3yg�]�����ҵ3��9yδ�?�ݺVְ���ǎ�o�ᕁ�f��r�9f8�?��˻9a���O��A6n�L��FS�F+	
��!�D��\��qb�*�`t�0���(O9WT��0�F%����TjC�8D��]��8Ϛ��|���.�l��{Syg�}��%�qm�,��쬨B�p��5�Λ��(�a�|����	�wA�槽�v��A�2"k��	C�MO.n^D�"�B�v� ��vu/�g�p\�}9�����M�(0�B��Tʱs�9&����WW�9��a�R��{=E����"�Ѽ�~��b�r�Q�޹Z�m�C�u��e���5��`f����{��}?��Z^�'e���rL�/�V���>���Q%Ukٓ�26�!�y����j��
\�m�p�Xw��z;�s�)�`k{CC.��>�/�@Q��>�>r����4��A ��lon�����aZEi@�����Q���W��+�S���ҚX�
�R�<�ˈ
!7[�D�6�G�f�Ngy�i4��Z�����D�5�Y�k�_��d��Jȋ=Ku(/˽~>^B��-����9�az/6��m���%%Xu-&Ї�;V��)4����o���7��z}�G6�"[�a�ـ�z�@}�Y^���G"/X���r�pl_��U��@ůUJ�_ms�h�}�!�	"{�(m_���jrd�1��|�����G���B��pga��[�BDELo����fN��/m}���Ѻ��A��a�W@DiA�%-�s|EU��8�S���M�?���ջ���������o()"�]1J�������]J-W��ɻ2�N�о����[�'qLs�m�[c�ӡ���1�r�ڋ�����N�嫔�]O��C_�R��
�����1
&�%�њw����	\�K�������9�ȧ�굧����k��u��W��/[���Z�����Dة�������7�Q���9f;߻@�劸��Pnn��K��_��ț�������YM���]`�E)��n�� G$ꥵF�DP���a��W� ��?�K
�;^�LQd0۠��7���\��-Kr�����*
�B�:���v�Z������ݽ��ĂJϜ�.��6:����Y S��}�U@L�[�$�A��W�MB�{0�/����n�j����t�����+�S��.e�J�%��Sq�
��[�N��7v·>7tEʁE����@����n �b��	��dl[9I�!/������^)���@4��J�$-��Q�8"��<�VW3��O�-Ȳ��1�F�2�Py^�_��q�����嗁��ET���<ɇ���=�����ΰ_2m� ������cu6�iG���q���"�^����]t�(+%��ٖφ�B*(�][ z�^Gm��K#\#
��"�iW3O ��92��Ykssn*b��5���p`�Û�L�ܖ����2�$4�_�Yq���4�v 7s��� S�}I}�����O�����e��ɡ[T�q�6�����.�E�c��#��\7k޳$�T}~z:�n8�����Arp/+��6���SX��	�����-��{�v=*����ԝ�LG�	�(Β�.Tw1p-�lvC��od���ʆ���㼗�|��9 ��G'��n����`�� ��ԭ-5��k61��X��H��f��(�J���hӭ�� ��@� �g̓/6�Xq����g����v�繩��[�p�U����ٟ�vL�\��P �������y�c���\��{��z�%�\[=�;�CR"����u`RmJ�Ǭ��&�c��g�"'��㥀X v�����Cơ�:AFӊ��-d>�U/y�4){/K��N�3���ؖ����G�J$��j��`D#%�~L���~��yZ�b+� �_�2��0�S4�'���α�<#�n1I4ke1%�z d�Q;�-�ő�&V���QT���,-
O^l��j�Q�q+^�S ���
������J%sT^�7`�Mbj��8ٛO���5�b}��|�yϛ��ҕ���3�C��2�R �46
�^X���o���WZ���ܡm�`����Ȁ&�1Qv:*t]��p�J���n�w~����u�7���D��m����	\���a!Wć�E#*��P��Jv?�`���$��jЗ��-Z���h�8h�Ib�Az$�/���X�:L��B�:O��$�c+�/��yn�uu���|_t8Y��#pT�����K�c�}��8>tM���C{7�[�{-���a�3v]��;��~&:���K�4Ӥ�5^΅�;�F�?�n���#��8ï�����56*�.��>Y~`-�x�T��*tNP�����`>uo����];Ց����:���"�I?� �%��.�EK��������΋rH��u���iϽ��4�'jv�a{��~�"S"����F���;ss�@;>G�)�oSʂ��B�Y�p�o�
����������\<�l��I_���]k��O,D��g�eP!��7<F�H�-��˾[:��867\u`٬19�E1#V���9�O0�b�F#��&�4,p����K{Rmp����ɋS��4��!����Jo� =:��yg��G�������y�d��/�Z�65qL"m�q�)� ��K�<97Q�1��~7���1�g|��f��`�(�� �)�r�sӼ�$Y����W0�mHFM�8B )R��Β"U3�1	]�,������JKH� �+��(�����7�O1T#O��Y� Y$���Џ��[a�n]H��'ZKPB5�j���6�������*+��:�Q��/:&7����n�,�%�R�<[~�pU�	�R�;דy�K���\����ٳ�k����C��m��pT"c*�!kc�1�l0t8]�-����}��+�{�]1jְ�d	����c/E�ؿ���U�v�~����e��Xa���T�=�F3��ͷ���͚y&�g��1���c]��,yН)?� 
��/�8k���Ҭe��AZn�U����1��h�J�[��޻[c���VL�HI��_��S)�e����v���G�7�
����ѻ���V�{ۥ2u�o�����[B��'T��((0��}e/3�"W���_q�`�3x�b�&lv[�k Ħ7%��y�p���T$�u���[S9�2)�=4&I��:�!���i�"^�C��9�����k�	1ibؽ��\Z䶗MI����h�@I����4xɶe����(�8���H/֒�H����~�!|w܀,?�GO7�Oy�e���7��/sk�0�ľLzC���	�4���S��TӤ�E�\~}ݼE���`����:��D��p�iv(�˰���
WeF氕q
2=+���]МF]-��w錶�77�c�/����gK�A���6�%�_����]D����/����؀o�>=�k0�����kt<j<��m�9�ܧ�v6���*�ᢇN��Ê�>����wh&3:Al��Q����zq���wɡ�Y���Qy;�O&,��<��yn���ZUi�Û�!���-n[h�����A��op�@b����P���q�����h��Ń`��@g�eR��$���'E�Df�qaiU�N.�l�w5�o��S;'>t�C�ͻt���wAZu��/�p@+���ET2��:PN� ���LEh�-oФ��[w[L�:����f��8��� .�;*�v;�	!�
����k�S�}aT�&��=@��A^QBW���SWس��W��
Ȏ��X�dS~h7vd%2�(�
�,Д`t�R0�p1�R�c9(�1f�`��FI4U�{o!�Ke���9��߉��"�9SA&d�񵍺k�ϣ#O��'� � �P��T��P:�+w�1W���O�q��Ů�^PU־�R�� ��ͥ�![�M� �1�|����Ԛ��9Gv�z�:XkV����l��z�8b}f��Esa|�VТ3�e�Êp�G�W��9�!Ɣ�h��#�Nz�D^
��Z��-��ͅ�� ���0��ɋX����b�X�