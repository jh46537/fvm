// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CNN70lIrnJmSwmjRy5Rwbl2qZQgsabsAcxAqUPplfk/2yI3DmiIDvMN9JPcurhw9
PSqhkhKECPOyWrkJ0Hvt1u18N8U2QRfvI6L5+9xufQBhBtNcgx6TtiOR/fNuQcCE
QmtwxFE+bRCj6iM8KAxdXjazMNAzQ24ZQj92d4rcgs4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 196112)
xP2ewCgFQSPWyA0smOa3OZHTaBpI2RXMs3vohGL7m4QzLt72c/XhM7yc1zec74B8
8AfkEQw3Nv+97GDwn+3qZm911BxxARLYsksRnnYgPuxt2QnNa5BmMpfQnJBlWqQL
MtCYpJgcIsNmxaw3fGcf8Pi21rPPjdImuqnhYFminKyEN7pH/NDOVq4dSi1RMxxF
53sXzhAAr15rRcMEsfQBU52H7rke2hukULODrjXcdsmHSLW7/YCagm6al7ZGWhFl
JFRdgzqPIBQNMj4Rs7RnL1BGEO48CyQ22nV5bkQ5MmyMODUuZttXJsiFH2qabNqF
T1gCaH/WoMQ/kE2hMZXEgbBRaHaEqq0ttJjfmI/iFwuyW5QkfDnjqk32+hlRFYYw
PHCtZ3kJo65WHsTzPps9N0ca+h4Q51qAM7yyeOi3TXgoy3YsiZc+0NzDLoGNBZDc
IpIDybjKqr7+pF27owqAZxTYRnpoBaBwf6Rt06O0VY4GoqL7yy4clgnjYMwwKEgX
iINaBIRjNNoUJ5AdC/DYqgLiO4mispknx7/N7uHhYF4VSdxIYPavONNuiDJKYtMB
z723YHI+rTHOHdnIYQSs4f8JxJtdU9nbKZpYKYVKyjSc/osdXZT6eR/tUXxwreNo
7CZcHYAcX85DtwQz6i8Hs8QcODlhQqsxcH/lFhIjKCtsJbw3BbE5wM5V2aW+J6cC
Wm5hXzCrHhpPf+pdm+oKblFLKsavQAhH3Ptyh6GhqC+u9pDp061AXebfpoyxMysd
fQQFIXg7vfpai6vTy7E1S+xc+u4dCUV/s188WixBx6iG87zyVc7XmH1s5cszRlA7
84P9FDZIuUPBQck/5Fced2hA8r4yr1if4qU2GyC9Z6uSq77QTSOoE8t2jWB0HDlI
q17gHsocgdARISQUpedS8qHPPjHQK5OLnQf1HZCKSR/lR2/SWg5c6TnRKgmu3UR7
mptGB93SnYiNjHquOCG7oJ7E6qSMFpmPGZsYRdvR8Sg+GTDMds2UNfacV5tE8qbP
TviIV2Pbo6RMlhJC/I2zIKe23zplWfHktZn+WJsb8A6ki8Vumq5wS+D24raAysbT
uZJIxtEXhvglGKwT/qRTBAzmDmAX8zDcUDZZl0Vj3lfS5QqXkil1UR+0/aHuHVqt
kQySpf475JZeQiUnR1+0lcURE0UtMKCmpOA6YDM8JMWXpChQTObmva57atzV9/ZW
cPbjjtU93e3zjwQaG3tKk69LmUBnKr8d/JO8dR6KcUA36TQOGbSxC0uQ8gKdrM65
pMjywlg9d1qK5ewKiD9ruX99nG2Q11O+9SvMHxZ0JHLI8k/B1yn0BuDgBx16Fwvl
TQWJcX4JCxQvhWhWPaFnvTFCRTsbuQfZBs1CTd2N6+rRZdCJjBt33N7451ZKa4pb
Wxa+PblGHqVgX9mI/SLyF2SFRQP6joSs1mlXLmbk/CLa69YUuSV6SOFPk2Z3Ctsm
M5OooDdgf1QBz94c5wwMC/aJUDeF+TVjIZTH1CfZqH/DitWxM7LgVSIDQpj8dXaJ
HJJHzJZwRs19ruH7DcHViHG7Vy1M6+CAVcHJ+yOkoRPrA4qVcVIUVihgSP45/a34
ruN7HhUYqAxFfHaeUoCa/sIlmFxBPzSP4Kni0KB+cZYsjyaG0oogndGboBbrHtst
Ok936WidKGxL6EX/qZlqYj1/CSAvcXJ8AMnGYEk3saF4Y99WLs7PPK773GN79nDu
mwrPVI/Lvj8ruS1LptDgkMgscKiH35dHzmFpPFFEAY6mK6muybfITtxbN5mnaD/+
2S2yfu3+pZ8MYyBpGg6aHkC3RVovPxqWZC7pishicKJG0O0utkH7MnYE0WJWk8Im
yD2C1g4PDHLhzHL02HgJLJSE0YAyUg7d9+jasJ+2QgFlR7wZQ/SH3WENWKm/lAl0
LZ++Gt/UsQLSK6nJZQrKl9cOF/o2gyo4rsgzESuPAA5Bsiyc+bKs1Lu9FhKbXNAc
FbiM9IyQPtpofTy+8c3KEi5my99gxUXnrwUbQgjTm+vQQ5LAvYAO/9MxeLx+FLy/
p/bH1mdgrjHyFaCIbLKRynV+7PcPyGGL3ZEFiGctCpvW+Cur++PoaRYg6IQayKw4
px7pDXr1m6XJO9GmdIsQqdnVnQsT3ufkQzwVbsauGCQJWk72O8XpF3bcao6De68q
AKDWE1dYaEEyvF5AZntu3dkCtCwLHqRgUQnbcIYBUXhb9AX3HEm1/wADfzh3IvNx
zL/X2VzxVOsrg26PYm4RzXbxaxAa2blxqI4kbp1eIOznwETkMWasePJ78BJCIxp6
2NtbUuKs/MMLS/DW0xcSt2rZXID3NQTgM4Yh/y4CFZ6QcgefwcQBXa+WCOgv4zkE
ef3eqSkSd9ZY3sH59kmuPuqkZfXAy20fLK8NUPqYznu2RbES3A39iZLCUjoWT+in
Ne4pLY4mdH+Qytyw873NsksyLEjJHtgKtkf9uSbgb78P+M7gJgIUiKkR3M+gg7Yl
xds5N0H72igGJZVK3YwvE90CJ36W7pncMAlpv/1KWVhdvegokhitXqLxu33m8RsC
tF1KCIdBrQ/AdElfxkHrVWXovDDl7vfsX7pvTaYSsNyTGqid44qf99tXmmKw+bk+
M4UQA3u9FlbbtzGfcNn8LcNp5R4oXaqLZMzilrAlnwHRICZz4GUVyM9uB7YuHJd+
gdKSKWpFlvVarjDuaUSRdBFs+wECg5+tWaaYTALLAyE+8YssiLCJYjFbEtKzW0pM
qJbb1sLNaPfJjh9tnsmX2aNgKAm14aYfNuMpy0v2lR0g0a36qyfDY1+DCcddGWr2
wQLcRz5uCfoODri5VU8DJNCj1HJQknYWMfPCarMG6zESiXELsTP/KSd0psDINjXs
o6aQv3dVAijptsnedMdZou1VfOqgJv78zmSrSjliQKNWp605DGt/p3fySS1sgpH9
8aE47xvpdzOMa4N6oYGbRWoivq55YqQS8KqBv/zOMnZKGCUc8eziqfCUaHLyO0Hp
EQcDGJt4dbMpVddbcP/q6S9qI4QNSfp6LuL2Ocea5pEk2aSNVDtATyDs/ZZ5hbqO
OliGWhXKHDoeYnE/5Gka74aGbXr0ecVussoxg2d6vRsBdfFRzdLjFJtIG+MWhVPV
4SFPRuzOKWwRR8/yHl2MxRFHUlW8frxXjKeeRXMu07NV1CLz4ORs17/DdtTitpwJ
eykpF49hjq+mnL5HINCENFx32v6N69eFeA5ntvzhMhkI5UlTS1cN4aog4Mwpf88U
HaDDEQxHp9YWvMKsZUr8cfAiaM7E/xbsyrI9PElUvNzcXSaWF1Qp4/2OOLAAWwpl
og/sLd9lhfsOVjl5jUIP4KuBOLIQV/xGuH7IEtKVclh8IzTB7xDqFiDa2O0EoEHB
b0LzLAFIuAWERpqJ78fL2dAU5GV2Zg50dXPpjNPX4AxdK5jaLbIJcZ+a/6J/ZTwY
tMgx1BXb6sFh7sl9wpB8bXDWGVJU0jpG2xLzM+vefeykTxolG6ceato4HvN9jDoP
oXI2Pg53+G35POPAAFUEX6vIXkSnaTOXfdAC5zn3+XcNkg8OVNm7xRbZCsYdgbkn
jco3VjAKAuNoGZ1k6HyVWJ5xLPrUIS3MuQgBsCQ3lfs9aJYeSVr5lOgowdhw/Taw
ae56pYOrmiZUf0J6YcZz9RxTaCeJEL3qRUAq6ancjIW/WEZIXuT4PMxnuhxGLsKG
wYfM3pPmfrQCh7SoDujkQDIyXUTTjX2c/bXDyFaemD3HW07R3N3PAnUDOd0HGyjH
1KhI+TgiKW+Zwz49KjPKDSFHdVA/IN/c2im1H8ko5wAhzMQ8YqcvGLy8wLojGKaj
SHvURrPETOzMEoXZdv+6vsoDJ125x9VYzPWq3Vuz3O7Vf1KMrt8ePLoiOAe2eW/5
YHkOKknmiECq3wFL0hPco5KN6qqCyonR1z9lVAaRsHqB0vcZmixlqYfM0pnrkFOA
hOL6geKxNYEnZysctUUbFAHjv3TIFeYulEBlsvGobZSyWehi3Tnu/IY0strPc2rE
A7wv+Sb8jU96SM0Jr+sGtdIdIjR8fKg9kjTc/Cyrm8L5mcwYTlSfj9aLOAmrEoN2
uKLiGgyWyVoDu8quv1h3u4Fs0rq5FKLzky6RA2w3+zJfbVbZK9s6uNqiBvhyz9SC
sAXeHagqMUFRBnfNDopXbS/p0PQY13qNW0Iic9Ye7kB4MGmSPTkRLewJQrFYB0Jy
J1GtoydO/f5y8gketNdbUlFI2PxAf1RuvH/vl3n39IZSNDRJzcQNIH5olBx0XjZn
O4gLxYo9o1QtVXXYZn/fdnaC08AXC4s/MVNR/oNhJAMpdwmH8SArXRiC76yKBDpg
RfJkcRI2f/QSoeNzazSKf5gEuBWYgLoXjtonBhqhkqjUfBMD7A0VFB1dFfGftlzs
GHq6fe80WPrlPyCwT1zgxAgDbTjtTK2tNb21UnWJlx454zfyWz3IcDjYuIf309qS
lgSvD9pZjUsEornIgqtR50HMLL6tFq0ihZP6UvPtW5EfZZEv5M+sQAARYhqYP2ak
ieAUp11iWOniQSHn3eOqu7VW5mpnYRPKVDWS2yfvHkEsPozzrfisgmZi/Fq8Zvy6
Jnd+cxv4qiNcHdTvfUZGQHR4/UZIcKxEds5SoGuWSNgPomPvtZNKwKD8UfnGm2+d
D9xzen4qtiF6Wt1rxY3Fte1rM6bpH1C0bE8079Zt41TvhE3W/KOVdyFM0a87wd8M
LswmNZPz8rcShrTkCO3OJNnmvh7KMj8VzrDalzPBFMCVnWYOoY29Sc/XHs3P/NFx
WHPKvhVdk03vWM2+5d5eQ9+87t2OOch4lrSEmLBvphfDZjC6v6PRKRMMhwZyrAID
xyhAikBdqfKn3HgNrt4NYnONROKzyozpW+d/CHtMl8VYZwqMn0ZJjNNqzQqT37yq
R42U1qBFGJLuigQ3YjZ+4IcgniP8fupK15LXllhUrFg6uYsOul+d4aDErn48OlEp
ARr/PyIiwkJt2/0L4pISMUsY/tOQWkUN1uWzDmhS7Y0jKgV/R/ScESPz76oJpNzD
J5lQz6yosAOCnSw8Ws2EwkWltwch33BBcRdA9hfTvT1Do3d8b/tlj8BraBnbb9dX
6YyLoBm1niMTBI6Oh+mggtYAvfvY9MtwCdSBuz3XEpcAu1IhLYmFFXRC6XY83HSB
Di7e0SWeIHj7vYslxrLyVdg5b6jcOz7A0k3EVghFCYOdaDDH5AzLI4mV+ixFGC9l
f5osv3k6evZ2qiconFckwVLT5AsJYl8QoTyvfDZxuByG0jkCtIQ+SzhYM4bNFJnl
PFJEevqG6HXTlwO8y/wbi6ECZLw6fvac32fHTceIgPDhnJ8d1yoUeY9THZgx2wqj
dWBDAKcXz/mx5Mhuf+jnWTsS5Aw25luX+iaWelWEQ1dTFZ3FPY+ENM/iUTqfcW+q
kaG/kN70nhpGTR+Mhu9Vsk4516uAXOSfzw0wmlSDpU5Nx0td1PS4eHXui6lf/80x
7RdUUr0kJr5Tm+QRM0pNOsCbJI43SZkJ4CODh8XIOz4a7gme1jS44D5m6IuZl3hq
oBApgOdsKFNhll3bUFtt47RqNURk40zPxQYd+exmMhCzWTpFuPkKJ3JgegDL3GsL
1nFyBk/j2R2EC3sjnXfDLc7pcj5Hq7FAHzoW0YrgHn5BeN4u3KW9DdzbP4wLVQcl
Vj/LvgwNnndQPcoME6XeaAWpKJKB5ZOdE+76M1aDdiYWSfYGjiryORoWcxgK510x
pglGFbq1WvUhOBc63mXcrLMLiRi4PPxRfhogD3xFEwkpNf/kS3iABuseHZJxz/gU
WhnAMLWHSZM6FWCp85nqC+OcPXvwTOKcSuom0Q1XAWGvmWJGAw9sFahcqAH9gG5w
a3QObrK86d1bSrOupaJHbjh2/UymOhh9WHm5MLjzC31hV3urfahmOTJGaXlWxGku
Yxq8rygQuPyFqN7jheDiQWie0qwnlNoBp4IYFLTA+Z9NGnJD/X7f1OLEme3wzuYu
DU78iEXN7ccUMgOOY3PannzyJQ9eguJMvLzR/+JwkBZbDLc7dP+qp+fw5+wRzLax
wOTWzBvS+T+P6yJ+ge5y343L87jF56yaUEDpGzO/qitk6ZoCL6z/4Sm4nNX8jM/b
3vzhiWTlZYEEl7EWuuwC/Psq7yBtZGxBVJA7X/v4tBBzlHpzyq3zxsYHHGqUTBhc
KcE4/dm7lDpgH3tsUObydkdGTw3ib9jh5ojNr5WKIGAl0wTx2Ia40SKjwq78ADgv
lFKwLOgEniTUCjGdUDJBINzhf78C53qIAcI2tN0t/JS8tpPhIeRPphunWCod/q4S
UdLk6gxIURHVUP1sX3k1wqs54cuSpuJO74weMj9pHr5KiO/m65rPDGUAfyc/WfZL
2vl7s8CcD63YUrqz+DaSEAtmcycyVfLOadlViQ+zN2btbpuvQB/uqJLUH37qo9zW
gsyTKsJ/e11S7hSB6AZ4mH3PNVSh7WATbs16CcgJkeyyPks/mpL+ox0bDRo700+F
fkmphn+Ods0/6DWAanCEak/M7KbAMnsrPjX2GxvY7fOFUJVtytjgOkbqrCfC+L9V
hZ1G2eI0RoiaiM9YP03rIVctsInzOvsT/m39cp2PFx80JCrAAaiGr6/lK2ydEAcT
KLdjjfFOYFYz6UFp7pQEE0otRq3+8HVi60+klcO+TKzyHhyvyYFeQcqSj1TqVMkq
Mnps7pQBz7M0yatSCFB9knzEd51rqDt9kT+u/l+nSk/yG759P9qsJU96bfhGBvmH
IpXRFAZv9yZoK6tCVPRICHCweFyYg5YvusLaKRh3TcrdC11uMQraplG0WSJgM0B+
SBsw/qjvD/H2+pLLU25AxsUAfWQ51SKIJFymAeOzalSevxGWdWzoyH5sZrSZtGIR
Iidwue+x9uLbSGqJ6K12qq6RPKksWwgt2bomNPmElg3KsMo+itF37vuqaKJZGnD1
sx0nQMCA3eJ1YIAYbmhsqZnUq/dODp0mxX9oG6Vb1KPvpNmJHRb9rLAugW9iql2Z
Df1QLIsxgeBv8kBMZH/7LIPd9x7ZmKFYbIuy8PboOOPG10zlrfrolxOHZp3jHKA5
mry45fTB/7n/jr49bFkQAyDyGvPpaCcqXDIZLIVYCF5OMc+u/DE7PyMkMrBLUiER
7nvPRbN44oBMNmOcXPdT8m2ewtMAx/e+Wn3Hz/ZOMa9vBdYFEWHAP2P7R8fMtjN1
mM1jdzgmCH8zh1Xd7KfzqM6ARKCv5IRPRgGQtHujOgNrTLCUMJb12dlhNnnLuVmr
AZDO0djUhCop9FTtjzA6x4AMpfZgkgQgTEzMZ2sEEXR2O0Ai6K9zUuwcQbqv4SRB
NBM1pPbt4Gis1dzpxn6HwTnN52XBBJLZND7vllUlM1edEa9QWfHNQj9KUJhIp1b0
q1ft4QZIgB940AXrmkvb5RYU3W/KsZxA3n4lpPvsMDScOXTu9xTqWwnmC+TlpEa2
PWvF/GPqjcUjR7PquiLHoGnBctQwkNASVF4r6ucw91OzkTxWdl7qweKSFKW2k1Aa
zk8Tfzo4bcPgJu8L0y6HxGiQVo9O6jdFdvDD0l9zN9d1MuAYFX/y2F7bJ6GNHfAm
joRr1nX/N7LmDgjWLW4HB/8Hkz4NeK/hXyekrDGwhm6RaIEIYDRz8lpcvJRgvTBv
YdFnpVXmEYniMkMcp4lIt1p2Mzmsd3ZUy1a3jERf1KLI2VEzC64iXRZR4VHy2aba
otaRaNAdFqwjKPCtAkTYp5TvCqqWUgy+9avqR1CG9SpIdpNsCNAZbxLYrWUeykKT
krN34ZMohTACxExjZIPk72OxQ94zd3xIMCvQ6jv9ri7CQ5VSfkzIjsk9dQ/2eQRH
qOxsHU40yV0fO3RLgNcqTVNcpROD6nFl8EDGEoe7FpkX0yu2LaeECDghl+kEfOnI
WY2jM3OBZb1JfYfNYF7JasAfNSC48VQiJcj99H3JBAwpXFnOC6E0GLe1V/Qmhoz8
/J/cvNYc1+1G8drYTg1OjT44Fq+BDCArM1RgecOwIRKT1A3lPnxciM+VwHcUukY+
yISxTZJ80ZcvlqautWcl+Qg4MI8upOpsKAXV+GGhAtZqHJypiud5yQQlC/Xh/7Vr
G0osIfFTzqmRK2VGUmv7BazDPoZav0tjJGvgI5K3UfNLuyV4ARQVmPRebtXPXgDn
C3UDpaBqXjTIo4HgsykzD77VMCEZ50lZaQVtFbh4rHIwF9VFjH2Vdua4byntDK2W
g1Dhs4i0Z+DbrIcRI/KfApzWlst4dAft3dlM0UsA+9I2wk6R3F2urO2bngotxTeN
ZO7AFJ5qUMYi9IPtN6/EkDoxbBesnFfx9nrvyx9xdYkicM9FfzeZdFXvXs/nJxCt
8+G5MV/l7nhSh2zg6XSWT0qMH/U0mQScz/0wH2FG6F3Xcre5nR84x68s35Fd0oXn
2+6h18gTsHfPYHzbY+HHe5N7yxJg+xiE6IVfxxoKtlAltwy4UjtsweBGdnb29HLV
Rllxh9Qs7NmPDfUwORqsaErIwaP2J2jUr4Hxkgg2ZuEstNJdQj1eCXg0r9HEFtn/
PoeAqYNk3BdTfppdx40CTydQfyR3c1+ax0HdWwEQJ+46ZS1asHy264kLKZ5Pa0+w
DCdsHwGokCPIcvjEtIlvSQ4gqqMMxSkIvN6AwtgaMUvBbgxn6D0SFwwKaA1Q3JQU
mXj0X/3eXxjZQechGt15pURzX3925+jM0aEtO77VM1gl6at9nn2q7M28N+oI9pGh
3zbThBCuERlwdCqidaU484yg3opsOwY+aTOR31vKjWxWe1adX3tMF7ck5BMkBdd1
z5LMFqyur22wDKbf+7gO8x8El3ob/tZtnB6M7wPskKYc8FEqmnoCTxP+kSTrU82M
CsxIJwOoAz35SvzjrQHM//FRqRX01x6Nng8JB4/BnIxVPp5fj/G5uaLrpYosxttG
+H3b8YZOLNgYb0zH3kNsP7lljkz0qURf4eHxlbUnQaS88umzKqH3cG0c2qjzAvQh
dvpZhBntAD8mzSMgIm+1NdbgyiGbuuNs1kHVdgaFObsj2sPhrZqAt4H0ZgWvodNi
3iFdKkUkG5FLkR44bHPjA+WEUJiaLEE6m0P9I9fPM7LgdDnZj43MvuQfAq/ZC2hu
gxLHgdabzTjsNo9Wm+Ok30QU8vQlJAGyyuO4zPk5pbmnDOUzMT54RqLy83+lhN/c
BRuyjVA9pMi7XkzHIuUxAYdNcUt4CMrTN8PBkpqqcl86e6npDg10+utOAO+HuDTy
qoXv4zCgadFUf/wtfkbosbeap6SdjCH47RHjfSTtMkERzGP6op2EIYAD09vx0itd
XctI0SWOzSbTYPv+TUJ5uRJffsAGoemzBWCok12IKZ/G1YOvI389jGcShwX7sHd2
ZyfwyEZwoLaETGkYBGHv6OlQ1Yhns4KfdTO4imXfJmIfl2BeZ2YospiWlWc14FeJ
CkpDbnOKd1ivi3OJ0oCv8JXXsLz4pZMoXjiqTIH7PmnCCFXLnpPR1LfJ+jbUrabL
d8SfogzN+ffvPzWZ5UT6yXVxzNzm5PQLsFpdeVAeQ8SXwL/NXBaLdGZsAkvGK7vH
M8YNtjT5V6s/LP9cBMQofftDafQiwnOF34fe0Ky3WjkaM+HDobme8/Yo8Fq+EV8o
4TCrf9fwS0mhcx/XC7D7u3ijTZcp5lME6eRBXh3QFiMgazpkbzmWdW/2H7BnASGU
CCNyr58Y/6Jclp6Ap7NqjvvXAAWyUBtExFZfdl22aueYzaSJqx9rzhBzoVRErdC/
mfdZh8cTN05n6AjpoQ+Zs4E1MXjkHOtqCcOR7v7YB1Dh24BAd6ZguEOnHaY7Chv5
Bb+5Xnu/oxx93nYPgoWHL3U1EycMVjqnBj7h5+g6UA8ovrGoi9xmR5In8jPL2U8D
AxCxi8rPaJC3mtQ5S8PORY5rYfZq+vLAxBolwB2fgqoUEnpnXeIMpS9XeShOvbM+
hg+KsJGwdJR4Ma5XYmVJ31R8rmHAQKEwGivLTbj1oh4OcO2KMQUpLVMMf+04lrRT
YWFqYSi1vJt8jscSulimduiIgU7vnBfJh3n0AU7N8+AgmMjtD+0zu1NhGHwyd3HU
Z/rH8jC9zpeQtEOzIKg4L9Sj5T1vVRbt4qsHaGJ1w0/L0y7KuS+KYWbdR1VWuYQS
zcdSUhVcBMqvA70Km7hoICHxavpFcL42TZP0/Z09wOBSA46xMYlzYqgE7S6bKrvD
MYnCkFBE6C/HZAlScgiYJzZRp4L4mSguzQFfHbKSNfwo/Cg/pEkOZG7khkiCOIci
YHWuQDRlswxd2RwNgg2H0RYE5GmJ1dRpYAx8VuvflgCvl9YppmSiwfxlBKQbmLMP
NlzMJXg6q9EvYj1RszsL2hLR7/uag8Im4jOLl5pgB4/SqCuSqia+Ksc3JnKJHcOX
R2Pjp2Tjn7KX6WDGNizcDtp2Tbpmr+cBndIsp/ZlE76UkCMA4Lv0o/dz85jnb+qq
slp5fnGC8FiDjp6IuEvazouhPE1zqj5Y1c1lFigU8zNv9fVTEHtcCkoZpxslrlBD
pWBU+IFjALru5Xe3CCLhBPGxFmcTYTApaD238pFCzQqG1Wbe9C3LXsbNUyqPfhZO
XxT0LZ4cVsWyjofRgM4G5OYbCJyPmKW7c+sRssU6e/oL3L3tNzj/wO083o1yjO0s
rIeRqSUKzY+oQGX8Zg9tPFO/zvws9gpXfRZdO2tfeBIZca/RTxwSC0LDKg8tSwOB
5xhH4FnogOG5cDPmOWz0iOieBkRytvDD/5U7WomX6pKKjyMoQhpGwlRo7QB7mmEo
rBw23PYAiJgDHWxi9gwop4kmCeAHfr/op/IU0VJrvdePOaYL3epMwLHq/LPcAo/S
mI7hCzWOlkb6dxZGTs4fhmVahkBVf71+xH37/S5fYIijyCUrTbZycP7aEbCGaWjy
V72ATm12YkwmqiOl43mlPIzYqPUxXepZBH4C9i+0ls/QSdNbGRLSiEB1C5yKqf4F
nJAig9NoxwEzcoayNP8mFf+xIi3LdeW4dlA0+52wcuIDOfPg72gLgpclxmYqR2W+
tvG9Cn0NPQ6wowmoNl2VhLB8KFvSzBjPLbaC1UCflklR7tAv1Uc3BMei942szYk8
/ckJ/HhIpuIF7a2xpIkVaSnqQCIVwUy/rXSeXuaVQTM27TcVwKfpuryU6baiejSR
s+oD7xGRxi0F3EhK0pBEVbtAeL8yM8RWiIuguB+Ecasc/k9V7nuxsl90MOKaoE9E
JNRQ0xI1i1cyED5EU6Q2lQceRZ3HBAZwAJLWQFbUhWNyW68JpWsmkUlE6Sd1sIul
fjbueZbHH4rKPK5EdB+A7dYanFyJfqYBZNtD4zg9+A8jwdl6msU3fhYtiIJbT4hq
kri3df++5cp5Dp0kb8bZ8tTCTz5C95LC9hQMqDNzMpDSXNZQpjWyiZ/cUKky10Am
jRh2WVyMAe+nMA++p0yRrabQM3C7hRe1PLsoFXgb0/ofCnD3WPkWvn2brq/m0DFg
3wfHJY/dbQXe6pEkAOkopF9RFtOKGu5yUIgkedtVIbh7F03QXUUMq9Il6uTIafhI
GVmwVuJzDP84aBVbqQkygZSn6f3+IuL+cIRRauSvnfJcZAsaxWdQzQjLSrJJuUjp
u+S/QtwQNJfFcBXm/1HqvJO1d62EsJ2n1tsMq0xgS+uvcbtccM7cFjIL/SR5QQQu
bRERYsnwQtbaTaZfJ0J0xH/Hd3W39Yik1PaX+wZ6HTNiI8m3Jmx/PCVvSmjF9hFY
oLgnZulyzsuwkGCD7UM0kchk8b4gd/b/S0SFHEbnP/LyuxS4yNh7mTvuuI+wLROp
X3D601F30CXQ70uC1yOP51r/1Ig1IOmiN3tkcITfX3JtyWDwlJmSwowV3Z1m2rfL
IGaZTSf7Uy4DaVbdnJdKEhLnEpUsNIn/IfB0xBbZraHFZPoKBAD3TkYPmCVtv3rA
bOc+sx9+GlNljb0JFGqmuVMZfdYSBlvur9IOpT698HSdXHnYSygMdVcXypERm43p
kUaPRpj8ebvGrHp05jNL0fNogkuqvOi6i7lkMZHqElFJMNECGOXdxd3MagfOrKVZ
m4zfDbfPg5tr1OgjlQJvuWK4bHsrQnf+rTkBrn87KCe0QUvEWqxLFmZ3IRGvAeSv
lNvOCJt76ur74gn46dgJ6LUZCq69M8/xMD2kFGEh2lHMXlX5bWrEbiy7D2zvAS++
teeknkIgMEOBR2mp0rNfX+x/0XSctQ3HKD7pTUksf0+0/JRqJlRSkoL679jFwe9T
zT/L7+z9vgjpspHNxmGXhHOj/ZC/LWjL6zVqjoXbyXId9sgWwTyDfPFn9YTidAIo
a7uup1KzQNOBASpxlKgvJfG0QUHqMhTAGSLHQIvx9wRLj/5k4AzPJM9mvLkJwHpY
cWXdoGpblqjkre8WE2Pmj7UQUqFFVurexUdanwMZPmwWyFj85xQp605fKR8Aj+4r
vmnrtIixgc5wiUTbNqF3lWYQ0UwBbrBkxTkMA//kPJPvbA2Hn4QnCBT0kzLrCLec
nmsvVxx/41XtkKhWk50L+X4U5s+WHmtPaD1PLpMQuaqt/LFyCtKxrWQDL4w48iOU
taeuNx7kOJ2PvZEQUADgDwS+4imp16+YSs3MFYgbL8HW/7uHOwVER68RUb9RtRRS
7oBaeRYfTHKPpiA9DHOelBTvZ+nF/WfFp7Hl6M+sJy0tmiAd59R+AtMxrwxYfop+
jnRbr6u1u5BsyQ2PVSObilKSwT9vtbHnXANK/WrduNxVEJT2T8UU+ahdqNiTO9Qu
fVh9+4SFcMuI+QH0Ni9UHe7cybHKtIdJ8hKYtTfqzVEP/VnY2BEftKN6neX69ugP
uwVRxap0PlmNniNMpxhQxycvumkUwgPbxPQ+7Epaij3CXPxtWHFufb3Twl783Moc
kdBl3A6EbLwfWRQGAh01XJSi8nKsbgpWzMhkPD3QRvAug+U7M/twbkkv8r/ZBwvO
ofRyyknyiQUfBaSRVfxC0LcNQz/wOLn9yJ9NoGNXyC0dckwyNGxe93PTvq0JgncY
EKy1gzsRuYsCeZKjCVbZMmP/kl4qI1+vhY5wBjTrUgJwe5Pj3KWDMKTZeBOFJx7D
iT1lmKdpi52r7LHyDZH5jp8NoCPtqS4Sqj+FNv1kgd+NePpIYfrtwcJV1TrjcyY3
XC7i4AAIpnGjfuIs1RTUXctAybacBoushb2Nc3K5ldzdTiiCD3H+4BnOiq4e0/V5
04Xp+HBCy8eNPESl8VQ5KDc10Cn1AZdaGEeoeJz0uGXayHDQ+LaT0yTAWzBQuhNN
MPMC8v+yIctmNLXF4LlfFHV7l+gRqhO3tP70bHUStAVyryL2mSY9pH5Wo373HPOm
eIRgtWC++03voGZllelzlLqkPEyqC9Zf0H8AQXfl3/xU0Bzt9OB5g2qk/JCJtHO3
tBQyxJjx/MpewEou4SFYrBsTFGROK2+CNnMPzqnRLa2YOhHUbXWYw/+3b7Uhwf7R
Y4S59hpbuZ4g0e59qj/EJBSw7msw7Fwl8G57pu8t6VJ/dRw0x99Up3UmVKEPW7Wg
H93+DabUKJhIXsid0uy+TpwsbRes56Ep08iyAJHRZrzCd0guMRMnpRO9KL7kKorn
2Uh9T5bmwtj/E2ZX7oKmo/LDWgEQMbXb55+uY+OGs8Gks7RAj+sW5cxbY9dmPwnp
wqpb6+eB6PcQPwH1jBXf1veKI9aqvIqH1DMw2u4ug6yz5avAgIkl44bxwjxjUEMj
v1akJljeW+ZphALu3zyjOdOPR9lSFrT5G8f1sWcj+lGdhnzYrMI00KqPZcNFlGp1
UzPmd8Ev5CLTJQIDFyzASzmOZzL/yUMwvLa1KmufME5kGmvVjilVQUrqsbQUFqyo
vguDbS2t/RzEFbBRGKPlaAmA1XQYqpNN5LI1hfZilZQQD0VELzk/Xsvg7FnrQshW
x4gmBtenwaQNIEeGrStw276eaZTg8D00q6aw4WWHBjsm5b+k9xVdz1gk3a3av+Iq
kYBQOmqjIfhjVc+MIn3zLgKvQhr3rHF1LO6zWJOKXIy2TeRdImx2Ww1xfGKAkmVN
Pv5hyUwb8BS3Zsv/NCyS8AzrvTKV8xXY0RjTYPjixyITTkaRziXxvW1KjSaIlPvW
pBpzvmKNvQgZVWu7o8I1UQnxs2jmWdVXTTKRpsgClelp0HEAfBP8OqzxhG9aZSsM
ENrnXAhkL3SgtVJX/vttRgWTt9WtUSHu2/9NI35LKdkHod4olYnDK3DnDuIfEWw6
GY+9Y4x5NRm3JgbJoR7T8xbRNHBstpFWBvo8lan7FQahgkD4ReKCKwcDkHDapN02
W3GH/TnirFVDrRSEUP+AuQHD6BTJ5BF4IqrW157AOFotScfqUmSvrpF1SijLQ0UD
66T+Cv+CHytyLWrGaplRdXtMiTLl/mIWdnyPlzEasKyIk+FwsEwg4sO88BmY0INH
Xqi0XFP52xVSN91dYDkKXHSrHHYXrMX+5FcAtvYg8VSO5oJzw/3rrTOUUe2CtcyS
08eLT4D6CfPqB/wc0/nhswcRWUna5Pbd1qAhXxzwS6D5wdSjXZFPHd6voo+1WZrX
vH4cSdm20oH1L454vM84Orv3A8OHyW4m52OEDC6dgrqm7325pASzfEqF/nLsLtqi
hY6Q6kN8R4sO5iEdrqmK7bJ+UdhYfINTnKXZus2DtlBtGQbO4maOCRNVJ148Ugit
kv1Kw3uZsFhvNC0ufCItfXqop7Owmg/aHnI1B/LC4SZeRgssaje2a7M0OXphAxKW
q8KI4a7jXKBLdXMG9Y4IoEP6HHwzQ2LkYwJl24p9BHCCmZwzwKuETLS8Y9H+KVym
mB1Fos563uFCOdIwPr8djmXVPpGB3ZxFcry1V5WzzKAf+ibiYQmVt79Mm79TY5qn
rCWSBmjDd49IpPRBWWuIS1CdpFgtUHdFNLYHPBo9Hc56jtzdnZb9dtGZJRWY+Z4W
BFGwhrv6+niP9TSLgCYlMb0kQ1jYvHD6a489MP12t65zHsmjcY21kVb6Z1jjB4pO
2zfwRnraaz0AJVHudemPxn1z3xvyDdxP3AVK+VUvkVM/NbaNY1/UVPLv4u2XZ83W
GUoB1vRehg0F8sQqHet2SqVD8WScLdaW2ciYvSPC3TXTgfDT5FZWck78wMIeLI9x
IDdveE3HwAyvnz8sq192HNLlPfYS/8N650WBIQPZW/lNEOGFSzLygKmMSz08XxKn
zJG3ryjJjamR7F7xaClf7auqWToSg18U6gGKxpGVyXOEMxvEOpI4zhkKdwELXaQZ
Mx7zayQbFL2PApf/fNYEz1u+bt80xufRFYf9veo/tqRm5geUMhgtKEMcZtV5BgJJ
8PnradQVjBknIUBC2uRpGWfFUwyjkmskiTT/nP7j+Cwsx+8mZUJztioFGccOAWvo
wb1FJZpjBJV4bmcvbU0VttIdWbIVYJFwb8yNRtyQ+VkYHqNj6PtCaGvfs7kuDlEQ
yW4jkmO1jT9+YzWQP5dCpTHr/vB+ySaqpMnBEn8RbTXcJF7e95hPQvM7hkSqp+4d
t8aV/cL2hLN3Vbn0K+EoMwlqcfIiU445VnlxXQVeHk2USmtz3VNAJ1TsarKbfb+O
UFpuztUHw0XDxcgY2qXC2srfFHrScq9pTPWxHP390qLoXPnKvhu1zNHBSR5i7jxH
c5CTBNd5uGOsa4edATgFQCeSh2VMs+nntsSLIKYjBrFWI2s6HN6s457apbzkbgmd
1Xz2q/079Dn2Yl0XLj3E4hNOAek+pIzHB3n342ewtBtCiKHEgkk+JBtOLclTopKF
9OsHbyLL1+fZf7AJ+rndVGxHUkm86EyKeNjgj1gLDmZWTDvaSrI4Msvr9ZxHWqwS
aeqyaZU7Wlp1zEjFOK9g3U7/utRRY+9Spp+LmwwotO0Mre8RFE6wKRCy7kVIF5T6
Yt7pHJ09NVOGNvjBlPTZxVjQiGw9Fhws/UteCpDl33DP+1bNZa/c0nRa5HEs0atn
3F0uxXuacfjaEeNLuDZmS3UHuXgHE0EIMg41GJPBsBbjms3Oh+ow+x4CdMahABD2
6ShMq4qUoCoAwVhL4Ne5L+xR1E7+ADmpM/caZ1kStVoX+Q5uMSpM4MxGN5aPz4z6
yYwWTMiLf816fp49MS4SBn8rp2pXMeIxrcMcBSQOu6k5rfCpitLHIHagclZWULjs
awbAVojySgXsAkRjATzYaOL9l2UxB+1hg7YfnR7Cw/1jlCM+11+JKRlql4P4RAYj
w9yLPhOp4lKobt1S8mmFQJSBojJzz2yExI9Z9H+ctZeW8oyXnDeqyDnGGfN7Y6dL
GTlhV1J150Y+uir9mgHA7LwwYY6mNiDeOmZppQq3xcRRd5WJcxNkGAN8LRd00gMb
R0dxyUK4VQ2GihCTVg3cPDV6miuSSu1sjh/+8HNL+9ToL3hioV4O8kO1hMR53V4o
iJ0TthfWLbjx6GtEUTXK91S+25FCYmMlV4BJUQrmhjHJ/Ct1dfDFvMf5p5M/OD7Y
pRanNfc/yx8nT7pHmwzmb7v/k5llwj3YCf4S+5xMTEBgm/fWWxdqyGFafR17CjJH
ki43pdfcZdaaIKEX+2VltZQ9D2LonfxVvJA3tXFJFeFMRTMxEQijP0JN1lWnSo6Z
pEYqff7bBm+bIGGozFGi556+mSQiEwE1fhGbUdqsjkQh75o6CVD6583ArEzEEvuU
9haXmXw4mUTvSSPPsST6EikviwmlTxdkj96kGmRp4hDDme406oj3ISg7d0I7IcTX
TA35kAV7pRyCSCg0jz1DvEcTzMx5TrYY7fPd3j6V/sYATsfELG59vhRXIEH4MSTA
aC8pXh2SMyAS5MerMRQcFvxH7/UYAxQjZGP2hB2qQMZNh7/ajDJKUfCP/bPCgj25
ljGVwAjhN5yil5dZvaH8mjNc2y6fNA79dRywve6q7/KvezwAhTTHqB/baz71/6ll
+gNuU2ZC8uXgH1MfihOkkVR5PNcaB1OF8/oTcfojwJHQRP9Ymvk3QVxQ2UCgV6zt
jzlry9nTvRZqsY2JKsnEJTFk3RWeKALGkqIUGEPP1raX3pjoeJ3MlY/yO5hJzDJU
KOmfzcxRzy1e1132UyiCwlARYExJUx27Eiz0/5WU5VTNAeFmnQRhy7g7J1E8T4a1
rjOYbHdLF1c6C0u+g9M8UPJKXXkVMMxbseBsztYkM/us3pOLtvz31+8IgFRmQFP3
AnCy8xvZKd94mkK6CwBEGMHQbb/lzxc13Cg8F+21Hj5U5WWe+iTqf8JWPUBxIOII
d0VpN2Hn+SUstekZYojhLrq8UL18x2zos+j3A5y9dEuKdmDhgYQlaSYhWS9DwESJ
MBp3CmRV2Mdf/apMD5Z4xAVNkdXrwdxLP/QhY7eCdPapBEJxihbsISkcBCZeh3+a
psoQ2BiZ3ftZHl/9gA5wl6AcUJA5ljQFi43um9Z3pQ1oGuHf7NPnUjPP2JNa5MN+
9I7hVLhxwVfoY8T7qM9wWoPMIAdUOhTuCXvqdRstxywiarXrUh9iguA2lRUHTF71
GdvlsHrCfNpO+VHc2zrRVt7TEOVi+8/Mu/QM00w9zkig+lIBKcVtgSmqpdH8lZ3T
vNysFJdQqRqyjcnnFCb/l654iUVZkoFqCTircQ3cSubcgU69Y4qpLgz7sI7JDVoe
hRHf0wp2Iz19j+w4Eq1S2sgLAXiM+0oDy6K6r+wV4JWIC/p2AgdNln2FvneluMR0
oF2cDeSoLi3KOFx17CMmfrrJRXQ959fNQibe4s/kmQ55Z3JucCWBaT1sHjXa8BKp
YRByg8tJviDh15A2PGfOB1g2K9SzG6QJ1g9fg2nBEOFeuDQDXhp8dENgf3AYfjNI
qcNaC4+QhMyMAjLKpSvu3xEPth35WxSnIhKweqRCqdoXKf1dONbQHvljAPxUFW8Y
cy3cjRRuHYCGwWnAtqRHZnajs0rqQ2Kbu1S6bCaZp/nd8LPqI0VNpobMGoWTa5pD
XWap6Y8wBdYQydN4LHkKbEH8/btFCPJx8aS/c6KIDNcoV5JA95p4+nkmO4z65bcZ
JLcS85P4Ko44wkwnvZ7t1dstfncIhFUjrw71E9Y1KoGyBxOeJ3i3Gvrp9xPQZBYS
ebF7Nyc/Ztt0Ho2bBwxAFNYNilEIQGnzOtIaSzcOjL9h6wT5CjNkCA/Re7cHkLNY
b074x7g6ueBAhyj77PyHoeGBhYwIamBr9p6u3kZLy54RxHZinAi6gy+c/SgLohxN
DcWlYb6Ill6RFE2VnI/GepETKJ9iVFstMx0+k9yrHSrJfWxMgT50MAtRZXCKfzbE
JFSCw8sDRNM011E7E5+HI+rVKTRAHztKqx28dZb5+R3mhpzvgZKHNdNUMMAhq8tM
3K9EjcyGtzU8KTWy953vXII6poYt2UauPjcjuVvfWLUmq0wQQNfYJmgPNkhI6jJT
2hUM36mQ/1HpVm4YIdYh2V8GaSqBH/kJNEuUcJod2JGIAvxFpjrlEI0Mcl/hvAOn
+cZ6QHTOZS3matURNXUWLpepnAzM12jBimYkMyBJu9ifTnnsHXYkaOhNeHeAVvh8
1JbreJcqVOW8fdrSa8shejjPwD9abdzGJPKN83xtDhkhCw2PgdUakum39tLGo488
CDq+VYooZ3u4ehKQiqNcCY9xar1F5FQ+Pl3o3ZPWrzquzPQOkk/AmKTgZU8fzRrZ
7ayxLyv4hwG5eVMLlFaL58BbhuU09s9EnaKUAv5LVhWvPagDwPBO5avr8jHUqpYT
vuLxUDmtrDoJgRGMUteZ4ItB9C91ZTDZ1oXS03xAAi4G9Br7x/3BnIylIlg8OvKM
DeJe2I3UjGd95E/swx3i3sITZUwWQ3pYbPFaO0KqCtS4oGH8gk3MRxZlQUwjTw0r
MtAS5JV+1ecjX+6dewVltIf4cHw7HCk9mLh1rghMlbQM9+40CHKhpMpkXMjkrerG
/2JtP4lX1fWOK0iUu1zeBSDc/wtRiqHzzjJHMDJJjG/idT4s9/vtFc1Ph8FOzjTP
BUB38/+FCNrzdw8eXMSQRQGA2jj5ocgEa/rJr05onScagP/CI6LokpweZaGrie/T
bL4PSmvvG1C45yMHvEb1o/xMHZot6vhUn8yEUrMvUj8oqayyj8fySRiTN/V5xlgM
nco6brADQ0/1TJBDx+da7vJtuCX1pruzP9KGIVlSp0vV5VOaA0xw/J4KYKrq5w8U
kyW2nBGsd2FiiaMmZdifnvOKJQ2QMwa6PKTnHk7DeG2707QP3p9Hw5eIlLxeAaTd
DRL1yNONhCKcqwpyuUx+7wyyclBBesXfzBWpMnkSNpioxTXRMAzc6BLeLMzHTGfN
eoR6HmsEbH8LKKImMd441gdcQ0opbWIaVuTAE3pS+5UKwxNz5MMHaLTE667SOWXR
0JCzbYsH6wB4D5FTcq7mTkCeY2Zk8ww63smFLRmEXFsPoW/csHvN7MnCbXXs2YB1
Sd28Ah94BRooZ02qR3ry83hXcd7W4c6X79F5V4RX1/OYhE8HIdrKv1a0jppn9adl
XMLaMq7ELJLrK5vXyGdWnn5wM/U47b6TmQ8W9z4XJ895mmgA2/3QiG58PU2AK56O
S9rhReWNZS+x06SWaQATCVDoKuuSpn7oEMGz/QXD8hDD8XQzYtc8zUACU+fh7qvs
Te3zKpB0IF/CABE13PSq1XSn482tsaXZusrNOKStLJ5DsJR45ubU2hHdZd1T/7IZ
zmPpbpklcDLOPh1qb6vb5Tbmv8eqsM5Xr7scc6Oy7nsSBsrmHcZMiHtdOMGnnTIw
oy2ysfzgZzLqWF1lDuFyy5XoAvRMHYO2EBPOtmSbEThcQZ7lWdCCa/VhXzyN+1Mt
O+a4Jh9fzOFQCXv9VSDupVncA56wWwmjjRexxqlYSsv5kFey8LjfXAUXMUH7Qq32
Lrs7ocIB4rBNofuSodM5jEMIy4YtyfptlAXq6NVv8kdTHKHmK1AbbWKqKlhC3gas
lxB2OUh7QgmQpbmoQ5Q8XKshcnM07MrBkKlEtqHEjs43Np9HB0oUOl+e3IBEqPqf
5I0ucdjK2/6QrDS7W8FOX55mD8xr+1c80dk0CQYdLw3+oiTjGX6qqPHMZvZ+USqR
+SR9umDtsfJpRM0ad38Vz6Nh5jD7REsHVihc0CSruHIZknqbn43sjoOBZrvm9db5
zfERs/GtXC16dMFtknaQZhHVlpqc/8/FT2+OT77mLfdMV0gZwViOFiCOiJn1dxLo
13cBp659oUgZasP9V+euGXno7ZamibZzROV/kcccnPcALm/exfhCFPTPVXonZoKb
3KYhjxfFwn/UC+mJyT7cc4gvwL+H6W0aXe1qVR6kTGPY2wfJYuwxVBI5rdPQmeZC
qkxbjqtBHkjTKdLySuuBXN7fsyWZqE6UUbXg8lPT2hwxTfyhdHtp+k8S4qv7/sTr
jqY0NDj2r1b5dx6607X07nEtj/LrMIt+53hkuoeq+V/gWG2LZJxMvBN66h3QaVFa
1280INxP9FVmFrEsIm+IrevOuymyt4pnNUbZKYlGQLOdIGWWMmuurt/rpyR2NfkM
rJCf04qjFMtE7R9Psa9eI581PnTgMFZKgLHJbrRxzqXaFDW0frXubgDMGeZGX5YQ
HoelNmip93mwsWjNVRzAzvuCmAx89xMJwzFBaJcaNovpgZV+5xO6YnpL3N5nHBR8
RPk5ErQagIwy7M8nu0eDuBEKSYwWFdy8VTyYMKm+7y6GmHOXy1bAmtQGSu9Ee9v8
cTjLkDJgmsXfE2OcuhBW3JZ+7PNPAg4hnyYpF0nATK3MGg3MYeAFVhNN4/a7YDjH
3z/akn6hUiaYE6fUcpybp54PhzN5g2Otg6fTnRREnNdogFYEJgHnw23Ff1lwfC0G
jxtRlAv9X0YjRNVm4wupEZ8lv8wFv/fvwAtoIFgHU27G9n0RP042B3e21eSJlyOO
se5rSyhiUumKxHUDRTKW8C0lUyU0pfUVn6c9fBdR6M9kuOGWkI9iqKjV5yCQvF5y
9+VqDidLisvt46+Gfz2h8hKgzqIOxi1vF1HBA4rc4o8dJwaVNp5P+XYJzGdOG6ND
u3kL45JaNeOhfSSFBd40TipPo/pTB4qVWYQEFSwZNY0hhWRL0oiTIECfdSebQQ6L
WDfPfncZI1gow7f538bM6olv3+Gfj5gW0L0baXOeRCyaEq24ZLh32JEsDZcBganC
ugkO0XQYgvyFcYXa4LmXhpKQFzoztBGYja0ZbehKVMQh6lbix1UAjosWU+kurOeC
E2HzXWYL1V1fqlMZB69rs2biIr1YWD9sYx6HLYAYap7kUnMVFpHyZu3gxZE9Kmo/
C34khDgr03b8RJXRsK61cUn7HDFRNBGVI8adXHDXY52MXB0HTtacvY1i79cciMJ3
/nchi3uZOAwz+yQHnmQgIobZZ/WGsx2g4t7xBsZT7Giv25FVs020wMDu+zEqKGOD
usqyjDXyJv66pQ8u4FHN2yWAHM5x2sap5EWhh/SQOXIrkFdBP53CAHIp4CSjIjcx
F8RtDoBwjhvBmxl4VzqOd+VnYXS6jfxtbiO6Qf/HY1iDqX3gmibUDP4usab5IGS9
r2yJyKGg+l2KUa8qaNH73JtLQy6xHsb7MJWQ8cKIrxbWJ6DYdG7exjud2goygmmt
Hg4KAWwa1S3MhIWzx29YK8nsbauOvv8rS0vyu8rEHB7fmrYdb03xzYyhiltrRwv8
zqPmolXaeax3GGoppPcUyli7daDvs18GxwFiOaDpqQXhsIwWKX+VIO068mxO0XnI
dIXE53/8ecMrMe3rZH75/ABeO3cJYLPe6K0/v0uNCtJZIs6u5HHKS1AsVI9ZNVEn
UsKlO7CTBJfRfWphOXg0qQ/HMavdQzu0EXkcNSDaxPRZJBJybvmczaooszzp6toP
KhxPevGfUb03WeOx5zLrocSXOshIthWl3AX5G62Dw7jCQLVlSvJUZRJ6IyQdjWvP
yzjq3ZdYmYWboeu2n1q+TnVvetnucueBjUc33cgV27UyaHUWZbqBvXIXXSx0Jqsp
VpyEDp/PmJUOqj2TI66tzcDP+WKjcsHhhwv0BZQPaP+5jiTYMbK4r8dEzsx2gh0+
UUypfu46mQksFkI84wxF9/jlDhOwkDAYwOsbEiqVu1P0b2ZKGxtSs33wZg9Jb2BA
kcD7JQSvWAoNYgwls74vFdTtahdZRJtWDWbDY1htNiRNph1BXe/2/KNCAB38bxsJ
KOSKPZp3xw0+MBGP1O/rMuA+uuloUsfnzZ7z46zytGFF0TeOGU2mtIYt6V9YOGiV
dSuBr0VFAIXFw9d1t/0G0G7dRRwpCOLKtaqjr9frsWPEyS5oaBX2QDnzLuUlx2GJ
s9LBfdiOGCuW7AFfZ2MVr5gJ5nuq7gADloxyoNP79FXHFeLSgyKXx8voSXEz+Hb3
xqGDzJh35/EH0VHEXhpsxtkwMLeT68CnqZcNm0QOZ5v6YP6Nxs/+X7EeMoJmhx3Y
5h24+Ob/R7WV3+IAP786gn1akirr44P6zk5Vij+CMFdIpQDO/eUifVT7+jQo78CE
DGTmV/CwMR545a4Q0uKWg1NPVp3kMxKft1REjJ63eWIUDwWAv2ECqnqYBL04I4mZ
Xr1qDNZ0IdXqpjNFb+h/bOlr/biRfHHFxV3aLh28c9pmHCyb0Blmp7YOLGryrSka
SnT/duJ11WlMBNVyCFomL8F7RrSQQWZE0YqYI8FU05Wm2SdtM39sX+TCmxElP1yu
ymY96tokdlZ3pBpS1BZXY+iW2w5CdY9r0bGmGQ/c2SH1OUUbX0hEz/MgUM+mSP7k
NuvJvI3HOD3HkHYF+BmLKtZMtz8n6LbhSCVx5CWz6L479RzlQUYam0w2SzbU/rmw
SSMiPj4/s8aloaPydt7A5r+oOi2S9Zqah5rSYVHdx79bQCSOxAHFauWzAmSbmUXz
4/y8LjsBcc0KQNsTn2sB496Dt4FOWm94aFaJ082d1icD8HotewRxSHcC+9FUp3yR
D4atC7lQyQPd1a1z2mrpHL8sPuAzygWIpVRVGi3uEWYWN5IFahrzaFl1oRTxP4Hi
0HKk4YHPm55bzQ30lrnt0+8rQY83vfDNSLrPk3M2RJ2JtbQFjj44kxQzyqDPSieR
24L/kUl/4ACm/JT38Mjpyyu/TNxArixkGmrKtswZr5yWh48+T9b14USLHVqCFWwF
TWt+BCwwuHqoq++9w4bVkpRoIfh3fbRAhKxRTtxBNY97ZtonKocts7Mj8QtstDD5
h3wt/hid+wWT1v4uUoIymnPRIWs8HCSQQ0dmoRLgC2wCBf3VunGm9d0A5Kotu9Sf
mALLGXJ5xOXjA0fEVp5EP6RtoH4nFgi84Z3c/BoyF5Z/mr68th80SyA9mvat2ATv
l8+hA24JHhSTTqsFfyk4BM/h1SXj0ZXePx1t2YeHBMps5Wb8uJi33bpsu4vh62Zc
s67KMqk+1TH88EfdvtEECBPGQdEHisj9zSwspuZpoeEq1JD+1AO/jcPsNSUtD88+
5SvwnoavaRv5F9t9lKvPKv/oHU4RuwHc5uZSuNHSsn6HIEAX5QhDgHyw4r6gmZ9I
cjrgzqr/n/ir1suVGy4jhqTSGJ8Qud0198e0SYnqnoJ/0XxLy2rx8TaOLfq1e3Sm
A+S6oRWP2FGm59SOFFrqTbV83fH4KidKBbzm4Li3uDruK7Olko0PogkemRtBGsnd
8BbPYOiCKxEBcIuOVsLnupNj8dmJBkajsO+greUigfmbjhSPJ4Kz6P3B8CKN79nN
32x84ugG3CwigxC76OmWTpNOpY1xZpBNE+sOHgbxLpibVdtuX0c/jTKeY5ac4kWW
JBOqxTVl4nQqLuWL9J3CbVGGnSfhxjaYeZ322lPZglYhMn8KHUYdYKIVwF6skSuU
ghame27awgKzYZ9xHMXd54LBlR6pZOjQLE3ODlfKqxM+aQkJWQxcxghZQP4+zkUk
QADZAS9DLrd9lILeVcmysHpNgbx3P9YSrQNyO6z92Tpp38v1/lKwxoBYATsZWUJp
7dT5pSR0jXFnpd3zyRGxGVrITzznk4+VD16y4uIO2d0AnyniDN9Oa2sIdtwjnzUy
t6MKxCckE1WqRQOpyb49VjU4cZAQh73GbfUSTplPc+gjjENQz7ClCp2Cv+6Y5RG0
mEMlaADD8vpeGYoigBKuTFpELFO6b+yS5jnf7M5nVqdsOeHU7VF9bfScUOcHvSsO
ijz9Wu0yXtNBDWSfeZcBGj844ovQaX1btKtaHoc0b58mXFSrOGVmefveQeX7W1Wc
qjihd5z0CizluZLbLfzoL5lvSTg8hH/yTtQ835ty5sosI4A9gTR0PcZ0w8+LwuE4
eLHyzPIf4PZnsHMCiL0rxFTw4epzeu01gR5mM/3juWpou2AjTqJPh1sfX/XzvVS8
m6qDnNv3GZ2MpwVVcsY70A2QRLS6up0GpR7+l+07xEfQV/5mgNekX7NMElB79m60
jrgzxCnyC0uGrvK3es9j8ofuFBHEpplLse4Lq131LjxVc4sVYKWGMNwa7HV5YDLo
UYx3xM/GqB7tO2gUFZUpwMWarDxo5RLCNQccxc5vj28ELcO4i0iefmPqRyYbm1rR
SFsWKJduaWZwIG7jemq8khFq8y0GCZ7tOvaewb/dFhx1AHa0FB0XVrM5xM20mkvh
NAVHeORziHfQhgbp4AjxTt6kheeLp8M3mEDuyfphTjkS0F7IhzPfUSsvEKSW2tcp
5M2UvTv2DKkudADDr8U7TWaoSokQ/rl/DQXXKkq8A39byvkE6IuOfMTYawrYKWxl
ZV0/f1VfbCHU2WhsMEo+h3DGbjxU373mSSgczhEdZQOmmiAzRZCIhpsficZLLlPL
S8dDK+jugKYndiRX1SJljVyisdqmNiAbmwMsDwrSPg5ADzhgOLe6zWIHcB5o5FWL
/34vcyJhUzaOlMfoaZdf619E9y2bH0nvgufLwhMqug2SAe4df2EYBPs/HD8vlkAM
tQdHYh8CPHnI/j4FVXN9eAL3Y+h7uLzyEGSc07d0kiTFysZEvbIQCd+LtRAkz4Dq
qziarcSIxa7WdjSwqmqirweu4of1ZCDcDN22xkESI0dsVy3hpHT1GhKu2LQ9IJT5
OG4XkUNuyCH0RR19sO+m9owbK0KUB46YehJlGjGBNcqvnM5/ETLWWRsPtMX0ZvLE
XiS5i2Us2D5l3Zzul50Z0kmrFKNS9Mti+wJcwemjioLxo8RrQT7kXy1QcxQfSl+/
lfMhYraj6IhU0EL2hRQL2RZWLQKNZrn5zo7KraZLCTIIQeTqDXCoOEZD4fQboW/q
B7bCVzJ8Qu1k9sNsEPURzzEbMCLE06mzKHzAv+jK1HWZkGN2zPc9dORrM0zon1KA
t2/z+7MNXXLMOn6k7tzp2PhTqruEnyQCv6afM9U3KKTHt5+9BOOb7HLXL8Y/5obp
RsHWEfx47RL/7lgXjsN3aCZp4O+/LQufI3LVpRNZiPmD+dvvoseDL8tLWt+SZHmS
cFbEZu2yYlwbCQAiTFZQohuxVUYTPsd3bnISsdNBNdnVm3y74RlDkKXktEZ6Yxr3
TvDMav0+5+nAHVQNjNazUQW1ANestdIb4TOgn5cz2eF9cEjq0z/2MQpSV1PqzrRG
91gWvF4tAAusQbFX3+aOrII9CmpbYQBUbPAQbLOqnB0GSAcD61A4vwbZ5dIDM4kZ
/D/rdHUpOwj9IZ/EFRCvc1jKagI6VWx+WHT19Hzt5xvSKSpadhZuzpM7oiSNONFc
bb+VgVsN8ld8wOy/5ZJrL8+kBA5/vE9KjLKEHvYUIUJhOd/wo3ZBvaEbtdhFEJpf
SqGmk4emTEnRJeROAUA0lKKhs2FwOKIVkN2FqA3zjqYRY3TClzkEQyzpR7fQEHU2
5iONTrIkNQkFwWRaMsWxI5fikEk1OCT145PWID79ZW0c7dqAIMivq5LxBlE+Site
EsGo/Yfq0IgW2ojPpwYv9d4cwlAfyRbeAZbGC+KNAPaKb5b5LgDM1GgBTTsoXBM+
bj4IgnrFd6QqiMFIT78vSL2PHT9m8YVLgw2PmqSrEYW83iR7Pxx5IRGUrOeTlyk6
V8+SHYSobyaYSTGB5H2cQilWyiQ5L4iJ8D+arm6LGn+pxCRfIgjyJ/jdUuSQ2Nho
+yQqsZb8CDomTHRZlO/ZwAjKRh3/Ar8tbtSMZ1boiqVWIBW4fZjeURnSuIuFw2Je
w4CeUYk/zV2Atk+/Xv0Ey51W4SPEi+Xyol5ehMCfjFWU0FGBphUA9m6j+hDhd/O7
YtEPEVMdkYnd4L3LAOkogBhUGVMSe+pl358szytg5DtpotT1to4dgmRPjpT50g5v
thMTRrl211cPw1u8H8C/Am6ncebVQUZR3OSvSay7n5rzAFOKq8YGetZ6U/4Ep/VE
IlSsL96p7gRngJot1EcDQndN5xTiYXOovwRXM326yp+sCdhHG/dzXexMpU4lHA+0
gM3kWjx+ZoejQv42p0J8qnnMyzS+6E5dPhX8dcBO9SkToaXhLPkmTqNqSJOfJGUK
JPrABK4rAJ+RN0o9+RXjGcslfTQ2yG/H+45erY8JfYu+JLiY4JqWzRV6cG2umU7h
AmyCiDYz5goCLEbOYRNwejE9ZIHYiuQkMEM2izEN3PGLDEVMe/5jfgXS4+hVPd/D
mscYwCK6M1D8GXhGsYnHCNtGLvoqD48tsyTK8N40Ptd63nhde/F1nVwBcsNjrpJ9
2UqayUSW1uVGm8iRVB34naUMjusLuYMwul2EWKhdoe25av7MaHKIWbEHVxdWGZKm
Uu1oF8+i8rpEGBvfV6oME0/taqUf6mD/hwmYN5Blvq7QBHvJhBmFGumADiv7g/PS
9RqVBBPR3jkB9KfLbcsea6oY7xVZ1StZ67uTQBHOHqhHChYKTCyg1mu9yMFULCKt
smaaQg1tY9HkUwogJ3Z2XNIpaWvz9iGFSZrzsRJZRF8rHxqqe4rL6U6evfCXR3MY
HqV3HDxpiFLfA8WR3v3sMnwgi4hug56C8FPLpTtKawABmnf7fizbrbOi8gbowHO9
FwcVHArV8o5TLZoTzNOmGNxbZ6CDOonF77+IS5jScvACwPCNpM0hpZBiZ5rkTERL
XvKl30jHYMoy2BM0Ok5DwyN0Kfn++tgFazXxn66ahrR/rFCs3Lt/zpd5f81VFNli
x64uMkxRBNJlADAkJxEvTvEyEZYoEbxvJP5WimXrvSitcyELLUUAG3ZalkI/+Bk2
tb7WeBtHjQ6zms+cbMDv7VTeQ0aYCmOn0coXIVWTQWjmILkVXTKOnoouYlwBSmf1
VekStqTJRv7dK0yDPo4caec0w9y7qss9o88sp3xeTKhnYa7soDny/qtyr5Y0Nm7k
+qDpqBku7IL3DJbMQTS1/DdyllKgEYDyK1WGhdhJTBSRYNathSCWtF0XaZFDkj58
YF2B/aWSof9Ran7S72jvO3R9BOaCSlmAe5PTIsDrK/XLlTL4dgbEOfqGvBXnxMZg
ICIihjRaW8IYDcUDZ68bPeQSJZIVvYubsR7kTDAxd8Uc4x9y5sNWu0/ctLqBlveo
SkN4nMOoBFhTsLmeQDE7unCZi1iexFefI63bL7E/JVNNet8ONjSf7Z5Px94JPgB5
m3FICn2lhg/rLhTpGHibycTxQ31dmVdfREvIblabeJU8eFeIbesR9jvTgM02TuU0
Xwq/oMdkBldYDr+8KVTI5BmNQ2RV5BhFFjJv+mNYqcjRo0j47VUkedHuSFicrQJT
4qif5ldlF+e7G/w1n773Xty4KJQUMzJBqMplSSal9Sq4mTOvvXBpIliQSsix8q9h
ORxxN6/9Dw98+K1wDDBrT6RU5TS7JJZJd145RIDackWI8slt6bYXCqgpN8u65Fsf
qUhPizZpwjXkOhIULjX4Nkap8moZEmZNRlM+kn2T6WpuGybl49W3kHhu1xPQj5ys
WBKJZy4CRlKSE6dkCoUzQevPVcGGYprXI2qFIIRYfKpWa/7Sms4VKY+tcM3etOkW
DdSHw8F5gRkTsTA6bapukKOKUdI0WxxwFRubRJXHS7nyx9RgeT75UzJUBcc7C2dn
mtS3v1PGeOqtUaDyja6NjhHBAoweuSimk4X3I7yIdYu1grgtm+QIpPxgsZ8j6ueR
WC2jnJsz0QKCyPsYvvBfJk6NLidUviKCtonCvwSC/ulMTPyuLqzBuhKuOAOp+k/T
15o/Aj06wfQDTW9kwlnI795j8RrsfH6O9jO4T8uQ43tLJJKmUIZ4O9FkbaYm1NY1
v0dQrOCoPL5mPvF73XaT81GpV+I5+Wk/+4dG4Gjil2zqaUhCo+C/KzW9H2OsAePG
YCLSDgVoMrs1ZJcza/5Kv4cLVF5wOvJIL0cGzFYljRReX67jPnMbaoCs1+o8wuRa
RNlW3ydoe4FzFMxnMtcC8XEC2s31zfHl9d4+O7Yu45BNCzH23kmWAo0I1VmIt14l
YAIrnZc716y+dNH+0fHYG09sOzRZzgw9Oij+UiWBfH3f2wi5NS7W5gPy3ai9EgOT
tQQjvGexb6AaaDZz1+KdHgp5oDemckQNZCASh0cRexIotjui+vJecAJbj1nQIHvr
YbToCaONwlROQtvZV8FrXLkEAFfUcVvGLNB8VXZDos/7w2t4rhdOw1QRzeCKkty0
D4qTFp1YlO4G6r6SUiFCBfUNqAV19wVBIud/YHaQUV/Nvwv0IP5RJWLMEwu0FBFh
hc83fpPFOFh4qNrA0FlXoDiJvqC0DCHrnGd9FiKGfp27ima8amWPihKZQJOhROuS
RdEB0otOnX80c6Q5ILZe7sPX56qFbdbMqEYosDzlYgkKyrH7iBKyem3HODWANEL6
xIAg1FDWhp/WxWP71+nnxTQHesDI98ebz9xc9F34mW/WNZSATsPK5SRASZeUlDUy
EmTE1ZJ5Bj15yt5+ivChNnH4/1rECRrXsBY+gcOvDeLOKL19ce83k4LHuASoBrsr
vA16rxhJvVQ2dgpnlrqd21aNhQAO5ztdtRGNFjVvkB++mRQ5DIjetB2ny5Ef2Xg2
TjFVHG+FR/uPBOhNYGZ9wSo6EqObr/CdNNRfkgghxHmW9BUuhOST6COK+A8hAVjR
mL3vxWK0gWogrgMvCa6xbpQVfGhB0U41t2zJOmdKSkAVkjAIEOCBpLwh2goL8y+/
GK90ziqZiTvi/mwF9nByoTV9vh77yACfS+hP1bPYvb5K+YI8aaQrWI4YnJ8dPWc/
1G5/P1oRgyYI+rfNzimnQN3G4tuZ/hKuGaSDZQeWBNCoC0RUc76LfWwl5+PGWZaC
5/ghFN1YVbyhJaybIIPXsqWuFTZ7Seqm0bMaWjjl759DEUWvfYm7WTj532U+X0eB
jeHoJKUCsbz9ASaRNQTb3q6QU7Cu1bppUvG6jgIQfoemTTfLsJeeeVTjHKZOylpw
c7gqm/cKvIRDsv2D6+9knluBkW4UkI3lQ2Ar6gyI70jCnwx6GYIglCX3jhN2/qTS
SldzOAHN6k7tDnTF9nsOAZsxjYr44nwJNaAsdzxvJT9THwptJxED5xzGKcWSUDXr
QR0MDYgKIN2McfO5KrujReS93SdMhfYojjXGF3ddjR/B08DHkqWyxO8FA5Y5bWUe
EjF0ugcj4OgovvZpqzSIbL3JDQlsLCT7VBxVT+tmXoIF8pKiPae995HxKwfy0dGq
gAUdViglX3SBd5WaHjmNoInCQQn3lzrcAxMneOIdLSFt2Ja68quyNuZ2vlU+kFGB
Ot5bP7BxYs1jhdDuDUdmU0QltCPRgjJZIuXfs5TOPIcwloXSBrd/PdFqms+H78H3
nuJtbTYC88rkbEiwiwxRqrwG+Lq8Hh/abJzFN63nEvHWws2DdMZdYpk19wIekTyV
CokqRnP1J0vObDE73y9TUMj2ZVyS4l4IFOrY85WAuxXoncm0Gz5TlOlL2WLF7cvP
MkvU7nDZu3JMCMT7QT2juziMK/sqF790Ibkz8sLW7cVx276yl7CE9zoqHbQBXlqF
rypkXuVln40ThoM5nVI2Q69RJ29UCLYI4O2mmemRsVeLCFDCi9scGyJDdj9kDfQZ
inDP7krPCoUN5QWkBWv+6h0Iag78Cg7Xez0HOqJQnZhu1GOeW0xnB0Dl88uUixGb
TJPNkZdkeMM4vFUav3/o/Xc2a+b6/cBZm2QtW8DlK3vJXn0JBpzafsPKCQuU5/F2
cTf7CUre9c/qV9Ed9TOiOdVjH5qgVB8RUVxDwQDvZK8hIGTLCmav9nXkNeiXEjwV
NvmTct8E3Z3Pyd/otFRnUru6U7Vfd16gVSUPlyj65U2g4EDI0cDid/6275HT873s
P5Zz/0WySXTfUANHMRX847ZvCC9uMvgCVHg+g2Cxn8NDky46SnclSnV2wIKHzjNN
fuJ9FtJ7fFXtBKZvjDhDQpH1+9oraqbB/rilloyXIWPBlIlQeS/drggpKViCpgMs
wh5UMM4luyX+R3CD9AYY1t64idZDNqffndRuIxXpEEYd5ZtSCLxehE398tfl9SF0
haCTsFhYr2eKIIaCgYWyoAsd9a2SI9Bn/eCb3eOUSdAvlHnnKayihy/gL+ntb1n6
TGpLwivNldWQ0Z7QBASuvIEXDOqY0jYaSLpLTVazwPrgrpMYVqjjsbgeamPSn9Y6
SI6cekfBmjgmWdJEAPzidKrNiNZsLvCVVVHOZIgfeV4d0LOAMByCFZMTt+xEBYJN
OZH6ZbqWQPoaTq+06bPpWo7T3TzqgfsAp93Ct4Bw3ADs0G6ukFrf5vgRwaqUvSg3
FOJy9nv1GKleUZmcTIpFLSTSFgC1KeVzLcDsWc6wsF2KVs2f3Ly1eUXAVTUjnKaF
DMlhvp3nXejv7ChHFbEUrYqJ5MEEXBkoN2LYNuwk9bbJG/1OrpDelZmuSRPRbikP
hC4S4rm1cNP80nfQiHjrskwONvE1fJmhPUG/kjJ1Azy4A7rvYyPpWz/rXcbvXWmc
UCGXidpQrmjZxhXxn3ObsLOGNpF80AgAn1Yda4hQbjV1l6JGRyN0mKlR9FPjF1uj
W8TMeCwbtErs8nVu02zwnd6e05ge749YCxHb3GYhZxkpmGyGgajDZAWSF96AAudY
FpC7fUrqQ6psQ8m7UJdN1bujz5i8uWhvYQMTv56o5bpae+lYX/yrLxUQoi2qMgIh
HZFG1erhXTtSB3Ydq8+S6i7heh7gKc/fDErniai2+j3iRVBroYNbD4g652hiK5Uc
u2EJRO5PM7ZybE1qfe7nmSNHVEmr+VO+esmW8Xk4UJqqcwh+0baQTLeWrZF6eE8J
39IlpNOcc5Fz8f5SkcfaHJ4KdPfadposOimBkUaWgb7N00p09Cb2/NIFQKOYfhE7
MxHofzwC3mnpCLyJCcQf7mi8xzE9gCYXbzPkzQzIzAU1g26Gq2FzDS4J1CPfwFWf
kD5vSRx0Fkwl8fk9G9gi33gNwvIlsui0XqiBrNxJgAshv7fA78dBs4xHARWyWA0t
15MtzoTMwKXTIQ11LbNYBSJZU6Vc9B3H1UHjlLngK/Cl2nxWR+3S8nyZ1fiH/ggU
fM5BPqYjB9EyBgKgFVugkscB8v/3dj4vDMQA0UwvAHSjU6d0TS7AT67C/2FXF0CN
Jld5clOu6PpUK52Uf8lGgi+O7M4JGtKZDYqtKUrOGmSQAGDqSgudF6IG1RGWXzQ6
sPv3ikBNnsHtSunBglBfsuo3rE9xxwSf8OIOMFgYrmvOszCXkrqeS/fAsNmy5Pbu
F3Sy5FeB4zxgkfktj2JoaTzA8ktbc/IpwTueGpdxtCKMtREHAzBuHRzLuFZlUFRP
eD3W4SJkQaHyNl32ub4JT3zJe6UMV5IYXSUmyJHkHPpcnW9zx8FxUpTCLiRvDvJd
jw/1gELQlBMAm67yDa2prRLJH08uaABDAMI3DT2yZ0KzFKRtF+hUUJ/tY0duPTq1
dHQEiLEATke5k7etcEFULnPJRyeblUC18sieOwXDhlPGwCT9WiqOhoYTpoxUaW4V
Vo8wKEmRXjhHk8838lxPHafvQYih+9zmkdxiI/8woGo+HFTll9FrcR6gyKRKYU0W
DzASqHkm2LfFNs4pTDFqJqwMU4MYWoyl8FqHszBGTHM1q/dVawURSWS8ZRQ5m19e
eLYZ+H5TxWc/L7iJMgUJZi3Fuhph35L/qsLOqDKS1ok02d3XFJtXXCaSnn/p1Vsx
xHO7rtuygVT4BNGotMZ1NnpmciShR3srhIg56JmUPaVet2Wr8aPEOKgtiscnZZlZ
ZEmCAmkErEKEgw4U7/pNDfPM8bFSmM76C0dNTB6ReKuS8jZ9HoY818Yi+Wo/UGDN
TJABe+TEaliRCOp36WduevY/lcLAGoq5uhRmgLOS+L+4E45spf0Mvt6E2GIp4I6D
1H2IxsyYZDlGSiW68ir07VWt+Vwme+w2K8acJKssdNWS6sB1iTuUaEiNHnPZlvYM
CX+OJVhr6WKAzRrS1My7rAv2BD7nhNT1kEJIVV5y4GjX9dHJ6csgk89eFPJoksmb
WSYIZLCvnnFtTO6cdM1EmMUWDz+1jvaHptKP+YmsP8McGLFvQ/yJHi2jIGcsCYsu
hFjm0fB9/tuBxRAElkLZ5TeMofY1NoPs+4XE6zJSkthYdUvGgozOJ19w7+vHybZV
BLlTD206ex/t9R1yuP9F6m/XNelkTl5w/fYjQRB6Yz1JuJkvgbgiQShsU3dZbd48
Y8WQy/0ntFq+MSPbvJeW9eXV0tOCbiwJVVqwAucQYxFbj6A0Yr9t6K5kqhP7nGw3
o5i3+/yAIZlPBP39n+qJ8h8EtpnzCwVwmc3bcE7L1TW+RAF6a5Z73WulItnTL2TY
cFCYbVa/VkGf/2AVgrWQOcNx0Gfg4cADkxGVsQzkxQ9R1SKtI+a+OPSx1ETUtqs0
G2l6TsCAxcIrj58AzfSs6CbIm1Jjzft/1TTpqIcdXcceVGlSxv5hNGqs7wQbcVS3
ASRY29g+Bsh9NmDWRgzNVcsb0HHZ8TGTkKYtm7YIGh7bUS1+DkXYzc6o6DfL1u/w
DQjP5jgQWEfBGvObF4vk4FSJzHb+oaiddQPC8AsM1ORj33+PpSDncQTMr/06n1dg
hmle+e/zDp8N0nU+pZG6H1mfvo13OI1D1ZGWHmWqPWVZeeOMq8AsgU1btQqNPUxs
cmRk0ZSzeufKlRi6w8vohbrQL4xlKG5ZSHwqbZstvCJmWA/GsOSg9fMh3GBtcyJ3
TR8t4gA1bD0SOdo7D1oz9/LXJBCu6rlSOEJhM5317QqVYgP4ixSMmp4NrT4+NuCP
eESmpaqcU9//9Pv/IMoAmmVTZESdSTY3Ehwyt1wqvRx1i0lpW7DDZ3b8PvrXUcNy
1iDi6KtshjGbxE0Tt+oBKm9vq8+SWh6rdvFpxXvtC5gw5gA1bThwo+KS1F0ruP2Y
a/wFugiMtsCtdNY6OiNPL4YpCUjlY7uS75+kjy72EZJal3A4wolmTsl291o8f1HG
6pqorySzr9XUNtokjTygg2CLYTiDhZU1EdmjsjyotlvhlWLkdESfxRTlBIAm7Vre
oO/gD0TLfy9Z0jemWIXt+nJLDjMlM1X9hJtob8zBPfDCmJ6N9Q7CCoeo+0COfDDF
dZZeUgu4n+2Za55mm4ZdCYnPezD/L9sJbqJ8qAhVAoWBeN9UqoGHs6A/8+ieY41T
Khi40INuoAD6GiJelNw9+PhIGd3L11OVwpe7W8c9H6MygCk02wJDyOD0Jw5FIZLK
px4S+hC7wNE4zvP9i3u+iH+5rTuWqYEDbROUD8FyzlBxPAT5IgGDfVgmNOx7htGQ
sqS+rxbw2Bd04kHEhqkF2skhqSsdgPbP/sbMWpm41JrYnE0nHkumsUcq7n3vFZbl
GjMlfX1DCA1hJdOP0UThn/2osmKNKvXTfw9bDwl2J2ccrTnOedZ1Ajp7aVVIzl4A
1ytpgwJg859dozWEkYRj5hc6ka5wU6hHLvMSiJtO4rvSF40zyyAwJTz+LeOzl/Yg
D9juTYfG95uR2i1tJfAd9Oz4oA1t4T3q0cSvDjvpXOAdar1PeXS1c4zPIoGAQzqO
K9+0lK6pJMOcxGuvqv7V/9OHly72JWlDfbCsW4z5yXi3ett76SbravIKBTruEtTh
5apJGMMBMzv7JCdaUOrs0iASSIkrD4bFEZ9QsG0NnZBRGfJs1+zAwHl6Lai2oYv2
mfaDQD4JBZdLM1/ht79X2i+pByCB7EJSelY1MoPhjnB5iBMruTaIULAoko/BpGkB
cEUV+zsyfqqU5ihIl6e0THgxltNPrEYXmuTaujkGkEE2/oHIEQTgC/aEm6wSUrMV
0xVgOxu1H31YqIIptTtZB0c9jW2/MKG/sdcDK2F6klKD0ACKXtMbuuxZUHEUpN7m
zsfamopF3RC+aeMBX+yjjKXrLQ8QodU36WYjn/M+zB4gsc6Shf2KXaLs8kEUAVQs
uGQt4vbA/M4aSWPwVpxl8PlBGMntCtnxWHZs1ENc4v7bMgNcLanE7qqhZCtVTtiv
lE7VTcl7UV0k9ws7/3V3Hp9kLC3GY2AXnND35ACoNs0bHcUQN+JDu/5otY3eS6ya
OVLLyqWr5ZudeY26B/nF5k58WWPH40vahTADZOIdeGaPtzqOOqMl2o0VFunMtZ7x
e4hcyj4sW6PdnBHmo0xD+PASD0JcnflH0H3hfGca9YqQNZJ8wGwXKCTCebfG+HCz
0Hug/Wzw2Yn9Df5neHlGm4I01++RULjItByA3+OzfxOoe8BKn8dX4CNF50Xj16cn
gZGVjqD0+0/aBbLAZhHoP0rzHc4Hugi7YpPhwAt/ab4fKlOJKITtiuWZVnLHLCoW
pmO086MkAgOQnfbYypo2MsTU1CU3GEuQ9C6HkRlTz6Q5Jd20j1oJjgCuTagIVULV
GBVIskluwx/3KgN/VvK5avZh8Blt36JuFs8bsBh5Ab2dHyBZcEbAdnd/kVZrddBC
NMt+ER63U///AzizVhLxGSVqTcz3wEObiEDSsfWco8aMp7zZIyR5G1IVRNa6E5s5
LgFLfVuMqqURqFciQD0hhLQUxucLt1f+3gtkyZ3zp4nhrZ6KJ511jr5xzC500l/c
UF5IZQploRSS/fvcqArebKr4FlIIwh0OuvkW/MWh0ckY5mSP3tXqK2UXo4/dcNDo
mETYhvvn0OKK+jJEDCl9hKzoKC3P6QYC3w1vDSg9YHjZsIz5OFRToqSyBzcz33rd
uufmYW8rHdCqZ00zXiPdh79cjx6h2De93+/YLfmLBrtQ/ofZKvh5kqc60OlZ0gl9
Y67U8YSQDuQiV0gwSGrPyR7/DGQ2VwMO5pifBBodoM3ayJO5i4z3YA6U4Vg1QjCa
LSKKf3WBAN+L735NPVwvvBsjqruNk2CaJoqvTmDqwfIWWopCFgsBWBBxA/mOcTNc
/W8UKrKH6CUxoE+vr1Y4lFQPRbtWJhgsM6eWwQHk5CDwPShoeJOhETsczkQ9U+JR
AvguqKpyDS46vcwcg2qPyM1HnHqGLEbBZzL4il+51YV5ZCtwE+7PoIv5U6wswzLh
Zzy7bMBeFtVzdtptwS19X6yqPgLZR34cm3h5wUj+4TrPTnT6pGuUoejPCmC8Qj5C
adHDhb+hU8Pj+3BTR1Leaq0wRuswDTVH0oqBaoG9ei1zur+WpPnp07yRavUCoIfE
wzZl6UhQUgxStZdZvlMnXZyjYyAifHTrnAkn5ieqFt1KyDM16pZfaO1ow+ihjuHn
16BGJA/h7Vh9v50xykSOphe5AnZKg/T8StFCvX4AZpCAgjsyd8aKygLKhTGYYB7h
1/9KrbQO7hsWFIXe1veJJvq/wm1PMgGGUK4vxImyqiNlTBynu9tG43rOlOiaMiNC
Wids5pBk58c+BsTlIiQEcbwyk78MlhNNARXuv1KP5T6LQaaTLV5mf3UyISZr/Pta
fGY/PlNV+b68pnuL6qdpodTZqYQKYOjiYDyivK+FF0QXPzDmCBR2ck4iM8yK7QiD
m9nN//Ltkjmjj8umbUYIY3q6s10MvWvlRSJ/kIPBJT2W/t16G0m/jeECBmwDUTEr
U20hhjbLBoHEOqOCejAyram07D/ZuECDzFyhi9tvOus6/KWaFUIdSUJKcJL9LCem
BAvHE+pVIaUQXTnjAoP9LIR1batXRpMLPJOzFLZTgdmtkaBM/VYy24epJ/3RNlXV
W8GBIweZ9nTOCGTgrG2djt/I4t3ztJ7GyO6Uqzk0dRkKyZkoowCI5yAjNbd3orza
vDapNempMvQGrfD/UuRYmfFN5dedQvmGYrAHOpjdBAA8m0d/KhQ83hUgEIl1qDxN
bOdKF0zgoffEzXWOc8rvByrIqRf6nLBkiGFMq3Aatc2NsyagjXsNv2d9Zdt6zyoW
sB7uCwCNFy04pyVqqeBDEhzqV2DnlNb9B2ywcd+h5UxBCIlzcEOW+xCkLhxyounZ
TQQBYbXXZpPE3bKGd/9ILEyM7mMn8VkCfz2GYG7+GyRsz0KeTSUBFGvpekeybxV6
USCMjnwRehxc5BsBUABG4JfH5uNCKYpVt+0gP9n2jte7vPw0FYtaa1O/SYjEMwiv
gbqiF2SsE6bzS+MK+/dCbPPk3ilUeGsmvBkVR+A+A0Q+arQ+fWPWhn8mIP1B8c8f
28slAR/yHCR4Sgr74Z+QNDVPW3VINvzi1vNjIAb5kSlLmRcepGsLsrw0UWkIhjkW
OEEet41l2/D9WNfZCR5hvpSwjyCSGuNHunl+FdpuBHokV1FG8ZyLIhZtBwRgH9Bt
bbMCOWy+0JRIsu4TjT6a6dpwyp7g7ViFayYpB4P+Rs7IzhnMHBXyTBwBMQuuyfPc
/B0fNky8xQqXjxWCxe7FHAqAeoby/VRUWFktGDMA6oaYX2Ukwecg0hke0GsrwfIV
4Ukic/cq5Dy2ukiQDXyRNqoH8s2KcpXvTBreMMfyDwzt4vmivd3M3KAMJhdyMTCP
vfZJsYQKwblzRKLCv/U/sB9sN1Su72Txz8D3f9tw/+YXqVlK13TALI1ImtAXxOjS
zT9xuE0Ty+gZ1wX7lk4Vzg9Nbdmzq8rrSpKAH/oN6Adl96xuGMiOk0KXGuX8cJSj
VWl0l426aIZLDGUyXSgDz1EwyU8a9WahxXMiMbjm7Xt9AbiuIDEJ2eHW9JmHktKQ
Vu7WMmaMvKiZKmZk2Z+71tTUccNnchvIpPWx9SZTxP3EPqIoauABmHjR8KDmkcNK
TyIT17g+pPV467jF9CoWoCbcnZMCkA2gpzbVJ3HyWsjMNsHILIjtLMFfkmEhMi92
I372LiTIeLSqlqtukYXK8iBlj3H1IRIxRfLaod3z+a+6hE7SJVzndE2HFuiRj7hr
jlhxAWoC/to7QQEcsNpsslodpWRYjIf2wKmgawSeLqfvkr6HE3AFwiWtj/EgvqiA
Q6ZMDbvwvF7Zmpx2KZBvfst7xbz9zDhZ7S5Y7kxawD/osfQnJ0K1M0vs6Q6Em4Bp
UUZVVyQ5rp4rO8Uxk7Zsv3b1+yOgkqCSAFNLLDjJD013uc3zhflgGw30YoXSUYHc
7WDzq1y6JT779fjXAMDbvLAH2H/uL5kDzZW+gc4QEiIuErguZi6moEbMIpw7zROg
gUFltwGlcRKLHCLFZCHOFHdWrLW4tCjVjclEQeWoFEkjfKL91CsabmJpEekDg6Iw
aTWdoVEYZZq57yVujg7XfTyN/i8SMv3xJeoQBtyYGSygOqN1l6ZeX0ymnBQh0EUE
CvnjaBlWPer66x4A1obQIg0Siflnz/NDpfqKlcfyb2BrwT7lIh++sGzGUD9LmqFT
ZY4M/ia4lTcu6qJrWhiQ/UTrVnHYt4un67+rCXSXWbbG0KrC/rEYFeIGkNccH+/C
35MmyDTajPEe2lQoAG/CjgGkRjCWqzsxvLdnOmu3iqNO4ZEpP0Xn+mSQ5lre1kvL
6s0uQDRwMe7v4TV9sZ6TdX7NmChYqklNzgyP5bZkocYEA3yoMpz4eiwVRqHoUaQY
gcFK1LJAvpZuIyvQ/Vxrbx7jAEjy0R+vFSpN65QcfRpPHXmiB1USmurBEO+1dmpe
7q9AD/c7nNQit8ddD3V5jmi6VJFBv3MHAUdp2NsE3hP4zugVF7NZob8xmRmVhNMt
pFULPoTu6lk2QbagpCqzabFDdhyiuFM8mlM2V5U2gnpYLcmq8x2pDap2vBxKmlRK
4y7k2xpF9Mnk5BEEEsC2X7q3RVl7EABugIUSRhfp05B9BfzUAKtl+J3VSfqs+PFs
1hkzJBwXJkBRh2CtaO4XG4JyXDg5vuEl89/CuM3TEhNKaRTjIfWG1gUMnNvmGy+1
z5tD9Fu9dcOoW9VvOKCpoGmnbpOfbIgVrx6RKctkwTWJHwUHxveOjwSX9KNIKIDW
9afkBfpQgXaQ9oC6gQlAJkrYVoZ+IVjuOD46Lg+XkAf6CRGrjEnLgOPfM1oTszKg
SxK3THMxqOn2rCYAhq5bgzc/BiVt6zC8aXTVKGyU/JCN3/QzbM4tYmmnHYwQgMRc
aBCCa8f0mwBGkYCEhzcDGZN4jYCvsK285bd7GrYlmF0/7VHGORDd6cWOMpPoGNXr
KPpOwjnNKC7GbXeiIlSvPDsixw0wF3tIfGQcO3AEOMsQ9PsrVMIA+p+c0wbciF5I
0NEPDTYx1cun72nWrjB2xeZU2VLFb9OCZQg3dJZa76vuh3jd+J09WIB43xYP1EwW
40J7o1nN0VOE6pFfrYSgvX1IyG+lKa8Xk5Jg+wpGgpGLLK0HMu3lDIPp8SPvTT5G
qqf76bD4aVMfl+rlzf2LKqbsWWfxeGKi4LoEoyzqEARDfQ4VVm9paJMDsBNJIJzp
aXXYoqggdwB4ABSUw0fwIElOgOiCffSzapU+DfqTAIs7xQE5hxVjLHWkM6zrWLIE
Tr/8NrtRUOmwriqBpfyoT+f4gF7i5ak5ImDw9uEj9rFb8kFWzC2DH6qx9xNktSg8
1beNdjx17f7B5Y9VKu919+XBMZzAMvICM6QxZz9DsSyB5r2heUxAhZrhk06lSQcf
5F78k0RRs+veQC7wT9xEzqj4gEhdPWOKQRRc8Ysd7gFUb12cTFGFI5rt067CcsXO
tQuXJ2xpBmgFEj6LGmtac9FLBuKio2lDjABjggwmFrCtZs9htb1CGNNsZIhGGUhh
dMEV3vdCnkHmK75iDkos7ycKQCWAdZ1JKgHvTY/c58MaqUMClfPckXZM04SP/hGa
7TjHNF+GBY2tiKiOOmsk5d94WUhsKQNMC+qkoH2ZSWrUTuJlLMoHrD+wjxvaFSrc
MLmfTP8zCXozkQCO7Kjz4voN+ZKDD6o0I+0dHQanfgU1MSbRr6jVoOLC+EOGaMJm
uv/gpJKGHkQL/HIhNCZqznd8bWm+idSx2L9YCYIBcMqMnesdPdbl04VRi7WJgyen
VCs/MrQfFqi7/OdRV23s+nPiqN5tPLl9vTl7PeUfTKdDBgkHmORDzCGTYLSnOBzS
7hrggZDuaeR0n/1zjWO1XupaBz+j7WWrSR+PbbSN4PoMPuBhwEbooiyT+qLZSlTw
oC0ZsYUDE90R+iuqRlQ30Pv3jqkgnN6sNSlJ0luy64901Ma/DW4YgaFAsgsTAx+m
OeYAZgvgkp48fZ+RyPEi7XDGbxlg5KO/vekkwCO4P41Y4asb17qzujhbslXpS35+
vgfIa/Ni6vX6SITZ/x6FACFQFS+nfqCBXTimqbOZoap3VzVwkDPgplMRBppLjHjE
vcAB90JDr+hIg/xYky/UC/Zt5Tjz5PqJT4yBtGIw0h4aZpRhDYIf8bYB+WKA/cJg
pVmcmdhDRqz3HRTfTC10xSigvg4BJcvsAtMbF96VLKLEtc9e8XVNFrZAz3gGCMZr
Wktl4gD286iSIbT8nUaJudGcKolizXPXTyei9tH79p+PZKn/Nc9Y18yTmi7AC3zb
FMa+RyyAQMGCEU+TXMfM5F6JvNKn9hVbKf3qx2FEobVqwkL50scqRnbT2h+DxfH3
fw/U78NcUlVFB3koYuDJsYtv+buiRtN+oDPQuCzl4GNHfPLRnb99gGvqBr45gMad
S4MMkJKujALMhYgJre7EqpIVBUnXE5PsmpVik/H+7DldsXnATqG3egUevFl/G42l
19qRUFiT2NFQx7tUBtiqws8/WNCnJj8+z84Dl8nYnXOlzME7Vvbhr3XELHYlqdv8
x3ZARAk2uEfhv4AnbZQ9X3UEwEGUY80RM+IZgVV/3jychugK04F+KdGIujtkyRC9
ItidTY3k3JMaTNMwl976Pvv5BNBadFIdBZ/g4IEPkpBUKpCTPj2kt8juC6VVhpjq
e+GFQcN2+zlZpsgNOQUFKuIh1IQfSk0FbFOnHN+m4fJYLJ6AmsB/p6SRe71gBZpN
gWhNE7bupEIqXIL2x7fiYLqo3cgpIGb6/cxtSnSq8mp6TtuoSgUE3aVGh7+6PweQ
0ZP8fwfQRj4qpO/dhXzlUKkO7Z4fKI4er63WDxHwko0BCaMiaRM7dzEDaWyvvLb9
6jumtrMptt2UuTw0AcFVseTKOaSByj5YQQ9msXpJDWYJWhSMGfiEmAT7k+ZWTBcA
bGyD0RqdJAs1DuioHD3W/5CDWJ1Ra4FsmFKlcZO5cyXvzjLX4dDuYgjFZxx49iVa
qCZMbSYUahn86JuqM9F9N7RBbHbH8oo7rYUywxHRg6GvayQtKjyX4WaA9N6tkiv6
dZmnBJWSf7jHdU1G3n5g3MtRA7WxusWf3zng17zqHLe6AGgzeYnYpkHDBiUA0f/o
XaK2p3YS/usUvPr/hDkzGSTflClDS0M4fZP7lyu21JEVcKMjey266Kw85I8gA76z
v58zPX5CTYHUF/K/5Op+0pqKDyPAiKwcrGdG3TxdVD83dsLw3sytixRRtXZbx4HG
STt7VZyFwajAqsrbUZ+/zZwH8zniTyI5eWcQbemMLB2t/EjOL3XOoGrceP0IlYRD
3tfGehbgZhpkKO1JpbYL8AoZt4Q4DO/r4PPqx4KWm8//8E+b5G+LXQ8N9QHOMc/A
dKDkzsvvr/cOWTP19qDkWeDswaJpROgs8TDpCLeLF+J9KhO+zgYiohxV91JkhS+W
M81IOjjFPJK8Iv52PzRae6ny/n7nbxIjkraLqrOLNGPnTevreD5fiA/F+S4TrB0/
O2zT7tmjbT6trJyfMEVVj1CtIuORUsM/qRC+rKnS0J8tk1kmvS/OEbwiOCIzgXcv
AU2jusI6izVxX3M3tzijQk7FG8b7xsuDblc9QcJJsmUxwIAxS0nJO1Q8MuQ2Bw39
Uk3uLJF9pQ2sZ11TuE7X304Cnzhbvn9WMV4dphPjx9+i9DOUiLwvvSLX88HD4Tuo
qE5zEDXeH8JDcKyyz1B4P0SC94SrepnB82B0AlNcxhR12G29ap+QyJIMtcIZX76e
9mS3EjCjxSKvzeb8uMT3rQ2TH1Q2alOBpP16C745gmQhHDRzY7RAt0gVKd7Ic9tl
t4whRDNks9ABbryjFQ+HA4tpHTch8rTvDqmk2Ftv5/1qnQfQUn9TyNbPFy75erSO
F91OsvDz/FGc0Msezj6M8IPreEasaQQ5KRGz3/DnErU+cS72wa8r7L5+PQocPRta
lATjCICBLN1DkZCz3m+1beUHUx2PHSzlFU1x71mN4eqJIW70so5FJVrtbnEvRysl
T7x08tSpBe90rjk7IEqtYsxFgcYUvzlmpSEjeNlfaxW0/8TbllHqt+oDEOQTvePf
QIpt9q7pgltuZUzTAoLFSiMxh1+gcMwpTvWL5CYKgDFK9FEOoLnwQyp91X51sh1k
RSeKwVJFMJcTa/tO2tC1fBAfJD8BTXCjeAuYMNnLbMGk24+ODS5B7R7lbFJeP6xp
NLOI7DXf6tzWLLSPSUkFuzKcTFWAUKypH+wTQ6K0+IoagvTM4FQlatFmbcVDpdXN
qRSvg2TpOMZhUwSZ5lvJ9LPQdiIGyaqPIC8c1rViN/ExfOnFE+NVL1+KrgT/n1P7
J+aErBT/JA36zvbD+3RDrlSGYb5/ZF9jdZRa+yRipNDZ8thizRyEcdrEGoc3VE3o
SZzl1dhCK3JSiiaK3t6URhYo9GFAbzby3EhZ9cPqAOsbMnExMqePfsm83ALUXv8v
FC/6kOAW/3kt0kQ0yxfkJ3cxVDDTJc1pYfxfRcpfE1BcJ0+waBOHOsx1Md1ytR9Q
QNbI0Pec939pjcWLYPdNDAeadA3o8+XWxZQtowxaQ1RsrnDJ7i7/JLp9q4+6Os/a
w3CMVUroJJdEx8WerdHkkFF+gnT14n7N44jAQm59z/othsYaI/G39mI8J7HKhk8H
OTZ3ppLNzKoJmRgMyBBnUs+7ptbGOE/qhnvQ3L8evih9EBgpbyQ/nBYMcVM2+mg8
27ZtiRsT9B2C8MhPfY2P5R9qQWeqb4s5KdRJFdTQy7IhDwFm7OLPibtjeNy0Zb4j
RiA2+FHZtvpkdd2kG6dq8qtEaSVYNHacRQxIYPGpr0Rot4r+Qf+1Kf2eH6fakM3+
44IorZY1yvXe3AyvRpS6amENfG5zfPZedk/oC6vGy5dsD1xKMWAGmYzV56jbaIWu
Xfk21kxQNkxO0aaauu5XZzBeHNwqqwRCMeo9r4AgymblLY/z/IBgRhVn9dojzH7J
AcqhBvLgW7K2SVQzEqK4DGKUsImKnTnuKShfuTvTdLh1I0dY/qN9BVBK8cBQswTs
A0GI9DZEXl/sJTMp0JfeaUw/05EuHBZI7Cb7cZzvTTtCY5WDXjQsB4uWl2RoLC/3
jdrQqlKhZcOkWALzsj6vv3Rw8ETUbgvRKwRatKHJKOP5mX594eFVC1UtvAooEom2
oYZiXq928Gac9fUT0Hor+ai6NRn7/zLNR8ldcuQ25G2QSSYe2J605jFmkZs+zUza
UzkJSQBuYbQC/XWYJ/ISXS1z+k4C52ZeoUavpCfRezNzYJfPeDZRJ0g1DEGfnYEy
rFhcsg18xC21+FC9nY5tsD1ipuKZbq0n4Wc6hyVuNBwQGNxp6gNJydlpMOEVkGo6
lee/DMSNzkS3ab6Gbu0ZZDfOcK1Qb24c8OX687YqdHPxmmv3a8jNJkmRsObjGtxv
YwxeO9PS6huMB79mBX7kN3TgMVNp5O6OYUzwZhNsliSrNTbQCvJitr/5Hcm2Qmt7
NEwOBe6bsZKBmbclKBTL4sWMWRMLE89E33y8Cz8GvLcAKSVMbiW9iJE5gbd2h1Ts
8N816uveqgb4/HdNT+p0RI5yYo8fZd/15gNubjN8sHEu8U7RcJCL931gb8rcz2b2
PwCyZsIhEaXTG62HqkVK1a5fZEa1INWydSLlyHGw8KCSs9A+8YZF7CTP818bkj8u
CcQo+ulZ8awoRo9bx4h6oJ4uSxQ9dQVEh9xs3DK/yPzxtkZO3Ffgg/lPQlVSGvOz
ObModcKf9lanWlhgbgXcezRqHS6t9D6OQmHXfEAkkmWaQfDgbGs1cPoSm4XWNY/V
oFXSccnSIhBnTUD+VJ1kpAZ87ml7URaAWjayqIEB9AHOwzetxlRipjU1G9PVnavO
sYVPahxc6lU5P20ZHZGQmnk39IGfaS0IAU45zjKLNGi6KBZodxKO31MJR3Vfu1ul
9eNUnXaGDs0kFLokMHzyvG1A6JujeeAKNB6WhTamyYTCiJ8XGjxoo37S6JSN97WT
KxQpQik3VqM1IrVVT9vZUIaSavYx9mAZUaFLziq1fcgIR8u2NcCM9zNCp9s/9Ewf
JQxr9n45t84myWea0fFATR0HsqXR6Aw6GHvR72TRbuhp5w+OVFjF115Inal2+BG+
pNi1fBk4/ArZEyjqVDW+iGEryAW2Rblw3/Txlpul5a05jRe6Y2B3kb4NdUac9aeD
NntN3UFXJCbnNV8KDG4cl5cKm1PwM0Q0D5h8ilTw/7lAs9kakAzTHS8bHPzyK7Fb
tmAANAb4NHQmeuaw5j5X3mmKBdsRzaZwTrndg+VTIJdst2ZPfjtQkx3aZ4+91Kz0
T8mQ1gmTawDtIqNH4I/DLeLIAT5wweWoXzu+Ufc9gGVAYJeIWyJvsurKSQVw7o00
YVy3nIp2sk6lT7rMpaO7GbLtMXU6rI0Sew9KvKaNOaCsSYaKhdWEHUmzbe9Dgpps
Dsi0PhZjwYHjEHhX3uG9C7+Be3ya7qwJhBT5OvjOdc0PB4NyxkkRyDmB+FKz4eEs
+Z9KoJK5XbWaCMytBj+TYkI9lzE2cag46VQtnY467WjtN4Vsb8FMnQkwKZbPUpHc
DTSwOM61tTylU635s6I/lhEDF1zK1yO0uiSLaVvcF4Ef7LdSUqVOsCloAefAHu+6
NMQfc1YvQsPB2Ml8/dTOmRqHlUAexEg03xx2EEHhGb7RSsKom6iSspJ2beTgOuRO
Vwebfl0j6msrjl5QWl87lJ3dDoUpleEr+ROPOa3G4vrqwllY2ihv6gDGL9xo9/Go
Y523XnVGCqAXnlUQjoIt8uw+1NN1kUT0gs2agMrVx8jIn1KUjATVlZiUKlQdOjAm
088K+9kN22ri5UT6gs1nZjQcDtz9IQ0AEaJziDyfiCjS+8nHy/pVsme/RbvM0/OW
K1sit27Hjd/Jq/wIMyLtkSTTj3ev7AYQe9uHRhvWie3vPBYqxzrrBN37BVcIalWA
kb2sRMPGlA63p35J7tNodNCAZmwkD2lwbo927qXUscTDxMDhspfvIaVT//qc6ZLG
YyrJ23HmtvWxCEdv+toX1xKvPVQAYyd2LrD0+dxcDT2LoTPATR9Q/2PrIxlRJDJ9
zsBJnWfEQOpkHKI1P8xUuZUuhcx8Eyi51nqpKvo2/eJQVw3r7GEg6sjo8rzNxH90
rwX2JxBquVG/92b6EhDjfmVW6ucN+2qMHw/5kgDG6OXVzY98MOuHhzZU1w7bTJaB
Xo/OA0LbV3vh3ZMkAbK9sJLRHEitRadC7FzxzlmhYDMtEx8QCdLZZzUm1jiKI4Mt
csOvHq1xzjkhkyL6xcoPuQpjuBSykFwJ4iB4sWToNmXGNMXGjyvXy61td11FUEOn
P4c2XWrzxMhj3niXGpWihSDd8NGYlzkcmGsp3zVMFaTvxigCY/ny2xcbvotVCTMT
yWILvX0f3KJ9+uSkVCpGUx3vyv7ygU2DXcSQpXoERVzWSQ4Rh4ObZL9YUtzWJFFc
2uc+mNX7c3sPAMy6gRxDK9hLtyCWz61umRelLsQxqs/o8OVWmRbXH0wIR78wQwf7
E0dHLMtqjV7PjG2R74F+U/Ux5gRi4Fj3udK5xawK4M8hc8L5PYBJN98zan3K4Avt
NKel1G61B9Tyf/kWMmtRKE8VdCB03DTvuj4J+1Idk8qce92pP659WwEuTfYMGT5d
5UyfA2JZEBNX5mZQ2HFh370UWJSQs8m8vKz1nJE1gE8ia17WVDtC/MTTIEidim/B
QT+R22odXMzts8+504qCdLjVRKP8jwBEvs7F/nGEqAaFdKXllowNYKGvB8Ya9AKM
2XndRFP2nEzD3gDDOWwwFxm/2tQOCjnenaX5f61l+1B0syJwwEJla4SqHyqhDKl3
IAMvZLnwG6e27Ptw2jg3W6XFsKRlJe2zYHHfIhGqI4PD+bOODFKi0Zc84uj+3cwU
7pbtioD7f69o2rugkbyNR66E2V9s+RdKs1g7MSL3f/YzwoHGcXa8hKq6ZhdHDqAh
Xf2eIDZOEDQcwbiW/ZWWZ/0mDHh2wzVsL+dyRb1v1hbnvMyNNZMoYDLkpjPLrsEa
n3eT2OMiV2WIa9JoVgCLyIOm8k5xWHaeG9diVS35WHMxhkTjk31lpFuqc0PKe7wL
oEKfL02Ki0z1JiN8Wmwvb2gQUbiKznpW5SJaZ9oWL1U7VrGEWcpifvYlONvIL7OK
yIYuZmjYVaaZS/Rhk8JbdYS0JMD262bGyRu7BbJgBN8pDLJ0Lza5M3eTH/YLYN4e
jVHemrgkl7kzyt+u78efYBiWLTgVcJWtPjMR7JZNFW/AAIyZLFiriSTqt4Cldd4d
u5xpVG2yLGcjBnF/1sltrVO+i8OVXSlwJ+y6IhJVJAbcEwH+Ix7r+1fR00qw35TO
RPznbNsareH5NbAVHbZTHP/DTd2awHyDRAtUFv8Q38AJv2DAGG9b9DAz5Ac+Zwl2
cLV+UPmNqauNzDajH6iFD84owoM6rsTu66AFpQ/XVpK1ddwk5ATD/sdhUHHdRb5G
NJsq74GwDvg9Bjm50eEWhShY2SSbosKLFhmA9HqiSK05YdaYK2kJGNTb6ZrvXtEp
yD/NCf/NWZLC+Zv5eDeOF/LQKWwof0dKqe/HtcE7Jk1/AUDfYsYmEPCqUWzvIPSs
oOo5IYIaW+VcIZiG3bP6FA9BZfqAMLy8SpRm7wrlyhlEI2XQvfOBp60vICqPrgzD
Tkvt0r6wA1/LLWNjWdFK/2mKI4GxZdaMVSVHQghl0a7+KOE7xz6vVUDEQrYajmx5
pExNT1fEVp9++Cx2NKoYEC+C3ZYpnxNU57dAhclcQ0o1js+in+8ymxo2QQpK1SQL
9DPaIEBhLX/y2z/mQ2522zHaczNJ44WBZDRG8gBPWFUrQA4mIzaD8kp3t+OROtGy
mbWWR42VIWZvZq9sVwBfY5Bm1ZKqGiL7+VKZ6doLg50GeGMzFN1W2YUrEE4xXjJ2
A9QaQaICp63NmCrCgWI+8gpBwV02aUFCF2KEDX0+XM5EEkJ5+ij3ooLiy3xrh5N6
8ymz15v4uMzWGbH9IDSPgwWvJaXVP4kKZg2H3iPf1rJwB89cTyVXMbr5AV4oyLyl
AJfusXgaEmmLvda1GyQemSNsHNRiNk+znQtbONRxQjw9ZcMLMnmaneGJWv830Ja+
RejOEKsscEhM0rB6noq83AnDY6AKKjpBZK9h+/PJ/3jUtxOPQKJwiMJdLEOK07do
QpER4prEBcFRdIfY9EMtwhOw4HHmwW/qJkuxaEi/EVL5PFMzy/dmYGKUgbets4ZM
5r2zCcZ0g0g12xav89iTpMUMF4rW+HHF7XYhHdWcj8pWVufJK9m6/Y8QXThNBpBV
XNxeGHlyxyohxXnzDu1FjVPXVl6cdYX9tDX5/C2hP/xZqpFY5dYVOoBJctCcxHdQ
NLANOOeosnSPcupr+7U68nCdEmzWPf6GV5GlSWSZ8nA/0aKQ1s+bqX0paTGMU66s
dILg4Aw7U1/DdiAEUspPQwntGSWphuO3E/MGzTC54LwD6W6OczLo+DGhHT1tWiWI
qqO24LmjksbbhVWC6GmcADKFQ6b3khUT5C4KZYWQDmf54dZOvfIVp4Hro8FuJF7W
rmX9zw/1dn94VOMOTw0x9uMcQVbzLoVnj93dnvskbCrlOaHi8SAig4nJaMXtVWwO
3MfmJRZEdtK1YnxBPNNCM7pBRoYTQyHziR/1QlL0zgUDX0xl5a51nVTWZ8CLfBj5
pw4yR4JcJ+WZXFObuFf4YsMMqbAkzhOizt1Q8CGO9FgDih6kRWg6H83hi1ouzf9i
r8nibWkhGKEuTDE6hbEiuJ/tCyeXTrKu4Cl5AqMNmKaODMT43NMisDFRuebO8L7Z
lU1ogKqXfVScul8deEPJYcH1+ONjQCg9R7e8grzDf71jk1uVLWO33AVXPTQbhm4H
oOAaYJ8AjBS2n3aTDAa9ejw9/qWpKZuI0mt4mg9ez3YeF3V1/XBpojIHVl9ZqPFn
D2HGT0ckmgbLfws6rrOmXemCs1M48pCdY5Fp+z37PVE8l68exRoEpwIWCnzZYODF
07nI7JVbe59k1VDwksOtqkDKq4QphryRtcDroRiFSZuyf5vS+F+1xSy/TUdW93vQ
9RFhzE3trd8BPTZLzEX/Oe30i2oHH04rfkoeL0QnMbSmQrbmKsAP0cMMm+j4kr10
o0QGvEMRJd0MCQy2smewqK+TPN42ZosCDCWKN1xru1bdQrr5n41W1Bl+qFKzTq1D
BqXaMUsV4Fj/mKijmiz48jq1xlW6JT9TaE6FSlWBsEa3RoK0lE5pMcG6JMiPkY+c
2nLjL4wcH3/jYyXsaOjXOcA5cfai82VhFQQVuECCNYFg1PUMV2iBI7B5DJuYtU73
R/R14h75Xq3Ms7nB0gsnJZSewaudGrKG+zXziCfNvpCTq/2mMqxhtRBlfmTJyT/0
we14U9BJgksNwxylw+FsihMup1kkjff+bS1CMsFj6mZnWcCGW9KkC/mN9GkjXT9y
H8K3reYfoA+qQJmknLpwDFX45gY4z5RqumqrXdtW/dgjLyv/DejHW/xBJJKN6dMU
Qazr2qlLGtwTMzab+n7AvOgAyQWqFJH6VwblKallrlj3nSy8me33LR4VbxFZn00q
XHoRDQIHmxFRcCN0X3KoDCtMOvuxVkHkGiDFNz3SihUYBc1j+/JxUeOc7qx0ThB4
1dWVQp9En6kHBsTl2lMcIPK+t/kDudugGuv52uVsazTSqQnLh0i4x2ZJWu7fc/Wd
DafuNACRjS/1YqaoJrehMhllXAisC1glbs7elIO55gYEeV4Plka/BL0aTjzlnDy7
D5MBdftSkLUg1nfy7oZuUS5UoMrav6YBDPwzXi1Ujax0ThyPKwsvOpfkJ7LmTqdB
ohUGNnU1Gc2C+T4pZmCqJprOBcLLZu3IpRF19tNoOQ6GwjOEZ6SjySNvIve9jyG4
NgZ6Dmj5iN6MpLhww3qTJzZMfCesmjkk5MCvN0o3HL1ofn+kd81+4P/CNxeTuNR2
qtGPq+PYE6+K6elSD3KMMD5hEPd/uK+6FBDWoISF/2lbX1QZzoMB1Jw+foZesEAQ
4hy2FlWIKxgRbIB+Jr/hYOj10rvuxw5Pk3nwTy58X4ttXyaWfo/QuGqOTp8nq71H
WC4Vt2sQL8SD4nl/6SPnlwoXhHHIBJ6fs2vOSBcDpsihETdGfGoPgUd8FL+JwRwC
N/V9bN5NVeB1Mp2KbKlr6tWQ3fqwPMWKRItGTqW1306fRBeiAjrsyEvCiSvJ8tet
DgQq3PTnEhCm2ZxKGvyqmjQXdO/j5qCBV5QebZI2M4kLpQ4RfSjH2OMSv7dS4Svk
Vni0LSY3valsHcLhSqnlNWbkHedlysHOwrCWVtz2Ke2Nud2nEhJBm2+E/oSACkUz
wHPwU+Ij38fWpUBrW9ge6GxBOgV/gfwXnWMsuT7KBWzz67mqKygXXXQHVWeG0i1J
MLuLQgX8Net7HSYfRxkCgqVah3GrRFy0zZVMQlTg1nNVCHfMnbkQSP+Ni6MfmPTj
LGC6E+ntCtIib2RBd7K66qJJRfRaFEut/gXxBjzWeSUZ6hW3b/ELwTJv2qUaQUfO
SRhv78EMNyNcqVlC4jODKS34aN0PMQGHPMQJJDOM6DBbrbZo9tZr/6NGMJtqR1ZN
u+b1Jm3mbIQoqhB/2okYKVF2PTQyM/W3Nc8amh+BT4TFdV+hexBspDG5zpdQXaHg
GfORTlmVvreagzLpmksXufiJUcsZbOlthz40pCmNPHD9XKcT5ikkRo/X6eYJRl1S
vTOViHTVD0OcAYiL8VBfp8BVO2ehQR1tK9axmz1+CN0DeZjk354oHjjvbcwe6swL
Wo/tPXwu9V5Lvh9hoEeiP4/eRZaZ6DXCz9iQqRLZZbt6k6DydMMvXv5l4O7WqByp
Ck3yJlZeDFV3DUnJAIPpiwtsoManqHMLJC/L+rCq0mmWFUd369e9O08vUjsZmdWU
jmNO7cIzbM5s1TVH/U7z/QuCGlUxjJzta9FPOLWGr1bdJ1rceLjhzzxUfeJqnNIY
u1TY+p9lZVRQOhggGq7rb30VweK/1wqZo4ZSbeKzBnmbPaWa+ZcN63wQkfiof37a
69Tn0dHCzIOoYdnu3IPDBrur7qLKDOYDnNFFZfgtPm2vCVTCUAMedTDT2pdcveP/
jjzkcKhCXTg4fVfekpMvQ3YzbTdqKpT232osZTEfoz17F3vOXYzaYG9PlSvKL9NA
5kt0rVx4NhsP0J8/2/74C5gMHlqVel4UebXBdq1w/Mmh56ZfEDpp5PeADoUQNVaY
6F7x27oJ8vCrF+spezZPQuwLkXdN61hFs6xgXD5MMYrnRsvXYbsM6kPBA/ntpLhL
SRgTVmGOiA9IvINr7fHCbVTMC8UX+6rDLRZabLwrnpgDRtjW+Ix2zyxPmq4Pcr+w
TdDZ+t4qNWG02CElqBgkae4fyfP6E1gOt1rOHEoHKIHGE+q2aWPOcjmGDcCFS+X6
MgCX+VLjrez9avsUIXlmqisWELqtmoieWT7Yrw+NG7+yLWukUH266FvdIgV39phZ
Wty2hzZBKQ7uJ4PMY+O6ww2tQdxUai0JmntytyjX8DVMeFRXGUq9S4UMTGek+6UK
0x08stZvzCz7nQpM9z1wOmt5V1wDSxbQFs0uWTLCqNWoXthFQivUIhPWV9/nMSPG
CeyLgXCRf7j/IbzVzD4Ul67HAOu/OpDxAdCpdDMBORQWa45sM2N3mDq/2t/GhSTy
WqYXcha5IcR9HYqKNv3moJVXGMZKdTC9vS+3BjY2o597WjYPbdSwDU6rj41H/+P4
WcMV/rcWlerPKrcg1y5/taK4oEH5W5XUaogaEZJxbbGBFwp0WcYRCFxJUjrNfPnI
+N93pJrMrPZzJ3SLEcihwHdkIuzS8PceNReGMKQUWdPh8Ngr4yyxUK5A3/qQDK5y
P0pM9cESQQvrTmN9wpGbamPldw1vra1W5bHZj5fj6q6F+f7GxTTg343/Q49EIE1e
MaJvVBXqvtuN0/r9w3l+SFLInPdYJ4iqhbgcZ5bcUTGoXCJMj3wtFnbAS2u2p59r
pmr7wRLi/M173FCr1ILp4pF8VMVls1f/nxwN/jce2ayz2lOvzm++22W4PSPrJgSZ
61uK0JlN2Zd4E2jF5I7W0n4kHK5lSklDhTec10XzM+V0lOsua0IyJhTc6Un/tINP
ys/BKDWsrI2biIp8H0d8M5nxOkMTsZHjo3RuL6ZHEx+OuIzsgCJL6PD94wpVHTYP
qvAX7bBIZcWAih4LiysBosKtQ9gX+MIGRmBb8TTY6bO9mhiB1Mw6OIWI+yXzppjt
232um+NFXF9pigL+pf3UhGXE9gkGTa3+9OhKOzKjfgYGh6O763KIvilamkQpAoix
2qImcIwR9F238Oznhata00q7qP7Q9XbGO8tHUrvXp5sU4dRIeLN82lON8pvp48HQ
n3xJGQpYsBk348u6Zd/K7WBcn1sfgD3NXZmymLdqukmyWjz5IxuYfPRrhyEIUOJw
RDrJeRRxZrniMIMEiXIRN/CK/7Yzr8bLKvjNiEZKQPlXVlJRPu18vMd7R+RxozWE
o/Ua7pmrnax9kYVTomkk3wkY/eeghe/gaHGv/x/U4vEoEYUrBjV/L2z2t3heoAM3
tGCM57lYMlfBuq+05Muaj20H8SKQCUcQYIrMoQPhUZXDTfW9lUPfaBr88KCJcXwk
qD8vcbzqdfvQ8C/gTaT++tjZcLgoMH4Pt5ACicKhjiMpeePXw0q6JZJ0yJg5niz5
cx3JrMphy0/ho0MQ6bNOhRlmlQJ7Cu9VuiRykon/RHh3Jrmq5RE7G9SONrR3HlJx
6Q4rsYueCPFG5Flvwosvnvd2n/OdlECB/eMxepksdL/mUgjGxKGLS22PNmCMxood
duYImRsYqjnCQsEB4EKryCodqeaOHO2qn2fw7SmrU+DnHqt1wEpwoXmduRkNkFOU
GKC4dudmH330VN041HfDv1gtn2U1cKC2sdBYI5HrogogktfGB+kKoC/3LjwjFM8h
ExuhTmG12QzGRdce6auKAAbODHeZVjAYrh5XPbPbjc6YIunsE7r6CdUQG/XRJee6
pr3qKxWcUpWYrKV1z6dDR1BhwJ82d4tYFFp0YzGZbcAhF/v6xyXpi7awA06VyWtR
WGdYyThSfD0phEXjvXi1EVwnqGgiRQmGc5eZf9Z46DdECefb7Iaa2UuqYqrVrv1b
9wXFhgpebxuOQxqTIvBgQNVJaAAwQEQPFA99x695XIwy/EB4sr+V4ksTjzfmS+oN
LMbID+hCadj/iizK2LXl1B7BjzKmkn/68QtsLhIFuuAgPFIkVEB/fiS0yUiszLaS
0j7wjESBjm5V/JCCxC+S0+hbIYDmdEK7n1ZgxuToeK4R3O6dzU1gP7eMEZelPXK2
C8Fy/C/tUBjMR/fuj4qbj/w6iUdenz7+IW0FY3TUfg1cjuaxqXaPAZjLqwG3srrC
zORGU3kVLuCC3zhysO6fEBvPxIGTxeFbsfllSiPq33gwMvkq7IYa2rhZYTLAgro7
/NL51EYx5JD21KdhVTdqSThWe5hbw4jbGfmUHR9OSsmHm3wa50vbQVpZvMXJb6Bz
Q2FwtwPwUVhXcCaJgE5m/VdXt8vxyt5B0HZ8PVkfCRaIBo+eC79nYhYXqYda4VbD
0n5h0YNVDgCvUp0//rimi2fr6VsjM4SSVHwlXkVLUR5+6d+3BZzFX1fjTcNFRRjd
x8HsKf61Ao9Jm6+OPDrW3GA+u8ICcqKiBQ5uDnMda97W2dZ7E87GRxTZxFOt78iv
/Fr50spwlQM2qFRAK78Vmj1r1jwUDSjeCevyf0nRo0MWsKOEEno2Tiszatr/ac8s
IraCd7QIspfisS093kmq03IU3D/AzZAx27T23YmH1fd1q9Mv4DxhjP5SuTS1zzku
tDo+ueY44epqpFj2oJACy96MQ3L3eq4mBXt5aiwZQlP4UIemKS7eEhmgx8AytOYp
LCw0qG+w04r2LwdYxWPA4hWH+9n8YmRfHsXrdlFPr3UI+JuuaiFXD8nea4ZFcR6k
ISNnsE3ya3X4M5ylVuXagEp2+Mv7raJ4ZsGUdG2HD73alYjLxfRq9u6I8yZFrAPu
bRAh+Z1eRnYPEsvr7e80E3ZYKXnbR4KKh6yiK0anbqXcSZXY+xreeofyVa3smsvi
csNsd/0+gQg9oU+uHrFLnRLT9CjMNwNc0Ooc1VJ6TUlUN02YfBnPcffxlK8xtIL2
1yLql3AG5cp9ZouYpyFcMZGUaI0D5CsVFlU9Xe2y+WGd2mFSouM79jOMlzbYBUuB
0hxKGHA7HkmycGMBvoBYJjuWuY4rjbVhI0T/61fwTW7gEqiCNYo4ZkmTWigFDxuZ
b90j+3NaIvLXx1puw927184vD9jpzDOERkQx/I3WCflzHKOwOL4qwiUWI+JFy7sy
bpDU1OlbYneyZQOynPV6efh2fnk6N2QggcM/pgHYIkR2M+g174D4SuTsY1uMySkB
HcY6D0Tyly7aO/fwCAkPs0uDboMErP0Q2AGBGnsWAJL3D5RkFWCayK0+oMZltHDR
V3uNjrPi1szXzr2qYIv2557AY/3mfkRgi+WZM8FtWWlXppCvnJS1/G510/DDW7m1
aQir8Cg3mUGD7Kk4uaP3Be1w57XQeSQU5D+RpmQ6U97bytymzW0CkIxYt8IkJAI3
p/awwPZ0cX5U8xMWaZFMNR1z5RO7zBb/mYRSJlToavAQGXj5Yjve34BBttsdzKG3
9thi0oAXTb6E70Ou/foIdUX7yUf5zCFuIu4xBYBzdsdmCyW1ddXWeZuXbcqws2vy
ZkXg52ZFPC6gAP2OBVp7mPgThI2BNjXWpCTX5Y3ivTST0G4Q1ucr69GntlAs5uyA
d8DpRME0NfEA1tJofC70MwDB9NAMt5YN5sKlEt452NGKX4OXnE5b0sPIU0jIKMBD
TLAvRFn47hrNcLA9xRyvyPBPGMiiPzUvSsbzGZCNfxyh/qf8wz7JjtDdcWmKsZB0
6FBA/FWK3oV9ec/638Kc0yFQp1dHCDSd+KxXrA3nuWBHCuE3cZhmmXnMllSZ1T5Z
yWypR8g/lGrhuxF0SqX9Cu8xUnCK1/GpSJvt3l3/2WKuSmptGWf4rUfV/avmpMoQ
TX/l/C17c2dn4qGtwG4Y0rh+1iAPWjKQBvzaQYvjcuEFqKRt+w2jbXuiDjYkSdRY
a1SCwaVzzpTMTm795Tnzjiq4cy/TGlxwn25WopjutJzlXVShgjQpdG/atnQXdjnt
CE5FJisq9cD3YMGPovZvxMacfAx/Qohq/lCV0hzYrMoXfwxwhPs0lDlUqnMbhaM2
du/w8hyZyCV1WFBoFD0FNU1XuJNGkAGK+3DIJ2an5BA0YdLnmrTmfFNUCOLWP8Us
RzkE2/+Lw/NQ2HuWLQs3/fBbXQKgnkYEIyQW/wz9N1YQ9AOEMseLXhCl2lT5E8Tu
cFOHh8s/kXqHGB246NxCxceQVN9ps39LxmPscIRYo3rG9tKqmElSa6gAMXu2USeH
fuyoh0ncA7kA373Zw02NiKCVeEc+MJ8DgSJzVvSP2eRuXQY6wl3euY0mH7n3tjt8
SmtsD1cjvVS+R7bxBOvyhLo45mLMyl7I8mSZQdWSIKcBP278bC9TVmJRTsbirLpo
/pSJeNnjr+9h1PzNvcnfk6elCeLdj5LrQK/zdVPHVq31s/Tuom7TAVHKZEaYMAiD
gnwtDmDv4nXEnfSDDD05lNl/wAeRz8CuD2+Ej22jSRmlD0zPRTxEtMO+gd5psu9Y
nBPt/0JtFMdBVg6FDLqkbTPT6cinuuT4L3oUcGT0HzOBuJOnRBiQhHTmKJky0b8l
o+JLf9q/uaZvacOEyH7puzB6p9VZpZwljdPDNfW75jFzyogpyHhtKlPq5/UYOXeu
X6UzK90KsaKsW9NlSdSRXxA9x74Dk0WU7iQwdAtm/VnEoU40C7TQBQvM0nnI3lQC
PEKoSzY8+8meDo5JUwExDqTuDqSH7XFN4Guqv14ydKSNWIFoGOLjjZIAtZNhHnvU
G30Ps/bbiSF0KMZeSqJEHdLRvJjV8gxix7ejQ2Jgaxj2cxoCiJ34savhLECkNTT3
TZxSR4i4mTeBSCRCXGrXujNTd/zeEbzIYdAxROoAabIDNxbpWd3YFbROY9SwEgrq
8y+lGi2HqHEkjkm4fYE7Ssi0lh8drTW56+rL61S8ms5TS/17xXcDpIDJFH16OmlH
IZkxzmvjuvh9LX2bfTMxZylMNAuFIavBVxKXC+6z2pY7jOFPDqsMeqznpbJgbDOS
CTeTe+tLWFRsa1Hq5CN+PwCzt+l7fESEZfkX37Ix6n3XNjCrbih26VFY1Ij76ffC
kQSg1ATI1F9NF7bk+aIFUXY+VSzhdLo/mX5Ihc6B2AdPL75KTEKzhBAbT8NgI7AH
cwG/bpIqW0XTysIiG2MH2GMrszhlR0fGf7MV3vVwK2afzfSUAvRz2k60k+OVIATN
WV8wnrhq63+9tYNW4UhkRM8H0m/iFj6d0azcLefJjI4bUMA4sk+zePyd0ZtIKGtP
nyxRIFtr+ofAWcPOoomCIJ+J6O+ywh3VSnj8l4mt3vkO4gmJ/vV9aeIwsldGctZp
M9nQorljuXTi2AdWh5Aq8sfeH6inceHHRNv/wQeOAnGeF+rddpHQ+zYxWHmM397D
SQ7lLXyFKjfDfaprmlsbp1hQA/gf0KTkSgg/4y1Q2tj4DnSVheZsBwLQdLJXQcRD
rF2em9j836W6PIPyOyv4dFXeSEVZkoA/iKMaofuZSAzatfARNsJtTobOjren/hdc
j/6FzyAtbPN+9EwPvnJ1NYaEGMYS6YOQ8fqtjUczOojax0iZtBq+U6HG2tAXhF49
6YByZaYSkQeHVB2Vj6qfPrJh+jhxmrynrpHBu9uxeVUgmblwhBQUsliNeGzCiK/r
XSEUZdqCZIH9lFnC0E/ahlHyjZJXYw8lPMYd1cc9G0YPVFRYdizUslkLdqz3GK71
GvB38woDHJgd11N2wQKBGPc8/Ar1eCEgVsVm/Nlja6Gy3Sjd2xZILdDZGuh+jV4V
JJE5yRh1tpZ8QjiBEcMh1xL1Ix+ELCK77cEdjeyCLTAGyBI5M0K0iEuUdMmqmpc+
BPSOq8w2PTXQ9hO9z0gD3DL9Ei3BxfMtBBAznxcFiHr2Uwq5nge/JbNTnuCk0Svy
HoDUjLoPxhNIAa76E16ww02xOrNp2n8bLfKsnkYIDtVSFQrSVX0+GBHlQAc0h9sL
3tUD8SJZWOtMldDATwPa3LR3mRK9sdQTUcHAlFtCoqkwxNGPJ9Y5lU+qDTUciuHz
bUpBQgM7YmQ6uimx2zkaeg81MGFAS4B+D8iJAxgyUzZvMdL6i3KxNzUpnn60Apm2
ww1QwtQvtbNQ2QtTYQ41XbkhcYgffB2Zj90pGlhnNDpO94bjb/MzhpBniYfaCXEA
VAliAjzL6+JuztXVadUXzXDJ+2CfZuAYeu9WafNiwUztAkcQQd4B/j9RB1VWxQ+1
K7uYiUsLbdS2PvS/If3irTHo4erxcOmQJAnG+rOFmRRLGHin/SiMRXScqk2ZFd1K
X4A9PRvUhbGg4gffPes1Ab0Te+cZvria1zrI8/6NQ7YeWypkUSkyMmPczOJTovk4
wIV5e6FmGlialJYGWpSaNVSEbJatu0Dnq2WT94+mr74Lo+gxq1sQdwqx8boL/Q1P
5wfNPmPStzd0/cZu7nczbqWi1ZWy9poiLkqvbWCCRznGTwUlI1EV59uxy+rbzoCA
GeqpIchOhhMNISt0fO70OCQfmKoMimQf3FnbSOe20v/4eC9x0mlb6Hs43cYHxUwe
FBfBkjJNppEmaHq8o9z5aVgYckBYqvuzwZSqOnOBv3WRztY6ZwQptLWnXnhmbC4S
ZkpuMH1ZQkSvdkzNPMCmid/2sB4ml6uJ1U0ozRdTv3Iv+AvaHGd2RbDLrsAEsTEX
OIfKBDt023++WCqUm7xgww2GVGAKVsOkz40oB2a2EcjzZXyKca9Kp3yBXfWuKX1a
gitqR2zDFdmpuR7EM/l8CuLV3LTZotiWBJAqRs/eH9o2uiN+SlQ0HGeqy0lgrI7s
PQ0ZuPU78Fyo13S5jABRqylHZqhJtdXqtKtrPv5kCGhWvwlUsNc+rctwapYjKisf
YI8vZUnMHrqo5gNP0/r46lu4vPpQhctBayPyVMBn4FO/jj80dHht75PBH1Oytijl
IxLu7Gp3sKlNqLDrbq4tHQ23a9u/gcmgUxQVbItEdzidFR4PPGFlE5L2Ggr4Yf/c
odtncR1irqTgpdZZ2w95r+PKiyx99bDhb6t2725IGoPDeyYNx+YvtN1uzLniutOg
mm0hh2ZzDL/oCSo7aEArfVe+gaCW0yRZ7zEDjmAS746Ff5TPMs+M+ArA7X27QONL
yXg024xnDyeVeav7XQCDAwt5vclcZIguon1fk2KRUVdnOoOu9SE+H8ybZ0e6NSPz
Xln8gubP1yzK4ROLfLxrLnl2UnH0L80jmo0UfDwJgpsb/xejPtCwwN0kEudcYEHZ
8/9H8Lm5jBgx63wBX5Vwpul4qnEgWpGQIBl6XVxGUFpt4CIu21fPsNH9bYPEqW6h
1xBYCqbZNCVFjr1f26teZ/iZNq8AHjaORCRVMBpPna570GzS+bPWva3nuB+M0uzo
/tMx5jN6QSxW/tIr2OtYQ2q5MZ2iuwYfz8vLnHcVTPv2FZXf5QX4MkjPk/JkAU8x
PSCwwFcXPytBuobnVssTdA2sdbHXbIIIoEike0q2s6kAm3g6XsENADUYmaI2LN71
9xb9SFBQybVEJc0Z3golYYkA4+RmPCAIT9BavLu+rLMBqBtpLj/pG3MtWanF6dCG
TYdcuarLb9ipndbxaFjcahRPu7LfK5GmqAaPZmYekQODE+MQzdUzHpGs9KyZxKOF
VvUxcFWPebbe86L7ytXhhQKDD51QfQwGPKAsZs8u27M55uQFuW/qs/f5DbDaTAeQ
hOTX0v7KjOUSHOV7w2Z1LrUvHUsAnUMfg0zjMozuv8PvTnE2GDybAV5HDjnI2Jtd
kcMlnLLHV1z6NOv7h//q0MVYytYheG0/N+wi5whVlOYS/GZ9oi4ECvBz77JMKE+4
rjnNoHY8/q7IYWzXBo60M/teu0SNH/UgvVDOd6w69hMvsURuiJkmLhKjEpl6UQfa
gyCiK3rqUO0fkp5snUWr2L3aBuwzKJ6fWwI0EB6mXuRygyBosb8wxXTW/VgvZvWr
VlRdfjrB7wJjuD8w14j3YZwYUAx+D4Tc0EydiLKoz3ulOfDlQvLJAntxhCXr5OBv
GRKQilZyHgoh70FA6SFoGRPFjxmUnTnNIiGWccj9lw5LOo26r+jxX3An6kOmTKgi
BOj9YOj/FTZ8oCso5TtET9GwhI5PNGSKlayTNty7uB/dtRz+EcZpOQ/zusVVBZOL
nriAXpRXb2RvxI7SW2v6OKR2uFr2a+oEp8KUvh5c5Az3B39074tygoopiJGyxno0
2ug95PiXmzHH+DVejpvhBSUFPLGTYUyXxWEhGOAgRU+F3+9ZOB5HbY4DNc9sL7uZ
iKPy5sbrdz3tlyHbcrJmH/ZsIX0Mi3z1ioJ3uXwSF51nHv8CCRIJN6b/eolrcm3X
k2tsXqqwecZWu68mt7aDYqm0v80Fojdkyv8oOse0MH/iTozolZtcXsqh8iTu3jEa
CLcvhCNePkGMCXaVgXkA4lF3gVAXq4LrCpU3t0IuNpU6fgoYZYb+ULYsxblsMYrF
W1l5DD4cu1WX6uWvW9NZpMO4GEOqW8eBZjHuX6EbbM7J1FQLSt96f84nafXuSBXR
AoFOKthxQBLvGyh6TJlxn9eM3V7WSou7ChFCCDWxD02EHN8yB51gZvO8wgndNHBR
Hsx4XkvJUsgYpsnpK2oqLy8d3w5aK4kBzyxLUsrFvSYgF+LlifzLqA1vFLrQeNbN
BeqsMelwVxyPaGrs2BtUjDtJXCcs+HdUNzKPsfZB/EhqzU0nMSDF0Z6rloJjVXx3
EfN/fqm5u/EFEHbUT6kvSkBNc0CH+MjV6Wd6ygzM7hnshCX6V0WIdVfUiPLZ3AEg
g1kM+4woyz9Iy51taK6As9PZTxLuH3upMW4c3TGJS2NqZsDCfyZ1aZ7grbvHKrml
9neB2g6ZJXojfr3SU7SBSA2luqsp0Msga5T0oRUbob7qxrg4208hRuGNZ7waweqN
KlhfdnUFFXFoWwCF05uSR/j38Yd8toKngyZq40SqpPZuSwUwJmcmB5J/dKaLNU0X
JBaN7vnklrX1U4JUf7sQI3p4vWAUt+2mljBHLGMNzk/gdmZ60uSyo5a7p2wPx1KX
dUGpRpDDlIdUi7PuJsE4qdjqemnQUfnNgJnwpXr7Qr8ZcHpyX7iTY2nvjn4eLvPg
cCPIgsWwTgqctBHoeeHEku4ey6OE0AqbpbIKbmLG1EVUdsz6rvoSccamLWwlDRbx
v0akLx3C2rFP5xEJf30sXCsnD8o+1w5hyiJ8SF8SZfWXSsIxxiI4PawRGDgyKwC5
Un2m17isxo2pigU65/T20O2Ikc+Nk5eZkFvQuXC6ivw5zJ1ihytxrOgyhcZEpY5u
EpY/p0lBrcTKjzJ34Z1mtuhJzildRuErd1ltMb0s02YarUvtpOJvQ+jRx6mgxGHg
xbVytF1Ud+7uAaP6dOoFtyd7SqyP4p7vABo9HfpYnimsSiDIw8f93WbGbzp624k4
juLccgbSj4x6EY0KoimEf4lIrpO+cQihSB0JjfdBmKort2pVLzF/F9DUHuVMDMGY
RPzvBSDFho9yR3Kip0VbrRfeHxyrf5YNrGVHGKPnH7MqFD7OVYiqQjzinFTNiux2
SUtT4OOOoBN1t7s/xJAgy+m5wwJH6VZejV2Ymc1pw2kiS7LK/ZI+i3h6iO2ugPan
Gt8jMBp7Qa56ChL3DqIJQV/J5BI41gdchp3TzMVkPiQSAAdgvSsAZcKpEncNeUu2
gj/Shw+qoGzkIiDoZMjnQrickL/UAjYn9epFQ/JdqCLn5YhQGTiJ2uJvQ5HC0ZIr
M24JyD+T9JLnemz8+wpaVEsXcBKUT/VbOZGHrgt2mPHNk23gKKYEk66BWBq+FPkb
qLyCWPCkRA4To3NOGUSiNO5zum+cYvJHu0s8yCSXL6w/y+kIijKuhXHYe2NllIiz
4tgbYVwjqB04CAIoh+/KO/F2osfk9DEcDU9uOTN8qr4bDC91qFKsM1QVHvGWiFui
KHHKx0VEU8/LxKQDiyXLFlLZ/rErzMuFuko5SxCOyf/AyhsG8BmEO/XIjSp+gK3W
G63RZcnd7wAZneJqLMqb36PaRpibIum/J+yxSr3h3g1jb22v8YcQDHHGrqjy3LKi
yx85C+ILAzm13lDwBGPmKTHLBkqmPtOsalHTI1XvVzqCB39WKyK0iKxtUbdyQJza
84mcSLtFwRqQWy5vIHkAyD4aTlKMAtY4EaFfqgQAfs0Qx8Ikqa59iwFvc/YcHQrb
tM+/T1T9FMX6rB+aKl1UpjaTVDhBhL3HRjfifNWOhahRLUZnhAmPcOa6925FXTK9
AWIUpU57NddLobzAuYCgUPhaxmRUVotiVJb4SU+JyUo2rF1KiqJE4+MRbn+kP1Y6
BHW/utSd/vnbjeOKoxS9hUy+2ak2h2myeYr/LHP8qJTOu+QrO8tCXa67/cywsPY2
5pA/TZSKv4tBxYU+IZYsJQghW/s/dWtY3NOATcgd0dRBmt6QvY/AO4KtmEGnADEL
LyUiLKxVxSwBmoaxBqTA+Z2PEyXAVX/ulJyjXjdbslSmwCPgAmNfs5V7EEuOswLC
0jfgUpwceOuGtfYSYDEB/drS3D6U4uDqgrrcw6gFJ2I3It//NZyxJQDaHdPP/xBa
wQx72Q9q02nsN4lROM63QPtOhcmagQ+lBcVALTcO3QZyNCmKOzYTz2sIGttuTljq
27E5aSZU2zGUSYuqQJ+GxIj+RmqdDh+tuCO7Q8cAVwBJuNy2JcTsFXLcI5rxoetZ
qglM+wafvor41w0LpXW01/2w6Fm6Zs5fKwIDI8FPdzHruJz/8da2o3o5hZk8RnZM
kBLCUvqgz5gFW6OuGswyAAhfggj7sFKRoFdZ0Wff79k54o7sQtCO7jwnHvOsyD06
/O4h1S+7EPTCl1GVxHDv7zp3aagaspBXSwYtbLTWf18oc64Ku1qcYKLUBKQKEAm+
2+mMA/vfcMWB3ZFr/4WR6W50Wjf/jCZY7ppMu1tOV/Yfiw6vWFmIvemU1nmssZq9
tGa1bRdKqGKlPoLW87YHOtl/VJvOXmkLT44ONG93OnJn2zoGL9kE8wNgrD7peCpU
AdcZNpAWcR8U3nzezwn8E/4iQf6OFfNxJYjRmk/c1stGi6mx6Zw9Ibq5a3Hu2EcM
g3fbti2E3YqOU478WbksPO7j+Z25/6cZzqHp+GgNFHoFcR4LdiVaG6ekk8EtM3pV
sA3aiRxx2z5jw763nbYoTFNgTJNtrV2hOYDhqiVeUXnkFKbyIlxGNXv+hnyzpZuI
NtlpoCYnl7taRYGpBchyl4BokH+6JcLzKUnGRbARficqyh1TGYHwd3fDUC8E3exq
+7wZ6KYj9zX4ve9qaHcqDS82qwMTIS0hFz9GlevJ4RU9z1VaaGl6RB0hLUOJMKC/
vISiQE8QAeLXhuBKvp2IvOnEsrKiz2PZqWD0FR4RZMHVqYOKNs+obeXulA2YtxNe
X+A2tyzpZJ56cPZlTHmziNgMoG3VcvMPoNbnnwG5QWvrO5r6RCK1G0+rND3lNJOg
M2CYQRQOjD0AvVKij2kJBRWI1lP9dP9dTiq236IILIl5wpoD054CvOS2ApIO3hX9
MrrwSUYo2czerAJHMcV3NRLYr/9KYZxNANL8MsnnJfSLAzFttCPp5ThYwqLuX2sC
TEFa3wODWe2I1VMoaCy2W/pIezW8KAJzWkjJtS+jHEbnQrEGNdw6/aHeZ/vXtb+M
E6SsMdZpVSUn+mf2bKB/RZr0kpDwLAiEGeBmRGi6XMJnj77BM2gI7eU0MyJbFsZ+
L0w+as6fH+/9+ov5pN8ZcBaqqioGI8AqUSSRiYT2HN9llkcJ6vsSVqWt6z7o7c2V
BpK2E36Vjb7KBWOuhNzhJ9RKmqUZrsn0jhOzENqbkhz/EuQtf8G5X22Rz6WwovhR
NXJE+vMMnIOnvmYUQoCG1CjEmsg6RSfgpX1V1Pfr5s68i9SsI9zlbIynf6YdAbrm
vu3Lm9sf+fCAIa0gqUreWT7Lj7B8fa+wjiSJc9/668uVPxrBNtgLARIwlpkduhFG
98htglpxnkli5ydAkhQ/6yMpujyWJhEkKlQdxQVuhhyEIuBikaEYox9NpanAw8UG
A9J+hRqJOEIsqCupyQyxnV0PfIMfMjsKWrXfuu3VXubp6WIvLwvHYnTShQXEbI3q
4n8vliWvY4o6qLvb9kOYn8xzYUGETBtuubU2wUZpyMsBEs/qpDoSdnPaII0Qp5XR
asQg2rH/Flaf4XHxFRr4mK1VdZJDpu4k+Kt+5vRomb+1lAyQSKvhn7AbMe/S6487
27uHwsf9NS3UkZmK2xXb10elAAWJvvWg9AyKMvjBbzIUyht7/TScvVxg2hQGkahp
SWuqkF8iKYHq3VS40ua3AZp+UFUJLlnqmWQZhltP5ec9LcvPDI3hk6k8tm2eJdfC
L8Uwoxvk/BwBDsGz2PJwpFqI3CPWJBgFVe10BUCjX5xigzDNoYk1M3WsLbJgYX9i
zvoimdNy2c/ETd0tPR3EfDvleyCOoWr47awPbk3PtqIsbtyxbQOhnZs011RYr+E3
/g8wN5UdQPp5JUkOKsgbBr0qe6gJPsF+zJs6KmWWCGPx/NNoAH4ol3oLZgZNkqw3
c51wkpOg7Sqdp4ZQ1jy8qEvdeHIQD7dkqL1wMMBtemloo9cvWgfKcDVKZNGsgbIZ
XvozGibI9UgRnPVVxlz5l0aTDKv4iyfQUjp5c0LDVwmptiI5RUDrrn83KOzLdBRP
ipWodEoMxBdx0NVCSfQ2vlqk1lh6QRxewvRHYISHUq/8b5yl1CeQU8p8hbVDMbgb
8IOUAx5/nssnxA9f70Si0dcs5hVogqpn/JpgYjWH/u/IKdf4XeQc5d4SvbqtOv+U
FGgv1/EyzkcP/herZ+7gBeSjeP4Da04le8g3QZHPVLX6/3EXng9jOjKPmdC4Bggb
ngZeXruSPNvE2pIuqaMpbMunebQZVYQXhu5d7TbJZEAJh1aYnUHrsD8d8/s8x+Xs
Y68mLlqlBoY+Bk37QsXIiBGn8Ir3fqXYWai1DPSITopOhrFB9ivEEmqeOjBoJ1+O
03elDdjQ00DQGxCIdWYHi3Y7KyukgDDK+sh1FIo5ZoKymVdJ3HTwenQhYXpfyISo
ENsYyW/4g4P8HxmmeGQSboe9QRgAqb96kREnNYIVH5ZQkyq91J2wZ3eAVOG8x7No
DoiiGUtitHkxzKUdJrwtVebsUXNwkBBe2vfhN3685FnqKWM6n4FB3nddDRaeu2eh
LZhcs6YoRngDXBpfQ8C0FB+fusO1GLIgiFzvO3V5uHu1toZqPVJbVuqH5By/Twij
2WHpt/GF/eJ5OdZ3Nwia+Qa4z3FkAy5ufYjEyMpY54qyFg5geEoGfDhL9lUgK9Ur
jZA1Spo0PvRG8vumcBeYhKkcgwGyYAfab4sT3TaCA1AWwsf+BpSBDclVpLAVnqiw
NCqv2Gyag1VI2Pg+0tJfgXGUhE3cKJTPmGSETcb3DocxwtpLux0O42eEllt6xHk5
MfhAZcdr8arCkCRcDJf47O/ykyh8vnRfGb26zYdLsLFgAR4qdoIxAEhE6d4vcAYD
AeY6dzo1BZ7O+zmPXq8V0Xuv1d+X/bsasfAMG7Dy4d0wla/BI7ci7EA/9PUVwiLd
ESfxaaXQ9BHMpOem+uyXU+tQE3Qjgnso3ptL6Hi0Ynaj7LnHqajuPL+5RqDxU91o
VOnSFeGFgJQP/0e81Ol+MS0CZcI3qlCejOA0HihFz3ybsTgYANDaZeKofNHmk/vz
UHXypGoRks40d/9tBYRQGDwJx26Pzz0ukg8ULCbfX/hDcKbYgfIqj2GNNIKXlfan
4yld0+954T94yh4wAP2IGRIIZMpur6WMdFm/FQNUaP6ntClAFZB2WUfY0r4JuRyi
EeRSm+O7/7AV7gR/QLTDGyyXJpeBXCxUYcmyWX4KFqEydfXLjywdFLDv+Cos4AmQ
paohSRcxb+VJhPUQsSd6VkNaQstqbHcY11b56HVeiLv5Q3P6G5HKaix1pNsYyrOw
LamCC49hW9NJ4/gh6E1B5AruRARw58eHz5sWGtDJ7BqXWyTcuGbmWYdp5mL02Sky
zgjV4km2hocwPLneCraIr/1ieQXsIkWu0ZQO4vJhh0lTjodqiL+t9uXEw8Ik6SUH
H9ESpimSkuhBnEjtzkpunxA2jQ+HdBvrEEdzIeYl5orZns+sGdTGVlY/ii6n7wAX
WErnefx3rP1DcJYabDQa1xvJNAs45vqnkPoz5N6SBDF2GnCtTFlaFJ3LrAT1PdgH
ZL5uBClnSJjgdj8pSGyMJ27fY8ptp5yOv7qS/3KgcLbkSdpTDzxJ0RtM9UKmoGNm
L4HKTw40zrctiJB//ioAnDSCk0v6gRx2STwMP+GSIorxao11He8QeYcNKHk6vEf3
5s5mWB27sOTBJgS6tR9gbOMmr0AGP3wE72xHaEVnHlYEMHZfsWLUR+4bpSuPjQFO
JIdcMl3XDaTROghmeqLQVXyY6atoCIht5AjkuYThxDPfSre2x4BDvaJjEN/iZUAf
dYRBAy8SOt14Z78ALbc54FH5YepGE6GCpL/QvW6rE0PhjQhpGoujWYZvpsUr5X36
6M1DwU6uX6BAcvsspaHioT2adVQ37vVD40e7tlVmf4qeEQtv7SkYBAKCnd1HO5B6
EGlQanLqU91lbnE3aNnuqPdKjHeAwm+/18S823sF/sJmTH75J1UHLB4bprleYi9L
OTQGiWuYn5su1qkL1YgeozoYV9OIVB0tcozDXJ/Udtj41SdENUiKOQqvkx/V38Eo
K5thUfr4zuGv8RvigO9T2GYteWlexyNrqi6LQZvoqAW8kERHFUaq85//Fy0nWbWL
/RHOVaeebnJZuA1FLf8mS/Zdz/oecdXWdA+DZx62FyDDkp27+k0o7dgumrQrT+TP
DplFuUoz/Pb6bc9iL38IsljKK68gh5pHqCybCI1fHvIaxfy6ktmRaoRS9DCpSmU9
Isy3Zxv79wQfnogQKrj4N9VH8btDkyIXnfM/b68KvkK61Md09Oi/Qu9Uu+N/M45Q
u2E4OoKtlAUrPgt4VPDNMT4EusrGKzK12tjWtoEJkRRIUFZZcj4nrOQqKJ710Xp/
orBJvqUje2eLlLFqM5hYCwpTge/jSqtbL0PYdEIgUn2+D7Af4345vXnlSxEG4JLp
mSVIsClUy6FORUpOU3JoNfFkqqOWit31zy1s5oFtg+NOdOfs/Bfgw8pnyvan3uk9
rfVk8tZSBoJEK+IAbEG3XPEA0mBnxW8zeryJa4L2kk/5esib6L9vEQ0AWQHiIRmm
DJOSDl0Yt7TNws74PsETxEBFNmagcxhwfip06IK+FkiLU1z1esUhM9kesnIl/I+A
pUJr7TfxP1ofAlIWWGv4OIb6Zdni2yXPmj6xPZMsQMTMON0lESBfUxMIDS9jU/ZP
cSR5c0oPiJIM/Tj6EsNo9VlvlZND8dF+SBstP0/y8s4N445NhQWCBc3q+3WReDwa
4WYIxmXn8N5/rIX3XFtxaEWDY6NTeZtMbx8HUkwokiS052M6XzIMpCMfTFdWNaLI
pE9YiRxF1VZ3D1SPS/Jx0M03xVBDyaWg+rLPOsy8Oh6ZiT+WT9dw0ndcnjNh57xC
AYIae6XKQ+uJmzFR2WZzZuloEJs2pjp9zAunkH2iB3gfEQ2WGadQZpHRnmfsIK7P
tVfFNVXq6U8h0XfZPhleXX7lQJx9yxoxsfAT9ejx35C6CrTpFmW5OHXeHHZco/+l
Xo/p7gBdR9bLlLstE0pdQUlUiQDfmxNcN+r7GCu9iUfGT8gB3g8wn4vh+oQjMAbP
RJzu+01xXhGvBrPwlD6K9f3o32l8FLpD6bZx0NaSPXdJtDYReXLp/3AgnIHCL7OK
9AqgzcljIf8wkLaXcPH8xCFxpxvWhfGgzi7gCSVrXNRApbRy5G9RVZZdbo5eod4w
KUbMcFp1q1VnrtT4p4Z83Z3BVJpYraSSK9WEd+ns8WQ0N2rybkSA4xugIYkRklGb
9ugcB3ozPmJlAA9tqljinOHfAhwg6i9Rgue/v/fvQqPOkKS2MuE9NpE14PIvkBJb
pskPmLXTlJpxyQPzeXj62Vdwe0qyv0isyO4yE0+dkwRvOrBwctK7n8e/qlne7Nqk
hR6foG4jLa73i9XM9klJFbRqVpomSaoMglMpgq5ec51GR0UA4m4Vw+WSkWGyB2b5
Q8ex7HGzWgqnpDMQGEhPwhZGeXnzNtZRyBtOi+sHW4BiXGfm+R2PTulrhuHM0aAu
33Ppr3gyDFnWEO+IgLLTJg35oXC60BvG+gHyA2betD+id6i/x5IptAcOaeIfLZBH
5tdciMuqULJoTNBpr0Ql9jxyz754EHwOFvyp+ZCyvqOXFgKLhs1cnspbXayGVjIE
lV8IZuEFKXnZcjqkP6JW4JrBGLliexURWVUzSH5yw/3SXtVMr2ciye0UZ2ZQcUGU
yj345a/gEx7C1jhPDFY+vOXYDPzry7vyT7ZyNTWkP8bde5AND0KC6efkdkdTu90h
oAW/hADvb16qew8yfNXU8ZI4DPMPNMb/C/mNesuU6dZA1bb0c/2GDoJ4N6nj2CVQ
/u1g6+41iGNrqmEmZDUXT4tTQBB02gGHwLyFy6o/Ru1dsdWmU9PxZCHprquh8dsV
zba812B+Ng5CKekpaR5qaz6q3hv5Za07GZuGFksbJtmdGuYqCLu2lgupLeoFKF6d
BLwEh7uaTGgABLnbq9LmMi1W6lFO9tCkvH4KFJk+Ok1ndlFOOH9aOh51kwW2uLM+
Z1lugiWXEWJPThocf6tAT3pwKuWNGqDiAzHEUsXzyfs/bNptHV1iFhAUlYJgMGGS
mL38mHWAuQdV0KQWP1DoHgryidnVKBe5wnSiSiqne+OyyhFxo2lLY6rM04Px11US
a94oUCVE0ZOEgGph0rb6AIb+MIxSpg87DmwQFnql2GFV5spVlGaeiqIh7AjfmwMz
6kYsajSmq7LrYwp/4yr7l02DvynKtZVrw/Byp/8v1d+Pv3W6DIic2Is7ES5qx7d+
tl/DXa+ooOd9cBpnCXrRyErPCvyqkIFMCWJ8UHa4Yncmi4Urag8YoluokqbQr6q6
ZrnjIwJ861zGxSSbW2lmkGmhGP+BcdvcwQAeu75X5SGx00yROj6n/Vhfwpxz6BA+
ilJZYvaeNY4d3WMJnoo4fDk3cE3M7GKVFQKQ/kqj6i2/6Jh8iq0pgjICzOOn+S8r
7v0VkDFAMrw1EYGVxx7P3fP4vWgsUYD7Y7UCDO3IUu2DhJbkd9EwkprcWGDdOp21
/G3MqIptXudMt20liOvElgSMa+kMJ0UOha9MOgEPKowk4502eQAuZhAn66yY7k8Y
RwoG9oH1WE3b5jpMfJs2dKv+UHBZDCYyFMO8bDQlD1qSMtW7c/xvDM1VGJlM/OCb
xqENdjwMI930pmAOgn5/88nYBSIhojo22Gj3nOqhslJeWFubhKPqIbGCBVzfxG32
aCvkXDXnMFG1ZBcjkwPjatPhUJRhTvKOPHumbzV/z6EroaE7SVcUMiVDoRFr9yLK
uqf5Ry7FtM/pAdcj2fg1VCjx9NiO0v+EyLoPw4FsNvxD9pX4E+/DILpf6nC4w5gL
oNFCPRFynGm5QdfSXlRSjula17Kz6HE5IbSHiRQMnvPlgIBZRZx4goQjQfVUabYn
yGNapIpbT+7DqJfHyAnrllYC5XNBuvGXRxtSU+cSuiGqu8lhiJAS25SUofnFxEv6
o10eU44PGiAxxwyEgDqiBegL9/I9OD9kvG7VJVUNiriUIUgvfGaPD8KcvU+1DBmZ
7fKEY8k29GShwMgvUut4HRLwrT5YfnGY8nJQiB1AjkoRiM6+VOU97OpczMhrwHqk
fw1HGdppu7sq7vfl6R+SudVS1DkyQIhbrEDFJwVi49xpFV/DRONP/rZWrsSEv0Oh
J4J+mEjVeiiF7Iv5YJ1E3SGWclm5WIzShnmWO4bfk9UfgkRyeKeqWA2RoNcoFZgU
0qRTNf1mURuJI/FkiJki8v1zXqwp+l20d0o0Uca4KhFqWwb/5JSEW0AqLkrsCZ+J
86MZIybkH6sf15yOHhE/OzYQmLaNmhxxA2j0IXppTt5HpaUZ+z1rHnAhzYegbOSf
iPSArYSD/KYUp6Oo2ItAc70qAk2DjeEtw2cw/rsS+6QJE3DEgHDeqAhoxs6ADH7M
4rFVYrEsVr9Uzu/va9ghGCkLBDc/cygBca9RMv2Cuxc5kN3bv0eo3TcT9+q1ErJx
I7ONHCJ7tPo+tejr9h4cwyRIXjaIqlAabBLEwO/AOhY9qChZSRmkE6S5QOCoOpaF
Y1oQhYEjqgf5Ot1pntAMFnsEZFwYih7aO240XWHC5v3YhztvhJ/6jAjoNh6kn2Xz
joRMOAPImS/Ku6mZU3l6xHEvj3MIJ2Y4qYUuHq6j7ggEedruQ5kVwePqgloFTYPU
6HcY+ooTUSxrCBsqo6kkJjEaMy9EsABt+wFCi5/4PgbIkcTGRmdmC66bQrpyrF67
RF7DqqUsoWk6tvjYrgbwRSTvLCzFwH3gLfEyl9quiTyQ0jOQ/Du5vK3/GCEEW2/n
C0fxk/01lYxe/BjLpZzb6ylmolM3Vj6HBQgvEraNsuKpEXI0UX8YENRj6pDMuEyN
z1PZUbbDzHLJGDWs51ICPoDwRXvCdwsS9GXPtHRf1bwAirw0dx7pd5FN/ObHj7Vd
PW4JZyIc0mIfSPtyDZEfY8NQXKpXg64YjdKkmT+yFs7V2Mb8TxA/BL3/MlAjBHtQ
ijw1SIOk7j/id0zwcNk2Jxw8h2AK/mUZFVuzWl/RfDJU8eOHWz5xYg69V5O6tmnc
T2Q4mUjWTNJEUHmhzQ2ZcKWi6pSlU9T050Bk8Kvg4mSO9Q0iR4WvllR6PXTPW/8N
4zmCnraoHdtaDPoprwGcDAo7nhN83Sa4cBr4yjKx+mvC2qiU1QG3I83KgiS28H5B
7r+fKaun7RcoMCa1S5193gxdZxSwlHNVY3eLpZirjrpZx6Jo6/8LiA953I9NrMnO
ZgfugU2Bqo5lO0WFkNelxL9MBVWlixIp3NErzWVpgqH3NJpsPH8YUpfVWXHzy3ct
r4AitLEjI6LV2YCoYrTgLR03KiIFKMBgWeRs1rze57BdW8D7R21J1sxkFmJkJvl0
n5tVNw/0g8QZ244jZOa5icZeMnMzqBD3GVOxc+2lBPAD0r/d5DYaCT/a4Qx4eGSS
BhyYwBLiD/nMT51AuVZ/8bfIan7IbLgmbWhRN7IRUG7V/WZCl5FwZ25SqodYQQZk
HRR36hmJSrJW5UEOL6OQuwxIH6FgMQgPsWR76WDXBzX2OBI2pEbBB1GS4pLnnfrt
LxUXCRSZkRxcGhWLqzPYtJlOHwYbI4UHPY6jpUQqb/v/dZALFIO00wTDtOrCVBH7
ziZgZ+xl0NIpmyQRFGIYu7EFNRzpEZP1DAdHaCz8rr3qGsslrwjF6dMyoHZUUK7f
rpVO7nffIy+W7YF54H8hyJ/xhBNZc6O6rKHPWLPfvMM1sKD/2aTJLfZnJJ6AUYpI
MKFD6tfmHbAZ1LWjGiwDOCKUuB2miqjqLIXcE4T4QidLihcPTMvdnSRGfdbEhnsA
RG2y8P5H9ZuBbRN6akJXR0uZ3FIGvW+VTQ10pGFya4HBsJZblORCYT7dmy26W07Z
kUurpItpJKPZuIw+ib1bp1QitXP9uyjqm2wa5jgXYZWsi9mxekRrYDi7vZvnBHVy
rsb90v4NG06ZpV8QEZR4Zi/V+wLZpVRbNqX8q7YtIrpxGKgIzjB70Eu4tk5cuL/J
h8dW7DLlYLoD7RSn5/oReZ3aVPgg1Z1p6rmJ6Ai0UptvmElDJqRm017YyZ0WPNWU
JiaB9RFDupXy4Ljg9nAsyqD6UmZij23ggXAMRZdCt45L8OITLJ+O3m1wL41644vI
Mh5nJE3R7BxH1AUAIA5mn+nFPFpwyx60t0UwK/1zKbSdHKfWMim6K6UAqG+hYaP5
2vb3obaWkcjh1XlFinT88XaObLnP7shWvx2OvPFscwIc2Ji22cXh0U0aZR/+V92N
NhyM7t+q0VqsvlmO1/qKcNCdjNbXy+AaaZoV0BovpGZ5BznEPIjygIwbMXN4PNv3
nFXG+1kl7FOuQUZ4rMqnKmNKijM6VCa8P6bPCLiC5/Vl7miN245jc/yDZ7FWLXu9
IXV9q2IGLryw/ChAlm8hGqinlMxR3xzehIS/t6uoESBV9BvMlEGXccst0bX7tYVz
HM1xcSBGxCLknylWzpIBFLzyH1SYmMOq9+q3pj49YiJPsyR4RMYUumLRZm67SM89
2fW0gKzMpbat1U6vtwUCMAMgG72vyZ6vir+NRPDhLdgiNW85s8lnpI+Kncqf6vmx
e/FCFMVqUPojOYrJ/5mCMsSpxzs8DUbRlCQ8vD/7MARt84vYxHR9C6bVqLIGEBRk
usyiKgNqgL3D0GH9MfMLl+t+Fer02Zz1uWADPbuOBJ19vdkvbkCbycwQO20gq7qq
FCIb8x9b1r5GvW2v4F+tTHhwqPOxPmys5woPgqaB6Gd55u6wyiif9cSsEp+Ydc03
OtbU1cDjCuJ+r4+QjHAxL0rZUX6zbVHxOQQJvzlPDYUd5F8Y7hy2SyE1mc1sTndB
j8Pv3ak7sgMgV2vjYzJD8G7uEcI/121OnCC4sNr7JnlFp2OBNjoFRXUhljztaS+g
yUVCJydZ7samCRurzvHgaYfDbHX7GCr9+9/2yJM26YIPL/hJYeX2bkt1bQSx+QTL
de1UHNcO+BimQggO/5ut6qR54TROvBpmUq4oT5+PKVAwgYfZBxaQ8UFD8KeThMIE
GX5FPvo1UK3sPTj3dABykvTOCcAyI6trJRPSbXdKOQ2ZdsY2VN3gdyBOT9VhwF+0
bTbhjFR3yTUzajmDq78j1SRnLATZ0iFZ9CduPoj4KeVy9dPCz4odvFVOckNIvO4I
AO6/cVB/m2K8KNxbgBXt1gn8UIFLAc4c5aTuHMPbrJ4KVewA4zHAIcdL00DrrWHc
fQD1sJ4f/pSGpEGkkAf0L0doGh9PgIGGK7arpbb8qtW7qc3nflrKera76sHukBL9
nTmXmV4xlxtL0VgKbxSWFwp6eIrDdVw8xCunSae/SGXA9H4c+/mAAxNCdAWtRWFh
+J/8ESPkwcdbQIiAb23gMDE/aaYfEZZ+vN5o4atYN6czA1wDqG0bh2c/pbd4kprR
N6MpL2W35Gad/SNveUds9OJ5wjXDNME7EgtONlnHrUcVsGTa/i3tewu62YaVaFU3
Of+mJUCi+VFuuA2RdlkeWyeLW7CCel5FaUM7nJan7IvbKL4V9caLAWtJU9zqUnZI
Mox+J2q9NU0VRTWaVJTMvBjeZMxDbXa4hIZaBZ2Zj7Ftxor2j1FBH7TJhiSY1XmK
lH7193HjBEYrTWnfk9Jeli9qUK70Lh6sm8NZr3RbPy3cNjXZ5iwkvd5JrwCUVXtT
sfUT6dcq/llvPYuibynJ1z2sslvQt+SQI98jWLNlzvw2mzJ0X+JuAoc3o44TGG8V
38SYoaDQxTJxuPyLcX9RVJMcBZjp23DpIcINKy/wnWl3/2DcOOGbT58utA+YSPaq
JpQD1Xc3fxi66sQgGYooTe4N64BB/vhsAXg8gEm7ygY0J2x6+tC/JJQ3MxZHFX0u
xzLTCO2jpjuVO+MF2aNQwWzrgUBsT4QV/QS2Hq8yZExRGev1w47OXz3VI/y2UEZ2
Yz5dbBhjD5b1P2X8VBTt1/KEGKdBzoYFsv/8YCQJ5GipUaFUtnKWI9YWqotWnWeI
zKwH0dNYGyeAcZwLgM968GdGtN42Kxydrk+WGohcngdkOTpVx2S/3pndP8dZ61+O
mONkwkgLca/eKHKI3YPTOeBPOSjxzmQFx/X9B4WNMfecyuqukaa4A4JI+gj/9uMl
ui/fUfQiIjszrqZcm3GHB+CsGTHJ7dYE/xU2wtWbVDkkUusi2zEDNK1n2y8/uGta
QPxFNueaRFYHyP6IUuoHuxiT3ugBzlqWNnU+vYx3xsJYfPGyKEIGMuPFLjYTWkG+
ocmPk/6+ejcFbogAjnyAc5uiYmDlMt0KlSYfL+XmMQGfOO7y0F58mXIpFNiNFH6S
xT7XY5GaOmG8G3ZZm/txoqQ6MiwSBzVBTbH5SQhepEcVFb+THGY8Qh20rmE+O0y8
elW70ADDFYFPFdAyClW8JEQZNTf/z5yzm2e3cq9o0Q5QQ9y6dmrY17ZA0uGHVwW0
YSlDTo3ZFlT0qqom+HTk08dBpJmXtVFA9AL8KsJRogCyA4TVu7CxDVjJFzuu1LTT
s4MU4Df1DcEmAzV+xeXf7+s2ShehiRVqtVII8amLkv4UvqnuLoUd8eqERJC0c6nk
au9R/KxX4EKuIyO5oNO95NTfVA9cL8rqJOTz1jm7olUstY1aN69FyYGlIIa6CXSo
dCtBMh+C391eJLQvSDbIgMuvtGE8KO50CyLSBccbiCEJy820ffukuwFOcGPljU8n
+lTl1xl4L0NM6SoFeMJ6xU2SGHKmzkzTzGI0TzdH/rcEEf06ndRG4d7w/SdYIa+6
wSCbWRyheJQxI69MjKTJkm9JWFCDx5ZVtD75XvZfz2zhrggGVNLNwTf8hxRiW1aD
XBfG5ihBGqEc4ZV+9GaUg+XU4PAUDY1YR/EuDtboQ2mUT/ujcUi9F9r2yC9rZwoZ
yZocnwgnjhv+0dyu7xDiMHUdbYk14Q3aQQwt0nc2Crh0gTgoJOb1C6m8i4sGmQh6
Oo0667VwvXumd/3NJhk39XcZ18Xw1NggIpsMcSx8RjzeQY9qJ6YUTrlW2siicsNW
hda7mID8nx/ngz4XvnPXzfsM/47yONLmb6Y4lSBPEOQQgQ5BQMAQIv+xb4+u5HcH
2NsZPZbuHk1KPkFS8FRy8JjeFclKOSUMbbnIa6ShGxjdcVyC7aLoKwqmZRcEQMcc
SMUk2WryWnbsacTJ4WZ06mzQXJnpDm6xAjOirSpCJ7VR70ToDh9yFhMAw26TFE26
+Tzlii3IU8Zzz1hnnht1Pr/5Wiy6tmQ/GZmZG6ku7ilojStxx0bNp/gEduzBO2TH
Tpup94mvLKZP4/xxXDZ0K0CWM85cVPtsfFfKn6qgbs8RTRl1q6+wzALSJ0U4Ogxk
X0DO7Y4kKFRCGI1MGhCdp6nUjqCHesfqmKvlDtIDJyQW2YHm6loIiFj04TnjnYKu
ybEmJ4c+mlAUtQtjDul9tbV6xRGfzOos4iUPnWPV/2vNLn6np5mLaCtbuJUbmz0C
lra4GUNC2D9sl5Ah9mSywFiw6lhJIvgEzXa+ipF1ceKcJPiOz8FohBbPiNEgj440
TJo7If2gAxIDDMDuL2Y6eytt0tG5rsqmBmsfm6OSy0Jv5wuOnZ0e0YihDwj8wo1T
qXY5mcNL/4eyrSsWHAAF/jDil4zMyAl8gdHW6QdpSsMMm28RmAVmoD+vYUtFDXP0
l64jh8BDM25VxJRw85AMRkiIgShLKMp4PL4CoxS2R2hdlg4YQUIFki+DSORgBQjV
jewc8tQYkHhgUH90JGkN6by3WGzVmC/YtCBsVacI1rmqnha+DvzvOubDvp3XowX6
e/Qi2k4JvIiQYbcSasTOQawSLkrzIy1MbZkecKXRWFdQdqO+CgttnaMhcWU6vP3G
GOZm/a3tpsjURAkHq9a9aIcy3RRB/Xed9V5G4cEHMhwK4V0ZRgyzwBzyNNUJ8mhf
ElZ0c0W7JzvUTRbh/NmcD9ISeVo+/0Ti+7JEA4rGjoJAYtb21nzNvHAg3vNbjnPD
vIz+hD865jhC41k0RQAxYY7xNP3TMS4fifrET0yDjrM5Et3QuNGu1hQH1KWUNA9Z
M0ERl/LFCEDE8pcdoqTbHylhI7kkLLmby8MM1ZrNVbf/5b4qbb6GomkO5WeOUdNC
pmbuqClf1f4L1Nfr4riP1BH57zPmWWSopgY/B5367blw6Tnb/A+VMFQ/B5frUgRn
Xj1bTHcaDLaTku2+fwMBWoCAbvgUZlLTFnvcUIMVEo91m9n2aBSsRvZ96RE2PNaa
SZgE7d9naZDLwk0R71GMezPZ9TutI4eg/sBeJf/zkMngUZ5Rk6CDSq2/YN0XWDoE
WacOljUxMJn4q8NZTcxtVJyHvA5kxwhvh05C0IGAsVIdE59POYuu8Y/bxoVQwJfO
epgveAtffU8l/zODEy7in6CDq78TPVG1YES8UY1tgEG8E8c/UKdY7M1f3PKaVFCS
B6VD54+CCC5yZY324KjNT4tUdhgSMBhg6SIT7GWKLI85FxMoRV6btRlG4rnrs0+/
2GeWoUygBjYEYiaacNxwLHegUsEYnh4/xqcdC7VMJOgm1d7xmy8hU+wl9kXT43fy
9NAFNLQ6+cARfRSxbMtBNRcSO2WS/RpJQgSd5KxbzgajpcX2SfJjJrxkahFoUgvr
Uj8lt2Pcl3qsWGPl17TH7zXKtvqfPCHz0WK2TBA2Avc+hUrEvvsHl556MSEWMeD6
UvP8XPKo2RPJ93GxlBeG+LAFYY+gJBclNvgFbp6664l+3itxus1lFMSDgMGb6Gqs
1Df8BC6MjDRpcfOo9/4a06jgceBw8pLKXpueZ31Vv81UHbJKBv9Y99ApRevtB52m
to9/StqAvXl9iv4PEeNu2PxAPDuhWnu67upa3KmuwNm+bBr2aCXUx8qVZhuICc7q
eSyQZm2kxfzof8cDfHqdkFrgLCfuQv2x4YuFbKvayHY9ncix29AZQS/06XxD759F
14IQcTMT8+D2oQXvkW5RDMR9/wF52O/aE7rn67fei66WbLKxKwbkQ1coNKZ9cyHc
1SBpV2DAD/zblcbseFUXSw3eRDn6gjP//4zNcZJxRfofC4YKeg0wpSj3dOhr3soY
MnBrtyj0CfC5A3PzPttBsTU+6yspVP8ZCcxp5wh1dwx0RFDYj7C1mNReBTJ/4k5w
TAj7ztTR2TnsW/9IoiAhS0Fm3pawKJRDz/SFKGoZNgW3EtsKGQN887r9g3KZ7dEN
w8fJrNgNISle1F1XMsLfuzjoBTudKZVvKjkPWtl0ezfbgH2eppBRy6KqHQyCXKSc
qu0FoLWuEDFtI024tbi9YIui1jY4EhiwSu116/kVXVQjlSGP3KDeqZybKhsvITo3
nVxi3BERnK5VF3v32BXNSU/G2pZ6fyQCIyod/zfnkvjl+DU6Q7cN+13hS9KT/xA2
iDzf2MuCA+PhJHA80gv3BvBr/nFiNWE8u9yymzdwGhwhgQIGGARvQuFNsThudiHv
2uPrNfJPtYp2eqDf00CkeTfYSU5ZafhVKmef5T61++E67O2xQqzPX5JmU2TyGHBM
pjBbHqJw8MIB0ho28TaHuUJOe3pEAlcGEZTMdc6603/rssp1yqhUFEsR4jHWCQ19
4mfce2NJKXId32WdQde1Y0RQvjLTGgHjjGZnSnnTWs42lPxe5vnHTQRvX8JuoCFm
MBV6GeKHKl0V+pK/kAOaYTDGlSkeE0pHTPhLVf6RnUagKN8bswcciNNQMbppjUZg
2iUh0d0xnkOOsHY5BPIIFjLLFiHkmaUo9+tImIMetBVx+ErMSBlgZ51sdD8Ieem5
HmuSdNX8e4j7upcP7DW/TRAyZh9+EqnFe4Rkv8PjwzL/XyPvK0LPIQ63DQqsLsHR
Wbla9BJwCEXvl7vYlkxoWdvuEYBgrg5RdT/QrTHJR3Y6TJPpxDe9qxlCyj6Z4hDe
ja031lc0LGQlxTbvH8xBGgU4dqosOSSa8Z/0ALkgLE+cHIglUzS6JnQymgIq6ksl
oQ3lIrxZR80IKU+6/sbQpo7GI3nQCxImjAwPPpJuiF4IwyMZm6EwYlZM/VN63xIz
/MxcKe9WwkKBp8NJCHjaTTaddwan8VMnjCD8aPGy8piQJSsb5C7uHcLh9eRnATKS
tmH9pPFwYwzNJngrtnado4F3wHRv399Xle69KXnEuqZi51HP3OrgMGTOcuHKqvjb
O6+cPgyDwD4KK1uv7SdfSDdy2Za8Ygh+rK9zblGZ5eoTKCgH+ORk6zogn6T04ME2
9hcga7/WrgDho3rHWJoNlxvFFZk0lRX2JqhqQHcznYOp9AOWRGOd1+6jjNQzjv9t
e0eTIozfIOGPhImpv/c/PgKzkdVmFBBZBhty2dRdIeiOKzBeFDGPIvhHMdciqblA
EWTxvIL86aOnb9tobuinwN+thk+kr+Ku1aC2rrNMZzgbaLd0fRghtIKfIzeHAwpp
rthUjJxjK14x31uN8lqHvkSIFIl5Q3Tnk/J7/F9aJASQAFyCVdvsW7AhSqlubMqP
ltPG22aUF86zVLRbIC0XVUvsVNGuztDyYn2f2+66p2fjzHYHV2lOoLasgWwojeUc
Opp6h4R9Xo/2NxKvfuL2AB7OrFlHpMhpu5E75tj8+M78Q+KNDoZrXjujkrL1+euY
hwSmO1BK48O2MKp+aHtdzf7EQFV7rrg8a3jTFFqS/oBHYdWbZXR/HgUmouyF1B3v
Mz+H9j1p6om7CdvVPDe2Hn/k3Jdr7LHnYxsjwLHnwc9TlK4Eaw8p+lmDbSqWsu6R
XNSP77R5egH8WWBPUqA4WW2kjY8K9vOYVi67JKt634Q4heHUNnMZE0EdLVFYBypa
x/ao81rNCMTVAtEmpWJGxh4YStRGQBeOxqwZJS3LCsOnBsUpoCGfi+Z6IKi2V9zB
HZjm2ZgqQsONc6JqyyY4kTPiPR/9Qqw6UQ8NsTi9SuVXFu/UWAgPTO/0rmCk6A59
wbnBL0h3bpxhnFtWVIlDzwCEC381PtMvsFmZwBVJtcCHcdA1wx+DndwH2AuEebck
iqPh7kZ7myMI/Q7t0fi1CX7Gxd+YtTkxYsBC3qE9gLsmSOv3iS/HtucJMhjxINRU
FX+MnPxUPUl3ukxkZiQQKfPXGMYMXwxRjBuJGUWnGeYGhPFCZ5hCMUgYH48iPT0B
mWtzcGNbkdjEaK5uPwQEiRDkF6jcDV9bQGUmBFKIuZ5EwkhZdp45pe94/z00dsgy
SIeX6YNkk++yrJZqSY3gZCRQGDDbSF80f6MDmkX6pYKDw2EHa8yShPoyo+EiKN9n
1MOYESZj+xuX1ZjjmX9qzapLHNz07/Ks+gl+0kvqgG273e/9QAzT8yGTDoJz877b
yn9tBk+ew8mqH3eEkYUkwMB09tjqAvUy+cN2vaEaI29s9fjNBEnBlA2PW6aRCZA+
ip5Jer7y3hfbj7SQGwcuGiLsLmdNPZQQrx8JD6T8kFedPB1V2Q0UOawk+pagV1n+
V7SBuvoowAXvXepI3oLz48Z1w8LDD4Kad8PabfSoDfI9V//UiHfZiCbnNHMGuixc
uOtmz5YSzZO3Ts0BwUW/qxoslL8gPcyFaGZ1+fOYLxjK2vVYXY4h2u6dbittEvDW
q8RqWJKbaEse5w+mL35gbQRP8H7XUlrqmlP9zF3KJAgqcCC4pKp2VfhT7e5vnJJ8
hj2R/mWR4uRLL8KJhR2/Zn/yin9QKnfdgDkxmCwxVTPTl0qn3KGIpnjxEAH2+40G
tW4Fsp5yuATOzCdJeMfMBrBaYCfgHskAlu8nDC5cHiFvL6rVzl+MJn2K++FIudyi
hvH9ToE3nJYCwizxlHcW2KfPwWBwTDDIIfSGp34gkYBZHgc509qLRzMLd9l0rMJ/
pxhBL8hnO05ioUR9sMWK5e8oAYZEmipboc9s062ytl9KQgFgpTI1o5G+s24TMm6b
3ucHAORajRdZ97o39uBfrWjNs0DlxMmaUrkVJqGLDLK+n4fh0fhmszyzqaFhy+4Z
KOgrSembAyOHcpeGw8ouwe44YdiXh7jWgh0vYVvcAZG/vV8e/y808swkv7B+Cf5+
/rixkwE8lCPZ6WwobhBG/Rf05tkuEZ1IUnsEASoDOXWUHLYteSRUVE0pkuUoQ84+
hz0rjNHEmOM/AipGKa+wh1/ZDUDaP8giprbdrdlFubQtWPDWen4/XwrtJdEbtojX
htqvNuUnYfIr9swaSv/LUheZ+eqYPvmtGNiVLqA97I3W80ECT/NQjtXlj68+5wjv
aNRFPbjQg00R+fHPrZLAmIH1GdwvyydZ+WgyTl7Xlpcu76EghXNL61Tj78EShDmh
IKHwHHJKrAGd4fVRd+lBKk1oBec+UNURL+PUC66lAtJNkzpvyaXku6ndwjn2HTjt
CmOsk01U54b6kh9krkEcY0J1412F5XCra7M7zpx0s+VHAxkVzXc7vK8+1nTuEjpo
J09QbOTYEGBQ0YWzDbMJXX9M3IfNPn/4921m9ao15pGoEk1yE7piF+lFsnfXyOnS
F59Fo0+6R5z4XIEwykBxpo6DUmmAXLx24jlCmsDD3AJ46s+Re7NC+2c1nxklpZ8U
LKQyE/xvOkIKuqAVnFmBHdHdISjWNZ1PsoS2CrDcSFu9inw8tHu/u7TAWK5y75dG
8/adrihj4gZ5Nz4Xgr9u8p0MlRxvpwkWglxWyyzSx7PngdBukW706KlQ1hj1nkLm
YTdJkTUkzehF8IaC/QH/lSnim1kuhC0IGR3pjTSrbbBrFqE0mjhF7AK6+hPWxYEC
tfOYxCtNWnkdG4SJrilevxM6PHJgHarqz1M9x5+X7M/0oNep4AdVZmpQUcNudIQW
y7RWCaf/Lb+1thfKaP9JhMz6PVqebLr14K29nwS8/s1yyOfQrI5owZ0Xo1eWu4QU
6YYhMXoxdjnxVRmXoE5Y/uW44vGQbHYvdJtwLIrOzjLIRd/tFdIEkHDCV+pa7V9u
OOQdZrsSFEVFrQ6xk42t3oSpahQwlToFcBfFPn68rFShPAXW+lHb+xsY+VXYuOKl
yIJdnKl+UbCpRjcrAMz3mvTkd5kLrvdCUFUIqoIVlbuZK63UqAqyiJ2b4cYnJOlw
+N6qOUa6LMVHCFvx6YD1Vs/BF/XnoKeP3MoxpUksU+PhXkcypC0eQ1saldWqzDz2
59vwBxwsDGdOrheenLZirw95jRJRS18obxAbR73WKdFwmQjSiabfM7HYM59NhbZt
w5JuWyXRsdPbio4pn6Jog4MXJgSiyS0SED1xuMa36Q0Y0eh2Qln0qaXVDNJBeum6
+qr+OSSjoYPqk1XGq5Glv8F2KiWqoQ+V/0FP+kFyA9sI0PgWokRi7j4W0DnF6hkM
9AvXeKT1z+j8Gdc9aG/jiVHGkyNK7pjImB+2tV2yxoxaDVUFyHZaB/L4ySuLTdMn
dcQ2iXyF+8kmqrYLM4GUM5kp8uPUuCWPASy3/TzEWPZr1msnXjm9bxXXgL4gmqOm
MmTP7H1DyNRJZG97Mb7iLfAhB8KakUy78vJd9HUZ8WFd+7SGj7XgMDmFFlC+mIRy
ehu2noCL5bjdGc14YJWzUaKewM7w7vUogFnqkmG15Kq3Oju2Lw2KoLVKrpcxDEuN
oUiqHlhMZGWi02Ae9+CqR8UBG66+gLVd8gjcCa0ST5/RNVGvScVsTn9fqpVA6KUo
/cYbHMI+N+b39nQDitSQM3879wzpsJ3J9+wqOAf3Ttsq625WHfkLkX+Nzjq5/DEc
xfuv14YwOqQJtjsu9JB31kl/IRh9EC/nYjrotwW/aisutaMGkFs+MbXKRWd0Jiwd
Rrs/uG5VNdHHB6XFF9cC39/TT2ccomCD4IqC6RvXz7H/2FEUfVw4g4HQIixEoYDU
Ecd7ALciYY1xbf6cPdb49mQAMhFjoFKmYQP2NrJzMTcYW/O0adm8EjHccC8UwFBB
4M0j+P5Mxvia0ihm4mhfk2+nSdsYQqng7kcE6SmZ6u0EMS0xsbT26H326jOmWxRJ
NyqWTieE1XmXkNGG5gxGL80xxqIvSJOGCWEWJTDAYtBxK4g2NQUSJMMmgSzqbmAo
m3lM8yoaOLJWBGp3o8IGb8vmv3JWiG0ekqU2IvjMG861ZvEJ9pIyVbKymFEPUG1B
uqvabyZTZ57IAhSIVk0xWkq0rFV4PSm8HA8eP5Ut0K+7Bv/HHFpZEvQyQapbK5nV
hprTJ6piJzzCZ0UELqjy+5ZSYIJXg1y8jhiqrl+EpKDha1/LaziEEMf+6PAIl+B2
JKq/gH9707u5UxfVYu/u77j6bsFcJg1/lWVAsmynEUZ8Ag91sEoTDf/Ru5jNd9ck
NkXoqxQ8BPv4uE2zeFnT1d8qvr8ezHhmbJ2t3eGnVN2A79rI1dpoYetBWNmjWP8c
ty0Lkd929lHpsT/ABEQmnKukCp2+HlZcundcVbHMArzUwKkGdKYUiqLRmWiDP9Sx
YN6+s5cQjFECNZzoe0AhxOAtxHGhqmmf5VUuDOZn48PS2GLwUzguLa328EXxmDzh
oRwyC0y0OqjgkqpS/KjGFhGJvQKG7ZimZoYNH53lTuQ0h9z1lFqQAdDN5SgC88Zf
oteYv1hQJ0aPA21KNrCGbd0Otg0DEAnvVg9pX9+Lx7o9rsL+i3tUzTC2vot6x8V2
a0tDxrh4MXOVAVz2Vd8oCCq1CVEAORL89AS6iqeqnIwUD1Cu5xTFkgJgA27leUak
r4kbB+o0wCS6icW+iNySc0cfU0i+KdAafqTGZy75EBhKZx23TNkcDajlnhqZzqw1
DBzQg1TiPfkMdxJ2d6cQ83GoScL/EnftnHD7bkLnlg26B9950Svn7qEwnx+Rad1K
OeHl/IUFJb3EdV8w48stcWq1HP6ZehJcPGDIMxh8XHzxmtooUJa9k4QbMRtpJAli
VrnbtHXI7I1tvJN5QQUcaeBty/FJ0n/HtD1VlMdA4AmyIi241V5H1AW08XtcO2WE
VDCdwlh82Ojt8kWbUoZdA0d/HjGYikHUqQTX7UTfncOB2UH7opi8qlYZ0aB8p9Xo
dwsJepQhungb/rhNLx34sMOxzwUfEoNqdb2enzAgLB/NAuEnsAvF7G8ya9L+dC3Y
C3QbLuuPxBFQIZAqAow6FGBksdvnOOqxxLQ6lmG5eKvl1+YLJGtN6kk/W2Z5WnbH
i2IltuUAnVSPe3h7q0L3DsF0S03mxwfKbuk9SX4BGRpHldcNnRf30M7uFoFBI6sh
wSIGSzk1jUYVoNazqLBD1EnOxByUmwBUK8T4I84Xn8f3B3bjKwa69gIJPyraN14L
urh4LKSAUrbaADQ0iCUHx3VIXtjZ0cl/6OFrsTSh7Q3RmkcMPzT6vjDSeYFApDmU
TCU/XLMa3MnkjS2MWR0snGtRCYbtQ7gNei7aRtcXYn3GOTQqxVpl+aw0kJ6afMaQ
8AUSGu8LsltRNBek5hb9ZGs4GskUAzNI5CQZQm/Gy64pleaklJNCw2wW3Mygjkdv
kP71tnfxnqKxb8dJJbAja2KCnEF/B3AWpe3o8mQFvinXnUl59jw9sCEiTLABew9t
uS9t+WboOzan8ftPnGR0LG1laIMq1ZbPZszvzMXQOijcp8JaljaEixD+Kv22tePB
MbehSKhinyg2bbA604nzwtCSsJNdb4S3IBnFOBup10/J8Ql3ac63RHRyGgVWWC/J
jl/KwbRosvMDIp2lyAl4581l/pf5+D3Bsdwz4/GUBZeU6pvRxsasT5F92iO9ikmU
N8J7TOqeo1X2Echd092lon3DHeZY6RWHJj07oD1fZFT0wN96PW+uCTr/r70IIFDA
xLRDIWIK+b32PNlMlV18vR4SqvPxCnMrzQ38FJMhY7ZTEd9Z537NntmTyc207r0g
ihOoL1W1Trk7uyZ2kSOl+jfgQTimhy3+2zzWD+dsSbgs4IvxDXZpILuGowbIdRVH
rX1xraXrbG9Tnf3sAcply8GtFEKSV4dUvBZwRvy30LXkVubFUWIV2y7FvGZ0ess8
TTDmBDL1Gmj11YOKkOyyUxD0qyHF1REbhjRhGdOFIVc788OcG2LrKwlxH5LLUBvU
pA4t1w+U1GTHCPrRfiMNyGYRVCbITGv/7StmVIn1arQULvv1aTB0wTZvPv/62l7U
h6mn+ThAlOLf4mh0g8aJnMB+kq5CZ+XvVX/XZ5jxvORLVnk/Z8/AOKxzD/+dzaU+
TF2V8BwlQAqvM47Gk46X8XQbdLRIadv7MUm1Ode+sBPrj/3BVwQNtLgXuCWSNXgi
J3HyeQs+wbU+2BTLixSI9yXYZlvYmGBks1U5BTTL/Z9MXDWNViF22Dve0WvqAXSl
OKPegMVAuqgk+bYi6qxT4bZU8GF+1K+uvW9p4RIvdpeYf9T74qK3fUG5gpjjULMg
C5ROD39GvtGPav9Gyu10fScxPOJ+ji3qLT6mLkqrJKEC3dHSTFg5bA+m6/zDtJtt
dqn0xiU3Y8q3NheiPsQIk82fWVVdcUzeIVeTcG1NXe4k5rQ9LeJFKsqU6E7d4z9K
s88x9s/gTEvM6N8Ii/2X0RjqfUOtttJVOh5HihD/+lIfN3VIxQ/lP3sZedu7SHEv
c62+/QDZXyT8Zz4T3JakCbpMwhFoNwBZ2gdREMVBJWCPIU6aW/95m1Iw8mje7di+
QSKukJsCsmJ2pdgLvj7ng6qFUqhT/8hV0YVkMu1vVS0ovXvjaPp+SpxYAC99s9zi
fR5IJQymuf4rk3CBrfWWXntY4TDd4RxH7aKQZVyQiEzOmfkeKDuKUpkCmn8ms5dp
0HmW3bqkzFUe/lSH/A4XE9f0jVmYgGS2tmcAcA7u9nWGw7UyJcNmf6Uy3waEW342
oc00eghI0hWLjdESNnp83kLxlIZPR5D5tSj2WqvHHDTHhXqsNnknZqLiQrbNvjI2
v7Mzd+FRC2sYL9FTNzmGGvp8GEI5QogQISoOnYNb1w1RPwL8xHsA78xbzBErM4+w
BBiRs9Wv0aHoVd52Of3EoFG4dPhKMivL0soar/c6p1TqCkaBwcw8v6jtmdmL6cpH
0TyTo2hUfDNE6Sgay11BqmpthfVtg/5i5t91wU+4kcSd3Rl6IZ4e6QiT/uM2PvNn
h9yjVZpMmQGlhOsuY0Gp6f5mJabvmtA4q7LRFQ6+NmFNvXXUEPVpi9kUlZfgSKEZ
9yRVCX5N9eBvkp8ru22QqQOu7WCXZqqF0G9RUrHs5AMTaC0PqsH+95/InaXAwPqT
6xGtu8B5kEF+9weHLxf+l8AaLCRCLhakFBMCKqcD5LtlNuz9BTgZaeOs/pOM5zWL
/x5fXWeWJ9U1MxqMYDwV/4Rzi0QVbdVMSlQ1Qe31LCDa1FfGDrRFUX3xzlcXUhWV
l7T581aw2enMXhZSOq/gITv0GlawtgFZXTWqHPGieajXDZeK9YLgrk3nLtQxpAMr
pkEkGjh0ySXG+yy/KHU8/bDRhuPXSc9G2tYo5NMHsoPXI9h1oec31XwPqrmINcA9
cVh6iLqsV+Fjj58RnAH6IR4ZKG2xAi04ctdYshdxM9rQUpT/lbvye7aF2exLlEyA
SUjpg8e+ghyhaT6J1pMDrvbJlW1cPG9emq7JQFYe/Kc0t0uKvYkEu0rMrgoMvF0c
7T2K3ISPDN+5zhBdrWDI4QdSb0lV1tWKpAggWYk69Qike826P9rzLZhmjwyItWQl
YZMqqd49Qnn3afMLanxhhNDyk4ykcc/rAKXlVq4rDWd9E3Mrv46PRjHAYpQjRNGj
CRp+uqwIEmRbCsk6suDW4EnDigPwz3eWCkMG5owuGQIrWuvd2XnCD3CS3VkLF6iv
PuU2fUHu/055BGSTskSs7UfutnNEkoVkGf/0IjIM1SLFc9y6fhkReJ046A6DWLFG
nLNdXfqbsH8PatzbSXHszXAlAlOCy+uAtdEYHdkbG4yKOq0D8fzKjsAZo/VGZ15m
7cUZJj6B4iXATZyAK52ggmAPX9WianNQp0wd8Sx31CeZBlmlyMRNYs9bsdvaT9/K
19TfI67Zckev07UlqPRlweGq8JtdJbeCvTeXEAyFVQggoAUmKDaiT9ef7FdQ6JiF
yDIc0rF7SRmJdl1zHfaTzmoSgY57Su4VvM1s7XTKmCaJxAk2noIa4i+kk+wuA8t5
u+66L908by4CcYjd/WsOPkM6qHs6vPvaxoJpSQcJBo0UK0VpzmMypij52YMJ6dh1
0nYHcW/iMGC/Hc+fggHlI9B7sjLiHBEh8NKsw1PZcAAHKI3XVggyCeS1exKALmf9
nWljsC1rTgEqXsdIzVsYucvL5MBoZB0O85AjCn+OOuboolEtnEQ8jOQGHaQYaQ15
KTnrPQI8ryPsjHvGpZXWSWjlRqMXAcA3AkNOckH0vyNk90CO+yTj/smaJTx94vZV
CuXZOMbXh+muuam1MfUiMZHcnOiv7cCMgG81ngESvuOgEseGQxm4fbJdz2MQABIW
KSkBeqppwjQtu53BQCTOrWqOjCfC3hhkOUmzmAVutCFPnUkR2ReKfcX6yGXxen7h
PE2SjZAfDWV6hC3cy5sfnWxrvDEgYY694U1f5pdchNbar/m1WEeXyRVhp6GWPyZz
/t71koEKRW+bbRsYXhViUMo4JyU6w0TeCKk3NNyvZLMIj9Si8J1zCkohWkQrFCbG
1LWJi/h0D77DPOcVIoiWGX3u1rCpBFW0v2+Ykzqke8aSuyLDP950BFEhBMcjxLQz
x9qsAMApJKOx3Zd3h0r+fg0VcnwHpf/mNzQX1tOrFUrZkN82DMtwSf5uosFJrPYO
cap7X2z3r1MC46y98+W6fyj9WSprePq04sZLrdY518ahDOCVekLMrHB+Ln1OWTNf
27fzdQY1IsTJMH7wOi+s+/LliHb8RvqvL3uSufo2PdP4CBmSKK1UeIm+GQoptpq8
jtm2yJyc91pAdKccDwNk4xCjxZi6V9u7wLY9rbnzLwGQ0Wy7GmuokmbyH1pibTvQ
WIRJpk4TEljEnsiHVUA+40GAy4KbcnHAhV6MAsM3L8FyqVqhII4i+SLCskzOkh7m
XjcPGM6h4EcQ0hTH2A4BGqbMNTLo5IOn7wKr8AUJXRdmQ9/GqAwpJ6gmGPv/TY/+
9mVFYbUBTKjlWjN8dL6YDrA2KiNdPRzsq+rr8B4ZztiXY2h7FXXqKqclAnw5ZC7U
8QgoAq4JzoY7DENAEEtyl11tex7RRsPm5XBrCUCeDA4Zvv4wUy+EorOcdrBOgBJ+
zoXJNoiHyDjD6vv0Td3XdMHeqTyYPjZZi2jm97BzZgWOA0OxM35heXx5DJQNcEGu
F9LX0v+gD3X5LQLKmZZS+kJJAaCNQ3RiCfjzkpuQR39rFnD1YqyYymKmFRqE7Cn/
A66Xqy23swuOwqiyYMSqdeLlX5mTItuZbbiSdbGKfrL+NMl0s9XMcHveepUVgJLH
h84g7nYvVZ8zTDby59+zQWgQPAnEuLhKtspu6nPYDFHjj0cgGnoBU4EaqiiW98QQ
ZzSO7WAlxE+O05SSge0nQWxVgRXktPgGXXOFs9Q6/83qYeg6ZkD8GExqvSqZsuqM
75EdCzf8XPG25mx+/U8vvL28uVRHJu1BSmrKl9RyIsPoYTfrxdvRWMg6VTyWoyjD
Og0S52aWa8LtnC6EOgJl5KEkxULWF1Yg22eFi5RwxUGYtZG0l59ykbpOG1BQAWoS
eCfBbXI1plvfpXKEJzE55dLt0R1s1GxDET46b1t5tzo5GAnUxxwzzThNY1Ybz047
16nyulcY3fDPh56lmWe71tutY+x4cnzsGaiEY/TuRm98yrPwyaJ/w67VGtGUE4hC
5PvoTi33C5n755zXEASZ6HnZALM7H0JA+nYmp1U9Dpnjy/BBFoh8JuEOMr/KHwQt
yctOGZrdbcl0jU1swiv4VDAmG0CpJtkMXTjVjmg05Yrss1LlK2IgdfdKunza7EIc
4vWzdGlUyRcVyCEqvOXrYUyKGUH7Bld7agGW2zf6HwITB5yV71tnKPfLeqxXpv7X
lSpCG0XrWFgmLY9u6jHXFEON2hzpGDRtGrcPh7R+RJIBKKjbuH+/32Wo4AuDwpzV
dmRSzbwGPfZxlB3M8G6krr7qz5+jcaMdgOklJMBkzIIddKD9ptcm0q1OkwZMWn7H
LNv6v6A/VZGEssayjyI+hO/cv36wPayIoYsm1wlUDAkfMmKS6Zm2L3k4venq63BI
0nrEEv76l8H0boEyUBuvF697o4HSsIzByOJG0tssWHMeBAfwlZbf77jDevjzPZKo
wHhBKxwmTx25pQ7e4IC9VE67QYTVrZl61IhOn05N/d0Fgn85rgY/27m4mmFuNLlO
41xz+b8xdXEAvfiOnqPTvi48LZoPTK8j1E0YUJtM9P66K619hHAxv86XPHv9SfQk
POLgHztfew3MiXY3FrBHHVGOKm4PMfmpOXWkSqmYVTTnn8cKDQF9/0O26FJJIgGC
iHUiv2jBTgcL0t1eHHIZhRuFj8RtI03mK1hW68fbE9CXCMR64BOzS9DrBtwnAkZJ
+jTn0Ab8T4NzqajhxtJbKW7pNSwlRnEuIkuPu2Q/C+6kGCMhG9ww8hw1jLZ2sDwE
XWkE1EzJUjyppeOW9ZZcN7UVWfaUmBUUxwZWjAEHF84I5U6PH/b1n7R1P6b7mBKP
gYrlX7EMa8ABX998QGkbG/T3LA+QhRBe0P0C+RAqfpU7/f0fsu6EYC+hSj+3SKl5
wAyV6AoC5OgKYY4vsnPpl1fIn6lb1b7ExGRsVaUwRApMT9F+eOzTDkgr+55qBk14
VBhLXDZHX47FGcFAUKoOZLMFFxS1jPQavn9lRLlQ1/Y/cvNFhB7ZU8VGKqX4bPWY
p1NHSQBFXzO39n53oyEs6kXvP847VlK5tlUUI7juivwemjLGaK0/iFI5IsFiWpNN
10DHuV6j9Uqm/snH1FFucKMK3hWfBdImjrbSyPEn013BiEpJcfryi0CskzHUFyiM
amr8mfYiGf6GE/VOkTRqHgpgGRnwG01YLmq9s9/qDy70aGqKa9LwE7wDp/PHyP7I
M2A0dkzt+NODrJLcJ7S5+HvwXSic8/K/uAHwGFuEG7KCSJ72xAPkjHeLtdIOzGWi
ShDPCyORBDrGZ4EuDn6SuMinxL/KDYeqh2r46cuUrjRXQB2pt0bKxTi1JfH3I1ld
/5r/N0soiv3EVOdrRgb0em8VNBsXPA7NWb5tzdXfhKlW09RNQ4uN8CT4aZI+/LvH
pdd3W2nUuMRxIy3FmumvUawftCxee12H0tgeOkVv2vE7TQgR5O8/f61B8NCCRPEn
T2qBWYk6QyDZdozJ3h1hi8cmnrxg66iWNeTwVt21nP26EvoLRNcTbqtmunTm7Qyh
AP4l5apYT3c6xP90TnsMjBlK0eQ+ELmhK7EctLKJzH9Dl5EPr6YzxcTuWxvgew6k
vX4mTagPC3eb542+xP4A0FE9f73XwtsIGFoej2E8Aw4ChJixIta6IcaEUy6dIciX
1/EXCcp+4c/IQHSmQw53etvunaJre34lu3j8DQEQ8bttmKbWy7WsCWgCyanICh1k
o7PVSuW3Y9n4kHxkFdXzTr5/fxrtUxJTitXsmybbwp6jSYK5z1QH8k0LZe2ftNQI
2i3Wfo36mhaInejbFn3B6V4YtAVZPbn7zCfrkbJhdUtEuXa2gyV/5lnd7Y1foSQl
84okVMlStj0Mikmn494rLyVZbHMj1m2OhbNT7thIR26NsVXaILzz0Ms9s/Z9MDkU
/SsrjQPJVTsT/C/xEEDRnFDROivWJFRAQew5gb6ZDw6BuKqL3rO7zYXyHymjNMTB
Cg77U+FFJTvyQT7yHZxCsKTJy4/Zjz6ritWSXWCemQtApXQlKLo+3zd6NKZiMCFY
x7xVoENOEQuaoySg9Ci/UYqQvV7mYCMJSPDJ/g1QANSW44fONXEePEsatgammr2X
UFNa5KxQcF7YT0+Xv5vkeGxbaW/rKMGvkRkgwtod+ZZ9QwkYYNGfGjXDW9iOK3qD
ehekF+b5hYo0/9uaa3Rojw6L5FmJaaoeGv4mjYK4Z36k8oxe0nwEscITR/JNRGWZ
bin3pgj/wHeyyKnqjaRlxwH7Dt3SvC5xBqFh7Nq6+hgKQAgN60q+nbolMY7Jqx0e
1LgovXnJPfmiXib4xeiEb0nJGwI1ImdPNflStHJA1nJzilrNmX64LaB2OW8k9T98
p/JGnqaOsKE4jv2RFXuVorjom5uhppgOt0cCLIHcJBEIgSDGEkI18LYWwo85tAED
PWgQ+AP+cGxhrL3VfYoxKjnf4VpiEbVUAvxyE/IQhHDGgpPGBamsDDx22PLUmYpX
BPzegV8utkaTyTvKRQje7qpkbx60onfTsPC6bl6ptGjVEv3CqI4csrKxv3v/K6VJ
17hCPvVAn4r/mlxCpdPxzyd8m08XYQ0N3dQAE9MpMZncNJJ+y4v7xnKamgkznCqo
oBRf3BPlInOqw/s7t0+lsHwbCRGS5a1wpb2WWDCqA3p6YWjmWsKl5Odnj1RXQ7vs
x5Ka/nPDInY0lCgsI6tkffQ8e+nDecPenEy3KOTNOBJWKWe099oEt0zTethh/tYG
Y++jxj1ajDRmxU1asLf8B51Hu86GftHeX7H6DJvAOvVtJxzNK8El4jmQvFJLMZvY
XtfeoqUl8kCHiPso7+MDPps8OleQhS+qbhFc5txgQjL9wmvbpeesqQ4rG1CcxSuD
roWwJFZFbXBH4nyW2gBFw/oKO3hs6tLWXvL/SAH1U3/e1gGM3WOG18KU1SPGAtk1
xOW2JslFUJgfqj5eM/aQhcFjoi3NKZiqK0e7aoNHZMzHDWb7XlzYwh0+kFx2ijNj
z09EdxqH0UqaqUUfI1/3LwGQArzwE6gmtqrAk8admR6Ti2SR8ySuZBH5AwzdT2G9
hkvyqyZFfz/qQfDVyr4n+MkXB7D+tgQcjpmA5rEvsPhrk5z6NUEpeZ2g1GlsgzMW
zSCmLUsEV3vsMoBAIS3ZIgzpVxc999zkYw1XEGaVxNvY2dm7TQ4mTmFgQE6qQkA6
TS9YqroO592xmyrUw8BxgWtF5ycRGe3XBRDrJl0FjHgk/S10N13rRrcjvKASogaA
K2PiAWQ9ZLqtF3H+hKesxudybdWpSf1epSBnfuoAZAap5DNG9W1HzclglJQjLhrt
wWMNSEoAxvcLA+QZ5vDvTPzpuPN3arMloK4lfts9HtIQ7N7S2syfLsK/MVGW5nbH
9YmZd/lmDCGMMVbxD5UoEJU5hC4fxfkxfgYIAH6xloYEB1F3GuVZ2dyFMPQmV3Q5
fBAOBQ/3QK+6FJ44WsZqtJ+gZpDkkDmC0X9aR68scr1WaVk0WvU7eoxAcxa2r0Qt
s8J4IiKZRbbgi+p6SKR+mU32C80BRayt2fo+1PYlo6M1ZpBR+aMHAfLmrmzMshJC
2j59GBEXfPQepmP9VabloAOwzdw7R7+gj6qRL8mirho4IYq6zTOWT0b2S8Q9UfHJ
J4KobgWMyZiWeB8tsovlRIo5dkAE8jGG7yxVug96lGk5ioZvtfyHK88NMVFWK4DF
0T8GZmmPc4ebrzjc+KXOKOS8cHqo7uKGrdmW2uFroA1o4vPBxXpkHIUqx+Z++ecv
/hLj5tQ8OopOgiIrIf1sobTcdRmS9VpCx39S1eY+Ob/p0yaaG3ItEq0razCbWt1z
kwE3zUT8Jh15omTRuArHjGbwoH/v5LzszdEl8793KnE2BEkurlilc05Xmfbcuy9+
9BK8LDfLmhBcvk659BD9o+8zkpTAoVpTlbOnjPx6kB/gMGF9AB4UzlWJPbwIipPc
aYc7ViooJIFeRJk3DaECfuFeaZQtg8nU4265oMp7M1P5XcXu3pDCNUBIKiCGSxtH
2CrChyrcGKHlyMJxIxMVbIsR67QC6tHdcmE2t6fOSevZfird8lSorVqXy0QE52PN
QHRaID363m7M3Iq1Jov09OZv7T290s5Fz/XLSzGvQxKG2TImWRG+fEGsFLGhVip9
/WkgoxspJD5GHcwOuRX87EqSZjUIpuyduPKrCBUOAK1kx8DNTIiYSmP20p/BonI3
kJ1rZvcSZhMt7EVI60u5MkF7FyD9nCpuWzcAFQUuCmBu7gwjMaIrJ6PwEV5+r8VG
WxYYL6olVYt7F38Ik57yMOCxpm6YVORoB2hLFxcEoUfLgfZMqy7mFeCbNaE7sxG9
G0OmZGtcpf1Ypll249xx/nniQXCO51MaWvTYo/ncdKh6OXGwLopHG1QyE5SELzKR
oWwJTR9JkYOGbOASk9/DeTgdxYYUVewoKOFn3oVNVPBZI+0+ogEu+WmO8Grgi5dF
sUtGtXDVTAcK1bPoSK+fXy22faaXO/ZqXTNz7xgbjRjnnuznfdZEhbbXEmTGyOve
0N68wn47bUvOsTctGrYFoL7vmO5aIfE5GW+/cz3Ih306gtdJYaM4qOyRqiVwfx9X
7mZ0Uusf3pPyiOjfQQZWFrKcOCkEpERNTFKlGxbpASuwlSpkEJNk1buf4h8ryN5S
YwV3xuP0fNHZnlPjiXsuUKAXpUPHv6OqAYBq9BTdRn0igZc/tic5bD6dCidrk51M
1lLypdMDW4ftFydDLWN5jDqaqcHpp+Q1xIZVcmjF3pGiHQajsYnHB6Pgzbi/NwG6
msXNIZ2Hiv8BxqwBvYmjwjQi/aoMJcGFlaYVtQh0udqrdebuHENuf5CG3qZwlKWQ
PUTA06jlMAhFku93fJBgauBkZ9gQeCa6oKfREhHPuv/gFD34vQVqtTxwuMF+Gccw
dYCiPGPlGwukffdVlpXf5MtVYoX0Pqt8bMzSh8/YFKODPCqqV73S62iScT/UVqL2
2gL+kW9++22mvi8uxxTOfukETnEFWp2G3HtXcC6OsCc5sTKMqIyYIWmItgAzx9M1
Hq8Qxqff+v6f/lawNQiTIDTxZSxcqV/iqhhVucVKx9+Ou4z4v9K/4wa8yg/IHBCe
OLfgMy/5wrqTq8y5Mqq8oed+adAhqbVY3zFojgzTZU4+xaJXStP1Z6vF+DY7bMv4
yHu2MLIDIzSfHdKZFVx8iNxqU3L04Njt1cv/pYwS4l1FWI7r3YQ6Xuf49d8RixEi
tiV/MDkRlgdLaOVnosCYDy4TPmf16t7T9xZAYMB8RbGJ4JDZXV/sJGGZ8DfdK4+d
0pTR2w6Aq83KpVwUotCCvCNOBhGjNvHXqjG7izejVN8SZkSYfajPPtUC2BAFYjrB
HxGIKcf/dS7t2ou/gZWvLVmkcaXKhlrNmAZeXBGx7dFm3xcDCg8SBDWvRvOq8VMC
oEu5IJB0Hz7Cm2cawuI7BFf6gCA054OC3QkBNVLM8jiDjxYgc9QzWIVReUCLRtDJ
5cHZ5sw5FSFyuoQiN/bU455VeFHSviDqva2GQFNQ69d7HN5nh7IbFbDGB5xuUFZa
tgGpTE8S/dFdPggeqx2vn5r3DBqckKtgRmzVkIqOOxRg62rIMMZmS8vcUwt6bq3+
4c1ojzK+6CrH4mXV8A2kCAxxzGimJg7yjMDKIxPIEkcEKN2qkfKC0DHawdpfzhto
oq43jYhLJkUnVyhygJG2bN6FIb6aXTTV2nYkonsz6tAdN9l9+AleaO2UNdMCBTXI
nDru2NuvBuxLtRBYL1n/gKme+I2d3WT93e99sylbrU9k/+KK40HhsHr8rkKymzQZ
AuE7qY6aLl8iRicrxxUiltMWepCqnDJUic1bTm0xhstiUY7Ve9L8l/XfiEkcpeMd
emcUIKRq7QGAxjbY6HaSvDU3Fkbxevpa89XsIkUkjiQt/e80arsCoVKDYOyY9lRM
/vanx3bF1RtZKQFrLB967ifbJ1n2FXJ7hgjUhyhLHVv5cOzkEDZvJCQ8JrakFwMM
ahswLR4/GuRNsaK6TuPOG1MadUdU4Dh3Q+YwlnJPG0iU8GhEk5iMJrbHOzFDfihi
jCyPT3QV73kdnBvbhAmbCYJfKrgnm9MTglwHSSNHmZPzyLVxzWUuvax0q/Gn1vYQ
tquDa4VQE9P8ssa2dvjOuHSZ5dov8cRLR3xQucdfy6rHEvLWyGCC2/4vH7Gpr4Ag
yG8HoIbecofTpdD7BIhaoB2891TFb6TU17DR1/2cVtCczjM1ygvmKLmWZEErrhq7
4+o4P4rxPbmQTc8sqHcasJ1Xj7PlPVVuRs62hDnsiA/Z5LqHlmIi6bn2eUQT/aKO
xLscHCr2xG4ISJ1gSResND2qedo4GqmmbU/5jqFRmp+hmVsYzY+REsOtwtRjoLtG
2p5mDJM2EWjapwwfpsti4unK+kY2L2+PJVUAL1A+i0Dm7g9aUfgeq8gYlkdqgKir
C24Dyigb+dzcxvjrBRShtIVeHVupBDaxgWnCcJvEUm5PeRws8uTdwd4gmqjerx6T
zMWT8AYfCSKlAfETWo7evI/HW2lt5/bzf70lPHkU/q9D5UKAp+EyNXwe8GHyZ8dN
1iwqIsANV1JVvu1D9GoHssEkrzqNgfGyhZlaDa69FZIiVAI1v33aI6ClEVw5wHu4
a/50KhdeYJ+W34oA0jNOM79hRkIvTow0eOgOyW3+h4Zu7Xhheh7QV6w7/aOfxOlW
+TXR3SCvtA5yOWFIrCxY6Zfq9U+fthlJor3orbpH7VBGhJG2Pj4iQysjTUiZj4M0
DmvulAJzbUyFvUEhvrdQECBx4jBCChOW+nM6/gNWztsFnviDEDKSmBfJoBC1xjkb
tgDSKld7Y8hcrMXII8hGK+Yova/5cLDYxBQajaN7XE2oRbTUwruPYTfI7wrQa17O
4mfy1vAjfUso1LPxsSM7VLTtG1ozvGlKQdpwMm1/gSWl8ARJsw2gPZV7W8UHk2Ek
jjh/ct912i1buH5+CV0A8AbGv8bZagy60QWeAXJ6heEre6eqE4gjRQMQEw/rEh46
g7Hzocuytk3Mw3aNW1UZIsgBxVR61/Cho3M98YYaVxh4l35sK1WeslDMcQ7VZAYw
cZeVYmHoRGw5v1PMAEy5Tx/wiQKgcmqHNkMAMliPv0soQAMt9Z4n6Y/maOZMHDh5
GOk8GsZnruudJmlbbDERMeZ5UZfopd4tAGygxidkdgyo5HRuK03qjnShB7509sUi
BoNQYtyDyRKzisDDvJ5io7kLkjAcmKrLpO18yXCsFcL/6NAorp2yT+qy0GhayyF+
N/lyRhU+vJWdVRGHcMMl7fqImH2G+1w3V5LVZi544kdRLp2vZIOd4Ebe9l2tDQm6
75C9apINWzX7ub22WxNDuauxTeq0HLhWM4T71kCWw58c2JbY0MJdd0lXqOkob+05
hk63vWu/dLqiHu96umQpbMH9tEOnwQbUqayXR5LIRzwWzVbDkRvvR0KfGZHlTQa4
PdGJmUeBR1ovTT7v/tDEDaWp05sfped74JWd136ULNBDqUVZ00/uTLQ5J7rlBbjw
CWmfzOcC/ZLN2ZkzmVHrzrHGASgB/E7hH62OUNAG/DnqtBs2AREck+BIQirpc5xr
9QXmELRqKUndpjpVCB3v4/ymmRFP659fVX9pV+9Li8EV+Q1kAbMgm4SAS3sPgOx4
+q9KTpCKVL2Kjv+a7kZnnkMpOA5X52GWXAiaEIX5XkpFyioEcwtcok+3qJSDZcS9
SUe6em25GSbelrlfKGvVXTS+juC07t9icpoo5bqDC5KrI4RxCOvITZbqRWGrRWUg
8UtuHW75Y5m+mV+2O/pSqM5vb5P3Nd2ltbK4uDEVal7KQvdUBWrs7nmzj3MOJu9n
fWaliU0qqup+GgVw7ROS0IKKZx6U9vjL5m+jQeuH/GSE+3eiD0hJjSrD4Xg0lIJy
E0TjfdwN7HRImp7gnaBIVa8AxSJHZ7hUjWpNbHVOcBUR0F+JWbSSNLlZnM0ubiSo
HBNeFkqqE6F96D2JUO7z/NuVdyx3IA+Ksqeif+6vM+K4H8yLpyn+GlV9+B7fW0rC
f8sKmJ7/+QkzhZlwJlKSyzwVXJEZYoTzWTnyI2oapu29zW1UHBHpR2kuS7z2CQ2V
vb1Do9BRJx7kLrbv9iecvQdSNNrB8gsRpoM4BjZ+xp8H3W25k3xMRwAquuM8mf2u
mWWbdMI0oLhTQ8NSceh57RuLxQMsCiNnJLC6HahLqr/33O+zEqzagIAYcym2+um4
fJ9BpJoQGH7ZiII3KCrtdSd0SerY0q4BkSPWhcO7KjJ2bR0PidmMsKxAKt0v8h3y
/aXUz7mRhWhUuHqxLM9s+r4BT5TAHRcKD5hh8qvvqzDnwCkf7qMyyvmzEjnrLjOS
rLqoROS4QfOdpSZsaRXO+u8zwvtEFWCmBUcKqF4TL9Jg+C+QcDpUp6K7ZalUTRsw
cQz3ByRAYc4wnU/I7bciqx0uhKVpuV7j572dN6JscMYR//GYYcz52Lp2G3Am71Zd
Jkx7nYNXwkZpcn1/fKhDCVADY5U2Kl7Nje7oM2UBPcBrELNvgnWK/NP0A99SeXek
6BimdO6HndrpBQIVT4IN6W4D1SQJZQVI8Qv0hlt8jR7fOVvrS1krmMMsYVGCjt9D
g2qHj1vtdTCR/zHXHUYFZH5J6noEyHM4zz7p3hI2sHAzCPkq0C9C9rxextPUdK62
QLIjcuUs2Q0xZ9JXBQco0GFhceEKAOCnbX8HqXBGivGopt4TeMjpm50xgAOnPa6E
2gLjXgySlqPuMVZBIQXRxYZUe/2sJNEWr0CGPWK9gNkQ8I5wbGHnZ/dhRNLXwA+I
byUVz1YqecX4/WtJaD1vuEHEa5VEXRRfTT2dsaEQ8wBa6V7/CjTlIOxTctdLFpL3
D9oCEAMf6/+rUvTuzOhAXv3ikZr2DTSswlgwK5Ch7/VKPuHhEjJ/FeQOa4cRVkK+
KeBGntW0aEY4Y4W0pL1ffXCVK2D/ed5D5a+Bqf73VQF+z7GJId6vCeixi9M/GoXF
XGcQabuje+C3G/1aHcnCL7ik5wmU3NefsvYc16P0TFUNMCUgGjApGtiOy5Zqp/t5
8MPDlLIZzLCUH2n2QxPBoDdsQ4deBqrNX0JE6yhJF2k24DnwfklJo3lsJITIea2W
Kmd66i8wJOTPLtLNLwDE/PDBygkoGWqAlCtY1c8f+oqFtDKhkVNkfIF4yZnNBd6j
lVYQF1fhZ4Puwx9SDXKden76MUEv/zYHkneT18V++FNJXY70xC8iiHpo7Opvvipg
CIZB6dN6SqdanZnCgnMMLqpanDTb6TEqkK2vgy3hrOgpJZUY/tn7a/DXQmmkIV8+
q84fn/OnifJJURNVMLUzbCNKzBuT9ZW3pSSc0BLtdEroH/Qh/vESU+eeD6LFllUi
crtweVrR5uQRauiZVcCG/EQoyKxmFHa+4fFxvGzyvdlWq+tsNRY8Z+D6kqPA51DN
MprZ9H99RBq2S3nsOkbc0mbISG3nKi0hoBzyNzUt6EFivRe1zk4kNVk3SFQqqUkL
5yKqcsFZQ/vAFokqCrC7XvE/afOJUEqbwtJpIHFUGo52BShzvmuCa87jAjbScMfw
mRf7eenL/RptYxvvwwSzxFDrqlmDdZZ7wpfLN1CYtkVRz/8yWojyERJqUjg2Is0c
pAu6rSV3IQAlxGqpWTiW4oupNDnqzFFJNC6doTEvFd7XqdgcpTu2fPm+EzwkDzdS
bCQaR6E79TXj7U8MG6fTN7TyoGtbYqHZiPPXYpTk9fdViu8/KW8i/8woBQAQA2kV
rbklkrXDHU+QBFMCrs6y1mQsR8fmjb2YLEQIqRTIzbxI70CItd7kpr34mEhKlzrS
s7AOTPMbjl/IpJcP8z7Rvm8QJLSulce+GfR8ltbzz8amj28W0x8Y50nDj4DV4XPP
mhVLEQTNArgNzMD6GoAvcjm3O1dp9dF5j/hsEo22XaFLQ+8cPWINRRKcr6clsugo
gxzgOfTd+Q+YDRbP7FijerbudYo6faLiegXaeC0coYnzPlRso4LUZ46/h2EbldO/
MCTI48K2HfaDMSeQqtGj+m5IpwE7EldF07JfhaIG0kMUiWDkZc32jjwvS2eskPvE
bSb1Rg7HZmzxRAI/8tf1Dj1YteofqJPSeIhdMFMXvS5jcH6Mz7Xev5W+FzNmDUpK
nnC6N1lNWf0NHduusLr+7W4WCjrW4inlLI3go6QaZSli8lRGADVMmnOFM3HRfcRu
HTFQTPl+uKD0WIvp+NFmTeGBcg110DenbEQJMZWmnqMnvVTS/UR5i89KCaWbmuE4
isRrmsFnDnMes/IxzejT/DXVhJ1b6v0ruGVwEhQU9GgmxTBYayFHpvdTc9Hxhzqt
sqW57xIyXvx5vVfxQM3L718Rg0C8Es5VrKakLqCdhFbKZ+zXbDFXhp9m+QnwihhM
YulcTbfJddcwcy/AeG4nuxdf30zhrYPdyGePX1S694ugRxVw/p+HLj6mlQ8aFKHo
AbLMVK8sGQN+ffbnaM/0nD5q0c5SfHRn6eqDjaD0nORbyH65iUv+PpOYU46RF7EX
dQrxMSQ/canJw0FpCOMAdswcBfBk9vyzH4rbvStMyiACRy1wb2pibMmsxUbDFzh3
X/FYC1ZC6ZAN4GjpwrT8BF9SGZNvIpPlAGUxeeEoeufjetVnINJUBMV8+CLWnhlY
13SuVhtWOL7r04FbAaQ2gDA90mx7DUg8PDSMXZCBwnV1ND8cZBF6hDuIsDOUEuNQ
sD72D5USp4tImFsYd59ZnZQc5geN3dLz9trN8bPNroIlxYa4o254NjcL00yZp+FD
d3xg7REOhNRN5kl+OptRJPU4gXeIUmeWve6hwVXE1h+4gf8v46xbXJL7+UR+01wj
wUX3onFfmypZj1VwY4HnAFi0T3muz/SgJReMg2hdpsEuDX/6UpRli2DnzavaGy0q
OCsnMIVZ4aDe9L4NN8f4cCYulvzZuG7jZElzCiI/tsgh7gTw2kMs/mUU3WStTmPq
l8sF7u4jgd+2Um1a+n2xNyhUPve8sAjO3rpeWUXVw3yo6W86n6c1Dj0FLUB3zXZC
JXTjCHxtEd1c/6r9Puq2XPyku23wwyrCoKpHK1v9F3zKp6nqgKavPrjgPD5gFejB
wtVNfOYbTlYTOtFOBGxTqZsjKwVe6VarxVvrpulrWQRHf57jMTIJ93HC5TrEuvYH
s80PuawoIlF6Kpq8XVRIYSn/c1M/1i8+pYMSoTq+49eUezNeRo4U+f1MTNaqG5BG
RBUFWv8JZHTk3o6ywGizWbnlmAI3Y7Dn9hWbz4y2h61iA8HHzJYujPEeSI04HNw0
3waEz25i64m+x9oo6ufHlmrYUElEz7e3tCC7A9PtBThLxOj3A2uZeWL9zVd5+mUx
eSBBHEmhFFdKPNRYkciZeoW1IWrR54gkjNltiO7o1Ww2WbWnrtObu8rfgtUol0B2
DJMe8QsTLW4jlm1Gjw/UQ0Xk0BKBt4DUf41jGqwcSWvKAEJqCGJq8m/cIVutEoOM
t4UcOKNx/IrdbQqBHfj9PKsTFviMkNgiutCup6HJHK9lvMscEkOWs8h23lj2lx9D
Acdhf5tQJ78LLQ2+9WSgMrbzjystKoyoxbZCXsFmQMgyXoLw1pnkP9yw2zxeEtVQ
l1rgNVT63Rw5DJgetLpKNgWAKgMcI4UWf3P9lTSpF6tFJpJilo1tkMzSKOf8dTux
giIVuoai877fP3nDttSFGCJe/rRre/5HIxdv4CIwmiW9V5b45FrtUnmhO4WzLCrt
ZabrSksS374iRak1ruDHpfM9fxsbrkSUhXGU1FQMA36tIIwVNlO7S/kgg3f6mR+y
xSAp1xfJ6kNUvAfAh/Ob73WcUcGHzUc/iwCErJ2015FWRI4NI4Wr6TUfuS6FQoKY
WDTFYgT0NgyrWxoTi6ggQPgpKVfhr3KT6NmtWdJEPWskqTf0nep1VOzDPgxV2R5Z
InBFUkfyTcy32P/lgqUvjclaClWkVRFACVwu4N8vY7a5i5zQpKr/gjIHSDqgOHI0
gUC2dBRPMYFrYJX3PWvw+KpBDKvtZIUQ2GftiHXglHeRQli+YIcAi0SMBwLqR2jN
nyan1JK+lREt3SNFfW14pGOeMdNZpklVZtKfXR9m1peluROD1yFYi1aieY9nyn7N
Hn51SFX2SDvsHD84NLnsB+tkDci2ECIIf0ceg2vMlQRmfRMwnnoVtDfS4PFm2vbE
50yDy2wZJMRZo4tdDQsiowrYn+OmV/CpIyHocDKLrvFMihI5i24D6hw6UwcSfxil
v0X1zkjLE7vmCeN99oM9yPduWXaQozeeT8GMGu344GIegvHeIvN43ubCDlwXWuWp
dWtvFfdQXErkJEboTZ/Ij+1868K3rwcPwzaheAWpf+ZydrKtZ0PluPgyxKDEwOuz
u3b9WQfaHF/FqPwCDFXlrC20wZpmbxVS1jC9oPw+0/pcYENqmSrVxHlFc7Az+Kdq
6rlK+p9nohpvZgPGfFkZ70XBxKCOojr12h8gxX8LqirNFPCAV0I8UuMl9AjL6wG+
15lxKR7ngAbpDFRdlWwpM9AXf9mrp8ZAi/AnHEOekdJ2KhrlMtCBDitPoeQu967E
NZH1X27+8riYxdy3jFqZl8mPWGNIMueIKORJ4wQH7lrErkwUIUojGiThrG7DcDmR
bxfC7cbFgAIUDke2luaCjjHGPfDa3sWn6YYV0VMeDO1H2ZNkeguXIT/Dl93pW+Ui
zFD37Ol2sBge0NlndpTGRVCPtoOtlVGKsmy71FtnwqKtLPrv19AmQQS2sZInHJGV
p5OldudKdE9BJpnJ4TiozxSXqyCYoLPmE7usmrF0vNftG+XP0rO2SDkhRTeRB+nx
GDeToypRz/JcGhtJyIJdmAuq9bBw/VcdGsfugSoPyzGIBItdPSTazHiPAlMOM0W/
EiHlPr/tpPTDSicYVFEuFLnyk6LE5Zyc8j9IR+2Ql7XZtNIp2ocLTiDgPRGW/Xqz
/eXvpYaQiRwCfb4TeBqug42rvr8+IlM/c9ugNrxjW79Qp+8SF+vig/SmFAQ3rvug
RAY4/ak4PvEeje0yM2SG4VIrVQmFxigBftxIJ6qDOq4w68jS3Wqlb5LGAE8P/v10
uOy0qznhUqyZMWh2mnNllC8z3auIUcT6f2ByS9NkP0TdfWLcjEj7sFvcQcoI0x6B
++rZybhxXOJ66veSK26OGi7eS0F7ad8mCg4liZmAxmHKfZm4TkOQbif2HLegV7q1
Vp1aa1FY3GWocoDasSg3eAmDcTDykRFD5iZyi1Qg9kOO8Cv1pVRPSMMfnm9Q6dMt
kk8JeWW6TIiGB3TaSZO1cgueaP+Xd27Y7RfHYauvDgR+5otEQqvYvrx1hKqugrAB
TNL3YUHjoUxkCdWajuhr4NpVQHvMiQ2NZceIHkPdHbblGzmKcHFhnyze+1rdhTPe
dHGlpHXQ/IxariQWDqsdJ3aG2ew4TLeaEKKaVzNvvDQ07S012uVIJsltJJeB+uAU
ZK+ioni0b88poUqZaiPxe0kfx3hkSBMdR0yhk4n1oIz8e71nv1OjHK0pr6HzbXUj
RaA75NjKCOIy+ew3Ovcr7Dzf4/btWtRTtdvsI1HXzHww7Thwu53WFLmqfFDsn2zg
Giz2eSqI1PPpa2U4LvNEuqnfMfRbOk/aRiw9x2FkpAqXggwtvN8CegHy3/cmUd3x
TY6gEWAG9UBTPnG/5QxGnhUmvXKCVUzkAIfwU/MpbCUIlB23NIiGE6bogZpv86Rd
8+F2DtlgRvy/AFcBFIAXK6Ti1l24j7aWwDBfGHmduPierN9/JC4cWG//wSXMuU5s
upjkisu8puZ2uyple85Wic8FgFAUBCKhuMwcts3OoAImSW+jMggDqTtX/N9ZP7Mo
g7G7ikrZyUYgQSrHLE6v8Q+iSjXnKHFLX326e0VtthhAp8jykPfDZZcA2X337G0L
zvSOs8xvycnfKd0fdJ3RCqlGaktTUY1O0XIgYcktmfNrSEe1c8E0upnN4Ilx+Uau
gcPVpPJ1uQz/8G3ygKOfDnLiJ6B6rQKKHzKhq3cJtkN1En/LlO52JCDAxuXcylZj
Z3G6R5Tav1POCupaBFoHZm4P3Wskd9rDcZJOoFzxPCjJ5g9akiScmjmE7B8gpCFN
9OSW91aH5qIEKRJZVk79+jbTrKowTK/ve+EaRGwpMj5zs/Bp985Av8a+/QDpV+Mj
NiRdYr4lMeXYrk6hAGv0XcLMaT5+fKkQKtryfGx+EiiIQJBwnGBE2/0ROLnTmc06
v4316fR15UFU3dHd2rDy/+hP3HRJcLq9Wjkcc55fM/UFJpTRGL3iCf/L8n+0zszv
IF+l7qPSfJ2BL4RksRJr7apw7jM7HxCuprry9HoxqIavavpulv7A50OlJrDch+Wx
cXz8UFCAlH57VZfbx5eWyvfNYkAaEFR6hw3P/qVgP3UtilHYAVweT2nzTxFNy1RU
DBSLUWQ3BGi9VvVGDZkg5mQ7sxFAalZN0yjdjwXCNheSRTDqD+NbQidoIc580YGa
mZLPtTGjTdbzg9rxHbW+hZom7KaRiiZnWozAf4gw/6VevlM5l3ly/UF7M92/pspP
tX1oyDigFpbyShqVjFBEZ1blhw717fCApVCNr2Mw0GPKHyxUq5/4r1TVLqlwBw9y
ojSABvrtAuugK6PzubqphJOZtRHQc6tKHKSF911gH1OBiMBiynKjbWnmVa6Nw5Mq
0lY7mxGS1BLCV90n8xVkNlLmcERwfYJW0sMTw2EzRxPAA85V+ZZu0/yUXqqiLkq3
7lGqC9O9HyftFLkkkryPp9lN+eVS6rwLOBAn/45UTaAXt21FcXRKwlRwS1AWUxFf
YXPhFfNFD/tf5ZS5IqYhcTpXbDkGQyH35xwTLMo3I3fGdD4cGkC/eurJeJOJjf9c
gDo6EZxkYYlcI1eUxU6RNtjLfMT6R95U/9sZ6I2ERQcBXfOPc98Uh/zGL/EouPaJ
/Mj8C8c4ZsRvWYG2w18oFlYlPffq8Di2CaGMexNFWvJjYGAJlya8N3G1hpb8YVaf
nwjz1Oy15iEq5V4UwZV8u5pYfHPRMhfRdDvT0iHezlD448+OVGBTZJfkPpc/2Q6j
uSXB2NrnqQ3AtoDYNVFEV0O5UuQyBZgV1H213dVoZVyhSW9S23/l75pkI+SY69nf
dvqPX3hYkFw8r2mFZjyGu8UP70HIbEy7/3eMdx0/BSsMRFcvHkLKocbneyORw37P
v7QL5PcZ+rgJmGfM/sEsMVL/EswayyXSIzEJHqjfM3yTAa/YHZIHAq4AT0gumXog
6mfILEvjWiJINhX6zhpkCzEyXbHLeVp+2p4VKspBzXa7kbW+p8+NnvpKgfLOWCwR
F9hjueknx4GGtR2eAc8JJEsJCQ+KKDqEM921XZSzn/4OwkhQo4KRECS32UG6XaSI
tk8qfrE6K6Nf4LXZyaKwOhGqjydI1fwaHVsoXRGAWiPntlTZKvWi++XguRkcf1j6
Ro/uO7A60Tq0I4UOOjj7KV1bN4gGFfNI4xZiA0y0I5o5kP2OUYvTxwdIg4aGZkEN
vQk+EkA2lJz2xaglm1bJYWEKJDnjn/7qD7BJDeTijr+PjcaOsE6HTTaUebYt/n9Z
aUY/rlWbGrclZ5T2FZXkROQkpLYofUS1vIjeaGoHYAMmL56WJIMisxWCPyt2AGpj
B81XFFakMzatJZYvdpIOM7vNoXB/U9OzpCkfmcM9rILfKqMvpgF7eJIdjWuF2D0H
RNWatJKcn1+ACySXfLejcmp7TY27D17wjPwG3HCTOUlJgnB3gEWoi/7F6E6lQ8nw
bsytzHqfsZHOX3w6KxIHHHE6AbrviKWJh2Z2+q8mU7aDNnR3qg6BtbSPJKNuEt59
jP0lUagDSuQW9/p1otwdxAUfME2uoGottPN63oFNHbPApAEIG9KsNb1m+oXiKK4B
vrmlR9RQEMpn8Bt7KaGfjqvSTKmxnsjlR9j2sBmgU27DVsnGZmwi5cj4gpx8P96R
0pGW9r8FzQHemuzS5oFVPLpvoyTzeclf0V5P8GIDfQ0H8ovm4XaNsyu6GL6CHIXV
7fL6YN+uwkd7SI9YxYJ8YKlRdyqeBLL9gTwskMNWM5AqOLC0D6wJYxsTz4wKP4Ac
SmOsFyw8UHQefCcOwM67p89VILjsFPfMxNEm7CWe8/x1HYtKZMefrXDYm6CxWtLs
gqu07/Tn1IQTB2bbjP16DHOBh1NoD5/V05aYWbR3A5iqwouoUkCFFWaRV9KAY2ax
4qaiKLde2C4YEkaiYEVO9OBMzvaibGzKDx1EpMehsVPD+q3C7TjqKVxmqSiZ3bN7
xq21tlyiAv606CnwWAlJZ75aedGjhavMUzsqu4787CALzzDsmbeG0YClKTABhSNz
zJF0FkpPdyyJ4QtWHezlV4UzhjbEKN5W59G30CYwAjSvpFSi4/a+I3SUcenhmaSk
Vvv4bRaRsGxiC4rjS9DlX/CXP1UwHFgKYKAO0rPUHlRVVnjOlnBY93a90XR4WkgF
cinxktceA4w0lOewxcmyLLg1MZoa/QD/5vDoviB1dAePENVpWc9kpKOBH1owJSYx
ZB/mm/+ZDhOr4zNHeEGz/GtrcTwhj/Ayip+GiydiHz+p5behEpOJdS+31wiChpVs
9ODA9Gk7HtHZS5Vtl9hNgZXMfH5U/2J7pk/iLP4oXo3yKjxStald7vVRbkBHqT7B
385LuRoGcm0/RYXu25qrNTY73pqGeQ8Fi2jBby1MeUey0qyzpSy30x5L4RnVQE5l
/4t0AXlXbp0F1q4dPzCaj0iEzdC6a/SbHoeiJZUnhw59W+9H117/I5FihcNrIg15
8x050ekPiHXTMlRVJJDoBixGXkLnKqbRHeh0QItQcYhp0qdg75Pj3lQNeCwhSglB
NcMMU1pcOJsHkfa2eAoHbT6vSiTmWrkR0KMu79RTUXPSeqS1RM5KUVWirk9Gp6tz
0z0/5Qf47dzItEU4sbfuLTjhKb5eNeEjGpZz4RdROm5xE5h1TpAcsEjv4ZnTGhDM
/yxn5owz/Nr3kE6R+romsW9YP9ToJr9WOdWFlJm0VTOLV/QWVm5PESKHgYYfeCUb
fBMSCkjedZFgtUfTr8YAsMlxx3U5Z2bpTPOE++93ZDkOczXEvUvENp50Jh/KWI5U
uzcdYl5pk8JlvypycBAsZmnNly66hRJEfAzFvs3xxuZMhkpkQa0j5OKqDPw0HEzC
W7utzcOhBwpQnd0aFO6OrOeNhxcEwvkdwl4VTbjyS+FRj+MNwAj0pCmmUlKHJotl
BwM0JPUulUMRlP17x6r95oUFoWLDH92XCLrsylHO1nNuRs2e8osGhDo9ZaPwRRbz
pXXngWTM9BgEIz+FogiZaN4y7uQIMkkeDlqCoY91KEC8mI15QOl5ZybP1W22DNGZ
sb62hsE5ew9tqJ7iJEYFD9r855v3W2iR94lSdQEWWmUosbA0ke8sUOMVq08J60ts
v2F7eKp+Cg13xYTKeNNUr/Mfjza6SOLuG5XzHdLXZv0SLNx32g9dkWmk629lHuIN
p4U8FOSoGgUzmmAU0H1xRPY4VQhQDeBCx18kkdRDIkUYLtCrp+NojF1Hf3e52cck
Hm1wnIgZZGTlC2PuHDp9SuVkUP/5olm6sYCtfYzvcFzovBvnVQhJoI4xnvSr5del
4FVPLdWuvYkkj6sRESC4Awnh3YvE5+Q20T5sa+XLq72L0gsL2ocUzPC0dxuOxskf
MaOVEkHNlaaRNwXBumOX3uDz7IzZ5kf/vFN7OsSFbALtWic9IkCd6MEq94cHtwjG
mHhPbpw7X4L1HPlss2LEaP/V7FkTlOc9zCFVF52ySCFj24iaJ4QHrxeFOuGmqubW
aVNmFyiboYGdudAC365iyJie8y7jm2coYg+v10KvdYlCCpOehjbKrw2y/OGvrlmS
FVfcA2HbLY7aLGkCSvrZ/sTryvxFnYZ6nRdpuNWmBsrDRYmB/m4N3K6GuhByXQ8M
oPmnU19JrgTAahsLW8gdY5vUCZJkQ30XnGQ+yWGndIXunfRX8VBOT5jNTyEXhTf8
9qxxX3tyRF+j6WFKiSHawLzcLwRLSVFpC9POxxW1dXWwv1Pq++wnSmSq23cX5ig/
cg+iIHk1W8FOUlN/KX9D9owxav8eMbVlf9vryiFDERr2Qf3fJEcZntEikJxz1KOs
+hhUbR7f3u3jkUQnsHOfC2sJ2NlJBZrfcfhKbulE/dJ+jLkZXJYIQE/GtLUtaZza
+tl1cX0/iMAJmH5ybN7ZLsjuTo4dqb1M4UdIeAbEk7TACSuVeuYvrXhjtppcESir
LwZHIYDKxFE4wQbJUJcwkZ036PATKZdO1rZIot9s7UzbhEm2Z5mJ65t+57/MDHK3
p5aDYsgOUwLoasGQl/ZLyVFZqsA16Rq1gxiSosBWknyAJCp2MHrgWh6wxQhvwH1C
UaeU7OatvlQ4ibxmknNZKRLm3fEFN9CZPZbUfSJaakR4eGpIW+/SwHXqWqAbZ0Yj
rPGjH4DLxG+shk2xlLXRoPfkEwUUw/OC3JF/lfccmc4BLUsy09hLzMDMxQvQa2ki
q2l4zyHrPzgwvrc/rFueGIpijwgeV/iit/A5B/6yup7uzOglip0Zf0VvGchRFIxJ
/H3aawtAwLKSU8um+xRcwzpzMAhMRtajkUEtIGJJgJxVP1vd7HYIGH73T3vDTZ/O
iiFcEtXYwmpSXckQZX8mJ1Q2NO3Sd/87iJHwCTfEU5AQjDjt5jhZGCzqG6RV7gTU
yxZLOk7+ZL/CDjfl7ziVbl6+MJj3DvVwjBy+jK1t3u10sdVHT1L5w8EVp1a20puk
ueQKqqMWh/57lHfqelIwbote8d5RA9szl3ntxDq7WakTTHGjLzCw5qnDA9zbT7lK
MJDwnXJboQ+WJx2R+8QemG/FF/g+PmNrjm4Pdv0TLt+hqQEbxkbKO8sg7FuIz782
TJZ+4PM9M11xQ6cXaxmllSqrhIC57NfWWCd6TYVBJ/IWDooVlMWDv08crSpUZpge
ZqjoUZZNQxu0SeiA4OYoQXjaYJG1Ae+HI5PHd08KZ8hEBa5y7W3szlcgPQJDqpFx
pzvNyNKS0y9B+eOAmRirQvBoX7o2fJ+emTMaizVRN1c0pdSXU0T4KsQxf8xZAwZr
Gj//PkysOVcVqFQzC0+OsZSiSNl8OtcYZSf1EJjlBPO8yixRZXR4ujz3a13h5ODA
SJAzsJIwVp9oDDma+LTiNuJVBGBunkjAXipbSYkOQ6q1p3/Exw7YJQ36i4WmApkk
UHrs8so7umtospT4iWrUyHmdge4SUVspf7NXw1PgQ2s4+AnFS5Us0GVJbiLwsNM1
2d0UvA9TEWNv8EthngtFgYriDLGRsIKRLfnlIG1Lu+MHWiO9tL5tdW58OTvnI32h
6uqVTg7ra2MWt7V3rioeB7DK/w36aDIfmq9mHlNXad1k3b3RlYfFRcCEqy+mpFJj
5ouwzkgWsjvu6xgFtJJBxvZasY2JXEjh1x8OZIOV6/aMnYvHXGiJli2OtLGolvJr
t6e8Vod8FOrtnvQxDj2VRi9pHtbDIlcCLyHVyQsGdCHz9sOOvTiLLu3Vl4h8g2nh
njAxU2yydbRgVmjK9VmFPoRzrorbSEOlY/5Urum5vNRoUCbuMxQJy8NMem/k14qo
1j8RyBrHNt+62wWDwjMsgBnAjmCVcKYdnT0+1APVnxyY6CXpjtnN2TT19D4rpOJs
PRhdObLlbGMHewyJf6jaKc7jXYPE5ac5Kt6eFeLBt9sAwMK9u022WAJCxCwumJNx
u6m9lE5IRpWBBtu0gyEKej7JuXi7p4ZnA1vw1PR0qkf2Wk8EQ4/JvtBB0ewSfKI2
/2IPv5Cvvhe9aEx/mwmL7Gp/OjIB95fhTUXTC8y1Rmlt972eSbbXgw8ktRHBt1qw
f6Qo+PlaVAXxparikRtxHXUTjEA+wr/ojiKuBg0RC2k4FDQDHsAqVCCQkMKJD6V9
Vlb3fL7KXEsNjo4PJmETsFjs4zVVKpB04Avpcl6/dQrSBqJGFpab+zFCTcylKb+v
WA9a3MH7t4kUr9aOffYKMmBGxzDX2T0gg3FRO1uEaR5MKxOIF/weYumJXAgtTr+w
LkMlSF2LHRbIb/uYZhFNSQJcSTnWZ3AGNgHYWw4V16885g0LAxWr8431QuYqVX+3
mudHgmPOmSwQmtQ+c8xqQKdWEU4WcEB+Gan7TVPGyBwjLWTf0pcxgRaTDFMpXLsi
W4oYFgesFcT3K6LF8bsEJsTP99W0punuC7SFtEYNDMuFoZwR5QIdBW9yRrs4EXda
/mGkY8JUiocRshxIPCnsfPDBxH9svDq/A7G0kw2S2WE6APn226WOmbT+A8H88Me2
O1HIRSf7LQjZWEimhRe2o50paRxkFuqytqVTLmF35u/z9Dc0eugBjEvAIp5nxVXA
8xh+s2+pjSMS/pyVX0MBgSsdZzGZkfOtorV2KJ8aM4Y6IXl1QrJmqy6Ifc/74U09
HsEsQQDb9KYHokZYrNtA4IEdrszG9+nLoV5mbMqc7tmz5cK9wnij0mxj3g5IbopR
zBpKvo80W3Tx7vXYWhu+so5GHkbZ9p+LqnlKxOqaumhMxn0L9wGJrWTY+o1FQ9Q8
mYqFdDutKZccKjyrptd4X+mS027Ly1klng16y0hPR6deGtM62WKM8zZcKbBgWG4n
KQ2AjvOsKcJx+IzwL29LrmXUU1BDXkKPbk9kAa+K5o7bA6Z5QkaE31NKs8IrWN+X
EbzdW/LfOdMMYccQd/rSgsTfRSsmNhezlUB7S4G6tFt/cnTNG3ZVgmBI1CeGbWSS
w603Ai2DhlPz5hhiMGCVmwTW/AJ9Ce6WxFqQOb+Dp+rA/nRMMKu5pi2NrzU8DSx9
cCMnUMfsMiA1KYyD2Y1ycgC1pFV2lVQ5WTEfJfPjpAfKesorwAxR1BVOJg5CW7LK
wEzy165lTjXVxjSCQ1eFNVUHpEt1Y7Kd7moY1XzRczoKVKRnjdXXw0ITn98wI/SA
nC9G9yBuvcjf3qDrXnnFBwU6nIFAOJ5urgLQce7qzmvm7MEHgrZduy5dmkt8N0+v
bx7opXYzGl/0pA8YfV4fEd8hm642MhUx3+yx4SaW6KZuq3Yz9PXHj5TSC8T45b6P
9ItX8f0hQFgcIwzhAI5dECvB/8ED9a7JjnE0n0BtLe3Uh5aaB8rilYflFazsTPCi
0LHPUZA2/EnFViWJ2Uh+11ILNEgBhHWvzwkase68yTbCprqarG3OlzFSfxxqjj3d
9UUmHbm1Jn06NBSbm0i/JHlR57CsYLRCsdDTUf2wADjm85V9Hn7WEQGQVGNkKfwQ
SeEpWHxmO5aHkobuiKIOMqOiLKEnwy1aaxz4ZS/I4e7pSn97pGValNHbY2lw+4r6
6b/awOoe2SY0yxd5y0spVWShbl8qJaC3ZVmlgzU98jWVP5GdDfbV/n1uNtUmHomW
AMIFBXqH57x4IiqNeHVwPpvlnGsFUcEWsS7GKNPjnoZteOuHf2s2GvpLinMWIL4E
Iv64hw3nUleOxjiDryTZ2KNdAkaqGFE3i0lDQAP2jXhAucRqV1y1TqcZiadmfLQT
gvLrxSIt4aHYjKd+aJqGlj/O+5tskF3OJ5i3jilsTT0hGvAmzpxVvyEa+mwD5Kd+
cBUfi/JfEYzgBX8zG2egeUjcyIB1Zq9huf2iwmR0l/7fDs7wFhh2OgxveYcQLFdU
isOOWsDI1FzGQ4navaJohSFywKpULUHy/QTxYdSVLkdV9/2JSd5OOjaCq4N/PoQA
7CUSYz/8K3W+e7WjpsK/tZXIWTxfBhn97kpAZwBvss7LV3i/sxu6xfp7Utm0EnHH
z2KOwKG4b+r6tDDor7vqfBo31HkWarP7DBDQ1ItcR3jhgLpC6ERHJol7DPxywukf
/6OMDWjN302j1IGWYG0k7hP6fnUq+HvW/UoIwIaEMZ3TWnflarPyPAQp4769cN/v
uOdWmJhHjgOP3RFPNVz3ccO7Fd/2lwSyxme+sJQv7kce5CMeyxgXfRMr2ka7AwYX
3toGOHOBXVUhfZoFvEKv4T6cqR46CcsMh49nlK4IsOokOFOS/WoAAveU2gkB9Ir4
rKw7vkWP7HktgmU9wUHaxAu/HXDgUJsCdh4yxBrKqqjCjzY2Ybyn16fjTUsKVW8U
Ifsdc2zzZKh2VYcByXMG7jjFseZB9mro+6pnWOJ4PAzOQTsRovJ+t40VNap5zhCc
/YrYI/RIysV3yftLTMRMHlDsJqZnm2mEH61blbFhqRxVGOsQxVBXD9vlrdXoiSbH
3yKxi30z8FdZEQ1ltq6U1jBdfjeiwjA+aQnwEsvaYK7VtSeVq+LKPIak/yjsKrf+
7gkKFWCJ2uekUUbjNG4J0xRwDV8YsJqcFSWfMagzhN16rrjOySRnq0BXL2ydL66S
8Vu3IgMJE0qQ8aDRh2+2RugUwhHe+tzHDUVn9GVigC9KjkzCi6fNqvEtb8vmFPoe
fs2IHlS6Ek2YcH8evqgzg0ivc4lg4i8PzFG3Od7YAWxORK7fFwEFUXlR4f83pZnX
PnJL9eCjTS6h9TGemwQYbakxID5C1dZqeqUDjPUDATp3Ot0E7ck2caBffQDNLzYz
MYQBJBNpN9u+NQEPLQ+UA5UjCbH2k/RU2dAESGs52JTKOXQxIxjwLtPrpbo6m7b8
2XwsghcWMYedB/e4p9wOad5uvxHy9Xghj394AZUHC/ly8cup01DBdoeo8WwSCyhJ
eRxTUUZDMedoR3UEGSnocFq+K28HaU4JDzftvsRnHw0Wl9bAz17EepMEFo8+bh30
1SyBUvMcr8Y/gPpuLlN0RaBpWNPSAS+oruoG+4Sjokds4IV1ua5x/AJYTN7jBx5d
o/aDJ6K1ffimijcalwR+3ZlFuBWyZWNwqSJWpt6Le5J0b0MZ81nbwuiHXeidlboJ
Z+F05mURGtGDMlnmFkAVZNyQvxz12HlxjNNqqwN7Q3yKCrexRjexFl9obQ7FJ7TB
9FG8dUw82+lAUyNP8mPYMv5xovHhZSXKB7DZFdZAiZXJPJAtdEWp22NLa0EjT2zS
NVDeSUwLWZCC3BhlUcPnZvmwwlWVXdaL74MxEElxyjM089UeA5Pq/JDvwXUOlBTe
gwgimLDFQmmWyskH1seLw67rqVQp3bCxbjkMfjJ4gZtD4c31faa3tRe4dijA5Vgi
ZvhItRX7ZhztQlli0Hg9ynLjppPaGMYbV40C7nkurZ3DqehhfR4w2YvX4KYxBpO3
8dctQerM7gMcP9DJ8blLwXOzQm7N7/Cs4S7j7GLsl0k3kQvLWVfEVqkc7XTG9SHT
xk89zmyx/1m8sYsqSULvq6NxD5xX1emUAKe0puGGEjjPftgwkSIFQeGwSKqp9pyi
9buwN8JjrSOw1vHT7V16aBy9gKT3hu0ooxW0wTKVqMT0UF6TYsayauPKk7tu7jg8
zewDG2SqitwyNHqvNNdCafZwAdrkiivxi+TE4+gZoZNGl2ZcQqgG1Hk/kX4Hiz6I
rX62YGi9RbiVn2CTFeSuDgURP4Mz8OdHUBGP268ZtHsFiulBjw9Qj9QHcXUddDjZ
OFw73nEGsFSEHNP2O2sMTy1gU8sXV3vf+Iayj5mqH/kKx5JqqBnQwhjyBpBM/Exw
9Ih2vraBLpCJy4k+5g+wTSdsGdDa9jAmpqcfdN2vRfCHBSKqcPYsMYeeNAI90BD8
KrlBBRFeBwhq3OGWfpTK9wEOQvJYcPbgk2VgmaRhcoCKggZ1hxqrNoj2IA1pRr0Y
g6HieQxZ6hLPKimrS5zdG5H05OtJaTdAYs1QwhQJjm1Vnngn+BcPgltNRh3ErFlP
SnPySrM1t06l5M0rDmQHbEgncRmtd0xdZMskPr2zY/nds4i01Q/WCQ/97JlyO11j
5tle1DWKnWHp2ytafoWYfZh6KXgWjbbGFr+Z0gaWGjouXHFbDxJ7y+K63YPLN97N
V7la11bT0GuwXX4p7nqTngI8uZo6lVsO6GDvUWOC9FV3EmSPXePDONKm0Xa28vJ6
OsjLjTFLLRTCm1n4OPbdbf6tzZVFpFSzlbOYE+1f3WODs5gY1WnKcAeEozY8w9AB
XSqoC+FJkReMmpDkyNFsBW1FziVJ8OEn5rFBcKiDKRkZ6d73VVH4miHymKFxRQm0
1rqJDy4ztFe+tipFrPwCn4/rKK2uT1MLoVhFsZlJtX+Mn07gAqDK+53Wc2GQBISp
xAeYyZgycaU+U5WX9SxtlWW4ktfgAr+VjgbASVxGP/5zzSgyFHaiB0cuEvDb+Sje
/zitQ+xn/Ny+N3lq/SUdJCiAJR+9CW02EtF1EIUOxZcdkpqYh1TeyiZnZrRI+5oe
9sV6yWZS/98RB0zZNJQFOFfCvDPWrsbnmCcYgUnKLPS++DsqCZMuhvbDqJoliY84
YUL6iC5S6LBuAQs0GxUmWn9s2iTBzWyx8nXixKn/ZpkONuZ6hpjg02JW+8fjRSH0
cOKoE7dpY3NxpS7Bid9thyPOsAb8dEeduZ1W/TbsrfdS447kAcdeAkYY0XQlW6qr
W3dBwRpBDy9K4Jxd/3hzWmOevUMKbePPmdkwaGICnk4PWeRbywKyGbg5lMwEj+Zb
9Bha5LPSFI7eDJe0QZp7kAUdAfJQV9Zfsi0JdoACnmiu0uoiFL5aHXqAJ/DVgyMv
v4otbaDZvC7S5y+Y8FsHMWmIqZJ08C2Vtt/gmpTrGtihjMyQMUELohAuFMWEwrjr
L1MQiKewSiShS4W00/XffyQ65jjQDqgYLew321SJf0vu8ItVEiZhHD4zLuiaFegy
ML2pn+NWgpNFj6pO3bI6GXIhJ5LDUoe5juL9nh6t/h8Qqw12rM/VygS2G0EZ5hVV
kkTa5uiGZqgs7sBVrK+VVlXQmbsCRIGm+MhEFbWquhp4lBHlHazU4olIZh8//nwT
Pm6ZS3mQ5haifw3FCzy8Fi7+UXMdN20iF4js+wKvMu4X6Q83Q1NkPRUE8qRrAVai
lM/SEr0Ja5kaYhSnETN/R9NuIfNCtLTaMaAFB3YXlOdi05aqs/iZhOSm96QUHESM
Cg3h94T0nSK1+gTl+yWqsALwt3Hsfz44p4KENFERrNgxFRdQpEv+4BSRD2nVLoiD
vLoMVSnEjJvaprDVTAHCPXZVWFuQYm3ayPc0Az0eDzrdBqP5WCQyi0/zRGaMAXVS
vaRP++/FQmQBYQssZJxgPoPwUD6p6J314B3UcQ8JJ3nPMqWCWLOi//K/PDPejYSV
k39tsYFGmX+Wmvf6c5b3V93Z9xe+ctWfXSdNBI7OFeLSdoIU9+5km6mZ4y7Mtg8o
ru502GLIJR8+ca40kFiHJueUBD7m9+zUhTBIrGaXhdO38JA4AZeAzRHXY8b+FXV+
MvaXKvPXITEmJ8GQK2vz59099Gprdo3LnXoS0RTDmgfwhCScBam3OsOYqdUqhA6v
khlhlvFhKYfENToIpor4LmVWPetgMUuydZD18yo+wYS+gCoVJdFDebZI3NcpdrsG
MBvBSyRIc2ihS2P5w6SN/KIbY2dgabY27/98XoaWvpXW7biumwwNxylbE6hHCloV
rmKgcXGDtE/L5FrFNO8xARS1tq398ZISiDwLPuQNsVuHT/vActgTKlqNpYEldBOL
iis1613yycVe4KZ2V46Ercd+8BNnWS+XsFARLLi3ogcVUPPKAEXFCrrgtz6hn49S
qSlXVbTsPETNoitEXGM4Qt5+yyOuGv8AQMAQrnj3pI13IQaZwE5wlKjpetUMwRA4
Hc+SbDXFcSd8ZT9tm2m8BEyUoCToaKdtmndMPPB4B5ygdvSdpLm0i9q6pTRm2pg8
55KsvyL8zIuQmuCFKvot3ohbeBbD/v1DDa+Tz1ASN5hRugkaYxq54eIHb4EOWJki
v1R3oMUIBY6IEYhGLWee+FSHR0Kh3Ba+9Pjp6GvwL2XEKG5lV+7TZq8waPGK3Mvc
JZwwVBFvysw4cXYy1i+mDQ06T651JuexvO77HOt0QOQXh/2iI8QznyT5P/z/y8d2
YpqKa70RJS+ccRbyuDKFHr0wVOeL6zMP7wRcNsiNRGt8WJRjRc6DLr6ZNF7p1USw
zLBqAhQqRqxBbQ3fJO18fJut3sB9/r75TzgMFkvV5RGeHpJaqwrnZni9fcCOMONk
j+8E7KnVQN+QhU5lLgrdEA/nP/K5DUl6yw1yySzK3qvIi3gsgE8MpkFxvzrzcn8Q
NaSaKnLdKKWk9YjOXl1Oq0AVm72WuLll8P1vah5VkXtWIbA+l0x5fS7HW5RdC4au
q0L6iS1fP71zjhInRWA/Bd/v6r+rpk12E52ySbtrN/TzkZCUBwLnBdjcGtjbQuM2
wuwE3vUDOAt+O4TwlpIrb6TgA5ipxWrmfIZVt6GUhpy6MkuA2eflqUv6QBg3NKu8
v2lA+HXvWr7Q3UNXogK/GGLVp4vtZu6FvarMb+zwOcc7WMX4Drwg6rB+z4MGmeWj
AumH50Xp16heErdD2st+e6p4jwpq/muR+TB8uKcojLhP4a0iWaI04uzicTSNAvr1
sHaMSNHN3iW1oGQ2lOiTLX3XkJRWIBM3Dp0nKud880Uyr7BjBcOn7fTAtLAtzHn8
F0T6kTwD81nDUwCe1f5WbvY1xOq2U4bp33fUOn2+wIVa3MI87xjG9QGrdrVH0N0c
jQqkokJNOR4hQE836qp98dw4Uwad5y1nE8KrQchtG1EZSEDRloYXVIPx5HG7QF2L
MpQJVmOU5xnigEbRzBjSR8+OFQey2ar0a8q7pSJyVPScsw7cnaPGXv2CRD3D8z0a
/DZ9OCS8nD4LmDR9YSU1ZHdX+zdlkx1oyAtiEqXJF9849UlAEX/9ctiNECCuYBu7
jvHOACkPxJLtd9w0JWI3L6Vnsjo0oLD1vZ+u6Frj5P0Mm68/8C5F5QamIGr3pzDI
p+qu3pXr4RZ9hYsSTCC+BbTHeClHVet4GxnR+viBBKp57+9rUNoTL3PyS1IfTZvK
Bg96rwLPyEDDGodGNDebMyX3AXPhsrgUvNY+fV/OqE+Grcj7h/zRd2syPu6hnd0F
pQyudRwp0gO1ckP5DcS9DRTggHzyPeRQBV00ibi4rmaoWQae6NkKn4uxUaDjX1d9
r3chiN20Jt1VTn4RDG/I0tat9iPETK4LtbTnVx7wf3clXQLXy91hFAauBZJDaOA9
sIm/iLtYcQPgciyxly5V36kRl4EPAc+05JX8AR5jfxwt2hyRFdfbBXyZzEgl+4li
WItly0w5Jru2TYEEh/hGYtcVgVh5EcgIvNFWna5eXWYbFj+5+aB0dxgyDs+t68zR
VObxtXFPOeCg7wMKvixpGWNin9dIwBlrGSdoqKde57NMjdXnhvwq++ZhdOHk0b8y
SWEkxyEY/iOwCR1yHQNXs7PpO4W3GuCAttnUR3PxU7Zoa/Y32Ba1J77mHv+y7mdv
gEJoYnt3RCyMAiu7iuuOJaOBpVDDWqD+nQsxUKVw+tESCpz+AsqaPZa8tJLCjDg5
Q5Omh2GXJRC6gJfO7+AYFD9PSH1E1Xl9GtSyR0WcLEl1byzA4lBiTmKQ5Lc6j6D8
Lrqk/ElMFPgzrZHP5FnlgpA38P///i4TSe62vogZBbHKU8aAJVMTgE/13tgYLdNl
rnZx91b+n6gqpZs4CvSkljS6hn5d/yTB4/dMuTApqnlioqJ2/aRzRE6Y8xjDueC0
y8O61AlVDOdug6WFdMld3VwrRPgQqkxme5aACDI0jLaCJgLNZmZ5u8eSzfwJbpEx
uWHhvLVfQJjo+dLkW+NB1uZjd0EU3zQstiJunWOJyimJZdEG8O5ZyYBx0gvY922G
/9w4DMvvrgs5lfaArGiNf/TdBUABCGPa8/uGTIfvUbx0A0SuV4BfthhN7lT4IV2c
HksBtW1/SaKbWJq1i9Q44OPP7rj2lET7i2VBmQ+jkwSoSS+qhXWjuphqIOa1J83t
eP9QoNGmU59PANxTZ/LZ8ZpLeLi7lRj3emJUkWATiVQjQ44FJvCKY6RrCmq1oh7S
QdByzgi3H6/yIbM/05SJyr5yXa6tFk0bnNA3U7h3g90VpO8PTQp1n1eQhPvzzQm9
djNYH30xUwir73b7jej2dRNbC8rbyPDx3d8tT9Fs9glo89mrdJ0J30erEui/sGH6
OfJtWEAQGQOF5C8x+s4mSJi9KT/agp6YhISN0lbyiNHkeF1/iwSEv9h17GsjfAyT
KH8ahiv4Jt4mkqSh22ctyZweCGgaDnsacrXzMD25eXfZHBUJ3V5KkAcZBDRP3ePW
PyKyUfaEZ5oi5NOmgrSBV2N1xQHFvNgMejn6UUtxdydhpZHHR2lyzb2ZpWQlASbP
YJBpBOXXjGL3a5txg4lb2Kb0oRuq0ww6bN/OQKKq/069h/An4NHQFM1J0rclk+X5
CuglYsmn2QGV9EczAPiDcrKkVNW5/upC8yWOc16G7GNuXT0LVoeZWdp45LkkEB+c
2wK2RY7t6kV4j1R/0n31Kx5vCau9wJBimO6etYpsw47xLvym9LDFhUefMEIW4u+M
xau0gxdqD9YxNBwLTtN1/sLSDgynQF6fNAkmijJnJufqZxPkdazBJZOM7/hcqpmI
UNuPOaD3FaIHJ7DgobzdmlM2NJcHdtySHmq6p5ZSD1OVGiD2FRAz24AtoEfdhoDP
HXq1SpyXKtRQs5D9Dou97ea/2qLxGTT6ntnz0RUI+1CyUIEg7xcc+zhlcERKjQBD
ev5J2g+jA3tTpyBwZF5C7ktPKXdWrFhV2e6s9xEJVdbtST71lAwKPIxyttd+FlIZ
BUq3UmoO9aImB5gY2FfstcAIlWkrH2KRUpmx3w9LRenlduD0krTiigbHRbbEkdQW
5xEPggi11tNeUU98+2bt4SOAwC4QqwjLTG2yk20PIUOtSE5TXeecw662/eOBjbDa
18tLYia7BxWkc+C9VK3p9van3lNq7gGax4xX4WeaaJDlBE1FiRGLOUgAAPqU9OP+
IzhYwQPEm/RXZ4v5NzA2QQ9y2DpVeJn0ZMkZpLIJhu+lnmaFcmblNy7JEuXnwCFb
fW6LlyfzZEtP8ahD/W/t9mKyhAsGOE6+YUlUgTOgRCv3/bhP1mlyklM51l7jQtb2
0pVAJIlkzf8DEUgYU5QHnQ62m63HgrcEs4tCx79k3fyOgse0bslHAzPXJwEqbXu7
Kkww+njzYaciWk83dPaRs+ZxYJ7nJNxe5VBpq5fIa+uKfL6iKxY7U+gVOENhkdxW
aj/P1zgGkl/Arkib7SUvg/2aVoueL8VNDdaCFb64Ul3xubZJ7EeWXGwU1X3CxX1D
M92pe3on+0RsN3dUyk8x7vevGBANpLZHZLcGUzsV5YgoUAf/2GgR+yFW7fGEPCWO
7aGZ7MAxmBy3FeYEBlFvy4PMI0SV1kJSQUo3T6qNIu9FC4hxwg2XiDIpyWkbpZZR
cRl1odTiJUDKfZPC2y4Q2etVa8UDGBNQfaDKiP3T5UcyYf/VKJX7NEJ7h+Wzwgto
2m2Kzna54osTlQMFqvPrLBMMjS+LS7gQRnXfs1gSTiBEet9g6OhVatkqG8l3An4M
JnnbRlAF3VnE5MDymrWAGl3fWU9Wm7HpL0B843JL+T+cNRuYVQkLNLgbqAH2sFK2
3oEWQMHc9pmNKFe2kqUwm8zWSb81wyGhCI9UxrYBjR2Cap8W3OISlCj+tVpuJsA9
WcKEq12LfQn1c4USeB5Pb7G1rH+FeW5G0tl1hr3hI1Zft6zDkb+bUYn7xM3uJzLV
3OoFoA221ZJlwdj7+0NMtA7jB7Bq7Assjp4AhzIqvWWZ2cdUU2oV/BD8GJhtQ2KA
xMmXG6yeXalBhCevEXcqOGr7MSAecIO0oAU5qU7aK6EYNHpPG152UT7LDP3uek2T
Rg3k1N5ERI34zCbMhC3IK7lvxvzYTWRd8FfH2zG3xfzyOKVl9o4g4ouHYGQdtW9E
wjq4SBOBOgAJ1pbUY4uW0FQPGZe5+mCN1LmhhQ9M0/SSj8eobhBQ0fM8tgrxPRoS
+IpQ4lUXCmRuWbexBj7jRnZ1q8T3Z3nRJadZg54Vryir3GTc8CSbfqTrim1dRkHo
yz/y7m1IB1+mfvdn0KzzPcI35XKbzT3zTbzCfcUvCFFVM0LjxKpMYJpOlq+mUFui
QR6TCOFGPNW2EdLqDvz2+8ojEoLOkYp8ZuZKjHBbwTtLOpkO/u+TEWVMWiy4X9HB
Vy3kipYe7vBSOsL0AhxyGm3w6ZroztFYq5Yqyj92y3wEU4gkBmeLMedmpsFM3Fnb
ImNAN/tFg8/L/unT5KcY/97mjFXWxXuIMhXJTWitkDVH0A84ujWBhZ60rab5BVFz
MeXgLlM85nyB7lU7wWKn8Qe6iI58tfJ8m+xIUCEdL8ObScbmueHQ34CbsTegcX+W
QwnwYOLCDzDfutuQZpZ11eKYDpt3a9aOut7BanWHRgfLXa7AKbVkrfw276cVjQu9
fIUM+ydRkFJJCPDf/jv43IicrmfoEdNSswxzZUqRjPX+R0bhJO2r0Dgy1NKvv89B
zzmeWs68gYYo2prk9TvQoW+h9CFcFRetecWzNdlS6semey9V32xS5+4GpUE/VjlQ
f5eNKSGMyiugB081Ay7GGzcnDQg+L0bIUHNSHAma78HujRVNQ843ZkeY6mNIPlWV
Ea/iT93iMEGH0opAFXwFDfkarPTOMqBcKVWdmGNT5dqWQ4JEAKhhW+tOF21vG+Sc
7I68VmzlqWpFa6RJToJQeHvkZHiUMX2Ip5LHYTbTIrfusxNgSSr80pg1qZNvQTeo
jnDQzXp+cUvJY/QvZBg0J2X65xMwdS/Nfxx7ZDNhdaf1kHH8e5h9nPZXhxKX7Raz
mHmrR3X7/jiZjxbmpxJsQ1d9rMnpxzlo9zRiyI+DLNyEHbx4OI0QP2LO852xA8S0
oVo/8d7cblCI3ZNageZFxqXntHLNuP1E/18pAdfAm0b8cZ4SH+4Es7TQ0HejFBh+
OYvzckDC8CRyrR6XDbpJOH8sWaVxNi6tsf04LmF8W8BDL6/mzgrNqiu8b1i7JJjf
FVdQ6m1FVZAPKJkQHvjOZsi44LkEQZiZbqZ4xgt5wuB6PHMbF5C3nmkzTPoaM+MT
lZbveBFagQIZwV3FhDpOLXdcDX7FuANP9UJeY43Op7tUuFRsYSnjrJEWuRZ0PBie
xQP7Uvu1wO0LxcJiDC0cQf4sI9acgKpYJ8s1jXyLobWk+A+D82+1OksmKi4TJ+Oi
+7xDFQ28E/mBZnPi0DdkA7kV73lTnb2KiGe5ssmA21WVnhHEHafdfMY6kJQNMDHL
O3FY8kl0j2lIP5gfQu5aJmQv0umsbz/mszCuUswaYQMXrdj0rTOBP4P22l1J1gQH
UzlSUJGmxZhYiGTexRqMwfsu7IreHqu5uJySnE+5DV8OW8QUEZYPUjkufV5XLu7F
rBx5Y+GdSUrKDIv5829olGZnIiPXkgRo82kvrRGmByREZ6hARdJJM42dSouNNHqk
alM7jGzZxUNDuepsZPLVgpXoNf6p2TxAUTJoAvdlO87/pkFzmwAPMx9FxuRFgZAL
gmvxK4D8xAiRbQ63X3Sxx9xGzJIB1ysGDXVXvpjiWGk/kgMYTvCrtayR1SsnnRNU
CAA/fTGcVcYnHWorUMzqplIbGRK0hSTPtJuOlJxrHmDHkhL69b5jumetS7nXTF6D
6WNQj9ILX1unuUahvSMY6qpFdD1cJgZCQRTroM9xAsgdTk3+yaA/1PVzDNuhvz7W
7GSBp54qRklI7CKjqUDBf+x9o+fu3jdsZ3u4xvJnAkIgao3GGuEFcP2XP9y8kRWR
4VFlpPTKAAI8vzRyYJIwiaaYL+lQAS2M/NY4dACtlmLbWxqXw5S0qc/K2K/xxI5T
vbcTF6NXocqvfS5cHBLpqOJOLp2bIm6xxd5dXgAV9Fu4NaBVPkQbvV/SmtqBq8VT
TI7yv212z/A0jJ49y2zn3cNGe7wIUY400JnaADAy0yrT7DEaX//DsgXMmfeQaBpW
DIeKS5buPj2ifmoCAktSL7sYBww0IQtyP4LT8dt1yOz8kxt4MgnmYxu0hLYLLx9X
YyPCyaFiwznsUVZTQbZGKUHWGLFGza7VkwGSrOTkHc4yxs+dvEfkQtZo8J8VLNph
8WfNGMvynrvI0TD6TjDPxkls5M7bk2cMCYxcmFU8ZNV9gO6jIDGVuQwAE65b/2B0
OQzT9I1B8n4NGUOctbVViWbz/UuOiaJhLVA11c/BQvEp35J0ZOnIxWWYYSHvmRiC
UTcCfiLirhqwKftZDKQryd8ZmKWaNe2iaXFtpTDrukQ6RZmAsn5+dKPhATb1xFKR
Lrz4jht1L659qLf2BpV/OsAHbCHLWqj+pgQTJloMjISduE8a7SjHHNaQCljx2+TJ
gOPOKiG0LCWR4s2rHWisHC2UCZ99uyWwoSPbHM7Cm+QdtUV/E3ruym7rBbmdCuuH
UhTQm5t4Zlv9nIaqrKuynpOMfSXAnQe1PqoXDl20vzAza1Sz11gv6SP4uJOBuiyS
1o6pQGi1G8qak46iV1l4fpBS/LEyQjJWjaZo61LIL+kxkVtZczn+QxHXBxRzu26I
DLBGFXf7nPsozqLI9KR5Zp8eXNZea7tIFz6ZYCwyUqsnd+99f6RBmPKPIZ6FeXVa
151ZzJswpHt/Om23kxWu58NukAlxfuVZth0aD4mkaC4ojE1sfaVSFeDmPqoKyGCI
31ji3b12w7xPzDaXJ4m5cxdvwBe59Fuzot+jhGY3nsRjqFtXKmgETEL7ev9xXVCy
zv4G7oFzj7mh2dsC+sV4braovD7N5pih5ME7wdMBbM7QFmNTNOMfvYc4/K71vZNC
88D27jIaUd6rqZM70n6zZ28p392FnCg3lQDJhadCsxCc7n0MhpJNhiEIe56/lS/0
8bOAFXb8Z8wz9pHCcTxKgptjNWpQi4NCOXmx6XrxuqpWGhDEOzUIVTqj1Z67WKcj
tTNNfcy7njpeEomiQHhlUASodLx8X4NJ2jT4ydgjIvBPhhFALnYTNbErJxw7tYbq
gjJkyVZdmODcZCmKzoM7s9wUo+40vy4o3Sjwwk3qi2+fLqCdTSi0xpjmWWc1E7xJ
QlNQVzhAzsGVMrMGO6QHJoIq9DOg99le8v45CIbewzro+t0wdzM9N6jHQzWujX1A
SqD53wxlXJ6XeI6B9guuJJIpZ61xHMsqfhIULG1mvv/fraFnyXHVJw6hI6ddFpTE
BV3ls63apjFptu0uO/ieAkWC0qSYEkofURgWaCTEPLv2RTZK3UHyKuH/2sAzKunI
GkiuBLOHpPfchesiChLsXI2crQ/ldHhdEQTUhcL2Y2YzKCEBz+44ZiU9tSXPpbwl
LofVUJ2y3kkgzFmpr0szAhJFkR86ZoFOCQ8lMRpCjN+Nx52ogviwbLxdPDf5prJJ
+tVAhThVdZeWqfm8MSZJwlQdPJOlIjvGWSZz1OMEgF3fPBBBO50NUozCrZmZb8Ue
/46k0Dv6VavixOoxlwxo3FMBiuO0U70kjcElqTx7HlhfQ0Bymg8IhzdZleshAx3R
4tOiqqjVwfCEBZPrNfr+QKENy+buSaYYd/802SOmk1EZb9hi0QdN4mRMb3s6T0V1
OdINoq0vtq4a2T6AcqQiFXRNxBJCFopbE/F87suDPPBmp7+AQ0LFk4DbFaRdq61F
RYCf1L9tz+PVnPVQRSAkawA4/xUiu6FPcHa3686mOkDM9SxKOGKZyGQQLCeXwOkW
N1MjzHEGhYEKT1qPJosPRpXNXbvUmRLK8uE9AZAsUKX+kkxvUsIVqUpIe+YOXJtL
fqb57osIa8hp+QAi3LgNNGNHXTOh4mmVpI3ZXW61yt6QAiy89UddViUbzz1vU9un
aYmy8Zq/e4/ugkCUfwqrNUY40WqLyBGEFheQRZdSx2eKT7eG0QuwkhiCcYf6Gu1v
P0tTkQBRWYz4Ee9Zdvm6WM2DWKyel1PLsXgW/vFQwoV+6opq8qrhUMLuGfr7GwbE
dluU7CJKF9EkMh5mDX7HqSzizpn7Rb6CDQPYBSpSCkE5kmFtQR6P8tPtJMWOIO2H
1wWYrbmiqgqAv2dPvDkpVjjQ078t6A/MjBU6yeLckUgx7W6Mh+PAMrcZAL3EgYV/
R5MyZ8N4tOAxIPg2B78aSr63ZB/PSgTVogtNGn10g/krREhvtIzSlj35SIbPvmDf
NGyC6EAwUarpNd+NcyNrfR4F5rvPYV+WazBXvI+ENIdCbb/qALTJUJtFYt5s0FbI
Rvafy5CHZeDVk8VzQY7ihnmWgA2E2v7QaNVgg+R5ebM4rK4nr5GI7Jlg8177ePRf
c9BGZ8NhXzCEVRJEJ+qYUpLku7wkc98OVUWXz32z1kZC6YvXL8jwgLDMHUnDohFO
kbv/uFJYUpybNXxsc0I1FxrrK6Yv4g3ZvBNjeJ8+lSFQ9GHnSDUi8tv5ED/u0C8H
5khZcZLG4tDgflDQpkcVWwMHWJJzIO0osi5cz0PnvaQEtG6axdOj4a6D4/NpiLfi
KoiKgT1zAbd5QgJ9vwuhX7oxvo5N2jpsvCzhxpcftLZyPdWzNQ+soQtjZLzfrzEr
3xgoGiN23JZm0uC3OkbDWk5FBaiCXnP8bxWeXGCCxN1iZE5E5tsMw9FKeuFDbshS
WCSucjl+WkU563sdNfnZegx4ZK0wJtVGEwtDGWJghgBbBG9se61u5gU5F1gIPwha
m12aeEHFuoaKZyfEIgb+L8iwV1yMuSwNZyaftyXhCHy5dvFXZ7cqgB69IITUixrD
bJH4TTsUa+rCOYiAFIiqk4LyLSEtK2FUY0cdBWni4s1md9csTzC/rsDuHB3a7fCh
2UlCrsv2j88tJdhTTaKELPRS04Ql925YxlErPgqOU57eJnv1YVhx3D0sv8bhs6ND
r4QqJ+8GxMubQei2b2pBIOpYKYrH5tpA9ylhnpy1Cm+8/Rbswqw+4ApX3JjXT/9o
g5kBrcfaQgguvqlyxnwI5eTnjiTjeq6T+q1qRo7gifwy8nQyIwN5cR9eOlWZMK+K
v9ePDLArHKo8IqQQKYmiY0AynMdbi/PVs/wGObP7amtv1S12wiuSQ/hOLSUkNfHR
frJvbfVYstfHNMxxEFFmXNb+ze7kMfT3SfjxBwnCisLjcnlcjSH+QJMrTld7ar3x
NRFvCT6MXTDcZPBpw76GoetRzAqK+asFIWHdlzq98zHcG92oA6UEhpIBao2OBYHj
jOlAnDqooRx8rG4xrANM5Wssn9/E/zdetGd+wUMEyIw9CNMIU6jnjL2TGks9UxZl
/yL4XEBFY8/Y64WP4EQKzFCDiMwTnGHQrWVNK7kcmUR9XRfYleFSAh2X0HDbdjrz
NiR8H/tbShOyRks/6k5+BZ5bF8IyiirRuH7WnYeP9MFo5/cDEil4vAjI48E0cV4D
60HwWzJTYrK8cfBLQOsXnRDkY29J2KVkXyCvkn+E+KkT4fXHhKYoDD8aOgx5Wxcn
JYUtZUMKbNTCZSri78bmhevrQoP8DA5/XsEpB2VRLNnzTi/QghDpQZ39zNVxGGdb
5zlKSoRe0KJk+B3Z4nAXt0NJbixqwnbHef1YXVrg9KqEBe2TusMN0uooTF7sHDDF
IW37yYd3aLWE8vV6ZWMH/LykzyTbtCwKQivUd/pD91DpQcQtYj5rM3sY2ENongWq
Q9raeMW9JvPXdZw35fZYqkYuvn5wUKsQAwF4v2gAFTYlWokPhH9uclGt75goKkVI
Ip8bR1N5BSSVR/yJAPr/ZMAJuzMgxooG3ggEQ3l6/42f1yw4/1R7acUlA5R2BgY0
NQVDSZRbGQ303TwG30RbURUweVefh1N3rFVGkL9kglyfpK0dy/63bhm5AAkgghXM
INhDuRTFngl/dhf4hyE+0ZlljmQa6WZOg+wUOpsV/5n+2vzQe8VPLh96KpSsUAWz
g9QmEikt7FCBCn0FkJTfYbXXA94i8Tqda3ovrv3m5GzAbOjLIjkZ3f7Iz+/AUsrg
74o2C5ngs5tKUc1xDpQT/xAmrnee3ioxAbVghIHRwsnLZkbr65wZJG2CGn++78+e
DbwKgPvBgCq/FJhC8QnLkWnk19/5xhjfO1Bv3GQC/7R7bh49u/fgvuAZAgyZy/rz
ayYeQGfsRe42lqYPMVuyU0s2R1ncReLPn2+BHXt//EMf5+yahLRzeBn2qW1jDboX
SdvUM3w+KIg9mI1nGNJ4bF4szJOBsgGMZpxddmKOp3gSwq7ccUS7poKWTzXI5eFH
+vgPF/F1NkPTXh1+iaQcVAeWXCELqDxt5qh1JfKLAyPFWPqFSJ/rQOz5Y41N6DGN
+u4x3aV/zG2jky9UGSwDEyxrF7+9O8bwnwUVCBQzpSm8Zdxo4NkyCtbWe6cEAKQ3
B3LNH66rJ+cvJ8sAV4Sa6dWVuGimXmQyiETDcBRuloZXvYQrio5BaVIIeNGbm/Yd
O9jmLOCUE41TrOiTLylg3cR+XaqDNtsjLX+9lBCFqZtgLSHM6U9V19YsmGFbTrs2
GLc5caUDXFci8NAAH3KfIi+MqIXEYbAUf2DzghQMNk66jFBsEuTo2FdMNcw847ZZ
XqOHLEOaY5wdAbfRQ0CTjv3ALH/e+xXUIhP4QRjjhvwjs4Qof9W7Dmrb6L32a5yO
Ve/Zu0YvZkS1vMbTzSgcEn5J9MaAbXl2SPEdsm6YNfOX+rcWfCmEtrrkZz63FBrz
pTOY0KeEvj8/rfC6MtFOTusTkLFuoQtoXJMdfxHXi21gkedgU6Lh45bYku+agGcB
wwj+XFGfi4U9Ui/v3mwRkJ4TluEuokev6PL3OC91VXKU3dKHjTIVUiYq46a+4V3B
pC8ZN8EIHchJyv6rVAjDsgjmxr+3lnCLoFnoLp7wWea1On7vvBr6C4ei4BNTpfvo
H0A4HYVjjCZFdAf1Q2VOM3ONTWlBxIm/yKY9JnHDxFc3JeQoIIaA39v3kC7Y2LuZ
6jQE/h/9NAspfhnoSljfmWn3f01leZ5UoAZVJxpBNNt6qRVY7oD7HHNclIT6GjTZ
1TB8H1JcNhSKMCx6o84xF/rX5uRv/wOPMEG56xJW3DC5KlSBy1gXKxkGo/KWK0/A
lDl1jXnpcO+iH6Fjn0DUXVBkqTkuLKOQWN2wAaJLGmbi2W+fe6ozTjvQLQh9fdPI
1mme2y4TOOYEk2nnCVms6FqOohATchBcgO1b/oF+5+cX47dJPjCFnqJID5LFhh+y
vy83GIGGwo7HyvWmPaj/P6g7Ujqpkcf5lq5h5wzXPkrXRuyjQ+TYvUuxcj1hCJLZ
xDfmjDLMcM3jLnSgNoK+26WhRBG0uD0yPs7V2x3QR8x7usTa0U4ZT+pa8F01HPn3
HSE4+71uRTDbCBowy0N8T/Amkh2YqTilUcSIEZB+nlin/spIvCrf0HV6cVxNH/JP
t2q2cNArYU42kVQKpZtxOorno4c/kGqBXsSj39WEPySNStCp3dD8rbSpApyc8N1i
OXwo/QuHLlKXUEroLlfLIryt4m6aVw2pmiGmabEzfl7hLp/4OK2rE0lVpNR4CdIU
ftOJ9odeLyjHxb7TBKsNK8PAPoBFSuNDyh4utIQgUUdDr/SIKAY9nkH9J2kLchBU
1jSUcPlq/zLRdtRnsoWk7ntPUkHr4oGKsbIKpI812ZkhSFuSCa54tMbywPItlDCN
tYFCUVGYs/n6zOpTExlDjUl4xLjsNlMJgJq9wfrt4MiNndK/7DLWh5jykzmcZf0v
xqVUOd87oaZFd+g+iZvx3jqCltoKaTvhhHkjFAKUfmnd+AWkOMU+dBMQuQEIE1dY
KhSPNGXAcyyJyqs7i+0vJ1Fkb3qYK+buju+1BFjn0ujfkMXD2VztknPLTelDHCtx
bJlGozHZyh/N/x5w8vhU6VOG/cttl7C/yOIpMh1EwOU8Aq6vftHs3JTln6Ad63wS
fHNqou3DLYYfOn9f0JDRgAQiFe0KtGiYvNmrMCJ19m/Iz1rQPD3LoCE8elGIHh3C
pOPjpNqDvYie18qbahacGP3FsiHakrVj7xZ8vHf2Be/eKuQSGOPkZFxqcKgt1dfC
JOuD7sIq2pvLzJGTE5ATjtZZayvdyX+OHO+yUBli29OUdC4jc4JYFcXq661oN9PY
8kNrkXqrO9rmZOf5joarR5kKTWvqOS5N7UL/e8Yz2nfM1H9yX41wvKrLPDCuKHlN
1nf7XP39ZwPCBkHfJ+r+hsyAIBaXQCMPiHwHVloO5e/YGDv+xjOX7Rdn/0YEbaat
ZUFMOEAlPBgKwTmZ9faycHWYsqUspCkunrcLJ+fZA9pcfB11CdX82Itm7YAK600U
bhhwbA2Tm205cZCu+eSb+snIMGRIg4i0FvaLbIKZTFLCIbgQ3+75xo8W7oJ5LadO
7Q8TDdC/Tw27D6z0UVymLCt4y2/zaiHOPxxZaDl+CeEl7sVzAhuiXjjMWx32SH0W
bDIJt5GacaF3UTlwMD+r8Pxp1pqSHOnBY1cpHPBV3bCddXKE69XZaMsg96r+3QeH
6DgtDO5PSB/lLyJIo1wxrK1UmlzlIX+kA6LK/0ZW+4hxLne7bnh+O3yoQ6MDNhzP
L0t1GlAvyoAkXhmnwo4tfYzsAFDe1zU10tHfb3MzYAP1VMP6gzqf3ZIfRb+AGt1N
G9JGIKMPDf+kvkS54RDGhIvtxPmepcFOn3jsT00ECoujQFjoj6+OwxwXmURmSUgV
Bqm+Fj17exi/upUmGhBIYDSU+AK5iVU5KuC1slfVu8YI9ufEJcY93ep1bph8rUeu
D0xHsPFJpsZzrXDT46ivSln1w0mQKe1eDIZWITm2BGvv9K3p6neuUZ9dMLbplhv4
msDUIwbfPZeFiMjkEmwwiE9tuVK7NQtKiU4XkRoFMyJmpdg1dDEMYd/eUqrYxjaE
8QUpmJTbYc7VbhtP5sMimEIcR6N1OIacBV8Qhs9pxXhmYGkQgUwDcQSCWAwI9J3z
V18+gB9A/G/JtUND6zZUAEI+hmCnAgY2uO5tWs5BkO+I8t1yL1oOAANeAjbIhSGE
kba3r6pRr6oDx83xTE/v3eW0YRHUKayeOF3PucO69R69NyS7jSvs9yhsp/vj1LmE
65kQFlzlWeI4LRim2x1qlgWFp0SQHGLn9JT+SpTmGx+Jdg7jyMFYYkA73MSWDK+W
FH36XWFi/vuOo4IByK3N1nWmmNz8jCCdXGc6+xgOZxeD/vW7++gRFUL91cRi3ANs
kjbXohp+A2eQKuNE82N20ynNaXMFym+Vl4vQvZdEYPLjaVkavnTrZs7lJepP4kIu
xOchvStGOSliK+aLi7Dv/+w6gMEqYYw1nKPV4AiRgOrShFoUdW4WRiFyjPuv2wE4
5kErXKYsKxPwfEEqYW/zoMwcuWI4su8TueiNeZTnkl5b5lr1fanf0p8MwUKvIqp2
rbbRp4ht7OUJo05yH81ysUqjtFQt8a47y9W7NmzFjzDUzcZsN3eGonMEB67f9ofY
wr3UB9h+m6Vlp2txlm0kObvOpmxAEDaBGX7eDDkZUZa8LFcJ8KwKW/+LNbCD1Sgs
ipG6RUNwSElq+okMrbX+8IzKDXxUZvsnQOBXb4VS3JjtMCWjHcMS80pSzCE7PxXx
8bsEDZ4mYUD+woV0clzPPJaniMMDdSIB95iARZtj8z/aJnCZ6Rgny1QOy77yyXFu
7qJVYQblnc5JX52BvnhMSSkmy/q/lS8sikB9H/Qz8zxwkChu9vwuU+vSzEgxplp+
anKxN+bqiKtZy3VofqUmz5oAh6XpQBdITX5fbZT94gpst3pIcV4HA8AiylSuyweo
KmQ209U8T4Eo7hyYoJVftMLJ0Al6agPDJ3azCepj+2xlDQhRgv0cirOlpKUJc7iA
DXeZK/icVVqeLhSmB7DrwAcVObrSa8CkC8X5u2IHTxQ/9O6bENJ3AO+RwlH9g/2x
YTNwhmVJRaFTd3N4rRKwqYSaAV8QJ4HX7jz6/5sGpD5+33U26EhK3tcYpDtNbhlP
o136yuK00GOombpunI+J6Sn5w4HYxcJOj2nZg/EIcZVL4ZyOoa7NSJFoAGU0z+rx
KJYjEhn8aMvvgL3luI8X42umqMqWOS09b4xTZI16Cpg69PslfUX0O7zCPy1l0QOr
niQo/ofAROofCJwkz/l8W1hZ2HYzxIgefWaCm2AdmibgAjVZFDlgUtHCVvhsjkQj
eT/gpod4f7Ll8vitCfEkVHJ6mFSjg6tNjueUzTiGqPhMTQAcWrrlUGSKqlA9TzrF
FTwX4942cGrZPYzPRf09W1je3CrHs32DWa0zF4ZcoAATbe9YuhlRbjlgNHiKbFR1
UowAsiQCCk4PhwKpf9yuTk2f8g1+gRsIw3lk1WQdcOOOeH+e01zJS37dBLS9Bvz9
A5iHeE+LZfeQAi5+/zB5cY0+uNSnJ5OqNa91kjnAa28yaU/irOLfwQTJXdAJn9lu
xliEwh7/9hun0JGMw6ZBzTEbBd6z6u0NMlzMEonsi+Up5VZNfRdpyXKI7li1YBTw
upqVk8Dcai3uMRAttl0Gl12U+57s+9WDRzO4PJ7WspxVGkJdXjdjMFm2xTaHjo31
cAcCYt/3phDigjSFpjb24H5BKqD0OE0NcX6NNRCPxYLpz1B55zj4OXRob3PMokFP
4llliKqYRrV0YJFOtEuiUtIk5pOjIavTlJ5iEQr6QB4q+W5LUVvOpGZAdPlMnunV
YN2+gRq+DRsnSEmRFRgC37Kk6FICA259smZwv31suos6WNwacbTCj7H0jPOa+gSC
kaWdk2WJXQ8lnbYZeTJLYeRbNsnc3HDtDJlhVaRK4TKBWrOAGYejm841EO6k11Kq
1DD9yS3Nar+89Z+pfP8lgeCWD37s3c1m8LPbR6N+NCOdd8ibchTYm4jPDC9LRDDd
XtCYBQsWzOsKz0LxfDm7Zc7Es3aZo2oBh7nwcFLRKsRgFj9+3L/JN/TSTVm3VKG5
vsJQPuxE5g+/rv41x22LUiI9Qa881HVZwrfPfCURKbUD08ZNjT8lHAfudE3CzOHV
uAOTFmqgvmoQ3D80BYeJKDPHoFEhBbZFU2itQwL7GEH+P5MQ6iG2huytteHwZRCu
o7oO2zMoXxOD+T1QjCGhaZQVhaaRGMBZVnPvawP4TYHoVML4Tr+V0P61nYPBlGBc
bDuAPgMSCGBiemLFpoHs4qDA38rdPFKAJrh199D/ycMO6ToL0oPXyFzFQr3+Pq2g
pSjAq2oTnR2FWDGL1FLDOARb21KqXNIzeJmeEHXHd/qMZVf8FuN31aumCOQbpTc/
sHJ/GBqnwxSyUY4rcjtRWdm8pFwXdLpdP9OhacDOtyOd2RLpQzisA4aWZ/dBw54D
lHgQgX+RCSAdY1DmeaSszMRog+/utbxsJbllhzFpHKHnIjSa/Z1/w0PKDDS36WjI
5DR3bWP+M78O1/LSsY/HJdTkAFBNGkXyOlJl6RRRcrAwiYlFxGr2clKHeWZkTpho
gFVvxWp4gYq/csIQTb6wHk6X1C8o8wFFVU1nDZDPX1UhW3n4stmNvRGFnxKyRHun
3gE1/zRagghz2GNGhIALWL8e29+PwEWBsSPs+JaBMJDbubWtuIGYf6JXZlF0MSMv
Kc88UaHlqJU3w0ML1AcpIGmU+szqibx+wzbWfinTuAEldG5sQaIEgWei0HladWo+
KLoMyH+QQTHV7fnuH5qcmbxPIxfGWd4OuUzdsWls5ZZyiXOFrm/XpUbS2a78UF6H
dmHjVykDpdne2aQG9cO5PN1eYiqNjgJaVXMDhYkZ9wqAmz0Gui+pZNc/taIwXByQ
SE2icrvq7nfL4mz/Y80hGBapztxZoKD/qnn5oI3ezZRCO03OgVhaku1CqQwjESyF
5M6B62zc1mGmVP0X9etmEEwb0EU4GYxiluupFD84vyMdqjGDgXWMBUOGvUYNgwCb
qWrQOKlYBNRzil1/HY3nwWM5UIw6jmYUv/TgjqAAlXTqhymVhy6H2Lt4cKcpb9QD
Bf8h8LyOh4vEA8VquJj83gM4gup0GcV8YEtqlLAej+xGXgEtqQ7zs6Og6z6XvCPb
ydMKqUkNNZOLOK5gYeO3Z2dnxSQ8HlirBbgKahIGxuIAtov5uyAuzvPX2fihOT0g
kZZI9TRTMWcfAPfAiRgsoF0OrCVHjWL6Ipyp6RDF3/Tt2+ZYxnQW/cdw4R9lsCTs
y2teUVKndp88xFvK3SLT4CG9t84QcQqYqakcKlNjUx1bcE5zGg7Ap8M/i7gJ1MBx
rkILtw58GPH5dgHJ9BOoW267gfe03xWWwvagw+HIuTZjouo1SxrzkhTrfyKVhMnW
AgETIdX/Ml48ooEDwkbXzMrjVOBhkF2bGAGq0YMU+CtqPi2UCGT2PqAy2gKPisz8
1oZGzCN1yNwfXHkcVEL4WZuUZ9UHYQ2lVdzBoCO+xihzqg2c5OpWTQY63Ai2u4yR
g9CK5rJyN59xGyi71eHOlmbbSeIb+9SsJiEnWGTKbRDdXxS3zZiG9qMttjEEqrSI
FqpPZzCy5fP7k3h2P7i1m9+26OCYJ52stv/wxUeM0a0VvpTIfKJt+X/8r4tSD4NH
xQC30hbHMGA4HyfXxTRpVwN8HgUzOC7zk76B+C1lTfK4OIOHidcKO3LELCJtgros
Wyr5qETpRntJbqW5L8BDYD4UWF73anH9UU0c10vvz9HsFupvRZKilwJSEZnRpT9S
Q/R/3iWn08TjQwfnRld9VF/thlUYeYKUhRvG6JKWz/8m/L0ZslIwGh97Advu3tmt
ogvHzRF+6BdlcCxpwW4IU1gZac1BGZWJp79zUtI86ZjtrmJJXbvJMcR8z7fInRSB
+8U+mSRhCL2Sr7vD3bhffSX+A4LGsUpKIt9wWuWdDVds+6geE3Z/UDUqnZiGqWw+
8i6vfvUgLC98Uh77hIcldmuavYZCfg5ih/EArKdP+FfveJNJ+4lMyHd9WkozdmCA
hto2DhQTOMLuLy6KiSk77uo5vffWYbRq+9N1mfUIHxdETmEGrZCY4wpBtVeqjczh
NS6Wac/EM35xNNJW9Py+2pF9WcJzM4PHSAvedKD3Mjus978zXGgQDEAJ7XaxBDKx
rgueV831kNm0b/bNESEJXLcBwhxw2RT+K9NBi1YRuxagUb6LWWcFpLKnYc9qZSwt
um1XSW1vIa5p59DOKlgbcjQTIxA/D/bvQFMsACmk44be3Xfcw/n+gNiUG7cUuXvi
mE0iAaF9S1Esnm4yoDPZnr/3i+yq64Zs24wViTSJW0c1EJJKDXRyQPyg+7pqRASa
+X25qjOPIQXEREWsIJnncDcojsU1XTo/WYS+EzRIcEvCMJDBwwu+30LVoJATgN7H
mUm4MlfFbqjuxagfouiEu3b6XPIIrVh55kPRyzCD8CmqFuqqmOgVtfh225CFqJzz
QUHP5qnWG33umjHrvZiWQ6y/jCtxQF9THYwhAmCYQqL4icRUjLcD+336JdlvoL6S
xb84GKspe0zlmDne5BxMjrbn2xH4cB7Z99XyH/PIzXTryxytL6rbCaHp1psWorjS
9rR+c9kpwdyo8og1Rq7eV1V0SYDwO9vkYAB4hJ6U1ibvpshl9EepHBndlK6zd7Gf
renh6Zxvzn7Wk2lf82yaHx0MyrpxJdv0tW+mshA83m5txeP3VyVWLvXO8Kc6l0EZ
2ZSb3qCpdp0/T/TC25gyV3/p6iGkQTNHCutpHkPJpyjCfnR4cSCtDswkCMZJrXCu
f5XaEIYAE08zZ8cU9Y24dRqwWDvvAacimT46ZOWeCu6uxSs9WhDq9u8p2SH1bdTy
oLQk+EnDu4JFyg9XS9WaNteOJ3/eXrnZWi2XPbTMmDDPVEMcMni4X6iTz7vJZhqv
zM4e3emXbgloN4wfSNtoNnB+p4ZckhuLmZk+mf4pMSFeT5Gu1EAde/U4OXPwDJL2
i5+dQnqTFpgNJEnmvnBGoeqrKcP+DOjITs0hE7+utuTuxUzTsl0mf6hhph99qXkV
QzbF3XhqMNrYHo3N/B5CActoEXdx/k7EN1fttFk1nf0acv0Bps/uHgn7FT2ke+k0
MgLRzuILC8ppJiNJtIj/vZsq8QBDZ+icwP/sYTmomfdCXzFdMGQprz5lPzTEB+fu
cklumvIfxJgUsIgpsdu6YRycWIAV1rCJoWTaD3Cl4f6/qix4V35+LgYCv/lj/t24
Zop62qfDVlIoUNxEK6aT0+RNiSSTWsae1Vx5M3f4GU1WW5DowqyvoGLnNcWGhtsS
rtbgc86CZj/kUb+dALirMU+QQEsmBHyBJD4I8abkyFiu2zsxGbZL5+Kpgpc/TEBO
Sf/2ShWYd1t0EQyMeJQnmv7m/qML3I+HttM/e+xUBiQhLtmOa5ZLQYyV2NeOcohF
owexxdD2kXrcIJgmzKuecXm9htt3L0hlr/J381Z6YiOxmV31m0gswINkGGJjRHEX
Z3hfyMFqY6ScrCbreXVk+Cz4b3nsBXAcHEnPmWgoc8qG9duEWv/PG7VMUeXuptCC
Ttaz/d2aS2bbeQ1vxhS0sUo945j4Cvn07PUR1TPLHB2+/vS33O8kGOfSHUkQegNF
q2IzuKRbpK3rDPtISc2t43VnYU8m0YKyc5ak/2TJAko/kMVcjHYzIEEJQ3yN311G
GIU9LLLSs6vCfWkP1Ls0IcLSK0/xwvAepIfGMyA91+0aMQSfW1wuJpmpMPc/cwKc
j41vfvY21t58vOp50YVlVl6n2oPhb0ozXj310gr+QVY/xbTE/an52WRJI93SDglR
0F7mHBaHQu/paNdU6RM4hwf0TSO/FcjttnjKdYmBhF7uRHxQg8/++2gwwU9wSouR
Bao1WvHFwV6GqnVhkncwcELlzcf9CgRTtw9k8LFmG8foY+MHYjLHQ512JuJisNLP
SKEINVfsMgpCFdp5kb+sF/McsMjHspagpPtdraVPhEi9Yrwl8dVKNXPWQg+qTFTp
Lgk1+lnMjektyIL1PcNEi0AhZlu7KyV1neDQI4TvzEvctkkxbToGta0i/nHvlrhG
4ibiEyykKoED4qbDeykld/jkPfGTqMC/1JQAHPyRx/xgWbMvJFJBrziseZikCfID
cq8YzOocaOjpvsIHGhfEHc/7UGIVUxorXtmLfhfvndbgPAkK6UVFE0jf9ZRV6p8h
EC7WATT7lK4cwz4K3P+i3a0j5Fj9K9va8XMpsAnGqH/kB/cAFXxPZPvNog1/IUVr
670drfW7LzkNhrB8qcGmIQk13NsfBj+ZwFNsZxejfsO2hn17sIHMW+yU4CYNLiEx
Ub56qZqcOADtvhjzxAIOZh1GbjqmLcOpPjX61Bciv8nwUmSsPAqX77oOr5zHiYF0
u4Hp5hmsHdtctOMVeYlXpdHeQoZrHJDe1LZCQQ1A8HOR1ubBPpKee29vCPDlKd02
CeNtqcWGi4gso3bD5xUs55Hg2cg0LDWcwH/RacNz4dPWRFRUNJvgQ+KfMpB2+w4t
2GJo/lXFkSz2i67NAJs5CH2NnIO28cWrvzQx7fpcOjXpatKe6/ytw6gaSgaz2v4M
oSY2/kdRF4wqCEwGUYtDWr9beTdiw6DMgGH8xn178s60lqM4+Qoblm3bSfFWopLb
MfRpFCLMR8Qcnxy+sA9qxdHaNB/0P6WPzn83fSd/CbwWWI0UDCLF7KWby9b5/wyA
bf4F7hYpZtyzAhdaDOOP0CunZCFo7oJuaY84vpVR1L1W4Z9wJ72tUjoQD8CGlfmm
W+RZIr9khxfXy+wK5ae8UGPTSU1eX1mXf6LgfPyWSzfIsLpaFLnCv2SMlPoWfwJQ
+NL7gXR521laAmcstFU+BN0vBV4QqPxGI+brDlTZ3cpyKWREwkXbYAxGY5tt4lag
thuSdc6PeI0Ly7lZkbY9aA7v+fmYzwo7FrGnBWPgja7fwCb2PMHHOdwYDHkLH0A2
wdRLU8Hd8cOTvRjhd2BSzFK+Xu17DrOqPDyvH5rDbtMLR49WXy0rFcwb3NNEOSji
rIOKVu4RyRfG+Ibs9aaTv/ZIMXRRiAhCzUVCZvfiuGNOqIegoWffjglfDoA6ayJ1
JHkBEiiaf+GKttDpyCDiVuyt96GIe71Xyt1tBfOvFzzBklZqkAAa6gPOrZRtMuS2
emnMG5Iagx2OzydJAo90zp05gucT/I0+SlIithR+50WHmvCxpM7mIWvZ5OE/FGJo
0+q2JoiOX14yraw6+/3HFrGaZFU0EPK7I5JIvzRcld2c3M8khn4N80JFN0BdEeE/
dfW6L2im05v/JISbXcxaU81YgnnPXfIjVHMRZrdpQVjercQqAeUKgRwThD9R5sXm
LSAwk9sCUv6HA80pI8qjBI5EoC0NSi/93HgpXKS4IKw83t3T3HEP505GyRYmHZ8F
u6usFxBuXufbJsmTt5CJ7nfynHkFjE4Lg+50W/2VtncWFcR/+Zow3EJjooLzf3TE
hyL88yU/p1ZOIPHbIWnx8FSzikHdjUKsXqaITe8IF5bxgBcQfWVZozix7P41g69N
KhRCSRTJTiFFBSQTEpelxww4lEb2iTBAsPh4mjGCXQkwerv1Itr+hRq0UxSd+mVR
Gblab5s2pelzSo5CjkjFI8JGE4fYx85GjY4g0EDBKKQrOb4kanm55uxoowDWbe2l
vkhqVjofEFp4MQp0cf9K9bZmyjc076Bu+UDvOYGnIs06Xs/ZFq3Tl9u1r29e/zIa
OBSKiPf8toQDYEdB+/VZgvQo8qsW0jJtU4kir/8xkslP7QOCVVWVt23QBfHJU3G2
My6/1rmo1yTpIE0QRJIp5pTFysmqgQ/31c+m20IxnfNJgrhMUipQkNWZyasE2eDC
41VEeFU4j+tXqMrdxXcAm2I/4YpTbe9ZR3vQg7EF75POpu6OAwaFteAO4hMfW2h9
fx2YsptNmP2rQyNLjSvwAOYiAbFfSyLPgoLHbIo2fTnmIrWnu1bjyAkEVmQIWBga
pBkY011Jj5JiTdWlBE1ZjDrZvEvFJa4lbVpc3O68uusnKsVwo+hX7yZJ3NKb3xug
bTK4jR64NqO1JpFo8J1QKpc716JfWnxhX80zux2XNpaHpE7XaCUn5RBBtWwIdfkN
CAGNqA32nwHW6v/L/Zo9eFuDv4YIGWBITvbKFlQHmOnlOPmVV/2g4dWJHG6/Ag2x
7Mzxbushk4RNpbEWfwMO57qIHcj2GVkP9gkmVXU8fPU38HgBC0RS3+bln+kC8u0m
xdQZgTPsaU9msiNsvYAswUWsHTvvMlpD2ceCGOgTBcNN4aAElJPpi9wGMZdeNa/O
bCN5916qqxyCoAxX8iz4ilrjMz6ZDMAkUBqxXWwedw+jMuxqwu2rC79tMsTalbsY
g6479nX54Ep9uxFvL+Y6+uqlNKLuJd3DF87TfZusbOMW4mA4XgHg4HG+hqJrP+Y0
puDz0LCvyqLSo/CuZDr+a/ibjv2jIkR4Y0mncywIArIBZ31TxvDY+tarsd8wBsY5
FhgHsTblK7Jd2VhJyDYOvzeHcuQTk2zYorFkjQk14H1VeqIbUw+EsI+Jg/WZo19A
RgiKHXKZmCKfK7pMiK4xVDZKyr7EuQk1xscZqmJ36c1aPdElfhpaYz3S0xpmNdad
4KFaqZs4eZ0Qw1wh7DPF9vMHExicfVWSazv7nZCpjoSYdkHC1x7PCaEfTTHGUN8q
2tNcW3UP3iL6oTm+RaLs2wcoVNeAjPK2bzVymRJXOFmdAjaThJQy9wEj5yLebNfe
hSC10NvMHsUs7ak3feH4SPHvF4tXRGh/oaM2rvGAEvPjGy754rCRoDRvkKbYkD+h
2KrJf0KHnfKoyEmZLxQqIMDKNPtbRryWPYPCSBPU7hxhB2gFpAxMaT4PyHcx+zxx
kHvm/znJlXa2DL4eDbWLkFM4MlCP4/iu1QTZRN48H2zcRcKwQiq9bntlMHnVXysl
ZfxjQpD0GxFyU80a+1vhnfBaZI2W5fCr2h35pYMohGRH65XnBR1Is4U5BGyKo0lA
x2ilnsWXae08bsXyJun2PasRwtgmMzARYoXgPU5b6JPpDD/ioQFQshwzSKyn6YR2
VCjFvpKfv0LI3UUHUXT6kLMrFaFidrBv+bg9EYu+nK7M+RptKtg3QdwzXM9EeXDO
S/tCWAX5wvezZM5LYJ2cm+y4psEKj22hzNzto7A2/qMKVm20RBSx91eSFTMiMpNc
6mXfGmnY939f5PwZif6c1MvA9Qi+StZYrQMm2HogmRSeHVY2qM1ZPaOJ9Bo3ClLG
yT0yIgU3ATfHzLr2fj6irfqXDwEqAWtg3c0xVTLGnrCiFMcBQZa3k0uyBbBQT4x0
wPSeBc6nCUz8rAnV3Hmb9GryYBbMg/yAy9uDE+wp4Uno533mVmOHlQIlJzL1QVML
kYUsjK4KYvOGUPMDh7vNFodjkPoyKHGVALBfU24A3YZTuBR6Rc+ds7sRWe/V2RcJ
jYO3+Imdwi3cFgabAFESoxgko0iBoED6BozRR35XZaCVEMCSR3ISEU7+Jh+C3GS/
h6sNuUZFzPBSDxoZgYNwc3HK3nzJ4tbkQZKKb2thF1WqV/an5VK0VmyRD3F575RR
byJeo8bzHMbg9Z69ZQmMOOszoAL7Mk/7xJULPNlCy72Z+Ldffg64kcmRyipbDhTR
BlGUZltiEPh+s7hD8JeKBTnQr7MIdyrSUbPQ/TNF/iKIA10+mbpblbbJDQgEPVis
hIoQIGZ/O/Wk7xDbnIodZPRSBcbzkbfWDM+OfVvIWQREhDmCN3X09iMneaACTR1r
nfEoRUBHTTWHbBR+tKUZj6zcdzaAikKP5DnJF7E5R7ArwyyqduVbAL6qVufXaZTE
zvK8rWQUh0EQoQjAtRGC6oflqxwrpINnVAkuv97PmYLFo4coctZbFZwdNwm+x4l1
CL9zoPl6UzeW0TO2SIqUc1sLwMMw+n4C3iDK+U8PnJ8WPwbenPRoO5+MTwu9aUZB
rC72b62o4ZJT5VgldchwobJaEBJUHISaCdIuXe7jBlQqm28scq9KBMO20zlfm+2P
eAS6twgWnaAzIZSCNCoHzQ7GFdTcJMMyikAArYX8qXZ5FWt8idSdEFlAVb8HSs0b
3fDdsXLwtvDX+4fUMu20fTlpshBjNvICCcS588Lr8TD5djO5VZMhuKvn3LFrucmk
ZzA2fn3c+cPXq+JCRmz5vf4fAUVRWSgSJy2ZPWE/k/GXpw75Lzh0lOt5joQWeUuV
j7LwsI8XhbTjNELv/aWOXNp8S5pK4cC/J1YOQNgARL+pIkp2xJ1RVV0qo74Q4Pfs
WjOBSRE1W6ezazZqIfCZvESDur1Wcw6+Fh8T7Cw+Q0EcRZ10zrlfc922sSdHZzcv
bYIwS5wOSUxwdvbDZRtMh+aB59r782Mz2QJEzqtOZuFJGLMrJm/UI7vx89wmNCKB
eEKWriTIlAYafrAnfNq5KGzO5ZRQljbmIaxToi1FC8wD+RlG7ZLQyjjEUlAi1jZw
agqz1yXlLhb+lM5m0+ip9SFuAoQg6d77K+lWWySt/IvlH1+0aCCzesiAdM1uQ9Ca
9NI6QeDmLKWwKZHmsRxyPG+r7Fl6P9blB/BUt6S3VQkwJyr3R4f5Bx1BCax9Yor/
F4xl1C6SyyBjgXj8JUJ4Zompf8MTRMKylfVz1WEzyBR3FJmK7TZhwXEljUBK2Ale
6hOXbOw3U9/+QkA5plgqMeKGnjt2WS1JI5LkDlyVxwA6TSR+QbSerb05rbcbEIUb
l+AhyYl3xQqth6rQwGB7Ue2sGUoI9wzkowQf4YxfPicRlF4p1oso56XxmmQtI9Hc
ZWIHhVxjJedBCu5RgU+OiQkb9s/1gTiVEqeEureuCKzd5IA340jPlF3MchxsfzSF
UxtcAcBujpgUqY5IaFnXxKS6dQ6A1Yqivzb+cBoQRzLbZDIc/K3YeaDYYSn16iFF
JDmHaZniT7bWfa4KxmkMhPhUigKvr/nCykcHmwChOXHWGH/VccU7oP2KJXAltAfj
PArWkg1s/S6twbaTBPJugHKQUDRBgHoAXYwr+3uhzK1wTkYBlLern92rqjkRRCCf
+6b7VaAHJ1gx+VeGV1nV7NxsMFOZ1L3jbrBIg0hF0Ujoup58S1mYpDy87J2A2cMR
zJY2jK+nfPi5FZd/2xXozRkwo8yVEYAaiaSvlR5QOusMAi9l1kblV2iIrz7t4hIT
ZzOBvBCrMNw4ptbVJMg0LgTgN0SQ5BRZmTN63P9Mi0rVkkRXLQF1T6mXwP377Q/R
aY6GWgxXFkkSOKxaLf6cxtOtIlcPn8ihZ/Li7dQW1LNIC7PbL+Rf6wWV4caV8tWb
AgEBqs1sJfZD6VnV3rMKOaO4eOflBM8GogGQ1egabPgDoMaz97b/HX2jASFWVi0a
vZz6xVki1em3P3sby5VvLoGPagquuzZR1toM5gSN8NcN9Ov2x7FSXmYXFQ8vga/D
BT9bBKXNJqh8lPkzstStUmP58yvl2slLawu+ikoP50xOIfkgGIQx240ay576jxUF
u4nTM7mMwpvrHjPsBDxbw0/zrdGkAzbsmXwJMbaYTky3fLFzJ4oweMWnKbOkqktk
SLDVD5RWnrkaOO3IXW+R0ZA5MZ9k+MmyzDiu3P0u6iM212A489jAighMmlS96Slb
pQkMdtl7tyd5v24qv29PPTyxqmIUUc1H1Mlb+22OJVGXO6VyQgS0KqLMjhtDLJjQ
daBykaRm3Kx+kIVGS277UpSHOoRACAz1wRd1pEc5xxBYRPCSSM3Z47tR1L3W662f
cILDvbOIRU4b8wb3dA4yiZUEvmGu1zQbKgvi5RicF29VjRmM5Lne+rHrD6/NEEUf
TZ0akIbfKAMhEvBBUbVUX6RGTeuXi0VEM46noLo4BMR0OxjbBGkfea/3frVa5WM0
NbU8tQrnuIN4UEvLFBWs6YO5Ohl92c7+95XQZ/iIe1dZc2uI0+Ne1MrFtSos3sqS
kQ/3iZPkKGctvsBhrGjnbqofK56/XAY5vfVrmsNENuyark+eI6E6hDuP+ZnbznfO
pNcuGX2gX/PQq35AAmKV41tnOq08g7Xvi9s4/2/nkTU1f0AWrWRXCNNliu7svHm5
FtSK+Cin1v7Nz/1p0Co1maxWYct9aZWogtH3ULFSA/chhBblCkO38aN210YBVrF3
/4xYIcPPY3PNVfXxioAk9sciFC/DxPezJDlHqeqKfcSMZFRd2MwLIMj/Tylvtu4Y
2PqgaGSM4kKMllryb6lyOwN56z8dBWbhIqLmRJlgkJb7ck6orsiWOzUQ/jDKoqNs
8TpLn15ZmMAbb9vk9FWZSKwYfaFGxcqfSH8YttZsu7+LNnhZbTv16CBszLN5dCbQ
DLylwUF6jDU+6Ivb/Qgd0rhriOzJPWfUJaEyRGAxluRiqjUYxwS5o2nNQqD4oEUG
BeP6hpJdVUSO4YoaEn2a996tweEz1zZXKxNQ23z0la9sMOlsbhiVU5nhPtNPbP9v
w/0+NpKN+1+kei5LeU7FKSPGFAoP8iS0mUhcHMjNFp0zNiL99nGxyAfAo+jXF4mR
JRnS8ERysvUvpd35O9o3e1l1LCybAOrA9oaGo+VxpCCgywpGyx50C2a6+01gtM2R
yyURJCyFlZgzO2DV67KWcuqBDBs9i39l5xgiJ529D9Xq2FXgKP3NI3N62itndV6r
83kXUS1/FuCleunfjrTkh3QriTBzy3pJjDaoD/oUmh4rRWpxpITFSDoAcpEjWdse
SIQLY0Yt/8K8PDXjxS2WrHnIes5ifvrYa057Lnggi4KnAgSPerr1TBpzGj/BVzGJ
7uCfYF6zHEdm9SInZUy8OGggxV5xYMAHFcEHB/kk0KJibPy2KcY0ZjvCunuNZCap
/kRVjaqK3kgGfo2Xc2DR1guy+6opiMGsnC9V3jvxVPIvTnoyFqL/GUghywXrCMjn
IZdNbdGv3sPULYRSTZWZGdOlfi8+SoEgnZfh7rGlsYndIGnVjHpYmCg/3FjjlSzr
aP5lvcGUT1hpsu+bcdlghlEJYwK1WfxS484XKzTkqydcrXCgUi8IBGsQV+cqb7id
cPe6QZsFDGyj2PZIpSwRieoEesuMODsWcn9yYM9q/tm9pqzwIWkbGX8XT2k057PK
SAbHONB6CVfye3b/VdnkbM86eWyTC3f/h96edKWGtKEGvNIDAzVgmqB4ClMr8Egs
GiYnfSc+WWHyL+XHhsrqMjc5IdP12dh8ZvzNhNFaCegKXNBMJFd5HHXRj0Rn2o8g
9kBK5IXlGvXP0MCTy/CRfesH4AzwzmruY2X+myHzbJb4ibfjFVGR9EFPK5ixaGlo
rh5BzNExkWslTdVEGnlH1LQ+OM2MnQo6AashaShJW5M5NLSPdNQepwZnZ7Vo0r3H
CniD1esM4spKQGpnMXsRvOJnFkCp8VkRpj9tWUxfkB+F9nLfWz6HZM3519pBINms
Nt2MWHd5zQzO3CAw8ZcG3BElTLrzzM6P6pWwlatnJrw8FIPpf4W2sSx0SbEKar8X
qz8dDSKJ++dq2vwzGAlca3gw39SQW0rqruTDv9rU6jrWoZgvq1OLLFqDWdCwiLm0
GGsmbW+73vHBJXmilDT1B1D7+sh4cfTd4+dYCftoKqLaJtY9KwjGw5h4wnOhN7x3
6TJ/TySfb3jxZnkgeGrc0k9U3kPkzT1FVdDvKZPtY4KFcAY9/67lgjy5tA/dY52f
OphtJoePcJiMwBHdjlacE1IFzSY7stjOMj6bqU7d/3IJfoVVqPhNXlAA+cRE3Xnq
LJUou9DTMM3n0/BluEwN8ht3kRtHQTtTU5kOeTx6kbwXnQTTmS6LlKFVR4RKhd6e
vnW4qGXXYCnnTSSc6+XUFC1z6kLRtrdUrtDnmESM3Bx7rNZim0ZU82sqT4uBdw+R
3NIGkQOI6G4uh/LaXZOON+SZouOOZ47FawARPxfsEL9UWmD61zm9ZdRh+oSpgRos
SHfuv0Ipuji37XcbF3gKN8B5UH2oy79bWKpa64rfZqEeDxiPEToMebhjW+PdFlUc
WtLTP/yatJWX6NJVO71QHP7iT6qfVIcKSSTOFPqfAHl1FGv6P6qeSGmCFc5B5srE
lH6nyVxQRtEwinS6HGhChYPE7xHOZgav4JVgro0r8Eg+xUP1RP9w5iOlLJusShj2
RSZwSPmon0omKIYf73h7JLQDSLbEysaN7tO7yYo/iDNoWaU3wGo1NST5COhv3Q9H
y5q9g9xPxgJqJ5r6s4x5zuNr5BLpkkXTIGfe4UKnJk742/3UD7S0a8gXjwfbqbYU
0/7JmTxOBKbWD7+bkKEyPNlzBVrGBC/Y69Z7iuq7vJM49B2ijghVFaFO0UXnm5FF
hQJdm/ynCT2NM5lH3P7Ra8zmWq2XP7pJyjuKG23MoAUibD651Eqa+dOxniydUgcS
3QOIt0HZyhuxlcTNpRfXrUvDsVQ3rcOAqfqNujz6PnbftiZ1swtw798GDL0Yqljw
mcFJEcT4wl34lPQzKlJ63JB6uQkCxzQdLxafETC77rSkMEH3o203FKUtimfkwyg9
WReR0XOwlF0x3ks8N4o+UHwEI2bc40Jtppj/XZ0ekMC+GJdUrbLrpxUXc5StZVow
jDThq7SXVBAoDSYzqZ/2+P4IbF6JO3QwH+MEunv7igW8fsTOtH1ZC36AGKnN6F/2
4S2QheiVTAycMNeihcg3plbxuI2cdbfrmFBFsT1nh/0/0TVyJscBhOGhlcYqzIys
MKzRZVJPVMk6g782XMwRnPcIcHTI/ZFWyrtMIqS5BWA7D7b+AZmUm/tMFTafKRDF
NLbw0cgDOMQgXA+L0hOG+EpUwhY34b2uLFaYXZIQMBTQZzgu6LtEt5XYlwYy1Q+g
+a32hOaAGarMIKXhTff0ecyUCWGmGthm+/kN/cJGJ8kaYVDojDpemgmlkhQlBq5K
dxMr0DfaF5+B4f0eQqxLsELteGygHCt7eZrmbFQAPrW34jGQGqrAhhrC6Qdkij4M
CH7KPC3AgHiLSQoqEy7HLud+wQHNCLCepH8H9VL3G8rIL94wnrbRa/EMDFwH7siM
5HDasKcWwcZWEowwWhj5mCZgFHVzBAk+xtMGa3H39/HLE70gQF3i9tr2ipbAH9h+
d+BRJJKJKqxIhOEQk9FSSZ0pNp84nTkyvKrseLhHgjHNtfFREzIM++m+GqoUcwFe
t0AxDRbZHV4AFmrgDeQatlM+dGWcXfWCrWC4/Hg8FxiZgfxBEpbj2iFero/cW6QZ
pqvc+bUY0n9/DL/DY++xedhe9EQHRafOY4lsDBFDb1wceMePkmn/WNQwKvXcBIc2
igIZHsUqiD/SDRhH/U5gDmgCeV7F0+FLbbc/jFRJR3UZe7W6HNN6J/GEsAHc95cI
GFU3Nyy5SctVo+CdKShMcZgE21jrxtdXh9BYB6txRnB0VtVjPpuYkmnAn07iFNhU
JR5QO+Ovl19vjY9X07CkQYKjLbhjmDIqYOKHBM4qSukGRgDYOvgB/Wh8h4H/ipDU
pZwUB9hAOWTZe3afyvaxAJL98WkASywIUILr7pVjou4M6HO9y9vVxlJrxzWr/LVm
m77LVl6fJjTXznz73CGxWW9WQxyKYnfIIT2Umcb4WFMGnGlh+ZJCdETv9U4ClD9q
BT60+9+bSmt75ZPyUsfkZ2g93Hov8TIyqnyTcTOpoggAP0uUt4wPQ0GKwD+kgK+C
L2qzkjg48ym/EIompy38B95o0f9Fj2v/yzjiMc14H5/OyCOXLaNSwHzh7g/kN91x
4z3Id6BMiFbHOnKScHk/nOg6Wt0bRlNFjjKTBTBnfwSlzj24lIIFWENzwn64xQCU
0V68Fyyfm/YYMpwGX2kPbPDTUUODSosSHIT3WKl5PuZXx9qQ2GXLArpMPl9F++vp
ZK3/LfccMTkNKzEmGSzwwyR7cogFEBkgd619PIP4vvrZa/oX5OkLeHmHZD8w+R/z
Y8RtHf5e4z05wqdCnQwqyE8YvqZnpHOPbuKMdx7T1yXC89n5dTOOxFb5TDffHUvw
ITgt1xMXx1TFk5v2MkDTPOiZ0rzmyTcLZhimcnVNb2qcFNBn7CtqGpmAjGIbm7cB
V/dkgwRV4tdjXocxnM3lZTLBgfHEURrHE9YjLXcxXgp1FopLcIzmTOOoUm4iJwiN
2tV8MYq3LLzGMZPWhde2jfugyHGbhqHC3js1DXM8rEFF1Jyil5xHIZcodJnGIu9k
WDR80tIVvYzknHSvMKpRym7Ywi7k/r8mb3h8HzBhmEoBXiFJpCike5N8YRJzl7Mu
Wx6/ZnpKKbFZSrELSH2fH+QGTQPHMV3uY0KQ6tZx3q0cLWNtuyBAuXJwtxAwnFTs
vAOMOp2T6edJPznrrqPL6dA8QW29L/G9wNlnNVnCYBrRDH1xjHO/MTUy8QQowY5j
iu4VuQIN0DSw6PTOLXlZArFEgq4/K2fx9+etrFKpgv8fcnl3cwrme3rG4UtKar7O
CE4cS6aR9XF5apTNOOwtwlPU64anjqQ+DEULUFviSVXUNdzVPDXy6bq4mL0r04Gd
5DugcmdVtyMbQUrSaRxFfhra5oKugjm1h2aq8LxDoF4zK6AHEpzkp1IBR9KYZv/7
imScxuz/NPjD5tYbokGOdp+3sHxRS9dsyl2Kkxdo14PG907Hav/4TXhtmAiiGXK3
8gywfp2ABcno7J/qmZ3+eJ9Lspe4tfWbTAFO3ff1RN3ck0fSCZcPZnwL3lxNwlDy
MO3N/m/voMHv8K0mnO8Tnd0uPKIZLIYFjKk3EaQaNCf/fe95TX6UkLc77rkqiHGs
x0PMRFZWTca8I0gkX9ovbjDib/arvinPf/+z1RD+dl/FG2O3EbxmqIzMHLdfDVK2
81VD2dG11F4FzFXVSi+wx0pYMak9R3aiVIk1OsUUPUqpxicKtJIYn9W5B2V6ehcC
BD5HJLlmF9GkZ+6cjxFVLsO38t/SGBWgnHLmf7Z+8xxj7a9moOGbjvefrfWGFkGm
jI9hQDlvvAE6W91k3UTqJQwZTQmCMQPxJ00AHNWY3ou5uEeMARLcFXjupuacOtTq
1aB2H3mVztDcr0aiLh491er+4gZXmXhAFQf2k9WElQtxYnmi27o7IbcxJWADltX+
Vt6tOQSpCyHWVOaE4KYQEvA8/nx/H2Xyi754aLXMOa8gNwny2/oNSUyYEti+br8E
nYFqNf9h84LkemEZI7+PA0QTGdpkk/+sJ8lTq7NdqB9N1a6HbtyCmOpO4EZUIbzO
SslsQojtsRzLmQ2A7+k1h4VnKIOdLrvs48vJnE9fku3taHbB3qNrfTpdgC/6UD9C
XJVSX0xWMMmBDiuFHt6QyaRQMyhSSqEVLka+hNQr9Ej4+oDIK89U0vr3qCO38L3o
kRWCeNwZbVqx/OqeZyPgmJiQCzO8eS6jo7pBRSynPvGoqL82Hsgdm4vruoFyGcUF
ruLbadOKIGEg/FvApxsB8hm+iPfFFgcGjyxZj2Pt/NkgMTc0V4OU49zNRi5VSGAP
Qnlbzf+vuiVIKLTNIUo7uvksDntNLzQzJJ28gZT4T4EzUwbuxbvEZuJ9jzRhUBbL
tNAUV3nrl6ocMi1YqBdo1rlx5eNufE3+FaY9M/XyG91TKKHiBPcx5o3tz2Mpt3MX
vCee9yz1XKLxyu+9kkzDGv/A+ZwDssREIPIlEANE7vzNHfCaZa+0ndEjXCKzUR4K
UsMUy/Q/Vryj4G61+i6YCVu55jZCojStHm/JIjgu2YAlozdgsk4VXIm2EJuYMs2f
rodFFrjFcMaUtF7KBGzMoBhHu8z1Zu+sm02UZ7qvBnkTjimOZ1FWG2R6NzhZv3C3
ftnD3YoLaUPbTWKYMuzP+luKkqs/iUC1ymTpxyCOYN6qsEAOH/p8YbaagtRDzgmM
MJpMWGl/aQ+lJqAMkX3Yjq12GoBw6pv+ecnDWkjm+nj/sSeij0pdDQJNQn65aDyQ
SdF0swzlx0caBJ5VlZ6itRNaSNnyCTqyMI+foTawjg96OFQuO0YYk8RhXjIQnq/G
KSuPsgfz9lzvl7UXszxzTdk+Eblrm5ZVyWDlFJ+xjGfbuP+BK7DSbZ76xBVnf5fs
/sXc0+TK7pm7tx/jU3V3KVmVDVcBNdD79Q9m2nFeeKbAeA1IhaSDf7wva1HeopSW
gqj0iOxo13nbEVNsk2sGCsZrUC7WNj+IvxpC0rPXCGQsQtMBrMVCEaU+PLD6rgYb
D8OD17/C53hxftzT376cFL2mpsPHn3+U30e9IEWVjsKcr7a8PjPIL1zbCgsM1NHB
p4tXu/vWOpLbNzWqCxspru52JuIG4Q/iXn8IQ9EdfK3G8pYmPwurcbwAyz4VfThj
qRdvp2ws6sc6aD5v0HCZ0spMo0yOxHDaPezQlMxQgAWEsgrPkZo/CwDZq7w48vq6
qHZLvOJVICiBDZA+Yn5f1QaNDRmfkeqmjm9o4vHEvp0KLQFLxubZ2T2tDCNXXZeW
k49QrRYadSamyHDdwJNGlLh0EWIT6LzRyBoLVGHeCJAbt+LbFF4UH+qWSIsCh/Gn
TvCLpGYsLLSLSeoyIMK+Vf0wGfGD5gpxP9WzdUoAy1A9NXRVp7CJfs67xdR1d3Rm
6DeQyBSWnrQiDygwgviwWB2CWcu11BTuCqoKkK1L6gkhTbrNEz7w+VyC6i6HOtUu
Ax7hJ3zhwuGYTFMDSVfJBcTikyLXm5BKCrmqrkPbnhFfpcvI1ad5xVCF2374V9Ke
A0RTZr/033svtuThvosGUUt9K28PZLgxWQpvjyuwJM6d9n5StSz+drEv8qpFgTUh
IrBV1cN9Wz7JlCm/z/xos8/vfvgy++REcyRdfE/7g3N5RV4sMylmaOpzry8U9n56
i22ZFfu/PH/bMHcmPAVoHczQHRYbXckBuTcn/kEILqLRkrladpVhDKSxPNOgKFIG
9t1cVkjdCJ57Bzgy0ourbgZjjDaP3AVJ7EPdgrGBGqOOSQVFimj5hk6D5WzryX6U
KgByygJSNVEiHhepMUT3FaG8wT5yBQCP+dkoEjGdierRm2zHZpwe7qa9vsPjVqxQ
rkGe1jdI7zRy5CLHJ4/cWuBm3wNzlatzpIc0Pr1Tnu6NXUhT9kSxhtB0gPeh2oBB
t5LeQsXGOw2q2EtA2WLWSu03knXXCyAdji3suTEp2VRvsyUjC6OBPea0rT26gBns
+p+D9OH1xcfw5aNCbWRk07QYu048eP8pwIkYVndg8OtBMnFX6pdUxxEw/BQ+QW/L
3ZAbntkyU+RZ01RvnEum9Wv2LTmG/jH17tOpuVMm4LbYe6F3sN3XuJK2DLLlI8mD
kJEgIr/tl1P1pd9yYb50UPFQMVfI2pAFG19MVkkg5hKNFxZjoJGYRJZoRuohUQth
bJAbeJuChL6JG2Ybbjv05mSm3iF856ydHt5YiplVMLwDtPaR0UXIFk+vQi4IVp6X
xk+jtzDW3tiSnkROq+V0dJSAOHEtEJoXg+nNTDuVSWtXYnHzt/+/fXkABjLxPJj3
qqzsY5vuhKjmYbDZz/je0raOuhnUdqJGme6D5WHnklcSuAOcOcj2LDcXAw2rgeLo
jpj4vcBx3d4SMsyuf6ht85OYPKPY1Gsq0U0Z/iCYK3wICr/6JxHWUslp8OP/S22j
I5FgKXvmXyuvT47S74pD1vylyjpMp+PG/0hbOQjON1kAc01GWgbZfEr79BbqxJ2k
L7RfSjMFauWzhFEDN96bec6gDFQipIE81MUavtpaRT/xm+WpohyeynTa+gE1OdrP
7moDFZdlc4slP1OmdgNht+7hXkcqm1f4W7EUXq4GrsOng2iKFfIqC3AxScdTR67K
5xgiolDmO0bJ7ISV+MMXX5VHqQUeSgc9GQ08bj6tMIHdf1rd2Fm8JOZnYOuzWIu6
i5DHngExsQtnR4AOw/y9rOnGIHyJbcJt/BZYYiq9g05n52Vj+h65dvTx7s+7v6P2
zOH314F2DXyzgKFXqh+vxwOjb8TFjCo8wK5jI+bnx/6CEfLrCocb4ryBiB5GQOs6
NorK4QFEcwbI02X2tOD2AQsMXkH1SbrziLz2bU17eWXB/c4TSPTbIP0YAXDYSbJG
nvaYWuJI2odYyLsCxqrdZJYd8k0SsX4eXlvFC2LzDO2kJwH7ezSio9V35XgdUKnr
7BK48ntmGqNduFNj9/Tl0nRiVNnCDbSaK5SsVAkfSMy8NhjKZ2ObSjlHfFPomVJd
9ZierjeTF2bBBhZccSZwxWYm+jsXh0+Rg2KtG+XibnwHPOeP3+6t15N5MLWpiZcu
badsBoCQBzh9tJTaPQhIjsqpvDahQNQxaJa0chpg1JqMv2YpGzTyyngAz9f//SGf
X8SaWBVx6rZ/PqDH54mhS/0ITL5SN5/pEiySkrrTcztKoU/InXcSt4EiRas08vb5
HHmxfNymdtneCkLcfvqa1RxF/QO3qk3/wCmQfCWKsEXfAnxelppBMRiOLSucnN72
OF0TL0qSB8ccyfH76hnY2pK2s2iwUH3Tr4vhwqnuI9WN+DGhx3VL3LAIGbAMWxMC
zyzCEYK8QNeh3RWmZCEwUgAHGNnv48NGrd5W4vl9/xkPdS/LdIvpE7jh6ab/x+W6
7WEX5tlx65lkJw/v+9OS3uV/fU5vD8W4kp4MbbUs0ZnSOQ+0Zk113ZYcaae4QhZI
+kojfA1uibdwW30D/L4VpeJjwQS11o1mIkvwKxYHWUXWpqEDWgtKHrrs31yHta3B
uQyHfLS3gta3yGUWxUwzn6f3n1+aTT2f+mKPrXmsr3oYtX58XHzzXDSGHLU/EXtS
4fpDt54fOE8xn6jDydoqBeFnLzz6qoDxfJhX2dZpbArg9rlJRnMBmEBKj/3rBJCt
zaosETxcCO5C6TkOq/KKgRFWdh0LpTLTFdrP5f6GC72N0azTZXVnjcadjbmEJY3m
nMYvG49IP7AyF7dSEu7XW4uWj1nkI6L9djwGHNeeu7YqPnxQQfWoOsZ09j/Qt/At
6WI5G3sAF2b95tReSpLW/8jxp9onW5NEDfhqCGKyRo/UcPADSbX1uOhVOCuyTEPN
qMkS0oeAZ8+AAoWPCf4TlUh7U5cx28rH4Af1Ol0NJawVvcVBgW32os01ZzAtztoQ
lp0AL+VL6xQu4x9EmVI/PmKYxcAe6Hrfh4gdnkXU2xxR3qFaf04ynOzTyxRphYN4
QO/HPTksbEXFUag7f8yBNy3kN5xWtNh38VbRwwb+ZR0Nb4EIVUjoEB9W9M09BeVl
z6IOG2BwvZCaiiYUR5Oajwtd8DNuaM5h+5Tj2Oqq0o7G2oFtQPM5oWh5f7RsMq+j
qviWR97lzO/Dvia9L5tbG1erXFU+JDZTmsNV0Cbg1qFY6yYir3NykQYg7j26sC5L
TiMsD8DOrV/LvuxiTEhRDKzZ2fFRzXV0QhOTazm+/Rrf+UVnRLcwdMANdqrp2Sld
5nXgi1+ZDlicxICXkqNXGrd9A1ri6elr8m2KF3W/1+d6qvZ2V3tL6wQMzP4zt3yl
kGPQpLcFysxidgLCRk/q5EZFEIpoY3y8rbwbQ52lbyS7wqIP09KMynvbNVwE596l
cevkA8cB7VF6xIXa060HKJpk1ffyzj7JsEVhv9Awq6b603X73QTZhovzKYm3iiUX
/rYgyuIJcsoQQTpSzQ/AQ9SHk+8tJArWFNf1Sc3xdxb6Po8rDTRkH93JUbWo51vy
tDNNOqN0HCFpn9bzEdPnIb3jn83BFOiKZ7WKTSXQIScNpljPslg1hXBQV7sAbY17
H5iCnlsnNpkuPBVjsChu7NHQSlYk/8WOdKvbyA02DXwuADJJS4nGj52X5BONaQm5
6ShWH4/Bj3TQ1h9UrbJIGDZhaQzet6YvuT6P8orAuRzwkVO41oRYF2k/P7QX7Izz
egNEVkzePT6htQE9WeSr618nJElvUmbrLssT207JpSEVajKwt/ugRPkIIzGizNQu
vEQXTKkmVdifgr8xgTlmb0GHdOWacror1YHf5uQdxRfDsFCq2oZOZ/1d010VPysd
Vj58dTOHy6arf7zwb+m4j4Td3A2R/k7R/wHk2rx1DvASmbqxdxelAAGXNSF3gjdB
JnRNddngKZMR+yW1cFSyEEM86SIabz1x++3BXNDWprEa/69mRjLe3PHSDPVsIwH4
5yND76RcYzQrX9Xqxc1WZxqc1lpYpmn0xIhSAzTAtYbPj2hwg/JxdRy2SuyxCFZu
e0WdFbV17uJqiJ/reWXa0ZxkICAQIkE98aaTHR+KeA0B9LzkEB0uZrONKjnmMRWx
hBdoXAKUU48qS242jF2gZ/5n8n+8vz0qvLNAhjmNucOZf3B3K0mKLLlNaIkE48R6
VKXW420IYBSlyHg2tEIjTOilW5kUwLwq6fMFqMB6JfGXUSD2vJ8aar8PtZp9jitI
lk4ZeumybgDyowXcWGIrahNyr7B6LpwhKyXml2rCfdq8bGpGY74B+I9+AEKN6zEC
R3/G1yEivivEXfWRI9Sshr2s+eKt2dHoILDilSwHVxhLXtjjaCRb4fssJY71HD/f
znhgd8mjm63VXoDm2zigPtEWXOfij38uayxG7gNEaeyjhDsweSwAiQfe7qk+MNXH
FFxGhGizu4Qz/NLUb5jwmQn9q3gBBBcI9t6c9MhipnTXBgvT04lsB0fnUNZbSqg1
7O6q8DeYmy7lL8WuVZb+tCwWkwAERnsyUVwbBu26WB4oWGCT4mg7XyN9kOlFBYYU
3uyiP1VeaF6rJdEO2umh+fifX4e4+dsYxWtYtUsWDGlNkArpbAE/M4enLsxtnx4E
n8qlhhRLqpVnuCRmFj1l+fP/rCR8+5Gbqm+qRDljEAO118Qa7gSDIxGG5mDsXOJp
oNcQGZjpkVt3iYdtWsobrfwpoWGIiPz0azjOwzSiBGcWay7niD6L6bwFnar7+AID
WlEDIIJl8IH4NNM8QJ+Aoa1kbgJP1fnm3dUwoFfiv9td9Krhd9dHnfKZ3livnNCY
AwW1Dhb46Cp49tAs1MQIG3d9ubBEXmpJpXJ4p/ySx8Zt1xtd6EYKnN2uCQw8OD8g
1kacNivigWS0rp87LwLVJhMRFGb+IC+bZ8tTzeHVSlJ6d8WcUqFvmSonD1pCmugm
UMyCwjvPlSbNNAnLr8GvS77Imjx3PaEG7UQrsAOiEGA7tv3dqp1sWxQKtlcnsQ+U
+bESB4i8c85YTXgkGzKtNhwNls3isOjNrRKI7pP/BOayujZ1/bOdAoShvw1hFgCP
71aqXtlGB3m1RUfdgvGilu3gZ31nuLpoJ/HYnwzIXgc+XI4ddSKH8JqCi7EPMWTs
pj3duaNN1kU04RH3Jw6jVeHZjBrizACmjV42ZOfDItz68xvyHomBO7M/bZ+xDQYZ
Oz8u6+hsWW0J1uHqNmIpHC/6PVkwSb+1pGGLZoesBXb8VSpn5iSGDRnjtZqOFCSk
GeUOaIxL5KHbfQWiN98nl3bwbpmGEhBr8JqJpjEVFJ9I3cB3PwLT2E+utXBSnCrF
QCbHua6uwoCpOXK2TzCYjljv5H6Gkzu7w63VwPH5qswDMzP1zgzVIW2cGxwsYsnn
+vnrCyFrxNFDW0wIao0X0rrvWWzrRS9mOC23fHuJDNtP+x+kuPJ5FGTKd/XMss4j
M8+IbyjO8VR1GdlYasZdENRgIjD4EeHRvUpzZDAjigZYWv7+wTzMsw0jwWmFGZqf
HVS5vV4DtJf59fN72On7YDQaecZmbS7AZ5koyx2/fV+hbD2VZmr4R8pQlcdeQCQP
Eyx/Bb40qlaT2YO/lgF62t64L8rJEksxwtOwYCdwdH6MIMkjhxXp4Ovdna02dlLS
Z+6/XFDKmWiL4bOFAo9G9LMjQnK5mi5YHA8mmv8Xap4T9EZcy76qNUsVG77vNrHk
9j4Gfsp5ugW8AfB0Ubdv5glmdbVBGyidOXisgUSwh4XxuZVRiTN5pGGYmRMIOhZz
T1jInf1wq7v29H/52PDMRQl/AM6JQxZgnHHpPlbCaY3eVvzYSbBDdLEa3vjh7N7o
hTCFscqCaX8Jx9hs1kxhKakE9WBX5nYR950/oo3X5jHIbA1VtGNTGRxU046Iu0fx
BHfVQYoB6u6TjJ11DMav+6FClpULExOlnShJJBXO6Jp48BwO2b4t4oiXy+f3ASes
Uy9vbixye45v7AxkmN6JY/50hYqJDdnfIKWDnj1rwYzXOk0de9Eosr+8AKEBtkNk
whiM8Ak9yEmZjfM0jZ2laQzLrO56n/ktnNKTEokpO5CATWq8GzEQJr25FBWdjuZk
Z3Fhay6bWrbiUM42kTeVeJkXT0iptIsscDXTzkQ4xO7WJaHdNvGysT6dGScfUkdP
G5wvbrl82QAjOgFpvxtSbCdEqeiy2ORBglM5vwS5lED358aaHRVNxlXyH8S+tSiw
Y0mkhiQ4M1waQ5O29J3TORJ+jwBypSfLbZmb6CsbmicESbDLWDogX3G9fVWyALL7
bhHDLTwDrawqbmF+Y0a2ZDiGj7Ix2sWh1rOCdou7BmKd9MsmhIv9pCa+wLsTcKen
fIbpSyBLF6MKOVO0kcOjb2cZiK2dfiYi4CFjpNvHe2HNKUares2wWMmwzH5EG+EP
DIg3TS79tySE8/QAA9rnfl2BGxdab8cMt9C3zj9VoEaZq9D6VCgM6cJ6QcnTeF+5
0FSV8DEpOa8DhVbIaLbB2VGnwy1jqvJe2dNRDc6tQ3BnTJxai+Dizryi/9QBUpgk
8UORb8KPNYh07gttE1H13gEvbnrAVWBwgJs2PKsM2A3YLYYgJp72JfAm+122jgSD
cYup6GiChqpddGOU5dn8oDQXfMqUEl7wWXPl6uA3eslycl6ENrdIUZSZ+V1xK2ym
NRXxh5PYyx1YKvfnYm6PL1zI5pI4AbQunwtgWl3Wkn/jIyukN6tO+yrDSKCivqfd
le1h5EB+S2ajK+gakgm5lBAlfzOa/4MAxnbACeUh7aB8al/+dvsELLGKFFXk29yq
V4+LWh/N5W0tF5aSme0tHrwwVCqh94RwLs+KGwmBx/uiTcxBIuP/kYY+Ow9zV8Fz
zJiuWPGh8PjEEG6cvcHEu0QohzyRu0YfgPEJj8TooUIJe90urfgQp1G9F3Jv71H9
VUH+8b7tb8uNbCEm3V6uKVh9Io4O7CdjZXcIsdcx4UiscQRl+3yIp2WhQKNbdNGu
oLZCjXEsIFDT+ICxSWUhMSB1gK1VZAI9rQOJgrA/IId47C1m4oJRKS5zgP0VI5BO
LXAfzy+G4O4z1FeAxwi52rhnVFuxgVhLeOzdPmRvf6IpPtrYoDjWx6Q5HIIj0k6d
6AELx6Pn3yPyIgL4ojq2Eu+p+Lrj3RTVUeuCQMXGj+3QoC2JESOmU6IMM3gsAEhd
fwSNdfbRT4+Zx8uxturyOVijl8muGJo3x5nPH1UQVLI0i0BSTDz5Sal2mTpgdUPd
DXMFVT1dkQpNWxMXsANLHYjfvXMSGTjnogaGiifhlQTy5S1NV5b0aliJsbx6g4rF
0CUvQ1trztlmHwyaOxMfA8ubxtgxylQVeOX30UGYp/YGF1Gi6hcTPB/q+KKb1YDc
c/yCqn14R03vpNSsWSfw8jOd3DNgu4XcgqhJwep9WJ+n7/tfFpAhynWCJFlsXvJM
WM6WslFZhj8CbEViUu6UMinvXoAS6B+IzFMTAfRMiF/1FYk7jN8zzzL/c6tTgsaQ
ukw6NjPJ+knMM90oQkq/ld9V1XzFZqfrO+48qXgnV5wdIm3/0tmnVpfyhWknR15K
1MLgwW8B7jlNGf1HnV3SaU+a4mybLCvrPUqatNc31Ji210SeS26gexcE2TQx65+l
iEB6/xdyIB8KToe2Fs2IvC/tRSFOWpz7KPAhqWowj3TrYpakxmZKOhQmjLMWGOtC
vVcYp/sb445r1IaYJ4e8+HQPULDhcf7eA/PW02w7pNYsrfWWxp1Na6ZR02jQi0Ua
PsckSgW3X+cFAThB8DyOGFpPosVJcJz8O6Xr+Rt+vWYq9YajBohfY3a+KNYYbpBc
jMPBrVmmxHCXKRhjPjBRZIXw0H6HPXBihM5H0uE96CvHx5KXcmjucgLtjqUTtvqZ
a8aYNRFLDVMNQJSBMPS5+awhrasOkFKuy38UEeQ3km8M4I5nwxqGF5GFWzgXFva1
buglaGTpG/hj1zJXwJ1LVCp3yis6Dho0Lxp5c3XQzAhcnnOlyJULuQrnpPRW4QWC
XrIUpcuKp4Dv20XM4xrZUBouRg7iS+7HYqvxmMvNk8WEF7glQdJ4n9/HOb8pi1SE
uupAkJ+NKpNPLjWeGKs0AwkSdgMk0MUAvTOuUKIO+M3AFYWBjvgS5effINW2DCCW
bqMzPFXS0z7g7fyIoXs9y3fH+5R2M2RGBtOJT2c8HE7d5zG43rVJLuKH4pTfwNyQ
fkQRVjudrNZn8+RQsE/wyzT8MFv4bm+ccjht+e4eNLE+YD4Ap4+T5deYQMVSIvnp
yk3zz2yhPADYeS8XPyVI7IGYujOdnP0mEULamNZHt94lXxeWLS9ZQ+jq6C14OAyB
bE3hndLUI1HlLjvqNvBnH2X34Aw8iXMMButqfn/pK0YiNgvJI1ZZG+bWtx+h7+00
6w+27swc6kICCKMV30rJNkh7JrtiARaSsZ9SA1QEvFw6E9fEsOcSJTUjIi65pEz/
/Pd+Rs6vZIDW9VuBLk8Ri3e/qb0v1uGgzYVNKxsEZ2OMv8Yy/U+rozbETqJsEN7M
m0HiBU/PsUIO//qE52L+4uZ235Dh9dL/t/CDOMCSYdj2ml0oyNeEX9xsiNjvWXHC
8X6rUGXMtUyd9UbEIS5GJo/dMM6XJSMkVdRieAkPoXaAqBH1EPVWvukKM/yzs5pF
xYnXlMKB8najt1IlqrRDyWRRdY3Zmbch4wpdLxGuvaJbRKSwg/x/ez/maV+3Zkxa
Lzt92DZVDStBeDtzK3WJmsjJvS7Hv6mpa6XHC0Gbv2A5j2/Z6alfCcGr6Xr25JGC
MOi1DH2LwAYQbwsdab61/QRBI75J9I9PDqYHZhFoZP8bO2jKFPZYDDTgRfgVgbgH
7U0P9aMSA7KlAq+ae0F+JB8R0sEbO+PKUJk60yFDlu7ukdXQsgJSDrWJKiblxj3n
FyUBrNBGUIUEtl4FT4x33tElYf/Ulur6xwbeBCxqnEq4mzQnzkSI2igdd0xuwVvL
SY0+aMkqYBs47zCre3nYoLWpzEjR2aGWRWitQ8ysXBzki1S6yAnSBsgTKs/EcDPV
uqkoxE2MYs7V9Q9PStRI3q1t+lxYWPwRX8oYNHhNeerQCWFWX9AceFVl6hA7C4W8
hsJ/mlPHI3es4Q74FhoPdeeaBYXJ0yJbUk4mkQ1qDSLNg/AMSjabahqDfCLBNVRp
cic3p3Cxu5MsRP17Tlyy4ev6q57/JnsTVZ8ZGLN9Sqq1atKzzlpdhvpcTeVg2Cw4
9t2pu2Sc8Hyz3qDEZs535Bap5ScPW2efwqJ+SjP4XiEy7Vevm4aGqAhkGfBtMySa
1Fbs/IM58vjmHqzBcrpVB89LMA9I38m0zsd5UJT/fSSxKycObF0Ney49YjjrryOL
wuiqx/AMif9tLDo0/DaqDfyrTEgukzoXZrwAQwdkmhvGU/7Ho4L9XLNGG9o6LoLh
xVMUj1lSDBQ/4c4QOpWpNdpLzvU29ZMPZwak2WlUU9lCQeB40ckVETL65ZP2AuaK
ViYMIrz6+9VtVfEIQ1mN2gvbFk4rgxZVAvtaZo2EQ+BkBzbVf+LkLJZuoRvnlQae
8VD1fe0Y6uJuOx4qhXw4MwrmvprEP2yvWPyNXM8veSMM6q6jVl5/TTyXlAdMET0m
SnsHRDWMyVuWYYJ46tfzr4PRbbikazzl8jGTf+CfokG+HDd7PkQq2xgkO7OyNJnD
0tDVtLtHqobXQ+M+sDYDfe1vl6gE9z3w/Le6TnFnj8qVEjiN9m1cRe/idYLlpqDA
uCm5ds65Iazg/j9lqdIPCZJSuHoa2UteaA0utXcgakJk9ovzZ0XuTGbGEUyt/qWZ
CPWgf0LVkbkVNnnUL63P2g4qbx62mIjfTMrtPmOEOl1GDk5Agdu4CxgB6xAWqEW/
b7lPhU854YQkABXeZYK/OluHWztBAlhrFsxVued620lltS9AEoTTrIxzyycGeKhj
U3c0T+Z5O2GFpI4vIc6XWp5rJuWuGmU5h+WdEeiLrSjH0ZLFmD1t2T24n6VQ3tmh
gAa2MveY58SdpFakxn8l4YoZFc6op1+BYK7Mm+RdZVFANbsxu/fihGYp125L3TDt
Z1HDUwESAXm2Lbt9T+vlVm89p7e3uDwyUOiBGpRq/8n4Z1RgK3tO1xwNXy0qYoJq
zZVOkfIx2SbP1HbXc8Pft/k7knxlc1T0jY5u4mv2qjrrM5CjZSIC0y852aZnuUAg
/4y+MlxQu3C2hPaEN0OhlTMJECfj14T9dUOuA9r8PoRbLSvMEDcev66KI7vgvU2j
2CErdKlOVvoC5ehsN4vYPrg9ort+iEL5R5QnaPy2gvgLFfttqTZk+wAyTo4MZhL6
ZWnxzCbRy5+5fxvWL3pebmEEbIOkMGVZSN4aerNdvZiQn+uvAdgJqhcAOT4rHopE
Mc1Hxij/L1hiArKihZUdjkjxoaO3oCSyWb3wjtqEAtq7xCXlXnGqmcvnBGK2D2wd
mMBfrzD8Dzoo0gOMetTQGDQs51/wGWXEyYkSZV3D/duR9Qlura/ptbEimVvZ9/9l
8f2FwT/MGjcLwWxjwLm1HSr7aB8k4I38+hkoMb7da9rx7ltUxwQXnCQ9CkP6oaCF
JPZ6C5i3s7eXfenn5+FLsif1TJ9HWNBN65OrAL3VJNYd9Cpg+MCthSudlyoAKRjE
O1ky+T7lk3ljixUhNGJ0HPURnOnpAFLN2Zn0pYC755K6yMVRne4/19elWvMRFP71
KlYbLCCD+pPO2vNH4SzI2shmix/xzaXFr9CmzU+cC+1xH9XyTaujVX4ns6yxxmEY
6IAS+BZH6erHLBiLffHaWA6HFQkFIduscmA9M45vqIZKLLAKoaJtZow5v1oOuI/6
2F73Rd373LaNtMQNkzw4OVSAOgwwafe0bw88kOSNL+PQHdqo0Qu3pUZQj8A1iFrm
rzmzarUI/OtBGabKGhwP6m5vFJX5f2tXCx5t9rTHE6CruxUcEJDGoIU/BZmgEC5I
cJ6DnD6Ho5UtxkP6CdIOWgsgfOxDaoGVhPI9yWJZCNN1SSCbo6ZEr3rIfn891+lT
kSr9o0kNV+6Q4k7VdO8+GEHYrMzA379ZWGUCZarxO/uz0IiOyCtcyVwPRIutxs3L
6Maba1eeZPPbZzABRmUPfud7Ta5qrW/Mpk5HPKceu6dofPUvm9dFL9XJYQl7CSN+
njwEJdWGvqv6iAwER8EfY+yFSHmZEmNxCiuRWR/3dFvE1SnYQvzqLeBM+xOFAaIQ
8GMOCt0yIg2OCHa6e0fL1DP4GV6ecxumnXYNAEx6mMx/6FIo8OacqDt7KFZ1WILb
4DOB9sXtjnWOVU1HHEhTBo1e0yY6OicQ99ZJl/MPIg7JBezS6pVZOa5GCV2Jc2GA
rI4NF/tgOwPUVjWs5mC+0QWMONvA9qf6X/KbCDN/+844QiiWpxQWXVgs8V8zH6/U
wIbkivB22JviGN3IiJw8ABDS6efGrYzExR3Vh5Lpkn0d1zhWqI3aYN6o/Jjj9gWf
ZznhEllbovbFPCXWYdbHQVpXmLD8eqeX/LWM/ByyHtr2/nnYENyR+1pPdj3/BPcl
hmHXVxkthRHC6v+2NpmsnKG6A8sI68C7LpAgDWaapM6coayrHoiCT0qiyBgsJ5PL
mmUSKJHxuBKySX+7tPTHlEW/1H5+BCwuYVVbq9quXicX8BmNH7I5731vdw/J1ygr
IG+0iv0YwOWFsV343TJu//Feyrtu13q4MDtM5jY0eKeqJTXU24iIOlJLKNETvM6q
rsfN9ZB8MN/T9+DJIZ+jctgSqFUXQWJ2Iyjnm+LZD1BmtImiibiUj5sWTyEdRs/b
GdwBe4Carp2WmZdwXH99/H0CmdXZBXGMndj0sRnEHupr6g5kyi9qAtZqY15EhjHb
uzcUXltNFCxW+pGOF+MgcKrgwf3byGAgJMNUrmRkQLp82M2uYXEZ0nAnCplnaGi3
jvOQfeHOxJZ+l7ZJZNJY1deoyOcv4aU5aoii3fLkcSyZYRPCA70iAEuT/1v2/6oR
Y7SSHSQke7uFKWxDVxA2iAye0mY/JX8KQ2NlgNu1viAksQMjdz47NzlCk59+hjwU
yuPUuuextwn39/3uO/H0+uNpjkDj2XzSepzQ1JgoaH4YpqNTlaOXzBwiturUky+V
F0F9/Sk7ZX+QmGUE56AeYFYC/vvmGexi5l9HwH3WEhd8/JxzZh9Ju/sjhlNDzF1i
XlfXVMp3ztg8qNP4uTb0ZS6lUHJ8mLCN8T8d+GuIK1uNJS14GqvWIUwDKoh8yr+t
oEx418npZT+BmLNPtm1NxdmJUWV7J+4ufZNQJVF/BKJL+frTPrtJ/7FrgDWuGIiq
HitzA5Hjdqqt6MuiRahYzt+4YiQYSm4Mi0MNKt3qPPBw31xDW1HTpWiEGIb1ZKat
SHr8gfzJy13LORZoAEO1DrFuP6qLJqrwnn38Kv7jAJ0QyDeCFCS5FfJH/iVYla5t
XEaOx808KY/38ecB1M9WaQY7XKrfFJgEKW6jEjpv3Nxz679Ad1OGoiQdS1PirAKC
QlsPACwUPUiM4oWSlMx+mfgQoEeIsU1JT27KcxEPB7WaYRjykxAu3hQytmAfdfAd
W8Jg8cFgIL2sxwMytHvt3B/XS+3/QLj96qSaHBAAUHSDDwZ4/WrFBRijbVsLIkeW
X22tqzGTdZaLdWOOcnnYefCcTiamPA69p7fB/fo44XiIAaR48BRoUKhcbap72P/Q
19qbSmMddwBS3jF6sZwT2VFmwEUJexTJzPj02pwu8COyR64I8OiAcs6FcYgSrCqq
s436kJCigvHLJFsNEV1toSPlNQr45hoeXwVwPy+rdP4rI9w22EM9WzzpraxWo/sL
fHKxgo5Gtt7GVNrXxyu3VFyCbjBp5wdqugVV0KdsvQm3Cf/Imd+i4UGxig/i/O3s
tATRDzrYR7amCM4qEcesnL4SMARdO7eqe8NvqfzpMeJjHNqwE9LANz8QX6W7asqg
xOZhKzkowQdwDXWfDBpVzcCi9UajaBrlLa5rO9TgccPBqLMwcTF3ta8eyMtMQ0I3
ngoMrb+XpE2znYO+eUcteykQu7GvaWi0p7JnEOEwn9PmEnCzkPNdYNZhGIIVetOK
7tNfdLBeiW4GHincSixNGIvYnAP0gHgdS3osHuPYS61ktZa1uLHqa7ESgKg2QwAG
umdk28q5V0n6WD7lpohsdSYLbWkkX4tV3KKpC5GKeyh+DHR5ki3XVfnHQxlBjcyc
zZUTcHdHzE2SkCLtucj+0KHqb8Ln0kxOydmhd7TPVpbxcGyqanSqFWR4kR5Kj/IK
CHZqQSr8zl8MWW8Sjomb9crMoD0f/VQCbEJg1AIGroemeoQI/i/JzL3BSuais3q9
DxRL0CeGa7sIQAnC7Wu4NMJGauuv/2SvTTEtIWbe4pHhsUETIOT+OeM75cIo1Or0
kQQiDUjnfpldjKO5/XODZp7vI9uXkCTp9N8Q3KMGAnDlIN1BFaOvzy4vfhZYt79k
1utpNKL6eHzChC4RS/MNvjQhWD9jA5ABl+cIUH/PPbMrevuxeeMidbHTpANo73po
+7iu6+7gdB7exEI0i43FKIH/2pBsiUGAcf8VoAOt5rfR9pCKfLFl8sidWYAEki5M
kI+Ev+2QrZDrIemkLnrTvcCcnMrEn9Ckk7t0PU7lWiJmb7xbN0GcnOYn8zQC8FS2
voifKiZa55jhZH70YCXBaJVfHeotZWWx3X41GuiA7vSrN6ItX3xHPl9XbtncD4qE
cZIX0yP2WtO2qoitUjCTZe4p40QcA/9S7T+tCUE3avxM+f7osDsNV6FpxzzQMeXP
Vc/YUCyps5TBOgVTQ/rPwICEyCtujLbTp+YsnpbouphDjQxxPV/xfL8eumE7/5fV
8nellzmZX43Rg9x1APf9ocqpHBS+FHgCPTjp8VXbKxqndy/lH9OQIO6vc7ERpEId
uLaebLmID1zZr5yIHPq6hS8dJXDTwpoXb513/MyMSiUXYZ1QjzO7D3E4ow0EZOGu
aj/GE/i5JS80MTMCV98BdSdkR2pXuTKrr9sgJpJAyDWiCO1gD6eZwHa6XSlF+LUw
uUQQ21ouA3y/p3dmEw/MtaaYaHhM1q24rLa4EdnqZMqTB6pTxamiR2LOtX4O8CRd
uQUwg6axLQ/nI6uLtqOVyE1Gh136N3Kl7cHD78rOW4YVcT8FRNmJLYlG8YeODaY7
DgDRWou4oqZDhhYafwiTt5+dvRHLfF9gqujdk5elei8Lbxh6KWehsMcg3J1q1neK
Z8muVDxZyPiKgqObtxXIunq+VJtdT2juv0MKW38YIjMdGHerJulUS65bUbPCqOEO
LFMz4ycyHTjgOr5KB3JysKPR9/64rLynEJwvQ61HaHNk5U74/TnLMcabYGvTCWj0
zApoJsP3zdl8ZmzCav89FQE9rdu1t+uXq98b0PHZz1Se1YOYV0NbOpzUrOYLWhjM
U//LZ38YspAtnqwnti/FlEOi/g+w1IZhXFj6tCgIDDtAtw73xul44CfaTaXra/Rp
oXeFHr5f27Td/xUVhQ/OanUpz3JxQQjpCRIeL6NfZ1wkH1xiHu9QDDleckCkce2m
IMziTrH0B9l75LuapYguZA9NhD9im6lLHhoMFFScIMtkBijueFMCM5D9TYryU5HA
GPg30d6QTJN0Pe93fqYMMu09TwD1s3h95YfV0RoZhA6BAmGk63lO6Jbs3b7NIjts
+sn8y/LfBGlA1z2Dt1Una0rCp8lgFZ01vOu4A4SPnW5p23eXKF0ZH3CHuPhoKc/5
Vn5OGXvkYERV0MaSkq09MEcXJmUoQzr4CsXGbU8/PyebGBKU0ffpUx22x/PbibJY
W/yOaOJ/FA7D+EL1FsSElWfkeRuwSIvYLFfBoI8oxOTJYkcwB56pLU6kolJKI+4g
RFu1geQVwxyq1i95XuaQkP0+Sb0GJb0f1k1xvqMslSdPHJzdfIjbYIpgU+n2HrqH
f3/qOoiOXPT0Nww7nGyynx8UqqvT7NgvlTQgcjf+g+qN2/7ipEoTDSKnl/NcGlPo
79DHFL9HbigR/WLuyzzjRm35DKPj8QzT5ABczDnf0nUP/eWbFg2g0LDAGBaJ6/5p
gLV1K4aCY+MaQFZGyumDxSWC85yhTUwKbF4WiMNefixmWqy8d0fBYFIL7E1RSdB0
CDgEH1rk7owI5ZRHuq9arJ/C5u7nGzkviz40i9vXI/iTXIId2TGn6lXWXo96CK4O
1aLbYkXZJEibQJtFWsWryaIhunKBjjPR9S2BmpFGBBZqU9IoNIP96NMA9brBzIgb
/k3vavHjLvXFuDEyv6yX9qVvjBNmP8KQceasKeMJtGKaat4gGZgyrdrY/DkCtlke
8i9lRqK4kXx/w9Fyu9CnQGGH52bMKkFAcZdBED4kQwSOIos236FzWl/J9CkPJ5SJ
nmOnXf+5bqiajju9q+q29HtO0zBIUHtc0OgabyYSVCWRG1JBMg2P7Kg+JJ2jiKzR
OUHMHv4C7ni/LV3mEuMwtKCAZZRy+HvY7Ou9vWw3BPomf3YopPMz9xN+NGDjEGzb
e1kR2yN5304539HQFCOSRWAbDkKv7kRg8feDtR8Hdg8+bjxdFR6ZTKv9wbAmkugv
kBaY1jDRZAOrr/i0U3mXAwW+cmSx+Ng33xg7G8QndlUk6xQDBPX6pfyELbxPjnUz
4ctAxBAqUD/COSUOQu6RlyXYr834v8ocnkyqIOYjB2uH3797VxzyQeWW0I5AiuOa
4YbcfW0pc2yH6LdL2iNu+TQOtEAs0QWgpY835w4wkB0Pdq8qcBDb1rcvltlBc9iQ
iYYFlme7bVf77sYoJmq/ACYDdft8cftW5Et2EHVfjTk4iBmWrUQLL1vgSkTXT3Q1
nNILh84teSn92MATnLrBcTacCWfJBQjNhPSEOnbemMzHWZlXDIRlExu+m2Ain+mo
K2ZrfBtYgPh+J6ZxkbeoGleJSjGsdTL42ycJ3uNFUTv4rANONvrwxcy5RFx4o7Cz
C0UR778+r/mCwnoM5iiEkk/xtffbGCp746uVMaGht2B0hLBzkScF4rc74clcmuyT
vULTf4E4ruXIY+vAGAwMI3Zo2JkDTc+Iw3w0/p2N8RcSudK3qjg7hGCakFJfvJ91
4Uyl8bxea6hLyFKkMc/71kfS2YfvzK8p+Lf8UdWIAKihNMck5FrSML5eCxm1X2Wz
+uQT19v+4EGwr4+qQpl9vToGJqZWv4Z4cJMW5N5xSm4VtJsUHD1S/K5mlnKjb7gR
iowWgpphTHmL7IQ3Qt5A6mHNU8bQsO/XrIF4mvrvazR71t3Tjhd1by04ChK25Lhl
GpYkR99iEcFvWMzhnu84Ql7F/8kswK9OhTfBc7EdkiQ7lv8XmnpoR6Z1N5lo7gT7
izx75Yhiy3GArzLBwGE+Oqcdbvntqohq32iesLwV1SKXEae7JmEYZI9TdxSDV7ou
CkH35AVDAyNiEjOFwXJJ/dFEMTz6zYFrmlyR77rZq/ifMnjXOBGegTRrFMEkovoR
/okms5MxnEsL2u/xlekrAPKMTZqVr1KX6skXMc6Rb0yeszWEd/HY6IBmXDnVQcLU
K0WGGj/bPyC+y34WKn0jcDo3EXkeT05NSTufpX00R5ZZ2kfxwId0SGh39zbMSqtR
s7+KKu0OREq0Qc+waTnl5XlmEXtF/GXmhEQ3N13D+UDaZhuowZHnQsgEUQ/iUi20
+JmOA5HbIkowDH9UOBne2bSoHvwRHAA736Lf5RY/6k7r/PMlZc8fMo4NJG53hmV5
C1/BUUsl6FQD98JtGaYRIFDe4xg2d7RFy4PNrJa7WzohWw9KUO4BGFoevqf/e1+T
3fYmtNBIfRi1rEioMjSAiTw4M1YnHebggSFOdPiBPHsz2GdcSCQFaFGdZnL37wdB
66nrsFdav3SzcNnJ9ebYYqYbKwGSX2C1x+/smG1l8iFjWhWqpouNwVEusutpum+x
5O4XSNe9m6ADIqX1/qudMiCW+S8PUSD3CYWIoKMlWPT4Xxr6iPiifFZGG/aqAdNZ
3m6e2g0b8krKc1D8XreDDXMGNY2qJZSbL40LgLGQhkHotywDuMlgXN7w3oNQRh3n
mkcedzDir3hNysh7PI6BywQjIxp8T9s4+n03Ov/i+wi6ht/Tr8AYoJMQf7fhTi7Y
xcKDOaYvHY5DmfLioaNsHN0sYhvnqRrWgF8+y66ltchXD+csiX839VD2RIqzRNSo
u5MTkaKgKYN2i/SO4X138ZDn5lF5S5KaULf8a/PwVpqSz2MLfUQypdeMVXKkX08Y
J6mzZx+ldYvtBXlaQEsexszIXXZkRffA1CIeeD+NevRrkgFeWNDNa0H0GUe+KwYl
1t63ZuJK+YNzug7E89SsfhKTYO0lFq4BxhKVZZDZurbwjey3NDLcZRX/CdfRvPM+
7eMHDzTYvKe3q0SycxFpifztv7JGg+La26ny+yocSpDgAFIFBroDg63vu8k+M0cW
Q4twDE/krLgEGyqCwlPfl/d0g1maWUWiD8uBOM8CD+rivDat3hN5JkANpj+bRocI
LhXi27fnrFLCLnZiZIYL1J87kscuUUyOQvnK04xZHaZ53+zE8iqSsQzCLxZRXxed
FiKN8Ae5bfc7NrX5gzyca1a0AmZYWAGkF0adIzonAi3r9BVI4HsS6hkGVMdm5O0X
H1+ztyHgW0LYaMDOPPGfh2XkZZJbwWnkhgEdF169B0DuZalNMgLJgEP+B4uE4IH/
810tyepyzQG2c/rl+VvCiNB2K1fFM0nAok821+iuC5n/5cSS3cW6DWx0rQt0nxA5
dVXK5oSZZ3bmo8wZOPAbZSMpf1RoLEjdGkmuru64XKouc6ZlLgXpPVXmNWN3Z8C/
hdjyTya7pELlle17BnSsbYVsTBxupPOejWB8iKqiUwZtYaeJtnO9hsrhVUgO5eN+
AWIV5EsOqI3QrXERYFAC+lShxTbPaFOvX6RvFfw+5j+UBofcSyXxoMb37cTZS4QQ
HPDWTq1qaoNTjGQCpri7QKkEsugHhgSo8bIJpX7GP+nSrfrFoP+DMnjTls63uuEt
qt1osfnl+BTNQyZAxI7kvonclMgSGTJZ2UHNyNLkrUlTllz2fvsoolR+t8Um0Phu
RIo3Mz1OJ90iFfbZJugP2uPQXnrkM9mnYThyC3GkqIpwxUnpqXXG6rkrECw/ksmb
5YZoxvjOq8+nSvunU1/Dgr9rGwZ52N17IyMgWiutI+xMSn9xsY09IZKrPTEHC+DI
+ak4mEdnwE3AVDeEVqdQBFHIZ1QtndHX/6OyKuAM0SjHSJLdKAd9kPujBpAogzzV
CUzNuZn6v4ixBUAxzjIU0AXSl7Z6xiXoT2wZ1xhFPqIyhfR1mufDLupZR97p9j6C
AmiLrPavVzAU7QrKRq++9lfeUB4JtGee0E4MTIjwz/rqqozAHq6kiuG+H0mR7yk/
MGGm4H8ilAn2a13xkbINK6ceqt7PXmG7Q3c+Ewp4zB+k/LoGWm6NFED6UdLYaZjG
UpEaapZsAS7mu4YXF73Z98I3UaM4DZ6qciF2ZCgvaq4PweXfV6kljm4/yCXQHZcX
QBq7Pcv6cGSzQZhQsbSKR1zFAeIywTvbztsQSdIzDEuJVABwNcbfLSLOoqp6vwEA
vXeCkoca9GTUYxu0NJv5E8RvIB3NXTpHq8/wzjEm290AIdUv1vL7Sla0NdfqSXMf
SY9eWdXPKgzys3kdZE8zxhvmc6C0HquOPUi5qjPHIYDIUWN4aPW84c+25r7eX0q1
+yUnMf2c9AXUm1bR1X1jVU2U3BnJCOaG53ZUWmJIv1BOw1s4RiAPaq/vdz3Ucjd7
0KxHEUuM+TKTaKHxlRsdLtd5xAnc2uDADr2IY2G63VvIlvLWw9hP4npkRZ9SHsjf
mumJsks8XvJ9VyMp6prgAoD5lcZgb6FM+PH3OTmMe1sqx3bP43BFBokXsN8Yvd25
iyB06oufUE0Al1ocUDxIex7q6hDl8HutP61QiL3RgQNBUEu6iEAWGVBDdxlE8zY1
kEO3V/PjSrXeaqlw0cRJDVP6WbjUMF60zKjmM3tCLgEBI8ZhQKJ/E6hOi27uOa7Y
8k7M2JXkAAGaf0SHXptT60K0iYknnosBe2bwiZBtjq5Y9qJdaz09lhBB08XiO3Td
6rcLHatYN5fvSXGUAl1VgdiHj963q/kVzNK/XVIDGmUTJukFA+koHXzUkE1VuAUj
CFL4/KLxt3WkHwx0VU840tYc428arjx6DD1U+F6C8Aam4HBEgdZLJVB97reHTCvw
B37Eu4cQpknDO50VrRrr9t0flR8HKep2WPpkptmz5hNN9vqSZfO4yKwg61yfutYy
IweQPpHN81R3bL0Qz71eLU86eXkVKIAjq4m/yj4O8mVUnHoByoYk08/dc/gis3CD
ApOUT2JLmZVdgsK7aNFUzuDW9bD3u9gbJH8jujEx7bgngwjvRR9cAQ75+RUPSYgr
AIWy2aidVvl5s/cKTqPMxpfSCcinH/gkBJHIO0X7G0Bun1NLB3ffkKN84b9k2ULu
2cY5iBK3vE2i68nr3c+sdt2UbzcLtG/A6PMff+vOhHw8mQh/tBWdYDmGKQUAUKQW
cx+18phuoC8sBK0WLC2/V1pRZ/7HYA6483zy2QU/ulh0sOJZIHGTWZ2ePDMb3Rry
iGrxc49iM+7SAKt4tyGaSM9hu90xbq0Oyp8wy8m1Q9gI+rKb1SFo5HEcY1Q2hYRQ
EyOHmkNzyo939UByQg1Ti2Jb06XPjLrBgAwj7kcWKkYfnJPv+HktbUW8SsN59Lll
XB3BxbWfAod8Y1MT37PWsHjeH8K0gEmFyFmKrnUO3phz36ngwB97D5PZPAkKd/Od
JeFycQ52w27nBEnI7u0o53u9PY9E2XJRQBMij7lTrOuC13tT66WUU9dO5qhh2B9w
0Btae0Ia9LMMmVaviYy+1JgyP7fD8e2tW4jidu7HzIalbtxpgUKPkmOiXtxkThlu
R7zPXgYc7s+0xiZeluS9EYnOkHzOfHUC+JOyRDEih3y2pU4Waaw5qnuA0vOB+Fbx
Me91w1htWEaTOgeATvIlmzwWvojeUyljba1lGmFv5ypA2a/bej0CbsRUnFz/nl4V
ca/Y6c7jwV3O9zTEIpYLnlMmZ++Xf1ZxRv1Nxvy0GLtQ6zrTHsbXvpNGPl6T2WOT
j7/jPmu6HDpqFJvjOxvyDUSQw9//hPwCVBpbl9VLaIY4Zxxx2QBuHmzLsLmCP0Gj
aT7HjjJoHyhCQ0kNi5bqMX8EHdD1K2j1UgqfD8qWBD34UD6DLo/MU+Pmy5JVR+V0
3ZyWO/mxRJ7cjeOLp8Vr3lv6BFM5v3rd0auqxC7mCiU+crmOnB7zJVsx0AZDkN/w
vYgv6qyftT6MNPi+zzCq6JwOl7mTQKnWLEom3rBCWI6UF5e7dsL1dPCI6rzn4B+T
UyKrhXAvuc8tZZUjsGPvKg5PH4Nsvx1RCRNDP9XrhWxC0YPGT365mV7/RaC6yxNn
1Gnad5+nJ/fT2nkrY05kc/mQ0BFqaSrISRQG99MPazNhRMBfN5ZJmDnzc+efT9f6
aRHrQn4mCCIULnvm0Ha736BrJSpUluNHq6/0ien2HPKUX3hrDziACBq1z3emhgRj
R2Tl/NJ0yiuvjHZ+NNAfML/tpGaSRRFW93ajpJFKUn07yN4iabQgk00Iw04YD3cQ
tA23nBnbNqP8hdMFSaDaarNhPGlgpjd1UJMN68F7WJRv8wrpxGsxnrtxNtOEDSK7
1ClMmEKrF2GoAi1WRg3MDi4ICcz6a/y7/ov+W/azLG6Xh8naHGOQbiW7QvgIU7e+
yW0mh8WH0AFlIbW+PZ3gRfJvXt/5bWH1+DqBcWiNEMZmTznT009OINL1blJJoySg
icZk0nXxo4t37zxViQjL44SgN2TxLxIVBsd714+AuJ0TbvnVMUw2oPxLxNHRQPX4
lwKfxgcxwfQnPK7wDYmwWFZgted0RNSY1qqtyyrwFLmc9E3G3eYcoBdeV2gIlmsN
7ZT23iLMRk8HO14BVV5UyEzGQs/mxyNBDztLVEybu9rl4fqqGvFhO+vfx0J4L9A7
MwOSk317dZYmU629w3uLLzydzJJ7poJGPAPT5pby+tiGmGYcyllYqMVAO+qdzhVN
shwO3yFOgotK9IIHEIwsi+l8/PjLrZdPxvMYegripDJVQuvcwBVQiLXzawIGZoeZ
FUBJ6pwocHIlE+X+jeDB1sNCjWfc3IoNaq2iJwoEKtzvHIvQZCNrVZuCo6D+nWVL
ydkpTh56iyPTiX4+/chm7MKpjmCIPPwHpzv0PLxgh+WV2UMeg38eMcdkNogy2KOO
jsGtJXIFYHGNwgqQCPwMcJHFObw4aG60Lm75CdTTa8NUwoX65llXKzrvQHSikvH/
yq+OoCN3y6lbCVNAGyRt2GPigG8ZKNrujhUQAwOSQBGBLwxDkfir48ZK0UXK813b
UMl2Uv6phN82JEqvlKHrEvy8GxfbgIlpF6QsJPxN9BBxe35zprJCpajEGDU9QLTD
OrQQJz2kK421SSbk+Z0SIlUyLHykB3pPM7TdOC6b5dPDfutKr2lYRnJqQGMZfvBc
AIGpyWpX+cT4/95ppXWieSAZyaskqCAKrZL0cLMp7AJjh4NfCSpq1QtBJ07ifUl4
SYjtJcZBtkpZ9zLySwoiWFTA8rcQyX7G6FZLYi3zhlLUAqCeJwSQRgIbwShSxSCQ
JokBJrXoQphzJjmLs/Gmsxz3Dy5nDv4CU8d47y5sFpRXuAHJ040sGeHMZD3jKzJ5
xlIoBhkPmmgoD5YdWXRr1hPQ5HFGDLN+Z35PkSwA4/lOlIPj/6sCPIbMPdxVPjBE
0Kiwr/kPdWvlaLDyxfEQc+pj3sWRK2wgvM3tfHlmyq7bVRnO2gKqioIAvMg82Qsn
jcKn9c6EvPbSGtpge3MhVfCINTrUtW/6Dk0p5PVlQpHa95kimxhJwtEhpHTkjxRD
qge8TGc2wJCyyIojFFWtv7BrSPKGZW9cUMPuwisRaVszDGWZS+8rJiDHlZvsiIdh
PFKfWsHzWg4iCeWlh+0la24eoWMtH/wGs99NgPE4bUlnwtatuidZBMs/DLZvQQ0T
bLAQDVwJs5pewLlsiT9A9z15SkuiA9nh6tQj8T33bVDcrDENeqnR+NxvZmHuvcrb
fsQp9FwQu1GX1qrH3oppeZxOKEcXexiA/g6AS7shFZNbDl+nz39WZ37TbhkjAFtD
5xXdLUREWGxRnTB7ejz9Sqjk6RIhv8RqbaLxwEnSdlHoRLn8rydiSJ6L+jJM0Df6
ultWRVrK06eI8sokzr8a1CV1jKIUaS8OAeKfhspWbgsOWVZyd+XMj70GrZYkMiOS
IeJVdOkSgc18P54rlGMSMEQwyJy6mUlSZ2QFicQG6r7S0RqZtTJwfdpZR1Pv3qSl
l6yvX/6KfJrmA+f+PeH97bqk4Jr8JmKfxpbmSoLegsc//vOYdCZ10dQw66qsSqCn
HFlMqGwnb5f1RXmdwedSiEIXeiimXqZqW0YpJ2bWt3Zsa+TUBbkFfid/cepAzp92
R/JsO2FfDYwFEmRnTOJNriCQzdC8dmNuqGzgblRgbmrdNPiXLSoKxBriv1AULyUy
2uj5uV39YYkFOQkwI+eAcSAEvpi1i1gXjKvmbp7G8AuEax5roXOM1L157Wm8LISe
wpf7aECYTFnMf52jI7fwm77NuZIJkFHqq0netEcgD0VH/vh7wvnJW3VFcnpSGiAc
lQ78YFYGODUJ75DP0nvvO7MezNeQmwaJvNXmXcTPQAScar1PigYIvLMlScPkSadF
1Fxa6GYsF2FcnoEsiTyTbi7Y9FBYDAWZYxFuyvLIPPKdgKUI48YdPs2TSqWCb/IC
5ArnXY2/6lztAFLvWlum2VSyyQ6uTNJMe+HFtnzz0wIryxCg58dPkWvrYvErTwLh
5+NYefUyD4r7cpcY+x0j7PG5HklDM46cPv8zvClnRPTY8/LCxtnDdziIU0UkqKGG
R8JQr6nOUvT/92lGWFTEFykCvdWn0LBRP8xye619j6ibnuNnJi9p1nOlFKSHFSfl
co9YIoYJvXiyVkYYwIVMnd43No9RliK5NyKec0MTKJQQbvofLGon6RuH9Z45YY0t
U7kH076afNJISyyBkhy/k7bNtQdsf6O0LrO48trpqLs1m/zyQjekfsr0TatLJocg
FraJiwREn14sItkdfLCiDeX1ak+jIhwa9VYJuHt20Egu8cw+bWVctuaQ22O8Y9/7
atBCtaIzktptgZ6Q/PrJKOZSYa09/FYlxmEjcXuI44LMMMZMKpWbyfCw3Fm4WI+E
K/BK3puGVIKvu8jyXY50dP38tOwyie2vO+RXxV8fxDHGtFeaROLVl8R1WZaY9woE
G/OqeghIcEm+CEU3nNduf6KEgdY7Aed0Qs9VcfjHtWpleBEL0CQvWPhy6WLiNG2V
+e/E0zA0oaUMw9K+OXTRS2aqXlsosO1u5+IaBXIgrotu12LXHzvslUDwY+caZcs6
xH4XcjblG/vyJ6Ood/4GBKmT0CeCsGHqeizz4/0SlYdGFLRIHpglJ7zwEQTT9OY8
YkTEmsaRF9VVJlFFOQTmUitEgji+fCHoKtcWfBYDdw8x7whX1fyAcR84Ht2pp9FA
mjsmWzJONQg92/DMH2Kb49VFHQcEDBLx863jSKCXRt37MoV2d8KrHwTdGI3TmmJu
L482PIXr6GrM4rMSbUM72hrGTL2yxMZCkL3lEodPVIW9IKbeS9QQoW/WLrD5FUhy
tQWQ2LJYvVBp1RiGBPeAfR5/+pVMRD6zDlVREH3vA8zyAPBSNFTBz0+SKQrOkABa
km5N0p6CmipDZzAFzGdm4zXZTbARKR/HRxxNU/cvPTZFaw639nNNtwEXsSFtJ5YQ
OrC6mm/zFLC4mISueYSjIXLPm+dfQAEGCUKPaMQsOjqWR/cUDBKtMTuPycdLTuwH
ilbbFXS6S/oHR3+0skdsNAz865Fs0wvXdqfl9mZ5SpRaqH8MwMhvAIQ0q/S4J5Ma
kNinuCNYqRHHWEfmmX73vvlLP7Cr1+CzPHyDgCQakhVsB9HJLVjTRHM9uyN2x5rJ
GEqohXYD6MsviE9npiXdOgB69YHH7ocC0JShWX5VUAtkfbkl/RZkSf0Zut1kH8g3
FSuwpnRKROASTZhkd778RCPTLZtme6jnqcdYQcUj8ugAHa4n9WlUgVJpQfp4zRsd
enfSzIlEID+Urz0ZSoyVWcxU5sLm2bZTDX4AacPKyoNMzcfbG6bYrHWy0PeO64lj
SYSH3p0ZWiWabq7d2KqOLzWABlTSRuOCv7G+1og7Cb0DpZn052U2Yc22kdMlIJbx
mTZ3uHztIjemE89pLzIjogegaZp19mrYfOo+nonzoNoO9F1a1ScoQLHLJTvqT7fJ
go8uVYt/miFjaeqryjn6OFwjOQx5c/wHxjym5fRBVRRVF/DscqQxyxbk3hxrUUhz
gCly+CDDQyTDQfcdZojXnr6OjZO6MvbQOW4lnIvKWgV9wIZ2w7BSLp+r1aG9bXvP
cT7hDzBoPlKsXm9S10PfnfQNJECCkuabf0g5ehxsNhigcNgqaOI1eaR5iwBU2P7R
pexyYkeRldFzVQa7hAcaAbegzq3Nf322X165I/Sbm2nOzdbfeL5vUGGP1rNdEYDt
soZjDP68hy2t+5ejbzs/nRK9w5p6AVag3YToa9CuJSFx8sp2PizjumR11xFECnIS
H6qXPfrVrmdseueiULucsxE5RWgytxqHGGtcjCB6aQbrzrkwtoLqvjlZZzgb0n95
7lmoYCuCwjM+tiMgT7OAX4QHRPKlEVyqjzOvSL8E1DV4PdwXg397qv0LledlHC2w
n7dCNjIOmf2TR8v5kyJKEOHWej4YSXMvzA7zdbwuru5L+kes7b5qnmwJJry34pzf
QeHeTnayWgN99pAs9sCMPsKuxWKImu78sJyEgHUXS9NsKfH2aqbu0e8ZRIHxZMUl
/837A/GCQMEdz6khytZgPc9RyT5Mo0fHwaRdTWfRwi7xmDZAFMDwHJqLeNI6AKno
PpSAjXKVquBPuz77OhQUa+89dGbId6EeUfoT0muo8dK0+L8eSQbmgTy1FvVRRBzh
sF1AprD85YVD5Rk3ijtOJVhknXVZ0woXTFB2qEyIvRU/RQL2DPbdvYLIOwbpal3r
/ODG5UNy7AAoIScpAYIP2JRCw5SbJhBQ9h/ShyrIJwFMkjSBcnHN090yWKfsyAnv
Q2QaG3H/DjniY3s5HyMVR+vsgpiBgxfEN7S8aRJjLw5B7O+PgBx+dXXUynJz4cdh
l5rtYxg8VuN3fS65G9NdBmLAey/YdK+4kejCPis/fzfkUe9AMXdMTOLQ9f5n/och
Nx+gu6/dDlVwM8MTb4els+bngKnGGuyCOinTIXjiy58RfSprdJhO97w8cEv38xrZ
W7ohFrKu2EG0CC2wQZZOHJATVji4GApte8FvaLjLDFMeH6MPmr1FFHZLPKbSMyMX
07PRSbVPo7nmM1w90swR55drNYi3VNkMWbhviv8Aa+6ORGbobUp6+/4PG9WqDPHr
9wMRuAEoW5I35zGQuaOoGqIDxJdKoHJgjg2LYku335iPjbNZVGugEWMu4iY3cGAR
D6u2fh9TOURF6c/zZH2Tk7ycaH/JrtPbi5uvEPh+vOFijrMvQEIPqki/T9OAh617
oobhwo9uY6XwgPd2J5behPelFouLNX9/N+XDdUbU/DuvjU3G6RZcDwkYvXcdYH7L
cSUtilDpxtQ+3kUiNZsKP+qw2gGKQsEeKJvzUf6PVkhDcSMMjza46LLEycbkqQJw
Mk12P8DRQRXQx9UBYfm7QEwRPxURUUkPJL9SOnOAYH+HEkpkwMuGckuleUWTpr8d
7GMKCpkskh1ZHXHcUzdYnUpRGK8Fu1lKNFxf43QSNeP1Sk8GxxLc+UhZ3fcmVAyp
MonFVPym+0GGxcSqQJ0aK5gDWn6Vzf/hmg/GdIxeEW5YJjSRlIIz/7prWSWv6yQx
xbAdUxUzN+3jTyslXqKlK2RNxMWr3ioKsfm3XWyddQu46Tva48kextaQfEoAIBh4
QWF9surtMnzpuDiyvnya1k7J6/LDprUqhbxTOO4rKQDu3UJx/eeA3/nPNqff5tNg
H4gWcVTTdZqHJaGpsSDbeWFwg/i6iscYyf2UaCRbMgvwFCVnjP65vWXT1Wj+nM2C
QgQDmICl87MTLZCEqD1kaHzS3ciylw77TpSI+IsQAlui+oyrmAemhghIdZwdAo0d
Q6h6GwGG2M/9vz00qFSbgbYAzXInt8Pc3OWXOxFPGTCSH2JWO/cldj1ShRDxsJ/A
V3pohgScDEYlttEn+ZXUVNzLhy+oAcIHjSwTQBkkbyQ/TrNKx3+PnPzOl7cPktrB
7sJCGfj/iMqMSIXDVbRaK3dhn/Ks+NAlrQF8KiUxwq5qZWxtduZpgArB1zLg82gQ
11HEgTadUKwDzskc/wWYzp7IxJMWGvq6+bcmul1R/t0zw5ktQCB1iPoSgn7w+nb6
QgigswmLDuN7KrF/CE1Hs1JBYdA3NOgmfvXzDxP7s1PqnHqdziKKjtEt9l8t+4Es
Ct5MLhmAnVdKrYXYHt4L9qhGiblVaNlA5J9XSVYTOwjkNF2rq9gLvvh0hcO4etls
f0ywvPvmy2kQ06Gai3BWuFzao5SZewCe0rh8MplLXkPRIOgd2ypvBgIF24tHwTyQ
Yo8joB9d3ZOq+iVzAChFfRx7q73h9/0+OI7cpHVAZekjzmLJz7cTsKHBGE3U0eBn
WxVIcDZPVba4aW6KVKnpXgARloHKieRqAh8aug8G/YEwL1x65Khw76nXAIeLBEhn
S5PQ8929TGGmDY9pPjbNbiizUpJPNoO5koGM+ipjqmllJhGN6OBSWhGbCKpSWSU1
kc2V4FOsXPp/1tXkpOYjXZFaEYlaQlrRF1YXOuFMYFzpvbvDgNhSaSDkbqBMWST5
nTlV+kpK+0aGdtV+8O7Z7YWAW1nLdMDPTVVyhSE6kcjJCDe0TAVQQ8M5F5ZLSxnm
C3WyEidMN5sTahre0F5mS4sKHke1bEJvIq82be5X0puw4SRmKO4eL0uiL7yDYNfn
qFLf/9QvtIQQzTKmmeHmd5jSsyJv5IK9A87h/6sDEnyIQSfahfjd+46FHNh+ytbe
mA8VwYeueiOEcYPYu6m8H2AxcteKfPveVKzABQ28UB+V935S1r3txNBHegIExVTz
dwnY/VQGYlVFXntWEQQzZY0EusawVkOqQerDgrak+yxLrNabrbpxzyyUq2CwQEze
Thu/EFSe25iBGelzDEyyg6CeG3qWdmg3QI3WnwQcBTKHdsl/9yaYxa1cv7umoy0q
UaUEgBEoZYbUeawYVKXym0QYhEclM4j0wzi76iWuqNHWcE8L9o/lBd1M8AGeKMXs
CU4xRX81YPJhxIT/0bwOnePsPt5lFFEk+bEIXO6kZ/fDgjlTCm60+eZhhuyDGF7B
txvpkj8OFzLXmG1GbRdankqcFEmro5pS91Z5bsHJfae9FyHojuVoPzZTayj+M/uA
HrWGCd8iGwcTeep5q45u/XH7/cuqbcGXBZ3Rd52bKjKi3YyjxOyByTKQEsM+eGYD
BplcCsVs5kuUgOZKQ9tCmP6Qwt56Cxe3Qlh4vwNUi3lmPNURVL8nbw2FspMbmmCO
+FzyMop/V8eElDqUzTmLRDe5xVeXCk38vzN8txTtUst2BxRmBVkBWN3K4M4zt+tO
Rz/CqJ1/heKrMDRtU+YjcpgYmcnC5LljgXnJ7yi281PveLjbxVSfB9OG4bvfuAFN
Zq0MBj3BKQmiNjTKzqO/KvzALwCNAidGsgO1DtdlkZGyZ8VYSfMeLDYP8OVgfKNL
RI84MeOcTKcLgEP4yc4iIt/jh15UFS7w0afk6sdpNAbseYvHv5Z4K1ff/2qN6T+V
HHeNobifTHKiGlBp0RGD5RFLOW7pC8VGB4AWYiVFMS5SU/9Ov+UgycU9PUAIUmDz
7pk650kya3/wgKW+Kl/QCTC5HORcFSRW0zayHt9JcPvKHW81fgsUjX81jwPf3vaJ
SPeYM6isrJkwHaamQ8MQxeK4qm/NITqitY51wKbgeHOH/9ZnWz5gjiTgtAlslIf1
02ImTI2opTf7cvcgPL9PAF1KP0Jl7k3/tYq91vCOSWxAL28+Q0XDlcocpMGcgXjV
h41qhk30nvzgkJvpvTjthxwuBoqiJPDFXd0VMdwjXfeRWSNzSTX88trIHHCidNgE
17/P5MtVRa7eyoiNwGw/sp5DGH6fL9WiKLi/x8m2qIiE5lgq2LqhN33beFxC4+sS
/Ovi5OSk3KpRzU6SeVjEeXRrKvG9LXzsrJDyUllLz2NKE7Bt9z4rWA3mKdU5dfc7
XtZSVu9Ma6cwSwI5gP6G3GxKp70TyTtT0BCPil+Eo47W8ufJ6UpSYQaxARJ8WCat
vP3fJp4Fy6PjDkU2CkC+T9JraOWRMCXUIru+IvKGLFQvEcLRpGYCkR5opMj1yKF8
Nsei1bZkTo6f+0zBRPqsBLNyjB79OB6+iNQ2IM2QIoXMTyUVWS3gmdPRRBgN7I6S
Xo1rKslJTP9awDiIlH1I1p049l5ax69np36FtNWQcijAygAzmEE84dzfcEY+tZbL
IvX50KwVa9NrPSDzEJgjLX/SkiNyMzc9ruOV/2CMLkzs1GaTOqzDLd5zRTTi3Ji9
C+sgm22kId85UTRgjCAOWfanhvIxePmWHTCGZZ2oyuIK9TKHIiTSiSAP0J4puSeJ
zl+oD8lT0OW5qVyY46+5l3KbNTwYlPpDmfT06BXKW1KazBY3YKHpVKsyz3qtKyZb
kfj4GyRsas6QK+d5r25iYT69tLK83NzaMgurYLioL2RBMuaYNci4ExxYnqIGyJ1P
y947N5v4VYE6OOMaruZ/eWi9Zoe3qN0Sdnjkb604uQl7hj+tllPv0HS0p26NAuNE
mknRzV3iiF7bSc4Dd0FIAlUht3LlJ2gMmhQIWLtjNhIMD9Tic5CjJZDgR9RZ2xW+
ND/hhdq+vYma/6/9uJYGJChiX7aKpDGA8SQps7hw3sXC4CRXED/UYmT3zCQMoa2k
41tf5QYk2t0t4MaUKtiIEh2MjOq4X9goOCb+/1QrkPyjRAqJSux8wZdIQMy85+Pm
Vau47lT+7yoD8x2TLpoylVXhvoHjUgBfI4O9Wg7faJyS5elrkNuU2Kh1TnPOWWsQ
CRGhGqWPPgikhZu7yc+HxtirSweeP5p/yYGYG9iNRiTczCngU+v4h1adonkXEJ5o
k+nwKYTe86piNHx0q2QKKrMHRwzov68dfPzTaHtvEkE1KZLci0xZTV6U2Hyl9RD6
gHhuTCJZloJTepJutJlxb+xk8D28N6P/T07xHZe6//QZUGmIAIcVck8LxigpY1iQ
KhRwhCMgxaKprK7lU6FxbvKpMCcJp4sCQuG78+v7Uman/P4y7lKie+or6nmyLEfj
PLghoikEJJ0AVM2J/8Ryn4ewKrClDaaxDyx6TL5Ci/qfYjHkBfAlneeR0h51XqtP
wjKE6teibOxqM9i9f7K+NECYBItKZv2vABHjiS/IBL7QfsAwyeeg/l9MT4wMFlYJ
OEqOP2+hrR6QwT64JFOVOjWePA0e5yDNhNrY0z1jU0YLZsoyUNpMKxgIljtq7SWM
yT3pLN+iRMcFh/qM8HfhIRABKw5l9EZUn1K5uHLdFe89nZ6YqBFfrMAADbY5S8R4
Xvg8Nnx7chJ4nbH1mIvZaYBrElSTAkQA1iTeP9FfwYqxt/36KaQs0Uv+qOY1yogn
x8a/W3qtdjdiidqjCNq+AQwI6cJGmXnwp2G0OFuoQu4sb4yamKBqZXLXaz5ViZML
Nvo+Z8JllE8jnDrL9ZrHktw3rQ5Iv/JuOpQRt2UKFe3u8hQsbkpg8rf2j5J1yp76
cDz6QS1J19thvOSgDUcvfA5qwv6Ii/p4IhDA02SVyUptzwTayr1e4q3wRI9hnUnD
xmV6U81EfQYCv/ttZUkcyClv7N5+Mg9mo1iyVYaL7JxM1KiPZ2MgF8IN/uJx0/Gj
XviPB+rrUCBjFBaT0kmnyAF0X2C4TEVgWq7IYvtW9y0tJW4SUhCq+BNYH3uZBmDx
5yvI8v6Mi9YiKA4qjVpxtf4yZ9G3pkq466s9y9+wwDTeo6yAPpBGh8Tolsb3NL4N
KsPb367zY3JrLqk7oc6bXgp0V2MoslniTNiM6z0UB+lUR5OjOGrnfFTqin97gkOy
p751CNRqsUWX7v1MvYqiUgU5GW3V85Mm21u6cSEff3c4Qm+hJwkko+KCZAswvTmk
RENwJ1pbfZ8/0lQ+ZhrAfK4V1fYLQB2E4x6g7eihUsQCJmH4xMOzwj8adLHz3VOY
W43hmn7m/OD4KcDkuQCEhIFCaylzXuuraGbLaGE1xB46vKV1e+iagCWz1uz/QEZO
575cNLVNuOTaphq7j0ZfTxN2/CWSXPOAFIZUBDhtJkF7hPEjhyiHSHHk8erV436Z
9gtyEQO1CbTiqR6R77eyxyiC7ilCEBEojW6yNtENVUK4YFrqELy8CYi5iXIUn6IV
UCLFs/lzG5cxWCXxB8njiTrlvkicCcwdLbCNrGaiNYBeU8DbtyPunb44e+V/fgWr
OPFp22pQ0YNb+MTnbJfKtmxpH3cfwy4Es9EbuOqWPfennuxhhcWCuZyAyrXXnh8u
mVGefCU00GLHU+qkkVtBiAYE8lCYD7XccuniyaFKdDGJ+h1+4tSEk2U/hqU9/RVL
/Xco4JtY2ZnmpbeiKavVPERPwenRBI6aCJtqCYMouVBTOM59JsPVrQgQVXUKGvsV
Cm3HxXbkb41UDEiQPO+DwZ55M+o5E3UNG9P+dlZvYNLs0evNvbLs2H5dAiie2Q3a
kqhbYzWhvelKK4KPmhWToZp0Jlm8PQgFMDOQudrxXLhOnGrWFyAKsXip2civ0O2Z
gapR62kH+xh3C2DdZC1wJyDNIJVyMpkEx4BXwUyqIOihm4VRWxy1wlT7qAyDK6i9
CBjN6MngL5HJS2SrTtFQgWLHutzOnAVIO2+SEg+ntsCr6g9Ji2+8CviRcS4ptN7z
kV0p/kj/z2Yc2tqI+DizdQkBgR4/6IfKmv0V3TzIFe11c1ENCNB6WKnA1WN6Kokz
svkuqufiBXRkumfBH7ivxRxajh/TNYL2RVD+vRv++Br0UpTTxHE9iZtwUpTJMEsP
HY5vXDJT2fDr6bnRaQwI9YB7/JZSgv+1+dRo9zXBJZOlEqIYQht4mEFe0jR/aBga
dATqwGkGGd0rX4gNvyrOx1G8Yf7XXYolI/HCeZr5oFh5aWWsY0Wlq7nMQg0zjn80
UGKFWzz6m90Z3Knanz0PZHsvhw8XPc+4M4PHPIiZCQvl0VFmLnKCt1JXoBGBIPAa
j7OnTaBR/Rd6nRibHTxuJ9NNWLt071IplLQTfCLkN63R1D3dMbpjPvSYYlQvBqbf
DO3ZLTI+bRVQ0qZfD7DJ3/SXdLzx9MkHCxMZAlFS19dMpPbyCQXQRRULO2B2XOdz
/R6HaCXi2/Uz64HA/rrcBYREn/0XN+a0YFMWftAAf4WgwcyimrN7VZq3c/LWbXlp
fKGpt6V6un5g9QVGRPZfCeH3KtX52337xxa6TuPpYrApCgMQ05h093hdvkApThSX
kniw9zVQJGZgF6jXLKeFrUAyRPIhMZqEHZo/Vlspf/nko3NDSrv4f5AXj8kqkdFK
3UoJFXNt53vGARqMBrWbsHQU7v5M3iK8glnHptx4zt8/HffKsDh+1GVIf4tK/JFu
0MdOSVobXtULAZRBPDjYwzNWkzYLJhPpBeVNIvztwPN7A6EwVRT7UIoXNRLlrtdE
q+qpfImI5uInfFwGJAA1l3w/aZJKCewJrlrXtIjyq440/ePEDDFUM2zUvssCc77D
Dcl9ucm8zogyvpsmJKTc5PvJKO0Rbh79gKpzq3oocsIRYPkklSRzOFYyTkS8YXX1
SwrfYgOPpmHi6wCJcjxrynM4b8b5e5dDueIU77OpFDUyX14npHw5Lc8ZfOJX1iSv
j5OJI4FsDxxYbTo8KC56BAlSRAXujap1xrRG57jwYeSdkd82Q8+dNCP4w12G45KI
dKYlRlxZ4tZ2eo1UtOKhN3I6MNtNxYSzdzjGAz5ussdLzUSox8hvaWxqip8lJ3oD
gORsRS/UizkvC60ytSO7L3wGKgaqg+d0G+eTNvNmaWlKqiJScPdmTtK3K9QNC5dg
j4Gwc5MylMcor8S0SPF4Ohp/9ex5hshntf2HL63EnuFUkaB1aepewIRtMvGuyJZO
jzERh+3mm229j4A9+0fuFdIDdZoTi4UkVNmDg92zscLmSuZF0x5vaOTspvK33s+E
r+R0QmuNPtyNnDjHAIkPApveAv8pO4QZSZw1XawvltU43aEihr73BUSHI/NvnRBI
Nef7tyyo4aQtR8DfiGhmjYIEwA1z+M2gUE3+dUJ2sShg6Yolznue42WD/xHLnLg/
7pCwXA8LkyniHJkuhVGeuCgf8V2Nv0eMX2XDhhwS9L85fK+70Fq2ngwNccp3yCTs
+2ua9D1t2pyvBm5dO7fAzHYJE3HYDdAI1y/OQPUmPozvTiIZU1pKNG9HjKjYXAmT
zPBcU9KUq7yXrtrKC/Wy0DXFVt8upycJV8SbqzNhEbNWIoZ01301mbS0L1AT8L2k
hcB2XSkeGm4A2e6MpiRos4ZiixW5xFRPBzdzeXqUzdlBx56tMUVoja5gnD/gc9gO
4+9/G7DKyKQcSgcL6PbPisP1T2fQuAvp+OFeNw06fFiyuoEJHhcGUaXjz0CMPILh
dDAMT2tguOw+vqxlQ2IxkBY82dVjax2vOdtelHVmeOplWbcKBK2Iq7AOMiHYgrmF
cFmi5tQQF7wNnB6+/tsHvyb4bvI3bxbEfFvqoBAdhHayYlJZlK5j9/gHnrJ3QaYv
849piRD/OWqjr49vlTpNk8NbHJagIgxiOt7DnxFg8mCGhPnCtPOWjBWkJe8ckwzN
5x7Mjq28Ofg7Gn113kKyMfx2JemmT94HEIhbTu1mc5TVz5jArLsBo93yR4wqa8kL
dpZuB/RHrzXOSsx5aNT+1CMDSJT+KG7qtgTmo00xnSjiBQv2ZAchAatUl29pzgrN
PLjemAfXXyEdulLxhCO8QaycXx0rVLXbrJUps5/UjNs302BpTXPawhXlmhiJVs7h
6nbPdmNd4zCcZ3SzDfxomgrmldsspUI8JmzC7wf/Tuc+4BUWmvnAM7U5xa6skkvC
XM7LVNS6pfljCPesYVmHBhfO2QFFpoySLvDff4Z09/Ah14rObmhD9F93Cvc/OcNR
+fr/XBsj03lTOL7LL6cVGbY5sb7fzXm58qlhYkdIrbUB9OkGgItkdv7ej/F5izpa
5sdWMvrZhIlW8zZogyplysQ2pEv69qYhCZ4WoeBXYbCIvyxqI2ailtrxawf9YX3z
/i6UMnkbQ4OT2GxE/v/NpEakVu1y7TmDxnjzad/bOmAPSRD/yaaHvcUl41xrY5mN
VnIZ2g9OykhBPZEU+9PPpDXjATvq9fISzMlsAmATP17kqfU0aeZJU6gg0DTV5nJf
+U0O4vOnW29h7FdcyRuJCVl+L7yAVgd+dOz6KBfuGvy3Y65i7AfgwJYPvmb2Esyw
T6g1NGhqZq61iRNzlXjeUASdoeSnxAjMcBQc5opYkFUdD+YxFtb4K/pABeziDeR0
DERDqVekdrmev/HwgLicBRi6l3te1e2KDppTilCcsIX5IK09FO7nv+HU+UF0ri78
/m31ysN6qukHoxudBx0G+EePtOVaLaPVBmEl5Bn7n18clJto7wT34n+vzpBqcKog
cK46Bg0hHUcgzeVm1tCual7n0+bawgOPvuQ5TokFtEMsw7NIod1yuEsuGRfNWTio
YcDYKikU/nA+PJzGvOM3HT3K7T5/p+EdLHowosCsEdEo86GpkWKapN0tXVNuBaiG
k9bCXkpNRrLkZ+fXsPqbsQcr0LwRgn5WGLng2BACdBDsthDMrcwzh+IWGn6eftEx
hE/PvfirJ2+AjtzKfrpOg77pJmEs6EVV8y01WPTzWRi2EWrgOnOS1GonD+wl5xFC
KMCc+pWpkYaO/jfcxi8KA2zRcVfv0hXURx5a8bEECX+3kWROMJWw72juFtVQtns9
RJx1FJxZ8/vnKwQxA6k+T1pqjmMXmUa58I2UCcmNLaZKwbqsApay72pq6SNi84uQ
Zs/BMeKA1iE4Kj1yuvgZXGep4QVxjOQs5JHk7f5VJwK7R2Q/3/Q+2lxzfszZj14o
OCwaqTVs+yfk5FeG94y98CtQW5tk55dQXIZFRsDIK+sHWtH0BXMzJtITAprp15mC
rXc31XMAapbpA6mVAdGrbDkEIOoTstg5PSvSDf98RwbZttGGI5NeU/w55PmqaGfb
KOtbnoGfUSaa/+hZdh1Vqk2AAufnxyiRrzKcc6P7Y+uF1pUvpmSQ6MhKVuRyEv8i
61K26eV3kUsZ/3puhaac/W2adIDkRPW/Zga7Rlw5lZU5M1U1/zgJ6LApwCO3J/wI
h0nSI8TGay7baTKEaCGDset5ovAXiMzl53YFyLyMdEvo+12XXF1iYdjHUM+r+vW/
rKoD+kcNSe8b0snRh6FOna1gO/NG4OjVWOXo6Qab71/hTwQkbs4si6cWUO0pUCYg
DRb8URsBh9fNa2tCrcUapeVCDG0iuSWBxZPbPupNhQ6Qfb6HONaHXfNCPaAzyVW2
yOqulF8AG9Gs9vhbwvj64kWSQkA7D67ysl5HZ5UzghWlCZwxLxaom27TmGk26MBU
IhxK8BOx4TXicKyywmveecPSO2gJ2ZJU3MwrWJH8OZ2l4SUE8kLiI/LcgwOm2XvM
6rEjJXiPX/Wd0JV5lWmkRpN5livZ/Mr2bA21JYLJ77lUpZSiOwt44n+J8vqw/TtI
lfrlPFwjqq1ZV09BfddavD6+USyZSfkZsg/Y2ByoZSY6Q+1DQXlmmlvNnzT5z9pQ
d9R1AEYkVs/RzTyd/yR54JKX2+svM8S0At7MrtWy2iUqkJSqiSxc/CuI4kvandCB
UcPoa+rXeAXUsOsGtic8ST958BPDf6rHTiQodG7Oq9CWCBzpJx73s2ZZqSJJoORn
93Z9feUPUQH7jZOYu4r9H94If50FgA9bvftqsTdEvPrn37coGUD6GUiOIPgLqnpc
CTdFmtRiAKE8gz/325+J4yq9FccPEqljsT5WtcDl1f7ODYUT54KTXBXUq/3/yUtW
slLvyAAFppAeMS5bZCQttco7u0xa3m4ljVud+EGHZ0Yr57mwtxRCL/Po4DGrxer9
ezmfEq8MYf99arpuNCulsa3erb1J9slVIhIeWg2ULsVa2sGF5zo+eNO/IqzaADQH
Nv0BP/jNQqcTYsQ5pYnDtcpmqjDwo639CkfHztlmZpprTE1rW5BOR6YRZ6Y+eipI
aMTN84Pb+DGbz1KoUNisnMSOQZXsXx8mXvUtBep80K7XBQHXNh/QO2BizMhJnFPm
cTD8N2yxclZm1znL+RtL00Vh663oZrlLDUN+Y1o8VOIVIVAVc7RV6UeeqhkYHhE8
Hxt/i3gEYE/c6ALmL2vpJTcPw3SYhIxcHVlg0tK8+NOPXlrwQGCtAYlq/mt1dmM+
KpYTGoPpOD8yoeERMaXtpjslSyOMxkxv4OxeDns+M7xkN1m2UrWY//mJDdc1aR1B
oMb4S97iNYyQD8ZHfcPq6Q/NSJl+jHupwRr9bqGfmvDaZPoHlbpXrSztpkAWL/z9
y+Kl/qT5UFo+3ZjpQyfb69EfzBtj/bkHOIDXC2Tx2pw7Fg5cJ3YXiwZJuJn1a4sm
KzWC+eKPP481EiJuDAmJIMNZT0SUdeaYja7qgbhihqw3xwLBCYonXsQKb3Q+Mbk6
Q0ZCi/4kFrU2daqcWSNokdi3qansHgQKBGPBLRRDs1z6o8wKrAQRgBEPAxM5LoAW
/Ha+8sYOTezmg71UBuisz4zW4T95dD3O4JZr1laVXLEzJftRZtzoRm5jHvvnInjx
kIw6sQs0ZClW1CfAaxN5bcL2sBseMS3g1DTQhfu5yWZa18sxWRGmZEFwptR0Mga6
CvxL9OJQ4OfLLyrr95h/y58wLf7Plg/23Ms21/xfjWvFMZ5JkEYm1IKTAjQyvUcG
yBE2LMnP1Fej4dlbPX0LXS30S/Om/Cj34SrTIxbUg1epfsMJd+T9ZZM+vVpNYNnm
TcmqXL/l273UKSPBIrkyedR9rgXZYVsCDRqdswu7eC8+xuXT+Kl6blmQM+TBchw8
RqcH6mOYgPkhKbXSgBUmkvLhKhMTTS6akjLuBrRrXxLfQl3YBipbxMPeU6BvvORS
EFxOlSPVamkBEEusvVHlvHaO389lE4jbeCMpRQtc6hRflGOjTjGHChyUfZEYum2g
/lqNVjYNVXOgAqY3fXDy7mlX0g7+InIRrBHxLovUm3AI8NZ4MK6WMlMLY5Rn1g7q
DIpHeYujHQRHTnef/9DOrCZgmHylHnwpTFYVjJtdNhPkBkuIgII8LNnVxUJIuZ74
+XNQYNJzTIg/EL50waxzBfaq4Vk6NQOIqQPzZKgOUzbLWkr4ulFnQIdTizYxn2f8
miM1F2YvClIi7ZIwavVtzpKj+UUNYx2EVbZDi+wKYTGhMOGH+nh9jB89jm88uKX+
rDa6097Btc+eDkj2Xe412TzaXKu82mL7eY7N8QEHMN5/NomCFvlpQddQmMH6TL/w
YDrDUX2vH2F5HyZbq/7FRBkVvrceRHUMzgnTeoSVyoFoxeI/OdygyoGKgvMNb/xF
W9DEvIThkI84to0Ie9JyCq3s4OrNMX7mrAttzMe99eDnw713AZLCWS6Fe9TrMbGp
rU5bqo2v4HC6QxpMVxoYsfv24qKTHWOExkmMNB+XH0Qi1tvggXXc5nKWluQt4Xd7
KqJkFP123lt8VT2A4Gwk2SQrgkR9l8AMQUMBBjzI0vdZvHrzVZnIKLlZv/Fzwwte
5Ht3ltfwpFFE3gnUreGN+m3S+0fkOiXSY8sxX8+0fqbCt7VCY/IYjZPljiN9rKLp
ZU5ks9eR3EBwBb4WQHYbdMIBpnydRSyySHXDe9Z5xBEeeID3KYdBRDiyKxzE3eWA
JmDGic7RdLFm/ryPeqiwuPnd2Wc+HIlQRbbVW7/vjyPq76Odh6DmbhOfFY+CSAHP
M/hI5hRHbP8/acHp8bX0k1BTnnnY72n76zEdXl9PcTs9nHg5rxTszzp89RvtNXzk
bycmLUBKIQEszSd+QTdFYEQJ5lKBTN3HU53BRE5zx/Y++WJTv6oZsRWKUaN9MI75
8VL9vyVXi8KNCTC9U8Sf6TM1AgQfYlLVIvjhQBJNUHS6w3abQ66/q1RuAVRM1Q3T
Ab0lzSUuhAwo4cNfbXMZsNFn/Y9rb7ToMH5pDah0/e+VdTtC5kKVd890EW6kRu+B
Q52bi5OlQyvl1StZin5AF+fD4R6pOZ1NEkf/Zggo1yp1xzhXEss9PXJuxwDUIJSY
LSu3RQL69zJQhI82UxNLcPw0CsIAn9F4Ljaw+qD23st6dGOHcbX5dEi/F18IgikJ
iuLMULjwtTTj3OAOtOyyMoNuoiHt+xFKl9kaOeCP5T3j22BT1wP1HbcDN6FiQ6i3
Mq22xRiWZho5Sd/Co+jE5vnBQAKgxAS7jNqy8vDRkAHlNQDgJrYuMxfGj8VUyYac
1c864nVLgLlcTOVuw39JkbrFzMiWIaP+OxVTHgz7WJvGbRjlGEJg9tU7rptWupO/
uJVBGW/piIq3heT7rn5vALCFFNokDa8YyQhfdDZJDz/i7LIFLCSPVjZVI7Y8NzsJ
ilWmJFY3vAb33gUavrUkXFLVk+27V/zzZ7nt/yivmxiTOMF0iWm4qczCCVCIQBsX
iVznG+XrjxAZqNNcS3plPqAw8I/HiLpBvww3VWCa2IVHL7c3/fvAS5J9Q/PUM9bt
NzMacv3571rHyGbOnpMBNM5QsDQp14RLS4zxHuNqQ4fmZgMoCnZiQ9LMWVuIwjpW
0R14OvNgDAU9ISkquVPHJOE5eSyG8/ELqx3JRwT367ig137Cdz3t6djcc04Xs6tA
yiI/PCY+/MkNt31Be6kDA91kR10gjuiTNHQDm2yIgpGuSxX5erGCdctGOwh3XYsI
ylAB6UU1Cvu+iPwfsBn6v8wJ2Dv+zLjQjDNY3Fy7a6nYoQsgoCbbK9Q3boRcxUgu
vH2HnyK9vI7+YHHtKPIbTzeG7HpnAbBn8UWBcztyd+HG8WJsSMlwL8TZYVp7HEp+
ZVohtT8kmfi9zeqw80zJ0goIOYrgbT26bYUS6Ie30RibIdF9HAhxR8qa3by0x0xV
t/BENeRiFDKLlyozGIs3afDc1X7JC9L2hEMP63wfRPRYe3KNhiJA4C02xnaOFGuC
Ql7rMma4mg+ePdARe+Jc1kn8YGt07wCnXg79VUDhxrB+XzP8SAFrLDEW6Ff3uUfr
3i+v3S5GccBan6aUguPZmOTeSvxZQ9xWa/QyTs/yJh/vDIwWwFhsothXldrzsBpV
Qp8xFgFwfMvFxkeoF3UzDaB7emowsBqIz+2mIM8UJTAxZBm5TmseM8lRMxHGtmDo
59QlAkwsXsTtrhT54kJ/crKYn/Vix7HcnRr9tOs8zRRoCty6MYv+m16xr5yqtxfJ
kvTwdfnKTMgEgx+JztxUmH+zoWCklRrVgjs5/VZHkdz3pMjIGdHQzv9SvI5Akexk
oE4DK7a5x6DP86F3x8iO3vNUQw5eom2PpneI0tRTT+QFaqvqk7JqrrFVrdQzDZBc
16Ox/erwKYGn2Zc5e9eU0W9Rj8ymT0U0Jcvra0dGHEELyWlk3MQLSDYTHfxZ75fe
OlnAX5qlqFkmexDul0LQzHjPIIeFwyA+nnqpA5dZkG53GeU7wj0NOgwiZ8qHJ4cL
XmYp89ehO+GSN/MNUw0j/Qwn+c1w9owNcPK6spioT60783B8toub9aIFcLd9/boW
D3/vu78Z1RLfnpSf1NWU/REBPDlA9OMFoUFDlXdmewV5JyDA3YCuz5ShGpClqBM+
2AzNwmAePgW9C8HVc3fbgKo7lGUFbhZWdJ9iDSREGO+a3WvTDdAHHTQu8u1uAu0M
X/CWQbdox0Uj1JCqK9o6xhlUCsisVISxHAww//122eZApFUx32MXaLt5RK9MBMal
pWcT1mlutuIJIeJWYAs+swo1xoD7dnwlog6BJ9ejZiuvU0VmA4mVXogafrUid5GZ
vYOcZRqTDIzywVQtoGBf19aaGKvQQNrEg3VXYt9sUlhWjNhadLfWovcRwoHquUQ+
kZ6dDtjJvCv16V3A69M3xcIvDUacFuc1PohOOKsJoIv46LBmD2k1gbCVB20bzK+M
UF0bTOHZVGQNulgRR3jA3fRtXp5TSVO119YB3+IIy4LX5EyKRaIsg0psBmThRxtt
7lzW3LBFX+mBjXlwSFjU5hbzXITVdWIktuytWs4ADbBS73zx+A1LxgAK/q676iiF
JCi8J64W6jAVj85nT2ZlR5kpp2WD1wW5LR0IrImNX+jsU01arQghvKLy6fZWZW9d
A9y+80s+Jl0a9uN8KSpq9uSLqs9wvjHo7UCeVQ6RSiokQPzBLPRA8PPphYIiLbeW
phHf2jJJ7hz2cUJEJx61HSiUPdC/CtiMbVBd0U68WnGhaGi63lnpVYJFqTKIaO73
XBk9AqZb8UUENaqRoZxMfno1vMzZMqGHPuBNq3L4G7RNtnw3uh5Phg79aRWNp2mT
gkbE6LQNtbMD1vJjUpMUUSgEKR17M6Wj0M6YFYCClZ3vtKUr+VzxXLRg2sr6uOXc
B9lj6Bz/62ZDGhmcKfXxHeFTsqOO5DZS98AhprU7nC1AVhhncvdiUUn/P0dGmV2A
4s6FO235EJ8lT8Qgg8rnF5zzPfEMXDyCaWJkNMKGR2LCH6Gvhm6VwXLPlIcDXy1g
nu9kucbqRiUW045S1zCIn9TMaptJm7MwF/wjaE4ajtC4z36YNgCiGigpY88JmwMz
cvd64arzbXZfZWAg10Nf2H0ZnnFG1P4OdVn1qAR09yPlIh+E8DV9nQ8VGq+8AB+E
p9oVCW5zu1xvDe5jMmoK8ST7QxBt5YsVzRFwCHsV/qwt8xKisWqEyhOKwmDvsuuq
jqsBbc4nCGXQp7ALKUW3O1eOAtXf+Ptwb4JLJ4GEwy90oxqST29//fewCfUb6giw
e+jxy/GjhW4OAPA31v4Z2DR3G2s0v1jnjzUZ6sGbrU/8uwjO7jaa25B1BOHQeogI
58VZ571SBJVmpB2pPag7rYVGLAbSnPkeQRldaBJawHznMOsokbb+n+Hj9/4ylyVR
W9w7KqmuyZdG9yul1Ihd1NPHX+DFoTob0vAGHGvc5lksfgjQwcv3I+bqLFdy16Ci
lj8NTkistAsUrpk2QYXPZPlhpBpXyJuthYw3XWomnEkiQQyBCKQ5uR79f5eV1jHy
sNbxtfuPdKVIfmI7+iv8LsF1ifKTf2CSNr//4XTh9fm7AeDjYNpH3LEODKX27flw
vAulGgPKwSqpEOpwKm/qiviN/BMMv60+JLTwFwNwzbaKhG09iAwlqTpcWn5IuoJg
PdyMOcZ4K2qCu/BYoTxzHA36MD5URJXJtChwIjiTnq5HquL2MmNlvmLpiFOJIGTT
xmBVLCQlW69ggel8HJovMDuYMqLeCcY5WJZ/GhLttTAsCTWvuJwgwZXthn2w278B
6RuE7CdAQu7YzPHEnDovDEz5AZfy02Jvhk7WlPVOA02qMImJCvWkgRfRSx37NwHC
kTfxcGcPAF7kDoyz5VphuPmrYKKTR9JYENmfXqAc5zo50s8EG053Ill+oejA5cyz
xN/r83BmBoHANU3SoyiCVcE81Ew/GarEU7bgEIceoPI6MXBBWIa+zqaErGakz0XC
frAAH9j9TTSlL5luD4SGEIybpdEii6l/bP6ZLUIJNUm8sqtnEVEREn7js2s4CE56
gYdneLI4mQF3b6wybAqDS7xemlZ8ekmidmvSrAj9tlGkysJmFDI0drHE2/RRNfMn
qsg7v8aFSgNseCQBdHD/zVDCzy08wlUL2+bpEobmQqcTAieKdWyVQQumOoBuSX37
hshlmna3GOsy6VhueUtaz6NAT9YWohLLbtkxtMHiPmvlQzXUa4HZ7kVO5+wSI3xV
dqyYHYr97AHGgiMoujApyR62D6NjMWSRCChoPDLeEbzQnJZTa6kMafaxDozORCmU
Pjg1RV9oBO3rxulf3eJdtrITd4VO6tsSmMIYFDtuxWqNOHm4xfgyBEBfmWim5iAb
43lHz9PyVnO3f63MqwGSR5G+mXWpSiTgY3BHXZzjvggWhfmASl1b1vnaFUxfmn5q
PwseNjZvIsOqpFGjbS0OAhoWD/kU5bxxU8lfEWRSwIXaJ5jNyPQ9a15HXmXYK33R
mzgdzDqBeUmodadQedeictJ+Vfb/xyCT9YogRAzLn58xKyAZ+QI5whVXDK5WXe3b
R3x59E6Ie9vtTq8s0ZTaqC/ZK/sZ+fTvKr/3wkO1M1aY6Xo7BO9BHM8KV8F4txRr
/mqpbjWDbkh9cVHRVi9ivE+QLyqkrBAJtsFezIAJzRfv6gjib61w6uqOyLhFp0tM
5fi6fXuxdoyZryLhtitAarkZJn+GJu2WLNZUr7nYiHJ/4bRC0FkUPACq2799SBl0
oMwFGR0fAXQi5adVAdrHHTFyqQM2XYAYcDrU6VFsZd5SIOP7WJBo95/Hy5ovKI7X
77r8o8eLIpXZtlsiPgLvb5AJq1+8BKm4LwTf8+b3Aok3Qcbni91j7/yG87QG8boa
gnYXxLpaa1vaeBekEObx4uyNmVzzhCVeJB4P0sUJgkd7NkcYgcenlEPePzQ4gcC2
1wLuo41K/iX5vq/Xl0mYNNtK6zPh+q9zVJRXzZKUDf3cinXubhjWl+o/9btgCbls
IgFCZjQHLP+cdEkGDL2m129SxE3biRCVh9I/k5GyQdinhuNg5DphCuwpxAe4tNRF
VkSi67PVPNTWFlLrd/8bHdVmv3LZmCekruopGKPj2xcHBO52n7h7X9D9ZPOxHtAc
kKzPEiEGpx0Vl9k67VWrue8v1KbB/yDqvhh3MHCw9M7TAnOPSHscIDPa3hwIUzBq
9xCEq2LuRT8jS67C0O297iH8Z4L/5uiYcnJ5ghIjANamldBmldbUlACNlPeobgE8
ReibFFvy8NJ9pZm1EKW08KvF0hp3brsbbjIlyfOk0Hto6N5DF3nW8UT79bOz8AAQ
m+l9SBsMG1Xy1uFqdZbkcCeGu1MyIcOhX++iZKITH8egJslsfxSce30+uY3JrjqB
aBQUkGP9Q39nhTMGknJmMqbG4s1rutJrGEqFucJRi1LOEUdN7f3IxpnnchBa5oUY
4XDtpCCj7ntKU6CZ/9e+1I8W1AxX5ewd2oFyu1n2OyIPjWMcHpqcEb285BxQjXBr
ZSqgUbwOWqoKMxNku4AmH4r9jkeD3f26jQ9IhvvQiRSg1/Xxg1lK/0o7ZzetIKxm
UAouNoqLeqPfE3vhq6qcQQIJCcfFOgukyarets7cK8y1RyCeOpmLZPf2drjRruG9
veqvJoUzOmbnX26CdWqxjDlxtLzPc0fbUxu5ylyBmBa7JQuGqg2mVb8Ql4Yzn63J
6TNAispZMOReYNmLE/7+hY2WTC610uCNUcNr4RT8nV6R37vvGa3ymNZn7Z5dYQid
+9FJ0IitcXv1ictO7I3wspYIsiLx6ArWr6Zid5/OCKOFY5JyK/5o0mKOoCcKzEap
id2CcJymnn3rJ9tV2OBldtnd10Or8g6CaROWOOSdJVjtMk2okZ1sy0nLX2B30Tl/
IQUv3ECHG4Z7rYBLyjzVtMETIVgD2thgC9XTOuH/4U8eD5Q01W0yqxJU7wwgwQqO
GVTZRQww958jfVL2Ci+9fwiaXngvKaJPoXs0MxT0TfUY3wHdDy800Yk8rAWDxcI7
wOn6QRg2WAvE0kniMR9xIjwVofnz/88H9u9Z1+CvhOHVYewpLDckurviuJLUTxWS
bt4CUkJyKni12heMd1m7Cl3vYoODSpUtTOLHU6sH2A0OwOTwrqUCtjtNWa6KijVb
1174DWEzJGpmRE7B9EMvMEx4xJyRirciBzOpQfqG9tIB3RB5Xpao7uLJxMpDxFPm
ipgBOJkzWCJ0+gVI6dcgDQeNJL85ZvvqinUQwqG9hREMXPHp+BwqfVd9Acg79cMy
S3U6guIKDw5hhFewzIyRs/115A5Q2RQ5ksH1vFSDIeXjtOHIROkoFFGv+M/9IJOU
GQqwhTg+OuZ3D3axiOKs0Az1MkmT/5N8iiFFxHjwmMgZG4bd0ZgcHrW7BOcX2vax
PeXg3ig3XwV0f+Q1nA7Ie6wZd93C8qjvJLrp2T1/Ta0poiz4KnUe6M6QmxgMHhnG
l1Yzkjr8K1zzGslFJMhEMG4d24ZosIDEhmkaMt33rMy2c7ST+RLcKx/k0NxUoMyX
hxcvdLYkdtCoZ8P28ArzYfHnYQp+XC1rYMxXZp988z5dECT5m3tN4tsA1srpCOiv
fJOhHl7j9x1pG23g0r9t6bBjjD3emVWsZZoljhMv0B5u2D4LIWXaEt5eO416emCw
7AylL5WROVaa9+6PXot591AIYzf028KBJIssYCqGewzvhpWN5olrSBcQ+1Nh9O8C
PDyxevghIrS9sqSvGBTHKm1u4e6lhP1leRT40xAg9rBDhcVSP3KHn3ybmGqbULFS
4FRFi4EmeuIHDHt8ZiqCfDBlQ/OdI8NqO2keXg/EKAKQnOSt6r/HGWRWAFrhhYsc
yKO3aFo/B7t5sHWroNAPIEgMipjBuksI/GZOhBYkyvizkE63Ds2FocZgR8to5ePW
y3Fae+/xeaUcftMuTXjyUvLqQQFyUHQxYfr1khYMgC8vUscqUSFFG1vuKfzT0Hzq
LThnsAdRu0zqHqU13f5m1K7lZ4menfiHNRgq6LjDBgmJnue32NFRrRS8zU1svu/t
yDc40/OSX97i4JhwWHEhuZ7P9YQ3S4RDBokE2NUN0UEc40Ps1i4a2H6m21pWhsc5
Pyvcr57Zglyy7tGJ+yMdR740zk/bWOH0omHXfPIgaFBIXfa3kwMUOuyAIpF0op9S
f2dPgxPxvhJWBciz8prcGKMIGw6Y2s83ricTdY786kgOPoPDBYuVj4S4GoaGcPxI
wTutRKWLP7JWuIcoYAy8GYSk4cfPGnXZX/+a3wc7OiZqK/ZRZ20j0BvRFVfv7SfA
SHl8dvLUrwwdeSQNov+Zg5r5i04KBdtmE184XqxZBG/On/DtSDI/hw7X9JBT1hXo
7ddxqaOy+oyt0eFL1fp1ZwwWEJlPXi1795qQsay1urjJen0OJxZEvZp4+yXlBBX2
dlkp+uuHR5+7fB3YGxcrJpDiYjfyPHQpjZUqigBV+iBJJ3NwSH7XKVEZ8k38N4XT
q6Ya7eeHz4r7SDKdCrOy3LAdnXiSpGtmMYoxZA3V8kAjDozpo7wv0WBl8FhlDOug
+HL/cAg5tlZpWt/dFG+wGKbO1PCZKxZd4ahbxjPYRWsG41/4/xt9wLHAY3egOLiY
tZsTg/wwBW1JaSNjX1YTueqPqSgOtLBMzdxrmQwmZp4CsmitVyHNI8kxpdYgJQ8l
JemTD93JpdqPih+uaxUI4QXFd8ymYt++nS2uKDkSdoS8mroLwUX6+4VMn1Xamywd
jTB2OM4cinzvEaly21+SMSTCYs4c57jIHQI9iVignKOAaUjIR0rThDstEBZEdkpB
J6PuiUUzdDjBLWLhtE3/p/5gO89F+17MIbtWwcft4c0ci8ps/no6SgJrUHqvkXQe
BU/p8DbP1UgGB0jp2hRzh/Bp6mf8Z0XB88B9AL5L3SnN2LSfwxSGbH+9NMDhlFUB
RGlzOeiHDgyjouwhacCzUF4eS2CIG5EcSOUBJJSglbS/HwhVx0Z6hFYIewCJoP85
Eh0uEyaYdyFFlgJaZZ1q3msvpn/MVR4NqPC5yiYc0CgkreA/0xcFwrgqD0m/KF2v
L/LghSjX+cmR4GpHpFITllldBPC4237+prUKgpZSVnChhNbwTBG9nhrVBeas8aHk
zOunftjbyK9UH2VvqfEul3Z+HMpyTJh5+db+Rk3Pz53JPXJVCIvA58iMV8QJ4Idx
Gp4mDK1ISDqzwAunsAkVmYZCTRegTDKLoQTy94oFpD7UKljVY3LTwt7OgXqeH38a
oD55NGTcztHFZRLE0BiaQrNjoxmlO9JkbQeFdf7mTlJCSEBkP4qPHt9drJlA+ezL
ye69X45sEH8vKW1TRMwWf3iA16upvjNKGlay2I2cUeKLdP45elGpbXFTtY/GgQXi
YZqGhNhnFkWVCL4hsUdi8tW2S7K7k1Q0/e2SWV2R+24SBW8MGRMdUklSooEM+rz2
9af937Nt0VUK+HNSdkXORramiEWAABs4T82TVdfENm8XKDOtzyyd9en2VAwjRzlw
qC4+Eh7mhR1a+9iybBJAp5tN6XVFLCUBNcjjgsx57xODT6Oh272K9/K8xGW2SlR0
LZ3bQeAvZF3+gc+U7xJR44hN/MKfJyjTfGtw5cWGBrtvvUWF6WBn5pnbalDJ61V1
Txh45bwZnF8/duqDdtn9J+RhC3MsS42ZOPk1QX4W0/m2pSA3fTtaLtNTQ6HvpAQH
xbHZg+MRfDN7PDKKtc9355MqGyRRGuiXIRZCa9lECJcVvGU9Jh/3nr+7COckAXPo
OwuWVwlc5AvB1E7f7x0NWXOVKWAPbHV0uywq//7lzgjLVTtMZCTi7QrhjU/vJtVu
VeHsjWRDM37PLAhPe77zgPrZkcSY0E6hDROKRvRXkHg1kuMhGX7bnokKSFgPNQmC
yDHdSZie+weToAkIoADZ0BP9Wfm8UcbDcwCNXsCDk9can6E5h0ADr1wksiZ0/bq8
OXbVtd4PFrI/CnLNthPM8+Arlf6IBaRzbNswSBTB00TYnNhH13p6NST3XRpurx/U
Iq7XDVg3NifYYZa1Zk4e5+CO3UCIUFVfrXQZGsoueqcYh7I6HyYtKY3Au2imMH42
PkgxK7dPJqshx7R4T79rXPEbj8poot54AenCIV3tzC4bWzdkt6/gUj7QZfSUE6rt
bJhLfxk2hVaKfEgQqEELuV+3w6sDI59Xi2PeEcT0n3XKaxRN2g6bPfwQNxNcH4rc
XiZK8qVgEVn80tdakAakINzGW2VmVa+XAlhx3hMe175AZmWuHEdf9hx3+a575CvG
M7PKsPemGeM+OXc/qeElc1XIzQ5gfLpaNdAKOlgqjXF3vWq+rbWhs4ef7LBmKlnZ
yataVv1nv7vv9obdDofEoHHrM7zI+9ceAVro/HI6MLT//hMb9PJ6L6MO+h7I31qA
cB6MFZUNbtA4pEqMOnLQcXISULeu0wgifxQYI5KVxCs88zoZcYZJJawnBSujQoLx
NJ+4jGADtHfkVyjbKq+e1M+DPSWXzcu174WyYdzOItYjPYE37upmo9WywsKv1Zqn
RUMTv2l4uPKoj4KczbS7LEbEp4uPF6y7cjo9QCPLfST6N0xMig4OXaTzrZPNAqIM
0nnY/kKxJVtDbZ85ccMwht/NQBB+BcMeOrzHDptnBplNOBUu49TdvMLjPVJ8zLp9
fRoyBkHjLs1sZteZIDIWxjoPIO6+8/cs9TpWQ/NANlq9kxuEA2bDpx/0kA3kXQ8F
j3MD1YaFGNKraMgrVU0A/BlWVQf7IfylaX4wAcl2nLMegQB+sYmRKAQJhiUgUQfW
KZqbxzq4DftTjBT+i1rCgT6M80pDfdRU9WoJN8aDa32kvcwtNarg4oF91sEMIB8C
CnJrUOep+0w6FOa1C5h/Hez1r7uVoA9mVwQ6/p94Sip0iiXXTQ3QTUTyF+CuDcMr
8NQ2gvfYsm23An5+UEcHTwXq93fWOoP+EjssuqfCafFeDD/VSkkV4c17+fQE8eEr
l9Xzi6I6FwYo0r5pUT3ga1ubFO0jrtpm1/L9XFhuKd9OxvOS1dR4LUibGlvMMrdR
gjo3UQTx9H+glmjRoJDEqgR0Lb1osQRtuKrBxAgK4zMQzDH8Rg/CII9MPOhtjxsc
covROsXClhOoLUTzDC8j1XOub+AqLYVpdcJUhT4ldgXyJDaD2zzJNogscVsD0G/b
OoD9JiOn3iy1/ft+KThWxCUYbNReGDprOoYtw0/54r0RCoTq3XMX5v24cv/YtrhG
IVjHqdvf4VVo4ESib7bvcjUvmqRdw8t5hnpA9m4vYvLm/PwahOhFNn8eTeGoeoBU
5f2A97d3gL61ov38v3oFRoAeA9nHGorBirZe53oYAQuBBz3FFW4bYde/b/qOHP5z
J9E7HmjhDgNsV0JIjpSnnHDPW+IpE0+Gwxf9Ok0VnlZ9sxd8hN64VjX5IygDxkJp
62ppgk5w/IpQ9/1/avF8Gn50tYG7M4fltqkPkzcuxir+v/lNH/W3tiuUPdoMSkPD
FYBzVExmaBOHNPUHJKiS8hXIMZZmtu8zTecsKxvNuEXaJ9zp6ojkDEFdx5ehT+T7
tPBdCtPAg1FhTmSUKaq2zzqhx/Y6+SFRnPSYhDbKnQtydtkw1vjdGMQ5WGI0KuEg
Vpmg3Y/ofGlqvT8/F4Kbx60ekzN1oEA77mQvO45wp2Gaa8vMLObWruUDWXKwOo9O
DGFxHTj4WhWSxS6/Zj6VLRr5pSNkB1EEOngRb5zyD3izVQL3Ld7RcXYK5hsMEyHb
S6fd/xLXAD6z+pxBmHD4XVL+Vd4xZlrYCPFMD6rUFClYIIimY5NRGuNVFriybfUX
ZuuZxVyO1VE+VY8CHC6EfMg1hAbyxXYOkM07l3t9b1MBvvXKIBK1M0wovoCoxgrQ
qLUIFrie2Ke6ILuY/PUYGBH53pJZ5DfqWiExxxWTpCMxb8MQFjhFsUwNNiG49WZ+
FxiI9DcPg3vIVQ4AkvSW58T1VHTvzoIj58dpakjeiSRdu1axu186PObO2CTdEBpu
27+DLMb6SLwVpUDhKDKhMauUlIfz2hrqbMnhPXcNS5tlRYy2tytRpavHDsBJldUc
BK/QF+8BxVuIkFX6tzrKrInRpCfv0VMcLTnIReE+aRWNPGYmZqafIGJg1YUzWWJE
ntOkqiHYjRaDMlJEkn9BpWuXuLUuEjZE9PpcUGpAJd5MUbq5bQgJ6PT8qx3W4uIj
FExkZQcsfajQfiKT8YM1KvGIWel2sfctqPrAUT9RnHubKLLilcA0PZFKBvBY2bjb
CPtRysnCVBlv5TeqTYNNb3jSr8QejeF3B/uygcYTAR6WFHXowVeZaAfK8SOTRSfL
SxikdRBTskHRu7slgfNP3GcdDRq54N5gnLyYM3xOWVVbXnBLDQG34xyJ3RQyMsHo
C5xiJ3C/9Ds9HGMVFqWYpnpfJj0TJdJlcmvjz6AH1bAXyCKvnIzBbva5QYM2n7oq
3OUkV6HvgANWcpFaVhx7Eqsr7xadXYDumzSgtAVxyyPgipxUEkSYIBAFKVxpQARC
Lgz+XHxKw7xp+XLoSrhVd0hgS7t3ZWoX8z2NL3FV9AsTnDFVOaQpCIjAjyFT0KI9
Zt9LgE2+ZsKrnsQtvR3GG/mDD54EXmRMBe2u4WN1vSUdg4fen90FcuDYvihKNYde
MXvUS5ib8y/rnjBgLOMJ7hQIZaWXz6Rz8w5C7EA1ykaAe/7aOPaV6QDk4aylaiJL
3Q9Eas8Qc1F1qrFj2fhBXlsuiW0GWhTbHuTwdNtwaBi0G3K4GHp7oeIbiUPbkt3T
yBFBy/4+5E5UFsm+72dQRWDL8+oPYpBHkt2fvvKWud2D7ffiqg3cGgAdEQRc/kEj
tEJCVWwY5Fwtvh3AkNSN6+bxxACZ5l9n9DH1zc+g7fBox02u3Igf9ySnM/Nt8lWW
alWiHqE0GXWmrRWjXzKbFKeuhp1XWNX6NBJ0vk0bGFOZ/St32ESbVmoeZYkpGYzJ
a7sCULLk5URL62USWHcwLhp1xtqO6chRBgMCjLTDc60FJDp7wQ2FiLMAfqb8+sUT
9O00UrlRKh4d1EuJoJP76bJLguA6qszM6t1PharrRIDk7IcexigNmQ+3BLk6C3h2
ywdJ0N77gmN0+Jq8MxqNZUWN2wCRuTTUxMlKFmv/y9ypAOCLSEz18reQu0rSjfqq
xVJgZMeT1kVmzufNotNLmTtqTvDPYW9xHSNKEmbP//HB9WBLxIYR0xaNXAclPVEP
53Rx7Yu2ELFGPwPoDheU6BQHbOtWswuwfmBvqL98L2dT/ZMgWLq196/5L0OTmSbV
GlCP4JTxpcDZDAGgnDojGAdw0xJH67u4LupnA9JlQpv172+fVUaor0MVsbAXPgFv
mPKr2esbHuL2+R2+KJeBm5Cz0Y51st9p+YusFcwfNqSiOAMF2lTpOPmd6F/WohIb
jOVBT1R2eylcXQG154Jj8TihS8IPkIKkUfVZwbcofXH8ZSD4Wj0wP0CcrjadR/xc
pcOIdC3cnssXv31XTtfJDqU222eGlgYdhwtHcahzNhzS1aNmMYj0fijXFqOXpJRo
jZrlPhjChHvSOm+B3CXNzl9rcWDiQUymuKVbeLAla1vfCT+OLRbPvMxlsCRQiwFx
FgreiTwedVClaP4MNJx2AG30V79e+WTwqISjjLzgmj+3/bCQoPuXWQnGQbhFu/ez
LQ3mxQk9u8ZRcOb3f8viJxQ5DOhlmMiYnGKn73BJMTxwzvwzWIeCL8d+rShr7vE0
UK9/7H//uAXLvOn6Ro4fqZy8vdsb2dVfJ/S3yf8NKHeLGjS0ihZlnXLxI5/X/Zc/
gWLDVyHu4lLI6NIkOWAxKTFwXwnyEvH5MhfgMo3vm8Mesx45lf+i3kruczG/Yzyp
56pEpmpMlInrz7icC82wnyX4/vq8jTvcL9hu0zxMHbGcq6ASOZCoQrHAqK7V3xim
Xqzh7NclFGGMUzSqAoJ6uwfVe6m+thscJUIBl4jFYYKs5K5K2dbTePWJJFqb0b02
VheaZ8EEwz71jKmnTlb1MVzWcT5PkgSTPRDHez55BNChCWFYoYm7wFnNB+sMsScj
ip5AMZXOlgGfOpgFbHYsjxu/0rb2iX0KTZuK+BTsczK+NG6k1Ze+4tSgwNE2WsN/
tg7cKEtAU0R84iyod+45/Lj03Pr6KFRXMUnOBiPLu9sfHO1Gwt2izbgBVX0gyLhH
5UJlsPQem2ykiK4i8KRu2quRM6EqqJyyxD4uXfKSi2VhGuUvURPFQX926nqU/ngM
yPxag/adm6NWNfdJVGiKnKHxZ2+t5TeAqATZ2ltjJfbPKvS9MVC2NRF/CRbDa1Ix
3XS8eKrgWU+7uw7F+aamfg7MO2piAgkQXrpS4rP1hDV4t+UbPNKPPtlJkYpnknMA
eYAAcbX29TXazZLsSruOVjTcLVQ36QWGetxItasOaHZewa7wp+NOZKK090qN8edO
sNN4oCbEZQ7VOrGCKWWrnk81eqgNUJyh2KdXTaoTf5ZpQAJnAzVwKljgNVfQQIzb
lwJvcvLj3dWcxVbBLZSugbrw5/tMlKsQrHVSfIqeDTdx5+p2F/w9A0zRw67o5VPa
8dnEc1Cg7XWwrKroT+FJjOzaQYBs6klKnVlEQ5C9wWI30V3N702bN3S9Z3+X4lL3
O+gqWvPbvTKbzbvV3OV0PWOPonY7DIYbJil/yNVn1j8affbsWcLIoMwaaih54+X7
9pr0yZEDgNYyO9gu90XyjhmgXZsMPqSre+Zgeo9C3PjuKQgvMy+srBGUcHFzgI4k
xpz1gq8eADZkyEOiui2nmS8rOjpVjFY/BdcjX76CSovi4Fuq9Ame3rGK0gLekkiA
vnMdcKFeJqBtNkGGqEUby2u2VaR2xvBaXp4WL6IFRVz6nTcK/0xNv62ko3lP8hr3
13gXQ5/cz3IkEn5fBdWo1JgfN3yT5OeM/TbMGOB6XmmVfPWF7BgycdnhX2dZurLR
mwTa1VtLlTor5/roqVYq0DDX71UqlG8EfDrst4L/es1vaknwBgT/VdFLBpRErxay
9HqoZIo/mao5/Hia9DczgS36lYS0o7/ixGTlwrM2oXHrFvZJoMKptGKXaVPM2oRl
x4W78wdRPUoYfqfM7Wn9nIERxudWJIqaWuwchoJq2+K1/xVw+6gatafccqlFQSLS
79egYQTngvuj/BEWi/cPQOZETLAzxWKMG5lWjtWSkTJ+HY5OZ8PYxGRF4Z1kHC4T
dWPcor9yKjBnRdSm0vFoj5nbReRDBjta4q4H9Ch0Zv8vdd7DD3CNfQo7F6TWQ+if
y3whd+MYEhzAfG4MwVqVcIh1qXrqKo8a8GGof3bOhQgllIpc6yK44Eg0GfSMQtm4
AbHKSGJgCJ1dBWbaYIfu//xWYDS53EoYlMKwrrPty1ll87qBr+cBa9PPNy9IP3ZE
nW2YsvHpWAauqQ8HnfGRdF8hzWQxZ3WVGO/4U09VM5ZZVkojKkk1cUgCCu7hnHim
oIsPPOqdjznVs+ClXmisgp4yQYROfpGS+N1a7B2c0bJjSEam3x6HO/tuZrA7d20M
sTkHF3FuksQq0h9AtAkxKb2OU+2IZw1HFpZsAvZmXw02zjMMp6n5Yyh463KHQ6c6
MxArg3CiYFl8FnJLhB+JsVR1SYhOj/oln9sPdWSnTzTaplulXqHT83LLwb0e9iri
mvvhNM/CKRJp9+G2DHIBoHMg7lhFHnmE0P7ogwpLyAHp3DacTq9/4+FxKvYitncl
Ji986nAGiiQzetNj2QnqaJJrgEhMUa6RM82umJ3Y9WLQA1bN27FpQinYiSu2u/U5
CpkvZAsiHdpDYsfdfPx0j7z6PYu9n1yHC2fr/esHmfOXYIaO/H3zoHd2Vxh861F+
mkpvVynUaDUrNkSSaOfDhgYYQ3zqr5chFLulBsdyi/ERmqa23FWOdP28yPWsHjhO
JeT4R8oSrJeNOs+IbpO1NFCOiYwRFsoCS0hL58MJu93zhaIzIkvt+IncFgKWFfJe
Jlrh4FZ1RMTKJ7GhzuTVd2Gly3niP+x8vVVvtaCpSXkl9OTtYrUQQaJ1JySPU1PM
JO4Me/uw4iIAu+QkTpSoSImi/I8U1HuGqfFhKOBJTrLmoYXCBYmJ14/GiFhXvSV/
+aliA+PNMgqP5EIhGw6gBPPxzCDnEiwv8D1TzPuHda22ws2ca1BlnhxZhNpsr5ni
6QJrQHpxNDZUjew/QxQKPA55BA6I2NSjJGRXkpFJsS9/8yTqG+g9G34tB/Zxs+b1
zFZ/tbwpX+XbiSdoytzEHHgC/XnRiUlVfCGI+oJaX2HVyVEimgSpdnFp0mzCjEIB
m7ZSPHTa+r42ugCMRnhGT0s/F/yoRafbsLHdz+qJV+XA/WC5u4m9EHRwiVmX/l7C
pVb7wAY/mOPMUady67bXkg7l35WUUc4Eil5jldDuyfEuQ3IbnnmtY4dlRNfhwM1q
c99QvzrTTaskLr96Y9rIV4gEA14BLjteKcjK5iQ6FBQUtXMAXuKoa0WGFMMuW8At
4pmQrWRk6OfSihFSNMCh0/gOCAQs1ZLtO0aTBbzLNP3cNiCNPzI9ifpsEY6aBxc4
14TeSVMuXQ7bp6NOJjcFHjLbJxiLGqj6ipiMyCJx7J1FODCgsse1hB+bFlc7+ltD
igkSLraL3b5nB45myDQ+LD0IyIF6GjayVkPN39BhejwjeCUP/8rYJiLUNaHWWFOI
drvWPY/ar2GBZydZvNFV8YjYFBktDA/fDmtKt/Aqp4Zk1EgJmUMbMpT4esz4KH55
RjfnP4XKfr0eCJwJaSmZQ3pSqb55ZuLMFmS3leoOcSCQaE6vb7snolmmhlIuIIKP
zrkvyWa+6NSb5Gemo4JM+B97nlz/pMNA5H0dQjIkZ4A5Czmr1b+Jj54zw6Fl+DUC
cR+u6gm5Dhr30ygblud3Vxs52snhyOIme5tIuf2K5ECdpNwGkIMZ+KZOVJ9QWHKh
RcZ2sIXukfzPjCoyUK4PKCQz+pCKukoyPdN8lTl2wZNk7PcjE93WL6cjlMeg9VAl
W2xyqVG4BPD6VjNMX87V3tU2OFBAQE8h3fnZNs3iqYE7ony7W/HmkLRlUtVOclbd
yGFjvokRFnTlVf4Q8wfHcwE5oeEE07u6I4eyBSpzIfmf8BeR2CSlhoQybmNqwn2Y
Utx9IF5KuJHy6P1Fyr8xEeQuo0P3yVHkvFWkkT7qxPmJzHVwy+8v5qUnUQmOkq5t
iuqoStcZUJM3RAeyiCxui2cz7b5g9oCxFuFByWW8UA4mkyVJamMx5yPdFtJ0+1VV
IUmkbjE/ze4YJJ4yP0FjHt5H/M55KOq5mOVRfkILtBBkBon0f2HndYZ0FbIjnZYc
FThl4r+vJt5FE82d/SoqKicoRhuH80QHCu0pxhSoZvRTsu4WxRcD38wAsfDXg9E8
OBGBA6R/EwH6C8pCEuSSRB6G/1UWqaRloo9tj7rCGHQLJc8kLL0ae0DXzaf9SarS
wL6nMGo0JKulRb+nZxwt8PsiQ9RVuzwAFoW15JqA5haFmoQJyrcD/VHKD56B39NH
rOSSP4POB6GGILtkLfSuud3uWttj/fmHY3f9wOz28e1zqhxPOH3/SCNe/tU5VsDk
wzU/z51cqa60rYAYaLtPBTp6JYdOaA8wJKgactogTaDNcMCNhwwV4yzjtzwaIy1i
vtbiF6t9GCLLcQl58H3JT5XANF1hNY4SE9e0zpicZgbKAKz3pF1CzThdK7LnICb9
ZefBhttP9LLnvr+sk4M2s8fHofMlUE2EkHkgfPtgQFr06aB3LAzOp8USGgksLLOF
Cusm6aUo6Hc71OOc8jhJvGu+t6TrZvM3350YBYTVlVgEREUxhJa4Nz50uZYFIeDu
Thjid6fNjfiEpgjkZ1HoJe0+x8OWVRabuBtIdY705q8aopFYpjM/DcXsvdpSf6OU
NKrpScSkyAvXcp05HUiB+hRAkcMOZwkYFW2tPe5AERodLybxc3977HnzNsSO4GXX
2uWOiyo7ElsgImK9yTF4fctzbAgHps3/gIKRNTwBJMqcrRqjer8dO+5J1saoeRSa
yGkRM1PCMUSEWG8E2VSEW9EYMHxIZ/FiBYyJemy0XRFyJM6l7ZKtAWtilGJoJZlb
f7ikFUF6ai1M8iCKUk1qogjxVBi1+UK89yk8KPZ4GrkGsbli9e827OdvDjfsqfT5
yCdBYOys0FYhzaYM7iuB+mEq0D1ApkWR5Xrk9CsQNGhDZq//i2DMgTRRuyjP573x
PzmctZnMHBT6N974HLbnSH1PK15uQOlC5OPIyTYBTCEu1fkj/Gk2JvKIUox6+HPR
MKt2rAA+Sx+ePHThNR4TYcNLYR484JZHYEyC9EpIBWBihCrHSfahRLimV0AzVkLW
f5idB/5RLSE8ef5sK7Y58zGXEKHSKPQt+eLMdE/4rOdQ2ycxg2Iw0DBqJe3ym93t
GWaMTWJtfXWgJ/WBT9MTfzixxruApYcfj8FdFlTU+wmDwEAosJLdROj+To1FtJNe
u21v2ovMap/3L7CtVGYtm+kdOLz/kuN2K58ad2Th6EA4OavSzDgS0MLWOlKxcTGq
hdaMaXpTx/xS3FWsbmi8jndWD1+8p/aiUJFzu2cJa8rTFgDxDzJCKwwm3TvuWS0L
Gh+CRdk5hgX4sWgkxViOt5Eo6hzegZH3fe1/3sqhFBSPFtVCx9V9yPPMeSk5dM20
dOgvvec/StNkHrjWMopUkIP17uuFkZ3IAIQoWKfDWF7vP0tIHxEH+I6uHgYKiWKU
tPgHT/ixqn0ecC8sajHg/C77k1IYOjRYZTxa/LID/2uVJm5HtUFdGLxtCrw+IZ0t
mXPV0IhimacQIkKHPQhsa1fTA/bCyKTjatb/hL/kT26HmniSVoYgzBazLFOHMvuH
LhueL1QsV7DmzebiHgaqBHaY5bChF4pwVMiDIh0sz/3oL1UAyrREIoOXg8Qi8Ih8
AY7UU6s/sYdTb1NGk8lHk/fafNOfeW3eGJe6yyY/41GsWWvKLAdIzlV6uuVWhMlJ
Ckg+bmDyXN1+6qpxZsispSGVPag70qvJ7ikBsd0k9dTsQQ/QzFwvTHjTyF9jNosS
UYoBaRfrQFRGBTykIXkDRHRkNVjWZVUXngErotpgLMRiwMdu/p+xvNemYg5eHF/6
Egu1YrxKiSosU0zgoLTMayENV2O5Lp6yZlD1u6U//DS5nsSZQLRoOuMLtgk1IWMJ
CXNlw/dt1N9sXIHtmTkHe2vDCv+YNWv/Ez0uWjUCUCXjTie7GzThkUeIpnEUlksq
xoZ7uJsDmX5wRRI8TTxZXpknw/ovkpPf2iB/OuoQnQQk69uuaYJeap/82VU6OqHp
q0rbrQG5g4ung4eCS0dOMpkbKCK08dj2yhP1Q3GdUpDnaA9DAUIyhKZRKfTUiw5l
MX7ULoklI+/W0caR0l/GvP0/C/wY6Grrnp5Ykm4QVnEAKcBTzvg1hNGROwaI8mhq
6Rgnl5OMBgBIqePOGu9EDaM+joHHGw4PKMcE+UXNf2EXlb2PZNZUD6NKtGkRNs/5
xfQO+JlbhUH6v61KkgOXp5ndZrOwvabtVHhWvqJEZrkrY88oQ0siYhsvT2MmwJpT
61kIinUop0fgRl2PLpjpibFiqlmpZ3dnLeyjdB9kjegeK15h/LP/XRrNO2SaZBg/
jJlHBVRCqDfJI9MxVoioAdhmrKn33vwA7fhFNzXqpN7Eb1R+L3+PUI4bN3xCsnlW
ShPla9rlrdK0Dx1fxS9jNGCTs1MzrNV8p9+GD7WfO+9J4nsUt4G9Ubtk5ehpoi7j
hX3G2/2jfDjeK2cMn3TnvrCA4lo1PxKGUEDQ3dSJi5RN3+7exD899fueclQeN2QY
sir4IwKyOsnOsq+WtWZ5YzvaGDwxdE0tlIs/wSpf5+OrqfccxhCurW697z41DFNt
Lnbe+Y2F5yI5t4qljlBLO+kLTCuraqJQ4DlwxCLflRAqGZ+lSYN4KpebXNvCwgwm
ISNm8HhCNeB7eUE/8BOnVVReg8chw5VW2liKZj6nM+bIwTy+bCX+iaKQZ0+EB+7O
yvnnqIprmkQJBQNfEQ16ONZOrkXeK5j2F6LpgpC6d1kaZphV5cZNpvkfdBYyZDpG
8HfUSRII0vsTMhb1PYenp3heDXeYp32NIMW8CFob8j51/oxu7Rf6Mt7/3LAMEw4e
FN6zOUeKlQss4FCor9gZEtplwsdjTStVUGxV0x/+TcLksGttKg2ms/LxAqqiHCUy
A4In1hhySf3HOphbgVwXCAPyh+mYpMM1buuJDvzgjmhgN6R9TKY4v6O5Sjji9PE1
GdfydtTcVVbX5gmc1guuFD5WVJgiBGiXinMpDMHg1GeYbfqhxQsTxzaAxlXL5MjM
9W6hnC1oqNPRWDLjE9kepdeXMMpjTJLGfnKbrbRSCy/ydA5f+a5nnwyX+h6wZkgo
raC52bSSB1Sev6Fqj/H04E+LvB+rmon/4tCqQ3L4QdWMRjwLVabvknBQZv/UmOeU
6OOTMQojrzUsBmei6nfxk2sym06mFDqMeXypqKrxp4rYHzp/Onp0yrp+dJyup7Z2
9ogQi+Q1cQ82hxuf4w+JL4ygTc0rXvwKDuQRwQATWfcxe5f11bi/KmCwKUeEvyWg
MQOqM+qsJCL9IFMYD+HjSkj4BuZho8IyOiLfRvvj0t9o9p08zNZN1a6JBw+ZvMcM
stl3Z0l8ZXxZfVbdWsuiwWCQDnMf2xX47X+vEV6C1YHwZW3Wu3CSlMVF51y89ccI
YAMy9/hdqEJp1map9S6ajmCW5SCRRczPEgxFJnZj2YSksKFExpQtWVbs8+BQfqbL
DItwilqriASPp7mWV2mNPMt8CjWTDfHEUPQ8lheMssTW/JkWtiVZDbXi+Ywuk4ig
HaOB5XKt7kvkM9AdkG4Yq8rVDK7nQX0Qnwy4blmTPLUs+AaZM6zwcYwaGqjTwJ9N
wt99/iWiGAlWZYpAgVrcRFQCz7sZFZWUYfsYWIlonLJSeEYzlq5IZS+Po3yIkX2n
TxhR0+2aplFLQyb3nqe0YEGmM3xiQ1kQtP4ENeVZ8dCdeMeqeKk2UMuEWCK1VBmq
IzVb5TZgkVVmCGhJxgkMi2taAM0nXyVneXLJq/rUP+ZR9oBxoII+ahXaDhPpzhxe
rhA/LeRw9DtVrw24QvwI2hEugT6PO4sa5w3sawgr1uNWleem6srwce0cCCBIt+xQ
Uq0J4GcAw2QYMqO0AoKAl8KCQbesYQAySasLWj9Drok6GZrm1SpDs2T6hEOoj/QW
uC7aa4+OxDPi21vP75/JXcdGiYdnhx7jvfFQPaxhU+MBkSn5C7Ou0Xz0FVA/v2Us
gh+U6ST5w7LrKI9Z41kRXWdz62cW63T/oL7KyxRDl9jE0Juzyapou/iylZzBpqtS
y7CXorH2fgGxBM0K1Q/PJ98yi1qtpEAHgdoozTUxjn7uFgtvkgx4MeN9OuvWhaix
ZozSMcwtTrK0tCSgkjDo/DAa7zWlZq+9GSfR49imuosRdzQFDjzuzqheEiwoeJzw
r5lBn8rBXN2oQa8+hAKIqEVnFwgJXcURyM1wvIeL2GspF+mOomW+v+DvnkFDDo4l
4tStWySUz9QFxxR9L0nFYgqBZEtSZFFEwFFRjL7GrdHgeiFbN93X1XoGppdV4unx
lZkiC3m/FCtoSGG2TNzWlABZi5esTA3Pd0LznQ7uECbzuAlsLHw5Ilb8JR458Hwu
YS2/+WzTOjG1Xh5AF3b++MXJd0p1b4LANf72UCaJ7FPS4n1gp7k//vBJvrJp7YQi
NJ7qSX7Z+1bOo8OQsR18E0qFtbQr0m9ZLCBMitzuddunLwpz2kb7fz9jYpgf2ruG
zO3e2i1AZ23ym+cSQi4cnNyC0UvGwDo/cSgmIkoJdFfeQKOOeBjOq8sHsML4lklx
idNRoeZIVJ/SFu0esF9wlmkaqp3tSB+PUjS0E2BYTI72Q3V/aRPtz4TQk7MVcrLP
OoDrSvx/8RszVs1TJDtogpGiBboDj5bfO6h8OfDDSahCXWouFKPbtDztn0Nl0ylK
FnGx0Ba58V8kEJHvD8rn2rBJAEz6548DxCAXRj9ZcQxktztFU00Vc2aA+y7z3gb5
LyWDuEHtwwAEFEWxCrWn6Dagp7VtQOgA+VuqkE3IsK9ZoGGF7xFLG6gbqWV3GFxF
GOmb3Lhabnfrh3eKTFcqual6nmR5gJ2V9nnW0TLI3vHiYgUHLzwgGNwyLh2ToKpU
tvI5eGgn3127clNakHx9xe9N3pZ8UmCVfHGqFEEqCjKhWZhTwsXdn4JSWNiEH6TG
0EGp/EEn1NTrqXgO5+jT8binVRf8O3Y/2KZAaIsiMRtk4L8REU39xOjETxhS+Ge0
B9iq+4bZjKVBqKT5YrFKO6UeJ/FC4tmSCJJpUXtEPQ1rXhYqxpG1DEx0oJaAs5A6
qwRlnjPHr3PO8bEnLRiAJGF5/zSVuONM1J4bJFgivEStYo4P8QcmM0IdbGMlIIft
FmaWV/+hDwAQUDEqTw4w1wJXkVTqQiavvAmaKxsPPBBdmpquuY1YxscjGPSDugux
kyCjEl0O15MwWSDk9199W+1OSsmSs0j87bXfPEVKLSHelZ1hyVagIipdl+W/wSsf
37cEBWZsI8RdDh2otjoxQ1Tes7GbyWct2+lyjsuRpYOLNLLUebcz6sNbF3z82F4T
vj1M1Nl6JVMsCc3mSS/vRaoCLEoVuMzR4/yhwQspMRB4mDr82VBBBVJyuj4RFvk+
qEwJXwzs70HacPDt+3+CSYwCttD3HeLjh01qfvq5s5CugY+XHr/unNtajqVYaGIQ
9Rbsy6d3rGgwR1o/0NK20RdNpQ6uPl4aANtPRfDn+OmvzZI4D+BWG3x+QU44QSfZ
TUPrmfM+IievPW8V632IxTrult4Qy0w973niactdb9/ZLm0nU9oLM9pzh5db9agI
0gwoQMpeeraQr/uDNxi2DXqG0Cu1wZy+TbdVOlgDLZsncOHkbOTRk2BNK0+1SKn4
HAyoq2bjHw47GNO/NcDIhhg6XVjnZqrfOhupBHoGp+h3NZrUNBE9XpnBn0JtNr3E
Aeq8KsEEWwKBHX6xnef++JMdGJBrBXn+faKvsFM7AMOp7SOpClIpHS3tB4qR93Xe
86p3y+2sODfoYpgW9CywiNk6tBNrgb99/Qo1R1DUH91wlg95fWZEE4OzscJqbOpL
oN0ydrzn4J184bjQNb0384ZSzKYzvQ1Y4IS8UTGhwynUFmioRqiT/yHQYRF/aTt/
kkMLI5d+yYHxbT7DHXp9CLaISp6tGH4UVE2LMAqg5MlC8WZiuxcI9VTd3+FpllH/
LEwM/1cSS439eYl0Jfq4nbpRUTupaua5eMq3f+EXs1/Z5JLLFXrPwFcs9ZF3cQXZ
fYKMR9/sV0gSZCiWLPOuwY7XbeyvFKOw9zqAqOQ+2E8GW002jdWG4pZrlzkxEzzD
cUUhBkb/82pDNVARtZnDutdFKBqfxV+4QhP/08qvUuNdCB+Bvmjgj/60L1XDpXa1
tFlD536dHk4NRnO54pz8tHRqgYIAuUHgPgLaYuaGX81s+ls4aQ7puRAeZdM6gNiU
9ZMpmBhBXfZ3kSaW/632L0ABidALSYOVLBKRfDPNL6bN1qEFMC7dXm4SshlVXD/3
aOzD8gDS3mtuO6a9f7sy9IPFQesfYG+3EMUCWDCO1dohaUhS9fPRexiaM1X7iEyw
jXxq4up4CsASIbBM5KxvyxTMFaEjAjWUlOXl9WbEqQM9FcO0URk3ukYAQnoY/noI
k4U6D14evzUCLPRhFB3/YXZj+efF0QAGe/VPzn/V5PgVodOFxOI24L1H2ARmBeBf
KkwvfZVVC3ntzElI0VsrH4p77qTjaizmEzJSa12TaRxb0flE17l3brPqiGMNXaQC
ywO7N3oUEzsfr/OXtr9MQEdF/dmgmAkJnhWSDRE/LGI7XsGs29m/dXiAaFUas8AN
d1BYC5xX1yvMMiIyafQshiCJ0kq9SbDXNQ4evJnCImUqTRkh6S2cMh4aEphNli97
Ny1R9kwiRMfP14i+/nv+cIUEhsJy/UMRVdtYJ6/+7oy+WL5IJgV93+cKS2Di1Yyh
oXg3IitKWiBjxgbBorW5HKfPPMzUBtNOWXJ0MHFSowJZNOjkg1wzit3MbQzIsUZd
/MIzL3aQcDuM1WWkwe3PgzvY/q78SLL62Z/SP7AoXNNoof9i6P2oZBF5XjVj4if9
5m0cFBJl6xjsZvsJ0eSiXLzCplKEbp3sliQR9jO26lmlt7lwDa6x9YoO6RpN0+pt
XmXhRRvEf+Hw/g40kzceuccQd7Yd7lQLT+S+471YKP2hsPirZqTAM8E0/YatvyUX
2Y3mUdl+IvoBhsmxpPbBdvD5To3yGiGyjXpPO+FSBzIe5UHcP6+eY6GHmIr8ZMMz
Aw0idoMG3fP0x9MwA/gA8BMnEVJmGaet7TExxLcCy81aY6gzZoo97FEnUdWWjUEP
+4aTvR9PpVgvCvhwVKJC+D1WsmMkDpVOfhbMTS6HN+zHj1040AkRHAI+y1SacVfR
VoLlIaWXSYhRwSHxTeHeuI0BdX59d44no28BM3pRfuXu7DELqhzQs1nJtJoGv1sV
Pa0/H3IUd+eGkLoSInDaq21tDFA4YMoWQZcww/+H61ZZoFdG+t3Q2kWiQJmfp4ym
x3hT1I7dI1wumUB/mCucfh76a+oKc6UIPjaMJ1LfNx2WerRoFN79lI1EOQjCv/WN
3wxCplDip5TD2Nz+tlHRb57AUmk/PBMRUSJ67i9gi/vKl8QfvNb4FQEBghff2oIL
SVis9tR7QTA1Dl04lqM6k/2flNLqy104yB6gdNjPPPywNLXyy0ujoJz2bPoKV28w
EvTQKGnX1+j/wwghHNqyeQbjlIlpFTk6fAkLMOyCEniCJjItbzrZ3Bq0QWfVhhy2
DDk5GkJ8/tA2on04oF3d62S4jjhQ4nBuu60BFejwm/wmAYT2JnMoWQHtRfbZ9W6G
eE5U6arc9oSC1n4aSlcNJj3fXxBZ8Q2qERCpcENf8uUG4v7pVfZWlNSwabiZ2Ih6
R69RqME38KuIFLC0j0Y7IvG3eBTsCIbRlh7K1JwzfLU+WHaSKD+s8T096Q3di9fp
ukBBoZoRS7F7A6XedWyOP13Vn2XnTfpboXmhU/yG1VNdLO67qxQbfmnFLGjjcAqg
ECAj9Cf2SZL4fczjLhSfiiTx8m7LiBir4+WurE+wububmiTkh1d8HZgwNIntVc4Y
7wlE0c4NGa1hPSbkfWcZZ2O2PKaEPgBNqKi3DedPh8Bdzvk6lWKYVaDUAl3DCHp1
LDJch/rSCIckBwRlcgzToY5G2VUgOlu3mrQBQvwsw0oK7mZj3yN9W4NkrdRjP9Rw
0keCtL9pwfz7uV5MSaSG80t5VupyMIhh59yKeLShvAKc8TuBEpUJikBAZuHWviCA
1GDf9Zv56g8Fk3LhczKZYclmm7HxIpyBExpLjgU3dj6bATfvTLzoJN8z8d/i9AHE
DS08qVVWg+36U8EG/cqh+gebY1OBF2eqiV7Ojh6canFUO31RHubtKyRB8urmhWbW
wxddm/qtpRXxqrHCGkf/zW7zTGBctgUSgzlUXQ0Y6RijTizrOy7PxTmCWYBUpdXD
nJrZZuNgguNT3GsokyZN5XQ+k+T+JgI6M3ufaJj/Ve0wbdFbEWw6ucvvubv5UWBn
iCX1aFyBnxOXi8DYWh6T3t0fH+E93ss5OXzkX83TpzumNH68dRwr2fPsf/r9E7Hs
qYB4xBLJwIFYmYWbjhwnLtjsfL605PY6LdCwBfbCNiV6E/nX0959cWwZ/60FKUOl
NavKW6AP7Qj5YdBxTLD5Qu+CL1DqI89l6/iEViiDK2jqvjn60Xa1io2Q205b3nel
LQbrJImThjWZla3kINo5vq8JW46cxJBqEMNTXRwxUUDpTEafFnFanzvr+rpUnZEG
wW9FCrfHV+wQJkXPuuFkvc3VAGjmtnxjJT943i8JZHYY97y8/M3VuokVk37nzWpb
d6JFYrKgCxhcyMzjeC11xyjsHwgYEhhg1E+X0Tchv/2SebPpHTL73hXvOiD/T45b
fHt5HX97ePkxZTOB7plks12dffCqmDl3xql83J5a2OvmYY2G3QtncZJ/6gilJ0Tr
9KsTdS6bmA/aXcR1j+xsvQP+PAbv8tHqn2iCJSeM/2vTXjKB5wuLmHWzj6tjhVrg
lH+88EZ9/0f1XODoPmLbONOj9KrNifHkrj8br4ZjpS+eoJ3d+BVX43cJ2Iv3nsZ7
i4Kx1Oz2pN1e4VKhYm+0ikelZ17E6l2CqlFTiH1zcg0d2qtKl84xwDLTYBB8cJms
pcrLr+bBTcNqV0kLpdgaDOkuxpJ9a8Y0ZuwYMLyCK+SZD9A9BG5TRGSI18ObAgtd
WWNBUebG/+9oxHq4EzDgvdcCH+OWzqg7ozg7HCUwrvXMt/cPCfCzTTgn3AxIQusk
RbJOuODbkfHQ49U32oKEPDsrh8czNbDTy7MCs5yYHbPWzOo6TlsPFdMohY1Q+GOY
AqeZ8LjlmuKXhgdcKraeuiEehKuUTHW2Kl84h5eZUGmvdi3hBmSp7g4TFukwsNzn
fmTVcCKmx9xSv503EwFu48UeI4H1ehLJrI9ak5Wl4EWlmwZzAXQsWAudzYZYFezj
qbg9/7AfsVL8kz5XU1jY2/YWx2tQjerjdoYh02foSM3XBspPtCo5D2MmcrZXuKm0
TXg2BpYJekwrAeNOc/Oy3sTc1googPpbIsqf+3EY+SVC4GH583nyf/9Gou1SF2+z
gujl6zCU37G/Z9SQupLC08DGCpm9SJhW7feAnLcanbaqjbHloSXgKiptvgtijoTg
P6Pe8OUwz2MFxl1C+S+AhrGKxkBCuOkgEhKlBmOYuTMInVMQMbVUvV85VWQ27Iti
u++jN/tVfUfO4fOWPRpHsjQd3MK5GydmM5cxDL8CCVmkFBldCiNKZBd0TDFn8Msm
/RA0XsMoGUNtplMwK8Jng5IjJKr9dLk6uuH7cn8s3vcAjZUbFOpCONYDsICqvIvO
B6SQaNv3lVg21cYonZT/i8YmWcNxHClgEkfj7suLrNiKw1AtmPDLqRizxZLjsuRV
Tlj58IJkNp3E/vD0ITKVSgWz2KH3OZf8oVOaQsdEFOFpuONhEbkym/3FvI9WIcoD
CC3vUw/UyUqTKmm4ItvsVel5JqyrFSUckNy+JNcO4LXK/HC5FM3BU+NB/BKsB0VO
/NPYdJhxiICzXiLepW9mPECFTiWXbbYl3iZuUK5JgoH1UcMewnldhBWpsULqXizY
nqyUGfF66Jx1B6jM/SsE/O3fPEtV/6wBEZkTBt95bzRZVhzfM59YEXuoLS180Gbn
sLnHpYJot0NQErWCMqOsfWXcfaVTnSYRSTcD+ypEU6/EnZqT5BjeVorYA10ZAfAI
1kUmTCc05tMzd30cOJnRpiGgY3ciPGXFfH9NWMwqXDnIVDj5sU7jmVI+l/qsHLcc
UbeAIM7e6UQ4XTLNWo4SM6h/TnJn083fZuVceWplzdtEG054A5MApJ7ljscYomId
tlpiE0BLAV1BDps1JC1SybqiGlBYmOa2k32+/xEy4ULg/a8Eaki0ngyMS16Qi4/V
7dUuWLGvFLAtjpRvJQ76WKs3nyjM1H3ovNgFJb40JMYSGsGmMskN0i6eUNTS6NOD
5OPN55qJgpJVlAOz8+LfkRJOxRFf6WTY18pNa5gzQ4Oq6b6oZVLHzKV9DJu8zkS+
AaQwR0ASrCqmADxO+APfuYUuLrkQrWsbS/lHlqlwms8V0E+jwlhtIBd2oSLBwA/D
Nn/3ggrJwqrmG17rlUsz+4KnLLHQfhV2oXu/rmHPxtlbTTnkTi5GDkrQcxbyti0M
LAeoYsyUlvj12nBYVgpEaKv+n9f7b1KqZaaTb3bwN/K/P+pT/yBDmrpKR1X14ku2
c4SFw5T8PidaokGGMABHcRHmZ0d9rfg0Tyk+QZKryXfQhPFtSiuNjmWee3yHna8u
Ujb3dOCAZIJEEszVhm8pPFJUKJvGQA61JvMfRvx+IM1JpYI6uZGrURJe1ZPXYBah
tQs4Gfvh5gn69WFgx5RGEfegt4OjGinKR0Fej0UdF8jSre+9jlZVJgWkp3dRVloS
cRBBNH5QSFPw7eAWuhb72EHaxE3nrjrj7DGW09cpSggz7CrGmwOjL6y9z9vbQ20w
f6IcRAfSP20aLOr0rQ1PX2mYBpMIOh/MPpsbmkMN3Zc+LUVys0A0OP1DoEpx09Y3
2OUw+Fidhsm3RjXQ1ET3WpWzTimhLAel3cKBSJpCUufEW0+0M71UDUPx7/2iRt9a
gI4+mzbS7/NknCjub6Dw4LMf3kZQgmCeb8vT0l2cL3QFVBhG2IhvyxJI80EZC4k7
ACp+QDA7yZEoiy3amhpMow1wubxGkkfZthqeO05xv+aqfRzbuwh6eW/GSFa/ZXSr
2WXOJX7ZXj9zc/x8dqQ9IudWVmM4QbrAuLgvC2wid1g07n0bant03wIj3FTWEXev
r8LVH2KT9GW4dIuvpLx3bTpadHRmxKj18meTtiaG1kuZOl1NCQOyFo4mX2+Zie3u
2OaVXHjJPaNwRWsDa0Glvq9SHwCI0atrXs33qWQE5COwgzKq+4V9G8rKUMJALrkj
aZIpfJW/2WHsKtLYn+bVZpsm2jh3r+PaV7WDtp+W6RtZNIHXR1SN9kCeqw5q7WBM
IbLPea6BIOERY5O2iFaxojWBNmvzQVvlqdcrqBkZm/7kkGomqKJnGKswXAuBpOba
wJs/VZYxAaqVNoh1xD3/L/eolzZ+PG0kskH/IYBqIhjqPXZzAaHdDLXKhJz18JM2
C41k8PuVP08vS0Apbq8A4R3TOB1r4+0il85d75q1/XC7zu0y7cK+K5lhGmrOMt4U
5FcFAeWeaJFNU1www8d/8phkdbfYsYiFHp9U9E0V9iyB43Dt0xALbXqq8zQAJZ/k
cqcc4UuSjsSU2kKYi5DwxC2PbU70ddGxoi0tMjOiDVmMxRK3EAqbmP29gTdOYlpD
5R3TrS/M9HY7CU+JvRBefohc/ApqOnS4qqk6TVaSGK7SULOXamwLq1K4yi2xS6nt
nUKRpDczEyVnxwQxvbcfqBUVezPiLDBKEdmEH1C8NwBstqRDXl8nlpg1NdPtUjgA
A2RRbKAsS534VxWcET4eEdlfxx0vTw62P128tjdHQDUvWjZc3GYc5DaueQnNmJVZ
un1PWdLbN7WYvlZCcEqzOIHGw48F5gjqH4iVxUthE3D6LBbHa1az/o5hcNOiIQTm
kgPZSGENijyqtrKLrCBesjwOGF+161uClUA698I8dR8PPyVvq56xQ3ClGBjSV7Lh
D9MYfalje8F6yD0YPvJai7k7d1cMjQ0XtgdTE47PoyleUDEVCaMiF4uC0thilpPp
ezL64/B03Ns/7/Q9yYKo4wu16+OT2WmNZPzA2KXksW8TqeLd75nccY1UB+XYUzMY
mAC5fMYSlHZiKBOK1XJjktyIQDxtkcjhkXy1AzhHI9Azz1rh7sVtMcAB3Qf7UlII
/GXO5GFJLDT+qWJ4CJnReuOQVUuc69y/d7LO4Xv0tC3opRdukndgLnTNfNppfB11
eSiCsfDUcCwJ62+gupACRf/05pYpEcpMitmVoU0sEbtPQHl7iB3lqXhhIDlzJh4o
QajgzmeYDAYoMqqTlqovT5mVAEDxANs9qCK/lOL75aO7i1KsKveD9NTImwTJDCYk
ZB2sX+XkKv/VX14JHGnY9yGTpD8p/WIhezNXRFuv6//y1ZVuZQ1ab63IVJffbNVN
1TNmPqukyoS5yY4iSFDKDbl3GqbvHsU90T2gsihr1GAKQx3+dUkHW+c0/jDtuHus
EvLoanz0QcCeBZS+lOFtW2FUxbXOrGmftbiLLCShDwnxQwAXVFFnLJyGOTDcr7YC
FPl9CSFJt3tBvqymot1iLqjIdZ7mohZYxeE5hfxr3riZmu4tEVz86Su+IVnBPVkj
PMTiJ0C54kmpQxvgLR39pKoXLxvV54Ujb+QNcHFMhj3SVf6nC1UwGbHu3fE4TJvA
viODCoBcko/Gvzb2sBaGokfPC34IgElkuvr7qrpSps4X5ycLa0xS1/Zwh44+rKNI
iZxxP+U2zf+g2Bnrn4h9RmjUwrDxTxgldT2by+UcobDpxfAnxNssUQ76UjwE8LnJ
MZYc4tLtXOXj3ulct2nCWHOpOwL230xJoM5iKPrKRc2b0HCx6QaHt1aVGB6on4jM
8TtC7UscZLqHcYSHzPJQbJG3jepcBe1iNxgrlsnR8bobrUtBKUs/7rel6OnlJbnf
c5QXIuyKMsOu0osdjQcykflzbKxuX1+PjheCXYMAO2NZqZGVM70uu07PU+rBfX7u
bMJzi1WTZayLWhBcPdyIcWjIAsZnBcZIrquOJyaYDM8yNgRuiaCFWq0Awkvgsxnx
GwzNqos+GkDmyjlrj9eM+5roXxmuVqAzRlejifXMjIc0vEzSq/irfxk7MT/9uvhC
rkrx09o8qgZYLYNyRfmQbkdxsRn6i9PKX+e1krPVLBG+Cxr0gK2YoGHnCjP5BY5C
bbv3TvuWxEprt06c3XA4ll98+FRy0Kc69aXzTAhsHhZgV2/dx+pYWZSVEhVo+fgO
gUzp+1KS1zo/Om+/WLCAxGKHL/kFOZroVhrKWsnSSNwJFCvuG5ajQ1WBJA10fT/m
JMBFZDe9dQlQRDOd4Bv71sMh+CVfHxl/Vsq6EMBYkZGITlcT10PPpsbrVNh9PC7P
8SQEno61VeM8NddyVLw91i2N9vWsCJ7+E86e/XiCHxco70TwE0QpH65wnQB0xIUT
EQM+/wrxJrp2FCqfYIOYlQ53wd/gkRndvV5EELtu3kd073I1Wj70IBcHfkEou8a5
uKXJYBIVCdUACn+wDt2tDqUgZ0UIxo5XTV4d//GzkxpN7pLswKxT61L4GG45tTyt
uEHD+17xilmiQdg/3S7edvWd5YxW/pWm34x4NzlTNc9HyL5kwHAB7Oah03lkzd38
j64PhJg1Xsxh+RQ5I63D7qyZqVWOGChqtSHKpac4SD4mU3IbqAbhA4Qkb/aiRVeb
IRYuC0f68lmvq4wcnFMUQLPAe6cU/oGC2j/tjHHC6QHvXirF6KeYdG+t5viSNi72
3LXzODG3Ukie8YpysDmZbPLYCaT5CvQb7kHJ1E6YadcFhaNMaACqY6thMWU3TuHy
ThbXS+HAKqLp+PAZQ4VM921kl+2XyL3tYLHzHpmLOwL8g1P8niCq1gZojdxQ2zQL
hV2BJoYlnMngGfYbbiYaVIpCDbAPDop65c0P0GlaL8NHgAUxn1pjD/N4I+jz8Sel
PmybT8jMKV+HyKdz66qjqoKyzaJWuZVXNSMivWttCQaEejU7+XRPmDET7mG2q8w+
1/QdkEE4LKS3igiMOsn1j94FuzmfQz9EUv3aV/m+ClZQEKZLVLgdEfMnS5lOBQeE
fYRqKW1OdZU4YpYzNFzuYv3XdW0mvLeG0X0hPR7CrG2Hvzmo2ZffT6f31ZJBVIvp
L3Iws0nfFH/2vlX5vs2g+YOz3f/+M5Lw4L6XqDuASFtgMeoEFGW3EnkB5uC66ydC
E/C7ZBVZ94anoDF7+OeNu9gpt9DA7H+DDQycOncfPEwha4B2t/0U0weiL4pH/eeb
/uHuuKEn1e1u/Y1Bs0kf6sji5Bdxb9YwNk+S77sJVI9gSaF6RZ0tRIsGsFCjmzyA
OPr2fMMgauj7nS+2FJZgUjFHjurVfP3+f70TrlxtExN9dtdJ1LAxjYYAGC+gzQf6
tyiSJBmdMozKO0/v0dbcWadbyyidEniFlyk+ufFDujWiIbcPgF/xC/nHaCMl4015
4GKcnN0JR0OA+KYZtW/v2y2H3vgkqYeiFYbQ2lGxKwBu2F5vezHb9swSFD4gkFgC
OjhSJpS98OqjcgZdOkB1zs0nonX7oWtYKNljEL566Ymrfxf7SEqTpu8Ll488FQfC
6xQIAyaRnrzaKEME4uQlZERfDpGtT9bRLMc8rCKVtLVKmQRCqsv/X3dbkxsViugV
JWXBkf/h3dFNFkVdjrfU7krV9Vz0hXKcku0bVmEu2cq0Og9J177/SFeF2hZhh/yE
6X0xoulJjT0bASF9qrk5+gaCDLq1cSg66UzlPRLWFLRG6ht2V46HWwf/arGQg+CF
FRo8yd9Dh1vbEeGp4cjVnEKerWqfCAFbiQTYWveSYiKklCMj7WgSPrPNAlcRByU8
BWY7U389o5EcitpayZkEavSY+xn4sOqvhs/kOsMkQopOLvQffXrRkP++n7XvATnj
JzGoHQW0+/ScHrlcZp/Ns41KKt/WNacRjmvEsYIJCg0uHjyc/i1IrY/mRr1YAtFw
jjTgNgXfK9dVcWobjMuJjVwVatld0L3fHA44bZGODChpHp3iQf4oa04lwVJasX6V
6KIDM4efyGG39hwWu/cwnxKgIcv/G6Jh38swFkjH/g430cyr+7GS7j5FeuqRPoq8
ilCOG9PjqmjYFOADx8nMdRPS+9kFDgA2eQJsG7fEfpWizuAZcqihLoLMJ/siASZq
9GV/xMU5kUFKsCYKyEz95lV6D+ysc32AIVgsGxFabb/dtZF3W7ubDSyHxFFvI8Fc
M8rSMnP8nDIWY2ZeqUiJ0gnuPyMxwwNaOZ4BVeWigj1sfG6W92EJ08XKvg2T7fkP
bafP29WIOztf264bEkQxVoZ+Ql+CIynjgC71gdRCiuGw2cv2tNla4WVodrlRb4eT
lFfwn7XT4v/DJOMygeyPnH6EUhP8Zptc+ocK5GyhgF9eDbzGw0j7Jx7Wq7jvtuSW
2WO8Vgky+4fIM1CJ1YEJHkG2KhXYq5d1Tp8c7zpUdlC1FlUBdVrHKU3Ax3MpAlsp
tuUvfk0+gKCtc6wvizudgUQuX6RWVZGU+GkbOBWOEBy41DdUdPdcdyRxfs9WQoyf
ATGDva2BfcWHnMV94CG/aNs2s3PPg3tO8P/pa3gMXeuRqqytgIkMBn44Wp5eNshr
TETLeQE5ncdTuhKHsMM9ai07S+oRW1PhD0Q82V+dvXxkkJ+nbg5BZfWbc1dQ6Vre
oIveWTo6qD7MS8dsDPXlxa2XPATsNB4jfcvSTF410ggv45lWyN14ihErc2OGNHkQ
iLs8iW7o9GSMNlzrJofrpKPoxLE4HWrJ1xrrZR9WBqpPjdFroeRnaZsSuCrvLtJb
vCcKMIZTVSGrbqMSQbXSk63i+IGJBy+57PS2TmUYFIWHCGNvOoXMNFXH9jNMQeLa
8wfwJQgX+jTET2J1R+ehg3RHMwR6HSIRs/BR3ozX2OiVSvon7xqMnMzYr1Be+XtW
6Y1SRUPn9nseI2tbHmy+ThlwPjR9bpOVOxAOc7Mu4ruLYon4EhxEaTxvD5DDmJkz
3tuWiKwABWbN+kxOjWcaCXX8Le7xFgzw4EhE6liGPwX7469V7b3A5l6lgJI33GCD
qFJHjgimpPfIqKz5hsNxgOBbHTdkkSyOI1aXX8PWPL3guCGZD4KsKQpMiHcsbmvP
84SFoWDUp7QO1HBRUHI1FMGLZKUxyG3TUDcKcdcSFl3m5ya03eRIfRYUf51psGjS
IuYn0x5/pthEaShqsUN4R4vkmLAWpp+jsQjO9xKGqRLhlKhnCytqgDKR832Yn9je
92aB+hPikuG9Zg+A5yxB/Xe/TYn2UDiN9XfhCapd2RwM3Q3e2PlBE9xDWR/6gwv2
oruPQBaRmqQ9Mdoio7rZPk6Jv3ehNFqwZaMYU/hGQc9IGniaeAiRLyOZ1Xte8dBM
jPG9v1khJW3Gji9H1m1ctNgJrAQBaV+Jtf4aZ8ZMCfbiiTD2isnb2UgtHbtDLb0m
bVyTrbpY2Uxa7GEKjc2IASyLYyZ7tHhhb39GjFbpf92wOm/NZO5Z4sZvgEBPzxRM
GxfBbfSYovV5PoW3o5bYOSQ9pUDSW2hoy6eGxjvvT96HwHrucqqN6Jd9vkx/pCti
sJgHZ+XfVLHnYzBOuiDH8X6+00ip6WlTVvNvqxum1mnpTtgDNKjW21CJt+nkN43h
RSCzaDW23+FilJqCWMghjuKN+3e9e5A02i3T65F3/ZHE2QzH+MjzWcUmBLpSGIEM
nX4XONSEuy2LP+kfcGG0L4d6zlOXI0LxnHmcEm0nQKwWaJpY6rUbz6nSW/PSuG/S
DRP50nGNdr0HwioA0xpUvOAIk21NW15jgYX3JlVSEYeZ9kE9ZPHY6KuPuuRyJxvz
qaIovQyR1ZBGBzmJfuirHc17A3ZxlMveR4Fq9Cbif0uzaEMsC6tWHHGZUmhbT8uO
qi+5qDfVZzwhjjRvv6GLzNOPNRgsFSeHi2Bj3YXnZy8J0FFaFhtH9WS2WJFxbJAI
klZbLYziVJIxnbYbExVPc99/kY+9WNBxgt8Pye6Wz+1bnZM5CGSWy7SC+aweMEcQ
vtVv8S9GO3xhbXYOGgRPp0nzhs1yseOFpuNVIBwWsPQJnmBqfHt3uSQmJKT6OvBs
IopPYB+yxdPY6E5pLHV4HiB4gIemirGrKEx+mpKQ0slwi/ZlwA6CnRA4h6Uh2adL
yMl8IxG5G9x3btwrFTGlhiuL07DtboaIX+7QJ6YxUKBZLLZayqHd4UdBUJJW+v5C
6aYg0Paxe+ylS6/7wxlgmrKCct0x1YrMybJmX/BqoW2Wnu1TU2R8MOJHIbBoTJxi
WvTRwtCdNs3w8UsUbhMkF0tKgaxrWoqyevB9392nnKSFic9QOnwnxuPf4uGtxMB2
XlY/s0C6ZFAHrvjI/GbAJw8Cxh7pQ/ygSrT8OBuNeKfpk9e+yBlXvQgI+DvGAt4n
huzfsqHLEjosDJFY9OhqiBKxo7FVbci3PZ/nkzo9X+Tb7t4b71fmyRuHU0sgWLse
JQ/JNDWpMF2/zMuq/4jd+BJxuI6iTZKuplE/c0Zd2Kr9CNHBYTRCSySNwxFtB9Rb
X1EG6tJ1dyXrDy7sYAYE0dXZlnd0jiW+m4VwGMdqFYPcnLVTbK0jsN7zxPgVhnJR
oK7BwOiAquO4YFH494Q3pQYWcGsKGJKuXFyPK4cl+msyZ6xzXzTTx5hpnSsKcxEk
TodLCvxOkzEkrJbO8E2P0s5idLxsgwufBKxhe9FbS0jOBHa1zSFDJoI4WXq0QJmT
C8EWPtCBhuO0xZt9sL4LLgVEiz7PBurL2w/OkNRLyqYxQbiT18sssdVX2wxm9RpJ
xEySXfHwnKermnMAR8rKg39Lrk1OQWB0V9tLJ1vRCDhyuaSIziGGPg2UJ+HAQONI
/lG5Tsczoly3xkzXMGRJaMpndp8fasF0D/SE6L6KXR8wTUVXij71XYi4MsG2W+HU
H/96JOjjkkpAbIpT7VLCADpk18c4m4jgf3mcghhNzdxq+p5VfNBBAxrhf4ETaK1V
c+Pzf8/7qWJZrgJ0cMf6pQbw6183JTcoLbUHHwEK7kEJ/RSAn/ObTX/RSz7DbUfm
g96wsPMCH8DVA28TeDvcy8mD5VcGLArcVjxv2RV8W366Qzvs67/No1rxOCdx7JBw
USHIQb+9HfYIywoMxkh/KcIGgCUX/Isni1sEnHhlgldhU0cKOa0PH+ZIRouV6F2P
cDh+j9WHtUH+Tk0cO/2ZZtjVLiNiasUiwzJ0PJPOucgjmAHOatcMHCYLbVwIhdyc
Uuz6BHG5sZ5M8SLkCPA3nSMHxWeX9OpXPNk6o21A6+5jUYaThjDFWt3ou9+jy8eE
WbvnJEPujgCCosZplxHBBD/DiFJ7CXtQZTXsWSaO5lxyYB58u7lT1FshzEAePHfR
4MV1MS1sZ58vaNx4m1vbFC8M6hCDY58Is3B7t1X5XPi4cqamzlbyTs1AaHhtBRDI
snIqkb+7bOvVlzT8oSicXma1nDvVrnjSCod/cez4CatbQQQ1Cx+rCmVmLQY0ZyzQ
xcwJ/iHZWqNY4jLR7FHjJKLpTZNSbqglrgTjqOngUOi1f5H/RbpipWecNXD9w+s8
ooZTlAzUSNOmpA8T/CTdED4DkClN5RiR791a3ok6BSG26LqncF6siTWuFIzFw2ki
V/IfFUMJzA5EWgWroN4kWdoOdCmixnSQXzXl6lBIIQwcu1zHvk6hkQKqkw249vnE
z+5yrdOZ5EQw5znsqtS5M3O5bg/O85MBRuTsi11QNF/h9L5rfHtn5RbL8RqoiQa1
Is04HG77z6I/1tmxyxHPXz2rl6FV+jVlI4aWNyGf7gNLlGwuM3cDKRSbZkNgXUJS
Sn/ufzdX6udpzTOyLuJM3YbEOFH00y7hXRU4FSskJb52TaYbklFflzwHkcWRgvKK
El8t8VlNETBTbobB/sUw/RP5Rjsa85Vyn0valPNphetwQ5n+9akOCIxLJY1jmUX3
yF16v7gxDg4mcNxC0+EmzvzAg2QYfavHS+1NijEy9drPlRw/8gPpr+2q7k4xfAtK
PyI8stn4Sn3VLngUNwFqGOlfEv0Hedqx6hCjgKoSf8G7b6Rvd3CkFX02kmcZ3DlP
9pJUqqr0dMrjbb4ZK9lTphjMQwVQwJ8Vm0Sg0RsXTYqYYHHwSw1MvkcBbQ1DSkM1
sXGkC08xRPJBKnSU8H38yEqZw7eaXHvB9B6E7KZiJlIC+1kSaD2WbaWoMmy3t7bt
DKDxQbJk4YZXw+T0mn8/6Z43Rgtwc6Hzv5aghoDD4CQdWY9T745CEuXPblIZLU8M
PXsZfMhaSVx61cDJrDPIAmN/FJTbu3oW6afvIro1+mLEerfug7OCzHKzvZ/fs4U5
XJL8QFn0C5IaoBfrSm5XlMw4X2Ozqi12FrNqHFRWFNK/ppUwPrsq40AcYwsuvTZT
U6i5RQ+HMR5JrKxRN4Y+ECskqZOpbKR4RXdbYj4eI9hoDoMqNttluHTajUrCkOSD
UzkSiMf0WQOCHAYo5ImBxEWfzasB9Ekfg14Rnn1lP8l0nFJh4OwW9GaYqbVwy/R3
vYO3TQpq5ofmPTzySGJN+VZmTyLdjNX+5cgu2yECJRW+xEaik0Ak36gYb0mRCHp+
S1CU6ANWsAwcL86YsLX0XQGfyRMjNDc5YTWos/Xk0KARMTwu+ocyvgI2aAs0eHG7
eJ6fxndsj314LMqpscUA6qHRwZuxln/p7QYsD2rpsafpvE+dTPg2ESjOJzpWvRVg
JYvIiIKaLctsyMs2YpuGZd6mciNPIPJrjmak5EP9sEbcjKJSb/Qno4BeWqM6asrw
qGIkSloOA1DgjL8R1+/ZWwOTYncgsdHwAniLI3mcaCYQwVfc9BXtMN0ntQNwGrTz
KYaYTcUPk8T5fuHzQvt8gLfxx32o2ylxXXNl6ngZiWIWZbBjNDXgf1fUjS9uVwRu
kqEvM6p/5/DwNASLXWuGSqQH1vN27HJEHnU/tvB9vktHYyAHfkucaue9rFurjB/p
u2y23KA5tgZlCRpHDC1ksNRTllWfav6XprzePV3Atxf7FIfzm8PcC+rts/UAuaGq
mXf7Vm3TjiUzsjMucHzlRkCk5OqoV4vFIOA82lGFE9O663YlLmPrp8NzZ00Ih0Sd
eNeP+VZ9q76cn86dYnBgrqZywEI2MqoshQGsa9J4SPtF6L7WL4rcPFEq2kVhKfX7
GhPp6ABXyMx7Vyrwbftk54z6tmip+JnPLoi43ICD5uAxSq9U7T4Em6S0DnVYcwmB
7nTaX/U0OzK+6jiNrLLFa4VJcwMBIeFkAcVnS8aWeJCr0Og6QG/Jz3toqjs2bVl/
TH3Xj26CbgafCgWzIpTWyThj1H78Xe5c/F75xMfVcZypE+JCAE9vf36W7FsckgCP
mAHG49qYfSwL41YTn4BkaNWRHkgi0LMwgewcKKE+efpF4A6/+AgkUyeP4cEyreSr
LAe50Qji+X6dVhkVELDJoVLa4ZNIZNK75QqlLpDU/tgwTtFztXaUm6GuAi095YeA
8PTUrH2fWW6piCcQdPDJ+ZMFmIO+yWzk7+tmlU7g9hvjjRdopCuo+icVu70UsARw
KmLwAMcafLWw85aYW+NVp/6nnVKFZ7slzfa73sS+aCZatNVIlpeEhzwsnEYZwCx4
zoyJ7BKPmuSNbRM7d9LPkmt+xrUOtAufy8rhQ6PpU+jUPdbOExKvBUUf4NQI2m7c
n4boBwhf2DKHMtG6kS8HVdfufhJHhIwWX+u6gtZGwR7tsbz0EusfDFIXBsy+/17L
6iKrc8Ic0PK1KCxtVnOMxL10oVgWPd8cHr5XI1vevshXljqKzE5Kbs9cPh/Pqif/
Yuf7EATAa/h394xE2swqCp8G1JncW5yKeF6wk77U6qFeJvtpbnfdpDbJGKRhruh6
LmXWNLP4/arSKgEqPSPaqkuUXXPG5WmRkjh+W+57yDyOVrsUTz5w8uLG0nZwFVq1
r6pCgh9cHoKkvwMiIgHwNUqrrIUjMnWXBp41DBwJX1NJhVSV2IVcaAj4tQI/AOxu
0xN51q/Nn1nQQvUOPdAKqwmX5UAkXSNhxJIpPBrqhwBmckxScIvjG/WB1dkBiqWV
l1i8NveB4GcI4IpAiLc3UjlP2ulAMSw0QauHZkEOl/+ITU1obJhtGgtvIMAIb0kX
i6+fI8lF6M9Lp/gjEx8jZXYbwns/hEuJqksuQpF9EDXktxQrn3+QMJtfEMGrJ0rt
0fqlxDCl3GE7gUNGupE2naJmJjHNFdMwzlwtXni9A4RSyfkVsMgHbWrFKE6+inuw
PqyYj1W70YcM7u6guYsbwCAqbs2FoU9WBkW81IGNMceCZA4NoyvJF8J5cN4G95or
TfFiVK4tg6JX2z55EgL6hDSk6hfLeujiCSGKCqX/0hZYEXutlJQMidGa1+g2jFBU
XAHSlJJHO9WeDrS3xOt9tDKMQ+vcjtAcbLsJrXIMuYzQUeZAUK8/v457fpk6t/53
9xVWICtI5YJKHylpg6d4c5QsCGrZzY4e40MNqODvLuf4uLUoIpEyHRbhIbbveyoa
pO7tp4Hm2UsCDaulPijDs242THkWeX1mT2C9VhqHhuF7EHQ495TsPmLklClzCuu1
NOBBC7SkImpzQlqfEqVQmJFtuDlqfJTvXZqeweYTqLMJl87bN1AxB+thVUXbK7/B
xt8Xq+j0265YnduQh4SpUttmVxzqyzEjdzO5GcNJMQaQwP4Ydm8oxdIFt/hljsHp
H4KIbHxeblX4jPPGQSH14QmH8P2z/OCmSrRrw+kjeurBPvh+A7tbvCpb1TdeVjWh
x0Tu1sES8TxDZF533W0K75eqPUcTy4qJpGBFWxFq/cOR69DTmPZUppiQnX3T8PwY
4h6H/K2/1OJJfcdGWvUjRMf5WXAfZVVB2gpP2O0M4DJuM+VvpNkJrSQKMu+SSH4H
X997XBwd6onkmhk335QVveVV24o0NfZ/e6ymBDZwfiUEaWCUykbEfGbudzqhNu2/
GYJWnkJaBjkE24snY6Y6vJ5rN7Pe5TwoubzY2tMuwiw4mysKk0JEDI9TXOoZYQ9O
HiUuCssdlFex1Cix/1qlaGwBi5rq3L6Z2aWQVkYdFfwGUt3foMQlopxv/Ti7w3wE
HcrBGKwCh1WNG2AkzpDhQodZLtsIUx4g9Ho/u2QzRBQsYmRHsbhVDZrtoOMx51t4
gcEblC7u3fHzhmGNyqjmAiqmx7HY9GiouiIJbqO72kGS/8K2G9b7niCcaSn/PRHF
kUJRjyzYKrgznRplDmMzMN9SgDG6V+zL8i+8vVW8pTkJ9oRfmljFiijN8fjCHLLc
599RLHd7PL2Mc90a7saQchhEhIjNR2X+mJLtim9KertwSn17wRxdVw8Gk9ne02VN
GJR6yvAPQZIO8fwKFs6X1N/rP7ALYqkZDzZdjnDrdzarTsfzZvqorUlA9B0L6GpB
ZCo8qE+bUXOsV598PUVaw4GZ8W7V0hKRmVgzdguiu4zFtSSQnr/OEUGijUKONSJs
hVvsv7CURDve20exYZLaMkSUzjBTadqraUFhk2Dl8gFYeRUuJiqJo5m+K9bhlSXR
0A7o75OuYDf1zb9WG9YggX5nUHcoi8LKIEvLXk/aUyhG9QmbjRUJhQGA/tdah3gd
2cFf0/B9r+8mXOk3v7Vc/S/DXBAzBPJ4F6aAW92dEnsDD7238OMnPTw+5F2E/8VH
+7N7c56b2fc+A2SyNDC/ofXh4K+qDQj0mCDvBVzd531KhusX+WLTodhk7h3jSRx/
u3i2ob2nFA3U0KpEXPAEgV1ZQk4CjS5kL+/S+o7X76mNX4EB2kVCk/TCqjXLo1N/
LrLTsqvndajZUB/tmVIJp0gnzBmztxT4IhV31NEciAXxO/VwKzZhB4RaWAs+s4uO
wooUGil5Dzs9CKI+TyMQWTy7x5N2ZW6zFOEvfC8kvWyA7mHNatxhLK2sYbhxJHVe
r1gaWmfM+aC/+Rn6L3DZNbDbQWoxdNkzNW5D6NfH2XTdNrQjUyj4LYF7Kq/uRYQC
9/ap57WFsziYfquQWScGVV3yfNuUiZbhLXwvp9psNPDp4KGn6SVVdV8tS1uVywQs
IlYlK3YKHsZzpo14a9k/AvluM+OLwg0JtpkO26ShcliW6+3E5AHPFk61jtDE3tj+
Cv8VG5r9cIfD0p4xyN2sayD6XuyPlD2kWDSAeVie7H9Ts/1nmrFdWBU/a1IZYphm
cb0OdVlrYnSM9nbRFLc1j3QwXVMht6bHAhG1Mpi8XhjRQ8SPeyo6a5rYAXsGdGId
5mZPi0MAeG5QdggYCzHey0xBZt3UAdmQ5tIieJbRmz1W3xZxQb7+qs0bmXCbVKC4
bVNrz6SUZ1vih6rbWDSqPXOQRUBfGiUZzI17Lm595I1zdn/FjEImVWi5glVaN4kc
bHynaCBN+0PhbqMJzDPM5kp+GhILQ32FUQ+S7N6QDJGXilWJ/R4WOgA2vaPnMA7j
TUjyLz6PvK0IgO60f7EFvOIpEAu4CzyxC9jKhhD4PQXR0YwmyZM+m7SjuMD/7O0V
xo3GSY5tvAIQmjw5vbQWHgX2Zi445z1rw2mcFgzxqFIHLYQ5rTf1DLE0fJkWISlZ
ABSUUXZGXTWalTVlSldMD9rYi4Ujr04vVylW6M+xH7PxSuNqe/3DDyF9Xx3k/jNW
+kB9u/6gAEJ+QOIB3Jssf6WnwQyvAarpFHFuHy9dWPLSXOozwfxcXfvsOekr6b3V
alRg4vGXR55+HcTG2eXd14aPIYbVCudLWHbtSONKn19fyMpRsj/SSmZCC/CNc0PK
iGfipPHqfE4jN2RKgydDIFUmU7cro6VfwjgbsYa+00R5JUAye/WQcI0ebM2p2Zvj
UnCOSVer6WXC1oz8j/GYGJT3ZPOenYRgLgc2+S8+0RlU9fLQ0iShKeEwOGFGVR9U
1C9BV6/Q9Ur60KFUxudFn0wIwJL/gzhwWozLFeaN71bYcSWhtdbUpT89igCayU5S
ePM2loy2clJua0BzCuEf+QIwYjOfddbl1UfWJ9ZdglHQrftknM1fN2WFmD/08HeG
QiBOoGlzLaNQ/sBU+8vk252GWxYHtGulIBHDQKxl0SfMeNfXYR8eNWW+YyEfmIqw
yo7WyqaB2lVt0iNX/OGIQxrRZ5jia9uWoQZR3F9Ut0sdqIvuCzX5ZCELQVfn6rZZ
kdM6+8XUwpoJuoJ1FyRw+Dg4YOATLsrISYRDBOigUgX1cU4EuPuRsZdspSeA9iQ9
7+BrXoLiv+OPZNtsvsno0Dru5bw+ruqBby+UUrRSzkp4FpHx+PSjueguTdD7FHKl
1NEWWoUirATKifIIklbhkX8kBIbWVBEaESLuwIspmKGyIgqj2UeZMZO7tW1gDCKe
cOyCzLDwacRVwf/PJqpqZc+UZ28ubl6yV1zf8Z0GCPXKQeaULYNc+lBcS+475yZ4
qfad3D26dBxY3ocu8Cxe2ThgaTvN1vVp+Ctmpj2qi92wVP558L7wJ0FaKJQ7bVxT
n4hrZCMuA78fv0Fs0sUw7FmWchiXoTipqw/678BomagxAZiSCcwMyK9PVS4qSH+c
BgP44Mb8hITwEZimtM7Gmr6WgvGMp+qwwENkHiKMk7nk5SFIYe9A5XO3+4sr8BWC
hf2lg4PGb5EDopI3D00Tp6l4vH6U3CQfKBSuDSYy/GNFamVEJSmJdEPFKQ6ei+Ve
0qgB3uKsqOYr4Bx3Qi0KNmjv6pgzwMre9YT6h9lfQvXHhRpRyvL3lCDlHWHL6/VQ
VOwBNvfwBi7SZmnkhHIQClcJnBjm0KKpDbmoZaFijQ2vvJ1dqVOmO7YHBIyeww8m
rHCp/M5dU9hkqZAr+Da4hQhObe/zBSx+aQ1iBjIcZuLfIjUjoGpsk+rRQI9sOSYA
P5/Ni+6hEyiHagLPZ4NwkAXodHJsGoXnXOil8HrOhOGzJ/z+1vsY0tp/H+97FGs1
IrlBQpjxtJ7Ha5bdXtCDSPFm47EtBi4GovvgNIFhngGw6KcayCbkTakpZxsh7AId
z9//Cu42o+a+mdzKkjE1dn1DQyMXwRmsTJv8bn9Lm0dh4FSfH7BMhUr0Tp6ANlPK
6amozjl+JmWII4HqTRPR95zU5imqqv8aO7UBccbqPwm5QvYNPlyCuNLYpysnRICb
1swkrAZtfjyku7CG6eWhSQ3rM/wKcSSD36CKLI+vxK6hQBhlkEPHRiBPAvBlUzA6
d+OWKjk99CmIwVW/hSCfURNfEckkH18JgNsAIeHT8VvxG/l55K3dHeKvzuJs6YAw
8Xi6v7XUMjEwcefGBDpgqaQABcxO6qFZstAtXuwixkIXX8qDDYaf/sRfh6BQQJGJ
RtiAOgiexkxgWzmAxAME/1snI9E+PO9l5l6hOcDvAFLNFb900njBeMHAnvcZh/rg
hmjzDjO7RyN/qkWIXN2bttL2qcOdMCOobc5Ze/vvMS3LIxSFPY3Q1/HLP0fBN5tC
ymWs0cMLhtmYKfNflJUSctw0O4IuA7EdRVkgF4y3pvDqtnWEc968Aj7lgCbgs3vK
PciSBeq/qR+ZGPN5+U9bMV/po0lhNUWAXTl760BzRwZi/5dFkLUzQ8rytnZJilYK
CdZxeKDRCdq/+jsWG+EcPo6eHhhrka4MiHWvGOPIMsFarpILWJplTo4YsuSA27DV
A3Tv9UK66IVpC4bMN4HGrKUTEWjHcY7idzltnwq11LxjsLbkRulr0HTcXLLjJiBW
qZeQiWj7Wk4W/7Mbrpy3GFvU4Ap4/13JRIyrnuITRaX0d/XaI1gUQASQfn6ayNta
qnsgABsh6PNhdP7QONF7aDuT0CrjWsj5mg/cTadP7ULdm59Ksfej9f/yaiVy6484
OxcaAHTTAZXoYJXNVw+s3/A2gPd3bNsXge4d5tNHLHWlBesWplTwRDu3X6ktQuFj
boY+z/+1FGU1P0BHdxTwPfkgkn72IgtHOP+mF6OgGINOGfVycO2sscAhNl5S+3Ku
zGS3DzP4VMFff4Ugs5lzGu/bXCavUzaOWw+9/e6tqvT0tJcp9b7N+T5/p3YU+9z/
Kvj7WUYqHFcT1PKsQIWU4h3eP6S5E3JvX6etHm/PzUYVe1ZsKqEChKr/lIzEa4oF
taYRzyvJ1VnHLQkP/BKYRQf3ygZXN/Ul2snjeUwrxf9PMS63hASfjoQCzTlb5EVB
YMPIRGB2K2eHabB8/SV7qrGW/rs6ZI4EJUY7QsGam0vEMzQoKncsGgTfDYy3cLwI
kFHXoTtSqAq9G5u9TJ/pkCWdMM3H9M9KK48XSdErpbWGNlabNo3gSYnz8qTd/peO
04Sg6QcizhTxEsBceVNiAb331O8aJOyydobalHMAulI6LrH270YNIHigttnk3PjE
7SKI330QzIRdfImD76N+0Yz1qSKpKkZ6U5JUEyUCqfPutJSebSDoaVz5p7tCp8Cp
KJZQUhFPzHmzac+Ms1hgEFsW6KG/T3cV9ht8iYCi9qtzOz3OYhsike3FiE4hl25v
emCWBpAWNVlAnr5BUSWcBCt+UcTdqANeTFjPJxFRjpgT52CXlgWeAOZS4V6q27uE
AyUVVg60202wdO0QH9Ckl5g+TrBItlVV1BNQEi362jCm8bvRSEcPTIVElMbKP4N+
dETflHQHHmhimLFgY90oFCKEVgf/6LswvS3lwbgiV1mypYpWmQY4EqmYQa5LH/Od
ao2ebh/svyj7TKzF6XqN3WnGaOXFOfVPYS/fPIYZajyLLUEVUkWVF9zyykek38p3
8tndej9GE32HQc4m4dXSMfzC9uMRTmHbdtryleb+yBer0wuB5LlYBjEz6KhJfy3n
O+Qc35wldLEG930YO4Hc1kfRzcOW7fr1XGkdpvOP2f388W+BCkLJ83f42J/nJnGz
/e1kbxYAWVgzqQ44t5aOcHfeHLq8pXAYV224r/zq9eG1lA7huQFYEAoBLZBjVIct
Gy/GAXX7Gvn2ki+vJCzPQN52cY5W+fh8W1zhdIFIqEHARmh1gPEtCauHPJ/EN0qo
48AslRMy52OOCmNPW3CIwXcK9W32qCdF3hvSO3tOi00VW7ERIpQCffbbSWWdcvcQ
Ghe2nHlmltqfeRIdoBgJmF2z42OPWYGyZnmCno3cFXrMWyKkOpV3XnauzG8rcXCt
sx0WNxh6sjMHsjstP4Hx7atsQuFTIHS0+RBHeAoBiOpC3h+3Af6IapII/GgRGlUI
a01be+XHf6saShafQdwpLLjgJWyZUsqGLiGL0qu+ui7FZROgisiJyE3r6OMOi4XJ
JgDLReF5Y5gFEtIx4tfWQQN7ROiIIISJd8DQFFwllQPLjRxF0ij2UcocRJjzgo4A
vgDDD3dLNHQMEDHQN2upbzaBPmaF7G40XMLoS1L3eAp5LDGDiDAbc0AgqSORg7DG
M0/eOgPFGBAhfCWc/0h8DpbRm6GyPKN5cWPkEIKInNTMaYb+HTLt82yGpJaanbgR
hNOIkIxsV2fVZUpjHbXGBF+iiegxZZUHkl6L2+a90G6Spg9dyV+V/XzNc3ld0M5Y
hQdZL7SKIMs8xGc27F8Un0to+pLIFm8D4Y3CcyhvcuZ8wjoxbaHAWnt3ghRxwgbs
O9GkMP38Sqe8i8RQ7u/olM56qJZh220YJ01UgCMQBK9vvXKnMmiuVRJaw7OvrMfd
c6KfeAILuCVAzLkX8vcqRtdFOwR28IE0khg3kyi+PQE1s3JBbumBdu1tns6mqW+R
nR/NwbDKaFlTV1O5/oxu5Oc132qc/YmpdNbB+GGoU5ZgkG9E05BhbsCAKcDFxzpZ
TVHOP5Lxlq8hzJNFxSgbnDCSQSTm1NJoRmPoQPWEVUU3eH3GwHkuYrZMd2KjV7HS
JzsA8ETGKVe2XAaKUMrHM5EzYrqLklV5pSxMuf93FRsR18+Ymj9rb+0Wv8P5mSGy
YpEPW/WD4TNjShayr+Xxcr+8GE9Pe42VwhEFg1KjgQBKfzGr1D0gtKthELCdvGyM
JFobAtlUabcrM97DkhCY1n1mhQhD/XXAOucPuRMrJ9HiaJnNlaiaA5EEZtLlihtD
CLqAKMsrYv75R2MugGozcmnmSNnQLuq3OP/nnB1SoQUkn3zEagkOQdkNkZDdbuFk
tH8NgRfdVWYJ35vjzfIcEn2dPcgy4ySd1BI62QsPZuyflnilILn+5BbzooDCj2hr
UGEA/ZFb7YNjs/+FaZktaYC48wr7GhmW+hFQhbvUqBqOgjlqtYjh5FH25FX097ck
4ikWEIXLDLy9qEpLZ9CEMtotY2787pK6Jtt1TygQ3/Yo5q36reuiggvQgPie5J8g
QU5TJWCViA0D92zYk9aAm7b+rfgH/TgkUleDXXaU91C4AEB1TJWfDJ0aRIMcsmnK
yDPOtTs3Rsn7qnrw0y45odA9m6mhdqrXio+w6VX4tKgC7ol0FZ/8KUOJ0o3nWcUM
ckPRKJ4rV8b5QbASKa4MX9w+Bj6B6zGR52wxN8RbwIKeeA+/228bioYbi4yf/fP1
xXzSBCohcLFehReG43pfxv5dp/a6fnPUFmbp6vQxKJdDXeC5vXAQ3VRucpDhMlml
J3QhgmFWCMbmC0YYe1S2p4ZRcPJ7ac5DXDe0l/st6FhcU+0b+Yui37uNPCLfp3hv
FO3wrXHYAzHR24G1nKuY4hf6+1MdVmcv+FBXDKkQrCX9BNMSQD/zNId+QLV6bQwJ
MEZgbu0GjeZtTFDnvpSAPtUhLTutGes5TlE8auxBIh5VCbRt7SxeStwrpO+UZxwr
tTViknh8C8eqW/igEoyzvV9k+A2pzpYEx6H5HOqEBvDnNOLyLY2975QOgeJ6fIYW
B9x6XvUTqBVP1ABxVrR7NlD0AnIy+IAOSaFsjCRevgqdI3aSb19+J6sy7jj9Fe+/
U8HBo7OXY8fYqlj3Gg4ldEpO+PKhjQBQXyDO/DVUZAohAgTxvjEixvZgz6bJQtCg
NkWEV8w1qsZAzlwZWUoD3f0NcLQhGdeAyN+kPlh/9s5LDspz+UWEfk20DdpjHhde
s3eacGMmqpVmQ7i/ENrU90DkBoOYPOzMm0Mwm3WEhRVJXzdQjHXMUedB2W9KmaV0
r/xdUGXboW8o+0eEnnLtHFLoEsdcF1TqFcbgL5pdhWhllPmZPuwFV1x6M0o2Khko
DCqenCoteVUAHBXQZdTlxsB0le1ykNadxHdUXBI+ZQNl8HmyfpZ4AU6Z+2YIxq87
3SLYY6IZnUpfb3pbUiMMbuOCOk3VQ2wDRsjEJ+Okxi6IgONWL/yTndhfDhjv7xSN
pXRGv9AnsHS2k6VCtpv5whLPjgfNSkGNYguGjGrbeWQY2uxu1gy1lY8EIMM1SxPL
doPKN4ak19/zr5mBH/uaTxC/0xOg1KTbeUVNAqN+mm3QBC9EvL3xvuzA2bKnA1oQ
KupvSIiiBTShrg7Zm4smFxLUussv7q3lpZ0H2wERhe6wd8sRv1I3aIFQ9P8IwWX8
Gk7JXne2ZJNW4QKP0NL7ZQnlSGMb20rXF7e+633tj8PccVtRd1LWbh1ndAtns8T3
9apEAPRG3tsGjaua8z2N22dSWS8DyyW9LEcOA6eiuvWMsvrN3A8AjC2mBHCOgvqS
ErQAvkyLySDI0XGds8WxYR5Lqi0fi1vX4dPBZmiGBapIeHXgQWSwv1ttgqwnoWE7
/Hlu7cFk/Gafeq9pLONKszXtkrg+UKNmcSxjiRsg1i+aZ2cTEoYdWuhBr+2Sgiq1
E7IpxmXT3IBduH594zXLZ/O5/eHaCBWg6dbYIxVMKM60JzU0gk0Te+bDuY7HCs3h
7kdaPnrsW3AfDkoSTGGZ3pOecMaTF39FRGcL74XhmaMlh1PjhA6B7yus0xn6W6Kg
1v/Y8YcPHUebG0GLDCryb4NQfUdNOk6XyCzkvM7hW4VhHn9Rt8fgKPA9rARmPWGt
XUEjrlHb/wgUoBYMDb4wFgsNV00TacCK22tBHOZsRgY7JPAGdedSg1hJyWgFR8Yg
H/DJtaM4kEH+Rga/0X7PrfkhG3+rfypXk35MMpsaE6G5q3TsiOienVcAssymqkks
s98cX2fa3zPEHTmPVTS+Dkapvsgr/RnCFXdP7PCnCmLIMWulgHbRYXkjztVaJxL3
BZsJ5xGvEzrkB7ATY23Bit0El/PBYZtoXe8MsCEygzQbJJrNnjksjptArGlks2Ny
qbka/rI8YcfjcfjCZ3AlTOWfUctS6l2nQJIObthLChNbghnUJB9NOrKeCywqTeJ0
RBnqNqZiuTpZUrWlTZ8WaP+QeFJrTaMlT4JWm6AHdYc+TsZl1AtYF/2naoOc9L7u
2fPTBMBwbcimqvIW6N93lo+b0OEQyaK+Sp3WXn8jKf1zjgzWB//OnkZeANSSzpf8
bnbDGAOAOli90j07VF8/xgsAzsYmQPmYgbOx3VmP4DDlx08dqRcIZZj590yC+r9z
haJz1doNQgrhR69/hZcoy2ga6o3XOuNPRXodaL/8LBiTtYZzXwzoTFmJxTy7CJne
BqTX9WuRVs+Wlixmu2pX9zQHLQ0NPlXgBElHS5BUzmRlLz4SCnZH31kbmjQ6JQey
69x4bSIE1M21Tjx7p+IjNDSdmfbzl6ac0ekXMWFrtoTJQcczGkpzOImZNnCQmty4
UUeeJQbuTE6+oM8l+U6cgWgv3QPlqNlJa+7FpQ/H2uxubFBpBrp7FaZdEKB8nFkk
f2kjMEgPkCqWzTz8CxwR3hJeml7eYlfhR2syyVnj3WxDu2bjEqQOc9c03DG1CiVb
+HvE68NIOuDnhubFOkE8D599vxCshMaU2rS3JCLvm9x5q7MQtvVcB8LJHEA6M2TE
vCE/UR8YJEjfzCvrBPBUd5XOWZH96/ZQaXgxkjoBHsVwvbyB2Uz2kSkRfWIA7a82
sQRPyCJAKz2rmghvyewWn281s9buNopxB85uX5UVbjxeXs6jle1NdfpVwYdcJYu6
pmNkhs1+JpzwJ0FkY3E2jnJZr8L7Oa/LbmyiHTB8UWjBjtuAM2P+JavJFr/7ov/E
XpRmDDc0QlngqjEUAp163JTym9iLVC7ExK4GPLsM+bsbDZf0ccGthr+7bDvgAr9k
bQq6/Vt/bvHxTPHBNmRp+2253XWYBD3oY1ujxuw3gn37VzxeuBEX1JRvd8B1FrJd
ofR56b+DSWiF7lE8EYXF1u8/8cPNuJfG8elHaxPvoao3jL752LtOGIdbnuSiW3AJ
YBpOle/6zJsUTLwk+uhFtX6e7SWmWRb5WaXA/RCRtoEvdY+l8G3qwmF7OD8dZBVn
ogBU3jx/bSBvLGbc0WwnruOjcM+AsVf0UiJt1ZJ7VNpEvP0dj+kXwvj9tHiiN2J+
QvIbGdVzZLZLu8+BCMalyHrIzHKS7CbGY7FiI4H3E3sxMBMgWrtez8LbWa7Jp7or
hg1zpy2xtedihsMKcrGoVNaRC7ghwjzkMdzkMRomfm5xvurutQurWxR+8VFXQoVe
feh7wfj5/EBsT/kcAUFDELaJkF1sZokrzhwAdI6tgHoy5KJcbE+jkXTC6X6cb0RQ
UPSpsIoe6JnN5lu2LyCfHQ7vzY6v1710L10bi4WkwqLFWXKL8vNEaBMIy4EZne1D
DTNzpKraRcGYfEM4GFIkFOVSrZHmKqnxzxSxz9BERZhOHQzTMVp/WicGljmGSXla
rSa3Ux65thymd9cdGqyJ7yvX05rIMoV/n8RAuisHvaKfDNWprBCv1q1hWFCr1asT
HgV1KoBr0mb0FYSyzj0vBviUFDah28tZTq1Egranbkw8T/tNfWw2Fav84pR579o0
fjjDOv9PgI501v4pU0Vh7OoIJO5C0AMhH61jqaGwk74MhmKZuGGxNMY+GydWXFEW
JmW3SuhavFto6XPKsU4GLBzMoD+kVI9c72lFu9sK6ThDEj33BajxGx/M7aJyblG5
hsgZ6fmAcIoW0ezpoORzICvjKky0q64G86pYQoXjVCDilucG+o0E+2EouFkYMiSS
D61udKbvS0yRzTCVO9kV1T7DlC1SEsm8givKHfobdVsGJ5tQBVXCodXy5XB6zItT
ERJGRz0/0eSOZTHHCBSMsiDJY2XDnrRISWpe9ek3cn2/9vLPDYJl0ZGHC/IrFcnl
BDraWlAkcpMyQi+SmaWaE0EA3WIzScT1vAN515RM2IMkCcBjh9jlq/zpY4qNKR85
JnTNRu2hVNy5vbyBqE78lOHxWcHi2zwKAaAzIXJW52X0w2ydmcCPXrwYtFhqsb7M
oadVTG0oNJWMGjMGdUpi1fYacSDP1vvcqFdLl2zbggMzD3FDVg+yJcYijzHRL7Gn
ie2MbAeHInH9b291i9cucZ0rFcl9NmiEY31s1EImJLaJ32rb69tKA5LYDKT+YHig
XWxKaMji4CI7P92fjr9lj/Xp7j2/PJ7nR6NEIH+IDVBeT2pL9q2BZtHJds7PXsM8
SmA+0RdyVUoIzRAx9K7VpzLdqio2h3RKK9fFVXsun9vPeIsWeaPrnbhWQc1umlx8
0s5RpI9UxcZit86As8e5n25wKXPlNd32Jcr/d5PF2SQylehFrmRKtUTSGmDCOVNs
x4vXVyapryRlbP6FFFHx5cy51ZoLa26KBQ2AMcPFKqphO9lj2v/wC+XZKdnLlN22
ESftucdC8gEz81Y6r154NvRoRuZ2kzAaWfEpMXiscXBC6RyCED7PgvpvieftldJ1
KXxp5wUNaFJbbdprBeW3A0ZOqeu4h9/1pL47t4K+VC/hBjh82/pZRtwGl9rfWbrL
22fY0xFuvPdTv82V4i8vHkJmrSzNQw7Yb96lp0dWyb+UBApiBKxhqk0l/dwFrob7
l1ZLGVlxb1SzYQILUgmBsVNBpVaOvzBpS5bQoE4wthuU/P09nEBPWG/o1+FqOY79
PYySBOmAsKcZVcI3qPiB4Y4HyyrcGYqv54pgW+ZZ8IZBbOenZqQ8Q8vEFk4ZswZQ
qTEwLs4sEU7snkvaAjRl5iClF8/xYysHSEyjLYeCyuOk1osoNVc2wy/ynG0VeFBH
RQb0zBB8D8ipKmLCetMrgbkBJ8vJgUD/pd2sD37W880uGcOR/UK+jkfkf4QZpmlo
jXmezODD53zj+7BQ23wdPnLhxuj+5D9JCOkgjkLDXHjKrn9KXDBIayj1gHM5YVDX
KhofBuxPwfPYjZQK26hP42g2LijlMjw6idZOZTo7DaQpEJuhBo6kETFLFikPnl6/
n63Z/x1G3CrEetPs8yLPU7I9i2XQlOSXR7Q0Yc5jmI4zzwRIJLCHnw3Vp+HEtkXv
FDkO6VeoFIZbEmKOUFpzmAs/HldW8jxn/sRE8ywoQI3t0RdynVFGMNYk2A6fKv2o
Tbr6lH/1VG5StR98kz2mCFlK1ZH4bUDAWI3oeSR6DELObXxT7C4RHnpQ4BQp5Hr/
3VjQKEb7IaS1aDj4z6/nsRajqDVwSNi2pfMTJhTwXKMgR/c11alFuqW/8mO7E41X
mr79wZ65HBbjbutLyK/v8ZyfzIpuOOrIRFXHRCMvPSuqTILLqFOKhoizHS6/0wT0
eCgh+ReF3vaiZotoM5/Ah4H3ikMeEhgdjzKs57jiWSsCWYMkA1syE0EZzcnM+23G
2ji8x5ohoilWDUSmeygyUJ5kkVnctFjlNT6uElXzB/oVUtZgou+tq8m+cgG12Gjy
hKF7jRmSkawRinbkLtkCl/6+nk7AyOco2s9mqAFNZSZdUz+98FHXskH0UE+d4K7w
Kvh4qYnyurfnMATNjhiJfZk3lDomif6P0iS6B2h4tPRM40oraBbJ4kFyeiqg2nqn
lOT7YRTAUbhOWau5TJqHL2wITqcuxUA7bm3AgsrRXWYRWR72mgU8jDWNxBlGB1e1
cER3VKN6rHpv7SLeGd80VV0yUPOpNGVV9yMsjjdAZmdumR4mdUe/MsAdhhDwWxTs
Oz02db3w+icghBNA3oPRXcek9gtDVf5KpbH4D0gokyZkReei6PEl0nalNewrZE0y
LV5gzMz3VfyG6X9kmRt2tyre7dNJMfmWtNgtcYjU2+nFHE04gqXOorINckha5nG4
aCyo7DYg6s4ZewtcRdpUPS6+uSjixjv9Zo4SMkhymYkepUx0zSV+i9rnuRDSe65Z
GavkTU6tVBEHzhWtKuU56kdJYxlCfw1EPJs/93/6zG5C8SIaPjsUuPoQW5pnioeW
N7L+SA7tH3NzFwEfDk3czEhqlFFo4y2K3TcBOf/19KAPk9CnDREMFZaxWgA8xvtu
SY1MNkcIgsq6crAyEEhe9IUrsgAx0po8sXSPDl6aCMHbra/LFJSHrJdhOK5GRARC
UYo1dU7w8wzxqmX3ZQqCjD3xzG3xZbS89LTWG5xhLjtD1j5vfJSmKt4J6nJicVNr
9vfKhlCXJkVsOyiuyavY1xSofdm2C3qxbO19h7TdK58n07WeTTdPqq7MmAsjKyVz
/eBYtH+xIJf4MytySIPKDW43JPSKzZeqQA7I4tFO50SfVXQlnbC5Rh8Ewewsgs9x
4sZ5Sz54owahpEHc16fGXSY0VyZC+2KbB27TduoOgNmFHSyiJTVCcxyw7qpb8UME
w6hnZuRnJthtYx2lyC8EA8F6zj9x9t+ukjf+xrXC7qEfaRd4UssKoKyplzhRjGsK
UhmK5IWjcloS6ooq/a2VwHw6u8HnAYeLpTVXinHoAtrq7hoec0TLD2AriD/p2bsa
fFfub7R+4jiO8p/zoLy73upy1S6ItuhV4WxApSk1XUJr0e7C7dmKxGOAhOAGoLFV
ZbnQzwOBXRYO8+sA1yLX3E1n3T7FZXcEToSv2JhGP7oXSazBnl+9WiNbf2tu3JKt
iN6xYy+Ql63twtn9UgpXeiZNY/0xktKvkT3uP2S2/sHelItPpvOBjjbxgYWTJTDo
U4JGRRuGCRUPMFPGzrH+tn/3SiLP6+OYyQklo4cuTcZvLBH6U05DP4UFxVJ19ZhH
TweUZLkeyhaZW18rP9FhnPeSnsSnAUcNGKg3i6uFzudOqgOm8lAaXdCnEQFt2BKu
oGeH8oi6ZDpEy+oNModVUL19k8iSRIzI/f2f5prY2i2FHEv3NASjeIyfvZS9DC6P
Pod/ib2fiWLPdIR6EOFsJbwMnnPkZQNiFHmRWkPih6s8DMXsHPlpG6CPCFoKhGjD
ybRKC8XTQlw8ugyavgsjLf/8+lw0Wcmm8Gy6gwF5alwopqR+AP6v7YT/pLU5YLA2
kvFpC9t+1Nh9EQgor58HR2GNdZAEV74OB3BLAk8kyB/7sa2EWunrL3wMFu7XHeGl
rCW3461aKwJD2S/R1z1/F+N3643Qdr0050EDbhnzzShcfrDhAB1Ah7h8R3Y2h0Nq
OUAHEqLxCABG74BS8X4jCM6+D+itQxGry7zpvHR0C2WKPe9QUE7tgwvBYSUBIxYR
oIYb+iukpeHd3Gys6ybPX9uldyYMrZpL4OrCu9oYeQQtBD59db0VMLMfTW8pA3Fh
U6ORgmUIutyPDuj177+qqvQUM9++LWqEyGXFlDLpxjvJRqwkdzwl5eitNBKcFAXd
NO8ge0dh1JeFKChihWdalMPnFV82Ryp/IsTm/mkpXh/56c4Ls6yWCbqNFrL4+wb3
76+nGMM8qs9VQtsg+Liqy+oP46CuTwayNWIRlf9WUhQdWrx2lO+f3KhwPtnn/YuW
ttkcgza3wqvuRKZkHpCMmGU1Zs/k867OG7b125/9mGJcFbCn9tkndxHA8bRy+xC4
V12E7EB6p1IdlgaC5TMbZs/AZnUehUo++Ay3DcQ29I6QoBlXOxwPvRKHXn3L8ex+
FzV4KSSFmcfOWdzuWg5X4PPANGyruqvB+KPAc3STZazqV30QUV6TkbrJOfkrYako
o/7DOuZEJpcGmcX8VF+sgyYu1+iA8evdu6BPE+JFRqkZDb+0CvUenTHUQ4/4lleH
zyrAjLo42GcdYeT1YNEBLaP9/TVUTZQBQ+8r3hk/4qoaCxdGDR+I5+FyLR4bsnxt
D40NaHV1iRn9FsU7hbS4SvwegczKq3/WGDHd5cLTY7d2KOh1V+GIteJPibJnMjqf
VR7et61CeudPtmFuKOwyCBUl5lbG30s+JhG1tuu2O6KSiZhXpgOX7uyMg0gE+RcF
pJqiMkPMUk5MSB2E3s3q1hlmPbgLTuYKrzdnMdEagxnxcqM3RFBYpG29tLLdJNug
a7ubFddtJEWE0bS6CEExMREDr+17tfwNEbEZ/pmm8rH8y+LOAVy1z0pvUC7Rp8bE
CN/okGYBK79D4olGrRkNzzNfNorRPIFYykP18CYE7M2/IMBalvJkYoo6AJxTmHgS
itnXVA5pMogMHmQ0d+xh0jzVIQDrtdhCR1REpQ8ZzJH74qZ4biuT/hUWyTHNeCtA
8Ci8VmreXUhB6owj8kQw1cVhbIjq7iPCoUjSuXD3hTdB9GYi3vWTMlsYl8OrWFtx
cLMUKFRdEjs8GYyQyDAXFYM+gPlb6lGBVI7xMXBZS4OH3hZOyzE4VL26CUS7qPET
aj19p2lc29QrJhUBglEWRF1nrJbxrX8d5jbEGtptUMFwLHaTPmvkp4YOfjmv1oIu
CLQAB/RLwKsFGRO0vA17MIdq4I65El/Ag7ZIsLZX7UVBi/QSN8qJRiSOO3kCSmMo
R6QUuDGwumIc2cwkTLgxIMFB+RUqcGOwueMYZ2f60RRia/0oVNZyQQi5d+ihPtfq
VbwgtZVv9BWWuKzM5e3Ph2T4+k9XIU11UDcn8qW1Ay9JJHVqU7bt3fKX/CsUTv+Q
5dS4F64tV4uKYJunNlKY+YUGhfHNZDNx+3vnDAuDlrnoP+zAhuTgxNoOAuMCSZdL
BRmdXXaklxISwTWm7lmFH9lwx6vjRduX7uzvhDVWLLO+BcDvkiOv8/hjkMSxMF9G
3UaLE41a598delCgfm7sukyUaJKbTzIV9F2Q25AAtZdyXbORTS0ek8AKieCP55JB
RkfgcIU8XDSblUlrZKd61T4oJdO/mh0LxezwcxutUZPUfJ4rMTTQxhZcpoCnBqY9
T3wLDAisq9YKrw5WYU6Yo6aUMagJ3mUIwbU6xhIlIPA1fRMNosTr/dSVoWWYcIZ0
sEIuJtRJKwi+wVVcoq1IoUSkdHWCmP53NErMtLoY3dvFIkalG60I9J/tZMi1xbh1
Gs9OjmUby68Sfev8K0ew82MyNZesauSah6in3brvQqqhmfaXPt63R1xw2dt5m41+
7c1/8M22mwI1EtsYEzgWzvgJKogNS/4RCC+atkfj/tsCPqV/7Lbd+ua65EPzfNPu
vhMfZtYTCyLlqSpTWo3Cb3UPcQ8C54oAPAYV+5Ck1mDgVjowm1GZ0b/EK+haQ1Pj
eW59aBhzkdP+MqCFovrvbHE5yyKwki850TKYMjl4DvkxwrfAXkBRZDARiwr96azr
aD9calerpwLKXOtFd0U1l0h/Lw0WO/6+FMfmAiczbCJ3gDvTiIwD6yrGrSTX9Sgh
J6Yc5citEbizuwt7cotTb09p8lLNcEkfrvorBg4akY6OXM6vfxzxHsTLpKrx4QRP
TmFmtcRHp1MsRXJDY3SyQZB3euzQ/c8dJWMXz5R0qv71fxpe2yHmJiKssTjSaux/
32IFpIWYIhWfLhWX0tCNsUl9jjEf5k3qwzmDmjguIENjYDUsSRXrFK6WFuE3RSv4
ZB0pERGChAToKBQpga8GDxcb/0UEvwe2oIzNOC/PCsVHoyqiByud/tyRVOL/qfhA
wSDRKTKABL9lwaYhRL86DpVHmnz23L+L1NEJl4hC63shlnHlxSnzRjbFIx1IxroK
nhC4f4qfjv87XmULjeFbrFodLH37+4E/bth5+czRe91EyXYpREPxdxLJZvGfxbkM
Zg8phNyyvRfl/9P+d0a5o3I8HrW7j7yL0k6n/eq4op97Jgq++eLovtzl/glfD9tx
GHxHKJ/r1sb/twX8a6ExKdKlTnqrD73eeDQWi0zMe8yavJKE8Y7Uy/aMPrUWLN8r
Dg+8f5V6zsW6KFtcHKMyMHhMB5WMcBT2Ypcw1qeXn0FzEcqSkCd5AFT5g2Tr7wqY
5bqKDckqy3t6IZ3a5GwbbQ1acB/8QYF91QTCYyK4E1XgEekdln9QnulUUpnn7yjS
NuC3No6qw72V8GURRM8R+TmNONmai+S6XJPI/QqJaO2oODTOfsOruEPFG/Th9NlA
x0SFQPalow9C/JjcGghtWYTEgxS4CqG1VMizoioUnEug+5FydIuxjzrSH2kZhgGv
V+PdhYZ3fEQkQrQgtqMfVvzMKtP+nAwSUqf6y3dW7hng+/1z21KzerwK+NImPCBt
trhl4ylPDZf41eBdUS34Q0WsqpAmDxcqzimaxFn5Op22HDuXy5ZK7auI5JEeXllC
cK55EjsRxKN+ohMj0qmRYbRaDNBIKMQHYJTrgv1UKRENVMeY0HMM8UrL+l4xdvhv
beuAUs987VOPJUDmKyeRcsp8QsyIuFh7hy6jh65Hcekp6RFEzdtP8kIAQ+/pd2EH
6UgGRQvTGAMBwv6UtyrkMua25uG3oYRAKZ57COssFqCEirLOEFMPKmec1mqFf4U1
sC/TOQh3VN4LkceDhCGRwAYu0lBF9szhxo7mcbniP+geUDprJVst+E1keIkkrZDa
Z95KflareO/Ugg9t92zB9d8SJQUWUk8kJcGLT5PWX+e13IEIO+8nuDHfrf8fbnLI
qCVQrVYyMUYO+fpgonp4KgKN06tP2yvTJ/LN7JEzr6h0zFi9ou1+Cm9ruQBWr0fN
WFjxjePwfzj7PTpvDu0LR3QpawMYJcEV6VAP4MsVIEdbAuFWj+hfN9kaiNC0K/Vu
3wysnDpecGXdKyABKSAbCZfNqJj7zuS0mdG/NgxamCWovnzCDGoWsfVtAcFurG+l
FWuF9iZb8N/clSxeJHgCVAAafqKd8sfyQMNcc6yo6ebJsAU0q5wiEcm03SyQ0emr
rrR9bWTtDPVEEXDxRfzDiN1S4xB6w8p3Lzv/5oyV4/Ma3fBI2X4EqM2iMjGQH+tG
Zc1kYcSmskJFrzvpMs8HrjuzrRVJapSzf+zxHeq0I16YQjU41RQTbEZZ8KlPGbha
MQeCKNpVw0AJQHWCa5WMu/Qxr+Q6QpVLgYSEmDAP1cZyXcWhTapDmoU5A+udCvb1
KrkHQhFlIeWrrjzdfnU4/uifiboe5j8TPMkQUxy70EYqWUnAhDES1P2sF6WLhBBR
Gf/g4YIF9hLdcUDHdb8yPc787KyK6wIlS4sqeUur4SNhjjRms8RQHIuIxO/U9CjB
jG2lLrhvqi4lT4ehs/FTPOY7PbrAbW0IAgQ8eqfEcCH/40dHdzmBomLAbCXocEIX
YIixNq+MsaVHt7is094X3ilnddN8shXGI/ale34CmJyf5O+7cVwOH61HwOMVYTJ6
bDBTt3eIy6P4SUazAWVibjRw5qUmeSPY7KXNEjuSczm3jWWOJSpdP/I8XkkuDhEd
tz1qaX53apQ5yn5NPbLaDs9ql0BqBLPsT1gYKT4gAsXxpPBqpl5cTtDVumCeZnR0
siz5MhbXLtjEkMRFYRY0tysncIwXgjieB4YANy6e0loDWYtFIJOU7I76JH30LJln
CjMeKrtippbdF7As3/CZT1WeIZcY7HUB8Zk1rC+YkVpJn54jwwYoTGydkULa4a2H
I7WmQ+tVHcYcDIDrWKWG/1Vyk7wF2QdWGMNSyk157WFJlCcx8nALU3rtiCeOzkFP
6qrBIaUbx/TaUG+dwlPB3rNys0C1H/rcXcE4ZQHFNwPjO8PTNGj6q6lznpwgphuK
2/6gJsJ1J0p0+56zjy5H4mYKRDQvtIan9opLKjwXcxVc15Bl/QpTgPM5TMT9f9Rd
lLgS9dRBNKf2L/u4sJVclfVYP9keP8M8K7sg35mLUOLKz1I5L1ZLlG6Zz8N+DoXT
lEcjzxTYk//YPmoNjL735S5Odx4c915v1eh5zT92PKDxWwbC2r7jZXRcMcbaR1L+
1O759oZQCWkLztzr123lbOvLbCWTC+PX6xzMIJrAVpkvlyp5SVR19o62CBqsQfoc
i7UFZ4nmHztbysa0ikJrwoYLMhFb64Dk8lhyQZA9xlQZcY8QWaHqwbyyJX0+SlIp
dBkACV60H6KTw6eEgNO5xJjpGdvtRcJbbJDQ3nPqJNjKcsUVZ0ixEXIFljUhIfXl
FTp18zxEEaJwN7Ua1/z8W5gayUqAmH4d6UdRpNW/lGMTRUc3rH/EnLm364H3v0C5
mEnaYYwmRx9kYqRK8qNAOtHOtN2a61PhoF+imPK4vF22lR0ogxt3iOrkWGv4lV8E
fEqVgn4NqQjLEZwHRlI7/d6AznDQ4LZWodmJunJclq2gsU5glmSRVpH7adc4BUO4
73bOnjatNQIXS96ktbiznPuGQ/p9QK2sKlChcTJAHuiMLCdsmyyt7rwbokN9xLc/
U6lxEF17fOS87pfX5WoKJzrTnLCWJjkeoZjqixFqG2+2mdgGg7BFJFA0nwrXNGyO
SD23haVl8yaZixeweOA+HlTmmGhg+USA/LPj0HdaCSsBkXci2HNTSZDGLFcsXNNZ
/l0NtR0eCqsK9KWElU7zEQr5A+A5giT2YzN0tPBpUE8YNunbYBmUu3Y7ng2L0S9J
g0PUtISp3sF3Q/ttKYIEFvh5HPHr0fVxinBbAj1ZyEa3Lzai5o66kH1kJHgdEHCi
p5d/1YCCabubZAbMrpTq5KaStzK5iMgKiJIfebQjA2/VN/fqEmlYMR5ceztmambv
tK0DLE+EbEO9/ZgQh8KD4ToDl8M0rtf6du4LuSNRblnABNSdIluZ8jtB5jcLpaZv
4vZ/cqXUYU5Mkh385G6NN2/Jx+yPxA55gI2ofBlHswGWIERHih6gKSLciB5ovxdb
wco8+8dRGzEYO2fCj+7xaVy1TYoIyGdRUQ29eBW5bqCmkZzkdAtuAaEf/cGyWTz4
RLfWE/bB3WqF4e/RDNxVr6jtDclk7ye+KVulN7jVcXMxDCPtYhuQcrpROQXeA66n
Guf9JoH3bdEI9KlTeZCRnGV+R0/2k4cO8Dmq4HhfsYur60D7SvnPpXZqYmivIX/u
r2aWLhC9SKT3ljg5lgf1zvfdFzA2eY59/wV8JzmHzGgA8d3D6Rd7JWeS3JFonuQ5
76ISctIm37B/aP4mgRZugkCMFNHua4NoXMbyVPou2/ayBiG9upC55enp9fGfwOzB
tFvF9BPss9h/PwicNCrLc84D2vQXGsf9wOo47NXkIk1zK2dBhah3T66H6acm9FeI
lsj5LyhO5dAwwkvIOXGk6tXhL+85wMyYPXbCUnofjoUrNbyQsuZsKrDmOJ6DERxC
RRUUZmquuvB+O1kNFEOuRFe5lk9j7UEj4cM6+EqdDVKJafAHAmyldNcblO4tm/Wz
kAE4gL6OaG38PIAD9oDbiOofEeWODua7icN2C1OglrsJ7ja7bdigHilFeH3cKBrM
5KsfskUvbQw2nOj8iVIyGRAfiqJJ19ecc0bbk+yZr/oYdr7/5uDsVJaUeDDXU7GS
saN6VmdbYtCIVduFbhx0nSRsT06kDSNL4Y5P5ZDwiP4okmBf2iyW6McEKnbrnDiU
ffthD+gCyYkxsZV9CERM0UEEC1dVDMJNwRVmnAxLBBqmHHceEF6NGqyI8sT5Y1uW
LkIpzoJGp/8kBf0KQkoHCDvCeQT39Uud/HMU/X4DRxazxD8n7PiZ598294Nk59GT
jNvwUy4sLQECtfyF0vn2e0bk1D1jNodUfYj4V/VuS0PVC/m1AHSPFtnrVHzysY6N
7+Z9RsqJyZ8RpAuqKtyhlrsqJg6zwdU4NbrY0dRaMOi0IPSPfF8SxV9+jq1XnM4Z
rQsGy0IVvTLZfhrMobHZVNz/IMt13NdoduplRO7kRJ03l00M+731OxFr7JS/JEp8
UbjQ7nOZkG4pFV3CL1Ca4+MqF5G4wxgQ+ltbxXFQ+UiuSjFy3ZBgKoTw2BdEMH37
8u2vul5TmqxLE4Pdjr88G3BqwK88CGEU7aqFfLTY0YibYx44g1qim38DePShOa51
0WJ09lA5e3TaXnJ1pQtp0cX6RAjo4sjmMFapak9F4ZoPBPVL3UC+LL5RgukcY3vO
CqTtwLqfTeP3EMXr64k6flikmrU3ta3jsUclq7q2ZUuZBzBVfEItmRJCvXiDcq9f
uGVIdEQLZt6PLaPsIkUcCXMPvAVxmVnm82Ms/TQi3uXGl+TJIgstgpU5e+1l12e4
/HFYhoZPbbQZnk6apqWaheNmtlqVEDGlnjN1ZACPTddYtQ/nNHODSV2TwHMZ4EBI
Joyop5J6X7emMvl8yAL5pxkxZldKd1rQSorphJlgd6Syo01S9pYEYd8hhJcipnlu
Sevly0+LmjQv1vWGj2eW6bVE2CS6LtQvPCCWFrSmxctjPZ3RDf7rMslcP+LU1D7T
yQRSVJ1xx33JJa1GcXqGul714g+Cx5mGOhxmuTZT6c63c2wiRItbVdvOOH4V8oEX
aaMkA/tmcGZ3EVzW6X+NLoIjA0CnFPIfmXQyQ3XxAVxGKi0lTsQTzPtJS+9b7yMq
4be1oMhTszX2X0eXLlpmfWkEiC5K1AgaaK6nriaAbtqt6zK9c7YvbXkeeYwbYz9B
rsDSRlxM0/3A4tgfFM2brJ3AC/I9MX4Lac89EiVX1lpy8S9bYaWziVfF7iZ6GcV6
i7M/x8QLyt4I725i2BeNSKasLav46h2G6uzpom0IZmsO7+sTzCLGqB1Lk8lF9tG7
I9VvPi82+m/CUtJD3RijrkiN3tsxcQY4bSwwhSVuz//Uxv3m5Y2MDnS+MTm46I4I
TsYqwTv05tTjICRkvJorsR9fADR6F1oiS1lEBxsNTAU819pHNjTMLteJQpgZ4djX
7WjFWUfh7Yjbsn0ZpWpFXGmUq1nP1VVpI1yXoGm3P73Z++CPQv6K6+tLzJIAMbh+
W07+LWiwKjFs1TtD1HgLkM/C+O/Zlj7gv9ENr0F07FgIftVeKfsWcRtTIxb+OFnr
5coZhk28KStlrOZx9R/YJqE4970zqhYrNt9BIVgjbBogDc/XDuCmhcdAJLwhDHFf
5/zAlRBgaxyHhwoWZMy21To52wvP/pXluwhlnLRNP4FTJxAsiRKBqX/H0pJauB6R
tJookdZAv9UfFzMcfmUdR0sdAjY/RTGzBdH2SRMxCe06JW8ZZdO+9tvX1ObY0oYZ
asvSvQ+XwMXMQTGy6ICtEQZf1yXMmL/yH0x/W1EdPuXfcIPqBrKCzwZ4UKoQdmk9
sbT0AzgGsqNuirIrbAFvZg/m73AyiUruKflcJrL4fCKe8eQJYKh3yldP2mrDJMZH
ecQILuHQPuCEonWQH05M/7FjTnwKzi5wYuWeM/tO5y4aTYXyIgD/yzLrLOpLuB0T
w5aAExrI3yDrK3X6vKI7Ogt9gStDTL4VlaEYchYJVE/1Ey33dEvvcnoO+vKorQoO
tUNSyfKjtPv+7Kz5TMWKnm9fLuzcPPiPyeEbykOT9KHf6rqR37rcgJM6Zs1kpmyY
0Wk855+TIUD3Mov1PMkJ9fZRZbb8B7nHilzdMm/w3SJwSaEKWlZbQbyUPcVDQ24T
JiqFDWTyBkICR2sfiAzfmO9pkSwMhtpjWriwNeVYWuAVVnFKUvUFU61NGQ1D2hBC
UyzDiZrlJwSdb7WN/26QYiz/4SNd8EsqnAV0j6ne9t83c+aWA1qb0rqswjsLt9fk
1OWilK9tAHSOm9i6WCXUU0XYYIWUH/Go3K6B+qccCkL8Nk+YCIbsLWmKSapiD66/
4YzM7+E4iBSS3Qk7ACt0kwSU4Z3NAO8ko/ElQzs1F16C1v5Icw6r6R9Kv6oWfsLX
7fEhhATb9iXjBiZXY1bySjapqn7PBvm9r9iNxwLqkf3Qczxj/I/vNWUj19p8DAn6
2QKb54l/68ILbnbJmku3XjTC0zNWDMO1pSUOpqAtGV1DKbA/pc6RzIvHDT2BWSGd
zpTPgfdpnEt6ic7nAY6vzvBVcBgBW2r6A3CXFxXZ+IbZzpu6dStO3SuIixLsiDRW
PBHCsZYNG/nH/Y/Bo4vL/5A3R+g88jvxHspY8LVpGbH1qDWiry7/vdkqyMTOKXvD
wckeBV2xlUbXEHzK0eVj7Rvq01T3stx3hzAFwsRksYvzLeOW5EKpWfI8jL6V7wJL
KEbPT58PQhsmWefjPkM1MeZRYu3pwrAvXkv7/86lUKf6uFKtRA7FrwgZWXqDHYLz
Yc+0JwlLR2uKt4xRiNplgudd2OL9sS+uJPsHASKnLdGzDkiB4/GMzmHxhnP3wnNy
okF5pkyN2NlkWSwP2Z5lyGBTANDOQiB5y+0Urv3/87Hs0A2T7j4OfHjiY4yPR0kw
ONzrOfGmyeoW1toANdH7O7z18DFAwvNvWBkwmOTP0PliWUuWCo8p/mrWhPiEJl68
3oAOW95m0zC+VfHzJYDUNcDf+t2lQsCHegikrkXbCztO5+XmOGxHm7HMcLXWzpzu
IkVzmN058AXQrGZ1NyZKo3RZ+xi9bO4IhK9zn78TR8lO21ccFbpTrkKZj8YcjmZA
iZAaomny3nUp06IIzSP+4X1EiVKv/Adb0UO4Md5po4L7gOAsBqZuQaFnMpZk75sN
BpH6JRPn+YyZRObn+Y9PGppbSdDXF/sBXaEvSGBA6787mj+1InpaE7GBta8hQFQb
Kw2KruPhOKD8FA0fNGL1ptlaYun1O5CNrHUBQSNoZZ+UcYMJ23q2RT6/l6EO1F2B
Yc2XogxuvEoebSgE+Hy+Yv/3spnkYrtobdDu56I4mVmz60PVFAw+CtXzwBLxRVmd
S3aT4QK3/HER2OyviiXtbO1HHnawD613i3bfTdCUPCuJRwVaadHtILIrLk+jGd/T
Dtdya++Io7duibjcByUetS5xMhzcEZbx9f5greEh1m4ks9Nbn3ypSfbuYaP0bYTb
LUti0tZOUa3IPhX+5QmRRzeMFxoeIUjgv5bzZMoDK4Rg3jS6ow6cXUqXA/5VrExO
gdfThPwV+UTvJZHj/DvwY8AUvnkpnUrYxEkxllK/A7GK+Qh9mvG9XFrx1ePGJZsQ
jsk7PGcYiqqdfiV6rqqr9e/nvMU6lDyyuMVjwJMJshw0jmA/djl+cBRlVGU/Ny+q
1/iZLyN+8ovtUwljXv2RDqm44iQuqTETfZWuP4VDAt1Db7XQO6+gmCf9ewMCL/VG
DjSOyA2F7fVbIhaa3khxi4SDq9mtW28qfpO/0rxCvRnvOmIELZYzQVSlJfnLqkD8
e2P/x02nZ43akemo82FbKfYwLeeV05LrJ/52L+H8yt50uxIIH1WSLr90UxFqIXEw
KTEcKn5bwqCRBUZMdll38o/eCXHH7CD1z+5/XGxjS0RSMvraUWjXOK1n6uOPUE49
iBsXSdwGb/0StOmhVUKXuPBiJfc1D2ICLpANR4+CkyYjG43rRKZkH2dfvpPiJCNn
zWqAm/wArZu7BupzA2+i/xb7h4x2F6ZefxQGodGEHqwbAhymxOTYFw3WvDtzSpQT
Ufga1zdc4tDuXIbm1HsvM3Ui9rElwNivguwMQQhUxfH9aXw6m8EY10stDgOF1UOn
hwf39jaWtGakl7+zz2KMziH6lap7KsYsE1toTNmRorwbkZmceJGlJrTfknb1DReQ
NEnHVpuxUDC0U2ZkaSCrPfQE5+CLAASMzm6LQ7qFH6gyyOC0LD1zVyomcm9ee5Lw
7sD3mrURCgHjCb8dDHWdiUO2hJXgedTWNoNa9ce6tvLljLXd1boiz0Tn2jvEIuxT
yQ9OCKnY3rQs9ekey9Mn2OcXIr2ZPve7j9QGcay8sxGjqmf4DRWvPYEUCWiaZ96X
tZTGlQA/h8f/DMEQhT5vbEkXopjokX4DZ2hWBMLNFgf7DHM2xDNo8JXysWoDZo2t
jWYrfDqsABWDC47J/TCKIvHYEo4QuN2ZiyecyUH9X6SDb1T1iaNNznRw+KP45DxM
/7XTsmENpniP+RNkAB7yy5V6KNFGS+OsfCXuX0ROautvIOUMRYPwxNzz5JaBV0X/
PTGX6lTtYDTldeErJu7woJpIsHeh5U8afzX9ZVto24m0/Enx0ArQgguH3OoZccAy
VEjnOmBQiMzHPsiyrHvGQ8M+tf+7m4lEd0n9pLhLbvTWLPMoL+JgMZSDmJpPWidz
RgON/TTQLFnlulNT4jjswqPnPIY8rgxArnS10wSkf13VeFTK4djf2QwmDEnf2HaX
+fi5yz6KwcVtZ/Cqjyp5QnLWbj9Mn7rFbkmgvSC1bDJHfN27l95+3G0mN4icbcGl
hZog1KiUd30hJRgLOevsRief3Opc9n33h6pp849u/SJ8tLlwJ7ACY6yT4hlMWK7M
CK6744d2kNANb8atcc5ipmfxi29dSpyp0c9ntgkj8LEiVu+V8IeTbGmUkg0u/dbz
l5pszKaQp1gRWTxV99HqQz/mQ6ZHPJRLGYd+drUbEPchY/bM70hiWaBx7YYWlQVC
Mr7cMgNwQ6m2QwurmZnKOfs48RgVqDopf0e+EZpkrSnQsEC5rRUEmfZ5aIcPT6KD
WxoxTb/0DL4G/jE4vSYl128ojKcgszW9vV5Rw9POyDYgZ1e/8dSICkLRyEWJBMGP
sX1vmynRWVc+eBE/jRbonrS/Sa6WTj+v9xSEFps4MiqQHwW6PSnM5dspC6fVQdo/
LQdIDoKBb8uSe7yBbnuYFMHM4DQ94lw11c7NSFjyWdTnJqRn9X8JfTlPCOUdN7kP
N/seVXyiM7vLz4xNC9oscoMYbTHuzm4XUOWtwwY+3ZGv/d3xpo+LXcStDPfZgiaq
gZoqGsN3CIxaZxx1WXOnkX3BGEOWVapHzvMHp8T2bJXsoOZ8plJC2s1g8talauxs
4hsnIElIK27fRd2267wdl0PSTAh77p0is/MbMjzBPPrge4AzXrYzML3tk9nZ95gq
vBmdpd6Dt/qgzN8BUCeGd3cRupJ0nnj2VrW4CIfhWfDVMKEYhsre5PlL1UucDFhl
03wdsUzjihtC+i6SbvJ+vrY1iWBN2aSN1rsc8LcNma98f/90N2b3wlPoC35RtZ3E
fcdhjPD0Bucqj8UIUwpaBBDS8lC62MYFmnsDSKwtJyxAQDKkrOVM6DtA/uTYFczU
rF8pI1/8Nn7sJeCTQYFusSafAIEoh6BFBOKQ+x3TdIG1SwdsxX7C+RX64H6gXk/A
danjPU/JdTyuP12xxuF24S7g7PX4qb8kn88gxCVwRl3itHq445Ah19KTZXwTuv+o
0PD1XmT13pb/WtEobO+vqTQ8oKk91NEFm1S/OlsUHnhuOEadZ5HlkDyPhK/MdI6y
gJSORV3JkKQ5B5cUkLg8nmy0AvC7GAj5FOmtHOu8D23JiWoNtuvrWE/AfEb7DvZ5
+BEz/Vh6O5C1r9ZjWGdNjWqvP++LYUYEMPVnBr1VnKILXu6w9FLanNbELpjSVB2o
W3myepd1XvCDIfCgqW7T7CM6fg3ET3Es+11xHdCRi5BOdskrjJfWIoB+AVgLuwga
XjdVLTmA89CPpvMBokCPZEbgtRPJ+/QjtPcececOg2QyGm0rgo6s+I+idqt0miWs
8UeuMxPwFgwKG2OIsVKnWO9g2dAhGyjY5lyC4dvSJV2P39+OvGN06QHzHSlbicYj
+9kRff4RvC+6qa2L8jfGVv0I1ONSUWlES8UMssVUxh3ILStMDNYX/nqSvhTc56bk
wBZIA+/vu2BLyvml1OxvrM6WQd6ZFxJPK8ayfwwSzwRpVD2D/XPpkZYrgB5wDC5N
Dr0efLuWpZn9M3Xw/VsGXQmrrztNEA7D3Be1BkCumSPcVXNU8sAJDhVaKhWL+L2u
Ejfwe85X4HmQrzsh11XQoeZ5sYPElaI5e+ifBg8VGqMYMnNcpXLqNmfTa0Ey9vYS
qX2hlTJxkAOPyoEdUO7ln3MeckpIOXtQdP4Xzxrg42YppCRgdWqiEiL4Qn+WTJCx
ocDe09I/C65CGgbJ77LD5a2pXaGwEURwkVu2cnFkU+tGkaYRLMlSsCeoXKHf7MyP
agxw/hx585UuFoKQ8yNIftfYL7icizqGkVRsx2ysh36ot80O9KET1VB7PntjKUyN
F2yCfYcaS83Veq+LtV3WN0c4vnu3qdDbW/Y/xO1/KUZpcifsAjcMpIsjG2ulVgaE
hurLqQJPoKBx+nmX+7HRpaRACuZNaCAHioBaiLAgT32JFUejKFI76W4p+w3IHxZ1
NBv75Ceh3gq/VcDm0Q/EiiQTZhhjqjCtWNIIduY9I62K0h+TjEoHaA+pxWkqpob/
429dvXsj6YLBFGfrsK4tgJi6DRKFSKFvNWVNI2r0SpCsqVNTYJUx2rt1nIFUmqME
LsW8lpTrJZkuz+ER9hUo6ikkjHY7ljsky+P/RWhvbNUG6dkkJ0xssBTimiU0Rjlv
Bpfa2Sfp9JJqZ5zvrQfU8x51eaqGqpEEVeWgereS/arlY7uxX8kQnZ5D8T+7X2rF
EgIKahJCFyVF/K0TtH277t4g2NuFRFKQ9pY9r1trnmAPasSSYEmmfP3KUSDUxRto
OLUJVDTvEDOzZK/Yhr+SlMyYC3kZom1MkhPYMMBEaJrnTrISEwJ95dyh0nO/HCI/
NcHcL+CS4Sx924YLIjaGoDobx0RWNIVl9WjX3o/f+oSR4v6NrfGc4JVspn+9WVRi
DreS+lQoLvWKO/E4PIcPIl+DdRZI55uiLlPx78V5qjYajM7Xq6r/hBuSl5/kzVl9
Vjn49NHFHr/2Re+hLWWAEZA5c6qgLT+9PNrC8WqeTI85Y3iaUHH+0WAxYQ5CLKAD
sqj1UCCJPm9myHO8EZyraFSftssXDJnUdxHZwfmdvb2yxHXKuOEK9rrQfsfoIVmh
DTjdr7HNqJ12EuRY8ayMbMkdVky5Bm6ZYvXLO5pML5VIhQCxrA6anLpuFpHkBbrZ
Xrz6+NMU4U/1lMNIDECoJx/DKYnZpy5STrdS5tOJFzFldbZWSM/kPtaDQlXUNeUQ
q9H8Kwbmbi0JUHVSNtuINAsqFCM6kKbTK09p2t+Jir6c9bD2dXuNH/Cq8D6HcrWd
7dtCp2Yi3bMugtkEEPIprZoCehSfaRSuLBzKyf4BghZkv+Lk5YuBEgD1s+8C0yZX
PhVR83n41fBMGR/MDw4PkVXytxrxCEdgpxA/NzRAVEVP+VeJon10X0NB1Oqo3rHR
99TFuwvmPwXA09+9bgHhgbxzET4LmVtEhiDmYqj3TELKa5fQreQSuC/9ELQdBFWb
zlaqijpSaahORp1Cd2Hsp0NdyBSYX13gjxKmOm60n/PqSTviVEvM+zzX6vmzzlg1
7m4KgEe460h4CjITmVKjTRSYJRkAMJzSUaZnDGTK4yQL3AchN6gP6MJQOz1pVz3e
8bl0t44HeUb+90GsRse4SUmCrHfleljmS2n+TuC5daB/gQdAANpCYfE5pSddXR2L
kWyl2kATbq/F599TNXuVZVuxEQfHfAmnTgvm+rvbhHeUX6cWYNiddQXwLuTVMMIy
gH9NICddtVKy2BMMHjAhCvPW6uXgjgndRZ+uWV20P2ndGc6adqAYbKjA5be4gLp4
L4p8Z3iTfKzrmDAzenZ/AbxPqaK3qhhEbJkNDK1W+IQ/RoCFgJuLgYuJoZX/v7fW
d+mvNyvgXgv2ROBjxy2tuGr6jRa9ytYOaSnzHtvpIIlju5DTh9eqLSs+PrvmM6Sp
7vWbOxFN16nn6BBSqVqznVM+HlPwywERuVWeIt3JEtsHNZG0mxWPUi9ssda1pruB
5m8w4AAPAYH+roTIgAdyMGOMZAyCdWPRKx7I1xK/+AyO4jWlopCUkXzXxlvs1brI
ZLWgGlLgrN4J5opBwLDBqiO3Bf4mVnlLY/1D5gIfgFVHQGiLrQoGt/GIq/UJIfgz
oOgRZvO5Sl7lVnAWeNvR0dDHXla4kElfqn+pYZUyUOkYY53svh/NZQtVIwNDfxPP
XRKoxvUrLQPlI8zHLRydrtYRRv9hCMCTVQlP+s0/pQrcRx1rWzwLv/CX/ARwpPwI
xoG8v4y6Fj9t3CCnvXGKNI7E5hd7bKTdRnqHCEsOo1kgzDabNZIF4L0uYQpyFS/G
Nebxg4IKZihF/Muiycp9aL66WXhgKLZOSjKx+scPx/WQWpnpLFAzMFzpLdLe1gW/
Ps5wVXqXx8uWOq9zxi08FLm2YwRNYYrwSXO7z82SzzNvpgSmSKqlwXj8x3snwN7w
ZsuEAiribEhUM9PH0d9UuFaMURGSNebMPibGyhP9btycRU66CWuHuT+a/xRwfsGV
D+TccNLFCkwIxpI3y1qtYt4i6n8HDpKwIcY6vYeWiPNwFcp/oRh7VrZIY4AqhpH+
UMp4cs3lCu6ahZFIzEDuv6nm7X1mTa4R9Ho1TXLB1Sk89QBvVj8An0Q+4PlXJ8H7
1W0HgmGvN+FNEZNHLHvdBUU/hO02DZ8CN7Ipvv0W4vExEuvPK41KbzRx0HhroROo
gSjooD1aKZQDRcmGnihpqs2MFaPg3pq/wE42iWfmSbR99TzP9OYTggq9hHiQcZsC
ndqORjd79hIt7i+bNYwPbFg4ArTwVNc2lJ6ggBZNL3+JWjiE3jQo8PeHU7N9qPZu
xnZr2OENV0Vn/bXGkqtZCF2vNamI2xrb0FP3UJrBQGpXDgKgItD6MeujuKd65K0n
IzsY36ti3THxxVCRG8bjEM54iiOUj0vSMcgYvFQDcTqvStZOX7VVxcoPgTpXI8jd
+tQZdY6n3e+vpG+HwsTLTl5cQa5zJDwbtOfe3gxJ/8ONepjpMEH5Bq50IMd+3IRh
SdYMsYyCj3z0qNU+QRJTn9KGwZkolDH+hq1DoNGII0q47RrvrOsXB0JbrjGCGC7C
6XBrb6xG9oEKwgR1Rd9z9ylN3b/bKvMtRRW9jbP8zKVBWSN0nNkjRvqJhHoVubu/
nFjB0hjnpOBvFUoTEH1FJPHKPMoWlJwn4hO7mRdOjfEIp0ItiYE0qy1CdBXQqhdB
RouwFro6fvzWT8cOHeu7Ov+aZv8fsnhJgx3z6SGNFK/7OCv3hgMswgrodepQJTTx
VOx+I0kSzpvDZsyIInuLSolfFAg9K8qR94HTQ3WK2VCd4iFtch+NB/E/Gp1UKzqY
baadvvvN66erMM/UxwLCy9NtgLqIBwOEdeMqk8oQ9tfJ/hlxbQsY4MdP/DPvYsZN
wf/02C3hBvd3PAcWXe5AuXWiIAfh4ef2lEhj89mPYfjH+/v27y179lxhEIVBMIZV
17sWAlqpgTT0nuqtGOllQrS6LpFFeHqVXCuLjkMlgA5/dHmHsVlyFlfThg1AsMi4
Ur54p6IPrnN/lrUeClxFUqHNYGjL/2t3CWRoEKwIBYoCp7DofXib0K7AaI1UiwXc
LxPQ32O/J8art7NEKyTjJ3JTkomWZp1H4B7GvCdNmwNnciEPW1qkrjcTgZSN5g/E
dkhNiNVJROLHUon4p/08K1An40F79Mo2W6YQLp0FiT9ptTp8Dq/HzRtwX5JpL/hF
hhrFugN0WBoHLvwBKY9unydfAF044mgH7hGKpkAYIsIfBCsqg3MM1O0sYP0yLf03
DCv9sC0wxFDztOXZoqKDL8cIM3zDmbqgzoQuiTm4ZCy4QmW55h1OXhi/JokQDVNi
wK6WAbqRsTyK7BW+6R6M/WffZLeulQktwB/yeV2rRYwO0Ykzne0wTblN/EV938sS
YuKtwRqZ1d1wjQCXPNfdY3aU+d2IbtYfzdzTsm0/EYwJatHUwjqQT4DEDao2fxRe
bt9xg+YFqvvGSrkavKDJaPs7tsyPcrfHDJtN1Rfja8uilxNkZMtew9BanlJcZlD0
4sS0AaFWgZNQEIMgbHO0d6LulTXk3MVv3MuCYIwQEx8KWBOPq0U4gFre0eI7BwHd
/gMBaLgPCZ/s94Hxq4f8QVlrRNWfZVFGdeBPU6bdba59JxuG6ChOLgEFq4cvwYB1
ObGtA3OazMA9iKIr1I6LWtZkIdnMZAMa6p+rGasuvSMU2XFdM/Sg4P6m26zYk6tu
gJaT1B7SGPaHzriS3oXyQ451eYw/yxWlRMLxK7yBHudE0f6W8r486LdYLDCSHuIA
+XfajZ5Hv2jHpGJeS8SFIaneGO72fMxKnKVY3ijYmkjkvY/DRSgo/sz+f/TnnwUF
5PSoTHL0XvPjNAyAdICcAxN59mLkcCMLCswcRdncQU/VO6McDK6nK2Gi7cairR0g
p9biWOUPukIs37psn7dlixQ2ktF2X6WwKJGQfdoMWIc+MO0k2HiKqoIYzpEndIj0
T3jftzFXHHzlk6vcX7kK3FKRytxF7ZRFX413CT8HuOs2tlLScKuGYqU8MMO/eoAV
ahdnzIdkjsP/ouYYbwXvjzY6yLj/5jrXEoaMGM4P+eReayZCCBfkjrhMfYiEID7g
bPEtfglJmLsf6K1mblP+htoFdwHwQxs4hpd0Tme2p3zLUn+GgYT2+L2sQOp86Pa8
6JQHwpUyHk22ECtz5qXZ0EKccWIXSN/X5TRBxUrCZJUNmyH0bAZzru4UEooelV7f
ep4Ls6J+/cxge3LfAsPJ58sEmq1LDS4g8F8C+Ov/95eFU3Uo5HEEt9pzJ0NgTY2S
4Kna0BpgODqqulip6gJZiCl4S9JXERLncEmqPNK3KMXYOYGG1jCaIWeWdajvEJad
nm5P1pyq4ReVLSDTCBBwEbTZoMHJ81M5xVG3Tt0KLKOmy7/PvPi6sKZ2dtzHzDzU
jkmDRvFUjn6uXLUSuEmiCQZrOgdeHrT5Gz4yuCwN8ivLgE3D5NscSXxhIWoITZX2
S2HHwRs1NdLbxV/7z9qY8vErWFHLTWcbEkFZk6YhcEE1tWeU0pKs5f6s5jkISkJx
OEneSZgVUB/6qrnP/xUw4nJzEOjO6CKto3b/dgNOM38lE15kp0DBoYZ9gSaBgksE
1AEP2aesYd3CV7M22AQ37dE55sX76sEG623Dm7ztDOe3xREIc8JXjOPC3gfwoiq5
xJh35uNF5tezcuEmSOg2UbFGkKrRKsz85+TIdVoWKTxj84cLrco0MK8tD8Wlkp46
aY0qP/DZ/gLzitO8p/XTeJ8+EFAuQiyUumdKaRIcK5EVd75C/OLJ3IwoGm53d+OK
guyc0Vz6liXxJWjgiB+cZbPCdEpjFK61JCcCR3tYVEE47rE3NV4q/tQuuJnyyCgu
y2SOfaMufDmgdbpNpezzB/VSQZd64kDDY13SjeDKzTGNJRB8dbKgL+fJvsV17oge
bntpIshxo+aWFgSI2M5rT+Lp57x4Nk9NLA1Y9zD4oY9/hnCUD1v+OAJkK625rr+v
jv4cbo9W1EQnY39H4d9FIa0dkLmdO84iai0QP1fHbpPEiZ76D+aw5P/OOjG9jbpj
qqNQZ+EnARul41yO8dKTU5jDALxruGRCR4CR3YmY5aussKjaXWkVp5R7T/ROnjAF
1T+kPWgNAoBYx0t72FQyVPgmXniOPEYEH/hAw0p+aj5ImWuI16AUIBUFULVtAki4
1Mpo9mafpYv3r8uRaBGkzCXEaOJv4RaE978VERvJR60vceSpNT4jF00NtiECqkc5
FzCP2GyYDHE90ZUf967HFJL4P34UM/OIJqzvTZBk5cMNJHj5IwhfOU2kRuubv3OA
TsqI8B9wIABUwVZpw3+/ekFiTPxPrUMWWnfc+xTuFGQ5m4vxk4owg3ODdqbrEeLK
ZMjS4qez9zaYwUdQIBf1dVzmOoT+P9TS2kP5ytJIwTfQzBkgq0moZYGHjFG9e7Ga
OWUqbugUJOo9c8F8kW/0oXfuks/O92PpGbVz9tv2GN9ET0cJhhdQusmB1/FymJ1A
b6JpyjGHKIgGjzvppVtoY6UEX34w/bZLhobQdjFwGSdTqGnCgCNPLyZ3eslg/JTO
6DH8rk+YVtblSE/D0U6XH/KLyQk5ZEM9OnfLM0j5G1X6RiI3X2Ne0OWRswiOVCgW
urMuz2Ya9ffZORaxihKZMC+pFkEkvzpOhAA/IjxJlc9fCcXcFnQKICDGsbpMegfs
v8W+O6dfK/xmBYNVZhEK2kNkyPqGW+t6snhosZ2413JEYbeuxbCAjHV9EAPgYgh5
i72U5x5MSs/gzvqqvXKZagAMI52nH67241RMfHOzGJWwc10Mq76fML6nOESMewOq
ZBEA38ShlVmfxkwDIwUazDRitsH0jNyPFz5i9VQ/Caa/x+5f9qUDIsVJ/N8Kz2jT
GHEDBww0D125NJ+HZ/w9e3SnghrHuYuGHRM3B6BJtmhZVCuHKPwo/H5PfyNXp7us
jL2crMhy0Os4MYz8jsbysiA4Exgeqjnnepwe0cWKRVdSSKsur/02BfDpwINt0Sq8
/9MWoGpDEUsbL4FxBON4SE2hdjTEVqIElYFieLT4VG/APkZvSM/GxpQCjDy4VNrr
C5titiSLSOvGlqoXAPDMVVdq2ONIHEwR+Wr22ZhWkvaE7DTrFU6YhOtvWN0qwgzn
hJA6eqwnMGixuffpvHC8cGv5YmTmVr+0Ij2eLjaJFlOh3y6hZSj0AChN1HcS4cmP
vDHQV0rZ5hw+Aw5InwX86hGBp1M6JqWK16FF1s89ISNxAPjpjtyFeSOP4b4/XXza
GtpmpF7td/GfoCpqmg5cQkfvGZ42IMIY/0fkla810S2TskRGYSqK5Mv67ZplKL49
ScwKxnold2BZt9yEVLALxUTQGljlq0FBe4J0XTKrx7v6+qiEUGgjxn+/0ACU1IkD
liRST72BCZK/n3Jfk+bWy6wEE8dCh0yUdyUay9dlVu6wBrtwc4rO/Qs9IC96/sop
Mqq2h5VAInFxqOH3yJ++ducxLgJXyOn2vUSBdv9tjPgIXzQs2aAhTRsKRUSObih+
RZJkoNIjiGyrR62wk6ComLHHWVJRdK0j80jzGDn6SdrWBy48yd7CuG7PFzRBEa7U
Gip2KPxpL2delkfcX0qWhA7TU2infiSyddAhGZpyMT1v8Dg5yrG2dW6wuAHTlGi8
A4JM4FgMGryAxijuxKpRSnw7uHy4kwhgGYt3HFUP847NGrWtpzDIs5MU5KfW0xe/
j7a1JFm+eXvQ9VO+aeFkj5xczxLeHHggBq/Smxrvh91Jm0lFHCYSycGemo4oJKxZ
sP6RFNC5wLH+GHLsyamyMPO9x9xtma1SpIp003uxYRzn2Lzj3ivz0dWFuDREh9u0
/cF2hYltYppNo8PAkXyZAaV+cQFNKNww0ezxmR+nAuFC7jy/16gyx+kMom6021p0
PWwxVxdjoK6QsWU6i8nUcH07QvvAyCyWT3cXWpJ58J3stZZhrocnwIurz/ShkjOP
RyrHYRrFQloSCsd+SVzkvFwerzHGokgb7+9CR+NDgW1Ia7YSpCgxrLXeqS/gZvOV
jI2Q8Ib8g9R4kk/hl17pxya9DRaogQvhIit5be5Mhq/fVKKLk8xPPlI3h/obUKKS
3cWZU4taj8YUCAiDYLrUq4QHiHgdhtw4q7drNBi7BCh66CjNYSeP2ho8PSlwP3RA
0C/8filt1um0qW4mobHkWUPpksLVJjaEJULCq1OjGiBwyfYgzUvoiJt4YV9iPgL/
c939NtLLsTVw5yU+cISTQ5p3tOidfmxgzbjJFfI5eqEtSzteQS5FtPxiNUjJHnvI
c1KzTQ9qoOzUyXdKKRJDNes76/j0D9VPszRxjOaxU5pjBGfByDKMnx6M2hxuwcfY
iA4SdTh8dOcjgZ37ROE4kKhYpW2XL7deK2bzGimez4RdWidXv70xU7lGn54AXQkd
YA9b0qkHdm/XPkM/e2BpaGehUp2iOh1QK0mAJpJ2c4pOMa4LySPXy1EfEeOtIgH1
Vpx6i9W7w2EYHtLdltOSYPihNc+pzTxS0OX7IYvrVgwI60BzZgtzgVPtaCWKUsRz
xsd7Q8jSepiXgjplnbd1mKFpsVUqX7/O7suMqnjW10C5NiA1iLddkGw/hni3J2OX
yyCY+DxXGlJjFO417IsLh723ik00hHmUgH5cH9fIuyvHSDLpiShVogZACaCYEXSK
SfSxuqPtlPVDskMsuIYOquRi37ejce8Ne9DyGZ1SEfryO7Nc5EtP/1uoJDwj6E2z
0AGwzWt9ZrMLrzo7sZNbA50o8OVKPm+6t/BYmPsZjdI2aaCmMLN5uM2g7Z6MouqQ
3qTZxmxtXVfwkUbtD5bNXyS6+fbZb4BRXFBIHEN4W2phMtR+5TdULXSp2s84Cb5L
kJ7ZyEhGpGqqLtbl075zDF6B0G5GG/bJu+KxaNaqSgnxfxiZkD03a9xX7SnZqpsy
3uWGGWNsAZB3C1GeSLdl6qL2gzuLLTgABex/7lXRiIwsZGp88uKIHH2MbcSzvl0W
t/HmbGi5DSdYU4oKiUt3xqKnW1ePuafHQ2mf0Qs8mkeJ5S/t4dngeXYgXB93LwGa
Rl1FTShpvkaDvDN+19EBp/0Lf5+mn7yomBBOPILG706EAt7a5MZsiOzVmaaYmUiG
sd6Yub7dPw+1vT4RZz7fBUsKUxZtFLYsdhPSrporPyl9hzILuifQYDOJy5GpIK7v
z9HrHdHnS6OACqK/fNqWfum82IP8b1l3irmkRoxOkh97W0hluEok3fcGXSyUxvpL
xsB22z+2usw+v1z2BWCgQ8lP8k0vWrtKcwnEckB749UU/ZTTN7wiluPo6Im3hR8b
tZwxOQgsZHUPrmnD2/NtsVjdIi5a73MB3Zylk31yL3ImxLXxXOc3qkGCIu/Lg45U
PrEHy/5dtiJ8WAul7HpeHxe4APn9G2xmzUnkNXwIWL8jS1IEEbOgZ/H3CjPdZD0L
ravDOWTb4Y2RGD857p6DhJ7OwzhZueO0QSpemlsuEsaC/LqzSiBI6IhE3+ZU4Lrg
dvky8YcNFtEMeXJcGFTkzBtdgybP2sm1J01RlXTYo5IYpT0lVpG8PBOq7H4K67Lt
yWUiSFVLZ73WsnHbGl3kGsBPzFvzWkEeq0ufM/tfqSMMy1MYYzQSR1iqHiKfvVwv
L8+mArSPG1jPmtAQAlZhadRxj8gYUVtCcmNap7Eb/Cf/1klSg8pUF/ABylh3tyPL
4DYBFh2o7QyOFnaRbwO2qH03QCs4KmG6jbtJrmXLObgZT8ipN0xRve6kS9rnnQRM
u7lNg5IK3uwK0rfdpYk5iu3W2n76t3vpJvl8Vd7PUZivqGHDOqJbHXOlrX2ftjp6
RsOnawp18vlI3JTPLz87VmTBQF5/jopRX/UPOTybrZ0A3CGaS6eJbAz2iR1Lf2rd
py7m+WvOy9efa37dhS6AqIvwyn9E28jfDdB7qT362fJfAhb+pqkAwXEzEvOpZqBi
Gg/0enEqCR7mJoY+eqkGAQh9RMGQoIwD9uTx94mS3SL6Kr/xvPhy9I02U7WEu1Ck
CvGjQixVL2IQir8bzP4V2BO9tZumpdxNSKbxxb/TTozM8t6x3Xowz6cYUhkpGXXt
LOGB13kbkvLNh9cquIzcgYrOB+43+CtJGa+FTUa2kYcyXCC890UGqAdtkbvmonv5
AknoFn/5Fqdu8NpSSnWA/0KR11iK3NtxNGKuZpgWUvDlyAkAdOXIVTqiZG3di1Ut
dFGRy0kISetxGScquh4No+eHe9SpSQWtp8mivlWfXqHWq7rSfFsZ9Scfraeoru5N
qS6kyvrJLd21J/rJ+eN16PkAHhBRdjH8aFpLlX2RAst7mnws2u1DyGLcbYrce03u
6tqa99c5ItPWuPfBujxfEIicJHvkameYVSWe+ypX+OlqNCMfTBTMvT4MrL9CJGaP
yrb/nyvvu4AnxhTfwCcKr73OdbcXXyn8sTna4q+mFAV+nvEUhsuw7cuJG0NCI5vP
t1tt4rVfHM79zJGk9rpugmo3ihAEmn3HCNaECdUKNgPKLNYtm785dy3vuXF2tXMW
9BcC7UBu6CBT8tMhWRPRF2x4SadMa6gVGJEp2zEOkT/7xkzjXjF0xAd2jSbGLsSH
klbRkIRE8yJSJHWLS+kXvDoV8QlZdEQ5PO+AnHtdtnIk0KVucZn7px8KzLNmzuER
w/wo1zXxV/gSOp37KWokEHgizDr7CxzVL7vPtFWIbqDh7/jqbbOWxzROKoj+n3Mg
35opP+J4uhWwI7aFDrDXanxjDaOrNw9piDfTzfEP6LV4f6lDlbitotWsVwZQ5cQf
I4z61NEGURF4BHDGITYF2snU0laQ64xOWqSFN+s2lr3S98fMeTCy06x9eL8UrioZ
rWUkPO2jHQRVbG0LUIYq9o84lct3yMwSjqw+RONzuIU8cJRZEUrftYAznsx3J4et
uWYwGroLui/W9sZlDM6w72gM2qzLj0yvgx58QHMkAGvqEfmAVotPsym6WS/FodJy
XN05O9GMQBxcdTJJy1xwSoYV2RyoRoPX/pbZF9XJI1ay5oTL98pADBbAX42VLKui
NFvI1BVEGa3rIDYKn/igslC18ImNlF23GQDBJnRawvt1UcBol5tgi8qmi9avduAZ
snTpvjt3BkFBIWrW+J8uCBfC5Tp0+5lnksw6W9Sr0JzHMxbRB1J5LTk3XPvqZ6B1
4MAvZwyZsch8CwVhoKoRkrpTqRS59nsJ35Qfo91rCXrmVJUgp4Sz2c24IIcnZmJI
nSIf83Mq2wcmG0gl6iA7SQAecAjigQH6rELrOS6pP5jKI+wQKwyLtcfUE0FhNumo
8zuMSxheGMTduOqY8tWj6nOxKQjFd8/Ujm41KFQYYo9ITL/P2UWIhDOO74l8xL2e
Y4Ic6mqQibj7TmtmuFBKVcxbmx8qVLXYEFnDqLLmTsA0kYeDiXLKZm8+uMc0vdm4
vwytCvNwUx932MWeKnPYf+ll061u+yn9ZJ1Zyg7+9Z6eaXV+HNTjLOcNxyPLRCPV
5MyfyVbihlWBZuQ6MRxTHQMhfGMdQ6x13cy5ZV/Mh0d/mmIvMjOb1I+Tw+dwgs72
OwFXA80SazMdlGm8rvrBYzCfrvAsjy0tslwRjLt8elgLE+0FxGg+R36PtgtI5t1S
zHL0Lb8mZaSJ6kCp/t+8byCDsJ9UzTR5MhNRp65APD5Na+WsF/XJhopG7pBmDu/j
emwP0yhe9M8j0aaAvUevLttuljuU6kTHfj23dGsLGvVL8+G2JZaFQQEzq4XnwZqv
BrE2PGNTZOCymaZ7S20bjenKpjryTc6zV0sc4B4A1iiFSMWgTnuyjVN0mqlxfPTV
FGIsGwxhN7to3HloXAeOILei4XT8vAXvoeqwxIxGCTXq4nhexPTK/afj8tZfj7or
2mnPn7yiWnWwB1CSlFLLK8lLj63o8+9H0YUMBiJY7fGWSVAd6phED3yNFo9rXYOx
RxtKQicDA4CF96HzXeO7JXwQxnG3u3fTB3OUeCAerZjDOcH+KT9iffxqnaGZGJwB
nc8kAbFuotq0v8vugV8srDIqKT/nS6CBpWnAkQFcDHJAbibpmM+gw7zRye+r2Zar
DA/Bj6lnp6aJUnY21khLJY/M8kCbP0k9CRzX7BNXTiCP479ok6PltI5n9YnR79Uo
iIZdidyR3DPaKRWGTG4xxIjqBXCOo23qRTS4TcEeiu/bptAtEsUrpnvDxqtu1n1F
mbUEX/2wbW0QgO8TiQEOOrJJ0944cOSvDzieWTNa0XbTU/15d+Be2m5feJfjHjJl
DLlzXYEWnDO7p2of7AeyWV3TREuhoSQZKk4megHyIos7zULzWLeAjA1WFdBHdWrS
vQFZO11FsQydfmSR5d0HwmrgxMMFT9kSxquqOm+igFR1a4LHlCHdOAR4b21NvVJp
j/LKI4oUM2lwkklU52HKmCLbdeHoBR9mUh8shwR7s0p0SHmfCQr7wgdpJyPn6T1x
QMIKC2Y7kLpnbjmKcwWIUQZqby9Zu7muolO3p5t5FdmDbyNFCWwnrljKd8DXPoRG
da69hi1rnSb9gFyLowEO/NWOIEFpxMSITHTKw1gvqAQQI6NMAIkjK39u8Le0Q1M7
bJkbY7kY0lH/dLwSxfxhiF/3C7afPWDcHFvX196OrfX7JNmo2WMAifJv8JLE/n6e
GyxdBTP5pmHlRDcKVQdIbOCLKbJBzPeVcREQrjciaLxDAQbz+QbFTVfrIZiT6+VZ
I+oPviE77jGAAbE6Q41MaaGw9/1MNw6IhnSZxyFgiIpynv0KYN1QqS8/ceJw2ZJc
0dHky5dOnGtVwMvkcBaIR9s2WEs48J9mNW8/uxlqEJWOE5F8VlD9dYcf9t0gOeFd
Jtq17xx/auWuIdRKEv8TBOU2NVC168unPAhasMI2XucjD7CcJK7kvFmfx8SU//Xh
MRZSRjNhK93is4/+uI75IpT7CZ1yZOppnJEFT2ANHxHZzZl3U/h9jNNBJmuHWHxh
hoHjZTUpIyD/tvjmPtebEL1k/j7uD3yguordkAM8sOV/wpPVpXxzBwVEy/605115
xv6R6g3/P7qpjZCnLvXwzn411fRg50vcPv4PK5LxOmduhE77FgVK0lYjbwwlXf8k
50GFJKtC4EFloEOhLYaIVlxNmb6/Qp7WaADDv1UAgRsC811ccqeqigUpY6RHNcnJ
DrKJZfAm+j10ZcnOXadUZZ6iErjSP8R4wG2KKp2vNTC9ExD4eRKmGNLFN2r6diIC
NHQxdR1Cs9zeaKjcYJxBC2X1aWdGgUhbBjFVfgSeRkLTK3cMVWSiEDOYLgAaXcwT
8KiooDRCBNLq2RkEUxAW4azV/uFOfPSqIPzrHSf8FyhmmlZmJlix6zARo00utlrF
F8xl5xX7ukazq8Wx0hjQAL0I7QavS4HwfYGSdpsY8RhsBs0VNyO17sCwciWaVIYo
oJ5HpbaaumJZcklKOByrED34SMluARTzCjwNpc1tOHiXqgwsgNgGuKlrXQOJrwVZ
45WLR6Nfj10hC8jDlWAG5Sy0/D0a8KI9RHg2AhR2JGG+yoZfkizWjP3KZNbdUhcJ
Df/9gKdzXPksJc/Dv514zhfauv4FoKcL8nqowLN0HxzlMHkhE01Fry5iuFpa1COV
SpTxkv4lCn2RFkbLatwgqgshvAny4zYFtMPjWvXJFbALTCOSISeOK+RLlF4mut4F
R8CH2XR9utDhck8bbqUFgGG5xb2INfHQn/8yGl5T6/P33/QgE7YT81kWC3Lp7XrG
oB1OjhRj082Ob3f180FovDNJguPqMI8xAPkazznUWvkeSrFZkTmno3ku2k3TIPkY
vP4N+SHL4o/zaWdqvHmfp6VH6Qun8dOWxqfjCg4zT2nukcJjJLUSoSwIsVi+MMir
5rBQpviGX0St1iZs+iwvQQEK+h701/ooPT6Qv7XNVgqWnLindTWILGb07ZvDD2Tv
l0BUy7K23bDuvpXsgEYOV5/U72Bg+Tyc7rAzH4DSfMvhYUwdVBar83jdj6m9IE6N
LSRQLptJnLUOCxAcH5vDAdjXkhaZoUAiHnZaLqdT52CF2PHSZdWvhZGRQb68K0Ud
QiaW6AJUp9x+sM0hpbZK6wSyke/FjWl7Or9KwrGagbBMHohdF+KAw18CqdZ1fxen
Aoq30IEPuYzkRVMGyu/uyuhM2S55OI/qxtcl9GZmv56L6ni1HWnlYixTKiMAui4h
Lra/zEEi9nsgFgfJuR754UrhEnAQNI+qbNYfd4S4Wj5Y215rrexOitVN4ykh9YLp
AhWRGKVqW5ijTQXSBn5sOz1QE+kzrBBoWuFRmLui+XTX0dhSmwK98UDTE7lIfZjZ
lx7oR7WRmMvvRrhSfLLVyeb4sXAAGFdWJkkQgVx+SgUF8+WXtIDsbaINDd7UAa4H
G8J0EVRbH8v4PPh8EuH29tQRZLJtMemP45TNKxwX2+fCPrSvY5eTeO9CSNUFn/2Z
UpO+i+XdBGsjzhTfJ1ipCeIvyz/T8p6K8f3tMza/vlvZ5yx52dTh3yp/BZlfi329
sS1pnQhMXKZGPz/lsTk61/G/tnoLT2GbPwlGCgwTb9CFFWWETuJjTI1eKDzuhhvT
xdeQ+Jha516aLT/VgOhv3BGVC9nJbGTD0g6RceSPr0xVecjjFPp/OaeJMRmINxp0
akWgaMXQ0zBrhcXICnE1hLRM8i5ApQvV3ex80rX8jdb0CKF8CA6y75ojUfxYGtM+
Mz/dSf3xPUNkhn1wpfW4NYDGtVvGHmYiehGS0hrZys2TXPPptz0JJONUI9Cc0Xf+
UVmGRAeQfEdm7mR4fS+XYcB/e7/agRGokWlEIcR2Dr/Q/1CWM5V2cEflrlSZIPys
X3sju1CIlscs6x5dFEbIOqqcCUYc7oqO2UMDRgggekrPtLt/LpQhyu+lNVKa702x
i9wiVNoju1lIWxyUEK0d17Op60IcH96+zYKwvVOEvqMuLtMJBam8t/Lh7GTpwfVv
YrIixXQ2RPbzOeUPRHEscoyBZLAivTig1G3/L9orLFY9736ve2fD8dWRP2fNoD90
2C5eX/7Fr5dZrrel94lFkAEn3+jKyb35QSGMRdIXSZRE/VMcvABcSycTSwXej1d1
5OaYMnRZGY9JQhFLBKWiFoV5+OiLCgkUPtNhkhQWH3irA9EtSu43R6Dyll2VyD0o
zdAuDgdsK1ja8JyIQbBZKQ3gDZ0X/EHqBBuEScb4+5YYOwMmYljk3YsvixdYft+s
fAkpmerylvM0YWN96XsTzx8wKy5XTlqLlN3x1jKl8yAEx0H5lfDQZlG2fVD/0RRb
qWsPebPxr0fwnO6yLzHTU9JDI+uRNHbLG7zgWTQAC9JEJ8AFE0N6ZIchhgIsoCYu
VijUgBA5vLEav/lwrXibGl/DSAQIoGgEje54h8Xg1NYcqVvoD6Gm0ub9n5OyBh2v
R9LYzoax6KY3AhS3jVCfwCou2wYu9zG7ePHd52cVEiRJ8mcUDm/mMlUFAQ4q5GgX
J18cWqEZ978Ucgy2F2r4YyQ5ZUFCteSU/PZs85UWo7Pvct57Fqny/Oz1FmbHjfNm
fKxzXU4ttF9h43KBobRyPSDd8KZTM3wozI6wV38Bol8KhlLt3g0XDd6/8Ej+3Iab
nlvgDX4J3TEHcdMYZthBNCPBQcsdceiOPJifXwWR6hxiTQtQrw2+IQ24PXAY1fZ1
pKjiFBair7BKJVE5rW0sBJj0Y9GdSy033z/mK3H0rLT239E9JbmgQHqErU/KehM2
ufugUQ0CPjx6ztglo1soUS1rJbabLkYXaBz2fz9NzZCGAVIck529wDQgJMrnIkJL
+qxwC+XKtS3AOEh3K1c0eK3ZdLNhR1VTXRHYqiwu+SCDGNOBu88Cp3xo0fTY+1e0
ROC+IVqQcTFzuyBxfXJoneM96VZUbtMSRXUtt7Zu3DMFf6CcmdACMzWZEiClAif/
msUvRaCQJHOyr3K4l7/2WINQsZ2efZurhol5elkTBtKw7/FAzrXZewWR6cO0D1tT
cbsbSjeQl1A/VPVC4z8pI/QkmmYM3zZwQ/fb1EzQbXABvkvvdzKU3bmssfk/Ucxq
MyEpTqT7OfXEqhuPovFqaHj/NOiiVxpXgumoRzEBkdS5218ukC61rVAVfaM3HUKL
KdpZo9bKfILyBmihXIBpyLP2LG0b/h0cQyoTh1yGFYjIPoLofATggA7hw4Mw708l
bndmWe1PrsGLPyQk7kI4y7DlPNyY51G8XSLyMt9+ZqKYXWezLDLyz1dYk0Jpd0es
MGLjk0YOmbm6zw5hwMeGczqb3OCsZ4yc2nZ/QZPSJ+6LB61JFfInoj0tuXqRVI8l
q1Po64EM+vCjh52eVp5CWh2cUYjS7f4DSNx/EGKaBSjU2FD/17N4kc2cnm6Enpke
Fm8Um+oQiRcBenpcdzJQCi7VbznP0ShrUxwBZt42Z7QTAKdwAJQZrHN010oh+WY3
Plw74eu+wvq2ozlJxFpXF4vmU92eF0FWJWUropJDoq3HjxjvDdwfFfmo/e+iSRXs
ttQXz4WJqmt6OiGpKB0TUJylRMMxtsqz+8RFXdPqRZ6/L+V1LfBRUnBwTv7fkh5T
PetTrOBih3Cbu2G2YSAGujhGrvW5eTKUmuFORBOnfKwgnHMfcW69Md4FdgtNAwGS
MCagpGOVRL8d0CTU5Y8eygcFpR6T7zT7aC9qnDsDpXJUs7ovWxXi8Z2pIofKi1Bd
yxWswTJjdYzB0MdetGirYWr7B5SwRB5xK6rIhj95/RNk9As63Uw/Bvl753jU3Y4K
lZqhNDcfLLz3R97JzbSiAbgfpUbQ4lxA8Dr6SRZTunSeA1/YE1Kldo/3I/TekjIk
aMxAsxFF2R8BqmXKNq1mB0eNUT5ISXQmirnA72DPSVJ+OzhZQqU0PexlBH/WTIaI
iCzC6AW/Ze8lqogU96v/3mVcIfqxi45CCoRPE4ffPL/UpTMAFpZUcbfNeihFOZx6
e2O1Ltq9vbHU+TlFrocDLJtIDkGNWP7/533KywYnMKPXIxyoh7TQwwAKgKTXFsJG
ldJedmPezR+KNs+VmO4T8IHHRmo6BZoHiOx0Nh0wGYzkPHW2du4SdHf9sidm5V34
t/WM/XBDjYCf4V8Qqq5C0AX6Nwp4Ia7ZQDcfmY9xg6qwWexomJL2AGEOwOzWkU/j
PFV9lv2t14B55isok40zIMGvSFAnouNficle+dDN4KI4bo5WKihjPhrv7ZBwN+xz
XygDRK6y3E6X8uhS/qWtzHFH0iSk5l5dWhud3PytJYO6dr8nOxa6anymKMvVReSZ
D9HSfS6FxiDmIxYOOsk0s9wHBOK2XXZU5aaFfn2pOD73NJkp8/UsIOG55PRNGdNU
woy1kd7w7HWS0xJhqtWULLtcS43BegCwKP2QmDaXHjkxWoY5O+jipz/jluPRfreo
4TKO6ZThllAqx8za8GHfHOQZKZT8c+L6uic0metuzxKQIZiwr+tvtIGAmq2/DJmf
BXwIMvU7SdO+Fz5pZzI9AzUJwu6CUzlwr7XC+jCbOMQnu8FOYU4xVk1XVarP68q/
2ofpaa+CSmE1ic+2LTKElQkwTa0IRQyf2nS+53VXT17VEA7fGHEKi+WKeQ6C39MP
l2aMgmEsQ3kvSja9VbwSl+4y4k9oZgEncLH6xqTotRVTQgTB61oGuGUUKMvD0Ocr
2Bs0GnfcqHKsgzEJcuvf+03Y+9E7X2IecXzXKt7xsQEh2wxPDC5flw1v3YF8lUey
gsVb3Mh5vlQUuwLYyqMzwkxncCSL6RyXb9KkKbPFyh1FUf9jwHsQEWNohYpDlTW9
LUmBpTYfMyQbpAw71KWDhh/smUc1BNbV6jNilXhDo268dU5ehlJGzxSZjpg+he1K
guX1ScF2zbUvekzAXdezly1yjHU9GF00nPo8Os8wg9YT9b635H4hGloVbfcxPJ1I
0tQvRm0zwqQVFTfwBXSPiAvA6UX9bsCuXJzabtmKPg2vGpKR+CE0UhtLijzuiA/K
tyl+C/n7XOZrAnO4iKsOKmaYurij18rBOAjbzDSa+YuCaMxntppoPt0+3oue9ygY
ZDBPcs+Chk6n5kVDVqatQsuDEB/L/jdyTj+iFNifB6ztCjpA85pnWY9buvHyM2yQ
gkETI5sub11erfL/aO4NbtNf5tT7h08ZJeFHBEZOHRur+3eAlwKVhMpM83mfnEa1
VqWeksJqQRvoOM+TGqXkEAJTqRAGA7hqNGPVqkLZpPsB18kO244au2D8bEQBrXWU
nTqgBbF273vV20HhKS8tTzMPjnVDfVE5VFW85LYbXmCEYrsw3s6TffS5M5pTNX37
iNyG0PFTsUlitcCohLVXPeQH/O5M0dg7mXskf21Bkz6JhB4ZNl4alB7ev0yt41hy
ZQe7paA1R4X4/9IGFA5wVR7ikRPiwvS3jI/SQ0Je3tF8B1Yg7mi31PPJzZvYiilM
E7C0EE/+iK7Rv3OE8S/m0HuzfaTVobEyorMO2pmb4l4AV+fL99iPRVBB+VtGfaQh
rJ+IxDJIcDeoMlqDjdO5jBI9X00n/grqjob96J5pPbgM1bW4+lSu4zM1xK2aEq5S
uIBp5ji9nVuWGMtTlnzqDJgKd6sAz8KVAifotysXiavuBYgYRBNH+SeAylRI3oZw
QdPDoH6SOw8ZdEHTHMIUwOak2uoEIxlJwlTDauSC3s/1gzFGGhxn2EhPmidH6WIW
RQUnMTvvBBUUC36ugCMUz0uqn55m+gX8qBTQdGiA89i+bugC11fvXk1wQD3jnw8H
bIlH3adcGpLWBDHZSlKHA+h7008/XJ2EZ1ogJtLwaA8FxoWmW8dvhZGLWWsT6LR6
pF9sLzpKN1z2PdFD8koM3dNwg2D8OClokeXOhJ7vNZCFAgNceqRwyx5TGL5hpbaw
eF4Sx4UzstpQfWdt6NZ2dnKYv5YU9T8bnPrf45m9sT1GO//ZTGu0wcerxoOHjyk6
e291Z+nuTWA4WQw+GMq6n5U3U2t2VwHHhKLGTZOGumm4P493KslP0G2i8jc1iyN1
LGDzg5UziVAMjd28ffiUBzyCUasiLNB4tfn8OFcKyKVPC9BdvTphxtDlCY+7llMW
0VSU6jXsNr/7KGIJ32jkx+msoHyf7QQmnarl2Hku6FHnVP24tIaRD/KaSWGKsU6b
cnIwn1RfKz/nLK4eLk90wVeOifipGqz2lQHxUtVVE/wY6oVMoXx167hlFPnUkfW0
OnOOXIrkAhz/dJ5x7fhubKpU2vv2IgUyexmmaOtqmis=
`pragma protect end_protected
