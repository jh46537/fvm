��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG�'���-v_�=@��*�S����k`��sj�a��ī����s�ޔ[�*
���|��kE���,���QK���R�-��-v��V|j�%itt�N�!�Sx�X�8��z'R���Ԝ�	����>2�)��<̈́_�w��Hz�(�Y�Y'1�7��]>�^=�k��g�KhY�ux���q�a�z~�M���U�]�MWi�~�k􍞴�%��X}�+�V۞ޱ�Ҝ0mD�i_"�����dT߈��zb���8�g�c�lw�H:Zv�/���J_��M1� 㤶k��E�({�j�#g�+�P�J�A��x��X�Ԫ]��bfv��*ɤ"��Ayش26��A�`�Nv}]Ѳ���)a��D7�,DR�����m��iW�b%���>�\�*��mOĲ��!���{ޥ|<������)H4�RF��	R����ե?�e�O�"(�~ұ 1�=�n��*tA��3�r�4;V��5i?���D���/��/�n������P{�${�b=��"��X@|���3����)��p���J>��[��*nF~j�368R��?`F_%J pX"���5@d!����3^u�/�2���V(����9�#�y�l�<�ke�
ѝ��|wW�gdƆoDHZ��֨~��K\�b�F�)��)�G���C��};UO�垘���@w|�gy{�Tf��z�gG����8a=N� ���Uܮ�v�;*<y B�pN=����v��R~��L�����@�һ2ĝ�!#���a��g����{^�z�l���poC�dDHݻ5������;&|Sn+b��Mx����L�b��v���E���[���`C.!�x�qp�r�<�O�K;b,�/v��ZX��w�r^�_k������@R�Խ�;8 i�������Y��3�������,�]o�%r�s�,8�-8���,n̪RV#�����~�KE�vea�Q~)U�"�LC4#E4cx������~Y>����=7�f�C�N���FٱdK�RT�*�}��u7��0Y�ْ�2� ����r;��&*PK�1E����p�a�k!FPs��Cm��p<p��I���޼⭊�9a�&~!���<��.�2F
ՋLy�hm���(ˋDi��{�sh�%��n�H�3F�Ju��M���`>s��ZСtL�xB�����W�V�z�+I�[N�F�heS�m�Q�Ӭ����Ey�/�Ҕ{����yҵ��c��w��(��p�˃:#;0������3�	���M�ؑ��x�����q�f�9��f��༴s�N�mJ=͈�����=�����nH+a1�m�4��q�<�r�ܬF��ejjĴ�� �-gb�g\�=�-v�&lQ;ؿ��Q����T��s�]��z�9�^�=���ر#XI�֘P���L��|
n���9��9u������ ]��'�4�����1A�V ���[�M �龭V���#�1&��x�q|���Kޝ&U�������O���"�]�c������V�b�CD�fw;3���9� k��3��a�~1�I���!cŔ ��]<�z�s��m:Y��W�0���L�]3�u\�]�Uyb4~����)��+�]I��r�Sޝ�A�\�N��� :�Of��
�IC_]Ё��\��(T������ֲ0ų>[�ħ�
Y��1<5�Ā�����>ZI��)�Z�)I�Ƹ�kq@1���Z��4�s�U���!4���U�B�����T�ͼ~&#'���O�܇��v`:�v�A�+�?�H�D[#�A��
�[^��e�>0��f�[pU�B���S\�eiF	���̚���A�%��q�b�X���"a*cuFu���{��Y�I]���P�3�?���3d���q����˘p�߀�\@�,�	�	K�����C�͚=������eX�Cb,jU��'���{�����I�����ֶ��w�j�꺱?b�1�1�BN-q�g1/�m����[��?�Bf�r�5I7��T�A!�t�����	��MI���s���E�"�Z9V�zr��0#�����*W��/�M9�\�zbK.���ѿ��f)^�/��Cƌ�����&L�*a'���f�v�� t��QR_����G��L�j!>�k��A9��ĮO�$�,� �3����~�ڐi�=0��B�{n�|�'�qF���,45ݺ�azS %�#�= ܘ!�(og���C@f�j�B����5�I_��SG����*W��R���1m���%�I ��e����.�!��/Z�N�O��.�3��M�4*��3*x3�ȹ퓔����z^].Ǫ��V�L���D�։>'�@c��f ��9}T]����NR���Ǫ�H��E0D4���}���ɠ���I�=�qͮ�{�fl���g��hRcT̳��6�8��PT,��|5��Z��!A]�J1��Y�.�J�����1�҅?
Y��Pg�5�֭����t#q��u�ǝ���+�\@d�,!�f^6�ɵ����E� 	��!\�L$U���^���?~g�[��Y�YS\����D�8b��Ib1�[�G�'ѮY2q����}q��3��HdZGi�RFZ�����S�?�'�u��\,�{H�SR��z �h�+�\�,�v�ʺ 8��3��@_�:&P�C��16�պ}#_@�3���\��Y���^����89|�Ek�ˏ�s,��6M0��^ˎt=��r�8�]��YXuS�7�x�7�&L��.{FN�9�ߒ�O���N�|@�Y��l���.nX#�aX� ��#cv����u-~�K�<3�‟fÜ�(⍘�)^B�leM����n�)��{���N��e�d:8MO��=�P@ZM�zǖ"�D���*�bjY@��zi^!�Z�~���ihrTߏ�����ĉ� ,&��p�j�W� -����q��+�[���6���z�M+)>�j� 3���,�#ʡI:K���J9��W�E�m@&2�6Q���)��T���#uVDs|�n�e�&zW��噱�^Z�d�wE�~I�_f�E���'�r�>�0	��̲
�(e���q�G!%��/��m�����K�%�3��[ְ%��̔�v����`���Ϝ�T��9�ʄ���84q5F�ş�8��U���X\��:�g��R!%�w#ea�g2��e��T�$f�T�a�M��{�K�A_��!�QR>ƿxWE��ar)<��(!��X��������W�����*띂�rA!����:4ɗ��uE�A����� ���F�+l�]WB���+���yDlH�'C%?}���@q�}C�W��*��Q�G���M =+����mk��;}3{���A�(akM�U�2���#�k�����D�l:*Q�5{����^����G�D��u�Z}\#���.쬞�G}��=k4�3Q$Y��&��y�� HM���Qd�FN��
��Z��h�Kp�Ĝz,��g RMz�dY`�!i�]k$�"	��9��lgZ��[�4���IkS���_JF����cI�HzTHm��O��4Ϝ7���r�o�-�;���ڇL���(,�w��a���|���(a��n��U����lrw@}��%D%�LK��8y:�8�C��E����+d���@�S���,c�%���>01S����?2(��00d�	5&��W֮@�c�l��ʋ�
���4�2߻�I	ɧ�J�&ց�7&�R��瑈P��>�kL3�����'�ėM�C3���<���?��ק��f�̲2������<H'^��Z*����^��鼡ܝ<��\tN��ʼ�Q�����#5X��N����O���zz/�愇;���-<S�#8*�'m�6~o���:6c�f���-��r�>�T�i�H�����"hrB��O_���� ����[����E�:����2�a)/v���Rf ��p�~.�lTO(PB'��%��iٍ����q�˅'�	�2(���!�q�����7�_w�O~"4ܒ ��1��\�LO����my�3(�)9�v�5N;P���^��`W�K���ƛJw�d���Z��˝�&�g�0�/����+,��.����kHs@:�������K�c�ͧj�X?p���7y��9�T�R��1�x����K30}�\���d�63/őj\ǭ�v�=/$�}�j�N���)�=p=oD����ᑱ�j�:�r��#?Ԁ k,�tz��ČcN�Xm�?r�
�ij�f�2bܼl2��l�5�����cʲ�5/��gJ�/X�cl�p:���EaX.{�.��,��`^��>�Ww*��%=��]���g�c�c��C��[��lwp�h�ecso�wtT���7:��C������ֽ�ԃ�W��Hߣkm���|@/С����d��|μ�[<;()/�˱��`ϳn��u,1�פm$��	YA�ã~�m��e��;|E����3�1R��s�Q�b.�sl�;hlbIK���� ��/�������t��y�V��qO����NΥ@ԧ���W`�S����A�J�%U�nZ{H�xD3�1�[�kY���o��g�jv�����̰�MD��f�k����RW*p�Fhȝ0k�UÜ�+ض$9�+%Ί�WD3��a��[S �pL[N���[�CD �����Q���K|�� ���&�	{���X&�E&�$�9�w�ek7	*�$�'N��)zN6� �!V�1h��9�Z0�e1����Ήu��#�pNf0No�n����d|鰃�3�,��͗Y��$�F4Â ��V	���M- ��~�h�_����7l��O���`�$ef){D`A����Pe�8�ը>6��Ij�T6��׍<#;וz�J���i���U��]M=t����i1����tu+��k(Q,7�X���Q� Hix�$L�%l"����YFH�5��0}�L�z�&b��9W\��ŗ�r�"�ű��w�ϩ��ٍ8PF�`-y�� ��;c"H�+Ɇ�U�t��o$Τ�f{�wJT��'��X�o�B��~lV�ȶ$�� ��z #g5W̤4�QAL:B���B�Y��Q0�(�Z,un��Ӹ�x1���K��@�9}a���  H+*�O�C��Y��aq��Pm"SAL>%����#Hq��U�J�+x���a�V���u���H*ØȤ����/wSÞî��g��;�x!��P�0�Pt�=�+����liT0 �E��8�a�{-�7��~�L��X�>���eF�<#�N� ��H�+���T �25>���J��-�#5����'����OݭnY���M��>%�⋐4"엑���^	���@��9��?���#�~]��������z�3���)GV�&�<���J%�n5>�[�m4hv�/����U���x�[\��Ur��^>.����.l�C�i��UG%�{�J:�B$��:�{�>B}���GN �i��dta�>}�ҟ����Om��QPN7���5��d̞H�^U�3ߓ_�$��e<).xbS	�e� ��zb���m��{� M�k�ǘ��R�( ���������ڂ�!�Νf�V��^!\ɯ`��A/���i��P2l��s��\�Ĉs;C���2�"�RV8��"���S�J���e�G��8:x<dg�'.��o8��[��֗�V�\�_KQ^J�t�1;�t�^��?y2���/��0ePh�vY��i�;f�YF˃÷T�Y�u2��T����+?	�6����(`�99�O�֠祁�d�igSF����Bץ#����<�,�#�z��#"��!3�թ��le_�$�f�X��g��
�F�(���T�)�b����o�ɯ�WZ�-t�qM&�g��8�6��x
a��W��D@ĦW:�$�o��j�Ġ6��2a~��Z��b��ħA<	\	�
d���I@{䓥:D�(2 6�d�ś���|/3EA�x ?=`�2��R�F"X5��w�l�v��?]R�F�3Cg^�n��J��40iM&�"v޹�h��1�^* ���c*�jC2��������.R��k�M�Z^nNBBދ�9��`�����[��f;���e#�L�XpPV�}+_O��)�	^6�	_o�#;���\T�������|��+��������|��mg���t}V�/џ(�/� m]�,�9���kўTV�􁝌�\z������WG�ѳ�����\��y��o�"�HMz�.���3���(:I�J�s���1�N�{�t�(���c��R�)���>��\�,�m��M6�"�C!T��ԭo�7 �5����LR��gM���6)��h��uЪGk�C�7�k�kq�v�e@a~+�N�M,c�8�Cy�h���n����ꉃi�@=�-�[�L��ɢ?�=j�}
E���B*��X��Z~�<�ّQ����h��}��TO�Pڞ˥�U�ԩ=S���x�����x9;.��:k��3\aJ�C�|ӽ��{��/��l���dy�{��Г�"re���Sݮ�	�Ddz��8����V3��Tl(8����;�'�#���lp�9p�31	<�	=�%�j͐��M���RzT���,?���S���¿��U��wgKc�t"X���L#4������A�Śg�j�t�-ݱ�C��H�y