// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UbcQw8ssfh/OsI7qLEVBaGApYvluWgpdgaiewRXhpyr9NkCXku56fi0Pg7WQOMcZ
oHM5c/zRX98wXBALCG2XVqS6tt24UKO9f9g56kzeTlmCUrjXq6hDa8qLCFcCnBOg
c5K+jhVJmbnOkElWzXjJEzSm4sSeSTPMgGUky+aaUyQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28016)
DaGq4oO/dwXvI7BIRr5h/4z3VvUDmDrigxCKbYT/tMyexkd/R2lJf5IKjMT8if2/
ODcdLHppeQOx5ainFlP0SVPWEd4AYT/iK1CLYbmICm6Nry7S6/+ZgCXuOXxGPcGp
1xVNUKT7hSasfcBBBdiwDOR7LxfJ+70ZL8lyGV5WlvPedTBwN5w+QPVFCBRfJoS/
vbP7ka/O5sSYvSzL2TJnZSFFW21l3Y/u+ZVEshsQVN46yQK3GjbyIqrIAuyxsYkv
RR+qRAclZpFadXR1J7ueuegl1nadt3PCOmRhAXHMsES0dXZDW6dtox4ePAtMUN8k
+hKZp6Kr6Ns1GM9/50KSjNoaT/UPlSB1OJqNNOypeizNemi++lkrk0R/j5O6fh/4
uccmBgMJquf8WwdW7l4YggwxWvELPc58L10IM/xbgYJ4v1coFegw9EbBISSbGrsO
4OxQ9taKwMlKi2xTM5a4szdAeiwcM/GryoiavfMCIQKBK9aFw9Oe2Q7XqHBCUkES
bQOn/h80UJfai/V2FSiYd5RVrn+3olpcpYAN7eaC1vDU34OzaI2Hn3/tZ3EIdu/k
sS4IWMu5fNMjLUU/FUs58UQD/vGVvL5Bp4BaQrcqQJBHsDvq3MYdWmJrnwTR8cki
qCtq0EZIaTSZrSfgsVuAGtxaQY9faBhOmzCFhCQhCWYZ/v7rzYs3UJ5THAgD+5yv
6qY7WF3jBE9zMsFWRrjMQspfeCuyW5B2k8Ns4kXeUWr9lcH2X6+ZgH8mC4dN3zrj
dPDIYNNITaggAvycuzskjDhhaR/8CUfjaisim6cJKuZPzLcsEDV1TRU/sDi9ZjAf
KjeJ1p9axGuEvX5sv/8ZZzjeksioIXjEiPHNACycUlCjNDhZJE9FyicEGCHN/PDm
j8J3PzBLF3lJ0afZObeajQFxSfcS3RTo5/aev2SEKZTw87t+cK201qWajnrwQLBj
WL4ak8HYjR0GaFwMsJ5lLeVxKbkzqEMj7MAdjj9fajc10N3vsXsGhLX4rClAUBqb
YYhNBtkikEnhldFdY8HaoSBDHzC8u8OYWStYqg78zOUSHHfMGtKgDiSS1T5Vn0sM
mL6uH5DmPjk1u7OA2feHKd8AWpnw1/2gUhElOqPwczeLNFeeyrum1bGhumhmbvC2
PJBZAurv5vtu/poVRO0hvTgG8mjh788rhVf379XRGd6RdWIJcAunxsxyp0VHCtFg
D7w/X7LUk+raTz1AmBUCcF6a1IH6eI9eFGeAGvTiTZFi0wCDqnwsTCgYdkM4ky5/
yFMRN4pqAS5EcWqOuMK7XVGYfIF21eNCOzzv3mc+C1MH1yJpVlhnL6XZfkbcH1BE
DaRPCrtd9U9K1kA2sO9Cu5R3NICSz98/n7f9fkk06mGksunplFi9dxAvrN+P0P7b
LfsrA5BiEIWVulyc0CCKeRCU9Bw5v+lKz68gq082WsTmsQF/ae3Z7DZOMNxDzXLt
sSkqkic1Tz+kbKqTI3o9hqQxvFf6yHLu6ixF2thVKFjKXRf0BhJ+jzs05ZBLa+we
cePkIHs8c+RLbRLmMJ7wq4ZXelwhWI0YImRNjUO71xI+W6t26WpqIAh+ff50IrxD
WLhoGUdEVUiHuXkR6a+vUVS1k+zbVWcmF7isblcjVE7sXJWlEojjwct0d+rJEMXI
jJnm0VuzPOhRV2a7eHAvRAK6yEr2TLFvxcR+4w473aBKuOkumZBaJEQu7DCrgRyT
a/BW3V/CygKgwD8n3Muig99PxUhidGGEvwGZt/1b07frd/UpNPm1SNUnbJ4YxbVY
GfNbpiWhw3qns/lchY2BaoLn/KHnnnx3IhqyiRA1VrS2dSGpQOZbWmSv0HEv9dfp
kSYSS00eV2O7wXiwhajc4Z1mIQsA5e7Q9unNnQp/Mdi4/OgTeT4LZ4XwGp236iWK
i1h1RHIscDHoJlSr5FJUscazWCkAmBEf094H9dj2G3mAPspDrWfiFjJZjyFHEUFK
531IKdcJFf7qsIRwVLdN6hYJTxL59M1I/Hloj4FxirqV87YSm06IL+jN2OGfUxM4
RsAo4rtKPRUbq3iN7BdzXbRtf8I1Q40U2BNOF5WjqdFXoe7TouiHEsr28cSKQF7F
VQiPq4W1Z1dfDiR+EXaveISAlapCpbEikVz/skqSChdaFVyRmcsjqslZeARxbSAr
DVTX3dCz6feszPp4wMCgrHDWs7HjIiNQtnQ52FgFs4LV6Ct4LhJEasNzhEncvpx3
zrlrpvOUdWxO0WxKrY0A7U7WokoEuk/Wm+/xctfw11iJwD6sMZ821wE/d0YV5VB+
78HW/GShNsif3zjuMiz3kij9qSIHf15HlmrEiNrT+TYKxv8JRj2sW7W1SjzvviKk
/3rKCdJZKAm/1rF48CTbgWGoml3T7vc9A8zZ433dYpZxvHRWgUz9ZOIMKFcj/IZT
Z+B4tg79Ir8wGt832ZddwfI4SW0UzuB4Pz/zsEgDkA06ASEu6XX1U+WE0eWQs87v
+bHwJOvY8Jh0qyG+H/ZC3gdbyTQbYqZ4RGe5XQMnL5c4qXS6l1iOBZZqC5FR+8XC
NAhTde67Q+iaYJrtRGKYsof09RjkdmWOkJNjBOeaIBxhEaVXu/3NKrR2l+xyYogq
6DuM/rEo0a8rdG1ExcwnS1RBXVQqYh9PX/4a5e1Hkk7fHbj3Ozw+O/Mv7w29ThAT
J4XVrYpL7YoO60zB84U1PT12SYVBQ5aWX+iCoDRoHTnv77rjlKeA5vkc6V5q1dSE
RE0QPJ4eJsCr0VUEkW81yT5SDZg7ulim6xnMs2FFfEKSKYV4ZqzJIxccOeodY0vJ
avx/jugD6RknX21s9YXGShqQFLkEd2DPQaGBDbQwWVM75PffYFGj2bzXu3StdRKm
eDkMYS95FHY/SBhOMOXfALS8UWVkuQHWF3YT+SRu0GAir/qaUa7vjiIfVXsjekhH
ERMgFiZfBA9BusigKiA/dmg4a0DNbM/yzT9F8stT+cczwdhDqXJqGQfJ6wCiM8EX
ODBRz+5NUFX2jddLrtTmJQN5ORKJMlmpAfhIOHVp7pyW57Err3+52AG0+jVOdDlD
eqQGQcHk+4HcGrVgrW/L4FebLIjbt0gCxeE6xXkdA012Ar8JI6a618pXgKSp7hCZ
Xf1NEBWAh1lQC9b0YZdhhtLSvYh2d+lObchIAeBVQP2hG0C4Ycz61uooXOLl8P31
IoYUB/57Iiaf+XSrjd5rXbOZn7eyQCtwiMM/HAcOGrGzg8j2sVDz5+MN98egTa6P
VIzzbJtyuoYvonaRSjk8sfCXN6xFlpXtbJK51A3jX6x2hXWed7gH4rY3fouJ4lr6
TqLQr05laukWJlWJq5SQuifoW2ShDpLbmntXnN2EAo9KEvlbgwHu5aeP8fHLNA4A
EZz90F9Q+i6MdjVtLY7646Qaj3rBhepK9Cui/ioAJ1jl4YqPz8DefeZXaXtwGDmo
mak9zMKhVNJXwhiNzf4yTp77tu2nWpZ9xd7OlMWvxEbYzGUkZy3cxx94Vpz+yV39
qqCvRrMmZifqR/dVJG9UEJb/YShPbaG5hg9A8M6rgYBNWL8oSw/xvRrucNDPbC5F
JtoxOxOJtkhsE03lHmuzvADfYcPO0CWBL9v8lZOW/Pv46FtD0cYc+8r9z4c41B6f
PGGiRTa0jrSc7kJvtxEseFWnZC8iNs1JBuwEq9hdVUUFZZsQj0lqX3m0RRzRt+vu
o5XRHumkf8JoJnA2ildnJVcp92Nyp7Ppx4VJ7JzI7fam3KxAo8uYxKQwRAJtDMQf
M6gNeqXjtVys5XiKEnfabZqKEPhIh+h4ozOFBDzEG8XrcwKIcKX9zkAkEiR02/3M
1rSi8R9lpOlRhyH0TmTMWHJZda+i6OCVDG72MlwfkBGDuH9ErzTFFxMm30AOTBzX
fUfe5ORx9UZ9QgjVv5d/LGf7SUUv3cP6JSeG7lpGDXNjMiNom0Arz8pPIpkkHdtd
WDJ9JLR9bp+JYzj3tOAgVCqcsyTUOrKLlHLOWYtKV+QoRtU+hFTb7ciQhnDJZ7aM
UYPmOIUajLNQiz3DssmXH2O6L2je+npLcSIn3aidpX+ItN40RHlaSPADKoh6R5hH
cqybQGh2keqeX/mzOVhd2ht1ZfB25iuWLIETLOwniUfzVh4vw+DY/LUT5aTEd66n
m8zYC2/RGROpzur2N3/fPIu/QjonK/4wMy+KH5UDLWHEfWQra4ok6auWo+YjP6Aw
ZjL7QF5gMnY5zSjytnJeVs/KIFmu3U9VFtIcoHbJWXAOMCChD/wp8CX+E/G6Ytoa
GJ5yo+msYajW6CzA1oOKAk4hs5V502DasVNz0VDU/tz+53+9c3oGSzOJHKoMrq+u
uvYy8a3Gt8mA47+KtcYd0HgtommWvACXL0LGGFrRASjclRv2mHcgc4Ji2D/FUThC
qpDEdGruE7BJ0qCdmdoXziikvTtx5ZB/rqKw6RFa3XKPWJH5vd8vYBsw7obwfoCt
WY6NXEa79m/RZon+l+/o8qlTJbF3SK9egCqf2Z3zpj7SCi0qTB9FHtpZwF/f69o9
FJbeQILH62FP7zoR8cZmc7mveWSG7e98Snm9LCmhXPrIKkLIURXz7NeBTH2V4RTm
xa5EUfdgkoozzuwvEV4loMhl5cJeyTLhKK91wse/Jv3R+kk89nh94V0MAAYZnJj5
EnaT62yAyFNUcmTqCFPel58OefrRMRuS5TH+RsjAQwjMuV7lM1cjO8n3eSbswghB
fuSGfIxl7v19m/apGzA6GyF9gr3s5YTn/3RB4483KmYD/tVbeRMWBQuP1UOux75U
71gUIImLWGASWnJVPYcGEs0e+OS8bDeWnampAVSNAO7uvAbzy59Sj+IHFPP6/Uro
7nSobccm31+/4kosnIFRYrRFJN7i5sORcnCuMhRov4KhzzFI7HngJNVoOUtflR+1
YyKBIhR4TAjbdUMLwJtFhH+GthvisEOVpOAFAVeCGCjJDsLQ09Dkk75od5ex4VIe
rPw5TFrF9E0SRJEJNNfO0VzV+asppgMjq7SkI7Td/ngwmH8bdy+iRYp4WpQplWk2
3AOWmYtv15jDhq/vh3dyz/Unosh1PjmK2KsoVYF1zpOpWQFV6YyFDZqzYCB1ND8m
lFnqJwsRYllv5d9XG7Al/DtbTrZNZgnF/FtmocEN/oaS/OrMkoQpVv65uP/JF+AU
ekVyyIQuEy7yP6KFPd6NU771JITxa84Lo9w0hdRL1x2azm7KYCrTvSWeOKkVIskn
tjuqAN62BXWe7KjAy701UtFUqi41/93z0aa6PhVr8Dn83JUgtnIpsXWMi10vomVx
B0iz6G0bX936yfXkl6C4VIabfcW/aYmXrqgfE40QjmmGy1F4WQBjQHEnhNnSy1GD
fZCCsSzsV2c6BYqw0Smzp00GDp3Yd4uVFLRinJ0nN1Kxa8GlrmySeXhJQSqNyBoE
eQXh051DxnqbBi86REfS5ve/2JYkj9EUrRAqELwh4GSUHFITckhSPDwHlcHKGdjc
kQmLQg4zigfQI4PoLWrLF4aRb5WgROdWqh/XFzZtf/m0Fg2auBbrIQiSYP/WZX4r
gzErcMxw1K2EXxd2r9isLQ2JeuCSl0H/l0RJc1EqxH5IBZ++bWoCYF3LZo9PO5Tz
NbIOkXL+d5I92OdM91IF8hC5I8PHZyVCy0bE4Kv84k7VdMUJPK4rWi15gHntvwSN
C51+HQdWBXsfNMWLDJruTAyf5TTW7djjXQPrHCpFmjSSYjpVwpm70njWJM/oZ8cA
w1iEaTC/Jrs3vBrenH7Oon9dsrNKDbmXsNS+U+eGVp5RW6gDBzvPwbaayAT0OtSU
n7ic3sLATeG/OkZXzozgrU/ALGKwrsPQ0eFtmWylpPdXBVDrN4e4V9MWHXqengpz
1J8i5Dv6htAXw6tHfBlLyl7EknR7qklfnbkqfl7n1IoOWmNHP0pM/W+kmsIZ+e3G
MD1S3HgoFf1wFq/STKnQs+hcj7Wba5ytMkM69CUojybm/7sVS4NEKZq7eTbjQBAz
W8SXL3/kMrS5x2J0lHo1/BPfGo4elSWD+iL/erD3yTfqLaK+IxZDcEBhCxSqGJuS
nFW0hYMACBLzaonF/1WlImZ+JCMBg+TsC/vK20+TxsIA0a7Tmduig+UIZ8W9fpbO
axRkvSmmQNeK5LaTVN85PWePP9E1Uy+Uh2+Gg8zeaqMDjASJrdL8FPmmK+teQ/oC
uZ2xMUFyRdnsZwOk27ylaFb0bC1jzAXDSYmJt1DZWy+D5hhn6sNydXxvMvexy3AP
KoLDRQfjzg1JTDvPZ1mVpam/1ldgsNHG598RJlkRu7fmzg49Cput+OBb/8ofHmrG
zyFjO/p8z2N3I2+YPllE9s5HmNuMmXFNAtPhgNXMdd7NXv3JbcfNyNnmKtNR+Wbl
OBcsdF2hnzNw/UP+J7K/VgAT5gQ6V4u8kvdsCWyrysJMSYOa9S4IS1pT31GXhnS3
Ao/xZ4uaGUvh9WiCv0p0tx1vHoHfTBvqhhpFrzUSl1nivaZvPUWZA/py3Hay9j0D
MaCm77GnSY0OYdvXE1Mf4VHhjpejDAyqWCGe9zlqOPR7krwo773987q/QJtFQh/4
GlyTW+nNSto2eqE4O8vu40xfgri/JPHObTO+3nU8hY3m5sCkA7L58GkPR6ZZ6Wi/
VbH0kOKH3Wc4Tf1JwkT/nL/k6CEqmlD8rbGgRBm0qsfjf4lIoR+G0MU4+XxVXDBp
Vtm8kaBLinr6cb59tiTsmbMIvxlpNIa4/GcQJqwZFt1HTxDCcKSSTVqCBK71xtix
/tk6OYqJsL9njPrLtPOTqdigIgFlCijDVeZOx9ksgdyB46vxWQO1Wk7oMRzWiQ2g
P+WMYWGw5jbHVaK1q7aV5YfJG/6vCO99Srnvt7QNR0SP2X1soN8Jsfp8RH/Ah7w2
fjpBrPIgCLfDY1hym7d10Eymw476jMSnE8KBn9dk+kaFAorr5ihEbWWdXySUPliW
9LWYTslmFslwrGjj+PVRPBONAUVCsj39MkL20x2V7efB+LWB2nFF/8k7JFRVC97W
f+OCVcliRnCfslhtrSArFqJckgFr9uDIWDMm5gU3qUtzbNHlKc/Nncn3+TGXbCk6
rMYHBLJhSe0IWRJYH+UbxW59hh3fgF7096SdrwdWbnbqHX4Fq+Lls4JMCRUivf9a
99mgDPzNKL5zGTgimyuC2y+iLKtRHOgXry3FQAKxkXLQp8ISxOo6P0OVPOWDadux
M/+ojLF3eY6tD4RMzqY1aftEuRL+GCOm2dcKEwTVa0pZBrnsltbxHlcon27LnBdF
9MLE+u9/fivVL099Fma9L0bhPrdduj9JZSePo06vExC0pP8cAYZygqggNe3pYaCw
/jUZWcHygR5QtBEkCh3MLaBHM0dzf4k6zaB7Uy/PieyPcLM1OjORW0yH5u2R7usp
+lJJXmeAxVB+3D339V+FwwxQkM89+nxpI6XBg/xEq/y/FhGzvt9zIK58Fur4Q+aa
+2d3lJz55CZmZk1YOiq+rUFOLtD46CIWwfLP8uLHygx0tRGE7d0C07A6m9+VEqnT
FsrNdy3Any1Smc3RxfeS4KuVmLdShVxp7Z36OK+nhE2zW1MfhhyZCLWYxX+2DuMj
JHEsqgUBIl5XULWQKOykpxAtyPTxQM3+5MVXS2E0MqlFQlO8/ZIr5IuEOW8/fJX5
5gVm5YlspexUi+HmdyQZd/vcTBF3DV5p6ZRFHXB0W4Fgsfw3Es1BNYHbu4bV0rwm
obf81wZyR+O68OVDfnqpWEignpuAfzfd1g90v3Z6jRL5vAqXGj8DHJTd107OzWyD
CkglBR6eUp99iuN5eK+boLFaRzs/a4JUpC09BEnAt3sYfGeNR2Q+DJMIyFqg9beS
+6fLBffHQfKTmfHdH2YvpjKwisW/detXLU2Ra9WRSjz5tCzP/W+6CpUphml3Tjzi
YoMOiVPR6WYt2g8cjoOrd1R8cgy2aLkkb7mtYDrwPbbm77IqeshACiv/Ux2wJJR1
pyCTym5b8WsKN/gS6oC1YgD6ww7X7u1feeUDZmDNjtbxKnrHJSdWA82zjm+xzM1T
WRgjogcG9XKvsknE5mlahlpokvhV0fpFhIPzfzJ8WeGU37Un0cjzSu07oG3zLpbw
KB8Qqzt754IT3FQv5vDUj5Nozz+8/4GTyV3Q2c8bYDHGy1DPRpSbKzZBKxoiLRb2
qjwLh+2t19La1LhoQ7TunglNvf6RpJa8ep5fxCNtbZQDVcapHppDn6z0Cr/IBpfc
+PBIjiXWSTQ1R++65+x3kpI2ZsJuTiJh69A2fEbTBJ2a5KDgIk5FrtEdqtfQaOW/
mCWY1JORu15m0+fK+xKWKtDc6vmo2cqIgZd/gj46Z1H6UvmK1QKcrLGx2MQOwWKa
v+eS0FASFYO1/955SwJyJQeGLwV6J/2K7bzcgP5HNtsc3HdgYRB/xNBN8V/Lj5F2
kuMRI6EZFLDV6n2LEzclnDmgsPb3GT7hV6AJm9tLAzLWZgD/AxCpZ2ggaHoj2wXw
lSwxD0yz5nRmc8dMV/0sxHOaN/jlFzorOUL9q44smgwQy5I+uqYNxgmqdK8wCXno
C5/W0O99f0oN2Z1e5ATIe4q5binuxrEO7F5UJhYO6LwuogHHEZI7xYUBuSvTYfws
z657ZBsgCnke89wuacqjyYZAI6gnzp0AeNpPpaafswJ/HEO7OZGQRjTxCK8IGP9k
byy0D2ubBP9/eV3FebPub0HTlApO16CBHKSqigQoMTuOVNqFYDd2DtLScQYT+blP
O0/MdWWPH10Q6OV73fUVZCU2Ef16e0/GWYXN+aTzKpifW7t0ofdGeeffG7NS0IiK
7dbgJiQC0uw65qRfbUPqNDu6f/uvCl88EjwpUN772WKpX11aInRpJYzXpgesj8by
PhPNaEQqOk7iIjWt9O1LepaF2dCWnfgmEw3NBM2xV5oLxQdWYCS1+r0NtgAKCnad
TqV2U3wQpvARTQLwpG9GYhgywGUXInhiumA+cjOG+QzAeiM7VM1EUI2MJuSptu59
T1vEbs5s9JmArTMhWggANwQ3vooER4QstoUfr/AM+E72ToOYTipCOaqWkzvzB0oX
bWu1bybBqKfwcUOR/9RoBSBPMJQjBtxNsqfVPEtXGPaLMIQpOYQsSj5UcXzDGyDV
Yh/TfHWcpovu8O+TMNHXHgRClznt8WP3grBtBpeD+cUqgyDYppfdS+ZAIJeqUeUw
tSrUOG9PlqmfH5ylj7gKZwneFjKHgoqhRlR6zbdbgs/bSHIRoM7woczdRBtqni9u
UXTLn5vRN5KxyGRowWpuaU18as/+1LvYBUMNWXXqjQ072Yfcm6GEIzUQw1k9j9ra
d7Y8FMY1BOIwXugBcbSJX1xoXNHgToQ8tnFRQPxGTj2VS4oLOjzmAvi3E8T5RTaJ
Gty/ED1OCOQkxpnHpqGPnGlpM/7y3yqsDy9uSxA6RyC44LCJa5IRpH8QtKTk71PY
gau7Pnth1Vpr3oHf4x4HGY/vQyP3tSskGbFW5zlORKhaxh5RCNDqDvSJpWTphuld
xk9Ml7zxwCZma5/d8kmloE4gTCLM0mbs2szrO2sF3jg0ynwkimA2YoVW/kAHkCCc
EcCoio8Qrl9D4Q6s31SFKJxymdNwTR2y+3qFdRR3omrGzQV+c+09ama6M78D5XRB
BqI0wWfUcZ+lOUFVagyelyQTtKOiuhOGh4Lrz5uR54JSacTD8GNCC43M6TyNAWHO
SAgt3gLuQV8vtviS+2r3ECGG4z8JY1DVBlTcer/UW7QtNC9Ie66HOmzBpS7NotSj
LKxUNy9vRkrPdrG0O5hAbhXLvvU48Bpw7baYRKcc7ghJc4hoXAiJr1IVSSG9xu6+
I4FLvINiT1AeRsUJTOQrBTNRwet6Z3awcFSoT9RlnBY9Gmf65oaUXEkr8KGN5b4b
PMX50munUH9Hz9fZPucRFbia5bA3EhUeoZTs92xM1nAToLvhSe8xWroCENUP1qIJ
OAfF34EiQUiZQM0StOwpeSIQ9qUAGWxmGB4TqLD/BuELti/JaLu40oIcBfkaZUGi
9MvRQYbtvuRXvh57eNxouuxH3tWwkkcPdNKFcNGNgjuUfIXd9GEC7X98rMun/xoM
Wj3EVUpFu2n27qRUg5ApbdUYu85Ub0Hsa4wzhM2oBzoBMD/EcEalY9YLcN74qwm0
rbcICrSg8Jv94t2a1wkMuBfGDrBvfzr1ySAmfuqP0T8iVfKCHMYIrMBdOANkA7fJ
zhnK2YM+qL8CqzImqvL00o31/TW+Aa7yfw3dG/Q+l0Ifkem8oyZcF/kby3GLgjZK
ZBLMU94zVQEk5Ky24h8aq7Jnm4DozxBP8fEqUxqzGg9hSUWJ5lSbmVjgN9Iac/zD
l3fXVa8u/lFielEMZ1tZ36+KAf/HsF0N6To57AXGuq0cXCkYEVfaqPkDyadrzQF8
RaypD3SuRfYB6sjsF1f2IdSZOb1qHbzdS+TZEsXJDbShhY5BMKoFvm48gzytRlHr
j/1mHVVeGEh1ZecWJgyzW7vC3AXfslnDt61VHeZ6ErCfUbiA4QcfRzfdclYxu29e
HB56rzTaacMEbxKgtDPSBLdQkOeoDcLwirnqALAcmTsDBbrkRGFymkMFZBtCQucM
/k65iaQFPoBeJoxLL0A47FlXlABLzV8Es4D/2MG37zTU0enwqjacKeePSyqvi+ar
7FA1pK7Ts3t+SwkYe6BdlZeKwK1qWUe1yVfLDyx6m9Unh0QIT4CO1vR2ym8UbKrp
8Ck3ZhvfaZvSX0G84fc1doa5QiCRRrzjCwWH+pzdZQTUEyB6w4tWndd3Ru0Z3FgX
uGAPQqMwLJtQhJKhfLUnLZtb0huCzsjS+zqIuun2nSbXcaUHJDyMJlKwNXYs6O/g
Zzj7pHagU97WNmOT2EzrAkbYlXzY/XHTxw7+4YeKj/0iVKuDwsdBrav1tg+NrUKz
I0RTA2q6i15A+doLRnxUFkzgd1E08FaW8iRH7kg0T5QbvuLh5vLgjxByj4+JjKvP
We6rrmeLBY08AFD0xQE/KJPxfjuA5vfHpGSDseGq4gKYsjnas8HM340b4CwGMWJu
fq+YDlvsAXUvFtJG5gbmDItLkVHrj63qn0oEq9zhVJtUgsYjJr8advxRjLHWuwol
hDz1KFKb76MMerj48fTgL7Pt4/FYq7bI7gUp9rDx+4qgZdfYWo8E+1ZfKGUtqjTZ
JaiCdnvA5Rw2vJ9y64eLgdu1s+5G0ODi9RPORFGCP5OzD0VuZ4TkOtsB0SOkXxmg
cyBKEjAKy3rBMSGJmOiIw+j93ZwKeSTxl7p8k7PtoeNHM3GN0EMM0h4Ut1ieFI57
wwWVmNJcAOChDr1dbC9Udyx0T8+ioOQ5pnVTccwFa1RJISmvWKAjInTCQsfiUK1u
wzgn5oz3m3KYnoDmfCj8HqlKaqJYKUpgu+HJzol0SVt/5t1v7VJRhsuRgZZLwHgW
El4iw8C3JgRpwZxq5mBXIZF42jinjIOFpy8Jz7233C895hwdIsNiiUhUUT6wKsXH
Gy9j2VqxMCT83Qeqr+ULc5kfA8hyv48JNS1GXveZ17x4/wO/4OWqqWLT64oHIPAp
6ZcBT8ifDOnik05fuSxLa21kYD0M1tYGqcQQm+9L4TZ0nCIX5u93prNmtsqyc8Ds
ARtwps3oFP4JZhjYIxJF5JdK+1VPYBOW8XMREOO4VA2Se8hloYkRgSNJHfQStrMx
CtL/mkDdi0hRM/YzJbtxopZohoXqxq3jlJYF9p946Pjr9dkYfH3mX5ZcdSFP64+S
yDDvOi5lZVHINwHtqIdRaAWJhoF8X9Iqwkiau1uPxElyWs8ssageBfKvE4N0SUKj
6cwix75RWC9GYpHMChrwd53hDkmxsm3bWd1a7LCd7nQh1sRRJXzOAPZ9atkgtTs8
4HprJmckFqFqRVDXCmaapiBQ1alCBn3IHZZifhqUPwAojNBGXRIyTSbEh7RJjYY8
qnFwOGZTCtX+cIn5bz9TgXWQ3zzxPfmwA69bSmqFdYALRvGlPYABVBL/YZl3Wm20
IcpsMzoBbEDsb0YmrWlOmLER4D8lCOdnchIMItpPKqST3N/Em2s4LIGwabfnwPLC
lp+m4sMk7AmK+BK1zWtDWJKSDw+uMEwn/FYbWt5S/BunFz6f4SF+Oo/wFatLF+Z4
xQQ1/SWx1ZW2MdfP6tHaz29j58nHLepPZ6e/hy2gCj0Ef+g6n3nid0g37YrQFa6Y
Wl7Dh9Wk2LonjcnhOZX1Wu82JbJk5X5Bq34nBbKHOBxUdhFIi9ma8ekZ2OplKtkQ
OufdXBBz0KaEFfuQrUkOD44rcyYlcGgZ74g7KBwj1Ff/KyaEtmH8s2U5RcvqRn9L
nMJVoPgCbwJ8gC8B1xD4Ikwchd6Td1ZtBVTnj69fAIVn2ZMh9EennpNzDALZqTG0
2rqXlDAZxCrbe0XinoSn+QvL61QlllXFYGOxPLhTCfMd5Xch6pCCxx6GiPd4l6Bc
msYGkmUaz6liXOrEU20e84kJ5tVBELnEZEfWQ2H6aS0nkDbk+LeNARC+nu7A7suj
FByDyDF+ENkcU99P30RjJTm+c948CmS9cRtvLw4uDYAcqW9H87d6ftL+EpB6Msh6
/9lF1tWfQjSoRSDLFi25IOqmmfjNy7Zxoy0G2NX/RsmiD4HhlU/d8IU5bzzpITQ7
C8LsiFe3u/RQW5BsrRG+wEsABq3LoRC2jBDtjioXAzA4FuqGCj9C7tBDxDn+yC7y
Ly8W91Ih1PrekhIfIqmURry88R/DP5bJ2gxX1GsbYrxdMzCDaXjNx1cEGvRdL3tD
ISPXZnwMJEPA0/mJkBIPjqQ0ZIiUGnelRnABhtmvrivUcz53dBj8M6WZE5IVh+oh
5CpguQAVlwSea95C5dIr5oITioOJxYMNYE7fQhNJNtMCRwqlWaxF8wuH+Y2msqxV
6rqvKHgSlpOV5TdVkZw7zw29JdHwlUd8bDA3CcZofiMI+lqkabN8hd+ZAj1XsPCK
fbFbBKmgn6G+HXsB+ei5eWzOyZk6xmbMVsHBlXLNR6UouA8RdJiOCvyRu9xjbMcB
AL+A47ce38xpwEO4ht/w2PMqBuvREB7gGQSiBWFS+gm5JwyMdJADeJ1p0QMLUciW
8UiMV5STPyvw3uDof9rSe/46H29LSDwQ/qVLQEiWc+ZyCPL0qvQCSS/doWEwu8MW
m1Q4++dLm1iRv0i2+XnEk4Gj/czn5Kna4enrIGQre9v31lhfIhFDVCPYp4q9OFyL
FBvb9TSE/T7T4GFqCDs0pgjp6rd89DFxHjWBGS4GiCxGOXYyqh2lYu3ioRmkiYRl
ut8AqzSulY/yQHYEb5Fa38/ya/yHF6eJgsiI+79xHweeEhWHNvYpedQDYEatFG8b
wjpsXCSEFJnwkRPUt5fjwgLCSSF1ETVaFcozOdyCGzc/OARRgFD/ZcgmWQTG+PT9
sKlezYpE/09qf70h74oJ/TxloIDrz1XoqVMXkUgEgOiSIWMw4HykZhchjHbQ88no
zsI7lPoiApMvNlwFlnEFszeeE0IWpdumCaNX0PSfptbfh6Z3QhYlqLK6MDuk64gB
MiVTbSfpH85ypAtEuBtnojaUwHr9oHD0R58iI+w0tTxcNBEy68ZSQG5Ad43gf6KI
MR/xlmSksnfg2ke3jj6Hw8KhoNlFJ2mU0WKbTqELClgPdy60LD4YUsg3dczh4nGJ
kjlc9xDwrEq5C+MXnrsfzTTGTGYqZjkOpCys4v4TL/QeLZQrIyew5o06YHJeIRDH
xoW2PGV9IcrnQmTLMXbUcifsS8msiV0U25v05QzTmxC6PI9gdxBX4A5E1bq0Mcjd
1c7K7Hp7qyaqKIdGpUs3cvMWPBexpNHr2+FSS4wYtWNLc2pJ262RZrHQLB5BX+ph
FwiHkH0Nz/OZ8EQIPtUoLqRMcVCMYXUyYo2YgoDiWHCwnko6y3fDXoXY5xbsTp1S
tgdXyRrcHGsZq8Ur8sRgLxb82nxPaqfrBLE2U/5AvwIPhuuQC4vW7qHUQT1xyN0z
d/+kMYrglXsqSUwQoIJtl8rpKIWJtD1LdnTCHGb9trFyKlGfTxJBEMPUR7EVmyZN
uOgYBRmxxuG77hNu7dCRtsmJBi+kAhDB9r9I+/DgtAXIqRpbld8WXrWuzZQCtkYJ
ma4UN6K8oI2Rf3kGzGlrBLRig1rL6mwd78z8/sb+q17qVz+sf21vx9Vfio8S2g9c
222sV7XW9gZdFlOECWUo4ScvSaX2+0JSDEKE/mbEbz7ogwQ9u2ALHGwpvER/AGXW
Y/lZ4kW1YqvNfV6UDHBFpG0kB0jyISBKPZ4dzK37lJFV3RKWvdnWxSTcbvWQxiIY
VSVoL9gFa/A3CUHQfvDxKM19iV5QP5edOIEF9uV49BabILXN2DhY7nLU3ljEQtZj
1LW0d+AOzazlnfSEugEIb0mepD0Uxc0mznB976oZ/nKSBHggXo21ZCC2dSCjABdJ
+FxpLOwmQLz7y8OitWRmL3BhP0hhxbpzEgtycaQnDx1IcZa7ahhfr7MFRv25gujB
iKRrwVEWyiybwQAXq3izosQtGBvVXRt28CVHVFH8gqqDzuvCAfI8LGJpITTcxPEN
Ya+WXHGGcePdewHMm34P0S0XzsXqds3ShPhFnNiGh4IEgN91gS7NVdd/S+/tDolc
T0zF6GHWuH73XvGFRx3/Q8alIxH1kIb8L1b9v/JdxIU+ALi7FVLZ7BfKEtdww/1L
E5MDpxP7wj+QJkmUkOPpzZWF/zGcrikLKfZEZt4XJyr6NQwzr6gT2VirdEHn8hrX
lIfaE+jsf7dLlKCKKuEKcSAywncywaFM9ERFrn2GZE1oAy54dYsIuQBgNY2g2lwT
a9N72aWExmEAXHCTpWzp2gQ8F7vwfNCQSjzzslrrO4mhDp/mQPE8FQ77fgsxhvve
cWb7I+KsRIpzPzDsHJaRPnkL5cnluuvVSswEYaF9ET99olu+3ueJeZ1KsgLkNx4T
JpNLgareHoDNcIrug/5TSTEJgupnsXp8Cijx0RjoHi3ydc1FoDuulvImcmO7nVBG
YczN0UMhbTh7Od4l4QJduH1IvZbu+5pRb4tYZXxGJPeTrxQj+MHl+mpMWm8P8X0j
95mjTLjhUlnO4jV0LN3J+KoAu5XxDtjpt/cT+y1z3C+S6l/UGP4VvmYY4KtqdXKn
p0caEkVp0qhdAQ40U1eftAFEEqlklP02zzg2qDco6U9OZNlFZwwQuAQhFNj8OtDZ
lHbtP94eRpFaXRk+Z8ywJ819VJEEqyO0cszDu8YKeDf0uJvL67ke8KsBkW//cLb7
7/DLyl57QBtPAiQJVtcfEkCIvcGnhuTmysSMBCUHSnKvf8pDa76274r4lUiBVsg4
oiFNQXNdRZWBWqhMX0gE0yDGFY9mNNoTG49yfQJfhQ42Sx8gAqDgZrq+dlcivQ09
KMQ2k35zZWRbz/z32KTz8/rzsnFpWfF6X/jWNtEcH/ucS2xSamSDeHcm77ZOMEmp
gA2DNwH5W+oW64asT+CtEKTMnLCwBuFNclSX+wr6c/o+SdNIA1NGDYLgEqfgbJi2
cRIbxL2zHG4Sk3fnTrGX+X3bL1/NfaN60JmxHDBMyKZ7Wx+f7ZEPem28SL2Sz5Mo
nCV82aNric9Wz0LuiCxwHspQGaOI/NWLJopBKjbT2R2zcKCa+KrieB4EjDdsXZ8T
U+9tPdStCrlgHkoaPcuSyuL4YfNpw+odk6yqnQuYkShU5V8i6rfAiwdKQ+QdU/jf
3RodZvcEGKBggrfW/FAnvDwJRAq+GhV7A/QdX2XWP1kMkd28zAqb1hVSQhIGQX10
4zL/XEcUkQldFXuGwJI7jbSgObr6/so0p3+wJvAYIt5dBTIjvaPbhAeQD6czEyOJ
EFKv0nHZ1XFpKvH7jtBjZIne/wr08koFqyDcWFwfJM2kDcMaxJEEgI3l9ruaxhUE
awVGMMkApbLqkh3gWpBEjbgY1RaWmKndlHmkDBkEdFOyMrwFf3yBypdAIZrDslSL
Av6JEg9/6wNC4qYpyqvMc/nTxt4qPhaoaVqwfEJVuq54A6SDArUu9HFj53MnyXEb
ACJ9rFJlZE4mFyhE7Tj9cLjPTQR9/lKDyA0clIML1GlbWr+0Kw2KGgfmMF8Ut55D
SesjtJTHKko1wTQ1k8D/hRHdPf8LqTCqP2cJQ8mmkjQE0OdPqEiyTah77F0Hdpkp
2wnQG9jWj/6mkl6+Fzy5LNe2eVsGpMIEGXp4hLU04wks9IU0DXhk+29H/3lQV3bs
7Q/lV1FEkPMTvI1+oOQQ2btEWW7EOZ3vQpmh2vf6tspCkG1/RZx1Zn5fKEyedP0B
7jMGwA/vYUjg7NmcAy0RmrD3H+DinvpcVL92jazi9g2KODxd36jMK8SpAopyFv1T
zIHpNSvTd0BrPZieeSLy7M1kAR86e8Kvth/LKO/n9Xl7JuEGU0t9CFbEE2O6TzCS
fnqHUcL677s/gBpC//F0YeLKpewBP2oZVBTewpAV0+kFRtAeG4nL5m60o7xDEitd
eG9tHJETbmvnRzNa1795elF4j8NszghRGnfC3pTXOK473/U5zfp17C8m1IAbb0Ig
Jtg8+DAoBZNjv01c4BTMkFj/15LMVGplbHiINUVSIcy5JQAVAhGovnFY7wOcIJqC
/xLka9DPN8wOenLR7E8kfZDtRyJAnZBZ7YOWYXP9fhvUEqFhFrf/rPa3+2FkHXEb
IjdOCGcjGEc+SJrxhZET1yghBG8KeeTfCVsSKz8K3PRlieXUCgLdR3TS6Kay3NSb
13vizKA/cjlF/rT5i2ytCE17/Ak6EdWVDzHDLOuIdhR/YZHjP11H/MdM4EhJ43cK
3A2aVdxSJhD7j1hypeLXws+ZxXu6/AqMGjR3az3UHGkm0dTT8GzB1VJYfxuuufPo
xspznCiviloAfD6Sp0pUsdhkNAbBQigSrVnfubaP6VEijH9P7OBHs8+I8bncOGND
24rd3FTZtA0rIjQ1Fqb1AGl4cs7MiK1HvQJTc6VsDFETg9RDpITQ6ji6ePnlvBUs
4QdFD5kBRO86vuxWA7nBBqhL5Be/Kzbni5R9uxFa6sNtFwJrOLCagwyGVoxWZEPa
lF0UZtXM9rlcA03DMA9+X34eVPtzebQiMG4paqo3/yFx9om9XyGk0quxTfkcJdhr
q3fs5llHK6yzfU976vnCnVMOZ6juUF/7IsNt7L84vx+Mx2FYbrns/Z0RZo5gDMcp
YDWR8jxBTMvBx+RMxB7hzfBAeqYtllmU1aOCKk/GNOjQYitUuoYLUdH+UqtiAnq+
jqIPwXrRVG5cgn3GxyZ7KjJi5CqcVpGmeuhMEIVwgNhx9v4pU2KxiqO0Nef0P3tC
1fUwAoX5Kctm9Pv9DbsHsEwtBKsTqcqrZd2V1EBQqam4/0aW6xph+0oqGVqTAjsL
ma9VNZ53jgFV35f2T2g0Sg/u9B9+du/H0GDm9Ft0sBRUTun5vtwZ5evDagTUfA9B
phWCsBbV15HNfMf/sxd2XX5VAlemJvam0Soasf7EnCgJlJg+xV73Gs+5PWJr/r1e
Ip5kdwJ//HhXuITtPZ/XAhRdvXKvhhjzIbObI2yP4d70YNC0JMLBv0t0RJIsLhdi
/3+/ibkWhOD6hffFSRM87zrwpdPO6bAI3oBaneGHcFT4wVHAD3xZBlZbgIb85oSB
VHcTjYwmhdnlRv+AyB6RneoXHEhGgkBvoI+pTkRCDnsXVrggFvxsOIsUnt42RSVl
5TvRU4NH2TRB7gnXTt7UUlyjz3eKu+X5v5unQS/OdyA5AetrWkQvA/iRCrExx938
XCu6AA9wNDHxRWg5q3ooY5BCtBSOrciKMY9Stxum9tFyWLs3USc55yeVhPmSJoPf
ZR3TTwTkawLnNtdrdVlXbNQW0dXmCbjUyLK2T83yAQaOsWXn4XTJ2Tz8j6HYutLT
a2fKnhXcPm+rcaXOw2pEcOIfwSTXjA4IpO46pHLPQGIzHwLcFWFqnJaZTo66zOuv
x4We4YeLX8X6saPf2Y9G1wBbXbnwXw7lE8/ZLgV80gdvJW5PI70ctIj+uOsHLfjJ
0DiewyGLZXHT1rgirVoPKo5y1M1HFPV65D8QhK+FShcGlntnlasjYsSE9P8DzP7U
vPQtSBEhHVn0kfIVfMzJYyAzJnwT0VSib6a1hEE0MkOy7YPaGjx919sezZjFEMZQ
ZLszSTMhVBupoyvSEI3EZfmDEqJpmb9OKtc7WxufSbM+uyk0guSntq8nrHXkoDju
qwU+SMrS8cCakhoQOonrElzK1xdSwm5a34I1nq+ynwdRCrloFrEAN0+OSnIApJA6
xakoBdF035Sl8JrBvMtYJqq2GDI7KxWm3sAtxMznnM8l+1da88M9QosONI/KeZ2J
oGJsUN6/dSQcmePem09Og4brBdq99COEFXZvjfHvPXd2Xc1sBWuohNs3KQreQv76
XHnlwa5HmWDQxQsGBDakLqxV3n+zo0ixHvBMTlzihJoAj4UWYSPhmsTUkcx+xxCi
8xtQ6lK8OMKvD7uUp2dm93gE9AZVRJadoKbwvCwwdgDqEaK6aIHLylKAWKeDAchW
9UR7wkCiHOoyCQmRNmWlBf3qrSzk1de9W5M8L7QVsGSG4KeA7Zcy4aoS7mxI1DIn
n7GLu00gxUfBbC75MdYFzdFh1/agRfT8QAy8epAIuA0aYuL4LhwOGB2KS+bRaTks
FQCrYyX3RZvquP/KPAvSlhRK3Rjv9gz5KoUBxzHyRgYrS8eecgElQE4b8RT42l8I
D7DLGfoAGl92YzsWz94rAEyuYXb6V02Hgox9fAdE4/p9Ql1UJ2ZJN9E4WzzET+Q3
yFhRHRpNdLAO/4BSRszrM1NiS/Jkah1k88Y+uzFi1+tEyC9sOPM0rsOIlavEN3ZV
u3MOh7geAXsmUKmW7/pnnCXMQSjuqDviIP71ckPWc42SmFCuMnC8zSj6uzaLspx1
dWRpbiGbd5RCr6nWNHNAqM/5L+uN2Vi0I/YWuMi+zpkGb9axUkS09PytvkuPPVY2
jKr+sNxtXfztsrux5fbhtpyIkbZEjKRDSVcs8YxxaYrD8P1udNJ7ETp7Ab+MpVTn
KU/K9aX8WqDWmghatq+N2m7OLjnDVIoo2PM4ezkgUexCrDJAyBwn7wDEB3oEBLTE
++YiUj4W+MxnlAZRZAsO7PjDWnNcmBLjDyJGfbxM1dk2U0GBn3/qLDPKcGauxEbY
s0BkDGVuo5TpUMi0yx1aAUfZaq4f0Ks4gdyssxxm62WvBGASSOIxMyV6aFog+itk
4O2xN8jeYIXfsw0ltXqEerwTFFBal/UH1rSCRZsvNCxkpZvsla8ZYqTX8ugeRlf8
XBPUbUmcPIGv3hxQRBOZe4s9e1nrJiSDVxvKZ1mrxAgBnuBXX3QhsFdWznl57m11
97TkHaqZoYNs6oJMQM+XSboT0i0/9o9z8wBF2FMHlmgRv50OzSm8YpaYvleJWfxa
1yxyakBwCeLz7D4li9j1eI6aXPNg3idVLmA1/SYmUshW1dhRsxNL56KJhBz64e7e
69HklFELXJw4e5oGp8J3z7oM2hXkrrYpD5QIhmke3aBLuBJq2Al6xmGPKz5FxKaX
L0BkaA/3cdWTlJUYvkGIRzqYYGRXov6xAGO1eyKgLtEEk8PToubF1vGkHIfDTog2
dWgYbe/Tb2qXC7p7mlRGBDMhxdbEi0hRetE5UtDqZw6gMhOTl68i+ozXmRomlkBg
ykpEGcKLraoGTrkvE0CLY88LMtuSFfyYjY3kLf1ggWWz+Btohz4MfdL71xcqzosa
THY8Pk1C+B2ovaF/M1kBDiZlrY95sp8E6pCLnSuduzQsAiIPk/3nDy0udeQmsbl6
ztsCLm+d2VJvG9gK4ZYHR7eDCGI0NkdK9gbkfSPWNiJ317DrWk+3heL1C3h2FzN1
5FqSH5Pftsve94rqNPVQmjTXWyGZspGtr2mZcixA9BZ4gVFTYobKSWcavfujjdei
aYUoh8+6gj8Ne+v27ztMidWfLMgHLSkd8OVEatIOCRG15QHe/nMQFwd9HA+Kdug8
Z4kxzQVEBCrKhgUpZ+7t5O6rhk3x/9+EowP4F/IBf/MCHctPyMkzacmZTzAIceN8
wsdrbiWitufAGRsz9vFPR17vNMitlWi3AI2bCWeF6AgNxOcGQ9lLqQzQG3S2G44h
XBjU+bgLpk4r7a5OPmvKx43V8lbl+Wp/R9hUvykw7hbibElCSoUIn8R/pbgARmAv
eHYPVJHrJrQzJjfIt/R8xTGqHW0AJSlxFzwSG9gmeeFw53hVNbwEVRk1YJ0neuB4
zp92k1YwmktNA/BtrlXnPmcIODb6C7pLeHy8fq7U6WTiQihSTy3YFs1iMZ7gGMFJ
QMK1RdFJxR3lk2bnR9YCxazW/xMPzCJ0lZxxBBMcF8HmF/Xk6ox/kLbn/2U2Zpti
nhwL5euZbdPW0KEAZ7SJ+1cr85MhDbuZkzNtWqwqNDy5F992vD69IKisYnUgwDcs
GcFJCXh7TSBagdjIGBtM0uYv/qKwfHzWzfuE+gjF3C8zPnxKrWZYich+zb1TlZCB
sMbISEslmwzqlsqFcGCt0/5JKrPTrDlLl5ps2WqSP0QyE/xx3U4+KQZD+ifxQTWM
a6v5DBuEOMvRI29CXXS+x6lEXRkqStGYT9Egh1xllQ6ztrzTybFOSK2FVE442lQr
RXG3MFuVhomTvfvTJrgNEDdbI7XeQ8KcpsoC7N6rU49HsU8boJ0pESWqwbyUPFEf
1mf3CwWrr8ZaDu5cW2dDRi4u+pFe/r61IVrboSESBC8BypsI3jqL3cgl5CmIxmMS
SmC0ZjqJxlCjp+0OOEbqg9og6/YvbW1npJHGx+DWJ60FRS3Ms/QCcSC0ftNWNiFJ
c2isqClhhbH8yB6oedkWiMwI23m4q8U7PtwJGXJ2fVUjvIm9Op8SoDB11JcrYacD
q+ySwVDTozse+8Xe42SyxpemXDrSYAT3zQ4/C/7QfOMGh4948g3OLvioMLHoAjA3
h00JSDih4Wp0EHdWx8iNJP77+Nhj1P5q8npqe01YODOpo0wbw4Hwjni5eryrnm6l
ehIYo/W2UR1heYREG10RrpzaGH3v7Iv5uv3V4OJTxqlMgVsQPaSej6+rpUKbVhr8
maiF8T4urJ0u86TxVe3nmXzE8jhRkxp7x8+zm32J2R2j5EzY50Aufq3ANSruRoLx
t9IOtNBTduiF5hH4rfKrmVdvvaGvuXgZVDn4HylkTDPXMh7NWBVL0ZTmF3oLoCiW
7QKTa+deKdKCVI5y+B/olFoatY5kSwAYqbJtwjwqPlrmGlIraMFQ3uN4MFR1vqAG
HLqbfH+fK4wBKeXY6Aj/9B5/prGWNaVJpJbFCto7+FzB64VGANsC6wAgJtOwlBhT
dyh2QXsF0a4QMahjTnhDDFOQIxDtELRVtSW2jMQ7rBEZjWrK3mYZdBIjdVGd1QnJ
Na6B80TngqHk43AvMvnfJIdDETi2IdB5gB5bbIBbM3HElBv/TClnlth5E5WhqklO
ghic4tjKeu6magHsEj5S3wQvsI7klgsPpDyG7xebamfg2/Jgwxeddl3BKSZ+L+vE
h14B9Sr1deIDrTg8sD+1f1ujKj4YktJEoDnNSkrtL5k324QcDcYlOONo1Prv7MEr
1Gf0BXC/7gnFU8Q4WobqBZYjQqBjadOeLN37Q6TW1OGUoZMHhCOapbkjBE6rxh33
KExEha4RMWmb2bpDy94pCCvbyBzj6hh6xTmz6FxFm1ZqsCQEz81CVx95/tNH5UfO
Wt3fgZ3XZXslIoDgAFo0UXvs39V/LbwkCJGTHbI1lLP7hu9Y9sV5F+6B+leump7/
loaLC3JnJ3kAVyzZ9g0NAWTL408IrqxKOWyqueOlaKJnaMUO6/jKP435W2MmNY+j
ba8ELyswoM1AFYYuPHwLr5T4XapMJfkNZ7zEN2/p3SrAlXFA/j5m4eLb7FJGeK6Q
kZLWjQbOwN0uuFn+ikJ9Sk0ZmC2AEZJymlitsxNpAhVdqybsiycZNOjCShremRo0
G1U5kI+2hihGR9QnRCTQmkDzm4JMYMn6lVu2zLwDE2GWrwnIE9AFY8zmm5vF+3ce
ibLoisdS29xfzIqJiH9CC3O3s+pwwFzRt+SgE9ZCeRZi8F93ZY8CONaYmcMeuzXt
JbdbzhR0D7o3ygoTegYBVUJD6aqdq+xvKN9cqwASGpbpoxei5LcI81fwyyqBC1iN
qOL0Rf5Z3lmc1pRcWe4mTZejuD31aMjDIlbXerfIzgWvbOPtC3Mh7WiEoT2k5ee5
Jl/NpNd3uT1h90nIjC51X+uZVJBjbqzn+tYN4QSQDvPNqCGeDAzY1U6+3gKXNMVb
K6fYSBvrfK+E004mG5SNlJj0Z6OrZTfBvzNC/isnrVmw3SQVexm12Aa1ssRk0SLK
221htqZ0D8KM9PvDN8a0vzjni5cgPxIJA02ZcbIB+AGNbkZci+vAjm2UTCTi2nu3
MbWo2XBsssryXJgskC40rdH8TuaIKY9ITrU7WdmS3GmunswUUfwIEqlrQHpCAHIO
cZbQd8LKPnv4gnFHpFr04RcLr8F2cetaXQAJdvE5Ju+wHhX2LOqFIrjyWXtmk0YK
AhIB4ocOFeN+We3WF/tT5dk5DFCbsSzov0bh+jLuXjPfmdX8rPU1w01Tw186DhPd
lW5XC8tYIu8+Kq5vYQCflKYgHw7HRP9SnKKonN2xO8H4deaBczG63mh8IfXHE0Oa
1xvmp5qstwfA7qhMHN2OpAHin5G6Nc7DzIjjcro8Ln0ZHwYhQHdIa0awMHx049Fz
thfO0qot18zuhzxy11PODNJao1UTT4aywx4zvofX7Lh55mkjrspHsMMoWr1edkco
e4UMfbwv2BQU6g2eyM77oyRrhyvEDUNQ9DSPrMF9hoSj+bbsvTxf2dDfnkXw8dl5
p255qmvdKgUOxcH/ZQcCqTM6OJylFLGBFEaCWNohHRRw9UPiIcJU3zGGJ7UYh2fA
VmqKggY1gk/sHoU8Bck068JTvTE1uYKGxj0EEnyKIeC6VWxw2OUXmAGIdGXhElX3
kE+sbOf4yX85pKbUfZmgmCo5sXfERsQSClgsStlgk4UiEbfR/L+uEGAKn2kRZjcE
e9s0nXWO4k5LO+L2Zpd0AijfJu3Tqfznbk9a7mF3YIDhPI8zqJXiXDhkLfWWOAhC
Wm+smtmA0CP1BEawRIJt8e+nFwuqkCecwlG8ia8cDBP8qtO0PSSwcdofEHTTCrXI
l1F+PDZiFz+eB2lEyCRkLTZJ3d4mBimHPAXrGPTBJnzk7HxXnhDnK1wcxO+8F2fT
lMFtktDB+7Okov3UtiKF9zHOZ73Ze/whsz5L+QUeIKnzdIiPoWw0tVQR5PTWlo6D
IaeCgOjkcaV8NWDIJIUrvdWQBCEPYsANVwOnPfMbceF5niHlqv2LEcGBbbqQlVd/
BxwR0ttOlh7KM9AZanx8YBpKGgGeiYFcq2W67Ekjvj0k0a/APAod1Hqq1LVZNLsJ
to5RbWLzXSZUmR+4/teD93U+Ouuq/yyi9fRBTg8lbf73k1lFEMKO7hPiLDTTNrRI
+bRgejoJW7GBliuOAQbl4KP8hX4EvkjC5LiIGWhnb6p3Uh0NeclPWf4NZEH72zAR
sKUmaK8GkhUASPKMUNjg1O+bIQmRKiwQAjCxwedwtIw8Zme/QoZRO8t86ErY08Vu
ppKNo9pguaj4sDbKvXhsI8EzrUi0U4+uKuQG5YlE3mllHwGL5V6PIZE3388Ef/SS
J+E3uZRtuQz1duCBHNT++JjdrHN6RRjVdIdrqAkxpEA8OnRO2DugE1NiyDGiK2G4
PWFCMJN2ZfG2f4a2Yrkc/pQ1kOQglGcpQEPT2d35xWE7HEIcRFbQKqtMwTBVz9KW
TDyzzf/eFqjozadb9WjS0RDwCalBykR05mGhLYD1XtLp/Y3sVYF8TrlFtyXSfc3w
QQjKkcUWHzGch64jhGnDP/hghSJfzxYRF3IHBjro4MwQAqvr5tw/GcrFck3RCpt9
M2D9Db/F+D8BURiXqAoVG7tOySjAFQzwBmTHvxiVsGLNJJGJ8ODq3aL2jsLplvYv
UfZ0Kk2JMmwzD5QUqdEdGJQkr1EWm7EoUqRNFMq/HwKAheqIM8oAzlSXWO7FCvwu
1XKQL4vV0iT95761VaU/nNiUUBUhRAW9TyY4+AGMXuwHeoBV+GpUc0Zwm/Jh9SgV
M933Ohrh/mh7LuJeK3OU4nARJbgDfCgOtampYfqBlrZHpWaGQ4qIIIZfOGRrSU8z
U5PWgiqUKlj3hxUKyxgDQoJGDBVwChUy2rZ7JrrEv3nkSn3coLkj1X+4THqrX9c2
05GSc5p8y7KWoPCl+165MD1QbJcoBhs/B/H9i39h3LFsYVWt9n5+v2bR/ofHQqyR
lYn4Mlmqae41vHxGG1p7GZChW8kW0mGslX+C3rvvmet3Pa8/L/JApHkGrcYutmJS
vo19rsXwRf+TUCdyck9U4JvFalGhoNDzhYhAs2twnfkxusLEQ516tPlruQDsud/A
W7VBxnOhf+ED5c98uVFRkK0+kCkItdkeybyaY9DFkev1fYMTvh6mcwbDygixneL0
zT2wcdK/7dLWjAJupxBksqOeLvSCubo1w8ceI4Y311m0DcYZwOnZqa6npRYAyc19
jNV4zBTL9euB1jk3uNeCPOBVeV1xm0qjYc7OV0NfDqBIIQtnGegATyujGmibDHUn
scjaG/htRDTL9t5uEZAVzScEb2FxLAZs01HEOfZEbcAXJUgMTmD+7QLeVFmhsnWw
3Js+kseYp96dFvNQ/8DJclu66CtdGHCuL5vM/Ibkupk3vydLjVANrDs7u61itY1P
s2OE8KzDdJg3X/f0NK+vOyUn4jP4kxX1WFEuL/GnhzopfjRdAV/fjWxMQ2hkosLg
KgIS7cmelWp0or/fw4/OAY1LBDdFvifK5PPfU5tHgOoVWvQOE4eHa2NQ8ftVNxB2
uTQ1kIHxKJXNjNtO7hu3TeAhSTw/uqp3b7i3sZLE22YmzZNfzLmKQRskv7M9AaQs
drPL+prNkIak5CSvUCe66fbd5wvFQKmX2wbxmZuEnaJdh6gEg3wLdlpKFtWmAR0W
AVKJjWGLCNOV9FVkNHCRagMQFFAbDiZ/WWEFWfimwHfnnOJiNEJor5EhDfE5Afia
klvLoriEN7Qddy2TzsZpN7/pCv39kwcTFZA0kXwX5bvSRjkUHxeOaKTrenExAXtm
SuY3W9kGkgyyftIl6y1UOZbD442TVpR6wyRlB7GwEQ0ym74a3y8n6aZ61BvCS5V1
X9LV8Jlc/i/WBMTyoBszrvyTwGON6SwcpUsQ03fmmIgBe7rmKMXILxf36hqBRt/g
mHxrsYO4pFjuR/JuWPz+8PnJ6Put06Laj5q4jpHVhuv/JYegZc+0DCLx7EtrQED8
KDqGoB0l391YKbGEDiT4xdlfTjZTL8KIiCCylO7XHFmTc5iLzZlWywsafpFj1bj9
WkWrultduMCJoYJu+aXwneax8q6lCYrFgPg1KoPt4PVgaerbCrmid9mDp7Gs9ODL
j9gO/67FOKfavdYrX3gMh4rOJqWXIcTp6meR0tr5k43cjT9gCbaka4NS3LcizWX6
m9l3LTxHZE2FmyBWDw8IRsl0gtOjNHV/x+PMLpLSZAKpRTN3hznjz8Ie5FPe8ukq
uuEdDTGJZeEmm11aIsznoIbpxVUA1FhZUz1wis7G9v0wNbhvcGL64IK/rQHhLjcA
9waCI31lkxELdXWm19FOrhXuf65/ZyaIj+empw7BgZhgqGol4xHvveMC/WGzIQVr
0daQLB87QpdVzOIZUvmsu8OmzV2CmfOgM/rfzt7hOFd8YPC9PZSqtZhLv0oBKSr6
Q4TsmaV0nXfE0o48VxDfMJFR2IZGONv8xyn/JeLVgmgJeD2zn1FDqTvdJUoyDd6b
ezGYOstnqOuf/63lIhw+G2Nou8xLrblZ7TcHGGU/boQVXmXiprZkHsMZNDiSt0P2
sp68kfbA2ZkaQg6I+R3wl5MinMgOqat8/CS3B4xuE4opZoMxiFpAg6iCipjDA1ji
I3HaA02a7z8YSYRLCxLZVYGOqbiHs8iHk9Rc4PQHniFnQsnc9B24Hp1+mWsPtzmk
sOjFrWvnHLARy5y/ucxYd2XW3KMwzGx0uJKOZ2NfOx/wyg64aNNuPdkiceod9yqG
g3dP2uzFkYYm1khNj3iWLh4jV0RWeHsc1ffCAiy9l6wJqOnrFnXCPBCvIqX9wjhn
lx78s37cq9GQKMIkVEbaJyiNryDt2VjDLw6WW4GH9Eaa91vNaC09KjOcAOacxZwP
hBZvSdj5QBITiS4YdmnV/UAp9ScaMKVl3CbFWsG3hSBrQw8h2Rooo35mQd7NWqAy
x76xMFnhytpymR6p24PcZwWeeM9EKd6kvZ5+MJBISl3hQTZWjaFqBXl5S7AI+6Lo
Rgw9NTuRbDXJkCJKgf0rkIYzkAPZ5MIB8gs9s850Pz3m4X9qDrv8MDMOQ7hFroSr
gLqE5ayDTSsVWDwMZCr9DkMqSFLU7xlU2bcPi31rwvPdk9ZEd53ekR8CqF5dj4z7
N5UK7Hg8WyzMU7cdYwHZqo3vrnFveG1NBwNpjvS+B4JisgiPZhSrrjk/9LcGR3HT
Udka5fPZuLvd9Nk8aOdMVRuwbiArFWQCsMJUY/7Ak0hHim0NViJgugkaV2GJ4WWu
nkC5boNUXGs4fRjagGYiEzpzKnMEXp9lX2oru+o2vDDmuqxJvhV/ZLy6U7G4SMoB
JYx3ECwxrRr/nUpeZVn0YPwxkfNCRfvKQPA8Pm01uG3nZ1BZajxWpX/30BpjKvR2
lmWkPkcl91lbT7YEKRqwxabWAeR2hHndhE8DIeDETFZ6Fzhf3F9GXJGQCRfNwVBW
Eg4nAeHpGdloYOmqpS0Gyw/R5RTCGVvuW3wmvLIZSROyBmegsZDPG9A8iKEc/6kj
Sg7epRYEin3NW4N4r0JF8RBzxhMWNRqU17RqUwqjJWw3Avg4EPNObI55RA2PTcyE
HypQNvfbhCkDQQFAfwhU251ZYdZldjgB0q4IBwxa7BZANTB7Bh/8XaCKcGShyJqW
bkwvqlMnj19n7/yyGQOmsTGP6SuLQLsCEkXlxZ6+FpBo66brLOf6z57EvKi97ptT
qAPIzRmVEQzyOxgkP/w2YPSFsHj6ZGSL+wj+SzPPB8gvcowpsSpRJqJ2coLKAk1m
KNa5MYx/gH5ZGbtq4OWqzEeHot555DT7zHmNS9XPjD2R3LsJR/J4zDd+ko6eCvVY
jdgYI5kzGTT+0z59Ec1lBdwwixHIpmXki0Jxi4CVx+cmqFT765/faETcEVa1YCX4
vZeE9DSubnenWNnaizXuj6poJLv8vgRZ2Hb0R4srnqUfVWKnEsqAJFcElKvAUaQZ
Is4/XfZ9dx0e3GmAulyrV0Ge6tgCUczcG/xiRwKwkl7APSUKpB/Hbpk34NNhBUOA
1ykmsENbEjv7kYHp2neWt8GtmJgPSLtTrAYEwk1ewA5b9x7sZC7LqQZKvzkcVkJt
5gM7mbK9GW2xk7Rp1kGUxr2A9k4Oau2VUzThUE4K6OtYBk8Tkp0Q4vfBT7hiKA8r
/Kak5PPNFeelmNcoG116g+Fyh+qWW7WBk/kKPvCYKNHGQUda2e2P2/gwueBuh08a
4awu+JVAX/SLzlgNXyQc0zoN3YADEinEjhEzZaUCKX6AtObAf0x2vHMu32n75CMy
Pk7XnWzHzPnA5UwGsJLm+OB2todX5PlAR/LnkQKFgPLMgvnJ/tJhiJtKmD+0W7az
RUECMC79quz6keHIaqj/cuK0NndFqvoVG3r+LsaiuqvnZ1z/3Hu/L/LGhaxLMuWx
AvdXXt+VgHfYb+LMZEmWkj81mZYOxuE9smn/M07iBJ5WT5L/Lqb/il7wW7//7yxD
fVvy7FKT/7AInaajNe6I6YI+AU2zg5NtwN+UIRWgWD6ab0ZIGTeAima8c2CisgUK
Yr0ROSpp/NHCymuKWv2KwM8YQNYN87KHtYT1K0lMENp9Xi7gvZqJYRKFObAa+Rbs
HhkzWzVWhFWI6//ryrteScRPSqKhve+h5xKT030Dmgr8Y1aDCEfXp7ovcjKg8vpL
Qz3EiZSUa7yZJs3J8sSp2EbVg2J3fRC84oYQhCSfbE49OMuQcv8pcCQTaQjo9ko9
0gBJlLik/AetmC0/oYFyVasDv1L9W/cbhxpDYDoqShU4dWiZghoAPWE1YL4L/yJ/
qKi5eljcfyQLyDKImlrEvz73EBIMMG5M8mDNRkxMCg/UEGK/4LOUqoMTBWRg5yby
raHixB1o/MJ33wI9u4QaSsWaXBbezKxLJKw3eqz4AjQ5osOppIl+UNSa7O+POtI/
7fuTjOlpMxx9kolT2BVAy2pcSfAthXJZyvRAMIJTw5X0FvPA2r6zHjP8WnMprpF3
GtUnB6ipb3REUKdotYD94DPkn7TFkaD0xhpOZcgONGmP4031apkcIZRbyzEVCtpK
0mwTuu1+b9WNIebTEukuXvgThyWZazpCXs/ySPfm3ViLwf6+BT0h+FD1Xr9PvcoL
2DZ35FZjR/ltdc5LI7GmhIk8oVF/G6CM3sZTo2OVflvR6P3qMtJdNMEnST9O2Q1Q
Oai0MZCg3CThk0aVXCErfWuewxCdDsPH+ivMJHujEwGU9Z4anaxI9thCGjJ35gir
qZBhzKwml7CEd37yYZNYOwO8eMb6DLa6HcCMtKxuB50zPoW1LSSVZUpLx2MZzvRJ
vRKO5gpT50xUwEKlpeaMPETDBeN9b97rIPsiHqxYLJ25r4w1M3wiYtfKkCmVfm3u
ryPGyt6gp7UDQAdN5BEkzlU/tDoeCxAJUSTFOf8y6gxn7rZZoBibbMZ7FHSru956
71tIRJBLI52VJ+LseO+rO3BXFvmkf4ZvGvPrHDp5uEBogWsLc9gS/QPZXYAb6AS0
XaHgOKRNgNS0WGMuctkszbaV3TcpoIK07PIH+JgExXxo+83th1gL/4D8uu5TdUn6
OkWR5G6NCOvL6QOzEdHTCtEbLwt9WwRMShXjiHS+UZ9O5ZTsFVm4jbhTwYntqmGN
hWJcun7F0UbEMLWgLiwd/yuX/Ex9o5mB2oni5Przy5bnPttR5qQCbEqypAuos/UD
7+9Xgzr/M0TrBmckCDyEw5TZjb7/8DnQCXeRngd7ZAFX0HDtri/A/Yq+PWI2qPRr
sTtON2NXLJinYzVKln/ygd9iwhmjXNcFYAup/M2MOKLRXjo5Hqg2+LxSfcRcyigv
EBac1QkcqODQQUqsmnAMmyOn4giCvNPFtgwHur3VuHyA9qByKnrU8Sy+EdSEMhLl
YFQMm9h0U8HrpwgDqhGfILekjXrfg8zZSmbaZG1dVm0KzdrNx2DjYjGAi/eotJBJ
8HletSpbph16J7r6DOzPWyYVKyvfytCkvngW7KgkOHORERNd/CTZY3T6KjVX1K9Z
ZxlEIdkSk4ymiu1bjQD4tdHuZzmo7Js9NIzR/uubAwn792XGs3bc3Re27RrTbxv7
UT3V46Sb54XC069K1LKbf2ibfYVvC3tVaEkMDP3AGBpDEcPwaG0ujm0cNWREN5yA
ef7ZGieKvtRiFL6Ag1/ExIrIJP9zs6E4JLX3RmNpZXo60qB9FSubEJbad8J3veU/
Na5Il+s6b5Ihkjei2VLg7uOo+4thvGMEACSiNk2IrNX8z3K5rD5WpT94zUjN2TlH
mk1Mhk8EY9LErjq7IXYE7M+JegX9sHc5nE1w3uBMyJjKTuA47/UoaFK23/yy/Sxv
UMqxpCEBUvgrg/9uVDYANwp5xoMynIcANlW+0JLeRuO6VfKEaATBxMz6G02gBzhk
O1CjnJAUOT9isc9RMdJDzeumjfe22KbllfBwxpBBCdoFfTQnRGRPrR3n99Js+dXX
PpmcMVVebDwXaIeq+ziDxZYbmVcb3dRJrmQJFvRjG4cmmQeq7gtbO6jXc8Eyx7sa
fKI7BrEEM/ilVB373dwRqSiryIQHK10le22otxj2/LzVhUqGCS66X8Qy1fZiV4uN
n4apjlJ7FQqYAvA0ClaT4VAXpSggXTMvNjZuBS/+r9oBBYMJswFT16tFY2d59nwW
0BIZEsNCv4mD08lND12UjXawlb1aEeW9rsPbvHBUNjt3eBNdWR5AYPRqiXL4C2+K
bQHrLI+FPtow93jbYGrlAx6YFrzRZDDTWB06HB/eovBDQdfA46fR9aTzjB3cM/de
jkGB1NeV3CsSoOSJeEfJDw5onpRjFmxIQtRk0dm2ganVLqjAojKmhjrEa8W4poOv
t2/D807XnQCPbMdugtcQUTaZKiMQErVxIkdIZQKL+fk96vR8Dz3utPXWOBoSDmDI
Ot5kl0x8mdC1JzIIFJWTl5fYN6QqTNo8e7+RRZjj7n5vYviYjeqg7RF1nBtH8xE2
rmHgruPdCAIH4vUY7mznX8FUsc00oIZLQU569e2lpHS023zVh9qFIErCserIlPGI
ReGJQ2QGKbnZXFxwCXkdh6OYP94lKAV1LaS3njhnjTxqXmN/J13WFsiV77XrUTM7
SRQ9vpcDSNdMoNV7b1fQuHFriKHoMnOJ2Qm/sSAdB2ZDkN0mjVC9FxdNH/H+pVek
dcUTlZyjiM5oT5eC1L+TrqwwmQJyNm/LIKkdKw9dFUXIf6pfaAasJypbA/d/bzDF
/EUdBheL3+EYs+FuY5vTN76tkl8eyLeqgZG+9t7Rf54Q4r0UYa9UOMmnOiYDWFK4
EhIibSeRwUTWzxu8h6bgzYXiA4k3U0pzjIDE0PoePZ/vMt8PP59w9cI24oWO9Ah8
IsghCBCQIu0E+fCearvEJY1qft6W3iUw5IyWicd9JccAkRHEfHUqcaVJQ6esWQax
TBKbiYk8fhOjxv4IFmsuPwBEvoXUAROGUWR5AvZ1acZkVbZT+Tfny2a/OREhqlDN
DPR1bV4pemB9ebSVP2XCn5wHr2b9fmr7aDNU2p584UuodtuI9TTJdwa/HLSZeqjJ
A4R8gNaq2sreR2wFTVZXupzVdCp+jzHMoaSUcKHCQI990FEYy7hd8jQU3jCkRkv+
EKDgvmrUuXnHSbLXzkM6w1GvCjMftIk0us9N0nyTwef5k5CbUjsc8h4SLOqTIz1U
ZYwunlZDTpGN3urNIgpTrQuaZ5iR6hWFgRiwaHnpo5stFpVdquacZAeq9+NXl2xQ
fwR+rBNolG4wkTSxgt4aXJaXCkknfK03SBFPt8aRbmVE1XS9cGN52+w+MLvtABfI
xk381m76yEnltFSDYrAXzJD2SZpX3zQdnemoVNutUZo+B3swGma0c9WfoQkg5sLq
06ohAwknEozbXM4S6a/fbiS010LWsL+KWz3heH08XAMyLf97Bv8DXw7AgUcaV1RQ
drDyGUs2E8dT5ru3IMC8GPkesLY6NOWPNlHHUkYaZDTHxMCKMpEIQEU0+XS8THCg
7an930U8mQjWKIxYbIQLhUc7Wg963bv0ZOJCp8m0CpOTS4P7gQX7CownCHzMlqit
m6SQUULdrsYNWi7XKH9Pv+foVGX4WovEx1rdsQIozIJnGLcTpZ9kAexIMMGV4J3b
Hec+6tm0XPBVHBlCsqync54BxNBFhd+3SiiPhsF+0T5C9gkoC8t9PBkqJHlSkPur
wmHIVzIioXskBOgjvou0/lF9Dkgj8lyZJ1jHOr0Jdnk6RqhziMkxeqn4AUYMv6jU
ka+is0qmXqGV6C/ZvVAZInVRHoWbtAix95LjCD3euvzyTQu1u2984KvwnyOKcdG+
vBFlCfMZfQPOhpYt/0z3EQxGcKCXWPpQ0CLZNuta9k+zwoSgKwe3ZipYNyItFCa5
5r/z1tjCFPm5ijYY36Z2aBqfpB0JKM+1jMBv5C2YHW5JD2AV27BaI6/wtrsLHWWt
5xTSpUQT8wOouWWJT6X8O+PFva6LtBH8NYflHA+jdz3fzPEqTQKKuN0QRB6N62/5
g2kNYRwh+vvEaEAraQoqPK7+jpIocPcS54cYScFNzDpq4vK2jL1wPNRELI8VRxz1
4ead08yfRaAX0Nh+wL+81Ev8r0RjsLeH02qGwUGKdydifTYXekrGIWgjNtouvQFH
45y83k8Lly5Hek+hIllwGJ2bUuUoDr0Il6Mq7+6ZIyiJp7dswx442Rn2NRcpY3AI
PLKl+uL5V/fi1e/+0y5UT3U0NFz22cr1AI+ZxsE9TzAmOHsNMjVT0Xqpv24Coy8O
NnEFR6rmCKGNdnUHScB47JydOYohofaUE8O3F3s/LIHCX3H4QQB0JfDJevD52u7Q
YXUMfJ9XDk7xarRhHM27dNbN439Tvvf2gQhfS8vJYVxS+366b2WtbHwWng4If7Ep
xXPS8V4g0+H+L3eb0tWH3EdBBZZCohNSEorFPnuYtJNw3nNFM6/TsDf9mdHCpw0z
/CFA6m4To/uRrUEcz6paWgZ/VAt2wzJ3ZLRYbptO3Ufc16tcQoBb4P5ZqEU5dts4
By5Y5vc/hohyY2wcjTdpk1LY70E70bycIUuafIPplT0WrnzMc8jlyCrBGLegHhCu
XGZaMhqF1dXm5iMGdoNOuQNF78ge2+DIRPDPTO5C6HOhJZZmhCnxNEkql3yhaP30
L3kzpi+gEixsy0TnU6hhiVFjaWqWbDBjaDUPl9lbPbMfNWuRDEvwOvsEK272r+RN
4GxDYkMvjl/hBDffE+0P5dSJ1Dca7stLisyKhP9FJEU3iWC7HCjjXqh+RSQGrh8v
uvOozP+BF3bD+PTPpsNmVHVJ62ea/5/5X0hRCUFAgGMPjZtoebzlRB5qyyQk9mYX
A3tjHFsdxZdxraoIJ2GnfR3YPQZuj4AqhjBBx/ahIxzYij3xeP2hXWorjNFn/PEM
Go7KXkKYP+Lkq19oYL8sRUCrUItiVlHndjbOMMcwkP0/rX8wpwwakv59G5LKgxMS
U5mZ4Qs0GnvWk1ZIEs9wcBTs5p7QA/aCYnTnE+bCqoPr2cJclapgcsSMjx5NI2sL
F0rxaUgoQjIv34MYMGiS8QR4cvzHQZnucTC7C6DMeajV15taDk+SLtC33vd0rYVV
qOHJgVxyYstBUuq1bO+25XknShUj4diMYn3A4AC4Di0EkZga0bAi3kF39TtkkatN
lXCbyT2E/QmvtX6X+6cZtgVoRHcpcFxwwQO7tzkAKakAyeTzNv1XMeq67MPQRlTL
hRWEGqwI4T7wmu9LIASKFnt0g1egyCkD9M7fEFuN+hW2ZZAUpU+IeGl3ELKCmVDl
DZN5ukEmQe2JPP1izY5MUvREE6xT0DZQCsqz7ZflBZQBTKciSAyLMcmeGbuOXW/w
+BslisQMyf3PtqpQvovex99s56QAZ8lGtWv1hQFXd9vLwXrKRM4WqCmdVNr/wvcf
2DuQtrakWFyTwDtZcfqLExANQvzNp8R4IuHVC0r2AMgTlMX+U25pckFyvW/PFAIn
9xhnoLF8OJUkC5C85E0kgYFZgeL+Gnv3HWGtxI8JkoTSG8QtOikepftBaa3PSt6X
1ddXwG3fmI+bjspChoWg/9tEwwfqdlrruzzZxo4g1d1v9Zn/NEJOkxLpEub81Ysz
2YJJhs3jQx9qFjMeJ/Txd0YIZrVveRU41uNlbVrZcDZtYkSXoU16YaejyNeU1fIw
QYjUBYV+c34YjtrHk2+tYyTv8WLqySRbYlm6EMkdPIW1FVbkRsNSmD0zE6zdeNu8
8KYdr8cSRnKrf33kU8NtEsKuOPpLqZgOY2D/1sZm9LycCuGRrMEL583kqGWMzWRG
nMhhq+AkTXoOZHSIEz0V2gbr32bPLRa+6LmOanfl6igcn9P5njD5eIAR5YMDYTwP
3ECRDwE2uj3XiOK7lnSdyOW5vbSMXtGh+0ri4rnT3nfQfW0+ibyIYpuMgiXgAGQN
9oYEn63pwHLGW10V0WPItHqVNcamPsm00AxaXlLOSdd9FCIgPTpLX7XsdiUifkD/
iLAY9amrQatSznHRgok/ViqTGT6ySrNidS86dmdVbMg7vOrjvynqSQDLda+JaWS8
pdFrVxvk8TYEgmNuF3aK+zPwq8bQjf6ZALN/zEhUdMXVsU3mG87+8/kf4MHtEcrr
Vyco7y2EWbDigRMTD38vvN6sDjCiSuXZlfUHNvjHUp3vbRbAlNrp/Qf4XDcUOwLZ
U2rVDihHV6b88GeRkesMNl75a1LJbFug5btXPFuRaiSQGRl0HuuSxYFJLSXvyXmF
dZcdHsFlQ7fZggjMwC2Zk5ByBmX6PVlT9O/JNSk2mzvYXEYB7Zc06K7fJrD9MOhu
22kFddKaaVN1cO9CmE8IDW2oq933FzJeZIKTgcVKAbuwgEU64ewRujUGcOZmwoWc
kqxhYhASEzxxhUTFR5fdwsAJtotrssXtCDV5LodtmFcR2e+zaSeu3/OH88e8hCXC
rLb/vj4Cts0zlXycVrqhE9SFMiz3K7eucTzs3fk0xK11gs/FNVmhDAs7rzLZiFJt
w+oLTFp3c5MYGjKqSAPvJjkgu4BFXyNZ2v/B2I5IJtH9G9M5duY+GrhzZVOvG6iy
hIbXe+0LoVDPhXIjdqYduIy1L6DOLizzyon6D7+1gBC9zzyfpHkxa62WqKlzpbt6
4Xzexzag2Tm5KQyGBTsSOgf12m7YHpp0UNmJ2ENpM/gUjPfk2fgOkVUzGFfiIiiU
4/l8kl0O0GBzhjA8JUaY2GNKOSwDusW0KB89+xPfokQCsMe6xiu+EiMTK4yDYdt4
xxRDYmq8SJ7Om6bj6ZqRLlJ+2NQkI9B0DCbU5lZwCYlB8HDKdMDd2vop6Nb/hoaC
pwdsYwif0xLl/c0107qI/KfKCEn7lM1I9LHh7V8OjY9wM2n6561k+g1UMxkvdLcA
B2aX0iiPhIq5Dd+ZDZe3wDAk/G+I5aQ/fQlDn/KQuuUYxkvwhfHkfvlTJFuglAc0
5ONEXO3Bh2mUQlifaBdsCSa1C+XpU7qk9NLq+QM/nT5BJgxztMGrSONmgukzvYDV
891gPgMVROdtpoPMhw7JPwnzkdrjmkydaISXPdqcYOMSwVUYA0jS9xgWqp6zmcJd
sub2shNdB+wq5MT8wECW6S65Zllr3iiVnUdyURxSVOptrO67zxmyl5Kma1rfFCcL
423duSwD5zx7jGvcY2uRAGEhG4UdO1Hk8TKAEFkJhOXzj5g2kVI/K1/kjW1ZWSDb
JaDtHJgNrS42aBon9hFJSSwfizRRgpr2rNuOGlSMGiGtt1fHPGa0jFsGSSt0L3Ez
jN8sKAHtjNGv+1whz5XOaTH3j9/xjlsyibvupiF5FtrTocVCZzoIWTLHsjTk2/gi
kHbG+G+TXYpPLPw5OFlxYKBWjsTVev5pH3Gu+J4uXX6kjCz8YQzxm2Busa9l88C4
mln/hB/kEPn88nLy++oW+G2etCDJ93bCFYnSpgRVznFQ0NJcq0/ruxKX7MzcF3d3
aEA0NvNaQIT9edVxNAQxmc1HoLGUWzRyxxLfvk3iePu9Pd/KuYDgZk8HlLum1uue
djkKsTluX/p8esEzdkjqpAaHXPHfCWL1GjIbNGi2dxtXuXfK0oDEjjCCUB5CUPKR
BnR1OOyvqsLjlWti2U8OFCpdgUcQhyApIomR1u0Tf6Ij+LKMS9l8fz1vg5kJjII1
oa1xxHqRXFxyMb/zZFTeRv93K0bCfzuD4jHO8W51u3VEgE2OkJcY1kOs2xB6664n
ABk/XChKkjNwJqcr0hZWAUYmfOneJwv6k5z1jF7UjDY268OB6uKE5ZaktRu17Ej5
hbe/UHOzfjo/eDH8Beu5llMUs8B5DLAWNQkvvoUl4O03n0PhPqdJNWn30fQgCfe6
fcPxZ82JGEO7lC09/vgZ2VEgatiw7XM7K9v3b/mD7ZDjreNMFDcu5SC6vBMPTJLu
sx8KkgumHnVlZkVR3e9TkGop9nBHd2mmjr9faRUsJjpahRUeTt+6R5i1+f2rpwTQ
jCnbJD9tSi1OE66N/AyFsSUo+EVHXm2DGWVrOSJef82T0Lhj9dDx0mSSpz5WYeFh
m0dHKkP/diLASoX1sbN+UZWyeWFGHKtHMxy4u+UuLTW8z0EW0tYb8UQ5N4490zYs
/4MIR5K9fpHsiJ7UOQpfbyNyFeZflhbiNslJ7zsahYNuvgfv8MUXXux8OFUkZEmo
O2YtG77vas2C+U548kRMgR0GNfjQ6elAE8ChobqnjRAPYJiS7tEdQdZUhBSkpa3R
rqEeyzWIca5s0NKdbae+aCMC4N3GoRTveoCKWz3iw7mlOyhKu9pPAhqx3TbVS/Ab
ZsfazYW05VuKwnBvtmNJFML+AgCwglaP4+xyAwIhokr0mEf0DKI+fYcFOurLFtiZ
1xA3oF+4EeRxduBROPUeMEnSocxnLEqbXibE65MIMKcv8/TixYFhmCH6XkoV5Jon
LVZbI3tfNaN1hYeKHZIAhJS36hxQAlYQcDp+Fc5/ePnlbUm/TWRixg3ktdkopve1
958iBCIo6Mgilsq0/d5YVCgur+8+YpEXj8G6JGLF9bKRHGaouDZRJlTpPltu2r9f
/P4JVF2UtSmR3/a1JiEGzUHeNC/bwhmFmmVnfWrXhq8yEgMffXX9bPSgiJ08Pb48
yYODw9/EJCZ0Y8c7mQcw0P1sFNY0D1wb5F+zaSnB4P+VCmKD5KGj5RNbPLWFSPGh
9jX6fmscxycy02ZcXLgzihOLsMJLGn8Nk7Dx9e40vbJm49vcXkVwmj64C3Zpnxph
OP2Clq+A9z/3z+VKsYokJzyRZilOXcbFjMfrBoFL+zljpLM/TlXyQZttSGDZq7qR
/nskUN6Jk4+jKwDZUySsafg2STwzUb6w7v074O1tP0A2kmsV3UvK+7XWsu3r6LPy
tEf/Nz4vyYCoBBGEckbNCCBatekHKkpenTedLYY444LKWm8TuS3mx8ptGsNi+8rx
9g9L0Wi0/H+9Dtx4TvJmCP5JcxxzLJA03DHswETZZe7Nwe2r9H/xY67OWvGZGOzJ
oLbwc/X7SrKJQNkl+ZfpGVQo9TmPNDhyrLzApOqfp1Nc7/dvaJmBx2j6dliyKT4z
+kz6ovQJ1r0iQscwTiPaOQv0LwZ3FFwMDRA6jZwNzVD0ue2CM+crglm3SHGzEC5M
Hr98o1B9lh20J2C53qtKf4q6iikTO2xMvjSsRTXsPz9S5bMT3nvoSTeL446DNRLj
+1Z6ubDJcNLLpFjmvqmhYzVN/QIxCjEOYGgBNnHmxmnsWm00wrI586r5qijabZpc
2wcPa+gmTabQFRgS7pOEdl3NJl+/oeCYT47j3Fej2WfvP3St+yJJmnPrCVBiYf4v
EtDhLiHo3DhV39rDbony5uAUfKdIvAguRcoqX4NnIPY5eik/giAwmDPriNWJrDmo
WzFfD8dHM8uh4jtX5ilm6TViM2kb76XbsQ/uJjxVHdg=
`pragma protect end_protected
