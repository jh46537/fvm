��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbԒx�#3 �2!����=8���:��/�/B�s��ރ�'l�����C���(Mr����7�r� ��#C��dLWN�)<	bU=��*�_B����:����c��DU�$+�'uR�T!��!���c]Q��������1��B؁	��Z�6��'kǜXq)�10L���%:Ԩ����+1�D������/%�H�v>a2�u�y�;D��b7�P��u�	�Y�#U��t�4xD��*�X;��.�RN��-m(״���z�]�V�$�ߠ�d֪��g�he��ͩ�@�9�7��=6���i�Z��K��b��U�:�2I��fX1t+��:���ڹ���ȍq���f͂�o�s�%��R���kƶ���pŊN-�4p
e��V����,�� ��RJ7YS1�V�w��<d1˹0�#��O�����O�M�p>����~�B-\�׬�W�aY�o����1p��Ȕ�w���d��Bo� ��@m3}1���t��!���G���'t"-eA�Tn^�&;]�. ���S�F�Na���{�Yr��6f��n�<aKJ��\z��.�-,i�sh�2�(���04����xm�0�Y4֯���$�0ָ�����>(i�F���Z��l�j�rMCG���Y�[�ij��:p%�dx�U7�aT���R|�J���=$�1M�S5� � d�>�H0-�"֖�J<4l�R�6�,��q��32�aE|t������ۜ�C���� �t:���s�U+T\�t��j�PRR��jb��aZm�Z��!t)�2{{%���5-�>��s����5R1��΃��o��DT�Ԑ�0?=����h#b7�<��L�ʆ	/4b�h�1nd��*R+��#��
E�Q"�����!݄�ˠ��v�K����K԰[�% ��n�Y �O&�c\:�%��&L-� ����H��
-$�.��9qE��L�ǢR@fb`bɥ8S9��yA�*�z^Ž�x�^X�_#;�x�ې۰P�)[�A�/��Q ����Q�^�M���k��x����"�R�V���-P�ӕ\����4(�O�<ݧ�]��;��I�����i�P�F��:��zs�&�C���D�nx�%]D')�<�@���=�S���b+�Ihv����S���HYUY�#���+7٣�V��P�}�,8������0�(��,6Q��%*�K�#��tG�Q�.,Y(+f��R�5�|��9��0�S��/�^�8+�0�H`�z�����PkƷAn��ҡL޶�Z]��ɣb���՜�H��$}մ�]g����,�7�d4������N�8W&w��TG[D����[�Ξg��� \\�*�
��B<��KwJ�f�����{��сEE��1j�;��6��(���/L�X�C��>$_��z�KҸ�?l�j������.�~5)\��*[b0e�{��w�x}�W��pl�Rۺ�7Ќ�l�m>�M�Z���پ|��������PK����tt�Ib-���w�&�C�t1TB>3�@g�I%	YI�w2mZ>]t�e�Hq`E6�6�H�R/�4�1�|�����N7���i-������(�u��{7���x?ح����r�y66�.˽a<)�5}d;o�:�.�:��J�K��FT�7�X�[��]=PC~I�\Y���M{��C>�O�j�rl�1�7��<�/�Biơf���&�����8I~�!��O��^�V��}/F~��:/l���B���F����
��Ӝ�_���ZB~#ءc��Ѐ"˿O �E�먝�:L\@(5�����24�3��djM��!sL�}��Tt:EJ�K��p0��H���S��1�p�l*��NRNő2�#}7�ܒH�gܱ֢�!.#$sG��֬�yX�F�J�����.��y
�S��­��r�������&��o1Ô)^�����4��`��X���/�l+N���<��xU{2nZ�=����O�(��#��z��a��XAr�ޞ���d��yMFZ�/K�S7Ҝ �8x�8Ȕ��6kG�����0W�E�<���bg��Ċ���g��Q��sE�B��\���<&D�4�v�N/7Ça�\˹#��+��:n�?*�� %xe3ݟn�	��;�󽪴!�,&Y>`�m5eUS5L�(V���
4�.��Ůgq�f2��*�Ǌ%���s1��`O�L������y�rT/Cԕ���F��/:鼡4��~�����f*��'� �؀���x���{9l/�%6~�rvW�/�R����0m��6�eE"@a���l���_�n��L<�7��������i�R�k\��7�;�M,���Z�J��=�dSEn����:��.=���"���J�ax]4��H��ш�4sc��,�]�
z,���(A���)ym���P���3�º�h��5�|��PH+nAq�Vw�#�o$�?;)H����ej)���䩌 ���'����i�s�U?,E?ay��#� �3�� I&~��᠕�x�ޱ|�$>͵�@g"�8���Wo:�#���{����	qB�5}u(��gI��� �ж� ����W�T���U��-:1�lD(��N!{94Y�SĘ>�dE���/��!ߟ=��#��D��fld�%�DPE�X���A}1E〱ӌ�k�mGk�`m�}���mrY
���{�O#��8�?w�R÷>���:��	�t		��G"a�>�:�Bܒ�Vd�����g �b�-#�ID썪�I�o�)�����]m��^�[�y=�g�;Y5'[Agf@��U�a��t7�,{1�%ֆ�����b�2(�m�U���j���ӹ>����:-�z�-���=K��g����
 ���&�Z�~�d�	j�]Ħ�T:Euk��T�s��+Eǘ��]~T�J�ױAQ�\QQ����g�g���X�u�,��&s�j�lA���^f��k�ްt�\� �)n�y�}�H�.��
R{��me/��*p�M�g�^�AD>R�x��zZ��ا�x#-c��HPͶ��;W:��゘�J�I��Rt\g�߱`�RO�1�+�6}&��)��*>��|}���8�i�_�I+x(�j�[S��'�+��G3S7�m���� ���q,��.;b�T�ۮa�n��'�Wo��D���^��)�b���	�������I1��ďsi��iP-n9���W����)Ʉh
��Є߿�H[5ҠJ�Cqi:�@��DJ~Ѫl�<MpG�&�6=��Co���q�f��ޑ�)qц \H����/9ԭ<Y�4S��0a+ᓒc�@ވ�i�%`�ڧ���rQ~B�i
2�M��ƈ���aT�]���}4|�%�-d�]��j��|�2��G۲�uڈɁ&���q���Ē�ٔ
$uS��p��+:8���4B��/kp}3ȩ��CKIM��fE�M$���L�}C�f��8��e�F���5�R������9$.'Mgc�{��fpN�gI��D]/{���%��,���Z�U�PF4܈��"~ȧ��C�e����ﭢ8�٭8�/ya��E:rqJ=5p�͵w���{6�?<�?�G� I���QM��aIX O���;̌w��,��mټ��R�]�u�,�{���7X���ngi�$憍���+tÔ�(�wq�� ��������
�ǴҼ�T�)��7<W�	�V`����%<n�K�K�� ����uE���\z���"U����i4D��H��,����ԩe�z���|�n%��z�>����:� s���
�!����e�b8E7�c������+��R�Z^/,�6�Q��B���ժ؎-~��[�+���dE�ߕ$�g�(�`���J��J�`c���܎d ��E�3�U�Q)>P����k��f5����X�k|'�INs���_�~(�I�l�vE��,��d����ڔwf�؍��\6�
������ڙ�Q��-�I2��4Y���;ƅ��I���ל�9�}%QtjTz�*o�F�t6�{���%K���%�g��u��Ew]e��IEa����$Йmh#wX����z:�_�t^�Z���i��h�Z'P5Ð� ӥ�&���ܘ��xC��d-0E��>&�B�������Bd�n��b�v�K4b�����k�ȉ?�ThVem��,&��M�b���AY�#I����
d1 �y TcЉ�i�i���⊫����1��ѯ��ֻw|��5�c�x��ʎ"�S
G� F�܂��7���Q���N����8Zpn��r���&��qFv�LM�OQ����|g��=����d�+���ϯ�����>��a4�_���e�	�/O(R��E'�!�:��X�wL�i�\~��5�3�Ç���if��@ԣ���K@4�>&&v{�ј��ʕ{�>PT�FaBq�H*T�j�j6ҙ�H�7N
��T�pAh$,9�H=$�c&��(�lM? �C���H�:19�O:�������bU��٦��׉�d˞p�-ܩx���p�*��g�JԀ贬6�;�&>���8E1�m�3l3����l<��pG�z��m�n��Aڻ]�@�f`V���o�"�A����Ժ��/s�<׵S'�������o�	���I��HjGd\,�*��uX��j� ����z��[�����O��d?bz&K�F.�]�T�s��t�yd�؎o76�Dަ��(�hU�r�ӊ�8���T6_�.ሩ���}�.�CJϓL�S����	�o�ߒ∔���^w>����(|kk�+p�2U/��ez�Ƶ�k�8�� m+��.�ɹ��n���Ղ�X��`����X�XFL�p������3�ٱ	g3�̺.�Yk�I#�ؚ�ϱ�j�kb��k_M��s �Ε��krq҃��2��\B�3;�F�Ǒ��d�la�.���$fo0*�Y�ܽ��p�.�3�/I1��4_�E���7�|�S.��S���h�đ*H@��%o�N�=�J������a�a��Yw �n]�w�b�t�G� yc���n�{b�$�#�����^��~��>��d�<i.)���z��[��R��k�d j�'d#ʁ�����ߙ�	���H�B��}������/��凯 ��#�R�����M��V�0L��ziV�@J?:�sSB�ƈPȼi^"������ψ}��A"�q�{��ɦB:#<��A���2���qg��}�N�ѫ�x*b�A��W�~�ծ�Q�Ґ6^�sN�c�*@�"����T��YU�^�w
_6�(�ܵ+��N���e�� ��U�I~۴��n,�ꪦ+�W�F�|������!�O)8�2�4</L����֔�<�F<��u>�a���k Uჶ&u�K��21js�+�b; GH~�&cxI5�
��de~`���)~�t,�e^���	�'��T��,W�W����twxg��~"'=�<f|�ñ~�9�ݺ �i^�t�)����a���H��<�<WN��A@2��cY�3� �"MN���ް�Ht�Xm�l�d�@���
��?��o:˸8,�?]s��F]��-w�!z8�ZQ%~���W��^�?�Ͱ1,�97td��tM*,,|lwK���a�E"ƅNo�@�,�J/R�'��%�y^w��~Z3z�a�<bV�	�᝻�Ġ�w[��W�
7_>��K=&�c�n(�w�ٰ�Wp�-��?�B��L7Iq.���?�|�0�W�1���6��)����U֣t쪯��r���-52� ³E.�	�~p ��8���"�q�̓k��Jpě�5��$�V�ѐ��/�����ma>�|����̋Ր���3��e�L������B?S�s��%�7��Y�{��2���K��C�˭�5�b���lw�A�9ʹ< "��C7s��c������d�?�)�V������C�i�`���vƀL�#h��<��"��2*g�!E?Hx�m&���i��.�Q��~]��)v[	O���*�3��~4ߨݢ�fPLh���ֱ���5N�tK��S���(>&�?�� �\�`�X���穙����NL$ h�K��u<��[�Dwlf�!Q,�$ck �VT=�M� cHG�	SI�E��X���k#��E{2�y�`i���դ����4���&�;���P�mM;2�����\F�F����3�"�16���S��!2���ڶ>�89�I�B/5��<3?"�de��Q�ƣd�M$�ͳ{�?ځ���Å��J�&��A��>h��%Ki(�kQ�Rm6��h�bXĩC�.��Ya�:82��ܬ|��z�Q�ʍt��o|͜��.��k�t�X�P
�@��O��ܲ��Wާ-R䵾�7HoK�l�E���N��ɜ�Pb?
�0j�i�qAR�6�^�+g7	��-��U�N;ȫ_zOq�NP��W��Z�r�44��-� �+oR��N�BЃa�Ȉ�;��Z��s�������Y5�_FO�b=��M�~��]�����ɧ �cXG��[�6y<�tW��{�A�!I �EE���"��>�=�^���yn�KJ�ɱf��'$�OHS�;l����Q��9?�'ڹ�+9]�wV�3��L+��kˊt�Jy��4��w���Z�/U�aH��U���l�M���m�b;�?D	}q�7���#����35�s΅S�������x%�G���c��-��NC@��TS������VB�>ɚk�9����+���Н�a�'���~�¾�rn	!��OISK���⡡N�::�zCEW7B�t�R�j�Qt�R��l�롓w��\��ҹ���K���΢M��8����3�0��wfL�:����i��d~�@h2qz���؊m���WW�5:��ˡ�ѻ �]f;2Ūx��^�A����o�N8�2BP�;�)cțg֫�#�_ȗ�E�.�@#�����Fd	��	l�v��sR�s�Axx,��|h�O��FmX�C�7�$����[ao�tpY�P��Vy�晲����=�"]B��D�[V�_8����xB,���x��T޺e���r�fKH���W7dLd��#q�N�2@6P�U.
�:�hL��kE�%�Ǧ1Qlw�	�̃=ށ��3�u��=x�;|�s��`���j�?���l�TT�Kљq=ϴ|��7b�!�p�d���/�LE �!A9�n!�E�3
�,l("����>���s0x�E���w�j~�L*���\/(��<�K����26ϮFA��ŭN��TmQ?)f�o2��f`���~Ϯzz�z��Z�i����������5�"�&��0�E��q_�
����4�zn�}ě�;��-v��e������т���!�M?��(��̼��"�]�H���nةwG5U�h �;/^C��.�I������	�w�m}�U�煍{u��<�������|۹�������]9���A?g_i�X���;{�n3m��0�G�S��'�w��Vj�l��!�T8���e��V�ކ)��I�Rw�%���e�R�-��Anܣ�t�`��/>���8A�ʂ@1g�cq�8I �F`jC�Iᗍ�����sZ�Pt����~ \=œ���n���1K����b�iI�5d.��ϋd��3�ϴ6O �iΙo}��z>Y�@UF�x�W=�Ç ;�*Mg��]����J���W˱���[C�@��o�F��Wd�1��!��BQ����;u71yt� ���R~ko\�0��j�4��������FlL���4Zk�B?E��yX��SU��<�+U����j^P$�:\6�C�$�Ȣ'��?c��j�"0s��	4��x6k��|8��a�	��дD�/~�-¨��	�J��P�Bp��k�)�ώ�w?�G1i ��00G?�����m�>��	�/z��RoN��ٖf�t��L��>vx�E2Ah,D\�ð�o=ʂ�"�H�E����l������K���t�� �W�Ue���g� t��Y�4��ɝ���_��=�K�<����6�0���R*6��	�ˮ~���sg���߃a�~3~�jύ~���e�1�6Ӹ4n:��ɹ�v�?�~��N�y���Qo�`�<>�!@r�n��5�8��Xiv'�{���<Mw��e$`�)\T=�%�Wp�����2/i��I9?�ݏ�afu�Twf�:����	Z4
�aHaN{Y�7
��NP�}��A��N/�g�G��g�H*i�؎?JdM�h#�
�����!;Á{�Cx�����ɲp�G�p"f?�9�@������e�*�l�(��$�6��p��v�ڰ����9������Gd ��|)����twp���|�G٠ᘳA�&uj���&N_���#Y�+�����^I!��oK�K�4l ��6}�i����KL�h�	��>�Du¦��A���?���7wY#-�l�x����u�f��<4bb�Gzz�X�~ީ�l�II�7�Y�^�������pϫ@����Q3�V눅]�HlJ���d�碆���Fk��R�ٟ��5D�+οQ���j�`"�nJ���b�L��ep��ܶ6]�ގG{vÜ��5���x�Wm���4x�O̶	Bm���I����i�)MgPK`�x����Z�[�� ,x�9�],�Jُ�f��hv~�I���ϒe�3r��_�L	]��N��5��(�?���O�]q������!�'c��Q����TI���J�k�D� �rdPw�q����7Z��R�r��z��)�׵#U�k�*	�qy�R�8�U��g/����,v˽W-�L�<g��އ����b)�ϯc��X`h�w��O�EoG��J�*�����8]Kv���)ʥ,A ,������7c�s��0���Q��^v��o)�k������sG&J�8�xU�B���Hk:&[�Ť��H���F���E^���Κ_[5�$���2����8��'�Ox�%��ab)ԅ�[��x�y�}����7�6���$��sR=F��{�"�}8�i���>��+Bn>dta�����#�_�J>�O�(h1%B�rt����!���=$���q�H��XIڇ*o��R�{^�.��f����I����l�?�pWi��R>B<�֥�yV�5B�4_ϗZ-�	yEl|��rnK�Ѡ�������
a&�G;�)%Y=��A�O�!��f���?^�'�9/�)dRǵ1�u����� y��aHj��
�q@^�W\g��"��T�r�;iHb��ޒ4��1g����_�~P��+�M�Nv��90/,�}���T�(���i��"�1����C�R�k|��Ĉ�2@�`h���lj�`	��c���^��ώ~o�Z�^����8����	sm��QO�F=@�ݿ$��{���j�c^e�!]-2�aĂ�\}��[�7�/���C�ڿZ��QYaw4|�M�p�A���a"����NW:�4��=|WV�B.cIhjh"�wA��WA����N���Ӹ+#��T����k���j�4��%�6���u펦��;��A��1��y�1,��}!+z��i'^�TD���{E�Ru3�%w��v�<x����_��`=n܄MO��Q�{���[ެH;n��bs��8���pع6��_Toz�����MR�s���Η϶����w	�y����=�T�c$�K+�w���v}"�{���jQ�|v�YQ��a`/�W�	ܷ8=�c+bTt���2��Urj!(�LJG�B�&/\���ߖeK������͋�k�Z���xia%q����"��ZS���b����K�������O;��/͎�LE-�S9��k�V��)o�h��?B\��̤03�@�-��h���Xӷs���4Y�~R��.�H�E��,����3	˅���BC�|;��|ofW�� ���"��"+ZK`��G��f2e9wA�՜�U��X�d�����Oq!�O�.�7P��Q��򩑧Z���f~.�&� :>"��0���~%�^Y$��v��w����`�ƭ��;�{��W��6\Ɇ�q'�z��m(���G n�R�*�`�?�!�
�Vj�T)5S&f;�_��NR��y��y�\(�e������(�N��\Ǖ���:ϳ M�~����ͱ}���i��#�-����Q����a�0��D�/��-�*���@����&v��U7@.JYB{�r��E���s!j1oVδ���H�?${�W�hL�n��.�^�4��$�jiH��g)l�Z���\);�e�g֣@A�"����̲�Vv�2��C�l}�q�|�h��m���ZY��v�ꟷ���I�p����
��[2�q��g�|.?�%F�Z7%��+$�gkh�`��]�@� xO�&'oU�H4Orb�.mj�!Z��D	�{;$�^�dU�w0ʝ)���߾�+���Qˮ�*£�q�J��t��=(�-���W��'`p����� !��f�(`��]+�~8�O*��5���k�tw��º�8p�Mr&�D
������ΘK)�m����r8z��6�-ח����N1�9���P�0i\�``�]�2�iO��3�$%�C@�b�� >�nS������O��
�',�E�R/�4��s�]���
=�2#J{7��8�J��+l��*VAdڥA��p�V�['�����S��:��RP���'Tt}��T����ܽ����-��Q�DZ�~ �y1�Y���c���);�u`KB�|q�$�Ƨ��e�W�!��9������SL���E��7��H
��md @���`l.N�_���N�[Ͳx�k0.��^E���^��A�o�i
P�-vr��%(��=�8g�|���sڠ˝P��ߙ��4�	&fו�ĥ��A�О#�Eу\�M3�'`+m���۸�&�$�+q͌�9��U	�J�u.��w ��?�;���Ԅ<l�4ӽ��J���A�1�$�Z����c�*c��[�8q��C[9��7�C<�G=C6�s���4M��m�[�x����kF����K���s[��[��g �����D�����)�j�[XC��<$H����M���t5���T���:�h�_��e6�3��	��Iq;�8��`��'�0�*����Dc�����z� �ەlüL�Pv��qxV� �uc�Y�}�7N#|8�Rv����$F��iϒC��7�mM�z�q��H�7�UT���� m�(ww��Q���U���iy�$~��0�;��Y˟rk9.]�f!q"0(�:wܤ?Z��6
����>6�捳ϣr�nX_��@oe���X��L���Z�En3ș}m럕�Mk�F�S`�1��2���>B4C�ydm���x&s��A�|qd>؆ń>�4Q,�"R9�F��1O+?��s������8�cҵ?�� �D�R2f���V����E��2�w���Sd��*�T�,�dx���7�Z����bҀm���3y��A�ųRM	U6t!?B���v/~���6H�A�ړ�U_��� �P�����s����x��u�uW���%�~��0C�i�/��w���bW�FVD�@4x�����X�z��'|΅9���%1�j���	}3�~��d��#�[��zጳӂ���nav�hH���Z�|����YJߓȦ����Y����og (
d����$�	���Y���\�ˮ��#�Ȕ���3>=���Msw.�����J�ƅ,�b�kp�8�(}{Lb��Q�#��)�݉% 3y��<e�/8V�zcd���v�b� ���T[�  �ԇ�Ȗ�B����o�&��!�;�1�Z��#d*��P�C^���4Z��_�^�{ӼW���S j���W�cE��!s$���<l�����AE�Ѽ���rI����Q�ܔi]��I�BV�Kr����Z��*	�9v�!��#�B�`�����Pg����*y�|H��$H�fn��mŨ�^���[�6p|_#3�QB̆��!��� R�5��TrDhkP�q��O���]xdS�^G�,��VxZ����aOe���)�<�>\_�w�R�=p�e�:�W��G@���r�B�f[�����wQ�AtX� 瑵/����9�����eyL�Q=588U�֋����f������9��Ո��?��"+y�k#�O���6D��b�&�v>�֒.���d���7,��m����>2�����5��x\�&K� F�g��KU�N̆����N q��?�b�����-|� )u�Eq\Yb`&ؑt/�PD�а�y�'���ݯ#&
؍LK�B��n��F<����k�_
� ? �S���:r:bH;�����_ܕ��88~S��mŔ$MX�#^b{��πF�W\L��g�qӜ��g�K+̐��8�cOW�L��d��:k�9�E� �Q5TψpWߞ��Ac_��F�=��pM8�P�/9����7B��4���2�hW�q��E�tCY��7��۠��!ro)��"k��I%�|̳���;�=���|�)�h|�����^��v�"�v��{�e�b�!��r����@N�RcNv�,��1=�*����=)���#�9ut��rc��(,���4�p�����;%>W3ɉh_���0��u�	|����x)xRY�~������6�ÿymG$G��:ou��Ϧl�f/��e3�	���M����4�_HpXz4�"�F<�%c��=����R��rI>}'ȄA2��!GҐ��;ߛMfy�tJB��%���
�����V.�*&��jЦ?)�rX�1��� ;5�G���T�˃��_�Iý���*�(�F׀{o}�M��9��Z��:[�ށ3	8�b+��Y���#x�[�����*�Z���B���^Kb�ʍ�'L��^�S�|ڳ��.K.�<��-͋�U�|v�L&h�Z��_����Ŭj�����M� IS�X��<�j쵋�mN�O<�$��/���j�3�X�n<��T�x�v�����/��@c���~w]D5J���܀�m��z��"�l3�|`{[�!ıǑ�ۢ��s�2�Q�q�Y�#�Ռ��ZXBca{�4!g%����w��X�3��Rf��®�˞R\�T _��~&�.��������E`-������[���
�C�6���oW�L��!��H��o/ѾvP��-H�C
��9^*�4T��]$8%
���)��[�n�f�i��U*�K5����;P��y�'n�m q|2 �}^�o�4��73x�$4����m����_�ؑךu� +U���}k^-үa(Ly��wL��:Ƙ�a���`U�/9;O�ӈ�+7���(J�Z�	��xC��x���! \�6+���6�r�L<Fv���ʨY��@���:��!]�.�
h��&���M��~�NU��:)�����}3����Z�4d�#j��?|��W�����e.1M�O�b��e��c��=�
�
nO�|Ԥ�z���sYT��3*�l��̤��
 m�L�h��>6�R*.�n%(ϗ� �"��O��o�W�a�KuZ>�%;��'
����4C�ь�{�~h/�N���4�`� ���$�,���}�T��F�ǶELԴkv*�oWь��|	U"�E�(܏��漏tvu5�87��U6��~�v:��)��ߵI���B��QH Kn@�ÿW�f�T��e!��~5>J0;��3Ā�Ɖk�n6ݻ�ш�Z�Z�!���a����
�I��V]'3�u�߆��-�z�����O��.��RMd.v��� �[���d���aY4_��|&�a"�0�5�jeR���:b�Q�Q����u�Cʚ�� H���S�ק�4�%�S�[_��4�5��=.i�0��Z�e-oݙ�!�u���WvZV�
��>%�l�Wm�U������!�VN���S�)V]`��)���xze^�:ꢥG�s4\��%�΍WO'z�r'y �ǭM[�T��uZ�K�>� ���qѸ���v��	e;��d7�#-rby�W��V�G��Iz��|�~^� .�j��:��������(�剦�bN�M}����j'�@��׋�Յ
�j׶]9�ɿ��֏T��.9�c��W}�@�6g0�����b�-RPX�;�G�����R߶Uh��\�BN����b�[�1\!����]�f�9C��`rN�=��Y�y&�KI��n��+]	M(��D
�W2'٢�K�E�y�_c��":��$d�.$?\t\�D"ǧ�ܳ\g�Ty�21f���z� vF�$�t:��4'h���dWj�]�J�s�f�5{\��W��<��vX�f�z��,T���D�}+�� Nk�(��/_�@?�a���`2Ⱥ��*f��[���s6��Մb�$͚R�q��p��J����kҒ���@�ɓ�����H���U����ȧ��l�%9R�Թ�)֣�Ү9����Y�U���T/W�0c+C˫+��eG1���l�Jر�V����>��Ҙ������\Ǳ�3w�=�����I�(`���6T��mA��6����OuZ��j0��i��tNQ[�k%�aye�3�֐Z�3\>F2���k�%����UVV }��am��Qã;�_9<1G�婸�Zc���P=x������X�ok��1
t�dc��Can��Vҝ�p�T���i�D�X�$�;R$�v��'P�8W*�=��LpS�d��P��h4�w���	��7m���� ��	x���Z�8�<��4��������6w�=X�L���i�uN0�nBV⠊*��J�T�6�
���!�O��D��p�(������n��駦P+,%�����֯A��2�ͭ�³-y��y�8�Ң�/;��$���c�lZ��|ʞ��;���E[�¯��^����{Y��~�E�]��z� �<��]c�d1 jqO)�q3<x��.�8v������K�-�� -Y ��4sर0���]�.|rG�����dqpy�d�:�<O�� �qa �ގl�,ܬ�1zSg��w$Q�� ?���L&�|?���4x2�F
^RЂ~�����/�_���hсK��Ok�2�ݤ�K`�� ��'�%�=���n�-���
�Ԝ""�1t i�����r�&W�n�\�#�yh�������q�5�5H��%��o�ᶶn���9[-]�ULjmC�{�]K�@�>�NeG���xB���y܁gJ�ߧBk +��㵑�/�l�?� �#�ƅ���)X��d�b���W�7�^�>��8��Nl��R�my훂M~��(�� _�@��#�:j���]�*R$&OЪ���Q@�YɜQ^9ȥ���}}��e�L��2BA����9m�v����BA� J�:̮͗#�դi�,U�S����i�n-�%�ot�]�`-��jw0�"+`�:��V����h�`��'���TJ��ú.���Ww��%�͋�t'�H�Tލ�^��˓������*�5��'I��n7���΋���[���4Qv�Ř	y�wߥ����z晥�]pS������#�����JQ����$ڱ	�G���%���F�M������G����vI������ݯ�&��%�I�'�Nލ)V��aV�h��xQ�0�X�yp�=`9�∬�֠_�"
%.0�9��6"�2�,�|�U��Η��XA�~�1bRyBg�N��q� ��;e�$����LA0$��V�1������S�蘐�7���L�p����������$DکN� V9U+�o�nz�����Xdn���ʉ�/���>�
�U��m�韫�V�
�*��<[��z� �H}��3 䇭M��ub4W�2ڣ��l^�^m���k�2����~�T�q}�Cb�¢TG�'����ʖC�%K?��(�Rl��`",�ʸ!���I��$)�����h��,�E�W��ͩY'i���"��aL*g(�і7����[�S�>����F�v+�V�����`凶 �;[�k�=�e��G V꣍mʷ�)�*�^rB�eh3��)ഊ(��q��3���0��r�ށ�/E�˛��9��(�(���5l��V�J��X�/6P��+�P�
�w��U��w�:�_��wڥW�Y�2�� !�ׄ�+�5�<	��[	X�(q����9P����A��oK��=j�]�� W� X��s�d��UdV�?�	��*��`n����#�R�!#�v�,���+��Xu��6�S�|�w��.A������9m�OD=��

�O�a� ��{���t�9���-��*tۡ��
C��Tl�����F3J�VnT�����x�]ji��\^ퟚ���tdqmU<�8C�4]<�|����p�d78~�UƱE�Xu�O����Ё�u�a��)��3D�s���p��;ul.dk�R�z�CU���M������,�����[ ��c��5��9��Vn�譛��a�b�Y�B�F~�j���4}�n�EƢ5k�`���xB��{�͗���׈�{RG�C&�����m�����)ly���%�ff�t���o�CR����D�c�$� e�󜯐�i��� �F0H�:��D�.�7�&�]հ��
��ytQ5ΘYU囫 �8Zm�Ԃ!&��c����Gn	���n� d6��)y9wn�V�?ŲG�q��}���V_���#$�H+�g���1�������R�Vg8�"����r�^�**�A�����Lf�F��Sv�Kſ\�+�u�7��=>1���]��>�pR�+����~"tR�W`��/��3����ٺ�ׯ�P�.%s�8��Z+�&�)� IV�5��m�[a_턍�:!�g����[Qm��ʳF�O}V"ޫ�Q11쯐aC�rJ�zÉr�eh�@�f5�����?M�"��[����A�i7�K�8%�p1��&�N�����>�+��6r������YLM��<y믉h��tT�R}����3g���6�T�?$h�ѦZ��du$ME�@2���Rn��|k�Tp��@��J�xޣ��u���ӆ��=�r���}�nH���9Ej�=��:����eF����
�������V5�>�<	�2���l�M �(RY�,nX�T�lpec���x�Q,=  �6N^H`̬6П��@��a��N䃜��7�z\C����me6��B9b���!��yȽ3A�3I��9����9GX�x]5���1:A�ѹ���y�ɫc���8Ű��S	5�>��yի}�j|�np<"��ƙ?�͕̏?�����J�|�]���Y�R��u\���)F�ah�!��^=�2ݼ�{��D���]�����6:_�B>W�����Aj��P��'U�>��:1��?�C2;(�`m���_��ƶO�h��S'��ɛ"�A}�����ь4����<��/,<ע5�� �ꢂO�o��� MV��ڸ���χ&�(X����|@ȩjX�?х3�T�=�����u֠�1g{�iu.@B ���d9j�遖�A�sx�w�Z�[kR$���'-�=�W<й�!l�Z0��hH݅��f�i���0H���(w?.�r�	]�*/H�R�@ט�o`��h��|݊X�^�J��rL������ؐ]%{(#|udS�dg_p��/�3��d<뀧2�6�:f��
�%�������-��
3�Ѯk����6�t��Td�!���눴eJw���H�g)�2\Yg�Ӂ}�pp��؈C3�/-u*�������z1!Â���Yyl��KaD(k�I����S�����@�#1,IPE�}3ٿ�9�^��g\���i�t�Eq���]>r4�D�_��K]��1v&;U)�I��X��Ó�`<�*�#�sД��k��$mߤ��l�����U�3a��vj�i+A(jd�;�P#�z%X��꛷$n���PG͍ulW*>�latHô�E}�8��<C`��}�\�F���kl���=�����HY��RHtМ�ѓ�K�:�W���/�sib�5�Q�����l�}�]�U�9�f8����l�G/y8&���uf�����W�f�1·)�2�d�^°���i�=oh��g���;�i$�Kb��Rj/��9·B�\i�VN���| M��@�|j"m���T��X�����2>&�s�|��%#�$��951��z��[��c5��Ll�f��t��2������ð�酟Ыq�x��J�	��-5�u���޷����G���f>��in6�'�U@95��S����8�l�H55�5����ʍؙ��UCnC���S���dWg�ŧ3R��Bٽ�������C@��j����]$���Z'N�/��:���� 7��0b9y����_��u��'Q�A/�i��HĦ��uwIݠ��q�-O�=�X��ۗ�����9�[����]�2*�y�v����n�����a�?�<F��d/��2X�r���+|��P� �aa3K����@ۨ&�x�}���ns��Cxdpl �ewDoX @a|6	��E�$����@O������R�g�g���D��9���Hh�LK�����f���Q�e01��~P�b����vZ,9;��ن��v�`�(6���a��s# \YN�����b�b��`p�5_Ҋ�m�p]��pp�y����}��!x�5�m+��oQ��^��փ>X�w�1E\���ί��A�v��!F��㨟�2�U>W�-�� ��sGq�S�:�.���t#-nY���rv9���㴏�ب�@�?e��?�/���6,�/��@���B}P�rk,���9�dx�����{W�TT��Ȣ�������Y���*\l�%�t�B����[�����ٖ��g��1\�1�︻�.�)D��c��S؀�2��0tt�u�k�8�V���& �
�� kA�\����^Z�8���)QzmΚ#5�d76��O�����8
du1���~��cG��A/�o�$祿�_}Q�K
9g�W���;��!8�c�#���$#(����^ܽ�v���7J��,� "ܖ�{C�5��@��ZϏY�1
�jW?�O�� ����?�1;v`��=�lE��z��.����7Z�f��,�	?jx�F��</�)�KLi��̳�c�K�X���9QQ2���SgEƂ�;��M�pl!g�C�W\��LM�^�K��DQ�����yU����Y��7�{>��~&�e��� d�����/��d�]�5=#��̇�&>�Z�гo
�Җ�U���CavXtSv�$vi�����~Fײ	�������
��J��3�u�,ž�����P �M���G��ˈ���n��go��_UaN�([�l�jo�xwr�Bc7�������{�5�(*������g>�T3ď$АحCR�f�D)��H��YyJ�����������W��H���C�g׭��	� Da�߻ ���1D�A����&Ϋ�w������A���Pte���̍4�������r9S���>��!���	�7JT�R�ZA��v���a��E60:1Q���� ���kegb�>f'GU�@���e�-�L63�k�8�<�X���}��;	��x��6A*z;���)#K���06_�N���I�ٌ���M��1��Q����8
G�sٮ��_�Җ�ďJ�]���3���1���� |�`qsJ�&�Z�Z���9ύ��J�c�5~e q��ߜ�Ej@�>�����JKS֨�Y�;)�GP���AU:��������>��5�[/��$�e�������>��|H��L�z��(�B-Q�|����hyb�F�D�l-r�(�L��k�^L]쳋{A�\�@���o`;�,�u��� �����o6y�ڮ_(K� 4�I��!70eP����G�=�3��f[�٦�^\��ovŇ���&��_�,����e% � �d����F��%���֦��'s���0PV�FS�׵�e
�g���x�T�͘��[L�d@I
F>���xtأ�o�f������m�� �D��pE�G�dZ�"T�1���ʼ�p9s*q�j��Y��Ě4j���QH�q�"��Wck	ڏ��źmakJ�UlS(�)�<��L&�_.(==c!Z�d ��"���QYb*�lׅ�q��T�t���!�.@nM����f]��[e��Z����"�u���w]	�@v|ɥ�W3S��Rrÿc_�?3%^��X��0�Yz�~����5�^���n�bI;���
p���p{?
� ����A�F�2�idgŬ���@��#�a<g�p�A���{0JM 9X��ۄ��.��ڪ<�ؗ���O�
m`[y��i�����v~������ꧬ��(�4�YʑW�Au׮��p��w`�z��(�A!˴jk���%����O��Ɍ��|\]q��O#��{��#�6\�ŏn������z�..)�a w�0I�&��H8�TMRpF"��%G}���ݘɓ���֣��"��~x�q#�g�]����u�HCJ��9�!T�l����_"�_�Cm�:}�Q{��;�Ҷ񕸹�d�h��4-�D�A,a>�������"�����Qm����y&4)X�]]M�.��`Č��qN��\�A?�2u�9c[h���\L?-s�\�]�V�fq.�m�嗰$ź�T��9�L@,�b�j��3y�4��������	gS��rI߄>��z4�J_������{���j����-=%0�ryQ��{=L�6�)䜙6�v�� a���e���E|�1�iĭ��ZMk\fN��P&1��M�{
e�h�zi� ����PD��!�<q�>��Z.��\�[�Z�*��}R�$��������h����_��V��r�l5�*��q�z��k@�n�p~���� ��W��r3����J�{��$���k�NQ��AU�|���^@���n�
b�l��b��uP�ɗ@����W(Xռ�ru���.S��u��5'�tH(9��FwW.~n��4[UK=J�O�Fd�.��]T�|���vD��_�%���kl~ۜ[��w���a���\4I����4^»e��g�(>���P�e���3�|o ������5��@m���wF�(� �JX�뺝�v?}8�7U"��:��(e��P���ԑ�r%cFH�{�7[̗f����o�1�����dc���i�~��x�p�/Ρ�|�ج�?��GVtQ�Z�j�'G��U���sm���=,'��CI�va��-W3���T�*���b�-�py�_��p�/�Oɘ�\�Β�r"��sg�㻄n��n߹S^f�pH�P���N����,��̓<��8��E�r;l�*��� ��MxB�h�Q�2xCT;�0!��I�x��6���+f��*Yt�p_���vGM[,��Օ4�9��9��A����H'knu��9d���O�����9$W���OT���߳�z<c+��'��"-"���v�,����X��:�A87��
y��tș�$:蓐����%�۪)�����07�@%�\z�,�S���[��+�X23^Wz��l��0!�.�C�vC�	����&}���M)��|˝�3a,P��e�AK��-���K�Mϲ���	��P$-��n��H�p�[�@��P�l9G#F���������)z=��T0�R���=�x�v�jM5����1Ġ<�&5Z�@�~Q!�x �m������_7��	|�)O�`E�x���!;
�� ;�]�٭V����po�Հ?T� Y'��y���Y���k.�.��B!M���w�[BE���[�����1�ΒY��ZB�Bg&u�G�U1`��+��+Ã�!�gzKuO�����\H�p�韙m�x�U�D��ؕkF�0��M��jʋ�k �_��گo����2Ps޴��4�$5y��5Ձ��D�X"�
�-�hP�9�ǎ�"_\c�ۧb�O���2�΁�B�̍9�u��+�̩��<,��<B��$��Fe�+c��{W��������u�O�F�o, %]��7-W�Z��3>b����?�~�+�
�~��ɐ%T��u3:�V|İ�k�>ʤK[����^�?ȅ阯ZV� s��ASx���V�[�/�äu�����D�RF��s#ˤ�dG_���-Vpeu7������	�n�`Ej7�9b^S������<=�˔qi*�����+Q��.�������V�1�����Ϫp�\�� �wU�c&f/d3�"g$�����Ղ�Y ~Օ�(.���?T�7թ�D��*�L+w�9�+�>i�"*�x���4ŬOoK��@�hAxSj��{v�N�E~�@/''b��b@QIH��eri���d���#��D�u�����71^� ,���Մf"�Ky0��WDX�n���)zO���n��po�\Qf%�����.��=oh��͉���;�Ir�@�i1A�:����ZSP��c���1[*�� ��������5��^ǵ=UZ�N��MD,	���~�D��@H�5�ЄY���,������7��C���'�9��M�a����l��� �
�����O�����QY���Ҳ�b�c���?�1�a��̣��u�n��%"<�����.)B�!ȃ	#<)��7o�cJ�����֪_;#�>{�CX��V@��t&��-<��礍!X��#)�$I�G��^�ŕD:X=�F�z����hݭݞyߩ�X�>�Q=6����q���L@�6���6�/�9�oV�Ƙ�	��БE