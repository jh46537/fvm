��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $Wժm�5m�ܚ0Y�@���W���[@v.ZX���B�n-%L?]��{�{B�k�1P!�5�������l�pE�X�Ս�m�h#�26�`f~7/ ��5�����`nB�/���i�/��Ip���M 㤱o?.M3��w���2	��� ��:]�����gzpW�5��a���>1���"\/����)�4�◫ͷ��0�8O�6$���i�vK@ ��:>�Z�>8�ߴ�8-�Q��	��������u�݀�5���</����>�S�1�������n�����!� q��D�t]oQ0�"F|y�P3�W���Gu���曐z�nj��n�b[��ȜM���7_�bF9K����GE��R��FY��T����Wxv�������@��"$q!�C*����O��.i�fS���?b��|qkr-k�8ns��˽k�}x���p�#��Uf2�k}3�6Y��7wD��"�F/�� :z��c��3p�	+S���Ee�����Ӟ3
�Y#sAԜ��1���WK��+�����^Ɉ��hRC��B��G�҇Rm��:i7`e�i����y���L�c��#qn�W��W�D���?Rg#y�<q��/1����v L�%h�%mV���:Q�����n"t#�x��j݅�Vv�ؾt>�^Te�0$A�S1>��{_Vrl�6���l[0���u����
�_e$�>_M>���F
��g0>����i֓�fX�%B۲�(�<	���	��@О��f����y`���M�o����3Q�>K��)�O�F�R0�1���9'/fೆzvE�m"O�M|�2�F=W���n8V�0�
��&��2MyO,�W���j��J.9R`|m�4eeK���	«�����<�3h ���� ����fs�>�㜣�{k�kG���������HP�Ӥ����,7V��ݞ��3̳SV˙�,�l�W�a��7�-��C#.@����'L���f�^A�ד�� <|�+y"��qDMA���d�Hv���!��=�$���8�q�� �����A�+ܙ�����&-d�⁧v�%��<T�*��>N��m�q�Έ^��Sf����~U���m��p�gJCO�o����G�B��������r�oQ����p�Ӥ�k��<����d�
ƹ;&ٻ��>J��`����"eG\����!64���MQ�8	Ԥ�xm�%%"�Z�������ikp]���8T- �L +#,���-�H�H)�s)k$9���lٴ�qkV��y"�̭VC���-�����*�1�otn��*�ǈdc����ţb�^ �;�1��-�v�QR[�z��?���X=�f������	�1�b�r+MI�^�3��@�[��h��PUKq���%`�-3)̀�mfC�җ�yf2GG�uHE����x����ፖ�o�����Ӕ����|[����vH%<Fzr3,����kB"�a��Q����-�X#�i�WF���6`�]���h��I�,9����Ez�,0R�w�Z��uf�/��2v`��Z��d#��.��K��