��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&e���g(�N�A����_t6P�N-v�l�)xC]����,�sd
�L�]��bSUO�k�q-L��6���x�H�+滑;_�;�_?m�oǮI����x����KyA�@�\�-lđm�L]��u�g�f����}�e��6rP�R�2��w$F� ����_��E�<�o��&	�^Z �������Q��v�Mϵ[v�s�4�R}��e�0�\�)"�����m�,)Y�[���:���#���އ{��:$�]���A�k�׮�tU��t�-d��~�o���-*/�N�PIq���\~�s3t�U����җ%� T�sQݐ;�v:�?���b������l@���}�_��Xy8 ��T|� ��o&�pӠ�Z�pw��}���4�λb3���7R�����}����?}Tf �0s��/F���� �$������Y���f��K1�%��NXR��3�`Ѯ����ց��G�:���-m�[a�~��9.��BE��H՜/Ay�[^o��lh[d������ʀ�m�7qf�m����I�����6��Ŋ2���	Ԥ���Q�Kp�È��	D�w����3�|�3e�M�)p�g4�U�܎ڀ�{�0�a-k���)�������{��E�)�]�J��0�c ��(ũ���?��P"U��w�QWc��D�$����>H�¡`���T;�r��.(	\s�#��0��5������C94j��H�x�7�*
�7�~��A@T��CYY�{
�H�ܦ�e���t�í���m�7W��� ��i�H��X�<�rړ5Q!�o�F$K[��O;�?�W�7+[��A��c)Щۊ��Wr�#�
�f
+������f�iH�>�{]9���T��چ��`��fF�(ۭ��l�W�+lU~X�"G�EѰª$�j+Ɍ��/�ŚK�hq��sEυ:�fe_�oay;P�����7[D̅�n��b�ć^�Nk����@c�}����pfL�.ߦ�� &$�\@*��do;���*F",�@s0'τ�3>�����	P���"�Ҟ`�m�Wɺ��&?�[g�1.�ը�a����nK9�[Q���ę��a�`����&W\��K{3�`��B�݀"�l���WMQH��a거�<˻���r_R�W�3�P�����@y�����o(���u���Yw=7�Ⴑ��>N�����d+"�2Ϻ��������ٟ{t^���(�s͢"[>�>`�W	n$�#�M�U8ն�g�����ʞ�,0Q9"�i�H-��X��A(s���ܰ���?ȼsǦ:��68��U�����q.��86�S���ˬ�����ӕ�݅}���1�����y��= 1<a���WM�,(��X�ʹ.'{Ή�<h�w�R-(&v&B��y!Zw�T���FAw���C?�[oři�s
�s�8�jƻs���Q�M0��>hE���c�$���(F�<�c;l3� �:���K@�TC�|<�E?\�����[p�XqG�R@���ԣ�[Ӏc_(N�9pw�I������n�,�M23����dnb|R\�u՞#=܂�fV'�җ�\;�{����^D�9��*ȎN%�)�Ż�����I�� 
vc⊾�@�����N�Б��vG���=b'�'Dq]z!�l���B�[Z;�&��x�}��{0Y��{�/��uF����Cc���m��d����:����^��Q�9h��+X-/�oTPa\�iPW�6�+`_HeP�K*�����rzx	����S'K$Nj8�<(u�!��t��r�ȗ̍�h�T�*$�P�X(ͽyj�x�j��dx�k^c�W5}"va|K/�;���x�2�xEg�֒�u�L{(XQ�Ӣ��0�Ѓ4����'�I�(�r_0����H��l�