��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B����d��:$�馈����Vj P�d�r���rO4�`O��A��4�k�Q��)k���E�Z_��r�Y��C[r2ҖUg(���`�S�L��Ȕ`�?"F^���w�r������m�6鿜�7��~} �(Ĥ�n�Pe��	 �cE/�ݭj]x{�s=�Q�BQ��T|��-.Q�p��.�o<��A��3���$���'9��	�"�.M����(s��?x� �'K�S����� �kfI�Ntd�J�G�1Y�Й���eRo��@�*5�g�!�M�l���f@�1�&fZ�S3˶凨�_����E�2q�YW|���"��,w�	L���J��N��H�m�rc�O��k�#���g�T	�@y���c��v�Vu;O��h�ʆ��gi�	[ƁLT}[,�i�,�a�WC�׸��Qf���S��/�����|�c���{��xI�;W�_�����~�� ���D4�7M�`�&��R�$~����R`:]����*���>�O�\L�}|7s�c��&��^��h��P��n���2؃/�s��8�h*�"�c�D�%����Eȝ3��:�9�4�ыrb%�ҿE�i2J�[;@�(H�z����2��ڂ����b2�����F�նmk$n�Q��O�GB>�V��(�B{�M����CN9�W�G�a�Y6�>x�����Cz�]��>WO�ːu����!�1��A5u��jLŊ-�8�(|�T`��1�>T,�Z��%~L�����
}�!��&j֤�BҐFw����Q�v����tNXj'-~�$�
�翾��*jR�D��;t��4͠���*ؒi�I���{%�On���͡"$��7U��>�D��!'�_�@a}�B����Xгq���5�`Yţ���zJ���A��+�q��b�6�����ÏM�Ŀ@K?�b�跇|�-�!�cu�\X�/p�I��J_��������hwR�C��ѤT���֔&�����!�Lŗ�<-����¤��hu3��	\����4v%�t�6�Bc����S	zqmt>#3�J��=m�i�:9U*�o.���n?����vN�o��G3ų�V�D�:���R��Z�;�^��(�ǡx�%+���ݪ8R�SwX�~�ڪ[�P��3ↄO�������{5	(q��`��(o��cBƌ9\4 -9�#������N%���陾��.�OԜk �7&k�]���3t=Ә���I=(���Fkx<?�(N�8H]�!:5�D��/S$�Uă�?++�m0'����?���V7VI�e!%�L�0�a!. �]��q�'�,N���΁��JyIo�:*	d�����'�b�����t�.�Ja����[��t���U�趯9I�S_)�R���� n����,b�C�L@@R��f1��j���R�f:.�:�BYJ�,W*^���PP���(�1�ȇv)Tp���Wli��gP���_P�S�?�T^�8�|�8y�8g�s�����ݤ��"�z� u�X��R��r��=�-$�$S׹��~�hS�v��(�Dr�w~���9�>�;� �z�9�An�$�k�к��>��S3��~T�w���\wŸ��a;��WX�O]hކ4y_!� �a����[x�� ��x��`�8���/_?��:�r��Ot"Zj5��1��	�vh���@�O�F��H�/�4�qo�h�ud��W�>gv����dz�H�%5<�����OIt\��ם؋�l�Բ�Ft�>O@$�	m^X��\���vm�:��	v�^奛�֥�fj��E��!��-!�ȧ3ǽ�f�T�1���n¦L���!��f��&2�k�S�R�8JC�#��'���$)��R;nj�+B� 
�b�4U�b����e�-]�8/=����Fb�gr�h��?��<�,��B^@���\]�
d��*��y& �d7s�N.��7ܩ��9�\�$P��:* 3��ɳp9��G�%{����2FJ�G�ep�U3�}@�I�x$�Ԝ��{~��!tzg�Ǔȸ�˨T�6���/9zn/�i�J����7ʱ&� Î�eEPxw~�~ä2_3|�S�m%bP?��;A_�j��h�A9,@-$>��df�zG��{O%�Q�ײnkb��U�[�!��s����4��������&�;�$�ԡ���ѹ��%pT{WO
l_�	6	�S�Q�b�%����(j����MX~�㕂�R�~��J�M�5��mM��u�w��;��tiD���QBŬ=��c�3�H��c[�2�CB���Y䔊	���}sW�?#<��N��_�ω8��t��R���C�J�6ԝH���{&���<�a�kH�]kXԛW���w����!����A@�ܧ��D��zp8�)lK)�K��ߴ_qe@Y�Q���KA� vj��J���I/�hm������&�@�2/��/Ng]�r���]@�aL>��I�h�a��OV�4��릱��e�p��%�s��y!�s�*ڇ�U���%������ߎ��$�l�u�瀧�VH{ '�mc��.��b�bx�(������vY���'V�"��E��\k2[�X�6'�ΦB)�V+�����o�)? z����ݼ)�'0ʃ���ɺ> m]�5���w%������!������C��	�l^^3��Y��,((a���7���4в@�k��f��S�������C�%#��A�w߁7fS��~�w�1$�|=K���i��C3���~�H��;
j:�W�էz�o!�ɾ�{рV���7��Ӗ�>�~xF��$~G.Z��f2���W<yyG�O4��X��El
�2���e� v��~/	K�\:-&W�b(��s_��ʐbؗ��g,��OY�O�9��I�i*�f�ٯ�.�/~.�E�<F)�@��w��bBʰ;�"�ɜQ�bFdޫ�C=Q@��e+�J�?J�Q��9��>ܵ����4�3��Ҽa�o��B;!�`���Ōз�w�Y�r"0��'c�{�+@�a{�b�T��:��0����h=�������Þ�s�I��V�AU_���t�.�tFcJ��t_e_8�*BޗΌ����^���%��������l�L8Y9'�{ˀy��@��\�_�Or�[m���|6����^�w�\�lY��ȫ����"��9y�=J�먨��8Q�CE��������qTZL���	B_����� �qb�@xl,�L�-��5Y]_����K���.8�N0H�q�v�� �-���al�r	$�.\p� ��D���,ő�؃:Ev�9�f�"e�����¶`	�}��d��F+�ֆ��?+�:P�<'�U�>^�����)�wB�no1�^�31)�}X����&����s��d�*�]j9�Ǹ�X$��XP��T��=��;��(��zL��d��/uq��?>���M碨�>��^p�㙛g$��)(��@��1f��%3V.�WI#��0eN[X�n��?|�Ky�Y�?-�^q��G|�؟���͍$lf1~�ǡ&8�<xg�W:P��qn(8�B
�t���
�/�ܲB̅s�f(�k�v*����T*�R�h�������>��:.�0���K��A$=��^�ܙn�)f����e7L����;9����G��;��z�Q.R��IH	�o۾�#�����G��t�Ӓ�������n	�a�� �����c�}Ʊ|�z������%�,3�w��0+3��Վl�/j����9q�{�Z������5����x$.���]y��!�TqhDG���G��4AH���]����r7��{��-//�� `���4���?��X0��n�/-l��SL�{Aa��y�����
��z7���O� ��_'jzl������>���٘I��Ɍu�E��ޙ���o����J{~��> ��߾B0]Z��}�H?#�ƴ鍤�6�dl�o�.X<���&^䟗��_W��6-�Ȏx=mM�� :����\����O��:DQ$+�V��ktgJk=����DM���#���a�+�&�L���W��ǖ�]΢P�E�77���c��ց�7
���G{�w
��W���A����  j>1{����'	Q���'عw��H��D{ͨ�	)f�������>'ZZ�z)<�ڌ��w:����;t�+ �Fj��4��&�I�;�%e*>���z�&�Ġ�1Ux=��_=[��ew�����&0��1e<Hw��ꀨ���NC����Ϊ�ߊ"����_�VcY�ک������^�)�%�hi��$$W# ��>���£�����6��(��\өL~c03уN����z k�m�~qE8�?z�Rp�S�GW�N��=��K�@^��	9Ӷ"��(��9�un��"��%� ]XiFӟ�zS�o�>�w�Kg�#��v+����v#��NV�^Jwr;כE�ɞqxI�ج ����j�u��ǫ攽�%{!��)��&[f�^#`ہ�A�e��ϓ3����/9�!��60��/�d�U���c"c|iR*R�������k�
縚�)��	�c�2b#�@�kʜ�`��EM뫗	P�,~O�gḂ�_I�?�:���V��Y�M9LNY-ROʀ�aA����]��6�ã�w��ir{U�]�L��bH�s���6%�4�X��M�r�҂���Aq��|j���$�jdƢE4.��.c~+�6F�\�ǩ0�u�s��ﴵ	P1~�V�߉�#>��2��ȁ&.�<A"z���:�I�ZX��<,0���� {�S�t4I,�E���N�����ŗ*U����J�7xGbT����4��a!���ꗡ.��Z�-0�++8��I� j]9~F:�>��A�K��d��l~�� �����2v���sEZ��#"��^z�K�l�^��3�1]OS����H�UO$ҿx�E��� v�W��|�#߽t�>�(l��G^]�z�s���S�V�m�_D�W�bfDq43w����`��q�@{:G�g{b��6�vJ�'u���hJ�ǓJ���Y����^����Z��U	��e��̥���B��/�]��_?Ȼ�I#)��� -���<���Riɮa��$�ߚ��~�D;t������72�W�5�,ӲϦ�;�}t,o�	f]&J��:�� іT�Ci�t5��B�l�U��LӧR���0�?��jW���"Ao~��ށ?qY�Q�G(t�_�*�:�V��$�ۊ�;rQpE9(��`DmQ�,�|��b$��3l\&x�(��>�8q�E櫾:��"�ݮ�Y$��Z�ǔ���SW^��G0��������+�K'��%��Ȳ0Jr�a�0֌ޱ}�����|�Ƃ��3a�}�[�ώG�t�'_�Y�����I~e�p':6���֩O��Y�5�s�O��3��"�L\����3,�9��[�MZ,�y4L��_Qۼ�\~m� 
n��h�Wv��!L��"�>y1k�~�/�GXӅ�lK�]�-?�_J����*��b���[������)��G*4�nK�QXrDDAC[�Lk�������YRkδҍk?)�$��ȚK�Fc7�\��:N%ߚ�
�ug��5�1��a�PH/ou�HK�M�e n�s�:�,2w�Kl�g�6`R�i�i{k�����Շ-�O��oȠ��Z�� wqB��QdA-idL]�n;(��9Y�6JO���Ůj^LFʽ�)�%�6�fHϻ�D/h�Wg��)� ��cJ'}��Cg�S`W�:���@���O�sY�;� �*���*nk��Y�T�ͶA��wP�㤚�p��St�=���_�m
�|�=#�@=q1��:-f��R�5������y����ׂ��
O��_7�,���Lk��x O�?|��0a�pP�iY�A4��P�X��-PC̟���V�v���[��E��wsP���^(Wr=���,���#�}���X.ވ��b�Ru�r�����N��Ԃ[1�U�I��",@��m$h�I|�Ɩ>��4 :Cs~���o�C�����ǥ뿧Ư��%��Gi��{6�>yUDC'��T��)cj�I ��Qƌ	�@"u^�?1��
j�"h ? N�Ma��j]<��r;ܖv{�4�aҭ��+������w�f��ݸ4ƞ����_�Y��R�����~�m��qM!m	|�,�^F2��L�cPd�A:���p�ÀQPKL�$J�W�tx,d� ��``̖�.�ZQ��k��~`����md�_
��Ǵ�<���U��ݪ6�Ԑ	�:�"��<nORZ����������t�W\cq;�B���7���Vm8�)��d�3�M�,�S�}۳L�v�F#���7� ��M�g�٤]��CKe�^:�υ�1�GЙ.kN����>"?�WR��8vʍ����oJtKĺ��A^����`;+m�g{A���Y�U��?X%�~>�>$��n��G��,o����\�Ot\�zYKg���Duy��"���2��MB�h�c�@؂�p�|L��6K�t*FGQ}����] � ���3���ո�k(�A�ǡ�^5�����Lc5�����T↩�����;����Z�ULA�^��#t[�N	�ń�w-�q�=}���a������ �y�S���˴�{��u����{#�.]�ϢM���7�E���ݜ�7�zR��t�M`�W��/T��s�DB�C��e�W��0��m�J�k��˾Z�
'�pz�:��ޘ� �>1���h2+��u3}�ؚX����@e��p���]�jҥ콭��yF"J\v���
֔�O�`I5���n9��s��T�%LorI�j�,L��*�)�Q�C�ǽ�(Ot{�[�TS��lr�Y)�~p��D~õC�3�A��?,���m��4����N�&� 0S���W}dh�5�+�m�A?1��7h����h���}th�\^Ѕ�/�㰯�U.�+|����:Ö�ur�f�O�q��:�����v��L�\t�G��&_
����,��u�|���U)e�ַOu��Z�
��r�f�|m7�s�8r�%����X!4�K�[~#���&i����v��V�3rE!��6tA}T�Qel��Aa�?&k{�t|����C��M�KG_���\W�ugR��&z0�V����.�Tx߲�'Le���6�Y	��`�*�g�n���=���&��V<0M��T�sm���_�T���>�o���{xs���?���0���o��޴�^X1w�vI��jѴT��[|�*=��hm�Jt�3��up�+�J��0z�I^�MZ�6E��xڑF��I`� �F};�1���T���r:N�dy�La�8�m}^}�,L��Ѭ��6�>��heEj|� �zk����I�$�"�H�Fh�&Gw{e9�U�ecO�633�t;�\���q���&L��lJ����b���$s_F;-_cOB&�4`9�����1,����̀��i�+m�����9@Į_�-��֌6�T�6🦲�B������I��vL��b �U��������|W��$�M-�;�K!��r����=G`W�z�C!X��e�`�+IQw�
��Ze$`KA�c�`!G$h�N�������{�#�[��j߮c��)u��4���.)pB�I�L��q�̈́i��}+d!5Fnۼ�3���8A�M&>�؛��؏~ƽ��Q����}
TQ��G�o��w��`\�b�SGb�G�D����"*��~�T��|y9�^�2+�[��ڨYK�%���ⶳ^��������e�e����4����3���1����&��b�6���Y$�X���s.}�qY�ia�31��æUI�7�n ,3�ʴFr�k'���?=߯������:r��'��5��H��C��o��✋���2#}-䔜L XN�|=��� .//ޔ�Y�[��)x�`�*��Q6���`�yZ5eQ���0*�[��g���#��Z%�Mo����X�`���<�ܦ?(�tNڽ��|}���.a�M��@������p���u�}���
������:���ް���P�#g��?� ���y��F�h��M܎���Z���;��%@� ��ٴ?��5����J�z�4<�qTL$dȫ<8�7�����w.	��$H�<1�z㨎��bȽz��Z������]�*��j�7�\����j�J6/���@n��)��/��j<��6���U��|�;����z�E6�boz)2�~O�����)��N