��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���r>n�W��0���g�}�aHzH�[=�/���hIo��:���D���ZǄSh�|uVYo��,xL+ �k&��=r��U2d�e'���#s$�1�r�xI?|d��a򆴋 <�,���_�v�;��U"���,��b�n�YN4�,$�c�ib�Yz�3��"k��$ΧHM[�7���!:6�1�s�_���&F��͈�T��<��T��}�a�y��=]�\'�cd��ۢ+����	�a��H�'�Q�[x�ImSO.o����I�%W{�ӝL��s�>z������ɬy��Ҥ�2�W�A)DӲ� ��*l0V�� �)�u^h,��R�?���&�Y�@���j���$:D�W'Ѵ��R��q5/"�x�
�6Ђkો�p�(�Z��:�A��x0	�
��~�1� �C�E�/�36nD\�t�g��.��ːVK��i>��U�I�R����3!̒����leF|Zr����b���Fax̊$K��~Ry.r�F$v��2E����DӇ�e��]�h��m\ˈ�S������S5.�.�s�Ww�źՙ�=�pcBJ޷kE`g�zb��Uc;�����?��DM~AVr�*��Ӿ�,��\�x���R��D&�5j�AcY��;X�G[%z�qJ�2폂ԋ0S�'��n�x�F�6��T�m���g�>�UK ��!�M�$�>kC_�`�+&*����+F���s|DK��t��� 3Ę/R�F	��;�:�,!S��k	��3T%D�+����W:,���:�e6������*�a�)Zd��G��R�}�Ӯ�a��B���O�j��d�NS>��Z�s���v2�C���u
T�������8��k�p۷�l���B�@���~�ӓ;�'�P�.
����5V�D���Ϧ�dH�x���R����x���O��.KlI�W�єo*~�Z7��3�o��-�������i)^���c��<��&@5��*��)/A�!'��f܊���ꪶ�S���|_Y�}�����#�ƑZ��s�;�{�>[(������]�ԈF7^��_��5/�n�4���B9��]�9��^�w�Cع[{����3 ��#u���t3���� ���G�`=���.ulC]���m�˗��ҥD��g�o�ݦR-�s����G+x
�C�O�$�������I��KV�_T*u�>ῠ�'DL��g����Y���9�����r�-?(.E�	7^���0
���.\{��S
���肞�!�V%�1�*`��?`,9�nXw��;�QZzJ2��;���$����H
��r&��+�� S=Bown`:F����_����f�N؅��p�DQ�ܺ�$�n�����f��L@eَ�R�<=j�Z�ˍ����-Bx������$�[�k�!ۯ��9b�g��B�yw	�2���$��-Z���j�4�"*���s�_
�#�X�������e}7dL��`<z��<4�;��T	X��;:Ŵ��]�_��1M�^Y#L�w��[S��{Z���
��1�%�Vv<RUL'G8���E�Gh��q�����d�<�ste�mZ� ��\U3~���5b�z��	W���@�컇K�/H
�?r�\cb�r�����k��h����[��Z��|�� M-}T(�
��,r�6%�3lշ"`���CPHVNQ�К�R��-�4ݍ.z0�}o����/W�?�׫ش��l{�h�Z��t����q��۔���ۮ�wq�4���0Z�fz�'c�h�@��B]�\�O�l�u�E=;��q�<k` �"�hu�x�N�f��9��cJ˞[�(gb���X�4!�As�'��Jw��|��8
:���R�.���V���̼�t@���Y�#&��)���y�)qF��$U���%.�zՂ�����4C��u����˽�=�|gn;}�P�v�Gt�znص���i�_�[�g��0�׽��L���o����%N>��ڃ�p�23���"��@����U��s�'�ث���=B$@|�d�;�B첓.Hk��"�wL� �g��LR��V���SS�������(��e"��(O���v�Ҹ)�*����x�y4ǥ@��w^���%
Z�C��5��Ĭ�B�W6��IX���=�����C�*�C2�@��@�U�(7�)�lhb 8��9k�V��vK�Ez�k�#�@�!��]���]&2�"�
W*������|J�g�AL�`�ڬ˧д���8�=��s v�Z����$�ei��;(�D�[{�Ӛ6@L�W�^j�3C��	��<#�R?Y�p=�~`�9
��l���_P؉�ܻ	xTKZ���n4UT�� ��:5� AgN��u��!\C/n�Ib����>k)�_ �Y���'��@�z����f��S���yH��K�EK�s󞲺�N�F�C�_
��L�I��B��r�wa�|Y%4]c���4H�Ǒvc���j��u�P�Kf�f���y�Rj90�O�`��y��oNt��-mT]�q�{.zl���>C�b~;�h��O�҃S�����׮�n	� �`�+͙�g����7��S�X�������=����bA��qv�6��E��j��CMG�� A8�C3���kox�pab"e�Jό�����-�n���o�����^Ͳ��mm�q��Z�Wܵ�>��>�A؟�6�;cg��.n(*rJ�*/�[2hፆ���V���5o�*o*���(�b���?�LJ�����=A���X�2��pW����$��pC=�x��ʘ���B߼�{ٓ���z�n��D.�h}�(�ѳR�Mm�� ��_П	pSY�@. ���r�ȕw�+*�HF4z����4�����gQ�Ɜ�:YQ:�u�����ܪj����~;A]ըcn���Ѿ��fڃ��:�E��n`#\t��v��"al-�g���^��[[g�2�>i���'RƦ�W������)��ᒫ�'�BLF�C�X�.A!$��|��1������E�� '��o!3g6p�:���N߃��Y���s�o@s�V��t����z�¤z@�1�3��/ҽ���nnRfz<	��$�����8i�me������Ã�R�wJ�_{O�;�[l���3�
���&��ߜu�S�{���S�wT��5�t�:AO�+jS��g��هa�i�83��~�(^u9 \|�>/���.�(Y�����t�FqO�;oY�QWT�ȟa;��#9�� ��I|�]�Tʦ&�e�C����QO3�7[��Ý��Z��~���'���/ �ߠK>rﷺMԎ�ݥ�]4���b �D�)K�hf�]�u�d존��Q�y���%g����y�>��1�=y�ϭ�SEit���������JE1�eC8�ːM����͙�:���{Hd����
(�'��D�2MeK������_�O���+��֮�/�0��2� �B��`�kjʵx��?�d�ӓe4~���e�4��m�d�	U��_yu�k����r>9fp��F����:!�M�syc�7V����o
����-!_u������K�~� /�����_�X7�\��d��#I�M��"[j�����FRR3kpe
�Y��~��|�(��H��i/�d��0hz�;�6N05�J0�A�m	�l�x�ٓF�b�:�h�nr�C
���3���܂S�����u�4Hh����¡�3�g���ű�K9^l�w�n1��o�Zi�K0P*���>�Y�n�_TI�Y�9�'�h�����Y�,ƪ�Ú��K<fS�z4h�e��_�ϧ����}T�B#&�%V��Vg-^�hWp�f��SW�R6f�ޑ�."0�+hgȆ����� "J�갢��������s�ʅ��v���=�S�U�qeT��
��%%��3���o���{�Spr����#�
&9]�	B��1�]����#�3-A3����A�x��f�!#�Hu-�6�G��*y�F�{ɂ�V��b�z��6�!�ܕP�|-I���Eo��Nt�P=lv&>��ղh�G��z��d�NO����`�K���`L)�1��� �O�9�7�3���I������o8c �| ����<���~��uE�ޙ,�a���hk�Z-���j/.9$�8f�ȑ�)�|��^
I��1F� L��n�!�=������R	��n9������m>�b�����:9T߷��$H?X�zb��#�cs���tpvb^+�pja:H�~Pq���p�Z��6"�z��"$�&d�r����{+���E�&K�B�w#H_�����o�ډ_���:O��gȶqv��~���--�Sx>y�AF�;�Rʞ���tA�����y��lĹ�QA{ݥn�Zkߧ��J큺.ԡ�'�!*�gRKx�8U�K�Z�؏[}�L���v~>�v���]�R�iNI�q��nB:�p,JA�E�:f�^la<S��w�^J������� �;���D��_�C��<)S�sc�5ٟ�o�aP�R�W� E~�Zg@J��l��m��s�$�ҋc��0JF��ѩiq��&<�k���2�A4����~�3��:2T���f�A�Ƅy��
��?W�~��#U��3m�zF2YED���%) ^:%bk8��)�Vq�l������H�g/�D�-x�@|fı+�S�G6�?sw3�E�;�;������Ad��1�����S ��x��BSc�葳�������7X�"�}���\5r�b�t�~�|����^�C2�^���3��$,�8^��ߢS!I��'jO�a0'O~?�Q��:�2���={g����r^�<L�{ƘD�ꣽ�sc�VN�F7K��AZ6�%_����#�ۧ	����<���Z+Ѥ7Z5T ���?���6y��T��5dɕ��[��()���*���{N���۶�}�7L���$DL�0�~R(�gU�͍���qr$Zv�6]���5w֭t�RT�8��r
�7꾷w��Y',83�)~S�,�9��+8�oV��N�L6rB�grIQ���N���@�mB�R�H�8��j����9�5��S>����%�A���ͱ�\�?�gөH�w�Z����,�뤥�a�� �ޒb�>\F9yQ�l�>���@���90/��Ʋu�o���'V����{[�>��ڲ�g�ڊ�y��5�R%���F��y���`�Wy;�F@K�@a���8aI�c��^�va�䱌F�Qi��`W��Fϥ+K�nĩ[�C�ϼ_��sg���e�����6�F.�qRO^��MYKΞ�h�s>s��h6�6���9u� �k m�s�*Ď*s���!^s���wn�s/��Rƈ �jc�}\J�א��	�34�v���>���ԡ�Y�C�=-��q�X�'1���_BϏ=��M�U	�^@mF��,m�?|���A��6NF�c��$�iϬ����O7y�q�8-/��
��2�F�*�$�r�7ݠ���Մ�Y�@+����T��4q�=C�`��V�4�Oφ��9&�]���\��ɀ?�?r��{�@h+�}
%���I�.�)��_�V|5�4�z�I�2��l2#�M��X>����/�5g#۠������#<V؍�X�����B4%ށ7�^!�$X�Fq]���I|����nZ�B�'��`��Jj�n��Y a�g���ݯK Ք�'gVЯV���P���ك�Z�q�$��T���E�FC�c+�\t8�R,�9���$4}]�� %���d~Q%Z+��������k�N�t��XV�+�wH�,5� ���8~���q���u����+�C�Lh8�^P���<9����	�#�N>�9�
���oU��|b]w�w*l`!�
G��_�| ���Z�9�#RM*���幢Z@���>dx�����Br)��T�O��W�
�܋ݚ��F�=��p��������>�Jk��a�F<�4QL�t��`'����kp`��Z�����.�ۖ�r������@
]�[��[���p�P�Ġ}�/<�wƒ�e�20�ӫC�ۇ�t&!�T^@�������z��Upd\�+��;�#�/�V����=wzG�L�"(��(]�ߔ��+4,m3x�A�˦�~@����95�Mʿ��쬪  �>̪k�u�)�1yd�TD/C��炏�@������Qq�+_��*/�͔c�P��t�ʀ�:K G��s28�m��a�I,���c�>�f�^S|և�I�8�f@�̓�6Ħ6�h����Y�r�u���Cޠ��_]��!�0��ˈ�٭Uq���k��'��*���-َ��î����)e�L=޿��/���V]
��)o���ܹ:"t�9C����C�|e�rJ��fV@����q?�~F����DJx����f#h�5�@Ѕ�d���R�T{5D��
Qn��m[�Kj�0�knb�@�̆9h�_���&HP��OM��f�ޱ�q8�x)�[Z�[��|ꨳ_ؠ��U'��E*U�M(��|���;>�M�!5�p�=�w�t2��m��h�{ٍ%�������A�^��_��7�8�9��A��55^�\�/��dI++�.�jK;���i48�6)>�e�	�$ٴ�\H/r���E{O��\��t3��@�+}5����e)���|as���*�$�Z����M��S����I���%�9� �D�"�)݁��X���8#vr3Q{���� �i�x*�����W�����-�04�1�Ԭ��>q����k�JZ^�d�l^�dD�c�s�2C�YރPgg<� �zz5�r> �~״�S,O���%V��:l��tv��}�R
���Iٕ&���ݪ#؞VsO���\�1l�AkD�s3�E�-_zfA��Ui���!鶹T!��!�A��}Iȝ�ѭ!�_�����Z3���/�R5�4� � ?lH"B»�~v�kb�cpr�@ʻ&yRSU����!!�:�~��|�^w���5��$6Rb7��a����B%�5�3���S�����!_I�MEQGq�RnZ�/���ߒ=���0^�ɨ�C,ʊ�m�,ħt��=�N&}�w��K��0�PS��^��9��3��=��+�V���'��Mߚ�!���4N�{5��3���ܴ�g06�6�v�-IƝ����A�_h��M�c�D�C�����:E4Nт�P&Y��b�LԳ/�2��G��<�Kq����IzWH�fc���Lh�]�� �b�{��9cD\8 �����,3'61��N'����7�C��1Q�;r0����~*4��?�I�_�<����}!\�b/��4Vs��N)��(���q�B�oG��	���J,�0�x�><�BQ	��[|�|/�OcO�PhŧxƱ7���	V�-�c�Cx(E"NU�c���Þ�ceخ���eFR�^2�$�jV.�0��n~��%�L�v��-$����A�)'�F\
0�RN��eo/rm������`_´�l��Yb�|���z�qѪ*-obzk� �,O�*�%f�J��S������ix�2������3��,A��wZs��@ĝ~8���J��ML>V�*I&i�͔��k|mK�b�o�I�PْHʨ���Q'�>"�ZI��~�W����TC75M*$oz�w�첩���\���'�5����f����Ё�93#����ֆed4L�C�fiNrEgs��f+��b J�ㆬ���N����c`��Y&yz�ى����4Gfn�8�k�ҡ�3I0��U�3jT�~����y9k\��ε���rD��%�������
l����,�,��(��G_�Ә6K��Lb��rM�?٩&���L������~,�^1)s��\d���)���9��[%Ƶ���ȳ�-�Lʄ�^b�oX�I%o�~���G3�(�=�-M�.��ULn�Ӆ�
I�_�i����߸���J�QGI������'*�'���\����nP�ح���5�A����W��@,�o	򥃻������.À������!@�nc����m��Dy�����x/X�U�&'�A
����>�YAL�S���Έ���VPh��4�oJ�����np�7�[i��L�,��΂��g@��g$��w��Qz�5��NX ��b�)汵|�/��^��^_��(��4-��gJ��&q7��ԧfa�{�d��א�^ʘt�o�q�5����' �BT�����!�>R=ĉr�Vz��>�P���m��,����3���:�"�%�mϸ�-"�Z�7�Oe4���nZ�v֑�Y���nS����|w���N��/k�̎����i'�Lf��m�L]���k%V��z�9.�( ��{f�R��0J0���?�ǟ7��dX��8GxUƑ4M��pD����jN�"go �v|�s
w�d���|=��M+wU�;�Ր$0�Ր�w��t��ZP�u�k�>89jD���g�P%�Ȇ˧(ˇ�LZ��4Lh�f���?����lf�ۺ
��{&Cv����/Fk�^�ˈ<��a!ih������;����P�h�q?;�.v��ul�To�̇�ٲqͻ�a���o=R�Z�{0��Q��S�
;��(�=~Z( z�'PR8@�BYsAG.��<����rI��P�mF
�aX��V���*FAJ��u�Sn� �� c�7���~�beT� #���K2q&��l����*lr�do�'���|\rz�]�N�x�йi������$�;��P��#�(?��=K(u�M�܏��TW�ՄB�w��5L�~|~!��L�T�m%�l�B�d �*J��<\�|R?�����1t�DQ�31	wi�b��L���t�uCs��+����$+�r��%&v��G�3�'�"�.�]DYk�ʀ�:DL��e��S
f���&�K"uso���.�Kl��}�}�ϳњ��{d�0q<1��0���6�0���D�����%T:�gI����5��μ��ˍe!-A���my�s'xb��C��Ù\E��Y�6�*(������ԋ����Qc`��-&�0����U�q3�)9?fE�-6�U
��%+R;��������b �l	�<yV�6N�2'.�йy�ߤ���$?��|�*����µ� ��J�qU &��y2o���F��[��������>�h��,.fn�Н6�ͥ���VS�x4!� V���D�V3;"��;o-����r��Qs�X	�ۮd�����=���?�6�vvg��>h5=t��Ҥ�����4�ǖ��r���l\)/d\��;��T�$t�{p1`��m�;��ja����1
6��)���S���JA����b�B�u�U���x��Ŝ 	�0��ЋSPAܲ��.�"s��k��}�m�3"��]LH��Z���@��b�+�y�B���Ak��P��~`\#�OŔ���g�<kIĆ�X{��f�?!g�|m�1nW�.&h%�B݄�����!,`A�)�k�v�[j��j���B+Վtcs	�NpO��߿@�3�Ne[9G14+�E��1+�f�A�j�
�@]�n��ې����R},kA/p1����޲lJ��t���,lJ�z�]��/��`p	lQ�CŔ�����qt��Z���� �@���h�DM��ӭ�J�[p4Eo#f�&��Ԧ�u�"���QQ>�����sdfL��J\G��,��������~��ƒa li
&��o�¹\Ke�.8��álm��=���@���}V�/���X"�bP6C`[���`���9rG�/  P�.}(���p[�v��_�:9������6�WҤ4}iң�|�dX���oC'�,�d���&Y� �9I4`�[�������ps�ؿ�x�BW���V��ߏ<�k��2����)�13�;C[.��ѹV;_u>#c���)�/�&LZ�6!����y�T��K�=��{e0hߗ�|.ɑ���+XCay���eA� ��7��]�nu{im4�W��v��+@υ��]�M��a[��;ҳ��Ձ���˳[� })a}��O�ߑY��q��F��In��H
�@��,��@���������A��x\���X���%�e�����@F�U�jO=l� ��Mߜ�� ���$M��@��h�uX�λ�4�'��$���?qqpδ����<�w��V���>K
��#k���/��cL�8���Ȫ0z�m����(�dg��88�Eo���y���Cw_)�xlÎ�f�=۫�݋�G��l��|*Ƞ+�'3�'��S@䭽TRa�H��1�w�aH�?<K�{�x�i&�=t�=����v���C_��	B8"�cv^ė����<��O7�&7�T��jZ2��%`��o���l;;���o	%r�|�F�;RԱd����p�������1�V��5�6G�DZ�{�QR�"�=#q[��p�B�^�����D�i:���F���M�:����g��_�@����~��6�_� V��,����X�,�t����T?��Mc��x�>7���.��]X��c [�Vbvw]��ܽ���Q������QYe�	^�%v�\R�fsm6ɔEN$��5�~KgX���yu����x���DlJ���H[���V��e i�Ky�1j��lv�}���I��w��� gQ3:�� Ze�4���ܶ!�2a�)�$L�(/��q�Fӎa�)<a��qQfa@/����<�qc�v�8 ��?2e=��.l���0�w�0�m���F�[.c�N]�˚�[ <pl�f-9ɲ)���3w�T�����_��>�"l���5rD���i��#�va��.mW�\l�g;��ԅ�S�+S������.D������G�0���XS�	�V:�A}*J��n�i�{�����P��Q�F	s]�f��fSYfy���+37,6_K�-�#s*��m!��*�q-��!����}��թ����/�V/xN�i�=$����pi����Ik� �c�Ts�_����^��I�������+�E<�q��v��Y"�*��q�p=P�����#�3F������9NLs��g��sZ�����K6{���yd� ��}Pޔʇ�Y�}�[3t��r��W}[���K�+At,JZ�D�$δ˩F�y�3����^|�:	�2��TV��/#����W�y�������1�RЇ=��t#e�`iB��l2���jhSGu�<�і���Ŭy���J�6�=!��+����R4M`�E��/�&�ś��)g��1$y9,On�����ΐ�_6$�Tc\��F�M�+�n���*���A���6���c�K����y�Зm$�\2S*Uj�°�Q�Eu��cw6��9�;���A;�롷�p!6�j�期�S�����2��Zv���i��_�p�}I.�p���5�[A�'<ʃLL5�3:A1���|)Ҝ�e:�,.J���M��;~S�4�è��rؚ���x�+��g3�7��rm�����7�-��K|^bztnFZ���q�g^[uC�=�P�ѐ5'/����oد��_��0["+���Un�����M���-��=��û�(��BڦhSQdHɴ��y��/��y�%���!�ؚ폔�!pMH&$x��7t�a��x4��Y�6�G�3#�G8��k���w�p]�w�Γ�&#O�/=n&���Ut<��yX}.?ق��j3_��5�Ȣ����ElTvɖ��jJKo#�"E!�8GW��j�7C���������c���r�`� �{K�F�:TF�P��������/�u3��ǯmVG$:C��2�.���m��W��F����#�����dZ�B����N5�F���X�h�R�n�3m�a���+��{���6�|�����/���Ap��(lZq<���f������[i�x\&����>�����c�C��l�w#��g!4Q&����OTμ���f�"�q�Q�q��>�z��W�(F��++H*r���؁��6������d�#�-?�pfl�,NÌ#�9ޛ-;�A���x�^�&Zǟ�Ж7�e�t'�W�%�y��2o�|���@!P���c;��V\A�x T��x	}�4��N19Nx/]=Q@OF,�&�5�Cd��邦�I�%����c��~�g� �MD��]���Q�Yl�>l.fe75wP�$㵣u~h)�ȫ�E>���.��v�ڏ1����a�՚+��@�o)�<q!��L�Л��K8 �~��Շ��.[�������h���bg�sьU����􇬉9r:-c
��z�ع+��hAN�����r2��L��a_^��(aDW��DA���*gq�1Y?* �T���bD�=�8e�~�c\T���[S�?���4�/��=�ZE]���@m��WL�ħ�#"�/��?y�c#Q�yw�tk�]�|�5`�)���>�Ҙ�)+M�"Wӵ̥<�w8�=D*^��1�bTx��BW���7�;f�ͷ�̑"�y�|���� -e��ڧwJ᢯j�-�eGڐ^-�\|�Ӑ[���%(���;q
�d�q��;�$A���.T�����++}s)�$#2���ѹ��n�`�G_�%{��[Nmu(
��Q�xL�X�(�ٹ�=���خQ�~Rc�>�eK����O���&���9\h�*�F㇇J-A�F=�BW,�J��u@B#���i{��������;uo��`G��L��%w�h0Q8hQUTK�"Ws��X�P����6�'��q��4��җ���Z,���!$��~��衇%	��Z�f��.���)�˸aj�0$u������Z�}�^�Ie	e�Q�Y�d��J4�/�P��5#���D�Lb�����Ig���z�b�t���i/����h��b�P��4X������h����<r��rv��b�;���3
� M�P��G��GO��3e�sQ^����3�9�	N G��_p�l�rw����S�D����p�z���e׫L8|�_�����7�Ѹ兊��`���-'o�ƤH�	�6�J���;�v�F�Ԕ�uZ5 3.�M��=9)gK~Em�e�K:-��O�nU:Kb�!A�v��H��x\�fv�9�{H�7o9����XT�X!&�y摰�Z{�sZ�N�5֛#4��7���5���"���`T�i���E�0��&d�=�
������� $�m�!����Z���Y��ϙۭ���7CB]X&ɶ����N�n����h�x>W�1���ӫ�Z������������#%����H}��z7���pE�5oR�iL �b��J�@���ǆ2%v�3���Ɇ��
��w��^�� �2_�j����$�S�	s��f#xl�`���7�{)����r�7��79���#p[���zN /����us�Vﳂ02,��̟>�j�9��D�j0Q���5;���د޶�稁����'j^��U/8A��X	)�������\���_�%��;��XBP��CS~K"g��������5�Wײ=�z?yP��ѓ�#�DU�d���l'����Mv<S�C��K�/��Ŭz��x���i�
�[�"H��i�ؕ���lwc��(_*L��.��c�9�r��ޜpX}������Q��5�D3�#�k�>�-�8�D��]M��@�@��	 7ۃ�y4r�w�<�|���\d�e����3��)'h�҂���e.&�
�Pљ��SW䴸#k�r�O�3H�vAԖ��u�Q�_�G;��V�%ER�k�{�fݖr��
���GѴr�)hTE����8S�g�e�X�ˈ��s�|j1a�����j2�z&�J�����lp�Msv�p��}+񒂺g��Y�LkM08�2/}�-3�]?���A�6|���'�� �� ���JEEߕ*��9*|+@s�htq �+�i��H�i�|��n3��f��o-��gD�j(7&�W�ih����h���oC�w�!N�߬�%����p5�*@Ǝ���NЎ�}1�"�`RQw�2@��X#��GJ�Be�&�E�����C����l��o,< ��x� x��o*Y6��q�Ï�Ab��@�|�ͩ@���%{����h��_���v̲��
������h�7�0�(t�X��,��U!p�Vn� $�I���{�m.�bô���}}=c	�nLA
Oe��2����L��]��S��������ڬ�X�%Ni��ݵ��I�E����r8��!Z`2.9�<��1�p�y��ղEDdE�_��P[�!���������}A���y�B/���a`CS�3&�'b�	���ݫ�K�W�������`�fg�r�I��#���Z�Y�F�Z�9� �W[�>;o�dK�l4�7N�s�Nn� җU�9]K�-X 1�L�y�>��Dp����;"���������Gߖ�����J_���Ӳ���CڴJe�G�5'P�(�W�Cd�����5ْ��ݍ��c!%�X����3�id֢�L��L�G+:Zq��aT\<�o�BnP;<
�@���P"������hz\#�g��!c�����CRA�rRM����
SB���7^T�$���8���E�M�2��	C='�HYb7 uj ��`��8I�&!�R�4e��اV�J��Zk�0�Ң��a�R�<��GO�umHg�8��'����F ���)b�^�ծr�v%CsefV��yxg�MI~�!�C�X��*����[�����]�����g$�xQe�)׽A����&��ɷK幑-���-!���t��HV�[���x=�2v�M���BdDU�o�01CΛ_�����|�或���?����͓z�Qg�����`��+$�)�����B#xX�"0�k��.�*���d5�#��4��D��1���(��d����(pM`T#k�2w��U�p2e7��"@{��+=�&�W���ܙsIU4��l�ډ̨c�/�@?��\&5My���J��-�$��ng��^ί�v�N:�XA���{İ�7l�V�m�q;;�G�����7`��B�_=͛�ȻHsM�j �5)Qd�p��[1)|u�a�[����z���cĭ�%��n,.S]]�c�|���_��ϧ�%��"����իG̵�p�8���b̨��I����-fs��[��R{��VU���%l�bz��
�P�(nՓ��w�@3Lk��	xu�k�&m_>�}S��*P)����g��R��ꮴa�C]�h�ߒ�Q����Vl�÷|���� �t������>
�6�h	l�Y�!�8'I��8��g�+����i%��#��d�rJ���J{H��9�Г������ Cn��u�sY�Pq�.T>�Θot�\�����3 �0���S����`�ǝ�c��j+�] W��M-������S�� `(��� ���.b~�+���23�_�e[����ūgt�Ɋ����{F�&ω^�@�=L݄�VV"1eѷ�$P��qy�����eߺ���	Uqɫ�d,�ri���h�8X�GR\�9�L),
�:�x
��i襼#]�w��Wt;�j[&���e�X�m�"<�sY����6τT���rJ��K�[�`GW�
}���� ty&#�}a�m~������@u�#b�xn�t@W�CT��ߙ��%�\�~���E��04~gw���	{��奇�t����=_M*b�Ӱ�OG�y��@�r��t�4�܇K� ��/;��E�@ "F�#�M��O�����r�6����~�17:��9��8�.�����n��
�y���^��m�(�$r ���Ew)�s�"��l�4¹
;���M\t��P���;5]$̩�������t�m�~�兼�E�߀�QViIJ�X/�d�d�0�a���ҽ�l�a�0u�_3��Hg���*��L�3C��s��k�$B�v*�D���;-2�� #�U�iw�w���=����IT��}C����8�$dw��`�f��[ج��Π��Hеr0�"����ͺC�<9F�M'x=��es�݁OH���X��im�q�tywk��\����á��\X���?ᏸJ�~��9G�ks����*O�M|.y�I-���݇~���"�Z&�t>��/͗��yb��X�$��c�D�֍�Z�|ޓ���w7��t	X�;&*��s��˖���n�/���\.Z	���ˮ����P��ky�5!M.��c���)^���l��%�p=/Y�u����8`��Չ(��?������]wVb����or	��V�с���ot����(n�.c'Ip�og���٧�-�R�	��ִx�����y$q��K��j�y���H�I:��g	���Y�a��}h��枑%�l\ω��|d󙿀`6���w7b�5�$H&L�9b�����7s;<4�)�~u#h��(��1���'��8$��6�$��1�]�t/���mٚ�c���9�&�z���l0���i���D�T_���>�z<^�Z!�;�y��C���������F�uvGQ�0or����Ks�;��ؠe�^~�v�F���x����f@�|�hX�B���ċ���
��W�q�U�I�y�H�s��ԯ�V�CtǮ����8"���h:5!��,�����#¦�D�жf�k���O���q�:�D���e��(�����
 �=Hx������;�f��:l�)|�������<���{�R^)��bHq�	�^�LYkm���}z�T��lP*T�㯬�L ��CR�"��=��9B��#�f�BE�X�T��1�P��������]��<Z�pe�dVC�����\X�IrnpC�	ݝ<~��Vˏ�ءb��C�ZH��J&���ap�K�gc�46n#���RH	�0$�dI�lU�u��DU͠ZL��[�~�����jBDn�~����b�;;�=G���~��>�0�O�5�y
�6z�k�`E�D�/���ә	|^M��5��z~�]�H
A��M�T��+G������ð������k�gN�q�����%��4Ex�fWC���;�=�����u�b�@	��8G���dV����i�4]�F����V�����ՠ��n�VP���� ��^Eԫ5��D;j6��1������^Xnc���G���aq���To'�+`��ڱm���k��N�;��zk�<���X��"��&u�^�������*6F�~�g�6}<�`�\
&�w6�#������5x����/���M�p+1�Xq�d����`-���� �0b
F�%�Ľ���r���U$���M�Dsn�"��\��u�/k��y�tĸЏ�) �h<Fc0aZj(*1�����Kj§l2�/��K�=jo���U$\��F��6��P$�U=�,]�@���A�*��Łd���H����5�+x�e��$Èl��P�Љ�K�M�(2�r��<S�L�#]�(Yń�;��G��Q�N���
j�%�v��n�/.c���<��[�z�����4{S���q[��*q��*,5�澗�80�����O�x��b}*�����Ck�x;	#��kWbD�jԇ�%���X��n�Uj�n������|�}`Ay�i�e��|�����2�7&��P�����x����#����_�t���z�Zx#��ʏ8p���	&<��@�%H�-wdL`�.�^�(._���</�
���sޗ�_k!cE�Uv���ꃑ�t�F;0���E���@5�&6�k{��*wᚕ�����c��)3�0B��p��C˵J����#��5X38�؎�k�_/ �*?w�aC�� Kh�i�G�b@��Y>�ug]��˸s��Q�n}n��*�4�q���$3����'�05����>r�>��~�̈�����9��x�A\���@��⚁�����픲�7�M�h,�(���8�\��s�qk�u������tF�p�N7fuߛ���+#(� o�h��R5�mBz[t�R6󠐥%O��`���H4�7	���Q4��T�Y^�O'P�M�^�:~@���9�U��5�~�wkgcjV�.� �DQ'3h�ѽ�8{�pm
7KO�$Љ�y�X_��h�*�P؝�('�ULՐu`�sM~y=�s��d�� ��FX������t՝~�p�_,��՞�62�U2�� �R���UL$���Z���+p-��b�w��fOoX�����Gb$�I���~Y�ʜi<��]AgTtz=ɬ���?%��SW3 �jJ��a}�K�NQ�t���D7��a��9~�Z!�,K�R�|(6o�8�$y�=HB;�ߒ�3�<k�����p�x)��Ep�2��u)�	��I�CC�P� �8����0�����?cQm�$����pU�74�rZ��QmC�c$NM;�t�oލ�z�p��9�[�J�(ۺ����S߇�{�F��qo���x�x�Áˈ�ľف�6C;��K�I��Y���X��U�=�d{�3�q�(;�?��k�R
2Q^d�ĘLwS���8 qz%�ʖQ�Q*�B���akH�9����Ns�lNhփ����6sJ��ל������}�`�������<�d�6.�Mch�~�Ժ��K�W�t~z-��ț�+��_r:T_a�v/�*7��z�g�Ul�ݢ��^cf�mO���q����Rx���t� L=�]�1%����( ��������[��c�d�6ݘX�>{>�Omt]�6j��!}�"<�[�)Ү^{�	�q��;`��jn�ѣ��������g{a��d)A�K�Q?��%ȱ�3f���!-��M���"�����Z��1,i�z���ʌ)�W�x�#�e��������%��Ă���BE
��	vt�qp�X!%�ϻ�N-a�L�IRlOv����E漧d6&L�%�`%��hx�ˬG��|t%���l�82�½Le�M��:�$�� �\6��}��fKv��2�,ʭ�t\��e�wM����K��i���d�C�6bʷ�Rɋ�wA��1߉���;���b�Φ7j�:P�u@u��}����7'�+��M.�\������HP��1���#���uςH�0iϪ�R�Jc��PQ�|�f}(.����������R/R,��;��������M�c'�3ڨ��0DE���A��ISP����73���d{ogҟG��.E��C��N��c�M��F@Q�x���
�=��C J�� � �P
���T'�!�+�E��8g���l�ԇ� РV�J����_��� �2��zֿ���5�K̸Ɉ�C1c<��M�(����rI��A�e���VZP�f.b�)O��,ѷe��D�n�P>�8�F>U��4)��1o��T�hY�i��+S�F��M�@���H������'R�]R
FN�T�U������ݾJo�� �VH�������>�ۮ��{]�8)��gL#@� P��b��9��'�^c��B����O�[��Mf�B>��8B^����ViN��r�#��VtY���iڴ6]��SO=B���FR�k�O<@�Wf��A���H�����d���pb����~��*�PP]�bMۆ�G��YEO�����d���	a�wg $�d㤛W�6��_c{w���W�~kt%lo�h7�V�i۶�(�7��L9�=��b����y�0J���[$�c���T ��>=���s���������0]÷l�^�1X�u>�(m�)�������F�*i��E~��Id�jm �{���!���%o��G�S�7���f�W��^�A~'���������u���k�y{�cE;婫��"����Q�H�����6&�(-�]���2�l�٢�^������_ Eʶr8�^��_�����s�:=Y�\MԼsm��U�'��)��O�@s���ǒ,��)糷��r����1�?N�Wt�{��F2(B8��k�yt
�H�f�n'����V���� ���9��>�gz	���!�z���H>��ʹ��@J-�^�|oJ�i��	��W:��I{���ɵ��!�u!�gC2����چ�29�)p%S�9/�SR�	��<X�9w����H8���%�z7��%R:5�������3���%R���v��{�~����M�r�/L�����1�. �/"<!Z�u=1��]������R
�(��G�}��ſ��n#q0�.�[h��t��iK���������ɬ� ��&��6+Ӄ;af��[�6�/ʤG��3���Q麤���n��KDp��,�ݏ �Nӎ~�x<�R�r":��-��/BҺ\�f��{�j"\�2O#K�]jU��K���*��>*�<i���Xx��m}-]q���#���o\��{�5���h�f0B�e�'؄G+Y�7��N���3�,7��d�����7uN�q'*��e��5�3�Z�q�)���9SQxM]3h�WzjZk��#Fvޭm�lgN��.��#�~�k�<���T�S�tz,� 3�|F�k��4+�O�E���i4z�c�G��h]:��7x!�tn&�z{��1r�~��R�WJ�d�IjT-���oǀ'+�i�}�Ԏ�6o�pQ�$�%~�.[���*���¶�ޫ�3���#ꅓX~�Rde�y�%�an�A�6��������=VX��`��j����N��{�f�}d�	�>��wfRZU7�K?�,z��C�iZ�;�>lo�)3�B#֕a)�J�o���ETq;	�O���`VB1�^)�����`-�ènIiW�Л��du�P�b�r?`i(�U�N�P���D��r;4Bma��p��/Pak�v�o'p�%R�,��R��M]������.�p��x`tA�Qe�U��ΰ���L�h����� �ו_��?D��kn��?ҿ-W ;�P1�3��`��#�x-S�Ը��iO!yq��>���O�K���*u��uM��I�T���өF<�j��$)y�2�����	T<{��Ej�[���^�x���D���]�MƅG'�2��P���°�0+;
���Ⱦ�GV
����d5��)-)���xY���jrkř<��3��(~Km'�0	`v^A��[{�NP�U�_4����!�%'$-�~ٌZ'�v����_��~&��4S����#P���E)���]�q?X��M�LD���0E�ntr�h~Ԟ�,E���F$�^��H=��a�I� .���5�w�>��L�����=h�B�mWK6���n�l�u��?ǘ}������J�<��U��ͣ�Q"mD�?v�1�z�
GW���B�y�}�_�F*g��Cc���A��A���$� k�X���ۤ�}B��G&�p5�E���HY���V�:���L��$��β_��i$�ٿ�1��2c��F��V���Z�r=�WY �?gdK��X�ؠ�t����}v3.=�=��ױz�4�8{��f�"�zH�L�xzCs�H4͖2ffNԝ�7ĭ�����^_[Qq�⡯̲N����߻�j���h��3�w�ݤ���y��9�de/yU��}B��K!�����}�-A�7'���/MY��:��c���!3���x�c�ɶ�VOs����������-Ȣ��@�.�h�Z�a2�.�.�X���I�,��_�t��&�2o�ї�[������K	��1t#w����Q�	?]�Nl�VH�e>�iw(�3�;�D9{���=�~�(Hݫ���r|i�����C�2H}G,X��0h���e\"�?�%A�LH�ˏ�!��8ƅ���.�b������o	����M^� u�2|>���>�N�_�&mF���"���Ηp��Up:�ƺD�74�����=9��eaD�
��Y~�-Y�.s'CA\PzX�Y�MwTG�)C��/���������#s*���uFs�#W����,�hM5$��w���M�C��-�~K&�q�.����<����i��9^l縞�LV��̈́^�h��*A^�%�H���g�%D�Gf�2�)����)Ci/H:�p�A��;��4�Ϧ���:8��T"���`aQ~p�n|��\Emr| =Y���Y���SHQ!u��S05�B���L�,᩠9�-��L�|���g�"9�E��>_l+ʔ�A�-�� $���0`�a]�tŻG����hB��d*�B�%4��G�n#�J|�yC@~o"�B>U�8��P~�3��e)�^^#@8�L�i�=RfY[y��\�f��K�i9"7���z�5�t/���@��dTBGn��0�����y��j_�N������	�����f�+��@e"�,���5�8gR�/e͡�R��/13J^���y�qL�$��79k/ u����O�����~�g�g��v�s�8A���tlD��Ԕټ�#%Tf���'v����-t��f�s!�=�;�c�3��˻ۥŁ�t��]���@_����o�o�--<�>���O��
㜄"�3"�����/����¤��w{5��*���m���1�R����%���X��2&>ì��M�2 �y���꒽*A%y��i*���:�Y7�w\���+BeI�Ͻ�0��CW����$8mv8Y�~�Y&����尪$T�s�зV�9"�c�H"�&Y���0�R�<������L2t�Ҝ����1�������C�����fvHu��QZ�;"��%q�F-� �)��gDr���8��,�$,���s���3,�u�LY2��3����c�X�G׼��i�_��[i�y6ɵ�!~�J^�	�e�
�nu��R��@�\;tM��)ң�䤤�����i�'+̢,�:<��j�!*�ȟ��)_rצ�k
��@��?4���yV;�5�P�U|&E�/n�@�g����z!5�9Os��}�������6?�V�
��g�j	X&C���x����+y�f�fyM;�[��x:Ṫ�]����w�`���d��?�=5Qސj���</ g��CD_^*?�s�
���q��2�6�ۣ�3l%�s5Ks�NE���c��0�|�k�
K��Dt��^@Eω;�P�-��v �F�浅I^+�-�^%ϴ���6L�[�ߺ��%n��m�1��ml���c�5�E�|�z�'�PLV�P߼y���?�����f�u���1^kB1ޥ���5\��Z���CE�~:Z�iv<�yC��0(�"i�K�^'@���"s_�6�nR`A�:�Ey�rm͂ceo�">�w� ���N�{�*D�k�tן{gI{��g��'�v�WCD�&��������C�����dH�H�}� ��w8�X��s�]���s8���"��20a����C�U��VY����,6ORw��<�ʻ��4Z��Td����I����s�oI(���C����6A�m0X�_L����p&���^��JD�}_�˿��8Z���>յ������JV��X�g�7��{/���vy����ɍ�5B�]	'w�����7�l�]J	gjEp/�ig�cJ<7}�mj�6�3,N�i�}ǿ�l�h7�h_uP��q`mKّ� -�Ur/U���ɁQc��r~�F��d�?�{���.���QN���a�F�j�_�.��Hs��r�J�(�d!K��x���>O�q�]YY�v��T�K�	��$�UN�_zqz���wa[[�,lv�e9�N;g��a��<@ ����(�����9�8C���,�*��E�RUp�B	�\46�TΑ׵���V�$�/�M���C�T���{��~C:)G�~�+�|�Ӌ�A�,��:�`2��<�E��1���x�H,
�ά�lk�B����v	�y�zP���z"������[�#�s�At�Kc�pA�e5�{@����.?<Q��ڲ�6��k��;R�����e{K�$zUIԊ�f?
i�\��J\z"�9~+�x��&&��s���u����Y��wF48�����]/[�Ni!��O�x":�%=�G߹�'|�i��//��&��\ɺ*&�>;�';jibKk�	���Ԅt�(�S�G��A�2����/귡��à,|���}�L���Z.g��ӽq}�X�S�����#��Q ���	����������j��9g�[�7�Ԡ�27!Hg6Aq�F�[��K=ˌhJ~r����.��/?d���H��Xe���B�AU_\3�Rh�	�+�Mt:�r�_c����鬛��S��l���n�TU�u#����9Bis��ѵA���]�fWXO�eB��PK׏���Um��� �6=R��*ש����[��\�|.3o���t�].�+Z�ft�V�s�d�]�,JZ��Jv���w? l���;r˥-�oF/�zڝ_0��⁧��E�P���-��7WF���B/��Ro�� �����M1��@�ZI���s� ?p���ױ^m�b2$������&z?����2|���'��[�t��eH�n�u�O����+��#x��w�劢ds�^dπc0�y�뺐��5�r�n��o��&��o�	��z�M
U9�v+y��Q{z�	{���o��dL��z�	����3��J����o���ee(T<���j�[��3���>��@z`	8)N�[����_w��|e���_��"������u�3�_�#sYv���e���=2�l`˭�8�h9�f���A��f��B��-���]9Ex4u����YG?�y]?N]n�$9�1r�1���Q�;�T���/8�»>[M�q���i��V�te���J��
:F�ND,��`�GЙ���`h�� &]Bm���0�$N�p!�x��¬�j7��m����q-!M"p2Cz	�^ms����G$M���Ԁ�5�^�^��,s��p;a�:�ڌ;P�6Aס�K~�����5���c��;��5�s=g�x� i��"�U�}R��B���22�\��T|�#.j�<�jK�2�Fp8J�ʌG�J�DX�'�xT�= ��#�:�oV(+W�7���̉�����	- �)�뭕��p
�_fV�W�|�z�X�f��H� 쁇��3�%��p�ڞ����#?�(�$���<�H:���ify0� _�e	S��m�G�6��cQ�7�~j#��5���@`}HX�;��V��X��'t�'�F�����ŢU���ץ�j\yT*R���҆�����ͭ���)�r�E0sT��������_�K��=�d�	����ԟ~�M(���)��$ٛ�����d}2o�҃3�;Q��PmY�\��"7���5sB|�����-P��Hn�	�ĬJh�v�^��l�2��tq�Ԕ ���:�e���6@���a�<c�eIj�����;a�KӲ�KH���Wn]��-"����V)�5����|�`2G0�:���R�'�1&ǣ�Y[~���_ç�Q�\;Q�V��K�@�.Y�WUաr�ğ�$��)u'(0@�s��ר���ť��K�W�|��X���mOS�Z�d戼9$H��o9~9]���M2��J_���C��zu ��ZU|�d�C�z`�2����+0�puz�Οь2L�!q��^4�;:-;Xki� Uxh�z؅@��j�K�@.Gɬ+7O\P})�E��.d[�;r����"� C��`Z�8����%�<��`U�A���q���w���<�|��xT74$G�����TXw�f��42b�p��]����5,jl��1e�V���ۜE�	m�^-�^�q)1d*�"�+1�쐠�(�uv_'J�~~� wa���Y���,�����桦�:S���1��g8�����kb�~�ez��wbm���6�ey0�u����@�Fp������6}|
A��e���ω��$���ؒ�<�K7	���Ʃ�ִ�vؚ�Ǖ�����Y^9OZ
���O�"���9�=NjO�z���r��S�%{��b��΄�?�o|����s�� ����Б(��u2��%jh��%�II��+�0�:{����6o������O7�e��/,�h�FW*������j6�+���'���Sd~#DL���Ujx�,H��ݟaI���!�=}�����_~�\��p[�	�=��N�� +]�)'�Џ#�0�WN0�y��m�Hn-/:R��kĂ�^#o����˰��#og�0$Y�x��2��m�� ��y��'Cϡ�D�����\�-�8ǜ�/�806����{�g\�)y���������n\�M�X�@u#5r=����1J��%��7�Z�b��K�����5,�}[�>�C�]&�w���i�� ���bY���dXH;u�g{�p:�9���-!�7����^)�QM9+k��8�3��`�7v\SK���W�!��FovReU0�X�Qv��3QZ�0����P9`̀e���Փ_�2}��ʐ)���"B�!�a�4�E~�y����p����E<���߾�!�K�1xt���ܒ�B��l'Wu˓��_̓֊*��c�̈́�9����T �e���#V���
�9ȫݦ<���^����3��I�3oeA����<��&�L�q3Pa ��½�n���6����^��C���$��9 �^ۖN���c�6�><��,U����4�
0'����$9is����[�k2Y|��%�!�^�~u��ř���6Dk{�t�Q:�g�/	�G
}�C�o�!��\����&Q�RׁK��At�4-�x��P=6F�{p><��S.+��l�f
��l���d���c�XQx����n��ĳF��4_��}C�{]e ��E��5�x���*�������:T[��,)Y���<	��p���E��HqN'e����V�b�o�GĒ��͸�u��ӂ2�c�����퀠+���0��=�'f��=*P��)��͸���ⷁ�s�fN���Ն���:W����kj�؟F�/� (=7����mˤ`/M���Z��RF䣡�;!�m�L�c��T���4q�t�Ĩ-�_�{��A�;�T���+�\�� 5�g�+��c� �«e3`INn^B0��E|R�n�C���O�&�۸�'�6C������$n����m?���D�����[+����&D"���L��0CZY�n������0��&��*�Ǧ���ω�bb	>��~~rY�������l��Q��)��FP8t{����кa��$��jQQ�xZ%Ok�F�b�ي���]c���A���	6�Q�X�Q&�(.�Y�i��Vc��y7�c�K#��հivc�p��4� �2t�W/\]\�����u����Urc�1�,~�lP�8���%ɁO�OQk��6@��E7µ����F�V,l�ɩ:ڊ��.����-sP�\a��?�$��!��^L�\uZr�����J!(��+����y6����{6b7�-�^���I9���ό��T{;��N��4��7���V����b���Cʣ�B�K�]�����y�˳d���a�MOԎE�m6���rD��a��lzr������h(�-s�'��y����5�}w��F/7�6z�6���3�Л�9�3)�����8��-n�O9nW����\ӌ9o ΟA�:v9�#ra��q���h:��P!��-�!����P[Opi�7���rx�Q
!���p�<�
J4�A�N��(\L���Z���!kgq�Lg����Ձ3I؏,�-n��Nb���xr���g���#�ꉳ/薢l�qHh$��5c�K	����m��߶$ ]ϛ���(�?^��/���E=� ��o���QB��t)�>�쳮����"qѐh��N_}�ݘ�����.)���n/U����M7�dCm�� �Y �|�h�ۢ�M�y��%i�ԟ?�ۓ��Rm�E��J��3���+��֠�L	�J��F�BTwM�Fk��ǙO�!��%�G"���?W�d;`�t��`�1Z�`�˥>��r���C����,b����j"�rؓ�Y�t�����U6z�t�k���\����b�:y�b���ռ^�cʱ�٨�0x?��X�	�A7~����q�es��
>Ѻ�6j%�pF��Iq\��yfӓ��ki�z�g=�xaX���s*�C�Nȶ� C)�m9ъ[Z��b����۝"�ݚ�5�=W��u�:4��#�@Anbe=�S7V��Y�qs�:�����T�I���$��.`�"L�7�����E+3�`��v�_H�_k�,
'���V���<5n&���m�`ר����؊�r5�C�J���t�Z4��Hp1im���=Dޙj;�u�WS"U�:O@'!\,�C׶�
"�yɍ�-�8�Jq%v�<lGt��,�.��dk���3�"x�uL��a�  �f�L�7j�.�.����k˸͸�U�u�q�Vj�k�2'�{�|�����3��X;�\�$�O��v(��D��ڹ�mr����b
O�js��p��N��%��\�B�]�M��Uz�螾K>P0c�9~p �����M�RW]�v�e*�~�v�ѧ7�=	c�٪V6dA�LG�5B*K���;Хı����E$��m{U�8f�i����p��c�q<�=؃Q⤎�����Oe��qYU�]t�<�o�D���&�/�`LX����|�^�,�*��,�[{"mC"j
ԵH��ll)�I�,$-WQD; N���'�X\R�[ᦋ��B$�L<�L�����%S0#�5B \>��M��V�J�ȍ�2��9hA���ٳ�_O�����K"�#u4��栥�G%El�3�� �(�z���0
�î	�P�{w͜���r�ӊ�y���"	�I���,3Ρ%I��l4�(����R�'�R؋�*�`���ɍ���������Gi�9����m�)��#)pJbG�I.��.ᤥ��]����ᑨv�t�e���h��%0�����Y�,J	�G�29�.q�K*��ƶ��d^`�����`�x"Ǚ�S]!����������p�6��~M?�fZ�g�=�C~\�Y:,Α�ǒ���5q}�ً\,D䍜s�*.�,��$3�����Vh��9NPa8`��" ��u�4!���3l���9^$�z�xB��Aq���������m��Ф�ۘ���F��|���6����s��"?sr�]��Y��0Y���-����*��ͤ��8���ք��G@��i�eC�3 {\@���(�3N�[���[���'S��d\�,-e�Y�1�Sܠo���T�E`���
	��َu�j����%޳��q�&C1�M�J2,�ӃRͬ�ء�|<浑QrOJ��A��*���3�<�;1�T	 ݧ]��)�}���!N \i��f׈Z'�DTfw�ɪ����f�+A<el%Gإ�~�V��Mְ<�<,&�e������\���aՓ1W��s����(��Xye��܀�4��9!�GI|�Ҹq}�p6�F��eJKXS�	"Y�Wol�|Q�vT��Nǹ��0����y��^�2�2V����=h�zz�p�Ò���O����.`�l#6)q�h�