��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���C1��
��4��$�6vW��a��9a�#E���}�k��?�|_(W]�?���D���޷��!�h.�:�p@�A�ҹ��mJ���=��jf���Y�\k�
=��of��.�>���ݞ���χh�s��W?׼t��=��ѥ� +}�B�}�M�.3�y�]��2��@�0p�o��H���p7X)���.���t��!s3\.�H��w�U��>�c��CK��^Z���OXW5�!XU,�K���/���;���[��ɗ�t$/���4�#�|��0�P�� ��5�n�E7x���)A���o��/#���?	p$��YOe�	�B�́Խ�0���H(�P0U�����wkT�N�$��(��jU�M)1	����g�*����ݻ�U!1��{�&0�^�|��"��ݠ��Y͝=��`��U��>��ڬ9:�^�X��U��ݲ[:5�j��(����cFk�̪���J�!G��l��PV�X53Ã*7:�v�x�e2���������h��La"�Xș�d*�l�JI]%�� ڦ=�����/���v������+}h
[:�#�q���әW����e����X/ؘo��_2Q����u�ھ�tsl����BR��SH+@S�ۯ�뎋w����}�M�53CZM3v4M�'&������dg���m�p�)�u���:�y��B���?�^���O6SSFӋ6�w3�'Y��DXM����>�c���_�nD6��6.�T��z�����_z6'o��F�o)5�C�TԵ?'�#�������,�-˶��� �ӥ�0�lTފ��i�����;�?�@}5��XT]7���7��f�\���ecer���/�r�!TcӒ)4v�'��h�Pԟ�a�-�W6rئf��PE�OVi2��=�o��fQi�]���n�����h��@��� A̓�gF�j`-��y��in��m�S���T�nh, �>�LP:ŗ_��$�v�x=���,�������3�ԟd��g�	��b��l�-HQp��L�ݍq�#��6��7�=�� ��-o�f�q���eP���d�E2���/�+�a�Y��,R�kx�PҗS�v��jk�ʷ���μ��Y'k�#��I7&����6 ���*u�����x���Zj`�s��(@��DU��%J�7��?��:2he-3���K��m\�/6TT,܌�p���0���zV��ȭ0�{��*��L�ȓ�L��{��')�Ė�$����}��h- �(u����S�gʄa����4�_�\��h�_�?�e�Ȇ-����^w��X�v m���Z���iϻ̙,������Ъ�Y���>,D���q$*�g��'v0_��^�����^���>����"��yB�gX��ø�Z���Ň���[�#��6��#�mq�^�[��J��M O*	�#����2R �i�ֵ%�Ѣ�+�:ȴ��ͺl-u?�m���c͙2/��g��@���m����V[T���H��l<-�`���>�gTd����Й�#�ju����˩�Ɗ~"�5��j��+OZn�R�K+�]aAݳ?����iF�Q�N�c�^��{����/��@�������T���D���ӈ饁�@Z�⹴�����"��*t�O�lp ��Gƿxzf0�5ϸ�F �Mv"��׀��wks)@�Op<�(A�x{�x�������b�qNE��9�M�8}��:B�DSn3v������-�w��Wy"6H�V��h.���2�(��|r����vzS*n�(�,� x����۟c�O�~��vKt*:T��Z�s���ˀ�XF^���N�������\y���8F��*����=ө	%t�z]0��p��sD��&�x���:$�1g�/IHb+�{}�V(G�����{ǯ\0(���ڲ��E{f��,C5�Q������̌�\E��Y�n��]��*���Z	eފ�ޢ�\�VW�>�%��NE�:��߱�
s	�e}��E��a"�D�d�n�oJ�����4nJ��7�i`п��΀
�� �1�{��djw�%�*%Ʃ����"�˪���f�˺��Nl� �u��m��KxK�h�����H@��%�yk5^r��~��۞���~=g-B���\�Z�m͝w���W��?�e��zg�Z�En���9�!�����c�)p�Ul������3kU�۰8q�p)�и��f�h~�hX� ;������0��m�M���k���:����O���O3��-^6Ӑ�V�V7О�!� �X����,Ӈ�� ���Ҕ����2� ���<\Z��6s2��l~\���*�����|���(K��ɶ�Y|K:�-GZWn��UR,��ǣN�7e5+�`��J�쀺��#��lt�6���O���Ϣ� E��&�F��̹1�����.�����y�]�r@��4��n�@��4��VC���J�]ZQ㚔��!��Y$��L�X`^��;53w��#}�ח�}�}{X�߸_�ccZ�䪎��,nvo�ϓ�R�zi2���tͱv��`����<D��}����{����j�BbFiw�I�z@cm�RL?�=��h.;7+b|��K	�� ���;��-�����;y��܂�o���\$�6FZ[uO�J�_B5��7�����Z��.��B��M�����aia�f�t���v'9��u��U�m�������pl swSs�;�&~��h�B��>_��������CkN6�D_ٺ���.�=C���0�G�@�l�u����UO��Ŵ�4@'�qO2ԇ����f_�����ZH�&�~E �`�A�w��A�7�󼊸R�����X��X�!�WNK{?P��Йʠ^H�!Ҳ|9����7/([���Z�X�~ԏ�`���ޫ�{Ӝ��FԀ�*�3
�B�׮��Yw�)����؁����� m����!�O 3��Ǌ{����+*ͪ�'�����k@`;@����4��x����-�\�����>�R�R7��:�WC��xr�]4��Qĉl�x��d2��0��$s(�+�HN�9����"���QO�V����n�Z� YaQ^��2H1w3��g=-�f���ٹjl?�p>��JcJ�t��y���A�=[v�~]"�O����Њ ����	Y�Ѷ�L�%I����T��8VF#�j)9ӥ�%[�'�~�	w��	������_���f�X�1<o�~u�K�O[��:��0B��w=G;>cv8��Ն����l�<�+[$�0\�A��g4���;����W�t���i:�>���|Y?�W"$Y��L��O�:��~�Ji���LnI�U7!,J���BTq��bkL������I��T��9Ѹ(�������l��1��e�O�FD�1 �D{S�f��6B{b��C>M\y���E�[\��(@Qk��T�����/S�0�p�C��Ȃ!�z��V�u�JF株��b��d�{�O�h�	���R@C����qŎ\���9�۞r��Iy_t�I��܈A<\}���������:��a��%�J�l\����{���r���'�`7yZ-��.��QY'��"N��*E�&k����@����q��J�pW���S�����`X�����,�S��s+M���v�h4�`�2_���H\5�L:���$�i�κ�pn�$Ρ�� �v:�V[�z�<�M��
&x���Z�V�zi���oa^��`.���^��j��E@�{X#���lW~��0o�l��'���P)�,}�Z�ݎ�f���O٥��ae�$@�/YtRhݱ�庡�1��K6��P�wia7���+ǦpOIgo�������zsy�i�~����?/��e�� I��K�2~�$�s�}���X��u�:�"�fw@�DYi�=nB���,��\op	z�65-)@�ӝ�D�/�f����:��ϊ)�;��4�U���?��t�0��{\M���";e*D	h\�\��;:f�4$<��F�����s�Kw�,Q�Fo��~�'�2����Ln[�a�}v*��FZ����
�L�'���K����aKircK�O������p��50|�|�ׅ��2Q�c�<j�]��R&s�1��a��9tSI�U41�W��,M����2B#��p�w�����c�}���t������k�@��%ZW�ֲ�
47[����D"U��R��ce��w�]O��x;U"����	�=E�N�zE?�%'����QW�bTD�>�����Ru;�V_�P=m&/\��i�l�@3?�T)v2��t2��\�����
��	���I����"e˶n%8l��s��>8A��HdP��	���� �n�cG!����ͯ����y��ns����i��S%U���O����%��N�&���9��;8~�ꟴv��ߕ�ȼ��h�(ז77�g�▿�LS�q)�f\�'���mU `���!jai�z����1-��0G-!�c�:>%�А
=?�[���ƶ�=�^kė[<���fkK&>��Ϟ�q,�ͳ�I�N,���u��%"碄Q�~,َ������o-�7Lv˒T_�k���D��LR������}�)pC��"���]ԣj��2K�o��(�̿4��ɰ��
����{���{���b�b]������)T�'�6A\��-���W��<�u:	אۋ���1SEv�S|� �򺘞AՂy��Dݪ��L[}|���E���ϑ=�t���C,kVhu�����9^���"~1�i d啋��!���b��%�˚�0�=Z<������ڦ�`�m�Sq~ B#���AO[��i�ۚ3ٽ�!m-F6�ɐ�sj�SZ���Su���Ky�12Wq�H�4�B"}�a7�3�ʂ��y�~b���Q@�:,�Ɠ
!�Hc$�pޮ��;��8��cAq�OkpYV�\c�r��/�@�v�?8rK7N�L�~?��h��h�y ��i_gWQ��Q�y������c��ѩ�%ɇK!PY�z���u�5�<xG�!^�j��g����u���
��-���y���i$�/�eg��+s��T��;K��=�^X�W�@�3;�gXr�[;���x ������4�ɺ�|1�槓v�N	��>�xr�f�:\�1�Y��q�N���i`'܍����2���q��|f�����'=��̐�����p�h1����׈+�Q����p�q_'#9S��B}�J�R�e���K,I�ɻฆ��=��(�%	�H�0m���_h������m�����4�/��̳��U���!���v�0��k{j(w�
�9y6�0ᷚ�[���տ����?�կD9'ɏ��S[M^c����ST�O(~�='V$�����]=��V�pm���"�JC�I���k�cH������w���-��� �z4�0"kzh�?E��łe�� �+Z�,(F���I8����f�ѷʛM�Mqw��/q�G��w��Z��k9��|y� ��]P!0��8�=I�
Ȼ��  H3!�(���ss�c�;y嗘¥��3�I�VQp`�z:����=���')�#~[������-aiI�����Ԗ{�v�3���F5���LR�u���K����_��o
��v�Kg�W���j!� -Yx�mQ�ʍ�6�P����[�^^\2.�|3L �$vs��[��� X-%����Ǘ��G�M)&Y�; �ϩC���.��W�$S�G�J��y�3����ږ
����N@�v��n��?�Q͢|���B��S�-r�F�2�_^�j0}� ��{	A%0}��ߎM���p�B�-��Ya�_�^H����)\�P5�ކA�r�9q����}���lt�Ol�u����M� 9��^�/{�7]�яW췢�)�b[��*�<�<�T8�9�|�Ӑ0H	OWH����d�p�>ݲ�\4 ?1��g��>���~���>����R�bW�7�a�����
U{D/�ڤ>	P�(�*�^�q8�*���iǼ"G��2���y���#���û#���h%��]}���ǧd���f�2R��E���o��E�4�����F����Pĭ�$8�s(�;�j��/*B��MT�ߦDs�،��ȴi&;FZ�ʽ^�Zd�F�#Z�*�kݵA�&����MϪ� �R�챑��ç����<���o�J��7�����𳅴�{^����e�R�o�n��=/�3��hFd L�1s��Pc�����ɦ��{s������!;�Fۤ2�W
~$/����3��G�a���E%3�����"��DX�8�*�i��
}+�VR��s m
TPN̓~s7�wr|�n��/���	^B;Ks9���1 9��S�)Z��-aj��T�,~\a~�����TϘ�����_��b2��ȍ�솙�n��$q������pug* ��5�v��9������;�_�W�r���@ ����C�Z��8��w��.d�dj
��gzW��ݾvo��e8J͠�be��p5�e�|J�k��z�i�J y��DpS_�]�jfR��"`�]{8WQ<L����4����'�8W�"'�k�I&ymn���������wۗ�q��X���L�w?e�lz���Fi~���a���g_ĵz"�נ�;'��"���,��j�N�H��;��Ny�6X�<x�8�tG�_[� �E_Ah��:n"���IsDg|��6%8�v5����[�i�A�V���fx�AV�9C��R�3�h�o���̓�x;VI���X�ԅ�)z@�а�.Mܘn�%�s`S5�6�At�7.�@��d��U��Z����b%�{lI�S�b�%}H47'f��M$4&�R y�JĠ�s:Cl�j QG�i�ة���-��6����d?�����?�D5���-��.H�d��
H����%��.o ���*.6w���-k���:���I��6���.�U�W&O�#�E����s�>�h��Լ���Q�c���jò��"��7Ul(sB&��ߢߋ���`L-`xύL���E�.-�����~k�+���Q�G��>y	@��Uw'���n�ʭ�:�L8�Ц�JӔ���k3�08{��6T� �,�N)�f��������P�K�b��BT�=:�$��r ���CL��éӖ��y������͚�K}�?�H9Rc6����ԝ&���U� ��cm�����DX~a��?G8�`���%Qv�ʯ�T�BÎ�\}�\0��7���[ek7G"@����~^��U��g��g^���g3�!��t��/����������	P��;���TA��y�SP�?1KQ��I^��-��ɺ��}�ȵ�gG1����"�9f�`1u�(�(#�;%.�����qR���F׏!:&�N�<Gat:NX�O��6j��\�U������o ¹7��.��n-݁���n��0��Az��-�_�9=?k�ۋ��n��H���T:)�$�o~���.
tO�{^���@�QJZ���3Wu=�n���=$��M�`��w��}�'�fw\P\h�j������|?}��U@�"L�X��;ìE8w<���uB�
ê`h�_� ww><6�
�ӿ��ŉ�6{ēO�JY�a	�^q��~E�Z��R�7���� �\�����]�H����������K�!�l������X�S���.���$��}i���#�Hu��r�ڡ�:�@�.���G�^�����r��� ڟ��Gr�?cWu��$����ū��<���q���Ύ�H��ˡ��fyP�˛����o����r�qI�n��^�6��V�]d:��`�t�I���U����Ó�aBuP���az��	z���e� ȚP����H��*T�����0��`��\����eY�U[z 泄z�l�IP�S���Ӿ�ތ���;���"��Zy��^[��ZdSv�R]g�\ۻ1�Ɗ�0����QO�4�9�v�^q��ZOO�`�Y�&�+'O��O-�w�3[AW�;��K���A�e�=+-�Y� 0ȦB�ڥ]]髪�.�,����[���rY���؛��N��H\��7����l��t�°�L} ��&�]�J5�t�����x�oS!H��W2Q���]	eVs�+��^Tmmn^��Ң�	H�E��e���j�����C]����Y� ��~m��������+(���+�ԑ��J���ٶ�Q)ޗ�Cs�R��6�f�RW�n!�r�K�.Xh�zr5S;�l'�^Q���f����F	$�͗��sփ�tK�C����:����7��Dp�d�Ȣ�H��Ma;��Q�nU�b�<�3j�D�=\��4T́�M�CW�i�t�Մjt4��74w>!�""��Q�g��?>�u�˸%2!�H2�~i�Ԗ,Ї�\!��-���\u'?�i&�9�qۦ��vϮ����q�n=��2ʺ�����n��m_]@����L�7G�7L�. ���H��%�jL7q�MЁ���W-Ed���jN����-�RRM���Ut��������[8Ťw���@�����$�E�㈈��=/�Ծ�D�^}��8n�6���8@������%'�w�h���m'�$��L-�/[1�Ɋ؁������956�G��=;�4wl�����2����۫@$>��7�TT�T���6�Ɗ��(*����'l	i����em
ҹ��m������Soȱ����i.�	�� �[�􀷙����'sk���-����k��!p��9N�")mf�7��k���O�3$|�ſ q���.
��v�1�|�*8�X!�B�#G"�_�\	�\�T��ͼ��������Ѡ�KG�k�D�*ÑЬ�L�q�i��u2������N$F'�N��p�$�؜� ��0'R�Zܾ�@��b ��vԱ�գv( #���Ar5�07�UI��J�Ze�F�2,'5�{I?����LD�&+⽆�y�2�,�㭅��R�_p��$���߀�=��v�֨���\��a5�4[	´��fx.].ek�N���R]K35��T����%�r���L��b+27�-�r��7��{�N7i�-̶xŞ��U�-MXK���)����s�#Cb�*���z�3�-�����~x��1��D���ŶM?�<?hN&_}l�>�[�?i�#a�iU2>d6�����M��1Vi�d���NT2k���_A_��ƧE/��	����a�>d�k1����	3#8ãȋo�ЗaI�z �6)�9M�xѱ�8�s\��Z��3��K�!�7-wMtB)�A���<jF����1��;Ç�AnJ�]�;B�Z�N��1�)��e.}D�3VZ���x�S���DeFkz�W���������Wn���:<e�;1��@�	}m�)>vfk~�B��0l��E�z4 ���M�U޳g��s����M ��2u�2��F���7^_U�-��~��4f�Q���e'U��<}��@�	.;ل�����m"p�~��[���	);U�NC3E/�[�IɑN	�X:��A�#�0Ih))ȃ��`)��	�OuQ�Ñ�`�K��A�]S��7s��1�Yu�A�X��_:�޴OH~��_�Ý�(��Mҡ�d�{�Ͳ�$�%1ޑ��w�(s��>�!0M�+T9eE��u�Ȧ�ωYCܯ6�m�_�te-٭�(	"�ڍW�*��u{P4���0Pu��5��%�+F����!���*l��(�b��GM�ZH�^�G��@�y0@�%"�(�6�a��]�/�.�R�ۿ��I���n,���(9plt<�'Θ3��qص�~��X�Yͷ<uk�X��0֫U��];R��0#�����WIZ��b�)�5|�ݩ���QI�.�` ��mll���cN7��O��ӟ���]`�����N�Hm�Z���ڥm�m\��=�@)���Xi�Yd�b	�ķ�\���oJр�>D�gY{oWv`��w'<G�U{�jf˦��/��H
�е����+������i[�j���Y�5s��#P��'M��(��.�T���x4gb=%I@b8X-�QF��P�!2����I$���S+��_w���d(e�|R��*���ʫ�}�pͺ���m�1�}H�n�/Y���D��B4gG_�#�B��1s�J9T��O�&]��Ut�Ay�Ӗ)�
WU���*�N8D^��4w͠���kſ.B����T%?C���j��� �|�,�Z9����=�9��2)�U��+^n.~ߖ�5�3�ϙ�K#*x�l���;�0H麍��ϙ'�͍.f�־较�wF�cjƥ�v
�NW }�q���>�����id��J�u���`�4T7�؅���#֯w>v���d;:��9�"�J�J1����Pb��F͟f/��a��_�ҽaآ:�W�[�n9V����X�}�Z:=!h"�]�v _I"������'��y�K�%74tgc_�}��,_W�K��m\�h'rL����R��c�,�Ji���@"�צ[��Z�k�2,�'� �]=̪��7��7tv�~_7+��C2��e�C}���utО��S
9��? ����X��
nh��p���	z�^��}^�cf�k��~��g�"����wI�5[`aW�}:����Î4Ḕ�]�w���I_�F�I��N-|�]��[D��	�k����r�{���/T�@-��<���~�I���a��%��#�����M�F�ِD�,pV����2��򂻹m YLV�������)m���?@V�H��	�~� A꽊���$R�{�W�׏AVx��t��!k>����ᤥ�!�%��C°�����|�MP܏�;�k���������G�f�w�s�W8dX�ܼ�^QBr�ػ����_2�Uƥ�g\-��c��Q6�y�˪$0��m�3������x{R��ۨl���=Cu�9"�Y)@*ؙn�A'��%P�m$ʉ���R��������t�9�,�y��D�n3���y�8J��a��>�!�"���%D؍�r�w��܃�l�繼�~]�:#@����"�կR�p�e9�k;x��77%�!�B ��GD�L&=:y����-�}ހ_��QYL*���[�㨱w�,�%4�@���V����zob�xpKWN�n9�5��#�C4�9�<E�+p� ��DIT��C!\�5�f}��S�W�tkyJ������?Ω�@��Y��9�]KJ�p���o�*�v˒u7]|��<A��y2������N�2�eo��]�I�X��T���-" ��+?��Ժ�tl�r�=�2[�ր��Z=��n�
������zM0�x��)��O��=��4�a�7l0V���e��枾����QWJ9zdy�=����
2G��q>�@݁3�	��;U˷�E���vxt��
�
j�� �7$3�/%�Qu'ߔ	����?C%�j����uZ;�L�R�D��X@\���S���63k�c�M��m*i2ͦ>%�֟�Z�~��\��t���&9Q,� ���V�l���\c(��@�I���fn��u�TD�Gy�R��x������sy(r�9K��~�����R�$w`����ˍY����
���if�e���$<BL?EO�3P:Cb�Ξk�P0�CY2�?P4�*���N)%{]jȃ|@��3-(C�s������g�Ś�לr?�BDj��=�*H������� JGx����]?��9�;��%_�h'�*��Y+/���o��)=bҙ�5� ��Μ���#����G�� �aͦe�^b�@bD�=�H��O�D��g�Ǵ�Y�M���z4�{˺8����`1^ɰ��l�|��֢L��� �������W�������NHo�����U^��\-�x$�yWv�/=��_%fD�5>	 �F?�k�hq���	�v-H,������!/��������F���@pj��g{tZ'�̑N3����SO��K���Ե;�s�$EK�*u�V�7:Cĉ}6~ήu�� ۰6{~.J���%�=At4����U�ԍz ��=Ļ��2#H�PI \K��b��Χe��@벰���fvb1~����#_�a�)�j�3�77(�L�H�2��	o��t���^&>�%xcp.�����ր3X)3�!��<N�,�R���A�&O�Y�����2g�d����p��켣X��A���*�.�N8�uY�Z�fO�TUJ������à���
%&K�� �t��<�,��7�6G N!���I�広¹g@f����^]r��� �;7�h�� Ӄp�C@��W�0���Nf5v.ʝ�H�G�����|���%��Gt�)����V7Jn�h>���0��48SCD�'�Ä�!>[��|u����_�e)�"�$&����򰴉XC[C'Eu��Xd]�r���/Ң�Ø��V��I�8�8�������B�1Wl�\� )}������B�<Ԇȫ�Ey"�?��tl�ER;�v.�Hcm�����L6�JW�U����-�9�tL�
�� 	މ�J��`gc��R�쇝��h�ӣ���.�#��/U�/�_�m�酴�� �.��s�ZU�"��X���:��)$�Q��z[)�ؾ;�X=�c��sJ,�A��~�C-R�,+-<5ۈ5��+2&��av��~ �q�� ���A/����A�q�Ճ%B�M��e-�f���ޫ�\M��!�Ӧ�j����O���t����V�`��XS�&ԕ�iݶ�x	��Cv�N�/���<nQV�����B3�X�+�8�!-�ː�|{gB�sQ��B� ^<�b��Ն��J�"f�wy���7��C)��ruc�G��TA#�)S���4yr8jmv� �G�G䰈�E�ïq��XH�Kס��P���Z΂O)�d�`ðQr���v��&�	B�`ؐ��n���m(I[��lo'ݢ�6�K�ll������1*%��T���6�Xo��FH7�4�褸�km+� ֔���x��&;�6��PJ�������M	�z-��RI����C+W �9^!wf�lsQB���H�;�<%��4�N%��L}=�8}-=��xX��T����1f9��?��F��?�l<c�I��`W���8��?�?x�)�u(j����UrN?�D�I* �;9d�wi��Hؤ��7&�vfj��f�U4�.`����xǷ��u�Es  `"�ŉ���`��H���ܽ �.�F������JZ7��y:'�],o�*Fޣ��#������S�~�ׁPѷ�oMh���s���:1��C����B�E:0�Z�8引�t���o1q�KN�A�S���>+h�E���SP&⹼we����6f��*:��曲i��|l�}��f�,ZXOs��㽓wț���]s)]�5�pU�r��ٸ�M*�ڿ}�bpD���I��R!����o�tP���J�:kt~>��w!.d� *�"`�þ�ɀ2T1䦒�}_�,�G����q�?����X7�}l�������O��K"�TrD����
�.�.�a��]k�����ޠ��>���~����Lbp��	�(��6>�5�u���@�Al���B�bH�rf�&A�(1����=e<])e�_o	�hK����;Uyh�
���H��C��s�s��!�9�\^�"����b��F�(���n�V�m�����W͚�hI�Kֹ�yM���3Ү�A�@��1�����a���t�����4��A�tT�ї߁=�G�S�>Tv������9+���/b�sW�YkP	c�RX"�bۀRB��%���=���P�|H�<�K� �;z >ңt������kPi�������	�.U�R�M��޹@l���Z��cְw4��.���Y�@V�t6��OQ5�a���c0�YqV#� �N+ϔ8��A��e���z&��2����2�Ϥ�&xl|B����kpc��:A=�V��M!CX����F_x�O�w����f^�EPf�2F����A(?~ec]TD�1.}�Qō�mS�MK�̥��� ]�M$\�hΟ�@Ь"��A~@�p��ts��{�D4�h�ʆ=f~�e�MBk�b��Q�HK�C`K�1%�K���Z�~�>��E���?�9�4+¶�l+�F��8���Z?�>D?�۰C:S|z�8���gu�E���'oem�m-�@�?�5��$?��YI���LL�̄G��6$��V-�=�j��M�����'�_��i��@�g+��ܼ5Rp��MA����۶3�CIO�\w��5�ֵ����Y(��Q���+���Y'�B�,N�QJ.L��ZO�Duc0��?�w�9�VD��E�xة/�ۭ��QP�<����q�ʦ���H�慂3�UO(
��Y���+���:e �`�ʴ����<������k��Aq*m��Մ�V8\9彠g 3�VP��~�CiSy�pW����Y���T��M��=X��N�d��:=SM��D��uR1�<�o�i��*j���
]�6�6t�U��_��(��)
�x9k�z�4fϱN�����Q��ٯ�'�8�����}%\֯�����#K��76���9/�l��2~�$�_��1(h�7M@k2�%���z;��V�t��@}���z�p�^	��J=�¹���&n��	�*�:4�9U��gh۱�y��L��?3�!`֠��u)ק�/x��>W�ᦅ�@���!yY�$����l�!;�+��u��u��+.��<���G��j��؊�8E�'�����m�X�ۯ�(p��t$��)�l�|>s0 �K'~�����@0�.?P*����3�����i�OO�e*�N�?���G��#��K��@�PT�H�Ai?���C9��<3?�(f�{����ONt�"B ��ؾ�]��9wᓧ���D%v�η�E�+�vF��k�]R$�;���КB ���4 ��N*�H�t���H��ힹݜl/k! +5��FAL�i��jlF�Z��j=)�:��29��d||��4/w���h�ڲ�|e&�s��ۻI�E��vl����b�y!��O�R�F�|�&�������P��C���d��-�?�T�䋺�4�g�[�A[�C����l�]J������
��ױ�V�#�T��ij�W$��\��X u�()�mR���P/*��!�����1��+�#)�yC�/z�跀�W �����lߍ�;�H����>_=A��9U3+�'�3(��G�G"���ڰ��c�I���;5���w&"�Tj�o=���}�� �5�o\��_�(�_��)����ξ�1pb__/k�/ptx�|�߳��}̌[XT�ǔ�p�-O�q�Ԓ��?�u5�D�b$��L�>��
�r�{��ĕ���8�;�����|TK�.R� �Z�\`�ò����u��??���9
�I�V�S��"m5g�dĶtƢ��L��60��^��G�n����X��d��G�����l봙����x�[���|��kiu�:�H�滿��P ě�"�.�UP!.�����"������u�~R�r~�H=�=�u����v�<�R�8��Mz�퍗 �.(��d�]ꒊL<���^(�N֐�ڜ��G�&5���$s�Mx��o�]��:����~���I߭؜2�`�'aBr]��(�$���lL�_�GS����nĲ�^��q�1�N`�	��sII������Ei�H1'�A%��!��8���%��rE�)@�����`R�����g��@�p>FC{R�9o=6���$E�T1P$�a��W9�7�c���Δ4&�5��l�ۂtg[�-�8)����u_q>~y�a8p@��꯲	"���x���1���}�M��=U�־J�J�=1��#�kT@R7~����7� ��V��+H�������˦C�4����1gκ0�\B��s�Aj�MǄ�n���y����Y�pQ�B;xX��%g,^�a�:&��]p˕��{�.8
>z�}-�g�:���5I��Fy=��o�o�Dn��$������>r��di�>�B�K��/��׌��v��U+�Ui�8�v�cD� ح�U�'U{���;����f�=H��L��n$����w�l7���播���.�h���e��TB�����	L��ڴ+����tP��eȒK%y�^	mU��ia�N�2l���N�:,���핉L�z8��X��eK�Y�+Jˌ���1�,�*1���)�{�:���X+����������S�w�~�r��H�o�
[W��F��O�Ώ?߇ŏ*�J���Lwu�i%�c��Fr����5:mu�35���$�S{���=I�c�\��m�J33�45nce���i�K�M�WMv��RL�x��LnW��%˰ |��Q�O�-Tr�ÆSw�8�Z���@8fu����-�-�XS�X�e��z{���w� LU�k~�Z�>�8vԉ��p��'+jL��3�b�D]��毌̯+ :��)=��
Q�a�I;0�@�/�I�mw�4�c��j�����ECU�5 ����T>��d�_�q6�� � �r�UE��6�7^�WB�jEq�M�����+��eW_��@Bٌ�:؂t�\��r���*X4yE�'H��t۵L��`�`H�k�åGP�3��5�:}V��I�(��u�G�W����=�ݱ�R��l�\�y��r��{B�Wۜ�S]%6^
�]k+�@��ڳ�i 0	����|	�o�����7ݠZ�?��P����W&����J2���23�FS?�U����2�c�_"���a�?���;������o�3��k�&�!G;`�x�!�Bf/O��q�+��:P��Q�N�9Q�8�Z�=�Op�g��b&1��B�YM>�C� ��YG&�{�ح��(fRZl���Ԧ�uK��ϧ��r��G0X=������o���8���$??����=t"�	�b��k�=g�b"B��n��s,r�����C�'_�k���<��Whu��>�9��L�+eR���b���Fk�ώ*`ю'�K* ����D�����l��Q����Hv�#���ؤ0.�����&htY�L��|}�~�}J��,V�������-��9,�h�
^���) j�d�	H��-K���-�By@��'������x��"��o�b�=��0�!��d���`��*�}�=�0���I�����_
�K}-���~L�g\ߪ�`�=�5�8R�*Y����z��G_��j�x@	L;�V9�d}�^U�}{��@�w׬0Pn��+�x����P7f��P<7���JNzM���$�F���YOg�q��X	�v *�d�f�z��^I��w��]ų�>K�$t�E��K�?�m�zWv��/s��3�i�}y�X�T`g6Y�F��?��Ua��yXp[��Z��{��}9	����G\�z���s�*m&��ޛ�v��^��r����ګ^�*Wj�ߟ���%�\,x�O4f&q�2�=4��k~33Mژ ���8�6[M�O B�������P�I������*t�o���Ѳ��x�C�g�I�#��<�6���I1��vtwY�W;q*�~+&�Z�a����>i�x?&u�M{ �}����i�kH�v�Qp��DQ�o8��ךCc4��Vm2ߤ���rN:���OW:��,MU����E�I�rt�vo͎7'�Q`���H����P�U�h�����A㖳>�W�7b�i���X�y�T�7G��u��\`��@������0A툐c��/n��?X1UU�s�=i�vn�@���)}u�#�Tǘ��Z|Hl��#"0D	��Wv��}�Yq�>a������Jn���J��|�ď�ŏ��S6v�5��.�+������9&M�������2u�����S��w>zVj�j0BY� � ?)���_͇�+�O�����<�j�}�@~�/�̫�趃'U�G��k;0*�����{�A?�[�?���;����#κ��s|�iI?���%Ѣ��_��rK�ه���m� }I\z��~N��w<�0U|wD���*�nl ���)V��\���JU�(�&�*)����h�P!�C�[�珖Klb ݹi2��9����^�!��m�co�ܯ����W׻v��,�7�A�I�i��m�X1��&!�6�gKj���R<�:�H����u.��:�:�y��LQ��s
J�:�* ����!�O_�p_[wB��>� F�#�@�"�ߺ8ie��Ā��w�{t�x��*�e\Qm�7R֭�hƮ�n�q� ���]�@�@I� oF���?�iuԋ���w�EX��M�e㘄(�\X�7sA�-�{�M���xʔ́y�