��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�ףe��	�A`�������K��xpO�e���ܭIb��]��͓�.� 7�>�9��L������f��KL}.�F�� �M(�����f��;�5�jG�0j�R�:,rK����AZ�3',�&X���E��L
�z�ʠ�����hF�L�}��x)A/���,�oӘ!�aO���`q����f�Vю�q�� HA+�h�	�����B\r$�
��r�����ǫ��9�Z�c���w�������,�F�#�"w�]���[8����Y��u9_TmFU��k"�IնA%+�W��z�h��-	��04����']s���?���?\<ߋ t"��附@N�U��s�9�B17�$+Zк~�|)KҸW�:,V�N��M$��&�qR�DR��yp���IW�+2b)�&w?4�����E�\O]#J58�O.t?�2j�t���U8�v�Bfh������m�*
 hQ{:��ebٷ��%z_lū2\� �F�s~4
a���꽧í*ː�̩�������]s'rϞ&־�l��y�Q�f�n� c鎬�Gf&���*~���R�vׯ]�����?_�U���p�z���Ȗ�eH����<�M#2���i֛��Q����{t�&rGĢ�̙O3s��^\������l)���K��<���hLx�:�_b���+	Pf�ɐ~������o����'%���������Z�*G\�<պ���'����Z{e8�4�����T.d.�f||������?N�{׎�� *'��Oa${��\^�JW���;.���(��G�6t���?��H|�Î.��k�Y�����)V��.F���/�S��7�=Ei��a6�l����}R�4u�N Y��1���ͳ:f�o�B4<�VT1�V�f��k�<�M������]��W�(��Q�5��az�d�R�k��D�@0ɍ�9d��|6�D��
�y�!���I� H�� '*���v^z�I��=r,�{�){�1��[�g�����>Wo��Q��I_���L^�/��$�A���KȀ��J%ې�v���A�?��t�!�<qq�b�	�t����2	�������M��IFG���Pv
e�y�eY�$[Ok�3Y�T�{N�H�z~e��
�Z��B���Aph�ë'�e���������.�ib+�-=�.�{��VWl���7RԹ��NZ�6A����F�&��q�GӮc{q)B�k���/?�e[�K����A�Z'Kر���An�1�.ۤdB�-5z-�Y��0��Ub,���Sa<)O�Ô�	��=�f��!�58o=���]�΂*��I�5?U�qT?���s�}�4{�A�L���j���ھ��u�<��J�;��b�u5ۭ~�D�)��� �U������p��rz���@B��^7��B�n�f��cT��/��f^i!��upA�ȕ���3Ux�쒼8_�[�;N��_�����Lsɦ�"��6��|���g�������>�Ƚ`=��%��sCP�˗a�%� >�	�9Tl��tL;���+~G�wh(Ê=
�e�!�G�ݑ6\°,{��*��+8�^G��7�7��j����m���5����W��]�ϻJd�<���c�p�\{�`�S޼���6���!<|�����4��2����bfb=�'�~�ވ�а���:��-5�^�������p��ֻ���9���g��R1�S�ڊ�������]������� ����(]6�͛5��8*����{�Aڼ�6١:�c�<6�8aj�`'��R_�2*�
���{/X�1eLJ�G��3����~�Ym��H��G��f%��ׅ�lA.C�M��F3�i�-�T���%r�폄"�虰א|�cWBכf0�X���zy~^*q��H�m�A�ژ-�H��"u���q,�V3�E��M�H�&r�啻�_b7�h~���%��;f�p[o���C��o��J����(R���nX�F��uۉQ����#�W�W�бQUp���z}��`�.E��q��ȳ �`�|�\F!�G�������MkR��� ���8f�r���g�ٗ�v��M�1���Q��W>�m����M5y*�4'�~�ɖ�?��Wg ��-��