��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbI��2��Ձ_N�RL��������lx�^6��ᗾ���V!���!�C���;s���S�b��PS�m��f�W���_QӔ���ų-�ؼ��j�R�<��bN���<#Oz�0x�2�j��`��پ�9����jt�`�tKȢ�ñ��H�x!q'�z#��eпO�%U\J�W���9���r�g�Cxy零L����_
ɏ���j	��
xS��􇾂u�=Iq���/��"�Ǯ�Ût��'7S�7�����e
Wvv+x����0�x�@-#��mbM��q@ H5C�@�����Ny��C�E7_��T���>M7�S�����B����k@���@t?޸ܬ(#�eLث�"�~_�5-ei�G��^�5��'�SFp�3�S���/j2����R`H��&��|r;�<Mo"#N��K��:��/H!r:J���`Nm�+"5�����x�	��Q�sw�Vha�<8(�� �QH��?�qHk���=OHQGRn��6�^�(ޏi+OҎ��@�0��n�R�Z��E݃d�kUY���Y��R���68'����_v�13P�P���9�N�.#��0�р@�$��X��W�t�	z<o~[8�#�,dO��{��eOϠ0A��u9 o[�o�)�n�[��,��ݓ�!�v���Ђ�����3��:ia�?Խ/u��`=�s�򍛕=�����2\٨]'Lt�Y�+P)�k��G��K�sIJO�U�R��S�re� ����J0V�ќI�@�o�"&�a�%�Y�c����L�g*k�o
8?������Y��g2���%��9A�(9h�~�_��XB��{�_����U|q;ŗ��16��@�Vb[d��T��f9*��^��㔶!���-3��uG ���0�����u�O�l��0%���/�Y�u��]��X�m�g1NbKӌ�x��ouM�������s�#��A-�f,Ե�-g���+&؂S�
�]#�� `g(_�2U8&�a�@�F�{QC�KH<s�St��\�O��鮩͏��#}�O+��|;^<��^xC�V�r�:fAnZtzC�[F��]��ph9B�E��I�YO~%+�����ᩇEwu����TR���r=�q7�G��NSNz��P�1#�.�?P�@�ѳL}1j���tw�C �M�J�k^w����3��N�<���g��s�3�MD'�3(�HhNB��!71�-����nk�$dƂ�}Q��۲�n�>6�̒>����j�"A/ޔ��E��S�4���ײQ��%��M���,@�Ϊ%5.U�d����x� �Ob�\B��,$�2�&��������J(���H.�,G�rܶ}�%:ʤ�y]g6j\�Ꮯ�N���6(�k�!�e���J2¿���QwDKu3ϸ���S�>�z'�KfM5%E
��A�y��*���ЩϷ�}��&,�/#���:K��q7y��`Z�Z������T�C'hO���c�O�z;K|�;�4��~ݗ�>����5"4xꎳ����+{]�e�l �[�O���0z.��d�#��=~�;�\o7dc�M��>D���G� [2Z�p��|R��爩|�{|/�{_~2�s|1`x�f���ڎq��,��2拌�f�
i�[��I���o�i����`i-HDyDȜ�w>��Zz�חn?fOpI��Ϗ"�6�*~m��o�:(�_|GOX17N�³,�6����y����T�c�W�����eN��ʙ����)S����i��Fbk&A��M4)�ǭh��%�T�vX���e  �+D����Q�b>������c��ĳ4�ϴÌ�Z��*NB�K�N4��qQ��S^���D�wN��M�B�V2�4�����W���zF��+�-P��ǵ�~ޢC̓��4��G�Y�t��-�nU7I�
�E�]�r�c�0SN?v`Ou*�X�F��8walj�&̀i3�ثN��fveD�\[K��Kۋ�Y(��qy��������#���ʓ��Z��p]ͮ�C3-��&)�sHV
�WϾ��G�\2�7��^ϊ�M`x	���=+TV�K�,�Z'X6~�f$囟=�b�����{X`�P\�|a`�]������u��x���_�ޘ }�`,��<�j� �th�1�Ne�R�2,Q�[�P��T���Y}��r>���׹G�s�>�.�X�"���\mƹ7 ���l��� vPJ��lD29�R<�lu�{�s̨�\;�UI�_!|�~Ӟfb�uZ�t��/ �6���(�B���=?G�����Z�����l
$쾥�u���e��v�GkK~xPc�̵�(~�ԙ���zC��O"��o���M�x$��@�X�Sܖ�[�`�\�	�����$�aD��G�4��P��~���R?Y6���z�^k�c�X����,E���v�ah����	�6��%[TE�_pq{���ݦQ���=�
R7�o���8D��IY.#��k��:l9@k�#���&h�@I������b���$H��qhm�,���'躑wqJ��5���'��|l��J�_z��Yh.ʑ�L�z�	��po�0�=�G�Xwk�塃��������-27^ڗ,���:h��\�K���j6���sf(l���\������6Q�*RB�rW��M6:������S�4�^'G���S��k"r��H5 ��~'�NL�d�� �r�h��1�c�Da�1<�����cַ=���APs��=��4^����u�����GCQ��6[c;np�؏� �2$뷀����R�� |�Q�-n������ܜ��|z�f��{Z�L���bx�� �sd�Z�/�4{C�l��p)q�O��E��m��ZGe�C ��1)��*my͸0s���n\�Ĭר�/�LO7�)Ə�C��5�K�]>�ʭ�\A���$>f�D��[��~�&{-�殠m�|,
��8j5�,x�����ɒ�F���0�a��՗Y�Y����ҭ�G�!�p|U�����Dz���X5��J~�g]�(J���կ7M�:l~'@i��;�!Ҩ\���n�:w�[�ሽFf}�#9�"/����n�-�$"��� ��1�yG/�
5�}��.!�x>��f0��&5���dq��6��g�Q�K"�Vک�
�!�!�tsƌ������e�[���9�08!�o���H�^	-���<=��ڥ+,1�ؓ�)!�2=g���Ѷ=������k8����9�+T3�ĭϸ����o)��.(�Rv(IS�flU��gHwʺ�6��?�O�_.���tD��K����LF��QE�\��!����"qL���I�v��2��B�C��9�ڧ^0HfٽB$G�I�N�c�������Ӆ������Cl�
X�*����J�;w�)7�9L�*%�0W8eV��̤�(���j�L�%����~����¯I*�)�iM� ���S�n�����-U���_g�O�M=P�WN ������t����Ц�7���#���cq2�ۈ��ר�K���r��U��Y�v����ݵ�"���Ϊz�Bs(��8����%#��G�&��X�S7�-X t#4 D���[�R��H6�,j�Ӂ�0���Y̿�79�8A��;i4G2WTH��O��m�\l��8׷�CY�h���aY�O��w�IU�O<<��,��e`g���{K�e�g�P&�f����M��z����&J�ܓ]�E�"k>�)!^��d-s�����sY�<��E+3�!�4���-���a�fKk9��9��������N�גPTp�ع���	u㛌(�9����)�(
�I]Mݙ7���$$ٖ�d0����L�+��ֳ2g|�a��w�ćX(��������49��O��e�Ks�,��oJ���k��Е�Kh��x�pdݷ�� q8\Nt�'��s�9�-�뀵�mM �e��O�F�<��J���y�߃�6cJ��6���[�#|8S�lKs?G�	qh�ذ�a�'l��]��Z&�8ʡ� �L��Ŕ����x�_�f���V��O4ۺ^�&��Č�����nc���V��dD�
gb� I���� ���Q�ϒ����;��hU�E~|�����RfūN�qy"��
/�$Be�)!|�8�g�"X��-TF�Q�o{�����4M��SIzk� MRE�ې}�|x�Nᦝ�S�alv�Q��3�!�ygjH�K�����4����2�-�Bc�� ���\|�1���3�L�;)�:�	����t�{Smν��]7`�Hq�H*c�|.w>$���*�\[��!�c��q�u>����Q�B�y�G㏠�B5F��DR�����,�����b�dd�"�<� �����W�f�e��}�'��8ŋ�U�7���pu!��~�*x�N��.���+k�&����T�1�!-7�$��Wk�녁��� �Eao|}�Ǟc4I<r��"d�h!���
=���b�<[S〡"H0��Ό�ʪt�9Bc�u����4]�z�whA��� f$=�J��E�@��[