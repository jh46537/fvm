��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ���>d���G���o���TOZd�A��-��+�A��#9	;_@�*h�[�k���p�>;�T�O��1[a���:����3_%k����!E_�^Z�J��\ǿ�g�]Z�@1��e�p�wp��'��P�ްc��A�����Kd�� J
x�C��F/yQ�ޤ&�wϓ�ڏ��(���p��Vq��FJVgx�)���lx��|h�2�C�P��&Ȥ�k�]�Ϡ;t�2�ͤ�`�{�Cz�������K!�#]�zjQ�PL�EL�j�0p?�3-��ğM񝳌
AႩ��P]Qf&M����H?�x�=W%K)�[�cE{��N���0v��j����5�����p�G�i��D�ȉ�S� �S*��NP�UO�	��ڡ;��wli-����/�C��^��Q&R��N6�y�0�*P���y
O#ܖ|5}�P���i[�-�LO��8H�	��^��N �Ew
:_U���~����T��F���Tw����vn�����u��3{�p<����볁_U&�7�Q�D��I?� �?���Daj�Z��s^4u[�b��C�W@�q1�o�1^�������#5��B�Ps;(�HF,���a��]@��R+��P�ZAAJ� i&�mA��d�cu�Y��Ey�g�|[�!���*������V�vgA(.�]�3�H����9��OB�����\go�ӏ����s�}�"E7�E�R3)��"�6�jd�-�hF�(#Qc=���g�M*��mp�Y��#���eK~i�Ǖ����:��!a�� y-����%SaR�YP�a޹����ioN\�a����ؼ7���fF#��x&����d���S؅�Mr_�Q����k�dM6NE������]2��kZ����F�s�R=5����6Ɋ �eF�%r��r�E��B�ɯ��A#��	�hL�D�_���2^�-��y$˱2M�������K  η���.�{�����S��4�iRuB���1������	:��!��!�����羪�+G�vZ���k�@�6f�rM���G�/[��',4�Z/Y����(�K���5��E�ٹ�֥�R�Y2��K�O^�b]7�Ug�ľ�3-�����@\���lO���mK1֐��8�}����V
Un��K���+?�L,G�=k�98?$c�&��k�9+�V7��A'���ZN̴rN����O��?�	� �x��*w�Ɓ�MI�r�B���W?Q��c���FW�����P�����=�l�EԋlrtwhHQ��4��M�!��]pMP���_�̦��=�����ￋ/��$�IJ;��A>mjz[l�t������@��+���`g�6(C�S%y}�(�o�b��(V�p���p!��-�0 ��c�}��FXm�D�c=]�+Wy��F�'�f�;~���P�t�����4q�L�>`��C�w�G��g��
0
�8�&�s�qw�D�	s�|l~������|�*e�l����1�gP/���c����������Ŕ�ȓ�%���AV�/�󑺨�a��-6�tdm��֧T�Zz�Ie�fllJ*��R���?]5�5^�}�_N�#N&;N�Ji�Ag��*�n�%�iyں�4��,�ƶ��1��S�r����nn��S�h[�o�I'���Ur�d�����m>4Y�N&TgB�	M��|2((6���c��5/]4�v�0>o�э���fK�eWթ���7�z���􋍿&e�gTW�<���:��@C&/����aK��2��������M&����L$-���B���I�U{�J|u���6�<٭:Wn�z���tZ>��!�dU��p�_�M�	@���C�7�z��^�ě~Q\��n;�:�.�n�Ջ=m��.KRb!�zSJ���DM~�Qd@��y�^���2��$w��_�
��$�DS�52p��t1m���,3t���H���qE��Z�@�ࢪ��$�a����5�R���09�!�&��z��o�_1���i$�	S��[D�����T]m�=��*��t��;1=�E'����㄁�W!/v|hvQ��x�t��=��J��j��=d�
���:8�H��4��8��-��ye����k���/P�Nƚ�WlŖ��y�p^�1m�{W��kC�lm<�rEG�^���;� ۑ6EB���J+�*߂2i��E�$���T�K�f�����r�
IBKu��� � wI��V���Uc��>/�����3�J�,�J�Gg�M�s���`_�~+�7���Z��.G=P:�B�o��'ʵ���o�=Y��7D||�<FDN��Qg� ��L��ԍC��;O�+w�o��ش`�gH6��]�����������łE>O~���5 �M}-�����8+�O�%�8�[�D���7tS=l1<	?H:�#u��늸ϫ��̓t�e�i1^��Cy�,i%�!�W�X�nc�Uq-�Z���0�֞dh��b<�}��yІ���tzƩH�_�þ�|��h�Ȉ�_�MW���Vg�d݌)�A����~�v�B���Xp9Y�Dµ��c]Ub��g���ۚ�+iP�N�hA�����⎋�<V������~̹$� �0B^.��W�V0�>͆�ћ�2Z�φ�Fˣ龑�fl��jK.�Bǈ�z�%���B5c��Iw��&� ����te.�W�"׶�Z��mI�-X���_��ôv������`�W� zf����u�q�Ƅ�[���	��/�G�2��6� ���X�p85�]�D�,̹�"^]0�a�Xk��"��h��F$F"v裤���5o��B�3���z?���]k�S�GICS$�`�/���z�&�p�)H�2X�Ž�'��΃u����M��$Y?џ��}[����g���"�Jp��*ZO����w]����@�z\\���w� "��Z�fL/�5��p����:կjQJ#m�C��
	������.f"��vQL���ذ�r��x�Y��e�D��⼍!�Mq�(H	n� /���Y¥�;Wx����Y#yT��)<k�s��s��v](�A:2�UI�L��^MD�c5�|�� �i�D8���Lm�w�@�_g7�I��u�_�S��iG���OI �Wը�ɸe4G��u�v�ԏ�xO�<�˺2��O_aZ@���%=Ĩn��:N�����c��4��*���kF��A�e�������ڣ�et�]���D� �pmQ�ga�<DSӑ�Xp�v��!�gW��X��б�뾴0���L���A�.0fT	�n[<��b�P��l���T�����~;L6�M0Y�K��N���k�i��b���aīkW�eO2�0��E��ג������ɏ+"����`5��RWm80��I�8=��S�֧z�A#z���%� ��s?�M���y,Qu�=u4eMTQm?x���+N��_\l�b���XU��o�U#μ��r��\8�J5�@38x�u��S�z����h���֋�Ϧ#��s/�T�g:��?�Jw���*`\UiIq��#�]�����5�x�
xp@����FI|�i��_�%"
~�w%P�iL�7\k\ggJY��c=� U�G�_^�:M �$Ԝ
�y��T1ݼ���@:P8�Y ���奻�h��u{����(�^� ^�f�s+L�3C�:@l~c��n �+�@r�u��?Lm&xΖ�-tʸ���Ғg�y|�T+geg�la�Pe��d"�j3�<�H��I�&���W����7�����.��v)� `� ���]�G_VCw H�|n8�DqKW��~¡O�v
iE��ͥ.4hZ�1T���!>p�9w$g搰�X���d���$G�c�QL� UzZ!��Z�A�t�N �R�n<�����N��s���"$c{�.�ɩ/����\�H�Sʔ�f���X�ҝ��o��	0�8�HT^�=�O0��:��}�0Yn��G�e�l¡������w����l�;y���T�\O�]�ed&��D�-�5�L;Z��U��
����_��/g���z����d�I�Nr׫D�9�P���3C��m��\�,�1z�@�+�#>r��('}5H���ڽr=~��R��b۟��#iR5X�=���(j��K>�\�`mK=�	�ڿ�T)�W�`4�Ȕ^�B?�32#I(A�N��d�������m=�6:���
�	�]!��Kڿ�6�.�'���' p���3�%���Jt���+��|G��'�2g6��4�Ժ�w�߼m�m�����F��f^�BJ���^���-���U?�=�ӭ���3Ȏ&���^N�����QV6�A䛚�����:��%��~�B�#į�^��,ʌ65EZu��(#E�޴��:�u�x-�Vj����gU��60��z�h#34��h��.���rk/$��"��i����h�����a�i���`m�7w������9�"�S�eF�+"шN����9���rrD�S]���^�M��6뮜2���=�0��xx�r�,�e��p*���d����t�W��g%��(�2�VA��	�5�u:��Y�D�ωS&�e;ޮ:U�����oI
V�1�����s^N���P�c��ws��B��N����붦n[����0I3����ft6=X:���Kλ�u7Z��m��Xk��!	��I�8:���k�l�y\�?:��V\�:�OMgj��x`���H	{s�V=�fE���j|ț��܉�Q�̈R�%�/m�U�s��-SRߑ��xhR�)�S�W~wY{n��ZB��ֹY�_@�E� 4q@�{�6t\���T8�7^�]��}
�j�����59���^�8�Y�a�E^{���s��D}���V�q2#�*IY�%9�K�T�@�[ u��.��u�אs���{��жC�CK��b�#(�R����E�х�d�;j���RȞ�M���jO�/9\�Z����T����}y�	�3ĽGY2���t���B���s���V=�텂1#����70���QR�=6�����Ե�X�{,j���0���/�b�s۔ҏ��?鶖�/��,��]�,랝þ8x��Q]�H��↗VB
�*ǿ�dnA �C�ϒo��^:{���=�;41ѯ�[!���QL�Q�t��;�wЦ�8o�nO�ٌ�J89��d�Z���da��2'���u|�H����凬i����}L��î$X�̐�B��n�c�?N�?���[#���6F���H�˶�v�~/-Ъ{��t�84���|�x�iqp{	���s��R9h${�X�C�}�XF�v�!�/
�K�u�FC1�#����
ޔ\�=2��>-$���L�P�\��U|Cj�����J�_�PWv_J�LE.65��U�)�>Sv�`��I���KMT�g����E�]���A���s�ҸY�W�A��a�U~�[^H-�Q�Q703�i�����,}�Y�S<�n�(�6V!'���UPa�kk���o=E|"�>(F���d�s>��ߠ�K{A��|��lu��Wڪ�$�$�-�>A�~J(@{(��8>1ϔH�HJ���c���K0?��kI��i����h0So����3p�3��%CX���Of`�P`A.u�)��|�V���l�r�{�+S���9)?���ۆ��/1p=L�訆�h��>;�G�џaR
��@8f2�6�t<Q�^g|J{:�06���Bd��3�#�.g"�nDxF76�E뎟�&��؄o�U�X�:���K_�L8���Ί�R��u�f��*�v��\�RDBL�v��m��ԃP�)�^:=��׭C�tg���]�%�RR׭]D���%���&���g|1�T���@��RMgf�����Iy6i��F_{��\S���=#�C�{��q�@�L������f��Og��q��W'�G���_���
�A�C��=�}�y����$'N�:���ۤ1�=F� �)d2EǸ�����zΈś��l������%S��k��*��q_��N���ll)����$=�A�~.���l��su�$��E�yѳ Ջ#ix�M����,Z�*%0bQ�$E��9���yU?
@�}]��B��,���2��x�]0ɟ$��v�pp���}��\r��!4��VUǜO�H�@rʀ��[cʸ�Ϳ���E;�^��� s}��{��387���u�����&zh���x�*��U|\���ñ���`�������)��Ə��ܾ?)D���+��o��f�X��vmz��	Q�4�=<��C<��&� \\pK�SՆT�ʶ�/l��V�i�/���d���iO^?�[��Q���B�#�WY^h�$�	澥�B��qp*�i
S��qkN���r����K��Yy cS*�~�g��Qm�Ɍ�Ǥ/��t�D"Iݖ�iEe��Ϩ?�ۇ=t����#= �@_<�%Ld�iJţn@�t��!ap���s|t;!<U�KH떐-�5�ym
j?tqU��ȟ,X�U5a%��?����͗`��k�p ��P�%VR�nP�����l�
�~f;xAՄfYW���a�����ξ�6����C��^�`�J��}��ʀ�c�AX��5ǬZ����@Q�?���,���kB�V\�Z�'*~�V'm._}���N�pz�).$�N�q�Lӂ� x&qV	���E���_��I�u�0sp\�@6��g�q��c"ބ� ���Q���Y���J�6�J�`��I���y����}�j3�ݮHz����Q�GB�O�t�^Imi�}�/�.�[��T���mbs���ѳ
�zt��$�c�ې%j�:沊�>Nf�N��܈[�N�#����;+$�HyWD�`�|���{]�"z�����pNo�e�G��:��I&	�ρ�%gvnoӳ�XI�j��^�'�u�ȨG����i�e�ұ���5��D[�z�ʆ��OXQ@�`�%�eg"HR[�/H�0)��@���<�<.g��#��#������=҃��r�MVT">8�S
_'�V�V�Ļ�y{(�>'r	�	���G�/�v��*�Y�3Ċ7��5�T4�5���r�]�-�|5�����=e2�i)pD/����p�8%�������#��^��}x��D�TZƺ���I��"�Y7���I�6�SC����hw1��Ӱ�%#]���_;���eR�� p��O��Y�d�׵��]���8����Z'&[�ix_e�^©�d��Sd2�m��������;"�p�,���->�ǣUf�8�C�981g��,1|�{���ߟod��m�:�v"�D��k�&�2�2|�i�\M�G^�}�19D�N�$#��|\�=����r�(V��<5m�c)!�v���XR�7ԩ�t`���ZF`�����v9ƫ[��a�QN�H����񃂅�L(������Zeۑ, ���O�/�K�m�������LW���PQ������ȡ���������b�sG���R׳Ϭk�ӈ?2��H<�4��N�Xp���gQ�Ռ�QJr��0}���`VS�lt)Z�k�V��ڈ�����RJ�u)�Vƅ�\!��#.�h��Xt&�`��BǠ��0�,����r�	F3�36�sĚd�'�$9�)")��l�O�IJJ�K�r�{waxRm��\vNx���p��h
zU/_�ۢ̻��Ći�#��D�"���o��_D��	\�К���ns���~���X��zC^����%h�.�Tu���G��L��|�$���t��N�,"$����,T��Z�p�(� N�ڷ"F�@5G l�>�c�8��|_5�y|DR����;�����r)V���D��k=8�O�l����1�?Ҷ8��N���-�Н�3&S6m��e���8U����=�b���f�ro0Řc��,uSܩ�ɓM�UE0�xS��tm̴k�r�`�n��:�}^@� Sܙa~��`���K���/�un��s#�ٓk@�@�����)T:��503'e�ί��vC\��P�ma`�v����xfP�4b%���w��!9����s%�Z�g��S8/�Hɝ*Ou߲�?xMg�Ɠ!��N��Z��SH�SM�(�2�4�Y���s샅�5�i�Y;�a��M�n���d�5n�ӆ��x�y�����iیi��P�y^1i�F;$A-�=��V��	cͷ=�lB(P
=��@�����!�؊�y�x��Q���Eq5�ؓ��4Z�������*��x
�����8�LZ����[9�~II�e�$j7��C���4���ص�R��w��7�!]_��c���&�
>�s	ۓI��g�'��Ƴl C;�� �b$����'�&�2a5���aЩeYk��W߅��=E����v���͑B=�d�����|���Q�ظpJ��ړ���yR�.�c��%u왔J�\M�m��� �Ʀ�8�	��H�D7�Ŋ�¹_q��DC��`����[h�=xYI��L��w�k������_�^o�*�E-D.>�is� b��0���e&�����c)'�T��'Ĕ�;����_v#-'#�ܨ�*�3tm%t���Ó�ŷ����X�]Bt���p��kx;3*O��ּ#�A�g�e�x5�q�����0Uw�j(x�JT����0c)���-�J:�m�x��s8)�w�����`��
������PiE1��r)���d0w��V<�߬47ɲ�����'�bP��-c��#�wS�T� ��(���,���Q�d� ګ�ޕd�
b�.qP�{�g�x��"Y,.���a�����J5��O�B,΢C����=�ݪ#��~2��r@��y�y/����K>I$�e��ܙ�bBؔ�� �qЍ�f*\c��o����(�L�x~�K)�Aᅘر}����_�:׷��D����4���=qg�>hxI�2���+�����ـ톛�'��V��{_a�>V��ɖ	d�&�a�D�5TD,df���֕��cu�q�������<�~mV�H���* �	� cKH�,R�%��I�²���t@�,@M�>���ON9ldg�94��[e=�0�)�O`��k�����u}@�Ӷ)D�'|�0#t�ӼL��h@��q��(�]�.T7��I�	�l�B���<ઊ~���{�a1�9*��!.m�ww�������j���r;�d¡�����~�9�̝�"3�@]���\>�Y��&�"U�6S�=�c��Ƈ�,v�#B�W��!�9Jܧ'�t�&�h�T�\�ӆ�[�i	�����ɀ�����4��.G*�@)�>S��I�_Á�	Ou&��N��
���}��T�a(�)���r�P��k���|�h�Ք4cM)#0pd>uPW��f:G��_1f`�s'�m&�<[v8��U��#-*�LS~rD	�:e��%�m���č2��3[�4���p""�/kj��E��H���%�\��C�~�p���=,�$F�!��0��8,�G�j����O�X9��$|tƐ]�ޅ�D�)G%�W�w�_�K���?�0��4��+y�&���yCeM��U6#5���.ݽt�FQ0nq�C5l짆�@�Z�^ ��:3��6:r�9*M8)�Mʵt.�J`V�s��=��R�m_�1����\��P;�2�O��6Y����H��@a�su;3;Qׁ��j	�ӛDA.�!ʆF痹��nѩYt�g��%Ј�+�ѱ�;�0�v1[9��8��zk�SZр��v�*!"l�����@�ꏾ��nϋ�Ԕg�"�V�JA��<8��Fv�ԥ=�����m>bQ6�4�����^����&���Q�~5�,O�M#�KV�4�m���!	ի�K�m���F����t�m>����v���mA�>�n�X�e� o��3=��	�&a�"��JԜo�wv��'	����׸�$��x��s�k% �����W�m9tT���SB��8��>!D�7��̢$>0�H���~������#�@&�	 �A�� V��&W?l��f��=6��n�>���Z�ޓ�VJ�v���|�����Aj��Oa�'2M�7����d0��fd�+D��`0�C�HHlN�ޘ`�Q_�U�d0\X�M�vzo/���eH6R@s��De�K�O��U<˯F��0��t����l�^�f�p]
��R��;b�ر��du@$�s�P�M�B��)����F�� �eP���j>��slX,�Q�m��*O�-Uɼ�4�Z����[aMϾU��<P�YY��+8���fSTϗZ]~��g?�+�CX�����!-����OĹ�/e�˔��UXvKX�kG�I7�L���p�~�T������*M�բ������R�S؉��D��]��a�˗.��B�M~�����,Mj��]�/��Z>���U��L������i��Hw�C�A�?��G-1��q��>�e����_s.#�ɦ1�1�,��d����G�H�y��g�F�)�n��2(�ut;<>��t
4��a���	Î��y��F����Om���E4�'��ɆX�W�TS{B���9��LI�ճ]0d��Mԭ-�$ܒ�j����&d)wݚ����eWl�S��s����|ޠ���Ō���mt� ��ܜ�Gp��#Ժ���R��ú$�k�7D�p��� �Ѥ	T�5��5c��P�ֆ�~�aYU�J����S@��C!T�w��� d'O��9�����g�>��X�K��]���%�c.H�U�g����$s���M^��y�b���粜�������aa��3@q�C��������)���.�ȋ�Y��a�`ZV�%���I<"�tV8ѝ ����Z��` ����$M� "lFO��O�֜$:V�׶�>���� ����&�z���0T�D�3�W��8z%[G�7��G����0�T�͟O�E8��14S
#TE~�L���]�Yϣ�f���������D�����p��e>`Ô�Xa���٣���X� ��Eo8�9=4g
P} |��O����k�PP�&�N�Z)�V�\�.gXX  pW��3]�9�O�)����c�<6�<�T?�|"C�t��2
�s	�v�f;v��B�o���19��m�����*Ə�7~�q�z����MQ�7�\����˾��2Z��������(C6���,{���Ϥ�FXZ���_ԫ�ӆ1c��)�y*W�ճ�_��4�6�9����GR�?J�$!�r+7�R��1"�G�Դ9E*��`��ױ�H�s�㪼\* ׻�ѳ��Z�R�)9wG��[���k\�v�"�)��Ϟ]I`z�]	�p-�K>m=���$� �s�*�%�Y<]��F_y�:��@�g����u� VG�d��[��{���t�M��
�C���C�pP
�af��;��b/>'_@t>V�<�إeG���]PP��ץváJ��P"��i�m�(ƍ��9�}��޿k<�f^B�i"j�lM!�LIM>�Tg���$_�Ĕ�$ĤZ�/�lMm�H�\�w|��J1=�G�NK��
թf�O�0�"��:�]}�P�%!(i�a�1��Kn��S��(sZ��3+2���P��I��No�sz�hЏ1�6�����Bo*�W4�]~�K��}�_X�P��h�js�T�1�V�)�hn�c��Z
��֢\h���[t���VlSp0(;��m�q�����9�b sqm���m�[����;�0ox�z�څ�S�@�P��T�[;�:8��d�%��8��Pt�oRk�F�aw�8�GA�
�w�%���	0&��O���(RM�޲~���@(��Ύ�퍵���P�սq�22X����f"�[�!t�_����:���K�VQj��N�Gt���n|4���m張���z&�A{<'�����{�.��|�1C�(�tZ	��"rw:[��u�H�+#����m�������*FlMJ�\�n��Rc�R$�:�%��yO/��-U��P��I/K�7�iIb�;#�ו�2q7i�LF�$P
٘�i(m_���ƫL���҃v;<�����y�wo�8�^%<z�~�/F~�I6����z���S&�H��)h�K�ғ���خ�q5q�\M�$#���r��g��:�lߔ@��r�X5��'X�Q�K���ص�x�	���s�����D����o����
�e�8E��h!�YE�N~v�+p�!*p�>�`J��Ά�:G��)�����C��)��l$��%tL6 򵰢Nr��r	��[��qӅ=N�Mk�s��{?-|���]9�#D�n������ʊU�t���� ]s܌O0R��l���_��;�>*8�.Gd[y�y
b�ŭ��cf؊�;�8X��Lh�i��`�Ε7.�vY[��� ET�sҿ?O�:�y�#�X�#�@Z�P�D��QcSL�C"���7�znb���a�P�kk]�e X�0X�t���tvy�i`5ާ�*�SZAs&���!��D�f<RK�g���
YF��q[q*��8CQ$C9�83?F����{I�)���~�����Y�>���αTh��띎�6_怵vu lQ0��l�(�t�����k�+b��=O���ez/�?C��@]����B�WN�՝Q.� $T�x��&����-��\���� �l>k|k$���].^�M�C8$N�{]��LKݑ��p�'�)���f�D�%Q������E����'�K���i���8�X��ʹ��A� �k���90�#��[{s>J)���V����2�v=��� ��w:��/�/NnPJA����<�.�$�ߖ���$�A �Q���$����W)���-�>�}����|��c-�!�g	�݌�Н��Q�?�N������1an[����%�^["v7bU�J-nn�	?Eɻ-yX?�D�X&�^Grֿ1�_H�l��[�_la�ɋ�|��O�JH�?�MDXU\��J�t~�9c�˰�����dbmĊ�H$�[B��K�u���@��|�Fx�.L�r�3���s��G~��F�l��i��O��E��Cy��qа�!���`���v�3�K�^�dp6��vc�]��i��2q9�ӸćxZ��}�]�h�/�m��,�>��]϶)�.����R���i=Ut��3�^���
]�t���$�_�&��f]J�$X��Z!�~��q!����r��P� !X�\n�M�y�![Ty�w�mY��kO�Ñ�l&�K8�E�Ϲu�xA-غ�}2��F���Ȫ������y}��f;�`�!�[�u�T@��K>�5Zҷ��6|�έ���
��m�(���r]���J��k��N����
hHw��ч<����R�z=)�x�>����H��D���_fA�=U.`�s,eŉ{�	���p�$-�L��R��d�p����}�'M�~�PLw�b��T��%� _T�̶�/��E��JI�a(4
�4"ee������@_�)X�-*��Gs�����9�&J�
x���~Ռ�k;ThG8X\�2���h�Qn�m` ���z�[��g�?�$1�IK��~r]aQ���^"��n<���A�z����#��'e��h�*�}�[�t��cIx�p��*�{��|��|���3Iҵ�����?-`��y~K Y茶�jr4����s�H��d�
9�L��K� �jt�؛2�!X��p1��pS��1$ۏJA��։�m�RSv�GI���)ۋX�+}��E������TWr�L��}C��� �H��i_<I'�*=f���ѺF�	H��U+��xp���K�:��K\Y4��GvCf�Aؕ殉���w�
��u�/$�*!C}6q�BIx�K��O�g�#�pOn�OxOn�da�1i"�A���ϵ���x �u��#��4�^x�[�g���tn��������0e
5Z�ϗd8������n�T^�h�5:b.�WT�1��,�3��KyuΖvHǋv���q^ ��v�^x�(m���F��nӀ��ݳ�q�E��3��8TI}�u �o�;�;�����Z%Gğ�b��R��;��7f����X�tt�[1/�ۥ�-1{D,iZؕ�Y��[_�Z������1�0��>�>	\j6t�i�x�������d����W���.q��~S^���k��k�➴͗��0�0�MM��`��fm�_M�v�/��,=;9e1�*��O�3���+-5��\�-�τ��S�������q���(�۸�pwU��,�[q,�SS,��	���VE�Vn������9촎޵��f�.K������(7w����Z�Y�:軓j�J�t7!���t<�~���;�58��`֡2X�X1���-�ߚ|��E���E�1e�)볆��4'��(M�̀VL�d�w#�șv["z<���r�����SO�Ҧ�������AC�	������Ƽ*QI�J���h5�	�C���}7�# �r�3�!W��{��A�'�m��ʖ�^I
�W��S�8��ir��
|`-'!3K�r̺��>gz83zԸ_���)a3�Vt賩�}�^��Hc��/x4YKKTyOǂ܅xsu�;"^(����?���=���@��iz��9���3kU�;b�N�0P��S;p?1�M:���{1�$b�g%]\i5��f���t��2�e`����w��G#�#F�R ��wz��龌c"�Is��f��I.�-�[Gw�Ɂ\,�&G��LE�~ �P����8�?����h�w%B^�Cd�����#	���C!]r��	L%��|h���QG�f6���U�}��T�y�(���$!�*�8�p �L�ET=L�͝�<]���<(���a�h}�� &������ư!k�Vh|jj�U��4����]�8��F(�]Nq��ǫ\��r[�ū~�@qk�
̨�bc���oؙG��}"Qo|��<3��2=�ĮE�'��AJ�-L����,at'�/�D,h�y�N�c�"�j�I
��!���ى5}6�� Ծn\��+�'Z˨N�t˧��=��Ů�3�)j����cnp-w�� �uJG_\s�E���!ƞ~���B����V�% ������_N�<��<��KNq:$:j���e	���TMD��l�EЬU�?y7v{�40�<�l���v��-�̝lʹ��	�s�bʸ�3+�ye*fI��@�<'Wg�⟳�W�Џ8A��]'@}���al�Z�.o&��.i�tx���d+�Q�_|A�e�_BPw�4���!b���OD�糐3 �-��m.q�J��R�Z<�H�#	�IlK���q
J�/(���������y������Ռ!��]V���TW`��E�B�h����wsxc��6����<{��[祹OB0q���Ʃ���J��"/xfU2��| 5�2r�{���7�@~wn7�:a"u�]��Qk��R!;>�[�\�E����Ƙ8�I�2z�5���(EpU��|Tcs߯x����1��t�x<li�6A�"fǄYL��l�����c�BY�������N�x��p�?A=�C[�[X�/j��݃��<~mZn�y�ټE��e{�ug����HI餬m�<6�+ezq,C���?c����˕�&�	���g�R�r�<�&�{�a��)�~ě������n|`U)�ʯ䇡*R@��a1�\7��Qu��� ��� 4��χ��#��'wc�[ 1�M,脡]����&��䅮b ������������$����؈&^�N��Z���Ѻ?�&0��'��w�B�8��F!�����q�C�]q���i}򵆏}��o^ȴ5�51� �]��,�V2D^y�[}(zφ��N�U��O������2�^��P�B\ks�PB�d���ܐ"y��M�����r�c��0�H�Nsv�s%n�ML���;g�Ᵽ,�W��9�t�D1W��V�'�#�b'Ѧ�����1؟"�0~�z��^2���ٲ�"� rٵ���w�������v�yQ`j���>T�/��TH�A�/T�B�@'����ۅ�� ����Y����u��3#�&zQ��@����|�c^�"#n�q����s��х@��Y�`i�szHJ��ɡpz��1��@w������G	�89�3�Ą&}�z�;
k�K�����}�P���h�O\�_.�Y��j�@�Ql\"ԭddݩ, ᦧ���I�۝�v*'��^'���A'g
 ��4��V�OY��@s�/�$.���1�#�:j�]�W���C��`�E%aG���K��$�{0$��Q 8t���3��n���qV^�=�,Iߡ��m����k�>8d̙��o��hI2�s=�"�%-��F��{��o���k�͌�ؖ���7���f%��TeIHQy��P�E�
s��8����&rȺEL̨ը	mS���!|�uN9~��*�r���R�v���~���AէS~3�/X�5���3�',d�����f����K��_��C����4���i�_��K����@q� �	a[+~�@�_+YS��ldT��\�����1���y�?�f�&���JB��ǹ��N'�.�>��Y�g�N
�	��{j�Ed�"nG��{�ӷ��0�U�*�5��� �lo�^p۔v뢧b�l�)������;
�lIؗ�9�T��,+�����$��@��1aU���3{�y���T��Y��M��P`8]�5ĭ������Y�0o�`E4�����&v����WއFRUK��&,5�u8W�nm��-i5Q �2Jx���z/8~HJ���.sV�=���w��A�+p��u���JNHD�V��}�j��A��:��3��I�y' ��ٓD��$���ڻpJ �� h�胍���{Y�Q�6�I�o�r���`kw�����f�S�>���/D�㼭��oa�E��-3�PȒ�|~������+CͶ���k�WL���1Pku��z�8�M�٤�-�h\%ºg�d�Az�uM��L�jsv�Q�f#��$K:w<�ʴ����_��I:�h ����!�ѻ�NL�e}�gz�jD2E�B��p�c�E��.��`�����5���@���(fq���w����� ��p���	��rd�4[&�A���,}c�x��� �R��_2����q�}?Ez7/�]�Q�!<�S��I��u~X�,�"�J#dl���Ni�-U����[lC��[��B=�&��y�5F�v���S���u���;a��C*��eŰYl~,��*���v���ޕz	&��E�ko����TP�����ʗ=�Ҫ�"��`���/?Qr$�Z1��L�Z���ͥ�*��Q�<R��T�>�09м��E��u�I�}�����N/I[n�k(�8��}L�,]�a��FbSU���N�;6-/t0$6f�{�D��n۹��E�kz Hk;ah��]#+�\���׆@x@�Yo�Z����/G���%�91��a��=�&m	l )���G���j:��-��Qz�68:|2���$^]c㺊�@�h|	�ɤ� 2����p�/	��1�4j�]�1�GZ��p����u��4N���E�m��h����=��EtX�j�E��9)�dM%����j<J�~��'X�ENa�9��l�����mN��ߴR���3�1��h�5��U�������X�`/��+�U������R�f�rJ��(zS��?�srr�jyza�x:����2�$����AS���F-m�<�mn�{+	P�-q|=<�g��VGwv�j��C]]9��Z�m@����"��Q�Vw|�p���5}]եC�6N8}�3g�OD��?��/P��r��鯠D�˩��o3��֙��=c����9��(�п��L�ܰ�K��ݣ0�"䫠�ϔ*�MT�T���q\�^�@�h���u����]XҼDrP���NX��JK��_�I���ܹ��F��c�Z�WkfX��&��	$b\����DCƽIlt�2M̦� ��-Z��$أ�6=珨'�\��J�O�֪�2p������GgF�*ώ�j�%^�Rb2{O��r|�#�PF q���~�_u�%��U��e�JHW~�$~����(-�=�n+v�g���Vȫ���#-��N�S\�GU�W�M���[R�cگ��t��[��U��}�Ϛ
�fkt�wc��1��x�b)�6��y�c�=��1N_�Ԡ|��！���W5�?P���O��<-Jps?�C���h�޻o������@����w'B��o3��������ѿk S]�ǭО�/dx��J�,�E�h(�����](𻔟�<,-�[o+�K)|�/@xW��M���g5�Q�p�����#4��uC�� 1P'�]a$���"�O�R��{��
�7�g��[06��C{D���t	��@pj\���H��������4"8/>���=�D��� �����E�g�#?Y��D���b=]k,��aa+K\�>��J2�l�0���L/��wX�l�ii�s��?8v���5�ͨs���]����ʞ� �q K
t��E�?pLMTQL�A�	1�>kt����G��.zu<��w�s=w�K�%��k�8�[��1��f�oÁMKD������S�i�n�᎗N�����P*w��U#%Vg�fAE[�}���v0B�H�A*;抧��O��K��Q&V׎e��]�MĐ��Jx��*a!����FPl'<Mc{�x�~~��e{9����G����~�!ï�����􏝉nz�1�3���s���Ʒ�vU���\���0�Ϋ�KA�~χ���k_'@�Xƶ���9�� ���E��D�$Jh�>y���I�&PQS?[�w�jc-2�T|��㛒���{g����H~�ݫ𸈩�j7Ϭ���(H��>�1��ezv~��?�7tO9p�	�7D�~�њ���B�|�4$�w�/�Z�L�Q����g��'`f�ƺ�n,5��7�0�qJv�$\l0,9���an�>���+�C'�ky]�ړ�1Y�*�p�T���D�5]z�$A��g�?�|he�pP���ʘ���{��t]-ϳjn�2���h\\�ǐ=H�I�D5�����L���TK��،ht���rͪ9����uֱݲ�a*-�&�0��'T�L6���׻fg4��+�dC�Nc�wnL��gj`R�:��(8�>�(׌��
����I]��������nuAri){���̭S��=��#9�s��A0�X�����w}1�YC�$F��^;weĂ�6���}:Zp��7$� vO`h�d|�	��t:��I��3���}�L�k����m,���.FS��^橉�4�Ϧ�Ip��J�E���b��3a�Z5�
�o�ʌ���Fv�e��	���v-�A�P0/h����
��4�u�W�az�|0�崷q�>��9�Se�W�?&�X����{q~C�{� e������HJ򐒯�l5&k��[�6	h�B����|��{��z�����C��̋�_LQX�^/��ZUBS��h�n{K��v��xN���e��ZD68�W2�:��e�X��Ð!W��MJ[&���Ϛ��o�<��_�Z�mύЗ�%G�t�Y�Q7KPy��C���Q�2�O���/lP��s�$�b��;�N�=�ʪZ�v��"I���f�͕qOT�I,�x;$�9��[��n̾��wd��c��)�Ji�z@n޳��2�ˇ���I0�=p/Y@?��������,n�(�>/���~��L �y��q�{��!���iq�Fæ��Ձf2����<�*��k���7xV���]3�����e'��c2�YP�o�g��
� +���D�d���������+/0�!B�sA�!&�sv��u��7��q[,p��s8;˶W�T�&2��*�g�[�GZ�RD.O����a��,^�n�;�t��&���.7�,WG����i|F5��B�1�S���X~#-�[�R��s���ƌb�{W�#� �_�R�Ziq~(X�y�cK7z��.^��z��~�b7n7���~�/�b߄�����C�A�Fe��Eb�$��&c}�n��G����6�?��bX�J��MÑ@P���1�-I"�%J�)�O�g��0"W�����w�݈T���xx��/l��}���1l苻�����e`�v��ȇ�?�p�S4���uH��z{���h%���MR���Ms��$��^��v4/���ll p\�0���{�D���Z�`���d�϶g)oC�P��z�Զ4�$��gz�o���$��V
}�L��ف�f8`��~t�	����j��k�'����,�~�՚�k�x�}�*a+!N��V����)@��"�8GB	��lnS��64=�:"�Ι�P��u蓟�s��Ґ��	�R���[��6�� ���ݥ?�N��xF�����P芈z��.l}��.y�G�!���s���$)�b�6	���+�b��>�W0�?W)V��'0x�W��i�IP��I���\��X���au=W��<S{u�_��]}O�4Jʸa������o�K��?�o�5qd�Q��}��רL?��)�MSX���?��o<�ML=�j;�����\M �/z�ܲ��������	r�?L�L�����9��Þ�d @��!�I�]dIyV�ah�g9GJ�Ŗu��ĮQhC��	)�qwtE�[ l�w��X����?H���&(n��u��L7|Y��3����V{y�!ܻb�j��
v~	s(��m�|��#���eB�w������{��BsKI�(4��ʾ�^�����B�TY�S�u���ꘕ�Rs���p^[X�����`=Y�.�Y��1�J�7���=}�>��l�����re��Y.���C2�Z�Dh�������y��qj�C��E-���5�&�Ԛe���l��y�z��.'��4�c��R(.�_��K���׵�l���OX����ŉK�P�'r�9�zcAh�����K	�A��#��+̼���E�y�0;^�����o�Vx-x� W﫞�$!�譞t�n����ŒMHO�3og|���!Lv�,&��:��b��m��$�{�ڶ����I����z�`%��v�g:�䆄�٥�Q��L
 ��W���� =�&>zQ�:)�Va�/�s����{���@]�`h直|���M͏|6y��3�kDN�������8@���;ص�D�+��Ҡw��x�@�p#�(���U� �O�v�+����jAƖ��i\ r[�py�N��Z�P��@�*hۯZ:�_�J�FQX�O��Tm��g�'&d���p�#�J�A�+���~�V�_n�5w@��S.�ߐ��sr���Ɍa2�+2��j,�+oH���Y��cGX)ZW������OudO��	]eY�M}Z7F��j,�o�o?t����gv�2�5S��z�eq�r����yX;���U(HF3�1-$�C+sM�a�P��.:0|��|4��p���,�����vV����[�Mx�_U�®�T����p���f��qH�V��6Rp�����~.&W�oj�Q<�޶�-v�e�}���Ӥ? �<ݒ�{�%����L�c�ѡ�*ykm���W��O�3q���zPŝ,����5{�V�%�}���c΢�8~�i�r���Qa9h����s�&��� ˕yj@°��e�-��V�7�K4mq��o�"?�ǥN婩��J`Z�I��b�i%"�f�������@�w:���*�;��ԕ�(��,J�����r�
� ޾���ߔvwF��a���Y��]f����31�G�����I�O���5�.I���g1��_I��_vO�	�΢5�#C���G�
{fUN!�j"�&Fu�5����v�����lHˣ.��q.j�R!q�0�����,����Wo���G�k6m4;�uu�R^C�AgQ��}�S�'�<��_	Mx�<�n��Qi�T1q���.�?��#�L-�2R�ӐCÄ��5�����^v#�͗D�Z�K�Bg�����[���?@s�ѤD}bƮ��.�ݶlA^���2��2>;}/-��/݌��_�lN��^�>qچ�GL-/���}�]H��T9:I����	�3!_��O	��=E�h`&�_g�ڋ�3���D�a����}����N�^����=�Np�ծST��%j4nx
��"(m��#$�V��Ƀ8 g����Z�O����������v���q�\�y>�6�Q!<Y"΃c<j�*r夦�(��54�\��=���m-Xq�#���� h=
YK����	��M�˯�����)�ӟK�+��\EF^ׁJR��V�uj#���$��se��h��Q�`)�K�e�C��ۉ����-�d�OP�Pz}�\��E^���v�tȞ?�������7w�C%�9\����c3����ׇ��>�U'��T)<�
<n�҃N�,�bt�ZRd�_�+���Y�(O9�{�mu��!�n�T̞)�"�e%���8V�;���c��L�wvM��.�K���NyzFăiI���b;;Z@�q^��@���,%o��~�c�� }������:~�,�鐴O�:�%b�F�9�K�N{�Y!.��O�d0N��:V0�x���"MF�l�R�����8������H��m 4�̍T��Z���^�L:��e�ݪ���kó�R�;r�!f����V*Z`T� �ߤf���w:��v�c����J.2*�D���~��胆�O+0�s��z[#N��A��O_X^M؋CV	N�	ם+�؄~+2��{]ê�.lM@ǭ�{d��4��F��]�"����ޛk%c��Z60(pP�v����ˎ��=�.x��X��G��+8%�A��{b7H�K\�@.�&p�)��}���d�&��	�3���_�7QW��MK	)B���M�W���Wo+-�j?�$��|	{�i-��7.�ҥ)��2�9Q�p��U��3x?8k���y������f���������ňY��K��IOcQ���*�z�V+q:Tz��X�=D�!
��,��סPsRz<�*x	;�B�����`GK����Y ����	�ke�-����(
��������OApqu�n�c�#b�#���~��E!$ɠL0��	7J[<\��@q�y<q���HY`��y��[G{�j����1��ը�eD�^���6⽿~�k�m�.~���c� ��Gl$��c�yI���������?�$�UdYf��b�I�tO�!L�@aP��W* ������lt�px��{�ރB��G�׆�r����;�BDUm�i�։4�y���,��TqP�.�td�=�덕��{���?>���@!5��j�n����ڃ΄���3���	}҇@Z����e����mV?�����Q��ZQ��5W�V/�11	g��Iz�Pfc)0�P��`����q�jUL��0�a��)�DV�],��,ݧ�ul�(�sR����K�i ?(���߉��l��\N�ŒȂP�5��B�Jo �C�����*��FU�ӷ��]�g�	q�	��>�@�PM*�"^Ka�Z����=O�g����X�CU��X-�W�N��X�0�'n��?����8��:���@/�̱Ii�J�},(N������j47��08��8��3�
��e�*-űw�f���_��%����j��� �*���̀$h�r�}�)4�%���]��Uч���)��������C2�K�Ňf�B3�����t�O��J�� �VO#�������a�j����%�Q�����IO���$��),�啽�k�
LVͬ��Y��nL�l)�mF������c��"�Y�zu"��f:c�'�4�fy���p��va�mp��3����΋�x��u��r�X�t��������)��S���� ��9v�'����.��!vJRz��x��e�Iw����k�z��h�3���A6�*��ՏM��^��1���<Ŝj�-<G�n����~���̀��D}#u�I�"���]ySxO�d�f�H?�	mt���>�Ƣ����|w9X��IU�ckf�q}25�~�����
H^�������\��-@��o�GcY���"A�/�yl�]��������Cj���D����AZ�k�2���3�J�/�|U��D}�k����H��$4��@��O�ɜݻ�����;���,����L�	7�? R��H�����ʥ,w�tCX���Mc(��N�=Y.5]��,����=�� �&w����
I�%w���8�� v&��@6rB2SV�6#Rt���l��)l�w��#z5��zP+>f���O�r���Ǒ�׸#��U���v�wWiΩ����U� �x�3�?��v��B�:M<����xV:��8���~B��(V�����~�2�;N� ��r��L��qL[�Gg�w��	�F�ƣ(*el�)�夝1���z�(�3CQt�D �5%���d��ς� {+|.H���Tҍ��&gI�pU XU<��>���j���G+F}�D�F#�ztn2?���(�l�7_��Sȅ��q l�J����l�M ʤ��X]S��$u��3�����x�zHrq_#a�`NZ�q�~��`6�����TU!���+�ϣ]�?,wOp�}QY�)��D��)G� ,�:ɖ�t�'K����P���J���N��� %�"}Ѧ?FS?�(�y`N���0�}�Z����)�U�����y^���E�7)coM;Y�{��7P����0���y��n��oG�?(Y��?i���9�z=���M��1�%�%�Ώ�ޅ���q�1�E[A_������+��9��#���`�қ�d�R�-�p2�>w�����BZ�X�s� _xcR�kYac��Gqoeo�Y�`�tu�[����\�P�7���2�F)7�p����7��~��
�f �JS�����yj㨈M"��X��g��S�i�O��b`'Ɛk3�����Ⱦ��$��i)ܗ_{�p���5F!���1���R; ��ݣ�2�vz�����a��� �	oh�G�`z_�k;��Z���<��:����kg������r\�pː���4�m��7�����N�L	ɀ�f�p���GW��|h@�:j���8d����r����;�hT�!P�]_ӬLI=�tk��2�We�����)�ގ<��	�ȅ
j+g5�w��G˙ŰI|��1�1�ҵw��l:@A?�a7a�r�N��-@{<Y6������]J�}9�O�)���
��k|
k�J�I����ܘ�[�eqEfVⱩ��r�O� �b3DG��|\b�R�)'"�1gכ��:��-��F�v�|���B��CXGm�D!>tk�r;�}E5�|=�U`����ٹ��U�
�0�3�G(��(Y���5�W�������U����)�#�f��t�꠴��N�4c���n����f�ފ����b��94y���/��}��^��̲ ��ڻFTyDUTq�����"d����J�Iк0,'~��'�Q4��������'��u�z�r��Sm�*�*�,��=xe�e��!��/'�%H5�����*I�����&d&�/� ߍ��UGm|�|J榯m��)K����� հj���(���KS:��H Y[���.j�]K�������A)���u���%�Y*�ݦX��c�����=��DD�Q�u�)��9����V�=�=iq�M�_jj�D� v� j�)��,�o��-g������&o��f�Y�->\��^���w�x�j�52OC	Q؈���'�)X�W�r6��/�m3�G�r�: |2A¯L�P�"ݜ���h����Wav�o{Z)~0����i	��,�x��$^y73*�YG�./���z����8��?L�����}WH�u��"U+xl
��B%���|;7.�C�	Ơ;"��jL)q��Q�;V*�+kdͿ�@������	�_�0��u=�GW"_�	��^����>��;��4q}�qfjc�b�F���f�͘�7�G�<@��7�>����*���y��(bw���L��(�v`A�)��x�@Rcmb���m��3"
	&ua���L+?D�d�d����Wu~8�NX�C~�Q�)�s�G�tZ�`GD�OL|�m�W"�(���6����31��3V��.����Pa�ܩQa�z���&#�VW������[-W@�}���7g���<��2�\�����n�q�4Wv�XF�2��[���-S���=Mr�q��¶Ȭ��={Vϸ݀9��'I'��|��
@�0 9��Q�C3�XxfT�+n��T���[�2*�)���P�>�AT�:�.��AIsl�(������w�s���=�![�X���u�^�
Kٶ֓�+M�	���*����g���G��A��)?���ie�0��z�~�� ��"d �&FC�8�HkIT	��p����dz�h5���U\{���Y��d��@�Ky����=�����\C��P�"8�P��~7���]OTv�uF��^�GpW��ͩ�[]�G�rmh�sk�ZFS�?|\X3�k��ĝ>I4=޳�Z��ЎF�L̆_Oe%o�Q��7FY�.��JD�DP�^}+� 4{�:�R־��J�AirQ#kd���0ADQ��g�o��M,"��=M���/
Y���hr"�b�ONz=��Hh,��$���J���m�u��`�;�0�G�6���L��vD[����y�ı�I��q��F�l�F��8ob��g��	��'�+�u,��ޖ(!:�?�ծMK<�&zX��ctcb^S4��ëP$�\V��-��]����οA������c��Ɣ0���ȤO��!.xMc�H�a����pCU�-��f�����
M�}4����d��M}�}�r�T87 7C�D]:�H p��3M�=�4�I5|ELy:/�����Y�Q"��z�i�5%�H�������ii������(���ݕ�Ǉ�_�8ݑ4p�����u�WO$F��@�dŞ#�y�L���;�Z5������7e4T�#�$�ԱfBr� j��#�,��U!R�C�M���ͻ��0��59��8�d2�w>r�����ұ�c�1'f���:��wb湎���)�[�2j�} 3�Af>@�ˌ(�	+p����~��f�D�b��$��!E��,�����62�yrG�S�M�UQVP4��y_X�~gXEi�vBqH?+]W��l�NSd5aw���I����k��'���/��Kq��f�Z�4P�}�-S�n��	F��������������?�JX�eZ)	OH�`����g>�u�w�w���B>�A:�	mt�Pq����Y����Ycn���-����ճ�$��z�Ѐ�YGv"Jq�"w��<���<8���"��G`���k����4nS� ��jH"�r���MD#MN1>1�`�ѥ�T��,Y��UW�P2�����1b��#Os��qh�ws��A�7ۡ�C�x���	Z�7�_e�;D}ҎE�D��^+7�wFV�p� ���N@w�Ո�WԃJ�<I��"�MwUH�֮4���
+%/��#D,Ei�J�6���H6ľ��������@���*6<#��p�]���ם�'pv�PId�No��^'��+X'�-��:"E�k������iZ���⍷�\�#8̾�i��M��V�?���ٟl�<��� xX����~��4���	��
�����rہ��� �0��`}M�9y@�����9�U�9�Z�ѕ���1���BPon�W����j�ޕ��H������G}�ݨŰ��?�X-��9\�';��[����4�V�®���Z�(���l��g��Z��{53@ �"�M9��<,&�	 �cd+��.�������m�
L�0@Q`����в�-c>��t�T�Б{�Sَ�/�����@�Ktc1����a������Ԅ��R��:��Y�?�C���V;����Vɹ�=�ߟs��@���P%eI�jA���N5 �0�3�&�K"��� ��z�����j���Z=���3�ǮFf�^iQl�@�ç+W�+��1��f19��f
O6�vK)�d�w�d3��5j�vؓt�?9?�NvL���%���dʙ�8��/��׌"䊙Imu��^��O��9�?@o6��YR���T�WtXm��$\������d;�G34 �{��4F�@8$���h8&� �f�2�d4�a�����W�KLV�@)��09��.,[��cf}�*�#�����d�J_Lk�q�{��O@��}�P�L��p{E#�>a\�@��ݚ��7w��\R����$)�6S�Ƨ�܈��s�_%��z!3���>�A�fC����"-���ޓbiY�c�>�/EC-�发�]�:�܆@��mr&^�$5��Z	`�f�(�a��0p�Ĩ�fM�Ju�K��p"�1��2��6B:@Ɵ*^��}l��!���{��R(ܰڼ�b&{Z���УA8HO;�m��8�NCDZ�"��n�*�@#��΋���������;;mȅ��x/r<(c:�����6�(����ވt��c�!Io��j#�ˎGPp���4TYO+��mihɯc�d�?�d-�c�u�	��ը�'�q�P-�#��;����3�Ulͩ�9�t�&(�pI_9`��92�ե.����kq3�,����;�m۰ړ�$f��Vޯ0���-{��@Z {��u�0�%Pni�/���������W~M�{u����S��t�L�E��,����T�匳��qY��Zz��#�-X��4�IА���0�wj` �>�:'�ǻ��v�_�dx�'w��hO��L�&&���K�'�B��
��Y��g,@�� �e}��C��20r�rxM ��v��p��%����X�gT��FHF�3a~D;\Tu��j�6$�h�Ⱥ���e�)o<l�+�P�ke��!�q�!��LE} 	uV���6��m�K�����-R�~��to���*Q5.>U<a���>��􎠮s�n��Ag�^���3E��(��k��t�+#e����B�軓��#�6��>H	,��w���dC�R��=#&w	�{��L������9��Z��|y���=)�)���K�-���׆��ǋ�^I#~�8�����낰Z��:؋'�7٫G�O���_�s*v^��
�u0�,Hgsr��D_EW�<���Y�u'f�Tsm�����_��_Dqm�3�P
�Ý�ry=��߹�^��ˮ��S���9�M'J3/y/p�~Y\�� ���>(0zCx��z� 7lPL�{�/
��/�����ա^��g�I�
�^�j���i�I�oLO3��7�q���9Ȗ���:�ɥ}�LLV��k�j���𤿔ua[?Y��P	�7��3))+����)ԼZOr����/��@^)qnv5\���U]���S�n�T�(9�D�A�k{5Ϡ6=K�0��}e��2�@�)n�pi:li����6.c�Op(u,nQ�L��ӓ�<:���#I�p\jH'����O.�X*s�d�莢�ʠ BO4�*J� =z�	��s0�mX�oA�(�x6��y���Cja�
@����LuIF����rm�����5�F�\�q1�[�?$�^n�j�;���Ekx~ɿ ^D��)��?��bK�I5���-�l5[Y:�� N�M1 ���, �q*�pðxt�`RH?8�0d`�6G�1~k'�7�~����kǇ����`%��_��w��"�'�/���kR�� ����x��޻쌇�o���L���I*1��_���__�13L$@/���Q��K�ɱ�\��_
�0��[�������g�l,�wp�^�H�] x����e�X�j��f'Z�)nP�.�4�ç�%S�F����c�0�gU�@:rMf����u�7�it}�FŻmRC9ʿ�ވ�}G��ZY�ѓ�fˍ�a�x�X��^!�n!��lo$�4�F��bIv4��D�c����s����D���t�Y|N�;�Fp ju"��h�IDW2�v���:Uq������Y��o2�8������U�_�N+@�� c�v讻6&���fxWHtgr��
�9�4��7�|�C�%�B�0���R�����*�M�E
��$O:����1�=D��6H�{KeI/)�M�o/�%*{f���N|6�k�AR@)���!�`@���5���SD��Cn+F�h���TB���=��B�𯶴v���l0��+��v�B�� ����K�p)G�Qo�_u�s�?�sa�u��Y?��+�/[���e?���ȲXF��<���]û��f3`scm_��범J�1�=��)���f{k����b(8a�<�a�E��]�\�����HV(>E���S�L�Ջ�0��䤡ŶHHQ'XO����C��ٔ�S�D)�,&�G��ʂ#Z Nκϙ�˂���P���z���9��޿ف���s����
9�64�P�Y��Z`Sj7�J�y���v����R���;9� ��\��sc���VT&=؎���p���Z`heJ�+Y�j|ޒdկ��qp��n�]b]�䣂i{�Ų7�c}�Z�X��6����Ij��V��6�,�<� ��+��) 9b���.]��z�P�\�,�[C[/L$d�ψ�	Xv�~�n+Um�y�,A=�W �K�hu'���KiQ7�ګH�Ŏ�<���ZuڊL���n"\ų�����@\���Ɩ��HtG�Vpo��%7ȨXSq
�@��!�SX�lq0t�}`����(��c2�>��(X�.ڂ�.��xyN�GL�`-�:̫>!v@.��R��!��
43����>��#Q)Ä �ѵ��-��?�`;OO�n�:Xq�՜�nmdVך4�^��᷵ٮ�O��%��MT�U݂u�s��F�U�	�%��S�w/%�=�Z�YA�(Ą�O+�`)�g��1�i�2&YU�Ǉò��9�I;bo��g\7vN �ͬqHaf�I��׀�&�A#^�h�J�o���I�3�@��;4g2~�9�KI~7#8��1A��Ǟl^!k�M�Fh��'�	��S�i�>��Ϝ �4�3�O�@i}���:�8(�1'��� +�S7"բKʸ�p�"�O�{����f����T;Y��έ�2q%dQE!\�W�i�����Gd���^�؎��ݻVw����b0'}D�dHE6%��S�XZgM��0�5��DLi0�5�����m":�/PŬ��x��� C��������_����S>��
(�O�%ޑV�\z���Z&ņ8�������Gz��~���K�(���{����(1E}3\b2�w#���JR�����V��V�#q�Q����-�4㨉���6�^t�e��J�ȅ;��e��\뢠}���E����/�j�I%��i����5]�8i��t����r�] h;�φ�|���J�BC��!�E����ݯzq�OÌ�.#S�]��0�#sk)���k$"��p^f��mzQ��_?+2��Av��y�[L��v��;��w�-J��]��E�@HF�]�����n.@̼�UG�������_����ٙt��'��t�9,��ͷ�����=�i��ӡ9�ŵM�sB���:�����ﺍY�J��o�4�����=�(ې��mt��e
����.o��ܿ#�ڍ�	�f	��'�庆J�l
��|pl]��9�a{&5T��t�}!�n�0����$��E��I3�3	���a�|x*�����U�.������?ѡ�2@g
�28üF}sw�a�M�x6, �4u�{ U���$�+�6���|������݉�K�_�S�����h�/fa��iB�G��Hp�� K$$H[��+1G���M�joYI��68;�۸��Q�_�o�Z�L�[�ϷL�n�K�8M7fmH�دh�PP+�R��Wޜc�T0p�*j�$t5�%E�\�xK?8h))�O������m�4��T۸D!!Sʨ`�4��t�;����%˧@VV|3F�&��\�dJ}�Ef�!�?H�'�����@�����ӕ��{k]B�LT��}aJ�^-!��x�<9t�G�Q�XE�x��24 �nf#k͝	��ʦ6�� B��L.����+O�h{���#QS�<P�_b����0����B@L�-q�_�{Ym�W�*.L+[�~_e`q �#L��1���ͷ�D���8B���r��dSU 1-��ݦ�'괅�Wh�H��킫 W�]v��y���K�����񜜅�)6%U���|�khKT��|~m�q���  G�`8�c��!H"��s��j�?�@�J�7��GE����Q.���.U\m��ƫƖ�^fd&Q9�E�~3M�����;�!'�8�d�j����e�	�0߻ _���O����VN�H��=���������¦*\)����OKda����0�9��zP���z��@��X\�p	g�]�$B�h	��p�"J*4�{���v���oS��j�1U/z�*�
6,w�����|��p�hp9�$��:m���l6״/vp����o
���M��I�4��@�����b3d[n�:qzxH�I&�i�yd�PTo�Lt?���(���Ϣ�����->�MQ�t���o��'h��ʿ��g����fԖiLU�pp�h�K���s��u������`&��S]Z�?W떐��?3n����[�=�����)�[(�qB�Q�ʒ$�n_�0�H?I��rE&j�3
�
�h��A�f��?E�!w&׊2��Ǜ{/��-��;k�x��p����,�����k�˞��bڲ U�m��y��5�Țk��%�����S�[�5)k���\vt�r��9Hg<�?-K1�R�s�T��"�~���o;����X�Y�A�G3����"�_+����x�]��b5�[q��ezP�:BH�لDQg&x ��l��W��� (?�����~2]�G���Ƕ;I�z��^~-z�<+{c�z������=N��9�2�4g��(���!0�l`�+P8OTB�۴�pW�ڪ>��m�`	�L�tU���� -��۷^M��=��n��gdF�	�EJA>��ɚtqos1�ci:{7J�+۫��޹��ә�Ö�L�\��i�"`�z�;t����/�щ� �#��x[r�[�oI����T�f�C�h!7<�[�MG���E2_rT�Z�͍ǧ�.x|��Kx��x\���(N)?�ݷ��i	�u*ܱ�R�3��Z���@�?L�P�:����?���������=�'����eH��@��56�S��R��L�����٫��$�Ξ��t9y��V[����F"k��Z����1Rq1�,�Ցh^�'>$W><��앿�Yv�AB��]�*��|nx�T��~$.�9�&��C��N�)�/D�zې��ϛ��cֲ̯�W��?��HLґ�8�!@���m���!6��8x����8�k#��T5ֵPx��$�O�bL��o
��RF��Gwo6�%�]1fsT�@aл�>ͨIh��ʲ}�D�������V{���	tz.^���*;l��;1v֜	���&Wā�=Z9)Z����yz��-��-�Lxy7��$nK���� �'?d���PY���n#���O74�޸͝oM�Cz#��GC�R`����*7�}Y�F0aN�����l���kU����80O�c�P�ߎk2�A _=}��{�h����W$M��#Q4b 	x��r�j���V4�hS���x;N����Hj�$8����j�{F���M��ˆ>e���V�H��V��qt�!ˋ���L��Z!F�vI��p��I�/������u�jw\��4Y��V�`���|��u4α���Di���M�=1P�@n��>�ِt�i�������Hj4�6~F�G"7��#��f�L�UOk��4�1�>�w�I����q�ͤ1�{!��>�W m������JKjяEsOp�
�T8�����82j0��l1���ѝ//�l���x��u�a鷽�d۟��sՅ R�D�N����h�*�'$�XN=q7���<s�h��!Q4�^���a�U,��X�����*���܏:���K�183�b�=��~��%z���T�VQ�B��[�@��$�+�=�D��X6�������|{����O2��>!���Y���
#��=���6}�3���9�<)�XtTx��Ĥ��N�.�5�3I�� 'QZ��-r�D���(��wζ{�i��<1�♚HZ�c�+�r[��l�U�MW6r#��tH����Hג�k:P'��61*�(�o�s[(�$�����"���[(�f��f/�*J�
VW��Ơ�.�I�Y`Kls
��q������y�r���n�à����9�8)db�����AHTx���o؇ǈX)�9�(",�4�SgI��0�L|{�X9�4Ɨ*���: �a-�9������0�pa��0�$�^��`�"���r��e��Pd�y���������L!��y��2j'r�*p�K�T]
)��v.�d�c��G��^;�y(4�]ꛗZ�<E��+��SF���]=�����)-���P�KQ��f��o���s���lS�ce��	���+	$E.�����4�g���^ �b����>��S���H�}$�U0-e��cN��>?�f�qJ�\ |��&��;���w�Hd�A'�2cy0ȗ�DG/���tV�}��eˮ部�I�$#Y��	���\�e��uҡ�Ql{Hf#`$"A�A�͙'A�Q��S��v�G���^o#a)P�wqVbJ&cke>s��na+iN�3��W=b��"�?��W��*�% �k�F��}�����*���{v�4IW������̀���
8$���a�[LެBjd�{0�ՀG�#�Pv}d�\SA�Π��%$L�w�^��JB��v��P&��6�9!9�ݕ�}i���W
�cqa�qz��-R;�<�=�X'K�Y�![5P������Y�V�ъ��g�cg�з��۝f֮���|�ʳA~h�_Dڴ4b�Y*�_�i�_��qn��+G6�%�5��`I|�z�gL߀�	�$�7=���
=)n��IQ4^SM]W�N�� ��������N�����]�}�"h�{_d�����a�ъjpa���j���'�K��g����r�/���+����X����ܗ,�w�Խ��F̱G��&�e��򯍊�,�O1�>�Z�iy�9�.M���5�e�~� �r�$�<B�B7:�"y�fCJ��7�.0:�2fq�f�C?�C��As�9�aE�\
�H�`� 1�.s��c_���X�]���˦ɺ4�z� ������K6�WGHf��P����e��P��{/�����tnz-�4r��C�An�'���~��Q `8���ͭ�tp�^�}�u*����>��e��y��;������A����ֻ=�4!��W�E��G!\ ﶸi l�L�@� �Gߑ?T�yW�G�l"VO����N��J��V4p?�d�ٚ�j��M�ێ�?|,ؐ����o5����򢦃s_�����	�*�S��Y<)7��g'UU�%79c���p�W.�}'-,�}��HJ�j����JW)n��9>�>�v~�1���ȿ9��2��`�+80aـ�����pU��q���u
�Ba	�����-S4Lfe�k�$/%;}��b%VJ���M=����:��cB+8>�"�$�NoH�TI^z&��S�0�x�tX2_��c�'�3���y�ͺ�@XO�8W���?��!��py�e=VYK� �	�]�u����@θ�*���eA�>Z�0�1��'P2�߾�=
�Rkij�w{ȷ����5%����$��'
�����Y�ǳ�)��|�����݌�8#�TH���k�b1�ɏ\�*q>�G���ٷ���&:��W�G�2��"��@s]y�z�6Tw �g�O��RQ��{�m)Oa!��r3P�y�C�~�j*A���kM�I����;kj�jl��{�_ujUg�25�1�����q�s1�Ax|���XS�B�x+G"!�:�+�j�3wc�G{���{���h&�p��ą����:�8�Z�5+��(�Ns�*.�%����x��q�[�m�QQA�HKTQ��r�� -F#/�����x�Te��1_�@L�0�����'J�C�)z ��%v��MJ�5~o1��O��b�26�(�x���0�XQ`����q�K����z�e.6�H�H���V�4�D�>�ᥔ1s���{��\j.��.��?�gb7a�d�`Ծ�5��N���[�.��`�h����V]+vux��