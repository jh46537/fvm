��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $WժAi�.��x�Q�{}�>�JA�����M�S
�-�J��l\��ҀD+�A&"e�X�w˲���g$�IJ�_R�	~fʜ+a�-������J#{U���q`���^D�]�r�G�B��y3�̑��&K�{��"]Ί�C�3)�������1f�)Dba�*��}Ćf��aw�����uncg�w+RK(Q/:�z��O,i�,��+6�����@/W{k����:�^B�a$J_s���	
�0P;��Tu�;������a��r=�SG�����4�c�
�%oYH~��|������Y<�;�K���L��U��6@7�ʦ�{�㗺���S��?��W�k�Q�@4������̏�c�q���!_6�C����,�Єؕ=sͤ-X�UB� ��=�<����<�O����2�u'
����fu�s��>���N34�bV��\�-��$Ho$�j�f�#q+���F��~W��s48��ŇJ��;�r�zz��A3L����.����B�6��+�����J�ns�a][}�k$9��k��Q�0�1r̼$"X�ە�4ym�EG2��h�#i�Y^���Z���" q�����n�\�*�-�e��!�u�s���0��V�_A42r�1�yBV� �#�L���^���T�h��0R��a���4���@e���+��E�Sƅ	�������p������HꢧyȐ����tx곖-,g爪�6O���� ���x�N�� ��] ��F�߾�nYo�M��,�y��/�nI��s$���l��E5Њ@���Y��1�z�4C�W1�c���V�LIi9�_b<פ�VJj�`����e����V�{Ӝ.�e�ߊ%�������SL�bi���ȩ�pF4��|G>�!�,���?�d�&֖�Y���fV��Cr��!���l~�VpA'�2�C��٫U�d ���"+�T���Ï�����1Go�yf���34?��;�� -y��@'=f�4c9gU��鷈xͨ������\�<�޼G~-�
�Y����~��b�[�\�,�lQʪdϙ�"ʝG``+��NV����,BC
YRģ��Ra �P�`Vb�2�>��6�FEv�@�c{�����=*�P�&Tza�41��_�]M$�6�����-�c��j���̍t�g�_ӭX�u��-4`
z��&}٦L�N�;��nw5��=]��4Dg-o��GE�Ԍ!y�������2���.�\��t�z5��:��ܿ�wT`S2������.�y�%@ڨ�A�6u,-`��g-�����:�ﰝ3�
����#�P�rL���c����š��nN�e�2��fr$.�cod\��R,�