��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�;<�T������8�l��s����v]��;�W��@U��9m[��d�����p����毲�F����XɹwRD�ۻ�|=�����-�V���T�Ԅ�AB�3�)T��6P^7$>Ƨ�#���`��z�'U�
�J7c�Z���*�g�U�cF@B"��1K���P�&�?26�҅:�X&l�U��S�]k~y/}��_#�j�|1n�a�B@d����@:0��gl6"'�m"M6 ��k�ܰ�M/ەs���Z�1�YOq�3)���`�{Z�i���]�}�<���'8Ь�Z\^��G��ߦ
�R�g�-LҖ?;+oȿ�B��_'�+\�EX��PxP�k�ݤ� ����q�%����$*��h�r��M{��������W
�	�! ���ܤ�[�G��Pf�tY{��N�\�3s�p� ��Rٶ�2��$��hW���4R�6;[�d�Ƃ7��4���]E H�3� o���Y��|d�p���������*���>��:�6h��/�0:�2k�}}�%�ih/ĜE���Ƥ�͵�M�Ke�>[��%�ɀ�๿ƄN��5���pT�>��B��6�2U%����3�d�EV��h�S�x���}�,A��W�8~�#�X:?#�=홁�$���X�s���"�+�2UX%�RP���>	�\bʡIw�2�7|>^t'�˫w  )��ug���R�����3��i�7#�M�FI����t%Ū�ɸ�7g��+_{+5�x�.���x�N�� ���9���(�g���x}3Q:�gی<���$a(ȨX��ܩ����!�R��asd�2��@��7��m,��U��i��YlZ�Ё���O%��_�A^b-��L��A��@����f�S��nwCv��$PgDQ�S�i��φC��`awl�?U�}L&���=aq���2�����<r���h�K^��KbMpv��jc�}=�H�%D�f�m'vP@���̒��7�za�`A���N��4N�:���ޟa�e�v��$�N٢������x����B=N��!�d�����Z.H8���o���LxU���@���n��dd��P��%�x}�_��SI��	�Y�&Hn)�3n��D�^�"\d����;��&DBm�� p��ز�	�dp�ׁS�o¾cs�3G�zf�mS�51��Lɇަ)�D������#s��Rp����>����ڟ+�e�`�/�[�����*��u�(	��"�������?��]!5L���sb�|��;~��[��x��)z��B��'����O̷�%�}���Zym�j�e��V�5w�������ނ��jI�A����w�ry �v���.��%��t�_�~鵣���(��φe��6�a�S�썾Q�_�tB��X���;�_F��Mݧy%R���w$x�|Yux�R���y�8�u����{Zڟ���܀k���KqC&)���rHg�O�����$�L��}�eh���yE���/Q&_B ��́]��,�6�����E��:�y��2M�f.�t1�
;��X�F9�?c3;zY�vI<�9��|��x����q{���C�r�%�Zg��^���:��=���H\]L��LC�I��"�OZ��a���f�4h�	�[	�@�ik_�	��;Nmj�p��ٻ��/��9�����GQ��?�n�zF#7��W
�����]�D㬘P?�Әgq�O���o�FOO��i[�h����צ����������D��@�,8Z.)Os���9k�;9c�@oAg.�'@��&
?B]��ꅯ� ��o��*(��uR\ ��8,[��*W���r�=��D��,��_��
U�s���c���)��7�B�g��^NOߺ��h}���u�gy[������z��ܭk�|�3�׆���3ߞi��o�䞊 Z���5�4�� ������lSr�X��s	��U�)����֧�v4%ms� p^%y�6�(��ʭ��/@��A��p�N�Z�#Γ��;�O�	Yl�r	}T�r��Z�.�h�;��h������c��裂k�kd�O�۝\q5^`ѫeU�A�O0S}���یRF�(�� ��}��&~͒:k��!|(�,�;S��5:���얹���$����  �
F����>��lߏ�P4�0*T�^$�}4����,י�E_5�H,"!����p�z��<,��F����{
����j�dӐV�)��bHI����9�'k��Yb��cz���0�� ��<����32n�jUu�)��B���x����1��j�rn a���,��>ɸ�����W)�5�y"E�E"LtۆM�CՑ0��sx-���V�˺��$_�5?I�H���X6�m�A�"#J�n�-b;�0��|��ҩM\9��Z�a`~�&r*�@�уm����S�?">�~��I�M�j��ߠ��	����Ǚ�\��,��m��[�'��{�_�ɗ�Ŷ�����e�w<8�${-ht�����ΏGM)�voh ;�Nh+��z�h1O`����Z4k�%&������5r�� ��S�4m���S�ˬI��Yj��4Wވ�5[Y'��5H$��</��;�A	md3�L<�̲����v�����M��<�f.=��V����HCjc�����������=cD�9Cw��
����A�A�2�"���7+!B��pFa���7ș6pʎ��_Z��v:�ȭ#�P,<c@5��R����=��\��Ö��X�ŷ�S]�>�+
~��ZD�.��d����bˀ�L�J�@8�]��_pg.n0R�V������ՉCn*�oj��8�V���d�:R�2�mj8�S�*/:!!�N��23%��������p�-,�m�ALp#j�?�Cϣd�N(("����;j���S�#5�Y}��R>�q���D9]��Pnk��F�d��5��J��i7�}%g���p��d��)חz�P�e :�;�'�:�<���������;cQ )O�}�z�tJ(J�n�#ְ�����j�>�C�������]��͖�j��n8��3���2�33�����6���,pgtXV���e4��z�<z4���4��|�UD�W�BN�
�g�$ڹ˄֪`̅���U�LH{IXj���r��M��C7�?�_L�@]H��,?��N=V�)o� ~��v�I��<B���	<�a"&meLt)c��<Y��.)ո���G֐o ����^jN2�{&��j�@�=�+.u��%����}�<�e���q�҅k=\����hc�~��Ryϸgd�Z5:�ᯎ#��3''�i�E��l���~�ߐ��i����}c�����
�,ٴ�O���;����{M;nsN[� +n�r$9EɅۘ�<G@U2ɪ6(����7��#j�[�X�\�}[2?����e�'�Yk!R����_�ۻ:2U���g��f���(�V��ˏd��h낗J��I5Scs;Vϼ�+}u��	N5�~^s�]u(��Wd'�i����ihX�  �%o�<�R�M��n��1�s�F�&�M׍$ֲ��2�ΎdV��1���ҍ��g�}gl��=oP�Nr�{����9�%\�zb����|���>R$��5y��n$�T��6钴��2y��B�"�38r{x��Ӈ��ŴC��m���V�l��'GK�oyr�Rڃ)~q�ٴ�I���5Y�l�H���+����n�l�>i���4^�BF	��κk���V{lJ	��go&����9�WeƵ�P��\i�j��N����C�4^�8a�
^����3�&���V�\���RQJXAఱK���힦D���XZB� \�}o�ᄻ훼u`^�1l}�	�$k��p����W���r�e1��\�@x%�<�W��:4H[����Dr��J*����'�4^t P��cF�ג%�[��Ay7�y
P��"9O!Z�y�.���y�UbA�=H����O˚������ơ��CrbS�S/-��K8?Rn��B���g��e��{DL�����b��U'�Z'� �R�H}7ʫ"�Ty�|V�Bx:�LB&��E٬0u�)d�ё5<���Ա<�����YBě�l0�b�en}�%A��}���>�V�Q_��T���qɌސ�]�.�� \͡���
i����D"x�(�=t�Z�d��UiU̡ ���F�i2n1�����"#@�ľo��} �y�ܬ���o����4 tB�[l TO��9pNZH4\Z>O�5#��`�JI���:�;~CPQ�6�g�H]�P�T����֣7 +��o&J`������߶-��j@Dۀp������f��T'���ەw�Q��b��5L�`�pT��Q�E�W�d�`nܕ�s�k[�ș�
*�,F??^�`�94���(~�%R,W�y���E@3[���5�/H�-M�1���K�Ư���Cea��Z�<g��s��W�s@���s��8/8�\���$(��߆��l@��g�b�����$=��tF5eS��h� �O/������\e�nHNwX�a,��^Ư���ޒ���.�����!�d�LsA��M���>AN�>�DH��՞���?�����{���\@�I᥉��4Ż�K������`0��2�n�ĕ��b�v���:����<��)�El�!A�����8�Ɍ�oW].���cl�|�j���{JG�䬱��h����h������ăB���AF����L��08��H��]W �J?�BB�V�H�~������Q��M�A���w��B��H��ٟƞ���!��&��;�$���Fp	��Ky�ԸH��+�nW�Cp� d$,����]�����P��{W�ڤ��V�;��0���skg�.����V�M촎WL�[K_���Z��񡨋��ձ�o��\7��kS~�C졹�k5����{89�
B�`&�g���n�uk��a�$����N�п`�ιp��H*GXԻT5�
+I+�'b�͊T<�@�T�[���"Z��!�4���i�˟����'<�����Md냅4�s�a	Q�;���$��OjƢ��-�A�OU��:����E������k~}��!
�S�;�}��X�8�kp�r���yi�j��p�JY�ڟ5��OIE[��z�c�!�4�����+�6��Z#�1&�ί�b7�%|]۫�ٯp�V��X��TX5�|d��OQwqa����S;�j6�ȳ����3��(��R~��[�#N�7H����ʾ���O��I���Yx���(��\�;*X�n�e�f��İ���]a��� ]�f`g�@Fc��S� `��svhS��(����#Rx��w� y���U9r) TSC�_�m��+��]	�Y����9T+EՑЇ��$����|f\j6�l�z�$,��}s�$��Yqr�S��0�%$�'22g诔3�6�+}�.]c�e}s�F�ľN	�n"OMۉ�k��?�6�;?���ހ�l���^S�O�y�8�l
jn*A��L��cA��l�T�H+:}�-��/	�GS4|J5�EP� L���\��=B���<>J��tj@�u���Y����95�<�_pO>���~D�F��I�K##�aCD��T��9D	_������1�+so�dkM��e�qnO��`�E ���gj����5:�2]Ћs��J�a�H�=�iu��Ly��乮�vwA"�خ�^�;%[���U���~b��w)�tiji��~+��&Ν���6��H<�BI	��*9�+�4�S,�fX�?��!��)�:�V�+yW뇈��b.��+��\1��:��v�m$+�8*�Z�[��Ntv�a���MM@g~��H�E�a=����>�8��S}E���s�t����R挹^v�;�'��:G�P���~��E|K���l3� ��E��E�K���?��k�-'�A�!Kn~ce0�+��9d7Ұ}�$�JѮ�	6���1c�^d=MG#�i�R��L���3���S3�Ӊ* �b+�h�.7��/�Yg�P�_M��C���j��6�y*�tb�h>�Z �#f] ���EFE��6��_�[�H�3�O�/���c��|s��Z������v�y��0��.q�PC�215�"t�m��Cs>�ux��4��S���	@�l�����ޥc���m��x�SzmAr*�n	5*m�ޱ>hրX����͝4�鹧g�0o���V 9P���IlK��Abj�hk@�Y�Q��Upu�4�(�sx��aH�uJv�ȶY�ZD>f��a`6N=C���`�:�pԐ)�Y�uyd����vt�#C��/+�(�`\�r��T�	T++�����G+}��&;[�6W�L��6(�#��jJ�?�w��j!��O��=[�o��ނ�!�i�/r,}��q�)y�_�v��ߪ[K�\W4~F��tz@�I��vٷa�O���J6����f�ٿ�������"�'L�;{�W3♡
���KWak�v� s�(���FA`�� �i���#9�YMT�v����Z�;���g��4����x��ey�����潘���rU�c�zM�9��@xe�l�6�CSq�c`�	����e���K]!���Ե.�.��%�GYAp2rY�r����Xv���ؕ-onr��P��