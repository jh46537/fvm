��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�ӿ�J����m�`�ϺT��^���D��$΍�`��ꈤ�ŕ�^�hT�9��<�{@���io�@�����}�Qm �r��*�g��_�U��I�?6�Ip�"�� �!�i�-_)0j�J��`�qr%�܆�(����xt���	�go ]~�(X.PD��e��啌�Lkc>O��ʂ��s��;����;����kEs�L-;��@�O�6���{l�[n�rXM�n�D���Y0�U_K�3�%��(U�B���Bg�+f����3�,oG��J4��;���ُ�ț]V?���W� �C �ĸ���b�3d�h��W��դ̟��U�nN	#�K �[���p[�j6����a V	~<�Փ0_�D���	7g��}7�]�����D���!.�Q���fk�?����'��5�V*��A��-��K%��# �$�'Zӯ����=���{�\7L�k�ڭ3���RA;x�]۱ � f���}��8(Г����h?
Bw�/S���#O.�_GZ$ܮ��o�����X������6o��1?b���{vu=�jI+�fӵ��©���K��܋$�H�K�V��5�H!��n�2X��,��x��*]��o����e�G*�G�&=�[]�
�L \N����c�y#�A��8���B�?�"�\�n�lW���������v�A�k��w��RߵF��{+��- -�0��LԽV�)�)�Z0�l�����Ǌ�9�Z{����)֪��-2F?�z���.j@kR����:�G�M�?*�]����ݥM{�u���w��_��-,��k��_����D�=_�﹌���=9������"�m�u�ep���S����c��5��͆=�^GE&�y��9n_f�}���)P�%N��tg�(1�[�K��`J�4f]�z2��{�O� v����|�������g���ڐw��H�gۿ�����Ǐ�R�n&��Lg��7Kv����Lq�Q�{[�a�y��4��u?e�ZY�qw,�p+ص����h�Ezѩ�'�HW;Ѿ�el9���a�,���<��9�Ӂ5��ȳ�N�Z��SY�W/Z�DL� �f_�M߇�'�ؾ�3QR��Sm�s:�b-�,^��3	�α~�T����ϟ��Q3���n��q!_�)�7J�\i�x��R�@7����ie'��a��[>�%��W�؂j<����\"����M�H�l=Z������4�+�\�����9ak+�
�Qa-�ł� ��z�*hx'#Պ�jZo�s�-Nn2�o�'�aVP�mS)J�Æ�66^ n9n�
��v9��ԛ����N,���H@}.���"�G����=�������砕���+��b�D&Ӯ�}��������Z��ڽ��o�O����ګ��X:�LK���¯u�l�N6v�rM󽋯}�
�aĚ ��d2}c��o0�o2����L�P2?����	�}����ޓ�1��j�z�<����������l��O��ǽ#=	)y�
1>��[l�����o��q���',-��ؼ�'8\����39�r���*E%Y@/�s2�0f�s�~�f~;�23�8��r
��<"k�ȏ�DT��$��_�ף	gM�҂X;_L�c3q�zo$-�ע���"��@Q����
�s�g�A�h
j�҃�WN�~�vBՌ����x�/�n�tec���x;��9)L��"rr�c�S�*c��'u�(m������ �4ik��e�)�I��>g�6��@�[7\�hB�����0HT�YR��A��W֟��.�[}
E>�S�ֵ���燻�)TI^&$����քTi+��V��1[g�hn]�<�P{��j�e����B�zM�� ����~���R���<�uxa
Dz�Ԟ�BZP�:�ӿ1��QКa��C�hN'4Ŕ�Cm�=5/�@C&�=8�|�l��h@/��~Gu���[���s�g�S��8�K��;h��*��׻��@�N(����m2��W�8�з�4]�c�0$Ɇ��e=���]�W�Fq(ν9�������Qݙ#c��f�*�`q�"͑����[�>��&���O�����cC���Baa�F�����r���/i&�׾��i�����.�������m��GRҨUxĴ�!X�G!�$�$à7?���
Y���c]�����K^Gtl-
�o��7R�