��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm����질�95J{۠�`\j��G�!�<�ց���&�l,�y�ʰ��D����&��ejP�4��:�D�BH�v�Y��0�����"J�������W�#0���1�Ay0����+�.��g��z��Peˇ�;.��㝨i`#��3K��o'ͪg4��T>׿?^Ti�j9`��j��#cu�����vJ���J�����|N(�on�@u��w(�������'9����'�(
Lh��*���ù7R!�߹O��l��~J�v�8U{�P�{י�-	�3M�b�s�O����	z\8�L���ĺ9�!y�9�R�$eH��>P���1�?*
2U���W5�҉���<B�vj�dW��j+am �Y�23�]�����;�K��Xl��!��]�(�S��Oe^���%��)=��x��@�@�@�WvF���d�➲��� \���"fK9�'8�}�|C���K�ԃ�u����SO�5j�rSU_?,��Q�����+��7}��}�ofX�{�g��4��؝~�g��v(�+�4K��0)�%X����[qZA�\�{��U/�;C���e��F����+���*t�?�dILY�_߆��w����֎�QEf�{�#9����
BR�q4��vr),�ӈ��_`��Ҁ����G�t�����ًx��*~{��,Lz�S����(�N�'�M"�՘s�uپ�%5��B�*!�*Fm�ư*%4|�b����▁wⶁ�����3$l�od���U�ԁ��B��.�ɬD�Y^�խ4�#��sg���.b�W�Ԅ�? *7.
�I�U�8ڳI~F|��`IN��Ym��X4po|IFڷ<�Z�L4KW��q5�;�;ҋ"#m
q޿���wm�Q����:�,m��NQ��d����/�����m��(~�S9����dX�W��5��uF;������S��e�<�� ���2=��t˺�r�P�~_���/�����!Jm��p}lԎ�~�:���pK������'QUl�DR�y��V=���W�-X�4�i�H���l㪀��;ǆ�#/��/�η�q,5�̓c�5G���~��U��݄��f�#ju�g	\�mR� �@	юQ$m��/}=E�Ha�)Qڒ���u1� �^#��&��H�U	V1�=��sV��^��7�	��a{b��gO�p�;�>��Y�4��&�^f����ܢ*ހ���\�:�_?�v n1��}�@�Hh���۲�\]�\�נ�hN����JM��蔻�(���z���dK�D��q�x��e/e� 5�!��E��j���ޯw,*�N(+�U#�EW�h%�ڦ�`@��a�l;�\�y�����4!b@���\��@h�0�}hጟ����Ρ�! ��a�ЕWM<$��_6b���j|�_�͌N9ך��G����):!��}D�xV���Y��w�3:@���\mM�jw� ��sJ7�B_��ðbf�b�Hvڦ�?��=^�I�%o������z���}Ϋ��,���}�i����I�ϑ��&�P������2,ź���y�>���Z�ǫ�r�xu�m�8LJ�����������f!q_�?�/*��B7�],ŗ�2o|��g��;G<��B'�̵x4��l���'���u��<�'������O����d5,�*�'O������-_FK����H�g� w��.h\Ƨ/�.��4�7d�h�b����旄@�6q�MGQ��;�,�$6�i��uc���&�̄��@p<��	�(R"�;[����'`nA@�H-����v� ��"�$�צ��U��ks��S�Zv���ʳ�`MjrV���bKv�帵$n��W�[��x��B	o���-m
��Fd9(3h����K�Jr�O�����[XWk��]=	y��F?Bg�ݗ"�e��鿋z#��sl�.�sF!*(/�|��N���'{��?�����%�j��3K39.��b����w�[�%�%d)���=īɾ֌!�*1:]mbr_}��'���Z��W}ل�����> Կ��v�d7�^�G�������zgJ�¿��.k�2���Bt .}:4J�o�_���ש�M����>�X+��݌�P����r�i��9P��N���F���#c��|�޳�ܠ�~ܟo� =�W��U����S;��FWB�S�sL���X*�aH{���Z)�<�TF8k��w��5|?=�&;/�^׬� a��A�f���
	�����ܒ͐(���z����(p���#�ϱH-p�e�ǫ����&ƪ�40���n�X�o�}�(faX���Հ��ADT'��n�����E�q6l�/{L����|��	����b��:�� _ܻ<�0��Rde��#��ޒ�K��k� �0��W�z���B�d�TպU�<�R�+"�v�y�e�sޛ�Vjݝ�N��u�\V����L�[٨֕<h`������)XG4'r����}8sܕ�3����2)����̿�5]��Qq�unc�����dH�/�O��3$�l���U%��6�5��"/L=��-��V3�/!�&�^�Ȁ"���M���o	�,��1�P�|ǵ7�<���1v"d�Zқ���kig�l��u�ݜ1�ɶ��N��U�C���~���r�7�N�r�*����0ϕ�u�^Z�ItP۫���]L�ѭ'w���t@�P�e�-��G��:�:&�S��1������|nk2�籟 :AԵ��7���L1[�w�n����������N���=����K��	L�[���!�}`��A'K(
O(`j�#��<x���Й��H�p�2��4�)<}�$�d����)����z� �k"��
���k�sճ~��Qa-qN U�x���o9�4^�!�^O�g�0�}���oZx{��x^��/���W��UG��65�w ��<�ש�Cɍ?�,��8�5��d�����EE�y�b�i�ʈ��]���$���y�oՅ󫐊R�FR��9�<�eb�K*����\�r��.[�=TC�ˋ3[d��1����r��";����O� "��=�u��{������L6@a���O@�������:�� "MҢ��2��z��.���B��:Û�@��{/+'�Z���V3���K{�J�MG�SM;*���a� 	u�FYM|�z#`	E�����-,�B�����!�Tr���U�]R&��8��<�����|謃����s*+M!T�Y᳨uw�y�9#��?�9p�!�5�7�6I��F.�dM�;F���^�*��"&�IG�+Cd�x�'�ߚ����@�)W� �<�����~$�J�d����w���ֳ_ܹN㯰/Ԭ�B�����N�%�uD_���RҮ;�#$y���hRBV'��	�I2�2��̀���A�n���kT"�^����A�Tj����[ٔr���#��V�Ӭ�4R�i��Y��"A?�p ��qjY���+���ɷ?�6|hr�Q��0�洙)޲�~���+F�W4S^#e�l0@!���3���>��������X�M�c���K��H#�)��D��D=^�e YŴo'G᫰��T"Xl�ۋ}E#kQܤ��t�J!�\49��T�6~���T��dqX
�
�3�4�b������~�l,���U�t�a��16��1-��5������@C_�j���:]�O�R����ew�W$���p>��8���/Z�K&�w/`PMnr�a�˳�'��dI��X9k�_'R%�e��e!������*�h�P'.��u�ߦ���D^���{F���ڢk��4g��z�d��8�͐���L(1j���CQ�Ad���\`�P�+3��8���Uv�VL�L��v�����{�z�k�"�݄C��Esx�ʾ`�n�|iY�:��Y�V�H��G��)!:1�v��B!17���HHc��R[#	��W��i���}�G��מ ρ��ir��Jn���V���e�tB#]��G�o���5��n̪Hlu;Ƣ؃��T^o�9R�9��Fe�<��X�G��̓��\+-%Jv6j�f���s�E���4\�<����;�YU+���}1�@3j��Q�mkQt�c�%���*��[rE��@��_ �?��V�+��{�~pg��Yٝ��B����.�5\�j{!���Z͡�>$�/���IWp�[��\�����G ��Ȫ/���q��W�m%<_��;^��.�,��"%�"t�������CEWt+�S����B��4>4AH"���~b�Ɵ'=��kQ��&?��޲�ޒ`i봑K�l~�g�H�䇂�|�!� ��Ƚ����rڟ=�.�M�p�c�>�2kW����K8-�����7 9 �#��f8l��A��R*��?e���m��6�0�S�c��Dڙ�&AI;�h����<� ]�����⁩q��^n��4m�0�f��4b������Y1 ��
v��fO��/p����a�mC����Ϸ��.����|�X�N�b��U'�����Q���a�y8�;L��J�ˀ+ND5��%,"�*�����{�ӳV�ǠQ���Vyw��,w��[�g�I����H�F�H��R461L�f������&/�G��`�B���zi\�jB�!En�m8�-�i
,9;=�:
�/FD�g,a�����NpY���'�F@��G�P<z>c����rFl�v�+�ܢ��[�h]�[LҢ��Ͼ��p���<3�'��]���M�!�K�B�l=���&����MF���!���I���u)6Yv'�z�����B�pi�׼�� �E��Vb�8T�:�'�!�%k�g$6��pv��"������j�a�m������L�G!ѝE�]d W}��o���w��ͮ���e_�|�d�^���eBk��f!#�4����OۢkX�\!�hh��mq���z�!�%�g*3��/�L��[�,�{@��\�_OM�$�B���h�]�UtH�c&&d������9�,�A>����1�8V'@7ð��	9���(p\%��I�h�/F=�AB�<�uU��D�[�������A꡼�ӽΏ�}�]Z2�
����n�ſ�ZѫL3�k�]t}���G��X|��+(��ۏ �����0E�MlТ�el`Z�&P��ۡ_��P7��3>�r����p^ -�h�Q4��� ��SZ�?�u-��qā����*#XZ��svШ'1��ޥʰP1e&�O@EN��D����G���9�@�6�p����c���m���)��R�sJ�����������р�*��[	�!�W�SQ����lc�y�̴�|+��$ߘ �'vN�\ϭ<�-���&��w�j<9�7�={��ʙk���2�guCB��ʡÕc�,53����&��}�#�I+gl�2�t�t���T��;��d�Զ?�Zk����K�Q�:���P4��с럋)�w<z������cK���G�R\s�����R~�RZ��$��(���x+�t0L�,�閸j�+�.�?���σ��Ger���xx�Im6-|��I�~(8�P���r��!��w\�B澠���X��)��/��K�e��6D�u��`�����| ���둑�ĔY��U��ŀ� =(i���Y4��3T0����*	[���TΟ����i�����je��� �|r�*�Y��hi� �>�y��"�2�CH�[�.'g�n�8�n@��B�{�E[��Pn�II*Ex�X�j^��HD<U��u�w�آ���q��9�[�D�n��?�Tp�D�>�^�|�'Qt�Ocʰx+�J�B��i���=?Y�r��E��j�T�~�"�=a!85lJ�#��0LA�V�ԡ]'���l��	�tt��F�P�X(B-sŰ��:��������ݓ\��E륻�$���j�/�u��2oB��u)
x\lC�pα�e�谓�S�o	5�J�W� 
�i���,k�4����Z��.���ʫQ�Ջ,D9����i'�5c/U�o�8~�v����{A��_�Sf��a�u����i�ϵ�\&n�������Dj�x�	F>t�'=�B�<��~��5�x�P�R�(��Nċ3�������ǰr�_���)<u����H��n2s*Ij���3`+��R�L�(��V��޴l�3k�9��P�X�͝�{�[��a�S��
�$��(	=��/i���A�4����J|����,�p	択�3����<c|�������ˍ�A�횳�Aq����c���B�s�aLAr��g�V�c}A���8�%�J0Ӣ����a�5�?�2�\}Aatl���@>����o�p<0�:��h5t�֜��Sϓc��o�%K�F=�-F+��.Úk��kP$���l�VI�`���F������<1�p������Q�r���
���G��@%%�h|�~1��ԫZ�@�DBt2YV7@MΔ�L�����.��*.��<�Zڨ���)�Z�J�a�F��l�t*��"p�"��@��]6��Q�W�q6�Z�~���T�8�@�}�W��"��3W_0r�E��'���Q�-�����<��Cd`�ck%q�l�װ���U?��e%�z�㻺�xA�B��rDRM�{��$�
��Nɼu������p'�E�Ho<͹G�:��8���v-����!KAwB@u�;�W\,���Q~*�e(*t�7litN�o(k%)����M������}�z�'��2���3=3���oA�E�i�fM|�:ƌ��Y�!b5*	���0ռ�bn�'�bR0}ڶjz\H�`̾ ������4��l���-�A�����e$ uH�U�Mz�g��a�����*��u��^������ lw �/� >/ak��Da��I2Cn(�B����pf;ͮ��J��x�[��8�8�������N�%5�I�>�ɦ�X�́~��N�m�i�-�[�.�P�9Żr0<C����W�32��ԗE
p�7�.���F�).�.2.R���ę �Ys/����Ƨ�;In[2�U;0Qu��k�YF���Sj�$����S�Ɋ�&�Գc����2�4#Sˇ �k[��p�o�b_i�R����x��{�8h>A`ER�W���&vh�S��b-��C�lw�	 J�$c���h�$� �W� ��)8����@����1�kD�Mc��gTQw)r%���=�9!�� `f���� �