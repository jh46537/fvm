��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�Nf����>qXQ�J�y�� �&��};��_�g���	�߃�:������p�x}ן7j�0x�	�wD��ފ�t��0�A����]dP���D�����8����Ֆ���K�w�<��R�q�2h�����'�� ���j|ئ q���4A�jq����<XV�0�rpƀ�)�UnT�Y(`�WN��!�o�H7zC#	��i������0&��v<L���MhBO^����&|�"Q\sn�uX��EN"�����f����9Ew�?ֶ�h5�t�kn[�ݝ2�Bn�8䋮dn�zuL�[�JB����Y#���3<��23�+�]�y
9����uw'��zr[�Q:.K���kRiS3�FP�'qc��?<?\��
���ȥ����E��(��U��<�40i�=���QPMcG��fO��O���������?8Y~�WPbWL� �MkM���6��\�'��u�_����ݠ���A����\�/O�C�2z�},b��l�ם,��I.m#Dι<\�-E�>�޿3�|>�F�J�Gv4�㱺T.�e�|q"u��9��{G���V�~��՞@Z�������@rK|g�~вȄVcۥ�v�h{�
�hL�n�B7���Pz7���̛�	S������L�,��ve��[}𱭊���y�g�<7�0��ƻ|\(MJ1��uG2L�:π<$ DdG�r��f�0��4�!��oe�J8�i4���BbL����D��K+)t�ĖT�7XhJ��bL�s�es�a��$6�R�By縀�%Ƴ������Фd�MuAaiǏF��YnL��a�㛏���w�1O�f��@��ں��ƌ��?L�6��1�=��i�x%0�E*�&^C�!�dV��å�DqtBCz���f�4��D�p��X�+�-t.oM�f�)�a��J�8A'9=��Nh�R;�D2�M:h[�碆n���5�zÁIU6�Ӣ`)*os��g3�|�xL�t�I*{�]W��#���ռq1�s�����	��� $j����b8�y&���Ι�����i�i���9�k �K=�S�YT�e�6B$��G�y3�d�N�h�8��*���f�;;%GzQ�WvÇ���=�z֐!�R�@b˹T�CX2�H]M�w�����6B��"��T	$_,����U2u��l~�tT���&jR�{�4Ά������8��#&z"�����,�P��`4'�,��}��Mc,5�(-��Dz��Gx٧�W��G	��0�,�/��S����	ܛ��"�D8�vG3�B�Ҳ91.Ȋ�0��0S�^�ka���� r�}���?1לkO� ����%i9�66���@槍P5�D� ����T�1/��ǡ��߼,УK,L.����%�'�[�9�����]��eܢ�i����l�t��5{}!��7n׎��YHa���`.X���C�}J�$��f�e��j`��}k��7s�X����]f�:��8��p q����u�9�H��D�/��y?+2��oz��H���A�5h,��'�����E��b+�]qպ�g��9�3��D6���<����6K��N�A�O��]J^��O0D��D����w�	��q�����B�yZ�!�@���=�_�dǟ�1%�^`�HoI�hե-��Zf�kВ����8�����⣚>:�*�8a�,��}In�腰�n���0^�
!0��_���K9�glpTD���$*ןL `�m��e��)�0x���P��<�Ɩ��]�C�%ї��c>uڜKO9�D���h�_ɰ���j�W����nW������@��Z�D_�e�ұ�xjN��mv4�(]A��o�;�P�]y�͖P&a��2ܣ�\��\k�i�Ldu��T��t;�.^L'�:�Oo����_����(�F6B��xE�@~Ӑo=�hu�60L�u�?��#E޽�N�L�=�;�r�7b�^$I�&� ;ո��s���B�k�;֞TDuY�Z]K���`�ƒPoF�c�~�ؗKۼ���v~ڹM+Ϝ��89��I�����䊒�4��5ݵ:����j���3��^���՝E�d6P����#μ]P�V5j��(�h�� ��W�: ��W���Fx����)T{�k� gx {'� �vh�;�華�����c