// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:43:21 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VupX5ZMpJ3aBQ7Hr890g7defBMXTqrJkinDN5iSNZAiuSCpBLNmRLOUwS+ln97eS
hJc7Rcoe71K2jLpu+7vtaEw90MHhRob9zXH64djpVnkw7QJuskpRvCTb4D2cod/p
klmNT1AWdQ8/BZrQ5vgLNVbSyiufAqCnE0HPqCliwuc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 35520)
ZIgZDIyOhV1N9pZ4AKBmxMNMDr1hPI9lY7ZZ5Nx8vQvUeHfDbCHLLBpCvzUzVGZl
RSIYcIAyTSmVfQNjTRIUhc4OBcCz+T9vk39emxyZZC7Ef67SxNfJSPpscFnL2Xr8
tLtSc5n161njSiTv1JDvW52XP7ADfuSJVJizjwT4A0UhYe3cvSWJDfLX6QGcIi/R
o02jCbFZJVL0wcw4i67ZcUNQ/HyDU50q/QalhjrMHYSOk5WrP6aShF8zVY1VXNE+
8cJ9JtuYRejx7f00m8JC3G6IGtdRgov5ImVg64BH+K20/PscFpmqyas1l6eF0p/p
XQ04QQueJXfngtWjCj5+MppYn+6qmttTNk6KXhuH0o8y6RU6Mha90YPQ6M3UQsSA
IjdfXDDzTN7enUA7OKSpTsCN9Tqbv+v3P9FpVEG6W6Z1B1tf38lBHx6VgSNdFg9K
9iaLfulconvIa1M/Jl6nvtwdTuSVyj28s1WHDSi1ZFMj9FPabkCBRAQ3Cc/yB1fK
uOnF50vOAvgfR6BHKXac52zIIc2Mv1CxPbn/Ftaqjzp2r7w4fjD7/p2DMTRzjWxi
AtIs7CR5w7G5pTp34Tfue59wA8V9onQeZF5EBa/Nwfsr8ew+mQz2yGj4eCH/C3vy
S5A8YPovhVGtkr1ip1TdHOX0oHNBq+7BP6Ue2Obj2n5VwXg21jXrSTRzeJOjibl7
FPrkvXXMyF/6v+L/u4pWnqJDFwAC5AZ6GjNcO310n91BvrUZsPHIl4LYEKzDprfc
Z3W1dFqg5uHHhbL2nnKJAg4vuqbSySbl6MKM0ZPoRLGVRsaRGQEilXEYXe0MI66t
EM7J9m0rbDXF8Ci4hXeAmf/LAG9qOXIkGwVWRM8nB6ZkbSd4g4zq7znNyWxFBrWN
M68+SPxQD5/O2uxWoBG1toYxz3bvF87+DD65d16E2DBbFrNq9/ExoWwoPlbCtRav
3Y3MzEeYb/bjCXLy6Bkm6gJzj6NihqUNNp2CQXpSo3kWtf9j5NMh0FVCrh7eB5Bs
zVFySSS67RGg7WsC4RjeJHfUBbd/S3oJivr94Jp+4unqpUCMc901tqii8HPb7fKk
mplhHgEksn55p0T99HbbA3uFxWxKoUvTPLiHvf2LLHaz6pmlliC4jUYG1qT9KUnG
imNg30Ed/mo6OMYiNrgpz8nlA72vgtAx3XgDQjot775pyiPnaNcu/fLAOPVaXPVV
Ex8amNHXdOD1k6/3A7AX9yV186XFiATC5pYFPaFZpmMgrgBeDRPVZPyo9xMs2nsK
UQmZhZZLywSsYqHGsjBFh5FTrx154ETSeWKs5NTj32XOuq7eDhr9z9a3nkLuwMdY
wFwP1I1gdA7jlLJeyQ2uUPFND6LKQSmzU3CtwwragjT89GOyO/rgRXhCzqYHlCQr
O0AmlkcdYg+NFa9ksiM8dyTfji87Ig2jV2SN6g+70hH7GC2brKwJzMa8/46W29bZ
GZes6/IWoJfviePzs4BQw15UBz5S2hdruG8+8j0Q0Gjuz8SvrJBhh77XLiOapUhe
/MsuDdW/R7d5xAIhBOXQ2WiKK7LhCFrdafRpU/nDzGB5fSBfW/ebtdAkuWniY1+m
Rrv5ed8k2zRp0mbDyiwe9sFsasurnLny121lbcLYhkgv8Lyz+XIE7jDDjWiTsA62
DcfHRpODdWmmgiP2+844n1gJ/7TFD17hh3Dz9unjDpSycy9bKx6kFm8z3BZ5Bdpl
7lrLgDAZNjlko1pAiHeZ/bD2YwkCZkPVbMxTeo+p/klejVn2xOXLrISpAR11i3nj
f2+5S5z/7g26b8ie0w6I10/b1sqFbJx+ZvQMV1i8gBTmSX8wU7FZypKqlA43UCox
t1WPIqWzIfDzSN7D+GuO5URzT6pqp6+rxmDRVc+7yuxf9nqd8JyU8ikq/+GbAgE7
6bu0l4Z2TrBJ+SZZTTR31TdfH4t5D4CIBZEFlKpcLbJykBiXX74oPcXoh1hTN7cd
cL523VCl3WLzaL9LlXgc+ckieaKMaTaARPiBD1fgjEwKQWwh4niEzHJyI4+fxhcK
U5mUq7WmK5iOGZioPxmB8Xh2PRZ/cEh45LgqTucNSPcWCPppbMiQ4GZrS4OjRZDc
1G7HVJcqhzD7wxf77itVwmlyc3DGaHyOGPd1+pEOfV61SKJID3khTM8UOMi+lj8A
ZNoLSqLrDPznOvD/mg+c7A7sXX6StJFdMme+nW44cg4b+M/wttdvUCbXAcfEGCZG
aICeeT7xmtnLxglXPweEK7/TyzjHZJ1LjNiBt5q/GRxhoL7fsVTPvNxatkIP2vga
cnOkaYujPIHnBbpBG/HWIkgCJcARsJVS99ikY3Ac0E6J3JBPzPmZnTMk2rO5p7RJ
qtw0oJgy2ljOA/cdx8WPGI1ZNmluxd4JD7RXXIjFYuqioSVXmTFOCU5W/dX3pHQR
2wKyWS0RJ7qgVaBrFDoV7cbU/WyNm93F0S/ofNQstf2miPWj6r4u9Pq01U+XKgJe
HWQO7bwVfYmoi9fCMCD2iDFy6LZ0fST8XQUJTvTgMcOacK2ivO8BpOMdavpU6RP/
gDrgaPun2BOmfUv03eSPSPx6ou9a5FpG0Jj2xYJjnVCMWysgkVgbGF0sEvbpduJc
l7E+zISGSj2/WJoA4RDaqfldbwW1GQPxZ7q/Gc9LzQ2v9Ka9PzQ+NibsqbWrcNXx
21OHln29tFU1rDaYAFQCv1D8akgktVH5X8Bp/mNFJmdLqEx00iA9Ikoqe4vL3JVH
QcfFY7C/I6Rb1gjumQYyZi6AzxSqonOsejwKX8wrJ66htjVQZFaRj9XPERI+v9ul
TfIMWcDlCxnLw9UgglzD/SzKvZUexU5YlvUJAbQINScn4gqZb6gDF9ABr7whnshC
e8GtJWuUa79yO0H0I2p/dHR3z51Y+T2/teRYHwbfqBhyWl0FDBSCYzpziKWZ0O+v
fM4VCUPoFuaXryxOSNIh1xDLKSpqIywoDDEEQ+LYeJCUwKbISqovbPnh584NJlk0
NY34oPK7BwSmf+DVvjpcRLx+CMLYtxpN2gu7sGH0uvuEnI7fwwzdRLkWfi0O2u4I
HlRyO5v0PrxxhpnITCJhZufpxHfRVs9GBQZl+IfnwOphlyH703canTS4eHbJsSd9
3a89SROwXl+uPNKA54KnKWu1VXNKAo6JluvbbbmxSx5iXxvUN6ivBwO/BYX5Kwpy
JX+8ZdZjReed1sPlpYoRHxpDSO14BuWGEJnfkJ1EU6yX9s3/7haE5KA0lXhgNBsK
T2Qyvd5xxfsX1cwk1PllIfXTvza959SmD0r8AsIt1/mJ2k7CgKyMInNr1r7+fac6
TSdKAF0+SGH+zQWK6qT8Ln1S9COOeayqtfqVyQHSCQnhfIk/VBLlPwAG3QI8b4FY
1ZC2TISd2vRR8POJWZyxYqDhk6/T6PbiSsJ1U93MPpWJQqGcYUUnrK3e5gdDlkIp
1n+qqrg1hjF8Fh6XPs4g+yifiUzrpjWnNlrFRGpIp2P2rFMTt00vyIfBRV5stBYD
Q9RbKc/MKrFQiXs7HZKI6fdz7U0zbjvtItlZTD8FI9/rhkGS+q15VWhv/tGxO+Pg
Ugbr9z9Z+++gXKgp9pTWo2KREjdCGold2sU6EMCkNjlM67Ub31v9/sRGvijJ41jI
cYeaNrT4Yp14ryFlof/iG5R80LbVMeTuXOPnSTKJ/lYpid+4MLpBiPvzXWIPI07i
3pdl5gRe+HIBbUOhMexBAILgs43GmyYdPKNiEokHAY6QGGFTX05HYJFakZpwHKF/
pqX3rStrO9DcvLGgU2S8Z3fF2uarsbXac+9YDNFjCT7YcCFoVA6ZARiFZ898H3VV
kqi+tUpcvCmE2hGJyYsQVYltQjDDMC4kpd4CIIw8FTwZh2gvmht4m4Peae/WlbmM
SqVINQ/PM/y0ME+IjHmHzyqJz6Nuke8jn0ipZccxW4n33ilaGO6yBZMDWOWvxQgp
og1qzPVXPgDJMdkCqqoiWKokqXVwkdgl6iXDJRYkyFeB9kPklri18XWe/XyfqUOH
CRnVnsYe7AzWN8nrhVkQO0dZ9X9WZH6AhqhdELseOnUlyT+X1JuDxL0/K39bpJnV
yeUG/ZDiHiupBEERtN25ongT3o8AdBDVNlqhNJ+/btMxmwyFeFhkpRkydT8HDbzx
kVkPuUfphHHAkZKIF6fuxoyaoMyA59Uq9VUiXC2Hbkz/Viv/INc2aJheoS6XdXSB
bck9caWOD24fU/MrQShPLcHEStBXAp8qBBu8DNywgm7aDv0dmgqwpxHw0L57Z4JI
JgCPUKDH6/tQTTzLq1grBrTL9ereYkRWH8bakpYOmT8GtCMM/ByJX6fAuZpSHhtF
FayZyXyLbWe6yguBeiF3anJcVIQwzcnY90CItyJu0wsCkw7fOIAhNgu92E60PqUo
OTaN9/fZmVBfaGNfXWLQBWuToENdA/s1RPAUkrTJrKXqxMDGYqTRqjQdxZ8iaPvf
oJZ75MMwbqWniYAaoJtkrAPmznGuy2OmwF6uiL6sNAlJVTTjUiKJyqtDjInRbSX6
+B6OfxHQajXeC1d6Xi4ZLUQhNl/9dNtz93p215Qw6CpAKd443bJ5e/ujAlwGUWnX
xlJzrGDkC49A6V/R7REfS1ZW1Gb4TRO7gMfyxin4nOgbEDXZ0oISm4JGcvy0Lokk
d8wOtITXVtDcFjQnOQY2Zd/q0xzQ+SlMR/t5NToZLiv/4nicMDeZlM9+ovBLM3nk
t1qw1UYCtZ6Wp2vC3cRV0W1sFzslxdGy6+Bl/LhAvEL3GXE22FQ8juGOaJd4GIg0
3L/QcOLw1gacudKWWT4QzVJ6cf2yheamw6tddEy+HtPkZtTXYYV/ut6TE3Wehoo3
UG4P88pZ2BE4DzMkVM17eYDq/m4pnQEd4hhe6Tvm13IsyunsTnRwl5RQ5DBA30fU
R3eKRaj36NwBdod6i4kCB3wyHySE75u+4sdIDaGFP5q6Qdsw+JUiR5Rtqiik6PSJ
1B9rhYg4cOn1kjSbVk20RuYvu3Xz4L0Bboc0DauwJG1XIgudJpdB5X2jfpXesKqc
soFo3rQel/62Wrr3OxykB1xf4CxsIqXbSvSAmjuru5lbuIOZkWiqtCgBKCiSK95j
BZV187+WahRjTxf9DDE/9TrYLOSHOOuGJXA7n3x3O1jw2mibcVxjXHK7W/jOEsrS
WFh4mYh/vdlBdkAlWvtFZ9u1TDS0A4ZBFB8SNAOC8qkvzx1WNqdBDa4buShKu0Np
kZ5rrldWf5BAkqt11GeR4CA0dqd7cIbzQgcJbb0oc4oUk/PEKfuFgne/jFdII9LF
Q5yIEKOX4g+cEbGd/DhzE9p4x6mcTi2JXOGRuCQEGViPzd8a7K9nx2vjVjGlsfzq
TERVkizyawdSJPqH+xONqld7guGIufqlZYoKzFuEuefiZlffJhJ4KQePqZUG/g//
0M3a7MZ6lnaZUMgSfJG0fsWrAjy0Er9BDqymfcP1WEw5KCqAfRyzH81+BsESEURE
un0cmApB/ul2y/BGbnJqxMNxmnDTVHPDvtABIHUMxrBpRGM40TiXiSK5AdB3Fmfz
gFf7Nm/1QSGFtHXQ+AQtnYXNSjPRUbY3s+qj2O1kglDfyglPVzaLRS7plmD+SP/r
A5S5FVjloFKuWx45OI9hRkL71rcPIGlM7gau1zevUdnbrHw/Y5ReU1ItcUg0Kwno
KW08UXk7aU/G5aY+ps8SUNtEjXlMUDDNbFR6sEYAj+fSUtulGy3XgGcoi7BCixCj
3MCqg78Co0Ub0qzOn0XX9Hl3iIAzBzE+dccuePq4CVM0LvAjVsnJqk8OJN8MUta5
TwZ0oJRprEfMHpUg916mpl/DSmc9YFaijyzNHbx/Xm13HiMjJS23iOACMJ8QPCqd
gBHx/HIdN9lhBsDMGvK7wvVD1JXFYL4NylfLrLIxhJuPIvLIm2pBoSy/Lirap0mL
3c9Yd6rT7kuVIWzUX70D3tOVgFnD0j2HJe0+gihMIdfC97VALmVBMlenw061nxyP
K/SMsHMAnsbng6uTmqPPuJ0ZO8qOu50eMpQkqa4btN2lTKpSg+DSGhQdm5KYvUOl
7GrbvNW6QVHVvgKvbGEpsQ00E8KuB8ftgHOzfbcc3dXo8pwSuDLDdtmrqi0+xxvO
KY9UFb5c2bouQjXRbHY9GNcr7PESv8qEO2QIDftCPupdLkeYEXdGbUofwYd4458P
hzTGfhygJ48qhUZeQzXe/rYErQFSlDCei9jJH2eT2ZNmufZSo1QaQIe3wNJ0Y8kN
ASy/oc+VKxgH89VpbnzEs763mhW9xB+he0xcE3WpphbWAuySdndrikRjNFo3X2ut
hP43acJBr+NHBc4PgdZko8t6gIq/hHSLsLIgp1sSIOhxupUtQq196a6mIglIsBcr
rIpA2jQJInm48av5frxVSB+qyPUQpl8YnL93dmXHgFPROqy43HA5HHfC8EZUSxzG
WM3x+IDNSgEUAO/q+S10vtn7WJ7AhEZSDmBaSJnxNiNDqV4qF6pBhYHnmUfrbsFJ
F5zibMqtkWdkWqMPxPhTUMZkNiKgx7oEmyxXTgH2A5mSJQdq8tnc5jIa5yBi75Y8
t6fV2uw7/40XHUa7ECMeRqzP8DHJMC9Fvax3FG2ZK/RU4Ls2w95v7n+r7LJ6r/h+
uE7luVtDHyix9Vp5DnvANgkKaqxJTt33/9pTpjn/1F+GISrOiMoufrO3zbeTRaTD
j5Y0NU4R+RdIC58wzVB0Rg54v7swHTjqCphEp9KtT12LHFl2kP3Y9frCE+t9hBbh
P+eGZ0Vj0A8Xy2aumhEpMRBUn80jvvuVYM3tFX+6WBtQCK6aIBubON1S/PweoVUm
pSsBmhcdxFGJ8Fi+fuSYMuvRoYyH4ghEkcXBnhy7ut8QJDt1DGTDNTiLvF21HJyB
l3ieypArI5fp4ws34a1hyNtspb/qAokyrBffu/MbWozgzI5/C0m5TMj3CNXuK4d0
exdO9QnhNBJtjF8dsZoWpYLZjyIwIt253iWFDnyqzjhYPQiaEwgE6+yh5wylWJq/
hhobmbuyX4P+PqM/XajOXjMw7Mr2EjiVccIp85XqjywUGycJd2ct+mY7lt/FEkoe
fbU92tdGj1XZqw6lH2lKDin1jRc/ICPojJ0lqz/9ITO+Iz+nqg+lhobhNplh3FYz
dRx7QXnugglZWWkwxEjmtaoZsPsrxZN5vksqKKkL5DO/JhSbekVEPwA3cm/WazP4
/5uev0ZJVI0lzGPxMYEoLc9pONar0Vvl3ATDYi5IXSn+FIV9VMEGbX8DqFD/QPvt
ZCxQd8xiz6WNI9A62zoAAcXo9D3NrpoNrygRWvXXbSkvumyeCFQpuSjk3UaHaIip
J8QYk8TzTSPszFVlO5mmKnEiMYcY4JiAfdEaCofce+iWl4bYEEH7rcndocS4n7xN
/BQwV1l+Ma2TEIbID6eT+GjUN5K642mSAp5JAU/HQwsBCMuUDqOQQrSK7FDihK+4
UQ5doAiDX0fJzNkOdWLGCRL82D5dp3cqC1coboNU5ZzhkH5CkykYMk9dMAqJS3Hf
pSuSprAUBvwpRQmHXWV2lkEwrDZPD54zRrC8MRrV6kTQdPe3S180ZDjaq5Y8v5O2
E7IpPSefwdhr3d+pk+KC9/a2UBfPmgU76Hj96DDLS/eUXA24aYYZdrfomEsOvJAn
46VSj9HkvHgFfKRKc5g6YmsnrVBo4VLVCfytr15iqZRNI+7pVXBN74mRfY79zOpZ
LC78KKTwbOGRTl58qyvFhUTYvCrcf5RhTBQGiwJW5dpsi8JoWc5LH46xjDM7IkgB
mxhUhKiBKVBsdgJE+DVgVljFXW+C9gtBVrSr/tpnj1IazxQs0nWdL472ieZlKzxA
Oq8bNmZn/isiAxXZeX02sxLwCSv7FBhjnFhaxL7SFdGzLz+0DQmj3QieZWPJc6LQ
anGSMAKhy/1pA2r2gx1vHKJeGnJYb3hAUWw0p4puAFyj4j3GJaKFYM9ZvfIF9N4C
rPz18RrGcf9MyZTCNx5ZMdP6wxAFKl2NY2kploI29LzuLybt9Kw+l3ov4cleTapO
z5um6OAz7acnLtUiJ4ArM+ZPFy7RR8Y3PkaGigkgc+PLsVYZSTuDiy3KE1mktNHh
uTmjDb7RTok3m9GLK+xRBvysQ23OL5vMKHptAwA8ZVZKaRCOdVuG8+uJtnI8H9cf
ocFJjvDx+YnrE0g/fktMPbZUkR0ZTTkpK6iV49ACuqQJ8alOUkZEHVk/it1yur9K
rNMC+BV7tMatsUmx4laCTSrkug/NXX6W1B9x7NZbZ7ZSah0V0pHLsI23OauyC/+p
qqRyD0F+6LTwgbR0/DVGgh6yg6Fnd/d83i5jpbhX3aohb+qfqJKw7kpOw2nWegZm
olKQf+orqRzVy+2ylfHsUtLz7B2hd21czmO1XCnZYUkO49z75dK/jydQnPLePrmg
4l94uXH4oRCFawyASnqdE7lfcBVWu/cESFix6dA9WafJwqxvkGrdmIAJ63q6AYt0
xzzln0uPc4IEuzUVfLj73jyfnDKYsl67sZ71OkbKeK9SXj93CpZf0AFvdcKVoMW5
SMv0S/rNso/2GUI966fSnRAa8OtX9OYJaZHfEZ5ZAgr+4ZoaPDdss2GlM1bUDJnl
yEDQAj14txVY2ITVMxtlqA86d2Mr8Lg7oStfhrkB9ligS+e8El31BpPvDJigLSSV
uyIEKrBdyu1IR9n2nGTCfWZd2TGTk/jI/+bwqIdkgxBX5JWAiirbNcLU/bJ9P8mI
g7965KrJcYB2O6e03KvYMH1mRzIkPLwvHOOOOMbY9IhHYehwsTlXi2H1b+29XmyF
+IWYHfidNvWGBBuFZpYbMTMFc33wY3FV14mlROuIyKN9hq/zS7kQy/7ZOD+pJgdl
f5aJOUju9KngvVKarsGVwdhZQznblZw7AiR6vUV/VoQ3Vdwe5o2+XJLpZaOdY+lL
Blm4RIyZEh13UbHu6Oy5ltkGDMxZml6i/TiJbOfIk2QRmYvGxG+9VdaTlhcE1Wrv
uOm957ZRZ4P+Wxo2Sy1ZQttnqlwTzlZT92YgFlKeffrZE1oW8yRVN3JLbDg8FflC
DniNd3q4tVzRX6VJI2ZG2LB6Wlyj366cZ0F77362GHn0Qqyw1uka0TqUxgwfF0CV
V7mnW84JjiNL2l4FDEfHI+ceg+IDKLNjziyQOI6cqwfTxakK83hfw9XZydb6d85d
1MR4yV6Q4XgBQJuAVR6brABcgwjp3eEn5vSvmqzx+Mv8/a187wxqsntJB4TD6IsT
3Jdfn6v4XxJDxch6A8w6f5Lxbx36YIrg0hTIYN5KNjqp8H9xZO+RLcUMwNiFesYH
YJvajCpx8sO+NcqqQOF6xkUOQQzIXOlTnWOIWSHpEkLrHht9fcYUvntvy2mtQni9
7TcUDkyRg6AwwlhlkhpSOU5CmyzO8J0FSfLcqOh2+lHVaUd0UCUPcUkppPv2wtVJ
28M+WKOZ0blDUqSLet2gZFN4aN/IBqzAsoWBc44XLBCnBFs5XxZWxFhCd//KGC3B
9Ex4+0TzB+iDbi2LVCOzvLMa//vMSzewJKnXFw9DE3mH6ZCG0C0Vi1nXRfrTtqlv
VnpHXA986twpJbSYw2ormy7yN/BQihC97+KvGkkLWNqWRippYpRZ5s4QSSZZGKe6
vpNb+u9D8DhHb4Q/lCZUMJtzPdLrAVbonpSqzjQijkBpMwGzet3255BviHlXRuC+
41DnjnGD+puXQaS70IzcPaBqCY+SRZsS6vxL/i0GKTMiFfQlPWsuVwyXx9qhQSpJ
Y2F3MiQYkV6pjiyhtYE6Ot6cmHN2hg/0tLYnF1d1WUoxr3kYkoK7FJd8IDFTKcNb
oCOcLzHMEjZnWPN5Os1to42YcShbTs8B4KJ3ydKFlBQmzLi3NzD0Q41PZKhx0WQO
HRkNNXqVJuZEYxIOwsRIEWq/1iEFk2xba8gSBER5rhzaSjqPLSCQj4z2Bj+Eo+V/
8d9/YdAt2zlTHNEZWfPr6GHppxNipeqovDB6KURPTfV3JiRB471lt3tt2ZioOpDw
dRnFUvsHHc6lawCUiKacrpcnSABnmHh8L7ShPJiTZpYijo/JdyRai14BekB3pL/3
TSvNmHK1D2cMIq2WNz8qJ6NPoEpQ9moK8TqEZd9U22gJym5PX7RfuudZH6IB7Bv8
r+BjBApRsOcHhP7aR0CzISWE4ZiPgOCkSzQoEzo5Sx3MTljrW1n3aQn4Z2yE7497
SG1ZD4I+lS7D+lnsLppyOwH/rKGqmuZYz0+1133+TxlWqRNf/XgY2JT9vjuB+M+o
vX4e8SMdG+Eosn/faZtHkQj3XQ1VuknCdlo4t9je1c+Rkc1zWrTrsfSHyB8kArKt
YeYBFrHn8gQ2hK3lzIp99YzmsRL/fmWIlnj3jVuTnKBfP0P5BdoEFy5PVQXkW/JO
S+yC7KyKJ2nnUh4d1c4y25/DfQ1Pp+3t+T0TpbWwpDMSuFPd76BdO0O+ZzDAadyk
BKD2HrwpHO054mJ+QnVoHNSSnBKML9kMFi4mR1rygu29zubA7AllKmt6PgN6pQ3r
QNlics3jyiCVUf/sznDrtlLv2Yh87JE1Km5w4TpqrZ1XdCST3ETEAQqnXNzfF9I8
l6z19oPTLF7wR/FtYws1OidK0bqBYnBrWTtYpiqo3AjiHwvm8D57x5DfELoLZo6S
o3FxAsX/boONoLU1OuNp37lXVAyKi9FgM/VXYB62NPHMLFu+PJAlRIgDDGyw+wGy
j21oYXtvsVAcJ590Act37/v15KSsNmSALbSYi5XH3NV5o4vaJ/oefJnW0hPfu2i6
Rz4KoNDTTBP04Prf6CUJ6omhaQShi2CQvL46lN+esY6/3j+neHs8oIKBjUDP1VOT
xJ2SUBw+oQlIAwdQqGbu8cp1iYUrHS4QiZZ7TXWUdv6MtqwDT9Iyrfi1aTcu8qgV
mNy01iN2/nA4eykSzrRxu6mu+CPUT6pfFCV8RQykjuuxByb2OTabApWSGbUAGy0k
W8P7hHTUwNc64lP9ChicHhWLWlZ4O3XeeoXL+rn6A8FXY6igRMfItq7k6e34oXQl
hyoLYPlSC9ciy978Rz/iKOdU6805G7vihauHv9PgcLQI0P7GkUm0jdOfKc5mYeBE
i225nIFH0SbVfX+kR4hMtMRt4CuM4a1ebYvVq039AR0V3Xos1BMu+Df4fRYzqwJT
Wil7EWE8XLErZjR9J//Gy9mhk6e5K1CtVIfCb71G+jizdu0g3HQVUBCUc5NiszCk
G9BSXgcqbacQpjDO9BzLoqZ5MfkiwT++DCfeEgKL6O7q5oIpUS1ycccMagD2Ghu3
+HqLGPPzbozi/83oAXtM7WV9OdP3NE4vFQoW//VZZ0BTHdw2qLSbEPgz819mwD2u
LwWO5ef2H+wXDTDubFce9Hb74pQ8SzoeDeaAHillvEgBSlXxoc4T5Luon8xwIX54
4YQ4u8cX7zqeu/VWP4tqNAW3pKVnkLzwHIZdKBuJCOlZpmw9uOljTsZcggnghlVo
GDnVqwvCcJGV6ebVsIcExxfzpLuVS3LVBoZSyoiPpceqlWHIRkXAqnhVcrel9/Ym
rr0Mn7B18fQwzBno08biNp5CPYWCueDhEUIK3J1PlayfI+OWB2LZuDn1NDHnB38y
lyH7WM55kUDj+C0PSj0E3aL5t2zi7EltP4cAnJ/PTfVMuuqKCEKrRhi4pq/1Yilr
Wyf+sYDWUVXXmXMOuYG7nJCKHa4ppS6693pE/UqL7Ux5An43UmS9+NyHzuMQuaP1
E9SM9aNRBEwY+bncmXU8gQHTCQjqKtSgrpTaGad67mnSUVLNaMUdZARVt4lpeUqj
J8ar1A+qQRPpqFPefwntxeRyEzCAIeMCxJ887WAEvkH8dPVCg6pAHsoiWuK0G9pP
uxPVbHvkBPhNMtD6bFWoSyEkcHmgnAP04acjBKHDYd6z4yOyLXGLVxAGzZsteIRR
vzMdyQ5xrA+54jHhTx4y/318KizCdcoOUTtAZ/eJzcV26thmwPkqACAiI8rxjjPE
g2YYXDsfVs6G07PLvSHHpQYbSZ1EhUbgnWPnNX2pb2GhDJ8verVIsBDFRqwONSBl
xHDcNCZxyHJZzcuUITCVWIfXPqfZQJ+YyrLhPxDyRpanTrkjD7QnkaSxpvH01zRn
74ZjE4zUoTIUCvB+YPbs5wiIbeeI3WUT8aJRWmEh6k2lMHCp+z7IfBi2y90FrWgL
spz12LoJrA/mz9mTBA6rSAE8Li/ZJ1liJsSImSn3NdzruorcuNCuABPHxvQlMKvT
Jezs5qWfLV9R+jDuwU6V+uLCi8u4MVgmMyA4EBB9Xwm/xsxR7gxl6VLTaPhRBiyZ
qJAJfOpdcHKAUy7Yd/dHnSNZLX6Baa9dYOSAZRQUNq1c3a0MqW/Bdh1IKyUuKHHo
lvYBcont1lMA+Ea2+6JThoUf59aabnjMF6KdiBVL0RXCDdlbrJbiuyNWvBHcJKQD
qfO6THUZFCiZ2zDNBXFFq2n4pcNpGYGlcRPJGAujX4kok1EmqanEzyBb67wUJplM
kgx1Cxs/IF8vd39seCHd4urvXop14ocT9saZgSDMkHawym6NpzspBwbZbZk5qLYk
gPDrqSNRF1Jk0XX0A0c+AQ8n4SPPEuKwMImYYrjgBGn2BwAlxxPhkTEspewEY7fC
4COqndfr+w8/eUdPhi4eQzvw9cHMuNsbBx/FJxgpnkhUJv+nIn8O5Yqf9048iXbE
vn63F+cUt7RuAMm/0lKqQvGLzHfLQLXXZPxzi+sBlsz1u1HGVCLkwIL3E+7oaB2+
uhlQVOY3FUjw6folXB3NZ2G1lLn2GEJZMi8SJ1gj0eFJVtp1aFATtjz8foUMQnNM
7zd4izy/mZyzPJs9ntCGeauwAbKF8gzPrjsIIwh1gsi8omkPmuG3Y9oi5tl6N0RB
mXfittw/3WG3UZG+dDVlcQMHaUw3UD/O+30dR1tbSIk1f5eLRV/kWNyagyhr6uRo
4HaoQCyZKoJMl55Nyv+fEp8GRkIKsk/UPRsNO6N3s9AYQqhSX8cEyZkcb5xTOpf8
pPUItulng4GhcqL25PEL/V3L23nJRVqnLlhMT1KY25XarfL3Won5VbhPgv0JoTo2
Wh4Bk3JNMO6gLY5FQEZ9mD/ds8bEpVfinsbsV45vnCPaB3waJv4XzqYNUXDfNwGO
zr7bak0B4VEkYgWeGyQ6InOnPMUfZuRrzveogi5v342PsOCmjYVaux9nxtbmEC0j
7nI4U4XsShxvZ4xBn6WJkDz9uhXYb4rQy7t1mjqiSKI+AZ/1cBN9AaH1QGudv6JV
csc3iUpsmuJZUBo3nCePDWJ2xq5gwdY5yEGuJliL8Lv12jBt9fa57ytz9prjDiwn
TQuZvA850LQbKTAHU6HL7E5g+x1TjaTs7180GMNX3VIBXw/Opb4T6c4/xEDvqsCa
dTZJiJt0gVUXPSVUV8EyTmEWpPrJ39r8L5SVQ8igJ5EesxMmdb27LOS87lo4Ea6d
yW8CQWlZV3UnnnK4od0bc+ZYD2xhuk9P/Ltp3oj8QmasZbA0+Rq2etfCo3A5rvz2
xQKQwG5K63MtAdVESaj7ev8vh1dQiZm1YQTtNIdJJrOWAAZ1BA3MEvIbWIpP12/9
UyedQqKjqAaknw+I1rd7G52nsS+1HYWbbKB4MEHKG1Egdfc+xyfXgoQFO+qK+nIg
ezwhOw3yhMfCPD20mv1l+Aj0PeGnixfIgH6XPiFq9OYQh7elrxA+i9g584C3xku+
7M+cJR4REQgvJxVnoSzdZn3CknqjwEj5+qxlfz9tsXuPdxKgpgLwbvLRa/OVuW0Y
8vua88l4KVdDX7wM7vk4ynlj0pzAkDd5jrjzw+Z6azD5egRvaP/OTnJHjHZoRfgL
BvdBSv8zjfuiM1MFGZDfRaT1VEm0xRt02MSaiy9h5i8yhwPQkEPiQNjWkz+SPaPv
dRoZe3J3+UK+XCwH4TVuszgSYtERdI5du66JSZN6fTn/esMkgmp2tGpf7Dqjc/lH
FL6Xe9clzV0y4YFyEtFdx2uwe2a5jlZLqZkFtvl3XWC51XSo2x8Xz/wKVs83khU/
eQRJ3Vt1aNKgipwNYkC8xo8leIioMKKAQzvbnBqRWr0ZIBFJsDRYvm8muPuKf/Ox
wHAeHNwis4vnBi2IKTSwby0mKbnBHlRIn1zR1voj5huU2/aOPdLdsRrUEIypbReS
SXktvUGSEIY2Rxp4VHEE+9CP4bFGoeHxTlNt9NWWnbUNPiKGlhGWCgZaCJd+G8TF
6gAusB45LQYiwPDx+GUTsf6WcDTntD2YxSLhBVxXyBSGoROcqQXazqwkvrdpFlG8
BVbtnKMXjfuFjDG5DuyS8z3NIH2afhUg8YGmTJQfFPajzHKV56esXW/4HQIdmRWV
HywncdxRo9VEC9qRFLJejqPcomtdF0/MF/JJoM7ruP5i9snbrUAYEQT91NhmR/Bg
lBJnShP/qlHcVdp2FgFPY72b6Q6AHoLnwy0vtmpvlQd85EcXp35VfHD/q4+LGN6F
2o+R1vLmu4Finmkvm3VNAlXv+0XYP55tyiVC0GS8zDxx3Jh5AIav+Ju2jixzNShc
aoaT4NWS24APZyS+3imTl5+cKNxzp22UNp5Nad4aHSQ7gdkySkBlURN/e/tiJPPb
MVwr5YZWFm6cqdh1fXABb5+bAc6AojzGRnE1yEAt/xO40JWOcR5bfxkHpKPd9sst
H5Vew9VSRDe8/9pouTs4zCJTzhrOY5qUAM/PVb8RHrQbYXONYnV1eGCTPn0AOHne
WChB93nZR1sdkpHMwth/pVu+BH14yRD3mwI7zv9xGQLzxhzwqVTM+Peg7DNhq+EW
R2Jn/NicneMQy31w7xbfVj1T8I5MPh3CSc4X0771+1sphsqItLBSjBjGc6/SDFgT
m2/51PGLsr5G+4TAedL4wB/YhB4cx6pvaaLOys6kby0vMROKbK/lDFlgHzFTgN1p
HSnnTRhW1bheGxxVKvgWnyJyah4CSjMm97SL53GpgZxykh809LioeROb9dKho2nn
jvVlm8Mdxfv+827CI8rDzCN+H/c6xEKzA5dLQT5kLKzeUfuXovU2WmkCStPNmcQV
jz5eRSiuzrSOrPEutD3LPE+vPL+03Jzmhh0jHEe1Yx49ZxKaWJOUFAy4HMGAt2AQ
g1ydtkL0aLYF4V2wpP3YeysVYk11F3RL7+fD+L2uSVeuQ2h+6ybpLZRAUt97ZxD4
2s8K+qsyuecu8sgnz7O+YB82Iroa1Z33sdh1EshaExPmAzNN1AeLOdiekFrb+S5E
APvseqwJjQChdevsW3wQLDbmxyDxNFYPTDKgRQDfbrtGFy5nhG9yhZnk2G2tLOo9
5MfcvO5OKGyfLzUGO/s/QG3c+yvI6u0tF2yCc/989gJraCqzp8fjqT1DNA3oxI2q
AlxN7uqsFx9GQSRVYxTZ2zJxqYFAJikn47T4JdLhnEAMXeLKlOG0Kk2WINFI2G0a
McM/EQZVfodOQINaG0SzLDdP6/2IR02qv0SqvgMamj8kqGbpY7XuEjZBhVrqCdZV
PPQTBqWk6oNryuxvYe2SaM8iSXm0Rm1FcMxSupnbhIcqD3gyY7wfure92YmTk/8h
u+jOpR22M/TofWDyGMY35MoBse3+l69uKwVtDktA6l3DQydWuD4KJfH1jka+MYfP
7Gbc2MHPbTE+9noqbHfqj7wEz2kt7sD0JMe3BWwolZX6Y8o7B40gExquK+fbQp9Y
ZYVMOW+kLzc3aH0jPlNwdQ6c6X2nBuD2N9JnJUig/yKnoQWmUQQQepYLD2mBFMjv
iPBV8VqJ68vjaH30+zJbspxJxXc9+UCyFHsUBqYUrRRxbDrkG8DlE/NObYOe8gup
0gIi8YbCCfFZVqyvW/LaRbEccontjI0p/NLuUSDlV00RKTQY9D3RRAvW7u3+922u
JNyLZAVO31B688bo0+H1FD4SvHZDLUR1Zf5tXg9l8oySMJNM3K3HOen6ByFxIErQ
C5E62zfuOtyWWsVQe0wZeeQbrsI1X394NmaatuL/Y88+3WaYVWDfuCMeGcO0J4XM
cSULwq4bUvfbhFehT/6jKdPJJM12x/0BH/UmOPBdAApGaO0nBa7ROqQIYyYeKteu
+rSl2oYTAM+HNsRgfiHCF1fL4ddcHbgK/fK9pqibD+Fsc/X+AigYROTC9RLdzjMa
8GroiilLBiSgqWU+gCW8RBgSQX/U24c3I9gxpHPJCQiySXJerxRRUlWkGHb8ziLs
efJ0tKGx44cLzgLACsI+nZkUCwhjTQOCNQivibnVQL1j8J8Ma9QJHDtqLDFAdn0l
S1HcpnR0cG4g4CShE0gEKNK+/SgfbkpSVvl/UqCBHuixuldAAegx/IexzsH/KwS+
mcZ43/WNt6YDvRgjn/XFhAuHpEYnD1WSXVac24trmCYB77DxXOHRcWwW2t7eezJN
oODoo0C1kq3tNMmr+ABNhzUpXe+WC/ta6+JKUyfyT/T4StJl/fs4bCnwhlvAxyv3
xPuA4Myl/4IKULnhSoDyXdFPJ1VNhvfnOvj04Pv1brLq+/lxX9NwGv5+Kr8STfzR
1P2O+oQKijYeaWGR8dSMe2yElvwnTUEMwqH6LdZHtEQtlhWE0m7OPKU2IBjjRXi6
8B0W9v6UgWyiWsNRY0LCDOMGonbnx32t2CdWaulFfcX01cjK5m+rSTSOFnsZNCwT
WePwTsG3Fddi1E4kfH0ws9a5mJXU92BbizVfNdk5FS2JB40g0+eUeH0/9BymHzEm
skqgxSV5YFAsqibWAz07X+mrc5UcHxWDUdJKUzwBYJDPYsuhzA1tsSNG5A+d8BH+
a0wgePZxputBTdNGfZ8xDMUe/S80E5HsGxheI1akLidRLqM65S+QnFPyA8BRMD3z
0vH5jAMoZ29nhnpGLW6esP1bLsjr6WhO/L6ON0dYkSdkCZZ4aS3OpveC9KEFqMi+
VzN8fDw84bIj//r9jmHP8dtJKRsW5K1I21mBfcw6AwsBN/xUj2dY3vHuGOYMU3s5
ydq1cgny6H0ZbXpdWD4CJx4RdHxw5ZgBaLEAeQ9HBc3mYcvah5SOP4YjA0Zk0/J1
DGQeliWJp0GNa4XgZHhTHgQ68jhFtLloSOtGeTI796fM12BGsZRQz8mbp2BvcZ0q
CMxAnSAQpdtmmm/gzvxgLmlUH7BmUkO32EyVDTPdtX4Gxm8r5GnkJlJfKnebq5E2
KgKsLeYT2zf0qwqLBNbb883cAO5rbWtVVvDWVNfvAUUMKjAdOArzCIW0LYbXJ2D+
4AsOPsyBRf/UqPhR1kNpx5gJ64EPt8MPXtG98qkg4i43MWY3xBEVk8EvWkR4X9iE
0MpOMwTIDBZdJWBIxB0ArDcs+VepSugAAJbKkL+uAk37MzJ9UgufownDWTdhXh6S
LRajIFESZc7TVRfAZ+LRp/X2O+/ZJTUVTwyJuVES59DqR1dC8p2gjsbscLjvF4vV
xBFAG0fyx+TlaVmW0pAIxoQEa9Wwm0nBIqBdMeLMShts1rkUyglF2CywPuF9inU3
I6VwbmXXAaoWX+q2S1anquW1XP2GP0VEYS/DBf/yQoQ/2byCU6Arwrp8+0hk7C4S
/XoEZCdif1KjAbGgofWDoQEy4mlXCNbpnJm7kd1jXzqa0axIUg3hrg7u8EDqaH+q
XwP3ko+GcBgyQAeTlZBP4BQeouC9f8Vu0OZfz/xFGz4ptLiFJppqWzj813Mf/+KF
rq2dCU9R8AnoiIJExPj3dZxtmIQ6mrlZLlrflwYEDdc7E5xtN/P0N/IggqBK3Jhd
Kk01oNhvKOVAlWDc9iRIwOGIeox4T0hnqu5mEFxX5LJSqRsh9ia5+pl8eu4Xg85V
J0iJFwbEY2ps75REcn/ABNWna+dE7MQF43hV5rpF4oYeUPexwngZB9ja10rXQWFi
3loRDGSPVisBF8IGBzDCpQHNIeWwOEAuVywR0CPENiHGUb8ZRs/0k6/NxQmIotJJ
xYy+TncFg7olgkTSNV4APDsgFi6xSYjgwZQHOle50NFZHyx2bRMsT7aF3+9PEiLt
bF/lYRHD2UUBo7IXh7SO47F2zV68iQzBsjpFUNVqtXz8mhBGcddthAP8yLYukq5X
W2+2M5ljJQROxtXdMbAobnsDxObtoeg63ijRDT0/AFV8zBFeCjhE2Q6MzJwwtAgC
ylAfU4GDeV4OTAV3/z9INxOK6vKt5Wou43nAz3BPJBSKmMsN8XmFiaBglYlbYANY
Jr312Lj2jCTzmVqZAeWQLPHwHlfzpjSBfvBgtj6vFb5jDP1hv8iLRxcvu5bcoKFU
U5SLPwlEYo1mWkj33T5UkCGIhSzLt4p6PUN61BzMYwvvSST37YxF36+YLNOZm9IF
xr3ytiOflztHllZPW1qdmOdiGyK5C5ULkiB+YKENubPl+EV/ULITJfZTlX9vFzjr
w5Gm2ljH7DwqdkT2pYtDY7bgRy8ySg2tupp/C1j11mDKCyFE5u3lWg1KJRH3VFJ0
SggkIf71ghtp/kjcjQph60WPwUVKRUOi0le+/mFnxANbEgO5r3uO+68BuNfXSlrv
FVZRY+vFD7wdXXecVMEKCTG/sklrMKrXNYkZQ6h81Hjk/3gRbp2aW0DZQxVhZcYx
w1eDjQGBZJL1WBBVR0E+2qUfxMcCDxex8TaDMgXp8j8PbrZkGRKBQX5TfRdB9CwM
VreXlqpHCENXwMFhUXmRUVSuoai1UT6n7XP2LxjqVRx0YZtk+UY/WFwcHhN1Veem
IhS7bCNIOV5XJ8IPFflduruDl82D8pX9YJ67nh9gCGtr+uwF09vhygcFaS0EEjcO
dJYJbioWdY6XExUJf/Ti3wCY4K8bD3cx72PVVm0n8Or1nSfNcGBhxXstfxSuQREy
nfG0qrHBgfH8lCETTxsofv8Yh1OnGpX4P/y81TQGxru6QXh2SUTPDFbgubxe12mI
ZlFWlXjo9c3+krXcEfnqrJjquERMaFrfT9vPutbGGz0qfO+bUAHgp6T14gjKB3Zy
hL9BkL6uYTZBfCcBikDsOpNhXKwvIIvm52hEqBuROvXkWsBkjUm6kXY6KsavUDYz
OVvUZbS2kxCpl/JMjxt3lQAp8nQTXs0tT0syG2nDmutA31xpp3DGtc1/Y60iFLPM
ScOHXMcttupRjGxAv+Y1kTDXmCjMX9IFGZDUrpLQjSs16+HO0So/VeObHsKEgUa1
WMmD6MUJVSUcw9SXHL8t9i3bM5EheEggdXqOD/X7mdgBHOxrsHBu+m+T5KiWQnJZ
EhOdJ/Xw3fN3uTeccChMgiQBlamqkc0HYGhxs/XXpqEvM0IMNxqgXLu5AH5UCSSh
kIHU/XGq6ocSxeCPl6S/a9rhBFwKOzMVaYEN7pBSzGG/ekHY9fPuGxWb8un/vCzn
bfhzjJOxoRXLNn4PF3Y5O0ck9QmlfMNR40OrzkdCMJaCCGzKvr8Boi3AK1m7nw7l
nWEuVIbD4Iv0QtmcoQAC484OMUM67gFe0APDiMGbWw1KrQLw5U/m8jhbMwhvvG0L
k9m7ClvG8PLsZc1JAC0DKUxLBm2wkAbHQTpRa/Lh4k9uQH+vMkyGgtX3wzfuVvFd
lseIzWnGk55Xe44/PL0opIgxMrGbZSBK1Z9NVPOrTKaC2IdVkAP9OXkiY57m+Bmy
KPk/Sm0afrCLsTfuIKq7nMRbZYoaVFRMaGgrtFAovyPeJS1UMcyHtnOjU1nyAQgi
4OoS5fDUEpoCf45DowrLXee7dBdRlXtPXTG5G83J+rDGozF2qKAGyrF1wWRrRI7c
nLGNaamY9RN1Mv7Cfrm2Z5oiaMyfyEHua7ktgWxIWmb0SvAuXAUlp6I+OUxics/O
pO+zzdFTAmmLyG6iZCxud1RHH/a4PV8Rrq6hgqfqxgEpsV39qN9pEeDNZMMvCfXl
MBZ0fsWz3svClMIKQ0VQTmRpBO3TNUdTGGBDd8tNBeD8aR2pp0LVnm/BOwwhelnu
xNgzhWb5SwnwWS/6WBGcWt3I9GaTY0atirgvKVy5xqCW6lP/rSiO7ZX99olClPmZ
bjgAo00vIOpMwWgkUwY8k3cgnBkXOSQ9yyxqx3Ym6ylSBJoKoCwH/lGWlwDQLFRI
b7gfBBUk4/UuPP6htNctsCRDWUfgLS96Zcazc36kRxfw35HejeqFYXBCK8d/RZNc
8QzxnECgCX1bH8EQ8SeGqv07c8UrTcEkbCFG/+eS1u4XhA4Mv91BDMqlsrbD8/GT
DWrMnbaJzsHT8UUQxCnCA6OMj9W6tFp6G6HHFAcVfzjW3Y7AOGSewjVbb2hihvZn
aHSuJnRYihlRZmA+cSfJKkbP3wd4w8BMubE2rRIGYvNL1JSm8r13RNr58uZWOUpz
LbuKVwJJEGB4883WugfCTjmmTtNcrKx+vlwzW81Sfsn6dyLg1qA12UtNukw5TjD/
VR1qTHbf8mtRI9RMFroMFWpIRverbkKclP0fbI7oZjZgK5T0EplAbcjhzqCqKbid
+gRUUlCaUt1ciWGgAKmWKF5dY9WIoBFTwoimB/s0QaqymrKOdjrvMpa0RbMBK4w5
TCQ5vNXe3GnUT5oTXkhvXrSFb+mPohxifUvHF0dVMBxy6pMNignGEttB+XC+MKQ/
JzERoIRobvaSd6VYcCwFucnlAh50S4A4Hqxyw7zXwE2I3N/wyosIRuPdI1p5KWII
/ocE9lGoUGIo0NqUUj8Y1lab0fdsW/Vc+MjJGYxYVU3OhYh23AdnEQN7TLoYDvlk
HkGnjaQy2fpVKKupo4GA/eRkO9H2HBDA9gljnHF6oxtxua1hsVjLJw3e2kzgefWq
WdgWd1TSquK38kK/pag0WK1dXvxF6kr7D3ELGqvOii0lALrVY0Ibbvc682ADNmxe
kIVVSUJtgvYjkKxCY5LJ2KfMGno5qb/Qq/ylo06CybpZguK1AIkr1PYDylVQMwS/
/LMN7F4vTazKLfPBTcG2cykNsBh0u7inDqKlnMQ7Pf/rBXxirERCCvQmUZ5f/CjZ
pA2B7IiAQRvR5FGSArF+0SMJzyQekxKbaawWiwu6pMJ1lq05epcqjBzq1MhG1HY4
4tdlu4msdcTYJZaS97n6C1e5kx/B7fpEJ9iQoBoL6Hr/cF2RPmu4q2ffBEdjzVuU
KjVMKZn2gq3M7CS2Db0oghznhz4Yj3DJMOHBUC85oOLPvDHonw5Jk8WkH7eB7HkG
Rdq2ibjCwnnIWQ4gCze/y2WZTmKy1oTlKohoWqam4kqaAgpIG4waPNUc5KhjRUuJ
N0+nwGayBjo3hb/p3+u1K5DMhs2CmYndBBwL9cav6vk0//1OyCP774WyU/cFA090
/sLSkolhYUY6o/Y/DcMFugBCiNm0sxVEE6JRMtFlFuayCsou5CpM4SA2pT5usP6j
Nedj88QkDP/t4VYtosQohKFSxuL7Acguaaly0mDSqulg8pv4AW31WZjpO9kWBtb5
sJssLgS7piLem9E+GUh8YheG2Ftlq+Vn9X3sBVrIbV5RkZ+enn1hRKoZk9nMxX/r
yup2QYHLvgCvleZDu2ZTIX5dqhLOBRdSK/PposRisv3e10Gfs2dRS+nr1BwLmC6w
AXsk0/LdDB6N3zMVTjN2bZdOM4WjlRfQQl5VcxEowVKsbcBqyi+slBQrZi2zBNSs
78VFN6CPQCDEkAQ9RBHblO4ey9EQfx8JobPVw2wf2wAhZ9Da0z4gLHd+oVTT1J30
lPnJvtH4/CsbLobWrS9hCC7PzKm71T0Iplbh4NJUFOgHTg2LaG9dvGzMZo+5Bv4f
pcY9fo5h+uJOB1rt3AeP8OMGA6Zfi0FLsGPlCtLiODBNycTgSeRUOMOInRidMSKD
3+D2yB7uyCuRK42peUv2XtKKZ/ZrAn9Ll+qGWPxStwxGQOOiAsvTAA7mRyQIV0Wo
kWhLLlHOUdz3QJx0/eieKX/UOs4tTDz7Zp+bCwtvK3WkLRVE52bI7hohRhH7SFbI
E+Q/0FHhzHCHtYVMFv6ItNjkWwKC5D7PJ99YaCKVfIPNOAOoYped0ppC/K+elpRX
q9smjdmL5aCvlLTHj9ESIrjst67hGx9RdyTWE6W1CZ2yXz2SFO3M/aaySgWZLVix
8PwWH4qZje86oIu4lWOpGtM7tf3oGfoDqVUovFRcnuAVQjV+NtYxgKadyvFD17Ef
2hPb4vWdQx6jCA6CcxHApwfdpzJr6KzsxeZGBdhwBi/c0d8uHMfY7L02SMzEZPwx
5OoiwJXcGna2XNd3QdJptHNwKl2Q9+wBwLkkDE/O9CyJZ2D2nrO7WhHYUNtuTr2X
0HqZC28EXoRTC2DZtIqyXQLL5GwQ/8nlK0CJIUDNrhe5G2I3M6eM+2XOnzkCjeJk
rAEbEcd1fFZKKupKRWWyufwMSvFx+AVAw1lzCtIpoWptcmURff+Gfr4t7MpukJru
3NvyV6kyScrFjRxHF0Uiu++vRQNcvTIjG3bWOvAUnbkB/wYF8rniJZ4jheSb7fYV
KNgSjk3e114QOCUaMNUTZMLt9nlfm8Q/eOjwR3wIwq30WA2S8uzp8GCNaGsAuRBa
rSw2m9DV5DHR2ClzoT1DoLIAhVC6uq3RX9nrsbId3A/XcHAk6k0kJM9Kz1TnT28e
EDNX3hmni5coqb1ky92rScZOeNbaISO8dGkebl0d5Wp3fy3lCPtCSzMpLPViSYaH
qAO1/93AhLon3dXXDp2Ndy5tE925GIW2X/ZwrZs8gnBBfRHEuayf5dY5686isRdd
dJE8KB97rQwCQmM9e53mNW8KCtmMKlinAMNZx+TzJy+zHHfL2XzRjfUrRfF2A7g9
2LtwkhnpsRmETvtXQzEEBfYwdhrqtdRtZvk8m/urYxRKpuxVZ4mlRVNECqJidiz1
PxRxyv9eEDygQ/lWWh85LchM1SRrPstuj4o3O2C7IoQdlGMLGCYNGOpCB1u8pxih
gCfYhsg+gTc6IkqZhOI536KARWvHaQg3rUOiD0KlczyL55y7WVv4ZB7j1G4YOiRo
o3QD9Xk2L6HhvH8kgjo2o2uAyRXkPXmdvfDBVNDGdVbkQio5ASnJasK6yg2U8jWf
XAZBwVTpg1xfEKr0+adlEx2Wg87pxMltB2eno9Domqfo2l1Q693gqHFpQgrOSmln
yWF77R+w8ZNJSU0N289HTiUj7eZvW3+4GGtGz5KqpeOer6DFs9wZM8zaYm6xWwdb
OoNaXPtnmdB00uidD3jzBbWZ1ClQi/KijttqAxJ57K+53d2enDgS+cG+f6xO6rlA
8JFgSRvzxFbP3h90pGoQHJ74D6CQ/2zLyrAPEQM62PqD155kqsT/XEADaSEffdH7
bTFbQ40btkvsnq3LuI3bB7cj35bu9vQmpAn5oh0FHMjtPMfQTSbA4y09NgMQDa9x
RVf0ASbk+PZ1GxMcJfm3VG+qIJOC6cdKdfW+5Iu7LpTuaaK49rwjCMrV/ZeBo4YD
JN/8lATkMwa5g8BtrM0cQv127HCiDpnd5gGKRbieb3lhQSBOB0wPMsibL0vFTi8J
PM7JQS358pI38TO28nYQsrcgwyyKdYG2P32/WpcA1ybAxVOw988JXzxNzPcz7frt
oeF7NVfJe2UgRP3pu1ptmJ1BgiHqDNxX/IDxz/Ik+VWUlPlewHgkde92jCMhUkFL
t8pgw3cEa0OkMFGlyRa4ssz2r/omVxO3pUso2NetSp3Ut/o0Z+Zg1p63Nnb8HxQ9
EIHNhbmJjqz+Ix0uG+XpHegrS/9wJ18BzebwT0+bHSYq9cPVC6BZITxMqvT3XqYQ
0JmAc485sMQuU7LVBO2cE/HIM5qp9TjC8MV8HdquThaaQmMH0RhRvEQcnRq5RRD+
KPV5VAz2sRPeRAU8CLigQYVnFBe5HQl1a6c4bnFyDu3wbixz++uJU9ClHAiB54Cx
zh7Ch4uHwBpetUs5hI25pYA80Kiiwn+DW4X+UWpqxKUZQTFJkngZMduC1U8fxCCZ
juA3PKmG6KxGLbZozy146PRKLNCKgurBpXi0d4+LdIwnYYyHD7Av5SwMdEWnFDL0
3Fly+9jdNtnRXa2Tf+9gmnhGNX760QdXcnaquNdGKVli5q58ode1ERe8QbX6sjCJ
bpbb7mv/WJy6N80Gb5zEYg5W8XEfjkJRUF9zYMncYnTt0+9C/PAfsLE4J+MbA8Wv
iisWXFr5gfudu8EMgvisQRod2OOt3hC7uA5Mg0NpqQ8Sj2upe3AaDBuWcR3ef3ZV
0P8SYGGkRJl7KAxeoADCuGWyvk3pX2x32BeeOGZhgo7AzkcWlessP8zfJwDeu9az
lgxfx6eaUockudrlBHqqZoCyByIHrZjWFxFZmjzsBIhiAXHBCq8dEP7jbuXxhKYc
yBvzonTC5vhF+SChfsQI8dLB8om1qojFJy8Zis/e56MJK7bPyDsXAI+eSLKl4yCP
a446Vy7JHKpHzkoQT+2Tic7Kcd8zR3UtAnPbzOfKMKCTpriQPBBxD497wVl0CZdv
LzuG4UibWP3/reiBsxKTCQuvloW1fDJ7PLYZ6Ib0K8DXJacu+bIirUdwD3sQXeQi
4YLBq1AeRqd9dmcrc7imofRs7FJHHiX2/cPRrx/ZVtPKavG4UkgEoiYfjXzUAp/U
jxenzO6C/weX+MnomHEudQdilFDzKd+I7pKMoCovQSU308EAT53ww8YXYHrFif3u
T2aR/MuMEEg+r2cM254k4wnhh8OlGz1EVq6njRVumFtGbLRO1CfNzjwidGpw+2ul
ssC8ce3HFPSc3ZqRl+VdFij82cZnJgloFyrIzXPG1PXdoqrfY8DYLhc+pe/jY0uB
3uSRnVWZSJD9Ng0JfvWOmMt+YiV81WLl4asOEV/hAeAraAkewp0invd1FW0/9gsk
iuirku8qvyCcdLfDNnv+nK3X0hG2q7slQei7ze9REJ72shlcNRtO6gLZ5GNI4T7O
N7oiONxuqeWYpyamU4ED8woSsbbsPNf6pa3qBlFXavzFZY9F7zjvIrVtnHxHeR+a
t8SXK+scq5ZlF3LjqQLC8kwccvWv68uNARcaElgmxUUK86G8Ox4v/bSS4ywQqWAd
F7JVHUZE3EAWf0ubLZVFo9aRIqIzN34tyKEMc0L+jxoZn0S2JYGr0TLyzJUhK6lj
n50fAxWtB3r2K90nlJpTYhz6bDNb9O3IFPTATuZQCwJvcI2DHVKMcrcWYBbIM/F3
PQDcGQ5OhyxHA06AArs0U4Z4aPur5yH2SXxDEWh89KgU2yc+fQRGE/6bnkUcWd+g
RqbqJSOO+px6Q8ikHS4f2SM1lKbyOX/jq+Ptr1dwAIyN4JPN5tPL2tipXT2+X/ab
lIhpOyEGFukgV+aO/kPE6Ja5dJPjFirci8/FeO/KSSUwDIIbwVccNYkV/m1mZoml
DZytBAKs26tD3DjjhNx89iEwJ2Tmp33zPfydU4AHi9VJjDAqW0F/fyphvPMlLwr4
ksk7er60bDA6kkg0x6zjlZgVVUmyF3JS4QjbYBE5jq0RSzbvfzPwmyMUITfmF2xc
pQL15LGdLFGZ4oUzNGAbY9PrLOWb3eFJ3sGewlUA78l+EP6wX9d+p1fVJugRn38H
gNlYSpx82ph+/slLiDvV/zSzuXmfwWPCaOaF3fAQhpMLWJ5BuKlp4/Njlm3zEW66
Vs5JSJvlwZyetvFZZw1025cpjpkjAX6N5TZX6PeBenHoP3ob2xhj6kQtX2tbNmN+
7L2XAopY4rZKj8TG4zLSDQx7Hc4guFo8gkIU6c9MGhfsbLUOADV9sMvs10cQJII3
UK2IeztAKG92fYSFxtPLiEq+xKpMt6b5woQ9P4B9AwBgz0ByjBtKuvx05ocNlRmZ
I/eZiAOoOlnmbiK4B6z24f3g/tbXqbRSME+bFAX7vfKkZfDQkhwVspUsskGGOyTP
HNZ4+tfUv1MQSrEcy3NRVwF69U642hmqKuahZ+bYNSSmxbHiSFa7FjxZzJZwhrHe
wWb86h19aeyBhVj2pma4zuOLUPZpKD73tolhOmMyb2UXSt3+HA1QhwUjHV/VhEOc
tPUW17qlhOmVT1vjBqzBaKvB5jvU6TNtp0mby+tSuH6gwakMC6exuUNJyqnNLKhc
yy+Dws6upd9v/bME3XTOGzaLUt0J8EkG8pmAYkKMvploP8yh2CVUXSZq72FznvxP
y63kOeX5vPYrBJ8c99G9AZQWx2Ntuy/rRIPoPbMdJ1sm4iE2HWlT3maepkH4be7J
/iK2erAFwkXQq5cGnE3/8boiuPcIfI7xBpSHoYp4HoH0MSqg5Em94wiPUQRX8klE
jzq8xuXxDkAyEg7sepUpDJbGKTJm4S3KyGXHycLeezDCHoVTnreGjw60apFLV2bt
vSZLNty3YcCsX5r0RxFNHotQV559EhONrYzCb8ONe0XZxZQY+Ci2rRPm0Kz+qxUm
1h91mffaPfD4c/8CI0HRl6wVYCHE+P3ViDCV4E6sl0VO1XuLNGlj0T+ZKYQhQjG9
Dm7htBKm/bPaYQzaiq6uKo24QFr1+AA3cAW5hdcASL0LVY6Owk06Wsz1FdIat/z+
g+YW06iIsdY7YcOxH0e7BS94UPkJaUebnI4T0x65kQ0ba0xFp1hgIhvCybqFYpqh
7nJYnuSeCx2F0322uJehDRz/o9vnYakybwgA4z0gG11vGP07sZffHugr1nB22iIi
cIE3j+qbTI5kzF83HH+VjJBVF275oJ9cjCGtBUJ1W6pUHiQzkXOISd/sL/U6rDen
PoWNQDfyoS+1EvBhlyzt6WpbGy+AxzjCR0FxoFst/fMViOA/hKB8gaqV4/ZDPDnI
mV7IWwP6PhW5B4PfcFa4szL3cCuVzwkbh70tC7XAcGz/giP4i/HzJTYtPlClrKel
wdxjnsDZCpsUaB61ItBR+mQNA/YgWSejeUJP2mHtc6htOKaPk4rFYhaEwot/ip0o
Mk56PwS8Y6oKuCrZbYctm+35UHo17wLmpXJwRJdKTetoUVb6VejrehbN7ywlI3t4
AyQHVHLMh3XDx3gqZ8FHskSNKjMhUF4UOMORXvCloXmoNPBclTlb0sN9eQUDe+ez
vUNPquGYbV2IHFpdadBWzqKp3kfKwOZXTnZ8sH6OGii1iijsMIKegTYPnL+maJzU
KcOiwtB1VZOeYdDTzwRahJp5McaWX8BeVWCA+IsCsad0IVGgSQvEd5vDZFch+nK1
93yZFExb6WPMIR5k+GRU0o6ZlVcczMgDVqTjXy3vlZzOJ5wtjqWm9YNqRjBLfqL9
gJtA0zKGv9V5bu8oyujqyv8juqpXtnw++lwl4nQpg+7DAk4QestrRELBTdmpkDqX
QAAgjffoEgXacgz31Zk+BuSIvBuHyG4Oxmyxizh+i30nMcFuwBQMB3cqKNukEJaC
7j3bA165MPeAbZ6USu5SfjJ3a0DmNygegwE9ijvzrlcEuQLSr4fFE5F3kayERS1K
fgpo7Y0vOTtNi8jWwUqn9j/1HGFnmD0TQp3Kp5UfUmEnLZlOUtKgFqVTDeLzQGFO
Cr5SrH7cBUB75l39Gz0vIguRKvX3lS/wQ59OzmXeadAsINAxtEK+ppE/JDQD7D1O
7BwgK4GIIF83/ehhYjuNEF5OsX7dCfYnUq2gTfUzwhQtyfEUNgYjVp25EOxxDOCX
FmM1oDtPnRyxEDVyqZXegn4fW6YisQqra8GNDmodbvDYM3mtKv2ym3Ag89QTAzSB
kLUnAKLlyyK4M0u3H+HzTEr2/HbgWurR/SicQ5s+ohzIYwJcfOIBPM8AqIrD8aUD
49TPuWik9WP5HFpC3EczFxfo1hLjGKLeUvc9TcXWhlEs9sGPR4AWVUTuFUKw4K8Z
Q96VC+8RZot2LWc42Omwlx+temZtGdqdzDUm0N+krbp0AkRNmF8V5tZn//A4pTfv
6qUp0h0WfKb9sXV26i1JoKpc0tc4/WzP7uHpiPLi/+Jbt+ENmNhq1Q1+aB2VsAA1
gxFR1m5/zif3rwdrJyfZI1eZRot4sXYiXSYn5LeIzxQbjjVZnAXnjPMUS1tmvLNU
3cIYkYZuoR+RzeJMSrQj8fknJuFqqC5JlubUthqZ0QjOFdGFAHoAT0DL9NmIbOpb
ZM5dy0PGbEhsY+R2IOVZObQ1DvN/B2JjicYccHahKZknnlWrxnhdztrL67El8ZUh
V1n31PdYbiSHxGqCC14oEeoLvqWcYS+Y61bH4ej4fVNVunxALGfo5T95VV+IkzZ9
c7U1wsUt76Z2IGIeb6BSQV9zteJTq8T1D9Eo0vE8VtwnWK+/z1WUsEQzZaW88685
s1ipCfkD0qFOdjkUqLy+Z5BvrMFTiYIGi2gh0fdj8kA6mjnxjuq4oFPXa77N5AI7
N7QAe+nbWh9jaaswPObGjTMRLFeQBMbk094iaVURVZGetgY0nY6dq5hQjXtVpsux
WbTb/dAOSWZfAsjnhHoRBBigKci9HNBtBpElca7F+/fKW+WCjI9gq9a77/cEyhVY
QdbMCLL1DUL21ZOtPXu0msbOLteGSppdHdYTwLOdVsyXfu4ENCuTI0w4JRWiZVBw
YtLNU4NwpuS0+J0MJ9gmfxsQI8cX2ZLUYxs+PYqbAT69PedQIjBmWVQTySgpz8L0
lkISgTaaq9+2kTbmvEE3nOERhP2n47nKejH7FBks3+gsDu+llCYV7IcHvMVm/tco
lupIs2zooymCRny0lrbpgugzmRD9zbCtzoQMsMF8MDdaZtVd+VvyItnoS2ebPDBo
4hbS4Ri/7oR7+Zf1b2sS2RLx1TxVZDnZu2X5+fJSr7QegxEmq0U89Nl8Jc+oRv6v
DjjpbKR5tZMSWa2QOlM/hS2u+uNykoo6zcHuOpAWS99Khb2jKITm+w/3NqBWT75W
uoM3UvJs7G36FqyfX2T+HS8c/6VNoB1gp309HxxH453Wra2X1NqZn2DvyNfm8r4a
YS26MHkc7+hf6v77wWrGX2nnINWd7F/9vEQ3a131JkAtSHv/6eUFYf9kjnq9qhuU
nRUX7dwYTerRsA8gxyD1kEXHXGu3TGMI8ZT94GdCtU+uzgFgYZN7B2IWi0lTvsL3
OrA+h5sKXKO2a/Ga0xqcCiLfSYgmobLlIX4Ekey2SWRw6zGCAX0Jt2dtkRAHm8kQ
DWrBCOgDjn6+Fri78nQ5hJIbqAsLhhXiXXO5VcUBQ+S1B7mfnXz0kGbwZ2RbPjsR
on0jmtqX7Q8DPIoT2fGCcq+3lwH5y59dbC8FJzWw1WdmE3dBhJGUAX6LlMHNrAY3
wmeK2UMjgLw6ey40fVVnDNkPP6qH04iUuanoB/36Q0SSs4onQssGvPFz2Tav8Fcy
VYon8TWi4mS7P2us0W7x4UQ6IclfQgdPil++JmMpAeO3Y24k7c/W4WD623otbFdE
1d+QzTFrRA/Rfo/GMJEik+fJPwTsM+lFVzfTAyW0vpCxREpivkrnivcasO2+bbnO
Hb8YoalrugOpAOySfOyEsHSTUFKJUA2vd1Y5N2uaXtipcczFxEmBUYYm6e4W7JKB
XcXaHoyk+vfsQkPy3jBQyQfxG6cyF/aMbryI2oosQR9T6zYPuRn/mcpCDwiGgKgE
hwER0BxVb33ZzjY003BhRkHblvCgTEbSUCFOMpSNLXlMJVdd43AJ3a2CUopz9FdX
l0Fho4nVQwMqVo1FxypW3wCn4+zbl8XlpjCFfZq4lIO/iRTSBk56AwgLFl9nv5BF
71j9lgU+WAwLnLi5r+GP7ZZurY9fg9nWQousp7k6jdzenmoyWDCgdB/px+jdjlxv
zvXIi+4DYDNe3XKMAHQQj3cUaqRg0IIUg5ZvljgxdaemXIBLHF8zINnmmwg/I/ds
9bn9M8XlIoZP8zlZAoGSRTjrNhQoxSXPJA9+SMGHDGuKOUPziR7sKhAkyYDLp+LP
LDlhC7klrrJrVT7TehMJ6cFiam/uUagC5hvZvbUS3eitbZo7/amV8dK2vhk15LbZ
oiNlRfhnFwYwEYFZQ8jkydE1CiyfAOwsHl3cSPvtydQ2yyK09KPrn3AbTFHrRIKS
JtxrL5pe7ZRCVIpLuHsC16GcFf9Ih2VDN9SvN4smDopqVBeU1gnejS2shnI2jZEH
ZijYjwlWvaQiKc1M3NpzyVIoy+3cNTKVl+De+rmkKTC4Msi+RHfURLLCGPm0bAXu
sIzUjHr+JfDYvy7MsQKCgalRipptS4tfJh2S6mR/xmMp7SshsOnA0/QhZ4U8VILO
BZ8qBDdCzJSWLbL0/LFl23gk3g117p/8IRX/8BkUK25nYm3RLGfnfQdl7p6AKNGN
Cdf/Uw3sPRfjTQO8YJzSU2BHYyXGzwrTBgJvWXeJNym48sfxnAx+LXGVJA+D2NVX
rNIEOw2gkiE1nqkADYQI+ZF1Zkli1cIAXgypTR/4niypo3MeAtov0OVJnYj8QFVZ
JiTURMEb4K6KrJFwt+muEUJJEEyjFus5oNy0L6LxOpWH/ednBIhCT5K8IOsu8Y+/
E4hJDf11X4w5ozcWDgsuHDZFrW0V64vin1GdmnwUpQQow13w4/IwLcQa+Jq22JRM
ygqAL8WK2dkjK33TwiZNNbhyZpkDbDXWhbgonCUNafoex3QW9sX1e9HBd0SxHwPD
4lnXgGhgGG996BsxjZJL2tz0SMZy9HW7upqg0TqGAIRuHckJk/B4SFQBGdXzPDx9
zVdFeIh1PZdNGFAP//pmst7wthmK37RJYPQ70j7UecHmyqMqlEyv6FChAPQNa68r
vZOZwt53RTAghODM4TNljTHZUIdBMntIVg9eNnLELDc5W0MyVXVc8sT6C/bXdJEQ
HBtTLNQi3mg2ZzyZSgu2yqHZdcfS32sjeBiG8cTe+fxQColKr1TzVnHLkO2XojAf
iZ/7qNXULPmr3XlQaIJBNUbk2TL9XB3dZDKJrPuB5iyZSyLt6PCRWNSDJtS6SExS
YmSHT67FM59vrRkNULE9F0CqLSUh8qWY/XT5sO17/76LElnlskLMsrRqSugcIpiv
G9cs5gYAOTkajO5xA9Ldkx96k9HQyVo3ILWl3P2DEGGKz8sqNPTnINhNN7/J9/+b
HafuEJWDW97QbufMB0Mw8eqOOCJh4UCZk0yl9tSOUuAIcyRss0sdrW8WR30HpL1A
I3UDcI1ZMYy5lVo3By4ED/9FVhrdGsXng0VvRKTENzt0yitKavFE5hDfwIMsfcpc
MVSFSwLSgAuX7puca6a3jBBEgmH0yS84jP8MrFE9PQ65dBEgHpvUMwnxFw74qMix
VkBCwUx6Mr50220JxWFGcCC0C72ghgzpAYswGPc16+tqwJJvRCeem11fCCXHByPI
Vlgj9t4mekPMLWNr//pG7FZyB17qIrz9vIU2ov8DnOKPJKhXuvniI502q2j9+/Zv
6KDaW4wO8eJ5C40ulC42pSmt+YbpViFiOE0gNOi88d7OJAfRubKnDSf8Rlj9aiGd
WeTabNgs2aKFBILoEijTK6MAFQIG8Ezkt9Fhk2JkDmtq98/rQhZ1gLgoPWy7Nwd5
eaDXSRBeik381CLJggxqiwbB9SiU2977Sji3BfMnK7wt10xM4BtvDGKAjje2sbd5
hbmw5xI+IXVTraeCjihhmWX9YqbMQmzZyzRkP94IFarxOysbPKLgZjn/Uni8M6Tf
nxp7DDfoiBsmUbc7Cc78vFIAJtq8UjydL3OcHsRVdIjwNviDn+55AW6cQktplPwO
RL6a5aNBO5jzZ/+25kigbEIWgJzgE5+VpslxGF2h+r23dq8uHN/B6jYR9AwXsdVY
Gh1C+7VF8AWV8/79WXvMDFzo00vH16X1jR561eqydVHvhneMGoY76PodKLlx0orB
5po3RuL/EtX5Lhq3R36yMwk7bNlLOuu0dk20HawiKN1h2nTFmjHeav3HmUMe3fMM
O9uXrwpYHpnBdnwB6sNhe1C0wbqoE7Ya8sCNI+r90G5fN9ND8HYR9XJwZNHFRNGM
+4MmfkXMtSzKkBZaNJKdbtnyggId8n5VScpzn4B8HN8+7Q+jwQcHNwL92vGkh+wS
KAorirtA5ZWpkDFrY4MpPzaCMnvhndVrpjCu6kn9xDk63ZBtb5DohwqJKUfNVQ8l
lS3v5Y3UGRw54NXJV5L1dQqNtRv0PbUsueXN+TWMU/p/KkZKVWkeJoeErHXNpGic
mUcno/+/hH/qrKuFkWI+zdTv8ueJkN950e3Ad+cVOvgC+g8vaUvxkpazUtzn/joz
klOHqUBOQfBvOGkiUmD4HLcinwktwDV/EzInKe+s3Gy5eP2tV61+i/3iqatvubMt
aAI3NFD0aOGuB1ERaJHYAGaouHbTUXNsQCjsUutCTbxUvr5oU/3FgbB3kZbUov1/
fm7fk4zhslt3Vv4ogL6fXPoQsmLzkiVeuIhbxFtVexR28wVNoYolb2ndEuBeSmwS
2887ZMXFzJVSEMdHpIYOV7b+sfjotDhLVdJ9VE6GjzrkDnOrrr0a6fn7Jol4qjND
jiAwM6vy8jy+laJtjoVM0esO7WeQDHHF/cFUuFQ/v1mSLRH2pvucI9o2yDdoI4TW
9WtKEGGDW7RBY1PiIzY+UYhUMHUHKiMYe67mLKpH2bp3B7Q2HIb0gT6UMD4muQMg
k1tH6fuo9eg2Z5+6grOz7m8iPTL1iIViA/rRXk64GEOcJr6GB0QmXw/MN0fCx4kG
m4KZjh5LGgYyebleypM6JW78rOrzkfScT4FXh/LXEoYR6clraFJY0q+/Gj97GnBG
WMi7tHrqY5E7Zar0enESpbekvmQkpt7AxEteHrv8PlyGnA19J8ZYXcZexXBa1LR6
9/Q5srpXsJor/etA0I0NP51cSpUe5qRXUYoQpHad1XrcJrD+LcWlref5rpR0+a+k
Q37MYucqJqerxXMl9JHnN8Ovfhko362U/Ur6o9xnAKcTQXh9/v8SeHcS5iSRa8ky
iutd8avpmt8Wg3s7o9jSJr7oK9Ro3IXCsVSNSBJP6rCt4PmUym7cl9g8d1d+V4lb
5v8YMVmdPTfr6GRTLAuduUmvlfgYZDt9xc0IwzCaFZ2+oH6gBR4zdyHwg8mcO1V5
mnkaQIRKaTmUs6MBnUH3nmVN64v8Cox6ONogKuEnv92D51kWZ8lV4HSbfVYXfnut
T3uIZ1xWyEz3wddfHfUiQHWU577sr4a03dCHzgZbTOXefbYhLPMY05HXzA0w5GlM
3qNRbOXnH8qyWaH7o+V/Xm6xhWVpIdlYc11/ems9cY6an0iWNnawFWDY7KpFb9nn
kjS7XlcGXbIMDjDYYtbcwfxp4ZFORq5KjKaLEagLOcVUaKjqQKs3MDTe3KwZRkVm
4kmsSSWWwSNGPqg3XKhsuAQUpO4b3FVNWEfVopLc333K2uTTnvhvn0rDi9zi9Trq
YIzDBs0wnQYZkzCje8NVltRRx1htLpio+M51ox+1dDkVA/Lc27gya9UAetglGNHH
ppePut3O7NOJsx7UpqsT4QbYGlSiAnlKl2iVK0SvEq87njJj4C5GIiuKoM8I4HIe
VnmNCzBdf3MgGxhSbvbm1n9gCrTupCh8yhoa6W4b7OjiPviqTCp5dBkRuOw5ryAU
6ZpXtV3NE5TQHmtbq3dPeXl6/t8Cfo+2fwjJFQgdwP+ctNSfMqe1vQSNnQz38CPn
78EDFZjj+954vPM7hVVnNi3uxdvmyc+iRBMqNLeYVNirDUstwmeTHGCzq4MQC8cf
seiStJjD2+p+YpfG3qgAl+oB3tRpQdVtnezidJEqtV7Fwy3YgmAQov6hSNsLhcp2
9FzYJJe0YUIES+EVtAv5fO/MRoXRIzBiUHc0iolIkhpN1TT4MhqarrBKcMJTXBsH
0sAvOAkfuzGE5EihoPmlWsLMLyc8tEANvGpBiDmfWXKSGhS8htrFPmZdxKR0PH0h
kye2WoRruWn4HmH+6pfkD8p0wZ0JVDLFe5xNB88mgOdqAE8XRJ2m3Lr5rtPrDuAH
3Ili7em3UflMBr4w6pEN7VH5dwOgd07dej12ukFt4EK6z9LBKESTfUblImtpeazI
qsc4qGY4rAak3qsGJVf6MTbAXODE61xBfMGXVToPWsvEzCACQnMHQrUNfTXFXq/b
0V/EF+WcvoOBRS134BFvg9w7esdhbYJcpESbk9ztfZWB7tzG6eeY3U2xGvV+678N
OVO5Iw2dwlb8S7v3wAfn46tYE1BJiAXsPX1hUAuvBhmf1VAVJeECJXeLHsPs6wzD
WGBQ0D3Lm5v02zLVMR62/d8YRLFlCfnEJyLigYzBMe0PQdMnM0HuAXGwgkt5zmXk
vxtqWwC4+Gs2ddGCwh8we9Z4gSN0T7+xRUHER7yYy4XJcH9Ck1mdXGFMIoiiZZZD
CMammR9v+ElgP9kRJtivQtXJedOsOmhatY1FTMSoRt8EMXgE0Xe9MRw0sQqbxUA9
SQk8p13rt30FPfe63qk33c192xMKwFXJwxxecag6M4ud7L/L+PxoX91hQ/jGCcwf
qZW3kSVluTQH1oxoLWcPik2LTHhBEKD56W3W6JmrZ/egKREFF+VFhhcSkyGYO24b
c/F4O3IKUHnBA8NlQ3tFGtEtuwook8S4TbclOgkGWjq5qH4J/AyE8PtJRMnWXjeZ
4EMsbkDDfcFaNtoo7HvG3TQLqeFbC5lJHTNLBbSGOei85IkqqSolYXZzbTOTRAmT
ymo8QcfZ6yvFQnEZbUY2352K3IGw1IFvjJJN4KywZcZ+gGs6ca9UCpl8Fk8PtYzw
GM52x9dIQfZOaeOO4SavLQfb2cL/q+TAQG5GI8kvL75pJbvQCUKmUezc7h9nnYvc
dh8eD3IySv63oqFMjciLxHAQZIV+cvyWxBssH0krfvcf88yAYQ3bmvTv5xe3LW+K
VLuK2H0/1/a3bVxoFCvxDTaKQz1q1FudPv5Nq15Xts34NPqWoppEnDi0QlEtyDBX
IW9OfFHjq+N0nMRxuwkhrDsQhb2G50KH1Z7QorSflck7ucv77c6y97V4hhCfEiUg
cjIDvBwWhaqhpy5FpPue90g7LUnbpCyeJXLfxbMzc7mu27j8exHRC/RJ4fS11/+2
QxHgTnEV5/8SJJDxpCwf89nYdoW1mCjhDBDc+UGzociVxXAIVHLjBhnqmxRv8MWQ
sJ6CS5OVb5D2NtMx8MlDyoMGVHnpCrHHfkJKZJayNqPKsFB3FwsBw8yuu/E+lzVK
GZg27q3ZyU0t0VXs4Z73Fry3jD/sGLY1dLzXbdO8Sm5WQi1Bq5TqiLNVSA3YS1Si
i9YMt2IbjfOlAcaiWR3U/rJhYHS8HjYOn1co0nmY/QTs/oAELO0fO0/3aevP8sEK
1Hjuf7jemYRXCovWY2OSlPA8rYly8bM91G5QtF/zNtsasRQdzss+qhKqmJj0TJya
WVWUi/pSkiLmGGi+1C1izFzqNxMN9x2yhm1/sj2wI5mr+ORRM8bBeqiIie/HpXp6
vrAKSTolf2ZV24RAFFvEuxuuBo5jYiLbh17upabLMr1ojep6733/h2HHHy8yY66C
f2PHyxPgOCJdRaGwV9dyWGp9z6FzXojQyeTNUkG4TBYfzTBCm6l5LzKGR3ZQzOKX
FEdt3WGr2qdnEFarSpYR3CscC0G9ZSqiRQYF625W6BRMHDixIRZUb06vGH75Z2UI
mg/fOrAPfY9E0jab0+jcbeBYsNX/U/iu/xj3liDs/e76nGiUOk7r8LrenehtmYPC
254vSuDYlxQRDk0e4Nl90mkGBUqTWfG2J9k4ClAgyu3lsBGWFldlgKx3NohF+Fjf
3teVqE+LjZNZ4uIFPRh5JQRG/9obkD9hgHI9GOY2Evh9ELdaXRfiuS6QXJGEbjbP
gBJt7cMtAatydwU2RSBezPGrgqeAyu7IegYyF/FbdneAuNl0E6zTPXAAj/WYDKBf
fBpLF+zm0BK30eDEvQHXimsLr9/vf2N16KoDS8WwEaZSSRBc3Q0ou1JR6fDZP/yL
ro0KJExu3ylkgz1y9+HCett2b/fI5HfP7grGhqP6HvLhf8gXLbxuBDuzhDGAFtSF
JnEUIQwYPDFas3tN8g1S8ZPkw0BWynewQL13V+RoemhfG3cjW9g5l/g4G5h5CbKM
0eK3kky46Jge7OlkQ3aLxQKfNacoPWT0tZrJWPNRt+OAOxD6e8jBAjkewPGo031H
3A3zvg1ClNHKvG1Ks7gAPWcGDiA18Qm6yqWeSc8oF2idXSkgeh/OFyGKtzaGexyK
kHp792uU44AQEPFeH5ovIZKCmnfqKNvqnThKeYMfBjr6v9mlSzshmm6nT80iWNp7
zXQG0FIsjtKheIm9OnrPx/VU7lsFbjoajn3gFjogBhzoVO81TlA+XGinA1sWyGNQ
3k2O0Hj8Or3cnYPdv5/aOYM7IlVd6Ty6jQdRCTyEAdqCR88NGPaGh93Mv/dkZTUt
IfW5wltIFAdzQfZ0rfFVasrLA4OcC/Ql9H5GQ7Cz8YUct9P/wKNZSJRAGTMBWR3N
J2AsExyR3ZY/m5Azj0CMsNXzSiWhZ0L6laSSXomRANC1QnXA8WGEJVIcy2vaUpv8
mZk/U42V4nKNW5rM0TRFsWHsnu7WVcm2Tk96lr6i+Lgn5ujFGqbues0mZPXw/9Jj
OeS+NSh8EYFMQLsM1so5Q7/Hdz6xqwdBRevb7O5sRPfHEwHq4nR+6P5NwjAbwGS3
eLS9LILHb0P21S58yRLF+HfG1UgfNwWGlulqKNb9cXfn5p8avdaylTD/4Q+OiPR4
uB7Xe/W0J7jSVxOoHS/kmL1kim5HqRxvjGO8VrrX23+Q8JQGzqdAdNz1l6APeDig
n91E4ljJAlY9d0pdA58EOARIzt3mBJjalbRm8AUslLzz72Ek9KRSJCPC/pR30bxy
KoK356G1EOGezSP8x1pYyBoAhZTsG56NiPai+z5HrbY58BHMDnapWIvGWKtRlxkN
3QDl+cJeXk+VMHrS0XpEdwAII4SJTJ/WOSVtGfUpbHMe1ITsr+NwbMsEJ1l8aZJw
JDwZRiraqAES15Rp6of3AMphNdMijTi2MEvbu2zv0dyYA4P0BvDX3u1vaRYkoq6W
vXgAq2qfPC5ixf33ATwPnAmivcepTfNWS07sQNQiGPiM8QiLSOIJdSqkKx9b/GF9
WX1zRYDXJz//aQsYHv75UlkekWrtLuKZW9Zl4x4gCBX61j8R2BTRo1Wy923UMkgZ
0FOVHjJCUUgAxLTYpH0C5pl3LTC8qpdON9VtEOXZil1nFkecDCyqDFXBtyQmiFq0
a+h3/tSUQrZZV5laWwgf03itGXWpIg2frw0tgla1CSijd/SK5dpj0IQko17mGpvx
HxXcUnuG9cTgDS08pkqNZZAMB5DMUOoL3QkAJ9IHNyV50NfUFUnkRaVtcEY6wS05
oz4bJqbH8Ix3SrRO/CwSn5CLsDfYSbNV9Uf87bZOeNnZqqeLHjIAsQkcfWb4ztN/
wcBYQBbQB2V43Dw4uhi4zhkmp63+2QVP9zYaRLNCnwLo4KM8XsXAQ1EPSwdQjr/5
t9E1ZVT5yP3UaygEgSeGYufIz9RGIIPSTEqGjimeAwnDR3wKT9futCk0iKovgEur
AAGBl0FlzvBYliNasqGS5Qy9arYQTlSaj6+ACG1gFHSOlveMNnYt9NW9vYsI3ram
6A6lh5RQn6oqwg0LzziVvevt4NJ9TeMJRTkQT4qEuNPsGDuOBA3cIikhw4XuRGAh
5NC3pGxISTaPcYRMO1J+mjhJHjucvZ97ihfmxC3+mlnkHyY7CMvcoBg4ZYMc+lsq
RHngApzNE3Xkw921rYmkyMMXtvW3VfgkBPtbA7RRYitGX5rAQwHOzwPM4lU/mty2
Zd10jo6yKgHjiAivoY2GR8to4sXQBg5csd/2XhigI1xECV6c4yTfZT2AWz/RiTt7
qFioQO6uqOeJshWTc6Uay98aXBVFZim64PvczKKYVT13vW7RVERzfX+kmH8hnGXr
fEmpfJzoDT/9VpzHTS+fA/bPeQeVt/17rgnL8e5WHEypEgsOiFDLkQ/EsGGKNy9R
oYb/z++ju7U5HKMYrQNWbxGqm7g4UYi4Pmwq8kF6IJXJfxd2RrBKZn501K9XRfZo
p4J2sEX00krT/np7sa2J0sl9Y6hoCyjRtiXFDrjvDtGZR6YFYX25u+C6b45Q8xMq
Icu8/P5tzLo3quW2DQ6vZaVmE8swB+sZLVVKjG373C+d+7fCnXjT9bkJbXDnq6bM
Mw9z0NvRRMddjpTyVHYfa9o3LbnNSgNaaCurYUrgIVSBuhBPsCWsW2F6DD2kCE+x
ef9DNuy1+uiOAVETLA4LD+bM9biSKYzmPm/M74ruvJfNn0nH3BsDQIpE0m1Zw+Em
l4kV42kpJ7tEfaIGxUhSw48FQniY4COGPeGs/x+foLJiBARmJzgDMQ/DZ4JLQtIK
Wr28FFb4B5/ofEvgNACIovR95Y4hvohndvC4tpCegTLSX5DDvgD36LOyJYAsOLSz
6KBXBcZWVvEWnz6B3UF2+OsfWTjWommJlhnHaQWC68RYzgP2Mcc4zq5wgvq0oae6
1tGIWCn5sdsa2ROEFTHs+l4jkj1X6TiI5cB/9lczYQKMTOAHlzVHuob7HTukm/3A
XpIOxQiLErQpgZhs/PtwaSbW3aee/SJNuj3Ehlam5hnjkM4s07crrypwamPGCI2D
+HcgIvvinmNMO6Ys7BNuYHRDJN9TpOd8nCEoNPGf1wQQNkJkbfDq0hLhUV7LMJAL
lGY+fFYitXUNjtP7LI2sYZBo+hWaGhNqAe2CBRTptoENNieqYKX7DpS5KNe0HOcT
as3eAMl7N9qUeCKFPVDw7kX8pX/Jrpy2qV9hrbSZGVQozUsxwkJ+ry0wOPBxUw8+
UWsU90+lI9e8564Mstl6CLQPI/gtcU3WkwImTAzvlvHHxRSo4KcNJxe4spn4Trww
9ZWE/M957GeCf8YdPqak0yA7vh5EwyosLPBQnn8J2DETk8Wz0LbwTOXN8G8XkTPl
xBo7j5SiOHuJkoB/V1PsGO+HYVmgCdOE1at7eEgy35ce6W0DF55Cl6JvRbmu06G8
9W4ESAuy37AInrXOgcaW6OfoUxAOz/pfRl0q3NQLOtTBbRSb1RPjrxsJV1xhWH8f
bNUFm1v4EjZQJ7w/nfRkF5vd74nHVT2Yf8I6hr2kBokv3vF/qDqOBKyo5tT6lSTt
wCvsphQ98aCyuFQsfDSpjttrXWUDUqK7WdPL4f11g8rf9GRZ0HRf+IuZQDqCHzbu
tJI3Ct63FrrRLwNJrFm/oudc1AjnWO04Nxl6kuJKl8AJB4dpRPrBxZlqjwjJiJ1g
Y+OeTxAPeWmqNTrbrHHTRRPBvUW5Jo9uv0uXFJBCB8tY3JJxhDtKWgULbuVctWv0
aqOiGPWaz8TD4hon1EzIUawKgt7V6lldkLYUh+Cvgxv89SWdgSGR3A5br83L71f4
k0y/QrweJx9K3CkbAzC+b7s+FHv4WjZ1U59mjVmrSCwAw6Zjb8KxAwDm9Y5QEbjh
CNPSOl2JwESfa3RUAsC4KM+yrRgZCVu4KxLLJarvmjsYrplZnYq1/ODT5/8fhHVS
pUmmkCFXam5FVFC97LOP1unUJo1aetkG7oSv0dOK6CKzhQlV9BRTCsHjwsv0A12w
EUEkoQwE1q379rcFbXvirWUKWm4IRt0sOAl7ThEpY//mmOYzLXTFWjpdEP4CeANE
eWU4DUkAlXzppZMRkMT5Tj0li3pu6f7YQZK3zM17Nxn8EYVngRMF76QzwKYGhFBS
Va5qg8oRHGdMWGG+8+GOESF5mMX3NSG4W1r/eXcExmrGXgMfzLhSihYsw2B0GIMO
fOaF3j1l1XlFkLh+o78YOxzKQA1e0/zk5derppAkuanqmdPWfvSv937oUqCaBOwm
UubJz93bvTOAgp3cZOsVJsNou+vktYNCCp0rULTofVKdAEtWFi4XkoHsLszDYkvu
wCe/c9K0bFBJxCcemGSpxrZ+fZQlO4K9L4Gm6FhyU1y6zIpLodTFCSBKJ9ke0td0
gzvvZfltgzBDlBh0wNCuFbDLI3jex3qq1x5NLRsp767tCZI0zo+RawxZ2VuW9S68
4s/bx+xpIbFSOxkjt1wkba85cmPRWyEG+rlvGmcVCG/3WN5nz6K496qW5KUW90rx
oeutBT5xMox6PsFEIUQ210u/5mvExULemioELT9fb9GtGX3SSZ39DnCyI7j4ir2W
/LjrjioOfCTerMFOcq130cEHjJWnXJxLj5zn8RSBmWNm/OmAAH2FEBL5E+paGTbb
rI7ZXLsx2nsu7w0Y4NnUzmwnJSdayxULUczptqZukQ4cvlBk2V9cXdKBlmAV7YdL
ciDo53WtSPotzeEiTmcdtS5Oma7j2qlYu5KhWSLa33zBz0KuLfimM43T1tM0Qhyl
zNjyV6kHSbPiRBg7IvPWnBuypgEZvLaOd+VDHNxfjAfjCyKttsWxlxk67KKYCWRR
4E6eyB1mm1qEvExXz5+1ZyphP4dihbH33Za1F4x1eq6PwjcwuctNAJ9+7hMXlt9v
+A9SK77teNNd92d6DA5nwrPivEauGx0dPgMNKfBAviKvQ5dOlQkUHYLl6gt13Ffy
D388A9rhf1y9TUfSC1ufIlwkdLh9ZbRwM0hMvRh411IBDCBCqOkYXcYv+ROND4EZ
WyeuPEbodTHj7pwaEkwa4iCLEE5dn1dnsHrP82fS97TDwY/UR3bY6m7GN3yXyhYs
StfeidduhwViHEaKq12++P1dVXpayz7Gi8w7FVv6fqjfOFteR4lcg5pTwFQ5nf51
lqZlxEdIQkw0vY6ovrtFPD0Oj/bTEoLmoATqBZSkDbeTNxIJIzfPAh0wmoxYIBL8
v5KZiC2umXaM58uu87fifJ0sCGRIQZ8uAEHwM0xnTIfYjPjkcQcLR2haW8coehik
QCABxLuPAQFHXVLH2Wia4eNwiVqAm1bLl009rwmWtKXl9aGja5RoE8COyk2CWkuE
dr0xJY4oNCMCGaNOc4vuZVracA+65vnrBfVg0UHiVNsD79tjdRHnr6WJ8D74GMTm
zlF3Z1MSj3TKvTaPxWke9IcFVBp8bRbrypNKA7h422zJakkcGyzWsqkh6YZS861y
dn8wY8sDVekEO2qZdlAulT0O4vzyTb9lhDEpIs6ccJEswyJAdwsEwVZybpAw35YY
nrZunjrHzo/vyoqW+tveRHb/8TwfTL7z1O5EB14mHSSvpONwAWkmxwNDkEledTo7
tq2i+0NezgDabda8aeZGosQoK3FRB3Ik5UzqrMon1ah5nL3+5friBPxkjqeOnI6g
ZusQAGbDwd22OATHsLJOpTzhPrkkWpEVSt1Bc0uFD6iDTk/h+JB9uI/nidE2fN6E
QDo3OID/k8RDWYjZOGZXcThiXJ4dndH9CdJO51i6XqTQsDG0DgPim0u5iaokNi5+
i0rNAYfI5k7bnA4BReEfNHAARYX+/ZvlmAXpdv3O+AQYN7lMeq9AuscsqQP7CSPN
VVKlCtmeYLOKTUeK8OjClnCqzddoGWlRhXLNZPfz0V+yWcrP41UFucFmSJ9gupzD
n/mXL2jQwWymyLeZPP6xFosRtvxT8fuq83Tt05mw7Seh8glYW2ILIXAG3RQxPYAv
tZbYlpaouoU7XmfV9Gf1nu3DjAOOtvFcOQ/qBGhBSlVk1K3D9xxPNbaZ2gL6Ba0F
hC+YkxKuU9EvliU3nXLXa0kHlxnGb8H+KBczYCmcPVnPXZHSOjkkXeSuo6Ia1tsJ
bFNuOYw6eDmSbosBPSKbuadw9tNhAUgd9db/no9r3q7uSLxN+FKqEZSGkEO5WFPh
LUue/1tUMsrnseIjmhAvOGIaIzs9jqzMMAA0DISfgwa0btx1kdYuG6QYhHvujRKd
OkPzDIskU1dAPNqE5gQ1YNEhcXlvpa7O1RNSpOpNRTdcuDHwB3/0uses53xO7A3N
wpZ2tdAsHgTim8NvZw5t7xVXKaz4KJi76HlyUVlZtkANXCx7LGTWXDINnBr1uWvo
94aobpbm2onAT0J4rCTayPj07PNi6DL0jrnXRX7Xny/glPvYqnX4vjPaxNs2QQ08
7evZp4hFBMgOvs7+XJs7ywoKkSpYyVfkJkymwt+lzNbQsveQpVgHdpsOkO7hP4CV
Xg0uOK5k9SFa1J0UGBpAvOWXtY8kO6EAjBl0XEJA+wOsLHxf/KH9MhWYnP1dOkyE
PTKyhpTm/oUeX+MVbsQW0fbey7zCrWf0xYxeC0HiLyd817ougrxGuHSp3zg0khuj
ewwsGMXLwQZvgc1ae0l5yvRAUpkw1tF50SWBGPFgmF0v0k6Yh5uiXRwVs8bDOr52
xfP3XJPIJ6cm5jaL+1eIThY0K7Fs/uqlFlClGwqjpR54MDazWZLp2vkh8aG5JxCh
GM8RHDb84aSkQtToNg+Ej8mNLCNvoCQZgYEoz4BZFovEw2NmbN1OGSMvMbpGJclQ
HvsQ6zknR5blws/+8ik+wriW/aMFujKWN0ozw96CyXVlddQ96YUh3yaU9G7xUIIJ
sh/PlHg/o0KMc9jPqsSkk0trb0SQ8X1W2pUKsbcI226o3EdDaoyRQ99ptNpw5f6z
18fDLN38bxzq81xaJGP497/6VwJcohghxOJWgIbGQdf3ekcXgWp+IugKELVvN9HK
bqf39muGOA6UXBXdaKWSfm6h9AorX2cpf9/PsLgvdkTgxL+emn+LipvHy4GaWzeW
kBIWxZ77A+sik2T6LWLwN8wZjREQOy/bihf13r+Qsz97GclnswYSAAU/gDUUGH2R
SCmQq3+npHGidf022d+ZMxgJ4xcaCgeoZsU/IWujrD/Pb+wjtdAkOdPK+bxNQkrT
5tfuUaK+x9o60qXccUaHgt8Su8+NO/Bxu3tjAozhElQIpv+QwyOJ1FLS/PM67k5y
LPIre/XVWdk1Y+X9kPGn60397AQORxNaJrCLPPNX8unTjtehs+SANNlEwhxBp+XK
jhf9Ti87juJo0yB5VBVWgHNKnSCKhmER5yiAXuutedQkBdB5NRC6YjmE4+HL44At
gz698AdJnenSlGAt2OBkGLBFBUY/GfAEIEAHxJcL5q1KmorKk6YQPvv1IUkkm26N
XpQfbEE1SVEABWye+vH5mCdmJ57BWor7lK+xVQ85AsAphOMj4q8b0pc48LOKhU5h
P8c3NBaP7L2nop/RF4ucd2kIG9gclDqhky/6IvnhpQOzpZmR3MFe4MrM0Tx1GYbv
exImnifcgyD94LEf8q1BLFwwwQwJxYiFIwi9ufGHefr+/HorOQUN/TUUDz/bcTLM
0ylbB/AZVOZKnOr6J9trAXyYWID38d5SwHfD/wFRjsO17VNbTU+qHOxcwkJnH5w8
BR38SrD/YZHMPexSctWIAhqXm3i6qGhgUYTkZHSviDXvrM1L4N5pBpHzttr7VUJP
MhTwdRe0Q/2ppJa0TUNgUu1KxpyyuoDTEjn3OdB1+4HkEVC1X/gmLKdhKuK57Wjc
oAsYc6gbEP70ZnPb/fgt3omBP3WhxUaS93Wao9iwHJhqhKPz61lgZxNFINRDPDcX
HwAbPSbC+MDdimiNu7ABNTPSYrfdRAhwccgtEczxtHq6LItDFZ3aUzu38dTzV6a1
gM173NU7847/JWxQNEwsPZkBdqCjxBLwxaY3XO2zC+d/keg8p7Ka+8YV4h1NrsS/
ygc9FVI4DwylkosuziR5Teq93oMYk0qkI0mp24VbIIt4A5wPcx8ZWcAAAxt2N75x
xCkEWSG2b4lm+u9OuhRYkRt6+4Gr+UOvq/8o7devnxzD1E8K7VJvvRdwVf5AhimD
KESVPzqhvC6Wiac6U2TcyBeRlZ3VGirD0KYzDi6+QoqhbtiwGexRwStjX0qmVq35
2eP8X3Cd67tyG5HFxBBsQJEi7qyj80ExHds8/Ql9dWnUPYlPglDBJnzFKbYfzr7y
IB+taa/B7i1gmG8rEKsen5uNutlXW5QXSAnCBk2PH5vp138Mh3xFlPF/5fw/xVu5
sqCb+rEMgAHglSMkdHDoEIA+Iz93Uwrx/4z3U+H0IDtUi8csb5ITin4CuOfSiKEI
M5xSfViC1aiom9RIytAsQTo2CX6kW8KmR7ChDiIvo7VI9jdjSz/YzhsWgK4AXPKW
VN0gtI6f3xU1XoHi/PnwUAohT9+Qq8rcWQGHjYzxWok5ykwK1HDG8V6TglTlAgxt
5eYi7iP3uXiF0Yn3iAssPbxqpWtYlsYMIAqLNGSL8LrMRZOAqzPmAAmLm89Ju6dw
g5NUn3cSJaiVy2keZUM6KI+7jjhVVXT8yH9po1vF/qp41BILlrslgLzilBKXPxfb
LHL+AGbIVqRrfgvtIA2prPGvJ/2Hr+lCa9jyZZFLoP+RuGLw+/xcoGqvw0DKI+ko
4Js5Igi6rkfccMs+300gBoGDP5h/ZMKoIao73YJKk/v8kY1iB2agXTXJgq0dx2bE
/il/W4txVfeUi2tY8zwK+H2O2j8y3kd3gZwiqbtB0Zn5xNk3SMzBiX26/1UL27vA
pWVk2HMYsMZRkcf011mtP0S7pfKbs4xCGrl7XWx+wRNWGA2CqqU8ZqeP/hT3g2kD
6svd0gSQbpI8FOsJRe2tyFow316h4EKK3ddNr32CRbGAhh9rk95SZYqAyrH6HEgm
a0FsyEhcgThX01jvk7xMBpQhqgXMQ//BbHpLWlnCQTyJHnvGnSLPgjJ0KsDF2lmL
43vQSz4Dms3b37QWI8VEhakEd1TYgn4PPXUT9IBXk8loaue06yrVtmve9UjZLTBE
Q5phTliy5A9N2nSB9dHYSv4+RN/wj/J8+DoQmYHcnV/a02GFm8AcGL8Yvu1Iry/s
5afU+OeVxGpEIjCiBCoxReNaR5wFtJ30wFhi6Sh3UoaK2XYCGfrt01HB85rA3Fdn
qztVOYkEetnsemHvilDCYAPDBnMOnsnNYDTU7SduYX8VRtYbqfWV6esVt1tlZT/A
gMqwSCOfoZvLN6QckhaNRYIPJDWIWrtTzjevi3+jTmgIEU/WDmld+E6Qxep6NxVs
ouVeX2MAjVz0JY5q6WUuvBGYaMD2HkSgpQSD59yWstZ9w1Esj/xy55lbHJych4Sf
/gZHc0nhff8rH8BMnEjiTzlMTSapUttbBbvCsXrt9juY5B6Oxr/qaaUSbALgsZB7
Aqcx11u0MJuUNdzWepNf+PjqiTpA9aDf7N2gbinihlRu/dEP3cb9Mr05tctUmuWZ
y+rb7SvcIh3zaxlg2UOkg1z7VGnk7Xk02ih8QHQDINYQ+gaTKEJISyppONXFiN3I
UfOUpczEHsuh87cxGsKW25va1NUmvxe3zQTy5X0eptx/+OKR85I31ylERqU3pwVl
9JgdrJMtZNn4szmPnkbv22l4T7wp++0Ltwj19AtcEHmeSGW6FrtCb1bKHvEtZ7Qr
FoCXGnpNoVAmE03FTWDsXECzazA/DMpVLaIWsanbH+lY14ycJ7rM/uJ+yeiH5p1/
7uhg8MBrdcSkxC8aBI2ebnH4z6fapYc+1C2FeeRgWGq+k6JmKJX9gfiLH2SxfnGO
OucTe1cKeV04GkRyhMF6p2/+vDO9eJYoagQBl5gDFZhp9XVxEtPBOcAjrbNNndqB
4A+gOecdMOylNwu1fEFcJYEnydPDHdXqab5Mhxte29EVzVgxIRF7yv4xBNjyhqWs
8VNB2qCDBUCcEFmPiWAoCdvpypKJhcIGLePHDLMGk3hEv5yfH411XW/zCa1ff4bi
SpwEfacASbvu9zEiHfz0f1gNICE0QT93vDIfKwui0N73lA65R8Ejvp5d/3RtHP5J
8haCqqFWsIb37VpiHvkpxyrqL48NOC1cyiYs9jLTQX1NQ0uHGTuWlliI/wlGErBa
SynbbJAq4jYiAqsSTotGAp5XUtQlI8QiHU8gX2bt+jJmjZozKYUbiFYUcKqrTb/9
1H3a1+Q5oFVf0ccFMQ5K2AUMOYkwJNYrHFYBjzeb2hdb6VdBt3hjSEMGtm0Qe5Tn
GDkCgRGEE/4O08K2fufveMUHMsu7MHOSwqGboMI8xjO61qOQN3+hpq0ARl2gt8IA
XDgjcq6xVRIuModhud3fBIb49uwhtCcAFlEzYebKNxNI9bMQeQ/A4M9Da2sfyaEu
fKKa2i7pjwqv/GbJlEI+aD2Bc0kudaoS+qfiZybJRo2/MlQ21HdMP9VE5gfbbzDt
TnyA84DiFlWYaOJT7e0/i/7gr1r8GZijuHoSFre6q3y2P3h9OQZvCznG8/WryV7g
wlnC7omXyqgg2AWVrNT7cyZcevnPMC9R1NrrqxLZvcm9BQFLnEKCmSQEqGtUxuYh
Z/V/YhggxWn/s5pneYz77/pDTV8aqscflFeTGO5HU6zOoCzT6EeRigr7/Pr6PGvB
gn+9U4c8b7MmV/Jo9QSRtEOlioyhz8qovJ2c2XsOccxwGUkhI0VeWQ+caoHzKv2M
e/gPMj07alFsEtbhCY6oL7xj8hqkH8NnHfzcr6rcJCNzTUrtBbhhAE3SWMDMh44R
tBzndkoVauciloKPO5Mh5IBtincqhhERgFfaj9WISJZ9iBTJva7O6YPXNRCxM1DX
EG88MpsUcj0kecpEXVnYCr1x/OWdJ59kuhPt2xOwZ9djAdRzJ2rB6PMHchHtDWH4
gYyw4tgEEWgoEHtWFC9uesI4lfI+lY/WE6g5uZDd/U0lkA4etzoDA9RKfLEzJr3u
TEr48FTOwc9skztZNCq5dos6+1T1FTQgjuEustu8ju/dJdt9BLNyUmDC8rQw8o83
vyjtfLnQsW0IBzuakA8Qt42ESi1vpmL6oqV1/nXcrwkZNFif2jCFXeiRTTVN/JW0
DedtkByWr3PwsA5dph8TjIpOAJ0alFkUrKA4FTZImMg1Adx6Dv5KM/pNkyhOXk7/
dT8MfLwNZZjA3Snlr6ZoIQmRxKO/WGPd6zAS6LT0b7La/3StrdEeOOsR2QdigXt4
JPvVpwfby7MZOBeAe4GYv9QRtEZr+PuvOzOw1/QgdXMkJJUOX7/0GR+ycdmEpwIQ
R1MLYpEHOSwUW+MuDFd0SiyMR2r5JR2GF/b8qSjiXJA2h6mnY38ZSqUf2NmB4kjB
SiSbQqllTMP9JW7NwLl594AWHsQBeZdzkRsQgMMK9mM0Hd2EEGR762p+YHl9w13P
vFNQN/WlKKOcNPhAgKP12HAgX8QGhNjaOIk5JgaMArbmKEuH8lerzLBPBwW5B8/G
QaTHldwr+UYXA9YWoXXfxMVnHxc1UPAENlaA8HLkor9ihWr3fPOuOfTij/YycZbH
1tcGlkWiyQQYkRyKNBgL7hETUkt874haFJmaVw78qiTzuDU796rahgvSwXVkmOX5
+AlDP1V61q9B0aDKNWo9z1MmQK+n//mAGLV6/XuDcpa7LFpVyLwiaCYsdbTEJEdc
KMHfiB/NVUaYtQYWF3o/FEylSWs1rQ05E1mfQUm+ziJIU5we5mi6BaEBpGc4cUJa
r7pTY2TV/KVzVdLdrQBumfv4Jsbd5bURr5N7NphBrId5IY+MeZ9vs70Tz6TguwjL
`pragma protect end_protected
