// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rhUHbMrWtyHjF1V+ygP8StDV79OH6ZccfudG4Q4wIaN7/CVlKG7JPkbw4IoNgDaE
wx0iaVgK3SL+qQ+U5gg8HfzZHGXuNKDzYpN8f2RGDOjDZFwr7ly62urrPYHjdCfg
Qh8urlokCwZc5ag5nA+1oWIq/IpbYIoWwnc0x3JOPGY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 59184)
tCtQxtClr4Imh9fP6vi2/JEaXh7BWetExmmPfswlzTUo+NFGXPvZ7jc2jnn2C0mB
oFkTtI/oxIGEX2wqlxtFc/so2claTIcw50clH3zVezoyStE9sAhb4GmtHVDq98sq
+IYCeWBEyiKh6yMMPU+wnmBnshqVf7CeDFBOvA1l+3rC3yWXbtNmvlWt5Uv9uHBd
bYXvVca4hiN+VTrzpB9mU/8IbwyC7x+BFs16fXD/KqJCFL6hwo6d66XUsXL5pdeH
OxSiqimik0UtzkDgEFGRqMVswP7FzWR3RlAQ7TyHh77JOK8t698JjwmX2HCDmob3
ytcNkYxLJbVRFEPcq/FaWEtKsBjKke75f3mofFi0YfN3uAEr/dfQFpsMAlrLpkfH
VihxoSwIVq/7QmwbfRv0StrjUnqIqBecOnMOXYndRLpW2OeUvhDJiJL0qfav89fv
Wt0p6QEQKYjhQy7fIuaN/zExDCmxhapxeol0FtSViae7RgWyLK8ObYKTBaFWmWDH
h2dP35cKo3tEh4OfGeovg7LapTkkIMKvEJxKaW3+7A3/9qy17V9S+ioSNfD6z0Gz
5SAHMJ1QLOZWS+pTH4K83XnnHjZ+ZUhovLvq1B9VjQlGivlguoWsFBiDU/C1KNst
UmYLpIXgc7yB/tJbNEgs8/W+dNDE9gYeRihmf49ycM2tmAXNL7FFFQHyrNx9Og2b
NVkzQe6yjN7rGMt8tUJNi4xE2h9pQ/JyBkmlv7pjmVX5nESJESHSHGvD0SZz2QWa
UiRqwCmcZ2MSB44ICaJ9mr6750yKLCBh4pv2uEnWtlD+1v9YVGzJoqGxBHUaZPgt
NTaSgwkm7HJFBwof0ChxyYvVOhSlS+fxL3JbzRvboX7rwJYx5k1FyxgDtL/EhiJK
9Lt/0aSupgJ+iTbUGUI7x9iJ2Lidtq95xHxCaWmRoqS1Z66nggoJAUY8JaHRy8yI
v8FdmfMg1YqEE1Waab28s7CFudPUI2aOr6Meg1HWA1QAvmGkjB4yrkuCVD0wdqZo
QXSQDKUPEZWsh+f+Km0oe+hezq2FaMqGgdpCA4sdPxPQlAMRgIn40u7+9Cpbfrxa
vguR/DQMHOJaBKs4efViSwLPVcfHQ/YY0oy9g0wntrAS7aDmQL8LsD4LPJiu8J8B
Jut18fE0K+C3iHMjQiRE/YE+X1NcBshguwmT6JEJ4FVLdalJpMvyyuh7SZasR1PA
g4yWz5KBUDo0hW1MMGA3L9REesX9H9qKERKL+q1ZpCDap/R4XBCUICmXgbMcfgog
I1U/ShPA2bAUlTDwhVolSiqbrKQ8LN6fvj8S5Cwh1SNfx3MMOxVKpyZS1M0YaeLC
GbEt9TlTicmSpTCmBMzMuykQ+oNnIQnoJWIszQ1zoepEzOhYNlqI9DJfbzbLxUqu
JawPw2KQJC4anAyjljDOT86ApyrypwvumPfngqimAwlKe8KLzd8bq+pKCsTDODfO
HMdzg30KyRNR8D5aMoOWbIGFolQH8T/BaMGWSItPvH69tXKJV7+1C1cbJwsGTK7R
ZtIjWsgbHiRe7VJa5FxGjZ4MerXKgiYZ1DKnANxNa8luu40ElMXSW6TSExY2S+MZ
d7PXGhku7aqUR2m9v8w+R0FLZ8kbmyn/nM+ZQQSeLjkAxgIOonFtJLehG7DWMchV
z55UMCSAuVd7oLYY1qwtI+2Xd1ILg1YlzZXelaAe3qSqVlIbq0371Z5H+5aiUW7a
kLKtVx3XWukSX8SQRTlpEJOh67ArwbcHxnhEwDJ/TXO5lUVsuimkMD27fCrOvgZ4
q9azxcgWS/TlONlRWGeZA2tH8sl2xklDhVMZl3nbI7DQSI28By6Fgai6XWkefdSZ
88RSAxFZ8sIVEk1XO259+1Nb5r2mjZExq5pe3DQcRmg+ZaX+3Jz8dnGf82ZTreDx
1cNUfTMJtyNo5RaL3+6P6nvI+wtp5cLoe+McnrqtTCh8sV0JdvLBZ4Zu3xlB7P/B
RTXpbupjcS8jxe6m/gn8i6r5S7BGRBD7jBP+fMQ+455x+1YnTDryDNRcLnt58atS
pkA3skg8qie3MaI6HNqX2mDPdjLSt2brvwGrm4YKHGCkYcoXgWZw1TYOeOcYawx9
gUQEi0impnotE0v+kMSDj+5Y8X7EQvNF21XtdIi8f7J1GCVPSAFbf9LjOaByYKKE
ofHfE/OTE87yfeiLQmG5npEMj3wH594BZ/7UVRclazrKYBL6aZDnSPIeEZU5vXLq
kU+BbOtjgZtpE5h+FWQS5Difpms6jxg9CJAVbNzEPcO1gZuoRGHXSKUfUZ0YGUiu
dlENK/+TcJERrDAaxtXlTcE5I1jyRoDZfSimYOjEOHkUe1l8GH/X1Dhi4RwglSKi
PFKA1Qad7I/gAu8hmILqXYjK4dR8acjmaJ2VVnrsQwXRyeWrRugkcDmMuKTmDoDE
42p5YEDsSzgomK6R00RL4IbjokLAjMa2I8dAQMMP1jVEzVQsNt9nrY5FJuATTtX4
6cWwQsxnCJbJ+Xt8CIuvJMJOa7cd0nhTUrAu404NNwahkS71eu8BDS52tJzrAxqe
iVmQRGgGkda1IC65w60HwRriErETb1ahnmQtEGWnCsunKgy5FWCbXTlRajrpbgZu
zvDntUvGtUNUw44doJxq+dQwdL0Wlyyq+iIpmwO9u2x7xr5rmwX81BDMMOLBxxm4
Q0qFcAokhQSFL+1TU4PCYTrp99NbO4CHtwFDDj93GHz6WELfccbN/RxdhKeQ7cxB
EyBYu3weLk6d2ooosMY9G65VmNC1HDV9mgk6u0GlUviZ2DJZaZfpwgXXhDOLIJHC
GSzUvaInM0NU4aVeuBvEw8jUnMAUxYRv14ebWFRhJ1mwBTnJztdyV7PuVsRCL7Ia
EOFzyaW5O10Y3p9SgMNDmo3Ii4r6/Zq6KyirX5a09Cb8WyKXmpBi59ZGF6DiwlvA
E6EQ98502QJYhxS0KjiVv9wXaqxprARPWLfB/3MCT7gvifC9QvNRgRBB8Sm2DRa2
HXGP9zocDk/VsiPFj5LWhq7czEolJ1lYKxMXEr61UtJP4PJqs5o0yQqKuw2lo69f
rnp+X4Ry0ypla6vt8rltyGAKy/aQHhtsZOr6n5XCsPVg0hmFJ8co6oIkDsmXRtSo
M/KJ2FCrAXuJcnUpT525O/DbpFIQSfLl5QHwKz01IDgKrStqbd/yZ/ukL3QS+toB
A7SS+33tZXBfmT2gH91yUI1RzrZIpGynvfTgJ5rn++TlK6DMMi9hGezcmlvky7ii
8/DyP6NDkR7YZEAwW13ENWMgZo9TAn2Wl3gbUkrKdh6kM17x4nsaYOxbinScoM3Z
rfxRIU1TGavlf9aAAL9XDyB6/xtOoQc74KYWdBjLCaVArKiFMVGZTgumE+6Eidgb
rT1vFOq8RiUedc4sPcwCcmreih+tdxDNBr83MvAOZcOCr391XWcJY7rE5JtzvzZf
KlyHIFQ/3zVVzHh3BU+LyLOyhJHWB0r23KTIL67lYyzA0DEe+x0Fn6JQp7Bq4q0v
EOP4GwkLJdQyTAVZntdMeO3MDeOFbS2P32o8bRxrY9hTL2USXpuFwrLBhtNE4ngP
n6BL48Wyv6/jzjEpn/D3sj3H+QXgyDE7g7niUOGOS+WSoaJkpsUgUuV4X5l+8X/4
Md4h191q3XIkRQ9FpwZ1IlonnCRA6flfEm0Vi1ZmX6ARNrpwKM8cXAqOjIUWuU7z
vQ6hKfgrqRAiQya303NJK291qD32oy+xAcaHHaDRljN2N+zt80Fk3/RZd3Xu8zvG
YbrEmCvk9z0CfH1/NVdc9OAhDy/ne0458Y2ELOZGs0QdNe/Yjd+BRZ/EhrYImFB1
3Z3Tjx9+RYteRug6pPQYxA402R881OShxEAvQXji90B0LlmTrzKMKSL8yVq7Vp6e
B5rbHo3yPB5+mbFzyf7TNlXNTUNuRezbEbg03E39zW3hgOssCPtDuzzPkEys1upS
HA2mFozZgYikCPshw8k0Wokqlv+DFbwL+vT0uFlGEaRcHuyT19G6RMp7Wn/isfum
MRIz6QFh/zXJCl/oSv9pemDZzWJp9eSdQNL/Rm1jTMXcWeZcgm4TMMoE8E8KUnw8
MYJeHyAi/aQgGO0XSrmglvUTyCJfgbOmV9aJZC01EzJTVf3dGoeSUNeaWOTCxvhq
q+jceFzzHIDVzWuLhrzVv3sANVtFGalWV4L97Bp2+thgaN7VgheP2h2twGV6yNa6
hBXcCo1lJrSTmK/B8d3zq43g5qFhiprKLCJP4YFSf/7B/88dX7LS3kyenv6fbLUb
1ndA9EIb4B+jjTth9e25haCugVq6PHNkFoe4FbGYX35QW949Qn8yY12z2cu7O+XA
IO3ki1NdqwqdhVwCdEqdWF80iZs7pX+81u51YpzmlO8ucspHYj5d7342w1MrwkYJ
ZcvvErVrGKU6tGQJ6VMbJX2M3U08Qee10F0MNEQuWyOpVCkvd0js4sqrDeh9Qpe/
aNQGOYAqM9tXsbKQzwFOhk3dZhiXcBoJYHNiLHKnnMGZd7DQUcc//UkUCKtgIHTt
rncaTUhumTJhPyZBz8ltjHQxEX5RaYv+O+7A4UyewnHQZOautmvYazUJXcIwKHPy
IvpI11rcxyPczb0u5KSwT1pgG1tk9wMt4fiXJ1cS9GjxOPXuNdAC5EdmyiOIdkME
1i6uYQFwPLQLEsOFXQUSBKlxIu8RwYt9u41PHHWhHTRo7S06rVhXJY4WZwF56tmC
w+p9GUNqyvAggk+iVU+7q5MfY+DNpMIP1cdNv2Kp2opzKw6/xHqEQYZNdZQqV0UQ
q3TNEzM6J8iLyZF7Ufe73gbKzz8rRLXvIKzc2B3h6m7Od1AZSMeFjE4v/BVfN3RU
4HHA1mSK1CFlJmXEhysaCcQpKEXF0mBwFY2llYiKKF5+CjkRk8CMb/8lVELcF3x9
Vv75p6v98QAw96KNMLdlG/wVuwLhWn+M3WWlRjyfo1E/8cJyPkx47zR528dDaCfJ
u9CycmCgt+OJjOxTB+eTQz5BwyQwK4yZzLqEzcivEtz0W4CoKrxgjp4ghzVXgxEP
VJCU2/nq5KR1PbXkRdKomIXVGKa5gxO6+9kIMVqo+uBhpktMhV9n5yUgrnO2DQMw
dHsI+/r7BjU3/CsZdCn4mabWjoGc1RPwve2iggTS3U1LaRjYzBUrfz+BQMDagZ0H
Wrg5MeBJOMYYoq0izPW1GQNNHu4LKl+4iwMH+x/yQV/8OQs9snZ4LbF+7XVadfNy
K0W504st40crHTLc5sduhuRkrGN6nTWn7QlAfBGHBa06GUzr4a0E7YwHA1VFgz5Y
JFwchP9FvbFN+J0DE2YBpFfElIQ99SCU2pSmV71Ryx+CMiUN2Tq1toSciuEBLTP2
Ks9lragl7XogkLIpGnOAU6srFr+SwhX0Sx7PViZ6cUZ5kWOhxdMyn+/x249ZdE+8
mKfw1imOKSKKlVi813tMInxsfpVcMXVoFPXA0y8rKHGhF6P8VH+x7zYF12mHbN2o
6PZWMVxwjgJEFel7OrH80fzYOmlSLA/Qy6+lyK+jScHJNn2fdeSzTOLLtTtbd1I3
GEJ/F7fNWzKq9MeNP8Y0s7SiePSfXWmYZo4m7awqpJ7iBTMnKPvpPaz32uJVs8d7
S6M5tfFbbYgPFgBlqLQbq+DOwV2bjnjEZt0nT/QwwaqkEa/FO4jdUYhc48P2Me5H
8SZ0wD+9WbDHXtEiiG6IBVeIn2ow6biqALOhLQz3zxJgXDm2/w3giWYwgk2KNaP2
oUZchFn1Ib/FTO2x9+z66zmP0XShwYI7szwcZmIuOeeDJtzAQ98g6KIexeAa8caS
VXlHAwCfbZQiOjB6LkboJAOd2UYZFJ1D9POpuHeglquR+DaLLIqNj54oLIjLYFsU
Z0sEHib8KnrVGvisLaGyQmv4aBOvY7sHXPlTQU7lp127U7rGL0uQgABWiEMzIalH
RMSQ1NCxhOLsgyQ7N1I3HsKvlQivz4kTncG6Qd4wCWb2zOdX8DDkRl7YjHFiPoNW
/8RFH936ZiLJY97aFWnHJSA2QO3F8x28TKei0kn1WDlAFCmMoLj680HJ2gLMdHJB
89wCL9+5q+Xq5EgDHAPjfroyARIfMPr5YGcDQxMKMVtUhENNrU8q1AwYMDmNFBTe
79YgApGfxzZCoUfAn+2Mpyq779PV270wMDEZoUoCAoo7/Xqk1foFr7LSuQNQZHGi
NPSGCVzokhri56aqZJ83AGX3iPtLhsAr+Wr9o/R+8q2gMNVm07Le0d/efVOuiEoA
dm2gv5OIpIJ//B14ZqStaOYR8H/AIyG1Hd/CEJWRcHWfmH+4bSmPUMmxrCq92l1g
Xjcc/XpvrRgPqoZGGT5JYGeyP8Itr0vNoThYnhgROdOyddXgzA5VGHl/kQpNkNzp
2h6UD27Nc0+BYG3ruysHujvf93m3KKeB0Mf9LxjW7+6Xlyyyz00DNULU6HWUDfpv
J24XdHhetz7kzgppquKCCzh3I1t2MQlL/dzk1Ki+PnFn/Rdl8IL1HYPRm7R+y4AY
0f9xlPA6X/e61pDcBVyjhc86mI+e3V9Z9YD73kSUDpQ/cmvfiTTogJo6hnsep4tJ
7ZFawL+j3kqRLsnm9k88v9zXRHc+cf+6XS1hyTRlpGbNMJPesl9JE7JVUl33wqIF
Z+qSBjQWctX+taUkxKeZjxb5zZW3IxWBddg/eUhL52/EzKQGSwqCJAcl2WzT5pJR
MaBZUlNtI5aesZZpBkPh3aciniJ49vS/xvMdF5m/ybbor1sCEgaYvb7FuOFQhgCh
rT4XWk/HBdGNawe4BDZxVGowfrH7CpV147oFm5x0h8qd5TFEt/mwMGpdlKU2tXKs
Y0RT2TkFpsjYZiwuxdyrJeeMr2EdfvfJMbiX9K51to0JzaMeOHI5uMUfo3Dikzg8
q/IZLEf9hnv+bkMWuxZDBs67O0dwCKwNWpbJhtwI66Eq0X7SpI36aQnMKKvS4tH5
rtwm+bYXXM7FKvPX3lsOKdhY8vXr5+6K9VafXQxz5EY8YRuKb0Q8f/sATXlmx/OG
n8rHtatIo/r3G7xyLR6hXRTJcAeKuMIaBX1V+ImI6jEUbKwxH/dTyJcxUbOlnAqv
8zppjnePN4xmuNBuhT2KfiP7Yng+YsgzeXXpdCArKi92VIdg/AtmJcD1FRkIjE4m
dwqqQyTkfin/wCHvZ8eI79uV2qovqXVovBsoDfuqZ20whVyZbMlmeFDpsYaTOdgZ
uilHWyMjIrAc+NH13pLBiPtXqw9/oDo50k7kbSvltBew5nNbDOjlh5yhLvLSNmKh
FEtyzPlxth+GSrvovug9f/hUAdo4O+MbIFkP1UNoR1+a2uuAegIdE16ElEvI53MT
p8Th999CHz0I8AM+k/POde/v4hLuPb6FWhwC0r3jlmuhtiGWtX4ClxS4Z3CegeCB
3jwt36SbsTxCT5n/PFFLArCPYsyBlBaveapL9/ozfXMlnrdyt5/zbDVMiQL7jvGm
Z+Lg40S3bY39YtysJl7aOc31d2u7pkYyC2RbChEr7g08OO6vwCnBA/VF3vgf47l3
oKBoZrURR5cXOKKzKOvgdkc3EWMBDrCyDnDVqnt7+VOHk52CVHkoWTOsHLQEEpba
ssFByIoiQYXxIUltvfPkjoH4rPBK7/cRdf++2zVrzgtcGZzKNsUDaNGFwYbiyaBZ
ZNSOzFPf9OoTXjzhfPbJjZ2Pe3FMfyoUsPdPEtyghglngq7SweljD+wSu4R80Ztw
jTY6qBOc3SbfRJKzkNWfZSjhgrPRDw9048kujlwi8gYv2WwqjhcOdTwA92Mo8IVu
VXY2FrNtXN9DtMoQIFuCPuFOUa9Tzbo6jvjDjOC7YOhjTF5r4sGnVePVnbhjDbyV
y4OpA3c6S1aFM5v/sDzJdxrlNc4aOA8lCv6U92xJ6zleZkOhftrDqNCW4D/AbWG1
WcGEKRc9VmSRdT9WdTUXPe07jzr5qkaOyMw/SnbDmbJp6dBO7jWVMF+8xhHjJAsb
+r/yonh16NqiyfQqgylnSUsFwdqQJqsKzA8sPTnhHgZCBqxjj6fYd+y1BcPYcAp/
FqHHchSZ3EmHRqCZdSFJVaYWY6VXzkr89rP9mzIatxA8N8Hq8V5vatxYs7kPZIK8
arGRQbrGovxJKb/lpMokz8Lo0DSYfUDTFiaCnFKCZm4AAMCbpImUYaHJnfcVVpsz
kT/DrLmEUg11TN8rGzT7LkyF/2gwzO25VduW4TjsqrEMfyfSP2qBLSDvSOcC1ker
KrULHByckJCS3sAMdkuO2hMIKbL+dzFKD5jYVNKobKa7tLeq4RVxJDQ5WTdhwyRv
s39ANoIzOAOzAG6JFNbIsfF5Z0VHzQ2xGcbBwCrUCLHAhw2ifb6M8RsNBmlE253J
qsRayfysLkVZMMlIRRpdNnn7iQdpgJCjp4l+AowOKWPs3a+04ZrvJdBWdx0JrkoO
B7lCT9am0czFqbBOYmPmfyv7k+/Qul8dTKWdg5sKMMqoImUY6ii2Kk+ydl1MlhnC
K0CJ9oPBxWoXBfEOp4OQUP5g14H/Rwze8oyh2zmST0EYg1VVlLbXo6cVnoB2Daxr
oWaBXvjKSA+I/qF9PeoBiOqNJn7KbqzPl3FWrxPzGS6SCrtuQuPQIOmVoa5DTEmV
swP4Kf9bBcWzwrYV82CHlQ3TA8l544o5AHTO99ybdwmx1qsIheh/cVfqO3q15qOY
uL0Q6wXWn4H1dQh3jYHpBzatouh59XCfcCtBB/6TjE3MEB7GZagJH30aK1De8VRX
0PuDIt753DrmhyYK3fspllPcI7Yx3eYkziIrMszxdjgVE3FOzMNz8eVhXe6Pvs1T
RjmkuSTmBAmvvLSP78AnQTSMh09D2av3f0Ct93qDO8EnuhSFp67oP9e4ODg5WhKD
qjTescd5MMLTjLbs2wHTZNPaboqqgkqZdXa0rJSNjL8rBIKkqs4QgNbFnuUtehJ7
AWFd1x+pBQa0oWzLrdgvjrClV9nuoNOZ7A+XlZDsTMymssDbAraQ6oH6MtkzJhIJ
EuvYxFFB/+z7Wjyc9r8+XNCzLJuzkpMBmdHXOL6XtwSqnLfcx0SdqG/AyH89bRx0
nLI/yHke0gs4GbXzx2v+0g9wmUErZ5S9NHW7mqjEMy3kJ2GeEt7mXydsjFm2QcHB
+ZURcjXaQDhil7R0MInCUEzjz0/Rdr4n7pqey3sLUiBYS8PEaoiSjuQQSvxjIhB1
zCNZLDxA06uluCLQaAHUd6LNwuu3Qd7zo37XIDg5VMrvF1/c7Di28Zl3hog0qFg7
zpe/j+Q25MQfjqyLHruHzJLxLWxvf/sktpuz9pP0wh3BFMmGZSXWIZpwR1RWT1MR
ePtrbMvasOFsGvTzVblu+3FmtqUYzn2pZOOSm5MWaMOrGrX549rSUv7zyUhImyxT
wLDBLDY/mmYfytyg/GQJZnjbm/BROf5qbMoMuSiayePyILCH3Lm/+tvNUg6P/8R/
Z6A4fzldbZhxjA7tj2lgJnknk2BHzOZbiyfeXU/4V/pr+5p1OleLOwqtD1jlgj3D
DLuBqpr/nR6Jua6MDFj93p1Sb9GcDNkCb33steSnNd7baJp395JK5auGh5jwnv7e
0g064A6rHQaNkApO8aN6U7a9fUGopMJZqXcy5JkuwXvH36VWhgSeRHUEjRhBo1YE
m+c/29emmbR65/cKrsAEYeQ2qn0l9tm+hPlBVfJZbqHqhIoBeGSdnj7JILr0LksV
c+cD1xHpAA9xoG394vPcjQ16lSCo5AzXtZLsTxF7mBhIovw6qHKJF4NX0xo1rSpK
v+FfHGC3na4o41z4UQvPu8g+WQF79rpK1hGOqAQNkFujszFzmR5pClwl9PiNIDE+
DvIJlkmQqZlbBVpKB5JdEJaUCvQRjiYxvVTnWQh/a9TcMAKrxWYSZG58Eq5bPjRg
74+SR36Dt+h9xBTem8h3VDZib8xcNY/77Eg/X1NhvmdSSaTViVha3SzFO2CscQ+E
V/A1S1v1rpi/EGLeh2bkso1r3/Z1uDXhpQLLMirvpiLwZn1e5ydLaIhZZ9AyzQdq
pwWjFNcGYsidTmtSeIMfCqtMxvcX7p6hWGYpP6mkhs/kzqa/BcGH2ozBJz45xCYK
SHRbDzJFXTJDt/Uqj4G2o/N2ZeIGlpBAfJHlu5UfWsmdu1x/fVx7mFs5IHLHRUHK
VewAE/wUYryPb84gY6XTRkXkXPzzOp/U0jH99zj6b8ctL6Zq6H1AsYAHlBlcEJyI
ZbUwZNgfaWBBPBc2e4yZ9xQ23lkD8U07a/uwd5ZnFbFWRvw654HMc41tfxir5IGg
c3pOlBWEruNZG2iHRb5zwhSLr/HTos2EmDGPlvQLPGbp314FMf2w0RgAWWTHEeOQ
Fz3tP6hf5Nepze1kiW8pKGMekrMkREWqVLQNqbPC7jbHmJ8dnsvny9tE7XAx3+1P
Q2VkmLjuEzLTqb3ahOco4cNYOmxwLuCJHBX7B2Ijt7Gw2fM8zHoxaas2plhBwe4m
FGCWabdFpL2jC9/SrBVpqxO4nIwRV9TfB8OLkkGdhVpGUZnvZUA1FicdWQNjj4a0
VX9bpe3x2ioWY1hHqdFcUhElGkm+GqtntG4xnXH3nW2/JzIfMy/+6Ydds5OD9/rV
enLbsroNHsvN6mTVvalhn/vURLA7g2XKujkwh2NaIpR9pjyTympTNH1716xsdUST
NY6wt43NwWuCEy99V0oJF5OsqyUtyyaAU+25UG3Tfu71+YlUOcYMsVGR7JIGuc+S
NTwNT62FESvIpOROZFYUhsqpf3ktIi6qFoJd68sNPHT8XTAK0Ma/xocqOBV+y9xK
92HYw8aFnZ338UzAxss33K2/Fx8byRVxIZyBaThDNNvQzaMwC3wz7LrqzHpZpnQC
naVpMbuNimap5wEei9VMOpg+XHrRh4An4kmF6ClLqK+7yeI+Mmq7OQ99ZD9DofAY
GpnQiypnw/uCvxVthmRdiqfLd235sxUAfs4LWx98R0eeeu+Cy9rRsqtTTSbtv8Wk
eAzHUUcnDmVZmJVFq/NZ95t4UX33kDr02CN5WmMrF22Ixll97NS5QV7L38ElZkK+
7LTUXjRig8KxeAoPpbMOkUThcOJ9qu4V/+Y2Lmrm42CXDm4bxnWaONz8pb0IO1OL
FYax6sijzFP95zVPalRUCN4GcaCg2AGqbk4qbfsUe8tbpJ1qFlw+6qEJ5vw4F4r2
1zwXJr2Lz0B1qjq8m8bi98oqMQD7VvFpxjZZexchRLEUSFTwXNhMsPlbL9Fftil1
rAaBCXdf5taCLDngsKX85L+O2velUSJJCFfDUqL4bbQH0+s/YlX5V5ecaCmm6O0c
mJDow0G998QVkQYDt4XroIHV+erdWDEGQ7ZTEoigz2gfVpa5QBSuYJ0O1LpKYB/Y
8heW0Z7BdFG5Sd4Fs51QojiNenQzBzf38cy9OEIZtfLJmxjtLlc9W83x/WTwoMpB
wbvr4Rr1l2GP0YYv4cfqa+Bzr6fHgwnXhWygwdjOvbvZx7IiKNGllv08K+7M48ue
RGpxZlp90cTqNTqul6B8yFo85NlW0dQn/RVgmLqTzvsEj/BS4TYLGOGKLIIH99tv
X6zewEcZPtUafw+fZOLsJH04aDY2+qBPcB39IoLynq6spBDkivrwEJl691atzE73
PCaFtiqXEgCPh4dAOjTJTwyzHFxFgxqATXRcPUGk4dtbsJBEr4SY65jYtWxpN1hP
yAv1J5Rd+ZY7PLj/VuMNfIXy0qO4XkPGEkrl1O/yWl0/zsFOFoOhaYm3SL84f9ap
jF1uiIZp6BZQ83/pTl0xvmobRc5zTgjlxzGqu8mgY/oSLk9OA/l8rZi5wh4ZHXhd
E/HA/BHOpwAZYi5ZgMy5ATDv3dj/X0Q0TkQu8AfGnZYHB8jegnKOeO/gtre291NE
/gIj4q6w4WirIpwNSrYlIetsEdYMYRy5f7MiPz3GR9NkaOL4RmX89VczNKkcxfdm
fBK5E1ZGq8d2ArP0zJSkBSywxYvTVI7wSj87TMiQY4xQVE1EswkY1JFOzbnBKw+c
SZpQbe0JDaGuUvl0bSo4Lz03h22LRmLR7kQsbDiMhDO5NLh3zkeaq2FH3wr9aNVP
904Wu//UE5llAuObjgLGiYdqE8UEmFLnGmLO6uoLZpNzWwyJGwSIFN0PZinaFTIe
uU+BQPcO85YTzb4Xbw+dwPIYX38o+fvQGXTY/T8ui3LNlLv16ALPbXUMkTUabMHk
iCpFuvyZtygzwrhWNV3diJoww6rtz9LJ/gvE5ypQGgRdoq28a6TG/MDxPB6Xmlwm
yvJuo3WnE8JpUIdlzLokS5grI4R1YImGgwXzP5ov+Gdw5RwEBwFkdL5nxqOQXdfd
BH1+uFzfiFZPmMhGBYnVy3jJvWCS7MHE6QBmqRmsQXpmg9sMwaI9XxS2QDB0RYKs
VHG8Uikaz89qILQhRYrSy4Okzp4rLJqf55w5h/1eF+IXmH7PmdMvo15tuZJu6i4o
tS/2/jUZVSVAee2r/d11qlhK193liOa+2SGzG9thNZyUEYJWVUXKvRyjdoFBSfoO
Fj2ZPrsy8yx1yqNN9rcp4bmkf9vYgUdGGSGjvqasjxAEBPX9KqIqHg3mvvv7u9qG
Us2yXVkxaEyfLtz4vkzPILP8RmauMYrGEpwMF4oNHn+hfb6FvGTWpAsHsa2Tl/zV
HC0oraL3FEzNo1BRKWtnYBtJLzdUUNASANZYvcC2dBguL2mqOYNqQMfaRL8zQHsN
2dqHcJSCYd34hRU/XPs92ASRZnggroRY1LFEPALhZvCd5w5+3UYDbj10EkULZa1H
RLCizJI5353HUT6hnW+a11AxfeNd5wH8li8hH9X5yIudwMMwY1yWEGPmS4rKT+/R
IoDidYqd/88kCvDS5NfCMKl570vjKXf8e28qlfxlGeELzhT4NqxXkRf4cfh8LXNM
5Xe5Dw/vdgDpCHa7Qntj6t6yb/L0ersc//u8fU4VFMohKZnoB2dmzRBfSWUm7msL
OlerX9jXMQMvgA5RS/52Ecm06XfC34RwNHWAWajcD64B1Z3DPFiK9MAJDENcijO3
KCkpSLvU2jykafuLW3R3ivtuqdbeMBDeKHZHY3h/ntqbqBwI6d5bBOwzEwXZVcZN
e1S8vxyD7iXUgylwggHolmltMhBRsw4+GHG6uDDFDO/AfB9n0QighXTQs2XBWyRz
uDuJ431XLJ1nlOU6KRD4C+fZk4wIj1mDRvkndRMny2GivvzFJQ66pTzuHcBqsrHA
Js9LYZqa5KjxaEtlRL6UYdZ09d3DoNflpNZVmaVKBLDSuepcZb4J6FzdrkLA1Ypf
52fXyXsW1OiNqUhQ0xbXZryIUJfJ+90q4SP21qI17AQVx56JKHbxM4E/70NbTz9r
+5ccfO7hbavIu8SoQAT5Rpcsgx/geFpG9ugRNDyBwUbssOCPaaRcULpJk0ft6cJz
k4kLACiLcZ3NpyRNSXM2rHEWMfZZ5OrW8oTcULJNArilI25MAHgdmFvoUpFfviEE
GxRv5WhWfzNAEeU/VDtLPKLN7MBqEKDSF+SmICchjKuzRukCGw6ffqePDQeJdOcU
UoS45/BIu8qCqAQtT6HAJ7sSV6erJL4iDhMwbY8i0dOJ+VTOZ9quHHO85jRW8fi8
z6uDJ+qBXS7q/8ZywdeoeTJVuUt6w+oldnEP8aIx3H9pFtq2xB/zyoE5KyQT+KPY
Rixr3eWof5zxTNCZO022/bCOTT2fvA2t8UVtq+XAP+UU+OfaTKEVcvGlzmDfs+hM
9Vk2JetNogcVte30zmXfWF3+RfsUzw1W5Bx5sKiHFKBG0AyY2gxtbhlrgGVrNI/n
WQYpDmqrVFHZyY5IFhFxdPJnKHNRMLk8FLw6vWkoyFa6MhnGOIkTgbBx69szrL7d
jZVYea7VNiFSSJNcyh0Q9RJtLMFh5OmF6H4N5fmlUniMnZCdiic4IFKtfTqCvdkm
14Zm8zwbQc5FVsZUUBlPOyOEVuW5HLxB7HKvbwqv6g2xBn3NQTjdbbXXXveJ6lPL
M5PA/kPY4dArRJv+wIhyc8sIoiUxlXG7YfzasrkYbqLrgLSVOdov1Y2ZzlvousIs
E7GPLSrs19COVygnDRQLc/hMa0EXnuOW5pRLux+i7t8hwRlmmABTSHBRFcnz+6t8
It4AnOCfgq3R5hJzlmfBrtwYq5psuHSt6qNqUENrZrWDcP8dKC61Y37O8ryL3YzB
QqcvZ8EdEVKDZd7WyhPWtXLq8bn5MldYdk5aOf3CpX7smFsSDhROHmUD4UOgl1GF
nNpqp4Hb0Yyv5Jp+mB2B+AcP1qgEHmOvZ1Ki3uytu3xxpwU22imWqhdZPdN3sNUW
XAbXxMtCitD9ekdKCVPmGz2E3XoNlFWCdeYlFk8qTvpBWPCvAXdhvXpBBi5G3c+q
uCQ37Zt6b1pDGFG2Ej2Y1JUQkG22cN31lr3gr+Mr/csnRjXaH27PStej/nZFnI9c
chdmYOzNp+1je9mjaq/WjyczSme4IuOwuZw8tB45+BeM+Z8S0bwx1L4eqeAkquK4
ctOdUBSFSkyZeMCaGVHa32WvOrDHknhBtUOGKzIm+sw5/+9tzQvC4T7M1JhlILP5
HZS/y9Jn6rwrRZhHbkbOWNi2QLM09bkcJBbzPOZ8Y8GSZLUS422qcziDFJOXaLMz
9UdNgi88XJ3v6liMRM3lt76qdWFsKrmU1D1S5flMBHqDAR6Tqx3a9EZgDBALLDkJ
C9UV0xHz279rGTRqeCoPqr4w9ELdH+mqoyteie03/h2f2u8KJTYC9//r68hJN0wS
l+oi26/RuqsABsS5WBocM884n1VMfGx57t9E0jh/cWELlE8qR/gPMSke6dCRpSH4
Nk4+zCfg1xS9P48Wtt9BjP131VSC9Epo3pmmuXw+oxLSR8f8BA6gP+xNmZfAdV6O
wMBor1fclfEIvh532aBu4Q7OXQm7ImNg2ZwvnAm4KZDZo1dcELjrwG5TsmHvOPlS
qvjEea+wp6QK/DEe7WJwQXofUic7aR19Jt3uDqtmf/9oxFC8YX/6gPbemREpWz5E
8neSotJf0JtZQq218hqLD5R6g0D4SeQOZI2Q6EDDAI+kh6EIzBAzAV53bowIbVlz
1Ty5hUdEU3VimLXn2hHjKtMq0K+aoqTPDXfWrEYl4UE3KVLYGOqSjM+DlvCJnrDk
Jjy3uhPunGDevohxBvegz0d626msjE9m+mqvkTZxEVsTvTDAqLbgscAXSQSRF4Qs
4stWyPsLskCaIVaD1yKRw3xwftpAOxl/XbzIM/Y7oP8F3SrY8/HcMDRxzPOuFhsr
tIoId75JYxI2Tnyw0AnvB90NofbiPUR51rafI2qBMd6tXHvjGsHsFqdTipiKXSR2
NA5iLb9I5BHYLYX/g+C2UyRSu0XtOFVUe0K/xPnZvmmAFu0pW20DjuhQISccl2m1
YTQIiZKU/ztfsRfEpYMvoWNxBn56F1/eB6qQJAUqIUArTdsoT9cLd/dMluBDp1fP
imE4VZbUQ5c1fyx0vebC1+cBedIyoWdAkJYa7hgYHzF9mmKzJ/Y0BiMFd+qlMuoC
hw+evv4s4HteZHoAYfL/NtvqQyN7CeeOTIDoFRAoEOvu+gEnPaPQ8bynm5JDA7bN
kTqKEXOg1e/j8/0sKzU8RTTnlIkLmnVhU88RN4knkSAa9vKcwROCJtcvu0qJ6+sf
mYGFUEYZomIQJosK+S/Mqk+8DL2hpPwvCbm7oPofeVIjlMTqaCH552atR0L7IAgo
9896/8xwdtTVQ52T5eOkge4puL4h8fkLEqFWcQNOd5+xEt3dppIaA/G07VdQRWZN
TF+5RTGgpjybpEYFI0z20/0ls9KnFkhInZ3liBeHgNPot47fL/no6P01onY8DqGC
hOwPGiSzx6WtrUIkpaOoef7umswlCE2BqqkkakfWGRFcXp3US6uZKph4cOykcLXi
Y9fPFbq2Ao2Sf/EKB7V8mm+5zlbPch5yA+ZQeA73IrIEN2FyNTPa67Em3Nyg5rkR
q4TJzkBv39sjmDfhsng9CDANbfYqwg+wADLv8gMNFK1oNNuZ4Yh+sZriJ3/J77c3
pyVDm08gk/0dlZlq/nhsRJ85RUuPi5LQn5ZFD5hYWnW3yIQdxobt3XFbWUlrzngv
VRc0kLHKXznbXN4sgAnQC23VRXM4qUc0Gkjm+8fK6i+L66KNm7qYabMhPf2peIOa
/BRkPGMMHfi2QvvugwKrVTo22eNjOkeXorkA6IwqjEz1MXjvNnGbX0ZmosMZ5XYh
hihKjXI6+vTDPddfZQm3b+Yao1J/2rVb3GEoThuKmZG4d+JIEOsweOpVvKdGF2/d
CY8b9rV+E+NJZi/mcPdQ2BDZvyrhG7km4OPhEPnefX8AR3JgnqletMNExJDT2Atp
naiT1b2pPBegfbA7ITE2rYzKe86Pw0RORerC1dVsJaAU/nMvEPnuOXsqBKNlY3Er
zatEbL/D29o8/Cwl3Hi/b9taxG5qmXBHEJ1iAux4NqU2sLad9wl6YFXl8ZZCAENO
/HHjc0xEBefMszb6kcxiFnOs3kOikyGNcfaFkIuN36OpZfI8CUzTrzlKji7QKhlM
WtVTNLz+zPNcLt47Mlcxs7oxkHkUIqUVZYrjFTWb9GrWrm2P7mvVMdmDdQsOkb9T
2x91jN1aVsD1B/XuEje6lA19L5OAoh5w/E6hE7YyVNeFhh4fLuvzKsGW1UI8qv2P
trL/J/VAsallxY1bMAwSATtgOj/Hb2GHatEAMDmS/FjaeoCJhhMsbQbeDS3bXqo8
iUQ88Q0O09Q4OP5zOYmIoNoD/+X0aLtgtQIBPKfBiEDcFnacDSOWxLsTRoN1kxIk
x0v33z22hhVFGz9i+dp8JJeje4RJwedMj4MSuYMyH0nf42chl3hcZAT51VfiEOl+
jBA8Vvk4PkDfUoWloDj9AEJ9SA51EsdjIrTlzGpTGloHVBfqfChDJW/t6cQF0LMc
fChGsEGMOJvypCheXTY1guA6R3JJvny0E50FyzPxUBmY9YJ/hBYNwIUYIYYzJZWe
tF0JFl4vRsDLNZ7K+6wsH50BjKYeLdsNj07sUX1BZcaZhNaVoB/+b0H+8UUXv6U/
sD7O8EdjigCgPTC1SdhUwncfHtYqNUMW2t3uX54dYuBSfl4Z2+ezhuffx3gqi9/l
2CkIGcam+ztHF+8UtRiXVl127LcIY7PultaCWzEni5FO+p8ZnoExAglNr21qis3m
p3s6QA5uVkVxl2GC9lp/pvOvQlc778DrcODBpJOdiBHOTHekvmuZv8E4JtlGjpb3
BvBW89cwJBkHWhQ7hVOlYD7Hoxb93MsQNcDcnPKwkbM0/vZlpcH46DOGNs1R1gf9
VcTSH6o4tRiHSc2W0Jr5WpwUqcB7OiWUIc5PI051xbt8H/oqZuvJXjr/YNPgkq6J
GqKkQ/iGnYaoD/5T6uopcJWWskvIV9RFTOZgl7Ko5+PQqorODaKLwrOKjSfrHd1j
uZDorDws0UWqE1Vw/Iio2cHqGfPA3msv2AVNi9LMUo7jQ5jfKa49e+XyyMNJfmKK
IyzZ0vX7Nf0AIqTXQHJXSonJc59ezQ8OMhVjU0m+cuxlrI8cTItNGkxSklqEOkm5
TRnsvQMasbOfJT+xIiex0bS+jkPXx7x87qMdS7IVr7jwSm02xn9V9pp5dz8ZFeDe
BkTTzz5++TX44hPAofqGkA4C76P8CBH2XIu8hqzGLgAIimBNa2a353bo/7nUWkwW
zGo+UIaKiMgWKa7acEKnDgh3QZ06SR7Xc2+WdFNf+07VsEi9t79N2k5YO6Xvp1zG
/AXaTSlf4L+HWxMC2h89+E7DyNpVA+bsnopv1D6OLganNu7tEJ0E4OWSoPm3aZ9t
c4M1usrE96jTy7T7GcF3JIcVbV5BaTK1r6z/ALkzNxvp8DKlY27C6ratsq7lRhVM
IhQSGcg7LWPH1RqujuYsnO0SHyp8153sp9H5sOy6OkSbe8P6wB1oZo3yA7xN0Sxj
2uG3BkOlbqn+YrwHjK22IYLwQAqnk5zTQae+gE4w2MZrjaN0pY5yZY7B6ovx0jdn
LKIdbKRB6YSOwFWlCa3kuUS4wVeOKUL8l7sxNV3IzhEHMHSWn8NMaZ9CTAY9MHZC
c0rKnMjblwTsI5MIMCjjYjm9U1P77fU28+uhMp+h0R+jMHYVrImr1Bsr/MmCdFi3
/BjoN4WfskPRU9AZ2yevbIMrzgPO84CJurQSnrJFEPc7a2vzIrybtv2qxc1Et7mB
37biDCWH74LMlHJin9HPhEkhRd0LLY/l3ScKflNc9Yn9YI53XimAxmDjTU5xmT3O
sXN0Uk7nD+dRvXt5l5LrtUl95Z67poJ9pf1zq/oJ8tBKNwShn6n98TXeMY/Y8O6m
1UthbYa8wK4JckaOQ1sjJj2ZKpmx2Ff44Q+9dQRzAd3NFQ7aYo9dJnMPZHFEw26i
36AzyDrEyBg/eU0I/HEZCeFEdZG0RSRyZIFlOkgA4byZBM1DUAZxnrlGu6hUI5KT
GbJLd4VJtuo/j32RKfQ9e8YfyzPP5/TZkrHAUjRMGC50AxnXCqXcLkLqNRmzGJU4
B6WN77TrfE7O96zC9mBS3D2Fu79YNo7IaRZlpu582aeCOm15QlMLMzarqmJm7y7P
1sxagS7fRpbW/xXa8NQNzalf4c8cs04HFBCdw0sc71ShaV4lLJQO6H+Iz0qZscKj
nFno3qAN0GxzqTIOLfNoOV+Ru8M1BBAp1jDFjm0TQBB+emURJMKLYtquxixbXJ9B
0/1op/ZE367SZEwz9272+QmjQCmsTJFINCuQaSN2Wnx8NVtOloVtNiYfQqtTN/iz
NDvqHnuc4woFmjikF6ZGgFMK3uZI1v/Pjow2QSoDOT2O0MEjLozRRDWrwl+XQfyT
dey4WejfeiKoPeZVhNhRFlWZanYJKtfYK9hSmmm84VmZguDNLXfeIp+6MmdmWDko
MK4TmZJM4uDiiFypnW1Vu7l8ckU+y4Ox3EmueklgX4AgLrrQxi8cq9HNyiVFfxyw
vu6AGXYZa+v5A75JxTUy4++QyTOdJlzOkIf7/tUEtsfL1vce8A2AiJ2h0rK0xd6g
DC6cT9HLDFvpNTqpmX12TAWBzr+lfTsv4OXCgeF/IeEGa+3Jiz6okE9XEkeoCfxM
tAzuqLfvcMzjYZJ0bhT2BZQMqgnEIrLk/9DNcLH6GSxmUcwCU5c2FDMBeUPIUsFz
UvS/9vyZDcNnurSJZvafBYbmtlML/pTHM25Xib5bJbZq1Y+iLJfBdSmwbGOy3n9S
LQZLkEzZAdk/3KZMfO5aAf+5/HF8k/3Cef9et2XFpgOl2HZGLRhrjv4RZfGrNtZd
tsKVb9uj1mR4udoWorzeEnK/4oLIlL7PbJnkbqjY4Sg24UIXHKfvolbroRt01Pk1
1BYeTqpHfjur7w8qP2ijMHGJTWAn+Uny8VM+TN3GxLPLAccnbUQRjv180hxEfjCi
FE9y/tVJBg7CJqCUMt+/cNbPzmK0enaAILhTTBXACrpv6aNIDLJSQUWUQpB5lFa8
ecmfW4NH0HwFWmmkjbD3kZbY9d3mc3ftgMBlL6rL9x7mT419DzyMIxfNMfLJVWY3
pi3J6gKLltxdmUTQuDanCcSWVmeNLzQ6fZJw0tgW01cU/ziY2owblYCCEpATmlS4
BvyV1XbqoTPbClyzvCzctBR24Bh8Rg2sY5zgeof9oDaBTDSMFInl2TJ7hZLpfUgp
1bG4VIUucS4Mtlb5MvVHhkrFwP1+0/c/L6J4n9WcBCZF8/A3tgHKh+TkqbKHLCHW
iZ+Z/vdYrFMQQ974i6uwTpIBVoeqlm/lZoTjUCt/pVJhzJyJbiG+qTxt71YVw5i/
xYTZwIXonp5D9LUmKiM1LbO4olz7brfQU72lNz2fS5EjAke6vGGp6cY398FBhgJW
kVGm7+g73kRYRfKZSoo6WFz1mp80TcJqvpuM4jLcrFBkJefrxt5KtsKHLTr4cg9J
qvkWVZYoX7aThr1+EVMGqQZXl2EIt6tP97V0cWqfviH244VRsH8YoCLuKxc0sUwH
tuvfhNY4WbNa+vg/iFsb1YlhkItyuZNaQuAkzS8wyA0rAcMXkDbWuHAFD7ggENdh
oWIZd/kh0Ki2Mh47nSQoSRAcUPzZH++yMfsk7q0z+xoUY5+Ix74rGe9eFpGcg0+z
e2ti7Xjddf2X2pi1QBz6tejSjsxJRPU1EUFSkjPLue5yHrFiD12jr6cou3RIoRan
AphwbrfHVWRq5ppcMZiHmvioHPuMJ5Eblggjw7cg6r0wv7xSU9Km86fmnXjDldeB
hXLmLOYuNnqBYmK3A/g+U9LPjBQ4Hq72gCfsryy4pWYT0WPze70mS1Z0nhRHWjdI
MrwHH0/ChUTE2R2yS+i0a1/awYt6aKK0Y/G6EI10dM1Drh0mpHS7t/KSvHhvHHRU
MdpkcSsegp7N6NIKBJJMTucn/OkQfT6YSB4lVn6JgQ6fC/3O/IZtDSiQh5iujnYs
7PS9Qrdlf+cJCQaJAK7mBwZcR0fvulC9nwE9C3x+GxNJXexuNdRN4pdN4VgPSfaG
bkeDDvpwTMssRlJ8gTR3TtXYZYFcdwC6Ru5V5qdlyOrDdsHWt0JyHofBhuyoibYR
YPJw+uN9F/NHJ3flGfN0/jd1kJIOPPH+8F4rygWNIIUWaxUOuZomxBNNiyjV8zkM
F/XSmxByDos6715kuQPnw6FlshiIyHMGQXfCzC8+Fxj6zV2TRx1iRCoW9krItUbm
lT2asgC9W/HjK4G1ALZuIq/5K+AcivTSRY2njJ7eVrm2JcVxHMJau8pIxnJu7Epf
zV2dYfjqzPfQGx4XMM7NmysOhgOBZaGwiqL/ZMTAK3HhVA+FOA9rS/byk0XwjIOg
ga3nf5fAllpUPJGIrJNY3i3EWCtzAvjiZZ5rCLw/vEO/g8YOHMJwvyuHYp2ddtH+
ZbO2FucPtx4OwxWWK2jgxz9UnoMd7Dr4QKNMAHhfxW2kfMbc8OuEmc7vI+zadZ1n
31X1OusnR3H9FeRW/jsy82aFAiSDMOJBV6Tfu+OAxRlo+xVMR8DTpym/98BDD5Vn
NsSjPP41XSvO3ajULUFea4oSbDiAXZ16PLUPzSFO/0oThlrSQIaigetXcWgYalVe
E6jaYa+atYVZqKFI2wxEO3sUClQVtvLc8VJUUsVRxqeHN5MOFije8ol3+b/48Sm/
uXC4SG5Bx8B71ARXaJE0TbARNupOuJSQ2e2+uSCDAj296pOj1bByHuPwUfQNAYgn
I/HQ/X5FlMNPVoBB4kr+nIEX+ecFTTJOOZc6LTl63oUZ/8VIXeFM/iat0RgPs97S
ayojC1oh6HONPUVlSex6wq1HoEzYsfjGvYIO1r286f2Ni1mJYc7vlc9PqQbXKLUP
Et2RgMbXNnH0xHR1ySJOO1H6G1496GwZutXby0LoTuuSeZk9iaLzfT9z2hIehcNn
C3xoOU2pwq3CsOfNLbj8kC9GO27VSQC/hutS3L2YzC6dErRzqXmHsApMudtleGD+
6arOWy3Fd0JfgwnEuM6SORfa0iWM65WDZoo0kmQoXec1RgiEiFohVbshqNDcv0HC
EZ+0f10QNhp/3pQGDRKhiKpEKoqkw47p7JuJ/8nWiqNZHLuhyzgEtrRegNetPfad
46pMD2vtGDjmez/YlvJYXbZWSzDfR6PUos1CnW0jxsUh/keRZ+4i8a6ycplJf8IC
Wuw6JWxvYzTIIi7zox1h8oSiP/MOpTW4/O2PznXxeia6UD/aImNoxzMhQA6+ugra
SHx+ehYqQuJyxoL/LYGxt1pM48y7ViR4uB3RDlFqkjrlg/4/+ymECUZaajAGy4P3
32T9ezHGFNnkhCmtPBCHy/9wkhSTPnQkp8w16v4e1AU7QKDrRtFfY/LoHzg2lRwq
xIDUARFOmgkuBZAH/mqRhwdfFFUrwdXF3wFbebl9DxalfDyug3f/w+KsamCNIQZ0
ZY1/PuMqvhLHwkMCNU2cPrpV1ZgT0A+eR3ApvGnuAW8HPCshFIMT5JDfbQEjxkgf
V6/AIlIeWs2AIhnLuKE137Z6QpZsQ9C7gLjckZKzCiHb9+f6rVwaVF0f3vR8u9oj
mvdZXAa6hdsxpbd/7Ns7xejKqNzLo8cvqGGy316KRKY6t5969W9QvR/Jjm+rvC9c
f4HM8otiMA6OT1oG4LkRgXt+ERxm7VYAiwnENLwQaHixZfc7LENwAcNf5a9z5Vvu
3Xili7kCOwyPXU4qFHwRR0YYMFWLQUmjoKKZupL7EukNX73mTjKuvX5FPppn2jfr
Ty6igjDcvjyA4ZjoGpUpJNZCkRb5kZXQgUna9y6kQNT9fBU8PP0cyPSXrwKQ5Bmu
E8MtIRpDopr0dYR9YBpeyfDpDfsK5M1gcJzPjJVLIZ1FDCDa/sZahyvprOKnF6D6
3KFoKfKFh846oJTkB0/VI2bwNYwR/jJ8JhqmhrAt0iFz6E5/cqziOabz3bpYYSPS
jM/7nZC7b4WDPvGnsDGlqDJML1as9a9cAJdX4b/U2SR0e/EPvBTwaGcPyrYQKOgH
luW+Mx1w/0SeXnsvKaw8DB5woTHhw8AuqwMGAsVOa/rxkE8RRnEd17io1USqvGfO
p0teBRST+Yq8p42PjDRqAMJ2gyOQNOirH7+KALeD1t/2j4vQ/S7kakRZXLrq1UCq
UOmUdpUnxoA0AHzrLEBDFj28ecGI6gE1FnZOp3FhDIpIYLKBQ4xqbVAsZRQ12BR9
3Dm2+dimuVobqPJMsUDDI9itezQbi1bUUeVyj+zqViubWryw3MVGosOkqNwLyTt3
PcnXE/0i1sUiltaDbeFvM7QHexKrm4yqcX0vqj55CFNW1+lZlOfJrsRR7AtGWhFG
DAwVIjruRQi/daLTGyCHhwbVg/RZYrSL5X86lpSz52aSi8nQPb1GeBRVkbPoM57D
mzt7wdvJw32Fak3hx3bDFjqmcnHPI/X7VFdGznMymCMwLivGHc5Y8akviJQKqZCW
egiXTmBnDR9WaEWutC/Liqo5KZrf05U+zI7xXfULnP4oBr8dJdw15zbveRif3mMc
B98F1qTB3T1pW2egndlGRpwdP2xiOd1SAH/d+PmVaVMyjIRpPn+8Husa39Sh4cOl
HVbabAkHzBmz/c/JO6MfYIUcCRse5cHWu4TO1DMAk9jZYlzsxreF4PcL/DDGW5z5
Jcyv/eLVqWuFJOz9qoBlu8fFNRKpq/5TZ5Y7u3rVFUJ+FYlC0wtH+AZQg8L9QF3Y
Ulzi4vppCOwPbpbfFv8wu6tgDw7+kfBN2H3WasJwTXDZ90gC+kYR/+EMIhZb1LM2
S65f/1Dkzh33fouCpJYci6y2QwIRy5Mo/ThysnnZRrhCoul2XMk6WAiH7yfg+P2N
z0We5ZqleNuoYQhElxV1q3i+V5H6gxRbUju3LP8LeoSIq60bJ0W/7An+d2Wg3lWJ
6tsM1xy3P8THzp/oKJU43jnDdxw/xb5nhk+JZAVtTltqbJO2UVHU/+QUcbiJDobd
G8k3fCmyEFtDBKUt8JBB2WavFh7TVrkkRfvrdVxAWJLZXBEA9XQ3NXMgQ5TaWhy+
y8N/5ZPhuFMQCCGup8FLLvny8KrxR3rXwMKpHigagE+Ak433FA70bVcNnY7VAvv3
2qpX65ZxzlfikKZgypaJiaan3yXW6UjTl2hUw/xlc5hxrqfUpKrFyQNAXXELxe0z
+SD3RHnoFMbq1BEFqD92g3cIBtPGemZL6rzsqK2TP2YHKYw3PQOCCLjDTuP9iLck
5lMxnYXc5bcanM257Qc+T6FfS/M39KQs/mbzPAbRBwJdpzSdmWQ7C+Lbh0I8hEZm
s4BWpEP9SwSNJ0m3njFeVDWQCQ1Al/FAsS4alzOXHm9+DASoc9np7wCdEP0SEqzP
VwOkXfFN4DDgCW2NkLOkc6tGemYwKXDVxA/GJDLeY69Umg+05L4IJpuo/K+WLkHo
RnYCexPnd3R6ce6ZHESWtZxwNZgJ+nNNKzHajLysI25vk4tHIeQ8OFaLmmqArTlJ
jSECONzmwzEPYHMU0oQtxkxf+aC8s9Z7Ub8CRp3t61MpBjDypmTWHyOEEOXicUxl
TlQBoEarzZuRmpw+CdUQf0Yn/myjapGec2+fnUvKIFY8H5PeejD4GT36KBf7jZlf
Ws9OFagJW6obo+iPn8zL/acWUD7EdOLuBnpFprgVgUFf4FPqK9WxORmqTc0+RNyY
qRu8+iUtFsDT45LjDGkP1X+9t27pn36GRS83jcxZpF2nSojH7ZSp0o97wPfeACrI
u6w/SKV3sY5xoOpJKbokKMoLHL8WIJJs4oYiUiFjFFyTZXlS2f4PNXZJ/LlIkdHT
jfepn+bjv6SFvOM+4OaST5XEA9EfknEL7SmK+Rro+rJ9SbCwduyyjtgiBbUyrU69
wnkd14FWsUWPtqFhlAyNWWMDeDTOuD11TTfjzVnZkP8NalzJFzkytPgusEyH19mU
cKrz3kZaTqCXOxrUQUDhiKN37biewi5fKwzpOSJvlIHIu18v8gGrix/K0APR3Gom
x7vgm3Nl51YTRSoS3moJ2NQ8oaaID1AjKfamho7CtKQb17/DvPqgst3L8txxy2Gd
7DSn0ZRmAHgWQvMdbjw0eLBDoHAUKgYQBsdXehhLwkGU9DaE/XgsBnRSpvJ7CAtJ
MJ/G+WLf2i6LDO/rrd+1kIgmo04UUAnqaiQ7OeQoWB2/ocj9HhnH5wBRbJYhZuQD
563kpeaXLGVm0LGY4weLnLXi6e9RxKimLnkCJcJnlHiQHvESAFqF/jEyhMdjFoPR
r3DYgNemhudEOD5sCn1/0TJFqrIuWsgOBYnIoGFpc4P6JzhEci0zMONAzHxMeFEU
QIZBaW8Jf3oeUIMus2B40x8XarwKpUxXtgn/Jx9kdkiB7uWBSPEwtcxz/Clh0AFb
AYtcIKx703WnDxLWsBaBavgLP+YBIrQsSfKzGiEBMQ2ox1MqTNLiWdPjAg0V6Q4g
fwXc+g9al6ACRg4uXZ7TopFAdBMAuJU7JusauWzHLmFjIBZjxzw8CCmO46xUSngo
cNDFuWWaW2VTUd76acRFU68gYWfmJH7ePr5Y3I0MI6/X8CUc9FXjZuV6sHwKyvae
MAaeBWIBiyZ7beN6T6FBytdjU0v+gwf/V/rv1YcHRsk5rV8oDZEhNBn/x+D8jsY0
EwOlqiqxXWd3nsW97FqhtFU4r+WfkCTMAYdRpyXhHpqYnN8rd4ibaCpUEU1ZHKuf
CBqsNxokiItQxPMujW9GX2IBZGdfL1h3/wkrbMqC0cM+wrnhrAltm2OjTTMDYTLO
XYR4Jr7ctiJwYWrwMJoPMI4LX0jPn5ReJBjgWjy91n5t64fAMERC4HVFVAxjM+W5
DljV9hHeI9iPchiwho3Zh59Dfzv2alrG1InUZEjeS5748BiqiRdMSt4oWn9zNLzL
kaLaGsyuOH0SVh0yF2LHvisiKtfO7NJ60zFEJ4fZyxxRRraxRU2fB50/cZgmkGFd
id5sJNnBhC3z8pdfQ2ALsVqTiX3BEAJgvsOmrcwbNSBoSy0X019W1mVxWrOGQMhY
6PWjCPJaQPbmmlzXL9aqvpDRBF+QDYdYEkT1diB9+wUT6kY+gLrbYfUwRnj+F9QZ
TMQqLQ++dqXy3Ph+cgvtNMHQ8Hyz2InUpCxBWFs8vPdG7OJYKwL04+GQF2SAvSTA
S90PkaBu0RLWppB29Z9YHZ79x9G/k5JuarsYDWMQlsmEHMH71V/djuk/+luxEcmW
KIi2BqdfXf6bEnOgquG2G7JLccCrdpqFjvaiVyI5gwcE0bH+d9dl/L5X+b7JMYCZ
gOI4H/fsV7JdfmZIwsumf1tuSNGH0FM13KeWLthSJP2tRNQkjkYrj8ghhc4HXJTF
SuKzKc5a0seJyaZ4JyDeslYZhhnmxmMuoPKfNFLIjJnXxIwe53T2mspwnuWSoxsB
VhKt5qn6h1dkjUw9ZviVCEnDrY/72dXPQKKUrb2aCWTI8zYFvMsXKpNyhQXDKdqq
LF9Upb850x2S2HpPDI7H8WECaGSXoiME00AP4jd4n3N9fljW1gKk6KUfOozpL5Ew
SgXKyTQQiFisYjecflJR1WOQk/OUFX2pdc7DbBufxx8LhsIpTYKpT7qp4WajrQNb
SLOQfBVXoNnT+TxFcWniRhMKXSD5vtz5SSsq6I0RmRuhWthLWRye+SYsWRCxEhDC
9iDzAZJZAbBfRKQ3AwBqovl53UsNw0dvJAbUdDLCV7g1DiIdOq38+NaCOZ65ra96
2p44F0+aDa7g3TMEUyZPnP2Uxi7WKZxZOdRCXTAL2W7lMnmkGvluKcx9gfoKfg5p
QWMdOfvI1Ah8kf+P582EQjOs/cPDvgWotB867TLoJbYSs53XIEF2QFMc5dOGHoag
YCXNJLVMcWhBhWXjm9X6KD0bULYqJbybM5pnWUOt8P4Mpcpko94ldE/JufKx/ngL
A93gEI0sirQfPrY+bA6Vl3Gx+loYpeqSHk80RTynYMu9Ja5SjmpW/qI6PSEIxhVj
F49dJXEB1aeJVhKt0S9LFdKUWEFldJt9B8CcYZKpb2FlMWYBWuPmtPRZyT3PqAja
7S2m+hQXQ3F44a82vQ2xGSr0VZ4v42O9lGGU9H+sk5VQoSNakR9sFs4Fq2lOhvVP
DPB/iGNTvC7ES1DGPOiqjSDaM44y0J6xUFvv8jgHaTFn6ip2wDzkgRMBfzLO6JW5
kQoHSTGqU9cLFNRiAPKx0YGZC1dA228i5sWzT827mle39SL2KROolXgGJeQ/4qDP
jY1STddrRFu0/teJPXjrNH2kAVrgSOqxlPcKZ8a9rh5PiacUEqFwTZeBqIB0JZsI
Nu6LuiEb3NwXL6EKr52lZfQhxz/Ep2Sn6tAKd70MaRY+IC8Q1m3U2Oropz/0F4HH
SuJOYw0WsgFxGv9t6DIwVfNhYW+i8EEcXygJVtkeIRnO6+WBe1VdVTzj1Bhux0na
6tR9CHhd6fS4RPclscL/2gCkInm7+xUCoQ/Sla90AE9IIUTDXKLrKrZJ4E1IVjLQ
QwLRS1kf3FObiI1t/J5uJOt2AU2k7++V8eZWwZPk8/XrKBBhr1HZEXtunMLq+Zcd
6zUIVyPGBMc/+O0Ziuqe+b9qX144plTAxEZPYmJGwaOGm8FdQEHNrdgrtFnm/OOK
8s6y08t/sYjNWyt+ZJ8YbDGj4gfokf9RAd+m+boZfJrNHvgc1RDT6dhHviNfw+f0
cPxYarcwBggLb69+dBPY0cu9KyCG8X8i9uJr2AtoOyk7KwKnhX020KzUeN6armeN
qKuO9F9gqUW/+ifGQ58Lt1vakYKZvli/5pYm5hSxStXpA/2sz2C6CpZ6Zg8jRe+r
ZUkwyTbqoevCtCFvUb89lR5nZh2ixweh60GpHmWWTnky+Uf+5PXReLLCJ1JjsP2D
+1Szu7r1LnYGzOdsTtgjZfgtADyg3OdFL+7XfxWxa+aBghWMTzqhLu4aQ+J3/Kqo
zMFhx+FLcRrJtygq9VCjzEagpsHeEdXiQ+iRdPQVidKDNzlxYJc2zJG48HS0APlw
LxpPftIxcAhXFxSTaYRLU9HjV0jIK3ZdjFKKUWffPGQkSZEgfti0+A5RndSI+vt9
bkxIdIAS/hlods+JjIa2zpvkfWTr7YzogHrbzQrKLJrYCbv6IczuwFXHjbOKOzOw
2Fshpk6xoJiLAJzKXMHuBgoefcwxhVa1JQdANPRNSc4Tf7aAM7Jz2CTGCJ46wpLl
csfcnfewlt22UMZIba2Pyz/1+vSpymZcLCQhpHzp/G7Oy4wDS5syq6RpdEBBD4PR
7z6CI2mus6i82X7ydidyZ3tYVuDRmRPENfDmEkgXnjBmHz5KV2UoUSBeek6C0T6I
NJhJfkgjbxRjJxYMUWywUZ6YhMQd79hmj3QltP44OXr5xvkTZJ0Sr0OjqpN57hST
oAIJIVxtATiy5eT3rtYnyW2DBAjb70so2kPGfGdVxkyLCtJFckW33wPF6BDdN5Bh
B4CVe/P4/vYp5ZQ55hydQ/QLVC1V3ZdTlT7fuvyQYggBjzT6Ev1IrswXlDDyj9YW
qc6m65vweqvgVwOgEWO1KQ7OgzOcmaymJQQ7uhin5HvB2CPOGzFWkF22hEfXj0Fy
3/SXPqANuCRKqRDNShENJw40C6GoUHLCM3Zyljv6ePZD8gv7uvLhntU5BzWXQY21
t4J+b9RxFgO3j5WtqR7UWQdoUFonwSNKaNz015UrxevUbi+2W10QwLAcYaKrMbXY
yCAg2KYpSKS0yPVpyMOaLuW3TG+KZGMdFGaBEUHsgcxmjAhPybT4G5Xy6lwQLumL
gv1UJvWAH4juYzjG7/tDHmhoifFgC1hJiWpuedoGri5AQTIAHsT+pd8ZNCuinumQ
kXxjxgMC/4CZJyRYjrexP5MEVYsFmGDRzUMwCzqjHvo0CsyAQ2fGwEdwM+xwT2CU
9tbnrgs7W5/YVBeMdE6OWTFANh2emXnPfoYYM5WY6ZE/bMkIkDSf9/DDAAQ4dlNj
lj0Ek20YZj6Kw0uuhmx/IuCNXXUHhlsZWAPtu71fl4J0PhhNVSV/a+QwEwTR5oXa
a7ba9+YqN1M192M3Z6BcAtmgZWy2Q4asibqKGX8rw0mOILd/Dma00g2mBE4S6PW5
o+s+4kST3I7VDFWzcRHCDDAjKqEM6ky90h9bc9LOuphQQ5IwL/DFUdSnNovhqijZ
moO9HTIaBRzqh2KHIaFgevbVlkvm/e5EIRisDExGdfd2UrTdMl3Jh6PkWGbvHFsF
hlGKjNIK2l+fNjhgrIpZrh/8Xxdvc/izysKPoFZOqF0cXy5jhZ1bk+YbzQt74SRn
5HAIPTPFHhPPVqKGcDizdvrMD86YBzpOXgRnzloFfU5dBBFAp8m9DIRi1aI0hT1t
tYC7tO9TLIZYzYddQaRhzYpTz1KUNPmZ+tu6McPIYKPB4RMn08RTowcWDyERR3/B
+swaEolB2FChbuqaQV8vdD/Itiq3H3Ro3Zc3kvKGzHjiAVNRg/j1A2JcZ1evI1J8
1Q2wd7qRKvpY2OViAJLc9NoUjDiQ5r/HqwP7mrU0N1ce+4Zhdr3pcKQ25rcd7wwu
QWUuMYfCmxDuhseL0E/bW1+QpQ/SaM/rT1ei20w0XmyFgOojkFw8mij9NC8Bq0yb
ij59uhOFNFdJAvBmplj36ceTSyUsFDESulILvKWsm8Ev4ITJF2jP0lGhjijnVh17
nHSs777cQA5yFqj1t9jw3HxbMoGhXskaNvvzD/YCuMz8wqnF8KzP+WN8UkR1eQcu
gCo/Z+Ck5E+SBG31qz7XmQdGsSYuYZYLLgmCUa8hUnabDm4xTSs/fTzd9sNy4HK9
rvjeEG8cgIROShdULvPLg1zKjyqFtkk8aXE2+et6Kx/8Yepr8Q3nk5lXMV1bgZmt
BD+pzZifKShEx+GK5pO0PlsjA/AuzSEkPRa1oUxxbm7K88q19PGPTIpGr88IPDar
3LG8UVSV0vOsp4ME0lbvnPw7G8AipdtYbKILLta9sHCRtA+K8qPoGopqWxet/ZsC
EQVdy4mCsOPquG6pVSrXA05Irax7sb94qm6sSG41MfJjnSK4hYhuuVpH9ePgLdEB
+JUp4VQTS1Pbhj2PxcR11BXgEcwkXXQ6DkPFSaIzEDyC2OHS+uhXySsZIdYuJ06K
5+SOSfONfNWGqxisYEdSsRyh3Jw5xwhAjpvOXvJEjQw8kqfl+BP34T/LZ5ZxLP+d
Hm/XanQQUhp4QNSjIHr1UeRjDajo4QINFQWzcXyLqx5in0k4DEY0xrn9ynAQq3CW
Hwz4g98oHLsdWIAgm/M9HCCp6jJGP/t7r6hLSnDOQJQNdDb5vHRZHjKxNqN6pEBJ
oF4v69aeKVU9XSj/W/1antt1E6tdbkS3vmqI62MI/yZZk0rhyANzxUfCXMF/+e2K
W8r9yaxq9ex50J8vTAt4FCGhTZ1hC5eTdyi9or/5rNd25Ik2eXXT5Mgd7q6GqCYN
ROtTolqEhl+vWJzByFsYmF7dx+b7sQYjNj53CtC3FT+33D3Y25+v/TLF+h+ZD8u8
sEKNZofZ/Qi4fT7ofaWNAtN2slhrirx1JLxbYUHosNuHshcz0/Px/brD/io0iygX
S96xTCqPfAZ+w9VSq3H1EBnWYUaD7zg+zBlN/4fi8tGoJTzU2xrLtJ5ZEsDLDhz9
915RpY+FiaHGSw3/MNMM4fDza0Ni7CKODgHRi6oUIahEcHLQUHqN44ZnjummRLo2
W1LEtgLqdAI3WaN7VybRtTlIqtS4IJ0ImrjPvViNmxDbLLcH57YXA+H4/7xVMJ5M
gbrnmvVr9a8q2MroOwnndk1qCWQks9oAMf3kpCiaxrjTmybSveddrfpdFfDp6Yr2
6q68csCERAVamw88ik4szd7Sc8HLtXO6Ss00c89vIleJxek4VgwP3/6r5iceX0Fw
ud8TL1UNfRNzQATOa86g8MQaZV9RKo58ZrydVtG/jJPl3CmGDk2X3HATx1sTU6jS
6PkTk5lWOqdXrH1UHo6259XxX28rjlHw7raUeg4SVT19g0M47l2EL53AzzPnd27s
p+GI3oEV2H6xqqpDSs6gpePHwdAgqeEJgwLnCq28FY5QpiNTcp8JHUL6UCK8WCpg
Ka47NLxcLXpQj+Ego3egT4dhIBz4wY/z6L/YAZkfSUgVMue5gS0v5M9Mx1zDqgmY
TB1qEErlNoDR+ibieOKhK7rPQyzVSBeg9oU5MbjZ2klzC1UKT8Vxum1Sm0UbAf19
8oytBKoQXxgr4foMYNH021LnrQcniRojD3z/Q9DG6csODue76IZ2FHUh0dQ96Mct
bWRm8OGYwpSzxm1dEjxaso98yPpcHjX01X7D6BbBLeEVXZNVTtosOmlnhOhdX4wK
9X2y290l+57htMYTUco2+bi1dv2RBA5ekoNAU3C3sZQMrQcLJ+qBZsAczMHURqs6
+yakHmyLKFwy9nrld613CV9bRSGBnQCiMUFOU6YAlIQFkJvEpcbxQJXYSJZEpkeN
CtXXJhNTIIynHvupAVBGWhDWMQaVqes46AYch5n17M3UITSiJPjUA5crSHfgEqTm
d2ICsVN5g6JdESkRMtBFe3dxZieW/XQrU9OAhSglw7cc6KD+vR8q/UHS0pIaiM5D
TQEzsecA3wcJS7UrdRLkqt2ak/rAsMiW0QICQoJgXwB4JjzaTymoDQ1HDHjXm2M6
FUP4l798UDzjflwyJgZ0/W0RaX6o3HStsOpBU0uW7cv2AXdCE08d5sbHxSPcPoUa
NFI0msN0v0S6/VXJF4XWcR+4x/cjFcpAHQmFIeczE9u91TKwBl2H853vNpmTzUUP
ZqBYSn83G4JkdRt0kTMOZ28MLgd6NlMon/7jRa8qVOwbp0eiqEaNcHaO6VrBXThV
L9b7zOil0vn35IIMz9Hay2VKod0wZDzJoy4E4cvK+MIUpr5osO0r3OFsFHNFoYLn
8twJhv+ouPKO6fzIYoDhyl+HB9wAJhdJ0/Oktf3Tw2aUdVBtShH7C6AFclIr4U9t
AxuXF2fn28/Z1TgKAwwFmwU694fYKrwHDBI55ILn3X8RTQlt5R65vMO7COMgKXXi
igVODYem9znWGHMmxX3pKhZlnxQ9pLiu+VN+ndNHx58jHbly/w6M0lF0jd4UqEmM
XMAC8OzOyRatQCn6+SwxGRJuRtkjsJRSdSfZ41ZfBxPj/TOCXtF1fv5s/S+h+mnN
OpmbbmXfcJ74E/fpWipt+6+mKLfwub1Icdgyuh3F3WBDXUMWwCKkMSobYPy9UBkt
vK5dizNcQtmkBt8VdFM36yf9uu1OmlB0QFX2PhR+vIpmgR+Gp/mIFhMnKwyyFef+
QjsM0yWOIzEC7BSEyOIOOx22hr+J9kPb5GCSoNcJHzyNi78Jfr2XN9jZNwvevx2H
Ge9/s0yBuTTrEHj0msqEj0PEcBT2rbk6smGmsPP5xPD16FMICcwDifeKGAb5hf2Y
aLmeX6q7zqMSPy7U9FyjNwH/g41GWQRn+1Xs0ytXTUoUrtOY3rewUwn5FAUrNOg1
EWX41mOjkJYtkElp058PI/bnIdbukb9VCocmwPtxHoxtruEs5uTIIiIKS33NLTax
oTiewC/iBAUVzqLV122lU0BslTEV3/niJYzxnqLHLDnwDLlE3SBvVVRw9I1TWEHy
6I6CDgiFA+athwu4ewjDu8gSIq3xr6VWhkT3WzlwDz5iQGysg3xmQOs6dtw2qcSs
ngpcgMzbvhtBbMYxzllYNh1T/1w379QSXXT8rqXp2Bk/b8ypQxxY5uRsUHGOfdxP
7xNxbROTzMlfqd6808LoEkDPoLI7ehRaJsMFXqB6E5oD7aZFtaDgvIQyf1yBZkfb
jHlgvsN410Hiu19FI6Mtly+LQirlZE88TwRd8M/C3OEhe6j6cmOPHnv62AYpTaTF
u97RdKqmhHn2LpMUtUuupYzDFiDsdFfi8kklNMoGSkNg29bZMd9zAFWHyQNkodot
H6F59k/xD7Obp0KoPyTGSnhoh3fIK8d2b9Jtdb5arF8VnrMltudQIeqrUfxtG6pR
ER6SImojfoUIRAyiyOR6GPCnutgc1PTCpjhAAaGEh2V2JULVqUGBiDSWul0MFGe0
Aa64RXbFn0dlm5QOqS5OjcfGZs/ZDkgyKL0dhmELuFVtY7tR/qzH26Qv9C3YiY9e
odh/Fq3JG+N2hNIer356m8zmi3E76tcknlF0A0c3Ek8c3iNlAbMxbH/lpMT6HYSc
eFibEdGRYAj6xfDJZKUjzYYtv+elsGrMyoXZ2grz9vi+tFNkGQdKYc+LJ0ImWI/M
O5ZphOnAyZeuJ/iaeWsyclMZh+wLXTXpaogzrbZO6bGUuW4PZ/CuUXhEthduIHAe
wZGwOKWl5wT9S8VlMGJeTNo/yqM4Oak2T0qXhy2xww7KEv8FcCqmsZwTIZd59XzD
F5HND9BTNulwDLpBUduH2pGJ8wdzSuNUcBX4C7EazLzBWgxfE9Txc7SE192/XaTd
1pZ3T/2HUhd77tsuVKEnjvIAUolhXSoacS1FIndl8pDhuoUbzmfA60+RdGHw8IS7
fsf6PYOZXIP7f0oUch65pRq1+uhpmS7SDjVDjP4/+BDjt63G6pc7fuhCh0FnCUEC
+fStsF5VNGUgJgqHvtcXiy1tw71MCA6OQKALdT2R34Mcwt2x1aJ8lwzIa5a0RVEr
5kcuK+ESeH7D3YgX1N7FIzaY2BakY19g/guSg9595ujo9KZj4oWDSyEDnbOobgeo
dHJNS6pXu/M7ynyVrY3hRZQ3na5fKVWJxOlBAPAbS/cxXJmhwE50Id231iQHFwWK
V84usCTeiixZwFvrGgCEsR2ThyYUsW54cIiWAVoE3o+BupSvfPKZptbF1IOfyfM+
yIOT/nERHsvwOO53o0wxE/968eFRRfhfJ+FzwwgxZadYTolABkTalzqeW3aFwrkp
uErDVt+zL1k31kzZKPZuxHhAnaINvsK3E70HVYBtu3bfvH9es9X00UkjdxKbDpSJ
5KpUnkIOn9zdMtvH6IzIFmcKYhHipujPetoaAU6skzglyvx+P/7bKYHLdYv8aMoI
eM/HqXBWAok9kcMOSopaJW0DoN1JBzoDrnpbEvsgu4r3EOHIqnR/b3yGnQJh3sX9
/rJkfVJ5OTVsmlOoePpHPa8PLsY6LoHcqphYx5LY7izEs+nhU+q8ujbtzCfvBxTz
ZMX53sFtwRb8YXUt1kcPE4e+EYE7NEr7M6utUA8RZcdpZS+qOLZuklBfCGnVlipR
br0IdDeUxakoxnTYJ+K7AaCB2DFqtHsE2vZgYua1QBWjob7vuRLU6Vfw1zx4Davi
P6J/FELIwreIMVF/FDA3smtsf8jU+1aUmFsOsC0Du3Muw8txI9wl7/5y8uXu0S9z
M4SQhGi93TU/qWJP7HFQz4I1Ocoa4IOWlBjD5yCMdrOABr56sUTF2PCssqC7OSth
uU0kwj47WKdt43rUbVR4Lq3wK0IWqvdVOy3uJ15sCnWeOjR5Ubb+q6qdbFlC+PQf
/4MX8TqoQQX/Nc4wMQlaCOxmBGeGxOb2CCk4jX57445hSJCfd/TBbPViToEIPdSj
CxVkSSvexdP35Ay1kBAyTd5tjwlfjqIOy4nGbFoF1JJUZJekLhhe1djDNlSgTaET
BrG7baJhtPb1BPFP1IsS3AwHyb12eD6rracKltvLfrtniFwkiJ//Uzf6tgnhuuBy
czgIsVeLZ7FQMmAIkXunrNa02U9jFLaAycfwoiog5MnaMs5DLHoCTO/bhwF+czMz
mwtlJ7OwXAjmYDwhLfxjFmosX78HbvdGP9gI2/KmSodYv4hak5XAiiiM65IGd6kS
VuEIixoZYHZ4X00rAhsgA3LjrISppk/OqVuBHULZhAx877qluVtp842+pUWnyWtT
dkV0S0xAGykLSZTriSqlBIIPTEwyLjKhvCAYlU2YRMWe8S8rYN/W2oXL19WU9+kQ
PK0aK9fG6VH5ChCjATXVT0aQ2WJpiR/6/+Y4aqjfOo3Nmbnm1A8gfkg92McwfthX
NuB/jfBqPIV3cIs/q3qlcHPpTnqquMRcCAaMMI2xHt4dmRsYpDA3dnxXcljiTOn2
3ANADLZ1jrTt9G020KDSQ/KVyvpOrGlP71fDGjx2ClBe1hOifCADX5IzTZ+27Dul
1PNCUcxFK155NKrpo90HzBeL867BUGKPddbA7+lI13cXNlqLcqDZBSYR4O4pCI0S
sHHf4msSAerz/mt0zPOoRxeeYiW4NqDlD6S8deVWb9aSecb7FEQJAgM/EJa927v0
krIcb8+YuF94TzDHY8LDRbIa7iMIHLDIGG4I09+0rmT00WOdEP0ftgCOPBqYvy1h
bkCw+48hEPzWHxBL8aOCszYqupkadnpz2pOD+kb/jPnoljbnLrtuVFrbU8pRHzsI
XXJ0XoG19j/yYwHu/1hiHeyxvdX1VY+L94C4o3pQXyFm9SsKEpPp3ZXNH5yLore6
STpLmZucmYpSE+y4ZEcGbf9X/z+BSMgGtgd2zvlr9e5Ek8rE7en6/jfQBWKSBspx
2CSEAupQD7wc37DJRIOIQOYTAPVb9AY/mkffJhMDTJh/pfMsbWtL8pR6HBcwH57i
V/R8qAcd11D4jODX9aDozOkj3XNDbvCugltpVaiVyH/ZakvFUr8UqNmPu8krndSG
OvjmL3p+yBCVE0qZMPjnUDJw7QiQlplJ0ZAWAn58Non64GSKCEK8ulq04REEUBEk
G6fe6RTWNHuZY5JR4HuVwMGVvFxGx8O+avJf5sJgkoja6ge1gxlNM0HPdwVBRKw8
NljN/xeHWo9HkvPHCgE66pgQL79RDqUvqVfTf8gYj3gVEWhZDJ8ASdIvQaJEK5EQ
2gMkOeBkAAL7BPDMbdbA6Hv5qAT9XR8UvaGcO0D4ZsXg+DVZdsxScB0T3SfUGjyt
y9GQhGco/MQYZ+QNNMx81Ujzbw06lyPIN594KwH0J71OJXjh8D6K9qpS/VmLc02i
DDLHGRUBrGVktg+iefsVraTE6rnddJTJJ+3TtvqGZK4dz8PNf3Ekl3UeiHmtJ9j7
kMYUaOuYG4q+m6efCkikzFF4UFrjWtSsTk6BZNqGC4Koa5wFimKrHzME+2Ktytrc
NRV1S2GRQydAea/LeCnI4CayqCLnj5akTLWYh3LuzlEwkkIufUc2CceYNq332cQl
Nd2LQ+IFqRfmuM+hA17E08lK6yP+i+ttA4ayRe9anLlb2F89hVeSx24pti1vrB5g
I7AIGYOm1nkNFiDorn610IC97m0Ubuo7c3fkmzMYGW4HsKZjpQXeYkJ2OEBwJvmk
Cf6Dk2u79MsWd5cXr9DtoELbj2Qjx94lwFBNxKhyjVSHENp/vj/D5g/wwmAh9Uu5
Es3X6tYRfZSdhNujLOvo06edSXctG1iNvWVNvqix/b/BWOIK78ooPxlAayne92el
TxsYqCG4cPnfLdi9LgfXZHLHYrZ1iRLrWbaMgWfbjagC/JJi7jVxGhgmDHP8eQEv
E/7aMXatK3Dk0NP52DTpNVD7XWJuxXXf5cCOMhe47K2Ic6LFiYpio/e3GMuem/Bw
zxsRsbDH5MtAmY1y709CfjPEP7TiNhSQWE7LPW2btA8kOF+4ee99Rs/1iXLxWOGi
ZvtFUDAnLOL7VWlGtJSxzQsrQ+07brfwiAojJ0K+Y3u7yOaJ6k5oS+BZoug/AqFD
VZRraop54Tefhf6gA8b5oY8Z0xoj0cLxhIoubsX3I5/kBW9Ox1R01aPIfYlVKS8A
GUKUINnR1s+LdOJgLUkF0oEfrdjUI/KQ8kQmpTZ6QTJSzULnvYoIEOBur63g4Whz
cUzxiYNwHp4oWo5rAU0ogAV9+a6o2jcefSxOQY6tuEltlQraqVdMfVp4EQ/tI1Nq
XWpmECbKknhrFbMzkb1UH7nck9/BhCpdpNUSI8nLO/XCSHs9uzIH6Qb1ocj4UHIi
TitOKip6VrUpeGqWHBeeTxgaFnfPosQ2gxZG1z7ACvecFhiE/cSsCvzdd6nQTZbK
8fmza/beRhYWElgk8rRWWVeaplb6sAIKBmWc89qLLVPTsHb+MB7ZlTfDDnuXP7W1
SMrq59rjUP8jt+DoJK9THfyf42d5xFylGbO1sWz3yAc+wkpt7iM3lh6c1CfwdTSK
xoOWyJvrRSXrsbYv6wFvATAwYe54/c66ObETJwtSuQ20jqk8uYHtwN06UuIE+R1q
QeEkAeOIie8GJicrvoknt7Ut1acgMSi9vdxBqKwPePxvYo07algU5dMtUXA3Oaf+
/UDM57Fdhq/gLwAYTN1Jz5Ci/1z4LEzyBDCWx8n/si52RoAZhhbUHfh5te5qipFp
1qE459rbpcalBH1gb5iHSZWqn4fi7DBNrHeBYW1jkRpIxt6713qaDLeKf2w78x7K
DlKv8zYbZuzb5GbaE0o01jzVtEJLP/wo/Xj6B7RJNZnELm0fC5UQV6epndC+5c0p
8o9wRBDc2Pkr1L9UoPdYmr/X3hGgrHKBQQw7W6q0YgXwkWkYpP1Uj/hRJPU9IjIE
pwNuJvSBewHtoshU5iku8BkDKCrKskn8WsIGhh/YlmWIZRTQzdbbcEQSa56qcqP/
wNVE3d0A2EWjJ8MZSlNVjJM8WBi6Zf/3SzXjMU84eZPCeHeAFw2ng0NBc9/ez3EC
BvaRkKzO+oTAGHPR5HTo5ip+C7qxi5OQPIGmFkJwjcr6a4BIpAy5daYdS0KB4NVI
RcqMI4jTw4ZQBIh9wXwa0Q95VSBpKq2bzM7qziioZFQ+T3pAWJEcU3RB6mKFW+Sj
XkmUD/u4IfD1vCiXlPZnBdu4HW9u5n2slQdTIr3HYVhe+EhGg5UcsV1Q9aNVZJFU
Bky+lLF0QjiePbfVRBCDD7S1PgqA6XseN+xmGsq9C+y3t61WDINy2CY44Swmiu9V
GNnFLnZMWPRlPVzxpZqIs1tn9DWGVLzwlwmMz58Esy7agZNlMwr5QzOJlYixEMMk
WmCrTTTjpxIW9FqxrTj1fsxqIAkcjxWQDQF0j1/8245UQaTeoIJ3XVjOocso3LDJ
aRFUKMGwGGdngm68mIeVkUyEsBYoL6GFcD2xNicMsxINzEdT4RO62WthifJbfT5P
WXWXXXyTeOrOzz7XBsbpgTr+dJmui1PBbYPBbkwsWCXV9SSuoc1WSGhfFkDz7sRa
bK1WUtM2i1FXemDqrxHaw6+7VzTQwL00tqbjbTo9ZNoUeuBfQv/tgsPP1LtMW223
yurnUfB8ZQsue1oFErYomI2XrT3fzJUaw8ptUJ94emusfYn3XrgESJP3hhiObAjo
e1vhslgvvNOvtPUTa0nWG4wKYyuJG3zdTsGzI+KIxOQs7kC9MDaq/tLXYFhGBqgn
Onp58z09u7KxZxRUtSMBjU2W+mPVyPLxVM+vZa0ktQZUOydfu/cR2i+YR7C8xesV
q/sfcZ26rQTKZ7Xt/qyOpu96bfMJBsh5NJMl3nsCKn0hJ5TkjjtV0z7oT5ZA7bwo
itqkgemJyxWSBP94xDOAXWMDPsoXic3YjQQR5nP9aqg4jGLwNWZKkMOPcx2TGHTl
GwzEXAM97QIeSoyPfiSpnZI2s5nARO1tVztSdedcAZXFndmNwC66YktUvZCjD1Zz
leaNq0T9e4jtgTAFQCBqQtQohF3NA2LHofFHzRagQd/TnNiSvaocOh5Cd1+YiG3z
TBCpMrl+PUSgan8AEjUZ7xf6WUDCOb2Zi6x9wHXfFUzT+5XRQX/0qnbJ8DZ0zVn0
m1InbEDfj51AeLCIsr6OPlDZXaV0hwuv25VFoXtC7XA/KMueHGfSC2B29PW86LX9
vPCBMgYOeqVOW42Fl6Cj8zcYbFmSoikS1OtF9IgAucemeyCB/avSy+KgWgnZA24P
fIpKrIidH2ax/KCJsYoObKXLkKcFewIL7TLjRNA65LQBbLIt89keOlg1p+CQKSCK
3sXR9tIDThZOFD3H2JO6LnJBgAMZkczF7l9s5H4Q8PjLivn1zb0nwQa87yoEjhC+
oRBYE2fTUuI9eIjqkOQhhzIMtfgF8wKeto2/yoyrgtROBgQUbDS3bPd5jgQ9Fnwi
KpLAM7w83z6J02wIaJAgwNEaxv0lxqRWBcBFRON7n5KwD4KHOo1vJ5SBBZqk5WRI
64wc3uELPXEFp6bfb7oP/MuV2/0/FK1mG1PFkpvIAX8wt2w7fpWHRwlWN90t4OdK
vpAX3ClMu1BCmuTQqL3gPagKCbp9AmTbdScInyHEBxhzThwko4JlBz7H6H2c8bVR
A9BLup1v5jU76eUD1Yz6Hw0XvTxuI3TL35xPkTUxpIEhMzt8NiN+RvE1bMJ2rftR
dgoA8LYLSqZ3VUqkm6FpkD6uYxMYh1OYG+o3nLPwqmbAFUzFoZXu9bnCZXRArdsb
hFtp7rTfGDsyltEpk/Gero3UKAsFQ4RRRZk4Lf6URoe8o0nJGflC76sU8cZSshJ7
W9vZsyTH80UbRuXsl3KiGTLXVrnKNWfQKuPwcOJ29vdsZ9GLeyXZxZCPBbX7j6dG
VsHr3kdT0CLtdfuXJQSY6r+0lQaIgIAWsqOvmaMXhisFSm0Z0pAzj7v1tpl4Q0AP
9eeVyblaxXGDL5dglY9Fbj6pEl1sxBs2sciLePn0BxVTLI0yADFj2PhKcUcJV60+
9xJvcNSYJAMCmYs6eImL879bcEd7kI1aODOCRhzp44uGqVenAv5EMNicQLvPUhJO
NEejEJ7UOTUAiTOp9I4k3cfNKuOqnhKmcX8EKMn9VLqhUjKWk7ZY7E+hgkbma3Aa
CXaMh1GNMWn9yA0oT1Fd+UHAapilIBdTyiOECUQPFxqI8WrsFA5EovSAYeOrmKWr
ReEWi9cuS6a57aK0qwWPfxKYvcb9Ob9EIGLueJJGbCHdZIgFngGxEjnsmXtSXG0w
JJKFA9bgLSXrFDmbQPcwRrBtDE0l0akIxVmXfXDp39zowrUb0vCg4fknuAfT0Zvk
JxyCYW/tNgRhhnSIJ0wFs6E+bb1EgmZMoWJ65oe/I4LjoNFKJnr4aj1lFac4FdRx
kstcHc+H4UAyHtThoNvMhIxgo/HZGc7y8Blcn98yaGkEqXT+HnpEk3i+tWs9jbRv
2RFrMcPhTno8tkmwBZnrpUUsT6ob15V5cU8rdYeMW941naRXvqsMKZWsHAdyMpl3
v9h+uKtLTvAL8gD/zbhyW+AASN/zMi6FZsjDdWTsXo8gUimJD9ojgVmS39FtdqrM
yQw8OXMHsi3RI+OGKZQ3a00PSgIaDUAq74m9Va+2RH+/ULkP/7dJ8ihsk2b3Q2w2
+dPfOpHSoTZW5jLR89gGBPYZUWpPla8i1lrJH8KsjEWv0bj7YB0vdL+eF1OGJFGI
bKW6c8gMt8UypjWctfgOAOTZAhb4hXmO/tQrVcUU6/mBLZHIzxhJmf3n4LWJOTFU
vLd5CJIadkzdj63X+SfT4LBdJ0UwVpWK4sLnVyW/IbwTBdD/rbJ1n2ccwyF28+ff
4JxRmf+I6A0zLq5dCRG4Bw040tjm/bBibr+FDNf6VTTBTduUhJ169/e5ojdxq7Tx
1p9YStxeEcTq9jKBAK4tlT5E6uX3QeFekjuPVUbgjC2VNc+lhtyR3+5x5jvvgeO0
cOzTHtp4NdlNz3+D9NG41TiKMwcRuGot5oj2Uo90rHTTmGRioiChETyqVVlxpJOW
Pvvt0zp+Zn0+MOcr9Hg0wNOIvz8F/aPxsYODwE03cgIK4F174n9Ybp8ob2SRonud
bRhFFFDI0NsAPqHTgxMAgH8gDaLJwQ79LQPGZxQjQmlSJiYKz15waQdSOO3D746C
HOKn5wfr4OJ7bVtuONDFA+ABRxW7fnVCzV3RYsYL27ZNz+ULXsLHn3sPovGiOBDd
90EPpTd+2R66ejFDcAgmdwknGR9b7/MTFcntD48dndjpFqQCkHShhvpl/aQ0UdFz
6pHuD0jB5E87CMWUV8Q4LYgTj2DeBamC9BbR4LgdYXZWc3Lai5Odm4vfllDuPy/m
LoWNQMRMQdT6l7BbUK5DO06K0caUGWSaqbLiZvI/1UKQaomkt/MQobufGsfmp3cY
qUKjgTP7YLl6eovCVaExY98oaPemdpES+aQ9E1F70fNdEn6pgtnphiSk8DU0U5X8
6ttQf5axt+zwQWV+X/Y8k16Aqy7t1mmvMDTu5xWbxSO59q5t5iwho1IRq+Yqiz1H
4bd3jbtknkysrX8h0cGLMpe9qGohJJQUGjNPQsfWvtkTUJeV3Mq3cjbIdXcuMD9N
4lxyi5NSfOqSgkUbzzDLnctd8rCYfQr3T9rzQbjKytdMOtLCrtAId98R225EoJLi
f3JG9Fng0PmEkRRw50ALJBdFl5P71TK8Qj9Lv2oLVBkS4/M+KfJ/EAVix4x5JROP
M/NEoVVg1GwGyWX4bninsaLG2IIiE59dOxL+UpK4d2l3BK7b/CNjLyeUXFxBiJFi
kV7ugvDC9L3i472MPomlPpK0jsfiUmQhWlj4fObx6Ag8zt17UlSEkA9PLyImrGu3
EZsPKXpadfRjr5RT7ZAOxEmuKL/BC6P5K3Y18auRYfFhFKsGShRSzceR6UFhQU03
w+WG4yfp591Rdwrpgie2YD5GZYdg+ceEi6qKK6QWkaAtqNsOFSdUOmdEZdOdJKjf
6R8jH65qklr8c9tvId5goFCI0Nv6JkwbrHTBbwM38gpy7Ar3d8Gx67fT8tKJK/pk
wwF4SN+RoWTdQqwFnpeiVi4EtMSadNbCh3Da12tap3z2xqctH8GByZSXgNYbmzlP
jQEN8OD1P7CWH3LtpwDULMQyQwfYd4qFLkzOFDVpe9QONwVFt2191+Mj0zrbWnuT
EkWPh2F5u3RdBmeRLyYGfVLKbJBaAt7cMYl2Z2XUt7j4KMzH1G75iXOMdhXYctRU
J8polVO5Rv3chkQmIa8Dh3252R1/vvlAvKXWe5FnDi8RfpmFJm1cSZwkOEBlfzjW
Gh1qsURXCUdnip125P4kkwHq5KqCoe/nQkyreKXgul3mJYiW2KkuqAeA8wzl73+V
To3NQwtNjwE0cp3ZFMZKZuvwPD12Mdf8vxu4kWQeg2XhHFIHRmZW5ndVUXlLG6iy
U318b0SZr1oNkejQdaCHVWakQEyZYghOXjOLL5AKAicQEyIQWQX9BXiB+HCwXgk0
yZgDNhqE+nVWOgiFZzbFZ7mcTh34qggnkdkNiCZykatKapGbEwrDZ0yC5jXu22Um
AzbCqs3/gj42aUK4i0KfVXmHUdIKQoRyh7uwNB7rMku7F+ssPYIgTvP/JyqT0oSC
OEo5i1c5GQFU0fqTyWkhHsbfDwcx2EYZt/B359pdmrDq/lPRU3HzHARd7s1ErL79
thpUZVJrPHP/7cQ+sPHDJmUybjs9hoMen07VKxd9RKOG/xSfpjs6E2WIbdcJU+Ph
2KtprKW6hO4wmJdVLBk7bBGlD4LM4oYBGf+MCVq3AfwDCOrXe0QOvvKkWZ7Se6XL
VnudneM8bbZQsNTlTg7VSZDVP89VpZM1KQdkXz574tD7aa4zDURLES7E4F4xfDUe
jbXQav0h61ByXETN7BIiAeCNcc/yB9vB/UrUtz+nD8Iwfdv4IyCIr6QP3Ca3P78B
nJL/+2WIBzkSpfoCQiKdtIERKQqjzygtyxfCuBmoUNfWqsFtRu05Lbo7ZjjepTVs
evWCHJ74np6MLRukHG9VRnWeEoUqdPEO8nBxx56Sd9vvkZgi4PYVmTgFmjFPInSC
j6rsJDbS5nkCYTRDCVCWVhu1To1XS+qfd7z6hb/UrN5iWiz4fJc6gyfN+O8KATxo
wAC7XNAnHQtHot4f5Ltncoovc/SOoq+qOkgtAE41ihSZ96o3NHYTUN5gOJ4rrUvg
XR2ApZUibQrxlzwtymVFo1jE1s14XDhaz4UsIaA7vLhrXtsMghoKSRQjPi1T8lAd
kRMQLW+NHrmohzjqBCbjvG5iT6nxuz45QYVC2QsL3zBvEumRoXgswCpjoJ5Qzx2W
Wli+iZZ0+pn8CIW3prYHoppSThnQVAmqtLkefn4wXmJeJp5XY2ieDWxr2DUuLOPT
P/jFKvA2cS5Rm3lGioNKeqLE5Bls/DUlfIOaLJqtD0KHMgxUqIJ2qSNjGOmuovCH
WDcG8klpl0AHl2mwrlmd5y9wf10o3xmEYmCodiosKa97363VBaq9V71elfLGvFCU
NcY8kf8e1iPydkrYKJXPzvKZryy+CsT680iqS70vhHGweDSJKov96iTk/H1LlAEA
Ato99xWMfTWxQSPeocn9UubGCedBm16WNjD6sNQcTtsKj+IVTF7TsjM7SgULDyDv
hacf2n2RsQLmx9z0JzFBE/cNQnmTjcSW/+GhCg8nSeepnt2zu6ygXMEVpQ6nRTXQ
9bjDrGwpDmgQmq/uqxUOfXReBvPK0c24IaKE7A+FAMvFUs4wEHjueTEOPQL4SU6j
t/C9nyw5DIg/dHcMG2RTNz/MM6x1BEDdHqvfq4QgRMxB91M4D95Q/0NQM5Ukoh03
kcKSIB8N2fkLcfR30KHrDZL+2N/81bOvNALa6GCXQnROgsg4OXdfztbeHCucrHoo
ngBG+zaDPOSDT1ndWv9FTlta/hVoSBZEcmgKm/BP8GQnWBv9FnqEURY8r4Qe64n6
Xjd/fmKiS9YxRdSzTqi/j5fBQcetnrm+jtrilGSBkCMb06dOdyKV3Hwq2I16Z8Ek
3/SJ2nqo9jwtk/f8RcMgstFXI1qHjgJcbOji50xlGsvKkYaAW9oF/GWNZQBqcZwg
9vLy8XIgP1XOjmm7LPEumLL2TOe9PsvQYqdreHbpJ3AefjjKvjR6BdvRPcS1nmRN
W79yv7ODx99UAfqeSjcgKVRQuhrndKo7LP8NVxL3pgrzA+SLMDc2nah1Wl//2OYL
nAbnKQ1GPeSow9fdZYUr9W30AL5gM8K3Tul4LPQs0MVMC3BJOV1loHGAvBoInm4K
GSws+qeyimj2w/7ZiepMEJ/NN4skvhheKFXYab0txEpMAFjGAJtKfloM9QeEwN0f
KXHcNb+3riH0bsuBSRH8R4YOozpGXivxh5i1sQjVKCQPqVEvXv562mCeTJfd5FVn
jYWj6Btpxve13ArvnrzMRq6KuHkpC9cjL1gh7anrefxorXbWKBxtn3Sfy0YUPJQy
lknSyaID+/VUgqhsSgtatEcKjB0sV+FVQCWxX3qqVpiE/6UV6IFZ+zBRKK4Ddtyy
i9nIEJ1k/fpb5UamSP4tJfW5Sk9Ab6seN6kqav+1l1Rd5oIgR7mjr5paYvrmiceY
t4xi+1Zddeb2cmXyrpPlud8rcm+c3IAskSi+wvFScBHjsVlIvsBwrwSNBYn/I3th
V/FAnjz2tvc1tBsNh7PYY+XxNgEuvPa8yvYJpy079TdfeBG4TnnzeQeneYbrogkp
8nFXX1mSNzWecEg/qsyF9rWua5EOD3NBmzGPnVM997YYB4y4sr4xX952SBmMA4Xw
gBO8UDd4ihArvwXhITZjooTuTTJPz3GzvUL1iVn5L/3n10/qS1HDpy+JpWVambrY
3uWoIakjpkJFxjmi3kK+7IlY0KqF96pw0iUBoAcHalijrlq0MDl/33C6KQGMeQqa
xrZzNtssf3W1vijfTX35Xe+8nN+ersjRB4soRiQAhG6ZmTmriLzjjLz0P7+YZkQR
Ggq/e7e9PpHa0xSRHo2hookatzRmhRxQQNfhYF6ff8jZ9tcvll7VG1VmXRgrc3PG
CQYXIE2KTsF9MDBL4NS560pwlo3EZiNoMabeuZ7cEfF6Li9HCH95O+ldEAXJo881
AHHYWtc1ASKrNHrbminQ6yEdvhAIXS32quHMikLm9Bn6HPdYOYteqcILd9gzVEJB
s2pewG7P/hG+eMNo0AuPvKsxKMLIs0ZrrD3Kwo6qjSO7fU04B9MFf+cgIS5/66hk
mX6WS0lbhLEum9PT4BoJvoRhGiNTTybh2IGWfH3h13/qZA3REc4+8ZAmUIK67zCc
k2+eba2SiMGMLWKLwuoG7W0MqTHoLOE5R1j2EU/whfOK2sXEkkXAb+5Mxy2VI7Wa
eandNbpMSg5HUaINKtXSOffzT1+u0NoRRAS8Csgm+ROKvAyNoDGKSs65pxXOYUPh
BuxB3bUczhxeE7xtbq36h2+3eZzOK1IZ0jGCh7CeVqGIKLHmPTUVKlLc5VTHy8DP
f13RCyjc5JSO14aTuxU2U+JYwtg8zPhhT6ysB4Z8MYZprrtAGXvf0sQfPW6kd45O
nJY0cjUtcoUd/MOdgH+vsvT3dErJFB8kiS28F0NVgUKkvpksmcctDOiIVD0GmqkV
cnmK4ybHswTHPRA9nDadiJAeWgq/lReAL0DaPBgFQxL17KZ04S+MGI7lzG3xMQAp
DBU0IReYCGo5NH7bJgvJIZkPD5JJMHqipW6uE8GiCEgV4YBCiKa68ngvbYDnlu6F
67/jrSVb48ldVp8etFR7UvQbRges+piIoI1iATW+L7hAJ6vjt5ySGjRag7588Mnh
TDjfGPdFKyFOQoQMljm0qylF3BIS5cHsXJ24QsBLR38y3noQ1/IauBuEaT0AUPbl
UvNN8yHvEluudW7uHWMEyWt5SujocyqzeCdTlPINsnEG1ZEn63F7MNLE0HuqRwBl
6+58oXbL3ZT6vjszutowV1dBtGxhLlRghMauEtKJBn2JhLhsg2r9sZn0UuwTSi7Y
Cfpn0X4Yvl+RzKKcQLcwTpyasaFkq5sLYcoR3l5As7Z2YgCoIvvIbiE6ZUQ2fT7V
POw29+3Gjw3XE9/s2NuuqVezV/oonSq1wcNGqxepp7zIPjzjRomLCZH1du2oSKa5
wZCUQllxnbJOBX5LxjVTv+Y6JEuaa1KZ1l7K9KZGE/hj5viSx85/yUzeMtVvuOOK
0useIHDYqIjCNIOnK+7woDlL4x2z9YIsSHZDQmmIFq31aAfU6XmcyQ4q9TXBQZxv
pwxlWPOWxih4ZkA6ECxR6922E3jPnzMnc3CULRF12kIjfHijFaRghGSTS/Em8Wbz
jDBYcZoZ2oczGkqDMELwXXmxBrCZWXlFyhnzBHsbB7nQR9KbPvtXj5HFC+zlJoXE
7raMGEMP5VUIYfVW6/aJgzhbtWOdsPzf9yWQm28UgL9H0VhtKgxgHIF5kGp++pS1
qBilBrYnms1LkJFXJ4hnopFoYZexBma1jHWicpk+tu9BSILthIubEiTUFVaAhXdy
uPw24PFxICMFsPPSUpgUp1qZABxDUbISjipvwpcF4kdrzJtdD5NjXyE/uy/dYxbG
fh6NVe83JINNqVAIrWt+XyfZlJo14J5PVBUlGbcvyDXwNiE9stN+hnD3VigCKglc
29U2kKGlyFBUMwhnh7cPu5EziDekMORm1jS+BwEMBr2AUrcEdgqW7cFmfgNRmYz5
/cPQslubIwsL7B2fGUzcgKJHfrt6x+Vn5dFFfIwuNhaTTPxK7y5K7VEBAnuZ1//A
tAcClLEsZeaEjymPFpyJVPloKiZnbwJErTw/Uv3VBrkNGEWr+g5tZFkAMzXjl2RU
zGgADfPQLrH5OmhqZmE++ue5WU4y10L0psrpOVqxLNCnBz2Z85edl93uB3rXD6V6
+h1nBOXX5P0OkW6xwdx4fIaaIYAs7naHJw40Y7SmMex4m4HKzHlkXRNEOX3bKVkY
dtR4rBHkWMDMYrBgqlOBigTZGdByZ6FndObAnREZZwkHptHJxvbsHqhXmwcg9Kok
oX7uV8klKJNk7hw8mp+ToIHi+0uKafttf2SlzCGPX9eyZcjhb3V4w5+GlIHJEnpP
0kNp9DaQ4eQcPDl4neaF9OKuhtoEVZ4ELZOqr257MhHW8xTI1NsmEvkH/y01SGEh
u6p2xZ4p0hW1VNzvNApLWiwFEDUY4KJJnb9xFkpivF2Ii29Eqt78Klkwz00pM8zp
dexQ5EdAgHFd1iqSSnQwsPgoJH0+uAkQviq78VRe9x/10DMeldTPLnZmok0x9gXs
Q7cuCr5RyCFHjqLRWdq2dE/b5SsZpE38SjakRO85RNyJ0BUEAChgxQDxNVOv/0+E
Go6Q1s5encbAl5dmMFzRJqlXNpd1saskr/74/8FT6du3lc6F7+C+L1MmrJMTchB0
j2vvpBvFJ8nCVbmgpLtqkdIQw1WlhR4YjH1kyC1UO76y+uGFDOG4mGiGfDBm2SkD
MlC2bIvO3QV07o3tErHVCX9byDZjpsqQdOMOvaNrtsMUHgFrwXunk95U1CImU5dC
Z9rtq6sOA1AQTMYw9tGwryXxO2uIZxAZSruP3pf+XPL4v9p6X0DUuDOEOIuk+kQH
kAyjtMWy8UwTpqEUj7H0+7IBJtrDtWu+ijBzmibKCAeDK6IvM2KI39bYr2Dbxtef
vHIy6bMgg/BdnNfH7LFMWCeD6/q3eiICmezmCo/rIEqO3mYZYpNwRF2EMC9fNlzl
vMRA/Z3CyQH89i+1SJB4OHt2zPlu87ucHfeIHUt1HWiQ40uJTBLkveNLxodrMzyG
atxwJy+ghe25LGDndEyZ8g2u84iBFfJjvU48w8mHL5rjqbk9NlbW2m0zIscVXUMV
k9QgsNN5AxGMZpRUMRx0zqVjiQ8kMvjCEgoOk/5gbrhIzcFqeQPt5MJ+tXjeGG6N
tezv04eGm5yGwpa6NEUGTHN6xsUn3H5341VdGRFdJnUIAnDsYVN+YFA8SDQs09cp
ErOSRymvVxTDOH+QTtL65ZcjZdAhIJxbVu9g80L6+v1OmxgejwejlbuZpUC1zX0l
PzjLeArlYKeKgO5Mb0fLn8MnkntrOGF4F8CVcVTb+FE70yfLJKULGiOwkU0bgxJX
mZMD/O0WUm9m0I71KBOhV+Q+x3nplUiS9kQhXNb/b9Xi6e0CqylIjLp2mkwfxQk6
zRTaugHJM7POYkioLyXWzCoW8FYLISij9ltBCoOvlUFQdU6ex2spAKIhaODev0GF
v4VR7PHVJXl+zUH4pauZM6PPBfWzxKwPErwnwV7Apcos3+iQV4oIQZelc9BAIFhV
OQ+T8meCx4ngCMKoTNMSKxHKC7xgPhmf+d+Ohb41RdEoYv3FS1dEmV970y6FxOzW
ZptpI+AN9CH5CXQu/fb1yFB8C/MUNPhRbiF0/rxEJmuvcGtCeA051IwafKoGfXZt
VQflwsk3e/89BFVkK3AAApM6eGnXDkD3qodX6kMiIXEOHxw9Oi64Nx/5gZ0+QYaf
OEImxXBssrAlKtWyMwTQwldAJTeVBVB5OzE2g2Mj0edNDXrhVlEVFbUSuLZ3XgXW
SpVGTOKG5zjyPq3kGQsaQFTwovFGrBQMiTI/3pA/xDvplSy807Ibd1RLui67LWSV
CAb5t0XDQBZVkrZI5FXL5UldAuJ/1R6gjPZzw7uMSGH3H+5efxrRphXNrUpjAWOY
Y5fdWVo6BJdsAuFYWouVnK2Kt2F7nH+yJv8eTYMlQidDyKm5us0gjLsJXlwpb4mR
vyY5OLsqZ8h37adG/KuCOl1sWKmolTmTS7MDdjI4uW840KbZhsqwphpHKFXIEKmd
r+5Vc3p0U0/Xq/c1gRrqcgbbYJfBjzDU00hwtA2wNL57iEL9X4wtTIZcHfa30hRO
RgUguCEW46pdoxs4JtMO5cPCekvtbc8lJREEgR0gMzdt0GnfOskciSvfyt9jNqtM
rOG1+ZJJgW3ThH+IDJeLZFL1MEyIWieVV7LGy1WY0bNGyAGF/wKNa16SJV31OQVL
/zuYkg8k8zoLBWqzYzhV9rscZBY39DQK+OczF6S1FUVpP7msn2JLd/QU4MiY4Orj
ODnF0o4/5HoaDpuUt/Q9x9UNGAWsKviiOhd2T2nwcSVB2ojF3jCVdF4roKkNkNUa
dcHXCDqp2vdyxE61yhgyEHZUZS9GlIyIP2Xt0AH9usD39w5KT4fg0DevM+y+7xgJ
d1fZKND44K81XupKWcOZvyHa2oEpplFqENC1/7wdi50sjPHRoghyDcscaLfY4MiM
uJ+32wjnyjXNI1cXDKY/v7mN98OrpW22+SrJZKuKlxaR5jG4vaJcodAd7zEBRiWx
BXTNuaRdjX1+l9g1EEtye6Nn1L899rJhWLxOkFRZ+vJiKf4nV3af+stYpa2gDASB
wnjkEK7kaEPJkrJ82/Xv0bkbaJ6mZxFy7RLLg6L7nbfNfe8pSRdCAuDnhZWMxdvw
Qfb60ImYLs5qQLHvxS29TiDwsR8WS+rN05X+DzmVsGEz4UATlI08dLjUmblONOBc
QS115aSBsYNH5H5o8VeoHkOQngA+33GS2S/3GoVWSmG24QSWC0AH8wB1/Kdy/l/v
uN+WpMKGi1UboYX5e0FeHz3sUA8GoRQ9qbRCC36BJlkdpYOMGFSKCxAqxVHlmIQX
GYFdEXirkXnFLWPc8IWxUDop1j32UQsUXd+a53l0MGZuc9+mJYuwfTq2UYnufXyx
5qDP3uCn3ruG5MwPUF6RNzhfYD/vRRRZW1K/VR86wHSp0NznhzxJsZBFk89jQTnB
eZwtaYUIQRMzVhicdIAn/Q3a8kewaL0S2K64brffgBggInwojFZqIQY1TQ4yzxWF
A77pMHbIJgDnXkp8udWxSeFdWMyrnqs1Fg9x2wnvueJ1CS0YrmybqVgqGC0XxwCQ
iMKxP1Wo+Z+MVOgyTJ3kKqZDfTHnjkYzOMyc7k/+X3VKxgfaP/tqlPL0D/pDskdO
2aZK9IPxKpG9hB9QMGETxHn673E9OarZw9ooXDeyO974FHXRUALaPo59ZGLMp9yc
PYNlQGS3/cylHA26w0xwJLR8BQuo1EgVYojewec6RLaZv97yQtXMn0HXtNuoufzG
Ej8Y+i0W9UOWPkfJep2k6JuXUCr0fWuo/e4Ym2Jspuz5sq1bCSWefECpzgoDDcAd
XxN2xepPll4n1vRBSkftEcr0I+dgA95VdvooQlulh3HKe93a59eD+uMe80JZvu9g
/c/FPy2HdQAzq+cikR10+VaVQfIH9Tn08p8Xnht0tW/lh4Rxw5jHbZ7+iuRv+0lk
aXxvMVf8kYnOASzavItFy2WRQWc02tQJgdzkcog7vGNVR06/st3RhQ6Rx1A2ZN9x
hdtwJoJ2owfqgsXBgxY09UeAWtrZlQ5A19Cd+3kdOfuiH/v6VkcMH9dR5rFV+mVJ
QiHVBhOt4k4jJEUl1+Pa7QWtwjMKm6lTSNtkmPaTZ6PU5HgeokD2AzMg8+VYLImU
8Qy/zTFDbvs9/iGnUm/hU5+HVWtBRE9LZD2WTOf4pZFwE4tQrbaCWLkqGoHnIfCD
wUWc3XHWCsDcxarBP+DjNlU9kIyI/cXRR5rrGjGIVizaQzOoYzSRln/bQ0SSgBgW
Tk9vxWBRMP5q6s9xoIgxetzql5LkVVyzvSPE6WVD/p0tuXyJjKo6Z01b3P6vlQR2
9Nhoqkltb9zHK9hgknnLQK0x6jAlTQOEGZa6WTu01EKofUUkiW1Y0yoTDO5Kq1n6
P2qIc3uXpT3JF9tzbCb0aLmlXqWbUAKZgW/i8TcKzDVctjX4j5eLGzUvjkpjqJO8
WsdLxccMKIsf4+BFjqiRn9Stl+tYFrqNO/nlDp6dvvSRq88B1G4algVo47bdl0l/
1SItcsHLc1iYzhwo0Q5ewhzh237udIa1PBTuPk7cu3U6po1cvg9ml6V4BUtR5MoC
gKiZjmd8TTlGzy8DM5WDYfiPomm2ZCRFhj/xB2wQKX8AqPWSeFcHXTquWk8OVOxI
bF+Md44rBPXBNYcd81lGGD/BTqAHdOZsVk+LBzjBrNI9dl793kWOXH8giBDzg814
geAd/k5dmxHxbyLtSzV5aLJrbJsMZUXjQrHz9IwIHNv1ORyAusfTTUJswOcHQxUH
IVyxV+/1a8jUvbiDaDnTavLGjfigmZZUtFHqA8cenOfMa8swANLDAFd+Ex2z0kyv
iRnxOCZihRkihlQBELJMhKtTkbpWAKRswa+Fjmxc9Aj1eHkpac5+jXbNLUKyPNQO
ydhsx8xbxHelGsFuQg7wE5DSlROEW/fkT21Xr7psSqpES7ul0mOzmVwj85qTo3B4
aWZ/X2Y73Ql04ezpNgKTFhrsASGMbHF+NU7TkM6EKmKAm86QS91FerZZwEZegpGs
lZ2z/5DhTn1TklJ/jkRg42EckyFKoULiBnnHTCekQG1cxfhb4okE8sfQAwxsxDgz
FfiZ5cJedzOFAqwB1s1IL8lLJ45l9oKB8Ue1SdQP8vGvNWgXaKYr3XrARUvhTrae
+ynwUrGCG+Uh3CYvbnWhFTJbUOXpOeMra+djYL9q+salfxtm+/QZRhoKM6ggnfZ9
HIf8aCTEdVoEAw6RmCdBQi7F67/W+t3wu11dsinG5pfD7sDltVsE5RGcGLMAbzR1
PIzUH/XoZ3o6is8qGPvkSdNrfoV3IMZnRjV7g1/hfiqJGEVx3MuLl2m2bdFhheuR
D9VasBzRK0279QRE2K3yucX4Qc6Fm5gp4Yknm/LDa2hQhutmoRm/h1zrHv6V6EfJ
qYcCJFOa6lF0JAL59WJcuTGJmT/1DzYR5+gVvDeD96CjBPybSdYEQseUh/fj6nrB
DwWOxr9D04c7lZgaGW0BqI0fUt5EZUbCXyBZHHy2UT3u5F3O6w0KRfApOMCJ9vTt
fpARZco+9BATsFEorF6O1bB1S6O927lo1ITYN1FICXg9v4+L9zTh61mCM2VAJxRc
QQ6Awif/P0gsQ9N7bWjXY5g8iYzQjzo2O4MUYESElQZdhJOVCYV0VpU9tj4N7Aq0
x1kR/Ws46GQnSWhXM88Yjw8U3TFjTDtUvF/h0tcmqIHhcyo2fg8GUTuf8sMJj6Le
v7YoQBrtwcQuGiaUyecMwPF+4dj3zjtRsOKgq4NvSCMMgnkZyzsop2FfKxXwaDzu
FjT/iNO7aldGBOo8O60BsysDHTJruF+X/0J2PTJYOK9FSS0lJ8JISZJzs0cRbU2/
NugrQnVCrbbDN5LdOf3gdiVZ/tnLnvWc9s7dj6XEZb23JD2gCwlVOWjzIYywSPEr
NOO7uRTV1pNioUZ7QEm9JLDH1U4eBF3qHXzHkUqGdho3DBvkR+3IctBahSwTEqD4
WQa37ArlLWIjZzuxO/+Kgdk/Bga6aL3z82VJYERlwYf45mjVAYIWCcgWRmBuLDhB
8ZiuVSryFCXdeD9KBdPAJu2JB5nG0Ht61peKAlUOWBt/QGdDnU2q6IV4J4aFPI1D
CqxVrS7aJkdArJ5W78VmMET2tdz9nxdM0Bkudw8XjCeOSlGr8BqZ5Lazp7C15phv
H5DSQX3LHsY46sei5VzCHGvySDtvfpRVZ8eKhPgZgfsmtFWMgRfcT7PIpQrqlkua
22eExCi2GFg/u27Qr3WGAjcbim+IC5aT6irEB/8LmYiGtzzOf9amqWl/kYgOK1qy
r/26FNrE+SbM6Lbv92zEcFlECqtxM7lg+dkeMS+kVcFyenNNR+qs1zuV2ygUeH1U
RcK5IN9e4SZzIih5utu6KQe727xXj2mdYt9DJTAETVDgw1uD3P03P37YtUNUZmA4
Xu0kW5Svffm7c0NeS1YJCLrsg8V2k4Tgt93mzcDUqMLZPxGla9doAzXzxApBPlFE
e44LuktKXnfWc/7DfvyHBv2WIRFhQXfPSCOIBT6wQLQEFFW+nOak4koZT/Wrnkng
Odo9KLOEIzCkCQ1iqBhbhtL2iI/UhyWoxDYEiOvfTnESVh6mRnLzbk0XzrxoDzuV
CzejrpWR+Kvx7LgYFLkoRDlRayV9pfWqdV5IIcNscGFDj2tqlUKNgZVxdlRSRR9X
TZ/YNwmzqxs9fARXq6EBAlCUjqrAxBAJ5qIneZrY5f8pf6YjVqxDcts+pn3R53SB
YusafFhJzj+clNsUqvPlj9jXgxdrjRLyx2UMrDepJ/WiF+f7zvMzGcbFXaEwaD7x
cOeswAWoyUQLekOxyBek+dSwCyVP7cnKAa3K4dGG0Vaz53F7lnBoEfMfByz7J1t4
V1CxpKC70OILIpMpM6bIdcTL/jh5WYTRPeOBtbyLvQ//+kca60ODp+fyVlOgWziF
FPLsqKJEDfVokOqCu19jJoOP8Ox4ouoTNPoe4cdjklLuee1BnHpqBfRQeeY0OUB2
Zc6IH/osYfWeps8rJ77BaY4Zh/lq0UMthkXLkWJ9TE0gp9bLBTJl/GImAYxNtkZO
tYbj8SOo4d1oVcEZdMeclRQb9UQDjKwMuSa9P83BwDJt4igtnnMo47blZyxfHeI8
KS5H444Ew+FUMWNKW+Adlhj9koBqlnv5TnTXaT/SG5hcVK7AJaPHokVp3QAFOYnN
uclS4MiLMWyyHorWlZ7xSatwuRJaPUlbYQORuPvjn6OVkkXJJaYWJDX8aFgUojj/
IuUIJdVlA3OzjhS4lFrvIkGiMWJizGyzLKvfGlaP2GS3LNEhCErW4MyS+IZ4Wm/B
0SWZeaE8Isg0SwJvNJoHAyTvmxIl0wS5vo3gqpGXBZCpmCPnHLdQ/lOvm2rMZf8V
fjtOrJaBC9va1AAwCxrW2DFtLcfs7TpprSJp/ZUesQ8MIAqM+/gDGgDdMn/GBUGA
oVrGBtMlDKgBqu2yzTf/Jr9zXPSBoQG8To1hmY2/pdGXKjhuXzOiTCGN1TKEJKJS
yjy9sM6vU1ASO8XxsEGrG9wzsgjhsO4cJ2gS9StTSgQ5dnr0hHKOi2uatHWRaJdy
TwsIw8vaZ2e2MTThObF9sGD8vHBu4sGUIBQEDfyElXnhC6oVwnGsE+QYuXhd+VIH
/XJvNvTi8o2DMdSO7J5jTA5J62eResxJvbnuOrt3KW8EUqmcmsuLWM9Jdfz1GXbm
u5r1k0Q+CfLjyrudNFnL88NXWOMZ9/5OLo6lIP6xHywyrBRCxzz99TkV6Vj63CW+
EO63pxA0LEI8D5Gqw7aMmoG66CO+8EhzX0paKbUvCmvAeEUkv9rtIalCHgyVk823
QS2OlIB9O6AOLXorVc/Jq1ziWre+hc9vj76wmhi1DDzdv7dN3MkGZh3dmlff1zcr
lKM7+414WBoqoxgEc2VSCNcfCCwvzW06qnRjDiTrTi+1/+lllYbUbUYvDG+fNe0W
mgdhONoZoCBfFdm7qiOha+DAJPQ6DUhDnEoKWKHSTkIhmMaQvuSJvX/UQVQYWItT
SaDS0+/ObYN6J/2ANcZ1Q7D9us4PLzi13c9rb5NeOlHWXx2IIzymhlrizoTCkQED
uVkmTFrDrm7y4FRoCGf7JJR2wrMzHcAU6uew8j0LifFhqAEX0KyeUojIt7kKGpOB
ytlrFwFaQa4zQVfMEAZWeTroUekmcJ11+zhvcp/7nj5GrX1AIQljrH7CWHIj6lU5
9+cx1Fk2VeYPom6QLX3g7iuQn7V6FZdtJslqEIwDHp16EPM35WkTJxZnWFjSta8H
B+xWqHr3bjulasobVicl49k7xqp0HLBH2e0JDtUgNoE7arUSS0FHxC6j+fW+xPv1
aXJF6vtfqgcO1JbILXlSW12+rULHOA63fNR6jMnIuIzzJk3A/4tRqhZELWrMf0xa
n99/ZBBcRapbKt8aYtT5tNjQ8LqxlJ3j5YMzBtAxMThhr7X4xFe/EHzlzKKGKK5o
t/Xe343JClP3y47cXUNHC6GVb570FvVHVaLiplNSFX8JyMLnFUjz5L9dBVb/Uhky
5UgvzK/DyZxyQf5tFh8HZoQH/eY/XBHftPtSOHH6YogK/L4+pF5by+zh+Lpyb2Yz
fA2w+6SK6H7jOnxNaiu0EuCsHy0BYjaQcizQ0TFQSNNJZQGzAY4W/mv6FVnaN6S4
fJn9DRYgZTCXOjm0G4CJl4sn8qsASXaXr8v70TiyGkKnpwwbRAXtiHI6ajtCdwnb
1JY6iqOrA5a4sTsiYV0O54igu8H4AA12xOPIXsmfPfDWZNXAnGo9/3sXQH9beqDb
vDeI0ZpPOI6vd0NbbWVV+lyu/chSD3dx2SqhoGdLnePRb661LEotcYRWIXzWJWX6
XwQpo9I19JxKk42KWWCmTQDtK0D3a0KFJSGFMXTsIJhezvqX13p7Hpew72UkWIOb
WfyOcZiN4cU3Q7I86P+uARQBFaRFQvbDfiDfXHT4sEUsdJ7AqmdBUiVXIbH1DzTQ
wmUkz5W+atsc07oV0bqLXZKz3+2Cp8Zq2A0YtJBB8e3DglEJnoB3kYvBsBM3y9lK
EOOi1/jQTccM9vPhSJDuRzKlRNF0x4xrXbhB9qx4JeiqCLjrxvMTL9SPuUjknP13
KzIEtJdogrO6IcDjghzc+gBaIlpTSVMgLBPtNX3uaV1IJ5keaMYReFxZy8sYwf0X
U9JbB/AuZk/vgOiqaii+aVFL/OEMOSkLk3UDeryeRQmbBLhymYv7e3YzobOGei7Y
M2+Uw6b+cWc+cmXsLSQCAlmltFNC3ZLqKhOQFKIIVrXOBl2iogorbNfCUnwJlLHJ
Y1U61Tp5j6NMdXq0k32+akj9RVlQzGj3ZulqXSycNxBTYCBZ/lTlf7m/UZhdGsHw
rLxqteyWEkbrncOnJT2/UgDOoCuhrymELkdhO8oLYDm/9ZKPCrpR/MJQrz8yQ1WL
bS1HqOW26fw+ntGcgfjxRw3I9ai/Vy3d1qXnbq0+zEaJmR7gP9DCxJN+IcJ9AgNK
kK1Vi878xDnoX2gXgvLZOxS9dmwDhw0AGAqqcA9Sr6uFz9My2c4d/JYNizzf6oZg
cHOqc0fDnyf8wecZ7Pjg1ODRAZBRLkY9tU0CxfD5Jeb/X10vYkg14Bv0IgzyK72L
R+anQbF1i2HzzHPQHQmW2TgTfHoAeIvriBGtFKghdmARjG28/ifoye3ADljCiL6D
RLWngKZDIUuA/qEFWPVB5jzKg+DypkhZloSn/w7lQWwI2QO0b+wLMjeRV5a+FoKb
kSQQgXWziER/OCKjn9WnAC7hyxSW7InB2U7MzoqRT0aCOR6N5eWCB3nG6vxB2LMF
+jJ0UHKdqoJRshfuOlInmCvsLNjNfDMe9Fvz3uoRNwCNPzJITGynA2QRr0eQ5xty
3BPqyhpHsI0GxqG0QOKS36yrTPefHGIoDD+1WJuD/Xc963Og1JEzr7efSrlbkN8m
WGYcxqce0Cp5bVdPDZCCVY8/Ig3JJMrM/MbOPssN+rrzBctvY/yfXeRNZrybVhXF
WO8dU1IhV58HIu173upTlaNg04uiNx/wEOn78ziZ+N+ou1F+doWAkHy6YlFPAz9G
EOxaVcaX3RtNH/0V2PFMuUOB3RcL2aZ7Z7KQGPrffV6Ju4o/lQHgVOp+gkHfr0gS
X0S3Ns7WIn4E6qSyaeLO6PdI+h2riMw+s8KTE5dAOztraNYVG5dX9K4bwoOWge5y
4aJLCko+pb4EPftY3672Za8tHJQQHdkqqmN7D8fn07iSlcbcY595nS3zICjoKi3n
z9eptSXf6B9TbyuJeWuIULEfHIOnvADkRAWkWTk9Fancw1ss4yLeSaEI78xvrA2v
bnTGgx0LOtcQP4b9CwnWzb77T64PxADq9tbINQGgPvv8+GlcKIuTqS9m16nuCQEH
lSUHM5JtRNYiKiW5BemL34ZeB9awFxJPPA6/V5//egJzqC0HbnsqeA5Jcz8jyPN3
6667LuadvE5D6N5ErJ4ESZY5S8htkll+5Fzm508a9Swjhy6R0RCKEEn8b9z+Uh17
tpwOrY7/VgZ3RGh/NbjwRysgejmV3F8uaMvC48qxgDkXjswOxdJxGUQ5rnEDGAEg
1OVI8y3s/pUUUniYjRAvgMkOLty2/5+Lp2lYzQJ1HcotdDnjoxOrXQaa+mBmkHfK
ZS66jWSb87oxhCF5I5i1TO3trRVi9dz80lJ9CKuoZK6KqirQ+NK62aBQIC7YoF80
8U72pdIBfsVXhrECNLFyp3Tk56y9Gjk0NFz4pJIZ3FAxI6bMeDVfpt40jK/sPsPR
CBlOGMjn6DEY7+IXhypZ+sQs7b5+MatO/nt/kg277VODA/KaVuT58kU+SveWiI++
VbhUYWO65f9Hz6/JFe6ySFsz103cWvGXT5wPR59qVUgTyzggeAt6PxzxJgRVgIFk
emAdKTgWcahunHrd945aykWQnklHxd1v+pqL4Bt6UmtU5+nG+urauvmpDwNEm9J3
4FYMx5OlQI3w2syq2IEx1aEr1ibrL6n1HTCl3z802kuSwrhRrbedUZm8YseukYDc
PG9oBptFYJrVNyfGb+GPDNFBwtSxX2+8EkJWY3ExYCzGYjcqnxiUYHqb67MKmbGo
qXQ4IqIVZbdWqMyiEwf+QbkasIGUr7DFi/oPG13RbsEHB8zokbRQhM1BnWZTYwYt
DyDFyA44Qx/e9Tn7TK9GJHNdwQ8i1VUUlK2d2NdkcQJFgJ9LY75Qtw497ccROtyz
q4Ena5k7hUZAVwOm2VTpg9mW1Hamdwbdf8+IpvnmpfyYfnDpG/mjGb0imA3O7ebr
69ALsLL6M2N4NrXnev+dgkHtyxIwDKZrT7AIiVo18DFOHijGN59k8kI6knVGuNqx
4qMRdlgWpE2jxycKmUeYuIH6n2uCuI6FhTNyZpZdlsjl4ITG6naBLZJHpIgP6JHa
TAZM0y10DSmc4XqvRwysbzE/eb8Q97V6Ifw5KQmzqKXeGZA7iY3nCSWDqQCRrNH/
bjup/OUIPP2vAVwH97kM8DqFZB7d8xTY7MvD+Fy263MrA18IEBThnOm8QylzxDpG
6MIZbrWPyVlUpUnWECpGjTdzyeBBUVNVpJ90PlaannfElGiI8EcW3OyJk0x8XYen
EohFb+H9BF7TECpqUdWY6Lx1ID1VXXlW9ZQnU4+LtubgR9X4v36pAhCTCJ/OjC4q
/GxiOH4Y1FOrNuqY4ahDRkg7YdMquCWG3Sze3/Btdb3ihZE/dsKTeCPNByaaFX9b
JWav4mb/ucgIPbm4bf9wx9EfvVP6m9HBS8+1UolmMh2LGI76MPqaf81aDxv346ln
RVJDNuor0uCmRHHaHAUnWz3Xc5Gg6+ZRvEkbEhLB3AhhIaui1S7LZX0fDnQz9BdD
es3VkfKNfoTC+DIeeqQUGWaLGdWVW0JGsBy3+jLI0/dmKdc1sHVUAyuQOSTQyVh2
Wa5r4CK+ekv/AIYWB+lYGLV8yYaMlwgyGGIKPDoROe/gqnHeEcg3Z9faGpiszjXv
ZONsq0AJmMFSQcKVgfRGQwgov/cyjSuMJ00s93/7aVjRyjHktYlgRp+Hc5jQzcZj
+L2dr9QkcOAG+2EQvY/ej6FAcM98R/+GunbetU5iaRIDeESoMry4A3wYCMRgmv4I
GS8vdyQn27X8dx/SR4DNaaOvAletY/2til+sT356HBazXuyEr7XXhtxxW13akXea
7zK7fgQweDYuh9HwjF/9ubbEYfk3ePPM4gjwbVQqCMM/l/3LKux3NCJ244COlBxl
Zp3o/J8pMiFilCcsPHpu8QIjFIncO0XI7YUt0at6o5s3wZr1JdCC8BaJKLhv6wIM
MbvMfoDwXcYO4yfEZuJCS4LTFRIlO75sFudeWsN+jsXvVFK2YiYFIXbSCvdo0ea+
eQ0ZQHRlhcfMZokho8OzqbaNJkINT6uKqZlapG6EPbeLbyfypg0ELee+fqmYmogz
91WTup128JzYZRYjW4+V/Q0aa37WMQ1j63PM/7+j96BHnOcWMQLVourz6fU9sRrW
/NqkfvmzXdLxW7Dxh3sZorI07HPjRNjJBJDlbogN3uzUjSUrbDHBDeuMygHJ2PRX
AgoK6aPxU66vB90IvcJlDsTI/tnXTX5CzB859cJgJ4v9daLFJdoQmIbUVx4K/9/I
CDmpUOwfx+eTdddbnorbRwyL6QxfepCG4Uvc+MDH0UjhDUgF2NAUfjUBNfO48PB7
kLqu0/PuWTq/0Irv+lfLbyw58pNnig94L5ZWFEaJabijBhmfp2T3xaMlutrLrAgq
ZD72X20UHpEmsL71nP7QbchSDUQaar1VG1hGbAjgrq0D4EMvBNeFcFM5yQgwY9BW
IzRcUl2fxjzVO7zkBcm76+rPVNVmqICxKqzqJwGopgmBnQq0eJ6bdQ0Gt4EVZIm0
JZgGauuy608SMDwBNXST0p7zaGTunfyqrXZWUjQlcnC62LfT7b0xFuykCCB/ifEY
tsbGGVzekQa9GK53TWylpCpDEaEVVoMT64Zw8yJESx7ph3JvXoov3zfeK9/Oj7OR
Cnka57O6dNXr7mPALziJa4RHNAxMpJNGI3Jpv2lPEfBBSV/WfrxYjEpQHIJ4HoTs
7VJMV02ffoz2SJY3VXVViU2bP+Du791yoQiOikVupy3UG5hpCtYqbRQbD7pdhWtY
My9j1g4YZsN22W1dTr1T4BCaw835dzUV07LW0Y6HEtCJmYC1nCh69T7CQnMkYBRC
c5df8DJNRYykGozzpJ7jDi7wn5fkuK36Tk5Mq8KW639SO0C4rfHs4n+SeZDLG8+C
mWSoLQPDmW2Orv83leDmL7pOOCrpjnbbkB4rLQVDUeMtq5yK37HjuqREtjjiVexY
7K3EDoKRUfu0dhQkC2OMYbiV4AGaz7hw6PbFScVwkmcoqy7zmi/NuiyxT3t9Qmzr
OkadZNE+WSkmDM/BsjSRSE6xrRBiG1vUrBkiKlnAFB1tQ/4CUgI5soA4wPd8MzU+
iAUkas36pJjx5kKA+dNzYnWn/spbPTDz2lypXkUuPv2G1OuKCXH9Fo7S8t06hDfQ
6zsFT53vjMOiGdUSoq0H2qk2i2ORwblOdRtCLBH6QOG5ww3sspkWwAwMYUdT71Ue
jFfKcJ3flHrO1epHmStuTznrIh16rrEbjpu5dhNF4ccZOKmdTua9UvZ3EN8ZRi5c
ZYO1MdqwHqlrvgNpAoQ0Y2c8H4aurFaUTW9Siv2euNX/KMDmZ05SsDdVq7cbjeoU
bLYFNS8JwrUyWMwuzaJVZmSrtGTKWYmo2Xp+d4uAuB+iWsfzkl6ic/7NT5OSa3xz
trp5ZX5a3QBOxObjhIeQWm2lVq1Nrsk1catBx4ri0wLAdw8rYcOAmZ3v/ghWC3Be
ipd2Rq2wVgFxDPpgmfr45qVYpaI5ope1drjOSb/zSA+3bJGK3Hkjk36JQ9DMAsYg
R/XuIkbkOD86qKUisHhCva7SIKSbkntIcXFkv9OYqg4j5iD8c/dNKSnlLAid/REy
BBAFuM+wyTjzENloKyRW5hfQxadtYPSvLxV2hXgdrermERyP35EeShv7dwge/uHU
+j1FPT4UiWZV/x6V6B+8J556r+8G9ATIdn1NijFxHScwXuMwhXsHWH6k3lj7+rh/
5JL157vnZpnaIoJQm0Vs1gmigZTgOGXvDLwx8w5Z9kX5FyMP72BTaGB7Gw3iKjDP
pVWOecdivSUoSEkvyvdci2RDBB9nx95iW+r8a63piBoR/wHY5uRftAGrNT6pUhbD
JMRSALnBaF+Y3ngOc+BJ8eOrOKGjT/J6bbAVKHoHYq9GkuKT7rVpYlujsxqS0/8l
3VuvY+U7m4ghGNzK07NrDs+F5WA+EYy16ggx+o/B3jMBSCmp2msNeag9HICso2B5
OuLr1Y0E9C6fY92L6bkq/dJG5lHIYPqpFPtbCQtndjDmyX2ggIa/akZpfGGhqkDd
z28k9nb/tCB555nZu4CXYRej3DNnp1ewNUXPvp6kFHtjknTnFnHhDyq76LaCaOSc
Kbzuk3MAlA10/W1NefYNRz2sox7t1qIf7Ja3zHaAMex6gQjl1DGjUqFvUuoiPL9Z
dHaogcyCS4J1yKtM5j49nZdDuwCBF4USslgIpR0FHyEeDEEWUJrxJXhLhEh+Zom9
QoRWToz4f4R4lELXm3S9i2jhHdtlSSWCVBmm9dnLKk+2DdJlbB20WHP73T722hUb
NYAGBNth9m1exVVL5I0jUw/QaRSzYEm6VdfNXWX8OT4wcowMz8pWN3LQyEN5tOb2
fC71+LP2fBdh8QiVav8R3Q5k1HMzHFvMFtb4f3dV1dZs0lBe5koi/DJdRY2AQFlk
mnP1RlLYa7hJ2tBcwWI8WI5pEt+Mc2dvwnz/kZF9v5OeGPKBEJt4+mUznalzf+po
ByB9b420b9QBrWT9nvyX7SYEk/wrH/BFiWQaK2rBm9mEHiFAx22ZvFboDU9Lpg6l
iV1mJoo/guSgkxtWg9/ZVDgPZmF4xp4qQPAQ3C204ijNfXM4d7Yp44bkLIWboTT2
506Z8GCjrt9YDGoKNmUpzDJhpesgEF9EG2Ee4Jr1GX5XcLFPaS59DXXvy2HkYuQd
svk6zpkO03fx7PTnekHs5OCo9pO018A7bt/jLgG/4WBXMsbjaj4Ft5fWVRxczyqR
DWd0RkvUuOLHjwBJ0giIyWAQwxKPybd+J1iDjfsD/j8CBUQVvaIixRNeHLuRYVZ3
voHZ93Z9rSmXH5giD+RwXdkwf0Wlh60wPDU/c+dEW8tST7qRpmWvpqHxPj6Q2n/E
feWqbXdbC08WtnUft2g4NK6qPTwIHMRYZ086HjPDlaV6F0dtV7RIy3I26pOs+Vgo
TmRUM/pLos9m3g7tvbF4md2rWtutdxEzH9cCnO4cPkVkYEaAB2Hxj0QpAo1VQL51
E5zT+M4Z19B6OEAQv7vk4A/b9GUg+pUQdpzx1qPdMM2o7ImmpW7f5vc2Vfao9Zsd
30a1acdhO8B4sh3AHA9Nkxgkvn4KH8TAXl/N4EdkhXTHkg6mYGgDcv989L6oHh2a
pO+lChQJHhqbK/faoMvNS5DMZHus0BMiqS9480AqrRF59ENNANN7JJk/Y6rruiNY
pompQbgaKBZXrbTOCCWilNxwzZlik8FMHlKSBOlgzgqsXhGNHu4cAkjcCddjvuPf
LQo1/yls6cqyXx4P/JBVuIj0hOnKnZX/ggv29VfeWtbOTm0K3W0yMalVo0pu0SpN
jq2fZcbH5a3ng81dOGlwxPba02ZRCCmTzIhYHCgqHwD+kHIRxPMBqG86dGWazKBg
3m9iiZNIbbMjzvE+pfX/QM4tjcGHQDIj2SV0DgKPWUwIIT+3AXgnSjJjcx2olSDK
jdSGbP1CfEkO78V5AtHvjHYoqHVAfXuXHR7GhS21cQVF0oB7bhDIKhRcnS9mCKmz
BXLNUEDZtXhT7NMwG0pZ5kapL9AUSq9tdP4v/YehyAtTqxb0e59ETuYWq6XjZafY
F7+FX4zR0HhtSzZGIoE5k74nHu0avecKdJcde0OTMXf9OuH4JmVmLO8rlzhGUq9v
NF9BVT9DJ+0VzQeGdYG4F9PzN7K3HTls/J8VsfD5rUbF+jCOyesWkFY7YQCXWtVx
wC437XvPfxgQfY+1TG0mpanLE6Qm2WWZj8/Qr5xmlza3U21u/qGfMitnR6mSF7Pg
Az8gaTRqVM3ibW5cKqD+fYOa3HpNR5bl0m3NMsUTR7n5YBNw2yFZJe6MibJh9LP3
BdksshVxJxkDxk13eS0UAPmOAW2lh4ZC+O8IcztJwuFMOrIgWDcfkg8y449vSCKN
0aLwpFmmM38O0yxIg48wW3OZKokBriBoaBE54cH2Y1y/7Akj3PTTVkySjQh5dM94
ABd3S1OYw78oTlJoRYdurQixiYMWt+n28SNuuVmVZ5GKjDQv0pYnJSVJ0+TB2mar
mtdHKAXqr/3iUyHchncAqT0/vglg1LB9M296vAKV6nhrnVIIDgfoTV8boZqIeerY
qQpQ31G6drau5rF8Qu2K2S2tS97Am3DrmV+X5OVmPT/4V8DKi6J+GlQylduJW9eB
GwLmGrH4/LGdpJw9V49qvUkrmLMtP6rwXSeSMogKKV+noO/6aG7yUGVWi08zh+BS
OSmhHxXyNGuwuy3tYprI/ktdyIMWbOSMjjCyvXzdXsKl6z/1lREy2so7nBwFG3qo
A5HfqX9hnZGf1Ogx+s9oPWWJMiMmB6ucnQ9EJZWz2T2oZA2AyxhT/cuciKL5gFYs
NugzYFXmg2nz1VWiRgGe+sqHiEdc4w1F6KJDWsDGYk6N8QB23w470zIh4Vo5xW9m
6Ff0D40eaxTbRn2k3nZvK5Q7vE4tQX4CQ0PJfIZldnoonZDmE3RRVULnogQMfIKk
CUpGC4KE6ZDTcBIxqRSwft1WFnszpDg71fVcC+811uHmaKwJRUuKRHdoTK/bbMiP
SsxPPGXUyMlKgCv+DG8BzvdAwkcMzQntYMi0+BLr5wL93OF1IaW90Lcq5yxRNvnB
p/CSlmTMFhG5cdm/2LiT5e81jhnqQkUullINd4XPm2NihDaemFjOYGsPW4hlSpFK
lccmcTr17d/J2qnKGB2I4qZpmalN3KaRNYox5JplisWysOTRJmIFHqS5QuOA+8PZ
7wfnpwEztJ4QZWZOz5NiAUROx7VZ7yAjNDCvdOUXn77fhInDKNulMyywRt9zFK/w
f9CbZzG57NVpk7cEiOzlSbC8gKTXbivsuhWUvtnt6ypxvQZ8RA07saKjInwky9Ki
umx/IlAqM089bJ1GRXxqRwh841q5VaJ9cDwdLl/zwIXT4BWzoMo6Y+P7/1TZuPyq
TF4qvUvYNcCklL9G9rp/H37q2pQ00V9FhVE+8smrsVdbbYrMLj38YNrXsPPKEGbl
FADHtyDZAD0tGIQQNJXpMvGjg0zmP3hCqmEpSaN1RGZ9aVam/HVDVlcouhL9yQbW
85JCIS68afscQ8V3pER7MEt1ACBdTF4CrhJqLaPf6mek9GU7eQH9yazgkCHnG+FO
xO3gMnqtD9ggMG3IJZXeg9lTl9NPizD575WUvMkR+CE5UcHSTi+cT7A9rOOlhoh7
eWenO7nwPa6GL7bRy5oy7XrW8iOEmPcaNVfSACkrBwzaa1FogqxN/rtHaGR2SH2X
OE24OChF/6AgP7uQqEfYbeEIkecwG4mBm7q8uD68g8cw/aD+OWOw/gxytwUykUeO
zG0hABaQYU09w5BAFAAe1Cm2q9caxS8z20cF/hwI1+2SP0327xiLMTCufJXRRaF6
eKc95ICeivtOKlX/x+UpB2iCWv7xJO6FD8cMeCaYyWzFEfddEch6/CPCgyReeO2/
Hft4ZFIMYf7lXZntzdFe0oX6wj7M+0MeEaxWsLvs57P5Eo05JBcV7zwDBKHoHQX9
wsYYxvhgKLgBQKMaR34rpPd2JkNA80h0/GiULWtffyDC78SBeq6KOqAzn4cPl6o1
MzyNvYQNrYvZI0Ty3bC0XpzvWhUuOsuyIbPSE7bhtsHOucrXOy09CKE8TeLKM4/W
5SZCjjJTPzIThbZVHBa3ym061qU/FHWR1SbJFRV0CyCELwJMgEJI8lqOwnyRz/t2
3+hB9javXo9n34XiTZRKwpu7oCyFOeyTmhqPG1a7K/9ZeFTrc+Y/53T22R0XveSk
8Id6OGFGi/l2HMu/FVXalF76Q+/dK3jtDbZnaBQL9RwxDI36iEj5DG5mYTuS6fVn
wT2TDTfT9edZtTTjBzXXPDSzI34hgik+mTN/RV625yxPlf78//l8f0aMZc6miu4X
+vTrmUa+FpkAX1CONdn4a44/81/p/gWeHU5i927UXEPotgzt5mmeZz+vk/CuCGu6
u7udPTdMY03mRvIDyHuyCa5fmfKi/RhXkznTxZHApGY0VDfTXJN2V0pldip9XySr
x8uOgx4jWx1osL6xq3ze6Hi0OVlAxxrjxffvPGF8jnQRybKsbo2XkfOKt02il/YT
/sc0Mh18qS9lePu11NxfWBaYATOssDr4MXcq2SyUTJ/m9+JZ3LKPfNFaWWZpgG+X
wM/1Vr+/46DX4s3PeaxMzeu+MvTHMBFzvFF5Qe7ZnwsWNeDvi81dRqqRcTnkRqW5
eGLTkL1iY5+dF8ylh80ugJEq3tZtpiU4F18fF8gA6Yvz3StUw8i0Zhx49b7NhWc9
f9ga3IzLR2pj6oteXK7Zlgb0ZThpk0QUbxK2o7raREIG54r9Ng8Rb0FwBGlzf6Nt
XNRfiVN4blDXxgVIwzG4lMXGZkdHlpFM59hnEHzQozUWvFtdtWuEYNjlMYl00XKJ
JRm0AZkZSSOEHolsCw8NdRmXFp5RQbwZelo5K9bGo7Gh1zrq4FpIEoTRm3T+kWXg
8iHNIGD6Ai5p3ElPEzOt6ME71qCDLIp5k9GM8ifpIVPuQN5yx7j66cE8XEDTweqT
pAmwZBGVeRqeFOxO53tC/MhvgcJf15vKD/nPL+kd8enjfGawcChyMDcmi7efNpn8
v2eyE5+zdV5aVCVxuDHZ88PO05cMxghVlZLdKDYoraODqDmH112oqg/jNIQs3V9c
dAenYSDcWVb3QpHscQKCGXeQfyxBVI6q7Pkwzcq/HqGDT9rCzfW5Rr7v+iclkGgQ
TyDeHnreWwR1pWTaGPM+Jv9aN3FijUo/8JmNHVDaYZHErUMVwWSHWjKyiFzwDgE/
Bjl69OWLoG0xNFH4LqxKdSuSZBuT/CDWeAzrB5T6qsHN4TgUOAKgzkIKOol2X8Ql
jv9iepbcMTS/xzijXp4M7eSGoPVahqQtUXIoCB+/5u3VUkeaJD/LHkoZy+96q+3P
6rlxgGBEZM+O7SKMl97m8zPtduETuSw82k1u4m8ZB+bA8z03slkA53sT/0sGDuXD
wIt5f+XjFJpj8TbA5y1vcBYko1/4CY+uTXNEXXf3w7Hwkafeun++NxQ/aF5vW4N+
/WxjsVqjlKFJ/iDKmO06JTn9Qqe+QQPs85E9UPlIpLPAbJJfoBa4P1gvUf7RbM/8
FWRuWzm62iLIawizprGg/20m+Cwt7UHbMYbfhHGchuQ4U8RAG/q7JtY//OKZSrJ9
31q7OSVYSCSveEJNs1OSgtvjEoGiU3ZZ8Ucf0ZUGrM8pr6Qd42x1rfAVmPUB5pg0
OVH3meH+Nz42iFbm3IYSuRjIMhFBwcL7qHvQSbnB6CYKEDoPP8uY1Ldlj07MLyLD
7J3rNUqAam4PIHCo9gDY3bOQorj+agQ4V3J/xPNCfAmJyS0Lb5oJTp/IJNA6JjjH
+YnGQnY0/Hw6MQNyYcjgbjh5u2S7KWWJ+XZH92SyaC0N6RD++XvxCj3et8LsJL5B
uNXuFguoNjrhFnKE+gBNQUZds2FGyMsbuRtLpVLIldYbW6ZVGKgBxuc6yQh9iAtt
l8mDZ3rzjd2J5+SZJ5p8Ci/I4vyLKHIdkRWxCVYwcSEcUJB5Yn/VxNs1eaqSdiO8
kXpHcsZWGVyp7U828Ip1VaqXerxeSpwnwRoxlpjfcJuJtixsWQLpBC2L5Oy9FgLP
joI2FdDM+aC+IJfuW50EgWXQagNXM9tJCX6RmXYSpnItyz9+KA8GyLdnL4TaneMK
RWFhQslTgNUJlZ1PIJqqtKVteSCc3JWbw2oJt1OnwhhgF8cmLEojZUY0EcTVHt2e
OTt6jVzdc0/CpgooR1G3b8xV7ocHxwSAjFR5nVLfhtc2gAbrbmj30lTwoBZA7Rea
O9kl3z7RMgzvjpCoRzTd6Chmpw74MQ7Cb6QI95noTFdlW1uPINvMyOKtTkc4/aBH
FPRS8JAjNdk1ehJhwMK0JAQUTQfgnT/yVoNh/DUpACgoManYMER1oMktxyGykHJ/
rd1K0zbhbQ4aR/ly9pYTAHp/7RXVlef6pPINQ5P0qAWZvYNgZSREOMQOEaW8AdS4
6wAanB6CGfa8W0IaeyxlbU1sTjx0uP6XrhzTsuHi4Un/bxzuh6xO+vkXYlYJuHES
bNxkTu0UfQFZzWQjCliz+NWgtQ44wQCOLpOGinLTUsOleiRqKjNJZo6++npPbvKi
2Cj1TjKzQ9puao503TDMYy/25CcmutVcI9H+Y1irUUGarZ7VssC7YSUFOFNtimu5
FZgOoRFc6s8JLX9OtdaopLxC5B8OZCriJRNHFNSNS0NP9wHdE5RJEyFyRKoPZMuW
dWnKHwMTehhG9iA1q6RdCTE82uWAHUcyATfL793bdGxqrwJ8e7h2i/zgJn96xMcM
9XlleqUE3bYDDTb7Kib8jHU1Qup8Hho8wbfkia5QVW8PHwJkql04G+zMFUq2Y3ug
s485vgknZlK6stfzFuvtPJ/ek4FESdEfJpE7gDUIYdguT3iYKCQVQlh8KVXyRXYQ
o5jrfBVd9P1B6kBA2LYj5lwFdsFaALuxNSJKy6RGmFqjSfzg/2CBehLKntA0kBnX
B6jcKhLzwfBTd9gJ+DAR7557bezb9GDSgJ9WPr+sMLpMcAMrPX16vRWumUoszFKV
xRR2n4cvEEptplHe+Q9tNg+0e7ffdPclARUU1mYTcNNifzt2NtczmM2Tmp9gIGAv
SOa4WH9cqT+A0ODmKc0OYmdmAWty3vEFwm6QwnyjJgsY8L57eo49248iYe7AVJlf
GYq5YXZpVwFaNqm9oq3yA99llABqBZXv7HjZU6dGUOk+QDKOlZThOzkICIaeWvT0
sloZCQLWBSAA3gHa5MSxM96Qd7HiaeYRoIlYRy8t8g+HnLpeUfRnq3POf9Q6OA0i
w5meNXL5NAms+Y2s5GR2prAMViavOn3tfKbeyoJufihDiSFhLwf447fuq+lsIyHP
LP1WEtPf0GYN7PtEcjx8R1bP1tO194mCWXZrZZGWjidNByFv64oH9AofjSHxjRMy
DaHVRaGOmFPi1t47oy0833dZhvC6DBu0gyaAaZFpU3+AvPUkm3dtcVUL2an+H+vh
KWF6MIn2o8pIkdjJjCJuqkgl3OJy30BnpBWkH82JTh22/tZrsiQ2OKAifumyYuHo
Fs5WJWG5695KcLfoKZbVXzgU8FQBqkvp+3W2NlYsUmsQFf08iLqp/Vz26VvQcgjs
3AeF4BYjT7yZwtreSxucZALBGfaJMIJ5/nEbaI8f883/ddCan6xDajBj3PP9uXvC
2nSDp/24m9ILpH9QyTDRRoFPc4fpL7H0YfUgPhVhzoG5k/8PiDlhSGiGeJ2eaRNA
PDCftDUe57WBVFc8PnoH7YRt1v6JWoRPr2BRE6sgwzy8PFsAxdxekxxyfuvUirmJ
+rebYGZ1mBl7eCSVr9I/Hsc1rbDW8FNezNkMWn6BuMXEC6OCCBXZdIk00/rCa6qZ
VHJWAVlvdRWe8rla/0G8MKbKVqO16jb67ZW5HgZPlgJ/AJAh5l9HIOinQv/exCZ1
yeFy50C6Xg9K3FmbkQaFs9x5IDXgwkqn4RB18u+G6bTl9EMa9nfTA1sFJYt4O9Aq
muNFPAJw5m7MOtfcfoUcTW1d94qWltXo6StRVEotFRRKalVf6s4sUuibSWOh16cP
TY9xXy9rYRs7U6PxvAu/m/8dXEunOQBVAGUSVOZlJ3pAki1nbwTUNBQRJvEpRikr
+6lwVhKffOcdeAyu4mqQdhU/8oIsxMZ7d3Ao1zSv4Iqd1OsWjnXjJ0zjMjlwe1Y2
MudXYEesiOtpPZh9p6Xdp1FR8zb+dOechwSWFZEzDrZs45kHZHpMVNywUYniwl3n
6FmRgbkIRgSgy7gMdRB5n9OTygl3rQvtT9AfoLIIExXP/xW+VWrd224C0v3WwLzQ
YaCDuQC9U5Fsq1e/SwbJ7CsE5Oici4AP7+U06wywNC96j4ECnPsI+0tN6Y3D0nfn
MQsytRV6nMsfibNve7gcyy54xMTR5RRLyAl13oaVrrSqlz1YXX67hbmonysIdolr
5OKdjSsNxv8GeHmU4TZhdglQVbpTysjj8oPN97gd8HQkedKMFcMG16i5TaHvo3fx
B7dzOLX6z+aknNYFJWSo/vIawhDLMZQYsWhchqBzOQmPESR0C3HariYk6DrL8nCL
oWENjN5PnJDg/9kdxZkQeTD9EPC0iFRbjSX5MJzp7xy7HL4VMfQvT2by6CQ6QSp+
G8yKkABdrCHH4WGmpU3METCwBkautrXVZ8NJmfSYFQYfsnBRq4Z/CN+f8kV4Bo8/
LClMP8z09NglURMnLY2nUErob18yOfE3HeDuM0JyEdnl/E9GiMBGRkson+PXwufs
a+pChRM7Ba7L6gBvQWdQY/SEYA99OH5WInGo7QCWi8SxX0fqiMOFoXz/jlfjNAbP
Y+I7x+hBvbxOepuoNafrC/HNNoRx82tsP09DY7Jm3fSNEZnCJWvOop1BpZB7zDfS
JYLG/TGVwx9PxzoXawG093t3fZGIq0SNfKLey/0yYqVJdZEUOXV1A6zCyjt5nntd
B6X1K6g1pandYhoiykoxx1bI6KJsV7kr7bs4Ri6OOGZwHVpAcw2ij9mEeSO4+zDl
RUE/f8l6tYrSxIggk2bXPlm08x6hhu2HHxSH8QUvhz2mJPhIdXRZHcThIlBBk5Qe
kSu1Ucepz48qgbp7bUMjvrsHBCvSUlPvCvc86QiqSKXljBsV2NkuE3WoTnq7WgJg
xmHoJezE3OSuUOiyuZ4ys3FCfUyFLS5Ean0+Lo0XBbeubNYw3O+4uFVHvK4XHumY
itbnU1R6yhwr8FwD7oAqeHlWXwxLnYKoxxsP/8BRaiDANrOytXrTWx/YKXGZ6ZA2
r6VWCUcdAcEc6hTJcIkYhb5OslbQjwFomcWwS8t9w2+tgR9L6EzQAlAhRV0saqep
RPpzdZmDzQ7S/NedIJAFCUEoByBXlP7HSkZcqk3+5QJqyMZVHwESfl25Bppqqedd
R/vS4fbwsw7hTx0kdiTBQHJH4cKCL74YA6zRnmR4/yx2XJbMqgMdtT1fqgRBSh0R
ykLydBa6WFD/fH0fNK0sarH/9+OWpBU/pip76oueVvJDn7gQ+8iVGvMNnZbK5OPz
LP3CUHHZZ8xBNU79dSmIfn+RrbfI0zrByB/TuY2XUrHKI8PZkgMohHhzNyjNIWp4
dQfKIIJVBzxGo2b9Vn0q+zAUVOfYOsr9rQQZctaXa10iyECUOK3ZZEu8mrtx2l9K
kJXgG1hk8k9aTuolJtX2pgeIrn8Xs22WWaub4UNj1hX1FO3ml3mB95k1NMzDFn0N
JuAujXQS3ONwFb05n0VoBW9ee57+pOlAD8w8hf37i1paDbm/jWY37FF799drLbGT
0fwtDXaRJbuypKBhTHh0zXMvdrT1YczHa8Vos9+brXh+buRpf2gcWk6VlZAHfDzi
LJIWlfvL5G3BXQAEhXsVwLdLtydPxxq8CnckY3uj5hGUyAglFkUn5rXypvpKTzvJ
wJp/2q22D4BfnK1Usy+8cq08s9bVy++Sh34DWReeq3M2/a+eoilhLAJaWa5PQn6B
DCA3adkMdk0ayWky1rpyPqJxgH+B//u0WymHbSS/8sCPzT0TkHdkkTzVdLLxuNIz
B1iX0ccfA/rOaGCtSqvTiRwfr7T86XJgP2RsZFqNFgau7gLLp1aWa12vOi2dblSt
ruPcVud36bAFZK/z1nEiir+d20NVLlW2AmRUxtH1vvJU7vuEmTDssFuZ7s6hGWCM
cunkZ2B+fw/dvegtp8KX4mrXzzlYmLwh0xQ7I+PMsAU7K/vnm9bD5r5xSjC9hllI
z4GBgo2Heis+XWMmiLacPjn2kI4j4fYbEWPp8T9i9tIMA6kFxH3fPYkSGwzeETgk
2EcNOr3ud0V/pkt94n0rUx8OHub6Nh8xAXxSwU2vZQq+LqPkwMoBvXF6zAdZkTor
Ixyln6oGz6FQ7Aza4ev21ZAQPG+9Ukco41+Pe2GdUfkBPT8pfHhHJFjyDDbIUKyR
MlMWc+FiqGVq5PlUOxj0p6QXNDic6DUmHcjgmC+F7+idxa1vb3ABwISx5BoaRfQt
5/3Ku4on1R4NlINUbG0WE8JBIYpz8XZmkFm9Y2BQN5wy3pATBm2nGPSaZINgN54C
445a7NgMgGPmBcZAlaxHyP7gt5z1L9p3tcpxcf6nKpUVM16kaOiwm+wUfZezSZzs
eQt31GDNZSF6mPwTNDvfgjwVirZmNW1j9HxoPe4yhyYKFkpTLC0ND2yJvilcm04i
EzA2PKwIWsnrrV3pS/OkkQ3O+fXPxZ+x8Go0f93X0EP6GfMJJiODQU2+rRHKn/qf
QgkmW8HG1rTM2GwhuELxU7HufOUTJcED32uGs3GCWI7PjodcRER7urrnUC7s7wrq
I4RCRlLgPy/B620KyYrreAXXrvfUDyZLasYw6o2Aoi6T/6hKoncWB5idIDlVU0+F
LyXsWkUK0UGH+wiQI8d22VroptyFqrq3azdHjv6U5yVYi80YTLrFhTvQ4vJQjILV
JttFscZ128Ktjvj78ADp8lmBZaW2W0g7ZdpKvrocuzkjCv13USsd0dazlwY4u8x8
FFb+K1yMhVZ6RVZ/t36pGFMOZNVwxeTzLVFNcSeMTMD3edDWe03qqPZZYYS85d3W
TgpVhkH2ivQm95ndxlCHsxpcBukhr0GmAwPXGLObMH6G5qfH+prIuZ76ANMHaxj0
LnTGwZ1BiG6gAfZkDk7Of46sqMNJ0xPnyCyn8q41TqhtleJXZKJWa7HwGfUe0uuW
+dc5H/6HOmLYXCZg66WxH6tPWSw/oXlBPSRb1RMgp9z94XHIY8CPiuc0usorKiin
O4YEVODKXVDLj/PsVvbEw/CHIvV+APmP2EwhrcJ8izlIHBNsfET9Ks+kWf6PrL6U
HMCntOyZEX7HsIjvG08o6AZ3odYskYvDVgFcpN9iYFFx9xh74bEfNBzuz3apGcCZ
jwnNJi43s11UtBa5iH4t8g1SB9ApiFA9jU/DvVjpKBFSnTkdaEAwMYpX2VBFGc1F
GfxEbVv1cYuJm0MGZrJXa1+lRiHOrFf97rllQLGWnXpBhlb6sb+gFXsVoxitmDxT
QuHo6MImF7xCVxEHvGRkiTW+B6D+NPfLc3HYe1PhJQBI28vvG8WuK7U8Uk4AD7mJ
UUKcmTvNZ40eeqQl0SQGQ3O1mYaSyoqJyTs1sjs/IScB2A8ftnU93GsLPc/mR2BQ
X0ccX/TEg35/QS1O5FG8kGtQZ2umxsDsY4t7D2RwmJqD6EJPvLO3w/qW274nn2ht
PbaUTvvBvWcyNi1nm51AdPvRud83009h9ZUs9wmXpGbIov+01Bk7pbWq2A6ap8RW
6lAp6T2v7j/GzBS9MFVdyZgS88U3l3jjVONcSvSbu5RI1q2cfUHfqi0OJEjhls1D
FcGS0/6C+wmlnGP6BCRQtnzWSH2wt6VzCVV2y+RmQUELKp/lWe1Pv7HDwrjzpSox
VRK3ci33eMDL/ncrAd4TZU6ejGl189g4WFXnvfcPhHX8Fv7bbXK64dFeeZsuoTd8
RHAHtEMQ3xXdfdxeg3Kdhr1OUOoNrFByYfj8MmyQiO7NGA1MDMbWJT06LwLobupe
7B6qcoLDoabzPwF3Y2NA80UX3CMUKaO3um9Q3QxdEeTzk6m1jvhfAK57fvzpG9X0
8PV0pt4wOL81C5pHiImUZm1oaNcXHuevyy+0WIHbemp6dINFeXom00P1d9nFb7PA
LEcQ/LjD7h48rcbBOWIdv7VGCpDl1UorXirTbQkn5FSTSwEED/eDrTd5N+6Mw+3A
f7oQ0DKAzgn/FaV592iMhORqehzOWHwTDXgPuQfVn6IKaz7VUHNq32zgUdBDyi6g
x0BhfoQcRTFIcsJNBZq0dmZzbfUC9Uur9oQeBMC1lVriYBFuSqU1znzJQc/EVNR9
LDM6PNLESMeb7ThOTxwqJ0DSQHLXt7OIPrpf9J7OuDiV7Iwa0hUe3Mqup1j1isJL
2NhtWZ5ZSZON6FLm2rnGmj3TcNrrD0BwJ2MW98V6rCZQGJtXUNR/y9cyywuPN0u6
0O0yAg73lk9ZljesFlvFX4ZgqAWwowTSRk97reoxU0XY2b+TFkr69djMW72jMiCf
PZzqXe+cl1IOKJHrCESPqJq+/ok3C8fY/GIrXPSyHOyYr5S2HXHj5zA0KZKe6n5+
UCKfN5hMjcUVm3MkM6HsfE8mLegV4KwvKXB9w65nCFNef/FiaJk1xGnfaEp+Zzwz
lWG0wpjazcO8tmC/5ijxwCdf2Ii+8DA3tTZGNSwYBNCoA/5bFzYOx7xgKBiINv7B
KlpyhQCrtTV7njLen8jT9HJVuBLnTscYdaVXZn8aOVkdBZM8byQ+1W0DmixZuyf9
6HNhqgUs1zFNdqmg4yYzIGfe2IPhNKct3v55kgK/IDpwDhkbzXfE6H2+X75iuSEg
o6YEReFVELAsESxzf7YJYDRSJj63IUCCd33T9Ru0ve2K9og0HS7O7O3+i08C7Orb
exExaTqrWsTwQ+K8kaGiRXwQvOmcKrtZU/Yr5xPL+9NhgtMtBKT0LeMAQdXtuwPD
Q8S9uXt/lf6qNi9FiBc+Pe0k/Iru9CdRaMxStB1BsFxH20yxdIHDc0iH4NWQa7Tb
8iBd//dw9wHsv+2IGCU3mtI9OZzRiYX87ogbu4HG+H5lPgXx6GXN9e1ne7c/THeM
r8/ba5TjgzLO5Cw/s+i7YfvMbd+qs14Yvr9i8RhtDd3/uer3NkKSllQgXZu6cMij
1R/XesXVdPIlUpVzfq8UGLnNVgd+Z/9T885HlU74ak5i2+IEdSsVzHaQJ6MG0N7e
xCrERb7l3QHvTcVhj9k2UYBq+HDz/xR5FdsUBhebnwXCz1uNMDhYehsSEqnwZO5a
9gbdqaj1PvFLDo5OHXBc658tC+RjuLI7aCunugbJjRGgOfWE3y3Pj737PN7PgEaw
2WScpQKAQLw9PY2EweFSh5ZQ13HzKAzcWV9cU2Lvh4kUG2+/5aPTr680KWM8iTLK
vbQadb61keuKuV95fHz8GqXGHdbSXJzhTlCWmgJU+x+F2FjMooNwsHhXnIe+SYKV
e9hs3J8I0dpjmFyPUcKrEqkz6HytF1jutM67W7BrALOuhavCJBhd7SUW+ojcKjqv
K0sNAlYTdz8efWqI4kedb6QTWW0BdQLHncYftKPWkRcZchRj+3LNPkqC5ekAYZwX
4nnx4jmGMpsEhBrFqKrVhtEdcNj8mgVSIxLXV78Pj513m421Ml7cNvyRYCtGplxf
KXN4WhY+B2D6H99sJes1yys6YQP8OTlh50ZWDYYuz0n+IxkTtFg+JTp8+Qsut5ba
3DrajGmM9/y5keESrNrTSaFY2xcQOP/fhXX+/fP7E6b/TBX+pt2Z2jM0UUFiJRkt
vKym2ihOzsVzFR1K8rdudFnpCb4E6v6omyYgg46DfRIJ4E/g8djqBLDFRxaVTVAe
bNKUZ5+KhpnZXf1lgSF7EnUyewRM5j3BWDXC7qvnwAJxIJ8oAzBGPwZDUwIc7j45
OtCOshhK5B/YhR/8O7CFAc6Ee1HcvzzlutXqG3wL8gBWfLt/aVLn5LmrPXE8o21e
lCtoeh7Hin4j+R1xVDmtZ6p47iJnZYMcUxtZyFgXuzMqJa+XJRTRHqmjk4jKEUL7
5qGmei3daYTog/0ftKYkQT/MJJhvZFyAZJSOP0Wyzl7lsi6R/WH0razBrjYr/V5N
TKZVm88GILucIC2CLDj5DGRtVy9q19csw7u4/Mjf5bZfYukvyRFBdj4G01NjMPab
XOBQ0EVOik//oYApwMc5pUDVzgI3ENOi8C0GsxnA/RSTDkEsHy0a/eWYdxooKzyy
+7gtibRCeW4SvglJRJ4HAs/5HDRprGUwFEyd/wPH5cDsZJKJp/h9xViD6+zywtiI
eZ8ZRp+fNBoeWOkQarnwm8KX5zDV6Ln6KIHleL9Uita/sfZ4eB7Ow9EqLd7i/Dou
oG0Xe9jN22HNtf2Swxvb8a8mCQiDUvchzJ102hhSgEPyFl4cncp+c3o0NAqUpQPF
bL9LNk9MYy1tSZu11XUy7Ju42KxTtV1wR5VcmG95IK0xTsDwjMh5Ja8SPSMk+1e/
atJueRwwL4Lq+cGCflZqDAqVnXoKiumOXuI53ZLhwKD150f5kkn3AxyBKpUYc28F
fE+HPYb082dUHWg3GWf4zky2HTGfV9cl5Gs0eXz66e0fe6pCxnGvsUuhbSHKjCNc
QPyl7sFIZs6ICQUtU+FgA1rrXyFPb4GFhYyUqMJuWcfY2k6M23jRC+uad+LY76Tu
kXooElKWa4Fz7cxFCbPlbnARwE0tGyOkJ1UHCcXUqjXHoAjwXuDNOMKZ4oO5xxvi
GGPVgwYQ/eNP6KvQbqMNhXTg80aVC+42WmtDVW5C7E3zn04UECPdYjss2n601t7K
wbGWa70c03GC17iyDtwJus1yAh33Wmq0HXbLFYKsp5oWgigZuXjNu/HMECpWB7jE
28sJNRjXmbJF2mxsBCkPOGWqhXJxeP9130jZCxou1U8Qs/NBfU/K0/Us3qH7B2d9
pRnDSu8Cm54+SYPNjttnIloPhqOCRCM1tE7orVbu+VtqCdezpGbTKqIoM8Cs5zHV
nIe/r8fYFl2BDf38oFCcnIOyzDVSYPeEviPy4aK1aSdJ1ZcT6AWdvv4AeoLpRCoV
mPD0ypXXPKedx1iLwJYZrUGLoN1MiEwKmeFvNqTc5xaIujVJ3a9kJX+haUize6io
J4pE4fj5joPVkRLRMskvkDh86eQlJf9IMtVFGmcc6BjWEHQdpUO6Pw4nI6KpGRo2
FQt9cb7VtNulErIZa/vgGn6pV3VHe6qz8x9b1CvLqRtU+FpqNzcxQjkNpaTorl2N
wBTWTIsjBgKp5XV/+q576KtE9at+GAOqk41kjWs3Kjr9FymsgCENymNcdt+aoX6i
F9XvLqmFsGG4O8DWodwvaLqVMcvOlqNvGKuaVgQq0CizGukmfJX90d4luCT1QwUk
1jqhYXJmqQFOLdUPvSGbj1WI+cNnmw1d8roCeGRjCUVIiIINIOsLBrZXs6e14xV5
3JP6awI34BWr47DPbivk6UF6iVl41/8GeIw+nl42C5+NOvaIhof9sRClZjPb3NSK
NZgW9AcYBqHF5MY0qZVFQXjOPFTYZPa9jmgedwRiJPnKurbx2xJiHQo66XzBpCcp
dU9gOXqcYWzxslA5YqIfRPlWPdk9i8ZfTbW35R2H7IzsASk8vk4A+4wuvTvLmmw4
HjWzeC4yqeZazKcENhReCg0Yd9teXn0pdySQNtyCI6gCpeE5HgslGK5EhEf6gp+1
Ud7YcmWwOYyc45+nZCLtnR1EZ8dEeeFMERkDJc4frS+WwvNQKx6CMSaq6uhuopKU
kV614LfcBPKhw//5RIKomBkYPisgHWVII3ZAVvBe8QptHUCsCug1Eg+O4u/7gPVR
o0jKZw0ITvssv5qIxUI/YAiOakK0Sg04sWqCDWTfKG4SWKK8Q8GoXfozZRIuas/Z
fn45mCYuckTd5dYel8AnfmwyOZ7vC1QjfOW3sMoeTHGO4RaduLbkPyRI7PPT36ZI
zBFrE4JY3+Hr7EJA5RFmc/K3kmlll4WDS5rJxcllkvSOF/NQnQIWkxeE4HDE397O
fdpps/L0xdVupiObxpuYjIebGg4t30eJtMYXfuzXoE91qlyXq0PF+f4LlbWRvTSX
fmkLjD4wIaDIN/itPH3njAv5gN+s+PfyIW0pDMyJ3FCFJXxeUgwNvf/j1vJcQ/tW
15nZ4qavKRlRE/2MKjbByJkV4c1AHs7bAfJxBhVopp2oVvw09dUBCFZb5GUxSvN5
g0p1gUo5Q323Y622d0c54qIxQhHX0mDt9ATq1fEejoPhyneDID4yYajluMNd0HYl
hC1s/di8xojf3N36silqE6BX0qZwOHGySiX9dthlymW1U4e0zNLdDZzqkbDfHgGF
hgRDFOWDvRMClM/VFyQPm0kk27YsDALGKPEvmqyM0J7UYqQjf9bgSJsIMz5YcSQS
MFmxY0+gjan+Lsvpu9UUNT/9pPsJsqiMMlOfOKrxECRmWAM5LbGuOzL/+v+POAjz
Uu7L2imX4us1FAbKw4XDt99DUQV2R+4ucySN+2+RWAoQMd60ji3PhpCVWyWMDag+
vA9wN4jvTvZ4wSuJ7hLJ/dLaXN0gbDoEWteKuduWhokVlzMs8OJgkYRwWdL1ImbU
+w72yCqnQyIhI2OZIyTazqr6EUDhUWl4CQCpwMfIuD1NzSx8k8KBBsgKjydKOkUR
ri5ulJeiFS6QcmVyRKyaNwUfOBrtFlv27gaNeH41hlGLil32j3nSFx31eLy9UvN1
D9WhcctQKzuxoNn6prD174ELOUL8SuQwmIy4P2buES0bYdxVGW8DsiE8VVG8k8do
PfASjDi8/HVfeYwNCUaqhZRfMcSihkEt7/a53hwWgc/ywSTSDiQmHWi600kH/NpY
VA3z72dvYJACXz765zfAEq2U92HrVkosb7M4pL6C7lFmbgBcYEAE4J+BFfaMz6Ur
ZOn5jeDuiLdVjhoTgr7zLvrDqHmWvMQ8U4yITFIy9BFyE9MtfLTl15wLrA/QLive
E90m9kvsYoj5s+77nbX08ufhw0OOK5bs6EkkOQJi2zTrpcLPea7MRKL3iK+F6gcb
e6AO39QCnDYN0Y5K+UhN4miy5PRLW7XLB0J8yqgJyS5IxKaivZjUQT4ZnNWg+ztu
43DHoZD2OMb4W5SpfYteKyOPU5PvChlcZIUyi6ICvlFBVKznSdr/XKxhBfwkk58c
SL9qTH4qgItNt0yBouzmH0GL/yEC83+WoS4hJshO4mPKZoyuuJQR5hOCrUU3WbEl
dMLHqxs7o4WcEPzJgUslUUrjaMqh9ayc+nAGgL9H2ueCBeyd+kVYADX6U0eeEIJC
d4keKhFXxNQBkzRgIuMiyprRgL9OL2V5Ic0k9nEYNFPu7XwN1MtvoMqHBbJLBVjW
oxc1c+UQF/gezd7OK4kl0Oyhad8KMFvJgMXYKN4MHaavLdoeFbZt7LzcgF64bTC7
uGGY3WNjcDUA0YTMoDShV95bVOSb60/Ly3ZjMuw9q/LUgDpWXHgWF4urTp8vvbCc
ltS7i0caOPinW0hKbc7dxUC9Va8+NGn/zp2uBmDNqgoNlsCnziHIBPMYZzaaAiBJ
31nqcwnnoMii+7UKQCq19HT9BZvOBvxhw2LFOzMjPW23dR/WY2jbhowZnoWB/hSV
NhOTs/neBJLYf65oh5//ZnINHmZ+fp6BXFlV53Fy96FNo7AvvgHYvjnstFzLLNht
5hiS5/emKT3laR7uno6ijlNA2D/wIV0DOKjbAU8xjuQsaodSCree0qZqRsJxb0Bl
S5YD7TarUiBKlZlLPlWyvHrrLLTnWz9yoBKgnbZC7mVSvlN61l2iSkRJ27Y2g549
HU+qTWBFlMMjGkNTE0bWa8ebDjH0ZwAlMhCwR61l3QoXGw7XetPZQdEOGkcfEEg5
XN6W8+ASvVLa8EXY4ZyXPfWWdZAnMswFhFErqSbgCdryCaT4kWoAqs5wJyhDIz1e
1dAVaZTD1ccI6CM5klbFAitoZ60oYb6SfIoAlZpyeyZWqPsGaFXYjqjBCPJU0tdY
mOMhaDJcOi3DUbReni+0DzXPUN0QWoT7UMNg4hFG6safypHr26hFbhXXiaPtl09b
CnK94Xshyf8GyMzqh4jpSLvbU8OGnhrf+tA7EDVhub6AOxWxBOfYEpAJd4ac8+sG
YOp9n4yWRsWQsMYgq4hRdDOostRL3SXVfYbHuVluMFi6E7JhhrwAgrepSWRQpsem
qHmb7IKSRbGX2dk53RNmBekWygIGryDp1cE85iUCEX7EIhbMRz6r1WdOpv2yzH/u
3uTrJLK4wDQBvNS+GBw1vS+qjCE5zmwh6ZnksxWK1Pb6WGXshd6GxHWeCJfDgqNG
gIr9uKWxWjMalPC1fOFtYPcm6LcNOiG3008RYtAYoZUmlhdD7pxjPo7wpn6HTsx9
XJ1dV4bAGL9jF3h1K1JqUQNix1GfxVsyTQSXU8p3aIUSkeACxzFcB3/zJcjpFcqo
4J4zkuUIhKKp8vr3wyDJavnE5horE9FEdcKMl5TWEWR7UzkEc3Fbid4qi06zukfk
0O2I/u5veGzJACQXdl1v/RopG07uET0lNcAFZ/T70Z1TpOalCtwIz2IdHxr4k6Gx
jZx2pMOtTPDuRCtl+F4y5Q45SxevgT8zhy6pm8qruKZAo+T3UIJpSdvQyqh/YDcs
ubLdOHyF5IfyXAUT1TgmjO+2TImDSRiQu6U2SPNPl3tbQhG3j12PKjDoLD944uZE
jg3avBfU6UHAc++3YGYtUMiGo0Gvjvo5a7wEJyJWzqmkqy9iNNUSUIqFGS8RBcAo
CjOc6MBQ42wZQubin0/eLjd5Kc1FQZwEaXnCY8sxB8NbJgQNW/lNy7PCMm19SBcG
BFDSfPXiSQXZoetqRzi+a/o7Bcl+wqHKSbrQmGxpU4lWoMZwYvX/SdT816PolT2W
NzdYhfAIP/Lz0BcXk083maPg2FuHYFKc+y656/GekfQBNhyAxGMzWHe7FZor9qAh
/ky79BH3JQjevkHjuMuW+QWk5XNYsWSJxqqceu6L8xLmovwz9rYJ6lorYnShn96a
JbqPCw79N1OPOisqFZHPgn6GhJw/YNT6uRJYtud1147MEcMDgQkqBCATlFH/CxJ+
JtjATK63OL0W4AN+YGCp05nA8e114R1s6vS13v/3q/6AmD3jaffGC87M15ICIXMY
sImU2rEArsJiueYpfNaIIrNieAy8V5XvE70Tj1SVdG1EA+swdAN08/670eRRMmjT
r5PPvPwOGLOfZw3PsnG/g1+i0WsMySWR3z7qXfX3iy/HR5YADzbqtVhEo7iGhFUs
b159+GTqYT4Au2+G9EY4w6iIQXYm7odK5yxQo5LFb+9vw+kJ1EhSvECPxyrpB/OX
t9QP4crbFGRItNct4UGaRpdJdzir5t/CvhpX19NLvJ1YGlEJsTzqI05ifOsQWtmk
Q4kNf0whvq/lSSA9hVNXwnAj+MOlwwDdPlV6DIvdiseij589Tt972i8dfNVLY2yd
`pragma protect end_protected
