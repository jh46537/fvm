��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�-No�?�j:C�]�;�%Q7�jZ䒦�xMd��7� ��Zw0�]���	�Ϲ���f�0{-���2�`虁j?w��؜DP�'��>������N��܃O���~�/n�1��x�6��p��f�g,v���"*�Aw����g��f|y,�1D�?z�-�h�Ï���N:��Bp��j�
�-k�g���N?��1��Fcq5)�jċ")�g�V��d\�N9H�*�ۡ���==u��Bt��.(	�$�7h�����D��ë��=��ʩ�  �D��%��NS���5�i����lP�Pݯ�@��Z$����s�ۦ �C��ZP{w��+d�gJ�ZS L}o��w�ޤ���
����x���I�J�З&�$�Ē�{��r޴�7�G�π�o�����%_�������.�����)ِz�.���8�f�E�P���du��Q��U�!e��Zy�<��@�֌�<ߔ��Q5��s�B����G�����9<{��0��e�@�q62P�l ���ݬ`ɫ�c�
 �
�Yً7v��_�N�1H{�c,� H'q?�*�������ô&��wn�ML#��,��3���O��:��[p��`�8B�1�}���U��O�4��s�~%]�+'\GG�_Ocv��(Q��(`��@�]^��G�Ab<��Wo���kh�e���+����<a�s��K�ȾXi�[Q]z��Vj4.�!��r�������F�ե�!�d۴ǲ3@k4�	����=jE��\9�Kx���gMO%��]��QX<[��@^�E�.9Ikӏ�3s��q��Gʳ#u�Z �"L���X?X*$ہ�8ĔE�4k҈z�5^�Q�9.xZ���C�#��jC�u�k�
ߡ/=1�S�[Kzq���a�%~��S(��+ff��n�;d����r���^���(������8��[ydW�{����2�����J7��z��U���i����)����9
�b�X0�Lo���b�,y����':~�����d�5��:/5Ƶ���H�����d�@S��3�����Ee�7kW�$�<*���,~!��+����W	��-�kR]=F��6���aw*x
�M�{��+_v+���1<�~m��p*�4C�ՙɵ�|�j�����L�5�m
)�+hAr�T;b�����{�s�����VaG�Y�0�����3�78`�r��<_��71w�[A�J�)227Ƶ��7D��U� �l~��`��U��VH��HQ�N^<��t�{G���"-/_��xL�BU��(�&v�*����X�@?yɍ�����VԽ���	���>Z�lxk�>���ۢK�	͢��yl���0vT�>Ä�8s�Ӿ 7p3w���Y, ��.�M�ľ������O�V�����#����N|br
�ׯF#��Y�V���E����'����)��(�h�Ci
����dsn�(RV��������a$�A\�M������
�ta�U/��(��Y2\Q*D��(�Uv^(�ZYx(�u?���MȨ�hH5�׊[�X��a�9��D
��0�~��ܥ���I���n�����訔���y_��ʍ8�P�.i�!�e�;��f��m잮*��PJN�i�Ŭ���}\
���/nR�0�)���@2�31�X!�)O@��|�9�_/�KD��tT��<ǟ���>�������3���H�H�K���7q(�nM�[o=J�XjBB�r�K{z[�3�hS�[����'"q�0��<���+3	�՟��_C���5r c3L��3I�9����nfI�����(/�}@�R�����%`Q+Fw���f<%_-0tFO>.�f^S2e�+U{��6"��1�u�H�hL�XƆ�ĵ�ʹ́�<}��eXF*:��g��w;�8�Vt�0��'"k��k��ab_On�r]+yNg�u�4,�>���h���l�EF��.R��x�Px����XvRR��lW�	?�KYv�#	�0H�='=�*�]	(9ɨ�)��1j������e?&�a2ż@��
a�\(M^�<&2�ik%W$)��
{	;��A��I�z-�"���:�O(y�O���-�������^C��]��� �6S�B�*{� ��`������Ա���$