// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:43:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d7XmH38+qDiXlh0aJ2Xc6nHG0g57DsZRuZIV+rWsK6vZOIFiHNVxaZPMIXqU44as
sLDWoDQiJMkI+ww6s03eNpV/EHsFT+be9X690Bp4mNJrUWkFFivtfxBywp0r3HxI
vRsrOQYIF+7rJQxYRr30GSG0dXjoR4tsIXZC1c8jMzs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2480)
SdW6/XWHJOwAi487/3LDbplGW2xy1o+a2V/+3lmKpzRzcsRq9zxd//VPhIwHTxf2
4M/RhPmGNb1jZETPWS4mOksbF56YbXRcTXdDneZ4O+DfDiG+cln0OAmdPm+68bh7
r3Ml8BI6vpZdY4MvA2BfXOm3mHfG8S+BWfypA7HJJIVz5uxth0N/uigbBU6+1Yvv
pfVi66nT/2HRT9y/+QD19ktiWcd7Wl48SHRI8aagORdVXIToheWbLU4SyU7sjOrb
pOA4/uhEa0dFMuZYoChWmW0uK5H9yBQffK13VAzZcxjX1N4w6H4/8DgeyqTHymmQ
wOqvWDeqxmMTVhDeaZ4ANw3RJ4+NwkmGFdgKGoJcEdeThTRIpeVmZNpo1sTtI0QG
emqNqYSTV+V/RJziRLbNxzJVdhjVx0/j9aEntpzGwR7iqBMT4YXwZLG2vnXLO5i1
Cnx41oJWizrmFwJMKnRZa3g74V73gc7ZU52tra07byyA4w4wZBhZwwTXnMwdMY0P
Y7fFl2z8gIGZxuTiCfw3izgsGw98FKtYca7iDNTR3FTdsEisw7K5d3vJvsTQE/oE
2W+WENjeMHPBugxSJeM/AYjd5h/eY2jh420tyzHJPXjmmBiHpIRjW/aHy4ltdz0K
QCRYxpugm36wBDlaikSAGEc/Y3KhdOgnRUb8JwQeTVPN0PtaJbca15ZDdmG70XB0
LF3g1K7fp2QU+P/NNXkj7HnE2jaUk5/elOo2Hi69exMNyWXJSYQNt7YyvtY06nJW
37fG0xdB8FF3qOcC/XFCMtyJjJ0aYdFBGIsPIPt/B69ce8Osl1VnmmgkPoH7JQa5
Z/yzJMG1ulgimZ3Hu8kZVHyzFGLhKRKznhN0gF8LF6PXLXS1e6yPXN2mxYzB8uGX
Otae8lTdxplcCklu3/zAlP7qfw6/SDiiQb55pHOET6+Wrc4Nwi1uuxUojI+5UGHk
9mvlhBx6LcylvzrwWbQNmRHtVWRtgSlKZnfLmbZdecr3vC56berhTw9+TG5vflpy
wcII2q1PibkfBiq8OGnngCJYIXkFhyDFHh8FTZWubfv3f5kHnk6mI0uuYxRcFqKz
n4sSffw//738y+3um4HluH7PfcXaCfHurWQr22GSdoQkE3Bi1RSHwQAr50ntaAxk
N3x4Fe1AtHghi7eJ6CD9EbrsOEt6Ck9LeFbKKcIEzO4HOjIWu5zEAthEs3eHE5Vd
zoOJMP2CW0lytmlFE/Re7Lb307g2MQcVL6xQU8wy01svx3iPWtyTtTrW0MofF4Ee
zkhzlZninUH3+DTCr5PIDo1liv/3eA54/GRK4aGvMb45O06eoHhyAeQrXldj2bnK
XduC/aWicR9wBLvgvhkqI3csRTP/nmRKwH2OpJ+5IIrKx5VxWXDzJUb1xVmnO4Dz
dlt7g2abpUpM4B4zKehDZrPSwzUgWDwjwIEYi6LMoMPMgxxUYPNryCR7fum8nwOc
p9S1c90uAbbYMAqlXewE+zjWSfIuXXYU/O/ReF6VdaMZqHKGcct9gO94vkOnS29N
7KuHAY9RRYSLqjaKff9woRnbLTW2weNBd6skUQvb8SR9xIOaPFnZQpUTSwIOyfKy
ScG4HsT+wh6ZMbO9nqZS/hpTjO8Ynm9YhnrpkIc0RRnPPvN/ywCVtppBDyliOf9e
AohUFMbPScqKnxXd7KCAS6w5H/m5P+bw98eYAmgnDQRyYqETk7VyNFL08uYCxXEk
ALxQ5xW5lApBgKEexxHEHcygJLuZx4oPx+u2ouRDFCZHhnakc9lClZIGAaTIAkCS
ciHzRpVW4ctT08TNl7j6/uc9DRI4Q8Dq9fbPx8uAzRllvejaFMRdRVxinx6C8+99
s9XC9JH2CmWNuk0nrLpfLIQ2Yk5BQkpPH74CK/a3iTso8Niwza9P3fexT/ibJENr
AZSScuyq4EpYYZM5xb7AbYoLqdvqKacW+CrVEg13XqgBynnf4IQlftiEvwc8eRg2
jgje8QdQf2m2XStd8WDC2cTCrRWrDcRPodg5ITvsY0tX8JoITMEDtZctVoZ7HQlh
xFGqYJ8nplH53yO2EXvLtKn3JPOHHgFtxrdHWmDGPjyVYG0QDmW9XzOQi3qsAsSG
xynF7xoWVEqeGBoXEpWLK0xUrcZtjupLqhkH7nqmR+HkS9Bz7+d4wLrDnrmBXoZW
pbRtZ/VJUbnRIpEv7tAeBqwQd3+hU/RJz9t00BoWuHgbWCOwUWuN0Cf4d58RXEaw
5hQBLc8ImEdXvC+fxQ7bZqXZjUlZ9dJRW5mii/VXaMzo5VdKBrLpjRsNnL9ehYb6
K4PKpiLUM7Uq+ISSIWXuPOXal42ljojICYcYLhEZtlwpxZ1xYjQNK2AQqYaI/4BI
bJoQDhmDok9wFYqvTLhRMk/Rj1DMJtyWSMsBsFaA71bBoGxLPYsIykZMaBveXqYx
FjZzuiRf588+2+38guVkfqNJWEllNRC8eoke/D9dfjG+z7P9wonpRJTHmQYoasf8
adVNWmP1eQmXMFJrr1+nG61fnN48eArk0Ooh7s9EHSz2LPMc0mglXhSoN9x8yb2q
w1AA0cXT5C2/hM//j3NKNGS1nmMiN6Ug/mf3up70MRJwRHamuP8ZXztBK3BUIAmq
fG4QwrORXGx7l2JY0PwLiv2nBp4SonVP/norhgrJodjBY5OFU4oJvmqcvQ8K/XVx
U7Rhntr7qPTp9gaK0rNXCVp8GQ1+f012d+2TSY89n90W7bttooVf69jJlsgkqUSS
nb36R4atR8Xc9+R8NhMnmJVVqJBDekajhlIKOiSZAsIqqWk5YKZA4NPnf7jnOHPz
VpcTaZ6BYv1IswAKCC9qwdSpK+o8gHgrNHo0IJDJ3ddoppzewcxeOlvhWMg4djuA
9dV+GxIUUschpzit8hcN8wo4nS6vpnrH/0ict9GK//agFwhn5ztqqSgpu4c4GDPD
r8S4gI42C10/rCzaBi8YfWmoVtYhU7IYGw4QJmgDzW+63k4P/wZOLJ5En/XpcYo2
qSgqsgVUheGpIVjsBqxmOUtVOr+SpNGnrzEY3/kCMKQ3yiJLDvMm7TsWikHiMAxu
RTuM3ddeDv0PRDmRx+74Q0XP28xCRKzJOCiu/ONkSh5CmEq5bVJy+e2djQTO1VAm
l6FwSOnD76VrR1ZpjNmMAVyTjAh8EmS7e3ohFCE4FThq4i6HjYb7PdGR6jHVvRUN
nP49DZwVNYa2/JfMeqoJS0JuQXlGSnaRlOh4cjg5NiE8mtNPcXAVtZLJgGyFBtRo
W62FSFE1cOzCKJ815EEq0npWIkKk90HVzndGWaeBc2k=
`pragma protect end_protected
