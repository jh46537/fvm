��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�-No�?�j:C�]�;�%Q7�jZ䒦�xM��P:���b;Ȋ������qDC��A��露W�RUa�X'wj��:��ݒ_�f��~āI��$n�~�б6���/ڠ���L����"��s�?�Σ4���(^��!�H�d�^p�t۟�a/`���X�D�AF?���������G`��_��"��FT���ٶQ���%�+kVw�xh�}�~��os�娂�U�����Vq��عs�;����U` ��A���0�Ϊ$fN�����Ԋ'�g�cWʹt��J��>��xV���֍?D2t(������`��FzH��s�3^ݔY�>,GU#��b�V@	�_��4̢5�^̊����[SER�����2�>Z�������%*�$vژQV���G2e� �ǣ�a2Fd���n���.��L��j2|�\(� ���QV�_�����ph~�K�=�WR@�s�E4k�=�����j4�6;�?��LtR��Q_&�'�-9��o��l�|z��Q�t��E�.�y�/`@F]O&�~K�r;�{�zC�K*���]�H��O��$��'���^p9�I�`;��tm���&�����9Il��
R��������Hv���P� 2�	�/Дa4�~Hfh"���tpp�oB'��1APy�2��"&-�T5ĺ���ȴ��l�ĥ�F�:q56)��=�����t�t%���׍���#�۠�Z��wQ5ɇ�c�E�{����7��-N2:�*2�k���gا�jiN�^����[a�Q���^���P���#MQ���o<�uhC�#8�P��s;R����< {p��1��5���HR�q+�����}W](]��pjP:�ފG�D���Huu��:^�Ȅ�Fpu�Z��a���W��P�8:�L*�͑��h���p��#U�6f�+D��Z�	�O�{��4P��M?�Xe��G5��V��o�����{��a����J���9�[HMr4�Īӿzվ� �04�2Y�3��Bs$ZCy��3���_��d(NT�8z�I��C�߰j����%��;�?P
�C�R;�? ����U ����*��^A�����iã���_/B{��r�µ��s>��\� �0~�}О-�S�z�Y�C(�z�_9@SU.���``��BC4V�E<T{PP�c���1{:�c������b0�bp �0��4��Ń�|$~ڡ��A���ʹ��zj�:�2Xh�:�=�y��upa>r�@���p�ĭ`�1���Flo�����-�%3�\�6[�)�Zf	>.`�v9!.��C�H�qE��"$���Ϙ_�g[�/]�o�Hؽ�{�I�"��1b,*���,4���ARrr(N�^\vS!�qt�{\�iu�8�h������ZU���ՉHW�wq�$�&F�t�E���G�F^7VC��˥�X�I�����ݼF�o�{����p#�{�0wz�r��V���c�����u6�50�G�1m���6n��JTf#����а���<ݶjq����z����+�n!��Q�n����0��=�re�O�Y��{�ق��/C���Ae����	����N��.&��}$�J�Mpst������0�� ]�A�x̂*:H�$�2g����&^s����H]�`q��7\'�p�����#�f� �yyhDf�ޮ�r�@��8�]F1� ��u� ��x�t������}���x�PM$��9Z�.�����Z,;��/�8��8_v���5�ݿ�V�dN9b�gJ��A�=ˡv]�����1:���Hj�g󹮎�];q������
D	 /z��g�}�w�p]hCaۘ�����R����w���>��f��˯�+�"�	��G<]�_n���H� ��}��p�g���s�Zv�D�W�6������*����b�.����	R�#3�*�Qx=��K�yk.Ń��V,���7BD ���ֲ����A����E���%zgOR+*k��: ;���o��j;Za0 "X�,���z7��c�\8�~y .�}Y��]���<����[L`�$��fw݁7�QnJ��!��ݧ��f��KN J�[��d�q��9�K����c�9c��p%�N���O0�����������4�