��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9�/L�I�Ea<h���	ԎUӸB�z��V�����T�T�<��N{��+����)�H�gt����M(�>_���:�'`N���wa�)��هQ�6X���,N˛,���LU�{!�x���qK�Y�=�w�▒�ґ,רv� �����za�Y%sP��%�|�&��=�U���_�Ql�o�9g�Ws,_/9ڍ�����Ce�2b��h��Uab��V��R�?�jaN�����Ιjb}���f;;Mr[S�*�=���`�E���Mu�����.?z0熯�A�"'�x6���锴"�9��V�wq�O�3��r"~�Õ	�3���pz�:f�*f��2`������I��C�e�i!���R*��
���᛿�1�����u6E�З/}�F��+�^<��=��r�%R]ihCy��Uýw��YO�i���t��`�2�|��]��:.A��I%� z,�ɊX���v��S�X�S��lSR�~+���F�ȡO�O�=�ZZ��k�x�@��OFs����)㐁�&�8`l7'&ܸ��J���׶�\ʚ�5��G�����jW6��דL�2���66G��ӐQщ7���Y���8�<{�u;��V>ٜv�d0T�"��������K
�_ѿi��4�E]N��@3+�$�1z��8����zC�f"�Zp	�l,��:Q�c���t:�4�O?��}��VF<�?!������,�6LY(j蜈�w�ؽ�C�C(j_�	����f�]v_��#��<�S��A��s�V��l�ի��j�S�]N�݋���N)F�KUf���&<>0"im���5!�5�f?�����JG.��>�t;1O�2���Bi_M�t�ER+���.�T*�����9^�B�J�Mg�� O{�<�d�K�I�3$��q�ҵh� �x�C����2sĥ������F����O8%9���W�v ����E�6�x�"�o	���TND 9pc:�<U�?&,c�E�%O_r�=/��%�5���`����5��}G(�R�c��@7^���Ŝܒf����QBt���`5�A�=k\�96!Ŵ� ^Kȃ�/&>�:'$�Z}MZ�E�?Okbk:� G�e�\�0`"�R.Mн�$��'-����f4b��N�O�~�]�7z�G���qL��E�Y��&L`�p����"��-����<B�3z&������T'�qw)GJ��T��}STٌ���*S�T��'��s5��o��+�9R�Q�^��E��R̈́��[�t���8S��Ad[VJƧ��>՞J�ĕ���su}�2����ֻM�	�)�����C�Rk��$J7���8���RH���4₞�X`��rt��2�����_ೀc|3�ց����hw|O㍉P������
���iOz�hE��YRV����B�$G���ig\"b� ����l&��3pD��-�D�2�悊�̉�1��jCQ��J�~��C�8;��h��o�@�k*���deq�m��V;�;{�
����(�
�]f��@O����5Ϳg��8OTQ{�w<ID��[ʝ#��;n5�k�C��N�$����0��{3���߹�xF`�w�[20�����dSd�7�b�0=�/����;p/qoϏ���!��J��y@��'M��02�HU�������ה+cۍ�\M+����&�If$1X��wK\��	6V�U2��m�u�J�������to�yD<�Yh� d�7͜b�͠���Z0Ю�.+SK�s��&����`�h��]s��p#��`�M0�jN���9\2��L?�Y��'+����{��À�WH�T~<�c���a�r�Ԧ#_�غ_�^�n�Qo�z)�Y�DX�_�<���߼�ɗ�������2j���
�"���	�8�(]�G���	��I�� �4�m�rV'E��7���х��1Vi�|����(
N�0Z:�'k����Q$��џ�_��D���d��2�qi�Df�C�שF���zM�r�98�􊠷f��>𬖐��e<���" Mu]���óW%8���9o*-��)w��W|��!Wz	R�Lh3���|Ƙ֋���ڭ�p�������8R��
�i�$��dc�Z�^+M� ��5ޓ��B[LJ�������,��j6n�sH���Ea�˜"�����g�a�[�1����Μ�G���<��O�"֮��P�D�F���
�	��]�M9��i��3����睮g��^ŨT� �+���l4]�7UC���äj�jX��>�~d���!��T-�5U-����!v���W��	�U,5 ���h����v|%G*�E��a	��i�e�@
lZ�$#�*��g����قwDT��<���4���<+<]o^r�-v�8��Ј��2�W���~�'�i����� ��*KTQ��w����T��w�͉G�Ӯv`Y����V��,ȼ���7`����z(.����c-G��C������i�1��=$��&W�+tV	V�����
��������rd{����%1Uah(�q���G�Ԇk�q�Uzv��H�bM(F�&��V�X��p�K� �A���mk[f�� ��{�=��9���rm�w��])�X���ْ2	�$�)�ԭd�����K�	x)3�z6�T��}ۻ��-n�0��h"<y�OfT�j�h��`��	���d�/x�ǡ_��Ŝ���bel"C�c���1�S&SP8���qO�B��$��9��&5��C�[����_~�k�<�#��xӗ�"�$Y�8�(ŗ����U�Z�|a���v\gD'�ohs�)���?��%�e�����X��dc�������3&
p���V��y�;�?�"f/!r��Av;�����'ږ*��i�}@�K]����܏3�t�S�l�Vu����{0�@���;Ty#�:\<9[�x�	�L�`�K���i8�s��A<IO��y&�Z������n���b-�c�"�`�e������v���M^驎�%����@1Lyrq'��^~�Ӆ�_���U���j� �["v�AI������Z��N9�('=��-�j����;S�gs�_��q�g�Y��ߚMT�ʠ!4 �m{p��J�2:��R���ܐc1�e$a9����4M"����oG��Sa�ϼ��nG4���/��L�C{��i��X��v�e�C �y
�ڙ)�pzSYTò��Ƶ�K�( �[�î%ۭ��C	�H��A�A����$f]���R`�\�JK��7��Қ7�pe9����N��f��Ai��r��?g��&!�(C�g j�0,+0�5����%m��*�U� ���z�e�9����;U_�s[yK���,?	�����%w[zl�qk��);�r����U\-1��%a�>Y�Lj'ܥj��Q}�}@��z��,�9G�����vB�I{:�8�"���3fJ�	���~�9��/.��UW�Ę��
��#��?fH]��9�K��Jz3p3l�fz��ޑIV���au���*��b��n)�Ze�K[��R��6�9�'��U,2�և[�]++;���ʷ���j3�Z�z"���tk3xG�d�_]T��M��T��5i
b	ԏ�׷�H�v��(Ѱk,��x��4�k�O{oD8A5l�F���C_1bMNy�ЉT^@Ξh�3�T� �
HCйF�U���Q8O'8��XP���ӯ�D���a�^<�ؾ��i����R���w�K��_�g΃u�k�/7�gJ��SS����� 7"����V�j~�95�!ޭ�����k�8���-}��e���}���f��J<�2;R�]�K�|�>��ߧGZ��YF�Z �M����)�^%���׿�m�����|6�B���4����[(1�)�����	�yf0�؞ ���|�|՜mq�t���t�0����Oh���vV����U��}���{�ɯ��A�zF� �ȋ��;��3b���L�����j<�����_?�d))n9�@�k�*e�]���Y�~�R���ޜ����v�'�+��AA�"�S^x��(&^�zA��)�iӧo|��
ˢY5�ݎ}��� Wm��K��	�I���/.{�����rw�g��6�w�m؞�O�_��7`��]�*�,bNQi �Cܭ��B�]��ȿ�LcL�X�oi'�� :�����l��F\��+KH�����o�#���Cj���3Ǭ�8�9n��>���c�@s�����ۖ�=d$=�%i�+�n�r�;���AG�J���P�K����͉�&[|������$�T�����1⋍��	@&�"v�83�y��趥�97J��'CĶ��TNT(�+�{3�r4DtrZ<W�a)<u�K�:0�\5+JR��B`���:��,S�ܷ�C��B�Jw�@��$/�H�=I ��y�=���D�O��W��*�J���.ف_q��ü��4kJ�q.a�L��C��̛��T��Y�p����>���u�h���vB��)t��-*�-�&Cq4H�D�և��u�7�t��GI�ּ��U��I�gk�2V�"8�3=�͡� d��W�nlZw��N���J���EL��@��U߱�Z(x��$�IE����v, �A���};��;�Қ��jM܎��ӊ� �܍zW��/���t����W�T?�P���P��͉w5�M'ǌ����-�ݻ��/b�ZJe�G�ÆS�F3]�+�z܋~���Zq�'��̤G�0J3�]s����Hߪ��k���7j�#<��e��!�Ѿ]!�]����X��	�R�1nO?$x���E��u��h����C��H��t
���Pβt�ܚ'&[�z<�"�D�=U�sJ�-���~b�����=��I���ɥa���֙ӭ��6��%?+�>�b�G�er]b�ai��H����N.��(�a��U.Su%ן" L��#��Œ~q�N	�VJ�Sz.��R-�i����NJ�i4J���#~ʹ<V��/'��6H��%NU�����+��ע_�%pi��C��@u�ʰ�AIX��b'��R�.���`��['��@#��9���;	!/�5w�^U,d!���n��j�X��z!�G��Q������2�'�tZ���k�פ�t�j�,0����u���G��
�����O�yE�/W��3��˷��-Ӿ�i��gb�N�Z�gj
������U��(���(*cn��L)�+[�n2��3�<���0L�3��&R��iu��E���=FM:����o���Ar���H�,?΁~.�n��y��N���:�ۊ#l�X�}����͐���Jv�Q�>UJL��n����lor?U��ao���=�&{��˄�Br�I�iI�"',sEO^�궇9Ъ�$?p>�|/n�p�0�S_�e�2�=��D�R�r2l�}AB�)���������̴�(��#���̔g�n�(Z�iƸ�+	���q"8b�7Awb��p ���+�0쩩8x�Ci���
�&9�C+�檧~l��q��U���5[������Q��xx�����I?�L5�&�����`Hs�k$@ZL?�q'Ì���e!/�@��_9f��U�sV����ϡ��Z����b��(�O�����J�]�	K�oÍ�Bt����װ�3�E�j�N�F��2� �x1�� ���x����X�-��oi�gZ�W����o��1prC�U�z���ͤE����x���k���llƃ��'?p!@��LD�J/X���n:;��o���m�@�{�!0"�q���د��Y�Db�"���� 2N��;�7*�~�Y��8�m�1���k�&��U�h�g��nJ��9"�����Wo0-�1��qBB$/؊u�r��N�sU8���4�[;s/z�*!����W�d����΢D��/���J���q��L��H��a��%��Է��Ƃ��@��*'�l�1ݽ��Y ��p����k�Q?M<��	�kZ��_rF
O�һ�h��R�s�����&_ۊ�h0��
&w�0�ե$3�MqY7v�EG���#J��J%H�?1�X���@�3TH�Y.���rZ��Hl��e )�o�u�Acހ�,;o�e���m5�i���:!ѡ<3���0��[�/���J,P��l��⽊��M�3JE83:��{��k(��,����(�b��u��}LPc���^����lZ��W܈=W}3'��\n��{`*ť����bi~,(J�>q�Ԟ�8́P���n!Β�wa'0t�P�93�	?�V;h	c�	��l���/9��q�})������"���%��k=�Za�������h�U5T�c5��UM�_��E�z�,�e�e������W��������nP6�{VL4�Wop�D�<q�}�HĂ�Q2���E��ZX���%6�����1��4��5HK��q�մ�&�GuU%����X�z־ǯ�`�C��� "�&C�	ʓSV���z��^/XXh��{`�5�j�V)�1�,)\2׌�r���@Ӗ��-~�B|�l;Mu�Oj�f]OE��gb�~��w02�Z�`ݽw�]�T"0��)���F����tP0W��ȇO �gS����5/��k}RO�i�Y�,��eH�2��f��KH��l�e�O���v�l��/̗iS�Q3��c]�5���Q>�}B�এ�� ����^TثZg��!t�!���ED��ޢښK�Od�n��,k��\|.w�����:��EMĳC���_�L���o��%��q"�}��"���\���~u�sf'��S��v���ef[.���	�q`��1���dC�$�p@� \471	����m���*e�0(��_��ߘ�+�2�z�����睬y����LX�`J�q����>��[�Z�./�5�<���F46��=x�[f\M'.�Y�faN�u��ɞ��p�x �|6RUxe�G�HS��.M���C�cm�S~��Pɩ���]b�.Tu��v�;��ɡd?����94��~Z����;�F�&�_E�SZ�(r�+cS�t�qdx��0�/�xwB��Ԩ�8�� 8'��O~�S���w���:$�6�����Q�ծ�?$E/�D����\z&��T,3�����O���i+�S�#�b��gNN�BɅ_��*L�.^�؏�'�q&����v�x�W��ˁ���� ;Y/��r4	:��t&k9`�J���Fj�˔�_=S�,ʑ~f��R8µ��ry�~Л����=f�������R�(����YN��*�
�_��|��O�[��N�~'ti� �O�7�]�2<�E������G4jz�c�̆�!$}�8�����rˏ����ʿwK�t�j*�NW*R��$��xZ�|���]@��j��-�A��RU�/����.B�d�:�����*��]��g�zz\�Uz9��
6�YT�
�A¤�[��R�1�������-���4E�?[�S ��o�|Ȍ��h-� �(	������j��^�t�E%��Z����Ϝ8�Tǭ6@��zP.9������P�m5;'�\�.3��9�����Ͽ6� 24:��Nv;��C������� ����y�[�$����ʠ���,])u�߫�1��c���r�X��΃Śr���6\�C �����C.��]�e��gx�p�N��m�>Αk�ff�xqt�L���B���h��� ���LӍ��jdh��0Y��:Ҁ�¬����2>�X.�4	�*�xFʈfx䒑��#�"�`c�v�l�u�$:V�:˭Fs?�ra��F��T�����L�����	�'�!� qBh����
��/�=��d�<�8E"�б��:�o�)�B���h�͛g��畘fDp%$���yM��κ�-�G�$`�]{��	5�)]�R�vj4�.���u�1��n6u��A�2 N�����5�_q3o>UJ
9��tN�!���)�8�(1:C�r�8���2�yWl?�Xy�P~��l�vfwH�!��T�]�����ȍp�|6#`M^V�f���>�h��vnR�R��B-��v�Ig�e�(�¦P��+��b�U3��@�jw�3�|+~� l$uS�u��Qm*:I:N�F�&ڣ���e)��W
�¶��7
�~:�br���ɣ� Hi��#az2��t*\khu�p�|�`�"��f"�(.���0�jr���p���U�K����޳��W��ZJ�ڭ$�p5��(�.z��vf}��!��E)bС
\q1Dc�#/^E8� �
?yD����acO3���gn��?tQh�^GQ�C�ܰ>>���0�Z�uߓn�ω�V/Ȧ�Y�����g[BKd�
P��4�9�.N~".��	�����!���T���lx�'Jy�q禱��J�'���C�#�6�0���P�!���x�+q���_���.�is�
v>Tu���|��)8\�6��Q��6x����VQ
?�%�m���f�Ĵ{;E�7�D�n�du̞NȐEbH�P|[հ�3w�2����z��0��|	eEk���1t�q�����P����W��
��c({HO�( 
�3	�(�n�~�M�r�"�mo���郴��Zx�U
�6���mA��xы������<M����僱˜^R�3�f����͗~��F���a�^w,3��42p�qJ�S���5��]�d�q��G���&]��Tz�إ�D�3B�:*������	���0�'B�P�Z��%�3eT�����*�<�f���mr�1�ϺGj"GȪȦ�w,"pC�D��-����m��j�E@���]
X��H;4Y"bo�;\F�U7�e쪆�>r�)�
oY�c����>$X�y��1��ԴdTq�e�n�ZՎ8i���Z�I%�]�.�b�!�'�y\d�Nnʞ�=�V���W��~:�'��ɜm�ԧyK#�A�H�a�y����O�	�X�C�ύ7w�j�Ы�G�pIcl;��q����_Œ�-2h��]$t���I����F� C�;�jS���26%c#�3���f�ԬH�V��t�H�h����<RI���>��f��t������M�	�"�	2�~1�o��M6�p�
1��2ɞ�]�j��: ��5�{Z_=�/������&m���s!��4��X6DZՕ���.�q�yQ���Vw% ��)C3��{A���0K�W�f��Ĺ��h�l�xIE=w��a��;��&¥ˠ�oίʚ��A4d��$�� 5Ր��3�H�f���`j(�`KǱ,�-���z��j�"8[qN���j��r0�	���*mz�C�h9�Ջ��$��PB��ň�X��0U�#X�גQ&؄�����]*�M%~����]�p�WE�sRv�N�0yX���D
��s��wC�����i�~�����F�3��#�?�?��>�t�M�� ���UfW-�՜kJ��mh��J`�k4kQ�Y8����IT���QV���T��M�6h�_[�>��*�4 ��|"�SEX׺�����|�?_l\f�Ai�rw����J%5�.��v����m^�����P���sT93�}`�&P�*�i�V��)w�E/a�h\Kd瘗��n8gJg�M��u)Q���uuO�TL�
�ҩ�/4��$�͕a�}�Kq��+C˕^�yk��*%���srX_�;�=2h'��)J���?h{m�tA����6,V���*K�n��=h>���}.����v����/�@꓿	ַ\Q�>����5H'rz�<{f-a�K�.gv�9M�W��<��j��\g����K����1�c�K���.�cW��p��Y��u�%���7�^J������h�'���/Ut���@�.oqC�U�'_�P����!�Bȝ�R{SJ$�C��U�! RX}�zۨ{�{��>��*��s�Lq�˩�G󚎣I�3n���X�q�Gs�/.��5�8ߩ���v�R�E��(��f#�)fT5m'%�s��;_�����Q߸r�����N��J*h�����[c���o�����\q��� ����&ܱN[�Y��տuS����HP���Y?����"�8}_X �5܌��`�m��l"*�+����N]�*������`��>�9W�sbV�#��8?8��Ȭ��E�/Q�(�⎋D��T�b0MA�6b�P��~=ݵ�����{�2��F���AsXE`f�
��G��c|�+��+ar�(G�����m�몾�j,X�4��V=��<�[�l��,.������,uq������CPHun;z���Q�P�o���������]X��L.1�J�"JPD)�bRf�M�v`�ۀ�XM��L�z*��w��.����EN�X?�β;=�����0м|uX�Wüh2���"M�Y�b�W�L���2y�=���J�`~*�:S�M�7��A��+Ds�_�e��fŬ#��
��ap�!����;O�!��ud,4��K�"��ތlY]�v��$4-�F�z� ���lՔ����C�ak�c T(�֝�� �ߦ}b݄>�'V45SD����{��Wش�<�V�r���%qT���	:^r�P��2���@�2��a׆���>&!X�=2����x*e��~�������W5FMlM�s�_�f���Wl����=Y���놺t$KxnH-�5�)�?���Y��<M���q���y� ��f�����M-�N��9��L�Ku�e����Iw�wze�LN��K���=ǎ����4�3��s��ffz@�9#�Õ�k�,�Ӣ�2�{/�h�ʹT��Yep�6�r�J8�6��(A-:�֓� q�)B+c1m`J��~�w�7r�T�/j)��<�{�.��=�Кr�jh��)C4����ٗ�^U����"[��݆����>9�k�a݊N�^B�!G�ũUȥ��^ :���b@��m���q�%�f��Iz�e�:z	q����7�<JHh\|��ڳ0�l��H1��?I6�g�q2��G�8�$5���<b�'��
�I jLX\K����hn:p��8��I��?H��@b<T��'g]��`�"dF-ӹ�WJ��X�������'��i8���%��{z��K�Z�~����F�Ɩ+k�_u($_�s�S�oQ�I���L�p��.�ڏj	`�:aU�����*��iq^�wbf��Ԡ��@�]b9ox7ɯa�-����-��+��c#�`
���~��]Жj��i`� ��:�m��9��6N'�@���#�P����Q���w޴�kDKu��H-Xp�(lc�["�ͩd����	������s}�.Y�U�r���8��msD�:_����:��4�dq�Q���m����"z����*�^���;��U�@�d�\>�U��I�KQ���!��)�یM�?�dF�n�/B��r���a|�],ॢ߬K
�To�� �Q ��*p��џC��dy�욜��9I��76l�V��p�e��`_;��,�Θn��r�P�$��ڗvQ��g3�&>���>q���3�+�Y��}��]���g�ÉM{^pl��2f8x� ���r��LɅ%�KI�0�K̑���b��~>�O�bIx�l�x�E�*J��zmg4�[�/�P�*�}%������ޙ�Ö��ݐP���m���U$0l�@8�%8�{�֛݃��IW�q��d�e	Ѐ��-�iSů��w9pK�T!�1�?m=���+���9�?R���ρ��A�tA�
[�v9\�kt*v��f�/י�MeX�װx����GO�T1{DrX2ø�����UPqdi �[���um�*^~�E�^��w��߈�D�ቑ��{�@�*�\�5��m�uK�wR�uꡪc��)�4̯���\�ؓ�g;����V&�ʧA����I���!2��H���u�,�id�rDZ����B�]�Y�G�^Q�Iq�E���tjUQ!��]ߐ�~�˯r]yaD�+�p����1-Z��i�̷'PevMr9p�ҏ�ƶ^�x1F]����*��PI�Mf�g��<����0�B��P�b�w"x�Wl��D!T�ReS�����mmj#X����f9�CB�O��$�\���o ��_5�􊁆�(_�ӎm�a��S(Pqew�n�T/ q�Tkxw��?��~���i��_��3�-6:'6�aR�G�h�mb�8 T���FmSϕx�\
+Y���rtb��w�|Ƚ������.Y Pr�߁���\`���3�u�/��<��A����D�n����L'�'�"��@��рWֳ2�=��]$ �S:�Nm(���;���x��G�+٘�����&j� ���oYpF�q?�z&�}��G�M����}�h�O�R�����͡�B��C�S5�x#�d4��-�u�J�?EP�̸wO�c,̿c�Ǭn����NQ4�S`�ݷq+f��c��DmH�%U���"�bu�%�C���e�'�����ղQ�|���I��8���3���Q�;�
�#Q-���Y
�"N��GQ��%&��*���2����M|��L�og��rؙ�=�w���u���D�Z��*	B.|����}�Gퟲ�PU�����h��,�,LI�@���갼�s�AGp� �Wfgu�k���0�r;�$���v���a�͌���'Ƀ��1�7�lɒO����Y��G��m�[��V3cِ��7%ޠQ�� �2sq��9�1��'����PRydK������S�G1���/�j}s�����y@����؇��G^=ʞ�� ���A�\�ʚm�`(���$a.m4�2�����]������Y������o�Z`�1���_�� @Q\õ����խQ�������u�|b�& ρP��c�S��n_��E���/�>Ra�G����(�CyDE9����q{�K�/�~�/ީfi�Z񲽠�X�0��I)"?�f�uqg���qh�(R��t�amX��(tV��������ȠQA.����I>��хa\z�p��?ݤ`����gU��a;���3���_�>����{��C4�T���{\^������d��Z�"�%Ñ��Z���V/LL7R���ѝb��T����I�H􆩛��/Լj���z3�^j6�z�Ў�D��;�ZA�W���H�V�.:��jt"�`XvL#ZE�[p*����P �:��������2-�k�m��+����!�z� �6��Q���I���������T/ΣѤ���Ъ��Yhn������ܢ�lYl���OT�0d+�p��$A	�u��x�8A���;:~p0"�lmI؍�����]���#����H�X�!:$�)�.?��ש�vyj�U����
>�k�5xV�LX�����0�O����?CT�0jKO�N��T*�%9�VJ��kR\�"2g�0��!��)��P�bD4�d�\����0�ɭ���F�w' N�lݲ�d�k�O���lO�%TƸ
~�\�?���Xx)��V��m]�1����������hc��>���m���~��yH�Z��k�<��d;�c�\��?�om�&m�s��]�
��L�DF�G�S�v��%N�'��c�!'+�_'n��j����^~nl�����I�Z�e
u*S�b����c��
'�F��H���dx�1ȇ����� �n L�a&M�����sY���k��
S' �`gCL&�Ӏ���"՚�2ug�ݭR���"��k�����j���^�~#�M�b5U#j+�g�[-	=���ɂ	�X���0�l����Kd�반M��R[?s����:;���y �! <T$	���(4�	`#�13(~�w[��{��K���Uuˆp[a���	��Na��*�������OS592�;�.�4!�˴.��I�u?l �$8<��L{���	�.�Q��ʚ����7 )[X���3��g�m]YӘ%�a�I���y1i�_ʐ�º=1�5����X�'�I�v���n�gɼ����v��'Lg�{D��[�Z1q+�]���S�5w�j�jCޚ�-қ�z��!Hv��M�:����Z�8᫤ȡsK��y'\G��@�t��d��܇��J�k�؎�!��>F�A%�?�Jf��	Ho�>��W�5!*Ǘ���QK�EU��pL0�z���x/Sa���)/��I����:"y	.X�aRlO��ڐ�6�r�F&��H0��A��fכ=�+��5�D���50h�C���-����a�����(�K��1R-;ީ1��Qw��UJ���ޖ��Mʅ�ZÉokn���%'�\��S1�!�k%?h�l����S�j5��A���ru]�,�(GJǋ�>�pX�8 �oa��~|�W�R��{�b�
�u�X�F
׀�T�t�T��ڱrq���5�.����A�=J7D�7�7bK���c�YBvH�k9_��� �uB�BA�v���"H�FMpN�dZ�kY�_��.`z^�O㳲���aXO�����SQ�|�!1|%�!������R���a=6�[xȜZ�s�S�L L�,3�zv��G(J������ظ$��h�+Q8���O��!��K��))��$���;ƀ\���|Yo�q��:�#�o��-^��D%v(Rj��*��yI��r�޸�Ի�)���S�BM�8��ӖHd�V�2П��H��>�G#Q�9o���V/����r9j�F�D�@{JQ�����l�`i�<;J86|X���Oe��d������m1?
ei��_�W�rTS�E;�1��OG���r�d5:?�dZ����D�-J5@��ZW.fZ�.��\��8��G:<�8��<���r�_�{��&]��C{ڦ�̈�wm���F�ĔC��:d��S!�v�Ř����|N��s�Q��uJB��ŏ�hQ"��K*Ҿ"/��A�6��p�]#�or���TŮ�����g�B��r��N�$�hAa/v�p�����