��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#�~�,o#��uIk�˥W��.��-Y�S~d~r�ԖP=�b�8��^4/��1�>����N�ژ{�L$�<�0����pw�j%.����q�#�i���ǋ�6�>�Y/k���[��V�w��d�� s't�"�G��6�?�*(�����F}�T���f�'��	6�+`�X�-7�]�qf��gg,Ň2�{;���r�`�OoG���<���Whs��H�äe�6�k�Z$�L,���p�Fs3�9.��fp�2<��w���c,���>.	�Ō�T��������
�{e@�^T.~�˟-��F�7se?��rc팙ɜN �qE/j4/���-u
��������l[��0
�^�w^p�n3����v d�ظ72;E���۹�|rY�(�Ǜ�Kt
�F��᪆G��ݨxO.%Ժ�Ѫ�V���
L�JIaM��3tIx�vg�AP"����$�ߔ]"
�E���أ�q�S�[;�߈y8Zp��*=���/q͘&��ȗ�|"����12m�N��5�۳'@BEvf_g�n�8wOVD<�*��������Ǘ⣲%ec��S�	P������b�\. J��^�����K��AWaP�Գb����R2����t^������/���%{� y	p��FQz���4�h龦��S�R��Ӟ�K���R���8N������]f�6>?���w��/e'[��?����S��xbX�]4��-b�=��n/%y$��6RR(�E�:�񽷷��Na~��6x�뗗���ȟ1�N��gd�kJ�w�Iy��@8fz��kayQ�:8�튣%��3`��1����A�[�^6
^I��8ʇP)�#�v�*TKm��Lלj�%�u1�7\y�#u�Jf�X3���0z8��a��V@�_��:Rs �MO�җP���X�͛6��6�R�5gv�h�V�a|���x��|�B���e����	����ɦ�{�rO��H�1�Tq�Ţc�D����$�݀����>�r�t��m��WT��4���%oZ�Q��g�S޹�EzQ���8��8^���9zT'ݰN���H�-2ڛS���E���N��ń#����` �<�Y��AlԂ�
�QϏ�V����:�q�[�v�1�R@�J��zR��K�m\Bʮ�yGT�<��#�Hc�|=P�:�J~|W5��&�����נ�o�������|k�.���<jw�6E��0j5��V�t��7��ʣzo]ۨ�.`0.����7]QF�C�P���F��Cmq�_��j�Y����������e�����4[A)3ވ�� �/9rٕ"GoGH�3Y&�*ì��J��F��EG)	�-�O����ޥ'��M�p�B1�e��a���q�E�Β���#t�WE.�+���K.iJ�	ˎ��k/vT�^��7����E2����	��Ę�H�	�K;��A�����Za;*��w|<�?�,C�CJ���o��-�..�=���8��U��R��8��T�����pD\X�Y�y�ў��l��Y�ս�G����l�.�nM�Z`g��,�7�F�ꜱ�L�m�t�@�Jj� 5�8�ER�I�\�XYT�L����Nz�m++E��naF��;Q��g�~����ZiE5�p��,,����R�8<*
a;����ݫv����'0���r�#g��^���hGTa?��~�XT'|���pӚ�yC�z�3z�$z~S,��I�Rr&g�D]�)�1��o��.��R����?H��g��RރG���ԁ�,}Ok(���o�z-v�E��~���D��l������ ]2�<4O��õ��	��چ�@��q ��v�H�ɧT^ALݲȎ�`�gg�
���z���M�D���}���mܸ�zgfROX�O�q<�����H�8lXd�$�Mx�ld��=<E`��9����_�6���R�;:���裟��t����,ꇷҲ���el�imiW�f~^�z��F
}�qG��?�&����`���GR�LE�(�R���Q6xF; �~Y��(��w��.fD�꟧�j��9f�A�3�pG��TX��=*zws��#�Aы�j�pyyx� %kf���C�5���aPW��x�%�2����e4�q]����FP�t�Mii��%4[�` �:Eῲ`�M�#�W�o����3
r���}�}C���8�o�	wB"e�c��*���?k�#a�ҋ�'��ﳫ[�,BˊWN1[����7����NcT��p��<�!��'�,��v�!�w��[��Р:ɁM[2H���3�����'�GJ��` =���3��ζf<�7|�k�˶��CqQEtY���7e.q}����6bIE��5Sss��F���J�im����g��
�2C@	9��5��ޜ�6�}�j��~�Ʊ3��GM3zK=6E�.�����<����3H�ڶ���ye����'/����&�[b��c \?�i˃��:�v/�|�����D�>�b_���rۙ����?�4�+���.s����91��E�IT�/�#����"������<yM��s��a�sl��gd�_�������!m^��jF"�������?d�ę���+Ğ��C0��e�<Q� .ǳ�shS?b;�ky��[�D�����QCb[�WE��K�߻��Yh����l�F��_=���q5kg���nO������AL��h�DMo�����P
B�ԑE��O�x7�w�bs��h���d�d�P����z���d��|�E�����.�j�_�U��I�5W��-vP� ���L~Km�j"��)�������Jv�C'��ha^�Nvd8:3���_
ޡv�G8ϲ�Q>�i�R��֜]�Փwm�
o{����M!�����NP0:p��r��t��::�Y����6S�H��d���[4��^&�ٞ���U��*�u��د�`�[��k�ŋ��{1;�!�f\W�ɒ�C�z9�� ��^sY����<om�/S����䱻p�@��%��9yƛ��'�����lA������=�@�4ߪ��g5�k�T�{�B>��e�i>#�E�w�E��L3=bN]��A�*/�sFG���c e�S��D/!���.���0�o@'�y�� ҍ�%4V�!l$�"����Q�k�����]߂H+��03(H$��,�RF��d��b��
��p'��
<��,��3�T �t���n�������q7*�V���Nڕ[��#�����u�G������N�c!�ϕhڟeV�4Oz�2ݿL��Ȭ.�(Ӫ������R��
dl��C���yVCRk����c��8�'�� �������)��d2�h!~�6����{i7xJJ������	E<so]H��Q��z�&f����L���.޼)#y�U��jOd�h��+CR��$\�w �+��L?q �>�p�d�d�ʬ��k���S��̦/x��^'�a��~Z�EŮ[|Ue��?��Z*�a����A�G��$Nm�*`ڴ/kD�$�BX�s�`)m�&��-F�?�55>�ڡ�6�<����8 �:B�����Y��^�2gB&�zK��چ�ڌ\1��%�ML\���-��C��r�q]
�*	�K-:�����F5�춯�&/�o�K���L�����s*q^ld'�s����ױ���{��p��jr�P�锊��@V�{2B�I�pcuhͿXO�H������v��vz�S�� �~���@���B��Dۇ�����.$g��X��S��ᝎb�R�8&��i��:P�;�#dW!L���T&Fџv-�I�M
�Y��	�SŮ��SU-+M�y�`?V^��	���q���u����y1.z*.7�MiP�; &p�˰�Ά�S\}t���dB8�xG���ɂN����vy;��.vj5<ׂR'v�sn�"nk��]D+&9L�}��_�#B>bw�%�a�����J9��T�Δs��,�����B=�|��CHSp�4�*�;d�|0,ߋԯ	<�(c6eu=���$'��%:������C�g�l]�iy��bS�Gͯ� m/�M��, �4&`��ŘJ�������Q��63�yQd	��Rn)��#5*:C��	����0�mo)�X���c+(uk����n̸^+��o�;���'�v�<Ms��k
X�$�ͼ0�jP���'˶�Umw-���^_�6�.�`G�,�E�:f���X�}i;K+= A}߷�	�>�Ic�>�s��Ò^d|����*哘r�\�e���/���ؑ.pV��n=u�m�����>�o������=��N'���4XJ�L�q�$:�p9żVύ��'�(��D��f���%�}� �ti�G��{�E��p�H6/�_C��?g�i���嵃�o���=h����O�;���,�-�8���΁ ��Rv��M���N�G}!D�=��,���mԮ�����˧�o0B'n6$�:����$ 
##�q�ĩ��.>�crDpv�݅����L�\���Z��z�G,����M'�zy��"�i�ӆ��]�&�ȯ�.��&dE�(W3r������ͰSھ�9m����A�֘�r�f�?��E'��V���Ą��$��"�]ǌ=)r���wa�郁�eQ6��8��t'3w�ߜ�bs2�9�>