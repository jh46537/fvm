��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb&�L�S��O������}�N���A���v���sF�؏/;�uFܸC��V��+��N��[0��5s�a���v����1�Q�$��n4&ͽb�MD��r\���F��E���5?/�Tr��o0��Fn��/+�V����>�z�����*!-��������3�ˤ�F���.�[.f),���5g��k�6�i����+�K�cϭ~&���؏���5n#�h��߽�$F�m5���<��{)�r���j]ۗ����O[N��I +=&m ��E}C�����d�2g���edq�Lh�A�B��J�F��=у���Ü�vak��w����9:0�h?G���~�+�ATs�=�+��M��P{ ��Y-U�3U@`a��8 ^J�����^@3��ė+��Sjv����sJs)lf8�sU#�Ȳ��3�w�L�P��1NN��^6�ڟ}_{Ie8�������/�q����m������=�`��̣V��u1߹"��C�bU���3#?��`�RW
�
�'�8�������rj���S���m�,m��H��k��?I*�y�҄�>-Μ��C�KW2]��^���O1#U�	i��c���!ӵx�#{
��h�G!��O��Y�He������� a�db�4ea@\��8=�듯�Вq�"�� �2#V�d�5&ۚ3��W<�Lx�4n]^+��Gn�S
F���L�w%͗��{��;�x�`�ů�T+u*!ԈV�'(5��g���9�2 ǝFHw�J��Mzҩ�����S�M����M]�3>�(���"Ifc髵��3�͹������y%I������-zPGd�ӻ���&\6���뻹9#Q�e�����L~Ҕ�5����'|�M��#�%�=�3�/�Â��1J|�,t�8����t�1��◖5�����)�k���Mu��dO���,�/aQ�i,a!;eu�k�?t�Y?U����5���9;tC�
��>hSg���t�B��E�j]�Xz^l�ipV������e3�*���U�`ճזCqW܄k+�՞;��v�I��&/�5��Ϛ�
��ԉ��H�S��"մ�z�6_= ��vc̛��z�*<�*�$r��@���A��U���3][~G>��2����������92�˔HN]��΃Y��h��n=r@P�Qu�,�fON�L��2���_��'�/����:]@`z8�<����:����o�?a���'xzß�8HI������*�s	8}��R�3F�1�`CNCգ,-'��ۂjz~���J��,K�S�m+?�]�c�����Az��F[��TnQ�le萏�mW������!{�{O<z[�4�A�	F*Ԁf{B����z�-� �2��"Y7��+9�\�.l�S�M��|�c� ge U�\7΀#بeyU��
��	1*:V�3�"ǰ�.�^bH���n��q�lhWϒ��"��b�`r�C5��>0
F1%!ۊR;��+� ��3#ī�/��t��%�Zh��m�I�����A�iTgJ���h<"�b�EN�+w6M}Y��4W%ԣ�`�)�X�i��bU3�z���ea�k���M��ϖ�J����/��6�c����i�1�[�È.9�]*W�cT�~��3�D�!t�U�t������'&Y�d�;��s;y�����<�v�<�x#��:��j��6Ѫ�eJn���h��z`!�����$�>