��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�X)�='�L�.|�w1�ށͧi���캆(��	�q�8���Y���X"*�(�ܜ�R��(�{a�������aW��	��3&�b�OV��_�Ej[飅)���X�t"Y�8A��g�:��]?>��yle'=g�n�c�~�|����a��ũ>:#�F�~�hj��!���/K��a�`r��]�}|Q�Y��[����;ku�ԝ���!�o�P�P2o�U��=�N�5ogbF�9\I�M]�ÌhMۂ�m�Y�A�^�,�Nx��<�W#�9��G��2��x���9��Ȃ1��\��C�A��3��gX�f���qbU^��C����=,Z�l��{�{=WJYc?��A��5��ۊч�[�̐ESS'�5��d��:%���p%�~AS�~9���je0s;w"�>�_���7]2�Y���6�2�#4�/��K
tg�� ��~�d��
�'���8�MҸ�7��{K�m<���{���h��V+��3q�a�q%!ޣ��̀za�~��!W?���|�	�͊j��x�"��9G2���3�e^������'5F��~E�W��w�9P�9V� ���먡&�/T�6�q7qƵ�;(w`��
��QO�m*��8���A��[�Ee�?����Z��*
S�y���ʥ1�J�-��-�	1�`x�A~�D~X�zD��H�[����Ţ��.��i��Hw��,��<#�AS��I~�R�����"�������A����,�I)����b��vk�dS�����t�6i�����k�J�w��աHȖ�ϗ�y�V3���ņ�š���̬�*<��Ә�[��u�D��=e4ٜ_0mV՚�ZR^lUn��=vw��U<���䨚|�x�t��_;we
���X	�Ӗ�0N=���Q�{�7b^J'��˫��C	���� �ALybT���4���I�[0������@[|�����Y�`h�)P����>�����i��~���&�����|�x�9h�Ϸ�%���U��r^:9-�W��1��YqGŅ�o:S�E#ʝ����RDW� �ɉ;z���K�C�L��X�=Ng�H�R�U3��6|(���/�J С��NQ�Cz�C��%/6t��B��� �`p%�4P�V|�O�E�ێ߯�vc	�Vʹs��k-�O��Ũۥt#���0�����_Jޣm:t��%��f��r
���xc7�"���!}����qG�=��E�(�=����b`��$x%�H<"�Ә�0����)��7-�W�d"1��'�Yk�D'�!]��;���W�����+ê�e��f|��N��$9��7c����`��E�|tx<r' �>��;[����k�Z쮩��/����Ζ�s��+R$+�� ���Q<#�����&�^�m�o�~&5�ӏ�;�RT�&��󐁢��G�4�.�!��ߜAyAs�z��N��8�i���06d�D�=��0��	��}m}A��dN��w���O���7���\�Z�3vZ�=���F��i��������^��D�lR���x�����2��V�K^>��cO��<�`;�̱К���&=������1�yW"n�?$����ʔZԞ��T
)��Y�f�R0�uue�=7��嶣���# M�d0�tF���vi%��4��U�>�����&F��+�F�bN�D3nG1�"�%�k[F� h�u�Qƃ@Zy��M��aƐ�v���.}������@����wY���"��[����O��g.�,;R��)���)TcZ��
��X��|G#����H��5E�ݪ@��
ܪ�[�	6���9�
�j�U�p�3�Z���@E�B�N����3�87Im���9�6}X�i0#�]�}� ��wŔ?��6�W3�/X`�.q;��:/!X�x�y����(:o8 Dͮb���!��H?���cA�M�aɔ�f��ސ�ӽq�~��a��?�u���zd�m�F�`'Y�<6���[Mn�)sz]6�?��@V�G�|�c �3��x(��<��)�׬]��J�PT�)ک�ee4�9��q$3O38XIWdb�S�eR���S+𜆲��W�(<7]u�M�Գ&��8̒���2-9�R)�x��:��q/�jT��-	']>��J�q$:۪��J�`i/����p��ˉ<�<�[B0ls�9���^�a�ec���
G}q�<�cd�S���C��,w��V�|����Ӫ����}�k:i4{�����D�$��h<4�gVYVڵ7��.<~(L��0[Li�±x�s�b�{�f�PVz�ȇ,q������_����Dz��	v�	�5Ľ�E�2<��Y���Ds���N0C`ZQ)�r�a펐j_v�5�����)��Y����cޒ7��(��|���6C���w� ����;�jN�����ylR;5��+·g2�?)��0�B%-(j޹E9����ɖ��ö�.��<��}($�Oj���i6zM�c�۫���k[����4}\?����X��Gs^�=t_�[ȷ��営'��d��ѷ��O�ݫ�ߧі@���yn�^��'9������?4�
?�/�h
e�+N%h�9p]!D�^My&��Y�tԭD��}$�K�L�z1����F����Z ��>	�)R	����hwk|���-��¦9#�,Q�4�_�A�%z��Ti۰��ea`�8P��(�{�V@=FH��k??����Fc�H