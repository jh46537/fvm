��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���a�%�sK��h���/a�y���v��=��w�����:�y$f�*,�RA\��S����ћW;�U���T�Ǔ�q�0`�eѓ^����8YU?to�Pb�I�����9���������:����l	�~�Y���)���L8�|m[P��Z�ј�79Ӄ���e<���_�����^�2�����
v��;�{a�<Vx3�-�����ٍ��/�[�mg������o2����@�m�e�?ኂ��l:g(Ozl8S
�-�CW�gF�5�դ����>��'K�:���ϵA��8�l��X�0S����b&�7�%)����!�h/Sq�㾴.��"��w[�Xe2�.ƿm�?�g0ۉ.�*9D��>[ˬ�?]#��m�g+��;��Lb�W%��"�����n�F�`��VW��th��Y*�1 ��a�|�!D�+�iN�>~ރ��r�E/0C*�ၴ�ҋL�����{�ӷ�[�<E���˕4� �T�Zڝ5m�g.^kbHz��v�pZ�<i��9�� �F�g`�X�ӂCCG��t�L�ɬ��f��2q�
X7Gqa#k��H)��"PU=D� X䊵�C�C�+��a1FR�MlL���kA����P-I�נ`��j�"X��o�Mu.�y�nkQ��;�⬲���K��ի��1���p��\���/�a����]��T�K�~�x��q.�)[��d�����m��`��ϐ; ����V%����OŲ�FS6��*UZ}�������ăK�I맏s�4u�>���ЎK�7���"X�����s���0p��q���<����}v"�]6q���v�I��?�\�v�a'�q�����:),��"V�,r*�-�.�(����f�<���$��)�K{�3)'("*�ɪ�t�҆
Y&�s8��'�������P�9�1�~�)v�:�"M�B�93�(.O�|��I�Rh�\��O�\Uٜ��~�&�o�6�=n�����T��W��v?�Y���\�ФD0�S��Eff�2��k�(-�� Y��[=��{>8�2d)_�Td�����L�t�?�d?9����t����+k��`>+z�l��K� ���������aV���m'<�@eO,�iL��n��D��QLꪂH�O蔿�&��U@}�;
�Fm*��ᐎ'�MS����-�C5`j�������q�|�R>Bn%��+&��Y�+uw7s���V֍zC^�t����	�ۨ:���?q?���k�-�D�/.C���V��qig
{�MχG�����:���i���)��`W�6�B``���+K�B��6j���}ZW�t���q�g�0�;,q-+5�4d��p�#2�q�u��I�}ET��bQ�RL�*�
��z�+}eRd�|l������t��g{/��$(�X�|���lb0��W?�Y��tԦ�.l�\�L���:ޡ ����f6�{H2-N5��eH����5޷,=��2�B�y�H�R�_���Z]:)/�������YR}xY�#=ݿ�C��b%+oÃ}s�"����WB�A��v/2��.��ߋ��y�t�*	^^K-:����GM�����Ko8i塰z���^HYvU#����'w��8�wT��S�s���6V^O��h�7V}	��v�v�|�/��YU�7���;�F�9�Va��'�űo�H�	�@�h��c�].�YwsWE���K��/�;���񉕘���G-�ٝ¬�!���e�t�]	�����Ѭ�ml�$_{�'�H�
.)�� k��J!���Y.ʼ��qm�/��P�k���e���S�ΨKV3Q5ox���t��E�*��Ų�}��zi_��ţ@%���\���Z
�Ð��
A��������g`�ᮨc��f`��¾�
�6 1�F��*��TI�e�\ǣ$;�H=��!���B���#2���h����o� �q��s�%A~z����"�)��,μ��lsG�+�j����#yJP]��R�j���ьk���I������=~/ySg�Z�mti�
C�}��Y��6�q\��%��ƪ����~8��6vy����LE��/�?��!�h������d]@L'I��l��<bT� &��?S8�1����u����i(��i���*5Y�|���@ �5�1C�C����ڸ�?d`��b?��S�Q��d����m�7U���%����f�<��zZ����ƛR�ޢ�@������y�o�r��5�(�cR;���s��aq�H�;{]�FG�H�f�/��DЙp��!&f�R�y��m�>[)�t㯵~) ��mہ]�M5D�����x�O��h�ӬֲM���Ω���mus;޼����ᛣ�E��3ɫ)=XRFY�C��jg�{�gl��G�"��F�ߛ��w�(��V��vO�}Y��oDx2&�sV�$O��r�-�w:��WC���b~�oX9�+W%�ܷ@���x�� �@k�-�����3rT����"�Kwqx?!��\O֔ӵ�d Ta�DGH�4O>��pt�i�i�1�}I�Iu�=f������X��w?���;��f;�"����&Z���N�:7��M�KED�lɤƸRu��.4�(u�ɇ�O���o)a��	�hV��Yj<�N"-�V±\w�'�s�����S�Ɵ�\�X�
�{��?�I�5Qg���xmv~@�,^��B�*.{GH�)BM9x�1�g"���0&�4RN��?ﾧ�adl��p�̤���5���
Q���A� w��0��$V_N��"Qk]%��}��پ�q1�t3�y��A'�
kV����r��\2�O:¦h!�|]s�����P�r����F_E�Ue�e�;��������D��J�>�4j��&�j�/��)	�*�ͯ�7�¾O"��I�3z��I�V��B�A?�F�)��OEц���i�f�{��8s����@-�Yq��75 ��!�8u+�:��HU�Z�-��C5�Z��k�sꊏ��L�H���������θ����TB`��6�|��/衱���\y�8�@GWv���t�:0�AC+.H,F��ג����g."c\l{|��~��>�ŕMN�k�R�����^��f`��F񱂀�cU=��F�����m*������rr�ۍư/��u�C)���`z:���jZ��2�!B�S
$��p�*U����zF��Ue���ldNGiNض�m����K�Ѫ$<?��՝R@j�����d1�"VE��;N,�{M;.�Gy��U0�����)T����LFV���V��~�V���.��ܘJ�ψ2�����`�J��%��������qZh`{�����"�U���P��
ZW�/XIX�E7�Q����h�,y4E�zOH�f�4kW��V�n���k�������b�8��E��)y<.๕?�uě��KM~�P��%]�l���'�w���_��¯NO��d U��:�9 XG�	w���\I��_eѡ���>�����]�r@V6�@�a�(���(3����7VJ�S������̈́_*	
�h,}ۇ��$<�lY�=��ɩ����w����C����p׏�Z���?�����!��WjZ�u-�[p��uL���>N�>���z�o�8�6����$�r��ȝ��L���c��Q��W�Sq�h��,s�F#H��@�̯�HYq���H\r9��޺�0yC�P
4p�:�t�}N�d:7<�ե�Y�e�	��
��D�p�^O�qC�g~�hQ3_	�3յp�!F#h�{�@f�H�q1�����WĔ�,�d^ ���Ji��Qe��z����X��}M��|kL�� m�w9����F$`'"���l�;�+�[f]���#��j$��~�V��Ҩ�.me��_A�IK�" ���2ԩ���0��2�怛[�0h���X��M�/�3�Y}4l`.����ih+�,���u�=����� �،����@F�8�1Et����1u�j��y+�`����� �����xv���̙r\��r�P�y��o���JG�	ֹuYOq�u8��s�?�	�[@V\��0[]zQ�s����j�_P s�n�tOR�'���#-��q�	C@�,=�͵A<������|��(����8DYp!���?U7A<��07���2�� ���)��T��U����&-�<��u
��)�,�0�ɧB��c��A������W�\�Z�7R|��z���>^�_��N�d���;ie��R��io΀�����@I3H�
l�ѷ]I��-h�sI~�(=\�E���Ý��M�F�X� a�t�W�]��_�������>�����w��'�a�Dم��!���;�װ�n	�����vxxz=d@bS���H���	�	�M�1,΅��]>���x�iڬJ&6]�t(;e՟�+�Ȁ�LP?7������w�ߟ�|���ӆ]�zq�?t׊�*WF{,�����+�����ffn,�̱��g^��K��a�����A�P`&��@�c�ú&$�B�jrFd��L�����0=<�C�sپ`3��6ؗ�un�z��{1��ͬ<�l��f]�b�{�[Y�ˏR.7�
'�k��T����k{��sP�bh�I�ENj��3����G��]h!N|���MqEN3`�	ϛ*���w�7U��V�d� �CJM!�C���f��"�o���V6zj�'��k��L�Zj����� W��P������\a��C/'�VZi� ߬��ٻ 8"��,#������0b�Pц�p/~��6]�W�y%ś�0�4���N@��@��;��l�]�p�R�I��#q�N��x��f��쯡�q�߉��J�t�~ה�͍	�=I��B��I,}zg�XA�77n�^�������#�� ��d��DSO���`��%�=��3�R��n������$��h�[v*B&�?�DLs�8��B@µMt�Pt�HZ�A�q�g Z&zg��9��X��M�c[��R2�~=0�������vR�E3W2�k�K�J���7,Lis��B�%�Ȓ�%��ښj��u�d������US`'	6�R���a�_mQ��wW���$��3��� l7�1c����V��[�|nq�,��ZtҢ��4W!��k����	��Dބ6 ޠ�I�[Zwt�u��:l��,�Ę�8;F��y��Xu4q��>�S3�<��ȼ�/��xWf7t9�����eǑ��߄{�E�.�&��Sb�&��3,�fa\>�RFe"ֶۓ��*
{~��r<r l�����⤠'�N�ݍP#�fo{rs���m����s^���FC�D�6�\BJ�;�ڱN<ѕ���j��z\@�|�T�����es(�P{Ҫ�,�\�!�˦��D��ZI��fn
 (�}>m�� ���[�ݜ9dی��w@��k˃{�	��>���2�f����9�n����ݧ&�;V-[��-����Z����ͳ"�.&J�;=�x7�z�>�_J�������ļ�����9���� (�-�,|�Z!"_��ۯiS���dH�<���*���*!�I>���W�KT"��W膝�+��ӯ�g��\�%.��cN��\�D��k�ȵ�7V���9z�Ơ��P���p�ͻ��i��T<�[�Y��1
f+�:���-i�N��rg��G�
_�[A;�)�)@&t"��9��L�fFg�א]���p�4�� �o��{���.�Q����0���%����w�Hү��8��(a*�S{ �K�Ex@\�mP����x�\7^�a����f���Җ�[Sʨ�a�T�( �����G!Hʽ�R�{[K}��4�91�`x7�3�|.�{���]��%�WIk�B,u���Tc�Z��7�����đ;�� �Y쑫>�@���� �.��8N���XU���֠��v�C� �/�kO���]s��L�M����HS�!	���<,�1�D���J�,��X������ʨ�Vy�ȍ�5����ZnG�2p�IOM�a�D� �� [X���Y�îA�c�ʄ�k�{���9aE�� ��	�%í��d	�C�Č+J��so�Y2υhy�y��k�e��0��E�":�q�.tvd*��{P
��U����C��.����58*NY�n�z�t �A̩Ѥ��pb7�a���,����(��ǖ	�üM��e~�.�����ۈ>Ƈ�33��?M�C[��o��ؐ0߅\
�V������iI_A}Z�������E������Jo!O�Bԍ�@��fȩyr��1�'U�юYHT~Jhd�� 7��Ea��j��aO��Ю9g�A�pjx�,�q��#�CՎU�q:ۦ%�F*���h������ B�L2���4�4�
��J3�ȫx>���A���ȩ4�
�%��G�	���.˼�V����P����P������l��A��M.��yu�s���A���W's\�^۠�&�݅�|����l\��%��5�>�ReXc�t.:������j�L�B�q��~�mG?Hţo]�e�Ee��L��/�`���I�7�]m}ԥ���Z^IK�?�ORBz�g��_�K��hirÆ	�N��;��k�|�|G��5�%�U�D�5�0%x���s�r�t�Q�qO]��Jk��ŒЮ�0�7"p�F�[��9_��������r�X'�*���H���!��Ĩ'��,�N�cq��GZ�C�rl�Z5�:}-Il�m�21`jg@��ǟ)a���z4&�ƛ��
��dn� ��k"���]$42� ���3��*�ܣ�P�*�H�0%��8���5w�����X; $:�R_Bݢ�1DN�EˑlUy�$�ec�iB\�.�����d&XP�=Ss-�e��]�?r��ȗ���Z<&�4�̵���&��<��)�4��:������^<ڙĮ�"���ü��eD6̩DG�j��Tw=����E�.?�"]�?9���U����_�?č������z�ɂ�JJ�>��yx}B���E*C��	��8������͹��8g����K�0���=��V�Eƈ^V]���kUfs<��5��c����ت-���E��1p�C;��)a����Fn��].6eY����K^@I=eY��6y�>�X0e�ַG��|������&M�$dZ��βQw�;~�ڞ;�P���l��Ĥ� �!RgM�Eg�H�1�Q�	��˻2	V��k����k�=��6��L%U/�w�P�^�V�<��ASƐ��w��t����`Řn�M��xk�Z�g)l�o�����Pmտ_�����Yb���]w~�:r�{�(��A�	}��?�9E���T��?8/ݭZ��S�\�nn���bP߱�l�M�p�� CT�Uz.���p�-�lL������x@�+�KC�=�y��j���a]S;<&d�}�i��"L�.M�'��+�u�gxA@mdq�A_��� STa:"bJhb�)�YԤk����6k�X�"�F���{�S��gHs�Q��!bD��P\����%Z�M� =_����9a�][�<&�������[j,p��k'?�nz�<G�dah9�3�Y|/^�tuȤ6��2�蟮���L�q���P5�L�~�cd�����b�3- F�=�H�v�&jᜂqIT>���*Zc�,�:�x�*�^�}�`�O�.�z�}(w���Fd�fуJ��/b����Cg�O>�J-B�V�(�m��Ă�������b`8��.I:�X�����B�#��̹A�����(�[�rkiu"AC����d��p�����­T���+b /(r@��!�v|ȉ��D|v�	υ�dG;g$'�h�A���~U��W�!E��<����P/���"'�p� �g>��g]&R���;�*�!����&F�B�	�u��k4j�O�j\i
��$�)�O�S3"�4��l�ϋ�O-��ҏ{�#�O7p�Pt*���<jM"2��X9������>�T;`$㗌"a?�8��?���Ą�I�+9��`�&�uJn�3º� ��$���nBբ��K�2���r�N#L	���r	򎰦�:2T:
y�g�>�7�#e�ٯ���ߒ#�ZLG�xщ���(�_� �����ht"�̗PO�/�~@mJ�]x�������XX�!�� QU�#�;����C�m��8�"TDAb��@�� ���ѭ�C�B�7�!�Ġ Ǣ���#�{=�\+���K�~DT�0����6��&�/�m`�/�L�p�Ȫ�n2ܲD�Ʀ
�۾[� B�w���)Ke$k	��l��ඳbv�J��;Lm�s]�i]��lPf�o�Qp�K�܋2Gz��Rt��J�, bR�W4*P��2:����&a\s6
������;N�~4������S��#�{)R�X suw��e|X@+�>���A1:��~���eb��Z�"�V!v"<n��gm���Ș�%N�Dl�M�P$�KF����F6��)�d�(�'��]�WP<Nf���ų)an��'�T$�;_�r�љ���F:�O6*A�MM�����뜹H���dIi�e����Dc���3r#�< c���"����6�'>��~qλX2/Ez��)�RK�C���Fx�"#��V:%���hd��':!�������r������0����s�_N��z~2r�:�yo�g��,�?���J��o%�l���>�H�l��S3�~�X�[���)���p����a�7�!e����pq'��D���GF@��+W8�9xPT	���5����6�(�w���&)�]v��L\���}e-?���%)v<l�I����׹RKI�ŉaaٍ��P�0��q9 ����ܑ��h����)m�i�g,��b�S7Ϟ��/y s���Rt����U���y^�i�*nr�B�{Ϧd�tƝ��d�9�ș&��C��0��/�lX����`��a�n#�<u9�҇[��Ei�3Ŧ|��؏�J�>K��ж���K@�N6�H��MI-���Ksm�$XtSٮwS�B�ɩ¯��L��^�/�����~��,ߗÒ���$�i�Q��o�*�YhQF,�c9� ��T��8ϕ����7=�Rb~������/w-L�O�w��9s~N4ɲ�Ρ����a��z��5iٓGb�5�q�BS��k8F��f��u�<��[~��>��E�e�t�;�8�p��wE��#�����s�����g^�%"���힂�0�Ƀ�k�L��F���CD������F�տ���_���ꦕ_�(��f������=��lr�:$:�|�酞�s>���z�h������;&G8��,^�D��]���T��1�W��� ���c¹�[֘De��{D<�kp�B�Nŏ���B�t@rs�}`��"9�.%RĦ%�;v�6�08���E� �B���� ^���W�<X@���el�_?�_ڂ��̦D*5dGp���X@M>/G4ԉ���+^%F$��LI.ʧ�mD��blz\`�R+n�k˞Y�U�ѨD4�A&�o�ex��*s�?f�0@��"m3"�0�����=��ߣZ��hB- xP~c"��՗	z���*UJ�f��ŏ+����� �$��.E���]�sr:QV�/��.�N&E��/ҁ��&�l�O�c	�@ц�ݚx�``��<�b�����J�������Z�]V����=E:���x�P]<��O5t)�5���˻o��"�8���a\��c)`��] �Xӿ�
G���P91)ZՁ�&2=�a�Ǽ6���>����T�x���T�-����X��ٗ_�C�0��[<��z�G���P ף���$Ӎ`��l�
�̴QS��1�pTf�V�"�h��
�$�2R�>t�`4xU�3�}�����rVz��L�z�(��/)�n��EdJ�G�I�ބ�t�@�J?���g�/.�ݐ���X���g�/���Ц\�U��Z���2O��7.��9l�Z�ʀ�0itSе�zR9O�'WA��O��I皠���*f��_��A��MT~��U�u"gj�/��Wu+:�BzM,�Sii,3;�-O�"g|A����*��=E�s��*M�R��fq��8g�%��Y�<�j?��~OA�%�-"�Ш�T������(6�g����	��(�l�"���Q,O��lE��/�--N�Fg����ݗL��Bh�TR��bp.#{$EM	�xƀ��J��2� �u��V�Y�����e��ad4��s_���R��&b�t�w��GEj^5(���=��լ��X���"PW�UL�";���@\�"�U�Q���Đ�[ףɄS)�������.
7��9m�,� /�X$w����G��"f=Z[����S�oag�y�°oN� �3z�	Q��\�R��s�`4����m��y�L�M��ںT��\R�[�p�35�{(�PU���z7�XwUə'�S[��LG�c�}�M���by��,+�~mS���_O|��}k��s>2?�?�Ky��k*v�|7n8*qVH! 5��<��To�"q�`dck���Po������*Lv�Z�)�̰�O�ik�@�B�b����r`�>51h훸1�fl�����%�2x��#��ZK��5�\��m�"xW���9�e�/��eq�"���(>�P�iI����QU&Мը�M�i����`�AR���TnH{|l޲� ��{�LD�Z���o� ��5 A��D���k���v��bvA?_Jz����xӑ'�\�W�0�����$MA�ߵ�e{Y�j��_Wx��,��1%)��K�;a��v�����E�cČk�S&�	���h�~��0P�;2������ƬN��t~�-�g��ƽqW���E���yEҬ`d�~����?f��Ѩ$�E��gM����Z�8�����B��Z5r�y2���G�u"�LP������Ff�Gk>����E0E�[mú9&D�����AQ�(�XGFU0ld#�Ե1;��E���p
!d�1V�oQ�̵$�˛�(��R�~X��f�Ӝ�1�6�kc�,�Q�c�@��3cy��H�
���ls�˲�����T �Y�/�D~l���!
KThm�8��\w�������S�<�R�^m��cP��"����i�����HX�^�zP"�����B���-���_�ռ�e�P�9�.�7��9-��He�D����b�p����˭=��<�����I+���H��p�铫o���E
�̳y.�f9�����`�۰j�ɸM���[켣"��u`�%5��Ű���7:-�c)��F��� A�uz9Ϊ色�6 >���j/��:��סkh�Y�NBJq?�{d�<�LC��d�Y��9�Ee���[�V��1-�{�V]���-�/���nZ:���<be�Q��T�,`PXB%c��'�K��?&�^U�m����`"۩�O' i��VI�=.c���ۓ8��>�#o��I.Vw���f�dZ�[�^��Ba�hŧW�qM>�����)iF��e���e�i1�Nʩ�o�Ӓ�D���M�8�gI �Ư�+Illx6�*t.��4�-�ӗ�=��z���&n�@�&z]iA�b"������W�"�</}�}��@!^����0-��J(��iG�����.�b�����'�Ҩ�S<fz;�5m���o��t��QI���(a��4���g��eZv�0�A�k�yCO�{>n�L"]�����G	���8�V(L�o�{�3��(u5�ŀB��봉&�x��sNܷvTK����l=�@�|�1$���tb���~������ ����ױ�� ���}ʰc0VN� Q�H'��_���'U��E�e� �����K��ۆ��=B���NJ83�Ղ�E����z��1k!*�8x  �|�㉰��ƙϿ�B9�731�� �^"Tx�UN9{؈.����uHB��:�3E�b�׺wDb�9i�wM&�LՖ1k��)=�ha��ru$Zi5��Q��v�F�g�J�RZ�����As��p��=�s|���b�e��rj�c1�[,t��������s����%HK�Gu!d���<�3�p(k��=F�//�