��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}���j �]�ȴS�����a <���v�D���YFJ�0w�Aq�'���ɫ�o���s��Ϭ�K��/�)���o����{l���yل�Nh��M�����j������m�%k�=t)�Z�T:�/�9�bM�U\Q�)�$zAS%)i�8��>8�U'Us<t���9D��޴@��Z&��9�d��q�˯����G��w��~�G���J�����'�>�Z��U��J�����Ő5�����/���G'!cvv^����!��>���q�U�L�O1��'},,��sf
�	͟5d�X6Zx�n0�d�`=�m���!�	Rnq�̋�NB�v׹����Z.I�r ��>��1se�v"b0��,wI��!Giwb ��<WW�:��	>U�"�^��1)�}t_��H�[���,e��Y�6fw��Q �=�9cg��JǱ��9�
[��g������/���ɺ�:aw���Jr{`Bm)`�k�}*5��"�!�PRR�i���Xz�Y�/���?mɀ�|^�[�>��{)��6?��S&ǌ;�hy(�[�J�����w3���]������u��^���Xgidh2!��K�������^.���ků�TL����!T���:Μ�l��<��C�y��C��=̔c�zB� "�'1u"Ⓥ��X�t�js�ZD�:���/W���N��:#��8�-{���a��#h{���j�p�F��4.G��'Q���X[~�	L�)�On�&�X�iX�b9O����ь��8���z.���-/��	D0@���Ho#��ي��r�#�"��!8�Լ�99�4L�{�˝���3�>�^p�	 Lkg�q���R�˰Deʷ10��"7r�;�c}��u��9j�q�ͨ0�D=`�@�|���A����!���xvgV3�ꃎ���՗
P흐�mʪG �a��j�W��K\|��pN0�>d�6�gN�Q���_�m.����OA���:�YЫ���d�^����oybz��-؄��_��V��M�]<�O�1���
�p�m���J�(��sj$|��X�H2�z}��j-:�b{�1J�05�i�pg�.�O�'h��3� y`7S/Ը?��xɠ������M�'����O�׍�t �&Ʌ�&"[o��lW�./0�� 8�2��(�j~c��$c����1��C��8�o��^p5��L���q#Q�?j�s�)<�ia3�9õ�4;���P���@�L�>��K_���Y��+&SwOd~�7�=��d��۩t<�v��|��Օ�\�����bh�F�ٹ�a�m�M�:+;��3��:��gz�xdf{1���)���It&y3N+4A'�m�DG��OZȚEM�\X��bF�� !s���C�EҠT<>����ϣ�0^��u�����f�9=�u;�ܩo��y�s���J.r4���k����A��� N��l����Q-k�j�b֯�޹eX��
 (NB�O�dl} ��#��<�5]:L���S�{7zzU�;���w㬖㤟}�&�k�iR�-�)��?vr�s��. ��5T����,ӿ*,h	l3��V1a����Z^Ǧ�
M@�O�����o��z��#�g�(;\�N�ծ�c����Th<q�M��E+(@�(F��Zު��N�v5v��~>e�U�s�;�|��\}wMl��x��<7nH����ɧ�{���k�(<�x�m�gЁ)��ǻ���<���ZY�8$���j���7�5�a���cx�y���YNN�&2��;�C��͘"�[h����
��*Iz���J̴h��T�d:	��W�*�vԦ�{G`��-��Ř:��C�m�Q	�-�ҳjk��K�a:�F����dv���!|o��1�0 �"Y��-���+��r�6o����$a�h[J#�P�
ggKI%
L4���D��Mk�6�C���U2H)ϋf-r�t쉍P��DIjv����Sy��⁊ݑ�nq����xe]!�N�}#JBl?��'�}�����p�'f�u�/�
�H&j�Ւ��
��;}�ㆽ�ߚ�;��KOŗ���17���h�v2y$N�SS��A�k��.�y[��Bf�䏋�h�θ���� |>���f�����cj��H��0/*?�?��=��t좫�=j9V'4��}MBP�"M�4�
�cD���|	���� w��9�P�Ԙ��5� ��`Y����12�;7�0��=��Ջ�fԅ[���]��a8�Ȋ�ۍu#�o"�>:��:�t�W�NP A�VW���I�^�*@|�j^vd�y�~��)]�Zmؽ��5�kY�q�����Qg�U��i��z�1v�0�����1e���m��@�!B�_����(�#*2�,>���.�Z�`��]U�.u�S�lvҋz����!g��݊�C�����i��_�%����ӌ����@,:'��	��'<�A���_=��L�|�Ɲr.Ws��L�p�t,&{dH�wlb�n&�q[�Wj�����73ӕ�}0s/��n��һ	qͳB�/uɛH3-"؇�ofV�f�j�� ]�j��畣^]b��{!�pO�s���TEފA�xh+��/q/�L���i�r���W�
�燴����:�=E
�m��C�ҿr�a��
&�4�:I�7{.��2+�xH��TC<x� ��'��M�q8N��+��;�6�@8D�O�lš���`���+p������dh~G�_}.r�$��C3C�n{'�WEd
�,t�?��8O`Ƞ:+��W��x� M�d�C�}��zĪ@�cYJ �y�%���|�:�+f~b}�.��(��>E�Db�i�����.p��ä_]�:	xP}@6
bw�g/c��V;;��g���/%$e�LjH����p�
�*�W��ۀo��Cm����)t���e���x�1s�NM��,���鹑��kkj��y1�	~�Ho`�t�w i{6xU��J�jD~����zb����!�\ܨ���ER������p�a��Э�zw:�~���2X w����I<t �iހ�y��p��h��H�W ����-��h~�(���EC���ѥp�GW�TN�\��j;�4��������h�|4�?߉����,k��d�V�A��0ݷ#�ݰ��$��ޙ��ͦ�wĆu/�2w�-O�� ����>B���3fg8�����E�7���3�)G�7�
��Ȳ�%S�3_��+-��Y�!�}-a�n1;9w��u ^�W-Zn�̟�.�K���HH��\g�Dk�:Zn�0"�x7ER��6��1z�Nu,�c�h��:�~y�M�����H��*��;m(?_�����IXO�wX����gD"�F���v;Q�m4������zQ�X,~��w|D�E�݃$�[.���+/u>��!��de&���q�d�}�g��2���Be�C�s6:d/Ӄ��StO��. ��I�����OP�){��lV��$4�3��"@k�r�)�:)T�,�� vj����֎�/�-�/�����7jX�dE<���:�&���]X��J��O�-����
,&��[V�_:
A�(�#����L~Z��0�$� 3��b+]���l�ıw����6��2Hwy�u���`�/�!}'K��X�R�p*K�cCU�+��|LT[D��T�52s|2D�n�Y�򊄈���Zf�S3#���+Y�����P]��K ��P��QX��L���|����>FeL���2�\���	����x��M��j���՛`��?߷V����׋Pg��d�d�/<��h�ƃJl��.������ֿ!��!���^)o��7)?u�3>x�*Ǧ8(���p"���N�?����s�7'^:��!�پ��������2V��?]T�$^�S���aQ�f7�<��C�Q�d�tςn�o�����xL������-0�G;-�����T�iY8���EFo/܅�1��	eU+Ɍa�myq������'�C�eh�������e�D���`�δL�\It��5���b{�`�2�����M0�f�� ���;3���w.��qʓhŁXk�z�q�֧�w����q8��{�L�r�"W�v�����('��zw�56�#q������f>i�ih�'�s=C�3�TH�gS�d	������dd#�o�^�m;��cO�՟��s�վ��c$6?	���v�;��D�%�V�?�n�<���I�9w!1>ֱY��~�����6Kd�舢�s4� M���cL���0���X�&z��]��*�V6��G�c�R|1�i���S�G��φ��Hn�h(����Ue�dv�D��	���\3����r:��]��������og��㬞������+,q��;��l��9`�~�}{����TA��}C<`��5l�*8E���t`�2C���G���:)���rn���{3�/O�ت���M�a�Xvǰ�ʲὅ��b(��\��F?�j�0����5.�
��W����3]�D�ԚTKѯ��~J�p�o?
6�ɦ#'��S�5}�q;eiO�ƛ
��S���DGbz~�ٳupxHY�ǍLs�\��E��:{�o��d��U�CqyD���p����'u�&�]�|MI1��{Z��x1��;���ͷ�9ɻ�CL�D�(
�V��Wbi�."YHa��셦�������a��tIh>��&w�����a?9��Q��z̗#��L�U�yF�Pd��Q��Yz?����fing�����wĹF��C��׺�\!�0_�0��~�^�˯h%L�Kk6�z�9\��E�V�x�o�Hv�?�]�%V���~�
���81��4 >������3��2~�j���Ò�[�\*�Wn72h=���(�R�k�D�3'$��m�𠵾#���@A��v�9^�I���5+WRD,��G��"���Q�9�Ո0zˬ���p������-�0�T�MF&J/1�A~"�t4��	�V�F�L8WV忦��ڼ�Rٿh�5�&K�"��-�8�I���갽}1����+�]�����ȼ���.�ڿ�q���$���4��*x!c��°�?�[�璴�/�gQ�g���3{��;��	;��S"�B]�q�8�eG AX/�WTo,����+�4]�!�����`�@�L�/Ն�{��B����o���D�
hCk�J{q;y���g1���YBvp�[�.�V�QX�.#<��
~#	l�Y���A�A'��wB�ۂ�#&H�8�$���%_rHHYPvS&f����~��g2��^�+P^<�X�P+��ؔ9�
�C`�I���SG,qg2.�n�N	'���b=�>�W�=�R��T���A35�Э٨�D���\� r��ե�������a�R�vJ��B0nD�u.�B+%��]����3"������*��-��������5C���볾��$d�<5�:MfN�]�|������ܭ/"|qԂ-*Ӷ����L�*���W�^�UV��d�Xݤ�t�����������{C��T��I��a.�kA����a�F�/Cx[i�`TÒ0��D���<Wt��hW���B��%��7ύ�P7A�� e98�|R����PU%�N{�I?Gn��a'� o�)K+��N���S��`��7 �*�Ʈ�4���#k4N���Q��D�NעxD	I��E L2��V���JT�V����Ƃ��S��	�������J=��ȓ'��p5�ܔ�1��䩚�jgj��1�u���n#���!��Ӧп0�Dc�s�z�����u�<uYe�#����(��(�Cg.a�q�ʴ�w�s�I�4�%�Kɥ�@�au�TVL]
��}s�wc����� �2ä�ὕ�7���Ҿ/��Nj���Jz�e��[�������Oڶ>U�r�S�R��G�L�t�ŀlshS���Y^�ae�j��O��r�4�o�d��2�(�+@U��`�3�n��H)�%/ҭI�E���mEE]�;�Z{o�VB�D��S�q�,�X���� ���?����K�le���W�k�fc�Yp��!�0D���|�b�r{��y=�OA�l�uԿ>pZ�����l� �Ħ�_$��P3{�k�q͠��=�+L~-�:M˾��I4NE�-���:nL�.�K�ݞ��I��&D��̹�{�������'hHd�"Ay)V�Mzs�ĒV<��6�8iN��ض;���]�F���80�����-�f� ������#�C:��7��P�$�jiM���X� _������o!��R�J����ߗGZ�n��C��q�/U��[�����A��Gh����o�O�|���Թy��r"�f#�ѩ�z�1y���~p<����zʏ?I,xy��"f�#�'a�Z<�O)��\ivm�X���+]i�ߛ<O6���k+d��Psf`Bo�5_�o0 `
/��a,đ���,k�����~�Q�6Y+*��><���,�3�7j�Ƅ�Sy�4�(V|�-��}Jf�`zkA(મ~{z�]�j�z����-����}�g@\.�3/}��\���1�.��\�t�\7�;v��j�\/�w����	��O芿�U�U'C�Jk�T���+�
�fgXJ_�
R��F��W
g��ŏ��[9;Eb��^˂G��P��'^� dKs��.�K�\h �_U}E����M�xs�q)�U ��Y4�(œ�5 �� \A���/��M0B��(�6{�Se��XJ��1����u��?���5a�!�6�I�p�9x&A��b��oJ)�͘6_R�����!�i�D�؃c�Ɯ���|i�Lb��Ë3}Q�+6i�Q��=R!�k�̈́_�}�"��]g�W��u�X�5�W�U� '�k"#$�K-> L���$�����l΄��ރo�Ǐ\8%=)�Ney����!���I�Z�/t��,S"��"�_Y6y��i_k� ;b�C�kӴ�+C�M��E��1�:�- ?L�;��(a(.EŜUyN �#L�P�9U�J���B��>�*���g��K}��+�D	t�����R�.�+BR�Ì��`�����8&���}���$�Q'�j�g��i�IW��k�Yw!0>A宧�����b��O�s&X�rѣ�x�C�|z������@cGtt�C_�����V�ò��`V�2��x�rbwn����V�(͈�t��ZQ3�Uzj�@�Aqx�����p2��FM��u���
�����d<!���2<E����VP�i���wu��ؓ#B�{%��Ъ4�|X7�y9��R퉚2yO��0�.��d�
SPPe;�E��)ž��h.�ki��E7v��2��/8����-�#2�z�j1���Γ=���Ht)��0F=�"Wm��:.���N���D�(e�6?��ji���0S�i�또6�m_��X�<m��sN�U�	E!�߅��$o/k~��a��FQ�0��2B�	�/��C���Q-�w->��.)f���I��c�To6��/�X���5���6�6dl!�s~"�=�TS��kcUT"��@`�{i�{?SV�p�w�Q~�7<\WE|�񛣛@g{桁}	o��A�Q��3l�]�{���S&?-��t����*w2�w��'�j��7��W5y�����IlY�\��O�ˉc�BR�CDPg
}��Ð}�DԱ9����]!C?.-=]��.��d<n=?��v�:{����H�{|u~5�e�ݻȗ��4E6�_��@�s@n@��3�8
�v��D�q�y�6��O��.���DL&�s�;���^L�Tו�,z> ��bE�ơ�g@�� �|S����_�_�Y�6wz@�j)�pzK�Oh5��Y�(�K�PZ	�����s��l�_� "��[�8�k���l
�c�HƏ  L��B.G��#�������H�C�)y0��lV�U"��j�?���)W!m��@S�K}�Њ�6�w����r�����hR��U�f�]�Gk]O�s�x��-�t�9k����ޤ�f���{"��<��i��Z�#�֋
!�.�Y�t�)&��a�\ӂ������!_�ZJ�(������;(n���  �#�ף�zbs���lb�������n�)��},<�U'dY1N��]�A��a�t}��WC:�ly���D�iz9~�"t����^�_9/�l��a�\�_��S�D�kN�#���l�,5�eE��l�I��eJr�����ڬ$Z�I +-ӂ���ĕ�����՗�c-�.�IQA��q�8s�e&�+9�}�	۲C�Dk[jg��e���JL	���2P!����)��e���n��4���"x�h��Ъn�쒕��Q���R�^=%n�u[�[⢙Qc,�Q��<�ahZd ���'A� r�+��{����.3��!_��&��}��N�*"Dz07ލ���l���B�i22�)xs	EK�]��L�h��M�;&�ܜ
��^�|Ȗ�������ۛ��f�QZ�bU;���[�eJ�m����k���9T�|���.8��BJ��e��ŏ	�IRX��DH�FRL\;
����Ww�9�I�z.�Vk͔�7��3wQ���#|Vx#3�3ȝ�����}|��ƣ�Ye�j�1�5
+�r�p��E���j���Vl�H��ȺL�㴦�S�����OU(�W�[s3]��Gfoſg�N�/L%R��I
��x�g�I`������U��ҿ�ƚ�.G�[�����9���V�D�u��V�s�(�ڬ�M���r���J�]>jTF�d��l�±cR������@+x�9T�#�����*���?�-!�W�Υ��ކ���a�"C'�;�
oBv|ɖ�uo�D��*+՛{(׾V�ZD�0�[H��P�g )lF+�²��|Ým�Ι9(aH�!��&�ہ����^��\����uQ��uJ*�0źbv���W;)�S����!�U�qi�֤�#�1U�j�fv0�e�3d�i�/o�UO�]�K,ﷻg�M�����j�r'� �y]p)��X|n�&BqV�՜3��j�B`d!���ʬ�e?쀏��\��gϺ��S8��@� �$�-�@���y�jA���W8 <ۄ��� }�|8g"5Sm95�0��/ĩX�E�`(T��m��틼�9L�)"�%�X��M��3d�Vw��>2�*o3�� s'�T��hWg>�R��8i����U�\���RFI������Yn����l/�>lC���um(�A��UO��6/a�(3�\�TBL#[�Ž=��H�����aK���Y[	����>G���	�����a���:�,Y~�}L\���0��IG��C3qf�g4~�L�	�6�A%K�/{�k1�5��w�3�dT&k���Ll��G?�+"��A�"h]��gjC?í}��?6iw���me|��pL��¬m9���4<m�#��,ޑq h���ݛj��ɳ�'�B�ͺ��<=�W.���[ �ÿ�t���R���+l�~NHƤ��C�d\3*�4>�c�����ߎ�/'i�*�M�B��vmw^1p�>M���ݝ��]C�fp����8~4�U6G�n\cn��ZbK������a$��,L�
D�\�-���B��uh`�R�B��9H�\���b��$����ӯ���ǥ*w�s�-P�<mj1����_�n?��C�q��^np�*4|�+�`���Pf� �zc�%I)ďŨ�ݥ]�gl��
�.b�&L��'A��[$ڛ��V�,U*����rѪ��Y��J|������F6
iJ����)��6��[CV[�=�Oߏ����Pɂk5j��s�߶7�-�,Ψ��#���䃔�V��c�cɿ=���w+S��گ�"��-X�.25(�8�	^e���£��ORЦ��<���'+�d ��ET&�Ǚ�s.^�` 5qIW���%��ha���0��0��Q��0�@J/;�;@����QS����X���&2��3S����1j9�W��c�wXe�r���u�7��ŝ�����␗TwJ��I,%��Lj�u�G{	�ɇ=�<=�V�h�(w��_��)ą�{�G��͐��G&v��,�)f��!]G)�(�ax <�uS�5�M��$>マ �Z�*��cK��Y�(Vὂ](>D�}4�E@.y�_+���)�S:��jn��M��D���{�ֳ\�Y
��ԫ}'#���vp(jX�	�hn��ޚ#@�¹��Ga?1}���3x?ID���u�Q�ߤ�x%��S��|��y%�1wi���i���|���i�U>�@�ʹ�q���e�+�w�/�C�W�q��\Гg���,(mƴ�LGl�,�~(�I�"�O>�n��x�7t��m�h��X�B~ =��85��5�	:{m��-��Pd�#�x�a�	��@������^o\��H��j-�����S`(���Lc���#�B1����}�<W��CM�CB��4hSc�@�i���ؑ�-�[���yG!&_0h�U���nL1�*���;��؃�-)�YLO�P�K�{Q� #<pi^��8A�0zl�v�	�ZU��7���h���:�&��rE�%Hg�.J�W���
��+q}��n��&�(Q���~�yx�f}���0Y���|�c6j�����y���*�H������W%E��s���b�&�7��D�]��E�9�,%2jg�����Q�hA�[ �Z�,�E�MM��������ᒮ��tU�E�,�6�5L�l�7&1�s'j���Ƙ܃.��T�m(���^��Lq�v,�;�Z��A 5����Y=r8���.s^���?v/Ț�0d�B��_:R� �����2�˲}���{�Vj�����x��S˟FPx��&T.J�MP�GF�%C��bsbgex2�U*+ns��'(A9��3_OzP�K|��ǻCR(�v�g�¡ݧZ�s���^^`y�&H%)�1��4gUO�8�[}J�+T5���8�5�"�x���Ȱ۬d��(t��K��e��"n]������}�̊l�x���Vp0A��8J+��_8�����u+�����Hlu����k	�O��W�a5������%p���O��Q�>?aM	2t�b�o��["`�aP!��eO��,��fa.Q%�L@���*�)��>$O@�r�t�������S>ٸǰY�9���!B`@7����F��!�|z	?f����u/ы|�nL۩K��}ZQ�̴޿�
�
m��xx�|��7�ګ(�`:�����C�$�N˽r��͊�V�9�`E��̋�i�ʐ6�)F���ߕ0m��܃��$�F�'�'��B�NC'�BZ��o?�����7ө���K�h��s�뻠aʶ�%	x�@vNc�����N��eӣ�&i����[]]���NZ?s�l������s�>���	�}2<�4�"�Q�ξ�"���f�q�j,��#��?�[�u/��]��������������}e�>�3�*��T�^��$�n��k�
��kgl��<�S��S��m=]g������!J�0�r�>����a���m��?@`b�	���i�ObY�`oF.=��>fl��a��d� L�P�d#ܔV( ���߼`R��B7�5�;g�Y%O�	|��ͬ�dT�{����e��h��+�=y7�F��'U���5
�������}�}���S�'�HM�Z��#im��G��v-�i��萍��^0Ҩ��?��5t2-QVN������+/��߉��ب�ջ���m���+
��m�MF��\�Z�=k�����t�3)��t���ʴ3c�t�����sEw,��5#4?�� 4��9�:QCמ�ܘ����x��y��)�����aN��ӐR*����#��A{
�)��E�o<�˻Y�sPd���T��V��i�92�4�*
X�jp���6dK�ݞ�Y�������B]�idri��9��<��K;��w��c�q�3"�l�z:�k��\�~J�/ǹ��B���'Y�_Q�X�ߪY.nV�p��t֣���bU1�<��t����$�òO�o:��I���R������<_�'�l�$`�GTab�>�I�;��Z	^��gZ�b�m#U����{f>'Ib��ʀ'�>byzK�57�:��������>�;�Sn���quo���g�vB�a�nC��Ƙ��I�LL��I�<Ԧ�C����+&��+�a��Y�N���jD�.��~{쵼�Ԟ�X֨��f��A��Fq�����*��V�D>�t��e�d�=�-Б]�/�f?Y:���o��r�(���u���2�P+���%���ĺWS3�i0y/��ˏ�$zv��AU.�nxxn-����T��f�8u�^�'���hp�=�"�Q�)�p�'R��n<M��H����^�R�lk��^xD��С�
�k%\�0g~nSʈaZ'$��������YcG�L?���|���{�i�TȤ/2-��h���8�h5��W��q].�V��O��c�I5���1`��=/�Y&h�:��j�Y;ģ�sċ�4�F��1� A�7O��Z��Лy=�R�)M�y�S�/�T��2Y6�/�0EO��������N_����x��_ѐ��uJ{O[�$�#��-����p�&�CF\E���&p��6)��G���@�?A !t��S�A�]�5�	���ROi�\��*����?�!�~Y�@#C�V{��� u��Mi�M��D�HܛOS�o湐����~�;'��I�+�� '�:2&c��K�֕�zl�h�D
ZG�oU^y�:a�	,���=���N]Zr0�c�(}��s��_���P������?d�~%i[$��YL++i��Ч���T	�����0g:j<(�ҒC���{x�d�Ô��v��g(!��ł}�z�������Y["O�J��k�Y01<��O��
���x�O��-�a�����7i���~��^�ҠƲt�ǖ�q�G:���i��Z����(���Q���_6V�/������rPhN��.�h�uʔ�����}I�<��Y;�m��ۧ�]�#ۅ���8����jޫ��aR�`G�2�ƨ`
�ʰ�H��6�p.�Q�!2�^(W��i?�� `�ILy������肼4_4v��*��B/E��I)b�g�*
n$��)��DS���s����������Ȥ�{1�����"ɪ�������!<�1��b�N�# 6Fɥ7�*�J�؋��WQ��2W�ZE�ہ�eΈ
��f���\*�8'�KD�/��k2~de�qO�Wa�ޟ����?{�K����XV_�%���X����S^�C_F��A�'�X�ShG���E�p�)¼�����!�d��uP������Cc���wVwN�C"�h����Aq����v}+�)�j�;|��em��=_� �5�۾�!+���-����>�.���;%"T���[-zdN��x���fI�<"��I;ˣ�,�������[_`,5`b{�����C${H������B8Х[�&<=���a�=Ș�ԇ�d�d��^bF��L�X;�S����bp��4�WOQ�E�ΐ8�j*���'.�ܫ$����}��gn���V�"�R~V%����[3u��y��W=�<�62�k�v�N?@Ӓ�`���b3�G��~��k�?lw{̅�V�o����&�6ZSvᙜ���﫨��W�Wm�gF
�-���DJ��<���P��d5������j�3>�M����9KS�BƽC9�25�����;�m���/fR����3�d�(�A�a��`�M5��瞫w��D=U�Kr�ah"� ��c�]���3���JL��9WU�$i�ɓYƳ�nk{�ʂk;�6ce�.�|f'"�<x�.q������#�ԗ!��!t�ԃ%��������
��e��mc��䇣{�|��X-{5�9�(�"��d����1lgM��B�2�J�VV0��[�.H��E�H�<q�7.�6ڑ������huMҔ�=Et�n�\}�k"Y'O&����! D���a�)��8����sW��ߑ�'ٍ�<�3%����l����2��m��Ġ�J����{'��w����o�e�Tӽ�KJ�+�᫺
�7�9�� r����v����Y��ggU���hX� ��{jVy;��n<�lq�T���@zɛ��DH�����\�@)+���VV#e�,G�c�,%�<�sڶZԐ���̛R�nDۼp�9�?�9�zK.@�)ZlDXς��该{�:����>��͗�Q�j	S��i�m3�{��x�?�,�oeE�Lӣ�K��We�u���AN��aʳ-���"}ݠT\�D�n
�%���"1�&�8jg~P����֢;�%Cɷ�t6��lvx�xRK�	� #�Ӱ_�^���SC[�X8��Q����cB ����/ڮ�/�ȩ}�IJB���u�a�;��,�>�\��H3)J�QT#t&�)��Z1K�A8	�-Hn�cT"[r����(M�_��-Zyt�������@��%�_�E;��1��*ό/��J��~��������;�7�4M����)��	aj=NKO?6c����7���*oE'�<�x�W��t20��.�N@j>u+�u�N֑�g�q9r�V�d���mQ�*hp$)T�K�r r� U!�b���j]	wkYY��{��q��|�Fp%�4���=�`̂���.�[4���GX�ϥ��r9:�@�=$�!�:̄e#,{A`�Ƕ�أ�̭ p�,�ea�	�٢���u�F�T%f��h]�Y�l0��eHyW�G-P��7�5�rU��\fMOT�b����z��� [��n,Ё��w��?I	i��@��Ecf*�l�2d�@I�/��w}<Qj�w.u�|�F�F�4�(�Z�}��.>�`�`���D<�q�<�dz�p ��*ڠFiI�?��<�9G��_�M�K�<`F���\&�̓ST�f�]SK�ו��gJ�3�Ot ��jE����c�e�[���m��W��?� �_���6]�8<�<j����Dك/@���7��mԋ�����u�ɓ�iM���	�'R�X��R��-]6�r��0���uG$jv���k����"o�P$l�P��h��5��prV]]�"�_>��Z4��(�!&�Xl�"�N;��2*J���RKEk�[�����k_��IY���e�w2����j����&�x�<V���D�cI8^U���8��"���Ap ��ǹ����%Jn��Г��\ﳻ�I+n��@��O08�/1|�E���}<�^�>��&̘)+��v�+tW���W�J��OB@%J"�fQ���I�R�*�~-�'&`��P�ί�)m�PAB�����¦q,KZ��'��R���R̉]����G�d�V֫f]5��Jsem���)�0իB/p��4���cE��R<�ۼ�*l���̘V9�p>�t{��=�:L-�Z�6r���bMs���!���|���V�����u��X���i���3�������=�g~�?� �-�s"a���;��U���r#������������+hgw�`���U���>�.�-[�a�H�8�cz"�]A�`@\��@��t�=z5��F���$�0��>B����"��� ���?{����� �5Oj�z'}�CPK�B�����L�Fa�.�/n\4���s����&tk�^�6�3w�fĝÐ��4��]$K���	�.Ի��^��ϒL��b��J����Q�r�4���d�T�5a�D.�w��si�U�*�D�eY��>�9ğ؅�4�ѳ�1��@��s�j����<�P�w<�Yi��.�&�L=�ҭfp7->�pO�]��9.�";�@��C�M�EZV���ΨPM���N��*�'��﷜�ێ�obȝŭ>��+V��&�Vx��"߀{����(V
Zm�n�&��@:��3%�6 ���%��D.2)�=�-7P#az���/��P�-:@����xvs��,�#��v�&�F^Jz�5^��P�G�l�d�j������YqdH?�\��tta����]!�TS1�j:��p��:�<±�7i��!9*����LL�c��8��5�)��^�r�z��#݃�WI�S�����DL6L=B��B ��n���Dxg�ng����6i�;rWЀ����[�vs5��cێ�Y$seD�I@��ZY������X,�g�ix�v,�4���Yz�V���&hU�3�����|�x����f:�ٯT��l ��=L�:+���1i�V𙕩�����[Hl�+�J�j�9H��S�{��@~��~R����� >��!G�n�0h>��o���}����ﮎ�R}�� )n�Z�UK�:B$*��p���'2�<�"�+G���Oӈگ� ���x{������3��qC�����E�b䠜��(}����1 s�:n�\6�~`�#9�W��d���@�&LW%�*��}8xE���i��p����.�矷вZlk�����7���wn�x�����tޛ����x|�;u~�i���8p�m�Ʈ��m�D��$t��.��
����`��52���:U2��b�#���J�j�r���@\Ion$DXt۲��'��T��:�a	

P��u����`�ϸ���	�O�\��c6%\aV>�`ꮶ����kF�0$�*0O��"@U�R��%��)�"��ON,Mb\#
񗉣���͢�Z�W=�$�b�;?�H�6fb_.L�"�\����-��^y-Gq�ݟ��ON���#����Z&B�~ٹ����c��4NF٘��1R	d�x���G��B���6Ӟ����_K�����Ag5�U����w�u
���l�M�\����X�C?��!��`0� �����&�r��@i�s��ȍ6}ј�#�r�jc=�S�m�$���4e��5q���Ɇ�i�=�t�I�^l�)w��?$��7ߦ�lb$��c0��b��^�K��;�MJ��HQ����Ӽ<�梥(�
��[�Mx���r�R8~@���� \X��"4�$�
 �K���b~�<��X����T���
r");N�mƓs�
���*�Ɣ,[��~�|c�pm�~�l� OQ����5k�� c˵�r� ])�)ࠖr8ԋCP�J�cu���#�����,ʪ_V|�ﴸ^�A}����@��V�E�F������`f��z�6Z�D��h~&F�+H�=Z5	��y�'�q���V����UW5Y=~�	�����=.��Is����6��	�2������q��>�ҹ�;�D,-I�~�|����QӆvU����G��6,kCL�νo>|�7c�
;�_ߒ�����,R�<�� B aE?�%�58-)�.'z�g�m,�(�Y�	���veM"l������;hx����M���:<8LJ�/܄Ja��^��>u�ͯ=���~��]����@���%�1��p��}-��GV�l�T�{\�ɋ�kV�f@�"�-Ss�DG(^����ԭ��d�+�<d��3�I���d����$��5V�<}��9$� �da|��6Bb�0������5ֻ���H��O�B�� zܾ�j���iw��o�a�rF��b$6�˔V]B�lz�Ym׋�09n�!����ĉq����o�2zr$-��Ӥ�����+��	�fԽ)P��u�e]2֯Z7��|4��j�ٌ�M��ڡ�U��YwJX;�\<8x�ц6�h�(����C�ő~Hgz;�49�⭿���<"wH�O�^kh�oX�h}��E+IbZ~�ir�xM�N����)rhg�i`.n1~�$a�[
/����:�xo�n���v�y�S�B�}�(K�ӏ�ʿ�W'���=m<�;f���'����>�^v��&���R횙���[t��,�x�hN�n����־�$�HP��9 �5Вh����s��م�f�����E�LH��P>�ҷ*��="<��O�%�;��
$,KV?<�^F?��4@j�Rܒ(��m��� �<�n%w��x\�[u�e���������0�sUfc(�q�I���8�*��Ʒl�couow��4���ֿ_ "�՟,��F�K���o�~W�54�hog�#��w(�FxN�yN�<c�:6[��|T��.X����(�u�}/M�1�E�$�ҍtpS�qe�:�'�L-�A�f�+����(A�����?�a�S��	�wZ���b��ɽ����K ��V��v:�GS̐ms��;�X�E��L�B	�3!s�+�l?�再i-X�R�$1��`�#���T�DQ#Hɔ��<L\V��x��v�l�..���HYN��]�ڈ+갫�==�~�ACmO�\U��SȤf*��C��vv����z2B�]��p���(b&�1��R��5���j��_��kP�5��4OM2�H�k��Cp�L�*Ý3"L��~F���zڍ��3��6���~�˼e�䁷��5��w{V[����PVv%zy�K��/�hzL�x�
J/#�z�Ete(ž
U�0��V)Q���B��H3�/G�ha|����%�nyM���|��[�n �&j*�@�[@� a��gw��I�|���Y7����o&��?�z<�$	�����L�)�e�j�s]�h��B�L!��s����j�7�7f/�����j��R�T:|/����}.�̤DD��n红��R5�U*[�P���@ߐ#�٭�Ϳny[$"��~z