��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2)��Tق[�	��5�Fy�
������~�}�Y����%�$Z����!�:�O���<�K�G�PVP"�H��TV��W��e��x��Da�	�����V�BK�*��s"C[v%�����Y�����N�ϑ�m2(ѲQ�q��kY\�籾q8_�IagSPvY�a�έ��7�IR�N�50�[�U��+�Uݥ]&�K�ٻگ��`�9/�Fp�cl��{,�?�ILʮ�B]��j�Ը��+��EFN�G��T��\��h�r�C�b��|�p�4r?�P_W���NY��Nm��K����_����5��i�I^���sC��y�&��Kڭ2�0�����}R$��X�NWF%�"fuD]��FJ�I�"K\��~�.B�f<���<���c�D�9�Q�Y	7J����͙��Z��uRX� M��94��sŤ�egE�x��_���C�OYu�)���ST</�@gTٲ^�a�w^	��1��{"�H�5��q�V�r�W�~&�>(��_W2\^?p��<)��RG��LsL8���XH��wr8K��2�JJ�Y�OE����f�t�ek�\�h.����'���Ȯ�1MAU�wGV�%td���2�Ӿ���.��n���	��?�ә'�M˪�G�aJ��"�� g]'�	�2����J�Ǭ�-��+Kwͅ]_'.)T'��~�8`��gs���&쌇��6!D���]i>Ow��?���Ba@�KPk[��ԋ�6��{xB��O��$�W#�ʨ�T�f_���x�3Y]�ޟ�a���/�^�6�rhn0C�^�h��_��J��F�4�'R�{�Y�h��KCc=`7��c��a��$���A�J�k�b�kL�$S��>����X���(��	��u2�q�?��l��~A->�v�AS�{1��o� BE���ak{+�U�\Vx��Xm�J{�B�yt�
��bO�=�١r���<���,Ȩ�8ڵa��j�w+�alz���Ze���r,���a�0?��X1k�T����O�Q���e��& W���vx]l��C���� 䘀HF:̞k{��灗}��)N�����c��SAj��&�Q��p��oN�P%Oz�V����Ym�8d�ۙ��#�!�X&s�g�t��y��׌�CV�Yu�̘`�G���G��3X��!���������~������b� ����⎮�6�� ����@�Ȯ��	>�,0	�}V�o��@��Pl�:�9?:��`c]��=!>!E�D��:���|o<���~�9���,��~U��I�ė��$2��I'kl��H��,"�T��-��d�f��I���Y������M�9�f[�U����kA�D�����I��㮦���KP���ܫ`����P�P���vb=�rr��L������
q)flM�S�w4a<�J�
�ѱ�ɂo�Bցޢ��I����u2��ތƚ�r�j�òU���p�YL3��Ѣ��93W�Y��eS��mx�1LgX쀍|�s��H0�sǘ\N����)2q����d2w}Q����'�ɖ�F�H���T�BPe�mU�dt��P J���f�mz��VyN��b��^�<ˉR�r�u8P�����cq?�T�� 8��F��m­D�6�K�\��5��?H���u�EKF�w֙���ԁ��'C�Xl��ƞ����-U����d��O��ޥk9C����55BwA.�e��q�U+���hS����sH�|��C��W��%Zpꔗe�Ū�������[�q��l$�QoHR�3|��E�Ʉ�v��qq��NU�}�#�42��i�mp��U*�Y�N��tx�8<��&�a�͠�m���/��9-�T���/)�L��� �f�~V�s��tb����dHC`�3��}%r�Ѱ{lAWx>
I���!$�G
'�u\��C���I�r�Z�P�h����F��:;�b�,h�A��־�Z4���h�zL���{U��|Kvl�Ӱ�.��O!�+^�O-#�r�})ݷ���6����Uq:�H��T����f��>l���r��Iv�����]�ϩ^���^߯�R�CjK��9�\1�>M�ϛ	O�iX����$��F�#�7R���>���W���pQ�(2Ԟ��&<ŭ�U��1����Z#w��Ȇ�,0� �LqD�����e�����t�C˭n�ӮV9o����A����Z��b�N;��^��V����QQ$��oH&�HLE0�T{���þ5g)�!'�F��1S��1��3�ɄO�O�U7��,k�j���w�=�=ߥVgBI�2��K�@�K���7�1A�(w�e�/<�:�={lQ�%��	*쓂
8�'��4;�J�	�EUL����OhFa�����7���\�Lk�ˉ�˥�q3`��e�1���
��Ԣ�I
�c���&�J07]6O	>*�*�X���S�>�v+�Y3z� y�JDO����FZ�"���ګ4}H����<V	��"Ծ�+��5��L����"�Uanh�R0<xrv��^5������{�-Pe�.3�+�u�Ys_g{�u�?q:Ry9|�W�\�/���� �׶�-%^EX���Gߓ�4��}]Dq�%�2��e�D�<h��'�G./�»֕���A���[��P�^��7���d��k�����G�HU%M�? ��=7�|�<t�����Tjv������C%���>8�ј��I��\8�:�.ouԇ:`��������W��Cre�x��.ܐ�G�C�m�兽<�8��0&Ɇ0d�e��!��I�7��)��x	�j�@����ă
V�w���y�,���a��%��5=���J�
ky���f�h�`J�}�G���Oo�a]u�R?#�e9�Ao���lC����]��V���A���S�
@Cgp�����@A��dw91P����h�*�q�j��:�	Qt���˴�;ӕ�H���zC$���˄M��S���u�?f���gQ��u5R�S`Y�Xu4���v�- 	�H��g��fm�{��V���,!/�/�R)p.�y$LH����@��))5J��
�p���]�x*�4�7b��Tǟ��}7��7l=.i��|Q�����D�6r�L"�U2��X��p�lx��U���I�4͇f�@�bq�r.��>2qM���'iJ/�b>�W܎ ���O�صYE������%%�P�����^��k�3�����r�����m�;˾K_��q��_ma�� 2����{&E;z�����:�[߯
�+���Dv�n[��J�Q�Z�1���j�����x*�DO��G�|��)]Z<9�L4aBS�d�w1��7���u<WR��J��관P��|�3��Ï���]����t��sd&�4e7�>җ��Etf� �m�g0An�&�.�b��SM;�m��=צּ��BA�&C�}��K�s�@�t;��:aZ�-�R������m$ޫ�a�d�ٳ���A�#��BD��>����$ŰK�k<ع���C���N�!���0T#�#�=��Q��V�K��4�t�x.�3�<�ļȧZ��jGZb�%�@y:��F�5�`�\��0RN�^�"A�Y>,A*#R^���jS���ͯF�,m!v�����Cjg���E���o5q*l�k��K�p]>̏[;uY��H�����P�j��z�&�u	�m��:�]�n�T99�̇��(��̋��S�LlJHZ��m�W��W�
C�r������VG��,��P��J�v͗*p��?�;k�Q�g�Ъ����&��Wc�� Q�h<�_�14ĊY)��;�M E�E�x��	�~�'��K��M���*	'Q
�6AS@]��C��ky����SX6�C�����|�F� �ΣH�ur�|ԓ��:8`�e�Se�V�8a.^æ��H񛓶ZS��e(�/ #����N3sy_��x�)vu�� Y�i@��,����pW4�"�X�r*�e��%��?l��Q�E�L����_
�Q�,�H�@��&6���D�ZO���:�Z�ːf�{��X����;��rɏ��(v����)��kf�ފ�U�(D!��?���h��G�`�������	9Z9� <�z��Fxs�*{T�֗��1�f�d�9�D5X���x�>���$MB���/�������2����(�eh\��9�t!s>^%�!����e2�,�M�����.�������4�B ư)�X'��C������e�ً��c�
��at�;_���#�R)9o��YFw�;6\D�t_�C���Б��*A(z�ŰN@��@O��f<�Q����#���q��c�{~ۀß��C�Ԧ� M �����,bTԅ�Q1���2;Y��
8�8	��6e�A�n��x����G\�Ƨ
��|�чj�TQю�3oT�?9+)b�mYo��ȑ���C.��>mS�/�d��,E~����#ˇ� F�Vf�C�#b�Xf���J<��4�6ú�ƞ=5qE�������T28������SF�5�:�["5����3 c̰�@W`i�i����o0��:k:v�M�Ze3{����94S-�5k{�8xPb�+�`X�⳿)� oy��k���f���2CMC���)9�X�O����~�R���<�=u���0�6չ|�R���E̪L�d��r���d�+#�$ 沽n���'S[��y��3n��ҿ��;X�SO]X�yc�=�5�!z_��ꋤg�ୀ���[�EM�#�fa�vz��_�
Oww�!�sz͡���\H:�5�@2��@n�Of��W����5Ӊ(�c���U�oHjKD�����-s�p���ؽ6�KC�ƒ�^Pb�v���~����Bў_`A|4��P&J�:�7L�;�@d��O��V��	΃���V)֠�kJЃ�Q$���7YU�uGj��pc����+6�ԁ�硭'៳ѡ��t(5�-ɵ��l"�Ǉ�|T�B����]У�?�@A���0K��V<��O4����.<O������?A��@U��Ge�WgBg�lg�z�=f���6���P)��a/�*��D�n�g�I��np��P8�7��<� ��B :{�1x�{��������;[��7oL�z����\�1Ѳn��}��ꈚA