��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�he�4����؃�d�m����Z�x�`o�1�}�}� ��
���}e5Jt�d�]�(�O������g{��q4��Z������ ������^���`�j�"&&�AO�'bu��� �?T�D�����ݵ�9��DK3a\����}����Ȑ�O K�м�Qݵ?�v��1�('#�u���
"�� ����%��\ɶ��=��	���F{�=��1_��TO�T�s�y*2�N���zז-pS�]Y
���q�w��}��X�;��Q�nD��XE�kQ8���5� ��}���P��A(��n�������=�y��C�a��3��J��Wόi4E.�Qn4j8,�t�Ч"��m����HFԝ��-�8��p!׌�Ĉ1p�򊍛$�1��3�8s�'P^iHU�)[!Az��g(�#������8���Y�w�x �g���y����g��k�QtS�X�~�hz�\���I���3�X����3v��>��q� ��	����8�#1��=�b����A�� T