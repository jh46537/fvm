��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħa�gU�]@)},����ע�>S�H���+ÏFfYc�A�*�0R4������h�֝�._$8Y&�Tx(wu�i�ٖT���ʂc���7/���Ň�C�����$����qyl[�k$�I|��Oj��P�a��*��x��j~W��ܶ�
�dQ�ä��q��Ai�E`?�Y��t�%���Y�L4/6Յ\Q��A��ƒ|��b@�5���G�(��U�Rk���F�}i	��S�U��sDh���Kv2e��R�O5eML٘	�h����	+rdW�,���v�!:e��S}��6��U?�:�$e+�)�s�|�PJ����	���FⳲ�ᇲ�_�D�r��i4�E���q|9)Ì���}C��mTuQOQ^��E�w1��yk�dB�#ۅD�ky�TN���+D�d��yh���\T�?u2��g�Y�r�����]Ww�"W��b�k��՗y����_ą��*N�ն�jew^���󳘡���4hM����C�x�h�5=�x��v�ޟ)	o��sɑ	b���];rR`?�y�$V�`K3��	i�B�FK0�S�Gyl(�� ��t��5�^���٥�;�]�����~�W
s+2�C��0$�~���=�0�4DD{Q�T�y��+�@���D��	�b�K�5�=*l� �����'{�,�@��6������Ya(}���-�|��G>m1�ES�T�R�H.ڔ���K��jUǲY�Ad��=�*��u�-�J�]�ʯ�����Njޟ/˨N�V�|�"�:J.�Y����jx�:��y%�!�155�NBL���������g�w��kx6$��*�W�g�J���{%"��H��D�F?V���"��c�O��a@^�8[�b��V�1Y��U��Ys������NN_��D� �3yU�y��m�sY��QA�qQ�֯�֕u�]#]0��fN�j���.R͋�lhɌ����
XFj�8��O.�\aQ��s�L;#���n���'�H��a+񎍱|�w��X���ĳ1�Zu��F<���CPㆵ}�3f$�
�\��>�����I�z�a6��	�ߜo;~2���AR�`2H/�M�քƭNr���K��یb0�̤�	-ؚ:��wX�i�Ѹ�M[�	�X6��h!������;�� ~�>H^����^h��������UדP���f~(�`���|�_�&q_�F6�~ƨ'[I�V���>L:���f��E�+��m��C�QQk�O��.CG�Z�)3��;'�A�e�Һ�a)~�?������e;o�(��"���+Ws��C�?�()�����|P�����3�x���'�*G�=����p��ĸR$�-8w�˚z���Y�������-��
�!q�K�7/&��8ή���ȵ�����ıƙ��j���3�\��V|��ڑ���7(�vk�*o4�K�e�M�N����}��A�a���[o���j�|�@�xܐpDU8C�0wtFUC��_��b���&��v��]1I/�.�����[d�-��-M���|����5��@��ܦ��(~�J�:��.Sp��^��{���w%:	�p��������g�-����7_�/"!D�x�w���ZXoO�:.���yF�[���&@'���'�.N��
���;�n[�838��eA�Aæ�B�}�����ڕ>��l}nݿ(S.!�Xf_��S����DǺnK��d�ȭ��[G�/xj�y3����^)�2#���×��b	� �.�{��:?�HwX9�9Ew-K��M#�K�|�!j�Z#���ĝNZ���`E��y��+j�g$i:�̲{�5�RGC��ݫ튞��<�X����隱�nMen��a��Y��b
Ͻ�ǴO�K$�2D�2��E?��Z[���M�X��-� �{�׍�\1	�/j�PC`Pj�`*Z��Q��[�®�� ֢���$��[I�x�K9�RVu��y��������~˳F�p�1�x��Ko��a��4��O&j5]��1l��Mpq>�ɐ'��Kw�Q��8�iѭ>�p�7���aT�d!a��@6v d�^�s1��@������Rv�O�g������sk�摈�'�^H.���wsr�N�jd8���$����"j����BI#R؅�}�◈�z��<	(u5Y�%�T�r��Ju������e����J��U�9��2ҭG)�i^�gΠQt�����({��y������UT�?�^�U�)��]a�k9��y��u����ɬ�����O�,gq�CI��y��!l����mL�!O�4�Y�/�lT�^���X6eY�q��=�⢛������8N$�#�y\U��]�+l�`��bu��?n_e'#s\��k��w�+lR����MPꞓ8A���N�]"��<���"��vX�{v�cs��pbjhZ�/�b���{�XTdӽ�ID�-���}�mP��k�NK�bһ�9*}�y��f���JJQ:��t_��B��"()ȩ��f�g�V��PA	�&�]��X�����\<���@��K�C�S"�߬��I�N ���.<�b�0/���iN�Ȟ��F׫ �I]�i6ȧS;��d��%���I&���;����t�?C0��(���E�P��jIj�h�;1~Z���.Bb�"�>���t�ѭ ��_-��(�׏i�z�n.��g >�Sh��ٸk�,�xYb���P��6u��%\{��h��AWǏ����,(��R��A#�9�V_i��/���Y�����&
9x/�������5��ay�D/��@2�+�[ᵼH�$�R ���O�k�iER�3;�]��|�Q��\%]U[ȑ�b����'{�z�����$��� &�>�Y�«�m0�щ\^�B��;".�)�_tg@qC�`	��KA�Q�.J#�:p ��>��K��S�/B�i�1��1la�:�U&G���$Q�oE���
���Z��)�tDZ��9�2tl��4�~S�Fq)����v��e��E̗Y�J��Tnd�Ƴ��UO�1�j-�����n��.�?�4x�Yc��L�WjG�;{��`�O7{��� �rj^+��Q�>��~�������,	W����q+������ݲs�*�o'@Zi�N�=c��ֈGQ����ʢ$��f��v�qFD�Vo�ڟ�_C��ˡcƤ|l��0L+k
p����9�����x`���P6��э^�w���� ���C��{V��hU@?�?�N_u��Wb��&b�8�V�ֲ_VUA��#�U@e9�w�xr׹�Ϯx���F�>���9!������C:�_������i��=����>z��C>^9��)(,u~�b-H	���N*ޒ�1iu�".�3_��l�V'N���?�uH�m�~�QU( �5�{�Y5�Vgm�V{��u(���)���tYb�Z?��*��J"U��_��Usw��i����:_We��=V�Fb�S�@4Ҟn/���:#�b��tD�I���_��Dv&�Q��߭�s�|Ib���C�We� ��(�&����׃My�n:=��[��:�bp��~��*�r�M6��mb��-Wf�-3b��|�/j�H�F�JJ?�!�U�N�q�6BvC�.L���鹐��]��on?���E���<��=����bW|ej�p+���߮�j�}�aWM���~	�B&a�B�J�1Y�Vk�Qf�8�{��#��V�	��S�˸�Z[��p.��=F��S�U����~ŉFx̯I�+�B�����L~H�������>�!�����\�7�k��R�8��j�s�Tz�g��VH,�L�^!��&�g��آG��RFv���$�µV�:P��@5����f��%J|��^m8J,ـ��P�\�u#�<[V�B��a�h��hQ��Ee�.���;�4���i��n�E	wث��3��j��>����/����3��fP�?=1�m�s��TV����6�0Β�����D鄦��99e���i��ىa^v}�;R�_��A��ޤ��E�EUH�k<�AU��7�w��F�z��;xޓah�.y��Z�>\rX=en�i@_�
}���r<(�
���� ��~
Hx�Pf��~񖓥�}�f�_��g�[ϩ�9�P
nM�&��l�y���K3���M}Z,*�|;��ݐ�1F�Bhy�d�bX'��X���kb@	>+��Ѓ),s^挠�B��T]d�?��K�/�īEWC�������Ks��(e�=D��/��H��+��,�Ys+�Y�@���A۫�t�
�~sԞSu�j!��QcVE$� ['7#M��+wf��ey&śX�t�$2Sߴ�����j�����RpY�" w9�>�Q��>Z��[���7���6�l��t��^i�~kT���NI�$sRd=!o���;(>����9������ԡ�Le���L��#�V�oY�{�ă<N�Z^��X�y�;��_s*%%;�p6��%��:q���ئ�f*�T��%���r�dp�:��n�ӑ[�O4�W)��qO-�Y��/�&^�\�
)Z��o�Hf�p�s���t#sii�\��U���&L��B��'�w��14*���)��J�;���g�`K�C�PVm��@E�C�]�'���u��^��\~��C����^WU�a�ԟi$�	(��r'Fq���_z�{�B�x�\8�gϵ���p^$�!_Բ<��0t4��o��aX	q�גP۫5�rN�J�q��q��ܳ+A;)'�V7�\Y�W�H�g ��K9�҈A��R(�S�\�Q0��g�snՖ1$Km�M�x������/܇f�{����H��7�T�eE10���c�,}��ܶc1op-��"0�e�����_��l��J{�$�S\�[ ����R��0zV�<��A��U،y���<��5|��G`��s�Tڅ.d/d���k_�(?��e�-�~q���nI)M�ZG�P_Aq������f�&�A�E���8��&r�pep���L�&'[C�+�DԮͼP},{�s��Rw��Q�C	�3�k����rS��g���L]g��(�Y��M�U�e|�&[fi_�`�YF�q�$�\�e�W뉗�˚�Wɰ����M��~$@�\���u�����&Be0����У~��*�;gm7�*���v!�_��%�z���u�0����$���U�_�lY9�b�#j]��A㥭�KΪe�0����n�(�ՄB�wo�6#5�u���8��S����W�=\B��3d�]�9����� O��q�Ұ�~���#�p��N�%ƚ!��z��Y|>ց�L�)v�����:�ay�o�\ph�Ĥ��A(����� �\K߈l3��u�*%����,"��"�t�=kZi�2��<:��R�#�V����ɉ��%=U��Tc���)땍����J� 7�����$3>xJ���	�&}����*��g��q:�tgW�TX����[@�ƹ��j��ݐ���>�@fb�M��5k��
�-	K��Q�8��A�`*!%�Un4"����*K��^wN6D�"�3w�f��Y�m�`�#�GU>L�
,��ώpæb�	�=f� UY+�T���E��.��W��W�A�PI����ܧasz�J���f�<�,��YTN���H)G�9�[�ke��q��In�JC�\�b#����Z�O�Y@?/�\K��/���t�`���j��8_��!7�=O�U�hX�XNd'�#)�"\Vo`Y;C��?j�*e�K�FHh�$�����Q�8s�$܃��k2Q�6Ne�%QWC����s�1Z�v8ؾѡ$�T��Ö^^٩T�IܶT�¡�?Ki>f~�9��J�=��zr�Jimw��{�j�pN��Y�%yB6�]�gg����L��!�f�8�b��?5iD���n�v^��m��͹U'�2T��Zag�������e5c�q��2�ܝ>)�f�U�X-��&#�)ha�&�8��;o�4���I�-���FZ�t�&�(ΰ�h�,j�=a(I3��淎h*�s	M���4"�; �~f��v~���,_�����4��%�ynYo�'�ǥEDT�cp���D��H	X�U�zg�QG#�j����ݲ�N��y�$��Z]�<y:� {�a��:A�ѭ�w�n�N�K�K�R�����6l���Tu�q��`t�"q:3��dE�,4��nԿ
�s!�:lFJ2�d���]��u��)���9��Cӫ�C����$�K�;eٖ�-%��UM��IAo?v��C���U��9¬���.�hmNt�f���&��<�*��A������H)�b�;�b}�i�up!PR�)��7��qd�*2��Tn�ڮ�B��*J�N��'5�L���\���ow��p��~�Tq�ܵ�����U�ɩ�9L���Ҹ��*����{�Դ�
KřzNwy ��B�W%�=�o	b�v���vF��wM����\���T<�w���Hu>��W��cA���c�{����dM�-tC�1���-t�p%��K��앺%ߋhװ̟����0���l���I(�A��Hb�m~R�)ΐ��(b�F3X�q�W[�&k���R�?�cJ&1�+�����<���HH�4���U�mW��������$�[�
o�����w{�UQ�`�*D��S���>����|+$�<�ѻ�gdw]W�Qwޢ��b����b��a�mU�I�߉pmX��z1�,ٹ�x���f�U���H�_Th&����iQ�k	H���G�(>��ߜ�g���M�km����BB����	>1l�
��(��Tw)EvS��8V��`�Db����߾��sV��x���TJ>�������XҳER�x�Ď�&�L������>%�q�vS �E����|�R%��=�d��X���p��QG��L<g�h8���f:ǯ�1_ly��SH%U2X-;��������p�ַgUb�,-5o-�G�e�y��lP�2|&����Q�B�q1H��
����Kjh�<�J֐T<���0�&�R�a9�p��I������&}�Q*�k�%i���g�N�L��
��[(Tg�� �?5{���1J�r�aB�9mܕ��W�ծ�y���cU� k����L��?h�ᰶ�KLTun��Tk�I�<� ��>�Lu �VW�u�@�O^�y����+��LW��D�Q��A�Ҫs��g+��+ӑ�1����`$�^�����1��O�78����C�M��~L'�o�q0hMǮ|�V7������^��A��J���n$���PT�r�f���y2ޗ���
Pa�WeÁ�繪� �x�l�O�.O�GKb��%E�뒱dq���z���q�ޏ��6[��@���!$g�EM"-�6�`JB��&;ޠD�We��.�=��T��k膭/L>:B����xH6ň}��F;�s�{_��y��-��;��J�[%u���T�QB4o�h���ph�d��S~+���l;ߥ2��ab�.D�l����@=H��1	H�D��6/����!~��l�`���-���Ԣ,�N�}�𨲮�����i��6��M��ȡ��#(��ړ����qj���v{U��)���6^Z�[����o&��{5�P�%�to��E#�{��S�2��\�?���ߣ�q���\�J0 �$]/:]�x�S�)��;�4|��3T&��G�� ��u���1��7<H,����4~�E��Ww}�[7�]S������CܕEѸlM76��%9����ҥo9�H���{���q��p��a��5o��RL�IkGz^H}���L6�!�`3��MB`�P�9���3�$�0�(q����N�z�?8R��(:�_�xH%�7����y�[����.�n^V*�Z�k���qJ��ˢ�9 M2<x��_*:�03��:7���D�U&�~{��"������g����(|hQ��YJ���Wތ[#Q0��Z�	�B�z�O�X����W�D��f�0QF��4s��A��f��C�K��-u��/'��U��S6�o�C���sB�� L�4S��?�t�
JR{��sÃ��qI`��J0�bO@����Ge�
`=l7$�#�b�r<|��#�R ^5B�y�����PP���}Q/���#c|3�>tX@���B����RDl�x,B�kj���+���s#�-����p]�Ǖ�D5��갌�V����*�"��;�{/�����mdzE� ���d�Kkv-�-.��%M����j����	C��e�/��hLŖ���Pm!�k��	&4�,��f���$���M�>ko�Uo�ڻ �%�����W����\�}�q���$l��t�#j�8�x�Å�a��� ԓð㣑�������.SyZ����~��9k��k���#�R>") *Qr�-#x{e`��RѼ���T#�?+�H^�߫��@��lc%Ė"� s�n�,?�	�xu��ګL{��O!Ȟ Z�O���[d���sfU;��"����r�4���	5%�iĠ��=Պm��k����N�tu��(���Y�N����OXB�7�>��H;<�ܫ����0{�()��F���aZ:�8�!��	�z��mY��d��%���UŇ�RN�=��<�!S��X��;E�`��'|;o�Q���/��6��(tS��,��ٟ��N����� �̿�������֓�mĽ�=�!���q)g�A����8��t!���>Mr�t�0`�6_�ƀ��$��8D��{(��2��pP凞�鿋�R�/�0�.4	�o��;F��EY�f�dh�'�B�i7i�f��fDb�8?��biah��tn��N�]E��+��B��.���ڗT�t���OFv���fY\��	q�2����k��1WN��:��;�,vӾ򵝈X�y2$�J��k�C����ـ�VR7����+ 0D31K7���k�Ԭ|t��VŇ��97��kˍ�`��Fݦ�(�a��M�r�z�ަ���p��e"c����Yo�����p@� �p��b��{^Y���&۽��.$}�kj�
:R_Q"5�|��׾��������S�&:��ҧp��r$ox��֚�#� fs��cGZ���eR�����L�N���0��,f��sXtX�����j~�k�����Bİ`Ȍu�$��ꙺrӢO������Q�������ǹ��v��ʻ���v��� d�A�e���ARn�>8�xmn�3t��x# 5����,��ʎp��27�7�z��մ~��#���"յ�!�/BUg3}�x02^�?��2~BB�a�F��_�������å����K���a*�5y��R���|�/�B��~y~��[�(+�Br:��*���I:���#�tƚM�cvs�5������L����jD�K�2�UN�̩��۷��V_��
h�]I�u)��l�,ڭJv�����}�SB�x�Jr4ZVQ����	�� �tm�:����R�q���ր����I��ԑ}�_�;m��A�#7\��ʘ��`/�f�OH����q����-y�eE#Zs=0%�l�5�iw���*꾈ӥz�§��v=�Y�)U�e��?K6Da���rM��]&f*�-��������8\wI3��ͥO�8���H��C�j�;�n8�Nus�r�#�����\ߝ�	I*]L�� ���cP�ÛHӵ��E�_��K"��9qT��Q���n��a�>/��]{���,ƫg�g9�5�w����wez���o�t>���q��ǘ�1�hy�h���/�vӖ.h�#o��P�i�&)[j�y��n����Ev��:0+����_�φh�ے���C|Mګs�����d�s�1+��>��Ls��y��r�_�d��lX�I~C�x5kq���0�䰭����˽Y,B5�',r3KΣ�,�������.�܆8���H� ��ނv�,Ϥ�[B����v�d�+�/��+lA����E�e��%�tE��k���X+��8뇩\ ���׾8�aioS����_�5*?+���襡v`٣�t���||�cd%Ԉ^jz0Lfb@} yk�ZB�=S�SU&�x�A<:(2��Cb�� �>���V	g�=ȹ�"�̄Ԣx^�hnc؎��F�4�xO�R�}�a��@ژF�� �JJ-Ӈ�|�����Ba���A"��%t����	�'fl�7��O�yN_py��o���-�*�����I�`�>}�|Ba:g��p1�lol��V�.�H�e���W�hf�M�`���1a�ydl�-��G]���Lu�v�TP����q=�YB'�����چ���;��`�w�X΋���y�Y{B*By���&j�fFl�ب#�ç��!��M��A���_4<߸��7�"���=�؉�RS���%$8���)9��0c}m����X s�c�6��>�x���w�b��M���&�ʥ���2���&�&H�CT���E3M7d*$7u��^���� ���,M�����P5E&����y�НN�����S���gK@{`-0��iܻ
O���v�R�t�O5}�2��uS�s�������㏀؟f���c$~�TNt#;l��o�=���ji���Vٯ��B?��������߶�S���{�6?�����Jɿ�c���G��񵑸h��*��X���� �9+�#�=�5�~��ZB_��[үd�y�"�%�M��Yj�%���6�#q@&;�O�����J�K�2�*p��ɞ�O��RƜ���,����i����}�y��Ӹ%�S�U)�?�֎9I�F�Y��c�B�/S8 �� �T�\�\����B��Xtu��i�>�ɸ�Uh��|Y]Pk]��a<y^��W� �R87�^��]�QN�; -��� ~ 'ǣ;l�M�H-��6_�7"V��Gc>��S�U��o�K{}9��$�2��<Ԧ4A/|�4��y� ���ާ�9Ң�"&3����}��6�x�K��Ȅ�lLb��N��H��47�5yŚ� `B���:����nK?��O�l�]'���W�Y�"��39jv~��@��i�-|Јy��'��&i�O�cW;�>#�T������6�q����ܾp�.�w:B>�@��5e��k�U�K��3�=���Ԋ�����=�����Nu�u�X���%Ps