��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM�
Ɨ�j18a�W@H&0PoΚ|$�;Z��l�)�
q6���J��/�ݎsroEL�����Q��:J��R��/�K�&Ʃ�rރ�*nަ�O������K��o��n�꾬\�8��F5�WF���k��B�3���u�Dt�yD_���]��x? ���\[�9�5�0oK{�9�P�Z� �S�Dx{�g��Y\��"�����;�6���S��g������N�8QV0���#o}���X�9+�� ��f�R���Y�@�Ok�n���mѦf��x��ìǍ�]�9�����Π�3Ϡ�7��ۢ<�$idُ��t��1�����
N�1��_91���e*�Ev��;\�m,{�Y��l��wO��ݮV�ǚ��-0w]59ѭ�="��|�F��c�k�+kb��W4M�k��+���d���k{5��5��C��G�)KH�1k����],��`I�[ف��wrp��HO֧}�Rk�:{�*I��ā��ؒ.�xE�%&��+:-�c��j���DE�1��P"��_q���V^�$�}(/
"~7�:VL���0I��<��s���|*���y�3"Z�����NaM/�	���3'=7,����.
ڷ#���K|�X���IB1��$�f����aR��«G�|�=�O4����;���S������t��*O�!H3�ݤ� D9|}P�dv-�m	��5�	Mx���9[�S�я�X�I8|n�y"F'gH�~������fj�S��vV���l���U�����7��J���*��_�ʝ)}r�.��>r��ގs�o)�"���Դ�3�G��pÀ���%,N��lR@�y?���`�5�5�< m��*��e~Y��bu���d�$k��	ޯ"�㞇���B}{�fl������Y�,�4��}g �����h��aa�Dw�L�H��w]�h���n�q�?�m]I���hzӥ{L0a������G�|�u���"k�X}��~~*._0��Ã��,|5�L��l�o��ʝ��������;[/c���w�\�B3����3Hk c����T^&��+:d�����^6�@���)�9|D���#���Ȃb���O,#�3��eв�X��7gg�/?"�iV�PY�XɰYeZi
[pZ����p�:�X�ص�i��v����lK!S,�H5H�gH��� ܪ}t�q��_?��aŋ�
��lw����Z��K9�E�A�6v��������#-���Jw`�2�'#���i��WKL�#6��Ta�9�ǃ�n&?y�=�gg��!��Gy�a/Ci�R�`��"�VN�Fɑ�J���I:��5���W����-��X��ۏ��+�2�d2"'����	�Y�r����'q�ŁM^
��޾����B
+.�lb��:�{5�r	]���5�X�@=ҵA\f��tM(d�)��/��6��X���J)�)%X�������b�,�$���^��[>���4��Orwc�c���C.D�)�A��	�2y[��4�0�J2�DҜ�1u�ɨ�,��ZMz݌oT����hX\{=כ���Gp+��6մ��,*a���>vA|(z�y�+k/&��c�y�,�c�#�T�v;;�s8�S,x$�nѯ�1��Q��΢uy�k���v���p�cpw5w�v^����B@]ix"'��
E�����M�c�}����(Ŵ0����	c�Ha���7��Lf����})w���>x�i) �o�<������}^�׼Nv7���W_.��)o'�0�͘<��$T�4��R�Ț�N	�k���/�6:���.זʈ��&uܨ�/|���A����u�}ߑ�����t��]p�镳����A<+�p�j�S<�����J��<�$�%�t�E�o|���$��h����ߙ|&�o�����8h,:��\#��]�/�rtV���/�ׁ�M�����&����2GX��u�U{k�#�/�t�)8M},���z���w+5Rþ�����%.�v���Q2�Z#���~�J7nbX�-�z�1����
/A<�Ώ�K�"��|?�.��2LU��Ɂ(��-�*G���D�n�����9ꔑ�����nP���Ea,^n���AdqcQ����KX�U�H����CU�7u7��m#kE�&�h��f\4>�U� ����?(�,�M�Ym�:�7�10~؛=�z�X�(|roO��@N��;��r$T���_��xW�c�j���33�r�HJ��Z���ע�� ��=�C���Ly��~�(�%H�����ީ���w�˥��"|�H�j�FyS]�z��J�˥s�内��Tڻ�?M�6V�y�� s
�p��8�r�2
t�'(Е6��.Q�2˳-4����=�Tʁ��2K�(7h8,�;�å��ڨ��dߚ��k����a��>����\6�ǧcm_��~Ps2�ÑT�=��cN�}�����r���o�[�]'Y��073M[d+���:��omp�c�H�Hq�1���
�3��;sB] ��0��##�y;A}
��R�~��\�����[TN��I<�-���y� iŠ�%�_�O�	V���[�G���<�V�]�@	v(Y� ����Q$�!N����Ρ�w&������y��z��p[C��&�a���ʎ�!��x�K�U�d4�O����"=���:��g�L�&���3��ak�*@���w�E�(��A+p]|�D�x]-��b��h��k�(�0����d�%7����d��x�h_iE����q��K<������}ڶ/���Κ�N�q�
 *��)�!�*�������2����",c��hm��x�cO(uG��
�����艽/���^s�PW
]���1�˸�2�[�ĴF%i�t���nP���΂�~�@���x��	�K�[��N���?�43[\�8���^���������<Ҡq���'�)L�vSq���;�x��t���4D��]ܯ�3���J�Eyd���H�����ͬ��~�8+���[%I������b쮶����b�zݙJ9%xV]�M�!�i���R��2%�=��V�K^����7����(9�I����f#������X�R�u��kv?�v� ��T0.e����b��ң�j�3Fd����x�bO�b`�	���V)���j49�h.��R�Fژ��Z�d���[SQ�S��z��ݗe�����g'�ثB|�N?f�29D�7���m�?2t�8W�Q����٬��� 
��A_��%C�}_(�-��������x)���X�l�r���DW�]o�:b>Tʹ^'�sбo �ug_J�v����^�<s>^�g3j���G��K�;�)�J*!u�� �.;Q�uG��hz�ۛj�B��(��P����qK��8�?�[�#��	~��:i?�f�j+0�O8Q�r��7��R���-z�d(�n%�۠88ꓢ�8K����T�I!�w��T��f㮯����C���T̚�"��8�'�.����([�W��$#�n�!���5�Ǭ����e�X(�*>���YY�M\�����g�a�("��d�%ir;g=%�.Ng- �0�z���'����̖8�����W���@�D�m����h��,��F�P�?K^�_��U�ߋNۮ�}r�,<A�q���ql������HKT�O�>L��/ɶ��2t��1�c�1/����+h��kn�*���Y����'�.�w��,B�.��FNd�B)`8ާ����p'�m
�̎i��>��$�0�gſ�q��UT��N�)
�ϯ]e����^��^��*�!/�[�Tg�L��Kw��R��Q	�k.� ��e��FȮ�\]�i��~��-��(��Ҥ�C��_�#&����rO\��f���b.�ʊ��Po��H�k�F3�#��z[ �/[UX�B�;�[�����311��1FB��;ڛ%�`�˱rr��;�߿�ā���o8�R��RQG��~���u�m$V��ͯTx�]�w�n���Y,'k����Slt�y�!w`��N�C�ê"�	�j�qj��}x�<(6���2Ƴ�4߼�Rps��.�	����&X=i�jt����ak�Ea���y<���R2�*��<�b{�W->��d�h��*7Tj8��Ċ�]U�8�N��P��Bw�{a�B�+�\�wg9r�F�k�@��/~�{��E�6{ �^�����?�����XbC#!�m��K���D�{+�������O%�[ܛ0��̩�$��|
4u���x��g�D}��%&⢲�g��/��$1�?.�}*�s�2D	�/#w���U�>��n�O��K�U��l��a�~����̸)�:�]l��ms�E>��)�}�1;�1*}�м�/�6�[�Z�'(<�����AS�\F#�N�������vѬ� 5(��� ��!A�kn8Um��l$�]�1,7K�v�w_�o�J����鬫��t���N����x�R�N� ���n��0�%�ɏ�����? V���{|ѝ����
�A������}�l�{(�����	ѐ{�}$��w�[�)�}��
2F��^�^r��$��0���f
wɟQ�[C�؆FJ���W������,��$T� AՊ�	'�6��D��$��Y����D	�߻������H�h�$�\�A�i�t/&������N����!j�E��G?��xj��Q[���IPL+��=� �n�`&ݙ��ݵ���@�:���e=?��3D�!]��[�O�V��z�6V#�Q��̑U�e�,O�R�F~)�vP��8~�k�L��y��]$�y&b[��2���PZ욹��y�4L�@)>����'�#�ch����Ҭ�=�϶���q��a0i�A��VAN���6K=� �c�{ ��=��A̵�CyJi�Q�f�-��Tqj�)�2�7�W@�y�&��������wZ.~��&��>1�f=�y���N���^���U�e���9���)M�ۭ-�!s��P��}�w����8�/���4;�_ �/�����x/��������CM��[%��R'��-EF����G|��<k7 �sv�)�O��k��T�j׀p���Ռc�t�b#)�5M_Mc$���}\n�-��^Fzȝ��Ξt����~�#B���k��ꚍ���������e>T½�7S��,^�6�}�$�h�l<c���\$R�����z}�A	�j��n�=�F!M��
<�6�x�����~���I6��h�$���s����5�0Ԡ������O��|�	$��q�m�v��� ��,��Uچ���̤�����xaJ�$��ZW�2��!�iO�B��k�y�t]�$�D��}VOA��|D��G�
��z��3����	BL��.�B�_	�E`�I-�Y�x�e95ar�i�(~H���ύ"p��3���R	�(昏|Pu��s���	S5X*�O7�=��i��(>GgLG������!FR`�-�!{�AQ�A��o�3ޠ�����x�V�yk�h���U�~o���5�i���߷��Ȕ��>����Oq�Ľd��|`O�Q��x������^Id#ò9d�6�e݋��-,9v(��Ӵc��'��+s�9��ɶ$�%��q�0�.?
��]��u7G;Brqkq
�lpU_�F`׷�"����Z>�t@�B�S��c�q�Y�����9�4:�䕴߄9�ɼ�!Y���#Wx)[��Ah���?-�HA���L�^����rґ��(%�q����΃���q�~�NΰO����̮���v���tI딆���b漆>��S��x�4R*3�	�e��;G��g�dC�Ȗ�t��HT�u"j��.�ן�TJ4�$6<��~���V�bCMX+��EF��1ܪ���{S��R�3��7X;��l�g �1c�#�*X,Jg����2b�B+uu�]5�����Wl\Q�j�U
8���e+����|q��Qܓ]=S���py�7��6Hj��'�7/@p��)y��r�� {�Q%�b�x�������8 �<W�Ӯ4�y^�	5��&N�f=e�7ip��y�$��t�Z��N���ծz�|z<�BԜcC�F)ǔ�K��nkb��6��6Vf5�G�c\�[P+F�c.GA]w�+��q�����$J~j(6ψ��Ҭ�� R|��ɺC�?q4��ߴ��!�I����rW,�1z�R�=?���Uyy���H~M�1������b>D�F�w�!x�h�>��u��Lc�s��m�|���=�g�O���̸Q LpXͶb5)��0e��P��]�(�A�V	�h�$>���W�,��5�'�b?0�=&�6����Ǎ�48W�gO��|�$E��QN�F�pR7TQR�i+����Wen�ⅿ�03Ei]���[��ώ�|r*-W]�4x��/H��	��LfQ8�������v�P?����X�����0�N�nݰ(���̌���B��G�17~�#�6dg��}AҬ���{�� ��	|���D���cZB�&m�\�g㺂͏Z8?���f�;s���@���\w�^cYJq�m�˟���T]��7rh�#����<R��U���MI���i�R|!4 �_/��&JF�
����(k"Bx��>7��:K��Փ�$��|�φ��͵;��9y԰���km@��n�����q��J,��='W)R��O�Гþ3FǜJ��Ca�K�B��?8n��:��D9�	�DC�e�[3vG�Sd5G���N�qK�
�x��2~x�G��x��U�'�wV|cW�9�$;,�ɔQ��L�ۃW;h	��X�<�+�©Ov�oq&%�����{�x��IM�É⹶�(�&U�vSݗ$�zo��`�?��{��O�`5x���K������x��ݢu[���w?.6�>\�낓חJ�W�s�¦5�8r�6�~�������]����6@�%2afn3ث+���D��<���)�K�og�ϧ�.������>�Zp��ӶGVG���i�J���v�0�,v��4��Y���M�H��0I� ژ���W���).�(�#�s C��P]'3��L��ZǾ9�Z���Q��i��[O?�J�?��x����-xOi�dz��.�rEzw֒E���s<rx��,�s��))�l(%QF�d�U`a���*1�T��d���(�)�<����-�h���F�7��T-��ܫn%�{(s�eK6�O\tUZFc���1c�^-�JD?������{D�walV �����Se��`���H�Ӧ�Z(n��o{���jnnxR &�c`^EX=j��P�A�{��"�c[�f�PE�Q�{_�	���}��f>g�*]�خ���2�W1���/�������ym}M�n���l��`�I�~������꼯�yR�~�X�RzJ� �w��G�1GM�/?.�򱙽�N�.t�bg7���Gj��$�䠴��A`S�Z� B��R�� �oԱ7�g�|W�ύ���p��Bw$�ۧ���䊙70��Vdhh�իG����2>��HX��O=�88��c+C�S�#7�`�q��lT��`�%���b���U��9�}$tc���Bq�;��ŃH0]����[_�~T"�0]��A��n����B������INT��s{�.s2��i�$�|�?��X�J�Gb�3rb����T��?z�H(��褐B��̿M� �~q /�w6� �I��¿��L�u^�pC�p�؄��;(�R��\oJ,�u�m��
�����JM�Еz𕩷�����%�G�C.A�3؃-�$�.5���
:,%C������l*��)�y���p
�s�=y)Ƀ���w�[w���k��D�Z�NE��(���S� ���E	n6�L~�ד��u�j9�'��_�W>,���WKZ ĞHrk�GWc��������gI�"������1
��q�� �@��!�٠Ԯ&��ҕ����>>��	g��;�o0u腮��o\�<dռ��O�r���l�s1�Q�/����GW�0X�O^�z�M
҃�^�C �;?0�Cn�,'R)�{��ھ��5'�-uD�ÑcG+6��<��]�^��A�;u��Uf�8���?�� <3���0�#�jdf]�xǜ��8�}�DN�H��x�L
�ǟ��y-��E��Q?e4|�y�H�����5r� ���:שͦ�� ���IԬ���s�ZL?��1U����[)RR"�,z�ϓ��	�g�Z��]fP�fi,j�2��}�s'L p�Z������L40��R�G�a��O����M䭣�Z(��?Yd��fGF-&>�j};�	�a�j��<���S��*�E��ː���9��Y�@:C�ꉇ�G	�q� @7��~2�s��d��?Բ�Q�)c����A����V��}&�Sg�81騾���B�������F��X�Zx,�L�3��f6/ʈ�S޸%q]	rԛ߸�/����5x�E�_�:�OO9 �+ԣ�	��Aj�h�
Գ"ºT�3]��P��*'^
j�{��B�U%?O/��_�B��w��-h�m400NC��| � ��"O���I:�pM���IMQ�?3-p���Yʄ�2�Z>n�hs���ZX�'E���Ը&�܁�t���:�N��c~�F�O���q�F��;��?8܉���p�]��_'���Be�����HK�8tl�JiE]��m�ؿ�z��ߖg�I������$ǝP9����n��cW�R�?�B�U���v���G���}��թ���%VtN�a��� 
TBX�����d���}��]E�(	����%��Jj�}�۬c��̓�4��8d;�u���Zn��������	Lk��N�8���\v�6u��l�~ʨ3��R!��(5��{���A#|ƗO53��0��䳸���]�
�-\,���@�p�ޖQ���帕��&�����!��9�LУ���M���# ���FW�=]��s��+�گ��ziK.c�;��&���[rBv�4��=1�1s�ꨙays�N���A�ƒ?"���i��Fd|��wb[[�R��%�T�Y�N%�6h��!U�ш۴A���j��/�4b-�Ng�:�)/�������,@� ��0ṫc�';;�e���@�O �[~y�&.n�y{tZaJ��gP�=o��qɦ�����}ܲ�)�K"#��"Į�]�3��3����y����VK+�K_�����MO��-�.l`����������t�=C	ժ��]z�lM5�����ȓ{��e����r�?�!�:Ch�1�m?f�����Er��+�\�䫏~��5n�D����^j�c�6yW���d��(&�L ����0m�@_Լ)`��>��|�n�_qU?�e,W$G$����7�x!OU��m`:f%��:���&5��@�.Ql���N�u����)��m3vq&�S׋��)ѳ��J�.:�#���(I&g�$��&t|o ۟�::]�y��$DQJQ��!���%^�ǐ����y�x��Ӛp�t�pa�wt/����R?�!?1q�~���N̮�wH�Z�R�����T�	VkFc&l�l�V�y��n:�(�B7�h���Bs�B��=��0���|P�$lU��qTk,�Hm	�F�`�~�U$����D��Dr���V�%O�ڹKc�xy�J.�L���f�1~�Q},Ȇ�G�f諰X�T��ׄ��0���|��AB(\���'����=0s�ҋ"Q,-���e��_���g�
��{�]g���]ҚMײnՖ��yq���S���12���p�ʶ�Jݷף&W36{�O������k�嗥v#��cCۀ��oT�yJX�1�e�C�����El��D��{����}xq�F�%���>&�K}��-0���m��qp�|��\��i�>�=2�
�a	�T��W���4�".ǯ]��L���!��sn�霡����!e�3ڦ�r�Xd�y�rRS��v�X�d�t�A_�2���o��}���۔���F#[��{���2~���K��,��]��v�B���M����0�k~���	PXo��fdd��>a�`>�����!��8w�\T~�'Bo`D���x���·j��:"������I�k���4>~�u�/(y&q1���OBO<����I���x=�a��*mEc��C��m������k�"��h�X��_�7Xw	8���d�W0Ǥ:-��c���0��:Q�+����z��@����;\�o-:��x���)��E4���������ꈌ�M��VH�^�F�	8p��L�r��.wٜ�S�