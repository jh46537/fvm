��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a�
�Ys����'Gc�$��@	[��%S)�8� �QA�� ��GI�=�Q�%� �q��j�C�(N��.�GH�����5�5�kj��&i�&���eJԧA��}Ic�>y�R0�������t��ªo�B&c.i!b��c����N�`<�\.����6�;i�U#YO���O�tᒢ���[�j�@�S��|"����������єo���z.?Fy�]��Y�}�;�����-���8Fpr��|U~�E������k��6�72G6�EFL�ũ �c[>��(�bg#P�z5u�[�|�g1�O*��H&�6��K�	�K@�����\1�c�
�еbU��0�k�4؏��A0�k�u_v��,�J����Ϋ"R��xw���L�h(B��sSPZ�ir��d�r��y�Y,�#���ڕ�=r>�`#M9z�!i���$��(�Nn�����2hk@$pK�?�����A���I������T���ۼv���@�Ěi��%a�� #��Endޘ����>�4X��;@�è�+0��MM��:��'���}v��a��%aN��p�M񃽥�G������=�܏3�\���%��^�\����<1�����F��$�ᡍ��<(��d�Y��.��G2��dJj"&���,+D������9�x6�oc|�ȗ\a�7�-R�V�x�YԎ�����b�B�|z�L�7$>Xw�3!����kR@!�LNCNjy�M8"�y���J˟�)H��w�r��(apI���slY4>=��*3p&�IB*��7iZ�/^���>���
'dl]$l6������������'����]:*>������G��,���4�L���pB�"��P�F���00�uL�.�kG�W�Qj�W�� ��O�c�g�-��oH��>�U����ݤ�B���_�bdC	%��.���l����/!��nǲ ;��
�O����r�����9p��K�OI#�m�	�{8(e�T�����8��#26����
���N{��"#0�C3K��\��Qd:X�Ly z�Ju�z�9��q��N�`EȔ-���1�s&���̯�qL��[���h�*�s�B����ݦ��/lO��0VMW]�:Q��#�2£wX˻��V�`�̄�^ B���Vꫭ�Y`�at:q4���k���Ӄ_\��jB��N�:���7_��Qf�{ONܞB��%?�I���]>.$�a�nB=8��P�{)�"���b����C��#l����HN���⇋=��n�톕R1�A9��@��SN�h�XO����i� G�ǭt�Y��sƬe��zn<0,u;��>F����ą�.	�^��J��fK��1R���unp[���q4�	}��r
u'��t%X(&�,��POQ
{>�wҁ��N��+�Hw3u��}����#����{$7��Q}3;�v����UY�������	R}�@�܊m���j��暹�8��/��S�|�D�4P|[��ެM.�1�|n�_	�ky�����*�������m���Y�c�}�P�q$���nD��S�U�TqZ+ߕ���#K��������az%7�Lh��V��b�F���F�GnC��.z{��ͽr�kU�!փ���Y'hH�_"�`��C�i1<%$��81��p��]�n��T$ժ�����պ`�k�`|Y�����vl�����J��O.�cW%�l�M����YF'ס�Ϡ��o��AA5m�������%�r���C��������{�L6e԰	O��:���+d�gUmM	�U? �4�I�t���vo�;F��/Hx姬8f�ЗwV�H�p�EC_ƝV�p���j+���k�K��{���Z�H����f�%�A���_�y���3#�k���^Y.~�<�Ci�''�Hj��֢�� {�۰`|��B��zw?l�u�:X�Z������3*��YM���yoI4تWX�� �	YBh|�5���&<"V��x�DX���ƃg'�ğ����7;5�/�}�b��J=-ڦ����C�,��QX�.��T�'$ ��Ù���7��t���ct�o���)2�Z��{���0E�´ɶ�F�1��b\�2�h��-�>�<�cGj
�\D�8>eI�j�?	�������G�
9�Q��(q���܇=	{�N��=����`�3����v�	a�-��<�ç��O�h
ޭ�M�����c�Ni"�(g>��0G���p�b��28��]�����9;�d�[3�tɸ7e V��6aq�.�c��:JD���?V��k!��K� �CƆ��W��Z"�f�Y��~6�����M^'���f�b��yƄ'Y�lG\L�a���2���6Ȩ!8�~R��'�nAZ�HiY�8���U�w��3�j�̿�ή�v�]��Ƶ��������ܸ3�~��v�N��-��*J���Z�
3���.a�B���&��B����j�e���#�fC���B΀�s&<�.՘��$���c��5����u��֩`zD�����!���J���~��
1ڞ��5A������!?��s��/�佮�:6����I�'���"�2�-l���Nm!�Y �t��nb��ܘI{c4�]��劥�9R8��w���G���'�$GE{�/�O��E��ȗcܕc�KJ��Q��"I[:8��k=M�d}�'�q,l�GW�"�SD�O�;k��N��]�f��;��'nz�H jv�	��6�V���;�e ՗�ORr��;5;��È+c�W���=]X�ߖ;;�C�:�Se:���j�	*?%X�c:��ԁP��;{R�lv�ىWӯ�~ű�K�	�#�ol5!�

"�p�$OJ��t�L��B�Ǡ|�"w0 c{��/�������<�)
�#o��*/@Kf4��T���/��Qj���=��Ķž�+L)yFRx����-�^�'��u���ώ������*�1�����R̨��4�g��ܾ��J�e�G+�"H�,�g'���U�UTd�`��|QY�}��s�����K�k�D3SZ,�}tm�(:�WDr�W������ OF�����x���e�)J7ߗ���)�"�6���� a�����[�>�����`�9��s��6��|���i�k? i�1�mɒ��5�	^i���9��[�vE���3\�� Ԙn�6D��8tXbU˳֪�h���H hR_?rfW���%Ҕ�Rɭ��:���r�Z\��\E�jq�=ꬪ��O�k�G9���Q[9�.)su��GR�'l?�Dٽ�qlDt�%�'P�I�O��$��z1�B���9,Ps�e
�]+��s�{�<A�U����;���ܘ�����J�k X�� b����]�Q�V��^�-�5�� ��7AG�ac��E�����6������څ�ko�?�������yh|m�C�n�9 �ճ{t'��(������L~Rt�{�>7��=X^<��%�dz
�Ç�z쳱��M���m).52S�ZmB�e�o�~�E�8Q���-Q�D��4 (b���O�4��+�b$.�AJ8��7	�_�;�,�N�v��]cg���Dԝ������Ī�T��N���`��([G�ko�9�#��//�qײ��]������e��nJr�VK��m��D8;rB(���Zj�^�ܴa��[�!r��:��n�c��,�]�H��.=���cx+��&�0�t��ɹ)�W�8�C���y]��l|�i��.!A�2@"E3�5B|C�6�
� Z��E4N6;�^���SD|D�����k_d+�Fb���M�g���J�'�>1���RR���u��9�`��ӄA� �Y�k�-<�׾�j�nmA�^]��IZ�3��$������8��u��g��z� ��:
���i@���c�k�]kel�.�� D�c�H^'��QJ @����~���K����7��޻3�JQ\�w�=���Ri���ÖG|��h1)л������ ���k�Z��$D�ߖ<6�n֦�ˌ�V�=;�L�Ɨ�9�)C.X��Ћ��X�>�;������G8wl�6��˗s̀��!m#�Z���SJ��(�{�<y�>�Ǒ�%f�M4y�	?0?߳��G��.$±�S��c+;��A)>,��_x�%��&�pU/-�0'�b�݁�p��H���>iY.��K�\���A��+#6��4�>�gt���a��]�����Aθu�����<��^��(�N'DB�y�58�̡$�@e�c�Ċ%I4VB�!�9#�Z�'#�o
a?�5*�}�;�@���f��1���uA�j+;=�����\�@��JN�O��{��I�u:����.�Z���ip��@T6�=_B��~��f��:���#�i�Ϛ\��v��Y��R��s.�����wJ$2��Q�$�F��ȭ�eʡ�/4b( y/��V$�c�R@W�E�J��`�t/n\��:�W_=��7�_��6�&Bg�!�>�y�d�X�m�˧E��B���Yw%�XU�N�����u�o���� ����C���s?1dcC����7n�υD_��7�7϶��Z5}���D�f�*���i��0�����G��,��Ƕ��e8+I<Ҵ��S) 1B��%ܗ����15�3prq�v���bm/��X"p��1�thp�o�n�dats�B�P�ғ�08;�y�L��W�Ō��.�lH#cZt\�m��*�tk-��ŝق�"7nL����}v���y�x�@�����m��?�ՙi6$f��|P���c֍y�8)=�.�4{h��.qʂ���1�؛��i7�-�y�#1�G!�s��weq=i�d����d�HE�~�e�w���Ci�# Z�2��i����{ǲ\�*�E\r�F��s�261}�M�+n[�V#�^2	h?й��]�Ć=\dQ�2�H�g1 h�'����гL����
nmf��q%��6�����=������OQx���u�������A��3^G��vFق
O��pȒI�>F�_�E�?��y_���	�ȍ$�:�9����0�;Z����˾:��O��g&^}��������[!bU�<s��
ot�9�G�WTy��p{�I��pR=��t���u^�y�_�����p�Jkh�@���q� ���L,R���P�6��E�J��Mz�u�~��F�D�m�]� ��[�ۗ��'+~t��*�z�������{�y�4sY��د�++�Ac\�K���N�#^���1O@�K�p�����Ϊ ��?h;Ӕ��`ik��I��,3Cl+�A+�S�Ą��k�ȣ4Ϲ �py:��Yk`���0;�+*�U��BpG���k��q���x��k��Rdʚ���`:��9��̃�(�� e������j�����|�l��Ɗf5����ƽ҉�U iG��xNaQ�;��r����&��Ɣ��:'�k���|Y0���$��3u�o��������7I�	 ����0�ãy��7��5�̇?��~�����'Vz�o�z�2`a��+1>�gv�G�s�ؽ{0��Bc�v3W�&�� ������/?i"Z�§E�e2��W����s	�2����Rn��QL�.5�2�VD�Ǯs��(j>B�UF���e�Ud�C