��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)������ɷ$neU�f�_�`@��8�����Y�c?����ؑ�#���W۪�v��5��3f���D~a����5-�i^� ��Ȃ�kt)xA9wѴ�4擃��k���n�.KG��9o\�D�UJ<���N��rgئ�,�)~���P40�xv�툒o��'K����9%|iU`��kA���M�!��:l��ak
���8��'  g�ߋ<�{�I��-A���E�#�����#��0�"nP��~ž�?�MO`�b�cW�����J�mBj�Jh櫝���(�s�M��7�ײ6���g�w�!]c ��V`jI�\�k�O�}!� PWv3J�ݦ���d8�%�Nh�/8���e���*g&��ES�ˍ��N3}=X��-
"V'@�)>y��?�\��&��V]^��2��d�XPc7��kN�L�]�aNx�1��r���4���������<��t�f���=�	Ӊy((}`+�m��.k��8(��{��6�X~�A0J�TU�6�-�(D+E���wX�g�� �H�ۍ��q�C�5�h�iD��Og*����lLbw����ota�6����m=���USl�> ��|]����!S�䇰m+~�Gl����U-��
��p+�[U�Vk��{ȕ#�҇h��Ov]"�(��<D?Br����!n�b�ܝ�Ky"�2��w�q�y��� ����>���:	��*�����(�Cf,�^����5��`��t�L<0S�,�^i���"��5T����Q�>�svs�(�iL�#���`�Tp���2`m�7��t_����F%���vO,��kt�-���sY��?�F d4��cM����]oFW>��t�ٔ�����qA�������̈�*���:XJ��?u�ʖ�tsMF9gq�Cݺ!�k+x-B6�ik�g�U�
4��wx7�w�[�%�"�����9��܂Q�y��&��*<T��h\�('��ti�iӽI͠c>]j'�����]��K��&8�$&J��H�Qp_�}K�Az)*����Ȃ-W�O{�5@���� ����|���6n�@��8�l��7��ˤ�KXarhhy�k�>H�N�ʫc
e=�T
����i�|�P��}�H�)Î��ӟ
�P!�V~EKx_#�_P��k�S[��!c#��V����^9Kfxroх�,��Z0΅��*�-?Vq����k�]X q�����P�3K5�	�a�Ʈ�?�/�o�^b}]Ӟ��$��o�	�&�~�Ѐ�1ojnB>�!�@��&;c�{Ѧ&�AS�2�ir(����l��������fӐ?�s�8��,���m��Pd���͙�GK�HӁ�;:1/o��s�
�w-vĖf����{3�gZ�����[zJ��G����>��hQ�-�����t�)H�nu�B�jأ$�׬#á|=D��Ȓe���u�5r+��n�!���=��������fp�n��]{��]�vA0�!4!�ך���-p3��ך`=�R��Vr8���#��2�C�]6+Q^4�'���F�-�	���Oz+����0�WV�{�qt�hT���V�Ղ��k&o�&����e��$?ѣ�7 �~�ֱ�:uKSk�)B��|�uܔgb�S5W�6���-�/�mowK���[1,%|�R�m��Cmh��M�;��c�z��5x22ֶ�Qq�L�6n5%��Y��'���V� ���.��K�5�F���攒̪�T�PX����S/��a�v33Q�i�kz$D��z�:�CL'�ȦhC?�|�zv����TMF�mv	Q%��w2\�*R!����'��h]<u�/w���%�n	9�;����}�-��T�f��P�fg��f�Q�c�4*
�2�N�����_0ŵf�. �H�`2�gkF���H�ى�J���f����X�j�OR���|0���qXz"��Ҕ�ưn`�$��#å��S󬞫���(�N;���3�(�2>������8�������_O��{��$Ǘ�FE�S���	F2�֨��a��������n���b�HF3�4Bˇ�cK��"Jj[t�%�W��9��ż�lh��H�P��11�=�9լ� �/t���
�N� �[��D���R�~�����h�u����|�PQ�P����c��k���e�\D5��۱�
�0�%ߏ9��6Z��g�Yu��3�,.a���ɬ^y�2S��*�(��G��`��>m��!�ߡ���Ȟ���6b�2�� ��$g���"��i{����-���f!�o(�ە��|�AK�k���N@:�H������=�5�ږ��>��E�?���pN7��C�z@�Qdn�p��+�6K9�l&è (�h��!�{�g�!(��bhF	�6�� ��|�^9���ɕ��`oUm�,�q�~��i%�nM�3��]E�/.l����Y�9"'�����K#�&������Ά
�F!��Y���W. ���J"��������e$���Tn���|F
��z�$�<4C��űx�N�|�W�ޤ:�w�)����'�L���Լ��Q������i�RTO�� ���/.T�*6R�<�Ca���
���X�A�-�<��=�9�
�v��I0|$߹�ptv�=��7oO�󟑻�E�������
ե/��d5I؀�O\�*;�^)�Q`|6o`d�
_��wm�BCgt�g��;}@��@�������eU=�!u��`���Na,HԚ��d�Sa6q:x��E�&e��gؿFqو�}5i}�&p�F@6�����h�48�6��w���qԣ�O�˙�P�qd|��B��ƽ�/+1�g��+)O>��I���9�"&UB� 4��뭐���|��xLE8B̀�+��Y�������R9�2*(�\�C(�E�.����B��VDo��ɦ(n�Ƃ��p�IU�ț|>(q��%�2��u���ccר�Mx�|�l-���%E�PN�L�[�����[k�Hd�/"�uԇ�S�3o��lUiJ��&C�j���q�./a�z�	��#�j-�":xt�a���橔�g��c@c����Y)����Ѳ;?v[���-)g��mh������h��L�B��/�X���������`�TU�-_��A���ߚkx���HO6�g�����*h�uAk��X�3i�)�X��Dâ�T�z	�	��n�%C����v���8�8�GLdp"Z+���a�<���pzl2sI� '�y<���(qo��BC�~=�rlZ��ж��C횢��۸}�I3$|�9P���B�-���6ؿ*3��J.�A;�~K����-����e��~G���E0��A�jH��?��3�̎b��)�~��b��~��`�C�Y��+���K����Nk��V�/��5�i��\2C���.=zK�ƞ��l����Ը�(�`^�7�h`О+����pge�\��p�r���j*Y�k�׹�D�i�ZH28р�O&l#hzb'�M��án��B��5��zj���sY~ʹ��xb�hZ@A�1<�;:�~�[�J�hl�i"���Lќ��������eï3+�v{�)�������7 �j�x�A��r-W�}8b���ErL:������G��`�ZK |* Y��+���-�3w�]�DA�S�4�U�nK��7�bDz������l}�ſ�Iw�D�s&��8/�5�Nn<�dE����\@��C��.X�ë�nV��/���3$�ƈu�7����� m��`��Kq���NC��"Gx)��H�d!J��6I܌�g^bzA���E��
%4��Z/J�y}V���q����3��OX#���!�'q�3W�h(��p=5��<L�\�_�E��|�����e�]S�t�8i����R�e�9�ZSTnX�L��[ׅh�+DS�P�-��IO��Gj���(�l�i��dL��v����e0_�Ō��8uX�x�/+Ȟ��}�/�r����8*���xp6w9ĴW�1�����Kd������ߊ�m�h�}��](���[���9~�
�hWIJ����HC�ܬ����8�3t�����,��#���i�Va�
Ҍg�*>B��0Y�5D�.�3j��m_�=k�{�t6������SbAFE�fs��F��6�j�S���Ă��c��zp���E_��e�U���I���u/P)Q�,�ɕq���.S�{ӿ�,�MN%p����Z>�/}�=��)X���<��t�/��ya2�X�j��^���}ﳿ�#S�&�(p����\Z)���^��W���ޢЀ�E�.(c�{�L}�ׇ��0�̚/�;�Gq�����,��X�.�M�V�K#9�~�M��.