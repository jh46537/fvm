��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%r�H��Nx����,����oʲ�>�R�}0��+Z�Ь�i\ߩ��p�|�mAl`��-@Ӟ�1��� Z�L��SH�W2"�2�Skʇ���8��ޕG��@r;G��w�<�"�"@y��1�N�T�j,��C��P3ev��3�゠��뚷|kƠ�^�jG/XP�<ʽ�E�7c�J�{݂���3�A��,x��|��Va���rb��a.��rd�U���v^�6����=�Z���L�~��QIPR����N=�����-���gX7N��&7���6e�� ���
K(t���v�;k]�y?�cD�
6_�	M]�lFx�r]��t�fc����\�6�!^0!�8_���q�A�ǒ�u��t��6Mu{�S�	�����h%�d�(Ҿ>��'�ǈ��;]���V����0 ������*B�!rb���e%�-�����Vc���̿�=~zD�ݶ�z�M�oSO@��!t�ƌb�+%;juRYݦ ����*+q4t��)s'Z~3��^8k������U��tU��kX��[�����;s����k�f���KG΃gQ�'lJƀC?eS�`t��f���
w�Wܡ�Fu��[�k��0S��u��Uo����~|���(ΦT��o�q6!X�~����-|�H�rR�[�Gw
6�S]��ٵ��L��PC��[S�� �:*mF���ArZ2�dƙ�l�hl����'{y��1qY�r���U	s��ҿ2dnvճ�Fָ���1@Đ��`W�7�����!3�7��p��	K�0�AaTy������o�Z_@D��-����E@�P���
ӱ�g����~}rw�R�/�l��[���8��k�X�����ώ�n�iF�l���f��
�>�A^�D��ւ_�����s��]�p����q��;�1����UX�S+GU�R\ϒ_.)� �υ����J_Va��"b�����3r_�V����0g5W1
(C����X��Ee�m\��<���O��<����c2/v
 �Z���鄸<�r8�M�M<].V	�H���,q";��/�0*|(Y�������?�У��˖�g��G7$ ��5R
�x>����W��pQ2�$�5����_S�X0`���&R�ZE���k�C��@x{����4R\uAl������1(�SO,�U�����V�a�#�f|�b�2�rET�����'F�-�z�2*%tP��0{:�D�K;�l�ٻz�v����q�-��:�S[�����'�}Ԉ��F�WM f1a����aG�F|Иwi���?��e����.�K�����Ծ�3�Wu3X�7԰�&�N�/暆�Fmt'f潥H7ս�=�Xvʼ3u�(�R-}v�[I��h�.��q%?��)�DD7j>2}(��VC<z��g�i81MA�+��i�6v�[���%l�n��(�ta0F�K��oF�s�����S�^
�Y{ar����"��E��Gs!����Dy�b<܍9���)tkFe�%��h�bI8Jr�GB��of�0�ڬ؎�gg�0G	�T����v�Ô[*N�u��ō���&N�!��z
�������]��fH\}��.c��F������&ٴu�qgg���M�;@V/�Z����bgPY�hM�{��+�~>�)���Be(4��6����&�/6�<.@?Pɑ��R\.K���?#(�c�t��K�j��nF�(#��Ykr�|��+C�5���������)I^t�qLk�q�I~��]�¯�SQ����<�<S���c��26x���E�g��aFɿvC������p��V`a5��)_�?�Q�LA��2���4�83\@.�댜,�j�G��T�|w�7AE��	��w|��m��7��,�Ovi,��9�x��]٘	��]8���Vg'8Z���:��Կb>�di7e��	ũ�#ߙ�s/�&�2�o�9����*_:��dJ[��5�}��+^~�k~l��t��*xc*ܐ�0<��:�x����a��)�?@�����e�R�Z�:ϔ����N @՞�SK�m�;ʖ�d=w��[������<�M�d"�t@=rCG0�1�m��2��vƠ� �91��,���W�	�p��c�A�Uf��YueL�N9���t*�d&�����O��	\ʱ��@*�%�Bj9�~�u����p��G�s�)�gϲ6�����1���7��0 L�T��>�ã]��iᓐMx�!`����hf�KR����(�o�$����U����ؕGZ�j��0��/6��ÛM��竼�M�O�Rs��V��_���*����c��z��D�a,���Rp�X��!�_B�Ou[E�x"3	����"�W�H^��	�565)^�)����9�r����b4$J���K '��G�:�=rse�9!4`�Zy�j�2����Yӏ��x�ʆ��U����ąO�{'���jl��>=҅�8��Phm"1�@�휾�	�:E�-:Y4o%t��{j�5C�Đ7�;`��e6�4�E�Su
Y �*$�]�}|�ͫ�&�'z����p�B;-ފ˰�iQ�	
��a��-�a4�I-�z�#�Ԡ9��0k�l6�.u��5d�]���ID�{	dNT��њ4��j���Fٙ��_��*O�f?���aqB��=���|����(@��0�A�����~�<� �ԞQ��3�w�u���
DN;�>��1C扪0�4���;T���V���F"7L3�b�v 4H����~�W)+�qJ�|I�=J�u�Y�ڟOg�6���I��	w��H�m�ig�K��L#� �%��/�r��g���+��gNϧ>DQ��
�)�/T�k=oR
d�C̲V^�2%#�'ϳS�"Q�eS��+�b���@	���ߑIm5�࣓�4�e
!
�b����i=�b�n{�NIJ��~��P f���ǞP5�gEbro�P��B�fO��]���=[Ĺ��¾M٭1���5Φ ��'`ճ���(������I1]��s*}���Ͷ3c|�R��h^�W����*7��CM��������՟~�&m������`��˽;���7�:r(��KTd��JW�y�y	�[K��[�|rgؗȓĩfs��w�cw�:� �xCM�%ȳ��y�~�p��;�� =��꩖�Э���7�r~���᮲%}+>	�e�C�;6�_���$q��]b��MF�bE�3Q�`<�=��ච��S7�o��1㽩��zS��.�_�^^k�a����ZDd�mT�ד*�#( U
��:�~V\mݤXDn�~}��Mk��7� [H��z�����L�[��75SラW�,(O<3��z��R�s������T��y����1J��,*>�y]i1��1(��S�8��"d�U=�'6�$��o��Z��y������W>2� t��<��c��>�:���� h��%�(��O����큇�����>,�i}�s�̒u,�S�������Xy������hr�{(�n�c!Ҁs���X�B�@����j�G����b�2��uQ��:'��O�Ep��9#��k�y8N�Zf��tJ%q���V�VJ��'��u���]r���MI$�p�ˤ�,�"栀�_"T&UR򑖈��y�m�*�Q���e�Ѻm�G�]�\��~����w�\�W8uZ�c
��e}|9
p)PɎq-�k8�ڲR�'���`U�>ꩿ����\��oG�ħ��Wʔm�!�6�BA�s6�N2h-�Z_�%�a1xX�^1
���~~F|��`M^������P(���~ ��)-��r�T��\��_|����x	��x�^��]V�qԤb�6� i�c�C����)��}�$������w���9�2��Y�W��ϑM$��K�~1��� *=��������f���9��4���C{��ۧ��Z���Ry`Z(��ipB�߽Xۑ���1g��?M�j����E� �ಈ��ݶ-�w�Cf穞OG��J�MG�>y#�B��L�'���T&m����yu�_�Ů�_��שs��O��b@�ĝ3��'H�O04Eu_�:O�D�f2J�f��D2��sl��}#�����<�x�}$�k�PW��ͳ?	؀?�sc�AOP���@͔":j#+�F\��.k�)�)l3/�}�X8��Z�����]������F~G�*C�������վ¸��{{�F�-V|iqKO�[�? ��n�mK:>W�z��{��y��e,�JaS=
��Ⱥ�gȈ�:�m��v�4���[�]��v!%���"6�$�X&��)���'�QX��`v���[:T�̋�=��{&"h|�$-�3��!�I*�UK3�r�F�v�l=K�A7�[���[9��s����0l�+�D��nmi��L�.V������^�c3��sI.͈�7���@v�[g&�Ɓ�k���f����� ��Hs\������B�/�4�)�-�螢}pIu���t�	GL-���"�=Ө^��4WaYU��PBL�v�c-�u��B�`dB��\,o�R���|[�j�bqR���99_>�
����+�q_�wVhL���q ��ر�l���Ut)&�!]H������q��P'iΐ!��u`�oأ��AY��뿢�$����\�綪ԃ��`h�nAQ�Y��`������t�)����V)|�9�^"[���f��Ax!�2C S�'���2����W$��`� &3����n����H��hǇ�J�S�D�.1�X=M ���!��>[��=��:�����vhBT��V�7�E*���(l�p�l�&���F�=���wQ���k:|\�.��dsN���߽߯Wi��VG����9���eq�e"��ݮ��~��ySf<�䕎%�M��Z` x:�Ú���Z�ܡ>�4w3 +wF21�64�u-����1I��8��2�s��tjD���$��?����J-���+�keE>	��o���d��8M�ġ�>�I����.�qi��&�ͦ�:l�T�n�u?�tQU���PO�[���>���N//��a)�U�Yw� c�������9?|�&5�O��|�F!�Y��ri$w�5�*pp�f��3�2�.���d�M���Y56��4�J��8��a��O�y�^�@�" ��٪f�wyS�'t�N�<~%�����..�i.�RR}�Ma	�k%S�_���� D%<9���S��ֱ�b@�;L���
�+�~�
�<��g��'<�'U��fm7~ ؊�4�����0w��~dC%M`s�9�H�_��y�Yw &՝���#�6x�)|s{>F�U�	��Al� ��NϢ�hQ�d�r;+��d��!dԁ���f~��&L��x:?�Қ�bS��龳S�
Q-2b([��d�Jz�u�&��G��M��ߛ.��o�6��q	�׵���&|*�[P<�.��{i�������i?s��k�u6�l�&0��?��=��_͎����{(jO��p��d/<�c�3D����)�H��kA�����>�sY	6<||��9�$å��ֻ��Xq������yj���{��B�ŋ�c� �O�	<��"�A�]�MG�f���pl���_}��T���`F����3Q���g���1�:��<S���Û�5�j,��t�I��?ig]�~���_�i� 3 ���r����Ρ�|p��?�-�P�+Ti͕�M_1o�W�m/���V�ۏ�}PE��	����K
J0=�K�b�F>b��	�5���t�{G �Oc�j~�
��4�ר��K2��䘀��է���B��.�����[�Ih��2��5�^9Bq���)���C�����D�	���
���O�aClL���HmqpM+:�B�%��Q3
)��wO�^:� >����<�0F��tB��x�T���e}�ށ&�ϴ� L�o"e�惌���8��,��A�J����@:$-F�5�^�Px�a���� )����F�[2��(Mڮ4]q�����o+Q��$��!Z�z>i�_0����h������]�}��Z��M1���g��#ր�������XN�2��m�,n�M��hmͦ�2�TbLڞD�IK�)ܸw��}��4���S�A�Eh\�&�n��y�z�ˣMd���� i}��ӄ2�߃�9��g�ҔJ*�-i�W��B�.έA�e�'r����>z��/%HO���2N���Q%��E8���"-�!�{+���B�`�S"RS-E o����L����rS�X^��t��ov!����?J���j��Ղh�Y1��⫫�K��Jl�6}<�a��0�MY��5q�R����	~ �]J��F�G��-�B�����ӵК�S��f����z�,+�RQ�xp�h�}�Ő`�b�>�9�Ԇ"Zt��"�E?>��7T�Yͭ�o��O� 5�B �Ơ��l���`�{�E�8�w���m&z��H�q����|,�Aj������v���摜�YP�;	PZ?���68���,��;.�9�	2��/я��3�+D�1E;�!���%�sb��
@��X� 'HE�P���$�Aw�'���A�����0��L���96�	�7;�ũ���=)�W�� ^)7�_�O�U�K��"{ 4oEgu���}6�Q�t���o�K�2A����^oH����n8��
U4.�#K��)-k+�XsϟƧ�R0�lR��X�Ň�l�$�׋����S�c��.T�j:�D=�� t�#��OZ�a��t��K��U�&����Yx�ͭf�vjP*��&ȴ��)z�)��"g���5 �K#L�݁/�6l�� r��>���R�� ���t�zޮ��S�Zp��] <8���ڑ�M�.nY�R��2��yR$ږ�/�r@ B$��o��bu��飺�Z��/;�U��}5Eu�ߚ�GW����dj��Ͷ�[��.tvd����5�o��{��"n�~`��!k��/k� a?k�Kw}�;�P��ȥ�G��`�g���E�4;r,���@8����(#���jv�m�Ħ5ax!Y���u��/%��s� |a�}�@;����`�h�R~]��6k�|���>�g��&��1����ia�'c�t$��X`F��O�|Q4�`�Umυ՞B��h��\b�y4&���@蒃�#�=�z��\s������xƋ�����aws�l�g9�u]ZK'����Pb*��s�1C��u����xR�?ah��8�,�:X�ǭ�7�f�&ϚՓ`7i�D�1
��)U~�ԱVն�XF����(4��Z|ɀO�%������x<S��=V}ZsM����	.��n��HʶL��-��I�X	і���	�}�EC�#��#� N	�%�8LJ$^�Ef������F��;�0����Y�d<Uz��߁C��N"»�5/΄�wR�C���ң4BƻM�z�[6v8jRMR^��ɤ���&S��Mz���b����̕��c�!�U�D���S} ��ū}:~�su��+s=6Q�yy���IHNu͂*��G�폥��^�'��뜓#��-�`��@-�^�Dn%�v�#��G�'ʖ\�`�B�띃�-�Uu��/omF�u�F�Qޕ-w�q��`��Я�x�Zp�[N&�$�9�ڊ�ڜ�0w�������ym�z�W��r~90�r�/�JǮYe��[���D��m�{��!�������?�)�5� ?x��h���|�)Y�q-0���8�������pޠ���)��:���\���>�z��-D}Ue�������( �rX[�hG�����g>ӵP��$2���~���`��`+�>��8�';l�m�j�p�"��`/$��r��ƣF"5ң��ѥTc�_��`�u��\ŝG�^��y��&c��s��+�K�����pv &ׄK��u�e�3�3e�Bg�K�[�f�~�?>�1��g3����Š+y�y�����f79S���a�۽g���P�I8�/N�Դ����l�8��1�F�(̊����;i�+���o��L&���j/���V���"���]���C� ���2�5��gXk׮������~0���&�y�a������ك�kũ=�_�x�Ք��4�t@o�B�����P�S���DjM���`eZK� ��K��.�����-U�я+22n�)`�d�*i�jE2\���g�D{J�ȃ��O�f��m�)K����J���D�K�7GE�l�KR����g�#=9����T���#6L1 �wMu��N�a����"����?��ȍ�4�kA����M#f�);��<���ȶ]z��i���3x���CW�2bQ&��έ�8F�9H�oq?�Be�h�/x�-f��KsI��t�8��l�u��\Ҷ�KB���;�x-�����u���YA� ψ�s�E�#Ko� %m1�$��uӆ!��@����nz4΍N���>(lwm�"GF�#E����l(�V/^eU�>�y9^��n�Tݹ������V�^��P�PQ�ׄ$�u�b����[�3�v##!M(�s�BjR�Ld�A;�Dk[V����)��P�Jd6}�y�̃#z��*|��%�~𵖛V��*�J���j��c5�k��X𩍕�ʠ�u��,��Ō<�[.���V�����sz��
�A˵��i2�3
�EH�z9��Xٓ&�:�3�bU&�e&�Q1��cA���~a`Q�]�2���~H5����`«ٰR� Y.7J<�j�5.��b?����)�����B��qN�;~%Y[,�j�uv�A�u��K7�)�x�OF��&�#�Y�2�;A��ۧ�3�^�W/��4m�RS���;�۷���Nك 	'����ȍ�>l��d����A�jX�ʡL�-�o\܍4ZS;V�ȿ;����;�����9�^W+7��-�����Z��%"K�,�TS]��
O.I�3r�+:�yTH�X5�9�{Wt ��pl^�������׈���� -39P�W�XDAңF7��|����s��� �G��{�Xp�L��5�4�Zf�3ߎJAݷz��ɪ�x�}�9� D�~%fye���.���P���/2�S�t���zrw�����_��O��
����䄞FR`[/�\P�+(��ۚ4^[��x��N��(�ų�c����}W��xE��e�f��r�Z����rѨNюu��H����w8��C���{�DlD��o���	�G�l��t_��>��3��_�C|�eq��R!��X/ZVh�I �܌?����J� ]���>�� ��r��m�������Z� B���!*�������s ������'] Rq��Z̦u�J��S�
�v�$��	x3��Qk�O"�Hܾ��Z`@ss�޴��z�%R�~�i%�&S�q�yd����=	�K��TN� Z��=�
���&Ϙ����ˈ�[����_���}�����ݟ�w�u�����ܥ�������w�-�A�dE�Frh�a�� *,�_����C�L�ԣNK���hn4�7ςӢ�w��Hd̗��g��^�{)�����tY��YԌ�<�4�.X�m�`˞�*��؂k���ȣ�=bҟ�Lv������"�;�FOi�;!i�^zB�^>S���&j-�́����AC��烖���=�G��# �U��Ozw�X������G���ݠy��������D.H��7�7j|E���Ŷ6VR�}�	�G}<F,k&�\�Bѧ�G����[�3ڞ��V�7u��J̐o�[�\��h���J�3_��83���������N�3�:��F�|�'m ��o�<9�q�-x�����PX���|b9]�L�-���n>�K?U��x�JI��͂[��X;Z]�h�'�P��xo<
N�g�HHI}��aXT�q�b}��|���g;�.	�@z��'¥�u�I�y��8���m;� A��Q�\g<�$�Ut�!����dX�s��,>��w)t!�ఌ���N���Y�O7t�^��~� �XK<�8�(��Ӱ�#�/^J�deY�7����A������5⫝�������a-[?��;Պ�Jg��y�Ć�Q �L��iA9���gq��^[.�S�\]L6��e�%�X�5hb��6�c�^�f����MIb�=���?�M8��u�a\`�1r�,�_~�c�J����t_�\�������$��G�Y�q�]�K� ��l^>c?dbI�C�p�˺L�ڌEJ��f�۸Y������i��M=D�
�� (�ƨR���[�;���
��큱F�SF+��T�0n"R�84%����)+]���$��}b4��	a���qՋ.?�<Zǅ����32�.3�<)��X�0��}m�<Lj�����38��OٕQ� ��l_<]�PC��[��Q��{���ë;���E�FoD���\r����[�l�fį��Ē�����yd���d�YO��|ی�9.�a�H��83P��I����D5��L.,�q��$����#���E��U4@��9S��F�ٳ��*����98�0�"��E��Y=y0��^t��	���v����P�f�f�/i_�v9��-������a6G=��9��Q1��4c�Ѫ��i���gt� �������'���H\
��LH������A�&�{+!�"��!�y����n��z�Ѱ��)g�t�z�xa���,��¡�ȒtR��NȖ9V�h����Ґ�lI^I���=o+PrE�%�w��CpZ����U�����G�,k����GR;���Sl��_u
���̑���jP�bNĝF6���`J�^���9Ɣc /3�Y��a1�"x�k�M ̾���$C0�Q���g
ݑn�d+#
�Tώ%���,�g�N��%xiK��Z�a�t���-�^NJ���]$�Vta�D�nx��/��r�{r����/m�<���N^Ooj���7�A���U�{&>E�Ï���攑�O���.�5eM �L�7~�	FTjdp����nnH�Y�YN$k��ޡ@�Ȃ�:!�T�w"J5+q,��ˮ�rȠ�x�Ѐ�+3�>
��5��vƔ��{�ߞ�j��
N��%��%��l ������x�������3�4��˔�"�ӭH��QU?�v@�5�-�y5C����C1�jE6n�����y�tFc��r�OL��8"sF�����9�n�