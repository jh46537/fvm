// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dZ22ocGN5ZHlOn86KOSrkre5QoV0HnWqoR/gRcSdq81nNV+UnTsE5UXdtQ8tnT1I
YJz/0jocc69nLHd9d0h7lbW1mN7zrV3gOchCiubk9NlbBGmLLOhwjLH42Wb3Eji4
mHlGbhqsh3FyxIqXocyiEIPVAy4bQkOapbAcsmTEtak=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 23952)
byC/YGX0e1uMn6pJqt8v7V0mNMk2dj4Xv0HnpL/HwuRtLjvOVkmoEecFzYbjjBOt
H3bBTVQ3qn7XnvhbDFbDMfrcy/jTeotp8WgMNL9bMDAgQGi+cPAQ/2VB/CSyRk1/
GNP6Q0mgygQWjHdbmbwZ3UG2nW9WJ3FwTAr5iuhmSiDfV280biQUdM0VQjE7c/yF
kRmW7zLOtu85HTPXbX/UDuD8xb4c3KMgHdXgoq9EPT0TDtFcAjdHj9tu5xZWRpDb
Rwb9vOsM1Q74uzDReF41JH0lDXs8sTy5L+Uo8b+EJjBA7s6djuMO1GxFlETB0L9/
vAI292Yvde8cRFiHYEYho2RkdlpiEUDALaK50W2ybf5Ejc7iUenEopVjkhlIPVh/
bkdBKT4N4Ef/UDsNF+0s+raeeNxSQeRkwsqFJwOWNJpTEY6PJKNPuc97aPWcGGsh
3vtFxsf1mrMnSfNCAkAE11o2M+oXF94mzZlmKDOLY78lSkuC4u1B77WWsp+JbCwQ
tmfLbJdHU4LCYs0HWuDZvgv8T708zo5CltqLYGtTAlObtSRGxGvMyafRxU8FXZkQ
fJN5KB8nA1bjkz96NkpFoF5auWQy2/lZ2HWo5bPXCMlQY4mFVqDFnr/+IY/hG31i
CX6SEhVopSIqqBTlpNTLRSL7fcwSJzTt3wEPejn5oo3++XrR/90CMZ0xUbzNKTxO
0wrOSScWYHx4HA7JHMnUWJBS0BcCwe/hJiG9Hcxd/OnsXTnxxV26SXcrIf6+ciRF
u7VM9y672PvYgU2UoI5DrDgV9nZ/PBUaj1hkCg9c7giqMpREoakZytgwQJ3R/jHn
ahDpYtt2jSlhEIUplRbSdEt44AvdFjYTUKLdikz+kYR2pqg12EnpUN6hA1TvUCXP
1iFxJ5wW5ZJCdwDDMoX0NoHVPHYgv9RQPwfASury3LoCUBltTWeaYZkEVR2Qj7bQ
XqZFWACTTDBerT8dr+qwDWrSoDKV0523GGCqb+0pGzgJnm7zKCA0F3BvDBVVbnyy
Q++LaGziP/Qn216Ey0/B9u4FOLKfU44HJSXE9jN2b2setViJjGj1Lnr8ftkC2pmb
r3DSoYB+JCfIJ3U1vbG9h3QhUMY2LA+iFLqEUpb45W43aAx42DUR8IpnspVsUt5n
FBRgRtWwNfPQnA1qwLv59DCf+o5VqH6EVZRlWMFbD60B8a+JETlRrHKBwBaRofrC
G+BXf3/3UOpkeKjfky6VCY+A3frw/Aok1r074K4fSYerE7xxwBMXVgm8G2PIForF
+iEX6Np79Th4/KZ2A3aMplZ6bRXj4XyTWGUqDa/gnQymDx5EqMlhaV4vmXMRH+nI
7/qBamG6zUd5sZO71cz6VjAwv7m/CCFljhfL7xVQOC0xVIeykSQG6wMjio993uA2
hJg4OlKUXkvZxPs9jv7nKFzu2myPiBKJHVj9R9R6q1LNyNa+9Jp8o/0evDBKOic1
8jQkgEtc4b7AJlccBU6jsyWcBpqsTnFTt27+8W3DkkFkuH/Qn20N8VA7XkWFwbjy
GIENVB23I+cX0FHMcxc0SvWnQ/K1OM1KqHW1fXYakG+Q4n9f88oW9R6KOyWw0Gsm
8VoM1rAJq6qMSRGU6nQ2lHN7ij8emu2jaKaL/TrXwGx2tnCSc+MfTCpyQIH/CC7i
YZpE0R9IkKB/mAJ0FrKvEWahNjrzrHaVBnJOrcJVwzxmWBg1P6tFGPBdBVuzmxuO
DTZRzCj7KjQJ+PClt1miOtnGId+zWveawe/z81fUnTPhkegKA2gdqgf3M7OADQ+2
rbpnKGBmtSAeKQgKSXyYxXvarwTSlmA1ahV9G2fE4uCz5OAjUR1h8zZUts0p2Gxt
6I6rvoQMQVSUfZ9yEV1Uwh2CXazdZS7INKu7kB968KFw2PqaWRCSf3pzj398SNTr
oRZDBZkzemg85SXErOwBHjG86qaUl0KMcA5z1fWlMtbGdRZQnk2BSxXZ5n33k8sT
q0Zed8lU41LYXd3Be9W8olD+dAWnk7Dr2DPdOPu/ugrLuLD7t1i4K4+VvsjBRH8k
Jutj8j4ryjwrzDtGZF4ARXkNH9yFEv8zHmY9MSnCf5w6DR2LM+DV/zEyT8mZJX9Y
UOqHvusqqZfeO/HZNQRaM7C1y/WFiWI6QgyREpQm4ka6cfBl3zAcqEPryd0PlsFr
T5WDYeDbRKDFxJr+w0OcH/OnHiU8Ztao2d0LHDJ9+60vrZaVMz59/KFyvXIA1IP9
AE6ctU0KYJvS4z0IB8COOXFNzOyyJbmaQMe/72IolxewZdXwnFoabSOGUgLrG8np
AC6T1nVsTLYNG53t4RznmiMhTDMociRbs1D8fgvv5GWXUfnbMV0Okn8zQVtPGtsR
vActfE9mFdaZjrR52GjHtxeRh8oos/gGp7AFSqvCJeKJU7lnG/sMbRFuSk/Q6Y8e
ZYt+T+dit3xS5a6fITnmxSwgF6Wj83G+IaoKDf2Agj8KxpgE2p99FpKkqC3on8nq
MD6fjvjL98fVFxs7d4QrBPrdpdYidXG4AFc7DaF7gWeVqasqRCOBo3vMjEtCnkiC
SKeJxm9NbKQEt2TIuXvoWtmI0VKGq8mogk7oen5iO3WYvCL/nk6BPUDhzOsJeiHO
atWg/KzHlahCqeOAcaGTKFG3H0q7iQqbHCZvF1gsNZy/t1NXVmkHvg/gpmBEvZnO
c1E0RJ/ukFA8ZvH10gNqL95jLWmnKVlGwDvPyxpGkI0+JDEhSgKH6gsFanu+tzE5
aVxd/Nj/BaEdS7+mUEg3s2q2NOY5rTDWGqm4OU/qkUOv1leNTiMPiF82mMRVivMg
BXhKiYQTrT5AE2B7m4vvJrQKcGdTMYEQq03My4F2wcITXjJewCK7yr0yW/1Hbzjs
wJtpny6vdv+kG+lw/BMvOtDgKW/QxTl3Q3lH8rtxwviKCdRrRCFrettRHgDedxYY
0ssCJdI0B/ni6zpUBsjp/wi/yqS5AaXNTnpJAdYPkdeXndB6mVEPeeoXk8dEsrsv
Odwn/7AJ9aVImug8x4rNlX0XxUtL618FkgiwuLQswutpTAoyHdR1KDS8rfBnYDOO
Bt17JHiKtIjbvolMzOz2z+wWJFJbVL9MhH1+J9c0pg8xZktCBSzD6WjR6wUuFaXK
FZtcCN7jrUv5TC4/o85VQO+VCOA9NfmOVU7OANoHex8KvInUn01qmD1Aurjxe5jS
NUhWb3GY8Lv6SQevS7oSfy6TqdCtPV0aI/L1Qe0JeEwbv4XtojEeM2QKYD8EdRy8
1V+3xIIJKP2gC7zsnwAph4XQ2j31nhHFIw6n3aeApFioEG0Q17cjaCQP5a7hysXJ
2qZUxcocCAr9J3Lc2aA1mF6J4PhwRS/Z2YQAZ8nMkv3GbJ+rlkamX03W5sH6CO8h
7z0Acx+Fb2NP8mDn8aI/vvgZpNjGsNmix6v41Pg0C55OkVCMWjIxXdnLyTvZPzkK
5srPeChtxgAgDM27LFG+F4SouFbUkSF3goKnujIA9IvT2soYgxBI8IdFm4Fk6qnP
M801ie5XTkmt6g7Qd4G1gUFU53F2DsdMmOHLTnIKhrISUTYWnJFvNdMfS2dNarLa
uKyazh9xohHwThEZi2N/y/zmZ/h7n/Ms7VARZccboEya6Few/1xGutXGoGmE7qI5
99SbUvYc9/gdC9B2f3d3kJeU2ZZbwP/PpPZD8pQOdQStWUAtaLLeYFlzQ7q517RA
+HQSJaqlWuBw6Y7/H6mNCwUTtLtD3Gv6mGde2aIlNrn4E/ZRxUKK6bD1KYikLWvU
LLjBaC1h53h6ni+KNMZ7YS4r3LzIPqZ5NNlBHFI8+4Pxvznxg4P5ZCdnNim0jomj
9HDLsqws1tBOgK1utct0q1VVHnXl+C5rhim8jyP1qPrsA7uCukXK6Rk9wfHoKqFz
Vgm4JOKWhPFksnuYVSzyNp+0gkkVmQlW0QsVl8E2t3h0DnSP5c6mpunKQAjN+J1P
9Ky7zDLCnku9oZMOdU/jouOPZy6XhD18/i7WcJVXyZr7MRKtLLUmcvzEzjFQqg4G
6G95NtcVG/tLjOniT2nU+RoXy7PRBKPtnVRn0OdwXkvQj1Rre5t7gVRNqswsmwN5
rjS0LLhOlP1LNI8pvu7rFSwqgx0eIUeKBruKRh+vk32nLRJF/jIFKHyUJ2zkYH2X
p903yQ98zwTT3Wpw6UrN/YA3UjIwLN+KGCc6avRtJ4StUxPiJ3t5X3rY2tNkZQS1
uOgRAooq/GYYsblJd9WV0AsKPIbnw20kiDw3ydUrKoG6Y23scxI8XLJ258LKZEvx
osS3o7oy+Iina3/rQSpbT2/CpTAo6j3rETfmF3rza5E1CApxEk/XX2NzG2N8Ftha
5kBchXQnaFL7WzxBJ9wFspsFOWEcIdzI2cOaZKUTvwKAZ0z9kQsbH4Un7d5fVUK9
1NvUg9UuV2L0ozh4IeLvB3RQz5mwCqw8uDR2ORGIeX+Robm+naPJ54+S8WZw2rZ3
gGFQt0W5AGhF1tPQ5nP90OH58GR+x/EbK5L8BnYPJBxRsDmbobmd4pPfxj9jgBKu
9Y/4bf+/DL6ICv6KTHim/gSFocUbDUjDzsszxjceRINWJ1ysWAvag+AbTWIfmjqC
K3xdBf+zcYJf/r6TgWTYH8hdkaPu61J8pxtcFgRzUK8WFXVBmBpveHXzT3Laq4Au
mJYFU7Y1Eph/J+R/lAObWL/r2YZau/UeqE3c29VIHD+CU+DY+AyxQMsghv7ZDTX6
80zS8u0JdHRSrq7PPZPdU9v2z2nqTvDPMbeeZmUye6n0I0D2F7hYReKmXCGo3ytM
UgqUl8J0GwdpLK53dpb6gBCgXSUJxy5E43MqiY/HSA0sWGE1bT6TOi7hdNa4t4D0
yX0Kua6Z7vD5gYDAE7qBbSqF1iy70Py4YoOqiC+MjMAUa9z91/TBhjmOte9nxaN1
Fg6ES5TmiW2EKu2FLe2EVhLnw4wtGnCVeUBdnKBVHDcEnHof2BvS92ujfCUgROuB
ZTKYPpbu4NZSfyHxM2ExiGw53T7KX/RChkQYISQubUSirkOs43sbTthR/aEUDnTy
oEeNluOuJcmGG5iFVS7aD7FiGZhqNMkEth+2gr2IyUQqE2IV1T9r/jGYJJGmwBoS
giJ34PzKTqKqASsXj+mB9uyWTzxvvKC1oqbsyvU74To7V5aPgYdkgZ6QByxg3vFv
qKGtBMEE3i7CgSmiByMMo2EXW9iDGEhUZ+zQA6o32HUe0BG2IMSz4fE77D0TIoaD
ZfaBqKMr4PrwdzIjnQo1IpplJ6I2FSqnmfM6fghKoUM2c8SxNoO5UMH2upAX4Bde
EdE6c30V6+JM7Lr7wJWnQ5HmBqo7U3AXsyF+bRtJjhnRnFFGogrA7R2RCh7Cj1II
1c9xp4ahz5zy0r0GJsWPu0lAMz0YbAHU1kyXEcxfHY4NpdoEIhXwC5bzlPlmSCRE
WLlcwSXnGAGxVhPRg6FvmxrqN4r/Y6e+ZIb/sbcMZOWlZLyOi1in8vWN6uBlbFmd
BvOwcNL5RZY42L4SZ3YIwugICM4+wjwxPbfNZsmaVddCbJx5ZRck5P4jXTam+Qj6
Di+0SFdV5prWvp7XECVbc+Oku40dRH6RQWomeQ069fOIwEv4EVXWnfsLon3Ih5v3
3XZY40hqvWVsoV+aZV1KAGk8lAYwXX/tmVSqoDGCsLxrxfMdrtU/Rwphdiwj0ZfZ
ECRX9PkI9zErXzmnktAN8L7EtU8ijcLfcNduz92+DidbCwGxY4oOLdCiJFsyfv2C
zG0Fa8Uacca++akOZaPS+J4iIBW4PmyljtRhXmidrovcBBOe/oWsx9KsR3PyigZ7
/NtgK4ku7Q+sGLVzV5mUvknyIpPiY7oVMV1IgI0eb9yuJIWgB1oSbcStc2bQjRQo
5pK5A7cY5PqHvvZPutf6k+3eAIcaWwcRZhlhJco8hDSl+AIz0tkAUnGnSRn7zOwD
TE1Fy6ovb5IkI+CA3kq7+bTJJQJ12rf3qGmcfJBwze72E0VpkeMt/aUgzFwVLWXs
FxhIYYhqlZILoLSqOtlDyM8UYgwKDjnZhIAs7ZtusKUOSMPOLjl8cOW/pc9jpfR3
j2m0u6jhLnrC6dSYQ9K4QaLRiSM17GqSQFjfVLgBA9E93tNXMTWVvRcdcr+BwtQF
KYRhYB2wvTUuDNkPF4FIFl1Fpn6z0n/WYROrSyrhWNyoO8micAXVffhVYCLVsTmo
76ZtLMeVQp/H34BWNyPa1FAGe7HCkxVQ4lPBYp0soSOqvBGPu6O/6F7/Z2CDisIq
UcBqO7evPZ6GMrnFW+mkGiK6oYCgB+Skz2nw0dl+nOST6VOHH8ndRe0d6B1O1k/x
OFjbBq4FCIOrgGvoMeW6itgCpb54QdK4Yc7CSaCyKw+XIpv74fq7uwYG6TAEVkOW
KipAOFwn/YPrwLQNSdyfqZSPvcfW+3rS9tY0ztolfnXF7bSNB61RCljNvcd4eyH2
7vriHkET4W0vUZh9GkF0vg072GEeWvI2PrwFE5rkNDYQDHIg7sbLu2A8MuQFpYha
aRxbBCvx1xEifFt1rGb4XGgHpZbGNqU0vU4nYeZNsGtCqhNttd5aExaoOs2njov0
KyCSdvlbBULSV2+XUA0TUCuZEIzdCutsFW+K5vSSMSxcKkk7OU+bdTgJXQ1J8rCz
LktXJHvP0uPt45aKM6Xq5opVZyauBTL6Hv+XDbe+sO55mZQ2pZyCMV2wMTMMnzqI
I/cW+SUnJplXe8jKM92iCJmumItERz3DUacarmiNXQ8XQwugpV/GT8K2WMoLvlsr
Lu3zqrJ1r4DIkL68cNxOYsjkZwp6L/95XYdVeZABzjo1LGA5+gex7ey6wZyxICWP
bf9GnUO/PPjmnTVK9NbClml/MyHjnV8CTutGRD/keiVnNzqcQpXr6VyIDgaLMrsJ
UOhYySbEexHWHKA8MxsfxLP1os6EoTQP7I9HwHY/4immlL5v2HENl7MMWIwKsxeF
mFdDjWXnc1XrPq8omiy0epD/3RX2jwpbrgv5Ij/vFCBvxJi+X3MaXxDfMFxYhKTi
sR/qPoxPL167r/z2ouVukgyzpsv6ErUbrD0iDIxPQOwgYkONcYRdKGZ0zudVRMdN
kHEYd/DxARH1UtkZxF3a5b0pdILOvLnFlyuJgtJNxE+6mHKQqErL0ueDtd6OGxiX
QMCo4QSOJ02yy38Clmyukelenouyqym+/BTQIYGcUwsMut/Oz/6ABCFFANlN94m4
9hJy6jNbMKc85DrxXjp29AnCLWsid1iKEswC8+4M2edNtQE/M6wrKaMNk3w+qSef
ikQADxuwo9RQvjShwjh4dTEXDGtQyHpe7RTrN2iCeNicP5nEEU/99/blnj1/c+rH
TOjJY79fCRrIsBsiiZ9p1/sLN2TSlHfmd21ySnjJYcHHWKx8gkc6gmWw4MYilbLe
nmdPQhGN6IzE3kGbdIFLfR3rGPI58vJ85gSnr5TDeUo5k1/rXqrtw/LP+WodjNyF
0uoo1jLX3dDLrKRxgaDGTDaGQnEKRNu5ShpJabnPBra1syik/wjj7dVzFYfQqBvk
e++EzhXJMcT+yZsWeJWBIaIDWt6f0MFi5UW/I8DDyXPjLOOuyHMUnaiADQt0yKTv
pWX121LVMxj60f5yZMpZaYlB/cZJ6Vb5IxCVuaXcBBojG8CI19eQwCf/jgw1u1xY
a5F1kGjveCM/cc94o69leW+ZpdSK6XSz30OMjAxH8vTJGgKPpnpC+XHr8/rZR2Mi
JuGbAnNROtHekij/Dnrum/Gx08cTJNDTJeyJedJYKe07SAnm9E+K8XNljgyeymc+
u2FrpEMPmRmGCXmgem4rmIlL5ym2rEnl+0QiS4FDUzYf7w94mvkIlqO7WUmmWAKU
t8inicQI+a5dDMx3srcK9GS0f2jGZgKLHemZ4TJRYiCJUmc9Ts6qG48ZUGfjqcNz
A++7BfZJcFWiarP7Howh9Td4E9/R2+Of0n+lLlQ4Lq6zO4kF/hAaohghHYYfCgNx
v4xuQNLWnrXqxbuo+thox4d/4MV8TXSkVHk5vZUv+3Q8RJ0jGA3BabXuZIHRqcSs
w6UsNARuXTU6n+DC9xror5DGzvw8FKfesajoH2/K8/J/0isJn/nALg9g/M+s4zCE
EEjjIrPwqt5bST/nH5HSAB0yF0E9bOIWzUi25IaPs2wKkKk3oQhj8HokuE5JHHjt
i473TSQSwR0J43Y3f1BdbJ5aT4KrPGS7FKJXNrycQzjfAudJZDMJ+s9iFs7EGOf5
hJUwlmGdwk2HBQpyypjih4WHiR8YH2hn1tk+35cfUm2136KhzIkM1qz5Qp+LcMdH
5TH0dbb2dTe4GInqOSNIAuUHNyULYtC/F3Ay4n1xi5fZRQkj04bOrI0ILpPhLrZ7
Kj6WRXtcqYLHH+PS26n0aIMWa6c/bdsg4jDkDI4fXQGtpoAJkRodS+TUuWvSP6C5
V+v146ztk8HpoY2s2nes58/Pc1oRQNwBAp2jl0Y1tkr+TLcxXbNxhszNmrAhXncv
W9dQ1GHO+sCfp5w36pHqpgCjbUf/fcLDUlwsLEASOyB89YeVceRlUu+cZ/3Qfjku
Xgp4PWyXYIJ8vvsJ9SlkIorOX6yeVRjZcpQnuwu0OCKslXV+2MdC9JtB29WOYi3b
R03/pwWdqdA8y5QIGoyQjQJtOXmNxrIylGhJ1BPu2Nrf0vOYPksjJc8vninhjZz9
pbonH6jENYBahm7mzEmctn2WkhVsG/HoIiRoFv6g/xoc9ZVN9xwpYkIgIy3E0sjp
jAordI13451htWCPhJ8vCrcBqOnp1+rB53t2CEu1JRvTCqOvignY5CMDBHymyaGk
WHlZRhqoq+HuZIswseQGcXMFjhmypjF2UJvYOYEvBoPUMW4hURGCh2rZDd0oWNE8
+4iS2zmGK2IWTaqsFfsiRU1RQZcaAVu1toV13Zukw9CUSGUzgWwljC2BlEMkLDQj
WszYZqBTrhXxsaxQFpun2FCzfktuFE5NbLefVZLj1mMb382Qw6Jt6QKSIIHi25D7
CjI9GBoanuR/X2k8Hq/gIway0Kf+6gDamEoFPVNzT8Zhe/cI5+J2I7TN9oz0qUjd
2iDJpHwCwia79cwztWjzKjBTcgeAW+d8GUXpPCa5JZNtrrqMPlxmN7pS0fPX9T85
+y6AYHPI6fGoIqs8zNTtpRHrbg+zid83Z0vaCs7Fw18POSilR0fipb3vtQUK5tyf
Mnd2rEch+52bgS452pLCkCFKZ2ZT/tm+jckVkhHjRVb4rAXiloOhoHFGqefwDdlM
Fw54YL9Q8B7HZr+6HN3pn/1tJ4gd3Q4MmMU7ELH8aH6JvDCWPo1Pd4Lp7iCe8Nsj
JcfIhlPipRlTUcC5R8QIX/ssPvdqYAAXbC0si/K9WQA1AhDYGBdMdQ4Z+4EzHmEo
vhb/O/zGmxqQVPLkYCojXFcKSSKpDIToOdjTpAYLZwa0zWUNY869SKEeIcQ5WlY0
FzCUIx9I0m4bKu4neKz5nZuyfc6wRGTrwTV/fwGrqX9eWuAGTBPv4wBEVwsOzb2m
3MoBgES9VYVJWbQ08aDWThQMmBCTrEzuXgKGyEMMwPxyZ0E0WNfhulNZk1F8H/ye
kQ5pDpJvXVfcNS5GySBP/IK03c63soR9zQwuYrzU5coVmazTqlq1k4Zp/f35p9UU
Z7aVzRAAjOLVBtlETACw6voDaMYT39yaHaj75ah/RpvpDhelVsCI9/iO91KtQ1Du
o43k2GXAjlkVNvPIx3y4VC48GuMZr4pHIzFTPiurtUIsiDraQZ5YkJI0tZ0f1M6l
vBVytnPJcDKabHMhjb+hH1YYUGFDMuddZjU/ALFE6s/VXZBXd2Os+W+lbFHoe8dP
xKOIUKgk8+FxyRB8S6WOuSH+6SGquMapzs2JIK6B3krDu63QCE0o81+dnYVzXhzr
ytCvg8Ua7j39LGg9osKf/opZgtBE4bcALkXeE52u4wCOQjA1Umad40dL99FJgkW6
jiZTO/s+iG95HyZBv765XBtnsuUSTx70ka305iMpeZUbjDwbizxj1z4vjPyaZZCU
Xcyekzc3mZZ3IjczfTNNBZr1f/i99CH/b9bWZPf0psLHcZUTM4muAf/VfDXe46FM
eqQZXdDO3cz/RkpFbKt36V5ouixtg7CtKblQjAInlma/rIYbitJzyZ/xLSRlVk4t
v+sJNq6q3eqPTHtQ7ZIj7oRm3ga+y/GNGA7NcEgYQ9w8yCJfvPwhJDbhO6P20z7U
AmqEUu+CfkdA+n2K7dslt9NRCqyirszo2RVKcDT+jwjD6sLrShaqBbDn8Ea2x6r8
0mxnP47B+ChO7oAZFLw5gVDvyVukr7P07Nr3cv5sJTEiuoDBnb4vt1rXtubdDgoc
kgz+Rt8ZcGVFFtoFuX6NfxqrscUrU4FS0SH1seDVF76ICgkMms6qBdexu4535CPT
03VztEzPDOlJ93Eumv0UjeNjut7nNpul3j6wEsSgwzzFm7JILjHctgJ0Yq+lJHRo
w/JT6pcQ3t7NahiNCdakZkWgszaNlAB5715G1gMZkNwTKBKszw+Q6l7PuSlVeAlz
OLEsJkoN2twK+m7oQ9p7knfNE3krolhP1pNDlvAveDtQrBDinU54yv9E+8QYzbut
tEEIEMqGkXuFTZRgcx+IItXzPYf+lxNNmegLJCZ9BS/QhHRRZuZACq/2mAySLHK3
87TxFIKOcG8Ib6e6fMlymPkJX8BI5+wAOQr0ZsqcKpCfHJI0N3JgXw1JfmOYfxPb
ma4fT4RgSxLxNmZHlJm3m7WqWJtt0W3OCMfRM79rFf4WJfjUrTREE7dj/rR9QO8e
zPJw2R1Rd+sVo2nroZUGzlD9SwO7qtMmnUI8MrjEW/Tfzwqt7fsHyM4ph0fir/YD
QSoAM17KTxFnRHVK25OtT0a0wI6Jk05zVqAXveRMa+7AnkWcTd8WCteXIR5GpAiX
kebeiCY2GpVUr6Unenqh2bwdXRrTgipV3ZpApCWN+va5kE9OwX6xBgm5UsVyy+5i
p+VzVVsQQ/hCZjeXjE4D4Muo2XFRbev9lFdn8PX8J4uJXg+ZB1TxdBpMISYTRwuJ
trJ0V/heHhXF37t20zil7N4/7SEHi7DujK4MoJzbRjXHr38AJzBD2vF9hYEXEhqp
59tL/vJxuZsH3Hh+RsaSbqZ3KuXKq/UE6VIwbGPFRnLGtqVglcY6CwDicpNolCEn
K23ojMvDIwNxl4jklPnJWP+UWmtdgNDAZxCS7skFOGrdVIFBgREUB0mTBMLmJoQf
KG3QD12PjgKVvtnDmjn6sBXNeQAU1zE+oIIhlM3AEft56hG4IBkBh4RewedgCHFN
WB/5/bhTKvAN3DtmVwrStMfOcvB1MS6gPpX04oCBWVzIoBZQ8GpE0ol2AfEeSXIu
wfZpbPzHFwpbReOqsEHcyJtrepwufap56XCxcvjQfOEDHMhp81T98lq+2IuDDS1r
E7y+vlcKoRNgGVjIGthnP2wj8L3UEcYYwHbO4H/IXC7J2NnjtrmHYyzAxsL8aKgJ
6vMY3+3VTmZX8OxjcqkSx32U81yfMZ38pauFyW/56Ex1hYOILpP8sZF/EvPSGsR1
/8A9+yXSKX3vbUMbYGXTMTz3vG3UWbw3PB33qbvzAYBsO5V/NL8I+Dd4gRo/qM/2
UA/Fk5g2HLvixe/F3B8oL6DeRQLpLikCUV0feJaCLzX+8GApZYJx0ZhDfhPE2G6y
3jkXIX4AQOGy6oWQwlQR7JU3ojtMgyo812jaL5SxAgnKunqtdbxtJ9TzC6Fhq5To
/EF9cX22t22xpHT6u96D+DSu349p5vqwt5R0JTuDoabchgymPOI4gusQciGQABIn
b1hztIu29A/CG9JbwN1kOjBbb5+LHTsOAuAkL9qHBZowXAmcIxa6Upqqb2yXRjPj
QKdCV4y6e+vMrXNDfJkKnX01NvJoJ1Ntmls7zN9fkV161eB5JvbdjhArzFTNYADs
9FGpNkSrxsmh+NwAAL2mSDcFSb8Aiaeql+0G3HPAY+7fIBwDYtYbtjNypFx0UAod
ren8aQiaj0Y38Kw4x6Sbb4Zoe3iD8UyuyfSsAQ91WI4wggN8RFLx/3pNLxO96Ad7
JC3U5+TNY8iM/1RqpSAaKyk33OIgDcVCHfOAXwYHyFECd99xCneuvedWqTT/VjBU
ZdqDAM9wo4fYaCDSvgaVIMDy7jQlKtYNfGOXC2mm7xg3FgobkKtFgrR8hZvXX+Y3
6DADEoxXCZsvRw9olhRF7hVNL0LI/PXjSDcQ6m9hjEkm3rdtYzwGytzB6Q39YXvY
gwk5nrLqMVqOdyhZ7/iLCJE/jBz7lICwstmfN5C19Upwd5riZCIoMLGTQ2IoGmRS
cq3xaIQS5ZNccbxVGWj49QX3WZROZYrHJX3wuwuPsvfoJdIZWmhWxCXs0jW0lcgD
3gln4cJbVXDmWCHQqptldzFiFUEkEIReUYOGIi3y7cel1IJZt6igZglk8XTu6Uod
jbjSgYQsO0GaJAACDcWjYhEwNUIJXzyfHhoWFDAU1G/KZJCma422lJoc2F9fKuzx
P/ih9oJOTXAqIfew1PrT06GF3LFLqcXZJ7Rt/bKFldHMF/pwCIv5rSVMfysQkkn+
P8u3waSk/P1OibSWaU+K12i9/sA+L4yPrM5j9s8Rti4Y5EKgHDEG1O3PWRXCKhn1
cisGBPA9uuTqTwpVkSOtZVTkWCZJYgwTeBhzMJCzbzA86Ro9Yfje2qlXcvEvIRxO
8UOC+p4N05cOPEPaaEvusGLcWnunUfpBe+ZtLB8AcQeG6YyAcwYRVc5cOCPhNuLK
AhiNgX0pEMp6vmZTIc28ETSqMPocvuMIAE0GCFTScLy6URNpuiMNE3C/6k0hGtLd
Yi+Q5qe8JZTNW2snzFHhL5nGX+x/bMK2wfQfG67C6LWy75AKfPNKbw4BxUsVbRrf
7MvS2i8X7x9ZYEMU64U25RNMELGwIoHSB/YzRBgxQbqYZa6EFPCu0JmY0GjJZvCJ
K5LXANwDTQ2pQMzpC6KGu/zFVBPKDPbrICIoDu7+zGBfSaGbhPjHyMTOHj7s6QCM
rxumC2c9A6DD4G/gjtQvCfICQFGqrCtMZDj+qDSBBKzCW5HJA0JNhdN71kvlyjkX
BRjTUnP435/kBvL7vKZrj0Pl+PQGbQnWcsZvrasfPSzZkZiTbUU+qifZy97Yg7q0
Mtah5CcUHw56M3yWfC/eeYRQV4kzJkHnyUhkxlA6BJjLhevArRA3eD7VwlrfBpPy
RpwoZB7/0b+uhLJKLxEkpPdL7NDALrEDA1J4xNehSl5cA/1hByEK4xAxtfIXj6KF
xbJFuCT6DAN9shu4sDASxyHwG433AOiCWDJi1jSvlTREy/WxSKhvjqEQBCo15gdA
ietPOsBJhZQy2dktmtDwJgpw5w677omCghTfbltxWZsn9K87fsoblblfzkYYeAR1
pxAP8L+cfXBv/0b7WATY7lRJH1tnWb8Qc/GsRu5vfOtE6GBQzW+1CI9dtX8ozKBo
StIZwxWm5ToS8/LGFSCyFZOog1AqcQop5Nadhlg+o/A6NGBRQmTlIi+Dmr3sSYSs
KfJGx2phKMg8WGQ8FsInbIOshglRMorF+lpjo8Y3H4PlzmI8A+44EjjKPyRSQg4/
NgNCU9e9fjCZSqH7aPJKhO0zRFHVL6H/VwwqTrp3B3nfnEopohyGO2NXtgBlxx1q
Nv3io5aHgG9vN2PtzUVdufJijuEwaqe8M9CEV8DGrh6b4fBP68VkzUZ8wY03xjiT
wtEBeYUPnEv+GEHba9sBK1hDKm3/ZChzgz2MMLUOF7v7kRPeQg0izAYi6iarnNGn
32FMPlHPeSrf6f54yh2HU4JPmSGuZauijdBwuepKNOxdhZMca0Tfflr4wfNK/8xn
tMM3yzg5GM/NHlnwbPd6y4penRvh46T264ew2pfr8Vs+c+798tWR0PlGEGWOOXzl
vjs24nNOOWLnS7al0w83rjGWjfPGlreTW9MSS5yMZLzwnja4wNKm2VeodMWjru1O
jNrBnxYpT9Bti/BO5K6nPGR9RFaEegtkxvqLeyX26DJzeoS7qOAsMuuig2Vqdgnk
5OSpF3PqMvwGDq+Ap5JpADXtCpmlXDXp0y8/vTsrn5ZjW8dPIMgXQUILcTvYXsMh
2ZurC1XTB7L2c5hKZJu2PikmsrBidMcIibQzxE45U0JcQV5Sr+zUwkUbN1dsNEJr
Iu8hr99R6le+q+Uw0b9uiJBQdX0s1s6kugZHdGJL3sssHCpjVuBbh+/kswntY7uB
bWy2+VwJq17lZ/Vhz4764v9p9ZqzsfgJjGx4EgaZtCsDemtlb05EVdrSbVmIHUGz
IBGMmxF0pvtmVFNic8aAejGdQvWII6L7Tqs6NNNFGYnGl3+3kjJSimz74XGT7d1Z
tn7acTODIpM/2OWzhDjdrdm1NhX2V0hiVUYRJtavfi+jqMRDFhlxq35pWfcSWFRk
5xdZZltKCIYsqjDMXREvWEOfqrcQ14yUPSNTSxJvWTVJm6OhzHgaKM4uZ1ehQ4Z5
Iba4E2ZjpkXuxtN57JvKS/bgGxpjkIAULZQH+wG7RpII5P6Pz2cRXzgVCPD4ZZ/i
19PbT9KVRx9G93MVh3S7ieqA/PzS51zIrqbmDoL3KGzqPqceZbcTkz/CfoxmhN4n
MYjHqd3cb3cBmVbyx3GUG/jNU4kOXQCj/Yo0R0TrggPZyTpgvD/icbnROpZn7K0i
ZdWvDZE4IqS0IHp3YUI+RrKxARpfv7oBauUv9LEkiy4gkJ6el1ubvZALd41CYSi+
gI2VdgP28tg/+EF2xbMU8BXMj7Q0t1uWw866J0k8wSsblIqeoALvKyzdtCegspHF
4SwjCwGDrAj0hU7xyGWb5h0SgSSTVPDDT5HMsj1z3YAUZH3aII7Gv/4jx2tm4gj2
4Pc0yEBkloEpJpA7TSsXghelh0FNc5RQE4Zm2huAZvtr6vgL+mdG8YFa58N3Yr6+
wkepsdgyCMvCpCcjQQ50Xpp05FIJBaiH5yCEdd0SHMMRp8Ab3T49qY2DRx4m3hdb
STTJjTCpD2LANebVbOub0nKXBeqhJeRVxWBnRgCmC6JynJw8+/GHKmZlrtJ3uDRj
/hefZ12OHXebHnZ/9zv77mrx06b6UGs3sORr14nLoGmkPFGGl3njDhqNbBs/r746
ayhuqpK/vLyNGB0hiGfUwIgouFhOyLWHnuv0zPI00rxDiFBMIGFBllsbvrXe60yf
z2Hjwm9dwPZcdmR/TgJB50zEcXm8sJzPECPJxlNybjssMaP6NvIn6NhBHmSFpwjx
gbdVPsTvVVXOgHtXgZH+LX3AzJA6YH9U9m4O21DQWCNozvHIS2N8fuVwt5ZuVmcP
p6EnuaoHkdzxUoFi5y3fd1zosQyuIHRZgDT+g7B51ZLNjhaX/L+DFmhQX4w7OfDb
tLyPZaNs9NaI4po5euA4B0dB046UmIHqCD8KD9W3ejHEbb4Si+fswDe21/FgWGxY
JbqNA4eVlUIFL6uOi3z9U+H0/45AYXs7/7IgEMniuzcUMCN/emdqr3YEgmzpvulF
gBcBHerFVUgOXVmWsy5496K9+e5g2aXnLSkysFcda8o6CHGnPuq9uT/ASzW8g7Ab
H1t3oViSUQk3YXTeK2Jw6uSv0gc0Bpc+WLyh2wBdERPntuWdGV7N/MtfwFwdoE/I
y4C7r37eMY4AAvp6C8FHBAqfMsx2+OSm8soU88gw6PWze3+2jBZ0gF9KBQq5WI37
ZbPUUvuYRsjtv8hnaiG90mKY2U0nHs/ZS/mlP9oZsJ8bsz6vuRRE0yjtuAKDRfy1
XJH8oTc98xDbmYH0VPGQLkLBeL2yRygT78ygYThqZnhTbtDJ5R5+JNotWJlcW+Oa
m5x+SV6OnetpD+ISOQPYv9hEZ9s6v4yppciKYavWOl3iy08D2MiOPD1+V52ecbDa
EcYDlVUfdck2HrpEUw09Vpe57WuSZwcirYCch5n1AD4eZ7O8/SJHCUJBllfh6GyQ
CsDn4uLdrAv0uFXA0it8RJGHIkL6kgKAon6zaiChYKhTNtB41Y2FunbNOSToNmf6
9IopcA3YPaexNwsrPf3mNKh1ibbIZAQzuZVMCxxAJB59N+Ht6LQS8dvKCMZevkHE
kRhO6vlMou86zfM6OY6gx6Vzu1qbX64O7k6e0kd6tncOq/YVnre9bxBZrtDJFJdQ
hDKGfer9eGmi6u45HDd99gjlSFkElimZA7wU9o4JN0jGzibDK3EIzC2+rXCqcwd9
QTxnOVSKQJCRQMfAc/Lu1Cx9dHNA31QkFrCigsphZeF+tk6I03d0i2oxilwzf/5Q
hmULxfFltIFUWwsDeisntc9pWKKvct7PuJq/7UoYbdHXUbm0jU4CCowdNhJnPYGF
3drH+qH59/NhrxY5+h5sNn0OGliWGEIuV4pBlFBFU51UpCf3Ns79a8UAv1JBwWU+
CuyqT7AWKc8VYDKXLAGRAhDZRbut8GuA40bSakMaG7zqSdIOVbZuN9R3mEWr1Fxy
whZer0bYlKLIAR/ykJKqit7Gln0KD9jLITlgLETs4v8uQ5VnTyavwWA6AidgV8Ew
FjUI62qAAltxCnEkSSCFYS2P1F9QG+ULH7W1DnI1UXNUcqO6Y/xbe2i8U4BnW0Sa
aafZl8jbdzvsh3g3xdxmNmRtzFYswv4orPEMWFVjBIWx1yMfk4i78Q0iBdKb8Lq/
RW+jNczW3fnKcT4M2mHqMUQpaR1NnZurCDMSIlgUC6gR+YiORJkomJKUP9fhK4pY
lcjdyVW5ExYb1AnL4WYRgH1VwfoSI9M6eL/WV8rT8anDpUeun+hU08cprsTdmEos
WPFKQgjL/unu8DomXKJHi/6+iYzsvL7ecy2avJ6snwPwGsr0xLikubA5k//eIq2a
Aav3c1yGmTNoSHYug+0GqbabwMRoNbM9Pc8VguYx0vhhCNOzTO0kby+n76w+FOch
fTNsytEIcakM/d1R92JN4CNAeUSXfXOm6SD83zIpUZKj7XMF+9XkECkCl4wHT+jF
hWNHR8+V/yEmwo/1J+nTx2hyEO2VEoqow9z4xMZv/HUrUw0WP0EIK17Rd0bfnthG
QX60+WJj3H19qc8t3zye3vsdVnjiwgp3MWRnFf2cFDQosnlNkm79fNSjZgd0EWLO
h96ZmkKZjYZpu+1xhYX7zLn9PHAcBbSvUShpIjgYMYlI+FhG7Gr345KCKoW0HZ4B
rKsthOdiqyuPVkVzw3wKQa6qdVQUTyrWBma3b1DotTx2KcSzBPpaguvy4foW/KKp
GjsqsCCLX6LW3zKwlfbtHqiS/GG+2AHKD1hsFnhNxEy9zG7DrvW5zPa0G+IeUEpk
JvoUpYXnGC6u51JZ8aMzKlnRB4iSxTE5hr8EAmB5na4q4NF5c2UwEJqCaBkHQotQ
C9BSQjJGsubc7Jc6bhmnLTR2e0TQHLdo4m8c+2fkRjYDLYgdVI+3zZPkDTeAu7Oo
2+WN2gxCTaMu3kPP3AsFCzn/8nGIuL3NtIUsdYObpnUEO+M5XJugUCiirFR30tdd
lJ7pml858IO8TJCCiuxpwb0gMYumw5MFlBCikpqmeVftGLNS8VTyNr7CfGESQwAn
Roa2FflQXkllfF+wvM7LOPHstswVBNxu1Ui5P2T0CqrTjJkrhBGBcNZUB7wAz/hy
As09z5ZPr2PD1S7TedKMqmA0h4nFSyQG1uLpm+xtJuGg+dsguGCXcRH9JTYqplPu
wN6FZeL7jB3xpmH2CLdIn2KDE4hyh4ZTRlgzUIjM/EgNJux9CSHvtGJGYiNNF0NY
fMGrxzHo0x+590bD0sFbQfimA+J+jknM6KFDh7Cc9I0g3hRW63wqAwMbhhh+/5qE
KpsR1XMq2Q5Rke1382IASLcylzWEOj2Ww5KK0BcG1S3ITbS2FReEnFhB+yj0wNOS
V5xaKDuBVtE1Ty3SD56+fozZ/H9deoKMNceTZRLrbhY9mMqM+n/QvERhm+cXo2qy
4VqPZBPpwR3Mr/A/HjK8nVncIrYcsDpeBDQb/RtL3wxbgFw1l81/bfPEkNaduASr
N8xJycrzuWrsMi6Iz9pod0UEFgDsn1v6B0w4eTn1n3VRS8Sx6/hJx2K0EOqMCGet
vVuyNTZNZAF1D5nnbWfEdGjCdLNxPdTfxdG/2E7HYxfwQsq2GqOpm7tZx6NCIDuo
pGhMkQ7qtvdGLNDR8hJmpC4HJtUSiUAvYe3a3u71OH95epbshV6I/yFKy+ejnZfA
k3odZbRysiYiijYjZKm1BiDr3WV5TZdEgVMmIoZ1Bl+4s0qVZHQmxWsOQCb5QGNT
iQ/1tzjWPjo7vQkaqpH4QAB7+MCXKP96ZWdqvaDRk70urE3E5cD88KnKjjSVNpTA
9u9sdD+xLny8Ig7Izb5VdLd7mVO5J3VIZ51LnMrtZa52W0odMj3QZnDFlRa2Ngry
mQ7atXdFMWBNs+J7biU+sFhBJayLMtC9x7e0V4LNRJuOTsJZCZVeb8s/FW6HuiV2
d1aLxebgYXM86Axl7fmTA4npDpOERo6+1d4iF29NjIAFQM+ybZio7Rf2tOnZ4BtO
qjTnDFwqzm1RxWVWFmpg7ZjzXuePpWScN70ualIqQGOfaXBBUzyEH0mjN61sVbV4
L+Q3zcU90J1j2xVsciql/II/scFQT6nyTaq8cayRkp0LXxADe8PmfPDWVo5eoKVf
bcUqCfMDGRw5PppzFD1EGh6RMGLnLX44rJPaKHUFzAcolqs3VzXA/E2t02ixnp95
tgSdXlNasvgD1e+ZOqgUA+JBz0oC85ycMHL/J62CIzfOO5346AwMrV4F7sFtRRdv
pi98gzPQgbeCIvW79azHP86G2RtUU0fpWEXUKc8zrkygYn3U1IQUGDAQgwzUJh29
MVBn3WWuDzPCKeRSKcQN4TTETx0f0RJ9C1qeTqk/eLGzN//sfCF8+yPuXoNtzdu3
WVqWQgAoyrFNW42Ax0ogIAe8t1Bi3C6Uf6B7cEOemuOVQh2a4BZak9cvfx6384H5
/CT9+mNcKwuUDbDguW7oFxUXyCYMAkLceqvg1x1FIl1e15pPIT95BYh65OV3ZWfK
E5GqjT5KwMdFRwce9j0LFTeH+qgn2b5loch2ls2PxLFUASx5UE8ZKQxVewEgCy8+
F8R89LM62CV/KqZhd+7UEsKHC2t0IazChemgLvx8sBZMa5UfQ/m1Bb9A3U/KWrM9
egnWxe2JJ0aRGG6wibpLzZrwn6ozK3g5jgiHxqWnhjHTiRcplBnaPDmkOeF6DA/Z
+b+mr3emVhk8jUa9ZqN/yxPWb/nBIV8RbGvlPA5z7tInT7JNq8qrb7JRCGLyCgfa
IyGbEmcGrbX1utEeDv+cqbqVgtI5YvD8XOKRxd7sUaPindCpiemnFmvOjfd/yfxd
yf/ejT6nfRS5Hi2v7/PAeAW3sJCKqIv3xgegQ7cefocLoomlxMWh5xgdMXLq3umI
ZpxlDk1IohKBm2GdoOB+aB/vxKLYF0cxChCm/JVu+tunDsT9WLaZwRwg+GN+4nS1
WAC+83QG8Xz8nL7rKwgFuY+IKhVFzBXvdCUV4zgV8dWMZjXKAQidWyvpUC48Slyj
xL0Qy0MDBUAxQvjWs3LZ1az34egalPpoLnfAUDDL1b9GDRBxGmOBPSvonFcRZ1VX
CvpyaPhtmTW4DdsIB6th3UdSooOtZGgVwiAx5Z1Nufw31nJ1+z3ZPEz7XqS6dDfz
9pTNGm/kC7ua9ZPPsXVrBBbR+/yLfa9vlnrT0sOnhwyc5fXE/F8oiJko2uvMuRPl
FeKQNR9/4XSgdutnWVpDddTXEO0WSoFwwDaxdVNycmWFmrrBYQ63rm9O9K9pKx8b
ndDyfnt8uXgX0y5Lp0I9GKW7zCE+sHwK3LhlCwCv2DShBVJaEbfQj9LtEzcS92Jo
x7DuMxTUpwyBARAq3qiZ6Ns0DAHVbSPIjPbi5fl6iy6N1ff+x6p2qywt9YAhE5iA
smZJEvBdAqW7n8Ry4yz+DNzOS986M6eo1BpA8pPSSlM+9Y+jRSSsfX4A/gW8GQS5
9GaqUmSkdd7Eg2lVyfgQt27+6d4versy9z8UU0JiFF3mRJ6Sahr6i7LJIVxRM5XL
KFZr2rjC1ySm/PSMwvwdlbKZ0JeedurpY9BSffeaLqNV5yUEIAz2/yIiiJv/Gjax
/SlCShIS8kMPRU0RlTGJRryYhMwJC/mu8LXxe7rWF6BYVyfjrWf+M+n82Ie06AIN
OFSuUmeZsATjxmy9asLzZzCQmQNuti9CY2W+wgBLzTjjiWuIuMGf9/j5W3CtEwnX
EASwIjbd/S1yNvH8MzI+SheOLybKVms0+CUJHy73noJZXgfznk/XbL7piif5hD8y
gFoS2SMq41d3BUSypK1OWdX3XQIvltdvzjtRpnt9axke4F0XHme0CyZsOsObRHvz
dsxcs8/HD5roB6GMm9vdZ5Yw9kcKyCAQ1IG3g/KLWizR1BTL1kB4eFvRgT4fkWbT
8EnWrbY2FInfgqyoRNzc/WTmVpDJ7E+unyS9o5sfTNWzYJGDRyyaLnG4TLmSDhEL
mKAyVlaSeUTdbw8jqGkTOjIjucIvlQZ8C/8rVK1XP78T3G4LZb/l0tRBmDfEPHE2
kEdFvRtjMfG5oMqBVIrQidSJqKBv7ICWSbap5bbaDmh3dE9ie98ZzEo5+h7n6fzv
JjVZ+kstETcQIPI+7q23SPJCPWKysecR4HeLv0ligZ79MzviYyHLuP/n9YiONQkY
6DnwLMHF99KUZjYBZ7LOZiq9VN6yuO0N38hFbjD/4UAbz9j9SxqLuyjp0Ba/J3TJ
yRbhSrl32itUlQzyHJwVWYc0+M5yLjGUF/O2/nejWZNN0yk8DIz9/tr/F0IkXLKy
7LefLhtiuxziE777ENJmWk1wL4SAL2be1pyT/KEEprHwiaPP5OrnQeyfnj8BqFeC
BQJ+2Y8uUt844HXUdt1VvDJhIC+7CsLWPlGZpRFjYvw48hVEpkuzN5A18kVqxDpw
THeLDyj3WxXV5WUCWLrHHh31CPtVXlaDpV1l7jPOJJqasUWQLpMOyBDF5nqT2Xwq
gTgROT+DLOCJg0Pce1ShXRZwhhCeaMsi9VLz5Z4XiTn76tI5hz88sw4nWT6sTwzY
B8T3wVcchor9ysi9G77YK0CrgoZ9H8g4T0xnh5z2NvzIFFMQ23xGqXHyIhzWFNpw
ovFPdk6roGsxvWYypxwAg3i4HgRxWzS9oCH/Q88W5RlH2wvu5XSO3TedwhuRf9AD
9lPYxIepoMtxXpDcv4k3UwcaFgoRAGy0U1aoKysmeuMVM0T0mrrZfLThtI03xpKl
W8g/HEXbJHLYw0HKAfUOrlrG98vrUhbaVQRBUDFrABCU6h0P2hhZjWYRsa1x+ENA
vaGaJlMnz/SEK0H+IYEgR7GAPCgWOoxAWsHg5Vw5ROVLGmGl8cJW0MSJhFEDqeMc
ouyMuqxijtlarbguSRyJbLUP/1RNgV4KxqRZlcQqdTJmV6KYZ/thnwsTtpyj/KDZ
6KLeeQZpBJrXbtLolv7xfx5U1ZP78xXSCb9wi1+bj+RgwI/JLIPzdHzv6oshX2Dx
q3WpiXpFz60eYxEQdgXdkXGWZyGFHs39xwp8X5VHe8QtLa2u58tn++Q5yx/W0buE
8C986Pu/JxKRcede2b9ZOa+qz86+GZP0MDLepqOKnHfUbOJNRZG5/mGLqJwKB8lY
MkZwdkMfMuG4C3sKyrOd3AqxEPFSmg8SaxhifWPTYpNld24OSLXQngfjBftaFkIw
Od89jxpcX9s5D5/Nv7Qk8Gtch/j2t437LYRFfeZ80MvjYaFWCL33x5KBBBJOxaYJ
DInf3L6lbM3/47nRB92Auowb/b2403Oxb5/WWTug1tXHmHNYAlFx+y6xqo+JL/uu
cBJdzCX9Lk42lOHQlWCo928qIl0IRklm+kAvj/iCRFnto+qBZarbVA5eDhlKZBMW
uRO4XvenPXVvfcbCKvyrH3qy4YwzbRtbHj1N5Ma0rf4b+p1CXcZSw0edUGdze0Ng
YL3K2VLDHk0jSioJtdtic9mbUjMHdy6NnccU/Re5nkK1/L//QkXwKW3yLc/J6bUU
4q49iFo8fURkmohxcMCHMNMkiKZz6GnZ7lCq0/svTaw35THR/xuZFPM6FCqMm6Gf
jjhr82H+bp+HEnyFLbSMUOQXHKC35nwE31XuqvxSZwGknvl7tx4dN9KnxebUwso+
dWno3+aifyk9LvLeuqPCXXD9YzY32tiC9GR/V8VWH9nCmdrCaZ/FL/hJcQEaPUn7
F8/r08VL1P867IljrJBw9AG5jRNZZAXrboXomfn6xqwidiBCJ/R3giAtuP8KkE9J
SartHpW40EW+a7L8MSHqybpbk+AOjTsS8nVFWY1NWfyMTdy7KL8u/QggjFTTOiMC
nu/sGyY2239UtZPgb2pDsupKfPOX2dDtGwvHe5Jm32DRTyyLwCd0WwZWkoT/8DJs
Xvt8fweJYbtbfs6FECn3vYOEauL14MrFGFXlUfP0ggmR8JrhZvcBpQjRUZe9Cohj
hZDCz3VY3glUFlrfiRsBY7BuZgmDp4pB9PfVAZgANLvMPX/ezx3qAHQcs358EHju
L1M4I7vB2GJJ6jdwYAqJbxDhRbgGodF7Z+URnbJBEZpGvtYYciN0NvEPWqlTRDAq
rY58h+jlDtAxIMvBKf+zcF8vC9J/Awb9jPndTfi+tbN/o4T0Cit+dvaX+zm/6npg
y/iuvHs01HbYKtdyGXDshpjcMOaiPL0AZ5khoPRgOoBoWqDFeIYQ8L36EYgzJh5o
nQpy+0CJtjPG4KLn2SDgdXm2w8uk5N8bVzhdeYufBxflUyHFSGfh+YD3olxhGW9N
7rTB5ocm8dp3r2X1LxCFpvUdw9oM5ybZk0Pbva4H6SQTBCYRFrACOVzjReJMRoZD
+dPxZgc0s9aQwfyLvxnX/dBw1/9WnDU8vLqyDlNPim+cesee7wLvDMaeZvgvy5tp
WolPOe3RtO+EqCOe53a30MFXO8Mjqxhpge0mTAXh9gbIlrBPsfmYMNNaNnjV/meo
nVHxIHxEO2UZVzib0wRpI3hH5fnJOTXJ1xeMHPtGt3I6zudbTVPxe7+QVhomDgSM
sSKGAlLw9phHbYzSOtach0Nzxze5K1ibV/8a+FAHQa2zjxaz07NomYleW0MjMRUM
i04Nas4XKtYlKOpYqN4P7q35UhSj/FPwMGEaCwpvW7zVHtxru3ZdXPyhPsABJiR0
+7sOGkzwg+xc31miUZLPwFIptZ4c5fA7m2zxGycSLXXHih6GNIuv5skbip5VB9SL
M3YM54aSpZTlDzaQ/OddxBXaxDJ0W8UZyiv5UKUrn1LwrHmWAbMhw4EJJDKGMXiU
M+qkZZT1DEO6jcxdt9LFNEpbLfFTguOXsd6OBI4DHoeyRVWLCffvkjjnhz70cJT0
QJzyeIokWGAgm2ouRZ9XM5vL+/EqYSm0tFie9H9AvM0/LsNjA3JAWQypdqhyOEYy
L3Ur50xhzhrO2ngqXP4F/rF+QMaZ7jR+La393ieZ3vlSyGiidOCUGQ7rxBaMOcZR
w/iTdCnqw5E4S2L4Nx6YqrDKkU5IFgCw/IrjP+RA4poJiC21hghy58XffhSbyjTh
bt+QPUG/ImztLzZLjB0EjOaiXVhcV7DubK0XAOQ2MNcZOqg7qJCjpsqw2r2Vxtnw
rauVImZ6Q5jHeScwzJHoQj1yT4wsQ+eRDGTXMIahV2XDsou+8eJaL6edW0uQ716w
MHjr7DzNe1u9SZtiWB0tP+YSLJRGRe0PFcIf4jX0QfPj366cxumbm18WKZOIi5Jd
mNyyL6wfxWIdeptLR2PeYbDIOQiNGqXfbibl8GyJd0vOCWCSBlOp6HDWjYU87cK7
SmdSXeK6ux6RI4nwxU/m9C2d180yIi5TIxNvQDq2vGamlvFRnmMhWKGwKRXmhOfv
cRvJDYgKPOr8plip81GSvZ23c6c+oIqvREOWyeGj1/qNkLCP6WIaq6zeyN4DnnMQ
JUBk1vqLcKThrsBeYRDvllofwT7wFfSFoXz3qF60LCtajoJ1i0b8tJsxIL8Qs4pj
//RqBKYluGtJsvcJ4Wvk2XW21XRVf/nM/PBPyiOU1IpUbIWtN4mCcqJw5PNY1S0k
k9X3b3OKmwUf4P3382+Tv1r8QChzqnPudQ9J16sGHuYPij5hBy9kvSMUCBdWxdBe
FX2q9K8YAYDVP0WuvHFj986wSb5j9QfJ/0poMQeeKH1j7PMArJlWEWJDEDlrm949
WbjOhf4cgZUIwkwhdy2caMhwfIdyZp7xsHvTFbefV+CcA81iAJ9CJOrO9MaxUslv
jKkKv49bY3+8eQTsBeLMgE+dZH2hQTxWYrNMyxpTwqaavfqwE8Lc35bt+61EWNJg
6FLmxmoNfFz3G8+MBDnNEWYyKOoyv3Igp6iHTPiCSSBnWG351bkSunY8SybmbwDt
b0o8qfOwGWHssk9/J+6eKaW71NrTcIUEd0yh3JMEcA+jubHPp4fde1TMYOErPotg
rx9aK7BYuqcOjq7mdW6BqrM9UucCmMBVBOwXZP5KXf0kAGum3gfxofBuxHhOQ+Mr
rH+ZTVJMf+IAmQAUDtPFRlJxxnO8yLynKc6IsV9nuCreITyhcXXlKDCRTQJGLzsz
mIYnO/oxVovQKyWSQ9VeiGhtOFYztFAdyCSwONYhimdIm33Kb7ufLFjSyqs/t2P3
jGk0PEC7E/AGwyMHXaWtX6E74LlK8VlWJANjP6++eMPI11UxwepPsBewfUQeqUZM
b/k83TnyKwcPZh3QwfCFHrVENEnaYLMyivI0knb+4T/bBJw5ce9X4ogOyjtctoA5
g6djTgh2e8aTqdSx8SVY7FxuuYcogZwNPXOyXn/hmdNWOfWWVeN8/HHaqOnwtCB9
sEVcaDeDBCIPKOi3+PKjCARktCH9bERTTOLBeW09ASAmGlDmwUBZm5EaX2hdStuY
M2Pmxp8tM6HMtN7sP03gCX1SSFd5icfiCk/BTaUfU1bwhsdEzoaGUOcHdISyydVE
FsmK5zuFTEUuLEwAGvJ8AIgwUrEPKUoJ27zGuEh11qUJ2Io1ZuHjI1Iw+sUUuWFw
t74o+i4BWTWz9eXjAfIx16K+5QWJyahp3h25qoPAuDDZCDK1qyz/K2lHKxQnFIyp
8/7DEm66/u4H3l+LqpNHjh+Z6hENGSVoslWg8gGlCFMr/KjEinJGTcSPppax0/B7
ZaS/glSBZn2WIDWEYm0kCGGo8c60Hgh8b78hIQhOcTcPZKxLo2YgndwZV/sAbu1j
jLfe0gV0r0LdNFSVHmNYiExyZBh0AMBNu7RqXKVR8uZGhUFkQLMOatLq11ATyQTS
ap/gzY4m42rJvvYh9EuLzN+JZe+bSIbMp6q9efu/yDFt86WwPPgmVPNGGAhcxhp0
vPBqkmOOh70nMoYsanb4K7g0YFl8J0UqqPfnTWlJCjuGmo1E94EuaFJmVcOvdpFJ
Y3XXQWd1MMKsgWcoII5mR9Zo7M/CFGQ7PLQTscFSEP9QBywBTxU+MYOc/I+O1e5o
Fco8Q26+neL8F3HWCgqo9e9HzjTFLNya+OPem8ejhMjSzOcuxs8waqdzkqrNrHCv
KHT5tEoy/rJNZp7DLdIRHe/oHFkfLFk2Dzo/mfgnvSYRfmn+ERHHm+QeZGsJW5T8
CbWKrwr3W1zkZsKFKs7WnMuiTVQeh6Ten58QchNYoPJMCGpUn5qERO6pQBGVv8tQ
3US6GdsvM0A/nePN/H3emgQWAbdcdVTi5xxM6FBb+wE6EUcaF1otpXO3fXlmE7gT
bktk4AjpDz66DHMx/b4kCrpeZvaQLDClhaV1DKcETD3OvCmFNE8AZnhG4y0ood2W
i7bBOOkGcEii1ly2hruBnQLqDK4pC7RD26gCXJEX/atEy3TSUEQo8EETGRVkRkDP
2fq7ZHkSsRx8VYYJfzSoa43yKHS0RQ3AVOTlIOgSQSUs+J/nWrmBGGmWvGXQ4Jed
bfFyehR03KU2fVIGSS4vSaf+H82LCyKL3A6l4D5BJgthhdYzRx+L/2lmey6DHLak
rJh+vdf7dc9rW5oZ73aqDM8PgWqy2I1jFKu77LDe0iKZIAxbDdwLFWiqYzxyiqzW
QyCN9UziebA4x5iZfGTfxwyHl1+nAXJf82NrR0JJpDZ77RHnItuSWg6+2mOkXwWk
U0JfHlk6qHs6IkI3F2gCzeMYSHsYeAj0THSHqdoc9btxv6Vcde52xw58zS/WT/2O
qgXxYWtncs7kM0M+MqG08fB6h4sXIL1AuuTN0AQaHJLY2NVFUyNDWD5JW55laayE
49HO8nw2zPMcUv6rwMyVLhBQ3LfRMissfNtAUvzl4AVjZx69/8xnX7Yi2h+v+gNO
5/iNPfh3svHOmNYzkt6z1IDtI3DlWkoT5dlltHKeIwIqkT0kl4w2tjqP+X5nlgJB
5vntODmAI5jiQWP23oXwTUSd9I5wM22aXp1ACarDHwLtCsrbIre+BCOWMTUszKCC
7bJrkeYx/gRMihkXaeFA0qUwLXE6uxUqRaff1rkAYRkwZrObGKSF41uJk7GijLo4
qd/mKMwMOF851wm2JQ7tmmCNVnqhsejaHGEP0xqKTRlkVwmIRIqdzEo+7ahhDutg
df/diOlv46bJvh6dG/zeGuiC4X+gfxs3b5WkkkYkXwKisaEVC5MxxC3P2iqI7IKP
j+w/QrGcLO0qYeLMMy+XdvpNxP4UF+2DG+3JL18ysMMTzY1hNGKKT5+Z8eU55nSP
AzfRNhVF7mFd7nLYrhdgaPJk1nT9kBJ2vygaJZUeWyUmVjbq9A1igJ+Xh7+v0BYi
vyZYo5kM2JiLhw1DttNRFB/Tu+xcbCrzvH+ZUqqH2BznM4ErICGXaSavG5UTYWfs
+I0ShJKVzp3Ll1UNZKuVHqYLe/lAiOUoS31Kh+UUJHO9NAROTNXNbisO6NH/kfFb
P61vu8dA2nBg1KsvOqpz9bjXdDmrTISynw6AMed5tHilaYcBviPx8QmfAqdsqfxJ
RH0jIce56ZTk+eUBEXHvoL4s+OIO1xi6ejHjPOp3TaK6p13kRUF3bg2esA9mUrux
4V1tCro3CYbqAlViQtvFSflMkrztxBb34la/0DS7Wl5llktJ13EnQo1KouJ1iSQm
T45EqWF4tHcaqQdK+pQXhtPiGpJYPX3KCadtObL+rjFNW5MevZ0DZ8oozW+xJ8OZ
5/cR1f7MP/U7YXq8e5ZLB22Z383SWnZOItZ1gD3faChPd1plnjaAfR4YW5Y7vUCh
btuUWloHHMfelNozTYccbzDWvfeMCcummfhiNhgl/3+7kk3WdmoGqBs62RRDC+pN
TBQiPdXoWNmh5xT3kQg9Zjj7++A+l2F/uSpTzKiQku4dgP196AOkvOOcoZOHmki0
WulyM/rJ6FoZdQ6VpGRVV//afb0rUAipSYdUSelirW58n+GzjQwGExn8Fm/e1uCq
A0W+uyJv9o/7yGevtxMoWEgGpivi8luMb+1xdal8mlsYhYUgGnq7U3dHujANys2p
hVLXmReRRiKC45Rw9iypxzD3jcfA7eiFZEXunfvastnTFMN8KvGEQNCo8l4TY9eI
/Dx3K4PRNa6yRKjH99jDKmYrmlbkG3Y6KbtmC/oK2Dyl/o5btdv197YgdRU1Fuw9
W5ngF0Cgd/4wIMCqdaWD2MHhhd8omD85LBfD32zzGxr4EpejsHR373k2qjjG0ANJ
Rsu2LPvTTD+/jhgexMnLAtMZACZYr5D4jUpwgMUMSOyxQA3pISmZalUuvn4v2tnd
xM6PIAN1i1LSlGN4tXwkj3VHeOv81hW7Kpx1VowVYk0XxwQiKnQfg7EvzMC5G1rL
91M9WQBZw32HFLIm8xo7WOBQndU7jHg6lLhbTv7a2bwHKvTvr/1ZwzAZ2/UKM0VI
L8ryR5+Ej6pBuF+dHT89jqruV4wkqmuce5RdfSR4VV262Uu1qV7RpV2u97BM/SJC
k7K0RrWw321Z3LH2aomMkE0zCzkeLfSPr1CArFER74jFWvALIv0oNwX/jyZH3JLa
1kcixvVqSY2FsrtuxCmjzajAe5N/FK/fn5ckWE+s0fMJqoTBI+W3GiXY755MyrFp
pyo/J11yyAMgBj4m3JOWNWl3ajFZzMhWB95ApkS/PuEMu+XnHs1giI7wtgDGbX12
jmViZRaDbe9eUb0uuGEb/iOVuHysIQZlIucf/e0scTBMDhSK6ARe8E1NH5YXdGpe
lFYctHBZO3uGF6WPkzw98f6CUzRgUxclGg3hiv7g01/XfJY9ZqDlI6QDAXlRZ7lg
ByodovujvTuxqmpV9CdPeNG4xpwQP3u6hHv0WglxJ/wUf/0dlPWmlrIeQc+/o+im
DZ23v7eDA2Zn/DDRrVQYW1STkqXna5luJB5I6hwlP02fZfq74fAewxpDgcawrJLh
dJ2l748UU2wTqKinXJsh98BspM9jhy6CYugvufxyNOw32yqzKLBsyRVWzYWJwxgX
ZnJ6MPpgATFSqnC1Hi/+VeqrthhxQJdOG+HbJK7XQGuwPHXOJERxhOQ6nN+3WnAF
Hi/fnx2vw/phq7xwuZxKIOlK+jraLewO7SplszZS3WcC/OUTke15S40oxII+HsM3
clrDzWPkwOsydfCr045XAt1uKF44cZbiHPDP3eVf/TBMvQ74uUajLNqywXpYuZSi
uFLlSsPEoON8+1SQSsW/4VbpB66mRESf1yJN3xbbqPnou/u1xXe8rISAUim7BqVV
4jqiS7JYICrEE+E/DCOH+Y0ZeU8YR+osEVPjidhn5qYEkJBKvkgClmTafUN+Xb8B
NU4bVDbd6K7llkA/uCfRjc9Y03f7wryff35d5g6NHyrrrPdvgFbzgTY1bKJSn94h
ug5vFYjhqL4TITnAk65E6VsKfRue5/OIF107oyeewLtjiheUsVERwPZOfrB9LR0B
9uvJp3qNJ+dU3n5swKGApch86ry48U5t9YLVbMPqCuuTIahvBvH46i9E0G58xoNT
ZSN6dxjaSd97IgN1QFFhHncYeIms6RGYYQEtNZTK3jWh0Iw4BfDC422VBTiMAIMI
o8F6AFRLKKDD0p4aQ+y5dhBrABUr/c+4/hjhJnN5KLAELwZQaYXANhcqqdasbPB5
HRIeC8A3hY9SixIzcG/j1FAEZhRikApHmMDIon0zYJxxRAZHCF+Bjf1TUqnBAor7
tTeB1tN05lmRF8Q1JbHy1QcavCXLaODQHVkWgPIsWUmQlaLGP1y6OTspUTCjCDFm
qAAfVdNXG4I8jcdQZ2eonWKFMdxVcbcQG3cGa7XZVOQUZefgqmd5Z2OZSEb6v9jw
skgSsClBDre8+I3uB4X8FsYHC+5ME01EI2XaLDuVjf7ePPRuuGf04exPNu7YZEvX
OFdZgVy9umGQM/2qRE9sFfqGnGBtS3wMSLuEohjresz1nN8FtPD54evlCHWwl1EQ
tLxBOMmBVRMf8EMueI9FMwuoV3eJQZMSxKNayHPAcztAcWIEN0+BsEC7om+qU+A5
dfu9djJBgjhVkHo697YQDb9hstFjwztTGaAIAwesE/rSUtoMgjS9B5IiRysjA2nl
+y98F7R7pvuQLQ7PtNpwVcwu0IYcCbNevGF8dXhhmsfY3wk16wXAm6n4+XVOLvVi
KuR4O8xKs7emMM3Lpl4nRhi9vw7T85/fkvTcihOQIJEgN+Tct1or0Pl06RBQocN/
rQ3r0unuiI71CloIoUOrXiXFn69TDXZOhkkIUKfcuREtsB/Cq3x5e8ouaJN/ANbx
q09sMAHB93c4m2N1r7z4zO/NOx6qDJml1wzUdk0W5c/uBPrsy3L1ekvjsJoWWAKi
cj+jZ3aTUuiuNDEhtqNeUEPR72DPHU/JNGZrvg9+J+OM0ROvV4XKDyj5tfL/3y/q
0bShGmLKw5XYYQIv/SEch3Fr2EM8P2m2nnQvdh8pSAmCxSR81vddbiJuIIymIUTO
cuUmmSQSDv8xIIWmcV/hbRDwngLu/u/gMAHDhcWUn/fTLbhrZh7sYTUtd6mxr6s8
HYKSi3miT/g5fRon4MP7R/LXWxjjCuJAwOMv2m1GJ26OuB/kAopa5OoyehY2uvuR
y3CoQsT3XbBP55Tm1lkU81blOWxRl62S708EBK17iJUNq04mBuzbEl8ttfgSEwQl
d6mtfqigBFyFM+nilTchhJyqAdL2om+yHmGDXVpA1hNVME0PA+5cJ0zEfqiJYYw7
s98dOBtTj169W4FTmBONLoZ+0KKeVj9iAWNpJ+TXnikQJerQ4mq2RXd+zTPc34pM
5qplnG3RBlljgqunZNV3peq4fPP4sAPJ+s1F74EJhVL83896g1a4A9eK/uq7JwmH
JY/hPBStu3MMTf/O5l0mbwX+iVvKLvDt8tTLhm2E/TTzqYo5WdNQh6/UWYQyKTVG
SZXLv7WGFSfQhpqwzNy62axcWsKiuB8sp/UjqQZcCvXIV6ZLZha4Uv7ieDHMK75p
dSUDLnqx7a8fOlBJYRuXQnEjCDq6yrdmImKh74OWF+ndblLa3oA/B4yXj/7nS0N+
rC3S+wKXNYU6CiJ6gQCdDuNi6PJNVZvlwnkqG+lbmhx+DbbsojqWWClS24tg/GZf
4fuxEzRdD8uHGSeMyTvaFgHWK/UACKeAE1a2PQWs+oAX8GtVd7+16b1TiRC45JhY
rLwHpFbPmhhKOv6V34d4iLZw9e9/cc7lBbWwnobkQWpToTGFVTaOP9A3XyUO+0VA
OuIFiS6t04nPNaC8V54RKiDU8enEkHyVaGHXtkrRAXPBBQjR34n5d+Zl4bLVE0sZ
ZUU4mTsK2IMZ9lMTj4zOHA4FmmfBdUUFl5p/40VsynFEAvoVZsLjKdoe0JDNZeZN
XlLLcnvka7x1opkL0Z9YsTadhdP6eNAsvcaOCvyuz5DhJek1YiNSjMy+2L3pwU5/
L8wYDWExqFTA3nuzSaSG5W41PCOLkEwNP6HZeiOk8tmH0VL5yItZQX9WWWuPgNzo
sdD5CIZXkuGGYvAkKxuV0OIOnKiVh1jTLP/LJYpv42a+tQr/y3gR1Fou+kjCVYpW
jOqd/SfTf/SVpOQSPSYFUsxUpXikGlKBEv0C1Qq1V5lIdvws9IuZym927bBgxpU2
vrxLuTeHZyLJUPb58jz9XFUkwkw76lWbggKM2NIE5vTAUG33igGRlMW5GkPrZqiP
e4RQC73+s6omMq8UyQwcS5UnWX8V7Hq7diwGLgQwAPLhQ9WtgTAEPQlpNI00xr2A
abG/RPXhw0K6xlwsQr7/AJin/uURJFDssMmuadPpy+zVHE1Ii2Zz6iYDdfLqUwas
QkufQmQzjQ82itlNaFrcFVH7NjEM0IcXIPNG2Dk7esRESvnu7fEgJQlDtFrJz4el
uckoqhnlA7Fu5EN1UWp/GF1sT/PscpCskEpH2D2VlyOZ2p4H5ER0elD0ajMaibp4
uJdfK5XZ9GtXIsPXgIyQm7x9vA3WKwVrtcfUyr7qCZ7rdLyM6xDKn9olouSmbOaJ
tZm4+8BBaWviiZevrqq4HXHb8R3QDxSgVW7GV222u67otflsra7GeraeboK27TyL
JlwYFhDQpFND8S7SGvCTfdPHf0DCNmubmxcsPifGn/02Py7zBpagg009FW55WWbw
zeG0v5JowQ1VqVgJz/6oweJxwvB6rKHApXkNw96BaJP2hZ2NTtZPy/LWtwBJuBdR
3ecDfBv3b5OnbOOQhlAs63Q39PaCeajBCC5SUNxFd5qOoKyWxycVu0Mg4GBwilrN
FwkrzZody+NTJiEtiDSIhRm1Sa7eZARXsH7CKFk3rqkhoCt++iWz7xgIO35jXkOx
Y1V+PkFqhobSthOm6frMz45Xn6G/GK67ieCFBfJcXQ0WeuR4c83184CesrTw1TlV
X3oOh5wapx1LBVPfjhZHrySUl1wVvlMD681uODet5Wup4dWR89mAXiJhzM1nsRp/
`pragma protect end_protected
