��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[v܎��⾍{m�@ީ�I�F�b�cb�J��`_K���Z��:�>�_n�t�W���cj�z��Z�`�3!�\l�x�|7�����˂!��� �!Th�)+����K�T+>��~D�j��(�C�L��@�|"�L��"�:�|�����.�A�`$c����"��p����',�MN(�f�"�o���|����N�U�X��iMY�ކ�-֋���uq��M����ʬ�,m|���+ȵ��j����?�}PmwJ9��������U��p'���V�!L/0�Jܤ���#3YՑ�DčY�;��X��KR@�жkBA��C�~SŞrS�Rh;�Z����fl��O���BRHi����a#V��7'��E�j�q�V��	��(��~Uuƶf��^ʹօ��*��Q��Y)��k]Kf6b�{�j|����v%C����2��)�M��*���o;	���N�%���y�Z4�SΐL�B�Ib5秮ZU-�����Q��?f�ea0ɑ7���<#<����Uڮ]�p|0_p��]���t64K���ƴ�ϓ1� 9�����oa��hP?jK��@��;�٨u=7v�G��V��.���i��\Oh^ʉb?�^��
�!j��0�nĐW�/q�e��N�48*;�}��+�Z��е��N��n@'6P���>�A�m�:0��f	�&!�T}�T�A�º�Q��*�k�3q��_:�f̪*��o��Y~�gH`1���[@bP>t��ڞ���H�>rc�97%k���vVx\���Qy�R\�t]F�	���t\&@$�����Q�Q��M3���r���L'Fޟr�=W.o�bK.����`����4[��,2>�J�� IE��R�i`�1܍&%SG�젉�w^q5�����&�D)�1�CQ������d;�(]�)S[/���F��3�pY7�x��� ��v�����l|���4^0��]����ό.��Q���lX�I���IQKr1��:Ajvz�ӆ����2զ�����5�]U�_�&b/VAu@Q{_
S�'E�^�O��K4EHL�I�dNzQL&T���w�����w�:��_מi>� �K����[�<�w�Z�/ì�~�ް��Q�i��G)�i��:�QT��ч΁�9Ŗ~�ϕp�!��ʘ��*E���.���g���'v�5�um8���M�����߷*�{͌}���c54,�5)�6X�)a|���P��b��# q���o�\�Ld�|�h;�����A%ϩ_Y��+n�b$����a��J��8��(,J%��#a�k-��b��n�#EΈ8y��,e+èQ�6��~�g	ma%a�V&�W�3�� � �D��b����o�.!U��׊�y�xј�kiVy�=��->Kt�´�;b��9?�5
K�E���݄�FrRP���G�(��S/��q%�����C>TD��A�&��!s���!��(�b�$�ݻ���0�r\��y*2��R(�%�$P�Ó+��A��C,�V�O��6G#|6�ܢ�uΡYI&ݸRt^*5��u�.��D�� e�p�{�������`�Ӿ��$�O�;=���񜵷����)^f�(o�aIt]���3j�+n]��8�E|vK ��.�u��E�\K�.W�Ҫ��>��`�{��6��
�i�����,�b,̀�֪y�Z��Ԋ5g�fb��;�]��V��=L��/-8y=�.��Jq�O�s�X�y�)��!���=ܶ. �����!Q�Tb�r]�6��QH��_����{]�u."9�);,Y��%�I �$�ɡ�Ar��!��O���Z=���5��C)�2h�jީN�d�p�yNL��_����s`Lo��>���|L�P���s�E�e/S�%Y���X���=V���E o+Rţ�{@�*؂*��u@��n,�"]��BVI@�^�o䶤2FR������Rl)��;1#�?�M�S������uK� ��'纬��nEq:���4�����,N>��p���Xt��UlV�؟�K�ms�곭5�մ3�cgd���ϢWrG��>S��;���R����~��q4apl���<Q����z�h��!�#L�o�z�6�<��v����������;���K	��㫹TX5\eW���QsƋ�N�;��Cw��Z]�R��O���\�V����X d�5��ܠ{T��ذ���ѫVQ�6%A�H��1�����/w��GlO6�h�O����n�G��r�x^��)t_��ߧB�[RG��gw�*[i�g�M�oc�
U�ἢ��p��%l�+���h���e���d7���=�=jU�R����»7 H%sY=s׹%��[j_:�A�*����@�h����v43T|��nb.ue"a5�2_$�GӦ�U���V�"�S��]c�;������0O�L�}�\h�TN��!�&𪗪�m��O��ۊ��dm��%G�QJ�׬A0���0A���h�p-"���g`�����N�6o��Q����U�t�{lf�s�HӼN��fPj籉�=Lۘ���,�����y��pnNB[�0P�.����<be��I?�a����d��nZ�,o  J��#n�O!K�T�_I���JX�%WV���x�?F��I#�K���,���:�㗃?Y,����d�V#�%��weUr=�h��#�'�k��aD�q"c��c�*c�6C��$�:;fx/dJp0��&Vt13��B� {���G/#�xI�u�[)�?q�;�{,�����_�R�
��7�Q���������}PO$���Sy:k3j�}��4H:�9�8������F�+�).�a���1���s��W(���2�����<������8��^3��a����=_��6"���L�\��݌_*�5j���҃���ɘ\�e
8����Y�R5��Z>,;���Vq�d˩"�	r������OB��Z���;� j}�_L�\�y�#۬��`O�c^�ƿ����7�%J�� }��	❚�mAؿ��a�=�;��V[o�"U��X[Vj 	l��"p;�8��d�
n��vc���ň����� �\�h����k��y�<y�a�����sMb� 7��\�^�΋��{�t�N�k���2�Ռ��RU='��-L��}\J�D���KL��͓^{/w�ԃ$��S���t��F�1��<�e�A��D��_���D���O�����Omw��&6����e�I��y�2�s��d��^�`�Aĳ����9�����>���f�;��L �!K#)�sc@NDA�,st|Pkc�$�Zy���ar�^��h��I8C����F��j��t�)�.<ߚ��pf#�O�Y��0���V�d�߾X\��MuXc��[�v�wC������OA�p9\���i�-�Ch�˼����:��b������gǐ7���B��-N�!�ɫ�]�����Uه��� Ԣ��=�=�s�_�O:Έ�[b�:�����es=%�W�`3��)�W♵|N�pL�U++�Y5��"X��#�E��91P��@JOm��b�{���'-�z��^Ю����-F�`�̤)�$}�X��X���y@���W�����D�	9L=K{;�tx��f�	�y���'��$ױф?�k�w���m=+�pQE=��u�%���7���qbMn��
- �d�U��k�7=)��W����zu���t1�KCW����P�K�<���3D�,⭢�[��챳�J7���d�d\*H�RF릶>���mӚ�0�8�U?�wM�Vg��^�[8�\b���"U٥{�N#[��78��T�����M=*������Q�b1"j�X3���ϛ�⁳8��
�t���1xjHz&6��P��هќ�-�6�)��+E��&�~���f��4��m�����l%*;�5�&�Q|�Į��g�̊�����t����-$ֳq�E$�{�o�}-�&��A��Y#��'�T��2HM�kW��]"�/���
��5�ݰ����!1-��Dq���[L���Ek	]�V�S�-D�Fc#��f"�Q�����6Q�/0��/9��-��bB�T����R�5�����y�<d����36��^``f3Y�9�B�a_/���3�C�L�+��y�"�&1nNA������"SV��6hO5��U
h�V'-'�&k���ُ��u�gg�M�|��ں���W���}�A$	������==9�0�n%~��er�[g`�ۨy�}"w�G����VE��v�KgQ�)N�Ǫ���Z��~q_����$в{SGp8�@�j��{&T�L$W�?˹�����n��zKH�hi�f�C�0D�9�c�B�/8�;��b���1ڶt�m�[>>�5.<�u�X�����P���"�Ox���R�{�=H���a.�"����x�V�v�[��;�P<�a,��Ph��}��| _�׺��c�!�oR��x?�2]�.p��|���'�@�<1�l)8c���|�콻�,˹{�%P"X�|/�}�������\����tbC}���0Y�n%%)�pB�,��n�iz�X�ԝ��F�����S�u�9���O���p�޵����{a�b�:.��c-9��po�x�ɕ������;M��#9�h��GQ��ʄTڽB]��DWoK*B���(
>�?&"Wr$ x�\�]�t'i�s���� t�Z�v����?�`No	O�8�_�Ke���(b�F`�C���1G�橓�X����>H���gO�/�a*�x���g�,;�������m�H�f�9QF�G�=�����-��N�5).�B��<]ًI��"���S�����S���t5m��u?M�Be���<���)W�N��]��_�+���Xlޗ:[J��ǍGo�3u�w1d�tZ�� lp�1>�}"z<a�Ț O�b��9iO<�v�gj��_/xU����I+��ҼN���h
�e�&!P �1����<`g�ugf�E�N�\K)�F����\�[�vN�5L�Fს,�M$<@���)�#��5&bV�X-����,�Q"�B[gqj�~�^�7�~�i5����Lo%�i�@������dL5��jxG`�̓ia ��hdx��$�y{�T�j����x�)t$ѭ����)��#/T����L����m.�2\�ɞ���D%ݗԠR�C4�E����u�=��4���ҳY)�vki��|r�k	��|\8x1�k9���ӎT� �Jge�� ��P�N���#���l���m�R	�v���Z��k�%�nk� ���e���7���ZҏZE��>��݀���Pv��U۞�_C��p|\�:��� ��Â��K��>���)�>�S��>�e��'5�����ۊzt�?���t�^�dE��	l�@��5���[:���4��Q��3Y4!3�n-3��ݫ;��i�s��m��T�rC}
Ǉ4XlS��f���@��k�Q�0��<<�����y#W�M]�� ��/]dfe�~�)�n-�Mô2p:έ�~_�I�B��Ttp�d ��R�N�(����Ͽ�t��r@ወs�z��,�',	�!�B�F�n!���PV	��Uq�ٖ�R�o��="���[V���h�J
OH�]��y��m�B�O��l?�Q���q5����$Z�bz�
pn��;�u���w�'O�s�2��>�9�L�y�H��O�٠�I���^A�R;��YX޼�!�,�J��BK�pC��Nn�3���͆�D�H��:z�aN��ym{vW�P#�r�-���1;E:C١��1��e�2n��*B&A	���i��CDed�������~��i��d�>%�#g�����Ԣp��E�p2l������QG)��X��s�<}ZL��wd|l��Z	��Ψ
���D��@���7��Sp���9��Э��.[+J�2���!��h)s�$��C!x)J�X��x��x_3����w��5�M�(��g(M���u�G*,�����(|�8a=HΌo����F����w���	�v"�K�$`cXĻ?X�S�i�G	q)*,�j�Wj�����W��fY��)\4!)��Y_/c=<�����d����J`Q�ٙ���i��7��$���:�Q¨�2r���Vډ^��-`ꝱ"D �U�h	����!?dm��[\9>�>*��+��Aut����ܴ1�j���\XE/ ����dV{��r�06�s��U���tk�$')��u�a�`{O�0���ч�-_��(��u�������8 �V��x���l/�V���$[X/�BJ�z��1`��U&�v�
����7��:˦�RQ Yy>� �:␊|�,�o���:���f�dNШ�s�,V�����E�;��@Spo&�Ir߭GǏ���#�[y�\��U�T
��-�=�]+|���|1m�*�Am�_{�gb�FRu���o>�Y��%���j�ZK+�o���-�Uݭ��c�����kbqҹ|�C���6�%�,-�� ڪ<=~��
5n�v*�V���l���ʙ6D%��;a���|�v�Mbdw3/�{hD<>�L�u�N]�M��]�]�Ղ֠���Z��Ո}b-�[Gy����&�gLKJd�rr�W���#K0���V�� G=ߓa���R���L�p����&�ʹ�|Ģ�AZ��vuZ���6���]�)��.���Z�Ÿ�9KD
�.���i$N����*���%!f���v�X�aĻ̳�Y�!��P��}�i�<�a	����D�^ٙD-X>�<N�*��$@�V�NiK�źLC$�0i���~l�[SMY��r���a��|�o�9(g#�kvDԵ��
�,K���ݪw&H+��@�i�m��6\��b}V�x[���Uv���8 �t�:{����UWˈ�*�5� $L-��7Ϋ��n�
����M�t�! �C��W2�������%՝Gk�ǩ1g�e	�������}�9/�� ƅH�]M�2sC��n�+Z�&i.�����N��AD|�=����{��G��J}�"MPSӯ�ƽYk	�i��O ��t���R?R����t�<%.Ml����Z`:�u�4+[?
ߑ�v��"t��2�[Ꞿ��.�ŝ����?Ǡ7���+�Ѿ�����w��?�i�so?�~��3"l78��'7[�I�fݭ^��k�b((-��h�2T*�<}���V���`��{�N)B�a�}!J�7t��9��"P�螮 �δ' r�Zf��^(�̈�����I��'�KM�����@�"GD��T 3 ���1�'�iW"S����Z>�f�r�)�)%8:0���w���) ��	��d��H�h�-�ͪ�� �d��_�ګw���2\�\-=
��:�1�3�]JmL����C+�����F��o�C�{\�pK���/`�W�!�tٚAu�ٙ���;��3eu|j��������$pܐebv��� ��^�/�?ш4P�� �Nj{FX�5��ݢ�,��S^�n$���11����D��y}�������V���!���6/��>����Q
�-�o���t�D��K'2{�0�\]7x��J��aKv�Rd�^şWw�5���$��[C�;2%wJ�QlX�W]�])�+K��x�eWM���1'�v��}��T��_-��IB��X��'���Y�(�P�`D6&�r-�9�pm����-��)�c1x��SP�S�}Z�݈bh3�ڑ'�&�~Fh��ǫIS�v\��� 1��{�'��m��|/!�)`i�DA�7�ऍ�~�T��/vϐ���wz�D�i?�D�p�>/1���/�Nm�:���RgZ�>�c9W������tbص���7j
~ΛnJJ�7Ώ��eeh0�����[˗v URT��c9%?�qu�X��ћ"蒵c�����ta����Kn��pZ]!�8��cA(&j��D��2���z��4ز����1��ŧ@��>x� �����^7��^��ml�e��M��5���Ԛ/t�y[� �L7|�'��js&���gl;�zs�� ´� 
�>��>{�߂ �ƛ��ě�_�_R�������X��&.��$0y-�����NZĝ5���03^��S ,�.���~8/�c�x�~+x�Oh�ag8�,f3�t:5q���˛�̤�G��i���ŷ�����P�z��
�AL��6T����]��7�P&�eҡ��}ʱ�z��|f���)�>�(�ʅP����C�u��{�z���)E�)o��fN���>%�!d�0��p�!���>��uQ2����D��Ǣ^�R�J��l�I7o�)q�~g�����^�oRl6�Yf�-zy��	N���T�>��(�h�u�7 #,�*=0�4	�.�#�g���6"|kb��;��D,�U�Hʾ"e�.���I8�e�'�-|����~(DyY�q9�e���sm�1{q�^����h��Y~&L�@7?M�v�˒���}�N�j�jR����)��"&�0������ <g�=��l:q�c�-)�:PF_�"ڽp�+����C�5p�Bأ�h���C���"�Nǹ!��V�]�CH������\�D���5iuꬕ|���;��
0��X	o[��ѕfg̪H��h����R�
����`��v	uH���<v����S,� \��>�n���\������p<i*:��x����M�'a,EHh���?!l�v�L�av+��+�,�
�!_0 ��`)X� #v���j�gh,BG;7|U��N˙���o�A{	��&����jA��A(6�a��7�����*;;{��T^3���PX��t|u�P��c)��H�u��:72��'ĸa�1�Y�Zx*������.B!.JRH�V�؛O�BkK�m�g(X�,��#�l
��\�?>�@�&�I��p�8j`Lb=?x�b��iw�3LH�"bg���O��l���������G�:�~���BJ��oU�B�KW"�_����unnr(�a��`�˫;_�wK��	�����ؙs��#���?�����D���M>Y	?/%}j)^�pr�?�4� a��U�A��-��xM��/"�XEq��l���+c��b6Z���@�UIP\�ݥ�h�xu�y�M�$��
�����UfaE���۬�h쐑�tΧ����-�J���I��|�
�*3'{ .ä*�]\�|ڍ�M��.�:�ֽ;�e����l���d����d�pI ���}Ù�r������)�8�y���0�tOH�Y���#1�:�GU�v�������k���ba�a-6 B����.@s2E�"`��E��/�N��Hm����";�|X\���5 |�����cQk��\�<���1!�O!��*�p<	���~��鉬�9X~\O�!��8����D���AP>TW�:��1!�V�T=�=>�)(HJ��P����.,*) ,�J��UL��mf��U�0x�CZh�?��H��_X��6�]�y�/�T�D�t�)�
g�*/��d�d��TX�fZ��d@�<IE��<G��ʴ�}��Ll��7�ۼjA�>r@Ƴ��[�*3�^. =_�b2�>ɽ0ܡ(^.X����bn��J��Ю�!�2��«�G�2���a������Ӊ��*�(��_��^%j��#�F���Q�wfW��w?��e��ph}}|��nd�/,]�IXλ[��u��P��a��u���>XXŤ{� �W~>��l�����ԝ�}�9�!�ə�N���w�4�9�1�@�Z��x^�5�4:0si! �~��x]�+Dh��u�H}�[�eU�Q4�r�Oڤq��u���z���߈��y�en�ƭ�Ό/{P8|�b�_8�+�d 3��AZp��枇\! :��2�/4���?܍��&"p�	?����H)O.��e��I�ݽVO\]�r`�嘅�直�h����ka��R4?Q.�]�����M5N��ᙂ�Fzd)�8.�9U��d�W����o)o���gE�٦s�X> �ݫ�"]G0�C�6��'G �ʈ��G�z�OhZY�U��)ٗm�Ft��e(�nN/��.O�{��ҙ|Wr�G�Iڎ]A2,@@|� K �mh�Gʇ�6MJ9��m����_H%�I����t�Ћ$�ZS�һ(u�:/|��jyݮ)�	����O���ZD<�M�S|�iI���7~��EtY�,�%7>�[tvZL=0���ء��5^^5�|���!��?���q���4�@UY����N�$L��ȫ�K՛ѯ=��:�Hqm h����9��V���^�8A��gI�ͮ"	�ֱ�n��iZ6�����Δ�S�!�>[�P�������ǽbPj���xR/�������[�aj��PGe~A):��/�;�D��$�S��Tw���S�Bk7���l�{-cM���_Z�h�VX���t,��i�|��uc���܌{��@#�w�'P�_}���B��3�{1�f#2���$��(G�bv�/B��ƾX�8�Y8%�8ɋ���#	�xu�q�l��6��W�ʏ<
s���`.v��k�]�|տ��*S��لa�]�3	�t�Ά���Ek�����d�l3q{�;a��=.J��	s��"
ϓ�#��𻉶k�LK�I_w���Ï��;�K6�2�ma�Ko`Ļα�r�X�3���hh����QgK��澙�,��XW���͔h��Kl�<�[�[&���R/��G�K
Q��L��0'��ީ�R�R���IG��	��[Ŗ%���_lR�ʸ8E���g���Ls�'�d[����	Q_9�ED�(�n^ �-]{h��7�i$�ޙ@���T��HE��ũ��7z�a�b�a�}&X�e�f�,�P�-i�O"�U��7Ø�݌�A]�D�l�3����EKWMC�h�J�8ٽ>^�}��͌p�h�(G
�~�jg�Iz�.�o��R����wG�����0����u����d|N��ٙϊ�:�G���J��y\���zM�������h����k6��T҂-������	P2a�����gB@p�+���Ő���bJr���#=�e�맇���Da�ń��7Q.��0�����Q-�r�MM�=����q�*�Vu��]��y5��n�7�ߎ��7 �o=I.����h��@��Ͱ~d�~�#��5D�
a�_Y~_L��&��(T�.����Ek�C��GĽ%64�Т-�>�w"�a��>2�=ƿ�n���E]��m�`g�0Ǭ"}�k���0��\]D�6?ܯe���*���"��������;�`��n�{��CE͵�E-�Q��b��CW��NJ�O�� e�++� 񕃸6B���0+��'�^�z�*���P)�S��[l�_M�z:9l� ���֙Z�'�k��s;ƒYD닉o����:��;"��~���~��3Q�zc(�^MU��O�,�9;����:��)sI��Ǵ�[l�"�Y?:���­�I�gaL4E�87�7`�6V����NC^�>KSL䦼p��^��wwcE�{��=�U"YH��5��5��J[*���b���`E&�A@��)� 0�%��#.��ի(��Huu�B_?�1Q(�v#:�H#8�&B��&�.>�8{��E�*�BU}�}�C�j�y/'�.	Ra;C��M�7�翞c|�����=@�`XH�a���2�jM�-	��<�.���&k9�*h�p0g+�`�2Hìu�h}z��u����>��g�,�b�g2�Ӝ���>��)��u���E��L/�Wt�|�8d���K%Y��@�ո@Ƴu��Z�7�!5"GL���K�$@AcR�3�ƻf�J�:_L�Sl��l�R5�Z3�	�LQ�7�Th[A�B��Ӂ�d�13ɗQ�e���C=a�:���l���ȨI��� d��jdza�ї�Nń1�n�1��E��$�\1c�UX	�,cXo�QLw��m���T1�G���*z�@�v ��MC�����y8c����Ej2�-��~F��MG�{p���P�㼷6f�2fکpw)G2r'T����h�f��"|-���f,{���-l��~4:�33
+ϳV��ʙNe���<h�-�E�%�<F���?��6R vqb�� ���ZW>k�����)@J��/�=%ؾ�������y'�fԣ|Qv��C5p�{Hj��$ͪ7��q�l�6�a,l"1-��Ѿ�'�iT�t��H8s�R?B�D<�L���\�?��2�fQ�����`�(5�����^Y���s�{�!�'$��PG�g#)�r���Y��(69VR^�?���`�+_k>7����Cs��e��oRUxQ}�L&wiH�7tt�V;�?����yŤ�"ip����H�HWj��-�m):o���d�K���Km��u�ϑQş�s@�&&#UDY��7hԩ!���+�miUdN�[_��boj?�f��{�L~��g'����6�K�j�$g�����8������܃��m.%m'0R9���z�C�p`%5ya�~����<��͙�.b9<�vF
�O-^�EÂ������V�m��W���ǻ��/6m��R�T,����#�]�V&h������`��%%(']���z�ybѰC�K��;=>m�)+����I�%?t^��5�|��T�R��뢗A�	Ko�v��}Qʘ���=R�����qI���p����}d�&�1��,�'+�U�_��vd��J�I��G����Q�~LbśJox=�&@SՑ��X�#(�saN���@�Uޠ`b=W���~G٘��ȟ�燺��u�Dr�i��%Kח�����f��;k��f�ӷ��H�\�å����L�ېj'�O�!]���%�} ߙ��m�qTz_u������3�~�UY���h�������@���E�F���Ђ�b��R����{oA������,Ƿ0_���X!H�g�ďt6h��]�c5_�8-���;���s%�^3J�s��@Z�4]�{4��^S+Ɔ��Z�rC���Ƴ;m�o����"	Ok.NAI���-̶����%�,���X@�F�4g!�\8_��
��~�����^�j�3R�w4�t�Zo��%+��OԿ�,>.�1d�[h��P}h�,�l�Y�Z�?��i0��ve������4�m�C�̭�7�oLeK��+�yz&
�}G��=1���M�[����2H}�J�(Q?[�������3�	�;(F;ȧ��j\�6;/�
���9bR��D�O	��
�8�ծ�o�$<�@?�F=������m-l��9�i�NU� ��p�4\i=t�u��KVTDl����M�,�4P�ʠX���ٜRXWT�s�s�c]֢�x� ��*�c�O�Tp�u�7�Y4W�c��+�|��.�0������av�"I-.S�{>l��ncQ���v\���M��^�qU�n��ެ�*�݉U�|��X@���v���M��O�V�7sK��i`�(�R���3M���{ӻ�߬��m��	�����<��$��l����jx�s<������	�]����.��GT�TION�cf� �	%̚|�8��gS�G2���7 ���a�M��d���M[{�˄FYa�7��ŌR�uhݡ"b����v�m�)���[�O��;x�~�=�%�[=�O��J�%B�z�oz���cy�lxC*A��l��g�x\���?1����2�O~����jA^k��d?��,m����ڇR5^Ƶ�m�']8:�}Kx�@�:����Ѣp
�:0a�_�Uߊ�'�����Ȩ
��((�Q����b;�!���􌔢.�h��|oz����Rw�J0�A�H�'�/3�L��p�J :�bf�~�[H����U6�D-��9�AߍM�)�@$&���ЬOtp�_�� �Q���O	b����V�r���b{�Y�P��6�"�x�\������yݑ�~=�	�z�q��X�4Lj����U��?�%-:bft�q|;�8�7;ZӉ��r�ґ	Pi�����rOE#3�E��r�8���I f����	�p���g�	R�vp�,9���&&4�����Fe����Z��	�<�,C�&��b+��:��@�>�A���С��"�݇s��Q>e3���,��n���/���,G+{���Ji袽��	�x$*b�L.�[V���'�б6÷U��-�5:Ql�1-f�Fk[iȝ�>X��L-����Ď��������T��R�٦`j��=!�[�6Wt<���)������E��.ϰ���Ͼx�N�-��z��5��<q�(!�|ڄ�X}	 �d��L�J0S�'R�]����TN���lt\灨JϤd���O�m��p�(��������  W��P�Ƒ�?l����3��c;Y���(qCCH�Ә���s���/!w��@l&�8��]��s¶6�aB��r�?/J��:B�&�]+�h���s����6�[��8�9*�9�����h�R�%��sR�E"�rd�7��>#�����1��u��em�򧉠���j�X�-��5Y��{m���zuQ�z�fA��1��	����C�?�ŝ��j��Q�2���5q�M,�Ң= ���7��	hQ�FOv�����+@e���=��K��k�tZ�	'7��)'ʩ�l�=%Ci�nDl0� ��Ա��	c�?����Z��fptjJ[ħ�!�_�S���y�JՂ�pMaf�Z�a�U��5�P�46�x���Oyv��g��C��sm�[��X�����4,��9o�v��ɛ�t���b(�����{9i������^�'���(%'�>��Z��h[���a:O�r)�;�W�3S�����.Խm+��>T5��O��������P��D�K�:�]�E~���ysR����.[�RS4�g�Jr#	/�Jg;������'ؒ$�V+EB8y׳9��j*�=)�������KS�+���k�u�ld����\O������4+�m�<UT͊��t>7�@��?&2�4����H�^P?b�G�Y�S��H�W��RՕl�a*��}B���tD�G����@�����Ρ�f�̇f5������-����ɱg������h/"Z'�rM�C�J�����W�m�'ߥ�S�h`����Q���������︾H[qx��"�t��B���7Ϊ+f�� e�l�0��'�Ҡ
t_$���?�b�������Qah&�;���a�{�Ⱦ�@���4�_Bm�x��2q�'*,\Hyn�W|e��'� r��7�-8ԫ]t�V�t�'�k���f;:d��r��W2��Xw4���~Z��$�BS��@�s�j�rGJ�`��v�Jop^�eG��+����)b�L���"k��ޞ�eT�>���%�j
oM��G"���9�&��pB� &�|���8<�P?+����4����T�vb�d�k��^���%R8���!K�6���Z��a�%�p��c�����m2�����Z�����6�k]s�ZK�A?p����Ӈ2>��"������XN�]^�)����<�������$�E���a`��+����y��@�j>�hpV|2���7�ow����b��C��Q�'�h�<Z�5(�M��k�2�fk D,�*=�ꬴ D|b{����u���޶>�\��_��꺀���)Tl�uAl�<���
��SQ��0�韭xe�������uxւ6X����yʻh�~񸍷��0Q1Ը���cXNC���1�mP��L��K�z6�OC��4P�������h��^�0�u�£��߁zᾭ�V����o�ڹ�����ԯ��Y�,�fB�}���o]�b�"���Q���]���s�<%d�c�g!����ݍ���SI�1'�d�fk�l)��ȋ�~�~l��V�4b�>�!�����D_-Z�eh�A݅L�p݁f��pĘsAg���m��3������-��q̈�_cʞ�:��z����:�^.\
h�*_V�Ǵ�k�8OR�����U<ԕ��C�C�xr�9�;��!��v�G���L��{�Lsr��@ߥ=c�`��0�v����f�|.
��"�?O�ؤ���Z�}.c�~'��;7�r"l/:�-Hr#����v����S�D~���{�=I���e��+d��'�*�;��(-[4�H�Q�(|�zE,q�?`��7��(׃��j��^	���3���i�>ް��u�!z�l�1>W��qԚ�����j� 3�������^j��,���/]����X��_�J��DGWu2�*�1Ol�����c%ݳ_���Ai���"͚@����2��c��q��z����au&���/d�[&��%���lQH�����j�8����4������V��@Gv���!2�J#iiP��]�����U͖k�?y�m����ͻ-��J7@8%ï���9�2G���[Zw�� ��"S�h��C�%�b�oEw�z~DM�4���uǳQ�5����
�y���qV�ŕ��/�Da�b�x�芩\5��=�_���Oc����b�'9]Rv�a�҂Y��Ώ�u���8�,f�����3L�n��.�/ �)�in��qn���#Tq��� ��2����L�x�ҷ낖\�V�̄�JaBv��1��2����+x�d����c#ii #6�@��.\�6Hq^�eLE�C������B�<� N=�s�������z_1d1fX��J�3|����8ae�	tf̧����_8�����<��������FlfC�G0��C�v��J}^OҘ*�Fӌ ��:MX�k�!/�c(M�n4�N�2V4*�/�p3����|���3�B<��O?�L�@T���Ho,�N�Z�B�Lh���2f�:�����|�
W%iI	]1�#��[zj��f��A��2��g��KW����n@���\'t����, #rH�fEH��7P�;+Şv�m	�B������{?k�4M(,�{m]q-y�M�R��<%+p��!��Fߠ1�j���bR�k�/�#y�?�#�#b��K`HǷ,���#G���������Au�x�L<�F�D�#=��
���O%)�pҼ�jtqU�R��{iUX�Y?��i�qo���AΓB�T���;[(�V�N"���&C�RQ=n���|\�x�C�G�!]I�k��h#��@�_zO��'Ч{J���<H4�#���	�FS��wh}����Wo�(M�YB���i�F �#��o�������&��KhRȒ�x"��l%J�ݨ掣�'��]!���\��$���L�G����/c-Z�,�pH�R8<�.U���4da��_��K�.Y��u(�����[t�oXI�2i�թ*�x@��S�LEj�^TnM�����*��}�9��S/~�f�����U&${�'�0d�z@��p��
qz0�~��)�ʾ�2/��@O�ͯ�����Ҍ�H=@���i�Ǭ)j�&YO�a�W���|6����/s��Qn��黒�Y���Z�y���~�_	J=e��k���F���'>K?GiQP�(�L�����~<oqը�F VlŻv&E�Ԑ��9i���NX�ߛ���̔�)ܯ;����Ѭ ;��0��d٩gT���^�E���p8)(!�c�ޫ�]�\��I���Ԅ��?|�/b�W��M�qQ���g�s g!G[}$�:z{i�k�p�����i�K���#,���N�H���'���S� �1^<�$�]�,�ƞw*i���Q��!��:V����\GT�� ��ɶ.<����'�[�+�;��2B�e���7v"Jw;P���I��].�"�SF�˗X���L��D'�<G����U�G)��	�$�RWe/��]�K�Yb:}3�k�)w7������X�71���8��c!c��F<�b29�'k��|\ɲ�N�2��ws+[9���z��X��%�O��"��X%V�=Ǜ(_�.��غ��w9M���.`%.�;����O��nx@g��xn����k�媜]�>beRѢ,���ݕ�0_Gk�]������I�	y�$��ˡ,p]��Ӕk;���f5�M�=�<�R���K��d�����"��q���K�5A�層�J�J��"��a��z�T��i���g���jg8����e@F9ѻ,���NR�jF�O|�G�>���ȹ߳۸!���7���kaA*��4���^�U��E�=�?x�Q�ra���Pk9��"��J����{٘���Z��\���D,��+�؎����ܸO��i�v^�^J�4��]X]�И�`�oR�_3��$k���x`:�8��#Ojh}T�El �8u���%��vSB^�����9@	 ������jeV��R�]�,��Y��ZV�ia�����"ױ%Gg�U	ĩ��-ݝ�q��;���e��iw2�uSo�5�`Kno���Zjh��&ŀ�wRK�+۷ |q8���ym�O���`�s�,���Z�����q�?XP.S���yN�R�[��5�S�N�V���n��˛�z�^�LA}"�"^�5�$!10MkV�z\��0��w�9)�_ײ��K�;�ךA~p(�� Թ5!�b�k���,��V�����
M��((/	�\����f0];�.T�I�+��j����d���[�9E`��\lR�ӈч�X��iv��-E�Cı�������w�k�@N5ɬM��G��`/����6���g�G����E5���R9����J21�䝂��C���}s�5uR��2��C$󼦚~�Z�����5/���H�=���i��b�Z2l���L��f}���⋺���$�y���&�^0E΋�{�P���H��2�z�3f��_�l��Rǂk��L�e	ds��r
��4l�d�AԅͰ�<��7�;\?<��+�U����k)9�#l���5��2�u���t!�/6�p��C9�����z��6�#.O�,R�ϫkRF���
ǰ�U��V��pY�}���%���9��0��Bg�|+���	1V���t-��1�x�c'����av\#rK՜$瞡sH0j�?�`2v�H�;y�F{ r����kV��]�����Q��C/�F�����>t�0�'Ǡ=Ҍ"��t��\̳J�'�N���E�ɡ��$�����B��M��P����$u��c]�a��NI@�kg.��.�u�u0�z>�J���'M$ދP�Y�]�B�_u+l�Y�Ua'v�qo����gqöz�d�6�m�z���[r%ZW�'�.�
�k7��)�E��!#�P?w�������J�N�:!����ѽ�Bm�3�$��Y`�Ⱥ��͌�.�w�f��%P���:Y��Mͦ_��<�ޣ*�-`��G}��co���@�]�R�a:�|N-���ew�n����]�@��"^Y�j�Y����R�y�Wl�z
|�X�سD�iH���|ѡRh��9��4R��t3ے��6ՙeT�2��,�"�$�='�(ے�:�'��Z�[��-o��ꦢ�Mf���j��#�lS��P[i~��`����Z���C���ݑ��ɀ\F�I	vg�V�X΍	R���~���B�B�m���>�xa`�ǒ��U��ʉ3��^:5��i1�8S��+#"u�ǏU�6̑a�Mˍ"�4��$߁�#��(i�#6_b����O�H�KT����.��.�w.3�ՖmL�-8�𡆜�d�
$�5����8mڪ�����lsu��'�o�R�:��P�)v�GN�R!��M��&�kŨ�D���De����h�-WYX&��Sg�B��\o�=C�rΕ�ɘ'l$S<��c�Q��ma�i ���������7�@�QҩkQd�k㩈�i9=8XQ��b���3Ɏ���b��C$GE�NXI��s�R=;5p3�n��c��~/:��ņ]2�V��.2��9l�ڵ�e��[�N��Vl���e�����^g�'���Q��&��}�^��v�=,Ɲ6'/�`�BF�V�����N�8�mr7|�@���@v(�}_U�U���j��S'S�p���JL��&�q�����2E��K����4�������"C����B�a���y��r�L��i )7�z�;����:I��Yr1Äox���+Ru_�k��y�y �B�ϒy�������=w"��Y��m����Bh��)�}e	h�&����g�B��<p��# [�F]�`mY4��^DD!I�}�0�Q���3-��е.[ҋ=Y�X���E�E��'w9h�`��;�s+��U��C���^�N�{���Q���}՛�M����)�.���e3�%/�� ��.��Y�56�l��~T{��ˎ������K���J�צb��T�8��!A��
�e��v!�h�Q��YF�����/���4-c�^��<ڊ�+p��/�6QQ6t鿲��}8gt�zf����@�`�3_@Qu؊n�$�T�Yȉ��J5?-�0�b�f����I�\�D�`C��>����,����֙�K���h�LI3i��e�5�} �,�'���^�l�l��T$�[������r�[��Шz	�Hxy����Uԁ��W���y�2�kMiᇣ��J���N��#���$kM!��d_q����$�zB 1O暪N=@� .B
s�%�OF�\&J|�ۻ��Z�o# �C�ѓ�׳۞�N�32��V�T��"�L�G<��N�6 /�K���{}|m�F��O�8*��Bg'Ӧ�J"�R�ڑd��'��~e��Sz�|���8�KБ%�������jID�I7�A�9=#i�\pFeo�v3�Ҳ�'��y�n�>pCz���#cw̵(����쒫���A����.(��x�4����=}�+��܉ߝG�{��\<�#5��t���r\EG�߀{û���3������|Q'�}�	���7q�i�^�o��\Y-�Q��U�9�׃��i����s���X��a{=4�KA\L$E���j�ߺ���}u��-u���w|�@��H�0+ϖ����E�.�千R��3���O��n	N	/�����xP¸.=-��/�2	���k��_��iJL/��}�70��X������Q1,�����H'�W�Mj�73��O	=6�H��G(�t�ƿ��������o(�Θ�P��e]���tK�+34#M��
q���۫�7�I��k����a�r���yG�LZ'+>4?H��,��`�à:c�/��(�c�4(�4� �t�VVl�j�TB�@�]/����U��
%7h&/�s�Oз�2r}��$�tx[�o�y�
<*r�:�1ľƶ1X��z�)h�٘�����f���%�T���
#!�YB���Utڋ�Ϭ/�Hلy`iu"
�_��}��4�!�s'��O�����-���,���-w�H(+e9B�߯F�v w=[Qĩp���� ��2�$V穜 Ѷ�5e	�� IOR61�):���V�Ol��F
?2k������ (�зo,B��?k�D.8`i#?��}Z-�ѱ�Ϡ�����'��WqyO-1ɣ�r��v��/������p�i^������U�@�uSWt�~�[��/|J�kʬ\E.���yO.���f��w��AEU�~O#��t\OǗ���M��u�3 ����K���˫,�5�_�tL<v���I�qP��KG�����[�o��M�wO{�ͳZ�?���[F�P���	'fhmy�oMj?�9(9�L��P=���ז������i��Tf�!����/�d���D$n�5_�N���.���UX�ڲ��7(��JO������7NO��� P5%_���f���d��%��kT?�GM��WT1�9}��B\���ǈIp=����J�U�Y���樖�K�9I�`�>T?[�F�Gp��q�����^�X���=��ݛ�8�R�zT��$���[*�8�U��1B���PhW_�5�n��wѥ�!�k�~�lC-h�)a�Hl�s6�obX���v�,�Aw����I��w�Օ��:p"/[�{�'�7��Z��CH/~1R���6�.	��yd�ov�T�Za0�a%��e ��9TATNk�_�p���i2y7�m�E93q����Aҙd�?!$�7׸M��*��sMR�K&����	�#]������{�����3"�Ѽ=�{+�r +��K����'�nK_��볩0ƺ"������R\�ac��q/3�x�β;u`�E[%�Ęfu�v��d�fJ�=���XG�A���-.r:VB�D*�fBJ m;��{6�Hg��W�}l�ey��p>���A�˫���N�u<�/����W2A� ?)ּ2���r o����\p9"�%R����t%P����ɟ��}X��Y>	A?zD��C:����=~�;�8Y�g�&I�p .�Q�M�����=��R^�[�W���~kpUOx�/������|�.��
 Aط�aɼ��;�O����0x��A��"S�
�Q��dT��m��/�;z�> ��p�c$�+OAs{����-h��7�.�S���.�,DI�,�����.m�Ry��-S6xa>2�T��<׻جB
�����o�9���8�.�,*m�o�z�_l���V����\��	bx'�5���"�HE�&z3Y������+9���8�Ij��+����r��rK4�1�5 ����6N��$����	���=��Q����?���N�
̳Bgb��1�⮌#�܊q����=�X69�|}��|��%c����{��=�L�XEa�l�'����q�Jȧq0��=��̽�I_�<FXJ<~�ˋ�j}���ᐼ@'9U�	�R0�m�M��o0`�$A��z�W���r���3N.ONIwʂJi�.���2S~�6wr�x�~Qt^����)�/	�L����)�aC���&��inTш��d�tg(w�
i�*z_�l���֩mG5�ñ��imN�׉�@���SʴG��]��A��ꠖ��Ŭ�d��tB�G���cj��MvR��