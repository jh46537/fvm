��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��ߨ�=�]	7�N�)3�M�Ρ� ��B
�i�k<֐�1(�/h�"�+r��ҏ�X�fИ`��6.[���L����Sg�$|����x���
����v�95|b�fUw��e#���`r�|�QZ3E�*��e$㩥�֢H.���a9��[��}h��P����{7DI�y*��f`�K�>BW�{�����z��<�	&u2��<��q-F�zB��0�t�c\��L��U�Z���T�u�o|^��G�)�=�d�so,�yr���o�L1/�%�o ��)X�A��f�H9=<~�/�f�ԑb��ޝ��X����3�5�_�O��AX��ˡr*`�}�1	��83pPR]�B~ƫ�ug�D����2�9� �����/E=4�pzD�<QCY^��}h[
KV �����{��g$_�_@�6��F��7c��m^�<E��v����|K9$y�jx�~8'�}�ȼ/�r=�w·��}[#�p�%�
����6�u��NY_��^]�%�Q~�)V���#q�ք31�hp�~V����A�hw ���p��R�׋m�N�w�t:)&�[��|��?��Bg;6X�Ʊ3�����u`�x��eAw�2+�����ï�{u���:���4J.��5UA��qj��������hg�T ��8l������Uu~+�6���%zxm��y���%CYL4��� �+>)/��6NQ��'��Qi�����=�9.�%���8KB/O��Y34'�bw�t{m�����1���	hg;�|�y9�/u�J�v��N��/�ñ����W����z�,>y�r�p��i����i=[�����(B_|�'����>%4���"�1����JDQ�fg3
��B՘~��\=Q]�dxCk:�|N��N����w�~�S.�FlB�	9Y��,���Vx��A�*O/vܹ�Y� �ش���,p�Hè�=cpL��>`�<�>�g2<�~����� �)A ����ƴ��k�|�:K�5��<�TG��乁���I�3E�F�������_��r�ܾ$,T��%0�>�I�BO��3o%��=�����}f˔=�j>9,@��M�{��YW��߂�<��x���8���:AS��|>��:J�oj�2�r���9!�Y��6�x���q\N3��?�lw�}o�q?�H�$w�Q>~i��M�XQ�ܗ�@`�w]��5)���j��kR��ԷBR�r��>��|0�"B�r_��Ĝ�r�<�3�s'�V��~�R��G�j�������H����Xr��3�rv�C�c�����(��~�^x]8K�h��	G�:�r��H�w7T��M�rҙ
B�5��D,�8R$R�ڟ;�Z�C���Ʃx��)��֔�YӠ��;i���� �� ����	������U��b�j��'D��
����[��*'�6�4L�� ��������JQ ��	]�aZ�1igF�񂫒�	��v�NN4yv����܃��pqNz����E\�P� �_-Q�Ă��+�%L4w'�]\����r`c�u>>��ʖ0j��+�Õ���"w�@��7�uR��G����jB��%q3&�e8�|+_/8�	nu�=+MHDt��QW!��;޺qCE�Y���
�@�W�l�L�O2Wk(���Z`���VK}yN땐�����n~i`��{ƙ�3�~�\�A0����Dc�%}ˎ8$α��,�ѩ!�d���$�����6
�8�����H\�H���(\��_\��X���c���P
��R���li��19R9KY�:�P���4Ucz��s]Jq��.�L{.M��2�@4����ұ]�U��%'��_���y�)Z����UC�,��@����f
?)M�Y\�g�kZ��W��bw:��oN����%���m	�(|щ�����-5@O���0bo�_l�_ZѶ��˃z��w�����i����v�}�#:kb��b8E�C ���6��������1'�V��?�L��i�k;?~��?w��������v�f�?T��T?M�Ж@_�&�pV�,�-J2u�`�~_����6DNp�l�B�lVϱ@��تW��p@ۢ@�(�]N6s���Q�N�)��)o��oD2J�*[��xH1���N!w��B
E��=�~���G���aI,6��;�5p (���R鋞��EʚW�e�2�*N�hs�����}�9��v�- R��An[�v�+�y$&I�)�1L
?�'�Gy�S��֡ժ�p�g�tw��v�j��9�[�&�^��/�_�jVCɤ���;���#L��!W,j
��2����,�oCg"J�?�xrt�
l�]���Շ.ALDh�Ӊ]��l��B݌ɠ��V��j�M�~��v�z~]�$0u�9�!��!�����������^]<�-�Yb80B�Sk{�a�V쑳V	O�*�n��o{'ռ�E�� ��N��i�C�e�Y���D�������2��z�8?�X�g!�c�0�%�_}&�Y�,;`he�j��k�U_b���O@�	�C�R��'��G=O���g�,��]�xj��K�yaֳE�Y�v� �	u$�{�Gr��L��r��++]s�|������2�2�]�{�]k±��	/����ωQ�Ku�lR$(xm_
Q�?����Ԍ���>���.�T�����w��	_ѫ%϶	�{=RJ��$�1�v�9�?A9�H��1�JK�֔��6Q�����WS�B0��Ks�lh���Yf�P��6�/�vT��:7���$UE�O;�`݉m<���D�E�JgA��D���&���R~�	�[#��=��PV.��Y0��֫��u���H��j����bwc���S)+oT�7A� 1��{v-�3ĥ�S��I2aB�56��+�U5ׁ�$k��W4���Ci~��w����⛭`����gŚ�S�Q��}x;��IO�@�I�Z���Lp���be�I�J��y	e�J�	�;���gGc��b"AJ�l� spVoá�v�7o�XL*����bݞ����2n�Y�@O����F�3�0I�W7�=���e��	 �tL��} �x�js9@�MS�9���]Ƹ��Px;�<̮��D`.�/��{�'ު�]��Y�k�K ��J��E��'q�6.7�����f�2| �k�)Sϋ�2��p$ˮ:�݊�_f�'_�D0�W��&�2HR��Cd�N ��b�9}��+4�FN���C�ڀ�d�[V�c�s�S,����C͸v�F�n���$"<�D�:8�c�Ǆ�r�����8��S�,�I;դ�c�N�,���wϻ�17P#�r��H��]E�v0�f>��;|�W�űҧqlה*�\\�6E ���IvM����h�'�	f�xk_+r0�_e0�`� ���1����+�Vj/h�Z�v�k��;�0|�����G4�3~:�(N9�g郏���pt\v�uX+
�l��!��f4B�� j09�ED$�]���Qׇ}�g�L(�O�,.j����ؤ��	W����5��i�)�W4�v��@%���M���q�	��i��Ob�ωd<��*}�@A},�ڎp�A��	�&��R� 
G�Ry�P"�d��6r�	]�@���'���b��:�&۴�!Wj���v�pH9�6u���	�-m&�b�����RBa.$b�1���N{��p��t�b���L�\/�cڼa�0��p@3�0v2t�HU�����p���#D�~Oͨ�k��ɧXH�	L��;��5Y +��(����$���X��"���0v�T�X�n��u�tJFヒ@;\Y�&=�~x��77lq��F=5�q�uMҮy�H��뀲u�#s¶0�K"� ���׽��O㜘�3:�V��3�����&"�o��,wE�^$W�F�"c��R�h����q��*|�!�5W�(!QR�"��;������A#�/(����/�ޏ&��$��./ZAP9#Nv �J����.��֤�?ߘ�j�$�T�D����=E���Rs�yt���S��9�eA�Gܞ��8��U�^(9&b�\���wja݅������D��X�;z��%��`�س\~2���A�R�9CPji��kԌP Wd�r�"	لIU��Xd:%������k~��S��ĕ{�T�.��YZ���/��]w��hW����]��,ΰ[���%�"O�¸������}69�k��h�O�D�B��.L�jj(��re�[�ff��	����e�z�%���Zo�����A��`�ޔ��f_����{F)K;��܎�JU�;�>hrF���3�+�D!�v0�,zK#���)�%.`3�d��@�.��������A��M̩iTpA�R�o��U�$�U ���Zʲ}��� �mt/�n+������DE��+�k��M����_�XeN�/�Q[o��T��D�;�Ji�����ȋ��Ĝa���Ƶ�������婘Z�V4�N�[��`I�=��d`xs>�Xb�L!
bh�砐�Z϶v�ݑ�M�{��Ȟ��������z�2ܚՓ�5�e�5�Qα��CL�܇!|��j.�i������C$�1��a��E@C������wŘ��ǆ%p0\���jf(UiBu~U�}��Y��w�T/9-@-��I5n�kuA{��"A���#1D��f�wJ�v���E���	 
H$I�#��fL�Jr��)������W��H0���Kj�xW;�ȮttO�{�
z��y����PA6IV��J�bp�*�XK\��bm6�Gk�F��PC��#䔙�ն��ˢkl��4�ʭ�S�	�����T��'t�)��VdO�i����e����@I,�BV)�q�J8��A0�N4V�'�Jdga��~+�=;y�=�UR+f�zeޥ���p�L�t(jw��'�T���n�]-�7��TڷV�=�_Af�>��"���F��Ւp*�����'Ie�LY�c�X H$9D�*A�}<.��sfvHñе�\^Ή�=-������[���� �\�����2�͹���?������M���5Wm6�e�֥��L��Pw�ш�x���۸sE���d\7C�M.�/TV���a���B�)�;�Z�i�վ��Ypƍ��E���di�Ώ	+��$~k���Kֈ$���f�`k
@��x0�҇u��wd>p�^ϧ�?�SěT�L������gslh\y��/ �}g���9h!�aV+�HA�*@}͈s��i��_�m�� �	J*+�we�"K�+HIW?eoکB�i�ؓ\=��������_zmaѧhc[*Gk
83t������E��srcZ�f����HGO���Ŋ��a��%���Qf��{���*3TԪ�8q���� ,��h�a��e�7�6܎�R���<
3IF����VGA��f�r/����.�X���·�3A��8�_CV�m,� ��VG:��
A�|L�t@�Q�F��
��Bt�x�8�m�n�N�kZ�[dK,���� �ې�0ll1Ͷ��˃�<���O�K�!M�(�l�`��.b�
�Fo�:��Õ�2��!�*U�g4��<���&\E~�
�3�>�;�T@��nİX~.��tݦ�Μ�lV���.����Ū�<�p�Cq
��F�%m�!��F�����d�I�X����Fb�a
�5�5���@�3d�H�IF�ŵD��q����x3�쒯@����ܐ�]v�;�7j�I9��,t￱�w_������)����k; ���re�h�D��$5�Xll���硜jB�-��ImX�>m܉�~E�>;�';P���~��+0U����ln)N(g�%�*�\��.w����j�oVDuZ�~����o���v+ODz����|�0�tjM���|D���Mַ����Z���}���C[�� \<��|�E�" �t�9��c��"c�艹�)��c�9��v� GA����ȍ�
.�;3ggY���D��/�Fv~[G�����J$5c �t<#���Y�&}�}w�_�rX�)����H)��{�v���7G��E
C��.n���-D󺀳8g }��6����љ��l���=_^|�$B\:t\6Ѳ�@P���ĨB��vb�ċ�L�!@�R�,�#u��1�Aw;���EK�y����/~�����LBo77{�%a�q�*1��;���r�l�H�#х�ͳ]2?n�0�wo��<��;iU�̥���E�6L,�Z��֬M���gjו��B:g�r���F��պR��$���Ƽ�e�����trFV��{���<
A���y��$�� 0.O�B ��{>���;Dn16c,~1��h����K:pn��K�<��|�ϼ)ho�T�����;t���/$�'��q�M�ʨ�:g��q}�"��3(��r2n��������* �d������W�[k�cՀ�N�;��Lΐ��v�q��Hx�U��	B��Z���=&�Lf�|w0����x=_U'��&W{��Ӫc�f/�M����4z};�C�Z�I���R����Z��V6�j��2�R�Z\	�xv[J,YI�f�����n�̹�+t��d`y�Qr�H��n����:`�����\�	$�|��t\7��2�v>�Q�Zfm�Qc�$Q`�^�P �j�]8���&<r�歴U���qa�l���Y��ŗ��Q���Ћ 2Z9���5���$�a:�c�D媈�ǜ���*������r�,���#�kp�����7\?�G���]�*iĒW×��&_�*�V.��髕�w�{[����.c$O��n�C12b�Ff���[?�JyR��E�c�鹨�W�#ur�A���ul�bZ�~� WHc'��W�X�ߝ��3�.�<(?x�E�F$�C_�\Y�gȤ���� �V�	?�1Z+7\��WWrdi*���:��O��y�)�8ZL	�%T�����4��'�;�Z9.�q���^�Dzh�1$�r��d�N_Sp��Ԕ��7: �T����h�t!E��5?��l'G��񦓓e0rI|��n�!>.-tؐ��e�xM�Ͽ.&�Z)-H��Nϐ�U�̦����Ɋ1�ŝ�x���6lx��)W[�]�N.�{|�~�O�F���NoBwv_ .l�4�4���!e�ȥc^%����Z�A��@���~47*���KިsVV]�8�1�t�㷿t�����G�8��#��O���Xf�|G�����ܩL
�d��U'��U_��ny���K�2O�F?�v��4�a꩗����jW�@�(�[�w�^<����Z�C]���Hw;|(��$:]q�~����Cz�nf�M'�j;�Q��hO������ٌ>�QǇ{g~��;�I�f#�gOE'!�؜�c��_��7>��|pl2 �юT4�� �R��Ҏ�$�@|Bޏ"��@�<T|���08�da/0�JeO�PJ&ɵ`�^V�ae%��"�3z)��7 9(25e-�-�ߩ���5�s�������j	;yL�����J�^�n���KC��Z�,9��coN�0v�	a�Ă'�ɜ�Ko1�sr�8�3�B=Ć