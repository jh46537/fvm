��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��)Y� �1�c�{�C�9	��܈Y!����lJF/C$d,�V�<�.
Ւ�-!S�h��n����X��ѢS�R#`�ǗG�ݠE^�^HQ�JDbs��:��y��I����@�1��'�1�Б�4۔�K�s�~�Y.3�L���G��6���<\�.�
�m�܇��Q�o�j�>�o���L0��8_����M5ZN阮(貹��.+z�9�Y�]}"t�(&{?���s3�!�ii�ߎ�u�+��S�,�mI�=G�/I� -�Ez���xp�󴽏�i7s�[��9���?�i���m:eT�!��W�T�Ì%P�Y�M7?(�V��ē7�=�@	��$����ֽD�(S٤�����|>
LmC�r}��?]c���r%����D=�����h֎�	)C��k���ˑ�;�,E8��5�'��竣sC������O�X�Ur��p9��W_~{����YF��:Y�>��{�hR�Z�Z�p������Ot_���GPrL���.o�����[���G�0��w��k�nf���p�"�i>[.ڜ���"�9!!_[�=Q������˙��s�?���U�n-�;�����ϙ.q�C0��Q4շ�kI�5>�E'h�_��UBE�Y;&V+	�������J�t4�:�D�n��9έ�l�-�p�ߣ?��ܨa.��o۱�DbJ�e2Khܼ$��f��[�T��|[q�a�4�>^T���C����?�]�bܟrO{<$�A�90\����T����J��d��w9�U^9�-[�_A4	�+�Z̃��ƻ�ݽ��n=�1Ԑ�k���D���)ـ҃GՓ�?v �ј�vu�/,�4Ɠ�T�&�+���Q�>�=�X�btvJ̹cܺ�����'I�!B�b$��ޓ�<��*�f�Ly�%fT���c�1J�9e�ltj+��%����q'���K)�]�qvlE21x(�K��hg��s���!��$HB��i����@\8H1|�|����$�I�}�\/yט�!<�(�����L�-���`w�P�+C\�L��v��%����@%$٧y�Th�;�<z��7��l)�x���t��{m� Xmh�����p;��2�B���V������]�T�F���5���X����W�yA�h���6�f�"�
��E��P��=�!ĺ@p_�Yl���W�I�	���"���B3���[O]/wt�>�o?��T�:����w�*��(�!�@����裬8d��p5^עt|K).m�Ix�=i��cs;ջ-�K���G�Oޭ��H�;�sV�"�"ݟ?8�=��O��Aɰn�ʀ�Ok�'6��9�������. ћ��}��/(�W
�oݬS᪩>����8�.���z��e�o�U��6�MN�C�GP�*�Y(&�C��6b���4�`�&��R^?V�l�Iw��Gt1��m8t7D�G�U;v-":hm�k�9 ��CKqf1i�<���y�G�I�'ጙ
hsDގ"�$�KW]�"[P��`���*s��kP�m}9O�1�	�EX��s��̪`���:�ʝyܲ�FM�u~v$�Ti1ãYw~� ��-��Y������8������A"ƻ3"�2���LI�6�T�6O!s`�+Ҡ�1��^���z�Q�z�;C�W���ఢ����������S���\��
V�ǯl��խ9Wi�!��Ph���􅹘=T�:��p ���*�	�Y� �*h
���D�E�F�7��X��P�*�1��$wy�)�G��(�;GŢb�i�9�葢�#,����}`*�PB�[�"�d���	�T���U��ɺnXU,�u��K��x�I^[�:A�
E�0	����W÷�22o�G�*o����ԅ%�G��D=!on�Wߋz�%iiu-�roC�X'���c,�y��Dsd�/���! �&��2bM�1��+����捏�y=:����T�"ap�5�G�1N��e �(;u;� �����$�Q�v���´���pT/L�p:�=B���A	7u�p��-K34����$Jvdc1�`Ъ{z�h��8g��`�3�f�fl�3��j�0Q�8\$w�h�-��'�dR�Y� Z���5E�,�e���¼��8ξ�V�	a�h	�����`W�fL�	��!r�������9^���F(�x��[���87��<� ����73w9�?�}FO���<��y���y�s#�����G��7ҽ�#���'o�`��H�&|����C�n�g�������'S��kUF�+c9cq��G��"�h2F�;�=����A.�!.��"#J���rAO�vF��S��!����6�����6\8�	{$����Q"~H�>4;�6���2��tp$R��L��D�&�{7}v0m]%�fH����[>?Q�x�	�4u�ǘ ��7ߪҬ���>MZ!�M�^�8�����c���R���n7U��D���H)��DX�	�iJ-��M{�&Bc~�2�m^�dɍ�o�j�&��N��YK�+]�C�|t�sf��Ц:�3��$�3���M�Q�[Ϳ��n2���QƔ���i�P�n�	��=��m���"��s��:��L�E�c�
��G��%A�������WƷ]�= :��c��*�-�:Ż�V"s���&�	"bA�����Ro��<j�̈́X�yV >����p��fO�F�ϕ�Vpq �(����z���j	�T߻@��z���F�-���F	��d���2����nKG�nAN{�s�f!���@�`��uj7D�pC�>��m"�q��E4Fٝ�,w?�y������Ӡ�t(=�A�A��ٸ�z5�Ú�^%<�HF�G��T��Ao��z[w��
o�-jo�?Is-O�ƕ�j�vrfxԗuc�ٸ��G<��s&���+�������2��Pݸ�o�S|�W���6gVm:H��u�ڠ�g����4�6�3�֊��C�n�W� ��Z��l�4Yg�O�Kױ�rƶ,}`�b~xݽZ<������N�ZQI��ɮ�@n�:�Z�d8�Hv�Q�)�l�)jպ<��$�������e�qfd��sL�H[��J����=Y�HL�u\ʝU �St ���7��BX�H�!Q ��(h M�Z�纽T�؋���^9�J'���[�N*C~"����X(��W��%T��	�8���񪃵"c���f�.B������9��?�J���P�h4t�R8�ƬH!A*3`����N(�W��k5�[Xwn�Q8M�؛F�rIc�sq��0��[��D���\>�K�٘z!���0��}�L=���K~��%���÷� &�k�'���)<F4�A�:����J�������wIBڨ������@�ر�,���/fd�(\J>�u��P&W���6�������q�S�TG�)��/���zDܿ�mJ3�}�����p��2l�[�K
�!�އ0�(.���c��R���:a`��2�[x
��5���4-�Ok�{���n7�S�`U�=�f�sQ�pQ���@�w�Q��z�!?�v�x�|@v��(� D?q|>��Xu���Z�.���j����]�ۉJ�7gh�5�$š+��
��}�TK3Q�}E��Hq����(ٮWڻ�J�#��#d�jd�%����V�
Ӌgd��w�$f<J-�%�\:��w�2�s�c}�Su�[�_��!��i,ac��E�R)Ɇ��3-��C[�
���١�v�)�\"��p�(���bW��Q־M�E g*DJO�I���ں�/�VB!"��Զ�f���;�|s�v�㍻�����D��|�\N�#"Ɇ{ٙ�N��f �!����?ϒ�Q�1#�0\O�t^���;���|���+K���ͬZ���R��ط=s������i'Y�O/֒Z�z��/�����芩*�G�n��9��'ú��S=���,X�=Bf8� ��$�A���l�i����ģawU{I��wlbnPy������ܼ���m�@�Z�P�{q��P�N��k3�X0�n���D��&�*� c�/8M٤%hN,���έh�!z��iR���Ppѹ
�����@��ǥ �~f7�J>�%RmE�$ �M^R�c,N|�c<�]�2��0�S���^�a�4D�+��+C�O��i���t�{�i&ԥv�}}N`@���'�4_�����}n�TP�����
�-�fM���36z˭�;�!ѕ4�_,�
[݌�!B�y�m�ˈ>7��<U���v%�e���5��Ϯ�����0��*���>x�q�HB���OQ�+�W�{�y=(B��R`�x��w`ÿY	73fp�L�)��.B�b�)n��?�(FaϽ"=��k�0�9��;󵺾����ӆ�a�w��@G�@f���F���X�G��TB1A�T�XuD:�!����6AP<���?�M�0��i�?�g\Qi�5@:8/��j�S�j��5fc�3	�N�'�!��\�nZ�����t�vP(.�[E	��OvӖ�=��ܑE�q��:��J�/� ��q���=��8��4	�4�r�9HM[��A%���z�M��9��2N8�̋�ڣ�]��9IH�m��=�H?ģ��ʃ�J���0���U�6�:��:�[Z1��Zyt�;>b���0b��2SK��� ��o$j��
	=d�C���j���tE�'��o��̶���������s���Ƀ�'�=��� ~���֥�\!�Ġ��k��/��A[=�&w���`����q��A�=x�L.��@�!|2-}v�P{hQ�+d��P����r���?��%�f���j�İP�l��F��?�}V�G�&s][���mb]��=]ۀz�������g��n3�8�Hk �^4��R���WLgD�d'IV]����$�8D܌B-�@����"����`t�'i�?��.)�g\'���q�
�/���j�:+t��l�O�4���*:���x����ۓ�"���k"ѻ*�&��/ɗG�E����s�2!\�F'��y:�1����Dd9d��q���f�z�b�;��!�ES�+�����U�[gP����Pjw� ��z��J7�)Ոj��z�
»O+Mjw�ݳ��.R�=Q�jYS:�)�\oM%2B���M*ϒM�I::����R]\���{m9��G��m:�8;�*���B���jOO
�[b�?X�[��pz@X�_F�{�s��&��4X'|��m�ڗ��y�qb*�9�,zd��V.#�
`f���F�Ϯ
6�c͚�gG��6�w�����Z\�BC��l�������=Z6N�v�L{a��e��A��.���j&�:��#+�:�����{T�~̬�&��,!p@-��j#��<z#��`mXŢY]U�0�ص�"ۮ�\PT�E'��
sm�ʪ��o�"1�!)sO��������5.]P�āW���n�?H���f���3���G�S�Ѣ�y����^�_ƱT��ձ��OR�2���;65��ŉ4&���{૑�<�_�<gQ[�r���o��\{�e���ګ�r��"k�22��	�P��k k�,�>{q�	h�֡RԴƳ��d�gʄ��L
��,��oPh���"I��KU�2�[1Ė��kvM�9�2'mՍ区ׄ9�$�h0��~�=�0'#�o�WxLqP��l�I��`�`�Y�Մ7ӭ�4��ħ��/w��0�Z����=���m�~��l� Eq��>���%�/�N�G#�LJ�g�y���S��C��K��=��$�.U�D\�'�[�/��H��=��)����"�	�>f�X���*����/��p|Lu���e�z��h�pF�HQ텣����/���&�5�<;��Y���2�b�m�U��7�˘5WA��a�{�迉m��`,��8�g���Ҿ���ss׎�Fg5U��� �}�H{����ۿ�F�W�Ħ|x�xf��qI�-eл�������+K\��T�g�v�R혎�.����]�%��/)��X�`���Y���V2ð�^�>SLۚ7�b��X�Q�*z�J|w�;5�p]S��U�|!5:<�|��=L_�\��s�/Cb�{�����E(\�&G�ȓQ7�L�����_& Q�㥖�"��M��Kr,.	�(�����t�k����m��L{5}����Y|�v��zZX�����`Z���m��$R��S޳��13JexX��3����I�{�A�{Sw����[h����\b\2%���E_�����|BR��&a�Ī�P�&��P~I���>��A>1��Yx�Қ�j�Qt���8W+�GTb����߯�F_�	��ч
�,6�~��J�2�+�
η�7��pE�E�o�l�7����D��#���Y'h-_H���W������n��>l��2/Z�ڣ��b�&N���t���!�HF ���u��ٍ�r:w6UQ�l-��̸Zs�w���;�a��cS����4�a���E#l�3�Z#1�Y%���z5Q�����Ie/M��{�9A<�;�ƣ\n�{�3����E�P�&�!\eK�Ќ�E�i�XB�R����_v�����o���������J��Mj�v�X�Ӫ�m)��\�+��O���	���~����h���y>m�v%b+4��6����N�X:�bw8���F}�oY:��u⚥U��R�W���£��c*t܍{�(a�*4�1(��K�QR�����`��M?B�[�r
עO�
1�CxB�E�Basc�CR���jD����uj��Q���6eͥ�^���WŽ�/r/�%�Q��<�]�{�`������G0�&�aL�G���bm�E�HY�F]�B�r7ʗ�4Î�S=�$o]F�h��?Ay�^���r.�!���Whp.�cHPE�)��9��O��+eK�g�7��?���1���.M��8Bi��P��;���C@��W"����J����J�<�ҥz]/�f��U�Bb�@,�O�|o�rA��h\m�JݛD|I�����X�M*id�?��H����J�ρ1+Y�&�J�{�� �P.˘J�����+:�m��ީR?��i�b!�,:�|�$+ٍq��r���Ub�؋�Ş��Y�Jr��8��\t��|�0��+�n9��+�.���C{Uc��p��C���C�o[����ނL�#��~���|O�����ב�J��Wלu�h�~g?�@����gYk�-�ҟO�0,��=�[�d$��ZG�ry`2a��K��nxN�~��d~u@����}����ħ(^M�n���y�D������/��Y�h�U�	�g�[q�� T4b��_'�Dk4��U����M}�a)d	�cྋ�����'eO+)�y�~.���z��RC�q��
O�� ,���<Bq ͡Qo�U���=��/��Cm���PL�dhǂo&���lC�����j	f�E�?�g�65p�#��[�	���P��N����J���[ �Zp��*��K��WzrT�é
�$�,M*5�\[�#�ס�r�'LR��'�F������ˠ���_Kj�Zm9_�t����Z��ׁ���@F����{����E��_
}�l�*�3���Jv����M�UX���d�O��F�J钅�
��%����c|��"� :�W�'ә~7�Vށ1qј�
��XZb�.m���d�v� Q�c_ZM޽�$��S� ����!��lOQ~_�i�^P����/o�;��;�%�A�d�qi�HD�-��x^	!�loI��.^�&u)fZ�h�w9z"�K�t��ꧨyI�0�n��UW��/�o7�rXc*z��q���=�cF߈$9��^λ���ҤBҩ=���e���<�fe���.ʥ4�)�x'TjD�6��7��+�ɴ��bI��l���>Tu�"�!f���&`ežh�nd"	~���B��:C&d�r�z�eF^�0J�%UF����##V�����0�҇�]�g�tK���j��;���z���Zf����Yٕ��JB4���*�{�Ȓ��~�I>c��e@jϿ�Ũ���W%��/Zo{��]Rn��`�����W9n�Oe2R2�Lgp�G4�&�H7����}���ɽ�I{����qV�q�?"�s|���oFl�ߧ�1i��{Ϛ��b�#M�R*����U�Rn����W�|� ,�2�Wg�4�=����(#B�w��:�	�����Z�lԦ��Wrbr��̪��ј;\)K�Y��M��q3b��=͢�8��-W4����w<H_��5(f��b<R�h�Gm��8P/�� 7�L��f�	ڞ�1�w�E�9f��%�����v��%�g��[a�@�y�ٲ3X!S���O/LjSO�焄���5�*@P�άie�is��Q��U���9 ��g	<3�k?z�Z�g�}E�>0�?Z���`�����TD�A5��S�#7�&���m�$�K�:�řS5I�������!i��U��.~��O���~��CO�,*����H�J�S��?��_�M1;#�Ф�MB�}��W�T��/i�|����e{\�p>1̇T�n&�)V��{(�@#�0g��W�m[�h٫�x[�S$.m�Ⱦ�-������[����Ӽ>��X�j���0��͚����>����K]J�3��f^��	;b����@*ζ�.6�1{G�\�v�������V霤��fXqX!�ii�ݍx$���؏�<�bߚp��PV����ʭ��{ar�Ekm�9���jEB����������{離���2t�P�l�����{J�
 �ůX���V9���np���`&�\d?�^�ͤ�{�#��a�ĂR��O,�׭���8��S�W����f��XOtA���ʏ�c�܋`]��F�N�����od��ތG�d��$7�M��i����h�x�+���|���m 䑝��,n
ڗF�Z�v�}�AN9��M�dPg";� ��}�e{��Í�BV����(TԌ��~��P��� ���&�-���t�Q�yx,]�Qz�ن��������r��)=���zB�p!�rՂP�wܮb㘘j���݄Fo�tb�+�X@p򓌎Q�lՄ�仚dd~�U�MA	�fϜ+沛l�"H�<g�ZW}o�l^#���E�}�zw�!d�� �5b�>�Z����jD�I���R�e�E�R���GqA4�nH�������V*]P���fV|�EfH������=8���[U��uRD�k�%]���m9˔���v�Ț�܄-���I�q�17�9���׎�5�'�T�R�?���C���[��#,jZ9��PhQ�;G^a�o����PH���B��0�zr�,9���}���ҩ������w�X*gr�����o��X�,)�����¡G}��g-/�TNk�,�@�M-.�����hN��;=3F���Ⱥ���}�����HtV|F�)i����M�ZKɐ�R���Vx�o@�#��{ƣDj�{��ْ��v$���<}	K���F+���,�{���~�g[��z��)�/g��AJ4��oUZ2�o[U���#��.K�S{y�c)��W�v����G�A�l$?'$��e:ն��O��<����Fua��L`Syg�qU�щ�TF��i����>paf^��l3l�
V喘`��(O�2��տK������:�A��+��5\�v�n4�&�a]!V)k�Pt�`8%xߧ|y[�Mx�\E+�(X��}�I��2�@,�@SM(\5�N�`%��A����7G.z"/�y�CT��\�$jfU�FQ�,�Tq�)ҳ�f�X'��3N���sA�Õ�$,0l�kƝ�[O���֯�37,9��R�YX�-eułD����u0T����.^�꾅�i��+"�u�#3���d�P����*�[��$fۙDӠ0l�)y{����Z�x߷#�i꘭�?X6ߖ��5�Ac缄�w����>�ç2
��1 c��-��^OA`]p'o��XC1��[%��z���T.E#�J��������8�Q�&Ĭ�`��؆��P+�8��z���\=�)Q�D��ְ��_�[R�WȤ��8v\�Q�K���fv�A qIu�������cs�G�����`����l�F�����T:�����N������I��m�n�#�PKJ��w�s��o��gK�xb��q��CQ��P`94���4�Z��&��n��aMSZ��g�$%�8�-@9]�4S*@��',"z�7D�uc�{&،a7p\j �x�*nK��)k)_���J�kpmxI�q|�ׁ�@���,�Km�(�q�g�BS��\6I�|Ij�!y� �w���A
�$2P�~�E�J�����|)�d�Rp�_��)v�k��@�z]�Dg���n$ģ�ak�$�t��0�{�$cb�Ɵ�