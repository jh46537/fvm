��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��_)��%%�.��D�ֹʮ��������7@��=�y���fA,AQ�GD'"��j���<x�H�I���9�|�� (�!�h�"�e#�~iN�}�ѕx�����6�5���֜�J!�)�+�af֑n�۫DFJ�L�,4l����.��Y5��s����7��U%�o�	���g���#�����ߗwR�TR��I�vxXD&�I�r?�9Z�c�
j[��@k�5��PL ����+�Y������^WhuyIz��Р�?�%T�ƽ�T�Pn@av���Gow]M>\+�����}(%��V���e"Y`e�.�B�Y+`-�Gِt$
�12$D��w����M��j]��1�'�n|Յpǆ��l���]���?=W���4L�
�����w>�e���r[�|��1
m�}6N��!��\O��$�>ߖˣ�;���
E3���)=N�˜Z�ܤ6&��XP4RD"'�~`]lo6���@i��	��4��}Þ%f�Ǳ &��D��w��V�����HT3�ۥϊ�?�9���%��G�]�&��ޙJ�*��2��z���I����� pDv�֬�!Y]e�ť�R)I�T�,�x�)="�!����u\����eX��`-�Gl.أ�	;��|��u��iV�`�Gv�{c�\B1)��r��y̇mtb��5[e.�}+\�q��D4�f8� ��A����h�e��h�̪�Xe1rCr}�B�bl5f��>�A.���o~,&n�^�9%��� E&��|x�!LTҽ��-�b:z�n�,�u�*go����±���U��?���5�=��鬔>��c(z���-k݅�O�N�c;�s0�}@���㆞�^��	��QPk1O��B�&e\����(D��۶*�K��­��@(�k2f�
��a�X�7)c��g�i��Ui?�D�ɪk{
GB��O��^nHD�m O���5geE! e�X.˾$B���|�͸��J|$��mz�.�J:2�U�Rcͯ2�]K������[dDw}�eQE�M,������/�]�w�%&2.m��i[#d�^�X"9X>�V��;zmf�".k*uy*�u�D�Ͽp��
>O����	��+�q���������������� u���O&B��]Dp�a4�]Ē�0���� �!�lz�ZRT~�.�}9	�A8���)k{K�4��*O\�,�����6�Q�쫼,I�A=C�VM�+j��%����A��U�AC �y�/Y�ͩY	E�=��M.��r�@D�-�a�Q�-�l�M���P��a4/���Dkw�����Pٷ׆��A�fPD�������g�?2~A
ȿ��C�ܝ���O��
s7ތVRGF!Kv�^7=���)�$��z
(5b���>88?�u�ȩ}0�ǅ��,�H`�b'LlN�.�F��:�/��[KJI��i� �ԅ�s@J�n������� _�z��!��&@擤<eƵ�VZ����7)xE9̓�؊D����❴�����^�sY�C���O5X-Fv���N��kV��Uሶ7:�@�y�I`C.�|#�����k�lyz:���q-d���|ʫ����*�2�[���v�z�ڴ\�XSE��M�m��}U�G�N�b��ml�v��=@R���&�T")��"�g�S�m�'/�ϔ�! ��	+�T�oL>�X�tO�[��+A�c�Oh������d�ux��[sWpaNR�(Ql����u2��Q��Vk�ڂ�\
�dق�<�ěh �!���33�Hcn9Ձ�F0�n�9���9Dmj��ʋ��qw ����3����.tt��%����.���ߴʷ�,@�72�$�y�[l�/7��E��{~�+}�"���9���%��K�ު�û�.�YŊ� �%�Q1	�֤��B��>Nм�쥥J���1��0�+އ��Y�d���X�V1��$�	��Liy �C���;�>�hgF�"��<L��9{�=�%ٿ�"��	��V4�K*3�~]����i�n��Y��9�����Nș7gmEL���%��(\ ���G��<�,��$i@I�vg�ikRp�n�l���V���ad���%�HE�US������ ��)*�����$5�#��O��B�%�@��;�47���];���(����{�)�%�U�/�b�;;o��]��YS�x�������u�<�t[
*���bQ+o�ID�=}Ѐ��4���er�o�����q�a_O�
1����QZ�ܻ�HJ�g��)�JM��=�V��̓\r�;��7��p��!f�������,?�f9�MT�Z�)�|�Ou���9O�>4���W^f��o��s���[�~�?��Σ\����}�խ!��n�<Z"�����)S��s�i���`=��v9N�zTG�j[R�8=`�����E�ڐ��J�OH�vź�=��<~X��c��$�\�e�Pt�_UZ�I@P�Mz�{Zt�;��8�'L������A�v6�d�V�`�[���چ��1�b���Ff����FMȊ�|n*�R��I�R���x�Nl�Mk7�(�9��6!t���X�D)�.Jz� �s�.L��u����&�z:��U.�вA���9�|�6����G�f.E��3���]� p|��ȡ=�/f<9�|>u@� �T#�gQ��]�3�1��.�v|c ����v�����?��	�d�2s�I}�G�E{gQ�4�w>5i~��sGRu���h������@�m��}��
�����<?��W���f������]MV}����(���h�DN\�\�I)��,)��B2������]�L"c���i�HJ�}������x�-8��a~G ����$*v���Y�,��R�`_��xvv�M%[���)����X��̰oв�IU���=���;ؽ����]���?a��4�_��4P�����!ث	��m%�x���!g���Y���qؤ�y�ou)�mj��L\٦�׹���QK9!AJe�����K��/覢W�vT`pA%w�Dɫ��|��̸����!&��4��/�$6Z��8~�����?ICOJ�����	V?�Z�}3/<#��Ymy���6{V9�/ �]��PSkMg+�l5*S�����覒�מN�ڰD�1>�N}�D$ �̈�E9Z�?���3۱9r��j��?=@�1��2��C�*y�b�5����>+P��u�+�e/�y��V�{j;AI�6�|G��p�V�|2'�ǝ��G-�2K��9b�*J�N{�kk���f)�p�)T$�/�p�eq��OW\,VW&*�EL��!�zӥ))�K�����TFh�y���BI��h�c��uȌ�Cw`kY�E��P�ǖ;��E�W+k�Qj����,'�M�L����T�F?K�@��G.��H�Q��t1��������wE�a8շ|�zUF��K���^0��;_U:���E�o
n��PJ�[��u)�
�! '��[�şX�h���k���A%�/	�`Y��}�|�įD�^��}�7��؃N���i�+���gXU :BoF8b�4�>������2n|w������0�BmC�����}�Al	p+T��r��}����Y{����Am������'�Y����	(�ǰa��9��,��>���
���ҕ���*j�� tpxN@L{.5�/zq�mI���+$5ox�04�-�UScSc�~)
o�"�4�8��R�oꊝݐI� .~8M{Z�Yj}!�ϰ[�^��S����N����#����T��	aǪ��y�����-{�Ż�9�پJ}+~�{�9�%�� �.���7�\�͹�p1�z�V�<��i��JwM�x ]�ԧ�)11u�˞�����#F/ �����M�*G>T���ҍ�\nvw�aϥ �0�� >IK�n1$�3"��"�����;��k������Y=
kJtqu�5��̦�z�Y3��"�&�z��}���J	4�VK���h5���q��Kp�REo�#�H�/6���q�lO�sV�Yo<��/���n�S�~�щ[�´ԅ�#W���_M��C� �j��K$Z�1Yo��	���G�ؿF�&~���L*rOB�f0�u��h�6���
0�mE=C���EQv&ܲ=�~ x���!��?��s���,P� N��f�X���2�UV�=��}Q�rQij��\{�N/ԥ��rw��ͶF�6�(�K�ڷ�'�y�u�{c�H�
*I�H��;~Ȉ|:�D[���;���|�������jbSAyŔH��t'�s�I��C����zMQ[����N��ͱ���d����(
�$��#y������N�jm���i�%���N6Bv�Ͽ�Zl���i��g�)�����}%��֫_�i��;n��~�Q�ĺEY�������l���O4��u(6r�j��k=�rY�B	����d��=���?�x�l���/�ڈ������Xɼ��j�P��~�c-P�wa�Hq��8�D�W>"��|��A�U�+<����e���v(�X�|�~3O���A6k����M.LJy�����ډg�m6ۍ��"U�8��zo���S˪��x|����b�#���w���f}��39�wȃA�M�#j]^a��A�NN�$�����A�fA�5@����9h��,�-kr�Y*
�=%�t��gC�<�vݽp޼Ṽ6ހC��*ܓ<�[4w���m���Q�AkMi/�C-tx��nb��fM�T NQ�`ɒ���I��:��v2�j���2�<��Z����gGyЋ[]��̓k��HT�!_�%��m8i<�������hة�WHw�
>���g�x���^*�\]�G�]8?�O)�h9���F���idVV.���E���?��Zc�/s�N�r��JE�uǁb�*�ܦ��%!e{qU���9X5zA8��}$��F�����kɊ�&!�j�b�s{.O�~r���Sd@d�/L��pyryH�'������ai@!��G�fW)X����_DW�����U��N�,�B�)�y�g�/hP\){�1oi�t0��q��!	^7P$����ש,]C�Ǽ�����jH8d �P3�ZQ�-��Ȫ��5��la����,���'�\/k�]T�'@%S� f�_?]r��urb�M�U��l]�n�����'�_>)�������Z��C�!��~���p�D�8���y���ĕ#F�:����Ia~[t���Q�+k�.��v��>  �bZH�e�|<�nSe���J�_cMX��kg��B���>t��ʉ �b>>�mf�|�΄��D{�nT��A��6��������hs�,�}R��W-6+Ih�ߔsJ�{1/<��Y�as�(n�/�i̬�����ް�K�i���ј��<W�&~iQ:��1Yk�nm�xաi�`��9#������lx�2��7��1h�
�<�Xy���H��/����/�غB{#|Ј�N��N�c�l�+�5�A�t�@B���� {�r�7�;D}d�l:p��S�:nN�j$���ΰ��24�w<��"Odc�!=:�e~��� D�CGx
�=�;�D�F�9H�ґ	,*�Em�m��C����A҅k�3r��ԅvs=h
��u�7�*57�/u�'f+u�]��#��xIhǥ��c�RgQ�r����7	����?֧2wu�_���j%���U)�t0ò�[�����xv}HOL���9���>�@V2��dy/)ܮ���. �v ��t�Í�l�"�Η<��Z�O �W�(�Z�I 8��f���[��ٹҊ3�v=~ͬ�e�K��K���.?o����&������S�{���"�DfO[����­��j�>�	�4~�.=0;�K0Be�Ј��y%ʉd��uvpޝ�dÞkPZ���,#�	m�]��bA���57��;'�0)�����O~Y��=>�=P?\e.�\|��AӾ���ͬ.��
�mj�-�=�	17�����#��[?�*�L�b6β��m�L��@��]���� '!ya�����,k��O����!�k��G�6n,CJuT�@kG3c(�?���h��s6K*@�c3�4�N�Q���t�t��m+}0�xh�=�aJ�U�<�D��7C���Ƣ����~c{���}a�5���S��4�)� ��\�Kj�z��G�enBbl�H�d {�]�)�������_���6�"��|Ln{��pj�Q90��e\@�3�kR�b[�ٖЛ�R�� �3��h
�����ƥh*%�=�+�س��n�ݓD������H��~!�Ϋ�I9�*>;n}�j0ԋ��~�0r�K@�8m^Ƨ�����51��D�#_6�Y~��k(�jß����zx~���o�+^�+��=aT��m��5)� S��oP���s��[�jk���7��)�f���H���n�ڇ�+V��iED����-Ёj��U�-Y5�NCG�\8 ¨�"��6�ɬ���Z�찗 �u��iG"��0)�ne۹��ւ��F���S�аF��d�u)ZYn8��;`O_۾-�G��V�{��jVq�B���_��Y_�Ǚc��� k^ݬ��]���@C��yd'Eҁ����ǫ5�P���6�J)g�x�����Ďn��g��g�7�X�V�o��|:ML���Ztf�� �l`�)��-`��i���6vb��R�gXk[�D
.-@�x/�ͨ=�_�Uт�E�gn&v�#-��Ӳ8�lR&R��j\^�h�)E�/���K�QE��fT�`�JS�?������������MR=VxH�E�۷�&J '��H����+�R�j��s�=��YzUT6֚66��E���i�}��6�Y . �g�@�.�Q�H\e�
�� Tb�.(��=�Nt����'/[���H˃º���]���R���qV3� %����l"[:P��~�-��u��6����!]Gơ��=�h�MZ���]PT�W{�f���I���=�\�����Ҵ���5���Yѕ�$�P}�����!��}@����Pp.T�v�^�B�ؖ�ˇ�x�@ʊ$�4
fك�4U��.��G�X�C�+{U�֜W.`�C҇<��[��Ɖ���N �D N^L�m��l��ǯ	��jA�є��+�Ȕ|��O��7���@�bvC�KFz�����*���'@'�uְDc�?�A��GWW�!;�"�C5��d!R ��d���� HE^�h��]g��N߻�}��'��8+T�' HW�֋o������.�����d��S�u��C�tCXo��uIo`z�TZ:~�$�������7 Jq�̜��ȴ>��Z���//����m�\��ܞ�0M����)X��7<0�o{�I0�6��M�*�6g/#�	n��O�xs&e&*�X��.8	��%��8�RR�n��#�S%��C��;(Yܳ����_o��(5Z��y�EY!�`���=��,�8�Gi6g��&��iIBW y��NS7!$<l�]iF=�S��n�k��C�����4��b��
U��;AJA���!ƈ��Ř���U������kN��C�+S�N��y�V	<(y�W��g+v%B��Лb�**k�riIp�����C#Q��YO�h]2�Nw|]?�`j�X,z	�9��3�O"�n��ff���_�o��9�а����w����>��4�I�+�H�0w��"��h~���$��oo	���vHLbQ�^s�} mcʓz�$^�Aң��Lձ�N(�.�&�j�Ύ���� b=˫ N��m������E��q�l�6Hm/� ,4��$�ox�·�7�i�|�4��������7��S�ab8���-ow^T�j5�ʆ8���wȘ{�7�^�2���T����/͐"�p�뤣�j7�R �v}�LUiz҆Y�E���6�f�AG�?��` h���<�Nw�`U8uy��f���$�]�����4�ż��ݎN^�?��0H�d �&�!4�֮��K^̌n$��]ǤP�']u��c��rh�+��ŗG��!5{=b��s����~����A�K�Ѐ��,q˯��!wՐc�����������K��C�n|G��TZ��y�nG����W���j{�<����WjK�{�7��tE��ug*�Ћ8��I���P%���!���҈AC��%Z0�9B�{��쓦��G�*V��p�c:��4�*�'O���(߱[7��4<$/N���5,��|/�A[��X��hInDI�u��B�X`�o}�,�-�h`��ĿvX\�4�o��e\X��i���901IpTN�S��� Z����7\�_)����x����<�{賥m{�4zK�	_�b;���x�qfc%���M�n��R�O�L��.�8k��� ��sq>i �s6�8R��k��}�V�\y���P��N�$Wp��~���Y	����G��׬-����0���hP'��BkT<ZM���Q�&�P�N+ ����>�Sk#�^���}�X޺�t�6�q;VRn�6nT I*��7@��Y�P���h��ƛ���_�>��+�Gd�¦]�C�����"���c=�R������T��M4��@P|��gR�ި�2e�({�L�"0F1�ݼ�M/�Ȕ����e:�x��&��[�8n&�`Z�,�"�X�������	��-�5�ic��IQ�7��leFp�킃N���E2t��믝���Nq��&��J��kj>�*���7돮���&>�z����nvx�1������C9�m���M1>&�K7s5�&R��{k����ӭ�*(׽S�E��0M�.�_�w������/�O��o��cj�`��]u�����0�$z���1��7V��Q��n�9��uۮb#&���Q����Tn>�&K�*i/P�5�3=.Mf�R�Z߿����������Md�+0��U).�4eZ}y��t%��͚���{sH�v�bd�x4,`�q�9UC4getq�����lND�������\�n�4�?<{;r3d$9���8<?��Vi� e|M0��[�������{6a�!CX�w3�2V�``�X���2�h5Ѕ��#���_'ChW�6����G*� 3d�,�*)�s��-%d����� ����O�M�jը��.�5_���Wu�+(���5}��'SY_�aW٘'caT�χC��T,f#`0fw�A)�B�����P ��g��+�M� L"��h0����L}[�K$,�q��Ŷ�qmJ��9̴�3�.�����
�S���(����d)I�,~eQ*�J�b,�����a_�Qd�~�3k;ݨ��A��w"
��J�+?>�3���#'�&7&���޳���N��i�3L+݀1�7�F�������~�x�v�E�!��<�J���j�{��TJI�U�l� ]�7�e
��{>!ʩ����R�ְ9ʂ��T,�.��B�\���0��q��R�aL@�.Հ�y6[ �~iI���+�/��HF��8hˌ��	`I�����s����y�-~U�F��� N�� *W��,>�
��/>���B�� .����G ������Bzq߆��3�"gm�9"�eC��ػ�j
���S����/���\�e8ƒ����_=9n�m�0�n���3��8�wK�GT�o�'��ak�Ɉ��3ˣ�rR)�V��i��Ƕ����FO�@���M�K�@]�R�_��Z�Og'���P.��r��|%>����1�a�=�]�����S� S�d�JO��H�8�����y����o�ց���*!��R	�\\�Y��<v��]�lU1���jX9�Z�s!)Y_��m:�v�ҥŴ�6�q&��*Q�'	��Z�ˍ!aN�����C*�6Ra��;�z>��~S횘QB���f��7 g�,{�t�o]�øE�c���o|��W{mr�B����q_i��7����o*�q/�Ī��"��Z�P�Tr�s�G/��4��D�W:��gE����ז�KѸ����~�5���B:Y 4n`��:1lB\�
5b)k���!�Ο�9�2)�j�����;�Z4�ˎ�-m�v��럯�E�		��DrHnge��t��ӂp$��
$�"d@���������@̬�LR)�i������_��dµ�|�M�g��+�6=�8�w!��Pa<��>�DX	 /�/��Ht^����������O�ʎqxa��{���!X�i�����/ f���u�'��Mr_J�n��ծM#D�0�ga�����fgA�N	 �İ�{���l�A	do�q��is�ω�UC.�Z96Vʋ��n�(�L`F�m���I(<�!�t�dL�n�u�������c�%V%1��ۺ0LP��ǋ�wD%پ�F����hS�Ey��o%�Eo�!7�nA�� �_^-�|���LМ��x��,�$�Dj�c8��/�j�!��כX��m�p �O�m+;zhSu��鮥G�9J�?�ǌs ��B3��;�@RaE�gFm�j�7(GNO�Rn��k7�S:��{m��\����JgwX�s3
�&������0����YL�kOE� ����:�,zN������֙��K:пa��A]�OLP�uXx���㋌I��#6@�1�m�����z�wld�w��A���Z�rRm���?�T,�a�\��3ǚ�ߤ }_�L�Xf��D�!�;�.��N��<0d�%���ƈ|p��s@��d�Uh=3o�>�����rv=�vx��t�-� ��&b�^�is�=9�#F���s<A��g��}1��l��0>�t�r�l�L�sp"�4�g@�?������A�սXd���S�(��e ���2�~p'h���MR{s�ֆM�l�49�9�M�)���O�^��a@7�탡��
J�{J��o�R��*ѱ��|�7���A��3��|�ƥ���L[	g������̏�b���;���$���4B��ymw �
�ߘ6���0���ǾL�[zz�����/�dw���&~9�r�('����`T��h3H����Z�!��q��*O��[$��rUUw�"�T�*�ѧ���E$��P������23��@E�x������f��h�S��a��p?�脨d���Q���|��Һ��YgT�젝���K��������Ƕ���(������" ����W�o�E[�$�YU��>�X!x�@7ܱ�|��F�;Vm�nPk�E�PKνL#����y����Ѿ��\�����(��M+Ni>xȒ�y�����%Sj��vE+oP��a�X�:y��3}.C� ,�9�W��Ǚ�-�g��3-޼�I�H���
YH>��k��%;?�rؙ��h���X4x�#>]a�r1ja�����VR�Z����� )��&�2&/��N�u��]>��G*����X��������?�+{�t1���_V���O������S�H�r�<�~��&�e:�2~W
b�HP
ٵdd�B��}?�dפ�R�Q���.���f��Z����"&���2����N��R��%���k0X4Y�ޞ:P
P�ei�_�1��}���	���Eb#�L���4F��� [~�f������94J��(	40/ǆ"��mH���`sځ����M0
B݂unR;�ĊE�U��#�n _}��~�����p/m �����Ri+Hy��^�b����d�W��"����d���o}:��7w�{���7�y�5]�-gР�8��n�Ի@�P���)	�W�h�Qs��7���P����^�ۄ��P�aWu��|�ȷ�F��jsD	{z$�'0�G�)�9����	 �)��@�/�E�.0X�x��/eI\��Q3�vJ�m��7|��m�y�Z�a�_
����#<tIgT���&��Ң2[�������Kmw�;D���k�%�mt������%C<�Q`l��3�F���{���nV��T��(���W���j��c���|��x�G��d�yFl�ۚ�+��ۨ݊�r�1*tdM��b�x�z��Qj8C��� �h�e��0���fm���umȵ��5B����6g�o����|{A��FW��.mN�^�d��JC[���1�g����`\yfß��d��6�Ś#<��K-���~�.�쮙E���x���3=C���VŃ���$h�Z�F���$x�xb%t��'�KT���1s�Eb?��<XG��[��<&}�f�o\<󙚇���ءڞ�����En.�ℛ$�dkrOA�a?��h�D>�TN�S��4�w[�)�l�MwmOe�mf�H8x{�2Ƶ��[���KM�N(Էvk\T��V����׎g4�L�� ��Q�>����uU�r�*���R��]V=![�G�/��o&�I���@��G�Ɲ��>�	 �uE��W��!s��t_�
�J
�lX�b�Z�A:K[�:�R�7$�_�������+�l��	���.ﾭm4��w�T�N�v�^�U�"�x�8����0"�ֻ07!��0V���%�KN���$t��M
5�.�*�$&�c��DJ��Z=�� a��ɳ('�^��s�qv{�$�f�*$��EU�b�>~�4���FPy��أb�]A�y���g���X�gx��1%?6]��O!�ݳ����j ��\"N����M��a5h��/=�}�Od�fg�Z��:�gY��_B%����!7�MxF�M��	̕N`B��$Ɋ2E��yG��0��*k�3Cs��h���
B�����Zi�'M�غ�8hfXXi9��|�h��L�[f;m-�'hi����"�^l � +�}5�b�G\�|�S!J#��H����\7����~u@�1��·@��/�^D����s�'�7*֤=(�x�{�NH��6��W��uZH�̀����tF 8E�yP{�W q��t�9a��.'����}����v�h#Kz��`M��x>�[�L�����R��욬S)A2?RF�@��ĩ�Z�m5j�V��W���'8��ޱ�#-d+�b��4٤@*�xk�>��]��Ŷ�gQ)"��Ss��țj
���gj�(I��J��2�����޳��3'cc�nϻ�jG��W >�B
3�5�I�zdS��V�5���.N���.�r��p��g[[=e��޽�`�g�s?������ذ�A�ro͸����C�1��������x1�ʯ����	c���_EIp@%�(��\�@�f�]���I<�.�M��+�==f�0����Fm8&����]9Q~��5�TC��Ԟ�1���+x�'�Wȴ�$���u������r,E��J���us�}7u$�Q�S�,���#����,þW7�-sⰿ��	��*�V����'���Sg�9�pK>�j��S�Wn�޸,;o�r���aS��HSma'�r�8�b���X�5�(� ��-1߾{~��XL�'�$�)��|�5�u0	�U�]�������[�T��,��f��ɫ��,I�ؖ4�Gn'��g��Q<�>L��D�xZ������q?����2�v|oK��>K&�1R�q�� �m=?/>;ck�Q�n�aN��'�h�	�V���d� |U��l�3#�U'0 '�-��56��H��i�%.@�ɪ/�S	�M�$U@�� ����M�y�Ռ��a祄�J:�Q�Q&A�4]�Na�{uZ�u?q+�6�eA��!��=��9�r����Q�� v0�-�8���B `��<�$�Q��{^.6��������A�k�ބ�2CDt�T~��LX#��Vߊ�u"��\SAj��}���,ݴ�cRĵtgux�G�F�{��-�x�P<����?�Cܓ��ʨq��n��V�h�Ж2�H5\#k��q��|\�j�u0��E�����Lmuq��)�Z	)`���]�-�Y��/t7ִ���w#t�<�M�R}�/G��:ev�)O���ޏ9���E�0��[Wu�Kf�ݜ^��h�H���vj�$X3����؛h{7��� �QpK�Z�@3xT�$
����Q�Ȯ�څl�~������҂6_ z���J'񤌛v��^0�moR�	��P�O"�u�꓎��wLO��P͸ �^���0�J4�#�S��T��ܦdG��d'A����0Z�	,�e��C�a�������m�F��*����1RR��a��<�;���߯�s��8�{@���
���[�����U>샔+�'�G�+x���N�K�B��0�2�9�.�B��ق���11�~����ی`\AԳ3�\Ly?�޾C X�^a�j�w��TqE|�E�'�U�䝑k�8�����lg"�Ve�RcR�c13��Z���
�>�4��%�Z�u�o�l	Dˉ�+���@��6X�d�>�50|mq׉�ƙx����B��)m�Duߊ��v��������"7�^���������G��Ƈ�SqOW�>���وq�քn&�c�+
�U 4O6HR��������=
�;]���|�_O�1�Ļ���m�b�����C(��,VB���Z�O#"�,�#��^TYH�{b nTT ���邃��v��Q�LlDx":SdR�/n	%�5nx��%����ǉP�[�v�J$�x�A�gXGwK��P�@����<���������!UF?��2�kk/.���@}��択�ͮ,�̑��'g�+��0�uЬ�|Sb�8�;�)<��h��2c;s}�2h��ç2b�������N�^��y@!I�#�K��P@��
k��F�73�uM�q>j�>W���0��1�y���y'�t��\h'��c��[��2F~�l5�J�V,����b�7̿澳d����m�uݶ�h��[�/��{\1]Ъ�)�O�����!G9�Q�Y)���(�����G6��Fa��;��Yi���*G����Y��_@�&7s��)�{n��O,�����k�z��s���+t��],�v=�H��^��$6��zU� ��Cw�[�?DY�����~��s`�Vd��X�ip�&ۛ���+^�u�6*1�ߟ��}4٦�-�N��w�\�h��@F��e�]`_�E����8	z��09[l^�^�������叓�&t ����o�e�NkF�b9~P�j	:xi����(��� '��Y�?�������H�����8y�v��fW���`��=*m}�OO�N*1;�� O,��(��<:�
��-�:m,+��^Z�2y5'!�Ո�]�����&Ժ�#N��9��]�����NE�fI-�ȟ���f�xP~e�8=$�x�yW���@?d�x�߹/��[[s$��?��^��`P%�_ܮԲ��ۄ2�Ȣ'�
����~��V/�/밾.�î�����6<x���`����%��*;&6f���_@��3��r� 0E�߀�a8E���r���MԼ���ݎ	H�`��fr�S�Q�"܈�Ғ����'}(uI�t#]��.�IWY[���X{�I��2x~���0Mb�m�n+����Ş�(���`���K���9�e�Se}�"R��k��6i ����_���=��x<�8R��4����De������^�������c^�Ð5�(!�	@W@�x9ݯ1kq��Ć�Ҥ��^%}۱�Б�]NgU!�H�@ԉ�?��`�A�Wb؏�M�W�+{b���u��S�[�(�ꍶ�]��>~&�{�;&$��1$�;mFx3A�x͈�4W���r�il'�Ge�
�{��R�yl��W��%%	��Xr�3:ə��]��M`�I��z�ʼ/~�l���8�)n3Ě��9�_��E��2�9tuVеЉ�B�ȆO�&8[��D�7�j	Κ���!�W�g�x��*镙`��GH*x�KEE"Vn�b�l��5�t-N)�#[�&-�8����|�� �\=�1'�7�q�sc7��BDߢ���fR0,��R擑YN�}���L�^mf�u �j�1%��(�D�],�+��i�A����t�^�!2�b5Ku����rU�����Gz�b��޹۲#��+��^�7/"P_�v���
I6�X�C$\Fqg6-�|��O�G�Y���X:��k5s��TX�Fh���Q�\�2��&���@���b��_��p}�+`�,2���@�i�������Kgٴ["�	}��,R)�Q�7�������i{�i�2x��R��n�E���x@��s�h��	��]���TL�e7Nʅ?�ͦP�,�X^�@�,��ʚm��t'�"��T����~p^ ��sGvl�4����9�N8� ���>*�	��r���a3� R���*���2[��E�#���Hǟ�H�SM��k�z�N㦱�}yF*�#m�R���\��L� �<�$��.�<o\T}�N�fW�D�t�֓&������{�
�X|���I��^�T������&��_ �l���W����3~�)!&�Y1A,�;^��};�� :���B��{7s���LɨW��Q�I�RT��ThX�vUVnVEq�p�A�?�@�-$�Z�J�XՒ@��G���Nm6\
2��sI�A�,8�ځ�~��n��P,�cݰ�jR�pB�YT,���HN�N4�S�����;5�N�H�{�g��v�\������L���]�4��B�4�#���	\���NKf�;F X�@�N;�4ē�<�d}wv~���d���?e�D�)^����#�TE��'e���N�F&+�>��č/��f���J��B#��(8�.�H�C�N��]�r�O���� !R��y��"g�P���=�ϳ���"�%��6$L&}���[��[�e{��ʘ��;��M�!a�*+t�̒ޟH�@�g�d�;-r�P� �9q��G~���8Ea�e�Z�#�m%�w9b�M��b�'���r���c� ����xWR[�m?t�u���{�v�A�O�}��M����ە)H���.��Ys�\J�J�2�G��LF~�������+�-nR腏9��9���^i�L��AmQiaaMg�b%�o����<�f����$�{,����/Ar���y�J�@S��)���q+N\�t�rp�����$��k�9���� ��=:d���+�G�I�N߂t��
>�C�N o*YQ ;+|1;؅z����V�'p���G~�k��E+�;l��|�XXŀJ7��Dfʢ�q��Y��g�C�<�"gA�uc���-8L��E�-�=HƗP�A�M!1��*7���������<�x��W�<k���ɫ��>$�����\��7Ŧ딍к�� �Eq0q���i���Ƭ a��J^�@u�����"T�
o��s�p�.̐8��prC�M��G�l;�3=u�\�iRpQ�G�#� �r��k��X�jW|�^_����
1u;/�	N�Ձ���p[���1to_���R��%�<�%� �LD�Vc����H�'� �9f�ٍ}��(�SR�������<  �&�^q�L_��/��r�q��$����u`9s�J"
!M�Q���s��"n��g?g�O�큦�ī��R�BpO���h�������Z.HS7�d*�;<C� �K��P��Ċ�P�u���s�;j��fw .0�(�?�Z�Szɔ�\W!�~��#]��H������ �w�����ÃX��m��D�M��Pܽ	�� "�_�L��"�tz��y�UP��9I/�^x�U���x襒l��H��Lؙ)�0�t�D��(b�m����cf�6�?��8<���u����@���/�(@�*�e����9TGYm��Z�1W��� K_z��?*����|��}#g�8��Ϧ�����P�)t�Cc�;u[���'Ḛj��-<�7(�ʢr%������g���>u��B� �7���� Z�툐)8�"���"��;x����W�GK�5��Ou>��9RF�\x]��SF5���h���d�]�$�z�C$�s��;0ggv��w�o<�*_l�ܒ�#��į����%��؊�$G{M��}��]�5_�I�ˣi�{S�j%��A�*�2�|hE2���h� �1Y��Ly�O���w5eP��'D��/a8�j����eW�m.m��w3���� t��f�������_�66K�Ǭj;�s@3L�����vr����Wl�A~cQ�����+�x39ؕ���6�[�35cV1��@`9��t%���#������H��U ;򽧟�-�{�9�'L����5Ϙ^%���%�m٥��&��$�՗�R��B�&��;��Gbݛ�<"U�"��4];q~�ښ�M��lY�K�b��\-���%�֪�ό�W�Kp31 Ƅ���/Ui#����JS��b�]����C���o��<z��d�`�3��V+j�`����ma�lm{���@�'t�ݷFL6��D�8�v5��:��QY�Aؔ7~����T�ꉗ�S{�q!�cF+u�fC����s�_
��ĥ��P�p1�`�!=�����3@���e��G�'Ii�U!Y��H�-����l��P�M��$D�����_WbiӨg%K�Lw!�ټ`�9�イʖ2P� 3�c]_�W )�Q��Pöm�-�Fa�$O�
tS�$�!�-��P9{�<=I����f�_1�B�Xۺ<�4EcP�����i���д�z'���Z���%��ˇ��σP5Hn�� ��aAL��<�k��t��qO=� z¢�M�̟�'�|��o@^��P� �#� ���n��]��۩����+;�P�<�{D@���`b��*��= Ȓ�¿TB֓��������)�D�1�U�S��p:�o�qD�)�%N������-d<�=��=�L�4 p��b"�V�|X�����i��brN�0U�6����[�*�'����r?�u���Tx �'zg}��0�K
9�w��Uh�m�8��k�\N��15��м*J�eki���&{%�������/>�����k���xR�|e���;��X��hzM}H�</�	��Xų.�JΙ����ę���b7/�7Sc�K:c�%�e����,�ӍnӃu<J��a��y����|a`�SC�	;7��l��دg�8�-q^J�%����hHݝ��,��(�`�hJ8T�M�-�6R�}��{����jS�cw��������QEg�8���C���D 	�+V�B,�����n\⃭�ras�%�]�ֿk�rpq�p�f�;Z_=!&���S
�NA��� ���;3ѥ�뒣B��/� ~F��u�����9���}QҾ���$�{�!�ֈ: Qs�����I���ś�Z�ϻ/WIG��������_�e�g��Cdhxjk�E<O�5k%�c��AF�`$���ǆG��_�S��aX��Ux�ޣ�	��z�d�\(�t����k���ٟ)����lǻc�[x!��(!�s�tt���$~�t=;�y�EW_�ケ�9K]�8�ͧ��f�`�ߠA�B/TR/�n��lv�}�]/#�s�j�<WԚ1��^�8���ö�!�5}u��M�}/�����l�<S���<˒2��ו�%��s�J��:z��ę(��J0sW��<8���~+�t��W�*�7�k�8K���@���z��	����#S(J��{�ֱ8}�}�	=�M4m� �\�z�-*�{Kӡ�h��s� ��̃�w{�,$���&mv��-����x�h�3?��L������V].�j��'x�!�b�-w�i[D�b3D�]�wZT��J}��h��fIȿƗ��RަA(�i�k$��MRV���.�%��ę�IE,�������	�]b̡�Q���'85���3�~洹O�:M쨋��0�b(	��Nl����]^��mY#XQ	/�*mqE��w Q���7�k޴R]
�(=�8rq��7��~xikB��{���#&9�͊z�\��L�]�u��,+��D�J�l|���"Y�vJty�EQC�g�k�S^���A�Z��	=y��W&t��yHu�j�@G(����o��0�+~��]��{���_*�~��~���Ƚ�S	nm�&��ݿ}'Z�C`�J�;֏㎻
�t�S��;�ZO�/x�>�p*�p�QQ�ir�!(g��A�S�����	��0y�d5�dD �!Q�!�a���U��l��Ԧ���vd���O|����Cڎ㹪� v�~����1B�o� ��2X�̡��֎Q����5kH�D�L���*~�BX3��V���[,��iı%,�,��:y�Qbjh��OϚ)F�? ����hmf�ˠ��W)�U�x~��-#J�ƛz	��%�T�������U0En���ȏC6�OV�|˓�0����1�����@}�5������j������<���;��CE��8G�6�O�x=*��|��j���KG��*�
j}��@�c�h��y��s����2ځ7؝����+��\��n��hc;S�	w �����Ig�ӂ��(�g:��}� ��e��bU�ҪE���6��Ϻ�ꘐp�Q 	�S׀�Z	�88�AG���+�YDxEխ#Ge0G��Y�
�r:s���b)c4*�_U"�`]�G�Պ���߅�����֪=��
��-�9F3�z(���'˕1ވ"���$�Si�Z�m���]�G���d��a (���]�͑��x�=z��FUm�����(�8w_ͶI-���l c�&O�1����$�Q7-�&��oqYT����q"���l�JN��v��bk�����������3�~a����l���`i��_5+D)6���%8k+���7��r�u�%݅Ք���AXU�R��q5��:c��<X�®��8ٟ��.aK�&ꏐ}��)kh�p����������� ���@�\�<��O���r*(XXm����)�b��C佞����2�,���hU�p���v@/�`���!h*Z�IE�'�-N�%;4`�A���Q�1{�@p�bd��+p4��T���,�\<D�&NY�iuj��j2_��C�%��Y~�0�9[T�SF�� �s���M�0�ڴ�X���ڣ�ה��]���K���3^\�{�Un�����V��gf��OB5�pes�9����������-��������(�n!/��I�8�j��s�)�6��L�umst�
!�� ���T*��I�����F��������#`�s�����!3�%h�E�X�zU������O~7�S T_QMek�1�WʿH)<��hE�@S�Ǌ���o"�!�.�Q׋�$Г��7�$&+Ѻ�>w����#��b��$��u�_�G�ֻm������?^G��
_.�U�'Ⱦ�Ò+�h��T���`�c�6��V����F�d2�ʗ�\E�LP��������~�K��9> �N)�͌T~Cw�VM�H.Y�f���#�.�r������yI�ѾE�81oK3e��i �h�Q�Q�_�2"�.! �ϸ{��Z�ٙӃ�O�����#1��R�ОsZ��Pr��:{��6͔8/�H5��D�:�W��Q:K���ߘ�oΨ���-�p,1gY+�;�S4g�Dӣ��"�Uu�Κp$&}�`��g$X�h�Mv¹�E�<Xx��
��r�FY�a���wfB�q�L<�38;�(�Ֆ*:���-'=Y�U3Bs������;�|Z��W_��w���.�T��+�Q!.+���@����y[�w��;�c_���ӽ�g���i>x�}}�?h�<���N���_	ߦ���W^��N݅N�	�Ӟ�"f���&9Ѫ�S$Z��0�Y*;OKP)b�r���	�T�oWn����q���7ٳ]����E����_��R���2����}2�@���Z!,DN����+.�3�@y��iI�3̥����@
�+�~��Z��d���+�H�m�Y�%��8���N(»v?=>MQ����Jm,��! �Ch���:c��D(�g�C�`	��g�h�R��V쨔=~��eu7S�i�vI�ұUih�O���YVrB���^�f�����<��k]`aNs�4�ۦ�(�-L�w�"��
�y?[���A(��dޗ��;|(0�v��VC��2CL��8���S��X6��"�Ďў�N�]��A�:
�F�'Y�"`��ɀ?ϔT� =�U��e�Xh8�m�v�)`�Ff/�g�(Αbv��I�Sk��a_D�����NkdWQ�)��U��^�o~���7)�A�l���]�1g\)E�,�]ޜ��SN��40��"�����L�����;��߬�v�P+�!���~���b��O l��)0訮���3�MT}�%|���#	�=D[���#:�� �U<};Md��n�8��'�o��Ԇ���X9V�#���gO�M�]����q��o�	��H��=�;������7ލLo�Lv����!ݯQ���{yR���[Н�j�AM 1=�׊Ď�0�^��ŵ�d�t�&����K/�gL�=	Ք�9��/�]�
(Òk �-�?w���&���P[�0/F���-�����򚒲zPC�|Hu���S��<[
��b?y�\��b	e�{&!:o�> 1���y¹bK4
���=#_�'������nh�J �=�'9���G����절-<�rltPE9!��x�522�Q�)�Lx{ ��	��?�qo@��c,���Е��j�cf�U�s�.e��KC4lׅ���M��d�[L�&��8�Yg�D�M���> �Z4|�d0�>��q�J^��U����0��@�(��Y�}V0�F4R�yh�����L�b8!�>�ʻ�{�!![�	ghC�q���n}����� �¡����zwa���:u&��t�3C�7�W���~�f縯A|�1�~k����wY���w$c����ܾ�(�L�Jy(��iBz�x#߸�y�6cQ��D�U���e��{��1
Wfpn
_�hm����L<���\��w䒿�șb�������[�O�?$��@
��b'���kr�Ԟ��\T���j�$���$�e�p�m	���q�f�0s�^�_K;��������M�OZ:��=��~d��1v`-��F�v��V�[W������0�J3ă�b���J���4L�)>�݆��������F�{�s�탇Sn�~�M��~�޿�+�52f2hw��é2�I�����(�������q�����A�}� �_�i�·8�-����0G�!NZ��Ad�r{G(��ZF�)]��F}���	ս��Q���r �U�<�3� ����� x�9�~No	!!��|^�<I��4����v*g~e��B�q��*˳[��{"n�@��$�ZMk��.Me���Z��k���2J�>� ��A�x�C �>K��1��;�?�!��C���o9�˖b�HM��r���Dzz�c�ʒ7�������ML�]�y�K|(�H9e� �f~&�<�g�����.�5K����?(.\o,�؛���W��Z�ڎ�+�Fk����:�,���|/h��>�dz+����Y�z��`7�#5�̥ͺ�_�[?f��2�6˕S��.|FrV���w�u5��D?�*Ca�x�l���b��k[�ħ�)!�8�)y����Tk�9��L�Pj��ٜ�iiȔW����5w%�Nc3����c�H��@����#��M���sU-���Zwƿ T�3��R�Ӑ�/i������^�+c~d>�La ��ӷL8��<P�3b���·2�2�B�8���vt�qt)�� �]&��M�2S�UrfTo�coJ�? k��V27�;x)�Hz��C<{�?�隀���twT	u�ax/vu7<Zd�V�`Nڭ�Ԗ��E�����)�s���m�q}�^�Fl^ڮ4��7�/�}�뙾�-w\�I�ϾK��Bm] �AZ �ډ8k9����@�]�����8�����Z[��rٴ?��D#ݗ͏./����]eJ[+�t� ��54Z����)WS���!�v����2�ѷ�o���c����VzB���: j^�m^�w�n�wx6���,��c҅�x>K<��0�H�Mf$ɕd�ԓ�]�[V%�I�O����Χ�˘��n��XYDB"��\��K��Y��o�0��C�
h�����vI�#��b���irX��f�>�}����=Ϙ�єZ_
W���Wq颦�<ix��;?Kl�6�Y?���Ө��Bb8LI$I�3����\z5�R���Ks�I4�\�U��4��o//���"K��o簦�mn�̭$���I����2C�:���S��	���M�<��y6%Q��U�L�M�@��}�����ɨ?��v��s�{w�[��7J�A���Igy��N���1ۻ��<-�@�W$�գlniQ�� ��?��z��6ۘT�cr�S��M� �1g7�#��̛*.Mh4ݰh8]�O<�J����q��0���n6ն�����.�JE4-<�V���`ĀW<�H�7����AP�2�y؟[��p�K��@��!��s�ho��0�;�1e������ꎚ����(���O�XZ�Ay>�qh�߰_�1s��>|:u��ޏ$�j+rn1�^�p�.YC��hYs*�ly�o����C��Qc���)k�����d���K�A8n3G��.$(��C#"��`���z"�T��!G��"��g�������R��Mp�@�&���W+�s�4��8��J���$,��-o(?�.F�|�����F����Y����d�@iKK=�ʢll�qF1z!Aş+a�����TXa���`�i����pt��,ۻ���m�wM��bR|u�,� �;��}q|[����f6X%y��Z�R˂!��z�n��ˎ���"(h��{�5��3%K��F%�L�L'!!AU�i	�}/p�l� ��+X���l�"~�X /e��+��^�N�;�-��i@0���Kn#P>�pn�YI�g�5vs�UJ�����F�?����x4�UͦRCE�ng�ұW.�Ά��ډ�y[<�cѴs'����
�q�FZ��K�ɷY��vE���?93�@^��j�U��ҏ&�4��v�ėz���4��T"E44�
%����~
�?�/���|(c0�,⧙*V�)r����z߾�F�g�RD�����e���UnH��]�����?rrĲH�6��#����% 	�a�"�.�.�J���D��p"׼@�,�~����e���� 2f3�{ڽȢ�v�#,�8_b��Q,'�~L�����~Ș��BYF7z�e�}��y�I0=�d�Q�G.�ݏԝ�Y-h.�N�iL������E���Bą0v���_�Oo��H{0�f0T2fTr�3B����\�#��X*���N�)*��Y��<�j���-��i�7d@�����Y��u5�����44�k�o�,<N�U8��>D� �4=��6�zR~0��-�r�(���/:(��I~�+�s��3���G���:1��`�����1'B�Ú�i�I=�X��d!�V�2�N�� ��#�Z�A����`�o���HRԆ��Vo[����8t�}l���(*�����'Q��t`�p����� �4ڢPu�3=R�uV����.Yٷ�ނ�-�~*0Q$�����/j2�벱~�nai>��N^�hZ��*���g�"}�!Պ��k,C�`�{�唜��#�FDh��Ltk.�F::0H���ٿ���!��Wkl@=���!�|�����+��1�l=��=��j6o.��C�{3E�(ɟr2-[E�h8���gU��"�?��O�\�qllC�/�y���Q.������y�D.g��'�=QV���GK��Q���������xC+!���r.�� a���QG���}0�7Y�`A�:{�0�����q%����~�Q�rH�2�
Y��BHN`�����{�Vp{.���}0����%R��(���@��"�Z��R�5�߷�^��q��Rļ@�$~�T��k�L6/w�>�;�]�Pg� �EL�іҠ�ND&é�Xo�ab$��٧��\����m��E�h�Sg���rO���Nݒ�v%��ʰ�<�H�"ą!̬�ɨ�]`_F�Ji"��(��a�1�u�����A�d�]���ʠ.�P%�Y�\+�����D�ꨖ�ľS9����,b��%��|wxu�R�o-d5���8��Qf���N���0E�;6�\�n��c����i��V�!��� K���LYj`�^�!!�WN�7�ߋ�R�aX���q��Y4�)��nMF=즵"���7�����PBD���GV���ꝣE:�v�@7�w��AB=N�KxɄ��2Z�#�`�2E˝[��G�-�BD1~�Q^^Z{]��Ƭ�\��r���c�w��D�Ѕ�k��]a�g<~��?^�� M�i��A�L���4ɽ�X+��ѻ�6��Ue��FS23�p���ro�ٖFi�{\��wt�p�B�F����!ĲL��-*�8
�H�#�:C��t�v�˺���!	�S�+|�ya�҇�I��O<,N�W�q1���D�nBbh�����ʛ<�D�A:c��n�����$��R�+p�z�F�[�	fO��e��u�>�Q!#���@��[��b$���$�R�yq�DB=��e�8_�O���R�
�בHz�K���`�3�r2�97�̼�ez�1�̰��\b�z���@�`�խm��2��?�g�e�Y������2�FӮ�Z�'���>�Cپ����sv��y�
���
���^����a#�
�I��أ��(�����}��naѫ?��Bu�S��D��]l"�d6I#����\y�	2��A����M���4��o�\��(U[�bρ<���d��}��!S%f�quK�69�ki�x�QX����F=�����s?���%���g'��P�b�|����Br�3��U��)���$D�ȸ;�����Cj�ć�S�y�6��k�i9rk�*���j]zQ<Lwl\���IA-!	�۶H��ʆ�K`��}��� �71B�T=�F�z��Y�$������[��a�����a�A�l��8zpj.�u̳�R�����W|�����+��ʤ��#gl<þ9l ��j��r�53_��L*��H���R��+��y����4�?�E�5��cL����,�}۰X3Z�}t�vW��bf�n7��z����=5��<�!� �����ɵٚj�����{?��N,z���+麷�̴��`*]�cr�it��u5�M�UT����o?Vx���٪��I'�<eu���cD�݂(�%��yB����I�xL6���̿L�-���i"g�!ЁH࠮�  =[k>��֚3(�4�OT�QL�R �3�s��6Bʳ*�q�M�Bj�mݩ�*�O�0~�$'��.��e�T�O�ew�-�o>#ת:����I��F
	P�N}ϫ��g�<�����є%��|���X�Ǟ�uW��}�%)X�4oГfC�Q؅���,�"�rY֩(�I9�ƨʎ8�Y��D������}0-h���Ɵ����k���A��.HN�k!5c�QYĲ���r�B]~3+��>k�)Q�@7D �-J�~᣿W�ڟnЊD��9f`�T�o����҅��f�w`����f�4~u���(H�*G]�Ɗ��k����
V�Ѻk��.�����TT[��F<}�������`�x9-*�Y./#R��J�YS:|T0�ѿ+�M9'��Z�7��o�4����(N\�΢�K�\�/@^�/��0�0�y��8��%8<���{�K����2m��^�E�G`�8�ʊ�΂z*�',�6���A8����!s