��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]ǂ��O��˰�	JL��	���md��{ Zn=�S��.p�Ћ(�k�V�\* �*�3�q��eUT�eW�k6~�_�hX�(Z�*0�5�\dX݆&!%l��}nYv=m"���NR���	
`�k�c4�Q|ʛj�2�=krP{،e�W�ׅ
�˟�I4D�P��Z����MZ�Q�"[{ %�cع�N�'w��`�(���jܥy6�G<�7��CX�ɟJ�JhU�z�[��BՑm��Y��e5�v��bi/~<�`�����z~ ďU�g�x�M�D���OV�����-%[\ǾI�-�RM'^g'�R���2�Zf��d�^��D$��f�\��<�*
o.h�-��
��M���ٿ��4�����;x�4d���*K�
�FdX�uC�k2���[I(� ��T�,�n
	]����0��i ����
���T�-�(���/��H�/cwMA�