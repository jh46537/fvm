��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�loa���u*3������~��
R�:\�K,�ǉ."�"˞\Gr����[p*��%Z0*�)1�S��Idt�r�'q�)t�#U/N��{ZA��/�-�tTc�z���lf�XdT�cS8�1��<��[Y�b_�`��A��8Z�_K�g��6�F&A]z,6�>�_�P�_����1���IA�dJ���Ē	�����O	5���f�%�͊o�lR:�$�`���G� � ��6cC��T�2n�S�OJD�r��J�L�OA�<Qdc�{�'u �}<�q���' *|��"�O@XC���RvHHT�$v�A$�׳@}��ڐrt�5UU��o��Y3�;a��:�[�����<�x���]�~������F�Sg!
�8*v���B�Ӎ Tߗkj3^Zx�C}��b��U�9\�9ިԷ!a-4Zʱ����������҄��V���SC��;�d�z
I�=4ו�Jn6�m��e=Q�#*�2e�e��pIj��]9\ޓ������}2Yb9l?�z�z�)RN�^ !��bG��R��TE7m��zDW_�uɺǹ�x)�x4(ow�K�ǫu�~���F�?�T��� �b,��
"��g��E�A-� �� ӣ�zu _��c�v4�?{���g���%�5���Q���wa���<A���jT�Sa�B�W&8��g����Ś�����SyS3.ų�=[m��"�M2u�vC�<<5���Z�"g�LʋI5�U��vD���.Ot����]��l��eve��/�p�ƫ�m�aO�&�x|����,�]��pߺ)�|fZ[�!sjcQQ�F3��T()���s���:��v�crpگ����*�̡�+5��{���F��ϩE08"�=�U� ]w�/���C��	�:~���$H~i�j��p�K\��#v�$� A�e�a>�v������RF,̃���K�� ���ԑ٨�Ƭb����JarM%��I�	%.�+ǵC�v�'q~�jJiS�f���
�8Z��'a�p6*[�����&y�}Js.�9�;}���t;�0��@�kѝ����� ��®Α��c9�΋�@M�M3�LD�����~mh�SɼR#y*�ݼ��++�Y�	�&#��;6��?�s�b?�ۈ�tD��I��y�)��O�N��y����7�blR�)���,0.�tn�����~v"�Y�����G'�#����d��'���̳�?D*������zH�{n{���z�j�6��ZY؟�����l�Ry�zI�PF� k�W����z���N�V ��˹��k�����HkD�;�o9�r�{U����72|q��bΙ���?`�O4a���kØ���e�(�AD����MG�������(�?�n��G����Mՠjr�P�,�ň���F�2EGR��=��$u��y�u��q�/�h�q#b�{c��U�$`k��븘\�����@Q���G?���]QOip��Ƒ�b\�*�*�Le�HZ3�
��V|�Y��;�z�k�D�`�^݆�{+-�&O�ڦ��K�7f�[k�ˇ�UW(-؎N�Oǔ�4�5����e����Z��%n���SQ��"�	�z��j�l��\$<�^����o�+O�0GtSC�y~�I�T�V�X�#��BC�9B�/���Y�}��e��wd/���t��:<� j��?��9��,&t�k �h��C�8�?�C� �+:}���4}*s}��K�J3
m�%;m�G�j��Cb�}���f�Ȑx�s��-dҦ���PR����������OmԡW]��G�q*�^�]�aiE��}�*2���)��\>obj��\����DcFs="_̓�c�V��R@τ��v�&2EH[�|��-�4��Pv�h���$�l<�$Y�~a�=Z��à~c`�����$�\;��/���ܤ�SSs���:o���y���Gr(>��i ������c�ȃI��a�X�B������ �cv#�?�ӥ��l��޹����^���Op�=�B���ϊ4���|�;��h'�	��jove�����l61���[�6�{�R�&һ� �'P�1�Dޓr!�a)Fƹ��j4��u@q�ƜO0 z5cȹ���@�ۧ'���;M!C�y�{m0�G<tE�`�g\ּ�-�q��ᑭs������j=@`S�ah2�����	�X$��5�ҭP��٩d��j��ZDt!]Mb�T�x��C�c���-Z�QG
%5�*��|�_��*� �N�j�5nj�\����{|hq�/�zq��DrMO^
�����i> .[�[�.�W��̰9��#�$bdji��}=��X����2�~��"
�$�a=�A&��ָͧy.����ޝW��Y�:�Hdcޡ^H� Jv�*�ZL���&!�6+�Y=�������\��JL�5���U�)��J�
�8��ֹ,�
�E���PD� � ���A͖=�P�� ���vG��)�H�V���ݣ�T�%RIԥ�	�v�iʔ��!�m�S���W�;�|9���NN��oCY�������x��y� Q�
}���B���Wu�w ���bUS��I~��X��cO�!�m<�!
�A�J��|��%����u�I�U��b��VZ�G��{@]U$&�Y'v��e�5��y��~�(�Z �^��`+�3�F����Sp�|={Cnf^��/��uh.dY�P�my�,O`{t�B��]f�{�JR���Zhs���̛|�x'n�m;��������0��"d�+28@.!����9�D��g)�Ze�N�?,�fe�_�zK�=�)�@k+Q/��WU�,H��X�݀�t���f��;xd�E�&�ݵ�5��6���K�-�m��[v�k��������^���~���M��2�T�9��{�O��?�q	ut|
�-��_W��-20�]cO����{�uY��;@��x��:^x.	@?>�����48!�������ӗB�������YRq߈ �	���b�bc�@�آV<n�_u��0��8�%��3wS�0�^������+M�;��Qt�d����ha�øO��
����#���M,gm�=ڛ$�q�-c�U��qc�{K�6!x.ҭ�+�7�Y/�A3O7���N^����.��V8�: dhs
'���N����S����gF4��&\s�C��Z�è=,*]�g.Ճ���z��fj�t:v�j*
i\���RǼ��ic�$��*%�k�(g�9��\Lxe�����������ծ�1kDF~�h/_�9b}l�����������JU�ݖ�%�m�M�}[!��
�it#oYEmb0w3�g�곛��Xt���=�|O�~K��p$��r���`�l׸�A�2D5���@��Ϋ�� �j���0���lY	3�'�GĀ[�?*���^\[lW|U��~#Ǥ���̲��gfê����N���J|:�kJZ��ʃTK0� 7�����8�?q�#�����K\�D�O�l	�8���7�4�M�S�a�
�B [2���
|�'�M���'q	MI>\e6�fyv-�Zi�S��:��\p�F������E]�
��s�Y�*��#�А����8x�άV~��e��8XX��7P�m���s���/�j_�:���B���Uf�⮍�)Q�U�oz�I{�p����Yy��|�����ǋh_�Fy��/�io�rPϊ���n�����Ŗ���fX̢Xgܳͮ�m?�]��I�wu�nٹ�=�f�?kS	5����c7�m7�J6��$�ǢZEޙ&]A�[	Ok�_�h�b�g�,��+h
���kB�B�و�`zE`@J}����B>�`R��K���Ng�S�G$�#.����nLp��~�Rf5[�Z[q8� q�#��S.U4E�T+�2��yp�B�Zt���"�f�����J;8�k��7�&��xh�N?�	��!6 UǮ����s�#��̸$3��KK�="jp;7&��ɨm��g���O������f=W!���N&Z��a����;aȢͣ�{
��[�(�<���4?��Q�£�ߵ ���̼x�}��m����Ϧ�>W�Bk�t����h��tD�)�e���I�}u�L�>w����ضѡqdb!�i�	ls�^�$SU���+�R�ԝ+�Nx��*SD�c��_���f��}�YX�������6w笵PEC�!��IK�"���C�[��������|S򷼁`���Vt���
^D�|� e�c	���D�v�&���i�B��&�uf����,��{^�^	k4Լy