��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm����질�95J{۠�`\j��G�!�<�ց���&�l,�y�ʰ��D����&��ejP�4��:�D�BH�v�Y��0�����"J�������W�#0���1�Ay0����+�.��g��z��Peˇ�;.��㝨i`#��3K��o'ͪg4��T>׿?^Ti�j9`��j��#cu�����vJ���J�����|N(�on�@u��w(�������'9����'�(
Lh��*���ù7R!�߹O��l��~J�v�8U{�P�{י�-	�3M�b�s�O����	z\8�L���ĺ9�!y�9�R�$eH��>P���1�?*
2U���W5�҉���<B�vj�dW��j+am �Y�23�]�����;�K��Xl��!��]�(�S��Oe^���%��)=��x��@�@�@�WvF���d�➲��� \���"fK9�'8�}�|C�8�z6�����6�@�L� *
G��)	\C�K���a��?'��ZW����C�j徚�<�<"2D�X|�YH�eA�O)2
�y�6Kҽj"����|aO�Y��� ����n��`W���y�5mf�~EϪ��x����H��̼h�nG�E��:��j�ȗ��2'����JWY�{��p���s}e}&3���I��k�7AG�{�1���1�3.{��
Q�#���z ���:0�O��q\K����,��p�״&�CZ�W����X�Q�k��}�!�Z[�N����X��̥ܒ�~>�m�t���3����ߨp^�~4�A��Y��iw�(�;�N#��T$�O�y�-Ew��T��D|(-r���o$e��C�J��9�.Æ$+O�N[u���^YT`s������P�ӳ�>��h&��O����pUU\�u3J�YX��}Giw����/�QW/Qi5�2�%p��y��ؠ0L{�}��D�cIb��R�t�;FwG�}B�h&ѻ����6��e�h�/���3��U?� �t،g�Y���7��=xe�$�,?��k�OH�aP���� bQ�TI��n��ݑ��.�'�춮6�c����T�ڞ��p�-5�Y 0�?�t�˫ɇG��oi�E�ޔ,/��P@����B�mD�,����)�Ӣ�(q�6�FBh/q��}�ȼ���I���?��q{̀�չ�p����qv�t`x�z7Nkf/��\�������_��.䭌��~�y�:7j AZcb�G��ҙs����cߝ]bT4�i�hB'�$���v��\��Lo�wEq���X�}8Qz>"�9�n���H�x愱`�s|�����`	�s�c4����7s����/ś0/��������|b�;Bg6���HQ�O�8���\��E�>��p*`]`M4uL9�^�+���q%wX���(쪔گ���z�����xF��[?����~��H\^��n�D��L��݁$W�戮g�Bz��v�#�B�g�����I@):Z�ڤ����wK���mW`�:�_�b?{��}�iL�����Q��6����Zl{b];1�%E#�������/@%
���i��9���h���G��Y���1�F���}4��T܂m�*�*��s�@�'��S{�<�;���<�W�*
|�K��<p�]����Zļm�ob�Ĵ�H����_}�]�|nU�l�N{��o՜�'HK�]T����_�W����JxU�G�Ua�/�9
���)e �1_��ό����wT�ANx��ж<��%����A��bΣ��b��p�X:@�7P�͡�0�2s<��}NR説7> W�.~|��f�rѴ��P�R/Wy2I��(č��p�(���50�l�WV��� h��*>l]�f��>f�݈L�6�1��T|_��gqЇmC��u�]J&���R����vƞ&5t �9�z=����,�]G�ME�l�u�R�	-�U|�N�B����琾���@9զ��� 0	3w-|7fO�	+�?2�Okn��V}3�#;=<�JO��y޻�O�In�	#��R��&��9��ȃ%)�i1rb#��7XOmЪ�Sw���u8�������Y��EK���po�\N������Q���u�b��vϪ�(6w�_�X�RTˍ��;�r�:�z:%d��
߼��d��)�e�;K8P�B �B��8���M�(�^1�����r8��fQ��v��RY�K�Mm���1�̴������/a��!���$ޯ&e\ Y�sC��k<��Qe]��̼�8 ,�nO�j|��;+�}f�e4P6��t�y�)�tm3 �.�a�_�5[/�-GG�}s,��W�z��d!EO�d5��|B�A����e�w��sH��7�F� o�A�h8-�J��rxJ��_/�n���+r5!�B���nqr6�s��̸۷f
�z�S��
������t=n��v�\o+��bE�{�\�/�Y0��aL�)!�\G�\�e����%(O/�pJ�����Q(	F��]�=(�q�@��g|��W�P�N�@���#����16⦈bȷ=�B��\=����f���b$�m߁�8n$�9 z؉g¹6�:��t��������XĪ�C��[Cp2|��Reh������mUZ�bUH�]�t3$�fgd��B{f��c�i{�)9�li�~�Xy����=}]�>���륥��5�Ǐ-�vf�6Wu�:��*�QXa>e�Z�~�*��w�V ����ʀ4L�����Āv9�]�$���c|��֣A��b��#��wA:�5SX��!:s�H*�/� ���4%y��g�}DN��<����1$��z���e�?�U.���� `��qg4�����YqZ�a�ۗ6�_��N�Zg6��3og�$h�c�8aY$l]N�`������� �����Oł����/����Q�t����)īC�6�g�G!��(]�kѤrtNNˏ���Ɩ)h�7��*��a废�fP�o�N"!m`�ʺQ(OR��v��ʕ��qE��/jY��y3���\�Jسz��=���[/r��C���&���T�j©���T׭�:��jI����TU�H���{�����7���Ύ�w�BM̯s�7�C����_��S�XhR�(�j"���»��;/� �IƘ��� %�0[�Z9���F�K�Y���H��jg#Zrh:6���l|�,0hhb^��g"$�{Mxa�v�!�AȤ�7�+M�}�� �E��^�d�	��2t��8=���m���d��y�ϔ����Z���@��6ͼ�-,��p�^?."���J��hg�nޡ�#��W.>CyR_q_�~��m�������{nK�/��Y����ԥH�g�{�ϯ�tUDGL�ʟ@E5�w07��t^b��$ᎎ A��ٳS�5��Q5U��O\L�8{A��y�T���Ap��u�z���a��CM5Y�9�aD��$��$Vm��:�p�Z?���j�f��L��-��� c]]��@Y;�pv��vUJ���;AR��hpu/�NwW4u�m��-����]���X<�/|M���Q��k�4A�Is�7���IU��=�0*A���&�Wt?8��r<r��j�h�oo4�<�٬d�<��^�>w���懏�aJq�E](��Xyv������y�q'x��*T�\�㟨c��ۀ�����B�hʟg��M1��% GG�0#�-�-�c'�Є(���\P��}+��� �~u]����G��ƸP���;��ڇ��*��~!�$H����c�w�-к��D��D�3<e�͙#s�A�M�0�k4�t�|�5=,���������G�]��{�b8���p�$��w�An����bȀ�R�e��f��ƞk�49~�^����]י���0l�������Β