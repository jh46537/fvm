��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�;<�T������8�l��s��MC��w���;���%6f#z�*�z�ѫ#X}��_��pV[ހ�W�W_�^�Ʉ�'�l�o9�<v	�H���d��et��-o�w[~�?Cf��`,�Z: �� �
����;]S>)����i`Ui#���_����Luk���J�= �0�[7����Z�5~)����-�C�! S6:���,.��V��6K:�#;;>��Ɲ�>ʼ �@{�(GoRRA@7�9�['
�~y^��l��t�#���2g�`8*7?�E�sc�F0���3�O���j�p�_��;n�];%�=C�C���J�3b���FȒ���qU�Cӄ^�� 4	.Hu�:9΢���(�X����V'��p|��䔃H+yu'L����91�o���"B�:���:���m��nq��L����gE2�n���ġ���Ԕ����^B{E��I�c�?��_�Er�H1@��}�Y���-��.`�g��"g�%��'x��Q�3Cd$(ʚ�oF�:��Aϒa!M�s�e��a�m�y�v�W�
�c���|�ڮx�ˎ�w�w���4�e y��Ve� Nؙa�m��TK��8� �a��+��c;w���ς9.ېq�Z (�3����.�h;@�T,��Zp(z�&PX�JI�/M��[���|:on�[�:��-�sc	�@�U�h �v (}�L�+�!Kt�&�[q�#�2(0J�E�hӿ�̀�PK����N܄�r�_<��[i�q\ ���$����֨T01���t�S0��ꏩ_Z�+"�!d�
��4��u��wΘ5c�UČ�Ǚw�h;,�](J�W������LS��i3�?΢���"��+×ة��DI��Aꀾ���w���~=Y����8�'q.f&���*]�! �`(:�a�I�1ƒ��J�=M�Mz�
�[����� �zʡ��^�E�!�j���OA���oZR!�#n���~m�'!r�K��<_�F>t-��nI+����q9�i��̍���r�7�6�	�J��@���j�^�w�;:�x�Ee0=n[@���ᅥ�Cdb���L
or,H=M��%�߹�R*K.M�Hz1i��4����u�#�Z���Q���zŇ��rb{��t�b�������P�FF�}�Q�����f)�v�_����I�͖X��b�%"�����=�9�ݸK�dr�z�w�
�ܤ�!���Mo��<)�u��[�%�`+�"t.UF�?ћ{�X8�O2���J��S�$5��r
�Ƥ�P�sg5F9e�|�/��*��:G�[4��kcݐ^ƿ�8�C���F�Q{�ء	LS���;\�[�*�n9�Ŧ-v�}\�s|���WҸӭ��Sÿ�.�j�Q��xb�H��}d��o���������K/�ofD���i��UC�8�s�	M�'.!�y�΁�m�hia��"r����`���9��,��?�nU�;�bl�tF����MEw���M4Gx?�bj�>ܨ�M	� s)b V��{y�So^�t�v!f@k{kU�97�)rq#'��6s;a7b�a�z^�$��H~`�׶q)F��o���C�/��ϥrU$�̲��kG����v4������Q:^��ފ�l���޶VF��ׄ��e�뜫�X���C�^���'���� ��?�K�ibW�:Os��A����9v\%�0�q X��ӎ�"+��T��~��W�����׺/����a ����R�LLE)@�DɩY��\C�l��i��V�[ J))2���� ���5��,�ӳ��e���PR�z'e>�D�����^��,�8�2,��z!Ve����)i��p�N�:����,M��kd�������}�!n�zq�[(��y�8��ec�u�Q����6�(@����2��?�J�Ў�� ��߾;Ηa������1���Z����<�o�Y/�@���4���Mk.h<�)P�V��"T�"Ǉ0�Y
�A�����<�Z�����K����c����5E��o���(��i96�}�R���"kM:*-ډ���;-�w�e�qF�E�ԍ?����]8��Y�M����j�,6�|�S!�ժG��@��!�L�u�����%=��+gK�0M�����*Qٗp/���a"������y ����Q|���l��s_?u�,#q�dX�b�\�{+ΜCwx�U��L��+1�+z�\�)kڕM�fm�E�t�&Ӹ*+ku@�� \��ׅ�7��p~���hH�m ��6�}D�9���hS���V9���e�C������TX=nxhJ��iǗ����&��Fa�Q�㱌����9�� �D��ƪ�.�{f��E9[֦�R2������_���*�mQ�t�Q����r����1_�Jzg�ʑu�y6�+��眻���pĀn!'�z[%�4%��4A��&�=#TW!��zB�.;�WC�+�y��X�1��Q�6!F���e���I�q�������/�[�qƶ�E���J�3�D�&�c�aM�ܣ�!Ц�+'�6�eV�.�	1fNK頝zD0�Xek�cc80���k�X"u�O5�km�97Z+�9	N?&����SD��?3M�TB<ѳ-�F��g���k�����ܼ�^ogZ.��az��~'F��q�]m��],Y2�\���!$�҆�FvgF��n@�(�ʡ�ױ���:�;74fȕc>����c]mʄRy�W6ʑ~ƪ��'#��M��+�B�����R{	*�)x(����%щ� ��z�%����Y�	w���z:v�+���1�uW����x�b �81�
wx§�5�������9>��喞Y�
��$�RI����(0W6�q�W/y�C���Q�4=,�F��Qdm�Y=&�Q������8��#{ӆ����m�g	��oe+�� R�y�Zj�g��#0s�������O ���5j���b��3?��g��Ǝ���*/r�����(��m=�&��פ����JE�կ]:N�����[�S� �6QG��D�LY����7(��B�?;���N�P��n���d@�K��Pp�k��v8�����?�P32Wi���fpP��U,|4�L�P�X�i�*��[ٽ|>�m��~�k���kEH';J �=�p?��l����	�@/�[�~]�[�U�긺R�E�pAUq�����[�MhyX�#f���Ĉ��y�h�따ļS�����R����u.�s�`f�\O@�Ϻ�,)����bKL�.�/,�S�<D�����w��>'9auN.�nŖ���ױ�̍�[g/흘��Hͳ�zB�9X�:�ML�V�`5��%=v��D�Q�C��!�.����4`M8K�4	[B�/�x_��\��z���o-G`��Ǡu_�֋,�yb�
�]��bi�R�9�G��B��9�Ԉ�&VaX�'� �#���S"7B����E�щ�P��B�JZK���("�z�ۢ�n�I8�ǹ�c�Ǜ��~��F�In�"�T�r}-�>����A8w������5Ց��73���i��1�`��6��M[��������׹�Eh��{՗��u��>c��:ɩ�4)���隟8�8dc��X�L��o�sU�t��^���|���jiڵ|��I�E��@\ʲ1�<Zmq�x�O�g��������t�*��~���	q����;܁��%P���rg��f"^'��#�&mo�7�z�x)��lC�p��e����6�֞�b�C��hmӕ�	�n���C*W"�d�g�����׮h�RB���>=�)-��m�Ɯj��a�>�k`o>c4$ޜ�a�З/3B~�t9m�u���2a���-*����d�;WI���pO�e.�6_p5� ?ŲA�˝y����e��ʱ��X��|x��Ӊ���S��]n!5����N�!dW���:�D#�D�(��288���� !������S��n��c����p!�����a/��M�XA"WU� |�G�4�g.����Dq���ץ@�8�5*Ͷ����$պl����첫�{l�5yq"��Kbbi/�$d��h�.��G.��XI�c�Z���P�P/y�R�"��ۚh6Q�ȱ�/���e2��B8W:
#��	�nE�����n�"�g<����o���n�S���S��m�����}3gbqj�E�sA⽖���̰Kk���V�d�1A9]���G���N��a7�&��_]�q�_��u�-�g��͟���}���
T�������m�3�NQ���i�����k�e�mU�J[�����ځ�o��؝�VX*�f�B�c?5���O'�5ǎc��B�%�55��$��V���#F{uq�Ӭ�����HR���~�f���@��ߎx��+��hj��)h��}-��Nc��F.~�7a����D"�!�{5��̎�m��5la��;^Ct��B+�O�+�ܨD���%��*����)��=<��������F̖"�Y$,c��P� �=��ӰS���?#���I3����5t���_Z��g�S�6���ifl<�wF����ݒl��]D(��|���xA(���Wڱ���K-v2��Y'7C/�Hf����u��#�B��.�l$>M=��v��"���,N~�.�
E�ˋq�Vk�3�ȗ��Ќ�Z�����Tꀝ6t�ګrd�旝w������U[@v�:�P �>���=A��AW�q����AB�L[�*�������o�?T~�i$	����]4�K�\���j+�0Quǩ��/��<T�*��d�q(ԫF'<v�M[NI�g���d���jg b���;
sxۺ|���ΜN���6v�@2������� ���]��6v����8�+�?X�`8v1��>Z�7�\x�:�+Uj��Ab�J]6�l� �#fQ-.��/ B��I�� �_�����m+V��=�]�6
���4#�`t*4\�ĕ�mf��gu�s�{@.�X��&���{&���7��f~q_�c����ݽs�LK>*z'�?��o,jD�|(B#zQ�W\̵0Fr�
Z��0���*