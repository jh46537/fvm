��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>��������ّ$�*X`F~�������><06�L���\�D>�WҎ�����r�.~O�I�V�X;w�G��ts��K�5���t�7��R��пr�.r���x{��}sbeq�XG|7 ��$�ڳ&�e
�=r�$��!錋"���ۆ[�8����lr���8Yi��9���eIE�(Z�)��VJ�j��?~�	��c��R�6���/�WC*��B�����-~��R���$=��&����O6�F�~gh��\P:�w�o"Z��{��ܪ-|$�EA���ٔ:�_JFJJ��S�B	*.�a�ꇔ�@�/~�WC(���&q����?��V~��A������(}�b	ѝu�%k!gŝ>�I8�s)�u{��>kp�Syʰ+�� 2����=��D~0.i4��SJ~��U�h��ERc;��@�p&)Aǳ)��� hU�`��ߨ��a�:m �7�8�M��h�E ��sY�"H�7�l <�~>��ʻ�[y�N	5�:�C`��`�g��u�,|��z'<�i��a!�|��25��0�Uf������e���Yxy4k�YZ>N��5@�߳�V�t����9(�6�$�S����}���;��)7qR+�Z	t:�D��yf�R@O�%C;\�1U]���7]֣�)�p�BU�-�f��F'��z�D��DovnN�y��Wڲ�)��k�3f��-nD���U�g�������9`�SE��́DU��:�z�J̫uѷ*n*$GOoǉ6�:��^��/��I�Wg�9e�����Z�%2'ї���Mh���j*�����o)Q��Ha<�0�SMܘ���ª��ߏ�()�9\J#ps��n��E�8�	�
@�X�V�=�./s�X�	QbtF�����-ԁ?���/��a�S�t��;��W�2�A���h����$^��{���>�t��ݙ4)'o��᭽���e�h�\�Ie����y�F��t���*"����(��ŎϊO�|��n�/Q�KM:Zq�zw�\��s�1�;�Y��#���[���a-�o��CkM1��u)L_q:����ΌBXJ���8J�>�*+�P�Y<镡��K0V`�mG�6;����莃@r
����1�\�t��`�dH1�k�c�+��t�Y�v¸���eN��ϼXN�Rp�?�)cǪ0�o�H�E�Т��U�%����.�t����0u�@�!k�M��4����k�b���������s��]@�j�����:�:Em�d�Qt���
�p�>c<�AhKX�)����Rak!�h9�H�A�2�ZV������%��S�V�z�3���x2�J���k����b8vU���_@�8��;c����� �a��?�U{�/}"�Qp��~/ں�����9�9�$��9:[�/����<q����QW���yB�X=M�� ^�����\ε�� ��.�M�o���!����	
o�l9�\��U�4
��������,O�
�Y�X��Dw���Kdn��S����ޙ�
j~|�M�kC@�C�y��s ��4�,�tf�y+3A�P�\x�BED2�i��W��0@�݃�#JK�"WNSt�g���8�.��Ԇtx�.����R%��,Nޞ ^7�Bp[��
�=�����0Џ	܁�Q��q�f�P˄"��rW���bP��aH������U�� ���@Ǵjz���!�F'��O��4���6�~Xw3��+��M�.�����N������� �~���5EVY�Dz���W��ϋB5�q`OYosL.*��:�,"(Y`�h�}0�)�N�'��͙-����2(����쒚a��f��po<J0��3��Q��3�[7�S��3�[�0T2����Ȏ؁d� @	�!JFoED+���Ǌ��Z�@[�,�M����e���Ρ�`~�[�Kp�hL�޷�Y2��u;��u��`�.'S���~R��zC�|E��'/��,����r3|7�����~���`���
a�0����4��Kv����{sH^��ɹz��$�N��5�~@� a�
�
(�N%Ϝ�B.~���i�~�#_�q5/�\�;��kEIޠ_���6��l��.�
�>y���L�Ֆ��i��dҧq�#���9V���I~�E~gW�L�r����qA9}���$wFt����[��#��o��L�*�,���|avR�p��"�{z�@���g�d�3�+;8"�S�_�ё��A=�D���d��6�Wʨ���	�����r��<�K��(l|��ǅ^�__|���@��9-75,a�s�ޥ�z������� w��9%a�7k)Ȫ&5S��X�
XFT�I��@;���cx���>8;J.f hI/h!Ɗ����Q��A�	���_L��Bai[T��ߕtp�Jp:�^XC���P�[Ӥo��:Cn�%��֙���\��}0�/vb;�����v���dqc�9ā2�:0�^��GKKU����}�
���G�|�c�Rǿ��)W���.�o�f	���?;޲tv�Å^�^'(i�_��DtՖޠ�ڸc#����e�����3�.U1��q�g�����`>��PS���4���~�^��:+�a�@_�(�sb����	D:Xܬe�x���՜������U߳�p�e��%�]#j!P�g�� 9J]FhG}=xzRi� (p�D�d$����d�0I��ι��Nf� BB�[��5h�F��q�JYQB�M"#J���0?6F�0o��(O��l��f�_�$��/
F�Jl�ۜ�^�-&ݥ�J��o4}pc�?��`u(��¬]�C��@t�Ff.���ޝ%sqx�ʰ��uo6@���T�p�=��.J�Z�nS���?�}M��o�y�VyA8Q����M��}X����1�|��jyno *B����۾��d;���5�F�E�_��x�D��B�U�~�6��lWL=�a y�����݉9J�G��a�g�e�E+h�$����~w�'��&���k��	���§J��{��XTk:����U?UI�ĸaD��aVG�Cp�[c�*r�u��$� ??�t��*�[x���#SH�J{d�tWX�oK��d��͸r8`z��S|나d��e��	 ;�'nk�����/˘Y�zpC��
��}S�{����6�;�s 0�d����ZX�0gsM�d���ͦ7SKh�+�{���q���K��Q����%,u��N����Cz֩�L8��?7(j�8��L�$�JQ��$0C��gǗe'��1�Md�7�y]�U��������@���.�1��C_��/�%�#���F�?d!!�U�B`RѪ'C�下i��<�	��+���3מ�'r�X��z鶸fJ�Z�w�0�~1�없b~+E�_���F�4c�P��'��b�m��9#�P{Bу�[�I����ڦ~v�)�խ�l��ٯ���ӹX6�a˵f��i�Ý�����kc�8S$��_N�τى���!آ3w���VF�G�\�	�t�۝_-d�O���;��Ф��OD���)�W]V�ӥSŌ�R���?hI�6,��-��>�Eg�' ��b�-@HF���>�h|�����������_E���{z�L#���^JuKIAI���8oC��jzN�ql���#���W݊�� {��Cޏ�����Ø��о�u�Rr��7��b+��m��Q	��ই;g9�O�b�Έ�����<��'�H����3��8R�O�m]����c��k��_�?���$�J����Kd�V� �O��_��
���E
_M��Ʌ�����t��k<��j��#��w+�3wOK��ne��Ѻ�٥ue���Ы�����7�$�\CYT=-�K��lN����h5G,7<z���>
���ǐ$�*M^:�8*�k��������SwU�m��g��8ݥ:���5���Ly�'����	��K�g�����4���_�	��f]v�`�T�k��Y֒���d�++�
���a�Ÿ]���M�ww��\��i����[�������F�Dh�D�+ת$��܊`�҇���w@<+�'E��X�h |4s�E~ȏ5�69��٧Rkg�Ʀ�\ĬũE~����V@��X~MX2r�/����nS`���J&�5�\0�Au9I��"��%���t�M�,?��Z����3��F+F��f6 v��uN��^��љ�N_J�K��˯6%ѡ����d��n�ee7�K��}&U=��>��!�zg�I\Uo%d�)\�DBJ_��3�s���;��6��0�WG3X��+������s�M����h�������a����\��*"$���'��m{��s���&Z�7O�x@���r
y1���Li�^�%eCީ��N4��MD/q�9�F�\�x�'����}��*����w�L��2xˇ��w��Ō0�F K�X��Ļ�QE#:s���f� �hqХ��-3p�^�Y� w�I���)"�����.ԟ�(�jÌ�0Ԛ��܆�Hz�8��ɀ���q�*��}&f�Y�Zm�3��σ<�*3�0{V��Cݑ������ ��#2�_���'%��h�MCyc��@�:�)��3��u��z� �-�h�fno��U��v{ܜ� ���[[���P+���A��t���<�s��$ �FW3�����=5��-�kx�2
k������#E��s7d{��Ȱv~�(��3x���a
N�Y�� X��n�f�U��6r2ѮD������{C��!9t�&�D��돠x\v�ֻh���X�HU!//������X���)�[ǟ͟���#w:*ذ��Ӻ�
�dY3Fа.�?*Ë�|V@9�:4�{�E*�n��x�/�e���� ~R��3�+���Hz�C�0�ǣ !��:�/~:$�A5�$K"e���Ԟ�2�2�5j���P&��ˀ��9�~�ׯ1X���a���M?!As�~�P%��ydˏ�~O^��C�r+�����4C�`�����+��>-L)�����B莈���
�0�w�G��n�u	(��f�k`������5��y�����\�'�0p��k�6�n�7y d_Iܶ��Jjk���c�i#�Y�9�t}��/�!���=*�1���}n6	VJ��f�mpH?eL���l�⑘=~��%7q
�p�m�>��f��U����6��Y!������.O�_���˿���?��gv'KŌt[�~�b�}8aRm���7Tg�N�[t|SL�m� :�cP}椞s�1�ʵ����5�|�M�xB�U9~!9��=��L�.�YІ ����Ɓ�"d��Рby!HC��o7�#�f��N��Y�$N^� <P'bǴo��%��>�C�2LzT���c���u���~��D�ri��ؐ��(C��>�� ��[+��Ll��s�l��)||q"�@)��̽�'V�d�9�Q�u�0�7u���D�X�]eF�n�t�������z	�i�t:�L��	l�3�S�.+]4,��g��C��4����m�/��ҝ@jP�P��O��o�:�֒ᠠty܇~ޣ�@���Ŕ��G���P�5��ܪ����W}V�ț���eɤM��)�]p1��ҡ�
*G ����U�<�/&�'��f_B�uț�œ�p(?�Q�sI��>�uឩ(J�<��ǌ����{o��t6�tEk��z-R���|JYk<N���$֗*�握7!��K������8o_:��t��O���� y?.�n��?�����wa�!؜��&,���Ai�� �?���_0�hhIY�_�ȯ0�r!*�!C���̈́��2!O?��m�"x#%�.ϩ�l7�Gק~@E���x`6��A�y˘������c��i�H�L��ا(V���+�Xt�1^n��V��]��b�I��Qc�߀8�uX�Ε��=�E�zړy�v�N�����`����/���[���@�b��-_f�X7������P�=[���XM��7J��h�g8����!�ˆR+�`ZJv�5D�S�m���N���B��h�pb�\"�116/M�F�/�h0z�뮅C<A��B�Xǫe���F�H�#b!��m�K���}��8�;�o�e�4����	=cHW�ΧX���I��A�JX�?�	@��XA.>H���9�����I��� /#),WaܣbG��w9���[�Rب��������o��>R��#���s�ݍޞ�R���G��YC}��B���L&�G�Rk�U�Y��UO��k
_��/�a���8�;�B�mh�{���4)y����_q5	���!ƌ�'h*/�� �PV�s~1���G$(~� �%��2�Sl�0�����vA�iM��*'��.��j��nS��!{���^,؝I����M��M^�'Zk�t����,~΄4h��&������
��Iv�$�����5>�d���#oJ�1�8�Kd �5�Z����x�č�c�e�NP.p�ڧ��h?�"��	O%�zQBU�QY��6�y{�g��u(��,y�{��@�c��[�ᣀ#�E΁���/�L4 �8��_��f4'��MJ�������Ug��IM�[���E1��}t'�� ybQP�5v1�m�S�9�P��C��[f��O_��z�^O��.==tW��VHk�"���A��t�A{H�0X�&z�����+]������&-���g����,O;e%�7��}��]����;ֈ�Z����$?�S��'�Gy��^�v=�|��^w�.8��wi�5Cm�?x	�|7�8�� �;=I���=���/��J��Fo��y����.tuc×No��!i�.�a4�D���a[+^�#�5�'9�ʓ'q"���b��ۼi�Z�խ[:��+�|rr���*.+�6<��Ǵ�D�/��x<ID�x��������X�z@_�x�R�;���h���&�����0�xL�. �K���	z�f���a�;*�(�}�����L:��_j�FIj�,�F�۷�G��anE�dR� ��g�D�VwC:�9�^&�g����H��U�r�(V);��:9*�R�[o����oT�@u������5�ؠ��}R�.��y'�Dٶ}�Z��6���M��ww۩��S�*��Z����1-�!7\�O�lzvu	���ޡ�"<8+;Nh�����9���h��-sǂF�{>�j^L��D�ކ8{�q�
�r�G�y�D�kgз6�� e�|6d����#�Ӄ��k�Ҡ���>�X�޼2���rt��ԫc�=�w 9H��.PU��b��(��?P�;�UT
���꽆'l)#�y�����n6Y�(�Tgߚ���6�?c� 
��X���+�,���nPq*�"���8��(hDQ"q��Zݑx1����+J�����1��`�[ԃ�[u]���¯y�}�۠���=���.�gy�0�um�yme�dz�B/w�Th0T`WOҸMՋ�E�ζ��_3��֜ UT#��~aQ�0K�]UO���,�Ê���X�KV*�}�s,z��#�����Bap����fP?+�ЧS�הY=�XY���Y�e�fA��tw��W�!ٝN�TiF�%�6��W�i֩=�>��[_;�*�VMQ}��78�+<2|["e&Y_߉�υ�����t��!0o��`
n���3Yh1a�)M���I���c(]ߵ�31�`�`�[��]��a�f��O�6t
I �;4�[	Lx^�\M�e$j���؋	�(���ْSE_ȯb} ��ݞ�������e;<�0�_���(��Z_%�	d�����]�^� �D<SD
�M����iz[�t�����?>�7ihҢF�[B�����wlo�E��2��.�\�B��Q�m���j�U�����T���/�ˬ)�6��v �ʞ�����ŷ/Y�*z+aQ(qYql�9�r/����M1RIs��x���SI�����p�a�W�������{��0�Ǘw��o7y((/�鞚[�L7?�W�]h�������㌵eѤ�E�/��&~LBm�[km����G�N��`�r�,nS�\����ү���ҩ���=��֙%��؛�fTV�(H��Jx�3D�0i��^��i��l���5F:Pv�>+§��1]��ܲQ�(Ƹ�!ܥ�q1_1�#�.E��VTBz��dLΣ�F�a@F���B�5����C\�r1��aP��O����ўm��&ˈ�2L�_`��T���O�O3��a�(�D���{�v��b9�Sq���S��2�0��3�c���ۍ$��Y� ���r?C����,����_F���
����;����)KA�����J�5�fxV��6f�L:�Mh��%*�