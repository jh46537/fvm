��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2˕@J��+���Qp}�ń�9�����k�ۖ&֬�%P��[-?�c���ƒ�GsQG��'��f�T�y(ԜX��;��0b]m�T��ID��l�J�H�'Zec�j�e�n�s^�
oWs���È��3�_\8s���$��#�า*]�\,���I�\��5���<v�*��0M8���e	+�%u�y��l�	}�sĥv�j>la���3G���[m���k��'CW����Q2��2��
'�d�x�j��C8��EL!'��@��U��N!	W~�Lɪ�@~-�	yM�L�;�IW"� ���U��4��M(�ѫ�G`�o��h���Ê. ؟,�%0�m�ܗ`Z!���.�>޹��ET(��;�J��̧�1ƭ�/��<j�4v�ʊfl��DJp�rf~
��G`#�H�ʅ&��*�İ�<Zd�am�R�^�aF���1SJzOKM��CM��]T�!�~6�E%赡�̑J����;m| �2G����$l��妑-�2(�c��$��˵��`���3��T�*�c��A�5ꊠ�Eg�Er�2�42 �;&�s��Y�f
;��8���$ߵQW�6pmN�i�"�|������$i �;�yB_Ֆ�ǈ�{�DE��\>-�)���jُ��n�@n�񎭂�,5q���5���hE78���	\	~��g����L���Z }�wZ�oy����~�{�ng�Ǖ�w'=6=w �5�ה8�biܬ{���bg)��A�$�Z.�޼]���/
��7̽���G�i'^LX�vXAyf84'$�V�D�D�ae9��#gn,yw����˟!-��<n��u�z$��p�"�MlV\�ϮM�K���O��S�NG�
D���Wf�~�\�d��+g( ukm�B|��AF����ɝz	�i�̪�V@�%<(*2�-m�qAj��C���~|%껛Fָk��,���[h#x&4-��uDS(6BX��U�jkiT��3Q�����(L���NS��㣏��H[��͜�c�� �Sw8ƾ�j�fB��x��u�I�9�¤��;�w�_̳�����Vc	\]>/�aJ1�n�#!Zd��F��>�
��'����x���Onk�_.���f��.ezz0t�2Z+3@M�v��4�9���SpD&ʲ��y��d Ю��������AS� �PWwezHW/=R����m�v�x�)H���9�'Bo$��R�[�����VQwQ����5)LP~q_���m�@H���6��t2��I�X �M�����Z`t' ���DT}o��;��\��ǟ,z|C7T(�x�^�n��[V�/R&��-��-}1-����Y�h�����~���4�
�����_�z'ι�L�	����܊���Q�R�.yO��6�P�=�F7��`<����4��A���>��)<1A��Rd-�m>ə��<\,C��y�@paܡ�2��5��)��h��Z%�+�Ue�{38f_�b�.ʬw ��y�X EJ�	ni��BI�J09��U���gS'�_7m1�c��<�逮���
�^{�����6D���*��E>@�H �g����@a�鼙�7j)�{� s@ ���҅^'�)Rڇ%�B��E�E
Տs{I*C~"w2�`���[`~b渱�'aK�L��/�E����W���R���b~�+D�'��~'�+����j�
�#��d�S�^�[�	�3��+�t�%Rt�=�T���hs�|��j�F��%:�k���"���'Aa�O\��e�a��5G"��OR*�mt�|���C�*� ���m�B۩��.�qm��s�"�p�\noxI�Y���[
r���D�bǆn_m,��`ff�s���$�9ؽ"M8��/EO���������"�t�H�8qk��/�!��I�S����te�� :�IA�*3f}9+N�9���ӹD�G-�Ȝ�*XdՉ�i~��b|���t<����Q�Ŧ�'�+�_m���[����	�1��[����	U	���B5�*���C\�w���L���{�2��</\3Dv���Ӳ�{��U����&5�����V*W�b��/6s�:�UH��߸?�f�,�6�g�A6���w"��$n��򶫅�:������NQi�)YQ)��+�:$�тҤ�ށm���n���5jU��^bj�Z�DiK��F��<���	����'Ʉ$ zZ��m+����#/j7�'��
)�%�V���j�<�r� θ UR�ʛı�_o��u�e�D�j-�6���<o�z|�,���+�%���RўUg���З1DT��%�����=�؇V��f[C��Tr��A;0�u�5W _}/\|>1kq��k_��m���ɯ�+�&r=n�bhRC�%0�8�\��,M�Glk)�Ȑ�
8fBs���+Al����ޅ��Ǟ�w�L��O�nn#G�	4���x�����<h�)�w'��^G�w�`˾�W�����(d�1����b�)ľ�)p9W٨`B`4ƈ��>m� f�` ���uk8cEC=�G�����J҄�ߴḁdrF���X�=ԃB����Ӻ�������SЩB=��	�I�*r�=�2�"���\p�@���#R_�Y�'S��d��`6��Ke��$��U�q΄�
3P������x(��/�Z�g�qu�O$�E+�ы�8&�E��5�KMmm�������j<k1>���=*���ξ��_#�p�@���R:O~�׃&H5�����M�=�X�W�u�â�n��:�?v�S��E��"�?�u�n[�M��W��I��-Y�as�t�
��M4�`��PO`+�"�uK�R���!��d�hE��C��ħ��>�)��mw{LOJ��°��Ew�l��"Y���M����%Aw�Ab�S����Fl3Vi�S���! s�~`PîG�V��i�]vl����nǬo�V�|�8r��nK��V�pl��	|�e=R�����=�Z���`AK��JZ�M�5۹.4TQ��]K��l|�3,�	�/�����g6I�=`���i�f��!RSUU����P.���{��_,V%]�Eɻ�%.�hPS�ƴ�Gb��WyiV�W�?DVw�1)Odۇ����e�q�P�GlX���U����ۦ��K��c����uQ@��}��|�w��J亅�6�G�H]�tZ��jG�^��s��\:{ϼ/��Q�X���%W-�;���\��g��ಀ�ѺbV���B�	�O�����ȱ�A��lʅ>����s��5Õȥ�����$a��c�y_�_��}�0����>�S.F���=��p�vF '�ulH����%s���]M��Tg����K1���V�"W��l�H����`kp�0d��YxQ ~R�Q6��q��a����Ģ�ҭ櫤�*A�r�cwM�&J�*�x)L�rݻ[�J�И{-�5N�*����+��p���R��2o�]ђ�W�椤3e���f߽�?��f�A�^�8�9du������d����ӦA2j߲���
{f /]L
Q��X������p�h[6�\�5tOҧ�-��K�ғ�y�cS����/���<��@�wV~P���a�}?�@�: ����V���K@���n�L�oQ��Ş�=�$3����_����_9e�i|�[#��Sc/��@C�&z���6��*�zv��|�*�܀�.v�:��@��ͦ��a�dغ��R�ʂB[q�v��������]0�9�e�.d[56�*W!'�2d{b`
�S!�i#���ԍ��(b��nlCc3-�Uy�{T�빁�Rq�Pg��Iy�u#o#��l�p9�
Ȓ(�����9e �M	�RjB��J��7���PO�%�[�A[j3b�x�R/΀� �� O�^Uw�n��7�@���{j�(�c}�5���+��>�)�X��{�/U�O��p�u�6��`��̍�En'�F�]��%�c�ϰ��q���y82M���e|Q��c���Z�E�A���M)�6r��Q�T��ə�.gZ�P�q:��`�g���*P�����LwJ��?wR��9?���%�otD_�A��y���U�p�Zv�>vM��䗤��ړ���+�\��P�	:aráu�\lU���G)���Be7h�,�1IA� ��v����E%\7���Z��,u���:��p��H�0��w�
��d��]�H��˝��;H(��D*����W��-.�^��R�T5a$���^���F�o����U(ؘ�0i���x��)�x�$]�Q9�vGgi;(�BW~������}�����,;A�y��sk�sK�<��|�i3l��6��R7�q����^����X�yETwvv��ى��� a��I��ʠMb}�a��9μ:D���%>o�2�i"c۔VD� v]�\q&�$q%��6<���Q9W�hS�Ꝣ��Lb[�[l]��)�yVU�TF��Ѧ��>��b�O��dV�Dw��SB�*��ñX�,�HA>t^�32Ƅ��zB��|�`�׺*��l*V�6����X#BKge
�i�an�i��W7v�	nY�?��o��."}p(L3TЦ|Cy�ۄ#�"���椴���9˷}L��f��.�%��͖���t+��D� �Ő(򁁳��N����-�ݱShC��:�V�EV��m�
]���6���.�l��4�U�K�R��/���K<���k�zIs�%�=���n�3����[1T��^������-L�E���V��e�hr����I�ו��:p��=/) J�Π	�|zTc"����;Л�W9�
$n<�Z>�N�5^��i����Aǆ�`��o�t�i�Z'̱[<�����F�W3�6[�A3Mf�N�k"�=��)Z8ݙ�ń�Pۅ��A\B���߶�(��Q���齫�6���W�*LҼ�ԹF1�$��;�3¶���'�d+������W��Ȳ����-wK�pA�m]�/*d�c@̶n�(�T��o�F�?�K��'�Ry���C"�SX�:���Ǚ�Ln�oC���Y����<N����~��}�nu��Y^G��/�"˂F�V/�@�~��]gr��\�h=�7����� ��@1������;Ӥ�уgk��q��࿧�|Zז��w�|^�ɴk��gَ6[6�b{�{]5{���~�Qb#�������8�zU��� w�j��\
Q.K��zhB�B�R`Q �,���n��D^�7�~/��_M${`�¢�<YTuG4�*�����?`01�Bt�gaҦ^{]�o���y[��/n�t�ޅG����#i�ޘ0�K66[UܮĽ��}8�ŕ�L
���V��MȦ� ��n��'�,*�u2�-U�Z��u(�|��W-�O��;�i�����jFԝ��q^=Mm��J/��!,3� ��kC'�'��`��>��m�d�z��s�{D��3 {f�@\B�n~���0M�"_���>'�͆�g�)K��wO: jJ�$���7���zd��^� �y["k�?+@�[�$o'$����T.A�Q�6!77�hV��_������\�k
�]�)�P <4�EĎ�2�@�R05[�Z<˒�䦳�$�Zq�-��v���<��lc����" x���K�?�!�g�y��G
�j��@v1C���'қ��z��÷E�#�BX�fuS����a�*����/W�x4��R�=12?D�J�Sє�	��+-��_g|�c�������E�ݬ��܅�]����*��\��֣+3u��:�������iъhB��Y;j�� �:\��ɫba.&ͯp+��xIlp'�� ^�ߑ�Q��|<k�m��Y��~
=(�0��ô�B*����]N����ZC59���	�&'2m�����DO��4���
��� ��A���"d �������R�1�Q�^��Z�l_�v�]��p�L��SkMP��/3�X�:�b�?R4M��<�w��ŏ�Q����@�E�_���3'IW����A�_Yj�t�'J���:zUZt�c߰����0c2�#>X��wƓc(�v�|�I$-����r|-���*���K����`@C�=x_Q�~�r�C���9�5wZ��_�Q�N��vS<�^X��	��V�_�mS� �I�٭�|inek�t1#E6׃U�Ŗ�CW!�qf W?#+R���H?��o<`�nr+z#Jhd0�k�n��_Vř0ꧺ�v�jv�����B��n�ܚ7�J�DY*3�,�9���8�ӂq ݓ@�k�|H�?Ȫcf�ꥍP�>��dd�@��R�����;�3���
�r� ��	��Y��Ų���H�1V�$�B]g�nf�'N�%���$�1X�`�6����9D24=}�M�(�������_1��]��la|p,����OLPu�D��kT��_:&NN�~���2�ħ��mg�c��9_p��'>�6���ˣ�$�M�t8�F������Ƃ�}[:�	e�]�M>����n���֛����Wt��c5˷���Ӌ�1�"�7�[i_vqېO��ި�t��[$׳C�}��1�ټC=��G$���~�<$��hO�|G��/��k�sԿ&���ϟ67wo?