// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U85b/x5gytqAyFF0UvO+brHiPGZ7wHiV3VtiLWle+AQwsI+NGE6l9oxumXrF34ZU
5Xd378Tcd9/SWH/pUs9myn/hDi/lcYnsFucb5u0RfyWTmUqZq8fD5U1kgk/ku3Wg
SQls5BMMnhfjR2nSG8dLtVRBSM/r63+BT4HYjMjssCg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12272)
l/FTNpiQbvBUkRtTIGUVjbWn/3cRvV+KiDDGP7uNS5QIB7zC/bwR7gMgph6dd4fQ
l8zRTZ9M2hwoqGoRGQOKlJkXr0cQIoVkz1bjavw6g+LbSDk9oPglERQ4NVXve3Eg
B7+15C/cMptZBqvXg+Vc4U174FNt28qGIhm5MDCyUqEOQdCVZT1nGMQhk5c2kCV0
b0nxKaPFugYenuYZQ1hZ/gCoH6VtLbq7vhmVhFJPWR3C5pAgsgJ42yyGvXwkqsG0
BKtayn6mHwNHk2wlI5/q2OsgHJoEHEOE/i1czlnUwyTnISDVvC8GMHxtszVJG7Dm
HB10KfxhSI01ctko7hJW+YGBjJyCD3avrtkj350AnfuOC+RgxrCLJNPpkTjUjRIM
FSa83hjKou6FX8qCMdAQZSChi7H4ENCc9REB8a89Sb7OU1anzbaKFrPB1eMhvBtU
72mhCDH4aLJvfgndCmNxe1+Lbwr1AF8YoIsg9Ac1kjbnwkPodCgV259i1jVB5C4a
YvjRFb39nbOWRbaE2MfhbPyAlBxEKCVRM3U4MbxTrGERYJaOES4G4Ygoz1XhmHmI
vBx3rKkDYOhMbnWOeNt16EdQK1h45X88y154uYk8EoqDYnL3VYNnli3Yy+qiqAjF
ACmRDrIzV6UcNDT626qbTJpLkc1RkItQgJopk3v5or+TyzRjSTG0miPT6bzX1YOM
OQxFVU4sGmLULK5xtOVzLG+ke1Q+7Vs8PkLc9huAW6jp1WsCjuSVXPnJXxEeno5d
nXps/OP3YpbVVUWI8MpJcoMTJBVcob7DcOj4j1BVJl5K6WcU/c5LKAvHb4jqfYUk
ljQhSHB4z0mJg7iyjWXkNdkJeIHn39MZR05iW22fULRqEna1nhtIJFSmPjNW8PrI
NIlsIkg7sU3HTD5C/DRIf5Uwirrq8+7oW2efgRiOARKJd7/uvXnSevr9Ms5op3Fc
fPA6NYR+m8kt0TP57kKNEWUWmWIr61CDu87srfTa0LRL8ybN1EZWum56htFxw7sn
bRak3rSHCz/0ao17430whK4/ThVyJm9P8J1z+15tWvpov/luat5JSBSoo5dAxjCj
3eUahZQolHW9tKyuG7Dbqy+dhrScKOJEqHyvjv+2I8WDb4qZvg2MFA521B6a5uY9
rR74cT35LwmFk71q9Cc0j1iLqL7fiORr4BCVPEepyGwZA87YiQ+85r8tUD6Bl6W3
O36/13IBJj48rOLfnzSt0/as0KfJ4um/H3vIp9B47+8JPE7/MvYMKgipyweo/9bQ
Yif3vKwFcxypgLXpctCaOUBhdyznYds5mCz7owLw8ENniP3T1FdMfOoXZyg3DZ1z
0ra3aRGgTWLbpr7Ks2H9jAQmQIPFAAhNT3zlxzYtDrrN+Hdxj5VGYSYjwMEVPlVQ
rdsGv0r65DI1HzhgTKG7MbGztGzbXIP873NfhKdR1JOXQYy7obP8/VNzrnNicLc9
xZ5Y5ZpMULf7kJ6EHPbwx4kfU/R5ebuFi93sg0yYlB7MBri2DjM6YAvGEeZ/l0SU
FCzwL1jTlfVDkVZy+qTYk6IrwS4Z1ApqhKBKwJuFuaJ9i1i4DgInLhZ/PEqrQjCo
Ou8BA8OtIyr4MNv01ggF0jyHBr1LFz/8+H8BFhhoUiqlb2G+aYe+P/Y+9mMiJS03
TDr4TfgukrqEIwRPnkCao+l8PGiSqgtdziuv9amLe67i7oXQiZHJnJ5u2tl841wb
TlY4v0+4OEdUGbFSK3p6wdcftsEa22Q/wG0l4smnZu/Al3wuhQ83jZkh3fW4Iw1B
oBqkMzJTQGewZHHaN4tDG+qymCtObiicJlmamYXSM+Rmu96UFLeX6Cp3U8we5+vU
He9jvhaE84WjLRbdmDAHAi7XCMj6CC8xNfIaS8IwjOWL7EVPGEK/TBcFG3XhhxEg
Az5zLraRTyOyRie2ZBpSOrGNWRnQeuIN1CWUJFrxcscoTqcnvV6Hulem+ljZrHad
Lq3uszx9VKYVH+NJ2zhlEXUKVJ4GnJ8RAFr/HD0Td2Tmfu/4x3Ghq9OWVKrVgXi1
Qat75BA0iqIjbxmWxEVfhdX3XnhUCZ411fF6O6Yk6+yDL05J3wTv2NTBNAP8otjS
jy8KtFssd0/+LJcy8KhJms9SfN1pHfVO6AfJWddhWg61p/LN5TfTfN2pgfWKs6lt
7xxQv9NMyccmxvDq9HsL26nEmXpCvbTykLzTZgjXhUPRmO913EVJq4cCn+lG4Qvj
BuTxwjqJ0zSy40XOa0qTpEFidYKCvC48vVBiqtfF4YyG50SC1LcbboaXtEjNDp/k
NigrDI6/YwWpa+f8SvpXdFYHtiGnil0FH/CGpJlhSSqaiUonM/+rNWbQhpUBFtMf
AF3uJbhcQvrerIPsxI9TGXiXticP+NtoBRDzDjJWgMBnRw0wMhNE9DV2xXJeQvj5
LdTAeUlBR1Y20+MdFo+cdm1KrgBkjhAwuRewIKEsi8ibcOlNGHkAwxxdODz7+rkE
6qzhmsEABd49OWUeZ366wlHuoUK03jqs2dB2x0K1dtAGqT5KbHIaihe+gMlwDlvl
edCZxhdEOyKRElDWB6JWj9rqYTidC3FtoO33XbE2sQzshjp7YPGZZ4hkomxupaF+
LVVdlo26LLCFb1Bvil7bhQOoKXoWrMM6CkmJ0y+v5zVAyGhLf8KLz/CqT/+++zEY
1keLLn+IddgNcDvYMAXwnn7A4cIbZHNmLVvmtwsL37uAhLKAG9weOfJBPk7Q8Svj
VZLYlZnEtr1TnAmiLrNaT7/+8HIWnEfdxSrAtcObH15o+SlhPQwslL5FU9ndgees
y40sXg8CNCkHeIMHMZ9zyzBK7/zhuq6uj4lP9YSlYV2D7+Mi3oiydMjJvo9lzqra
NZrNCnXNAQCepkW30QtD4LRoQ64PWjiOXg7t4Vsvu/3vEhg2TVU+fYOYlgJKSd9U
+LC9AfpLjdXzOSD17bk1+eGgS0R+j+VWQ3cRoxYi4b4APeCpl2Z+175Qq4upTpQk
ZpJTea2fxxlBH4+j8wQvGxY+oHmb8naH7wP3NcxZBvudd9/pnvZhRgn55yCF2+1k
u7XHy9jmConbSr9pT3cxP6EVTtAYD1Caxy2DxnI1NxODeNjkvSw6CtVL+c1XdqBr
nNmkzmdPEkZ0wPemRqtgiXq/kEGiGEAOFHrb1cCFXPhQvQ8Kp93wSgQLbHiXj8H6
UuTuCAfjdLLB9TgdFt0lfInUnxf0RmQBsjNffdS51vIusqJI4kvfiCI7SNiDITW4
/SlB5PLjzRV5aYYPFTyNYqewUkLBOrhiq1AwbC5c8KOIvbvxZawLwdGbUIiDiOtW
8iKmuwmaMB/nAQoKwDrpmjreDrx4EZsUDn3YKi6uvIKAsd0qr3JsThctnVd8ZK+7
5ewCwgjJZwcGSjvo7GQWOfGKGkyWM16GSWROF/HWxTEGwdEJiD95r5PekS5nQWRU
y2z5PG6guKX3dujEibSJHHtUmj9Purj7iUrlhq2SipIFJnmoGqb7YZxiFwPiRuNH
3UvdVJtjFZBvl9z8DR2v5QSfRsvUKxW1WvNjrmjCHiJ7puEVu9i6a7UWC5WBAGhO
wMs9vHUgsrxAmgrvZ93OjqS4hYGyoM8NYMiJ+3nduC9e81n/HP4ur8Ra9qDLf9tn
xb9WUwLTbWyBr5773GZGlM0BeL1cHnAsBgV0wVMvh2ebOYT2kSP98UlDSBbvhX0y
4fTlq9iOSQYzNor8ZhI4NcxD4YL6UWh9/qQM9JNgKdYu7ZZiMpDpgpmbpBrIV68O
2xViaEkXIsSh2B9wA+u4IaolfnkTCvRF/FyT+ndpsiRnq0fqUwtat/8D83ZZa4GC
BkwiZ/R8WY8bYO2fzAIS/zJykZHa7wUNPeouwIl62seUwU5i913mzwMLmnmr3wUI
ksmGAiagK2sOKhyfzFVz4JDax4EVcSfpQHnTQTdF+2Hk0DMsYC2waaifLNVr/bLF
OlulEYzpZWN0bqmrpeu2ZQ9MkwHZJPQCaeTJgSgKTLOxdG8Dah1G+eOqMiFxlEvU
ahQzEHT3zjmwK0b7dU959F5dRQCAhd8hG9dKlbg8wC6tgUt+1przwx1hP2+qN7Z6
ppPeTLsoGdTJjYu2eKBXhq0kaTHL76VMXBN6y2EXWWPHlDOpOlu71FfN/d8qKDaa
raHNDqCsz1ZTPjHr3qFL7eYR8BjXhtPI/ZogDQqz+plDMi51r2M+KrTHKa7Sn4mG
LY4mM6ooEZ52+q5sH/WrIjJMnmHZ46HyQL19Ju6utu2kKtVHIFMn9r5vMT7kLbnu
GNRwWdDi6R3e/2pev8Yj6hbQw3Hnq/MK5wuTwQIDeDTtAsbWRa5RQX/UXBxZ3uGq
Zhlb90ULCeP3Hwvk6xDMoYXHvFh6iZp8Q99UwhjYj/AKif+Bz/qr0B11y5zlTuJ5
yzQpSH5MK4ik4Gah4RAwkm4zFdv++cKq+4J1KSNy3dJgFd8yM0tX9QrkWcuFoiS/
UkJkhsC6dUo/HdyoxVHm79MMp6+uG1AN1IK1PfwV59lsYPKd+GTjZ2nZaD30Nrp5
qn9as+qaza6+GCatnpvtAQxyIUSwz17CTidx9poN0GQpLlPn8VqISKyk2s/kXUH2
6b1f/2i071Po75b78XSCN2SFrjA/peXJl3BmEA1Nz4oP912JeJQD5BLAyvd2cLiT
FsH2wgFfa8B0DidTO/l6SKsV8w5Ao2IN6owXkmAat1i/Yzo4GT1qXMcA34psmFZV
OBBkxW7dG1yqZoY0TWBjvsBJ+fSkx82AeJOpcAIN+9fN1z5GxBWFJkhMfrEha7Yi
BrY4OTxfdwLLieJjIDm0IVUkz5hp4dFmSwcU4x81fr6jL+t0b2ZUMNIqTN5SSYaL
/w388rV7Z8AjapwZN35elUUKgwh3QaRUTqlCj2BDV4K6uFeqjvtx7nDkiCDgD2HF
jYJkdLxKnS8EsuAUxp2bzPYjpiMArFu/png2gHr2xfsy6OKJVgfkYL2xTVv7bYTw
NPFQyyDb5OQ/bXCxiMwjXITNbuLH6ET9MxzIqTcxKhRGSiJWRU1WhBNNoi1oDUOE
Qf+FiRx4noVV0gEnC+TOc/dO4lwN/p0ta95dxptTQalOFJGIIf8HL03JpcUzNKf8
+76p/HPXMjFGOPFrbucLjksvKLD6k2VKjZyuV2Gs8Z5GpIZ0B3EFCGSLqxas2aPR
pInca+dSIuc3SFXB+VI9w/zql6uecxo0zAClwUeYZx9Vf6aIPAzjjSbxLS0+EsVJ
eE+Zy4v0R+2Q3+HQr3RniD/g0INZWQT8AWK/nUze1rwhDpDo1es/PClrdgMAsjfE
OBHQStUSwSwu0MgG41IfijhPrAO6j6OGTQEpCsk3Uqfpddza+9/SzqoBEZgLZ+WM
4EmrAHPvcRB1dLkkt7eGBdrsL5f6C+7TAUJR1EdYXd94YGH5ZCOQcl6YSQDQGYkA
/7tC+TcFG8ylpKpFS6ccNAyKqqD0qMZVcNrXnQHuywcOYhZnpbfMMWTdtaLQ2emh
D3PYJRh8BO2blGo6aNY+rJ2yJkrRFupLDvZ5QUucsXs9YokCji1cWSmVVV0pOdAR
wdXQPHxo8+5wp//K7oAwmaGol/ejK95Sqa7GtZ9+WG5MBI/nofGKCvHUJLPQCpXJ
X1h7sHJUFAjUK6rMdx+gmDPlhkzE3aweMdcdu90hr/pyddu3VqbHyaCqBucGk76u
AMXiH38YwtW3311gRHZ5XgegyVvxLdoirEbzoH9rZbUvY09jDKFQW+N7aLWmBQzI
kU0K9nPJBkzPQvYx/2WHfyp6FxN9q+A54gPwcczJZpscnBoBtC+pu6JkI23xTbok
ErfWEIfcf7EjKgmqm0JKBKGNea/BsF3O1QeW7/Gh6JX0uo75UEnGw/n8C4UOmW3k
RdNjjapQPn4+rJrtNnLG3RWF9wQXb+KJzXFsTIVOCxvdSRcFjyY66KD0ESHtLX6G
T54EadN0FDXhWKc2nd7Jhk96SfC42HdQQJXtU6gwvbXumvdoOv6OZEpYMtH1qgg0
e1/AAtPbWPAHCfy1n3m4w3+7ATOVgOK6GBWrMxyx+LDWYzpe9XFqknd+/N9Bpd1L
0Mt3rhLlZO40hKqRgqeJqTluDwmef5Q+nW8vbGu+X9JyW9XDcH9lCPIm9aiKpZYl
vHinSKqJyo79aEmnE2ydY7FzEbPX+rL/c0J6+y4uoXkTWO0sXbwuB3ShckZ0czRO
o9IMVo4I+/EjnzPX58HEGQJnBC8yK3jrVuokM3/JDqfZS1SOwhZH2zPyZQZMEZ8g
IYhhJ0rrxPNPn/ocn3HplVxu8yJSouxsmUIBwhB9bodle9MC8sAwblArjYb/4r20
B7gA6wfw246gLYCIDemFkbuPlkKz95A6B4vS+CGkEXPHzsyJihgfUZVHPsWDivjK
nM3vM4cT0g2/GrWBURsiTJ/x1uwQWPoZUrmNayqtiUT2zIe4RmzBh+Bj5K8v0WL9
iKIDzDfBCEDzutPBf3YFpWMm54n3Fjsry3PjK2hDIof5vdEThPKwrHVEHYhSd1/4
OLai7Rq5Hg1ssgdTiSD4wVcaK5YGcCfPr69uj48Eb/gUmyBu/2IF8ZgD0pbyr1Cv
f2Leu5NTHVKO3EW+pw1hUgrb22D4Qn+UDYJtAbKPVwJPN2AsxilxT11xABxduKZX
y6kEimoXwtcDf+J4tbd9I82uEPo6ie2c1q7/f7gcmyvLn0mI0M2J2W20/nq3ug7V
MwYNFbQe7OGwxGblsNR7H0iVzh62MVbruaQE8tQfEmyzk0HwS2P4SU+LnhEmNX1W
9Btm9v79DsFGKASi/LFPnsGoh4dRSMYRed8tdn99HXkiDwxkx2D/94Bhyx5tYD9S
CP67daSu4vVoFbFMahHIWWPQFp3yUqf6ymtV2nje4pmrktfRYL/1kLILPRd8GOSQ
kMimW+fVcg+PsZUHXTdOFzNHw5ZxMSOSPm96QAnc5m18U8ciqt3BIjI+N9gAvQFO
AsKuKIGC1p5SPon2m09aoGoGBzhTW2aEdIBmWZwphsAPe2Yy2CFsyYHwjw3cm/71
VBXhfwdmZZ+3Kr1QT0TNzsZvUAB1fAlCAkyHNjXighNhpgPps1lKEr18JKLB0veo
TZYlwDajs86KxTOtm0abHRozhBTRiiv9eMQesSdKPGZD105Q8RgSZST9+bRVg9mO
Jk1qU2Tdv+xBgUwxbG1b/o43dQL90s4OoznBR3iorbeTtzWXTqdqiE5+iovTQAbl
t5UWXsRYzSIzzlAwYAtT5wR/Wj6TAUpExErctEIAii/fMF8CjS6kqFR+AnbaiUml
mYsOKKJy1MKSrM2J6q0s9EcZgyU6haKvzVsjABYZOCxE51dlLmMfFuN82YTqW/zA
Zy3k+2/XkZUNPHUkdR+AqjRBDkk+Fvf3LVPXfAweElnEUtmGE3QPIallEt9aQQF1
YS11kgEAu864Xa/yjyu5vc11ZRwUC86zlwCOdnAmzcAKYVsmDFrqP7EhuiW5IAZz
eVFIadyMnsmZnv0QB1vRqaGxavqQXi4mxf6FjKrnpu6PngiIXW6lq+FAHlO65M3x
+e+8NbmJa4YxDw3NY6NOOz26EBrF74iM4Kc3cTBoLCEhPoOXFxW7IqKMztuNGytr
Z43qhMgvdSP7kAtyqQTRr81jha5pG/zsgSAb4QP0/cxaA2rejfXd4QW8LbjzVuRJ
kkTgctxX97gFmAmEBHPjP/fEHdcJLtBkGfSrD+vacHgD5n4eAvEdOy1X+gBR1YaV
COhoDfa9VKme0kG2VbjnooBgJwlhGKbf4g1CpAUQ+akJxx6E3aQp2A0Ntg2Ch19b
aFOAM/i8GzXHo2shJXVQgTM9SOttPPqVn62AFTmbxvH/3goPVerhERuxe2fT1Uic
8gEseBjWm5IqBcrGKdDP3kUmcTefFVybnQLEWng/swbiCm+LPd09cn0YFy2LFuuH
dxm+Od9tqYYYmUPRV/0N7qbMQxLD0GGX00eRQT8q7V0iS84ADyQe6ujeUb1f7Ail
2pnDjIr8p8E+rMoMB4gPn1p1uagqrgm0sMWPSmlLUi+IFlOZfYaiwmi2mk1k8ZU0
RksOLOkYclRhmZNNKpQXg90F4RyL84sM2KZbVnT3rzNVg2fSgZjU1EXOiiFDT/PF
a4jK3eQykEuD5K6GnwL1UWZga5MTxheMqRp7k3DPeFz2pMEaJ4ilYlEHmBft/PRS
zL4d/Orq/CYl+PikbhWXsdz4hjNe2od3umL8SIF5YR5pbvBaRWxpsjhDrozhKGjy
51zItNfJh36Go/ar6v9O8CBF8YSjAH9kQGO9/oEARV8z0MsJLylUetauwtxAZL5o
Po5H2UVae6XvjN3EoStV6gr/AiuihLzuKDSQLFGRkk2aLSnQUpW0DJQvQLVRoRIw
2shXVofF7O1veIOUFQ2xHt3Ryw2IglhI6zV2G36+ccTlAqbeL4htGxj8Q9UIAoGA
7BsWO3IrqG01OGlGZSgpGngs3O7EfjZFWoHRcu/YcUQhLdE5UNjbj6DF1ADZKnPU
WcIXAq8WVS5LmTEL+LxbeZYYZlpnjVjSAWWM3w4HXBO4XdG+7a41StNoAyYtPVij
cHlGi4QfElLTuZzEyR7yV3Ekm5JU6NFyldvDdfRs0prl5XQwRQ0ZieT5gjc5c+9e
MoMssA+4a5kd/zvodkhmlj3DDEaLLmIl7yFh5p8gTt0jxHmrHpCP8XIne44Gb3pL
Oi4TE8a+oRnvDFT7VJTCmX+PZil0LoQ87gKA1COS64vis8T16ToPDTF+O5G87dIj
WSNGnRTCy8Tc6nkjsHQVCrhQFx1lQFGFshzuuq8pT1vyAWt7IiAcKYUpGDxtjwvK
0BMu08K96YEiuI0yOo5cVvt/AHa2bPDE/8pVXdZCF+Qb0Av4upevAIcEC+MHIgG0
wErH3QHAARfbBFNzk9w6rosvkpyNfsSYCQaeaPBr/gc9yi4RTs5MJKsQyKHNRfCd
idBCBfVzFI5LkKYvwIH+ccwbmol/KnWskG6idBhvIQqglKdHy5sfFUbjK/pe7jum
9U144JaaoYAlRNmsQ3TCBn8kt2NuN2Iwrunna3KOAq7R5jToZa5rfJFggfYCc8EY
TVa/DGBqfX0VOMl6WWF9i5L/gOeygNHZhNjA6nAaV8pSP9SvNVtau6tKh0L05Hcq
KMyjT+C7Z4fCx0WuUcb0CE9SnhlllFmSUcil9HapVArUM/M5dS2pKnFbceMYTCcr
HAGRO4mtvJWPFbggaxBZmiHST3JDkmjRm/9AGsvhRxByRbDjWvz75G/46XbRQ6iC
E20ABTeiJfmnIagHJtThkPf1bGB2matbAfG82AO8PH4dOQc1JAvgRG1Hb6r22gQI
vLEqxirxgboAXNVB3oKLeQGUn3puuAmIdUcjhK1w6/FHn8pPtFHi2jJUtekYOHFC
9xUeXORA5E0vG3/U+gMpfNPi1M3OBEI3o3MAigen12wWV6pH+ddF3wZE6Fhrfgqw
ahOkTtR4zEuvCkjppdhiDVkUcrt7SuXDzU4Kv4jdYc5ZYQP6hgywi/xJUuColDuO
htNeew3OcEXYMotWzUSZ8htpsCsnfgSKkheVUTuYevLfBH0+yn272Eth7VjQwRtT
Wb5N/lMSh/WAcyLMiBCUtKqBN/e5Y3fYrCzgs8J1QWUDme2kIbQL32lwVJBJY0Gm
qmBNHDk1UyNeEcSJK2AO/mA6CsvLiJLvfpJT1iO2J0JwHxLMvQb8C7MFvPQrRjNp
Wmw01P68ZPTyDQxX4lse/aWf/3HRG3FQAWAIZkJLHR9sn8D1TipEfiC9qQm+GhqO
ZRvbPufNk5fzyJ+7qdVPFOvkexcpSnyNEzUqiGgP9S5rCMnCB5FEhSjStlMUC/DC
fBtscUc/+cBBS539p60tLvbi47oJOC/Pzsf9znpJJHNppCFzr2+9Tvf2g7mTOoiT
EDZvTDex6ZQzmAssCbIOYzOP6ip7D9NxQwJabR01nQfqzLve+E3NzIhHgl3XDo5W
2MoK8QA6zRK9C+bYy3LLeXlb4BlJVuZzH7sd277PqSAT1SkfvS5+ZuWJlQNe/JYn
EmJqWCANfDoEbg15cZ1R/CaPn59DC+G+VpguztVJVx0NN3UVO/FzUx9Sr7rFIRRy
/8MPrDAeU0HTsNQqnySirf/KbcDZso7O/irGq1jxxgbt+cyin16u9bOgg2IfFGAU
lNnhE+HBfDoAhjKxvpP6DQbUqct12vd5w13S4QDYHQMPBk62e+PkZfQyydnCKKaL
zzwVhDVtfTAPLnjpHKiGMCBmkFYpheIcJ/s7PRorXTW9bT8Aql6NHch1tUydpO6Z
QhvQ9ZX5a1qItv5sE5Y/6KYBBQyHojDQDUScepkxSIsDKdw8IXFmaoy4hVxIdXbZ
KpEtSB2UKlX0FEo16WlX3YfMK/rBMxmsjnFgh9QjNFFOhWyrfEzZNzOKacXYsRZh
zI9jVN4ZMXigIYgoq4xscCzAhxGE1w3yXfzO5rmYZVu2coTNyAa3aAGCV6YFqtz7
N5x9dXxjF7OncdpqeIqc4kQjGUipCA4vME26Cy2EiGhA9M3nBGJpGS5BDJkVTcRv
ShB4r7yEKUHxxpubQJNYxC0bXVOWMd6BQ6VckJicAzcZDUIG/9hqucj96NcrtyJB
n49PIYceG1+bib44/Nz1uKArAWf+FuuFSq05dAVBr5BmPWU6e+XJuPXcPsuspWWE
I/k+iFo/lFrOOfDXHuuS50+3Y7pMDGM1r2Te1C1MANzfVolV86QpDNr6bosXlc10
WMtwwRUcFU63czMVPuxkTuYXmQn7ftqrh3MXdr8/ERfmwKWYd2ZBHNLTCeHofcRn
Ka/x6DwI4mtt1o5Ay6MzyWel/Wp7X/pSYqv0Nf8KRmq9CAJLGd1xe/3mUZj2E4pf
nwzSHS+IXaWz0zyNtm4FyfQxTgvAHZMJuux5FqNQ9vBel0kcOqoRXmTZyaCywwcc
g8LDXGFMMYDzCv8P2EgxWgQwp/QcY/+v9PHvgtJC8s7u1ZbLJ60Jex8O0yvBuDlr
lfvTTtQ17YQafkfba1PlB/9Ird6kcBDNOpylVRa6Liz9V/KiFTRUr3KQtFEVGdX3
5vix2fXazaGh0gtfeJfZx6oyaKJeExiYsQtiI/rnZ7Ar1qEn555CsLTGmAfc7uKJ
aSuEtJQR8+1K/iv0UudSpUncwJanNZ/hePBGTiIONyuUU7QNply3DshTj22VPlEv
xfyeNZ2g96dSMT0dcVP9ZfGZ0yIubcO4MKXR4ZvU8jfEmu1S1MNHRSqyKLAMREBZ
OrGAmDYz2Cmt0xR8Sy0bYeyIzsW0m3rBpdCD3Og8eTqAekr9/hC9QkUxjoSomFKH
MmEiexJLVIljcszQCSWPJwCfUV0ssG5Q4c+2VkmaQ4An2+k9Diw7yhMSayGUshWu
puYrvFIAvc2kAqJdRv6tE5V11kn4YNhek7iMNSweWGV+u+qL5Wreu1tvgkiOpTcx
eKaZ7jlaZdrExOVxD7E6kTU0KsHU3PYuWuUnQQluGZe+gRqANZ24yrEvE+XXXUue
Eg5W1RKLU0n3+ROeISOMjz1r2Y6p/Zo4q9NJH+flaYBkE+BpxPobnLAHo1b2WHHf
2E+zUGIYQ3uRJ//6gwTZ4v0PIJcVVyb4QaPft+Di3AgV2P6R/c5lM4QhJ+TRTT8t
CH+YA72EGLArZG1arFHyxTIzrztFkr925AofGA0pRpQz453zRUQJP9mvILaHJPbG
ifwwt4Ec+Yldw4+Cena3kZBWEBPVMGXJQcGddkZme3KqCLBNVl5sgjYK5rIhfeS3
4PEBI8CtGemLczZ81R3e2eLRFKN1ZhhmRvRn9gCfAhg8bR/i8R8qA5mmF72E3cF/
hXHmsfQBjfRC2Q/V7ROdfqJuiZXQgIPviRzOr0c0MhCYFoAZLvTqSJ+77v+l+gJT
EOZ91sYEHAOJkGJupDunm8hgNrDy0ds4qMm4oXDzKyIFId22HoLZ8Tcsl53irpn6
nvt0zcBj+kcDKzEG9Y4aRL0IO0dyBKdHa2x4g19laNmZmBCGrkkAOU1b/B0LhMDO
YNQGG7SQKomiOHl0JKD9ZoU9NTdTPYX8ERT/zl2CsrmSKNa75nhaJvMd5By/E76l
TT08iAVvU5YJy1QqeWbMR77AW1wJflRuqjwZstz1SnHFMYsfar/XLc0Fp9Qq1Y9V
MKxMEMoRjqjtUu7zpHkdV6KoQnGVkb5Zi0Z+cf/DfnA+X2qJRFriya0GuTMQeSAi
CKGJwQUb2ZquX/mVQn0g8b7wy0mNXVJKa2pMSGtOOa6zawlSDUYMltVTk/xt1sO4
ao4VK+kjU80D4L2GpzgW4uZLrS+1bhcHHChyiWV1oPWgcvbWoTs/NqY+tH65lHAf
SxcpN4fgOHACZEfQwoW6+ybfK7WJCkhIQUWghFMYM3zntC01R7WStgOgEDGpKdqt
uqXNoCpjl6YhO9Uw18x1Qe2TVPkqLpl+F2RtFNQd4+jEBD1kegmmcoasYZv/8kLk
iNzRZti+s3teZPjyJ6f0n+NUCidfSqbCS0BuQBUpdlibFxoTpsCPAREsG63UdS+p
SysMxC3D7tk+pUjbQTzWX44unbUmTYszgeXnZDZ9BGKVLoRcf2X744e+D/CnbE0g
JzJa5CRyLkdTQxO3v8zEVUZZuIHBbBS/XL16N8LbX3s8aZ8hmxitNcUyvYgAltOI
NcG80JNbdD/4N82FcV1YsCpv4EG6ecmj1blcDtCepwcI9o0rK0YqOaOJNrhLLS1c
h7lLJN2Oyb+I4cjZST/BYMHoP0q+a70PDgq4czkt7KtGgh7mBb+jh84TlQby/sWQ
KlTNMmeXrmeebaD/ONv5pc1xypw9mHEkWibhJNEi/Ur21zeBH/HGWCTz00b35eNC
GZURlhLROmnRc8gGeyYt6N8KNrxwE/0z9nZNm3JcZAIASIzyweVHUY14ZCNYMipx
94RitM8zjsp/CKKwSFoTicfcYfVjYvZCWUACr3xGptxMkPx6aUO/HUaa0tqt6GaW
kk+GocrsBBxBphZjigveRxOQfbXGDHB1iy77i1VDADugm7WXehx44pmxkZohCNTR
MNHIUVZKSEeB3I6gfM4uAm0kYNYxnIEmR9CZOkraHopfTAHJMhvRVNCFmKasKUNc
cy+efYH5b+5sz4x5rYxkE7qp7LsY7aNqbe6ShmcKdn5d4bUHWg04mW5qkAPjKJZx
HdyQ8vNxCE1Mx6hlFS7B+KdhXTpHS9QnymdFPGOdphtmjYH2xwQazwn1ZqcYtIUq
P3muJbU0eSWX9+Bc0orNiEpDbTi/Uue4k1pskNXAWUpTO0uJJp2KuMs5DObGvzx0
B6jd0M4wCu91wlMqQgtM00UGUYBkT9CUI7a6UgSDhnEdHOUlzm4EvMY1UDmK/ns7
TFJdyrqKTnmfbZPmncbYVyJny115vIs+5D+L1KWJ1ujaNuN1xWZEssauVuHB1Y1I
uN1517NM6gM2kOQcvKspl+aosb4+0x3IQSKkuV3+m1ZqPjtY0jQ4n/4bd1DaI+ix
oErQwyXLy0difuyz2IyBeDUEG1woPLwgdLeIzhbsKk/9/8Icck923SF3PmR3Yx/Q
Lst9eylqqSH5V2MHdqIMABvIayZDQvWeh+7dZjN4OncfaeuhTHFLlt8lDQ8wwxYh
24f6hVJwcrMJUW63qZIBeIKZRmND/JxPpHURWpAeS/jYG/HICzg8tUoSc9nZensH
tJf/aygM4y7V6WzkWM4j82cubwrtiy4Plr9nb65FlhZHf4Ylxw1PEK4RwNHZU9ln
NdU18NVD/jN9FYYaJpxyLpcdqOksQthLQZ+EHh69SSx0PXhqye3CXzcSsfQL5No+
Iw5uK9VPmR16WzfQpusGMCo9oIAaXMrfo/UyZoGryZTeBT/f+oe0e5ZH4h6dI5gS
g7o6hg/ONQqHUoa8lKg5pcj0w9tN8qGzgURArq+c6iD7TLmZbSlCb3vc5xp9sD30
dnF+lNxSFzosRazU/dTZeoPZ4vNP3GKvCV39QyCC/lKNp2NjAESnCTU9c/hyyve8
nsYZd4uZMbZtJbCCpbJtGnI+Eys7V83oiLWFXNmksoHJIMBMthWoIRwyLLCBylne
dQhKqDcd2z8uL4SSisjwIko2h3oTnVDjBfWOFttdZpLxOzvc6qGMqesW8XIi0h97
Ucx6tj0BqveFdxUYkenLupru2qohm9T9izeDQaXsY8zsjResd8TXjNoCrd5GCxUv
BmmdqBNxq4EMRG5Ka4/tNelQvzBtqAsITCPhnICqY7EaoXSpvokgNv8LUAFSP+tZ
K6F7CDUnG3UOzH08AhgWN3UwQuah4Q8Ii+nLtPvSk+V7Wnok0nmjdxCMAZkT+S9x
4BBW65cqjRq381tRrQqemAr3V8pXX5kwbYNbANVABl0iEEWlmL880XpEtgUd4dUg
5J6T6Dl5M7SfPwejJZzf9AorReo57TvraRQb/+wOTvOjlmXo/toiWNKuO3iSrQwb
sQ4fcfMuzBidCto00Y3TKkK9zrtqg+qdNUjM2iLS6rTlix114mEJAuc8Hk+z3Mn9
uTccS8A0/3LDuDPHFIbQuBTUnoDZgtAya8se+GJT1wjccJ/Nkegh7MV+uv3Bcra7
rKUJmEIbFri5qQJIWNdDizPW/2NpeOxGg+NczERkv9f3Gtx8IQnnR1m8VmihsxaO
V/WYaJYAQxnyh3th51ucBl2omKSAYp8DNtyM4BL6QqwSMHV4OKFB8hb2I0IysnHv
7K9KqsqEso5c6TQ5/6NHn7YacqtiTpnyVtBHwfZs7HG6nOb47CCYRWNzN4s3cOYR
z43oJ5KmUO6Wagwz89PEwpXIl75/ojOgKLBhPAIISMoBngnPpFUqVV9tkmhrusRG
4V51RBKrBYhXKutUaBBYLZ/C4Hwg933xgaTaAbk4xn3OAfK3YCyFNeWmuLrdyGqY
FbBBHtFbPGInegU4SrmGBNNpE7XMkZHz3W0r+gEsVPViyDpgJe4jS1w5yHzwao5j
4Dnvk/RjqM0AHRSuUy5RlK3cVOW3gCWw/lKjcuyZCdfAtdLOsOaj8mLdihqWdUE7
8r/a/0VeJBNlZLynRAnRjPzdoLtk/QA890itVSoI0XKRSi6+8BorvX+Hd39K5DUi
yIxn065v2Yn2n+edlOZc06onL0qCQZRiQgUTOuWD2iUMlIkq1R4fLITcId1EyS/a
5fr1/QzBpqo75jAtlO5ZIe5loT4e1oRRktFUOzilBf1UmxzXYtDfpoxy0g2PB79I
DXZWye2NfxKes4qOiIDYNcmDuQBQ1EU9NSweUWk7DN1RfpStpSsXRXFwmWlGawP2
u4k3cpw11uD0KqDbBMOebJE0hz7a1hChj0hg3cOGzUMbSCH7StHxaMgCYnRwTsBo
FBAKN3wjpdxlo9Vr/JmyxcsajvMGdMVeOCwKLNm+IVO7K0NzbokeuHA3I0rX7+b6
vtHKGT97U+gs5bi0zWYxvpe550szyOOxm/rGeEqupkblFfyAKttKIuNg/57Lz7vL
pAxnD0SiCuI5BVNQ8TD1g6Gq+zzZGT/VnZFROquq28k7f5+ufzLG+rNMMb0BC5yY
eaN9w7UiTMb3vifXl4/YohmsS7LSAW5UCFkfjEESTeoY7cxtCWCval1eR754/hju
d44i2ElLFAsQmtyKRSiMLm2/TYIaUQikn9WASz2FE5E8vlR8aJvr8GROBgRJrju+
QjImkv3Q4SriZilL64alVuXLfjlbNUYbRXDgZ1R6XbPCP9VfR1h4DoYqT76ublAK
mnUK+IV1EBSNswTxRU8y3iqNqFMHcokR4enatzEvQjV5De5OnB02+FznyLsf1rbX
bqY/lYY8VroOZAtiKRrO02XjJX8Zx3hLaiA8gwJaWiRi1Pl/votjAkucRkyzhZ7T
TQ+x9uhFwOHsArUCQ2sEooZGOrXg2MKNUaBcnTrpBkNNAoWBALVJ4YLgHg0EjYE7
6s71XDcuz1C1Nmj4okacpDSKfdWCtClpxAIt9uJbGo19wldJ7q+R/wCZJNfDr0pl
95VTbcMZRaowYAHCOyBiOAjNrItcRHJ9nR1nyMq5ApQix7Hhws3o4H52Fdzxl3YC
t436AGa6Ofdd3VKgBM56O8k06u6BmsZSEw+dR9MWbYkHbyLX6uIh06UoMu4WREmN
sw9nlzrG/rH/5LyjM1jTCQHuaZ1D35jaXd2rEd8AByju0ZS0RjGmEW7aVAEU5r3Y
JC/4MMy4YLLQnRDGKzsOAAOFm7gsmsXAwmboLhM5GuwC+DvJGJdFnZYega4Zp1X0
5Uo4sSBdnntjMAUkHV2U6CDiSwyOFozjuCagOM6iOLyHURInBxrYlkkJoHWVAdqG
RoOik9cADpRxwtwXvZpswuZca/f13XciKazeZwYzMrI=
`pragma protect end_protected
