��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbI��2��Ձ_N�RL��������lx�^6���-9�D�ߞK�`h2��Ɇ�"�ud� O��D���	����{�H� R���C��4ȸv���ð�A
�NsV���l����/��x'4"����������E0��H��c�x%�֓�[ן�I����N
5�L�Ly>�y�ފG
OC[b�ز�!��q|u;<��V���a��>2tq�-V��	zY42�0y:2:�e���B�C�[�4r�[���È}H0Y
Ly]%	yS��������=|ԇC,�FʐhZ��*/�,��3|١�������A���euцG9��0TaS��:��#�*��L���Q��JVD��O��X�������@�(�m�A����!3���Y-O*�#�X��*F�V`M�/{^$�Xn�p�h?�A`�^I�ݣ�-8oNۗjp5*6rO�Fod�@�g��AQr�`n��3����?x$T�;�89�'�tԸ�rR M,=�ոg��94'���r�;
`�f�p�e)5q٠����E@�4����5k̪4�"�;��s��T=5k�.��S�᠜��=g�U=��hn�<ZW�d%~��p��� ��Χ�1��bj�X!֑5�q	.�T�ux��I�u�y�|�_�N��1v�X���h;�k=w1J��'	X weN�2vs��Lλ��=x«�[�@��䪋��T</������`��.8.T�L{~�����7�X�9���S&If�I����N��}�n�0:&'z�3Xɤ����赟c� ֻ�{��/X��?���#����J�S�]#���hP�͘|;��H��Ul�8��ZD�1���h{�ż�̣q��q)�m���{�$����f�K�?�B=tO�z!�0�dz�#tzK�t�	Yժ�����^�\�9S81�����u��k�V��/��if3�2�'	z2�K��f���A<���HBA��]Q3��*#<_��b��i�˧��K�ڗ�sH�ܿ�8?Q�2k}v
+�,�*�;��p{F/��פZ�q��
�if��Hp;1���z�;�
2��}�/:q7M�{r��՝[�2�
3�D0�����L�/�h~+���N���r�B����c����ηq�aad����WU�@w%N�ʦ�u���Θ��w�59�]me��T�܄rFӱ�C����o�����;߆d��|�>��{vY��������8�
���,��̅I��,�S���La��+'���&׸V���ȅ$Uw��m+����<ص�;��J�����ټ������4�m��Fϴ�#c�r�B0?e���x'�,�&�2�8���KF�U*}�"n��L ��Ua���U�$ٹ�zw���
�q%�-��/�??9R���IL���w�1��4���O1�_�Y�wW�=d� <}7�ҝ�B�40���I��i[��7�,@��UD�v�0�}�/zC�a>5`U�n3�0���4;9f���{�$�"�� _�;�y����>(���Z��5]�,��=��|:���˻��`����8��-��Y�[b���g�6����_�_+"���(ԚwWx~V�b�'Q�J\8�{������?�i��<��3G��2�}C+jM�S��X(�*��
�0M��͋$[s�o�e���ќ�RfҬ^� R4�^^<M[%��
Z͓u�Xx���(Dl��!�f�.��/�x{�OqV\�C�	�hťd�R�`a%T��kWl���L����̞����>
6t]�,��D�t�����gF]Ja	ɄH5�S2+Iղ��Ja��?j&�l����s52q#9��utL�I�w܍ۤ��y�{�|QP֎7�1j�8��`iߥ�w�+(P�a�1d���� ��xsVMI��F�1��Q���~�����v�͵\�vЎ�a����6)cxYSH�)�U�6���N�(�d�&����
����'s�`�6�t˟����QWʢp�3�+]�AsNp��&ڠ�S�v%3��Zu#B]�Vg�4K�.��KuD+�䦓��G����v��,4ޏA�L���^zГ����k�؆n6���ВZ*HΫ�P{4��z�. _A� �Ԧ�5�, �@e�����-��g	򇀴\*�C&=�2r�T�ѣ"�Y9�Vlᘙg+7F=�