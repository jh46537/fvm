��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V����i�E��qd<���2���U���ǵ� ?��K��D��,����W�������:w��|�� )���%�c��L�~&k1�љ[s�o�������@�
�+�۶�����1�LR��XI�c��x�υ�$W��N�(�Y�j�KfE�u~�kKPy���=�-�U��ݽ8ި�Q���\u*)�����ȼ'z������?��;�4�p�&ۤ�'��y|���A� �;����N������f/-%216�@D����g���z�=	��E��<ƕ����L�q25oQ�Ӿ��K��[�1�Cߟ'�u�a����ij�N�o���׸��'���z���߽2�|v.Cf[�Lh~���7x��a�Z�0��=D'��K���)���`N:�
3��Q�b���;��(E�;��3,��Ly�k�5H������y�ADG2�x7��)y�g�+�5ԋ�`�`�D���tl�3Oxo_��3i'.W�@M��r�.0�l��``�}�%�ɤ�'3�ݫص�n��Gz��f�x]��6>h���w���%Z�U0�k$P�kz)�4�*��k���H$��T����-�^;fN���j��l�����
���� �vw����x��,k_f�L�PY��_� )Қ��{�p�~,A�G���Z����'�4.ȅ�x��E%��6�*����F�!��ݕ��*�x�F��BVv�ʔ�Чv���5��4h�਌uDD~����Z����.|�cR��wgfs�}�4uB�!��K��[�U�x�]u"�6�X�0T8�-Ə���F��ahI_4(��~-�N]��krXic�G9t]/�%���&���F>�6��sQ���K,[>'* ���ǿ2:iE���\��Vޒ0�;����dyJ["¢�7c�!�0���1��E�v��?�{�-{�44�E�5��JD��(^�!dw�k'@��C��lt��Ȓ0���\G	c!"0[X�\�U��"\���]��w=Ƣ�y��NmH���
��sַ֙��&y��5���W 1F_u ��}l�k_��^~�Q���SSs
1��jNS��e$���vD���[Z1�O�bT����n@U��J����I�K�3B��:��s����s�VXB]�%���S\W�F~�~�$L=I�o*�� ��i9'u�薲�|����<V@��7ϱT�Ǚ#c}]�S��OD)>�����e�~T�O=: 5t����t�#V؛�O� Y!�j�M����F���u[I��~,��t��}�~��2P"����+���S��)�gs�����P��A�\�o���̞e�\�(�?�x�To�ΑX�u�a����00RxDs��-4��G�JW҅D�{xn��K������,3OYG���e"�q�"
*A�=��܍֛�v�^*]���ׯ�afg�7�>C�d���B<�@�`+l�ns�R���4��_��e 	�=L�i��l}'fCaF&6�?�����8;��w�2�*�g�aZb�Xs�D���#��S	�Ȩ�c�I���9,�97���!���q���8\�}�#������	�P$h(�(�93��);���{ǩB� �)�a��tG���_v�!TY��DΗ�7ʒ�wI��c�bPj���ST϶Z��:t�I��8��gl"�*��g��qp7L����%s���J�.d��G�
|ò3�?|w'�|�T�Y�?��d�^,Pq�\����<*,p&L�-r�G�u�K��\g\t��18�����g0܈�(��*�^`��������>�U|���n���*c� �6T�D���$�P��Z��R�YlKm̛<H�Y�d�4gDw�'��R�o��JW:g�w�c���z,�Dc}8���O�I�O5M�%�FNs�Ε��yn+j�d�[֡�C�63�TX�P�USYO�Fn���@G����KT2�DS٠�:b�"c�S��Q��)�_�Z�+�	���55I�(�؅�����x��#3�\dD�:n�ɋ�I13]B��x���6�Խ�b'ɮa��T�mـ�DB|8�/OQ�"q�m���K��4��#[�lj�O����\?ո ��pl���x���O�tRI��L,����!f��Wm�-�@/����y
���f�5S+�
ӽNլ{�֭HcL~c�����F���+��gƟ�.k��Xp'�uʌ��P�O��͋!�J.g��<jx�1f�V������',�5�j�E�E��� �.���f20��kF��"���>nm�J�rþ���l����/o�c�I]P;�6��h�mM�Ȅò��ku�I�F_[���챿�o��V�qy��ȵ�	�*��tpI�qE�ݷRܩ㒔�f���� ����NcL��@�F�3���	+���:d�4}���>V	�4�?p�����!W�}"/�Û3!���,�3y���uFs��~h��az�j"vT(� !Գ-�R���W�%��/m�=�i�Y
4'�^\tn}ݲ.U��^0�x� fK�
�OB �bu��9^>a����M���������J��:�?�g������\�w$_iYA����g�}HƩ�/`��<��|�N�(D�<�t�}1U5��s��~�����c�	��Y�>�S�w'^f���ak��X��t��2kG�h��C�3H9��+9'� �+.c�vIh� B���X͚T�ת*_EBEf3�68I����Qp�=Fsq��t�[[�H>�����D�o�)1�k�e����~l�Ւ�����A�"0]L���qg��V�[b�p�� �=�@��_���ƲK�Fo�����{��$v���,������6���w�Z����>~�I�=gBaݨ2,6o8�χ-�n�Kp�������!�մ���p�r�㡰<�ؚ��/���	S�Q��O���#���{���E�wy����F��z��S>
o��'0�:��+���
�8�;M����$n!�����->(�-��op��QM�Ο�mN��TG��ǮT��x��҉�o�"~J�	�4�B:���v�(�1E��i�p���CgS4�~Ak���i�IK�K�Q��� 7>���?��$��p���KP���`�8��3l�jy�A§���i�A�����L`�����s�T�ݹhKpq����S,r6���#^����F'ϑ����x�@zK����ت����[����{�hB8u�J�ov��H ��^
��Q����Ϸ'�����N�Y~\�hۍ�̋��Ҁ�J7��D6�rб�8�ǂ�~������<,�0�<�l*E�aҊe��0�������/��g��(`0��x��Ij)�z^�ƌ���ST��J[~�M&wn��ڋ��I��H8�ixe�_����H$����l��ظ:� ��p&��g��Y����c�@Z֦K�ⲯ��wo����:�~rvl~@@��y�>�Ś�������8��'���ɿ�}��_H5j��ϣ�~��F��2������Ll1|^H$�y�P=���K����z&���9gB��j��
ٓ�B���&�"�^���r@_�<*W��G,(�,rS�j���&c�(�+��������Un���{�1xg��/�����B`������s�Ԗ���b�q�-!׿<������H��M��O(Q\1%9]3v"�`��%ɇM�n�/,�n��t!`�+|�@�ZvA䗿�ؤ�X�R���(E�`NUϳJ����}!�~kή��w�ɠ��\���r��o4HBg��7U�a���xA����ݶ1�)�H���K��x��ӹ/�}(��j#_�Х��;,���[�հwZ��m�!1ؼ�H�����]0�LD:�:�dQ�U�������]+�z�z���b^?.����T���j)��W���~@���m�J��n+��V��rr�#�J�^���=�j̢���T\�kO��DuAXc���StA�Ȯ��s3!',Dz�X���S�9�z��?wE��B��O�̍iƉ8z?��� ��c��S� 1���x���B��(�^KgG�������C:x����Kڅ�F���b�X�Ym��q0�뤝�<[�e�M;���.rUʼ�T��{	3��@�n��~��IN�iM���V�lKn��������J��ϊ��$O�r�ߵ.�O�r!;;�*��Bc�D+>�J�_�ֵLs�nD>�7��k���;�1�7�KE�(-�� k��Da��4�e�bQ	�v.�&����9J1T�e�ى!�ҧ3�0�(�G@%4�[P3M ;>,�:��gZPA�
��g4c�:�+!���X�|��Џ+���0J�h<��d�9gb�����I��J;��x`T`�ZrS{�e�KƤ�5��R��(F˂�?�T��Q�ߣ�cr��r�@�F앚5͕փƱ��fi�"��u��O?���㻽�x7��6�֫0@�u�B�@F�aT�2���L���l{��}���WZZ�8 �T��N
]e�}�[���!N�_�[|p����Q�֑�g�?�����j킒P�B�VJqs���4��X��C88�ƀ{0�ۚl���&�b y�]������]��|S{��}߉p'��©������9���SiHE���$ꌸ��"�Ӈ�T���+cz3�WRK?��h|t�:_���hr��K��l[���s��'𳶝��{�n��J�}�	FL|MI��S:*��{��cb�]$���;.�mW��q����R�d>D�O�6yAS�o�|�y�q�6�ՠ�kĄ�_T��=��	 !5hX	ڐ�[8k\|�\�dg�����v�&Bq��X�{���#Dk�[T������1beU�l�Qt�-[j"x	�� �Sj'�:��Q��2�/b�oH��T"�����n�����k�x4���m����M��7��AT��٠o�1�$Xӧ�JA"��Q���l{k�/f�����sK�4���'���&^��c�ȷz��X�rұ"^��.���q̳�3͢��4�����9�W�o(�z|v=��n���bP/��Y�ޝp��j�hXZxlҭuVq �}<��Ab;w�ŗ�b�����f�W�� M�U�u>���#��x^%^�R ��	�b�/^oޑFm�*���q<���(b�T	�N3�mz�߄l&��Q�l"��̩�0��Z�����P�a���A�˧`�o����NPʵ�ի�4��d�����o@Zr� ��4��^��9f)�z��[����Gr����=�e5dGs�>�?��8VzA�����$���3[�B�u����ߦ��<�������_bO	*Ϳ2Svjm�	O��L!ۃɵ,�٘��$'_�%'�]�o_�3�;��Mh/��2%��-���F��?-�'�w<�_��� ��g�c-:�P��bV/��Vn�>�5.Wy�=�~n�S�����ۚ������<���u��R)���1��8�?Y���C󐞷��e[!�($'Z۰�x�����v���;!)�����(��^)��t��Bjg��c�Մ����
a��nc\]�bv�nr1�/�,�J(���%/�e���&#'gp�A�͆%*�{�U�0U,c��Zh�f7��P�Zs&8�E{��t�E�ijQ�Yu��,�02s.��
�OI��X�~�\��żwj�\sw���P�R �B�`0{,<ԱL���v�Ԥ߆�Th<w�G������xз	V���r�3��Bo&S�Ay<�����Z�W���x���QЄ�P�_T�Ș;x�_�W��սa�\�\;x�������M�t�~ݝM/�^�E��9�o��%�'š�O6K���"�b��$�Iv�7.۬³È�dW5͜�w�$�0���=�e��)�v�Թ�v#9w�:�J��6�g	���Koo��ڧ]���S���s,0��g�d	�G?��G���8Ă($��#-6}�]Ԍ3���_h_���h��i�Ơjѭ}T#
_�X�E�����Y��3W<��J9� ��B>B�k��[��'������&%-�G���FQ�wZ�O�M�n>��������нJ��7] �|�;����K�ʌp����H���+��Q�9W�8������-���4�D�����tm<7e�`\e`9f|4�0�"����)9���P>�v`�QF��R�ReC9��:͝A�c�-��@����I��v.p���HG"k����2,��?�"ۊ).ڡ��zUV)�WS~���+�bc}�����E��ml5��?lw��d"�pt��¤M��Ĵ��+�����Tmҥ�j�;;�
�s1&���9j���Ad'�����r����WP gG��ʶ�t�5)@׼�c0bJn�p�Ydڂ�/wi�R^����}�7IA��|'�v	������.�O�F@A���1%�
�o���e�r6�cS������Xs��$p��:Zijێ��N�7	�bb�Z=�D���a��-#�3A� gI{�x����Y��	8�&$�(k�6�ށ`�>����i|h3gjHn�݅Lt�m�桱6���1����Qf�4���Mʫ�w��(N�̜|n�AP4Klzw%{��QM�R��&���'P�Խ�u�z^����v����P�����5�R]���M�8I�:?(�i�-��h���U���ҴR��i���xI��E>�~�a#�fj6��.�P�[�S�|��z�9� 6����K�#L{6���*���
��c)D$��01{���V״#,�eC]��4�H�]��<_���*�{�0E�G��unG���ɮ3SǏAA����\���ڽ����|��sd��d/Ǡ<w<�EC����4��&T�R
�.˽U;J�����=VH���s��u��eb?�W�V%�QR�m���~q����"���2�!��阍a�eg(F�>&?�7�_��;�M=��+Tˉ�L�dD����"�4�Ў;sE�)U#\��#��8c@RW(˼��̋��b��r��'�6��~����w�e�*����v����ف9~�$3�t������2g�R.?��Lz#��d)l�X�g�S�&a���/����wN,ɔȥ+�]3��(��'"�f��h]���~�;�2�:���� �q��GWb
�4��7&�/�-ҽ2���KjK�yS�����HN�Bo�l���o	= u��U@��.��m/ҩu��[���)<��&�68��f�:�@���Z)5ں��aī�s �~h���.��7��
�	��ې� 8�ǭ�
�m�
�"Z&r��,�����T���ط��%,�d%�j�Z5bs�h�����#)�Z�!ğ'q���k���9�����%S��[m���n?�݃�K���D@_����
o9@d���~\V?9� �=�#��J����3�J<f1����>�"&�J˘[ns�DQ��9�d����;��)"0#�(5��pbql�p��{��d�u�� �t��b�L�"������xުhg�1$��K�=4XYy��vQ/U�	8��+�g��d��ao�r�m�������Rb�h(Y��R%�xa*��)��ÿCT�O9V���֕<��;��77��vvU��-,��/"�Z�TBk��>���~�ڝ��W?{`-w���I�?j4�y�n��(��O ��5p�О�w)�^�x)s�l찢��!��X��-O�w,����t̃!�.;r�~��)��nTM荽p�z��dZ w6�<3���I�C�(��kU�P���e�)0ӆ9�`�?�����M�	��<�1��?�~���N�_��.����gX�jNdru &?�f_��u[~f��%=���(-���ޗ9zO:���w��z�����*눱����3K���*�3'�.��z �<S����ay��St{�Ɗ`��,��>� i�p�a=?�?����M�b�����^_[ƙE������q��Q7�d�Ҥ�ӿb�I�ՙ�eeՉ�uhs(I�i�M{���2ᶾ�����Gۘ�p��DaN�����/�Ri��𴟖����C��!]p���[�<� >1)"B��/���K�92�z���^4s�~*��a����'�cB^��HV �\�0r>���G�w�2:�o��p��-��>6�?�B&<��#3'u�0�"w2m��@gS6�E:���TO����YL
����F�ܵ&�A�-�!�=���4�3�x%WQ���`+
��j�]��	��C�_�r���ǿC�dO��D��Jt����Y"4rs<}�[�������Dٺ�p�9�|wz,K�h�����g
!����;+��[ܣ?$��h,Y��᭳��J��鸱�����C7��o���]'��k�C��<��7�����P�53�t��5��\!u:����6��÷�}X�I�q�P���Ϊ�@��lr�"�(w������&M��[�7�$�ċ=�5y7���x�R�4-��Z#::p�4]�O*�=���~�A��D�����:� �7��O:n6<���H�b�L�vџr�\��J�`��b9���ܕ��t����4��Ip{6��>�)�g&E�q�nItJȡ��ڵ�6gou!j�/��)��#K����[�����C�]c.���V���ԃ	lE��
�Xa�|�a�E��z�t�6��+��t2!:#iFk L��ʹ�x�MI�@rQ7w�!��`h��n������ɕ��,{��N&���Z���M���-��ͦ+R��hҡm�Ԅo��g��S=�{�y::��<�*c��x=f�����M���;���֏Oh�=}�+Z��c#�pj��3���*��;�RO�u�@�����;y�5�$��#?��]{/��j��q�\`<6�^��gI����)����G��sw��㤣s�~&�ۥ��(g�ɾ�Ge�����1L`�\�B�-�� =�L�q�.uD��s�H#���Oyo��Q`g�Ǎ�rK��<Ma�dJ��Q9
���NjXi�WxP����u<��Z�w�(Y�sS\��5%�vn�|��ź���3��䀶��̤:4n�f�W�w�?���do��m�e���{z���)Os�O0ր���-~���J�
}���2M0��q���E�t��
�`v����d���"c�e�������E=��&{x�g"��M+6�vK�V��^����+K��X�L�\#ͻ�ӈ� M�@�*#��*V7�\��j�����%�tr� ��	V^��̡�-vI��!�d��n����R�
��@Q_O�m|���w��0Z�	/�{AQg���眥_�x����Ռ�Fs"" I'��ȅ�2�P~E%��� ��?���!����i����n!^{����	��Og�!0y�n���N��� ݪã�Qj�q�h��`�g�-<�~�KmR�-�������u�u3�jQ���Dnt`�;���y�O��;	U?Y^�y�$O:�,%��.�ڨ�Ćx����O j��2q-@.��3Fd��NT�hIoh!�Z,��q����4f��'JL�>ʂ��P�$�+���z5޳��l�(��c����`�b{*�O]P*�]rj{3����U~(t�8&�r33vFM���?���p�1jv=�1ҕX��o��<u�7+"�2[��U���X:&���$� ��K�6 �E�xJ����C�*�v*�M*'�Ӗ$l��5�o���UEqg�?��t��uN�G���"��)�����_����vt&D����p��r�'��/�gC��4�I&
���/�Ҷu+�[�J��U�ah�w�5y���`�g����@E��M�7�M�;U�(��q`�8�� -?wt2e���dl� �-"^2)�ӗ��A�Ʊ^�c��G:�Y�#@�l��AW���zϐ.�b��ݞ7��brT�K�W�+�;�|)(�Z�vB@����׀ ��"Y�Ym�� �ej��5�x��B�i���	�����S�"p��=T,@]���G����i>,_���-i���x��GQ�(j�.�u$�K�8��rK�b�A�%5�)��.�ѩ^Ut}��B�������������c�t$O�j��L��<�z�(jg+�"�)}�_�e��lܮ�W�J��M+�X�5n��PK�U�~ik�b �����C�s����b�U�,�����Lg^�����:�+.e������8�H؍TMf5U��?������ڙ���,|?��`�D2�gK����"��,�p"� ���%���H|�t��&)�-r���5h���[������L��A����n�Ih���D����^̇ʏ��J��$f��,�"�C,��I���}H�0�(Z��,cL��h�؍zLdmK���z���� 2���YJ��}���"��o�Jq�&�E|�\LJ�2��D�� �,��_B��e|P�-��~���!\�4��!\eA��t	��O�2t�X �.`��o�9����i�tA@�$��6��&�*c�&�U��c��;`»�V��jG��#Z��}�g��U����pJ�	jG9MM�@�Ԡ��:44�_0,��a�ٮ5n�t<W/9�|�JU��tTu3ƋӬJ&���A�Mr����A[29.|����V����3��+I�)�tT��m�g�}z�����V�j�B�b���<�2D&P�Pu`��@�%M?N�+���,;O-�`�J'�a��d3l}���ai�R���q��)#yv׹d�)�pn��ȃ�S� B��xPJP�P�n��	E�s�8��௉jg`B�>]��\C.��\��Y�z�E���0��9N6���.���a���[C������e��K�o2��~�9�'����M��A�"]jU��ӜX�;x%��Ǯ�`�q���R�e ��d�k�\_�7�#cJ��uaR^;�u{H�\j��.����#t��V�U���y��c�7�R}\/\ط����d���'Iq͓�������6GF�ѐ�0qX�5v���K����۷	���䝪�>ʽU�u��&�q�c"�U��`�[Ns)vd{��i��u�����_�L�\gZڄ��`��i&CH��������c �b�HK��;�a��2��@[93A�
��$1�l���ȝ��sW�1�w��8/j���8�񒶼[���9�-{X>N�F�kl��S��Ӥ=�W����|lg[ -���w�b�gXz�S�e�$\>Y �X�����&碯�s�|���"�
�Ť�o�A����%�r�Ƹ��8c�6�!�Ub(X�9Vk��%Z]#w�_��l�$�v	9TH����q'��2�(�{F����k��������f0.?�X ��I�,��0E�o|�O;
N��ɣ��9}��b�m�t5A�(=L8qm:ܵ�W����Ç�_r�d���vksY�0%p��3��k�QOw��X�:C���ŪM%�h5��A��P� `��)*06)�?���s>��1	K�,V�KƲ01�f��(�A{U�D�woZN��r��Q�M/߭�K�a�/��9Q��%`�������z��u,�{ME<0�"�:&b��#��'��]$�IH�KG�j�]��VO��+b>�5��Ϳ�s�H��OD����Ĉ���"����>���1�ZD�oV��ekn�E�����܁nd��Hh�1 )��uݱ�N��_�����=燡����/����:A�Ħ��b*~>d��s�Z�����F���Kk@C��`��)��F�e��E�j�z�'��k��B�]����d���i���rR�N��X�/��q5�z*Ě�ϭ�v�� ��0T<�>����^�?��SM�Oxgh�{��^