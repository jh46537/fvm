��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħa�gU�]@)},����ע�����0v����)m;xH�|}��[?���`7"I7��>6Ɏ��b�P��6�8��A�H��0M`
ي*�鸆�k��r�6
��q>����dj�iSK�InoR �%�<<=,[���vT6�Z^�>�z�$Lӱ���F�扑e��yR��Զ�,����
�UP�b�P~J��3t�-O@r�(_>zb�����0�QrE��bO"[%��%�}˹���u�+�T�5��O4~{\�C]?�oH�H�yB�%��3�A�2�dyɒ�^@��� #T�b�@�BF+'�h��0��E�!X�hȈ"^&�Z��)�3v����|�+�IZW�&X׳m�ݑ��=a���@���Ɲ1�6<P?��P���[��=l�T �N�4L"�������"��T�+P1����d�y'��SR!J��ֿ蕷�`���C��S/�D�^<ư��觟��y�f"������~���:0?�#�-:@�W��4�Y�` ��t�V�-���t�].
f�I�Moŭ��6t��-�WP�d�V���^� 6�;m���͡Lv�BG>�Y�o_�m�?��܂���\�'n�ҵ{a%�Bk钤��W�	FѰ��<y�e���..<����w-��`A:�����,�JG��?��2N<gf|)�T���׃���2��H�ߊKZs<�cq!��R�qn
m���"���6�����]���F>V@)��ۀ�a���j	ݑ�a�cS�ٞ�izT_hVe����0��|�����z�t@�B6�ya�ч��b�R���_�=A�dY���|�c8J����<��q��<n��Ǧb���#U;-�
�G���M��$H��������֋��F4����Zܣ2t��vѢ�����itU�57���!����QJ�Qp�g��V�^G�2c~�'�F<�(�Y�Z6g�ig���
��6�4�$�fE�!-����O��B�K��:�RYO�7وe]ND��!�@>��))�AH�Kh/-�����v��Z�(�����_22�g,R�<��9���1�>E���"���D%w��ͥ�P�_|�Z��8������J��lv������
M���[�@���)��P����N(���`;$�S�fLP��Gg���<W�J���FWj߃jQc�3� ���h�N �xD���跊�4�$��O#�@ªw:}��c��[�g�!~U���ҥ��(8�z�+�'Qa'�\M.�}$T�
_�>]�|�Ͳ�T��G^�{gv	�\~GD-��0o�����+��[�w��]W���[0R ��i�._����f�]��S�&b�5�U����k�n�tפya}g; l<%;\����<8'�&��zj*_!G(YH�(�شݤR��43a���v�� &��̈́���CB#��L��w��
*P���� ����I�ZX	S]PcWw-#��F�BU�d^w���z�f���2����p�:jB���u4��]�ǁ�6�fźҿ��Q���y�?�,�9H�aWQ���W=td24J{�/o�~J<�ʤ��o�߽Y�̊R�ݺ`J�P�g�C%�K��W)XZ��4�Ը�w���{�):�!:V�0�욘Y��c��!3�ʂZ�Y8�W~���$;�L