��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[4 �����W<�"h	5�=uk�eb1ٌQ��W+�n>�I�Vmi��Q)k�|>����k]��T��qJ	��4Q�7� S���^�<7<�9>:��N+��Ś���:C�Jv�&T����j��/���=��LK>l{��)�'[x=JHhcY�'\�:sR�G��;ֹ�$�.� �Ъ�����F7X�Ƞ�:�Vv�O�ːʟ�2_�Q�/Q���]1�ؑi��_�cF�rFi��o'þ�`٫⡂���r�?��
%v�z�`&��.[$%��d��77{�X���/�Y�y���C����� � �ł������#�=fVu�o�F=<��"�E�V��rܟRz�f�����߲n��ZL���k0��ҽ�qs~[m�(~)H�Pa��E��ixt�:���|��aF"=`�?l��pf*v��rN{�b�s�(Ce������P/9k�����1��ܨ���4GZ.�/UhSX�^x��&y��	����uҲ�.�RP����a�1}��&	�ؔ<E��%���c�䐨��5�ʓ[K������&7���mo��1��rc	�d�Y(���R�����!'KVe�o�L�mI6 �b(�N\n'�1�jۑ�c�!:{�՜C1��vXSDԡ��eF�PQ+�1�h���(2����_�X9�9~�M+���u� ���*"��Q?�z�'���r7��&R�S��.o�u�S��߂.{��`[I�QB?�x��9P �ݶ�Sڏ��oS�M#�:߇h����)Σy�MT0���>����T��t�s��2|;`ۂ�ϔ�2|���ʦ���:� p�vOzLƗJ)����A:�g�ȏk��*O����W�Lg~^��j�X)�m}�Hd]')q�PfhX��l2Z!�}����t�
H%IB��=J�����!�];�\	4q�U�w@_��&��`��K
*	ع��s���Bhh���H���D���Eu���C��h�&�!�Ιe_Psm�5.��^`�=M�iKN6ɲ(8��I�X�P�P���B5���.~K�f�h�*�o��*�J��+��g�����ʦ���2a���87Ղ���K�Q����r��P��d�tF�I�7�D�j��9���
&��#�ʴ;b`g,�+Z�O��+`!�� QSR5�EP�V�G�>�Ns�M�Cc&2҄��h��;�!��;��p֦�n;w&|}���&�+��]��� ��ώ�v"�j����a��uduN�يc��#)&wY�'dĢ�o�3��e�U�q;*�-@C4J]xf�:铌]vQ_�
&)�4�x�HH%��ֱ,�g�T#&(s�ͮ��$��5u��ix�tbk�;?l4�,�/K��>�q:[z���ǭ����@�&�*��0~�� }����A�w�D��ل()�6W�5���a��Z��y�1��餇�����Fe��1�g��}7������pXm���:����m؄6�����{�0��CZ��DRnE�q�ɭ��~�� ��@�34$+����;7%��vem�rN���#p=y�L�c+���dDh�g ����C.�3=g/G�q��7:�ej�[gPC�$��CIY�ڎH�֜�%F�5=Nȭ��ی�s<%��Ơ�<��N͐�HtY�Äm6h]_�X�oi^��>H#FZY ig��Ay~�!3mDs P}��~M0��I��w��NL����� �v25��;�c䶼��hp{���&� &��߶�����Q����(|� %�V��ݳ�R3r�88uH�M���2�X�d��!˃2 ��6oP��7x�y��d�:ǮH��m��`0�>��s/�(3������v0��l��rB/O�J)�[Պ�zՙ9�i�"��F�	w�� #�Io1/�4��c�o�pWS���0wG��\.!l�!艱�o6��\#@�����A[�@Ɓ+�vYu�L	d�Mt�F8�9G���!�7,�6�0)N�AxGU�]��?ň�= 3����Y3=��3��#��� ����q/C����� x Ԏ��Ͻ�;Q�"#h�����<-��n؂������Mұ����H����^�'g�s{�!�G*a����ҞL��+�M8	�`��o���WLd6eց��Z�A�9 ����� �&��.Ha킆:�C�9)��(�Q�6'>/����tֈ8x�����َ�af�������Q�7�r��F$��0B镜�$C��a��X`���C��JwaL����l��Ok :I�b��eG�f�bc�<�o�e&�	<c�m�'N�E	��K-���O��tk��f#��(Y�7#�v��,y�i1
� �o�B�&C�ԅ�J�ެ�Wv^\vS����]�{�!��"���SF��S�B��v���c�ؙ3W��Q��2�x]��N�����+�ˉR����K�(T���첆�����>�-V�D0h���prJZӭb�����eK�ɐ�$0b�|�q�E����G!4xh~+XD������)oe�- �֋�J젼\I����Տ�@��}./W3��_���	��.�;�|����RebdzZ�`�X�EY�?���ؙ�D�a"<�x�/�x��OŨ�V���/�*j�6�F�TX��z��ha�-��T�t5��y��ADim.b���K��Q|ɘ-�`5ޔ�R��(6Fi�LU��
DRn1�r -%�v�'��e
(E�HGnJQ��#�B�`��r69�R�Jb����Jn��,�("�~�ƇG5���
x�:�֬ѥny>�0��Ο��|7��Jܲ��#m�+�؟�x�9�����V��:!�z�x�,g��h�`R���`������ң����N3w�s������A�tV�a���xE�x��}��,��NH�9�-�U�U�۪���%k7��s'�L@������(	���O2;/cC�B�3@�������֑i:�^c�-8�F��|����v�9���!�s�(�i�.A�-Ѓ݌�d-!��j��SN���SlG�֥p>@�eq�e�&V�Y���Jp��y0�܁��"��QW��R�i`Dو`rX��{��n�9��i�a���a��&���u\ݙO|�'?jX���mYc��(�0�IgP��>d,V������8KV,�,ڿ你yr2�'��6���M�E{��	)�yp�҃zU˻G��N��XK�5�ђ�;D�U�j�	8-�Fa����qق�4�@g>%A��4	@���}҉��ǙM��� m�4d�4�v�z-���]z��lv�9_���xR(Z@(�@��5�;��\�� 8����d�+�MR��R8ANK%]`�;��BB6�*���#`Z�ɯΨ�I(�0���#�|+~�N�2��Uo�v�
\{m�$7�8AP��o�����#[q��]Ř��rY��d�(�$M�T�A�	P�,�3��b��Ī�BG�]��lj9���Od�k�����T��:��$��v�2�7�L���¥�	�p$�$�ݱ�*>6���{8�l<��΃�H�T:��+B޼�F�q ��+�-Cy*aO�+�c�~G/�1h��mF�vp̹�2dR���$�TYIb ��B)�=�b��w�鿅������O�G:ZV�3�ZbgrV�dG�4��5��^�ժ��:�W �^�Q�95�ת�i��fb�h�P�jz�$�t�:'쀓եw=���%����ڞΏN
U7(I�����w�����X�h��X��<Knr��N�=�ǌ�F��kMN�/bFK��!N�T i�jb\�Y���e�r��jDb*&��i�k����{������q��)�u#����0rvԇ9e@��xɭŪO%G�5�3��`�[gTVJF�MX0�g�XTI
�xN��,�L��G�˿���+�w�?:�}%tr-��yq�]}��NW1�z:�� ��>�m��l���MӬt�i���.�֔n/i�ۃ���
Y�[�YO��ހ�Z�L1 ^B.<�#Z i��PxT�-U�3����A������ad/=0�X:�Ôcn���G4� ��M�2
��а�*��Z4Y�"�qwp�b����4�l���=)��䶫�����q�y���pN���3�<Q^m��:�by��h K��(n������'�R�9���v�Z
�2xh�zBq9���>j�xȝ?eb�x^�U��U)�.J��˃�u�Yd;|�� ��[���C,�A��;����@���0��z���f�u�?���'3��?�����;�j���^d��5�?k�Fk|b�* 8�(�c��|p�K?W+K�+P(�[�=�>�o�i�I���r�=G��]".�p1��wm�~3�r�@�:k*�w���m�5��Hn2��c�L��� Y�1�P�g1��b�{�z�����5��/
Ƙ?q,�h�쌯���?HG($�P���PpD����٤�K9��d��7%��� d���Hf~Xs�-��Y�sņ��C���,��o"�)�q�_����^���Q�NC�,�͎!���[p�����-�M���A�(�"(juƾ��.��#1_���L]�
���j���m��=����m̒5e	ˉͱ�?�����6]n��p&��J����Pq�@\�>x�L��4��e�)Ƀ�]�g��ʢ�\٭0�a)6��*�G�[,����b
E5���[��&�Y�H�VǟA#�Uy�<\��:�i�=�=�Oԑ#��f/- �/��Y0�K�qz�w����;�f�l��đb1|��U(ގ�S.B���0���y|g�g��l�,ЫC|��*s��?U�ݡb�1�٩�r׶�@o�Qf�X��@��_�p<>Y)A*��$��L����tʞ���[�9H���m)�ߔL~"���ڬG-�6���ҽk	Ÿ1��ҥ����(8�{� ���5C��V�G�z�7��Գq�8(s����=҅��łB����0Ky� �������l�g u�
��LK����a@���SM������l|&�����{��������F�`�Ѕ������[]F���V��C�.�,éw�?�0	�j0�����w�	G�^�\���]�ͫa��?E�M�څ��K�����4k{�K-�kz��"t@D�����0�u�Is�E�Q	c��49�|�0�ئ���|��ۉ�,'[4:��e �PxW�� �a�ˉ��j�MP�$����C��kPv�X�V-�S�����:������G��Kd�x�S��Y�uz��2�W�ߦ=D�2���v.�5�w��N�*ۉ|4��2g���%|��
�`��Ҕc��������
�����UT�&8|%�|��a��]FA�ѭOQ�!�B,����_��=�J���n|u�򆐯�(,��{׍���]��^�}�����3�9�H��ӏ�L� <׸-Wq�(�]�>�!6��:1U��ͪě9`��Urf�#�R@��=4�֩��@n���5hzl�
�'�R����Ŭ;�z�������6^�m����� N_�����t0`㣖�/���ؖ�M�!Y��SO��6��B�u�a�,���s2��xip|J��_v�D��*����{�)Uj��a�=h�6�D�����Y��*N��ɞ��MOܣ�︪�E�f�*����N�IߌR�us]��]=����r�rzT�-�B���m�#�=�j�ڷ�G��)n��h �dߨ�7)Hi�k�J�B���OYU*�$  ��Q�M��Ur���Pѡ�!@g��&PS��V���c7IqwXt�����)2"@�Jl�f)��g�|��[Iv0��yD@h\���%���$/#罨`>�����B@_F؟����T>D9�� ��)����:�����[8�mM`�L������V�3vZ;�&X�qӔ��#�����J�}�\|��[�O>&�#��+kO,^��(�W��[�`j�lhw.��L}@��Xu2���az��i^m�4�kMû�o��������T�}z�����M��6��X�>��� Ԍ�g�7�A/hAY�;��d��À�]R�w��2z<6�1㳷� ���_՗�����_��tښ47=�J<�@���������|���Gc
3O�~�InV�b������>��_ʔ�������x��%���/�%�(�	�ݘBɍXx�
���o�y,�w���-��&\��]��_��4^щ¹�p(�M�jF��N�K����&��!E��/�t����&�"��HWRg�[�ne����I�.�>��%'	;��}m+vkM5Er|�V��.ƥph���W��ME��C-�,ǃ'J��wIJ��k�<�n�T0���9�ubc�vk�l�M/fM����i�}�z�>2~y����hĘ2��r{ɝ}o:$�i;}����ݮgl�jښ�x�k�����P"������\�~��֭SX{]��*��,���>�VHK��E(1��0Od�$"����! >�_���OOL��> ��מ�,�=�zثpq��ci�#xCjٍ�)�]�䳰p`Ys�kJ�U�)J��T)��Q�/� �A��D�ՌT�e�"�����a&Q�Ͷ"�z:��UǣÒg��n���O��g��)[��{bg�$ͽb�I�7U��"ZXĺ��n&�e�
ڣ������?�u�c���Rb5f�gd��!u���*�;ݣ��j���Ǟ).��-~�c�	3�~oT�vG9Vk-��,�)w)��*��2��Ǆ�jK�	�1PbH����ՆeEVxy�;��
��|W��܉�3�Ie�)Z̡H,�n�i��v�Ml�2��K���X��@̠Qﮉ������u���2[���cA���9sE_��)�^Q���f���IЩ�NO W�]�t�?���-�;�ZZ�^M����R�[k�����)x��5��Y�I���������J�Y��c]��c5^�����!kñ�M.h�<��u-It[��0Pӭ��4�����]a/����a�#������%���S��+E��<4�������򕶈�.%cx�/w0�-�%R�n� �
��]{#�x��+��PST�z�/ix|���#Y*L�:��OG��>B��K;#a�?�B߇;JNTg��jBo��J����͈h�JP�Ӆ���x�;�ty��.�E6!����ͤ�w뷵(?E� ];NW����N<�A�!���N� �6���W� �sɋ,֐5e(�c�?�b��SZ���'��J��=��P=��5�9K�lY�N�N�:
�ɔR�B�O!��=�]�-��J��?����W[eX���R1kV���6�я1"���NW
��-�^ ����}��e��!��

H�Qi����Yj��Ķ��pF��2��&�wD�ӻॵ�?�Y+�O�$8�o��	�d��2���ŸG�/�I���h�� ��y�E|�l\���P� ݑ�Ju�z�h0�'�AH &DB���\��z	�Ͼ�����v�oO���s����袝%&� ���m��͋�B�7��8��s��������x��S��7���1"��i���)�d�?5|�"[f�!/���6��#�a>��O|���-%|euoᗀ�鐋�L˨�?�k��M\Ȭ�4�PԪk�>���o��:B�{�(�U�;x?W�������������(��|��L��i�C<�v�=Oa���i��w|$�B�����l6�	k35a6�f��N��>o	9љ����&�`]>_X��T*��r��S�����)�N��J7�q���x�Q�>�AD��JdT!�[��Zo�Q��9��GL��h��N�l0Xt#�V�l�
a�1bzE\��)��FKuV�+6Y����%\"���'�E�xP�M!#��w�����edH����|r?��A����m��P�k0AՃ�d8�{���d�,��۾^k�s���$�IpJ�΁q�_�;�W�עhd�"X�&m����U�N������qP��Y䆯��l@E `*FGd��F��5�d3u� ����6L��12<槊qgA�w���ƨi'����W�Q���.̟]֯��fN�%��Y�TL�u��/�i������ UN
�?����tvݯ^)Rh�\ى٭�'�sƼ~��b��h�������G]�"���Z�vSfV	Q�LI&���߱�<�VT��<Z�|��p'�	���N��i��R�)�--c�a��:MZMH�3��_��� �l����1�e����x~ą���)�DNk��4�An;Q��S��_#!������ky﹋i�3>��񞈬�P%�������T2��Q@���I�4�&���f36>�bQʆG�t��Zj%Z3戗{�0�ez���l����\�},�k�V^�%U�"�@��$��f������e�������� o�>ܶ�bC��l�X�R8���ς�q�?���@R�'��G��dQB�b�vj8�0���9 ����I�ȟJ��V�* �c�Ft�q[���}�"?�7{���Y���z��/����cneP�������[W��/CN�4 ����6�tr@�l��|��i	�=�hhl�������9$��.u�O}���*/���IWl}��b91Ź��+�-1���\��xb��k�x+���r��~�x�|Ihι�9��Vi2[UEH�.�=C����
Q���gWIJό�$ϗ�h�)q�J,~�lL=Dy�J�*�xdx�}��Y�O|��E�9�4�i۰�S��K
ϛ��E]鱦R&�|����Hgp�.�$-�_���p]��p����״�����ƧJ�.�ڈ�;*������
��am����A3�r��-*�JWk���;%kZlv����&İ��p%TpG�G�gb�ϗ4��T� �)M��z�o�O}��t#�L?�Ͽ	q�;�	߯�,����'���H�pW5yND��W�z�z�GӁ��� ��(g�nwMq%\t�&����B�Q�Ye�XԂ:ƒ�M�t��wI��qz\.u%ѵ�˴����tP�@�����="�%9f�S�ʹ�x����2	5;9�RZ���
��8N�k���-�}; bNF�g3�nfxܡ�*�u�~a�޻�n�S��aU�rz�"�x��c_�B�k��k��s��I���b��������:T��<U�6d�����yXD6KIş���C5�d>��4i��T=}|�Xሔc��"��E�N��:��E����.���x:�����.��O�@�;qs��ӘɁ)��v��7[rD�w��"�p�M͌a�B���$)xE_Mػd�crN��K��ſH��wzʮ�]�2=s<�܍}�����Dy0m���OAć�*ە���0���{�ˡh������8^�~*1ίH&�xg�1̋����%\i=��r�z_F��/�����ŭ:��P4��ݞ���=��G����:��jl�ݾ[#���<��ж#�/&d�(Z�TH<�t��&�K�����e1��|ULL��\އ�ȨXHG6�_�ãLf�}-,.!'�zi$8@B.2���.�nm	��9׾ՠ�i^��Q��h�Ț�:��c�q���p���!TwiQ��ɕc�+k{�ᙪ9y!ﭵ����6�L�]�b�S�s�Uv��Ȣ�bG��k�D��D�#=�w����M[�=_$�bn�Q�]�u)�4��#d�}�
��Y䨯^�1���=��^,�1�y	a����xJ�@�%�:�@�Lc���p��/��]���ޙo��@�k�Q�KNF�\�{�yz���1��h���/oyн�����E����1Ǌ�� eH�N4,K�nq��:g�<���y�c|5\C�H⻙4BN����҇=�a.��;�备}�%��Kiס���o;���� W9R��}��Z���2�C� �ȧE�*�s��>o)-aÈ�
�u��p�^�|Y��T���zcs���O���7�p�#ҫZ�O�\u�Y�c����7K��r��DU7�P(�3 K|��׾��KuNi8[����/,�3����D[;�@�L��_+��&���$ab�SP��aTw��)�-zso"�@(ߋ�E؅Ѡ�}�ȆIA%�uZ�L�J�Vz�gS�Y��|�o5Ñ�0
� 5P.��.k�ug���H����f�u!�Bm uC��L�V!"%3�eB�/X���� ���6��Dk��hH-Cw�ā�lw�9�CRԷ�t�k���}�z�L�N{͒��;Y��+���F&lNс ���.�P%���b��0�a�����VV�݆��w�ì��U�K]�uX
BJ*B��4�2Q�!��������#�L��6\�^�
@z%U��T÷ Q��*)��L`D%������A����{�k�YX���?{Ԏ���u��m��|X�"-}�
X�sER���Zp��K�(>4I��ir�|��J9��	rG4 �<�:T$�I�P%)�f��e ���?�h~a;*6�rR�j8i��M.����F�Yݧ�k���vpLI}������-ܕ�.��0�7�X��f�����'�زU���I{��0�kL�Q{���:n��̇�Z\SS����h⹢�(@U�N�!�.#�h:��9�p&�M\���{��ܤ��p�3�m���di@+_e@�=��O1�刅U�~T{+��j��8��RK)� �5X��X�{s/�_Ql�E��kq�u镆��d�Yd���\왝�v~�ښO�z���<�l���
�sw ���j���������M������c!����a���J����W׶f��c�'����&��em����Х�y�Y|)2�Ur����+�z��H���Q4+�z��v����]��I+'�{��Zr8������)��y��
�y�R��h��5�	ꈽ�?`w"
H��q��`�������4�*����v��%��oX���-�W�o�Z?����.�P�3q$�s)����t	���{#"bu,�P�>��rbs��V�B։�[(S�1
>���`��1r���,��8�3Qӳ��V@�VuG�NY+����c�D���(,Na߁�=���+������R�m]�^��ΙlY6���9����d/$UT&��ѹm�Ba�����_�ƃBW��vD7ք� ��M����^(؆fC�:+��
r7Ř��"�@1!����V��S4%�
^"܊]
 �[!���0�@r�����Q@ ���56.7
M�Q�OO�3���j�]d! �|���I��r�9�Ń�5����'��@����;|�0E��]��VM�Α�SK&F�B�`�$Ň	�*_��i�E�W�f�(�P����C1݉�}hh��1��\cF-��Q������H���S�(
nȄ��5}��#�e��$Ϩ�H��C��h�ŽoS)����&�S�I����M�������0��<������R�K�+)����ϙS_���� �oG.ߟd9� �a{��]�@me`�hT���&e�J����c��K�_x��I��j:qE����v��D�h��
���e�v��ES�AM6���B���f�8�d:U�j���L��q��4�A�>����1xR�*�%���|�Tvԭ�S�а �k�q�S�jbi�ގ�"E�*�P����nm��]Qs�v^hω�gz�Ww6�e��}��2t��V�u���+&9�?VXi
V=�L�ʺ-���=�ߗ�,ym�H>?Y�������tBr޿08�J�IҦ(t�B�\�(��?��1���H	4�P钾��T7�o���!U�zZ��W?�D0C§��]���í�B��-��X<����]�	�D]�g������
 }|� ~,%�&M'OU�oW#�5�i�ˑ��Z�	P;�g��{��s:�9r��;z�?�t]�"�:�W�*��t���<XpJ�J�����ϑx�x���z��A�u*���Y��1�̴	.������K*�V�o��xY���B� [���s�-���rq���I?�u���jTf�'�w�MTy�GI+`QJˬgܥ��LL��r��(���8S!e������o]q<��N˫{���
N��
���-8�EW~��ƅ�V��7U�R\�4�?�ǭ˧WI�O%rX�?�������7w@z6Ǆ�Ѱ��JI�y3b��+�������u�����d�@�����}��+�{jل_�n<�m����^��5�y2.+�@G��{#�6ܿ<�k���
gX3�*�sB����alz�A[w ������Fub>�v���|l��@C�k�Q�� �zY<}�{%M��b�����t("�6g�� ��\���Q�hS��˂� �@1@�>/��ג��4���Z8L���GB* ����M��D@X��t��	���p�uz�z�rN,JǊeBxCh�(�d�]�f�o�F~�>i8�oD�l8��^Ļ��޻�d6�ڤ�~�a���M�0b�C��;Jc@��y�U�,�F�`�)�*g���*�pjL��˞q{Թ٩W���ɻK����&YF8�̊U��$�=�j���AP`�Z�m��x�;I] R�0hQz7W��C��G������ʃ@�����	�ٌ�� �6�pj���b�c	Q��A��XZ-���i�۔�4[q������%>��(��1t43{MĻ/m.����[C����ɔ�M�y�B���Tp�y�>��{�C��zs�8n���7��<���e�R�g魩��A�ok�p��,�s��*�ا��#�/^�Cnj5�[i"z�&X$�m%~{��I��n���7����\2{:q�%WD�w��m���❛�2�+@;T�W%N�UY��	iQ�,���^
���9�b�se}�Ć��Q����*mVUs��x�'�n��p��B�� QPɳ7fw����|ڪA�j��$��:�V�5�u�)xDF
��üu�Ǌ=ڏ��D�|@]��~6�	�I=&�#�VAu2�yuء�O'b������,���:�E ����@�:�X֎%��
�b���O��f�G�Fg �G��b����*u9�D�Z�ڿ?5S�,����� ��"L6�O���RW���o��:���j��SF8B�`�S*4��F��Lq��l��dH�s(�OA�Ȃ��IX|�5���]��'�E�!�Kw������K�"��+�+��x;7KWI[��O�)'�' ݸ�z,Ka�H��^��(:,��H��Npe�4]L}�
����.��O��*��b�ha[�d��]�<�wVC�O�:�sLs7ͻvE��l;�[�I1c��o�}cKT;����~�&���A�o��	@�}�������<W� 3!W�Q?iՂ�dӆU{�G*�q�ۗǽ��ҳ<@�#�!����27��s��}�:д�
27��W_T��Q�^�i��ў�KZ����L���,�mmP�l��]$
f1s�����d�+&ųs�(���Wd�ԅ�lZ'�M�MR�#�@)�9��
�:GӚ�M�$��+��4����;	CQ
T��Ꮈ���B%V�1���mNlq�1r���l	SS�/�����ǹ����c�3�@��E�p*��Co+��g9�#۲�Ʒ�W�������2�#������7��IƲ.X�A���������Θ�jo�IY� cB�QByS���>��
(�6~<g���Ls��������?|�A��1�X8d�{R_�ۨ�u�X�,����L�ix�z!N�<��7��@Rе�̐l�vAr���*��$ㄱd�����s��&6���.<��q���1����+U���f��cu���GM��1�SZ�xD
m��_V@2Y��\��w��>b-�e��h$W�$3�5��S���$���{��*ƥ����;�\Ս��ƌ}��D/%EL��l���A��NS�Rc��sn�I�� :rH+^�o	z�{}�]���#�h �IJb:I��m��Fj\W�`�d,@���1ה[�����7ֶ��Y���iG���NˡE|/��P{����,���}�QI-�K�D�f�4�h�r���	5�����^%WU�<f�b����<Z�<^!�i�>� �(6LH<9���{v5�6,`F`59����0��T�4q 	8
�8�&^w#�T�Z�z�q?���\���@�%=)�~=����o����BmJ`��r�?�ǊI������?�O��
�b�wz�H�IU.�6=��khQ�6�
��4���δ���FM�+oqmR�6��h�f'��O�4o�����-�_l�0�&�C�C������
���T��]����0v����.�J�����9�s�6���z�XEF�-J��`,"X��=(Y&�_h��J�uj��&)�Ƥ�ӯ���i��� �`��we�Ӳ$�!��fݜ�����^�W��Xq[����2��^�ij�]U4�Oyw�ޒ�,�l�ƞtzx,�j�V�m~yW ��M�Ox�#��������N���2@f�\�!Wl�����i���·�q&�" (`3���԰o&�R�V<X���5���}\�,���#�C)~�j��g3�d��&�6�I����6y���z�-Dc E�@~�cl��/�l�^�����*���#Ug�?���lI,>wKlb���w�0̷����2�U��[�GO^&��"�\I}z�g_1���Ѱ����ˍl>�>0�Y_ ;�vS��OW�E�&v١��"=wg��Õ��o�y�2��OF/[f�/�)v;��zIP�˜(�c�"Ff$�>��'p��y'�S>)Z�|/kz�}�;��B�{!�G�����E�m�oY�:R�>�} �MB6��gK��H��i���`�ʞ��p��mwx6�פ���t�9[:J&��֥ ����y�6"��T��bɨ0��	�'n�>���`=Wv�
k�L�l����u
�_*-��@��[Bn��!�j�R=~2��u	�rМ�G��$�x�MzPU�m��n�$�#�v��%��+WF�h{��_�X0��q��,����T�1�ߪ�0t_Eտ�.�.��/�����?��[�L=n���u8Q��y�N4<�	������ouA��KO�o�@�7�҂J��}�?�/U#����wZŵ��'N���皃�s�){��������r�۶�[~-/�x�^2.{�tזGs�B���� �1h>�T�*�\�L�	�$� ���tj���E�J�G��Y���`ClP�y��!$�#4�L]��*�;��]@����H��}�0䦲�J�F���u����&���M[��X��@u��� ���N��da%-#T(��m+$�:��'�#)� �<�G$�ꋼ�6:��T���*;�D{Vz�<lܖ���k}���B�2t�t~[E�l�l��o4���t$�@�}HoD[�2�?өA�"�S�Bߡ<���+i�ȁ��q-����U%5w]zL����.��G!�Kp��>K�1w��{S,ǿ?� �O9�	�F�VV�k��������	�>�^Dg痎��RT)ĸ�&���R���`p��uGhx��H�+7�I��D��e�m�0�S>1bTɓ������`�RS����м���JT�Y�j��3^a)Ǖ�45E �/sg[��v���@aX�.���?���U���n�e�m���ֶ�l���°�?mfӠ���>ǀV�3�pm`��J�F'6�ۖUb`���a�"��ӓh�����1
��A��7!E�W'\j~<�[��Q|�h���\��X���
�Dm���%X_��
������	���V�(&����0���[ ��ՂM�ω����6�W4�n'G�]�ob�E�sÆ�"�%~��cܛ�O� ġ�!&��!�����g�]5��(1>ܾF�V�2�g�LT�;I��Wo&��qοk��Pݓ���n\�N�~���V��yf�)����m��$��o��i��S},L�K�F��\�HAO��I��1�c�Y�Cޝ�9^��u0���nD��Ђ{�P����qYx�C�P7Qj� ��	��t���k>'<�?�r9��I��hs�_�4�:�caa/��A�941�jf�
�M���^0��Ȧay����lޢ'=;�I5z�z�0�YO��w�u2$rhʥ>��X���� ���H�]�6Č�~���_��L��ǥ�Q��<A��;%����� J��'�(�H�p���@4����F2|x��i�,��]5Q�"��z��c:S"�1�?�䏔�ʥ�Bg�c�V�P�P��n�E�1��py���	����n1yu%ǀt��p�mӣ�`޻%��c�Bߠ1Q�q 
�/��Pa.+��4�����qo褦[���̬��5��*��'�6 |h�;���������=�U���]/����y��".����K��`>xً�A���w����u#��j*�w(��Xy���2�'�<�X_nZ+�#�S�!�k ,-?�����s3�eE<! F_���Ϻ:����U�`"��쪱-�O{�W�'ٴ��(�R�ӷ��C8�]`��-��s����V�g
�ۯ&3�n��Bq�`�Wp=#��q6�cX/�س�r܋-l,�/&�Ϲ����Ӱ­<�PҰ�X��z<�*Ć�}����8�7_;^x�;��c�lq9��;�1m�"7���3�強��a�Z�f�֎�x�;g��PV�P�$>�Xt�SR�/sgtkpK�)Rt�!:ʅHU��.e���6!+:儇�"?�([^�σı�������ȹ7 ,_k� �n �r��S(m�vf/:9`�@��i��c]pJ̘$���N��p}ij�Z H#Pn6���e���B�܍��|���6y)�;��m�rҎ:����j��%��N���B�$hY�e����o���g������}��p��g۠2����<��{����Ӄ�f��"a松�����f^�� �"��Y����q.���d�l�PߡG��9xU�� v��1�E]�^���ė����\ 1I���UjJ`	'�oX=n���!�
�[]ⱀ��,�S�lx��: �*�
Tc�2�Ѭ����Q ��r���c*�sɱmʥߚw)�*D/�����u�y�Vm�3��g�a�3^ܱە��s�T�C����!��=�����d��Ec�t��&lEg��ڴ���Ӛ���S�;`d�/���qB�ˀ��>y ��X��@n��nn�*�sH����A� nj�����۩a���#I���o3]Ȱ�R��S%J矓-�LF6���J��P�����e��gY����G'3�^�e`4C�\����DK���L�+���9ڸ/�z��>v7�F�a7)!�t�W�|\i����/��2!K3��]9G���G�G�j���<�����L�/?�X�h�y�Wp�
Q/}�2�4�򴵢.5kĘh%<y��ۭ��H��&W�o�&_Sg�aȫ:�^� ���ey"�q�j.�	���[嗠�E��t߉���:
Iu( �^��A2��q��cC��BΩqPad�w�i�R�������Xc*�҂�jtI�e����e���+�U���%�NBs`�ߚW0��Ƽ��Ru��5ե#L�t{X�C��T�N��9���,t>��VI+�����NO0�"H�S��B��z�#��G$)o�����~5@�m�6��G�3�DɔE[a������W�@04x��K�e�o���Lp�:ߙ�8B�~<��$Sa��U���ݦX�)�Q0\-q&Q��AˠqX���k��Q�$�1�ϐf!leU��N$/f (A�{�<Ӆ�o�ՙi��yr�_�#�Py�u��9K��i7xh�l �9d.S4��B������ic����qڼ�H�C�Km�4��?��l�1~4ǢN���(���@�����u.��6V|���PK��8�BiɅ����+nE����纡��S�h^�)q��S"�5�E�=��1v��V[���~��6��M�2�_ơ����S�\�tp���<B��>��s�uz�(O-����9���="�{LD�UY��e�7aI8���4����c;r~8��z���	ëz�&�����y�@�7�� �i�V=����}���*�`���m�N!莆=DZ��	T�O��:�$잏'T�iv�7�X�q�/w�'J8�cN�ȊJ�:���"H��i\�E��!�}��R`�U_C�.v$�e�-�K��ŭ�\����"���=/ԇ��W>ye�=�������:�x[�&K�Q�p��샒kiH����>�-�Y�W���V1����5�b*�<ng�M����Y����׮�W��W������2rf7��"�p�U=�c�ܡ��s��~MmP]a�I�réks�tx���j�CUf<��$�Ԅ]`&L�83�|z��s����{��H��w�+�q0��8sa�U1n�e{��R+�J��xӑ �5~���cv�_�}c}Y�?��1�5L7Me�ES�����fD���f��Z211�F��L'�4Ү_>@�I��K���0Y��O�S���W��KC�
�FYza�8�������0�v�NA
a��z���k{�r(�@
s���4R��@�A8�|kچ߀��q�BO�s��+�
׸������9-�m{�Ri��FG /U] ���N����3D2ҲH,-�*���hY�3�1�KQcK�(�+����zR��!9���QY��hM�P0�s:�ϫ����D^��T	��ۘ1x�Qw)�|TK�e��my8P��X*��V�S�!բ譮z�s�b��& �q:�W�(~T�9mn��̐%�ʊsD|'��W����>0���f��AP���x
����[צ`-��Ṵ�<@�88b%�p���#��hA���OT��T��?����CӺ_�mnК�@=s�������v�l��	���������������7�vb=�����(\c3��[�U�p@��l����/�/gA�@J����1�,畍}ps����4���a��=/	�m9��������#�[,�$��D&���z�q�8115��w�
v|:�M��X����X�In`��E�l�4�1�޸�����u�����rk��st#fH�?��L���j�pc+G�<�3dy����I���JGV/H�����`����3��Z�����4L�i�H_5	Զ��G�$2a$�g���nк����$L��EqXl��	&t^T�-�
�xZq�]�,b�͑|1�?ҷ��Fbn�Qȇ�
	�	�8�kr."���@$i<�8?l?p�G v,V�S�;����"�,Et�ȏ�7�,o��s�]��y&���Oh�~J�%�"�f;8WO�/{}��zZ\�yiN�h$�-�� �������#P�<���c�z�������3�j2;�Ζ��XK��T�@�1�^vYY�w��4�C�����ٝ�2Q��a�z���r5�����#J;8�\ǈAT��<,�d�o͛�d4cz��p�,�=��E�\)`$	��q����U*��n7 ) ��{9�=�����Lg>[jx�xci$}M�ܞU��v�5������t��!����x��Wҁ���G#�~�����fm;g���
5!D���6�ve�oy���
m�>�-	��n�F�ȁsZ�AL,¿j���[}�DtcR�{%E�A�Xh?u�"��^� <kG;)fq���ǧ��|ơ���+>V�� ��k���$ڣ��)N+x�������<���&.�e��g�i�?�_��R܍p�"HP�-���DyO}K���q�Z�9���6�P��y�s�r�v����5��1��%]pO#��`��^*�
0����勉bvd�������uUl�Yt������v�>�j��ڙ`M�{��U�ʸ7W��* `�o'���pHIw{����A��cwx�<������%L��SL�5�W4/��H�0��<XI���y6���=�_3g�gxoҴu���U'�n�ӲC��\��{�bh��=jA�E���Y�ǿ_|�_�	�;��-�;}�ݥ�����`�?�9�I�!��38t�T*�fj:��7�X��T1��,'\�e���;�H��%����]+W<s���$�9_�.q�}b�N�*1v���eX�ă�4[�SR�����p���\���q���g4�Z�0�����r�%�w;�$⳺w�!��O�y5o�|����#f��åQ��F4y-\t��lθ���F��1���.g�jk��K�N�x1:�F�����"�AZ�Ls�:�m�l��_������mK,9My�U��Fm;v	���Ic�R��}�/�6Q�9�	|<�w3��Ԣ�cj��J4z5
�Y^�O~��K-n�[�����K6R����E!!b�#��<ܱ���o�'f��P�2��-�Y'���^d��*���0��\� ��ur薤48-�i㵴�I��S\��@J"`�`n�q�d��X3��w�ё�Tl�8�V�f*�!	3xW9
�?pϭ�@PL</?��9ό>��w߷�X�jaTJD���TZu�MX���{��2>���H�+"#�I�P���+��`-�s�*�{�e����:�0^V���<m�?r�*���1΢ǪX�����JA�+���U\�n��n3h�w]�ꖸ��W�!]�����s�i���,�Gj/�KI�0Y�WD�q���0W�+�G��Lx_]�=
ѳ��7�l�K��SȾ	��R�Ϋi�Ý.��ӌѲ���)������.���)c�����;T#<uT�%�7a|M��J]/h`�s������n�6�$p�&x?�P�cA��k�B��s =ͱ�'���oH�<�|�Cm�Ѽ�qqb�#:~�%4$[H��:lg��-g�P@��x�i��z��&G�)�vXtX=���|��6\Nb��3�;�l�6s���h������^�Kſ�%�	�[*�.�{�ބ�dX�RH��5���!�q@)I�i�J.x�T�.V�Ύ ���Iv��Ѱ>Q�%V_���W�A�ѥ��G���0,"�_�d�-���cyy�� �&>���xߖ�� J���e�=��e�7�!G�G�H�}w��)&L�;����ݡ���q�Z����Hʜ9��T��9��/��ub������r���� ΋�?rU�k� ��� fKs����y3�����`.�e'��g������e��2TA�Lb�H�~.N&��1gWQ���5���`>nm���P�Ը�f�f��v�Oހv�Bpǟ�mH� �h���&'��-�n������ ��EX��9f�(ቪ�#k9p����������a0���ļ[�ws��&4\����G8�v�����:��Ɂq�6qj��Ȝ+H����}*�f�v��#��)m���I2#^���^�3��*l�,��s�)��Z�	h�~]"�4a_s!5��,�W�#�{TR�"B����
����[��
c'ڈ�l+����O]  ����Y�(�KN��	�4����73���
;rf��&f�P�q�-��㴖�F^��PX�1L�P')��� ש�E&�AI-�-1^E���;��X-%F5Q���!����0�# �ɽ�>d��XFc�GP���g��h�A����,��i���V{%���.��[V��Ếl������"LV�tE�jTX�v��-K8 �'/&T����/���P��Ǔ�
э�ȝݾ������s��>U�K�N�r�Y+�dv$*a�	�� ,lU%ȡ �k�+k���h������^�������$�`Y����,8Ag�#���rg��ln�4���8���16��W����� ^k�3�/��e��Lͬ:|>�3��Hs�]6��\$ّ)�E;fJ^��J��� fծÄ�CV�ki����t��1��Ӓ�ږǠ�C"��D�-�E|n7d��ָ�������B���O4��	p(6�7��C��^zsI�㹾T������R����V<�mpU�ʮ5��z���ɪ� �>�~E�Ȑ���"=OA�uXfISڙ���(z����� �S�0�A�H��N��)q8�z�zVO"A0�;_VѻW�,��0(َ�[F\T�[ss�Տ�.0b�G��Ko����	h�c5
i)n*���T����t�	�X�AU���K�'x�.@gr�� �ڼ�*�.���z���%��Q�zE��WD ���l:�l��L,~?+lj�P�	򝒍֮~7ě��d�k�I��q�X��Y�=:�\�^���q�����}.�Z>( �4V�Z#���M�R�ȋ�>��v&6���$�0�hBV�zjTAG��Mټ�F��;��;��p$��
CCJ3�Ǌ�j�D_��1��c^3��kEDr��+�c
��w\���c����<�>���YcR>��=Ch`;lQ�ӊ�*o�	AG��V�Ge�0֧����x5���W�C�[�cl�]2��r�x�ŧ�ݙk�$�e���yðwx~3L�R��8�)�oH��{�� ����!g���O&���=���Uc�δ�MN\i�vD/�%e�(����<���d�6�k�߷Ҫer�_�З�����҄A���x�8�~k^��"ַ(Tp�\���;��9J�.�Y�[�Ђ�=w»6�Q݋͍|�:�,5���zb�I�?�>ש�nc��������F݁��������^��m���$�} z���0-;���I�.��� �;l	����@@�Fg��3bg��sgL��w(I5�-�<���Vy�Dj"y�Z��N^3�+.������t�?J��.=H���_�	��$nb�:��z{�J�ŭs����@���kMd9ה}��M���I����q��)0��,~:�_�%�֞l�r7kMtY3�`T�J��ӥ`]����s޴�;~��S���в!���ǡ��yЮ��Q�1
�@�ϻPM�ά��zi��V��@�f+V³ׇ�1��(Z��mJ�VԖ�P�G2{����g����Q�g�X2v~T��H_�����َ�S�[��x�Ͻ !��z���C��`6���3��fl5:��$Efc����5*�R`���A@�"�x ;�OA�1�@�}�����"B@��Ƨܑ���
4��P��F,r�hF��I��H�j"��~�����E�޴������D��_�3����ެ�-����M���lU��% Q�5�aA~�\R�񾒵%��C��R��8����[R�lj��A��"K7�*-l�BR��s��im��b�::�Wq�8KQ|#���0R��
���5�p���?��l��,\�ΐ�nvn)�A?�/����דl(��Y�Aj��u/w�vՒx<��z�8��E/^�%�Er���rQ4�1����3��U��(z�c�G.l��5��9 �w��^�q�se��վ6wLFћ��;���,�.A���}���|���f��F1sy�����x��S��q%�����̏�n[.��H��T\
����79.7�	k�l�p����]�����&�'�x:󦐇Q��� 0y�"��.��}%�����p��V��DQh�ֲ�4���8����2�]�q�i��u~VIC/E�v�P�u�~�b�z�w��Ly����k�4$�Q�m�F�{m:1�Le��dQ����c�L�N$��-^�%��\���A�۰d��)��>�P��t@k�a�yp�^��c)��ӱp��m�z��GgUn�;����OWs��ɓM�w�Q�D���}r+�ب Ϋ�q�%ʻtL�:��H|���)�E�7{K�����2����!��t��l'"M�]*?�0n��F�E��-�J��IE����Y�_JC{Wu�F��E }��P�!Rl�Rcb��h�n��ʠ{����_RFI�n��~�����='D��/͹��cZ�Eש��Bh ��F9h�j_c�<.�h.yx��u#�D������j^�5>$<C�S���!E߳�K&ˢ 
���E�P,��� ؟W�X3��8@���V��*,LYR�I��>�Ҧޭl�O��UD� * s�@���T�v��'���gSi�h��A�P���@!����R\eSWo�YA��g!rǑq��}~�����/���n�~�zjo�p* �*��k�����6j�8�l$F2;��]T2��l-"���8�) �� ���0m,+�T�%W����v�9?Bi|z��ꔩdK8Y��7:Ʊ��;��B7��mp��X��Za��Q��O�]���|D�0���N\R��G�fbæǑ���l�1��ěV���:�?W����O��5�E�-f�H� �Q�j4��WocӪ�C%�}�HX�T�`��� ;PX�ѹr���.�Z������⁝���kfn�~~~й�	�*Λ��7�*�cg�~=�	�Ѯ�2������Z��U3����2�[�SG\�U��A�<�ǔO�	�خ�6��z�>��� W7�5�:����\����>�,l'��Eؽ�דLL�~�2�x_\��=��ӗ�����қ�0Sэ�~.��*�5�k�$���~P+�?��f�D�{�\%���~�Qr[��2_rU�'ܕ��g����e�x)1M�U������`Ys�@-6m)mZT��~-�pŤ`[�	�s���u?+c�OQ�u��~��-�F&1P�@�������Ʃ�X_��f��>ѱ;�jy�Ri��ݗ�[r��q�J-��z�ԍY�O���_��
�$��TX����iޝ���0��%cU�Quu��MK���:Y�ƈ��A�� #]�}�ԕs��8��'lm���K�����*(�4c%;� �����Oy��y��S�n���Ȫ��}�����N�MN&0�5e����,cv�!-8�����R�r5���2�Y����M��H�bd��n�q��L�JO��v�8��]�Mm�4?��?Cc�Q��t�#v`7ޅK/692��ş��!I���~��g�w � 
�C�er:�[d~z���8�d�x�bm$��=AyY,D��u��|@�R,����3ȸ�?�͂[z��jBb4)�=V�D,ڽ�M���~�ڿ�!�22'j԰�>���P̺��!Uz��W9����3xطy�]���s�u��|��C�ځ\P�d�
�L΂����u��0Z�v{�g�ȭ%���$�b�;^a��v$:Z�%�
#:��!&ݳ�m�x�����t�!�_|�:�
����d���z�����wv��i<Ʃ�����c��г�.8�@��j+ΠJ3,�p�f��&�PIM��3f���yzM��������{ ��ަ0�4<e�6�9�S0噞�9]\J�.����=�h����"w�Y��Uy�n� �ٌ}P+ԛ���òD:W*�sM����tI��yCQi��Н��3���9��i�ޤBh�+���A�cQ5I����u�#X8�q>�(�ɱ۲j��A-�N}�c+ԧ x��R�۬����|�X��#4�V���4���<j�I�M��x�л�z�;����H3W���%�R$^�T���,ܿ-�7���W�~V]��G��]�=�2���l���~��w.��S_P��2�AJ�UìBt*�|ǶIF�"����������ƒ��H{҆e{a���a��l'��[��@��J˙���+�A���z*?w��G��o<|�>i#��	��qR�1���j��0Q���1�)+���.k��W�U�m��D��W�Vd�������.��%3,���:���ָ��C�^ ��'��l��ځ��QG�C
,����)G��.ZWQ����
v����?H���+]��Z��!,�bΞ��*}3��,���T_���臼��(Oi,��14?���3�lj�|J�'+�h��ƙ#URL1�A�p1|��eLa��|�%��9���>����e#�O+�=C���x�P����~%�
c���K���מC��C�i?��:=���=�e������Q]�9���VD�x� =;�_�f�!��`������ҏ��3�c$�!ͫX��Ǫ�+����.��oM���q��{��ae��2?��EV/��zh{J��B�9�"��I"�&.���w�M��������:�F�-�}U��]=L�d��%Q�ۋ���a}SU$ ����N��;S��H��v��ec$D�q'��.�:��(��iq38�C��Mvi<�����ok՛�4i+̬�bH��x;x]I:-힕�f��@�����@��b^�������jZz K������f�	�i]��.���k�����:�?��O��鐧��W
�R��QU�Ҧ��OUS"8�,��>�젅vp4�� Ѱv�ġ:�����J�.�Bu4q�GGX0֫�����(��ZF��I�H�Y��CN|t�ڿ�*_є
ņ�,�\�*�k6�����e5��^S�ȣP�f53��g�K1��z��X>�Z\@i����O[~�4�%��@�E6S~�1�1�����N��m+��	'Y)v�1#B�_���Ps����' 6��gR���2K˛p������8p���{z�x�������~>�h@-Fw����Ñ��.V,�9�ׄ�sm�=�,����뵌ޱ�ЇLXG9q����Vn5؇�엘��e�D�Y�q[z���6��������05�߮��i@�	tU7�/�1U�_���!����cn�D+�%n80_p�'9r	�����o8	�/�����&�69?E�9�H�����'�`8�X�5ɀ-�!ӵEAF���T�s��cͳ�m�}H-�H�o9k5���բ�kq�	�{Q���w�Y9'�~l������O=�ꎐS�*ŵ<��+<E�0��z|���AC����.!�rjl�	W��%ŢW
W>�3A�@R�2�p����������.���m�;Hp��O.r���ב84g�d�3[���t�bDmv%��-��K��dYk�k?�{g����J4�@��q�n�R	3-�}s+�q	�G�jȘ�¯�<��<��󱖩�)�U����<:F�F#_���,w�� |v+�qM���g�:�Dbd��9���|<>�����#���|2RD�p};�fH�VG��d��&� މ�OO�H��e-& p]N�Vʕ�A�hܵ��$�1����7@6�	����o�
��@��v��=^�Er��sd��F��G�d\?��8X������}v|�vN+��H6{����#�䃸<| � �ʄ|��'��<|`f���I��	E`8��b ��%z�Ѩ�O�>+a���b�KG�N���q4�y�`<K(�V;0x�40���k�
��h�;q(��J�=\�w1�~><����\O�o�w��,�%�-��C�(��5Z隙�{5����? ��a^�B��R��C9���գ�'��h������3�p���E�ω�/w�����5N�ôoɝ׀�.f�!;E��6��O���,�������-9�Ғ��:��C��j�=;�s����7����Ա2��v�ґ�O�t�ﴃOx��z-wS|����u�7ɪG�&�oA��5¹{�U��M���/(4�0YZ�wD��j��2x�	���׋��D�:��~��h8Y"�d'��R�s@gLa�,��O�?Ek��=1�E쉰܋���%[!����%��sPyiu;_5ř�&�)p3�t��1r}����E�kF�zI��Ñ�81�4Z����2pǢ�a$
�q��]��s%B��OD���2Y��dX�ZRH7������JS���#���YTpEz�ʌ�qns�_���=e���BM��&'�ʔor���Q ����	,/^��6�@��g�D;�>W�>��KK��Ӛڪi�����_8+>a�����J�U���-<a���/]�dQʭ�'`咱;a�,��R�O�:Uta�K������y�2�+��o�eх���|Ћ���h��q��	g0��[�,�H��/�W���zË"YV� ��zAAubw<�a��o�����w���ӠѴH�Z���HB _>%0��9�����=B 5L�=�1�����[���]0N��W�~�&<'�a.�Ǘ̚�\ i����h��WH��j�9���)%�ҳs��?/����/5v��I#�ջk#�W6�� a~������H\A<��6�~��ǒ;Xw'`X؎@�HSN�}y��@!�!�AηR WL#�B8�av��[�wY��Z����J����49+��vE��6ڳ�/�M��D��H$�*Y,ʟ��ˀ	��g�+�Ge�4%��5^I�ɜ���V��bE��������yܥ��S&e{����0�;"�o\U����ƦQ��S�8g������Q�ac�C��|#�:�A.������	�I�;Bg	��W^z.ߍ�>*�CP@ORC�0gǁs��T:xR�R�����T�soF%X��K��o�r�j�zm���k{~8���Y�����g'ֻ}W\�0Ů�z�!��⢕fP�oLӫlE�c��X���a<����Ǟ������,97�LX�I������"��)��M���9�e�r���� A�kr���R���4����tsh��pr	��|��lr#�*�
$�
�Z�����)|��F1
F�>����j�&�6	J��+.^��Z���Ibx絪�$j�V�f�z��|W�iı�����)A1u5���O�l���X�kH��J�3�/�%^8/^�p���s�Go�=�c>�L�~CG�<k,x�����ʥZM��Ƽ�<�t��Ip�\t~2�` 0^���@��<�r���Ţ�&%]
=��2KE�ù��8�wp�ChZKf;8�0$k���:����^.�O5����')7r��.in��8��2����6.՚�-���/i�,���N\AED�Y�7����	���3�0�)����v/����C�!Ο�/�i��M�+�a�	�7jY���).���^�U�j���S��{�{<z���q`R� xO9��U� ����jS�@O�Z8��r�t�.~)��6e�M&rє��n�%��Y�4�9RS[��� Nio�(hšf���#8��59bs�*��S�g=2��nj�{�wB�3�K�&N�~�Ue!��֏�u��uݠ���8~@%=2"��h�tT��~����J����R�q�������v�.���#c<����b�w�Of�������I�*�H�Ť�]w���͍�#��>5�i� Ɋj����;<4�wћߗ�>o3y�;\��O8p2�^�8ǌOc�03z��D#m��Slt>��^�֣<te���@�3d�5գʁܐ&�P���qw2��<�b�?�u��^�D��"�-g�7s?���x��vm�'�7;��(�z!�TɈ��|���$��x,�=�@*���k9��H�]����b�+.	*���}��vȅ�i-��Nh��;s����qD��J�=c�@ѵ?&��ˠ��#��omY���b
����G�Ҍ�7v�Y��d���eN;��IJ���x���o��_�c�-nN��wL�#�.30�[d��@�Sɽ�5����&� �4%���K1|��esV��kS�φ���;���r��"���X�����ђw,�缅j��P%LH�s��`�q�cl��[H��F�I6����<=�j����Fe\� b��$8�ф!�c�i�!obqkBܶ[����K���N��M��'��U�U�r��'�9��m ��/J&r��G�^KE 5��Vj/�ꗅq5�6
>e}��^u�p}X��i���C���(�n�H���m,�~��k.�t�O� ��JL��S�f1��J[?�|k+ޣv���}A��t�*O|_��jŊ(��{�([�23O_�9�d0��m�1��������nl[��S9-[��ý%�~CD�c~�i��镍�X{��t1l�'[�=��0,[V����]�n�Q\;�h�p}���4���Y�"��I���\�U��C��������,���'�R**W����ͺh]�	��os��3 �Q�Ĥ8(�T�]5é�ir{���t�c.���7,V�9�w�'�r����i0�jGwK����Be��;&�1<d9���3��}��W�>ٲS�"��:%��ճ�u�Fn��c�3�JU!��ɢ^������J�B��f��
����{D��;T:��1��7"��PG]���.?��먝��;���.\��h�I���t��XvPw�я3,a�'�n��w[�_(m��x�EI:un�AGf�_�Xqf�	~�h\&��c��ih.��� ��jF���gtO;�#>r)43;�5CUv2
*�2Z��m��c�P��Κ�қ�3�+�m'��
�J/3�=^9N�X���ǂ#OxX0������۶��Ȭ$��\wx���	,�)y�[���t��RJ�s>X:�\&ߨ[��x� P�Ƨ֞+�Kݧv����s��Z|ؔ`��������+���/K��wz�	_F�L�b�y'CQ�NP�@��|g`�^���ZU,�n��"��i�$���m9�*G�V*TZ=*��c�1÷G,Uk�j�Eh�
���ihVFBZ�C5�?߷��qO �k�U��<<LT��_߀���7:Y1���3h��ٖf�P��2鯅_]�-�����E��b�Ę�������z�÷ſ��|���M�]�vG�Y�P������Ľ�JSzx ���¤��*��
�����Mr��������.�d;ѿ8;a� ���E�(�%)��u(N�U~A
�,�mC
���}��	�U�_��&��M2l"�̦���9�u���f�M����$_*�Nf�|�T��TI�I��tѹ@d�O巴
޹"���O:1x�'��U�W��6�Hү�pL�>2j{7��3�"߰��'�y����׃����K0�&x2�c�ǫ��
��N�w,�r�t�Xݼ���҅���vy�gOd����D�%;��=SF�D�Uz��� m�'U,���0	/�ߟ�����?�)<���X=�Cu�@�m�8�YU|g��a��VI-�De��\&.1��hW�XP��������ʍ�T(=�gQʠ]M�iɐ�� @�A�
9/�X�%xx b��B�V%����-���,S�0�,���	\�����������s3`�=�~�7v
�@]�|k@�������Y���j��pc��,u�=2�ZÙ��/䮧���Z�ZưM��-��m36G����%�#x@�{N�ò�Ow�-��`=eƨ���-��妏�����	�@Q"1�9���j4��Ē�"�d!�Uw6�3Y��'�X�=�����?ķ����Hx���-I_�����*�
��"�5	)"��?� R۟����)�_6G��PJ֐r�Hʁ7���C�����q�/MoK�[l��%ДS¾��?���D��)�J_�I�nv���$Y��[dzQ��4��il����?����ڃ_����Ƽ^��β45| Qc�S��̹�U`g�����Q5���V�t�h�.�.>���ȸ^��%�E�&{נ|IÚ�#�4?���ٴ]�vp�� �٨���5݂)_*�姥�"t
��K|�D��U�YUܾ���97�IN�����ne�c�ג��js�@���(Ǭ�%k,2�����#\s;����em��%���[h��l��z��T�&(:}5��"���������y�zx=���+����a^�m�����?L1�`��gOa�0���yP��$��L�X��x{#��R�m"����Ӌ(����+ b���U����ksџ�="��F	eP9�*��������>Ģ�:����������y�!���J�v��)�L}`��5nn��1��?G6�C�Ȏ}�ژ3f�5��ۑ1�UL���xt��r�)h12�z��E�d��Ō�:����!�˩N�NH��5؜pO�3<�d0�Q�v��QkI��b5�
0a��+�I[V�u,�|���B�|�*�r�SsV��zM�D���V� |�cZS�͛癴>#Ʉ ޠ���$�ڭe�in�s�3Ȋ�:`y�ⴈ��C�u�f1D+��6x�#Y�z�D����1 ��k*��v�d[�+�je����yo���mN���g\oI-�I_`��I����r�wm�nPy5�,	\��4�fl�I+frB��A�z��i\�Y^��|b�a������7E���	9�h�oWeVud��j����Rl�q0w���<�~3\��18}E(��)��)Q��f�bnI�Ф�o��݄O�揄_�R7��kՄ�u�㳞V���y.by �����vcr�d`��LS�a�D�\r����/� rč�C� N�5�uF��}�L�>��v,h+MPύ��U�N���Q�{�ӣR�ES�ud�;��C����ئ�VM��(5�y'ѧQ��0��k����-]�(�$��5�N�G�{�{��u㣿�����|��*"(��VO��q�LCl)ל�	�Tf�G/b~Ջq�c�gݟ��Om=��y��M����s�%}���'�9C���%	ܔ:ݗ���;Nto6_�[�d=�:C}�8�a|sE��y��������>�8ȝw�"��<_J=e�픋�{aa�h$ʘ/�9׬e�k�>3jJ^��`�q�&)�;1����]��Q�I�a�\��t�s��	����{-n�=J�H8m��D�����ZS��fݩ��l���EmR,���`���1�<Cn�ѐw��,�;x��!~߰)��<�B{���	H��J�9��gY�¼a��;2_������]�Gt`�M\O���J���'g��u_D�u�^��*�6@m�aF>Z�?$a�XO}�=~�����`-�W��W+�`1�ܩ�pҹ�vչ�u�8�ˍ�k���f$�"��/'���
8��굒�@�z�g��?pr)�f�[2����GL���K�2tR�j#���\�*�)�?f�A����I��SBi>�&u��
~���_! �A^X�>w���ሷ�
�l�~�C|��|8\��l�'3�v�-y�=�Zpn�k��=��p!��(�3���)̡;Sx��m����+��_e1E������t��Ia��@!�7�찗$�k�mZ���a!���G>��j\+��-�Vu�̱���s������P���Y��?�&ʗ|/���1r��A䰗]�2a@oSCgV���ɮ���g*���w��L�q�t�/���6�T���{|Z�R?��ɟ*��#e^l���b.��$T��>$#�:j�>�<)[��.�e��s|d��vyZ�(oJP�7+I>�Y̝�'?��CWާ��XW %O]�ݘ'w�7{�ھփ��?]#��ܙ�E)J'�$��y=��^OBW'}�'�I���"3��/�Cw��~�z#��uK��O'��[�,:�Ձ`��i�(��X�S�瓺�}�1C�P�KTc ��U���#, nڀĤ:ey�I?�$5_/@�ڧ�P�T��b!���f�fP�K���������'0jAu�$�+t��{���l`A¤r!�Ғ��nk�D�pTB|�S�����֚E� y��W5���'N��'(gAMÔ��f*�ig��Z� g���x!>g��K-�����?��BLE�/�X'����/Q&��c�k]��j?]Х����D��*T��mg�Qډb�c��p���T������`�SU�?��ߗ��Q=��	��ŌHU�>`u�lx/v�PVG+1�ll7����͔{�k`��&��������|�'�%��rՈ���rEY�&�x�X��#��hC��u�G�
Y���ȶ��J�Lv����"%X�ٜ(��5�N�Q׸��m�4�4ɇ�;�V"w�`�@,�F��|*#4!�$�R��.0�O��6p�vl=�&�$������tۘ�s7����#�/�{7�)��T��<
m�\�&K��#2��Z�����V7��.����+�9�by�̿ڏ��BV�e)_W	�;*��x
99�NM�Rb�Kt����HPo)/5X�HyH4E���+��e�F�Jp���Y��\"�N�kmW�v��O�	�e�P߳�����	F_>�C��8�(���q	�yy��1�,Ǯ��^�L�wg���w�C�Bӷ8lC��j.z��RKSh�����2d��8����0�-�Vi]։�I+�{�@��z=����G�S�,
��!Ȫ����.On^Fd�~��p&���֘g<�D2<�=\��u�%�_6�	��%�xB]��;� �d׏��f���H@R���mx���&��Ђ>��ɰp��fU�-�� ���Յ�����\%�n���H[����*;T6`���{��TB��7���A�P�g"Y�s<Vw������6�)@���MJq��CN���9�G3	Z�I|�d�q{T~lPXAq)S�]�S]���R�߼t��	�4���,
������a���@	�gO��^N�ҋ�h�uE�ZΜ�N�f��EF�쵰��]^����_� @�R�}�X"%�ޏ���Ys�%��f�-��?����}�ioԿ@i-����M�ܽ�C�� /�O����ܿ��yV�.�s��!C����nu��ƿLb��KE��[�"D���6�[�:_ ����̄���EV>c�|^8�G�K�j4N�d0����Kg������ƕ�E����J
���r�/�X�pJˆH��jU���3�s���A��R���������?�۰�0v�|̫�x_������{#�k  �+�e�D��ң��^�]V�s'H��I��0�z5�U��M��Q^9ڵ�7����n�%��h3��*\��i`M�me[:��<�d���� ^f&���Q�l����C��OÕ����+P��f4Ќɦ�L���KIǩYD�Hp�n�q4%*��g��$�Cc�8��I���p��a$����Cܰ���O'�q!�4��H�����&�g/ܙ���`�2b�f�wtK�OR�"�vj� G��_M�qMe�=O�n�R���mf�����4�p�Y1�63�> 8�޿:Pj���i.N��_�8/M�L��s�,LĪc�i����(�����VBDN�e��� t^yZJ�6��V�=G;��*Do��	�:<r�.�vz�#m!�)�	R�d�ac�/�Xq��6�#�)���}żUK�"���+1}�n�Ѣ-0*��.ca��V��4���jr�*�M�ؤ@Qm��a��9�\�����+�s_J)2޴��p/����=��+)�Y3�i�I�L&Z(Q�b�zy��]rQ�`�8ގO�+H��E�:��9��i��[6��S�s�ˣ��\g��㻴�&�$�x�/	_�y-`M�>H�E�n|�ˮ=h��N&q%������DMC��NL��˜àYj���
	��M��Ǧ�iU�	d[S(��Xp�5Rp���ϊRB�/��^}�%}W����(�D:���x��6m�Q�~'P��e~D�|�NF�%������[2����|ҍ:��d>�l�C���7�a�J);ks��0�SVlQ�/�q�aGH�����G@���kGF�m�¾�8L��gy���o%U!Ii�Co$EXAw�[�v�1ӬU�8e�Yϲ�8 �f��솝eؠ2��f��9*����E^P�i�i���e�uYr!
�P�D[/E35�ݓ��X&�e�_�6��c�]gE��e���~�祜�k���/+���<�*m���K0������Xy���&N�N$}F�9��?��5��|���I[��j䦄��dh]���(�&�$N��%_H�#m󘎊]!T��q~��$`�<����2���VۗI��<��x���_@��RB�ú��~~=���L �tǀ��c��񿎭]�J�g"o8��S��׷�ѐ��N�T�HR2c�� ����iܸ����m�tڛ܈f��£n�j����>_����yFO�J���U��s�j�E�!`$��K Y�+'�٫<�����2N# ��X��܍b���''�����t����dZu}�1
$H�T��)�)�n�q5����$<��l0�5W��y���z
.� ��Aj�)�"_��s��)u���u�O!�]��m��dB���;kj3���r����+��4�gOq7j��zń������"LE�ob6Q�G����T�Rp�,@
n�i��q��&}4i�hQ!|��1��L�7ȖG1A\��a؃���K�Yߟ�0M��yf�s0��k��H��د���ۘ*�>>/���21���D���B�j/`�9�37����c�kv�Fmx����X5	ͱ�> ��:vLZ���B�-$ދ7G7��Y���.����6d�j}����Yf�)@��JJ�G�mu�s��|�֊G��(����QQ��lb��2���4�z�l�@I}j�CF�`T����X��̫�1�,�O�H�0�D����ɒ��᪳�q�Lz��dT����E}f�N!���?�5}����'p����P��g�H�0�5Ac����9��7e2�q��5[�L-�z|��pe�+h�������	e}O,��p0pj{�	�F���%f6H7���5����L���kg"<����)���7��������Z�W�����{,8��v��Bd0�n0e�`�UqՎ�����ѾLTt
��K��Q��6�B�u\����Њ^��w>Jѻ�é+E[���O蹽�M��]H]�D�y��?��Ł�sA�8nG ǝ�?��iS�*Lo��VSR"X(�MH�0C·h��=��L|$�$��]�1��1U*� Cr���~p�:�@�Ja;��ͱ{D�X!i��d(R��	i��XDH�F�!��ч�ϩ�,#T�~�z�8 �ю�<����o�a�ϒEX�O�k�j��˜�����Y�W7�ӵ)��L��+U�z��2�r5̈́W8�w��T�̟��| 37\�n̔b�C�!�n�a���6�N�It�&i�4�+��)iS4�
a�@O���q���N�US����{�c����ܚQ�^�l�v��(539�)����L�.!���G����=���b��z��h)��Mŭ��ƳX�i+�쵉��Ao)c"V0��`��B�Ňu5mp�2����u�V�"���ۖa:�L*;\�r��^�,$�.$�D=P���*���mr�g����작0��S�EPw��7�Wj�~���'�6�zI��J��^k�����F>�|]������h7��u���8I�BS�Zj6�8�l�5"%��=�����O�,��� �L�	H�n6!"����ss\�gDv�gP�8X?��g��ڞ%}'�b����==&Z֣��в�o�{�czpɨ��mYgف1�y3��r�F�
c~�5�P
j �����|6z��w����-�$�j�Q(G,J��#nWA��������!ϰa���<VV�$s��t�-�-��[PZ��A���I�K2౩�67�F�<�Tx�p=���O�#�MK����>�}�)�Ŝ�僒�'��.��$��+�~���/�y��U�/
9�/D�1�r���d��2�q �`a,t�3�'��}�6o/p��&Y�x�C�{j4q�5��%Օ��"�xNTf$�>�_�i��z&�_��>�(Vw�����.$�ɛ�A�z(�O��4͔W��LD<*&���Ȱ�T��ɒ�3��k��N�ڢ0
^�J����K��U�^��z*ع+��&We5Նx�+\ �{��a��
�T�/i՛! ΂�����Ɓ�yM7����d����!Ӗ��NC���q�!�ϦB�Zz�T��0���d��
C��t�5!�+A���������?KN,������C���w�VM�=��������/��[e��
��x�/r3����W�)=K�Lk�S(>��h�&k-��}�b���0`�3��욋��t������򞒮_o�5=Tq=������sa��M8�ƪ����PPh��C9�s��M����avl��3�7�v�4T�kHS?�����r�N�y(G��HF�.�z ��!>\x!| :����,��gCi3��4[m�5M��ߥh�_��¿6�&�<�_�v�;�V�m��*1ZK��p�pc��A$�Š卜o��x�8�����^b)r����؟֢E��+m�� ��8���x�+�vF���.�*�[���ֆ[����%Q�g�aN4�k=�	t����P��y�b�S�v�}̎k�o��8����$#��ϫ�>�B��b��`�e}��[,e�';פ�'r�ϼ�������ᥧ�/1�VSC��f�>LG��o���
Zb�N�r�گ>�V��1��0Y׺>�4_�y��*7��P�{���:���O)𴦰���N[��f�b�GG$�l�,z�f�)ٔ�6=�{ոGɈ_nr`�]�-�S4U�7F�:����j�"f��DJP�$�hm5^��%�`��xRn/�����f��v��ӛ��8g�KjJ�}ۑv�LI��T���P.5�ů|�8s���=%��|����C�eb[h.�c7�u���<�^��ϙ�i�������^J�D�+�W�2U��sÇ�3u�tc͠|k�.�J��h�q�DF�=�xm�"t�Ez���w�/VXC��n�1��AQ5������E��8ۏ�$C+٩�����B�ׅ4�f��P��$�wP2I� $�Ip��{��X���I�a,��^2��\����w��9�hi���^����/�	��Kĵ������׊ĳK,��`���ш�d�J���	�9�p\)WG�U�) �Jy�sО@	�T�}�B������{�k<P dQ��nA�(����q3�86D�{\��~�f��k���M���N_f������Ϥ|A�>��މs�j<@(u
��> ��t��%Ό�fj���:�7�k=�X�*�DҺd̡ٚ�/|=i3(�"�b	!�*tv%5��_��!W�?�F�}��]6���L���?�<݃��/	�le����r����u�ׇ���u�j��D9�����A��Q[-��F��m�u�Ht�~51N�>9���_r$�*�=_�d��ʠ-x���ux�d�ͅ~���k-�������Fŋ�h$��_ -���x��(��N���㵷��� �u���,�ַ^D
�+�2��?s�V���Nv��t���yuɃο�s��B�I����KR����o*��ef����~�R0�2���4v����"4S.C���yp	P�����+�Z��3���p�
 _���D�[��f3nj*<t�.�E�k�SՂ>��^����}�Ā������K�������5���D��|��{J��f��J. ~zޛ���_�D{%�5�V9�1\�BDý���1o
k�3��[tEB��Á���X��h������b ^�K�ƹ�����zq1]]~,��X��*��s��A�RYM{�(�w�7Q�������3?��M�]�����7|
a��(^�W���ep$0%��I��j�jVA�a��u�3Ox	uW��	�����:���׋�~o"�Ih�
DU6\"��L�)�����짢{��v��,L���lN��V$���-Ծ�������Z>Ji���>����u�{���z��!�C�-�gp������>3����l���<��g� ��U�6-	����]('Dl��a�UD6y�*�v��St(2���cGN*:u�5�8�N(���YnZ�u�|�����Y@��&"v�폜��w���67"6ñ���*�h����o��ƂG�E4�(����/:-G�U��*�� �-�����`�މ�c�,���ym*�K�� ���}�Ï�Q'�n�,�O��jA:�y5L&3���S@��M\?k��3g�G>b�S�͓V�.�P$3���J�&��錶�"�p{��\��y����z�����h�ݾC�������pYa���G�Y�,���ʏ1���!O|���n����b<�ɡ�1��* ��/ �l�`S�k/_�v�f����?��!V�֣�G'NI�
Ԡ"�4�	���4 �+KmA��V��y�=�����0Xa-�lH���c�rǮ �������n��~��J̵_u�'���̝;�&�D�a��*4�ȺZ��ܣS�G6?�;�6/�Gd�vv|�ۣ��mz���dɿ��×L�����h���M�Joe�4�lV��*r���Zc��7��$�{�%9*�u�
���}m����nx�u��W�M�m8Ɯ��MtC13�I�?A�{�!�$�<ϯ�l��'��g_���N/[x�����R��x���,���-�,�-�+<)8��������G����6ԅ��1�>���k�48���9@�VD��C����v?S�[�M�C[`f޲��}~�1n�E@�Q^H�aҽ3���ؽ��l�����_���۞C�r�ΆQTO�[��R4ʭ��X�ևZ�uScU�d�(e�;*��5��T�+ڷ�'d���UȱZ��N�D165�"���}�LQ��-h���O�e���$�0��њ�(&��/���J���>zg^���\�L�x1W�0�+sS{�/���h���*x�ڮ���9�I2�2uh7�BY�Jtχ�1�������$u��1�����hbc��*{E���[�ܫ���=*�A�h�&�wW�xߵNdX��d��n$+��E���M����bbS_���8�N�k�
Qf�G�a�6�d�˯��.��ά�>X����0U���&��h}�:�!o�.�WF;@�_�N&昻ӐP�f�ߓ��]p�