��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���q����f'����U�S-Կ���Q@B	�Pv��IYgD#@5�gF/����|�����L��9;�̜8�=�6�Ө�m�@����)t�z���0t�x�z�]���m*'�� �~���td8(sa9�7����G�v0ԡ����0 6��u:��m=�׫$uS*�V`�bd(g�����D��J���c7h�k��z�����Tb�9v�{������|�=4�+Ǖ�o	�ٴw����HfI����\%i�5����8qq��>_b�h��a���$�Lu7vE��y
h��D*��d���؍�:��+�i�Wtb����D�sh�92S�X�Lݳ���?�m�p秘�����!�z�60�A�c�R��{yE���44c�G6�����+
��.���	�֘�l+�(E2���d.���Bd;�v�l��P.�E�3�19�?��ſw2�D��s\HAS�%�Z�|���Y��쉨�R���)���g@�P�|��6&��W�1T&���9��:bl6��g��3���Av�F����#'�C��s����7��
��pք۸�U!Z�S���q�(~i�t�DA�(�u�Q�f�Nt4��4����7�Ұ��7�r�:���a��@�M-�G'�0��4Q�C����_���tf�������<<lv�쫙R@(5?W�#vw��g�K�U���o���eq�74����.N&��L�)�бU9^{�U�}}D	P�2_{I�{�[j��H;F�dc��-��� ��U�A0�=Y�g�K��&�-j)�a���{L��9�"��7tِ��zS �<�i 4�b��q����E���N���߸�>g��?㸪����#K�`��a�l��,�`���Z�Mo��H���x���1�*Ơ�Z��V$�o�6c���{v�Ɯ��bZ�/��`:24�j2?<7�]�dx�9�3�Uu�1Y
A�~9�*T�ʴw�n!�$(�>�����s�}���E�o�U��X<��I`�Y����>uRE�\�\܎`�����;�>�f��Sf��!T��\�S����8��o��h.M�L.Ctu!��7Wl��"�5��`ٛ!^K�C���ʤ��N�?��t�u��cJլ:7�@��Bd�2K��_X�/��Ig�E/D(���a������P�wg>�h�YC�,S�`���o�����%��z8�T֋Ө8H�Q�֡r$L�U<�V�/�i���^ "��[�h[If��Gy���;��v�ȗ}��W���@@l@�#�<�ktbm2 e���$���RQ|�z%2��� 
���t���;w/�H%��Dp� I����J�S�xXI��Ǿ{�0n��w�˗>Ds��F`ج���!���F0�����*Y�k �(���'Q��ɬ���$*J�Nbz�C����d��{���㕔�w��X���n�0�������Be�:���6��z�l.B�%�-����
��^�Ϲ�Wz�����e�͸�nEw�=*��Yx����JA��e�EQf���C4x0�P�0f�\ԣ5�fn���uBg��LiU��^�!�X�>q%~T8ޔINSw{�s\�ꜹ����xt�=�C�O�Ut={_��K�@Է��v����R��g�ShmM���V�d@{�\�U���8�pL����ɃP���j����T҅�L4�ay���!Ț��9�!`f�Y�T�������Z��aZ�/�<�L�C���r6��|�S�%+�pC"�%@��략��`��c���w�b.=@�,�i|4T?��$��֋��︛]x�>!7���h!uP4���:�;�#X�x#1w���:U�u��]���Q�D�D��9�2�_ɼqIXW��.���po�!}A�XG��萦�;�cf���,�}F2�M
QDũă��efC��i�[5*l�}�?� �GNK�����q�;?W��_7uc\N1�I �a���ۼ��K�}�!S{����^�f��7�wv�����֝�&a ���Zv���[��.6������:j��xacX{��(�GRS�L��6�����zì��������V��;F���w��J����|��0� r�;�b���:���H�b�u;Gi��p&�)�ط+	!�`��:_3�/�{��I��ע�Id���A��k�����*�C^2��{f�ī�o2�,�p�#�9e�&;O������
i�ʬN$Dk��'�N�g�%���F2��B�ъ���=��0�ؐD��"$�>�Z�壟Ɇ�$�*S1�~�-n*3�b��q7
�q���������V��l�q"� ^5P�1I%���iF�%����*��Ch��qc���B��Jo:Ⱦ�m���7�0���v.VL��=�+!��� ��x5��ӏK^L6�%L����7� U%>�J��_dM5	�)���h�	����Vc�-F�Z˥�ܒ�18���uc��8Ft(�v�h�Ͽ�
���Ib��G����	2��;@��*��ތA��р��)�;n-)�&#MGk���󆵩E�w�!�ڹ���PO�[��t�R������$T�i��\E>{� _pP��IF��G4���X6��[�q>�φ�sU� 2����D�6�L�a ��77p�ԋR��>��6���a1����:�gD��&9<$R�]������B}�����[N*tXK��z�N�Z'��������i׽(J���$�)�w�;�