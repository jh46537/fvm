��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���q����f'����U�S-Կ���Q@B	�Pv�˖�(b���h\��4��9���6�)ʃ���������Vt۽�.0D�m�6D�R6��pQu)8cI�-�"��<���`
�qHKzǃ�=w-�@}	t�2nz�t[ޭ���l�cGl%��|�,�����n�����6B7���';��%a<(�9]��v���\�^u��IWO'�n+��%!�����X����t&��� ]w��I�Uņ��#�ۨ��9�O�"�SOu)�qZ�7Q��S�jS4h�dGf��J \z$�&syѮS63۸�
��'�oc��-�����^����A��uU�������S����_�䁕������s~~�O��u�����}�
o-���ћ0���5KEY��CxWD�r�Ovo?%��lSêKD�O��S���Kh�*z[bͷv��R����*r��$/����75�����}VFu�UK�뼖�����y>;�n�\�Tu��o*�i��]��C���,As�Y����m|�&�e��Ϗk.zn���8~t� ����X4� $lulq���$��	��5bjM�W�՟�­�����1�q�����*�R<�G���ԃ��}�D�9e2N
�z��M�L����Q�R�����g����S3��!��q �v�M��L�x���kD�c%��|P�z�|8]9=�n�e	i�M%�:��������E:Q�|�T�^��ū.�`fHn��i��w�s���D�.�]f���L$e���o4�Bo>ǁ�Hk�h�<[R ��r&���]�[4?��-�-aQ���T���M8�}�U���\��XIu���¼}	$M.�[�c�u
@O�ܜ��*y��/V��ZI�fỴ^����lsIm����J,�|��1�Ԛ��p�,nu��ם��&I,ax�k�{2y�8�� �B�'�*�2:�#2�w7
�-�]�~ۡ�GX��yu���gdr��Fl�>ܕoD$�$_kW0�Y��~��;�5p
�R��� &��@��N]��J=ә}Z��c�oc�Òhq�6E��m�,���`�R"%:|�Op�m.r�r�{VB�3T ,+_PA���7����l�<�y�Y�K�>9\d�(�ۼ㐷�Gm�ΰ��Y���i���xo�_�b|b�g���I�@���x��oP��]'��Jb�:+���-�@>�7w�:����:�BI_,0�+��"��(Z�T�%'�,���z��*�U��pШ�.��o���aŨ����,={��Vω�G4�3qĂR��?��r`ZL�*� {i��渼�R�H^>���| n�-��8��g�ܮ'�F�'�����&!�	�Wl��{B�:a�M΁�קX�����i}�����L�g�+k��˹��EsZ�Vƹ�	��- @S7�c�T�q'ͭ,��#J7���D�]��
�u]���y�`���f���`w�q��n@  Y-`kw�>6�1m)
�+�Ile�E6���	[E�TU"<*��}�������Fd�ן3T�T~��B�KX�8n<����6�`s*��Q7����+������Eq���/�5�N�D��З���LQ@��:�Z���,w�K��0ܮU��Kň�^<߁��k;�A�x<f�k�d&;�����&aS��e���C��ϗ�����Z튎�,�v	M�	ӱ��%��2�K��|z8���KR����P�O�-%�"l�J�i+�*va=��K��|�o��A��;�Ds��J�}>I��ϒ�V�K�"�ʾ���v��^Z�%���X9ǧ���|�ҍU9Q$�e�� o�nhQJ�Y&S�#�Q��ơ�F�O�-��>����"#�~�W�/ ���������1#O#L��6&'��Zx�WA����!v�^/���k�J}er'ؗ�AأC�ZR��O�0q=�O��q9�=��r��1��Bg6�ʅn0����>�H�ƿd�}Z5�rL��ν~O_}�,���vr-���P�r�V��Ĉ�O���+ZƓ?J�i�N6������[RV5���r�t�X�rK:����1�f6����'�A, ��jP^^�(���}L��US�H
����^�f���4J�Iܝqn��z��={�K�eL���i Y�l��͚�5uJx���x������:�"3��A��HQS��+���+�D��IGOѣ����T��+Z�3ʃ�yݓ40ÏK+��P=&@Il1v��ݔػ���T,�j1SGfQ�M�(9nji����o�eX,�{���cP��\΀Yą��w޴	Ԉ�~�'�U��O���8��=o1L�>�l����1Ο��M�c�|��XQ�+�tʟ���Yy�՜�۵c�E�hv;�xQ�zh1����&��D�UD�3����$�����-Y�S»F^�C��Y��ι�(�����B1��L��xU�oy,����HF�����1k���?���,/��m24�X�[��Æ]���CCi�A-X�ʽߐpDl�/k�c���	�ݗ���&�jP��m'(�}p�hu~�M2��p�F�A;�ߙw�=�a!�f�l�T�c�sN�9���{���������{?J�>�L��Tu<PV���ʬ&lD���SU�%�0;�}g�u�w������H]bQ����"��S�r:�8sL��'J�QI��;G�v�[^$�F����+KAHz�-q �\O��?�9����H-4H����4=U��̻��g���S*kr��ƨ������ ?�il���?X�L�b/rt^����u���'�Hw�^[['�):܏�R��t�r}�}�^r��5�-ZI����<��]J��)�^UJ��0���K���F�Ѭ
N��l	�n��֋
��󹳀'�� �5�*M+n���	`�ߋ��p����ģĎ�^hH�T�
�$V�O�O~�u'��1�찞p��by�٢��� [\xs�?[�P� �$�$>�z�=���]��p���d3��fE��Xx�np Ȁ>�JNx�ƞ�����yeU�d���诇	26j�2t�r�)�x��%�h�!X�_;�����5���|Dl�����1�5�]t�� �����/������:U�$Z<���"�XRB��޵������'�#
D�*�MvQ9��Bh�Y�¶I����zi�NB�8zJ"�e+B�*�c���%u"�_��K�(�'���疟���up�OZ�חH>H�@nA�x$^�ק��Z���7����
F��_0o��Jb�&���>��%�����";4�#%�g��!�7L5s
-����U�i���L���_1���?�!R�S��?>��h�ms�O�~	�p�