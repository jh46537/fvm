��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&+��^el햱\�9U\J8�nl���0�%PҪ�M���V?��� =��9��Z���x���qHtIC����*D6�qL<�@�:%���"��Im$�G	�a�_b~%'^��JP�x�֛��6�x����{�$Z�ca�����MU�&uږ�m�pS����8���I�n4JY�-�Rc�<�+=I%BY��P����P_�Z�H$j����""����q�}��,�|��=�M��!IËp��3�s�An�:�̙�8"ب��qږ;��9�ڬƫ&��uP��~D�|�q��/	-,5A߈:�~e�eV��������]�Pzn���3�6-��;���1�/1p�SꞀh3�	2�����H�괹��6��E����%	�d;��8u��uʗ���%��P@�&�P�*��ڰ���70I��:����
�����W�AcӰ(:��z���P�T�P�Yb�G �j��1vaK<�0k,Yឝ���o%Z��#�O�m]���R86,�)�j#лU�m�qEX�0���o7�����Ǹ0BZh�����^	'$����_���+�����bNp��%-o��kX��{^)��h�#'i��/���W��.�]@�;���[��ا[ۚ��1� b�~�1މ�Q]G^��݅��ɿL�<�$a9�7*ɠ��*Ti�l���<�h_NVD4�X2T�=���r������W�$Ƀ�k�=*��6�	G��j��.��|�5�)T�v��s�JNu�t�F�<����"�zU����s<�+;~��k��k�,��{�����"�,Hv9�$^�0g�Ԛw����$�&�{�Ǘ]kֻ���b�z/��̽K2�a�a<3ʠ�iї���t�+�,MΧb�!��.a�L x]�����^�fm��;��)�Q�Z�⡏�1
[�<r� ��`��K�Zw��o
����=����Qy A�1��LO�`s�uH@�#�6UO�ݧoQkS,���*i�r�\;�-v%9���'�p�a�U@��Y�G�guq�@q+?'O$|���E���a������5���_};>w����=�G��a�Mm#��+p�q�{����V&�����C�F�T�����|Ok:Sm���n�N�	�O�lN���|B����,�����r(<��6���(��
��f�
�J��p㻸!V�'丽 �}��g�Mw�!�v�����N48vD�ۼ}���,vI3{�xr�~.+n�)�������a�jtm����r��t�G��ɗl��_��W���SZO��5#��׿W#�:�&�=ۢ0���x9gz�8�H3]�l���ߐ˦Ƌ���1<����4�T8Tdz�'E�P'�j�d�R��U��=��w�.K�[�È���	j����5t����$t����W�8�[_Imt,v�sI50X0����e�B�8M�@��xVH3��>���w�r8�M�����Bꢱ��־�1��y�3�����RE8P�6t���k~}V;� ����	�8�	 � ��@觭���5���@��hT�K,'����\m%e�fl�����p����L2IĹ�l�O_
����ǚ�	�l�H	0�évH�,ob�v��?�A0�0Ji�D���q��3R�m�q?*��wqvgI-6>W�.�y�AS�Y"�Y9�F��C8\�F\���i��ɆF��8r���=K٩a(��zLP���pg������M�S^�D����Y]��x�=��+���C��D�F��8�>a������ZQ}8�yJ�W�JHx̎���`�x�a6��[R�@�.$(e�q�!5��ӀA�R8rph�yX|[��~��B}�։G�b��6�`D�=���%�������Ɩ�<o���Y��{YR�2�7� w`D��p�딱 +d���sۈo�#�;p��#[������K��}w%�p菜�ʴ�2i�X��HǾ4����Z�3Ey/a���孪����4.H�L<˝��:���}�i�Ð��������C�Z���+h��7�s y�����TmI|�J)��>I�.}Q9�%.:z�������,D���j5����X?��$̴�ؐ}���ԗ�!ȸ�o'"�,�#�C?j�����n	t�s��3��
�}��&�cq7��H�?�(�+ك�ڒ1 Ԧ}CՓ� !M�X����x����|*����ᒡ�����!�x��4^$O�iW��#�D���N{�Mmg�IG�W�%Ml�qQ�В��E���ϕw�(�s��{9� k���5zf���W:/a���?�g�����;�YO�p"�ao6����`���.� ���/��E9�'���|.�o�gi95?<���ٍ�K���Nv�wq#g�L��D@���ӳ��CϾ�Ӊml�~j��8��Vtr,�ƿ�����u�Ia�ӑn��� Y1�P��=��+�:,���