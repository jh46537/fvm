��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��V-�@m��Yx�W����A�.�ƋB8/dq�4z
��&�Lj��7(.n���{�֚�]C��e4F���7��7=5�G��m�L8��)�smھ"VJu�&�RCW�O�#~kP�_�u	�{!':/4c�� ���mP8��:��^��L�s�bH_I�L��Gv�\IBj!��f���jq�<���0*�)Q�������Ol<B���'�D~M%������v���K�>�(l�U��GdֻM<�ܙJ���	w����ǯ?����`�@p��U�6l�ۓ@̿	X�@�����i�M��@� �Q>T}n\���6��V�ZA�k�l�A���$`�0ѣM_>9�Z(��	`�� ɬ��t)K`����갘�B���81sO���QI9��@�<�sn�2$}y�
�;��o���C�*��ύ�r�&�m�j�P.��~�'/�}2���;g�rV .Ib0��y����\�۟�����t��S����lv���}�['Q�D'}���Oß�+	�D�&�=h�t���ܗY�y{6�!�7����#�(aGR�z����^}hF́����b�)+�#Um/�3T��Bwyc֐�jS"�����9W�U !����p�|N��1�h���?Ml�oB��W��ʚLz;$���4M���˻Vl�8�{�@ډÄ2J`�᧼��w����F����y�7uւ#��W�&#KУ$�;�L=��������٭���@���r�-W=3л��P|�N��풄�T���,��(��{
Ͳ��rɥ���q��n�����Y��I��&�C��b�Y�>}� "��II�,2���L,�5V@d�(?CK�-�u���>Qa��tz�&Lp\ʈ����ܑ��$�����!��5nV1X�s�"�1��N�5 0*���/���SL�(t�_G�x܁-���289'O4$<�S�^�V�����;[���F�ۃ?F��4��{��5Y�(�������/W�<q4��!�ٵ�>+�􀼰j�ty��n���;�_��H��a�;-2�0ԎY��t��D�`Ja��0�$��ѿ��q��!-�����8�G*%=�	gz��a��M������	�������K��G���T�"�����rRs�-�z)����F��W�@l�m�8B���v��	�;��,��z�d�!` �?����:T9�o2Иx�&�Z?���^��V�Vv��(0���a��ۘ߉�>DuI�)�Z@��@��������c_Hf��d����`6�<�!����;��v�ű3��`������"xvX��V�E�Bҥ��W��H"0>uEC��Ü�َ~<�����*�pյ�>o��ڶu�aU�Ku��J�'k�v4�U%�q�Vq�RB����Jި�~�?�"��� n[���7����t�5뿺C�ב��&��5��Jnw��L)S��i��<���Ԓt��~9��d3f���}jG���?�7(,!����-�d�����EOZ���k�*S���Yr
|܉}c�RﾳV�N{Xhc���~s�R�ɝ�;P����na@1���^������u��e7rg�E�F��LH�X9 ]^��y�e�W�.�����?�6P�XN@}����.�Ķ��y���h2��1So�H
������<�^H�v�p۫cά�i�X�Ox������ˠ�7Z�2�L���ɞ��^�5:0i���[�űQ�u���ˏ4I����X�mw�/�"�0e�)cW0)����#T�O_o������z���F��fu�:�)j�F���w�y\�u#rh+���^}T`�uΈu@ݠ�=�=��8�+G9&	�~������1�=�Ko9��{2�e����S����;W�hj
���n1�h%*�|�A/F^cS3i�H�~[��F~!+0����<���IV��Ǻ�A�I���-�eM�g*z���N���FJ�2�|���>�G\$Z��î�An��S��N�A��H��2?8�p�G�C���(�&(��z�/�$�.3�Aq:�^ժ����y���d^+P^�Ɨ�i��Q>+͚&���Q'Ad�%�PT��|f�'[����x��6n(y��j��p̰I��}?����.'co�hN0���ƃ�!�DM&j{�sM��=`�W!�f�J���E^����O�%p~Q��<!NƟ�����Ά2��?�gT�I/Y��Ryٶ�!���TZ�Vv��s��P+��-�"<�ze
o�8��hV^I�*S)��؉�'Y2�F��r1�f4t�K�ҭ����;G6�7�Z�ˆQ��۫	7AS�0�3ɩ�ȅ��	��b�ڏݙ#�;��ԣ� �� 1Y�.K���ݾl��6ܤ�7���Yx�3 J�f�;���֒�7�A���C9�x
��`����0Ȇ�����(�
�!oP�b�F4��Lt� N<0�i��m�J����Gk޸w(�c���P�4���� 6�r��Ve�	��nߩX���ٖz�⥝��D�.5�|�9��
&'Qì��E���P�5i�����A���:@��m���W��}O*&����U���.V������u7c�4K:�� ��Ȫ��m<��CW5��X�����({i�|��j������ ��K��k�TVl$�Uz%�͌pl��4�O�g��d
m�O�aX���n�M��uN?�������V�k�����.�r�����
����I�5Վ��쨪��4��ԃ�cW�[�L O��o�?�V�����c����`%Y��3
��k��{�K<3�|�HB��~d�AZ�(F��CL��_U/z1�n+/R@��0Ѹqc��	>�Gut Q�{{�ҁ?<�Cq0���Ov��G-�q�|�x 4L��|'W�m&2�b���������f��m&2�$��afX������fg��֌�$"���p�D�c��u`�^ƀ����VEm,i�'�rD����v��PZ4&�wCRxMl;��즖�၉Bsr���b�j�%�W��f�`��S5[�NS��m���;|�4G�x���΃��h���gu��r�����C?��ƶ�u�~�*l��N���ă�̬��'�[���Ӄ��l��w���A.5���o��u�;J/�egV#�;��#��T���]�+�dW~l�����"(-^Uc��.�)��:����]@W��M�H�B�D�MY���0�n�I�I��Ɠ/i ��7�R�������a�a]|�����S���|3wPJQê��k��_!+`��� J*�qoȫ쾝/��<M�{fN-�Z�B��"��eH�i�-5�t�z���]?��a��6<F�t�Pⱊuۿ��Mn��yi1,v���̗��c������g��O���D�L\�23����Y�9͖���[Vz����^�5�zdߤ2��.%~8Ah��4�5��Ȱ�@;�7S1$ĀI�Ȗ�k৔����)e���>%����31�h�^�r�
���#qEܾA]�p��}�`��}���3[���WT�R� ͽLr���U�q�pq�`��q���,�j@O{==,p�$N�_<���&���,���f��DM�u�8��|�'cڔ�ͬ��� t���U7�l�ω����A��T_Ll�>�\&nU4����7�א	^Q͸�f/����~C����/4N�! ��19���s���4e����Я��r ��$x�!�{���V	�B�������Dn^j_�qxbT	������}١i;��Ĳ���e	7�w�J���J�̾i�eD�lW� H��N���C��**1~~mGLt�%�����m�M�vռp����`6a}0І@��7\�L�����l�rǙ`տ}��� b�-�	�P_ Uw\����:.]ʭlBƑ��ɚ�Ԋ"n���ԝq�RoÉL�q� O.S۾e�+<�h�{fF�xU�4���r��E�.�c�o/&��Z��+G�L�ǑblՄ~�d�S7���-��4��������a87YA�/4=�5Jv}�I�9k\p㞻�Ƙ�x Q�҆���Ѱ:��mO��7�E����MO��F��rS�F�~ӏ7N��]i����W�K�	DY����3I�(�6��/�,�$��nv�@9��Z��az�[�͹ZNzk�+y�웂c��:�d�I"rj>�}w��'�i���K n`{)~^�5�+&
�Tƍ�zm\5�ME��j���Ǭ�����e�?xP(��`ÚkT,L�Ys"���u�6��`՞�k虋ar=w��CT7���E��U`�p�AdZ�U��~������4ʻ�S��L�E\ȾoJ`J��T�ø�N=�u�=�sJ2qMu[����{�� j~�baZF����xS�Eibmy�Ta�� ��:'%�۪��16'iW�(?�	1����h9�\��~Մ�3�<��Uٜ������G�e�6*W)�ݫO�5��h�里v�j�r�+ ��&v��~� �M<QD�*F��*a��\&�8!�)!
�}r��c( �xpQ���Hs���"V���d;��� ���XN
��E�������Q|���5so��i�e>�nb����o�$�@��l��k���_G�G)~����A�8�;D@|1�e/e�-p�0c�昌Cz�2�MF���?m!YV��Tgx#����Do$U�&i��B�\3W�?�Ǟ�3�ɤ�=�6�s61�G��}�x���o�3i�o?w�u��N��	�̽�����mZQƬ>�JI�[�nr��C0;:L�4�t�~+i�2�HlC�����G˲�y(�2�c�H���v���()�L3�"ۥ5+��#�}"^9y^�9{�]raW=f �v{��!�Kߑ��u�
�"����7Ƭ� �Z�H,R��LN�f>ވ�YY�hI������(&J��:W՟���3d�|U�j�ʙ�������d��	�S� ����]��x�Fǝ�:�.�W�+��y;R�TT3"X�%�z�u�@}�*�O�1\��y��0���jw����6��S��?n�2�l淋t�m�Y���qSn�A��Z�'t�W��)�Ҹ�{q�Wn���fGH��$6kd==�@ �Z�����Q��H�|s�I��"���������W����`"�/BV;����ř?����ӥ�=p�r/�_��hzB��K�ڊ����f3)����~ .xT�H>�~a��<b��T	U����Z��[�cFZ3늹�?.���:�m����Y��P�*1�~�M����[?��M����Β��ױ��zp�i���7.��Y/�,!5%C��c�ĘAk��ė�G;�dD�f�4η��a���t�g�+SLVs��n@k����Q}T���*l���㇈��'���j��F�I/hRo~�N�� 4@�o��������/R���wR� -H�ȸ��٩͗v9U�~���s���D���Z-��z�r�<!%���@���	�	e�x����Sm )�@�T��w�u�>�������]� ���f;��((������O2���t�CI������V����Z��A��y�5O{�Ipr�5���pLD�N<��K ��Ɛ>3���_<���(ҋ��N}L��D�?=PN<��4H��[Z �{=L�!T�i�����bn�ey��W��j�
9��
�%d�`ބ����)[v�d��on�}���y�qė������3����ĝR�]�w
�m|��^凜��{��ŢB�jxo%�;-H�|u�F�R�(�������.�!�j�:��9F��e}�<p}�E�d���HN;=��˅�[�B�t��v�L�|�n��uמŸ"d�A�kƅ?��g ���]t&P�_	���'�]M��J�hfc���X&pj#��a1z(���7��Alg��Ab�l������H5[\��:�;�W]9��O�oyW9�tz,�D/.�Y��u�P�T�9@��ZD�U�	7����P.���v�(��	�,�/x�+i�ao+ݾ�W���%W���ȗZH0U\���[�` 7L_�,p#u��,VSx�}ٙ������ZVY�?�zhQ�d	���0�%V/�����4t -���5��qy}�	��?�9�I,-�����N�QPwp��A�/��x��^j��t#����g� b��c���~��$~�'2��X�(M��U�}�gmh�j8�/QW<�u(����S�.�� �09��A4��~���~춹��d����!�7�m*�9��W�]�W��������tN/cW&Yk���Yv��VKŠ)�IڐÀk(�d-�|r�䒨�F��+k��a�XΩդ%�J��ԁf��|���NI�u�/5�֒Oz�l4��o���q�&��[wk�A�.?[I�Jk�����W�JX�2 ��M����=��r�����b��¢�$q�C{��m�a>s�c�.���b<|�� ����%l~
�r�cN뭐Dn�o�lHr
�u�0 U�i�0Zw���m2�]pל�	�ݭ�$)����v�X]�'�~h�d�y��K_݌L����x��L}��ۨ��%[j�o�>�-��U�U�≡r��<d���x���+,��դ�c�ݞ^^�{�ħ��}.��{���#���Y��Q�{��q��`�,?㗤�l���Y��?���2��v���c���G��+y��Ʃ27�����&X�"��Z�z�]b��0/jBD|bVQ��W��H�2D���q���T��Ȑ�	Ud���4�فp�-��-�F�le�/�Z�q|g�趟��n�i�ot}�5<ya����0��h�jv�#��՘C3׷ �o�}��вh8�v;������ȷ����ܤ�
�rZ(aɘ#��ۆ1�����Erm�.�>#1�ZR�<(߬,k�8L�,A�I��8��G�;;q��d�S6>��qCJ`z�r��7y�����e��ӛ�����Z83,!m�w�8��YKU��m˃��C�pW%7�b:ݮE�S��V��)T9����C�L z��Z��KL��%�U���')�T��Q�p���)�l�.�