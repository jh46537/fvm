��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�+�3����C�vmػ0ɋA�
n�7v�%6oj����T7?�Pc<+;F�]A�`��ӫo���\{�DR�^�k��W~��^ U�RS}n�J�ThiR#�ﬞ�/_X�:E�P�5?y��QNB��Kp���{:���_2�t��8lf����qwm������.�`�*9��rpf��,N^Z�$桷%R�y�)(� k�$� ��uz{�?�K|�jr��O��mL�QY�vR|y�#e7WX2<%�_���F̑tVҨ�1O�0���xS��=�^�e�b�u���޸)1��*���!	>�3�W6��E�Q�4���(a�1���.{���Bz� /�h�@��u���x����^�D$���VW8�8���p�U�|A�� P~��f���)oI� 싯��G���2���4��$,�D��Y�>[��9�!Y�݀��z��3���X4A͓����B����,�m�}k�I����s;-v�g�;�,��k/�ʡ�Ǚ�W��T�-�\���]Ȅ�x����+Y+%�AmF7��Γ���A�4�4�Mx��+�A�b;���ãD�8��>^��8q��7������I-gX�	�rܶ�r�^7#itL�����IU���,/��E)#5&�>�Wq`�|a��8b��B,An�pr�PQ�H�	ȱ����~�h��{�i���}+�	���<��YkĩG��wf�@&7��U\�I;<���*Q���囅�F��V�N��T.[u�p�G6�uZ\�)k�lNY�S�Q��rK���R���B&A���ƫ��]U�}:E�䩡3�� ���l�wF� l�o~Z�C	^��^?W����%�\��,6M�Ma�H}Ӣ���̉OK�i�v�b�&̇���`4u�ɹ�s}�m4u�����5���?�7eG���
<�q�h��u��L9_q}H�Me#�R=�Ϙ�J�נ�3�C�{�d�`����e��7�&i�A�="f���=B�4%o1|2���!��]�g�k�Zۥ�'0$���u爺>��́2 ؙ��:���ha�C��a�o�_��]��26	s�94Qu�9̌8�Jk�_̫Z�\z=����@�#��r�6�92
�qh�H�U��8�1�g`|9����
m�[|8����qx�	�Q���<�gjQ?�z�~ep�WB��c52e�vF��?��3��.�8i�-�́Rۜ�؟�=A�j������j���z�/A�EmK}�Q++�^������ 3[�oɳ��6i���F3Q��A���쀻>�}ީ�ط���1�/7�[���@d6J�^�Qo����ֵ��j}+6�j��Q�'�9��KƆ7QYXOn�lň�P0���	����%��j�1� ���r�>:	2��9�W�!>֓���d�{ב.  9����4����)�̛��'�Dղl�qZ�Vx�������,$�ӳZ����!������{�*�A���D�*tȋ5�8���p0��)\bG�ܨ0a�B��b8�l��YH���m��b ÕJD���S��1�S ��Y"F8۴�P�������nC&PQ��$�*eL��`0��� qW,���&��J婌<�O��_w�b��<1�	Ք^����:�F �i�|h�W��p ��<M�;T�bCQ�p�޽��Q��0kh7�,�[�M��0n	��"�.��o����?���>X��)� ���-� |�'
�6h��Y�[I=N��gZQ\�����v����Ҭߍ;��2p�� �W7�nH��������p�cPa�Y.��Z�-k(E��w*\��(�::3S�bJU�_����Bt��r%��u>���]����S��@roy�4[Y(��ڡm��p+zh�ɀ)D:5o�7�Z�&�?��54���>w��`(���䟗>^�����v[p~Ұ �]�"J%g��3�q���9G��O�B�[6�>�����������U$Ve����s�s��U���9������U�p�^s����
�[��z��5AҐ71�`�勨����|�qk�������|P5 �D|�������2��0b���i'oI$Ɖ6��/P��5����Fj�oYJ�öj4y�Z�CJ-Ʉi�-�e߿��l,�Mi�g6(�j6�0ъ�W�]�D)���|e!�h�[��W�~� ?��b4(��\?}f�ge����Z�c���C�*�=���=9ݮ��i����b
���,Ǒ|�53��p�n.f�?n:۔%��GƤ��8v�y�$�
ڂ�#��8�oxuA<��en��#���LM5���LX�{04�ì?����(6}��nnKъ��a�X`��%{J�c���P4�Ek���}�0�%� ��ճ]-�\�L�dG������7t�"}�uis�#X�ʊ��������#��,�6F��VQ1�J�J�
��c�\v)k�b1Ȋ��a����c�}�ێ��l��{���[�ӢU�k��&�7�<���{F�0�����v��\��4)��F&G�Eq��!�J0�[(�Hd�E�^Hq|8��-Ơy[��A=�!��(��K�[\��h|�cI`�+�[����F�oD�$�;�=���,�s�c�蟿2=0�^�I���#�����O��k<�ɜ$��-�[�ɵF�v����@��c�R�J�0����3�e�nװ^>ߨV�e��@Pd�CI���BVp��q�/
��g�B6���)B��̭K�_�>η2=JI~sUH��O�"����w�V�pJ"x�M��� �*�1���*nl����|t�?ǐ!�M`)@-��N�����(�>�2�h��}���Y*�\�?%����v/���T#�F��9&��P��q2�<��vn��e)afn9L�Y��r�Q�������8;�-;�So�q3�ϴ:l���b��hC$���ܑJp���H� /�����e:&>b�s�qk��!x<'��� �(:<�I�{��R����s=)jxiO�bȔ}6!rB��nv���UIQ[���/�mB��Fj֖������g�K�ng�ꌒ��H3z=6ǈYO䚗]���q�сK�FQ�Z܏��T�"�=�ۈ����v
G����b�:t2��E��?���;o2�1�������v����*��t���']��d��z�.�+�f�(��h�_C�]�f���4Ӂ�|3�����`\}�3]I�S(�(�3���ЗȗBxL�$�
�5[#�tu1��ɒ"�ez0�'���ގ�@�L!� ���'~C*Ϫs�&���z/��M[�콭����B����{����g������
@ �������� �o��ī%�;��c3+<aZ�J�����ѯ�l�"�[�S��P�*ɐ��Fb��$hm���8}_>B�p���N56F�&R�7�rf_�s"�2n<s�BPed��8��^���鋱2?n%�Gq�<
�߸��xX�����q�I�� -��82]��K��J��_�y�t"{P{9Ӽ����1�,F�@E���|y)p�l��n��d���z�/�vAnN
�UI^�3t]X36Z� �|`��]'��Ng���%�*���������C (.	��^B�,wӸ�>��ǫ$Z?'��Exd���l���3UX+�p6;�� H�B�'�"3.�1��%�V��uk|�Bm@�p�'����R��j9����6L�t�&v�>2����s-�@tm���OB��j�!8�oe=����U"@3�nv�������rr�8$�lҤ�p�%���o�"e3O`�����h�NO�Rj躵�H���8�*$8FCU��&x�=_	�@�f����3p��$��x3��.��#1$�u%�/74R:7$��z�*��o=��m�̣�@��#
�Ѷ�=G��j�A)�8��Mq�k��7� �h�=���W�\Ot����Jې���H��`�L#���Ӣ) {��TR����م蟮����F��u3�$�
1�P�?{[_�p�"�D�e _75�Q�
d:�y��\�$�GV�{�D���/��A ���x�d�I͛Luɀ�'f��H������$]�y��
�k��
v�~�W�)�E]��^Hj�qRqb�,�D���<�=��-��,`G����ך���ϣ[���u���cs��k4漒@�?A����9���5n�u�
�$�q�{k��J�����2�Α͛���=�ʵ�yC~ł뱒�J�����	�4�����+�ɥt�~VO|����"����F�at�Y�y:��^"�yVo*�@xܐAr��!(��5��է��O��O�:H��H�����ʳ�a�|APhr��,t���FV1B_q"V�O/�����>ǆf�9UF�4�	z�Eg�YGAS�ݠ��J�HY�� �3�E�=�f�2-�{�����S����	6��2>�4�&�kAĐq 4�##!����Zze���TySG	�G{�*��b����q,�M���B�{$`a7�Ҕ���=�FZ2ѫY���M;%���a��:�횸)���U>4�E��Ϡ��$����U�]�kd�v�-3v������{y�6�nw�Y-K�Y����� "j�5�O�\�}�(�����(@���y�z�������� �T��
�+!y�@��&�o���bv8�6�;x�U��/�[����ʺ��I6�.T�r�}m$��`���FSo��������E�ƔBU�=���>�7�as����l���\�a����M#�|@����E0�R�8�ʹ�y��[�|��P�m�aܶ1�i`	�%k����COB���m�V"�a�yM�v�Z>M�d�&�M%�;� �s�!��׋L���	�2����kE8@-0��i�Ϫۨ �K�-`�YF�������O\�F@	i�ۦo�S��!x;W�'������&$��w�^|�<!�/�RAׂ̕��Q9:B#RV��/?qz��o�F�:��1�m �J�X�� �〨�"bfТ�g���s��il��ɍp�4�q;�ؤ����b»���U��\��,,	+l�O��4�qfz�Y�5����A*���d�o{�)ϯb}Ca�>g͔5�-�X�wo�-�e��m�3s�uQѝ��R�H�]��</p*W��f)�����m�	B/�5�xm枵']&���+ZIʽXaY�/���M��0��id<U�ԗX��V�yT�M`����3�Y��hk�25���p�ՠ	�0����(���*�M�n�"��"i�T��5�y�b	�>ȇ�S_��A���m� ��n]N�9���?`8�4���Z��,k�rV�\i"
�n��-M�g�������*ؤ[LWOآ��@"�Y����q�-�u�xtAe��Ј�b� 4����|ؾ�/���ٯA��-`vU�F�s��jqW["b�Qt�������SD[�{�}�y�6�"��y�c����E� Fs�n��?�})ʖi�U�
�>9�h��R�;��>9����*6����hkoޫ`�$ƪ��d��P��q�1������{�_�����Ig.���4�đW���[���['��k���eO�"}>E�>߽M �9�ڂ�-�($��:��P��t�q�-����=r��,O���'k�&ٍ=����3���J��E[Z(� qT7Y�~���t�C��F`������*��cvOO���P��^�76�XO�]�|:�4RҨ̿�a������f�dV�G��_�h����,� on�LbR�����=O�X��Aa8mjh�b��p��_�k��Ĳ�I} �K�X�-�bq��ߛ�Af�՚�z�x��U��
��
�흞����o�{�i�iЋ���.,�$�������0v����U���<0J���dr�l���:,�q���PH��Y��K�r�T�ӏՄw��]M�́=�TǏ�
�,��*?�J�����;=qp8�{p���w�&�H!�օrdGK�a���bi�6Fn1�r]#ټv�c	g�&J�*VCa9�h7F��B�<Y'�j�pP��2 ����.�j}��~[<DQAK{�}Z�p1��h�g�:��� �d�'#-+�mx/KJ����1񳋻1�^GP�HNښn��� ָs�:c?�����{F���)��$��ơ��^�+���������|^�wLU���r��@�==�t�VP.��r�ƽ��Ӿ��MH)��/�̬�ׅ`�fr��]�	\ �Px�J��®W���q���dN�ǩ�R��=z��LjB|���e8m�bx0�b��(:�P���#[��Y���i��+v�Tc��߂*�G�����8wK�F���k�Z�Oߧ�>I�l��nĺ�;A�}.%E�ַ�$(@��OK��c�zk���V�$�I3ՠ��MT��Q���ҹ�أ���4���N$,��(�������t�H,<���s�U>r�ٴ[m���֖/�b�c���@�9Vt�i$s��\���/|`���3��	��5;�9��P���FgD�=(��J>	��p��Ȇ���B�A����ݽ4n���p2�a�%NxJ�L�.�sI��@� `�0#�Q�&����$�0����˾���u0Vi����Ճ�����3�5��<0��N@/�a��r!X�+٭�,R�$
�b�
b8ZME���+2�g���k>'����q��F�3����*2��|��&$pޙ �M��\��^��� ]�%궭��F���9�#�\�­��f�]+�Z�� ���ܩ=��H��L�D��l��x�;)�z��`�����l��82�Al�2w����(�C�p:�����8^<� ^q5��Qo�����.go�f�10����
�Y���W<
�Y.�Z�ZO���@HW���@ݝ85�c�J��qW�΁�!�a�z�v��둌�DZMV�k�{��ϭ����I�4mއ���K��u��Ħ����^�;��ބ��>@|k���L������r\�Ќ���=��)�q� Ý��F��>���B��9}b�$�3�P\�PY;������[K��<V�}ըX~`���l9F�+���ص��j[��g�4��w�\12��`�[�c��}R7O��p%��5y��U\�����u������v�lh&cވ��$#�})COj�k�-�k_�b���4>���e�Z�P����wY.����[�j�C,�k�9n�ǲl��.��9���6#s�#�k��<D|���]��m�ŕ{6���8��s���Å� SD"���H�{M����~B]�l;�'a,O�h]���[����j���B!�t�F5C�SS.>��>P��	8@�q*A&&��ry��S��!�~�5�"�YN�LI
#�hm�J@#� yuL�%�c�9��ț�<�RP��0_�Y�ӵ3AkB8�z�k6Q����k1�?����L��M,hΘ��*��;�^�H��Bϊ5}<c�K������vFפM{�m�����T>��.���T�ಽ�����W߅� SȎk���;�jZ���kj���0�SH"��[s��)�neR��ȃ���<��x*�kW��v{�1�Y��D�Al���wc�F-�����XF� ߑP1j��\/�����@!��M?�35V�p���D^\���|���˘5���ţ����\��b�"���3��FZ
�<�����@�&�w�)r�ߟ����EU$���5P��>r�GԾ�C�U�/W�d@`{�:��+�<�h)��FY���ܵ��g�P������Bi�v��p!��nwJ :ld)EoMrq������
tin�T�uoN=�4��DB�/��f_,�~��R���(���JYI�+�*���/��~����WEΠu� u�3�����8-k�!�GD�������̆��1ʏ�g7'�m�bKL䆢Y�,��:�C]>�#n��m�P�ч}���5��Mj9����Ўf��+�N��෾�qy�SvZ[�Y��l�r�	�TT`�zU���%��y��CQ�E�]����(�uh(6���5X�K؊m�G�����I���2P�tx^x���]�8>\��p��ꕢ9��A�M���KT{�$����sL�]���E�֐N�Z����j"߽k#�J#��*c8v�=D�˳��	+�q�_z���V?�5O�m�%	�<��c>��ǋ}�mcX�(ӏT�.M"qb� �@�`b%v�D�[eh�Q�ԋ������G�W����κ�mD034#S�"ق�7ﷱ���s���{7��8:=L�'��@��үC~�l�����g(���_S��;{�UoN���_�	�V���O/�-�W��_q�u�����Ʉ(��+�zY˅�<��"�G�o�Ѱ���~e�Ȭ_^�c��X�>w#Y���!�2D��2�#�hܠ����u޻�Bp��_.���I�9hI����7!L�.i,���0�W�_ŧ�m@#�h���z�UTq��q��$
�=��pn���:9}�z����J���ʟn�@$�P��?�k�ۈ�.W5fǳGiЫ߂M�z��]p�Sa�AK�=J"�9L�!����f�7���F����"���;�e�M˔§��F)V	���:���8�� 5�5��{��4]�$zJEz�SI7�u�9�y5�&�F�S&��w����53��pT6f������.���0,7��ӨK���۫;����t.�Z��'�	����	1K,jY�͑@��˩	��4����Q��YɄ�6��0�zi��r�q�_�mW�)��!��_�Uv�;?*�̻"�cW��j��G��qJ�R��~bc](��צ!Z��O��Ǣ�`��$4��\nIg����(��f��&�l�l�g��g�DS�Q(�dx=�*v� �k^�P[y�����0s'�poY�{�eO�����\��~�6\���Fw��	��3z������}��_T(�)s��va9�:@���ꤶ���c#������S3�{e_��(�������`�rL��Zė[�j[\a��%�"a��ɠ��ʮ3Omge�}��,l+��)o��֝������e�8;=�gQCj�8���\[�������rAvihW���)�uў"^�#�~Gb�8T ��F!��`,ؽ�/��AkG�0u-.��������M��K���n�%S�%=.�~�O�L�fga�.�|�u&W�xp՝:��q.a	�9À���ecHP�g�ܻ��@�ϛ.�٬���>*dc����F�@��� 0=�Tx�^�~�A��B ۲�k@0�~G9�2f��)�i�<�a��{���M�\@C���\ճ�L-�M��Z�ޓ�/��Pq���t5�� �/�>�-V>腑��g[�l����K�V�+Cv͜E�+NY�#&�@��qi)*�?�6�����gI��e�}�/^О�%O,r�������D��AO ��n�������2�߾�q�Vv�z�J�4�ꦣw*��V����?�2[�AL��ds�82���D�;��>�0|�f'��׃���B�($I������	�u8�6���H�L��6y�_�y'���R�����U�NM�]ݼ�ɭS0��e9E<\�N�$z6�/�4��7��������1A!�:x�"o;����K2O���2�ә,;7W���:rW�w�wr�9�p��Q�贆��zb�,�����c3����o�B'2���F`lLȒs�O�Gp ��8[���0��0�]wg�9]�G6�Řo�c�>^�oO��Joͨ.	9��_<�5�/4u��v�?���J�S��ցx�j�Ɏm� ���'ye�@���Rj����1�<��3!G����x��m8}�_��C�z_3Ɂ	PK�7����;	�_�u�
v��E�����ġ|�fj�Z���/�Mb�5v8vL����<W��\�!�TYLg�n�浕e9I���F�0����Ap��U�J��jň�䏖��A�G��[�@gHG5o���Eb0O�S���q�iv�*�s��h��u���]J�ͱ��)�P���1�(��S̢����P��{�Z�u��}�b��X�Ө ��� ���ُ�OR�P��	������g(o�l��1�4~
�������E���$��-�V�dK��v���k�4�6��ծ^�)��񙃰d��6�w�@�w�,�D[�p±+'4Ǖc�f.°kT�g�GF�w� ��Y=_���r�;�S�q,y���6/e�v���\ex-��4W�����e2�}���,~ȫ{�� ����ո��B�h`�ȽS����/�I�s�9O�'r8�z�(�~�i{�X7�Y��5��1�*��'1m��}��*p�ms�'/������y���LOm��s���j���i�05H���rM��/7r����VE�I�p�$�Z��cE��T�N�I�%ꗁ+&����Kc!�F��v}����cT���X��3˹��k+sgɄ��h�p�B�������f�'F�c_�7�z�!ijQ�2�j"p�c��1_)�-���B8'2���Q���MoI-���8bs*����z�˫�m�����B0�t`��/I�_&�x�iKQ'#�{C%L�
V���W��gw�������������񝲴�d&�j5;��Z�#
�,��*����>!B���g�$� ݮ�ʆ/�Йj@C�u9���Z<X��@�@*X�	��Iլ�b{*��7�F\�'tU
j	��$]����7�Hd���7�ID��\r���W�[�׽y$&�͓zdp�y�/&C<�pD*�Ȥ�v���Igp�`�M^]��&[n�T�B�ị�eؽe��e�c#���?:����b���P%5�0�0���e��d�R.�P��wg��z��J�:��y c���Zwil�	�T#�/ˤ
�X������b�>I�(PMjpjS2�Q�7�+b�{<��s�U����K�,[�&X[@�(�Wbe����}����h�XG���g������ՑA��(J��U�uc�?]A��ֿ�c#�}���q�����
ή���No�oؒ ��/%���ޫ�Wt}��PmmD��+\��u����3Q4}�����a�K �XtN j]�[�{��c��������M��������v���b�[q�Q*�u�RxN>CYd�RɴzxxJ�pA���`B��=�ֆ[r������m
�Ү݉���m�N����伭�Lr�����YT�`��n9���O
�������1G@�Svv���H�\&�E�T�hd��pX+;uK�2X��T�����6}�y�bSC&��~�y<͍�(�F߸(�c�6"�p�h���7�{�Ym�RZժ4!ʷ���z�����5�r`��̶m�F�0�����E$^�t���Tz�>�����\����}gXʠ�cG@�����ܨ��`+�O�+����۔��0�Z[�f�!ި�?jS� 7\���#= d�����rD,P��}{4A{,���b��~ٮ-<�sLH~޷�boEb�
Dikˏ.�`^����5z� �������  ƌ'V���$�P�*>�N�ظ�pr@�5���K�Jmy/��4����p���w.��>�����o\zw�_�&��o�Ӕg�h�p�2��i�P6�I�5�<́NH��'��	�̐���J����➞��91�}�%�|�_Fb��ޱ�t5E^)+!�ƽ=����oj{#�e�8�����J9hl�8��k��J6�����g�J�����G0��``�S�q��AFfh�͒JT0��+l�o��� �;ݠd�'v7:Bm]���!��8C:����w�2!!�բ����3�D*���9�*հU\�S�؈����|��g���vu>�4���V�]����J�OJ��ct N��@G�tr1N��y�!��_�6����-���3�vO�m<E�	*A-y=t ���o���$�Ǒ�j�w/�8��2�y���յM 7ַ~��\ԋJ!t����T<�Y��r\i�s���)�q��������� /Ҳ�H��_ F������֎0ld��P�̣�BM-�>a{�(yL����w���)>���0H�NX���H*�����Z�g_zk�G���?����2�_�Y�H�k0ms�8�K	,L�P���;E���R��,�uI��M>4�1|UD��R6�Oōz���7��-c�_�D��˫���t��9��N�x�Xk%�=��e���M᷿��ׅI����}Ω�)n˟�LR�Dtɓ������0�]�����k�s��+D�)��
q�(�|��FLF4�DS�AI"���j�����;�`@%�E+."�-6'ɴ���w��]��x�/�:*�42�bػ�ڶ�>�ƌ'�RA�>�W�K�M#�*��da���ݛ$#��*� �����Eֺ,
[Dv��!q����0s.3�h�8|�Q�WH�J��l:���ƯFN�FbP�@�x�r�&��mp��b�n�<�ʎ,)�}��J生R���!Ǥ�)��Jco:�F��!�c.#[�L�� =Q"���7שh%���ugދ�������v��~�SC�gP�i}'��O{K��LY�-�6�b�-A�l?�oo�L��l#�/�5�Mj����g��y�Qq :A>_o/�T�g�o2�yy=)�CW�����:�a
Z�W��9�mQ���r �s�*��i�@����geZ��G���1��J�"��^.f��8]�2�G��K�8���7�ig�i�x�Β�pE��� ����B�S<3q�>R���zA=Z&�ŏ� %������nfJ6�g�1�ê	��SX��	��w�1�u��+W���z���b��[9�9�QzG(�;���G�xj���1��r��`.9lf��Q��v���(���.��迎e�hkن?�+s���a��TJ}���m(��E����۟+ ۑ�XÛ�T;��[<��;Zp;��D�I,`�v�b�ޕ������È�Vc�o�p�=-����q&��40�V��Q���"�9%�D��m��E�wp}�k�4����᠍@.?��jy��9�����<c �o��3ϙ]o���@!��\��Ƃ�˘e%��bf��n��Oc��\U_k���Ŭ�r�Ǻ�j��l��t}4G���!��w^c={p�Z�AX5R�_U�!�D������� ���F�>��QI�����UR���;��i~�T����� ���<��o��h��ȲC�BRޗ��<"��8k|/w��_w�n	�	�ࡻ�ċy'��t��ZX~��Z$�=l�50�p���� S�u�\OjeW�u��a���1+B�"rߍ���3��I��������� �d�:yH�%�Zp�8�B$H�w���:te�gc�����&�*�=�95��u(b�:��7v�Ԧ��P]���RX�A���.L ��?S�ߺ�zV�e~�,�AwDq״V�����u@��N��f�@)�#��#f�M"�7�o� X����ܾ��ɉ�S�3�F��g;%���q���y���{���xOS:������Z��/[�4�I��s��9��|8����?�mE�
�pL�ۡx���uN��
���h��R�W�*H�t{�h@���fR�d<:�� �iq�u���}�{���^a?���GF�1Y�0��-y�l���"m߲�]a�B�,���� ��ݢJȭ��TnQ��;��8�j�G���F�Z���I������ԩ�8�:�W#��QaG����g���ʣ��na;���f�p��F'����#��qD?sNC%�szf����4�@�V�'V�z�`�a�"���Kvi�����|�[��0�����z�`P��Z�M��٦`���~�q�x��PY�Ҹސ�=����Y�y�G�>�l�ao����[�ZG^�.��	\��
�ܟ��8�J��ws�jA5��h��QDw�v�5�q�k���bㄒ����w܈NO�)�뻆^�S�]Ϸ+�<;ԗp��n"���΅ˏ.z�1�A1��1����k����y����,��c�������8u���{���B�0Se�;�$w�o4�4��תj����A�(��g�P������HUv���JB���!�cK�q���"��5&{;Ͱ�$��8��қC�@�I��<�Y�j ӊO8[y���D'?�L�7�~&�)��BB�o�H!T�LB�X�.Ǌe$��H��rs���D6dsk6�PGaB�1u������91���\���Wԋ�^����D�y�£<n�{Q�P��(:Taw���/��Q�𦪾���b ����3�Q�i^n*�P�m����!}]�χ2_��?JAX��T���ܤ���:����ġ��bݔ?��w%��9(��=e�L�爖x���K�v!�l�p��7�5��]��<����{[�C�nMo�#��=�����H4�a2��k-@�޿?�QVyV[7p4���
q��b�@���>%���6�+�.��f�U�����@��Ģ��hew�D�D��x�߲��q:=_�U��g� Fp�����L�WB����Hݐ��9�ג7]#��;����5��P��V��(u����]UsS�b��2\���.y�5��+�0ru�ִ��K9��|x�}k��Nm}���O4Cȉ-�f�U�;�B/C�n���`C�&z�	s"���y"�I�<�i2:�����f7O���0,N�B���(���>ؑ}��ӀRGU�[�	R{
�>t�Q筯Qj|���{$0�s����ࠆ�N�& Xu|pU���_`up�b��WN(��t��iu�~<h�!�옛Ǚq���k�c���֬D���FVZw�8#��}�c��Ȕb¬rG�����O������^�k�T�K]E��i>�"��t(3�g�2Z#:&���{tO�s�R��bc�����矽m�����uRj ��e��}=#�a��+DOAO:C�]- �M<۸�cd���i�r���N&@==B���r��!���@:�YV@@a��=�`�*�afߙ￪%��RYi����%�s�S�������bs2᧌�3�C.5*�m���S�7��ԋz�~2K�o�K�a�Em�"�+3������-f�j�!DB��d���j��e�� t.k� ���Ɠ�k�f�#Ge
q5)3���SEk����,�U��o�U���������q�Jj$�xFkD�,�z�DA��/8�m�z�޶k�A�w�e� 3��G��i@�o~m�> ����b˂��R�����ox��N-��%Z�Y�D@�n�ޢ���#��]�D�=]��J��Ǳj�h�j�>I��p��S:3�o�]�~�W�?�lK�2�9��mԷ-�\mL_�'��P��~�g���(�l���+��"Jc/��*A�%�����W��[�` .��3���c��X�Q]���h�o�'B�׭�@v�k������#;� w�ԗ�OJ�DF�Pb�����}������Nt�DDQ��1(o�u�M�����$�u�#��,��b��O��$^~z�?��NB�L�k
}�&CF�ڦ���q��(l-$��*Ԋ.�E'G���ka�.�V~���m���̦^����(�wX�Y��Xv���2���k�~*O��Z<�"��������j��R׭�nPp�~q��L��˩��uPy~���v���b�6�י��+�������6�Wp�*�;񶴺��DL"���U�I�ӥ��D���A��0��Y����)gf A�8�1�<�)���ɣ(f�d�^���,�f��(b�`9Ĝ�I��>����ڸ��)����<X��s�Y�(X����D��5�'Q�fq@q��,��o[f�[�<'�� Fҗ��=x��Yi�qƒ7޹v�� M����l��W�ك^�AYҏ�|z��m��z��#�<�k��F`4�C�:=ԡ�>#�?��5�q�/��y&ϭ��n���/��-]�p3���x��{#�旽��+�X\���a��$
2N?y`�\�>�d9���[�i7I����Y>�W����Y���C�5���/I*�.�F,o��,4��S��$��V������
`�[{[�}A9���G�hX�O�zl٫=���a.�,�#�39�Ta膭(�z%��T��8g�S/�א���|��R�p^�c1�C����X��j���i�J4��b�j�zx���e�{���ft�e��9j��|ѕ����ʹ�0��ʫ�@s����S#��ǁ�+-�~[Ԏ3;��3�|��N�$�.D�֢x����J��ӌOl�2��Cu�yE�Ɗ�4�с�}��ݨјb�̯�y�3��T�䐆&�|���#N�@����y�7�i&
"���W�j� D�E��
�ے��F"^�a2��$JS���A���Z/X�oo[����H3"�K`k�U��2�aB�n"��3m�}��gH��Z+s�׀��$�:i��*|-a#��Dyׁbт��ާ�h���-Y"'7�!� ������X��ջm���C$D�Dn3ņg��|�4�}���`[n�e k%�m���iY~+f�9ƅf!��שIB�z�[�)e��qG��2c�96���C���xn���ڄ��=�P��ΫH,V';��pwі�r�A���i����R3t`B��!���{ΩXn�V)mo��cn�:k�+\˲����w,YG��U�O�ꭘ��6�*��I@��5��W^ӝ��x�9
��a~���/�b�Gu��;��|���w"���"7�u�A}��̛���$r��׀"fqej�.�vq~��u���\_-"��x��y���Sg�,��O�oR8"Ҟ'���y�S�0(�wf�b�ZH�ޟ�گE�e�O�Ax=�"ȇ�6Z5<�֍�l}���C�\��B�ѝ�4�(S&ˢ�q(��.�~]��6̢k�>>��GA��
���/D��V ��l���@h�MH����n��\R�P����u�w��i�iT�\dn����SF]�YC��15�<��^��4=7��U�+*Bޜ�ȼn:}�3�E'� :v��
S�|�\8��,�e�y���.AG��S*�v亱�7�R����.�A�Ƥs�7�ƱR�n�?IP �
��c;�;��z���hn��1�be:��>R�Z��C�NZY}�fr������̴)�����,E�ݣ�\P2@ha�}c��^��ykp��Igh�N��G
�����S	/G��?�)-��tO�b�_����m,7ܖ��43*Rr�ox)ׅ���&L6�&�zqhyc�dvj�RtF�	BܺT��d�>����R��߯\uz�����$Ī#@iÌL����XE����p�M���~j��a���`��Ֆ�m�-s�v��lg��/�=���sR,x�<�j����Y5��)(�)B�ͅ.F�=Z��2<��b`����,�Z�x����1X��w�E�]��j�Q��h.�#U�X��*�ͩ+�������g5��r�ǫ?2���b)uah�U��E�\��]�Rۀ,��+<��a� 8$S��yq������DR�Fw�5i��-���RS �ޚ�V�tl����c�ҟ$�^F��N	�iUx#�(l ]u���eZע��M?������:�rQ�9�>�.�i��?��q���*G��s�P���K���������ض�7+R[�ᘾ�����a�,�l�6��-:����/-PH �ƭ���&�$%��!�\��E�\x�S����Ĥ����!���o8��Am�Zm�H���GG���9� `N?�,�b;�<|O�v��	M��P>RZ{@��9�~⨶f�� ��3�̷���k�$ f����]sr�����X�~-�ÿBah5�d��A>+v����b�,����h���dL�O�t{�T�.�`���$Jo*�u�7���>j���5Q1}*͚���(|�I+c��l"a��fϸ-�<�̲YٛI���S��d&"Ә� цZ۶NĞ5&+���K�:����n~��J�_p��=�T�?8�ؒ�^켧�|�l��UT��s�W�q.ӷ�<�vi:�����:#�{z��u8:�ڱ"�o��3C����U�&@��p�Q�x���Reml?�`cj�_ �T�dQ��!�'��%$��		!�d��<��x:Ek�D1�t�x�]r3��h�ّ$��䃢�ha�8n��Dվd�~j�[�Wl,�\�*�`���5�Ƒ��6�ˀ2z�c�(u�և���+�h���{GV/s�~OL�D��~�����E�������F���:׭
��lip(0H���r̘��u B��A�x`9ɱ���
A�KM������*?��t3Nm�=&�=��w��Pr�l�2�F���!6�f�/WH۹�Z�T��#�=Z��;����5j@�U�,l-��2��B&(l�������s8�5��p�|��x���f�NL��F�->�N��?.`I�,Ys�O�g}�k�m�q�����H2��%����������Z	e�5�mU���	�an��n��Nٲ�7�%DϚetl���n2hL
H�����i�S6��Tg��\X;��ͺF�,g���ㅮ#E�B:gR"�n�S�ttr��q��?i4�}��k)�l^ZO��5����ՌMB�ǝV)`:�F�N�_Q=�pb5�V;���G�ArseZJ�-��)��E�^d;�CO �H����0]��r���ՖW �O?�o�*'�	�\�Q�wOP���Ɣ>5���i`��6�DGd�g_i���!$j�ۊ1yQ��򐫊q�u�R���%�����ddr6u:�W���QN�WG��;����Y-��l�@1��nӿ�j��}�'�\����0�Q�kTΚ�l��8�V�S���QT06�0Z&�T�Cx���V,�ؒƹ��r���y�t����E��7Mhb��9���P�v��FWm�<L�����b��t���k���z!7��e�3WP��bp���8���fEE��>�VӇ;�EK�:O��؏Vv%M��x`�z�9��1/�����Æd�!��d74zra^�x��oBo	&��o#�@��� �We��?Q��Ѷ�I��7^H�Hk<4t�7�손�xE0��ŏ*4�,um����Z����+SJ�ـz�����僗������;6F�r5�	�Ν���V'w�I���!^n[�Z79���b�<���u�2Џ��}2C'���|/�������⩴=����?�w�n�@M	��"��7M��z:���P��'a(�a��W.|����S'�g�7k�M���I��橆�����^�M��f�q��-�s�J*Q'�f:Cw2�r�/<*��LCEM�����iާ�C����P��	����p��3I��\t.�j��j��Ę}�c�&k��,4v�/�)�?��4V���#T���L��D�*�R\�X�ރ3䙦eߏ������۪�����,<r��o��B�%碢S�,:�����4vtS�^ޡd�UP��jl���(WK��H������"�ڒWO���X�ۛ���#9�A/��[x�1S߂�'�z���R%�+.�C��K�,�o�i��<�;Ƴ���>T���z����Q���X!�Z���t���`�&<x�N������P���$G��g����^��l���h��+"���߇�jǍ~�xҀ�%ʴQ �N����8�@R������[�*��0��kE�D�?a�������W�1�(��Gڤ'�~�E�i��"���O}�O���k�x�nD,${!vdK��f�� MK��3UU���J�kb�97���s�0��R��.�	��%��	���k�c�{|B�r�.=.RO|u�v��]9So��=~���e���&}�`�b�-���-�3}V5����\'4��~�0�8{2l�I�3!�X�޺�	�k�o���k�G���'��]�l/}��D��eOݗL�{���h��	o%"�ߍ��Y���A���xs�������b����2�����.��K����@�C(�Ē|� }�pK��͹vb�ؾg�5o��@�A���?�`�:�݄8.��
��33���h��K)!�%�3%Q�WNZ��{�5z�Dl ~���9u�2���qO�-yk0�/�ԏ�\������K�˗���k4\�8G�g�P����|�
��"�C2�ep�v�^Y��>5C����
x�r���,�+��=&E��d�x���;@x�2C���F��d@F��Y�~���Y@s6��&z�eB��2C	S�c8�����*S��H�lIފ���'=m��4�|���<^�����Q�"D'�I��ZN����_����@������!�p�YS�
J������$�4���q� �)>7|#�"bF@�����ɺ��8�s��	V�qU�c�U��Z�O�׏���0_L�*�����^���b�
�q+'l�t��/�׏���I3��_�;�M����*��'(��������������5�&Ԣ�(�1��OT�<G���b��@����ֺN�oчOG��_?�^��u�r����R�Ћ��=i���&�c�zd��V�����z�a��p���lr���ua�f��H>i���Y�����u4��S4�ωB�%[����������q�j���X����?�'��D�&�Q<��V7��!U&9�'N櫫v�c�09���ܬ����w�*�̓[�7�jgI�Ó8��0���d��32=/\d����[�@4|~k�k�*���� t��pS[p�  S��z���u�Zh���ؓ�V���f��'E͔Q�v�\���(�QdY\>'�*�"$�1��_Q�∥(�>��]���7�k(C�+L�\�#��פ��L)7N�yg)��>�q@�x���4� �I�N��a��^e���s���2:��[���N�O&q�D�+�u�^z�I��l��\�LoMf���9�>=��od���eI�VGq���r	�����T_zB\sS���L�S�-�Jԫ���w�9���.+��M�5�ߧ|�	m@]�*ð��(�u�꟭�W���6 �-�/ÈZ��Dp(}����*�d���dl�H$��4ͼ0[;�ˎ�%3Zkz�v;���ĺ����p6�R��Q�J0V�S�\���G5g�ѡ���`j�������'����p��V���@#r�1=�8�q40r�#������
j+��c/
a�TT_Ј�ۇ�9t��g��
Ĳ�����������f��]/C�*�~!A�C}m-͖U5O@!zJ?��E���^ʱ�Y����΁�y������l��E���kuȔ���,��`�q��h��8:�:W��7q��Ҥ�+�3!z�����Bj�d:	cB-�=��0��pk��I�9�Ң�0�{�0���Po���V�b�B�".�C7D �1?��LIтXZ,.�?L��z���tD�����.�>9��4^4\�:��
��Z�S�ǋ��#�(����Ҷ[��ȮF�kp�s�Q/-S�:nuȈW��>�ĝ�;~%�%v���憁�X�}f[�s�'T�K����',����]��+H������~A�_:�����?��?����9�զO��9�/��Cu�"X�?����4���9�B���	�h~�t�O9� ��#f�ŤK0K��yO���m�u^`����s[T7F9c�eX!r0F%%�Cuq{���ׇ�ǯʐ� bI�n�O��Ʈk�=n�P�?�+�,�I^V���� * �ejϚ���29��_�͒���T���x,p�Op���מ
z�����_X��ܼIB�a��_~�=����C� S��/�mY�{-�)�"W�"�\辅�;�o ��K�}�*��/)sG�	��3�5!�5���8�G��&�,�il� p��ʑ|�x}r4뱥�ηVJ�8	����I_I�tNb��s\�^*�}C�����(6;xr�������J���Kq4���J�ym9-(���Z�Q�_���a�tѤH/~֝��Kx�F(@���i��J��S�+Ϙ}�)�W~ 4�V�&�]4���QH���p��<�d�Duś&/+�>��<}ˀ��1aݓ����碨{�UtʕM�`��Tfsȅ�W-�-����d�
��8��m���>ڟޓ�?9~Հ��^��nx:�C�?�y�p���U1}��H�B/�&�,g�_�2J�!�ΛF�����E��4�JM��{�&ڇK�h�4��qm
����Ln���[�`#��ڑD��:-G �!�7���I,f{����~�n������ ��i�j)��k�?�����2O`a�	or'Y7��['&[7�-��Wd2eX�~��;n0�k�mt�`�N�����䉦�h����҈d��CA��X�_�ϛ;��b�
�"���}�tH%1:5ܺߩ#�}_��%�,s��X���A�$�E�F�LU�/��H���5��/�l��.��a��c��F�-L,���JD�.�����(vPN�v��SXQ26h�5��	n&Z4M �g�j����i٢�m��qVU�UU�Օو��c��L#��W}�)a�����!>�z�t@��[��/�ڦX��q�uR�b����#��9���2��H�9f�Dgs���Z�yJ��n'a,�A�)ՙ�sӳ�Á�7��n��u��A�/��f=�n��d��\��n��uU�V]E��F|���]2�f�f��M������p)�ókM��������4��h�A	��	Jd�r�z�h9Uh�6�P�"�Ci�4�mi���"�u�C�'q�5.�Ι��9��WI�i;���#�,�N-�G�X`���j�qj&D�o��	�?���A���;�u�A��G�� vFn����zH��k\��� 4�?�-��R~���޾�n-MKʃ8<_�
�Yע���9�mԉ��2D��1[=5�oq?���u���
ғ?C�<��Kw�u�!� ѭ���9h��.���g���w��[d���=B�Bo��P��T)A8��ЯFՌ��P	F���5�uّ`*z£*�n���*L�u%�K�*����L��D%l@��ݗ��J��N2���+���ӛJW�?�Xej��>.1O����O�-˞$�b_�$ٿl�J��|��R?[!H%4Гe�l�� �Ua�P��D��P���/�X'qK	���k��*��� �j�q�Co:����W��Y���k���\)��)��K��i���*�C���;�Ŕ'a���ˮ0��P���2u\ -%� �0���-�.zƠ��6�sO~��F��ܷG��垱$�".BJ�E�ͤa�X�:�����9щ���F�O��_B=�Ld�� p�w5+i�!̅s�Rn��x��T�n�̻�q�Eg!|�aD�U���2[H��J�(��AG�3�nji��9z�*|jBi��w�i��7�Y8�6_S��ޠ�X�b��˞C�ÁZ&%a�F�;m�<͝qT�O�F&�A���ׅ��-�N�^�1+U���@��;Wg�3���4�n��9�����N�gA�S>��q���jϖu�{��/o��S�3��̃B���̍V�a���(����%T��;�|1����4��f�&�+O��U�m�>�Fv�Xӿ�R=h#����s�ᱴ!��������wu?�!ǆ����!K�֕���TX��j��G�W���ph,U�u1[yv��0{�H�C[9UŰ	"�F��cB��X;'/fIl��w.N�!ޢwH���Ϫs��_�T@uQ�0��G��rH��m��իa֮�g�9�|^���:��g�+Ն*������M�J�LQ��a+ʟ9W=hw���πEvb����^�)( �U���nV˹k��4�E@���-�u%S���ex�g�kC!�ڔ�RL��u����'�k]����=��A÷pT���ji��G2�qB]�9)4�7	�>L�>���̔nKP�Lh�
9�^�puP>�%`���4N{�$�*	�����\�d��0����Ű�ذɓ"14$VP�p�>��-�P�7�����bW;�8J��iǌc���|�{C���d[=o������t�}�]ퟵ~x��&�:��V�U�x�Fd��Rk��s�'%����L2'*��/kJ`Gػ���@�\MUb�4� ��Е�5�s��w�;�K�D�37�Ib��r.�~u���^%��6��������x��\d���B��aN�l�vӼ��^A��<��oU�B�Eb,���6�@�Xm��QP�zk�x�x��yv����?I�%�y գ�}j�_v��c��7*�'��]"�u8*�O�+*C߶S���jC�9�]H,(��([F=� ���Ωd.���S�~�ym��U/8�+eb�ֿ:	���-&C�ة�*8�iV��B����h�x�~*j�1d����?� �|
y�VȖ��nQ��{5k�*�7���_�.8Ü�|��B}�F�d���O�&����=yf������j��[�䰋������������q�F[���m�I`Ds��3��n�G�#p���c�؝�O��C8��[���74B!n+u:�]o���,�Fc�#帆:CC+�����=+1��:������նˁ�M�REZU|�����	�F7����(I	1ӭ+~�ybz�W�(�e�0[񜡍g��mWd���F�\"����C��{(�=�A(A_�i���J]�.����G��OhIM�0�� I7n)�0�N���R%M\��[y m�M�e�7�r��I�=z��4��a�o$��͌���`ϕ=6tN����dI0�������n�1B.��X�46��a�a��'��{���MI���i�w�Cٕ+(jC�y�x������`:��^�U�ג��pY�jˣ��sT�}���t����r+�O��b��j#2"���G�%�uxdo�pd��kޫ43d01����?�ٛ�6�U&j��X�ѣϦ&�L�0�8��z2���n.��#�Py����^qߨ����#�D���C������2ݰb���U�^������sp�EOR��ce;�	��u�\׳<0詵�7�H0��:�*���Rt�U
4��Kㆹ�@˃�[�X�z�R,VD��TF�@��؈ ���U�	р=�<��#]��={���ҟz~��/m�O��ùi�fį���P/#�:J�/kȊ�����QV�d���ؠX��TZ��|��&uO���*��=�9h���H"��sTe���MR�[P���N��l�H���mDB�<��z9�A����̊���U��Rw.����!�����0�.��΀e��wiנ��L|R�P!h�̨���w�ѓ�x���+��A��z�D����?k��џ/K� ӄ���b]v@��(����<�
Ҝ����O����<vkS�F�z{]Q|��yC�M����Kɘ��+(
���ϳ��P_�(�����e��P�O�k��^⎜��\�Judl��.[n����z����W>��K["��=濬#��$j �6��Ĉ�?!�6&�}��'>���
`�%)a��|�6;IG��z�Ğsn�������K}9�MO�+�:*Bsp�Ь�#O��I�nc9:Z����L6�h���� �Os1�M��&P;�@�L�!���g��L}O{���R3��k�0(�� ;�Մ=q|4t0��2*��\##8s�=��\Ļ3��H����n>�S�u��)���j��iUQB�H֢�r���p�~���%+w���q�Zu�*�]�d�7��܊� [bIA���lHwfYO��3"��4.����0������O���N"���q�H#ޒ��{-����^Rɋ�m�dB�j� 6�Ɛ���딌D:��ׯ�u1�؅���r����$��6�Q�9&\pf��C�"�V�l�ssl����R��	�"] x"���p�b#�_�]��rTg����_�o��	�5�;Y��ϵ/��P*{���#pw�C���nӉ�� ��V�3A��Ck�<�d
P-�w���֧����<Vjz��2�6ExCf]iz�<L�e���_�ӄgO����|������PP�$�.w���n�@U0D�[XS{ͯ�P��D�6{~D8���2t3Ҫ��Q��G��U�+�{�
U������o���)Dm�������� ؝ ���k
%�J�4R˂����m���}8�v�A�/����g[��ߺ��գ�I�ʾ4,n�L(��G������8���Q��� R�1�
������A�
��0|��1A���xeU�^v	��a�i����/麔O�k��:�u؊�~�Đ[:ñ�%Q��Q�*��Dyv"@vGn��uA��"b���}!�l��;���C�خ�[K]�D-&�"�Z ��87c����ֹ�
�H�v�u�Y�5	��V�%���0m
KyR�	Fm���#�fc]C�>�u��K����aqˮ,�1CTo���ݖ��&]gP���r�����=����+�l ���=9��aMT�J"�I���O���U�{�����0���![[��z�CCъ	�$2* �⢩60�$Cҧ��7J���X7��e���9\"I	yY�Ro'b�!�:��"�̀������j�t��Gʕ�ݤ˳�1+��ƍ�>���Z���nj��m��#������
����OG��..�bg�,O����w�1ǎ��U����#K=;���FA�ć�A����9�i/�K���s� X��u�J3�u|<��a�
[��Q�����a%�Y
���}?� o{�l61���G��R!u5�ep(?F�~��J��vp0g`��II���ym��$��V��?-ԆC��S%4�ÈO8b*�d��BB��g�������y��(:�N7'��]\��歫��M�Ǻp�ߝ�mGN���t����ѥ={4��<7���(|\]d���B��`R��x��vw�F��\���O(*0�-L����C��¹�tL0=�������7U�v�j!4�ǫ-��������A�N7���ٶCˬd��.ҁ���&��ɫ+�S���Q�p��_����"ّ�m�ȾRzeI��J
��y�A�zz�,I<�{c���s<��FZw_��&>U8$��ǋE�����$�Ph�lPff��鹘�G"4��B�d�_]�W�����ՠ�����b��Y�����%R���P�����>7Z��'V<و�N��F�I|80���SN���2��f!?xp�MV˘�k�c�_ހ�]Xt�k_��Rf�K��b�:Z��'K0����ʀ�3�bn�z��=�����C�3����`�Sm��f���f��ea1<�s���9��Ż��O���^��T��8�@����v�����h4�g
$�b��]-Ʈ��4���C�<��������� Z��Dut
,	���TA[c�p=�K|�L��-+����m��+b.}D�G{c�R����^�-�[Xs@^���dI��'�_���[s�'�0ԟ��Ԍ �ƍc���q��U�(�]sf�n����5%�e�*�,`>��cOK��q�	=��o�W9���������5"�KY��

 ��0�s��b��5�y�%�zRZ4-?	�|/�������0 �Nބ�Tl�߹�s��n�� ���k4&�~�r0v�![�̏3��w7(M�)ʐ���-N4F�����A?h�9$$r�aw<V�T���$;���?��@p2RF�5�FbN�m��l�\l��������k(�v��h,��;�Î)����M���X>6 ��/��7�hv}Q�����O�0$R|j�U��f�Wa��^�-��a)�>6Z*�c�f��T�|݂!�5�˫u^e��b�2gH2<
�l�,�/d'��rm�(�����^	k P�	��Cu�ik'��=9R��Q�����ڈ��5��=��U`�m=]�IE��IB��R�6���-c�[`bB X�N�<m>�}oldw�}R���<*���ܠM���1��+�����U>���a;��H���	�;~|gv �>U�C�g
8�0��Ձ=k���4���<S|_��Q�\�PvR��	��ր�F�k?i�eu����v����q%/��$���}�S\f����@��B���0X�L����n�f�Q�o8y�����x�1u)�z5+�,��l�\�#uJ�5 x�W�)_qԖ�DfF�LJD/�Sͨ�H�1͑8u���tcU稶	9��C�g�r�l���T��Qc,\�Է�g3�<+�,>U���,q��k��+��rC_%���"ԝ�sҁ���7�n(�z�(;n���N�RF2������v�LtP�"�T���VT����	{�k#�� ��z�3��5���Ijg$J�������0r`���)��(+�:���x�s0Z#����N_B �&�k�4V����p�@F���)3\ ����U��1ؕO� �[O��J�y�֢�ě�P����6?'�f�M���$d��e�oR�R�ە�e�j�.�q��R�q<��mj��o�qxJ�(V� ��$�8a��1�)\6�Җ���F��֠�ʘv|���Sy�'�݅�R\Y���M'��ʶ�'�y`M�Yy����j��ޡ��.�A���4� �Vj�^ǰ:{����(�MW̯;x�:`LKcx����*�m좛�二�9#���m�s�Ui]1�Fu��[m�7�>:�}Lk����%P�Cݢ=B�̊PTrZi� DY�s$�8)�p�3*N�y��h �Ab��� ?���K�O䁄����l�`���{>9�s?Ix_�Fx�l�Kg2�d�<y#���N�[��B��G��;SȀ�W���6ɬ�-P�`�0s���&@\��vU4�KfIa�e��~}B|��⹭�D>^|�K��e�R�2;X����\���vEk��*��z�2˺�^=ꈗ���!�L\l��4
xö�:n�j]�E��#�*k�Y�\qx�.�_��D�X��C���oDD�����f�b�ǕaQ�X�l\!ᖭ$tt� �;���)��Yk���h��8K�̑���e[�{�M�Շj�L�d�p}���P�4xç�L��l�p�[p��j����J�CFsB��@sҮB�^C�4��Q�q}�(��@�v<7���>4?,}�Ų�!�S�7�J�6�vm��eB�.t���S�^�Z0QmW�G����T�.A��i�4�U��b����৬W9o\��&H����۞��3dL���Ǩ�"<&m��~��T�R-D�ŇTυ������wVº̍��kZ�����*�3�G^n`�+U�ggї~��������Չ�n9G�*������$׮ߍ��r��oɶ4�~�������J��P~wpϥ��O�[�E9�����`��b