��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"�jI�gɐr	�51;.�0*����]N�.i��J�ۓ����Uld`�⼂o=��q�L���^NS���<�_GXy-c�w�j9a��r�n��[ج�ŋ��pR) �qu}�Ot��v�n��� ��Ķ��޸YB}Y�`F�r+����$��:�+ŠFA#s�S���ȱ�k�hhm�h3��Z�vJ���Đ�q�3��l ��-�E�a#0a�2�L�mJ�ý��ce#vPE�bm��q��z�����r#}q���\8/Dbu��n�*�vo��G0�W�F��� ���
���4���������NQ� �c���-V��<���3�x���`d*J��D�tQ�Ii]�#�P�C�z� Z6����AV|"9��--��	�W`����HO�W����.��z�,m����������ʕ���cG[���#�,�{�9��h��lJ��"��2?q�W�
&�e��D�_s���Yk]B�n0�8b�Ax]�����5�d���?ê��b7;�δ�>���
2������T�B�<?i<���dT�+aŞ����:�q8Rw�9jM�D��o�?�^GB�jo���b���$�t &����>rRT7$�_39��GA%\	
H�6	'̉=��7x��G�x1�wqa�^WoB�P~�I�dϫ��ji�6Y�֒�)�0��~�*��l������"��)��x%���㉎�������t$f�m(Q�l]����'�<�0W�($�3C��b,3�N�3���Gۓe�uX��呃=f����)���d�p&~�r_l7�E�X'IF��	��n�D��>��Q1�[�91L�r��}�Y��飡���T!�m���N�FI�?��+���ɁF7��,ˤ=����3q�5;]�%`�*���e��7u���bSFz��9�Hڑ�6����F�U�i�$x�˵�.`+`[����2���h��&���ҭd�X��&귫r��
�=�i���A�uAD'��93�M�g�s�z��P�/�0�Y�X��	��	��7F�==kV_VU�S�[cf�9�3�|�q�>��(���? ���-$N8qvA�۞L���Kr��z�X�cP�25���.�̓�)l�Y6��� �؅�}i+�\ǥ%93Cyʜy����<���B	I�s�Dߞ�s���
!$��(W։�����O2:�&�+��A^�/���~�$� �d�6,���d%�*�/>����̃Y7��h�;���9&%��*t��-[����l�sM���ʀ���-�w(����b�M\L���E���H-�'���~xVF�V��_�i#i���ʆ ��IFӇSX�^�=vV/��pv�w���RG�ђV��%��!=���	��� g��x��$G\xy`<�W�sȖ���U�RR�e�lls���RtU��2E*}x�r��{���F��;���H���Tq<w����������[7��P�^��ŭ�.�Z�:C��uU�o�ZܸXL�U�ڹ0�S	�#/#	��wE<l��� �*1�9���weSr�d�a)�a�,_�t��m6W���Z����	(�t�{��i8yr/p,���.|��Y.ޱ{V90k��m�����D>'N��S
>-$>c�1$���#�꿗Wq���2��� ��Lc+e�QP��-�x�����}$d?�_x�-�'sO��r:� D���819r�%��7U���I�xwc�X/�d�w���/�q5
r�G�S,Њ��I_���z��9�����DiS�:�i��#W�_��$j?�nIPŉXD.N����}����I�	b�=�������Pq���=����Í�����������z�M���\6&��:c�~���į�_8k��|@�D�ٸ@��tba�$HX�ǔ�������S�<F�N��d =��t�.�[��&F+�M!�Z��N���\��P�띐�� ����x�ι��]=nqT`⧔���kYS?�*�+�.�cJ圸B����8�GZ�mck������j�L�.�c�M�L���O�f*��pm_�b1��u�#$&`�P��C��U�I�]F����[�{���5v(U_�7,V ���_���'���!�>��F�Pv@]��K��"���q��<9H`/�ɲ�;�6`q�<NOjo�C+ۉ�лK?4)�i��)�ӥ����8<w�G��C9�@s5)�Yz�k��ܙ��kʈ1�"��N=}˨`�.u��v��vT�R�.��F��̉m_F�18��_YA|�b��&p3&�Z����c����� `�󪆠�;�������+X�bw��I�J�-=-� Era���w0��;��2E��0��@=�]N�+Ώ��Rf�	���@�]NÏ?��f� jq�_�g�|���_��_"�ɟ�X9��;�
���o�Ǥn�=��Ȝ�P°�[١_d�;�9��8��ဢ0����%`��xh'r��ށ��xI�{S��Iq���f�w<��tf-�;�RI�ck�e��t�Y��''đ5�<����Fտ%�EW�!�������/Ɋ@kK���`L�;4��r��vū��a�t_| TN�E' _�����C	:�4Z�p���ta*�=t%@8��ٍ�I��V�5A�h�m�]�i���:/��m� Z|���|�h<�2@�r�#�:~�����$��:+����T�5ۮx%������U>C���yi�@��7A���Q�HbP���h07����R���/Yh�H�li"Լ�L�Q����[�Lj�כ� �ݑHjl�&`��u�ɘ��6�-��VOA`1�������a�a1aR��{��X�h�6?���F6�zh�tTƀ(�0�ۅQ[$�Nt���b
cC��ӵW9�h�:#:���۳����ol7!�hA��|!`L�#j�M��ҌB�>;!u�.���@v����� �t���'n�0���c~͸sI�b�?�*$k$�D��]~e�����r�q<�s�2b3�lK9�P �d�NF�ݤ63�R�/w�̻w�Xɥ!)z���8#�.�cmB��x�@�3z��+L+=8e�Wոԗn+�Ƽ����.=�i���+�ɲ�o�$g��.��7-b�яπ7��
ך
�vn�\m�B��X��e�'\ηǛ�զ�	'G�VTJ�R�)���s֑�6>'-{�	$Ϲ��E�*M� ���䵳Ό_m���Vy����ڪ8*ZL����Iѫ%{ℵC�uV�2�G�e�>(�F%.��\Kx�[��1'����`2(�R�X�%�L�xx��r-G[0�����Q3O��a۞ yj���oȢV�Js�.�uh���
R.c�V���ķ�N�c���ð�N�S��'��x]Bf����[�5��#L�rl�����⑿�\q�v%u!����mU[���/S�Ӗ%M&�Q��:�8n�,�pJ� )$�0t�3GH�B	!{?m�y���2�8�M݂�:��\I�P���7|�����t��8�!�k[��[��>�S�g]�A��!��nWE��;�8�P����ՖZ���/T�Y�Y���F=����f��}��b�>�ڿ+�f�� ��G8`g��ڌ�6R{�4��F<��G��TPʕ@����G��J���/�v�[��c�%��ʆP}+�&p3�WY�|�݆D��hw$��K��p_��V���v�2~�JT��+�+H�v�%�����Y��Q�x��1�K(Cu020쮑��$1(>��N�~�t ȳ^
�!��V�Ўtt�0��swy0;G/paK&�.��R����Ͽ�ѧ�e�K�*pe�)�����׈�1��,����}�iP&1�~��۱�5%uJE�W	� ƻuLH�����&�79+ 35��P|�v�@�L�Hb�5�z��ؔ{�J�����D��3�|�M�H�lN�� �/��5K9Dՠ/��u��������(�I�a��üBB�G׫S��?���TF1_���y��,�)�B�]���7�6{��ƃ��5�lȣ3/nٍ�ǝS���O H�r��k�"�w�^ڈa�^!P��������ɧ���l5ZVTv���܏\�a�ي���2
g�_�����Љ��E�;��S\Co�=�ev�+J��H<g����]2���k���(C��4Cy�{}��!�hv��Bxօ�P��,$�<�naK��:&a���܌�mE���E��d�x��c��1�R�*�Ӌ9���J<,eZ�-���8HfRR��F����kr�&
�}���$��3?�a�T����-[���y�hd�����&l�%���	�H���[6��tt)����F�f9҉EA��dJ�����=Vf��-rso�k�4a�� [�q�閝�6�4��� �����Bk]S �u�c�����P�6a�J��I@vr�=5lʌ_�q��Е��uj{��Te�������Ȅ�A�C¼�j�j|�w�