��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9��m������G|S7���X� b�=Z�Q��6�;�L`{��JԴ��k�]lW�<ʣ�pJ.͵,���Fz�ԃ����v*H��Y�ݯT�H>RSw�I($��W��K�S�ڬ�d�H��]n^	M�[���|l�̇�GL��`-��bc�|Z�5��ЮQb��Fp؉���@gȖZ�Oa8����qy�Ut�_F��� �	�IV]EY��b$X���|l�!W��jI�IM��$qW̮"�d�L����$Nz�!{��1����?� �(�.��V��U1�m�c3.n"r8�E�7Ꮖ�-��>�\��eZ��3y�X���%=��+���F�/0ou���':�_�Gk�țÒ��CΞ���_CЧ�����;N룿^oɫB��	)`i�ǁ*T�'�����K'�9����M4��HC_}-�.;��8�71��ɭݿB�8��h��5{炼¢=K��#��� �n��^�<� y����P�W�(�g~|΂>D��Y��N~
�Վ�s }�=}?"��p�B���
��{L(�O+�
�fe��&z5kM�9��|�a24X��U�O�g�$�gM�L��
���]m&�BK��\s[ݻ�_z�4����y�I�
M-\Ɛ}��N�y�ztT�*A��n��N,L��1U0��7/r�08�Ԏ������(�$F
o �$�rbt��3/���n'�^�N�\\���A>�1�U���e���S]�w;jR/���n<S�X_�����0*��M8K7��!F4J@�]�f��
���k"^��ǐ]!uGi�V�k+	�y췃JX'1~٩��ޡ�k3a򝇫�|+E���a&D:5)E�Z#	�9>��S�����/D��Z.}I���H'Z����[jSKZ�@7�3h�v}��+�E{���礅��iB���A�4�n�p�/��m5��K�d��*w3�;͊)M���K�������<����m&��
�ʡ�}���`v��:5r���5ˮw5���_�@�2�{2_p�i�"��BB�[P�e��P���]�KxoΞ^��kKd�ԁ�{�@�M��mu	Ab;�
Ӆʄ�l����:U���OW��E*v�l��?l�h��_�>ʼ����s��R��A�����$Qf�V�%��Kyh�g?;�uA-��� �q�U�Z��#�Sv0����2�]u��-A��@�<��z��]�̂��CZ�E�����+c��9&8�RA_fz���iQS���a���˛�J�����|�)~9N�'Ć�=:��٬�\@���K�2�=�m=R��{����Y[��B�_I%|�����v�=L�j�.Cw/8�\F�U9��fQ	�аC�M�T(dl��D`E�:�d��i��4=��
K]��^�F3$�mH�aQ�|:��<UѮH���{d�u�H�9�Q���V\q��U]�A�H�Svm^H$1�a��d�ZfC=�����	��gT�D�xW�1d�K{�
g�TɜeY��/L���`O���0��&��p*�L����3�6�N`r��P���{{%a�� ���]u��ǵH3�f���l�p�;�@G��Hdͧy_�^5O}72¹h\{}w��By�4�5+y�����R:7l��>,���TDk"�ǨNs������pėNN�~6��cCy�M�8L���4Ԓ��Z���Y�	��w�dU�Q��j��\�ɫ����U7(���͸=�$aY�䓓�Nh�/�嬕|�Bs�?��ɡ��!���'�x���#��T����Դ$ؿ�N��ɮ�3y�K1͕�t3���G��O���޼B�%3�z��?}f����fP������k���)\j�KS�{���k�t�OĂ�9c� �IE����wg-q��!kJ{;D��R���R���Me����,��|dW�2�*�`��@�&]��8��� %S
f�,�(��8t��"���M����t��ZQ��l��W�u�e�::4��m��ב�l��5o쪙R�m��GԂ���� `i���tq�� �z�)M����kպ��F�}D�H�o�C�3VXe�������3oX�Nj0���)��c}eͥ�����g�%��6=v��b�]}�*��د��S���C��7���ѱ��i�7 0L�[j
��