��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<�Qҽ�������v+u��/�T����i�Y�h>d���7	&��m|�hK�#U�7QA�7�P^��N�џK7d���7sT����A�c�58�8�{r{���@&;Z��̶�HS�#4��ᐔ	���i��nm4YiE���[b�L��!��&�Ei$��ζ��y=�R�Ԅ��[����H��i\h��0�e�x�w �H��t��=�㩍���a%�����Z=��� �_��]��`�� �eA�x�I-Ki��h��~��R������D�X����;��������)*x�5I۰��k�A7�1���W�k0W��<7�C���1JQ�p��u��`���G4��^�ip�0��4%���pJU���m@3�x�^�� (.zh�� �@z����1W���:x�f�3�6_PI\��c������6G�<�@���ҕ�kc?2��
'����֟��*.�c����4 8;����%m`��%N��٦��%CL[���4�3g:Z�PP��f���]$?�5��C����n�"4&wO�j��u$� p��-���j��7�#K���o��g������� ��$q�)�����'�t6>����q~[OX�-��B�%7�*�Z�Ӧ�uƳ	�H[�K�)��`���[�Q0�����5�LzY��\
Ao�	uu�<�IC��~��sd�ԚYa`�WNJ�{ns�*lGY*��:�Y�w\7����WH���l��]�R�S��'I��zI�"f�w 6���AO	���[��%[k&;���;u�iKAuN�4qX���Y@_De"�o��m�4�r
�^B�y�Џ�M���z�P�cd�k��ce�m��Ə^�������~��a���C�Mv0d���)Ee1b5�8ܸ=�v����[�ں6㺡�َc�ʗ��ӡb�N�>��s�����|v|+��@��@��|/���HoQ�㫐���؞�����SJ�*�i���E���u+�L����@`��S4c��y�ZR�8O�E�Dn��x��AM8�v$�V���]����V�XI����e_�v����2�G@�6�`t��g�G8�@�E�?{�T�K%�-�`^qK0*r�����g��
���2]����6��S�+�)�Tp�}�2)��d�u~΀)Ɩ���$�I�?�?�[؛?iJ`C�{E�)Rnn�����8��>	��9�Q&4�Ⱦ�y�1�߽�	�s�4L[ L,엂�j?��� J�Gk$�@��Ѯ@�d�띦��&̧]M��2���T2��1*Ve��C��kx�a�
_>1}S�f�_Ih!�u.��ɴ	�uՙ���u�y�-�W�����A�_�rr��F����҅�^�D���_���/@��©X�!0�Q�2`�8�;m� s�.�g�k��U��@���v�=X_�	&12J-9�E�aFQ��	ٻ?*��2��ʙ�p38������?�����#�d�9�>�@:�Of`��ۉ�A�P�5��Y�0�9&��}S\���1i����n�V��s*��@��蟲L�� ��d.>=H����o�}T��./�2N�6��>9F�@��V���9�d1D=�Os����˩Rp�'��G�Eت}�E���������A�(�0)װ������#��M�]�qW�g�7ǋ���s�z�T����Z1�9�r��:b1��׹ k�����ď�Ұ�#{qB�Uf���tφ �VU𣽂��0d<����בϵ>Y{��O:15x���h����2�a�D��F�"��cu3&�$V�S�Y��s?eN�*ھ���k�ۄ��?a@O������xCm��/V���f����(������E	p�Ək�L�_�I+u�lT��L/���
gH����$[�>��U�|��q��r�{��̢U�����l��Xv)������S{��M9�j߀b��2�����3	Nl�Q�b�H������pmZc�[L!���'����S휭�O� {W�g�̃+#�Ft�ufr��ĕpC�_���t��uSL��o�Ng��6���񄝱�����ݟ���W
����sM<���������juV�R�ZW��	��I˙��L�_k����ų��q�WO|�I�(/jB�K�NX���hjb�l�cku�K�84��Ry�xY���hq�$�:����tX����=#kf�إ�S�8O9vp;s��˴#�����=&���\M�. ���E�3�P��?� $��]����Cϊ���Ē��A�<.򫅫+~%t��V���Q�k�>���"��(�n\"�ܬ��i���Th���U��&}}�E�K�k��s�ٲs��$��N@(�8�u��4l [�F��"��=pjEV)F�s�ߙ	0�&�./k���� �Y�nw��q<^Cf�/��>�)R3�H�Yv��ή�AT�����? ���Q��r���(ܣ�7է�d��%c&R�p{zzbae�m��ҢHP�*\�&MyY]���v�ۃ3���2)�N^cH��KQ�jtbJ �\�H�� =��&�t�3Py�r�� �a��"�X������ɑ����j��INb��(ɖoJ�	:e0����*�<�Z��Ƕˣ$m��0��D��M3v�k�k�r�Ckߤ��߁ǫ��#z�R�%#r�
�w]@�p(n�ϣw��԰Z��|���S4�ҤW�h��MJ-��lѷ��O V�d�-�݃$R(�؈Vq[`N�2��;�r�H�"CU70t�`����N^c"� E�_�5p�y�u�SQ�_t���4Ԧ�^��N�"=2sM�A�N@���K#T����o ۧ�Q
u����}�����\�Os��EX p���;������J��2��*v��&�F�����_\)����v)F�J�|z��8���^�'H"z~����8Zm%?0)�����G�(�"6C �}ۤ�'�
�wz�e����XCHd8=��`�.�w���4�W�Ԥ�?��8N�m<��4^\WMbJ1��$} X���fy`�}p��`B+����:�Vn���>ײ�*P�?V��ӷ�#�3�܇���3L/�w�����-��"�,ҫ���N6ʵ��!���u�EǊ@�U2M�j[2���f����"��@��o,����a=�Z0�T��F�0 �3������	��Oa @�f�=�*ܠ�vaw���_%��?2�+&�wJB:�?�ʹB�WĿ�)�S n����[�@��V�^��ʕ�J~��؛�*lZ�oByK*����97xܣ�j�FATvu��R�3ӑ�>@{@P��h�&Ȋ(�g��EW22ɝ�RCR.��]�Ɗ�h'p���'n�K
�3ß��pB��@�w%2Ʌ��}Ä���f3,� �y�$�ҨZI��kO�|���tB⸳|����`(�iuiT�qO"����C/E������a�3b�E�X���J����!ا%x:��F�*��.a$���=���xe�?�������ֺ��>B	�hg3 �l�,%G��P8�Ӟ�0Yio��`�$��M�������k� qw���ϑ������]@V+"�ԇqkT�����'���������߳<j]�J�8ú�51��D������=D�)�f˄����*��ЊnfLN���E�CD�ƨ�*�\���S��;�ݮ�Ha����c5�?(��W ��{�u���c�`��	Qi��z(�U
���N�5��Y��c��ֹ�M��"y(|9��L�Q 8��K��q��,�^8��(�#o�ܜ�"'΋����ku�Z4-""�f`2�TA��S�_�Kq�mz][rn�w^�V��QD�O���tn��?ԕ�z	Y�g�T��_�!�/�߻
��FL��N�����Fc�'S�B4<�P	y��G�\����	:Yjp���#=� ӻ����u9����$C�����ކr� {������/��x�/���r�9M�B�W���QQE2H�X���x��XÐ��](�"e;�c��	�$u�>}�	�E���k�Q��n�+(jA���#޼�?��|�.�fT��,}#�1��M���?�]3sި��劃����IcA�_��8=Y`iH�ua��P�b����Z�. G)�� �"�B�c��N2��u�J�0iY�'�cO~���sy�#����5պ����&��\Þ��0pn�Ӧ� � b��V�h��S�,]��Ļ䯟|��r� ��@a_����M��(��I��zB`�h�A� GG���i���]���J��0@{���T�{c�o�$�J���Y�t��;�a�/�hù� ���O�aظV�+F���`5l���Iz��S�/�#�fw y���(p%�?����)���s(��o�^�kK><���#�z@�!�f��Eeb<������v���p#�k��;���[�Y2��N���/Z�.߿��@\���5�E�>M)P�r�^�ar#,9t����R{}�7�1�,�I���z�2�\�-��iE�,�V=N�%�M�pؚ�P�Y{*�*0��`��ٕ�N�~Q]�1m��X�T��YCD�<K�m��R䖯�NN�泎֮N�%��@���?�c-=G��F�ݴ�<�"� �w�əsx����%�L���c�s�R iē�+#EH�����4������t�Ӧ��I�'[�8�'�نs����n�fN���)�L�����)�Z�� A��r_亦Óbˮ�:x6�@KAC�l�e�ޣ�V����w��u6M����|�&>��h��`�aE��hR�#+T�p��kI��-Y�_��]�#~V�rl�ڋ��2z������៽�v^JMo���Y슡��N��f��Q�G�P�/]3���р?O�?ժKo�׼2E��m�~�g¡���o�ΰ�7�ގ\�5߲h��N���#w��,1Xִ���|�m�V���ϒ��ɯ߬�!3����YTR_E�rQ-�/��{�=��eS���f�]�}���7;#x(q��߇JHtdT<t�~�q+�ƕ��{�^�w������icg�������Գ��b2��l���<:.O�A#dW���'�''C�O�xu�\1F0�+F+��'�Z�\ڛaFK�g.�0�l��:���	�����u��ѤPh�
�{�ؒ���OglJ�M������	���<���4��\a�!d�È�\=����J'�5:=ۉo�	l���-��Лj���<P�d@<���5�N�M�xϤH]�Ѿ�����pyEB�dc���Ay˛��2���V�Bi!s2�!�B>�Ӳ.�Lt�޶2��|h#S�]�%|��lA��۝?��G���)�~��ԓ~	�����+ƝM�}6��We�kW�R�yP���&
w�ݗC���G�)�6�ڀ+�0����a�ucpN�=�W��A�9��*!�K4��i���ؕ��#�ߗw�~'�g�+�3����Pw.;d�!� f{�i�5�=�Fl����M�=h$�2��	�,�����Jg=��Y�3��K���"�u�yv���F��97<�ԕsu�K��<"��ۙ��LN8��?T�=M���o�������l��t*�����A��N^M=��Q��ֵ(����[�3.`�`	��5$h,_����U�b��)��.`hs�`%Տxn�av <k�~��7/� �9v�F����b%�0��m�;ku�Ȼ�h�-�H�@p����pq�w����~Omq�oӈ-���b���C�xq��pɋI������O������X�4io>�vxb�{J�F"�F�:o�aع�z��L�̐����a���($Rk��o�^ ��n!��;� ɞ�
���@�������ʓ�	zZ��I�P~����V�i���Iˎ�Qc�S��I�3����R���IU���d�Kd��L�l��۲��ȋ�I����Y�.��.�o籵r�N���Va��c��߀X�G_��v&�/G'v���#�V�X���[���6�i�C�[C�b�~���EGU��"i�D�dЦ���i�4+YP�>�y�'�w�(԰�c1Tn�S]���Օ�%���֥,1qY��Vu�G��q=��%�Mj$�6�BC�uE!������&��r��I��%�����zַU����[�:�H�����8������g
F��M9���G1cCf�������.<,۵ⱍ%�N�9�6jT.�K�t�?C*�o�����J�4�n��%��3���6<����(Ǘ�'��/+�#"���7}O���L~v�t�r�8�9��)	}�������ݷG+�=s����>����SL��v{�b��o�`L��~̝.ƭ��>{�h��Z�㮷��kw^:�(;ϗ�v�]K.���)1�z1I��^[Z�w}V�w��b���qh�D[�^�E��4!�.:;$��@�r��_�%���sK<d�>�m� ����0d�	A38[�f�Ո�GJ��'~��-RH�S�z�Z6.u��������~�jƢ	���#���P�Є8�-�;�o}���`���!�#����j,�O5EΘ�*;7yl���`0r��#ۘ��D�z���񁯮M�]�Ur'���V�lq��W��j��D4DX��m]�}dz+G�N��Gg�!܍'�Iy`D���Ÿ��������97{�FM��R���\�^_,��k��C���J�0�(�L���X�?���~i�>Nަ��V����[G�~V~-��8�[���"'���B��u��E�apP������3T�����:���k���>�J�]�S��M`3�.Me�G�"�	�G��fp�U}�D�����Ӎ����@��+������݀�fWL�H�7�a|G�����]SZM$�q5\�)!�b��!��}�q��r!�H�S׆
��_�	*��\�:���$�P�O6U�E�uu��Ռ"�+�6`B�x�֡�8�i!b������-Y �/i0W����g�i�g��υ)�nK%�:V|1��jak��!��,QL;ƞQ)�C��?�o�n%^�_�u>���1ɩ�o+��I(#�t��5��P"��5&�ho��� �d@��ٖ�I-|�0�Bd�aV��PFGX9K ]�r䢱}�oFZ;H��jc��1M��VYb2 	�D�F�bU1i�ԥ/�=1�h1�>-T%����9.�E�'��E�|7f"z�BB��cQ����kn�_'ݾ�T�";�.~z������J!_���d�%$S)7*2V������0��洛b W��ۼ	��T��l��������5s��5��oJU�|�^��X��
�gs��� a��x�x�r��2Y���t��sP|U�7�����'4��M4�xhԑ3c�U�qc�$^a��x���.��	I%�ix̱��� P��|�1�#������5%��`<�q
߸E���v�mUQ5�e�<t���㫿Ô�3�s-��¨�����)���T������:�8�QCd�k�U #}_�yL�'���{A�%??9��뒲*�2�o�yL6XU"�B�K][9���J�X�}`�ɯ�oG�e&ט���F���`|l3Vck�e��ϖ/�뫩��D��6�oCH�X:�jw��@ݘP��j�����R�����cXn�I�ԡ-��p�#+���W�E�a}���C�\��t6{ۖ�l�q��U� �Uu/XoӺ_��q�)����`�FH��!�H��h�I����:��mƷ�pƕi�f'ڎ@�zp����d��C��r(����hQ�`���*M��ö=�:�N2ҋ�Mf�D���
t1s��ڗ"6�}ˠuM���4�:$w�N��+C�s*��Г]F1d��H����p�
S��r�!�!�V��h�|ʍ3�й���uh�$��z7D#%�6�FE6BA���@�h�-��3��ۗ_��<��ٟ���A�?&B����C�>~U�%"ѯ-��"�S0�He�+��D7JH��`���]i���	�eQ�"��X�`����݊�����/e"�w4��F
����_.�]/��L� �^�a4 �����7��	�:D�u��͸8Xg��D��߈_|�׊�c�L��n4)39R��B��)K}C�@o���ƽX[˒T�v�&��O�JHz,�!�ڮ$���
�G����.��X� B�4��n�:�{���Fe/����d�P9c�HH�.<��1�AM�\��^�����&}��kT��«���)L;V�*�5-P0sI������z*�٢�� �a���v0����KQ�!W�AP]}��Uj5���x����^��@�E��C)�`:vLG�8�4�,A��-����Z�"�a�6;�(p�8)��5$�%����9}gQ{s,?�E$L|>B'S�K3�fx~�K��m�[88���UhH�c���D|̌�f�P��>h������`5�؆��0
I�`y1d������ӣ�7|=�ǭ�W��Q.�+\��RGgUPN%�zQ�{�~U��
�����,ߛ��]>�7P�����w�}S.��R.���(���61{�O����
�*[ok��+�Y}<�g۳�;�Y�3�)WLmچ�@L����
i<�ȬȤPZ�kE�Q�B}0��bYmv/��%��>��-�B ����FY���/�.��ٮgf%Lxw���E��ۤY0&��[����uk-�vQ�����H����u�i����u�tu~.�b�}3��w���ܺ�Y�����J�ʅ�F���Nm]h�}�z�� u@��Zd�.��O��Ȍ�bD�X����p��U?�<� �.��2�:4S[n
�l�T��s`���e�\Y@;T�x5��.#Ih�K
M�)�	����G�N¦�l�Dv�Q@��ߦ�U�.[����	��*���H���5"3/#/�aAU�h���x4>;6%�h��R�h],�a>����N��Π����&x�#�����I&���̪y,�'_�ADh5C��61�B;�cQGdfT �c>��nBJ��]�*����g�O��;�e�g@��֕����h�̺LX�wY�5��

ȁ$�W*�Ks	Ѥ��~nFn�QV��g�Ǆ�5��̵p2��{S�#��8�"!��<� '��������	xz�"=~D���͎�n����g�82e�'w�O��e�J~�d��Wsj�z�:Kel�,*SܓA�Y�]t@�3���)0�Uy �fVj�O��6�����O�Fs��(_��\7��u��퇯/�>6es!Y%�0q��}����bp��W ΁��~��� g�d���?tb.�%XA$d�ӊ]��@�fVDvkcb)��'�wI����o:f���7j���^J���#�������3���@f��k��E��j�;���qH?vE��;��(�����1�%0��������{��K�厲�Gi&\l]�m�Y?'}�u�S��=5�kS�/���%���q@u!N�8�1'h�"C�ï�P�-Fn��ҌZI��{��rÁ�7E��;�����fE�=�
Њ�z
q����+0V<h�Hjy�����2ŚhJ�k�<�a�f(�Z�x�a�K��͢QnV��亁tv�C捹�����2q�:�pզ����ݷO5=�,�V�TjbL��/��h+��5�3��ED虺⡨��Z��w��3N��Y�6�ߛ�$l0���l�X��FzA��I���7~D���:d*NH�!�[�DD����y(�]�FS��q�<��mci��=&�ځ�wf]�V��;�qV�bF�4(�Y+,�A:˗@\)ɞ��n�Ӡ��A6�gD^��C<"4���6�l d�y护�dJ���ZV�lM{#�e��@�%�m���s�@-�/�c��u���z	V�K�Uܛ�Nƴ�$���4߄38�F��zٔ��a�-�ު1_��տn�ȹ`�L-%���#��5�������W]/J�g�*�5�W���])7�����\q@�� ��}f��`�w�n���</��ԜU�N��tW��;q;$^�.|���9�e�f���
�/q��o�7}��ہ�x߻a��ٽ
�ۜ���
}��Lڧ���{P��ca�z�O�g<ƌ~�O��6̏��y�Q��{p2~�ha?b��\z[�C����-��(�����9R��ś)l�)p9�(�=��&�z&.1
P= [W���N�-��_u��^�+1�?l���W�:¢z�(-�"G�ߦ#ڄ���A���?�g�#�D)Upn\1}幖��[-�ͮ�]dB���+��D2��A2�u����}��ia��|���Z�0��QftUN["[:n�����y�, }HҶ9O���0��ڀ��~�qv��r���Z�o��J���_���'�q�}D� � /�n	�u���9���zs��ژo��5y���U�
���ʨgK������!
�E��щ��&<ѩP&}nY���Y��T�o�G�P��,<���2M;'�Je���,�ώ�j�N=>�Iq��!�>y�ڇ�-\Č�65�<�c��zjIy�$�Oc[B��X���r�@P�B�pJ�Z,���AeU['�.����o,i]]^�Ѕ�(ɰ�5u2���?��u��W�*���.�q�� ]�ۦ��z~TC@�m�@�*�w`�SgQcwK ��`���]r����FZ��J���<�I~�]�:F�2���]���tl���6%��Q�F���_>ݣ�H�Bh��1NC�K\1k��@��T��-�U3i�e��y$�[��٩޵E�l�f\�zK#��f{]6n64���V�7�ˌ�I�x�2�ML��IA�Q��/.K߅��!⽂��?���(�A��OT)S��}�����9��f`�T<���`$ӱ��q��ٰ%�}�͍�(Ĩ͢#&aN��<e ����L��_X��mY y��Y;��u%�R���▗x�J��r�H1ƹ.[��Z�2��o�ko����_m(PXMPXW!�W��]Ms9���m<��-�s����. �o���=��������ou�o�������n��V�bp�Kg�n�B��,��RݰvI���O)��PKl��MJGn
��6��[�օ�����'o3����i�"ۭ<�Hfh(ba��%E$鹄~�9c�0��#�U#2߹_�/ G/(Tח��!ڦ��u��V�K���$zmδ_���l8E��-��52�
���v����K]` @)�&W �j�^�xP��p�ύ�L|�دڢ��'���+~�A��)$`&����W��f����g���~0��A���5k�5E�<s.v~�E%�p�)����p_�>2�h�2�k����<F�)m�����kL�"�%&sG��K�b���l9���¨,
���V�x�&�|�������M�^
�k�N�6�|�E�d�Q��iQ�`�S�ց�dO�S|Y�dϛ��N�k��Y���f�����q�O�Q����І���C���7�1�_�yS�Nq�h�2J���t:��К���sq{>�*w��Ʃ(=eOCn{2���x�1s�P\��zzV+��<0�lN���Q��`�L{|�p��V������d����F��qIb�7��� &���	D2�O����F���H�!��^�ǯ��G	�{�O�����%�T�X!$dm;k��u��TE�r$�ݱ+��J	Y�])����>��L��
b�?G���8���[��Ư��^�Ռ
�XL�;)n�����S#�����z����G�.�0|E��To@QZ���}��2�PG�K2k����X�N���t��.$�o�1�mJ�N���e�+��O��C��j��7T�v�6�"��s)�Eo��Bt׌�&����k�!E���d�K��]sk���n�U=o�/lma0Xh=6'H��5�� �tQ�� �Ʉ?�*h}6�`�v7�b�����WO�/�l��۬U6�c�V�Ӂvѩpp����f}~\T�w���u�]���	�伹��
�a�6lJL���s�'�*\�ڏ9 E����ۇ^~nng���v{{���	�:��*�GV��@�߁f�5�>�:�'U��de��#�P�v�E��v������ �c�p��b�w�rs��iÿ/��h���`��0�/F�xT�}M.4!d[��)�j�ހ-j(����)�b�}���\��c��R��؇�������<�"6�]Zʯ3!%9Ót���®�{6�-���]�#�c��
��&N�n��pCH��T \���Ȉ�g���^���ܩg��W�7?3O���52��c���t��3YѶ�d�
s�ݘ�eU��r�=YMҏV��Z�J.+��O��S�ES��`Am��=U�����b�|�8@�|mgW�:�׌ւ5�f���Y:A�!˫k�Z%�����ЦXb�Cm�=Eɻ,I ͘��I/��M^n�/*�O�V1mv�S�ς�(�O�ԬKdž���xS��)�t� �������Brxq�2���'5�*��������p�3�٣N]�J�Z�P��l<}��Ll�m}������{
���m%��t>y�/�$�F p����=MC,?��h�����Ѭ����VcZ��l.o�%E���=P���OH��/:��bu��u*�V�\��?B�˦���g���r�uݽ�:�^��;A��c�OV����#��خ�iH\���8<�DM�h�@]%��kt�����HW+����qN�\>x'���Z�_�������q>�뵀^ha��M�����k��H:�����*�}I�x�N�V�f�Tiס2b���l[��Y]�16r�O���sE���4C����iųߩ��g�J���ƣ(�/�u��P2A�S�D]PK��+s&�'�{��a6�j�V�"5U�h�j��;���6<q�)l�(rMj�ͭye���]���p�"��Eާ<Q��&t<��P���ܞ���u�7&j���클�,�Ǩ�bB?�=p�r���+@w��xk����Z������x����C��X�"h,�h��D����	mL�#"2ڵ&��ʮ�Z� �p�N5�/��c��'ISSf�+��;���~�E�OK7U�dZ}Gt<������{.h��zt�1�| �f#��I��2
 �֕A[̶?�} �z�P��N̠�_K�"�9�g��{o�3�Y�c���7e����b����G-0����8'���{�u/"6�� �v	>t����&�=`1u*<࡛��^��q�x@��'l��ib����El�x�g˄�_�� �������i#|���)>�R�D٘����������oY����]�F�^���`E,6�ȁ�ª��x\�����5�k/���
&�gE��;>r�bj�`���.*�3�~���#�w�
���PN���p�������#P�88����=��Nϲ�38��ޗ�����j-�}d/m�F��#C��QW��V,t(�Q�"�/���~����>H�rd�ڣ=��p��1ۨ���f����E��<h��y�#n��{N�1�>��xŕ���{��GN,ɀ1h�~�n'rD�����E��M;^-��}lo��yD@(� �];�&T �g1�ⴈv`��/#uC=�6�F�Y��;{9�t޻\�T�B�tJ(J 3��1��ې	��ަh����˰C�"+(�i�J0�@���,��>a�m���:쉕�v N
��-�b�w�!�Xb%�'�o7�	|\�Y;�lo?���R�$,m���'��5qM�O�e�C��x�x����B���L�R��b,�ڽ4����o��V��/��Z��U?�o8�n��Qa-�J�1�T������p���w�Mq�A<!�(�ʅ�T���?�ʩ%(7� u���+ݩ�*%h;� �F�J@-���d�c^#��BE��]��k�mx�7�<�V)A����?��i��]gN�s�r����*�( �>�l���%K�5h� �y**f�?eɸOƽ�w3~J����7�S9�M�`|���T�֝�ʵ�9;-�+p����W�'�[7	R��m�O�i���"N��Gu���H����ҨRH����|Bk�cd)��.S�8G
�(0�/&,�-2�S�t�Ȱ�8�4���ϗ��v ǐ-2@��5�7�M�{ޛ�;�.���F�<䕭���_�=na�:��x��5������r�-��E�\Ų�`�? ��Xb�aw������z�!�ܺ��Q>���m]�x�q;a�g�R�{�'�d+�j�y1��u�� ��x>��beL�z�TR~�hb���V�z��yF+�No��E�'��� ����n2�0p%O��v�[k�D].�X�M�b�k�'w�Ƿ�t�$>�X����;��n��"�.��;�Q�S�{�f�}�V'�b�j��w���/�м�M���t����e`�jd�Ҕ� �
��B��9i&?
�Z{&��!�u3��x!R�j�v"1͡����r�<�Ggivc���7յ��0��	�_mx�F�x�J�=��>�׮�D,�o &έ@��8)~��
��?1����!%#2��:��	��R[#�_;�wfA�}��{��Z(ǔݮ���p�,�q����)�fk���n_7��gR��?,6U�P;uj`�'FVػ��"*���C�O��U�-�7�7���p?l�Ƒ��t6U(Ȧ?.Z�Ge�ӧ^t� i��e���|K����)��p�i��A�k����~"�B�2��YN��=BB6�߉^@7 #OQ-Uh|�+s!ͺ}��ڍ�'.H���0�!JII�/1���jB{�n��c�߆���>ޖ�������^��z2�rNr��'����|�����靍���~g����`���?��7�=C�
��Iҿ�����!�;Ə��"�}~`�0�b��X�}-�(K���q��q!퉋C�H�Y�����ǩ��Vo|,0|(�h-L����kgَx��P-��'l���NM����)��R��1��~27v���򖼻�S��)���$���&(��� ���le��ș�ք�96 uL�A]q���_��`�z�YB��+
��q���<WB����=E�I&V�1�<j����H�1p��}z���l��N� ����i5M�������H�����$�tJ2q���+���X:����Kxl�BbF�#��;d�dq�@.a�+J��);�����P�o怜���h �D%K#�1`&m*�,��\Y�o@~,��Poa� �)R_����I��7�N�i'�yV�4�4��W��ޚ�����<�뺱�d����֫���/)�#M�^�z�ks(�z�޸4�}OD���r��;f��-�7	H	9��?��P��ԮD�y�*6"~��)"�>��Y�V�9F��r�9����w�;.�+�����Q�h;<)J��x��՞e�53@VQ5���˃��`̌o���f�=f8hm�	���,q�� ��
�5{udZjs�s�P���N@��E}���(�<Q%�d�ω�	�K�1�ZF�OˍB��=��O�Nv��&�ap+|����������x�Ӥ^�����|���v��<9:��Am<[a��e�|����M#*+�tU�A��e��Z7�q�_�s��!~�z��1��"Q��O}E��7�R�~�9�Xo�7`>l�ʸ��n�F�?5SO��%+Y���_~�V��u�w֥y�@��̾���@���h��p�Mc����Td��JP��c�8_�:Q��������: �jbOuM����+z����i� �bX�2Q���x�*�D�P���nE�w2�	j	��IHP�6FqQjg�l�X'�3�muTI���]$�Wax8�b����=AS�xr0ή��˄$^�&���-͖d�%ܹ��YM��p��������pS4��6 ������G@{xh���
�&�˹��l�b-(�4N�יn$p�MI�A�A��]O�F��w��5��|��O��;��Lw#�%BCHao�z�uk�Џ
y6�� -����r˲�J��*\�)�\L!�;�7��`�������k�G�fZ���-P�8���
�C�m��ҞF��}���YP�W���4 �-��&��^jَ�`�|b >���vtYJy���HN���)T����T����ۣд�j&4(R�VX�rcHI��9���e���]�%Hi6|-�hV�����YD�2��Y_����]Px{+p`<��F�D6����q%�;S���Ϸߠ���u�R���zS�`�5Jͷ|avg���q�V��ų��Fo�W����oTM�NL�5��2��Z��L�P�ˇ�#�+s�ࢀJ����~��|TߏzuD��ٽaҟ2E�TL]�C��fLH�K�|�8.JB����I_f��R���s.L�$^�!�G>i�V=�c��d��a�j�@�$ת?�i��Y]��VЬ���2V�)�Dj������}�K���]����S=d�?eޞz̾�쐶�L`Wүz���4Q�A��̠ �iLw4O��S�=[�C(�쮝�챊؉��\Z�>Y�	,�{��i������Q0'�M"|��q�r �⺝��xzD��*Y�%�"H��);���~ʤm��8�B���~}��C�˔�A����lЊ+o�#��8�VT�л;����bQE��x]����$��L��Ⱥӄ̐~������["����a��Ä�[�����嗕h�Rđ���&�{ʴvt��̍e<9��0��F�RJ�%,l�Ƚ��!�!�_��3}[�o�}}���wW�05� ��_�><}6.� �(��5��B�v��Q���-�=�u@���\�K4�6�v-$�@b�_/=���G��/�!�?�#���$PP�Lk'L-�JPx��7z���1be{o��<G�G��6Շ��%*7�(�`'fj�O����"zj����RU��3K�v�b���2�Z��t,�[rk�W@u��Io+�&R%m�{�@�?��#bv:��i�n6>��|O��"����rR�������OK�Ү<O��+�V�G�h�-��,���jC[,�c	"��/��1x"����E	D�jLc�:aj�W~כֿK��� iu)�3;�͂0|l*R͚'�)�eyǠ������3-"��rZw�]���èe-0���:��7�S��q��qr��~W�/�]=bLl���Ӫ���@S��țG���!�����>��9�	���ezMLCm���P�<�B��0�r�:����5b��g�37�G=��&�G� ��i��\�|���ZAg���Ge�:�)���[s��^�H�k��CL��IND�F��D}��	�8b�B����R����NӉ�ef���?T";5�3f�F�{$&���OI�R�wk���O�d��i��)�j?����
v�V��Bnp =�	��"�%�Zl�F7�ü�p�w�Wa��9�PRh��	�L᭧�����5?�&V�����	y'�FM��<$
��Z��bkE��:o��\54�ɀ��}����g��bdΓ��L7��6�`X��޻:����/ >d��B��>H��+h���c��<��<�EC���1�I�l>��M�� ��@���>�4�8��Q���Ǥ}�V���,u`�*k�h�K