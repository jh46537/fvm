��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>��������ّ$�*X`F~�������><06�L���\�D>�WҎ�����r�.~O�I�V�X;w�G��ts��K�5���t�7��R��пr�.r���x{��}sbeq�XG|7 ��$�ڳ&�e
�=r�$��!錋"���ۆ[�8����lr���8Yi��9���eIE�(Z�)��VJ�j��?~�	��c��R�6���/�WC*��B�����-~��R���$=��&����O6�F�~gh��\P:�w�o"Z��{��ܪ-|$�EA���ٔ:�_JFJJ��S�B	*.�a�ꇔ�@�/~�WC(���&q����?��V~��A������(}�b	ѝu�%k!gŝ>�I8�s)�u{��>kp�Syʰ+�� 2����=��D~0.i4��SJ~��U�h��ERc;��@�p&)Aǳ)��� hU�`��ߨ��a��A"��++<�QE�Fc��4���=���8��~A.�i6!C�������H�����!JKs# 0&[����-�w�j�4׵�SE{]�~+��%P�*��xmH�\������/��xX���'�G�����˙
�8|"�[A\�zf�1���vdQ�6rQ���l5h�7꛻��f�*e�M�i�_�E���I�.���9��R|��M�'tǼR���_sE�m�rK]�����\{�PY��{@z��FqS�xo�����kn�ef-��/�_���ͼ�������![>5�cv���P�W���6w1Y���I�ٲ�8!��WAe�x!w\�R�O��{����ʨ�0�9Bh,��ij�w���,6ee#��+��4t㊇��0�dƘ�(H>|��N����c�(��j$FN�Qֳl7S,�+�8��?ۙA�~��tL8mI�z���k=-_�t�����BJD�� ��yp8�-K8˅�ί�2�f�V�9�e�ͼ�p]F�N�/F��=K��ާ��J�G�,�| F������ ㊔,�0�Bڠ���ǋ���>�M0���[VJ��98o��x���8 *-1���oI�@,�P��a6H�)'�bԔؠO���N:,��$`�05�];W
C%njC�$��=���f�j��xu�<��+��̊�#E"U`�����u�K>e��OrZ�����!W-�9uQ���s�}�M�$x�tT k@��jx��;K�f8N<~?Y�*hֲ�����w�YBʶ>�x��v�P=�1�@S�T�w�a�Ө�g�ã����V������;h��Ji�Y`C�.%����G,�{�3�n��C<�?@�	 ��0�qCb�#y��#�_nZ�/JR�1~!���̂(J�T]�L���R�P�;$�M������_��V&`*W��P%�^��	M�rc�mS�N!�a��~SC`Zk�o:�!�V������E�_1	t��\�b.�m�+M���uNל$VN{@+̝��{����,td�0�;-8F;��H���,��eP%As��s`n&0�U:��$m�'�S�/�k"'(�w��d�t�I� (*�:d&|����[���GB[d!u���m-�F7T@��o�L�k�%X�(>Ne4Qn2;�����0s�+�O�"��SVt��u�U��(�/�^P��t���E?/b	�j-��t/WmZZ��#(���u����m�*;�H�KQ�>��N�9��Bڏ5Z_�ӊp� (�>�S�	��p�"�u?Fj�� �#[(��3�n�^�1No#�*ܔ�H��!e�4=�����T���'�̕:������Pwω�,� �<�x��v�p�T��<����D����-�~�pTK.g1Ża�/��۰��Y����1J���4�@µ�{�zOv���+�4$ ��30�GA���oS�����P��:�H��:k��RJq4�f�Q�
���M鐦���4�^�k��?=sFsNl����^bKL��3��7�3�=J�A��x}_���w���`Ҋ1��=�Q�����BK�~� j�{��Sq+�U�N��B���a��ye˒��
���e����7Kn���0�cS�-�Āl&z����J� �e+V1��k�J�a@��bG�M��RG0[_zz:)mlJ,��?��Mk	�M�}����%ʏ�p���x����W`Om�i)��-���J�?j��������N�6���(�L����x�W�����q����0��9!e�Ay�.�l������	amQQ'��+�$��g3�Zg���ݹB�9�Ɗ��ݣf;I�t�NgK(A�4���-������ϙ���yU�z��2.�����������!9Xz?���&�H�.p?�&�@���"eBn��OVqH�3@�k$��{����Y�����P+�)��m��;n	7�|=��x�}b@_�7
�[�_���fݒ��U�e�$*CV6O&�Ԁ-y2M�`�)���̌���@#�m)_�����E��=�"��޻��XoS��HTa�RN�
g#��.91����"B�at*�Ŵ l
'��-��Nc��>/_�
�,�s������9(r�}���)駪 ��r�5���:g*+�c���.����㧮�EVh�n���f	��ZZ�0��Z��/X�]8���j0r�t	�ˇ�C�JݞBn}�mغ��w���������Xa��5�GPLw<:��z��Gˁ��yH�ȷe[>[���B�>���޲2�kY��R훱�:=�(��`���f�o�S'ub�޵i�l��'=.6���ĥ�Z3LÀQ���+���ba6mÄ�cVA,����L�����~A���E�0n�]L����/)F��q	���K�J��IR����M��L���̎]���0Y�2�C�� HӘ��	{؂�Z�)�;�A�o�R����x���ZUB�iPB�g��<�Y*#���E@H'��^��q��1vJre��!�H����)������XoU�dj��,������V<X���Q��Y���R��"|�l@ׇ8'Mj7��b龴q��1B��i�%F�=��m��X�F/�jqX:����)�q�YaϠ��
3��IS�/7��io��v?9�}�m������ٌsz"Ddaqaɀj��G�DюVtSl��/�K�ر��	-Ə�t�;+J�z8B6W�7����1;LG��w�mv��D��7.�uSJ{D�(�k��,�[#����,Z�J���D��!��KgCU(��]�E+,����os�ģ��G!��Wmi.�^ZׁX���7/�s<�Y,ܘT�s�z?���NY��-���UW�>Kd~Y&t��TuЩ3����g<�B��PI#A�R�hӢ�S�%��oD��мH�|�Gs�d<�s�]M��؊Q�qڔ�Bo�vE�JMɦ��|���߫�?�f��r]�'N��M5�K�����w�������H ��|���:*������֧7�s ֏��Pzb�*Yl�#}Ρ��z`��7�{B4�Z��-��{�n�PW���8w�#�*:3����D�*_M��Mb\���y�`Z��Ԓ�p�|3��f���R_�z�6�1�#M!�c��UpH�tJ;ݻ����C�{a��=�/U�Fr�x��2h�a6|@�S������Ё�JG�;��A��]g�&w(S�Lo�<'���[�=��9�5���2�I��6�i'Po�� lw�8��9�EI�� V�ؔ&
�{}�dB�f���
Y
�ٶ��'I� �����Z��`�i�wvΏ=�����g�af�}ϟB���tcq�vm�:Y�S�N�.��(7V�ؒ��9�L�6u����J����Mŷ�����V�z�5�դZ*�$d
��[���4�t� ~� N�B����Jǟh�*0����Pګ�=n'�~�$�Yx�KE/A��[�"�#w}�wڠ�s��7NC�zƒ��z(��܋�s�jCM���I��ԕ�ܢ$ء)̸��w�zw��BJ�bgG��7<MXN�hn��`kW���*1)�a^y��Ckj�gZ���+ �Z�~lP;���=n$���6v�eb�y3c�����"~�4���RV���PUm	}ϊ�^�����ڌ]/3L���N�U�t�h����֎�qɀv��I��7���Ls
%[�%N���hG�Qi��n|3^�3�R��5�8�gQ���f]צ��#)NJh�Dߏ�]K2�,���쩻,�r�.�u�	�#�)�9�bY�	s���W���y4�"1�W�[�����Ĝ��[(%�K��'�ƥ_���E�-�.�t����"E�R�e7L�p@�&��ƿx�n�" �����u�J�xqYk1l�-F��Z��@H���.����*Ep��Y��aυ�^�������H4f�r��u�`���h��l*�s��2҄�݊��>�8F� ��25��$(/�xkS%���HQqc���R�����F��C~<��g,a$=$����)s��/~��L��t��/�m=���7����.�;�_��m� ��"�5W6�f&�%���Օq&r�upN
e��u�"LC�5��nrp8),g���]��w�4M�P��j�7�뺵X��Z~��-��i:_���_��O��C|ݩA�:�r�!�I�x7$s��Ɗ^?�vY}]1N��$��gm�l��?����@T9/N�q���<Q�",����ݨ4{1���ƅ�.g̯!�7�s�0���q@G�N�PR�؋�+�2��U�G-F��#�5)_G�_��\�N9���c�G��|8J&�V��UʙE{����l��c�t�,ר%�/D蛖��w�YT��-}�m���aK�I$Kh�U�Ie��Ư�i�RՍ	<���?ޡ!�����`�	��B	�5�����|:Q��4ُ6�}�gA0��c�ǙZ�Mrǉq��Y� �Ew��tmd�wb�N�N�AG��{	���)��K�GiR���߆�����ŨDDAM���k�:�������H�v"�Q0�T�=4ӋڞG��rH�5�]�|�D1~��K�ؾl��w�96ns~����X����-u�\9�"�D��xc�u'S#(�>��-a;
� o.�����k�������]쇎t��p!����r/4�����v%O�.6*J� ē��ʙޖ���>#��7F��~M�0ͩbæ�� ~����Z3��?l9���>&�e�,��������la��i�_����:D��b{�H�������ށ��E4��x�5��W��{�ڬ}�B���׸��>w>�K $�y�3�p�L�֛c >9א<r>Wͦr]��N���ѿ��� �hW����z�	��~�	9�|��T&g-z�.=i��݊�KÄP�X�d��	q�t����yol+Q�y��/�������Z������bȤ�) Ģ����r�u_r�ĴlP[q�#�T��@�mh`��~g�P�O]ǔ�2k�2)C�g]���f�S�}��y[U�N�������`����V�U�bە_�T�gѵd0�o����c��(��ջ���V�q��2jD�d��"����^Îsy:ŜZ$����'Hu��T<���8%�M�/S����u
u�2�<»b�Ã��~DMw��ͼ����5����1
"_p�(����&K�ײ��ֲ-}��6~�~x-������o����d������Dg�tv�ґ����M?&g�
V��w�#Wq���R�J�Tz�g����ӦPZ������|C�b�g�^��$7�$lx�2J="�a���@�V�<�2<�o
5�&9��v+7*��Q4��˧��ma�8��)���$�-�/,Ì�(_�&�Cb:0����"����
qL��mg�9�� ��*��H�\t<���k�� ��Q���ޥ�#�O����M�+_x�4�O�\1�S�
��BX9���{���#�uϫ.����\+.cl��5K7fߦ���0��|��Ft<~�Ħ�MWly`�M��t�C��K.(�چ�\��M�s��n�QW��Ӳ1Ѧ��q���m��M��\vs��Jb���-���G�A�K��j���Fbfo�e�_h}Z���d��
���} ��w-S5M�\��ȴ#���2�gILUQ�L�x��MC�P����w(������" , �:3)�М��#~�`����Z���9�򍶫o#AZ���Ү���­YEr�LI_�A�
�C�nG�������vS��JF���j'�$Ϛ~�A݉r����0.+cE�^��!�Z�Jd�p��/�X�>↹�3���/��s��g�ZR�x��'�7�+�f����ő,�?'`�⢗�ߚ:�����~B��j�Mz�y��b�\�<֡[�N~"�d���o�F���Sn�R ��C�����A@�!#�h��L��q�ߏۍ��0_���*8��
Q��Kj�����/4���Z�f��%ŷ;�2��w"*`ܻ|���F-�K��C�$�ƺW�5�������H��뱂�߃x:,L}�HP�K�Q������ǟ��,�<^/�^����P�YCEP�� �Ci�ʯ�`'�F �*DL���E���y͗A0U&��,���m�\�8^FpyS!?��f�^o{�K���;���N���[��-~��`���;[�����*Ko�8^rR�]��"Dc���y�F ��L��8<>Q��1R��l�F��d&�h��D�Ƒ�)�_�C8����#�o�=���k����2� nR����&�W�Fҝ�~G��tZ�)���c�Ƃ�̕}��I����$�3�i�e=k?pD������Xkңɯ��Ak�c�,9d�?�ys��ꥑ�5���j�����0�Xsa�#S���V���pj?�)K8B�.�j�y� �ŷ�v4"��8�)�k6��ELG��*�Hڄ���~�>�l�+�0	15_|�r�ق�<����q��s�����GC=�	&A76 <Ew�d�k��ƈI˚P%Q��x\�������PG�a�}��@\-@4q
e3.qa@�o9]���7{}c�;O�����������[�t�2Y� �`��t��]<��vwC�E��2���4��|=��ڤ�0�"�x>���[<�^4�`9��w|�v�ء��]9��L
�c�хá9֘��~l��n&*���Q�Ug���js\�\h��h���aǍYڞ2����ۄ|O^jʴ��O�)���cO�h.my���u+J�E���7�����t%�9{�W�F{]|��H_�F�p-yܓz�F��Ujaj�wI�C�lP�I`&u.g�� �\0J��E��uD�����8Q��B�B3�����ehC}k֞��5'�Pk�i�5���_�=����ğ~��a�&o��U	6 8GU������)�y�ӌ7� ����$�T��o��=�aF�/0!r>�D�7'��?b���_��-��_{<-6^P�s*q=����W�-X��ڽOX-*~��N���q���}�rq�ǟ��uu�W6C��ێ�l��,�$�M˪x�h��J�:2�Dֆ���������4��8K��[G�����:f���a�E�Np���͂{����l�s��gץ^F�Z 2�&�R��dQ������RNvڗZa
t�c|	�Oh(�'��h�c��@S�C؁y��l�Q:�;�P�a�����5G@Y��f�iC��[m�T���xƋf��ax���A����(j5������U^�c����`�� `;$�Z��T�\\�{ׄ�Gfi�ؐR)��4h��`��U'g��yͨ܃��۞�eU�D Q�\��D���Յ��e[��p�
�*�E�ή��VzL$�s��'�f��.�Dمoe�gW(Mv�=�T��v�&�99H|�q'���r�4�󧵦��aG�7�5����j�����rU�%���:�]�,ɇ$�n�r���ʺ��iC�\¸K��"!jB� 8�4#^H(LNַ�~�`���du�5Z4�7v�2)��$�E�W��1�p��=E��Z�j����2��Et��X�vQ\��6���3���
i1�/�2ix����dXH�I3�/�'��	���OW�} 	M��Ŗ߯Z��	I�Wp�Z���h~ �����3�Hec������m��O06a����+JTHS�z�`��N�bF=�n���'��*��A4��=�x�p�w���9>M��S[wE'˕��#��H竟���	iT��y�NC�7!���yT�(���B-��0�T�'��@�&�!͕�P�L��9�fz��<��g�
��|��ދ��N��z��i��'�6����Kkot+�x���"@����M?j�BC��})Џ揠�j�)��D>��\�zdAA*[5�m@�4l*\i
�N����K�X�r��&���!�4ݐH&����P����&��/z�|�^��7d!.�B�e���2K)��q� �$����d
j �N�ˑ��%[-"��?,��n7�
�$�۩�Xˀ9M�GD�3��m.\b�#�[�F�bS�GLWd��A��h^-m^q�YSJk���X�%��O�|�]6ګ� ~MQ���߬rgW� &-�\��Mh���PvzQL'����q���Z�3�+J��#���Wr� �Ufz����T�&���>�#��:�@T��9-�E62+O �n*��Ø�gEx��e9^m� &ت��ۅ2o+��rd	���؆�%Qi.z�J�#0�짩�3M�o+�)k��Ag���1?TU��q��~ųB���[|���>H�Y��k{�ȽS
9`�{�JbGm_�㗟���
#�
����;���$ ��C�T��M;�����И����	l��	h0pQ�T����l�s܋��^K���ct�X�	��.��U�L�x����h%�8�@I*�m�R�>�d�R�ݬ@���rMI��k9���B�l�	���D.f��D��������q��'�w^Dc����������Ѝxm��j�NRp/�՟�L*�ar'���Av�*�0A��3{��˧ Y�ȍ10	���{� ��wf:�(>՚PF���w���~I$[�1�](����v|o�L�̰���NS��Fr�bΜ�k�:?\�"��[L&�J����T�����;�G��C�u��ȭ��ƨ��0}�S��(���	���^;�Mk�c�p�F���Rz�8R�����uN��S���P��H+��}_)����|&���<�G�:�-���g���S����I˴kf����Nۥ�I$��8,���$�,%��+eEkȞ�����G�ѡ����͢��^�c��2؅�I�a�5������IY�߂��E�g��ܩD)� �C&�ը$�_)>�>C���7��8���^rOd�N[Q �tι����qt��%�ɍa�DW�A�&�1T?�ImE'Z��D�ȯs�΢���� z^����S�=�|q��f�DٳX݋P�%�	ز�e��6�k�⼀&OO��F
����9(�y�X<N���� {�k��CuwT䦫�F<.Wo,�O��{���o��?.����ف��^��K� Xa�O��G��뒘Ju�y1c�,�+��m�h�0r����@���m)øu�����5�O4��~S�M��`Yy�~�#�Vs#�b�n`07���jo`���ݭ3�)�{��Z�[�X�z�ЙY��f��*h�Gi�%ˑ��F�5gZ����Y2�3n�8 ������_��ٚ-+����=�޸�hϮ9bO�(iP~$�� *��7�JY�KFH�ō�r>0lA[ �l���@-�B_�J׽T�@�C����tL�yy��-���O،�jJ��3P�<^,�,M��Ԇ�,.�%�9c�DbeS4��o-��˒t �a ��R[.1��� �����R/�\�r3�Cf���%�.�'�[�6�(~т�	��A�t��]4'��@��ԕ8e8�,��*|��Ja!T��&��KX����{0?-&Qv/���vW��v/�/T[nK�H��?�ed	�r���#�=�z�]ƺ�����3����9h���K�����S����W@ �Nxb5���/V��@w�s�@ו���a[mog�̃֠x)�s��\� �+����r"3�*�![�9w�Yz�í�=~�R82?�O0����q�C��6*1�Ө\�-֭7��<�o+'����m'��:nlRK�/`&ۂ��6K:�Z��_)��0ןpG��lH�:��|���6L�*(�������Q>Tсg�,�ቫ��)�e2P�%���$�zǥ*�y��V�_;�=�m�$ݥ5������K��~���_����N@
O�� _΀ #Y8�\�s��ܗ��R<Bǁ���!���[�ށD�,�q戙�M�����|^������ ��k��Uݿ[��;��'�	 ��R����CO�{��@�ϤA���5��&�yF�L�O"�}f2zs��7�\t�<'�Ց$�ڧ�g�.q�U�S2��U���t��sŇ�&r�<tQ8T�Vқ�Z��e�)RÙ��/>uj��N��b��*+ֽT?H�mR��O؃I�ZQ%������b3�N��1o�]�ʿ��Eqx`���Qu�h�����{ ���Z�vۆ���O;k�TQ�d�D/����$��n8���?lyŇ�j�6a3$HRN�w�}56��Vh�Έz�[`� ��B���{��}8�Ԋ����A�n�'f���5e������2�k��[ ���6��C��F=��)��x�zӢiQ�1FU�	�RJ�bM��] }ae	�-�8�6��^�N��g��kly��*g�K}���"�En��(�j��~V�NrW�:c���t03�=��UE&ۼK�-�+?Ej����pK`��Z*5�l��xJ��q�8�u��.�J�	��NR��=g(	W����qc��P;?ӆ3Urߏ��d!�]{�.��?��J�1����jp�@���>�\�7RЎG�l��g�T���j��x��n !3s�����U'g8::�h��S0�����l�Ō��pƕ�GW��j)�#�#)�7O��]:�1��u���:9�������v�kg��P������ÇC��ގ���X����4g�T6/u�G}��-Ν<#)9]y��{:��^�6�J=���H�H��N��Y>\d�Ԍ�վ��by�%ӑ9л~
�-��cc��Ih2�b����$�׸�$~���J��O�Z$�jU�1��w�Ecc��OVO[w��� ̦��`^�e�a.'�F�zT��*Y��.&��p7����I8����P�j1~�JN��L��#H'&�Oi���D�����kN^��(B�֑k.�/��22&�ثG�O��n� 2`���22W�`�AgfL�қ�-�A�s�{��n��o�X����D���Ќ�Q��W��Q'Yk�ҀC>A�"���\�4lԮW�"G3H��1X�k��0�$ޝ؉�z����K$��s�l�cia"2���8�<J���6��\�����톊>�����c3�~>W��� ��<ِЍe�`Oaqf�ư%�����n����E�$	�$lh0Xͦ0�r���%�r`��������C����=�^#�n�)BO4��7��*sI�Y��9�H(ة�J�Sg`T�O�'�@�r��WRemާPY�������>���ys֕!�-D�}������$;��{���%���Di�ZՠՂ����~����0�¦�|F�-Z.��y�{�U�)�5�gk⨜2��&F�W"R���q������Q�/zѶ#�6�D)�4�es�\NTs����Xۀ7I����ܼR'wGm��vM5�q6O�P&!�dO��Á���z��(1U���iI����9=Ҿ����UK���V���w���m�X��:%��	g�"O����L��^gc}\�Q.���*l������+�����ClH4
�^�L���g�Z;�v�]�T �t��1Eً
u�XE�y��:����˙��OF�AB��9u��P���z)|���B�T
]P=�������p�ֆ�%���K�����,�^�)�G^i�UiF𣨋��e�C�4�pn*�|�6���ԃE��
TÈ��"J�B;Mo�M��y(��@�%YӛX��xt���Ù<��}���37[�6��5,�։�%�˺������'fĆ���AA��5�
Szb`��D���h�q5�]�p��l��f
��q�4m"��ta�H�`����e\��#e67F�Pz@V�\��|�h�� ̄�AY�����Le�/�a�<}k�7�y"3���/2C�<�m�8�0Os�ޗ�F3�u���	ڎNV0�@�kَ	Z�`�\Ȩk��{9}I�[���Zm��5��3�����Cb���#�w���I\o���v�Ρ���:b�`0|�*M��tM%iQO_�/F|Ue6����^;� �4|����5��A&�T�R̋���	�Q�ꀎ��E����bd�ꛚ�Z���Oa�v`�Cђ��V B]z��^uI�ē��#	��;f��>�����T��ZB����<��̆��v�����q�_��(�[��$���2�Y�8�|��5#�-��1Xx�8�ji%m���q�Z��[$�%�T^�hc�pէM}�x�!�t�'��_H�6�[4�?45��]��2ppwn(��K�~�4Zgּ�&JQ���`npZ�*_7���I����4��,2��C�ه�d!V�I�w5���������2�lQܘ�S�X����~-Ȱ��')�(P�yɉ�=��W��0��5��������D	�~yf�>X���V���<.�?=[�Mss::��*�j�����6N�.����� n-����$3[4�u��m�[�����2��m�}|n �Tl�����[qNPs�[M��;	e�	��sF�2z��V'�7�D����vr`�~�X��6�R���[J��?�X)�	�s9<��b�PzS=��M[A�@S27.�Hwc���R�>hPS-�k���lu��V�� 10�og����xB@5���C79a}�#v���n��\��N�2G��9}�c`���@%��Ȓ�L;py��ѥyZP7N׭�N>J	�)�Cc_K0��'m�z�'QKK��/�L�	� �(�z�xu>�3�Hk-uf[c _Y�|aX��{�X�St���^ʧ$�C!�w���E�æh�xB�B�):Ǳ�V�TcViOaJ�"􋚲�X�1��_|=�]�b���<c|~�1�\d�m��<V<fO)���M�4�ҹ@�Z�CӅ'�.����7��`����K=u�V$ނ��/rjLq�DW5�l�
@��\���ć�ܞJH�W>�7�}���߹r�h*lK���O	����]�e��պP�r%e<�p��x�`*���	�.k��NQ[Llɖ��Nn�P;s��>#d�5v�	`
�qܼׁܜf�"꘭r�R���W0��E$��S��w��Ap�x���e�Yn�@�L��S��?3�O���DJ�!��k��5쒞��W�8K��m�\����Z��l@���Ú�#ۂ��!U	�還6VI2�ȝ�z�z�h���F)n��+��9~��SFr��X;��&U��%�5!��Ȇ�y���Q��?C��sB��A�JL ����xt;7:i�|ʤª��DO})a/�b�g!!B�W�@�I��n:W�G��,�(ѹ��\Q��F$1&xSE�`o(kZ@��3�]�lm�a��s7{�'�n�����8Oև6��5m�����>+��s��;�Su�h-^��[�f����Ј��7�#�{C3x���Ղf��mw3~���#�.�"���^���Ek��/-�]��Qz7
V`�IJl��8��,�S?dS{pԎ�y��˪oT�v�)�,��]	hX^�j[��L�����ѥ��A��p=-����:���N�cƁo��Gr�@����$㹭c�:�Ҡi�O��lh��K���DP�S�U{W��FK�O�8t����=��m0�%#$����?�y�v�o*�Õ����I��Ҵ�׹=��_W�#F���Җ��m�(bv�4Ө��ߓMn.\4��S���0P���m<������3@��}�"Q�o��s��G���yd�vĥ�H�'���^�	{`G &���7�/&�
��j�6SZN����o�?���;����D�6�{�
4���L�^*3���Ň�6��WB<��e��]0���SGW�,-5���_�̩F��PO[؅�=!�r����g?��%� �ryC#
G%7+��H9���|gF�n� 3�n�*'!)hh����@�C�ߎ���#	��S8���,��h���b�Ľ���ח��
��cgw�Y�=�,�Eo���M���]@_pe0��p��V���k�b:�L�P2�!ٟpf�Ȅ-HnX}ܼ�\���`�O$T��¸�C=�1�ˁ��x�5���}���ui��T
�\f�>�k؅�J_��}������5�����J�sm�
iY�V�ݗ	
,//���v���A�âa��!���G0���88(G2,��f��C"��m�A�I��5�1� �A��M��2i��� �2D֗����QZDyaIǑ۱�t4��p<���,�s��1=��N=zn�]�J��D�́�z�w	�+h� &��G�i@�6'm<���Āf���::�b���HO��o�ՋRj�)�>�P��ĸ�2>����_wy��
b���g,��IE�h�o�[K'c����������Ax��.�~"�#4'�|TY��ۮ�������*$�­ʄ|l��l�R� ��"�R��:u�p����(���@��¦o�&�~��[��Pv�Ŧc#~e���&�3��;�o֗
��>���Mq��$L�6NH�}<\H�{a|`f9呈���U�QԴSҀ
��g���[��~K�g+���'N4Df�~ �����?���O>�ڴfC�7��5�Jr��t<F��J�'�;��3��L;X։�2�*?�~�-�؄S{�CGm�4:��f�H���p�u}��<�~{f?�
'�K$+���l;�	a�l�I4B�P�嶠���f�SK0�4�֌L����Sܢ�x�mW|�:�Fўen��|�TҸ�s��� ��(��
��Wx�������3X8ɛ����ƈ�5 ��	�4����L��%��;g˶��2ܛ:! ��Ry@+�@��>-#����t=�����l�8��	��P��{��X�h�V��;n���p1��SeG{Pq5|7�G7�V��=W.�z��a&+��$E�[pŰ��j���Ci��DS�g+
H�7yGg� �a� ȵa�= -C�S�	�ֹ�@J��NB��	G)�)���l��Δy4M��mc#�v�g�@�zN����f���;�,�u����@��Z�@l)�9{x�c�-]������aM��a�����>�g'�&C��s3�Z5~��ґ��̋��jX_Z:�����~�p]ygb�����:GDbc��a�N·�EzӸ�B�����Ҳ�b&܆�a��kk���a��R�^�;�9���-�&7c����x�Ҕ߀��"��#�by:�*�$:u��p���u���j��:|�i����,6G�Y��I�z|�������lf��/؇ϻ��H�B�
u��e�R&�$��nKGVp):0�e�j������(�^��|�=�6��W%ϔ�O����x"hA-�w_�Y�ƽ�kz��n[�9�Z��"�&�Ƕ��d���c�-'\Ce:2V B�L^3��-����+��D�������)�恅� xLl�7s��4<�G��j�l�U�Jqټ�< ��sNɔqsK�C��H蹠^�<�;����И*ϝs��E	��	�ܑ���r�|�(i}aj�{���<�L���+p^Rݪ��l ��j�w��8[`� X�#x�2ߥI��.L��E�2E�L߭���g�v�+QTx�F�ʓ���;k�y�K��������D���*<z� u����h}�z.��Q��=5{���y�+vO,���2�4B-,\- ru"��ց�>��Y��,Z��һC��Ҏ���� Z(f�I�p`�������MU=�K�``m��a� P��y��X�P��J��fy(�V��WȚH-������`�v0o /#�a̋�������h8�d#���N�6��)��J<$�M/F ���������y����g����=�I�ÑR��2����}A;��q��Zʲ]����<�Q��rF���d�#�>�]�s�H�u��$6����6%�k�M��fs�Ih]X�갦�M�k��x�L�k��Q�>oRz���F��	��֎�y��p��u)��f��fP�6�U��_tlQ��@��Ld`��6ṔPB3�
@"{R%T9 ޝMR��hL�U��R��\vc`����������dNyW"�����P�58���#6��6���OM�1߿��)*�3T�<�Ki����F{K(Ћ5.Q�����%�a���I�a����]!+CoFR,�箨 ��K�~��5�W�tpb�ӎ勽\.�E�0��հ��E2Qĳ�I�I*
�D���0�Wb�O'���퓪��mc�W7`�N'
���c왱M��V��f/j���V����iVt�<���9�A!����çd�1@�w^�M�CH�͞&��;����A[r�����i��3vl끘<�%jƌ%��\��;���
C�m75uwOgWf�ꝡ��D��2�6H:Mg�g%��4��)��/���@Ep''��~D�ԇ�X�[�"�1+��q�es���͂.�)�>g3��'���
�JɃ��i�8�$�����%H7�0Y����B�{�gBYZ|���7u�*�\D��������B3[y�d}\>K�|���Zd���B��8�g5�Rt�����Rt�� ���*������H�.�4��F`�M�(>RՖ�����Hw@�=��v�hԢ����!W��u 0�K*�?w�2B}(�a׈<e�v�uJ�w�ӧb�	?����'��2\vE�Y�RT�/Yガ��UgH�����oFd8�%Q��!ܡ���$7�Ќ��-����30��D�xÔ�9a7-`�����B���v7�xp�X'�t��U��8��&-:yŕi־�\Gc~�����_cr�r�N�#[������0੯	���� d�t�����K�\{�Q+��Q|�G�
���~��O�!�L�,6�C�y^�Ġ&�<�"����FCh.v�ДP���: ̛P�_�㸥˶x��@��������
NZ[��4F3:*K�>nJ��BBl�Ԟ�1��ŝ�_���f�K�x{��]TA��j�� /t�ک�v���t44/�ZO�ijnh����[>ޮ��m�O�"li�!�l���"�����m�-�X=�ac��b�kp�Z���l,�?�y�U�>����{�7�E���=X��� s��)h]����n������T�h���� ���r	����:[�A/����'v�Ʊ��sx�ĩ@b���Ӷ�:)��	t���ٞ׿5�m,�/%=�9A�$=t j�t��M�6+W?e����[��B��HA�h+�4�Q��Cm￐`����
6P�b�m*��������Z�OT�m�1����$�^w��v��4�US�
�I?uz�vo4ew��I��\hLJ���V.������E��eM�����g���'���td�P2Ǡ�;��=Z�O��p�<Y�*�9&K]��5��J^6d��*Y����JBi[(��|�N��Y����>��K��T�Z�� ��09P���?]j��˸E�ǯ���!#�Õ�<�|�@��[�È�.��-ޔ��a�Yj�"Q�����	t_/w�w	Q�{CKJ�%�Ўx��������۩���j`�I#o�����A���	�j���2�{�8��2��+%��,���t��rT9+�Y쑆��3Cu�g����� .lū�:�[�|��Jz[�l�"�׆�u$8�wx����z�[��A�����Ky��\�B��L�7��W�7���Gh]^�ZV=�B~Z!UuT�MSW�9�?�~�S����HN�߬?��Cfq"nI��7~��c9fe&6��_ m��XY�e��8|�z��Ң'�s�g�n�M����|J� ��XO1�?aᒎ8�{ٲ�	�SM~#P>�ߗ�6������5\v�`.*L�������at�����a�� ��-����J  Չ�� Q.�e�3�FJ�?=�|�D`ۺ�g�G��;e���q����/eW�.�\���k"j�5��T�lE��x^�{Z�8��z�]b4�/R��9j�K�H27��聦/\��2���`DO�Q��ȼ�ԋ+T$cG����<���uD�����ʃ�������w��������b�������f/S�hӊy�[7��-��< #�#n=����)[><K;w��I���r����]��g{����H���m,�iu�:VgI��68�c]�@��{����z��(�/Y]Q�d��nJ��<���#M5;Z�q �9��RU)��ao��I|��6�,�1a�*D56��F��m���9�ߝ^�M�y~بƟ�񂄕٬Q�1�#ˀ�+�u���;�k�ɥ.͸C/l��j5<Hx]9�
�Z�ĘA��6gH���\���p�^I���Ż*����?�-Pp�%g�3�{���i0C��='��Hk�N�%�_bD����ۮ.�]���9%)�W�k����q<�y�:
$Ts�� �:Y<W�e���ޭZa?uX�;�x��i%�]�U�A�B��j�B�;�<=�ˠ'a�6i��f�wa��ީ@a3ָ�;����B�@u5�+v�5��웜�$@�-p�×}�������π���`!�)*g����d�І�B�3���G���?��N�iBR�yi���5ےȫ�4�� �`q�c��؈9".��'��:�KX�򴉶��TH�ͦ�i�3��cOW���WLA��ۜ��ܠ�>`�����Ġ����l�)�\w�~ 4v'�F��-�F΁=�\��;S�.�Y��˸���7�!9��wD��L\���)�����(�ŕRo�jFA�gx<\�_��?��=��g�G�.�p��	I�S��c_Ŋ�:t�=��S
�6W�#CnKF�d`2��;��5}�ֱ>0�}긲���]ӕ� ��s���x%{"j�Z��9�Z
� �#On(���h��-���S��f�^����x��N�)�꽍�R�J!`���ZlE���^���.Z�tA$�uq�D�5Dgq%y�.�JڹF�"/���JK'���%�;�?�\c�A���#/eFҨC"ߧ'E[���n�e�a�s�;v�x���)�r�}�����O?�V���R��K���s�H� �O%�@i:��D)V葾}��u�1�g}���ž�@�J�Cp��?E�@�>�i[��#��������+Te0�K��m���i�:�/پ|�s�OeZ�+�t+�"t��K�V/v�:v�/�v�.?Bm<�%0{if����?%LWt��i%6�ou��{���f^���;�X����d������Cn<�>�X�|t�CpA��pŦ?N��޾�o�r1��$:���n��R��4��E��+T�u�bNً1^�O��ɛ�KX�-	��j-��hg�^��}��'�}V`p�z���L�����EUK�Z!��,�O�� ����q�qoSz}�����A�=�U�}�y��{���~C��2'#��=���.j�o#*:��!� OZ�\��국���9�����A��k�"f�x�) ^'��y��ж�8R>��oF�@�M{t�E�B*�]�[P��N�ڣ������M���{y�=	J�=�S�*���ɶ��HV�_΀D��~��ac����h�y�E떮'�N-׸L����3p�>���_ �S@#/'EQTX٢ �u�GM��Ot�(=���S�yn"���Ɛ#�'���h�Y���і6�`�CY��@`|��t#�6��
"�t�Io�U�;�WN�*)��BO��^΀z&7'୔����pnʊ?L��'O2X���R��v���-�k����?���LK'�1_;~\%1�4(wC5RM3Or�~X�������&;��3�C9{����Nw�l�u��B���f�Ck���H7	��zl�ү��.������F�l�}!$�w��B�^���r>-��&$2`��BZ��F�q���Wc�ʋ�x�D� b�2�f'��>�m���N�(̥��G���d@�J�cY38p��2D?-
ޑGqcr���\��K�o'��+4�$�i����㖄�6_]w�N#������j,�֪�p�C��f�+��ڥH����:�>\���ۧ!�m{i� �	Ҵr�D��I��)��#6���=k�j���1}�X����1�vv9$3�yV�_��p�v�9O����t苣[ٝO�핈��A �*�z���c��T�,9ƝRrp��v�O&[t�9�ĸ FL]���C\�5���5TM��z�;�	���PӇ��`I��y���3!w�S�mgxK�q�1�9?8�3��'�M�,���d�p�`�(��ߖ�݇U׽V6���L�L��Ϣ������u�m�CU��0��]�1�w��Ĭ�#H�u�0W<�O}�����@h&��0MN�6����f~��w�Ul���\^E�/ܴ�����^�,�Q$�J�)y�0[e&/*��
�OH���6j�Iw��C�FiN[O���w��7�;I|O��G'�1�z�&H�H�XX�N�����:.!�I&@��X���g�+�a/1��0��R?j�y�d��5�)���B��ET��ܺ�n��iO`�Eס͎�-Vr����K?Wf��?H _.w���ОW[K�x���g�ȍzL��Is`��ͼ%��H	��Mf�]�}9U�M��'�S�D�O����b��#j�%6JJ���&B�>�J�&��\�~H�$9`:��[��ʿ�m+w� �H6h������V+)��-�ح��J��8sy�7~I�����^􇑛���Xj���� �;n�gy$�#Rha�SUC_+�|�N�m-I���Ù�uG^��*U�u�SE՜a����1�|V'�A���j��N�&�����&x���R��5!�+9���8:��t�}bN��B�[��%�cv=l�9����%F���%�0�Ga�����XÑoq�����?�����>1ݵb�� ƺ��GK"|ZqZ?�B���	�B����8z���%�5p������98E�s�����(w��t(s!�[�>�R�I�87JAՁ.Rtc����6A��e�t�C�y�7�pL�l��HDڮX"�Y�{c�0­ђUV��k�]���Ŏ��vN�f�P��8/Gݜ/4�
j�H`�V�,fW�W�7Q�@<����2#�~����k֢�x����i��i��!_�~(aqt��C̴H�i}��}]ݧ _1���f!'�P�*x������<aF/?p��tvLi��rA����"�;��&���}��.ھ�ݰq��mk�D�=���Z������!�zc�7$���lwu�1C���y{�<H���=�i!�XJ��T����H�k���N���8sθ��*�A���U1�4�B��'�b�GX����l0͜z�&�\��x�l��ngM�s����;�64'��'���K�#s��6I99c��x(I���bM�£�ݎo��}%�a�@����u���f��.X�R,_Cw_^D��Z�34[c�m�a�ҷ�v��h}�����ns})�	.��pⓛ�-�bv��xt�r�D��`#Ѕ�ӵ`Z�hJ�~j~�
�zL͜5ֶ]ЯM�l�9؃��O�<9
���g��{����u1����3Rĩ �]?��l��4�i0薲5u�w#F��,��t��.�n�; �G��%���1�k�a�c������i~F`�1�4B��s�S�/�Tj��d�H�o�1T�1�kℓn�YCa8���`�l�Y�ex��r�u�էu����ֵ`����̈́x���t'~������x�� �--��[;c�L0��N�!L���E�T�o,����e�+�(mn&HG`y���nvXN�i"	Ӿp��v2��)�2�)�T@��� x���і���4��PW�������[5Rq^��?�����P��ot�$�B�<��a�U���iقb��~L���Z������p�F��Wn�{s ��CFf1$�_���Qz��@�iuk'��/V�G�e�:�Ǭ�0cQ�M��������!���tq��VY������,� ��YC׊����l)����yY�V��8���"U %�������E���b�.0�u�p
nO���2E^e0b������w�<g�ǲr�sN�m�-�`{�SX��ضfK�.�c>�̀�퉂����zĚ�C��y��@��x��; �c�k� ^�_c^�z}�x�"�σ��9���%D�B�u���c��:o�3S�|�E�@�A�ҍ�P���3x�E5ћո��W^��C�8\I.k��)�@
�%�>B
��F��)]̉$����/ђ�gӬ1�֜C�xd��U��R6��K-�sqƻ��rI3F(�^z� &$,I�|��n�8�'�!��1��ދ;s��<!YC�/i6�ޠI/��6K5��j�(R��
�Gc�ZDK����-�������g��c��1�,id���C1�(�J���?S^��i����y��n�3�Ŭfuf��Po2`��ݧ�3?ӊ�Cf=�޽�V�60���2Ui�w��AU���D��s��Q׋��#ـ��u炸�G �R����Z����:�\!�B}��;)FR������_%�� ��a� p����x�'q��]d�4B�O_D��L8�Up��6n�v��s3�TRX���D����U�.����"�`Z���2 �6RY2^��Q��%`M+Ņ6�:+h�:4��
Ӈjh��@}0����C���իg�`���1:���>�,�\����Hb���2�b�-+X�SJ�)%Uw\t�H�Gi�	��&ܶX�|L!���F�ۻ��Bt���`�h�����{���r�v���-H�}�L3t�S(�OS2� ����`-�1�|�O5�E��#<#$Ex,�g�U2py�0� ��;����4��X�T���0Hb�4��l[]k�d�5��L��<i¦��ĺ��k2]u	�95J�8�Җ[X'F�{
��W"�4�
1���{�s^`�i���@0BQR��2_^8�<�/:���#K����;��},x"��F_�jG]k�~�dZ(���'���z�1�@/A|��  ���
��&���:��O�0/�<�d���s᧦�����Y�jV�,_�Q��`4������i�=����Q��c���4B��� �}-cֿ8�.�.����7��1��?��Jpҋ�M��H�Z*ܐ�"#}-E 2�˜l�̸I�����g_��-�\�&��(H�@�a@��z�a	]o���}��x;� )�:S =;'t�b�m���N4S���*�^��:kP���B�����b���D9��UqA��s��X{B+��Qy��a�����j��X$�Z(�������b��N����MT�+���e�Td_a�&F�'
9Ha��Z���\ Ś;�ɭ����]�h\%�	�aΖׂt�Zw O�����h
����s���R΄��3��[���M��+x>�[(�HH������P��侕b,2u'�Cy�J�KL8b������dq�+�����Aw�e:{�#�H-����\J5��;fz��
*^	��t?�.��.�������?ƃ��Uv�t�|R	���qk�
��M:	��ƠGi2ނ��	���h!ʤWov��g�x�~i,4�R�Mnґ�EWt�}Y~�lg/Y̏ �B�������h��ӑ�F!�n���&���U?��/��x�.�(�@�����*�śr?|H�R�����#�6��D�ٶ ]�y[#�Vr!���=l���:W邆�4��?�m�O��Bn��OA=r|�5C�E�by����h�9ᒅ��uR�F����V���P���N<3��{]Z7�"��j��6�u4k�]?��
��?+L��X�f�e	~_�$l��]y� X��8��vc�P��U7��@�q�u5�>�q��^�E��4�$�I�W}-�o�m���6d7��n|�F��zJ�ıJ��lj{DW��*���$�"��r����a��	���o娋�2�D*E�"ݛ�r��+�-(c��-B>\���k��։��El��(�ڈ��`H�$*3"�!������vmo���Ս2�t�]�Y�Ί�j���v�JPW8� ���Ԓs�	h�aˎ�tX�\��f^r�&�{'@�>��f����"X�y)IR�Z5zC���#q1�� ���$P��"�v���E~��Nb�1���-�D��a�B�'�D�iO-D�;��O7ǹ_��Ә}W���j�礬�]J�W?k�ɓ��7��F/��l~'3�5XU�X=�?�o��< j	�wq�C���6* K·�'�&HHP�P='�U[-V��<���ș5k�����Ro�zG=��pc�8���ߏ��Ѿ�������]���+�%O�NhN����h��9�k0�꼺`@y�����.,�.d�+�B�5I�DB,�����VO�R��'��ǚ�\=w�<��̞�`U��H���JãtԩK�G�"��Q�ƫL:P��r��I��mqm� �)���oTW2�@KS?_��Mp�H�aF{*Q-Z�b��(oHŪ��Q� ���v-fV{���r��fjP{��o�w�U�v�+5,� )��D2OeJ������K�i@Є�Ru�i��_&Ù��a�{���=�F��k:4xGȸ\��L#LlN��$�o�/�+�������%P�4׷���l��X�,��%�b\�ï���9�!ԅ�a�@9��aY�1újuU�=2�OӖ��z����#��5�l;i6�H�QCI�5���2����r�S|��:�fV�c���o�G0DV2�F'��B����q�W�(���]1��H@!�N�p��
�;��ҍ���5�YSVڪs���.�b�-m���B��1�;���k�2;�0�6r��ǔ{���Q�Q�Ç�Ԋ����O/||J[|*e�)X����;��$���)�E��*���v{]ܚ��7S�]��7RT�+��Z���+� A�%�NMz��`� ��'Vh9�}�f�hT�3���J�7}C�⡚-��-CX��1���673},��q�~�(������a�/�U|i�E��\d��0�i:Ww�-��Oյ�j�l&�[កO$����N�)N � ���
,��Q���V�7�g}���;��5��П�T֝8�gO����Y`����h⶘NX}�$Z�0|ECS��˳>bz������(��>X��vP�N-�l:�ZȨ���Â��#,�����wB'CX3��:p~��5��x�S:��P�A_{E��ͨ�|m*�Sx�K{���Ϲt����@�h�X��Xz8a��HJخ˱PjD��Er�)�2�t��#��-��Ji�d�9�����=��f./�B8m~�*��&k+9|�s'A��ɺ��VJC�{غ�?�F�?>���E���Fkڶ�k�nßx|2#2W��TG��OQ�</U^'��>z�p#D�H�����&4��f��m4:�����_�:��]���W��ЈQ-����BWBW���Ъ�?�{5�zx�uHqs�6���$B�����M�|�����[X5B�i�Ѧ��D:!�:�c��O��U߇2�_�d8pBx,U䗾���Úg�W3��2��V��*T�u�}�]fml�n�cR)ꆐ�I$]���	�:d�����p�e�n�R2ӝ�N���v�K3�<�lI)[՝.{��.N��s@�Q[o��րr������FK��x�%-.>KA�D�3X��ک�
 �����J�{�:�W��r#���v�Ph ���L�~�m�8)�G�vH�5�YIY��9��6����	����b��0K�v>��x{��V,���7����-�$�B����J������j?b��^_�>�o㸦��`�&��ؔV�x�V�ƣ�{�m�k�q���g�YB��6j�NIPW-�4�(�yf�#M�J�c5yf6�����������������!�l���Sx�?����.�<��?�x��ޑ��­.4�74|Ula���H�W���C���-ܴl��&�A�X�콶L���L���}�=/��ό:Ҵ%	�e�Vy(,u�ڏY�8'&Ȇ5�KPSе�ƨ�P���Q��u�C9\�����U���ޞ�f�̾z"���U�g���04z�pY���X�T*Yq�c�6tzh�B�7�^@�J{c.� b�d|�l�l,�]�.\E�憎TT#Y����:����+���o�.��u
�}?A
�.�܏T���Pb0|@ی���	�z��ivY+
���II�����d�}�ę�/��b��
��1�c�����ul��xn�����$�����y�?
9Ya�g�D��X��Ev��.�G g1��ޛ|����q|K�����/�S�N��4,���sR�O�;����1eP�.?.��eZSd�Y	��	2&X+%���^�#�d�����.��cS=$�a~H�f��������Q�J��nU�����b<��5��Q~�}X��~N���3^N:�$P2��A�g�_�/��#�R�<��$
齃� ��-m�Sx��CT���Z<��Q���~fxJ����l�Pi�{DE`t*�w�w^�)t�⍔Q,��t���q�o�W����Av���(V�xTJ���#��nrK	_U���ykz`g�ۯj���sM�hK��:@IU����Da�-�IQh��:Ef���K_�u	<��~j𻉃r@��[Q�&ɃP�ҭ^�|�A��]�*E,��.�k��&�Hӭ