��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�;<�T������8�l��s�������{^o��;�cm�D������L2��h�$��I�`��'�a�gF�`�Dǘ��T-*]v����ִ?x������
R^%M�����%��r�~�G�/?EV:�(b�����L�`u� �=<��yy �Ny�OQ�U�&\�~���GI�d�:�n�J^�G�F��Z�ۧ��^*雇��N&��P^�@���y���.��w�feɷ���Y��䆔
P�j�Z��F<��I���;����1��頋��4��|�g(�!Ƞʥ���j�|��6�}�s����@Sk�ĩH 	�C1��[{U��]��u��D��XqwC���
@'�����zv_%T'^�:l>��,o�����g0��o�O�e�'rW�Ђ�t�̜
� U'���Y>��q��8�-c	RϠWC�!	6�k�4m��:��i��wo��=O��i��j���
b"�a*�5lX֭N'Ft?�̕e!ʳ1j�[D�ɫH:8A�\8	�(U�`L����]���)kD���[)h��U�����2���sӆf��G�:�R*�˚ b�T�z'��O�;��G���n�'���T¡W�8�?G��eц|b?�akб�#l�f*�ٯK��~$`zR5��h�R%:�B��|�6tGΘ��"�&lUj�<B�qF7WG��s#F���ѝ��7Y5QF�I��a։���m$���C�c���ϲ��ꩽ*����{JD�G������צ]AA�y�KdvV p�M"D�BU?�x�P��y�����d����>*���B�q�oh
v|�1e�սv�T`�J�E��#�f���������ՠ������\�;����+~b��Z��Y��:�>~�_z��?p[B��ś}�_�ҡ�)�[�����*X��0S³8D�ww6��2�Z'����ē���B%}��r6��z%k&��jG�m��<�"��b㶰^�h�����+�U�.�����dm�z"q�'����p�̀|7�M�>�7p^ߕ��1v�;A�=E*zm���S�]��Ş;���Cl=�R�-�[8�sz|��n�|�纠#"[0�wdI+�8�ļ�ݣR��6���	�+"VAͥ�����le�-��!
p~��+>{�?����zHx��1Põn7x��p0��4��ܕ�[9��r�~ؙ�i��z=F���c���.+{LԺ�׏�N[�Q�{����a��rR����Y�NP8�X�dPmƴ*]g��4!L��"
|�!V��'�<��1�<�9����f���,�̕ZW�r�<�E=�����2�z"����X�.�[�J֏��3�yy�=���p����;
����K�ږ��مY�	1D�\�YI�7P�܍���C.r�"�I�E��1�H��-��*�}�%|�$�'�o	�ǯ�LA�X=E�9�ɪ�"�v#Y�o�՜5M�nũ��~g���H��X�r��`�O�y 0���^[�-�����G�"|^��I-�~�� �=>y�}߄W,��6���V*(���-j:P��uL.��^gI�x&�>��p����ϰ���&v&Գc�f�H�)c���%:u�Z��Uݸ~���+ZBa-m'��z(�Ͼ;
�:^���h������" Ja��ӕ<���<�P�K+���yI�M������a92���P��Gx�vZ ���P�F$T���|�5%�2���XY�gߴ ��ܧ��7D�b��nK��g���:���~�_K`:������p4ʣ�+��:+��T�p����a�@'�DENi���S��Se5���xpA��V�'�� q�7�VE�J.����H6��ʍ1Yx=�o\�fhv��� E�"ܤ�/^�����ځ�$WOO���>�I��>�(��r���u��%�%Qf�O���I��<�fˠZ������P����[o��m��{b��/�����/_[EGӸ�13JX�b���LW(�5���-�qi�re�h=̰S���\�C�����W�44�q�a�6wl�YCpR��0���7�H@���9X"�?X(`y�A�X�-~�^C<3&��~�1��v��WE`Q����u�z��}��~�O�Pe�p�QXa�j�w�hO	�N��������t�&��H(�7 .،��j�4�#E5f������ȮQ�y��\Q���������#�!����}��ؑ��ZaS:�2\3m�"�����{�.�^"l��YV4Ls�jz�o/""4�Gt�e7e��s�Ѐ���Ц,fK�D�ڜ��H�DȼGg�^w�엱=�#{ �HJ ��JO��N��� DS�7}6�H�5,!Ɓ���$v���������?������f:5lcW���6A\��"����~���w�BZ	��;�G�NnP{9���aR{GF�xQ�m�"a�N�=��2���F
�A9a��s���XřAе7�\OՇ�X;� �>���7��vg@h�2�⯏�\4�|�q�pɞ"�b\���^R�X/��@��*�µE��zqF�&�I��~z��2�c�i>�C\�Z؇�*'�%�(�YE6�X 7ŪHY�0��3M�v�	:�����a26/��l�DD/���/���v\�v��̿$��R���bo��7b�1X����X!{v�!��*��G����D�[d�x�B5���%��_�TP�B�I4Ϝ�������T@�!՘i}@pO��w�y�4%B�e2M�z�X�q']��F�+��6���(��^��a��r��~bu:�p�wq�J>3��� �'1�J�E�}^�)�����TDi�P7�K�^SM������}��p~P��f������!� ������R�ȃΟn�>�]s��G`��_d��!:^&���GMy���]��U��.���&=��Gr�e�fV��n�\��Y2�1Kk�����F�[����a��x����]�m:n��k+��&�?3�����'ݷ�_���5�9g�d1�ڼU'}�23�#�e��X�]N|	����v�j�=��%�C����S r�v`�q�./	�c�t��J�6���� JE����j���!�oC��J�թ|鎒�_�s�_�	�>�hQ=�GG�p5*\5�/�&��f\5�cj��ic>�0���
���@����q��{����������~��ι���R� 8�LQ��לa�EӃR��4���Ry�p 7Y��AR������l� �gᐌp��"I����Or�OT
��ī�0Do�62��8;�%�7F_P�~�/5Zײ��ԟpջEV��S�.�^{�_�4���L��������ƾ���9e�x�Yx����M��̐�
�k�gZ�Yi+�=�WN&�"��6FVr6oY"�vxq��
�S;�꠾eW�r�[�R!�?5/XF�?��i,�� sK������踦�*8J:<:��r�yd��5t@�� >/:��o5���}~0��4!��NO�{\>�H�,�O��I����g�T�)��Ж�` �C��{.�@n��17�z'������P��m��W��T"}��Fķ���e%����׍��K��a�|^t��v|���7�[����\L��^�x4O�S�u�Wf-�-�]�=p1�GV���@5y&FQ�\�x%��u�H�8�:�.�.������e����R��X���W�b����ݒ��"��x)3����{Þe����Ē�\e�d?��*�������i.i~�[Q�x�}���q����ى��~���e:���|�S�NQAB��8΂Y?夤���i4:���:g+�M=�Q*�\�Kɯֹ\XOYpVx0�fY2tqu�j�P�ݖ|��N���2u�B�<�2O\�ii�4��Ge�SŚ!��ȼ�IoۚhO�Pnum���M���"Ծ����c��Qg=,�֞-T�ѹ����kC��@*���Q�}a0�a�%󑀕B��^D�vܨ���`�G/�d�ݖ�	��(�·r����%j9q6��zc�'/����0/�)�BO��!�hV�w�[K�rǗ�^2JZ-)95�����:��6�w޼�(kY������N�ɒ�׵����U�1��F-�{��7�wͥ-���);[�c�I�a�Ι�im6� h�60_#7{�G ���-ň.6�'g*V�4C�]����L��w`3����<��2Ѣ�3D
;?�8~s�e��A���k=�$YSR�v���E�x��|,#��A.%�F��)�D+בyۨ5����AP!\|E�e�h
��,xabV��`=�*�԰2?E�ñ�XT�����2jP=)� �R�����v��xЅ�A��/�:t�h�S��|�fq1�I�G�E�F�O1���;��m��o�O�FX�'N�?W����]�B)��0��8�5�cP��X����2�V!��=�=oƂR5��/���^'?e�4�G�ɫ�?������@����N7��\�$@Ǿ?�nQ�Į�nZ�Z��r�-�i=�:K��������*;D��#��n&�/�<��Ζ$�`�u�ĎAM�:BC��h�����!2��o�����E���|�
�~(1Rn�_6��6�.#����
/�����0>��W �q1$��T��}�Y�>�	?n�6gQ�sG�-Tn_r� ��e5A*տ�M����;������n���2��R�[�Yo�b���M`�%61�H�/a�\����E'����A��!S5��ȑT��<��Mvg�8������Ez���R���B��� *�p�WYg����ԇM"�z��y�lK�o,$��еN�o�>;�䬆�Vx������a�����^q�_ۏT$��9��W�!�����5&�صfH�`���@���=��?Uu~!�(F�|U�B%,*L�v��C}�,��|C$�طC"8����D1�]1�2���|��U�g��x���om$��K�
×aB�M������0���b���+iQ7漊�����+la�qq�0p7\�ӗ��"��)��k{��/�� l��Wpؘ�3�V�p�F>�|��EE�����!-w�6{}_�6J�JF�=_�x�N���&�z6���	�o������q�,[��,���z��Q^���	�&�Qc^�D���mq�h�n���P�$����Bp�L|