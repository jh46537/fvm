��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C��_�+��+��^���vZ�r�Ln�ҤpVCQ>˧6�C���_���Sa��#�Y�ϝ[f*�1�G�&ʤ�\��v��%�w�)@=�Z�:��4�9�U ?�� �DW� �	0��W�Vc���/��xlN�(':*�1����6g�}S Q=� &��˅.̗;%D	��Wddf8��.�l����r$q��^t����р���*Νn5;��KN�c(�,�~��z�It*8T�WX��������O��W�^��>��!
ȟ���&Jz��Q[�8�E��!�t,����ꪨh��G;L$�L�@�ȡ@�b�+�y%�v`Y�`��c/)M\%���n{��K�-�� H���O���g✄�Q�,�#��j�.�����k��׀��[�����غcj��� �2��F�`�mGf�Z��Ν:������ze���h�;����뻟;����d��<(p�op�6�&����K��_���K������UZ��l���v�Qq�f_w�"��/N���Y�uL@4O��v�A��a�:)"4��CS�la�0E,$���J8	��>,�qo����u���}��n?�L�콝-�:�5�>�����f��{~�/���HIF��oq`����8��2�;by㘖\�Y�}ے��3ж?����q�t��]	���уs�UW�VU�� ��ɷ�d۝��Ap���4!�8����m�Kv�n��B���8I6����S�$����|� �a9)�~��{ �?E���t`�T��d�x��3��	�D����� �=S�c�A�5g�ΗG�.(Cn�S��kBD_������cE?(��c�O2��{������
��;��"�@+�'ߗ�_8?�� �n$[=��.ȏ!���dhz*w�+���{��y�G�I@�XPkp�҃ݛ��u�B���VE%��k�G��T&t���OdO�vtC��5)�_CP�C�@T4a/�֙����l�y㯅�Z,�ݿɣq�I^eU��`t��C|-���2M���=�m��(���]��+����$���D�p2�Z�����e<�o��Q}���pƆ%�^��F ��h��������m-X?�E�t�+l�u�Ji5_W=	Կ	�My�w�P��k�"���t8|�1UL��Z
��U*,V����8��ޠ����5�E��Oe2�)��5�%�I��R����0��~/�Q�?H�RuIe�PB���I-�Rq��cM��v����
8x񠛖����r�4��56�al<'�d�Wm�A��c��@�^���?O2Nb�A*v�[7�~�%�HEW��|#�JCԏ��j�~V#��R�һAB����-��{���\aQ��!��8�g��݊kȥ�s��Aۧ~�el���O��]�!~*hju����T>̬v���v�[���g�楾��z�,N6�&�5��E����o��nE�;׺+��P�y
�����a��'�RHKN#�G}�ϛ$T���j�ߚ�{�6���X�m�H�Oƍό�%@L],��V �)��:_��A�ꡓIg��tG�hȑĢ�sm���9&O?�}Ω��+\�wG��o���I:��R˕�- #q yME�s:��$�J���vs>˔�P�v5�֭�J�����T�ެݝ�!j!,�"�?3�I�Pjp�E�� 罯tu�4