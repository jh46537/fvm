��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{�I1�+��:�M�cg�D���-6�8�oC�Kߚ)=P"�O���#t�M���S�k�5��֎����HA	��v4:R.W�9c��1�_}J�r��zM�X!̰%`�{6�pRH�]4��.���`T%P"�:���?�_�,�peB(�b:��̢���8W�����6�GzM������Vnޛ��ĭ�O�P�T]��[�24G$:߅H��v����H��S���0��e�&��P62ī��W	�a�=Y"Q��A��l`���O���8ԋ�	�V�@\č����E1�b�Ϸ����ͅ��W�K˗)�5�L�XL��`-��m�m�ۯΕaa�+7����:��>U+pj��+p'h�w��O}cG��*w5Xy|�o+�H�Jh�C$(�Pb�2�O�͎��ù�4�W�Bv.������'+�g ½	{���j����ي����W����us�̝��5Z):���H�C�.�8����^2Z��R�B���ޔ�_Hfd�e �z�Nq�����`�8�m�Ղ?�����3��v3>C6)!��l��,b���\2���K.����l�ר�-��K�-6r�i�`-Z9?�"��i��!�Wv��E&�?��A�x�����}�AeJt���$F�]H!&���m��	cy:Q$�!�K�S�bEq�3!"3�h(������[p��#��|A���|�+�X�df�K.����2�Q:��:p����#q�f���g��/V)�>�[d[.�T��"�돋�_�-��I��+C����*��V�pn4��/o�W���E1mr�Q<���(#cY!���vW�3����.D 
�%�c������;�!��ݹH�����U��PU������پf��| ��Q�+u�m�O#��ąLi�nh��)Z���y�>�%ػ�5Ϣ�s%.�5��lQ����G�-�P�\�����bܸߐg�tݞ�ɢIw1�D�1��JjW�����F̻��n���Y�.F� �7�z�r��M����#`^ G%|�FR^�c�v-�C	Q�h����z6�p�ݛ�tȂ �~��g-��^�3CtKݎ��H+s�4��!�(�G>��7���G3d���	�\�iS�Ri���"V!�V�����쮮PP�E
�a*lS���mO�����j��6�0������R�YN���W�#8�nq���t^ʭ:��Pi,�z։�áN���c�2u�.��^�ʠ=b�x��5RB
(|��S��P~uވKRR�+.����z��^���p�3�.�؂��a�$��]��\'���o&��g�l>�~�Tw&�ڜ�Tf��E�lp�32Q�<ԝ�+��Ŝ9}�։L�Њ��ӧ<����.ձ����\΍E�")��Itc#�=?�&��?)ۙ�|!��gnsE������;���ܪ�͟�|�
F״��
��a�������0\CU= ������R�^R$��&������G��aI|�ۈ�b=j|]��("x�7�6bP�W���W����_�� 0�PH����E.�u.�N&�[��=sv�Hi<��é�y���y�_9��`O���8"B��4�#c��D���{}�D]�+����r�������A��˥��L���kt9�����l��0; �^zu���c�hJgE�13[� hş�N�� �l� w�Ϣ6'	�X�e4����;E%t�QEK����R�E��7ma����&���S���$�M�{͇��ս4z�X���zצz���	��>���X���'\�~S��MO}X\�w��	HO݁ʂz���4��V��`�;��85���n�&N<\�i��v��S<	���?�SA2�&K�`�K74�����{���q�i����2�d���g>��s2���І݂qҩ�༤�-�~x0���V4��V`Hm�>�v�t*S��4�m��g/��.��Q^�W�����b0�*�#,�I�2� �2�X�tٓ�����hrJ�{sj�R�PL�Fۨ%2t�J�D����Yo�|pN7un�9�����buwd����yi_Uh�3 OJ�/S�K�[�VY/�nz�ׯ�У����~j�'_�P��G���qӗ���>h��P���C��X?pe-������r{",$�� ���	e�%����}��m�:a�mV:l���e']t���io�q����ڬͼnF�"�0�A:=$�Z�C�Z ��5�U0?ԏu��̞���}x �ט{li�������tQ־�Hը��Fg�%G�샍���Y��&��쫕��!�T�[�b�DmW��:\�
O��fqD5�G�)t�;����Q>+&#m#A�T�9>]Q��Q��l3��Vs��x��M/@ܴs��Ɯ���&��iI����Ԋd:F��&А��L�7�|�)���R�&���Gd¨���9G�H�����Y8� ��GU6�#"*������!�V��,�'�YSN����� ߫��B�e�|�}vZ|�u����<�a�=�zB@*�/v��'���� 3}�rV�}�ʙ��E^f����UA0HwH�B섣����:��ՙ��zL�а�8 Ԁa�ɂ.�B_�`��E�e�`����cZeMH����TF͆OQ�GF���KA�:�5��E��w{f�IR`i��d�z|��ogW�!�����j�1��`�%q�D /iy[��:@�7	��1	���mT'_4<��"��%!��3�͊��j��s\'�`��{8#�N��M�i߿���D��`��>r��A�3O05��H"��*=U�p�	�p�φ5
�H���8����1�kZяz��iq�!KD���{���XGY����2�i���X�� ڟ#$x�|�E-����#9lyN��2Pĩ�����ܼpV�>n	t�oԧ���#�}��KuP��|���_~rW _��2]4-��C� a�!DI{Ws�� x�̍A�B�h44�}(��$�N�z�G�#����8v�C<��jR��ͤ��I�@-F�\g�4(+8���#)OS���D��1qRQ��ȵ�d��ŪC��BV�E�+�Y1H�K��� �]����M�v�[SO�jGq��� ն�5n�}��Ҥ���P�s�ͯ�ܶ?l��{�ܦ�d�E��'Ja�'���}�G|�`��1O�����X��h��ٞ🨄�ҽ��թ"�od��}�hlI� !��^X/�|�S��Q<L])��z�4��
Z����9���3��*�ܓЀ��h���<��y��Ks��G���j��hP�)�k��_���y�� E��t}�.q�K�3c\2g�C� ���&;Pjf��a�w��Yz���З��[��{��l�1 !���g;hP(�JDʊ{��u����T�T_�͎���g%n�@rJ�x���v�S0C�B3����ҍ(i�_�0������p��]ٮ/�{�a��2EjQ$�ө�R��-��=@{@� �����$1÷9 (�����:$ҔA�Ŗ#������q�< �m>@�-$�3�1��wL�x��d���.�ӣ �4�ӯ������Z.WEx�yb���& R��D�Ӹ5�r���`�?F�޴�a���r)�ct=R���BE-�.�D����q��@C4�-T6�2�x�މ{�M��rA��+݃ ?֑"`6"������%
z�(���gTx�tU�(f��t4I߸�Њ���n���{j����]�Vl���7�YSzwGㄑ�M�xbYQ���;�n�.7R(>�F7�pg����p��@� D=�"�&�@����#(3��=x�)zQ)J����C-���X~��@J��38�䤤C:��}~��f�d�ʾ�?��(�X �	��1�e��`��l�AC@dFT�<*I4$NEE>��2�IAB/W��ky�0�wt���E�-�u�zoHD�Q�̀�����q��d�E�b�T����hIf�����/B�Y�o(�z	�`}&\CC�s5��6�M<ca�beOٸBڈZ�aֆ��8�Q���f�i���얛��Qtw5b(o��{�I &��2���}����W�3G�Aqk'���7L��bl�,�жW'h�=z�&�l�J����O$�B�,���mTx'��}	^�$73��^���8u�B����1�	�h8�َgF|��H�o�/:`�RH��?�t��o�޴�]p���u��<ͺ�0�l���)�W�;����{�Ƭ"��W �v0���T��D��g�MJ�u�4
�h�4Wϟk��k�7���xPf,���4$���v"�/͗:Mk�����a'~Ŝ�_	�]>��cm�Fz��w�7?��[�+7�-̗��M�O��ux�y��ޝ�G��o��_�/f�V=��w4my�47�B��m�3�sS�ҍu��
֛I"_I���@,�ک�����v�w��L@�বҝ\-��t^2`�����H��k�dm��ј���S�C>����Pb�\`� .D�`�]|��"���Y�F)oyK��F�� ti2�L���9�,�.0L� (SX��������r'���)AYn�6��J���x#o_��Q��d���2�|h�<]\m������oc����H��ɮ��o"&����o#>���-+kMC!��ܺÉ�Jƣ�-ȫ��UR���Zm^�w
���d7���0M���/	����H�79Й��v(,�+������7b����H�,�b�G�f)s4,���O]�-�ie��1��"^�n��{�!�
(���6�I��N'��u�?�D�f=����ZTqF�a��Xu9�iI���;I?�(��Ⱦ��J�l'C�Zt�?��+��&=< \z�|�����]<�/J�/s���� U��`�d���/W�d���Ǫ�kI�(lr�#�Qy� � �	W�N�F�KZ��e��V� ���1�b�U���}�C5�[�A?=ͭԙj%��X��%:R�#�ϯ���Octs�y�-��$X6p���o@ U����Ba���x��Y�{�� �zߓ/�175�}8�=������X�䲠:0j^���i9'�w��q��r3r����3�Ά4
r6dc��+8���qü�d
�Ga���{�u"
��:�����]��M_�
���D�e��	1��t�L�#`�dQ0R 0]$v�d�b�f|>-�7���mGwE�h+(�q��J[,ݨ����ߩS�OסQ��=*C*h�p�=hi�d����iQ��A���,iW�Yvrf�+�2�� �" ���n�Z�៷5�SC��1���:��Kg�It1LR�r�1M��9���K��>k�(��_Gd^��n>,t���1����i��l�$'���h���&)���?�8�oA�^�$M�{��>7g�d]�)/�i���Ji�55*�'Q<��T���]U�md+ڼC����-�ߚ6��K-}�)��"�5y��@�v�&���$��V3ą�w_u��4u#�HR�u���R�C�dJu�bl#�-�5��;����,+�[�XY���qcf�AƲ��Zi"��2޵��3I�=��ӡ���������j�6� ��L��V���~\�6i컺v��xͻ��z'���y9b��x�C�3�aE
������x� ���*�l����Li��Ɲr�G�<�͔A.��u��p΅� �]����"�wJ��7y;^�9�+�ͭ]L�Qy�O��}j4s�| 6/WA��:���(�W��c̐e"�r%� ������Q��W�ɣ�bBX}�3I���	ڻ%? �~�c*z���z)C���J���ǩ҅/{# �n֋}<+� �ڕye��3*��G~Q�T"��9����:� ������,~��l�I~�~{U�F�ek��b�`�A,LC��q�^j�xf�n��6�Y6'J���N��,���+�F�M�`��cKm��?\'0P��D��Mv��$q`��(���G\�F��=cW �\UZ�d�؉�plQ����dyW)b�=��]ۼ�kl�5�:���m��ßWj���7���k�%�Ο[/��7_��F�N�I��'��!�΅�ԭ(��c�W�x`��p���}5W�Z"^��kԘbA�:@�*_Җo=F����"@��⧉}�����Jzw�b]�sO�٠h�_���q�(��y����a�?�I���*?C6M�4�x2=O�M0m�a���b���:�n%OW&�
~wfe�b�q������%R�M�}�~kݥ9���2�xӌ�󣦒��T��=P�I5ޠ]�q�9	�p�+�2D�g�٦ b��C���Bz�>�,�/r��sc�f �yj�CI��ޑ���z���N��G-֝T��@n�����+��w�(���hzM?-4��}���'#j#���j��X|/1u��]�e����9�V  Ke,
4���fC&���8u�\6�Ƿ�I��*�|��z�Y�?�yL9�W��B:�~�Py�`!�j)59Qn.�PʑןI��m���I�}bt\ s���ŵ�8����6h���aUUc!h���$�J����Kv�3����!,�ۃ.x��{]��x�q�s�;���i��3k�w�=~�Y;�0�w���6U Ԅ��1�T:��^$g)��7���ǁF�f�����}yL#�X�U�^8��}�� ��"�=�,�_��Q_��y��:�C�]buVj��yf�zI�嶕�,H{A�y/|d��eA� $(�AĜ/B��)pJ�u׮��Ϙ��C���~�~����鴌%M�>F�������Ho���t�sÊ!�h��N&��`�$X�[��^��0/
�<-ud��w�	��vSb�oȳ-��׏�o������ugW3��P���I�������O��.u��xG8δ���;�H����!����UGz��?���}�GFر�E�u�k]�ػ55�<�+?�7�_H`Ҋ�yqLz<�]�z��C[H�8>���q�ȕ��I3euȆ�vi)IX���"�^_�l���k��5�e�\�V�Ȭ7�62@�-yiïo�l �s��
�"��9�A��n��
*�E�ء#�J��E�A��������h�'w��{���z��ߴ��)�@�|�'	�=�"	"�#�襘{���c퉔5Y�f�8��	�~��O�����;���4��{C��� �[�?�8}����j���,�<�)^ Z��H�}`5|��V�}���9H���w�#��%3��
�h��s�ސ�����D�;�RH�4.������xaM���;:�~��-�o�����@k�D�`�_Y�c^���赜�>�|�>�e��E��Ⱥ9���H	1$��>�L�w�̇Y뚎��'�P"-�:/}�w�ld"&�#,B>���`�)J�O9���3h��VQojM|o@��#T�u����
��n�ޖ+
t'!]�^����(����F�rMn�s���B�����K�#m�q�H�`q�ͨ]��#U>��e�̰�i�R�.0Ѐ����^l�I]�h�=0�o�qD�x2cv��.Tk��}X'�G�؊؄©���|}#�e����8��[��W��j=��Jآ6��#��b@�Q^�g�����H�&��}�R'���t��a31�=(Q�'�lK���P/�<��"�rÏ���~��!�����4J�>νH�9d�g79����%G`��4�"��d��RS�n���s����7��"�5��Ylr���^˶����Dlq�6�lj���'?���\�<�c<i��t�W��h20�U���`z:D���ȄG%�Ү.��M�C��blX��4� '�-�(�2�&khb���ucZ�ڿ���pW�a���*"�>�l�y�/z\�j%m�$`S�������Xv��N��X ��-�]D�/2�LF0�>���c^�#@��
���X����
jsK��=�=<�or�za�H� �/�	��*��}��Nj�rS��ޓ3�[Tc�A[Lw�j�e:�:�t�J/�iy�7����%L�����f�K�-�����%�L(H�.>"�9��2i	ƨI��?�e��R,�~�rM�lR�F��o���5�
̭I�b�V�3�+�NČ5X��&�xN�i�=4�j��6!$W��!c� Y�1'
PK��[InR�!�󚑊�a(H��o��d�Zˑb'>"4��������j%�ԇ��CK�O�:��Y��$�d���=�V��]2�kn7����4�Q>gq
B��=.���d���i��]�.��~�S|q%P0_Q�߼Bs����H�hv��w�����^0�e�r	��!B	����U�ŕ<&L�
�d��@�6���L�P�`g�CW������~���]:��B��۬f
>�����䆆�����H�h�c���)E����d�)�1$�I�υ��e�sEҞ!�u�=���z��V�7m�h?z�A!W�fF�{ �M\�#���.�J�ͰFF$0v���,ђ׀̃`�u��0��j8!}x���i�!wͽ>p{לd	!ߙ�/0�z�A� ���?n��p����w��)��6�\��9�t��9�Fp*���|�A?9���hWN	�uՈ�cp�C��m�`�����|a-�V�����丠{5K�S�Y�ߎ�]�E��HS4��T��z��P�ҋh��&�we�MSi���'� ���l�`�E��,�5��	o���̮�st�:Y�u��FYvd�S��4��2���Y��i&���]�@А��m4�dG���R���-��:�(u(J��ɫ�5l�g�H1%�/�`q�r����9��ll�%�ZG��jR ��Xס�Ev�& �O�TZy����n}�L�c�l���I���E5�09�BHǝ��`ws���>�$�� ��A�v�τ�:���� C�ʅq'�w�Bk�FH����^\H<m3�/�u��o.��aԴ�a�צt��	�W�d�+Q@�BI��T pM�]f@+����!6���m�A��(D3������":N2�g���۸"L�Z1F/�~sG����(!��)����!�wc`\�h�F��E�%g�Mj��,G�4�:�+P�K���;�oܮw���p�+�h�7;�ڐ�lX�V�ے��&���ˤ��y+)�YG
l�r��'�ԃ����`�5g~�#TL`��_�ɧZ�Q\�g|�(�1��f��G�"P��$�ʠ�-UvX�$�$6g��ZF���.��Ö�r{-���>��9�Z�&���	;^A~Y����Y�򑉱8[�E.��q�� �Dh.
	��v�"i�V.��Hg����݁Z8p,�~.GM�W�riQ�?��~�v�Z�xn��]��
A�� �΀b.ej71�rGҜ^ˣ�H�B��,��*��!>#�N?*�����7�Iy��x�T0ֆ�|�b�tyI�H"��^"g�� �F��Ra6�0�]��9��$d>��"������x�����T��7AU��`��t�ƍ�s���ٓnɕ�c�����M
`|"V">��^)���&�-�i0FH��$?�7��w��!Y@ɓb<��Q������G��y��8��͛xʔ{�HwtޯX�E� s- 0��A��|g��!�~�E�d��eQ5[�Y�T��e�(z�1lRpH�TE�»D'@�������)��c�ZF�\�dYZQ�3t]=%Z�n���^d�y��
��a�Q��	�	��)����t֦T��%��GW,��uF�zzG�;
�q���j��'����f���(t��c���(����f����eh�=Qg �~�:�5��/Pf����LTފ�r���..v�a�i��O�"H��^�{<� n�'�ķ`����ļ��_�����!:3z��e��qYG�hBH���Iy�7�	KOk��W�t�;ZZ"bL��:�tJ'>NX
a�'����K�z3�ΗrR���`��&�&^� �.����$P��'N_�[Uֽ_�S�@k���c���v��-k����ݶn�K�\�-U+�ir�����OM<�+�g<�j�G�z�6S�QT�\,(�tfOb&�$sr'�f*�޳x�M+�aX�V�� ��6}Dȳ7v�U�7L�h��d��(�-9�p�;�� ��w~ی����LH��>뮤򏼆�9�we � JL�2Z�!���(��	��i���	"�N�}�G S��}|t�_$[��Y�8�'}�-�o�x��U��%�����t�H�-�k��6�;�b�%� ���[=�L�QK��Æ2®��+)��KM��.�0��C�#Ɯ凉#3O�|��)J�̈́=&gtCuc�#���z��/v������Q��pP����B�%_�s�[8�(�*�W�4�&��A���� $�@��]O���i<�