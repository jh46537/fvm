��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��J��Ǯy{{͂�[��N��������]m�ˈ=g$k�n^v�{.��ʠ,�{������ld|N�u��v$�R�i�f�,Y���v��w@H�o�v�w[OC���UQI���&����RF�-�5_spU8��Ʊ���������k+�(��P�{e݅3�S��0��醆�a�p��ڧ{3�n	��?m*��uuTB���1����r-sG"ة��oE�P�pO����N��;woїc�	����aћ����#��,��O�����Vg��= v�ﴌo�ǭ/���9N�[��Xsr���%(Xy� C:>��o��*�c1x�͠�҈����������x1:���C��ɂ�a��ܱ�\���I���M����A �eNY#|d���������e�j'��k�X{�h�Eʐ��Fmg���b��p߲t5Y-輮�>�����c\Ӓ��=g�vhò�>�U��O4"�ӹ��O�*�P��*��l��h`��iF�
�W?X���]���Z4R�@C=.7P�]�6�]�U�jo�	1��D�-��J��J*��vӊ\��NR[>/q�u���)a��pa(�3�u���OF�J=)N���O�S��Ȓ&��U!q�_�p�pA �L��^���'��O��7� ����I&5~��:����|����U�.��,��>(��\���1g:���ܘ�E��@���{P;Z<�k���ȩ�dM��l���.���Ũ�������-�B'\Y{���� 1����T�$k�گ�DW�q�f�z�y��V˗�3������j��������23v���1��1y�Z�_Y�\"�U澹<�	nzEJ]�6��L)�|8�GI��W��,f�lqx��x��<��X̠�U�Ym���Z5�f8R.FϳC��Y�����~ɦ�|;˗u*p�<�R�����i�]$ar�ĮI�m_�K��᥽'$�������{�t|�a��<�~����g�l��y�&R,��BR��.��$��)U��TU�(�W/$V`�*r�n�!�44A$���
�-��3�U�GL�����z��7:�������A�,�q��Q:NiV�p�d4� ���ޓaLBg�k�e�����fD��x��a|B��i���3x����6)_y	�#��ˈ����������
�Q���n���YUv'�U�����~��Z�_�^5"1J3b �v��
0~퇷�b%I�m5
Dh�`Q���Ӳ����)/���Z��5��pf��%e�vŸ��Y	RA����rS���L���'��Hx�J�0�M�G��c�����<�i#���>�Ʃ��G��<�l�_ vkϕ%�W��t=�=��>cv��4T�_����󐌙Bx�k��y^��h=��>��h�r�}����gICpM�Dg�m]J�8>�x��!j�nk\v�~46+(UTlY	Y���U��V��p_�����;/�Xd���t
��Т��䬹�v������NҊ�7,����m��d���7i����b�5b:=u�Y�r܂c��#ssZ�o���Z҃,��/=~��v��gG�\�y&��m�}�LL�ȱ��H_Î*}!���Q���RPQ!$�}^�B��fӡl��#P��.�h`�>T�߳���i�9���l�q,�����0iIS��Ci�� {�c����*]�|�H\���^�~�W��6��4��B�.�.d���JҕVy�鿫Q��+ҼÖ���%������M�a�m*���h�[ �l��,��+�8e���\3	!6/em�|Q���|�A��?����vY>���B#�	|�Gc��ʶ�Y�}@� 7W�۷�+1X��[�� �Y��9��E�5�>áEy����$�J��M�h����s�"��aFw���W��>�i��H5-(�)C��d�gv�΃��<�9̶xI��/��5�mR9)�=�k?���5
�!^�ׅ�,��,	^�-��Q.EyI��r��&/���0�cA��lt�UZFXA�aUM��H������$�_,�%�j�T ��Lp��,R#�4�F���2��щP*���;�5��N)o��N�S���� ι���j��+��Ml�튽��<�$�!�,�V����+�T:p�5Kv�+W6�iXʆ6P��N�A��Q�����;��$]���ʰK�g��P关���`�
�Ζ*�����Nq` ���j������.L� �{FV�魌]D��Ȃ�!�ʍ��p�t�c�F�5s�5%�qh��s����.��\�% ���nE����
�n1/�<rG��D�c�5��xP�ᗱ�"���|��l�}�~q56	�u�:�g��Ģ��2��8F������|�Z��Dˇ�a�j�I�6��ۻhw�Fr4��옿vM�N����U����*CuQ~���9UI�s,wgrxp���^�ٻt��֯9E���~1�! �7|W��9R|���M_�ϒb8��ԢL��8����K#}-ɂ�kh:���꫖j�-��#����ϫS]'s�%��!�> ҪB���)U1�����E\�"�9q�E�K䔢/:;�H��#�&���e�Q/�Q�Ur�<�.��v7��T��HV�;J?�H*-e|؇%�G�6�闞1���6�l�'�٫���1��"B���'����G�Ofヷ��J�v7t;F_�~B�H*B���k�l����@�[d��r�=�&���B����Q�D:����
M�c��7�.��]�5�lC�K�`��[I���5�B�-�=�2�1l�Q��4��'�U0j��$W��rgJ�QU�)z��m.�ԯ�I6e6?Ճ4�`1���6����p�h�A��S9o���[�lǙ�.h�F��N�E�x$���2�12YEo�=/�DD�9�I٪燎q��n3�1����	7kU��8E�E\;;˓�����տ	`�Ag��!:g�t
�U2X���ْ�lW��g~�r��D�t7qj筏���N�R~]eW{����A㗨Kqx	ǆ�����/�GR�:��q��rd!HC��2�u
|;�1/����� �
.r*�@����>znn] �fc3��Q>���5��?���3%ټsC�N�����ѧ��0�2;
��M�N�,`�L��E��qa.ݹ��)�i�c����n5p�g2�#3�%���k��e�t���Eh�	�@��J�X,�d�jY�<�Z�?ns_3�f�ד[F.��B�^Ƙ���lԔ�)�aj�0کJ|V}�>�/�9Ӗ��[@=��F$7��u�K�|qCq ��?']@Y8^0I���9A�c�� �R��Z��~���iw����<�yj���:ݪ|�On����o�m�zL���y�a�� �����G��q�S��
vH}�F����I�Mv.�#��)����6
�D�h�Zr� �N�W���6h(�&���,knn���Ĕ@�-Ū�dVd}�t��LRѧ��w�)������[5�t*"3OωCY�NR	�������*8D�8cg%v,�.5�k���OuJ�Dy�MH��j��f�&r��;.�!��Ц��f�K@㐁��"�Yv���%����Ǝ[ 	�?�NZ�]��4�%y)�?m��� �!�(3�9�X�d^�P���k���)ԋ�:�S����8��&�H�8hʣ@��'����ёB=�8�9�]�	��֩�Ě]��a^������mV&``��׏���!j�u�E��g4��g�]����b��f�t�n���8��/M��ꊏaZ��̻�J�����г&PNɢ��,��p��� ��C�`�7Z@��B]�1ж�f�ٍQ�=^�U�m5Kx�o��-�#���1$�Z���B�|�&������u�>yV�����3���O��UH��E<�ȷ��%t�Yv�����
p(�B��HT�C((}v.�|�.�z�
�w;`e�q�@�)�Zk�g�b�L��KΊ[����.��v�r�L��n������e�QQC� NgQ��;�6�[�,	�#�7zΝ�<`4�/�o�4C�4�f��3_��xHE�.
�=qBWw-�{����1�ѵI��܀S��c;F��C2x����S�Be����&l!�����]��C��Fm�����%u*2+Ũ�oT�PnJk�$�.}p�x� W�L�n�d������NEĿ���T�L��_^)p�Cy%��,�5?��aI?�����0M����aY�AI�\�	)\2�>��K�o��;jX�Op�Q�@9�G�%�~Jn$�0�@�ķ���@��1/��йZoD��n��F�H��.ș7Q(dY�[n�{�X���A�͓1�-����|���S���9�NB$��&���o�U;ﱆ���k�z��#U�N��,|G���h�1��T-pX�AN�:�e)��|7&��0�bnTd��7�b[�?�*�������҃�{q�̳�d�N���l��XE�o:�P
�%��j�k���p�zݬ��,�@�]�j�@֮�������]﨏���*�G=x�
���_¥Pь�v=!�#������v���*6�W������?<�~��Ƙ������/q��3�|��]ݘݨ\-f��|�B�j����Z��:����D��S����|���|��I��%��9�
�₎?aAVt�֌
cq4���8Y�����R�v��#� :�V�H�=P�Y)^J��ol3�����E�B[}v�`�@�7(�*�@��h:H��yGZ��}�n��q�S�1%��H�B�+*��R��:��M_@��d�����u�E��; �S�9Bߜ0��8�HY�|[��#����Jaȋ�hD�}H���!��X��NNQ�pR�D��0���`rZ�D����(`;�Q��Q�=�_��Q[�J����O����@�MMN��x�Vu5h��*\1j��{�m$�����SL�nK���A����sO`2��ø�~h���� �
�0�e��oΕ��������WpX���n��P/�<�$h�,<w+�i~��L�HP%G��Z�� g�zԯw�#�5����'�P��R��("�8)<q��3�n�)��;�x�FI�??yMk����g;��޶6z ���'_�X3��ق�7˛3�a�(4����ݡ����|����X�Y[��թ]��X�Ir��k]K�Y��]���	�@@�5�]@�X'ςV�&��P�Iz�"�}mi �$El�dG#1�7 �Q���!�//���C�^��<�����Gs9	Bۥ�`}���m ���T$��a�Y�eO����;\��6�4>Q������	xn��DM�9�G�����Å.���^�5��I��7�;�������O �v*���5B9��}�D���k�!��dߧ_�DQ_�p�K� O��#��=�5w@~�qD"�}<�N�E�Q���7� c~�`�
SnyG�t%-�hځ�����n���}��7�߀1�
�f���^Lm8�҈�p��^}� *M���-^\9�}	j4���� ����v�"�dvѥ���5���h��!/�&��C�0v����Ѩ�yN�w1�K�(�q��t��ɥ�G�n��So'B纏�Q�:F{W�f�Dư��=#0a�t$��G�j�Ε]	c[�C�=R�9q�ՙk�u����Z��n�YoRď�L��0�6z�E1�c8X��|}gc^����f*��7�h>�m/�B%Q}V��NN���H��E����6̲�%$�GX�p��~r��Jf�n���d4Q���qB ��M� ��ls�1�k��������m�eJA��X��"-BC8{�X��'�H���,����ٵp`y/b����������&R����Vڮb@%��Z�$���(z������㓤J>|�-����Z�&��K��G��=�U�`�2��r���c�K�\K�r�_�9FQ�~;�!W��eo�%��%�f`.��ɞR���˿s��:C�vZ��Xc���U��o��pY<�v�(ʠ��I�ՙ�B��]���.ʘ����=R=�$���M.n>��K|��!F4kF���E��𢼓18���o���^�<L�AӠ�y���j��u��a��#�K��_x�tس�C�k����oL Am^�J0��\T�S�"�'G�Y�~PS,|�Q�<w�
����n���O��6��c;s�@�7��6�<�r�����E��D��Z|�yz��p�n=Y�4����(#����n�h|�?%;#8��u,�
#o �k]�Fh �^��8OZj��3�4���+h �9Zi+l���-�7�Z����U0�E�
�ё���|4��U9Qfȫ��"H�1FcĆp�ߐ[�V�W��ƜDfM��!�cq<�ک�:�#'��_q�����ێ�� ����И;����.�W��vE=ny��[w��� ���ֽg���]�]��~g	��2�CT�	���^f?.�2�ﲁ��L(�9�1�����|8����sw�^���l��	��įx�A��r']�>���+D���--=OhdbQ���kj��A;��B{��b����KQmqy�sl����QO�c�d���
<nu X������,�O�:���ݱ6Gf܆Щw�o %gr�D_CC���ށJ�A��Sllh2N�h��f�8$�\�a�&9�FN�93y^��/H����D��{��]2��`�@y4硽�/Լ�?�������Y�1�5������$���d �z�t��������V������dn��� �����,ݰ���W*3E>�*8)���!�s9���M��<}�/5���
:�_17�D�P!����4�hU���v���9��$99���jc� @��슆���"a�~R��M��P��b�oe�Z���`7*�mM�4o��bx�p�����?r&�CK :4��ő����5&�N�3m&�Z:y!��ӄz���<T���M<:�d;��2�H�������w�����:�!QvN^�K���N�D)@x��B�j�)�
��Cq�4XW�`:����@V"����૭9
h1 ��b��y��qE�7��R�".���O۟��^�2TQ;�X�c���*��-8�d��	���a�>�9g��N�
S
��k�3r� Q�2���'<^��<x�S[�����2��Zj�FZ�1�#(�g��S�NǠ�FcD@*�`"0o��/z% ;��l�9��y�b!y�6��!���R!��&Z�uf�Φ�CD<�,�ӌd��H4N� ߻�O���{~	}���{Z%�;���8�;c�ۗ�m������+Z��2�>A�I�f���4��O����0�@¦{[���u���p'��f���t��:�B�r^�<���>m1�[� ��hu�pD�:=B�ag���,��{f���J���y���!���9�q���o���	�����5���u��{z�g���Y�_)=0`�<��LF됊�|f�V5��̹�&��<����hz�R�΁au�툓��B��z�(�F�2`8�D�<Y�+��=�qO�\<���q��XO��j��\�	�u���*��҇�4;�9���V;��9=�l�[�g�����?�e�{;$�.��x,����!1�J����Ӹ6U���Ыe�pF�4`�Y[(��}�R�7(|�.:��j*�E�JH�Iu�����p�l�Jj��q�@��l|0����܃u�����UT��f%��DS��7i��-��#v@d�/Hu�|1#ۥ����3�ms���\X8��u�g��>�}2���a�)x����b�����䧺�2>���u���D�����(�N�I(�$�,��]�iiiq�Lq߀$6឴h>��4��8�ͽ��9�R�Χ���/��q�<�Cr�]��M'J����X�O0�<�ĮV��]]����k4��E_�	��_��*�H�s���{���μp�����
3�8GT�w(:������Y6��M���L/Z�̬�YW<E��]��1q�x��I������\�CP�����;7�t�KЧj����BTq?G�tKw�1�k�^ ����Y��-��C؋��h���o�?�']U�FkP�R�D�� ��������Z�l���סw�3F�ZF!�p.��d��Dn|�L�������m��M��S/6���T׀�)���#�E�f�f�}�c�{{1.�o9NL�];��}��4�{��mOǡE�0����{y�d'�AZ�������6�nH_4�}cM�����[�ݫUyt|sEP���
�iF5Ł��$t�g�	��}�;�����*`:3?���{*=X+b��K�rZ��EںJ��
wQj�H@�v���)
����������u��T�v��?g�e�i3�Ԋ.IY[�������LX��p5y�__Q�zB������*�OG�^�B�S�F;�"@�R�Iu2�`!��Y����_�V9���hZ�8�����9��K����=|��0�ϻʱ[�z���#�V�P�^�(�Q�p#[�|���R��!����C�:&ǎ�OJ�{��p�CH~d:��]�~ ]r�kb71�K�ɫmy��H�k�jذ�XX���6���q�4&�t��Z�����%p-<�3C���Y�15�k�$o8�ʰj�2��l��Ս��d�_ӤP�7��f|~,��R���A���_ԧ(C�:|zO~
��Y��r�@��OT�c���''f}�gy԰��j1U���o�`Z>��ذôԯ���	���q!�'D)=���8���~��q���wʽi���O�h 5�ri�����6�cN�}F�@�X�/���=��75F���	U\�Y���2z|��M���yϞ.�B���&Ͳ.>�v���KM\ z��)�aĞ�;Ν*��K����v�]�mR�c
�x������G�I��+�/v��5�� �z	 M,ȜB��ֈ%G�t�]bƑ�Sr�1G�7�3L�*�v`C�$��ND����C���+�iulr���)m�`�$=2)�����n,wp��������WQ*f�o�L�k
�+$<�Jr䪔����"��!`sAYk���z�^�Ӌ?�|Z�=�GOJ��4�^�=A%�h�#��"0I���A�	�S	Z�O1K�{Jn�>$%��q�V�-){��}9���V��&NTQ�D�w\��fn�w
�/�@n�,�4�uf��'����'8��hcsK�~�L>OyP~���	>�(���\���C��ﾴ�p��l�y5���~p֌�D����;�������D�n=s�W r�u���8k��l-����Ԓ@�!�l<A^m�g>�7�"B�o˔sv�{�Zvz���/a��R�:�3H�]�nW��g�{���9q�2L��8gT���P�A��U��̫�_�V�/��q ��RA��]_��n6XQ{��A8�k@�T�Py�u�|ڗ�KF�C8I�4y��E�<6(�a������qWX�ǭ%��D6�S�4�[��$rOū'ܑmϹ΍�ϡ8������Y��Sˮ�e7ū>{>K��Sʸ4cl�yZO��5�<�+P�kv��Ϡ+]�@�sq��Z�\K	�֎K'�3B1�?A@��9j��m�'5�yv��8��i�b�ky@
$ڗ��2�W"So'@����b͇�Y���m�j�����Ρq�V���V,�{�=�r	�PM�^����;�w�C`�W3��*b�Z)����xzn�ނ6C%��p����5�~��󐔗����%�"&��̍�c�c��S�����C!V�o�KU��Ʊ	ڏ�9H�!���X�0�L����G��g�k����_�tO�Q��4;��Pi-�P-��I��/����D�>^����ZtL� \��6"�+<�B�R��y����C(spP��ǳ�'D�@m�J�@it�!�q���^�{�yL�nYg��NݬZ*�Q�>������y��J�'��	�\f�GH�a�gZ��S�Fʸ1�e��|F�@-�)�����0��M/����YR��R�V��yi��V&��+f�Mw���tTJ"��b��8����h&-�|Jq��5.TG't��PY��Be!�`���8^�mM�)$�=�#H����ܺ#Ů[�Q��޼�VG�N�1ˀT~C�-��O���hѫ3+�C��Y����"�I%�xh�=c*iՅ
�4�B��~ҥ�ް�3�QL�<^-��7�ƶ:�U�"w���C��>H

˲��D�/�BN������؊���4(���D����x��۟�G�(���F�4-N�R���ݠ����a	dyL�NLٙvǄ��1"�V�;f�Ff��m/Q�˷Q��KxO��ro��Q�*|���rA�!�Q�%D��:�Ux@U���5�W�9��i&h�ǿĒm�V���&����Ȉ�C5c�3�!t> �G�������eۊw�n����r,`�JL�[ޱ���18�/o��]�y&��z�^L<K�c����Uq�'	w�9�7��FC��#���Y���q��{=p��c��Z�N/��È�7@E6�{BDk͟{&n	����V���t���t�Ixeڡh �g�Ҡ��҂�FZS�Kr����v�w�H��Y�zj1�����֋��~T�7G�j��@I��)j�t�З[��^:���)3��`��>Fzw�=�,�i�ŷ�F:�7}�#�NÆC�#����54�̓V�ވ+m�k��I=�A�.]��k�8�{#dA	�����W޸� �Uh�ĚR�&M�L5Յ>>)o��G-�qo��@&w����9��J.�f�iT�k��7(���dȜI,&����/�[�≟�pdcJz�1 T���G\�o�[�>M?�� �go�����w:��%3�AO��o �*pck��DџWY;���f={�Qc��'(+�V7�D�g�l���r�R�z��d����a��QF�� T$Q���,�c�ZTs8j�J�*��ҙH��:lF>^u��=����5����`�}���G4Wy�bQ�CA5���8��u3F��]��Q�K��)j�Y�#����Ų=���-��(���C�;hC��M��h��t0����n�Q$��H|/�ɵN��%�l�Icdc@4�u���^��ߚl��n���&#V�S�|ބi���jb�8 !��欎��v��7����a�2����kQ���-*M�����+�bD�n�;z)��#ֱaV�5������öw�HZ���ѐ��Q����T�L����Fҧ�D����Q�j��)�0�B�U���^<t�Ì�#���˹�:�u6x��焃uz1}#V��4�Ċ�~q��"�'DhE��r�'3�퀸�$�6�*�9E���Ey�u����?�˰��O�C�iE��멺��΍{u���RX�G2�,��g���G�Y�,���U�+jn|�u��oN��
yRL�"s�h ����P�sl$���x���Io4��͌���FFc��yR����I��^���x<�|��|��[\�<f��X�%�[ɬ@��'��3fz�]ôq@,=�p�1��L�?�1�m��'q���P�53��i�r4��;�o�T2�I�
��\M����W��Z�q�bT�=��yުM������6}�E�5�KH�;_ Y�j��~��ˌ���f���꧖���¯V����l�ܜ�l]�cX�[ֲUK���+w���0��E�O��~�!�~��>N����ة5�Ȝg�ԬP���>n����2���`��*�����K|�s�! ����_7"����<ܮS�v��6� �h�U�ht�5���2D���E_l��K��_�^�	i�Z-��
L
h�ɋZ�rr�7� �p&�|ʨ7K� �#��f��%�+�����z_6)�Rz����x�m<��8��R5q�kN�:?�{���km��)�� ҕ	=�
��$Ȱ�`ˉ�)��]����.I�������P�ҥ^���h����t!��K�"T�VއU'8�PB�L""D���k;�q��+r����1Q�ک���ɧ~(���D�O߾B �z!��Et-����֏���/\��c��p�FY��3F.�r/ޛPB���d6�aK�0D6�]١C	��3�_CPY(��ǰrh�+n6�7�ޝ�Z'���-������eA��hD�EP>~�6[��N*t=1���&�����[ ��y7D�Ų�G�L)\���S\��`�zP(-$1͗��Q�K:3�:S�i�ms�[3�,7�����ÄQ]Ġ�|
<�6]�_���468�،����.{I�|�X?$��ꓺ�e�Ge+xxU���I�\'�/e�y�R��J?#�X�����U��Ygo�׎ӅRk2����Ld��뛚�%�B+�a��@���S0��~.u�WHڴ}V�W��rJ�";F��ЊtB-���O� (�=E�B�7��b",gD6i.4��O���Ma&X�2��(h����ZUTl��L��D��'�dE<�*�5Z���6ߐ��734PP�˥�����9� }��(����0�M��j�w@��{'�B���ry�2����� hXt�"Z��sf};+�U��tܒ@]RR�%,�r�T\��~�r�!�C��0ۺ>���3}�a��}���$bA���K�__��������"��
�rRC%R�R�.����RЗY51ʦ����߬��+FB�|�n`�!�Eғ�h)�q�`�����M���L<G�ѷ)�PrZ�=��vm�E;�즴��HcD$<vk��Ŏ��@���y��9)����a�Eq�)7����b��m+R�����j1�}g��(I�ja��2I?��Ʊ}D~�sԻ`��"� ��Lr4`��O-)�Բ��GK�}c�sV���Yn)Z;B߀j"������#~��Ou8B����n��H�<�@�6JŦ���C6�˄�:`�vЄ�5~-\Iӿ7��-UH��
�r+V����R8�i���B�Jt�q�=sV���&vc�oc�#!咙���=r� u1�� �8��3��J��;�q�Y��a�ݦ;f�����hC����P��h�-��h�A*}�+s�/��N/@��g�d
�3��
����]��8.�[��ͦ����=%G�/�z�-�<�u��ݮ���h�U��U31 �14`a�ƈ��D�M��p߃L��K��p��T[v��4�N+��vC�9֓��՗+%G;���.��@���޻�E�6����?���=����*�}�ѫ�7�n�`�D��؀��0�� �����wu/6oʃ�m�5
�����%P0��S@O�C-"���MD�#�?��dx�Z�Au_��A�(�"h9/���`x�A[�w���2v'�����{�1��%$�qK�����ź�5O���P��*��.�i=xY<I�G�Б�4�|��NԚ~�%ÒT��-M�?��1���Mb{.{�Wp���6;ځ7���2,�e�\���7{�C_�˳���v<�At�E:DkPv�Gb�e*��s}?������;����lz3_HK�|^i�f��D�-�wR,��1�$Εʕ��J�X;IDH��Q��n���hv\o�sR��dW�h����L	u�#F�Ӧ^�VY��V�h�i���������b��<x�b@�<=�I�WS+J����(��j��¶n�/B�Tح6��T�_��\�Uk'd)���Xt�#�3d�&�*���3k�I.�vѝ�<�t��O;�6H�
�XPs���>4B6:�Wk	�f)@�v���B訰ܘ>�c_X�a��Ը�5�
�ʅ��,
�߬�|�2f�g�J���~RU;�xE.�d,�f	�8h5Bw�R�&���~@��w
�lV�i�y񸛁t�a�*BL�:�S�܏�d�]�o����.?���T���`äTW��?�S���
	�����E!�u�9v0���1�<F��9g�=8owե��3?6�A�..a)msq����E &�5{�=9�a,s�&�t�c�_I��+��pye �ᨇ 6�8����㘩G q'o�k�s���ܸ�D�v�)�lD*ʧG�P|�]qnHr�2Y�?4n��Z�"I�}kK�9_!�R�(�O��4�v�L��PI�����+cs� ���c֏�׺F�*�	B�~Թ}�0?�`6I��*��2�DI��+���'�IN�;�C9)� �8T�ZiT�1즄7FbHw-s��*Byj�92�s�:c��<0צ��n�HK�JO�$3��&]\��.ꈫ�cu��<�r��x,lxR�)C��2L�ɤ��P�>�)��(h������o�k�\&M�#O���F�����i��`I������@V]nr���9.*\!��}��Mh�W��&@vAm�z�j8)�T�:�NUI��\49e*_e�$Y�o�#��Ig��6�}k��왔���T��<�g'V/����S\�0��	�_���o;�h�}���ֻ����㏰�Q��"���{Y��~G��N�j�џP +\1�A0q��d�����ƫt��V	�栳:u�P�.�[%��ߍX}L�z���*E1��;�1��Y���8�;ZG��!�r������Wj�8F�$r�0D�y��>�pnf���8ٴZT�r��U������e!]��@�8H���/n	4I�H����23��+���J�_uk�!�Rl�����2'�π�B����tP��K:�����c8Ȯ��j ��F�gME�d�緅���)n��#l�gS2��]��,N�����i�K��H��:�]b�xj��B���+)'j 5$�kyG��pP����f�鬲���_~��0�L��k8���w/��BI�U�,>L�|�y�8Nrp<��e�A[�$�D�`t?���`�����#�y�$�J]Na���.)�u����]��P�F:�	���o� �&ͼ����O��G�z!��@Mo�J�H>QC�pz�ڽ��0�İ;��bV
.`S@	���IJHM3�p���fĀ�U�|_��u�?���Ɏ��mYC+�.�	���1j|���zͺ-:[	T�`���$�ڷC7����A:�-<���	��e���gM� ����gS$n Z+��ؙ���T���_rzB���H�Z��̰��{ÜL�A��cR�3rh4Q[x�M�b�$|>��M�EȪ��,�l%�>�(|�}%V��2����|x��;�ell���<c8sw?�̧^��[x#����㳍$�p��9��SXP��/�(��+SK�ԁ/�����z}b�~E|����^�H,����"٫l��'��6�J�D�9X{�:Y��u�T�)jkp��AL�2�Y{��-�u�ZF�Ec�^S#�R�g�ĳ�*'�w�wꉀ󫕄�(%��&�`ݒ*�u��伝�,s����������a�*�Z�k6+K�0jJ�˷#��
C˃�hz��H��۞R0�)�Z��)����[)
�K0�
�^�7��@�
A���,0zS�wHl��;]���,�J���Rſn�5^X{߀:��G %�����-��+鮻�$t-�_߭�3ou ��>�x �Qe�e�"pNԜ �S�U����(�C��E
 qķ$��­B��0;d���{c��y~N��,�r��n�ɺ����9m%�0�+["��r��Gk��pӱ�-���9�L�]��?;�.#��<}��o�3�?�DsT�~�GO2�>�D3�ヌ+�)�ʋ���O�͐���t�