��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<?';S2s"|��������>�A=�L��'I �.�:��T*�����/���1=Ȃ"�vEh�RTAP�����a�iG��6�9Aԓ��,㊃��;Dp�y���\aޗ6e��NH��l�8����(�[ ��L�����3����%X�!��ܿT�j��8ȸ�I:���B5��>���ivH�#"��D��D#�fP�*��Mה�"�;���0����є���-�@��s��_���%��C0 ɛ������g.K�gЖ'�9��+؄��Aה��c��arn��/|��y9� B/%�;<�Ғ�!؅S�I�Tw>�[�3u�X�D���R)< !,F��33�%Anc��m�¡{RSf��6���]p�|/�ș��&؋v�O@�3q�_�x�`(Vc�ʋn�yn�8��x�s�����l�m�ќ�e#Cb�����'�"������v���W.���?�Ĝ�f䬩#׿о�����"�:�\`����$��� �5k�g������غ�q޿����V���X�N[2:��3�V=���9c#\�_�0�m���$��7?�F ����]W�A����_��E�0vP8��-��Ġ�~^	Y`Z徍�fi�ړzO
 :����|������h�)���{�_����%0笩�rȳ�q��8	2Fgn�>KɌ��@�����9�	N� 2 �b�~�ۀ�$|�r.��^�Hicw����eu<<�V �	�C��?EC5�����ф57m�7͛�����3O����0`��&`�ï0su���O
�l�N���.���d�0�4r�^�l�c��+�q<հm�n�q@����bm��4�>�M�tT�n��6?���D#�����F��0�����~��/p��� h�La�S�t�]�YV��X)�ZDx��6�Jo>.�(MY����F*}�3�dS8LZ��<���'��1{��I3���RL1��M�a���7�?�"!e�jx�� ��]�O��Վ ��@� ���g��ąL	�)�ģT�"{ "�@U^�B ������R��#�m'-�6Kj�%bКn�7?��y;��nU�Q�

�F�/JY����� �v9x��M/P�����4ZSGi|u{R�<������Q; * gzMߦ�Q�{�I�5h��T��W${0@���B�[SiHmʥ�#tN4�L��� �|6�6k��e�	�` U���m�@hŐ0�K撞�緐�&)����?�K8,�H�f��X��H���`>��C���``���{��
̃dI��@�V�X��f?�w+
����TS�����H5���ZC$�L3�$�����h��x�@�yN�w��590
O q����B�!gcC<!׾c\u��_X}U*6��y��g�f��jW��HoK~�d���NKPEC�(7�QR��kvD����C'~	��XG�4���-�[;ݙ-z��ɔ�G�c�:�G��Ϣ�$��y`A?\>�0���m{Ѵ/q`ގ�&��3�.�zݴ��]�� y���p3�8!pZkF[��p�\ޘ2θ �P��x�ݳ/܃2�}�'w�����cERӼ��^�Fp�"�g�N��@���O�9F�wΫ�
qK�Ի�$Ϧ����VI�
�!ձb��M ����x��*���ch���2p5�35���V+��������&�08�S��-� �l�����e�@9�N���]�̨l�|� ��6��(;W�`���q�)$O�O	�IU�&Xs=�x�Ѓ�V�ςs�>�����y����e:���&��۩�V��åċ��\o��
�`��O5m8n��R�FI����FF��T�6ȏoʦn�U��[H���Ÿw��"K9�Rm��d���p��nf[^��n[��&�փ"�/��f*	��/�䶾���?g��b�W�k!�S'�5�ՐjE��-]�(<ږ�}Iw�����@���*W�MX��F��Φi�ÿ3Y;��"���tq�0L��+4k� P�7���|�x^{N�(k�t �eF�j�:B���xS�����L�W�x�4�Q�ܕ'����N�>f�*�9�!�@U�pBX�@�v��QܨS^,B�F��.!PA�$_��Ww��*�lma�<&�g!'��ZؐĶ�r�*l@x�U���TK��[&�'2>WOp�s�p�B��a=���s��J�-��O�9]������PH�J	s&Z]�����c�sY,��R4Z��-��R N]����/~0�,�E�DX�ķ��$���~ǱE��7��.L�|��ٜ��'�n�&h?u��Y�P�]�rI�(B���a.77��i@^���I�ls��Y�5>�>�^�����A�q4��u�)��r�gƑweT���Ďn����)f�(��Uh�o���Si�����,���< �_�sfW��[{�}VԆcTn��R�hc*ɍG�P1��Ďc|'JmrS7�ąI��1��s/�Wq�{�8����LN,����%���T��$�Ǵ���h�Xn�*��O0JI]���Pۤs�_���Ӵ*dsdj�'J�I�>F�c��ʸ��l�~�g֓j�T����;j����T�bi�����]��>����D��e��o�x��;I{W���`���;8*�h��e%	75�Q/�zOu@T��JF�!�r,B�K�D�h�tR�	�YC��l)�� ~	�]X!�߬��A[?�%�&���ots��ϛ�7ߦ�gn�#h(q݊��.�m���߁�0���mz
�X{H���8�N 7ٜ*f��݇t~��I0�3��z�P�C���Yw{�2��;Ԏ)%<i)����LQ�}K���s7#mhi�)��y��犐�x;�h�ub�`���VmH4\��^���Tz{a���z�쌉[�5��ё[��WX#B�@_h���������.:nB�:m�.��
�q�c2��i.�=�O�q�6R�ȓ���U���`F����y������ׄ�;q���J�Jyt�O���W4fm���!��&�8H���b߹7l)+���;�I��w��\v��
v͸*�ܱ�'���5,��v3��^d�����q���Fцi^��=�����i/Q���5�vW8�|Oԯ���,D�ZQ��U�'͓CJ��C �㭊��@�1�5�����>�y��meO5_�h�u4���P����y�=
�K��x� �Z���u����)���Q�i����3������I+���(���~k|��>��~�rg�e�RΒII��\��/h1�@9�\�b�YW��B=&�<�����\���n������J�ҡG(��.�O)��SW1e� ��ǎ�\��z�i��CZ�/D%��`@�5D�1Z��a�Kr�@9u��v-*�������"gى:�n{��n�t�[��V�͠�tu6�$[�b��ψh�g��[��QNF3l�;`�V¥����9���������/,��Eƕ�<��7e��c�F�e�wd�d��N��6\ Nj#�D���I��o^S�^�d��Rq�2�I6�}�V���&�d�*>������������%!̷7�h��R���*���'O�������6Y�W�ǫ������U0T���&��#_URn0���XyĆ�ֹ{���[	Z��?���E+ ]�Q���47���W�e�CӪꈉW�ƹ��y�@|���x(�J�ÿ�f��=A�v<��-�rb4_a�3�*e�n�J�q9AE��ߜ��
�j��F�%?�f�������VXv�='��1%�$�h�?��(�~n"Y�o�������9%$�V�'  Z�M� 4lF�����3kh�}}���m��S��"5��IuVfs�ޟ�Zn5]q�'���]��!|Em��*���"Kb쌽٣��&bp���=�i"�-�z�Q��FU�h��?̼�
����w=m������?A�'X���F��k�����|�^9�q�&��X)�tI�F�t-��h6�	$v��c�^����z���(g2�h�/�G�P߈���S�ߓ�1����-�H������>�A�&
]�`�S��N��O���b������/<-UR�@q��7honk�k,W�
3!���=ڼPe�M��EN�,��������K����}���&����B۶¦�xV��89�c������׮/���4oߊꊺáƓ�l2MdC�`w�z��X����w��-s�]v���ɅS@_|�!=y��������zx�A��H�ج8<�#p���N�q=�q��.�C&)�[�������+!<6��I����#�oaּgE�M��6�	���J2%Cr�q�r����}lȗum5U�ۮ	$���ș�2��;yf^*�wK>�������.�-����$�u?��w��I�}<���,R�Ԧ�bxOX�M�I�
�	�F���>��u��*y^'����r�ަq�U�E��&�����s��i��z����'�`�!�={�l��6����c�;�8���]�{��!����+�Q#��.������%�\[��D��w.��ʑU���,���[��4�K+8+�)�o���y<����n�Y|�vό���-K��a�-J+0�-�A7L���|J/�1�1TX�Ϻ��Lq��E%�&�u�]1��<������l�0g�N�>P ���?Ɩb1�b~Pp�>X��t�47ސ D�0Ң�ҥ |\C��⥗d5xm]3|0V�q�?��f\��C+�?�R
�娌ȥ��������8I㑉�_փ����N�sZ���@2C����ϯ�p-B�31�$O܇M]f:���h��.��c��ֲM+��-6�@0�'��0%k�5O�P�i��aj�u$o)�����R��%��ap�l��ъ�&�S�a�����5\�`���ͻ���!�)�>��?���vc�n;��x`�j_�w�֡�%�=/~B�s��m��Q��Ïs﴾:7�WQ��=���8���=8�"5Q4��e6��ؒ&�*��e�#�:�!����W~;����q4�����ED��i��9�d$��]�������3��6J�Ml��*��N9��j��]�fq-7%2�Y*b�R\�3����%��E���:�佺�{ʳ�F7�%��"�A�/s�\<|ch�{ƛ3��$���O�V僞g�� �\��z�`�J�W	"z�H{"��J������$�e���C�v�!����Y��m=
��23�KB��w����W�
���JՇ^��Q�%NM=��W�n����0vX��3�)1���N<Р�����;	^@w7�vz�1yV��Q���ݼchȘ�jlK����)��d�m���E�����"#����ҳb��5���,�,���u��}��C�2��,� ޷�ƵW>&�$�E��y㎏���ˬ�y��7gO+s"�.Bm�yܨ*��ߙ�~����a�94wO3��S���e�N�^M�H�1Ҿ�p�̮0�����#���$�<i�3�E����5y408�w�v��W����C�~��'_ĲM��J����'���xH�/_�R��ApLnd��..�Xu�%Һ��J�i�7�T�o�Ǘ�J5���V��m�y�vۛ!g7CU&�}�����ӀҐ62յ��s����qQ г��F�vV�Š�䫮��Ң�_��u�d��2�@ЬM;`���6t�L 6m�~�����+V��Y�}�(:D~�)�DB`[h�n"���‗�%���<m=3JNW=�v Wy���))"�Y��G�㨰�L˩\�m����$3U��IA�}�A��AКށ�0*�y�3�'*A��~�C�Z�u+)��vwL�2�3E��4,�bz�������/�;�jܒow7�~�̋E6:J�GԔnʲ��h�%�F�9zQR/sR �vh+b֊mF���Y�[��ݒndf�,�yn�
��_|!2��9�Mn��@9(�*A���5gw�qy�gX�f���L��>��0I�J����aj�|BE��\"��Ƀ+r�F�4�ȃ�twL�6i�'�Vk�k0����g�>�>cU��we���
�x�����YH�?�a/��Oq�2y�&��Ҁ�Cx|֌R�Q�ɹ�r�PE{_��w��K!�^nsW�)��_���i�T��4v�t�֛f��[����*DD
=H,�J��Lp����)�_d�Jl������D��-��KH�D�$�t�M��Q�;_���z PX��~������
v�Q�&�0&�ݦ�"vQ4�hHS��®�d-^W�uSU�=X�{&-D��É�p����Y�@�#����U��z&b�^f)lt�<W_��2����
��,�'��]�$���k ����nPBPP^gđƐG����]���J�=�h�,uzzn�"�����`�&
��$by/o��N���%�f'�&��A��hS�9������5''�
Z�a��P��O���+��q��bx�"���Y�	�eA�7�ۡ�1��,��f����������i���>��[K�d�Z1��/���D�y���z�
4�[?i��2�Y����7�����#;�
�o��bH>�+�0N��=�K�1�;6�!x[�D���E�!��?W
��Vp��L,1��g'���2N��0&?����E�6�<�f�|������\��Mq�zfpO i�k+7����,�L-��O(N��]C��򷛯���ekہވ��ke�q���~��"��^�ķ@�ѵ^�� C<�T0Jn�l�R}�W�D�{Jn=K�d�4V���ū�L��J3l�Z�����<q��G)=�o�ŭ�W��J�T�s�c�h*�Tk�Y|�A/�'2�S�1�P�k�A�N�`0NϜ�!���N>����]o#�(��F�6K�W�.i˿V:^�A�`��:z5k����W�.>ma5�f��V&��qX3�iC�3�D��b��C|?��R�$n2d�2i��!<�w3\O1� �I�Dݘ�Z����5��ڔ��
�SE��`bE�Z���j)�(���#j�w^��N`vL���n��S��E�Z%�S�;�NaR.,�?9�[9-����I���.���R���^>�u��1�FtX`�/�2	�u�h��6��D'j��-.Y��<ٮD>��&��ʳ�3A�<������GN��?:��;�EQR�m���0=��%��Iq�F�%��ka�M%�+���ZG���ʦ���>�R��lP��R��+π�v�N�_�[;�ko�S�IB�	�]C#3��	��Զ-[��o��Fr&������*=.4��	� ���G��Z��	�&�o�Y.Y�Ч*9��)}�N��[���9�ѨbP�z|�rm�Su�v��T��R[��p�:p��2���^�	��dH[�\0J�Xø��ѡ��=rjK��S�Z��*�����rV�6 ���h����h��$k���ބ��~_��ؘIw%H��>��%�pQ��Ԃ����`�@�;QT+ۭ�����[���1�)�0��5S|�ؔi,��b8����2��}�ޣS` {v���@l�n���ͧ��cq��b�e�$Y�(K)��գ6�oΧ�4�� ��	��m�K�x�jM^$KC!B2��w�^��|LR����!r^�.T6��`�~B�h�	�$�:��߃��0�L���׽P	�&��Ƒ��B9���h�����2!Cw#v�P݊Fb���*�ĳջ� 9��rݑHr����`O�<�����Su>��0��\�n+�᩹���0��
������`��䠍uh����/��^��9'�,��]���9�q5
(��^��Sn�/�!��3η��e��#h
��uI��+�TH��3/w�#;;����MdEߣc2�J�\H����.=f|q0N�U-�OpN,�^,���7��7Ӳ�$�C~��Y�F�i���8ͨ���Ǘۊ^Jo��w�239��|á�P9���dPQ〹�+7k�~D��y�"��Np�k�%"hvH�5l^n7(L3Ww��9d��ٔ[�Z2.R����d2#}�@k�Y�&\�%֓�X�}#XJ�^�
R�x�$�j��a�e�!ue��k�I�a�`f8Ѐ���S��b)�����]��:��X�)1&h�*�ePћ��F�k�Y��Q�L�7�.̪6�4��
g+�5k����`Y�^H�`R9�P�DEy�ʗ2u�vhH^>L:�Va?e�Q{klAE�W�s٩΅6>�@/���Y��\���L;3�5x&��b:�b��E�c�.Z;�苽�c¸��=��Ih��^�"�#֋���z����f�~�tC�XQ���}��p�,\��KV������l:���y��ю�%iF+P�nf"��*�%��ނ
Tʼ���c�J�G3�����59酇���~n�0IE����R���
�B)Y G�!��{�0�Gr,	�~c p�����Qdodw؀Zb�{#+��!���3�]�d{�	rs�4\�Q�L��`�F�{"�.ۊyAW���iW�K��wwd���2+��w�t�)K�p5
��un�v��-t�����R��`E�zR�������Z��=�Y�Ȧ#�=��T޸e@�׺d���ppS6���t�2�㚠�| P�<5�ṱ����U�㴟<Lr0�A��mW򺄵֟VE�f��0���{��ǻH�z~; ��Z� 	*y�n#��4�SQ�{��V3S}S͖����c�E%��qh�/s2f�ND����z�H>��rzq�Q]�x���=��mTy��e`�+lb*���\f���t� ��h���a���w#�[W.��*(�'"�)XOо�I����0�N�c���G�4��m��}:R�=eM�5S�V�;as5?so�Ă,�6B>I�I��Qvv�.i��&�i�֊������tH "��ؿ��3p�tA��4������"���D��>g���t��@R��O|���俼��@R�fp�H�s�l�n��̪is�R�xz�Nb�}�O<z�L�^o¾�/�����w2���s�t5[�{պ�U�z䆺�򔒕���f�Թ��>	�̀ٶZ�jU�����mF6(gZ�D���WpK����&w����d[<�޲�r멎����ږKō���f�8v0���x|9h��;��F���� �^��.Ҭ�ϱhi!�h�圐�f����3��|���T���[߹(~i���(�����h1��2?�V�5?���^�ht�+~�y�"K-v�\Kމ���F��ͮ(A��}��L3�71+� yw���