��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a��S]/�k�q�&�S;�YX���LҮX���iZ���""ԈZ���ރ"b2h��ke�k�Qǀ3x}��m/r��PM��%&;s"�X�x��<Z��tˇ}�-�Sn��t�	��V������"��l���B�	�Kq�0�p��^��\��f�U'����}��x�)�ۍ��K�,׮��i5_�%[�Π�>��ڐI����p@*e�����f��m�:lh�{<��ix����&�4WB}9	�|+Rfh���T�Q��d��/�K��#�3������g�ئ�w�4�5��:o�zO��vh�w�J�#?��r%Cb��4
����	7o�>�ֱc�	/��w/�� �?�����V+���G��o�X�-2S�	�ݹ8k�F?��׸��Ý�5�$v�V��:��`�+§y��<�����Y(D�aQVѱ�|`4���w�����Pl�[@�
Ѐ���R_�������h!���i����f5��8t6Q�̡2��4��%�r.y�
i�s,Ld�����]w�q���퍔'��?FB��Nȋ��'�.�s�O�$�!1&ﺨ,����vm���zj�+[�h[��/Mx���P�ݛm���J��j���jS[n�CENW�"9-�];�mwv!�𗝡��S�F3[4���F�un{v_�4������'�{ΝV_�_�y�fcc�/s��1��~\)�%���,}�G>>�q �v_9&U����G8����X~�ƽ�J�ĥ��؏��*�|�d����	R[��8(��H[�ecT`�#xzF"�J�p{����=��Ӄea��>����!�o��,&#���nPV�TX�;AH�(��/�\N{�0�6v���R�,�|�]�b}3(q3'<��r[;Xm���G�4�ƥ�]��ZyZV��=z��P`�W!Crnt
���qho�޾�Y��v�ΖZ�t�9�cj�P5/1���Zb1V�X�C`�.�:o���,�uDBB���@�t(p�����R�X�u>��̃S�Do�ӵd�W��r9)<�<��G,,@��8ѧ���:���R�y���I=�.��V�(y�l���vG��\�]��e������d��q�s��?��T���q��M�7�qg ����F0;7IV�����4�M�n��<��%��"�b�fJ�⢴X���
�W��pI�D�w4ʉH��7n��)I����=g����hP���D��3d�Aa
c���U�2��w���ܹ��H�Ij�V�>�J��[mD�Dǳ�'�8����Q�f�E���S滽���)堙P}�����s�c�U������� ɷ�h���G��wfF�gG6��>_� �\V����/7"�k�L��k��!���E��	�ppx��d��F��Jܤi�]���2 m���[�tō�LJ��S���c���jj���������Ƥ��筿+���P)$��<����i�ՉM�xzP����a�ǵ5�:��-����d�)Ė0�e$�ȵ��-�[O�d�Gh���ٰV檜��饝<?�H~JVG��������Ý���'ο�%]<���(�v� �p��S�@y��� �Mє���٫�-olP����H�3Y���������Ƽ#>�	0�<�?͖nd���R�Pͪ�%x������1�s����$X���J�]L�^/H�Z��së�U�Zw.{H�<~P�)���$�(~�vB����!���vr�z�q����u��k�R���{�{��*����y���"_{����T؝�@j��LgM�llr�3�t�@		�$���6���p�3껕w&���|g�I��v��A2Y�L�Iޔ��Iv]�23۴�v0��\�RԬ,�������P������-� �)�P��#v�O�Md�-"�Ծ��S�,PSq�HsD �6hL���V��z����P�:���9,��{뉌Ͻ*f�U�����"��e1���ٻ޿Ȅ��Q�brW4>�vyy�o�<t*�3� w����Yd�YN&9�BL����Ůs�P*�1{����}��Uw�F�w�<��8����$�T�9�|�o�~�4驵��Bd4�Nʈ�+޳	褗��j�B�@�S�<qBR��3_�xC�����AZ���A2J�s������2�.��^Z(�����C��ۂʏ$0��?�a�s��h�B±�B��5��J�d"��U�`��˔?/�n�ǝm��w?�N��sq�f��������T$���4��y�V�a2�)�W���<�M�3�֟��X `� ܋�F�M����}�ۉk�J�	g�S���m?���[uo�{�/�;w}���"�1T�����<�.̓�BAJ�(��S���(�X���?���1r���n�v���sߡ��O��CBT�7v�ȋ��7��H��V}�[����'=F�KΝ����v�3�5���;%T
���B�"�=Āk��zKeᚩ�| b�W���UR�n��Bs���xŒ��#,�S{��C-��;`��H�T�B���R+�� M��������wQa��zQ{L�4��#ʮ�]��`g1)��5慸�u��Cs	Hu-
/xP%=k�]��^7y��"�zT�\Jh���7|�N -zT$�n�^w���̂�󼦟���sϽ�R�t�le�
��)�����0�w�(����+������4�����b$kt���/%ð?�Mo�c
�sV�_�슗z��xl��oo�r�\.�cvT�x��w����g4��&x��%��L�}|O]�q�1��G��c����[ppO�����n���Z�?��3I`��"�Y�}���[8EC<-�&f�]�i�h*��{�Bh:�9���8'�u��5G��Sl*�\��e�EF��C�����_�z���>VB~E������7>�%�{5)�؟���Qk����`.rq��ܘ�4�������2�,~ŵ���M��Ȕ�������X�!����C_�u�wK d��~��g��_��4(��^�|qQx���a��Ǧ���`��d���=`Z�1G(L��;�=R���g/��&-���f�l�Ĥ+;�N>�V�o�eC�-fgB�ΰ,�ٞDB��Y�;봇$��(���L^���L�ԥ�y��Z�;9���(8��֚��Q�=i:h<��Fx'ɠ�n�`�+NO����&��)*G�z?�����k��c�W:����6���h~��M�хB�����iz��I3CG�������"���i1B��3Q�����~z�@�,�@Z[  �����ia!�L�����P7�����}0Bs�2Qn�®�������������	sO9|T.�)�=.ε��XӅ>J��������胎�~h��O��V�C>�2�>d�7G��X:��<������7�\P�����A�2t9��ij��9K�5��i^\�z�:FI��z+4��t#�A��qzպ��ǧ۞��&�	a�ɦ�5B
_))�g%���7*Bu	ܼ+!г��G���}���N���#Ӱ+�9�#S��Tã��?��Ȉ�U����ޗ�1uń_�t.��t8"��̐ Q��}��Jz(�-~�`��w=�z��M��v꿲���L�^���h�gU��)���N������j2z�W?��f^���sߦL;��Z�Cք�����]W�{���D3�������ns�E��)���4�n5X���n�R��Ħu���[���VA*�(g6���X�M	�^f�19/�[HZT��t>d<f�����d�j�Q�� ��H$���l�4�a8��@� �d�ny�e�ᢞ8��G�i������3������\��&Q�xF�7���rҪ���OQUd�{
�*I騏��»8I�T%~��3�|�&K�?v�Ɋ���w^��=cc�����%^ )�LHU���)熔eRV�'g��[Q̮�f��K!P0=$�\{�^ͱ\��{�1�u���l��X2%+m5�7���N����H���E�\�x�K��b<�� �u��r@�_�1��;�ݓ�nc��Z�lg���D�� �ђ$��$]P��7]�hx����O�#HA
˼ZdJ
��Ua��j�����vD6<�܂����������L����y �pq��\�d(;A��|��#�*����y�݃_Z���5=C�N���TJm^X�Dn�i����g��ߧ�-�3�<��@W�ͳ<��xoBr��SӔ�=�Dk%��}�E�c�[�֗q�'�͹�;�*8���C�l��[<�>T�wpI�H�]PH�Pڡjun����q���E�a����§w`"���3ʍ�gWy!�Ai�{쩕����A�ץd�&�	$o��.P�,<�O���3�d�mU�"dn��&���|(�D!�MCSF�[(J��vp�<�E�GE1T����M��iڶ�u��z�>-���n����#v�G*k�I�Ƴ�6�_6�VM���m��Q�[�⾒ﳱpK�Y�8s4�{p���8Y}�s�e�K�A�r�j78�<��MW}K� ��Y�T{�ͽ}�9���+�9:S��^�::��}�>h�LM� Jj]�~Br�1N��{ޭ	�eg���\_���Y:��7����1�#p�iV�;$��m,r����͗C%��ㄿ���FA���\�1ʛ����R�(��ceֱ�#�᱇��6W�'6�wy"|�I5��y�%��{��Agǒ�! �/�sJ>{���z�"�����q[�����w��u�/i*A�Z�6�ڱ�M�,:�?A��<$�ќ�PGz���	\�~��e����#�����������`!i�?�J���C4D�A8��k�ɱ�����Rwro&phD��~�����} M��n2��ˎ���M�+��;�Ÿ�U����~T�����#1t�#3:���E��r,�ҳ���;(S��f���Q�AME�6z���`���̶}}Y������8�,���oD�9�ƲUz�4P��)�����3��J����������M�U���8����