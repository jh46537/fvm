��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@���C�X�-.c~cX:�,�B�Gq8z����� e]�OTS/�vh�Ѧj��c.Hx����:B�yjdz #�Q?�HXJ,'��1��F+��X�n)b�O���iA�S!0��M�.Oi]|Ц�ܚxx��0� �i1i~t�td��DK%��s�b��ܸĔ)JS@���A}DZ�5m���ז��6���0�|������{U��m��ڷL�0a������-��R�u{Cm"Tz>�Wu��&��Q��<H��{ޣOY����QzZ����1b��s>P�i��EQ{Է�t�N��|��6���:�մ�����/�kp��Y3v�i��Z�/LR�1�_����L�_����chd�Oۭ�;�3l�k��L$�#���F,�>���VO���;Xv��j�:B#ʰ�2�Sŗ/�Tё�����}*���%��{ڷH�>�r0G%+E�#���e�/�Rz��,M�v��9����?�*��n������h=�U�=�!��U.�d�XѨMÛ�ou���}�sÍ��%�"�ݖ��ꍏG&U��<\8���h{)X5/]�ޯ�66�j���e�w�.�MY�ȩ�o�ab���[���?�{)?Կ�^���q�V���5�!�KZ8�cJ���}�QZ̵"��5�����,ML~�8���#I>+�(�oV52πR��U~����O�ĵf6KG������D��pD���o���n�k\��6�|��V��x�a�e�A���6����߸�7�e�% �Dw9����~�h�`�����g]�秔r��g?��J��I,	���È_��Y����=($����*5��I1�BTb6 �����Q���f�������N@�9,
d�{eY�Ò�/�U�Di��a�\��`�/7(C۸=�D������lH������.�/�>z����'����b�.!x�#�9�#h�j�*z�z�e�b��3�,8m����N��f����J;P���s��� a3��g�&�g(�G��獣����@�����}B�*���-Ur��/G��e�t��A�S�scu��7����	�����m���Mƚ_n����h؅�P��* BNec�N�Qp2ϥ�y��~�l)�n���<�}��É2Z�DY���ױ�s��L0�y:oa[���z`��Z%ʼ3�0$#�������lꆄ�y?�NF��>��:�bh(p����W���r���O�{�PH��Vm�G�W��C'�$a�M�R�V����,�^>us�B믫TَEq��Yٲ�ү��\�r0'�����"6IH��H4��S�7Ź�T)�*��k9��.@���q��+F��h����<_ДkEBz��6}ǑX��4w~m��e���p��u��q0���^�r�d�6�"A�9lJ:��ٔ��QC��~'��R������\:x} ��~�y4��Z�4u�-�G��o�8�f��M����1�Cƿ��O�����T�,8A}6��6��]��'1:�A����s����b%��7���roC�F��{"���=f�m��F7��%�ZJד�"$�y��������}�G�Z����E��Kђ��G��������,�>���FJ�57&�}פH��I�
��}�N��/ڹ�*��@����,p�zr���uD����JO�d`�������c߅}%K_�=ܑ�[~�wW!��φd�y���9��{�� I����O�K���̀pTD�3
��e<��������KH]�	{RmE�%lF8k|r�#Z<���}��o�����l�yCΉ��E�K�	ȍ�q�E>�j6)��vm��V �ȼ����+�1�Y;/3s�e�[���s��Z������(�*���+5;�^�I1aZ��Q�q��Z��ǷgtC���6�W��ʪž����ƾ�l�$�%3�Z&K�]MGE�:u?��[��BW�d�x�o�b_�y�v�GʷỊ|��f7�����	}�@`%�a������7�U�8Ȓhp���t�����ӄ�E	
�{} @��u~{Ɠ8yvAa���W�]��������>D������Ǽ#�!�@�a:l �ظ��s^���9�#AQ��~^����y��&��[t