// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:40 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R6dKhuaGenrLT0KfOhvD9kEFsjJW7NjdYAmhRn1FjaL4918dEfkIhNhtAyFYNFE3
FQS8MRKJ76fLPmm2DVnCF8HyxW0/paipvSIxW6NhuCiuULcX0Wk6TapJ21bhRQON
tgWRbqPCnpvPpUKu1i7LEusdAIyAWe4u7qccsa9SQCk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21872)
qek9LtaoaxolOwBRL6iBj97AQph+BbVSGZ4vI37yviKdAbaLYEOsedG088aIaAGl
WllTQUADQ7O+0obVdd3KRtTMkSwMQGFi/QR0IJw0LhFkUR+jF3WeGHfmC7HMOQ6N
ugxzKCqiahsaGnwA14OOH75DVHuZY1O1zT74hgG0N6I6dl1Ko0UPikSnT2zDj9fW
AzOeZG7c3Z1IzxzEK4tsyMk55dDKgKFw64w+x7Zr8qNfUTZCJbJPN73mdjBUxuq6
1Rs0uRMzqsmc1DncW/KyIVyoqQv9P/Tbo9x1HYH85yGXSP9CbOF6CsLBb2GWAnlO
o15n9Oq4/rH4jEG9FnSHlQB7+C7+nwTvLbE2XtqFh5lv2h91MXnoJ29ecLPwYOJe
U6j0ceUqAT4HAw05aTDhSYza/gAfd8pH0LwyTR/QjNjbY1JWk6Wis9S4ooqqH2KU
ToUNDXWGcyVuBsX0XswDXreLvuhVRnd/lHG16BkJntc4s0gFDztZSzWXgD8B87SH
wQH4Hddz7vo+R0gtfQDjdC7vCMa+KDW4sHn1AzNnars5gfr7YUp1GDzbXMKOxbne
UiAaS+Y3aL3OdWtRskqm0uKCwRDrJ9T5iga6tVjSdWuAJNZeCC68V8vsKvos0rza
QBjLu46vE3yfC59etBD1CDjZIVygUoNl0FAwLkYgAKdyLmBifDeJ7GBa6dKv+fqR
zMTf6xdl5JSQMPY1eMQgjCy0IkQBjWSLph1jR/bQjCOfVqK/YEjDguNokbM/srp8
9Nv4tuZTVsrBgQyN94jfA73ODV+MFrACpAyATtaP8bgT/bdN08U9dqqNOL6gPqds
fO318yoenIn/8gs+Apif4do6/i4+IZZKsa1dmsG89/lhGLIqD///D/AaZTZqk3Ef
79v1VRUobdLieI5KQiN0y4/WkyuPeD6b8DB460Ev7ch27UqWFyNywa+V/Ea9fdLp
Eth1NCiJ6N4iTkM2iXoh12OfooHR5VZlRgw2aM4D9/4e+soBvryL65J2lqx1yoIm
1GXdHCjxmjmK1dJObs6r8s1GGJJ9tOaLqQJZp1uEKzYhaViFO3LOoVFKNIOotZZz
xvymE2qI+BNQH/A5sUJVDTQThFoyD1hrfqDJOUq+tFcYl53YLhRZDsesKSQf1arQ
Vg7dzC65NEtNzVJH0W9a9VIg1+BvQyvyukB452rteaVE2vLMk2cuIwpKK8MqF9Iu
V7eaLQSskNB5c9Z1658eDYivdYc2pzP4LGoDnb9SZs6rgOoc4XeSqs52udpsKy7D
VjIiyOJ6LNusWQFY2LC7tcMClSbqp7jhD5Pe9KFYjGxH6sTgmiFyj8lKb1q2LPPr
cEY2ZlvwOEA+L1g+AilrnuAgrY9aL9Zl9Xd/xG+ZoSSAPXW2m4UBP8jGFivOYM9J
BIW1GZLjLMOITb12QmPAhxXEtsUF8YafkunPXWD9dGi2+9NdNz7VZMW9sqaF5RCC
Ea7dUeoRVWEvL97LvQb0UbPiNKXW6cO1KNlKnAPSDfNkIhneHg+jRZ0CVzHqaNDC
GtKVmtZyBMY5nrZfzs7DF7nDGFhEHMWHnqaJuD64adgXwGYNtSmqRmYuYjY6SVCA
dW7x1HfcTmj2iKKoICjulPkHOY65Lq8FiX3bGhvHuDEYcnwRSR+0DSJ5DzZtK/gP
BKvdpKFf2zZ7qFgOVU5erd7dSjavpt3vec8HeGBsuq7sAzIsjf6dHCVfkeCOuEuw
SCggR4vRhhAIlzvvHnJhFhMMs+4mxQEvN2XQPQNrPDSVHdkA5KwubYUBkk4zWMxx
XBfJ5HTvZkLoxUObM2hyXDqvVYGwgCFVz11Xmg1Whb2t4abFBmzBMVXFsNpV8noB
i604GdamUn2VTioEVu9MZaeS4zHDalUsnqf4Ias+8Jt+/J8WZDUOVAN/IKz7OgNx
LglFStEgSCdLsfnOz+MXesC0AqkvtD9MLXFpHntDsgan7cGm1Vh3Yhy7IEeUGkVn
LJ4J5z33l8uUmpQIzTUDbdO6UxeejsBngj2QUThSWIPm845zqhXrYSq+CFOw4/yS
9D/PV9K1KA87xnRV7YXH7wt18X7bI66pD7kSs8c2gOUpOQWnNRaRcnZZVHSbm30C
SQnY4thnM6/emWXWFdJmQ/uOvAwYj5DWL5QN5pP/LXc0LsBy9QHW8Utd/qiX9nME
FaOUetXDFALGaCK8HnhrOX4FyHZYNB+4tqxdVSKv32B8L77nTS7HtxJP1ieplgkY
nsst7efqtGyt71X1OqeVRqw+yuTb1tK6oEJ5nOXrVHI0crqOxh8r+9n/0K6nWDzw
Bh49UfF+XuYn49xvtvXtKbksP5kh8W/HoBnkVLy8s4tRTBzZm4EI0IhCYxz7o5Dg
Zj7tzKfUUpdHl7jxze7MTTNly6vFgAQoHoWrKq3S0wGZ6COSydBWKY/Gs1HpAOzF
TW88tOaRTQVPAgNnzzN0LvOFQkw/7cdAx6iU9znLhLD9spia98nzyDYc4zKIoYgC
8Z3cuUEWc5sdk2wjk/rWObOHdlK6IxYTPfCawK76EBTwLrJaIK2vCF42AAQrfdTS
WZsgLrQNIBmMoEh5wolT+HFf7BghBs+teXUtVVTI5QK1FV6nY4A6uP3wHBZudgtS
Pqhy+aCMo0FjN3wjJHnexaDB06zF5XqewKGAo389OBoTV5VC/T2uNNQw5iIYVLU8
qnffUYLiSRjYvt+3ZT5IZL4VgQoCZWpiw+QHNyHxkXsh6FDHUQf2+pZ2IMbAWdOG
Ytn5OGtPOT5vR/AMaA4/G0sb5RCS3ABeFH2bUhjDxUF2QlKwIobUaLpmirqmBMrr
B98eL8SEusHCuSDXb7hkL2qSue71Bf17cBN3dhQSBjoaZWgLZZSMd+n2gz7y0u3a
dt3Fy5F0y2YDhWPtlE9hDvI+r51a8eewgjZzNLlkNyYasaTvwaFeMlJZMYb1Q8nW
L0YmdoLGazk/6QDlHdEePJH5O7D6ZWlDQvROfuQEC2mZEAMTYGbff2mKaLE1LZct
ycHEWGb5Jc4OM6wksxCit1l9l4ed77Fv2KLvNzW5QHWNj+wCD8db2v0P6mAqDg8x
v7PDZhgiLQxHLYEzcDxdJfKq3nnp1vr8X7txrghhHoRHckd0MMsQNsII1Z9WiJwK
ObjKcZN+En5dk1CewGbVC3phpSjT86TC3vgLRNiXEIGW+3dydzXBQOL4r9mkrOLm
yq+sY6g3XDYd5NZpHRdP4cNi4FK8BzPPwYJ+5OwFmpsy0BRP06MpUZAPKwcyRLeq
/+QN071X27HQ0fYwjweZ4tv7c2eNUOXMKPO5hwaTww+OVOcN3Wnjdkl6gNvPK5V5
NpudvcAbXtMuCnixcP20V82q4UTZ/CQf0UBCJpPOXiGquzN0wUMnWMqbQDFHXw6s
JwQX+4nnFxuGv1eCGruoQ99RI8tbDtslIY6YaAMFnwkShfdagZx86OAieoMLBZNZ
EoDb+nMdea6Dz8mP+xfJmERuY9EahxcxJjvSWWpdc4tcYyjVokerFuXndzsLw84j
I0+0JauO8DMPEw7XcoeF79upzTIIEl22zcT/s78+OHNpmI/18vaBozow3Tagj9SD
QV668hs/jmNPImtY+mcme8QY80h8LbQtEZa06gt/8I4YrBrPDsfqSOpFpX1W4hu4
Ajfl4Q7jBWHS7O24S69tHXVamv48tu9jpmhdfe2jzFDave6iRJRDTlEVIPht42Xi
3DHtgt5Tsy8hDRV26rR6W0W47FTi7M2NDfdNvhadWOdFdCFWkg13O6gFhazSwAy2
HlEiNoj1fp5UxrkhAaECa3qTI82eRLHU9PTW0FPmIxj29cfLjzsswe5ekBdkx1/C
1wdOzBur/9yXFYMR/9moKUsUsRXBRPP8ZcdhWBgqPwMmFKAjgicTiXCo+Q5m2x+7
++WHsrLsOCtCLOcV8Bo4Vb6Uc6Q6Csr9/RVTBVzUNZ/6kG/cN+IdXyeuS6kUBRVl
b/qvEXprcMUobdYHKbLI23/RLU8tuo/Xz4HU3Xblgxt7gW+ZhJTvJ5W7pNNlYaPI
oqBGE6BrYgHgX9fYr8vh5xh58uXMdxDpg28XuGKr0kjrxME9CH9MJigblw5EMcYo
2aCVAumDzqehpQxyyu1zLFradUnONzqjjQhK+JclUNCHSuShvfBIgR/n4U9vqeDl
iY6w1B4zlBrCg3RaWnr2oO2gxfBDVzr2twaBmzfqcVZ8twsQ/KWf+JuqPYqNuDNO
6gkwboTJxt1q98drxYFAci0L9iKLVbAmWcZKJ7XwTeN108pbTX9H3lpZyRZ2GUWg
xC0/xaSdT+p7QAL8fk0jH9dAAYFSwpj73Olr+qRLu9+6R7rZvkK67sarG/cpJuda
ih105Iasw6SiuFYIESOhQ0A5fZ6vMOtz7ejrefDzg02i5COh08GJZE0/40XYPxjg
4DHY0OKzHkngX97XTSLe0sQMzQuhazTAIdySMvyQExolxGR7WyXVhBZoFOFp06m5
IdpTTRd0oBN/Arsvdeca5mAW931peqNKEjdcKKea3+ax/FAHMMIV0N7d0fSV1dLK
p/PmQDdCOBN5RDXtzg3Id+dvXPY8NG2huYjci1rHEIWZiBGvC5vPyYWj6/JvOyH2
es2KjEf2PEYmV0wD/PEGFOLepKY6WLTnEgDOUWy9fb9j5uq3o3GOj2tJC7pyGXnM
01lpVEMEk+2I2UVamebLAB6llmHTeQvksgaZcoFEg3ZvUpCfqa30XgtemD8J1qWZ
1ZlwxxgiFUQ9DeX2x6olouqqwMIwBn5BhcWAkTrI8qQoswqgSkxxnvhh676/FFb1
CL9LhPGGqjYpDeMCPdGkYnP5jYvQ1H5pSuZugbW+kDfPFOPk2SsUF8RtEFVxnVzl
sXGwuXvuHkOQkIIXIGSv2m4ysTcFQWTqZjg1+YyiKdxoX8qinSjj2dT4d3K0EY3a
C/XFhK9CfP6R3Avv3A8CJqW3UWPd+Owt0alN6c7jqgL2sTmzSiFVl8rFPcGYtR5e
5X8rPHPork4OegL6rbLNiuEHolfmtwckEA2vL6Nqhpci9XxehNzHZmJiZlHviNSp
yfE/S0a3IWEyO818P2xWhM2DuydCv2bohMKSMlBN7MkVdC9tdBnxuqwSjQ7QtH8F
vQtkUc3nv0HIpAewKwDu8qhu5LqCWff4r9k5A4GoiUPX9X3IQF2m4oef2YIJH3mD
/KtQAp5Ca3FjnLnmqG/qZn9v3n4+pT0hqKB8HAaHTKoA0OEa6hQOv3iXyrqF9J/n
DzEzcmnmpPjAgQbUY8tpvJVErPH+w6fCTfT7nTeAMvWx4igbVk+sHMG4RIXAi3sv
h3OnQ45oUyyBSuh3ckY6rJhtbrzGUgbXX4UEBMA06S2ybcWhXHUKZ0UYu+pefkkB
ewN0zQQ2ejMomQ4i48K+hQWS63CRGUuT03uOindKFp5ceW4LKSM94iZaf7WQSh4i
HawRo+ry1nmUr21ByZhLosdtepDE9/k9B48VO311EkMj8YoKDHZnbTl1Ij2V7Ppz
w70PKUcSHJDiwhBkMSC4gv5Yns2WrcX5fZtaFX0NC4vnng1tfzioKZbDforBpqae
BrHmjoTCKqh3JAt2/8QY3HjR6k+ZjNGYgmnXVeBowmH4um3Kma91AXxDNZmqJo+I
sm7RQPWMNWAWB0qUw7OV+1lCeo/O7b5LgxXNcGImvnig2A0NrEVrdZfHkjJ7uLbv
Y9dBd5XRuEmlJx3LTDx9+7bRo5i1QQKChzYmVA7B4CdMl5FzljC95jbR54LV5r6o
ZKdnH1W1sVCIwBsEhLRoOfaipJDEkmfRcxxEiNwa0+Rsw+yCfMZSdxyAWgcFNiOG
6pImcI1L4Jsjaz/iekiU9WA1YwFUQmneREYcPfvwixKJLNoPFSpuLOMWVJRX/vSx
fw93KzWK99vL341XZj6GK7VgrX3IujAUikSIzJLKne5OI0j6Lu67gaHTHCWxEXEb
OWIKmPR6qYAeRxQYKhrnVzj5TLlNT4rHhbCVqI/p49Ty71zNXe/adxEUCZaTYsWl
kEsCr21X5cyYkyQHKEBm2wtuV2nikHEd3QR11Lt/HZpC5inpTTouJGvpMkZ6yWvi
Z7zNwuZZd87X/GmTdTYHNezFTfGnGxsNefiOcTft63rtsnKeUdqVRWlcljarRa/1
PCpaLflYLYxcymb7psrUZBeljPsRjvqbR21SecahRAwjo7gDWunWqn6xaVn/vWZX
xVe5Fb9cbWmL42p/xYMRTZ++ir1qVyKGmjTtHjZvEFE2frgNvXobxIJsEPLok1UX
67pqxzIaLM4Zpn4klqTsASK+G3pZ/RBaZknAUbUQMNNQO4Lr++5TqLdMrKddqRwL
E+Eb5eMkB+tLfPEMQNzsZFdqVRF1p+46ixhK4oikOfLj/UHRv6YsGJNaF4FG7E8P
wj+9mqMOdQ2ipPsr8kmp/1tGecHD/9qpjURI1xrvkQM7/+RhiQJxL7xPNxk5u6Ve
M+TH8KDign3M5J5XAk7Pzu1YJVHNliab+JScDcPH8gCyoMJ1EUOd/BUHy7fQrVbZ
R2e4fAeMjHiKD/dDqM0zjTC5mQ9QZijhxlP7uoLWkGBK8aory1TC5gddA2uHgHGu
UphotCgKZX0urNx6wxY6EhzWgOn0B7mf2wclivuU0sU8nE0OHLqpx/w+fJ9+ihrl
raVNVMrwci7JiT8e2AYWyC07yERK2SVbVndnrY8EjXL4wzgLWSS4MM++VEsS2O2U
qa4ETNktQmOiBlaWObTTYAaa/o+VC8j58xFYNFvT9V+f98+6p3V3eIHSxvhGQmqu
40f9QnzLYTSEagzz+HpqoJzayOge60aBnV1GF6AQmxCkbq1Odn9K4ZFA4E44jgbC
nkEHIYjE/4qjgA6dZ1o9XdMbL5xWkBpF3medZtbIEe+KKi1PbKpdCiErqsVPNylw
WCdt2Uh/Ay/tIwyj4z1o1fRfHqB5Rm28DBoewvfWGg+XvESpaVL7INzW7+CuRVsF
jNmIRA1g+lTKvmJ1AAL2cTnhFAH+cnKHgXPqOUHKy4L5xesQ4h8T55sD2zaI2ayi
PUd1I33cOpjf7QvZlkSPPvoYe6bi2ZA3JQF2J3hKQtHhS7ADadk1s1vk36SUexNZ
C9eohzgibz0wrlX2JIEgvifRC5CilWYx0vke1BQaFMVGD7cyQsX9Ko600KBTMqL4
/6CtFS59D8WWksbHME0DV3ZLad5CF9svMSrKTz/VobB7p4hDnEzzJWc4uUK+BI16
GurYTRf15BI0VIdc5SlnFeAfoyu57gRPy5kYeFMq7Vap8Uyb+fKQc/nvAtGetKZ9
q2t0cSYdpyqcEBG0VDTSVCL6sEDCleGwODOrG5zZH7UVdfChvpa/FBmbairw9xWt
1BvMXh9vq5xw4TorkFLWS6mHaZNaQ6UfvR5mmyMeufPuut35J6he8eEslLkHBlSa
RKhT5ID8PQ8hwLps21HYO7s6TGFb/GnqT8U9+fA5Q+icabwmHtvQbIhXfx3dRd23
jFm8zkubEEO1X6fQ1o3+aJ2lgpz33YfPVAkeuEDoWouyUJh8KRp0KH9JscOVV30W
uVMxB1C9ARr58Q3QPh2STW1hfB13WuS/UrAKtqS9Jc3UieKuF+jbq27fsVp8T4Dg
umO9M4xhwkUGGdBT4tkcwKgYqODl1p+p0HSD2X0uaI+4Wa7NvWLb4SuFkyy9GJXe
EqXFlNSGScxpuoWFwQya6S9AhBLmJqcPyWQofE22IrWrhZQc7msLFdrBljQT5cA2
tr2sXtQYrANWRI3BVgK9zN/Mmxk8UslvZoLtMhjH1g+/aNcnc8hEicLhEfon5eGQ
psQ2nvOaBYh0KAc9LHFPFXzGqGA7HDBS1A2HwtQkeZQzUuHDF4OxhsWk5dYIY0Lo
S/q27qQ1Ycr1lYpBy5pvLuX1VHMIOmQY3/Fe6nAZwBMaCOdnOJo1GMGb/2sJk3jl
iBlRpA5hbT3tg5AOg63Ob1KTlQEfW51KWrVG5UAF1vqmdpHnTMFrfQJEe9rBu+MQ
351Un0TtFXP/o7pyw90ez0w/ad8xrIAplKgDFzyWeilF6hYM6HIEQosDX5JPmAQW
DNmnFVa9TPL3FB5mb1IHnmSIWHsqBW0APN3J8sKsSHl/qQ9YqRmDDWU/MBQsppAh
z0KvzjjNsYBftEqIOE+i5HD+Iyk9zthEDVwGCoHgAx7XbWB48SdyHxvrlKQcO+9q
gJs6t4MnxdibsllSyIN70KgwzIE5pLBxuNVHvnqt4NqLQ6INuE9kV89ot6Jqs7SD
Ni1nZeECxTsY+umaGqGQHUt0TM+qhz1KgOWj+Dsj43vSQsjFcPcvQGHNg9vMTF5K
nYaAZE5TNzl0iCWzJQZ0MAqJb5o/D2VMVhZOvdsEk7SwJsZU4abro0thtGDxn9dU
1+Ed2ML47iMkd3znmviBgCUKp9eXgua7P+DLkh4xmXVEhWovlO13LcrPpKKzCQPm
pXCnsf+FrVGuHLauyzhdoJVg/8VN0xCB88+qXDN+g87CDtH4Y/5zCSIKDXuIyPSD
WmYxZvrh1+1MViZi8ZGpNJMyNfKnv6kdUsBPzSODmdYgwTVVTTS+0N4KJwOX5qhP
2Thd8HR6SVdWvUqF9R7PVq2BMwEii4gVyrzDosWW6Vaby+d/TW84KsDWbmN9P3p8
uP1t2W+3hqEP1VMAJP2LhyqofAYfuHrAzznXrHOX1OBxV+0r5xfjy95BV+n4CbY+
WTencOq1jV9t6lYkPOpjsNrJv4n9V2XZzzrFeTe1jbGNRX49bKbYNLzfsr8SB7DD
2SCz3P5iCCa2bzTUND61N4Hpcu6qHBLXwZ1Bl9a4/8f24KSckXlgT/qVA3kA8oOR
2F7bJTFnK9XaVemiSWsDxEunNPzTDo3+jWtJoBnJPKiOWEo4hIcZFQO5qMfgUVMI
j9ICOgTj09e6cwKszDEI3oIIqAFQHGrB76vRkA1dL0ViqRb4nZ8jvKSTgaUOUXtt
qNaccGyN4sR33x4sL+K4b4gcV6UVhrf9lRK6OrjMqyr0WbsWC0sglMuycSY1J9A6
SZ6vkorhW+AvZKHXeujlWViIyL7RnEyzsrymA4+Ea7jggE6cxn8TuAKD6TCHMQGY
Jz2QI2m+Pjsrhh+OGR0rwbhVQ+CJ0aTF46W7KPS03Sn0wPP55d7H6miSClBKpduZ
tGEkS5aGdeWdgRNDqCc5y79Zgh83XKP0yvgkBySRSddmoZxX8qiBR/qLur0/+1Fn
SDCH+zGmjoMM02hT51Nbps9W5y7FqIQ6gJ/nk+iGSOciWXA7GvqnOmhstrBIuGQ4
awVfinbjS1ViaUOnHMDQ1ZCHDf2j8D5tN7ioR5kD5THH0LVUPu6SW7GdeoBe2MG6
+u1sCe2PjWyKGtheftbWrTTFa80xU+4erMaSwqrUyFwwXc9DCacu85l6wlzDVzFy
oMVpmaQv5fcUDE09x5tiXpNYia0jZJz/QZ4t6Ti6EUgTywk4UK2uKcauGi4VxAew
7V7quHclC+sXCb4ShzQ0QKwGfDU37tb0iQraDH1nYTmtBOA5BOJgUqPA0Bgge//A
rLtU9RFcAw1IGsk8HFQld5RJ3MBxFbsg2pA6humAaQ3KtZOxz6mSCxxRMfiagWQq
axzxHt9gp3azXFVZnzySWgy8rzgMcFR8irZMZhx8Pb/J0iIpk4z7aFtLfNpditS0
6bykdl0ZRDnuXuEZmDW49AFvAvHWy+LplO/a8GfXfR1iFGrZUFNP1W6U/AOhLWuy
JsZI/WV7ytI3ruyA6XG3Z+lSqfXCrt82/vH8IMMWPxej9Bp2Tww1lrGE2MCTxOim
ynX3Mq3hG2bxIbjChkPyP0CqJpdDlJqsC+WWp1O77BYaCoRjul6h0d0XO2ESjYut
EHiyhr9fx9bwGULuucIIBXaU3BCCaLszkujIsNRpg7Gp9mUYB8eeSwDp4lim+qAB
spuLlHA2Uqe8Jy+F0LEihZh+R33Se6xyFN5Rn2pAoHxR/Mtwicb1EQn8/Nx3pckV
9cwQ1gL890xr/YODfbyQnLCIisz9RH/nHa6KEUINCjjetLKqyrAbK/UKey9aydik
NlBvbL52xwDVBV6IOagUcq9DA1DrF7Ff3oZpM0KScVIEqSvIqVds7MqvhA0Dco5b
xRykyOrPhy51QqVahu4Vxs5WTVNmTLpxSuVv84jhmXa/SCiR9eqRhGPeV4f6+Ay5
FWL7VIg5Vrvy4Xs2G2p1Zjrmf85hb6axqF10ErFbXfH4j2HWqfM0nK3ccBS5xJXs
lAxWBM/zdrnYlHQ5KKRrNfWbHFdhwnuWnNZcuLvjy2FpbuckoFeSxAusVT+iyAia
8GIQO2ksdXnT7Xe65NpbHZH1rBaITgZBVBEniHzuw3tLgLBnmV2tcwWPKiSQAWEM
YnoYzk6lDYi3aJ+jOxK+m9f7rKHIcCCGwIgIYTrVMIEkHZbzBJ8r8yXvTITmBSft
9MEHM+aUzsDFCHWZcsCOi6fnI5FXOXOl2KBN2xVhB5+QeVzywOWrONMbj3uVS0D4
/DRMXxz7XNtAxRr5On9dMFaa4O+WRbwLSBlQJJlH5rKJuJoSkru7u14nT4FzaYnn
Iuf6ACiMKRCKvyXThM9Zqj2OvOu7+fdJOUOyBbQ45RJ/lx76B0E3PDIdTx7EbiuE
udfwwWr1UPUvx1zxuX/9F2HaxJ2/VMmH5ZyWxuoY4x1iAkZUoq+1FjKvPYjNpA4o
rQKZVAnk9hwAbFux1P2Nl1VT0EAQQ8jM9lNvXmIch4GaBQf2KKA400/G2W1InARy
iFquM5uUvVaGaCbd/3rohNNWBft376egzTvpg3OJ615OBjVEo01xZQ+77Hrb6e/H
1E0IZF0SCON6NyNUICj7KZYKx5FQ1zMhZiST4aOicpNWDYasYozmdULaQfrVraf6
kZx0JEjvlBT53s46l56UClFBIVZmWvQ50bbdL2iFBb74vETK2NFYj4Lx3ilOvaTE
cSyF40waVlc2YfF10DwT6nz0miH1x5c+uAkUGnpk4Th+cXN5sOHdQN4dUyovGL7m
/jsR+DyhItnk+897X3oCQkTWY8zS6Ea/Od3pxkqGKyj3S2qcX5jkiMIWGNQ/enKp
aPIK11Wn5JmdVcHcWmTCU3mDIn8RjFy3uyEPiSfWBQGO3Qo6wUHjdHo1mTXj91Zi
GLGclPMugfTg0mMQN6s+ZTHU2FTY56Thfy6cO3/MWSxpftnQviVAD8rOXvhpEidg
RIKdfVCVrRH6gEDab8OXORbqQgeZPObGKV8HrX+BUz9/LgnLL5zUxjmVq5xtqw10
z+EiclDXKp/UxmvM0E5ere5pQr2B8m9/bBNTaFC5iqgMwHyqsTmfT03+iM0iFIuU
+PLUMtDfUqvz5NNKs/hjN/+LYSyOFKE3eJPxA03BgMrkzaVHYhvrwV6btyMywEQN
k+FMiCxPKK4EMuhP4OCxSi326ypUMXTMgG4FD/hNjofhVKOUYGHYMcy4j11P4V8r
8v1ukuJi28qiNWFh5GMqb8tL3HkqwXY7TO+0kHuOg9ebkAzIG8v0RtPe+XQlVjUs
oBhIiNfJZWIH4dGuCwq7ozNq5DK17Pl1aZE6nff7sGKWBxJyMvSrN7uahKXo9lTx
IenhIahD+vF6WC9pUcsNNP3Ay44zE9LlH4bTxkoopcdwz1EUBkCyT65Oytj4LnSD
13XM/vsSoKLPOJI5puJCduKqwxiHjgtM6aFRifq+dD9wmoDIq6IFLotIA4B6BUu3
5yi2MjpiRDuYqvJ3W/WJhezZGpMn3A/IXTQc8493ellHKtYWtC9ikV04GUz6cnVQ
8tHJftP6L1EkGj+wq1vDs1LLsiPNB80hDvcM5xYZxR/ZnfxgMujkrJk8xH5afd4V
lWoXzpvs+GeZOJ1kJXuB1+Yl9oWT893HVCj1PpNACODyeJTeShGcEiOwH7lA3uCP
1yR3TFNdhF0djbbOgXhZvSHmS7UyvOMd5kD5tSno/acQOoENNYPAttM1VxGYrqlH
zUvIH3hrzyq0iqJ+AxSeMIJxz79ME96Ql1+GvHnNem/fqSxHkyHDHi6f03mWM3kf
OFGdS/EUki0bzW7PqekXGBubh7Ra2PZVkmKMjO0QMUSUclAhoZ1d0T2Lers0ZPG4
oaJ6B01mLpUd/ZHj7qt/p9O4D4MV2KpHR4iWFusHIqQJS6FbEbs3EpIX7KNWqgqU
tMTEfL7gkxZXU5QQIbOR9mi028qcUgJagjzJWE77sdi4GRCgOSjVk//eIdk5VIGC
rTUPYLa6wwYPTCg/G95VPapxWhhNonfTWW9wO8TBWKZH9S9pjbi8MTemuwBdWauG
Nn1epBscAG69WU4yYZVbzWA5V01ow8+KkLgTetiQEFS3xDVjMcPUqmIM4IXlaFmX
Zb/ej3YMcAI0jatP/1Uk5vazbEvBKwBxkEG0Rc22ST7NEuOBT8Ol3y9eJhwzm17o
APcP08nC+xXDtc98T9wsETRmkgcEvFJgoYFnmZXUCK7aj1WWQuIt3znWBxcF2ih/
Ggv8k5cS1osqisB7cDYrPLSu1o894IpUiZTeXvrSQAr/PORbU7B/CGIz9wH0V/0+
F779E6OMOkiyo2MOEvtmiH5L1ory7KNfG9L1RUXMxzTCDWQQWIsYmJLU46znTk3r
BO8LhJjA9nOA1LFqc+3IEMgQEi9gxa/qKY4ElrdelSAO/T9znd1vHjnnNedeN7ji
yJWR8ZOunCjpYFBCQOiFIr4Jf14mhkEHkXyHfG/d2MW3NsAy+1NaQ51/YdzgpZPv
cTXhLWORS9nVwyEnuEjzO8MRYEVLcjtPk6LURm7CXAArrBcpSDxQ9+2Kup3aS9f5
+U8YePo5z9wcdKs5hOij+/C6kwHDP3LMKkthBkeYgM1BhJZ108gyIUO4Lp77naR4
VREgFawbm8nFEZvcnQa3y+zuwr0YZtLjJyRUfbQNlTQJW8/cGcNgNiaXUPGqoW2f
oMa04NQvar/jcU9c/+VOmbWwB3NIEqchALRyStbvyBops26mAGKrSrupoqzd8D6l
mJ3AbPeWfgwYAYrdrixU5zmIYxAU1dFdvlXxnQeGm/DF/Resu4/5s8Lrr0eokTV6
5O9JRTCr2uq09i9YPfZFG6QnSi+HqAUqY2C76lw2FNlW3tmnMqPVSgEZBt4mBHqX
d15dCuztiRbPbBtLkAlrSal82ZJkfHrUYoZRqSYTcUtlICjEJRmxY54JUDZV2hWc
z3AMo/hvVL41pPwCQ095lAIa+alAdPWPbOO6j+/Yn49xWtWK/slsxtrtC2Abcdq2
7DKYeV/PemWgIEMLh2eIYbCwuAwX2iew88aDq97LzWn4Kat4oPYjxRzNoRgt8Vk+
D/4XJKRVPBMjizCOBbGZ+IukhWYokcZA7igOifcNU0E+WcenKJBgLFkdBNJMpQDi
AvaQO0C4Av0P47uWvNihxjKJzXIaYX5jM6zxYDyHHk5DZmiMIMDcxE6Ts2oR4wyh
v6nWRmqnBgmIZUXa0AycO+YJMqvKRfKyBVgzpIbOzhLRhSkqh7p1tfIpBvcmVZaX
O2jO1S3tDzlQYkvSbskxSR+5H6AhtTDrEPrGeho705eqOK8UCNIJO1qatmw3SAZc
HlyPrHfhUlzZg8yvRJPFrjCnu8DZBhGcO1Ki8Hj5GFtl+hYKAjF+ZkwQcFGgiOIu
67zy0p3hXelHWKzhQQHLmQ9pfUOtsm6bD1mi1FTU72x2ARTyjvGhwKoypDSdAMF3
tH9OuCjyx1JempvopRPe7FcUzxsQ1isoU8NLeNzFdtl5keBVEkHIAj//Be6FYvAp
1cCaEFrvnVl9wlJGHP6Ja1/tdfYm1wfvbgbJMfjBWn5jfxxo9G5Gfqkeazu/XYxd
FP0eofEBawtPvKCA12BIlEY419+oPqIvyIodMVBiiAZK30WLO1da7++o0t7c+8Ua
c5IZ+Qq3yr3LFjP+ZiQtZKyklrmizU4JJ8Qi0wvOxAs6TNaiSiOQGMNFYn9FTGsx
gNzgjaRNdDowDEuv2Gd0QNluozrduWMAyhjxYYiEDLtBBlioacyWFEPdVsUKg+Yz
XGjt3E552uhfUGQPkr5MeJsBvmA7zfwKNt6XELXYjjKMzU+potEpsmtf6aC0WSh3
Dr9zMDn+UpKPy3eTaUEPMZueYwseArYQpAh7LFqarW70x/aw2d/RdLCtRFy89crE
k1jDQBoluBn24R+VDG3wKED4dJ/k85vfhXGIF1nswJ6UHuP7l/d77vdvRY/K3Zp6
XtAiSFLnyBf4Wa3v4O4wBcTGO6LMmFg2kK/FyAOg7zaUS7Zsk8Pbu+S0Q7PEa6QK
NjgGij2Eej/X1cIN0E6RC1SRvkUbVCGvlvg1ZCSmFJQLrK141tlChCFsuacdJ1SU
OxRs+eOcmhBoXB31/x5u7gMh7011HV7tOi4zt9OHg7S8IFutPr0vkIBqSUSRfFHU
8eIyeKds5E0yw8ZyZhtfoUbaodjCHWsw8qOyVMcektQGWUD13Q+TIwbnmticCgUR
rh0b0I6pjoXE7GY8oR7DLNJk33Nj77TXcpBm8eqUT4beAviLr8MttIWDLB5/fj5V
HJi0M5rK90qeoQ5X9Vm7xmNWPEamgdYPfeo0TpznpXYU+rDCvGbHbiudlBp6WDB0
epA+A0nQzmU+kju8J8EpVNNLW7J46jE/WktdEg+dKz9dz1ks6N+g7ys4nxUb5eM1
nYY1LONTbbUOpWUcA+zq4eWBme9+A1kDVazPsvOSeUU02jjauQ0GbfmbLco0hdms
mAnvfK4cIsNq62vtKvZ+xPfJDOCNqYEXpQHF4szVclM8M8ZbCe6ByQ7ia8rr7Nij
g9vZBvmSvjDQMO1tviTuGJXTzZu5BkBu00/Byi6fttGod8o56EeHNdZMdoXRWlpX
uUOGLJvrBCSnODAxubaTxXsaxVfp+CjgsBB/GEJfmdFw1N6d4GAeMV8JJU3OffBw
XmphYC8wvOC5ejRyInWTpiGs58LAcyXRmzde8EHwhdLtul2xGUCAPpEeAE1DrhPP
IRgvx+hN2nycyOhS5ed1yDrAiH2+gSJS1zNNG76KhtxvU9TvrSXCRJcfMBcaG3QC
+Wm7o5TLfX5ITks5SshMr0gwUOsWokDxXU+O+XeCwMwOk/aN8VKxk90abNww5xk4
5clsxxvvt3x7LCpd+46pAMqVucpLc7/qaFfaTGM6FQwPjJdrG3i90ropRo1pMFWP
cqScmtDrE09Jfim0J5SbpoORj891n7jmf2dFmXzdv79EMGbgZgkbTvw7L+JGWDRM
x3QsG50RTm4sp0uzvMy1FbCxQtcMX+NjuKAierxjAbJyinp1wGOwbfK74ZWq2rzA
Lp2Qh+uYUlGz9egFgd9snpt1RPflOcdV+FcQ8vZXh5oMtAq0a37t3zRw5dUASBiV
Bq1WGvNP/bbDD7ErZ4q6mSjk6Q+d91fbpW2R4w7yRq2dGfgmTZQ0xKDPNy2VOceO
I8gDjxj8JoryzuTPztb4aJnZGYG3YurvB17BY77mpBZlwHMJcEtnMacSqZxpV2SS
iee3YQVk70QurvyxTUi46frbKiMK2yRZtbZTiajsj6WCZZ35cJk3py0EvvFtBb9C
2g+WBCGG8PtHIeRLK/Ihp1SsCGNHLB6nAT5YL8VpIrewQmsQG9nXm6G8we3I+cHU
45eLRgiHd7nMuienwdHs5fWEA+WkluB0VkhPNlnVjY980VsfiCH8Rxvuok9p2dPb
bR4CGEiAwRgjnB7K9sRAtWjbj3RXf1O16JtcKaGVjRX49bKfEmicmYwv3ZEBTm0z
5KDL83BNc2V/9dNqy7EtSNsPrlP7NwDODc6nUBdJov+bMMSH9UqHYROojKKOZHkA
c1dtq2I+H6zjNjsKO1UnAABMFZRpubfWhnC4vzIzmNUfzmqHgBU7EocFoROYrzhL
NXv8HV2JeNl2qC0wtetlyZTfQLqhY/S1maW8+AXgR6l69aNyocQfLhRb1SA1yZr2
lcw7zZyoRpJa9POi3jkiR0eUZBrdYgS5FO8SPCiXbQqaNM2HL8viuiemFZR/aoIA
ZuANFSOwbHFeTLuOu29DDTDoZqgP6SxBTHBCcTH0e4AKjZid5Z6M+sDNDTkewTTW
5pW/uRiQCFQL9YiswMAZiJMdNyFt1/N6OwHo143JQqzjaQAQcKne8XQ3k1vA50t2
AzVLSoftn4yCbruuI9ZkxjhXz6PWdC7aaoMNdLvWibYMRj+RaCqHh3d+0HqvE+q1
katayEx72vdag9u0fC4hLeUEuFyCc2Wd3xBqURkkRUIaOkX2tsG0CNf1bzmoy0G3
fCG6qO+nus1uG5mVWtnBYTAs4GisdAEjc+ZVppqeeWI1NiZ3ukrloxv5kz/zLpsB
jlMRbf2ylwBroP+q9X9UINWB1Av50okmSgpnPBbFipXdESmDzcXxVOV+X7RGfinA
69fQs5MIOjXYzBXaps6QNKnwEI5GTIg2AM1YjMPZCMMKQ54PgPr8rLX7s2Pq494S
t7SVIEFOUFdqlhgl87IX6Wyrsp1KxE1gtBD9BJkxM/xiZJMMHZwoCPyj/Iyy8FPq
OHKVu4hGV6PeJq+4nFZ0vPeGUF0btuSZlcThIqI2zyQWFgdOrjfqVWv3werx6RYE
BB/9fZRmVFrQWpDE89LmSAJGZyDRrhkuJ+SQqawPNod8KOmFXtobZr50iZ164+Fx
/kzBR1dusz6QKUN4/jOrXRtxT5egixUPvkF8907+FgWGnPIGxDXLyQXEi6HwPN6/
rLP8gp7greq9PvxYbVx82z0WzSben4wpc+2SrFJd+Ql+R+qYV+khuVB5P2dFBldT
mt35rMtFgqVU41FCNoIwgiiz+C5CR6GpKQBNT3Ikd0IEeCBpzxcDabWmMCOujpwu
WnSSXE8xxkE9TBAMqD3sHk8NgGQlEPCo8vnovzrV5S/FlIK1ds4DnUA37MUQg4SD
pbD8c+cdxNJKBEx1t1FURTec1Ssw4+tiV6b7uYidhxPgiZ2z+vknH6M2tVsyTlEo
a/+Sid0L0gUKFTqx14uAK2D8cfqqGZxRVDJNB9kNOuXKn1J0d96ZsQgt8cbXLheo
L6eNZmJpTKgaIzBmnsBU+vIz/zXl/tcqNTCFT7efL14gZFnHfQTRawhEVfjrBbFe
WM/8Acercbn8hBxkpJU9Uwzsr7sHkXQLKyeVlhs//xeodm7uHG7Xvpv4WHI/vxwP
h2e0/luyyNQ/g6nzh0oLTsPmdbQie7xNTrxXHdvq6WrDPtxdcAbDIt0RUannE2fB
i9/TARUw1EsAUGktSUT2L0aUAq0o5joSNyO+v0RWDGM0w5IxLmHXEmKJ9XLBvYMg
oab4xo8+zpfR13bQ8L9l5HmKXGphKrWab4s/PKJky7Iv9snqaSS0rR4oQLYDivvw
4keRN0MVA9isRCofgMJBABX74A4sip1I1SKlxzXnNxwjH0qCoSvYSMT5vhlvKR6G
+qtPGKMMBpxd/QjZAdTHO6LHs03Ko75UAXqnGh/1uavjTg0DBclQqqFuCy0MpTLp
hNr7q/yYbxlL0NpP6xVyoFOGrKSzwMsSuWHWT1+wsFyUVm/TahGqYFSLO8TFDEPa
oVOtiWAdOT0Pf9m6cM0HR6TeU/I8ESIjUdVEEW0FNokrzP94szlI3aHT0bKocyWu
re6U6p+Kn77wIyeBeRDK98HeCnuDPYw7qEia5SqNdgZFpAQo9+Hobf2s9xNNC0xU
N6AHfMZPSoc2U5HMIeWF+7t37ySLZTlOihLQfVlHkN2w9CNIQcYcmpExHPmC1BRS
cIBEdrzN2sTvaiMMB+/C7c8n7Vwp0QzukOj9BRwqEYCmSZg9kBOyD3AUdtq+iVdJ
Y2mqqvBbCSAXwy94zKqVIkUviisR5RwPs2MEL/ul2ULuG6/CZkqrH2D5u0Kwm8zj
qNAzs52aM4AEsEmxCX3mdFne33vMuIUkImZysWEog7B5S+9tEDIwu32C1mHG6JuV
Xf80j2YeskUbxGRNJT+IfM9H6ONCB0lYNoxdtoAxd1BKS8HhYUPm2nwrcJCrK3cr
BAvfmeqoa/aeEb7s4WRwkBHbCn9dO67LRfLUMOu7MfJv+OjloF788Mjb1KIS1BQc
yHjeIO9nNSXKm0OW/kpDvk0t4D6g3qvmFJgarrvC40wVkqXvjdpAi6y1ZN/EYFmO
5P/IsQRQQkoAxri2mmN1PuqY7OZiZICzYI45U5gcGCBMmAMSfSqajr0I6MjfFR3C
I6ovTrSIFW6I/gGIGHp6YvCZZeLG7WAZmFgwL8Ger+YwAoNsIv/ABR7rkeXA669h
v21FGsnNFUJ+gu6lfBo79xWnSTK5xa7IvG34Mpdrd4HrKMWJst2ql2P1ca1qrQcG
Yp6pfVauEx51P7uK4jDZD//8PhUDB3hrhyZrXYCXu0aEsVNfoBoNIhy3V98Hrd3+
7D769UW06yBNbPz21uvr/mQ5fpkyLvnTs3StfCviuQv7188WvBMHlrXHWDgRTcAr
CMKpcGs2C3qWiZ7ADcVAymGA8rph3OAEzHvr/Q/QYPvX5lEaTJGxLJ7/JUlTNvWh
8tWhUAOWod++/uflZMncxeHzap0KKNPknsMCTLSxPz/fMN6kUzkVqU8CKZqYLKsh
iNWreTxjC3OSWIWlLrw/svAy0wTJrOT8tNDhkaAfdgbo924illcoO3FEJbmJJzak
UAt9HFEueQDoDovEH1gsPe+1USthGUVtR1mT+XrAqjEKJP81/VzeVvgfcv3qGwTc
xSoWENOYvZw2sLiXidyg+MOJZzxtNmCsB796YO2uI7P8kl1RZmeaKNOClJnM0pqZ
KGiTvnCWPT2Hcl3wvp6OXleZlq27jJPdX7NXa6kF9Lro7QNzNJueV/wMsnJxhikP
horc4W+6uM77U/wJ1U0xDaPtN8uZCNx/FRfT0fUCwnpUav0X3zGH2mQ5VTz6iFNm
28CMyT4HaXxjREMQhebCpU7cOe84qbc/KaAjxOozqzO+9d5cIb8P+pnbJUJDLTp/
yEJJN5fHfRwX8K8BTcawNuU2/BpcUSSAEy5YVM68DtzpSqgSTmU8p1hIqDbmLVrH
IcPDYVAuET2pdU8I147Alap+9mcseQwHKSKV23GrKru3YKtjGBaBmS47BKICCiN5
QobdjFH37LXf6Iq35hwbBpi3gNaVJp8CGsHggl1aN/s4kEwf+MrNm0EeYollPCxm
hp5FWRPTijSVcXDBlMtz6PZkO2kGqmUu6ZXVWyXy6pq7/fuB7tSF0d+ahHJP7A41
AyQWT/hojfWlhfp9Nwc8BAtOtXgrGVw5DTcgXy8gMmpZ5NxgW68h6x/ShPleofnf
0OkGdrY0gLGP+oF/xN0+XE+GjCxM4UEv4xnq6vy1iylB2g67pgwvzVHUXgqHZdie
an8Z5rUqECNB6LyjwFDn5K3PKHdisyBqCHxvkcTElsGfsM2xOa1Msd9dC6HdSsmf
cmpGfCSu+UzozNK5wjTvJzTla84Sjn+4KNObQ0xOC8oxLf+bTG0qJAm6RdofkydJ
qH01Y9BZLZNs8IA686B4iUeGvodL480i/aS763yZa6cJTk4WSIMynlRYgHKFihqK
/RO1G1LxhPlfzGUf2hls3lxzVaZoHXQcf13+otXMy+cUhCnGoN3lX4+N+xt+Gscq
3SkKRce9vauebrZorTJZCjcbAUn3J0lRWBssCQeXkE9h3BLD0Ki2cozJszQ9J/jU
ez9poiWwtB5VscKoSSASS3cnPn9bwgvL2LuuJQ1W9p8eVXcQNnHpaKxKO1WrR3jc
hg+RGssp3aAUsT1FDVdbRax5Qz0pEZY3TsATFBZn4YznVYv0Hij32pWfwUd7/i/5
3Fs3tkAOevanBBJz9RzwMsT+uPBWSa6ZkBKx8i/atq7tRPzzLjd5AoWOceT6OLlT
yjv87BJXDQq7fJQYa/1DvVE9bZByVvX/v9BHsn0ewW5Z/C3xDa/V2hSiKXgnMGEE
ezuGTNIg30WdrntuNGm+uDEmEZt2hdbmST9c8J9tiwQ/RmNUQ6fo954MVZbnh0Yj
36oUiZb0+sVm5QiEAySbGWEn26fzz0kOcWS3FN3CwVIAaDiIXRJUjsLz28S882hb
3oQqH5gPcQE97bYlDar4417x47uQ7hWIN5XpMrcw8G8N5zHkK6xb1YgNN3mWqi8Q
3UGSbMy4XOl0VXbaiCLchGDWE7vgdKTFSmPyFwmTO6yfAzQWehMTeTCdYtYEVL+B
A4WL6giKG/HWpMcf4xFRFNH3UkppX4W/SyjUFbf/9oAFlYeB8tDb7Vno79/5HLVn
PbcVzrANYf/ahvTeiHnhksvlB9GlhVyWOq2Tx+hYfr/wcwTS1cjFCgxDBl+F32Kw
Po30x+Ln81U1g1czUBaQY+W84PyeyGaEJW9lSzdV2D+KqeSfZfiXK6uO2TxcvU58
pLVO0HBMLGVtahN/CB4LuOFf0v1fz0bNr2ZstKTSuHC8YuuIs61i9R8cSSEVZq6F
5vz6YEWw1n+OB3amsZJX6FxyCcLaRVdeUe77s/KT1tycgvOYpI9TZOze1eSb1Cc8
1H+hG7bkpOx4mt42b567nuBEHtGLuND/4CklPVD7WSc+sW/t86tuO701kVLh8llA
I29fCojFt5ZrAXf1Y+1GAoXRGN9Bjr/NcDpgV/k5qbROmuJgAdipk/pU2lL8VSxk
rUuVDaZvRNusY7IquJzrsl1C9GWI0DaCR5CSpvnPOtm7Tp8SiPaC50l++RZXa7CM
QYBgEBOTRehiD6v2+NahOeKiWwkz5mo5j8cxjbHQzMyvh1RzOox1o5ofX5Kn/LyO
IAyM1gh+IXWhQXM417dfF9FMHIChu9uFKxAz6g0RkydEMMrJ/x3okseUVHOXNI0V
CGO8HFKDtg5sCKrkKroq28XqYQGFIr0bM2/vUGgizvZibVB6VbwSnGHtRNFJfBuV
uc5bVBZo2oHwcJj0hdzBtn951qFCcpPfu/opWjxaDuI8PhM89u86AgkWB6JMQ46T
cDoskMs6bjsIkxBgwTPgtlAAjYb4Qnej1r/iC8RF/oGnO4awJGz6tupXcJi4yoNH
LaCxXRuvp8MowEdIFkt0DAyr01I7RgKCvAKEdygG1IPcwQAnTkK21wvX+/IjRHCj
Z4Jevh+W760a43x6NtBqhvH7uIfgRmjWbn6W4i1pMWFboYldEJh55WtrBgDEJHbH
5YVRTqSeL/qhLhTH7EiZez9Ui1+Vmx9gzgtPE601Wpxsv321BL8kQaHNDWNKdYep
oh8y4eg3n5jxiB+6zbge0HrrpPohp56PEjm0OgJvZ61TN6PDp6ypGK8/OqrbRQKU
PZXNeY4gLbHIWYdIUpa5zfs7XhP2OwiofPLJmGGCOtvu+6fsXht8xRwiW3mliEg6
MlC4RWFHNy9mqHWOS0a/WUZ3/zH4gJqjVLAr7pEzKDak1/jUePZzmM6+QoZ5u66l
DYTBhQCm1LDcC5k7ucKfwVYrDR2/HKLoi3dh7eBcpwQ8tkP8Qz9oU4zzDsDpTsYK
9Su80ji5sBmuSnFNDVw2Un88hRFsQEH9yusMAtacK+ouQ7x7ptoV2eW4iKawgPmO
7lVRal98cnUgQQwkwk8UOWYxkZRJ4xlMI+0IMrr8hqaKPU3G5HgWj5owLpu2TPSz
Hl3d+6AhJO1e4YJ5irMBTj3KyVcx5vP0Sq5+7URxJ0zN7Gcp5M7Ehgq6ElMu1TrN
o5TT4Nbl9AbPSuLApymE1iNryVLVyu1pyU/YDbGzGHU4G9TfCsxKcAmFdgnGJBjN
eDuX9ccnuZZNIBQxbOV7VKxonwSAC35hOda8qn4dPNLKXnsnKTqLJDxQeVmBnicL
ztQjZ9ZmheuCuDo6sai3A5haCldmKf3SMNofEuk/Fl90R//yHNt6fypER3Z2G70g
iknan3uouMNfofmoEBTyUlT1WWeK6qKrx8ZLna+jIYgw5nmyUzJdCCvUxqueMf1d
ZWQq0fhZJVHp0WkfQW68OXmhmdag+BG/toIK9KxNLjlEYKMQ4qNSNkNTKy9zQiex
YyPvIQDLhNIma3YbalLVaS/POg7BzVRus9WcAexf8UyOwfnYxyTX/gX290XNKPR6
Ju5ousTq4Z9wlgMGR5rubrvvvEmF1nRS0ByEhTFfc0zYSw3WkvgfYqZR4Vh7nUZ6
SaDsct22AGC4aA6iucIZEMJyg1K9dHjkymRQFLQwmBpNSXc6vSv8d4ZXeYbvjKuu
wI7QvcD43YPVL9X8aFRqdwi4uJqJZxs4J5zuFzqSYzJRCMoaBfGGOhUPesEmk1xc
yIST7PSpyTheO3bd/KyRViN25c0eoB74ZUs8Rb3NjV7cwqoZlBGPueol/uucKPG8
h2NYVkKLkGmucQZwZvD7tD+8fIGKoUzWFJVWC/6PXGdQV45XXsVZS0bW3a5ACwKP
77RqcLbjt0kpCH3DUdHetpJrNzc05S+gWlXBfssXXl59/Y01zfruW7MVqS6xYBTl
hWb0wnNgW6SWFISOJD//E2A0+r56vnLMpZPaiXeXRDAO+7LS4GrtA7mGee4LmEXW
rTFSN0cMbK41VvXHMFnPuoW1dqnu2TSCi1M6EL2G0MS70LIMHDipbwqiaGurSSET
sVDTTTo7i0skQNZdj6vywOL04s1NO320mtrk93RSY2VTpA2PNL0Rc63LHwwuascw
IwDvQZFoziYnwRASNLPsDfjA2clSegaIPPc+L7plr8rJgsLgxiMoyqnbjrAsPUxU
fB5DOqhrLZ1o8S4hc5q6W551JLuFxbyRMsN+JxPGEZ/A3ubuyPL+ij+pwGxqUdKz
90G68kRX0fc0tRY3kIR8iugAwOVSd2JjwMDR/aeusj8lneAGJH7b6vKCgxz8nekw
1HRl0b4BVLtkvn4YCUhk6MjlziF2Q9z5Du0mvuu4NBLPSwIe9X1Ql1Kkste580oZ
+lg68nU61g4dUQT44ta0w88fa7eeOR1qAOoWFmMjfz/snbd7OUzpfpZNDk8CLr5L
ZOR+o/wYBJm63UwAppRkuAp5V+vvOtrQt0nP5FxYdVcS26fCLofmo6+t1VjrxzKn
LAixk8WJyP9L8/gvK7B3leVvWYCSaK0kMHbf/LtkkPcQNXg0YFJXk55Mp7ZZ6x4X
Gus8RgkjUVE81gRqhv+rhUWy8Y0t/hZ/iVOiSymam2IVtVdt6SoINdVR+0te1jqM
+6oJ8vlr3s1nZRD77MgM1EYEZ5RDDgkZQDA59W7CrGlKrQ+FsLDxUUq9hk3WppiV
t7AKsl0HpuJz32CbFNxSUoGgygrNWtqjOInlF/nCfjiHKujs2sJltflBGxIbcbbQ
NNs7FjrFw/F+ZYen61DiaJ+qN8i49qDDLHM+7fzVwCWXtL0BJiy3DCke8AhV/oFz
r7CoIZLOPW1JP2ZCtgGPwItgfciT4ZborylvV3ErUm1UyFmlffzKCMq1BAXDZvBf
aFWcptrVwZ+otkFXVlZpvHvepbABzyejMMIMIFXwxbBM18JHa+ijYthIxN7Qe5Zt
NrUijfX9hr4SMzktl8YrE43jboLqHvSmkypolw4Ts6gSVfsKA5SvJX/DF9ceP6QK
D188KxVBt3MqvyG3yVTwcDW3dhkJeDlobI2W5qH/rvYLFezP52yrnEVHcYsARU7T
WZ/8a+lF0QkNBJUIdD/oW0A8bR4YngipbaOJxapRZCwnPo9izZ7ZNadWU+KdaTSz
Csu4a7Sx6xeN5jS+zhnOlv/rRNKQVp4t+pEJOG/DScowYd4yQlf51tLNZJjRM27w
JtDsRFmjIFH0d9gDieXEDzO6XU3m6FQEzRcPORjQv0stMXmJcnFpNXw6sl87WgsX
8138PmN44eBVL3316ApJF8u7Kz22uACsmdnURTq60q0FJOOUo7bqhf4qxtFpawC5
CgAb6sEDcZU4NBpkIuNfRrpDmSgcyeXVPKNFBPUhq7+TnOmRhXtsl3Ar4OlibsUM
j7JveIKp8c6pHshfnj8YsnWa7apbrZYPUVwQBniMQLNXedZbUFI/Ofavqa41S44J
jmMHixRzIHujSUoj/RQAl51UvvEpL4ufy1uvHa57+rQD6pVwQelZeTVgWb+pLf5K
AV6cSgLI8XAK9RbX2yiDzLENGme+KjYy4eLKZjBgh5ZhGPDBuDNStxYFTn0q+ctC
B7k+EERFbGPqpY2DbP7sUWV+0tqa/ToLBaK2sXdVtEywCBRVz2fYpdnYV30ewjmx
yFc4xeosxUaxiY+YEzExewWn7c/XjP3/qxaGEWfNqUgOYDTz7DXG7/MD2FN0YxDu
AWIXG9LI0XmaiIfD5DIxuh4EbkRuXZOeh5qhEpoIBZuoI9fdORGo5rBkapFXxBA4
+v1yNWdEcTMq09T8hpPDlZmmeid4hWx+UynqZps8nwiuxNOjsU9ElwmJSbCo0HIY
SCxgYSRSnJHE7/jppAd/KeOw/ggQbRRh9ylbXmYj28NDmvyoeJNPfm4mI2BFHgw5
P5NHWVKtYWhHeVnI2aVLlt6VPadej4NcKkX5sF7GcTF8V+z7ghsmQSbTKZYLtLCs
lfOr4ataReYX9wjaJHEQ+7uh5MTd15o3u3ycsmKycAGpq6rWstwVay33pbqpdZse
O4Gta4eernnQw3UYSX7AE6JCWFuq3BGaC5TshfR/cLqDPbMpZY2Cw8GKAVURsJhQ
VS5IXAtMNYAAQuCGLjA9zdhq8QyVjX+v4b6vMpBP+kgypgyajuXo5wGlkRYTRYaR
KSPZuCcvtMWFInWaOdMRk6XraFRCWQ1EM9TQ9bFWpJnay5FZiKcJS0JT4lrOlerc
Bh32fERo16CNdbVFAySYoNtVVHq6kmx57LHPZ7sGT7z4yu/bgENzJOcbXfxGeM6N
qk7nyA/7Ay6eiJwSsLB4B+WJFxTzt+c7iAhmW9Knr5rtJZ2rvT/NV8FmFWkMkuG1
ptQp7ftHc0YX0lyWajanQ63ux3hn27jAkKQNKJXXKL/GHj3E4f3eCTcwhsNINFlR
Od7dO2Nc4CWnFBGRssQaMOcuLuunPFIXK+UWJDFcHYFqYkh7Uk3jx7kbEcpJvQCp
R01+T7Es0qvFxAqihHWj4UOmsF9KPPzVbKi+QYkWVo2u/R2fpbab7Ww39+khee7e
o9QJM/+y9blI+QiqXjctxLlM5L8NJhBrWdxCkan30LRewPSgvi8yFZpd3aiyak7n
uSOiDHhPa46ZWwsaZ1t5uhiJ1OnihlA3e1BdEZrmbfwaP/6gIbgJgH8t7znOsVo2
i4CIYugmvSxDrh+lExrscDWsAoywy0M7TCFL5iersbIhGRrP1WE2aGcShGkItkVT
wjtFpMbREp/MwykUMN3OUdAEcVw/YsVsf4XciNXp7Cp0DeDpNR7o7fBpmFXGsSWz
sleNS87XCUdlqvB00A+NgyveFacyItEUZ7i8YfSSDjudn0OOGmPAnhNpylYrtMdI
3iWYdwqslWmZeHcwB75njIbw5MI+W16WzGP8NJacjMD95oanvmufBnaoewNvO7ok
O9XI8y+dPlNrZjgYXDZZ5xPG68KY5Ei8PbrwGodkJPVLng7aphlKSFBr76uSc91t
tiHR85rEddvcnhMkhn4WZShLE6R0ZaYDwERE3qI6rlLOUuHLRzfRep1JivVbJD5j
yuhvZP4JqH4TzM3Bgzdtcl1EP4+gDJ8hHnTdFYvjixKbLii24WEj9rC7q1cZbiTL
Qx9udI1J6CfEYTrQGNRqaIT7x1W0fg+wzwFLZOdv5MZcyOnBblqkODJULBd0AR+X
GlPPLfSghMnTvX6zzntQzi+DciVzJ1lGDajA/DUG6mWiiYCoTYlQMSxVVxQWgIr2
noBTaqPg2tpXyr7KJ4pxlPRCIL1+frYtaGdRIwtmLBW09LvggkNa7x9/FglDXrS5
qXTmqUKBFD6Ttp0KK1VY9zloH1Q1dufipoQUmngZRZed1/3CWzO2HvlrgA8bFOFS
kYGcvTKcMsNWF2o1z+MY4sAx0TK6+EEpmMhAZjrtJm+H7O1JhSFad2UBcFXJ1Uve
/FrOt52UjzRUnLIteM3xMu8HBWrcwz+9kTY+auHaKXuZZvZkRHaLdwnvouao8X4h
GtpwAh56GTGw8NXsq1uYiadWvguzL6o4+BA4LOQsqi2wE17Nqrjqqwf6yN2XbJ2r
pyZNUyLyR4QJrYWIfbtA/G5StW65WTAEeI9qcIG3HaKl95ZxzWIR7ePQ0xdS7Hy8
g1Mqc71jLZMrb2pBowYzyh8y1Kq8eNvP2bvgvZ7DRDSmETixzjEJViETFZD7SSWS
ZjOskbnwAs25NI3nK+8J1/af6w8KVmjiPlfFWw6Du32+Oq0yY0J+q4/hgjXxJXKW
oYQO1YszxC/K9ePKgndDLsqbQyZ1xfweXwZajT12yxO1oAnCTl7NICLSxz6oh5vS
UgRiEPthSlBwWdl/r3gDFmPQi57v0VvkSTBQlnJ7DE4l3X1fACzW2bJuMR+S2KmW
A+napz5AAfuw4/qOE0/gWKego62KncRQESM+sEPy8pt26CMER+XIG4uCY9Zni0p1
NLrdfUKiAOJJNet0Z9VmtA3KfsWCE2pztHYus4K9bs8/rZfmPQcHhXZi4ryf5QEV
8OfNkwjnyMBJINfyhFIIEtbpKNfndHBIApdShdxMCkzl9jTPiX6/aYjM6rLj1dWq
aEgsGJRPkW8e6JL3mawYUEbKqvHv1mhveHTOi0ANaOnxnpDnUDeD615mlgYDjYLn
kveJfYiDc9cLnKd1zJ+BvPzYqPA+xpIEP+SFzrEHF+Trq6TwI/wSvNkGWDQNj3sw
jNnlN5z1/2ZYxdm9uGVqaCsG3VD4MehytEb/8mpUGfc0AruS8aLrL1DWqsygN1Ob
PdeCxEFiY7nevi52lvtYXSlXHRrWH5a2vg4/nwdB9BnK0vLR5nVvFxMRM5+bInY3
cQRAN/56yBKSKcxcWOgL4cR/buvZFoUBh6FQsij6iXwdRQkeD59EQL7cQFUl6vXd
vXMpSrP1u4RdjoKLgUvnh2mvwhZWnjtO8xriB+yBdoLHMqwK8hx0pNOArGYDXHQw
5JW9QYOJyGFK2v1ig06WKYn0Rs+ETN5/TmHBjEZ0xiMJyNhJysS/GWkkO1wcNyB1
web1pqa5PvqpX/7oWh05fUpcI2enYAAAWpT87IIUVfpmSe2ZASEZbgHV8CNtUQ8G
kyMcpTD0S0lRaRvUZXsAXbhpwrDWG6RRDUipofT2+UMXDOS4NUIKRV+8dSGoLf/V
R9XYC9/USEb4rziw+o8mJP0LA572tlcgBO9R/lZaqRomQeKNh1tzdpVfp9c2OqBw
SVLrPVhjDcnJWmsKIRAZ2iSBuxS33jSl8qYCoMYvKfqJy4DL+wR+RdypTw9Fswx3
EDrxSGEa0AHwtxY3vWs5LHRmOn8IW/an+GSvGrjbtZfBe5O8koINm0rq/icopHKv
uwotnuhiwcC95QJwo7g8014xrx11stRxKdw5WuLXC2ih69IvLBBJJJpoqXmsoJ++
0mFNOmNyvYoN0OHMJoYVPgtfXfSxA9K1qsw4hB0DQNeZhazpgs76/iaV+/3qEfZb
lKRjIWTwxcBvluyR4+Jjjar4MtGelcVJzAGSCVYsP6NjmGes4iPecO2MU1ySvReQ
2U2o8eA09QLKy6Bv5yQSs0Yn+C6aAWYfcHKDs9eYxhOYaUfPJa/2ZKDxR6lGXzOi
HScgvPCmET6nmhXnD9rzIrrV5k3vSJQiUMZw6oohsRajgEwF0nwjyIC/YLdDZIJy
fImLBEr32ppCLpiYi9X5qk9WV69JCJCV2zmuLIcppamLt3tt0cwobPMW33QPqCdl
rq/rxKhGvwZLxLRt/sY9F0+US3fmYXoTJLuz/6guICugLuo3aaezqjalarGEtCiY
Q0J9xyF2R6Ve0htEOrytXRdn2CtJQPbRhiWD3lEUQUIsb/SoiwEbitCVKwjNb28Q
6KRNUkkr+FqFEwrYgDL/Q8HnmuJtzn4t34DLZ304HigxWqZUEDpKVAoJnLH6j3TX
3tpQU6g6JCBGU9ZeBltyGPXUcZVxmWnItoXkiqcu3NzWyj77fa3EKl2UElKDxvMG
Ugi8g9Ua2a4szLi5k+pp5RACVd1ALozBFr8QO7SJkNBCDhmyTjod04bo2RfqR4H5
074QgufpnDwbbmCqd30hgPChb24lvpSUBuCGkgSD4s4sk6lb5z1ryhTa+QpqBhsI
OVJN5WbzlEL5dtVuZLb6Ih5PC076jgXWUwPVEnj3pe+ngVgdBjCzpKajDYGA+VyV
yyLoY1qWLzvF2dmnYvd2cOADqDiQK/P0rgofFqMRLQDutroLI3BUEVXrJ0TDlhRn
njZpVlrKsIv1UFr60r8eINJLO795GvRogbEbrOvigFAC3sYtnYvaJFPTvtUKeWea
EGnnmJOcJL+qGxU1ZEvTXZlG6V0R4D53wZMgxwQTJyO14TQ0fdbRAW3OvHuFjbwb
b/Kwhrxybk41Z3AnJC9kuIN+RDQE3gGT6837vsv/53ykQW9KG8iCj8RP9QfhpazU
AaZhNpPhpZc7OpkYNKVTeB6e2UV9F4aRcrK146GW7xpV48xBAgWB6D9WR87rrgy1
VbKWf5DyIX1utA4T0Ru4UTnKCzVHdYk5jKbc6YeMA7HwDLRJoJFYZ03IXL1IpCDh
2w3nA4dIIfLq2GGTU2Acz4vLyxifXRbvMzKd3f6Xs6zYgU+9VFGkhwTOq/DZz8Ms
IP8HKBh5DpQ/Iu2uT4GQePEwpthoVfgch9z9JmRFIRadniXKyFSad2iYlYKMZOqI
/N0hK0svsUl0ge1Uc7rbsNCD02lv/fzaxSTY8946Pwl53/3uYSGJ/OAFfYR9R7uj
MQoffGqX/DgAaRoo5pvOLsfDDIABC63KBwyReqFvdIHhYpydCLJRFEL9UuJ1B77N
TLDEVcgzl0kxk0Rl6A4NQjGyGKc3Tzx6L+5rt4A8FiEAFzqfKkrUQjKT6kjutPj4
Kvd8y9PGYM9IEkKN1eX0B6a0DqmYsn9SvT3Cq4WBkxLEQQ2qamO+5RcLLoFzfAKQ
vTXkR/ZsBYK6pYgyQDCB2KFHWY0DPA83FpsSJxXR4/GCfC3UD4no5zOrHmBsKka6
Ya2SfQW3zBlHOf6VGY/vYWLQS/5EG1vSCnwk6ypPjcgQoo+bhYsc6MKDsCoYcMyU
ora5eGC0Mj8a4NbWE5zgiAmfh3herPL6fdCHZKmscPp3o0K9+ndzm4f0XmWJ0mur
ysjuV+9tWoYzfHNyCh+F0COpnWdC6dmhYQqxoJFGTeY=
`pragma protect end_protected
