��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI���!qp�6ht����B;dv
�[�܈
�/���t�!HO;���;��.$?�'�-#ܨ��q�X `*Ƈ'�e,��Sg�Bno~����1���V�0HA�=/�c�����)7!/2�����&��������N��Қ	Z�G�i؈�7ХP��^��S�T���4a��I����Zp^�B���,��1�W�؂���K�U��=k{�LcF���)��Idᦿ�_�Jy�����d��iN"����#�,^F"��.P�P�����9���})��ւ}�?�T��;_O�@0�|&���7cgKD��PD��댜2�.��%`:N���n�@�8�ݘ55{�K�l��߆,��`QJ���ɘV��kF�B��+]�4E�`�8�`�-��a$�$$�.~T������n`-*k���_�il�
�J��j�E�@��z5�o�v�ix��yK<��s}�F��x��Cn�$�"��u?�����c�<*��u��GI��:p���P��IDL���0uAf�t.�����G�چ�����_rǖ4�Z�Ϋ� D~%�Q�IM=�6������b�6R诩�a���!�T�fm�!@���VU��R��1��N~�x,xB:�c��А,R���#W���©�fIk ��xɲ�z2���Tl�xSW�g���JIe��OHb|��dvN1��~���fP��������{��Υ�������*~�#���f^f���k����U�EV#�Y��+�)_x��^3��eL��No@q4$u=|kҠi(��[��]��;_�]��AY���>+��I7kn��$�Bv�����}q?/pa傘&Eu2"-S�{]�Iv�Fr�5��}��H޿	T�ٴ�ڌ&�u����k��ь�Y�`��`e�ÈT��Вh�`q!6�WWڶ�_5t`һ���Q�a[��_�&�P���U}w�o�e[Y�K�%H�W��=�ģ �x�)3YS�������$SJ��|��s��L��C͒��c�$;�s_/o+�!���J`�����=��d�-���N	�N=S�!�\����˙|���:��H�d��x��5�j{�M��D����Qrs7��s2�։tt#���r�""��z]�u:��l^����Zq�
���uov@Ktी�H���(�+�B��HyGҪI���7CY��N��y�A����r�Pה�M�U5Xy|D�Y�WxPF�*���jqw����ט�0V��Z)��y<���⽛�M?�]�5���x��D��D�޹���.�i�ċ4dTl�.��*C�I씁���ZZo�OS������0��x�7v��Nh}n�t�Ͼ�<�*Q�"u�)���Q���ᇆ��.E��ts�
���:j#E��s�:[���������ZCNzG����B"�5���?JdR�W|@��qv:��U�E�7�'�Ԋ����B����\/�u�s�T#(�p�	��܂P�����D�����7�-�+p0^�� Y1�C+�����)���m��P�����5���S�FdX <�lm��ⱪ��-M-n�?3��!�J��@LN�RB�C�"bf�v�B�dy6�@1ۡD��.G�ql�W�1E���
�M��_v��B�6�h%PZ�)����;�;�|�K#����|�J5F���ᤡ���Έ�����#8�z�>\����ɾ�p] (heZ� 8У�Jށ=r���e[�D�2Hb�΍��s]��+<a4���6�����M�J=����>$���Vt�S'7��Du�3�o^�u ��d��a���|�H�=c[��G����}�ϝr"�:`��k�66��7��:'پ�iu���&J<�ʔ�������Z�֢vq����b�G��"S8��vB��b�b�r�)�fE��K���	�
��)/u� ���2q��熠O������i���R2��1|���JГ���t	�K�&"�p>�)pL"�L��5^�X�kӛi�x�mfi��	��I�⬩Q}Po�.�+e=�[as?;B�H�C�rUؕs�L��7W��u��iШ���D��-a�����q��\�̴������c�d!�'5Jz�R(�h��n�\A
u+�za��.�pPV�����w *�'�����y}.��(o�XI�|���yC�d�1RA���巳�E�b��"�Us�D2�����Ɲ��0�i��twz}dTb��N$N��7���h&��4ۣ_�t �;�,�u��j U�ţ�q�ŝ,�l}�8Q�vZ�7?/N��ܶ��ڟ��Y��.��V��vvL�}�Z���2���}��輾��]}�w-̈��؈dRb���W;�xىkLЙ����zd�/�ا!1]�aE�`ΫW[-ч&��+Id\�>�Io>5L��u4B̾���zܟתrt�	C�Fb���9�58#��P