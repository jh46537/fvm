��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ5,��kF��#��o`�Ylw�ve�ѹ{�S��@Лk�(5 ��#,�NN���)	7��Z����(iQ�|�Pr�b�j'�����j?Ɠ��OJ�$nr頑�I�N�����X�4�R�q	�8�*��D�6�o���4ss�X���M����+8ޑ��7�_6��0��j���ȇEga���gO� �>a�.&(JBl�j����y\+���^��c�Y	�P;�Z9C�	�$�Í=����qg�Rz���kIE�D>�^���0l_��K-#�Ii&T���Јv�s�a��-����'��Ŝ���rH���W�������z�Ѭ��$.8�,���gm[R���,F����g5V����#h�����Y�r'�s�qޚ
OmR}0�"d�/��N�3���������b\�$�S�C�#�/�J�����ES_~M������=v���7����]�4LCU��Cq(e�)6d�'�3IG��A=���Ʃ`��ӵ�u���x�".����v�� "W���R-��9]�]���2cP�3Mޚ@��U:I�=T����(ѸՌ��O\p=w���(z���]5se�����5��3�0u*F7�����D�up����1�M���&����Z�I��q���x���<�Y�o��e�>�U�X��G0��m��HC,k�k�	��K�^��Y�b��[G�5�g�@b3�����Rg��͹Uo���9��5ެN���r�0�:'���0�F��b|�c]=�+���{Tk���0�A�j�hn�7A�"�=�VC�����g��|��TT��c���^6��\I;��ۿ��K`��Y�����t�ܳ��+�Ar�[�� �96P2��ի�r�F�'�;��)�37�؝D��)O���S�}%�wn�P��{��Y}��͒����1��7�[{����B.�;�2^Vw�SXD��^��Bm��Ac`�'��ɝ@�!�>�l\K}wr>��lj�`"U��;��cPXX�O�G�B�.L��a�o�{�ڴI��5[2��^�`=�XĆ�:7۸���	<��U�p��)�Hdt�ºr�����؉�Ԅ<J�F���4M���,�E5��DLe i��rO��0�Y}���Uo���z� ��IR�̔�ڕ���`��G`⫽�?�'! Wv�0Z�5U� e�L3�٣Ǘ��%��V.N�Rr���H�n��D�|�B�נV;٪���������1}!qr�k��Ãti�E����[տ#�;Z��
�	�K�*S�c�/F�LT�$�PV�D߫)���(?{-\=���3�q�����2�� �@)�����#��k=Dp_~�Kn��Cm�U��8U�tk�L�4�Ő�u�e�]��j�HpsMEI�"�������%G�u�=��u������>�����<Wث���Լ�Σ����j	ʀ	9q/a������@�9�Ut;u\��fVO��V�����<��~�w�������S�`>�^|d���b@�z���Gh���Z�8x�Jw�8lI�C<��*�����Z�Z�h�2w��W����*�S2����~��<I�D'���aI-O��,�]�p��5?�%�d�|������7Ϛ�'�?��O�ӕS�,ߥ4��sA~���P����