��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�	�O���|�Kv�_e�|g�w@?"����W� �5���_� b��d���b��*���k����z��汥Fv���-T b�^ۮ4y��5�X|�{���{l�m�#&�|���^a�$�� m*�2�0ƸI��ii8�>�R�������09C��}[�"�A��  �oޜ��䳠�p�*j�=VUF@8��4d��z&ʱ��áDD�]H��Ȇ�_Ӛ-�L����!/���?�#����cu�j���R�F�k��h��x���:$��cGhrDվ~��`\�H��Rd�)�̸��=�tNҺ��J�JӸ,������Y==Tl	ۀF/U��Nf���Ųa܋� �M�	���i�|F'}/�^�q�����4�-+�puD<�O��7��?�0�C���= u6����Cb_}/k��ϭ�F��Nz���h�cj�SGD]�;_��W#���#*)sܹ!�l��mD��A�>��u�i8���m�t��Ņ\;�j����f��{�Q?���@�Rʂ��A�7 ���Y��g��=��`��uz&\DڍG�<��V�*W.�H�ߵ%��H��?5��s�d���ޔ���: �����lQ��-t�Ҋ��7cT��f}ʏɎ`A:�ݼ��d�Ӹ-�f|�Ɖ��E����Ȗ�z"sّq���I��
��x\�qs���ƥ�[H)��3�Ԏ�ͷ� ��Y�u4�y�� |P�E��"f��f�
U ���m9;�JUD=; ����)GU�S��%���m���*֞*E�?6nЭ}��=����R�EH�,9�&ma���'��w�D\�'?V����rI.����d�\P����x���1d�
%�o͗-�&͓�y�w�@�^MŪ�����^��ؓ2��ύ�F'�.�V	�^Gz��[�аm+s�Z�K��f|���ˏ�������Q��b�=�S�tU�1������j'��Iwi����P��I�XZ�~�#�H4�8^'��Э���*:d���C�.�1��+�{a���C\��\Ͷd�!X��Äk��G��ԅ�lb��gQ��`���"uX�׀�:�/�)Z���gUȮ��E��Z�0pJ���5�i�S��U�J��cQ.r�_�(�X%S@Tqa��:0�lǱS�F�OK��L��.[
�B�KH�W��l�v	����	`~������7�E#��J�Q1�ašn��eƀ�������e�gґF>LJkK�w� �5�A��g��t)o���X� v�-h��>�>D�K)i�d���g�q����tYr6�]���&d�n�_�&J��vt������kf�"ΛY�����X�Ca���c��B8%��FN9Úpo���!��*����<O=I�򷲤})f���`(�k��(�;_��vT�z Z��\I��>W�k7�v(��m�o��A�;>c�`��w|��=�5A"A��ꂨ��i��:��꾙�t�?٥��sN��*���Eq7j�@�8(��x.�ʋ�<��Q_>˻��n�����@��l.�"�BS;��K5,�F�2}�L+\	�$�!�z�,�k�S��v	��'��܊��;��vΦ��[�FXF.w���w!���/j�K�41�B�q�<�����f�9fd>a@�eJ#��Ϩ5QeP����~��Z6�A �G:̱�8��b��0�:n0z�ի1O����=���x�U�;oz�L�e������0M�7��@�l�.w��[0��"7T��G��Gꈞj$�!�tPk/����I�>�t��PkΡ$ǘ����ݿ54��E�� ڙ�W�� ����o6��.�)�E&����P<aA��+��U��Mǽ�!�)tot �KG��߼njt�#/�x�ޚD:��� :ސ"��m:}���z�QvG/#>�'�[A�t�1�Z��@��]�{�0����L�@e��i�C�h�ɶ�� �/{;/�D��}p.}ǩR>�p[��`r�v��������Ht�R������/��G쳈�q��v�U�$T&�?2�~3)���$�r�N�N-`�eb�� �A4wr|R9#��0@��pG�W�ׂ2дc�n�s�Lu�m�l����TVss��k^f��_����=o�s+'�����}�Ǳ��:N��t�! �k�z�}����Z��K���u)k/ΎJa�������EE�5��J�P�� 7H�}q�H:�"s���c��@�!�	)�H�:z_sg�2u�'�Z�xyY��l`Ѷ���+��_˄���� NU��*S��?��'�(T��T�L`��P	v(K�%�zC%�[��OE��^J�"N%: ObMH'��w�f%9�|�{���A�浓P�ٹVR��:��j�"�/Qn+�ӣR+P�P��/m��1�Nz
�����j �#�����Q�:Ř�I������3+isӸp�i��Ɉ<#�w��몵��;q?�?���Í�''�c���*g�T����Mª���nn��	�]%��*���z�/�%=3|��c�������b�> �"�<���5I�7�R�q>������A��x#�U�vyzv�����
A�~.�\��������S���� p������c�s���Ī�_����+H�������id��?�c�H[�Qڨ ��`�.���F��,ؿ�j�i�}��g�_��-�A��7n_��2�uգ8�Ѻ{�a�{߃h��/����-�r�Y�t��F�F_��/�'Դn\N���	s_[0���T���b��dSD�z��k$s����e��;
Ib�]I���d=̈ő�" |���]":9#�U��.��vߚ������<�*�:�V�/6�()�IBG�����ydٌ���7X���߼�OV+}�8ł��EShX"��,�CB������=����o�;���q��x��=f
������M'�s�e	!�V0������2�`%�RD�ٟ8�� ��Z�W���=�)9	 m��/�)��I=�#[L-6�6ϴ�/MT�k�+����!�j��K���BgS�6b*���ה'���pm�<v�>k�u��P>j*@D�wR��X�)�Lae�q�*n�56�_����q5�-2H6��ٺ)��U�����*M=s8�Kn�Z9|O�n�x��dO2E8�Xl:ǞI�PD�NJI��tI�ed�)x��V@mi2q�8�u���$e���6@�ɒ�7����U�>�.��|���?�%�ߙ�(.�����`6���h���z������ZJ��Z`jO��`�4Q�W�����cdv�5��|����^��ދ���)�� U��+��)�����&�x z��J�t�!�H�����3_�NCo��ь�9�X :a���K�z�~#
��6�ɞ�8�.*Н�F{b������z��� !���a�ģЩ�B�X�芖�,�K��?�������_d��ް'IML��JBH��!덲��i4��|r{
�(Eh�
�����5�j�� R|]T��)Qq��b����i33�R���Y��F�V$5|ٞ4�P�wG>����j��3q|�W���|��|A��0߇��eը�W����]U�w�ۓ�K(��UǢ����B��=!2�t�V2t�O�;��,����e�	��"&$��c���\�(Nآ1Ȳz���1|��J�� �@voxj��곿�!�����5͛�u1G^�P��f�L���m �]������/?i�X�$�9�Y_�bK�j4X�zl��ñ��s��r�Ʃ��A�l!��RP��҄����g)�3S����o�v��h�V82�D�! bE�!�K���۹�%�1I��ߚ�t6@���㒣���.�A���qOO�T�G�&��ni���*���m��/3�eaL�Ōz�Z��8:��y����~�����M{3��6�Տ4�����{A��NY�U#��(�f|5�IG� C���XqF��̰�����7,�m,X3��@�U�&�=�C46����'���?3��n��
> (\����>�8E#c����E�ɯ%����`�6�߈ʁ��!��JWQ`�<EK[�>�m|6����!aV����St ν��b��߬�BM
����ɗTm�SB�w��:��ۡ�
RY�[� �� H���f!7�:l�����}'���f�ݎ�}��Dr�{k~�;ֆ��t����ܪ���1��ӓv��mD%쵒ĭyc�hG�cotR�+��c��}޹�\2���3T��YOn<�EY�r��/���%'�%ٹˊU
�u�K��ԑ߱���p�2�Ob���Y\�y,�|��[FSx��ZrsϤ�U��֟;�ٍ��2
,E'#�Pb�l�>��09�F���a�P
�T��xD��^R���g�S��������E�Bc7�"���(�RtF�Qa ����F�He3i᫊�ٔ�Q"�����>#>78q�����e��4��J�Ҫ�LY� ǝ��+z���X�v���iC1cw*�
�I{K���ɣ��k��zƚ�Oƶ��\ɔ�I�23G�<����̊���̭v$�^�P�s4?Εz1ʏX�ݷ�ZjGc��rʚ����J�f�?(f���ϸ��>@nm��,Zg��2n��`a���X���믁:At�eĖ<�-ӿ%oj%�/�s_�/<�
�5��W�(������TFȰ�B=G�[�5�l�:���流g�P�l���+��,�:�ˠ�;,�	l�Z�EZn����;��G�e1M����_��=���\ @���~�)��p�^�KY7(Æ���m��G���:BB�5B]�5=�I���{ו���Q~'�A�dp��W5��y�ue�+`Q���;~þO��%"ۯ�#�����"ȵ���d������t<��s*eJ�8���N�\�"=,�{=���=���M�b��7?e)_#�Xsㄿ�Ֆ�H/����V����f�)"��h��ۯn��i�[W�"\�*"�a�ⰳM� %)oQV_�2+�6��r �՚wo���0��-�xx�U�6?-5n����#@`bJ&��8gQ�W�Z
������\b�=ȰWQw�����"uA��?���K�Z��GM�CN����p��y�9v�4<���4J���� ��reЪsC��z<�(LgT��I�