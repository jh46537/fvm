��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM�
Ɨ�j18a�W@H&0PoΚ|$�;Z��l�)Gh�V B*��f���@1o ��-:�"W[<����Q��.�Le�B-�S1&pbQ]�}�H�a�{VAG�-Ŵ��ܺ�PaS��鏫9�#�z�)eG������tY�$��Ё���~��Ή�$�U���J	�!'�[�p�Ş<��3Q�1-X�8D��29	h�t�4�}~�&�o�o����lp���l��|����oM���fr�����yv����:�b��L�L��8�ާr�Jqw(:�f������4
���cg�MG/}7~#A/��Q�)�ei��
�;g��MM���`{�2�/�v^b �V{����,(^��d��6�L(�/|�m�������8VvM�d�NM�@)�z�	oi�|'폕�^l[5I�6�V�^]_Sy7�>I,�ƺs�ypkj۷AROX��z8??r����~W�V��v�*�2���ã��_]""�*�Q��3��� 4��lG�n�2�Q���x>�t-PĔ��[z9 +�k_ĕW�kH�?�(o
<��bJ��+_ٯ0�륯B7�1���f��md	����\�$���0H����E��܍�S2�2
0t�������6[�$��.�vx$k��6��:,M)���;�s�38�\c>���O�H��������.�G�{���2<��B��M�`����d����˫�2D�+">K-^�Wڭj�X��v��g#�,��d�W�n"r6ցq�;�x�)zמ鸇g9?e��WLhb����e�諦rB��6|��0�!��t����u��[���|��n�a��KpQ)�oFl퓔���A֨�C�c��)�pn�E�o�-�e(��<
�_k�~��4�O9�=�=����k�zz�$�Hqh��[i�X��TS��Fc�����z�2z�p��*mh
��T��Uڥd7+O��a0/���ى�ňQ5#�2h=��}�&��1�n�A`R/W���N\��m������ƣ�A�D�`1 ��0�,	DEM��	��[=���x`���9uV�g3Q�#��/��q�;��zWW��n�S%å\�!P}���8��K����~��t���R���
��;S����X���֎m �J:�$�U�}��(Ð���{�4����(�a���
L��t�
-�V�P7\%o���X�2����&��hH�~��[ޟNy:�-<�s�[�Yu�����֥4+ǊF ��޿�M�ai�O{��:4+�[��m�cº�A��H�Bw���^ �t���\����&�DfY!*-3�Y��"�7d?�� C^��>��sm�pxҵ�q�|��2�hS�o����us^�fKP����r"S��3=��If�*���e,���p��-)�a��얷��6l�y_�]�D��#>�$��b ,`���{�} �$�u��$}*�SbŴ.!>���g��m��x9���O���)m3�&�j��U��h�Нt���t�\�^��o�8>Ă;��n���nƖ1�yW�E��.���m�Irt�1��=A0�b�V�?(�[n�4���3e����#X�k�V��9�%v�k��9>��N�pς�hש�=��&��u&m�q�V���JQ�{�a�]����D���nT�*��-�0
j���ؽ�.��