��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,��F�X|�ע��R$�O���J	c���1<KQ�0=��!�n]2QJ�ta|zI��s�.�ŧ80qб�W�1;Y��Vu�B�@3(����H�?��{�����zԻd-c���]�`E�W�~��f�W��c-����"�@pG*�����CYC����޲v��&�2��[�9)�����l�wZ�c0$��"��"k�a�R���pǭ�R3�=:�2f��<���g�&�x��n���[嬋��^�M�d�?U���n_?6��l��� %����7GE��$�������ys�~�u�5~�,'��FU�g6G�ȩ9�^�ʓ��feQL9��t��o��R�W�"��Xi��xF��'��c�=$*��͠��(�%�<*�cz�{A��β��Vui�����P��?��A�t�U�\+\���;Ձ���$��q����K))�D�/���lA쩏!� �T<��Q �<ņVS�aY�)�d�G�����a�=����$�� ��J}���oQ.��$u�-[ͨ�{YݹT���)[ �)��Vu���6գ��&]���ϴq�$�w+�pǬY'��ge5	�X����U�2!F72AR'��$:��۩���7���m����c��fQ��zz]��4R��ac�;^�D�Ce�Xh[/�q�TYBm��`�b윳����ء$�ߘi�s#��p��%{|\���*2�v�<hp���E��>�`S�Bt�
�ڴ���lLv�����F%�����K���z�Y�%���㹀���㬀V<g�����uC�}�>��\�rD�7��ʐU̵�[�0i��L)��Hh�Xｇ�a�
a]�0fr�~	�לΈ�����s�� H\���\xR��|6G.��'���YLS�(�% �Տ�{�\G�P1�<�0�"֨�ңkF�D�ղ�3��@�U�/S�<i,ܡ#K��f��Ȟ.��3K�א��01�ꃓ�L�Y�,��~"� ��U��1�P��W��֔��snb���v�t��d��d�a"B�E��d��Y��`-�KWu&���r������o���Ou��h�(s�|v3:Pāˢ���-�[;^� zU�(�>�m$�~��~K��h��D��^_Lc2�6���l�*�P��J�ޙ b�,��O���鏫'2^�"�֖�Yjt(�����D�T���\�,�.����<'ſ�����2���Xnx�S��^۽#D�x�90ȏU�n��i.l��z�^o�������E=�0:ug�/��1RS{��똉`Ӝ%�*�V{mf���7V@�)z��t�ie)ڟ�%v�Vc��I�[�, ���RNe��l��u4^#�)6۱�4h�%�f���>���n6�<��S���Z�F�(W���L�c�2���i材=��)/�M��h�wPZ��;�R�t�Z�ۤl�ԆU�sC��{�|���q��@f�̀H�9� D�m���d<��a�pO;�>cV�I|[�;?���	��i��<�F�R+��O�Ec*o�'�?W�Ƽ8�ՒMQ��X�lUuce��ꥲQ�uZ��<Fڪ<���9ۛzP�Ig�I�z��O�ӎ�P�N24��V"�Oa�*�\�a5���?nGOl��4W�PMyíN��SТoK��18W_�����t�:��G8��D	Gҧl]�𕙞�+m��s-�k6� �{��;u���h`y���Ew�ARj_,C���^���ć�_{�!_%) P��*�����v'�W��3�����G�W��?u\�b��<[�m��IŎ��4k2��	�T�Ow9�}ߙ���jRzM2$/>
Ryd�R��*Ud"Y.�|}R��@��q-0!����Q��O'��|^ZB�c�/�~|��x��Q/��8	�����c���8�O�(��V('�~�����j瑗I�%b��/����_z�I��;���Qu���(�@e1�q%�'B���Z��܂�¯ٍBja
��&0���X��,�����q��z�u�� ��tsWp=��D��®M �(�Ϯqxm����+dM��ɗ�.�g��/��e-	B�i�r���5C�R��h �]��ss��uv��n���~��T� �)� �'y仂��~����b��l_�q��?��"�P���С|3cHg[��{���Az�1g8T�_������}��T��1s�Y�nv$�+��A��1:�^��F�e<�m,$>�����,=Z-& |q��U�� wh�u��}"�:�
��E�E��Όn+��ƅ��>X��[��׺����NlP M[�&��x������d�Vo�����n!0�1-?�-�R{V��Rv���g�S�
Q��BUHP�Z��;�?M��r��%Ѯ��s�w�C�Q��ɨX�e-
�B����6E*�!�b���*}{!
y�C�ޟ����W���6s�7�a �џ9OA����Z��Jo���5Q�5.�S-#�K��`��[��T��,�=}ٍ�4���;��rvO�((��_oJ&�fjo>��=�BUC��n+!3H!�T������l���O=KZ�+=6�7�S�:c���%QQ""f�Nd��?�m�����֍��߸M��;!����Ǉ�~'�@}����	/����5^��|���_1�Fg��E:�na�3��f��n���?@ΦU�������6af8D�#)�3>�iq�'��kG!���g�ʙ~]_gUn�a�l��Ro|��l�%��
�ɿ����ݷn�/�t�i��@\�_m����,��Qm�暷[�^�T��S�Q
ҥ����]P7��=�!���[ �@�qrN�m?�h-������=�%���f�뢁PO�k4l���o�J^��c)��9$S��)�����jD �ht�u�|Z���K��z�!�ۈ���t8/}a/�T[
�Y=x���˘:�L�;��M�l���>*ݮ��eti�tʷ l����7_��!�V1y�/q+VQ7bS6�gn��N��w��g�Q+�ok]�)����	���eWgd B׽�Óm�4�m� �Y� !�fi�7��@��9����O�xgCĒR-���9�}�G�J�j���a����S�3�H��t��3��E0a��g�t=�?�q��,���n�j���֖��4CfL�d�6Ul_�S|�g
r���F�MT�qo�^߫ه��Tvh�p�]g_2l-a�2��'��3=j�6u�$[Ø�v��DoU7��\&g�������b�mq�@���8� ��o%K;GE"���%	^�-�JP���k�]^{���Y}+W^�0�<��ѽ�^�oo�U��0k�$�WF���\����t]*4�]�f9V���	����E����!�CC7�#�.�X�؎>V�!KM��h�rB" RI}Y״�G����M�Z�=��M�?k()����GW�N3Yny��*1T�ܬ�*��l��\b�钟
���W�O��l�oRQjcc_�@��#a#g��_�0`��drA��x��&m��k�����LT�B�IS,�R�w�/��{2�TI/��T�x����>�a`;^q�Y�5���
.r� 4_T�⯱��-�{������_�$P�ʆC(m��i�\�M�K #D%Tr<�4>Ƀb��8���f�D狵t JTs�&4�S+���N�~�ݳ����z�2�s�YV�nS�#��2������X��
`MM��f�h�}t����F�c�e�gT��J�%v2a�le�n���{�(Xt��q���q�ܤ��
֧�� eW���٧o�����EGQ̀S1icW�8����h�Jc���ʂ�1JN1%h��י��T��4��T�.%w�I�{��d��wg�qg���� �m蟨��؂%c�]�,��kh�B�G̣�ܻu`���{�������g�3���ĐJA>��EP�~&C4�����@����`��~?�A=����7�N�6��r�zξL���\d2��2G�����f����)
T��:d},㓅F4C�aӪ,#��UV�{�c�hYc�ז�,�5�-��S��(���Ջf@�����cM�DP�t �xLغ����ᢱ�L�3l|%��T�����:� �p5�.�3DQ�����TGzH�����v��֩��"�W�!]��.DL]!zР?Ⓘ���X��j	�a:�;1���\>�c�x�*�l�ӒF����2�%Tg����� C��6�!���=���ъj,�F�t��W}�:���x�wn$��h����6��EaV��"fn��Vȡ�2���$�51;Rjv�~쥠7�f�z��Go<T�#F��a��	�|I���*���Ez����6d����S�|��d��� j6ƛ����\�_�������p5!|��jI��v&rs"�L��#��V��IE�A��VqVp�����Щ-<�^�7W��`^p�Gw0�s:L>��-ER ���
P��O��cs2��3�B��g&� �|�-�tb?�	 �E����*���Sm7�y��q����S&I�*Q����v�)��w�V=M��<p�|��K�gH|�����3��ֻ�W��[�,�!���?&4"��R�X�<X�mv�K�5�t�|C9$G3n�FO���,3�g�yx:W�:��L!�ԗ[��b N�e�=5s�'�}�EV�KL	7'��o@�?�,exs�i�aEjaTJP��iJ���vI�w�5`2iW�sՄ<X~��f��@�_�re40`Z���O��KM@=B@�#ˢ�
�v�C��f�^�!��qq�|.н �%Ɩe�
�)ԟ �^��z�ĩH<��Q�G#�^=��1��Հ�3�؀�C|�,�"��2�(��A���IӇ	O�>� [�`߻�Rzt�Lu��^�f�n�&Z�	@){��������AS��{�fn�F�SQd%HW�o�'j�=��KOp�㾂q�kr�nD골įI/��𣁈�������@���o�[P��̈́'�ԷJzɏ"�!f9�
K�S%��T�B2���r��a��ѳ[d�o��J�WQo�JQ|r�f	� I����!�J$����L��(���{��X�O�6wuM�;�P�k$7nƍ4F��ė��