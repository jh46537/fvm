��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�]d�L=3	w5��?�N��A-�5�P����B�[���훋�^b�sG(�dt�.KR��:z��X�X�8,E��c��DA��G���\�9��=�����*z?��'�]?�VUv�.���Ԩ0���L�sB�Ξ�U;�[�B����gM�1�·܅�̵�$����Q��^����W�M5�}�<`}�]مڦx�|KW��(`G=2[�'J��m����5�E�0�d�ܩT�I�f�[9���wt��f>�eo��k��F�����Z�jz1���(�+־876�����O��|"��Y݄v ��#�<�;�dWZ3wP��3�Λ�v����6ě�M6Ш]� �ಳ \��+��1��U������
����$8b� 0h�H%˂��>�cxf�T=qE�Dʱy�B���	��cS��4���f#�72 ̨�Sa9���;.�,�b�:_�X;��<_���)o.x,F�t䪫"���	�8`}�5�l|���s#9�T-&�͹Ǣ�����>%zhDa���M���ǒ�T��	R��#�ݍ��[cw�*��tI���Z/�ަ�Y�Ӊr�����)�C��s�:���$�7t���}��eV>�doa��)|��2��e�O r�r@s}�o� �i���j�y��0�% ����	�7F.?S�.k�=�
93۟��1>/�@o�o�C�~����RS����ݤ	e6�c��7�(�]���w�Oh��E�~�:�"!�_�ª���w�gĵ�ŧ'���9"o1��������uχ�,���;�H��l��ޛ*��}/qDA��w���&�BvT=�M�&���Pz�d�U��t$ϩ�`���F%��g�8_Fh=��H�S�60xJ��f��1�D3I�X0W�XM���B�cx���l�I����d9�z`�+��b,!mfTx�{�_|�E�q��L&5�8����;0��n���cUo��7��1%�)W4��T�Q�[����j�sI>�1��AP9a�t����Z��(i�b@t>*L�9�lw�s�xPL�<ۺ# 퉄i� ɇ*��<y/�Jǽ���	-gN��������|��J��ӦV��كE��d��E���+�>Xs���H}��jI�"�E�TW��s���l��L{8��T�*�e����`�� ����t��3�����ȏ�%$�>��jE����]� {���|�� ��S�c��Ԍ
��{�Xt�3�U����?�s�b:����aa�� hƽ��Us@�T-�6�5� ̓R�$L�e�R��$z�}�1�(D3� .���h�T���K��Ɵ�VN^���������ש��W9�84 ��R)�$H�9�T�b��T)����/�k�f��/v���\>Oc?�쭙BK���D�,��7:�G8�5���V�p�1Uh/ﾯ�!����â�<oY]�o���]�K��7�A���S�Yy��ˢy(6�`t�~�~�|���<"�qK���2�i8^���_��6Ǥ�mhT��
��E����V�v(k�CWu��e&��E�nC6NF��q�tp�߽�>4l�诵	�$���2���⃺��[���)���������5���,ڷt���=�]�]C��D)����@~������kӦ��f�%w�ᯝ�8�x?���1'�_ �f�u�*��g�Y��y����J!-�PT��C��Z&��t;�o��6a�r:��ن�n'�w�|�[�6}�`E��C	�K�~s��ISd��ݰ������e���2��2m��a2>�1���y�Z,��J|,�nI� 0[�^[�}e ���N�kI���<��B�
�Z�طV�k �d��������ذ_n�p%�7#8X'��ŮO�� /�(n�	���{ZR�ڌ�(hXW���>t��7��cD�-�t����-�RT�2CI'��]��"7-K��F��G&���CMM���f���9<���^ޯg[#�2� ����eԍ��>�T3���0�JUG�1셞�4��N��&h��6m:��5�:��B�p�}��eQ>&���
1Ko��sY�)S[�K9�!�`f��爛����}o?4\�] E7޽�����ʬjb�h�JE�
�/�������.�q�>f�M�smC�+��MG�u���ӿ Zj/5A�y�囄��L*(_o�׹F_����f�$[>Pp�W��]Au�[m����c|�ު���%���# �"1��d�'l!.���Ϛk��C�v��@��^�	���t�%�e��ʓ
�l�o�!�95|dTK�I��nr��d�?�gW�OF(�Ҙ+�L�&e�!b��z;v��f7�����|��%7��B�G�&�8��@Y	Qe綯�?w��+L'��/�4��#�n{*#	R����<>:#�}�;���qҨ�(�3�l�+A��p�p��7R;l.�~���; Ї�?h�c�a�x�ҊK$�V�Ό&}ۑA1� 7���CN���<FE��Ѩ;;�6���Ի�M�AL�E�h�|���Fk�x���)h���$=^�5�SL��I���#:�Y�0ҏ6p_� �F����3j��Y�)\��~V�J��V�p��|�ZL��[�F��nQ�[�c�SkA�3��_�B�\�	���|��{�ej"�8���{ӫ@�	q�@������˷�b{�N��)Q�K����`��Cb�)��˄��n�mU�G.����Z|��-ӧ �2c����~��0��C����ɄY�Ҧч�E=�Y~�0�����]4;�ń��#Wٹ����Dn<G7�W�U ��L�Ւ:���!�Y��1�8J�mP����G۠��m��B��,RF];��iStpC����%_�q�eEt>���W��䱴��g�ļ�W���6�m<���H]����[jL�n��Vz�4f�DX��Ċ�����1�����,���c44�R�GY�����D"S�A�`�9ݲ�d��xt �R\QR<��Fu  j\��qs�?� ��{ch����|R����Ǧ԰/�a�W��vr����D�g	�U]O �����h�n��&�F3���V�B!��΢'�������4u����F�G��5#�Un�$��{���_���D���x�ȱ��Q�����0�_����!�㇨+<Mֆ��O4�,����7�Nq��l�*<��+Л��"3��2�&��f*(��9�vY'p��GD���dݝ�M2��S@�::����!�y���dך{0gw�=7��,�4~���Yek� �s��N��;����JW�?^�����" c��n��g�)����n����?�Zk��Z��B⿭������>�J����jZ.�������3|��9d�z�u�!�W>�DQ+-S��9����!c�[Ժ�90�+wb�oD���|N�!Z<�v����Y�	ع )tVN�B+k�Op�:�z���r5K�)���)ǟ��2`�?��4����r�O�<mH�趦�;�H Y��rQkT�v�h[�+J_ij�2(�plJ���6l(OL�jO_��dn0�<�Rkϋ!���C3��&ނ���[
r1�VB��-@:���/��ƙ�uc�z��nU�֒��8���s���^�AU��鯊)N|�n~�<�";dpf����1d��t!0��$6�T�\�L��
4��0i�Rg���?x���85�Ӷt��V���I������2]�>���Z��NN���T"�9��u}���پ\�>��,����X���.'H��.�e���oO{?#�t1���S� �#Z��3P�s�c�:�٬	��3�	�&���"���T���v#N�U8�-b3蠉��+�Qܡ����lqO'@`��߄١M^Z-�Cr���^��!��,|�-QK� ����s�� �p�,?�f|��3,���2Ѷ^��%}s���9i����3��Ƣ�Ʋ�*�,�+�rd��x���ϼ���{=��*A�������/"����L�uCd�ٌ��?���\�x�ጅ^���+	ߔ��z�D���y~=yB�����zlas���QR��w1��|�\�p���(�yZ'�FS*YjTs��h�3W���l��TcŊ��]2%"�D 	���6�����j?��v��XV�:�L}WH!�ɳjr�n��^�����������Wo�����n��]��o~�t��$��(ɬi�*��
��q�-����F%���cָ�w3Z��Iq�cl�,I���L�!H7jEw�N���ˊ�dJ)c� t �f��ͪ%��]SN�X��^�
�M�܄'��A�21�{H:�?��,���޻=�McB���4�fr��X�c�K�_��폭�FSVZb�w?�'�����(�[@���L�t�aHd��M�ھv6�rV"=8D(�ZA����)2�ߐΕ����+��*�$KYM�B�К�����a��N���̢!8+ٮ�C;0̰�v���-$/�#j;߬4�U���4N�Z��h2�M6�y̬��H�^�ۃ�X�=��8��Pz$+)�����l���G*�]��<�n �],}�Ҿ��p�b�+3WVp��z�i4������Ua�I��Z���B-��ߩA��j2��zJ��m�m�5z�ƽ!>�FLғ�f��Ѻ��Y����@�>:?�UI��Dck��7TF�� K��A�i$M�Dr�[�mh�)V���n�M��R-L��9\�?\}�,��)W��C�OӦIMc,H;����R��[�x��T���w`p�0t�h��g��g��d$�����bn}��%K�^���*����@�E��b]��Y�+CAlC4y]��߶(�А�x
s�H�^��n�G� &�T֥ ���>��"�R����p��ß[ ���B7J����w����-|�y��A����m��@Dam��z�7n����)�%�����H���5]ӓ�'��+��tq�T:yY�<l7�Yt�o%�){�Tz���m;�:�}�1�'&CO����w$�� �j})�d��������,��`"�Q���H&�����gDĕ�����u���^L�Aj�ܿQ1W
 4�}���4X�jD)��Ho�Zܡj.���g�eZnO�pθD]�����w�7��w�s�i�#���f)���:"l����cCU1�#R!m�\q#} A$�`_����Ku<C�x��=]�_�.^��+�a7���I��Ձ���E�������
	��?�폹p���Y:��̐�f�L�Ya)͢�� Μ������ʖ� 9Ut��3r_$���!��|��+zL����b�d>ǭ�EO��ݒ�<a&�Q�互���o�w��ܭ^q8\1Q���+/^;��$<�ô�vC"?n
K���� ��eBuf�o�}�, b�j򹥂hc���{�v�ƣ��[?�+9���]�뤽���*ܶ�i��Z �R~Ǳy"�ٮT�pn;��OV�JV䅲ġ�~
��:���H�̓@�+�������nS����ӔO��B����,��`��`�
WF�go�E5�W�q�rØ��j۵��g&��D�W�{>�t����:K��Z ���l�ǻ��8��λr!�%V�IF��v��:�<�;��ZT
h@@�/tƜU.����ݢ{|q����כڜ�ۣݠ�T*��1΂p|��iBq��P�d�V������[3R5���� �z����?uC�kX��Й��;��=��X7��Q"����a�-M������`qVkŧ:�e�+�֐�9@��C��d��?1U�F�к�ٌ��
��Ww��V�5Y�Q���i���%�s�������
*_sQ�
���C�cS.0�/���bSp�٤m��F灨��n;�F?_���"g;./�ޜ����u�u��D��z���l �a	PٵjdW�tum��aC���Y�o<�g�D}�e���5������r���[�0��¾i���'��C	s�R�?:WՅ�f�=�����Ԓ�|!yx�7d�����bI%pX��A��8�}�W����z��5t\�E�y�Rw��#Y(6�y�2��5��b��#��P�|o�;.v��^���fJ���1$b�j�O-?Z�e�#���?�<l�8�"�O����p��� x1yn�ꉲI�sa���,�
>�>� ���0�a�`����������6��..[S��7\ܧ#"t>�ks��������B{]���7����i�!"��W��u�$����:߇�K�+� L'����Ko�M��x1 'f�G�)Y1OCRq5�%��Ra|B泧�S�hMؙx�ġ÷�����3Z#�ퟳrt�?
:�&V�ŗf�j���9����� �x7p'Z䬨���T�_�T:����%���_��7�ph�x���B��0;r�ɳa2%�vZy�9Ϲ!m�IU�}��e�{���<�R�va�'5�Bh��kˍ�zEnRъǆc1�OG��U	k��n�w�zkjtg��<Ȣ�V�I\$����� �ԝj�ꨚ1n��bE@���k�؋�
HV%m�����Hzl/�)p�	u4�ހ��Q�)23�\��e�c��
4L���!�<;�ѢM"�L��נ��)|���W)[JZ�1�3����vr���cg�d'�]Ț��.mØ���t�����o"=_���M�nF��9 ��#qZ^�i�Vt_V���{���p�0�́O���(30�~����y��j��ţ�S�f�gd�@{��]{r!F�����0�/\�ɴ�qz�т+8���6HDY^�5�U4������g��_41������?���E��w��n�w�W9T�Z������� 63_�Dx.���W��i ��������7�C�	k������Ȯ0�~����6ې��X�7ʋ,`�� 2�#ӣ�`;�h:^�H!�(��c�b�'�P��6��i`����>a���r`F�s�`�E�U�"*��ځ�q��4;���}�j��|�4j�n��U�ұ\��tu:�$`s�������w����>&Gӛ�ۯM�'ɹv��քk���%1Ma��5�X�:��� �]�������q=$�Go�]��LE�Uj|OC����t( P�y ���'��׎*� ��' s�O�6���C)�,#����@�$!G'(�J2ʐ���?kP��^�t�#����D����.�n���9�L�R�T��P��\��* ���	�O���&�<�Dst�|�"G�%֐G_�7�*���ѡu�is�'�s��ˢ��o{=a��� �.v���͊�Ok�F>%-GUqN(�7�Owi�1���G�j��E��"M��NK&��ab/Y�����ט&5I��ᇯ��š����D>�%㊵~�I���3YР�2T��� �xb�	~.B5�L���)��Ҫ���S��C;����}�S��A�uA�_�1�E�!Xԡ0Ds��,zɛ<�Ȃ��;�I9�X �X��)��+� 
�M�7����p�pS�+�t)L8d�z�He��=6	p�n�W��O,t���>�<����W����iIsA����ǦF�+�����]T�u�Z�,�,jz�Q$�]m�R�V��1ұ��?6�A�"�����n}�z�W�_��lc�D�	�#s]bxG����/5$oo+�G"?�)~�T�$�k�������6T�N\��FzN�����|�ڴ�^C�@lwl~�v��gd��s��"P�8�����a���h`M���;����L��� (�o.`i��=j	�И�
B����o�h_�-����{L��}�`Z� r��]>�좂ym���&�I��DY^��,qS�K�eݶv@A�� �����}?94���RF����2�����^���5��g��r!"�Q��f�ެ��[�V�nYI��IB��z��ķy��`^X��²y���i���ޑ6e��A����eY�:J��E���_�-|����$��t�W�v�R�m�,V�D)w�V��9��!�I��,t	s�}����ÀᏡ���B,�	z�:�*K>G����O�9�e\V�;�8�LE���I���i��3��O�,S�t��j��]�"]JP�}��ð�f3��b���W�ڻO��=�H��	6l��Ŷ�Gn��e�W�tR\DB��C�_<*�R��-7"��M���(�3�i��`�«`ـֿ�ב�-�[�|a9���*��p�A�̈́r���t�P���9��i�TG�@�)R��?ʿ���c��}�8��.k��P��t�dBL�>Ƴ^Ls�eT����HT�Q��)���t�
F���`�]HN	=p��u� ^>%�`����5�5U�-�u�q����Z|����䌵�+WM]�-��
f�����3(��a��.�Pފ,w��(]e��z8(�Ѽe��,��'b�<ؘ�e�f ���]�+�4��m!i_��9r�z�OK֖�P�u�t<��Lw�ZZ�w-�\H�`�SD��������9��L;�O�!L�L)ܑ�%��7_v$����w�N���YS�ȘW���}R��V�`��o�-����~��G��t{?Wv�nZ(�ES��;�_�+��� )��L|��h	,��II��j�����$��]<+��t�G��"�a��-5l����� �N�uD;U�l\�b_��-����U%�\��:���E�wb�ez]��Lv�lf�.Ӷ���6����z	���)h]\}���T'T���v��H��+hK=@̷�(g*�e@BR���n�yGM暨��� E�QF6-*�8����㘍xh���V(:�2�"}$�v5��9���=}
o�l����)�%��ѣ���#�Shp��w;�H�(�9P"����m<Ѵ=k��iqx�P�5y�F�p҈�cr>�D�	��8���5��9-dyb��@zE��6���>yD�a�����՞�gf�ݾ͵���ƉX��c���JS�
;*b\�qza�J�o4�PҖdQr�\dtX?q�E#[G�4A�y5�ewK��-Sm����'�sFm��
|)W]@+���wSId�`�;���Ù�@�r�L0nō�#�j��yK�AN7ծ��ȥKRCG�M]d��yID��G�����hѲIb1�8��J����{Y��)�p"%��o��M*�x��ta��@�u�������ev�
��>#�����m}�Zp� lrq����
)�k�K*��Y���t^���X�|0_�;p���'{��,T?
w����j�ءC�F���w�{�EE2A�+�p��-?+��m�*O:n���B��"���h|l�oGH�	a {�_>�X�X��o�YLx��v� �;[j�SrS�S�������J>�fƂ��Q2�'�p�%K�����r��Z݇�N8�eurXa2m5�=\�[Ks��s&C�I<�Y�k&�|G�IJ�e�C�����l1�|4��	@~�=�c�]��yAlg�OTí��1�)PϹ`�/�a�'�
bk6�j�MZayW����m�Z"�����VC��}[�ٴ42Ƙ��GQ�
}\a}s�N�b>������	,�M��%���Q�ڴ�i?�&��+<�o�V`���wۃ����Q܄������0Y����oFO>����
J�������+�\s�(e	z\���>B��J�V�'1�H@T�TR~OixYpr���x4���^c��'��q�?��0��<}��f*JO��%�&�o�b��j뾜��Y�U�ܤ�Ԏ�B��##�S1I&�׌%����v��o3r��kz��=��oճP�:�V^�%�tZ`Π�Wb�Ǝ@$	`*R����W�e��s��|͊~7	�8�8̓X�
�Mdj[*����R;�]߳ig�ǧY�-CP�?$�Kf�&�A^���۬�q}OT0�>�"'�P���¡���1j��e�o�U�&\��r�}`w���J�������u�7�Wp�+����xۺ�*�F+"=��Vk�&zcl�E�6�A;Q��|,���r��8�[����m<)P�_�ٖ���J��ʤ���,1"�P�I�]��u�����7�$��4� ���7I��&�Ɲk�b��o�����A��ȓ��:[����:VL2�m�+�����xF�_@rfʚ����Jg>��軙�+?��7��3�4\^�$� �ɍ�![��|�ş�N�JR?�+-�v��[p�c8Ţ.�Rd�z�:�] r�@�o��p����|�n|��-I��6Q�A��ݦ!��"�=w_Ȯm�y��ѡ���r�U��o���*�a�K�q����/&�Å����ҍ(xZ��	_<	�#��}iKr,�xd,��h�d��Oq	�b���z�Ky�]pd�<������
|7�BZvs�dp���V�]o���p���E�M�K:���(�"EJ}X*�����5�����ޠD3�i���l�����=Ž6���sX�����pJ���˿���~@~���m�6f ����A�&��TI�"�'��F��i#:S!�x�p���>`д��9kRׁe�-�c��R)��9'�`�L{�[�� �g��R��$���
V`�����ÒKzF�r� J2�"��VR�w�('hpE�v�eOz�FR9��]����M�����e'�K�L6�f��F$m�w�?��H��ڑ����!ѡ��@�A<Ø��Z��N�m�t���[��g��5qBo�湞U(�=Ŧ�\��+��@`IEe׊�wb�醂cC��Mm^�M�@<0(��R{�ζ��x�|P���Qy�gA�"�4�b~��?��85d�X:~���'��t����F
��M���0�VU�aK���e���&MO�EY�<����pG5�����#~�����$a�ws�f�ቘqF�=�@v2k��`�`&�t�@��*�)�߉�ɟj���@g��A6��I���M6`�V�d��7zA9a�M
F��gϢ��N�0�i�Kn ��lˈ��2�L��>rC��w��haQ���'@�˺0\3��m���ڡB�j�n�Y[K\qt<����LO[��>�7@r3����=ӑ�7�o���4z��~i�4�!��������W������1����Uqw�p7�({y���-� �b���;CČo	��-�����~�R2#���@$(b�b ���d�^��cn<��҇�V��\��0�0rT�A�~&K#S��fbA�_O��ϥi8���R���ȫ�8�Q�����  ?���0�U|e���=�@��(�8`����\�&�U�f���(>Y�*F$_�\�_���G���C��t;����߬���[�W�CPD���7�ih5� �深w�9T"{|�0~�����Jl�Qq��4�1�
��G͸|s�`dKH؃��C+@��ިp���c�+�2M�j5���� xh\4P�.o虉ZXˈ|Lwx���ZTޣ9�0m��p�g�	�8��(��6'$��юet�f���ZI���gh�㷀'���2��� �&� ��ȁ�ňG��(cQ#�A���"�+�2��rQ��D�9����b�6ͅ0���H�������Lc?%/K��V�>�TA�1�x�P���_�N�7"*����ٴM�a롕9?t3vd{��xjT�PC��cϧD�0����Ȁ\��j���/��R`�2�D��.)��$}>]Tpɪ��?ྍY����n/�(U_�3�T��~�q��<Ư��CX�9^u&ʎ��w��la�~�#8���(���
[4N'�������idc�/��P�F��.�V �fA[_��`�"���ڏA��Z��99��+�k2�>З;x�����[�5��,�z@��Z�s�KSI����]4�r�C}�j���]3��"lY�r!T�"Pi"r��!Ў�
꼎�J,�j������Ͱ�[��>!��E��Vȑ��ߢ#�ރT��fuv���,��Xz�q�����5��ϻj^�*z�2���	��|��8�	S&����F��Xz6�~	��N�P�t����')�j����Ԕ8�Up�����~W&5���q��=]��?�?A��/������)}yMI��U5�	�r�יF�"�E�y���u`C��K0�����h�� �J�QX5�h�c���6LD�̅���ġ@m���oΑ�oR׆�B$�Ĩ-(R Q�[�t=qH@@��]�ՖښU�� ��6{�T>��zl���4╯���%^9}~�_����"���}$^H�P�-��;l\B�;�|��*A��F�f�8�Cb�'�����W��/�'-�+K��݄T��Ig(R݁n�sw�ƜiFcC��Q|v\M���0Ư�ؘ;���r@���@s������{g�c���w�vt����Î %,���1tq�(g���r�D0����`?�P���A�1N��IC2��)Kz��(��$#��!�"	n��#- �ܼ��H����`�-�%g��:���i�b:(������QN�Nr5@������q��&���k�J,��<�۫�Ӯ#��{W�@��߶F�cg�x�Y}��q4����`��Mu�M�G-PhL(%Ly�N�@�C�BʐV��E����0���l	N�<�g�|[�A��[��Qw=%~zKl�!���ӏ$/����nxv�K�dč��jM�W>����Ue�����&hH���|���؎>�X	�2�I+�凛�Co��$��1�G��lr@<��@��vCT�*<uT6���~"L�c�j\TdJ���X:;����?�'zw���FKOs�y����'�/�v�\�MSټ̾����9�6�
�'\@�:�qWL��r���.�6�����yPjA���W�v�X��=E���@:�/�ԥ��-�NK+�AH�{읉m�L�,�y��$]�����n��x��?�g�z
���u���QJ��*�xJ`�v��^:N
��R�IX@�b�R	�˟K&Y�X*]H|�A�J����[;���2~΅�t�Tz�mI�:�8�s�?���㛟����y!v��sd����z������1�"�!܇��HT�D)i�X�5��˛QI���4L�)g�>&W� ����:u{���@�2fD���)� �ғ�9\�L>]p�x���͵7X���e�7^}�Γm/�����s�WfĨ������8|��9��Uf
�yI��Q$c?���՛��ju6d�ᛘR�&-�*#t~��<�v�4#Q��X�8c�ofs�/N!1ֻH��չ�^ڎ���(�6�[IZ�f�W��;�C*���Hp�Z���a�ِ�7�лO����u��r�ק�ۘ/��<�!½��~u����K����&Yw�Z,kY��8wwG��_��Ҹ�?��@Ni��|� x�MO	��P�At
6�u�Y/@�%�b����J�8��_+��W�Q���&^�7$�R�����4��AL-廩����b��A��wh��Hv�B$���-����J���`<09��:L_��������kr5"t�h4PG�,���U��Y_T�v���G��_���f����tZ�]�7�.|����	��i'�D�D��o��tl�� jŔ���0��)S�t�L}�:��pN e���d��X�àzx�/9�&8f�Ȇyf�H������J�H���8�|����P��@�GZ�� ���[Mp'��C��pJrϘ�]�b]X�����_��3jՃ��P`&��ԫ��Da��|?��9.�ᗛ7@M�_�a�>��\F!{���o��Ɵ4Y�R�u����	�+�����$��N/�nJ�L(v)"u���$5���LZ,r�w�*���n:qQ�i��yƊ�DN1H�Q��/I�ݚ�^p�)��D����9�r�t�$n�\'H��� ��p��5>Ob�u��K<��B?����Ul��`�W1p�E	Wv�-�G�u����jF=�t[�2� x.`C㩛��=�i6s�ǂFAiT�)^uo}�G���B�A��ch��GM��7b���F/���g>\�fMR��?j�ۆM�=�%[I�ά�31	O`���^˵Q�+�X��y	L��)v\���ɭ�P>�����׹a�Ӕz���KX����z�ݕ���	c���6����
.t��������J�zM=@��ݟ��\�~r^�A c�̦�ṿR��둥��<I�ES� (kn�Z� Y�<fX:O+YqK��Ц��%|E��6��G���TI� �ۼ�/ɓ�l��X�>c%)��"�i�K۪����,��=Õ&:uD����ǐ�a�Ǫa��/d�le����n�4g�X�D̑���v���J_�nj#*V,�^>R�߭)[�0�6��³���}1��ߴ
a �4�e�/v��
����ź������pr-?��P�b�J��	��vb�v����#F.�����BO�0���].�d�r�<r��L�ݶo�#N�[�aکKT<@��A�1��:�y?��D�*�&��6{I�zd�N�)k���\ {��/�����$G�^,e���S����!���e�$uu�-��LV��'�1>֓����ݳA�\��L�.�C�Y�E-�=�L��$ډ�]�"֗p��	�9�V^���[�(�cd�d�\W���h�f����-I�gn1���.g�Cyw��U�3���@-e'�Qlr��y�X!��7����5ލw��Ӈ��l�=_��窬��e�N��
5�R3{���������>-}���hͤ���S؀�uf��5(�n}!�OUv���5�V��-S���d+Bi�����M2�ץ���"�5�Z�s�����o#�%�ؓo[��U)9ܞʆa�&�h��͚J,�~/��f?�d��GH�3l�:��I�X���]B�)<�Z�D��J	���~�O�%�#N��񤍮��Z���*t��,V꓅������-�[C�K�v�Mzg��H{�	�rv�X\�C��	=���]\�uN�W�x��"�e�O0U9!���TO�|.�o=��hG��h�_�=h���P��?��L"eՒ��e9!�5�M��-ѱ\{�GN]����u�o��pD��پR��:O�xu�߼Z�ܙ�>�<��Od�N�=�C��x�>w�C0WŶ) b��ή�|H�'*T��XB[r����M͋�MkVaS�	 ���.�&)�I��~0E�M�x����}7�