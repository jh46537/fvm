��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{MEi$ ���ݬ��Bj,����vSl��f����:VT�k�}�N��z��u�T
M
����PQ*Ma�Y�ω������"�� @$���{x��.���\���C���e�o����{�DM�>���Y��/f�'��C�Co.���qEzfC.�Ӥr��s������B_D�N��W����Ƈ1o+�a��ː�k��:G�?0�W<��@��~����;���F���$s&C��*A�9�-ͼ�������b�:�DQ�d��W{Ҏ1�;,�����b��>��C����-�)Wka,Ÿ'�`,ϕ�aWv�F%�s\���lb����ܓ`k��;�8�0T ���q�&�Xc�i(sӁ��!�]ϭ�Ey�S�m_�>�"�\�~)ך͈�y`
��X�o���i֏���^gAlt�&+H"�l$_�=�?Th���D�� =�8����+e^[~3�:�]��<qh�n��E�&n�����qn�]l(�ŏa �s�MW<�3�5��_�?��{�7�� L�CeA>^��(���ueO���r>s��AO̵ڰ�m1b�*�©�~��^�XR}�7E�XC�y��)��\�8�� ED���5�Ӄ��I=��Κ���v֮\2>�x�C��=xy�N�d}q{/�1�������f��-V��K ��J%�༽�<�8��l�{O׶*.��`�D������Wz��&"�� �+?� 0��8�z��s[����)ĵ��a2�����j'�Q׵^p{��mz�k%cy��F��#ϣI}>���.���c���Ѻ�`bƵ'�V��
�����.V� 1�d�֐F19}B-Ut��ݧy�� �f$1n�t[q�e�]�z�ǥ��ӈ��<�8�D�R��
>�g��l��O9�?؍��JCO��aw�ds'�
�T��uT��7�Xh\U�i!:�l�h�&v�4jr��l���>�I���#<���X�F Ε!'���ǃ���f@��q��%��u���/�hm7=�\��wepd�L���/`M@z [�2�U���I����`�� )rƁ�C��So���f��fC/d������8��Yءt�����]�"�1�_p|UF��;���E�ƃMͼ�}�Zy��y�O�ym�j�|��!���T�yL�Y��2?)ؔ3�z�M�Cɶ)� &(q�%��z%�D���̰�7$kƷ���S��/| K�s�
�\��$&:�w����s�;u��|�ꬓ��q�?�䨐�������*�A����$l�-����0�ҽ�bc"US�ezƀd����S�CR���,��hqV�;Z����.�=O7S���b���"�Q���;���p�匔朰��\����A�#{bt�f�Nd4��� 0�G��	q��9��OS	˯W)�qk�/�CT��� X��Q���Y�}.�|9&Z�[+�=��H����d�Eb�2U���D-���Mz~�a碯�ky�ƞ�N��o%���y����}y0��qk�gm�:A��ahh�j�R𦏣�t<�KDF��z~�^қ>���v�,��>�������<�Hl���;��ɬ*Į���u�97֧Ů��2ʕ���Xgե�J���"M�k}6(��� nۺ��Q��R���3+t	�5�BE_N�`k�.5�"4Zj�8�*�(굚ڼ3��
{s���5�D.���u{�/�p�dC)dZ����|�y9�C��C�k�lq��T'���D���������Gy��S��Hy� %�-���&!l��]�siq����]h6�O��%#M^H� �bT��n��N�2O�8��e�:L��O�t;�W�pE��ٽ`� �r��YB���9��w�`2U�$�7��?@Ik�f�MH�n.�MpA��� @)��y��C�y$���4@��T6j��_t?P
V�]��7V���B�X��e@��:+����aź�$����3�-z>� �HS;h8�x���՛���)d����R�{Y��>?�?����ٖ'�xJ\�(��#��J�����4�l�"�ZtjDz�/nc�+������@�ȑ[c�l1��o��?=��%��i�;̵���g�� �M*�=�S���V�Ē�q�Axw��`\����2,����H��{��/��OZ(�������",L,c�!]S���\{�ڒ�K����VI�k�8��Ps��4-`}
7`?�l�j�@���Jȭ#�CJ����~C��e�6@
�&ٴrpM3�P 4p�Wa�[��܌S�D{�'��(DZ�h����3���3g(������3��T�Y~'�d�r
AB�P��$��֒�'XԦ«������;��zB��z׵��<�׿Nw�;��e�����f�Eh�#@��K"��պ�QP]������3wҥ��!��"�n� W�k3s��Z�g�vLaW��\%�G0�x*��@��{�,�H�½.�s��K�� �vn��gߚ���09?\�7����#�jPZ
ƅ�)NO�#[�p�~�p�ఀz�S�W�͂G ϴ,�@�U�) W�Vƅ5`+��@~������	R��f/��N�;y��!fx�ë����������M�bM�.UO�fƟ%q�6=w�ʶѕ��V���\L���:��$�;{jM��[A����Ƒ�RĒ�+��8m�3�6���-8�	-kh�3���� O���|R��R_e|t��}���3�����ȋ�}�	��B���jɢ�^��V