��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}����W�![��J�n��=���_�*�?&	i̎�.��e����J{U�8o��k����"�F�s3�C(�m������+9�2�&^�[�xFuk�c�������-���F������ŞO�u�?�n�Ӫv8$���b	y�M8��!W�63�j`m
�>��Rx�Q<��Oȡ�L�ЖNf4�T NRə*8bf���JS;�:qڔu�Q�H���F)��z_�����%�U�8:!*�h��	n6.��M��^I� �)NU�0�~�yc�.F�C����}����^҆4n1����[�lP/�a�0�mAi\�Y��(�P4H���m�=)`B5�ʠ'���*�>o�xz@������r�dk�Π�h{�5B�:���F_?Ȑ�Z�44�=�G���l�u~L���l^.����@V�0�Q���S�df��-��柁x:v`�<-�w�<���fl��v�b�]�� G��
������ӧ��ǣ`��f���i��?�V���L${��p|.��*��Ie��-�W����
��y|��B ���{�]��h(6�(z�d'�me�9iUdڨ�gDE
��zWE��xb��<q��n��B��55���}�ŧ�Tg}Z�ܫʛt�E��8qs�R�J07R�8FN����C^>��|���9'����@'U#m�8����r��	��x��w2�Azt��%90��dsix'z���]����);�^c��[yp�,3� ��"�LTT?j�L�@Z~���q0GKU�޵��`�U�~*?�RR�����\�W;io��3�݄�s�A�&�����������/yAG�}��^�w�H������i��g.ܸ(�֭�7�s�>�c����/�GT1d[x5r�Kaᘏo�4^�l�~�+�sIvj�q
�N/��<;�F�z�/ߨ��;:���ˊGp[�F�)�(-����*�G�U
g�n6�^�HEf8K����-W^��rct�d��N6 _���ԕ<P]~��7�p΂��91y�R8�~�)��6ވ-U�{UDg�Pڮï��tʴ�҃�M��ƈ�����#��{��;�&T�
"ܙ��H�"�O���$jF���jrO_��iw<8�1�O���w��� ��$��5J�?�dO��n�I��,b���/Bv�N���H/ݻ���u�(�K;u�{,Jr�QQ��L��8��7�?��G��V�?��*9�ZXe��F9!����_B���t��z��y�В�$��'��	L���^C����O+��[�YJӢ�g`:!s1�zXջI�'��t���=k�-�*�'.����2(5u4�M�V2L��I{�(&(~��v^^��̐��_Y��'�"Ta��Ћ^�/�u�A"x[�ٰ��#^Yh�ń�;���%��ϳ���O�L�����|b]��� �ww��`�Fee�E%n�0������Nel6�ڈS�������v�8(�n�V���e����Dtz���3a�'��w�_ JJe��նgb�*�x�o����;��a}�|6%�bB��G���cv�T����Oky���n����͓V�[�U���Ul�����D�.�}.y�#�q�y���zAF�ƌ�u�	��搜	��&�z��>Q�G	��s�ɜ9*M��ˮU�J���p�y��N�L�g�<_@Au�m8\���!7���=k���z��1ARD�3��j�Ś��]稞�Gy]k�9���������H���+�J�W_���:�W������+��}�/9�W��s�ؙ���?dDW����)��ZSl��ݨv�gg�2�+��ݙ��YC܆���ILzM�<M�h�M,�W�Z�n*�<]���g�;�Sm��?U	�d�� `�eFiN!&}1�v1�g�����mF�y�·���T�@"#����?��C&�0RJ^_��~�(I"����s6�v��ȚM��u��J,w�D@��\��^وB�$7m��,��+�7ޑ�D��]2�>�� �:)�.�0}lU��I���41�İZ8�:;.a(���m�N�3��X̑�_xY<�C�9�@3��?H�� 8`�g$�xc�EɅ�%�8AN�o�GBwt�"h5�ѥJTb�U��o]A��L�l��,#zK�gB�܁���Y菠��1��$���������n]�Z��?ůw��ciwE������G��3�i����u�� �d�h��II���O��+�bj�%�!$k�6�ݫ+��� ��S��!Z�Cm��Q�p�8Z�W����+}�{�ȴUH2�RFA�.�,�H	eZ���֐����(x��D�s���Zp��w� ?��Uv��)�5a��V��xa##vsζ&�(޷����W�pz�'�ʆ�e�;��A��B���B�GY��PD��J$��Ί���YC�x���[T��gR�J5'T0?-[�P� �.�6I��ߛ]�g�r��o�j�DC�L/�����Tj��� ��Kn �:��oJ�e�ܪ�n�E����<�1jq������\+�A2bUi�Y�"BE��5��`�#-�fz��Lw�����B��V�ZɊ�v\1U��o��cy�ݲ^�Z}�UW{�Bl�+�B�G�f��`��K�| �h���ut�\~礈�����_2��a��5uD��,4'�.o���r����ܒ�&��_H�IG>)21]���W�+���u�8m���\���q�����eRbA�����̳���{�
���d��;�=)�|��M�ǒ�s�ᱍwH�Bd�I��N��	e5j��o�t��;�O&�=`륃<bV�u��?0i�L��!ҭ�b���K�����^~+��e�y��`�1<�y'�b���Y�Epb��M���t���X&T&��)P�1�Ze�E3�zO&����_�0���G~Wh�-��%�*p�at�	_�L8��tᏑ^֤�3t��ZW���'Y�1Ը�'*2E��^�Ĉ����g�|,�7��K���{r4"��('�����/�Zﰆ�&�t$�|�N����¢0�z��1��+�f���,Ceo]e�q�*Jug�'������y�@E箿�O/D�q+�z�h�G�A��9yk*N1��b�?��>/t�*<���12ŭ
�©�{�����;Z����1�W<�����n*�m~���p�"·��
DTt��-�%x�B/ATq(\�Ni_�kv�3k���:i�@���_}�J��2`-�l�Ɵ�r�a��g+�RaQ#���g����#㢗gL2�D����p��D��7K^BPO���X,�=,�Y��߈��^���p[�r�R����z��(��6:�Z��RC�Z�7�*ь�5�'�ۙm_&2����sAI�AWw����b�.&q�����ؒ��04���۔*��.s6�54�+�0y�]]''�M J4��ˬ����X9v	8���@fŇ�*��%;�j�áNr̫�2���5�,�i?u'=�Z1���)����)۫�W�CCX�N\~�F� a��9��������y��)')*��jF�w����è����}���J@A���Tg��W��b�E�Ԏ6eWՆes0�IK�C�������#�?��7d�6�X�MiG�0w�n�Ge�������m3��/~H&7�d��#��pF�Gr�^I,�0̅\��f�8��j���b��-�U��/�r!M$�Ôt���[r�?,nNC��h�<�٣�Qw�n��1�GJk�Dq6�"��=N1>�����M��Z�a/44T��Z��C� 8%�H������"�v�p͑�+��U���.�
~�W�*o��!������Q�� e~�4��4����d�A�����\xdQ�)0��l��a�ЦˆۚǮ�H6:��\�n/38ch�{� �5�'��O��z��P�r��O���T�V�0ݢ�<��8�+�NJ��%+p�@}��}��ei���.P������K�U�0��c����=���0�>^áM�����S�䳼^^��mM�Y���w�/���ᓚ��Tܓ��aHu�8zyd?������Y�8�5xr ��e|:,Yi�C�4��2g	9�L~���K��9�7�Ģ2����t��hxI3����JBr��o��f�jO�� ����<	�lW�wb���,��a{�B�4n���7��/z�����t2}Y�w���u�<S=z�䑮��
�Wt���c`�JN�y��%� Ic�L� JW���kW+%?�?3P]�.Mx����*�ғ8z�V�aǇ8�M�KN�lВ��Y+=�{q���a�縐���(��]��v�Rf"�^��и�l�	;�v�gX�j�S��zP��.d��-���4,�>f�qu�	m��!��]�Q�7L�x.�� �V��.��N��a�*w�x�?�!�� !��!�H-fR�O:3��(Qc�q��^����/'.�y�z�Q�j��@Su��r�w�{Nu�=�DK�.���m�~2�Lm��������W;�R�	5쎱�T����-]�҄�m������&����=�j�TD�F~�L,����-��i�����Ng���Lj_����Zh̷�*tT+�t��]��;��r��ݙ��Bs��N$]��Vj}��X������}z�\*�����]�R�(�L#�Su�D�����C�TjX�I���yZN���H�3^3[�g�,]_��	�b��*�m�,��� �m-��۞J�t8�^�D|��z8A��G$)h�;m,iBs]m���<�E<
�:��6yE ��M9��E>?JW�+�����(Ԃ^�M�|ҰS�*�1��>�<}��y�9غ?5f`���B�z�I$�
o��*�M����t�ޡ�`��7:�I�3��=cz7�����m��5J3����;�b�U�G"s_�4I�޹�Zg5���,��ݝ_
���Hj�i�/M�aަ[�1�M�]����Z| 6ǯ5ch�x2 U�������V�Cʤ�3��ν]���[���W��Ԝc�Q<<� ���u�q��2u�-��r��\{"Ԭғ�[WC�Ѩ�W�V��,0xz��0��7���By'�YV�R����@����p����(���0P0�!{���AB̎�����1� 7Ƒé���u_'���V�JK��T�3�����ށ�����d���l6ܶ��8�6mЕ�3�!yo�R�𽜒4�W�[���FD7�֥J�@!(k��q"���L��S$�As\�Z���`ER\A ��_�s���d�@�ǥ"�J}���a
�Ō|l�p:�k
i�2�h"{���f��3�5M��3��\��Ѫ:������k�qx�@���!��x�XQ#>�L�Rg)>Gn��՗UT��A��@���p43������ɰ����-Նc��16��@�A��f�|t��cU��qq	�$�گzm�fҺ��|���ms[��_��/l8��u"S"5��`W|���.F������?_�S�C�9�(|R��~ƌ���U-\:��C�����T���T�kb�d�����}���4��ܻ�o��ʌh��ܾ�����tRsY���TI+{�u�^ꯖ��o/8�b��*炏�N񿻢�ԡ��hvc#���92�ɠo�Y�����f��1�$S��P�� �b�6B�7ӟo�*�ߎ��K�\@�Bc��%���>����Hfɿ������������"�̩y���9H_�Ʀ��9�Oi��4_�I^�c\kc2�i$A*�=>:h�~�KŜf�e}������.�oo����C�-t�ɉ���u�����燐��1�'�@=��zS��J�_�K�g/sJn
� j��S͜Fi{�q�7�PA�e��8SsH�Y�j"��*���=��H�{����$��9G�l^�1�6��ݧ荢Ps�JP����R[KǥƲ�Ǎ�s&pr��5��_t��c�gD_�G	E2I|?3x(rB����% +��	�F-냪XQ�4H�ʈ$�d�5ђ����Lzb��?��k?�]�RQ�NF7*���@2���ڱ5=R�N��-A�1df��&sߑ���#�}w�V� }v>K!�t������<	\:���YgH��	��W��tL~��lC�V����Ѥʁ�Ғ,����z��r(�����G�����:��1�M��To9��%��	���떾���<�u��^g���g1��zd�y�>�E������� ~��>��0��՞_6:��|
��$T̠?`�/����!��*��hE���-, �q2%8t9����C��\Q�H����su��=DОDu��D�A����\Bܝ�>���nw~LR�r�^��m*|5CPBvN�iP��p��h�G���`���&hu��������T��Z�>���ˢ0c@�	}���p���Rq��[|���c?�Xx��_�ZB�slv_Y��K�.Q���F����l���G��̦��6�R�B�ڙ�LQT��E2%����
^QH���`7pK�zʳ�N�� �$�fl�k����̀�Տ��>�ʋ��D��ױc�c�W.ec���V�O��j�do1>��,:��a�2�)�����E�t��r��_(�00캀��`S�r�[Qr+2٢ '!9���!����� m������5yi{���e� ��f7�f�E+[���a�̇��:�h��#IU�{���;U�{=�c. u��ϐ�{�~�Ʀx����q���]S�_P|LU������3��D����y�+Ņ���Qy�G{9cN4F/��C��'r�ש�#���C��SW����YY{��W�s���������sZ8� o��C��jߝ` �΂��<C���>ݷ�	�C�8�b����٦��E��?f=q��'^���a7��ȳA�1�M6��GvvT�t=��_Vj$m ��.A;ж��p!0��p�?kT���|�.��2�>-��ȫ]��K���2�ؽ������j��d ��4���耟z���	| 9���e�0:�|��r6̠h������K���`�3��|r�e��3� ��_���u6�E:U���S����̜Ӽ���Xpg�)��t�i�&�'��ū\x�o����{���y�)g�aҞ��&R�Sg��U��";����2�1�,!2��0�;���%����d&�z��3����Z��53