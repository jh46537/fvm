��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�ӿ�J���I43n�l�Yt���U5
�
הH,�Kȑr*d�
+��ѐ� 9���?�#��i����b���0�Qj�Wl�P�s rk�����a(��-9��1�����݂�8�aS���W���2Y(�Q�٭Ȉ,H�x������cq7N�����&E���P*��>�Hm��H�^H�2s��Ԉ�� �w���~s��d��,8�g;�+փ)U�%��eS|���㙫�廨x��l�[A�,�lHm��vޓҺ�椨g�$
�+��h�0�V�"��ވq(uQ�#�'U~��UL��F��o��(�R&��F��+	�&��VK�@�=}Fc���|��yh|����"���&�\\���-O!s�G?`�1��]7:�J��J'���x�X��(�-��}��c�;��9~�?��a�I�w\:�7g0�rS����J	��%wW�b��=*��w��l����.�����CB$;����v$������-�,u��!��B���2�E��q'�ӽ�*�O��'�B�����N�a��I֧��g>B�x���v�/�}��0��:�fxB�g?��p�.ŕs�]��q��n���B�At�$�+,@�<7_���*�>�������Zf(��߯�x�.c\jhxG5]�Q!.����v��� 2�V�|Pmi	�	L�������4X����]�$�:Iǯ^[<x��;>x<��fm�Hk-�\��QԠBG`�!������J5s�Rze�	%���b�zB|�c'R�4Rwˤ\p}�q��?s'��u[Y�xV�"��ڇX�EK\Cј�H��{qn� �>��	���No;
�Z7�0����־Xnp�s<]��:>�@���\h����3%��{�&l��C��� �Ә+�X{��"�&
�8���m ;~����x����.�{^RJ�����r���>L�VLP���N��n���{Yr�!q�}#VJķtg-�IAlE�l�娤�Bj?���]�Pl�Z_�w�� sk#2�(3�Zt0��)KAv����p�ۛ��ʩ�*a靴<�v�}�����C��4LTo��pZ9�h�}�Z��D��`lpZԙw��pv
CZ|�2�8v]�W�+.��P�M�8͛��s�F�GHVd�g1D��"M�\�XM(Z�
Ľ�Y �U�rt�2��j@���Ғ�5��v�p	u1���H�]�b�
�J�M��U��LF�+����$��>�ӟE��nP}�����#:�qU���M6z�$D��1l:ez�Y��]�Ԛ���h	8�w+�����Y<6�P���ӂ�mw���jK�.�f�ˬᾠ&x4�u�JNz��se��'��a������<rpÎ�61��%�;s�V��ǜ�w@-&R�VCJ���o��{8�	��tL�RgY�%">J����e�~#U�GZ�W��xE�x܇��;���r�`-��r��0�~�~���)��A�p(,����q�j����h�HJMMY�US�m�naoh����A�;��%�i��ɿ�Y=���g���R�����j&&���5�� ��.{�ڵj]��Q���գ�}����@[��HX�˯�p�����4.�24�kz�+����
Ql8�ǼP�:�{�67�i"��R����5�8=���v����[��'T�hU9p�lAy���C�z�ܧ|��]yqk!�:ZC�2VW��4&T`M���v,�����&}����! ���G����@�ǥ8ɤ
�m�hT���Χ3�ku]d��_,E�*7BdH�쌋G-�6< ��A�AeA*�?Ƚ�Bd�Xy�2LC-'X�����O3S�&�.#7����d\a4>G���q�+�|cN{ �x,�)#,�f ,�1[k;H?��d�-!����R�r�D��!��E������|;�ǃ�|���I��y�X����#�|1CD��fdX�xZ̤u��r֌�����a���&��<0��L"�/F��f�C���pb��d��j?.\�R5r�,�|���0����+��K���Hw�y���L�Q8�\���z�����
��i5��ˋͲ�!�Y������k�c�.ܱ~u��#3���
����Y���
�J��u�lU�b ��8$�U���!��'��uv�.���c����ܧ����a������A�Q،*#�qd��z�}���%����I�>�"�����}�h`L�U�ݻt�n!����ڲ�V�R`�H`Q�x����f`���@�H']LK����"�ǱL���q�Ze=@@��i[)����cv�e��=D{շ~���X������ũ��~��'���?�$s�D��	��=�@ӵ7���wV��ߘ�wj�7,�v`�<�.������#���H�d��7>�VC��T���q�Фjv���RH�p�Hx>Z,�$*��5�*�Ü���'�
Hȱ;�:q� ��1m/:�7���>����n��7��+i�{�v�N}�`=,+�H �'�t"bY�L�w�D�n�8�<���ж��.�-~֚�C�Y!v��(އY�뗏���L�( �ps�;S���GeD	po�ys�.K��cAh�
-���٢+\�ϓ[�xeƳN�AŜ3&�%�7�B�i�m�9�r����
|���Q�R��?C�Q��r�9�L�OY|�3�zW��Z�H*&�:�Å�;{��=����AY:�^�����k�1~%�Dnh�®g������%r>TA����u:���c�,�.\9����O�膓E�9G���=�,�[�/9^��a?����MR��3�T�gW����
~F�B��O�JGt��Tl�{�\˚��X.?HF/Uֆ=�J�n?Z�+����{�f�,k�u�*1�S��,�Sg�(����f$�ΧƐRk6���œ���/b�'�RO�܃�n��� �Y�F�lF��Wr43�t�� fd���|Υ�c�?���YXu�Z�����N�ޅQ{��+&� )���Ə��r
ҽX� ��Tx�ȩOf���ֲ�x�~���Pf#/Ho�d��pj���@ .:;մ2���wsݞ��E�l[�CP��qطn|�v&��SϬ�����R�����<�5ݏ9g��&U]܋g��S%�N�Dx|�[�cu4z���_�!�ů9�>�#k�oͻ�+�-�k������8���A0.�P�&�+��O�����NsyָnA�&�5z�TpBM�G�Y�Co�)1ڟo�
�R����g-�W�|�sҜH��-z��fL�!��W�&-A|��l���wVl�F��Ǻ+C�7���si��KR���}�U��%Eιe��S_ ,b��CJZ�g��@j,�5�������aK%���ô<$iC.i����]e� q����r�ʍR1��{��K��ux4O������qu����q��p�l;[,����J���2l���+Z3��~�-└�>�֣sbݪL@Dm\��&]���OS�4���`�]A�� ����o�D?C`7^�C�Z?��۲æ�K�}���/O�	�S�B�M�����*�P�#�V̐��k�n@ ����M��U)�C��	���dk�Oc_� �	�T�wj}���=��`ėpU�ui/�=z�!���Hh��}ʺ�dZtMf��Y��}c�+���T:��z��ᣔ,�N&.׾�>Eì��ѥ��ݢ�:?��6C���5yЇg?���|�p����ߓ���I�F,��k>_���T_\PbI]o&�&;T(�a��`���l�y=i��'���9Alb�"�E����*fc�������ߓ*n�:���7{�C���,��
[91��"	N��q�u��
���:O����j��v�C�0�h���Y`/��̀G�/yJ�u�:q	j���[J;xw��=�{lVMp&=��U���%��,KIj~���'|"Rd螡��R��`�v/aM&B:2�HR�j�Mn����~�1�!��iOۥe�TQ��!Ȋ�79I���:}�N�MC�1�W4>4�1f=`�k��������5�-�%\#W�Md��6���1T�$��"]��J"]�^�.�o$��;�����Zլ��&}b��=��f�Vg9�!tS�i�F�?|[���R�: �(�%j5/J�1�,���q�^I�DL/�q�@ͼK�=�����jCF`��_��3?uW�!��V����9��O��y'������t�)޶u4��H��r�}t��p�$K�&;H��4N�8���Ţ��]#K�g�t�S�9=eQ��51�،�ô���J���]Ҷ��}Sz j#�"�i�6'yp