��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�c���G�J�,=N�{�P.�*�@�&��^[��Ԇ�Ă�#�a��� u!��;*ջ�2��n��:#7��l��8����k�D��"3rd+���]��*�a���7�a�W�Ce�L������ ��5u���#��)�g���=!5�g]4�y��t�/�Y��Kw"������u�J�M&
Rܾ�a=�;�D�.[9>��_2�j)���&��%O���b�R#([��%x�E��8[���i��xh Z�ulN�"m*��5ߡ��!���ʛ(k���=���&�}�n	�i��8�=�(=��>چ�����[��/��#�qĪ�7�������m�훓((IF�YZy�r�z}G,mJ��&���\�}ֲ�n��i���*u#R�c� �zP�Lr�U��]o���� J���Y�\�J��_ա叫�#�/��1��":0jO]�T�F~���?r�c$,����Ti�o^��f���eq�d��U[/���s������h~ߌ�o'�%v�j9���sY����2D� -�'%��Sn��x���}{<
��i���y�+N�i��.�w)B����&�`�ܜ�ۮdA��@���԰g�TF[ņ�Z�W�y��t�3�����jC��� �Ջ����4��S�/s�w�,��b��u�ƶ�>��ґtչ�J���F%��j���`���C�3	��@A�#��|���H�E̚n�s�ワ3.���lrӂ�|Q~�]��]�\!��F0�݁ʃ���Z5�;.Aw�� q���p� V�N#���m�R��6���~���R�t���[�0R�Z�aK&.�>����?f����!?��$:a'�/)�P�~w�@��z�G�g	9a�8�F�!Y����U6�<��#������ş�Y��Gٍ2-F0��eJ���XݓJ�a��dgT������� ��1�!z,�g�
�"��2��1�|�kOEV�TZ��e&S[��n�S��� �d@\�E�3����&w̜E����+^A�9,�)��������.T�^5N��8j��{:/����
�d^��U��N{�{��ҩ��I��Rǀ$Ɯ!�M�b!��~��
��Wy?�g�����[��)���lj]�.f�Q�������(AD"�d�*D5��v��rv��+����B���v��թ��� ��)���9�åCC�!��JfU�%�.1�`����nNf3�Ʉi�=���kH�� ���U��%`
e�R�} v�~Ǐ6��dq��wΤt���.υ���֣���gIM�B�r���I��|��]��0̾F����4r���>�������LS�.��@��NY\��`����0�{6��L/��QJ��uv D���&��8�8Hڑ�%�
)Xףּ۽�搬�A�6�:3��$��џ�ʀ��Ov:m)H��,M�:�Ι*�~/����!���CQ�����c�|.l�����1	!Zy�r��DE7���r]�\�"}E�Rˡ�K�#9	HP��Q`w��78=G�G��+u{��i��p?�6U�E+�&|KJ���6���pշ}G��>fc�f����m�+�z���j�b��A��D܆� 55� |��M��t���a��>�K�h�[Ed�*�DO�Q�����8��6�9�[�s��"`t1�є]e�aC-����81�t{�^JM��� �t��C� D �H�j��\�\4g��KP�E�'�X�J՟:8+�N�D��Z�r)��8����]u�-AEW#�^�6+cHx��N߲k�968;OR2n�*)�q�3�<�����$*����	�np�_�=[���AF�~rC��sƹjBjB�Vn�*b�)� +���¯w�/D�b�����H;sh,�}2L>�;�ȩ����̵U��y`�q�L�{�aͼ)j�+��A{3T��ſ7=��)(�e]l%�2�wt�~L�xq/Lo���(<�d�y��'�gP*��K�h����y1��������"�|t��vC���J���WqE��N��#d�I�#(�4���6��=U�+��T���aE�s��bw�]�T(��S_�M��"^'����Ѓ�bP[xኤ�zװ�/�,U�5�w�D$�CG�Y�ƕy�< p-
=�;cJ��gI�Y��q3��IA*�8t~���"�6,0���6�e��!�ka.=ZHv��5Щ^���J�pp���>*���XeQ����d.�4X�߉�Z��5J��U	���K����Ē_V��G �07J{�BpH��p~J��P���bQSP�2C!����z��$C]*�[gD?��ڋ�(�pn۾���������B=��b_�-���G�\Z����=y��̻��X���S���	��l�c�F���c�t����o�ב����h6?�[3�A�UYT�n����W��KH�)]���p:�nE��Ԣ�I�����]�⠬_J_`�Ēg���A���F@8��ڝQ��Ȕ�4�9�zz �6-��It�`�F��牤������b_kIPh�N�����k���X���-��z��s�zn�B�Oo1�d]�|{�Us@�j)T�0�(���T�YKMI��n�2c(8��D{e2e`y�.,�����(�ovr���ђ��pO�v�h���6{p���`�����m+Ա�o�� ���h�9�#��-�=N\U�fo��EG�2[1�;���nڲ�UX���ZA�ct������n��	��)������OFߞ�
ҝ�d!�s:|�~�W���s�O_����})����_�7R����E�d,�c��3��F�{��P�{������'|r��s0����ߩ���k�>��7}B�pu�p4�J�&A3���)Q��ILѲO�,�kc�Y����8���Ƴ��wb�m�� �F¡A�S����u=�O��
�z'��?W:�:�'s\2O3`�C���D=>��1?&V�&�'��lL��5��$}���D��$���w.{7S!"Ec����KI�Hk*r~�R��Y�������Dḅ�b|�����n^?(��C�0ݙ�t��Q�N2��
�'r*۱0S�	���HA����|��'����������G���y�ౝ-��� ���N�Y��n~-&�z�h�gp���1`˄�����)�A)�19�K��6J�K;~�[��9Z��Eu��x�(m��[��4�� ���X}�,�;�p�Zl�n��F��c��8�yt8vކlى�Uv�p6O���pH��RߦǍdr��>��W��DU�����v%��e��_h��`�#�nҨ_��*+}��i���Y�s�x���fzʝ���W �^��"���=��;i�zc��hP���h��?����������=wF4����W
X�.���3X�s0��2O���h�����K�P�&\��%JkbY5�CX����;^�7Fm
.����jw(T���@`q?��#���f�l��|	��d�譮;����]ʌ훌ęO\�8��g+���G@������L|�>6��#��*uCoqP��-_N� �{���C�
W&��Rϕ��[�c��zU������=�B�N3�u!S���\b�U�4�RƘiZ�r����Q]'�$O����������x|� �3�� %$w�HG�U5"��`��H�l�Ű�T!�H-6<� �|T���kk��%e��\��
F����q��vY�KJ�*n��t;�e>�d�[��E�>���"��w�s���Ur�}���#���d"�y!OUc�넽&p���<5����������6���L��L�� =��R�jj��=�#�8�._%��t�r۞��%�x_����|�kZC?uo����9pH���`�'�Tׂn� ��H���ևz���������������	�jO�I���&)`�9��I�?��=�6"n�h��M�Nn���VO��N�0�BesQ+ق�t�8�0�Y~���VKF�%�K2����6O���NM\~}7-P=�[��Vs����U*D�~��J���$|c4w�Jb��+X�|Q Vi�z�jQ�u��B����B8d�;	%��/�`-�}${�/���%u�_�W���S�j}bg�d]��2��i�Z��x*;i�+\Æ�w�yK�-K?j�R3.��}-(�;"����/�SW2~�^IPwHU<��6�&v��b+��r$��I�0l�v����?3~�k|�y3V�����$Xjv���?YG�"lr5�N�6i>mZ�\6��#�~�I�\@��5�k��t��@�f.�,>�t�ͪ�ޟ*G_�� �k�?ith ����٪��r�\� t^)F�g-Q������;����6�?/�����q;PŔ�������>KY5�!'�TJ5$\e�� ��3��ֹ�O~�tA�
���G�Aϗ��9��������3�d3��W����-�4h=\�2y��#;X-���1 Q��%�R_����?�&�1,�npx�6ŏ�Q�z�4��z����J��S3�]����b��#m�[�]WWΟn�߯6����{�~8��� �,�*�w*�4�p��Y)Ť���;�G�`vW�O��x���,�(��Ns�8>���~��.�Q<`ԙJ����S�5���k�p��V���(^2>��� 8(�_�E�w�:����ݿ.�:��pS�f<���(^ ��Ҵ�����ai�vʿqB㴿|W�~hO��nFO�ć�	;+�5��i,�Qė��V :����t+��~�菝fPM�uZܫ��%��h>	?k!�ql����A7Q�|����ov���zx=�����l�| ��1��k��__s�P%"�O���m��Au�b��:|�+[[���[�o�2�ˊ9HF�=���n�>����x��w����2��b��l��2��;�D
Go��X��}���e�^�EH�c�Fޚ��|�姚�qTGYZ7��˹�+�'�|�I?�B%�_}$0���~����װ�F>���
R�V014Vr�̃��hgPE����ﯥΤ�nWm8[��3-�2�
z���c�E�-g$ 4�����0ԯ\��UhG���=��ИG��G�Z+�eѭ�h���N�ٮ���^=�q)\?�$Ū�6T��K�*ڋT�P@wB�����ڣ�nֱ��M��L�]����\�(CY��g���t�_;.6o��f�q�����G�*0�q�@����U9�އ�E�� ��Y݇���W����k�qmY�,d<�v�j��_(�zE)�xRTw"��:����U~���?�Ѯ��YERQp��.�	�%��n)�7�e�+ɒ.���@��E�mb̜���~G�7�}L<N%8ah�#��G/j���m����4B�ni'�ʘD�}�agd�V��oƾ� �X4��5�	A6����&l��!T����3��Q��D�˶û�N�U�U;��/�1�̬k`�J���눭R�/��Hy?�Z�\4�g��H�9���B�p]l�cfCe V�~AW+�b�SҌ�"��9}�P����kZ�_Gr�
����{4p�p0N�b�
��y�$7vY�	R��P�K)>�L��\�W���<Ǧ�
�b5U�}~ؓ�Hz���BW;V�M_7
���J�k��
E�2N�I�k@8�\�;pN������s��ǆ��(��Di�аG�`�M�){�7u��R;�5ٻ�?ą=�mq#J����^l�O�^꿎��+8���?q���Q�1�q�2���p�jVEw�(�+�خ��=o�WڒAh��D'2���*�������E�w����X,�bʮѽ��%��%m�;{��ԲL��0�ؚ;�OȖQ$����t�4��A�W�SQ�W��*`�H��K��r/P�l+,��S���BA�^?���Y��Ft~ó�Ujn��E��v/"Gt7U��'@���J��rxjT�������<\5e7��vge����3b�l�`GZl�R�d)D�jiw��SA�&J�<��a=�3>��c����{L䫳6�j��}C�O����7�ߞ��Ԛ3I�hE����T5����Jy�3<.%D�?p�g0�c�t������=-�e�8j��1���~�j��R�=���nɝ�1���0�����H���}��/���-o��hy�"����<�Mz��h�1���Q�'��;���m�6|��EZ�[A�業�ݟ{�X��@���Z�@��l��$\���
7�8�D9x��]��� �n�	�z:��<�`�� �n �Q`��I�9B?u�S��^M�wu��k �m]��n���J�ܬT뗮���45Q�@�&�v��D`Oe�l����z{��y�H� I�D�_��`�L�%�_��M8��!x��+���q`5l�����
jNo��KD<Ga�1��F�/ߒL�����)?S�j Ii����i��E�d���j��l�k�S��euLZ�y����k]�` �&+yi��5s��ᖢ�Zi��Wm��N��s8�k7>qcL����(ǃE6�i�~`��ȼm��%���Z���1H���Jo�Fk�F֠��5�l/lf��%�t+Q��"��6
�̍���RY��������M�14_[�3��5-�~�JWR��5���2��\�!�3��"�#f`�􅑶$�Ζ:�-�@So���褢�5�4l~K�e�����	�Λ�/���[�_��(0���Z�6��!�܏�x��3�aCBj�y7$#�ۈ+�a�x���X�P'JQD��m&��j���F��������$=�-vM0+�