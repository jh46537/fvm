��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� �� R͝���c�	���)es"[��é�#�‍?t���4�5!S�TP��k�$��  ��y�྄ !۶��Xe���a2"��Y�������-�ރY���x��$HDA���)k��'� nA�4TM�w�3M�G��`Zß��(^����G�ŧ ��sMT�ġ�8&�F_t�3!%�)o��(�
�Z�g"K�z����&F��Z2��G��E����H��J�,����2�V��Z,���"������+uP��1Žɥ����vm#pI#��7��Ѷ��F,6��+˸�\V�3�9������̦�Xk���Q�F|\閮^��eN.��8;�F��d�D�C�W��2��N�4�\$��y�]Q�cEN#��s���$��sO�GIF�c�U���������?TJ>�*�[�>:@����KN~�#��{���X��S��N�[	�Ó��ލ��(���~��$@*d����U���<E.1!�3��a �`X
�*��&.��F�/ Ƽ�J��Q\= ��%E�H��R�W��@��h>�CB�O��;�"��^ϼ��NI�y",$~�[>e^��V�q�-�������D�(FG4��11q�5���S��+�ҳ��`�mV�VQ�66q:7�aBO�؝;�7/�T�ۯ�T�rA��%�Z6v �S��j��gj��9Y��w�*�szA��l�|G����ݢ9B-*@i�^Fl=�@�+�/X�����*FW`R�f�k=��B�o�(��S[��d!`]g����a�uo��;�)gcފ��Шa�Z�Gs#	T�@}��3ژ��
6Եvm>�]a⟷
�?�T�s�w���l�����O����S�	�s�x������!'���}\a�,3����`"����r?�dNF~���R}�̯dA�:0_�(@x؋Λvtu����\�f���mJ�fp�8��r�ΡuEy��P�v�L��&��&R�F�;�
p�/�{IG��E���I�\�F���FirJ�x��('��	����L�1~Ҹ���i�Uq���Ѱ�l��� ��TğWUP���z�7~ۆ������E�Ӹ�(��z�ј��[Be-Q��F�`,6�@,il�崔6bhro	�9c\�m!�U����J���xn0��i��i7�r^8{}��Wa5�,��Ex8#Wn6tѧz0be5.p�����Sa��AO�&�X6�Y�=*	x����y�ˀ<�Z`�)ϕ�6��)�X_�|���~�2���b�(1��FaS�bP�s:�RqbU��-&n?v����������I)�LsD�^Y�2܊f�J�I\�U2T�Ԅů������o��ap^�=?\H`L��ڰ9�E�m�t�� �-P� �+��;n �h��:MƗ�����up1�SDR���J:�I���1t�����-�Jwܒ��x��5{����
�����ґ9�M����@�x��k))��rTK/��L|	ӆIC��d:5�b�������o��~Y��G��k��0@�[��W��C8�y�?>̙$փ�i�	��ou��XR�A&h�����b��ٗ)_�����r�|��5h��x~�}�(��"�.����SH����	P�CJۭ٭b�p��i��%H�7�-8��i2�bAb�˛�(����Q����KQ��f��3�T�
��(��QGt��%ٯ�9ϒO�WN����0�6�p{gD2�g�泦7�B�7����s��`�Q}�B��U�����8>�f�@XV�j�H+AJ��K�@�Ao�w1G���>�9$Ei�:�շ:��¨H+�N�*��,u���%e[�s����_��'�_wOIJ����Q؀���kw��C��Jq���8����e��}�����Q��P^���=�$#"��n���Ws�eŽ�R�qS�����<�fϚLsڴ�|4��+P'alҙ��4cO'Cs\T�/�&�vxu>��XM�o%ˌE=Q�2:������5�^Jg4ýul���#��y*^y �j4̋t��YG1��!Xp�A<�)*l�����%�5�@-Y�����)� Ie�S%z�[��[]�����v� #�bR��3�Fb�w�n�Σ��#0g��q�Hh�&!eT ��%��FD�+5Ճ����;������η�x !нb��� �5P�^����	�Ho���0��!&
�N��>r׿��w��ܴ��YK�f6��'U0����8����3`�8�1Y�ۿ(/ԭ+�P���  ����R�
O�#�[�X��K1k��b��M�R&�ov�z0��[�a��QFmbv�)) ё���tev_O�r./.X�nC�k?�~�.�]U�2��@�`%�0���Q��Y$ϚH�
���w�
r�0��;@=�"�E����J�j:Z#l�4+��!�.x�3�_q�����c�tpgM�h?���T�8oS���$�N�2!����1s�������in�����T>���J�o� *[����ڨ��{��j�!k��x7�������a��]:"�ͻH��/&�U���Z,<�Pb�M[׀�d�C/Ε�up_�zH��X����d�l(�{.�uY�.��2T6��)<��WE�7M��E��]��>���W6e�y�:H�0.�|9�^A/��	�;��X�Mr�,�8-�J��p��Ųk6�����	#:e ��T�x
��9�~�m�~|�q���>L�A ݙb_S:����c?�"`�剓�	럿%��h]U�n�a�S��F��/n��:�10:6)���������۶��9o3�9 ��B�:��ct��ǖ'�+�_W�3_��fV�/0L�Y|��p��u*ڻg��ԃGF>'O��o�p��L��^�n�p��%�n`鳜^��-��r���gkt�@���^�7�)�9�-��Uڞ�/F��A0�!c�`Ef�=}+�t��J7��Yjo���W{h+��D:��8ӧ=��$�f�( o�q��d��|�?���K�%S��2���,V��5���l��]�d��|�{�%�H�����La�YЊ�f��L��zw��y�;������U���J^f��>��ƿs4��(^�fɄ���K"1��K�wSF�ꀟ�(�u�9�s�ml�c�$��C� t���/�2+zpK��S���εG��2l��h��*N
Hs��Ԩb�\P�ޤH���`��d�3e�1�}��֫ZI���ˍf؟���!��D���?�N���j�����@^Sp�~t%�X(��7������[�yU�2�7�����������a��4~#���|��ٿ���;�`-�I�:�d��r�M�Q$,A���:�2ڸ���om�âyĠ]k�uS[�ɴظ�4~���x�vs��-uD�V��K��`�^�y�xIL���u��%hX�I�E��z�P�b���K�ů���e��y�p���;Ʈ��8�]������,��~��Btk�'�����T���{������ 0`����{n���ڏL|�����w>���4+�ͶW��j>��o
_�v�:������L~��&2PM�����n�4 Q�� eB�1�!?�Ex��b^y��Q��,ʵ�#�{&�U-�=sB���4l^�R��Fiݬ��� ҋd;ks@O�組N�9�ɕ0vC��	֕��I^�SS8�;�Jt[di�Xm��0�rF�cmE~�2G9R����i�c�>+u�lމ��j�kS>h�ZVǑ=�&��rWf����;zX+V*���:��Ԍ5��qa����d�: J�i�F��D��
ͥ�� �`����%�j�;�y�'c$��5���j�L��S΅�!R��{z)�+r����
]�sϸ��g;�N.o��@������dȓ����QrG�ѯ.��d���!>���4[���ӏ���
p��PX���1��\�;��e�1X'�%��U��w����^Cԃ@���&��Ԭ��`�pPVR��`,!a���|QłZ����X��$�n|q�Qi �M�b�j�#��E�@���p@�FX�Z�X��M.=l����Z���!�Z!Lr�F�!�o;\$��3�O[t3�H;E�K�⡸�Z�C�