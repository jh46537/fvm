��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�`��L�o��<�T��u_T2�MA�l�PӁ=QA����9��_����C$dvp�q��˭��|c�y-������5�1/��5��Z^�� X ����d_Y!��K� �B�SAk����S�ܖ��N
�֝�wHcl��q�JU��������p���J_�L:�'�v���'&��>��f�Xݴ"�Q�1�int�G��ULZ��8�5U�ϡ�2|w��
�Z�>��o�м)��P�f�N}�0��b4�9���-b*�N#k^�+{�w�4oܚ�#��@u�->��r'�@	Xb�7��Q~���U���9˂�>f�z��{�#��o�L��r�֖�=�i���3P�k�ƽ�8��@tj�'�2Ʒ|S�V,PO���57��d��Gyb��bd��!�چZ$�i,*�߂B�hZ,6
,�ɏ��kI����P��D��;c@��|Q� �.�ռ��-�)�>��?���륹ҭkm	kt�@���u����������9���[��B�O�|���D#K��[�"��z�ӭ��d2��]1p�����H�>�_��
Sޮy����F%��DUu|�ί���[�p��3�y@)w�"F�� �$����mciв�9�Q� <��\/��=��1o�hh��/&����gN@.Q�E�����b�żu�a��.Ũ1`�$�{����4K��[�~���q�1|v,Y��Yy��ۿ*���vƫsc@!� u_d/~d��|�1R鷯���w)�v��
�4)Ҽ�L�#�ы}���
΅*OI%�13W�F������ɗ���~����i|`�Ǻ�P���[�6��Pw���|u�BU~�c�;�<��"q7W:2T��Z̈́6�v0lS�v���'�$���1���^.���p���Y�ْ\0V@~M'��G�.��+���䃰m��e��:��X� 姁?��X�������S��1Z�ɶ@X�kǴ*$�@����gYb?%VN�Qhe[G8��ypʩUu ��КZdqq��O���S�aH�n4�� W����m_�DyIm�z�: 'D����e�ɼ��]Z���,� �]�����e�u�6907�%��yٓƮ����yX%�� ��Oܢ��mL��).R'�\c�H)L�j94�[��V��Q
Q� ���7��%�<1����W��O�Wn���dY�O(�9�j��b��np����~�ݻ^fP�&C]jl�Y����;��f����� m�#sȭ[��,h��\X���Q���(�B�B�4���{�^�������T3-���\Y㉀��r]}���j
�\h�@3}�c/y�H �������Vkh�ᾨJN �E(�6�BX����e�eNh�xyn����s���KWI�=m�����\P5OD�C��o	��g	����K�H���i�N�~�}L�<z:Ϋ1IT�c1W9��
���_�P���X٭	Y-=n�q8�΁�bYT��_������z�D�~�9f��+w�xM�L�mu����XG�_�)�X�VR�@�������ŉ]=�{#���sw�Vs4�L��n姁	tc�DhU��]� |�׵36�,C�'�] P��R�%���bc�{r�v"��������-��K�X��}��0O0�?KP��'���AS8�~���s���y
��"��;���V1���g۴�~mz�M�#|gic�J���?�+1,�CL����p%��� ā�xz��s�A�O�t>)KJh�|V:�}*�����ϖ���X����-}��K��+��
dm������`9=A��Efؤ�n���,	D��(�!�m���ۄ�/,m���O�\7Hy�|Z�����%#.sU�qm�7��V��u��C
�/%�~ɉ[��`W���{�r���8��jF�S~����S&8�Bq6sb�Gt_ֺ����%���uqn;h��kg��Y��p��2�Ѵ��R�)�/�`��Oh�mm}J�����%V���g|�q�geu�(��K��c�8����@�;v�9�����1�}�t=&����nD��랟��W����t3��ȹ~�۟\��P@^IL������];����;�K��Ѕ�\�e.ׇQ�:�ϭ����5��BȆѾ�A�z'� �Ӣd��!���5��P�N�k�ۆ��d�o�F����\�G��cˌ ���9��=E�b���7������;}W�C�l���b�S���dN3�sPw��ͤ��d�<NΞ����=������J�> AM���F�Ip�{�틈w$U�뗖y�^T�I4&��2�(i�|�.'���3x4DT��Y��T����vv�ъ�:Tkg�ۻ�t'�����;������9e��(��	2�Q�9gf����J������|]j��,b���!�]�)��!�N�n��lp[���Ci��e"^OʥQ�c�Ԇ���,�����B=�峿۪Z�'��4.����E@B{�[���˿�kƸϰA�E���� :�9����*2�����'�� ,��,��Z�h�w:V�$w��~�BўD[9G������.���R�>A��ES��טܟ�9B��;��R��__ߝ�4���'p-|V�f6,dd�&Ό=��c�6o��o5���UX�~��[����!t؅�ɺ�b7\�\x׳zH�ͫ5�Z�tf9���)��Ι%�rQf^:X*x�T�J �hYv��Gou."��F�om�l_���8���oBz�