// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
W9h3GeaGx0aF4xP0c2DIrgpe5/ej2R24m4AHXRcqvuILzYl1GcV660wi4dQxnflZ
OtWUh2x5riZ0QJLHce4sJElArX3MP9y88O8Z8qhD1Jj1pq5oBPg34IUl3YSJJ8CO
dzJUAgrhXr6pFZKdppb1CGYELdi73OVNbGiQRiyRDfc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
pHYgdLW8B8XKH5dLgkpInw4QwfH4N9S463Io5piStCnGlW8foaAGtbz7thlXW2iU
NCPxIpc9SuM5ZunU7rT5ecarYEnhsZ4DAuJdA9Bi7tnlSRclHPY/JJ32TZSKHyBd
oPIps57GAyelrQ6MHyDSUu1B2vbNYV39x2T5yeIpzICGsNP3TqgX/uTjw1hz6ohy
OIG/qLbvhWRXaCBCuoic1uTy9OKKvsqorcLK6i7SfHnbetSwSwE9R0VuSsAGPj6e
f9gVPj7YcakAZrRBDM769JmndjbUxTUHinYoq/ZjTR9oDBHJUIsnK0qSnxPsHu74
40zcajfYbTI0IxXAav7yRxz6bC1/vJI3XWSZx7osjb6GFDA4GJOtHxmilAGFbnu4
EIsn7OSalRvY+gspm3iR2dWw7Z7Rs3n5ZeIcP9MdrBE9dG+wEckysIsyTaToCYzc
BoWHoKv3W/bX5GMKUHXn4QitNvCU/JQ//dF/w9x40zrd3FhLX1O9lni6xggMd67/
CCT/FA6qBtFdsXE3a1M4OCzFOCqx13ReM5de7GrVhtlGxvuiVKrp7/VVMGg5vNai
O1eKWm+VG0Q/z2KeT1XGyMO/KlJ5Y2mgRG3ILxSq3ROXxfF8subn8ED+A6sNbTRg
TYfPWRci8iqKVSWz3P+A426jImDScXBaHGORQSKFQa9owWypPCzEIHIcYEwJGeit
LhROFBLJvgrNYqwHOavqVvmhEVX3b9drilNsONUc6xzVlUG8+392ieAKSyNALDx6
751XPKmuwYGJFJhxyg+yILfJe+R0L70jFJiKbMQ+PrzQ0H9oxzS5Hb11I7RbKUHu
SNVO24V30yw+0CHvEd/7BXoKzUfr/9sHozDcmfpb8dpCUXWgjb5a11cSUQJSrbB0
SGxG4K6+pBOVMgV5LieaABYEAG0gIg0reMsc7431CmdQInCpCSpO4wnNDOsNjjiO
NnVtqVDa2m4HVcj6VDNy8EWiLbBr+YKAHMoWtIdK+EkPTCkjcyeFXYKJLYy9aY+v
jiEsehT5s9aUOodk2pW17H5parDpxSB06rTbQLqkkw6aGtmIfsavUcx6XQVZL+I1
UDABD8REg64d5wTZ4IHwx+QEBhV0y2ev6DCJHmaB+whbmi/g1YbExBdS+evRmqXc
TDFBIR/hhJxmI6OfuurWjkN4zZJgVbMevOiCTVcFvFZT4ogbCPYzoxmJCQ4j7ICn
gDhYdURCbi3MLF4xDjYMZUbjWDD44Awpv/cy7Q+89NCwBmxr0fCoWkpNDt4B8ZZv
ZC5kb6pDpieNqYIVFmGpRwRwJxbJzR22dOcThJnh5JdtQvnLkqUzrz9C13814F4Y
k8nlr2DmMpZAb1Gi8kb5b0eWcYbGlHktEu5O5TV45p+AUmb/udhdyGJ5Qeuy0Ji/
BZkSrkdyiGaUoV42XtdPSGZqhJsfdBpZBTFxAD7h+1V7W2AU+gnnRZg1R0HNjaB/
ACENfAzIy6pJ5sDbZlLWjy5H0q1A9d/YQjKnqHtwnCJjJKzUnLN5Sxfx4Ssi5ELQ
oAKN+4OVWF8Cg4SqLo4xC33OF/qr7vfnMZkM1JfQxAGAX8s0Sc05TMkByUkSZrUm
E/daI1RqXGJOmv6SAUA9cNBgSXPQNY0vr5wx+20Wd0/Z9WG4UpwaI/89dDEpEpkw
me51IdZg6H6YClHhTbkXta5W7q6cfN/AXcysJWlFpXoHwr4m1HfijDyez2X3CZwA
fjAlh0a0f4PxvPVSAAuoAHLRJLyvKahfJqipeYVSArJ9j6CaOMc5znIMX8mKZHoU
YNUQyH0jXnTlCpny0vsbzUjcyPC0ngtFVBxRwiEpzypa2dnepw5ppOsVBY8R61jZ
cNbtQnfCCLa31WltYOgbqXOle2Ji6uSHkKnVAOUT82DqN3mcAI3C9xgNtRWyjwpC
xWAHG+JSmZP4YqqV1zuc4FK1nIJrB8J3s8M77xyy0nJS6q1NMJNUylju7+H0Cqdp
/X6Y9e5VkRfeSd6l1nei0KTayknDETdIpNYeR6MujKVik7SHKDJCJtfZ/UvdGPE8
fgbXY3Csouf+JKIJjEci/Ci0Cg+Gg4rYzk+MImL9uB1LutcM76z3KnCqrtF5kcQW
ivK3q/zd4/In8nKOb3hauTYK5EZxOYfnh1y0O7nNfYSozgBRB7B3AmlEV+/+f2v4
em4h+tHWZLjEX/GjADcBtyXQWq11dN/11psyAoDCG9Ehp+ZV8EnPe+1l7yUo9SZS
ElL+odNaQWL8kiDv69xHjMZeicN4nnZU3+Eg09Gy17fNsNSd3Cvx/lqopUMgVPlo
ZfHwLt2Scb9TvpZGPDtP3N4DZKJstb6jX6APJASmA1nI2yF8yqjb0H79YylVxVfp
Ie3E/vv7mGC29UGvgELD/TKrCp9Zs10rubAOlawIAP+jsfzY8MpJpQzepFSuirNP
0u76LE9trOaHvrUASJG6lgC2M9/iJI3VRR4PiWH2i6nQhutR+teaqHvnG98yILVD
bJfG6+e5H4WCtRYbLI8+aGKx2AfED+gUmy9d8SZw4FxA+1NKRiZ6eaIXhFZPO385
kLmQ9ais+ART0un/LUB6aVIySg1uXGyqyFmXP+c6zqQy+7Gj7DsLKbZ0JYVh9xfu
z2hOCqiA1pb7kqaHOnz/3cRC3KUZ2dCavwYiAX1kENO6qYryX1aiokKhuovkSMzl
lTpIS5EzR4V5kanUXFvMj/r5yyh3gyV7irCkTvmdqKFS3T7/xUSdBE6ukmXJROsP
KXvIIumEPWSPiwUIfRRc9D+kJ+Gqfb8lfoWocuxBAaBaZ2Q0wDFyvuulJqWnU3T6
NBLFvIXe13JumOUfLPv1nwlaHHmb0iPG6vkCWPIFwiGVtLi1e5kgyC6Pjd9KrN24
CH7SuNAiqE//TIIibTJygF/adMnWcZeA0TLUEir8hOPV20d509U5+cfxGPY6PK7e
OLjcJeDiArVU2G7GvgwboObs/6Eu8Y50ljPW4x0mTqRH/2lY9MSMTtG53ElcgmFg
CWwmgmWO+/8gz871R14ExbJKk0anLG9Xv67qPv1Qq1cptupNfvdS75Q9JDOueKge
mtLLl81KYHXM7/rpON8T+nc7brsJXJvDPutWN9f5++IZwk7/DPuMJURsRkT6lO9w
jzZ5rA2VncsmkIt86gSv8wKgfZdWLB3LA53M0we049Y99CO1qHQozuA4oeYNp7LY
nioRbqk+ccjDwsaNFL91vwFnlrQTidc/7rG+vJjcP3wX7JNTBMQQ43QBrbB4pm9V
iyEA99z+MHiPINbih9ndXIv7cy20JsigSBvhIUtkKnoIZ7vUrP+1drKSWjKW1e9P
lbAjeLRT3ocTeQ/nJKMvm3RFLyRIh1ncgUmpK9NSRX+wNiZjHoWD/UY5N38aMAhI
lLW11KP/dWLZXXEAt2t4wU9o0gYAOlT4WgLwtfKLn6Nylyx4I9Lw8bSZquOmHMvF
ftnurhLl2n4DLnWI0kcPWcvU5GZ9XSL5UMd4PJbh9iJ8CUFaF4n3fmlgKnuYHHp6
Aaof4ec8n10hSrvICJc+iPue0ACk0N2t4BsSlZMyCTalxZF8YqAI51mCiqD+CW3z
wHBogAjrOnUrMSXDcPaHDRs1GoFm1hWT5KstVL6h7tJ12OO72a6D9q1D4Pv8MFOQ
2IrIbwe/LsXKUuVQcoUcQbSqK8OecTjrZItooeF6iO2LbLhiRo3sc45MQ1nfqbow
aQt9eVSZhlLpEktkBdiPfVc2yHkRH134liNVk9znV+bns3IwpqKiZDse7nfOMxHM
KcuIpqFBLQeQSaIME19aBkC+vtcGh6ZtrxlJ6S+56o13akRQV40rlisBhS3/gO8I
BSW5BoPgGI7FsiF6vd+50nDlAvYU682VmfTOxDM6GqjZ3+S4rsWhrwZWD+X4MnVK
h5aotQjlXxmCPE0cE6VwV2DvQeXhItKJnDIcF+/AEF1SUC59JItqFSGmXgMSXZD7
AJ7ngP9T38xgJy8qFECisiMvzpDW30uiOzCe/4PCG3F2qca74IpehPrkLziHNq2W
GkoU5ifTadq8H64CBScjo1jhBl1x7lXBsNbyskbhmwkEKL5uZkZUI1E7d0jaPKDx
mRG3a+AeSSOpru2u7l8UswkkjxPNvx1d7PUPKnUO78UBZjYAtLIxRBLWPxmEYVf4
fu7cPMWTkBpWYSlRy4QZLDuPVk/ElKjk3+QaacNPeTttZ5WmbOZQb7ip/N0fzCNq
Nj7rT7yWhBLWSV8R/BCO9HVh6La/uIIAKtfQ3AbjjvOYFQuTOZkgij1AeZtUr8Q2
WZ0lc29wuBPRO8hFyBRWDCLtprQp2SvEfFrBJWqivvqHfxTv2lCFZarxVyjKy9cZ
+0Xpb6mPUxOKyKunkMfOK0cgPzzvc4zqqFoq8jKLk5rO84uwIeYYJyYPLocnQgux
IzCOaFVGMyU5jj5y7lp8uL0+BBKhuXCRy9MZP22QrINCvKSd+N1Ia66waZILDeDU
S4tQyD/81cxYEbhhdSrySHYiogWpXmlBAV2aEajoXNDh5NM5F3xxXBwb1Pw73oL0
7tLQJngm6pP+PFWNhCylMSwoJcz0vs1VV/z0iybXX/1XkzF+Th8a0/NxCiFzAD45
W+zqdESRi2z2j19pCMZJIT/VDfGeCOzp4HEZDgMQpw6NafY5/NBkHqHVdmvxYiDr
EEdnC/8+ro3/ECFSDLfW2kSjsDUDLaLdiX5F5by6vxoDTZidDYxPyq2ZDN49tVAy
pBg2HBNR2k7Ofmk08eDeXJ2JJoRTFUMqT59+mm2Eup5xeIYHBco5lYtuk9PzF+aQ
G70QprhyVd81D0KDkn/NpRJxL25nC6PUFX1AhUYIfs20KuG3wySC+OH1IYn/Y+kP
hPyKru8/C2SY0JMlVKlBRhuX+DAW2cg+W/HUHm8+RpbVdeL3xRezjhRmYheuC6gw
TARLES+dE0Ruey0ZPUt2QrEddCN/coXVUOYrUpJY+yq0kJG18UoMwme0WacZhp6y
L4oEbXpTm20vj3D3Xi67TBUEiyjRAk4IDXGi5xQaE/NwTCss+aGY/q1kYgQpPffF
6pGAvUDxgY9Ej85lr2avAb6219p125cOcP7BMoA4qpFSB3CiV0yuQBZJySxwBiwm
OMmgdFQQ1q7BBCn4tyF2N0VDW1FsruiokT30jWZkTJPO3AhguPjEnl0SgfWBtFY1
ZWwJnpPG0NC78lq1/7DVTldeFoaJ0DX/TmViy5LOHX5EV7PnUZsied7hzULRXFOS
TAd+kRQyeaxPsT151GYuv6uG6HI9d4PLWVfmSzOcyd9ydY4EFrNe59bLv8s41yuv
EuQfAaOBbgy6z1D+su7S3eNn6NPtYPR3JmseUVHGQhs/uCCYHcsXPugkR3xjw2UQ
eKIoiaQO6MyyrMEmDEW/ZET6+06vFM/iCXKfaDr7Ty3syJwk7E64bF2pWxE8r8SW
BlJv9GwD5Ek6DS+Nf5/m4pRuRNQStatpnC0hJFsZ2jqAHC+/S7FUzn/VtWgkXFkv
4oQCT6FfsEKMOxkdA3nrXezWDXEtzfaAi7OpbdHghNukP98mlcoc8LlhkcX2h+j7
9GWnQi4wRAQK6BvRnzwghEI0JEdHpZjNmsHq/7+fijtEv7hgWcPiTBXzLdHm9hsL
AIQEPn9FPiERyDv7f8CACTSNvTQ1togITIg96RGgxvQk3iYzmUNRNCpgwUiWPCEf
VPGuFF4jHrRM3WvBdkmFTdYl3x/Cj5NFrC2UkKhnFzw9qW3WU5KrQT0VB8aAQSC6
LmVEoTH3aYK9QuLT4okQZ2BvSwKyxse7E93cJBpOW9AznQwbwz+V+97+CHZdB+6Y
ahkwfy+5l12CHaGwKDbsbSVZW5bw22imooyaFrkoLKdhddZVfhIN7zydJD8OjStC
e6jlDHF1LREsx6aqeJsxBhd/qH2CYENVNv01ZIizfTpLv1sKesRiZvLfri8QKVCj
imyVQnJhuFZeZz3hgQIdHLCwJRvh3lIK2IYlGEkkn2us2959u5CZrIWeNu79kZuE
byWiu2YrfYIrBPZqf2Aj2bs020uzZCr6nMRK/OrOR+Po8d6Fp44Jj6gEJ1+u9nZw
y7D4wIRJdsISuz0OO6VK3O28mgzOKkAEeIn+3s9O6s+sxFIig4eeL5Oa9bNbVjoD
+yW4CVGNvqBwkenxZmeQEB/eeAHkZYO1ZxlAzkQ/zHFhd9jDTZ2x0KT3UroSPB/j
+MpFh2lfdCDFEXstvoi60m6cRQ49wonx4H4NGghjJlZ0XYCtvX+O6w+rVjwylXTO
tZnJoum/OrupKv2LUP4uubIWzWTZrCGXngx9Su0RgmNAbd1xHmuRMrQ0B0hrtiVk
ADAQ0UIddMw7NPxD4P3k7wBGG2b1tUqiWAq5JLrTI4u1LYslbXlyGXXDLFmjQ3kF
s8udiHnN8kKZuSVLkMzf+QLk8bXtp4zDwI0+dGIsgYklIfRyeHymoCzA0+A4TyCk
/0zwWrOUcQ2WwoW6IanbHoLLBWj+8adXbiviWW9qsk4R3feH9/qlUs0cv94UTyHA
D76p08P+9UtMeQE3EFCX9f4M3PT35SNo8C/wu9bMpvaLxbkbs8ftPPuJuIQiD0WE
8uZSlkIxHc4g5SIzBcXknVAz2/Gq5brCOqugyQLxDwYkl1YbZWyEK6ugJmFx0Nmx
5O2rHTJYhfZqomk7TzjW/3gJEWp+8N4jIiLiwjm6QGIDe8Ojg4JlAN4oB9ti25NU
L7h6yPAsqJu5GSynH+l4A2d64fNo5zZw04tlkaqobiuRpAwI7Xh34tlyRt7Js4Wk
lGHxlGj13t83XsQvoYoqmi5qHcQ82EB4XdsN2iFCdRVqCMwyIr0UxG8g95ds/up3
nxFtBU8cTlOKjzBwIfqoajfR1cOblAl53nDD/xyEZVgTV4ZLGeWt4reCtJstqtEE
tjg0pYini1rjTjXuEAdneYhJzvktTj4Iqb1ZNv/1VSIZcOmyHVIs4QBsg8fuYyL5
HgXzB86oNYwN9oUi5V0gBj1hN1EfB8knUjBJyqW1LzFs840CITcCMGfKPRiyz8NQ
2niSGKCn2FUit2ki+vz4VuO3SwnxomCtVgp7Bxi4ddP8/NRks3d2ScqCFZxrYH8H
6FBmm/iAAEss0pdk7Mvoph8wKhGoTsapBxpreyviW87ULsuD8HRkBnIdRcJtZaAH
8QjsmIxyNoNklIyzDbfup0KKZhFsAruptKL+o1mOTrvJxXVkpo9MEobgnD4Y7wX4
XQRe/Xl6Y9tMpCffGa8keb6/2C8XCMDttI96/1AVffbj5a+nt3THKJ5+rd1kXBDy
kyNIhe3KegafQbUqRHlwFwC9pkxv05FDWJasXWMQIEjjrX/Tnwayk35+CKRQWZke
4IhF27eI1FqMvisw/czE5A8BLEhhNc9ngfx5ITsO3nNwd0prPeGDIlVqINzdZ3XF
8hVf1i/mbpV0K0+6t+QZkUpUwuJ5kzC17XLLwAwT/obeoTSatAYuEzejM1IX+zoW
30iciwzI6DydiER5oUZ1sDYcnYOTeRD/6DAyopukHU3JkWef5t9K52rXTOJ2Ne51
0OzkEsTAshs/u7JeoG0K//7S6bJXx3Fi1yW+RZ5bMxXYJ6P48YLwTuaI5EQQnyEs
LT1XbB5+K1Pn7ilXGRiURQxGAMtn14+Z/Y+d8ZB7pH7mAu5Mll9iNXR0EsgK9ok6
DdTQoZINP7SI9UNpugdWjuOh92xgko4LRoutaUW8ae5Lpf9EfpGqGC58F3zSBYfj
WedCdSLK5EydtiulWnDlaUCwRRMI/+j4TV3FOAts1fa6Jo8iaAiiTIl0d0DVZCpd
X3MPezop2fzPiLaOwdzUG2yNwz7qtxfbmo95vRRKwacdtbdt6yWw6SA16S6ZtaU1
ID8raA2y5/62ZZ/CmjF7bGE5i0ZVOyjAfQxTZfvDkhHFru8Vj5vyT+Ky6e3W4Rur
x0y2tHEaPstwWFoSVXZip3QM6+L82vjzmjQZLLU8lLbg34F0zDgKeHePCbTYAnVg
RfU9pu42ob9GOEttCVyXurGPt7/j51pYP3Y8TbL/PW/6USy15DptVQbITvYkWdoM
VIQ6+q/VFFgnB7YbUbe8IK78Ctloe4JFZPiEPHQeM3Z2uINf25JEdEu6GnX1yEvN
+zSjsRAdbZk1OrtkeQvc5NpedEdFaQBPNaPNs68tofdWkHFjXU7jk90A3TTh/MDn
zseNbonDXwxOOxSSJREm2lQYgDO0Bfz8QVo5RWVp0T7Naguu9uyY9VUNZSaw2Pa9
cOMK+XD3iIvhGSdqEJANYThiKg1wUayTlc63sc8Z8JD/4+XR4lq6hFVJzAvIWx+H
Fkk6tqlM8HqC9BoelVh9vnPmAB7YwLfsHbzXc7MgqSdRzZaXpnKDb7Iv9kl+KblM
0SndKno3B3UEqa9/HtePk63Q+/Hl8FNIewkI156e9MNup9NZCrOVRQXqXAUKpFFt
`pragma protect end_protected
