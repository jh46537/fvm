// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gvsFbAuPZUUQD7jEBZOGgZuqGKjTOEl5vlDQ/qf4N3WXZkXqxXeLO6FJPOnlmwvs
07LhCKAqU9aEO1OJI6a+e1R7gOPz3R6TZZrLXWcQLgPsrHLG9V3mUsBfCwsbRGOy
PHM6ZHg4OgCbQtmCzOUu6uxrajMtsLvoXood6kDD9hE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22400)
kIxTiSURB4Eev+NDdF9WuSXrBwFG89PJxecmWXTKwaoGhz1J21OzR3Ir64xalR+J
QetdkvXfE3BQGXTJ+niAmLSMgSXKBmsOIBmhg0mpFq0hHliTV4RkIiCEduJS8K3b
eUN2evNigO+SOnkIyeVxXeWeAN/ETKC8P9/4pjOrCu5PFPDDwVVIRO5w64vT2F/h
mIP1Mcy83WicY6AfrJuN6J1s/7qhBDBMwiuSUnGPllfveF4UwZPh1Bmvssuwvrl6
vV2tQhPmMJdKGfo+k+qxsKff7Lo3AelQXb53WYyYSdYEdcKHZIaOvtetwPHoQSgU
nMxSYKJr7DQ1ZsuaA6XA9vbLA+QMTlGuvO94Mp8VXdYMmSTM48rhrwJRK6j66Eb6
ilnvjgtphIpb+i3qAhUmbjkzJSnOVQGiW45+LfrnikGhfSIzFMCvKK6lYFRWEZQ1
kB5MP2QPGVoEl1nzZ3POwoF5wTnp3VLJNLtjvnD/oTPlifV2bXiLez/yPFXsZb1A
a6++T9jHjkIYL6GB/TYv5NFCslkc+q/a6uBX4ROLwclCNUc6RPDfHBsSlI+gqN+r
GE21cjSDh16Uso9T3QjAWl2Kb+tG95M9b6oYuwxykmLw+6OkBVRLBn3Y4Y3TBMec
Kiig4NrS6z3CBLAsuucV9PAlpQGblzJHvz6H9w0E8KbXRboa/z/Ipx8mKTL+QQ0j
mNexCumARpOJrSRN+OyAIZSGUGtcreZPhyBfWHMgOEcHrXSnREUfJVBoPXRZShlj
Bwd7Iw2ZnSPSjWF07o5OuEPnAub3o1sbiHNS1PyAUFIQFvfm7zBFkHM23E1JHEEv
km1klrK2qDkV020aBHBz7pe27K6sf4XJoPca0J5du7/u2jJ1ij80vA2TAQG6pi+h
GyUBmBbzwZqOVzg4TngnT2/o9GGIH+ive+w65TsQ1Sr6XJj/UNiwBaGAHW/mhXUX
gdzqH9ano+N2HwWd0xY5+hQ0gT+v2OEAlgFibZZ1+isBQLS3OuuL7UMCHdJnzWzW
JXTs3wm/LWLnryQqK3ebvnAE91ayd+eHRIJg5svPX/QaEL1uPiklsUnCLaE193ex
weCRqVL1fkIFR48FqVcRhsGNOftXkpw6BwnYh8VLa07xqbkXd8OsY2CCsQ4rusGi
NRs0nDKWltcSt9UMtl/8E45dNrP8h7h/WBmGdeRuT0dLd3LPD6/qA0HKQoigV3h2
+43wDE2CXhelemhEk8kRsWDPCifoBkHq0qL1hOh/WWy++DfcCjylpxsnNE0SGE9t
qzStqn3kmgyo0pKO0rUY00WmeEnbJ/4mFD7U37zULMLiyoEpgkITwSRwhrt2HdN/
OnDQQ+Ia0u/V54vksFrKkZERdVlhmcZMknbuybpAzx2O+hVds/sws5aFxGem+ygm
+T56HS00d+YNr5kynPgZJy7ZIR2zu/R9syUUIEy9FFqsqmi6J9DHp9+RyYN0xLTD
CVDDAgxNampmmceyUFnAwIlkdQBP6+PSdZ2IJvJhQ9a2UTzirBId+nCtp4JvChv6
ZxGm7bHk3VKS82XEedLb+/oIDP0jxRpBISJGMhPiRLi9o+4b9xil8Grrwai8594b
U8GJUeEzLngDP1Oj/ip57HCUfj0bJBTvr4QSL2KrUwzKDxmtlTxTolq6eKUVW+YC
Wm32+hl+LCB0dfT8JkHFsRB0yed1+kGrMdsTVF+kX3So2RIRllQQEHgQOpjEtpbN
coAxIKtMtYLrtlgfg2rv28ePOY+juhzmK9FMoV51iRw4FR1CI2kAF4VzD6/E6z1P
RBiRb3VzF8/VsL1QvtcneH9DErCee31QbXJ+mE/zVEvLOHjwiZLSxuS3LzfnJ76h
Mji6XnUmyzJkCu7OnTvjCHDNxABW6eZHlphg8Q6Wy6R4k0ZmBvm93k4p7xnZulwU
AC/yf1hG9DP8S6K6LGtOEq23drLgtKUurIyU1W/98jEHVxvooose/dvADi0X3cFx
djlfuXJogZptLOjaZlkN5Kemp1cnmV96jh1HBckRvaeCm/AlIuytvvFf0OkiJ5/E
+VTataY//kafMXB6KZu4eefz0WWw7BV4J2cnURU1GvaFkt2zgXdVff8LIZc2LgA6
q5hl8T9tL8vMrdoQ9+nxCcS6o6/eJC8NikcYv5VYDfS52bmixSv+Ryp4vD1foftd
X0tifWvXFV+EgYi6OeARsum4w3nm5TSHe/WprgabcC2tDQmd9olBCTo5MVbjUC1N
NJU2gRnkBEUo15Dr/Fvm6YXGIw9VD6kCb4eUiOHyOfOG8K1Cnj1aNCfsut8LP2HV
3gO8nUYR0rlp6dlTLSs87qUVhDG5+E27IoB9/UWzWOsqLUP/ItKBVy6indVafOdX
8G36tyL58+yLrYURhfNhvAxGzD/QZQSD/iiP+T7pT/iBrU8CpuPLPjbWI1iqSHV7
4xeCETaZfmHmbusAXCFAxwyYaicimreSezcT13I5hYF7rcTcajdOpBMYJu2MEk2I
YNtDSz83kmrmFHaTczblojDcgK9wNY9pYe1qimI7c5blklSrCXen1KfHynwhLljP
uv+t6jVon+DPNZMbCA+TgzrQ1+pHyGg5pp9uXQiTuHDJdT92M+uibNh8vVg0htFv
4Ss+TsrSVXDvPZlNKGL3nT3/+crJs3fUucXOE2DDOS8fruI1HOT7PrvPTatQDdYi
NyifRS2dT3G2GXxTIblYS0iYh5cSjv5gkSseLP/ynasM7CThW2vTUJZjwwNtx4Le
J7IuYTPn1x3tkhEUBO/Ez07/w7Py6gDzywl9sVNECYzCEWf+PbtAPNLnhBCM/wng
W2nMG1AtPqNx9ogHZNnFJHVXEDxgtt1LFbmyipgkl0cFQ+eHmHrap6GZgHk3/9oe
aDOxn5aXUrkx+7QoLS/1ueX4lliu0R7rQeMR78vxr0HUwjJK6DVgWUeufzgaoOb8
4AbXQ864GuyXThfo7YECTRq5wWwh8h7Ce8/zscC2RpM5XMEEsfjWBCDkfCCmhTZq
SoWWUsLsGid+9oSIFQejHW50ZgjHrXfPWOcCGRbJ68QGNf/PEvnKOGNDSTDW4Bob
m2UujgyTnS294KBHiFG5WBsDOWhszXBqTuklP+jlKr0M7PvRz9A4JJDwlr7ulsEv
oFp2SMpaZYpJgjPxDlXnIvIA8TyV+a0EEqp9H822TmX24Mm623vycqYDhb0OTrlF
q/3lDO6bUAz0GzVO6SrQ+zA7T+buk0LMluhm9VUmX/d5pdUyWD6pTYnwbNURnLiB
qs9bszPd9E2k6Udg973RqTkxShUh7cNyTOdquj+RA7faPuJlYDmfpKp28bHggrex
t3xw3zkgNWdYUtMhV1hl+qP9XjCaYhxh062MbbqoeOfHZcW2vfLtg7JmdMMwPCba
zJT82zwN/pEwuItNaK7BBK99orXBZO3bUba/Yx6WHL4pK0EHCX8EUG+OcyU5K/LS
NnY1tOP53Q0GdHEYX8oS1FVdveT2blSwpzKqBAdZotKtmDfMtNwXUK5rTVueW4qa
S8yb34wVNx+qTbnpAU93J2vayVpN7z7f3rJzPxScJ5Fa8HmhcmxNwUr8siJuj6W9
VXqbJ9/pvbmyVotQnTppyAaRXj/1khui4i+Ioc1cdbsXldRsfi8fd9U+5X0+z1xH
c17Emqk+K8h8XPYNxpo/OeXvIjE7EpkBShyWNttF4FHqVLw2YspBVJkRTZPv8jlD
nFVDPgObmuTLCLfmCba5dH7IsOn+4F8xWYhBw0O7NT7dJ2ZP3tfxjgDeu1Cvt+p4
/IBxtEDvOJg3x94631kPdedzB8aO14egNYqzure4a1EOymB3sw62jB62WjHOC3k6
xHJ61Wu1dBM/Z6Vk0jwypwrT0Fe8QFVHGpT3RRyi7a2/zUsMXDLPY7kfTqXcw1S9
U2eExGIrrQ9mRSIKcttEYNDMZT10mags+Ulv6wWvklwwsOjmTopNLw1RUPleuWOg
h6gw+CskCWhzv7t+LL9i9OYXIzS+1JdF9xnCTbn9VMw+j+exMLC46S7hB+X/f0Kb
B7SCmCETrJ6fM/wxtBHiuozXSbgMmEY2MmayMtxCO5gSk9dKM0fezZyn+00y25ba
eCnaMq54RzdFvhIg5QhZzZoEOnjUdQupcFJ1df71gOAkbgJbKXVBYkIkP7sjOPc2
Zc5nYdwYcBUbw8opX6NC/jBbHBOOr1ju+mOTguCjVNksohFq0+4xXd2DI9XV63kG
emWIjR0SO0LaKz3U0psITaG26Mb8pzs0URKoC19Ylc8E6E9p2jUGayN8mnsQ+Onz
neldNznKvSAnDgX4YrGXnR3pbIn33OvuSfee44rUGcjuUqsmVq2lPyPs09G8fvXM
HUdWh+dGALCdCBtwHhLQOXCDhDugZyAoeK6J+KVhHzq6A0oW7J9dMzklDjcVFFsX
KPZjQEdJWUgVW0PJOCb0Z9N6MwnSGLoRpiCamlF4MgNiij4KNw4NDIaua78q98KQ
4rggkComiicbpPnfP0B0RRzdeW9guynjOyGix0IGi98FU567FaTBsFLkdR5hsXhX
12wlZBR2JNS2i5ZnxHSY85TTq1O2upa9FU54IGqIwijiYHDWk5QxovJNKhRDkJdq
/0RB1+C3HI29T4cAwkntt1Xb655uxiOwZrknvWNBt4Xc65bPXM+4WGdFCa+4D3t1
phsczhlcdH2TkYwxCc0CmjtMfN3pkIZhdZio1xbhDQVLnoMUDaMpw8PJSCl1ktsm
xxrtqwY8G6YV7HhLp1ZpgpANAOSWd2DFw9iu5NBKlcSiw+7gys0QLwycOJkIW8Fn
GmWcM9ctGrcdNXGx0PfRltzGjZbcjK4oBN922nIR0daosGSMvJRDunxKxhoDTYIa
upb40norlvFAUnhI2mqXBGad5Q9Bp1/km+qcGXDl1ruHVuZyxHm0Kxjt5Oc3UJzT
pg4KRDpZ2XSc8PSgKisMVRWmrjjJimffOvcv9j8pd3Zpe8w9A9zKEnROPjVT2CKm
YY29h1t1+dRg+TnQDWZIbJeMZ+w+9HfCGDs2goiLzGHc8HYpWQRe+LK26a5KGLtK
mVIJq2Jc+cSzK8Fuk7OO74sVxlqjwu1TUQadbnaxPvJ+7bL7Yf3rwopL888GcTuw
4PhlECz63gz7oRirqZr0FlQIKyvqfQLPhiz5rrFRLcGw+kOwZcv7T7NxNonniIQX
4qf/AX+9BnAPa3RrDvKZCJs69baA3cp3osrlUaR12A/4UOyMY1G2QS2h+p4hUy7J
qJZv6s650jVr2ezmEi7QJpkuT+jpgSzslryFvBDVZz5ZWV3XTP6XwBbvrlpuWTot
9GyTVXJd5ttIh760BYfBf7ymEFItYvrzRJMWZ4bKasbCC58uzYfBlookVAxDrkKp
j7+5dnoSlN4K+Rx7WbLp8rTj9+C5MMx/ke5+IaDIzr4Zou8qMWm0qkJJwOu9aA8S
TWYlNdis6ViulObcZ6nWIUTpI0kWoFt5BoTTOSQY7WPMtoFshC5xktI86yMzC+7b
crt9G/vndL2C1UiqQdzHX5rU3qffHmVXUdU1+LXgep+iHfHeV8W7LHKVR1xJ0reL
j5/UsoPgyJ74DQuQ3ohtC1KmJCzAjlKjUh1CxdbYWpqbKYNXKfCQRMBPYgwfU9l3
OZJerXNQ5V3b6LRTly8xESejWhn5crO0Ega2CMj51flh1aDl4MO02Dg5HoiJRGbL
V+RzKGgxzvxV5ZftUgVgijV7ol/m7tgNeLGrbt2waVjgcjdgRH2O5/ijPTqb2NDb
3qJzQDHscSoUiNwHBRlsmA76PVEKhzSs1iTQ+IKnVdklN7B5Nw5Ycv4VTwRPwlsa
ms70q1ArBzuK2XI40FWuUtW7BUiAHGhb/ig2ebZzACZJ+Xvjirf4t9oH2iCwE9Ki
EnrFtkWu2owhujsYlbkVJSvCxwWZsiZB+y0GwGJ/5HfHFHylypllvhgayefx6nWp
32yxgaErJf10HOscKtbgxqsoT2ta0SOQL2vLsutt6yHyyAxDmyJYgt9krzdy9kN/
1ZP3GPwhL2Opf30IAN0DPw6e9oiArh61Ac5CILr78W6NRL9CxAj/H7XZO5ZNHwTn
+ltQWMsPfVll5v29Z9jFuBXJSuntBNMKsVTn4q2HAoPlhja2zGfa5vBeP3iozACl
nk8OX/1iiCwpicWPhPizXSlzSvBD8Ka4De1omLwyCTcPx3SHttT4Gi5Fw341buo9
9Ny8Q4k+XEGPhGehJqVnYjR85l1uVnxB75pIkYUyAT5q7jN5/HSTpThQlBAq/pAt
nqoM7Nxul4BRYzMSuGnN2vXki2fqfZWAFER7kdY2ZekYdZfUWgrj3iF3Wyb3Oy81
eMsWEJ01M+BDxeDK78gbZemz2pZ0r9NUytMVMvcT6LjeiqfV4CTZVbMU0A6XubCk
BK6J5OwAG3KIVSUmz8uhhDaV/AEWwKTt9gwwApMwHSU8H3TUFAhGzTRgfQ0nMBNS
YBWCvbMFEADFXf7YRMBCZ50SmO3Q68TH6qdUndmfI48iKtbm1wlDgXtHVTde9g9o
JvI/NNv5jV00gOs0M9Y8aNc7iN2jQJMCZ9AW7ChtHzrKRVZwnC/GBGR0AXd158/r
aPCm+Gl40S9gcYCpZHKbFNg74CoSiNAewri8hm0DgYbNsO8kC3JKgaUJ3ZUJP6DJ
pJ9pMJxDH0OXj2czPwguGZFjoojKdkHBxtH64TJlDTPbB3kryZWfjk9XYldvGOaG
lbS1q5VcgjC/KvkgM8Tm1dUIki0k4h5T9vXd4EI2k90eK2ijxXmiyVKAufJ+1K6e
oKkIVvZPRdHYfNeNOLpSjpIjaa/kLem+aJjXr+hTkl1cBdjgHbHS/9Rg+PdkEgUV
mwbGIhM0aycJpsGXiE7Xa5F/hXcT8gH3+/wjOTXSFksaX6NS1jkXxBeuwteeoIpv
hx1u5/124iUypP6FUKD1wLC5DO0O8EJIn0QNDJECcraUJTJ5d9ruEYsOu/XefWUf
3dg9XsrRkpUdQSouE6ZUB0QUzdi1qcfoeUFaRUDJ/qgnNl+qsUYzw2+e4g45mSWn
oC+q8RGUOsDTuzb2CfVQ6BY1p8ciYJo4VreEJ6jVoUbyjCw8WdgGCAIfn/v9TP1w
xAyh4FQXyuX+6VBALVai74ZRdd93BjCAB3V/JZvj+sr1GZcQAJMLKQtQy9HmukkE
cIMn24ABRUZZ31TQdusrKW7QwtQc0w8DA+AgC1wrHdCl5MQAlTFc0P+uVN90Vhp3
ileNzaptQ7F8pU6rSS9y22eC2/DoX5WhSCybD1ocaRNT+ozEbgY3xo/xzvtjP5Ap
kDafnS8o4+MCENkZ6JiqpX4PsdghfXCCS2UJxmaa9fhoIQYFj2OgL62gsL2dxx4k
p1V9nhLNNGRzhokakBPAhcY3pXDXWvZN8qYv2VE3cpBgqGXII9AmeEirI6n83UoH
g7hRYn/kpazqyRdK4fCSiPn2MqoECVjsAUlNmwl09Oe1SSaG8jiilGhg2GYWATcB
h293P6khBkoj1ufEnYVTcRnv0lJCqdM866xoPjo9GZIEe581286utDLfvZfgT8H4
s0SpPh6WtwrI6I5vjyxKzBL5Ae7J7zye1yXhg8kX3871u/e/F6bZT8R147UZHbud
EMYQ7+7huYifVcbbkfq0F4PSR+66tq8NPoVzfQeLNl3iXo7UDdixrqfVv5+QumiP
bVHuBRC63tFD6t/7P+h9TBtTsH6vWSXdfvqZHeIHDxeTmN8mg22ZFqFDPbmZDC5G
OsL+784hLfEmKdziQz6CC0AtmrjV9bfkxNX9P3ondkfbjK7YZObA6gLLQ5b3xLL0
0t9u6PQiHCSkPcdwU3Bc13vsafHRkQwJFU2C7Fg9dYcGZcs6xYc+lkMQkOaCx2Lw
KDbN5DlzhHMpNkWNu4GeU60x77X0DVJNKgP1gaOBoirOofQe6GXCCsXK007rpb9a
9RoYXgKEGK/ZfaegBII970UViYrB9Pa+Is/gAiwDVHxcUuZ3yFuQ84OmySB8qimv
qiURnWT5fGNj7f7Kc93IWN0urZwN7A8+3QAWAoK6fpot3+AhEOqgrVAl3lUGeaMH
UAkPWxt4iSLMLD/D7eIKaGGUDzuKDvtkw0HLcKjRyTrj93gPEOAME0ykzt8RhNrh
N5xAWqOHMv1tSCEqQf41+5Wr9tsdviCmBzyqG0OKV4OM2RYB5R+Wh603nrlE6MGA
OaLoXornvRpB5T3DbEN1jTtZcqQ88uJceFAqInb5WJVMB71U+HssYgoJmz2xBSlO
pnCmsj9cbzZfRN+VPz0tQ0miUH+JN7eLJwHcExv7YePFcLJM2Lc+lEHl+Nf5bFyi
or7+5PtRlbAhsbBmdapFn7UEQftszqrhhq5mMOlkCY87RrLB8yYECIscVROUAm0m
9fQ5PQzLWKH149JyWMWIiwbi1XL5lvbC+iSZZmxfaThfbNXkx/ubVzaK1vGFILiR
A7nWv59glZukSWag5lhngSXCX9W67FXr3tZ4BdbnlORODx4a4Sd+/4+6MS0u7Hhb
ceIXxfz2V/7IChnhrj2WipHw7+0LQwowOxkoiS4zpYpVUCgy6GpVyrIJf1IDnWS4
+sT2NPVe5ax7lRVa8ILk82/OxU6bEzsKEk3Y0rYtXTx0/SG7PSEhMJpgX6fgzL/q
UbOkRVJWzmZPbUKla56yzhLFOv6dZe/OjN5N8N96KCllpcLZv+d3j9hdTptUP3W/
ZecHQbHzuiMWnveeGE0238B8w3o4lR76rwN04pnymaDW+9acltQarMQir+fRn3BE
PrpQ+re/MwQg6app/hB6UKGz4hz8YDiNLZ2hGl0xtXiR71F+YgeI2ji++DJZQfdd
Ieaspif5lgFSEB2tRj01AbEFxD+BhJn+mjrgpDEvcYR1XWbr5Wxha4lcdhmT/SHC
Q9x7/rAF9kDSxEymIszdZaY2tGC3ImqhacPFiIEIFBiozZhtIhAWrbDFscKsSrS9
2I1l3q6SaFv5WBTu2J/blJH/g1QVukE5vbRMX9bm83xeJ5t7HVZR1xmw//DvIQgC
jvx8Q/xE7OPBJt41f6M3y5FVMHTGIXgOLZeWBx4Zw00kvScA1da5L397WS/VECuc
NPn2YM/ZTcnb9p8LY9VvvcE4B/8nDhV8p4wh6S9tXORAGt7egrBMGUKZ6HagVUvu
W5TELaNFxyn7AvMRzCnkuGLyHNyFFbqf9nPFp1UDZekrBsjYlLXWtlzYEGlut8/e
8fZZnidCkTGJAGhuFs7EZG91t4qXL2g8FGm/VRbRBX+yuZQxcoAWtPKCTJdotlLp
d/yHo7C2VLMXdh9xlLatqopPJW55IAiNCEd5v7ItnAjo2xQDdH2gGKrpRQaorDQ6
o2xZxwd2qUrk6zfPtXkU8c7dXL0GHp+Dv/DhlUIoeD9wSuKZ18MCKqdnpLy5abmw
ZC/g0Qk+oGM/xXSFJJ8IR0WrRhmY2mOQ6iHbub8AxNh+pSdD0HctC0930xCh3w+D
e8g9S61LdKoy4FFD27cw2dDMve+7NVqQSYqyljMaP+3lJIMFEMCbMpUnLzIvwgAZ
hMaeWb1VhdkjkITBurBxc5IHiX3pohVY85oPoaYHiDltvthGOTF9AZhpOPdvAdmC
357LYikXjF4d79q+JztFDH8inUKHp95fAtjWXpScmcvQOCwjdmAbAIHEK8kTD21i
6rrzvRGIe3HaWm3By4KSXxXLSlQIDQjIvQBaAuJLJrp/0X1q++mrrKM7d6tEd28z
PKiayPOAd47OPIRE5oPoQwI5tcugERhlJ2cD/dQY0LJ7M6RfbLobVVfXEFgkhN81
8irO9rm50fWohuBchp18PjvxR10RIzRIQQjkKW76TsZWKTx7zjWArNjErbswCY3T
7/sNhWeVtVjmwIraAmBy6p25WeEXVMSIoxYZ8hy/iABfvqzcovX5XxKifnXPNjHG
UltJqJGtIMuklhRiMtlb3YmEIAu0hnHFkiQjUKpapdTgQD0iaNarEAd2vKwkaH/7
pW7I+pLVqscxVgMuty4eDRg2VsOp0PkMsi8mX+jd1fUF/+tMb7y8eD7rd3wI+LPe
imDi0gVVPKhk0Ij696NQkxKcxgForUwyyFX+nJpbFJMPlwvIDqCxZ/xAiBv2xnHY
vKD9oesty7LwE2kDkrBrIBH6uQcWSls4kKz31kLfVgZ5XB1cdU/8a+BqQoOnvUzZ
v2NrMip2ObaYhixD6b2eKFINGc4G16pn5TffP2xXQyb+oyb8AV86RPldL8byGLcG
bHS5Br/8q100zg7sgot1SsMbvXTR20CfueQOYZg+APNi+GCpw9HBCOb6vNQcVStx
qYuLoKcowvvCEgdSXD0AfiS1YVlmdg7huuh5tat9Db7ia73cqc3AQAA/TyJJxr74
PQrpRcnbDFOuFRMZlKi985gwX+DkxiTJflNCuQLm00osXCGPofChnFodWZsHz4vr
q3kHQtMXXvtHyKVmGtPGGcKpvKsj3qnY+SEmrxfxzxiYH/rETBnxudqS4MQoLXeG
sym4fsDFcxVLEKne6tkGmMkwH6M4M48cXZUA7Qz2BwbaEkJNGfhPr45X7DPkcN/X
4CkUJVC4ijcePswIHg/2i7HMsU5j3tR1iDki9gRBB/Lr+3hiXrDSEsVt9LzzpyBZ
sRhbkdVYoigey1YuRgznSbSrFtTKWKyf9yJxbzP0SD1XxSXywnBydiDtJSe9AqEA
nr7XktKZ+mi3V9iQoNMfpSujSHDH7ClpRBhw/F1PJdKamS+ePvcRDcRl+ONOL4CD
UxqyNK0hGmvQC1YTmUyDbYWUAIXSQGv56Yv8TtHWcaMnPgA9M0D0DV8Lhxx/M08g
VvR+0mEBcG5OY+KbB+S+lOhDWXYJd1jPltv1+gVmLCS8QQBuQs4wL5rqFA/UlkO3
PYJZ2Imr/xEr6vtBYLBhv0FKGhHVhMLARy40m3/jdXYvLvIKpWuAli6clXDdLKMH
9kACCQdCtbOW9dPe5xicImu9e8Ai03TEL+ypgIYgI2UfgQG+w1+EFZ64SehqThGq
TWrT/31cDD7ed9RDG5YPS/4nDWjGqLghn7teUjfJap5JG24rle1LkBhQCS0fBC+r
OLlOoQPYgLliMTVBqTt54hcLidO17s2U24XOvZgSWSR0vxhS16/QMC0Mhw20Jkni
cMI14pZggPPKJc5eOhnExUOdTyXIF2O+PsDZQMqXxqB6jZr4BBkfuDVTNwZosfjK
gVAqR8FC3jpWNcOcAXuLpASLCVHZPZLhzFGLdNQ5OW5fTp0CisfJHIOGu/EqoiWJ
/N2IQuVRvgAegoEQuvIMMXzI+hMHTy+uDvoKe3NAsGipYuY/8W7gfZjl7oCsAHRp
+1OUDnyN0o2EFNzCqBptY9I7DgT1OmCilPnOVSg3IZk+W7TzyWa/QjODTlX7FYot
mJKNYD7i2W8x/cHbB1mw0O/uzKiWibHQolDSH+QxIplfVeuzlyi1RHQXDcetF9Si
stm/auNhwWeT0HMD9NwsnaTr0TB/AOpD8sthpm8w2zLtKL2P1GTNGvL0LdxZGA5w
XH82MtMSnBz8d8XLkAKYPstDYvbHgVx2NyFSxLk3wWFOFdq0VK6RctkCPKICG3Cc
du1m7IR9oLUdQBsXSLl1qUCvDAJIEJ+rGlLe/8LpwbrmmOqMgY5JjHinCVFfJMUz
vGCB14/ZZhwr5oP+m/5cMO0myRV3wsC9npvfDyd5zOj2JZHsJFxGK+5hRyG/nBH8
j8xH1uoqqBxBll4/s+a9CDt+JiIJiWTSjfWYPuyEbgZo4iMQ8v1sIpNATKnQNN2F
7dAGJEIWa1RpxyEhdFZR9PZMbDtI1B9TjUdwNwmIH+SYwSE7zdg5ONoZuxlw2u+Q
YPfVA0JzMb5ZVIgcpiZ4bdVqJB2KlqmPLqsS26fwh1WktxZdywb0RRwk1TIcNwYM
SL+fDbTaym8AhiQXLsAOA1axL4cFYW0fQ/DH3KX5sy2scN6mFrumOC1blOXru9ep
QfYYgth5bVLF8vIzUwQ/YiEKYO+euhH6N9Ba4BL7UeQqJK/Yc/Cn9OD/zHO5CGTf
cnlG19HI7NAhyOwx+OnE+vUU0SisDQtzqz8qSMdtSDbJaJOFqmmR333azcCJSPvh
Znjta6g6BzJP71VhkJFobUPOcN3r5GODgoOAH2HIMh4ydT06aVmOwUsoweE1f5yN
8XKsJ+oVKVnpHrxIGVhCWM/2zf/PaANTstXUREOR18wYor5FLCw0tq53ZwuXklx+
3dW21CBg1M+qnzzxIPhLxXB9oJC1Nc/DkQFQt5VDIMMN/NdRAt6cly39e73ydWFl
CoLQWvUID0+JJ9Vi+Nwnq6jhxeGSj31S3ux7HKlgXRdXWClHZYp0XG8RIg0S9vhy
SreS2IgCzmZB3iW1VurV4hcVsqpqyWmcPv32B7vvA8Ym3c65PPGRUN56VXp7T/xq
r5Xx3Fe+Hqd3dIXtnBBbHP1jWb7Ecp366w4l9Ty/PigJLdW5y06TOFajaiEYueGK
fPPitS7sb/vlYHbr30vwajppIByRMEaurUa8jmbqVFXb34qFroOAdMe//pwg2jVB
+QDngNDcEV2T6erOWMiq1yokJUoBe3EvH1Teab8Oc83W0XaZ3ETwBNP1shjR8rAu
0eqgwtmKcKpIKENRgxDt8AtO98Tk20YCMosep3lTGEnZ2z2NgHpoyTSwD5iKrp95
u/ODvqm7yhWfmgZBscCLnScyZ80y9m3TPBvFyK5PlmLT7DBYXNfYZlJhm6YjAb8z
lSU4TCLczan9m7FDg6BVF6uq5MiRRySEw5nHTlrnMP8YNIuWK92at8xSd+hhQfNb
gbIbZjABDS3WMd5E03xX4GOt96gU1dhKARXEgKaYRs9hIb4OnWfIKfyEAnobwYcY
mtoEngEBGEHxwXd0vJ0V3/36/21O+PDlOPMMcJu6lBOCknz+5K1NLsodmHAkyhhU
FxbaRBklgns+4hL4ngUmlCCA1t90LkHYJsTp7wMiQHGKY+sD5dh6erfqpLDu0FkC
ZQlEKoBezALAT2dNM58lJN5bpsE6FXO7KFHDog/5YfqpGk/RPe6ltm6pBYtPk1Y9
k1bExGVO1ijaWj6IPLRhqkNH+yc/FQPZAlMf/VL2H8YfW/QVLMzSWuI9tj/tb4kx
w1d9iHsxZKFnz8gAhzw8kpjLw4aNnOIjQI04L+w7iEZKRlewP14Qw6/g9wy+ltlt
chy8z7+CX0+nBwwYRZPs2A/4OTK8ezniXPZ3u5GAu5Xh1IdcCpPDHMav0+932iYh
LVLRRqPH+JK6B+qLG/e0L8HbzJ1bFnR6WrPtSh/SKZf5fcfI4Lg4ArYQsHqP8mkb
zQcnPUpHZ+YTM3wORx2wf2J9EVoVtZoj1F26sD4h8BSp2SSd+Twzfp4ph9terKPv
kDhX0ADg/I6BTGBnXvecfqDLcrEiQJVvlMmvE0TSKMn4IiZr+BUheqjCjnRYlAGF
0LC4bDuW5yG55NePrJ1efiBIiAXvnIdftveyloRKHIVAMj+T30/qVbuW2F1Q2cll
RhQym5NXrMMdFkC5a8lEaHEb4u+2KWWwReKqc+K9F++ioZes56DudINEtHS6IlDs
xWXv6XyjpCPQCWC36hg75mgrXOurEFpVgpET0m7mNy2l5LBa1WPkwQVng0vZQEmk
Y+iBjsKYtt6uraR5jhZJjwbayTtA0KAc7A7/D7YflUQV80CYyKURWk4Etmf3Y9tC
PhsB1tMM2SFCBtG0oBGHmVc9VUSSbWYBQMFTv1qaugwOIym9kEco98sAS5/MqRfy
zwrCmAocsdETAIQqXljLqIvF0oN4ADgrUiMGoZAmU7dIPJqfQN5CDqtQG7r0+CF0
yn1Jk7/ai2BS3gOpX0hZM9QELV6FayOHQ54uHwKFFI6wNyrh+8zAqLxEgdTePsLh
ZQb65Ii2K5+ZzkLROpciJBQe3Ju0lw7aWLM6QHSmSdQHpK80BFOpOUwImov3gYVW
8Jkird/krUyh11gVIu+w2xAmK31mYVDS8ZgOTlzpaY0TFwidwBwaScjXkBA4pff2
5csur8QvwW6rUxAWK+71nPDzhvZmHOLrmtO43kSvhCDIfTF2RUcSP1kyJxOHbr56
UsuSGHxo6CL5QX2C1VqSFUVMOLQjrcjtodXNLS6k2H2nzn6Z0vM508e/3Z/ASEvg
GkHRuzPn5hBXQ4GurlnSkoUOSjYtip//Lmp5fAvAXlP+pJSI6QEX4ixrBgFSErZH
D1H3RF6j3jCkn+7kuT5XuOynUpobFjotNMs9C/g1/VOY8TyjLN03d+AcFxdOKPbk
DRdOyrSMNAg9Pijeoc7OYbordzLi6tk6cj0TZZ0693FTlk16FYjN6zJVb+g9eqy/
SXvjVNL0gM57OKVPS4PVkCpwNcx88zCfDpngcb16/C2RuKJeQReyEoOskVShL7Ev
8RqoSEPVTIA1oJ/EY3WT8/1sxrsy7suEZopZ+Cb0AIPon+nYx92IIihXYxvAsRDk
X3MIoSt3yABJUjQ1+EBewqW1wv5reiJZgPtqQU+F6bmYM/1omxdQBsjsyMNTYYNx
jFP/SWGoKqcjOTjKAoFznkiQAmK71Te7manf4shYGtPj9J5CrBN+HcTy6MOtuBJ0
ef/wi/tsqHDlGo/qNi468jUc3hC7O3K4tcWqvc9xTDNdQ1+aWY4TngG7bvVn81Xx
JQF/HNEtzDyUyx7Ovk3MXO6x4OfsOeuzn9xgK4FF/CtqpsNyT+DVhLzYNzI7qPH3
Q5TMURt067iccvDNjwuUshJF46dMhJpuMiL3C9EXAdAmn6MwDOJk0VU7jJp1oeda
D1ZVQQjvyJqtQsHbhyFto2XTPTsVnYOAzNMvQeWOTYj72j38L5h2oWacRdVyd56X
kkQ9nLTe5/4QDWzzkKSPgd5QRpDXTBwA7CyZ+5vvBZamnBv2ADsHfhOxG3+mbRI/
THu7r0Cn89I2+ErLr0liWTnEnT6jy1cTVJdhUuypUTpsJJ97f/wdqhKKuPo7A0Do
PrRe7M77ct+OB3uR5rTEmi8cXTdR3XuT6eVQs0pWo7irBq143mpT9352J4VinWvH
KdZVP5IUPeJLHVRensZwRqR5Krl1m/8rY9fJZmv/QdOfTHEyaTgkbxYp6cpQyFgY
nii5wg30hFnJ/W4+MXuadtK/9PIRGeGSMI75FywDz59vWpN7fR1a8SmshbvdwKEY
PHZPTVxTh1MlVPPH5gLVu1UVgli3UjHid+mfZ5uoIT4UXZAXXcWem/v1nddKpxXA
Q/nyTMh2HAlkFPJbQOYfudJ2ogki4/3KM4NSAyohE/AytA+XtOPetO2MXapJ6LhF
e9cU2/0pRlIc1wAF5A7lGBKfYelNH7LcZRqSwbAsbNykjOzSZXpv/U4ERxYlE8K3
kT44vizMpox50nUdtgmDkmWM9KiNV2h993g5Rbzb9Q1+a/QNJEB1w9EqlF2lGr7d
77yAQhn6AioCQ27v+HGTvn3/OzMq6WblxUx0hqfTwJHZXcq3/+DKzoAQjCDLlu1k
MGfDniuHFE+yzzX2T5FsIop9iSWw9B6lCZx5EVtAdqwiB5YxBjsgNATQLZIiD0Om
XlO2k/pOamKrQEusN85bH+ZE4LoBCjvrYCxIGEprYilVCaIsz7SIhPc0xWhggbpm
5ZpzCZjCQahw/03YDmGvaQVLblfcQkDbKBOM3oaRoi+a7i8bU+ZBPcxh3Qd7Ojpa
0EV9YPhiL+OayQynNsA1rn06dh04fmRvv0VQHGwoh9q45talTp4KJv0SIhJ+uFaI
rQRdXGQfPUipmXsxeqa3u0oE2l6dVvMYU+nyJ+6rBEO24a7azqKmkpGqcaQALHbS
8G7QdEHjHWRYUI5Y/ruUeFTFxjNJYQm1nC8k/J9LhhHm5CQ4jKgAHJPa76yp99gf
6P8S6/hw/r4ByHurITOea08rGWi+3mZsMChpVaUImFBGHs+txIZfr6mYUL+CEGis
37c4ZuGssakdqLyE9tOg+gO41O9nZvZ53MJnobHJxgo8/0I+w5AaqLEJyGKZwDQz
3W0Y+ggYdcOkfnFpFSK5wlxOq1fOL1vIvtx2ZHgEqWxD4KmiKHKEJKB92gaXH5dD
DbiC4oN++YCP3SbYe9Sm7LF3GJfHpG7hpKEp9f5t9SIEI0brG0eKcHLbfTuew64o
fmJliEFjUCot0XmELCXLY4dx0oLcH9knoKCg0aWB6YMI5ZhvGmwSntdCbMYO/oI2
oOGwFEQY2N01a7CntYgBEL19RH8Wf4FBLtlRAdh8t5Lf5yZt8hbz80ioox+Wcudi
4mO1pOgjK51E5qkp5qjzEMEsshBfsrSKEabKBaiPJ/rvb0+uxEgHa+i5Gj6OgTTc
IM606oCZ9lvecPR9dnJ6iEBkL4OrGOFpIy1Wy/bv+zZ7xYEzc0EH4v9IyP58git0
nt4b8Eqw7ehQ9fM53ZXUtdoTTiVsk52P+0+d5bkxzZXgmxhzmLs9U5icGV6JTzVI
1A1taFr0ZrL4Ie6WXfbPq4wUqzVgPu0lApvmkBVAtgEDTtWFU5a/jCCT0jXd9xii
xw1Ab5eqBTDewGfWDNIMzqatQYGDj24toQhmWrbVFBaSgbM9XdfC14YbbiJQTzkX
J16FrH3jPJ4hFf9oGzun8XFTOcDRaT8EiqYulr7r+P6nMIiwBlhwJXHY0KD2HRmI
LucpfEekZT+edcw2aZacvljosTmrl74uKY2ab9NC3FWR151YQ5HEtDbMYypVSFYJ
y5Km9fML7ZSP6hJg1nDk7DcKm/4sOJPzarJYfQziLUCWyZeAEI308PtuVA5l24hC
9MhQQIWb0dUEmCKLYiWpsqRU3pko0mnzw1ycvdEiAw4SBiefKJsrgSeLs5Z2HZK8
aWF1jJzlcNJ2ewMTvVeaIDsO34/2no2DC0HCncycXjoWf+GETQHjQxubzNui/wkr
mBMchwLDIzfYXCHDyY0o2IyOvayB/NmSqbgha1HlG0vMEvRJCaSQsTh22CZ8UB5G
XvwtunUYtZcm/U9ay81gFKdH9mlxsZ2AWPmfDYOKMf3PWRdWNeFOPnZQaMYfljth
l9uInxasXF0lh8BYwQBqLhyt2QivK9FKxxg2ATLYojkRVk6ttDFLo7QUgbctCfpw
HfG8uN55+un/lq4L6lsngg9RMaZ/sVp9GjQPKs7IyrNBInEBWOCiQNi7LMERLQOn
5/KejIe1U/sggOnwmRB3rMLUOmVr359X0PwxmDPgyBdPi0c5QY+npwMD+yROA7lV
FWrb8e6vRuOf8+vcwplJUKS6Y3CDPlVkWkKY9T3CdifKChVfgTsHjcKK6VNpDcEG
lHWCZdpRNBbxx5uqVfUGEI1xkk9JezdO+QAA48gSnecpWHWzKmg1kzwyt2YNjAFW
FU8PDJpBao8nEFKvZFoRzC5Txy1xGu3EyqBAcjA3D2i/Xn8MG9SZgED+rhiQEwSb
GgHe0H+tzL8qfUWSHJgzjSqdHMZ/t9eukDnJJ8ptB1yU76R2hoqqzUgBU3CK4rOG
Ypt7ta5LGJc7J74mcNRsVFJiWlHBBScPIW1M06tJt7WkaOG3RVx7RKUzPBQLp795
l/32oCMqH/WqTDpm7P3aLzq2IkzUgQsxYjSXfRLRmEfAQjG4dO4LtvH3vNvZc/bB
2EnA1bDEHuC0dRYdkF2PUN9bnPamZOI5dfEF9ASZYYBKTJIPy6qqDx7g5sUtT/sJ
so0FWw/wWQlU5eKJ0AAQA5adLeSuwGD+caX5gQ8HUr4ADVJww0ezj8KazUM4TFpN
0MBv4CMGbhA1ZgoBqhXe3JU/8DPU/+UojcaI0lUmsZp6pe+8LvIMvN9CJLNXIRht
sHyUI8FHe7keDMV5nREfB9dWa2kfc9ZD6zfBVd0Jx4YGmuwFYqKAB43/osyoiGte
8HxhpNnlHsFGsrqrejtousI8RP3hn8rlQ8et2qukSuIKRi5yYEAzGaU3xOdRoIhN
+N+Ktb5N4Ah756hV2LWxC8JLtqa8qSUOb+2nVWPfqfZ9AzJUTKx9Lt1AeXCUQ+iz
TWKAMM7FCI8zXC1mKSbFusrctxf6O7FIReTW05UTvCGCtLUHjkROnyaAQ7sAZlWZ
f5lg6FKRdmL8h7j4nD/3b8QmF6f50fx0o/mFrufL6IKlmm092qDQ+p50182UPXuH
w6DovQWbOH8TK1R79q2YAqpVVIsYS7eTVEw0KjZGVH6VfZbQTbCq5eJuQjJ+dHpI
AeyHmYitqVPqFxzuGW4lMKjIJkKBgUKFV5FmnmNNWw65QoQORRm4VB2YE3CjafIC
9Sgby2GInHZXmm6F0JBApSXGhEQ+roNNM0qEMZAZ5WbBMwNnuOMkuPvtjLGOTP16
nfXmdvPTGzIhVs/aAyGgJcSCOOEOQih5QboYBNQdBXHWrIJ23zdDIrVbMUzZqNCN
k79vL7SivbXwv8VqLR1AJRU2GMVIL3d6GYO+tK7Huil6CSj6BXLf2UBE1YvEREjl
VWE7hte0XXUX7TJ/o781SPhdHNPlX5U35yv1sb1eLDhIz0/LdckqoUotVjzj9MdD
VatpdgIALbuEENJscaqnKKc9ahNMSoMmzjhd8rWZ9li1sslFBcxNhDFHz3Ow4kju
/GYeHcssTlJiJXV5mzI3clC1NSbsatalnnK7nD8CtZEV3YHpKQHcom0rXm+5V7U3
9dQo7GETZV45AyBHaKcvi9puHDjOT1ihkyZlageMrqzYoT9EMpmfiQE2r9TtMh9S
xZraCBsz2HAstbNDlnq62+BF8EOq3g3gaLoD5tieGOk28mkv+GjHTKx6mq/kDoTR
XSGAQMbww/LMmdMLBW1X0msHNXbkU5x8yntcXtx1A4NyS2JWXB579qqoetCx0Dr6
fuHo5PI0lXc5O62RQN/XvUtzRfFD3iDUHzmr7f5mj4hoJ0ewaRudiXep9Mn65kwM
HIyPZG8HW7Y6q2MsGEI84izKdD7CdPMqVuCCljB1gfdh0qLJRNxg4a6z8WY6sohW
CuYsa1sgkryeEnvTagafGqAH6SbwJjfigQdu6dKyDz+j9hMaRq0nAIizMQix4PLs
tDUmrNaqFl5ULclyaDRSYcZHTptf903Qfjg9GLq+ePt8EyDL57MuSfNOAgzNKQ42
hp57i+y8szLY9dhtwLMiomhrjHny+kExGYUwWCaAzubsJTqzCHRbw97v3KTx1ZoR
6x3d20vF7o62ZBssGZcy6M4A8m8tw8clJbOLdjyAx9fjrC1i3PUDqCDSvoyL7dyO
ZNR8Zm919l2CneWmqD+Bms8OsscxgI2l1IwAY688nK/bD4B2oxTBYSTLooMhT1Al
+KyJKSduOJr2pEx34ENxMEgKCwdSg1MFv8gsgO2L1TnMSm/jfJE0nS1zoUXOWc2q
F5hlSPwicSkdpN8HwvxxVLoeerv9gwH6idSP/Cg/z7OtLcv/NrGMynHCkcu5ksxn
8UHf2yCyDA3ntxfQy23HP4xZNap3VIBYuZVAh+C4qPP+8KrIJXzPxKB6LhM32xVd
I+fsNKTZYXFA2vbLcuzLD5yMwV5dG9vKXHszxo2I62mi8RDRx4HRYr5LDr+y0zyi
r5FD/i+AlgnSo09z7UNOZSHTeZ1d5FoKAqmrlf5gW/JiaenegeRphtGbj2PuGiYk
lYU+OjF44c/gMvWDT+w9rw7qCIjJCsYqCdbWNeczDLc+PFLP6Inw9Fj4LgYksbGg
qh4K60bHvt3OdAhwFHmrwM0dCCruLRq8QmNlJIJ4cmjRKegpRCfsUBfqw+HsyDV2
6mvjkdApV26iKITZ3OvPofxg8qcxy+OI7t0LO1b/aR4o2v3TgVOG3YLgzeXE+yoE
TQ2rLM0gKay0cAiEK+kuxJfO7C/QF1AZakJmDVT++A+2N7ScdM/p35UQcGmTqdOU
yIkYu9skDN/hrP+VJ28017JDiFSJ1bu6O/CRYDJvOw7l2kzzhWWFQgD5dSbOvDY4
R6ighQZ0s20FqjK+YTkfl+hXgrYiduQxupitxFOhmVCxtO0JODcuVSkAFLoEHMqq
un7dk3BnnHn/f25GVko19BPZkp6E37yO7MxYVg9GMuUjwKWA8zuW+WTwm1RudFYk
RgbudE3bUjZPgpzzfTbwEhn7/f+w8mXvgPNksfNfPa29I1XOcrywIrROf+VDFprQ
NLcs/v2V4/weRS2DcAms6VuqlHvggJyDH07Wa14f6ruBZWF1dfbLiMDjQlrY685C
YERfSEWswD6rBFijFLS3eOyQx81MisV6oeMAPuwmmiVbNubSgUvYH3k812OAwAKU
IE5KcwsTdXgEtDVB0WzksePvCkQkFvNAmBSHSwpaXcnXFH9t+6qicbxb8SlsRNTF
Y6Mh2DXPCN5+bzbNj8nzdNOVRndR0zzmlJRFE8D2AD2Px7UkMNgmbdPfxCOn2w4V
YaXYRiOymlcjNaG/l7dDEpjYZKemLZu5GBlcY/NAPo+YjC9xZElmkeMCnGTGP+v1
IP/CgzPEqjNLoY7oP3UsayjIEeAPODfUUXorLrvD/T3QGYt3BehKLWkn1+l0WxHA
T3TPPsGQQPd4gLawFysJk4S1n+VVD1xo7smiWVhR0KHVTY4z3+bQ5DyBgLWZmv8z
dFW6bM4QYqtWFmTjEBtm+yR5HvyeiwWAiAR1swpSsuuul/1yRNDFpCHog/2owFJw
AL5RDC2nVZoHhhiYQM9fM3/5JVKUt3wxMB/B9QwVpqioL6D+PtJyWb/iMyeHONhS
HYYjILW7/QXapMnDkIoxehcPUn4jqN1r3mLzI01HNfmVhMUfGJU6UmrSklFc5Txp
4d6mJc58zJ+55eGkpcvC5NFg2LHOYeEmfeeo6FjFGewr/n/L1+XZBQjngBhi6SXM
G2PSppshzMQ4KY6zwVR0fkdqrIbV+LsRzmWLoU0ZtoCd6HP1bEm6IFId+q1ETIJH
ABy6Lsez4Z5/HUzm72Q4MjO2dH5mLgjYqDgoiZLKfU5V0gXaLCZAlN0yZYKlY88W
fx70pjcY7b3CyewyVkUEDuacR78vy7k+aF6wZ2Pc1F3flgdqIzrQV27GCxCsf5GX
7vPu9Ejj2/IAsHmsbNaBwSNMY+Dod9USX3GYcUSa33oFZvjBto5qHKeMm0xk620a
GrfLbCFdMAciYnZCxtWSYRe4ngK3N0rpKriyLKROsBbvgRRYkT4KuhZ71hWHBVU8
32N7CMU5ZqTnRa1xcEn6Ym0jVBhjpcpMVW6mYZuSbNwLxRWdpl+1JUOOYe3g0VN1
b4fSF24PsOz1fKQANKJ9NpodgH3VhNvUYiB3Mxk8GWhUppiqavSxEunxwXv7KOVd
bYJdV2ZPfYMRInVuwXR+vS4zHl/N7YNfaOnehcz2VuHYcUlWRMrfk4HEuXZI7HNi
Kd1a3WwcOB33Qwg9eiIY0H72Q9oMk/gxFyFOTSwU4to+jZBOGaFGypb5GfVI35eF
vbrCScBgTmNb5/Xwj19sgVFVdxkMsb2rm0AkLzmk9v3GgVIm7rAo/txjPmUuU7J+
Xcif986FdQJ/aM3qgMCefWS0tkfUlPE0zxOW/xTHUCMjSfh1Bj3+aShXGJIgSVcU
+t9e2+cddd52iX7lApzsCtOQaoKAGFoDZdIJQSLmUTvLNY4bOJ3p1pqKmHtuK+z6
OSGVm74+6LmM+ASiMvtPxoChTEzH85FjY8FGdKjixCEztus/9ETGKfim6SZEnI2C
UFsb2RPxufAmhvMB3lETK0fD60c6wGrHRn55qHAlRIECYrygpIvmO/oOzqzYqu5G
ojRIZZ00hy0px6cAYbR5KA5UuSMT9dhTAkguHNjziD2Se6CJEo8cBYtKG++hr5fU
hMJ+Pmy4xcUKL0HsJbtTvr7x1ia7jHsl4XwgeidBIo4kOFdkMODhgWyz97h7FamO
r+pZK0glUUBbf9tS0WXDIkXcfJ8goZPaw5mm31a5UCdBGtVqSvO5qtNo7XmZcDHf
2a2pSvYSLtxYyNyzP6BE8xSuS00UhDx3UMhYWmemba6b334lVuAQNsh2IlY0tndQ
JXO3Y9vwGK8r1O07HfOqYGkydAyYE+Ehe5NEL/+WUQ2CsREoYRRcoAJ14FISawZA
14tog8Vakk+L3kpA1JCoyTQ/Z4FsuHY0rLIY+nCUKvdsIthyTDsOIwSeWQrpKCPw
Fo7CQyglXcBC42dkl7Y5kRxz8S+5z8OmRYOGBHdRKWwyQuwr61bIfnu+WDp5XzHK
WzGxx3eM9oqg4Uo3LCMySwyb31wKO3rfeKgEHSkm1kZBxDFDiwGtyp8Vj1AKd+s3
t2ZOsLPh+QIiKEWL6/pE+kS7aF3zFhZcH4qNfoOCxGhhwe6+XCBsu1imd0Jq98de
gpgPprs3vMuPWF3aig7jGBLSv8J5wQASF3bSZ8X9gtwpXTWid9+Iz6Bu43aREmxE
6Vkv79JK4YULcx0P8avEM5zay0/BBRybTps9mJ3/ROmshb4eOyyh0KiKIglotghW
4zyQKhHx8RxdqEcRk5cNo3CKV/zEPjmwSHwaLnrlXZiysWukkPr9jl/qVs2oxttJ
xMQXnWb/XwrsACp/7IRCibb2aGZ8VI1qvkiwy6xmwdkQWGx2QcOohExGanMOltz+
Rl+/lPTrYaT+D9B+W6G3JXyxDkbOfnEXQNtMm1DvmGmM+JEE084dEa7LWDyaIq/1
GnfAghKTkFNaJokTiZwQy35SqSYCAPJ+ALtoKAqN/n4ORaK/MZyySXbAXh9mQfwL
sxSNcxs1UykYrClbZucp6hw2CEEPeTCKet3ON65BDReTFWSTuxQ0R9k7U71Ocz6f
rN3ETjKF6uO/OXzNMpHUtuCdZvQh7soQS2jGqxmN8rqgICIEidUhsmu8mmuXBNAJ
ab8Yfe+IeL8SqjbX1BN0PvaRF8YfeVXFi9uwH54bRr/5vEqcMiwRiaJxKi9dkoQg
Fhr1fRhfLiLlZw+rMtlgOwcL8pDkOl2CcUw6WYkCqrL9NXNJGTbnrYijMvzPUEBR
cBAQMR2q4orfVYVDK6j6bBZgT1bTJB4ZK/e/jzxguXp6glNL/V3T7v+8gWN6IuoF
Gk/Y3NzOJz0OgbqjRMLo96X96xS24Pe4TWibYVDvnCwwlucOJXlB7Yxbu+pFzo+n
uIKhVJizJegPz6Abu1rwN7i+pOUS2c8bkuYez6czwQ8KorTWKUZDVPfvOAZgLX8t
r5CB5f6HGiC3UEJSBNJbf1yzrKQwK6HgoFUmwT67ZTyCejNYGJz5koQbb1LK73tJ
ZzVfxYigIFPXYfFdn6J3p2Wkfsl55ecMeUipOynQbEsLHE0v6X1IMh4gGnsdP1Zn
/NRaqL22WQftGdXEzeXG21AFUe9ADXJwlhKTCl4YtteHB0ahxaf2rUu8viucaZi0
wshvsOywPnA+ztbVsJaziyfrkRCJxrPkqLcUc+C6RSJPs8na0MkOpxTP3/dYofE/
0JQZs0PBw/MC1NDqt3GM/0DxEtqjmVrPXCEOkvq+uCeMgF3CvnwxvQ9T00pSr4yu
nvi2t6BxG/Sud/BgKQLbO7mlbpA9XJDItTC+Y7upkttOyM/PUB8jXnyfdUFtRBTB
Mw+vUhFkiUs+mAMDH9bb6ZVTpxjtnijn2MiPdqE6qJXCOySPnzoGtCMKfSc1M4b5
ImDImMtBjEinxyoy4Sm1D3zcp/eTcZvjcYeVNQtarvO7CRVFCiLkUuDXMskfUr1H
SYFNIgpF0qeGwRYER+K+sgYtt7H5EAwbe4kIfbYBgyaKZehyIyFojguDJeF11I9F
PqpMxDgs5kqcjQ/0SzXkdxF/X+J9SHf4o7NVO8unrWffuabp7fduO1jcM3b3SUuo
ScMAeN8inPbFaXSL+ApZxCG8LDp8FXV7HjEFdIfNfE4JH4WiClVDngzauvlszIDv
lwF63D25XnExQ0cYHysYZ0qNi0+E0WaujvGGWulbXI4H0a4bv0EqFM2CTolCZdUM
26YtgvsIRsNsD9Sq37MJG3Ed9sPADUN1scYz93/Cfm8lwXY0S2jAEm2nxMmIhksB
fomKAbm8q3fjX49cauR2D/R9SCTNXbA5vmUJ6Wo5sy2TPNpyZ9yA6mchWO3uwbHF
RtRK0euZO4VOAO5a9OZfYHTk3wUFexuHtnrak7IBx7tm8feec03MkTGMNmSlJobe
h7p1kc2QkOCU4PotQ1gjvT/lhSvoEFdTSKs1rv2t+Yb/OyBNNNwCB8TcPQX/aYp4
4TjBWye8tAvSpXyjauFpR6Eq614Bg6zAetu7u3ogfVc7kHsI8y0Vu4kg5tfQ0vaa
9AZDEm7ay+fY6evuLUauImagZS/8Ae2xq4OYb0FNIn3z0Q6S3K30UQyvd/VVeIey
GkSIbe3uHONt5tsD+wpn9l6JRET0G9B80Hux36npYYqRluviFu2jgyaQmV3LLQj3
ei3YP01bij0jZ7TbCBRQ3WMLG9C6Q3xiVFsxxE3x4evQoYXBcyOeEvDev2NYNCXX
M+Vv2lStOPz10jV5xk//FYD5eo646CwsxqInR6uS50KJ4DO8bxslGd6/FAmx5g4l
vHTll2wmyJI4zFJEiCGB/5j6P938JGa6eOA6qoVZ1E/OSpuyL5z8N2Mn6fOMH8Ns
8UTNstqJVh627ntJbxS9DHyJbseQazM007g6Sxf0IE7/gOxZhgz6BctL13f4eT5S
mJCCcKLOh62KvGsEiqvNjfAv7UGnGZAkp7At0YoL3cZTwrtBkoTWhkv+qCyX1PVa
ddAxTjGUbdOmxzVbiXzgUjPp8p/BLVXqEQYUVKEgr6/HxjL8yHbPKx84LkuuFGoZ
q6HRR8EdqcTfDUWTWUDAdFEUVUnNv3SyuZUmtBgOYAGcVE1x6rwZiN2nHcBxL6/b
f99j6BlzRmrKZpQG4yqCTAe5hbPVpIAL+BZ56B4QUY1nN0Gb3LCsQjA6oJfoDOfh
fTtPGcqZXpAlT+Ge5ua60LPf8h200TMcX6AAfy/le4kUyfraCMlhysICWC4aCnOC
e6UKEfHqxFCfZgZJEVa1J2VJzfuqYxNRpsfuORtex0yfGOV+CbbctlvBnPT/PPeb
R6/80MOKSOxmpjjMIPQl8mvLq0ECXILM4vBtQfUbYBV4R75F5NfEvJwTAkkHxo1y
wed08yCfWGcPQ4bD5vletH0RXEsYz/W4by4zH1Rc2VwjxUvIyMA4vqAhs5CkeWRm
kN8JnjZmiS/zRSzBUpEyWmHk9aIF1AlArBExzI/x4M+UpuHkdiBeIrGagcmtGc8O
bW9iWrYRqr9cDKfqm4qgg2Csej4/QPrqg7x/DKol/osqg1m+SEaDy0FwJNwzjH0O
/eDEBkw9iIv+3v093rDoFf3b2LqIYhwbNlKyIoAPvHZcPgaTY34kXmM5u6gEa0JZ
JU+JWqDz4RQfUNIaUHf3dxmrCON466zCYWnnvRqIqZBQuE0JkaUM802lmgJibn2n
l0KijnJodpoSoQwPh2LVZ/buVToVVDLDWZMcekCQTKxCx4Qw2QT+NfTIzjeMJF6o
bAxhE9VQjGMMTD2qKfgGmokvyafggSrp7lg5DhKPldau8qGbvvUACUolQLsH3aVR
9BwiUzLiybwNS6v8B9EzDDjzW/IQiNCvq6VW6rxsRKTYxkYRJAKmqLyb6OHrGQPV
s3TcOoosxwt68Ttyfa/MeZUFCl1rAxN6RWrEHoVHBiAz8kHgrlHgVn91RKz/Sd/z
iqDmS4zpPMqLnmBFo603M8sJH7FASCk5NbhgUa6bRHGbSbECkvDk2DGyM1Q9Op9L
xxrjTfp1Kwqt6/86X1XSSfsmWjLUIBsYBY9EnRqaK7mq2zmIfkufJN0LJ0A++Ex6
xdnRvtzyAgiM/Pp5RRIVDKz3tK+U6d9he94rujdgJbw/Pe/kb0RAxs+Ha+qXELq0
MhpUXWsw7a/A52w9j89bYJnr72drj1lPrxyqqta3EXgzF80AD5K5DfjBeGJ38Wcq
bZeTF4XnWRBTrkLUQXQ8tlK+D7QiU7SkahxtokVe5mFK0tKdooJVtfJHoNCIHAm8
nIXKrBbjW0GHSokJhSRUGq+8kt5F8uqBpTwc28Kgw84vLxR+/BOiiKdru84SLLZ5
YBsXAHHk//9Z3rKwu8AVhr/RYY+i1yi8ADIXBR7rBWpPrGtrOweEYlxYcqpB8Oy1
I0ikP84jmuIYC4FGz+f+7y6mswkTNWRoMFJRl5P/kFQQknRDDjLyETELpl/5K+TN
9R8ifnk0f1XAi2JcbhhXhU+yilAV5LB61LB0N+K7dylvrJJZVGP69RtxG5fWHliN
EL6UrBdEilBB/LYqTM+3Ztf5Ah5/fBwpVqDtnnaqt0tobUj9ohIiJlbgxx9NknSl
kUvq+XjStdGHQvqieBWqsuz9pLR4pOOQn5E2z/zdEQodqIM2S6FA1Ud2UeM3aYnI
nZE9hd8XSaTmAg7MPEMqE6qETeG8JTe1SrRkZJCFLzqnVwC8XBlFC7BMuGuGJxgr
wr6l4mDxD3Q0VyE+bkinwqQQkmJOuIrvSnJI5yAgYPUcKIpDMJXQ8Kx4M61ur2Sq
Q3/bvNr9yiexN4u2prxnj5bBUBz/H/gEVdzS3EeJtTSdClaffbo2gvb0tY0nFiUW
FNXOD3JgJc70Lg5RdU6QLJNUVpqvMzihnOA9Aha7yK9Wc36yPBi7nhwIKWNzZjLZ
PHIx2T+4q/V1rwOcFr9+8wrWx7icVo2tSuLhgOllwsTcZRs+s5kRHXrDWZhA3R8h
b/kQYpBa/+2pyXtAymbTPl4TuymRoTR8xfwIFDwLrUJ2SziKb7KMU1ZogjtfINaH
9kCZnAoEkjp5NYMidwnnR8RQx+lG6atW2JJD4XV8pwodRS276Tx/N0KhJHsJ6fMk
1654IxQM3i7ptA4qvHJaw+rs215mQnqApPnlbDYpjzkcWpHz2RvVe6pD7z55N4MV
p7ZFsfwpMIg/9gg+n7G5kAuBxg2BrttLDbb3HfmIrxy25SzA8WZMYxCETI1ePdVr
52LYzY8Ruzj2MmFeiLu14zJSFsAVHPZ8kh1sVHwj7sMA6AFK8u993zRO0PN+3WkS
NoCNmIDPhQumAfCOWXGSXyNGEGsev8kTv6pL0qsFETPHyFWuS9KaW732PtNuj0zx
146w1LtfbO66yVbxQLDGU42UaLz+mnc/eEoBvPqszoJVBr/JfPP9wG00GZqtBb3Z
5q2sD1p3FrBvdbPCBY+7sW0wNCNAWDZSvJmyBT02mzvhySaVtb4zWJqtD/Azw0D6
VTrOa55xqle7bTZQSkGSm3Ksziisn/CXTLTmQPCDTxjlBok6vt2h9OJekFj3xrnR
qoXQvX203Z6Nv2TzvZjlCSxI5ILGND1U+FDXnEfIEnyJyhHOyvPTw783ew0tj0JM
VJnmOIaVKkFTdIUkLUFjN645QJZh1ytj4/zt/AF39FymmndChPDxaUq5HSTozd85
qRa0zjEK94hCLhejsHtxz9QQwqiWR9/kkLvrvSKjEoCjE0N2Itd5CzcAO6SsB2a8
1Ri+qjIHRyonZrpTbsj5CGOLQmrElbGgNXeo6Ncjeqkxgf6qKqW8W9XjZlPhlTbU
QzSxOSZDOjY0ID2J/tI1yMwaJwzJykNe0GnQ8DS/paoHUQ8zzf+cDOn7F0xVml8+
ium2hEeZn+wUTlxhI/dvtDh4eh3FWWLsEtePhGGZ5kpFZ10x7WVJFu/nBpPCtyuB
IdM38bZ5ohVXR+24XUNX21U+2W3X0GrucsbfgzJpg1DEBj+oxBsk3HfJGXtj+yn1
3vWQX4OoN2toriA5hRPF27DAUr5fxLiBLfEuI6XUncUlstAQnXapxSUcSxUE0Ehn
8hZTmH0WZnNaKNNns3RETAfUPlPRt573oHPUN8TbB0QL4YKzSL8uWeLshbKpVHr/
A4PHn9feNTYUWKYkskIObdk7+/o2QA83ZHeJGXsV+gHkJFGxUGgyuRP1Z78rljOn
y5CR8H7S//NatcvEGzHadM4H4AZPdlbxoh85PtoOvBXVPg0wW5eiCTOzmAdo1R+j
kgq9oOvupSiIDg8hyGeOO2R8QLBRqPhhIWwtF8JVIb3dyLaprHCm19kcfc2XExo3
bHRZsMXLIu2lqMQXJ0Fh4sy0jMejTgRNBchm1dpFMDivy0+Gkw6cXyDgTFJVuB9k
7Q00rgND/8XsIlcYK3ql/uZ72v8D+/7SU/HT+df3/QT7pp9baXSFlblFbFlU4kp/
q3zAoRIbAoUqz8H1JJYOHHIlApVMmssENky5onI/VuIkTsP9KGCkcg+fMAoRREAY
gGhZcYT4WrRkhCG+Rn50q6/I6NtghYdWIDnjbZj1293rzBPJEwLyUhiZV9kshZlr
MXSx2FssdBD8ukzGk1DIfsYKCj1Tt8EoWnCVPPHwL9MaJLTMKY6OhAThDaRxehNT
s3E3yVvfeByiqL2Ou6p4bZ/gTiFpwVlOlGVNlc1jmDEoIQm4+S8Kl3KvMCWwO4kA
Mv74mnvuZWgL977PV8++mlB/si7oEU8EtOQJslyzl7A55OmONuSKBGepnk3rYz8q
Z8/BwL3ALb3q8hUflHNialSv+ozepfBUyDGf2CQx4+JFul8oWsKOS73TNPs1CKHd
8lw+ZirKzN1uqkeEi8SZ8r3zADYzq1yL30nr6ix0vQZT288FlGLvPQsFS1vo5eBE
8zvAAxGfy91RxzQLYPzpjnGM6dIlagysqkOmKRRxFkRr2h6yo4455k7PfVD6/L2q
ohf0aIhExN87cOjFmqLkf3Y0a8FQuInrBS45pX8DAAzHqxqfAFNhYvmY6uiMqd5x
ciZp6WVjJ3I6GfdWo538v472U+l0P/aSIarcbmcHXYs6TD9X8l1tpwulNPZZEI8x
S+VPg83LPL7txOEMTDcrnrkpdrr6mdGsHVapRySrjsT7M/fHQLZobpPWPQ80UhpF
HWpBxlRWbGPqQ9UeteKvbXsEp0OZO+CEwdkwRRJGZ0cJb9Axo9ij2zH31gpMloT0
N5XCrbIz8QU+U0d98KbztqKazEBFfVssIS8s8WJH/5QKK5ZBvGkoX+VMAYEeZbhB
GuZfu9cjhK4VDx3TWc3p/zpYxGcmcx+7EGE90nblkYBaF/7As5xiOixX9DokcZCm
qLgCto1s+EyMPrNB8+4oq6JaR+hSXKS16TD0rCdYqufxPjd2yIWDA27t1yJibPkm
h3GYGgYyvJVdAGzSZtEnrm+Yz00GWpMV73gsDeO589JWwk70BPbblDZLAGuOJkq3
3Lbxv8ZCABLjakOmYhfGUo8lptU1CcMVo7HVb2uCfywom59W+eXhQIvJwaXlCqGa
s5xVmX99G8Vvx+vXeQO+W2lsgwsLyeo/DER5P15Mu2qxmJTw2K/M3eQKqNXGBEWJ
JVQVX6nBn43Gj6BHu8iMaaDQkqpbC8+AzIC2ZrMXOOPP/c/+U8bWA3De5r0fNHZl
wLFYxlEOa8w9DXLNZlBHASDpiFwJUk3zoD1hPCLC7HhLnlzn+ZCB+zIEjT7+IhzH
+KjRJ9L12AQZj8tB8UzPovfyTEFZVl2Vyy4gqF1mCWEQKb5IJBNrdNJb7qhSKEWo
3uJFmYH35Ddlc6356NLC3phUUo/wem7XdP1hcKd++gku81FxCzD799FB0kAAJLvq
LMQHriStl4B/1VihhrcLHu2VTvlq7LF82VHXJXKG11rIUDB9f9S+9muCDKLL0P08
Tau7LjY8dD/MRh/BwcC4aflmLBsCP3/F/3QoPcoUocji+s2CuKOq5zDKU0GPfWeL
pZYcHxk74U1gQj4EA/hqoV6+xQ/i3syBkDpxkHOMVJQT2CqdML1OazisJa7rx+Hl
RgRlrf48GxoQgJG1a4K/Y05zpY/jNbbn5fLnnpmv5fwIFL0zOwnRQryE4WQu90zE
2rRZjVpOtfAC0q7W9OVSmqYfhAhuCK5h2FFzGih4z9Z1bOuY4yYEhCB8R8U80Hab
LSET50kZSsA2A9j6mCkMVDjiONUMKhTY7FhwyPqrv74=
`pragma protect end_protected
