��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��`Qi4�)�q���+�������Q��
����s���d@�0O��xW��-2�a�J�}H���q4=�H��]�+�Ԡ�k�`��࿫��͕.P�� L��QY����O��I���_w,xkP���pD���JBD說@l�19`2�w5h��� 6����bթ�}]���s���E^�5B�E���ZN�>jr��I�["k���a ��v���ռЖ�Z��~ҧ>5�l��L�4��x�X��V�	�ANcy� y�E��s��h;f��[�DY6�y�p�l7H8ҝ���7�k�^ �58�u�U^�N��`�D_b}��*d Բ�tGO����~}P���3T<�&��7�e2u�~�g#Y���,��=R����`c�8��֪;�Ӏ�l�3� S<p���>(u�]`�ܝzCւp���q�&��ß':��,0%��.�V�� .!�ݒP�����<����VPb��~�����R_�f0?]:R�kh%<��d����ǳ�pk駇�$|h8�3�xw� (�_��������g"Ă��HJg�R4X ���=���W�pP,(���H���K:]���ړ�]�
y��2J}-~>C�:,�7��.g�챙���(F�T�Җ�H|~MǤH �2����:����/�3�Ù�uױ#z5���J���Y�;�Q���|a�1�űe2�z�1]�$	��3@��I1�OM0cOzK��`
h��X�T�8��&��.K�{��Y=����Y_��g�9�D,��Ph֪>A�$�T�$�[�BZ���$�agZh�EJh\�i�ʠVr�s�Jt*� !�G�m&��NI�#QF*���b&�*}��
����s�FY§*����1 �U� j�tY���퓽W�}�s��f���C�	��A|�.� 0�GՏq��כ�*�^���Yd �u��%�0��#�h�y9���7��@���V���H֚^�EM8�8��%����15�V��R�p�M�:���r��:��s&�_"?�%q���JlI�����w�����ǿa4��L1��G���WF?F�9�<M-�4	`U���O�X��x���}�.�1ar�����(=lΒ��]��h�|��>F��B��RB��i���!���ör�nz"�_h��m�d��C>�~V�ԅ[iw�|�����P����:_|�/��oT3ƈ��;g�JN'��*wϲ(V	*c��B�U"����Ѐ7�>�7l���#KB�~\��t����f�|L�~�k���]�<:�dx���r�¸��f�ۯ�&�� ���١*bLUL�����(�ŀ~s��:�夜�T t���L��T���]�C��:����AS;�M�#zS����ʀ�p�)�Qr�z䁦�R%������3�[�2��겮(�Q�p��ܯ��cy6ЩAZD�R�˺�^���P,�r��K�	 IrOw���C|r>RL��H���b�&<�U���%V��r5A'����?!���e7� �Ἴ�n$�_���.|�R
߇��t�&��QQra�m�~M}�q-fJ�����E���̏�:���F��fH�t���m���XU�¯�� .�b�w<��H���Q� A�eG�O?p�}�
�;�<G`�2�OC���������*e�N���,��i�9Va���'?_;�w��[� ����j�?r'�Ԏ.Ǿdb��`�Z��(�T�Ej�w���L�z,��t���h�
��R�	���x�%m���v ���&���?�K/����m����@>@p���Ut�>�"��`w��g���Oe�V_^�#�e�dH�B��8]��+�w���?`s�I#.�XZz�'uWۯ�;�^�o�B�No������]�rPE[�,�����ޛY��	�ni�6�}��7$O�8&�e��5G���􀸭2L"��F:�$4A�%�C!�D+xz.�9=���#=8%<�go��M�2����D(��pb��S��<e���!t�O��G)\��)-D�rg�@C+��IT��>�T��Ф������z�����dg��5��j�(�l6 Tzo�E�+Yo	�Y�I�7�w����!1*���Ia��{
�i%Gy��}��Tt<����5�b+�`lt"��G�#��ć��d$~ف�H�U�vV<M��b��&3��3z�$��(S^%���?F��e� �q���q�t~wC1C�ʖ�~+˦BMK���e! ͱ�*�>8Af��Nb$�g��� ��k��ȼ��Q����5���&�f��n*k�f>�|����6P,E�f:��s~d	M(0]�d���-eZU��I��?Y5�yK�5JB��ڸ)F{�(5m�Y��������猋�q.�r8J|\�aq�J'�1�3Փ.�&�)4y�F7`���e�b�o9�����F�j�j�:��X�O����TY,=���yI��F�@x�c�����ȝ�LM������g#1S�|��q�������6�.���ҝ3����m+2t�i9���1Ȇ��!� �r�j��q�I�ڳu6��#�2Q ��8��' c)
m�������FW��ǒ"L4��bd�gZm`m^�zQƽ�����z��t3?�|��x��'8�$�zˈ.:s�dv�	Z%��~�,�gs	KYL����C�����κ�޴"�bm�zV���I; ����fW!��4E�5��!ـ����e��		7���ZpC�TV��Z8�h~�ء�*��ѣĝ���+����\�5�?�="��d�tx�H�tlh8̮�:� l�w��5�?ލ[neG��G7qJR8���#���=?����q�H��L�P_r��	��̸�'�"~;���>d{�I0�x�|�"w	s�>��EЄu�\K}%�e��l|w5
Ag*�����hi��yS�y�*X�h��9�%�g�)aBܻ!
U�3��@���I�Ss�*ĠXz pg�rw>�Ͷ�������wv�d,�_I���a��-1kɰ�٤Z�嗸��]ʏ.�5���"9yG��ݫj	Ĥ�z�Xt?\���ˈW��<A����r�6?��u
=�B\i��2x�,4��Y�ᯘ;`.k��e�dH'4�y�-����{*��Lu_��>��ؕ��J�'��~����~����d�)���q�[�=�{%ToR��M�%�#`Y�Y�k�o�ߌ�v�0H����Z`2��b
oՐ��O~��b�x+�qė�����l��ы�h�=�@zY�RmN�LVHj�|���A����=C�f)fT^� i����O��ɁV�tI�@fH�wW]'
�(���"�([�G�o������Qq!Y��Vi8mQ�	�Ɗ�G�)3LX�|��B��O�������-���>�0+�J"��k�r1�A��xFY�N�������]ؽ�	2�/�I�{Xf�錘�#�����*7�_Wi�*¿1��iW�豨��+<���z�J��.�T��Ǚ��/�_pX\�2Z��g�����,�TE3�T/���v�5�1��LybHu�v�9M᜾�I�x�wu����,��"��>Q���
Q�6t����-u�Z��c?.�R���Sgy�l��EU�HO�*����U�W��1�$������lw/��mZ_�٬yqW��,ڸ�;��xh�O�B4�,��jP�w��Q.�h�V�|%�Z_��>������X9���e�M_}\;R���Єa���ž�ۅ(cӾ�@4(+�p��)X���(�����{��9&%��W����,X�V�"*��h<Wf8��.������8"%���4�[�6T�������Jra
[�_��~?�����b(�Ǥ�j����k�gm�`�#msw[f&+���QF�7�(ef��Z�Թ�*v�yx���}�s�l�zF�g�mT��7�����4}�4���GǦRFY2����B�է�*�@�昺�
���r�Y�X]����^�e?u�?q�A=R�

>1���x��d �9'ל�щ|~��cc��;�Bu��/��k���H���{����x2E�fT%o# �H�lC$
_�d�̙�1��p�ڌ���6"
��鸊4V���q�B���xT�[��������w��F�V$��fs'�"HvjY�L{��_�>��}	MV�猕F�o��@E�*	��e�D��/�=G��G'r��� ��X�o���[��գ*Q��I��ܰz��Y|��:���Lhգ5��7��"��Ms��W�L&i[�Q��F؟�����r!_j�C�.�Ɔs\A��(S�c	_(���+�P6��]�wH����U<sZ^L�=�g��G-	kD}����S���<G��PqG�����q|�\V��س�t[�bgUb6|V����������n%OG[�y��0�.�a�x]�1���R$dIo�-q��l��7��5�û�.TU2<;ͱ ��S� 9��!Idm����};8f�Џ�O�� �=��Pk�%
E�����.n�7�C�ƾetR��d!4��]�'�鷕��8�ZW�8��
�測u�D'l��L��L/���W���[�|uT�4��v΀�,�>5���~��R@آ��w&6��3�ef�b!:]4�x����ػ������ZPr�v���m����Iƶ U
s�����R��l4��6Y[� ��=���4R��/���,+�F�[L����a�!��ztI��Mu�B�%����f�����fP�/�JU<��[G��8�w�R2
}c��X�A����^5Gz�o�m�w�>=< ӛk�R�~��rr�惛���!R8���L���k�"�2v{Ov럆B�}}HՀ�䱰S���[�lb�T�2�|;�[�Ϸ�Ce&"߯Z�m#�݄׺>���V^��jc��9K�p�gdo+n	a�5?T�ў:�;�ND��0f �A�!�Ur���eW����Z�L�S2H�*��B��@�'�
�g�y�K�<T[TT]v�L@P��r_ B�����73�
���_�I��c?�04P���(�Ξ�	]�QZ}�^x�Vtm� )R/h�4ńe�\�U�Bݞ�St�jl4��M��պ�<!�K���|����g��^�:&��?�� N�m�_��Ş�M��GKGY���頎sKV�2�C�G�n�	�iu�{͑��J]���3�,@֘2�%��'M�iy��J�,/��⾘|`i5�&˙����8�$���[��"�86�VU{`9����}�;Nc��A����<�Nk�h��v��j&Ư{=t��m_L�̕��4�G�����z��a!z�b|p��'e�g�Џ�cή���#H!�tMU���i܁�����F��ax�g��4���q躥�p�|���,W�#��7�>���}��r��qc?�%]ÊW��Ҥ?�C���Z0U��I�.�{��Z9���&�8�S���.a����F���^�dd|��:t��D<%4�l�-,`�PJG�ğQE\%Ze,�=z�3!Y)(���u�t�ѵI{�m���_�f���#U�3���=<��End"mxm�Gr�$�$�+�Ҿt����st��E꼦�L>�}��OPF�0]��Ӽ'j  0a*:	�G���� �.Ѿ��	��F�O�������UI���{��眺��כ,l]J�,u��ݶNQi� �*A���>���?�]�Toi`E=)`G`#���gW�����Y�O�h�~�����*�&��.M��)�Z}��R���u��<!f��g폊�����
�-�:Ğcr`�Օ��R�\PT�I��Zk����Ө���sT���G?;F�<�G��ނ9��^��S7�\��W��$%���	=�ce��5�$�aT13>�����z�zҌP�z��2;h��[���Be�yE��x��ʴ���o v^��M^����������M{g��������A��qF��Ys@�w5t��|K]܈
��ւ�ru���w���BФ9���-۹�n%L�!ǴQU���0�=[�y쯰X����}�Co�OSޥ#�5�v��a���T-� DD4�?�i�#'�����ׄ���x��6�YeL@�[���Bg�"��,��.$|n�C��1!��TB�N�_���$뗼�b"L�a��O��l�^�/ѥ{�[�N;c0`Ax��Hg'�F\{�ف钨��Q�&W����N>`���l���q�sG�O��#�2Օ1�0����>�׎L�E)����75�D��	�;�m�TC��s��b��y�hHB
տ��d�&��6I�%��97;�K�;�!����8-]���
[��_/�I�w"�Z\�I���zb����,{�Q�3���xk�.�g�z�ݩ�i�HG#T�V����u~�vA��ڶ�E3�?�����)T�ۗa�>��̚0%�UN���-�����$`<��G�8w[AO�,)tY�[0�`4~�����
2��Y-��@�k0oE�'�\��d��^��_8��@`��Y�5�1����)�r|K�7�@/i�?g��8���@DU+=��}��e!	� G��_���ф��:(��\���	�/��IK�,�@h����>�� �.��I�H��g��Ȑ
�������8Z޲�l�`�3/���5��y���lC�5<LIN:š��W��p��;/��5��ys�s���bY�:���H��<�)���0��%3f�20�I�V�Nx(�c���5+�%'��o�q�ձ�$X>ӱ�(L��SӨ:�׍�^h��S���L��n�\����P��+�Q�����t�h::])��FFPD��V(@Bd�.T��pr��B�?�(?k�h��d��m��3W�1|��i�t��1�kU�.�9���j��"��P$b7�A�H��Mڊn��cg�' z�y<t�I��H�P�>^N��[��[|a�޾�O7�X���&^6�`K�ҍ���p#d������ֈ�kF&Z��yH��U��yEC~*�A����I�Oo����c����w9���-�a ɠk9%���S�LcpBx�6!i\Y{:L�X,T�u��� ��}��w�b4���+`a�{�
+��+��Sf�S;Fo�^�Ɣk�[�I�̔�h��֔����a�v��l�'؆�.m&eT�"��G��[����McE�p���I�@���)q
4��/@ҡT��ֶ�Dy,b� عo]g�/��2�aA��u���}�TÒ��FPo���`!�{��)����Hu���q���	)�h�t��p"�2۝�����&S�獘Yc�5F$���FTd:�3�x,-��IQn�Y�=�	�%�9�����Mj�[�ͨ�>HB>?K�!�����y\�Ր���>�F^����eIs��VM�$!� h(6ї��q�ӈ�A�z��f7Ir�������8�~�T�6V^6�}T�(�%>�z�\ô"���Z���P��X	� ��l��dC���y+'	Z=�ƠF������t��s}�=B�o�S��	��T}�#���'{1���� ��O�g���@�f�?Y�pd��<�Z��\�� �����1�}9����������Ul)�~��A�|�c:��X�Lz���j�ѭ��J�����{0b�z@_�qY�ۉ���`1�_�b�˃	�_�;+�Xw<*�"=j̉����ֲ���	���bh��X��ы��{��7־5Py���Cdy�L
���\���5X��9�%'V��OZD8�����p��C�����g�B�g��+f��s�b�"<j���f��1W�Ǡ6�Ɣ���߰.e��kqڑ���� ĥ'�]]z>��U�i/�4x����c�3L��i�D���B������-��^JEūV1i��iOd��Qf��z�0��a���&ź�׆8���\��*�L�:�M�"�蒭��1E�T-Ǝږ�&�r$� � =r�ݭs�>syX��0��-�������9I��#D��r<�j�v_D��_y�F���;�*l��GhƱ��Ʉ��(�ܠw�|�L|��y��ƚ0A�>�gbB��.T�
REā��3,3op��h���.�v��X��3�Η)Z�����#KK:��B�������YMń�ɗ,
�[��i���nb���@��m� YW7�d�_����"�0���?���D�j�̨B��6�^�t�lS�^����>\����%ξt�5b��h2��r��Ԃ}�n`f*����Y���v o5����[ʫ���9�� ��R����PN�� =�+�%@��e�dD�޸��l�SƢ<0�d���RS_{�/Ġ'�j�Pg��i>k�PoA�B��F���s�4w"�:�qn���G���'���bS��1��SӘ� 9Jwp
��>M��B~�)��|1��J��j1$�5Qj����Cq�'
tEB�QTm�|*Q�ڻ�S�v���	<�:<8��JZ�P��PGhly*{F9�T�jMT����V��2�͸�d'*b�2�}j"=35� _��2z�.�.]^��m`�B���_�A(��~A\58���Ҳ�<'!�>�\���_!j���Sl�$��}�d��Q�F�D���22@\�a@$�f��.Թ[�G�Ms.�Fȑ�e.���\0y��26P�s�4��._���)Y�3�Gd� %	! h1���Cnw�V�����C�������%��yCf���}��qzBͽԳK�M��9Yr�G$����.�Ic��)�^?w?>}� ][{�	O�T�x>�;�,1�ʙH��Yd\�d�9�f0z�Ǐ�c��U���&o�f��p	%7oQ�ߔ ��P�|Q?��5����z��P]�7�~yD��Ƒ�\ϗ妋�ꭝ�Ĭ��9bd�*��}�z�=��R�	���^��v�}���&��ķ���D�L�����Sޏ<��Ɩ���ު!��2�����Y)��	D;��2,%:k)�Wb�&ҁ�Ey�-)�,/i�!�_ү3��_a"ob��H�CWJw��Ѝ�����F��b���dl_J�#9m5ΛO��|2q%��5����kВ(�B���H���n��QLl�}ם��N��&߶ڸ��&�|؋/�WtGw��݁��0��Q�i������Hǅ�r�4���E�T�'Y��� ��bZ]�|,��i}���Y��PF,����:=\���4A{�6����W&� ������B8���/��eq���/5�4���#��H��Qh�,IgK՟��~>�+AQr�ǘ3���bM el|Ǽ�ѩ�Ln<\k�i�����-�d<��v�e�C`[(#CR9}�=��y�E��\�SR��F�j��)����!���[�y�枹T/�z܅z>4����)�>AL�!q�O��fU��4���
r�@Q*�� �W��Xj�z!���B� ���Y�����Ȉ���_�Z:}#//Y�De�i0n�Ш�}�=��YBm7���dz�آ��1����葇��IK���$���>l �»7��tO�J��V��VA��#�mQ�����A})8`H����=�	?�!�w�#(nw��j�Ml����}x�n�21�]P;/��4�A��a%K� ���\(��,1�����eA��Ω�fck̮��:�X)��V��25��QK�;t?�D�a�Z;����3��zw��c�E�T~J�e*�CN��'�D'��~а�(�(�J�&��c�5�3ޖ/�hF�֑�n�0�Ա�}p�rC;�	����qw���U�!�E�`��?�i����
�>{��C����JM%x�%�����WlhFm �/=N�����-oa^�X�L�ֲ��""]�>�#
����%E���@~�/��5���R���L���x��(�@�e�EB��-²Y���#~.��A�����2��v�n�E�6]PO�D��~J��#�Tz�,�e~G����=9H���|Q"��I�&���IK"�S�"m���ʫ<�%;[o�&�=������1�1�O�93�������'�uǥ�+n���տ"/���X@��?��VX޽�ur�4�a��	��@����Wc>��/0��Lס�c���/ck�����U���n8�i.ϸ)ܭ���f��L�&�M�H�3s��e�9Q�3ϰ��S,��b�l�C���,h'���r;�lk�gS]��S���oycU�{̵
���}Kq,�h"�U�!@�*t#D�%T����.�`x�C����+)+b+�o�|�L�3_�I������`��gt���7��n��(��ѭK@��n��?I�G[u�kCƹ���r��_Z�}����N�Ȋ�L�Qqa
zC�,�m%��M��=f,#��T��B#��N��f��]TF3_��t�!t�UK��3 pP�
�5�&�e���v��@���fd����}��5�[�Ry���mTV������*���?�� Ix�����!��>t�:��=�����9.���"�j��*���_tP���NƵZ��c���ݼ�If�0���6���n��C陴��9��Z3G�;�,<84��?`M#m�i]]xpw>D��Ƴn;�����`��Cat������Z�}:a3O�k��A����b��4�XcvA3��BU��&$�6;M'	S$-Z�]����|ۢ���A�S�f'���c}{�
���k��qm���D�b���δcyC˅�����[�2���S�2U��+����E�Z�l����������k�s��"]�7�D������ٴmw�"5>�!���6X!�
�����$�%3��܁�'�'����$V�+�R�%�'uvr$��ɷ��f�өZ�~����LN���^�W�D������-�l����f/���ȉ|;�,���NG�03=Q(�p��S�рc���:m3$�l�D����f` +i.�h9 ��=�ި����,8#D�v~�{�q��h��Ɗ�iV�=8F������v��(�!�.���4�H9C� �r����X��P����0B�Y�f�K6x���N�4{I��T�:_���X�sx�
�vI�(���`R*mM����Ȁ�d���1��ɴb�����Ȅ�gaW��Yz��D�Ӣ�~|�o�l�=�$�p��g�Sˤcb�"��R�o(���?��ѫ�(�M��MVr�c���}�.�.'���n�����)��0m���{�W���6�e�A���^������}�VF��>����D��q+��~�R��:i?��6b��TJ�;��W���:p��JS�_ǩ��D����.4��e�'4�Q�
��ӓt/WܴLЭ�9m0�܇hմ�}	e�<�� ����"&�KE����)f���co�3�����,����|9xM��A�&� <�f`�ݡ�?r>͙�7�`�UgRҹu@��[sŃd\�]N6�c���N<Ѯ	���(��r��lR�z�R	����D��Ѷ��BvSqe�	@��b�ư³�� Խ��'d{C	�eNxss�3�i9�EE��;<,�m[��'�2�����la��H�d��v������<�=�@�dHI)��[��*������f���0��Ph#后���zz}��?�z���d����W��Q���wv+�>��1)2�S3��=�`q�i�&�hAb�Z�s���r�e�&����A� ��C�%Wi�\��0ஂN\�����FH��\���)d?es�����xd��xF2`d�E3���0ӱ���Wo*��Q���;��	K:L:��%�͋}v4���q�EN�Z�����x�>J���aJ��]��
��@��E���(���Q����	H����4;��ŢO�Ɣ��4ڙ�EE&�ήQb~{�'�ܖW����i^N
�Ώ��S����Ј{��L����I"�:�T��Rֽ���sXH��~�C~V��ޣ�cY`�W`�F��)ya��L�;�@_0\�������%����mp�>WN��3{$�'v����[}�.��,�n��]ϡ3��G�`ĉ�6�/�� ���W��n��H�y߯}��0��V�M	�7N�7�@{�`�b��_Z�����"�&���3pa7�j0�6�.�\�X��>�� Sv݄�ު7G�e��Y9���h�)2*EGp"y5O����/X��*�͚$z�Lvh�b*�<��Rg�f�z�O���%�eO;�h�GM���'Tiu�wY�-O��w�*��Љ-����VanK<O&˔Cņw���#�#>Po�W/���y��N��ۨ?�?We�Q���˖;TX�`����:�|�Xĳ+��|��L1I?Ŋ���2z���{#��?	�=C�N���R'B��R�v%`w���v���4������i�"���a�'x��'��n��t>�w<�x��۹�G�A�*v��0:��3�'�����	RVgA����������+�B��h)b����=*���1�n3o�~��&�j��f�?ƀ��G%�c_�Z���e��c�s�-�Ѹ��2����/�:�;c6�qf�l�e�T���z�����-��7�#�,!PnR��[�ݣ���$��y�b2c~}[)@*�d|k[��	��)�i��E A����`�[�D�}���:��m� �9�z����$��M��?���h�� ���w��X�xoa�}f)��%[�)a�����/h-5�oO�	1��|?p�^(���G͚���sΗyIrֱ��/�O���mG�M��wk�u�3�VI��Z.���AK7 ?��``6	�B����EN�L�ܣ�u�U�bP���$�e�ݚ6T��d4�/��ّ�7���N�}�D8n��`��fz몀kS�!��&��&~oL�"b8���?`�M����u��}�hL�;=cݺ���7h��
^>��F�@կ�G��z��W	UKۑHU�Y�o����@��6��\�����|�F-���zK_p|���.\��ek�[:�>��-9����l��L"��'���=
������u�)�-�Ղȁ5e�?�V��D�{&`s����ey�/�S�]���5����S=}�,�THB%g��8���ҥ?��/����$�m	�j�	ȃWV�~�%:BT�����.�L~�:���UM��; g@WX{�φﳶ��t�\v�	���� 2xX?�!��SlRk��O3[��:l5��;��*G��%K]��i�4���MG�D�^{��,��4�Y�q��R��*G��@�����S�b��ܛ�Igݬ<�N������#�jǷ�G��8<y���U@���b���m�c����FX��t�V#��DZ�� ��^�1D��B�q��e'�3�Ac(�[�r��F`h�s4._y̟�Q�~D@1W���7���n7YA=�� FuV]G��\�N	���=�,�B�W�&��Dq��|`֛Q�1V�M�[�и��O�Y�?n 	���n���R�����_i�N0��c�[�����,|�{G+=���M��1�MI�mB����]�)&�wL�Ѻ�C�ek�lSJ|U3m�rR2�N�u��ªλ�6���DIi�+��ϣT� Af�J�����oovf$�hx*yP��|1e�5(���Fá��M�3f׃��\��v.$E���ˊ�7�7E�&��1��,7]WAw�����l�� ��e�Eՙ�5��c)���c������m�a(�mN2v*��S�h���Pl��ϒiD�NP���_I�}9s~�G_��d�$��]��J�MWIGn�0��g�#��/o.�{X=��1�Njk�S	O�F"���s~y���%c�q�kQ�b��z�~�1��ڱ�,hh�ws�%�y�Ԥ�i-0ȼc�Y�~��&Ƶ�2����Xs4������3��j@E���c�`���/A9��@<sU����!i��V���~�-%�ﷂ|ȃOq�7�Y�;�7���f�k2������j�	8v��]�%��Za��$y��o��c�b�b��VD�`3~��-j�Ye�GC���<�g��<�G �E�B�ɚ���W�VR�յ�;�p�����*6�	�Pֲ�'0ɺ	�[_��W+��G��Q����y�o�u��>ޕ\k�LV��RH�� ʀ��Ɏ뎘�L�2���1�t�V-X���� P
Xvl�f�#�d3�$��7
�m8��������J�V@�(#2g}��Ռ��䔉����+m>M������AćUԴ.��z	C�@،tVJ����T� �n-���3sG�v��}�ʅ�����6��z���ՉU�FV���A@/��8e�Rw�%���z��_~�4h�g�9��0��\O�nC	�d���ئ�{qP;��z�v�T:�>J��Zw"y�7�h٩kE$�Z�Z��j#]�#�����u����� �`#�A±���7�Mz~:��c�C��"�s�:(�9b�]zLi�G��^�vUKx�4}��>kdҤ1fT{)�!�ne�B�U�U��[ʞs����NC2G@��6���04��9�u�*˾��u��D
Ϊ?�U���evq��t�	iqZI��4�i�T�H,�T|���vV�Nʄ1�D2�ҵu��Dfl�a׿��+`8������ۦ���"DJ���s O�Sj�Q��b�g�r`�����$��n��.Z�s�?���ǝ�F,Λ/�x�� �r���'n"}����D��`�+J-�O�zZ?nos����vqi�^�g�r����>�_9)�Fۭ�_�#����<e�q�
<R?|��ϨV=�q�&�+d�j?�W�� ?j�R��^�yp��&�0���zF;(���2ƊP�
���74c��9�KԊ�춦�T�xn�Z:�${z�	��q���~r漅����L
�y�e��] �����	п��������;�F��g�F�oX� r׶��璁;������9l�?L�έ��߯�r+o�<�~�j.���L�X�����&Dck~g_A���iX�f!��G�G	��F�pQ�*	�2�ݺ'���I�Y��
V�G\*��	�g�f8D���+���حΩ6X�r֌��ye���ɍ����$��M�}#��:'O|*%&�6�vϦ)��q��yk���s
�s9�n�rY��P�>W�~���h����c�gu7�� h�1����Z�?�KZ��u:c�N- I�u�qyiZ���Z�v�C�F��1q�M�7fTk�]��G��U噂MN�}4Ԯ�_`��9�Y�����%0�}j���&?U����+?��W�q}�Ã�O�2��%�MK��Ks3W�>L��b�}l��:z�:[�IR"��H�A\�zc2��6�;�}Bޏ���ah��ߟǆ�����G O���8t�O�3*�mԛ�V������+*�ɢ�����5��]�ٲ!�@��;@z`}y���	ۨرM���J��!�-uI��EɋJ��/��KG����Ő�֩� [�C�\���1�mh�Ƙ�n�śT;�}$|��X�2�h\��g�B/5�&%HSy	����	ɯh��~cA�CXW�5�#Ҍ���o�zb�6/y��.=um���D���t���Ƴ�˜�6w7
X7�~�8yu�,`���$J�<wy1�Mİ�I��m!g�GͲ=��}}H���!4�mB�V���ߔ�r_�x󇞄��2��L��2��?�����!�����zB��}��T߂C.|J��'�	q�p���K��^˩I͔�h	�&x��/p�`Y֭�c@ɘ!�)3�y?���;~�N0�7k�#�ګ���]�2axuЖ�𷐽�sp��YZ�7[�T��Y.f�����ީ���S�J����7�n8��,�^�H�O2�o�T�|��]���_|�=��@,;G�K�, r~`7��24+�R�N@~8�L���g��i�
���]s�~[�P�(KIv�f��1��\�}�)��m�I:�߬��xv��Mwj��G�V9����m�K�롤h��װ�JRv�Wu���O��H���Rx���+u0��ۗ�P�^�+\�U"�n�����0�������(G�ai7�C�nfn/%y�(�ʢA�AWY��V�W�T�sn��I^���n�ņ�A�W�WW�8��a��Q<���2�*[�db܀a����R�+�L�Dj՘5i/[�K/"^��9s��uR劗�z�����J������Ɉ��Y՗;��*���d�P�������c	�ʜ.��l�Q})��C\:�v!�����!Ō<\�i���X֕�:�x5�oў����;8�*8I7�ʩ]��| ����#�	:y���Q,Ma�7���2��)�p�vp��:Ɵ�@��z���
f.�vK�/�����U�,��Jj���xu(��~������j�9BW/����y�Yz��ʚPk.ci+��g"(D�'�mtB��r7�Y<�<�Bu^�+84��k~�z�r�~ �:��KmJ,���R�jo��0�s��1S��K�\�_Jq��{�O�<����l���.����{��H�����nV;&�a]Nv\-�=�3
���-Q� ��R����cRr�Y�E�c���f���B����5�ؚW�����^eS��c �(�PǑ�C��d��V<$���E:3S\�m�k�̧'�L7�j��d�5�Ww�|��@h�9�<�F��r��7��O ,�y0Z���p�p�K�-
Ӈ7�}�qJH���Ӌt^�gS��!���;�vA"@[Wp���^:>����f?\��p��QB��hQ��,����QEh]������yz5|�,��;4D~'�+��?���}l���}WB��d-��g�gɽ� .t�I����j4қ�\���1���DE�Ⱦ��P%8@��޽<�h|�I�I�P�BvfUB~�3`5��(���=���A�Ap���P�AƐ/�h'iW{��}��7�����(��zE�#,�ž��\���f#.�~MHtt������/�Z����`1����w��W4�EP��&�X��U��z�y4,C�mт�m���uCE�	�/�AC�D2V�@��܄��l8�gd��giʝ�c%w��?��wԨBl� @��>U���p
�1�����f��޼�n��|�F����簝3���J�5B褹�⤺�����t�iGA?8�{Bc���#:�Sf7k[����֯�Q}�n@g���lU �V����3.ĳ�{LH+�Ԑ^�a; "|	�7�L22�5�i��%��^ ���+y�����Jw3����C�pqj2��b��}�|%β��0 q�cgBE�nenu�3MK��ޡH`wD��}cH�o�?3��/�N/���E��
�4���.)�U;^���!�4�Џx:u}�O�i�K��)u��w".���X�G_>��W��0�2{���&K�u[��9*���i�F�ѵ��>qUZ�����@�
4Q'���&^<d ����"-��A�fleKr�	g&�����.��#� ��d�)*`U]AO���P����A���B#�B=����gE7Y����n��Y����A��Ca�e���s�Kn��ZD�e&����2���g�{(,g0�p÷2~��]��fV�]G�d}�O�`�+�?�z|�@*Nx�ocn�2y�^)���E񈔝���xa�޲/fr�n 癥n����C�zK������k.�}8��͈<�������
F�VVwVH��LDE��|?Qh�BQ���⩡Q�Q��b�J����8����g��4 ��
иc�!��{���c!Ur���J:���H�㴾m~����`>���k��y�_;!�2��"��t.H��Rg��@�H�M+Խ��0'$s�,�3|��h�y#��c-�	/�Sed�AS��9ƕ�R0��q�����,#����`���;Ih/ ʼ��`�*�J"{+�ZY�-�*칒r�ОR���˒ok�觻)�mռ��[��BkAȬ�^��r!�`Y�|��@��&�ܞ�UV#�J�:*< �%K����!"12����t���
��1���?��[2zS��/��y�'f������r���FZ���yDB	�(�i����6'�W�]J���6D�*lH�pw��I�G~�c��E��!=醡1\r�{��)h� 
qv���)M�E�/�	mq��yB ��	I]`w�)SCS�)�p�����m�)��cV,��k���~��"j^�4��f�h_��@��5�6�c�vt:�-?�e*l_Ϟ����Mv{��`�n�-M9��]\)2��^��fa�ވ6y͍���#�T@��@r�s�����P R^�[�gTi9�,��ٖG��9[7n���Ҍ���B�]%�6]L{	��B ��-�9��t��cwj;M$��ɘ��딡�|���Y�vzm�Vƣ[��{�9_��>Y��K?T�t��&�fN�8jy�tA 3ꡘ���T$��6:�@��;����9끫4�<`�Dܳ���ޟ��\�%o��f9X#Geh�W�B���7��!�5(w�5��|
*��u���*�A=�����,�G�x;~�5�si�oja��F�i��֔9G�p��-4�*.�r�;��r�\��&���ʤP&�����\�,᪤�˗f�y���\��[�I]j?�|�BW%����L*����u�D�{��E�����G���"NҎ�&�NPXhs	�?C��G�e��8����P����	�ڏ���T�3�}����0���9FP:�8��ns@��8���x'2t&�E���C�H�ssU���+u� ��HU��6�fx�P����nQ�u^��P�jaL�"H�8_��s��w�
3��哤��T�����PP�#��T�(e�ȇKr�˫*n�8�T�éI��o�9���Z�Z�����t�/�Qy�j��R�f"��S-s��)�)��<��/m�nz�ޜ씄����#��ll�(�B��'UR��O��m���]���S��-/�4�2�n��C�91�t��5�x_d�-�c� �����Xgr(}f3�t�|�PG&W�b�:؊����CrN��3�l��/�:�����J��/l����Ua�o��ZG0�5��#����Ht2�X�F��N-�H���H1=�Z""]������c����QW�C��*d�X!�\���/�I�W�}i)e:�"pl1-��+�C���h ����*g/Hn��
)�vYNVL[\��"=����8��1��d���7'd̅��A1�(��Ì����'�u���Q�i!�xQ�PY�Eǝe����P��^�f}2w!�br��b��K"���V�)7P,+�ƍ���Iqu���55����WO�����fè��=�����k!j
d���T�t�=��n�ٝ�`߾��	�]�O>6Rm�����t��į j����pI�iā�Ln�B�H��'_�?e�[+������� E���N�(���F���`;~z8�b=��y�!me�)�H4��R? ��"�3K��-X/��7!�+A��2$rg�Z-�8���{��o����0jr6[D8��> l�BÏ�a��,�"���;����G�/u���_���wP�2b����=�UN�9 +f���
� ��c�D�LX60����\!87Z	N!DG\�܉e`Ȍ�m;C՜51�]q�Z)��T7�:���s��N�k��m�jpo�ː��΂`S8���Ѳ8'�x�'m�.��$�K�"��6k���}���jΤX�	m�1T\�s#@��a��U�x���`o� O�PG���I��)h/5��\,�SNrN^�dDiQH]�y�a�`3Vo��*��i5�܍�UO�r�foH�� ^5CK��Jyv�m���z��r&�&G&c���l�[�Y��<#�9��`i�d&ؕG�����,���4x��ed�g��8�tj!5����y������~,���S;��Ҫڎ���\�	[k>R˨�a��C���?z�')��L��ϵ��iВW#�M��[�nyR�s��NP��+����d2Sa�h�;ٷ����g�KF��c*My.��{4HI��(�1��[OѻF&���R�u|=v������U�W�n��y��l�pn��=��ڢ�X$��\�5:��2�NM����~��ۥ�$g!���wP���;����n��9{w�[���}��J�z�u����ʓ�Y����N�_ܐ� =��(��l�����$�\	ۧ�C6e�����?(����G�K(��_���n����qzz��Vz�a�\��
4j��2.��q��#��ɚ����R���'L��c-e�պ�3Yz=��]��`!k�[�AW�R\�rTg�ӾI�,"R�FK�Z.67��7v�7��ɷhp�9Y��K!DRM|��D�����`@�1_h2�b��U�����+�J ���?�L���N
�|Ȭ,���Q��e"E21'��O��5�-�AV�)zZ��#� \&G���j+�y�c�7s����e�!-�p�KϦ�,��ݩ�Ň�o�*�lʖ��.4|�N�,��9��2ES,�1�*Q:����Z�'�$���vQ`'tX�٦Քz]����T�_�o�4�
6�g(�(�^3�qP���M���|FsX��#����Oe=��a8���@�F�^��e�F}��(D��bm��㽐��#���W��s-F���B��m�}�U�E�5is� f�9`�V���p$D��G!�R��Mw��\N�[�)�seݦ'L�S��>��Ib{+M�E�ʿ���a��~����~{_��~�8��Э� ���%DLrĀ�#�!B�1�d[%�𼰠�q�=b�<՗?�fǬ'b�����Rݾyr�F�#������_8�Q�'�aeM+Z������+�+]�^���&i`.(�� �3��]�X{��?��J�/&�����"կ(�Mɘ�jx/|������اnJay�w�dd�9��Ղi?2�,��@'V��t�i ��
7�e�\8��P����<�$�r���b���C��H� ����yF9Wk��\�<���S?_�/G�����X�s{��J��t�/�-�(����(�������baP��3�CTS��n�tb�P�7f�m"=�D��##��������r�k� L ca��]���d�H��y���j�N�O6)im�Z��X�a��)�3W��}ob�]�o����K.W���h,~J��U��XL�eĝ�p����3�ĭǮG����H_��&�<\:%���ϣ��<���h;{��pd�"i1~@,r.&�[���u�	�I��UӘ�k�*���֌7D���������m���/��vJ�{X��<9t�p��w~��U�[q�������Ɩ4�"��\���Mn����H}2�b����Gzx �9�az�#��!�>�U�������E��8��"%`\.�~wZ��J�`��6��$ɺ�{�$<*��83�h�g5��F��ǒ������z���1#d�$q~G�C��ۉ����K��Z����ɜS�V�t>���.�߫�C�o���I�E�zFÉbj$V7���gD3-��߰�ŵ��U� E\XS��|�R�!�Zì�E/�5V�g��v�>hG�����C'����	|ۼ�	u1��0��ӑ��9	^L��v�n:��u���YQ.��/cW[���+�\��g�P�]6��;�?QWנc3�ܮ۟�&i�-���p�T���՝�Ǣ����LF�aꙁ�k�p�d�c&mv�eA֎['�s\�����7\k��QV;=����њ@��B�vθ-�ZV�����8����Ζ6�]�DD3X��P��s�U���~A[�Y.E�gL�Ϩ�[Y���I���/y����®�N�	H���� ��J�)i7Y�6���6�%疌\[H�'F��"4�L4W�������0pul�si����#��������JY���d��W���ꮬk|�¹ek�7�K�Y%����[�T%��9�.,tM��z$*�>��*d�>�'� ��y����B�Pl}5�{���23�[��n�H#r�PnZ_k0/b7ä�=���c`nb���_y�����/�H����_�P��CoB�t͗��b�Jm%g �'X<�H ��J+A)����(����/������J� .��
s�w�a3�R`Y-lVzŝ]��l<�'��-�E&�N������a��u��c��#X}0����k8���u*�ݟ�bT�cH跍&)I�m&�sײXeO�ǟ�� �!�
=�����8�Eq���{�V�8�^6$>��A�������An�<���.��ƥd��Yt�h?����bm�=�u޹M��f�Z�g4f�,x�%6�����̃AU�Δ����-�>k�*`��>��{3c�e/2(	�$^A�G�:H�=Ҟ��!/�Qt�UQ1BH�P��t"�n|*�|Q�?�g��B�C�3+ǍNK�o�������y��Y�d`���HJ'$Q�|���|��q�Q�Rr�v';N|���F����@	�#R� 1ΌS����
�,Ƃ+h��B���Ɩ�&3�_8Tѣ��~	��u���D�8����ݠ걲K"& L>sC��=������ �I���c?[�r�ʿc;E �y)�Ĺ��zO�c9������e��e�{�z�k�C��� K�����Z/��)Cu�lv�"����~ܔ��|qU�\��".����̍X#��2��>��g���M�c�܂�A��b�ث�Ȫɚp)�V圧�VW�HbU��@�hGna�G����}'��4�/!Z�\TP4i���ٶG!_�ҧ�>��<s�.s�
�	Ǌs��,/��plW��H��P�Y��~���I�:�O"������Q������+��.��=���}�i�� C���>�?93��Ƙc
Ǐ	;�>�E�Q��^��'��{�~�����c��W��'R�d�(J�Lu�۬�������6ٛt��Z�k�e����+�&�!E6`�z����I��W&�u�JS��<�#*���[gd���Cr�p �ȯ��:�
@��%SK�}���x��W��O7
��(`�D�
�Ql\΄scs����@|��]�>�	eC&>��m1k�5��R�6�G�C<XUn�bn�ؼ1ET.[S�\�&͓��W	j�/0{��~�>Ҡ^Cd�E����mw�!�qAT�-��vj}����Hb���f6��#�<���Cl�w�V�E�q5R�!��K���!�\��|�;O�,!V&��W��\����˻�K=;�f�w O��`mc}Ӄ ���!��!����Q�Xa�`�4�7G���S+�`���L���{�ȗ[c���mr�Y�\�ǆ*4/o����O@|�`]��%�>����k�@~��@��g��A�N�s*)������U/�eȼPfqy����V	����Ҹ��C�� �Jq�g}���G~�aGp�%��[��P����H,��N���̂7�n�K��Y��\j�W�Y,�-5�g0��NJc*�޴��$���ub����3_��gC�z{Ԗ��Ik�Je�3L��������@|e��>6u��ty�	Zp�{��ޅ�s��� ���EJ,<��ͬ�0�3��2�оۑ�b& +�ʋ3��]%h�Ye.�[χx%?r\��!ߊ�~4����dgE��ч���Z���	�2N��{�KD���!�����5*�4��h�<쓓��1�z@z.�ױ��.�O���{���Ъҋ��\��Ym>[��ڦ��Y�鋛�[�R��?.�w�Uˏ�C�ZR@���G i��7� p&
��~'���Nb��B%���k��^x��>cl�K�S�UC�� �����X:6T�D��j�� �
Y�n���Ϗoc#��7����͍�s�k߻A.���-�ST[و����.8��y��\0�Nzن2u�X�uD�aSk��!��(fD�������H����ۭ����%����n��A:���w�`A(���:M��\����f"r������|K�/V�5���$+/�ކ��
QN"o��
NГ���#<0�"Ά�_�s�}�z�k���pz�����jj�q�Țw� �-�ݣ�Z����|:vwt�3ҳ�$Ȭ�5�rU��h�Y�̵#�\V���'�2$d�X8�s_�(�B�ǧpP�d��6>ݲ�.l+}*��-�M���U������ 竉�����<�D�'��V�)�ᕪ��J�6�g�[�"FL1^��x���Ȧ;.���!����Gh��>Bg;�r���Þ7H�z�V¾�f{p�A���z�63�W�(���~��Ƞ�7�o��qK3.�+�D
�k��6�v����CWKt�GaZnXu�8w�5g4����>�G�g�O�Or>��z7RtT�ӄ�����r�!+�L���NN�7�%M��9v<�8����u���%evx6����Z][�R3n�M[(��B#�B�i�ب���P�����)8�g)�<	�g��>�Q�.Gϰ�?���(�����+��{�(���д�Q�
����)����^l�
 �\߄��b���hRE.��[�hd���2�6��}��e�攥�2�:>-+s/߾��������@�v�@��ȳ�.ʄ���g���w:d�����ڂ qS�h��o�)�b��^[x�+;�����,���z\�]�&��s��S��m�l%�����H�rcw1���WfSw���&0�)�~on;�oxw�D*we4.Z���Mci��Ԛ�m���aGr���[�)N �� ��ʨ��~t�4��!�r��z� \u�T1���R�y�%B�e� ��^��X�[�/F��������c�1��ŭ4]�"���τ��x��˽��6k��ߙ�f�9t�'��N�7�%��o��9uꒌq�p�7���V�7�F���v����s������(���H^��Z��i�o ]�X��I)c.�Gū~�w�Ź���z"��������T��F����A�QM�1��w��l:�4��fWC�hL�d�BM}�r����M�P_	�Y�yܛ�5��eS��IU���n��j����!E=v����;Ig$�UTt���@$�g�)�&K7<�vY����Ƚ�F��R������R��q`uw��R�ݼ��D���mU�1���r*�:�ҮW��v��9	��c��n�`r�,�c$�C�&8\C��������/�������N�CZJ{��*���gf�cuQ{�u!4��C@��w�Ȯsn��1n]�<��4_Ϝ��\���}�ոx�($U&)��h�؂�5���	�<ZT�^�[[<�1��(�r���G.Ì��˱��~�j
�F;;v���e��~�t\�$��{J(�^�Ky�n��"�l�/�k&�z[n2a�HD}��_��ނ���qj����7�[�,9݈H��y�Y9[L��R���s쑢�(���sG��n����!b��oϓ�~x���#0W6��0�E/(Pt˝�߹1����I��_��9������x�<�[̬
����>'d(NS\�<��o���݃v���1���Hj�✖�fr�0�}���R� �GcE$ ����"2��/��>Ҥ֖X�]o$���.�T���Ӵ$��ۛ}�k{����p��
��l &�XW����K�p2����М'�TЎ��%�Sռ[�� ��"vi8�}��<��!�;����O��qpN���ܳ�+���s?��qbx�1���N�eM^(��!�t�E,�Ҋ��	R���&��1O���h?��\J��;�f��^N�ڨ	u
���\��yx?Wm3�-�;`��捗�P��/�z����c��X�aB,m����)������K�<H��`�%ux4�&8�ni�y��uwt̘�4���2D�q�UG�ӟd��>��m�7����w	4�
;[w�hW �6A�����J���4H�"�?��U�ۤ���j�f���T�YUvۉ`��( ��
�+��Q^��*��؟��C%ԃ�9]�.� Uxn/���U �e�N�#XXh�QO R�ީ;���Q�P`	��@z�e�0/�o&E��0vꝕ�E� τ5�6�k�<[�b R�� ҄����Uѓ,�c��#�ٙ)��u�������9�Y�{�/Х�D=6qp�p��
���=-�}����?�?cJǀ̺��D��P7�z����o>M��Չ����#�u�*����1,hX�����vtGw��"��=-�� �x��}�s�Ǵ��,BY���U�~���3�($��aT�n��Jѻ���]��4�6���*e4�8�,H��c^��''@;kK4(�?df\,�_�<��~����0��gN\��(.<�kE{�.j��A��� `?ү�}���^���`���	��b���,���L�4�;zg�^i�$�\�gTs`�����.� BH�+���>.0�ތ䢿�2^��i����3\m:%~���>�n���X\;���9�f�\��ԃ�<9���:sု��H�|�'��^���G�}�,�N���(mO�+}�a�L��;�z�Q�B��1;	 3��N*C�Đb7w'գ�:�����4k�)Jxj�Φ]Q8Z��o����p�3�q�u���N�E~�}"P�E��]��/t
?K�}Tr���\/�_�؈T0'PG��O1;W��Xם�������f?.^[��1TVÅT�	��(���7��`�'mJ�C�Y���h׿�F�i��o����J-���:s�˒۸
.�Km�综��m���L:L���o�3�P�zi*��pP���uth��>ώ�,A�+t]�9u��Rꘒz��邗�=�gLO�G�W��5�LP�1��],h�N�H�U�j�{�~y����kll�i���ʉ1vm��)Sp觟ƊU�?�	�x��\�7�@vچ/���ٺZ&xة̙u�q8�lS�ţ�T"۬˜߳"ܿ?g�H,�U�:<��!_UR�^����I:�ʐ.}�����!�@A�-{�9,5'�3�%ƶ_��l�0l�P'�"�F:7����n�>J�i4�c#a3�H!�A���.�k�WR�#�?��q+�>�߂���c�'8����G��K�<�M����D�1%�#n�Aܸh��[F�����?L��/�}�k��q����s�@������ccǆH�������Et�k=�K����X�j��:p9"~��BM�i)iU"q�\{�$������@��2�Ne����\����]�bګg`�'ÚM���F�b��T��u=�)	�k����+�%��b��迪V��*���l�
��;��X�>7m��@��Oc՘�5�'�;���z�4��ʕp���;�_�D�r?w?��c4��к��ю�f5A �$���������/PG�)�������2��e��G�/R�J�=P[����_��g�?�y������|Gv`T�ű#�G�e̫�a���A:���`�HQ>�g�cS^���G��>�=���~!�Bਝ�W��3�
��������;/KE���!���|��t{8;�֍(
��o-�f�Ƌ�S�������Z�:|�8����[cR�u��9��H�0t�i<�I���5X�c����EԱ�M|[��0�=`�	�����L����]p�Dn�`�,Q�TS4���-F�nO��O�)��P��
wD���o[2�ْ��0Oｓ��D��X�P�5�dy����p�!����+��n��Gt�h�5_�
�G/��M���-f�Xhv�U"c��"�?p��s���C�I;��G���a�fy3[�<�}��E���M,Շ��[���I �����&2vE2�'�JȂ��ۿp[�Gr�,�;�+p���oH��ҿ~����'���}�-����Nv��`G��d͐�~��®��fI�� c%_������!�������p�y!=i�:��L�0N���_}Q�~�k���8Q�߈U�(��y5��ģ͒���Bj��4{��|���3�\��a�cy���U��#�{0 ��w�F�C3m�EG��?�����I��}+��N�������t�p��3R���D�~��U�dYݧ��x���׬��hya���� �)��m,���Z��͐�R<��"5s���g�c-��O��ތ 
(����r),!�g��ɀ+�S�?�4�QM���f�U�8B�X�Q����we��[p�KŻ�=��Έ�@�?�]�e&�g]ر�L����'-��4m&��Kx͸"߃�&�� �UԌ�N�`�%>(qx��:��������=�l�,̲�cp�Gm/��t��)$��W�u݉��c�U�*8#�u<T�t͸F֖���0	Ruq�]_e�C)�^�8���_Q��~��r(���*۬�T�s�L �ț�6�T��@�;Q��@�!�`6����<���PFf��l��O˦��'�fuⷌ3�AA��#������2\U�0Z���)���4e]Js�ј t���^�)��� ��f� �vp������ɺ�[�oA��;zTx�a0=�,h��a�\P��\�
��}Ap��W�L�m���ܳ|LzT���h@��TagQ�z��1��?��.(�|�{��U�b�`�*ҋ�$�����r�<�ۣ,6彥���`��ҝx���sz�nB� vk~.jX4�K�S����}J�\B"K�9�l��� #��b����7Z��U"#YV�%�4�f�*6���m2�r/s�/=����N�L�\E��i�vܧ��0Y�>��a��E��ګ��*mg��̥_)'��3����f~��<�jn��ֽQ����%����=��Њ�����q�ݘe�Ϻ>3-�!�=�4`�D�W��(���՝�-���[��
����EW~�/����o��s%�F�����	���ؗ�4��՟k*����`�S6��-F���*���7���9��"��t'l��*�[̾���Z��|���>a'PV���7HjES�� ���X�2�J��Fv�����^����e�s���ܵw�@���a}��V4�:FG�kƒ#��h8b�� �,
��}��M�V��J���_l
a�h����J��覍�������@SK��8���3��hkgx� ��#�7!�+���3L�#w"u�)O�dщ��X-�<\����O��纱���a��;���G<}зB�~d!�S]�#���E!đ�����a�2�9
L�M�CDK��"M�gwg�M
��e�*o�Q�Q��?K��W�Cg������=��:�2@h6ߺ6�!�/ʼ*_��>�w��S��E��3\�ơ�C�[�g�������W���e�V�t�!�w��R��5�zvS�!��gI�Vg�D��3�`��6�����Lm���־zL��龢1��9I:%O�DjUU N����=��Q��v�ò��r8����6q|���pH�)��=<^������@��Qi�6���6 B�y�x��$�#����X�V�EI[�9Cj�+4?�ґ�r�xK0�l?��v-� B&g��^Xq�3��W�X�Kjs�X�9��'�煴�L����Z�K�R��}3�6y���Y�����Z����-zQr5t��������\ګ�p��ը"-G�h�.Vy��q>`�k�{d�1��MW��p���f����4gmyc-�9=A��]~��C<$��=I9-g��h�[B�x�q?����%a�(O��Fkqn)��
*�^�����8�pe^�w�?_�ɾn���̅:������>�
���K��y�b�N�mr��1Q��l�`s��>���W���
l��d�O5�H{BRx���]�E+���Є���o*w!���!��%�j�q�NMX+�E�|�;��ؕ����)�=�C.D���)"�_��R~<��Q����$2��sH��v�5Ω���2�`�Ҧ��c�������s%�����������s��[Ȱ��>��6[k#>�ƅZ��^�i���&:�n/������cƎ(��`i�anܕʇd ��Q�t��B兑�a�����@�_W��.���Q��<l'fuث�of�E��Hԃo5�2+�5���ٚ]ů�̊c~����~ѝۭ.h�������T��O�z(�$hiu�iFзi���R�Nd�rK��1��R#�o������Kݫ�A�N��P{�pO@o@ ����Y�)��ܶI�,h�����3�\=q^�ku5
$V��D�\J�3ߦ�(�#�$�z�%����ZU���w��*ɠO�8��d���IY���������V��('��^���.�/�V�9Ǜts�C�����ɦ��b&�^���N"��.��X����dk%�K}�9'�BBf���d���$"p�������|I��3ڒ���3�m�����+��AD���N�w��ڐtNEm�4?ZE�8�A�cRml{�����RT����$�\@�J��[���8�TO`���W�g���@�w��'·��]�u�bK��١W�ӣ�;�=��#y�=L?�pЮ����}J����N�a�Po���a�1&����?c`�&,χ��+s-��K�7���t���[�+~~���ĺ�N�G7FP0�8�Ru�+)q��>?��jQ���Y4qs4M��bM֞s�y�{��12u�NO�~~�r��s{����Q�,�ʄt�R�����7��LN��7������/��K���֘
0�&B;ogt��X6cͥ>I� ���-k��	-�7�KR�����%1�Xo��8��ʂ��c����7Q��՚��⛪�5V��ߊ`C���2\�SVu��T|!�,i/�۳�3�!�ǷHy��>eS�kӓC8o�Rʘ�ި�\�X��ͯG[�]�פ�K�4����7�i�j(K�bPIϹ�+�#G
Ɣ^�p|�<�&Q�;��g���G�Β��U���P�{:W�r��^S�ʞI吣M��{$��C�V5ٸ��N�
����IRO8����L=�����R���:��΅ 㞀/�V� 2=&]��R|P��
�2_:d���p#`k��kMW�lu�"�^�d.!Un���Tdۢ�1�P��*�J�8�7p,]� 鏞>�u���򡮜���m���F띥��#�PX:�:Z���:�>�u�(>">1�C���n�s:i�d��o���w�m��x�b��O�Kv����`��7�D]5���6�v��;Z�2Gxc�& ��%C4��ʬ��&�ֿ=6�{�Tp �b�J���zԗh�Z��n��}Ƭ���"p��x���Z�Ӎ��5" ��<�ǔ�
�H��9Շ��M[ZK=�ń�^�cC�6ߊB��E��[���[L{��>�n �����:Vh%B�m;1Hd�F���HA{�di6v!cعEP�/��*�d,�ZXL8̽6�3�#���u�IEڜ	���:TvK�~똿ےd<�&=j�o�6Z�wܛK��F�%�-y�՗���g���~�l�-wf�ݜ�ƹf�86b�[�~���fƔ����1�s���A�������Ŀ��x���)�1W6@^����f0x�ЂϗAӸI/��G�g��`��b+߱��Km�T�#>b��g�)���f�xy��(��� f�[��T�V �=��ͯ���9σ�����dVB�!7�*2�Tf��PU��-�0�Ļ��;�_-��$��y�V���A9�;6�1�����CL�|��/���ˊ�z���!3�}����O��z�u+�!a��Z�%�e�=J �n�Ju��G�mс��Ǻ����&|���+k�BȞE�+q�f�K�X��%�~6UY���,Ly���Sg!�&d|g`_榓`�!��P.��Y��/�^�΢A;9+�P�+��
��/��ŕ:�bޜ]��1l���Y��F��ت���25��JCe=�����(�q|��ֹA�����m�G~?)���`���N!���m2�%�{ƛ�EF�������L]�� 3tnizɊ5�9�/59i��)��%�X���
�T�����w퍠�����JY�+^T}�L\��X��EB�ċ�)��Ǜ�c1�g�|W�bT�\8̲*��:�-��0��z�o�KU��X�ɵ�b�� ��B�*]#��-t�4�mh͠q�g+�MH����g�$������PQ�g��p��p��\w�"�*�C�
m��醙�T��z�I�O���n�c&���VI=]9��,��i}l� Eܠc�po8�Z�,�H}�,�� j���!����l�f��O���d����֢�@ֻ�#N��l�N��mw�H�B+����K�-�f�'��&���*�ղ�=�T�2>q�R.<�`��w�zt�� 㝮TU5�Wi��$|_��r��i�ԋ�l��u:��sM�p	�����A�z7�ߒl=�Ww'%���W(��q~��u
�I�<(���5~�*����l3W,��<2��ڟR�f������:�!�c�HhÀ槬~P �P܈#�0(6{�u}�� X����_E[�G��Lm�'@���:�Y�!�,�s�O�4P�����t�k���˾U�Gd�̌�\݂{�K(~��]���&�#jžپ6�	�����UxƷ|i��z��(�[�%Z�{�f����>�g�ޤ��:ŪQ��5gUg�xSA;2���)�y�j��r�eK��^�����*X��T Pۏ��\M�mY����8��<�3���8؇�Z�Q]�.w�]{�I=p��"��Bd��Y;��kc1x-��_i��OR��N�5Ô�<F�_#�Y��d�٥��1�T��9�|��8҃pA/�%��U�]/�!��lN%ol�1���;9�c���W��m������]NVEFP߈EL����Hx�����&%�V$4A��r�Ԝ�	 ri�2y���g��[�$1�O	�p]V�c
������T��<5#xA\���F]�yA����:hc���mA!Q38K��%R�b��9�d�Hn"*z�(��	�X`B��կ�o���3%Nx�sg���AZ��A���� �ojQ�'���0��=l�pw+ &�
K��K`M#�y-s��I+�!��[�b�Z�%��z�:7��@�}?�~��}�%���/��C(q	�'a��� 6�/�O6��^���:W��h'�����������o/!�4���/�a-�]��&���<�E���;H���z�׊�~��-�h=
(�� 
��[�p���ĩK�߻ձ�d���h�E�!͐��b� �F��r�5����C�E���/H�6���d/��AG��t�E�G��/���!�@x͒�K�$�O�V�� R;���-v��>�F<�C+����R�nI,2���FZ!ů�w��+�a��Mr��X�`�3i�$����~Iw \[]��6)S�G��
�:�n[lȔ��U�C�wR�J���Ȟ����n����e�ʲ%r�p�A�`I��	�44��CuM�2�2��p�h��vWyM��l�K���fUcdM�n�-�ä��-�\1�q�d��eq���V	�������Y�fBgط��������2?HC�Q{֯n*\�����\�/�_ڹ�;:����O��7S���Q����YΣA1K��Ռ��t]��[�j:�������2:-�;�[���i��j����k^4�5��"x2R/�y�7��,:���NR���'���js�Q9�^�PZ7�	��F$.���̺�5+�P�b;Q��A���2� ^D��X�̨�br���^�A+ �;0����(0��5�����GU�<"�D��xu����b�=��&8�q�1��<d4nnK�M�!fH�؃�hl��G=��UBm��'�G�	�?��l��QbJ8��ߺX�=D�˷ſ�uP��vn^8v���$��?��������aؑ��U�4��[]�t?P1�U�#�;:��-"B���n��M�ze}�F�kJr�&l4���G'~V�{�z��r3w��G�:�
�H�^����-&X��ɲ�)��ܞ�<Y��	����<����qA�q�O_]E���A�������js1v�N�7Nیv<N"(��$M�#�1h@?�{��5xY,X���馊x�ds�9�r����L��yV����b��qJ�^J��|'5qq��CE��t��i��(fk�q1�ܣc�U�ݤy�~o�b��T��1�<�� cF����%�*��! *6!t �����7Z��Ȁ���9�R|�/�ض\p9� 5�*K���!�`��<�Ʊ�ŒT|���:���v.���W�Π��s���r�gVز6�xw��J+����G©�Y�u0��[Q����h���%�m>Ƥ55�5�2�-[>5��ٰ'�x��~��3�$:`��;�^���]|�;�p�e$Z����bO<�\���Ā�:��J��+_�	�֞���GF)*0�p��f���M��rId^��dȮ��34	�!���˻�9[�S6�I��ǌ(o��y�a��<C�:��X$�����A�u�:<����^� 9I.m{O���]��I�
o{e�)5Ig�^`��n�$�m>)-�.c��}��nVR������ɢ< �����S�Y���}�j',6O4kV�G���`��5��@�fQ��:a���(�Sc5�{���6�Ѳb0��H&�7J��;��;�A2b�`�J�1������QlL��nGuZ�@6ja�y�����t�#���H�yۍ���~l�m�6�o��o��A>��?@�Ƭ+6�%�5������3WU�	`���ǱiЈ�Ԓ7  �����T���C�����AH�5�h�&غ6��T4�kڇ[+��>�
% V�^A�9#�BD
Q����M�6׾/"[w[5f!�����@��3 ���w����i�D˾�Ӽ�m���lC^�؂S�����\kdq!w��a�Y���ξUa��H�PE��	~S�����Q �
�S��%qqK��������<(�h!���pΫ����ڬI�R_���ҋo-N�F?C|Ԟ���~�*�مy��'��!�ӡ��ʄk�QT.Gh݅1r���H�3k��KH��3�f^�����Ví��&��*����&���ǆF�(d렡��o�bdsgsX��Ȟɐ���1ߥ�~mĕ�7��B�/���n7���e�IY��>�_2��ㇴ_{������ˊ����]�H��>����ݘ>�M��L��
�AAH�"�	��n���/(�6�����G3k*ܦZ�����>���1a9`��b;G�dG�X����9��
d�BR��0�:��ʮ�-S�;E�=�7b�}�FJ�g]DI@���v
�8�}�A���k;$P��}p=��w9?������"q�2D��
	zpi\%�$p�� �&���P�Y̐]T�ں�?%'SMX�bvD��n5��ٿ�P3����_(6S�3�j(�aMÂ� ��/d��Hq�հx���V|>37�7!��g�>6u���a�"�(x�n���v���B��]�I}�䥾b-N���M�rAj�g��A|��% ��T����!�\������	v�~e�xj�]Ng.cbEu�h)z�EtH�9�P8����Aχ�A�cae9�o��r�T~�nj�[,��Z~Z�UP�{}�G=���������d��]؉a�*���ha�LЋO[U��"$A9Ə�ME"0H��Y�J�wA��yQsv샔���. ��=v9"6L����^ 󄅄:o��Q��Un4�^6D�"+?(RP�H�2g0W�q'!�$}^`�1֟��Q�W�_����ۛ����O�_�^�D�^�����q|иd�����s�Љ���C)�3�	���*��j��9�@�Qg�1K�K0
�����\��+kB՟s'��ok�u#e���||�2u�n��n�?@���u�����`��?F������� �X�۵��1�:��J�t}sf���ҡ-)y��+98���J�P�lcUK�W��MR��z���O����Ґ )Ki��'��[��}	Ԫy-uo��`xZ4oJ��$��mĥ[Eĵlhz� �-�Ự�pʝ#�A�"�	u:�^n'Z�a���q��Դ#;}�OJI|-{�~'�󶹁����ؒ'�Pked��Qo�1�XV���gYM�1Ȼ"��b��U���Ld�p��R%���f�~z�m�GZ}���=��}�)�8'XO���o��^AПkl��G�i��
ivz9:1Q~��j۽*G�S����( �ғ�37�TRѱ�P�pq.HB=�1�O�1t��Cs���,����uD5�6<TG��/�y�nnӀo���h��J�L���u��h^w�����BV_X/������k�U+�¢�?���I}�:@������%;�7���:�QC��_*��(!
Sa`
�(!��uoj�	|�`����+�W�=O|�5J�GK��k�x�Ԁ(P�U��#�t-�����4m/cgn�װ�u�ʚn x�,e���@���� �EX�+�=�5��R��Ť�P�Vʸe����༏��a��隼M枲
� &�~�Ba�E.s�xG`V���{A�j���*���R-BJ봾^i}�nj��M,���JL�%A��R0�n�1G�d$�<~~\�9J��ؚȞ�x�m�&i�D��(��Y�e�_{+R��Ѥ�lw��O�"cm���%�m��8��2��93��=+؛r��b͂9.׮Dڨ�+��nӫ�h8���%Y%�e�`�]�`�'�
�ؤ*$:�xh�`���j���$+�$���E���'�$�Nń.�],7d�TY*Кu��Ct��6-����6�\.Y:�|HN9Q�,'�P9>\�J��9x�C��^)���b��MNP�t��5N��+�s��U��&4�S$yz␢�GM_d�Z��2�-���ݫ��Ѕ_D�G��	,T�S�ƿ��"��>�`U�wX�����<��8��D�(�1VT�6	ۯ��B{m�I�Gy�{�[��*�s��?�`�� l��6v_ �a�Zi�*C/��~;Oy��:1���x��0�̽x�.�R�'��F�G�8�B�9��Z�����[6���"	�;�$Б�6���x��g[ޖ_V��d��n������r�*��fu־���S3��(:�'�W:*EA3�TW�B��˘nb���r��J���X���J&�>J�����8L��aٟ���7��X,���C�U�i�y�4��?ˎ�3b��/����S֫��:'Y�4)�H6���z��]����E���l�^6�>�zݯC�����4]�=V�]]i���� ��<�w�R��&�	SwW���_b�~8�,hCƋ��G�_༆�~ʧ����?_�aش�͑z��˫xŻĝc�;Ne�	�+!8v�����n�{-����_�T=�����ŢsEOQ�}�������V�t �xO4�f7|���ʬ��i¬���V�����[���^P� d�=A�s!��2-����Y}&��z'z���=F�DP��d����Mh�]c&�%m!�;d`�N5��y�"u�%�؂�@M��� x��X���0�&��w~�7�1��#ں��4�r[�Z�0�2����h�E��>�>M����D��ÒϨ�yn
���pHf.i5�o��#�|�r����>�eD�
�p; {�\7K�ҴW�M�5�;�Ox2�����?��p�s�JwXhz�~�x,�QT��IN�e�[���?�4�3Yx��u��E����牣b�/}�+�8��d��O7�{�*��[8J�j�����|IG��q�
OgA�I��y��&k3���{�L\,�%t$ �ovy�^����q��TmO jÝ�#�ן�9���wn̍tK/ˡY?��2]���d����)IR��?�E�-���>������7�3ό��p[I6�:"�;��Ĺ�WfM���h~~/��G�H�K�܀+�?P���¾3�:�+0�;�y��t���ٳ
�h;�%�7���ce�~��9
ú(�����Y.�Q�4C�Gw���h��-�_@EA�u�h)�Qo#�#�g)I�n�Elc�qk�E���3�D9�>�����Xo��S��4�Ocb1�ƸU��"�
�H^��=y�v����Z�md���`�UL�DJ\�P�u�5�+��)#�W5�b�ֻEx�?�rrH�}PM����l���{����v�B�F���[�PUD���i���`5 ��5=�i�}Q��
��H '��٬G=H�+�h?��l���E;��~Ʀ{{�5A�Pe�����R�!Z���|�j�_����|]�l�:ۑl�+��=�ԛ/�v� ����T�u�Ss��3*Pc5��%w��J����yz�ip�)1`�p����U4�OT�_*iTk�O�Z����|.�����mn�H$j�]v��-�a�(E��Z����9����|Ω�օ �ً�}��[�o�u1��t��`r�ɂlբ���W�&q��Kx3h\m��5l��O��k^�S�V���ߢnĚ>{�=��A�CY������p��i�#��B�"ͺT{�V��(n�)�����/�"0�<���'V��2�r�B�3��/j�u��b��0E�M?{�P�%8��B�^=�z�	b����
1|�h�`�]� Y;�{��	�N����i���Mi���36C0u��.�+�����,@:���;$s߇�I�;`��`o�4R��YK��$�0�"��˃&�	��|��������,>��:�R�oEt��6�>Q����$���}?(��Z�F�v�HN ���OS���������c�w�gy��m��V�c6��guݑ��M������2�P9쳶MIG��F�Q/s&��g���|hv�\<�zW�<����͛rv��LR�颮P\X�����!���h�AM�MjHLP]�|�	�5&��8b��?�39]A��R��V��Ǟ~� ���}��#�7׋����`���s O{qFnO�L�%'ĚI���|�E�$����w�z�f)3��=v&I�#X����$kQë5Q8����$�Aɘ*�����\L� W��et}���VΉ)4%�D�+��F]�������������
��cѯC�7v7C��^B�ͬ21�ȃ���)aGx������J��>�H�ֵ�%����T�À]�($p]�b����i��͝�1���e�{N�r^s�s�>��v�~�i5��5���j&#��>/"�A���Kpa"�-���5$��Y�P�c�0��)��r]]bh�%T�e�����<9v5�'d?��Bc�#B�DX1�zOXG�4$���[�[�Ef\�2�� 1Jy����6��T�c]i���YTs'��31�"��1㯅�����IX���пy:��振���yg �@<I+�_g��þ�W�@5����+���F���@}��Cަ<�����\�A`�D��)���A�V�3�'�<W
m�{{&<KK����T�O��8�-~g�24��؇N�%���v���Z��I(^e�}���ڤ��W��WxǷ����e�;ȋ1���е����x�l[n��("vwY ׸b^\�[n7� L�!Ǟ�;��	aX��U�#vY��t�R	����Q��2�]I]ta�X�Ù�hr#�S9<��2�I/*H��5c}d�n���.Ӥ@f�e!�d�z�}Ϛ_EWz�%R�� n㖉v@��t���U����@7��VԢ�A��:k���4��3٪���d�>�`��u��GL4]�ȳ��fbh�i!L@���(�cr�.Û��8�fE�u�Q���Q�g�%K�:���B"�d�"Q���h���Kp%��rÌ.��D��|U9ӣ2�|6�y�rJJ�z;_����P�`�q��;SQ�;�?�8eE��58�Na�ۥ�e{�T7<�hK���nvw{�8丐㞃t2�s�F�F�;��e�z�_}� �~�q��xo�3͗��ڥ䉒e�T$D峻�z2c�»�U/��h��OX��	Ǡ����uɞ��)�?�[X)a�O7��;49����\:��Y��� �@{9L/�J(�����'��v�B� b�'��LԲz�<�P��ExO!>R�͚4}9CiVF����\��V `$õ�3��ڥ4/uվ����^ec*��]�0����b��07�#P���i@�o���j�g�a�o�֊t��[h�)H�x&D����M��%�����sU��ܑ>H�:���Ns$n��^��Г�}��%}���	i����ޤ��P鷈/>*A
���WJBӯ�H��M�E�!$5�<0���B�ڂ <�d������~f	��CƲ����0^����'�e��}Wm6��N��X� �HHX)W��}xXQhPrQ�r��e�^�ނ�C���e�`�.�<�Q���k��5�if>q�v�����-�8Z���!��u��mA�̮��a|�:/�]q�خ`�9�@���5@B�p\r�y*���Q��(����B:jR��{"flc��lzZV�!dc@O[�+�/���\�g~�	�_5����''��Tsw\�C �v��"�����[eWv��%[�2��0勝U�1@J/��1-�g�-��>xaW���@A[�$�J���e��[���� *��@����[�r���J���c��$����F�s�ڮ���k��`t�a)ʐ>�N��Q��X�B�	�,"�>��}l�LYa5p֦r\:xgq�[��W�2�Qᩱ4�Sc����1u|�q��d1���k)
*Y*goիׅ�&�[�_�����E�=�
�%u���),&o���9��9[l~�7�c,x�[����"1{*���r�M��|�������Mx���]z�'�=�/��i�}c� {�Ք雖⩝k|���f>F�lI��̍|�Cta��E�2��|��6yv����䪻�������]����շ�gQ]�Č*X�#{+Ƥ����1�����TV�(B?��i��G����s��-����	�V��"�OH?�{�#�+0�o�Lf绿+�w�Ņ=ކ�b��$�t%�1(�>�����6�~U�՘R���<n]���S�ؖ9f5F�Ѡ�i�Nb�PI^��&�e�"��e���-�`:	0��YP�WEi�Bh�̘l,*&��a{�n�z��b���IGщ�ٝ���W�{9�\Y�-қ��v����\Ƨ���M��C�enh}�����	Cv���Q������&���Zy���̀�?���S��ùm���.9���a"7`@Q�]z�=S��Z)N���c,�$��	�i����?�D�.5a�|�'Oo�� ��qב��#NVI� ���b_PS�K�~�Y{�#_�9Lb����������;���?��2�4H�eQTZ2��Z��,�Й���kq��`9����1�+�a�ִ��Fjh_��-�h�P�����^T��>�Y��V��Q���y?#�\��-ʸ���Y7y��,����x�u�`�R��&1{���ӣXuh��E�L�M�/��֒��.�����=[�Y�aJ�׵�!oy�U@=6��=Dj���xq�{����/Uռ#g�	�c*I�&�e"Q+�q�-%��,��k��!��������^տ���c�K�u�=<B�m&�`z���v܊n�N=w�޲�G7>P���`�<�X����O���~�m4���n�-~�����ҒM˨�V�m,��OZV��k0�)j�嘤g��2�"��x~8 J�X]�|�T��X^g�;�y�JLBP⥯ ��U0[�2�%@<g�^�]�+|�ίrQ��<��IQ��h�8[�0v����yuyO@�����3�+���E���!9�m�W���T�H
��׷�N 	�ܽ���8�Q
�O#�Fb�%��%v���='��k:,hcП��$}��:N����[ɵ�]��$-yE�a� �ň��E�:���"�LH�?�S�&�H�lk]�_&�c^i�\0-i��
YxI��{�t"�G0.j�ma��b`k�O��mH��i�=�Nx�#D[�o�{���(h�
4$uo��RC\)>��@E�ʲvH�<}[n�0!�kr
3l�9Vnh�ˇ�h�����w���(~Y�������d��c΢@�,�s�ȝ��x_�hA��f�����;��^i��Ԉ$��`e-i�B�R�U����͏�O%=܀�)��Rn=L��k������Q���:�b=�5�b1F7P�0��50���p��g��G�����	0�*
	�w��������W��ͣ"�V��?�#n�� �NQ�@�����Y�� "%'����5N�4�'_�#����
q��D-��wC�tr1�#5H�{D�Q;���7u�P���=»?=gC����dxk��u+�U�a5�����㇤�(k�NY�z`��D�L��tǬ3��7���$)��HT#|�gi��yZKS@�����㟷B�9S�q��%A�����wh���YG�ZϬ��s#W,�^y��a���$o����u��4{c���e.�=���(	�+�9#�f|TsI�X�G�R$=�9c��'�VG@Ab_ʈE��k��&�(�i������a��%`�a����k�5L���i�h�H��+)��(n8ӾPcLr�7�\YRm�[��L�d`U��u�CS�=�ƿoQ�JH�?��ԙdpu�l�\;�| V��J��1��6U�>��|�D�I2��f%��*��"MF��[0�u�n�i!u���r��=�RM� ƞ��d��sH1��� �Hea	����/�<���dg6������}NQ���q��OrWF��s�ZFkD\!ʻ��y��P˻��D#첆�p����?�4xo�{n]���Əx��0m��G��K4���Z�7b=�Mg�ט��7qX��GCrj�ʱ`���N	���Z��b�����'Dg�Z6ȥ�v�R�!�O�ӆ��_s2CeH��h]H��t��#ڣ͝51DA�h��&������A��OG=���'W�' F��Ӏ �<"�+���+��ɋ3�0���FLw�����>;w�㦒�#ʯid�Ϧ�,ʤI@[�,�c���Bb;�Y\S��`U��>iv��1������_��M:;5w/��3�~;�-&�U������"���Y+�2P�e�g�$�Ĳ4��]S����Y�5	��at1�Ao���Q`�����	����C~(	�v�8,wӌm:�����ś$}�P!L�k)�9��}=U�V��ul���;@��?i��3�5b�h�h��Hw�X	n1�'t1�rGI�+�wC��.;0��� W^h�`
$�[1�?�3�ova�=�m6"���Ѫ)Ŕ�������ۻ��ވAl�fh�v��gk"
~LV�5r�Rd�L	%��)�s���`��חS��ZH	�c�lLv?㹩>;��]��Kz�Edbz�|��J�<>F�9�n=UP�Y�E4�/���`m�n���Ly�1u���.{Hu����P���s�D�b��c&�s4*	��`����b��;� �SĔR0G���-���z3s� ���&i��eo���b����:c����lV��1Գ��-�D_�����U�c�����*��(�.@���a�Jq����ͺO
 �2[��D]�A�@:�D�� 
Ǉ% �}�P~���9�d\Bϲ�<Ydʧvj�{�|VX�gj>s���9��Q�V�F~@�k��5��������l�"ٜ]�������o�;|�֤�V<��ٵ�fK��nX��k��9b7��	ǫS�3�We�c?+�]y>}b,�\'e���5�-��X��L����I�?�G�Duz�7��ŎʿP��j�Y�$_<1
��{Iǖ��_�̶�p��V64��ؿ��f��G+\�V(����VBS"Q��XS��6�������o�CR}?�W,6�\�����o�۳{>嘜m�G'��k�N�c�-I7^"X3ˁiS�h[J3�wnDő�':a$9�-�Ԍ��<�dLe���k�N���/�2���2Q��Ĭb,}*3P,��ό�|*&�������e��O��X��̙��o<��\�V��Q�j@�_r~��ۯ���
�A91��0E�q�0H~q$����{��O���&�;w��j����V��%�c"h��K��^qT)B���������x����Ҁ�TYL��/+�ק�� ف�@��y��6��H�w	��y��ۣ�Y��`�,���<�4��j�w�'̌8�yϱ+b��:�:ϬR�^���Q�o�^3_��	�0��dKm���ꨊ빍@�
8��ideʞJ+��Y�eI�]B��B�NR.�Չ����r*���ax(G�����,�N�϶�%Y�_rp_z�;�����#�;!s�c�\1o���4 �����������吭|�M�r��K��1�VRB��
�gg�	�ʓT(/����o�3lB������k����	lL�U~JǶ��""é=`�H�0�;�PS���R3�� ƪ$�񪵭�'l~����e��+��gnl�Б}V�46_\<��q�.�z���Q[�V� +n?�5����_�HB��ݶF��Ð���{�|�:!װ@��$�]�{@���b�A��3ҙ7d5/��ڭU_���-�����L �b�5�D2B3�6�nY90d���1S2;,,Hd��
7mz�E�#Ue��{�	^��x0B�^03�Y��W�M��� �'�t6�
J{�;�2u�$g*��d#BT0s���λL��,	��C��xT�"c�2;�[�f~X��pҙ�&A�}N�zT�k��.v	%��9��'�>SU�"=�}��*0��c��7JBǨਠ솪���
��f�*m��q���R���H*a,z<�|�2]��T�^�UUQ���!ʸ��mVt��b��`� ��������n7٘i��/ch���r��M�;8ʼ(^�&�E1{�=�,�wڣQ�mor/ [�>|VMuu�4D�����?�o��/p_恣��G��RK_�%��u�L�*�}' �E��~��3[Y�p��ee=����ƭB���x���~~f6�D��ڜ%siW3�]�w+8n�q��4��M
��9��6�N#�C���5�#���I�>1����Pk�R�6y\�ر'�j�i��E?������`/�-�f������G{�4��J�p�/b�3�*�,E����=����p+��q�7%�Nm�q�Tp��~���&i)�����s� G�J5&kY�)����oφ�s�1�wZ쿅�z� �3(� ��7
t��]��񕍞R]&}�PI.�*2�ьc���ˊ�&�ǅ�ԱG>	��r?VV�$�<��5�_�:@3�&�6y��౎��]�ןV[_Bma��͛A��_�S�D�Lb��+�=���7�4�N� �[Gܿ�����v�lx��WT�aq=Uv���\F1"#��c^/�z����
��'����CIC�.���ȓ�f;���,@$oex�]��Ty�������l/2�h���i:�3�j����=!�wL��}
�Ͼ��E�1�v�y��[#�2�rČi�f��z�ۅ����L�U�[��?Kg(%,��������eC�����w����Uq���V�vO#pӉ8�J�ה|Y%;��"K�|]��y~��������P�Ǒ�}Du�Z���9-�R_�Zq�����d��H�ᖝJh�oy>�����3����3��g+�>Yd`�/�O*5r�	��t� 1SF�u[�G�x�} �g �4i�z+���i{�#$E&��%bs6�U��M�Y���4��D�Ӡ�n��c}�鶄��6Sv M��H���_Q������GG�K���*f�h���V�Ņ�f�^��-�:]�l�Ř�w= -b����a$źp��f�\��X��^)���5����ۊ�Ӗ<Ec�a�xR 7�Z-/����a�Z���n��)����(��v�����:�k��2Q�|�V����CC�Qհ�OR�Ss�NZ|�e��;��gO�IV.��qSw����j�a��S������O�k�X��0O(z�Ê)��;�yqV��'8�����.��mP"�O��Q� zL{8�Y.�<���Y}f�Fv�[�&;ſ�<��	�(h~��2�=�x����!t\^lp��%�t[E���h���@1x�,�X�fq�~f#�����&�0�����+\�nķO߯ljʲ�J@f:	eR�28��e�������XV'���+{ʿ�i�byy����N"}�(��ɪ�l	y������}|�d����C�}���0�_d�X+�O���4CH���� ^36G	��3:�?Oƅ�Ph#����8D��B��=�A��Jҳ��Z��y�D�E��pݟ��� 	���v�@H�Q�W���=Saw�!&���y�������!>��ɜV����w��>���攣�y= �c���#6}��G�Bm���=^�ӭ{�d����U�?�� ���'�S��k��S��5��c���%��Z|���gڹ���W֭u�'�3������D r�$���6�t�C�X8SG�TK+E�PV(�-"�@���2��~5>i�R~-DAj�M]J��v�r���(�%���;j�?�
����%=��~[���d�:N��]j�[�2�Sx�J�@���l�lnym�a�N	�8���~�C��U�|3����M-eR�D�#4:�,�Q�<���[�.U�Ѿ��/�d�'C��"6{�3ګ����O1}��7���?�Y�]$gVV�u��pӷ�N�c2����e���4��p
�C15����鞗t���/��F��:��Jd�txB��U��> c�>�B��
�Ӕ��/�&9�$��a?�oY�ģ�&3aݻ
(�hK&�B2�!�[�	~�����[���ZN)�]�EW;?��-�z]���V��$����4���OUѫ�d��W�[�9�c��ՍȁOh��$��r{t���XZ������R�~�3�U��PwLK�%��w�*I�
��8�v�c!l�ߪ�`�]�CO�:`(�&:��_;�S��k�x;�n�:�R?u��:
��Q@ �
<��8R��̡Bj����cA'�-���؋o#N���g��a�ɀ� ��z����JY�.C�-<M��
_G�H�N�O�b$þ�$+�bv�ŕ�Z�^c�YE���p��t�ͳ�-���g��&�ƀCu_��\�+c��!��V10"}М�qie��4��h�[�b�l��YLhVPɼc;m|�O���m~iC	�8�,哓˒������]����eP4���#a� �o��]��7k� �� Oa�~pczϒSJVŮ�i��%ڜ�@����|З�+�Z?<��uI��Vg�(�S0��a�(C(�� 1��a%7) G��q�'ڴȉM�#~� �aD�a�jr=��tܕ����xT�C��ƃ�t�͸�p�
�h��5�qa�E	�L��$�:�X]WPK̝�?v��r����ͻ��dU/�}Ћ�}w�X�۠��2;%%�'TI� ~Ir>C��,:"y����N:e��v�:E�F��@D�Ś�Z�v�Bc��WE�T�8������p�G����Or�^���f���_I�ad>}���j�<�H*����Z��&D�\"9�v{M3�)���^F�ą�-td�>�X�Mᱯ@/1ɓ]��>�r*۱�}Aoٟ)"��[~t�yT��`���'l��0I��t�!�8�a9�.���3q���]�GD�U�����VG|$]z����d�#M��48�o:�ix��zbt�}�E8�P�h����m'�%�Rޝ�'�l��A���J<h�b�A�IjAw�`&a'�Lh[�n��n<\ִ!���\�Q��?~Np�!L@�V�\g1��I]\���V�P�h6����_-�J&��å�.��&c�b����i����uȧŸ���ù��t����M-�8�q#l�v>�]�{�/�_1pmjN}��"ڦ��
;�{[�ߠ�{�u�jLQ��i���gg��@�dɊ��9�l���?����^'pU=}VX�j�2>�]!x⣖�0�R�:p1\s�z�(�?v���VZ�o�S�nBm��������45��"ck�@h	��DU�cB�b��B�L�2��9�z��<�^�|�n��Z�_����ڂ�Xٻ\��	(�B[L�[��^�x�_���0!���� U���!׷D�01�qiϛ|Hou�fD2�מ��$�^�B�t���`P�z�|1�Zuu�aT ��k��0K?�&x>MS�4A<��]�.�K����.>h΢.(�����2�����.2��x�<�Wɀ��cg��N���7$����5�f�"<�rv��+{��z����f놼	T��(�o�b@`rq�p�1�n/�jsv�i�%�s�<짳m�U�i{�ݯ�JMֻ���8b?T��`�@�f;��1�+r$=�3R���ݐ��Os��cP3��G'�ɭw�����oِ���.�e<˴�f�@;G�\Q�vf�{�D�`%�x��a kS|Ƴh�W�;x�V���M`��c"�~����k�� �.J>�T!�h��< CH��+��Զw�H`X��9�)<1FK
$uB�����#��\%=�-5�"+�K��ЬT��Ȣ�H�6����MŃ��������Ng� r�̿է���s�S`	�CIQ�RQ'�դ5��?��m�j4)��X/���1LV�Ҕ��(,~Щl++���[�4���V{��3O���C�S�2._��-V�jC�/���y���?kL����*bߩ�t��!���8w��.��)���W=U�oq��?�;�l��(O�b�_�:}�C�:�`sT��a!���p���+i�e�}�1b� aG�DB�^P��P
���/���*}�__��1�Je��s`L��r��C=����TL�A���[�£�!���@��=<xۉG��M廿%αN�EA���Ve���s��4�M9�ߋw�
�Oa9���	5&-��(d:���3�#�f&� ���W����g�X�xV�-����gQ9�׌.gF�$W��4�*ӏ(��#�����{~։��h1�#Th�.5o<hnO��i�J|��~�	Gs1z�������9_5�p'v��*�.� z�fL�!�zQ5�3	S9�з��3-I�� ��Ds�'����X��w��!fR�*�K�4ѣŜ@�b[)��'0M2�*4I�v_ng�%	������:�T��D���y�ҕ|�ӛK����s�^���BB����e0Ar6�EHZ{�p���aq��.�s���<�C$�vw.Y�#ޭn��dv����֌��b�����AT���P�qМ������^{�O��d��	��m���B�V�F.)^�]�gP�pLt��5�
I���L� ��$K#_����|�����8���&�r4Ì53U �m@��@މ��/{�Da�Yخ�+����`�N+�ܥ��T����p�(�.��󠺕ȱֻ�hg�+ؾ�� K"��'�!��yJ��I�i��
�I���	��m�фQl-xG�N�"�KD����	���;�Y��zE|fm��,A����ո���i�]S���v�f����{?U&�'[��\'�m��/�����ZĹC�f�͍X�$G�9������*����hⰠ;6�_�Gw����t���i�*_�����02�!�(D��A�v�|c��$�󵤦��H ���a��Tٵ��������H��a`+F_�c������e^D���Mns]��������AC]^�b����b¨^J∢R�T�>p���6l����Bf_;E�����[��1<u��BA�x��Rq��a��l*������׆���"��W���[H��1�%IΑz��"�J�:}B���T��9��uLk盀\J{��8�+�����X~)�%�/���V4n�SU�<���y︭Δט�A��CC�-�/�o��!
@H�Y#�� ��ͩ}�#)��F�D1�nt��*���	����
v�'p�s��Ίݬ
Y�?���Ww�V����穚`i�����8mmzd�NJ}��ȩ����W�FDqԗ��g��'�F�['%�	6R�a����zq�����.� ݊ۼ��OS����o��-pՒ���J\D(�K-d�K��%'g��[9���&�8�P̮��U�ɧ�G�|Svo;�a�h�	R7�?3���S^�I"8s�BBa�e;�M8HU�L�!��f��@Z���z�VN���'�a؅�%�kK}��H�ЀW��;��r;n��-5X�K�d6Ce�lZ�|R�`Ì���@z�4I�ˬl��$FC�:'����*w�$í�ͤCd6�	�rc������6 GX��u��-E =��kY�}��UY\�:ŸT�>r,���$ȿV1oaTN,��WT�U��t�.\��������;���b�Kk�/�`����%'�� wķ�$}�3_�>i�7t������y��5��Ӭf��Qq����3�`��h����aL������2K]��}�u!��0�m�Ƙ@D�y=H�3A@f��8�*AIZI���;u���:,ud�2�̐ҝ#�ED���W:l�x�K�LR2m�x+G�o?�6���
7��0����XwJ��g�"�im,R7����B�5�jg�(����Qܾ:��m��;L��E&^�Uthd�R���"�%e��������^�\7��	���J	�(��*튥�Ձe�$�B	N�u��X��˕=]�RA�I2���Q�%��_�"i)?���>8�&<�^B��$&��ڃ��؎�w���cW��4�%սo2�$MI���mqE�W��)�1��&����%�*�|�n���٬e�;�����o7>�	U7Q-��w���nq
҃��p���`��@�5�m���H����W÷��e�bC��@1Ԟ8�ވ�������M��F��[d��̍j�Q�<�+�l=�L��� ��w&��p��l(� .e��j��@72�5�qF���k{��+��:�^�F�~끑�6���Wkx���x@!����t�)3�6�h�N-aǡ8}o�C�,�����Y�h��zX,M��y?�<%��	���A�r)�
���v��;Fs�����ޚ�V~Akh�E$�B �
74-���amCʱ�?�Cjn�J���C���@�Q(�7��/���/6F��Ʉ=m�ڂI�_`k���\�����2�/u�{�R����ôPLu
�!�Q�f�6�h����nE�j��ʃ��=qE�̼�G��vX?Hl �P��y�j��v���Ȇ�yQ+��B��q���X���$��`��:� �P����S|1�wot����_Du4F��֖\r�T(Fp��*Ըk<��~UN�H��ƏE=�63�5�!bt����d*wޡo�Ӹ���-�p�{����A�M��� � !xB�׎`����Z��~.�?p8۳�Q���%^ϭ*��#QIuHW��E-�Z��(2@m2T|ˮ�>%�U�:4~[�G�p� ;T&h�@������U�
�'Zq_@�K
=U/n�^�\��uIE;�j��>�^C���*,Y;�$A�5�G�s|dPm�u�.�@fP����md���������J[^����F-<����� yW/��듁������'#.g�s*��f_� �L�2�^4�öא%�
(͙ڃ���9��)��O����X�K}�~�S;/�HZ7;�SA� B��E����1޳��|�;Iί��F x��CD.��Ӝ�b�r������&ș=&2M�=PC����al����
�y諮�Bރ�u�[U��R��zR�ܼ E8&�f��&J4���A]Q�gz;3RA8��h�����E[G��Xx`��g��Q��^�9����+e�n�C���QM�	�Є��D�7S8P�M�M}_5H�[� �8YP����&�U�y����Sϒ������{�Al\�%.	t
�c�|i��:���(��&lS�.�����B̠��R ��Z4� ��;��ػ�������b�az���7��(&p02���;�|Q�?��=�E�hՌ�0o;Ҹ�>��ZTҏ��\����	���Z�0&H��uE�߭����I�:j��wvF�8"'�ʎ��d���m�l����v��(r�B���~�_�c��L��:�ܻK��J�>u�O#���A:x�m��A,�!��������t��Q�胵�ԭ�h��;���]PP\J�1�S	���&�A�@���:�߁����sMH��AV2r��E&��F�)4>����Ȑ�w�C�X��������
^�Ja,_`�zq孳�Lsu�f��}tpE@����w�w�$^�5+�H�B�T˷�!�����!�)�U�&d;ɀ�Qu�LA\�-���{utQ i��?Y�;@��
J�R�^�e �w��K}�������M�{x�b>�`O������ᅼ�H���*��g��UӯOU�kp��a��xY��C`���P�6�/˼qj�j�޴�a��o�SҾi�t�Q����8��ee)B���>L]��;'M����$��y��@��Nz����1Kp�.Lս�7��r�%���ŗ4Ԩw-�X��Ӷt���?���x�*�}��u�ؚf��#)����A�\����N;�j�B%�
�nn�L�Y0eX���ZE�M�u��<+T�:�ה�Ѳ��o��DvV�-T�485�岠��gm�D���5/l�q�g��$\�G���VW8H5��O��>��G% �W�Ռ�E>�%y�=�33����l���j���!�ũq�,TQo;]T|��6����zz�F�cz�S#�����by�a����剮�Bx�i��;r �@�̃�\�,�FrQ
��]Su�R|��Kjo����ۻ�;�r�켕0v�Gq�s�����)� �&F�p�2��KQ:���32�����3����`3z�z~��Y��+�CO���v�J!V
�I|��0�ׁ����x���"�GE���D����B�?E�`ڙ�.��Vk�0zq���`���w��[����fV�4D�u�Gi;��s�[)����J5�Fќ˞��d���W�t���J:��h��?���	��
�Dλ�w�ri��O�Z�T�u�yc�.����	!���^�d�:0�� �����5)���6b��m�'�5����6)�q?.�f��\�4���lA�':�ke�k�)��RYF)>�p�Y��,���ԣUG(9�t��pV�i�ݿ-%!��Hr�?��s�xi�t���A��	�+".���)�*����V6��I��әħ������	p�E ۮ���^|8W|����/ZHU�6��Ѥ��fO;�+y�l�dvIiƯc��
3	�v :�^��5
��fnᲛfns��T!D�j ��3Jǜ�$�M�
J:���sk��i&��(9�{&a��kg�?�=�"˭������Z>1 |j�g+~�C��ED;v(��j"D��^��V�}�Ђ�ǌ�
>��aP��5��/���/!����㞋mE�u�?O)�M�|���u�)��3�K���:��
O�L�+u�$���/�΅%@��Ä�X_����}��Ya@����9j�tQ7S�/i�",nH<�)���d=��ߘ���A�@��)ͰN�ð&�w����-/�bM�^sm���㷐d8w-΃�4��,$16���T/+6H誘�V�r���9 �H#!�׉o��#'ݞ�%'�D��pG�#	m��B4�)��9��
�4�`U!���Hg���fj�_VYR��M���Ch�!~'#5�/#�.Sg^��뷀����^���iƩ@�:���Y�GΖ��w#�y���D1l����?z�t6Vt!a�86H˪�^�{�.�� M��X�	7HR��lq��lC��2�Un���	��y�]P<���#�	��o�Cܯoޕ��,�8���5"�<�&��>�������0)�g;���7�g�a)�l��8�>E�Ш<�a��3ު��WY`Ah�}��o�E��A��|�� ��\1jD��Ӆ�T�}�t?-���c�r���o������[���CQ����46���a&Gʊ��K&��b����}p5 �<��C�Y���M&��ż��-!uw���)g>J��������N�X7A�^��g@����ֶ4E����癃廪#.��#y�(ʑ[wX�U� �A�q)zV<�9jR`��j�r+��?�o�f����
��f�H�+[�R���bS/��T3�\aZ���?��r,"J���e��	rGu&5���(�9����ua���lC+����B:	46 Slں=���7 �5����i�.���'�]��!��ڧ�}wk�n5��)c722��n�\�z��A�hf�9M[�Wjp���'Bpl\��ȅ�റU�FJ���v���0*�$�A��@~6�o�sj����α�(}���4��'!
�V:p�/���q֧j��_���-Z������A�\�=H�-�M��v�3�6��M�k�Sq�'Y��t����=��6�R@����p'fa�U~��
_�ߦ'U���	�Z��"�ո,9����>EI����������a'y2�JGJW�ɦU�/���b�+b� G(�f8aP�94�|�h���O ��4��"a�8B�.��׆J�����XQ&��L���Կ0Qs䕝��.�@5��7�Y*��/~��_A�� ��8D4{}��ס��x�R�-���f�@ړ}�DX+�4�j�kO[&6ȿO*�O���&m�A	�5N���ճ��ؑ�������@��u�Wz#��sh�?f��nЩ�܉����DE<��`+�K�>�d ��D��ҧ���Qh���%+�]�B僐���N�$p��0��~�%�J�:��D~ˁ�z�|�H�1,lA��q�un���}��(җ~L�=aE�e�UHdooO5~��Lk�����
�7�����j����\Q7w�I�aN��d�l��O8��5@g��}��� �#Z�F�JPN�|�V�r�y3/Ǆ���ނ��d�@��Ç�(�gW�E��F����$d�o1<#�������LT�\\�
�s�7�$�(	��h4�JjF#��"�w�����^T�"�����$i����Z!�r7^	b{�<QP�,ag]�/�\Eʙ�n�j��soR��y���e��<�z��#�?r�R���� {�%<e=�������p�riP>vY=_̏��y{�����n�.E8�,n�����R���8�����ex�_r>R��[B�E����ˏ��2�X���)�������0�LX���LE��,x!ű��qx��3vZa��b������ B8���P�b.^Jy�� n�B��q����?���]x�b�D����x�ӫ��b� �J,�5ٝ�/j��M�<�Y�tǶ3���+���g�JG��;��ţ�k�0�qn#�g>5���I
��%�W�4c�������z��}HgeG�+��bŋqpcKkE+������Y�fvU��@����Jw]Qm:ܸF�(L�2ּF���Y"�w7�'=O��U�0�L$U�[!7f#U�����S�@�N�����?���_V�
��9�B�AB�Y�9��|��V�l��mYYp�m�͙���v'��)��9����p6����B�_5�-(ܼ^˙��>�,�� 9�r�h�.5��ݞ�iu@֤ݛ���w�|�yQ�s8����{���Tӈˉ�N^ ת�Y�WtǸ�d��ғ@�R���e�o1P"�\E����xΆ�L���?J)�!-��$�������o>���ɳ��R����UP�lT�G�4��3��[?{��+�S$V�G��EzOJw��n(\�Ә�ֱ��f`=+��i��m��<��b�u�F��}VN��h{������c�A�� ������ �ūy�Q�����
��9�>��'DM&�r	Z|UMh�y3Վ�C�������7�f��n'��� �c�%�ޒ5fuvwT�ߺH�@h4�X_�R��5`����>���&�re�A�z� ��W�Ѓ���������GX�,��m��s?�$�K�ug�����������G��V^�:7j_�Ƅ?7}��m��%�B���\Ҧ֕9��V�+ڔ�N`
]�Ke�$J�_�Ǝi�=��偑�v�_�,��G�V�(�߽~=�����*�p�Q ��C�� c&��h3MҎ�EC)4I���8ё��,]S;ҍ���u�w���ͬ|Wv����?�Y�]�"��	���6أ�2��@��l\��5��Qs�m��#�;50�E��:j�)��������?TSy�d3o�p{ė�N.S�kP�80�ǅ�=�-up5q/­��}n�"�m$;���l�K�9��ȗ��W�tXs����|h\1�p�\ǐ�x(�0U�l����FfU�)�;[:��Q�y?5T�ǵw�b��Xe��K���G�*a�� Zm8+g$-O�����)q��ٍz{���g���m&,uҎ�Ç��{6F\
x�A�άG=u9�2�K�/��8��?��D���؛�EN4��)�ý��m׹=���O���B����k't�{SR[�0j�K�aQ�cU����U�+�ۤ�z�{��r����c2���c�' ܳPN�(�@���D��]�t�N��J� q�N�m!?��~X��ƷE�K����/�q��c-9V*�:��7v����{]�#�"C�|�W�:��h\�	�jK���Q�Fs@�{��rV;7�ΦP�I�'��k෍�e�&������gj�+�2�+�~)AT���N3�/��4_X�*mVݖ��2�����m!�*;�!����������fB�<�Ǒ[R��'=��T/�4U�ɚ�_�y��7���
�j�%=�Aö�0�L��{Z��zoK�R)��9�GK��5��mS��q�c���txz��\9����U
=_�jAt�ͫ\�=�|� ���ED��������ãF�θ������$7�m�x��e٘�֘T��c���b��~�#�	?����3�ö�C]�5�&��0v�2��k�����[�=�j�w�ˍf��~��S�O�;��7I�!nc���C)����������h�}s���`�xA���W��L�E����✃�@E�@�@,I�=F9,�?|�ֻ��@�Km0,(
U�2q��	P(W�R��q�f�M��=��fu�p��<��z��ByK�8��H�aª��c�$�A�\�Zr&oQlN{����5]G;�ۺ=$�C#���"���x�vV�%�i� ��E��fψ�R'��i5r4?��[*~�O#���*"�5��q�P���fg��X<�Pm��V�>���Mz�EFB�~߂&zYM��( ��Y�ǮnX��&������UXa�mO�{T��~��̦�<r��K>�*�</}�Tr����|�B6�߿LH��g%�D95e4 �'��͠��Z�d�tzs�Z�D?�A������:bW�����DF:qjb1��DpF����^�9��Ɯ%A�C���P��|]b�\����p��vL����q���9 �0��l[��8#xg�$ɎOzpj�6�u<m�(i�ש[x�.�,���]�m��C}�!�_��lacnS�e7�XY��.��A�DoS0%��vڳT?����m�N���sS@o>�|��mH��q�gU�םTR�%%d����6�)�{�:��Xmv�ǚK�9�F1�B��������f~��{��r_�:,�/s�v���)E�]� _���C��Yߔ����s���1��N�B���3��{��rc`�D�P慡��v���Z��@�v�C����pv���C%�ѰE5��>3��y(tt���'s֒+�,��%6���^�K����h{�~θ�}.��#T.���W�)b�UAy�y��Yc��h��1y��U-\��3���1�C��^��X)�ű��#B�*�R32�:ğ�_������V����S2���j�y�H�D9��{a���
3n���CbՊ��~��_��9Ugy����ڀ�q)U�w�W)��))�;s�w�U[{��o�VC�~��n���O]��xuȍ�#kv��^���Ԝ�_c泼��������XX�L��Y-�%Yzl�_��Ҳ9�b���?�h�(��+�	��v������ �b6jq�C�)�Sc��=b�S'xQ�MӾ�k��,|����}��P���g�q��b��s"�M|���*�a:R$�b9S%���}M�%#:�`Ϝ����@5\9�T']'�]�S1\̰Q�p5�~W�:5Y2�����9�f*ՒJ�u.�N�\�
�C��T�J�l9_�|釼n��k�X���Z�"���<I�/�j3ݳ�*�$��[q���X��e!����oE�o
�G�'���)�T}�kYE$H4ؠ�<��ٔ\<=D��)1��r�s��6���wZ��AY
�W]��fT�F�,�Z�������K�ʦ�����O��а��Ԝ��*�zu�����>!�CB��?���1���O���6�V��%+%���8P̶֓SѲ[����S�7i wD-1�4�"E���9�bcw����K%-�0(����dW��6��-�+[@�����sJD��-$ȵ�i�KY��nBa�l,��������H륙K�����$Q9�<h��jyj�vޮ�`���&!�}�p�7#��p���L��PJ�a���|��d0�K�O����=��c@J����Z#�W�	+>���3 �X��s�+��"�
�uv��H�5S��>��.c���i���\ae�dnr����Ѿ�I�M]�|)�U��*��I��*N�#H�$��L�3�,�k���|y�z��g28��<�fw�M��h1ŦP~������7[�+��X�g���f���p蛜.Ϫ��gw�mC���.2m;H�
����H�9��$C\�DEY�Cyv!-�{%��XS>U�Li��,��R?1SE�����d��.�1����??y�v-��k�G�vqt��&�x�.�X�8ȑ%tJӨ2r�-���Zyt�8޹�ީOǂ�õ��L���d�g�{�����O����Ӹ��zU{fBD=��R2^	*i7�30� �V���m��0���7�kVjG��}�dX��ؗF�H �[pr�UKZ��?���#M��{��dm��#Zp��B>\��.�����b0d��T���7���N��V�e�{\ɚ�Dm�jQTO��H�׏8*5H}z�P��C��#��ʫacE6���(��3 ���	X7�
�j��N�j��,�Yc���#46N���dG�.��:������pV.�J�zk���Q.<�h�䆺Gn%p��r5�nM���[����_�t%d�d�q/��Z��l��6��u��z���}��+�da�<�,����~��a}vI��F����q��LE�7�[�I��XiJp���h":#���m�hn���L���?���2z\�v�2�{���)p�f/���f$_U=Db(.Pn��{�*�|K~?&L}�̐>��T��ȏ��>���8X<���5(�r��Q!*�:v2|��S;w3�Na��OȒ��:G/܌G��\?�	�ϑ�>Vw��$�X�c�CEn؏K��z�L���}0�tw��<e�s~}�F�ɬ=I���l�� �(]1�%��vE4169:}0�S ���H�#�k	q��?��	�eZ܃wF,������R���Z�����/rw�{Q�!�{���78�{����GGgz���?OW`����<�Uz-ߋBN�,�Ȍ�l��Qňpda"%����S��C��p#���.�ބ|l�ڥS���M"�8�o�=��S�R,�! �����Mf�_�q�2f�e��� �z�ZP�ͤd�� !W#��^*� e�с�GC&�h�A��	jR�/�p@-����;*�q�C��|�X��*��N6�䴅�Wwhv�LIk>��
������{����;�x�8.�vV,�%^|`Z�y�@�~����pFª�L���p'�$=�z��*1�&�?lOo+�*EU�J�úAަh�����TzK+���5��T�ַc�#�
����s5c�W�[,or�?J�jS��눔=�pgM�ˮG���N�NN
+&�P��@���vR���؛�ز�u�GG\��ǱB�]���i��.�%"뭔��0C����z���g�T�r��y���>W��cPK�!^'$ܟ���-��4����y�z���ꗘdd���gM�{��`�.�r��7�c5�cF��#(�h��:�Њ����GC��sv0�+V��������F�l`*&��E`C��
2='��l�w�����M96�g3� �5����|�1Z��0�UR�Wm , i ������#�Q�d�Ţ>2�b@!?28�:�A_jC���9g�.s�����a�k�$��g��ﰮ cY�b,��[��&1&�5��W2w�K&�դ���):����S�u�G'bm���=�UBW�~g���mO��5���Հ�wD��ٳz����f2�g���dQ��ysV���j;��9���
��.��;���.��Mu�W�8��z�?+a.����I;��R�f�s�)�[�LN[�J⃍M5v�-k�t���}t1ZYlim���2D�R�ػ�F��DW�ۇ�{h�0���@��H-��T,!�*Ӱ���� �t�YS�k�x!h&4����id�^j�7��2��dZ(��-����ˊ����8[T�ӎU��p?~�ad??���ʐܟ��M�/��l��_}.�f.#��0�t�]ǀ@>,y���%����2��l���J�����*_��{�5��x�������S����ˇ�����BjQ-�r��'���Epɨ�7Ie��d�3ش��doc,��[����QoH���މw��S�`�����ؐǤ�-�v����K�%~|�|W�xV*U0Z�(�������R��7e|#��W��W��<+b�a���'Xq��q!������x�SkaNnw}n:X#zS�X������H�L)��_���_��-��$�?����5v�b)	)���V;���[������}�����a�ΰc���VEϙ�S������~a�(�i�����_�>V$|��V�Y>c<�f�I���@����Z���w�/�[3�[d;�m�|刓z[|$C�Τm��BBӧ�nzex��_�}�}p�6�/��)��
��s��I=��W���3
�tm>�̜�i��S�
��D�pZj��⪯>�0�%��4rt%C�JX�D��b��n�x`���]�Cw3C3���gX������(ў�.)�s�a=^3 ������J_ª��9�8�j�Tp�i���"�,;~�7"���v#����h�`W���(?TJ�&8��Sq�������x��&���$`�0� ��`:�&��j�t��*	��Tt �Z��K{S��;@[,������l���)��+g N@��6>�r*�'Ob"j�'�[��i�O�Fu�X�҄��,����:���+~1a��nw�$}�ї �n�*�v��ͷ��e�#��>7��\���B�M���i����wǼ�CsB?]��l\�IC�tB���BX��9��+���|aT���8}�f�v(��1�7�6��m���UoF�!��$n�Wy��)u;��Y��^#aH�ᐰXe�t�� M�q��2w_����V�Ș�\�[�/�0�BW�m�!���@����[�U��<&�b�r?n5-;��tj���s�dZ7(���$�&?%�tEx�otD�7I�A��RڮqH��(\��ⅲh�\��S�ެ���`���]w��7� OL�ڪ�,��.�T�8`W{kN�<���I�"���3݉)��]��!�����#�_���V�R;PJ����K��J0e�n�腾r╹W� I���J�7S���'�Z�3m��QfAh8�a���_�eX7l�	��1B���c��T�d���Y�yx�50X�``2/��n\��앵϶y��@��E{ʷ9P�o�����ϣ֭XVp�A��s�n{h�C��-�(c#��)x�
س�0�x9 ߊ�1s�5�h6[��R�,\A�Ţ��ҙ�=���UewJ�gvŗ�.E� e,.e�׾-�qrp�a����w���A�ש�2�C?��`�����,I}�� ǹOӨFl��`������A���_B�V���L�o���	A���vΜ�J����q���ps�aE��%���Q���(MW���?㴼p�2����(�	�O�"�'{!z�B6W�^�N�n�W�����xmCH�m�)��/�q@W7 EБ�:����W�����ٰ���3�Rc �;���'1�y��M2�f�lh��!<fHݓO�K�-ᆝ���Θ��Bh,��J�tAK˗�ZsE�u�i�L��T�Z�l�Q	�g��a��L�Qh �&�0F�l`�F�_�ͧ�P瑮����'	Z��p��~��@%տ$��oj�K��9A��fî���4T^g��0��a������J���{l���O��D#�����洝&�H:�J�!n������r��<{Hx&���I��b ޕ�%�i_x��#(�~vB>��ܗ� -B���_[�cRY�/;vD�6��ri2�/�?m��j8�,K��
����|��8�%a?q0a�>�a�����Έ��,����Jb�êO��VDoR����^�G�F)�B�W1k��ػ�<�H�=�5��Bʲ9��S�/�[�(�����s
�@L�]���N?�p���ّS�B�߆Rje����DZ8n1p3�+�7�JL���xg��]�~ͪ�^-r#�'8��+�발,U��VK�s)�(�����DJ6���d��6c�8�j�%�O��W����Z.s�����3Ѵf�w^0o�YM3��4&U�nr^ϸs� ���u壔R��ظ;��3����O��).�h�&@Oj�*Z��J�+*Agx;3��~:���뾄t����ؓ\׬�Ε���t���=��L����9�0֣���X����w�}V� �8˗�*Sk��vqW�k�u�_�����z?|�A���<�^��1������6��@K��ϑ����L��T��ʋ����L�7r�;m��g�BY`P3g��R`���;�k(�G`;=h@�C�z�>��Q��8���C��C~ �1��Q��}�އ�o>�]ȾvG6�ѐ"���C�(Mc�_�a�z}6��Bd3�\�I��u�����+ǜ}�k�J+���AM���E>oP���qM��O
��.Ȉ�
ȎS3F-=t�?�uȘBɢ��->6{�����l�kK���>Ec�~����?RW2���I��y���L��|
V@���dn������h�jX�ҍ��FJ\Cx2�<x�ty��Wj�]_�e>�g�F:��,,vW_m6+��7iV�JS��VF{��Ju����ւ+,^�� �h�{'G�AꬳɌ+�x�t}��٥NA��l@���qn�k��QPh6�ne�x:�������v}G-+�E^�b������GS�&����^MR�.��x��x��`�Ĩ�F[eR�J^氨�纾�Ύ��kM�13�9Uq3�!�G/H��ˁ��� W�/�!6�{a�)4S(��H����y�:��%�a ^�k�M�d�SPs(�ӂS��D�<s�#;N�o���C/M�EϢ�\^1����4�<vn���b����u���68O(��(�7�\.���%�cx,wk�E�Ue�9je�#���1��,�Ր���4+9R|t��ԑje� �L�z��5&�x�&�1K�
~�7�GM�EU�f�/+3�cZ��(M��Ҳ>b�ք�d��E���J_�D����T^jI�߉T���=�����Z��B:�������lĶ��;-�����1��0�jshϢ�|�����1�#���H��\�C�|�M�Hd�ڿ��/����^���wm}:X�!��8���X��@�d �����D�ā��9�z���������.��Ouw}���򠝫�-p0m�r6���rD�-#n���X����2"DÚ"�1W�l98�T���|!c�ί�r�A�M�.���6e�\�މ\�q����K�o�fUu��5����EГ�`{��[��}+~�۰�Df�p� �����i�(��$~���Ḫ�	H6� ��� Е����#J>���w	t�i�t���B,�s�M�B�#H����}LI{�Onkϩ��63��
,q?��U�� 
J^z��v	K���h@%��8b�6���n٧��  �0��S]�:��6��ڇ���fl2&�?g��p���Oh�x���N�0[W�&P@��~����aɞ�4��0�lX��o���M�/�b��X�}8�����?�r�z#�M�8�u�:����!�Ѧtj���CeT���e:��Il-�\�5vW0�9��y�X	?�P!)L��n���0��N~�OhM�'�Vn�o/�����hs��_��7��ߕ�EO����
���ĉ�>��l���{�L	d¡C���n�3�΍?�'�<x��>�Ca���'W��Ym�)��զ=(?�6����O��u�7���_�ʳO���o!�">T2�@�Ź�J��ڨ����i��������ã)qr���/�o��D�g�ι�"d{H�Գ �Dh�x-�!s1�MH+XQ����/�<�*�b�3��� i�_�������O��b�V	��փҁ�З`�l5s��8EbV�t�Gd�w�؉Gj~�G����5^�n�xj��3poF�� ���;>+���
��m,��ڛf>*O�NI�o��6��@.�1�p����ي>���1�F��v�}�O�Cb�7��t~�=�����L���8]X����*.K�׹Q¿}^��m~�L�qi��~Խ���[��Z�q�K��\�+�����Io�sl�G�t7Fr��x f��)��ʾ,b��*T�ɑ��0n��C=�dɨ�񌯕�el��i��n�DLM}��l+#�ɉ<*Ɵ���8!DV��%�;���4�2���ϼJ���C EA��%N��);��Uc�GR(x4K���$ ���bj'����	�D�VuV#��f�۹�4��A�@���d�E"��g�X
/����Q�*7�e4��u���z���%�]�z�)g$�ԏM���Ϣ�h�!���.�"?�F����l���m��՜���|c��l�D�5mA. ���!��Z�^9����E.�������*��uk
��)}!�_d���s}N��kh�$g�N�� +[���'��(~�30m���3��x�R�m�K&�%ṗ���Ld�I�\a��bA�p�1&��ڃΪ� ��E����龂��cTG�����P���ZU,:�\���I����±�N>U.�B�97ߌ�HT�0�n7�E���f(�7��L1�$A��eR�b��+�è7;��e�I����/��=�":z�Ϛ��}�ŭ�uN��8�9����Ƀ�q��u�� XE>�ViE��>U�c��zmi}��8�P��>�!}u㕡���mP����!���8i��\�`��m�l��i�B��D�jRF}��c��O#�h��y���y�����bx�/�[��O�Q!�s!�ɭ#�S�Y�#����*����(�E���X�(8v�'�	"��t̅,F�(�ñ��`���2��y�/���=���.@��DH�{(��5���j3�rLɚ:vz>�i�Ab�ir�z�}!}��	�d��&�R����B��=u|�\��6�,����;\U%�W� ���g���k�)�]��7|S���
��#h�����Q��: oXU�T��}u���0�g�+�Ѝ��I(�����F'�xO�Q�"�I���n��X��ik�>L�}�	(1� �{A-K��9�g��|=�q�dKC+&W��ϘK�3�+�^3��/7^��1[Gr���:�b O���2�Ӕ���c�7�[N��F@Ǆ4�k�j�(�C�,��gNMZ�e�i�R��?}��'V��Og^��8&�cPh�c%`"a���1{��v�Я8�U\����_	��#z$O&iM��l���U�A?�B�A��ɸm��o�ݎ�	�I���6� |��8j��M��ܵ�����G�u�:�b�2:e���崡M�;!� z��8�q>ubd�sO1ɭ'� ����֜�� �j54�R�K$�"OE�Z΅#�1��<4���� фv�ڃ��L�I�V3$wB��^Ah�+����G��l�d�8�2�MK.�*�@Bb����cRN6����ҭ~��ˇ�:Hok�U�0��\<&��d��	>�=:6���Q'U�~-��g=�T�M��� p@%��Ԃ'��A٪�P�$[�b0����5k�-�`L�� *��,� �s��u�AOcbș*Ry� CO���#EMp�ôWL�l�ZG�"Hm[-�B�
��G]�0V���?�y��ȷ���-�(��'L��I��������0F�Dl��6�o��`s�O1
G�QL�3��5�.��an��s�y�h�ŖeqGУp��G ��[�K�*�t�Mn,�;H�2wO�wZ醋\��;rsŰ��pw'CBo�t	jf�0�%,;�/�NlX�4	����?�Y-�>��?�z=��*����$�ż�
_�\�&����KE=�#޽%�x(?�S����|���(��|�h�In��dΫ����ߛ	��F�![/`���M�h�0ܒ�����L#�P���;��-��1
�\[�IX�B�Ƚ@**�.�I���Л79b�n��/���JT=�����iY���*�/_3�\�[9uQ��:��?nfn@q���!��]#�s�6�B1�9f��n�� ����q���
��\*�M61�I�8�>��lZQz�B�{��qHtr�:� �����E�Yu���E�@�g�4�?�,�*�T��s�½9�#N���Ez6e��	�������t~�y{��dܯi��M�aS�;J��х��>���sN�*�����1c�'aK�pt�<� ���a<·��P��*�~4�����pccU8�o�8����R�R,�wI�N;�Й#`v�Yj�J�S�f}�o 4�qQv��~k��n�:p-�i��ix��8$���s��*��4Y�j��coõ�S$�ʌ��_�u��"q��^*�ZG��]Î�x@J_��F��rJ ����QW82ͫ�L�ij���X؂�jY�nv$�sW1.����P�7�E&�ǩ�?�4~���V	� �?���X��b&�v����r�0߸A~�h7F^w����i�m�*��k>�?���˜ڞA}�.���,3t��d���Lk��צ��tb_��m������Q����+P�=��w�2�#�?9n�Q�Iy��8���V~$b�)E���up���t'�n�J��C� :���$������%�y��	�e��TCt�ǃ����e)Z�}`66ѸF������%b�eh�U��ac"��@}@�2��Os,����'��V�M�-�v��:��c5�rÖ��X#��`�iξ`?U�d�m�1N�N:Q k2n	�o)�_	Н5����і�i�É.H;Ƞ�,${~¶�,�)
G�?\C�'�'�y��<����H���!�v��k7�ܼ�z�;ˈ��ަ���T�^�|��:��\��E|�ty��\�D������"Yt�@	&K,��.��G.t3�=�H�����3��K֪a���T1#x3�<��LAꛏ�
�vA�g��pGW����1F()e#����	�3�ˊ�_*%N���/���rk��ԇ��Ф� �U6���+8��
gro���,�`�,n���ʛR)4����6�:�h����&%@H��3M�m�C/b���
��8�R��RMo�'��	��9,�m���6�i�A.UK���Xi7V�,�Β+ݫ�u9Jt� �3eF�-&��߶��)��{�o��N� v��B���.p_�T�\U��8l��b��d�P�|7�*��B�3��:�+DQ���RPGk��ɓ=f}�7���N3���D;/V@��G_U����3m����5���j���i��s/�.$p�XQ�#B`��ѧ��:�c�d��4�u
�w�@��W���3���`�4a��E�S��W� Ј/4�+�TȠ�o!Q����=�1��8 ��}1��(��g1&?��zC�j�u<�	�'��Xf�����]l��~-�!+6�ʞ{���`���{�`P�'�{Lm����`�;�5`S¹�I`B�@��˱���Xv��`Y���3�dP�L]e��z���Vb_�=�MrN��a��&���h��	�~F��N=,{c������Oz*��2N�=�:�ԻN��R3���v{���O<`��T��$���a+4��3�d#�MKg��?z^f�,a{�f��-�*�0>�~{��u�?�lj���h�X�C�I�����3㈯"|*=�x}e��>�g�|+��
oq`T��Q�t �f?�_"�,�ǚ��g��Њ�"2�)�NH�����J���|�PԹ&k�+%]H?fJBT郩~��@�k��=�����0�!�t��wM�ȱ�7%�+� D���k:D��v�p
cR��E6��Lg
�y,��Y������1H/ND�������q=����Q"�ݴ-�I��G��g�Ώ�t'A��:������kh
jP�Ql�����G��,X�۽��jl9$33K�.��2�,�E� }�@�f���[�[tje�x�G��|�����]S6�F��\U,Hl����@x柑wm������?��U���գ��0���eTK�C���@� �M�C*-I��FB��+.	��k��f�gϘ@�I��|~�;r�7L�f�;Z�/?���.�!�t���?�?#�4Q'�zr��LGU��J�0�m�`�k�S��=}�{k�~��v����C�gT�]�
R�L���P#<n d������.t���@Z�6w���,���F�.����%f��C<���ˬQI[f��;�c�_*�_}�I9B�u��.�_���yO���M�� ��Üq"���\��v��e��J��V�+U��g���t��8Ơ�	��	��Z{���SXk�����]����n s�s�"6<|Kf�!�D����qE@����:���zWB��WeJ�������_�-l��m����F����3���F��0Z�86�!�̅|��R���(������Tϱ18FĞɖ���w����p;ݹ�"��AdB!�
����{�M�=�{�'qPJqkST���s$F6�Euk��ϱ)�ou�%�S��F�U{��t?�隣b*Rc-�}��t@��`�ϣ*�-����9�����#@U��3���ew��L����h���v���0w5"����m�´�	<FzK���������RRRR��@9Nc�b ��O��
p�`+I��٥հØ�q�/lUd'߫1�p�}Q5ZE����� ��3$a�:�&��y��}�肍jǽ7*��f=g���g�Gݺ�=�q{�]�b`�h�;�Ue^z���Z2s�F�\��%��������;�'0�N��+��k_�F\����&�0J�E�*�!�\R�D�T��J���-*!�^	���V����ꥫj�?��ٕ�f�+�9^4��p!�O<�}&�ʜ5>����������)��R[��u���z%�\���(�F��@��mcV|��C
*bu�eU��ٯ]^np��1�Ŝ� �ѱ��d�c?�v@FT*���/%1��WDQ�!ҧ `\�"�	����(��pG��/0w���Jjњ�V�݁+�A��A���s�_{�)��v%��d�C)���>گ(�����a�yh��P6o�����VT�L`qJ��E��� ����qg<��ߛ;l�Y:h��&\���S�Hk��z�m���a��6����_䐇���+�����.��G����������$�N
DI���ܺ�T�HpzJ�P�1A��gGx��zʡ���@LG�/�Xɳ���1�h�tK�C�;�=[�S۵}���~�tɗ9s�u�Z��vu9oP�7+��$���U�(,�mV8h�*~�W;�E@��E0�Ub�� ��8�VL�5���B-��/&��;<��n��S����M��ӌ�/�YOn�.u*�R'����nx��xV0�s��,X��WDHzۀ7q4ǝ{M�c����}�,�����'�#y�	��c�� z����[GY$1P@>6z�+������h��5��:L�a�2�令!�F����	���5�!���]Ԇ0���=���4�n���d�:�Gi	�z٦���u�3ɪ(���6����Ә\u6��9�����u�+���PQ�H�j�������yh��t=��?S�Ξu�����&����n�U���w�ZZ�F��aY��G;C�q�}�&F��)�V�)ٰ����vV�aNջ��t�2q�J�)����*W21uv��7�r���p֮�!�K��s�9Md�g���9�Z~¯~�%������X0G~��L	��wJj2����t��Qd�'�y-j�_���	|�x����X�D\��ӹ�۵�ҋn ���­�o��f�}U�����G,A����O=}`����X�Q�w�Hڳ�՞��gh�#�!�Ef!��f�ox�����ƽV�x��B�����Թ��%�_k�l�����L���3�rd�������_�>o6`3�7 @���),�Eݷ�C���1��6@����
Z��X������cXppt��ו�����2�G��I�
���-X���8[Y.'H�M0�0}y�(ZTAA�v�)���]c��zeg�:EL;ICn��2_+��/�;]و2�ئf���|s=K�gji�*�\"��G���6T�Zj�3#j>� p������ ����&�����"쎪��b'ֈE�o�����$�����I)�/�������4�ȇ���Ui�%�b3��V����
W�H5Gae�/�n|ؼdeâ(��|`:�������h@��`�!�a�1�%�#�]��a'|NS���;��z9@�l���^�
���>�R��̺'À�G
z�R��x{�?� �b����h��
��Xz�n�Z8�V���	�(Ehg��«԰J��E]��M]�w��2�(�,��3�b+^�Z�c�ʄꚤ���/��Ԃ"ooL��`p��'�~p�y?2�1z�<�e㑐��Q�<mG�gw����,Ȋ��n�g#G��TT@��%��7=g{y*=���O'l�!����I���F:��������弭��EݯQ^$̶��ߟ���܃�[iw�G��_3�e��u��쭬��I.温}�k�&���l�,ο����~YW%���w7�6+��L�	��q����mX�~4�^�j�>}Ab+h��6�?�N"�lR^��+O��a1ߒ��ؚõo�A��9�a�2L0i���ah�Y���,l�E��FG���
0*gיe��綑��@g�-\>��?���n�MT�-׬vq�BK)5N�~�^>��(��=t��b��U��Ս}(��t�a(:��7�P����K��:l�.gf�6��1�-�V�94�`c�)7V���v.��U(*�ے�X���Qu]���}���r��i�і���U�|+��)���n�MBu���oN��'��$���`�V<��Juz��TV~�%~!g�c�H��j3���l%]�ܷl��~�H�R���{��Ez$@���^<#�V yIM�օ�y@w��'��l��0C��-�-�������6�89Y�s�3��m{���0PN��"��!a�<~����*�u_�J_q�*�&['��>m����Z�ᮺ���E���.�݄)�@{�kq�'=
������㽞$_s9��i�3�m��IQ "fr�d�7���a����d� �,��4�+i���FY� ���5g#�c���$�h��_���ǫF��E��6&�!����M�)�{;S��%#�(g�E�K	L��æ����\f��D˰QO%BL�ϼ��Ug2V�N�ħ��R��/��%`6�[���Fai��y�A�^�Me�3.�|&��������y�� ����pY��WM��������B�[R{np�d������E�6e��O+���=�H�T��o������i��Яr�M��� �m���#�EY����z�R��;����ý�f�/F��'��P�*d4���+o	=Y	���9؜}\�S: m��q"�����f�����+L��|��ֆ�1=�ϝ��yN����©��dK�W��nQ6��gq�kh�W��Ki�)mS���2Ћ����k�y�Q$���o�+�T����G�1��y*�ÖЉW	1���T����4�#eo�Z ̢���0�����&�^����������x�-\͖_]����U[0��T1uI���P&0�L�������%�}<h�_c&*�K|��ʛH�����U{�<�������Q~������Hm���'�=��à�Ms���W��Ӏ�9B<�f��9Nf@HM�cK�ݭ������Ũĥ��^;���Wk�G�W�8�Gg,Z����n�N�3�kU��y���/˧���{�W��v#����Q����`�4Ά��T��c�GL��y�Ԡ-U���Uq�\��H��&
%P���N�H�qD��H��6���H���g=$]��S�h�2�@Rc�x/�d��=����8� oF	�_��b5�ĜWO�m@��Ґ�#��]#'�cxҤ�C��𵙖~	m��V+��i���s�h�k{���w��I�\L���6�㮋���`yx�S}������٠���8s���	�^W�I���&\1pdR`{�B����i��C�b��Z?u̜�?)+��'M!�f���;rG|�Р� ����������l?��Vb���\A�Ҷ�^�z����wښ&V=�5���NldpSR��q'.��!���O)��/�U�O{%�r���ad�Py9���su}������鴓,�s���1_%�Hm�~&}zZ.ň`����ɽ�n$�"_�c���Ѷ��>x���j(����d*�ޠ�<Y���P� ��V_J�90��K=�`��ھmR�������\r/�#j���B�x���i�f�ZUS@ޛ�ɡ"]pĺ�� "`�JE�R��V%(�&P,��]ff���?O� �ਜ%1:�*��$#��-��?b�'Q���o	��'�Ї�й[5�u�.�,���.��'9rT#PF_
f���8iԃ�SK�;�(�߱a1��$�Ҽk��D�#�R�Yd>+*��,��7�N�ߓ�T7rr���"�6�����T	K�0@!=H��$Yp�+]qo�v���I��������Ԇx�S ,����@�>���ӎ;W�I�������,��	��a�yp+�"�vq)�
��c��?X���1j�T��C�Gz���Q�@��fuV���Me��_���o��?J��fE��1�&N�Q�Wk�ľ���w�?�:�Ċ[�9�	����`5QX��M؈�4Q+GX�y��>� ����Q9n+k���b���Q�yC�ϹᦵF�G���E�#�Ip�,���tn����ª�+mN��r���x���C�-�{�j�%C=�Xʘ4o���htnȤtj�D1!k-@����z��#�ݜ<�MjL8���ԧ<��e�S�6=���G��0�p�cvm"�v��:�乢��������#��q_����6׋�u��X�����E}�V�E-�xד���&pz�XP���B����T�d�7�OL�U��,�>�}C'���v��u^��A&�˻�E�Ԥ��z��ηf:�� �S�T
�ce��ߖ%���q�<H�z<4����/�C��_#v��)�O{�x�n�ը���R����NV���ݥ:�����~V�9e���h�#0�������b�K{\͢�WbҜA��s�9���ԣī����nX�)u�3�����܇cU�_0�e�!-~�\}e�95h���ܸ���e�Ȳc?�cg �B�7�A���3ElS�٠��,�*��x���_�������{I���^K~��Z%Φȷ�hy�����:z��Sm�cP O�a1���z^n��3N�4���]�]�S��8%�F�{GC-\0�<1�lV��<��SS64�.M)M��2!ۛ�̵�-��lG����A2~1Y/�������8��2wV� Z]f����鈕-���-�!OQfr��@-��j�
�F���K �4�	���G<���w���n�x���f��s$C�d�a>��,#��U��L���F�'+�� ����m�F�_�ŧ�������û��,��iQ��^}uE���;��xC��4+��;��+�a��s����@	p'�+ȍ�����K�m�'��[��~��R���t�ъF�Qk��G��4]I��N��3ז7��"I��Z?h7ݔ��J�;�֘CJ�Tv��4�xA���8��zm?�q��#w�����5�|���CkkN=�E��̯�>���Z�1jRF���l����(�l����\C>�7�h&T�W���;&D�xP�&:��(բ����>}�@���f�EZ��$��z�J{Ƴ�T��4� �z��:�,�h��{Q��;��J�-����8k��.>�(|83�b������ q����m�UVO��'�cDgw�.v��$6�ޭ�|-�a�飫��H�Sb�#�Κq��熫�(xm*L�7�x�}W����1�ZW�T�=������7�2�CI-�P(�"8K�(n����C4 $��/߭*��z� X���c?�����A�A�XB>X�u-�D:/�3F�PV������D]��f
����|��ZN]B �<��+LP�ѝ�÷��O�5��a<����<���9�:1��'�Mv�����q]���`pPc�8�Tz*�V���M�����/�36Q�r[��!G#+d�^��7�(,XJ �e8���S����enϏ�;)�5����j������F�נ�l��U.dGͷ<̫1s�����~�计��&Cz.�Lt�_B#���"R �Hy7)l<�e����u�fڵ��ؖu�
�d�ma������7��	�����#�u�',�PxP;���^V [�2��J@�$@M�C�Hw��ۘT��d*T��x��`�����[�J�~S�{���B`���٦ ��{�@�	}�ڟ2������Vj�]�$f���aY#��b�L$t{M�^mo�jؑ��rA�>��9��O�Q>0��:�i��rd���B�O��2��d����l�,�,�9w)��A*M��;��ָ�/ف��bde�L,J�`/��W�Y�ɇ;Y���L`4�؅UlݾƎݘ�����&O~���%n�L�>Դ�x��5U�2��#��_9�� @�)�z� 9�Z�� ��Ye ǃ��E��=����]m8S1�Gv�k�}>(uq\���}0��W.����^���\~S6�s��5w�c^9?�q*�qU��?��B�l����A�ra�f@�̔��f"Ҭ2���C���B���h�I�H8)h���]���قjaPZU�O(��Q;i�~U�������=�4��-�8��д�Q��Ogw���}��/f]�Z�=��j�B���W��b�hA ĐW�);?P��G�qSi�S�sz^�;����AP�H`�3Yt.��PrG��_�b��Գq�|i��Væ��}�P��� \��.���`�N]m���}�贮���޲Cd��'n�q|��~R�8]�򿌳��l����R�h�����B2}�^�����8R�s���c����O�T�3h��%] ��LqJ��/�F��t��� ���З�qKSau��"��ź�l_�
�B�}k���-N��b���'�a��kA}�ˉ�&21u��ٖK����m$�kn��u���@r�?�-@�P��[ؙ'��M��D�b:ƞto�����t�J{�ylH������^:\�!:/�$+����^�S8~�dò(�gA�.-��h�	�V��:�y|`rř�}A�dS0|.#������.���Eǩ���Dl�W�� ��J��&�E׸ز�'c�́�O��L��\z		�w|7��he���:������<�t�w�~�<�Y��cw�J�ߪ����"I�������δ��>퇂�vp�o	�5k�03�b3|�Ro
�d:"���~n������$+֋roU��y��o@�\��mvh3_�1
gEV�vTۧu��1��p�'���!���>\-rɖDD��:)ߑ�42���EL� zଷ�3���b�>7S@w5�RFh'?�8o�8_7�� ��ǒxVH��M"f�v���TT��2>Oi?W����DZz(�qE��%��~c��x�GAz^lt��l^�2�`�y�-�lJY�ۃ�}/��ܕڣEb�=)��[�W�ԑ���D��T|�3s����b>�C�``��T2�k
G�C�Ur8�{�`P�C<�n�Oa��D�� l����oG��+Ť��������ZM>Ú��ܤ�{4��������8H�������� ��2t��x���KJfZ�cc96��&\���Ϛ}�L8c9a��o|�NN`�!��7��VR}!$��/�g���꽲��<�L'�K��b
�!��!-�A���K��/#��Fo���͏W���ϵ����O��r�$ҟ׌fݰȷ�3+hIP��xC�����W�0�d?/�*�+K�A"��kc�:OQ��Y�S}t�������q�%����1�HzgSUQv	u+���E�jd&��j��R��V��x��A��(0�E��:N�r(;���z7�x0,�-����߅�"��z'��<y�	���p��{�mֻ�43�6mR�v,����_�7�fh<��5���Z�s+%-|��D�&� Z��3$�Z��fe0^�&�/�>r(���ߩ`xx�<<r����bKgDY!�3�s>�xo�2.b���:]$;�e�Mf/�90��n�+�t��4�C7���j���S�a&Hl
�y�N��Rc�VEEy�cSZ��|y�%'̣X�xG$6��ӏO�I�o��	�`5��f��������CZ������9Y������4���K�u�L�� k"��F��1�r��Ƶ;���:,8a�t�Z��Pٍm��$Ir��Z������3��6{�b��g3��y�]ɄGk�����~D���Tv  �M���:���p���n��w=I=B�;�FI5��%��v}�5__��s�*�<�J�� a�'4��-�^��c�8���F���%sE%�%/�P|�=�TQ2��ꅘ'֑z�7��cH6��ћL�����cʟ���r�kzcvX�^BHm�!q$#Yzi��O2&:�>m�v��I�\�܆��H	�l�*A7����y�yo-s���R��@�;�G�������#����-0�9�#ҟ��lk�.Y��2xp��5��A�U�1 �~ZD�/����&��_Z���=l��2F�t;��}T��?�|%Hj�`�6n�ͫ�j� �Qu{�1��:q���v3��5Y�P�|{����=�:pk�Շ,�f,�gy5�����񱋷�ǚ� U?3�h���.~�cR��)����7S}2UT "��?�1Y4*�2GQmT`��a�
>NN��㳾�'��v&���Co2|ɐ�ǯb�9!����v쥙>)�% ����ݪF����ࣸ�u�=4$�q:�J�$8�]��W����f�N5�pA9]e*�|���ݵ͸��@�v�)�����?9�H8�5�5�!nP
r�#_��k����_�x}B��~��g�듧����N'�҃,��n�e5���ќۚAd�fKf�:3��3����i2d-,9�J'z�\�n���"|���Ы�XF'c�$.��0�� 2�\^9�iTg(��)Z� $���g�>��l&��BK)ptŎTm�_���+�r��w�l�@��9v���7���8��%���/'�}HS�㌚��Jg!�!�˴݉�`�^
���䲼��Ǵ�5���sr�7|�tuj*"�$a���~�!���&\�����:�gG(,4�-� v�i�<m!��*]B@�̊�L7mԇ�M_�E����T[P]�.]�r)�M$�����$A61:,�;F�`�ϱ��և]�͊��u ��}ʂ�s���yI��,�f�.ׁ4����!,os�7%,�������o����Ę��`��R(4��}~�Yvo�5wy��gЗ��r�c��W����0?-#�����|9��`���aCA?�"ö�v�3�G3��9�2�U�ۻ��.��s���Mj�P�ŧ"��c��TX&y!���k��/�s�)�	Ȃ�3���c}�GِSYЗu��GQ.�D����6r���~�]���/V&"0�Q5R�Yd���ϡ��t"g(��c�����MC��D䴓&��Q��;:�M!�؆֫
n� zp?FPo�Ʈȭ�-�\SQ�D�(;�Aw���iR�`� KI����X�����?�����lQ� ���8=��a.�j�&�α���������Ƴ&m�`k�.!���ӶV�����;��Y�����'~�4̹+c ��Ŷgx�\���Fw���rP��Zpm@T|d�p�|ɠ{�Q0LMn�P-���YYP=]����U'���H�8�"���{��>���;���l�\P�"��WPc���
Ta�` �i?S6�(�uh����f.nсid�����$����ͰXs
�<kXs�~ T'�������$I�Wj�9F�]<E��r����f�
�2(Wޙ��4�>۵f,�m����	-Z�cP����z#�OS-��xe	��1�G͆QꌾШ�� h�Ӡ��c��M�r/�E�1�ݦŃ�l�r�C�J��|��a:�j��y�Ȉ�ror�d&q�D�G*K�RT�BJQr������$��*&�R��L8��c?͛YD��:?+�Qϲ>�C��a�)nQMb���������,S�s�l��Ͷ��;�q?N�z6R�)�	���;�����Ҡ��o��qv����9vb�`��a��tVhU��Wו�X(��n��<��؇�!7x�/f`6�I�}���wE�eIx�����%/s7��Ս��VPn�"�)h�]�
]�Z�L�}�*m`YIh2���|��Nb�m}�2���*{��h\�_#g����|ʗ>��3�;F�>l<��?U��P�0�S�d�@��e�=J�:��a�M��~X^�T�su��{*�g��`�=���V?;"Ѱo�4�K*�+��a��Q�F􋱀9Bq���I?q������9t
����P?��R$D�����i#y����d��բ�ga!�ta,�PcS����r°� � 2e�M���U�Y#@���!�^�lךT
� �U��P���.i#� U,���ԜwR6d�Yak?-%�bw���tӳp ���d�*�e���4~ �7*^��G�r�z���kuǓ1�ēG���s�F������/fH(�(����(�
Oɸ��hJ��#2�������xW�X��뫛��J/q��_�{���!�B�=��á���¿�va��v�7�'��()1I�U���_��}c������)$Ԇ��+�_ֿ�w�x8Iqɐ)v~p����z���lsD����=�;R�
ѧ`;M���8���TD�M/�/pq&��d#3���qƒ�(�oo4A��Q�2����C���W�ԧ(e�-�nވ����^+=f�a�7r��C|ʪS��׋T�&���$YA�H�W:ki�>�\waǠ��?�ޖ6� s �P}���m�pH����@�ϝ�L�}h�87�SpV��:�o���
��([�-�|j�E��=4֩�Gk���a��-��n��Gߪ'���$��c8����U�妿W�w��''�	��R�vK{�~�����o��o"{�Q�~ر�W,�'��� ���]�e�.XV�ԏ�w�3�QFJ+��Ĝ
�t-xJ�0~!#��͇�;4.���xfǭA�?/�}�S�O�ؚN*��|V�
(h�E�~ ��-���t��16_y��Z6��kaȌm�6_�n�t�mdC�%3�-=ģ�Fr�q�z���]k�M�p�F"`̛���D1��F"v����d��L~ �i�����Ƴ����k���ć��ո��w�u(�:/�>�.�$�ڀ��]�Ζ'��+��N^�ɻ�h��z��c����t�Fx{�<�0A<e��D	�!��[�	2%��,�mƟ�����F��-/	��2�����M�������)? l5�(��A��W;��s/�k��b���P����4�ӂ��/�))֋�l��>�X�us������ʱfU��R�b�
BC�vh��4���y���LL��\�_��{��l�{�xF�s�R�n�X�Y�O;��&l$�l�-����\�xE꼑�+�Oz���uo���l�%�y���?�톅Vm3�!�_jW]
T��~&�τ�MD�mѓy"CN�&�sn*�'�/"n����\��r.½3��]���e�^���K��`��Ӑ����1�z���x��ו-�h㢏z�(F�^����Eƫ�<m%��ͪ�M���p�\A}:t$r��ص��d&~��W������l����DF��l��B����H'��h���k'1��c����b���K��=�rӞ	�2c�Zz;|]�ȣɋ�z�|��tm�b7,�@娾���� i7'9�uI�����H���2���4_g�P�R�w�PA��$o��3�5��g�l?�=s��U|�b>)���hY��)�z��q��˿q%~�:E��J�9�p�A�9�i��T���x��W���Ly�����kS�ǯ�1��3^Ap0��F�1�B���'>^g��E����`��0���1��.*���D�U]�Dߖv6EBKs\W[^�6|#���u�]=��b�.4�#��5,/n���>������R�.��I���l���M�>���"����!`�����-h����8PK�u��tE��v��r�i�����]�7f$�6�S�P�@��6��a�'�t\>)�~�K�/^+�qY|O
0�g���"|�(L5�cIKW���V� d�<E�r珀��&7Z�{�UL�8���:�cQȬ	7��l����*zs�Fƺ?�
޵�*_"�RXWɔ��\5��4�����ޫo5lǰ5t�Y���W�Z-0U��oG#�����a���Z1	ϥ��֐��wT} ����CG'��M��n�� g��O�@b�}YA�ko�s�[��c��	�<���5�=��Rq�,j��|��,@O`Z���ϻ�y�x�B��F"幱5qH녕<~�f��E�c-�a%DH���Q�o��w�;LYǧ@��	(q�e��Y��۰2X�F�x��+��?�&�Kf!�x`��O�f��`�W?�T��^�k�J�KGZ9�/sҤ�ҕ�lJX�vr��g�w�2le݊��9��K�g�9z)}L魀_C���>�W��HF?c���@=�h`����g�-�~7�n�O�н�ֺ|����5��|��(�J̊hE�e)��I�̋<ܭ��Q{�m�D��$T8����`�N��vp	ڕ�j��H����m;�:%K��\H��l��ԃ
*���,--��k,I:�+T�DH?�z��Ԇb~s.�Qhٷ�S��8���lX��Nt����R�_�cg�ߦ �K��� �k�Xr<�%�t����FuM�������2�)>�?Жİ��v��w}{^��B�66R��p("����
��3�d7�����cI����2ś��,�ӣ�>#"m�����ε*��E�5Y����FE�_�A?�����`8�rI�����g��ʸ��WR.�����K�m�b�k'�r����T R9�,���;��gu��$7_C#���@��[]��߱u�U�h���l<%ŉ	��ҩ����z5yT��f[��ǟ��M`��:t�Q*�݇��7tY�8A�(��)�k|�ɢ��;��k�-~�	������l"i�]��ip�����qM�k�m��4�ay�L���jF&0[�7\��
)0 n ho=�u�7�dO5�R�Y�*Fr�����R���>�����e���� ��E�k���e^�:������[�:������ݧS�fu�����L��O�3��]����q��]�kg����k�E���Ib��`5��|щf?=�����p-��!��g��Ø�������d�)<���Z����|���T)��7
���D6.|X\��Mj��-��:�����~�����0u�E2� OSK>�� g_���)�[~�Is1��mz6,��S��!
���P��-� ��)�p<ohS���v]�f�o���oy�빪�|�sƅ;�+"ve$A�3����-�(vʓ��"qB"cWl�P�g@�Rc'6h�5�?c�Fr���L�e�Ϲ�c�CF�Ў+��v�0=�e2"��P��|<����?����m�^�)�W�6��P�@m�]zɢw���w��%�-M�٨�t��pʛ���ڹ^)ק�N�}��}�I
�@�g.�q$:����~]��M
�o�?�P��)�-I;x����;�.5-j�@�7�k6�j�v)ș׈�3�g�8�#��q��a����g>.����TT��q��a�ȿ�w&Hj�_��f�n�R�U��@�ڤ��"aV�U�5��G�S��*2���V��Q�u�&7V�V;�=���{�vI����UF��:E�RA�bƩ|�>g<(�G*�ռx�hAMI�ER)5��٠�^Ry^5���;�w��K��h���
��'�R#���HX�.�6�W^`�����&E�ZgT���PP��yxF�����tó�$���3�+nV�b*�dU�+�n�m���Y�/u�z�}c�:z��!L1�^�����P���H-�
�k�������}m���hA�/��do��I�6G<���G<�&�!2��p��@K��y��A(��{�ja��OY+�)��{�Y�
!�0>��0�>?�m��/;��N���.�,^�5Ae_�Bu4>��*r[�/�����v{��F�[4�� A'�i�W[qpj@v�-��W*�>�Ǟ��oy��E��ؼ�e�e�ʤ3 ߿���q;U����.i���-$�5C�ѭC&l]OP�#n�*����J�|��h:Ǔ��l��,�D��B���em�	L����+[aF0F�+'���W�@q�t���Z��E��3<���H�DOCn;�L&Wֹ�%'�?E& �;p�)>ux>���*��K�����PI�O����������82?�(���@/���䗭���NC�����R\I@e�\3���ǁ�(*�7�C&����CQ������L�[g���R��F���X�����tqu�"��ϲ���C�\Lc�F��d�߾��� �
���*�Ή��e-�<Y0���! Y;�"6
iDP�[Z�*&�a!��4B�̔������?���m�Z���٦�t�ǀ�Z�)4���m���AF`40��y���Lw��A_iu]�9�瘧<
N���i�H��o��6z K�hF�:4	���w�ܢ��7S%�6��v#���.F1�@w;�����&½4�6�l`N�% �:�~0�����㢸�-Q�E����E����*��[��}�H?��r=�x�`�[O�U�(���6�%tM�T��_5��gD�+�:�3�<^���b�1D��G+�|��4��TW��1A�;����Hs*� i�U�9�T?��a@��%���^K����i��ACP�:�S���wgt��I-�ӈ�ws�OH��9A�9��KA��A[fR�7��|�n��]u�=O���o�߸-z9+��Z?�; >S�I!��RG���[`WʰRe�Q'�IT�e�7�F�}�e����V�W
En�����5�AM	�<r~V�5ʽ�0><�.괌�ţ�G�\z�/��&������`��f��#�����!?lu���kT���dq֢#ӗf�(���W�"��iI\���`eya�J�o�_M�<O��-��7��秨dE �?��°���Nu%��e�®u(�G�vg��HbN�̏�?ҧ�>hc��\"�X��:(.k�L)�k��{��^����ǅ�K���z��ߍ�ݛr]f%�	�B߻g@P�<�e�o��@a�� ��R� ow����һ~�$W�,��D��6�Ȱ�ت�n��I&�ҧ�4Bg"�-�&��	0��+"I_�"?�%&��J[�:`�'b2�r�7þKo� �D�PW�Q�H��*Q�-4��bu�-��*N�w�p��w��Z		��D����{��Rˈ-(mn�R�^����[���{Å�YX�����t�0
6p"8O*(�h>l�f�2���y�h���W�d���_Wȃ��S�!n���lW(������`�h����a���y�4��Y�)�Ò87��C����ʫY�X�A���*"�g���pT
$��|8iM���Y����� ܃�^g�s(p����'�6l�%~�X���㺝�+�V�������c��	�XG�K��qQ����i��"�>���]��P�pÜ|4  �y��RϮ=�᳒�I7��\ļ���x�
�O�%����`�SϓW��[`Ѩ/ѕ�Z�n,�7�r����Ѥg�I7�L�D��t��0!��e�=�$�7B�4��+c���oE�ӓ���0�p�-4!0���T�;e}��!fc��.�fO9�UL��ɜC�ծ^�!�r}��V�����e��9NV'K�E_��[+�5�i�7v`��.�فcC�N��B�Spu�@KP�^D뭹n�@V<��<���'U:B�]���|ݖZR�m�|��3�+��i�H$�&��Õ��j���c}k\B"1�O�g�o,�l�8�����r�섋��絳�� �w_),l�u�t���<b�v���|R;�su�������o���h�PuĔd�k�����ie,Fr���<J&��������ȍ�4���4\�'~��.�s2�%>��V��Q��):�^ii(zc'��Z�W��4��T�'���x��ΦP��YF��ܐ�Ո�RmĢ�;!l�[DQ	��OY�r��F"��iҵ�8�+�bz�5��DL�-|���ʙ��I~P�A.�<���ʔ����+ƀ��<1���X����!O���<J+�ȼ 4�zw�j�������(��	{����"A�Ϩ��/�A�4zs/�~(��Uhk��R����?�+�VFv�0�bӽ����uE������H�+G1����������d�L��$�\�-H4�Fuq_�7L1��imX��*�٤~s�VDT^ѢՌ�ݓ�2 ��K��|������	���%�=�3Zi$Q�*o��ؽ;��;�WEq�Ɛ��h���e�o<�m]��狴Yo�e��.ٯ�\���Y��^db}h���7�2�E8�]�/�|��ut|%2� 0/� h���Q�G(�u�l����%��t�x�s5�S�Mt'��#G��n���J�MW�֤a�^��A�<QMG_R�h�"T���>A�A�G�%� �t���}s�fbP��A˘��*���e��ۏw7*��4Y�h/���ޙ��,�9'��!�m���\=�8^W`0�F�����Wb]m�$����?8��:wo�I�od�6`�D�?�����k�;����J�,<�->��Vອ[�=���������h3���pE/UԨ��3$��S>��S�x���>O�:c(��v��ޢg`kh?(=��v
t��`����x�۬�C�����_U�v�!s���"(��3fؚ�z���$��p�����i��Hn�6lFR�	��S���='�8�\`�K���P�x�7�*�!	�@�c0��\�H��P�f��L/�C��ciR��cw} ��ai'U��5M�<����p�g�9����i�J����#)	ɹt����a���/ �3��S��=�Z�1��AF��օ���O`f'������F�*c &$���s^4�|b�"�&�g�����NjCi��W�䔠����f�|��a�M@��J�^=JS'	<�7i��\����z�ZQ�a�&9"*L���2�[a����O�\�˲ǫ��ͩ��0�`�}ς���# ��/m��""��"S��HT�
��~��u�� �;/c`���H�nR�����t����8J�*
��}�Ht���Ħ26�PsR.��d^�m��|���N���	����ԞKP��Lf��|: (�L��Y�0t�m��X*?C�/�LPh:�6��1t�v�N�uU�;�P������:�nU�5=�@�*�Vy����U.BÕ_(�ʼM�)Z�GD�[��;��>i|��+8���>E-*��Bq�3f��E���<[7؍
Ӷ����{\�v���K��r������n�4-W8HA�!r�mʦZ&��č�#Df��b�d{q(��o�������!^X��Q�&ylӶaʏ�n�F��X���hqM��Vyo��
��L~�ǎN�[!6�ۏUu3��	X�~�@���ut��'#N�[5��om%����U� )q��I�!��� OΎ�����+��H�p��+�7,�4�ь�.�Ek����ѻ欰x��	Bj`jh�����=��E�C�fH���0���,?���k�����<��#�'^S�p� d\�� �+�G���ɡ"�coۍ�tm��������2���};�je� ���/�f �cE�u9l�pC�/K���9�v�(�U�����-K��XV��E�|03��a6$�0M�%`�`��J�AHn��Y�q��v~ҋ��E<x+��"�ݔ ie�Ы��~Q���Yn��5-��9B��9<]*b�Ix&^�� (�^��qnF�U��
H�ыҭW��G�ނW�����)������=�ґO��M�5��y���l���|�vj�6�rjB�Ͽ��^`>��9�{4	����c����*���R/Tna'󴊤|�<��@�����pv�#�����M-�{��B�+���(4���M��LV�c�
SP��7���������N�gPQ�Jַ�h�T�!V���NFI���$�}�~"�1�Ϡ�w������ܛ���0.°CD�];�n�W;��Z/�q�
���c5�S���(��2����̒k/��t;k4c��a��<��4��N���<�Sr�&/!pO1��c��3���{~A�]��1�3�}��=�5,�{����g����98B��dm5۠ڟ���]z�Z�o�t͹�E&�+���r���,��ń���u�<w�g�T�R7E5���p,<���Qԧ��Y�)� �x�o�HF4���
�H_j�v7��}�|K�T�qi ��.�oC;|k,ߢ5+��$���vB��ۼ����P:?Z�Ku�������ZՋ�3�!>�H|'BX�R_�z��a��E�#�A�6����|@9�3@[��ٕ=X�d#3P��	C�_�ɱIՕm>T;$�>�p��$��n��n��$^˙偬ϓ0�W �!�w����NVM
��$�Ć�10N�*,[[����+I���.�,����CaO������cnN��4��!��j~UX>fh�QDu�?e"#��?��H,P�o�d�3!Hۦ��F�|��0E5���s"Z�MDs`�E'��E$��B��@��� W��CU&�� �/K&�~1)���_��:������T�[�������0���h˜
Bf��3���SJ�P}�h\0�oB�IVVi�_L_��&� g{�*S��0�;³��-e�X�����1*ۧ��uZ��Nl
z��-�A4���P����:̮5�֟�ũ����|�0;�hg|ߪa��k�� R|&W=Al�e9���&¦Rߪ��t4�֐���6M�hf�'��C�	µv�B�M���$�4�3j%�at]��U��3.D�~�Sd�gx��]��qH�����ru���A ��?�z��
�CN��x�Hv4��8��K��M����h`3��^�8���2İg�E]����k���H���y-��ymxsMc�[i;xN9��[HkH	k@K~�J������bX�W	���6S
D��۽$`�b�F�$
����	'��}����Zv;#F�i3X�[t��u[_�
A��dL�XgO��)|X���7)����CtJ�u�E\����A�I�P�T��TK���������тw��U�ԝ:_�J @4��k�)�<npÌnmKg�0��r��a�$ۡQO�i�a������	���D�C���C-R�£��,6�(Z;��Ću����s�@��r�V�?���:���4M�� �&�:�.����W._�a��X��r�{Ǝ0���T��e<�{M���Ö�-��O!��?�a^��u`uJ����������7������M�ދ`}�&	�,�r�1��h�I#�b�	).� ��3=Y�&�p�ǝ?��ܸ1:v���R��5۾+Q��x��5Q9�D�x�$BO��M@��|S�kH�D�7�K�� �:�ld���f7��ߦG�30�L�,Ǹ2�9�>|i�G�|q('RM$�V<44��#��	Y�R�7���=�#�$�>[���*��N|��cmT�oi��Y?/􌧽~�������(���L\q��#��o%�j�.KUp�,O;
���?y�2 ��?ꉒ+�17X��ܤ���� q��x(���i���u@ ��G��L.��Cx��7�3;
�z�#���|$�Í�J��/?sX��{�3�py�����Q�����G���^@��������,S������J�OO��i����eu����0:n�p[߶B&�lOr��.��H�K�mU A9�4:r\+ ���o��^����Ʀ�7�0��"�IQ��P�b�im�=��@��_�����̒[��^����xes��};���S��9u�	o�(�7��������cc�nO�挍��mv����&Ҩ�̼n��:��g-UHfӖ����&��)����|�xӃaћ�׀�:�ǽ\�U�4�Hk��Y�L����i
��K����ͼ�/���6}c&�e�&�IO*Y8���mN����Ħ�w�0cx2�s�nD��D��IN�e��2�_F�>妙��'V}GW�5wwsz�&�UI�}�隻�
[���^V��}>����']�+��*^���~�i)��q�}j+��J��\��ꈷ;�;�&�[Vf4���lQ�I#*Y�M���/�Y�{��c����Y��4��Z��C���ȁn��t,�%���?)�F��O�Z��ZZ��J�NP�c�ƍȼ�r#*��=����j�w�q���+䗄[����[,��_~e�q
G�;s�]V7��+�a0b]�n�7k�Y#tC�)F�F���5/��Z� �Ͷ)�dU�**���g��t`@��NG��Sn��MYMd��V�1�����gm���h���a�����U����e�{�'��e�<��}�����3G�؈�4O��W�^*_��acW������I"$a�����a�K�aa�U�xJ��;-�&�FmL�@5L��׎w-lX�F�t����/���N�+�|Hxws%l��2�	�k��	v�̤�4�	�D����&�t5V�t�$O�+c}�Y^�ىwڍ�s�Ǆ��:�aֵp^G �0ND�gl��	dA�v�����޼d�md�Ǩ�ߗ-3$���sC<��<A��J����H��br�;3K���.E!�@����w�E�����E��G�`��+�_qd��]�e8��P> ����֪���/esL�ё�a�G4��������aO���3FG�*V����i^��۷n���,	{�[�c_��� �3���
���K�:��]/R�T�X���E,�[��'&��4'Ղ���Y��m\C�`vH5�
��b�fAIL�G�J�6����y�ʭ�	�1�1���3�X����e��I�$��j�cӊ��N��oR�}/U,,a]�$����[���S5QS�M�P�*��SR�.�b�����BF���=)��E�Fx�0a�$l�]��Q騡��ko�n9e�tk��r�U��ΰ
���Js4DF f�Z�a@ �֩2 ���x8�m�r��H�g�y��t�� QI��p�c�|�&v5^���PxƊ>z
����iY��4���<���z/���e{��\�b�[d�r�fٵ��2b�5��_Q �ֆ�{<��Z[����{�������{w�D!�;=l *j-b��J2"`�l�����{��T�w��ٿ)LL'�6ܲ�I��>�5��s�� �l�2���H<S���~.��Y������4�g�r���Յ��ƭ;�;-�|��9�{��h��В`A���e[�f��`:�^63uV��Y�$I�W]ӟ	�Wr$b��m@�m�O`S��|R�bvF���C�C`aS*��(��3��#0��?�5� ��8���9ł�3fc��^D�»��{ؤ��ߞN�#�0��-4�����|�fif�h4���8�g�Z��Ţ���&�W�KLa�1/ǄqH{���u���n^Q=����'�M�i�QN-1̥k�i����'$����M�j����Se4��̓�ܢ^��hI����cy��M���bkuR��L�}/o͟�'g�/�r��$]��ہ}�ٲ� ����=%bN���V�b����aE���b��h>���m�?�V`z��8aq�p���.t>�-���K��S���vi���*���+��9�ٜv�o�C{ԁ�Q5S]n�C�Z{�whO�2������Ԣ_�G�]&M3X���`b�s��FLQ�	i���8�_�y,^���m2A��ɵL�)�ꋭLkj�2a�J��+�?���\=�!��.�i�R���v��?���o�}`�[�
�rU���e��>�y��R���(�9�b=]]z�����|�k�|�$p���\�t0��}�	C_V0t�0 �C��W^��v�2��ɚ�	�7�mVىSc�����F}������t��8���O�O���d��-/�FZ�+�&i栎�r��-�����ax�3�u��}����ՄU7�sb��V��J7 j��ðG-������F�[�*�Z�B9<� �	TuZCc/4R8��9�]�t ��J�5FCw���|\���ʮQ%wZ���X�Ҝ`����� N���J?D^�ޯ��WI3��e�u��d�a\{�
pxj��FS/vhOX���ʱ�\�$��B�R��� G��p��A�gR
��a�/��^M�	v�=&�pg���eG&<МX��~�_�AE�M�X)UX�[����#3��bØQ�@�V�dg;�7�R-ՈT}h�M���nWni�3�ȃ����X(_1��b�e��A�-��Ba(b| �>��t���}֫�B�̸"7V��F�!����bfcvC��8�q�M5t�.�Hh��*d���R��2����N��E22��h�=�n��̡4�����C��8_;��;���|v�Tj0�G@�JX�fn�m�����)�a���>qNu�na�`7�|$RT:����q��RI��T����������������Ց9�%G�ce�R
����j���ċ^��",�]S��u�ً�Eu��h�nw�d�g%��	�C���Q�\*�W>�59���l��+v�M��)D���=-3�/H�[�~mR�����vL�~`i��!5��|m�)H�
p�yR�#��]�t�$Ǡ��>����h_ۅے;H��K�oȅ+h�v�˒��-����\v���,��n����+���7	7���)'��9���_�<�ϝ	Cݩ�U����)Mey$l<�w�L���nr������y7&�|��E�ޒ�	� ��9#`�m�� bSۗ	,8����yG���w�I�T'�c0<�d�o�P���:��-pNk뭢�M|�h���@ۮ��#g�s"o�ѽ�
 ��X����W&��^�HKPH�v�%A��0�h���Ԓ/2��<���ӛ�ԒMaffTz�<���X�pՑz�JA�j���D�W"�C�]\����⋮�H��_@<Ƚ��R�"�:�p<(y���&�{s�凵�cN�Q�ڹM�'���f���~c}�ͣ��e:A�O��)�I�b��ү
|�^�S��3��dA.�@7�I��ZZ�I��n�W�������;ľ�kBQ�wVX%�Mc�^�L ��1+ta��>F����J�k��萀|0�V���w�z>�d����쉠R��"5*0�����%�6p_�܍����h� �zR�)0�B��ܾ��K>T��`��̼U,W���;�pp4[���y����`}��Y���(����7Z����C<��R;���x�;~u7M'��ٲN	��("��`l����j��j�[y¥O j$˄��}���ڒa,�ҕ��)����_�2�t�A���'�g�6P��@����S�R.��������~2T_"��.*�᭡��Sݡ���
��~�$6%��zЦ�m������Bq�g�~�Eߟ�p��y��a��\Nci)7�lR�~]���&S����*�}�����54J��Ȣ�.w5u�j�W��n�w�[l��br�ӬH>��r�*�4 PDY�r�:޺L t��mn��(���ϙ �f3.A!�]���:��4p�O:�-8űB��F�l�Ǽ�0�bw|�;��k�Ƌ��Ҍ��BY'�9�E���xN�麬�-�vL��E�Tt��������*a� �����
�q�K꓀d����M��w��K�22{9�B;��] ��S��`3e���.����[{X��喤m���ӏ���W��e l=�f�ͭ���/�(���%Ox��$f�d4�����ܰʱ���e��Y�^�B_|�Za$�S{�9���E �̅�����J�d�Y�~�Czh�A1rCĎs�;
�V�����JE7V����UD�v� ��uc�$j�	�[���؏�$)�����"��G�����M���	�P�n�Tӓ�rl�rP��Fīk#uuӏw���O]K���3'�ŏ��6;6Gx��`�`c����SKq�تs�;S�d�w&ໄe���|Qӧz
�.D����xjoU_ei���s_��(%�QXH��	W_��Y���့͞q1N[�D�I�q|���+���é������f+�yt|�^�#���m!�<�y֘��<��>T.�0�{�,Z�ۅ��C�d��$��Z��׬J�W`"��
�����a��F���t�ףlm��[��w���e{:N��N�Y��� ]}��>�	�1q��W�b��2�W+�[-�N=:���/��O5�\��D�%�45mX}��t��D����Io�Z6}2�0>������G-�@u�?��ҁ_��?{t��Ȅ� �ש!���+�}V�u�Qɧ6�#aZ\��vh���(�����{7V���-^�-���j3]wv��_]��HA�p6�Q�����O��o���Q�7#�i@'�#��م�؄��t��!.�݂ UX�:01����o���Nh��Ţ��ʢ|�s^q0���bS��%Z���oh��Em���@U�C[Ćrt?�����`P�ݨ�������Q�­̱�o"w)ţ:1�����c����ZR|���v<�=�=�i��Cv��T��]I-#���*�����I���� ��8��"�k����b��z�9�7��H��f�]
\h��bZ�)1NZjeĻI�����J��c��J�κx�;WjMQ����c�@S?�xrA��G�F���ߣq���w�_6�ܵQ\Z�Z/2�b�=L �p�]Yz*���6����\������r[�i���%��(��F-؍�!u1>��.����[6YAё����8�[��Jx�L���N�x�w�Lٵ �����9�>�O�H��o-p��I���,�23d'�r����f���Y��(m��?�6���V"n�G�t�Z@�\��k�涞. �n�TW���<��3����P�,;c�k9���V;$�]������f#x>y	@N�AQ���`gZ���V�A?4��d�ǫd���^������M2l�eG�5��k�2�-��չ�[������г��m�t��6�1�"��ҼR�3vF.1=gտg�z��t:ҝ���3c���=���fߌ����2�����?��u���|��R��a���J�?x�6��8�_q�M�۵Ǭf������n���J������[�H�R��Ͼ:%b�c���n*tJ<���A�QǪ������JG����P���^��]b�抚n�^�`��e�Ť+�+v7?�Ш�`@H�N����LF�3��a�t�f/#�X���m�6{Yws�97�������s�I;zR�8Q�r/�迋1�b�6�LY@G������V���R��͕��;�?��cVCR��o�{�O�V�fA�j�n��� �4S����B#|:�����-��-��}�Ad9j��/L�����G--�]��FA�'�lM7�u�~�m���&L�x(j��j,���r���B*�5�k���������|�����Ӏ�B�o2��}��Q1�, �F/`oP<�cq���h`������xP�[5��^��h��=eK�<���L�Oժ�����;��Ԑ����[WQbI�����x��?��}����r���z����E��`�9a���`��?K����ٶ��-�
V1F���w�@=�}���>]Ӂc�١9WzGv܍�L�pVKM�*>�y	]�q'�HW5; ؍�/A���h������5�^�����ڔ�{��xp��) }�>-��P������X��9g��{{�����҉�h������j������`��Eb#�|�Y�E�>��䷟�ROZhT���L�r��(�a"!�!���%�o���Kz;�t��u�X��R�d*�ަ⿶4�٩��0��zL��.��%\�c�������@		��ԋ^DdƬ�)�iyoR}�/�9��
v��lT�M�	Ŷ�ג#�_�w�	���,�߱��q��2>������AOP�;u\��U"ԄМr�]:J:��ɝ%O�Vǋq��rEZӁ%x��e�x�p-��d�4u�m�;m�:Y=0��Z�#����u��3x�����ota��5�sjz����4�(չs�^����yv�����M�Qf�ģ��)�FMs�y���`�Y��o}�Nn�2S3`�'k�WŻ"�1qꫬ[B�0`)�/�L��ex:Κ����
U��rY8#	T@�#'U	$��z;��9��J���[��,k����|qAJY�j1�%�	�
a��Uv3y���/(�`�J�eb�	�{E�7�Z�ꎶ��:��s|Ih�jb���i�>��IZz����jI]gfdbE�.��|읾49�yқ���+����,����1�/K{q%<���D�
t��L�lX�6��@u��?>CjИ[W���'�tg�1�]����"��{:�Ɗ���k�'�{����ӯ �A����8��;J �]�j���F�P�)e5p�ߩ��]���ڈN8�T��d�I�^v��O�\u�Ǚ����Q�'#4YZ���5���Oip�lt�XG�^(����>������b���������ud<�#�����1#P�`0�֪$�>�)b�Gՙ�E�+��V���J����lo����s���8�P3��3��k\�p���K�D���Q�,�=ckz�A�M��z��@;[�D���3J:s�㗼�P��@��N�wi�S���k���9�&l�BU3���D�͠��xuK׿��#�)�K�R���1&N�Q`���cy�4-J�#g$�HHs�-~�)&�$F]��X��n?d�p
)�C߸]|BE���k��̀�;�'Oױ��a�m�U���<�6�G��4k��6��^`���&M���Ҁ�_�g
�0n��sS����#�����ƫ�>�N޺M��5��Zr�b��=>�@�y�XcC_��3�jU�iv̴�������{�Bvy�Ϲ�8Qr,U��Wc݊$��  ���mBFp��3v?n�#e��n���Q�zV�� ��g#ij��q`!?#�-0ETg�8�s�9Ww1_�*%)������U��dKq����8F�����7�Er��픵\���^��tz	��X�+T���^��_�j���\�\��@����W��]�:��щM�ZK}3���X�e�j�7g����.8~
��w̋e�l*���F���VR\��"M�[r�T�,����t��D��A�	}�� ��z[���;?$34�P��g^.�0��	��_	F~S�bP��ۛE�4|����dA��G�w"2�H��}8�-r�E 	m�~ét�Q�n��t��&�t����>>m��<rS��䡧��;��/|��']���_;s�=�80A���&��bc������ko�C*>��#V/΄:P�͘ݰ�T��t˂u�]Ĭs�*���9+Q\�i]`��+�Պ)�k�8�;u7���pH��/	(O��M�x9�Ҕ�V�$W��Վ�1���tu���[(q,r� tn kD���] U#2�ކ��dJ�� Ԍ �&JZń�p��<��?t����4Zq6>���g{u���J'�e�.) �"N*T�f߅���|}Ok��˩DJKP��8CD��OY�2.�3XB� ֎�X��SmA�E��>�D·�d=�GMm�5���32��J�Q�.�a��'!�#��a�E{�t��K��)Z���޴d7�[Z������R����*����g�A�=I>�L?m�$:�`�2���d���)��+h����F�E���4@b�!b,H 
��s�t����������L�]fc�����c���Z�BSR����q�\L��>�$nXfNbO��,�	x���F�D�g����*���>U���X3�8�0�Y�3��lg2S�و����;�w���Q{���K��D���	8UW�("l��ֵpj����}������E�}��l�����O�(����o�y�	���G໎����?mݬt[�܎���
�9�V���i�׳��"{�-Y:�yӆ.ʮ�`A/	A�c
�;��'��Ty�ѵ��$,�͉��� �`|u�6�Ϳj"��Z�U:~���-b1�4�X�u0���k�gp/�����t�Mf�)������M���- �Kٲ1��{�����4Z�tt��)�w�����{
[~���*�p�b�>�Z|B�x��$u����F�l'�l,�e& a��QMiH���!���(��o� v�OB����>�G^�ƨ:�>:�4��x�����{��]K-�P�貶~�����Hn^85Gfu���FxC�BL����:WH�h#s`�a[p@x�x�� Vf�V��)h�tP�6}�h���!bmjQ#K8e��pG�w�R�= ��j����su*�=b�$��!C�9�E�6�'|�m����p8uU��~����d�K��K��ó�՘k?v�j��)�lϖg⿖׋�����_8ь��U��@�|�y]�]g��u7*QR�տ��\���&� ہ�U���3s���3B�����^ڢ{U�m�u��0�O0��E����5����v�z�=F���H�&\���> A���۔戩�� ��t��T�zOf�"���M���k���bאdbg��}d�&�_�H�h����ayDQ��c/�j?����*s�|еO~�����-(䚼��u��B:����ȭ;������G;�q�*�h)B&�)�Ѱ!�J\��Buun���Ԣ"��I}z�m��\�6���ł�d~��Ҍ�:�)�LNCKD�Y�D����>�����`ʿ��p%��'d��L��uR���u$ܓ3�A��b-�
"^7T�Q<F;��5U���3_���Ga�C,0���D�?����Qš��*�	����)d�B��p�o�tԔk����N�� ^E�I2��Ũ���Yi�Uڠ�B�O��SY���s-QӺ�Sf�#!	�Y��0�ru|~v(#~\�4�;��R���bK���u$`�]��u�ͥ�9���䍓
����C��zHKZ2;��o�~&0�+��9r{'cm�]+>`� @J���N���Ԓ�'��r�ꓪ[q>D*(�9լH_)vc�W������{))&�v��8f�`��ۿ`؏�����3�{EI<5�f�.c���;áo���p����+�+���S_@%ĨL��� 9:�3���T��8�/���y��M����W~!��V�b��m�@G�*�x�2� =�)BL����fܖ��IVZfr����<�;�:\�c.�W�0|��%̌���1�-����?bᑐ��QK�On��r+R�EjA����p�|v0�q��B��~�Aٚ\�N$��,�XR �ֽ�����G��9i#���J�P��T��&�{�$1ώa�������u��g�Σw{G*��V��<ƺ��G�gc�U~�^Qaǰ�������I�R1�����*a��@0��#�`�o�;g�'�f�Bm��e��eM�	�oՉR���k$��"��G���]���UR53�WV�'W�[5��Q�=����d�l��s�O�Z[;X�$�B��2�"�	��VU�,އL��M >w��$3���!���&��Ә�S%��������/�(tGBB��{<��j)��U� .�x� W��v����d1�S�����3���Z���3��K�i����GQ���Z�_^�E��Lݜ�&{o!��i�fz�=��Q)�E��H�n�4:ДA��\W��G(��B�`�w8���;�.'lߗV�R*�(�mQ�5�g�VW�����GH���O������d��&rC�ف�c����M�3<��W����߳Vho�C$C��,��{��l��t[*��3���2ڒ{V���g�	3�J4�����(XH}f�zBvN�L]����W����UUkh�-(�������]()��\-�W�np��<?x�Q��o[?j6��Bb�����ʿ�F/��.�d][S�}��Jϓ6z2����H����}�|l��O��I��Y�W�_D0��ї�p�e�UE&\��G�*�?���Fa�2��TUs�9$�A���#�ڷ���3�{��W����Ō`U�����z�Y�?���1�7��z�bW��9?�Ȩ�Z���k/�G�rE��ߘ��kv<���V�ݞv�|������jӮ8c��7eI��qjT��eڴ�t��<1+���̫z,EJ+J�Th3p+� hSu�̹��"�M��Oȹ���V����k���	v�|���%�#�=�<��p�t^L+V��F2ߡZܬ[�G������pL�H�|��y�Z��	�(�7Éh/��8���N$�� y�B�+r ��ٱRh��s��r�j�p�T� |Mu� ��x&�|���Lb��B�	���<�I�*:��Nr饽�U��t���ƗW��K%�f�+^�[&��u�Ͻ�gD�
Ċ�I�uO�<ؿ{�t���ނѕ1ݎ a��B&��3_�DF��F���C�,	��ZЌ9o��+7�4V8�*�Tߍ�u%KY�&�؎M�g�`�rGO�ı́꒽��@�'X��O�YR�ˣ��f��8@@��\k���@s<1�/����L��F���F�56uq�.�{s����h��f�#,J���p9�/#'ȉҏ��GE<��$����I�;K���K�)��%��v��ҩ8�`b=��yyr��[q��	~ >p�QW�i�賋�:H�z��]��DR�e֖p����rsu>ߐd	�"Vں,���_��hJt�����^3Z{���+G�F�n�#��Yʦ��H�j �'J�� ���(�b�����p3�_x���S}7h�sf�&:ϲɓP'�*!& �!r�/�;K���ԆǍH�ҙ���)!�����X��Md���U�n�z��݃ږ��L�|)|�^
���l3Y�6ʑV�7VjH�,5u�K���9��F���qaVhH�+¹�cS�Kc'���6�}�w���]l���7�k�nf�gL��0b5�R��DE��f{ �V*J�\9F:(���^�i��ȰIQ���cC.��A�B$�3Z8��Fa�G��c01{���@łL�T��	ƚ�m��?ϰo�?�����rd�6B�6KM v���v˕�����~k�H}r�_l�ͧ�, ���G��Gn��?}�;��D-�N�-3�5��~�ꇏ�OX�7M5�փ�g�6��Ra��h�۶X��x���߬���%K�9���VA+Rj��ł�(;.T�P^J c��M1�$�g���?ۑ��\d�K3d��V�ܞ.ޖL'�c%�a����.]�#l��k9
���\��������f� ��x���	����i�fA
��w<��5.�R��7X�;���m�j��,�ΙO��rK5��	ch�F��,���� {���]{���x�1_���]$@�e�%�����#T��)�IA��+�ͥO���N��oe�b{�jm�Eم��'@�F^�H����	�l0^ٝ��Ӗ!Ɲ�V3֮�������^	��ё*�=�N�[����� ��Zufia��X�8	y2nD��~���,H5�Sb_u3̀��m�/Y�Ak�Q�uad�f�Ha�o�	�
�#힔 �l�-���8`�K��$?��!ͦEe�y/ܕCes�s��4$=<����9:������ݻ�q )|O�Vz7+��u��S=X�R"dq(޹�a�d��|o�,���?D
��$t�C�i--�&�n�0�4,"hlص �P�U��S3��.�P�\ª����̲ু��	��#?�i6�����a[�sM~��j��6��Q����ƭ��xb�1��C�?�4+9��`�?�@�-���ڟ8 �W[�`r�xV�	9I�b�ʜ	HW����xј62�!�K��cм4c骄�ޗ�V@����O��]�ѭ7�d鶟������:d�;����K�Q�Vi���"����pƟ�cL�s[�(m�l7NN���lX��*�dr%&����B����~��������E$I��ľ��Rc��%
�J~��-��׎�	��[�f(1W��I���P���lE�����*�b���p p^K�Nt�A�~���&`���Y'�\ʔ��L�&�5P�d
����#/s~�9�vܪ�/V���v�Ռ�yv7�f�(�����0@�z���t{~h�)`���S��〈Ȕ>�'Eؠ��aI[�������k_��@8��+F�^B��'�\��0�������c�x��I�<�;GŌ3����ǎ�د�c�K�1,��h�(�ď��q=s�7�T �R=��L.�O��j	�,��Z��oN\8��ӊѠ�@1�w���?4�s02JwW�~�G�\l,F�O���"�`��(�v�\a����@��#S�꧹���Vm�\��E� %ߠ��X��;��VA��~j�<7.
���m;?�g�d0`Vs��}������|i������n�#`�F2�2�83��"�q����y��ZSr���O�+tPb��z3��nUz#����xW՛y���>��J\����?�/&��mPiݱ㛔U@��Rz�	pX0n������Ap�0e|]h��~���?���l4T�p�Oo��n�R�+F,��c{��������x�L&�������c*�������U��G.�<��y��zR*���fIC��9�[�{����\p�f	��;5k	_��V�$ɗ��/�φ�1d}f[� ��??�m;I�p�w���vJ6X)�ˆ>	�<�hkt��Ȭ��>��5@�_P��.0Ƌ�h'��8���MC �
�?$Ho=$tCO�/]���Jx�#=/'�x�Y��A2$�_�&�2�I�%dېu"~Ep+C���0;M���ʏ��Fb�h��zb[�4q��{}0=ռn��f�M��ҏh(�t+ݗ'Hn=g<g.�	��X��<=�#J7X".�v<���@�dCbe�R?�WPj����ɬ�F5�'X�1��7|L��k6�4��f�,0܌E��Zʱ�Fs#AH���ՄW��uI���&[�(3H��8*�\�K��$�c�}��FA-H�c�B�Q䪁Jkh��zT�x;�N�!͊������^���]���6�R�`�P���Di�w�����J�|���!�V8�DH~�H$Z�þ:�� \:s����q�d4��$�z��c�0����T(f=��Mw�nꉘ������r�:^�2.�p<�?P�P1;�(;g�Z��X�t]���hrJ���,TώxH#�:���cq�$� v�C�:�OO�q��`�+m��.�>�o{>0���]�#K�͓�C��r�?��QRs:6���oa�����9"��*1"���P�v�ְ���8�[,e�tI�m+˾'� �lӌ�O���b:)]f�@߆�P��N��4ˎ�X�!���u��#:�0�3V���N�9�b3�t���M=�^�>��j�����eݎr&8�󵚥���a����fu�r:��w߾.*%'�\�x�3���K����m�T��T�2+��@V������zz�[6�����Q���+H�i�ӷ`�:Jɪ=*�&<�>f����0d��2����{�i��98=!�����N��w R�aN<��UQ�~�2O�K�K40ʷ���aS�*%+�F�J>�k�"7����a��� |��6����f�YGS�[:�d��$<�=��Z>�N?��`�D�ߙ>�S�� a�R}���p��z�'q��Ν]G0�n��J�����TQ� b|�c�-��0E�����Ǆ�sh	�n��m��r��fQ����fF�-�w����KwO�?�远�z���	�pm��R���l9
��QX��^.������=~4�������C���?���r�'5����I��W��+�=�!zK��Q��&����0�@��F���څ�V�z�b��x���v��
,�� m�]�� ���1�T�)�P�'#���,>��I^�t�J�;}��9*�2�ӓ5{{�*0��,[l��S�YD��5ͭc���"��3���b�-�T%S�*C~��b��Lo��`��J��B�Y�$�!|P.\P(D8�5*]�a^��H.,�3G��s(�C"������{m��U����J���������hh�9�o��"�a�^���ᐟv�J�^�ۍ�@�P���H��jXI[��n�K5�tj����Yb�}2�,�1� $��#�=�7�Z�Fz�9ֈ.��΁��J�8[-��z�a=ۜXn��8yȝRs��h���Z����ul��5t�>�苽PFhuё�
�9�Y�S�^e���§��Y�E��s�xV��P��w�q/��?�����:4p��iN��� ��QMY��/�0��~Z�Ez����GRS���g(��40��	�G�e����0%l�X����|����e�|a��N�آah���BSl@��d�]��7%�ψ3�:�����F�'|��},І�2t�}�{�a���+��__��oH�X��N�Ƿ�Ŧ���N4���]�P��w �����;@����Lߓ��ZZ�`�%�z����-4vR�[=��'�H(��!$�����C����v�aJU�s+`f��a�K>9^o: i���ͨyd�T��:�0Ւ�s�,���^������%D�DA��%�e��!-���sO?��x(����ǈ�{ݯP�J�~N#PD��$�gΔ�2��F)�}����iy��2�p��5m̙4�E��*���yl�.�]�J<�JwE�Vf��7��A(�d�v��5g��'B���Ź�̀��2��p*�O�F��1�IPȸQU�a�>��}�Y�kn}�M+n��Hm{�f�K��-��	`�Xbut|�gT15��r$���,��x���\�Mc��T�g�E�Է��M���?�k'�C�m���wዲ���<U�Wa���LF$���:�:K��u ��5�ws���b%,=�w�P�ٕ7���ޱU�~0�1���[��eϽ�P�4oq��.%�s��etWnj�NT'�щj�3�<���ù�n������Q6���F���q��2����[\��[��{���j�le���D(5��At�t�����'��iҏ�*q�v^lF��p��ˮ���OԢ��R�6�6�)�6p���#O�����oHe���3���[Vc�`�^�(k(�wH�\�s��{�CTS�rK�O�K���!��T.��=�3 ���84��e��A7"�)=r��+��`�Tk�w�I9(���AW걱�D�ǏV ���eVB�W�K��.� |�m�>��
��+�-+KF���XKۋ�/��Bx^�}��e�/�Y �&Ƅd��v�/�Tn�mu��J�cǚ��T�l�7k�D!w�y�(�P��em>Uk�}��(�'��x�3��.��Yq�x��!x�U�4I_�-��C�cj���VT-\�=���*��G-�
jʘsf�}o��QL~���+ z�0�Iͽ<ԋh T���R��,� ��T@�Qg@Jr�E&��d�-�prN�T�����K0�2��x��V�zz�$t�U�+�	t�R�d���::xe�e�d�kʸ�?�y��dx���'���Zi��ÎA��FB��g����A���0�H�8���h���L�b}��xg�2 �Z�m����(?�_"���RĽv��>zr���Mm�B8�>�\jif�`��`���VW���~{��#����]����C}����Qu/���u������U)y�/)���)9Y]r�ֿ5U?	s��Cד����pK�Š��e>�t�pSឨ@'�2n-+)���nޓ\a'OF���w���𯶲����(6�B����O�c�i�P։�z�18�#�R��l�3^"�ш��P��#^�w��叞A�=�J҄rY��u��c���Oc��3�b6�ƱNC���"`"&D�r	����%�4�t￥O{���؃%�n7�	)�0��Q)"�����fj9���-��4���,���D*?�G:�7؁A�0���'p����3,�5!�$As�^��q,vtxt���*Z��l�x�Y�����THtӨ��B�X�Np��!/�^&$~G��['�� r�����i��qf��!{O~���V�[�2\�I�i���Mvy���� �U��5|i�l��|�wm��)�K%1!~�1���4�:%�&�X%��m~J���c�c����@ɕ�� �/Na�Ћma������%���څ3�כ���Z��%�k"�w|�h4q|cL9S߭JZ�m�������@��,!��3s�D�d���f1��ϩ8g�
Ru��S�q�K&���+A�I�[Pyi疉�<���tv!��q[��a]z�43M�}�Oa��dc���Jf�]�7N�7��8�1��(�z���������,�vHRi�x~] �eh��"c�s&�SY���,x�4��$à���C�*������1;W��f�@��Yy�ޓBW��AX��Թu@͖oӥ͒	��b�=J��<���*��,�uZ�{�'a��R(!�w�����ʡ?�z�A�f�ٻ����w"��Y�}������R,>BA;p���,�ħ�\P����r�ʐ��O �%�%�Ѝ^�N��e�5FM�Z_h��0e`E�f�uY@����$�a�����|*_|���u7�����Q]$�T=,02�U8���f'zH ���a����;1����n��.��ϝ&
�"vg?�˪Ќ��g�茤֥͎�N�T�y5d#Yw�\9V}���k3��S������{�&7�\���C�f��E�@YIH� �Y�C����w�	 A/����y��+�s?���<�9,�W-���6�1���7$x��~�IuO\Bx8	�0Bk$�e����ǆ>�����٥�V�����Q�e��a��y^����[�(q��E&��MK�|�G��|������ز�O�	���Ri�N�%�2zD�� �A����lE�͠�X~�%՟������E�j�WrEa���wC�z�q}�gop�Tn�ʲ�g!:ג��=�S⛁3޽��hG+W7�g���IHtV��]x�$�4��vf�t�wiᢸ��^������Z�̸�M�F\ؐ �4�&��~�3��?NSS���	4j��9Lf=7��wa�,c+��?��iJ���{R����߯�#;"T���񘔿-����`"���q(+��=^��R���"�n?vP�B��2�x�����4M�b�=��6���Z�lH͖"t�1S|U��6t��@��v6�2�6u0����
�o��tR��xs!F+\:~�Qb��?���@�:�NS����\,3�#��gA����h!m\k��<X��K�D��2G��8��ϴWp�N�E���8U/���$7��j�܉�,�G�h���b;x/g��b+X��;�D�un�Ulb����t�b�NW��zWphrJ�&�O���E/��2H4w��W���"mn�ʉ��ɩϣN���'�M�.�VdvJ�~5��b�Ś���	�ܝ�f'R�TvR�%�xZ�-2����S��L�Ԉʃ�ѵ�\���j�&amP��0U1HӲ���"=Wc��3��Nǒ5�R�Q˕�a�ĂT�ŷ��հX&x��L�ʹ��1�ϸ��L!�]%�DTZL�lU�ߚ&T�d�if�7�x�;u�1G^yߜD!X���R?I