// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:50 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N0AnmtlMKLg+5CTc3XfwpSB9ze95bkpAqZqDa0f6GbasZi6Y23rsBlrrqrL6YwOO
2SuKzaANMcKBOs3j5youx6RSp/Pt0BCp7wrV5tXkcO/ofX0/qZxJyw4qCWQilLML
8YztlCh4XNcxa/OmQHDN+eD5SeDxzVJys7coJseeO1w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6144)
6jgMRil42vhZ5YGAo5wVCry2bRJuR7wPjNVNOCNLewftR/jLuHxKTA73olZ4b1Xu
bPr14RKrPuM0jxshG2T+X1VDsf8WtvC1wvduZHswORSpqyEXGi9yJ1yDh4uYSB65
oYzAszt8GYMjMivDkyRzJHqEr71J8q8QehHi+8gAkM/U3pXFAA96lfoqn8bn5NCZ
RaUQMHqzCnU+eCbYz8oJcWiCpbzEcH/C5lAWEAUYSdgd3U01yFmcxK4SrvDQ6v+i
KBamkXBXzajiWh6l8HaiPkfNQ5LpQAtB8cUnP530j4IFGyVFWi+wPJ3BS13vYrVY
9qWYqFFTeqDc45UsXCJyJeqv0Zh3+3dwyoFPnACCno1Bag6cfVxfmZns7qp3pLu5
0A5uH6PYUdAFMfn6uJzyLIC7dLy8NaGj3OxLmKNdxcXP7jj/jvNxpoDcGuQuhQ2T
JZsxJ7PLfEnYjRY60D/tCLMHAjJbxvYmgH2HYL70bMRd+BNZI9QeXewvg4IAyDeC
DBVsV+UfDn2C1XRG3faxDHpzn9gIqWZGFwKXguosFVDtcD8PzXlPEGLwhcawC6b0
W0ovKmgsoxLzXPU2WMwrG3wuYdvr9j0jYBaIMnPixoWac/nuRVB/3Dh725UAQlOH
eIcKLKEtnbJDomAXREksOTlPS4To8SPzqMD69zG11TRe9K/ZfGmVUu8Tsk2HwajU
d2bnhECT8JarHeuudzRFZLj8lUB4lpkYFW0p/7eSf4TDHwBycmWhSy+Lw0g/3oaf
ZoAd3IL/Wsusuu1IrlQxScPIIXQfJalIDGBVbwbcdnLvAhRyuFnWuPVvIplxyfla
wAVPM3mtUVLIzFSiwNue4SWMVkSrPmkyol2unAr4FMwn0gMj4iFbnE58gVcTA5hv
fJCb2qp1grpXf/d1wF+89CreJaUwQxH4Nmg8qsYER4ehRDQ3jMWaZDkAe6p6vwH6
RNkqRa+nAT0rqz80ebEWZpacDuzv/Lr40kuFZcWtaR9zM88IswvUidtpH8ZwYm6a
8lYs5kq1DzvhqGwLZ1Ym+RvQ1QbtL18mWhOZtizucNpFxI26znvx6qOHl/GziW+Q
W7YS8Cslm1mkmq2fDsgkb7oM/n/DKrgZOVGKMR5ryz3dk2WoEZCysKpts6H+H2PG
dtu+hTsmefyiPGHarm8HPrMk4pSRCX3EQ0WxogEeuYv03rFSN6ZckH7EnAREBUnl
eZmlpdNkGxrGrylhMwrZf0v/2tK7jYUR/ZuFPF9jlR7VvhNqK27hNt7TRTdu4dBU
ZXx8JP6VngaW4aktIPDuyQiz9PLChZNsE4UNTGU1bLyHg/mcMr8Kxcc400dNJ7av
LEtcctPHcKfNu5rwDirn1ZVCmzna5Ga6cW54idzSUh1rx3d0ERv7oMY9QfH+ji4K
AUpPk/LJUos4ikgxK6PlEbGw2h9+FqyfXYAdwLXL+RkUfRBQjejLxgt5HlKUxaH/
X0QYwDe/TStb8pYvFC4iigdyqwRVl9A8xyFPh+9M7i9gxcgBVrocw5NYeMcagBHn
YnIO0pZwWGP6DJNnDAfG4dS3k+73C45/90tC/Rf/HicgKMcjXPDE/LAtL0ddF7FI
BGwthZr3xAE5NWDALak4xFHk2mnAUGfQh2euTcylBmD6/sabVcoKrgwE6Qe67vwu
veLnU4TnQEAgkmQNAkWQxXMyaxVIDo19ZDruP3AnuzQyJdQkZk+2FynnJEGM3iPv
jAERPl5hC4liNp8RUPX8U0VL1UWoYKJspINlw3A6ZcSFUFcdOkPgm9IbLSYEQ6TQ
0FJeLvo5LGp7fiqdfPIotmkoC1gCoX2yLuFPBYlBFgT5fuVVNMFhmAC7sJ/gtSFY
M/02nBSFfzXL1XC0wCdAXShJBHrHZQA2Q2sNE6+aWGZf1NVGF+ONAv9kJbxL0bjU
ZVAiubYAODF5kli+b9u1gRyfY+j7595JjjjxECxLlG4yHfyGqOQQ9Y2ujMVtnBQA
xw7QX+rHuXmzSXhp8TttvITznFxWjWi54PRJQBL0DovsA+ovSVOB3CZKxOqLXLZa
LWhbkVKDY9GhxYVUAm7CBkHzzrsj/KJEEZpYPKbxuP+8iSrYdPgcWIXQ+xsY9/rn
3qkGjXv92eT+JbnlsuuzFk8Onxk5Ow5jPcPFM3y6uuzjuO2n9tfTttTG8lSC3rLy
XhDnLubcGyPrd4cCuZKbSZAQaqK3ypsqOkqOfRLIXgcsOhVmBe50VQwHE0tXK6nb
A493NBQeppCPIN4pPQkVOZs76sP1v8uyOsJfOXO7w6mkaUawNK2Fjk0N0qyJknVM
9yj6eU3LvxOG1ua5h5jmx9W6aslTj+0YHYChhl1t++MeKRyzmCrW/y6SZMnbZ/h9
NZzCSKXNpBKiYyAfkcoQesk4f5A1Jk14yqCbASR5dgLbG1SXFP6/kjydqDCANGw0
GnkLIzsT23qeiPyfao/sOSiy/C0RbQJAQ+JiuvngEk8Q/y4rMOR3ub3PoTn0tO59
dWIgZZVfQ5U0sizej50fiXHK9o2dQy3VB+LyleO3lu4/ha+tLNiMdYlG74sox+V0
+iINnuWbegHivfXrloaKPvVaSQQifk2qcuNstcLN8ErBUcRblqom/DqhbvJxTzNj
2PNVDFVv6yO6P1uUf9vFkYdXds9SkKReQhOFv9DLaCUqu6+eGID12C3N2hN41F0D
bPMyrZ1s7gplyUaKxu6BnBUB9ryaeQfu9o882JRWBKT/bO72Hw71PduOtqINC1cQ
2q4yowdYHcJVF2w70uYup6s/5RiGRQCdeMVEIKLtwgRaO5cTMMwbXPmUnS6VmgXc
iRx2FH2ca0gRNr/9D87DbjXTP8IKzoa5CURAyHTg5vSoFkFmfEq0jH+tR8qADvan
ZmLxG+kVkT6U3mxX2X34XHJORjTvi0rxxz5LO0Nqma09wTh4oAMKG0zbw9wJla5X
yR7J2B00nmhgt/tWUIxx+cSr5QN9JkuiLe5a2KFWcxUEdQd8OwxSsnQEedAOSZ0e
SGslKR5KIYq3oAJAIo7LInz8R4z8Gq3eJlWGD5NivhIUZgr9ImXL2QY8m3DmFbHM
I6rugQbrrnps7YJM0BpPWoQXfe5gPMvZTCiiR6Q5apQDofQKJTqCzKvi9GmkO5u7
RLPuVJgV3qBxxY770rtyp+3k/fNkeHVjsjFttRvoul3t98w95IQJEsXNyOieEJmv
pDcNycHh3oqGGdG29h7q15LVtxFuW0wzjIJLttbMnPY6Z0UvSO9G+kvbU6Gl1OOS
j6Ic6kLPwTmwXckq2a4xPvqM8yPKAE+ocGCbYaf2p9GpiVouvE2ZiWktaNV2EGew
y75nW+hcgwBfLzSm2CvWZmWgR3djSgPYMp5eJdAtEXudhFnn2gY7E0iPIsAd7am3
Fvg60/yCJCj3RTnAEtmHuMsEyraGxh20A1Lf4p6nKEy2YDY+r0WMaMsuF16hqjID
y3mnxirh3SxphogRlC/PFj3le9EbKRCc5aBkGkYhHfo1QOVqY3KgQQ4+tMKQULHW
L0lCu1UhZirzlxi45MqnVX2En6oRhTDliTLPLsaPgGz6hEAecL3v+Rxb81PqnB28
vFnlbZ2uj4aPoIjOMK5T6RPXVQz/1aZkIXn8SY9L4AHTzICMK2BD/QDwH4lOxUJh
K30UpcG4/EGDq9VIU7vIRCt/UAgXzIEF+EthAEwSa2uEDpj6SLiDBLGIx2BnrQ2r
ZPjViP3t+kdAmPinDhnq/GwTZ+1DoBkrrlXtTHG+WLZEzRY2BZbKQyHvFsjqU5Cr
XBaqRt+EO96HFgRPt6PUcUucrQJYvx6f+BzI1Hb4uJ659gaX18MvoqtOqagIpR9P
bJhCpMaxGME5NxE2lgCDNTenXExNHMoAQSlxk3Kole8ODUOWdwyvkc7dZBLo4FlS
mQ8JWcAoWwBzJlOKpmeBLyJlTmuvLcFhdxbLi/t4xIZPIGmTGzr1rA8hcmyYLRt2
EabpxMu1TYJj3ftdBWZse9VcfV2Bc889/pfHyDnZ5abBLUEGP6h3W3JLgrEjpxAf
Y3It/nY8pWPsluvGFJAM1xJWsYMOr54wMbXTitJPRbnQsrH3o3UakRymh5G1EzGB
RfsjapqgnTliFjlX82flhTCKk9iBs2FRowL69heL1hkjnF/eiSg/QT8U0dX11hQP
SEmYEhvc3Xt+EB/cwwLDRCZe8RdSy9WeHcXRy6GLiFqLeN4755EfV8kIYipy1Adc
nxMlq6U8BeN7Dh9tIXizNdhKFcwV20gDWbsJWF0gz2sM48Ua4v8HdwBftLSD8AON
XQdGXFdfCW8GQ017Jmhgc89BPL0mb8kUYhDsrGa5jPFi6e4Xya3sKWHUUgLVWNtN
StJhC+uPXna+ckhBncKBniSaWE+S6plIF7ggFjLEamMk1D2bl/fjNyOqSbpQsPuf
1bf6A8mEyYEc5GSw3EwYlcguJQxxqSvqMVPiKs8G+KlW9PdpjZ9YB07W/cz8dcwz
WNLtvUiFMsruLwN2x4YV/zINBlV6rTK3x22ZG1G6PMhseXIMBy7ZqM2p/hnlvSTo
5EsZ5ziFf40ggaKzNy2dDW0BuU5ITs7eRRz7EMMobau+5raZxkqqXny73uI5gEdl
TwOuhr95Ua4CFZR3btvBnzMaiWF0JH7PHYMtXLC+T3KQp6t1L9fQB+kObqpf6jWY
8IuHoZ5RTxegXPcb2bnQxSd9Z0D29P1wISmUR2Y/RQ77PYf9AmPAylhUppKnlL+D
FLmsi7quaXZgmh6Ix2pcYPGkh53oiudoXO3yJbyl37Uw/5L2ICI52zzykA1UXPJS
scCWWviitF3YO9uQdMJwTc96N50yXK955RXrFBzPW6MZfM/Q3KZBIvy6IdlktB/T
j9wC7MLFDvyzZJ9vrsAl2TkT2w5cpC67ZTxBVNxDT+jp81gyuTC0ltbNYBhCV4wB
G2R/a4qSDpF15bdd8bEstVMVvhuVyv8FnCD2F7JvG0o9BMy39LZZzeZMGfA0oYix
gS9lsDO4UeYcz2IrDAVN+HVxbCPvLu8m1NCRik/CGdpjMz5RJGp4my3dilC4Ssfe
S24Y4BUim2bzvK9td24o4+Yy/qMiWUmpkJUWiOLZ7uDyE9YvlIb9iPXRp5mXnEHh
ZI/D3LIRaOjNFHa1Fj3corRuZUqvao+E0cqutflLKeuSWyEFVOXnDEjRxn1E018J
WgNt9OiY7ec9AgUKF2bCjXb5nazEe/6TA9oJ3vbvNtieLYFWQVYveqAmv6Egxbkh
KFVq9N24fYveX+uu2dsiKg9jDa2M8iqJVbaz2Oo/bEog/UgI8l1qXvbUq+lfNlJP
Z5zZjJhN2b5+kBHXGT9gTiShxptPgqbSRX6w6GtL3jHZeQy2zn2TE7pCHFbSKOFE
/WsD2eOfF3vdzBrXhFJ9pWhN5SAuERs+lh5gmoEMX7SA1l2o5QrohdvfDNcNNa2+
7/N64NJqX8Itv1BLxdRekDnjOnXLIplfPle4d3h0uH/j+AjEMfJWJc1RrGFz8Vtk
8OYRgXlVGKOKhvqzKaK9SIDG+sSh21l9Fdn4Y1Pj4ubL1j6uWvOfknUgyqXbSM/a
DesT1QaixOnzcgeiOJfEBYiQKYN2JcoqaYvjMgKhUMIWYmb2knVe4BUl4iFfwrJP
p7FbX5F05ifGwqJU/j9LO3NpYYdpeyAiaNd1+OcLN9twBXdcuT4R0pOaNEvU+00A
bltW74/09tH3syaomUqQFuirhFdZIlw5dtzBT9zRozk7++eICRe2FMYg8nPQFmJF
6s0fQybGI/Lq98VMghiJ1z5raXs8DUE1cOELlw77elGRD5IZrJxOYe+Iv2I3Y/6E
zeHOaS+n9X2E8rI+vhwOD1Ba85XL9KNHRWP42lcWtrSNUwtvem/BVIbLpl35PUsu
SVpocqNTuJ3wT+yJjxGAcnRUo5mYBR6DS/dNYvAmBpdV7hF+GKwBIvI1jnxlqumI
B4Bdg169g+BRlZf3TZsx+5Sh0Qyhwt/V+nWU7HSzt3CvqkTuuH91P5qY35h+bcDR
QKBR2sIwx/ty/u/5YfjQZ+jpeA/xmcuV2+A9Sm6VIL33Lf5rWV4m7eZlS9YU/WJU
J/HVVpnkXFnMLZRMPKwe4jJHfKKzLKKascUfNkNZVQH8Z7MO7bzcbeQDyeFy8hwk
3tMX0nLaS/mVbcznONub9pPoh6gWbyLdw0L6Jbw8AJdveXdxNjWMF2QLAmCWIMnQ
u4310lHMLYfUeoTFP2lX/5XoL0ERaaLqDm9zEmCsjBADXaIL/Fs0keCwh/42X2x7
I7RcmVkWiEllu6PwWCBUmPqLJVSfkGFldNHznhifTwlHtNaVuuspCqLmi4BEJRD6
isqCyB5W/thERoNYvBusBdJjfo3k99iZ3QSzmCR5yqbnS/AtHUEJg88cmek09R4u
aFw6IvGDb048Rlc8+SJS/JlmvPqeIjvI/oGlukbM8SG5C3vKL5WvP/Efh4dzhW9O
ikfomBCDBl1ouAdNzZfsfGS/HmjdzdZVGD2JXykTQ5I8kBw7It1WGdsA8wODF5wN
KPP38Qqr9fV3cOA4EyB0AM2kN5x1Ru6kcmQpahoq2pCwnAje5wqPmsIPCdd0xz19
3AT8Fxnx5KyxiJ0B/110KqZErdd8wVShapkCqTbfWWaErAlAT7pVuY8IftgwwqiU
O0zE6d07Ef5Xs+3UafhQg/PaR+QMnbzuqI6UYPaFoNoayLW0b8uH1FmW0MEOZ/Ts
j8tk1uqAiCaFEx6S0qaANE5ZFlY9Ma7NYRpHCvE4Zf9ACwt9AZyhfL98Zop3L8RY
mHtAkaHtuklD+teom3mqaj6srdyqMH0Y3jxbQoseWv3e1ma2X70HOCydt8e+rvl2
b2Y877UZl9d3iE39OvPKBm1pQi/OfBhPh86Hv2H2DENP+7ANIlobhIuZeRRNsfCh
8H2uM3/b7pPUICRQ+AvuvjhwYNfcB4JPvfYMGLFgJlZvGLVvlZh87Ps5LUpKpPL0
UrIvPlGyq8LRDzvD7qoINROjigl4V/i4XH33EfoI8G6KqB9RgrChFAzdnhs0ZCGF
VcGXZLOT9vbgHv6js6ygekVpoR0BF9jJCEqpPMvv3fG5QIqrl8q+IL+PvW4w0jD5
6gS0yTNAVSb0SjCX7igUCKUMcLXeQZTsZl4Hoi8vWqaJkqGVnACyBaDm6hvstGNH
1ErYl9T7XDQCVN8fovbC2rHxfPqeDC3HRZ1b9D00CO5Te90qP320IIz1sjpnZ6xL
T0/QD+Kg1dmgLl3e9A3N+Mne43kWXRPS4xAvlGTstJWBsAM7is8rLBUxKA8UQD4d
J8JleUQBLZyOVQqz/igf1n5jYL6/c7SdPUIXESUj93N1/7izZEuwzCZwQiYI0Mhm
KjoUV7GnlWUyfLQ0dWKOxTrcNdQs0GGbhAi3em4ACkht3tS8tAuq7nL5cxy8QHZJ
H7zhYOdRVn9t9nib8iuZX/lNvnlwU37htZQ4mFQ2kPceITd1dL2aMr8Klh5Rf6TH
F4dOGe5zjr9hzvk10bipxt9kqE+cGCsJurS9md4BRT0GLqoocun6rdIVkS/olZ9c
Cn+eIfbtol2luP0pnxTf4fKGEQWzvtAXWqQEuYTYUfbZ5t39ECxemtpbaAKrfDr4
yY0m52HwlaJwMyrSSiibuyGigHaAOluCTUxOqeGSkbAEnTkHI7E06Y412CX1fVek
3L+rZNhQP/E3HUdzbdjagmlP71Lx1jI4ZPcjajvrkf1PHVk6Y8gqO963bSJRKz/n
VHsDJsZnxe3NSxxyaZtWYkrZsMKA3IWt87Bg/XIDRZkCJ5kipAzuc7ziNVDe2uwA
ziCHz2e9Oxmbg9Wg+WI+BZ2PvxnTo7/Omu96ZxoQgdkbYSnFzurh6WQjZmpIcj+Z
muyBZr2cPV/wyVMyhFm+EPGWTH+te0zTyzaOyiTa1/oyfGzJx0XeVDPKLPW4NdPI
jsENkB2w4JExAU8HoB7uO5lpkmeCliaqHOGAKfz1z0lBv5vEB8ZJWcqY2fXMD47t
EXACcoc4oRwu3+FIWxskJ/91Tm09zadgbbu2Zr2zA6T+NAW55/FIfqMgqm/iZm60
F79gNLBTlw1cysSMnyv2zMYkAoWD0jVsGMGQgFedtitHYJmKHTiDsMXVAePyk2C3
UPmip1zZJHc3WadRHmmRo2tI4bkAsrN19kPSWnUP8yeTDkOmmsQRcn9SyPsx4IS6
`pragma protect end_protected
