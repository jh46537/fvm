��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbʤR�,
���O� ����X�C�Scbe���\�} UR2���pSnܒ�%i<�xY8י�#%L��f�ў��Q�����g2��ug�ƞr:h�"�FʞK�?��K΁�ٱ�[�'��\��K�q*Y�J�=��ը ��9,�:_�RC�L�%�i�~��CLM2B�*�(0H���S�u�bS�K?��y���fq�U�d��p�I���ɹ��Huˤ�g�;�^i�g�=v'f���B�=⦯��B���컱̲7��]�__�0p]����O�E�P�8)����`�9<�6�q�� :/*2����m�b4X�P�h��[{ɪ3�����`U�Ŧ�U3�UH%D�`�m�p�A/Vm��>昩�X�i�G��_��oU�����XB�(�������i�('V/����$��j�3��#�Ua?@lF��6��5��(/'��]���������Md�j5�h` g���j�L������;v�醈�#|^��tC�@��g�'�����:eǅ0�M-���'--�k!Vn������O�;�4��k��1�12�`���6�#D�s=�G9V�t]������^*��>��	;j��⻲@5���a]�шM\�Hh<&�S�3��+�<�f�!�
�C �ѩ�3�஑Y�Qn�*�=�%�V��QD5�vU��Шd�}=65Z���k=미�+O��GW����aX��5M�d�� ��W<>i�q�AsK�N���-U�睸l墉T̷9"NHk#_����qSnaJ �tql�;��I�}���1�R��-R����9�u�E�H�����Z��;)�,ikH�i#�7�c��
w���cG�:7�&���"��n?�'�œ����H�-|����K�xk5·GS5��-f���.]��wݹ*��=.w���Ŋ`<\3���^���D�©dW\������f���d��ìbL&A9����5S�XQ5��1>��ˢ��
8�֢���#��@�si��>?L#�8aD�;�U-}�)�.����$,���wisF���kJ9 �;��q�p�����$���"�A��Ń��p�L���k��>Ǆ�C�ߧ�Q�]%�S:�>��E�X��\�;5�e�����������t�����[N�WY� ���#WQ�8}�a=>,D0�%�`Jz��������;���π����|�"Pt�d�3��BMi���s� $i���pK�))	5H�ø�W'�}�"��}&����^�
�3Q�M:&~��^�:��ծB<�8���V�㮈ӵG�%R����T+�^�0e��t}�;�X���"AN`<�ުX�����[u�<�6�x9YlY9��-��i��F�oHh�+00/$[�F���A��6�'|��d��Eo�(vdcz��\O�\��*_A
�d���(]n%!O��d�%�N={��|	BS�~�H���x��^�Q��״]����zv���9��ln�l���F��[�]/ ?�Y����6�F#*ׇ:?+�C��/i�a�M��U���A��k��W�R�s�� V{y�2�9MrV
T�0��'Rx��}��c��\PBl��+��c�������u):|W��c<x�D�$ʮxp&��<�p��Tӏ-S���?���9j%}�睚,���}����I����q�"��X3��f�j�k�%&�������"h'P��|q�:Ť�3zE��^g�w@V�т�NJ�ux5��o!G�"zB�k�W�[�±�)��٧km�{Ս͍��TB��o��
χ��`�*�6��5d��S!gl�����~��C뺑1Ld�����ó��˵d�?���Cq��d¹�#��;$A���6)Mg�gD�m> �-hY�����aBj�>����|Q͖Չo�trX���(2������mer���e;�]�*�\���8Z�t!ч�	PR~$�䟽�4���d��N|+�.�����h#���8ő�2Cב|T&x��T_�s�n�pP��A��x1� �@_u1��LI������q�g,y�G\^�!&���'�t.�q����u���I�-�='�+�oRToʳ��ӞH呒?�!��l��,�2;���d��i�eβ#<կ7����.N	R\�$���Jշ	����]��#�.�#�#�^�a.��G����@v��wh��.���{�-<Kwn�
o��4t|:�l��k�P%�>��%�.9�N0��`uU��_��������]e�&^wh�e�ɳ�(��@�{٥�ʹ	�)�d�-����t�:�`��x�����u��P�6�v�3S�ϺƲ�ۓ���=yU�oş�g:Q#$6˲iJ�WӉ�A6	����ܦ���"��ۨ5Э��(���/B�wКY��Qx��)!��$��\׶`,O��B�Jl��e��ti�j�`W=cUo�����=�����#��Ǳ�lֺ���,&(��u� ��8�;%�QZ����Oo����j��
KΤ��3��al���x�t���~��1�p)���Tn��E�FzB�l8--4X囥s}V$�����F���][�1pl�U+��-��	%KQ�d����\c��>��?�Q�%V4ƻ�h�)Q�Ɛ��(�=�@/hg*Ϲ�S�ZH"+����\�1�-0���B�i^I8��^� ����U�J7J� :���Y�k�dp^��VQh�M��Uш)�F��,61A�R)8�z�߁X�v[�\�5he�EXD��;��Q��>���.�r�FS�$`zm%���H᠄�J�P���Z��M��9�/���������!+�P��6�N��
0XK�/rY=(�����v�����1�1
ߊ3̡���m����P���W`������5xW�Ȇ�%��:��n󉙺�ˬ�@F8�Fn�5]�d���@r�U��F�M�i��0j�;����y%.�h��P� �_��9,�E.�03pW�&nX�c�E'ek�v{M����gA�Z>�����R�h#��k�T-K�q�w��i�E�q�ʫEk=�5p,����m@!B7ޛ~In ?⥟�GFp���N�R�)�.a@�U���_��0�2� u���U�v�e��f俄Nݽ��/M!:�Y|,���lPhՍT�Sf6�����ĉ�s��9���.˴�\�٬�z����)���l�X?T�u�95�W�����5W�.��X�Zţ��g�t,㹆s��HAkf/t�s^�R֨��ߍ����y�U$撅���Z���V���j���c��`W����oh�~doH�=g`7�,6���4���;�����g������>�[P��NV�[�	���M�c�I��ɵW(@z器ܱ�����3��[d�H��tSg%'~/gʙ�U��O�D��,���H��ݦM��Lǜ�f�T�P0mL$�ĺ�����;��m�<[����~� �ki�/%)���@��54f�E�R�����-����E�����<[
��-g�CBcL-�~Q�%͠�d���H�EHNs�^���f�XEp�Fxc�?�=m��u�8n��r���A쬻�d��o����{B�����}Ta.�Ƕc�;��`0"$��k0�4�����lx�I��C�W
`�6,�(ڡ߶�3�����I��fI4]��̿��6��!�@0g>�eߪJ
��F~� MCS�o���/��Xi�q̺,�t��M��ܳ/���VE�$�!�!ى"���G��}� Z*�<B�p��4��kTN_��@�a�Z0�"��F����\��R�ؔ�⯛�P:�j���jIW��T�G����6yܾ�aΞ�-�Ĭ���N��j`=e7@)_���4�i�?;�bi<R��L�;h�f�'�}�����ڜo�LJ��5���]6�H���WgS'�.���u0���B�͐-��M�����v�`Zz�����vt�xm���N��)G�ʨBD\�Wv�DK��v��:v��	�D|�OQ�Ɍ����Mxd��� zA"����s��;4��y�P�e�.^Q�$�"�˫s�73�B�|CxI�qGw c�Q�]�\�||��I0�ZjS6�%2ZJ�ąl�����R���V�Pt���"y� �KR���_i����\�����[�m6-z開��N����g���\�e��'n�?�+�c>��Nw���m����8@��?s�{��� o*7t	d�{u^���<�Q���A`{s<�硸�d�H�	��K��*�O�$4�j�-a��LP�c%U�^l�H?�\���%�.K=�[����H�LH�PBG�_�gi��Y���")S@�r�	�IE�d�h�k�4����`�������+��}���RX"���N�.4�_�X���*�)%��M^|}G�Whɡ]�x(����r�cx�c (���9�s�!��ȗ�'r_w?3��KP�XY
�l� ���)M1�әά>�V�2C|���p�o��n�����U�_m�c+�G]^�_Y��۞�_7F��~-Y��0іU�{C���R�U�0��g(6C=�в▵^��K�ϊt���|�F�MU��bC�vX�}3yK�Č��wI�\�����+�\��?3��,*HcO��ë��mP9���zp�n�H�ڊ�+�����H �j�TVr8���*�ͳ�x�A�&���@�����s�H�s��/�����BR������n�_���Q���'��!���L�^ X��Ĺ���M�Y�_n[%T �/gT �Wy_��:?�8�6D����l��K��~�2�9���*��B���rQ�Q�_�cN$@|�u4���S.0�t�S)h
�|�4-�Q�]N.=�]�����?�咤[�:ԧd>��*/pQ�l�o� *�.���+����� V�D�׳���:��V����z�Hs��eڗ�O/�,��NN��M%>$���Q�g��K.=9���`��z�c��S }|b�, �@~�)JYW��O����7�׽�d� ;����+�=<���W��i�&D���K��
/����@���(Y�&ʮ�a4��F R��O�ȉ�'X(Y�>�h?ǘ4kA�/�o�G�:�{����Z�d�ֹ7��{"Z�-���-w�gA~N�����1GӺ�f"3��������u|�X��d��t�L�{IM퍕ׯ��j=�!�= ��n����j�V���Q�@�S���G#�u������V��)��:����]�#v��|皲�y��Mp�c3	ִ�7��Ȏ������q�*,��o'rE�����(p��~$ ���~��#~��o/dyV���<�j��