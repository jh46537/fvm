// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:07 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ihXcIbh6Oti52zE9rm6+0DwVi8hzR+BiCaiG8s+r4HDf/OFvEUFO7ESc4BbOGJMH
BxqZDVdycb3pOTvCjoTV2s5FV4Z8KunLuA6Wih7Da0WGK3fTHEnIYx/IUN/tqlZr
NYrWk4oDJi2RS1FsBn+qL0VkuoWPgVqKiy8zP/USAGk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25696)
RQo5H+7MVHHAh+lgxzhUFMCz9TAjbKkf1x84hTnj8tnQ3/3mxVlgEzR/HpVhVwpD
smXmARR5hyK21MNYJpM8Eas0HJweq5Xj8wcDlsaZIXFwixlhv4yIWz9BBkyuJFNA
qrOBVPg1fQvWnwBnvSOi5DVgEB4fQxNmX0Ie39EBRZRLLTyzbaMEDZFz2Crbp3AJ
6TIMqa7Aved/N9/jcO7gjtjcnbPFGLa8sSDerToeOEGbyHWuzS2I3Avj2uLrVB79
dh4K75NPFS5o10jrtiymF2bq7q8rpyv4lPdaaxKa5Qv5CoN74AuZXVv+S5eXeDqm
hKxMG5Gc8mxUCsDAyh0/AF5+55RCbvAZCG34vCGQRu1Eba5/Sk2aW4e6lUJzCzYK
7VeMtUzmKTWsBSSc+BBq5ikSZRJPkF1mRQV2pd2MMpqlhXMpYzxiUHUQQBWrAz7K
lC7wf8oieOEMU0SqDW78EpvuTRIzsLphf0mRzI4WIjlmP2KYXiJNAodOT/rnsgO9
ZZYLr5yvOIcJ7UZhPXCs1TfajQYKNMmpp6bAh9R5cIHEH1YGF7fgTyiSNPmqqSLe
/kHEbPExRaMt9YIGVf7f0dePvd0wC/siuWgr17w752tjlvKQ+PbT9jhRpd9kv/IV
jH48PPrAxEIcAhM36AO+ZlH56Y8KKQLbPub3mAHWMj3Jc/5s2PxBOdTda3RHgkTJ
zlO59qbne3rB4jTJ75op75+XN8hqqrIqXnSHlZ2IcnJUsMKMJOoYIGAURzyZ0lbz
AlJTE13ZD0CGMP7pqkyRSbpymG0S/IDdTU+W6OB0jK9YCNizSpIYN7IY7zzrm+EP
5ndNgRYJD8ZEsm+/U4VaMkLiASvhNuxLrMGEOiPNzZLJosZfPV9HtKnUxVc/grDq
bdfS+E/J8fGtVUN/c0Y6B55XCP1bgg9WZ8vhmWan4eZ8eoC9c4rB2yKmUIExMYL0
0BQrx6BvgPLH5deSD5zeYi1mQg5nujYPDKoBYetDcdb/bHJKMsW5+I0acdUYrOOc
cpcd+ibz5MbWaErjcx226XgXES727GTQtL/ndgEczhWmRUbqhniUdJb/QgEU/k8e
ZMGvtQ5k7km206f58LhRF/Xhc4rkHa9bo/lUl/E03ghjpyyqTaX6bC4sFGvYLUDN
q2Dk73LBnX1qeuPdZtXIbNtDvFk4pMbYrHZ4uK1Rt8eHFp4L/90OosHpnmvp4y8G
mhc1efPgst5gqhi972q+7hh4SuPKg5vCe+2B7xb0jkT7DH/GiBxfTM5+G4Sz0+v4
o6UuRzDNL2iys/kRIgRBZ0pj76ddDPSoNy49+LrYqxwD3X2/8CD+qkvulW3bq9ZJ
DDYjqHgbt9QbMl38/pA//ojgVYdeCOEQgN0h0fibaXu10y6+aaL2vISL0SWwbv1r
fqPn1fozcCe0QW/CHjgs2niIVRvsuTuROmbGKze/7RGEg1DhM3Cutp300XDDRS+L
kE+3UkmklXsk7JFrSvuvY7l+anMX7J2lvOeABP+jQfhgHbIuYhKd3YSqr/bdGt9r
3ayy2ewJKZ4/Bx+d219bgH4rkS5AoGPcCj53Dq5UA/mBJBj05bnFyBAfyNSSq+tm
sxzpuh7zvqLFD66BaRFEfjbhlt/ofXQdk1jUpETdozgZgVzKbTkIMOPRsfwgldhU
oZRks0sQ5rYzfgLQV85LVtfQm8OtKHhtLfXUs36RyFlfj7m+5mDVEjS3gQAncqVn
D4nFzorBZIe9BGbqnQN/oP+Ij9eXhEI9rXUOgdTtFdkar3Dp2bCPfFWlNct6Rl4l
UaevJCfs4vQut1CAjW0+TN+mDNk7J/0imUSE+rHZ/mz8AgoepGy+UEBRH26Y+KC+
j6TLzc8vijDUNDzeIfA1UXjTehBFHDaTAc4tDx5YKdCVBPVur1m7QjCUj3INTaYE
fwyG8NtTK7TsY27VqvJ+9Hzv7H9BXxlv2tQKUK/ai09nuA19cR0zjV1PaydFWO9B
WmdSWb61z72VV8zqfnwRcZEBBBQ+3o8HCTp79B8FN/F0UZN+X5SRrafGL8OymWQ+
33jHCHQYHHX2KbcKs9NkqBQ7B0ZgovMUOqB/l5dMmZ+ZzNqUBZK1fEWwyNdBrkCx
9QxHBXrzs7iJauQMsfTZmO1CfP+8ll6xMgOjYEyyJRutfiH2R63sfB+ZWoi6iZzm
E09es3q0aYe/Zt21n2fxSaMJ09db6S26oiM9mLOGKXmRdlKW6/3muRm9/sBS1Yby
fBoqZ3BKzrF9/7G9UMJ0p7NVQplMb0AN/bUTz3a5pqsbvXuesIUCvMxc05YE8mmN
ahqfDRlaVu8JqQB5abvwV/+oLrcPTcmTiHx0usbkvdsWupjoZmAjQHIClGCXMmyL
/fLx7TXrqy3NW+mypwG8cp7gnBZbFwx7O/KAb8ILhJeVmpO2Tm4lXXMyJAA3AEKg
zF4/58Q2lxCVInrqRvfQY2l41X61A6okkWuNN6XUT91voO/uX5iaxfonMOiGzUDn
A4wrAgP/P7ls7FJsWqGMIDATI9WG+V58LQIQ+OZgZJkDBaYhhsIuMrA/7tD7nvlB
ozjEvIln4C5D6LHt933ZbV/nc/tqjB7UmeS33QaNSQjpaNUU+d+RJC9XlckRLjRa
q5C5rvMSkmWeauuSrK1zOAb33/wpeDxhvSeA97qxxk6Ma1rq6lPpRsRsA8TjbZEh
R6aY4T1ewqx8NoegrndAXShbWJKkHJw9yxlzuf6mCwfUpkMpryxOKAyzGlV6HG2n
nggCWZJR2KEflGzMA24LrABht13rZCd3TU1ygFoLmJGqe7mia1qnbKlgZwP0gXGS
mhCxnwnSiKuMZd7fuvA1/iUxjltgd2NIa1L6SEcnjdGb/o/TWylYNB7Z69ZrkHp/
818HppmFJQyWdKUj2F2fY0swNamXtOSLsP3K2mA9Yt0bOT1p2tKKSHc3D18IYsJA
10KUUtMdKCHrgtyMRszFhFYWqh7vVY9pg5uw42bP99zsCcasYHmxC+J44cZ2t0iO
9jx3kZF9eV6BTAO8qZmOZgmwyxG6Nc7Iq4IGW6103XQFHaKUNlCJQAL1cBf0e4Jr
wgG2KK/L3EwW/E67vY/qtf8rIvpoZMXLegt7o62j2bYxwJsuSos2hL0q8NBl5E3T
jOqkhIkQvW7oLiNog4ziYYZO8A4eEPmE94yYddo3sKd8ZnV4eZlgLgxkm1auxoOi
9Dny+1Ff0QmNB3OsN1gLdCpV3iiwcFz52OVKZRVFgQsH7R0oVDn1iz+ZvDQ7Xhdf
tu3eGmyBN+xMc4CbibVHw9DlvYHbcfw+H5JZX6o+1sZ9f07z91UGpMem3debfENM
Z3JIQEWQCOZwC+TYINTaBJBJalvtYC3lEx+Q0oc3L5M30ZYmjypd0M2TaDfbp8OI
H9CCH9pOdNkYiMxLjlscNINudv4Owz1TzQSzSgCqyTS3rzZdMaTQKVfDiyXxLA5h
mVNqroQ5pptxjPM7PVTp8PaqKv6VFzgrtb9LmDqNwz/xYdvt1xiyfxdaOJZX+kVa
EbitR8wH/R2j00B9yYLB5lBeEqoc59eDpF0Pq3qNKP0BRoMmJGXI87sQNQAIK5Re
9KMhJpKOd0B4cyWtAtvAYrhcw0QFpVKWUN9+vkm4+G8GqS89fVstp0fBzTV0i9Dp
S/t+AIG5GLcNWqaogMNB5KcRs1gTtAMZtFhIm4+lhca4ZzhkkBlKqVmrjygvGyjy
2QW/C/oy1E/chrtb3gaFDRiELIan17ndRkNjFdkxjPCHEvYLvv25kLl6Df49bdxX
4c4+sdy2YSlAJaIGb9Q/QZb1rE7pX8fVLQ/KayTSSAhfwoMgmUBQ2XSmCDn7ZFd8
ZhoMeJPGzR+VbgxZe4OmUnAjpkfFgBErB8u7eOZiSOm5KVtvco6yLMl7FFgTg9C9
AbHcutV9dzzHFwYgrbqUbbgbJrmOkhhWmUpqCOMOBCqzu4wceY4Xxx3FHyQ95nfm
IIuTIOhLcKXAO2HV52V5LUO7lO1TTWEHvXgUz0qqxGUsxPXalSj+FU/z1fLCx/Sf
SVsHBqsdfa8dwEfhPCTpYlLjnznNBojMQuPSBbMyQnBI8Tzb4hbohgDwVnFz5vgw
+NJvM5bBbqg2Lm3ugeIIsVpNC3HWiENfcT2B3WMIQFsJW3jtq1mPJ7EpsQR3K77+
0haKaYGCVVRE2xHanPnFi87sPp4c2V1Hbt+RS2zE4pQJVif1UACCkz73PFX9rBok
Sw+Z5y3VNJ0Atc4Fpq4lBcfXCl2ni2eaw2umfpIQfsBMRxxBCmkLc5jW6WwZ07/P
6L0uDV7dwaEpwaRWxgzcFfRN7ZjH0u5PL8Fw+bXLcN5gtd/mfqmbLLmEhnc+Ut7m
2WF9WH31bk/vyXr1dwX/qYUahN+PRnYtX+EuYYyftQKGSuHUDGwLS1xWmiJn0Qvn
Pp9vx4VJvnpmOGYtovodMFTSYyLX0v1rfH8BAW+/7fScYMg0QX/rleMc9Fd+TRhD
kwUFw9qRUhBZjbXEI7S/cCy8e05iwN6x9zpTJ5TFWgOrxyxuDs+RUL5Ad9qKcC48
TGSYmOUTMfuaS9MpjO9gd87osmoi+TQE4XOdVUPjXUXnwpb/OwPdOeihH9fQMt3K
d7NJ6lLYUQuIWeMgAUA3ls/om+MBDHqcCQUWTpa6WWYESiSCBpHfNJ3yNryLwntP
k/9C5p+uIAC1OZeJM2LD1ykRzsB+fwbkTWGIEnkTzl2L687stPo/k6Nndd5m3EUP
cH2StVLQSsW9c2Hb1m4V3tbmGcsJjGtK/F5qQasvjwIdoP/vhAmOqZxH98kGhAz3
Gfw7mM8GbWfMHu944Jx3v01tLCDMMSZKoi1HZy8daMVn3nSQjN2pN0zgyMQZK1oq
kw/tefoPd87RE6x74IYzxbeuFptoNGVkuSLnH3IfnwbqKlbxHVT9Lknehd47if7s
Skhq4F4GL5pjT0gcrG0nFw1OcelMNBN2sspn2AHJ3nF7knAJQyhmecxAsrsrCker
L051sCYzQKvz+ef0UxgeKJxVOy6+AN8Eu1uh2gtUvQmLFBErA2h4MCnV1lFDW+BO
O3ByhgLe7dVxgjDvuCBcTdAMFuZWw2prVQ60xo08QDIhLxvlu/htm3FgKHPpqRY0
J4m/JN4TffPjwdt6WgtMeG39ZrGwcI1MJWw04vfknYOA3qq8Y3adn3VpHZnJEOdb
GKJzHx3fsKk9StlP3TRVs/C/w9InBfOIYTjHSLTVyGX4CnTojE9LbCnXIBwqdtCN
NrVixXu1u0MPvRwDeiazkuwRQXHPX7IgzSwQ7RUFM+5c4TvD64010se7gWFsVohy
2UnOigN1XZJpRP+u4Gc7qlfHcbQRTeUlW5OEXASrrj0rma4m3U9QTKX/WfZ/6vmH
3fd3RcOW+YxDC8iGXc2srvmt914EnFyBEje7gESGlCB7s3Sa7cqqpCTQWfO2Baop
tbrtzbVGKLxWTfCU4q+BQ63Y7Xp09GZqPOl5NkjiK3gVZWLnsGdpbEMce5Tq4haz
mMkY+C0mkOnlZRs8bLGSHFvfG/KaUJiqnx38jeOBocnIc20ZafgPivhYzPNoAk2w
dgPCSL3STGwysXo/UvyJ1AWfa0/C1cHERRyrbNrb3NogIOFvSVPwL80T189EI/cW
2oCWyLL2Cj0itDAaxiSFUa/rMAXTwUUeD3s9u1m/6149peYz664lrmFeEGO6Eili
UxNomP/zzpvPOq36qkoWbC72W4LoJ0IFPYfPp5c53l1HHdokBX6r+3QsOmjgLwYB
mfMpLtFZT8zSwJaviujwHMKeA0xGodwhw4OIYSWKuMVk9RDZ2o4xz1tQ9VFsP88X
EZ40ukuq4CWK3K2v0zi700b2Nxf4nNut8lRkzaLpPUg5817FAchkZ6dkKCbszlM2
YfQEFpUWBBLaErzyC4L5Mq3YP25tE+3IbdFf6NI010LbIPmSXHe+DhgstV7hwQgZ
XYA7On6/u2CsDirBGYkNucRye43MUdVmEvbKy+ePKBWZKH0QW5Ewerke9SlZK+E8
lnAK4XbbbCG7zmlrt2cmmETj4dMWJRkxfZ4eF3HDz3TsWoWUQ9bAUSATNftagiDH
977lUdbhjz4FrnTcNZMp293dkodsHvIZKOU718vsdpqb3kkwvdL9dqEMR1WJAnrm
xE/V7NAyr3uQgLqB+SGg3QTHk0xUhke1VnE1mI65fm49lkfZM4e+y25xjuciWAto
8dVIOr3592WWWFgbKM0EAh5ty6mDXUwrThpDxyr6yrOVtVVabc+b8+rxDz8CQF5c
On7JNsyYWcH3vderhTUmGiaW723avAeRahG9G1jC94dYHZ0jfTt8D4REyfyC6uYu
cWaLX0estGELsC0g8wECAde6wdqZvgEgsu4lNhzusl/eAxD4vYy4rogrqFQfuUkP
oJdzpsLA2XFsAXai4BVup0phk1ZW3/xOYNMyzdqKEdeNu+6TC9C3y7zUOLdbELS9
8cIwer3fRT4DWa7ptSuXsUq4Llxw2Kfkhoz1GgDx8+fN3woWMAVFQIlrK8IROH4n
2hbuKxXtfF9ImCmjsNvkSiDgfxJqo05vVi8CHHwzpWbLCoiv3LGwR3NRd1uMz2BE
av4XjEPPA+/8gnnBCO3ZycaoHLTQEKeo8ZiBbBQ4pas7wlUf5qvRInncow2alD/o
IpIdrtqH3OXJVqhlz9a5JmzjblCWVbM5FzWrRzVeQ9ZkAbFXqzk75I1/hwZ9UeOC
bYea1zCx9UZIidT2SAvvuVLKdbgr/dh7+9Ev+72t/nrFeH1Gr/VBUNbzKsWGdFRA
d8PboQwpOzKdJz53nHfKrTjwJNPxP39kHw0SJKEzzMr1FVNxkaF0aczAqxXixn+3
X0GndA9PlC7jfGzMoxNW0ruHr0Ra6oOoC7ufDGpzx5ZJIrE+j8SP6Y/2zFobRfmy
v1S35rNpcLfzDP3Ll1ATVXzM4bjXM9Ul4m78k7L5Cr1T+mL48zBWIRToE4L6dOAs
jZgtD+fMuxlbUq7TYswXMn9G1M48EQWJsmGHNQWqsYauGwHV9+EMvuuKz/6Xm5gV
HRRjkt+nHVcqrQc7LvOC2mbyEwgK7IZ/MxP1oso0VFL3AOltaIN3Txm47DFLW6xf
iAXO+4EhR6LH6pfm6ZAqWclKSw1fn5jROPhnoeJk/xV6dxke8ATh+pRZkdAG+EwP
4/x/G0PsfKhr03KQO07+FNvxWQpwQR2IiM+Bn71KQzjm3FC8A7aoUYVJo+LX7mXo
P1XnvXC41twsnXSA+vLgOxZfe2MVlF+O1rZtreLcsthM5v3cMUalUdYziVGg3JYd
KD7OuosMstAKcxUr+Ra0wIsj1zH8XGNAXOG5OsVnTvqgjd3CJCUw8oC6+F6dm4V5
ui9thW5mB2Nr2unMjjFLrq8g+LhRwGfyiRTFIfZU5Q6Ac8yLmefUKz7J+gUZVfV3
ZaiNb8i6HslIMWOPIHx/X79aqLHiV87xh0r2aE9kvN+FkwvBDopwSpSi2HRvvqXQ
9UozL0MgCwtYQ9VGTzMED4ZIaj5nqakdmYbR+2Z4XmkZtR2hBqDr2X35WkPN5p/p
HPItVi5GnLjD8rwQg/0QdoOmejM5tkr0ewGWHo3RJqsVD9OQB3YYgJtn4SnDLc+0
WE2szg509GJXU/tiwFnzBunnK8Ou5s6e7Jh4eeI8z0sqY9mPd/rVslrDSwLUVv4g
XC7/mbLJn0jmS93nkVfP1aPQ1/1ypZgvl42a0+r/QPtX5la8ekUGPFpMHsVKF/ay
boQcMZM7LyTaP64puwD8W96rEC+GnGO7AdSBuFGdMVzgmWgJz7GTHXjdAdQ+k82q
eAVQjfej7gRVj3Xqz+ReAF3+H0D7VdKSSmkI1dgIkmYrI8dbmAa6T51BLtUTjfge
TArHGQpeRsbYqBdO7bTE92bLuSasKE3tQF+bihtMRtkZSZ4EWuFkOnyDK5DzeHaa
viDLD8gHcyMizloO14Gy3mk8fsWM1FGzv5tR/xKap7osy0LtmBVP/jtV+uDvUnYw
6purc3BRZqokox8Y6dLE2ohLy8e170L4tey6GqTq8ub7v/fGbRzqUwkYyGE0IzQz
5BpXR+bjpAcxpuZxU+IKP2oTYtW6S3nD5wxXYZ6if5Ez2RoS9YLljcllBqPddYcg
Tsvd/PSFkWWHasZG1wejApvvlpTDXOV+9otoc51VmUdc2XuDao7u/xOg3JJwq8ki
3+ozT3LLWpC0XssCZps+J2pucug3k3SREksM6Q0GAHMvJ+WUUhXqJvOH7iLSzzsP
VRltfrwogp+tvyxyCaQEapR1jwp1ADhDRavjD+P43LCGd2IDhFpJALt1+btyT/iu
dCPqAFAaUk48hWmx8JikUUpJ1wyXUEpC+SHP+HKOoNzbESt5T2eO/hoUxK2tof5r
6IwBGVoMkZ1WvGQQHdYs56Gb2dOBklXDcR98MZc+twH5TYeBZfJDKOKQouFtb54F
rhUO0Km4r9dIW69vD3AramYrUHrrFNqEFA410HsELF0ZmELSw4JoXbEK8u+xd5ph
I7XBBndzqEHyXkYWE9jyOKPjm51cYQr1LuZLNCaiVc3z4Oj+eOc7ZJPPar4FBptS
pm8e6ztn21Ol8TJB41kk7g4MAQQnvbATK93PZsrNm9b6vY7q5Af5a/h2JyhWNadk
m3xUxIbFkgfwpQMMwB9DNM9Q/j52OJY7ckhkxDgkhHJ3F3FhIhs+xNXpRixjeYyh
a2VLkC5Yl9JmAoPTcIE48Ro6iX8uZt5zEr2Q93IHT3DhQCSveGWsVrkAephqPmO3
RKovj6mDWSxmYwOCtR8jv2+y37i4EklZRTyJ6g4K2tmPSaLK41CPAAm5aCTyPQV7
4YGUxEttHcFP/ke+smTYCRpNfdnXrnWyx4yNh0R8vwGPv/xEK/vmoTGaHu7cb5FE
ETRmSn5ljo5l8RQEO4ZzfzME9GWSobYlr22DAB8pVuM1F5u9JWXA0flWTo2j4Mfe
E/iIAgZd/pyw6n5zeCCWn1TTJJWyuwLCGZuIuxhpKglRKXqE50w4jt2jnymr9w33
BxSy0XockXVQBX9wUxlm8AmYkDr7KEytF7FBfVwWxPSngACktHhcPDB4Svfr4TcB
3a6j41oWG24UlQBFCflBPCUMrmjMrE0LCAuLpTrdq3q6M072sFLHzeWnTi/uLM0N
dsEFLRhS2w7g6qg9qk+TSxb8RItB6ZHWF+oPZ9VZy6WuSh1XAOorJKsCINtG3YZC
aTA9vO4c0WZRs/7HpJ2TbcdPQGcMtWsKhtGxF1ifgus8/Qm/x85Xo/q9H0hrVKzY
HEJ4QGqZmxOt0hDpViU8eEs3mEmjfMFgB0podp3FCxB/1zp4KEMTkzRdPdKaPTGu
HmwsGNX5ntNHS+OWEOdMkY++OXaxSQfPkUFydUm5XmxtiNmj0290zCO16hTxzwO+
f3sVGXQUCpHir5wM/e8FiUy9Q3W9LGFu/g0aobSFbPcG1asLC8ZsCmFwKFoKe3wL
F7ahKPvgmlahrIQQH1Xm/yM85WZ40uWey63zC0E/oQj7OLVOWGZikrYbHlYYdA/2
t2S7UYMEpvieXizgIml2iE3PaEc6fCNCUc4SG0y7yEKZK77bTwcu+fRppkLlHP/B
A1C8SCkqh6LX70X3gBEMGtfID5zke/TB3xjok05t69nxE7YIKYeYc9MlW3rF5YfX
pi/Oml6LypkyQ4vkl7bmr51o/+nYOq9ZUQw9dX3bRhfJOMP3ihB5QmKFo8yzxEZO
+xIBkyxPRHozGvU0yD59InJJokyWJE62vmFHJTz5AYNz9pxd/JHarh+2NzGihVp2
KKDuwX39b+D0ZPswj3hnxUQ1js0fphB+dGFrx7mDN19JFI4EulTLGBUIsmUlJL3o
KV4vSMUUQSFtx0kCwueZShsj3w+41W7G4ozD7ce8NOynkdb8yRzQKMU/yBC6eKqL
vqaGLA3A6nnZVFmZjcu1UmBBo342FRW0jecBiu0U+tLABKt8Urbq8sf8CUJsvF6Y
9oBx4x/R71TE/JKqyj9sUlCotdGA0wRtZgywxJ//9wE5SczMzpExGMarFl1bbXoF
7L5wC/oL6eiGM0ld0pkEhaapl5zZSBBfGgngq+ATlv/Rvc0yV4eikuzGDsVSySyq
Jv+wb1s0OJwn8pPyqVijwZDBMmO3QYXikQlfSMgaeVa9cMQpgfCrDoJd5nVUKufF
NpqxR23+CuK2nWwQzCHc7PwsEg08JhGjprVVOkOAI9rKvi6vQ0J3yrdhtpASIdBq
MaPUcwfanETyjB2m4Gm0xoeiz+/1mSEyJhzB3PxieaHv7NFopIwLTjt4uOgWdNlE
m6hEVreS0kfBBM73Amc96Wpxd2ItRxJUZoJVGw3JnSHAOIjqI0W0AhA6S4fknf66
TEWFqRJmkwXHKPr5Di25fU1yFEuRV8Zl9a9rF/THyJJXISJHqJaGQK+2fcb3YFxc
eGJel6sTMLGHmpcIVhoKDDKvDgKmKQYsCsZlRPxyyiKnFtPcBnX5COk3MG+Z2jXr
o6ShzNKbUXNyv3d2spDOPkgbXWWaPrTGImHCFz7WLp0GXJTEYCrvv+Dkg/OW5BDx
ukvoPmSNdujiUh5A9IPTPWY2dnnjMauyykwvTVHXRNj2x9FZzMixfzXaZx64TdBq
SrRmwgeoRPUzRYixsnYUSr02YA3nVANVnQSHIPZ36oPj/zRx9pqZMIm7nh9w5Bcf
Xmkdzc3vYlMLN9ynNK54DLhN1UB1YEalX3oDO6Z3/AGI7n6OJCAK+/40FOgGtGE1
HENixAma84JykzIxs3iwYdmGaSEMyaRPrMQVh125+3SSSazII7Bx8m3ctaKEOA9A
X8nN/cq7RTIE/aHF6DYCJ+9DndOIKjSVM+zm1mtyDkGVwAejkFNPXnM/msMsT5Uj
3xYBGrcmaFFMTVlM2WG57VYsvVHqblT58UbdytgRAxZlrfnU720BbSM9Db+R/0Ul
kQpphnEFA60U+878lOfCzwBEHVSi3jgPYVAwmVNd+IjnM/Jr0ztG0hE/7829d1Ue
NJq1EHTzY28luPgugU8b5E6i4GT5FD9NwG3hHn/37UG2c/UuD2YXWym6MJKt63hL
kXTGdjdOPW0xFdloNMG0nkAgUnAa14Qh90B8rdJRdKEtIQcO5AzGDFeeePGiRUDo
aYfnyabfC8lCik/4FniXYwsMgjrTDp7DWGK/a+Cx+tKZjElSrI1maVuRQKNoFWUY
A5eEid2AgXm30b4UVnPkwpHjMq13WC+AvG689sOwDEhS0VUptL8ZatW68qK3RUJW
AmW1rkIY+NqXSWlrf5fyWKhMlUAN82bHkJnLmf7sKtz4xEiiyea+E0mBza5K4FvH
jAWLFLFzYQXwXJiLORpgaJpyW88XACYYCt22Eq9Q/8j1jHUPRfIj4BOAlmoHQtz4
OS/SG70RQaDbxoVTVOMRc6s1C0OQTT5xjWQybbhZwupusGbz6Af79neEPiw2VcYo
B6WbmoCvWqiLMxrQ84qc3dKO62wfDpYdlS0ZsDYGHht0DCpWKLhKRwBnoA6DUCbH
7IaiG0C+wkqSiVxeFg7EqmrZlCQuX/c6chw3oJkRzEY3pOUxb0K7o4kJY1Jf+AXS
LJspcRcV+agdnII43WNatWWnEpCG6TFRH95A9FWeRKjLXfJut6WOaCPgSswDohC3
D9SgRUzk2hIdaS0xle9NQjUcNmsGiE9GUAsh1VYYw+9YLfGzE+4ad3feSQOSjcv4
QQA5GvQEX1typ9PbTN9MWSDsMa6ERbJHtlu23Bjq09fOcm0UGsctbky0wXJpjlbx
tzVXOlu1J0R1Ys2/hDcYh5bOFv2LOo7qCXbg3R+nzrKPjPxricqhh1vco8i92d/S
9I7moQvkk/bErsRw3FTmwBhU/QLio00eiIKtZv2jCYvlznzwJFBw+CpFhvdHKkXP
UzD8YT4ivi9saDWyfsITPkZ6yZmm6sAtbpVhrX7TjuZ2LnzslwacAh7rMdlftH59
cfUAu6RRUwGi5heX5XNzsJfebbKzE8rFOgUuh1zJja/iC3y+h9oq/CIT5mHEU3Mc
SUFgoxcLc48EvvH1mXDhR2KZRMiTZVp5d8nabv8ysnbnwCg0ovkYTb9szdZuGE9+
KjrXd0/qDtgBrPadM6IxVq12W1SwaFCugOX6XDtY+LFl/Ea9tmJvswYLUkiXbS/a
oO0u594dSNxWCjJW3updKcHsoNISGjsXfukXcB25B4j3aChdKt7dao4WPQujJ7/H
dlnYlJMkNpNmrtbukqQr7zdn4G7dbJBg/nDG9CeFGCq5qT+QsC+kg+FCZHWYw+H5
c+lRA5tNxzdBMqi3cj2BV8CJeBBA4vdFYA1hLQ/W7rn8AuMi9xp/Z6PaPWE1lLFK
itonpbCgDP6wIIp7y/CD1SqxsT6Xxjsa/tKhBg6rJF8gEm11BFnAbnxQdgCqecbO
7fraU+dzKPSCZYzcL52hg8EU0cLwh9hzkpdCpVjSPrfulMD48+UhjW06X7Ds1dyz
ybrB1ek8z2IvHkCJFmhluvHsHyCuFGjB5ozLhhFdhp1DoGgu4BLBz86x+aFVmNrI
RFWAFZMHMBHsiZAYIZBOrw23Xo29kS1OuZB5XVHPVSV1BdmntX3IGa+MgyZNCrok
c6oE6hsuAWXZEUUHMmHUTMXP56/gT+0rv1gAOZu4BTHpxSrM3wSwumTQ3RKJLBTi
potCJwyZ9IdKqoZy5xsNLVLWkjX3LBaNFYJuTSnqz/B9EpbGWg5z/htKJij4mmk2
UzvvU3EXHj5y3q23J6EfX8KTXiTDbsPq6LvCSz3Yi1NSsBI+5YsaQfRrPiDEuwHE
EIB5C6D+zzXtlSWav+zu1TOsuDAudWGbDD9oX0u8/fmyCRa/ky7Z2ghlhchaD6ZR
RwzSz0Br1uSTorut0xOXKnfgdSAUgdBOv4U9m/fBz5r3rpjxNsJZKd/l8Xcne3Ve
Fm1tGJxfyLoEJHXsl4qUbrfAMvNrNRf6vLzeFYYEjCFiL+gEG9NZ/NnExNuOAVdH
nH4H36XHbH9eWzmOuDYc70RDIfg+rJ4i6gNLj2+IgAUuJnuETRP8FSRxprdHY7AB
YgmX7IF2z4TyO5W2kTY1DzRIzJgTKvbd7/v8rpRvrxot/7jKHB+gOCwYJHBOUZEg
fDHhXFtjOZG+w6/psUleO7+/CEY6SoqoA0CRHMCEQF/O5RS97hVZKbA13nYT8NTt
xt4d8d6rbIhIp3pn7M5woUQf1xyWL2egdilSrEStT4ANDCfgeOzwhMlsYwqTvzaz
U94cnri6G8UmjQCyv5N28+yzC73dMUT4QLfjUSt8WBJsIrbyt1s6CJUfEcW6px4P
wToh12Vb8fXpKBWewt+RkU5UUewQ0h7dTFb17mEHSbzm5syWWs0HOlzVG1pS6YK7
nFlw5qegtIKUsX2Y/oExkmZnL734KAY8PxLmjSIRWOhLv9Mi55nshO3UFkcOYtD4
t7LwFWBb6Gf8Bxs6JJ8HuIlPp0vlu+vjJc6mOnxyjLI58z088V8x0B5GDMl6Mza6
NOzupBM65oiRNMHW/LVaS/4paKNAlGL1FSf8dGX3TuMy2cwSrEpzLrNd2Hbnsf4s
azOgj4YZKk+UvYJaVsSece8pMnY9+cZbJwm5qxnBmV+WL0IVs8opFdCGiQmpF7Xy
OqcYWxfjZXgLRcSinh35GYZYYHr15asyLYpPAePiF2qsZ06fDEZ1Zg75jiftZQdi
f6uY6RUvF4TmGJOdyWzBFaJMDT9IXcFKTDE9uIHB/iWZm54kGKKe+S4NvGvB/fXL
Tkg9iXDStp4qROnFY86uyFmTEJQw9n9NaD3XuwcQI1lYsAJm0rjC9pPUwMeSqXlB
Cx6JNkIKHhBO9zAVL8bUtHKbccnEZakezZ0Z9hAOxJvI+iFkbkOjqep6oHFKNTmF
1s3ymCSAreODWWXdJcdTrdDTWn5+wAQdE3neWJes05f+K++TjXvi7WWuCm30F5WW
gGaKgveoLkE29FAf6P62JIL8mrm06ogJ85jdh6zmsvNfpVUVTuNx98Kk/WsRct8U
ZIHBmNYEIDQeKtoPj02OltvJoPEGTjgACQA76LkaOPyH+x6CU/lKZrehFlRz3hPk
2w8SCqvpSLxALJiNVEuUhsuUkPSsI6laEi5JI9XJFmdqj09InIEDjhCsoNCMkmrR
0O4XgcxGzuoccfgpEx2kxe1yEa35dPkPgrFRJ2U1LBfThnOLRRNjCh1WTGm4DERS
5sEFDBf/gHpfrJ+SKlgYijzlHsOLWHh740jz8O5XdWTyDZCPJSvIYwtb07Rkkojm
yeZNpf4K+AoVUhLoU1dY6harRZlFcDq6zsgs2HpWfMURhKBElRji8DvcFP+dD7sL
4AOe1mbMkWILNjZVdcQuo239q9IIodEWvMlOhpG7FW02SlQQhK2HclFMrl9jYY+7
cPowfsc3rDRIictdFCpDyUnMm7CWIQXXKW8L5o7rMw6PsutZBYk0nQTiPHHiEkRr
JY3/vfR1avGBCTqIpfNoBr9wWMRqhTha0mcL28nXRWHYoSiRp5aGLMuYpUzUbWmu
J18cUMv3JecAZQKWWl2tZbZDJblmcS6N/IYFLFnLdvBx/vjsMwfUqNBgM4C8FKMo
fsk6xsh8PPnTBGxSUzxv7eTDVTXEFAUNsc2IgnJN00uS3nSqCSoRH6pm2re97N/z
OgYJHhHrYFofytaG8DOlHta8Wbe0gqm+OX6Mm8eZD/eSfgBEqKm5udrSWlOHZZfA
tOVdErHQ4SFXsacUUP4d0oX7Fn1ksCYQry41i+JZOoez6Bc2DZpDqs3FMpwwtXtN
CmXukszaRV1In4GU00vkAIxv3yFbibg6rFCigV477fkkVc07CKoPPVHc+jYN2Y1c
s0stYWr/N9E69a8Qw6C886tHyldq6maHdR0kuJUtfKz0Phb0cmfjuAPIbq0SrVNI
SOro4QxNDgGl147IQJDSJpAsq840J/+m/Mk+LVJbxuMj4tcH0il5T4bIf2+YUwDI
vi447dHpUsZgdwCuzlOipYO6FuwGOfzNezYwwf4j/dCvon8IcL4ZQThbPDqzk7sj
WtnjK+roDW+MTMSxf26DStlgfEfP4/3Pqr0eHah9FkLY5FtOJEmVedNrFo//N8xM
IvhlBV7d9yJqHFvhH22/lZgnlRATk7CcIDbAJMT+FzpKBPmCBFNgkrHBB/wiCK1S
Qs/5q28mYhRBvZ0J4VgjAghnV8F/AkJy+T5Wx7VJBzry6iSI2OriJeYkRpi2TV22
1cZ4RuCI0N+CAoJgvk02pAsZuiSYme4TkGFzAtH4Po2EysWQeXqgxiECo2NsGHfx
YAjAlWnR8c5DaseZDewvC5d1aZvYNryXOpbuBDBVTKelY/C+NIsD/dHFSU/5TVtc
JYi1/1VyjZu273cR1TZVKwKLV1yvsCs9WvYMmT+PkftzKlh7UdY6OTU6/9uc9WBr
lGdBfM7VZQoh80MBTqJgnRonZEe6DcHlTZDGWz/hF7jny6hGr6Koy/PneFYiZbEY
+2WN6G/Fhp9t3GDD5V2jD4A502bPyHVf2iPvS1onOnR/miwNB59dqv01pf0fpngN
3I8AXyMsb3tczlSiuWC3OZ/ArnopySEQnuAVZvOokTSJ/Vz28qMuW5lyIsW9p1pV
oZrQXeuM8/0059ctOreakI0GBCJFYBghGDHVE9DkQ9ECUmX0KYEIkYwFI1lktKgD
4lrz1JEoLL02y56FkimE9klWgR5GeA4UaI4/aA4JHbQYktY+Jt6MavjW356k2MfP
vlOON2IinCiqPS5o64TCJqPQc27XwCSj6LYTdz1IXUjHJoPQBGmK3dx41ol0pvLW
8fBJ74w8L/aEh9vVXH9WLGCnZbATVfki52LXnk7kPLuEQFjHdGu0M7f698SbyxWh
cEGXAi3SxziHsor+c2dT0eqrkUYW/xVbDr2uZpaNMcWALj58IgVk5vnVAJbkrmJj
8SIDZ6I8uwm+JEqJMNIIaYLzZjzo2V3LZ6svwK9ihLrlxhsfbQPXKSU9LG3l3KnT
K/h93m1ONp9AgE4Kv/QFt0wPLeQUW8oB41ZWqFuN8ZP4XgbWLE4kXMIZRknrGMJ2
ZX8w5HIXLax7CgL4BNJFqoxy0QM9tJwXZqjO3bMo33ryDONmFR0DE7pcB4WNati9
MNJADfuxpf2YgkO0f1GZoIwVGHy5zueRU8a+U1SZeDtQlgj0SY6GXbjmM7lgvZTb
d3jlth6/XsViHMcbTsMDOHRGSg13Yj+qfgSVCUR4bF1KlQ6ZF/Pu2/Qs2XXUc7gg
u3PAoHZaME1PPEOWr9LZ7JEScI5ZGMzMdw2ldMSDzwg7EmTfAZITJpKaiXdNOmbh
nQDvzJavI281N35mgqE5QiXKMLAXzZ8nAFOhBzSuUr5uUdq7cy/fgOulhBOfM4zy
w5/2GaK/GLJz+yEJ8resRstgTXEs2OTmRqTBfZEIvVGzb73XoHMBSKu6d+MDqtX4
CrmNPEIe2VKeRlMjym62tlHVb2ML9sr7e/KkgVLv7lEe78XJc+STvLSvy3AwtMbc
sJivJ28vUs1bPSVm13stQDa8wfz8HkWOBP68y3ifODoTECifMT69BJInPv7u77/+
8uJZxarkk14DjK2cnXD3DBO85kRSsnmKYDw/kd+q8ePaHd6KnHSyzHSSaAvNPt8q
43VOsijY5B3TXAaJsCVFkj8M3gp9wnL20snaUnfIECuhRI8+zj+j31Rer0R1L0sh
t0acMhO14UrepGvCB88zwBCx1IFv3AvvxKXf1ti9GD0s+Kwb61RmbYvntdsvcs84
9Bi44nP+WnYJyMYaaakz5HgD2pe57S99bsS2OeTIUf2S0Un+XoTmrJYKgNgMbzS3
CERpSj58WWqc7utmdM5OjDj670sCkAxrbDTQYseQ2nfn00d5/yKS3HoP50i5L/3T
mXDtVmP06/V20zou6RHCboCSUyy3vlUg/Z6vtf2AWKT/30w7ICPZ3XZXUeBC0vUL
t+QVobD2WSwmH7TTHptOjYHxUo0bS6BVX8DxxFNcdEHiEc/Q7H//oPFnqdEf0thj
HtbCp5IrRj82JeysOnbwrbBYOKkpio2m3HEja8nw+qHRuElirCU34QKAiGxHq9dy
AKXWVUP0qNvcgZRXRYNP4uS3wKc+jXVv5VQSc63V7en+pNlkG12829HMs89wjCsA
d4/3B8eGZJYOi177g6zuX5fLAZmDqKEy5K9vOsx3OCTeGr1lHULN4aTe9JNrcD40
j1c3rw+/DcKT8HkLpo48j7zFdlwaJHNTyTIq4DlHoBTWCXi45oAFgN+AOIkMnCIN
1AovkpZRdjvO1bVj8v/d4DpuTuQ+J9Pzw/qN5PRzyh3+YwP44LZhLSiZ5E98Tz7g
44M3msYwiaW2lQdKzgAz/0/y3+8sL34d1fHacEAkXSgCHXIx5Z4Q6v1i1rvi2LlW
2Bqqaa2MRqpQ6QEhwJqC65oulE4XosOBlcuzk011nKRJDA0fxW21ml7xe0PDP4dF
I5gQGLfOK33bBDkfMmKYYt2sZOXgNw8hmueyoZUZ8D2ODTNP++rkrNCl/gyRvdty
FFtlEHA2T5nbJ8Xmhpb6lYgmzEkzTlWTMoywisbbhJnmfDqBzG9soanQ12M0b1ZF
aYzHbLZDex48BNx4zVRxrYv65slQm9TuQg3xIx4yOr/V6+TN8V7e0lOlovDlCyVK
zHyI8fXeRQbq0llQFV2DwcpPMS2B4LM6PGee9KOevQ92GRWaPobOVAP725ZHDSqe
K9LvaRCS0W6PieCVkAh8lnJCnhJPYlaj0fc+nWEBgx6IuNOrMlfgff8MCeJuc0yq
XxYLsHe0u4kHyQ1Yqdb53ga55Jgtkitd3WDALQYfNM/H6Hfc6qAFJ1lirwkvv3cM
2IrZMc6KYQbMGNhsdVIQZgii5vr2f1Id4HMGRBNCpYVh0zWk1qoTX1szgNoBbWHh
oQ9oW3/5awTKYfAtE+x6/kurCkqeqzoptkC81gdKiZtaxHpbdfKV8uNdkoUG21vZ
b2H3++cS/+VrntmadGd/Ktp19uE/SJ93ZC7a2yeiJ4RSND+vawabFu0VX4lwWiJg
oAnYYY0uNQKc/gWCfxSgC+8flRXtlESmsBhSJGVXWxbh/Wyn6/iZzSuNCCeerCPU
4odbVDIslBw1/MkxWv/ML6NHRKjLOZwdBAglSQ2mQ6pTep9kFfmp9hVclJmHH26x
136/obFFr9Zan//NH5Fe7+NcxRdcYdVf2ZYze04cI1+x6xSEAzNV89d+4wuGNH9Q
SWod82q2UlL0MWet9m5EgPoKhCtHoZbAudq/zD0aImeaonLw1IOggWyXbUoSPMHt
kCcfxC4+LeDUmgWJhphV56+4yWZGpICnFSmPscimo4efr8s0d8Jpkajs6jPrS5NK
xlRD6GdyXoWPMSv5hx5s8MmutDVr+GpEiMQGnXbCKgx/H/Qyvw+WBoPCrltk+DP8
LyGryT/tsn4utyzZbbz/9pcasq7cz2R7LPTadXGf2HGsyYzSf6otmn43kmh7TQbx
8/bX2RaD7LbbEKncIMhjlkh30qbb0G/Hj7qYXZfYokJnXI26gm7Na0JzPdOdF23l
Ijo+FbXqFonXLcSIUzYKKE3adm4J0K6AM8tAMX6kT1YeKslK3jVK7fCiBOm0RYPs
UyGVVkwckakUMM5SdsHBtBZ7RrP671fxAELZYtt6gytgFH81mU3U5zP2vbvqCuCX
1fhmfI9jMvRiAIzlv2ltvPVQvXNgKeZPG8q9vX8WVZHaH9Gqzi2Jv2IbgMk/8PBt
xsb/RBNv+8IY7OOqz435FTgLpYiBURnNgBWKxJz3fftj1VTyc1aOzBpfsLqe/IB0
SKHkVFeT64EB52dWQHIRCfN+UhyKReRUj54oxrRyDrIzn6YJvFm2u3Om/HS2+S2V
mSs8JqKlecp5qjZt1AX5ys7nDL8H6MUuEbFJpt/3GCLeE2niNtjPDeYuwCTyF9kZ
cV4tDj6dsQLJcRCp0zmhHm3EdqyaSwrChLRJe2WpfrrSPNRuW0dioKgp2RPvtoAk
OvvMY8fTTx2y3cbR1cjDc65sdpr89o9/UupLJqjwP78CRhfZ7C8qJqxt+b7nbwBH
YPVgYYJn2vqAgUYjiO5EondmfFgMPg5y6XPkR2FVUqCvfNL8VP9c/YKQXOzomny+
Gy5AsXHdS5TKjEAxP6BLYl2p31kPziAXasTXlygCHh+ImGeAHOumGOeC11K/wlDt
rL5fp+N9/OYDwvWiJOK7pD76qy/FTmZOlCeavqm4oG3PQd/FkWzM8ioQVxSltdOU
1n64IC5cQJq3PSabuSg5cScWy19KL8VDIJUj/Gy2nViQPSAEDRnowIulTKfVkji0
anqIMY+HbdkRL9OVrmcxnaF9BVKY/nSNmCrE6GRrpE5Pe9UA7iUGo0OunGANM6Gl
w5dEt4i9+IFP/4ujBFjfMVlG5kbNeioztlZ0cJubOJUZFOhJJUiu2IbPk5kvExrJ
U3aKLpAYaDL7l1oqEhiPm5mjenu/c26486tXgFB9/AWuC+OrYt6+hSpM57H8nGkl
B04VcJHhDXGoabw4A3XJh0Mzq3NwciIll+3bWIhcEEc0DTsiUpaGdU68HV8THKx5
3FduAgVqjvTmUeC+yutgYtxdYSQyoz+AuytRdp4No9l6Yi0FU5PWLORVroucEO6V
JJUE+vjFjO3RnCHQcddt2xY0gqMcjx+Kq/wLV1quSbYHYTsTArLRzzuspYwL7Pz5
YkDpXhtyJDYiXuv3lvkP+8BrIrQH0d0gp8YVSJPF2VoqgRmZLzALLsE3o7Q+Q53Q
T79sgVFLTDUZ4AZuJAY2rswYd6eVae26JS1dRhDD+w3V8FJY5Vg+GbD7SMi/ksZW
R4q6zz4R2M2e2drN/vJ+3z/kLkgCe8o3l8XWgtfEC/yCq4AzV6cFLosg4uJGHnpX
bSjtWP4Wp+rA27gkeYtbyYoly8Y0G4A8Y0Qib1OxX2ISD4J0pceXKjaczCekJz/s
dm10pZ7S9Dglb5EPh6DMbTV7LCo99dtTw9g9rhZ/3kSi8Ff7hJlYdVizJCp1HZSG
9dmd9Vnks3RjZlwJdJFQmRzaNuV1F1os7PJyvtJR47cbEq5G2A9TB25qL45rGFMl
3YlCpt6sa8vIuIswORXUq7OQfRiMjufSq/uNc3UxZk9JJ6AFcSxQ5C0a4v+0MOer
T8ZXkxoCaHCk3v497cc+BjZMZeJMQhPiRunuowoWXQmKBM4p3iOn/PXj+E9lEzs+
V+/M3gHDO8PCWKyXdgpT/CnYE5IpqOGcUxiLz7V2p7aj/Sxbm7Yj9wRTr6AUZCPq
kzOPPcNkT1t8pzDiOnvF2pz2xDQbuiTTuFeFwCyIN4+LgU4Yun2zjTAQBlk7NLEA
M2MX4CG9PM8ym6czuVTeZRuIWOfQj8aEb67DerHSz29SrsqG4v5+3nkbUzfEO/JO
/5lhfCrQ5rqk/g+QqHeRVZ/w4Eqs2/ULXGRgu15qiJo2huloTmDNwsAOYyr/Dakj
AVIj/aKqrkAq5GF96pTZhVH+6JFFAxM0BQktDpNIA/grLAIq/pdGOADkxXHUTq78
RJf2M25Gej5svgp2E7uUpicBgW+5qgALfMsaFA906T1vnQMZhvW66SlizGgGIJ5i
747Sfx2CfCjBOpiU42y9eEL+WzrZ7FhfvmeiPUW4yjIpKXaLhJpDiUDgOzqqTfXk
exNRC1I1gVqgyplP12GtGH/VQb+Ed5kukzK3lFiYMqy5HnE4rV5IAp0B5Kwgg6Qc
n3Szo2AGPYPB4nk3JBZobvFuwwOtTeoDnIaU2A3L1YDkNhvgnXbIt4CvZKHDQI6D
lATYjLrGDw2oHU7Uxa+zaC6ncOFxgob1/XK7bQFXc/7qiv9hfaUtaisPhfFLoBir
PxfdiFRwDzYrN5ChUY0WjnzjY9GzoztZq4Jveru9a2wkpUHSB7qu13NRy19BMEAp
erSpbYEEX5AkvR7JkkyrfCXyxjKfjtYDQ20Jaex9NYOG9E9ZbYDc78ucFAJN0WNH
LmBMh1iRi1q6XbVH7HftCrYBsughID8Q/SL1XeSVJnyiPkfFrh/PXKFU+GAMu1Xr
4mIBrsFR11iND/223z4SWmH2eltNGRj8c6+pVkBaneEgGmE8J11Va8OZCOs8k4kN
T5uljs3caeceswdaoaMXsvjMZ2fjEQ8Bqv/UywfYA/9exRVtOaSNVHXwBbjF1660
OmaCWO2N/Jb2sq4WJyj3PPUlU6pN1EpGUPMc0GBH6O2Kqf4rdlyqeGk/fTY8Zdin
BIsWYhvaqHqHajg1fY7XmtRvB7HKEzWGNTh6m6qOCk9FdwBcm7RMBjJFVhxbTp4Z
E5iH3ltX9htG48frwxB33TpYjkUtNWgDSnonjQfkpcWra89dtwImS9QXRXQpmoYe
ebaE7OWA7uygQDs3rzmXusRFjNvrW3Vm9AHfm//uJLQWF8Zm2CrScemd1Jm89wvU
eZV36cPJpJJ1CvAX5rsE7GavL6z+jmz8x268Qf6Y2ADC70xnYfVLYso/n61gQyXY
ZedtfWv0lJZqY9PZ1U0Z43oEl3mdIoSesHFSEadOB/K4L39jk54JoNbpruJbmER9
1bkzaUjKwYsDKhPKzzrnA4vtojyxzXrneAJSQ5hanqD0sv7ZMfGpMLn1yAS4LQDS
uEtBwCXCcvGryElr8obvzbO7iOV8qM7I7AZNJaNaW45WYTEojoWBp8bqdtHSFrDr
79VU7/xEPnCI3tXW0As4Q49/csh0SPx9KPRm+A4+5XwZQOPUwaYj7+jmKOCbDPpE
A7g+UiqLIvLloFOFF1KPgpasIxB/wn36Twb+1P6Pgi09ruUhJxyT7pHP3lGi2giK
YyFQYN5Vr5BkzkBZc+I9bfw7hvVabpfKect+WETnkrW+0ZErELVUPhyFD8EaLvTn
BNUAWZF44BMQFEaF7WXeDh+G1ALc6NzrfpogHU82e0nKD+0J01Kf7Rc+oozIq/FI
ZP2XG1VYDvYvZ6cWRw0/YcZnmkju8HR3VyyXnYDSHvDc5PtHcHleB8utWMvPOVCG
A6b4qRsOA1alHs9dmjxVlriL/JtJXF32dAgBJne7d/sI16JWpTY6ZW1MNrEUqy40
G1yA4TptXm3aIEgDD82a/kXYsIG3DMoDG5Ek8n+Sf82lU8y5h4Gs98GITQMAP0W2
Oy7vtaR0bD7qr6xpA4TlvL33lweOHxQbZQpFz4ktXMDW5zdTw/sBp+PTcIkOJs0O
+7oy6BKNG9ZdjbkFu+PQznXVgCeEcfa7rvxbcobbNj1ORh4x+dYzqKQZ0w1cWT6v
1wKr+lAwkklPN9tMK+4644v7ZCeFtxX7Ehup9zC7oOBH1qe87F8VE3uMBl8vejSG
8cgKzic/b1MMxzPgfQVmfln/uUQE2P+vMLzBIVpatM80n1sR2GtJkeSMiRigjVUT
h4s1l69lRbAxRwB7dNlaf61ma5lJdS4KfkPDz1x8IoGJFFsaqkt8QWTE1VbUYUmI
oYgbKO7TBEpis2aqyjFFR4dF5JwkQSLu6MmzcSRq+BFNJMp0vW5g2SQoDYwdZG0d
5FvlcPH6gLlvrbdMGx20FP+aTGJ5y7tE9MgEFZ32tJPnpR+Ojhu5rREtk0m4I+76
XaYHb/1RfwnaaKuvwOQFZzslcIpO34Oh9ayd+706ZjfgSIxn6vtVASOD29HtN/G4
pSI8vLKeg0gSUM3kAr9mwDQ4ZBBJkcf3MKZ0GRN+RbvmS84Et8zdZ4WqVVMbMwB/
rfOcAdzjnXmyd01jvA1OTJpuPHXkmjEKVE5WILA+us7C5tDUyrf9kNPaNUbTw0sZ
oW/B8oXxeZBC4pdCM6podNOMdAWEqhgjjjWSr8SAwGYp7xx2CINmxlB+43ZWvjK1
OFcoaluo+4/JcmxIv0fUh3ITLMfSunf0tdL7VKNcvUijmvpirVgF9D7dWsGnBAoc
Z8iGbdWEOgQEtDlHVJOCKU6+zXQ+yNdL2iExzHwvVM8VUMK1zdI7VaurkckLiqdt
0WBeNPBtDEjUTNfLjx5oRga//NuxeO8I7lk85v6yFWx9N2Rn/bLxciAYZPe476+s
veYrmm3Wu5o7a7vMm3jBMoSNLO3M3dKofOd5D3+OaJ9LsHxeL5PcGdpKupcbuNmo
/TQ62JSs5PNz5IzgiplJfrHLiuQP9zeR0cLdF+HLzmKM0Hmhx1zhogGVITZEiBzB
OMSywWIIAhDzu+4Dz976JNTeZtvudvvTR4tXMmiextAsyZlwkXK4ZDki1A0lqvpV
1K/KzJN3loY9Ci5NuxZ06LYJyD21RjiOFPtLBp3DVXDKCjhQ11UmcS9qfIJhqLUI
Au7r3FlBZ6zJsAqtO0OdN8ReenNCXQXxQvTZ3LpKmjrK+qQ/y7wY8aNF+pI0m6G8
TsDVuAXA/Y+pzByp6VtT0hRjjmGK+aDFefHrxOx8POSTumaDkanb0cA3ztGgR1KU
Qom5RpftXXBoXf6UeqbTVa4auMmOjR5GM9zsMH/aANKEuYyNtFF/Uv6WJ9qQ0Fno
wRi6B09AKoi5acfzXL2SLoylOwt1u8c2ngZl3nglQOiBzk1Gj3efMrYtaronwxka
EQil8PwE7yVQqoUvtQzjn+hHHxsD0Vi5WtAE0XG7ac/kTI8mc3EuRa5awNA+8hmT
wEK+16rQ7j6K/gtEKhyamqkRbv9BWHxjF8VqftA1UUJg69B2DHEGokZ/Rv3JuBU2
mTlDu7W1y8ClG15oPyhD/imH2c/n1QF+0q5rID0ESbLF37YY9M0b/hGQw7otfHAK
4wsIREBsUBa/FiU+7CrZruYOqzMKP+Gpxhec1AJar9wlus3N4HErt/jvwLsmA9YH
8yfSfVQwB577jd6YDChiN5QXTUePU8bLvurRpXq+HCxKzStMAZTu4p0xD1vpJ4OY
GwvjOEmH5MoVvru4tVBdn+rKiKEh/7LmjZoMx1f58pcK0+ajE5ws8sGwX/Rr21P6
A8yNJAgo90teRs6rXV2fFg/h3OUPA91vQ4vCohzqibteypQRNCyVVnKkxjBlrYoV
5L2293K3SeSJNJDo+KICSRGugeiZvVOQmFHWhee7/mwhpL1LESxUYlwC4zZSMpav
TUjL1I3I1Nm/N1UHmq6+IgNjDjrB7gkt6LyiH17G1Rf9xjF+pI8fRBpZReVeyYKU
pIobU3voNORbbr3ERqHXxBHyzt/AjqzYe6MC5617dxDfjv21T6qb0o8RVMNHzMT0
GWGgXp5jawngsoiBrrKfarTBAr67coMKowxv8uHC5hQngXJkdBYOK9t2+gX/+mnl
sgeA4jH6iiTCQY2PA36GtE5EeZR3SObUjnZzaBBXHPrQaq29LVVW7xN+rFyqe9PD
HYtgxQd6Y+v6KMoBUrKPWXKM3pkSixxQyATSxp5hwQjH2Qa5ljbID+XsR1qFyMtR
vgAabSO12h+WKViUxYLYzTX5pwqadftchy6mzcxszdv2tnEp5g1DbZo6uiZtHGtR
ZC/snJq7YLAiGaZtcEiDDSzjEl/pYAo2zzpzLwsHxF34LL9S51pwHXSAhfmZFLHO
EQPR5T9dOLUX4n67C0aSasGiBdyx6u/JQ9mgDXBjfhgUVveyOFlsRn0gmoyONlnO
lm0eOckTTHxUJXExMvvEBVSpOBOjrQsG83TPoeKZEDxr8TUVQp7llTmehf266Yck
kXGOf1DdzQcZe10OtrV33UX/xgwZKzUypkic8App2abxR3tHz9gf98a1enmom8bR
UWtvpnUJJqiIH3EhouQbOQkGEdmSeZmaigcWx/oB9PN7SJ6BWk2MyzcayUdn4nw4
YurLDPq6a+BTN3erqY3LrPmwx3gt27X0nxCvoJaliwIC/MDRhAxuogSHJQt7+G6e
4bZRytKbL8s7Lt/mPnOMIKq4S0D7Y/9561gwvX27M/pVlR5dL+Jpldq2OJckTdmS
ys/ak9JlQDTH/15ns8N40bUdGRexXp1kAkOMG7EeDUZw9X62BJIpHXr52mM1ZLgg
CPwYMIpKr7f3tmIUOM7YSYSTfT9cfp/47vZs51yAtk2UJi+V6f6+qR/8PWmxVlJK
hcuAuFdLLtvH/rUWQdT7bZ6kPppeKEQb0syudDw2Ppde9MC54c5yHhr8Y1mRavcJ
D7qFsjP7i7EbqWoLZ2DRjqTOcTIivSrxN8WsYvvNUo8cWaxa0LuykFbyZm9yF5C4
j89XDb0bUEtLFr07w33d+ZKeFJgK3QxTr5Z92I6VoJ45PJqOiNP7vcfuKKn4/WGW
s8ZoI0yJtuGGyHIFGpHdLLaLJqCyT/fedyttyvA4AaudO5hzwOdOcJx1l9ODfwOq
/QzDAMsgNd2Dwp6h0RggmI8uhQPC22JevEGLgVOFQM3DLOA+hElTa3UEC8ZV1RwO
OnrdfFWSqaRWXlK4fKVFmettB467bQjbF/O/xeRKBPyEJyvj+ZRPG8JQ7foiI3u8
Oe9AyQ4QJ9//pml1IJyB9adBxzJESkdygBscVXlgcrG38dTAdMU2xnqYWW6RmwjU
iVaMH3CSJrUuGRQZOS8MrkriZ8EPSPtKjBMi0Yw9Xl0am0GqtbqA+68Psfwq3vtW
gtp9DSZc50FLPsQ7YXARrte81rV0VckL9FIYsO6CV6upgs3wjIgOX5b27CKNE2Iu
nNkaCSaZW/Mlpo9spZ6xBMPuFTZJBnEyUcjWhX9G8jSrEtKr8EibfLUtPatFmqwH
SkTBRRE/YPJQwLTTXAwLm5AXVDMpCVyy8dVTFH6Ik/6F1y4bAw4YqpXrgdAzl8Ut
hLvHnpwFK+z0ufRxf3WwDDaxDtdUP/bqKuoVdj7rLK1nGYgZ8MTtiTnmuMSCJOcb
EfGcaeDRvw3OGggymoe8Se6H4iI9iSZXRam6Mo7yIS5k1JfGluKl+SwTm8UlXuTz
ePPeeFjBVbmM+ff+WisIcigQ0khehNXvUfPfiyI5qVPH44/se7Ztc8BH/XtciWCB
jHCamPFUxyBZrwkdgblwQsfxCD+xpJgmWYJ85x9XC30Vk32xMM9nJCszbCTARq2W
I9oYqR+LxTy1kje+G2auB6BBOJbiJ//Q2DMJHjlVPuphU3FaHMW4yTNNmLBVCeOB
8nePEWj/Avaf4JStWqRqs8l1+Z+7FKfXlosStW1Dwp5BAgLxSs04hZcjZWAbOAMU
IaPOiWPKqonqr/thKLCYld4P42iIKpnDAAbHI8IEirFBer4w8nY7s9YtpzHN8KLf
zCFOUVWYz0l6BzRE3J19e7FmwpkqOtObeBntGPOtkokmRRqOFHSYD4QJ6Cnfhdiw
Z5J7ZJxbx5GmVskt/scdPpGM15FerX3iUlaqc+Yk5cM3OysguTgFLOfLL1WUvYIG
0BApw0eanoC09zxsfJv2at5+v/B2UJAmgN1hXWKpHjxBIe6eZFrdJXbKK8UTLN7+
BLQ4wRglu9fBbxMGC1SYN3+xnNSfg+CW1ZSZXbISYW9amjgXgjo7kGfnVud0/cTW
VB0smDEL0ur62CcPSh7TPqbvwCcvOf1OMA8ube3a0AINFGZOZFKZ0FRCuypFB7uq
7Ar03rD87g4z+RyabPykzfSJKzWVTnidyryuZ5qpYpMP7WBejl1LGTTwkPNI126Y
5eAopWn1UvQgmgDIjffk69tWofTt5MrS7frReQWHBoNvuc2xlz2uT3etVRsO9v6e
03LF4nctT438cP2JfQaMa+O+R+9q3XnOlMM0Q/IgGQVKLGDNVoaDvZLvPYvBgREw
Tg4aEOGRjOEHCyWkpXMkk6d4ky3btZVf8nzcgfHQFLayqthvH0K1jCABjnkEN/ZT
sxMa073UPe6NZ6lRVTIO8bcz+D4p08dyzViYDZ1lL+FQNN0tXT5FBxwxRqKbuEUf
t2e7ZahWZinIgQspOIojuVaGmxfNeKQkzjdfjb+pA+tnQoTksUvrJNbz6zwSaKKd
j9+W/lx35AgrySKtgoRHWH4/Fgrw2COzGT+vFHFD/w2qmuwxjC/OJaMrqNVC7/xR
l3hQckYPLAk7ZyM75t9YjcJdlmd9KxA5wdXO7G85YEfOUMdO7ZLD5Eu2s7/cTdPZ
qVHhJz5rolxGS3UpeoL/7KWH85kiJvF33vA8xPMBR9BSyszKAR6DslfzQOttn9Ov
HRJKLGfbREyDecNPzA5d5LXOUWTgcqB9n1LoCHVpmdFMt9gNt2Wn8Ib2f2a2ncNY
j2ryXLBtkqWLTY6EZ2IJ50NGd/WTGI6HXb2EqGeQ68A2LlbaWhbWFc3RWOeasqng
MFDysmb8Q2+CG19m7Jz9/+AdYnxKnirzzL6CF4o9ZruOQzxwYdhAFUXo/JaXRTFD
KCYZ+HYd0/fkaoaUyghlTUgjHHeZE8Ss0fCYOelIGclcQ0Fr6rll4y3kTECKeQr4
W5VyAmdZmqAkXxmjdQX+eb4etm8i2XLFMztk5UujNP+P41PNwF0YSwhhqYflVy8l
O0S1NApiHQhBcSB0O5VLcBeNauljHUwWug1wbQR2VoFN/adJLBzeqrPgyHctdGSM
/eT4GPE8FbHDO6Bw5vob+42N6EcRhPTrVa2SMV4Xxj+r++2FWLkIMYrKdVEm55cl
Axks8kYCLEmpnCIZcwXiePcvnv4pSdwe2xe7vNZ6yG7KkZfN6w0gl8RuYBahabqm
FVdilD2Bf4TfQ5xZ6oEUbmFuNxDY1UB1KQIABELNL0JeDvR3NX3CD7dO8HEd9Wjs
qgjsZPdDZ6VAfsb6V5VAMWOiz7SwkB1FlH95ERiknGM6aj7ltfMvtfF1d3WW4Th3
mYVCPMWFkH2BnEGQLDfoRQHam+5jZjC8O0NznJKs3KgoHEHYYajmHX2+wWiP3Smo
eWhP/m/b1tivDBcbEKKpW/dDMD7a0IPIB0FdVnR0Z2ReyosArblI/Gt0na1JWpBh
n3wz6c+89pkwBrvGQC2DVaGDOuIqUZJh0GjpBn0gN7+KCbWeCHYwvXKOnWR7QUTF
rqkWXMc/Qofq1/5SARQoVD62qCKcfnG/jLquk2v5i9f+5pcc1A9AcS2UZL/ROxIn
mOXqGfWaZFze+UUC51CJMYhzKQoQGQipYt27hVCmAWS5YGnCfMCIifTehP3Sj/fX
6czZVAbHpYOaGH/oERvAFA9mX0Tytp1gsR/M94/rjrgaXsh6wiz6oBUDJXbd+kxm
EAdbnFl0QWuVO0gYbuyN8WnbBXQ5Wh8pLzzO0Zp1end7u4XyOwqHbwRm4Do7Kl39
pax/PlFWTXnhMkYyFGtp0fo4xb1GM2i0hMn2C/N0KuLOovQlplVujrZ1cM19NUxp
FB7pVJ2PZgAjky+DLG8CwgSx9xq+fenftI3XTXcEWPIwyJ6h7ss0Hy3XuRioSMp/
Z0vBVcZ6FQZhUSBBBtiWCrN93zkN5FeKckJpBjlP5glerC1KDCovzQpSGqkY2H5G
EXRY18mV97k1sB9AeipndcAB9It8v1rGfC7VdRmnzeo1kSfPTXVKFIS0+j0GSJKk
TO4l0C5WSER4EHMuCfowAw9hawxOhMrs5RsHqb7CxUuWnhP4D1IGwHyyx86VHZvj
txrUM1xQ1TNzd4Z+AxWCtCoh0u/1cFKPMhZPs5YCuDRmWs/BUbW/A2WYdPwq/yuE
8HBVQPju4oi9FujN9B4724ypSpTWJYoF+lmpdzhiACew7a29bk/nCINExc/zLarx
g0uyE4+IBWXBBLeJ8NRR31z+cFG7kYI4brQ4vPJJDNLj0Dh4xdUN6C2MUEI507ub
kcLAFb1h6iToeaIawV+9z80jhWBDhLDfE/na4vrLnYLdbv2PN+izj9eRKl+jthQs
l+dRXMqQ0MThhUzp8LiVwvDpVmSe5fyzAzJ0A1g9EzjPngTyGgP0hlfTR8Bg+qi3
pfYv4K9uPKUZDpJqcU2SRpRKI4e+WohggMOlSUi/+WeHRrKnECw2db15S6cWv8fN
ZBF8Alb6dZVrFp1DvMyuslpmHYE65UcH+lEKjJQ6zdlzfi1JP5uYsGwA8d4ajfhv
m0og8AK7QV6WzG0JI7GOO1IQ5fzXoC2wmeOgcIvtyLrT6hnWHgUn++ijVFkjf1RR
Q1FGvYlJgIfwZFL5HjYRAEE2BQdhVqn0PzhaZUSb+DslriZIKD4kQaldvQQjj0Cg
Oq7xc1igomxKVP+IMVZz5cWekZl7cg9b8oepegWvM7b9oOiVQjW6mIiWdC/ugYLT
UYTaQLItvrPbysA9Rt3gWuvqmvAprcdZ2gY1tExEAVsyX07upSQCg/gMU9fx41uJ
zWIziMzoYsjD5L2YQNDL/Pm+11Yp7TeUHKJNI0HTGl4nJl/vhNPQh5i+nN+RxSy2
xgogCopLzaXoE2VqaiwQPhh5eCHJAzu0DKRtq3kpOiWnDF2vlVIjpfj4dvi4ZmwN
tysqtH57jAs9+dhfbe8ksq5QI/T5IJVXTJ0gBo6rix06iglFZBA9W2t3+gmHLXiA
/vXhhyKbwQORR24hrYL6bRakEsyNZIoTH/Zt9ak5PGuDvAXejzeVRCAqomoVEeVH
2vryeYXeMcAMMX6my57SPzCWoWlLsIJ5NIH3KLm9HFo8SWPXIksXOiBwi3V2WJWI
EmGTsUnIJYGhz2Xg7iV/sOihLj8ozwhTBgA9aH/9Wah+q6IxLIgP5Vl5gKIU4c/R
GttTn6aDrKxAbZTtpD9oXUEx4wU05zhY4nkzB83bO5N9CU/o1/6IWmLx/M17vmRS
0Vsu31pVB07jwS/GHEUePrI0CILZv70FoBNfFdvQY+ieK02uRbDuyr3c1OEOEUSZ
QcY6jLecjy8dtoKgdFnXxkhEYMtFlwTtrQyYSMPdX1LxjeXxQ+8MeIEtLoRwa8u2
XMIH3E6+ccWZWDFGHDI7wpyGX88LRb+th5PXtR9y6TuepRoM/AVEtM5nIGW/9BE+
r1jH1pXtZaBPWq4deCDfqbFzuHUMLslCAuPm2/6ks/vZHff7+GNSPRhLKt6wJAmt
rTf3asgho2TKRiBWcfD3LyUMeQqKzTM1SIt9yXtl6/X4g81WFktunSXsUXIMC/bK
Pr/7zHSqkVcoqrHqtp/P+MzU9ewYMDZG2q46zfkjaJapudvfNS7TAfAI1RNKGS9a
rXfc/WpIaP7jQ3QlW3PI3qV0KHBDhCZosrj8/uRd/xi6dYVQ7AUYzsDH7xBiwHtL
XPhjL6lL0CnuiKR6hH/TnWUU1OHODrMT+cbJ2CSWJJD8E+bmQHnHliGqRfPfks0P
cLn3BeH7y9Wn91JIVJkyVwkMyw+hFJsISFdcKRIbi/kbyk8bqTob/+G/tmlnMsN6
lsujlt7RAL5E8A9TaLXOLQbmqxHMuJImINcFthjk/aGzKTH3mqdRm+pUmTtE9APm
7XtyW9bHcmTbBaMZZaVNTXvyadshgXlNwSUYJEbaQHRFeNHscVPAXGr+Z75+DmtF
tkjBU3ZYeJwBHT2R59X91IUv966k8cRPjbbX12wZmWfXQFuddJDzcBdJR9OgOem+
xrozy24FWf08IvpS/zCb7WjIPwBlWAV6zCDnWqQj32rry6Tj/O5XzLDHHaPixbh9
cKpwLlaniVL8e97KWZmcMKmejTTFqNSluGfcjdmqOllVn18IgaE5/IZOIaePG6Ak
DbeJG4r9AZWgXd/1DBLEG1aHAs0tQ32D01GGItKJR40xjJ0gl8LIrIrNo/+pcKu9
RP6v7GoVCpH/JEeCy+dTuLcOSKVz7JWN1iYSCSV+66Qr0Gp1Ne34+NGFs+SNr6B2
SBL2cASfMxooqs3pwOqOLy3T1bHAykEZxe7PRb+GGAWqGaP+JomtpBHkUuYCGVRk
1RqXxO7Vwp+xrMn9qA8ImVFFw58luPPgJOCbeZkzUHyWIv+0CuNquuMnCCisyGZm
EcTRbrB7+za3KMrtA+jOdNBE0goVUE8DYorenxI5afEj6fmAMZ/Jp1Ev6cM72hWP
7Q5WeGvYOIiqUNwuBANZ8c+cMRmD3ZZR0hEbXRgzzkWs24dkKTfQtrQrRuPuqwWr
hI9tEQyf4L9wZFPNHcUC2emDZH9o2GGBFqgwymR91C9+YmB/Nxs1zbmcM7ji9eiR
0J6sDSJImBfcozfF+lL5H9TtK6QXeJGv9Fj6005PuSJYDERACWUKcDXcMm3Y2kfP
COO1ZwwYrSIKPbKod/2lVEvjK+nKp8ry2ITDgkZHGYNYCuPKF7To0h92ggHNfMGI
zbed/KBVd3pvDafTN/KfVOxCifie4vMPtEUKOgufN0F0Tn2YT1+zvMzOm9tSeIA+
Y2iXUqZq6npLLA6cdHQTvt3bQRBSH/l5gC+kSUjQ3r7pIbRzfEokZjNISyYAr0Pc
pxPReuAytAvS1sGFVQhlif30tuoKYwbGtHe9EfEa//fTfZDoGsm7pg7rnykh0CBY
4HWX6ujQc31Y98Diqz2LzyzWGqEFtojFORIm4pzeAx9mnHEGOCOsz0+/KLAT6/8d
TbCYu9GkGVYSUtwE0KOBG2NrWyVzn95DftU74ru/+MdLD8DS5N1qWsVXm/enSH19
X9lEqKB5nmpnBLD+xmFTvFhEdFPosrHJ7C4irbycr1nX0nwKhSc8LtLQNXOlkBu0
WLN0scbjZCduDqs2y7sRLci+cnRXMJ1peBeVhwRN2v44dlwlG32KnFHYbybKBeZL
Z8sYGilBsLV/8V4oFKfqIv5c4bbdZ1Y9k8UvbAa3qOgzlT2QyO2dvecP21F1d5RJ
Pom5eHAA8HyFBfNzDO92ppOFTMoFwmZK1sRoJvcdkwXbnvHMW7Es2ld9OqNeTd4z
cZ2ak+UburJBefRV8ih8lViZwXmXc2qgEXt/oJGAsxzodeJ574zDW8Il8aG1EpiR
RxKZUbfo4Lv4jb9I3P9VIGBpBcx/Mp8D5AnwvANkNdzBJTAD6m3VFAwNxG/hftNM
i9KqjY4LER7+FMYRMkKydXV8hE0PIoceI8Ea/Tep958Uha+Rwm7uOtr5/hCz90Uc
2IUr7K5peIavzQDeC8QpL7C+F+U72X4ijkuWbvAIr/5pYD3cqu30v7IlOmd25sUN
JJjoXubs9DhkuuIlqO1/5OCXxGlzmVNpmbPsRPF6nHlrYQYIUgR+CkZ9tfHofnRS
lXzwhWstlRGHs0L6EzLq1/dTV7cLGu89VzyKlWVY0j4plkKj32lDXJi8bp9rcovX
8lKrpqfSVoxNeIKHacVHr+CDGO0C1B9ISEfrYFNr5N2mfEswzJ4+V+FazsIYiB2e
R8OmfyzM2Zxp2GKJsLG80RjMzRnKd3yVrX+dbkO4QNVjhJlr+5Lx9wZSkm01I3Cn
Y93yfPOx8oP92SrrRcv43SEdc3nU8OtH+9MvWBdvCcKuea2lX/QZxPneX5rgniE7
0blrZFRZuQMdThWtqI88zszapzkilmWb3CS5C15eweMWvyC7PitxZoalH9Fg/tdX
rsOuoHv0CJv5GwXWSA28X8bpnEuhGKG4YL//kZ1JKKXkw9b0418av9kkc+ci9/ur
XHKUhp0Izu+tTz4MbHSKXFjmnuAalC4f/e2rnhHX0Dkd4APrappUpDSdC/j7OlA+
f6SM1KRJs2U+71b1SDecY3oSFTivnZ4b9LPRkBIkbRAZJilBwQtDeOBPLrvsE1eM
u1Cwk4xf97ZvSadvgAZtokOHIKs3CvC3hpz7wRQsZlTFyOokgQ/7t9M/lyRfL/XT
yPLxyEGNXu+czahxsIJGq9mZK187CbF1uGx8xZoUgejc0d5lEjLJNxGY5XNJGRFR
rRm7Y2/gzbqrWH1vGWEQag9EMttectaUUdMqMEyq5b/zN0iQSjCGBSUdVTpeOAQ9
u+DByE2+me4AJDM8I46URP0+PwpLbYOf35DoCRrUfmvRTlOY9r8BA/fN7gFLJTfF
wscDiNVaxEcGZHLtevuH/hwjV6WaIlLRbBK2ad1PwncG5RNP6ste5hbKmdXV5UJP
ZO9TVAFlPzEVVKXExNfnnecL8N62rHDJ6yGnHGf190DPTl4vlmUVufSpJplqCkew
cloM6ENDy/Yufwdc1+mR4RakWZCBLQvJTDnZ0hfQF3BOH4x2nN9oB+4eal+MyAoc
CXIb1ICyv2fv5WJQoSkqYNXvLTodPxBCfpt1Ly5+GIj5xwLmahYHujr/iGoRttPh
NLpNuOhLmAMWPP99er5iBaL+jEEHXtxsJD16F0sfXC2kiJq9xaRr8WcpPfAxxJP0
97N3l0qv4YsGQZXTDHDKl7F/JamgAuulqEnkIwtTDrlxhyXwRtIjX7ZKQ1s4EdXM
4d7GSOvjrEhi+Fpvl9H9xUqROkxdzUWa1K6y1XKp6Dj/MLFVpQvJArnRbr0sGONt
429Sv0j1wrqgAYarKA15/7C+4pAQd85Ckc9UQY+wVp3SURvDXhaMLgVGp4g5mOo3
AJ7DDN4SHhYUb5CNbKtiJjzZKsGpgrhA8tl+jcjtsr/d1yRnmc4NP4pBlvAjCiRl
kP+PEjjUYCDtvA/Gt1Huj61qmwWd3Ctw1Z80TuNt+NfmnrhlItPTfyNfVXndw55o
UL+7skh7OTrJ/FfZuyP8VTJb6jenABxYDI2OFEHq9Hof4gGDkKi56mE1Zdv4Txux
UovawNiySsxUtyRESUcW/65gLh5nh+xgBx5N/gaw3tMCzwyqjyYq662JUfPq88cG
0k5m+UXwLnImDy/ZtXoX+1g1lxrdwMB32VwDJAAHQxDaMMUoaEPijOY7Z766PYP9
euH2slGk0MrxU+oAfWLO+CKN1pTRwZsOxZ1lDW0Z83YeUi9ofczWPdWVTj4alkY1
noMIf89ZU05A3hJXPD8pQW2bos+WMynbhDkJVGS7eUul55Nw9ASIKWFhF7Os0Ove
leXYlB7jxL5Xn1eBjpWFA9pD2ZixIwQiRaQTkY0Qt6GYXaKaz5RDYtdoCFqXTvCi
JVGQqbKeX90f6hy5CgFPaMJq4AAURAvWiOWoU1y3nFFiuZyk/qIDac7PC7IHjAFX
w1FAvNNgg77VrfQS2bxMxLsBlE3MU8s7i/j3cUWsPVmYykKY4wkdwKbZ7WCZWh6e
ajwbKXon5G2eOn21tMhxL+mTTBtDTXlddKjzSX5KETqAzj5bh247A+qid/i1Brfp
NiSI+FMSjYaJ0j0p03zIzd/Aw8WyziXww2Q5Pn0sot/maQng1gCsytessf6W+wBQ
9QMKuMOduZn217I7RQ5rKR6tT6FGIjn5UswFFMmm1gpxx6TPOyVJkjZbMCW9YU8z
FVKiCqeJ27Sz0PBClnl8Q2xmMXfe6hVPIIzWvqkHd71ZPDudell4z8J91IkovNaA
avhUiabRHea3Zudd6k3EOmeiZi6iRJJ+goRfwbzCJB9l86n4R4n3itpcx9BThF30
/iHc3y0ec6UkMN7rGzo0eA==
`pragma protect end_protected
