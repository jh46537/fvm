��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���;0���[��q�N/[85��1d�nޭ�!oX!�ذ��p�ޥ�4��^H��*��i�f�m����l��&�<�]\�8e�44���k�t�CЇ�+Y����^���($�?�`�\!��?>���l3�d%�	�]�_�J��^���׿G����y4����bI���Ѣ �4�L�:�,nmE��HHDJٰ��B��A/Y��́\MD{�+��<�Fb˖,�r�I �����$^�tL v�z�ڥ(������k4zV�%Vd\�l�̽��b6��C<�������2�	��ډ#�X���sYag�v	M�¥�.���9��䴘
0����m�}d������W�R�S<�V�j4I0ҙ�fd���K�]�іn��$]��z����}�7�O`��r\]1E%! ��)�)ua�(x�= :��i�(�1 �0�/=:�lr�R��� �/��H̸ߵި~�M�50U��Noգ�,؄]|D��?X�R�z<j��_Զ����N���s�!r����I���Fj�nwH��2}/�n �}_#��P��ҸR���7�)�wR0����C��|��_�c��y*�T�K�D�ƭ|{�د6�Kq����GJ�����QiIHcPw2���}x�
�`���N	�'�����B�
>�<������,���|��4B)S(!e�a9!��U�W�@ ��4�L���ʀ9����#�&ذb�e��Rt��3�^y>���4I���m?�@��@�0&��T�+'�w�6S��j����ș��bk"D�љ�WC)�MrG*�7�=�g��0N�9������E�RLT~�0�|3�5��
����'͆��1Ԥ��I�PT6Z�Vf6z���^&��:S����!_s�@>�&��[�$ ��&�֜�`]W���� �]������I{�s�#��d��J����Bn�˓i�+����5Ut�Nw��aP ����*���^YR,"^��g����9�s���Y;"'�?h0*q�E�ʀP�~��b( �9Q7��J���W��wNI�B���z�������r!}O��z]Qx0�!���RP�5%}M�Ms���H�����A��|�e��J����B��YnDu#l�@
倴J��4<����M�Ii��4��0�M�SkE�t{+oP�iY��(���碫���A)�^�}�~�zwXa$��9|@|Q*NK���o+���`���Z�/V���>n�>�m��N�Vs�A�4�M�5��A��f�޷�:G-;68����8Ңٕi�@	�$!��,�
�}�@��>J
�s깤\f�����P?h�\�~�`N�P��ϰw��՞�������*ab���N%���1��{^�N��"X�E3��&4�x�ߜH�=5�?/>�~��%A!�@b]��9���$<8�yU�ZW@�i�yG+a%.7J��rB<G6�7��[\��Š�~��֪ҙ�B��Y���R?�z`Pv!�6���w[D,u"�ւ��tP%D��=�E��A�g ��0F��o2�U��K~2�umH�$J� 9ސ-"ǫ)S׍��4�g�}�*�8|��S-���E��+�?x%r�U� ��h\X\$	���F�FIՄ��7��A� =�aS!wVG! ���pr��7"�s�;�Vex����M�N�`�df����Gj��bץN���^%5�c����-��.C��#7�Ȏ��S)������*iT5HFx�i�-�h	T�����R#$夁]�̋/��;|=Z�CN�`���.��A~��7�����_5�y`��R���f�ٷZg�02b�e�l�l}�-}�t.��B`EZ��w�B���� �ж�GS��T��j��O���In�j>亳m`�2G�n���X�7W��1^Z��F=��h�J���B䤗W~Q ̚P��ѝ=��(Qk���&�(�����������[�_R���TH��S(r`!y�����H
��~&�����	�r��2��g��-����,^���>���S���������F��t�=_�XM��� �5��	��㰗�]FO����P��6�iA���z�vj�k1#Ⱦ�@�e*M�/DY�M\p�+�yQ"��Vdxcy+@*;��	GT���|��(l���X�����^?#�������L!�b �>a�	�8��=�s^��|����a�����,���In�S��*j+����7��K_>0���.7-g�`CXtޟ*2��z���/��Z�0\�{6�p��1g>}�Z��E���z�ہ�����(�[Ã�@�7�ݢR}R��M�J�Bע�j����뎾�~��+-�~.b1��/
���`�ت03}mE����]H�P�<�"?�_�s ��!���0D�x&x�烬��A���)�l�Yk�m����	Q�,1���o��yO��z���#e輍��|ϯ��n�6_癄W�[8����Z}wB���C! ��a߀��ލ�4e����ne�HHX�-~�����+w%�}+�_DX��=�4�I�&��
�i,��pɒ[�^K��VnN�٩��Տ|0'�#���@�qn�����C�ՃD���s����;�(<��;]� _�I�Y�	��OK���햖��`�+WH���#��,pFz����>���Nb�x���1M�i���D���w��^��n�\i�t���(�5������4$d<�&cj�9cJ����ɘl�K��"�oP���q�_2�ﲙ�5Z߲�Y�T�y79U�
��ū+�v#)s�`�>��f��Y����	h�C��<�p�wQ����lV����g� dyqLh�K��V$uuk������Qq��ӌ>
����M�ֽ�m��ŋ�n2�=��[�d��fu��q���'�?�2I�c@F{O��fwm� ����q��d(��źS|߰�sʚ�=ק�ڜ��t6mU�A�b����CRt�	����wc���
0���ߔNY�H	������+��@�L8U����M�
w�PnՃ��99�5gC�����Q����#y�Л=^塑~lS�-x�(���Է���u}6ڋ� U�צ	Z�"���Y��|3�ħ�Qg�`�oE{5�ق��Jڇ`N~�9�����p���Z�LPt�0kp�MA�`�����1���cS���[�ny1�{h���,��1gd�!]Qi��=��J|0�>9�Z�.����M�0u���T�05)I�Hv��J�Wo�);�o�NSaJy��#s�8Ꭺ���c�<S��������"l@�ʨ�>�OW6cE�h\PJӒ�G�ş߅�te�k}r���'��&���dz�:���ʬջ�QM�8c��� ����f��+���������ihm�VV|�����E5�a�m���
k@4���鉦�M�� O��(f��y����W� ���eX�d�	��wq_�V���#����Cj��Hb=>�r�v5x�Ż#6$��g�]����5n�BIڻ�{#6���"�$c%k&+��?[��k�������"����C���w���v-�Y�HN���m��dĝ�&���V�^����^�^@���Fu��j���iJ��|�7&���&8Ld�%���ML=U4?�;��7H�b�^��۳�E�����x�t(��EzY���^��%�ۋ݀���;�4�mZ���l�F�j�آ� ��x}�W�}����7�Ŝ&�,�rby�o �+���]�̐�4ݐ�\Z}P��_�x�^��(u��@_���ӓ0m��xm�g��5�u���\(��z (�z��m�8Rg[\]�,�P�"���޲��Z��ԙ�&g��I�q�<�eog��Gу�$&l@G$�0�/�msnOք14G	�;�/@j"�:H�Ug�6�x�+sH.�[�l�Ыϒ�� g���œ�),L>��{t{M�$,MzW�q5m@�H����/T	VQ �ɞi�GUƈ��=Ȥ�[��v}�I;�����Ǥ���oDp��ȟ�N;�֤ٵ����Y�R��ee�`����d
���H GQ6}>|�y�� k���pC���΄�,}�����Ùa ��j�G������V�!�;_��/��y�__6ށ�n��Ek��}���UQ1?^��2���N���#;'�J��s���x	.��Ьr�yF~��@����䚒=';�vv�n��fh�l,�.ހt���y\Ν����9�s�uY��u>�A�X7�熑�7B�*����~�,@ �����,-d1{��j��8����S�C6�Tvk�Q����(�TU>�?�ZA���`��e)�J��{���*ؙeb��y�&U��e
�Lf���[�3���(Χ�m�
�@�ؕ)O]YٴZ���y�N�F�4�YmV?Ś=Y�	���#D>[{`�{x<�S@Ǧ����f�v�Y?�P`�����wi�4�U��T��w�&�(��r�}]��5�p�F�_���e��ޟ�l�F���%�<�;p�G�7Y�c������-��(���Z�ih�� ���v�e���n�����u3MZ�h�X4�/�����-7p��i�Q�?y�o���/jbJ�m���)�;�xR�;?��{b��^�m�^sl�+�?�tս�8���<
&�B� �6h:�Ԧ�%䥍���<�0�tb��tV@��n.�$��=���
�b~�l��%`��)���wJQ��1~[7���D���P#�D�Täd¬�y�X0Ц���ăZe�J��<W���?�g�
���ǌ����j��m3������[ć1I���D>��:�����j����$����G��6&jL����z:�S��7�rI�V�r�QH�ps�����oĥ�ݪr��bJ�Oo�I�0�ι]k��|�Y�*d�-R�̍v�O)}zoDŀ�CĲ��7�@Yv�ª��n�ϋ��Ks��\K1�᧵�;�{&�Bdt2����2��F���jy��e�j��&����W�\,���
���خEt���x�	�o\_"�h��S{^wVǌ��hBp�)0u�v,�H�^M��Gd�s֊[8JV5k�EX�Mh��d�@e��f_+;|��֛���rb��J*m'#�!H���<LȨ�1�Ig���j�#k� �J���8���ش��:�Ĵ�|�ThzV_����JR��N-��G�����Ny�u=�_��{A��2����'�Q��89�f�_b#�AMа����Ƞ�#�p�U\�S��`��DC�!��֥d�&�h�ۡH/��G�c�2`i��2��fg�����.2u���];m쯡��&Va�*��Y�%3����3�kâ�G�e�OCz����)G�?�6̓8�{�VsO���'�|�*/��r�-�o@��	ڭuG��P6���t��o�"�O����M.4�+�O�!pm��ɳ���I���#����Z���¨�lR5ё���~}b���^^�e�&�0+����LxGg,E2����1J����mY��2fG9�u;;P�n�^�4��Kڅ�42M�w�������@nM����3�2e�/���ݎ��1�LS���e�HY��j!o�N5�uT@�Z�!<���FG+�ؚ�eY���=��ip//	�<T�M�1�����G,��٢�i�(~=I�H����+cɠ��O!�p�H�{�B��fgGK/5(˟��H��&��qP�ys �tA�[���}��}Ś�sn�ic	�s�J��@�>���$��ߏq�X� Z�n��my��Gp*E��9�>+�����^+S�u���mf�f9��q�"�[��Mt�H�mSɢ&�<%��wCS�)J����i���l��>hWkn<&�VL������z R�  T���v�;I��9-
�؅$�{>i�ݘ]�r���y�tS�����c�D������p�㵹���)�"��g4eJR(;+�g�q���ñ�&�f�)�B'U�b�5�,��j>.b9)�=mD]����SH����fe0#b�;8Oޙ*���oinВIwysg�rj[��v�Nf���T��Nb��ׅ3-ѐ&���l�s�L��?�Vg�R�����r7�_����
N�C��^@�xp�Բ.�z+��1�o��Qy��@S@f�C���s��W�Ĉ�5M<~H�j�s�r��R@�{<$���r%ޞ�KV-�d���T�Lڄ��S(SZ���U!e��q2Ǔ�8G�V-ǐ������?W��
�6����=�F쐍[��/�ڤ:^�<M��TGj�'F5G�Z	ج�j�·��4T�|��'� ��t4_��6��Π~*f�ޥ[��m-�\p���l��_�����x]�s$	��#|d��'��i�`�a��0R68�֠��wd��仧��Ǫ"V�<���r�#r2/���,�P�p�]����ZW������;W^�}Ex��u�]����fg���u1�����+"�Y@�Q�.�i��os�J1���j�<Vw\�Wz
� v�"$y(@��>��Q�?,N�%e�1��מj}[l�S,�9�������_`M��!
��6W*�S�m�m���ﳢv�o����:��#	;4�4vS�G	VGO��%~Nn����"��}�|���_���5�7uFUDp��dUC+� �<�s��_֕��G��mD��{����nC����iOj�[�]��1���/��o�q���?�xvp!�2��{t�
���8��`�eW��H��a볩�c�$��u�k�C��!/����uVj���$X�� +.}���� ���ɩ�5Nw ;�8?sZb�<��q2��|�[Cσ���Hd��o ����j=�9hЮ�|^���i�f�֑���{ƥK&j��͎\�֔��&ʅ՝�m1�U���z�$�(�v++�J��u�+Q�t���ǲ�KC1و�_�^9�З��0D�n��VЋ�k�UHh��������ǟ+�
�� r]��XC�ӷ�>TB�Bv��0�S���q�73󓂊FP޲I4��eyA��3�.�a��N�6��Ƨ:���7iP���}?���:�!�ji�����M�,�sR!Y4��Rg�[/P_��<xst��z#��Ya�:��{�bDS�+��.�[�v�drew�)���_�˸���VSAsE�[��=�������&��_+R���o��<g�
��B���0b\��7/�Ş��"0aE�s3,%rƑA0�H���[! J�6R׸q�e,����[��ΡB� _��S�\J��Q0H��UP�8)=[�x��	�`�D���z�����k��LX7^,�rJŨ�/൬H�w!�q� �C/�o|6�6�ޔ!�[�<��%o%��!���0�Y\1{>*��!�er�gh뵱�Hr}S�1� dXB�V5uV����7��a:��%����o���Ѐm5̢�(o��{��h����V���Bl��l2@2��HHk}��G������c�B�
SaF�Q��wߜIS��(�-�8�X��b�k�L?j�(F��0%Z9��zz=j@ǘB��6��.�]HބQ@�Y\&9�;���0��,q�eZ�wj��_'Fԛ�a9��HsJ�'?�z�"�E�������~^�&'�L�1�B�T@$Xaٛ��я�y�S��n�d�dQ����l�� �EZyM�=;�	k�Q�=�W	���l5�L5���Hr.�V!V48r�~���0�RXeq�+�u��K�{Q}-������q2����u̥�0������	�u*��V�C�>9����׿.~7�YA�]��l��䮔	��:�wTOp`��T�at@n��3�Z��oDؓ:��c�q�����,�%�"W��{��@V%�z���s�1��\��	�Z�s����+q�U�=ǉm~��Kz�ON�9;�����1�<� ��D�x�iB%m�&��0"D⡓���.���`A5r��U�T2/���^��(0�â��w6r�����|� ���D���یe78^�D��'y"��|�l1:v��~0���^`���%���U�(���q�x]"5��jZۥ�,�7���xp�_��.�Z$�s��}6*_>
"��+�<~�Eϳ�� �Q^���4e���3
��c_�m:���w��f$㻣��OY�����T���C�v���"��٫:e
����ĭY|<yY�p����wS) ���M�h������[��Syx�����	��Ӽd9��;9QbK�cZdm�m�=�r>p�ňr�N?*�0�	���+y¶y����U����|F$(a��%����(���6Xe��_��=�~�|�0P���	�?�T�]��|\��pPrg�Ԩ�v��^�w�9ϧ"�mA`���do(elZ�����
�����6z��0;�W����G`�8.��M���/ 0Ή�k�P�A6/n���ͪܞ��m�a�]bR��/Wv��cw4z%� �s��lW��\�R!s�����m�Qj
�+׏v�^T�T�T##��*�<�E�9�C��.�=|t_!<�X�G	�����k�o�?_��Fg��Ԕ�n���ܬ�X�@٭�<e���xYy)���7���Q�h�6
~�LA��dg}�%k��,�D�W��ȇ׍�;k\v,�Gv�0��L��%+�dQF/�K��[�⍲�^�K*w�s�`F:��먽��$e�|��f��
����5}�M�e~���T����B�r��E�&h_�E&<�Y��lQK�:�8<7������S�����)��V`Ⱦ�WǦQ����۾|Ĭ�\�;��Ǹ�s?`X2�U��F{"��H�~�	����wkbgX�B�Xˍ���+/���Wr|!��.QGbq�l#5_�7��$����i�۟v1\ޝg_�t�����V{� ���%��F�on
�"K*:�2R G>������
,���)�<8QW�,�*t�A8�����9&C�r	�R{��D��m���	G;�ɏ(|���rr2�>�'��,9f�X,�/X�����Sw��^�t����9n�ҷB/�ވ���
՝~����閲��ݣv�INl,�I����p({s�a���q���B:�qx"�TT��)׭U2�0{8��u<���;b�IXk�T1�`1R��d>�Lώzv\UyQ���W�u���V����Oq���a��ph+�����b�D%B����	v>h��*���!JOVї9i@܌�හF1�\�gVD���E��Vl�'ǖd84�!^ax�Eʄ�&�)�&���r6Q-���x�5�aZy�����)�p�w�^�ጋ���~�s}}Ǣ��'%xP��;��l�V��N�l̵G�cSoj�_ ��ԇ�-!��Z�.Ob��¯8�  �W`W*On�n#iC]��i(M�	��k�*K|ǈX�ȤÏe���ǭ6j=���ר��w!+jLۿ�`	5�	ϗ#v9��ڱ3�M;)5@�$U���n�P�b!�JɈ�y���h/6id�k{����$T����o�e��p>�#-#?r#M^J����P-C���I�L3�H,�a�$v���9�®A�����1�:oE-6-Ʋ&V�̘3���G�=��Խ
�1j��;�Z�LZ�H�F:���������s�?��<��q�:��-f���ae��g*�H4f6K�#;�ݱ������qFa�~x�3 �������6q\����"�䒨i�����K=��̨<���N�ι�m~7v;��`z�q�7��&��U�^aU�$���;B������K�I����B�X}66@u��E_[�G�՟P������%��xWt�iPx�M֓��i?�x�r�����ݤ܎�k`º[�^h/@�@hN�M�\��4��.,^�~& �ʘCf����nj�8"!*)C;�k�|׀�S;���������)��*y�DA��P����VU~a���f����@j�f��7ا?1'��T	s�~�0.�:0n�<}�H��5�|Qe.`U�nH�O�Cy�B�:&P�15i[�ԎDW9���ɢ�0���B^�f�BX��p�?�E�J����8�b(�358`um٦G����u��ώ,?ɰTF��l�a�Z
O�����z��X��t]�z�:���h���X�]���y0А�����^�}Ȋs��,�%J��I�	e��wT4�M�f�X��Ǔ��A���A�s[���ת5_c�1 �l����޾2�ISf�ƱQZ�"}U�61��K�[����1�'�/�i��/Y�F�P4��H,(�8�<��<	���R���/
gpy�R�ޭ�j��]�9jV�<?��2J f��b������6]R&�72��Q��]S����%�ҷ�ss+�a�.�4q���9>ɺ��~� �4�$���QB(���̟�{�����wcD�M��&���X�P��}�˽��O���cpD1ɢ����^>�:UbW�N]�4����V��T�iT��f5EѸI/��T{e��(��Ɣ�{ZJ��i��Slq�`��E����BW:�d��v/"�B8\(�$#w�d�c&~���]�T�]�E�]Ձ�~kzmj�����n2���pA%��+����話�����BO�

�Vx��@�z7�g��&�SI�2�I|n�3g��k	����a�-�e���������p��p�����:H�<��Se>�C8+5��q��2������c��/'����U#�6���)κ�\�V�,*!��L5���:�R,��1z=�7[�8\Mm[n����-�q-VtD��J������G��3� ��K�Q��vIx~u��J�r�M	0��&!}�8��'�p�r����f�E]҄3E�+���жm=�9�.^����7dۯu��/H?�Ep�{����~r�#��P���Bv\��c�3B�iv#�J�`h���4Gu9�380Ж�|�@�l�.g�%"G>q�k!ŜqcA�*�6����\��m��
g�3�M�%0��m\�8 :r(@�/����z:؆���g�P©@��2.o$�:?�s�Wbϕ|�畜�$��e�&����3���"�SW�3Q<���Q0E9��D��Ǭ�i뷗��cZ
�#!Q)UEuS��l��1��_���	��Ι8�]�"�C
S3	[���	�����;����S�`���cB�v���ˁe}����4W�N�>��qR��S���<�v��8�jQ����5�#����u�n1F�G���K�3��Bt��A�x*+(�OX��6�C, ������qv��&��ui�nNM0�q�Q�B���0��t�#����2Hs���)7�0^��Ʋ�iQ9R��� B�<Nǜs
� i�<2���� �=3쟒x�o�Ԝ�\��ӕ!��D�]�d�q]���4M�(4��c�����X%���抖dlW\GF\+����m�ؿ����F0D� ���T~��$�5�nq֑��LӇ��	D����̞�W�u��0l��U�.��e�r>>��%V4��Źy��W]�R(%���"꩒���G���u���X�ø����cͿ/�_��i��<bf�ǿ>-,t呝�$p��h{��o'�Y	��+
A�&>�ۃ�da�d*0Y��@&��.�P����:{J�A'��s�|7o�ҲI�%P$�@R�v�3?F�=e����}R��v��V�Sp��.�
i���x�t�tVP�S_�U�D��!Q^�ד��F���ń�X��3������K-�9�wʻ)<����I5Z?7z�Z3��|��>&YR�{8����
m�G�c�������1 �|A�����`;��4�M8!� �(�����9���R|Q�-�7�j�b��%j�59*&�H� q�2��7��$׏�7/�����xh�SŻ����9��-�C����P%Wk�S?Xs*=S?<�tmϒ:��y��ViY�������o^��0��h�97���3qz���M̳[u���ȓZ���MC��5�Y�<��V�����J�¡-!�$_i�$��_cbN�t��\����]����������`��Vh��Z����H,����F��AeX���ݿ)M��eDN���k\ǣ�_�-�͝GB�s�Q�z��r�u�H{���xx��a�i��J#�c=��J�<w��M�y��px�}3����J��7���d��\oN��d?N��|��@�����{�f��Z��,!VL���*�1��t˵
���q� =��xpɍz)�y�9g!!����r{k�0�N��V� !��(��G�@��lλ5��}�9���gΎM�I����E��]s��]�<1�DR��r>WH��Z�;�D˯ڏ�^)V��iR�դ]t��
�b$� ��̈�⛳��j���\����v��5�Z�yO=�f~t�����X������+�s��!���q�8z��o������k���<�������]CM7B�����oA|���(��f����FB�]eul��0����!xOݐ��&���n���qbNVfzXPi1_�&�4Y|�j
�r���ݬr��+g7GtT!y~�Ir�%:�wdK��<��V}���!P�� �	����7m��%�Q63�5F��C	���.��j��������vQ�<�Qc�+�����Sd��*|�$��{3�ΑW9��:�<�F#H��>����X�b���՝�xՁt2�)�To��m�3��3xG������o�qP@,��9H��o�+ߪl��V����M ��A����K�4U��/�w�'����J���c;!�2Q#Ƈ��Ư��a+��`��&�x�5�yx$��i9��=��6��'��ZKwَ�s-}p�d/qA�1n��%�� %;��)UW>#"4�M�Вߐ������A�l��)��f'D��F^��<��{��י�z�+}�6�����shX2�_pUj+���p�'�b�_F��'K9U�	!�q�I�����/�hN�<�\^|�M�![���u��a��![:��>�AITM��ǧ�CJB���g����o:s��$���@�R��)s`]�jN�.���5Z��U�/�ȴ]e�e}�M�U��� 6����َ�F�ضS�Y�3���[ن)U�a�f�pF�7��f�k��7�Ң�/�Q���U��]r�S����*�^c5��\J�s�G��g_�� �U`k�l%wV�ќo��P{��r�_>�vR��nʟ��&��?ד����=�e��\��}z�i�)��@;�BY�Y�a�� �H[۹�5/��4�w�&�a���D�l���$��,��"��sO튕b#UWp�R�z��,e�y�h��"�+��>1�l:P_���iA�Q����ÑN ��	- �4�R���2�:)8�u�مQ*=��ϫPnzQ���<��#���o�$�Zq�k���4�K�5!�ɖ� d��Qœ3�=;����Í�4�X},�rj���H2�򎪣�ֆ�|%�Ɉ�����C�p��o~b�0zQT�z� ����L
����3��s���΍�,մ7�����f0���
VV���uG��H����ݛhV�-3EZkDc��:u��w�v�'�rR������:���p�q�_���q㝻G���b`�b��N6Ϧ�x�%^��*�w
��C�6tC<�.R�H���J��o ��c�'HuK�oZ'v�5�?S2���1n��Q��M}D�v��z�5�u.y�*��v�8�#���!���Y����,;�jR�arS[m�~f=������g238�����@�\m�1Z��O)�;���'�����7�i(�ϱO�j㥝5<���dj%8)Y"����_��3 �z�/8��}���S�WS0�+ȩA�'R�O�}���G��!;�#T�m�S
�x�q<����x
�Wc��I���ea9}�<Ӌ�Z}|��^�HÎ�g:������$��/�g3���|�|4����'=4������XG��;X�io���"��������]g�(�x�R��|/�-<kWB��c3BU�n���5�q�L7�����ldG�Ez��3㰁�s:�L�R-���=�O��۞'��TUU���W�.z,�����e�+,C��n���7�֓e�$�}����e��t��](5g�a'n=�;���Q�ꓢ��"�ZS�o�K)H�NKHs�i+|��c~��,�f+ue����)`�c���#Zv�ء?t&��,)T��}L]9���CN���.Ěp;���Vz�z�c�!�F��vT�P�*�X�gTb{q�ܾ���v��HOQ�v�`dѦOj�?��,����[W�_nTj]\�ѣIL�c��a���1�^7`K�w�	�����LXan.�35M������_�-�y(r�$���ZPe�)˃�Z�s��g�N��T�0��Ķ�L�7�	ټ��d�v��u*�`��?8۵=)��s�ϵ�'���������b`�������,���u��B�Tϸ�Ws�!�v.�(VQn�,l���H��z�� �����/[��6���V=	�r��;.���n�~��1#/�XF5����wǄ��%���/�Fw�S��O�8���um5��2�KV�H��H�,.~qÍ.9�"�%qV��oYxP �9�G�s��Q����oH���Ju���8�8�u�La�.��X�1�a�='�{%��A�w#�M��7!�|�n�,���m��y����0�2?��d̺,r�)YIg5�X� X������O���� ^.��@|�*�:��p����	�8&�l��,��(z�iq:���'~�����އ�*A$C?0��Q�3��Ȣ��z�E�� ���Ag��#������#�h��)�m2��FGZC+P��WA(������t�oV�8�g�]tm�s\0a�'.��7|��3v~��9HØS�ү?&�:�	C�#����y%dWFx�[�gH�iy�-���:Y�Y���=�~� ��=�Ps̅���*b�����B�O�}���sY�ÿ�x���&���톱ɚ�z�°]k㷝�sQ��^G6�Uΰ7I���:^A��X~aą5�����,BcU`���<�ޝ^��f�;��t���`��_Aq ����(*w{� �A5��4�(ߥp6�)t�Ғˇ �9��� ��NK[��<�3&ʻ%so׺b�O�:�IuQ�*楹"k�b����L�@ᑑ��s�����s��ՌG�X�<Ǯl��|�.���	u�iy�}[��4F��j�&:���{o�2�^j݇X5ޖ�-&��~>n��JW�vY A�!��_ޞ��f?l��+�S1j�P�V�N�.)��p�a��v7�AV��t����=�ȹ ��ص�����W5P�X����ۉ��9?��s�l�uQ��:=9���k~+��y�8��nyA�:D�-
j~CS��L�9����8���ύ��gu�1ϸ��MٜL��y����I��g�Y��	a���؜�\�t�_�W��9���3������k+���M�zaE�E+���A�<�z����P����)���ڴ~0�:-��x:�K����IJ�[�{窉�ݰ��o�v۳Jq
2�d6e��]�2�?	�#T��G}�-�w�;��(�;�zZ3lG>��<�4��B*��e>���^�����&2��mͳ�>7I�	�W���Ŀ�>50��� N2�;����-���I
�i�<�}�[�I�!��Ҵ������+pr����;�Ahn!�8��Wf4�%�ф1����-`Jzu$�1��Uk��p��%���E�y�٠go<d	��k5�ʿ:����Te�w}!�-4�H��(�q*�״�
�ʈi�ٮ|���w�X�@½��Ex�+ӬB�k���>�c�Fŀl�e���y���<7Z�*E�c"2w�� ���Q�u�j��	?�4C�j.FIn?گ����_��L���I��"�r�3wҷP��Hf{(��H�O����H�}�,��K��¨�7|�5��Žc�z�q�K�G���x*��@��`�pu-�
bB��f�h�]����ߦ�N�n�]*��)�k]8�C�4��p��$;[#�i6:P�/;6.;?���l�W��O�|̺T��������y�E�l�CԲ*�0d��Q�t&�=�=
��~R��Q�l7�X������x��hR����*�qE�*��6?�8vgm����~����f���S������]S�L*�8�II?�Y��>E����$2:�w'��b�;�`F��i�N�����1��(�;(T�;\J=Ԗ|��� k��I�k�z�0E��)��K��n_������� (��y�J�2��a���xj�]u;:�]��D