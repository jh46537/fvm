��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{�.Ѱ�!�C�8f���A?���<zj4<����R� �{a���<�t�q��|l<ч�˸xc+
�f�A	.�hЩX��Z��&���@no~)RxU�A/	���c�b����jW�ߩ�X)�h��	94�8�X�R��,�λ��u��|���c�!�|j�6%r�Ԯ�������R��� ����f�m��w�d��Z�kL1�z�உJ=z|��X�� c]�� ��A9�b�����cx��KU�K���S���:Xuߍ� �\;��N?��N�����,�9���	"�u�U~+�X߿� 4�J�b˫�N&2\�d��Gߵ�YJDR�D�%���rw��j��5�YIJ�x��
�O��r^��:,�$���F��w ���^\ǖ�I��S߃
D�t;�[������dU�P1 ���"��S�˪�-óSAY&�$�����=��ө���
�4��4�+�7�2�#�Q�O�ڭMY��m�+��p/yS�ɴ���c�ݽ�x������5�-����S|zUJ�fFW└d���sg�������`C��?�x��M�V�%\��wq����l����t2dG���}(!Ҷ+��TcX}-Tc��R�w }o8��z<2&8P��#�̀n`|4��v-۰
B�a�g�f�(�_��O}��g0.2��\��}��繞rm�+*�}	��s�_��!>�����|�U���a��M)-V͛�җlg����蔝ݺ�$*�d%�LDb/Ru��Vʚ�iQ_2�����m�J쁳FkI��1!����F�b�g�5����'�h}�^�]T��@� :#/U�ؓ��׳A�j�,3Ѻ�	���N�ؾ���8r�N�b�MI��~x�Rݜ��)�p�,I8�P��*���멭��e�z��J�����h�ZB�����)d8��Y��׫PSq��4K�9\��OK_�m&�[�l��׃�����C�)U�o��b�?܉��xs� Thf��@`#pb�h��E�6d��)�ğ�ē���s�K�7 yH�Gr�[�,�TD0�O)۸ ��K�`H�Ԛ��s��L/�y^{�եJ+�־x�����D�`d0�� 붂Q���N]�_}ø��b�.z�x�lBKйA�T��Sy�[5���@_���gN^�[�y�SÌ^u��--����V�>iu8_�QHi[:YK'�;ZfI!!���F�'��ѳ*#��#������Kq�0�;��1��l���=��}���4aL{N|]qG*"X߫���tI�! Znx���ܲ�	�hyA��f\
�bƩ�?��|㎷'�,
|�4H �/Rp��,C�g��Ʀ�8�a1D2�8U �<�L3N�U�PU�=M��B:��^`j=��D��hX3J; �8}����a��0[�]>,�	0	H�s��(�vT�x�H�H�� �YZJ[v�⍊�A1KL?6�T�j�cD�ܙ*f,/͜܄5�m��K��d��o_t�nM�}TU&��y�7�z󊬍��~�_i��A�V/l���D:���+aE$�X�S�o��w>��.���b��&�r7S���D�Zk7�'�������e};���W�M�G,�jvR�]��@���YU��/S<,t٠Vm��L�:#�

�߷<8-�᚛��D	-��3��I�D���u}�_�~�,�zRt�]{ЭI�=�z2D��5�]�X�v�؟=G y�˃�(�]+�0h���6�5s����;��{;3�uL�<�.� E�Ή�� ��s� _a����"��Fb�%�X�P~�̉&=��0�Ͳ^�&�{��I�@�_����'��c��	�b��n0<9Q��^/�y�_FZ���M�����5E������&`Ux���{�kG�mT�-9"X��h߀"���Rf��T�B,tU-�9)�i���J�H�Y�I�	O�}yo���)�]�^f�F|��t����LXeH\K�����U�p�*��;��N��6h-�R�Oy�jB�L�o����헜�3��D��t�c���.��ICBFD~$r�¿sU��H��lΗ�y�+Ti��(ߕĤb��+�ŸWʧ�V����O]=����Q�G��Z��`��������0ȋ����/�?\l���B����l_=
t-��ˤ�w� �@�EU����1oVZ�+��,wB���=�������=�[a���'M�D�&�����
��97Y����c̤��P�`w�#�`c�{#��W|�L_p���0�*�rt�������PMM�!e�[ �s x?�&��9�|LI��l�s��uH������O���8�.�ٍ���~>ݗg��)�_"c9�-�)�~���/�~ t��R�>���(eY��F89dp�X�|���I���R{��W����&�G��&M.J�I�� =N+�Gb�_q-�*��2�Ջ��̣Gm�9�&}2�Қ#��Bz�_e[2dT�`We�<T3o?E��W��/sئ &(��l�zC�c�5<��ۗZs�}��J7p6x�?[l~�g�im�a^ҬNk ��%�s#��Pw;���2گQ��@!���t�=��m�x*� ����������j��ǪG7�|H�y����U��gk=������3v=s9�!���cY�F�~�����M+~O@ŐɖV�_�sK�m�Q)�S�(сQ�
�Gyzᮥ#��N�_U�S�h��?���Sm2
::���`@jm"��SlC9�ԭ���e�F��z.r�[�l�?�q_��t���Z�T�sz�P�_����W�uF%�$4��\ų�֚DO�J�m ���Y�W׶&T+��5V}e9�Ѹ�>p��W���7׿�ϫjQ�I�r����P�y�hCw�6ER��M�&u���6�Р�"BE�ٽN�&�����k��F�{�� ����fO��?_�=Ѻ9��`��(��`�%K�2e��b.�)��Ip�����VOӸ���W ��2 #�"sh��N֊�O��������EK��oވ%�Y��7�^��"�S=���Tl"�k*��2^����?|	b]�����8`U�td� �tNh�l�Г��ڗ��=j���OkN	̺lO�J�a�H��nѬ��ʎ5��ry��^M��T�Y\%�#�	ܲ������A�j��'X^g{��D�Н6�3
��/ ��AJ^�q9jo�i�H$={H��k��C��(8������n*үγ!Q�����5U���0}���H�,�0*v ����d�R�%���������5�����C�>^���e\�� c8+�fo��.z��ܣ��&�