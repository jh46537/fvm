��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����ő2D�=C[�6-��$�C�š��m�Q6�P�h`{�Rk9�����0�	��X|?���^�r�ܲ��^қ
�j�)��a_�߇X��5���k�W�3K�����6t�R��4�<q�� S>�Tj5M������W˅��ޝ�m��F�WhN��Igj�������řg�4Eo���w$	6��8��0&�f)�;ܜ0]�%����/x+|u IQ%J���`\�~�
�_�n��G��BL��u(�x��$#�D:/�ȯi��@���i���(�, ���]pͿ�%Z|��K�H*���B4(�R�#Z�f�Иx����T����/?��y��3ׁ���	�e���q������O(#ŷ���^�҉�6T_��ĢnpeUG�����p&�$X���� �sj����D�u9,��`6�<����H�~g�K����$�>��f�D���e&���p:���q,�n���<�sCd�k�:-� ��Q�5/��^���vW�:m�3G+M9T\��|m!TFbB�|&k�EŸ�^G6􈟇w�-d ���$]�I���9�N*oKW��)�ykn}�Vh��9P�x,�s`���Y�P� ���
"Eh}�)�g.�؈�5�۶�s߮�NW�aҚ�W9vq%%��x���j�ؓ�����0F�����_��<s��؞E1G��-"�Y?�N��v�`�(E���{��U�}� �o*ؓ�@n�|h�}ބ���7L���{�|���7iqV���4�-&_��%��-MW\�6(my��s�Hw�+�q��T	�7�X����7O[!�����n�k�m1("P��6w�λٖ�̩�����!L�{�"*7�@��߇���S<�"��p����3�S���Z
,�l\,��ܛ����;H�WA9 xq]L�*�v��%>?�v���<t�V^�����q�_�y2�˧b_���f7f����i�e�b��0ߪ�hp���Tn{����L���h�*`~��� 5���Hq��6����S��Nn�Nf��V X��\��)�/u�x8il�����堊�M������Ý��6�ϻ�NE�[�@���N���OR�I���F��K�o:_�0�H9fpx:�b��V�|���G�R��0���Hf��N�U��QuF2#��������1����d?g�ܛv%���9s���2��	`�����q«�W)���8v�:�LV����f�6����W3�1�8�G4��3�G#D�(b�_;�i���	5m�6V'fTt�U�	�O��w�/	�&��y���:k+��m�o�=�~�����3v��N]s�wD3�'k�1y�_�/��3�p�o�������LN� /CR6Y"�=jAk� �E[���_��Fm}�A����ȗ�lAz}���(���(�V��v���%��K��I��k�5��uoU�W��,�
��k�`�"�-M����h8I~����Ju>Ϯ�"OL�K�ޤ$g�א�-ot��������'���Vu��*��Ė*�Por��JY�v�j�
[�ȷ�d
���M��_��zd7��E�=�y��<;�g��V_}=fB,��0o�xX:ۼ�D���IY�Y�N����߄Ѩ��n�0�Ko2��_�ETZ����V~y�>�s����A?k������@^u�r?A�iߣ�V����>$�2�jy�,�%��O`0��)
��� ���(�Y�݋�M�M��,����*�0u�^ap�-W)C7�
���-�nK�I^Ժ]���&Vp��1���ׇMiǗc!��eK=~y�z
>�*.�2���͢njIoĎO���r��di����%�e��.u�dB�ǝ��dj�4��=�o����v����;�C����r�NI;3�|���
�x�cF�5g���}i�YcB�&�! ��;��Y� �\>���F:$;�՚ۋ�~^pH�)ǱNۊtLq>�7M%�^���7h�k>[N� �x��bCѮ	�HJ�3�@���}M�C�	�ي��*�F�aV-�c�@���A4�<�P-�Erpmղ�1�FN,6�Vk6�;r9K�T���j(�����7l�O/e�V���?=����W�#]@b�y}����/"�Ɛ^uh��'R�\�K�ۦ��/I1�~�Ԇ�c�PgJ��Uv�R��u��_���&�'Um��M9�z�+���p�O`��Z��N�I�ձh�u�`t�z���|��V����4{�BQ��P��j�{~R�Z�ZW�� Y�� �=F;|����r�} ���V_��6`��Ѯg�B!<����6��(�/�W�*<��x��o��q�OK�s��7UJiP4�G}�^)(��+��P{��Mk��G�d�Q��\n`c���=&�:����+��}��s��W�M�߾msھ��c�\H�H*X�XR8��AsnZ :n���h��V��;]�;��4� ����R�)�����=�?��:�H�������-"�3Ш�� 2&)Q���S[�������_)���
ub'S�Cf��,9����t��MF�%�"��a�,���H�I����c����:NcT�RLQ�Vz���H���ݟZ��uW��:f�u��=�\l�������>�=������ږ^�S-W?�y�t�0�!/��m�Ar�~HY�����"������g�\�V��o1Gy�l��d�v]��e=�Y��D�uw��#<+���rc-3�,�j��sΖɎ�n$�+�����p%��Io1x1hF!۲bf�$���h+�k�~c�d�˕���)H���0{ �������c��<�� ��qx~3!�;Z˦�f|���&0�'�I0ȑ��������������P�
��u#8��+���]&I3Y:�.���21UP;~DI�cc��I�bp�L1=�lUK���>��K�[	���#
r��i�{���h\8�d��;%���P9Ƅ>���PhK���<��x[�Аr�hA|�dTZfC��S�JL�#�IY��e�_�H��%D�`�NO߫�?hs#�i[�9�晨�-�/��>��]	��&�Fܝ�"��72��Gۛ��+U	��ٝ����h&�\�� �����<O���&wj$j^Ex� �>Cԃf7��=�n�
	��-�X�䄻4	�U����(���E���q��� ���΋���=��X��݅nҩļT?&o}�,k������%@,�~9�k��T*أBS�!_�$����{�zK���Sn|�W4���iQ>?�5]���H��O�/�<��b�פ&�=��}�νd��8S"Q�6ȼ�=�ջ�{
��#�:�I��#˷!�7���'�������X����;���2�h/ŵ9�4��������w��E/����A�K [��ǴY�Lo[$���柢!X���/��PLdȵ�������y�h�QaXj-���~�0_p�ҹ���k@'�bq����H��R�Wv�
�����N?*W�}A�ǯ��������U���z$�NXH������!�.����im�Ziφ�݁�d�7j�>�Y��f�k�h$cQ�b2�LG�l�G�s��A;/��ǬPb0�㉱p���@�{��
pĝ�Co�L0�������o�8IM�N&�ݺ5؄# �e{�r_����>M`�䳒�,-k4�������!�Q����00�]	?V��pya(!�i�p�Ŋf\���Db['Omc�Y��1E�����f*����Ѧ����LFX^�G���"a|�aԳm�Ύ��y�׎�%.�)��ٚby���� D�i�o��Mj�!����}-:j���c��|���Hl�>�4Yò�p=Ot�<�1�wQ��1�'4'��R6��t���� Q� �m8&�f�@�*�Ix^V��%��BH���N�;\�"�c�c��f&z=��7kj����&�Fo�}���qȒ��'x:��^C��Zz+��[�܃~b�S�s�f:F.U<���7��1v*�M�e����-"[]���
u��T!��͝99������#�55��9�!+�#���󩚒:�+Yu�t8�:�'2�6
}�t��|�����*"V���/�eu�w�/��@� �{Y��7f�o@�v
٬���|B�W4g�^b�w�Yh�`*��{f����W6�g�";O�d���)棚�8�0��u�Z�|���Hgh�Y�� R�t�_fdf�ě}��I��{U�&D3#�n��1�?�>�h��e\�R�o��kٸ�YAD�aG[�E��6�v�