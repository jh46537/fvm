��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��V-�@m��Yx�W����'�4v0΀�A���^���*�u�I�\y#ȵ@N��u�q��m�XD3]�,{��_j���_�<���,w����i�{��z����o�ʷ��a��c�ڏ���J_�25R��c��+u+��P2fD��H�=Wg	qgB�H:�8��4:��0� ��x���cDoߍ0z��M|�:�3�; D,���Ͽ�0���`�Y]�F�
:	_���VSL�]G�r�N5�VT�	f�ޮ4�=2ٳ���K;5�8����k*.�tT�5����j//�F��HfcHg��IGd�?��L�12���P��U%���J�3�[�{�l+}��
v�X�� [�	Oߧ^�?��]�R�Rĺ:Rc�{u������g�'T�ew�&��)>�?���Y6N<�Bhj�z.���TQ[�Rj]&8Z�˟�$��D�`NLg�Ħ���"h��hg�E�#/Ţ�M#�F܆��,�+�r#�P�3Hy��n�
S��<���mLs%��?g����C��$���bbn���+��舔���*�����&xT����U�����4 �o�lJ�}�d�@-��~��|qo�Ϻ��Rb����f�lTw_�F(|��y�jx�y鋥���5���z��E>�L�@��N��`���(6�J���zl�rH�-ج��(�������C��C�a٥{FF	�DH��e��;�0���x�7�v+p��O�N<{�������=���oK7ri�*е�"Ձ�S�n`�R~���b���v�Lu)�o�Z����	�ѻ-��8t�µGB7;� �ȏ�`�K'�M�F�5/_�ctȩْ�ʧ8"\1Q`*��4�:3�gG*h��@g�%K��a�K���6��Ook�{�9�mIw����C�B.m�o�|��%&��[���MR7�mMǪ�m�_K~��a�ۍ� g#�Gz(
�J����6Y��W�H�X��r�+\j	2HU��K�,]�0v2�;���9��^7]O�x�U߅���p��Z&a?$��c�*nK��5�j�� $��6��p��� ���f��Ζ��N�w�*��tA�Y��NH�@�v."�'V��y��%��Râ� �/c4v��"O7W�kwz?��I.$�va�TEh.!�-X��q��v�*����=��-?�-�2�Ԋ��g�W� Z)SH�� <��V �y�BJz2�@Z��
�����oA�wi�f�l����ɕ�����	(HG�t�1��9�ꈀ{ a�+ZV0��m�����S3�M7:����J��6���(�� u�"G/~�U����>	�_;���_�g� x�q���]1 �38>e��~Q�Z㛮`�)+-����-��A�.�&��rH��r�H�,���n�ط�u�ܘ�8+��J��n�Fx���0~'ǓV��)pޫZ'��WV���`l4D)zw�i�H��d��$�N�6U����nlN�q�[��28�^-ol�8jV�Z��e^�[(�л�g7e����@[�Q2
y���B��ß�[s�R���z��l`��w/��A^B9v1��PI�2��m����,�9�I'�SF粚�K|ǹ���#D%�ݙ
I]�J��%����C����u�<�o�Y��(*��;�٪+:�U��s��HH�xf��P�َ7q����^���p����TGLP�mGPz:���,�[���W����б��e����+l�|����*:;��a;y������ �Q5��tg�tڴ���[.~�A��gEc��el/�e��Md�ʀb r��4y������)�?yl�}��&���8��Ӝ>+�?�����\>m2R��-y�'�C��v��J��}^�U�/�C�|k�T��Q+������+)���;T�p;2���k�&���=��]ja��RP���cv���!��X+V��>��*�YtS�1�.��3X�O��N뵍K�Ke������r��(�`�D3�eGA���[,r֔��� \�GFi��]J},�w9ؙ�<j�tˀ-J����i�1��>q�"���Ա��H~��k1<�R����H�5ˠ�
W��j$67���.��"�Ս�����.s!p�r�x������,V��>^�B�60��x�|���.���1]��舆�͓��" 3�w���������ҵS}/ɇ�â��X�e�[Tĩ��/��6~M/) ��X\}ad���ܔ���rX�!0&��&þ#-�g�*�Y�|,���}%���	0��Ӳ[v����[�V?�Ŋ�d����ɥ���Fe��ZQ3wIN����� �!���J(���%킧���@ѫg���T��	 o���<�5���5�V�(�8����:�Fjo��c�a�9���(�,��ݡ�f�
����Wl�Um�C{�-P�����4t���&�H0�(qՍq��'#m����:kx]V�(43z��l����@�[A�$����P�վ�T�Nt�gO���F�L��|�4	s����Y����-�L��?.�����T�(����s '?���yJ�d������m��qG�D1��h���[ ����˭�a����צ���|��4E/v�ՈJ� ��c{o�eh��Q�sE&V���'w$�E�10/#|<$.���<�k�w��!�D����z?i�_ ��|�
��l�� ��!`��!(c��ȱe]Wq��#��%b��X�S^Km�K�,1�1�}�~x�>�t�(m ��p�����:61v6�!N��a+P�:X>>}��m@IP k�0%��š��U)���9�Q���'kv�Yw/r�TQ�,RXaMc�^�H)��i��ظD�9���!Z��b1t�pU$ !����φ=8"}i��7�>�^b)�0��Xm$5�T����H���X����>��*����&���1 {T��r��0�F��lY$eU��[[�?]ǂgA\?�ٝWٝh0���h���{&$�X�jrS�q�B��U�&�z�4C�sszT��3�\��t���cg�^��]J�`�@�P߉��lg&Hf��4����8��mo���K�Nd�)�fL�E���9�����Ϫ
��m�E�����C>g���[�"�h\��������vy�ƣ��q���MS�F�5�3�E}�����f6�N�9�$pBE~�'I��q~�\n���˯rg�@��.�E*
�f��<j�BH�@��v����3��z�J	�-�]�>I�g�
A�ӣ��dN^m�6x�hnLwz��tӻuE����� ��G�bs�f����O�]�l����1R��,뺣���MYX��O���I(�e1A^������!�^KȘW��W~����D_�CB�]I�h˿���Y�/�&�"D�.���5�n�4(�X\n�vl�\����������2���	?�+F�q��6���Hw��v��!q�PQ����nw���cec!�������.u���b���ڬ�HS�rA�0��!����I�A�O�(��/��jAK<Pu�c��m���5�g��%K�I�)�9�p�鐏�CEdg�X	�ub��E,��L>k���8U���̼K��9q�lc��.����A����nA�
�o��߱���(	�z&��+�xM��d��8D�>a�/Du��������C8���ҫy�������p��q�Gh��>���N�8o[Le*Y
�XϜ៊����T�;�Q����J��sF���*�A�eo>N99�V0W"ff���i��˯K3[�L�>��]�U���� ���w^����Q�ɪs#�oE�z߆�i�ln����0!h'�5����`����:sAЯ'��)�C	�������Ҙ!~�C���]����V�ձ�����>�_��N��o�p�Y�e�,�t�y����ZLK1ރ�����S�e��ޕۂT�j�,�H?eU�H�I�.�=��xL���b��l@wtia�`�oB�	̨oD��ة<�.�������O
}�#T�q����$����+{�:����[^ #5d���ƘT��Duc̐�>�jx���R�g�ʹ��l�*1���ث"��k�NA9�)U^9�j@�2��o�������$)O]۰B� c}�HSi��ܻ��2&��_s�Ϡ�:�P�1x��ϋ.�����>f�n�w � c[��ǱK�W��#�B�
�M��x ��A���L6bs}������>�##���A��W>��3����(����`J��]M�7�D�I�uIڡ? �
^��.�o�|��ZCC��1���k���6֎B��2v��1��!>i���V�»J�xAk��]u��f�L��6�����k*{e	�ױIWv�	��ʼ
wn��e.y<���kX~x/�S�T��*#��b�ֆ�ł������%I���0`=IK}f�x�#�R�"ѩ2����.M����7�`�<Ni���`cD�a����q��Z��2J/�ˣ'
0��(�{��/	��`���kp��Б��"�Pn��&�-�]��Ӥ��tă��,�36����'��$�!C�f�B3��]�
cZ���F��B
,�Bv��� oE�e�<@��R��6"��ΔWѧ�Ck����r�dY���;�i/F^���ư�O����{��W�d*/��\HuD^�6�40�F)E&�����K���[&�� �Θ��G����9-ۀ\��7�'�t@��f<Ů�4��B�A�vN����1�l��n�;�	�m�D5 r��O��bܷ�xւ���A�PM�C��Y��C��f�#6��;�㖥��l�Ō�y��	�"8��8��-c{!���Hl�,�� ރ)��H][1��XB�oS�\6D?Q���bTU����k���;�aWb���C��Aa&�)9��֚��Ew]&�/��i=I���R12L�B���Y��	��Sm�-C�	M��R�y"�oܺ�@Z���'}�,c��s�H�M����Q���1���N�O���O�P
Æn0\���ӱk����T�^dh��u�[�K~�qQ�%�-����xYդ7�%���j�iT�~-��a�� ���g�^y��<h�س~���i�)'1=H�|�i�'��T�E,�V$��?/:Oe�{�3LDU�s*�b�G��XU;k��X{2AL��3Ͽ�ʒ;�mç��S&��}�t��O��9���Z.���ˋ��Y�*s�>�Ö�4*@�[ᩚXd��f�'l]��V앆4�A�s�D�NN$�:�<�f_��]�8I�$8�^���q���qNL���}�Z�1R��k�d�I�И,�G�Gd-`f��&�uK��O���e���GI�.cXz�7$]��%�_9��-Js���]��z��]s�\_�YW`�J9x�(�~5�A���XꞼ*E9M̄z_s%L�Ku3����A@m��'�6�
�cnՋ:"�[�)�zW=7+� H$�$J �WÅ�����N�L��?ܬ{��8��%����O�����.�km���^�8�NI�ýXG�!G*G$w4�+��a,�@5`���w��HY�?����d�@
��a�^��«�r��>� �0��pp���x����^�9w�Svpy���	m`�s�͖I��? F,x��\��kt�i'���E�fC*˄*�[���V��ڭW�8�8�l`��j��rL�N�금ȁ��~a�bZL�':�������)��@�MC
�dB*d�c���4粶�)�Xz��_��u�rS����8��;5�̝���9�=%x�[3ks��w����&£>x�0DŰ4� ڒ�eN������A����&sfQ�)�WV����fE�u�Vc_ED�4����٣�A���V�c��\)=�N��֐���e��F���t��)�6 ��ϝTWJ�WΎ+%vS��ұW:��,6���V;,�Ekq�����GַE�mN]P�^	~o��ZlB�ZY�aGQ����I^o��s���?��:+�������V�j�4iN5�1;`�%���3� �H	���8���	-X�[�����N����M�V��<��J�Q����f��Դ��M�Q�
�ƿ��ݖ�3u�FKGAfU��k���@Q� �=��	πJd���.'�=�W/�����U�)�F�[_i�� $��lxqxl2U�H��(�,�$g��8��ò'י^h4�4ޚ�Z�#/���\SKp���)��-n���ԁ��.��&�E�E�Ǔ��,&�iP�Xl�7ί�P��֕�X��.zڟXz�^��O�сN~wd!���������j-q&BL4� ����x��lQط0���gQݳ,�&��C����JZ��a�j~C�}�l}v�ə]�b���;܄'��qH&HR!9fY�����rC������Nj�)y��*�����Coe�t�'!L��@	��1y(d$�1�Xn�Y�e8�?hg��c�E��"E�b��	�^�m���q�qg����r�L��������e�5�~~\���\#�F7�8�?��K}a,ՙ|�QP���6���s>dQ�'�ے����=�I���c�|��ck�