��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9���!���s ��o\y\�-=.ɖ44V����G���(XjK��K�ךR�é(�>�Д��ڳ�ZA3�G��[ʛ�= ��"�
0��c^��ˤ2ed	:Nd�@h����[w}����ڷ�W.�.�ZWݝ�eRe8�^X���vԟ;y��y����.y9�0���<��i2����e��� �d��7�\d�V�4@8���CB��8�^NM���
Z=e��w���e��,���ր�m}�wA�P�п��sIj>��;�r�n�F�>5�����׼��7 A��}�I���8,"�?߽)��q(�yK�6k��gv{=�0�.��3�f��>��l˦�� C����b�^�qS��� ��Iwq�-���4�!��>M���Rɾ+Y$�z����>�a�YZ^�#��U;)��D�\�'����%���Um�x�Dֺ��^@pۻ�Ĥ�22Z�D!%��E�Tq��W��G_���~I�Q�Y�J,�N��7F�gQك�BI!�c�a�a7.��ā!�{C���W��ge��u	m���A��%3D#B޿:��޾��~\:+��1�X���pF<5��2�U�u1ړl?<�+��5���Sy�`5�����L�x�	�*B0��̘�:"�L�Ɂa���{v��8�_��D$�"G�v����j0dȆ��G7��/H����3@��K��\�)��fy�t�g����\��'R�F����ud��sV�ۗ��ϑ��Z:����P�x�:��E���V#����l�	y]����JM6Py���R�'(׬��6d@e@(BÎSl�Z�ԯ�D�>7�'7�՟G�ڝZ5^�"=�шś����W���al��C����R^�y�>��C&�uR9�J9��;���ߨ����vN� �q���N��Xռ@�U$�tX�xmԛ�>�����|�Aެs�����e �0�B�	���7�����X��ȇX@n�&q���U-�̀H��A*j�)�D.�/�P��PT5��p�{�!%0�' ��)H�L�L��QX��Va�-���:Q��x�>��L��r/�V�������(�q�X,�6������C�ew� (��"x�?�e�L�-�tD9����>�\ͮ7�N^v��F4�p��xVUUs�`��
6���f��=kDH;�07D�m��c˗w�䥻�u�e�EG�r��@	[>]C��OEs�t�"Cwjm�u}E���Ŗnʉj�����ML�mZ�M�q�����u��6���nW���8�
O|:�-Zg���7_F���׷@������ �{Ӝ�>`�5<�����v�',]�F01���b3��H�����	���р������Ti� -�z������"��_�t��\�i����e�p�[�!kT�R���Mpw�D�9�hJj�s�����*��s{A(��"1�H�Qr�ɺux�5��hfY�%/���.�;��=�ም���(i��r`wo�=L��9�kF(I-����%�e�����ጱv��;��iI�=?��}r��/��vB&�-*5�ȕ�q6 ����f�d��f��j�*�+�K=,�nP�%�p�2K�;g�Q�~�&PD����j���b�oic�|פꋢ�$�^1$"|��<W0^mAI�G��%PE�m��7ղ���M[?P+�73�o�p���R���)+Ӕ4m�f�L�Qă�� 	��Ýۊ'.v3+�iM��p��HW�;g`�XPLO���l������糭�0b���d���-V����)o��Ҿ�d�{<����yv$�U�����K��g?F2���ѻ]^-�
/���E7��^p6��!@����&f:I.��=�M�R���B��q��`ꀴ\�,r�>x�S���o�&5�6�bVO�Æ��TW���������㿋�)Q��bh�ǼO���k+CcAFL����r���:־-QS`]R��CZ7�q�6a�&�6Z��<�V�J�f�Ӌ˗e;+=o�6Y�8@�j;�è��;�Sm��%#Րg�\5J�B�7�Y��1Ι��n�Fs��4Z��,3Wj����2#�z>��G��x�(�}<��#��+�r��;ݙ9b���f��Y�U���Q �<> ;�7R���ͺ��v��~?��^��ռ�J]�$�a_��e�,gn�a��6��n����l�<K��PR,��k�(^�J*��hx�����ś���2o��'�S��m 1�A�8>�š�7:u�H�AT]`?g������ڕNT��`*��O.��Bs h:�����%\#�+���K���|e".u�]u�b5����0�u�$/ۨ�Tm�ݐ�|{�.�>c5���S��qt	)0�J/*\,p�G��y0�6����Ʋ&�R�]�}���o v8����x>���8�r}�D}X�5L��;�(cZ'�HZ�U�Wz�>-�>��F��V�G�������yp���5�C�h|h��G���_��5(�R�[�� Q�p��4��ro�����q%�-Z�֪o�z)���w_0Љ4ʑ��f��F��{[�?�W�0��#��@��!v�(�N�+����vH�7�ޱ�I��Ӱ�s��A"�-�
�/��8?-�b.��4��ock7���#�4PZ8�13���܈��GXn��?�ܦ�\�H��%�a�
Z��	 j��3z�t˃���ɠ�h�쭙Y,S��`��XQ��߳��:̎<c�V�`�>~+����	�Tc:�I��`Pvw�7��H6����}sEm����\���i��`���H/A�{��#zQ�$��I6�5�jc��|�TA�Q���xA���,8[�3��l���Ө���8:�=7�����<�����N�H##���	u�gI�ҋ�b@_���r�^�(�;�F�L��x����/�t����d�Sz��t�PPp�|E�T�Z�gZBnf7 �d�F"(:-�� �]P1���8�!�D@�5����T��FDf�p��=�_�k�y�\����a{کn��U��%`4�j��D��mP��H*Q��M����� {O;�2NN| f�)Q�4�y���R���|c�d�'�� ��0�r��M�Nz	��
�	���q���	5���M7�ff	`�O���q~?�z�e!��.Xj�'/��ρ)6)��z�q?%m{g�\�Z�_���,�m.�4�G�}����TO,Tn�[���!���4��,�~�(�Nv�164���)��e�� �1���Jl�6,g���d�8Z84�>1��T��<M����{c!��6g\HW�߿�1a?ڃ_0��RO��,
�e�dn��z )�,��I����l��c��s��bI�u�Hv�;���UCJ��0`�l�Y����/��;g�%��VDx�E�i�m�K��"��5���εu�aA㱛l2	�����o���/��M>ԓ�``s�FتT�sg�<<Cp�<���>zk<�D#��r����Ο���?�e-~\IB��:3�.��;l�e��&��rd>� ��ڍ�4(��O�BB=X��˧k�!��$ 2f]���jȪ� ��U�@��{R���yiA��dmj����~�:6x��ǐi�_����9�<�������%'��thi[.�e�`V@�H�ko���Β��k��F����$�g���Z���ľ����RO�*��9k��4Q�#�󕝢F�VVӋ7:�7y��K�����i� �.U�h�'�m� �YxM�&��J�Ez��0������nE�3��P����E�k��#�S�����Kn)����$+/Ǡ��2����|!�ˋ��W&�i��G�]��aX�����U�z�I���}[���W+�F�	ql��q¨�Z�:����?.SP�l�vo�=Lp<G.�s!)ЁI@������ݓ2!�v�%+�{��U��)����x��a�y.K���G6'tK᭴�&I��hz��p+��M�p��6m��/g��eƯ�ɐ�����b��:Li�|#�W���w�lܹ���u���dBN���h0��d��5�wYe�<?O����G7��a�;�H��1Ȅ+R)2�����h�/��{�|��u�2��ì)?��k�P@Gxg�K�k�X*����>xq涄h�l�e>��B�"�,��7��/���my�Z�A@�la�y�t�zBMN8q�H%���TP^���_�D]�+[I�Se�\�ci���'aeK�PB(%�����M���Ӫ��%��*#,n��OP/��j�q|�=��<>��ʉ8��^U�>@υ����J���W���&�����jO�X���	����HwܤK�3��yg���T��
�O�Ԟ�{l"g�����.�}��63'�~6^��-���Kj�ػ�6ym_4�U��F��9�
S=���|�PH̎�ro�/���e�)�N�m�W��V� ���B�(�j^�"��K� ���S���M"��2����O�dr�LpC9?����F.W�h�h�E?���&�U^�n�_{�P-�-�Øy����&�Ϩ5t��3�vZ�X]��e똍>f�WL�Mޅ�7~�߂����W�j�C� �0.� �	��/�]�e�J4�R
�b/�xݵ�=��
�b��MԘ�_ �/X�5��韌/"�����\�R��/�i2u˕~��(�óK\`������M��&I.ܶ!�OH�l����6j����A)v�<��@���b��X<!�5ڽ'P;�1{'���i��+��B�Ee�($��~����H_�X�%��;�i$y�l��ChY��y&kx��.�u�Ji����=�����9yNŔ
�P\��EYB}�S��	9�C¼-�S�n�g�Rq���hC�����3дS�ܹ��Yy�^�1�O,��9�͏���8��\wːd^		����� ���՗�n)�9����e�`�v�3��C�O�3w'����L��q��W�eK�s��W���vsiA�?0!�g�!�V��n�/��RZ�����m� ���];3&�3�ϒpFl`�W��7"�|C��תW*j���M&�P��$�������^u�e�Q*[�$��������2��Uy���K����E������� -4�q��G�W�w�Y�S�`/������U��{�*�	,���|�G���|��g�P��j�|(�����M��e0ơȬz��GL�^����j��/����<LS�����T Js�6��|��'+�D��$�*���)<'�Pk�����qd#���h��-�M��.��[��@��+�]�L�hp�<������:ï�,2{!Cۡ�+9�ܣ���%�4�y#u��b�� ��9�8�hmt�j�Ԝ�>�İ���0�!���$��H�/!����D��wQaW�8�z�Qx��x�������8qN����r���