��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>��������ّ$�*X`F~�������><06�L���\�D>�WҎ�����r�.~O�I�V�X;w�G��ts��K�5���t�7��R��пr�.r���x{��}sbeq�XG|7 ��$�ڳ&�e
�=r�$��!錋"���ۆ[�8����lr���8Yi��9���eIE�(Z�)��VJ�j��?~�	��c��R�6���/�WC*��B�����-~��R���$=��&����O6�F�~gh��\P:�w�o"Z��{��ܪ-|$�EA���ٔ:�_JFJJ��S�B	*.�a�ꇔ�@�/~�WC(���&q����?��V~��A������(}�b	ѝu�%k!gŝ>�I8�s)�u{��>kp�Syʰ+�� 2����=��D~0.i4��SJ~��U�h��ERc;��@�p&)Aǳ)��� hU�`��ߨ��a�r��_x�gU���$Esb3A�_��_9��dũ)d�)�2|�>hӘ���s���M'���ϩ;���,��R�)����tQ�W`xY�2�*S+:�#w)X��5�N������қ�Ӱ.P�`���PdnE���R}�>)��7�K��i����#�CbeRC=��%����V������w��2���sh�=�F��q楕���7�
?"�������Bx�����쁁���N�q��A�.ƫ�ҥh�Emj|�3�#�8xuT΅8�(�d�&���:���[�J]!�Y��<J8-/�J5Ü
����Ǻx�x%8��Wy�X�����g�Z�)��{0IX���{(���}����dq�폠����"d<�"���m=�>ų^�'���m���eY�P��tj���絣<"�ĂK��2�e����j�>��^`�M%B��½v��Đ*R�;�����yF��˻@mg�L�gF��|��v,ɔ,w=y҇���>l{~m�-L:���D�@��3�tn2�DA�z��y���1y�,Z�t�\`����ԛ�9����)�21�z��Ќ���@K_%6'���-�6�����!���$ez��Z�]��%�B�d%�_@��;˻6WaxXA�/Z��蛺��Ik�����D�7��"���B�����Ⱥ5vCV���Т�U�|��e,��i,"�di��L6XT�a����t�9nNu
x4�c6�r���ΚE��>/o�t�˨3~ħ[>������S&W1��М$!���t����3�7
�.��d)uIg�f��~�_�t�*�K�	����r\3<{�.��,�����1�����k��v��ۤ��/d����f.�Z�Q�6yx1?�IѬ��[�^��7��g]��������)�O�
����"P�4����d��WŇ�)�9S�!�A���T+��
' �-a���1�N�O�ׅҷ(���֢k4	���`l͞*�܁���<�nC����|���sL�A�e�H�}1�����d��$�
�_��x�$�� �C0&,�"�e��$ -���K�����e#�{.����\��NC�����em�х=�`�#�XM�Q���t�"#�
�Pe8�b�A$����	��ǍH�F���t�4~㈵�ž'�M,\��JD����|Ȍ���OE�~��:�������ba�����jjM+O�Xo1lM9�	x���Cޒ�����n+'{�WS�!N�:˵��-kX��~�Ϻ.>���ጙY�Q�U�r�(�T�/ߪ#=bPů�eS,-�OYO��W����9d���(�&u�y2�F����ô5�����m��D�y�.O��*Cb��6G���ᣍ�ς�Y+0�g�x�)�y�HTiG��b*��4��}g�sW^�j*�"H()6���}�>vOI���{@D��D� СC0�&o���]C|����ۄ<Ɵ
2p����?��Up�	���b�L������/�ؖ�9ktj��	��9FJ�,�E �bm@����n5Q��P���Nx�� �ψ��������ܯ]j��B���s?W[YK燂@�����d�$�L� /����7|�YZ:�+uҤ�F��<�(�n�$��d��j��%ƅ~�ڻS�WJ��	(n��Bҧ�F��t �����[���&$Z �4ƹ̼L����Q�>��ɏ���h��.�-�s���s���fLU�W4�)\"�V>����vN��_UZ�0�[���{�N�~�������MQܔ�4G>x�t�/}�.lA���g-g7 ±�].Jt�`Pb�G�����_��RZ`�|���5�t��ymL6<`Ө�������z ��CkJ�ِ�����������+K���Qo�5w��|���'2��qSϾO��.л98W�N�$��:�C!�sq*D�S��D�	���8@��`	�� �|ف18q�W�D�j.>2�y(����$|�;ۘw�a��V����^��>�Y�NC�S�u���ҢSu��K�%��P��d)�!�L�҈r�4�p"�K��4ƴq)���I�d	��KߤW��H���H�k��㛉�Bud�5��N�t���g�f`e\���ꢦ�'
M�|����n�i-��}$�V��v�ajC�\�#��B>����1�%.��T���-�wGB�����Zj�|�����3?��r[Yj��S4�8�Qc�xw�5J�a�Ƴw���ǋ��r[�$0��R=%ZR�Ɓ��ˣ��&�0wf��\��_*(?>>��D���<�i��a���i�?����L,o��T+SQw��>6���,��\�6��7�;=��[���)����H��c����X{���G�b6�ܭ������,�n��6�����-�QY�����*� W��w���A�j�6	:O�[!��\N�v#"�{�s�]�t��x��Y&P aIBe,|r7% ���>qx��Wo�B~���?g��}�%�w�v��V��@�Y��&1�(ܝw*������.>�Yr���m�R�:�z)+�C�,?;�?<)O���%�����p���1��(��:H�ah�;���ri�,���j�VM��K)��I��1���^��'W0RsH�*��3�ã�5��a�<�@��nc0[����e2���-��p�=`5f��s���w�Τļ�~%D�X��6�0��c�`'o�;���3+=��'[�6i�j�Mhh�wǿؠ)�֝>튇��8)f�P�:�m;���q��1Z��)���.a8x�J��h��~1��]q�3�/n�\a��Fq��V�iɸ�V�2U�i+���6Aw��H�M�>��d��52!��o�&��F�}�8��r��C	�'���4~cLO��:��	�쀸R��Q��;������s4(k�(b��c�H5}z�L!�d䑿r�L��-^�H��H�I�6��W/��)ŉ�J!�������.�M����tX}�p�$�w<��&m���� o;��Z�z���`pE ���&W�y��ի�����"B�s��,��E@� l%���Ļ%5�|�p��sqU��T�M@׶+����?�؂��1��^2(��Oqj���h�J7!��${����Ȑ-�v�ȴ~|E��|���)'ۯ�p�K��Mo�,IAvf3K�z�&i�ȹ'G�-��E[Unm�J�l��� }5�j�y���0e}NZ��h�ά��{^b<|��x�{�7��7�,u�m�h�gG��K� ��z=�\5+Ɲ#4A�s/ľX�Α&}UY��Dz��X�mƼ�I��^��f~�' /�.>/�#^H������'���T�Ì��~�ĬRaL�.�	��	�pp#��\Wh����:;c55���7Smx�}J+\cZ��dA�t��k�:*�Ռ"����V:�b�qQ��R��y򥏃���?��o�K�MH�����\�ԚS�=�����[}b�o0>�Np��f&�*��X��8�$��~���M�Ő�`���] ��y��4z��-"�؟o"m5:��M��<}�@�[=|���jY�ǫ����/�؍W����n�Λ���oC��#狷 Q�X�������S���`��?�-u݌��y���rzM()��x�j��N���+_���Mݼ� U!&m��".G%�YȚ�� f��z�3��o�xZ���K<}[G�j'�J���o�����WrJ�!�D;L�&'<�O�=3���-e_*t�m��:o���	���iɃ�>�00F� ��74�"��٠���kF�Ē$w@��1K��E.����� ��ܫi�_u���ݤ4�����ǚ�s�ј��B���U��&��ǥ��Z�d��}�W��Qdi5�� sc�7P*&F�����r?�'�[�HB�Ft(���������@s
�{�3�2�p����v�Lnm�q:�" �/��K���J?F�I�g\�B0����/��D�sW��ꚩ��ȸ� R��(+Ѭ-�{�π����w4.a���!�v�W�^��;KB֯�脈�Pb���<��'Lyc�uN 'w���'�B��u����>��� ���YWK�df��������4�x�������(l�	{i�f���~�����C^�~��$v�Z��'g�C+�fM诊o*#!T[�Ys��#�1ٟ,L�Ϟ��ko�g���b�!��:`�:vN���,���<�� 3�h!yI�R���E�[9)��c$������6�6,�~� �!	�\v�P�ZKT	z��25�()O��~��d ��9MɃŲl�����Kf�dJ�γ��������M�m���k��  ��j^��m�@k��D���u�L�w);&N8#�+M�!p��')Q�k��su�[�f�3j�j'�W��94��;SS%!r���k��e"�Dw��7.:�թT����.�X?�:.Y�Ţ 8+f��٨J\b�>Ә3�*�a��XnxNV�M�^[��TU@���?��N����=��� �M���sa�b��K�o<h��U�e���-x��즦y��~HĤ0��#����8hl��1���/���@d!�Hk�T�-H0�
YZ�iG*�}ux|���]}�ܢ�>��b3��b��y�+dU��[0��{ٓ���;��8�E���˭_\���>-�%}�p����󤐼��Hם����T��C��_�SH��j�7|�W��E����Θ`��\��7j�C��;�.�'\
E��~$^F�[{���8���A��t�*���?|.��~�y��cj��d�L�c=��j�2�*�oW н�{o`� ���mlsZh"���[$��{�	iD4��ޜ~�UM�H�z\�Xf�X� �nB*:������L�ALt2d.���Ͳ[)SFiG�~�����/#2��F�^��.��R�0-�A���I�g�k�d��\���^���kk���+�";m���t��"$�8�g�Z�5���
У�`�R��쟃�Kb5~!�(�"��-R��8�k�᝼�o�f��J�d�P>C����0�]����s��]�{J���+�0����*�j��N��$e|lj�6���p��R��B�C�5���?9��P�T=�|���ޗ}����]O!��!]��]�٣ܟ��������r�BY�������o1�`�V
��i_ho�Q��+��r�	�'m�3\����\�X��X�8[h��X,;��c�ھ����}�����"���ғ���"|�Ț0��L��m:̫M���}Fy���(W�@�MF��L�����_ѣt�5�.;�Y�{2��l�>�N��?�.��,Gt�����=����;��34:�)�/G���疴�:q(?�����혣��3���8�IU8�!rW�%!�"�9m���̞ݶ���a�_��Wn��;��M�F�2i��A|�C�EA��������t�Z>n��S�:V�|,|i��s�ϛ��i}PA����C�/��`�J�Վ3��u����j�r�[A��j!�o�#�0�(��N��h�eGµ�D��j7W��D���+�r�41'�5d����qǡ��'T$�,o
DB�;$�	Wwi�B"�z�f�������h�6��b�����]�$X-b̋U6����[\q�X 3"D�%�U�ҋ�H;������k��B9��V���'k�l�"��&�q�>���J��;E9x6�8k���F��<rSB���)�K�O@܋��O9�a�~K�g,�z��j���,���mJ���x���J��ԑ�5�o�)��p[��/����$e_����!�Et;N+�V����x
d�> ��^ ����t~��T�2l�������i�'.H�U��=
�h������_�Q�j���­��	M9���
�i#�&+��Wh��X�pui�E�"i ����Eps*�0=�Z~*���J9�S�Fp�������Jj�e��4Yn��m`�[���հ�5i��[��C����8-f����G���x?&�2$ ܨ�0�Z<MTk� ������Sʦǈ�D#h��>s�ah���s��5��y�=Yla�ľyD��
t��s���be�{����c�]7�C�pk�:�͘�)�M���k�Vf����af��,�)��ȭ_g��{	������}ΔZ��������' ��R�h{֬�x�ߠ�����o�-��mq_� DNtQ�K��0��o�.A<�<��6ˮD���5v�#��D�b�En�*�z���D~<���揕�+ ����y�֨|�
O��,:���R�1C���HN��bpDC�͐����U��m�8�!�@�
�I��n!�$d7�$���u*7��*�-?t�����e�9�t��@��#�wB��kѽ�$G<�oM�t+4ߏC��^ڔ��OD���1��+�:���o̐�>Z�w�w��� A�`ɪ���<Ѭ����|�N}�<*Ŀ�d��.��X��/�-M�`$�"r�	��؊ԁ7�VD5�ˀ�T�n��;;�c~�eE��u_7��d��	[F�w�Ab բ1.�-�hҥ�ot�8�O]��䝈��$+߱$�ʩ1Н�1��!��K#����)FK�WeCu�Fo��N�_|>��������y�o��I�i����P�N�rL/{,�Bb赠(���o���4Si6��8\qΪ�j���=���P�a�TyP�-ݝ0�����R��d�&�Fn�W�0
�I�j&l^u�v�`�Gٱ�W���@�����C�C�w���q�qf+��0��3(^B)�X�  ���o��N���E����"�$dv�@6� "�[
�dN��4�4��.x���%���J�7����8�� m�/�f�����n����`ajy���Y�
���5�b7��q�ꢍ�Pe���M]��l	��Z�:�Z��|�́z�z�B�'��3�/ΥH���|5"��X���mg��Uf\�o�z)�I�в��+'�P�FL!y������`Y�)�,9��3/r`eȭ�m�k�A�|���J�Ɩ��u�.{�R	����o�����u�=� �����#G���1����l�]~�5i�ijn�ۊ\\.����+�����)I�_����JJ�-7�f��R�]�?�uT���" �N��}� ��~��!�n<q�BTv X�������n�j˞̕��nD�/��F�b�����m�5��!Rn)kU�ߪ��m]o�7W��,�V�C(��U�p���K��u�"��c�Y�I�d����4w�{$ȑ��#
�2Wa��Џ���(�6��}���%����5jx�Od�+�����
�� �;{���_��h�D�"�W���d�_�8:�aS�.9��"����ZY� |j�9,��?��f���kq�L�#�vyt�P'G�^΋�K�X@�ܛ����A�>Q?1��L�_��^'��;�S�f����;�{c^m��^䈦D�ۥ������W-��z�_{F�f����mI���%�S��|1�ؐr�_��,~�9��7�� �}V�d+7���h�E�8�������;�z��}�QY�n��Z��V�E��OL7xy��;�1��LU����g��ƱOJ=�\�Q����g�b<C�t$@wu�T�5+LN@G7��rM�(�>�gd���}�ȱ��>��Q�i�jl��*�v��5�)#�H��� Ab<c����JRW��F�P����G��]��$U���m����JlHU�������h��5}Cl�Bz0&R�b�ۥ��3]�P��V;�.�{�m������$�%���g=n� a<��d]C� �w��d����