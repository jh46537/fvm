��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��x� �u J䇰`#����������T�jCQ����f�}�<rcb���]�E*C�:�8T�=���2%�O�r��?Q����������c�X.�������
/�Y���O�23N.�Lu��/��8b��}�q�o�m��t%�q�o��Eϩ�6���A�_֓DۢQ������c���W�m�[l�w����ҩ���WL�� ��=ohSM�[ݏ|�P<w=ee��g���>>4!r\3M(�ǆ�Q f�0�����ݾL0��S�(E��k��ƪj��RC�>���I�B������K�����03dlu�l"��"�u,oR���l�ի$�S��A�������^��~�����"m0�u����	���c�ώ-�z�1)����e��~�T>]��C�Xa��.�ܓ~d����(�y%�6Ոf�����0 ����N�)C?�K�ە�����yd8	H�jT��?��c��V7�����@��Qu���8��*�}��;N;��?mW����g�T���i�ޫ��u�Jt��d�ީ���l�Y���I�J�x:��rM(�܊�^�dɘ�-�d!F��~;D؋#紆����0m�椣��5�ɕ�tՙa� �E�u?���*.��f���Pg����q��q�:��9��(������ (vd��X�H�R�|_U-���Am������'�<��OH�{0�@�H��F���ԡ�2�gޢ9��.����9�-�ܫ	\!	��������Y~P��1����K)��\+�HJ��,������{���ე��`�&�y��
�v>�3v�T�I����Ķ��~K�P�zQ4��/F�`Ϊ}7�����`w��]�]D���_����wW*"�N_�~mXlSZ>�4�ڒng.�nj�Awj�HP�(��m����A��X���.vO݀˙u�P_��6�m	��ە^n�0�4��s�>���w_�l^��Bҿ	D� %�'<��)v��p_!g3���Q:=�sI|:��ęK���x�YQ༜��>��+AĔ� R1��ǘ˜�����f����]°j�LC*�'FP�U�1ݣ(���C��4x�U�u�i�DV�[V�[?_*�Zku?M!<o(!u#G��D��z6Ɓ�&-H�^��9%vy8�zA�$Po:r-�g�q,�":� �.i�[�t�ٔ���f�P��3�i4襳���LƲd��{5e��B68q������A�j����S�<H~�F�*j�Te������ss�,��ǅර����I�J��eKɪ�L�yQ�R����]���7�DH����u�;�������[>�$*���u�(�OA 3���~���v�����;:~���9�:�Q_���C:i�@��ݤ�X-� hR�m�����Y��%�]��H��ԛ,=o��_��}d�����c6�D2"6��|?nJ��ՠ��w��?��f�f�AN��E��(�q�+����7sf�V�BA�+��:�Vȿ)�
�!q)&k���9�<"'��Hٮ�-��e�� ��gъ��*�n >^�~��W�o�w#�����<�����Sw��`�9����ӜR��^k��>��$ ���V?� �[UM��q�rtz�������0��@���Oi��:�#|ϩ���4���XދƦ|}\���h�k�׳8#���e�����e�x]�.��ٽ�ҿAo;i̼�uZ����$FR2�PV�+ݗ��JP_��c��7n�k-U%�Q��גb�R}��V�+@ص���Ԙq�6����D�����+fn��E|e+�n	O��	'����R�j���å�;\V�N���T�A�i�sLW�(&-3���Ϩ��mh!��>5�OZ���UL *χL愶{�4�Bi�!��9��<�m���%<�F�>ɊH�PGZ���t�V�������_�@{�-(����"�}�S�9�
��ę@,�@�2��ɽ*f���˭Qǟ������,^[��rݎ�5:;lx%�e��qt��]�Z,umc �������s�MRW�J}��{C(*� ��K����ϔ�d�ȏp'0#��h`�Ȉs+�V!����^��b�Q8��57�f��=�`��iҡi#i�x��Dq�1td�s	�� �]��Y�g?�@� �:�����v�;��Ūν�_��� Q!�u�'�Yӝ���Q��� w�}H9�i�+��pN�Xy���#�v���-�G)Ag�硍�X��#�HC%�0}�$��x��X���ȫ'�d�H�l��n�\��iڭǍi�4n������k�-2���sx�'<
�@o���;D����?�%tᎹ��X�6(^Qj�w;�x������i�H�Ӗ�p_6J�ǋ@x9�sE�=N��Y�}Q����{z"���N�f%|V�Vɒy�JրK(�
��d�2�K�Ăؾb�I2���r�!�uJ(�������������p��+'�ť;������@�����C��:#>쭨��&��jI����Q�i��hC�9]�{�H/k�X�Q��,�R��|4b=Az
���:x�t�leLAFZa�N��%;���3hڳ�SR�6�u��t%����G��E�5����>^�o�a�����+��WS���7���rZ�){#�������iG
3/�z�q�]?z�ٙ��2���}�ۄ	�2��	M8��u�RXp|u�ԥ�ǃ
���
-ҏ
I#u�d��̷�kb�qdy�`+,��	7���`2�ծc=0�9��V���Ԣ�An#���M���,�ӿX���d}\�0n#�	:��sFUK�Zٟ+�jXt#���O������D������l��}�����V�i�4�)#��ݝ��ǙNw�҆w���F�&�x�@��r��7�]"/�0kK1lF�X�Z��Z«㊟�N����e̅jN��)Fa)Y���D0�VQ��hڈL�&x0�7B��)Zb�UPqxO���oDL���\��,���p��H��ō���+X�B�{���wV���Om>"�f�'�?D�Ά�#V�wH�q
���y��
=p~ε-�J�����"��d�����q�P~�dW*��u���"Sg�^O/��� �)G`*�#���Nt����7�I���'^��ͭ��)Za�-;=����d��\�h�ۿ�M���&�ac�ɝ���]�TI`�%B@FҐ,�+&�꘲��"�G@��_x�fܛ9q�"Y9���?�6�WF)*�E9T䗆P,��)(��m*���U�	���;L���r�`�l�Y;��e�ѽ�2O��F���f��u���u1 �g��(k�G}z��D��T�I+�k&$&C�N@�W��SC�VDS��n^ꊦ�L@��������G��D҈���;����"����1F����;/�8�1��t�i���[�4�~��F�/-��Mg$��^��v���_P��U-�RpX]X�{ FB�wP�eWQ3�֟ݝc�'a6LA[�h��A��CWP4	���sLA<��pn7x���UIӐ�����r�?�B���`��^��2��,���q���D��4��-Jq3\�@��/�V����� >D%Y�;�!�5�Ei_���0AB��4�6&�����Bc�b)�>����3������Zzm�D����Gh�G��J<��}�|N�u6�N���� �E�j5�������� /F���ґ���B�xC�ȉ�x����P^H������#A��h�o�!h �gD��i��Nn�}����5��)���pR͞Ne��2 ��jg�^��3��jw�gN4 瑽��#fԆ�����+��;
G������%e�s���Pr�#D���=2ZϜt�	�0%"���"�{� A�+�D���̈́����@�)"����mc��6��-q��E	�(Յ�SS��߷�ԃ���_"�Jtm�E�Vz�ۿ�k��X"ӌ/��-D�`����WF�DadU1�@ y^)�!ʵN"&���$7����s�X�q�i����J3y�M�т�[Ħ��&~�	,��wj�ZK��hC�͈KE84D��}��*��s%�?���
B��N��lv{����*NH��q����X���=�n�Q�;%d���.��<�(�C	�v|�?��Q;�E�)Y�s����$��� ��q���ϔc`��!�������S���:�=s�8l�B��� WoAO����s���Ʈpk�@�и�C�n��j{�'}ȫ��V���mn�ڌ4w�TIF���8�!�O��m���WPm��p�[*_�E��,���DXAR�+ S�THg����<�|���L����K��z�fAR�bD%Hr�L'����]�]����i�T->?���~�Oq����>�i��m�}�'4ˀx�� �z���¬��%	U��{?iLQ�~���I�E��w�i���GhT�{tH��"h3��`ҩ�3���k�j���^W#���1��2俾\D��^*<	��ݝ�v�O8n���c�