��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���� 6�:$���mQ�$��z��˙Y��ˍΣq�N�5sd%[s�����a�=�F,�9�z䮴+��e9�xh������"��s���\2%t���o����	���y!��}l�[}�{Ҁ�^~Yo�}k�&C/af�+�Έ!Y�����.�@��µc�P���Pn {���}�+�NupYH���_:P��A1+���n� ���K��,��Ǉ��\�д�E�(��71a�N�c8�k.�ᨃF�LoK�T=	�p��v}���o�;oM���|����l��o��^��k�)��m�4�ǿ�#.�;�+ILϚM}1����E��^*�xe�>|�x&��f�V"��,ߓ��@��c�4�p�&��*��Z^R|�oa�#_K��P:��~5� �/E�n0m�跼`�-�"�W�
���TĿ���׸-��~��JV@:#m<�.	Px/FQ�?��������%|���ݴp���<����~S���X��ǂ�j�Ө��gW�x(�:`ɛ��3���3]�܊��$*�S�t/�~�~Da��������*/�+�,�G�!�z�Ž��8�U��$���|q��s	Z.�Z��~�	�&Ѩ=���@�RM���������eĤ'�^���5�lT�����s j�	��z�9;�OFDW�8.���9`"s�_q24<=��ѽd%ߤeA��E�:v�
��HF����譼S�������4��K�;|���flV��C�A1�S9w{'��KQdۥ�R�x���Уt���u��˯[�##�z�FGU0�y�ɀ&��Å M�9c.���nl�&�	�qU�!q6�X���$�CѡRJ(0 8T���p�}���*�B䈶#k�*���@ �T�v�Zs'Q�ϒf��	�*�*8��ҍޤ\��(x��`>�<:�\���l�x�}���B���x����L-3�n�%ң�}����6��B�$�bն,��|eZ�XP4گ=@�!.e�[Ǐ�'�&���X��״�ˊ�q�[�Tmg�sx �����-ȑ7=�s��O!qq�^;k7���2��@J5����S��yZ���{�������Nϱ�q)�t��ۍf���|sJ����f��yTu"��웘H �ȹ05��T���!�?+k�,0�� #�;B0Z�iw_T���z.��}��A�j�P���8���Ȃ-��s�_Ɨu��O���ߜG\�L3�9��j��Hi�oRJA/4_3z��,��v�(S7�Y�Bzk��=��͏k�1Z��e�`VZ�$)5%�9}}�<�v�� ��0�!��X�&��	����)"_�c+�/�ޥ�qD��9�RL�;@:\��᪴]���;I��� ���Ky��i�x�.+0a�����M��#�GE�z��Bjp�a;wl�ǥcE�ĩ�l�I���B쫡�����3���Ⱉ&'��ix�~�֟��	FCVO^�@P���Y�o���T�yU�V48]q�\T��3©���t��\��=�/�r��C~c��@W>�5��e�X����0�9 3�h<[�V��F����2�	��,��"F�)��g�@�Eb��'������O��hٗe�D+���P0�ܣ�%�.����]�l�0�ڝ�dvp�4ߓ��u�*̝I@�..�E�Y�gC"�*ۊ�#}% �[@�P��3����N��&���Fo�WxSa�(��G�Z�[�c?�m�C!��R1�,����wMhϑ�*���I(
��UZ���ܢ�U�,zs����6«�M���Kq�p���<���
��)��`ᩊ˨�]�m��MN�7k���6O��ל��G�����Ai���/�M��?�A�����VY��,���]��ϭ*�d7�~!�"J4�c�t&����T_�Pc���8��S��
� �:��q%�gq�-��9�b�6mH#h�|��"I4��h*b
�qwڝ�'���綱�?��=`����zהg��ͅC���r�y���j�b��#�|n��#"l��TF���[|%�& ��D��� a���B������ɕ��n�d	Jy�Q�����yg�f�v+bꙡ��W]��]"y�Sy�v]�W�镴��ji�J��?��P (��YMn�ZQ�)8I�XJ[�������W K09A8�R� �[J����(w����=ŭ�ͽ�Q�����$��dm-y���s�v����0yZ��lW2�˭4J���#��(�;�8C��5��I�2EO�;~PI����FKE��wԣ)Z�O�}fi(��ۺ���]d�'�������lr�����c�r��qbt
�Ϸ�0�8PWg0�c��W���4�m"��;��h���%F}_� 3Q�P���|�b���>n6�Ӝ��)a=�\�5f�e��D��\00�� P�T���\�֨��f�6�A���y��$�(�p����p(q�^�;O��.	j<ѣɏ�̝5�U*C��$��
u�s-Xdya���w���'���e�&�������S�Ƈ�̎�Y'��z�d�^��	%�ܗ�Au}uNA���
�fc���c�Xn�!����-�^�y�P�L���Z���O��fa�~�O�8Ki�l���X!�e&�a�hԝ�[K�굸p��.[����.%qTؔV���a���|��\�kG�:��e�be��2��l1�A����q#�0 iE�S�!\2�N� ^敉�j�m.���j��3Q��+�g�1$
��C��n�xĂ&�p�i5����QR�vA��ҟ�ƥ��k��Ҩ��^����"K�f