��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{�J	�'=����5I=�%	ڛ��v�o�o$��D:$�=1�=��L9��)+�>x�P�ߘ?Nc�v�'��;Xq������c����ڢ�������r-�s���R��V�����o�dS��^g��\Q�)��D<�|��� �9h�����J8��T8k����?ڌl�6T��a� 
G���q��%T5!l�T� mξ{2X˺��i���0��Z.�O߭:�B��P�v�'�.ؘ�f���Cve=]נF4�c˄�s"� Cd�Ѫ�[*���^����ގ�9�A�Ѿ��D�?F�8�>�{�k)�'��R�åwobfD%O�H%5��.mɾ������b;�u�%jZ�yyg}��-�_�\�M�+c~H����q��R��Y1����׻�<M	�,Q?8:W@���k��|8A5��>�����WjJ�YC�)�B�l�`��H�2�Б��	�FSFOEs2�K���}<Z�@�Q}��xٻ��ĥ��ܟ�|%�IQ���{O���y�|��Ӽ�^n�o���R���da�y3;�~gEB?��Th-���b�G�ܷ�����k@��j7�([Z�o����n6}�+�Y�z�ʊ�[>¿�XX)2���[��x�0��ndc8��s��sv%��ЧM%R��)��.Q.Et��y�[� ��\��z�A�T����HL�؈�#i���[Đl�P#�9 �,�y�����05�XEȽ�j��g#r��1
��-	�u�4�[��]�MI���]��ON�<�����	�u˃D<!��W��^>��q%�cl�I�[���$�ლ�~Z?�I�K�� ���ޭ�
�~��fx]Z�K���uX�/2o�5-��H��u@�����N��\ݟ.[�O~�>�%�X�tn�^���wN>>��l5��,�QJ* \�e�ވ��2�:��1�ᶢ�)z#�0/��]�
HmJ�{�N`���>�#��.��������?��z�� �����q�/I6ME��n
CS��1tѕ&Cb ��Z�ٖ%��؍>mF���B�)eM0�K�,i\�v>g�謁.�����1�S�^v		]��K��XQ�l������]c�[F�y����+:��M�=�V?�19��g��-�*��&
���:Ŏ~�����S���b�F|�
�>_DI���!@�$a
-V���Hs�`����~����-�����(t�8&~�t�$\Ɍ��$�#��x�l2:A5���7>X���L�u�%spΩ=�(��@p�D|3F[�t>[��5�uE��He��LY�5�`�SWG�Ԯ)f(n��It�c����̊	a���ߪV��q�_Q���k�x��g��o��g�@U�Y(��2���������Z�?iL�%M�B�G�?hM ��R�vչ�j�6����%��������^���U5�!8��H�S(��7v:�ٰ��R��V���]fЀ�!l1�����K��0�~YQ���G!�{��o�J�*qj3D�(�Tnۍ�v��lf¼�W5�HWP<��r͌+�l�=b�K7ka_!ӿ�L@d��ꙧ~�a���4��� �^�T��28�&64nʖ����C��}�9�7dM�]4M�,��������
=r�1�&���k�5 y9����o��̿C�:܉Km4��di�d��SO�9���0�i��wѝ��kz��l�CRd<$yQ[��!E���R�q��Lۋ��-�5�����S
�=�cd���[UH cGz���W�ҁ O.Jb./ՠ��:<?qJ:���a�(�*�0�#�"���!���a��8���"3.c �Z��iY���_�݋Gw(����m�Ea\:�v�7����'��N�s�yv�f�߄`QI�����*vP�t	A�˴�b2"���.���ԩY�}�#<ka.��0R� M�R�����Z�I��6q�vP\m;��b}�7���E��H3�[�z�ח���r�S���E�X � G	��g�2�� >�Jb��%�T�19���ڼ
�]�{��@�&�'����a���--=����������ށF����� �{�9	�@��������T;��L�pp���b͢\T���c���U��ɯ[e?�(y�W��_,w	(7�]��c�