// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tNGBSy41csZjylSouFmaQ2uVTlg/Xm2bpmI87eQrLUsbz/9ToCpJXCJQmdS094Dk
k0SDYyLUhe1QmqPrbY4nfdXsbF2CmpYxFcl9nzZ4Nz5QtmDvseY8rdHAOVM+v6H5
ACmHU7kofS12yhoJJdPiP2q2FWl70diqargSiu+tiMA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11920)
8vwLByBk2wdIfSaX99ZcObF9zo1Oxp/AOdAyVodKvWE4VdCvjaY2uWjnOxOmuDqp
5aRl7OR7VN+C13ZVc/buO4rW3QHN7fK2d2I/BL1xkdIsNT8zD/fkrgHT/G3/LePm
wGMv5Sn94fy8CvhQPp5IVyWoB6NnLUgWlrRdYZRhFNfRAG6SWCGUZtMM4/ngL+TD
MSt5iTst29yW1oBmHXjxNL0/lFOAGRoHJf5eBJRLPandtNV3rypenmX8V7jEqTX0
MCvvo96Z8nM/vH/FYnvQqKeglz9VtfxSI7Frm7/g9ItWrJqbUo0CHztbfbNQGaoQ
tst2HDbBAXT7ZAlsufb9ZhmhE+KcvhVLb1CWgfbu8BLoxFnKVOJqk3HfnF7d7BWh
Ar5mB5ziLQKT9OGWOOywZd8i3SKgnU78cRApHOL/CXIAEY8Te4oaUicYjyyaXN0c
UhzAXwEHxpsDCUcA/+I7nUXfCi8KccojmbKZ5tbRLYr0nE236cCbzgPaBFOt8b0j
ocJTQt7RNf+EQjdkfUt+gB6RIX/qZK5h+eOZQpHHtPujVGjCsB7vcRAOy1raotup
p2v29PmEnzrDDOx+iqiFaiTtonedeYPExKLFnwnFnCJxOJqGI6hjEkYYa3fyvVSL
irER57uw0pBZp+ePakSnZ4a3yQnXHSW/yYBa/5I2pRe0AcYEi9NPgD3xqhzzmqM5
Iv1j6TXxOzYUQVcjpeb0CI/rhxxWGhBmuH2Jv95cxChGXpeZIoNBImx0juicE6nn
YqYLPoFFwtUDDZhrH6jCCtEk8toMZUI3mf9cHbVzXDDFI4BQV5Ql6qEycidHQw/l
QebruI/GcB2GTL1O139G2EaRx60HtL1oaqP32yxqOPGbhC3V93ZYVg1H87m0kkfl
MVmyr8pGY8ZxUTqHUf1r5sxXCar4J3jKEupouH+XWiTh7hkktYQNew/kX/1cwmPz
vPdoDNzc/YoJ89etE2IhRg6L+9GcMqBMfFxbwaX89WvQbeAE1gyyztsDEbrBl5FS
dXwgp0S9pyDogwGtnSDUZmv8SKLhY7QegfcwxoXGbEOVgZYPkzyJIhoOy3KmFy72
GakeiSIiRkOEVPWRCM1t1EXMnfSc78nJ2VlQBuVOHqQRJxzPJwNKATuF+XzBEXdz
bAuFb+4KJp2jmuoRJT//EOPMzEFN4rhKMlgZxSkaStGfgvND1+1kD/ctA9IkYTVj
qu1xgyPPlbsn8px708NHLo4Gkb4x2V3RYMqPkn6y09pTs0W4iEwPaL6tfKxgxWWB
wQq4HRoRAJ7MX2c2It24chlENI97F7UhK29qqHzUX/gS8K4kjtGwaMomaeIRwjvD
OviBukWCvz19YNTYPwHdVHhRN0K3QjEbkZ5ZFRnSiwUJFvkazHeRiamSrOnO7lWl
iaSr6iDpVQIsWM8hD+NuptTNBtyzV4GvT/rEvR1ntvQw3cZK1LxtEuv50y/UWYUQ
BaLcDTgmLb8WmpRJf1q3YHeV6CrIXcVvE9v5dLB2nF/drbygnl01NL97N4kXoAkB
5CxbHXvjRCrB8ysDEBsSoagOHKTeNkSzfV+EVtbUNaUvASXo6mNRZLupdUh1O+Zc
NQEHVpsewVRG8zNhgSDriRpB+zMhP3OFWqm+pzAxIKcdrGzfqqr8k7ManlaGMfAc
4wLN9HhSY+oio735DE3lifvbnIBMPT4WHk+Uj1R0s5YVnMguHnfqHAzgJmkhck5C
UueiqZIKJ5/8u/sLD/iyeaJdezgQSUnzXdgk1OZ5txq4KZQinmBIoUjoQMO9xV0p
cmIPo0dDI4w9/ywyMBjdaqZqyYxMAbKEEpA/iAhLColGAnn5iW/0YJ8Fnis2MFXu
1To71hNRXOhXgEsVRmeI2Be8+ZJw6t9IUl7ekrDt1obVXJLUcnS95g2cqqvfZ0te
Ix2vlphCTaCb9jaiCuJhgtPBM7opIOV4BDxWXv7Y11NoXstCOftRXm4QpcznmR+A
30n1KLz9Hn0p9J6igr2KKNbE5FZvmBxHq3rmrfizIvtg+F/BsySUnCRoQ9F0gK+t
6a+Py7uVpwcg9oRm8z62D0UkNQnFhfqzUgjyikvD/x6LfzqkfKMFMjFvkyKVPYQc
lwZj5lPXxuGqPYUFo6Uhtu7C5zjov08i8rHD3Fl4df0NkiLtzgvYk3TfZRa5F9Ak
qUeafxrgGc7ZxeGGV18IhLmTCbCrvqNjelGmdc5D78baR6ptQrQF0fpEihgyWbGg
/E3H7V6VAheDomBjrg05HvdRy43twKvvbz+8tdcUhc+yKPK93xDD5uATABSKjhLC
cLt4/HFAenbTxDaGb28CSzx2WGfQkV/UO/c69bjNUJjaFDPkXflCn4tOwHteNBTO
QlBZ9CObWWywATwXSjzLQGn1Ts8Vr8Y1MsuyoOKKK0cmUGj03ivjc7NwRqlrpcRZ
Qpx3PSTjjaZTfYF2vqYY3iXyl+qs0OrSdhsKhL9+xoIAzsbQRLjQPp0UXIBUmW2m
+SaTu4HkPj59XLZFeu8/yTv3ol5Q/0LCg9MXkjnDvUvzG8bh3rhFtCWTzxQmo5sE
sY+410nzubVSkWQh7m1YZIiVdssVdgBYiSmX3MOfGwfIDMgVRQvcOlYgGAbvjwnS
3LNgIkApDh2y7MPKwyQSb1cQhJR3CinQCxACZEZ957WE0YVD5er5Nc7LLS/K/9G+
jN5mgkhDo9iAGR3kGft7Ac1C7sEcr/yLRLP4kHD0/Dw3EvfqZd8XQYUAWUx85Jyl
xY1Z0eTpzvZ/NaIgSmtoEw8I1bK0eL4GdvDJJ2KtTldXDE/eQXVTvxYMrfoo/7o1
gtFUXzmvJstRYDIXVBOB0BzjYFZoofnwa7lWr/Z4+50LKMd75tVxmpDX6HwMsmX5
E8a/MmXSAp0yo1qhgFH4UY4YcM9rtOd9wR/Jeeeh2tgnIRCUh5QsE1nfyTG5tBkj
3dgVpzeiGdwp1mGRowftu7EnHU5GezfauhfJKfBWcQlhdQKq0AIt6ME82WFkif92
CTazJuE3EuOqMrNGXXtkE1xUeEybr7zfZwmXUzOq1PvnDsVsVvXLz91pk5iobh5J
GhM9PcW7hJfhMn7V9fbNHNAn4SuaSMej4qZ0ghZc+hXxMD7JxS5tJBXy+byzY0+k
apuE9HBK+Vwh4oRpoYoemEFaHc/z4h58BjTB1H2QYCq0jdsiNLl5pBcRsMLFdjmh
OFEMYl3YAwenOKQQZ/WBoyoX7z2YD+2LvRRdvsQu/n/G/WOUdAtWjsithb8GYBrd
welfn33Q5PD7JjVZznkjM36RVVQNZUvo5vzBMNk8s7Q60nCSkQ5ftYR9T0aAxyiK
diF3SRWIh3c9jsTNfDulmf7l0bOPzxx5jwPa0etKN9i/9IsoSPfbBRcTQiTOFBWH
C88hx1QvqU+5GXtwzOFIBc4kwBtzhF3Gj5+mEtCBwslSckAxFSrEuzSzJkDs+s02
W8flDszVzU3kZosIIqdkIMgh7+z1+3dvXZQYalnopz+xBErM5cDqyM65viPaKfmC
x8Gvp25jk4AkvyJoDIxHmmgDfL+rXO9jkVL+yTug7xHsz5jl5TSr6YTJcVv9/vq8
+EWUQgrqfF3Db5uIWUKwi0/90f746GG1Z02DK1DEuMpEF828Ew6MOcEi0uvO6CMq
lcoFf9VwjPXl5nee/x2A6hVuYHYIZ/VK+X9eg8yIxhlwJcB29d5Z6C8D7+5JJNy4
axNE2Wfy6ulJnhGA5+0FZD4s9vE5/ws/e+KNBUnFzqUbkDhv3Ef0U7TMZibJpnR3
D8+6vA9SB8dwmX/5Q7/ulRasXe57Gm+smmY7pjY920mVHF28+Fs0Zdf04SXpwCLX
WBLdF3pt2mNwHjlwFBVvHRgq3L4r46qFmRiXWC7gBSZMLgOOv+Hj1yiBlikClsQp
ht6N0mdOVgf4fAkIGEdnpg8s+i0jw4s+6LEUs1/Hy6KslE8SSycaQfZUQ48io/DQ
HqlgGuWKmXQxm7aLBBY3pgsFRZw8sFXv22DpMMoUcW66drkZBxmLAwsinsRz1XBi
QCH94+U8lkLsjqHFY2/h258mSsUYy0LBXnpDmIg6TDnMyVYX5w0tPp1OhGRBVUIk
lHqn9LMsoZfI1xFEgOwJhReiHaKVl7jaUqXoTOq4fF2WL4XbdMO5UQ8DPTxBDcTU
girGQzsaUxg6or85/bedIu1kLQz9lXABuZs40xZBOZMT/Byqo3OCf30rjPdxb2l5
yaUFoTpp5NZ4CynriTB9x9OHcqAxQqoee0Ob533JhQEImsUlF9ORQVAeyy6sd1UG
LzJEiNW3nuQJzXU8+/5oWHsUy09mVYFEt4V0xX7vEpJYWSWC6LumPEwWGFNOmK47
16UKIktzshjz1Np7FsA9MHZIDsxaUTvUSXw8ySIn/M5HT+vx0pQWu04CvRkCV9Nv
0VL/oxwHFwV+3tKDEQeKcW5Roo6tY6DR/HfAZVOoPTcFqMIKNN6YGbDC5k0Bna7b
vp6GPNiWglV13xW/f5oT/DnVk8BfYLil6Li67FRldmOw0HgFIaCfL7dOZ2YF3cPL
/vHjsss41BKa1hvTvx0z8C1x57pvlCir6TsY09eyfVwi2GK9ZHLvhiM/XWC2NmMR
HPdPfgU/SjRI7PKzc5lKgs/3UZn/RmwmLmB8vUYB3P6pDu3dRTVYvCpy2BOdVTY1
XPz3qpqSn6X3qKx0tHQfzLeYWGPHc3qEDBebpFjFQXSGxn5PHh3/H6ue2lY9MmL6
VI1gUI3AohcK2AkddSkp5jQpG8uyDo//EcCsRshtLdK4EeNef5j7pM38bfS5oq/H
wOIGLXyXtxoUpHlxwXVHLs83//NWT444pi6gGWAsw9i5AvJD+QOPpDG1ZNBTE99u
3P+0P0KsGX7jThBPE8C3Op8gT4xWLm9VwQY83VH197xabd38T8gYiZo2hR5UsVVL
F8L9arcqLB9Fl8oYtDKMaKKpDMp3k4t0JzSOk6uScmeYhsCSNjWD93YNCGywgXmQ
HPKG+/3D/ptAcZFaiIAfMDPNo3yF2dJrZjdboE8Zdikttb3sFOrzKwjCLxGUV987
ax9GzL+mO7nqXMHuFkRg2pYtB4C3L28aEQrgy+giReL3f5fk0tLC2zqyBYRJIUCO
UOlRv8kjlsLh0HoYL9ODPTSSDRyhHffihflsH/1F1RUWnFB9HYTdZJ969r2/ccD4
eHZiCI4XX4SI0x0eq2eBdD/qB3S7hYF03BmdDaZId9lVzqjvtqF4Z3fg+aHDMZyG
VhVb+HOzCdD0Hh0AEiAv1J8/PgYgILN5T3166QTF2JuoWW2hrI0Dyk+r5aE76mmb
3PumfeTG0vGv3kQkPgbDaT3z+hvjMymuJD+TXSwLWHs6sToJKWACLwbMdyvlEr4z
pNYBylDg+C2fcYco9pl7JN9rqVz7zWC40P1JqfBlRva4RI2n7N1YMEo18xehZr5T
mBWHcMNYH++EuLQTkR9K/9YepnQJYSglGfRXCYAUT+qKly8VXsnF1TE6kZbDiJz9
zT8jwwdBqd/SVkbGOkvASXwy6HAz/BlyjpElqPNn0IwQp3uOqB20048o6zBLewBl
3VcV3z2UVPuuHM0s6JxR9qxahZ1FLifl/9rG2ZXT8wsPDcFPLmPk54nq3ERGwVBZ
aQuvseU9aa2grS5s/2QoInjUhi02aKl7SgmQKeg1XyBzTGT+Cm+dZwZKmPOGs+qx
VfKNcAgbPgU361NJ/6DryeWESerCljz5LVqb03LvtsAXj+P0q9AldDBoSTX9RkNv
Giow+ewY+6iRvBnB9jYggRisT3cD5QohDwouozEDImrKUSRHfCjtll2GbXge8r+B
dwtwKpwphy8O+pRv/rz0YzBVPMYrVaANvkSrU9zHBTOoKmumUfLZryHbFfflrz0t
gERGDT3yyImEfbtcIZPSLXGCCTWVlzrTeKYJtbC/q5kbB+oHyeN2ITYWRigBD71W
5zOqBOMOz6H8eEIoguFFDfEkVMDNEhBNcq8cVZWoRCEUWOw7i9g9Cph75dazo/Uw
5OtJrJXSaaBEqP47N0tdrGvQCdTybW/ZGsAbJomPzJyNlU+0RRK0cvuZh7fl+Qa0
KBQJBi8lj6eZ+nmt4kSAz4qg7IPHLl1+fLioij5mqpQYpsfJkXW+D6OSGzrRC9Kl
W2ovV7vrrvMvwo9mmNfB4CJlSsW5GUbkiug4TR20ByCmAtPagfgl7mNNuv5yU4oO
TftIJPQyrhxN7m5Cy4idJQf+EDoiZciqerKvgWnIT7WSULukvZQ3Z50Wwx/lIAJf
mW65D8if2eFMsqy4qV5s9rI9sdAo9QXI+EyU0eleFRRgmGqWdG4CBfa/17xTG7Px
kDoubpu1oJDzDddXPxV26d0TMkzC1CGcgR5S+v7i5okKysQKaFxM+Hx+6of882wI
Mk6la25Q0zqxx+BnGYGwmY6fhriuC6ADM2Px9gKdOaWxjPhpCUDMFuIS4dVHaZUf
vn5vsdWiMpUnpxdrxHuHWIKxoWCOq0BUj7OeEmzN+uD+UIFxNVlhVTMHZHtQlGLD
IMUZ4CMgG74Y50bfKLBkYo8Fsub8WTbdWP6ZRNfjkl+3iY7q0+ddMNYzr3slUuFy
+jqQ69rEY4RtFBidebdtcMmJJfqZk8Z5ah6X7PIB1Eqh3nyPGBngpOpMWj5XFBKV
3LqRHMJEcfbq8OGUW7DVdYeFvlPW/NPfbtiU7Gd9LP5ze4lqNJdmDOvDQgqewqL6
KW6I1UWZzb7Tbd7DMxWBgpKGjXcsRQ2u8oxa0JYRpWC5ehpBzRsTZdppY0X3QhMr
pN7w+tHEImBXXskmRdOX5uuKqZ5PNv4p+sPUDNzv0gBaq/u73vl6iVUp6cryQ3aH
YgK7GyXF5MmDdYjsITXvcMNVqzATTD29YFyRxs04tBnEMsQ9cdjCJt+f61uW6yxv
EGWkJO1SZAr+an1/eCeZT1oJfzMCtLoRLjW5H8X/4O4H0Tt4c9SYEpWs7OoLUh9O
6lTq7V5PLPRTlpW9ca8dlryzmDrFoeKkjEh6EYsHZ2noS92//pOHm2yYwaxomc8W
UEsXS+XiRnDKZzyp+bMZe51ljmUkfu5KRFRihMdk1MtlWfyp1hCGHq3LUs4g2Hl4
JJdUrHfD6L62nyjj1FURSUarsTMtfg2Rfofn6SKCFxka+hB2StHDuRAl2Ls6ycU8
Zk2zZdYZtfuRJcc5pKmwpVD9VMtfES315O4ChBuPJOWC0gDyPles7vej81WYg4vK
UoC8zQ8klU1Ax9+865fVFGBHanvljtcrgei4CxOn6qzR1mCGD/PXljzrz9E2S3Nq
Pm137+XqQ6zsXTtybHVK4mpLbvCr2In6ioCHkvR5odb2kWDZ+UxiC3WZQinLUZmG
SxPpnw7k0Phi6TCQwc0owaE6tNhHWQT6SH6aWquE/Y7H9Q+clxlizFMhmsea4aQJ
eaJRpUVEHdzGVOX6MinzPWkRjDB7Rt8Gx/BqevTMaHoDjuU1BHHoEYqlVdoF+Azn
z70j2+B0F5VsUpcQHpkDMIuUjcQJMAbdG0wEKnoxqWd8zAoFu+ttfjW80Omd4dkn
LeVu8xmjSuBwrFPL0SJnwqsyg1PBRtWimGOLTqJo0NGCpPVSuNobCB4yi/60+ANE
YHaZF/Bd+rSQ83d8WXXWXVcth/FY7WbjKFUUZB6vf5qhm1bxsbKw0Jjj93bAlwX2
1lSsHWKo5q8RrTCSrYU+Dw5j8a6ORqrwTmSXGtdV6acitbV/aExAIfouXBcmCVlA
1BTGMujaab30UXPcvsxPTfx6Z1S2bugvAITIE292OBOajKpYffmmSIymKxx6mVDI
d8qQph2162Uaqk7IBmPborBvVrAFTA2Kal2BjtA9TG1rDWtf0ECKxdvohys+Ss2A
er4njyOS55C/bkOrrEB6E+oDH4H2ItBV6z16qaCARzyfNoribQOdALJ7XO1gPnPN
BXQQXk+sQ8eXdOJZoG/DNVE27KsVEpUeNi5rQZphpYuSXXBLllVdtgm9Y2D0lMrx
WT0zWU/Xts3uV1tKV6wqe0ZB2KyjSqx8qA9E9ls5F7ya8X0XzvUmD3MPohwdaNoq
pooMsRQ9AKN25r8BfgjJx+U6jmr010XQojnqZWts2W+4+Q3+OXeMSp/fqCkiVdPp
mgTI1daj9wvUFT+xXGSbm9/b0i/6kZGrVO/JUclpI7TwDQ35DSZeNsASM9lJwUnC
GudxbNSP2bJo5aRdFkOQVPqGSjzifQZ3mHaTBcgjisAUoBS6JQ9o2aEXhmEhtlYS
asDa8w9BC02r/SJuLHf7anCBvVT6Vx5DCknxiUs/nktGTkHW2fvR9oKK0ygzxaZG
ziMdH8DiyHLQP3G5CRZq/buSW+rf0GYJLR8VCVNSs6LRtJMiJ48hjcxKL9Oq/4cU
4btUc57bFQjGx9MLLFe9lDLFgyfhvHrXlVJhPZvdi8Fba1QYqToT6abjsVtWiNug
vL/2jftotMFHyvJud4hVANJV7mi78srI347rrHsogU5OtnUq2mlpziNMa95/EtyR
wUkCYW2pu9g2JHfsD/rN/pKSVCCsY8fU4sORFgV/UB5rEvs98UPHqW5c7Py6YinG
q3cJd50ACZ+S7yE0uBfLDkv2ZdNhvlQU1HKLoRRMgPr1wFrJT7/HGzM7+kp5k5i8
Ebi6udtRPfETv43FArBCvIhngYv/kG5IUhNn7JHZqgWL7NMt2bp3fIKwuehX2Qsu
e8uzZQye+NEWQN3CJQRfeetxKzFm64r8PB8EquIeiLPjy27aOG0UX/gmrXZGb3Bn
WUZIEeS0APrNUpxLb5vDATL0jZ/+9IRUPuwGr2WT8B7O/wiJaVN3H68NFQLwKkOp
ffJfkIUuytjhEbMM3L2E5gLX+LOm8L5UgHzryuV1o4Dw8FH02mndHvRR6R+WfNFD
jtP01vdwjzDSIEZ3cqGT6yJL9lpE2xE2gqttRJ+LwwBATLEZumropd4nlJnMBH8z
nNjazTF042I8KfYR8A4fUW8BplG3C2DBXlj3uEOncH5pay98r77E+XAaiojSvZRE
4+wvCHaWX8xRcyEqnl4QwJOLQxuJ9l0UNhp6S1UZm3OgRB58+aBWzsrTw+0j4DTv
RYurMKjYJ/gavKdXHY0WN41TMzT7v7ozUC11XF+DhkHYuOe+E20P+Y30Q4FVLeBG
rSSC0NCakwUNHLqkAhcmt5LASECFBqg9QSNdQwGzk5hTJRg7kqzfRRq2F4Gh54Ys
rRYGQ1UrcTfz51QXXWSvfL4/AkjfRRJOIHmx/mORu/TtGCldtXw/LFGTi8hFtQN3
vUwgxHiyuoycv2cYr/OTqe9g8C+FvUpDWvGyltbKmI7j1Xyl/m19OI0NMlZLSwiP
JB7nP1YVxv5lepnOuntBCD8deEQwUj8FmXfnrwYQap8Tq/FCcYV9fM+prFPJTWkP
oi6pKIoBNp43fxTMQpMwJVnSRzaN0/jATZ58rJWc4oZ2BA4qWs3OGA59qOLYnILa
M/dWDaJKszfQVR8rg4vZF1X2SlpFpGRogqmXsqH+rAqKX8Cv1AHnMtEKpfcudhN1
IiaAGoHtGhnwYbRfE1UD+ll4XeBYRJ1GtqN+7Oh0Ygm2EmVdJ0fERuvz5+Z3guV+
XM9rZbeeu6fDvyOCF/E0vrGub/A76eh8Y1OTDJDBynzXSxBe8eASLr8uiTA1wCSO
vgYfm6uuP65FhGOFn3Cm1AMRaZJgDZM9K5QQGJqqWI5qTRRSoSi9QOZ3SqskimIm
HX+J4EFXb8jbkWX1N0m18AC9/6tyG7F7PQ9CQpiSOq9huJLx7Y7n1FX9nGpN76mg
uF7xWt5TMXxFxjZdGpGAzEeNrwwwcyx608Xof1dASVJqKNjgWM5EZxtceDq2wZCn
HXyKICaJ3Pwb0AsvEoI75G6NZslODlz+IBSJuoQe5nFO1eefHRr5JvGs6oUeUEdf
MX3wQFT5Hhi8WiDxNrQqPivyPdykQ+WwBhFXWH49aT9pMsHhfWzz7GVTGQq7L/s9
VbU3mrhpdqcGqjXcwHr+tFqmIad+dhxxmhNwwTkKoWqe1uyAi1KAEZWp6qQzZH6u
02PJ38Hhe4A0+qnleV6rESL8k0XWK1PFOv4aqeC+pCgKci+eqcqB2Xr3Pxf5zmAT
AFdz80C+SxewTrE8JOFF9fjWKCbzoxh3Ft9tSYpC3hHj5QCgxCMjhdBYaRbTDhb6
bbyWdqfv/whbdoBb348sRUhasl+yqsUby1brUfflqz7/nFusGIna2pYPDMimdGoB
HREi+yizl7PpeH0Ebiw0c4Tzf8jf3bDlAfrw4B4NVxN89uaYj4nLDbRBym6vIRH0
pexGKifdsg7kRimVus+IM/UcnxyHsgHH2TRld/Ma4QRXasdjw71hZAhj799+0wR7
BxmT5GBmjqdnOxRNQuHt+WutPXM9O7EaJbi4dQDaatUwZwNgY2ryq8pIK0Bg5PeP
ZhSnqMFDqCQn06X9gc4ldkvOyR8+8lKpO6PdSKRrFJ9r35YWXiMwbSo2SJSVTwAG
jXDqiFYGye3IGsgVa3yblDg5G20DWSaNoJOHxRcgidCr3bJqmY4kyX9VYrVoQith
JTlP9/i1D4a6OrkuY0rPyRQamavAggeLCLmWQlDr2/bki9DMt1vUN+qbUnvTiSVT
2mIzOrGJGbDc5/AUvyNpRWAWVocuZqp3br3yVByS0E+eriASMiwukUa6KqXLCB8P
aDvy0+XlkX/oZy8PzjzhEhyf7+oxANYOOSYDiLTbDVg7h75sSGpljg11pth2dJL0
bapyo4jSZN+M8Y0K+BIGkJT5le1LXyV8oIuRwFmYblmxFpMT1a+ILzYy8qWKEFX0
4XCiiYjU2WooETBNixI6hGAdXq5zCOuY2l3zDQlnoY2pzGQSMsH0PTugqq6JeBJt
mCmAoxHF5v3kNti4r4iWLmQeiZ/VEsh2kS63WqzUBzMZvERdDNGrPVOr0ZcH49hR
rYwzCpqnNKi3e8FVWwss3tqNKreKgTGxDyTnQzJ9hxK2PbL6XUJfSwz3e+tSMNgv
Mq+xcxs1h6qqtl9N/+Uy8e9j72ME/9KlS2joC1zlSI+RgQ81ULml51DW8H0UTk8t
N2oLcDNn292ZYzWAlxkXqxbdptOl1UA+l2slUhmAm2ZLA82Ol9ApWf95lTqnQuh3
b+E87+AnJK+qb9995VnfIj0uVAIDc2K+m/bu96nZxaDpq47K8Od+i81Dg5iJQbJR
+vyoKTl5IpBdEYwAWlJWWxcB1tKPY0R6X6dIGuLxD/UP5RYetWj91MqhcWL01kdi
daM7EwRhnL5ac7bInS8wHSgfyTzfhSazxg4WOR9v/JzwkCFpR4qdcmCI1FLHcsOX
SCQdtsGzyfssLgb2iAOsWHGdkhwu4n+LLEM3ayhlidZAzfUISDmbXc/M383FKRnH
YDv33KoicQ4cYdXu0I3AXIRTKhFPFpV+i8l0P5gWIuv7RnNpMyUYmfrbjyodxOe+
Ir/NrYO1kcAfi2SumqZhpv7ExYvgVuQu6kwzPrtVP9qmmyVDw63t3zBlvMEjlnwD
DdEjW/HMmKOYgEzdoMBmEgmRUluO3zJcS6vO+rT4Ucwd2x65blUjIwKsMjQ427tb
xcmL8oN4MvLPPunmSz51nm3VBtvzSTexVPd4oZCCELLZ1i6qjEqgJ6HDG9RDjAnD
f20oybuUrow69GaJx4/UD9EUPygEwSXSpb2576oXKQzxDWO0b3fyW0VXWLzXzVpI
Qzhtpg+n7NgqCkxWSsHZ6g4xJU/YjMjTtUQbRnULtVSageADFQJV/E53HMzxAauN
JdbhbgL/hYab3215p0aB0Ao6dKyyVHyFFBMBex9slp7KfJ67zJs6KLbRu77jX2kA
+YNhqqr2X5Ui7FeG76Wpj24VlQ8N1i3Lrj747ZQWIfMOGTJ3J+3EvJlhYUL1nERF
OttZ7oQGe7Bv5zweDUH5YpTJlOjor6RDIFJjYxsCz93wYZz2t0vDUib4/79ZwnCc
5z5niz9o+0amHG1ABNbKTtArPElnZQovc5g/zTJZejTckLpUFh3OLRrJsCet99y5
mdG0VZ4gMntnww55WhBxKrHJRUsbrpnliexPb38Yt7iKep50+TrgzBxBRHYBPfWX
Jeg9KFUFbnZpjIASjnxDYTqCre1RsleGSVfukaf4oANVX8qEAraW2HadCZGtfiPa
6r1RPgJ+qViy4YAwgYJlKMH9ZkQehHPSTuDESE744aB6aak3UTLFn97aQ6uXY3hB
ok4K/idGvczCXD9TDJJ5h34i3QNLCP/BHafAsmYtehfdE2w+fgOugRurG7leu3vm
F4xaK6MbzMAImGfAuk9BJBmGisopiL2oZXv03WJwKsehCSsojBLLLDjkC5su5usE
9L+4/hf8PXiwjiWQ+vmvSG/uqHmlXQMtLvyt3bzzy84mNuiewNb36VkSsb/H8yln
cHmLgTYyKAIxeZvB9G7ctq81E8ZWnaUk09oL6fhpWZ2ApOrDvt70M/Q8nVdWzOFP
ksyKYGY3SwyzWlfvEQF/OeE5+NVCUe0mAQwbwm6DfLgbDGZmyWkGwwl096miDvYQ
Fz299MXB2KXYDK1FD37kW07PFanazrlFjYjgVWLX99aTEGVtSFV1NbabTuKO12Bu
MS4hxSHRVx73WhoM5PKEFmMeu1tIscGyzXlz+sys/8m5X9RUgY5PX8fzqMLB2y0h
Gj98KAMMSS6qUCrxtiBwq71b/n63pXJ3AHcy3O8XPU/WEHd/vUyWqTsZ82PyaVpD
SBY2VusgsRWD6zfwu5GQ5pPHxXVL+83vFp9zkwz7BiyQAovmhyuRJDqpoWtsSkTW
G7vGdXqnGaUyehX9Fl6m4R272ylPW83iBvG2w0BIiBXwYsScx9j505Hzg6O6TyN+
jAJiEAl4GyznwPRJl6cBe2VZ+UJknJchhIJgA1E7+9YEBB3ttQ2W9+tmq7O2LCG0
disV+W00nII7FArTGLYfjZa9oiOL8Zaj2hS12Vmm9DAwmg06DhI2tB9E6zMD83cr
JANiHZLm/tvjBdBGPJT8LmRwXhGW2sP/xLGht7DmbMSHXq2nAWpy3R5ousVtS132
YL/V36D5gU72uHrnOU+90O0UKX0Z1oGQFfQlAEur+Sy/Maoda3V9Rp61JAw0Ed5g
01gBGwKQ4xjk3czeed65hYdo8obDAfv4g1gR9RoXAzPBaml4LGs5GM4g2j8PAmHs
ZdVw5KrSAIEegvArgk8cqoNiMnBYCFDU0Q688E7aOzzRnJW9r4mBj8lQCUXQNiYq
3ybla2V1p9wT0Li6MsnotLJJTkzTQ/B5wfQKiyytrPUG5+XGI0Ysq1J9u2PmUOt3
ne0h5AqfgeedbYowVGNrRz40cmsn3er8+hyjq0z07XtRpb2HNonZlMacZb2TcBns
tvmibMKiWt1wKTcu2Z0Qj8Eyc/ndvaJ5Sdqeiw9CZXp8QoujXx43owfYM3mgAIit
h5udVxCHswnXyHh0YachTXEApRaMhSgqKyxD7Cy9AwCYlB1mqkAeiDE1/AyaLoEo
zA7eKrJ5gT4r52Y+QYWaeB0Frn9wa5VHxPsIpcFvTTMqHTqBd+YbfpnGSWIiLwed
wkjrufoP02EQHbeYdCm2mm2WiY4rmPBdJmXf7ux3DcUZpfgyLcbpyas6BDXmOmwh
KIdolRlXV7o1ROf1kkLt/93wyRUHfk7VTSKm8ekwttQZjXUbUSnF2mfMEYUJU7ba
kT+avnIKO62QuLTwElrh8g+QIOI5rD+4dGKF7R3CED6Bwt2xXGGO0bq3o8PsJ6rS
Kuah5GaAoRYuO+tkW7IFV+6rNq3qZgObtS0lzFrh8XD/3eigysPcZGWe/Myyxnzb
3U3GjGXl6KK5ZlRb6MD8trjpAh/Fo49VM3A2G/OjcW8u2IF8JD63DtoGjobWKPQp
qQioAkIELpbfIjxcd0Q7Bd+VbpOsdTE1/kZS31kWkR/4LdZqgEbaSzR4idZixldy
jUp0cYj+H4RfXf1VIgUJT1zCcRCQIFIzAvG+81zajVXHzlHEM+FuJd3k89FOiSa9
IJRPJ8JMUqGKcAIEaSin9l3AMcc/e32KjX+qIOu9ktPna/w0uSnPePkociFBBfNW
Z3f/20UMpVUbFZ5KqaN1dK5ivya3UFU6gx+2PpbGaLRMbjnay+b6oGTZ+rkWSjko
Qs9ZowkcCI7KXC4p1hQMBy5eWp7O/Q8BAu3cc05EW8sEQVQv3wu9kxvIVzdGlXFC
vRiWkQFKEby+fx/bdHBlRcL8c4A2WMI25MOcy/rPeKeER5IxsqksXpIWgtsQUwQo
V+nBQXz5UHoLCKtBRhO5omyxmIlKoeC2/IxuPDTDW3pWqTkMegK/5iFTarVClla8
latinh7fWnFVnLgLC4bpJC+1nJDAjwAQVQ49SQCCaJTaZDHU2pMCgaTlOVPJy0oi
+2OBX1A8DaHDW8/b+PY6tc2V/vrIqEl5I+tH+XLTVTife61pCCXIIlfomELqQc3R
VRzIC1HKSSQaE1Wzn5QzQe1D+H9uBZaIQpMY9R+LDpdh2p5lBtmIgVeMLN1H2j6z
MDjH284aY2wLgE1rjvmTZRQ9dn3o4Wlbp8Yq6Edymf5LOkKr6FMvqmU7xTZeoHlq
RWdLpnXUaWA7Qn6Hg4BF6f3weGkVBT3DMOjtveQSNvz4oYUeDOtOu9aCX/22VuI8
SxA2EtX5usy9ZhUmcLWsYQcL5WWdbTN4WZh3Ig2Ys0srbPKtW7TnweLEccp6qFyv
vlev5nJyom9Ipd63+7yT5c6AjOy4kavxeUR0tX8bz10WyEub31QIjegjwshnagW+
IOOsoPUNN4BOmXaefmjg7Ja8en74daRU7XiAeVsDBvydJSqkcT+Pq91t3MI/OISi
AGdFkITl9APh2yulE3NxdAtET4m6jOKrzPpI+VRS00bjwjg5aLiCv9KQ6ga6RAyJ
XZliIjkxPv6B+Gmjn4EGHt23dqNR20eqVFf63l8vpUSRpPlSW4Atzvx3m0IZ0Pxm
ee7dl8gBX2zaymb+d6dD2wbp/TBewI70VzK1HFU6Ihv+cnIB4d4lQYn54DO+kDM1
RlyqGy/lCkXtANCIOAxh6hj2QkYBKyrpoOeJjPTFsAauZy6D4IC9pUb4E1N/Oquc
BsqTJUQHsrGXtOLbOlqtBS8lgilG7r9ALI2Yxx9yvhkzr+NqgBeh0YGvdOKOjVLr
izJ/lSP8tKd5PoztDpNdyyMS1oWQceHjSbf1kKP1BrepPMypYeC6XF6sDwCi57Tc
7rOWxz3TckmxPpspXs0bcJiV1GTp6TPwsqIARd/w3Y3lXY4CK88UPQZY9tfCNeZ5
z45sDDbPjDI8geYaUrgDjpYzWAxLWD5qI9SU1GERUG0R6B3FjZ8m3IPOMFct5aIU
JFP2mgctx4MukFRXM8pCCwA1VmYIgiF6BLr00c6qWtObsT/porDdE4ybHcitU3nx
5Dt3QGj7KJ+ZGzeHYATTTUE+fN0XIUMFyfMsntTNKOk6Be8L9p7ZLqSZOCAQ1f5l
1kgt5cdIfoEL6MLheFMeMm63BR3Sdt07+tDQTU3hxC4pNQlhn2YjidJT+7UrOwt/
cuUv5BUyYbw8+ZbKLnloLeZtCN25IPG0mqEDhPyRfnKq33oUtqw1vOXdbWQ75DHy
XFQ7B9dNG/6rfubVdU0Ti7lZqYln8EcZiBzraFZSKKWwDoFBn1PtYpKtP6QfBWED
EbGQhba7aaoVBVWvXvR9zC2wDPy4a6e9Sm4jJFgBNC1rG/0EkyG0fluv/2KqPuhi
CBzupHaP1uNSggBgeQdZf0EuONDEpzRDrAv/vMR4RgjckSVKvcg/KHXp7HDWPIiz
id+PmvSqivZwPqvZzijJh5ymGKORn7eL/Ai/HwfmlhU1/VIAux7SXYr4RtFbNnCB
lJX+40yd/G08CXo2UyMMyQ==
`pragma protect end_protected
