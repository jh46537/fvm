// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:37 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SzYQH7ZeGXdV5Nwc51bCP1k6auYOwsEarBT8LB1IYqj2Njt+IrmN9nyYi+SOGE4/
JmR5DSu23AOA6b6vxzyAVbcb2Gb/Nx1DzBtiwFvCdngsjgNK9s2Y1BdK0UwNF6o3
8Lcc2kVU2a891rT3oPslmu66BfRVaks0nih8Xh0+ZCM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7296)
Ij0SUiK+8Amutyq9e8Z23LoJiAGF4YP6WADZORp8dV/MtCyCIX2Z8PZb+E3YcGxs
BVywmkKlngzMSu0y3QCxfnBo9GftXvTluxnlUzP/pH4P444QhjxcybPjBBD/dlEA
dd0STWo6zlY+r/DMrn0KGE9moRShN1pGoH7wOsTXy7Nu5ISerrnwF2M+c+7ncs55
KjrNlhpdQo9PX+07n4PMXWpgvZplLjNh5sa5FGjkaigRG4nkg4N4VOv/WmANkzBM
wIYS40Mg/WhB7QnBG33y3JbVmfawrms11kqoyEHzRuBMuaMxeX2EveszrHcgnDHa
v93x47bzws/Cxgs/oPcHIv6YsnoFySGcbnJkm3mmQqyv9eVg1R3Ncrpqzs2RfBQH
l941ebM5jkoXRy4O62+1FNfh2q5NUtKomC47zQXpX1F6qtw54vIEB8ejtS32g5yq
2libvsbRxVPwq95XTuF9W0R5oPVf3vqqTwL0wrPb7Kzu4AFin8kNa2alCCv5a/oI
fxyC3mxKnpEB/jKG8iMU1rwWmT95xYvpC439laaD0251282l/qesXob+yCvxdnQe
Q/oFL91b7A8EBAtPQ8HqpCMjLee49i737w0Gy+iDM7ruBioqmBa/tjKtQs+lp7AL
5wYjPBoxfxtptHflgHS0TJMVMMdpooO/0/POK00Wu/nNIg4tbiQOO7RiueGC/B3e
mLUVPexlYMDNezNEqUGguqAKGP5Q4BausVSTEJejazaXJGETVzJiG6kgLNcoOjuG
DaA15OhJ1zDYTqgLG/sI1KSIzFHrUMhuHdNgRNC6JvrPoJeJr/FkteefkEM/afjm
i9eRxGzoTW3YF2nrCp7NyEUd86G0axc3/cwZSuYxxuGrjzvRl4Ocx/Q/JZsOieRb
XRUsdz+ffWDDMIlkRiCjGhxpsZpD2qs6wmNYu/js9mmiczWYmLknI/0MdPjL8UlC
1ZelQC4feYRAZFdGayEPUAI5/qgVXUNyxy0uPMZDvARblvarAEEd5z1p6GxW6enl
U/NZh34unzM3+yvjP+mdwknUES3/F2XCQ4Gf4oMuguBWyh/oyJ7ZUKMRP9bKRh1B
5g/3H/FuSz65KmFNa4u9k+kXJs8eIaf9UNpjSxOc/lvbleoiRJQbuNCRhqogZ5pp
Sfkisd5U65Kvw0zyBaa8L3rCMRhEzFpNAxN9WKkBqJkdyg6I6QxF/YhMlVlSxaO6
lOcJYs1HTjCqn9Z40IGKf0juAb75qz6z770mvVSmb3+jyXkLoaS09/s1O+6bPy9Q
VVSD1fMFqisuDKzdxkn79EpPp42B0mutLznRhg9cOJ1+BflyT5F9OC32JuYQXX8y
zEVM0jIlPmwbJuS/+cSXG0QNaNlobZxRDTAISE8vOlrO211pX2GmagZwjN8tTCW6
kIZkPoy8cSERF+yfRc55pthXJCBd2ibhL0wZJw5LOGfwI9UnYQwjtyZtlP0pHO3w
YEJdtFh8SqHOTM2los6mdHVumVPl7uE3DbergDpl4LL834moxz4c2+pD9qu4301V
ItZZ+YImgJqrrQkklY7LVMYGm9Nz72zk9WOvzchB0kKzd8YwWWFb4nPHp7aNPGJg
y5hf+4spmgifM5WvqpxGEefAP8NVSGMViP6PE+2tglFsbrmQue+4Qri0HAK6kiV2
tDGrh0q1xYpi5mKha2Xzqvi1UO8+Lzk2YvQvJ8fJITIxCMx1AG59UGslaWZz980N
W7NQk3Be9ZOOBzuvNeyINGyQEXupYGr1Ee5bZVFkeLNnWBRTP8519Sqo2r4dvAZ6
9l4vwKf8DYAo0nRZ7UDvuRKmfiZ3mHGPaSuK5gRMhq5rS5R/H9QYQDOVCZhnjmEz
5BggGX/UvPYerQFHmXCYkS1lBfK0x9MjxANA4LyUmYW5l+CtZu01zpF1Sc1dua13
AXKqHoQgtZrG3N+eFbLvxVJLrfo7koNYaU/IYgC/tjtrkHszXhRJMBoDmLFL6w1O
SWfiW3PzmbKqK1va6vgIdcvAWCQAB3GJp8GaacC3v9z+kFdN1r3rFRhO5r6Y6SlC
j43wMzLRmAMmeiG/n9j24SOmgyP/GSYDTJTQMnIyH/u7IWJ9qY/+E0mjVC6sj6aK
nHn8T2uUbu/Tkp77QKm4NlSE6sO+UKmaLlPsy3RXM0eyZEe+C0C3CHTLM9RWkJ5H
2K0vvjV15eLdzwm+NzS/g54l5315uAx/GqG6KzXJeTyV70Lv1KRl7LfloOkIjLSs
8tICvcctyYKfpNXnPgOaY1MKxF4GHP6EQ1zWxugXsmgqUNSLeZo6vE6bRtqXneEV
DwfmZhDHULW1kBamhDtb7vbi+MVE2A3uD+uaJqG4IZlBEPI0p2p5hBrUR+cnym56
COvy1LchFmAiZufvdOVLKqTHD4SaLtv/OJyEXkMYp4fw+szZsW4/rxUqs8zUDBIG
xf05j5FjQf+gAJ1RW3AnVvxcQV8Fqtsr4itigmfJyaUC6qW2aNucZzmQ8hivFMBC
yHa2o33DB5vRsFzS86Nzwdi4DcUTWTrufUbbEbyuG5nGEqP3xmJTGtRfRqEp7S+G
VjBukdO1oJInAK+5MET0HzGv+sG+g/lwBod1bHJMf+wQTX4jcUwF0cakDoLZDQrV
kN1KMSW38guwl5CgyVhzp+8irnSV7794/a2YtOkWoVyfsB0CvqUILurmZshlc9Lu
h2ZRAthlsObkmxreU2X5GuwYtBzpeUvGaihldVdXMznzhYcSnWJOLkPs7wbTjdVI
JlMCYHvOjd/FoLfMR7jWpFLnj/q31EmMTqE/ZGiZZ+ZpcTLdqgqWm1uc8oQ3vK1j
0KEWq4aILiAiF/b51IAEM2gbCWS5Wq+kYNEM8uWzbzBuY2z5VHdfFI94Oi4KCwcA
8W6QpCgNLNt/tvdp6cQrKRdbV5xT/QOxwoy4hzKG8bnGd43wrO+uAy+mtvxdG4wk
PrCDAeBA8UYKFtiVkgq3TtoEdfJQyM/gjVy6ob8uRdFcW+IeyEiJkb6CvLtUOTmM
a9RY/h/YCPjUD5t8XsL7FrPFBOsE5czVQYuhWbqXEQ97zofyIdCbxsdPHp35pBOu
JNFvFWH8IjkIK9EwRv5wIBVapr5fj0loa1PQqwyqf2HS2Emb8dorOuRRwY/o+Ov0
Wswtjg7sfjrPf2BI3z1XMAhdDvuhWCpjnWh7GQY6ax2Qub8wqPCIjiB5qmyV9gZa
sRju9dG/JwP3THmdOE5vnR/BkO4v65Ms42xIeSwyMbnuGY3tfWyBgqJnd4qhecoL
5utNNL4vw6PP2ZaOBdcpXdwcaJkTM+1FFWnt/I3LT7g9eHcnOC8fpxZJ7vm2x6JQ
kg0Fu+YpuvjD2qIXMrMnDnjvI0i5YqyQvs1seXn0uobR/JioP1Wrktn2fmHeiDR+
jXSn+b8OYqdKpVXoRd0PUEfDtgZcPZH8qspu2a97/kBmuPMzw/J5hvutHQAW4P2L
Iw7gRk8gycTvCOjeLIZI0E3cVVC4rls0gcYFQ9dlKdp5q99dIufBArR+MgbyIf+Q
UQwjNcV5kPmUyk09xBoPleFSqSMGBQaaq+CsbOZxy0GJGJ9FfiCsUq5WCDQNb+z+
QiNYviDOjNXRNSijOdF5Vv8m87fHFNoK/VSK3Kata7kElWelku3xWKKmfUFfUIBE
hhb6tXw0prNHPr8r7DsOFV+qyNH1c48MNFh/mTmbMmjji/W3wxo9wMOipXTE1gGO
OK9zHj51LXos2YDTIXDUGCwbS1JzM99TqSqwE7zZBIltATTF+t4JPwhiYLAj7eoL
dwBQJVnucsiOeGRbVFIJZnNSGBmMt2BZxd1q1hhbLnXvyuF0NCMzCLnvTFDSpr85
62ekczh1M6ZSPQDedHEinSji+VEyqeVdP1p/OssECsZ8lts+PwKHtH9Hn6K3HMF1
CjW0i+EsmkoTeyoSQE0TsmZcet7cuctRg+eCCra6AS+AeRok7Ga+5GmGVIR03HVo
bbVlM1tv79Da4KEC5Tmc93Asuz+7s4B+BO2NqUP0x3/KW/HGFzuR4vPx72f2VtYA
dfmpPZHIdZLvJjH0B3fc3hUEizDGGXfuh1CWLRG6TlI8FFL3pMSmT8AOzqFzO7BU
L8/aFpgPeIXAGWRl6KEThCw2pZ7waYR6YPsHHdkpYL0VwZDZS3tKQVZ9dzQByoFn
ySnkHmIrxko7hHL+ZpsbniB5Pk59O6bUiYyp9wWCGmeWzpj86pH6uySFxFlvm/mO
WYgwOeHqpdbcvHy0X+ESEIuSJbUiRwqVLMtbsgD5SHmkyTsYjFtXT0jDm7ckYkKy
9Fml7rXxBIM50eqOyuM+j4gs+yxaiBEFKbVdeaA+aUSh3v14IEYitcY+olV0PJ7g
eOFUKYh6sfWAsUdH/zbnVH2lq0m2pdUnnJRJkaOZczJp2aejmOZFNVS4WK7VjAFs
14K6qwmtIomgJduOubwUm1Nx+vn4VTovFW2aZwQFS557U0aLt0BfWli/FbJaOU68
T4NUPPXF4TK5uOOK4mMgAraysCQzRAiBLwYqTxC2qT6Arj93m5sXFayOvw17jtzq
8jwTzLgXNNIwdnQbiVflzeE5VBeHjlFXaV/6UBmeETdz8xRNKMTvl9613hgCzJHj
2KNZdoyBsdsaW14DSBhAcwz3z6kcE7f0TZb1uUreZGAXBwcfGEaMvJfqyJiFso8z
uYrbJ7ODmxz3JT4L0yXZN++KPPQaQhYO3GG+5MS2lcFBKCNok/kIBnF3DLIZpNlh
b5gBiJeEVHLkutB84pY6H6b0YS9tUuOOAGBv4v7nThAh7N6bCJEsQBPn4gmCU5ct
4rmYYM+hiH/VaMGtAxXAg0Ll+QDYwY/ryqicNuoF+BYWMsqvrHiyyV5yxgDKUImC
3gq5VZyLNcxAuLIla7vCODItfuVJyb7/d8dLSg4YqHhduGrSQpkUaPquXiBthVfC
2MiIMXInGbRLFIeL6C98gn+jirHR7PJWY9eheIsslpGAQGx5Zb22toR2s1AvGyld
+LFTOmWz874MYL7nYY6XlVBPy1/2pFnSw+knFiW7tCVlGqolDGPlv/5HMtpCVxa9
7GpTYA8kaLZgg2a6oaWvtFsRNi2nGB6GvPWvlMXGbbVdyXk37RgjP/Krpvuiujvv
wX0lodX6zoWvcGhlNsbT4CUJFG3mx8xqUoWZaRrEuWlHLSawfIsfvvtdEKLzKJ+j
viZ2sG446Dk0+TttDYXXVfzKvfr1+SwqnbuTeRrHJppQFl8DWn1Vtgs6uKCML52R
6K9BI+VXF0Yk/jnbHtr3hHBnNWRO2KzO+UfwgR2TRi71vZ5h1w3wqxngT+b4RroL
uzaer6IIOvdouzzX76E9k3msBFo89bfUk57mnf1RQLYKZohb7AlK4MCijlklQ+04
QxwE/AYMGJtXj8f6//DP75G8w/r+Qqo/Nvsj0E5V5Jr7EEBk2qY4uJGUi+MEBhRj
iW9YFuDAiUmkvKE3sSG4Xs8P5dsggU0+IOsVd7TGTbsGVXeby8+mhilZyXIkB1uU
YDyhyrn9JfRQkJoXy7YuHKLF+I+lJK7YBA1SN0gnEBtcWWhldOMtOPvim3xYSP9u
aaMDqyUK8IWzOWjsGew+QsaOUKbYxTzRaoGzV/V/UpTXJexwbXaUy6Uib3BD11l8
LgnFi9YFWAuquATVR8OMn9xaHVp5HC94rCwPjU4cAUcEqtWkwjYZu/Bt0/0ZAt5o
jwcv2JU+PuKyy17IWsfnEAR/zwbDZkWqimXOOwZq2jCfVIUmAlvK+QS4Qe8IjOO2
7P6bP/b5VtGhr0efnzYE/r/haOWZicRg/EyVRBlnPIpIa5epb6B18LuIGD+Nfyuz
jEYDb0xI1cuW0VoXvm3+y2DxD6yglz4MvKpKE4hwNMtL9qyDVEuqr/BP2XqGvmGv
+DclZ1LVWcPBT9cJ+0Kuilnv2MGr/VEPJkh4QL8vI5mXptvWEwxohGDXS2AC/BRi
7lUPtzgbRBHUem861yKf62N0oET5CdL+jrQAPnN/Sb3CZC9S7PjGnAY+S4hrtQMA
nSayeeNDRBPXplS6rXw3A2662ni/FzkWlrhjwbsQbDjW0Ip2xV03P+hMthV5IIvO
sTkTPpGBP+oB7nPdUiF5k++AFwApx8zDnuDFLur5AG413AuksAz6QfP4K3rpRefN
JvLG863kJ6A/RVsQVft4OifumvG+mBO1tMldwmsZ6YJ/fYCOx8vPSO7Et+93XhQB
f1NUsnDs0RTa0uC4N+N3sR6/OIiz2IWb2vuY6D74trjw2SSQNndU6uXwY2rBCnF6
v/CJddrqdkp3IrjU0s/1gsRBHUqQGIylmIk87/WJH+0TJ+QnzkaAdcja9X6Atlbs
ZGGc55pOStlf1ZlpOJHeTtrnZ8aE6Y6HSHVCf/obL3iHghlA++xhd9kJQ1VBZvMg
WnnojBLkz3BGcvG8tQeyxPZqQZ90PnQ4Qm3Vvhs67NteOoGSl5ZuOuI1F2rNlyYg
8pFFUt2NjNRrg8JP2IoR23RvGMLnKZ+LVicAKt1LHM6lRM+sEipqbJ+j1jwcz5jc
USLN6D1A/vc6ZxBVxD5I+s/GfKq5HL52K2dalI9Y+Ds9T7abinC2jyB5eoCXt/zX
qYIHU9V27rifDXjcNFnWL8TU+/uSkD//CNJI3EyyRJ2OQ7O13Bnm2Lihp8r4kbMR
jEa0i42WR8l87aQJSb5MvpzktfkqO98e6Bt67ACzby4TPHDKc/9XDuVoKWvhV5u8
0IqS7kyomCs9t4MdDaez4UrkFkwaxJ57x+5e4ghMMauiW79injW6rmpIt67pITkl
4U4ng88pokKt/BtrZ3a24k4Y39lZcVu/cmBnqbN6jUwq+4uXMsyX57HUuiV+Eunj
e9i2qN/amVPnnwa5rJKlTQP+WudcYCKG1eBamA34RzeMwIANxUGDWf68Fwa10nlf
sQtwIeoZ+NF9RSEdQWweoM6sTGDGeWCoqAzkixHEocX8DMjlRcsX/JNReROEBvUO
la2e54Lil3/LXgp1nq/XCISpMh9QLEeA75+vFE9nnm0JGJYKbfjECXta9KMZWQA1
FGtaNDcWAoBhrqZBC4gvMdE5jDk/cqrCKJ0ZaZWM7tQiJmEd0yVuMrsiKkN0x+Q3
qW4lZ9xJ59QzN4UN00sNPyziSaJDIxAvBpK1DchoXK9ZV/TXLdC4n68tgWHjexU0
Qz2g+eQoCHk3fNO52Gp18ltvJfvTx1PiCGqgMmqPw95eEbbVcISKsoMXAFvpy6U7
NcWNIrO/FDJSByx1oHyBLxE3yc9oRNxPx4NL8FGavxQhqhHBhqQ2G2JvIHRf8qxU
q65U/V0AM5VCISUhmbR8jiaC7ciamAZL/1na6YuCo9bqgDowUzIgfx3MPq9dR0ro
DiRJiUXJsCD6S2+kDjbuMUKU3B/2kWxBnwYScVhE2Ss6iByEVvJHBkosqcHUl+13
CEWcdcE0boRe9F9n6MgV6oH5eE/BOmXVfNktVxN5JhbpevqrDricPFaGmK1f9Tth
067e+dE88ymjs3QjUTIRraTgDHclsWJHjN24yB3iogjn8PXRT3Cx141BjUk49Zc3
XOTDg5fJ9/B2fMiaUxmRh8WycYwdTaF1x0ZyqbBL2Kl0ItylO+T3lwd3jYP8laUJ
jgKgl6eOgQUxUnpNS28Sf7nYmecYzc+K8clflTYuoebr+LoYEPJn3t4kp+UsvKK4
aaWFbzWWUSELXJvH/EjQeq/u0gxd930mjNHdYu+ooJEGloPTbbkU7paS6AWhBM5w
sLBvUxbrW7bePY+om0tDDqJk0nuc0wMg7t9anlef1JMONWijgYqAsgmBhFBHciQE
kfmpcXh9hgq4Wl1bYUxPouPRiuGDcnxN4z5VojTOihvcIBm1hOlc80eFFrMHj4Bn
Cf6fcQ5h4yKEUyOFlzGrZR2n0sGMEp+EtgEu1B5NHmwencs5Ldr6rO8UF5WKxttO
+F8tTsOPy7MXyj3yL/pKozByTlAcrNjhtB96/GfM9klEeaV7v1cMrSX5ojqM08mI
e6zvPpH+gXJR+YPqBe866gXf2ofaoGuAU0l4KTgyEtTmn47ddJ423IEWc1U4wp1K
QAKt0fOpkexJuJUSeFrOwZc+iO/NHcCXY4I6L8ZX/aZnNkimfgFl5yMHKKo/9q3V
XQ1icprTDvknH65/s0JElrBuSGYVV8qU9gX3WVGaZuAdAp8m8G1kscU+726XeFYO
eLXeuyydc7nwGxvrIiNHMexz3u8czsYKA6FZ4tpnzJOx6oHbD34xBjYX1Exj6ta2
d3GgJhcpgGbQ8LaE/QkY5aKR/47TG8ytNFn1+sPrKF144FX65kn0Vs08zjczbWwg
y3zIdxcL1SNHdJhW1mpOxAAZJUMX7vxnHCVAV8jdpzqGfUrP6EW0E59lf+U76IwO
2IkU+T1jIQ9o+4qf/DpMoox3gQMLiD0nWGi6DgUXFyz4z26R3NPwqF/sHtdm3Gg9
zb/h7azTNBpbfRsJ8ZYmWmnor+JsanzlLIIQ+sSra+N1LRYTbiJS8OUDwIVP7cDg
f2Im7nIl28LuEiWAozMOMiIyNXxa9M6LfLFDcLSw3uDrN+ybRtg3UwqRJ0NdVjtp
kDKUPUUWlSMmkeZ9lNf3tFeKC3TEkCOZ/pJ5dFs7Sb1SKT+8Sk6oI+/hFL7WHME5
oR0RSwv5ckrbvYBXhWbTAPmmyfDgaArGznhSDVwAzDCN3TWd3qGUb6U4fc16hc4v
7l3CVFkGX/AFSpLr1mK3gDgSFKVGaBiAN4DiA08Bv2BWGgRBOGWEN8edpSruR9zl
zIJe/QLXPlqzlryFtsR/jyDIanWmENySq/G+TO2+Y5TxIz6ANpXoPGjjMXd6yKhe
UZ795uQYDDTYBHtHUiR4YhJsl0++AfatStF2qiXpw90+X2eMLo9ep7aYoNUxD7lx
4yvyOmjBhiG6IrKgF46j3RjfVLDpUj9a5HV0jaTCbBEBalyHGv4fSCkRCSl90aIz
U2qazOzJWCvjWTvJ0P3bteImFE7vboToe9h8Hi5dd4RNv+V2xCmqwwefXJTasIzy
7ymDuRtuzYB4hQ4NhnN92GFN9I/5YO3VHOeSc5AvgTpYf1/W8PzX/4gezMmAbJv6
A3bPlVJz6j1btuceXL9FV47Y/Xjy4Lsp1tSr0FZtK7nx/4SFhbqKOjflFtgo1Pnz
oeueCh4LKIltzvWnns/1XFVRS/fjEpXqZ7pCNS+bOKGCRDFCF8/z2IcrfTwX/cPB
uNB7+xXPR6Xu5iXG+pXhI2JhA8L67RcJQL5ZasDBW1jcf8bQpqJpPMyELF7Mj1SW
TEUrPhJGgBfPejjcCG61DQGHg6PQlOQF1vk6o4ETqaLDlg0emrF4G+aVGzIBXgV6
rVtVKEBchEWLkaPYcYbOwTvSwh/DscHPsnT7fb8LF64YGZwm/ag/aa2m8NbvI226
LzPWWAtq9tNvzNK+6S/vAl6E94dMyzq3X51jl6A4pHlKRCO4bZ7aBAH6PKUlU776
nk8IsnT2C4M5E0nx37dfQou/ubXnE35Y2ohiuB+ZRXdVNltm4WBM8FGTej2sq9St
q3IoUoktsIbcUX9EY3KmjTadTmvfURXybrj9FMT0nXIwV6h0wh6tX+NzF7UHelsx
levD7OLb8fpqNKLn0IsnxuSJNM8pR65ea8/CuQy94wcjYZBn6n7bP+K+WE+fGtJT
MnQfJnEjorYE7DfU+GJWdgEmFkqKXSM18KyPU07Mv0w6Hz6PbnkgQyIoWCrmFbA4
`pragma protect end_protected
