��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}�����°ȣVZ>@�#�����QW�|�i����#JM[fsW�Cu�6�9��U�?��#�+�r4�B}�a�+�M MF�"Ҳ��"txOX���q�I22J�{�|㹨�3�x�w?�Pbx��Ԋ�;NK�	��[�\��H�@�.��y�GPS���A��,�V�l��O��8bz����>�@�-��7������M)���yg?$g,��R�wΕ���z�`�O��ogW���~�j[L@�ɗ�/W�qp�����8)f��x+Q��_���ޜ���q��&�v�89c������>��QN[��p�-���睌OЈ��>k�+�ף*�U�M+��Z�wS�<n��6�J�ݢ0Ɗcl{ ?�H�����_��I�^�V����>.�pt�ʚ5�Sr�K;�g�\��}B�T. R4���j��}5*�F��(U�)M�-�
ah��*'���r���?@�F��*��?�;Z�� �ܫ��I⳻�4����Ӑ�k�������;��f/3:�Lgx���ZQy= ���$�y�_�he�t�&�a��I�K��V�XQ}}� ��,��wYݮ�i��x�t)�����(ū@5�Sa+
ަi��t��A!�:�k�u\'L߾��:�?�"e�m1��,�����E"���v7�T����1W��q#6K.�[2����'�%����@2Z5���2"(�ب�;fY���M�를z ���{��T#����àA-È�E�N7���lZ�f#�U0��ÊF:��
�H�5,��)�ʦ���A���rT��X7�bEw[�Ů}���������_�:�4�t�CC������?_��kj�b"֔<����p�i���œ���+�Ǳ�V�cT?1ߔ.�#����Mf;cޏ?%��Mr/���w$1�H`��_��l�E��0F����g�;�tOH`%���! ��g��8TT #�ڶ�����Y�\���P���/G��ק��Z� �97���T∙f�!όK�D��l��iŪw,|"�]�DwVi��u��I��F���T����Ќ��A�p>�?��.I��>:�y����[�z��Z_P�4� 9�ؕ��A�x�i�� ��|>;V��ɕu9�|2@8=�뾇p45¿���m L:)c:n�W=��rP�6��a+~[)w�P�:� ����B��2,m����nw�=��%NB���G#w��v� ����n��AwG/Z�dm#�O�̗�.�L�w�Iy2�k��Z�'!ʳ��g'�{�D�D��?����+WS�3gl(�a=���M>lW�	�"Rp�.�>!lm焮����l�{գ-G�I���%��57H�0)~�XS��0��vv� L=�֜�B�t[�%���������?u��(-D�eqn���d�4�c���z32��Pe� ��b�bi��8���K-��'�y�u&5Qh�RH(�h�z�s�K�d�J���t���/��>C��S"U��c�x�E��r-f�
cO�
�j�*�?�y�o݆Y`PVGD�[<7����8IS�����Y�*o��;�����6��|��UuSݧ�o�
�{���YW�;F��]A�ZY����<��iG�(	����
&����Υ���S�ׂ�	&�z�~3�U<�M��4�ƣ�a!W�>��������� o�[WhףiՆ����F;�?��QEg�/rB(a�,ؘ"`��KġR@��3S�d���y�>���mPOL�0�1� �6�/���!J�JV:�IP����J�������aG�"�;��fq�0N�Q��ja2������K���<W��S�c~TU�K�~1(G�w�J$����g���0&G��J��/���#��K���e��1��h��FuY�>_�ڱC۱��i_q(W%�۾����1�h�rHYp�a��W_�(w]�Y>�Ǣ��I+[����3�Z��e[� ��� ���ݘ(oyQ��Q����M��i_�c�N��\r[���ie��K�#;a��X	�}���ḻwh��9�Ӆc���5�CPI{p�]�F�Yf�n���6����{Dr�Lp���͉�^?��/��L��O:qhf�V�w��rO����6�X���u�Z�kQw.����gYS5*Z���OVlMďY9Lk� h"�~?�kwD��P��ŉ.T�������P��MBP϶���F��D�Ί���-�r��������	�݇��-���Ւ--��k����t~��̕�+M�^&��y�U���i[���"�09����_�s�?�w��A����{0W��/�j%��'�W�G��il�������&XH	9_[�:w�~�!�k�ȯ�0�c�jZ1n�!���O��������[6ܳ=u2Ρ��Y��l�_Y�[�s�0�+��(p���p�\��SĚ$���D#��H�&A�*Js��ՂM�Q�܅E��d�+�u��:�����"Y���u��l0Hf����z�o{%~��}�DC�c3[�������l��H��DQH����wK���V4��Ėh72^o�h������I������Qu�p�p�-��ʚS/P���l��*,$M�n"�2����}D�I�C��}bv,�к�GL_��Wjjƛ�M�u�І����e����[�?�$/ U9�G��p���/!Q�=���68�(C\'���X�sa�xA~�Dj����ҫ^�d�M�"I"�V(VnAN�56�sV%���~)9����Fl2���'��@a~!:���=���	{���U�P5W�������s9a?>@���E���V�e/0ȆW=,���E������gr�̕�b'�R��N�4��LLU�R*��d��|�z�˲��Դ0��xPW'�uLp=J���[��K�c/�JY��O��w����E�4o�I�,��S&<��'?�oy�o+���	j�Z�z9G*���6v$�(PL��}��A~ai��l̴2#�6��݅���7\�P,;�jA���/kn��QY����Nҁ���|��˗i7�>6]�Y��C�J��@����+�#V6���#Q��nt�;2VfS"�Η8@q�5q�(��VҲ�ڏ�E�E�.B-W��ȦW�i�[7���>;�﷊���E�����ce��d)���p�{X�n?�'�&j�$�E�
N}Z���Ny����u't��0���dq{j��W⮻п�B�GSjjtp}>��P '�����d  �of5�n�(�l'>m���K���Ҥ�W
�-��t�n���t)"� X��u�SMa�ٝ6��KE0:��UH�� ̑�.J���۠�'`�����{Q|7�<�R�z�i�O���j�N�sk·i��.T�×}�I��.��JR,.���u$^�03���`ya�1p~$x�UvӪ)��M�԰2{겅Њ�s�k[����<=�6�}R�^��M�����;�f���*l=�a�����咫T�_����	P��U���@y�g{�Kz4�E��$�/���2��7�Է�O����%�O�R�[�$x�L���q�!nC�"�И�bLM� _�5�A��+'Z�;��Z�� ���m=p��YuǛ�ß�,E6܈ـ�[��ۼ���a�\ű!���JFR�:v�ϲ����X�+���:�dp�?\��BO�jLd`����u73��rk*tn)�aBT-0�t��`����6�ڗ�`�폇M�D��;�I�������J�"���\��,f�ǆ�`h�$����t�	Ŗ�4�V�	��	V�m��n)R�Ze��ʄ[7������S7N��0|�i�4�p��2���B�pr��|2����d~���^ݠ��5�D�
ov��K������j��X�\x'3�GA?5�ö�QX��������`9l������r���M D[�����B�Ok��;Ҝr�T�������<0�k�K�Rk)7�m�0�x�$Uj%:�,goB��^^u�E�	x��Ȋ�ʣVP�m�S�"[���q�8#�<�Lp󷀿��!o � B�4��m��������N�>8��єc�e�ʘv6�a�pnE��n���P!�M��M<&ݷ�Q��X�nΒ����d��ג�s+�ʬ�Y:�Hf���ە��c��Kܨ?Z=�g~#V ��@񐴽�f(�^�{k3����x�]PZ�������7�����-���}���|P5���H+C�1É�R����A,/\����.6ܦ�s������l��4��(t���Ά����{�@$\Q�c�����l�2^��4�����(���U��x���Z!��4����7��i�˪�Sį�?���rc�w�4��[�r
O��J�!��w�&�G��6=N��3v�M���:&k�:fقr�_���o�����	Z,�Ez�5��cb�����Z����d�0�Y�%aE{����� �����L���ұR���ӔR��!V0����^/L1���J��g�� �v;�"�|���N��(}9]�f���]�p{�H���Z83R�YP���^t��d��s.}%l�7�j��朷��z�{�O�z&�ވ<!�Z�H��$�ӆK�����M����I���F!�z
|��-D�M�
�����*�;����Q&k^6Jy�"�&���^��2��!t�H�Da���p]Z�|�E�<�_?�_1Iڍ /���r���SU�7���=�y��S�8W��%\�J-g [��6w�u��3��r��&�.MV��W,d��}}�R�_W�0�ݓ�-R����n�J0����|d�8sE�b��6� ������n�Z��1QV�MO+M��G&�P�  눥�t����V���!~�d���@WiL� �[�t��<��s�2�Q�]f����'K�+�瞷u�����*�R�? *��Sg�5����C k,�6"D74�D�vӸ�Ŝ;k�dq	���x�d�M�����FWW� 0Omvߠ@ԏ8��sq���Ӏ碣��k�����1;���L�*�.��2���MUI-I����-�!�/�9�n�r|8���S2V�ԑq��}�ڒ�w������>9��i�ݮ;�:HmD�]@�@a?X���)�_�	%@un{�<����-��(��?�m��KRߨ.�OϏS�/�������z�rۧ���ռ�]o��0 ����΀�ߧy�u�@��.j®ΉL`����o�H��X�v~�g�ټ�3�w/��Dwڱ~��@�^��L��oN�.Ez�"M��lFLҾ~�D{F�";K1d �;�.��,��W����0�q���[�U�G�.k6�IY}fUM�Y� שPt$9ÂP��C�uJ]�����#c=!�Q��++��Et�����d!B�nC�K����v`���8+��Y��d��E/���%<��Wixg��0�t�\��ǉ>p'
C��=��o�%�C��^�w�=�p�����a���H��Ɠ�߱8?Q�y$$��d�/�>�~�m��Ԟ���MIN�8�j[�[5]���3A8Fu(�è-�w�M+�Ƚ���oG�?��Q��^��4	��aMǘ���:���X���y�(�x�j^�����3
��69BT�P�uZ�������"0��_]��*OG�����_OZ�*K��q�x}�uq�-�4<.��
�ʖu���}$�""J!�g��d=GZ��m����,?v��B0���S�^��U2�L��&L��#��H��X��C#��Q�>ҍX;ɨ�~<7���3���x�SP����NT�g�#���ؒ��r%��������.��3".@��)�a� ��+C��U�W�x�^�DA��ӗ����#�+ ��1J!W���u�R�<4ќ1����yN��c�m�7N�z߽����B�e:�$ 9�W�瞷Z�
�z�/qж&�|i6�m�ce��Ί]b@�����g@ A��,L�l���Š0u���w��GP�n;y������L��K �!��X�C,���ă�j�֏�'؛=�}�J�4l��av�(�G���$�~T���!O���8�6ꑠ+�FϹ+�g
�f�~{<|�������;��)����\�]�ZdO{��� �1�E�JM�����M�������|Pa�놀L��1}���q���Zo�$�W�Y]K�+9��D��������(]K�a�5���i
���%*�pOT�ۧUﱸ��uM��5�W��|��]����fT|?�bz'�5��Q��̨,�z��#�k�4�q"?�xЍ1�i?��܉45�|�LC:����zl~Ŋ�sF�'��U�<���߷f��\���u�RO�ǩ����rX#��4����b�$���