��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�u㎺��` }
.uJ����4��s[�����+	�E�FL<�j)w�vۭ��$Vf�DK�;D��ۯMI�ͱ�Y���yb�M(��Yv�ՍD����S�}�w��O���iO�e�b�s�-�������	y��@��a2��`���^�Y��$��-��^6ؗ�n����r!��r�������c�����w=� 	=�WB�.|.�S}�@��	ҫ�:��� /�h(T�F��������@�05m�G+;����7S��ș�/Og�Y6��:����N�����K���#��up~�Knt�*��aՍ$h�u k=<�Z_�U`�#:-R+۞��v������3�`3�5��\�������s���}Q^=<cpք���Z����<�D�yt:ɜ�-��/�]��~>�o9k����@6;uxys����l�~�q��Ҋ���(���i��K{k�iz!�-�u�@}q�u�����[�g�+Ee6�ǘH����W-�'B�-�ȈW����2���D(ܻZ���g�q�IE__��T��C�B������HI�*'\3u�wn�u�<��$�DG������"���sӃ����tu�3�����'+��ԧ�k
�<)�A�������x��9�a��{te`m�Ap�����x�\\�R۾���`!�v�hLk��R_km�\bh�Z-����|<QP&"��]�:����}U*h��MMy5ݧ;9k�T�T)&B��[�٭?�s7d�$�*�(�j�_.��)��b[Ǿ�d��_�d��k�m�Cue3�jH��8�h��_m蛳*mSsF��q#��a3�#��Ed����c�*�jb��(��SN��3�����	��0���h�zq�z4�l�,}��k�匝��E6��ͨ���1u�y��5uV��L���z�TW������A�\���L�B:|ʂ^��W��Б�<��N�-_���+���!d�
�~� Kx�t�<;b'�q� ������4�|�u%d
#��]�,���I��Il�\m�3b�Ы�>P��2��R�7L�c]�DFp��ZP
���@�w�Z��+{��G�Od�Wz]�=<�a� �J�xXE�(��l��n��ӻ1e�ݯ|��w�p/��D%�Xb!6�B|�!f6c�
��~�A9aD�"'r�D��G����0*�3�娗S f��'�`���?��y��bB�Re~�;X���w-���J�[�wF����ilњ?o5!ve��y�P)x��2�l}i&K�;	)�۴ue��Ӡ���Ƹ{Ɲ��2���kO�4�Bl(E��q�@Dn�������i�"����Z��m��:>+���M4��>�x�J��,����bgJpz�oQ�^;��=��o?���޽�wThN������So���N�Ә���b,�Z��$l/P�Z�C+k�x����!K<K���.>��)!ަ��6|@ha��yka����!�<@ԕ,��B���9&2��I��`��H���k|���������,���vj����݃q�3�k��G$����v��N���K$f+�dQ+r��R�o[5j�vƵ��'Sh��juEq;:�6�jn/��������jG!~��C��Dӳl�g�%���e�/+�������|7d8f^M'Nȡ]'�q�]��*�X|�W�?�n��B ��&�
��H�v�,��"�i6���%��Lo�K��DS�7�s�[憼f,� P5��c�\v(��բZByAsoШ��� � )�2�닣�	��+��h1��J��z�3�����=5���Y�f�ײh����	m�C�Җ@v[_4���V2�R,%��J&���ܗ\�WxH�<� (�u�C|�0����̾b�JWVv�YƊ\��5�d�@�;{�j9�I1W6��2�J��������7�����IY�L�}��8;�L��jJ?SeޗV��M���DR�� H� {� X�:�@����Q��_ H�j�f井Bc55�)���Na��:k����y��n�g���ץN����T춖?�
�	z *�����wj���q��'�k����}m2��U��	*oQҨ�W!!N�y}�r��Bm*!z#��*�<b����������Q��Xc3m��I��
�RP�^��"!2%"o�Q�B��-F{��=����Jv�1���նW�ºA�Ơ�(ߙ}��:sJ�P�m�O8l
����6v��/�mH��+�G�#S#s�	I���� _�������.,��$Uk�k\�au�j?N\�g#��{-Ƚ�퇿��~Cx�8hi���)�G���#=��x��aCĥ5uf�?Ak�l�:C��8�ѐ9�*M}t�~{�m�� �\^:)<��N֞Mɋ�3p��l�ùu.�j9T�r���f����t�N��%J�),w�xmR���]��� �J��l��Y�i�q;%�-{l�k���5�FZ'2��<Z�p���-N������64�06���q�o^ӥ>���� w����0>C��'uI� ��S��z-�ڱ��p�O��xD�n�%F�Y�ij
�hg� x���L�;j�Ī`�>d�]�"��.˃s�s��<���
��i����i5��B�uF���D���7o�;��@|�r�g�	�t�Lּ�l�z�7'���\L��!@82�|W���n�ШDч�PÁ�$)�?���u]8��k�.x��?��5�v\���G1ӫKK���Xi��,H�)���F8������^�C��{&�?�U�����$�����Ma}���W������6ض˶��!�;$���ٴ��J8��\�XE��(R���e��H��@&4v
%�A{XѹP�P�j��#��j�D5Q �+/���]�ObvZ�=\]p=N.Z]~VB�׿Ɛ5�̈_�D�Wc/P��d)�Vt�7S��1�y����>�[��j*��������rP��I�l��t����9<r:(t��L\�C�c���]����EV�� B��Zq��&x���ԗ�j?_�����\��b!H�~q`�����Ԣ+��E�^
+ܠs��`��j��oH�Q���Vq6���CC�8]���x-	�w�R����FۡP�ffC�<蔅��In�b��8�i��N���a�ӳ��l���޾7�"'�h:vzӮ4���܏X���oQ�IjzT[	�}��jy!���΍�md�=!e�|�|�`�r�v%�����MR"�~����T�|eP�5�l��:n�P��'����6
s	�/����|���i��;���H)��M��:H�5�q�,����;Ё�P��,�@�������e)Q�y�$�Sw�2��-XQɤ7��}�O�����9����L-�0���͞�lz2�w�w�r7��-���E��N�L�#�AY^}�i�מ�!�K=����Zj; g���[m��n�uL�x�Z�ɩ��oF{.<.��-���l�6cm�<�?Њ��O�Q4�L�����q�'Rq��Yw�A�=QMz��s�Tw�}�j~N��U�H< J��}M��s �\gN�>��\R[��Ul,˱��K��@�ou��jNt�u͎�8��uv0�q�z�����o�C�T��(v���O����D�����R `��	�n'M��%mJ�bǜI??��˘gyl6�wo�1�*؉y��kJ��xPK��&��n%n����@m�M\���I����PM5kc�黺ěh��;�Y�~"������i�A!���Z�-��N����&<����Y�T����)o�#%�u밳�i��?y0��:��1 谑�A���7&��<�� �X�����!m{�<��X6\�aS
�p-���>�C�ɞUo��p���nӷ���	xD|M�<�p��م�$�%����%*Y!�	�$�s��h�g}O���S0�<�#��)�{�ŵ� Tͅ-�L��p� p蜏*���zJ�CV�h�z��y8��DX�?�h'�D��J�����]ÿ�D��&`Rpk4'v�/ȭ�DD��l��ߠF�8X��O�Ƕ=m���d1���k���ݘ��y �>@T�}ᴴ�Զ��8�'u��b�f�(��Bَ!�����"hR���a��eٓ�]�r6p0Qh� ��٭�%:k5�Y��Ժ����6[3�Q%����e�[#�O�����a^h�C�V����XN�!�φ�L�ɲh���Z���/�:Ђ���+���oO;o�~ԯ�1��ƟJ��|(��&A1c=�\��<���P_�X�<2�3�"o��D�d� tX�g��`����b��j���1�-pM��\��n��������cd��2� �M��v��^�ۘ��ʦB����S[r�ё����	��1�V�"�%i��q�d]`<���nG�"�(�HK�TB�f�/�'�m�3��F���c��:l����>�{]�`��&-����z����:k��7r��]����񨲩��r�;�q[��L���N�B��	YK�f�~1�O1'JbS��d����4U;jz"��>��1�F�Ǎk����d�-�8 r=��3tL��@���N�~���W�{R��B��[�mw��<���_�0�"�z�a˧x�a��òUMё[�m3ة��h�I',�dj�3wBo���T�au ���`1�[��k�'�C	��B8w{2b�Y��M	E��aQ��4��"/�O�ɪ�ޢ�xN��d �83����;[�v�ڃ���˰�Z_�ɐ�����ϙ����\���Zg#����QIc/��A�2�s�g~D`o�����])�H��t!����=]�*�_B
�nmI���ۈ:q�Mn�?�^��"��eC�>������g��t�M�����*�T�ϡ9�I��f�[�ཌ�F3�׈�!{im	}<�C ����}a��qr\]K������aw�i����y��]��?��s+ʢY�.g5}$O��m]CG�y �m��.�bՌ��~�u��4��I�Eqb�*��v�p���OGg� k<8���ʂ��>�]��$�֗��#%yn~}�9�n�.<��D0��I�$����+�n)㨧  `8_ު�$bɇd��z�v�(J}�v:%��IC��M����J4VL�>/�+��=��hm��p���j�����(̛E��PXwVzn�5Ҭ�l�s�5�4ڀN'fE��~�t�(���j?�7�gb��UT{� �Fwp�v�ho gH4��rݮ����G�q
&�!a�}�K�t?pk�[]ys��Ϟ����c]��N9�_aG7� }��ݯ��ߑ���ۇ\DD�3�����0��*����������n�.���8�uI(P8�>m��ց蜜ԓ�
k��b߻���*�W��-e��ٺy���Uq�R$܁Pb@|�����HkK���/X�f&P�m��T'���`�!;�=��h��VUׇ��UG��a1v}�Cm�Tҝȋ� v�H@GpE���ð�_�AȠ�<�q��L-L����ώqT׬��`M(������*bYl�vJqmӷ��P�}I�!;��Nf��v� *R��Z�W
.�E���w�i�c��6!CHӛ�h�ǫ�c�[��i�Ȃn���T�\�]�cj�X.q��^9��ᬻlI�B���jj��3A?�=l%o R3wٻ���F�9c>��'���X�M*�h_�e�GzZѶ�˚�@�y�ԁ����_����O7VI'B٧� H�q��nı�1�JԐ��0��,�$c0C�5o�!�삍����g���ER��EH�)�;%�'�U�f�|����uLM�RQ�e��lc�#��#�(�FV�-niV�è��_��F��>X��~d<�qb���;]t*M���sų ׈�>�%L����՜|��|&�]Tf��W��M��eE��w�V�?�*�EOP)ҏ\AG?�
\45ʗf���|w�G{�>�+:������d�(�>�a��+�F�;��\�{+��Ѵ��g'}�TH�тa����|���fB���z�9��K�j8�4t��@���S������X�;��:j�:32���?������>ʃ�8�`�ЗӽE���-N!��7��^�:��<���le�ǫ��e�P�Z�'�����L�C��U:0�p��ţ*�KE Fz��8Q�:t�m(���F��J�[������8�y]�K���r�����^��/��-©xa�e��P�G����Kt��,Y.2Cب�sr�ƴ|�\����i�O5��R�N�2��{�>���S¥Jތ3cWy/QP�8�r�uH��n��:�V�%
AeZh�i^м��Kʝ9�8E6�prEH1eV����[�չ�w�`2<.�Aj:^��5��7FQ���u�Z]�U[����y�u�T0a]P��@aSt���i��p�z!,��<d��\�.���;�6`,3X�X�Gj�*v��߇L�'��x	�	����o�"��JȔ&f/<�����)�����d��v�0���1>�Z2c���1m�M�9����R!����f�M�n�����뙞4f�S�Xt�i�*�b;��w�U��p����+5nd�=�\dG�D����}L�"���5��I��S��Ќ5Ӧ��|�g��+"�`<�#\H�1vS��dm q�y+���)`"�����5 �����)�f����mo��d��i�	�L6��wˢev\3�����.��$7>��N�n�	P�
�ڨ�1)�^E��y-[0V\��Uk�h{����P.1�T�-�2Ot{�&�i���N�:H;�<����1 @3C��f���\�F����]/�U���� �Ș^�(8/��}�o`�R$�~e>�[�:O�Yb�*���)�ZP�m�
���eXC?XڽM��t�BvJTF����Fp��z77~�89�FJk��������\ۍz혗!
9�9iz?ko~�I�jG�K�g�ڏ[��qBS��Pk�`�K<̅P[��-5������R�#W754l�]��2_�$�թ��5�cL9�q��P_R�/Va�pp����Ǔ�H��[@��0{��>�����,���kno�V�D��\u�]K6)`K%��{�MY��ר�x�iO��V��M�Z�7�$r�_/�-�n�Tiu�

{���2~n^�|o��!P�Ũ���(�M�D�^�b����@Di@� ���H�+���$��ڐ�c~>�HF7���b�mU֟���n< P)�e¾K�4�֎�|��"�R.JJ��>�u~�UG7�3	������g�*��S�f5���
#w"�u��a)�:�wX�ЙbHX9��v�,���t��s�]�l��M��7�c�қ�.�_�؀j�3~�,`^Ԩ&��Vyv����Ȱ*�-�5N��7}�b c��#����th�(\4�I���*a���Ֆ��Α���y])���Xa@^��@b#���BZ�����ɉ�����D�
��J�q	� ?򝳘b1CS��)-�m��A}8 ���.woR&
�b��?�Nk�._�ZC�	���5�:�n������d"��y�u�&����ET�.=�3�q{��ְPbE��W
���#}����LCY51s*r�'o���_����Z�y�t����gn��W���-׶����e�Sd1��U��n����+��dLf˺�.�l��vw����QD`v�}�� YE�����xM�k��K�eP�|FtV�a4��Zn����v�O]cu�!���Y��9��"k����jS  ��9�6��py�bԀ��W�fэ뇀*\��	��0n��{�M&��\LW��&1\�7�t(��r[��C�6���Q3:�[�Y�Nn�/|��D��D[�l��#��k����{Ԉ^�����D�.L����?�6�i�!r�ڀF�kG�}��.���f
Z�<���!գ��(����Y��8��`fB ��U�`@U�.�R�kA�V��S�Od���`�޹w]��3�
LL�y��S,�)r�!�.�����K!z�p�/�7{�@�ɢWa��'R2�@�d�h*V5U~�AJ���~SQ���ۇpt�v�A=���8�H��U�#e�&#�<��� P�}Su %ϖ@�����,,�WrV�Fq`Yoh�.�&T�O��y�:.�k���xF^
��D���ê���/���4��7M ����y�O$��@%h��lq6��!v.~����V�R�0�]�O�~��.�"���t3��<��A��)�!�(t���ı��̛�q��)�.ڞ��l�M|:�8�+bs�'������
T8��jh��&�9:s^���_^�n��f���f���m��>�n�֒��q�Y�F�E�;�6�˶�~�nH�Sp�=3Z9I���ZT8�n�"|�A�ڀ��ߎb� 46�=��]�Sȏ�bk�����BKhT7�o7�Nx	��y�k�y"����2;w�C��t��!�ܻ'��ثo�ܢ3y�v9�E|ؘ������g�@���������0�s[اN�/)bvH�)�#������D�Nw�0�����3P����U)�N�{O��x��"�z#��&Ax�ے����I�<�_���r���N����6g<c?�}��tX���7F��ڃ@�����X�RU>d0(��:�lK��ߧ���-��k2p5N\*�R�Ɓ��9p���
*�����a�@��Wl-�"�_�RF��?=�T-�7T����"��JB�5Z���T�Kg�@?9 ���0�8��R.�`z@�'��kƋ�ϒ�(B�F����
�HL�6��K� lŹC��b��;���z	�R������A�ȊsA��ʩ�$�,��*��@�E��53��إ�P)��"U��t6dH	�FbHr������QL�;T	>g4���	ZS]9=Q�߭f�o�c��I�����wE�В��ü��/u <"���`���X5٧�Cp@�xicv�;��=�)��|vG����FV\�w���(���!���L/��S���������qSR~�}+��L�u/����|7��Q�+R�_V_��1U� |y3�7��r[ą��E� ����5s�3Q4�Y��VI*�}��k�<�BУ�7ex�O��(�i�WJ�Aփs��*�=�xD呴)x���ꉄ�=5M	(P�\� �K}��!�'�����ګͮ�rt 	�����۫�����i�hr�&�ێ	
��?�zd�%t�n�۩sZ�ý�D3~ڸ�Z7��嚵�e6��P)ı=�V�� ���t�{�爫QF�q4�B:�2�h����%Tm���$�p'P��u�z5��	 ����Zw���b�T���c��QZ��
9@�Ю�B=u(�<6�M��7l��M��N�"��]�_�©l�\Hz���F�!"������\�<�$.�O�V�q�(̏|��ik���	���e���V9(�N�g�gG���;EE����G]o���U��f��)�:��ǳ%3W4�DC8(wkj��c:C;^Uԥ=]	�����؝d�̗L��>�{����Bz��GU�G�8a{���V��K:q��k�{�F&b��z[Pˉ&Kv����g9���ފ�~=�2ّ 9C��J�����q=�H����C�Q����.�.j�ۧ�)ԅ��V�M,6�����"��A���Ɣ����U�8�%[F�������e�"{� α���`>�Qt�y]��8� �q��J�.�G�q�����6�3A�x��pȹ�Ι��f���gKe)�UHk�R$i[��Y�����d��0�ݺ�#�|[����j����cmg�mG�����ĞŘ.��yGǷq���'37*��=Y� Q��k��M(5���οS>f4�)�_G�H�Jc�ET�	\L28c]�u�*ịv<��|��H.(�FO7����<G,5*ޝ���tv�+�~QƲ��6�P�������1�t�5MH"c�&�2>N�/D�ɮ�5w%��ڬ�ǠlLpخ�	��!��� a7>��3���S��N`����1R����Ȳ��b#uR��)�~��Ք�%���������HG��K%���սY�}Vև���'��"��e�� F�y��1�v��=����������R5��ݭ�{����$��u���"?�"��@<IsZ����k��KpJ���$ق��]�l�����H�
M�ٍ��V�߅j�����\�)��z���Xd���+F/܍��lO���x�%�g^Յi��K�C.<�<�ǒ��^��U'��|��Lr��p�!���0�ӈܜk�P�6c��0s����{�ҪǛ!�\�]+��z�����-v[8q�ǈ$�(�-V>�(���$.�Ϻ����uTb�@W�0��)�:�cP������nҙ�s�M)��TW��U�K�L�9V��Ar(��+�p�i����P���	��=dh��˷��c؆��2U��q~.K�ХQ�#��:�����b}z��#�AG^7���	�]�:��Fݹ�^�K��ie��ȋM��H���RLI��'�7��$r���w�2�6��������t�2��T[�؟���]�[$��2l��c�y�a6*�����X�� ע;��C�w��=#�2��U��	���=G����h�w�vrj��*���K����� 3>�nL�M��N(��4{��w���Nc��Z�5W���D4�X>9�Ub^�J�[�ל���ݥ�Z
�$��t��w�"�-��n�$1"����/	�%b?�����	Yc��z�S�����d��Y8��F�Y��"�0�_�O<�#�����S�]_zb�(���ed�\s c.�f�4S���24��M*MxtUx)G���୍*1�Kq-��05��8��f�V1�?x��C� pT����<���}p�᰸c��\�
=�ԇ�����1�`�J��h��	��'�J�>�S>���xk��@��v�.�����ר��$����#����z�V��U<�7HF���ح�	�>,�?�]�m�>d����V��x%��c�l2g�r�^f�mw�h袄>�F�3nϷ�U%����u�`�3,��<�Y����4w�����fn+�Q@x��l��/���Nu+	&���W�**q�g�])t�k&�jk��'��ľJg���!���i�?�o����*10�8F�2��
6���#�M�ճ�%�LEH�v=^o]�̩�-��Q]���"p֤e=��� C��F���!�/*�L���fT&cK2԰]��@{(q���T(��Q���.�{�/�]�W�(&��{�WTq���N�7-�:�Μ,rB��d��7NW.����TE�`��J1M��@0}8�d�p/p�_���6��^I�{6倦�a��}�h>����x!��ݫ�Ǉ�,�uRG����r��.W�i_�t@\X `�R��LS�I�*?��@���__�V{ET�J<�	zd�GUW��(qвhB@��$BJsx
?�l7(����Ԕ"����nF�����"(�5�m-�a��8yr��ӻi��ߵ�V1˸�-A	��X���`�rú��A\�	҆{��>0���W���.-�o.	MN�X��=��-@��a��� �Ŏ�E��%�5Z���|mu~����H/�����wsuO!�9c&�:�#`6a�x,�b�O!��Nс6�i�Z�l]���s+�fw�M|h�^ԙ�8C�Q1k$D�r���vke �n�԰G���"��d�@Ta�>���b0�x�J~��Ŭ�7ڣ�nc��^9�"��eI�S6'����]`\(%�X����;Q�*����.�;g�?�'D�D��\<�O#��2td#�+��]=7fd��U(R��:��7N�V��pT"t|�����/��#��޼�������ͽ u�W�i�+T�H�=C�Ջ���x���k�r��.�Q�<�uu���3��(���������:�J�i���)�DvM;3Z
������ �d=xq3YKP�SZ(�ʛ�i�r{�x��"]���찥�?�/�96�x��"��l5bX]�@)��jW���g��3��S�1���K��k��X�̢����K�w����"�p�:�bc�[��=*��V�q���*���1��'~�L>CH7�We��FA�b0���e+=�ɂے������Y3���r��4� a"+<�;&_���).��Չ�\zs�o(p1:�@�R��;(�x��e�u�J��Iw�O-�5����ͱ�f?��o�co�F�q/VC�ӫ�ܪ����r����q���-������L�@6�����alW�+�QԽ������+_�%�C�v��y�@ 1���be��4U{J]��ԃ�^�u����kꀶ�4���e{�fq|�u��=��;��L��Ri�O<�j�y�>��b&xj�{\ �^(n�|t�|��géP.���:&�<.��E�;y�����g_K�'w����;���
&�3�h�_�^��B`"�h��3����PK���lYK��-L�鰜�i���C�^]��֖�K4L.��*����m�ap�XX=�ϔ�I-��6ws-8*剿z�U͇ckhd*�Z!�T���<!�"�Y|�e�@G<�x�����P��c �O���NLa=��EĘ��~���
k�	^�C�L�y>Â��!f�Wގ��;3N���.ע�稐�&�ê�~����P&�k�<Rp��Y�Jx�!zƇ� �y�1���hq�n�\�����<��Z+�A�