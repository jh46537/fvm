��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}���E�G
.��j�y�G�>_��#�!�@x�6Z5\�"��t^��lٴ[�G����Y; $��юpE��
����]�Rm�v��l�(E�}	ނ�Eۍ������-�WMI�@6��a�^>�=�A�l�}�o�-����q�V(�N�m��.`+������LlX%�vZm�^[ e6������qj�vv!NC7�s�J!���{~n����1W�҉�x��jPK�`�Qё<�(*YȤ�PT_�vWG�'����ߘeR��mv�(��&&��l��|,��;U���F�6��GHm��9!?[����*�T􇸫['�����e-I��u-[a{�
8�l���������`�?%�=��Z� ���~�SJ��o̓�Ù�	��5�)����ȅ�y���N�k�!�Q?$����� ����:=�
]!��-��u� T	�p�zt���R H���>���ſ[�N�z�H2��[,�	,(8�VH���w��"Y��o�櫏]��=j����n�b3LXQb�݈�]��'-Rt0�̴�>�L-�-85u|�5p��e�/��T�A9������&b��̴*aeK���^��H�j��p��W���_}��9��)�/09y_�����YI�Q&-�v��z�#��d-vZ|`E2-�vSE0+i�К�߷��U����8ˢ�9��g���5o�{e�����+?��7{i�g�I#� �� ���.�ߐ1� �����sZO�Y�u9�Ɗd�)]Pǃ2�XT�(s�0��%NC�J�'`S���Y�u� �������g�mf/�,��[ʌ��z��F���B������,�Jf�Mq��p6"�dn�Cu��S��|���B��Fr�u�^��	6�R�d>�'���,g,�u�U�=t��[�~��*ۙ�n�x3+��Z�h� ��4�5���)E|h��.8����!����!��=�Ax	� Е�mSڃO�\V:� ��Fe`�W�������K��EDT�Fc�����mP��4�P����z��(R�c�p���-}���A��7��	�M�^�6�\-K�e�u��u����V�mTh&��Ll�2�(LO�O a���\XW�O�7�����
�Ȝ���g�aX�鲙��f���'��IƷK|C����%*'դ�r�d�q�	�6ֈg ��ˋ�T���C�(�r��#Q�����\ v�'-�9Z��K���fV�Xa�O)V)+�"�)���q���t���s���%�x�#4.�SPd� ��c����Cp�|p\���D���/g�
���<�i\�)����2,�__�:�>��>_��~��O-ށ��e�|շ_��Y2Cɀ�GU�Y�}r�Y(����5$��oZ(�K�o���H���Mo�m�s��3���+��{�ڥ�����qi����I�-J����jڣ�ѭsp�m=@vn%����e��?��a�	D.��Y�'��8aޙ�*�j*=o`-��}}��$;B�x+:؟(�3�"��/�Yz�4�7���'�'L�U�D�3Xa�F����*��L�������Ne�Y��?k� S�H�	�(Cf�kc��\�by���oB��G:��mT2����^4KTH�;��A����C�}�('������,]ױg�\K�����2��XQ�^�'g4k��8NZ(z_ќ���cy���I�q��b����;�y +�xۣ�����Has�rϩlQ�T�EB�CPC�����˩�ד)q�},��̻�Sz_����V^�0�+A��7+�Ƌ4-��n;qc}U7��W15�GNrH�<�ƥIΊ1��/�h0eF~*�/#k�<��a�Rʑ�-�`�G�x��T��(7=/�2���$�HzϘpt�(cʤ�㧃�x�a���K�<�[Zo<Y��Z&�BZJ�� �_�@:��5������a��B���R��c\LH�K{�(~Asj���a!_�8�%���%�iU��Q�$IRl�(�M|�xAƔ����nݤ�I�m�u)Kv��n�q���Hs�����WT'ṂC���|k��i��J_+�b2�e(���B���T�ѵ����e��q�����zk�~�*X
�+�9���04�-�	�]�x�s�~ �̃���᯹l��d���a8�¶�?��̧��#��ÊyY���"'��'9����	�/y����X��M4̌3�`cz�����/-9���:1�I*���V��F��K���4|���錐���{�G�*�@���Ϊ�96� E�8�8j��ᚻ�:�`A����ݤ�m��@}.��aũ�;j���O� #��3B�i'�kò��
�`@y,9��u��x`��$)�u�ш��mg��E:�����I�CʞH��T��zM�kѦ����	���ң�J�;��
�2�ٜ�o��IؗLyn�x�����V�<q }�5 �f�99�o�6>8O���0�7} �k˃�4ؗ}���FB��=�3֌PI[�J���YK��q��Qg�-�Nﷲ ?�s��	ޜ�N��#���]`�T�W����Z��M��t�M����E �)O���1Z��KRR»̎8�w����n̆O�����a����|#KEg��M�.�E��jF�i�"�� }��9c .�7�iMD>+[`.�[	�
x^��kɀ�ڡ3sl�)RH�#A������R1 ~`�}�QI���8Hҳ�jI��ROM4u�%T`g[��r��#�n?K1�6�I�mg������=�w�'k�^ o�Cɫ�j�UMn�w��\S�ۜ�n�� �k�~�׭�ybؼ�t��@h�'a \���\��t�LN�nV�1��OS�*K��)FK���*]:$��JFΪ��;z$i��&u��V�V�����J�����Z�̃��$+ՅUH)���W�
��F82���VV��䲿�)�kX���ao9��v�hMG ��-�xG3�́�Z��)Q�`�˽_	9��͐>����?��?#w[���OnIݝ�9�&�K�I^E�Iُs/����V�Ћ�&�;�cL�a	�Ly����S�qv��!�4�+�u��&�
�:B���l��L������I��0�>n�
���Q4��J��)&�o�c��*��7�N�.Zy�߉G�=�^4x%�f2�0�(w�@Q6��	C���Pq����'��s�z��5�j%�%-���T��w����A��6�&p�D���3mG��k1��䤫PS�����zY�(W������ax�A
ی�>��*�DM�P���yq��짇d�%���_
Ը�����+��1�3@=Bz<&��WQe���`���E& [ �CD+�x�����X}��WU���:j�jv�L�����W�r�e{��e����� L8�T�^�(� T�����?�s�S񪛆��{��`ᓎ���`��������Q�M�x�R|fe�1?���y�=@/|5 G��U�״�.�:^���M�P�����4���:� �"��}L�;�P��n7���c����D�i������X���[��0K]G.l�-����0@{�:�E�DETl���s�S67��7ixB�z@1�p��MH��~T}�
�Vw�����xc�����y+
�Y�(����`��d� ���s�8�M�S㻯�}[ͼz�a�G`�W�@�)������F	}cf�DU�'��@��͉�`Qa��s��8I^�L�$3~������c�b?k����'�k ��`42'�2t�d���(��v���s24O�9�u{���Ε�wl=�41c�{6�k�g��vG�^v������ne=�@�d����N�75Z<�ٞ�aQK��j�?�W7v���b\�q�*)Uj*���R:]���HɎ"Y�/����R���k���LHҖ��#i�*����/��}35r�LY��R�B�<y�P����0ǾzH��^��$z�;8%�&��p�#g�r�忴�>�gWrt�"f&#ƞ��NA�'@�?P���aՁ�вxBTZ���T�fv$w �a���#y�>����ev�߅���F�h��H�&�q��݀���T��
���ֺ��$�"�]�Q>Xh�FN�B@ˋ�XLh��o��3���{F�4N�k�eN�Gd�çûmhD7�t߶����N��j��f�Y���Ƚ3tZ0�[�-�iz�/�p���ܺS��i>d�G #�k��%.������z��|�tK�n����I�Ϭ������ԗ�����,�VB݌׵��+�˵[���Ԃ�?ފo"ݣ����������
�X�d�?��"k!�#)�`�˴M@N��A3���̒Q�&��1	B��c�N\ÌߪҴ��}��Sg���7/n�"M2�j
��X8�6(�iW�Go��ܥ=*q�8������k�kYԻ)�v!�Ì<��,�oy�X!��>h�YW���CFl�E,�����@�s/���<b��\���3�f�̭SdFP�t7�Wl.d|Y�e����_��ȡ�1@Ʉ����"�U$Ψp�� ��_+�Jr
0��@�z/�^9p�_�5��Q��(G$&����gtdÔXY��\��P��j,��Z���6k�]$:�,�ؓvY�A��P�I7&+��L����.όvT~t�L��֨?����,���ձ?�Z�W7b��q��%^�$ƈ��V�����-l������5�腰�&(a2v���x�~"��?��ű�L�pr2�[��E��a#�J.������U�U.�cF�R���J��9����r�H��T�y��,/l9�����$`����K�`H�oin��-���[Jk����6����I����Y4v��"f��
6.9�ƣ���榫#Ԋ�b`��O	/��X7q�m�h���?#�=n�n�e�� p7&Vmf��̄��v����(���'T�,]1R��9~ ���y�ZTq,�_��´�O��{�X6�d�d����o ��N?.�O�����
JBI��ѧ�r���#OHi^�����N,J�#a�Id���E�(l��F��+S��G'��P��zj/[���1ޭr&h�f��AE.��ߢ���J�A~�^Pt ,�v2MuȾ60�TK���K�+SQ�@RD��ǁ�%���B��H�<��[�Q���j���Q΁A�ۜ��6��ܛ���ㄤ=�|e:�Wh�S!E�����e�A��[Q��oAV��?@�[�/4}�����M����������i�KUSs����](t�1�(7���ū->�-7t�-Jq&�]�E'�7�P���LK)/���Ɵ�YG{���j�Dw�~Y�z�D�Gyl?�]c;�c|�
#��P��˩�UE�Qɫ��I�w�c~rK�2�}���5 ���D� �)09�r]��5!ݷIǆ�i��<�Q�G�d.�xh3	Zo��Q��OwQ$BVK�aֻ\��.����` f��̏;��K�v���vL�ykYF>G�%>�Fv5�F����̲Wq�����	 `/Q�~_Wla�i暀U�%�Q܈�nA��Ĉ�����sHЁ���0e^�ۉ2���#3Y�*w$�-X�o�`��ѻ	�
Y����C*>Y��oB��_/���n��	쁍��@{Ts偣���R���3��`_lKC�5���RA��I���deD2}�sQz��?LZ5a�KG`||=3����eW�����G���q�Cv�0������joQ����t_����O�&:/Zx2˻_��۲K�Z������ ���8 p��_��?fAٲ(����6�?���t$)uo2 ��4��)#B	�^��ĭ�j�%��a�4�*���Ԓ0��O�*���9��*G�����^	Z�'��n�1�;yzK��j���cۧ2c�M�?!�w,ի	 ˶MwF>�ڑG�ٕ���2�?nx�:d}d���x�̑m����+��ЬF�Z�;m��\4 �y��z��vP��j(�&�v5ZGy��1猁U�Չ�bd�X:��hl��ځ�m���h��8�둡5U�W6
�&�It��C�7���J@U9��#o</����7���Fa�fç�1J�E*@�S�P��<h���2�;���S������`�쁷����\+q/D|��e���Xm���O0"c��ƅ��d�<�ͽ��nX7j*����[]Duj�m���w9��5�$㷆w�n%n |�z@��].8&�ד���Z���GM~�D�I_�_(��`(9�K��y���;	]��
��\*�dK�ڮ�)�i��/���v$�`&�^�
%�Q���*S"�Ӧƪ��l�p.Ю�+'p�I{:f���!�E�ng
�Ӗt�e�.R�]����; �CK����|3�E7!9�'8(��~�axt@U�n�ȴpW��d"����~8�\���h�������݆�I�4	s�;����=�L�@HŚPH#�a9��˽,�:�,��o��<���'�5�V�@�]}��=����2F�h���6J,�������0Q[ p��Rr8�Bu�.�x���E�t1���TSo�Vy��,@��rS�_�!l��16Lm@ς��"r�Q�f�:��@,�γ� �R�/�j����{��<�~�����R��x��͢��v���`h��¥o��U��c�<�H��!��G�]��q15�r%�NNP�I�]?J�d<�����u�P�@-�/xn^���˙@�R��1c2��s������/pa�a�FŮŸ��U{>H�f��e��b���OT	����˥�R�C���;%�����g)-t���"��ͷ�����Dwx1�Ie`3vN�4����/�o�纞�T�du��i�9~��韨 w���;\<�9\B'����"r\�; d/�����e��"ǜ����C�g��S8�n)�l�R�����tMP�3�7���|�C=s9��$��Ä�����P4P���ªe�x*O�Ah�_L����/4q'��0 �|xCZ|;�?�<
rhoY�g��sQQ,�|#�H�������p���,�I���ªn$�PSx�f��Rxņ�_6���9�;�Y����.�E?#��	Yo���/�e���W���U�2#2�u��9��-.m��g�)���O�w'n��4j,�Q��1��t�E�w�0\�����S�96��iŠPF
��t*M�� z.��T)�=�0q��8n_��l��X;֟�Ϟ�KR[�D���r
0E�^�Kj��o¶~�'�\��2S���p ���(���Z���S�h�]���efA7�I��|�K�&R]�BN�)Y)J"��gH��X��.0��	�u]}�K:��!ϊ�2W�O����O�	^0x*.��NQ�6)L2�c=1���l_���0��/�Oz��+y�X3�C�@�4�gq��d�X]���I)~������ٍ�Բ"ׄ"��l��8�]�-��W㰇@DFy�s�Yp�3O^���������"R檐d*�:��*�{޶�+���@n���p{5��K�k�=A�š|{}rѯLaF3�~N���xf�p�%	�p��o�a8D�߽����U�Obғ�/jE1W�M�\϶s�q�Vs�=4�]�h/�G�n��gx[��U��1�`��0�P�ɌÑž]ԻZі��b�pg�$�&��l+�"6Ҙ��)���,�1��\���YS"�D:3�̃wU'a��	�W�m�`rj�L˻����߯�+�e���7�w���?wvb�]찌��xV���� E�)� �|.o�KaQ�6Z�p*�`>�9|p^��>d�	ݩb��E���SMZU���1P�X1H�8&��L�/(i�|�$���B��q+��y�A i[^s5 �"۰��e��,��\t���:b!�Ņ�r) .PEL�Ә1$T�!V�|':��G{K��77>t��������H��7�'D�rc�>���>�i� �	._�"m��r���ˍв���9 ��C�/�A�a� ka5N)>�A�i����-)���_@`�o���![��)�oǍȍ�:n��/��p�ݩZ�Q�P��[$��$þ��3�<"�Y�i{v&U�������H3 �1Ɔ���2�ۋ����v�zX.��Z 2�h��pȣΛhG��h$*�p��o[=7��H(���I��v��k�
����L)H�y��<*=�-]��U�Q"�!������!�?��-J�a�k]�4j����U�
����i��~���g�}Ȼ��_��]2a,z6���RU���vD;���l���T�ណ�^��?8�?i��ο�ko��¤�k�7MW1��oS�[�]Į�4��<������ӥ�4��~����tH�6���z��6P�&�2q��L�T�a"G��K��T�n�S�rmO�=��Hu9����-v �U��g�������#�zp���5;�AC�(=B�{ғ�W���7��E6ߓ(��}Y����^I1��Ra��-�w
u�!�D�zV:`#�w�U�i�-@q<P[�~uWy[^����`~-^�M�#���O==��w�vԀ����ڳ|��� ��wk��F��j�}G���AG��.?�97Q&51S�K"8{��.8���|J>��:ƬM���M=��"7�A����؋w�����_C�-��RS鞂��n�)]g-.�#���-v���V"� >d�U�V ��U�i$ն*���o)�Q`�&�׮6 ?cX0������1r�4%����15~����~�%������Pf���Xki�`�BFg�5�586�lr._=W���t�ϣ���$���s�$r\�P�!�B�q�8|�>&T���P��hǐ�D|�Ò�h�����.����u��,b�;���p�! #l�?9H��]���G7:��T(E=�I?��.0�!'O\����BY�/�yC�VX�]$7X�}ӈXPlL5h����I̒���v�N��?֞�@7W+���0 ���!e�S��V��ckfZL�h`��_�J���*��Gs�}ۙ�D�'�r���is����Ol8bO\>p��[�l�h\��+�����Q��smW���~тh$B/H�JG*��Cl�b����eo���P�K�g_��(�bR7,ST�N5)Y"�,\@�N����B�д2̋�@s��q���1�uQm�.ߨ�BX�oL_F�Eg���z#l���DNă�F8��3'{i������Ԃi1�UI�`֑�L�#%��g�{�A�(d���$�����hO�C�=_��nRS���a�[��Nri���Zz��篙P���L��x"M.-�'�q��'�,M)JfZ�rXdBQ���_���wg@�E���0��+�Ʒ��2��. -T��,��}+�ؖ��9dy��1�K0����E�%w���N��B����L!���|؎B�	�E{C����Ca $�}�V/�r,�d��C^�f�%fsDg�����{���AkW�E��*���/&X��ӌc��@��«��{�=�9dU0�C^�f(,�I��h-�kщ�b&�J�B�~\P7XSl
�7���If]�Qx�G�{�0�b���鮌��6C�V���S�����!(Q��:V<,��]�R���s��K�{7(�
���6���Fk��4���h��q�@�r�I�k���z��7;����w���Ba�7�`X���s�[R����k���T�x$�i�����/7
xH^�n�����Xb���Ȱw�ܑ�4���93��ӌ�s��TQ�C0̕9â}(4�-T]���㐸���������	us��ɠHF88�F�^�JՐ��+)�T���H���Y�q[#�����X�j�5gƽ螰�Y>-$)���L��J���t��&_�*ֺ,��$ ~��HW:�\a���E����+|;�S1|�E��;�jY�@��=�$D�4���vy٠f�Ֆ�w�[���p�Ғ{�#BI��L-R�w�X����|���H9� ����3��Ix�7���#k�
==��}B%raK�&�?E�<'ji�����&��l�Q�I��e��z�[|S���� k%�9Z��Fb҃9����P벶�������\���0�5c�Ubc���@�
�������m������H�a��g0y���o��G�cM�#r}:���a�^F�߳��Ā@5�-�ktHУ�Q҂V�u9C��R�e����V�/MM�z�͛���.
�^��Į ˵*�{�7�9�+��i�G�d�W	��m��K�Q��RA�T��6Iډ�������mg6�/�3�������JJ�t�àX��c���s0�'L�]�h�I���FAd���ӘOA���s����
G_;Ib��卂��-��u�K��ǿ����[�ߍ�����q W3L����b����d��>�L]��_/���/�v�1���@l	
"C�\�����W�i�i'����o�+6�����ϥ���;��9?n^vw���z	��⑐����ُ���	��J ԭQ0TY޺��J�^���z6��b�/C/�P������z��+��NB_
;m�)����'%���S�ʧ�Z>��l��ar�lq%[��$͌G�MQ� ��g������4�`��r��ih���)_�����@�$��P}N��0�7���z�����Si��q��n�>O��|_8�~����%�01_����{�'6'3�4h�R,��W��1_P��>�U d9<"L����7�s��LO�.h�$N&+���vo����O ����q`,��d��{'@�Ը��Hb��Ƽ�a���=�xn4?��Y�h*�����R�_y�ʠ΃�*ؗ��	�QԊ�\��5ih��X��!�}R�U��.�tE;{�� 䝠����sWq��`�u�Jʫ(b�w��&b،y!@@��FNt��E��l����7�v���4�TIH'��Z�UL�����̸�=Y�$���!��}3���V��vd[y�`�O��Uv�Cf�d�-�+��~{}�w��pW:�L[(��l���q�e�֧���>��&�
��W����p|AC�/^����4t!:g��S��:*����G�=:�4J|qX�$S6�Ѯ�>b�/�$���Gॐik��������/x�e(�`��
 �s��������l:θ�kъX����ȹ�99º���Wь���OJ�f0��2�D�^���|E�eq�sdk��Ƙ<�)Ǆ��=f{_�-v����!u�E[�C�I��1��X��A��%�����o�t�vn�D�>��)�Q�glTP�����Br��%�K�xGb4����To����`�xh���<MNU�V�TDi�T�~�mMsB݊4	)RU���oV�Ѿ^�eF!5���li8�h�C�����S���N�`�]loaY����g���?G%BzWY<�^�m�K��΄����K�m�����-^1)��c���x'���YǨ<����3��V;5g��0�;�ޟ�(�����3���~&��п��Q�\!�%z3�X>���<���5��Ͱ=�fh�9C���_"y�xn.G��1PYe���u�@>�O�0��/�FZ����]qo�{r���So�B�<�#̾�mHrǉܬx��⏌a�,����!����Ka��t�޽����^���{2�V��/�-]��?��9ݮ�;���35 ^bϹ�O'U�*�:U�vSm�tX�6̠�K]@:�'W+S�l����!��/�ړЉ_�����7n��;KEb$��|u��A�Ed��M�d-P�����W�U/~��r���}�1P��j;WG'��ϖ��~4o�8;aFW��Z2:�����8��&.+�(�?R:���
��\MwO[B��C{�%
���u�|ri�g��mc�M�ݾ��7��	�>�#ٹ��e�.�+]j�>�	���cF�S��Uv�o%������1-�������/�g	x�)<cO�5��̃N�ّ��7Vꠃ�Go�("�m�/CY=��P ��&9_�ϙ7���"�y}��zWA9�X�2ʶYKU�V�Q�a����G��f��GV-��q�-?����di�N%��<��g��m�т���]���A0aڇ�����z��Đ�A���4�@8"mO��K���R��h��dU"���:�}��geG}9�R��/gv���wQ �Y�\�Շ[T��P���r�}�H�0z�Ҭx*F�	�l0_��e���`���#���!����C3��lq���hP�_?�0=�u�ý�s�ć��s�9�Y�Ldn	~4��D ������C*H��g�9(e�l�j!<�����Y$e��{��Ǿ��ȱ��V�i(*-�� ա�^Dj9�K�[ƅ��R&��*GA1�P}y	��2��Ո<1�>��z�x�8I�H��0�yN���t�DXv_�n'������н��k�ɂ�`�����",.��j���Ito�b	v�3�/ن��ڸ�49U���B1]za�*]~Zj��2�))r/�5>����/�dm_Q���r�mʗ���@i�+�8&	��z3�ͧ7�2A�D��1o�Vs"��as�P~D��4�TO�D-�F���[��
nS�ȅOMz�i��y/(��X��	H��� Sx�"��R��-_pYʅ��a#��&�nv<bH�_@ p�vbQ"q����j��zk*c���1��"]%�1}U��E ���'���N�:��(C��,s*���M�U#y���~%q j� T[�������E�M1ޚ�=a�����n�Y��S��J���^Gэ��Qm~X%�&�s��Y>�+Z�Kj�@�v��D�4�Q��,�爢6a�?f-z��p�i�G-؛+3��H$��5���fy��k�I@yj%n���X�����`�ٗw�+G�^o���@�����vW���N#+�2��O|܅Z����ө�`�rQ�9g�em=p<J�4�T��Ie�����Pf9����'}p�k5A�`�`Uw��]�rՍ�8���9+�H�Υ �
�O3��Gӱ(n�T��c��d���RĚ����ǅ�=U)�?�j����)d��n��t/�m(�/�뜸+Ӣ�c�x��-tRx��F�["j����d*��R�7���u�V;�Y�m�	p�0ܶ�՝7U{8�F'����wu3|������|�
sZ@AH��vX:)m\\�U���NpUJVQ� $T�G0����'ĺ�z���C�=�����|�2PK�1c �>}�r5@�ˊT�i2O7�mj����X��Y6��R�H�ה�8�$��k�4x���W�n:��#m� 2 ՒrԆԊޔH�uwG��"��(�{Βo_y��5 r����[������*�:.� �o�s��%	�]�G�� &9�����]�x��}�hem��y���0�z!*p.�dbK�)�'00�J��5щ�% �8+>\]
��mK��z\z�P�f�Br���Tŏ�61n��4;�L[�J��ܜ���g!M��E�A�L�� �-Q���S����^qOj���6�)���'�)@˵���kH	�)}�}�">�d���G��fO+�-=���I�@���"�v�iF�vێ�����;�+}ڐ��\�.�����=�b�C�k��9�k��QƉ-�a-Z��>��(���Ҩ}#"ٿ�
>P`Ҥ��6��S���LgoQ�>�Cl����Ks�����W��DŊ�2!Kщ��� �fK�M���4u8o+b����4�Xk��0������n������dX%Z1yu�y}�6:
�)�❔�o�,F6B����7D�\�ɪ� ݃Jq9P]�۔���`���m����a�/r�_C��OБ�qQ���B٩6�wD+a�Xg� �T��BY� b8��A$(���T�W�.f��<+�k�Tw �Sύ��YB��oBzLa]�w�]b4�-tI�͖}Kq��ץ5��7��\W��&����(J<�h�ȻW�ҳ6u�g�C<`F�@HL���k�*E+�R�I;9��v�{LM'ZF[��Z�����:�%k�:���?��R�ja��P�k���$�*A��$������u�q�K���'Fbj���!�J���� ���u}��Jw_f��JG��Z�[o���^F�b^��Z��Q�{��p��D,�6���⨭�ݥV�F�j��	_���="x�}����t�\y��y=/v�Vl$K��yUTcO��Y��J������;
�t@�Y�)�
�R�z�G��)��� f�!��>*�.8���	tX��O!'|��7�gL{g��q	�w�jt������m|4���� ����Vn�գ(�#�����un�9��}����1�M�#s R�����T=�!�j'Gp���P�f_��iP�hx�����yo�	�\Q54%���f��/$�)�{ID� �8�򠁽�b�����Z�	+�r�\��1�	#�o�Y�
ߠf�Ɋ�/�j8�.7���W��v�	��ҳz�J�J\>�*�2��)�f�\�-#/�B�H%�Β}_�V�CT�̽'�M~�} s	����%���F!;�~e�s�+GלF��b�"�n�`(�s��!�Ï(ᚨ,#Z�go1ü~�D�\^|�9�k�ʥ{��R�}[^�.�r��0�6< �C�4 M���ٰЪ�� ��U��:	i{K�ߪ cm�yb;h��4�V����!�R�X�QN�CM7+��9�N�X8�(��޸a,R��UPj����_謑H�`8G+��$P�$I����+�˩�3�h�p��F%2a��N=J��8��B/F�:#'�{�P~���u]�Iz�,�Ѭ�+��F��6-�?���2X�D��1�E���  H�9�Mz��gsQ�8�G��K�p��w��dMX�gӭ�k���x$D�3j$��k�g�AX�;j��I�5�V�"I �lB~
.|v�r%L@���m:7��aA+�Td� 5����^�֢��	�� ,:ve�%�I�'��I��^�q�Nu=����N��c���������������)b��G}��9B�x�x��y���n~����m|9	Խ��Y-�����:�D�gV�������Y��F?������$�Ƀ����	�BY�Iz-��<0����NH��*UP�%C�)��G�-�Px/�X�çn������!���	m��#7s�!��x7(�_q��}��o�ːǨJ�+ALVLi ^��MV�[�G������L*x�՗S;���k�O�fdr�Ăt�
�T�'��"��D�q��\N�u06X@qEJ��5����GZ��eS����3�x��9�S�|�
�0��T�=t?���zkB����3C'Q�?�	����-d\�g�X�M	(�ϊ�E<�`:�:y�f"��,_�ʯ?:��u%������[tEp�ī���]'Qm���h'�����t.A����w��o��a����2r�w�p~��.Lİ���3����=�5>�N#������j��#�	V�]9l���V1ҿ�?3m��Ԩ�m���P^�;CC�4^{wS^�d�kߪ@�k�3�e2}���)Uj�T\���������+d5$��a�p^�
wG �	��`Y{���`W��
/0�@��1#JK��:k��|9Zm�������5�w*���� we����J~�u��^?A�k(}g�Cg�%�7�J��4Idv"f)��9�	Ge4��U��W[�&@����������`����'�:�d���/��ᒨ+ �~N��f���HʪKM�z�bLw����o/h��U�D����G����wp:����vkR�[����\ ��މ��3<����c��z����ǀq6z�P���E|v��F�z�#������K]�'�^7v6y#�p�=�?x?�b?��k����2F���tV�k��9*
y@���xߕ���fL��*���pk���Y"#�Ă6L}uQ��X�Q_�%��q>�v�~�(��qZx�ϵ|�H4Wo�21�2R9�n�����D�:�<-7���CR)��'/l: �NK
Rk�0��r4#��yY?�Ŷ@>�!����y��byC�>8�M��Bo%��Vڧ���i5qK���4�y�v"dc\b�������9 ��' �m�BQ��n�.�6{�1ԗ�5�~��t�-L;?Oh�+6H���Ą�A�ve���0�C������_m��uһ�dE*闁TՃ��m$si��]5O���}:mF�$u1ĭ��KnW��>����ӆ9�F̔�{����xlq�`�H�Mt��Xj�d�W�F�`�n؂(e2��+�rUZz�<��"`.�V��qF��ĸ(a���3��r�,<"V�3$l��(B��`I��l�a.�=��}E��{�l���n��/d9�_C��ޛp�)��ߧ�bb6x����r������N��n:�C�F�� ���Zo����XF���O�-ȋR.?>缎��E�i��M�ƭ���X-	*���7���wzY���A�i����?�.?���7)g�b0ai	X�L��%�,m�TJ���険���O�JW������+Wn)o]ħ�5e�N<7����8R�nM�߲D�9���B'G$NXT��3���[Z�?�zs�YR/@Y�'��:� U�a��[�ҩO��q�a�8U(��r)g�e���Ql �M��������p���ʃ�,�z�.���QAi������rF�
�=Pby�D�����ƹD�)���a�;�!fZ���(�\��h���2���_vF�vq�  �rm�Y[CuȆ�&��T{�tὂ �4��}6m���3�є��R�g�R&a3(9n`�m�8��ѢQu�QB��\b`Д���T�[+)@QL
v�a��#W�@C����3���č��M�h& G49�R�m?����Ǌ�Ek���3�-i>U����Ns�ZK=f]D'5D߿<taFQ0f<�,{�'�,w���q�q҃�O����۶LܡwY%��7h�,m׬4���UY�ovj��w���*-�|��EaG��H�#$��zm�;�VC{���n��S<�pdM������.sd���i��xrV�	"���xs�ѵ�ֹT��,Z<��P���3�+q���:��*�x��RV�R�� >c6 �Y�����0�^���qC݈��
�Q��8�!�0l�q�G!:�}�˾m���f��m�Bg��m�d�����9m��+@�I�}<�t��S���T��7:_��LZK3��`�	�p��%��v�@�UR=�ۏ��}7�N���/sH$F�9#V���4Y���N+���0�&��*d!�`�jH'��+�e�UE5��Խl�h1F{j�Vuj���1E��]�$YKC�y��U�@2|݁�|�Z`��ο��%E��py�"gi[�'#sN?o�����lp"���<w0qb�" , DY�Ǻ�hf���'��xP̏G5U�ø��iNa?Ϡt�p7��"�6L;~JX�:�x2� �>栱lQ\�8�nP���A0�F���ϑ���l�ɛ×���>n6 �@�}�X!V��0��=�i����llx������D`�4��K�I??�<���V�S?I��Ѫp�ͷ7ƚ��Z��&Z��j%c��Ku"Va�	�n�qA|M��37aT�������R4?�47�ѽ��o��3�.�I1:�e����/����3�����^��㲂�v�&�x��y�b�{�弳˜A�V�����ј��Z*��v��r��0Ľ�Ny���3�5R��׵��ئ*,M�j���5e�TDc�.�0�XMQ��ۉ�`�6#d9@�7�[�A��I7R�<���Ծ�����T.�?�]o�W��jf�*���0���R�:�;����3�ar+��ɕ2��X�q��_y#���g3W@�|�A6LwH�7)ƀ{�~$*U��!����Ф��	�T�	������G�-���Gh��) ���W��4�మŘ��Q����U�#������ M$��!.�nJ���ץ�~_�V�J��Z5:�4(�nD�?���|�m(���~D����К&���{i#��a_|2$������	{8���հ�T.�n�����������|���w	��*33�y{�M|�8p��8���U1 ����D�*�Qhkm����R-���'�	���j��ؘ����X .�݋��`	�I%��T6�2��	�y~Ե����������ۉʡ���������R;%�H�x����j
9,���N~� ����PA{\����M*��0��*9o�g�:����B���)O|�bL�:��+n���%��/\�O��A	'P�j��`�
3��!h���<Z�d۔a\Z穪���ײ{����&�%�3`�/<L��e�����a�c!v�$1v/]�M'�0z�׼;Z���p� �3�� 	ʉ�lrP�c`�� �ݬ��a�uHd�1৆������y|#ꭞki.5�@Q�py V��q�������l.�z�m ��؈�� ǒ��n`��ͳha2�.B��Q�~������sν�s�jBpq�<k�����D��.���k�r+kO�>��v����G5�M��s��.�6���a�6%���_1�r�g�R��>L�,w6ME=Ύ8�h����*6o����Xh�l5OY�}�h����
~�潯�C��s��L`z���?��]�<��*�x�_��q��(ؽ����sXwQ;>��s,��H�$�@�U@���l8t�X9s��W�6�{h��*g̬J8w�-Kn̺X=~���a�vU;a�2�>m�ѷ�A�g��8�XL�@T1��VF��l��k�ʘ��U���t.�B�+��Kl�Y���񟂡�Sŝ5��D13�L3ՠso%(�U�)�����n��
��&ܢ>:�½�T��]T͊b� n:��L�ڃ��N��TF
���������!�V%J[�N3�H��0��e���M(���3�c����x���#���$U�4M!џ,���S��Z�[L"�(���EH%���:J��(���4��;@DCb��x�>�$���T�ۥS����**y���Q.PoED:i
^��FQ��_N�۽p�)�2�;Zc�K|���R�0�a~�>1ʴL0e�L��T
����q*�ʇ�wUT+`�$Ĉ��������c͒s?&��^��NΛ�ţ8b�ܘgyf�/J)�%ï�b9E�"Dk^��H�j&�`�m4~��;�Fk.|o8�XYX��;��ދ��Y�g� �񪞮&Q�F/
䱁3#=���M6����D���hA�� H%��?ص �P�.�C�S��IY�]fb�+o2FI�(ӎ�4�v�G�!�j)KP�)ȹq��h�B`� ʂJXn �����g��Ӭ�ɪϝ��|n�2�5)xp疄�#NVS��� ���x:�m��i�	�n�zҰ�sՕ����Ǳh��^�x����zj	��o���d5�����0,�Wt��_k�zӆL�{p�ą���w)��1��Qn>��JW�\TgK|Q���ǏH&`؟��?a��c�]Fi	�;��C���E�$��84�t)�b(Ҹ�*gv�Q�h&i���&��L������o�.��^�r�;ۊZh�Ͳ�����ׁ���>�(�J��BN��3���6��YL!#��������Μq[��N�V��Ub'���'&�ImEvc����\�^�@�0v�jT AV|f��{��˅O���%y�9i1�o/���S9�c"O�˫XH��sȇ|f �C��KbV�1�a�p �����ȏ�S76�jvn#���[�F�����!х:��d�K�Ri�H�i�]T}�V�IQ5.���5㲯��.3��x�ׄ7��z<0Ѭ5�vy<��?<��ֺ:eV1B��6��~y�T`d�v-р�8h@��oψ#�\ ��F�,A�}�	�Kض-��ݏ�lEeY��^S_\�Y�XK�o����&�U*@�)��e5�9��	��q�%7]�ns�9����A����Vg����0�eJ���fƈ�mem�Lcz
���^�r��=�rAs����s�~���
�Dbvĺ	�q2����I��F%�c08!s��a�2|��K�A�e~	�ƅ�����c������M4%`���#s(�]J�%��u��3�ɕ�\sc��$��޷<��0��]c�i ��L�#���w���pP�1�7���h�B҉s��I�����5E�Q{f|�(e5�gL9�-�F&J�7凶fX�.��R�Q�Kʆ9�%�#
9���j����{��=��O�@Ry4[>iS����9�od=��L�V}�G�dz�Pyh��Bj�"5�ӕ�E�}�;"����&4$��m�
�7�,�X��\�*�y!ƛ�K�mc��\L6��aJ��sԭ=����X��)	a�A�^f`���`c�2{��vX�����m�*9�1�%�&���EI�o���v��]�0�DK��@��T
 ���|	V����.��;zg��ᆌ�0*:�\��:@l�,����J���W�!k�7V8���6�|ox���/���ca��J�[�T&�Tt�0|Q��7����?��y*�ʶ/�����V���Lw��;KR�1�2�M�X���l^v��Z?c��po���v��
&]�/#��1���Wכ�p��IW��񦾶��˧5^�Q/"w�}��c]_�l��^����w_����㓖�* X���NvF�}��'������,:�j��,;�2���q0���2��`�Թ�Rѩ��@�D��$�_�ӺA_�ق7%<�4C�o�t�_�TX�����e[Ϡ-��-�;x�����@�Q)f񴑱YR��7�*�31�K[�������@(�S�3��l�Ib�:�>�y��COiQw��Ξ�;��Z��}%;�����_��wA�7��?�m���� %�5�����I��#/�Oji��-T|_J�*������I㔾��g8�������_�؜70��XA�)ܿ��y
���B�*�j�QBY���@C���H�B�b�ג�^���$�F�3��|z�$�Z�&���Q���9 �^�S9G��(��vjX�I�$ɑj�GX�ǩp�����AH0���^@�e��|�R�Y��QEb������~%�V�T%tS����u��~L@��Q���&/F�|c�L�x�8*�`N�e��r2>�f�w 4&�b��Qs�$��B>����y�1*��������#j��]�K���MI�:]�@07j'�/���A%f����ۓ7�.\քRV�͢'N��	H`���'��P��q�C.eq`�j����p~[C�MK���_��噿����S��Y�uS*�C��j"��;�h|�c1�,}LR���YX-��$���Fr7$�z;�{7K|f�b�G �m#C&�O��)$��P0l� Qt5Γ�<�j?�Umm,������S#��������W�-}�ς���N�J1�i���J�p� �Y�P<�R�#F���I�:8�}��hC?8-�0��aW2d���Pz�h=����l!]#*�R.���r+���9���[[ϱf���ba��Rh��7R��(�|�����?Ŋ��0Z?Ɯ�$ ����XﳬXEQ��.�F�?�6�o��B�7Jڅ�ԛ,{�M�����^�32#{�?(`E|�V�ݛI70�J��c̙���Sa�	w����P��6��� ��󕙞��
O٬���	"&p��#�����wE /{Hrz0��~D.������r~Q<%�*�S�2@��C\w��~U���gL�K��W@;9{48�&C$)����2[)�3�-�T�����s��Iņa�'͵F(�'�ě�m�0[�t��_+A~<=f�7E���B�T�/X,��T-��Vհ��S�5�VQ#�"�����h^~�$}�ݿ�M ���̴󣊄�Ӊ_@���Mpf5(�	��[��T-�uE?fɚt
e�Hatg��i��>�%}���$������4��a�.O�5?�?PA?!*$�cG5e�?�_� =���V�l�_�j:u�a���j�X�y�#��Q�L/:#Ǥ�2X4v�Q�5�4GcxA�l����IxM���%Z��gw�N���mbo�x.?�{$e�!h����5�xNz�F�Ty@�������#S}���4�9��T�~Y����Xؽ�_��([ ��K�DX� ���Qqt�*�X���أ�b�KQ���Ȗ�D�����ۿ��a��A
9���oR'Մ�n\�E��"x�B��NcU��(��)��\ٶOv|s,dôoD�.M񔫩6z�Pf�ㄞ��Bi2��w���&�d�|Ȓ3X�3*K>����xF@�tS�n�C��)p�thZ�y5ӂ�Sv�S����|���x��a�q�t��i^��Yu]�Գ,��<�A[.��]N�jh��w3#�%g��*�6��J�g�??�A]��ާhQ�N��9c�Ps��`~��%a�<��7��:���\����"��� َ�Ὑ�̢���9�e��#4�PM�O��^���y���k[�Vv��ŔW�󊗧��D����\m�_C�W?o�<ɾRlq�˕�����/�]j��ojLH�T���(��婫�&;l$GP)h�hpY��'=QTd;��腰P]�nշs�j�u�QDGF��m6����w�^� ���~j����G},}XxFH!�O\N��,8�öke���E��"a�עwic����U�1��5��-L�!F,<�9$����l���-�>����Vf����F2���n�3L��e7@����ΑT��_�� ��Y���@a]h���F��7��.�Nٽ3���,9,��!�i
��<��q�����&qhW/�-"��ςW���DxT�~~�K��P��%�0 E%1�M>	�/y2_Vᱶ��	FL/�|WQr�BT��E�jw�z&ˏ���Q��m�|%�I�٪�A�Df��?��p�ո7WxQ��X�a�r��6�9��k���Gb�>��L��
ZMT!Ɨ��粐=�u�.�;bh���	N@+K��G[Ͽ�i�|����jH��=�}��c7�z�3�[�)����~�9�U�U��v.��u�z��T��S�"Š'��ZkźC�3k�ZB���M+S����<�Q�D�3rm���\[X�������$�@��1OV�y�F��R� �B~��ʵFPp/Ѓ�ф���o8���._��u�����9O�ڼ%��+0��gƜM�P�z[��ϭ
s���\=�����ئ�t�|_�V���H%����n�!���N�N�1�*�h��Dk1�����������1�ί���_'[v��s����K�\D� ���v���ӝ��lRy���C��m'�QL/[�u�;�x�8B5~�ĘAh���X���M1��
ҿ8�H`�T5�`��+��{�6�O��"nK>������7Oʭ��j�x�C�B�E���$�&��T7�l��N��(�3r�'챢V#^XI�������D�LC��c��w'��}h[�}��s��w��/�!��Uńh�Т�Y���~Q$0��%�k��%JI�R;!w&׽�Z۫��dvs{MЍ�e�Sژh�N��M~b�
DФg\��6qg%�+Ԓ6�\��8'��%E��d��0/s��"�>x�V=���;�v,I�S���-�Y��ָj�%$�8ˑ�����Ъ�r�?�.%{}YX�F��l]���$��5�.�k�0�i&n�[�_ঘ�0R��u�񝞊!��7�Vy�@̝li�Ȃ���%S\*u�Q��0�V�A2Kad���������?8��6�}��yrFNMS�%ix�r��f��\'�_ �ɜ��`�p��5	"�q���|���;y �掣d�.~���7L%E��D@��?�H�b�Lzh'���+�`��� ���7�g?������3��\u�Pct�}��
����'���M;�����h:��h��&N	�ݦ�j��|W���ӇL��y
��T�v4����w��6"��U�������F4���h=��$�[�#H~{}	5��O��Y�3��	~m<��hAK�UD�_IB�p���؋��<R��e�}���a��H����\"p�%f]�@���[�?(�S��#~�+d�@D��>��q慞�D2�|Y���ԡ�>內J�I�ۨz�4��;dm	��x��@LC)�+��g�P<�R����2oo���9H��EI�k�����O�������.b�y�m4w�8��C�Pl�Z�YM�j��Ve�L��LZ���g�¡�]]!�L��k���O���hfG2 f,n�G�����O���%��A��(5��!����{X�١�>�$ʎ��5�9�Tӡ��8����2���g��`ej�g��>0����(S^��ՒV��6/!M���>W^߈m-\&�D�T��y���Î_.w&��b�g��B��8�@�;����K���g��\�`���t��������qG^cW}�3N�!1�3@��a�6����!Wf��I {I,�hy�	t+��[]��~�2a�$N�3M��4�:��Ӓ�)$.�`�D�Jo[v�&�n��{���A�:���]P@$=��bdW�����C-H�� Ë��
��
r/���85�Tb�&-�e��n��t���Ӷ��x(gA�b)�U΁�3�߇�^Fs�%���&�[~�z���:��y�ί��ˍ�]V�R��t>���>R�L<l�6 ���x�?lÏE$�U�4���Y��/������4k�{�9r4�z���~2%@�3_s:B�UML�qՇ�kz���T�xo��䱬&�Q+]��U����%ԉ$�K�A���
�3+g(��-����/]� $�}]�$��=�Ep��y�B�vg1��^d�+z����2�9wa3vVI�����=�Ok���\	��_�n(���CW��ddF�}��:��}�ݹ�I$��:r7�H��3?>��B�h���r!�p6NN���s�k�v[�TTЎ(t�'#c�~�6�41/і�=V2;�|�8�G%�m�MN�V��<+�Pb��9ot��ܴ~�Q#����Y/U�Zpʧ�Z���>P��{�p�7�O"�GF6�A+�ܟ�n�U<Ќ6I_���uP}�`8�aC0^�/$H�	`�*-����`�Pf�����!�ԥ�/Y+J���{��~}��r��HOŤ,+���$ob��6��6��L_9B�@���O?/I`�7\�l�+��y�^04�����3�g�L��K�LN`�Ӻ�7��J\ne��q_z:I� 2�#|���75<7� Z���m�[_�ks�{;!�!�zmK�zR6�{#��L`��o�=궑���}�3�V9� ����í�� ȑ�m.u�Lzco���Ԓ>�LO��x&�;�\n�17m�5F�>-Ss��m:@z���s�%�����fn�6�
?�_��G��u���$��O,�p�. p�s)Ć� �mr��W4���W_��X�C�j��<�*=�>�g������X�Pq�e������H
��8���}q�^����9.�^6��~8�ۀ���g앢��f������� P*G�W���m�~{�K�~��⶗]�m��y"DD�3T����揉�p�M�ח v������������{\x�,��lQ' D������Z0S
�!�V�E�j��N*-��z���[>O����w��R�����t���
bL�_^�TzOg�������㐧C�݂^���^;�7~�TF�Щht�:[m�5Sw�l�x��,jvt�|K�өa���m?n����ѷ�_�Ӡ�H��~n�p>-���Tf��R1�-J>1R�C�R��=(���RM���y{3��g�@*	��"�\�b�jD�AWÍ;�C1o��F�T�.�u����o��b8��r]���t�'D9ל�S�V.~��0+!�DT�lpC�EF��|�I:��1�ĝ��l߲V�$��H����-;�'P��c�YZ�&�\9�'��G΍������KL����*Uf��0��E�������L��mWG�?��6����:Y{[)4�ᇣ�>ˮ�{����sK/�P>��/�����Ћ�/�d�nZ�/�8��㤰j�ݓ	Ok\�.�s�#�B?)v�O�rO���l� ��夭�
L՜v]��RI<�����-j݌��>�&�.�3Zv����q��T�1'Y��*L�D���/UKO]�1Zl2O?�Eq/�-u9Hf���v�;�u:��Y�{}~��� 9&n��.���c�N��0��%�!_%vU���V�l��p�|��<��D;כ��s
��Ϡ�����}��k�5��	�a�SW��0r��pF��skx�����p��dj��_�GpS>e��� /����Y��#i�����Ds���㓑�cZ	�(w�\S�����׽9����j�G,��������qл�稿�Jd&C�����=ǗI�K�x
�j�]���<���E4a�p����1�zܕ�>��V��8�R�;��=.��܃�^eGI���Y�(Ep�xL^r�x�䬉��<���xLoA'w�q�G��_��&8�4!���)���vU� < K�ΐV�}���%�����מg]3u]1u*?��d/uA������:��ĉ��C�mΫ��@�7���*h�GI��(�� ��nC:}������S��b�Q�a3Mv陼�ϔQ�8JVic[��Ts��9�R�{N����}Z`!�%��;���-�x�!�i#	�����_��0���&��d%�ku �`��Gә����_�#:3Nّ�'f��~	��/��Ds)��4������G��L��5�q��N�l"#��?J��I���j����&�s:�E�	�]A����|�	r���F|(_2uj��3`˹T��������R���ͼ1��?(�
ÿ�Ͼ����o��gP��t�ި�F���]�d`F~�7�WS������4�ayF,~'��QjEK�k�Jb��u��8��C��h�~�b;E(��cUf�p+��O��u̮͊����EKƸ�qۦ�϶e�,P+��>�(�G�e[7�-�We)���}��/w7VZ'2E5�Q��ac���%�Nr�N���=ٽ����x�r�9�@&��}�6ϱ/4��%)B����Ф���ك�]ր'z�m$B�F�Nϋ����D���%V�\�^�aH��I�����a* �MI<�n�=˞=�>ɾ{��ݑ�u����̪��Ķ-0���Ӫ;�z��Tz��!o�Q{��"��z��=�V@����9w}y���ba)3�κF�%���r��eB�:��R���#��9�n[D�'/��p80Hzq�8�/��nԒ	�5·���b����i�&�2��V_z|=݇O�a'���Bj D��S��]j��$P�P�蕯4˜_D��ԙ��2��yNP��n�����HNq��ڿ �y��,N�$��#����֭��4��eWܔ���" Ʊ��;[�r})�ںд���fg�`�B!����nG���b?�\���{��Io7���o~M�Nh��f�vസy�<��v�'�5
��Ra{jmc<�&�����&��s� ���B?��<��UN�A�7��:�������@�|�R�N	�S3���k�L?C�1�7b�IDU)�DY/�i�
괂��G,���U�d�1>���Nr�;Vg`�Sm�ΗV��ʙ�^��3�I�H 
��� �C��T����VBeB,Q�,��6o�:!K=��5�?	�^Srs]ku:�EF�9��������KV��w#NS^�2�13G`��i1W[CZȣī+�{������بf���:)>�w�:^�D���=�����&-Hr��:�I$r%@1\��y?:�n�)��!����EL˿���Q~��}K,�^'V�:�W6�-A(���7A����7���%jsLe�Sϡ6�kU,��DɣDww5 �TU�i��YE�#i��ǰ;|��NV-�b꜐���Sf�'�����0�h�g0&q7u�G6:I72�&��\G�����g"Ŝ���P�i��#�h��SXi�W��ON�lb�����������}q<��U�����o�z6ZC��B"Ng�������Y0W ɰ$�7�&%��a��9��H�K�Q5�a�lAQ6?�G�?�(�M8D/�k�iD
�[c]�o�k(���]����*\���'�Oĵ����K?�(�/e�^����VƏSR�5Aۺ飝������lꠡ�a+˭G��$����쓆, E�/+�ӂ'C0Ka��M�.�]��.tg�叐��a����K���L��I�f�%v?�t-�u���J���He��k� �M3��~�Ȣ���|!��q&������R5������	&xqLv#�υt��z|�m ���74�Tƨ�5�%��F��ȥ�Ɂ,�3��)� ���Y�_��aV/�6�_H�*�Q��i	�E����^3V�#����	�U�X0����B�a��}�{i�$FuR����ky A��퐣Jɶ��`�Q�ǵS�Hcӥ�0`��L�Z �ٳ@��B��7��xEC�r&4O�iٓ˶Z�U�D7�O��_����W�Tx�m��X1��h���~�_L?�v��0ߟ@�5t�Sޤ�4Q�RQ�� z�q�)��O�1�b
DcCPV�p?M;Ð� )�}�� Y:��h`D��S��f����qc�6�7�(9?����r%�8�s#�j�BM��d0�Ҕ/��:�x:z�u��f�s�ø\�4q����َx�ҿv(Y���tlщ �}%'.��:���X���q���b�)T��X<\ ��rΔ���"�Q��?<ڣY�4E��.Ƥ�87:����ə�E�Z�ǜ��Rl[�r��:{�JI�y��ӟ��i��*ba��9$窉,�{඾mZ�6���xڋ�x�}w��2pn)��տ�ˮ�3�Ш3�y����gɠ�5���;���>�`65�ʚ�B���R�5 Xph�S��F����~�|D���0YmE�)��a�:��c��{1�э��-Б����0��t��7\/����Q$'�����#�PċKICJ�f��1�H�^��f[J�.�S�\�g�rS���Ӝi�J{�~�f��hqgj��i�]B�I'�Xvׯ�����e`rN,m��<�C�n��`6����̙q��cu��p��]c�Tt�ܴ��'�h�,�U߃E	ݾ�B!��$&N,�7s~���>�P����f:�<���ޟ��L��.g�m�v�9;�������ewA p�QZ����)L��h ���{m�l���|Z^��)�P��+(��$����;��[����x�%*�p�M6�r��'��ovI��vw�\\���D� C+�����g��������|dja�S;P��~��D&���&{$��:�a6���	^����2c5��bV�ct�"*�k�u�x�
�s�X��d�^��+���sEQ��8�k�EY�VsHT�	?)�dهn����#��j�+2�A�tLb�c��?��#�.V/X���)·��'��͞@d鍳��r	�`X[n���|԰u��.+��<�{��R!w*D�U����t�"3�cj.�uh���¨�4��b�܁�����jV6_P�n�.���|�}�ӡ�5Hp��j+�xȝD=�L���� {d�v�`��%0qM�{��a{�3��~~��!�J}�bT�T�?�s���L;�;�vԲ�*T{�`g9�:;��别 �]aB&�M�ܟ��.��JS6�eKz��ϡ&�Y�T��؎.�zz}Z	�噪�&'��m�tN^y�/�VK�IZ�֜���e�Y�􅀕W�/���_�֨�FN�l����\�4���S�~Q��GHh�=b��J�kc����~��U��ݰ��q������lːِ��h�Ӻ���3r�sԩy�Ο�d*�~j�/�F.��9�YlK��?��nbW��.^F����u��ipb�_�L�;���59�8�y�4�S��ߊ��z�M�!I�ݵ�o� n���ʫ�a�B���~���C?��ߨ�L��鼰�S�6șJ��a���<��SyݼT�A�xh� ,�ה8,�9�݇�n�Y����A��J��A'*_��\l�]"rX�ފ|�v��z�;1���09cK^�`� �1A,K�|����sq?�w)����Sut���h	��Pۅ�Vd�����|TG_��܍�-Kjܧ9�1d(�P�s��!=�k/����oˍ�����?��Q{/�ewZ��M9�`�6�AvP�'�[&�SRN�Yl*EU�:B0��U{�=�?/��X�g��:T�ˠNf躙D.Y���S��<\�Ͽa"�[ۂnF�J[]|��h펎f ����V��k�'	\@2(�z�
]���ңD�i����oi�����k�'�^g����i�8��t
Y4���¸������A�Q���vkGUy)A��˰O����n�K"�1/MN-�n�`�J�ZJ�[K��K���	,=���)����@2�W2�0LZ,���JyWz�Y_aO�A�����UeF؅U�1�i���4���f�s��ن���
f渣�H0�"��;�T֬Uv���YW%�q ˃k6ˍQɗ�����ͺU��P'1�9y�]��dTK�WX���|�!��4��3_�&��Q���5����ڌT>����4�VC���Wr��y�3S�����k�]��3U��QJH>W	I<x�\W�Z�������l����.���tQ��
T�Z}�
p|��$�MhJxr�v��|�8	���T�e�ۼO��Tb��z��G>k�qQ8�B;U���sȦ��4�b�@/��>fm​���_j���ws5b�����šjL?�Q�d�:�1�l���?�{��^��y�wk��&ȩt�Ñl�ԕ=��40)w��`��_���Ԡ�x@�NM$q58�7ܞB�6$�y��<gu Z�c�2=���l��63kι�F� �,�(vd���������k�+I����Sc�#:����B��m�	6s���ַd����0��Ob7d�m<3	��� I�w^��&�lRf�DƆգ3��H�z���*'6TPˈ�w�¬?�mY ���!:�-8=pȽ/���Ac�;WN\7]/P9̗Д��m���Ý�Y��>�&M��oi�H�1J���SmG?5���Y4���U��eB��O1QnZ�,�e6C����=I��$}}w�m��27-P�e��"����Kt���N)oՖ;\팄�b/��^)yӭl�K�hw�<L�3�2K��{̩]��''�=6?Rf�h (�>� ��d�˚H��:Z�<���<q4Jd��G�U�7EO���{���%�q�����{`��v�D/�5�����=�ub�'�h�*��#4n���j�Rp�-9}��	zG��� ���W�~\f�k�P/j;g�(�u�T����>�Ӽ����)�\�sV�@��a��Hw�JcӇo���\�����_��(�2K0s�>����4�����0�bgd�0���������w#G7v��W�+K2=�^��hq�AuԒW� �]��4w�S������Z=#�e�E�%J��T���1�r��bj�D�IZb\��#u���-ny���PM�I:=��d'U�|�Bi��B�3�4� ���Z
G��l�Ҁ����3�w���05ٙij��&�E�fQ�8�I����7��9��? �]VPX�.|���Gcj5x��cv�wF?N6����փ2��ˉ�}6���?�x���rC+�X���k���u:9�Œ�ޚ8���~�
�e`:�P!ͻ��(Z�G�ف�ܥ_�M�����3ԥ�~
!��@l6�������#�q�Mo�}�� �c0��ϛ�>cv|/��H*Z�z�ܻ��Y����ݠ�l�_�!�>N���zvv]��T�� 85���z���Nnj@����
�Y�E�r�ڦ��g�.�IFM8�8eN�9 -���ChH�%�1Y �I\��vr'�˓ȑ�DA2���wŭ��dNK{��)�N� g��!�@v�-,�VU�+!��7.��*� �� ��)`�L
|x?7��-q��퓁%=Z�)�Џ��@Ni��	Q����Cx���,����=�뼱�a�wSB�M����N�	Q���!b�Dm��}*&v�����)�d�$V5g���k����C�ZL!�Gݨ�w��+�.�w�7��ᩒz����>��F�5UN���@^h�9�R��8A�9�#��Byx��O��`ׄ�v j8
!�C��J'�'��3	:{��gy�|�ɦ(=�nJJ��F��w�M'l��KXfBDc���	��� ���ˋ9�t�]x�z����'�W�y�]r9f�jjֆI1+�6@D!u�Ѭ�w`�m����\�g�̧�)��a�I��G�1�7�4��<R�s�E�M[��u#ػd* �?Δ(d���!B���������?aTn����8s�Gp| ���-qĉ��h��/�/��cH�Y��@���?��o���%�������\Wq}&y������t���1o�D����`א�F�,�
R��^�ɴ>h�Ǉ�@c��_��+�=٫0z�V�$M�����m���Tz�E{O�8L����;�!������Ai-G�4��C-s�VPZ��}`���wN}�����h7��O��#�n@�s�gvQX���VT�S0��g6;e��@jG�Ռ�#�8{풶nϖ�}�I��@Q"�۹�u=Gh�@>^�Z$o��h�)%d���h6ꛢ���{�I�< ����/�_�B��1B�(Zm萫.���b
�U(�?��cK�%պ���w���P��/-b����g����1�tXh.����9g����c�t��
�H�*��ι��f���u�l�t��3V��V&4�XH��Ǡ����mO)!�Ŗ�Z<74Л�3J�,��7E�\�(_�(2��V*��|�"F�. ����K�*��\�|�����cЊ�0���aT>�P?�TC��a��O�_nHb����c�{�2H�bw�tC+#RE�GM��Q��Wh��	�N�BM>pT%��4��{�g_</T�Y�d1��O��!9-�\وN�7�I׺0ޯ��땞�j��@E�!T�`ۥ��7p��[�1�l?�#��d��|S�J��>���9`����ru\����ߊs3,����$���1���LR�ds�h�~������	�Qy#I@�9mL��*]��Ŏ�����Zr.����sT�c>C`��M@͹�)Y������M�m��������e:96V���o���^����Z��Nh�� 3J�潥�W�N��'3��xg�n#'4�{rj�:6esj�О��Y;2����S���HĆݴ�^7-�H��l\L�t��Ok2���#��/_�����>����FW���vp�f-�!Ԧ����c�
{��v�~�4�ͪr�ݩ(��k���+����M�� =�/�ܮi��3����Dx�Y�I�pd��6�ҿ X�r|�R�J�}�2�%g��g�	���i�t\P��x�vǡL:�P��$��蚁L���S��WS�22V�K�5��X?��(���(�;������
?'�Ϗ'������y�mE=z���7K�Ӵᕞ����Y[���vص�(���^��t��Z\�b@�w?v�h���m�V;̍��}\�Sh�r�����v{I��Zc[>�H��v�7B���v��H�~�H��&9�����"�����4�|ZQ[	Bcr�A
��P{����'�&��#>���'s��b`Aw�kuq	7�m�#���f!F2VA��Qd���hw��4��-�|�̄K�� �퉰Q*����z���b��`�vr�n*�����d��t�Q�*O\�����G�VEB94�#����3�kU�]笡�cMS(u�L`l���/N�azR����;�G9f^�A@��UaA:�rq\�v�6�ݢ�܍��Ȓ7�m���	+����@��X��.z�r�аi�G}<m�B��E�XQ7ʵ����FY��y��"̏�Ik���k���=�ww�g?�m����l���w�2��1�8�h˶��s8|s���!⮴�A�f�{~"{ӯHs�>���2�D�W�='!�O%�+�a7������*_� ���zubA!'7�c��_v��;E������7<o%�5ʫ�	5��U?v�>�
���P<�7���dX�7
��g�|ü��ߧU�+��~e�;dS�">;��_eA�k�A����J�M�g���UW��͍{�R<�',����*��ͣ�<�-΂$�{Q`�;��gZ�Z�73`lbF�����q�����hS�^,/=��]��=[6��
3��=�(��7U�4����][��������Zw[�Z9�>t�c_�!L�-A�A����x�{+��sJ䪏з����[A�$�kf8}��������;�Ƀ�P� ��\���L�Jx��&͆���3��w�"�,�����F�c��^����SYk?.�Q��̇Loޖ�1F:�.:� Q`�#7ET�W�����R\�8Hz{���|8Bm�y�}�p�F��Z�H�����2Am��?<,�9�3�M{�v�|p�
0Ȋ�Tq�l�Mp�M�)��,^���1>G�(A���Q����&ڡ߉ciMU���PِK[��p��	�r{8yնV]5h
n�p%�5M�0��X#и�@ᑠ.�6�*���r�/��ge�r`���uhj4�d��q�M����r"��4�C񲜝c?o��m���i������T��瑴-m��� ���HJՃ��v�@���%s<1���R�c/�5ak���_0�g�n-�r��kTc���iF[{z� ����]ųY��~lʹe�o��n Y\��{md�}>��`ĝ'��Ǌ���*���r^�J�3!��<{uy�ak���L�0y���Ks�}���/��q��bE4����-���'PW�)�a�t��T=(&�;0|hY�vS�� ��e���?ڄƉ�oC�^����;�kوrf�u�3��Ջ��B2�.�ag�#�8�GU'C�D �ę�ؙ����-���1`�_>K_�]� =����mڛ1�'���Rd�͓�*�jHe=��eK)�A�d��8(��Lw�#y�sL(�<o u��K.H{��'9U*u�c<G3��nIs�`y��'����%ۃ���^%B��\��L��|�U�I����t�B�;C�� D0'b1Ϲ��ÿ�e\AJ1o����u95K��m߸1G���:GW4��b�nA��w�8�Z1 �N��� ���n �^b��&��]�ո���,H�X�;t]�udEZ�&��0�{�αwc�sʪ��z��㆟VM�Ǉ�5}M�������$����\�Л��K���wJ$�����%��j�3���NE[u�(u��
�t�-���{ ( ������3 z�������L����Y��=Cf�ۗ�/]Q���-d� �yC+����\GW��>w��Mٹ�VgV7g��
I{��D�>�0�Ƿ53s��q.�,{�r�#�O��-�ݱ	�k��}�kR��g�p�JW����ʤ��W��)Sk�y�"�c6e`ى~��	�N�������%��A��Ww�u��oW�ˠ�-��],Ge�Y��Q�)�z��#��@���+�n͎П�?z�o[vP@4H㕝U���݃�d����)��l5�	Q�3�Wܞ~ͽ%� �����۬"㘮�<����jR�߸�1������=�ͽ�H����9�'.����	�&V-�AVt�S��:�'am=��KH�U�����:�Gf���}��ٿ����W�T�j@M_q=,^|�%�	y��K���E�X�D�K~�}���]���b�f^.��4������]�����y�"��u�L����߳��_wY�hg� ~V~�;A�6Y:H�F���i�Q� ��D���s\�ҋ!t�!����6�e1ҩbO�Z���4礤��O]��,[����~»ƚb�Pv��xJ�M�jn����!�|��T��ĭn�E��V�̹l��d��af�,���a8�/��{��o��MP��e8������>��ɑ��-�2�[�+No�6�e�􉝮0��r�ְ�\����?���w.�6����\�g�J1g�����yxV���X���E�2B���=�?�D�X�G�g��N7��G����k�}�K|}r%uX��SN|�;Ih��ѝ��S�c�H5Tn�B�o�cV��Zy�^�v�0-�k��*f���K{�L<�}����[Fɒ9[���a��;�t(��q<=Ïxg��ʏK]	I;����~l��Es6��<sj��!Y������������q��J9����P���U.�X��s\�'�Ć�=��꾓{y۳��㐫�Ζ
k��ٶ�Z��م���w�N/�xMoM��~�d���}�5����I@���������{+�}6dB�|D��1"��"�,�������	)mՐ��S]�@���ø\h�+7P\�������#���=���o� �(���/K��Y9�e��I�d��"�ҊLE����"'���t�c&h�uU��s���TcR7˙�vPO����6i���C4����F%��#}�(�Z�*?���D��v��&H�cc�$M:��6|U�rTp߹a ����
7���H��2���1�m9?܌�j�.��~GⳀ��n�s�lə65P�#ClgϦ��`l�a��sa_���<Ŭ�M�,y~��1qn1�s�4i�y8|�>GE��9��aj�m�SЋ�'�ty�%E�rMGD@�w�sHkR�F�-��Q�0�FU�IAʋo,γ�ƭ�o��U��9}�:h_�MX��[!�(}�>RD*�W�����c�Q����<ә$r�G�׵@����a���ѐ@!R�.�b̿�=<�C�Qxm��|X��d� ��u�i�Œ���>��S)=>|Jp�o�:[�#~'���n2�MK��*{^ ��� ��v��7f@�+�b���1q�����`ϤC�?X�J_�>O��0!Htܩ������?�<m���Y��pg~��9\����tP����,�v'�(K�J����Ǟ�=L�2l��O"v�]�r6�Ęj�
z��! 5�K��n~����<z�B[�Z6�7�W�U�!m1
��.�x=�=�}��W�� �t��<\���_(�����s���x}$.X9��t�[��N���p��qX��� ��,�=�ߣ����׺�%��秛�	�؋�`\ �{G�/B�B���OM��G� ���C]L~�}�^T!"[/6���,N	�Wq
z'��(�ll0��;�$7��Fi���X1���$�� �-|��,����V�v� ⫵�n��O���Ǥtg�������,%��]������ �@s��װE;��F����� ��[�8�p��r���r�RZ.}��`�����k-�\�T�`b_x�v����  
���>��ޱM��0��T�k3)�\=�U-���(�U�I�4v4~��=����6�ϞI���_ �m(']A���Gg�NL��[��7��X҃��r��"R籪��B�m��*%�Pv�h&K���ғ�3t��c{�Wl�r9��FL�!��25%#��j�pI�`S��hL�����[w�WaEQ�w��9eڣN�J+A��x�
L�٬�|DU�!��q���]o�����Y\l��e0ڼ^p�V�y>��w��q�ծ�{ =���i��j�\X�iN�n�a'@�����+V�b9l�J�4Э6�dky����3�OR�y(�㷒�KJ������f�_#U,��)���%4��q��������+u�ޝ��!���^3�6vt	O��A�"4L���v� �0z�t��&�&w��v���hK��Ȟ+�Tǘ.�m2{Ӊ"����|�I�Xr��q}H�p� LD�p(d��/վ��1�R�o ��Π�� ���4I�f}(��p��>�gyJ�����X��[�gf~�7��	1zxtcÙ��4�&i��#���T�
�v�<O��,�B�����d�'��c��l�C��t�"��۷i�[��9_���3��ʥ�\֣��(�	�I6�����+��e�T@됃T��A��/�`x0�ki[-����5;i�mV���}-ߒ��K>q�:9}��LE�.�-�.�lyU�A���'�*�<>�x�d;/�N`E7�"�Lsk�a�s�&��8�م�I�� S��i��N�n�����a2xG���m<�����p�5`�i6���u��Ë���X�-�Ȁ!.�hF16͊M�\AD��uU���%ا��4�Z���gö4� E�)Z����hg��da�t����z���\�;劎_��2��CPܮ)��/��9
�6Oޙ����4���*��]�w���F�k^���
j�������Rn��o\G���H ���p@;p} �^�	����۱���������9D�0j�0���=�(��.��v���H5�0E�I뎸��W�p�]ޙ� Fآܷ$) T�����<�B_?��w����GNT��~3��H��]�zR�7P�4���: ��!Q��Fa5һu+�:_�����qޘ>ތ\��m��#2��O	_t��fZ�NH�Gq3�~�?�<�\ӿ���'�A�;[�K=}Ng��)MEB�TK//�ԉ7��[,��2��J��� ���H�<j�/;�����z�(D�;�|���~n�J ����iyB�Z<���j�ڂ�YN�j��� i���&\�_�3�����2�,-��E��]�|��7��ms�!��-opTO��n�z�Va���*�"�.9�c�8Ha���h���yf5��B����W�05�������0�A����E�Did_���j~>����hMȄ�'��z����zq��[ �dXiy��M"�S�_��k�n�X�ݵ�Gn2͏K'�#�Ȯ��	��cHf_Ƨ��]���T�xIû�.3iOW���!MN4k���>Iٷ<�w�"��1�����L1��@���o��B�����%�{g��8�k)��AP��&�"~D{2R�� n�� -���Rz:�_�>����!,��%S@��Z�-�f���S' �c�z��������	++��^i�7=QE<]��z�cY2�r�O��vHch4"��oR�g�Ɩ>ދ�u����w�DT7\;
�'"�z��*�EH}�<�}mV|��w���ПO7��0"$X�A&����ӅW�5f��@`i,�^ϰ��zf�X�8�L���O4�X-�����=���o�65���fJ����o{*,�#���K��H!�d�%q��K:�Nɷ[8#ž���m�l��@�p���;�a��"qSr��WD��h�g��D�0=�`�+����1�;xW?�zH*�{Hꏵ��vQTF�4��"M)܈��v?��.���p�\�V�\ �.t���/}=�0N��q#�����t����!�ec�/�3�i��m��e'�}�Fri#nv���ı��� 5&*�ט�Fxe!7v�g=�A��u)�R��L�^Q�e���7����=;�_j�&��
� 8z�!��$�����J�<^��
؄R��,eT�n�Jm�����;PD��C!AN�_s]��E�M֋=̫N��l��R zKӂZ��x�*���M��q�`�ߒ�d��;�O$t]��[f+���C���v��JCg�7��%N��A!��~`�OQē#���b�hcp0� 4��fe;����7ac>��qb�:�%Z�gY6�2 |��סvt�m׎C��o,mg�ͺL7�e[�#��(�سR�~���m���n�M��<�A�NVty�5�(��dۡ4�����Z\�$3�ύ��m��M��XZ�G��wD��m-O7��}���UW�A��}��HGx5�ӝf懐����~��f=w�%S�=pz�F�����i �}�;������苓�����+��²f����<;����~�^? ���8�y��k���3���7����P|�	�#5��"�D�����3��2�x0:��C�zPh%����������_p���ؗ��uy�A�J�Q��"�S�IE'�΀�6�4A�����I@&�B���_I+�����y=��+�ӑ毑G�B݃F�r7��Xpf{�
~��mrHٴ9���0�v��f���PV�_����~(�]�V��t���Gߚ"����Q$h�g8i�Q��������߆d��{���+�E��Q4��f��戗6F^*&\�P�_��K��Hk�S�������~N1���Q7���^:ǟ��'^�N�pg��
���Z����Eu��S�2Ab����3(�mpV4�ע{�4�%�o�y�h��\V,7[�sӽ������>��a�S��
�x���5����FS��&�H�ٌ�+��p��'�$���+rt�g�|.TU?��rh�jQJ��v\j����1;��b��$��.��t8�c'��LrF_��Q�c�ȵ��>�	tL-��z=���..���`6�/���b;1�����):�
$�k)�p�x�06%����^��B�|>�7u���Ej��ͩGKNh�2�����[x=�1~W���c���h�k�G�̥D�7$t`1|S/���Q= ���͞��=�������l#JV�j������κ�@�r��C��ej��|N�:ưb%�8y��xC`�4����Y�Ԉ[b�zh)��Q������XO��H)��lȳ*椀�N�>8�)��Z'�	��'���NR'.b���L[���0�@2~�Ja[���-6Iq��8��ӽ���c�.�������)�[�]:Ģ��@_&t:ΌǑ8ݘ�bS�E�.���M�v���܂��ٱ+��!M�>�F�Z��Ȟ$��F�V��o����Tէ�,��lҩqϹ���^�@+�6"v&��D��Nʄѥ�"��L�+nt(��C�q�|�m��6�����95j=���	_n�XU\hn�T�G��7U�|�ÑBa��^Є��r�۸�d�t6cKY��6b��10V���0���'bl.�Sn�O��~�Tl�Bǧ��1"`�)\;F�Ľ�4�K������ W;)��j��K��d\}���|�z)�5A�fB�g^�r�g�^�����-Yx�+u��\.l�W(�H��F�?�a�>U�,��TSs��^`+�{:�C���f�郮�����Qj�c�y������z]C�Sp%��U�ޗ��`��0 )��	#F#�K9�s�E�G��7Ok���'��Z����+���C˛���'{3*��S^�sq�p@Ĭ	���z�W��jlH�����~�6
�T�81T1H����':U�:=�99���hf˚�yj��y��*2�~�M��=7�b�f7��D�����0dv�&���N@�Y�[�{_zUJ�Q�'F�%o!c�E[Ҟ�o�XV����D�<�T'o�$C�>��C�M���^�X�x�����\��܄p։�ti"����O��s�m�ȅ���S�� .Ǎm��g���K�ofD���Vs�ߠ�;�^s��E����c���#8�����%�%�A�blm����|¬QK�<��9�e=�TEb�w��Z���*G�v_�ŭ؃yPy���ClZ��Ad�v�r�]EII��vrK�F{l}���"s��F�X��IN��kRms����������"�Xg��GFf}���.���+�0l����c�d�7é���[�i"l��zZ-	�=�<�9_��=;��a��m;�h�e�� �"�u��t�Eg��2�N=Jܚ���4�Q_~��BY��m���*Gws���e^�̳�2b<��0�p9�Mp4ͦ6�$�D�#z��^�� �*,�+C��N$O�$męO���SO���Mׯ��H���7~_���0/�Z\_�C���-��M�.t����Q�ܭ�R�=g�Ȝe��㍇!����#����&�����Rʃ�&�(�=h�oz�R���H#עN� j��p���A?����� �t�M�JP%<�&�Y��4�R�zk �4����?Ո;Ӏ�l��LoE��K�{�N����^��3L��4d{%�!��ī˞�)��MɗH	���7��~����j�#�v�� �ޑ�uyA� �+�; |���8�Hc�
�{U�����%V������)�9��ۤ����j0�`����P�TD�0����B~�������t�\�6�0x��JΏ�j.!.�������jI*+��ӱQ��6a8	��1b{\2T9������$�_�&sB?�'[�-^������섍/��!\���6��#=;�A�^ĹɗYe.����k�b����ua�㥌��� �yݧG���e����"��9��}��u���q��in���Ș0T=@�[�ʠ�?�qv�+PK2`�g�Ϋ��X:-75��`"��Dg�x#�u�r.O_���^�̓N�XL	�QW�v�G'k=�u��B\����<�|^˨3��K�Q��p�:�Prl*$�i,�����_�!��Dc�p6�&���R66ҫ2�u�oR$6`uz�LE��3v�ze#Z#�7,$R��U$��~y��q�4�_Ի�w~�ց^6Sw/6�D���7j8��o$_U��Vf]�	-��qdP��t�Y���3K�XD��#֦��!�h���w\��0@q R����dm���؞��&PUN�oN��P��
)"���1�������!L�
L��!u)i��1F�<�S�hVe=�<�s���'CN-&$�=�;�%>����qT�%e�É�.NY��oa�h2�=�3�zH�b3~@-�:��Թ���(�u�^I���5|�6�-y�P�D��\�X) 4����î��x���K&R�''M��$R�oc��
i<�J����0fߐP�\2�l`y��A�Π޺�'���9��)��BZ�q�mWdۃ8)җr��$E���g5�ʒ�$�~L�^-/��9Cp,�uN��s��[��j	P:C j���ys�R`* �^%�]J_�P��h�3�U�Նc�}u���)���	�R�j����r]Kk��B��hc��vj��d�Q\^��Y�( @5�а՟���۴R����*[��3��y��O�[I��Y|)0f�'�d��"��z��=���G��6h^k�@Q�(�����J�r��xw���ˍ��w�s���Y�!���M{��Qz���������j�ڥ�T�3�pv���3�;��ф6x��g^���Zq]��h��2�,A��nm�͜c���x�1����H�&9`n�Z�	j4��^a��!�}����r6/J�g��8�S�d�B���cg�ܳ��`�D�\��I~��h��=���@񲆋��k�0�vjRc�,��]��kȆ�ic�`"�Ȑub�_^/��� �"�q��u[�d:T����nP���V�L��|�	�����#�˺�LA�Bt�Pu�n����@g����.��B*���'��{��g�C�Yj����7�k�e@�%���c	 ��2:���j�H�����K�AÁ,��ph7/���0����m��w�K����_�릕�K�v��K	C�0&��οA��C�nѶ���:`��R�MP���}��fgrZ���<��뚾�{v�vT�S�B��!������рh�j�V��E3�
`X��8
K>W���FzHuO6pp2�Y��0uf_56c����n��ʍÚ�ހ����+���������S��b���r�3�ʦsL�<ƓH�J\�n޼^�˖�),7�JN+)г��U��w�4]J����Z8\~�VR��P�\;�~��դ�жE�i�����SUׁ��y�("���ЕZ�ÙhV��(&�A�� q�T/k�b�T-�Y]{)q*4����gs��5��Z��7|���_�.p��q1�g��+$���;��S5~}�t����Kݮ*�����:H�X�8Yaj/jK�����yd�;�1�a~i��*b{{?fa��n�Ac��KH���P��r�ř�,�V���&R�d��!����.)���=��Qh�i�Z�C���$?����֌�=y�Ti���N=��$R���H�@��������6ݵ�+��k���	��*������&$��=	\�->81P,�J������p=�	�nK�U����)6ԛv�xT��C��zn_Y�3aռ�p���?�j�C��,�6�g=D��E��n�������n%�FNlA �1�A����@�{؉�"�	b���{/ ��i��OW6�&����V�;6�A"sg�.��"��h�y��zP�Cx��=c�{�ܝ��D��"!P��#>ҟѩTÛH�Ṇk�p��1��\]�5{9�2�ȶ&��T�Rr��kǰ�B� �/ݻ��س���j¼_�Fb- �4K��I5ի,�J��ͦ[z~��P����L�'U��/�v� z4Q�?`�}�@�y��v�$<nv���a�%O��E�QO�W<07x��|�<3O��2>4'�2˹Eu�{j8C�*��1����\�0X"<�_#76P�}��C���Z�v\G�����C���,�Ikmv|5�Օ����~y"p�N��f�Ɏ�������r@5B<}�Ξ��$�!r4�U�Y/�
�bƖ��S� sl����7v�����l'�L�AD�P1=A�p�$�nJ0�I�YS�^�K]z����/1�"yXa_��_Ƃ=�>������u_�L��p�h�м��G3�<��m>1i�Ȑ���z-;�֗��;�)
�*�����J��<k�QfR�y�W��Q���Bם�B�k��;���_��ִ�,DN������ܴ�O?��e;wO�-�๒���,�
�`&X�ǁ�H��L}·+21�Lp0v�ur�CҔ�֪��m��CaR~*S����s��Ξ�������V��Aߡd����$��M�}B���n�8c�h��|n�.TP�����1p���`M��k.5n�A󈭘?{��k�i��3R0Ȩ�������s;�{�6µv>]��ޤ����73�4!��9�1��RΔ'Յ���������R���Y)�i���� k��F��,ˎ�t*eL� r�r^y��>�;'�GvvC�M�U���l�Y\4�Ҋv�r�����-g

Lu--^�Z�%�x�p�_ʭ�<��!F
V�=��-�<���<LֿA���7ެ��͢�k$p��?��#L�ݦ�z2,p���>@�e3�U<�QdY��� �b���6��65������:^$CI7oŹ�=]M�ɧ&��Hq��!0R)f6~�$l;1�_/�3�p�ѻ?*���n���}���n�%�����,����U�}�{�R��٢��y��N��Ԙ������;xǧ�m��<X�X2jh��ӆ^�*��{ñ�7���0��aG��A$&Aw�*lѥ���9��4r@�l�`p$n�;�D�Q��9�8���y][)0�%ż��#5N(
t�'DQbZ��>*Ob�vw}j��}��鍐��������� @��RM`������֣l(�.�H
�t����U �)qA��^�`mb�1A�f1}���{�w\��D����y
)E�?u�;���[��Ē���.{9eK�ݘ}@��J�V�N��VM��}��� 'AL%��i���(%�tM�,v�%n�x���|2+�>�;;���U1��:���7��_J"��7��ϳ~�rmvDh�T��S.��-�B^A,��,�mG�(������"�.{�#i���f`���T��=0<@�>�����%@������QR����?߇ӀĊ~�����V �	���uu���9ĉ�t"wF���`~~،�W7�Bv�;���J%����: Svg'��[�b�*��P}e�9-B�Jb��H�y]�m��^߾e�uc�@� �+�x)+��Gf��-N �����B:;���[��1fE����M��C���j�+"�ۏ
��۫oU�w3����Y��'���\=ujo
T��(3�F����h����%M� +&c7���oiky��Ք��)�����D��
ɪۣ0���-�Ռ��ӱW�:"�th��ՙ�2���rv���д]p7x3ʦ(�M�
�	��6N~z��%'!��R�;p5�vB��x��\�|���c���*d�H��m�g*��3��DUXkb�]��D�B(�I�2�JR�ϲˡ��� a����P#ΥL�}�ՠ�;|����T,�8��F~�Wډ_��P�˖�q�����޷.[��d(/��+}wT3�/��5����u+�<~[�4�&gL��OH,3X�HTMk)�VI؜���?�)js�8T9	]���n��TI�Y/G�6)�]�g����
��&����⽹��b{_��W��-N[�M���_TW���l�7�^��0e�#�
˙X�j���˺)R�B1��s�<i�@��k���C�>	�rzlݟ�g8�Ӟ��ʎ�����r}���� %$A��Ncٝ�������O0cq��} IKI���D�o������#�fF!/6D����Ƃz��^W�7	h�͕���Y:ie��T���,��7��Ϥ�e����I�! )ɔ����	n{��/�U6�>�}rV��{|D���$�����}Vl�8�Q�`��8
l�_��sAY���7�1�a���7��Ҏ ���4�k̴�͍m����&��3o7��ؼ{т�(����<'�2&zfG��$}1����+����b�͜�4S:�L�n�V��~l��Y�[�U��LVu���/l�������W8h=��K���CQxn~+p5A�D=��7��@��x��޵zz4wFJG���ip��APT|����ũ1j��%݄pe8���m�q�zE2���h/�ʦ�ni@�{V6Rj�H��J����%�6��E�͕-,�o��T������#.����
��-Z5%Ua�^O��
)I��uO�.,c�=��,S�y;�$�M�[��y2�������գ�gy�5ǻ���J�!�%�B�D������6C,�7xՐ�+���ĵ 8�.�NA�SI�m8~�F�^v�F�� рVWL�BZ�H%�ܡd�<�e����E$�-j/��bs@�̰��h��r
��A=$�Y���&��X���rRU��<��i��sR�	'��T5d�t��/ �L������.d��L��`��X���`;��!;�`_��h�:�l>h������X��-�JR4��+Ȅ��N���2�e�q2�\ �7����T�3}=���b*N
z�����@�E���DWj6���k��w�z=���+��.i
�-�4q{�)�3�2c��P,K^&�ȯ A2c���\pk;aӡCՆ�G-ht�$~�B���G.�"��)���D=��:�	����E���.P��^���&.X�I�e���a��m-���s�A��:�#�W��)�6h��Y�R���Ӑ�3��'��fm�y���D�3TO�'���HU9l��]ʏG��*�� �T�Q��ś=;�pWZ'Ur�ؙh�/��F !E�3�D�M�˧q�?j�"2�߳W���.�<bw*�8QwqڪS1Õ�e�����1+���$� �#��F�wsZGj��y	��ӓ4��:��⼂1��X��?����<��ʦ�v�E��G3>ȹd�O��Q2�r@^iF��*x�I>�V�ټz����o��(02�a��vN�	M��|47a�-��*�L�m���ǁ\Tj\��hxA����ZIa��mXL������;��i�.�*���
H㢧`o��2�:�;�ti[�O3'�_z�s�Rs�V'�hb��p��U�ɉw_}�w?�du�ԻO�.a��."�\��f|A~�1���d~��A+e� ��,d��I��C���e�%��'v�d�W7	�������G�|��,b�( �'�a���a/o��e�����x�Ѝ������$�<��)0o{�@�hS�yJf�e��.$-VHEт~�!�@
��m��-�p���~�]�U,��"���t�5�)�yȢč�W(9q�(I}�iy�L����I+��NƋ�e:�p�U�|��ƭ���ͶA+jur�GQ嶬�9�E�m�͌��@L$���ҷKz���	dw�e]�SR���8�<��a1�B������#�t�]wR�����A�r�m���>|�|۩;�i����(1{ϜL,����zQb E�:a�B-�Q�a/�ٺ�����50ɭ-� �RV�HȟB�Zo�v�S�s|���#����/�\4��~�I]Q��D���B���~���ɰb��"+�'�a��@��/�̖:r����
UO-�����n�������A�Z�d��dc N�=�\�鮮��s����-M�ַK���X�*
*dw��`�.� $,�Cy)�ևt��E�v����1�����g8��A ��S(Rv�d���%�U�%4�Y�9l���GOR#��:3�Q�)^���lp�܁�?!�.�W�?���W8I>QD�>���W '?�:nB�+#�7#`ڄH���\uW�����h����7-ПUf1Q��M'��Y��4�h��"H+�L������;�,����ϋHY�(����`��_���w�T��&�v�Nʾ�?��j"��L U����'Qn5|�هY� ����Ү�YJ�S6��o�i0ptR5e*���a��zO(c�tm���NK&37��bY���i��40��ط�q_�A����� �A���\̜;�����l�͇T�Y��)������0~TÀ#�⇎~� S?�J�W�a4?A�ߧ���j�G@E�S�y;@vd��6xDP3���ta͋��̱��3bk|s@;�qH{|�m.+u)�d�쒄?a�>ܖ�=��߱�M�
Je����H�A�%jF2/_Kq� �E�MՈFl �0̵�m��W���/��W��P�Rl��Z�����Q"ڮ��?C.DL���Y�Ջ��0Ar����+8��"�\�ߢ�L 2��8(۵?�.��(`�!c�2)���Ҩ�@�i�bT����I��#�,�)C27���JsC�Ɍr���H����VƸJd����tK�:���������TNsYkjF�Sվ���k�{��r��TW�<$��C��z��myNcd����Ɲ#V�@�Y��O�1r��Ox0�� J}%�\�b���ОW��{H �ky��u2��M?�Q���.����&��LXq��	�����Q�m0Xu����W}���PK�V)R�l��Z��XTQ���-\�L��m��$-���{� 꺋����˺�M|^��M�"Q�>Ub��YR)]���v���� e���f$�>]>�:'���8��� ~��|�j��*N%u��s�]�bKX�LK�9Wr���R���\�)IP��j��}������<D��ҽ��n�7��e9ϔ�o
����^�|�I�4��
����)��Φ��a!�J^1v����0����6rB�n,��Z��Ak�˝�.z��&�3$Y�B��
�O�.J��|�*h��yA��8�7Zs%0���U��ܲo�m��;ҍ��'�!OX�P����U+���;��i���T%g�hBi.�MV%��� ��TlR�o���
 7ӏ�}Q����ƌ�a��S��C`��u������mO��
�>�����œ��w��G�^I�FH��קO�r|T~٠?�~ � $�P#��"}|�s���	p7{��o+�E�bZcAT�e�U�}w�hY���׃O��rU�1�˃���QZ��r">��g�D���M���c��}B��H��!Q��<���<0�i���|Zf����Z$��#��!��/�n~�pBid�
C'}��OD�Dpx�z"�� tJ̊;�28}V�n�ƂR@���,��~�9U�j:��Sq]!ǅzp�q�i�����TB��7�ө�)Li�9�D�����(27e ���3��/g��E��Yk�گ���2����R�9{���dK���r��(̃�P�&�J$��@� �C"�*c{�#.�g.��-�Ĭq�����C��~�K�ħ�t��@5��v�*�#�a�`o�۲!��ߩom^&'�ۮ>`ؕ�����{oU9�)ːNfz���E���BB	�'�.���X�V|%:�;ox� � �@��~�M(~[�K��I�E�� ���&�W��V�-�8ũG�N�"1�E��O�����^u:z���_��zl���� �`�&�t�I�e����r� "D��p��a߽�^_Gi��]b �A~��j���{�� �6��Nt����J���N���t���$�|AQ�@� �gC�[s-�}*�'��͘C��+^3W�hA]�x�*y����sxR=�mx���q~3�r�T��+#����$��8�_vV�~5Yr�ݔ����ʾ�D��\Y���!��S��/�w��7j�kb0�ۭשO��j�W��]F���P���}Ք�-�k�r�d�v-5E����&
�5i.��H7�������H�$�29��?��d6��Y��tiLY�O�
��J��z�x�y[�2�(��ԚTq���r�;����4j�;�r5�"���V�D��� ���}T���6�26��xΡzL��T�O����"��ȥR�S���F�#��031Z�a��N���*�쿑c1������'?�P,�X"h{�P~Q�&\ޫ�7��3ٵ+�hSLד������'�dX{�ugi��%\�
�����/�����u�o�����(^H�	]I�\+�������$��O�5����hV��H��x�F�F[�;����/Ǔ/�r��2.��[�t�M+-"����g!�~{�Tƣ
�
��F�`[ѝl'0D�͉���r�M�����.�@r�K�1��� �BF�Aɻ�B����S��R%�č�*����MA�k5�T�4�b!A��8�w��B�S�²���÷b�
+���>	ߝ��{K��٠��&~PQ ғ�M̈C�z���M�ZՓ<'�vX�N2��� �BA
�Lޞ� ������D�\d8� 7��Y��<�lZ_s���!&̍��� ��'gN��G[��f��Lʸ5�gP�������m� WR�^��Q*"����\���.(8�_�+C�i��B�hFR$Rp����ɨ	}\�����д	�Wb?qbquФ5�2�b�\n'Xiu����b�xP���󡏞˓�9_�=aq��>i2�ײBh)����ԧ:;���h��:~������z�g��G�[UXxbfT�b'��3�tはϣ�[**mO���iL�����d��&�"`��oSK�KsX����h��w!�,oR�Z����ae��?A�]_!�(��OTs%����]�К�ab��늅T&k����*����T� ���_� ndb�"w6���1w����v.R^H]٦�O����~ߘ��s�e�;�=鱤�W��]���2
{�5�5�
m����=���:��`I��ס�]��{V��9�4{�*�[�v��!RJ:��5&���ܛkv@�ȗ��+�F��M�
��4��/Ӯ֯!�b�Pz���١�$��=�GeP��i�09�����G���ą:ش��[9�N��ĶZ���v�I�C�i�
����*݂���N՘��f�/E}��F��;�2]F/�
:"4xcG�,3�:KGx6s@��1������E�av�v�j�=yuTS��A�^���^P ��Fq�_���jYv�\�G�#�&<*�/������]�}N^5<��Ã�k"�f@�������6�!���>�����
�)�>�[�J�6����*S��0��ӷ�"�A���t�./�{ ��r����-�A���џ��t��:��M�b�4#,U�����R�@F�2��5��?u�����&�k3 �����^e�v�v,XI�y�"C�M&�D�f��Ѫi�G�*�y�����5�W@������)`�0����:a���<3�!�qC 0��%��*9��x�w�GY�B#�l���s�������S���7˷�D�>R!K0����9$�?�Qy�0�ƅF���#7�n�l�!���ׄ�^91���H�y��?Nn� j02O�S'7���G�����۔��	<�'Ղ�#��ΰN�q-��@^�u���\HW#����4>!�۳=���t[�T�UEsÄ�ƕ�3�6��QU�.0LX���ǐ�Cv�2r��W�P;Y��Q(�<�������(x�#�9L����T���\χ�FFY��,�N�:g	�ߘ��#~��r!��(:�1y���r�&F�+��?�w��=����l��Q����̯]�����J�z/	�њ���(��$��!f���G>O��7FvB�R���O�^�C¢�CP�y<#d	u9�vjM5�B��X6Pʏ����͊Wc�HPǨ���/�?7��H3�]Q���Zh���� aP�"F\����$0E3����L;2�M@P8�Ǌ��;�O�ԡ��L��A�\�v�z��K��*����p������������r�u��PD\�;h��0��x����������f�;־K4�e�����'�r��M�S�����+�ș���ÅT��Ђ�{��m]ӭ�����B����Yl�����Ƞ"��W[�0@��Ϥ\���亽�qb�����H���ޑ��)�s�9�ͅÐō��$��f�_^m�*�kN���ת�gi/x�(B�C��\�o8�U��<e���������b��y� );���VP'��4�}߅�\
yK��'���Pd_ 5ډۻv,3+}��C$0j�H����o��u�CP������r��f�J�F�����Q��AoA�����N���4���PurL��o4+o�Z�r`H�r`�L�k@���C6��	���[�eL�ĕ�i�Q=�,��ҀM8O {H"�K����.a2Y֍]��A@eV�_.������e�˭�A���%!�e�XcW1)]�<q{1�dl�kT�c��~�����	A̭��=��MxW����)��������v+�yZ�����3+,*ޓ2e*P/��]��z
k|vAW$�G^�~<�ui�r�7p�4>_�δ)��lCZ��nl?U.pS��m�o��W�*s��x��To�����L���*K2�rc&Ǖ�Ə��>�J
#Nt�4z��6p��5|L��Cy�9c�����It����xI�qY�y^�	)��)��<-^��2�l ��� .X���f[�(jx�hݕ|{*��k��O"�ae�9.���"2[���Θ�� jg�����C��:��=�?Ra���S�~�خ��Mh��>����zv�N�v�/;K���MR�&{�&���;�����ā+^ni4}��L�5��I��$]�4���k�l�J
:]�~\�ym���)���ҟ�P��a�J��C��L���e�Χ��`1F���&rߕ�Ŷ_����鵷�����5���,&2�F8OC��Ǜq@Č+�y�u���<����QI�8�,H����O�����qW�]Pex%�䵢K�Q�z�:(a�Xk�ȫ����T�
��N��X����(���VO�4�&3��{冴QV�M3>��- �1�T��E���*xyi�] �-=c'!w�Q,��Y�����6����/�	�cA��ӱ����[��d���!Ǵ֑H�(�l͕��lWK�K&F9�Drp��5������Q}��Lt�*~x����>�� �}=��Բ�2v��K���C�������4��s���o<#c����1%�����R���#g~����wA63����l���Xߪ��
t���s��?)KB9�fHnݔ8���AcW��$�;�i-��F��CŴh�ԭ4璧JBw�\¢�"Ǒ
0 �w_�2�tЬ��22"��fuf��ً����W
A�ۂ��o�@�+ ۻ�tl�sAb��࢏��j<��0՞Yq9�1������8H ��/�	�b�q�>�B��B�;�9ϞZ�������������(_�hטD�4^%�Van��bS��Ǖ�~eq���Ht��ɥD����-��oY�yO���N	@���A������M,�*2��"�|�gE73�`��t�֏VU�I<���X�P1������ט���qq���j�}�0q����3`����h�G�9A��buK.b%�.�ɑSO�D�|<E�+��2l��G�ײ����ޜ�A�WqC�b�I�T�/�)6��f�ܟ������x"|2�Q$V�߁�Now�H��y�}ڋ�Wv���p2��;��H@�jf��p ��������@6��2��0���kv��-bG�}��qB�����d�3J �"㼉��t�P��2P�u�;�௩��'��4��/91���z�U+�p��vAS�AR<��(�ߊy��%�E���`mi`�2S�v����fo�4�[V�)��O)�<��+U�%�Rq=;rƸQ2��S�}%y�/}��������E����1Ƽ��Zw�c:"�@�$���Tca��ˇ��
*a&I�p�EG�eyn~Ӽ�G}��0l��6�d��H1,�*F���@�QG�Be�[�� ��U��/KY�m���fz�� Ta��~L0���帅�2H^����������u��t2�xh�m�1\���Y�=�f�'����Hʂ���W�y�x�6'�l�0��*�`�	�����������Oډ���b�P�����χ��n{��_\��	�dV͊Y�>�kɡK'����8�+�G�d�aɼ�&��&f���7��O]oF#E0S�*)e�����إ�8܉C+��0!���p�����Q��m��]w)�8�����`��H֚�ן¥Oe�TZ��<�Jfu��6Y��NU�����[Eډ(�b�TI����m޽P{��=��y�]UƜz|=����%P!��K�L��2.�E�M�s�ð�iib�w}a98,�k'��H�4L���zR�,��'7_�����Av�i�������_��z١I�:�JqU �n���CD��Z��ʚh a����(��ta;Ŀ�}��[�
�Y��=�����k|�TޑTl���{�ĖI��������Kٌ5{�O��5qZE�]�R�L���ņ�.�tw�TЧg,��fy�\J�? 3lW�����h� ����`��m��.i��v$j.��ʿ��E�J�]R����{D���)i3��*���[6y�?I!|-7�'ۿ��5;�5���xIE�a�^2^s����!�u���+��������c�Կ�6��뛑���u,w$z{�3����6"_���!!9,;�1քf�es6��v,U]��tߋd�O8B�z��wCe`v��Iݚ���r#V,�/o�e:�����blm���jK�Ț�*���CIez�4�X���*�7ԕW$���P����҅�F������j`�@���7м�O���=���L�~d�j[�xW��U����Zh�����ݝ��kx8����QTд��D��+�.>і���0�n��Oag��`ɢ�&���f�ߴ�t2L�V7�F7��/`-�!�Xk&�K!�>x>����ޗt�V���F�X~�6�	4�n���H_ʍ�x�A�ݢ�rަ *Zl��T��Ẃ��M+�SQt����y���C|y5�ݫ��c�����ھ�1%�t����q�N�5ď�����o$Y�C+�} +