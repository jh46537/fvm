��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{MEi$ �:r������]	�������퟾�hfS6]�p��
� k4�[���i|-v���]���ڦN�_���8C�v����mΟ��xi$8du�CG�g�,��zg[W
���1Xw��/8⑫��O����QL�tp PE��մ̭.�~*�{ǌ{��?蒿G �s��TM��L5|�������t
$@��Z�����p����<-
+F�!��B�%���^v��炅9o~�7c���7B�W�W)s��po��V-�H1�,*Ǡ��OC�����s1�{���J9�(�O�@��H���ɑ���C�~��Z>�xU>��C�;�'����N�Խ��T�U�x�W�Q�'�6�-k�<�!M����N�V����ߙ�/�W�p=�+� E#�P��:����X@/�-�[����;$hF�����>�\�(e�4�;�������U�֍T���xzW�c��1������� #~�2�g��8���7I���;���L�����)`����MM��ѷ�wQ�Y7���E���H	�^�ʮ0O���Hp���7y�Q������r5�N��:� �3�~*J9L���@/O�V������"#����걥N��)å�GKG�I4�TͪC_�)RY��\@��#��.�ة�m��E5�WfBJ�9r���^�m�OvB�6;6�
x���E��p:"��+���@.^���1$W���!��w�p�Vpq�o��xck��|�;��,�y,.ĹC�Y��f#��Ǹ>v���]��Lnsg^���$���x���h4�Tf%����W��!����P���*+o�ԇv�c�����!2!�}K1��W��xyBq�3�yZ�,������N��o�8�uH�EO�`!�>Xs*�7��k.��{�����m�lr^dF���8e�ďF��L�&�?���wD��tQçT�hH�p&���ǀqRd�:gH�43�38�X����U��AAfMk�������@�Y� "+o�!��sT�#oM�L���SC^
�R���?�>�N�0 �E:�D��w�YA�G-A��Tyoy�jh���������X��h�qz9
�gp�	�v��Ħ�ѥ&�Ur7��䀼7
/�o�o�%�P���?1�Ŀ�|	��]0ZF��j�dսn
�ؒ�F�����FOYh�(��i�YS$d��֌V�|!�LlzTk=&']��� x�o.�%��.DQt	��.�zf8��U�7�Ө��A�k'*�����&��n�uc�g,�Jm��\��4��1��@cȋt�Ev'6��>�Yk~������dg��=�N����-��O��;73� �H\��b��3b\�y}j�D��/2��OV��n�!�h�!
|��;AZ�" ��8�]'?���77��D������>�Q��X�,ٺ�FƇW�������s\���q��<�k��b;!^H$3"c|��r��N����HMj����q+�ޚB�P!B�Բ�� �>�?�ng�ѭC%�ړ�\�����-l��I�|�����qDUV8��'}M�{�A�Z�䷗gڨHzPo���Y� �<���?RJ";�p�S�u�vE8"�7�2��f�E� w���xq��~���ڶ[���_�������ב�������,̌b2����SLd#W36������a�_��� �7�x�"�#�#:�"��-�F�È�H,g#�ڜ/7��#��z�,T��E��x$u?&���ºi;��4�pe�	�S�(8�߶S{L�'ZÑkE���\�fv"�=�rd���|Pz�����9�9&�t�^�7�BU�R��X�Y��9��v�Cϴ����G��j_o�~5���J����5��>Q���>c ������9`/}MzOcz��j�zvօ�a�jq��y=��$WK�}���ν�gs,p�U�x��2	�-AAT=�̓�S�8Zޢ5���_Y�xh��0wڳ�^������ώ�׫�D0���E�Ùy}v}�(�q�2�Z�������m)\��M�+���lZH�������1e{[}�*�[:Hh�"{Z�H�!Ǡb&�t:7C��LS�(:�Q~��쯹@�,�E�ivTسi>�9z��.���n9�	@�,b��|��W��t vM{��m�M��٩4M�2���]�-xO �y����FX#L-:�2f�^�������2��-}� !����pa	��5�4E��B�5/Ԣ'CHl�Kǃ��e��kq���3�1����r�^`&�f2�i��5ֶm�����R�!49�`,� aVH�*���)U@5�vo k����~�cY
[ֱ��.�̐]u�,#7��
|d���5������h ���FЯ�"xV��c=w]I��d��E�u��m=��v�>��P�#�(�7��=bH��躐�<D���9�������I{g��t�w@g6�_��tm���tK]���(�[�(�]�aY���N�0i�֎I1MIy�~��C+�2w�\*�P��L���0��8���Ͷ�~b���Q�<��uu��l����g�Kpf1w,�>�/=T�&��H7N��޻5�E�n5��N?�Xhx��c�����Y�@(d,Z"��E�`�W���wm��	��M�y�ފX��$.
�tp�D�_i��K�}{_����5ŭT��'G�d�,�m2��|��𾡺v�h�O���E��5&7�ɲI#�3@��"�3�З�EW�I9�/����� ����Ա