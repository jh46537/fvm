��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C��_�+��+��^���vZ�r�Ln��5��[��S�g��g�	O�R�����=h'K�H:���e�]���oF��Z9Ԛ���e� ���NL��տ���"�̒�miɥ��Zu����+�ۨ:��:: �\���"�u6��y���uϮ�;~EJ%�@C��n�T���Ҿ�s2�ɲm��Wvh(U��u7�Z�������!�?֮裫�p-} �l��"r*@�+����쉋 a�qB�Lw\��C=�ݽ�0�.����I�"�u}��h���a��^[,l����;J�}����~��+���1F�[08��p�G$.2_��ғ#�쥯2ϗ2�J�����L.s�~����*�D߲e��+���̝o~���֫ ���a�xׄ�o`��db���>���3�Z��)ig�w_���Ym�m��H�Y��.�v��w'r*�t�����ĺ�����⍠�2���,B��L����&�0��K�����ڎ�����-07�Jt��(��o{ s��m�:w�� ��z�8cvm$=�Tc:6јEEN�>�*]�G]�(j���
5��[�4yr5;�%$��&��ܪ<&Kd����g�WX�`��>,rI�>��#��i�\��,����+ ?ў:[P�t���q�&��%�� )~7JW�k�ct�� ��F��YM�c��g�
���k����$!������6kãtG/�����B��<"g��M��� T�츧�"��W[\b��q�����&s�Kp$#*�)���C2�;x5������=�1��+h���w"�� 9	G'���C����K>I��{0MZ�pD�<XtSj��T@ٓ~\������2��?�"u��}ݷ3��kD�8�tm�&���D��:���W���̈�����;;��Rb�]G2莈U6K�/�V����x�Ol���XXҍ� ��&��� ��` ���C?�M(��d�LY���b�)�V
��Uz��usQ�ѩ���qlVdO��g\��hW�,�;c�p�������R�N�#�6��r���ĽuV��_[C/L9�a)>���������b���^yl̶�p2*�K�&�fL07��Ʀ�uN���J��7�"9$�T	k���D�gp��yė�(������F����)|��`�ӹM"�ٺ��t~���� dӴ�_
��JA�PH,GIt��X� �.�|���,[�7nI��� � xg��H����U� �x��揧(�H+:������!�%wR�+�U¾�f�d�X�É�5������&��~=�$N��-\���LR�,E:V����@h倷��y�W,]Q��ȞgF�׻eT�8�|�8���c��v6];��{��c����+&T+�ެ��5��#9�­����C�`k �;�X]�f ��KPQXW�>^4dܣ�����<Fv��)Zl^	cR�gƵIM҄�鮴q��5/E��R�3��꾢sÈ���B�����wq��� <���wR��'����ȵ�v�@G���.�J�{��\"4C1���&�x��%֌Z`�F+j�a�O��	���LLWA��'��.�5����k>b��}���ʔ�X"S�\�s:�uM�$�^��;'Ū����0�����g���w ����xz���ם�ިǂ.E����nqd:�%
	C�n�2����4%���X�	��y��㏧iy�=��1&�t�F� ���hT��IJ�"�Lԁ�t�ӡ�����T��j�&'�4l18�o���~���4��o��qOZ��2��d'{��Ը�����:�K0���|F͍�C�^bΌ��D3�[���ۅ-{ȓDSl�� �;C}�p�8R���t~%�I#�z����TU'n���y���L`���[q�'4���g�u�>-�t�DARa��d�tKo��=�+zKZn��BK�@�7D|W���q/4�9羼K*WLU�l�iQ3�a�)�Irg���f1ͅB�6��^������%]��tW������
%�ד �����mLp�R��~��L��J;UC��وl��5@����J�f���Q��F��*�h�LO����#@��u�^y�SAC�� s�YT��ܡ��(t��t7W[���6@�M�t�j���T!W�I����Ӛ��°�^������/�=ϢcK���+lm�d�m�6n�0�C�g�%R�Uf���n�n
~���?��NUk��؏��zT�H���"�"����*�Ȥ���D�W�	ʑ���p;u(�&4A�܍ �r�\�N"kιm�#�А�nJx�KT�FRnv�]��C
�����^_�S�c6	z��{u9�o\�"//Ԏ�d�d�%�ؼ�)��r)"�C2�D��څ�H�������ƫ7�q��(���}��{�,�G�k�W�Ч,I�����3�V�!O�\��F�G�ȳ�c����U�,�~%!�Z��]:��N��ŝ��$8�)rN#���%�E��I���%��{�Z^O#���)��;�R�/�1G��,K��`���qS�XeZ�X�{���:+��&$�P����c���a*Xf�yW-���h?�+���Bml�_^8@��O_��w/x=o/o�M�wQ�ڻm�Ăw)<�}"��X�lڳM�'ԁ�٭�Ū�\9��?��퍮�#�p&&�,�š��'=��#�T��ҝ���_��Q�������I�39i���o�euP�A�퀞�0R�����.X=$�9F���0ʻ(h�歲>��k�� u������D�i�l�����u#�"��r�H,�Z��#ϓ��6�K��y,y4Em#j�d�١)��GW��0$�6rl'�C4�5�R�T�3��0ג��A��1����
�<	�;xUf�G.������|ym��b�p6��{rՀ�[ǖ7�GKxs�- T3 ��_`�W��Z��)���,At]A�� ��3�+.����R�w9������J����	T7�O�dU(� >qq.�õӌy� /� r�bgC�2'������z�>դV���@%��}�6��Ҵ`�
�|����U�ox���������˱�#��:~�={"�'�]�����ع���I�Օ|ê���C˅�u�e}!��L�1���.FwטfN���}���x[����įD��R�Ź;�� �I]_C|lm��,+W\=�_�8�����
�� lhEj�*���D�u޿3O��@f�����?|(%dfDX5��i2GϺ#󶎬����oE��Q��Zr�A�l ��;5l���a�s��|sy���j�����T�c�A�%�ѭ��p_�̵W"F����؉��+1�@�l'W����cx ��q�*Kc��C�O�,\�9�XX+,<A��O�11֦�����A��R�i��ܴB\q�CYT���I�����?����7�:A��t	JŨ��Zە[�?]~O�{��7����OϾ�e�(D���& ��1J�}������F�TȓQ�,!Z0Ͳ��E�KA�M�rE?��o�"?l����v>35N̓�3���z���~@����m�6��)����j��QLVȝ	�ϼT6��U�T�b��Ap#P�(t��=�}�1\��gv�.3t���׊ir���>婫L�_Nrx��g���c�"����x%�Dx���2�������!̈́<i��;��U��$R;���X�����@��p� xNe������I�^����"�;�Jݣjz>�8u����-�7�r�	?��c;��[OL5n�cX��At��p,���I�
�M`e����D��i`;�"��Kd�#���R�rU�nA�.Ё�'[*�y:�A#�E=I��TU�R��O�Gi��5�:zȠ�*�9h�K��زդG��,����S�4���0ə�<�A�\-�������{���[-�'��� *m��+���_��`O8o���|9@�H\�jX{��AeLћ��`}*�]�3��=cM�����%~���2z���?B8��:�48(��ayv+�-�(�>t��Ck�k��>�g�BW܉�����>��|���hmN	����&y��g�Y�ʔ�����f�ȿ���<V��q��fA�1���|"<!�s����E�xG�d���K=�{#��i[�����}�I����^�哦�O��(���`,I+�}��Ps�C��@�[s�ԱP?�D�}J�8WQ��G'�`L�<#�*�}G�R$�E=��(\�h���u�h�5�*w�g�k�%hg�R>�p�t��;f���36��\�k��, ��}�G���z�"�OP�QX�u�9�X�E���Mѽ���,�d�/�&�tq����r�[ %���	�TF{b�'��Q�}��i?������m�8�����uV��3��~X�.�,����&t]�c!�@"�'�p�k Zr��q�V^��Vת^Z���t͝�l�
��4 77�W,� J�j+�X�0o_�0��>��%D�ҥ����j��a�_�~c|5#���/��A����N梶�����:�N��R!�_�*����3@�ﴕHe!Dn9[�P���L��D������lfы?�N���`S�oL���yx��/�)i�/	�����C�xt�_w�/.������-�Ա�1$Px���(6U��X~kuQ!��U�I�NWͫ-L!�2눕�;���e�!�sP������:�y瀹��-P���~I����.��_��58M�d����K���B�x`�[�l���ΦW��z�����%�,A�R�*��QqЙ>��I+/;CU!?߶8?5��Y\�WJ��o�9b#wSv����V�M-M�u��F�hg4ǭ[ �씯���b�r�1�9��XW��|_]&騗P���.U�����x�ו���n�����ƙ�ixB8�{Vyo�SN�dӰ��*P
�2uk�y���l��R�wP��q�2>�/h�O@���7W��(L�ˍ^��U<IA���;�R�G��4@�J�m��g����+�j}���j�s&�_�iƙ@�����[�$	�s��8M�x���Y�/T��|�,���eٱ˩:��13D�;ںNӏ� �� ���g��x-��se:<�ѥ��~d�әK:���m�?$}X�\-W�`����AG��)d@m��+@0����3���n&�>�84�l�k]�sBG��"�ހ �(�Hq��4�R"n@9;��
 �W/Y��Z�D�w=�S,��+��}"7�J7������x��+�R���&�v���Y4�jo��M�`��������� ����vwA���,�A�� Յ8�����̳t�l��i�8��`f�	%�NS�tG����!�t�Ɲ­���x�Ο�~�.�>�抲3�;,�>O������ ��`x�$���9�Z���Ňl�ꖏ#hu�F[A�0�?X�4|H�E�ݷ��k�+U��=���T��&���¦��N��]�G
���l����s9^N�6����8�m������.�W��LP�m�3g�+J�[f&�a �Gч��C���t����!��V�@"�ŷ��
{���`���b�#��S0
y���M�0W,����}������|g�<�H�:X/'Fg�!|Mk�2�-�������G\�O��oI.�Mj�����k�Hs:O+Ύ�X��x����
�Ӈ�T���u)4غ�)b��YM�خ���W��+a�gxN[��a8��%�M["�*?_����N�)�1���q��%���-E�S��=�Ka�r����̃�����f��'����gZ�W{*�SX��Q�ZwzN;p&\/�H�FE��x�X�����.S��s1���V�f��">����(�(�ҧ�}.��$Ю�\�)�^���A�~�&7�L�1���7����L�N�s����8e�8��U(�)RӼ�[���7����YM-�S�QE��AdR�{װ�^"*5�/�	
��O̵Nu�/Hi�%mrK��Ɇ��L��.D&�J%�u܋Dd���h�瘱��*)�6����89�i@|u F��ħź���6��!+�����Z}tr�n�.�;|�Kw$�r�y���t�#5PE���d�����F�	��i�pP����D���\�u��Z��^"��)+��~"s�p�i�1�c^��2%&[6Ȕ�F������W
������	�$��F�u�E�p�q8v�r3�W+�Ci��p`6�����xt�R9޿=����1a���du�&�k�B�<QsĽ�&&sU�vO\�Fxu�G�Lր�Uy.]���qr��>�C,��t����z��sSVm�S`C��Týj��EN�!���O�䗇Q�72�۱�Q��j����5}��H��ȭ�\ʍ�_:��to�\������2A-�M�$��$M,��9��"n �����L�4қ��*�`X�f�8� y�^枴K&�;��P���#�|��ɂK�V�=��cu<�4�ث���3��<&Q*ס��-_íW�c}�~�� ���u��¶�u%��U(e'Z��j��\�߯�2K3��!�y�p��`k%`�G� L����	u��Z�35[TU5��9�0��-iw3/3y����y����@[g���"V;��P2e|4�����8����1�)�;�p[����(��]}���n����#Ϯ@��0�CԜ���� �#@�p��$�cB��a.�;�x�1����Υ#��OS��4����8�J�[e'��#�&�T�Opg��*�y�p�P�yH�[m�q;2�/�z6�S*�J_���k��v�A�E!��X�Y�"E)m{"!X[��6%���Ez�4"O��k 0f�����'�tĉ���I���}���C"���*�	�7�RIW��m�ه�3~�##L�\�WO����
��>�����Υָ,�N;�Ҕ��(����}�8�vȂ^!"\�PBh�/j5C�d�p*SW��?ȸ���q�|8(�[3�4��72�IV�Y�� �;��Bt)�=Ck�^����|'dI[�H���#�ڎ��|��� r90ϼťP�op��ۋs7	�/�9*�\�J���1_߯�Di�p�C\��9{����9�UU�}�5{+�o�6eo���(��%����vm��ti���]����w�������H�T ����Wő�;��Y��A��ʇ�$d������R�@�X��#�y;�Р�<��B�9�h��]������G{�(�u�i4�C��q�m�ҋ���2*LF�pv��\����D+��{4���z�� �!Z�����s���/~� rO�-����=8�Mw�vǤ��v>�"#��-�[��shUgZ�#�����q�?> �eo����e�(���I�0��f�g���i����u�q��g�X�Ow���gFp��3�t���k��[�$��2=B�z���j�2��t>��"+fζ��>̟��W�2�gT��]8���ߗ��%���ѩy���ޮxH/����w�?b��+�1
	��@99:Z�� 6��e���r]���|�)dk/�g��Sׂ�0T��)tm{_n�a΀��"�nV&����$Rd�b�D(j4����l�eW��R}�)Z��Y�Q�cy��p���f�,�GW�:s9þ9c[�p����}Ut�B]��af�d ��f�_Ld��9��!Fs����pɥ�֤�Ӗ��(J|�Fw���X#^��L��SR����NRp��:�fH�b(���l��W���)i�m�:���|?��u&'Y� (B-`D���ǘ������e��ˡ�Q
�""��@>�F�hV��6CΥ�:��x��A�%p U�t����χ#i�f*9P�7H?*M�}�T$�
Ol�7a�K;,�]_E���K 8Q���O�76١��5����b}�jJW����T|�w⒎C�b$t�M�G����uv�Ds�2�)[�<=F�f��(�o^W�*	L���ʾ�<���hTS�bat%�����X��ŋ�� �E>�Y`���z(���zA��û֍���A.qW/�����2�mG�vF.	y��"�r�N����go����0�H���HbT��Y̺.<"o�!k����;:�����=�髨Ji�&��ѷ>�
C�I�)(q��[Ƈ�-�T�B]Q@�馲wJ�C�5Wv�V�%=It
G�qV��Э���7�P?��d�A��v�W�\�����2-16� ����u*�FCt�ϳ�Bg��Ν/q��Λ=���'@�S�LmD���V\�M�5��7o4�׽÷�Tү,�^�L�"���2������/�����)L��mGKg1%�����ƻ\��:�v���P�]���
>��3�B������������*l�1�Mh�	H&�(bT;���o�9]�6T��àhX��>�t|��&e��0�k�y�q�`Zd�D-�%>W�o����̛M�2��C�Q�����b�ك����L�]��+��i�j��o��f�P�'����5�h���ao�aT�6;�U,V������r���W���w�O�V��GE����K(S�R��L�Lݣ���j�Lm<�M3������U�P��vLNm�-�JL�zP�?��r����-�R�雅��_`��|�uշ-��kj���pb��{;mq��:=G��(r!�\�U\��0��B5i�l�������&"�څ�Q�0�r��5�+EJ�WP	[	�/�BE'ex�R�3�0'E��p
���lL$��S�RÅ����tH��M��"�16ſ �HLz�p��b`�Z���1_&��h�T)<��SQ���Z�M��;�x���� ����式<�Kq�?Y�����m��Hl���)�W�TJ����V�g�C���O���{�\�F��M$�b�"�4��t�}���z!Za�t")�}vB D;��L��u���r��5mb�#��$&�){��F���Y�`-��w�K�=�3R�CYB�pe�����Mߺ�KE��U��Z��������y���r�T������f�J�_8kӑ�{ �Ɇ�}�!���+����j:�K�,���]�"�@'(A��p�l�eY�FA�]va���$�fA�W��8�dU?������$O1�cE-�CБ�-���6�0!簞��9ju���%aPZp�k�ж��d�kr s�ܹ�pYu�;)���m�������eg����0Ϫ�vX�s�.�b����c�<Ο�\Lǋ*޺�e�u5�R���JHN	B>�'gHJ�����P��_%��5���tHօ�X����˗hWZ�_l����%/!�!.��C�膃����s�މ*y�����?q_�O/?�7g�S�椒�K'I��!+ ����˦��aޤ���;a�fF�������W��p��%r���8=�D���J;�,Cd�zد叢���w�����iDWN�8F��%�%�I=�zE�5a* d��~��+;1O&�k6/��͒H�%O�J�~���Ic���G���]��n�4��G�L-	�̜
��E
ņ�}x���.\�v��-+<��'&��хd𠪿4��Ĉ7�4��Ŭ}%j�xA���8m���b�]5�d�6���K��Zm��2���Fz6����
���ˈ��A�����a���Ƌ��-����m�F���j���G�x���Ԉ2��$=��5D���F�n_�>�ܑW��T|d�:/��[�=F#�ݟ� %<��(���W�/T��Bt�U+��`9�^T����@)��~\^�����|���n_s
v(��R�F=��I�����5��Y��qi��B���E�碛O�_bJ��W�4�	a��V�B���r����)���v��f�V�>�ף��x\;�:��~�;���e��]�3a�=�-����X��ao�e��F�U{����a��5}��u�s|�X�IaNh4�M~F���9�����g���rh�Z��T��g!�HB3�*��R�m��D���4�=��<Q�ꙋ�����$$��Ë���rmV� ��� r`Hy`��!F��m�|�Ep��4*"�- �8m�����^�s�����Wf�*1�.�wVn1��]_����ji
vaH��β��hB���HF���6m*m�Py��T��sn<eA3\ȯ�i�����C��Z������`k�?��$z6d(j4s�LwjXb���)������{�U56w���$�m��L��/��v>u�{�(r�8�S�R9K�1�k���@�0�����:������]E�����;��m��A=����Q0���B;�G���OYy�pX^���fK\݋-�9�/�|@��V�L0B�)���a[�y�ߝ aTt�|��ic˅_���s�9Y�ԋ���F�rev��@��*g��*e���-��?�Q]�Nv�.(���⥭8��mZo��81�d���0m�^���?FvP(S{���k6&����r��&��$0��}?W[
8c��Y�N�����8�5��p!��+���?y�eG܎�?V�	��U23n6m �,�(`!�7���CCC�/�ζ
ZJ ohWF�ף��P1OI�v&��I��lR����:N{��"V�O:�]q�	#���$��'x����v)�}��M������D9��T��TJ'�&��[n�z��e<����:�aF�\������v�D�:�x�#�T �9�Wo�԰�w�6�i�($��#�N�%��-^6���H�&~,9uW���roz<!)E>�R�Xx���&la�ʕ ����k>}[%!�l����մ[���ko/=U9C�N�ó���J@b�t���g½��t=�K��r�7w<��;��_��4��@~*I�(�̄��c�ç`�1�gS�ŕ��,�95��;šv��h;	o@�#jb�:�薗[����#�5��h{�͆_�w�zH��/o�KeGp���H���Wd�L��<���T�e�F��z�n�|Ŝ��]2��+�o�P�5�~��h��|:)��v�Y��v����X1 �a:�z�`�BI�+v��r1$��K�4��>IL���O�O��m�!pNy;�k�Ɩs�������Ԝ��rPoi(-?��[V��A���LJh�5h�;puO]0Ɔ���x��R�.�~�LN� k�H|�B��d,jTŪn��bukǆX�B�w���įt�q,(� ��