��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb&�L�S��O�e�m��R��4d|�}�si��S�!xx�UFMD��u/�Ef���p�V��C�:�k<�#��I��`*򆺐[о���)�l���c�Y�z�H���s�#~��ȿ���
���]y&A�f"���N�HL0'ө������-�y����� ĭN���>y-H�a�`��Q8�.��ۈ]`��ޜ��#���9�\��l�IYO!!�� �Y��P��Q��XIkLjБ����[�{�+��\4�{
	�:1v����-Re;|_�p�R^�k]�K��_�!%4xu�0$þGtuO'gݥp�_�!��*�Ŏ�^��*��)
����YO���CW�w0�߃f�,v��;V�si�	���7�qf�/�g&��d�%�tR�4Sx��?�Zp�#~u1�k�Pq�m-P?�S���N�'c�+�4�>�,A��=A�e�3[*�7 �o ���E;��zpGl+N֬\���ل�O[
�"[K����'s0a���}�YMWIUh�p�J"R���e&�n������d�_I�>����`�[�o�)T�G+_�	ۡyu#>��|�M�-�:Ϸsm��8{��f&��fn�b,���,����
#���4�����'(	� <嚜��)%�����(B�����Ϗ�TuM;+��;W��a�A6�h�ga�[);t��Zo�%�<L�������b|oP�D�@��*����:z����#�Ĺ�	5x��ce�n1F�^�Y�I�I���߻���r����bă�}�>�^���/��I�^4k���̋������op;�#������5���¾rn��ͅ�WIHf[(͌���ˎQ�=i]iO��7���B���Oku��K(Y�Y�E�T��$��q�E��N��օ H������e5�2.�����6肛� R`���+��<�!h�š(&�w/^�b���`�`��2�F�8+钟%N6�D��f.����q�zg0�F��t�O����0�Ԧ�ب��,yX��~���0�/����z�yJ�(H�� g�sc{���d���������E�"�V:��$z)�[]�-������u	��aW�:�d"DV��({�����Q��UO<��U��N��M��=A�D
�ۯ����|�#�1�Ō��c��}ϢA���i�����u����V�6��3���
P���h5vS�,�B�n���b�qU��+v�k�dE��Z�3I��+(3�9|�QM�NU\�b�wn�2H� ��&��"��@����S�=�=ϓ�,z���}:�{7{hA�o�k�
vE���v�<�`-HR�����=_�5��94�$4ý��~�-vj�K����})-_��N�%��0��)H1��"�j	�k�&!a�S��bD�n6�Wb��p�6�M޲s<�Ê��:�h,	
��������z��%9���H��q�w��Z�yޒHo�ԾlZ"b�2��4�
l��P�O"k8��DE��bw#Z��,�3b�K�$���k�(�8�DY#ܵy���!������jL�,V&���C��V�# BTp-�^�*n���o�\oNJ��>J�[�`��q��I})���ag�_�7�ͮG�>NT|w��ؠ:��MPк��?G���U�u����q���v[��!�O���/Yۨ?�Ꝩh|}d�C��8V����;�fN�HB6�M �ƅ����	�z�Ý|q]����X��	j-I�7s�y�R��@+��r�yUH�0ؖ��t�Kn[r4��GR^e����t�c��j�n�%E�8�9u��ew��d�.|�3�����}Y�:�`�oe`��0�6�:���Wr���gjq/PT�b
����j5���� NA.���X��M�r�Y�4�+&.� �����ť�\k{�	>���g�Gp�h�sri �ݙ(��߉az�rT���d�%Ӯ1x�������!��+P���G8�6t�7�u��N��4��70�njv��w��{�N3K4t�8~de��[9����n�M3�B-��U`�����(���M!4�՟�/EvS��2U,[�j4:k_���W�����%܅�	�^Q��c�K�[�حϬ�`_gW -r�|�{M,�2�@�q�X�({�n�6��� Պ�p�0
�r��� ����;G1�vH��ے��f��C�Y����y�"��d$���