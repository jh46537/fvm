��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9��m������G|S7���X� b�=Z�Q�WR��-��+�q�5I�kh�7��y|x�Ev�}5餀Xs����c<FVyԊ0�g�M�8����.�t=��������,r��6�����1���PW���-�:��s�C���d-Jx��꒞|<����@naY� I~��;ÀlFc�Q��N�}�č���ێ���?�[�|���ae�f�[XĂ5ޛJ�]{mff��V�l����h,�ZG��,��%���E'�5eF�>�!%�kTnhB��o��6���4i��W.L��"���OY�����[mh�YK�Q̷��WF[5���f��>�ՠ��1]c�2|_���q����v��I���XN9D�ڿ�A��_.�1���rP�b�Ј_�A:?,�<"0^��X�^=;.�����N��(`���_�ECga��?���>���1���E�9L��0b����&���٠��⪴6<��/�����i�%�Ix6��4D�Ȼ���W<bg����jH����ϴ�n�e�W�-��q@Fd�U����c��s��v?��I�@��;�΋��i����(�?�C v:��X�)�Q�ѝ��:��i�����Gy�����]8F@����?%9�B5����r�p��C�p	k�E�=am���D�\��׹&IL��N _N8w��|���f�˖�'!/ѧ�i��R?�%i������<��`��K�d�߳��i�%w�h�=��o&��z��Dhd��v9|8Τ��*���g�x�+r��� v�mR^+Ezt�(%�ռM�'n�K�\RCx��hTơ,��l����G�hP����� �w4�eh,JA��x��{��:��2Ɏ?=0A��%1�lѩv�#�9��k_�:��U�Ҫ6�|��z&����ԅe
s�[��@��NՙdG�/��2��6OR���B!v���2�d��Dq�Jt��
����&���I�A*OQ�X�1X~v><�jEqFV�̽��-]�j����	�!�o8�a�`����DX��5(e)߱Ԭ��\"�#fT��ҭ�� 
���2mN8㳮�j�Y:
:[�E۩7r�?��\�L"�o�µ�\sک�e�#.������B4u	g��ƨ���kh��=�e��k*As�"ϏidCʫ��Y׽=U���?����o;���µ�ěf҆#�`�%W�6Ȃп��]�y�<�%�QN{�wm� �Q�!��y�i�!�zI�:"�$��0�Ӭ<1i�
e��}peY���Y])�CR)E�F&�G��׼�)8�[F=h�vy^v@lVae�eO�c�I,?�HH��)o{]�,�'��ʏt��~c��)���cR>h�?U���R����0c��g,c��&r5
 }#D1���HS�NHeן�n�E
4�4�9Or�n���)7ʇ=L���٤����"�5�io�f�Mkа��T�d>�����v�B!�Sh�VE��W�=�	U���V�Flm����;�G�1�W�s�ʸI%֊�n�EhL�d�ō�r�r��`l��EDaJ?rZ�G3�C���O��T�d���B'�6��x�K��gGj�qI�3BGn]�71��`��!th0-_\�-�Ub�}�����&�}!�2��>��:��9�,��8�2޵Q�si�O5�?�V�;�^V��*� ּ�[�{�V����D���	Qjfd�(��t5�&��Ǿ����?��A�X��ӎ�c�d&���C���O1�s���ep�h� ��Z+S�% $3�@����R���,��2�g(����=f�}w�����Ԧ��b��b�S�wY�b� �
��T�Ck�9�ʷb���7��Hj��zSL|N�� 9�u�P�q�8W�ΔS�� ���E��̲M��aZ�3��͈a٢6ر��XDG�$X��	߀S�:>Џ}6�45�[4��<�S	��IR-O��d��N7��^���kϰ�VF��q�b���O��c^����%�3ZK,�����]�}�r� ��� ��N��d�����塤9#G�` 2 ���ܭ�p1N��;>i���Sf:�j�@ы� �GvC<q<|��ʕHq� s�<}��;$���� In��"Oj�fݔZ	�F� <��y ۃ����$=��D�.�����u��K�� 1��F7�	��K?���.p�\�V\ޥM�b��^�\� gThR�Tg��S��x9�9�!��+��Q��nv���]ы��O;]	�U�3�?"����T.v�U�617���+����J|��h�m�a���m���=g1�`kٵ�a�-��<ʁ��y�%s�9��@}fP�`��n;e��l��{�%)��U)�ɭF�F�Λ7rx�˧
��1�J���z3�r6Pv�0�.b�f)#��5���[����I7���O���z=ƴj{~;��((*U��W��5��jxK�`Qɶ.TJ] �� ^q
#������w�g7��]��
�_��"���bW�c��Q�5HߝC�߯�]���|�bhkV��-\cB�ߟ�j��3��rw�����i��1jg�7�
%g�,,�7ڛPVn���"�>���,*a$Qn�׹����P��J���M|�ʍ"^6�)^d��ӛ@�6R�co[�T���f�4Xg�y��b��+x4��Es)Kzo�5�ɼ�â՞�Q٣��&��T��^���_��P�z�y�w��6 �mik�s�]�B	ڹ�\-$��u|0>#{�[��jr"b�{�l�'������j:;��Y@�s
.�yW��� $T?[� �L8s���b��=�@��(�E��+!��XFǳH����W�~M��b3�c��V�&�DMw�Ӛ��t\aUK�<k;)��8R�sm]d��yM����Kn����oI|X9�E =}�B�B�O���}ڸ���H�t��Mu�X�-8�N�	����,r{M�i˳��[X���~s`X\/#K���Y�i����V��I�֟��&8ceF8���B���� b�~M����VZ�S�^@Z(� ǙI{�xBQ���o�°y��z0����e�Ǉ���}v͌���-S߂��غ\�d�M�4G��.��'e�6��V�����aJ���4���(�hZ�wJ��^]��4,�*~1�K�=��Ֆ�b@	)��Ϯs5#jz�I���[���P"�-�� �)�A)���j��g��U�
�ƀ[�(+Ϟ�a�Rg㱊Ͷur�������^+��q��8��/�r��p2� �"���E�,h/�tz�U���bODO����������|��Z+�f�4�8�iA	�Ăo��?h?�6�Uv����jjH�Ï�}iȰ�L5�pf�=���R1WS� ٭7��n�˸:�4_˜������[.z���RԛQ�_�������qp�މ���ǸJ9#:����X��<K�dp�N̕�"Y�d�}�c���L�p�S�e;�֫����;�^�Sd�tN8�;���=6��.�	H���I�U�N��D4�Ö�}��u6w�K]̽ud�U��6ר�B�^�XnNb�k�5����/k��O��h��ǔ�x,xA����QR��e�k-"��~ �q�BK�T$�S�%V�cB�r=C��c.��*�t��[���M~7Yw�p�#NG&���<�C�~�����sQ��?�r�&��黲ؐ�-��Ad���L�0���m��eҢHI����ye�d�oIu$�)d���E��Y��;�N�OE<&+��wV���{
����7tY��3��H������$
�� �
���ZM��+{���xK�zz���B�Tɷ/�@;N�6f��ߞ�Ts�`u0���JqQ�? Ȉ�\b�1ZW/�U ���ԧ�ZuK���x^M+%\5 ����k�l��#��w����xb�y�o�##���#�+4���m���`� �GP0P�0R��U +#��@
y|7���D�����Ɨ:p��+����@�	����p���~�ʲ���P�����?�+}Ք�f��b5��}��3�tp۰ǩ���#�o�`���<V���e����8#���ϊq(����\?��뫦�j��z���?����u�f��	��^+������9������3g��8��.�`����+�(Hu%]l�st$�2��"�/��p\�ͯ����D�W�.�l��6�G���a��ƅZk��*h���1���	��P�[�n����/e7٣����s�&�h\PJL��=?=Ƿ:�������e����i�����({j]�L�t�#��X,/M�� ��l���c�0�D�u��4O�{ӎ(5�e';`���	��݇?�[�q��d=f]7S�jV;޳r�O�k�0��h�DqJИ|��K�ըj�,�(M@ß����F����{�JŊ�y��_���*q�#�=�)�����g�|h��܋/�
+8b�=���a�����Y�Lt.�0��X<���[�eM��3����(�7KQ���n�J� }�����ְ�ƾ���k�08D��f123d�~GЛa�>p�(;��`;x26Ԭ
:��U`���]
�L��k�pylxg(�VU�$�Z��q�ز�ˍ�g�b�$,�~�^�L�������-%s�6h�l����)������ݫz��%��Z��u����jsmu�Wu	�&�L���-; ��;�?$��<L"=�wx\U���?�?��B��n�8��
����t��p(1�u
�1�j�4.����6ڎ�g`���P�h��9��Eظم�(�p�+�QO{��MRh��E�/�i;�!�^�Q���a�ƒB�=�cs�|1�����q�א�<�F������Ap�<���pr@;��U��Mzy�*��;��_KX�T��Amb�\V6�0�DK�`2�}^�f�2O�p{�Xy��#OSU�i�*^���F����>H�N��M7�I�syЃHG���6�������Rh�E���<J��њ�W�CV�g��h��>��	�����+a)D!�ve�F��*���_j���B��``Ϝ^ ax+ć.�|ƚ�uw�PtC
�d�%�V�g@�Ap���3�i�H�9�g��.�A�2�0F�}�8'��,$����M�; �Q��I�A�n2����GM�:��A��٥�ؑ�Q�͠�r><圠G#ͤEo��