��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���a�%�sK��h���/a�y���v��=��w�����:�y$f�*,�RA\��S����ћW;�U���T�Ǔ�q�0`�eѓ^����8YU?to�Pb�I�����9���������:����l	�~�Y���)���L8�|m[P��Z�ј�79Ӄ���e<���_�����^�2�����
v��;�{a�<Vx3�-�����ٍ��/�[�mg������o2����@�m�e�?ኂ��l:g(Ozl8S
�-�CW�gF�5�դ����>��'K�:���ϵA��8�l��X�0S����b&�7�%)����!�h/Sq�㾴.��"��w[�Xe2�.ƿm�?�g0ۉ.�*9D��>[ˬ�?]#��m�g+��;��Lb�W%��"�����n�F�`��VW��th��Y*�1 ��a�|�!D�+�iN��,����p:
>�qC�Y2+�0q[<)�����;^�c��E����6�A6�\d� u���T�j���qM��������?�``�����[�G3w3���Ie�OE�̎U���|f'�v��^�ɢ�Ԓ@q� ��bV���F��5���%��<�2�d}f�������ڱ��)��(N�)=��<� �i��<�t7����b���Ԫm�i�b���x��]%���شu;[vz��r^%s7���k^�h�4��es�k��T���?΅����+-5d�BK��䇆Y�zsME\���)����������V6Et}̯�\�Jp�<L2�q��=�'���^.?��Wo:�f�<gf�����{�l�^�1*f3�y%X��_�4Q*i=��,ZI�C�M.$q}VȀ��x�R�ϙ����H#�k+H�%z�7�1kX�(�]���ʸ�C�O�y=?�Dv@�dz&!��H�K>2�Q�Քh�S���<�`�����wȟ�~���ׄ)�s��z�q�~Z��D4י�����K�5/p��+����swv��ܲ���ޜ��9���Hkgި^�A�d ��C�eS�k�
KY�v��^��Ǩ�� >�y��E�v_���AT=�X�]YQ�`[Xn��Ż��},k�c�Z��X��"��%�����p/Ҋ�z�*�KӲ�_���0Ҋ�%��?M��X�-c2�n�d�48'����c��n�ز��� �g�N]���Z�l�̓�$��wK�X�\N//ϋV�PXOE�?W\��d�	������ˇ;����	� �V�ԏ�#dˠ�ߑ\��d >[�����v����7p�ֳ�u2�B�F�F�¾�w��Ȍ�8�t��Ѥ
�����s��Mt������O���]RG�Q��WD�
R�F���ؚ���b�t)�&��-ӻ��>��!xt>Ls�\��3��Xۣ�G^|R�S��J�7ol��(����u�*���eEj��ꕫuE�MJ��Q|����2�\�М�d�0/}A��)\섞��r:֦���V���S#�7C6��ͣ��/h��gO��V�X͹+J ���{)"��|�\j(X㗤��!/k��`�^�&�l4Ӊ/[�Pa�� axW��/�)ۋ��¥�X�k4��X�ͦ�}�6�u�e�v��3�}gb����,>���0&�L�e���'?��3�o�!5������t���f-;�ʝp~ 2�z.|rN�^�1���	�&%�>c4�jݟ�3��hd(5� ��vJ�,�&5���0'a�=헬�|P��8�4��x8\�	����R]2�� <�� �z��_h�*V4�J�RCn�-�-:�m�΃V���/�e>6X���IX��m2;�]��1@v�)�QD�32a�ޱ�@q6�=��� �4�A� �>Fi��va�ș�|.H,nԕ�=���]�0�gT��L� �sU�B~*�0�X`�@�@*�J�uj#���`%���v_�#J�Nӿŷ���cJ����;��9�ۮ-��*��G����4�Ks3�i�랓��[��'�=��oӬ�.Z�fq�K�@w�b��ʑq|���UM����շ�N��o��Ē�x�n�� ���*P�4M�ک������#͑ϼ����g��� � �j�������|__�f>s_����?����p�d�٤����^|(��&�� �&N��3�2�~�Z�� :(��x'�.��	W���)T�AԦz��0����_>z�n�C��'�-]S+�S�<S��������+c�$I-���t&|�@�I��_zoNQX�Д��r�$���jd%��&��ξ=��-Z��ׯ7�륤�5� ��t��r��ה����r��g�sK��<_������sYe}�xX�Ӗ���}Y����&&�r���S��3u��/_`�^�UՋ5�tu}U_���g<8��b6>����%�D��ֆN��b7z��F7<��T#� ���03��9�e}��W���ԽBH7 F�eÝS�W#�f/
|�Jڷ�����}\�&�*؋�h+���..^8�j�AfE�p:�,\�Z � j�U'����uA��N�	|<:.�1��/d�;vF�0�w�m�O�(D�nl3����b����� Mֈs3��G��.� Fգ_!���X���!Nb�°d��4H�T��sJdLMvC)v]� הߋZ���I�te�pn%d���kp*��o�2�\7�3H^5.���'�if)4p1`~�֯���K4��"�kX�M��xK5�c̈�u�e��Pg�����̞&���[MN�/:��R4���G6c��H���[ڗ�������]���d_�\/_�CEy��*��`��)өY����u�h18xͮ��q�sڑ ��Ϋ\�ٸ�{��GP5�w �t&�J=G�^̊��2���W��g�M��G��.���~,	�����<ֿ\=O䂡;�y�Z�[�D)!������=�@kz��4*�[���0�L.�ʁ�X��'�jp֭�1�-AǼ<�R�B�M��h�	����+N-s��t�qhM�nɰ�h��P_6�_!�h��0xM7�[����ثy�kCg5�|'���'�t,NmK���[ij�o4\_#��D���l+�aE�����J��Sm�M�.�2����4v87��cu�̀���.�ʏ��p�b���Q��*�J������`�%��L��E�Ib[!1[�������	J0Q� �����t��MX�I�
��V�"��0U,�r��]=Zsݶ��*�ᵼs���>p���L�s�T���sc� l���Q��zy܁B]0��~�T|D��c�b��<+kS��d&��݀1_}c/o�uyz9�'�E��t��lE�i���)w+)�*9b�%��υ�Z�ؽ�k����n,g��B����&��ؗ�A�4� �� �<�1}d�}xFm�-e��|��Rޔ����z�#���d��]��%RD�b�N�ԩkc�`:o�J��@�4���"?&�]s�d5�G�>�?'e���΃a�'Q:�t���p9)����Q�� 7@�Š)���g�Ӓҷ�M���Xŷ+�-�w\=�#���� 8����!�j�_��T��g��u��X�~Ӥa�Vn���-��|�,P��_R�~�L�عD̪U�7�]�Mom�G��`��z����Ug|�����%]Gi���cm�kx�=�LM�K��7L"��4�������"at�����-$��J靣Y��	��Slw�ƌ�{F�DF5NZ����P�5j���|e���0}�J���J���}(�	�T����-�`D��&/j1�rj1/�1�?}���+Z��ў��#�̓�S�%�]�^<�`�o^d`��,�'*�A*#��o���8�����ܡ��[qQ{=���@l��.ٷ�
�䯥;۰DD�TI~���Q�٢v[�K®E�b�7�ȓ���V�0d�e�#`���#"�E,Ja\�	�kPo\ޤK�<�J).z�gp;-��X}D��y�:S'�����ΦdN�~],Q�Gi����#�ID�,��6�_.�r�1 ��m�p(�$����b�Y6��#�>C8U���r+�ul{(�M�|�㑚�7�8�ձS���!��x?��˖o�w�����Vmc-�ܕnC��D���A˚U)g���'�sI5�3}<I�YT�;)�Ef??7<��٤�����.�8acF0K�>�����r��;���Ѓ.�i!�@|�-}Q�WP�a��B�����𶳯D�5�h�y��s�/����k�7��/�:n����Q]H���7+�E�D�Џ܉K�s��JTK@�L�SH�&���5�6!}��q�u��A�@�V��+MM�6_��叐����r�q���ܞb�]��}����>�Nq�IW��iiZe	� �T���{m��I?�<�\��������H���
�ͳNԬ�6��Y�d�^��� *S��3��3����|��I��� �H;9?�h�������˼��z�ȼ�m_�!3�
�}��QE�L�������p^�%�!+��L�����L�t���WFݒ�u�$MtƉ��IS���SN����O��I�X�xL�6���0�- D���o���⌍9%�ۖ�a*�u�V<2/��R�Ͷ����[�	�(e��7V��̄;�vȞ{-r5��
����ap0�19%��8�A$�I]���p�tr@[]���� ��;憿�u�|YӢ��/Ih5tŀ�O��^$uc6����2��|�"����Ӡ_z���Nq^���)��U���wi�����5�	6Jѯ�CW��tF���Đ��ԞR���jmK-e:��x>��wh�f���Ԁ��	���b���I���d�2Ǘ������{���i� �
)'Z��n"])�S��0Kg^A+	�见�~�&�!�n�H������D.����@=#�o �w0�9��s����ʴ�0�H0����w�nx@�"L]������t�3/�}}Ε#9���+?�8`���{$2����V>� 
���j�ԣ#�U�-x����dᮔ���Y�����1��]��}om�̉�&ȶ��Vw�j�C�v� ��ނ}}�&��u=A�ssE?ۑ=ELw8�9o,]����0��؈])�RJ.���Y� 4�ߍTƼP�'�����+/,��]e�sU���I����d�l�CbR�$���gøA�n��7�_���
�2�9���-�i����s�s�u���R�
����mS7�~��R_�f�=�V1jjB��,��˸�^+�pȰs c}��a)�k��}'�gb�cP�4=��;�ȩ4,�<�tV��Gm��M0\Yt����z�N?��-ߏ�9̌����6My(z��C߁�rхP����� 6;h8��Y(/
�g�JP.8hG�Ų�+x%q7E�c�P�ܬ/ǳ�29"�D��A�hQ��H+ۓ�n�1d�kG���r�} ���ڋt�"�\�t���ыb=`�XY<�0)X��0�I{O������'v�6�%H��ti|�N�<:��S��t��'�\�y����DɣSP�"8�~#/e�#���T,�j?�ƾJ�)���b�/L��_�P��1t�M�Z�x��n;]�gP��?��b,�ԏA�a]9�Ϳ���p1X�܏�E�pc4(xNtT `j�.H#����]�6xuHOm��}��<�3�~�)�Jd�Ip������轤�H|������I~���	�H���zO�8�鑒X�Y��U��8�i�C�r\���Ү��0���ƞW�F����Ō҅�Q���c��,\��i��#�yW�Ya�͹ FC���Ĭ�7 ���U����+����"yQ[�r~��r|��1K�����NϢ�"�ک,�n�)����W9%$��XX�̱�(_����Զ�C�g�="��;i�t%�E�lΞŻ*����9�NՉX}��߰H�:2���'GoiAq4�� 7�+��aI�Āu���6���2<�e�7�
y�A�
���nS�j��!O�5C��?��^�,���~c���we��C�Ð�k[1��I��_`MG��b��5��8Et>��uu+���gy��z��;4��\�	���A��rL�Q�� )��!���8�ƅ�K�<)8	3^NI
��o��Ze����y�`�s�ˤ����Pw���n(2���AM�##��-_���%�j��Bo#l�Ŋ|3zO�m뾘�O�GD�p9�� T��E�}�
�T^rc�Z��~�G��Ô�Ë�вӑ5�oa�fxlnp�c��Ɗ����d2�Pk<o�Oޤ�,{��ܟ�"��9��uU���+�(�����/���^�������@��O|�jc����=�A����+Z�3�p�5~f�5p�5D�L�C�dTyЃ)��R۲��ʇ;�@z��@����b�W�B�in�6��hT#��N���S��Ď$G�e���;U��¥/�W���W��N�:o�a�u�(g3a�����r��Ȃ�m�����	��P��r�}�8���F�:q�Z]D�Y��r����AKW��AZ�s����L��5��ݑ��R�^ɟ\��|�̇���5v!����������!5y'J���w��[�%|:Pu��Rb55��:Q �Z�����A�8�_\�e� �(y�t1Ol:@�o���m�q�(Ql�:��!(�������._���pb��"6�oC�:�*��3�_ڟ���Ú/���b�I��"W�r����wk�"s^I�W�=8��y�Wz�证m�j�q���}���!���m��,��{��is	�k�`_�2��f�ьw�6��ұ��L@2�U�/7���fa�,v��t���2q@|�T���`J��vܑ�P%�Px��]ȥؒC�tPu�ޯ�����y�1X�/i�s��V��ME�[l���w�bU�4��f%����!-o���Q�M���k��EHz`��Xh��*����F3�68�xr�|+S�Ȍ4V
4[��h�
.�*�����rJ0����y��]�>��ez`��x���['כ�J�zO�a��*<+xq܌b|��֔��+@9��9�?QU=QnT�;C���z�J�~u#��j�*�P7t�����և�p��j��!��/�9;��2M�C��)e�W����ݦ�����
���qUr� ��B�������ܝ^���$�ѴQ�3�n�۷�R�\��+ި1Y�����,��Z���\F��sA����o�i'��URf�`ʔ����-��U�-�8�$�-�Oº(����8��w��P�VK�~��ċ����8������\�����4p���G%��OQ?L]��Ҷ[:&;v��Z}n�x>�/�Rш��h*Q�I�7~�����R��k�K���%ź����A7tͤT{��Q�`V
XV�KC�y C��P��S�Tc��>U�k��-f�\�#��X)X�q0����|��-%K����	)�"�h�\%#F���ju�E�<��c����N���Q9U,V�la�);�����:�0��y��%Q��HOԔ��\���<��8���S�Q+|�7uT�~*���¾�k��*`R��7�I��,Ҍ��+�%��rao�|Gp�[��Q0++\,�{�^9Hrz�#��ؿ%��h-�4��pPIR�VŎ	<gm ��W+��E ]0��|�nT%���~��7�9+�ױ���Тw�wSYǻ�l6I(�C�����ݠ��-�u%!����Rvc����1�Ѭ$ Ӹ��~�XQ4ݠ�LM���wRR�N�41e�g-�H��EKV>;f����x�<(�`en�Am1EI���^��Ko����x� � s:�xR�ￆ��4Fu���L3�t���_�-` 
�}L/��W'��١o�35~<�b���b�Y4�X�[��Hlѱ]�蓓Z	+p�G%�=T�2}�S5t�����ޝ�{3�1;�����JX��$����` �+�?Wh`)>�ݫ
���иV��G�jp`�\����L����*8���ӫs����,3��@z:b�\��3#�]�A߽
�OB�/����M|.�� B�X�W�������n���k]��gO>� (�XV^TQ�ObgK*�Jbc�ܤ���t �	u��Z�f��)��H��RW�(�لq9�u�՞��\�p�&d�g�"}֙[�3��9��z;��k*?}���>"ܮ��2�1�J���~�33VR�g.W�y�l6�
}!�'���L]U��Plр�k�N=*��2�p>'�)�l�����!��3a?�d�X"�8�i"9�O�������@O��*3g�r�nԃ 7������&����c���.��VH�T��W�:�=b#q�r��O�0�b��C���Ԥ�.��[σGM���r��3��ظ��Ůa�:.E�˒�q��-�d�CI�Ƒ�r�g�D� Z��,��L���egX��q���l���19��]ˀ�{x����d����/�N%�Y��m�y�HF����}