��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{��3ts6�vD�������T�̓C.�(��*����g��R(�����2���+Y<p���O �d!.8��A	���7A~�?�as,3�S��[�x�L�������D�KU-����@-溈��AA_^88C���>���0J�)�/��H­����F;�󛑒�X�tvOIB��j�T���|:��L�t�+:v�]���<�nl��ݲ&��c��6�Dw���O��,��",��_�F7tJz\u�
��C�s�T���{�aK��i��}6w�W8�oo����qT'�*�]�1�c-Ќ���?�ϡ��̚�5n���(������a����u�D��9^���l�3�/�'D%�zOHư�Ҫ��O24N�l�;"d�k�/L,��5�.:�������ceH�j��
 5�Yd�R)6a��!��L��nY�yص(�}�0Θ����y��q�,[��V��)�K�׌5G�a���~�n����]����?�J_%��������`�HW��`��Ɔ�������Ős@�����o)��E�(��f��Fd���F����<^}�>����o��>tY�;=y��iW��c�l������B���T?�q�d����p74��1���!������o��ڽg@F������y�������c���n��7�v�aW�
���|��2
<|���$ȹ�¸_�B�~��zn�$x��e|�g	���.@�����4qOG��u��-IC�AVc��3p����X����	�K����F��&F0�9��acؑ�h$0�)���iʿ��8�n�󸢏P��5������
� _�1���,�83�7�N��Ϯ�v��1 ��I�����2İ�J<�Wia�B��j��N�v#��,�\ͭa���G���H�H��P��h"�����c��Nw�7�������e͎�Z}�sL�:3�Hb��W-g}��"'�j�3�q�6|w ��T����9�W����,��l����̣�Z�1��T�H�VX0x�~_�2�+�X�ѿA��e���%ieס�Nd�X!�!���M�>�g!�:��-��m�ѵ��d��}�b�8���ջ<_�7,"O���Ra�;��#��-��������2�N�q�J���C$Ӫ�]�E�}����n�Q��#�W:fj��b=;�e��m�z)$����CO~��8���ȩ,�3�b	� ~�o�8 ��?��NF�l��5#��@k���Sn,o��+[�M.+6�j��{Nd���$�r�a� F�
T	�h�eL���N.�,�s�S�|̬Az�RK�|�=2�V5#��nӣ�]�#9f1pwl%��B�3�c@���Ê�+t����;�����.�IVE�/�	�9���r�������[SDw��; �W��5Zt!q,��77.���]?֥�ҫ�����/�@��b�e�_h�����V����,'���)��l$�4z0��<�^�G<+��!Q��O��E$�-��B���z�/��ݮ�A���z2-p0�D���y�����[����z@�^I����Km�	����@=[Wns��s��8�
��Hb�tW�|$�AU:�`jj	�i�2���v��n�e^��T�Ƕ%�� 5͘ο�B�+3�2'�43��Dg���ut	F)Q�l�J��*ɍ{|Հ\��T��\�x݉����]W?K=��y�p~U�{0o�'j�We�nh%�kGplЇ:	,:#p��^��q���+	������2� p�Z��x,>6+�s=�n���r��/��)�l&���؃TZ��gco^����������h�cX��	��Ҩ1�e-A�aT��x+�hˍM�^";�k���F��N_�L���o�{4�~[u���+�@�i���cb.����n���u�1�`��xs��C�A�)WxDHH�v;k�Ñ���j'�Y���M�+,��dV=�N�S n��a��Vۼ'o�3���u����V��N�cUt�~,5�/����ީ���܇1���v��J(����3�rm���զs����I�SH���Q!�z��-���e��zHET�[���#ۦE�S������1������>�gIa�f*"G�VP�k6Y]�?��$M��%cy�&2x�q����G�h�� t@G~y�j3Xi!�iY�Cη����K{fΑ C����reĜ'3�x%��q���@;
e���=sCm񓠷+�6��ۀb�Oavt�{"Q��0���Z�-��~I_=���^)�����VҘ9=`�����E|���aIq8��+:c�p�ވaF�=hl�1�#{���������Z�C09#(�n
7��2�N��h#�I#4�q�u?�+�{�S�k|����L�Ƒ5 ��a�6��g��`�׭�%�;�P� �}�[����'j��'�!�`�vT�]�DĽ���>.٠�2 �JO(����%���#		,��DqPՇ�J�wyI����0'���s'.[�S�x�M���xǞ+5���ޗ9yq��w��U �D��gk8S��dt��E�b�E�z��	I�æ����V�<�{����f]	����w68�`*eFj�yC��N��c��mgBb| �s2�	�*�L�7o���Wqz�ڐٗfڴ��[U24V5kv���״�V����=B�����%ei��,�R@�_!%��juX����:Hٶ��T�'�}z;���t�%@�a�{֔`���\��:��D,��` �c���(%��g�8.���}�k,Nx�����MH�����ºǇՇ����{Od�"lG/��$��&�[��I�R��^��ɗ�;	l�2���f���m�EۯK9E���\ޙ��I�y.ʤ�['�>sؗ�S�7�SB��\I���U��h�MC4�҃Z�lS�l��\�	"��k&��-�R Gx^5<���Q���,nO�zbvGo�X���UP��ؾ�0������!���Y��Obp�i���T��Ԯ�=*�IU@+�.�)^2uwDA;����f��.��A��4Q�X�q��'�����U����WB����Xjx88�x�cC���t�����[�^,t��{��2�>�?��7�Ȱ�P%�����q8@�Hi��u�"�|nhun��G�k� ����Y���v������ipz�)���,Tj��Ѹd#}����**�u���3��QU�7j��$5��J/�F����|?Ǆ4G'����.N��(qx�8{���爰F����^϶�ʄ�H<N���	k2���
 ߼Ɣ��S����0�Qw�:�^�e�7���*mV��g�j��vZ��K���*Df{Om���������p�9����z��M�p���@�eP��O0�Y&#"��Y] �Z�w�Ȃļ�Qd_��Q�*)�7C�ݛ�a�>�ʚK��K�"M��]X��	��-��;'�4#Śzh���A]���������]��[V���ӋC��[7� \i	]�z�0�N��� �L�v�����T���Il�=��P��IQ�į��^(D��Ĭ��;�:��8>�O~֕���º#��$0Q�����04?�qg���)hc6��"��$Ӓpz)ݏG+kCO����6�S�C�����65{K��wI�ˋ��uK�]p.����������c����M�d��0jd�W��F���R
K������z�z�̕u�s��(H9p���J��͒@��.�A3�$�V��.7V���n�v�I�B�P�6w����:`�VU����c��yW-���r��X���)iq�(�=����[�X�V5�\�uM�M�4S�aw�i#���Zs�n4g$��byzǩ3>�4��G���DN+�`q�iU��2$�5�qhߐx[�Sy��0��z�<�A�OK�~�yQ���RRk��i�Hb��!4k��A+�m�:��ʷ
��a ��(~��=���Kt�Y���,J._޽جp��u8���7g����}����m�6�\�(��#�c�LʩI@bZ��`�;����y5����|�C�X������g���X�53�P�C&,q�B�s量s�0Q^��FG���q+�����G[\�M=.���UM;�]�BϨGlbL���O������J��?Ce�]4�1d�ugN��ќ��K���������M�n�*�MH|�R� W�>d ]��6	�f�K޴5֢����}���p4���V�4��+l/Ƀ�)0j]�Jg4���;�A��H{��#ȷ����/���T��W�&�+=��0�W;������*�Dl3��/��%Rֽe�� X8�g}D0�s�
�[2�O�<I�r�u�3�mҒ�j{l�&�]�d�x��������y}�i.��r�Na,�ך��Z�׹�G���7l�G�˰�2���"v�r8v5z�`!�,����-H��ն筏�=�񚬮�
�j��c|ڮ�3b�x��7�`�t;/�{��bd�J·B�#<�J�ѵ�b�
�(�������<k���c�`c�e��,�oM0��zc4��ߙ���m��K�5TR��y�֨�T���$pMV��`�V�� }0��-Q;qٱ;� �����҅DKa~��]RJ� T�̃��l��I�8�%I@�&��.>�du�[�����x�?��Xd�Jǘ�k6_�ج�}M@��~A-�T�LE?dCMh���MH�{�e����
����}3�ʹ��U��qn��-VWd�
7㩏^�1b�-�)?P8*v�H��@��x�;�D,�4Y�[�";�w'��v�No�>��w�u�qH�]c
������ �gİ�����tm���ݏ�tJ3����L<np�I��S�sk��MȜC,2�fT#�-`��|��fxF���;�����CP}u:�Z����	zu��%��
��݀[�����d.ߡ}OK�!�N0�3~�Ҽ���y����h~���td��3}^rފ�Zq��O5l.IAlY���O[S�L���Վg���j�/��m�]��S����M�Y5��{���FH����������%q�� ç��W�"!5�jK��&%À+�F���{�P� �uO݂9�U���hk+�6� �������B�V\�`�O�I�c�����$��$��8��(8�i^��xڝ��lJ��B,%�j�]�!��pESs�&��B(>�uI�ҧ���ִ���n�{�x1|��LgD�hvK�vR�����J�r`:DFBn!�J���K��` CK�O�� �Ȼ6�|)$���#o��ba�3Z�i1��+n�w��O>K����Q�cϫ��X��쭰Z��D��@}��4x1zP%��ԩ����}�Q�.����)^ 
�+�?���Mц�o�jָ�����^
<��M��	���K�u B,��x��1�J����t#\j���Y�������l:�� ڶ��g5�8�ݛ+P��������D���e�kFZ?�~�����Μ�ӗMg��f�!�;=�QϺf��5pDuNT �z�x���.]��A��x*s�UD~|�ɒ���8���,�9�Y���Go+e�1�<�s�sd�&�7�]�P%l_: ��eI��}?�V�����s����[-M]h��yU%�������.%xa$�|少�~#ڠIm��]5�T{y��c��F,p}�K����S][��'DH�헚��M�&r�.�R�0�s��ф_`��$%����r8KBu��+
5�����v�^�[��V�&��¦��r�	նD�3���B}�^L7�8�b����w� y�V�5��Z'�Ь��u��,�gz�U3*_��Y¸�q�Q��Ť��>"1�SL%��1���&n��4��c�R �9T��K,�j�c�]��F7�J��~��> ����5x��c�y�a���[[��+�"��*af�.�tY��>S.Bp_�t�ڢ	�f��H}�湏�)��z�|ie��V��(��B�������b�!�<����T��I����B��&I
u��D3��������)^��@P��+��L݄�y���rHHjeh��<�:o�C���%��]<�A`so��- n�>� �h|_Y�Q�<�x��78焍u������O,1��j&����3�͞�3���N��5_�n���љIzO�.�"��ܶ�4��fژbf
�Ώ)R9>���wh��%�Xijo�����RY|�c�YJ���xލ��(�С��(yN�����^?'r�3����lu$�*��N�q���
RA3����zmЅ/��ݿs�F�]Xz�7���kjcP�Q�n������h�N��f]��\
�f���g��z})�c-����IG�4�ILv!��dƳ�
��'<�K�)X^A�I7�Qy���� ��:#*T�vd�O}j��V��/�1`�3�r���QG�^�~(&K������[�J%T�±�Oq�	��	-�ڛ�bg��\�
�	~���E�F֧���lP��c�A�J�d0��l f5���^������}����]Rp����������ϸR����d{��n)��-����~qf7	��%V�ށL��L��ћĭ�������1S��B�q����S4����/��[��˶���Hm5�x����Q�Z�����EcWo��פ/�Vc�I�&fO|��������Y�����Ţ..�O�;�ֻ�':�q��u`�1��ޏ3�׹��wSe��=MCz�y�8�ܿ=*p@��JI�q�Y�wn��?a�����t�êK�� ��z��Ոa#��Mb�Ӯ��J�[<dq���f��t%*o%@��j�wa'T�IlD�4�X2_���8&Mn�5͊Ǽ�?�����J��K�����,m�9a;|�%�}��s긘ǖ���
�@|��Í�d2"G��~Bp�(�-�SOH�ξ��9���d�.�26M�t�Fn��?K� $f�T(�hWr��w�����_V�/�H��l6�����Ҁp�GgH���O�{�i�5�}?�ob)_t\��*��q����6��&~�򅥗�vX�_�c�/��v��/D�f�`.vݼ.�����7}��5��)�
�w$���@X�r�*�83��V��y�������pJ@Y�^㔰k��&���6�v��ϣ�M��D��1٩+�{��QbU�/7���F7�F����7�O��<� ~��w'[O�O�u���7��E���H��*!�8��r	A�).�=[rZ��TT0��>���P�VQ��5B� t�zþ{9�pSF$&����grܙ[�Mzã�k��3k�4rEG8ѵ��p�c�_	����IHxF?��5��V)���ht�������^;�U)ӻ�i��ḯ���i Y��[�_���l��&���HY"HB��ũ�t�~�|��Ȼ CǎT�����$�LJ	�^�U��{�7�Q^h�3\��,(��4l�	�>^A��^%�>�//�o-r��i�v.3��2�
TĈ�8|�r�����h*�L0�\�1�!�x�'�f�HHr�����*�J䫔
����	��ٶ�P�� 
���W���8,i	x�ly�m�
lQ[k�:�>�C��҈J�@�㖑F��n(��U�{�v�oe�T�W���<�md���h���=��5,�Ƹ�P���f�u���z�OÇYts�!�VMC�܆��
'
���󭐣�K��q����<7Y�性'w�a���p�A��Au��:�)��;nK�.�l��)!s�I����L�R�X�[�M&�Y5[l�!_�7�@��&_���*/:`�HX�l��IW��
�0��y$��(E�cT�dT���F.�&ĥi[��l����Fn���A��whQFnM���-uoʈ<U4oQ`�� �[��6l�Z#Aq��÷�z8�=�3��`<���B]ϟ=�����\? ��%F���-���`뇢-�w�_�G]�	�q9AX��g�_s���w��c�J�1,37��Y	�Sq}?��~��dK��AГ�)�9+�-��٧�l r��P{Y��Vmn�����D�+����F�]-���=%өJ�~������'W_�Rg'$
��)��P@�E�&�Y�G�3�=ۅĥ����h#۴ܦ�_*�،���Z�G%�מGS7�g;��Z�,i��H����b��j�kF ��	�
A�Xc�1Y��<Hi&�z�-5N�#���s��Q�Zo*�9)rH�5/Օ!J���iU�
� �����j�}A�;���fhQ��:ɢ��V�jp�w�ǡgdA���?~kE��u:*T��R�
<ʹ�J[���^�L�睅�������� ���=2��3g�?�3�C�V�M��נ_�F����m?�L�iQZɏ�?�q$�r$��6/6B�d�~j��!��Qu~)(T��Ҵ��"?9?�5	1;������NW�'wB$t@�.�.n��IHQ'���n�,��_5b�������!�E��]������|�MaA��Nб ��#>4�V��&'@�R�/~	�4�d� �� 6ݹ�cq���-x�,yB����aߨ$(\�D�˞k���6��R��Sg��O ݍP��x�1���)Ӯ��J܇m$�|ȷ9im�	��d�5��_˨=�D�ʿ�C�6��I�? �v~6$ĕ�ʶ~!=��2����oe(��L��.�ĨtR���dx_ީ���W���s{V/���fg{Ox-k�p�Yr+���D�R�Uk�|�?qFW���ܴS?9Ar�E�C�SC���� �<]I����]5�D�b &��P�N��Y���`��pD���၍b���$G��i��J�B�8�����p�C1����0�lϷ�V�����$�S^F؂����[��I,}��Wڊw��˷*� FU�ëTUr����줷��ǎ�h��s�P�
@����)�<a�sMץS!, QH�N��`�����E�5��w�V�].�9��a�vK}��ҟ�Ǆد�W[K����DM3��>�K(r�$��N�y�XLD����eu0�o;6m7h5���B��!)��E��[u�"�9n��zh����~J]�)=0���+���.��3��mv �h'��<Z��#ib�_Zp����pB�{���.�|�2~u�J��$Y��M�r�t�L�İ�%���d�^�'������sO��<�����ѻ�@�9Q��H�\'���]�GeZ��'h"�&X�(i�`��l=ԙ���Y���?��C<D���i�5A>3wc���Eh=I��{��ߙq��/�#���3�lU��6���� pyU"�s�oc��4�Y�u��gc�ӳgM������ߣ��=�)�y�l�M���i<����jK���B��L��m����g@�}��8�����a�ц�#�ha��$���{ �z�{�8c� �oe��h��~�-�X�����B�1��Z0C���Y��N��޾Φ���#Tj��,��@㏉���A�����kPk�'� � ��T���ٰ�6R8í��"(�?���F ���[�|�=O���^���j1r�z��;v?�sr�����T�}@�^���������N؊��4�Wq]Dl]���a@���ۺ��2���%_�0��^g�*1k��:��������_ش��GR�^�Ha�
�'�-�sW�v8��I����/���_5�(Yu���[�a(�4�>?y<��1��z��6�U�W1!�ڈtE�I�C+�]��o~k�V!>]p뒫��x{Rl/�������|f�7�$v[�ء��l~6ƥL[�ϟ�3PP�p�C�@ڱ�x�.�-9�N��Z�7/S-��it�Zi��	o���xF�HY��E�Y�=xv:)�&�d�T�U݅�e��$�ܑ��n� ��ݜ�^��x�tM4�;��̟ە��}+�vt8��[��2/�Hʶ˾�d���	�] ���Eb]�/�s�\���>��9�����J�>>�v�Ճ`=��
�E���|4U�<$�
H3���0��9emf؞K	)A.;0�;�[:1{��U/;Sֶ��7�x:�����j�[1���OGJ��vTx����aM�E[z���w�P�)i������DH-w"���prd1~~��M㑦At�=��ʹ�QS>dT73c�G�C����(��#i�x�!��tM����f�W���'��d�QC�����ʬ��ޯ�ڈ
��Db=:��EO��a�/�\����>EH����?�6B<�� �@%m�k��0���aG�x�`���d�,%�������a��_W �V�e���,�aQnsB��$��u&}���8z����5
����x��:o[ 4	���#���D`���� ��_.XB=��#0�z�YP�$�C�>Hjc�%,��Y�n�!0)�6� �#�t����ٰ��c:[�O�����~��aI36���%�3��X�L�&	#���Xh�{�������S���3��k���Q�����.)��g�Z@-�)�V��pKƕ���A�+ZQ�᯴w��6)q��AI;�����(�N�*v����'<�|���-}���~y��밧�ѥ�/��*�?��]�ή�/*}9�*}v�e�R��X+4�3����7=�LS���ڒ;y�C��t�b�L(�t��Q��Ӓ����Gr�Z�=.�`v�\\���C��d�ҷ�6Ň�2����D�Vy퀎��1#}	9��{��ЗcgO�׿����sM�l|���r54�D)vV5x�"�m�5K\H�Ռ(��v�3C�'y���ݨ'�YǈGE������Bh���Hu��8����7aT���]�ǹ6ҢbDa1�`���խ�d@�l�ޓoM$M�}�ݓ��O[�?	с���֜8e�!�����N4pw��ŗ�,��=o#�)������"�d$��<����G��?m�(�fZ��N �b�����v��xP#`����	����CN2��Ia��k�4k&�u��:+r�|�~P�R���xd+�kQ;Q�0SL޷X~�lj�`ף�~�-���YH�>"����7�k�R�P���HP
�q��Fh����d�G'o��d��1p��PQ�^�����a�:	rsё+�9#T���f�gY��#�q��by��Y�b�'���v���<���J�&�A���>�����Z�9$���P�Ɔ�qy J��h��`��4��s�Z���V���Mfǐ'wJj��|���oh�6:��|�����,�������i)��rU�s�4bn�Z��~�`u�(�ì�8AG�����$#�L�}�$ﾔSBH�6���(x��7��P�R�q%k8��BN
��
���\���HnOcB仢��v�ϳ�M���,��EͶ�|ĳ�����c����b�����x����%3��T�����u�/���
�W\ĐpЮ�w�����b!�X��7�Dʸ��CB�"(��c&O���)�.�v��1�SmMzQ�kA�=�[Sge\��o�"D��H�g�ɏ�(�'7���"�x�[EhJ��|
 @K���֔�>Q�u�Ej�tLv�i�������R�+�B��v��rD7������* ����ܝ�#a���M���kA�+Q}�u?��ל���r��l��Jd��@���4��C8R"�X��϶]Y�hۢ�d1 G��0�7�1%�F�lk;%�8:W��i���ޯ����r�F�~:U�����v	�����<��fa��}V>p�2{�Ұo�T	P3I�3�O�-xb��B�(�� �d/�DS��;5ɍ&��UɆ�rw- 3M���ݤK4�u檕��o��33���a��Wg�rP��>B5�f6�P�)��W�@�>n8�\/ح����b�٦�:		�
�y�t����N���,��#� gĶ�6@����(�@��f��'/m�sP�����D�4G�<;��ۏM���)�".^_��|���~Y�Lf�};c39y8�X��]�.#qҗ�i<�G ݑO��T��>ٍ�LF79g����s�$�] �mxU�Jk��F^�����=k��v[ǖ������%(�,;4D�6��A�q�;sةV@D8�= Zz�vB��L��!�{^�D����4Z,�$� ?:��!f��̮��,¿z�C�/=/j�C��{��}#E�cpܫ/6'N-��hnf��h}�x�s|��8�z&vGW{���� ۋ.��NF���� ��h�,�k���q,,f����a�?n��O�O�Rd[��֐}&$���6�!cYR��3L4�e��aMO�K��ż����
�):�X�AAƻf���?�Ùel�-.7}����}�z|v]Ҍ7dy��n�8� �U�a1d��R(ͧX�|�A?K,k�Z���������S
i}-�q�8,,2�/�SL��NRg�k����tr����ǳT[�M?b�),Թ�YH�B�C�_�����m�� ��#꼲��d�Yp}T@�(x��#�9~��@�����𪡪M$�!L�%���������.��@����N)Y��>O�_��CE3�C5��c�J�l,��d'��OfBi�����9!/G�tF s�f'x���jX�7,yn��Ҩ�M|ըh<�e;V57ku�����Bߴ2M��Ⱦ��V�߯�"U����ϻ��g���kH�p�[')�bU⑉���.�z�<UZ������Z!>	��{32NƑ4�� >�$b+.�~�T�yv�hʺ�fD�Y�>�ˀ�j
U`��a�]��T�j|�D��>�}&q������C��̎����̭m��' 7�x(�g�g���;�7|�����N�ewp��`�ׯ���lJփ���p�wp�j]%���)ι17��ǃE /P���ͪC!��5Y�۞���������K:*D�<8�MkVa�q���mm��$҇{�j��C�~2g�$$�[H�G��`Z������m��rz6`ԧ/ۺ����G��6�{�"�hW.oѓ�׎�I�S�y+�>��W��lM�=����˘5�<
�ʃ@�pt�_�Q�3h�'�V�PN�c���F-5���6<�2�o蠻����?�yq���qxo��6V�2j�4"���r+k�Ñ��egDK��~E�����z}�^_HE�԰ݪ6O�Y#?�VO��׭��+*^~���Udd %s�M~�ߜ�Cw�H�2�̧�@��'!�j�ʠ*#jm{1y@�ͲKM�;��O�x4�v��9��m��dw������涣��y�ɿ٭�Eb� S��?���BO��1�����q�S��X�,�靳7x�
����`�6�|�)�a���_͇�Pv��t^Mې��s=�iD���L�P���]�����U�;���y��h0R�m�����̬�A��Ы�C���{ u݀Ԉ*��ǟ��[��v.%�� ���*E���M��NY�3��5={�.��\1�iT��*i���+��^�؏��&�e�����t0�c����M?X��ErN�n�`�_�"�^/Уm�wL]�uʲ-]�Z�����m�vh���(��0�t&�VD��C*�o$��� F�h�ͥ�H�_X �;r+Tj�L���)�!^"r�[@Q҉?O��]b���W���䷱�tRbT��JrN�>O�̩���\�#�E���U�0~���7�����1N|�x�! ⏒8��V΢��@��m�1. %~�J���Hb*����a�h\��Ɉ�#?�z�i�0x���/��L����-U�������	o �3��˵�h�!�mͼ.	���;�P�&�r��[Tn���{-�;����) &Q�j!��|�~;�Gu0�� ��S1�6M�o 4l�31����T������Y�1�����ecZC�^`]�S���շ�,���e��V�rI�o�Ca���B�g�jT�+����zr��F�m�D�[/afƿ.�~	��F�Hߵ�Δ'̇��/��z��["���;'��O��6OJG����o8��E�;�g��SM���J�$6��5 Ծ��Bev�$�I�9y�����(��H��]�4'�a~��s;��������3e*��U	��4���-f�<;Z���<�c}r�)ֈ~M��,�؅��!�u{{��]��>���)�L����G5B�O~R�J`d!͆G������ סۉE��M���2?���/�X.��0\��"�h,�&rF��tfS��O���s���f�>;�dܘ������՚R=�)%)un�kCY�A���c��A�׷b��L2�a��e��bS���"qC�̊�qk��։���L {g]��{ڛ��0\~�!e�卞�
�?��]��xt���Ƨ\ eJΝ���ay4َUMC
`2��d���'����v@���{��l�"
ΐ�@��C&��n���(+��m�� �z"�~��c���̿� ��ԉ�fSIM�]VL�W����m��vR�����	A"#�ʰ���)��Ù�QƂn��B�r�=6� �ې����a9�0O���I�R�m-��6�zDm��n��"3v�<[��������Ah�A[d"�=�v���!���-���h8Y��N�X��Й2x�u�i����:)�skμB/
f1��+@^�a+����IlB�q��z�l�D�"9�g���.s �i#1�����Q��gRX`j�/���RO�u��k�yB#�)��攴�2�<߯�9��p�y����hn�����~K����-��1+
N67*��l��:������H"�Ҽ���L�(⿻y�ǉ3�*N��s?]<Jk$�S#�֠=��,;UЧ�ǆ���t!9:pmy'3�:7Q"�*���4�t�qRT]fŅ2B����6��(�iL60����{�Q��jC�l�H��������#h�ӌ&l��x���<~�!"�A�?�u�<�w��:�M��O��PcԾ9��Y����(�S{2E?�����\�7�X>{��WX2�ܓ���P�c]�&C�o@<hL�KM<%@5���V0.r2t�v��>τ:z@ygx��3����S{�U��:G+�� �p.���)��v��US�hm��4s�,��"nG��w��|d�dQ9/�
�&�`��?����I
?樫~�����<0!��`�|�aG�P�\�K��B�/�j��p0����E�ސ���d������uc�Ӈ�Kb�GF_��S��b�K"P��z�,��8�٦]����R�p�'�.>	6� �On��v�`�O���t�h~2!<9Ȇ;3�٘t���k�T=sTݼ��;���$O=>���Uz��lT�}&:�}��}]�X�nOo|��r֗B��F_H�c.S[}�3&�<� \����f�:"��ٻ=�Ȑzo|��9���D43�aشt�"o��c��@�Ǒ������a(����q���mև�5:��X�d�����z�0(�_��1��^�`��k�p/�a���D�_�L3�C z�:C�Ο�\%\ÃQ:h�oڍ��.���x��/�'[�Ŷ
9��N"ǓL �,ЏӀ��-r�'��A���7�dU�c8��5��r�H�8|�2<ş��ċ�pA�?[U�+0�0��j����&�2Z��ds��[�Ik��pfi�*��n1:���
l�P:�;!!���������a&}Jd6���I&p�y���~<�B�Ȣ�>fvS�����E����sk��m����.����$�|�����L~Sk�Ōñ���@f_)澯��mv�!dp'D���b�O��0G�ޢY &���pk��O��$���_a����ެ%2nu�Oiu9�>I�]��S���E�s<M�{L%¦p�Z���S���2�0B���&�q`��٠����5����&��U�\�\�
�SATX�Ku�m[I�H31ʗm㏆41G30�曊���ͺ�M.��C!�uP8��}a�;ƹ��N�Y|��2� ��#Ⰼgو�=��tC�@���$͜��
�\.B�� ��3JK(��B����2Yz��{�&�H����sZf�hi��p�~wr��*R��E�����|grM��:�Ve���O(B��5,����L<x��XOj��u߹���~�f�Җ2��ʗ��G~���Ք^�`��ϋ�>� ޶�I�dp���3�fU�b(����ucK�����XR�7M9ƣ�����ʛn{5,�
��;�Mي�o�~����FLx3�� �k/Uk�^���e2Q�%e?��y!,�dտ+�DYkQpq7-�5��,����Z����Yd������z�"�$Ո"B�=@*̇�;����cD3F�����bO���pI��zt��&j������YG)�W��M�vJY�?��6yq*)��PWF��Za��ma�u�܉�����k�7֝r�]sP��|rio8˼�橺��'��+�X�1�'��C�f��0Z�,�^��d�?�i���z<��S�L��A��F�{8�_tw�?	����l ��#��}Y�m|럆OVI�f4���.k�!��ٲ��	�uv+�֧H0��w/:�39��N�s��[�k�ѡ����>�UF���-���袖TIK/�l˄�{�:�ǈIEmqsb\ѡ����_M��r�iC~�a�gGښ��3�E.�z��m�l�V�7q}������Z7����sS�������8�2�k �"��q�&�m�+^N�㾧��MnU ?vB�V�[�ַx�F� s斲϶��qT���ixw�'��3]IIŻ�D�^9�h���j�\��&J�(6� ?��|4�$ӣ������cqP�?Y�-͖��3�`����L�I�r���]o!�U#!�⿐+�-A=�Sjh�K���A.|q�k�[owK�9; M��:6���E���њ�Ұ�� ���g�3a�ѥNA�a�k���>'��k�O2�w��3`d�K��Q�4=Hz_��a��Q�����)�j�����~���pX�#XRk��q���%���[�����39a���<+S�f�kڬ?�'2+�@���p9<�
Y�OQY�AH�#�s��!��H��r��=W���7�@5�g�>iC~����<�=y�ʓ_=�A�g����U����;R�9 �^}z+��O��� ��v�W���sH���> .�M3�c�������[�n��<	��M���:1�6T�"��(��+o8�6捀a%��`ڡС�Ғ���3�[��ںae�b[$ڂƭ�OOB=����Mz�(�Ȫ:�� ��u�GPoS\���˙�0}��$$D�s�>�T�3�<�h�k)4=�צk~���Vr�H��W5�N���^�!)�'��@��\ؤ�������k�4e�z�ce���^�Ze�}�T���Z?ziW-�����^wK��q�5ͮ?l]�e����c�,?�x�����.t����ї�rZ�K��a�j�{ÿ�h�2����.ȹ92h��Z�H�J�� Fp�I�Qu����P� �YJ�1�+b`�h�XD��e"P�� �����@�����]<���rV���!hVSFl����D�v�{X��F��p3z|~�Iy�8-s'�T��+��OeK"�i�'l����/���^��A�F�������	�m|�V��c�����x�L��}m�8��QL���:)ZO����UdW���Bt��J�:����3;��">���{���Я��~���jv�+�2��O����zC�>��C	rf�Ѻ�ûe��W�P���^t"�1˖@p�HjK�ٻԏ(l�X��G\M�@S��F����V�7MLg�Ov��}�c�,�riq�~�qAj/a��<����ר�o���G����6] Zid���뒱"x�9K�m��d�?(ie2vŅ獳��N8)8Q�����.�lB���;b�S���;����$��A�p�E�:Zcw/r�->��(�1y�L�\��:��ڋ|<o@W��b��mڼ�F����%7�"�����G�B:��]����&w�<��"�
��<�ѱq�9Qc>���[��5vr:�������7�[�\�j�G��H��i�RI�L1���xR3�y��x�*gT6bDGhG�S�H1 �ྰu%㠄��X4��������![�S˲���?��U���s ՛��P�|�uzp�-�5����ā�L����	�r}�N�W5��&���������9�/Iu�|C�Hʹ��
eƱ�N|&%�]ߴ��Z�[E^=�N�ڴqTY,<���'�I��p���"
+� ����2�T20��͟?i_����(S��7Y��`�RZ�z1��.#����������l�@�h���-�u�����8�zR-j�q'�n�z�n]���A�O��P�;��QN�N�V�.��^�e�i:j�bR&}�^�}���p�0��w��r����>�GWw�w+����w���)�_a�r�e\-����7�+��O��l��J���}^ː&�^�4�~���p�B��c)
2�X���