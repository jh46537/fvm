��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0����>�P@�:��N���F�Q}���=��P� ����T�3��E�!by��3�Yn'�S�y��T��P^�3y�E��pzwiّ������l_w��
�5/Iӽ3ݖ�#C�����պ��o��ۗ�}L�-�ѥ��&4�u��5J��v*:��A�S�ƃ���Jg�qS?cZe��W���y�*/Q�"'�`�"�"u�f#�pd��xaN�D6h����� �~U�.�u����%���OÈ�^D$?����O�6P�H��퇱(��pM��,�`j����5O���_<� ���;R��#� ��v*�1O����(�񎜈s�xQl\T�K�=�YB��ȪՌ��vL�^�~�m��G;�M�T�AZZ�C!G�k�@-���s4��{�ʾ���`vI˓_���:S�~�]t��1�W��2M��Z40N�b��?|�ر�G�@/f��q��i>��2�
>C�ʏ���s/�oc�L�9�DTH6�2&������-@�$���2p����|��L��ѾC���2gg.������n8ן�2��L?2x�����M�
�U����|�g-	1�ˤ����=2���o���/��6�{D�в�# ��
/ ���t����]-�}��O��G|�iBi�r"q	P_�J2��28b�HЯ.1pRj�ݳ�"���É�9p���HY�׸���
�!d���@��%�>λ�A&�v�r�xPȍ~v��>;���fOTx*��´���=44c�L���W7�.ݿ����%�hmC�VH�<z�[/����VE+bj�Y=LDh�wu7�t���&-Y����7��4�z��S��m��A�`�(�$�Rp�MA��Dܶ3�%r:��=�� ݣ8DS�Fj\+��87~��Fҟ6���
%]�@fn]Pi7�[��P�n�5�TN�c�q '\���̙So�胙�o�Wz��cW+jꊶ�
;�-u�&t�������BD�����&�*��q�&0�Asʌ%Pwn(�F�[�^��b))��6Un��<ly����d_v-W9$QsZ���B�/	��5�����r����\, �gi�y�A�s��Gd{<���	p�1��M�E5�x)��f�Дf�_����n�:�Io�J�{�U�r'5X �E6�-6o4�^����+���}b�!ytT��n+�����	n���]U"%q�%�^��M�^�f�9![G{�����y[g�<��+��G��_2���֮&V����dҾ������Y��]n��s�BK��q�*G��{6�<Y�P!��a 5f�[�0��Rt��xy�!qV���DQ�)`u<���:��	���a[��D��i�`7ּ�����&�l��p�?�7pu�{3U��dFw���5��u?��Mc+E�B�9�>�+Gr�O6M�1ܵ#Xk��g[��gq����i�"�?ȩ����P�����ĸ�_�@%�i������v�6���e;}rC�X�l��N��n��{��M�l�PfLAQdÆpE}p1;��vo�B�huDO;��.&�{�g�i�4��8,,T͌\�����,��l|-�v$[j����G�����.�K�͐}� �<Қ��0�M.
R�P�ݛ��#Ӗ�9��!�c��	��,��:�G�����!�I]��-xq��eF�T�	z��qH�ǁг{nwB�-_�O��;D�?rۢ��.��~Ž�Z�����h�h�W����y��GȻ���&�iO
�7޲0a�l�D��dt���/ Y-z�o�.D�d�ۇ��(��� �
[��_�!�;`��T�S\=�)A�ǥB_I2o�I�x&W�Y�����G���ۑ�f�թ��6�:CFn�ƼDnD�Ү����F�ᦧSk�c�M5���]���.���=�e�OzU�T��<��F���^(�J����˷2a�|�|,�*s�Z~���D��h�Y�	S��R"�c���w�
�zq%�/�^��ux[���z�1X�N�b����]�
��1�ik�[ ����ho͛3��Ǫ�i�Vơ؃��;�������'�5QJ�>�ΰ�7y�WA��T��Yf8+�Ȕ�]|3���@dEz�;q],�|���