��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����u���y��O?��u���
���XI�����e�����Z|��<��@N�B���dK�s���Y|�0�����H���-���6S����+v>3g?��a�u�8�1k���t՝�5� �8ؾ�T�n�T2�DjD�^扷>,,��?���m�B�fP٤�h�驲o%Hۉ��_-� +S~_�j����m�Rr(@6µž����ƹ]/���Q��)��e2�q���Q}@(sZ��\@6:�̤* m�����Y����U+����0u��QP����x[�����W�^A�OR��O��r�qG����6��s�`�@�qZ�3�����ah�RoѺ�@]��>��H��|���>+O-Y�!����(�������J�ڄ��+�#3�I�@S�)i��j��*��XG�T�emr��
�[��h)�y#A����
���v4.�hLmA��� ����#��~���\-���:gÄ6]�$�͍�db�IJ�������X�[�����wG����]�c�#p5ϊ6+��~}�/�b^�S6>"%f����F�7�9{�l�ٝ�~�< g�ddH�EI2P�!�9ټ8���0%p�g2�S�D3�¬m�a�2��1V���-���@��~Gq��1��W?�C�ؗ,ER�hN�<��l1�/�����EO�C�6���T���o�\Y���К���,�X�s��Tpfa�k�_����s_����@K������-*0�S��^wUA@�@��9ع�֩���]�ty���E�j��a��f�s{�hP�Y���"Gߧ����q�?ʁAa 3�������G[�f���S�lv�����]��5��E��ƹ�N��l9T�Y�Ś���eALs�'��=�Td��~e��*!9D�I���_@�%�����`����k|s؁S��^H*~���FH��h��&���T��V.y��W�n���h�8�ݭӗ��
���aY����UN�����=\0e���� ���%������
��� �PJIյ�o��G�M��J�{��9�1�jd<~���b=��Q�����?E:��\��+��	�`�xs��'�a �{�&�G61rE�t~��AJK��U�O�,��c�u�Tkv�a�~X�r��n=A�y�/l@(��F�Ut�@�(R���Й�S��G��$��_Y��)��W-��F7�v#���XK���I�!��$�Z���uz���@��%R�s��(�7�]W���t�@h4�P��1����X���f>]ȑP`�^��qK=�ջ��˫�_��z�za�l�ϳ�i�j�q�c%��z|�j���������Ņ9��H��XL��a pY�sA��~��H,n��#0n��S�"�\? �V6FZ=���)@Ȗ��LV���~ �cBQ���E�Aul��:��h=�ܜ�ާf�;�UVr���=������Ettm�/�ȝ�o��B(h�c�!��������U�v��(b}��@��n%ߖ�M��-挕�i?�i�'�ٲl�%�=<� �IY�J��9��+���<ô֏+��M������2�(�jc]1D�y�17aB�(:Jb�4}���i��������u�!���Q����D�(k�QV�	y��A��f��?��\W��%���?]͜��n-ׇx$��c�~}���q�C�Z�RF�~J�͟<��,̸�Q�tj���<T�oL�����P8#�������� _)Š&Ȧ�#�d|`x��1�+�.߁,�#p��N);AXc�����|�N�`@xsf�9����]��Ǭ�����FĈY�w�ϬM+�}o?�;���T{N���_}�]P�Ã~�ƕ���)W� �O�7��G��A
�H�0�_��+S�8��v�`��ӈ�Ã�Z�TT�f�-�H,Ԧ��	�}m����\��=����)<Y�2]�Iί�}�	=����['�l�����K��k���Ir��^�CV���+����?�L��B�Dc�=��`�o��^�z��P�1�]�#M#H[��H���q�� ��G7<���T��\/_��b�로���9o���^~��l(u�
���cg�?Z�vT�R�Oje��>7�\���9vP��`&�ZDK`:���Sn���n+	�8�ō�W0�:�/����xw5���� �76��wm�
���o�"��\�R%I{[�H�j��3�⦩�0���Ɋ��)"�~pR�-B	�{��>l.���:�_t ���2��m`��hU�z�h�h8�5ƴ��2����b���wd���3(U,��T���/�H,�!�9/�cǢ�ǘp��͉-�x �|Oq����Z��ˉ	E������]����9�/��yr<?�M���=4������]�Yo
���uGl�q��=ptHR�Pý1���2�ܷ5�B�C�Q9��r+�⅔X��+��$�3��쵬~�J���RǛ-g���tG*�+s����A��\��IE�	�XJ�Ime�)���3@�7߯A�r�"��~~�/��{@/�wg��,�/)� L�rܧ�b�fޣ�GdN`���^ө�����R�O���e�{b@�=���ѻ6d�t�Oe�6iY��U���WlP�p���U���x���["	g��큺�%P#ֱR�e8ݙ�2CV����A:V�&�)n�鈻����ŉ��V�%� j����@�8�TXI��kxaHi���|�%��P_q�I��R�q2~�u�P�y��4х#�*���Yngׂ9���������J�wI���\��J��ƞFq9-�Z��y��bWdKd����ͪG���[��E;�[
j�V�US�ʌ�6)hW�'��?)Fѯ�����`�C�۱���h�rxj�+�U��}�pC��dF��!a�8�M��6�l?��?ٜ�{I�Զّ��kA�*sNb�Op�K{bW`.�Kd��/]���\�[��x7Rc����E'�R�8���u-��-�^�i�"&�#߉���j7�E���+��T��6V�����%~�e=۰xh�ר���]���V���Z��+��������.�Mj��bp��Ӑ�2x�9؆��<��b��iyհ��F^����wˊ���y~Ɵ)sxgQ����E�~�c����%�|`�C��ţÊ|ml�~�
FA�9.�Û�'�2wxua����jS�4A�!��¤��:8�BN�ɓ �I��������	Ƹ1�tz���>�2~f�7_� =?D6b�:|�T���,��mK�=c�x�_���9�԰������TcF�H#����-lj�r�\�%:����ϫ��q�ί-}؝�2�.�p,��[V{F{�>�9��f0�&�^Z8���5f���E߰��Yo9�
�Q�{]�Eyf�5�Mr4X}a 貽-fOf,^"9���Q�Æ�,B[�`h/����ߖ�"W(����'�6��>)�[��Yuۋ����a�G�Ѓ'��W�a��P�`m�4�f����xEҤrRcn厛�#��e0fΊ�~_��E�(s�2d�E��*lsR�������y�ջ��ڱQ-�����Ұ]d�Oǵu��V��o)pþ��_X<�;kf����&�x��ЫoE,7�#o2v)��TM�I����Q����e`ٜ��`hA�;�ygJz.��v��ܙ9DE�̖KT��+�a=��8�p�iz�Ç	ǁO_�M�_�5$o9��(iԪ����o�s�T�>)1�Ѻ4'K�Tt�i�/�穹�} ��R	Q��%���H��朕�Y�H���Ir9�j�9�oRÀr�1���(4!:H��&�rkn6 Q�7��������v=��aW�2n�M+z�+�Kt�^;�$*�H �+T �H�
� k����M����ߍ��솞�,��ԯR��R���-�N�;!���p�Իn��I��e(D�k�J�D�T���˸��w����F��+���8;K�Ϝsչ�!�Ѿ1~;�X��;w#���0���}f�:Ty1�A_�?}:BGƻ�r���^�qۗ��{M��+�J�V���CZ �I�T�B�`�_M�j��/D�
��1�Iu���{���
�(�4=tEYS�P
���v;��]4�i����Oa����ǥ�O��V��@V.�@�b���W:�F�lU�˟�N�%�w*~.��s�&9F�bfe�\��Ҷw6��@�4��V�<KB�ߊ����}ǀ�z�i+��T�O�����s
�%bL3
�ߙ��"�7�`�O.a�ۣpÑ�sI�'���'9���(g��@}s�_[��Ty;�,�����Q1y�q���ftUE�*I� -p����F9���)��U����S0@���P>y�B��,��|�2H�Ş�vz�I��x����C8��Ӈ�a3�뒈"0u�mQZS�د8OK����0��Q��{�mS��9��~	|�%�P��KZ���JF�������);���?�
L-��3�[�d���N�=���(kA�}����^a��}���f:��c�J�.l>�v�u{(s�H������|tls��)����c��9��T�j�D�U0���i�=�Od�=VL;�N>8��F��cv�C{���%dC���*��y��&M3���k]�j'V�l�k]ᾢx���)<SJ�d��S+�*QsyM��H�fe��yPPK6\� ��@����tꐛ��ϳ�H3Y��\D1����
|
}(e��h�o*b��I�pi[���=xz�y:0��]�_���]��Ŀd��?�	�=�_m�*�a5��:�$+��qA�-���1��
���6���U�YY/Cw|8qr.��x�3ͻ̜�.��.�9�RHm� h|�*�%��Ճf���u��i6�ڠ����,}HI"�?�-%��T�TL!^��.$�`5��<�g+_i�^ww�l���r�����I��8D�w>�<
B��:eL�@���{�=���[Y�mi�Gy@R-^h�V��	�2ݭS����G?�'�|�E9�	ό�`cr4�0����q(��C��܂�_��s}�)Hh��5&^�� �6�[���64�0��k�S2�&���d2�g��b�"�!%ϥ�@���l�#_AC��������/�m�j�.�������HAq�fr��1�n�s�7���A�ZJu�vyd� ��Y߄^)߇}�R��6q�ބ_Y"|�5�ch�DT��Wo��s��-��Y���E�% KëY��R��!��L$Y�G��*�bz33ȡ����s>3�f~�$b�+���y(�7��9?S#�$�9l`���N�Ѱ~����A!��}���mgbN�����J���F������F`���)(�KL�R|���/M�H,�(Y������޸��t�,�e_msI>�ۡ������r`��л�#�������� �L���7���|]���I<�������\��l*%�Fe��\9�x1� IMT1$0�_�/�g��r�kL�?����,�=�q�IL�u^�P��Q��I��3��x �������J�]r�\`��BS�l�Cl�����|Y���LMK\h��R�y�2�������+4,g��D�2�Nw��jz���M2��Y�`W��>�Ŗ�
����d�m���)<�Κ�</e��p{}"��DW�9�Tn���V�]����(�^zY6^kϻ����͆ǩ��+Qb���'0p�([B�	)���)R��h#W�g�������0R�]8h�Ya�}�+=U,N6.e�T����f�N;5$�N��2H��c-1��;ޭ���ycAv�J�B��-�s���&{���xvF�Gi��%������3���V˰�I�^��D�m�顜Lv��*�=��	�pĦP]�/�޺GdU�X�� ��Ņ�6���ts�t|�N�k��+�N\�����8��*����8�BNl皘�g�02�٠�+T9��_�8�Dm�k�z�m ����2E�)�>f�s�J=HK{y��j�g��� �:ox6��*׬/���
q�8�Y�/m�N��w^`���j(T�,��mӅڢ[�+��S�a���㌅�����L�(�}��SWZPZ��*�*l".��G���j���~x�
P�ui�R|���~�bG�S�����ɀ�/s�6��2�d��ܡ�[��~����D�nMZ��(����s���¤/�/�v��Z�'�Κm��X�qM���H�)P���=�G�}&_�����e{o܄Rb�K,��E����6N}Fe��/�+s#[!�Z`j�o@@R��ΉO���qgC�o-Y��ki���gxR�DE#B�ƽ��n p �J��+\u�B7j�W�"P�k
r"G�ҼF�(�ϖWқvq��ғb���r��Y��G�}[��ۊ}�}0��V�$7��Xg�p4@t7���\�p2���[�G�˝[cݓ8�)��:�y�8ŧ&]U���H*R��l׾�2�ѯN�y���{����;q�����l=
�8�2VL9�y�&���Eq��q�[�?�G�$��������f2����0w�Q�Dk�z�ؘRe�iɣ�v��*�h$e�+E���٪�KB�� �{ =efD��5��O�d��\�K%�ld����03�˝�[_x�Y$X��؏�6�b�Qd��r$���6U4�_J�ån���S�fA�ܢ{�l�\3�R5��w@�tm�T!J|����"2�b�0`��4k��,E�=<�ե���c?,qQYI�R��fs��^�6�ckI���d�r+�\h���k�s?� !t��B�������f�e�U&5�o�q�B^C����ƀb��Pƶ�m�rNLpiE�VV�ď�iY�:��i�\a&�Y/�;m�N1��H�0������)h��W�<�El�g���K���f��И��@=ۄL�N�7�]�PzPs6sVF���1��
qu��(�[Z��M��:�c�� z�F�k/�S�l��'r�3�b�o.ʌ�!�n3d��֧�e|x�ˢ���gO�:$��Y��u��Nq;V�H�ʾ(eO��m�AA&7�V��~���@o�Б�����_L�ᛯw��l%u\�����fT"����®$���z����>�eC+@�������Gg^R�I�S�A��C�Q��c������<�]�ڳ�Jv�c�_&Ժ�%D �1{\�[W��2qu��z�դ�B���Ҳ���S|��&/gt�+�G|NJ]?J� g��P�5M��Z�W���NHX�Ce�|5x�$��-^J��L���HЬ G��d65�����%k���ׅ˨���3��#�X=w���6[z�*&��߾K6�׃i�����6޺��^�m���Q�v���H/��
k_���Vn]�G��Bv'����3`�b*@�K��@	�C��[���<�Q+%��3��d���o���Xu�ˇ������]���D�3�Gj¬fꪆ������=�4γ�s͂���]6��Z�
`- vH4�B*��� P�ϐj�Q����W��6�m��]�&.�s����DIq���B"��)��dI��M]��e�����>z�f�_���}4̲0[������L�t�*��8!�א�i���������2�Ƀ֖gbt=c�t�l��
~����u}���5�À]�%�ײ!� �i75"�Z���鼆�^�.�Hk�$J�yW�(wȿ�.�T�t��h����D�Y�!S=�.E�F�2
ID�%�I�PF.+M�	_�r���힘�b�{��Rx����B�$Q�o��˰���d�O�r? �'��BN����L��_�}���n�|��C��� ������:��u��.�H��cGb�(�7����Mj���1�ڈv�k�	��&m|����F^Md�M�"���[�%~G����-�'�2�=,�&Qh�bg��`\cd�2/���a6 ���~h!�(a��T�Ek�%s�IX�T��gM�Kȧ��j�TɠDд���X�YI���J0��Α+�ѹ:e'��S�jը�؍��o�:0.lWUsl�	�#��~{+h:��rvz*���c���N���I#� (����}u	+�)f�d�xu�'��[>��Qe��n�5m���T�!v�`Y�r�d孓Ox��C�.'-���� ���s��JNv�� ����
�=�����q�(�����6�t
���f�P~���V7�v��?����^&�mp�0�oh�1�|�9�K������Iw{�.zf@��7�3oN�̛���(!$V�{�훤?ʇ����QJ}k��w=U8� �h��mQhlҹ���\4�=N��r"��uM#�^R��W�o'��YJ��u��*���	A	��Sx����Og��*lý��|}A��^�Ϛņs�5�/G��nR���Y��?��t�5�e9r�{����8�l���!"èkaV�[a�?�;2ƶ���bl�^Y@Y/�CWI,p�&;�^8`��2K������,˔��#�O��^�]�U��{�kCW!��,���c�": X���CW�x��C#%F�J����`��)��"�u@����j��j�װu�(���(.�!�M]���X��D%�8j$n���n��1���7�A_�}P�ݜ�VX��jG�I��.��e�_�"��$�} d��E�����s���\(�;X ~/gl�ϳIc��|���y�(���)���b�,���ޒ���{!�
H���G{�X_�N�2�����Ȃ,���o�K����8���dv8L
V�t�T��Fg�蒔�x-�O�E�$p�y����4H���nb�r<�U�V�����﹎�L\��J�΄���W��3"Ȟ³����Jli�l7��Է��v�URxxN³����
��~4��c$��� U]��b:����|(ڲ����)rn3?R\�ȷ�>��_�����!ZE� J�a���5�V������[�k��`C���^{�M1��9���#�$;��H�������ޛ_����!�c$��鋦G���u�n�����e�Cׇē5P���i��`�E1f�~A�:�:4yc3����"C�N��9���J�����a����vO��꤮�R������?�DY��;�^8e\�3ٓ��1���r�ß�=2�`�(3�4�T�Z��n��,�Js���?����/�FZ�+9q5ڱ����j��B�#�4��B�&�kM�gXv^TcGP_���lR��2����Eb�Z��Z�m��rF���L-�{��\�R�=:W m�~M\J�)P�[E\;�I���.�vX�x�T���O�vכd�^�X�Lo����ݞߒ���6P��[��BG~��f�0��RqT"\�9���N���r�g��x�L����	��$�7Fh��mW���A�I��&�N�X^'C=�r���_�a�0S5�m^m�L���Yݓ��T��{W~̊��a"��<q�aE������nCT]U�4�
#�Y�v�jfz��0�Kǳfɧ��:���d�H gƧ�׫޵��3���sl��>��zy!��V��6�q~�� >�7po״���� ��6�]-�?�н��*]���3���ROR ����K��W;2\Q�6�<�c�OF�O�
/<A����>��tn��gK��n*��s��@cJ��f*e�!�f�b�|�C;ӮQt��T�>R{��1۫xd�^\��Z��\l��0(��mi���Rg�?4sH��8>����;)������ʢ{�\6�%D�ͮޅ�O������_˥aAΕz%'�\2� ����'�
N��*�u��DGM�R�����v�zF� ���}�	Ɩd���1�v����Q"��{0Y��g�"��r|MLߩ��'��.ж���X�Mh�a�X��ׂ�!^�Y��'�$a;�g>�!��]�+����i�@�t�����h.�rv���%߷R�4�v�w��w�|�A�d�)J�7�~�pp�ń-�)0�oS=���Az����Vm ����=
[Sc���±4��[7���TS�w�ʻy�����w,\�Z�覭���>��������^���TT`lr�~��;��KcLw�zK��c��4��&���W3:�"~�ؔ`��!����J̏��	��;}�;!h�p�5�.b3�X^"s�x��z�c#7�.�-Y�=�ܦ	c�0�!���X���H�5u/�\�^l�պ��Վ���GR��1�"=ֆX'p����UZᆓ��ՃF��ߐT	v��L���3��dY��f��=�
Mƪ��^��J���+����-%�����0�����U�s�ܫ;�ʚ�����eb��y9�4௓� ����щжSAC����A�*o�X���z+����:��b�P��#�x>�_ <�EVX�=*��7ً-��<s���`A�\�|��޽r��rV�*$��`����&Q�@d���a�z��� *�1��� ҆Mu{H������v��ٟH<I$5:4Y��F���o��B��=�{�|g*�"{���&_?�Ȩ^D�Ȱ߿�O���%l��,��i<��xĽjS��3�n	��]�+�ǢXXVC2�;{iS10���b��D���t/�3��D��5]�r���Vp�C��lso0��Ʌ ��A��'�*}M�����Q7ȏ��"ZN^��ǐ�r�AU7�����
�*%�T���A�	�\J����^ut>AAMx:u��.�I	�?�>N+�E����Z�ے�u��wfU�
̴ȟ_/�	ǐ�v�ܒ���!�?���������B�J���s�� ��G����]��I�M-7K����?A��Y`��JޟY��q�\ ��"Ƿfu���z�SdI�,k�T:yޛ���n�47����Ž�Wk�ƕҭ��nL���-9Ί)�k�U� �W޹)꒟NpD{V&�bM[�i;d�u��ϏBN�V!��"�}\}����-�����n����,���]=S��"�[���yh,�C��.��ƭ������.�[���F��J�*�.���@2�5$SK.�f���Z��Z�%��[
�?�%t桝ŝV+ᷪ�#ec�c����J�1�\�%�Gm�1R(gy,�)�\|t&��i��U����A���-A ?�dd�|���o#��v�l�Db�|�j��ԍz�^�������FL��	�D��(�yL�mh+��\�<���&(�`B�%�0�������hsfa�]�g���5�8���z�
�C9���!8AY�[�� ��j��#I.t'Ң*����J��J�_gyb(�X3�T�버���;���[Hf�����-6�l9�qY����A�HØ2����"�0�2Z�nU/�}GM�;��m1�:C��!�Kd��6�;fP��n��C���nĹ䟯�V`�)`���$�,P8�=�1"��+�x�1�$E��*��j<H���I��ո��d'+:�`��j����>u����'^���)0b.ʁk긲�d%�:���l�tn֯��Ij�<�<�%{-M�{BX�Fs�~>-�.f�b����C��>j<�X�82��m�;B�v�@���Y��ߵ-M�.0YS����I ���!UZ>(�u��y�7?�B/���kQ`�{��9��h�>�T�G������@�����V�3 �+PO�� -~؅ �@V~K��[��(�8(�W��i�$O׉N?�`�ب-�;��tq�5:�C*�4��o����_5x�+hΙ�<U��|�m&V���5~#e>,���j:�u1�����q:Ck�lC�G����m�a��j@���M僷�	Y&�wX*I����a�mRKj�SkX�����b�2���C5�~�}�tuIw&f|��p�{�"pO�6��%w���`�9��O�^�HzG�F���	Nn2s�ey��
6x/,#-G���=1���h�i#^���Ԣ�1I%�ƺf0����3�'���+;�d'M�rG��7d���