��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�%��bh���p}Î�C#u4����M�	N�s�$\�L��6u���jTЦ����X�����k>�G@�`��뉛>�����MIF�f__���>AN�(����.����G@h�]�%@ܥ������U���X|�m.G���Ɏ�`�����t�笮�9kW���auh�	oD���EV�<4�+㵻����#��X����6���l��˃��5Z��t�M�:a�3��_�pI���va�c5��j�N��l�PY����i�Ed �:�Wfb�.I���h�����H �'_�ŀ�
�/'��u:0AV��i8����Ev�?rڧ������ԭN�k��ɡ8vv�VĮi�j����W��o�.�E-_�Qiȸ �3��� 	0$�}�G��Fi�w&~K)�{];�x������h���&�abϚ���c��,.�|�<��:�яZ�F�m�9N����?�M�N�˅��D ���B��E���jy{��tpF=��L�g���X�(�����:�[�����zT=}A��=@Q5p���qp��)��
(Ԋ��M�U�JBQR���3�~��~�sNE�'��E����� &������߽c�y�Ju��c�S0o&��>�MT�^a>2D�4f��:� ����G�u�[hO�S� ,�[9Z�R2`p�i���L��%���2���%\6�[�a�h�\X�t�|��F;�Kry"^�+Ӵ�c徳�������c,M~�����y���m���=�v��'���s���u������*��:f��}������Fodi<�����S���	ߡ���م�Bd6�~�������w��hsd��pNu��.;������S�C��!v�c��4�F1�a�B��<���ʈ�R��{ȵFva�חY�7��'���sز�}c�.Q��"�R������E,-WD���x��(ǝ�M���n�^KN�Q��f�2����(&o�< �T�񻸋G�Y)�/�Rb0<=Q��θ����.1[��.�8��r
k5j#}~}�Q!�X^�������_wR�:0�|-�7���/��o�-$�ݛ��B����Zd��k�mx��K�\(�r�����x�����]%A��G�}U���zf	�D��Nx<j�9�Bq��y��8XM�D5n0��)�d3&�wɄo*�G��<e��TZY�$+��Ez�A/s\�>A6�H��tx��&�5�UT7��]b�~檕Կrx֎�ǣ�m	HW��| 2+yI�����~�*�������3�X�Ir;"(��8�#@�+�rу���C�o)M!J.��w^h�����w��2�5}z3S����:v�,�t3$���A@�n
h����
[vD$�(O�g`=@z���fb�k��y�Z�>eWi-�J���z~tI�C�Q��sͺe5�'떻}��cM��ux�"������i�ׂ4�^d���[׹z��ē9�����QlL�9�-�;@]��v��׼�������F�,��)(S7ĺ�A��c��+D;�A�����Vtτy$	������	s�mpQ�<���À����d��z�[����b��몣rj��pQ<���8�5-��کx�U�~�)0�Լ��f�������%���#����f�2ib#¨UF]s3� H#5h+h�(������:h~I.ɺ�K�b��*�L�(h�f��=|����x^r��o2�������b��ꫨ��J�۟����e��],پC���c��,
f�-8}���6�Y��V 5d\	O�K�7\a�\�?��>��γ�6w[%��"5ѳ5V���"�-a�e*u0�o�%�a��uJ��P4!�=h*,L<�;��a��(Z$b&