��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���tǐ-a�Z��e�l+�H�uW�Љ��Lk�p�@}5�[o�Hݤ|����j�{38��/qlW04\h"��=7P��2.��[��,~�����d���4�o��3%��!�:���&��G�Q5FJ���H�(�m���G	.��I�I�_���]�r(1��k��0��h�&��b��j�����Ǘ�g6Ԥ�f��*��9dS�>}᝟�i�C�C�����Ó�����RǬ�]�BU�����po7(gP�ݴrsе�7�V���~'�u�=��Y��<�(�;?}��Q2_�����-N6�R;SK8�n#1�d��0R*h%]6@�Kp� #�|�S�nj�C���� ,`�T��m7��O볻�ʗ���lUw�{�\�����pL����@��pEkR։��h�����,�Bf}'}'zM�����mm�=F���=
⮅��s��Z���
��=s���߇�Y��3Qm�R3��5�
�-~�f`��S������"��9k�?�@��M`�)�xE&�a����`s�:��`$�=J ��u"%�{E+)���j��%���!�I���Rnr�t����Ȍ�4L{��,Q�����l���GZ4V�~��/ 4�| �쮱|%��I�Υt��3�wRm�������"7�h#��F��Z����%F�sp���+V)�6��ڵ?�*�{?�kr�L���ciK�u"~m����
��D�i$S�FAe+��t�V ���!�����4qP�ި�&��ַ W���F_�j�	��p����4i��wK]���Vܭ��C$���Z}�)Wp�9E4@���7���}A�:h=�����:�4E=�e����;k���=��/�oY��;�,
��K �Uå�E@�����͈ϋ��o�@3%���X�l����ţO���ÐWH��� �#��Q5���v�a�����^>�g��,��^IV�k9hC��T����7d�����I"ư4w��Uti��<�g�݉C������� a������W��R���1,����.��>8 �&�b��Es�x>� ����8��@SEH�+� VSlRt���I�f:I@���uk��%)k����T�!l1ڝ���UjZo5*H��,ρ;NB�*�`F�����Rµ�ܵ7<��e$�G�$�\i2N0��˹�\�#��a>���VCn��hU^�oE��Th�F�����K��G�Ə7!:A�C{NN����Z��hڶ��G��⸃T
��eE���ׅ�WE�}(̭�Ke莲SV�Tj�J���&�!��_r�e�HPr(֌h�+'��ޣ�R����go}B���ty��Ye����aqB���$��6���V��MQq�[��-Cb�y�U�P�A�wz  ��Vl귄C�e|�v=�T�ў���J�x�S̀�ջ�v@�G]7h���P~}_�/Y�A�2heXsz%-2�l�� �Az7<.�M��Έ�Y���O�Xw����S
\	X�P�k��ƨ�Tt�i-�<�h���Cgo�	|.d��"DCPF�{K����᷵~pv�#�+9��j�w���Z_�҉�=�*�$���vc�J[Ϟ�"����积4hZ!�����t�	�����^~�xa���=1�4��-wQ8�L4Bs�W����]��sHW��z�ë��$��e�!��bbu1�	*��>��-��jv��*	�t�X_Q�$Y�����C�#j3 �� �(��*��=����]r_��d{���������}o5Y�m����l�Md���8�^�����b͠>Ҙ�<�}��7ݢ�Ɋ���\7�3R1�e�dJ��Ph�.|�g�gB5d�c�����t`�
��I7�\��v{������@^d�ltin��w^~RЫ�:��ж�p��a�t�~'l%U�<�ϙ���8#U������/���h+�A|;p��]����������#8�����9u�yQ�$%4ϟ*Me����צp�J`s�$n�a:~� ��g���%��8 �8�J���&��9�{0Hv���暾R�b=�K鉣#@;�~OR*#��U{��7�<yJ�!&�:4?���W���I���K�j�ҍ�f�"/U�1xF�=|%L
]�a@�ْ���tph��螑�Ou�{Z�W��΅临����Ա��"�|��@Q�����տ�AN`��I3]��0��x4JXCc�~�g��_���8C��l=��O��b7�P�e�Ӎr���PH~9�������ޥ*67� B�Sm("(��@2��"ŗ>^fO4:v1j�HF��*O����N�e`��Ftܻ�%b�����\EO~��Yw��ML�L�#q�V�:_�o�z��fq9�U���N�rr�H�WW�Yd���ڒp;e�󔌇@��9@���[߱�G�������-����o��.%ȗ��2�o�Hc�P��3=���k���Y՜V}�p�]ѭ��E����D�N��U#���ZXf֖s~�f�BL}o��<�p\�QKIB;�,��p�n�AEy|�`G6W}s4W)��b��B�`	���vOǔ����;1�*��]��Elȍ�$ ����Р����ljt%���r��]�(F�x����3�L�n0H`��I&d�&t�5«(3)�������n�_P�����d��(�sM��_��Au�w��p-�D�!�R�h�wg`N+���
�~}�+|>W���H��?�8�ej��՗�~T�˾�w��?oxb��d���K�^@�5Eřjf�ґ+�������X�S���OV'
}��9/ В��Mx�3f�����d��ݤ��Hq�+G�Xr7[d�Ǫo| ��%�u�H��ƈw*gvk,	!��Lރ�ő������հ���l��!����uuO��Zԅ{tE�`�`�,����H�����iN�8@��A\��T9_��Y����(�c���m[����ݢ���dl:�9<�YM�%���X��CA�����^qc�%���ip6ꆆ�!8���fߣ}Ri�H�B�we�$�f�1��[�_Ŕ�DVµ�U�y���W�up��"�?� D���߹���2��B�8��[E�33�����Q>7h��;H������-��jg�9�	��L�s!Z�j�/�~`[��0
�ڱE.�n�)+��jm��V�G���>a��s{_�?j|D�<)��x���
�rA�S����n�l�_�g������5���Ź�+�����#g?�_ƭ���p��4��s�U�{rq>�����z�s*UHE��Ŷ�yx�ȣ�$D=�U��G�k�����N=���[Y�
�uf�?.G��zn�<]�y�k�9�gP}��Q��xt��b��wo胫��7�C{�-- ���{n���z(��T�QS��-��%dx�$*��h�,�����]�LW��z�iZ8#�/�x+�9Ԓ��~Q�0F�X�.�_�>�B)��3�x��9��@$�!�'�so\(j�ø�|��YZk7����mI��������g�=dA$ض|�Q�^cQc�����nmp6�N��y��Ι N�9.DB猠f�w������*$e���4�b���fֆY�c>����6Kd���u$�h.Ai��0W������o��8�G,O��fר;�ܱ:�k�js��v�l�o�s���P��D���6�(�rN����J�Q'���=#��|��:Q�b ޘ�����vo�:_9S);�R}�Hv�\5�>�C����e �Y��i�"�#�k��sZP��?�?3c�MJq Կ�҆U>�Um�}JLs6V��r�IuM`��7��T���bꥅ�x��H� �Q��U�3"�M����3P\��E��f!`�,�5������e;1�⫞~�Y��O� �Qj�Rq5���1�3

��\�~��M����ߘ�\��1�-��_9ঘ$=���NZM��+�~�۝%3%���'���7 *� t�������9����|����ǅ3�8��ݒ���Y����k~�K��<��Xth498e�$i�i��W���	z% 37u.�zH���F��]в�B����	�-y�#������!��*�U����A�"7Y�F�� �H�;6+�b6&�z��n��ρ��a����1=���k��I�s-�#��-Ti������I�����d��	��gx7X�����b�iy8GDL�#���j�d�+���i��܌(�j*�;z���iT��!�`%d�c��e�)pC�^����V;�HK�|Er�9x1��A�a��M�0|��%,zy��/�1�Z�-'�(�y�Ы��;�n*>��\|�V˾6��8�:�K�=��*�I}ה�@ǥXN��Lߏ=P~�g9��<ʴ�&
]P�(�z��]~m{�w��rv�z���w�:_��3㩔1O`��3TÃq��c�8�SZtX���v�N\����a�"8����<t���΄�8�
�E����6Q:�$��� �mg+�d�����D{��[{}�C�~�j&&S#U4}�"��@�.���AnW����=
X�Y����!�嶤�ҫY��ދ�.�����
���\��Q�7��.Z闅Q�֬�&��qEO�hx�WB췷�?��JGѳ�<��{��Z򔺵���G<	����͌G����&:�N���e.�NC{��5����=��5&��L ,�ћ?A!�I*�=��^&D-F����Y�d����ݱG�QTY�B���9��N��!Rܥ�K���&қS,���rD��3��
T��Yt/KNx��F�q�XIdq��[ǧj����!6H�z������B�)�q~Q�����_T�:�Wǜ��rw~J�9C�1�<�5�B$��}O��g��á�����	wc����De�y���:�vɇ{�%�mE*\7�mkc��Eп��;N���餍����`!xzI&a,X�|�lfFP���q��e[듉ֳD��-+��,5h��j	�گ��EE�-�&*�E��`�����앚�tɏ�qO��_�
&b@��5@�2�,m������t���IcϻI��O���Kq���D}�G����y= ^'�c��ݔ@ô���U�ǥpDR�L��٣`{h��ܓ����K2|�zE���J�q#ҟy�@25���):�����yM!��\�+I�o�����f>��Zװ�1�lÙ�`��wL�,p5������y����
���[P�ؒ<O�N�E���}�ۂ��Z%�[f��G�y�