��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#���gXݤ��$pp�{�:�'k୸�i��8vY%�E��&�Р�r)M�8���RAW\1�Lˡb\�&\�*�^^i�ٍ��,���=JZ���������#��VDx�O���aK���%t���e})7��2SR�{�'��M�|�:��}^�~����r\(7I�ڝ�MZ���t{�o�dgd�dV�'����4W�1n&�!�e+�\u�5�_W�e�|9�+ƥ�4151��Ѻ�§x��e��g��ɤ��|^]��i�M��(�`Z� +�͉N	�2� :�
g��[����O�(�xL�n	_�!��m'R�U��k�zl<�Ym�sWE�1au�j�P"@�ۿ_ջ��XQՙ�$����z�[��0.�ryi-�b�ܷ�V��G*��7��AmC��ל۳���/4��9�c���ɥL�|{_�j`)^p�:�ק\��M�IIGGΐ��9����i�w �^:txi;PQ�~��1�R�+]��?g�l��J�hT֎��V�,�T5f֑ �KQ_��j�\K�$��zjr�z���鲽J�Y*@�ס�*�Y���u2���%����H�~��[d8}� TM4�l}b�le$���ʫ�5.<�M^��׈�NԘ�O���G@OI9��F����O|pŇ���7˙�ڪ��kh0��]��>�!N. �nc,y���XG0��5Y�LWU������qa�s��u���WsmS��;x[�Q�:Q�� B�����ūr\�w-�h�I3?y߽��,?��** "�'��^P墺dQ�_q��L���1:��m`�����fϩP���pAA�����!k�z��q(��G:���:z3��Ɩ@��%/�n��EP����V'h��UG��Y��h��O'^�׹�`g�� �y<�<�8��{G��s���6VN���l�G����喻Ӷ�e<���(Q> �3�Րطio)���d�'��z�k!�^���ف?�TD�9i�bE# =->$��{S��F=����4"��}�^�p�=(/��$i�"��{2y�ͼ5����вj��K|����؞e��u�ǧ�U6{�%��y�rU$*�&�'$���T^<��4�?gf���>�H@yZ��'�	�3I�qc��ݾ�{�ظa�ݵ�"�����@�6�
�0��z�_�::�{"�v@g��k�ڃ��<��n�9�j�0���� �0�NNl�xlUڀ��9\J}4��B/JᒲBb�4}��)��Fo>�-�<]�k��$W���w���Y�DR����X}�IG�lrrj�S��ͿLl�r��s��'2��c>xpH���	m�	/ǎ=2�]T7�$�Gm�x�e*^2��]K؜z{eM�e�im	!T����$�ӆ��<C8$�6�����;� �-,7~u�e0%��R����j2��5�٣l���_���e�+��n�?�����U�$����7&#�7�\��ӧ���c�'�8{���I��@�W�C�b�f-�|"��4����Q�hm�e��zQhţ��qPU���W.�5 /�x�P��ت�H2�H����	?%��Ѓ1.QQ��}����`��ZP!f��&h���	�j��s;�Β�2�����xl"9yp>�q����Fu��f�P!���nڮ���}	`�+�X���������6� ��!Ś�l[�2)�D3���T�|* .���-�N�q�;T@�|��s�!�����`%9�.TG6p,[�'�+|�@+_Zl���w\�5u�Dh�F2܌^N.ly��I-�\�\s�B�Ε.!��Z��(euo�q��o��D@A�w�*mS�e��� ��Ea��pX^�pD��s�<����n 9�B���gg�߿�wNI�3� oj����[[A���݅�[�0�M S�T�ܸ���`�q��@�dLu1^��<�� 5�A�\ڳ�6����hj�[�F/<�]ې yg���oh�oBi_ێ���G��O��6M�|�
�ն_8l���o��z��\�Be<w	Hp��m-�u�8�|\�k����n!����w�`lâ&j�%ЪDk��������^�D�s�ϴʝ"���%�	c����=�"�����/,��:^�����en�T~*�f=��9靦�z:)rf��~i/��g����>��K����-N�-��K���2�+(:M�bYת)S0��1�dE<��V��g��[㢑DʑC���9��=� ɍ�c�K�綮D</�̙�4:� B��sNE~�vD[#!���Ь��h�6�9Qӑ]� ������s	�E�u*��WR�}&Fw��wEۮJ|�|͕��%��+����T�5����R�
2����h�z,5��m��vX��G�N�����e�0"\Fy|��-���t���Nz���2�j�Z��`�B۾??{Z}jb���P׋O々�7���o��l��:��a��G*�h.��3	q2���ݳ����kL��	iw�|�?H���d �!kwٕIՇ�;����Ak��M��NPXT	滽p^�������f��*ג7�jP(��n�m�*�8��P)�(�':���Y��Z�`MI6�{���T����
�W[X�u#�h��&,n��
c��o,`j����1��k[������ưj˓ ����M���9�l�h�CL���5ZP��*�V��D����Z�g����Sw������FScE�f���_��qY
rC�Y��S�
�bm�+�B�m7X�{�aq��p�|�o��F���a.��p ʠEFv�ϡ��jl�7��U�w%������	;\p������"ۏ~�հ k:�Yoq=��O״��o��|0#�S����w��Oғ��㸿;9W�u��Y���0z���(���1_ı�27�����ah�q�'A������b$�(�󌈃{��T���~Kѯ�dɆ�=���fiH��a/�`�i"���W��N���a��W��`�\��K��~v<B*��-�������^�r'=u�;�eq���4y�aT��t��ႁw��ԍ�r�����d��"��3B��?a��)���L��w�}�=�����Y�Ø ��TҼ��M���)���w��h�*������v
�ndj��F=a
���߱�GS��b�U.��f�����A��Y�ba��)W��a��<��c�d m�dƙ�t�r�q�v��m�?�CD-�0�r�c��D��c�:��ڔ�].�?�9��_*b�;A�>E��hv�p�i��	�G�����d�H��� ���_ �՜3W�!σ�$G��7A��M|F{�d����ǅ>�(g���vI�nr��˕S<~φ����:���@���\�òq���ކV���=�J.|�?l�=cȖ���iS����tV��)1��p�g����zhW[�s���.�0I"��������Y��R���g��\z�����Z�#�t6;�i^��L�~z��»p�L�&pO�M>�,����ɂ�Lb:��r�� ��Pҏg�yŏ�0�_<
�N��F����f����&�=F	�n���D=���\=����-�C�~曋 ��=H�ސKtL���=DAԹ(:���gc���v 	��|n�����H�L�����r���<Kx��t:�Ҝ��F:	6��
��ט�}އ��wb6-���ɻ9T3)=#�3�pП�F���)���%{,8~�k��]���`V�5�-;���s�C
i�d)�2�'I~!��
��{g�k�繵���N�٬���,-ej�=C�
	=2ۄ�¯N�W��A�t@hi���q�2)��3�tx���k�*�bЪ�Z*��_�i�����+��(wL����/z���6E)H����3{�s�x�݉��o�
����T@5�q�8�nxEN�!����4�<�2Fy���WZ.���t?�������[��i�H�W��ٔ�G�Sԋ��[&�����V��F��0��K��`�#������{>�X��H��%җ�塓�Qі#cLץUx E#e��.nb�˹�K�?��ZY�a}��+���a�D�;5�h��c��1Z�e���>�U�x�!{�2Y

L!Yŕy��c�|C�⑨p<��,���K��j����3s�X˽��R+��X���_5M�U./�hv\�D��8��#_ZSX�YEs�����\��T����Q�����^��NB��D���.�E��\�qiv�C0١��E���Ȅ��O0I��p�l�P`[���� �w�D\w�} �	k\Y�R``�HZ����Tb��O�b 
U�2=��	w�>Y�I������ZG;�r���H�~��W� �7�:��K��F�9+k���Td&K���'���lvrZ	B�f��h$�����'�0���zXML1揻�B��(v��:�C���	�������[�@�&�_��Z=��8h��)�',�� �TR�F��2O��0�3�*��O��r�G<�����G�_L~�� aLU|��VF J�^j��\��jW۾��羲���l��l����\3�7��>C˷���[y��ז��WP7�р15���-o���I�"������7G2�?�W{�\�g�4KRFHЛ�X�H�J+��Y��0����?+q*��d���)wh�qK�f��n��$d%���O�28;�hi�:�P@�_��pN-4�L�]�����{2�Ҙ�k�Ts��_I9�_�vZy�d��/O��nъ��Ĉ,� ��~���/o K�������&'0l~����L;��뜲�A5���~xϚ��y���)�L�yXΒ��$X�C�V"'5#��YG��"����W2�4����Q�	*g8PwuID��I˪�#&�k��)BȐ��p�鼖5��!�`"���H�M�����:&9io�a��'i��/C\8e���5��Am�r}O�"B5ʚ3���W�r����;Ksl���ǋe�G0z���$G+;j�q���l�� �c
��y��