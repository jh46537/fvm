��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ� g�I��Jw=���c#hN�j(r�y��l��έJݬn�1�Hs�P�fy:�����gl�����y���NE���J�S���r�B"�?�a]xD>�G��,��#�ô��h J��"|6e���${oT����f�L��-������L�;٦���O��0q_����We�f����@��52?m[�-oZKc_��*����)�fA��7���p1��Z����C��u�,�$�-�8��z�̤��QOS�i�2���y14�W��E��B�l�St)��܁tᤌ�6����c�gO8��q]�"!���Pg��p������w0vwM"���I�T�h���[�b�vӤ[\�c��-x�X�����r��X��4�:�:?:�4è�Q� %�X�%�-�U�a&��qJ���M�C���ߕҚ)���7J�H��=E���������������[&R@�eD1>����z�����l��-7��t�=��7l�ۙ�e��=M�➸�ԫ���C7���%�q�/�d�މD�C�
-�Eh�������Tt�˝���Txѱ��7�ӹ�f��}o	�h���`��o��Q<��ns�Ȣi���;3�	d���L����׮A��8�꼴K�c�h"���`9���w����r?���-���IV`z�x�G�w��w�Y��rj#�C�30�)W�&Ⲅ�΃�W~���nO'�Y��	(���y�����Xh�m:)q	��ȼ�(n�E�[M�a��f��#��e8@:�&�"�4�K�Pv��3l�X�+�PJ�ܥ��P���J�	K��O����}Ҍ���cT����4�eB�#�� %�{����/�i�.�|�Bap��U�L0{���hn�bl	����`"���A8�2sL�>���1>�D��;��	�����+i����ϒ�@9��Du{���z�� z����3��U��߯Z�v�a6�a=���l�Uv���"ܒ���K�
 r�Y`���}�Jo�a��8�<b������o�[���:�f4�����6r��5)f5�P%*�b,�����x��cF���kȖ��i�yZ�Qhr�[�r�_�'�&�
���;�^��Y����B�k�~��SS����������}T��'l�A�P���^U����[kg[ߟna��$����5�]|�	����p�h/v&w,YQ����;�\_�iZ*�Z�R��j�p2�s���K���{��*�i_�_��n�������@����e�~H�*4��jY�����N.B�s�P�*v�.�,H_$����t��DO&�	�,�C/�޲h���>)��W|�����s%b��&�Q�5�7U[R�n�/�|��k'_ ���c����=��a��!P���f��-�N�4v�}Ȯي����H4�[�G>$�f��Ayw�Y7jCsɌET���DB��Ck��	[<HS�oVӇ� lR����J�i�3y�����f�]?�m��u�ܬ������>��Ld%�#�T*�E�᠊L6j��\�G��L���uw�P�m�C'���,��u'��������4
	�aΩ��+td��y�(�!Ci� <?O ,V�#�����v=q�%�uiѣ\�����}�߀�NU���7?p�s~4ʞ�D���=���C�