��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzG&jI�#�a�_{�3*�
#�%��F���+ٸ� ��E��K<D��NS�Z(��e�8�6� <�ESO��r� �>� )��N�*}-�m��>�	�$�z�t�H��eR<�A͛ve>�3�_P��D��'E�;�������Yf�Bg��.�w��_o_��TT��'��0'P���<�<8���b�������OH�3v!/��/;4�p�{4:I(��~��Q7�#�:���%��8Z�n
�D���ٙ��Er��$&�P*�d�#�6:� J)��7�/��g_�!��𝯴�O���r�����Iݼ�Mj'�D�P} ҆b~���}��m�hS�[���sJ��6S��e1���%���ŇTr�R
�h��&���A�E�meTU'U�q��
5���L@�}� s��R���Іi�G\%]��q����t�u�wQT��\�CdN���(/uu�n2Z����$(�`��(�����T-����c��U��f#�V=�Q��/�zz������0�K1؛�Fv���h����0� ����P�Z��H2v���Մ8Oʸ�����ʛL�6��٩ȥ=p����!��->qB����7ӣ%zC@sM���M�U���S?/0�9[9Z~Ex�t�ð�Cd&��H�D�K`��!�YHy~��k��Hg!���t��:�▢LAP��W4�
�!��Le
#bk�`���qY�"c�m�����`ZhJ�NJT'b]��	�#�� m/eJ��eͷt���}d��f�dy"=k&���d��r.�5_�o!��`"��LUu�.`���q�_>�F��{�nmg5����l\�Fؾ�`�v��]J���&b%�5��Ϥn3M�ʂ�����4 ���S+�FM��,�C�"�JK�FB�@�iɮ�T���������3�K�/Q�7>;�K�7�t��k���%��v;efI�mf�����&4�=S��i��\�~@f#