��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	�����'Ri�g��
�&v�/�'&r�j�U��
?��A���Hg���Ѥ#��3&;��V���9�C�}-	����-�+��%���aa�[�>�;_ĭW"�<`2,���E�0��P����xs?�l�M%����N��������zj����dſ��}G�����y��"ċ+Ϋ"I��|:��8r�<�d���s����%���]���?�x�;�}^��P�&^)l�Q���(k�t��0w_ͦ��F��̍���8L�������x#�K>�7�N�{:�8�9��f�ܫ�ܾ_n�$2V?�������hIw�j<8xڀ��Z��u�s^SJ9�|i���$�>"�\���?�r�t�zCi��Q��5�����N�^���M�S�!�%N9��f�(
ɀbv���3��NJ�7��Q�ˍ�(%�����V9\/����>���B|����T28#"�YpI�k���9�e����v��za��7&���Eh-�Qg��x��k  Ɏ��\˒ŚY��t�c�-��ƃ �����q��y��b����$nf�7�S��lȷ%ZT@qj����z�bL�b�h���Ǳp�o�1���P%��RD'����vyD鋤]RV����I��R���i����nnP��ؕB�R=����U@N��}�E$"3�$�E����>�[�k�1Z�&�P�r�B2���K	��s�W���X���H���f���Va�.[�.Wa�K� ��X�H��$��EԻ���>,'u��B�W+0҉���^b׉J�~�����`�O�I����?�t����Ȯǃ7?M��V��fm� Fm>�8(N�GWh¦8<5d�U��N@j!q�p��2}ಔ��!D��8����y��r��dҥ�;K�d�����H��uV����E����b�.���ˁ�!K|��sOx	��s��-�7f��O�:�qkZr�#ى�}��2�Q�5�����e�{����3F`���E��m��߽_j�Ҵ¦�Fy�@�H�b��.Rw%9���$�)
a��q0֬Z�)Y��3"}u��c��J�L�H����Qس������;��v2��v���^�t���{܌�<���R��[����y$��V���v�p}� tCjw�ދ\�o��A�j(]�'���T^1����:$�tESE}i���9&Xt������³&�	xݤ0�F���#��� �*(������-��ɉX �cBF�Č4��?�=�V�i�>�C�Ct-��Q���F����LI�b�E6-�xW,l�^����F�·�:�V�|����XY=��T�ȅ(�����_N�g��=���Cg��4F�C8�m �9���ΰ�������o�0
�oz(X��V���1q0�p�k�������pwࣰ4kO; LI5������m�^S�tv�e���i��h%��]k��i�R���*&Z����/�ɰ`xƎ0�厁񆊷Ѐ} ��1ͰlI�\��M��3��la�yT���!��.������w���HQ革�QG�0F�y1��w����\�Y)�8�����̇�ac�Q���B���������<����?�ׁ�f%����Q�A���1���'mL��Wj�'����^[�H�e���٠�k:�C쳠u��䯥�m���M�1X"G
��V0�o�cOBg�����W����Ѥ��Z4p{�݃3#B�o�Q��$�q��Ye����i	�(����8���n+���>�9t�8Q���˽�5��˴����J~-��rp�?��H3�a#-�E �Ƿ�+RJ���໽�/� �;}�8/�m�%�o��
�t���˧AZK):9ȏ��D�å��5TQ�I�Ð�\���a�o{��v��bh�����7��c�Y��Ԭ]�����E����$��D������X�X��jxs��m��&ї	x���%#�%#��̓�)��m"��S���RxU�/_�D��5E����w�닩��WT7��p�{[��e/"��p��3��IHy#:s����`��Iy�v��;3f��.K6�.�A�{��TN�y'F�d��������3Q(?���#�c�>�F���&A�~n��s��<vg�ΈZ�Y�]H�8�;f������ѳ��D�f�����,���n����R��4��[N���:4v��fo�8U��Z�1�Q����0��
ە��@g�+g	�u�=�c��B��W�3�h�2ť0��@x��\��dk��o?�-R����I�L��5��������]�zI9i82�x��^e"8S+C�D�RS6�("��B��\�C[��$���ِ�)���-2�������̩�:]D�}����y{��2 ���\��'�8���UEx�H�{ԾxYN6�=*�ݲ���c��)�m��~�n]�N/ײ�����A%��\�!Y��N�z.̈́e�Z	!�P�vr����<�ru�G�{�Y���,���f�ez��b���{���k��cS�*�QR�
�A7Ҧw�'���s�� 7օ�~G��pp��12�t�ƛ�u��������(�S���y>��_�XP�;K���;�I��Qa
���/�]0��/C�E>�u�����"�臼qE�V������Arjmgy��E;@�V��F��%�����$"/sr�2qR:���J��x!�޽� �d]�,�*)6#�!	�9��>�%���BS�]���I�x��(��-�L��6�;��d�*,�L~�4�P,�Mwi��e~�7�>_/�P�6�n�X�<�2�6���[��HS8�Z�7�� ��~e%���S�=ĸ�
mѴĠ�,y�����^p6����^�H%xcL���u��a�ll,Уo�t��
��4w����8��f�q'�>�pK��q̚�K6x�I:#L��J#FJ����LZdR�*
��2B|Ajy!��J{�^D��7�H�Db�"�:X|h>:9p����Vq�kvJ6��S�v�#n֥%�`�}���v�,\V�N���͜%��g��l�#Y��DK�����<5�����Cϡp�p��9ȯ7U�����*�����Uʇ@�\���1i��Њ@�w'� �]p+���`�ٌ�4��.�p�W�iH��&W�Q9�n}����.�q��xQ_�F���f�Uy��Vb�/a-�m��
�鮘̍�r� *������\T(�6�SV'�e\c\�Ҁ��Z ���}�%]�	N�M�Wa���$�m�~7p~�G�tI��h���P���B�t��u٣��U	vF��2U �)�����W��������z�	F$'u:�x��R�*�z{�c�!m	�􂗼n���'�xf:���a��C�E��y�N�n�a��y���P;H�Aes1H�2¤y�[�k���t���F�lsx���!�m�Q�;S��F�ZCH;K�FM�i��F!c��a�a�Q��'[[%��N��Z�$b���Z�c�g���j ��`[��ժ^�U����4�OB� +S]�!��k��m����҃��x-��s[�dԶ@���@�@��lES
�c�~Z����{�i]�Ȥ�Y)nV������Z�4�І(�� �
E��^D��~VF�9
����C�����_-��K
d֗�Qw���D(�4���v؅�M��:Ŝǂ\!=�pPU"5�.��κ;/�M��5�
/�A^��̨3}��#(~1%u=qT6���jِU�Y{��f*�/a�Q�PJR:�:u4��1���`����+K3D3�QZ>�R�r6���[�f�A(Ε҂�:8����720�6\Ҭ��x��i~c�!��5x�6CP~�ǿ��i��éA<Q�k�㸋�P+�Ն�X�\���\��` �P�~��Y�s3	1����Y�n��O�7�=��؍��0�����S,���mU�b��e��ڶ=3��[;⹱���G�K}��Ia��%��<b���c���@��]��GgF*U��i͔�,;����yo����E��G&1ԱK���E���K���'�3I|�']����à{I��b��<�sѣqܺCM���s+�( ���n�6xs
�VxD�/p9^�b�:v΀��x�X!(�q5��ay�M���mH9E��Z:��yr���)���u�uL!�&��4��e�6�_:V��M�u�v��S2�� ���r!� �E�#S�\`��W{�"z�3y@f^�T5re@��Gt���[e�.�}�؅���-�3�^��uZK
sOd�u3HwPS5w���b�Ou~�,��k�Q[�O���O��)���m��2�
(=𽄴L�|.9�mW)7���>�m��TK�T�qǏ��w��"=9�3��z���2"��B̵�`B@J��0��g�h2�a�u�a��xTce�,_������Jt���G���
���4;��2S9ƌ��]��T���