��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)���LB�o��Q��'iT��OH�� ����d�;c��e��+>r(M��5��q�Kx��p��i@��F{\�@���
����۵� k[�+����N榜 �^ �ق�{�h ��=��YYB��Y�"U'�V̅�ϻE�ݕ@�v\2E[b�pM3\��P���cΞY��׎���a!�]`��$Sk�s�ͱ2�E��1�[�����5dFV|��6$�>>W��=;��qf�O��0ˀ�K��JZ du�p���ӶטE���>���KH��.ޅa:D����^�{Ɠ��=�ST���W�K��F�ᥗ�pK���(�����ac��c��J&����1g������,{=rб����y�ϡ������?�k��a�(3�[�L�mP������M�n��g�S�a�r4J./b���IE���ހ���� P\� ���[��!�K2)�SC�]&�>��S�a�+�p
���n����7d4�Ug� �ӎ��
N��Uڪ�,�r��%�I�U��]�%��P��.3L��p�sy>:���Ōz�]�$�]1P�9��9�c��5~���_�h=�GӤ~����[`N��#͊�C@������t���"78*���ZԆ�����!�5w8�8��p�y@ˤ}n�ݒ���%^��%!:��,%T+"����R���d�֟��{$���z�k����s"�r8��{%q�L��#��Q�+cu�崞��Ss��2��^�e�F�dmΘV�ǔ�A[A�gO��E��0C4�W�@'x�lZ{���+s(�l3�WZ��π#�4��Q��
��
%�R�]���K�N-�7��,c�93��;�~c�4�Ϋ����U��x����Z*�|�����D{Ò�X��͒/9_�ay���l@ �ܧ!�S��i��������37aA�zB���
�7 ��4zYؤ���d�����~�L�D7�8��D���!B�v�ZJc��?��_��:�	�3ڌP��%" �υ���@(͚������
�?�b�La�Φc}��9���"禖	fr�G$�_唟�'�l���o�=���r�-=�������>.D��}a��u�{����c���@����J+�� �
�P����������4�]�*(�K�K�`����E��%G�w�C��	��ki
��^��Q����kDa+z%�_�x��BO	��;����/�	�V��/�#Zc�����+,� R����F��m ,���1�_R\�c:e����Qi�营]~%�O�+�ި}8�y���N7^�����?O��Kv�;�)�"h]�v�Na |c8u�n�P��7JU���%(�n�g3��a����ͼb ��^|G�3\�is�GF��=�QU����:A���4-�9��os�Gt��F��n�d��8�E��j�Ћ�Mj�NDS��_�F�V��St�s�&޽�|o%��~��e_��dVù�H���
�mnX)	J��R"[�H���.�I�4[�C�\�%������M
F2|�j ��h6��}ȣCw�� N�-��d�c��U�/U���7�X���v���5a:Mv^��689 ���莙�EO�	1�|�9��F�zzN��2����f��l��P%�L��.G7����N�`ykE������N�W�zbs٪O������b,`��J��D7�V����>3l&�WX^�ǹ����Bǲ�`��&���+�F�����O<�@Y��/<=��|��:�1$�䰋�8�?�Xim�7b�7f�	'[�78�'"�'_�����9�6���ˇH���0&�.�FB�&��#���H� �+p�sA�.� ��Φߕ�$��uF�MK+�c�d_����y�f�8�}C	��u{����-t���s��g��b�T���ȇ�h�%�cY�B��m�,g��v =�|u�	tߟ;kR��ι�a�d��BQ��Tg�ص_�s2q���I7�������3^>���R������/�~�Ŧ��!�@A�{md�A�򳟹�/ }���G�U=HV�t�º1��V�Rs�|q"����k$��%�u����g����6L�ڝ]������� e�p(����$J�1o=������h�V��'�
�(2�����1�Ïh�yn-ݡ�yr$�����k�u~m��f�����o��*��a��SR�a�%�M�8d|V���[.:ʆ�M�����v*��I��Q���~�1$«w�x�@����ߞ�sw(T�﹛=W��������9�q�޻�4ؾ����#m�'?� �z2y		�xzn������[�������A�;�T�Q��F����F��Bž�Br0����y�֑*L6�>Ye�����������@���DC��L	�	��Um���E}	S`�3~|�,��B$�|��k�lr_t���-t|N�$�b��d#gu��%�h2*�(�z�݂����&,0�#���P�k��޷D\1������2�C�pS�AN �����%�WF9�J�2�����O���W��?�2;�a��A��z��έ`��뭗֎'�3�;4e�;�z/�7��s�r	��X{�hF�mb��s�KA,��YB��q��!˲��`�=y�^�n}P����m��8:��ۦh�ԧ�L�sKwK�4�'9�J��ےd��S��� ��O���M�1������QO%k$�Ci�o9�䓳�i�U�L�/T8��B���Ƙ�'W�:���Q� �Zﵸ#��Ա�|!�3R�:?#��:Q5�/�Ɛ��������+2�._?Hc[�4:���>��w�4an�m X��ڒn>�z�ݹ�P�0����M�<d���A�G�ou��;�h��I��y �O�h�L��~bfe�Vl�- ̪2�&2�qg�C�V��hN���K�N,b���FtK7_����>	�y��P���;�"�o�t:���0�]u������r"V�!��*�.��]yX�����Y��@vjm���Cm��|J���K��\�(`��W,+�,#�v��F�y�����M�cǀ��l��J[�P2�ڣ�˄�������;Ȥ��fo��ߑ��7.WV�2���-�����1���l�:v
��@�k��L�8��l!g�Tg�T4E�#��L�U�hT���Kbr�WA`;�1��7�_*[)�8y����#ƠSX�����"�qL� c��s�?��?���V����U2�ýG�Z���l�;�}��3�{��~�W*0C�f�Q�U�-Ʊ�����ñ7<�0MfG҆lZ����aKIu�`i8<Ӳp�\�?�-`>��" K�y�'1m��W�.V?��sk��y�^�=a�v���f &��y�q���H�IɄ��<e��=�[�q5t���!���c���������6ݘʬ�$��V2Bw���u�55�4��P���x�(�$0[q� !��)�O����QM"7��d�u*$�Ssr�<�&��W�aD��.mkWV .�a�������P�>xo�c{����X=���G��\��"VF�.?� ϰ�]?(CCް&��u|򝄦$ݒ!�YZ%����B ��oy�V[���|ƅ)��U8M7ו$b�'Ĳ�$�~j
J��=��@�'�_O�i/Y=i�&��&���?�8��n}���4(���)�-��.V �CswtYC��O;u,H���i���y;��8	��Hy?T��04��З!���'b�;j��2p�|6�|���S1��������:�G[Y��� ��J�!Η��Ϩ�J�4�5������욭SA����[�:�6��S�PI���p���R���t��h��VP�:�R^�M���������q��r��';ɪ}���;���X�z�˩��]668 V:?G��̓�]T1O�����J�'@��1�Jʖ]7JD�ǮDp*p�?#9�;��_(�T�~:��㚓A���S��7��=��|�bJ�@�>9�غ.�T�!@V�>Z��B3�%��{Z(f���<ET����;\|\����n��'sF�kوr��"�%�Wz�XzT?�Ek���]��ΨL���,���hJ�&ުd�;k?��#bA��BH ���>�ꌝo���[
�N�y�b�'�0cI4��6��8k�1���#Ix�o�Y��]H��ʨ�QL�2^�hS�`�.���vD0��#%�8��Ò��/��m>0��a�V��������;�PΓ�-X���4]IJ�g�zKvc��ˁ6_�{ X���=eu�9{��5����$S�.�V��gč�%׭�M,>���VF<��Ew�|�3�#U�{��J=��&纅��h+����_���a�f�Ӄ����"�XKs���i��;4G�M �U��y�Yw��8�!����E��[�HA1n/���8 l!.�0`�_�)���\>_��x�63�H!O�An��<a~cA܉�U�>*��w�1�y�gZv��y�>���o9(��v2����%U#4,tmum�����c���#���sv���-�rGjAx9��°7��d������k�J��^`��q�e�(��s�����a_Ω}w�Cc��6�3��w�\K�*㺗�������]���И!�e@�@:�d�-�V�"M�9(��5��Ґ(��c��Lm�*����)6�zt�t���/�+##��%��:�(G�(�#Em�Aͨ��R0���v���VN����T|}�C�����?{�[��\�jH�-Mb����d���!+(;Y!O�_�W���A}�^|���I�8���C��x&m���ߺfL�Ч� �UM���^��A���7ύsu8xl\��	bY4�����#��75P�o�����)��YM�t�^t�a[Q�ke�(Y��3`e�T}���E�[V�d�$�??��6n�E<��;x�P]���Б@#�Q_�w�M�!tkW��"}L��Rd�߶��S�}&�-�A�Jcp�c�8,�2/���|p��G����K�ekC��a�%:�$C����5�����bh:�-��n�Z�g��t�O����*e|.j�Ø(]I��r�De�ȓ���+}zx���D�ףv�6y�I(�y�bH��B)ь ��6y��}�X1wM�5ԛk5��;l�Β\�ab.�'�k^�yT�ɝ�҇_�n����h<mOW:FhA�aI������/�f���Tj�[8W,xk\��$i&A��<�J�3{+k$.�1昿�F.%�S,KYoLq��>'��.R�'﨧�[6�'�BG������>x��?�S����)���nû��9�tUլ��O��f�=<�K�ŋ����_qo��T��T���eI*���f�f���C�^K�^dv����]9�Dh���Xj�,���O��ǐ���n3%<�4�V��Q���籀�]�4��^oI�̕Q�߼�%�^Z�k.�7:��\���t�9� B�K�O�.����L��n���Q��p���0���U� �פ�H�#�z�{N۰���j�=��j#�$������|�h�8�\G%���|2A�j#٠�cEO��]c�u�:hZ�V�� f\i
�����sO�_oL�U����T$Bm�&�D��Րgݫi��`�+��{u�=��2��<F�X(�A�����X���uq��BEu�e������6K}(��O�������;�aj(��
�]WAYu��ae/�ߥ�e}bg ���7y^�A���I����,�Ude�Ό�2k�usiN�%k��<?��#�&�P��U��%(jḆ��� �������U=�>���
����w�C��[?�@��P ��O��%p�7��N���[�&ƝQ�D��>xA�6_�}�I �Έca�N�nk�=33���3W]�y,��T����������~�k:'��uB��Y�S��o�k��o��Y�� ���ړ�
�]"R9&���Vl;�}��s*�!U/v6·Օ@����5E�\$rK�na.�;�/�p��@����3��+��\o���v+?=b�>׭���!X�S��@���H.�(���"���U�l�ŏ��w����YGc`�\}�"��*�y}���V��Z�M��n���L��K,�9zlűb�Xz�4%�1 xt��D�kT׊��O�P,��f������ªQ{�W���g�eX��{
�>r�X�I���d��-��>�v��iIY��Z�D���%���z�~�(���& GVx�-���W~e��EM����_!:,t��Z�Ӧmt��:c��Sm�ݬ��Ze��2��T��D���7�Y�Q7�f�c� NR�/�G��w������J;]��sF����P����V����RIT���M�<J�I>!bs@՘GNyn�q6oŎ�I���}g�eZ�`6��V��()xƀ{��\GQC�K|w[p^�%J�eӧ6��m)n[�eJq����Ǟ�Gy���#�p�m'/c��e���j���eto�����Bk�XyM����߂:���sk@2i!i0�����أ����_���L���'I.��)��κ��RE#J]h�\5�'�K��*_��(�+A�*��u)'�xe"���Wwl�Hq�g�NM/\�e��)a_�(L���r��˰A�򏔎M,�͕�o�;6�r�,֍չY���Q��W:}���SQ��#�n�R��=n�R�ru�`v�|�v�,/��jRV[zM|;zp^����)���^.R�Pd�(ҥ�"���G �����^a�ϲfw����T ��"�6�Ǝ�"V�����(S4;W���g˧�Қx�� �B����!��J�4�^��b�Ӈri�:��$]9_5IH��<s��:�_�G��oL�޴Y�Vp*ZWFL2w� �%���6�%�t���+���<�C�Z�U�$����yW���d������A^�W)���T Z�����\��5\�dإ1Ü%W�f�ĬH���P]���"���NӺ�	Q��%,���.�=�5d���E�b�=�a6��ĺNς���bMFB��3���dX��}a��;�Z�/���/ߓ�cXV��s������s�0ԓ��l��
� ��"t��;9s�q�@�mU�e`ť1�'&��+(��ąE؝��� �@M�E$%NJ5������v�L��.v{�^�V�r5��N�t�;B��O:�O�� :e�)_YDw6�~.���HIsY ��*1=�:ʈ�f��hܷ�_�l�1�	�ĝ��FZhN��5�M��Ľ�o7��"��e�K�C�eT�Ψ2�}�H2vڊ�K��"J��:����i�͹rQw{�n<-�q˼����糕	�$�op�eL�D��O�c�
t�0I��6���ӓO��������D�Tg��"䕹Go5m?&�ۭ1Z�/���"�n�c#heM�IF�T�b�Ds`��qћ��9D��b���W�L��r٢GSٹ�_�|��JB�6c^�P�����m��4p{Ɨ��q�h���g-��/H"B`�ĞK�u9�D��B9ǽ=,Uߣ�r_�?ϥ�,!3{��_�*�|��@4n���H�_��ESO��@R�Ax�=A}����gͱ_�=�A)p��k$�J3^gd�i���*��,����>ײ�#�Fi}����[�JA�O�4\"/	��G�=��ڞ���7�oJ�����_M�?jd��;�%jo�i�F� v�qn!�C��fZ,�𶢓���� ~:� �\ST��VOM�i�ⵅ���G����L�w�17�m/��U�O�����8��S�o�Dlk�9	�D&6�J�)]ؾ�$���<�T�fK:�Ш����*���<E��������9��9�F|\�����,ILa�-�i��q%�����\v��Bږ���<���%�`���|�?wU~�X*NuA��0PR,�cdZ�tK���	H�a�f�9Z[�o���-��,�Ƈ�E��h�G�ï��Ϯ�����1�����p�fO����-@�Ufr�����~Zl�)������z֘���e��ΔM�E��
�?�S "Rl舘����*�~�j7H8(�	���!�����W���M�
�)Sq(p�yS����z=��`Bp�
K��� �I*��Ew�L�x�����O�<0HX���'��k�q?j��b��-�O	�[b�A�E�
���/m��`�����m|;�J{��;��o��~7���I�����+���;%(_4E���f[���v-��g����b�k7Ĝ���v��"gCiǆ�yQɽJ�,��K��{��ZQ�U��Kbf2�B��}kH��^�n���b��Ԁ΄ۛd��3@r!��rT�gQ;:����qm����,=&J�XH'yT�;?�d�:�^wX���f#ʜ�Ȋef��ko/H��d�|q
��^�}e�C��0��>��ɐ�m�v��]%�B�Rh5
eEV�t��Xi����f`��e�E}#�;���
�J�P��*��p�r����ٯV��o�\~b'��>6կ�!gtT�g�S��/�iH�S\�Z�
��q��4�5M����oт�wt�~3J�^sTb��R�A�e�1���;9X��{��S���_�Lr��ǄKe�GI-kN�5��B�mw�J��|E�N�=ySq���L� Ge���+���G�_P4����@�Ė� Z�Da�x��o7%씹��pR%��}�b̖�%��+E�Ms,�=�I�H����d��Ѐ��E�D�\��N�ؔ`G�p"��a�O�J��E� ޹V��LJ�[Q��˴��<�SUv��1-a��Gǁ[�x`�,��h$���x8�,)6M/�������B�ȵxْK���Em҈S@q~d�B\�|�>���c�g^64%%TA~���p備��H|.l���o���A�T���túڥ����"�^L�X���@*�W�9�ڻL��
�Y��cq�š�4���XDG�ߴ��r6�g����7��s�;�I �h`cMA�,r#�l�t ��-��뺎����_L��U��]����de��3�.�V��ē����(�F��5*<8@ⷅ���,y��ą�����9��2.cx�j8v���?�a��/j]V,6n�I�Ed���qw�(����Xܔ��j���}�:- ��I�>��� �][%ly󇯬��$�b0a��*J���K���vβ>-�oz\v��M���g��jG�
X
�	�9H5*���`�
������|�v�4��O)ǡX��%Qz�%,��O�?��6���(���Qj�^�(-�K�]�����-����7)��ZGE.�k�i�A�v�4���xT૞�7�(�U���;�� ���6����'��%��w�3<�W�g����B�O����^�����VfwP������+X5Q�-.�_+�w�翜�M�+𗁞�!�fG}ȽHr�^��\Zm;b�=�u���^$�܊�D��<�ԧ �Tv�o`�E ��qK�i�1�&3��l!Z�������S�k����=�QȤ�E���<�b�����Q�}�����Z�"�N�ꀦ߃�㕲���E��8Ec����T�����ZQ$�C`�.���2�l�ą���2��P��|�r�ةѕ�1�����#:gN͜~�v�k�W����b�\A{�c$���D!�UT\Q��^�tG,<l�J���Qv�t(+� ̜�2 � ���&�6QH��ߚ�ص���1�������.��j�����y����T��X���&O��}c�[�9��c���t`'_�dr����W(�C(��6�)JZ�O�m��=�&4x[g�J�,��~զt�^/����U�����á���<`0ᵹ⃨�E ӧD��Web���Oh�e��d�f8%�Cū�p�؈ނ�\�DX�*oZ�8f���@��G,,�K�Jr� �,���)�S@������#�{��y1}�Me���R,Âh����'j��RL�P*��O�W����GL��)��c�n�i��p�鰃�[`��CF1�ض�u0�V���]��M
�%{�|�2�Ͻ94��_z
�we8�$�Bۋ�$�OH�qˈP�<:�
�#������Ƶ1����6�M��~E_a��:ZagA�]���W�#�ԅ���=\�`�%W�;#HI�g��|���`(J�� MUsl
q����O@l��;��H�Lу�"�T<�!2�OI���
��2�|CgR�.KyۿyRʣ�}�{�G|V��}�jGd�/�z�)�$<3�_��
"(2/��kf��d���NQ�U6��H����-y_an���5�����'��������:%��7(�	"IIM�o�lg��ci=f��J��n�=)Y
ct=4��G���w0�Q����ۖ0�*�3f��Z_�Q��F���ՠ��#Pd�ӱ2�?�t�&���؃[8'�� 3����p]ͭ�u���4n��9�L�8@��k�����i�7�����1��<Ҽζw�9C1�J�}�ڧ���N�xpP\?Px��H�z�
��ide�4�y2���D'��j,~�����+�y7�3@��Ja߈$��R4��U�R���b31�����c��L��$+��G����|��	<��z��1�0�k$�N�t{��p)��r\@���d~&*���N�`C�uy歡i����,"%�ow�|c�(��J�?ۂ�Gh�i?��H:�K���XX��g�B9˳�V������#���#��,�0Y��{C����\$�D��=����WQ@joC����Wzub3�p7!��wJh�C�\�S���	�U6��J �X�	b8�d
nE�;Y�|�-:��4�� E�'v[�kE��4�J�h���[��V� �e���c�-�� C�l�	|e���Q������1�RY<L/ʏ暇�J�A�}z ��j
}����|�n쎖��C��Q��¥�>|�@7�&���AO8���!՞���&j���m��r3ʅ|`+f�|K�R\����T�p�_I��5��A�猀�����'��G� �WK��46gZ� <�-�f�X0@���5m@m�n��I��X�&2g��pQ�Q	�v7�n>rV�8v84 ��$�>��H`�`��;�bo}�@oD(�� 0 #S���#3�֠��:� ��ӺCnZ� /�&* Xr$��0^Wd��k:��z1jÆ(k1i�"��ճvw?�qL����$��dSL+wԧ��޹1jt"z'�p�q���_�icA��I1���BfE�|��Nxy+N��z��w	Sb)�)�^��j�dCIAݬFx�hn�6�vw`׈wo��*��F��$L���r�N�>d~���O݅}x)HF�վܿ�v=+=�RV�K�Q݁�ڋ��X�w�<ks}�̵���a;%��9�¡*x��l�'�d�'���>���`j�-c���P�
�LP�����c2j�X(�b�����\�5����`�֯���1C�\�卍#S>~Қ�ϩ=? ����#���tn��OA�9N\=;�j`�J�_����+�0�	��ꪙ;|�祄J�QP'���L�x�A�%Q�q	�9�	C����\�md�|�W��4�N��[x�	"�Ы���e/z`��)鰝�����x�-�a��+%�zԱИ����Ba��nM#����<�cDC�N�.��bg{>;�nTļ�x�a��Ƴ&�K��B�y�Y)��O�۲�ᆡ~���6��)�1���v��]�A���[�l�*��R����R�r����j�k�Nw.֧�?�as#��ҩ�u$���u
%K�(���5�����6���u{xK
���J��t�S��^��w�w+�.=�A�a�E�(�"�]�H��z��k�����g� �J�R��BU[Xܩ c��E�����ы���tS
�  ����-�´բ�HU�x�꼖l	�g{�3�3@��y!��|V�sÿ���g2��ӧLy$�9������d��;�|ι�p���و���~]^Y�ɡO�7�� u���?6��*��1W����`*��n)�AD�<@#�E�mLp�cy5�qh�K���N�$I� �ɒ7W�s�cV$3��5<�m1�!����+���[�F��P1�6�����lz`�i�&��آD|��Z�4��ǭQ��XaӔӘ�!3:J�( ����<�ܥ�y?w�q���IR�I}t$�!^`%s�ɨ&7H^]mҋ��(�%=�����q�&�h�|���xB���������J'��ԝ3}'E��Oŵ&��S;�OKƴ�o���>��rcc�08�r�`��G��zɂ0\~���׆���n�(]�G�ra_F����7 Ys�k��@�����:Ѭ0�g���%OU?Fe�ħ�Q_ʰ^#����ЧDi���12�:xL��(�ad3�^�=�.�a�u1˰+����^�NA/�e�i>���Z�Uc3� ]{��"�Q��$�)^��%��K �D�L�4e3]y,ڈ�K�ź6Z�:�.h�S�VM^���8L��cN�l�J� �k����`����-v���sC����xp�M,EM��8�H4�L,~�}�~�)ξ��� ��Mb��`��=��)���0=g9���=�
�]YL�q�D�B�a�񝟄7�6�>G��~�+ĝ,�DP�]��a�ķȽ1-Q�/m�����՛VV�/L�=z]����Q��WJ�;[�W��Z����ܬ��㈥�Q���XE �.ŉ��;��o,;�w"�	�R��3�3�p��(:�{"Pj.� ��#[}3vN���7�a�p�>�	�@U�y�����H������ܟ�^C�<K��K����@ÂHqf!��0/�3h�i�0�9k����z���?�m\Q���q�u�+���,���:��X����c�c�SV3s�4�si`!�oF�B;��/�wF����Ņ��6���t�\�I����>�B���xA�0�C�J^:�/�Y�mg�q�d*a�|U�m�}HY-��� mU?��.�7a����I�����d#�x����%�Z�!���"�+>V�?���>ܞ*�_�=~� "�� ���g.�%��	�[����?�y�8=�~<��+�	��T�Ѷ�-��)��8��cA4�7Z�F� �{L�� b����d�aQ�a�Tj�c7;�j�<=�����|���$�ڥ�����)B�d�U�� E��*�,E��k�o�>�@@�}~��N��ܓ�!��<�WuA$#�;�1�QԾ'���l��R �Rrh�Vͣ����`��ԫ/���|9vb����r��M� �_D�{6:�BVb�T��������*�m�v�J�?�si�[q=gy�Ҍ.��\z�Ns	�ZS�g�$,yZ4byBz��x~�$�s	��G�K�"ZC�X< �)�����G$'F�D���|c`:���]܅Vĭo��;�c��P���n�!����l�BF��PW��Z��� �I&~��X�=6��SV�i��l��5��'զhL<��^�Yy�oG�����쏈	��[�'\�2�P!��E�SY��3s�5�f߬�QR�(�vr��C�B����TH���Έ�hpmϷK]����*��$���x��0���8s/Z��
�����	F$���䠶
L䵯������ �#�~��d|ԙ�luTpzG0�lWW�b�x�0_�Edi�Ͻ%�MK��p���4�AN�% �?<S3��騳;P@�Ő��d���Qk�}�-��h�8[��Z������N�Z%U�0�J(U�XhD�?M�����+O�Fjt�M��{����u	�8R�:7�s��j�B��`�]�l:«�E��b+��"sT��mCaf��P�ڴ���m���ڪ�&�pi�[���U$c/��5�wi�_F�WB�T��?�2�-�,��¬�I�F%v#�f�V+�ȣ���@3�I���hJ�V��K³������r�=L�OJ)dZz��>�5Gb ���Jk�~t�,��J3��7i�u�8�ćwYK��΄ۅS�<��"kj;ye���M�-
��F+�4D���uY&�:vk��O�ʷ=���ڱ���c�����Y���0��h��b!���N��z�.}�k��~u��E��y[���
��� J7���M��_yյ�u=�N���N��g}���E��xB�AY4_��tGP�2b�#@����r�ОK@Uǥz��ߡm<�]$�����^��3����	�p�?ڹW�a�����hy�n�x��fI3S���X"�A�����C|?3QC{�
��y�W�D��r��̾~"�����nz`�H�V���E�(VJ�jP
�{��&YG�����������g�5��4�-3sJ�XFu(���:>�ns��p+�����.%#}t_5���H���۶��r�q:�Я�\;b'S�0��T�y��$�=�6��
����9I�Q���*��UZ��V���5U-�:7R�TKI�G�#i��U����Y�ܞ<ư�I8պ5j$¼�R4�c�T(����th�9�B7��Bn�U�C��<(�^����/k�s�Tl�87<
5�h"�j�͙��Hy�R�,���UVQ�MJ��b�#�����t)4:FNdK
�ʂho���=�E4=X�2��7�L��4+b��*&N�̉��~�d`vU�O^-j���k��A��J,X���r
�؝G^����~�}�M|�|�y��1+�{�:{�������>�P���4���	�U�-��R�I�X�o��TXV}��� oO��=�1Lyk��3n��v���п�*��a�[:����u ,pa�=��i�9��p��ި�q���	�K�@���[�+b���I�R�CQ��޵ѥ��PpزBP� 7�Ѳ[v%Q��5|�@��� v6��O��lm�ɲ������iCfT���w.���O��H�y��Ӣ+}U��Jh
�N�
Ǚ���n��Q�##>�<�^�����	��5-K��5:���C!���^޾e2��qQ^HK�dC7�b k^K��R����g6��1�a��%��u.�DP�4~	TD|�
I�X�W����ߢhp���&��w���rD4����;� 0ȩ!S���g`�1��{b�0��YJ�/�����>�8�^��V���e�#^���H�
[14���˴�hiu��uC�!��0�F�	��w�dS��HhOE�Kl^���D^$����C浐S���d�@��H?�/g6���|kD`�7
c��)S�b�?���&ةD���nϬ����ޘa�H���urp�d���������q$F��K�G�;����1��>f�<a��j+7k���i��]N�O��B�/�l_�F�V0�����[��`����b����J��Rh[��!�߇�Y�NI�_E����$�8�b�݇��m2Ζ=D!�]�o~���8z\�,9y9�䈲%Á�i���>H;���?�WmMrΏ��dkN�D7T�+@�d�z���o\~{��,��r��PH��l��<Š�<ӥ��dxu�-j�G���Ň����y'�?�����vikq�=!0����tzu��ї�hC����I	�M=���H�߬#���.���X��i�*��|��-6�����<9��h&%�o!K����+�V�-A�Rn0˄I�-�a��:Q�m�[�በ�	sDp1��������������<s9 ;�N, �UiM�;�7BPM�����0c�#\PJS(BH�f t�"D^���Oi��u�8$�����B�e����L���k����L3z�ɨ�c��a�N* (�$�@8���ů�3�/tx�ǎ�Jd	���b�ZO�HH��L���@e3t�[~c�~��º ��Z�y���}��k�t����F�^� �'m�mնW�b�3a"ܩc���<���p��u�����^�,����uq��l��zPO�i�o�!��{�4�-���`�OZZO��v�6�r-.��8�Hw���<��LhҿL���<�Hu_��F��s\\(�����ȂR�����!�Tp�1g\f�d.�>�dy���#���mד�	�.Tt L9X%J���C���Ѥ�<�J��loR/m� �N�݃�q�A?�L?�,�5���	��e��_�Q<9h��.�WW�{���o��[��I,��D�9��Ė�5���h�`�]��f~htK�/&~�>� ࢙���`E�Τ�J']O7���m��PlO�٬ڹ�)q��=͛�H1�4�s�Y�Z�%�7�>m�r�%������LD�A��-�y�)��_�6ia�W3�V�ښ�����ˤy���|�l���Y��.�fN�V�������A/��(�yƶ�	~8�C����7u[;�Ckohu�`���ʇ��!��(ͱm<�Ԫ1���[h�1��8�SB�R�-+��C�x`�cU�Zg��r������� o��x�(�@<7�sWȮ���5�C���m*�GQ�
�f-����H�	й��14�%i��#4l��f������&2�]�cD4�9��/'��pb�P��ｷu;pI�bfy�=a 7�eM�tb�^����l�D͖���-w����2���`�* �G6�\�j�����B>~�HT�,jtc�BLx�^����q�5��x��-'��9����V���\ԁU��k�Y���Ydh�)�s�*���o%�m1��!�<�x�.�;fr:��x��5�pꏪ�Xx,�MY�2M}� ����#�ׅ$�_l
�Z�MW�&�]����m� K&�!��s;�s�I�L����<���ݑ#�ieGV����i�m���8��9��Z�ƀ؄f�%���Y7f��{�g��l�~�J�`�њي���UD�#�˱�����2�b�ϼ�7YTZ_O�p��G[��RK�%��u���A ����Ѐ
�`|�B�R'�]��s��
ZSUsi/$�rg@�U��%��Lg��qV|\�$�Ȍ�����F@��9����M�TEC���A�P[B��)�D��O���s��P~�i�?k慭��^����ezZ֐�#5�rq*��L�&)w تq�����0� ��G&�S?�3��6%v��*����������c�ub�88�F�U%=6�\�i�#x�-�T˱�!z$����y���ͥ��
|��گ@.ۛ�풔_��8jL��OS�6���S��R����d��Q9�K�fH�`TQ����dM�5��e/�%��a�[z�����k��W��ϟ���Ĉ�lJ`�ٿ Ej�j�sYǧ�L6���1��\#�L4����c��n���■����0қ��ì�s�l��ҿ$D�+���c/8�QV�q���Ο������s�����8|M�Y����j���O�'���8�G!P^�;lٜ"�K2��]�>-o/ܖ�=m�l��3�����g  O}�H��}�6�4��\h&]XD�b�eЮ��[�q�\O��f��C�Dgו�f����eu�zP�_�|K����j���`�	:�;�X^�ki�N�ޑq7<w�o$;��ה�62�J�$ʝ��aɽF��ϲ��#�����n�'{�ƩHQ������"�f�����ܖp�+��Y���1�����+��􇑘z�\�T�Q./!�g4��3�R��p̗�޷>1=b��b���Y����'�OS��)L�3�rzG<6R[�k���MT)(�o)�Zn[.>hX�6�-�xK��H2e�h&��8G�]�!چ���7�T P2L�M��gK��n0ρ��E�u^v���|M������nu��E�9?��t3۪tl4��'p6D��˲�cjۊ�D�������AJ���W�G��lud������%����.��e[B��3�s/v>6.)4ci��ƈ���1\�~v8���Tќuv̡�;R�h��v��)w" ���S�����5B~�;���RcC5؅�e�HJ��Pl��O���:��=�0�w3]���o݄g���I����0�T�#�)�4a/G��Tj������-������d5�k�|����̨˲�Nj2k)���.�FVe�Y�*��ꗑ�U�����>�.�S4yc�D����`�@�Xi�S�L)�My�.;�&#�2""}�co^�ё���2�����xg�w���|~H�,J�ś:�ߠ���(�g�;��`a<��lD�o�M����`����u�RM��ۑ�kf���kz�h$���$V��TkXje���+�/?�c+O��	��Ť��i�0�؆��Z$f��Ql���Q�b�p�$'�9���㨪u�9>g�>�:,��ع!��Gq1�C8x@�yM/l�,x=O��O�~}i����@�w[Th�iU�~��0�$휎��8Ao�1�=F�dS�Z.�}P�'���Ա6��n�f���cHP�s`D*��p`X��')'�y˅[d����N�xs�ʞ.�5,��
���s��nP��~��(�tv�I����k�2���F%���9hlV��wjϭc7��Wh/#��b��ME���O��0JVm��_��0�6���ZZu��`���`���e�r5b�̌yE�Y��P�RܟG�t��'4�R#��H��w���BznҼo)9\$|C�t3K�5�m�;a��S|��D���a�8���g��2%�/t��G��a��`��)o�e��T���[���S&�ևrx���'�x�5e~��v��D��p��G�֒r=Sr�����V4{�GI-�&t�K���&�㙤��O��h��0�6}��p���+�2WN�.�����>�f���ϯ���Ա8����!�wf�R���eE�����_��REt�)+��*=n
j�Sv�Od/a�~K�� W�9&�v��J�����cm��&m���%옧b�t4U�����:�e������fu��ͨ�+�z�D�hUؚZ��i���"�&򱪍���x�L�`��j,���ӗ�l�:V�6�e�K��8�\�ة_���p��MJ�{�%u4��O��US���P���%⓶�����!�2\ FϜ1�ͦ��s��{Bb}W����$���r��H�-:`=5Tu�1����]2m�	*�ogBjKs+9ws�ƦVc��I~�[��"���oT�l�
�ím��J��	�.�5~�ޓ�*�f�3�a���볐�'������@��`��/c((3YW�Th�b��	li ��6Q�)'5�i@�\�j{i?�gj��6��i.���㉵ �\��j�v%)���gr��X����52X^���}�:��(�ݐT���	)��4nh�!�h�5�]je�x�B�Áh |;�(0��{>�y7&�MDX���]̻�)]�hQ���p�J�
u��1�eD�e3�`dJj�(�)��uN��G +�l��c1�y���Z)��wlay�N�Oe����%o����0��)n�3�7ǽ7<��#yW?sn"��\Z�ݚ��h��ǆ1k��1+��iwM��O�+8��{��Q�5������*^���7��n��M?����.;��'WЗ�3۷�����庌�$ߌ{	�G�yM��٤��.8f\��A|��gV=ގ-)v��i	���s��s?��giB� ӂ��H���ڡ�|&W��l��W���� B���jmu5��w�&�Y/
߼q����%���0x}gh��u@ �t\,�:��	�J����Yƣ��A�e]��q��k�x�!7`@˝��=yP��0�!: ��U�K��r�/2�ܥ��8�Sf��Ux���� �l�mp�ꘉ@��-ωt�ơ�.���.*_Q�\A���c�*�8u��ym��mg
4B���n�l�{�G�$��O]1�6Q챆�{j�M�AQ�Z�R�27fbK�3�put������!A:�U���˄,�;3U�d�L3tA~��ko���$ޢG�5E��ڝ�zYy��(�p���]�7�@�n!�sX�@ǔ��<)�1��Ś�%S�`�fe�^�/�}gR��s���K�*�K�m;VE��aL���v�f�{O"{ڟE�W(��Q�.��c()�j���i��}&q� �WBf�X���L	�$RJ?���bX�(�`a>*Դ����Jԣ�\�s17��1�r�`���0�� ژ��62#+�x�"%l��8B���
wC{Ɩ��$��?�?��ٕ�����k��G�G� ׫�Rq�yc�s�F�����$��fD��/ّ>3D*����?�Ej��x�O�<�Vc))N.]�^�؃(q���޽Щ��|�,uΣ�[���w�"
q�ۼR�`�K{}������0N{�f��� đ�yp

r���D�Oj�3I��.�(�������j^�$%���y��q���}��&�1Z'���0���NVN_,>]-�e#����a���R�G.N*�:Ք�g]��Aq{M4Зw�����n��<��Nč�x����R�S<��h�X-�<#��$r���ʹɃ� һ�����a<�m+v�%��?�
L���J������XW9ApX����Ԫ:�����5�X�C-��I�:�`7�N���tCTld�V�|�Q+��P~,J�[���C��k�������j����,��{d/t}���4�*ɂ����7�-�𻒢uMcf��F��7)8w��*H3�9��
�m( ��; ��(�� ��ò��'ڊ�Z�(˭�?1��>�:F�	�	��
X�Z��DW��z�T�\�X�K"Ϡ�{��ΰ���d{�k?�D��h��ޅ��I$ ��b+$NgX�Tbn�*���bǛ��g�}�0�WO.��YV<(p��.>w��^\y+�5������P�CT2�/R�/�^\�m^�L�v����k,��}�]���Lz߲}zf�7�R��0p��Wrh<�;5M��n�eb��=�rQ�3�%�+[{���}pz�_� .'
] �5��B6��G�3�Ҭ& ���(��d)�Rv��.��t�+�^Y3�̛zB۱TտN��λ\mk7A�5���}�h�����F��X%�He
�]X��y�CQ㝋�ʐB������l�����I�䙶#D�;����#
���
�#j ��
5�\����/~��)�l�+I4�������y� ]/
��C���g�? B)�:��B���%�d�E|5�Ơ��*��(l�Y�R
�F��)a;^wL�x�˼L�<�r�
o.�͑8���} K�O��F�����9\��w>`��� ��@��m$h�r��jd��#�X���"��nܼQ< $L�?ܒ�����B��� �8���[!�`��F�M�v�#jǬ6��Է�uS�,9�H��,��:A�X����ЫuM�Q�F��g���[:��9Q�5�s�dp�mm9�~�D۹�������U����!�d�ŋ���ؿf�O:�zۭ��M�ҚTh���� ��O����eE�w�T�Ac��������AJy�c�'���RG#Ql���f��ȕ�8U�|��k���!��L������ƽ�.������.�T7fM��s�-�2��kC�j}�:f7�3��J�	�Y
d��S� �F�?a泆:)".ثʕv��/+i�N�������:OO$ۯn�Jlv��_�t4�ii��犸Օ$�֞ G�'z�}l�W$�Gӑ|��;�7����^^�}k��q��k4۷�K�6\)_��d?�Iod6V��g�g�,j�Y�$/�qe\��q���3�V��%��i� ��j���7�$��1|��!�:��DO
���?Ym_d����O/S��;��� P5���}W�'�$,�)rZ6j�t�����C�� kuX�9k�%E��$P]����
�6ZF�"��w�r�);j7i�������4���"�d�U�3pl�UW��K�Bt(dH'7��Sdk�+�k�ڥ����e�4j.�n�����En2�	A1�7���������'���0��Y��{�� +��UT��e�$$<�^����W�N�ا�`_�k��
f��C�{i��K�n���R�`��څ-`�}_}���=�L
vp�i�za���Dk���!TD��J8�n(3�H�8��,�֘�u�d�i⺒���#�b8>��DaWr��>��Ν��&_�]��ط3��w�F�ϒ�3������7�8��[��ǧ�`9��J}�������i)����Mv-�<�T�k�3r>�݇'�H��A4��16��B*��7v��BmҖ�`Io����2'�_{�m�5�7y�p|❫��.�I��J#����k<�[3/O	$����=8�{<(;���G�������vn� .�/��*O[^bݻ���t�2D���hF��r�2G��낗���8F�n�mu
��ٿ����`ô5;��D"p8-����g(&J��P�N�ƊN�����
?�SH��.�ϝ�l_��\����������Sw'��y�W�"��	�|J�YU0lJ����ǉ�G��yپN��B�[��9:DX-�r��q3�F�n�'�= � x�D�}~a�嚂�oy�	�G�c�>����fY����ø,�F��OD�r��Y.-F5�D��+_f*��pb�'�`!+�`7�X�
*<e�mg{�Zc���3X�� +�ۻ��%�@��H�b���W�΂E�Auǰ��XD3�I��z�Y!�3��ǵmZn�]�L �.����53��(;��Śk8�K&��Nzb���ZQ��a�ç�Κ��Q�]�Y�;�7C�����%��g�X�?�M�f��Z�f�/�S� lG�y܉s?:��j�ލ�o���;h�	#�v�K�z�cU��/�K�.�/�s�u�8M���]Qj�P+Hd�7�Y���U��`cY����XwL����N�҄�fIH�؞M�������Ǖ�[��h�_�X�$��uLB��o?��mh����ؗ�(����Lς'紓)D�X�#�ñP3�d0�}N��^��Ǜ�0�OG���w0t���o4����=��z�îS+9,=Y��'���
����Z���d��SkJ��K����%�w}���[���
qau�y[a蚷=�p�gj�鞦�k��&.��D��MUA�&�!R�	�Tw��%^ɔ�ႈ�V-���m��W4���g���AD�R�][6�dZ��C)=}���ނ�H���NZOwA~����b䊟UBl�f"����c�J1ڴ���SO�Y�c�@M��):��y`�}E6��|�Z���P<��W$���+�@jtJ�ΐ�� k'��{4�n���P���O.*�S�zeL��L�6范d/�U־�f(�>����ٶ�^p�����Uz� �}�0"c|wB%����&���s����}�y��I�}������ߊ�~��Z�H�f= �B���Q�Y���O�z�;*�Br-�D�{D8�
���.T��rꦌNe;�4��K:mF�P�W<�2)d�c�yY���$Q,����N��'��Ǵk�GQ��9��8�X�_yon�.�$!02���O�璔����������I8�������Tt��J��j���l�ݣ���a���{|���n�[�Ɇ��rv=� ?{,q��p��E���M�ߝ-����V9���NF65�6�7�?j�$O��h�����ZsrzP	�ء�5T1R|�Җ�7��`ߡ���*F=$B�牚6�q2Z�RE���v��'��y�slbQ_`���A%L�c	���|��@�[��G�hJ+l�!
�RL�Bnb̊{�q�D�v�R�28�9�h��ᖺ���.x�q�M�)M�:<���~6fzt�x�;�~�s�3ٱ�~<�I��J}�z~s�g+�(դ�������;�tUd7G7��!by�T�p���0��<���'��4���?Fy�/�}m0+e*�n4i�(}�*O3�Dp��~�#�|t� ��*_�>� d����
5�D�i��j��@J���.p��#mԗ44Ҩ���4�lJ+�g����&��$�kw[mMS_�߉N�:��]�^O���rܐ�pli��M�����<Y?�yiMz��e�M�Y-!,H�`?4��k�P�ʶ����{��;��<iaT}����]���zM�g�"�S���}5$d{kk���K��
��'{��4)0�Yi���;]i?�Yg�3�`�Gĉ�ٴ�*�n���H �=!?b�g��b�l�\F��t�Gv�_XH�S���A*D6���4{���k>@�3
��.�Z�QVI���c�������y ���#�m���r��:�H�i���(���/EK�`�m���a��d�w�X_X�ɻ����W��4���j��v��"�����<�#�@'"�,���R�; O!�3�釭�f~�{�&`�64�$�^$��� ��y�X�-�OK6���8 ����h�z �HX5cL�l�bY�Po��R��_p��RˀH�����2���@�F�|�l^)~q���	�)�\M��!��h����?�/����>�&�qo4��On�$6��p~XD�$�A�)CD-� )�1P��\�K*Y3@TW?�hS*�"c��O^�5����jzZ'�՜�$Bu8L�k��a�U0%��$VUȜV�0 s�po ɩ;���R.\�s�f����Un��Ƒ���±��S3hW�ٻ���y���P�_�d��~T���eA���𠱿?1�_�:��&>�������X���� 2=�� "{+/ Y��B�+��Ų$�Y�B�dH����b;�*�Eڍ���������mG)2-AE�B�2��S=k�	�س|Di1�C���&¨�t�j{�ρ�7� ��F�zN��{<c��E8B�,*m�]92�>�a�q�1oO.�a���]�Q��+=P+80[0C�c�|�T�:K��}�i;;�45}�SNb��P�X�_p�[�8rR:�]���&1�(�c��DLl�;TZ����'��7�_��0}����_U��-�+�?���0Av4�49�h��Z'��2�>��(8��<u��.���$j���߆i���X��rZ!3d�h�vѦV���&��3v�[����Q�H��@IT<��K{�^J���7݃з�s��Í
E@ WD�A14Q��֫9�<�q��:8���s�a��C%ra�z�8�禡�ع]���2g ��:r�����*�c,F�ۑ^s+�m,gS0�B��<��'�T���'6a�(�e�'/T��r�P�	So,��#����P��������N��Db��`K��x!��{����n�$�_:TK��8�d��e���Ӟ����t��L3�$]O�����jM������6ۗ��ď]Q�7����E�P#-��ے>�!��zl��^�"/qų'Ӽ�\z[��V��ǡ�RU@�Q�?0Y_u���	p�w��RI�U�0�<��¢�
*"G\���Py̛�&�uI�
=g��l^�^�q�F�(L�Hښ���'5%��Ӂ�,��FRm��x��4=����_r�[��b���l�2�ՔwB�Xިu�L��i�c m�c&���6C�"I��-A� �}��`Ž���I�9?|6X�b�5�Fϭu�x�!�5;��}�j��x��bC[�཈�~/t��F���kY)��F���,�y��T��)Q+��SpP��p�
�%:��N�Y�Ҫ>�Su)	�!Dy4�����|�L1_K�C��?lEj,╇�y��r��� ,^N<���~[��s����W(�j�3��Ԡ2�J�J���������9y�Y��f6kֽ�x�G�� �Q̬���U�؂e�&�2��	#�s/��u�~�
��y~���6��헎��-(���|hY����s��uH�dx +�9�p�������gI���z��4D� ���^bK��c�.!�?�V�-+~�s�O��΢̤��4(�໥��)��f�b*#�R��:�J;;��%���Ewb�2i�[��>,>��4-5��nX}Y�P���}���V��S�f���bC��5"�$����0X��Cf�ͧ�N�R:׹9[����J��@%I�߳�{4O=�t>anC�Y��zi1�%��a�'��u@�F�B]�������y:�YEQ�&,Q�T6 ����[
�@�)���uG[-	�7t%�A�u�'٭6q��tiN�yH�I��֧�u6����Y���̺�3Kr�@�d��Ew�q�*a)�Q�pz�(�C4s���$�ފ��+ٽi��Q�������l2�DE���b�S>V*~�G{����_=� �<q�9�,�"�g�׌oz递N��Eɨ��8����ϳ�j�N�
�nEFէ^j���Wd4`��Ѭ���8��2={EѓB���ˋ#���򪲵1EǞ���4�l|��d�iv%0�i��ǝpd��X�"��!EX��Z���hT�	SGN?�~�V��l̙����Qp T?͘:|]`^�����h�?QM���t/!,�`���Z��s�CØސ
��$Vv�J �R��ЏbE�����G8��tu��Aw9&�H��\
���-��A��M�@��,�'��z��p�X	�����^�����I�1{S@�C��牼N�|4�Q+o�c3���2�d��7\�P6�)E����f0]k|oTEC���2�m	r�OT ���$��\�Q�DTB ̵��A`��ѻ>B.c��eXwi.�="�!D)4:���*��eӗAFC�py`]xs])��1���@9=��9�Go�Q�3�jz��ws���?5R����AƜU9�d�n&a�ᏛI�]V��z��P��s�+���A�}P���֓�zm�O]��mꋍD��zr���_�L�a�qr5��Q�f��cR�D��jH&���d��u'&0빿��o��[� ��܇i��2���5��:G�'w��ؤ����>kB�E���"�jԵq*�����-�8��B0l���^�L��ս�w��]�M��7�S�H6U�zK��O@[�� &>!�S�iQ�F1 ���?���=��M'�5G�ѷx�+Ƹ@�+�G�#�M ��_��v�(;����x_�l,Hݐ�AJ�j^>��I���Gu�<��ѥ�mI�\���#u��$�ߛJ)�S1q����	e:�z�����6��O��a�� #��WߪQi������G��=8�n_g%�:�:���� J9
��`5�炝�wم�}�]�u���8K����EY�
��^�V�:F�$��x�l*�I@�M�(儴D�3��g�m.f5�
O&�������Rρ2��Vwl��HJ}��)�Z]��Ö�*7QL���{;���q12Ϫ-�V)�1�h7z3����AN� ���,�v�&��������L�K+b�V��,^�o�e$c�>A�Ud��f�f$����J���FD놽�ƙ@:�
ō��ݱJ5���TD���q�ɞ	��3�����׵x���o����;6�A��!I�\�9؞�;|'�R<�f	��˅y�L��$RASR��;�#~�	���GR�}4�D�G�}
8��#EF5�����m�BMϐ�B,ab/��ؚ�yx5'M�@�9�32�'?~��Q��#Ǐ�:�t��k��e�g����>�1���{�Dpį��XV,�K�,aj�nYp��bq�^�xh�0���k�K�q"�
�Ԫ���w:�]�2�)ǉ���)f�\� H���<9Æ��!�"\��q�I�l,��Ν�Ч�5BW�_{������5��|{�;+,�쁎A�Z��A}|��� �Cē����ս�p"t�<����H��o���k�`�r���B����'D�$�����v�oꝊ�|H�7� �u:����i��Ie���b�OS��P��]~J�v�w���0�H!ɋ�Q0�S�`VTѨ����Ħ�E����F�q���x�3B�:.O5�x�����Rl��ԟ-9u	���Gf(���0#��O����4����m�pz���$��s�6�L"K��gj����*{%�ؤgj��k���7��]a�a��)��RU-;�H*{�_�/�k&)ԩQ��>$Hx~F&�H��[C�=?���4�-�H�ZF�剈B��Ϟ�'�'�Y���5���jPպ�?FL4#�_a��X�֓$���.�ƊY��N@�\p>��vD&��Yl��V��2Y�d
o
*��2 !ip��	��j�PԻ���;��H��� ����޳r�հ��tbz��a���	��lI��e�~X�_`�U�pG��T��e�\���~�!�@9gr�w��?��o��Vp�����.�u<Q��9����{Y� ��~�YNs���h�vQ��0+�}N����xt_]��N�Gt�W�D�|��O��cV�s�����"lŎ?��:��-��2��o`2��pֆX�������R=�C2���	,���T��V?xc3��\{9n�Ʋ�j��U6�tg��DT���@&H�N�~��uu��3	<�S8Ջ��}Wƹ���!_����y̻��շ���s��Y�����P6f�
���18B��Ri+�n:���pd�_��_�5�y��lM9(ml�k�'�@�cl��V\=G�z:<�ʤzC�V�2�����D.״��ɴ�i�Fvk�s5�;�����eɸ"j�$��{����X��1�?
[� �IX��铵h�Tyb�	Ts��{�ٟ�;p%z�4�2������k�W�11���O��)N
ID��5�2P^aqh獵�l�G�ݧrA�UԸߟ�>��o���G~&���վ�[�,�kPv���b�jivj�.��,Z��{;C�������?UQ<Jo�p'�)��a���XX��p?魈9Y���D�4S`!Ph6���T����<I��������ۡ�eb��[};Q"ݰ%)&�	�x9�&블IH��&��~q�����oz�dc����Z�?����YeU��h6�?��A0�=F
����*տLT��ů@@����6Y��1���u���}�ӝB��%c_���9~��B�m�<u�DƤ	״v�rRٝ�W�*ƐAR�ǁ���cr3O@��1�1�XfO@ ���W�|�Qɬ�e�9����i��FG����ȼ-��(��]����5&+��2�q����N'�-���<; �.���X��������V��؀�769�(/@������:,�v7N<�zŅ�
��P�:�����Z��GNq �YL2x����2����y�����"jO��y�$Im&��.�]l�^<�[J�����UMA�|���:V/��!_&0(S�$���d�v��D�����I�����b7���z ��Gzz
H|�tU�Ö���cO�,�.�)�ݳ���b�Ἐ����KJ~�v��7�M=>�X�W{'��\� �|).N�,�46xFX8_|^�#N��ܒV�h/$��B&����Yk� t��i/\�����gzł�t蕎WyMYN��Rk�7^�q� �M��>|�6=.�agv"���76Ɇ�x�r�v+|�fR�
 ��#q!{t��f�X�O��2&����td-kP�G?\�̥�1�;�i���8�	Tk^�u�?��R,�.��D����-�l#Q5 鿨H�������;��O�~�0� ���Y�6F��Th�`�'��ok�U�dY�.Hc�7��7��e �8ߜx#�@��
xA{�
�%�����]*y�_VM��lE���� ��4��֩Sp�4��a�3�[�Hal>�6l�v`�&]�����*!�ߥ7�k�tVf��o�>t�_iic��L	����5<;{6xI�霽'mH�VFaC񤴟�3�����3����]+�dF�2�(�t~��a0�G����ě��g���N��7��ʋ�Ń#��y.z�H�H{HE�����l���r(R�~�/~���E����:�P�	J,�Gi���t`ph�`P���\ٟs��X�5�)`yZ�ë�" ����,?<��� 6���y��+{lq��_c����=fޱ�Pm�k�@�i�8d�w�6��w�N�^O%:HfB%۶gBSt=�6��]�Ap{C�9��% ���9Eм|W=�p�f�SbY�oݰ�=�o(^v�ۈ0�A�h���jH�0��V;"���ʣv)�/�X������ZsK��<?B��J4�5 o#�����LQf����:7�b�����pa7�%�#q��]�(�:�Fd1(����b:_?}`/�ZڠR8nʓ���՟��}]��^Ir��|z��v१Vs��`EA�~�Jt�8���%��q�1h��a��W�HD����T)��{�j�&��Xi"��p�_Px�h��
�c6�Q�y��5�
���Q�u�0Q<�䪴~�l�}]���v+!�����ĢnH{/$)W�D���p�T�Q�E���tW���WN��|�����R��u.T"<M
��
x��h�*�ʈZ�^"������/I�2 ��W��MP�rV���2����x��ҟ�T���������b��|uv�',I)�Top���M;���\�^o�p�(L�@[�!V'�`)�:�#ú�X���ҎAp��T�
�LS�*�ҹ�YY0O���P���L�MJ�(�y��e'���ȍ%>f;�V]3�)�=���~}ս����أg38��7���P`�Q���[��z(�<���]	���<����N�&M��K��ŶaxL��w��_��\'^;��X��H"6�e�&vݝ�zms_E#-�9�B��hw���^{�"Y����
{VN�A��ɪ���m8����XBZ�8��'Aw��}x�i�V*��@��krq�t���)�Z���J�s��٣�ZGL�v�[:~4�xdXZ_��b���v��u*���.�6� G;�����3�I�^ڎ�����S���R��aP�z���h�$[nԥ�*D�b���m	g�#&��!��ω5��Y��+�%G4޲��ݷЋ�m�H~:1���*�u� g2^a*p��y�d����`���.�R����>�`���%�ǐש@-u�ǚ1�Vm*<T���}z(1��,��x4K/�����)|�Ăw�5�W�!�S���Oڥ3��D���;��J���C=�eT�[�-7�����Ln�m�� �ͣ�iP��r޲�]��G��dtN��4��ȟF�9��i�%���B�u��4��d�f�pG�o��#Ao8޶}��*	51���,���E����p��&��v��7�c�e�/ �ؓ���5\�a���8��u��,���4*��zd�=u5+���F�8�\����'A���b<�JAM?US%��,�6�P�'}WoKz����{&�tJ֌�Ǔ�io�Sۧٺ�8�W\��6c]�	pv��f�j[�%O���&�ǎ�|/�vg��
�X�(05dF�݌,�`9���d�C��@-m����LTu"�6r�Q-�w�m~ĈMљ��4�������_���8�"�j�,4��p����b�IH��Y����3���ְj�q	6J�\"��F^�p�7p�O�urr1�)Wu@F���Z�nI(<�f|4	!N�t�}�w���Zh�I�zć��
�F^���r�(�K^�ʳp�Yq���[�Q�nY�q5��H\�O��0T��dA�gH.����ap����V<�f���8�'���dǄo�A�@����
�zm�uT�d�'��\k�jcAZ�X��\z�͚���M�	.�"�ȟ���Gd�n�`��?i�V)S^~@=�Er���y�ڍD^-���t;��@���xe��a[�]z3Ӝ�
v u5�^��g	��k��,bq2����M�6@��W�I��6*]�-ol�l_Ba0��Uȟ�s���EȳX´� d�@�~ȱO�cNa�M?le�[��7�TD�_=�)�+�п?�r�c��&vj��B��^�w�n��X���n���5�,�ւ: �`/�T���!'c!h���kjW�=���$7j���}V+U�RXx;z�j�f@Y�%���J?(~!��7'Ю��Z�!{-i�Ď�a�������O���<M�c�ٕpL;��g�I��Fk{�s�U��r�[M���_�//BN�2�:���%;f�I��c���p�۳L�7c"B��j��ɊZ����ۍ6��Q������u���bo�m?���׵�7-���Xcv���w�j����	#�q�Z����d
�H��`�/��9�y�zy-z�Mz"�^Y�O(�Z�9��!�.��'ӡ�2OC(V�+��C_,�fi���k��P�g�t1E�#+6���	oܨ�����(��.#�V_��t���묋��A��r��BЃ�_'�v;�kI~רS����o��)�iFR�^f9x�"Y�f�H�دa�y��h��-LBZ+Ɲl�2��;��*|4�~�'v�)DgAsq�_��HTp��"�[�o���c��t^��Ց���{�'��{�.䧇�LeI����	oQS%�7V#����U��]�<��qЈ��� [ ��(�&�Q	Cn�Jԑ�L#ҏ��aKb�[�������B���å��K�qT;Q;����*�Ĺ���X�2��r��Z5+>��FόYŶS�a���e��'nfڛAŌ&�5�$�l��h�tļ���K�T:4���t�ULA�+��]Rq^;fk��(U�����p�b9�Nvl<Ť)�!�ҵ֍j4D-Mc���6oF
<0�ݲlV�O�(�0/eP�����3!���;_��n��2#�bv"��Ŝ�Nr�zLᅢ�����8.|'[�6M3��q�];3���>����]�0j�\<}IV��Si�-�#�ժ���2�)�5�[L�:F���85�$�l٧2Vtzv� �O� �6{Lw�]�S=q��]o\�xpim����+��!��;��p��g�GIj�Ǻ�w�N'�b�ܞ�������e\Kb�{����{D�4�a�S6��Sk0���G? ���