��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*�����W51R�@0`�T���-\pǩ��ߵ�P�����a�\^6+F.�L��=2h!���N��$I��}a�<W#�0Y*'�����v�3�֋/�dL��;د�5��ﹼ�`���@~��h�}�R2��Dh�a�{f/4��Xyt/<ܔ�P�H����	���Y��������I�Ȣ����jc1&���(���$���!�lz��A�����!%��.��$��$���y[�� �u�8&j�W�(IM��t�(�Bį2ӷ�>	e�~���t�:��"�ín	�E�TZ��U�l�˞as���!Ļ���la`O�H�m<K�7�1u;���-�5kA"����?���b�J�ϫ~ݒZK+Y��2׷n�}X��ɤ&�C�檳���g��OFY�`3o	N>=���d�/ж����؛S�|�Vڊ[�=�	��t�g$�����o�<�p��P��Sd.����l�-Jy�)ra��_y�(�k�Au��������4���X&50蟎ʪg�d�|�|�y��,�%�����Ug ��y|.���L	�h����97�*%���yEZ�e�oZ�i��'GU*^Ӆ�g��]��Wa���i�a~(��*��7�O�μ'�B���uP�=w�2��ǘ.G�"~H��I�R��;�p�-2�	z]�>Y:�E�<�C r�rDd�k�F$QfF������CYh�� �|-�N�F��6�f�k���У�v��(v�sUo�����P �F�/yZ�����Y�2�L������Q ��(�� n���z��]��\@��hg1���g��v��̕�4Y�(�a�=�)xA����jۭ�8 #H�M^�+�Y�����1]����
�.��z��#ނ$V�}�+p�������#�;�
ziڵ;T�O�>�[2)V%��8��Z��<��`X���G��h����@�0e��u|%TJ�1J(g��[,ž���n��`��ht��h�$|����L]߮Q2�"�2���~�cjIO�MQї�Xnwtt����E��}#�>k������������,���nE��C�מ��
��.W�I����{J�o�R�.G������ .�Z���F~�#� �|�Y�B�E{<������EI@2�����O�'/S$�Ji�a�!�6}ڰ `��'a�&��Bv���������܌
F�V�>ݝ+�(;?��G�p�F�塻������  0mm���D#��Y
4=t%�#���Ui���7��1��[�d�J/%��45�Ɍ�d��j�&Ե�	�0+VY�g��'����BW��pҔ��y
�^�}����(o;u�z-ֿ=kLd� o�t����-fG�v���6l�W(պ�Z �ħ�=�HFWgO-�
F��$:4l�OV�qĭ�i_LCO
���>�n8e�4-T�*>�P�Z��s6y���;��5F��3[M��̘���B��m]��h�ubd�d���t@�*�Ii:_yls�}���;Z	�o��r� \b85z2S���������Ě�"(&'��y:���ա��:�0�4 �(�c�U������?u��1�Q�5��|�F(��{�m�'���4��74SS	)3�AMr��k�>�[��c{{�l��>�?d��h��Cғ����l�N�����HM����(�h(��H{`������k؇���������4��-��-P钝�O.�\�� �k��!�K�Cz�/WV���ɟ�����fT�A
�V���e�`�o��2Y�e�B!�hVb�:e�� z�e�g�����~�r���讝vނ�������y/�s�r���w�`w5J����(1�N|��$�F�M��	���]��as��@nA]Ϊ�!� �Y�W#�v7$+��x�n��w��\�#2S0;�&�_�Y16���9�p&)�����{``�r&��Ю$���rIu��U�UuO:�g��<
��5*?��t�L��E7����ν1��q�÷#0����[���A�8�wnr�SU���U�`{�t�փ�`*�,M�k� ��v�?�kgq� ���df��ch>�P�<;��=�A(��շD=��U�<k�*���(�'����A�oj�;���~r���~��G��awWg�9�i7��"��`Ӹ��4�"���u�_�����>�Ms�ﱖg/nN�!��yP���a_��P���X�2`J�'~���0b)-(�*�A��� ��˚��J�
����W�P�^��l�Vi�J�	�Ϩ�_���n#��&�P�^<��m��Wޫ����y�􎼱1u]�װ�x�����Jvߊ�{�M�'ɧ�r�:/��%]Q�����ᐠ�F%n��;O�Ƹ��ӧ�Ku��Iڝ��e��`f��C� ��!��L����Jw.�ND"T�HKi���}̈Db���[Ւj��+k������*Ŝ��C|�g�\�Z��6O����Y�v��>�PR�Ek�U*�;@_ᵓ�5Nj�����ec@q]ӽ�C�{
��	Ӓ�PR�*���a���Ξ���8�k ;H����� �$"_0�R�F�\����\S��Q}��T�BdO�M:�-�����dR�P���Xc��XS�� \}�$ߞ������:xeW+�{�m/?�`��w���PL�2�s=��t��k.f�������?!�z��ݒ�� ��O������{�ݲ��G஖�����sf)�H�3�"t�' ;Pԑ������Q��!��q��UB��r	�?�_�Bk����#l�=YՑ2��A҈�e��u
;*S�s���/�A�j��[��z�Os�i���?�,x�}��Tw���܎KV����L� ��-&y=�w#P�sB�+�1�`~����	�h��%Y�͞���1F��G����;�f=^�3��܂97}
r��$��
lVPR�%!d�j3Z�6��VF1mV*"،)z�'�v~-��3���.N��v4��L�\��D�n�r�v𕜜�E"Xz|�?�á����WcX'�*j5����� ڸXBӕ~����Ą�w�.
��;��i�[��ڪ!h����^5Zs��e>�!�l����G�aZ�G3 (�^���(%�I�0t���4���N�.�~ĶJ~QH�q���_����bP����g�U���d�	K����S�7!�|S�ʭ
�A6��#�q.�I�FG<P�"�Ǎ�z�KL>WB�5�*�ZG��S'� �n|o��	M�r�b����,nq�䱧���z�.x	p�cb&�n@��
K%���Ҝ���U���7e.��؋�:C��<���[��K�$,�K��X�������n�DH��Z�!��M�Yy7��� :��=C�!ғҞއpH��I�#>wDl��ã��w�8��W�Z���w��N-�\�u� �g��";V��7���m����n9���N�	�[mR��ZR%tٳ�Gf�B�)�Iz���g��UQ>��>Y&��Ϲ7I�9������H5�zjs���V���2H�{��jF��t�b�$m�;�&F���{�1�u��:l|�B���cMx�n��� �0�c��z�]�v���_��h/����Mԭ���>���f/����8�T��=/U��T��4��T���*�2�l�x�'��m�� t������d-������rKDz'�����������3�X�`\�c>�n2��RGK~���S����J8nM����Δm|���)vIG��zv~E��ؖ�܊���d�����p�B�J��~��?S?/\�=*�~��$��(�՝5M%���Y��Y��7�6���^a����[A�r�п���q6b��R�=hs8�ku��Mr�R�.��`��=,ϕs�I6�Z�Y������^β�k0��+�7�ቾ�`+z��"���:ˉ��b��g�I�Yd�N� ��ᐰ/���q�=�����s�Һ5]
X�>Y����^NI����Ñ�+2��Z3\�.q�)A�Ǔe|����N���A�w�]b����N��NOt�O�/'ӟ��蕯*D;�"��^h�xD;jPb�`!E�A���<����&�GC�!���ף�����q*4�g�IL"`p)݃��{��s@J�LiN�ڏ�z�`��U"5QB��e��'����Ǫ���4}Z��+2�QK\���r���>����ې��1gS4�a��fK6#P��R� �o㏎���_�j�c��n �sQP����Z}8/���WE\�@���@"�dkg�aϡ	����@�W����!���n��Q���=���;<���Ŏ�)~B�k�n��yt���w&f�Hl	�t���|�����1fT�Z��Tݷ�b�b�&������<>����T�i��c�+���.����M lg�b�2B�	���`���P:<^˰x�C�*��.D�M�aW�3x�ʘ3S���M�؛�ѸV��cלnl��Z���������PSl�ʨ�H�0�dh�g��K������:����m#��3 n��G9����"�]�J@��ӯ=������j��n�T���5���GƶE	`�"q&vF�%���0��W�
�x��H�Ct�L����f���4_'�0���>
�tv#�(� T���*����	������ 6a9qҺ�l6I0�mE�V�y���d:�2ȇ�A*���	��������Q�Ҕi`هgz���Ug���O`3r�v�ˣ4���ۄR��� q��r��EꮲG9zmP�A��Y(�o��}�k�c~�^aذ��R ���.�H�e�X�Gs�!�F�X��Z�g���9�,�������h%�`��4��K�&����+*A����x�	��a˨��Χ�`��8�~TA�ܞ�Q�n��H�[�C���_�ό��U��3����Ɖ�{OU���sTXj1U� >#B��`?iD���-{��B�W�7P��]��}��Az
EI��A�% k��	I�%����C��2K;����Ȣ\�]T��>Tƞ,Ϊ�;U0Z?
k����t�%��4�U�F֩ u�t7ܫ�AU��4��+�9������-м�j_��B����