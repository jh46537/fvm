��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{ϫ�*#qxi�6f���z�#JA3b���?���f����>7�+�������9ʮ�����������-&��!Hì_C��X�Cf�F#VDJ8���Kޜl�zQ{�t����!�����K�z�3Ek�L
��'��O9w��G�d��n�s�����rG��+�t�[!���i���o�=e���)ا�߅�U*�X�d�/,Ԥ���׊���<�TLF/k���S��U��BD�;�+X�*�o�d��fȿ��h������ ɓ�ķ��i��@X�m�+^u�7I��>��ɧ(U&�Ϸ�&z���|��{�gB�f*r%=h��A�6���R	�86)91�I�1Q\�o���^[_�BѤ�uH)�|�R�zɗ����QXxU�2��l@����;|>�<� ��Ǩ���Iђ� Ź~LN������-X�����	P�3�6a#�O��rz޷7 �dT%���
D����V�cB�?J!|)�j�x!^Ш@�~]�������^*_YD�P����Sw�ё��Rk����Ě8�v]�j!?3�Ea;a��z8?�}��^�}3^C</�ɍQJ���Џ�$��R��C���{iHjjx�pt��D{ҭ��� ���!����:{�ޚ��0����6pk���L�H�~%��zU<�nˋ�4V������~�	*����po�^��}��
����Ʌshs�LG����~F�yw��p�C�M"��5:��Y���^bʢ��
*Nx� \ ��e���T3Tb|U���q��)�"-vb�Z�NT?�HK2Y&��.*CV�\�-��<�A���>~ܑ�ԃ�X)-6j8��ٝ������S�3�g,;���C=h]K�3�q(;��`�&�b���9)��/ٸ�7g�ơgئ�M78�$�A������ 149���Sram2Ŀ�ކ�`�'K���.��$�@��+,*�Rs�F�ݶ{b�R���,l)^lQS@��O��kJ�m$綫w,F�J@����͏���a�l�U����2��ޱ,���m�:w'c%��`�4}Օ_
m���Lu�
u@�]�⮙�{Ⱦ�{�@~@V]�L�"��_������o�ͤ*DḐ��ށ��Q�aU�:�D��I�=6�ʚ;�b�)��ݎ[�AigB��Ӧ&��M��ND��j��6�5�p�Θ� �d(�*eW���qj��G����3���.�߁@���%�v��?��i����!vsa�M`�bQo��o̼c���=����Y
�H���,4�d`=���k�]�c�}&dK���k�O�ϴ'�fz1�/(=�����mˍ�`%������23�\���l�"�
�">�A��Vꪾt83	נ����"(K��]>dJ�-���T}�A�.=���V$�h�Iz��c7;�W�p1o�	$y�6�E��F��ŠI �9��6�� �@c=��^��:n�ZZs�/�,|��?c�/���C:/�P�#{�;���q(�uF$:��gJ��)���3爐Va�/ޢ�]��=7��q\�Gͤ[�目W�B	��{r`c�|7M]��B����
���`j.� �U��x__P-�o��#D#���#q�����>i:�,��jz}��|����W�����<��6wzn �d���0�hU��7���M1��.�bD���-(��@�enP����X�mz��*��S|+��I~j�<����T����0�7��/9p4�^�D$:!��m���x����zse+�L�{^�Ɩ������O�����:~o������.A�GՂ=^�^�
�"�-��ɦ%6̱;W�I`���n�"��o ��8���G^SHn�{��ǉe�TIL���ӫN���S���pt���Q��,+�@��� w�/�o03z� �CK����V_k�-�'T��4ԱG����-�/F�6��̦�׾}��rן�x��EkM���D�˓av�:i�kSˑn�	�өTu(`�)j�+�k��3��-�fR@S�p���I��������e��sa#���*���U�����a0�dm�د�r���O���THt.����/�w����ǭ�=�qqJ֣��� fn�:�������ЁO,����LT�4�s�5'��~1�U���
=����.DG_�_�c@���pm�1�*�i���*��� �!xG�t�{�'���5��"WH_�V5�1�A}�.�ժ*iB�d��/��z\D>q_�:�1t�%f~k}�N���T}l���}X�������uAK_�����M���AP�l�|�sep��]��&ȴL���u4,,欍S���7�zQ�Ϝ�JZb�S)k��X0=uۗ}�?�-j01�G���F��w�t������S�,c" ������S��}��P���A\���^�]�D���GDU�~���Z���5.d�k�Il�J3X��Zʞ\�o�L/\|�8��)��E���f>D��zIj��5I\>HRmu�я4�HU���D�R$R�5I�a�����Ʉ�^�����Oہ�&27/|��h�U�P�1�x�4�;N $FI����"~Շ��}�Xȧ�A鯌��s�T2��j���H��[�I����9I�2Dz�q��\Q�}���!fX�rn~"��I�A�,]*9t��]���	M�b �4z?^S��N��w`�/�Ď��Hr
wo��3'����M� ���[��s��ɟ�?2�wjn��.�y�L���$�!L��chC�[��Z5(��}��t�.�F�b�:>�N�4�$'�b��VKY�����7�{1�g�ז�m�?}�4��<��n����OzD�g������݇ƶ:����#NIg�iogrxAO��EW����>�"xߚ\5�9c���KJŦ��ؤ�(
<�+���+/��@kp4o�Iy��Po�I���q���5�D��������~Թ5)
Β�-�Y��F�H{{��K0(W3ZY�G��MHڊd=���Ͼ�g�[��5��w>�