��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�u㎺��` }
.uJ��@DJ�_߿x\b��tV�./�������3%���d���*��5q,�S��I^���.�%�<~fi��O:����\��=zg/�҂�[�ˎ��sא�&7�	�'��W��j��$
�-��� ��'��c^���[��Df��BGa�����6��D����.L��R���` ��D��_lCӪ�B��]��N�]f
0�B��/Od撕����3�y|G�۳J�e}���J�:�Z� ��_t�Ꮽ��d���Y�:}��R$p�z���#�R��Q�p�6�vJ�z�J`LB����	��h�qƗ��8�{fղ���� ��o)�����i��fp��ֹ�LZ
_���C�'~�pm����H��߶>��慕�1�3Fl�p�ƠTrUj�O�{�U�>HaD�g�Q����(X�㥕|�Z�8DUcj��>�ώ���T �I�i9y��0
Q�f��=�CМ�k��j���B�-����rid��M���Jqsa��82����z��񫢪��2��O�eof�jt��������C�����y���w��ʁM�|- si�����KH7y���\�c�wd��2;��ܑ7��>_�;!���ww�!����~�d���$�E�:�u4�cn�X���L}��h�J���7�]y![mV��,5�I�ngA�����w[V�a��F"ѩ�ER������m)�B˾��%XU9q]�坁X����J�L�5S��ϋn9$Z�=�4N��������ay1�۩fН������܉�����JYv0Mứ^��}���T�`�h,m�+&�^'"�5�K�T�?��0�U�lU��٥,'�� 2�B���jd���Q�	�T�d�F�)�M���f�������?�sΉΩ��>g�[l�۾�A�M|��$�%K�W*�z�f��b��D6ws�-�R9v8��R:~���ml��e㝽ۢ怃d���cT0*�{��@�o=������`'�C31�r���E�wx�|5�M���)��L�	]VF��}J^k=a	��v}�jW�������g���Rc�-�����w��ߞ����n�9x,1��X�%B�}���$�0����m�X�_�u�=��5�"֞/�Z'��9�����W���#a&Xk�>^Ƹ\~��S���\�5��g��|{��������D�1n�Ɵ���{aB�V�g��G�m��ȶ�%�T��?|�|��dT]F\��,Vs%��=gfQ~<���2"�Mc�H��և)�i��|���1@_PYZ	�f�u@���4V���L6&۲[dhD`,⒜�c�h)`�q`=��PK�&�C5~\��Ԧ[�m\Z���IO��n�ӿ���ne-*���l��^�Ezӣfl�q���݋�D~�)�l����-���~j���(���*֬�����?�-�~ϙa&4Ðw�^�	c�{_´^ҳ���b�MOH��N��u*W|<�(z���Y�y�|��f���m�!TxQ�Q��!sQ���7�4D��kh\$���Yw��fշτ�<�TB���yT��D��Ή"���٩ϻ0�G!	'����2;�B�ί���(}a�Y���;4*�Q�|�-��\~FA�h6��7:�ςͨ%O����qz�}�3>	�q��ۜ�4X��`,bKIۘ���}��x��;Y������Kڧ��/?���'t�޲YLǫI�i�a�k,�QH�Ћ'�u����b/e(�eL�v� 92y�x��>���h�7i�M��ePJ�E�*�6����э'���I/@+V��z&����4���m��K��}��.Z�e(������y���eԅ��3���w�~z��`���x~�A K��G�g��
��A�0�2�b7p�ȅ�&`'f/7�Px�D�ڟ������W�oE�3>�G�\<�!����Ƶ-l����8F�*�>X�{񬿬�c{�(��a��~#W�N������zjT���?z������Y\���P�S#2�l%��H�Q���o0�K"���p�g�N������P����▴أFm�e��Hǥ'�������m��D�Vn��Iѿ��K[C��W���
Hh=+��(D:�'�LI�^����ׇ�ΰc�9E3}�P��6;3K�Dџ�2��&F�9�� ���+�/@�ƙ�c(���$���ff��8�p�xB��^�N��P�˗B��J���d�~�:W�}�$@�`(0W���m�B�/51p8�'N��Ǵ	��oޭ��%�*֜�癧���CGBZ��z�!�*v(�=i�f��#���+�`���їY~��������(f^br���D��hN�*�];�&I���L/=�~��Y������$?l�\��^�E�>��=6X�0C�v�gȾK��H���o`7����ku\sͰ2}�cns�Լ]����[���m%9t�����!��w*�`�,mGqk�L.����?���xoM�> ��~{�j ��L�`��G�l�
�bDΣ�u�=x�V������G�e'!84[�e��̙���(�`���ܱ�M_�S[�l!���N���y�������o��u.ZtުK_#	����\�{��3A�����(@a��!El��I�*B���A�a-�NFښ�Anȳ�*�������/Lt��C�w���P�F�!G���"{U�8��I�|���=�j���t0q��<�EJ���(��bQ�3L�ِ�����3���0��w��zvh�,��v�Za�4A�H�6���i	ߕ�Iנ�v��'T0A7�~_���	���d��\���&֊�J��?x���˷P�s�T"3��0gy�BY��#���	`h��{�2bʸ���e��d�=�^���d�d������g�.]9��F��P��V�ՠ���qt�T?|�ӲZ���}�Ї)�Y��ª�j[���|E��aeÒ���:9�l�$[���/� �x�л���������{$#h�2 �,�׳?h��m��ҿ[$�y#�ڎ�t��G|����%l`�-̏���N�?��	�Ա[�{y����ّ��=&�A�ׁ��4}z�J���7N-��p�]՜'���b@ꡟ��(��1����F�3!r��������a�RG�I�W�8�,j2��r������9��]L�a�*0�@�qu�4��-�'iۯ��!Ebj!��5l��K1�jD���>�xF��ED��h��FF�c��E����E�g���~rIʢ;r^#��4���Q�ANO��ou�k$3�G�B�����c��?qG&�D��i��� �s^
C�[�:�/}��?�_���;=�u����K��
I{�M��[S�ӻ<�}[a:�x���	2��o�'�����`��X�=k��a��Fv��?�a�qd���V�|]x(t =�k��q��.��9d&tT�@ǘ��ܼ�R.�"���.���JX��8y>���Q��`��+�I7�	�s~�3��[�w��+�i�XɤI����4s�'7<�Z͡�M�1�a�|H�g�)��#z$��}8��wPj����=�#W����-y�2�^����h`�4�/�i����l܀`�l1�'�F�0/SV4���5p�H��3;�QU��5�0��+�Q0��kȑ�˒ujr�}��"޲������}9j舌]���DѳԎY���&PP@�������>����#]�Q].��D0��2ػV[	;x�ĕ=�ҝ�G~�l����ۛ���j$a��)�`���cS(�z�j)����`�vN�X�ұK=����ᐴ�K�f��-ч}�n��4��̕U�!]�Ƚs���E�FK����	�0{w�seP� �x/�!��D	�����ȼG�i5�X7ċ�]��y�y���l]���"���m�����)�@�+1�D	D����`3�%?�g�h|�Q�����]]��X��E�_��% �Ȓ����)�Xc�(v�b��w𘍀r�g��_(�C������ϣ��"��zM��HX��J��C��n	Q�-��a�=SN\y�eH4)Y�����Չ~Y�XL��%�{F��Л�VY	���Z�e 0�D$�\���wi��g�7y�Ҧ�<�)�w4��'�/I|�4	���[�<�[�VUZӺQWk`@�� �˟�QK���<_�Ϲݣ��]��㲆����UvbP�\��uw^�2(�KN��[���-���5���� qh
!�*��G���5�Wq�=GS�4�W�To����6�w�|; ��s 9@�t4�o�,:�%�Z'�8D����\a�P�qĨ	�ɻWT��XWI�_���>��J�b�1��p���c\'�����������7� 2	����@�%w_m����<��½JT�ˆ�CZf��Q򷖹��FĤ�V�)&�P���ّ
����d��`�Ֆ�N�C�B�g���Ⱥ�%�
{q�bi�G��u"�������Fpf���`�;��c#	�X>KAQh»<]z����y?d�ydg�.��9���(c&0��8N	ԣ��d���w�ux�{r;��D������C9?� #9(9ɤ�xUZ{��u4&� itK%vW X�'�����	�JN�r�l��L�[Ч� ��µ���~,>�?{��5	W1�ٺh��!>ޜcW�K'��[��z[^�W0G}?c��Q	O� 1���k�C�C*�BrKt:Eo�q�� �t��ގ��B���(//;l]�Ɩ�7?��K�.]��S|<��<���<��d�	:yj	���q
k�2��X�u�B�|��3��;ay°����#�QO�(��Յ-+��5P��~?rc�?��֊�7��*�^�_� �������q���2�D��7��0L<���Y��zq#衑�;F�vԩ�Ho8��H��g�1v)_��1�H���6$Z�o���#�tT��ꂬ�1g�}�}�?b٘N H#�����ް���j�CZ��x�C� l�4�t��ڡN�R7�9�JE�����va��\��uz�M�1�8���E
��K�ƕ�%4��)��;���:B)̠�IL����i\8�j]L�1�H��	�WD��:���G�GMWΑ�#��-���J�mڙ�o��J�\���3*,�����,o�=~�&m���X77̟�!9ł�.�3���v��#i=Ei�0U�!�Lz�`#�,�{�cӒDFp������o��3�	B.GQ~�#�#FS3u��E��C��S"���p9������l{o��#�i`�c�f[d�pO'j�����`��an��i�՚����z�-��无FO:/���B5��;C��Yq�ž[8)b�:^�Aa���2'ڞ��}�����"=�Z�M�8�9W�?�{�������%,m}Mj�| l������sXC��~A���/5C�^�h\M�6��A���	)c978x��w���C�&�9@f/�C��7�����%H/��ʪu�X�&W�0�s"��1N]�p�����M") E�0�������$�䧊�n�P~�o�u�d�t]%�EYT�m���Yk')I�ٙ��1%���)�7��3+qI:��h�J�$�ʼxy�b��~�@�p�ڠg/yU��%@X9��ǩ6C ����8<���O�\"�&�t�מ=[���~(��#z�h��եb��ߥRNC���X����2vN�X߫�5{��A���A�4���a�:$�A�+�t�
�'����k.���T �G�ߚ#�<g�X�	�N���}#�r����L^�:S��c*ܒ��`�$d��ܰE��Q��3�D$�k��V0։��KԵv��*j���)�o��{۲��P��eA>?�J��&������W�XA
��e���{�۳��i����1'�<�K��-~�J���z7~kl��U�r�#/*fz��|�vD���}�9�,@�`�L6��$���7=��;�r7T� �<7R��@Q���K��D��L�XՆ��J6P�!@L�L`KF�'�F��R2��B)F� n������E<3�+��Û�%���I|�Ã�Ǉi��e�/0���]^�{�ۻ �L(�oR������ǂ�4��W!6uN
��^3��D� �����xG}s�ů۶�M%�P�p��t��J�J��K�ۄl|�m��=$q�-b�-=�ܖM���a/v�g�W�5�P���oK@�V��-G]��^�KFm�E8��ݥ'����it�I�m��F�4�ŭv���QVH�F$�%"����NÈ�d/��SJ�h獓�]�Y^`�|T�����Kn���m�b(��>��Į�שD����ؖkC�.ɮ�p��b�Wٴ�U��4����S)�=R��GA��3�P)�)�Љ ���A7�V�	�_��m�)X�)�D/{
�h�?�ۨ�y{?�y��X�EW)g�R��6��Q@��)��]�X���n��2Xo�� �wd�0p ��v��E@�MH(���S����YG�M���9z��A��{��r�)��`IM��mI�(����e�4OG��t��f��S��p�
���l�i��66�rc�hS�(׆��g7:�|[��ܝ�]-�/%���f�Q�������}�*5,�	�
S��w�q�k!�����#����2��=�p~�3�"V��:���}'�X�%N�a�8�*3��j�w�b�"gꊵ���n3���&�X��v�Nk*:����H-f'fl�*���������Q�7n���-�M(��ݯh^M=�@��/!��*SU@=9���t4�.S��sE���âT���8�>���
.]
hW2d(�����	E��K���KA�	�׉S�ȧ{W�hY �R|�(���+O��&o�tXU�-fX�=J+�2���0�/�������ºJ�.ܮY�a�PU1(l�>� ��]�FA��������J�C������y�Z�7�O��&��@��Q���Eƍ�Q/�oˉ�Nم׀�MD%*��KOP�sK~,623��5���G4Ą:��ɜ@�U}2r�Lc�0=�BX<��){�N�uZ��i��T�n����G����Աa��)��	.|�l��}�-ݗ�ut�I
2���#��?�������U~�0��3�>C���!���Պ.��n���\���s`J�����^.�d�aՁ����3#��-Û���*�q�H�F̖,*��Ud8�Vި�љ���,��.���ҥ�vV�ۓ������ö~M��K��H����HU���S�Y��Ĺ
����T�ΰ58<��Q�<A��b��	�I������Co��f���ڱ��Ef�������[E�k�>�<�zb�Og,�ʯWc4��D𶋙�1}������v)$��*����v�-k�+��H�y��یԜX1�چ��L��ڃ�J,\���u�Iy�>Y�O�.:��mbJ���ya���%�J�L.�Q�i!U�Qm����jO�^] �w O�-8OPr�0؛�^@6H;�wc  �*�Ss�$ͦ�A�_zŖ
��?�t�,���x��j^���=���P���.��<���%G@�
���S0j!���e��[�����e&L,�n���� �][�َ`��8Z7��Xa,-�,R�Ə��e����t��8�k!xQ�b�p �[���'oh'�5�ܚѺR��z�5�ؕ<VV��8cl=��Z�!u/������K�[e�S�{&���w�Y@�*�=���K�7�R�)Uc�\Bn��RPsD�zq�y~8��:��d�V�k�TP��}xR�Z��\U��8
�&�b�6�ӟ3��LgL=+P�h��)�!L(�WU��p�����;I,�[S����01�4�j��JY�����6)��+�`��'�j�/��㝌t���G�D(�b�k��r<����.��O=��k֑�����L��j)~���yA�mf����������P�M]�(,r�CۜW��R��U�&�K����{K���/�v@ۏ�C+w8|���s0 "��С�#.[������"UvpaQ�g1�@Z�X��ϼń?�b�������4w�}gq�`]��J�r��ˢ����2�����G�����$�'e��X���sF�\��w]\?r��OW]{̮@$$�>�n≁������@B��H=�>�j8m�����z,��rE�����>��<�s��ټ0��6�;�V�VP���c��LZ�)9W�+��D̵����s25�q��d���͊�;p���f�g�*7�m�T�u�}��hM�4 ���u���1���g(�
�2��T��U�ǓO���(*cj��v"؍��30� 7rFݪG+�줖�s���ƻ��_�_�k�Ķ\��ϩk�̟7��X>oqk.N<6*BM\+,�QQ)�`��.�g gr�D_� ��ժ���s������I�����^%!�񋖄��J�B�[0Q��6+f7C��H�>�B�QU�?H������4���C��'��I�sDy���ٱ�u�Kr(S%�L�W��A�G쾯��ݏO�j�������������yi���~i�C��P��B��P�8چ��:Y[��a�w2`�i����bq:&=����{&J٘&�~�%��Ի��W�A�h K[/�Am���,�p�S��ak6R��l+=���mk DKAR/4^�Po�-<$�/�BA���rt{]��ёW�&5�>���`�p�������s�Á:��F�k=�@����T~~$1E-�K��+A��4�?5x����K�x�Ř�6ʨ���ڵ3��=n~F��������T���z�N���'H�fD���1�ſ{6)���4>U�P"�j�����j�(0�3+b��"B�@��УT�����f�	sn�@��`KWjnѲ��HZ�g9�:	0�芚�s���t&���=�	]���#�3�սi�ܛ[M,U`P��J�!(n)FCv+�V������|<���l5�2%|�%��+��=M��1q�T�	b`w��I����a-��O@�ڳ�rt__L�1A�u4�L@@��t��&ϐ���:$����WB����R��ʄx���Jz�&lms;�Ob�s(���Y�>�����;E8j� ��*Wg;I�-��?�J�kC�N����*��h��MKst�OÙ����VP1.���D�	R^I��>q�٥��hS��)��s�� px����w�:�@��?�*�����Q<�]�X#�r�Ox2�M�'�í��Ă8Rb�"��>�׵ε�YL���p�:�D�őp9}�U�:�*�ՠ��E ���Ti�W���c�B �fӔL�`"�$~�r�Kp-q�ż��� J�2�,J��աL�����t-)����y���-�� �(&8b?�T���p	#s�L0)ečƸIA㧟��?�J�ʆө$J������,e����Ų*�T\�L�]�d-Kz���WSI�֤p�q��IWL���5��G���ʷV����C�O!�G�2V���͵v(M�4�4�(�Z�uj^fd�� ϵ��D&�L��;�W(���T�ݰ8Ol("�;�g�s�����0my�b�<�������R���`�!�k~�t�p��Bf����lt��r�m�՟�v���έ�q�����I(	�f��3핥�
!�BW�=@s