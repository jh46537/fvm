��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�%>��1(-fR�6��Oؽȏ�)���V��L����W�H靠�Й�t�SO��.|��0�M%�}�eߋ��O�	������Dt�!]��ݐ����p�H�B�ݾJ/��\�/�)$�yU
�e���5DI��ka�����!y��u/Cv/��'f���?�����Q4�n戤껁�����o�|�B�������>ܩ�FbH�}����z��b��9�2?.��|��oMS݅y��e��Җ�W=ͺ�G�������y �e�~A(o�����^M�-::���YчV��:Ơ�Ͷ
ؾg���iѻzH|:̠���B�0�����#�,���4�� �'��7�.���L�\j��~���̶sϯ,���~�_7D
a�(S����+(�3'2�?'��AJ�Xk��z}R�Ւ���k��|���*�+jh����?��!�{BZ5���,��n�`@PTHxǘwgU,=O��0�G��f��Hu�(��c�sH���?8t�ǻAo��Ϩ����1s�Bx���6�$D���(H;Xh��Y�������t�������N��/�q�X�D�ex����j���d	]��n+��4�yQ��ro�E�a��ӄi0H�^���S #��	ECɩ���0֩�����[�WG�����H譾����1��l���ޏ��O/,�Q���@������L����ao|���y�D]�>u����6Ϛ�OGW�������}�>�1�?�k�?
�B�]{�ZƂ��:�]������v)�e��_q��k��ru��*:;�,2�!���j6�~m�zP<Ly���Q��;��֖�����>�P���T���ʯ��|:��ʝ�{�hV��ʖL�U�{`7b8�Z�I��?0���"l����`iG;���BI�k}~�+�$w���x�he�>��/�C�Y)�o�޻J��ȶ��x`9�5�:�����g�=�ﱋ��Qr��Ƽ>��o��;MC�cwI&]�b*(}����^W&b^F�^�)�"�R����ˇ'��E41/eFig��:Q�ÆyL�w�����+��y[�a")4��}'#�M�"t��.�h����=�ձ�GuN���9�]��J6@����@��n���ǈ����t��.������1���Bj1�������Ő���Y��2"�4%7F4XiXI�?6���V}/���ȝh�s�^�[�@ (9�]*����6,C��8ĕ�qT�Z[֯�� ���+��#[g�\&�m�% � ���ί�(���J�)&b�ܯ��5����Cs���x\�P��U"�q���X? �����- �Ԫ�~�ɭ6j��7f�%��!_7g	@�c�=�"K���6��&��q��nLe
��\�ԝ2L���V@��w���3c��ӕņa��z�TL��w��:x��Se�P���Kg	��(�TjX1,I7�R�� �%RaF��p�6��4���yj,��x���y5�h�?0X�}����N#f/]�o"�{�sQAy� w%�*�6�s�������N�X�&��U�p	)�gbbM��r�Ǚ��F�Kh<A9
S�a�wPH�������&�a�t�kY�8�6=i�H@��/I�EjF�����X��z��G���%�u���7�q�UP��)z��0�PȭL�z����$
��K^�!}V��j� K����v��U�Π���^��_u	��o��h��/���m��s�T0��'2y�F��`	h7�^�+0���We�,����Nf�h�űC��������]�O��B>tA+pG��h��/A��(�ӑ�p2r�U�O~S:�����D�*�N�f�E|��^�C��,C"�	o��ة#��Ȫ�yhSw�پ3SF��Z'����`1�"�������?(�g-X�eIv?Ϯ?�:V����ȒU~@݌;�1���0���wR�4�@�1�����	�Ҭ|T�~qi]8�tt6�M�L��+�2J�5�G�F�}$�z�D($�� FV�𐚲0� �T�)h$>~@�Q����/׹�R=�l']�]���K=1uo2�b�D�ʠ�x����䯓�D���HW��2����.I����ڵ�,��u����k�3�ǘ�T���QƵ����}�	�ܨ�7�1��i~��v�K�Ͼc�����E�ӗE�+M��R���V��J��9�g�����E����P�s)�g�"o;����s��h����k`y޻$:�&��7�W�ݪ�����̗�Y�h�NJ�c,�Z�;l���WLE�W�{��W�%1�$Q��اYi*w�F�d���?83qL�V>�Z�w�ӈ�7�	^��\m\C�R�/�P�+�;�L��0U
�Q>���jRw[[��K�`���������;�X��i��Q(qU+�6��P��5[�
3o���nF��t�ԫ+�N�?'�:��K�mO@ �c����+V$b� �n�����%�4­PG[c�ۀq���8,�p����1T�4|��J�y���j-<���t�b�;�pl�%&<�[�i�'�a��ԕ�.�ŽA�Pz~^Xh�ɽ����?>ϵ	o����L��F�=p��C�be"7�юJ��I02C÷c
�o^�.L�^Lc���USk��>�
���P�|�%V����A���P#^(M-�i>yWBg�p��ե�&N/����&��D��EU��� :?���}����yۦ��F�|���}�_v=�D	[���jK(��J�N����7�6�
J\U��	�m��`�'{q�tgA�;EJhޛg�ʒx�eJ�K3I47�A�!��	Kٛ��C�!6i	��9��U�^E(簹�a���C� �a�3��Z��V&�셿�����N| �f��I�}ϥK�w?yFa�� "}�M�(�g���Б�ZUXn�����Y���^�r����ܽ�}�Xj[��R�L�d���#ωyf�/��/�� ���Б��R�#'4{�X���M��JЊ&PeV�܃����n�qrGm���))�����j4gDa�����$�#""�^������H����������a݋���c��f(q��k�����%��������brw8��5��p������Gا�������9ACh,G�p;��f& �!W���d��@���H�
������q-d$Z����s{�~&�~�
aq��B#�H�`� ��6J�>������1�/��Wx��MWxMV�ȓ��OD�K���ű� ƹ��gJV�I�|�s+�E�b$AI�қ�`�l�G#��ѵ�^�� ꋙ�Qt#�x��zz
(���.��$U��Wal�ܘ�	�6~7���פ�/'A��ǲg��q��h�9�@[P��0 >��`�s��y�р�s^��gx�Y�� %5��{H=��'ɪ��E�>�Nc{oJ�C�}�a�ީu���F,T�V�׀m�G�+k�v�������+Yâ?��r�*V�{cp�Oo��HS�˛sn�����_��i N�y�Q蘜��e�Y9��'����+�1��߾�+�~wx�BiT;2U��- ����ŋs��	�Oă�.�w7���TzJ=��s�M#�_R���U��æ�"�{�j�4�#�s~��X9���	�?��fj�Պ:9�2�ۅ�G���uź�ٲ�\ZR\��`&���n!��UCrB��d?C�_6s��� *0�Y�pz��oKI^���U��f�r�������2)��kA�껀
��Y#g�B��y�C�W9���bA�D|��FK%t9	��_;y��7oQ4������!3�j�[s�r*4z��=����=�]�Y���Y� _NB��Kb��][�}��IQv�!��W�ng.�Ц�6�4�`'�?FV����2�f� ^eɒ~B���R�=���w4�&R��wm6���(ɠq�D�@�{��]�����8P���	��/�Q;�4�+G��������o��>v�؝Ԁ��M�<����G�&������:������Bp+*I��WG3޶,�B;]�JO=���{���g^��f7�������F��E�!� '?��Pc!��fA��Y@I�J���??:���&n��)4���e��Is!���+���V�4dl0��5M����߼dX�L`F���wֿ�y�H���\kD�K�F�c��W�p�ڽY-\'c&�,҉��䠄;[�����[̾ɋWe�k�/=u7���!�:J7?I7�ns�WN��L�"�(ϴ�:�wmu�$��|m0�jU`�Ȍf�̈
�$A�؟�g� ����n��_BN�'���\���R��#�~�q�N9���a���D�h�J��M?}�<mO�_%�]Qp,(r�u2��q��S�X���ɢ>�0s6Ύ�74�o�A�����%"�S1�Ct��\k��A��jʛ9���(��_�N򄛴��vw��'�2�֟d@�=	�5�#kr��P�o�VϗԤw��P���l,4ҷ�D��j�L@�jpݞ,އ �z���J��8	��۾>ϗQz��U�_��o��"?&T
<�����E�[=7�YmOら���E�ĥ���p ���5�s�[2MF�7$>b���BCӂ�}���+�ދ"��3��4W�w��hZ�������zZqE5<�EC��S����Q�8��C�u�ˉ#s`����v���L�:D���G��Bf�ѕ��?������������l��r�c"�"��,޷�{v���!֑fLwu�`Y���Zam�%��$������.C�k��9t��pKj^0���+O��*;���B������.����R�
��t���v\�R���5��a\�6�ԄyJ�cȌ���Hl�:R�Fn��Ը��~�F��E��1.D�e�VR��1�������85{�Ņ�{��d݈���d�2|?
q�<��doQ�+�YZ�1��K�g���b�3�`�pk�B�^��|�
��O�L�?�pO���@k��|t��Fm�>'n�X�_g|�W�&2��a��W5��HK��2r�'�O�|�A��;F6�<`]x����E@j����\|�DA+(��m>�$;�b����֏�A�;
S��8���>�ȗ��󠠌]�w"� #�D�wI<��w��b��n%tx�By�I%ZI�� ��`;�Q�D-�R����%�'d`y=`�Πt��E�����6y�sV���Zv�;��q<�o
���&mS�ɻD���J��r9 �'�TW>q��'s�0 y	�oq-� �^Wc������m�5��s1����߷'�R��H�	�x�دW�u˩��L���o�q����+apӈ�^el����aLp�k^qZ��(uDLk�x 49豟�a��HY�Jwf`�RP�jf�v)?+�m/�(T�Q@�6