��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B����d��:$�馈����Vj P�d�r���rO4�`O��A��4�k�Q��)k���E�Z_��r�Y��C[r2ҖUg(���`�S�L��Ȕ`�?"F^���w�r������m�6鿜�7��~} �(Ĥ�n�Pe��	 �cE/�ݭj]x{�s=�Q�BQ��T|��-.Q�p��.�o<��A��3���$���'9��	�"�.M����(s��?x� �'K�S����� �kfI�Ntd�J�G�1Y�Й���eRo��@�*5�g�!�M�l���f@�1�&fZ�S3˶凨�_����E�2q�YW|���"��,w�	L���J��N��H�m�rc�O��k�#���g�T	�@y���c��v�Vu;O��h�ʆ��gi�	[ƁLT}[,�i�,�a�WC�׸��Qf���S��/�����|�c��TY��S�v�Xp�z�)h�g�gb���ҵ�9д?efZ�eBp�x�$"k)#�.���{����ZΡ�縀%u��"N��S &�l#�,=��#��M(W�n��;'W���ƴ�.��~t��bS̝I����?����1(�+���\S.��Cjz�� ,�݌�DOX[	ɴ[�PC�O)�%PK�io���#��~�����+N9��Z�UJ�Wo�D�7�ԱBY5�O`��!�V�Ʌ3�v��i����3��=�~8O;ϡ�e-������s�x�~_�ί4F֖Y�z�ޘ����� �z��(���[|
��'�8���C칐s�<T^c#���������m��5srBg�W�������s��5�O�tec���Jn.yE��9:��IkPv L�,��;Ni��Dtڍ��Xvb�R?VNj�(C^I�w�V�?J�2G�)�0��v��|!�O���3!-򽺪48�	� Q>F\��x�zk��� b;�g�����ZP�_�
�������ǚ�bW�&S^��˦w?�[�t����v�h^�|�9u4�����r���ǚ��|�F��/�d�$Օ�m��98�ʻ9���Hd>�D%�_���5�O������"�cс败�(�_u�XAR����K�#zo���K�'	��7����:b��X��w�<��%�W{ؕTg2:�A��R
��� /G�(��Pe�Y�(�u���\;�����g��a,7A����N)G�N�.M�Y3M��'hD|�M����
$�*;���2�ОγV8�
�H6�����K������U��j�0'�����^��i�$?�j����9?��3�u�9���8{3��\=����=�CK|r�y9p��� X�VB]�W��ɜ��Z���
����>��)�Z�o�"�:�C�z($�y�[��D��	~�����}-��mM�P��G��u5�r�����������ࠬ�2�W,I�wXa<y���h�.��RnC9%y2�������U�bψ$��п!x�4j92�3��I�D����F���>:��3�k}�}��]��ŌZ���6�.d���z��\�d��T���;�8�V���3~�EU�K�s��q��~�\7@�y؀~�����TOտ���׎)�+[�[�к-l��� !��f�fd�>���`��g<��O�+�\TA0(�{r��k�=Ei*G����$��5:^o��`,�r�|�%��,(����^G�_%�6k���Y�<��}С�k�E���V��ޱu�=�ҭ )��H}JQ��9������H?�D��lK)�o�dX![?�����-�2>ўzԇ*`����9�\U�w
�1|����d���9V:�K�+��h���0$]������p���Q8��.<�6��kD�][T���b(������JG	r�d�y[Fw���mI�]+�WR�K֧hr��@��l�ڵ�]cF3N����>H��A���Qm�/"p+��e�$�d<XlC
�!2�cI;����F���{"��7���^�Q��Q����7�Ç˧YowCJ��@`�R�L�Q�ͯ��F5�4�߯�Q��Fgme���ٚߵU������A�?��NuzM�i�+#�� |��[7�`G+
���I�j�7tƗ���M�nG�㧡vuHe󚒽�{2����
�{�d��dP"E�{|%���7�,*����]�3��Y���S�z���w� �zP.6�b^���ט�aq~�2 �����W�� f�
k�=��I5w�k���%،V��⡠
��_�5�?m�[�[6S.�IN��f�l��z������<^��f�����b�X�K*K}=���9�*�2����UeA%2�r ]%>w=�u��lUB���2�����yA�4��>o�SM�o��O�O9wD��H^E��;�.փ�z� �v��[>�.��Կ�6�Ǣ�;K~U#��>�B�����R@zc��Ĺy�B9-��'����U�
}¢���B_J��.̋(뎨*�CX_�F� k�f�0#1�B�g�o$���H��	����Fj���UY����ۦq�<[ן[�����&����w	�PC\U�� {�j �N�'��$��ll�Q�L�4�����:�ȯ�ܫC.>v������U�X߯�����~�Ȕ�r����2џ�w��Y�s�Ff9G��t��}{G�<@�(o��H��=>[T_�1�+l����2tbҥ��%s�����=/bTb���+�����x�+S�5&T-��=�r�z~�ڞ2�|��ƅ�4]�yAJP�}�������+����%!М%4^�w2�߰��l%'̥P��c��an��m�+z��+�P�|盱�O�ֺin
�k���T���ć	M;%BE͂S 05�_y�R�׮ #�<?#�q	����z���E�7��({�i`��)��,�ǰ�決6?H#�;[Y$�7���
7���ab��{�[��+z�<%d�����9��R@���B�k�g#VҚO~�!H�`N��ɲ�R���Ҫw��js
z���K�p�N���NKi�!���9ȁ���:1Z򿽬ػ��/�5���P�N���&{�z� WȈbw9*�F�o�>՗��X���E�f�B[��H�-��~���>څ�	a�n�(�G ���bn�DN�1��Kqcͣ��!c	G1)6��҆a�.�*P��'���&ӉAj�,��k׹�uB�k>[�^����H<�%��uE-m:����6�p��DJo#F��]�Y�����Qf���.��*����{���B�jH^d}ֽ.w������`JO闲�K-f�ed�4� �eIn�(.$�#g�l�������˧�������WV�Z��n2V:�:ao��>PYż4����6�IB։�!�I�A'XQ��4Q ��[��f���Sݟ����`c�T�S4�k�N��4H)��b���C+�-Ig�w�}����v%+T��޲-'�s�KV"���#YR<���=�"Ż9q�����Q��u��*�=C���ߦڊ���GS|��C0+���=�Ό��ip,]p��~ݎ��-	����2�I��g#�_�{�3e�s�jhe.�6s�Qpg�A0�o}Y��k0��Œ;4�w���R�O��0�&�5�����IώB�gE\��2��*�n�L��0PBDN�0aT�!��w@���V?�7VlI����jt�+�1O����)<�0�nWc�x����iXHd`���zb���C�N�r�0g�@��οhR�RFrHA*Qzf���L� �,��|�ԭ���pm�OoqA�)�.�@��L�=j�6��<̤,��y��W�媂��A�i�X�>C���G@eOl%��i���y�;h�ŖI�Z� ��$�	�0���a*RL��g��uS�~�*|�n�|��>~�ҺQ��n���s��>�sr��~n���Me�X�����9�,b!��\��L1fbDZ��Wi� ����]��Pl��̖RV�Z�l�����N��$�էXۣ���T[�$�J�[�1��p����l~�$�4S�֩-���ʦ�
d��'w�8��C���u PG���#�~`2���WJ�.Ed��te�&)����k�3��k*�%y�3SǙo'4Nm���;�?��Rq(%eKi�C�c����t@d�	8~�����T\�Zu!��b��������!���-Hda�z�H8ږ@ �&\��$L!���o������"?��Z:�\���Gi�T;��B�z������ �C$�V�F�c��s���hj�E��������бb"e��Oy��7�O�B���X��`R��ŸB���c�R�ՠ12������׋#�����Xz?��9-����u�����U����tCT
�~>Hx��	�L��V���*���b����n��Xx�e�� A>*����:"�*�Q �f�	��BK( �φB�� 
<u��bh9���;m ΃c�0�81�"�����$)c�z�\)';�S!o94��7 �f��p����V*
sDg�BCI�K�B�_St-D��7��4f�.���O&��՚,gJu��W}Ţ��}B���>��?Aq�P�B�TUCgBֱ]�U;���HE�X
��Ѹg)y� ު/n��]����%�R��@���c {��������5�0�<{{RK�rQ�F\�C}�>��Z�·�?�~&��ޞ�u�/zPGT�4DC\lC>�]���:T��ŊL��Z�k-����d�D����}���bu��$`�k�ӻΚ����������	Z�=,վ��d	��4`L�\)W�J���=�ªS��]B�Y�@�ҝ�����g(@MTG$*0�ع�V�/��W� �����ծ)3~���G�b�d���T���*�B;~4�n7.~�2�h"�hA�@���a" �'��`¸�
ر����&e��V������� �ǫt����m
�U�ud|��n�E���aE>NY���3P�Z	��x�$#?��*M�����[O�[uH�hm3O�r�j�bl��Lj������F� 8Q�}h��;�.Z�f�C���l=��d��RG�݉ҽ����!�r���v9����Q�����}Ŋo,0 8vU�1G��n��q�^���fU��${ܴ�=q[�P�`�V��Bn���l�:1��_�/#,}:`J���#��P�v�! ��7����	_���*�����jF��a����Ż�ޚM��_�t
�w'�ɖ�UklW��1W��t�c�l��X¾2N��Fˮ�4�N"�"B!�G3����Bd�Y`�d>�t�>	�zs\kp��u�)3:v��_m9��X	G(�۴? /��Ŝ4��uG��{�W;���_�j�����b>�%N�m�b�E�N�5�R:��5VA��`��!t�r��@e�:�'��}��m���8�*�>w�qw��"��7<Md<1�Pˈ/
���*���R}k�1+���Y�t��jA:���bUjEL�rv餭����B9�����n*
�onI ��d��K#����[�V���W�-�j�= �8��}#��i۳1m4D�c��]լ^j����;(���M	��1Z�,������]!=�P ��L1�����z0�b�	,�4өE�c�lb�[ހ3:AS+V� �i*��L��֝��K��Ꮫ��H)q_���򾢤4��F(퍇�O{��6�:��͡h���0Cl[���v}�`ԅ�-�;��V�>��!�i$�n��r9�"��Ƿ��B*L�\�zq;{�4y5K�<V��QLI��XF��AuШ,�SϿ��^�K�|և�-Tǂ�I�u�J�G`�9k��X3��ӗ�����mQ��n�{k��\�Tn��2�.�|/'O[^�H#>�[��v�>��5Xډ�i-Wg�����T_e�I;d.��b��M�����:]�*�G�������'��T� ��KC=��HmgV���K��"���iɼ���}����K����7�2�%M)��	�hs�0Ľ|9Nb�1p	�V#<e��=���` 迌'�֗�̓u�ՃERM����d�MW�����(�ߨ��ӮmDwk�L^	� m<�"V�x�V�ͭ��Y���!�)I�ѧ�u�PX��CL-��u�Y?��4�{�Nm��c���Q���7��$n��Pc-��=�y��T;H��-y0!ˣS}9��8�?Љ�;�&kA��=,38tP�$PvA���C�;XW�DbY�ܵ�|J�5�~-SQ%㱙J1�ڝ]#� �,���I^Am{���~��`ߠ�O�匫�k�Y��"2o�9��T����^5?���z�\�"���*kuz��1��_F�����ɽJ�
s��%\\`R��X���%��[���/o��¨����,��i��y��a/  �1���5�bͨ&Ţ��dD��G�v˫S�z���g�&�i��S3�ջl;4z�?1_���Q1�]A,�2�'����`����ᴃ2�c�2��3��Ko����V-3�	&oH�˯�S�X�^;��X����Eԑv_���}���i���@����וm2�g���-5�'ZV�tݴR5"��qO��Z�i1�3?�A�
�U]�Jmb�P�1}_o�Y����I��Ûȁ�mq	i�uo1��]	ޒ�H�Y��گZ������;^�)�����������0�����w�͞I*:G^]^�4��t�6�g�Щ\0'���)�{��WH�or6�׹;rӦM˸����4���7u��l^���Cz0�ɀ�^�&k%���7�w�iܵ{/}^�1��M��#>�`���v��Xȍ�zR�B�ܲ�*�����C{��/ek
q0虜��o��$���tE|f7��(��#q><aϼ�ϒ�?O&�l�����V�����c.-��3p���C����c�0(Pb�/�lMvX���*Pq��Sh���T$~v }�;�OP���}�)O�����.y䶟��c��|`����[���ir��1*�ƪ*?������Y��Y}�
c�bNV.�hC�p�'��zќu��N�F��J��j��^Q���G�I�0:\�M����C�%IPpW�4I^פ�ĥ4��
t�{���{F9Z��k�W�d�Vy8���S*�2+�����.��~��Ɂ��N `bOt��ͦr�wd�W�����Ah��F��t�k�(*�=f! ͜A4�H!�0�>�����*�y9�i��\$dS�Z'��!F杻7˱.e�^t)��[W�?�*�L!�ZGk.�4�@!�����d_$��o����4�.i��+�'ާ����Դ�)��@�6ʰ�K �[Y����3K�V^* �|%2	Q�+��O$����X٤��w3�i��0۽�c��D2��n�%��`���P�~`���u�@�����������A~���Y�b��#(©&���3��~����9	���Y �N����{�������澅��d���ESt�����C#�g��'��@��q�g��[k���: ]�`�?Ұ�9k�Y;����o`j�dɢĲ]���_�δc*�8(�S�m	�T���q�|�����j�GLږ�/5t��vLHXÑ.� ሔ{���N8^ݓ�sջnԹ1Y��d"�#;�K��	!��un:Q��!�"�s��NȥuSZmNN���h:W������[�&�k�Y��
]U�!��r�D❉n��[>\�u��n�t<u) ����n&P�g(Ĝr&�l�U�Z|O�7��	8�w��듈��Jv<�wR�C�-�=!��=�B0��.�y?e�R��ɫ.�N��P����Wa��73�E,����*;<�S�)�?�q����pM���5]�iq�>�ݯ�f��t�!�"ec,��!a���z�&��3�jϣ؀��ٿ�|6�=�&~��]O)e?��Z?�/���p=�@/P[�6܀�{�X(
����װ����u��#3_�.���� ���!K0��$�C3�{ߠ&���*�绝��A��6���@~�M,>
���5��hJ��Կ��l�+��_��n��̷�v�N�ι���h�gz�k��19?�sB��d��XH��0��wi�T�R{W�=j3lݫ�rQ���% �-G��Z��KO�ͫ�fG���o��֑3Z�a�8�<�����O 9{���s�ʑ��=1�Y~Qk��[�4�p���q4���e��/2����̴Wl�{�ʈf���oI�ϓ�=3v6l���S��8��'��p�=�?����7�g0�T4^���}p�K���x�GAnv�4sr�M$ʚ1���;�p�Ϙ�8gH�겸w�+�#�aO��M���ɢ VOQ f���WR�Q��fCź�ҚL�l"^��+S*�.�V���F�l��ӯU3�2� �P��%~�[|����a���ǋ<<TǱÓ0x#��$�ں�ƭ� �xl����/�=YίG��ck*u�<�א�8���]3��Fh���y�r�*��� �`H\GF		� %��}&�	GOq-�^���4<8�w�$�F�D�	/�Q���k�n����}hN+�W�����dH����~�.�+쩅�_:33�-%ff
��Ԭ�`���$ _�a������3�eV~�ғ�Сu����q�S`|��(��F�h͈Zl���j�h���K�y �?;5r�_%��e�w�<�zI,�>-�x���`g��_Op=��[Ð�1��)#��Ѐ�^ΐ*d��VY!H ��D��.F)l���\��om�[��=mj-s</}5n]�9)�B
?�V3�>�j�I�D��F"�*����W��r8T�d��j'�TpfR�P���ԟojx��ӷ�ی�Z����u�%�{�"4�0���ܴ1k�<A��S��,���~Ms�VT��X�S�*�#��'E4>��U=Ap�"7�=��ϼkk�n���|��;m��/��u���R�G3VH�_�&r�j�������qoIjé�K���i���V�� =��v�� ���Ī�t
J+*C���6�bo۠T|-��w�y�݈"�Xf9�[YIw$`�"��R�'�HA������JE��}l��Em��i%V R���Ϡ����ca��t�����>��?ǯב�_t2~1����,�/�	�MR���R�ldҡ����u#�(��3q��#K*
A���J���Z�#nE��	�㨁�@���m|��~	�+��;�K��F�WB*�� ��$0�ƪ�����������$�*v~`�m��$D)+�L*0%��T�k�R�Q|vm�O�>ÙN��W�H��ql�����ǟ�^�7*���V��[1��	F��@ʈ��x��+����ZV�HPj�ua��B��9z{j
�"rZc�	d��'��愑��#2���[�~b��q�'x��iz#��!�=\8,`���v�\�7��'��:�7qY��{�`8��>Jnþ�r
*ZF~������W�5�Ǆ�w���	 
�dV4��~Pڦ�Z9z�1�F��?q��]�=����f���m����G���Λ�FA{����������ej*�:��"X0§w���R��oU��%����R��#�MI��6cÂ���A��S�)�.ڔ�[�����,c�D���(v�GՃ5�d�♒��1܉���rjG)�xK�!i������Ō����j�;�[K��b06�G�~�Le��EN�z�9-n�U4Z��q^}�
�z�ctn��s�Z8e#Q���iϪ�i"^�LI�ǳ6r(�.G۠;��z��7S�fQ��&�/'��.���E;�z�u64���'J�$c}�yP	M?�ͳ�޵�۶���8��-����}3'˩b��S�5Y%�5��#�cb#�d���������v�}eUI��W�̨m% ?�@�Ō�}׻T�NN�9��4�"�绲衈a�/h#��ˏD���4h��5�.Q�I-F����<�!ϯn��j�a���v��4f�\�|#�gX�ȞO8R�^�B��~�p���4�	�ְS���*U�%�ʶd���Ep1Љ�=���ζ���$�d1;������t7�uq����Q8-�p���?�K��C2xy�\����^��7�;�?�<���)�0��ju��m١��$[�<g�Ƒ;ܶZ��3�B�"�.�X��Y;Y.;?�L�J(���K��ou��18���J��$�KO��_�k��QK�`�#�F�i�x�2jM��Sځ����Mb3'h~zL��v�����S݅9~Ϣ�
�H�RB5��Pf�����fz%L��Y|�^�\�Cn����bM.g7�RH-�V����$��5����Z��M���{��LH*��3$��jA�.�U�D*�P�Y`ə]pX�����f��@1<��H4ks����n�������ԶCO>����zI���"��d��?RD�0H���HK=�*$��vY#�w4���ן��Pƕ�O$��,IT^>A!����IY�UN$QY�f%�x�pИع�,�׼�_9#�+�ʉ
�q���)�i'�6�Z���b~��0��f6������ԯ�1��\�l��зmp��^S�D;�(��"r��S�_B��}��n��˘��ʌ�3���P�&�#�����F�ljI�
������1̓S����V���mֱż�vK�1�E��U'�����&{N[�T4��T��00}inx���Q^���)��Zu�V~���>����O��.�����U�Ғs�q\BS�:$^R�e�$)��x�J3 ;"�0�:�q�>��F�b½F�'�`�v�v���f��h�:q[p��iv��q.�����V��;���{�CZ���Yp�/�����H�8��<�?���JȨ�6�މO{�eCx����6�G���'�:��N���c;,Ko2��˪�?�u�V� B-��A\�_���u�Wrh'��y꣩��$| X���;��un�w_mK��E�mVW�J�j7y�!�!�#�|py-�>	�4���;���{�o���t}��YL�C�Vs��#����4rb��Sſ�9��s/$	���>lb�@},^�o�miH٦e0�RQ7^t\ٌ�a�늠�>Ǉ'H��j��Ŕ�K?�edۣq.mD���2V��
�x��Ɓd-6`P��O^�C��rP8Dz5��Y����¡s���� AL�3˖�ͨqU�P76s��c=.aO�?�Âd��)`j�즖��*l&�UW\4�*0^���� �R� ������I���}4[��R�=a)�c=�u8Y�(@��I�'��LM{	o:	È��k'�z¤�<	��(�+��`0}uI't����g�tp�O}]?^w�,��ª#n���|����4V�����..����y���O|��"j͓��m{�qj�ǻ�N�N�<Pϧ�!�
�j�h���I:��]�K��q\&GL�-�j�����&�˸Fi���k廨uv�v�Ӥ��%���h�~"�8|f�W>��Cx��������8��w��6��.䩹����@�39����&�).z�� �0�m@y��/z�_���vG� ��ѵqOU�+^�7�o�<A�!�[��^�F�S��fӰmO�����׷lд�-i�nZA�����'ξɪ��ʞ@����P�䕓Q�M*��
�;�ty�j|��/�1A������dm�n�0k�Am������X�7��M��k�ngp?�F��iE�������N�j��EԿ�/�)�Y���@���N�}������#����.2��q/!TH����K؊Ұt��/Q�dv�I,$�+X�G*F����@@�I)��D��%��J_�r<�:����+1ۿ�������C��i��aV���
wǭ���5��H�<�,�%�{�4o༿�)I���P~�Z.Z�
�����0�6qqP��т
�^ ��qs�`r9͉6@ސ�H
�;��[a�;@u��Mm�

ܲR��b�<�v5"�L��`���Gӹ��%��m�YD��s�Opnݨ�%C���ʉ6#&)%��+�YC��pY�4�od^�N]�_�|����
XoT��U�թ��4.DQA�!�MF����8F���\h><˽K�nN�qD*������^�>�3}���A�0|$%��+���|@Ŷ�-Gy<�G,��N��Ol�VK�Du�K*i!��&���]��! ���N@V���� ��'�w�J�&Ȫ��~F���"�zΉk�tE]~� �m;C��� 7�I���P�nЃ��2yG�K�K'm�(d��8ڃai�fZ����l�:�dk�x=�N�ů�/5z���9g�<_����q�l6����D��o9h?�;�Q�w�@�w�At�h(O6�?[3���~{�4x�S�o�
�#��vV�:��]�l�'���\����3�����u�U,�I&��B���K���:@�nf�Јw���	Lw��f�L��SZ�b����BF��1����\��TWT�������C������9����G�_�J�#0 `0�&y˺�S����4P����>3��!�{��\���Xqi�5[���/Οݗ�E���dj9�m�i���3@m>�U*�C���ϩ�f_��ß�)W�<�򙋵 ����a��SAP�f2��}���ZNB#7������d���G���ߑ�c���=����.ꁜB���Қ�J�
�bC�5�8���#a�������M���~�%�5��!YK>�� ���fe�1�����UJ.iKC�Lh0��|���]�����Y���N;�� р�M��ig@I��;^�X�Y��!���o
�j������@��4���Қ]�V0������W�����'�H_�O�p�aY)��n��]=`7�h����(X�Wb�2W(l���F�׸��0�7�qOz_%�,�1i�w+`���(ٍ\R�rQ�W(x+�|�͑���Bd���Ġ��Mb���-�
�T�U�O��YǠ#u1��e-c\�m��1D2�-��������>���Q�Ɩk2״ۧ���r�cHQA,Os��&^};���yɄLUG�>pU>�,Z�)u���v���(�w8x!�G�r�0��vC:XI��B"�cQGuX�:��m��������Ӭ�V���3Ig�'A�  .K/w�s�p��ҫ=|��u�E���h�D��N}�<U��R0ʕ
iD�f�J~؜�j�����H��!�(`Ztݣ��	�☇O��b��~ƚ�@�������.	�_o|��WX�˿{���v��ym�ެ"M|!kqK��dmB0��HO����e�I� �v�yJo��́r�&M�%,;����e��º_'��7עϾ|��P(M�\1<����#hޡA��y�'�p9�|����L���S}��e���Ѹ��4�c���ԕ��`ߺ[
�*�i|�U,���s�
z����X�߀�2Pը�y��UB	���!������MQֱ�>)T�p�@4�,Q��vt��I��!,,}V�R��2�����7ĺkm�:1��5�6�<���i%G�:�R��j4>�QM��U�4��ᅺ]�]ѓjvj��$�'q��Qc��0�I,\;�sǙ�ȣ��!ߺ�w� Q
nL�!�f�w�ϗ�+E6_��5�[�]����m9�56U'CϜ�+�c��l�(.���O;H�{)�6.���R�,*Xv@i;��{��~Xcj���@bg�����2��o��Ki�����H��Q�S:���\��n����Ed�ֆ6AXp�*����]-	�,�F�VՎ\�Q�z- r^
k��W�e1�j�E~d?o��Ä!OӐ���+T/�G���q)�	�GSdF���wu�Up�Ԙ�{�eQҜ;��>��B+�rσ��zT�I�(���%�yh7Pq�$������a�Z�-��~����/�h������̂�˙�=��� [d��J��?LzwCl�(1��29��O��f����5����+f�h�5礇	�q��Sw���@������#�vk(�fM(;\}�K*�8(� �(A�$�Ũz�+�	����פ��д\�(r�i&�&O~�~�ZYf�5H����55< �l�E�)���h+A�/��&gP�S�Om���.�s�y?:&f�}�F���ɴ��;Ov1��4��	�%D�������h�U���&v�g�ˁ���K!��P���� ? ���R�V�Њ�*}[;�gqn��~�v�q*�_P��G����mP@���	���7/�$r�*��\���:i%Z��?[�Q��y�:Ύ"��Q`HQ]����7>���ki��0~禔V��҈���I'2���h �F�W���k�����!y&J��D\���x�i{c����ң4���T��
�	��ۏF�Q�W#���a�H�X������Y��f��G����AC�L��U4��(#Wo�ޗ �c�Cx��y�D}`O��l%u�Z�=V��9�,񭓲The�2��M�j�:T�t׻����������(�������b)N��;���v��z�����w��y���4��l���AQI��-�������9[�[6���7���e�#	�b7Ƨ�����T���+tny����6�v�P��{�[��J���L�;�^�#G���������!��2vA�ǗL��[���p��;�~¦�`�2{I�ZɐCe�(k����a����0��z��U׾�>@7�H����:Z�I��6廱�"鎒����T�ܹ�B���z��
����;E[V�:oK���u�F��Pca�n$_�0ʣ׼�z�o,���a�f�6���c�j�)���/RNB���iU_�z����`��^x޷� �M����6\�!8�ph�ճ�1�6-[u�>l�����IMI[���iMfr���Nm)>Hn�ƨ
��y��p"' ��__a��R�����ec\3�l7V�P�81d��/C�������a�Jb2�+��q^/�$˪y��gF��U�g���x�E�o���s��3pE6����p,Pk4E����A�R�2{��N6C�������ytz�;�������H���:^���@}s�\bP��ȸղp�%3Ps��j�/d��H}`��Ǵ�VdX��>��m��b`5I7��9.wwI�Gs�	guZ}.�+�j8�
��73;����.����3��T	])�֩��Oz8{��1�w��U�&{u���X���h��9؛�����)�8����k�Q��m��i̷ό����G�O�}TѴB�cb`����*Y�bHy�N0E����;������iS�)�_Uy�O2m�#*C�2pq#���ޖ��院��#��fW±~�r�rع�{���~	-�ࠃ'j����u�X������Q�2�`� ����@�@c���ph��=O���_�J��N	7&=�������~���JV�/=c�-��{��"����n���P�k��5KB�ԙ'�;R�"�%C@��1��I��}Cl7PS2�%R���ȸ��'vӈ��x������܈��j0�����k��Ӆb���LjS3��e4��։��*��d{J��@STO*;��(9��GI(�?ֿ�����z��D���5h).YVfl s�l�X9���R[��`V�޼�qz���2BaߪA|�_�,4�NҤ;,1�����%�w�a���W�s*�B��)I�۸�[9Ił-B9u#�'m��tǚ�Pبr�3������)L}}�#{�.&V�jy�����2���r�6y�)m����1.Q�%��^U�y�Pq�0��mwR�E��}�M!1�K����]���g*O���6F���G�������G���,�@F�O����J�xm��6ke�r -������v	�Z�B�������w�k'u�`U�Ӻ�	ɪ�A��t�D���(=�<GO:D9��x�j��ן������{�xb5��s'#�� N�RaM��?�C��M`��TQ��CϘ��C����if6�rs�����I�,��ÿ`��Qb�Y�dE�菫��
�(Ja��ġa����|��l_.(E�L���t��:@҃6���Ţ_��&�`�A��f�����Q�!!��ē��@*�i��=�8.���Y�9��xw�'Hp{��,5�U��k["�����,�����M�.|"����q��>�F��f��Lꀢ�剀��5h�.G4��s���9��L%�i'�m�hoKH]Yؼ
�DV
�1��m(�Rv%��xU�:��x>l�z��O�����d�;�w�M�A�ҙ���R�Bl�`�����%Wj9Dڀ���
/�s@U��s�|��C�`�HӃq��5���8#��zo^�E�FW���$� O���B�b�׊w��fw��z=1�#������T X��_[���}ۛ�`g��yT|���z�88�0�v�6d8u�+>5j��Ư��i�8#T�)S��%dז6Y3t\iF�h����="�a��q�/�P�2'
qZ(�vp �/r��x���*�pj(�!Wz��5���<U���lf� m�4���u�6R��Cz���VɁ��{�������˞J}�UVdv]n&��"dW �W��jT���Ԁ��1��\��p���'QNk� ~���P����@�ln�1�
�-^�B)����{K�{GM�U�J�RQ�U� �7[���*9�q�����I��<�<7= ��$sb
_�o�wV,^xԤ�gl�pM,fn?`v��m���QL�� tD�v-Sb6X@3�S���y��%1����ʆu��Q�"'�D6��{���]7-��)؀�"U��b��9�!K�jS���A *������@k��?T(3>��RP���D׉����70}W�ACe�r�d#"JLz���9��Ux��o4k�W���&��5�RW辏,��Q�IM(����f�֩������#��D�u�麎n6z����	�b��>�݇�J��K���R_�g�%l?�������2`�0X��L�H�9,m�������i!)lL�g�1�Ō�E��;��,B���_�j8�CG�84`}8�^��6�{o������5��o��c�}�
9b]�-�:x��t�X�/p	i��U"h����;�$N���m��s��X�!־���V�>
��Q����"W:(�5�&C�םF���@&���t�
Y�J�w��ە��t����Ǔn*��F/�w�����?2&8h��i��h�(��]�?{��+oi��#�s�#Q����x�L3B�7�sU7�ԙ��Wg�!-����44�#�q��e�) ��X�g���H낱r��m�Ub�\u�N^JY�jrq��r݃#��tӿ:��J�)���>�!I��vs�Y*Z��7`��B@���>~>ɵ;�g\pJ +R�S��W��G�|xA�8��9��L���3��O5T��[t�1�`��b]���zk�.�rt� V���le�[�0.� ��Yrͼ����mo*�N2`�#WÇ�o�����B��H*���H���ZM�5��#�B�4s7Cs��E�dz�!���(���գ�x6ψe��~ˈ����>"�8\���y�y��{�aCo��Rx�%�d9Jw�	�꘺�&]"X!�q	-,J���>����K�n�Q�)��i��#��>,�S����tRȀ��ۢ����5�$=���]i���5]x��A�]g�ȝ�����F	��Qw +(� P��˕F�j]��V)O��P5�����AR��m���X��SĖ�dc�"�0Ѱ�fd�w��ܰߒ�C�T\d�:Q��n��31"�D�������[�.>og�0Ou�W����h�Y��7He�����q˅���f�o ��D��k�����Uя�����,��HO$���G=����iq����̑��8?׬�!�.؍Y0ܙ�!�"����6mB��;�U��ЫEYM(@�qy�]]��dX Tj�(ן��	Q�8s��|6�k'[�!�
�,�-$�\c�X#��Ŝ�rD7�qx��up�\��`�p�zXNS!�vĻU-��D�G��^Z.lΡe�v����*�݆	�H(�M\�A"�k�.@7�<�QG��h�N�׬^&���*�DK� I����1����t�kn�⢿�9mt:x�`���;�x����6��	�/`j+-TS�Qˍ��E���cԾ�X3���=;-5.�4E�,�[�GI�&��9+��E+�M�J������ڤ4b]=m
�8�����]��A�ǰ%Z��m��\�����mJ��|��t|�~a��ד�D �j�)� ��>��w��C��\.��"h=6`R�~_��� O)��_{l>��»1�O#�>�%��8�V�+3���y�f�Q��eU�� 8������C�q��d� ���^�
Z[�܌����*V��5�|!!�<&�����5?��.���<�}~���� oX�:��Mo?�q	3�ȚH��"N/�$�e_����q!S,�;�SH��eȋ�{cA@/%���e*j����r��
���\�:k��W����7��5eF��6,�'�X��t��W�pݧ���oQ�5�-Oʏ.!&J�����PX��8mfnu�_�	�Ǌ+r�����[VQ��Ӊ�7�)P^�4�Z���tU�t�OD�r�`��Y��86�P�^�`I�1��1=�����<,����G&6+m�Y� ³Q�C����$��3�20��r$�?ޤ���������K�R��C��	wj�v���A,+�L� yEJ2h-��B��	�-���@K�X��h6 �=4��YU�P.���74�3V��=�K霘������++{�C�[��gt-�=F"��gW���҈-����J=��ɍ���W���)P1���2�Xա��l�����m���1�N�a�ތ���^�](h[�!V��7c�_��P�a|-�H����5n������;�T�$��oa�zp+Z���S�C^%w�����V���C>�7�:���������G&��[�[����Y�Q��&-s��U������+y���|���t=�e��a���߶Ul������~Ui\J�ÝE�.�e�R.C}`���,��g�M�{�B���H���NB�Q�!ƌ�PD��ԝp4_w���05�8td�����u9���`�Ҭ����h"c��,��*������X���07o���>>�	�r�)�2�Hg/q�5QD�o�D�w�׽����(<@_F��򑩳s��zZ�S�	7v�)��s�b�o��@*̥L.��j��%�Z�P@\����6ANLt��g�	@;�2���j�c5W�R_l�����R�x��}2���ܔs	|e�7[;��/y�1W\��9�(��O�<�-c�,�5ų#E�hpRW�u'5�����?��Kb��'�y"L�����}
�9��.R�-���:�g0C��=C5I�n��������L�-0(q*��T ���h�;�l��=.���o�nɟ�6o7u���'O����̙e�,�T�(g�\�b�7�HU���*}ʆB�A����ӭHa�U�ދ��M���v.S�O�7Hݱ�+��js|,)I)򳖼�O8)8�Tl,�V�);��R�^�a�Q�W�(0U~���d��ޛ�)�3�p�їZ���z*�cٟ�:�Ӎ�c�#X��e�5�f�r�K;f����U��Q����z�i^o��E��$��/Ȁ��V'�r&*��ԣ�E�Jg�+���E]hQ`]�.��r���s��5ߑG�h����҅$I��j��]�1kuĺ��+�8�Ȕ^v-����
P�4%��c����%9����� f�v��J��{�򶒤���V!�T�j����p	�d�#�|tV�o���$��AU�!����)�_���v.c����Fs�ɇ�Gܬ�b��?h�$�3<�^�5 6]�r�[`VC�|��g*�i�uhpvks�7�r�*���A#Y_F�Tz-�C3�y�a��! �P��H�g�;���f����3T@�"AAfE����Z3�PA��^E�EQ�q7���Os�? }@��N&�邴ە�����6A.x���u� �U��AʉI���z���2���0��^�eH�%[��z�2792�f�=��~ɠ�	v��SG���
#c�# ��Ƒ�C�]��C��ݫ޶t\�G������Wp�`L����wѷ-$���oǿDD:A��9�N��<�sd�L��/X���G��ҥ��q�݋�r V�"j9��� XF�4`����zÍ}���Pq&9���Ol/�����b�Cq	�	 �G �{�G�D��K�@m���#+ved�xY��}�:}a���G�������O�yzW��qS�]�^p�㱳���X����>Rv�������k=Җ�{�W�G��z�z��ƻdP��5��.�d�,����^���n.���-�'��u��t6i�徧K������Ӵ�o}��F�y{�#T��0�����q��̍Z��<"���|� �P��ʥ���ϡ����z8S���`����	���8:]�G>��);�t׶�'�������~Ǘ������!����1����bL�hX�O�P���w��Y �<���d�cV_$o}��u�-�:��]�Z[_�� q�U���M�WV�
���%x_6�5�I�VP��ۚ�Q��ky<��Y�&���n�ݫ�_8�a:�����paB	*�L��iEw�αc�4�Oaub��|I8:�˾�9z�ူ9'�{�H�zM��GR�?X���+>I�`��F�r?Lh49��a�?)7��,~S�r&ꗳ�}�6����Zya��1�z�\�9�K�ҎM\�c����c�J"���<v����%�>����^\��:�rZ⚁v�3r��s���(ř>F�h~_.A_��S!�mv�����3�>l�U6�t�#���\�$>��ב
�T�kRoU�����l�ٺ��n����o$PKq��1�T=<�t��1��{��t�I[.!�A��/�� �ڃ�v��r6�z�3�nƮA�U=�H��n�r��ܐ6�2�4B�ad&�׃�F�(���v���1�\��2$B��#�*�\�l,k>ے��� 1��zȅ���i1�����[��k�i��2Ծ|"����ũR��8��V��b����h���|�_>F���� /�%`�%QjC�'(���n���'�T�ܝ�t�q���n���2L��������LHeV�8�����`
��m�	�(�Y�_��'�'}�w����ԯ=0 �:zq�wp�����1�^7Qʇe^{�P���m}�E��iU$��0�d�2hQ�%�}n�� �M╮uÓ&v�u�,cN��zV�lE0n
U-{+�����c��|��»�zɞ���Q��R��vN���֠$,��r �K��k��������
\�	�3`B�o}�"m���;2�&��z$K��o�7�V5s�B�����yߐS�`ؒ�u�L]�eq�5�sL䙯�[s%}J����� F+@�;��%a�Ǒ�����G��r$?�/�����fɽ�׳D���*�U�M̌�Wj�ͦ�]T�����b����A�1��R-I;N�|��A��?S�N.����B�X.�C���y�50C �}܎�D&(�áԒ�'��S��4�Z/(LA�'E����\h�Z�����P��|e��|����WDif�@�G����{LVy���s���V�@IZ�SQB�o3$�V�)�5��uJ����'P4���t<�%T�ئ�>���h��4���8�5�Ծ-{*���OOa�9~�	�ܦ�C��\kGk���K{-6U ��T���L�
������b��D׼sx��Mw5�}���w�%��}�܋��㳇_P�~���4p��\t1Ő�6�P]�|��� ����L"|_�����*];��K�~n����F����v6 Ũ�%����ȗ��r��Dy\)&΁dL8y_�6:cYn�x[(Q�0�e�xj���.��Fй`��l����^o�M���ܢ���Ǘm�T���c�y<47]������˼0�F_���ވ��#&E]f�im� �X�/�z^Gt߆�S�������g�f�K��i|zU����t��)7j��|�1\��d�
�#��J���А��5��.���foI� ��C�,�T�׸-�U����<�D}�u��;�s��)���c2U-7���x�51> ߧ�ٟ�Qo$�[ƀ�.��>�93�D*7(�j�	x/���2�}�b8uUi��C	�X��48��=,`�ɞF���s���[���Jz�(��19"��|sL��ޟT��S�����ZM�hp�f@��+촡Q\o���Њn�|�Xr&���P+a��ffZ[�SK� G�]w[�:�mHg��B�Հ���m�=0�ù��s)|@^��%�5�[�`w�_�����T<
f�n����㽋py��I=��0k�����ܼ�.�ŗD'��,�X F{l���9�}�̿q0��Q5�8V���ߢg^��K�?�؈ga��g ���3~i�G�b�nv�n��O>kڳ�a_H��C��t>�Csm�0��;���6�����{�6�z��v+9���Q*֥3����*e9㒡��`������D�e���'4w���-c�`������y؂����O!ogǸ�,��IK-��A,P9� X�{%�x}�@�&�u�$w|�Sӡ[���O��b.�>WN��[�mD.��L��H��
��˺Ҽ�P�մ��ŕBR;ɺ1��3-h�����Ϙb�F�T B��N�m�t����ѐԷ[�ݧ���2��]�<�2�0��h��&t�U�|��7N� ]�����a�Ɔ����~��r��j����@˞=�ec��w"i@�K{v�����'c@9�W����AU�pSĺ�ޜi�v��3�e�I���Qq��.IjXj7��������P���d��C��t�����+��.w���{�۔¶�W��'��xӬ[+�M:��J#j5�Il�0<6��/�:y�v��X�f\'���|ra�pH��Ԟp��Ư �=^���3(�3ܽm耫�Pa���8���]����P&�km��۞��m��1T�bV7Y����A{/��:$ G���؉���!e4'�����{�8"��k|�/g�+i�j!�#y��1�%��&T�Ґ�sAA.fE*��}o�d�z�M(����g�]�D�ݺ0x�	|
-A$ɦ�<߫�P�c�j�hN���ڄ�fpD4���6�YL�E����,ٕ3�W�,�K��a,�?��U��gH)7��#l���;�Q����Y���pn �6���5�uwZQ�,�2�mӗM�5ɗ[n��QP�d�؟�g��X����i��6��l�n9�6�>Pn�����A�:[Nf��Q� W��Er����w���"p+�_�9���d������,��#J:B*��,/���G�����x�(N_�gF~ߙފ�
�0%����w�xߞ���/��kͯ���F���Zʺ3]���:�B�����N��$����	6V���=T�cw-��8�ޞ
�Ŗ��4���u��6BSp��7�?�eנ�FlG�;�{��1�U�^
�'B[���f��ak�Mw��*�H�Z�\�0��{+�qt�B���4΍X�0�R��&�ⶠҦK]����(���g�C�W���]�BK��x� �j��|t�(�/ͥB�״���1��0P�ok;�L#HZ�Z��X�S�p!�U�%n�9\z�ep5���љ�k*.�e\�.I��;��tD�,�j�j�#������k� yS$J�0�]q�/F9H�Q�CU-�#)���������L
:��_	�f�=��̪����R��d�ų���������)�O�� ��mٹ�Dz�B�������ƺ�+�=�]>'&5��'35��2a(6*�{N�-z�:�u	3���[ѫ���k�`�����;�*0���y4���C�����jIr+��a	����.���6~���aZ��o��k����� �$�P��w����,7	i���T�t�8�Lo�4�Ay*�B���%ٍ�$��&+;��ť��*����(����+%XW�l�
�<�h�c8�ɽ�dF�-
��R3;;Kn�v�\���q 4�>������@�rq�cT���psX��s���.��5座��O_���c�z�F����bV���e8��Q�7��{158?_T��I�v��d�Q��=*&�e� $h�[�������R�U�9Wu�<���L{?��'/c���r;�b����� q��X6NɶՍ���1�)���:�*	۹�'��A��Zx^q7H��������axP&<��ۈ�3,���r�ۥX�E��o��N�d
���>D��Q�A��6(�d^�3#E��S&�������b�w>�_Q��k�1?�ʀI*5�<�La�k��G�(���z������H'��vʟ�e�$w�c�,QJ8�$�ݭ\8����%DT���CȽ�wpO40�������
��>��W�o���e꼞�r��-�D����n�]�[bf�I�in"����$ךрY��~<"`��ʦ�CN�x�,[o���)C��ȶ}�ʰ���}"�?�U�l*�G\)���V)?A+@f���0*��{hͦ׿AϿYz�*�7���GK��� �������Cp��cG����1`^����PW
_��Ͳ�(�˙F���C���(ք`n���Ř�ҿ�uS�f^��Kt���u�u��uv��j���t���B�ʒV�l�7%�0G3�]v�X��)e�q��~��d\��7J��?�!����΀�tz�jA2s��s7D��̞/�AcBD����:�S�Lh�2�u����2�6 �� u%��nY'����7f���W��~x ���L�Q���1� -�{�C7i���>�Nc�]\�����^zK3�Fpm�xFE��s�_��>ۻ;���ƙF矙x���P�\��;A�]��o+zmN�l�;3�f�6�gf��5����L�BT~�{7PH�,�<<�P<��ܪ1�҉��]#0�K���&n;�2�Ţ6j��T!9��O�7,��J�"YiO�i��e<S��^�������Y��"F�QN,<zѳ�S�����X_{�Uq�M�wc��.O�����1\}纳���EY�A�h���ǰ-�5�Oc.59J��ƍ�mx6?s�4gj�*\r�����?W�^�f����aT�ͽ�\iA���;��
�0^g"��;&�'�b���E��?��B������:"o��˻G��ߔ�������DH9g�,
��F:��d1���,yj�*�P��[ie�-�^�R���xwh/Y��°Cơ1��fそ�(�nB1�����&�G�ŧ�J-paB�a�\^��k���[x��5��k����:��E��i�׸trN�s���hb��\�EB�e�٤�ۆ� ����Zʐ:52�pFG?;� >���q`���螿(�qH������\�	4}_E��5��~������j��jFo�ky�Dz��鄪o���E�
�5+̣�9�yآ&�V���+�w�lR��^���-~E�%p�x#�e��븬�!b&ܙ��E鰹� ���c�������ӧ���ǿԢ�����T�Y��{U�y�;JpC7X��ˢ�
yƉ�9BiY\֫�6 N��I�v��j�'E�1	��y�=X�����u�J�A��H�>k��T�y7S������+c�O��G]�r�X����؈d���o���Kߌ��m_��H=��򫒙�)�i�
�Ȑd�6p��k��i7�>�?_M!��&z9�b�|�Y����$n�����Ex	9� ��j-%qHX�+�L��&�= �/T�_��C�����m.w�č�2+ܨ��4��!���T�P�X/`�b_��9~M<�
O��Ox:-�{Q���l�� ���[�%�+�`\��/ӧB��&�*|�%�`c����S��*M�-1Z%1�a���M��K�mbl!*6�/���"yI� T	�#�t�N[о��g��Q��-��MlzY0����p훳$�B	�x�U:1TZ~�sxq��XDYↆ�g���{	��� x=<��0Quu@��� R�3�JU��P�oܱ5�Z��ı��h\����:Ŋ�dt�@���pI^9�����O	�����r���~V�]�;�`&u ���$���
W�TD�������T=�IG�rH�qnk�p4���QD�(��ކ�G��>˗��M��y����|��xk�L"˸�`�����g�u��$�嚉5�BW�&W���<�\�\J��E5��2逭N6 N�^R��o&P���_CL�9"��1¡��ļ4�W�if�z��׏�7����4�
��}yW�|���m`ei�(�E�F�h<6���LᾹ��C������o��z���풃��l6���	��|t8v_�	N��Mώf�r��wx�/1�/�����S�o.�8�׍�Ɇ4N�����v�y���~�ԿNӕ�K"��P2�Y2�Gmٶ}۽Є���ے��HsQ��`��_Տ9�+�����6�f��V%%q��n��0��9:��,��*��!^�/H-A�Q�<��vS4���PvNd4.��X�<h�7�����x*�d6�������ǍWCj�C0M��9pd�?D2T;��"er��#�c1�rPg/��Z_�Rh�Є���� Z7������(�߰�p�
-r/���l�9`�o "��)�-����<�WA����E�3Jۏ��J�&<��tڑ�ѣ�(�J� 7��Z2�_D������&U�_�̜�t�d��v��:g��/�^��A�=K��	� X��VI��R�hf��T��R���������&Φ���W��&�0a�P�F�
�1+�;s����aG\X��}mO|ҿ��!���'��?���c��)����,Z�����q
{��O8
���2|���mJ���%�T6,�7��ӕ��Z)�G �%�\��g��Ȩ@�4��k9�k�>Q�O(uO\����pCq�a��E�{wE1}�Jz�MDNviʡ9�Iߘ�MFT��d-VB�G��Y}GX;�5��l�����I{��֐�{*��1O"� t�s�>�毹w>x��|~��t>p~Z�ة�[dգR��{/)�8��M����uұ�jR���\@������:�_k�\��y�,��:e��J�?ؘ�E&��ʞ��]%c[���zO�d�~�����⊌�5-�ެ[1h�u����7���[�,�f2h����!�3ԋۻZ�CW�g�r�4��|8�~��	�7����%���ny�?->�P�,_�	i�RC�2@^G`+T�
cճ��M'��a��V���pf���/�O���[�M��ރHH�������sKC� ~��>_z:�i7d{e�7)Rcwq�PJ��>t�Z"�I�[���Xb�V�G,U���Tk��Pņ|��_,aͦ�}>A~��,P����d�dO�
��^����-��T���ڵh`�H�ͫ�=BbLe�v?�a�-wk+cA\�����p晨{�63��oBb�����}�_��E���$�l=I����^����ծ��S�l�r��.�
�ۭ) �@g\Fk�����9�&ԡ��y�S�oG!�I �q�0遲\ F��2V�U.�̩h��r�7]�P[��D����B�q��2����h�+ſO�����`ј�2.к���)q�h�Ӳ�~=7_�*�Ō+��ՠ�P���{���[V�ب��kw3�+�}�S��d���L �3� �^�����K��ڗ!"Tv��^����{׬����w����"3�թ+����r����G�+�6��r`��Yc���*~��C��2��L!x"!�w.�\G���Yشu��n�FL��;A��){�->��.{��������w� ���	P���D�� 5�˳c�bm�]�>]0�'>����B���*4���G��j�b4�kϤ��`>	�U �Y񛭈�ew�ࢾ�T1�GQ#�k}�[
{N������ X�>>�rKMz�v��JBFoH�ٺ� ��ܻ8y��#{s���+GM��艽1bR�)Y�a��#��_ȿ)5)O��T@�H5C���*�PuC}E�,��L�g�a��[�.n�+ԆX�d�M���L˟.�K7�D��	���o\��6y�z8c��ZCpf�O����z��BG+�լ�Lt�����3���с�FsA�����_^��%ZD��T7���3�BO&@퀙,S�����{�P�dp��z���,�ju�����.L	V�Nt+��Ă�9�i2�����dZA�%ϱ�s�.���8�^k���*���hR��p����ɑ]�Ĳ����̮(������j��l�z��[�Z	P(��Syu<1!Ek��W`j��_@aԱ��^���z0; c<�oe���tz@A�$�{�+K(��#���er�vb�W�8%�D������p�M��wՋ�{f�6OǟM�i~Im"��#��6�A�~�n+�D*��#��e�:b��5:��?˗�)N����Q���ʹ1�D8�\�U3w��T�?(?R��������_�E��d��Ƣ��>-� u86f���(�dc-����!u��mG��h��2���? �+��?���P�e��|L0�����T�>�^WӽPpC��7Q���T�5H�󡰁��^cF���g�9�9�	�Ơ���߼I��U�O����,	�%���1�j�����Z�����1��V
x�V��
�%Xd<���r��=�yYa�:�/��u9�ţ
a���X���"�|�D�Q�Q:[j��q�UdD@:�R�`4���_��7~v䔌/�[.[���d������|"-��u����D�!9�i)N��A�ݽ����k?���:��2�tVo�VkN��S:0Ԡw8����:�f	�5�����"@��Q8Qz���<������OL���}�������+����O�۲>��|��'R�3}J�j��Ry��ik�fKSȪ�n��)���=/R�oO�:�/pm4c&`�x)����T��^Ro���ōy��\+M#�k���^�Zk�!G�LI��9:�=�����ƈx�T���(H�8.?E���
�!6kjbas?6�]�a��P͢Y�"���W��Yx��؏&M���!+���5!�����Sx1�BQ�c>�|2#�������},8�Hj���F�<����9�x��d�)��6i�_��?���~7v�ұq^��W
Mכ;��q��h38&Y�yǩ)6��gK��b�UIj�YF�y�h�Φ�9ދ�J��<�v���C1m�t(JCZK������浚�bɷɛ8�}���2�'<��7DN�.S��4*�s5��m8 S��J�~�k��ކ����ۃ�[���'cv�k-�5��v�����L�' E�q�1�L�|~"���יL�-9!��3��٦,w�
�'y����j�Q�ڀ���I7�����x��L�f����Dl����zY0Q��hؖ�B��S_�!�����u:���=u����A˓]M�1:<#�����T܅��~��I�^X%���K�}B�kĻ	��k���d4�1����"df�/���ؗ�,d�_W�d�&)�?���x��!���슶Q�/��	v��T�����k�܃���.A�H�tmk�('���6
^)p][/��r��9%IMWU6��u%�D��N�w�J#�G�O>s	�h@����#�w��}M��kT��&۝�N!v�J�����L�)��Fc{#nl|$e	�Zq��M���zo�Z n��2rd��G���D{;�����:�*2vG��b�Fu��/t��kyQA�uY�'h�����K/���s���3&`��(�Y0lq�
��-OJ���v�6��Jқb`��gE�.��{���vuq�G1��7P���Z�Np����"���K�4�l��cVN��E!�t������}v�T#5:�ikɹ�����*���8�k���0~�/�П�4&m�
�c�Lq���[�����N����TC^~�����ut֕yR<|�AMI�&���+�/�H%������c��fO�֓�j�+�-0�����Ɣ̣b;𴺎^�m��J����x%�pF�����>�%�m�~o����	]��b<猪��ip��3&���ۻ7Au�)	6�{`r7����N@���5~[��QK^1"�9��_�hBg5�z�̹�D�q��<W̟�U���i��^` �3�K�R�����>G�h��i&�c�VF���&+t�������.��Y0�;��tO���CL����i�Z�@6Q�3zKP)k:���^���@����P:r��$	:Ҩ'-�X^�T�M2im�a�Q�*�+�He���ToVnk���G`=@�EV����t6��D����{�b#�%d�)�S/?���)��%kgi�p��{~U�����%�(���+��9�;Z�^ ���)U�8:,���0� ��/zѶ�d��L��?�;cUm������3���TRN�xa-�^�>�aLj,J��~�b��{p\��Q������l	=��N�z~&R����̛7�4w��e�ag�/�
~sn�@�?3=�o�9��,M����%�����Ӥ�#Ȏ�}�����X�i���ł]�/[����LU�����
�׆��m�u�0��lV�%k������G�a�6$�I�wI���0����d�2��8'���`۳�V�ܣ�s*E50n��b桪mx�Kp�H5�6ƭr@��E�$\�%�@J��D(y�|ոM�W��]���0l�%�r���E�ō�+h�c��u\��J�pHX�o����@\� �dߡ�D�D��~^NBt�\<JW-�.����b�:��G^�(hk����u���~f�$�<�0E���X�����ī>JM�2��:���4PZ!S������i��\��V&rr8s�K�K�,��=fq_�����#��<@0������׋�P}�yA�O��~['�����t����\�6�Y �pKTbfc�G�5�-�Z�7gc���ʯД����	�-ig���޶��0W\p�D���S^�њ�|WMX1�=���Wեq�!I�z�A���mk�Ft^$8�g��eY���%�YTo�(���oۂ���,J�k)��O��5i٧�zh�W� am���^�q=i��BE7�~eXc���l��-�/���b��ר�1��~H�ў�@����,¹��y�~)����)��q���)l���V(�"
��LV��V�zjbA?��s7#��6N�k���t�w=g��j��?��yuæu7��ލd�ߌ�"9G�rƬ�Օe�o}�X�eC��ժ�5Q��O���"�e���+G�t�?��W*ߗ^�r�V�E��֋&[��-=�y^I����<t}\	C���H%��ؑsM����'d3�W�������J�o��|ae�О��1�.���R�\��Y���nQR�j���T��0<'n��Xg���[6c��-�JKxܙ�U7>(HA�OB���8XFX3�W��sUY��_aD�%�,��R��%��J��c��Q����D�4�}��d�ts���-�Q�	)��vб �׼�?{��R@�}�\-2�r$��̀x�ӄ	��6��"�4>�u�Cޓ5sC������G�i���1"K$�1<��S4(�W�On�b�ƜWkI��L$��p��c�͢�Y��Z�O~�.=vB�\���7Nҷ7�"���<�P��N��{Q�[z��6��i�����p��ZW�����,�GM4�<C��ԑ�7�0B㨾"V�2��;'_o��� U�O�.�F�u���f۟���B���2tS]33�@ ��)e�)�yK��ru6��f�|��w��ޓ/|hX`"�seq��N�#�i����8�m�/��2@�y�w�w�
hƊ�k�!J��i��90��+��FP�����9�fS8j��u�:�2/��2Ծ��,N�~e�ǈ�����*V؋Er��iMa��Z�R�m�]޹,�X[xW����M�e��Y����1���Б(���B~��3W�ǜ�ة|��&�:!�Bq�Zw$KG᯳]�+�S��
��!lPe�0h��k���AXo\���n�L�������R@�s�s7���?��x:|�Fu�.��q�� �Nًuk"f�<Hx����̸,�L�zs���BQw�[b(�j�[�r�G�40/Si�ߔ�2s�2 ^�T(����u�%�tn��~pdK�<JI.u�1����/H>N!Y�i��o�͐2��6jup�
:��v'�(d��Ԇ�ؔ��s�?G�S~.�+`-��Ty
)��Ǜ��о|�^�O׀l^#wc��C�ቈ�bӉ����7�p�5�l7G�ƦXb�5���U$�}�*I"W�$*�s�֡#�gL�q?}���/O,c�^iN�G�j5���|é� e5Tv頂r�g�ѯ�d���8S�%~�E	Zz0s�J�gܖ���*�v8���Nuh�y)jİ�9&x	���	E�pcW1'wm��'� da����"t�N��8��Z�"F�\������g�5q$R%W-pY�2PnH	���[��B�����u�i#"de�P/L�\_Ӄ��"��I���0]�_:�A���-�pY`�Qz�⁙0�������A)�5T�k�ex��t))W�+K��_O����i:�`׭���B��2ȭ/a���g9ZO�X�+�ȼS��Ha��!Plde�}���F���1zM/��(� q�M���ZC�9�|;�� ��%��QQNj�xx��f�2�Y[��y���>�cʁ��|��s�Ź����^$�e�����
D+j�?�Td�[�4��:թ�����&�b�`���"PU۵A�t��Wy�K���d��ޏy�h�?��� �ʋ�]zr�h�=���Pv!l�o:�C�A��i���E���?<[g���ZYI�Q"�V��I�pp',^J�ͳ�j���J���R��M�rr@�#�! z"�.�P��Y�C(���'>��zz�m���8�*Dt
z�-a���6Z_���!z՛��/x@���E�q*�o�3:9S �䥿y�����	�F6�jU�|>+O�ʧ�����'%K�V��@j槶Y��ňa��\}���G�~=a!�TmH�������9!�� 6�tAASWْ��ԅ�4�8�ū	��"��N�>�"��v@����;��}�&�ȥ������i1�;��Im��1�4Mͣ�C�^�F��,結o0]	��(��L�{*�a�8�bj�93Xkc�%��1RŅ�=�{����4����?�!Ck��2u2�Tsz��4��jQ�H�R-:�7���X|�^;b]f9���y*@��KF���
���D��`�_[�|?�$|3����b�n�ED��ӓ�N�c뵟���n�26�U����b�-��L@zN��8�'�F.b���t*	7oǵ����:R)\-Sʗ�)�ˈs.�T6�G�-+�Trș4��re����9E���x(^3�� d�~���㲑���!Ƃ8�e��x!�֨ܤˍ~&=��t�\ix�}9;&�'�Xx��j�ܳ{Z�m!�l�0y�4�A��eT
��S_'�.��Y����]N�mB)�P:S�� ap�$i����j�"y�!P3���n���2���@eW#�6�@d�彎sNa�eSx��t+x�G���K��Y��Hޮ���ҧ�b��A��D���چ�y%=�GcWP�]�l��N����&�&[Fc��.��ޛk�]C����ɦri����jϖo�Q�5� �LL�dn@׈�gm:�k+vG�S�.�Т�0�("ޜhN�d>f7dKl��|�XDtw�'�O�1��7E��*�9��'4W�	��`�&,����Z�s �#ͺ���7.l�y6< :����-�mU6���g���H~���n���0$�j�;G��q��v#,kȽ�+�C�wq�8�4�8��Ì�^"p�,F�y1���F9Mh��_R���`x	�cvb�}W<J2�o����Xk��D�'j��63a~F��g4��� ��$ 2�OkK~�`��y�l"��
Q�$�*�O7.z>���a��^*v�0����e1EաD<_�	��D�r�C��N"��d[�.V�ߥ�M7�k`�|&��ג >6���-E>�Sa�x��UN�o?�hUn'EPv�(�L�?qI��a�^Q�����X"=^i����E����iT:��m�c(�A��� ᾃTDc�)N�	�n����-}���Y+�`yV_5 �뾝~�S0O���ݻ,jh4>	�Y:�\׎7� {Nys����ms�����I�>��h�Ilh\��c'�gy�8�*�G4��Gb��{�U+rV�qX��C%V�7�yus�sDX
���~;�#��.�m�=G@�ŗw�˛/{����ɍX����̬�����|r�Y,;H�O�	;|H���i����Z��U�W�@�+U�ܫqA��p"���q!�X)g�"#�<6%'�%-��s@	:�@{i����.I�ZyE�=�n�dJ0}A7�^���T����RA�T��7�4S^��������i�2H2Ȝ@&؂��ƽ7E��K�A�z��̇�41�����gm�%��Q4�
^��#�xY<��e�@SfPb1�ۓ�hA���T�s�J��V���<�گphU���7�ˀe�����/��ǔ+칅�>�T�@����3�^bu��/:�C���_�<�GF�n�=6�G���.��Ȅ����_�{�$�g��bv�?�����9�
)?X~�K@�'��TӜ's����ꂄ�ܪ^������t�>��u�-a���CX�V��-��o�q�&�qq���]; mx�pC-�k�^TP'�r� �����D ��2 ���'��Wz��Y�9�v�8�M����s�;�}7	.���Z��8�N��4Q@�FK1��EK,=QĽ�u�-�O�3̓���ӹ�[�}cJ;ۤ�����B��~9���Ey\u:&�ۦ9�=^��=S[�8e,;N�i8V�<V3����DwhUasB�x�E��:T�V��U�7���b����OW�j��K�6�R@��p��鞯m���`��6^�$�ʰ�D��)��K�?�&0K��a�h�UyQ�J�
A�"4tï�8�\����!j`�+?iE֋~���sqK|+{�or�����M���#��d6"s`Uʒ ����wb�f��f�
d����̱����%z�)~X�����(r�=�$FN�Dj~�*����gY3���gC�`Z	�J97�z�,\3��6�" zH3u��Q_Stj�Ų��i���R��a���j�*�F��?e
4m*�֦�@_ʼ�9����r�^�q�b�P���{���p�3Ǜ8.3�f�-v[����6GC�'A}�[u5̰���?F�ҟ�<e�}<�z|�+P���R5�J�z)
O/ k*��Z��̏h���y�xA+��7� �atN=^�@R��[`�qV�;O��Q��W��V�������Kb?�Ε� �^��Qx�c����(���5�&��D.No[��/��U�`�'��PG�H��},H��[��*b��t�,�hLh e�p�?tM�堠i�6�tK�L7]�D�C����Q�ʣ�_�@��n_B�Ԧ�{	�P&�TS˛F������l�)ȧ���&*Da��j|A26��	ˬ>��������N�CQ��	�ME�a�6I�r�|��D��;�d�ds@�mfb<x2*����=���O��g�7e!!T�򽳛`!�Όdm�6��/���e�H�k��|M�7R��髂=~ɺ�����}u�qyƅ����t
3T��!S1,�6k��fS\���c���W��2�[�W�_����)���� s�1i�r�ʜ��5KS��l��yѢkM�V�:�r�iX�q���/�^~�B� �Jx�I�|�de�{;n���,V��i�d5e�	u�Q��Sn��6���X�A���C*��]�hL�<>��u!��X0��>'�ݠ���l��� 97�}�T��zW]H �?_���_��~��c�~,L_�7�zƶ����V?C���θ�ހQ�Ъ�a�3�t�����>ۋ'���3�r��}B�%J7-�*�1{�U�7�����>үB!Ȭ�R�IC�q�h>5j"�姹u�J� ��4$�+X��0�+ �ǧ�Gx�1s�OD�8c��w�+�!�����̱f97xIǼ�/V�7}AQ�&�9�F�G֩B�YR�+k��R�tR0S��<��s�/lE�,Wr��'7���l���~��g�o\̠���%�����g�C�\������-85�~��b�X?����	J.��:[%>^����U!���.ߓI���_	�(&Ί�ߒ|�pȾ� �2��V�˒�P@�t�֘ݰ�mi��,B����t�rP��ծT������Z��;�V��qu/;�5�!ĮE��>3�_\�,'c�|=��@�^�|�}�TG�xG��S�ix�������V�h�GC\nf<�r
�j9�Ͱ�3c����N�\����]��v(�mp�ƃ��~/f��_����?�5����X��P�<>��t�11���.o��ASq&!`���e�����?����UL�r�%^r�Ӡ�
�#r"H��7�'��t�9D�����v���x���6�<�ڎ�=�	�m`�[�xJ��"5.a�Kj�������b�0E�.�+��6�B�ә��MgH�M}�)��3'�7���<xT��Ë�'ʛ�jG=nrj�Մ�8��q>귌�}��U�$-�f���a�!�����G�1os�m�
v��F�����Aj��Wo��JU��n�a����6ZsK�mȇ����߄�is<���㊱8�R\G*��mD�W�; &�jS��9�]d�g����'��+:�����4�X�Dukե/ڱ#���M��ĘH�?ܣ��]CW��H;9Z�}=j�X�i%�Q옯�NouX����wAr�%�x���^^�7K�������p|4�M�O� �*���c1bpSWr�L�A�ٛ!��7��F?�ޡ�ęs���Z�����$�0�:*4��:�	�ȉ�K���M[)֛P��9��^�$I1���#�1���ml��R�"��k{�6	�}ua3�n3�E:ǭ�T�ċ|��V���\��,��q���Y��K��S��e譙'��0&YO
9$�q�q��-a�Ktm}��s�棑�Yn%�EI,hPј^>���9ڦ&dv�-��fFሂ���}�oK�<�����k"�$u%E����6�:/������IP�p�ɹô���z�A{�ƺϪ�v����@����P�Ǻ�Vuo�M�޸�ux%��UɎ|]T��V�WI�#�J
"�C�,����F3��z7qALRķؗ#�t�p�M���ax���a��� C�i�Sm�r�$9]�s�l�(���������?)]���s����.���	P��y!X0;�������)�u�4{�����&�ȟ���}/����Fo��BY��"Q�̓9�_WSp)%�̵#�z	Β���9#��3L���C�#{�Q��A����(��Y0��3��a�1�I-q��KFiS$3�לϨvh������t, �V_n��GǦ���DG�4�j�<6�$�� ��5��(yi ~|h����)� �Ħy�y�N!���S%3	�֫��p�b���.pK�:�A��{?1��sE-�x��d,mf� O�e.�xXJ����n,h˙Pd:�&�l^��������1z9H�V��V��%^�W(zO�W�8ʧ%I��޾�.�Lq��Q��Ǚ&=���Tf�������>S�J��W�U=*9��;}r9�./�ӫ�ѓ���vC�#!�K.Fi)����Y��Hő�pQ�p�)�➗�pT?��Ju"�s�/��`H��i��^�lA�䡜� d3K���}q��չ��b��B�i���Q0C��+����nr��,\hW�
`.�>m�`"���` ����7W����6�/ C��ž���r{jo�0sT�f$����b���)xKR�;ާf�ܿ5��:�Ɠ���n���t#_��@��Pe����|)�(�Ơqƌ� ���=�ԘhtY�����#���.o����f.Y�ۘ�J��^����$��]|�KQh��H��h�Q@����������+n�����u�CZ��vY9���������i��f��\6=�>�A����=F���t����S�� �q���߁�K�M3R�=j$�H�'��J\_�Œ�DH ��ɼ�xq<��+�,��վ#*�c0�̉���C�l`�~��/����� 5?�{	��j��� O�#z���XX����zV;�E�1��|�/5= ��PiU��XtLcxv���#�x�*!�->�h��ZԜ<	-�L'����MU�c�9�6~Y+N�p���[3���&���Zu�����$Z�|��$,�P	�
�ŌH'f�3C67{5�����c3�}w�"%ע�i�A"��
"��7��������F{S��W�G,a#���7q�֦�ymLx��ry"{�b�`���;�Kj1R���������L4�?��.�6L#݇�#�	���g���
�	+��3�V� u;�"}��~��2�L��%�^9�ǥ<c_�� �r;����jTŮ	<�E(�����Ԉ]D�$�6��L��A�!\Z�z��v����+k_��\z���茏t
.��&D#5�����\Y�g��8�2ip9��i��9��P�?^�c���}�iX�?�4��_4��Ƒٛ��֜Q���ʙ>g6�6H% ��Wmc� Ȓ��&n�c������&e>�Q������z���9��e��- �����kDf�Z��-T}��8B�8sܷ<��]��4�\+�t�^<e�Z2t�z�fѝru��� �rAS�K��$N�b@S�7'�q�6<f�4�RX���[������G���ވw��ޔ�<���򠢤C�r�ޘ����oH�;]�կ��OY�k����X��|(�'�M
��ep�v֍��躯� �y��#s��]#'4ф���Y1h�� =(���W�^>G�<k��k#<��nc��A6�
�	�����(����@�O�h#B Y�T�}ĭ�	5ug���i_���SϨ�-wН�*� Ȥ4���a��?�ܯ���t���R���`*�m�W��gں���C�pZY�֌P1����
�6�(t���IV� ���p�U$�i0CU�ӛ	9ը�o�8����Ĭ��AI���
�/Ƀ0)�o�V������{�+�4F����`)��A�����e�,�j�=;�?�n�4oe]��(�A�(m���o��W='�d�J��� Qw�BBϰ9��\�A��S��5~�s��e�.tIt�����3&��}	+gd�\��em Zk����J�!5�\�9$m��U*����+���U덫�f�tp�>�Fh!!] �@��'w�`�9�{�گ�7)�k�s������I�ᤸF_�c��*��h��Z�֖W�Q����I��%���pt������"������z����A�R_���X�Bt�\܇���g��aca�Pl��EDTF�'�$��o ~��
��Z;d��E���U�Z�r�v]�U��!�����۽��w ��*��a5i5����ъ����@�<|�15�镍�L���u&KA���� !�8�Kx���~X��\�J���:묢'W���Y��:|�%cҕT9��YB<��A��[�KF���S�|�f��&z|�^�C;�`�ԶID��n��4�&�� 󵰅����Xr���4z���[&��W"��I�O�����J�{��b�"V�XQ����;l�o$�7�� j�ɜOp��0��bE���R���Iz���C����8��.�	U�D�Jt�oL#�<oȕ�eǑw��7w�b�o�lXvFp�E8`%������7��|*�dW��M����ʠ��є�R�"�tm^��B�m�� ���L��{K��/s#YpW�Cs�y��a�m@1�u���PNg8a	�c���	y7���c�F09����^�}��n��6a���r�m�ľ ��C�&�D�����6�����G�,ʪ���4"MP߮�X�ԊJ������;h� �����b�pt
���v.D�Ƽ0d�(���)O��\d��{ހ�3ٍ������
ju)�~/������3�\j�.�8������~����b&	����0��O��O�Z�R�MƵ� L���b��	�Bg��Of��R*��x�8��us��^���8�Q0(����9%6f�pv�iY)	0C�?l�]Sn+'.a$���Ήj�c���[/�z)�|Mn��=
+݄.Z�lS�*"�~����'.g�ݼ�ʻ��r0��dG�ջ0o��ݒ�s��i�7!̈́�{��r����~�T+>j@J��*���ZBZW�gXm��lur�oQ6�}���eD�O����1����@(r�q�~��e*�Q�p9�1RT�q�����
����RQ�_X�f	mTl�h!�d��<ʴ3,�T:�y��?�v(��n�4N����� ��H@�R1�ms�!L�:�,B� "ZI�џ!�~۶I���3��ƞ�A7�fKs��GP��E�e�閊c3���o0�ߨ�|��F"\�_�4e&������P+%���f��+u?A�#�x��(���ቐϔA����i'ʕ_��U}(��$~��C�/@CuD���������L�˂~��@��b�f~_�7���[Ǳ����8v�"���3�%�qP�n"��k�0~�⋢zU:F��-G����.׹�r���y;�P��H�2��H��1f��&�.y�P���(�ݫ�[xeyF�|"�D�.��wLY�i�� ��+�ǀ�C;\A�6��'t芷Z�I������*\�b6��t�G[�B
��{�g5"(��#SS��T8+�ve_b�m�-��Gc�)�[�_��&��i�^G-��J��wM{|
z�D�T��x�̛�Vt�=MI\Ҍ���r��i�T�f�7	%�Ш�~�0*O��"��\�7���VJ���Eh
w?�EM���`�Oİ)�#(YR6wl5��<�TŜ�	��NdTQbQ4���D�����΃�������XN��	[������yo,k�噙�v�u��U]�/x
�z%���.V%	�)]Mj�����:��Q�tZo�i�����@o�1�"�Rp��W�f�O�B�͇��Z�.�e?�N�q^��R��S>���=�s�Q��?~�<}����Q.��B���"���UeG�D`D���G�h�t�v�ĄG�2٢Y�%"j&������_s2n�ڌl��������h0�����������6eK<��<ꎤ��	o��5�9��眑����� ��_m94�]�	i��f�<_?\V��ഠ,y�ңx�致������k��������3�P��v1F:9�^�K,R�Q��J �k�ȍ����u>xg	�50f)Stq��V�k�z���	�2v,�&c�N��R��{q��\�q�]�NWNw}̵;�5ڡ��ν������Y5�p_���[���uɗJo�&��?;�@9-g��G5
�PJXS!Vo��+a���w����b���aV?����M!Z26�];C:p-F�³��� �똖�u�,�Q�"�/!�k(q�S�ڒ��$�y��a4�򀓡���5����ԫ޼�+5�I���͟{�\��@��v4�'�C/�0;�`�YhwH�	��D���1�+�%�R�ȿ��w��f�����§g><U�S��T�uY�-mZ	�������H��e�$f_O8����v0�	<w9��p8�k�4��H�2/{�����FZ�pg*m	g����W�Vy����ֲ)k*7�~�L07�D���>r	�k�h����9����(�q��H��M��Z|K�!��/3U+No�o�m�����˭l�6I�|��qD����eS#��Ftho���	͘�S}i�4�26S���E����1��C�b���sZ��/��~�:<Q��*����Ek0G"rJ�b�C�r����ri#+�����c��0i�I���S�8X�[�\���r�㞖|%�X�I�A����dN�[�X�AL�8�!�QЌ�i������,�}�~���M�)k�I3�pJ�t�\ew�aM����ؔ��xҚPͻ=��������Ҁ���=
���%���)P¢���@L���)��M�P}���#+U: ���Q��@�A+E�	{a����[u�Z�VNѭ_�`Y�����X�(���w]@3B�U��j87?�����VCJ�֬�ɚ�MF�#̜B7Qo��K)� �9@�샕Fh�b�qnFF��(�d5$U~�g���"�o�S�8)ÊOVv�,w,��|�[^��M���M �k~�*�Qz�"�M��=���1[����󭫒��AWrL653eqy�]>�M��\��ݯx)��q��!��7��&=;2|�m3iN�Ó�T�r^0�x��OJ\�ׇ�m����5�_wU��Ls�^���;���7Y0�
K�\��r��#=�kO�3ǦJ�Δ�4��/���oˍ&F�`��I�����e�[�2�s�Ξ�5��mJ�|$͆P�st%�^8W�LŚ]6>=��	��R����dΓ������g�1���^�*�*�fSx���/,I_�#��DK4��Yn�%X���=�J�A� Zl�!�qh�zK�g� �1KH�;DG��%*��I���{���"��GIcG�V��[����J P�(%��5�f&v�i
Q�U�H��j7LR�vsr��{.z1���af�����$_9Fg�c��2L�����$l���#W�W2Ae�������W�񀰂ZM����3��M��Zˌ6#��(��~^�u�,]��-�uQ����IX�V{�F����h<j����:U�r�(j���Su�hX%TFE8݆��a���9��Z�VHS�-�`�%��0��*�ʊXq1�����S8����� ��0YI�^I�ߣX<P�[Ì����S�JF��-w�Lq]L0�7���r���V'�U�Ye{��� _
O����suV�������-�A�[ž#*(����i0����E�),����jM�u�v�k�jz�]�t�/��,0)��O��K8� ��
�cNp�&Ɉ���z�1�:'Z�J�^{(��� ���_���1ғN��}	�8ʒ����^�a̅!�g���Z�"e�!(7A����N�C�"@ȉ���x�7��by5ARO!io�;+Ȝ�Gd�Z� ��8���FN?��tEٞ��h�Wt�!�p$�����s�a�^�L���$9U��P}�A��ʹ�,ʔg���s��Ǧ�*)�_����G��-㛺I��T���m	6��Y
U°�~�.�w�@<Y@+�	�-�LӁ���'k�}�ϯ5k�+��$]>�g��������D��Z�AB���+�!yz���0_�|��d�����r�@�2.�k���,��.�^�}ȡ����-�����㩛c�Zm���	����ha�Y�|���mw�>�,��9�e)�	�y�E'�}&6�l���	k�b�F�J��߾`vA��XS�֕�wn���.���0�qy�z�J_�Mc�.Z�D����C�`�i>���iR�!�[,r��3�������7�?J}����*��ŜC}�QJ|�H"���JQ0p[1��E� �ܧ�������[&no۹E���ּ�0�!��H�"����6Q��QX���0��� 
��1V�U��-�K��H�E
��p�KԹ����Z������Y���E��8Sò��X?�,����q>ؿ�6=�̰|U��<��n�{5�(v��'_}
���˱�aɣ��A
g���_?N�^��2��l�x��BΞ}�Le9��|h�l.��=�����Sn�F/��ұ[������g�O�����
XU��ڠ=�d�2�8��s怱�ph��y��^�au=�JT ���a-H��S):m���4�t/@�����ѹx�Y6w�{p�w��]��S�`�,nmZN�L�;�(	��_~Hk['�9	���?�,e�a���0� ��Z-c�tQ�X]BZ�� �d����n����}�lG��xĭ/���P�u�w?�a9���Z
p�?���S��e��*�kw��ZA\�uBd���aV(�=�3���$�lHXƲg�\����6�K"�sa�B��\#1���DX�,����ȟj[���7�;8�g��|B\D�Z��^ׂp��I��&�7b]v�xri5���ӊ		�z��ӌ�ԏ+�j�DVvy��U~^���Y�!�4�q�6���� g��:R��t�r�r�G��5>]�P�kgV��r�nJB����vI�U:wq�xNGĄcH�g�]�Ɣ�^�y�����£��|9����2�b��F�p�t����e��)�s�O���E����U�*U:&�{0rA���.�3�Bn\��58��:���4�/"� ᤾�L������F�0^.�j�n�E��	�q�=+;e3cSO)��c(dM�<~ 9Y���>�1���\��@Cpʥ���`�.��Yp�Z�v��{�a��Q6r/S�t� 25�%8-�(f8
�1d;>�5��-�)k���孄מ}�9[���ߩ�⽂��/����w5���V�v9Y�?��gWS���i)NI,�5BN�!��x"��#Yn�|��ȏ����E[��EO�剿
���|"���Qy��J	��,m$���4S�9�w m�n��:��h;��WV���!�ɩ)�/��ў.����N�o�4R,��}��VK�I�9�{d!H�[�C0�����:��h��{��w�a��\�j�����Y&FL5�y��<8,M�}��x@vC9�����Sfz����,���&p�����̓�l$���ى�a�N��ls_X@���^^��X{���ȭ��ʏ/�K��ŷr��$�j�.e��ʲ��N�_&��N]��\v�w�ZA�i8�rY���`���\�x��Ô�!��_'��[����g���}��\��#�fO���ͨ"ý=ju���;Ϊr�פ�
�#q�Ԫo��]�c	�Z���?��^��M'��smw��b_�Ok���O�j#�ޝ	��e�i�j�ɦUY�L���ƌ��V}B*���*�� `!L��a�c��ǅ.Fsu
'�;F�8�^���{\`���Ba9�S��֤�Z����ȳ`l��}?�=�ĳ�j�R�O��_O����rO����!-h�3�
Am#RP�Hf���>�P�R�SP%��?w��{E��*]�D�:OG�>�{�|j��,�)��� �?}��n7��K��S���Nhmz������2�	��K��}H��嫰;�~���
�&���0��B�o{�BM�.iX<�u��`#(�C��_��_Q�v�l�CNA�������e�F��!w��q�=d�*-�����H6+C��A�RM�m)�q3,�>:,������#U�SV��a��p�uC(�f;�)�3�����,Ab(�C=o�U�v������ɏ��oq}�C6�|�&f��ϕS�8�e��N�����a�Q�w� �~����o��%���^��_�@��l�*���)����Ns���\�Dy
�]9��m��7���nj�xY�"N�/Ύ�uR��$:��@:����-%�Q�`pa�����Z�m^���0����F�
�~g�tr��+�dV�rp�M~�=u�0y a����]MY7�o�_�Q�lE��_��نW�J8B9Ū�D^�O���uz|��I�V��4��$32FBt�bv�&����Sa�sB*��z���Ukfm���Y}�~8����i'��_�`����ip9%g���u��͚����g
��4!���*yw~��;�l�-T�BzKe�᪄��;��I�>��i��@N(h,./���x"Mǋ����8�yy`o!lAvV]��*���{�=b��z�_�(+7��5��k�V�) �2)����M�����ѐ",���A��ZOm�ٟX����K��l����A붢\m�MW�T�l�Vd�g�
�}\�g��mW�Ʈ։ڳN�K�x �.�����:��쟾J���V�vR�׳���e:�0JSBǒ&�)�~�����3iy�qH^��Xb�����F���߅�*�:k��A�)�^_�p�� ��mB�=��q2q���(�2�D��Tv����zS3ïi�̣{����T�Ș��@��.�����'��V	� ����A�)�wtB$ܐ�Z��c��v�����j}ో	�V�6Z��9� 8[*$����rA�h^ Z��+���C�y&���k����8`��vY�^P��9Z�U����pt���	S'&%�,T�Yש�Rc�\��j�p,���Z�!@}��K���Ϙ2kZ�mR��rPF����Q�(JEhm[h��w�k��7�;��W8pA�=[Q��}Q��<�T��1�n&`Z�>`��?	�=� �yȿ׺ ��̏�b�Tp���l�G��d�@�G%�I�������!���{�w��*Z��E�ijF.l>��͑��*ޜ�{R � $��+�{;X[7�xu�+6 FZ��j�f�D'I�T��i��I�o�5n_��l���u"�c�㶝Xu�|@{)�H%*"�����>IΗ�7.���N�:���{��*��U�'M��jBa��yy��ɎY/�H�"�0N?�D��(����7;`+(nUX�t�پ��`�煹�S�w�G�ri��ȼX��Z�;W�}D�\�����{�ׂ'+/�a��q���'�I�櫰(�/p�O|
�Z�_��� �K�����B��4@j�c���g��mMF�wX��{E?�62��Y�I����f6�|���]c,Lv@���m��V]YeH��{2;��]vD�bR���?&���6�Y.FM벲��Cf�<���ۨ=��hnv�T��d�E�NZ�AV�z�oj�t{�~՜�;k���n!rK'�hJ)��E�8ȕ�qU�I�Q��s8��5{��C�y-U�/����:"p��9۠�7oQ�������u�`( �o����-��m˦�U����n����k 员�����x1#ᝂg���S/��R���$�%V�K\�Tr����z�S� ѹ��ƏPW��L���+�����M�)D�XL�4���㧯�lTaqͣ����_Y-���o��P����1yz�����PVY�ކ��2N�(����r)K��nú���Jj@����oT����-@"��٧b ���|�����c�h�)��u�Je�k�)�~L��+�<X}��FB&U���| �gf��V�������{�/�NV����+T���o�5�[LԳXC�	���%E��j�7h�����~�wa;��f9�u���	����A�A>�צH��0���ȫ�<h��Xr��nAB	UY�,H�u�7w���u�/��r���0�z#��Z�=J�W��#��Nۋ��l���F,֦P��I��Y�QS,�}��뾁�M.�,S��cr��3��Kb���������v�dF� ���NH�r��B�ږ^v�nOX��%�O���ԩ���Cb5ڜ�,/���U:���Z�+E���(Ņy�ֿ��L�t]�u�/�F�v��1X݌�j&��!�7�&��m�zwzm%�e���";?C�j��L�F��O�AO���x���@P>�Z]m$���>9�Q8%�����8���+�r��J���a�b�����6��nQ.T�z�)�Ν�^���`�;#�W U]��.�:��nt�9�-�j�Z�P�R<���-�0'!��|p�]���<N���P�v[���ٔIP�� �W͢]bؿI?�ҝn��{�a�a��	�B��d� �<^#l��X��G2�D�uL���q���y�	���޹�V�K�^�G��z�����O�w����,��'b��_ �p5��X���a�s��X+g��\PᎤ�B�X�yI�@�V���|N׫�����8�2s�I�ĵ%)M"�z�<,KSH�b������zZTIq��j< �g�`��f
o�f��o����u1�c��!�D�8f�{ݚH}���.�����GmS��k0~��hwvǊgq����e�d06)z4�~�����/��2�8�f�JQ�O6> ,�]���EB �g�u�+X0�p�*��^P[���^vޅ���(�g�,��-m!e��ȃ�I4A���1��@����	��3��w�na���ŀ�;����g��cD%��OwQ�Z/���	���j��QNHv&��,gu[gVnl��׻�8�$������wLq��h0&z��;�
XEla���{��� �?,���*�>mqq�X�	uaN�otQ�q�b����5�3cQڿʡR���]��W�b6��YrH��DL9���a�:�=H�;������r�Ps���z����m�-�W�̢�e@��=!�ݙ�#\h^㳁���	G�����a!_>���% ���]�Y��#)�^��=$x$���V�ny�Ҝ�#�D����7�U�7�A��S�Gq"�~bmq��6*L\���־�\%�j�6`&��D�r2"<9��(f-,��K�z+���ua�2�Zda^P���B�
�󝓽�b���/eˇ���9��n0мE��x���f���81%�T�6��u6q�����cUQ&���C�g�*-�j4��Гq�	E�<[E����4�*�0�e���@T�vz��t]o�oY���ʁ]EX�.�Z
�����w���̞��;`��K�Բx�ܺ͢q��߀PR�Q�)��%�N�:a:\�r�XЃ����Z�C��
uZ\�]�F��P��f�K��������,ι�xO�x�YE#��D�4��G,{���Ohأ�m��H� �����t+����d�١M3�^�Z��&;t�9?�Z!%d?e�v�8Z�~K3�Ëe,꜌�l1�7��bR���d���'x�^pr��ݘRl�F ������FQ��=c��2 襝��[P���H���g26�ŃR?C�7rc�5f(ޯf3��^�N�8T���+u�n��k�C�V��O 1)g4�'6ȇQݨ4����+P|��G)-�e#������
�5�d*��}�M�g�c9B,��U�/k��^;E�v+��H�s�-G? �q���W0-
Q��z�!�W��6b���v@�P�a�%O�!�����r6x	s�+P>,J��	k�]��3�iA� ��G�,�x�T�8���_��ˎ��->��G9��RW?�9I	���J+9\�6����úӑ~Lza.J����!81|�]�������oQ����\N����~	���u�zy@6d�L��1o�Xd�7��D�'���c?Fk�OB���9q>��>�$o`�� �&�W���I�.&����-�S%Eam�_�F�}dg��=���Mֲ�/
^�I��w�f@��Rp��N�Ιb{_�RĔ�i܀�&]f�O������3�KD>�:꾟�F��Y�OW-��W�ɣ]
�����'�喉{|U#,�RZ�x5�#<%�ۭ�ض��Q��)�(��^�ɀ�2cl���L�-,ˎ� ���<}��8+0J���H���5,�Ⰴf�-3	Z������<FOb���h{��Iwމ�>� ♒S;_p3�+���R:*���K{��jZ㊔���۠:�`фN�8�ig����p�Cy��v�Ǚ-ǲȮc�O�r�?�����x�T W"�R���MZ=br��Y���LW�G+��c�v��Āv� 5�t���ڎׯ�+�Gc��:��ɳw�Va���֣7)8&��	?��3M���f� �Ū�D�r�l�nsщt���b7�7GA�Q\�V1���{	�R!�?��9�2N�0{t��0�p���|�,z�1*���oo�_�0���YR�|�J��V���(��/Z��U�X;�����xJt�1h7��p�1��lk=ב%k����̷��ľ�ܿxe��q��~Q��=F���<��� U����*�hkV�0�oqpx�Ag�Y�2��@���Y���"���)�C�ʪͩq���u;�����=���}H�:���7����������6�ʒ�T;ˢ��*-����n^.`q��h_��:VP�?�����Ǣ3�S;�����B��K�~A���y(B 7 ��<��j`"�1�%���8<ey_i��s-m��آ�+�O�n�m�P��b��y�Y���Yv1Ak��`S�'����
=��D�oA����NM*��Y��=ەZ5��)I�"���*�z��L'mZ�f��m��b��⬍mt�������LcM�B�z)���EA��)�/:ܾ~�ڮ�E-Y��Oω�V��I�2���U,�ms�����cH���@�r��z�9Xr���֚��-`r��Z�GG��_v�������@����j�y�ǐ���*����4w�>���vƈ=n�;�!����Xf��Q������Hj:?��2�74��F	��1��y,%�}��Ҁ�B��ͣhg��=}��9ߖS�9�}�ܵ��Ȏ�������H4gC�򦢕mG�q>d��9b���|�Fq�*�ȏ��<�IZ���Z���w��L5�Q�W�>t��jl~�:�r!���F��7<���d�E��˯]�hT�[p��${D!^�Ѭ?��kCW�H�c�������W[��M��y'$��I�7D�p��E�h���f��7�����kn���!s4���Om'�+?�*�9+5�Z��i�����!^�O�J���u]�&!7Gڋ��B�`����U��GW�E����Op�����rOX���]o:�����%E�]d��������0Ϩ�9�n>Y1
�A�7�,��Y/(t�˳A6tx^|I|�ߋ�Jܝv�E�.BYZ��쒯£7�ʮe�M�顈y�:����Bd�,������)�Օ2mܪ�u�@����?�R0�����)��آhz��k�;?�'>6k/K_s	Co8a��G��|�Js�8�L��U��!�:�`�F礎�Y�Oc�����E�Ie2��&���������P�8���T:VbB�h��ë́���(�&W���:����L��� ��m3�l�Z9HaaB��	Q7=�d���6�R��<e�W�$�����80�y�ͳ�o#�Ռ*dd7��RvY?�8=k���������]�9����VD�9/��+�z�Pk�"��	R4��K>)��xm�nZ�Kl�� 7p�B�UT@�R�0��F�?�u�(��yQ� �����jX�u<-���n��Z�x{��@G��s�k�s�?��+���9GL�"�7G@Ƽ,��eo�c\��(�y�䤴-~���qȏl�VM�S��*z�	��_n�}���ם_a?�W��!q�$�wL��<v��)��l<��p2�������D!�Y�'L1��v�C�`�(�_h����d�1��(���A�N�����D���+�S�>�L�m��������鵔g��rn�������|��`�W����#smƐ{TizN����
Va�/��Y����fY01��-��������>��b�Cf@?,r#9�b�j���S�!"��h|�����'�w��K��dȩ������/0X���֛u� f�CN��/���p�gS¥�̀S̕����g~`�%����B�m����ɱ��*ymx�����H���:�����S�oC�u��V�(!}4��I�J���&��#�����1L��K�'O$o��<�g\tF�L�� �Q>:����6�޼��aEC.y�m�1�_���٥��b���Ǭ~�H~��cJ�~j�"�dPe��<&�b��TVT�4e�����(h�. Q��h�$M�ỹ_���&�fe��j�D+�(-�dl�MmE
9��Z�hEu�%����� �T�Q�74b�ҴS�`�O�7Q�~�����Ր��Ǉfi�5�qC��^��Z��0p���d�lY�(Q�*j�I���7R�v��hm��١8W&͒�Ud��Y秗�Ri�$x^:L}�a��k.;�.ZO���_�#^�}x]OyP���m��Ȥ�^dk].��Lw���'3�t�����@"���`dXMI/����WYM�Ϯ�@p��J
{�+F_m0�=a64J�3U@!.:�H�hڹx� ���|@�=�A�0�4�����s0r8�c��5W��]l�Ȑ�ڐ2��h%���rɒ��U�	D���1�Ƨ��;t�2�c��1�0�JH����d�ӈ8E��G����RH*2�"?Ѭ�OT��ʵ�S��P��,I7�o.{�wl��)FCOS�����^��������C�
�&�ۣ�*��犎�.Är�&A�~�oy=��*���P	R������4S�&kd���n`YjV�df\^����v�)��j�w�L���������R��A;(cZ�5�L����O%a4@��Z�G�P��OQh��?skUkwwy�SR�gم|�2f�R6��~��`U�G� �ײF*9S�u�e�m����ͮOAv2��ͭ �߅������ﰖ&�G:G�h�i';3c�;�Ӣ~�ŀ��ww�@^���:��-���y���-�rXX#���U#A�s>t@���3��ِ"50��\l��\�A�˲��F�����I�T|YϺ�*us������h��W?��Gؙ��Q��N�{E������b`!�Z� ��*y���"c�(2p�т)>.�V�� �:���`��IN@�������$e����0Pu(A�*�e�_�@lU����J"�W����Obh碡��[z9�8�L���8�ޠ�`Z}�����Pty.����E����T���?�=�V�6�����<�ӄ���BU���'��g�֗P �	}���䨫[g�T���W��y�ʤE'���K��5���EM�\��O3B��g����j����a��6�At�D4��k6@�C}� ]���nKEu������\���}g�+@D�r#N�I:�p����o��{$���ݮj)��h��l*2t�����q��j[y��`a�ke{{��9�A2�����A|��
f;�H<�Z��\8ꖛ��lw�s�v��!`�S��l�b�~ZX���W$KG:�A�\��Я���<��]���Ά@�6�rs�ȻruAѥ�h$G;�2� ����Fp�(`�6��t5���l?[FL�婎���� ~Re#�v'>�A�'�{��:;m���]���o=���f&Ve��u��L�+�?R����L��*��Pz8����T�|�� &�d.�^m��+��p�b�Џ������*򳮡�������l�+� �0<�bO���`�Mfmh���FC��Zo���I+Jbɪ�^��O�7���({�BծcյA���ʗ�a�'�2
�\�����8��X;����Қ=@D?T#�kW8�,b���o.�?��|�p�$��{��`��y���Vn���m�@�2�3�����%?f����%�ͮ�:Ŋ�sRY���s	(K��<�Y���@�dˢ�m|�C��8�	!1r��;�f7k��_cZ\'B�d,����{Z_�V	6g�ϕ8�2	/T�_��kb��\X`�����.j�� o�Y�Z��B�=*��U�4|}w�1*�v���9n]�{0�ECC[.�wS:����v���:z ����iς�T�� I�QTƌ�۳q _CIZ�����L,��G=)��<�`c@9�����5�����]u=�jڛ�l%��iO��)d8�zN�4~���f��H1&� 	�r����D��>�0���0G�pq����ȩ��XDd"��!�m����Ll�]��0�4�y�a���$��9���ȏ����GI%��Vɰ@j��~Gr�����8�l�p=(���-G~��`�R�e�SHL�֍����/,�9R��1����т�;q��Tb_ωP���WyO_3+�%v�*���a`��Ⱥ�g�CM����*�����BOh���󦢧�b�j=�*�t~�1��(%�\����O��jv,�=6������A�+>�N�5}8�{i�K9�BH��?� ���ܑc� �?��6ɧ5�� ,qV�cEqw��Ѐ�C��1*�K��&��7�4o�岧m��:����2
��`�>�ԫ�*rK�6<�����kQ�Aw�_؜�tƁu`���R}-��i��/�߾�QS ��A �
�+��
�?gTybEЛ���S�7�&%C�������eFΣt�o�X"驈	��9��m�o t�G�~��b��'��&<���^1���#zq�Nu\|��OL׸���r���ⲳ0��Z��#֡|�P�i��Z︇97�*�Kc�.=�s��Z͝@G���z�k@��(8��6�͡��m�{�s�~lA���JGΎ�ɶ���x&�lrي��Nj��-�B#��i!��3Һo㫃��y{�8sH+pnM��%����s�i�gw�>�t��+tf(�h���>�O�i��J3�d�5.��*�DՍ��+*�]�y�;��-��|���:���x�ԭI��Y�{�S]6#�?pֳ��,�w�BM1�ɖ=F�}�<MO�.���7�{���!��ِ\�>
���z�G�r�(��V�'��\%^ۓ�F?b��7��p����i���ףxR�� ��H����T�/ڰ�i)�~t���W��ܠ<����N�)���	ߔۦ�fY�ST���Ņ�څ�4�_eYR�{���"�ե?���9i�t��and���_��s.�ϧ3��*_S�g����_��������6�W\��~���N�9�V�Ɇ؝�{���w��v��8�`�=	���,�W���t،}��;�-�֌�51i��qP��F��([����E�A8=�BB���j��#���T�;�{���3dJ~�j��.�����Ԁ!a~f	�=�n�=��#�G��ʱV��<vi��n�Y����v�b��#�\���#�L����]6�g�T3a��E�ъh�5��)*}��dx�I���d��-֍{�)�N|��i՟�;&&R������@����_ݰ��f)D���l_T�7-X�I1��k�A�S��k�n�\����fv"�o�׳�r��t�Mb�Gq� �q��o�5�vZ�����:�ϙ�8M��r���'�kk�+S� #���t���~8���짻 �@`���hsc9��~yF�u�Nfu��=��*a ~�7���U��:��Pc�(#�Ii�IH���t�_̰����.b�L�?=����������E�:���!A ���Y�q�0� ;[S㋯n��]���\�Gɬ4���j0�fj�w�R`�im�Æ�hR����(0����
VV[�5<��+Q=T�
1���bL��m�g��5'7�,�Z�_����������0���$��\5�\��r4����m�y�u���Apr��E-��Ғ�?�`�I*�ck�9?z�a���زN	U<�ӛܯ&�LD�͡l����
�~�.59i��$~pX�pG��w^�wd�/��:�߈ǂ*�����?*�y���{2���F��~����(�f��!^%��N�F��1��Ţ_J�9ِÇ�9���y=^x9šC��r���#0S�ꚗpS%��l )�,_�
?�-�Kn��~�6S�aU�N����'8��\����6'�`nX�k��v��h�)9�lѫc|�\�=��ۡV�����]5��Y��� �k�I1�#|��+����b��'B���Jt�L����E����?�KYc��<�@o�8�gc��8\UR��IrO����k�E0?�TX[��u;=C�����'�n�O�*��e���~�%� X>7�8��$vy���A�����6W[���gA�(��a�J��z��k����
�78&i-}!J"��q��?��y��#c7�6�L���5U���L��M�Ɩ�. wi*�`�;)!��y,�mhKC�z��;-���Gh�Nq��2+����Pf3}�Z0���ؿ+����q�X�3���(�Tt (mšeΑ��Zy��|�N��HI3o' �v���Y e��Z��B�n]f�x$���zX��PN��� ?��8nt��c.�j��f0qߨ��ōE�Y�ŵ�
#d�s{�s�2��OS�=�� !�Ԋ.6�[����%���_�E��I�1���᪦�$,��)ؘ=��i[B��Y:w|��$^���5v�d�>�}o�S��_�9�P<�x5�=H�2�m"�O������6�O��,s,Hv��O$hyR�Ǜ��Nri~.���'
�B��q�f�S�LE`�}�_\ur�w/�a���eJ8.0���N�QQ3�
U�o�8��j�)�p�<w����s4G���]ê�L�����a5oq�j�>�E�v��J�SǲL��u�����B1�|@i�s�#�$�3�j&Tq��`]Qw�w�9���H��kfM����jC���o���Ʈ=~*3�4B�H�;�<c�Ts�`B	�z�UP��WgK�u�����uv��������t݃�;�̄��������f��
�Az(��S3컢R\�E�f�m���9X�G.����5�`|A;�m�ɦy��R.���<�ĹA�Y��՝q+�Og���F��Mb�>�&ި�v[̪4��"�t�;���9��l0�)��Ul��#��"��w"C�X�
�'��+H�m��ĭ���$_:��h(}�(�E0�y�JКQ�"��W�<=E�6e&���%�2J��h��gI&��JT��	ٺ�'i2�f����a��� ���\+��LuP�N�Fq��1��g�C4@��5�Qw��;l}n�d�J�<m�Q2�2ns������jA��~/�	E�J��.�r����i���r����'��?kkrA���6�FWj�� ?^Ϋ��j�,3��e�)�[�+5�݊��JG��:�~'��o�H�R>	HϦ�2�v�)9q�g�\��mR(�������J� ���Q�� �#��޻Hc{��u�4����L�O=?z��(����ڰ. �7�rP���t~�GM�dy?+��F�h�o2_�~Xb���up�OZ�9N@Cws�Dp���P�n�h�)������,]'=dApב;�i�X�ޝ�9�3�����^�Q%<:g(��c�m�<u�:�H �� ����k������Eȝ��g�+&����� �j���E�A�c%���� �^�c��BE8�u`S:;6l�;q?]����W��9%���d6}^��OZߨfu�V_,VS0��б�
�e0}����^�mR�W���ϭ�NF���(�hO�Lz*UT�WDJ�1w�ڳ��K��r�->p�t�Xf"�b3F����%���D�0jDu!z~Q��X��ւ,ɂ�
�n�/���{�O���U�Qs9)����s�XՐ�:·�|(5��7A��p�߫U\|}�Y�$l��"Į|�t=��kK�r��#�;*�~�Ss����ػn����.�O�=�ٗ@ʱ+��Ùѫ��E0ĳ�'�=�<�t������ I�)������!<�!k�x8���P=>�P�͒��Q�9!�]��h�<����	E.���F�uA2+�@�s6��jq��^"���OeT���,�p'����	�]�pC��!9
n�������ڙ�4Y
�#s�sPz$�qY����H/�5�K�T�e��c\ܮ���^��֤`^�'�`�]��d��qCrMx(F��o��^��ANZր��.i�v�>>ۚ�,�� %mh�!��V�z�sl6UL�����!u=b	û?Cܨ� n�u�{��*�{̋����ʧr�;4۾t a���:Rf@������f����-��r�]��}�R�+9���9)��&U��s�����I��k��/�����'w�v�&�G*5��dbT?ղ%�3����%^�آ8C��R_$|y�t�B�����T�tc����Gs�֤�g�E�1ߟǳF"di���P�[:ň�^�q��lK�&���q�ePo�����y�oT�5t���2\�v��l=.���^�=4��3��J	�����7M��
^�p��=�^Ƙ6;�I���]�Ȱ���AhLH��T�uHi�����)L������p�D �r�;�7����:"X>��swVه O�w"���>���x��m�`��@Z�H6���a�j��/V ��豖{�����9�v���sڢ��f�.�e�kJ�pSrP)�R;����]j��v��T�S�h�t�ܐ�GS��|(f�>�TR  ��׵e�Y9�\JIBpO^6�s=�EwH"�
cJ{Q�j�A+��]�\����[�z�h�}H�,Ռ�B�����j:�j�W��x�A�Qu����A�~�4�@�r��'|�Z�n�ܪ�$�j4���)3���/F�m� ������%�{��ϊ|$�}��q7�;{Zs}�bp�������U��#��H��<ya9Tr����|W��8i:K+�O�8mg˖��c���33�����nu7�q��s�$��	�Xу�}Z�}��7����-���Iƍ�.�M�x��{t�9�>��:s�y���943�
���Y�(�Q�8���'�ؠ�����U� �M
�艅(*���a�f�%M�k�Ы�:���F6w���q��,@�cF8�#���4���&�Km�{|���-���6l <lK�9�4iI�.O�j	��3� ���	(oɼ�6�-<jG2�h�lE7.Cj8�b��E6���'�|���X�n*^�Mv`�,��������ʵ<#��#�8�фd%���g֟}w��v���1�mzQZ���/k�uF�D����!@B�s�]�r3G1v\�F�'��F�!����]i�]�z�(g�Ug���|M����Ha�$H����X��Yq��B��0U��C�8$(��X�鬤�z,��*O��ÂP��.�#���|G@���4E�`=*�:�a�E^���Ou�$WqQ�#���$�^w�)֌��p��|��K��[B�	8ы���m��4ɨ~��B�i$&D�V����G\D1�r�/�8����YS�TI����Q���v�_��yf<{��7�SJ.�G���^��C6s/���Ɍ�cέo��O�^�'��f��@w�E�z%O/	P��Ҥ4�=fz�K-T�|�����VT. %ݲH�N���'&l ',��WL��q$$| �Y�����2�'b�"��u�[a�1��k�E���m�T�d�j���h�lӝe�� ��6����k
}�܃<��RK��{��y��t����ו���jC��^6���ٞ�x-{�N;��h�����	p��͋�� ���Z3�Ml��f��Fg��Ʀ�ˑ��e
H�ÿ]K�() 3��������9�:�!���R,6����|Qp����xkZ��������u�|vf��9�D���M��ݑ�nۢk��G{t�I���ڠ.�C���˫�dl��"�cd�06A�|O���䥄���	B�[��3~K�<tr�%XI�G�a�_
ʇK
T��Nc�K?���`|b���8?Bk�:������8�HN�Y��G���O%�!�$FU1x��X#i�;AdB��G/�E����n��x>Y�291��˞�:G�h�t���!>7ap�3L�eW�X
�S_{aE����B�m���/�[	rDK~��e��7��v80�7��e�1V�f� b����

�|H��}��`�+���H���/�.E��C�-f=�00�h�)�b��Y�>t\����j/-ݔ]�ŽȒ���J��������R63ɔP��Dv��D�B3j.�Q�r�~�VV�Le�z����.�|�V ޘC�
Yc1��q�Ӳ�����!>�n��h�
��BPn��%���U�����uӝ�Z�6�W@�
Y��ȭI�hÃ�_A��059G�dO��O%
2��l?�!<��!\�D�Qd��%�@�J�YN�X~}�z :���H�L�9b����h�|�
$(���\Q�D�NS���+�-T8�?U)���Μ���$�%�����}늶F,�L�m� ��-e.���������~FM>��z�B��� /����}��U���e��kCʒS�EԍR��P��}�~�y(/��OV�Ƙ]  e5����
�-�RRb"-K�~<VY�:�y�2zcjeZk��|���O33\���ª���F_[���ّg�D���ߺf�^h���n����D`�:���ʰ��c� ��U�xK�c&�1� �^!L��ɼ�>�*yB��jSw��]�N�7
�C�;�v���ѝ&Z��X<E��f��|6��B��U5��a�p[��~��q��W �)���7K�^�ZʹIKebi`�:��;�7���4�]X�\H'W3��@�B�Oپ�(Ԝ.jlfg�����H}f��&�k���g���K���B�R�# .B^��ϸ��,�h��Hxq �� ථu�:	��#�u)>�y`�ԣ�I��s|�?���|z\�W������mk	*Lx�$s���`�M[���+6v��� +�֔HP�j
��l�kׁΕ�Ůvk?�J�ۚy�m	�nN!��x$�x����'&WN>���7�2�]�F86���&�e�����˶[?VW���������NI�ω�M\����.+�b~
e������j�!X��<k5�O�4q�G�/���BE�F��{II5<Q<a#�j$���!��C�L�uq�Qy�����a�:��=�.�圤\�:�ϗ6v��4�H��7Ћ�?�&XΑ	u��%�]�%+��s{
��6����(Rت{H��uR��ahJ2��)���|ķ��Q�y|�l0ͱ�m�.|�,�y��}��<��zu�<C�G�N���t��T5!4K�!O�<�l&��O����Ҽ�ya��ɒ��̷�\��$��� A����]�x��T`�	K�a�[Ry�c��Ԧ9�!;�Xu%��� ="�OS�8�A�*�Q��4^�� >�5��t/^u/:��x1·�&������ ����t�{���DP���4F��P]��l������0����9�D:)��c���4�����o)V�������������}Z�j�ũ!AX0*��f��E ���=�'��G�����5�d��?�kD����`s��I\:��W�|/�����m^v���ܴ�[Q;�<& �.�J�,��� �Í�a��18N_�'|=�	Ԣ�D�Rx�y�r3�l_�줈�R�W"�:���Ѿ<ޣ��0�7{��3S[��.�PՅ �HZ �g�>A���%)��8$������"����/Ʊ�MW�v��R��/ҿ8I2�/R�Ǧv{J�T��M�1\ �V\XV]���/�9k�
[�Z���~���1e�ӷH����{�k-�_I�*�������yĖȭBd��P��XC�i��J�yh8g��pb(��|� ��U������-3�/t���˔U�Fj�5���Z^"��򙟪W�N��#hO[X@r�e���p�#Ѿ�p�j�����J�ǔN�2}����㠈i�}���lW��^�l���h�B0�����ts�j�p	�D�ZR��1+i���I���\�	��Bf��A瀱�yX)F��30jY5