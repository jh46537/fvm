��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�\W� u(�=@=ͺ��*"%S<E�E��r�YY�HPb
�^����S��E�P��62�xk6���xL�\Rꟿ �>�F�#!�T��'�����H�X��NX�A���wچ?�t��RP��߫�y�cM?����`� �{��q�W5�l��pؑxߜ�<�B�Z"�7��J3�.q��9a.��,5Q��cb���L�?����#�-��d�~�5wY�q�nV��i��Ω��g���UvG���-R:��7��p!^	��ʁ-�����oQE���b휇��J_�����W{rV5�9T.3�w�2�����|���;�u�A�f�aLނD�r������00�6A�N�����(񆔣2ı�=܀��r��$T1%�7��ɎJGg{R��ԑu�,��I�.*���p�.6��	6aR���.�f�Xp�@�"p�k������/pAy�Z��"y�M�!-3��sŁ�VB~X`�zg���[T.�rGÂ�٦T�bK���tU�&��u�!�-?���(���P�i��*�W����A���Jh_s��he:wm׀FH�@�4
�1,)s�WLG����Z�I8_<�BOPz�0ϕ����
ď���vp��k,0��x�K�3wn���.�h�x��u��D�D��a��3��Ăe�#�Lw����3ͫ�q�~�CaY��Yq�ӠiY8��{;����ŧ�Pea�@ꏳ�h��u��Ns`pzU� p�>�Ĳ��װ�����͵|@ޣ��g�R�Q��5��Q�|r��7VzM�7��*�(�߯HT\�q�w�e��,���W�ODA�ף��3�aK��:TWW�!�D@+7������`�DXI���+�aĐ��zp>�S�t5���*�M�b��`~՟����ޮ�J�����&��H��0:�c,t��͔ȝ�����Q5�cü!���lJǮ���Dʢ`4��?g��T����d���\�u�y�l�L���Zq�e�x(	�M2�a��Ӡ��P�O���ٌ����	�Y�o#Ğ9V�h05,Mr)��#�-�$�]A4VZ�a�/���S�����|�vVZ4O@�D�_�ϰ$���̊m�ȍ\�2��Y�"sԏ���zԲ�'H}�~y���Ct�S�׮�ji�뵬�d��9I����磆eI?oI�u��ŏ?Ƕ2���F-L�L�Gc�\�[�ؖ�%���q|��"+����JY:��B]��Ti��3f�n],Qh5]�څ�0���='���!_?0��+�R���d���5B�:�By���F�5F�Ⱦd-3>D6�U��*/֏$+,C񧥀a,ʂAR�Ӡ"�J�"UR�0��63O[�����������f`٥П��@��c�[�C�@rD����uy���=�/��g����%���T�q��	t�b$#%;m�f��p��rm���ĸ����,홊>��2�VI�k�1��.�mr�3` a8��14�	�ݺO��H��s�
U�&��+��xz�s�=��0hЎ�S5���H@,�3:����de�C���}â�h��R=��v�t2��ݽ�~�p���~�J��7���9@�N/GK^HpQ��g*Ռ�{O���ǟN���P�_S��˲���\����F`�7�� 2�0�r���!�Й͝�s`:�9�O.�9E�錐�34� �� F<��7�(X��"�\��hI�� �-<[P�Ģ]c	��R���"B}�r!���2�	��*M�*@&ΐ���a����{�BQg[N<Җ��Û�A�5�6(���b[J�~�mܵ�*�+����7�f�'laШG�ץn@
���p��"��M����}/�W��3D�`��5��C�^z��á$��\r��ON!���7�\Ud��=�W!I�;�}�V��ۢ8Ӎ�Gv���z���z�R�
י
 z��1^��C�՝{E���.@�׺j������E�8%oŕ��o�隳̹�(t� 'V|jP���R��Rx��j�cq��*��m��1��߯-�2&:��V�D������|@�\��I��}�HOg/g5�nA�W��!}!e�c�:+���n��U@ ��UOZɘ�e��7ޝih����/55���g�g��.����JZ�λ3ʯ�;�����E"Sݔm��-�t�8v��M�s����]��NW��|��^Ubt)S/V��B�A��r6 �h�{��N�h６��3�Z�p�m��dW{G�c�%�*�FL��� ә��:������.�J(K����5���}%�22[�EH@��k�(a�K-Q3B��I�F���$�(v��]��T����������܌��!��� ���\i?~��WQ-	a퉨�&Ҭm=��� 2��6�J�[���bη���ehoq�V��t�o&�����3�����O]����]Koгo$M��Y2�=��9{�]y�!�� �^��)xk��4h����N��B�!^�����a2�Ë��p�U
��*��iԥf�*C{7�.����b�s��7�h�[]�)u�����ykis+@������1B�~Φ��:�h�~Y(�;�g���6��H֢-�r��I+��io� �W��8j�����B?x/�cO�'WA�̂~�����jw���O�0@��Z[�&�!����-LI��v�[5B��S�v�ho)L�D�%�W��<������lOy��Z���%��]U*'G�q�"��Tz���؅q���Sv�i"2�3 M-�n�:��/oQ�.����j/�Ҙ�P��"/��|��>�M@��"�>�%+wDK�@�σ�-6�Ԕ[�y�mV���]���QX
�����T�>�|A��T1�Ğ��uOd.��o�m������A�a���*��[��_�)����j:��2��O�X��i�:~-Z{��\�ĿO<[E�P�v�r�6r/��ըU�T8�d��~T=�^�;�2b�ƹcuRy��� �ET�V��]�h������$t�0$\i�V��k��q�����%��U���2�`�;0M���|�wn������׎0���z��� N��j�̰�Ua��c8$/nyV�� ?迩����<��t���`�M�tv���0뛻ވ�X�x��x��+X�-����:�S��H����?rS��)�+�ՍY�>�W=FNܞV5���݆<��nX��Z\���Bѿ-��L`ILtUzk���x��9<�G�� |kA���Y�[�	`t��q�.����t�3�?��2�7�g�Z�R��o���%���@W��(�@쎞��H�F�R�σ���YO��L�O�K*l��e�Z�b��	�#��X.��Y	!a8�+���+1�Gm�C�̈́�;��F$�}��Kq�@u|�hTf/Pg\z st��M�ӧ�dQ��ݷ��w�	���9�@!��C�X���pT�s��F� j�Z���:Q�W�8�v�w1�m�"m9=�}�m���>e=C&�������~Ą���✥��E�5+Ӎ�ޠ�2s����6k��G.����81�ߊ]Z��2��W�	1��m�y���i�%]��2����m~!G�
;�X(6�Be	uox�_�Ґ��h��Y��e���u)QHfh3�.��)��j�7�5E�&=8����� ���i�t���~N�'<�G�}��09�I��������y���)�QH�}6�XO�VgC�z˘W�%�܂=4��L�Zך�0ܵ1iY���ތK<~�q��[(�>��ӊ2�\���äRn�,|��>���-���8�W Y���QZ x�����W��.�Ԋ��voL�C��jW� *P���K:�*kP������»���k=�"�ʦ�����
�S�m,V����ڝ�7e_�,gU�H��6��T^��kp{����NV#��9	�^�1�Њ2)�A���u�<���W���^
&��4����{���:��m��mtd~�+�:#�Z6h���ZS>��٩����y�z܇`o����i��%>#3����XJ^=M�&Va�+����ۼ�Q����2x��� �O�[�k�Y�����v����KX҈:�����I)�L7�z��;щ �*r�2.��`�*�H�]�v�GKW+�&����=���s�I��_&+��+2�Ë�����o|u�X+`s����_��4���/y�����xV濬je���2���ˍ2OK�G��1$ʈ�ҥW�m�ͲYt;0'x��d�Uc�?�`�CVl��C3X<��bs!W�O>�*?��k�X6��Q<�f$�O?�	�wR�؎�'X���qy�'�����8ԯUG+Aۈ�<wH@8��&��ֺQ�����=�f�~q
z&,/P韮���{u/Ӷ�K����f��zƐ�� ��Uhy�W9<#�cl�z���~���@I|�3�G,�j��!�b�Mj<._q#&3"щ�0I�ڦ1����Β�( �[��Ԭ��&�:���^��F���Lȯy���9>嗠,��-�Lr@6�c���-A�;�����ﮆZS,�9��{�ޞ`FD�ɉ�	�I�]p�EK#�.�Bؼ�}�� a-W��JA���K!��f�I�t�z�Q�A��T�re�)3{іvM��?,&��I��лH����"��J��Q"Ae���m��!9Ӯ�j�4�Ib6}�	Sg�
���� ���0�����평@�|��'�����G��������U���� �j�?p��u"9Ȑ���f��߅�b5K��K�r9�wA��/Q�WA��I0%Í����H����K���9�:�@wD�S
�U*��(�\X�����.��� ܇�y���*���������V]����N���~PG�E�#�C
Ѹ�+.[Q?��4������j�5�qr���> �Ĩ\w��]M���4c��Y�,���3�bh]��j��9/�L�
 YӃ��HV�Ӗ���j���3d*f^��]�B_t�oNX��5T�Qv��g
������ZN&����+X)kW���Q�*��x�],
�XA�1pb��U�<���	��v5;�