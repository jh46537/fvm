��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����i��;ݏ+��ↂ0�?�ceR
k�&��;T/�h��HKIw�|��&3.��Ů��p�!Q���i(�+��gX]����\G��/"�TDV
x; ��*���1$���'�os�G́�C2�:>�r��]�#A��]F�~?:6�,Ӱ������4;Y-�����|��U]�Ԝ���6&F,O���*Tkt�Zzڠ6]�ޢ5m�IS��Z䝤����VX��@)���t�I��Ml�k�{F^��-���2#��q릍@�BF(S��:�����jm�â.]"�	�i�,��Z��GU�՗��5�P�N���Lh�����	"���>�֞=]Kd����;�'��D�Yj���I��Kv���R�]���}
�jD�Kh-��W��M�� 	����eD��p���.��8�O���lD�Wa2]8)�b�;p![��5E���I6�����>FN�,5��y��zo�����f�_p)���P�Ey������0~$��^F<)أl�Ϥ��uvLi�9���~�B�pQ��9��>�_��/�:��H��R��G�MZ޳�h�i��Nt���4
F��2�T��ƣ��7nݨP�,�Zh�T���i�
����b�~
�`��+����e��
j"`5e����}���<%��H���h�8ו��:���w��(��ᤃ���Ԗ���;x��K]� ;�L��~j���g^��j2e�h�+Wb�0�KH1��[!����u�A�b0U�ԵJ��X�gi�&t�6�K=�p/h���}���˷��S~�q�ѻ_��@��C���M��`_���f454BR�����JLM��t��� ���u��=�V��θJ��8�پ*~�WD��nI���2��v�����E���Ë$�o�������e>>+��{��KU�lhe)��M)��Z2��k�z0WS��������T�R`|X�M'��jYh���_�a�;B@J`EgƑL�sdMsˈ�Mn,� �/i]�K��41v\yD;��P��M.�J�'�9��{��K���>�1����Ձ�N�m+��$G���E)���dphFS���	g	�K�O��YO��|gx�$tGd�c ?�M��3S1,L���"�C��PBW\���`N��St;Öpq��m�*5p\�#�v+�4�'�V�ʣ�,L�졤�xyZC^��L��
Ǐ����̈́xp��yxw~�s�8�h�qK�N�yRXtm)]�9�?��nS�v��F��^竔H��Rx�H�}҈y$��B��bf��?�N�($p9��^r��2�d�|��M�!��E�CLQ���Hf=Z��r�����c��T�9�0�	[��Y$6x7�	^3�6�0e��?Ji�1<.�*�0�q���f�O��͟�5��O0|�Wٲ��@#�6j K*���"�Fx;[���#PFc�G��}�/?�St�Q����Q�1�2�B1��<,�q��^�F�����U��g������yѺò���s�C��+Ƥ`�;E�Hq��"+*��P��g"Dv[�p�H�u�u0�ߍV�OZ�_ƄѤ�L0d�?�x;հ�m�`A*�7�Q�@��z�KM�*c��ؒ��ؒ���_�`d �v��,��-Z�jGN�
�PiH�/'�ݏ��g�%~ob_�U�Cd���yt����H�ଽ�����?ں*��u4�'�(��7�?�������Źz��Z�Պ�E� �1�yn�:�ax���0��4�U}хD*����m#��
T���/�Xry���-'k�_M>C
�åI>w�F=zȖw}'Ab!�#)���ic |����k6
T=�lh0�_�MB��Id̙k��`r�N�Xaxi8��M����;���(Ht�'�}���+w#�h\�9�1����s�F����EZ48WF��1{,"� ��#�L���X�'MJ��j;��ZZ@��8�Z+����[s�J��7iX@ќcUJ,	��"Z*&4����R^g�*�Qr1�@u�A�w����J��n&i��Ǉ�$������������Ln��d���f�S�S�H��/R�4΢l-�0�_�<�(�������C�"�6l#�
������þ���E��F\�W�F���Q�|!�yn�;��NC��i���Y�VH/u�q�S�J�hPi�T
:��w�n\����~�Х�֝�4�A=�tZ,��
�a�ȩu�Q�|>�|���G��b5�<�B�.����:#�Xehd�������dB�@�� �L�m�߮�uU]�|sd��Q�a�ꬨ��/</�TM��F<��'��ʰD�p��ڇ�Y��*T�-�|= ��o��4E�����u�Q���AC޷7�Q;H1���rj�	tEta���]�U��༽�e�yK\��Y�?<0��F-_�n3����w�����7�3�Xȗd�9�ylX[*aIx�۫�	��8����Ur�̙�Q�!y%���pj_�����ӡi�.3��E�k�L7g��n��z�N���) �g��}ʆ&p*�oU�|GP8�:m�>�>��Z�V�3��d`��kQ՞;�&�vU9�3V�T����3/������Ac�\#�7B�M���x2�ԡ��v�o�ddU�>��r��4q
W�~�A��� ��2F���!W�B�1��^P������|��Y�DY�]چ��\�%���w`  H�oT/W�32�ӆ��T߅����2՚E��^
x�v��{b۲�7���򍞧}���O���5��e����lk�}�
Â�i$z�|έ��Z�K+���V��X�'m�p?G��W��M�Y���0�WQo��'��?��ox�c�P��KCo}�f0=��,"�>�e2�(�bW�C��fhO��� K�v�އ��X�D�ż�� �$,���i;V�r%��_]UC��n��r�0|�<*�]
��킓D���
�JE��J�h%p� ���3󢨮:Ć1���]*V`���[�����-�� ����ad���" Q^��t�p��,l7|M�A��@��aB�~�}���l�q�q���d���Jz��Q�=R��U���E��}�s�Qp;�V �n�Ip��B���O�60F���Zjy�i$�^�x�L��M�Q����e0a�]6��ƿ����d:2�=S٬��L_����`�����-�&�e���
����k��>��o���h�5,Mf=���8�I��u�K2{%��6��ӱ�L��[[�إr,�p��K�+_�JV�9�W�� Z5u�����E���g�,f	�����dd���ף��1��,�g�Z ���@�$h= (ŏ����v�hq��c���� �{���ocݷ,�]c ��	g�v��L3�ٞ�{�h�~a���m���X8�:��K=\\��I�G2��f�m�6�![c��d�ԛ���jq3��k�ˀ�h�w��%�[K:>���e�Nfe���1v�X�s��d�L�U�a�z�a��ݒ�V���"��
k�!�N	��"8�~�Uv�yOs"!�챬yd��0��e�o�?K�Γ�T�6��-��+`�<,A�nW=���U�Q"k/21Ta�	y\��WK�W?���M=�"J�ZèWS����u����k覎fes9��V{��N�������Ÿ�����?��� ���!Z��#ϒ�Ϥ���m�&�Rz�t�cn!�EG�^��DN?g���#h���̹& �_R*�۶�j*LT�0f���d&�J���7s�Df�r��]��bn����	t�E������8���`��V� ����`���M;-Ö���&|������A}�W?������y���N���7��4��}��%��D�4
�����3�r�����t�Ԩ�Jpz,�� $ْ�⬅�>�Fs����C��w}`�����"H}�*���?�ů�Y�rL�e�]���r� �M��d�P��X�-x��3Râ7,�V����)ruil��S�q��x����a��ׇ�ʭ��f���'���F:�-��(%�o��0q
�)����,<uC��|�n��G8�E��FfK_A��ਇ�(kOq�L�[��ĩ�j�6)��ֿ���kCqVxtӂ���� j�5=��9���bA	�x����CØ�K���R��3���}}����p}�o�ފT�B'���)>5K�kSR�f�b5��&K�8�H���&îo�%������dN*K9��u�
$���;�ޚe2|2��{��6HV�1���GNkGh���	Y���Q<�j�r���*EW�.-�����뗪����KOv��ʵ�&!��6�:�
����YKc�)�}ͺ����_/[��{6<~�='龄!�t㒝)/e��߷3	���5� ��J�ݒwk��(��w �[4�1ք&`��e�/I�Q�Nr,fP����������� ���Sl���R�p����<����o�����-qU	�&�M�V��f����+D����$|( r�21�JDq
����$�E�d�?˷l���B����|UI�����$w;w���{�G��=T��������*b*��u��L�9+0�^�dE����A�q2Vlz���%_�2��^b�0~�R��F!��n`p�H+�!3��]�qn�`����M�6��R�U��crI�LFYw�y�\���ah���L<�����А_����"vl dOq�]��iI^�?�m2*�G���m:�zV�п�Lf-������[���q���\��WK�J�٤c��|����0��5�͋���q�<7=^��)Z=�uL�D�:�M�h�q^c1�!b����1$���1D�/ ���.h�F�A|#�XU��MԸo��P��q���5�ɠݠc��� �h�3����#f�g"�t�����ۆ�$	�k��gPR��[T
��K�}߄�Rg����0VOF?n���|���?��+b�m�~�+�T%.�E�R�T��q����cÒ���v�M�j�H}V?kO���C��.��	���q�;�D�ŢeSl�k�~��cnaV�������_^�(��4�u�Z��d-�hi{�n��Ryof����g�S���7�#%�*{�~tmw����b)�Yl�6E��4���!H�ʍ$��rg�5��H��U���-�ꈝ80L|��;;�g�YKg�A�)A5����Wj^��_��q��U�V~�@&�Y����=8��m��������H�h'���m��z���V����&9T��-En6yq� *���B� &S�� �V!a��xp:� �qg����7Y��_���G_|i�}2��V�G�|z�늑��meW���X�F�O8��	(5v��vƑz��\��=V�*<`!��r-�D��L���f��Q�72c�ݓ�8�mp��HeUO8��1<����H�96�~,�=f��ps�~"c��$5�`a݋LV�W����|Gt��`�\��w�i_2W){��C�!��������N<0A�� w{��E?6Kƣ@k��������M
J����|4=d�h��WH�WC��i�_}@��3{��	����D���zLd�ދ�Y]]V�m1*9kF��JCn��|�߾)�R��1]�u[�/^��Ԃ��2�w��T��9�=B�!�T��X��`��C�̕�F(TXҌAԘ�<��n�]�3��Mr����(]/�'��o"�{_��l���҇o���(�8u`��)ʖ��<�ޣ��~�SjkZu6]��#n~�mP?��\��0�'X�t3�f�P�#e���:c|r��!갨�&	�_�78���J�IBJ�S
q����� �j�稸k<U�{�ܡ��7+m�1� 5~l�+�ƙʃQ�b|(�����[���k�IƎ ��w�w�B,�]d�\�5D"2�,�M�3��'�4(;��0c��TEYvl0�~z��Ϥ�LX&]1 �����t��>�7r�vT��������}~�
�e��u�v�	������4���5L�ݾ��:;��֏1K���PM��ˊ�d�J������7��D���;m�ccI�^a� ��P�o�NtЇFb�e��8q]��Fd���p.�@rS9�*�J�~OӬ$��X�W�#����r�,�7��m�upX�C�g�$�� g%�K�a�1 =J��%dq\k��H�sA��xtE3æ�us�M�B���#�4�M%r1�Lh�M���:�"��ՠ���=W�Bp����:������1|�W�k�K P���GN{1����o�.��ak&0����N�*c��
�*}�!����O����"�>��]���M)PU�t	ރGf�Z����;W�D�Јvr�̮ɛ�&��:��	��G,�+R�m*q���53ɕ��Ŝ6�}	l���aM� |ݔVn������8�Dv��6yfΕ)P���{��n�%�%��8��;�g#.�bގ���{��z�]�j��_:$�]�3L��K�!
Sa*��b�z���F3�!�+LpRq�������ĩ'63��~Ip1#�{�� �Ԥ��F+2:�^��[�̹�骞J�]Ԡ��A�&%?�oj!�Do�	%���|b�@�#V�6�����G <W�?ދlPU_d��BaO&Q;�W依ʈZ���d��<43A*��ç�y$Gӯ��on�
υW�M���Ä]7 �@[em|W��E=�/�KtA�(�q T������C.k ����n���|C�Js�� �a]����X��:�C�6�X̰�V�_��"�_Fe��~ނ�3�Uh�̟d쌞_�#`Z�M{�>:��i��wdu?.rֻenL�:�rk{�|���Q�Q2���Q�vN6�,��u�S�0����� ����8��{�����y��g'G�\��)�ta@��!��6A:��i�m!Xɠ��F?GW��G%�k�a}WJ4���
_h�n%�'�W�@*)&m��5�6>p���M�H�Q�cQb>�j!���O�2D]��ơ��<{2���2�<x�8����L�M�uW�w9� L>�0� շrg��2�=��D	��#��I��7�]j�[ �y��17R��m��:T��PSv���khF1K����&���*2�����q(��<��D�+���E3҉��34]��5f�׌^bu��ȧ���xV��j0��r�K$&�n�6]f֚���E���g�\��(�N��I��[��veZGb�G��쥲� ��ق�d�\cΘ\��/k�LJ�*�J�G�`SRvF2�=o7�:���ܛTe�^M�)��M ���T�����(���(��J��Q7���^Ԣ	���1���䈀��u���W�W���	]�axArk�MSbc��ST�^��`S����a.(a��n��d��_2�Em�*z�Qx�>���j�:*���N���xJO�jV�e��7�Z<��Պ0�+LB�x�$#�b�V:"���	j��8l��gl\�)T�E��R��U�}k� �Dg��`f.o�tBAԵ>�_â�p
&%}3�Z5�l��ËEy�$!��-�+Fc%�l:XER�({� ;�C+���.�+��[��9}��@���
�^v	���Z-�t���|܏-�L7���ĥm��un{��Nd2�ܦx����]�jߢ����a<F���"�����4���D�����X�?a�QvG��w��aN����1�Ɠ@ż?]�gt�&�;�ܧ��i��6� oc:�'��Y��>�`�m�ݖ�_Hz��������3:v��|1�[������e<#���B��H��9����?��${�eonH�z�!!��w�%��R��'\a�϶���کn���d�9M�o'��1��:�bm<z���Mt���fwC-�@��o\<�x�!��%<��&��<�G��5z�I^XP�~V��b�{�D�ÉB����xI�Jcȼ��-P�K�gZ��n-����21�vVF�!��ed�+�k�wM�O�r�ۻ)NLJ��^f�$��pjn�;�!�G..Gl�"�)*�U#���o�(���M�YD?ֱw?U1L�;t��A<�=-H�d�7I�ւ0��SS�?�/gO�N�)�1�	2}k�=e
)@���ղ_�z.�c�Q�l�O��0�K#2N�0f���7/��Y���f7b&,"20�'�g�����e�ږ�q�򹑬�fYdL��<�v��/��ϭ�w[H�=~ �@��~�`_��
���d�;����:�����E�u䆥Cw�u/�;�P�P�Ɉ�vB������egg.OE���j�2���|J~����*�ݓ�^�� L�����$=JJ�F�4b4m3$���O	.i���6��n�"{a%�Qm�9O^�$��
eo.�T�CRt�N�
����l�d^Jm)=S6p /9�.��`!9(T�1h��<��2�:��~^K���I&麬t�qT��j�`$C׫�hf��)��a
5+o�cЎe��
Zj�wq�ߏ�"i��cLj��U���lזa���N�&R����[���B�C�ſW�:��g�F�>z�ӁgX�i�N�u�R�IOF(3��1c��7w�/?�=�ՌOq�Aj�g�#8y�Zfi�,�����"xB�O����R���5��1����T�{�Z)ѡ[&�ᐘ��`�5ߋ\l�r��>4n)�;�rXRÍ�}�L�@���";� ����"� �B�L���Gm�-lGҀ�	�'��Q�i�xu���$9;��^����-�{�"2��D��3 i<o�氚j	��d��[T�J�*��Y�Rm@�Xy K{����.0�q��G}\�B,�����n��&&5h\�O�e��_�Ə��ٛ0�z�ch�5�-?d�Y��P����_r�=ꩈ`2ݓc�G@�9 �K�(l�c��k*�&�"U�x�&x����؞�ܯ�����!{"�x@�o�w� �r�˩� \�� �P��"�^M˵l�;	�;�����M�\�	;U��8�N��m��2O�lD���� ��5<���e���.�s��h�YV�(S�*Ѣ���L���8����q��%���)ʬ��#W]U�*�� [R�ָ�f��,���A�R�>mHt�*�)#��}qKZ�v�t̓HC����3��C컈�nѵc̆u���MK
��9�Ԉ�� ���[�Ȏb��1{�.*�4��[�y0��hq��(E')mYb3@�̓z0[�t�A2,���mL���>>���_����Iva"o0�]J˩hj���=��o1����pw�y۬Àr�ؚ�~P�������x����Oź�+}����&�����&4 q���sj�_rg�'�i���\�
VEr1{?(r��
 ��r�e���15l풒�R*���i�#�|�o�A��2%��=e/�a2uȌ��,����K�%;�f䨓kY�Hx�������hW�:����*Εu�q���R���D�O&�`��n�Cy&�`�X�uO�Ld� �e��r�P't;	�"M�d<�eڼq�@:����((��R�6油w2��7qn�גF�*��z@��I��5A)��儀���cj�r)��>ǙB�F�m�����c�7;�;y��C��D��ר�?6�_U��R�U��o�my�R�!MO��-��K�t�g`I�D�N6�u�T��y(�����1�~J��t���UU�q�t���b�	����M�]1�{��7�t�J�;���:s�\ݹJ�Vͤg�>ɦ��O?�(NK����z�
 n�#���X@����N(!c���F+:)�����0�EV��*�4
�����.��#�ǫ�h��0F�g*Õ�y�����9��[?�L��EY���7����Z�hL�27�P�f�d��mB���Mj�@�Q�02ܒ9�s;h�ߌ�ΖRJ�6�z�I��_�Er���(��z;��3�Hc��2!b�o������S(0��)���k���E�+N5��4)�W��\����^��8��ޞ{>F�غ�+�!(��,���%�~�D"�y�~ob��]��g��L��L:���ה�A�#�m��]�?��$f�LЇ�OË�C0���i�g$p(���G�HH_�8L�����^��#����q������2�?��$��uAf[��G*+�yP{����D�ή7ݼYma̥;l��	��1y���yFTn�ϧ����޺7���G�Ѻ�\�p|3�g�����B��vB�����^���#��a�-�%�ށ@B��$3��%5I��@�
���A/c�\�m��k��yC��B����)x�j�f+�ꀈ[���xaq��/�^C�!;��'<$�ѱr[1I1��Jc�]y�?��������ɱ�������x"i���>��}�n肭�2p
<$�D�5������f��q�,��*�EV���^/�n)//6���.������ 9�	�iX,��P
��;����S-�̭��IU�,��P�Wp8�/ԝ�\�����7����E<�U�N�&H��d�c] ���E�;�K�hf=�6q���?�A�>��+��m�`P���q.��Q�l��FoܨT o����6��Gk�� D�Ȱ����]F<������u���Ó�&7g� I��g����x�a S�Ch�c�Q�+��0�LMO]9���C���ga	�D�`�#K>#f�N��sW�	a]��Uڥd,��e��c�đM���<j��6���jٷ�{1JC�*K�>�zf���^�6ͽ�2[փ����Kz��Z��ſ\��r�-C�,ܛ�_,!�1��_����Tia(��f�����F�ӵ�#:DQa�����7�}VA��U�ٕh�
y�������\ �F�v�k1�d8�"j�d����E���Q\��Y2}[�m�a@��t{��Ӑ��C$�$]�c.���d|���{X�Yѱ�.���ba�^?���`��a���z��_���ė�ఴoK�g�5��[[�����H�^!���*2|pJ�f)��X0�����}�\ ��<
���a�Hs�j�
�'˹Z��z�X��ρ��Z��$���_~C��н��C)��L%�ڛ�L��)�������f7W��>
�Sg�%�0F�<�L�uR���P�#�J��g�J�YϷ9����Q�ߌ}����9;�f��� &n%gcZK3ґz����F�S���qק4�{]��'�C)�Մ��
� �ɚ��4iߐ!�VY���9fd���Eӝ�aż����vSr����W�F�/�z��R��p[�9U8�q�7 [ Cw�r=&��⎈;�m;�����k���t\h����*��M�W� ��;��p1��F�#=���})=�[�N#�=��Բ��~��������~g��IC�( �&u5�Z�E����+��	�|��0�O���_�g �l�U���:�hf�w��}"��S�Xc�p�Y\��T�+���b���V���5���Q�x�W��,�,m6F���K�����ɢ}jr��*������G��åF�#Y�7���E�?]����E��`x +G����M�Ec�y%jg��i9�VP��av��]TT�x�ioࠜ0Y���;�(���yJ5�kNKΡ6���KrVo��:(jx�f��;�#LSz~r�o\�� �;{m������B��i�q�W;��������n��m;yW������E�iĸ!��z�1�����6��.�fw�T��"�8�+��)\J����>�2���!�d��^^Q���\Ѣ��:6ۭ��]u��(����<���S���n�柣��}?�6G��z�%����7��2���Ltb���2	q0HK�#��A�>��y����sR�_��P��1�@n��(OS6Dț��E���%���H��|R(��-7�2�5��I����(0���]�$q�i� J}���(v�F�%p�٬��f�����xu��s��WX� �΃]���9�����+Ã�Մ$6y���
�s4���	~���g)��.����cC�uzPmG��4�WN׈6FOM�;-W����v��$;/���w_#���;5��:7� )�WH�FK��ч��x�ĭ�/h�<����A>z��Oɏ"��m�rls��Q
�Y�����h�*d~ �A��!z�)��i���}$|�-��.��M�� с����t#��c^[�z� A�~��(%�9%I�C8 oT5_��ٻy�6�hO�ĪX����0-F�)�ol���3ª��R�,s��rtTa�S~,+��9��TY���w�Q֨�;�8ɩ��"l=��%��O)W�Lm�MP·�9�+�>洷��5%�\` �$�Ԃ���R���N���e�8mv��R �D�90�[�Y���<�r�~l��S���~ЂNH?|Lh�k�(,_Ka�lx�Vf�u�]�
#�yr.7@`��='j������D��$���;���!�a���+���:9f�@��c��^E-I�o���g��7c��2�7]�feˇ��v��qퟎL�y�`�,�W|�=Qͫ�
@2IÚ1��knwȪ�l������� h��5J��O�4x�h����:�0L���-���b��lY|�sB��0@ih���#��\aw��2y�?�Vg,�Hr�^�>�M�G��<}��7��2`��<35s�cH���0�a����a��X�/N������c�AJ�6�*=��އ���1���a�zgI]0X�OÞm��ux�+ �W�Y�X����ppb��ʫ����G���Ʌ�xTf�q5b"�P� �W�<�f�йLE��QP1�a�I�ě���:��)��|Y��� �mҰ8�D��GI7��`l�	��yZȘ�W�(��G�/�	ړ?��_���
�W����)�GbF��O	����
�$ʰS� �����m���(f�t~B�����eQ�gs�m#�d������� �h�g��r��$KQ������'��^C��.���۽󣘵,�0�㵖��b9�#�H�
��� J
Ѵ���_պ7�&!�.�	�� ����V޲���DDU��X`�� �����4[]�'�L����Bd$��	���4�r2A����"K
#���k��6�Tp?�L�|Q�.�ɲ�-Vږ&'�>$��D���9�z���Ds*�t<��ƕ�b�Ë������<\��3�7J4 ZO!w.�������z�V/8��(A�y�u,^�<�ե�6l��[By`}J��ڸ��'�ܘ5�o}c�'�s���[�?����D��$
�5������ �:a�4��	��sp&-K�mHKfE��&�g��;,jF�V��@Q���*�ƞsO�YZ-s<�U?��t`@Ӛ�d���S���6�8������΅*d$0p�[)9L�pQk��N�]�5�Ȱ���b����M[�<��ъ6�h����vɰE����
X�ى����+y���`�>�Z_1/,Ϡ�;��?��XQ@����\�O,��}.��=y7\����@�x�C���|�����$I��OF}LO�Ǆ�d 2��A�Ҵ�;u�܋l�%�$Ƞ�����Y���}=<w?k7S��x�����s7&�?1Z�	����rS9��6�Y���{ģu[31�����H��B���:
!��E����ޝ�&h���[�,q2���Y����^�;�쮩IZ��F��j�C�z{�bHo'd!�q{�ej��V��F��%�=���*�왣����^͛q�b�Q�t8*o�F�1�l~z�x�N�3�.���� ���3ǒ��<�$�z�>YC0z��x��h5�����8ZT��/K\��uo*r;D��񷨠f��Р�J�a��U{�5A�� s� #�|@`����팇.z���?����P캙;����1ߚ���@Z"s3.�h�/�Yl��É�{�j�r��?���roK��	Ey*`�K����+��/"���Ǯ9^�<��&/�{-M;��7����|�Jv���:��H����XD����ͪ�EZ�/�p�Ik+3�ѦXh�-jt�3~c�0!�MɘL�c���2��=i l+������z1:Q3?�ۯ��I�Ԅ:T/�+��^=����g�#�J	����Kȡ�aB���M�ߗ	�O�W��-.$���*rG�J�Ɛ���_g"1I��ai��;GnK�Z�a\�P�M��L�D�|
����"�2a�!� A���$���{��T�V�h����wo�16�.P�soC3-���.�Y,�JI��+x�	
6}^}�9Ww��X%-�N�r��ȱ�'k!>������B���FPބ�Pi�4�`;�����3�G��v�	�vH�����N��`iqR�eI�!*���)�<B_@_�O{��`��V���� �{�
�:��v	S�j�&NUP�Ș���� �:^���r��s���]p����Z�pUMWŃ��Ȫ��X��bֱ�"$9!8�'B�_n��I� =-�����Q+��1�<,{���O~n�Y��������wV�ɶ7�Ҧ�	f�3`V���2U�>�`+�b
An#�vtʤ3l:0�o��;]|E��П�O�I�ꜤBÁ[��������dF�G,���YF�GA'���^��n�S������
��ޣ�(S�/��������E�`oՄ}�
�a�e�uVee���\��>��S/�\���N��gT"M�chv��V�[��l������L�99檣2���C*g�mR��y�����M�?̴X��v�0����lИ�੐��</�N���(�<���D��T�Ԍ��0y� d����xU(5\4%r�n	_i���޺�6<X�@(wp���ѧU
k�1~<W�`k�3��o���m���?�7Y���nlB]]E�=2�_��n�7$�n���*]�^��1�hy�]w6~�uB�	�U��[�`�~�iݨ���E�Zl�ΑWز*eDvr\J?�����W�c��"�(�P���ݴ�V���%Xl'?��U=�[F25x�^�J�~�Z#���OТ���I�gL��O�E+�z~d��(i�����!~���)W� ���E�2�-�����>%���ú���d�����JS���X���j�I���*�[�h�㻙�8�P������A��d\���O�Ą$��p]�x%� :`7�7��̅����dd��P
��#�c24V,�u�s�7�*�r��[��[�M�[���Q	�	J�t���3�,��př�`�]&��@؝��̨=�Rf������:>x�k9���PS���Ԟ���{+Y�q�o���7#�`~����3K��Z>���c0�t&���hO�oM��I�\k����N	<��S�(a���E���9`��O�A�C8B/Y��LYf�F �Ŷ;��C&���E��h�#*��.�ÌB#�>����ED�ן*,�&Nɮ��l}���4  qķ���1?�r��-*�)�9Y �N�m�k�Щȸj�oH��7��#6 8`><$��qDc����iq����\=�E҆�	sm��d�|��u;"��P�5���PiS�I�}qGUe�I?B/M3��M���U��4m�ʄ�M�JgAy�j��lTٕ1��x�g�^�����IU����v���_<)���N����`�9�U��$����J�Vl���=ڹ����������
�`Bv\W�w\V�Ǉ�+���%��� �L��ީ��� ��7��|ס�&c �z�>�8��ekM�L����	��Nյ_Pi�A/�zG��jb^�h������99�����~3/L4/vx�4�7��H����@���f�O�G𹚄Tbs��W�(��>���|-�Y�e=/�6�΅V$e�+eww��Y4y�^���1���"����qj#����L��APu�k�E��!ٟ|������1��z�Wt�d�����A�{O~˼:j!�Ý�_�V�R1��Ц$�7m�n���P�X6?r~�q���Pǋ?F��6��9���[
����]>���N[Z!�� sL@������M#�_6�b�����,����B���mT�}W\�^�:PM;A�� Jm8��Ȇ�������B-4��
\e�x�D�WG���W�σg��72>˰)4���nD!����4��=����-��g&��� ��#�+��o��R���h٣<�Lu��!�Y���y�]��ҏ*�PKz0<�|jE���+���׎D���#�Ǟ���(�	��\]6��/9��l��kPo?�����5����T($el�"��ޖ���T���� �
V~6y%�6�m�NJfN��6�� �ȐaT�Ař�V^L��>0\�:��um(ҜL�Zd��ۇ��m�T"�Y'a;7���(5��Y�E�>��SE�]�s_/����t�8�>�h^g����7((	G��x_��]b(s�_�P��#(
��|�#0�9����9	�~J���7�	��8Օ��*`�T��9���<�u}����Ǩg��V���W�0§˷EoA���:�$��������*��J�wM�V�Zz����Z֝�?42�`�_�㐕i
�ߛ��"����'�D��Մo���2���w����ӵ_kS|݌�PS���S[[�����-f�:<';;����rx�����[�v��<�-����,~�@��{Q����1|�����!2�^�-L��V��]�3k�DXmWw�g}j��B�^U�8h?bh|��U:��N��\8��h�� �ۆ=׭�@�hh��g���eԛ���P�Q���m�9Gp(_,��\y6k��>/Y��[y��B���3���5��h�琐w[��h�RO����+ʦ�+Cua}9�|�l�)P�iEIet�����G)���V�&��9>z�W��-d���h4B`	@�)|W߉Xi��A>U��<|fd_G��+���+�U�b16טQ�=t�\&����8��$��s���NX*WǼ����H����6���)�h}|J��ϑ��=�$N��y�ј�	R% �u���uC�5V�{����*)����k�YYv�������P��Z'g��qL�tLjD�aD}c��90�x�u�m�Z���x���I��{n�L��fm#`�{�k�E��P-b7t�����\�q����5�LUn{���Q�n��*-.
���o����e�x�j��Ԫ(jz���ϗX�S.�M�&��2�����i��1s-[��3��SC��)���)��}�cڑX+/�Y��ˬh<��Gvk����v�l�Nfi	����Bg|J�KT��Z`D3��i#�W<�W�(�X?V�-�ts��~!�-�~y�G�t���x���2i�m�(��97����.�<��\z�Ԏ.�닪2��^GE����`��Ħ'�h͔�����,6E� �<�􁔟-AF�(3?�����0E[�� ��E��(�j����x����i���FNh��&���@���r�B!�)WHL�ﳷ�e�dks<��E����`|�6�;����`�l�������Z!1�ߥ:B0=GEX��w�?���K[�`xZ�W���&�A�,�qh@U�
#Km�^�AA�b�Y�&�
�3f��_������Pk�̑x��놙��'������_���I�y�Ӱ,��+�:නL�읝��^-J������02Ó�=��"�p�Un����SzZ��2Z��4���-��t���6b	?�i+��Ԫ$��N
Sx0��t��M��;�i/�¬�Ʃ�5hq�Gx�0�ݤ9��s�Ui��[!��z�j�Y��\��@�XW|�$UF����&�����zN��㡷t���3Y;�c�:g\�9��T궓Irݰi�+,\Qn����F�rg��Q;�����䤤5�wM��N��"�.3�q4�Y��
Z)�g�1�zk�s����C4mj`��"��}y�q>�����U�@��{�e�<��?�B�W��X����Ӵj�'�_o�{�{�X�s+��u��WO���^�Ef0���Ť�(�I�).�<ŷn���X�x�om(�f�����98O���D�7i��eå�<}���4�P�E:W,ا�>�{*��Qy? �~H��<5�%�1������s�M�.K��&��G�I�/�w���D��@R��O-�O)��"²��0���l��]:�}�H �����sƔ\lY��v�t;��y���JQ?fni�u3?�@cL�$UA3i�St���U倕�H/�F43Oy�	l)�n�"����tn����h
<�5�C�'�ٍcl���L�����"�X�|>��X�"ȓ��߳���z�*�Q+��s��g�w1�b@l���=qg=CW�^<Fꆇ6@�bM�Ԩ��R�&6��c37\�5�uk@���J���4�oZ7V!����ɰ��+V�i*�"Q���i?�&�Qq��D�a��,����ju1O��;U"�����B���F�Ҹ�q�i�C��4�;G���lrڹ��.E.�|��B�r���+H}�2�
�	ttp�vbA/�����	�#}��W��s��{�3��tI�ʣ��7��>�i�����g̷Y�*HDL�~�r�V9�����YG���݃`��������1G`����!Y�w+?]e���|��ԗ�������i\1j��}��c�I������]��6�`\�����%�}{�Ⱦ)�LMkC(^��E��מ��܈�E>��&8��fa嵯�=	�+`(7�DG�
�I8��$˅ڻA&�9��˔��&o��f�K�ZI5ĥ��|p<r�Rp$W�M�����=�4��_�p�[	��X[��2�p����@�R�����,ӿ��n�uSIMJ,`��Xlj���N(D@c�@� x����ݢ�iь�j�5i~2
qpyE���^�~�G*���S�n�����:�%����Ԇ��%5廆��p@�0�K�7gG�`�ڃt?�:_nlQ$v�`���(�@���~�R�W��a��x���""1:*U�b��'�E�vpi��d�<]�-2�J�v�bө×7��UNg �w��3!�#C蚞���]��t^�<۸!s��[ן-z��M��re��sS�i�z�U�z٭Y�>L��Ru֝��_�?���F[謡T��k*���*ЍoF��ݠ��S&m-6O*�8z�VA5�Y%};����[�޽����ǂ�*�tzLV�F�s�O�V�v�E�1f�>�!?Ϝ@�\m�Ri�b\�. ��驞R�կ�(ȵo9Ǥ<�^��i�kϢ� �����
,~�����5r�<X��(
#��},�����t�ڤ��+/_���	?ܻa�r�_dP�c_��J���]�0�?9�������f.΢�Ƕ�d����P��O珌ȃb�[�ea�l�+T_J�]��C�n�^�۰����-���a|��i��mxm]	��_TC�*w��#�&ʝTy�IZ�-D������d���0)y�VG����ٜ͑^!kx��"k44jfj��h�B(=>�b�ֈ�5Bu<�3��';��3��;D��@Ȩ����A2�N9�8�Jx~k�:p��H��#T����wS��c$�J	�U��)��� 3���	yqr�,�v�ċ�UD�/�1D��(#�:�^Fw��q�ڭ��Y\lb��އ��
+�bZ�TIun����Yg��	hjM�����d����?K�Ѽ.戾��Lc�J+�������g| ���$5x>�l�3�β�}ӎi��^�`������ͨU��E0:�I:s�a�g�1c��p�e^�d���7,=ٗZ���O,�y���gL�*8M5��lkF?�=��'zk0m�v֪�X������(`۶�V���H��c�s �B^�HЈp,�p� �\c�x�T�Z��v��r�����Y��$�me��MMf��HAٽy�M�r��d��M����W�{_}��@�������pdQG��[���1|��?�K�h$������^JB��mpS$~��1�f'��pc5�`-"�_8�p�ǊU�p��� �oy�1%s��ᣁN�Uû�ӗ�Z�U�����'�D׃e�@,D0��C��h�w�6	�x_'U��a�)1�	!%\	�5�V�Do-.l���|�C�U��Z߽� �ʇ񉍤3�03�&+X�H7�)����}�*f��G��b�0]1������r_�}���";�� M��M8����x�׸�x��v��~��M2���P,T��`��&gZQ;-��}]��Y]L����7���0|P�r	�[�
g�rC�k�;�*�i�S�[k�bµ�ę�_������V�̑N���+'�n��'���:;#  �J�����?:��=7�m,}�/?Ls��n[ �`�&�Z��N~�)��w(��"zk�K���A)�f�@�GC�\�wM�|Rt�k�NPy�Q/#3]=�����������/�Z�Q�9���[��M�2���J̻����Ɇ�(�+|�W�s�t~���M�r�~҉d�_�h�G�R��t������R��o�ߺX6k�fv�OOEQ-���N�cX����|��A��<C�P�HFx�Dߠo(�GQgY,�1��1l��ӟ����*2�;"���sʙі1,8,�����䙁5� t���/�\��൮<�� _=�kN�Q��Y��7<'5���� ǵ�Tp��,�i��ܹs���(JRz�n��+�Q�Եh���󫄩$���DNKHF��C�> my�ޔ+�rh������O����dX��W�lMX��^��@'��}ϗ��8���/x�%��:ۮBr��(��'7��=qF�]���j�|/�\SA�|R��[�\��j#����9�Ԅ͵���N���[�^�ٴ�o�wf"8�a��.���
�*ԻgQ���9*]�6�Y��8_�V�f�T{O�%>�3��ްs&�-ۻ��7��O'B�̥G�)dx'h×�s[u5ٍs:+w�00j�e��#�f�«��!;��)7?�����+��ݔ�Y3��r�p����KH6j��jjB'B��
�����r�u���T������C�-
����:�?)~��|�Ö��[��4<�����Vޅ� 3�������̊��B>y��d����9�K�b�`�~��̚5	Vx���[�������f��X>�{0�bъ����.0{npK~�w��>0�ܽ�W?�U�Ć����3@"v����Gx�\��6����C7���m���� )=�:�}�6�kNW񙼯VP(z���7�1�A()��՟���D�
R�/�CNc42*��"pFgm��Y_E��1��V���l�tz��&�vO�7�8�n�3�
N������ w��+��y�R����$�ˠqj�N���:�ܻ�C"2��IEI�'��)/U�&,p	%2h]�<���6���H2ŕ���YX�bY�~F�z�(Yu)���t���d6k
+�i;�'��!�f����0�2�`��o��c��)�j)�Z��� �h�Yӊ�㼁e���ѹ�(��v���	N�.3±���I�+��PP�};�02�t
J��q�W㴅��9Xl��Qŀ���zy�-/f�~����.��_��M��X!̌M���˛�E��>j�עQb�dE"r- O��1?�}�Z`z��ea� ��*~.��Sg�N�t6F���§ |%A�,�n�����E��*/��M<Y��"�[jc�ʩ�88T�U��x �ؖji:���n�Y7 'c�\y�"Sa��AK��kQ��t[t��a��#��~��F�/�"�Fk�� 	̀$�Fѓ�-`��ɂ�]���d�7 ���-�[�z�����ج	9�O��>�FY>�l8Y�ݏ�mak�����Z�(�r
LB��E�ܰWv^1�1���|�F�����u՛D<��d�J��p��z��&�/���A�FY����ىj����=�x�ʮ�J��q#��d���S.��� ��P��ܠ�}�Ǒ���ݼ��?�k���� ��?ऱY�÷Zc�N���g���
,�Y6�^�$�u��MI�3Њ�^����4nnOw�А��N�v���sc끿��ĉ����ͥ��1{Nv��V�\c��A��>��2=w[EV�7�:��KB��u˃����G�<�;��:�fr�& �[z|t5툪X��pS׭�Lk͛(['�3MO�Eu^kJ��0�B���0�ϵ��7/�F�hc�)z �Ho˲j��ځ�Dc\��T����xi�����*�`@��b���WMè��lA��{����H�ҸŞ,z���űS�'S
�Bx@����4�4��|宒�n�#JHy�~�9*1=��:���^��W�(IyWu@�- 6�)D'��lbJ7�a
��	gj<B�Ҷw��e�S��S�.���(�5�l����q�����1f�ڮ���+�Ynʺ�h�=vCn�K=ew����[U��� 8KO���dkSui�.�8����|�/�M�:v���V����l�	�R�}_۠�%�t���6М�e�Ī��Ã�j��m�!Z����׃b8������f���b�M��^�_�CBE-)��[�2҇d�z�MG��HΞ�s��7�~��-ɬj�WX��f����l/pO���,]�8-�����q����e�d��1-gKd��R����g�h.��G�ր�me�e�9�� ���E�j� ���U�a��7��a�Z��4]ɡ]˙�b+���x��Q�Q}�m��=���
[j�0,5v�" �>o�o)��&>u�<uOZs��ȸ��i�\�s_��b��7����CkJ�`��n��I�¹
��@�-6��$!x�;6ǖե6��E�QK��'Z�B[��O���鏿?��$PR��f�2��yq��H��_w~�b�-�~I\�Ug�?>�9>�1��Mk��c4r)���W�=���\��B�&}�/P�v-'�7��{����K؟�{��Z��g��SJ���j+2E�|�X|�����}n8�����p������"&�6��f[���C��C���˕ź�� }�����\�<�
�P�ł]����P�6����0�I�tp�"OO_��P�#����,�W%�0�!^.�l�O��
�/	�*b��Ea��Kʂ��$�ծ�H���ck�T��=�=�̪@�E�>�鸄�u���	��t=%��;���	��<���S�Q1� �b�U�fn<W����g�3�%�r'9as8u3%JͲ�5'� -�[�P�-���4@�OD�B���ܤ���,~n��xs�����f�6����8���<rZ����Z!�}�8E�m̈���1���?��ny�'�Z(S�����5#+(�_���_�ȴ���}�ӭF�����c�.�m^;��������Y�PJ�3����y}�p�[t8���gXjc6_��Y�|h�=h���?H5�.�*������掅QO4; sw���T��	�E1@��K?[�����7"�G*�X껵�D�.}�d���U7��c��0%�e?����A��}�$���K>�v:|�{mw6�J�2I��܏���*�����G�d����1� ��� ȝFؓ���o�u<*�(:�����P�����	�ލ����Yw8�Bx���2�q&���&(%�ԧ�^.���rY�����C8$�P"�߂�Q��`<OM�6(�N��q�2���Bc�f��r��������^��A��4Q�s�T�73�D���/�m�Y��)����NiQ��Y�����d/��@w\�k�Sᖺ>�u�L)��F�q�X�ڧ��0�?2\�=͟��RčXt�-��<y���hG/�j����Щ���I-��I�{ĶMUv��1UG��r�����0���w��OA�%]��|!3�WG��!���s^�f��4<�y�6�^���0u��`�I�6�A���͑��8Vo��&��\������M|W{�����ܷ�Rh!�l�Sg!ch=EX���(����,�m�t��j�h+Xߣ�E |"�c�?�h�-گ1!�R���>K�4׆�W�c���Ų)mBM�NA${����2!��,�ףWJqe`��_J^�#-�B�:^���.�\�V?[�� y�@�of=aJt�\�N��S~pf�r�����X>W�N�t6tAa��|{Gt%1�B͠�*WRƱw�`����M�������6��_�.̟�ʒo\(,��~���������(м�2�]�Ь����,�y����	3��Aۙ�y� �5���
gd��sG�)�}OY/��_���JW�9�u�n菶,r65��k�8�i��(��"̴}խ���匊0��7�moʹ�\q�St�+u���S���TlS��Bƅ����r`Vdnq��=���J\�L���I��V����k긴W���A�G  ��{j��.���� ���n���=��Q�m�?�$�`�ū����%����6g�僦��``J��2��!��pP*�=��`�]}���\���z*P#j	�l�*�`�Q� dY,,�����x���ؔ_�4%#���ed
����j�ծ��v����JKcn �tΞk ��C�<G�쇚d����~&��@��)Ra���o.nc���d���Z��W�%�h}0ichҁ�x�� ���F����ƽ�1q�� K8Z+K�01��j�n�Ht���w�T2���E:/ej>2M�s�{�x�A^@��s���Z�����L0�@/�R��Wɶ�D.��C(�̬�B4��,��Z&ˆ8d�p91����2&8�Ce�(�;�B����8ѱ��{>����	k��o�>ªm(}l�mH����+Q��h�5H-]���ׄEj�-��C��.���&�༜;Ԉ.h	��xb�LHm8�J���L06v���׿1�%��+��W{<�����2n����|�P�=��'-@�W!�#����$^�fG����vo���Vi����E��)�Ś.��X?kMZ�YA�+q�/��f����bJx������}qC�s���XxyWι����Ϊ�6!��{u��z)2!��sl��ƨ�Y������n$b���[�u�m��+7��ɔ�M�$����4�V�|,�_�b��,�/5��ϴ;}���y7���q3��lX�2v�vV4���;}>��r8�%׏�pro��U��e\m*#��ySOX�� �u�_�h�k.
z�~ճ���|m#	}�W�t�Ey��W$'1�X�d�`Dy,�[���.����d�_�XZ�����ޢ��r!�g� ��?��W�\!�d�I=[~O	�W=�Q���,��Μ�h�uA���*pB*c�S\T�WI�22�#obbo^�u  PEM]r����v^�U�a'p�3|�r��)�?�݀�`���X���6��-�p��=r5�!1��2#���@]���g���(N�y�����$y���+{ldg�ی�t4 uҠB�M7se�} F)ݴ�/��rឧ[?�3U[2GI�/@�R�ޛ�̜�I	)�s��Z�#y�
5ݤ�.[�F������l�ÀS��s�$�d���L?!l��Q	\/�T�����%u�D޽X�_�3<�+�M��F8��@��k��޺��2��b4���Pe�φ�*��q&�Q��ĳ<۲#�Q�0�ֿ6|��zL{�T�2��]��V�H�{"���[��^4�����Jiv��M}��N?�g0��P�Q{Z��H��6,��RP��)���B/ ����F��U$��t���N��;W������2�W��\?�뀇Bw���ɢw �Ἄ���6����aI�l"Q���A��c�Ҹln��H�0qTS�(��M�m]����u�zd�4���\v�D�=�8��YE�9�V��5�h��?b`:2��������	�4Aw�����Uobs<�c�z	�)����6��K+�F�+IJ�,�UB�;R��LA���l�	�0L�v��w统r�y6��Br���pL�↼�2��A�P��A����T���/!�o�En\�����K��UNe�UJ��3����k-0��`�����Ǣi(�-�c��d�W$�9m�=�lL�a��x��n���@�g�5���:ZC͸($� U���
���FAv���3ZA[���W�nʚ>���h	�X�g�g��x�����Qx4�
8$�6I(�ȅ��ҹ������l�k4Rl��
Ŀ6t.e���o�#�&uP����w�86��z������9V7�~����0~�Z	��km��/��&�3GY�σ�\L���,Fmq��؊G6�w�1�"a>��6�o���hGp���E8p�q-�&�'��(vzO8�6[=��A|�x]�2 ȏ� �%]�J�gח*��G�:�_��n����;)��"���l̸�:$�8K�ɣf᳈��2��iwB� �2����$׾��ok���I1�/�z]^mv��q�d����߼�S9,q��Y.q �b�9W��I�K6�T�1���ic����%����dr~*�iQs��j���X6�.�=۶�Ur�ս�Y�p���
B�C����!�2�m�<G}��x�7��6�����G�y�����Tc/#�%6,���U�tW�ȍA\����BDt��v޳�U�KH���^G�M"|�Zo.M���L�Yv;�Z�r��ڰ��X���	hFq}�z���M��Nk\�vr^s�~x۹��`�a4��4J��6�����GÃpHp�(p�S	���'Ub�:`��j�4��}+,Y4E�{��XJ��k�`U !�/�ׁuQ���o���k=�7vd�≶�/���s_��+����x�ԋ1����=h�v�� �ꙮa3TpV1���a�y�j����s0Px��L�Jά�m�PsϽ�;r�T&aP�����1ӥ�_�rq�GE�pI���_�p�O�[�����o����iWS_�(,��!��Ꝧ��]�7� �`�;�6��_��>($�:Q��5�:�c�ɋ��П�?Y+ڂ	��j�4�>�u���6�H��WR�ĳ���C�L�y�z��{�Z�-^cFѲҰ��O��In4����c�6��W��p�B���r�ڒ�m~�(��)Us-M��X�O���;7P��IeB��MR��S3-�U�6����j�����]���P$����-�w<��4؞�P�0���3>jY�Ȋ$5:�����/�!� L���E^�8�q�q����9�����s� ���W��`���m�ig8�k��S�ݭ��VIȏ�����x�y�<LU%�:8e�{o�!��˪���;	�8�y׭��jhd�C�6^ҵ=�ɚNӉ<�3�f����(8ƫS�[�s(Ts��ͧr.M]VAeYS�'L�{�X|��J���<�&G��ny)�b�ҬX�65�D�#Tm�U��ґ(�G{��4����+��,�PRmO|�*�v?[��1�h�9��X����j�`�}�����W�8��n��.}���=������� �?��\n%��O-�B=�i�!�ݮ��� ���e�����,1�Iכ��-�Q�l�F	�e{�D"�=���K��e��)b�(LDĂ�)��%�_Ha���`�dt�#������o�&8��s�	�a�蹈�U��Я�$�t�P�s&���ř�Md��;I�c�v"��P4���1� ?EcNH�����H[�rޖ��r>3i�ڲe_�"?f�n�:��m*0J&��Q�ھ�vk{3cz��a��w�g�K��(�~U��ʃw��N���̀e668���9�WP�|������T���H#C�+j�%���ƅ��$*\�������>ϴF���&��9��M�[9i����(�#�X�oa��H
��^��#.'���%@+D�n����b;�������VG���}6��|��Gh�u)��g�d�~�l��j�xLJ��6K��tg�����sEޏ�� �=�վ_֎ǉq��T������x�}L���C��ё�L�a9iEl(F����j��έ���{�+}~Т�&A-ܜCf��k��$'w�0����±	����	ktY�s��A�y#f�|S�`���'r6➺P�n�a�U����.����܋�U������$���1���@|��9ö��A�i��j6&;��H���p���t�^֢׷i�l�(oMw��ӻ���|�7I��P93z�1 X�W�vZu�z]9y�@f�jئ梱;f2?��5�ϯW�b%��\zZ~�k��KP���~r���n�"�E�)��8i��ho�}��b��^O��(��v��<�g�MI��������Wix>�䰷�6/Xyg����@����}�y�l��b(?uUb�q��d7�mV�e��z���r�����í�)W6X��s�	�җԉ���#�C����B$��1�E�ώ>����b�ן�0Z<6T�V���{��,['}'�|p�#1�z�)���8��&u \�h���\p����P&��>^Jئ]�i�7PG��>��Ǭ
���p��oi]�"��'�A��oAM��
����9R@��!۷1	��qֳ��¼�r
�0z[����ZW8��b��8!F��	�}<�[��6U�A���LJт[ć�'ć��e�C�2��	���Tf�%�t��1K�e8�×�-��<h^��F�J�U`-�ǄXQ���Q"S2�C����v�V+�zb/Θ�Q��V�����j��\�)���
f�SB�H�A1Bt�*���_6^Nyr�#��]��F����gv͝�êmȒ��t��+������8��������bB���C�����A�����>g�Da�aeLR�Pa��ذ<p��z���]�0{2q�1]١3�V��a>tѺ�Q������0��n��]�����1�m��%�����yl1Ԛ��(�q*Y���W�Ʒ� o �K�1B�݅,���TK��I[�������5�\6�z'�?~��S8�9>��T��
o�[��AMH_&
���޴�G��<u0ٸ%;�q��x�:���(I6��AbO��nݖ�����8�����i���V�� 2����H�Es�]x�mւ2�3&�	wo��ʅ-��Sh��u�6X�� 
��# d͇�z��2�u�!X�Է-�w���}�Ĺ����m���'0Y: o@�@�-GCqDP7Jp�ٺ=+���Y�A*�<��toi�՝l�`v����\����^�
�Ys�gIOt��k|իG���I��`��K�KP,�3o�����:�+��5���)ohj������3]�|j�WQ�T���%=�gp�/'�����{Xv����{|��:㡲�����=�'= W-�����6/�v�8y{��:C��h�d<�{v��[H��oŠ����(EKeBZ��ь�?7TVƂ8tx[������5ؘ�w@�|�84�9>I�4.�}��:���Eq�R�|f�G� 
�K��X�)�>���w� 6(f4,�u��+�[,�N��dS
�a��d�:<=�����,��M���fcAM+ ��+oR�<�B�[�X�w}ȶ��5~���SΗ���^��"����:�D����$���{�Q$���˥-��R1�U��jX�O���s渏������������h/D��p*��V���Ѯ���srL�α�ם9��k���F$ǖZ�lr�ƞ�4+�*>�)�(��΂��?�eZ!Tr�������<_�T+��	�g�%�J�&G��2���(��_d�s��5��P	al����`g�V���c/�lK�UĚK�x����w)$-|J�-�� ����hA��iܕK�b�ц��m�Xau�;GLJ�"�Hsd�������z�ɦrS�d�iBa��`ٳ�O��Ѣ�v��R��9#*C/���nҹ�6���.	Nk��4��7���Ay�VL|�Xb�g�3���؄�hTe��К�s�n^�0�@!�cVP���=�aSB�e+���N��4�����Z��m�1��+4�l�LVfI��:��ZH9D:.�fB�++�����^�kN�e�k���;s����ݯ\"�.�7���ͨ��>�^��˼2\�`1�nIVz	A��rP�*��.4'�LgQK�2\}��9=�o�6�z��m~�|�<~�$2��Zk��C�Il ~aV��Ѭ��B!��R�����>�C�u5�z��;��Lq'{�f��r(�3U���S�4ڶlb:
"�p�G,j4�$�>��M�G]_��h�MM�q� #.V��|K�n<�^8( ����t�T �	n�n��qc��}@iB<�Ѡ�SĢ�׀�NT7C=�)IvEs"��!��,�4:��j�9X7���5(R�(���IԪ<�(lX�1?��KZ������虴]|)G��\�6k�[���R�M�r �n
�!)#�R�;}-ɕ3�w�kn��{������q�����^��Ý�N�u���RQ�);��)�Nf3�@��6A��6�7}�_�(4f�*쑍u|��mz��,�=�r���Bp�8�e�v��f��;�a. �ub�ߠbtKUi^�5`OU��R#����ZH�!�/����QUe��,�!,�A��P�a=�E1[c�M�FJ�"7�j��:�O%'���xU�&Mt��mL[���9�8he�����}�4S���&�֋ٹG��z����_?d�,L��˙�h���/�U�z�i���W�9�_t������g���-����_�C�f�YF/NÅ�Ь���\�2̊��K�-�z,$� !���c�:�:�E#nc4}@Z�w�is���#	�釧C�rƥ:!�
�
&PW�V"	����8���6��Z" ���5��Uq�=-���5��k�a�1�I��Dڦ�$�T�8'��{T0S��(0���/�Rɒ/[���JM�G���M���k��ȸؗ�K�i8�g�f���x�(< my|C��#�/Cx`��v��*�!��,�y'<�� �+�!�D53k]/s�����{���֩���oV!�M7Y�E$�ۣ3��6ٯ]Nq-e��n������i�|�2V��Y�*Y?b�	0��1��H��5G����{=�{D�>�?�+дo�5�q��E�'s\�������(I�)�D����_��T����0���ݏ�u�Bp"R:d�j5�u�;���~������q
��r���~zcԉ���]� �~��2�?X"6�������u�N�8���lhPX+X��
�O�u���n��4���p���!��!��p��)���ܡ���<�)S��f��&��o�6�Y�ך��%V�ᵖg���oh�\l�z@��a�R�h�>��|M'�{��1\k�>���B���CR�y`p�*�N����JB�������{!�fS�r�f+B��G�<��EԂ��(5�����
qKQ�;[h4έk�Gr���W&bm/��W��B+4�xW0C�K���j�)��W#��ڴ]�iχ�_ș���G&�7x/���S��>ɋ�՜-�x�J��4~텕DgS<�*������Yhx�z8c�G���s$6e���Y�< �s�t�`�X�=B�_^H���Ջ�gX�,rx��fy�T��UB?��5�)�\$X`*X��m�O2�^��oOe���KsR�_lÝ���!7��jު����yF燊�&�B����<�