��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb0(����	�,�
f���M��*4%����Іo��"�#�+�ϳ��⊁��Oh;݉_g4V^i[�൝�q%Rf��͠�xN&y:E�X���o��?��K��lbAޘx��<�Q� ��#��-�G0�ύ%����T-�s?�	���v��q%�����ҧ����%(Ǧ"-^ڡt������O�yMe7]�t"ϋ(l���F'e� ���� ��+-KJ^�d��H�fo9�آ�TgI�Նt���7��-�+������5N1��s�
�{��������u��f�J^ԝW��5M�M��K�T����^i�P˝8��0v���)q܄O����3o'HQ��(~�,������Z(C�kc�r���++���h�&��̈Ք4bD�5way4�R��i�l��V�u�]�)��t(��ċ�n�����Iϓ2'�j��qWꚎ�sN�[�F�\�����o�	Ĵ��yH�]P5%vµ&��ǬI� fIK���sF^	�7	�{�$�~b��wi9#��j!VoЀ�"�q���U��q���=�*��#%/�<�f:�A�9�U�p�N�h�5�ӄ!�<�"~��\���˗���B�n8�aedܘJ[Nˢ��.Ư��X1�RQT�e�I�ci���Y��M=���˪���Px��7%���l,Z��-V y�!¡o{�F0��2J���./�U@�tD|�қ�VU8�ŏz�Pa����=�3�����厣�7m�_�}�!�1�T�Uw2�K��χX��]�֧����*�:��F��0H�#��w
|��Z�"�,�H��I��]v��D�V����*곒����M����q�>.g�3�Q"������O�L+�
	��p�	|F��8�k���gߕ��
VYn�0P]��Y`�X�B=57��5z���9�W�2�چ�VK5L3X�ߗǀ�G'��u&�&�B�8���Ѝ
x����>�Uw�	Mۃ�z�)�����'Y����z��=�<qWPƜ}�A�a��(��K҉�i:"O)��aZP�"�#Q����j��޵��EX�>�U��e+.�]틺�ѫvjzz
���>�L��Oy r�]��I=�����l���QS��H0̻�7�Z{fb0kIp�_܍Z��Y
tJ���1 ?N��.&�c)��� ��`��+�/������eE}k ��s�2@_���5`��d�Q�n-��h�$�-lqZـ;�}�����!�}!
�uI5÷�Ņ��x�s-��GP�q�o�E߅������(�:�(�}�a14���l�a飻׍��T�c���}���B�O�}�������� L(�H3�yZ�a��1w/*~�	���eٿs^L"�є��^"�����z�~-KT�ӵ@`��|-Q���rۏ���~-�[�_)�����Y$�(���Q��VAϖP�ǟ�rk�q~�)+��P9�o�!�t�T�F���[�<z'i2�z曡=�U���w��f����Qh2X�xt���Q}ڄR�|������F���#�8P�1WK2�H<T�����_b�C�A�wW���|�r`�J�8� őrlĽ�lvAq�7���҈0�Q�5��r��B2θ�b6j�J=:{z�P�Ju�����d����t]�-���.���-Ѧ�l�&h>��D~�Y�}�Bjv����\P%��+M�O�;?)���K(���G�PέxP�3A�]�@��b_7�`)+m5�!;��+ӽ����s�ڧ!\�Y�>j��!}>kK0����t�rw֖�u Z�:.@$璧 �:ȉZZ����35�cnj23���=M�����q3�k����V�P
tt�&Uܻ���@�wJ"�/��i�9Ylc4�e<_��x-��9%���B��`���ٓx��|s�B�H��V$9������i����{j�D����"��[�x, |�%��Q��A~�vp���%�Sa-��ʢ<��ݿ�v�a��A@V��k:����u ړ �R�B;]s��H��ף6��j_�ޱ]U��	���=��.��"=�j���.�+v��˔�"Ҧ4��%��BzL�÷�m���Ҕ�&�Ů H�X�?��	a�I=)@P-a��s�*����i
��k��}�+�i��6WMW/���&�V�f��ג)�p�����i?z6�[��h�Vy��4�2zD[5��MsPT��[ݶ���w�����[.��w�pJ�t��$�yYp��,V� yD�E�Te�=C:T�1��K��E��<+vT�3!>���I[��!�v\�rN����6�"��2W#�<�L;���ר��JU�H��=�t�s�����X�T���e�lEג��E�e��~��qXt��0�$�f	�d~�$`[g.6�:) �r������0�9Sn�'a-y��;���q�ֹ�ȯ��2ڭuE���M���JY����A���V�dg'�d�k
-�?�W��]���-\o�Wxe��<2�]oZʊ_g;<��05���AH՚�B��	��t{.�<b��&#	�9w�@0?Yv�:'��H�ř��O�)x�`m�W'�ϘU�:c���?�[�֞{v�xQ��=�Liq
�Y99�`������3�v  ���_/�YCZ�����/t=U9J�1�ڄW�-�gO�W8-Z>TU{�;3�������G�w��;,�D;�aL�"�X�
�U�"C:Z,f����V=A�����m�W�%�W���� ��<(�K �чF�]5�)Km�����1�u�6=������vbQ�߬�T����U��wX����x���h^�:W��5��+���N�V��J�����;��� i�et�V�:�Aog�O��י�Z6�w�^�A��D�&i|5!Q`%ؓ`���<� �v�,5�|�9�%
���x@R�pT6C>sVpM BDu�2�3�e-	���iY�2\μiouu��y1vO��[J�HK���؈�0%ž˲�%}C����z�䛿n��E]�95��hA� ��v�r��O���GbI"nw���?b2��μetBr�F�9iQR����V����g�:Y�	'�}0(&Z3�r��Hb��n�즑�f���?@ٯDg��<j�Z��FŐB�.�%HуnW
ɝ�9�M�۪��ʓ*M����c��]i�������O~�^C�-8'v�1o'�^��`w�@ܺ֝daj�q�Hb�$�p4��A����%�ʩ�6��j��bU���V�w�0(68�a���o�N@~��
����ζ��=��.ly��K�$�$Pf�X��E���.��߁�@�8	.���.���a�7b�RP�����:O۞�����yd�	1z_f�j��4�K�HK��B~�nG@a�ǭ�+��m6�����>�ێN��bέ�q���[�/�SB&��u��Be
�T�w��toO?����9f���;��6��$���tT�dTE@7vdF���U"�mR㯛��c9��v�Pjs��!%oUqԣ�'rn���.�<I��s����x�
��3����,ߍ�E�
fR�2-?D!��:h�0l0��=o�<�&�&g���;�3�`�:_M-��ڑ��	�M�؏�j�8��"�[�������l�Q<�I�+��Z�YPb�5xD����b%�bLy4���	�p9�"���k߫<�f
�%�3l�c�F���p���k��d#��~YP|�x,�a�R�*�u��)�o�M�����-X�n��FֱeK���a�&��1�X���3�N����� Xl0H?S�䦘�Z�Ã��4��;�'���,���9R&�U+l��hjQ_���B��J����WN�v ����F�!+�J�x^��"����f��כGLVrE� ]״�N���`�w[-jD)6qQ���r�o;�����]X�����қ���L�hI�Z�F�)� �ˣ���/�w���T�ZT/1e'Y����ˈ��s3, >W!�z�K�`��qs�2BS�����5	_DQJ��E�G�n0��E�"UG3lsr°ʈ��d�E����I�����`�䈁����
�nꟃ@�F�}p��2��I��=@�Ɓ�F1�s��VS��7�L^X�,\U�Խ4������eu�����Z�S���7�����>K����'���D��5���hS�N5ҥ���)G��<*)L�{2��U��
0 w���Y�B�ҖH��W*�o�}�v�Yy�QN�=
���Zm~x�q�#%���++1��#�[}{}�b
L�)%+����J#��%1ܸ�<BN�+�D�6j��+luO�H�G�e�@}�0��)P̙ZJ�?)�B'�ztaL�ȩqnf��� �u�'[�e�vt[�����?��o��U���ҝ��m#l����|�e��U�i��c�ߧ;*U��"4P�u�� 4%�V�ss��b;T�������p+RS�}���K��ꯇo���㕭�}R^�mu�V��"��L[�8����g�%�a�/����Y�.9�G� |��|��tJG��#5Ҁ]��5�BT���q)����j"q��<G\1�]y��U����f� �f�2��䵺^���_�8i��N��:�A��"�iد�A�X�8�g97��� ٺV� !��s��J6� ��g�LO9����_��Q���A����Y�I����Ko���T��p|��q�Q
fa}T�/�!���D
Y�������8��D�"e� Ae՜½B)_�{�l(.�U_�ݫ_���:Y9wRV���qɚ���j�#AY��{{��r�z��F*���"\�E�E�M�F*�����Fn��u��% Օ�Q0N�)����0�����+��L%������Y���������6�
ru]*{�p���W���w�V~��b�N�48�B3(!�%#J�Y�V���{p�w6��l{%����d�9&�
u��Olb�R06V�c���p ��`J��^B%պ�'� ��J��������QI�.U���]�[G������4����g͟%�Ʃ�,ү!G�A��1�-�����6�}�2ߢ`-��W~�!)7F�o�š$�n��欬�-�@tbf�&#�d�A�u�`�N���W$�+,��b��Ϡ�w�^��ms��h���({��/&����ѽ+>^��R��~�wo%���Ur�����r�#?���s3"]57�l���P�LWŻƵ��{;�/"�]�U�%�a�Ty?}��t'��t�*��<��2,�U�%:^bγ_dF���|*nc��n�%ʵg��4���j���.��x5����	�IO�V��#���YZ��/��&�"�� �u���N4U����]���5	']#60��C��i��'��|��4Q#ߪfaFtZ�=X㊆�GP�V����7��̰ӓ!ҳ۸"e�͚"���E 6àBc��i(�i	���aݪ[��O����?��M�r����#��Ht1lW��֋9V�<���,� L��U L]��#ƺ��,Ԇ�vZ��A3m�4]�ѓ�+@Z���![D��U���s�R$����V)���ˇ��X�29t�{���t�!y�,v��3�(i��	��&D��3>$3 �}�؜��^�?�)4E��vOރ�D�.�=������ҩRX�]�~����}z��*��n��$�������� �qA}�"n5W��_пm�eI^~���E�8��!f�������҂6ƽ�bvTD�5~?J��څ@�46�Q�T�|���|��Y� �0��97H
atE$���Y�8$�"��v�MuYx�V�����������,��4�8m5�
����X�|/������������!�{�Y�v�����Z������%�?�#�B�7 ��g5�?�����O8��w���Ai���I�e��(�����w���*$��;�����YZ-�4���D�K$
R�v�{a��!U�D�j�P
Q[�ӫ�
}�a;y�>�VŻ:��{�^l�!-6�8�ñ�,W��v�Z����we�#��R/b�=�����R��}�^	,fAy�|�@`B���a�Yy�	P4��{ߊ�R���}���g}�u@����T�8Iz�v^��BV�e�$�i#|f���/Ҳ��D�"��!MD�^����J�����J
�|�@}���S� Ω��d[8��n��o2*�m��,K��@�����e)I�jE�1�e�Q��x[���O�V�>��G-c��3$j��}�y�T���wTTTUudD5��2ND�:o�"0�*~�?-��ju/0c��/^R�4��'a��z��|/��=�W��]�0��*R��G��)�!ېѭ��_��6NV*��G���I'��~+���#)�0����� z_םFC蝺���u�6�X�c%�:Ŧ(KQ~��P�M&�X��ϖ��体�,��_C���Zo��6�Z��i�������=1�h����������1+��H�����am];��t(���^�D�;�Z�i�>7��g��U�{�8�k�}<gkJ	;{�U�͢�����D��~<�0��.��,G?˒�i�Mq�9��5��n���~ ���F��#7�8Yȍ�{]ο��w�S�$F�3���@�<�X�ѓ�)n]�2�M�B�E�6'5D��\;@�>`��+:��J5���^x4�s���(ˮ�D�#�^HTd��^� �+1�w��G.{�~'
A>d!8E����#H�Z�>�q����#���_Y~Z��cZ{�)��I�*�=�����+f�+Ew���(��Ǆ���b?�HY�!�ٰO�7���@�D����$:�[船�{�`	��>���"y%_�y�U(�U�.q9g�OM��7fc�J�3�y
�Ԥ��3&g�EQ�]�Vt�Z�TH�X�y���3���1̮��3VCQbr��Yo��Df�z��o�"hيF+	�^�k�"+�#���a�x��J��;�,�H{D�
@���D7 h��S9���(22�Xqw��M�b�(Q�Ζ��!r�:�������۔B�����i��?FA4�,��P��ׇ<U��g|0M䧐� xU�ɝQs�l6?,���)�8��D��x>m3#��NGgEM'���Z��РQNcS��JM��=���]�Eޮ"/�5���V��4 6�B�&�����8� ��&���C�o��3M��N<�o����<��QM���=�ٮoL���j?��V����Dߞ�\B����[{^�!��&���1B��s
	b��KF˯4 $&�����끢���sn��8	,[��O�Y�������:���7���]�J���U�k������I-ʔڍ갠�+�+�Z��<�D��+���VQ�����J�	&��!UL*�/�pf٨�=Ɛܩ	�;��.?'��o.�Q�3 WC7��i������L��*Q%��r4�O�D����֟W(d�n���JN{�Ad|n������?ҳ��j -�d����������1�4�
"�gW�6t�����7I{�!TL͸C��<��n~$,"�NcWQ��u�b�b᜻��nJ2@�-�����2_����s{G3�db�A/��'�t�|.g:2����9p��@�my��.���U��0�^�΁��o��_)M���F�)��l>����f�͌�hJI�z�z��7�5~��S��ր�0��_��"jy\;Xf+����3�C�qr��J�+k�G���×��!YҬ�{f)�H�jƿ���o:~�
�ٴ�P���.c3]E�[�� �z9B��W0J�Ý�"03�5a��C[��~�E
��o9���i���OK��RB���mJ?ץ�b��#	�7��7=����o2dH6ޡ���R��ƅ˕��Y��!K��'��kД�T`����b*�t����髓8㎿og���;Yuц�R�< �1?t�kI�|����/v��s>(�
_uW
�;��0��o��2�Vi4���X*N��.p5n� �$��Q-�v�eD5�s�����Ye�������}��V=i34��0��37���hC�VY�œ�d��7�����TPw�*:p������ȘWtO]����j�y����vL`�P���`�B��Z<Bm5�O�}�JϤ�b���,Y��\�h�xD��7J��B�JYD�F��5f�n>�������m��0�M'��`�Mӊ�X���3|���N�fc���Q�!�e:�������l�Ԩ��Ԫ<�8o&�%���7�fե��3�:w�b��ό�X5N�դ��^tx !�Lk���v�hooI
���L(�6E�$��$��A��y��d�����W��˺f#��d����wS�'DЅ�
E��b3[��#��u�M��w��Oð<�M�;�� �E�J�8���p�?����V�͙�wKX�HX��)�ȊF�:�D󊇐�gh�]�j����Sה/�d7�c�#ef�C��2���9&����er���eN�I*�lDd�����X�=9��;�:.2�UA���LcRT�{��/�G����C�r.�o�l��˭��۔JF�A <Z	 lN�/�.�A�@uZ�V
�!��_,,d쁲�g}�uJ~��a�0���0��?��CL�4��adg*�GB3L���9�D��0BO`�5}.l
�0�>��̓�R���v�o�V>S랛���$V��>i��NM��^ܕ}�c �e���S�4�h��zm[�r� ����ж��~K�P���O2�ܺ?�w�jUZ� ����{\���N��;�kY7k�5������:ъEXˑ��Fs�	zH~�H�DM���r���������d��fR�S�M�XR���K� dۨOz��,�~c:l��C���멲ߒ��L �\U %��KG�N���!�pb}��ݪ6��2�����lf���3���%ˤ�ð�[�n]��5���r?4��:z�� ie�H�O����q�f
)]!#�%�&�$*&��ιV���6�_��¶�7�)H2���S�_[��8�v��X���4"B�nЋ-�{��s���j�ٯ�X�-�cH����H_�p���&���t'^�!��h��L=/��<�M30�fM�~=��/#�C���F�a�3*	9�;5�Pgi�W:]k?#y h��R�^KF��U�I=^K���|�w���Z�`E�<!�� �����gbF�>������*TO��Lj��1,�ɶ]��Q޿B��L�䭓��6DR�"ڎn]�9�`�D�cO�������޿�̸�iS��e�~ ���=S�i����B2`�c��Z`̡�x�D��ӫ���Nc�Ӷ#[�b�F��Ü��H��@���j���J�a�DQ<�G���oÍ�,����]�s������Gy�+�Hw|�a�1/4�k�SA�S�JP�Va�(�)o�+b��}��~�3�k�
S�����*�<��A���:4�j�5+Zd[M��o��Թ�KX��X�ƞ��_\�I�B�Dg���� �V��X��,�5��X�A2uʹL�׺"�HmB?��d�|�����֢�"�O2z�oz Pc�#���Cs7�%a~4�����2�k���}����h@/��뙊�Z~e�])+��M_BBC1Mu*]������V"���@�G_te�WO���xM��8~�}�f��	0���j��7��W6�c�x����� 4ZU��ׅ��`,�.Q����<��=y��kp��!z��>��u�����*z��(Z;N~�ͤ����5�I����I�y��qF��q���)�NzQ3}����s�\](ͻ3W3���#�|KT	}bQo�-f�u�g#�=�(�qn7��}ⓧ��+}B�]7�p���)��UO�
(=VA�޲1`(�[NNai�����rP��o����d���-��'��[_/�b�Ծ��o�n�]E��^l���b��¯[xأ�V�a�5WT�O_����Rd
�.��;v��#9�#��_�:L�]�x�|A���EφJ�;oyt��z�i�P���~,�e��tu9�k�7]�K7��]���44'[[xIN�H���]���b���N"V��9�O L�lLI�W5��#��ȝ�@�{�`��y��DH���0�o��=�En z�������ގgN=Ft������ �_L�y:��ٖ	����̓g󨆫�ϞNyQej�(q�$
2�z��x��s������+Z�����
t��0aU��ܱC�u�w�ǰ[w1�ﰒ����/|k�fT��-۵��
���q��$4|�=����{9*��V]���$8WnuA!���B�M�4�W�z�vſ`����׎l�둍nq��k9P��Q�]R���>_�7�ȎX3)����(#��b�1.5��f}=xBl�J��wN� g���F俽���1�?�'����"�WK��j���E�BX*�������N���z�? �S����^���#��O�a�hl��B�X����p�[�Dge;�i�0SS�Ȉ>�f�i�	 |��c�UMt^��y��Ltթ/�e*8��:��ץ�����Q�Pi9�����F�sa8����\��(��X�mkj�m|P*�d��}���a�G��簡֝;d��9���_�mt��ݚt����mk�v8J���/<��\\���O�fBc���`�ڨf.�����Wp��rЅM�i�^Z�%1����Ts�B�W�vE��EK�No&��ާ`����[���C<�f�8�E_���}[���6^��������Gӫ@W��MN���ΜO�,a,�y�U���S���� ��O�cm�k�<�(�;ˆ �h�Y�i9��!������Bܝ��v�V�w�e"��;�>Q��k�;���TD��	����<���뜸Bd*���I}����㏏-���f�&kթ�T��" 
T���"�h!���={�-���k�"��b��>G��R:��I��4��+��<�U��Ww���(��e��fx%\��Jbq� ����sT��+�"�����J��kSd⫻�d�ƀ�v^�q�755о�l0U00�h��1DЋ�i��Y�g���]9��;�j�d�s�����s�J�aS��F�e.P(G�5E(&��QI
6�i]ż��dB@��ʃk����!,uBȗ��"�E�	�Amh�}�D��&A��9uD����^��f cl�ܯ4A���^<���E��'�nxU�qD!��#�g��m�>�e�����ܼ-�v]��_8�*��b�hE������aXV�ma�)^8�2�S�&�:�oy«���{B����׳M�6�$���Yo�����Ղ��6���%��r��ľ����E$��7KA4�`��o�x&V�+��nmu:�yM��:���k-k�I��@��эsi�5�i:2�}�Y�t�*��Z�{����6�7��|%�8�=P��o«_��2
3;���RQ��P�ʄ�
,�.sfǦ��a@��;�n��Gv :���C�g�V
�Xzq��3�/r>�;��uᦱSމ5��+;�&�-}�x[�0-1���%P��h���O}�]�/��!�(�T+0���<�3���?�)����Ia�"��H�c�b�\�5�-�~9��{)�F胓�zp�>�|n�]��Q�!g��d�j��X��T+k]���]�E/�0Bãy",nA6V2���$��=d6��Aw���v�_���Գ6x�-�
�=��DhBLQ��A��#���q��YQ4N"|e"Ga�ʑÙo����#z�s���bh�����X�Qw�"�k,߳o��TX�5 �����j����"MPf>���ch��W!�5V����	R�l�k�\��%�5dg)��dT�}Vd`�p)U��z�:	��5�Z�o0��X;�RD�0���8W	�9��71��%`��7�:<�"�rd��[��~
k�. ��G�a� GWm-�@̈n�a��<����$�OA,*Y��7�$�V/η�>9���{p-����k
�_+�O�_�q���Č�h�]��-��\A�M�(b�zb�ڠ�b(|�����K�ۥ��"<�첳��'D�
�W� "X� 8GhHk�Q#�o�-�+�{}�"]>�j�������I����F[؈�E'��8�R�$Ӗ�jD(�*f�@�̏V���(��S`������ c�C��W��D�#�AO1�iQ?�Md=M�k���Z
+�{1�q��� ǚ��d]+�z�,j���fu����O|Fo������~�̏Z�0��I�g=
}�*��+;�^���G���n`4�R�B���n{8)�`��-�M��>ŋE�H�t�<G	W�eh!@9-P�4�[�=yz�${ۄ��w��<��HI��"��ɏ]�@���;�ۗ#Ӟ����^g𔈧��Vi�$y�t���C�+��L�S��U���uh���n�J�.7��V��L}.}ؐ�����#���xM��n��goC�K�s}�p�W�!�2��ݵ�utY�'�EF�%��1	��䡼E��jp���<;�
|�G�=��G�Ԍ�f�=6l�M1�s0�y-��< ��əO�םF��_����Ҋlu�DR��D\���D� ����$����o�g�,��x�14��f���u����֪\�'��k�@^�xִ�R�Yr'�y��2��C��@�>��{lWcj��OF06�B-:�c��ɢh�Leb���c�s�����ӵ���:�L�-f,��� u<_=L�[��!aGN��pf�[�a��T,�;���}0��d��/.8��Ή����1w� /$�����������O���	�Q^��i8d4߂Km�{�5�($W�ݩP��Kx����<��u	��ɦA��IKM�
����|��@I����K$q�;[mQ��K��K��7�M�� k��fbq��Y���q`F�2�}�)f�k|hfR�<�2�,�s�޿F��#t�>������ryc=!q��J"��>�C�T�*'4 9�8��d(-�,�?�6�׶�Xm��[y�!S$�N��u]D��@`jmnn {sZ���z� �W,���m�ۧ`P0�d���ҟ=L�i��p���<+�9`ۜ݋O��g[� �m&x�y���9a�ͅ�x8�!sT-�>^
�\ �����%vm������l��zD� �����\+�1�ϊ�C�b%y&˂�c�́��!sK���~�6����}�� ��S %��:N|.�>�R��e���3`�7ƪr�<����܍�p4�Z��EQ��4�X��vd��A�A�7Z�4������Ƕ{�(�T'y� ��O*k��a�W�q,*^�?z-��I��� �>{��Q�k�M/��C���/��˺jk~�2x�*0Z�&�݂� Ҭ�#����(k`�^���(_��ʹ ��#���~\=x�᳧���{ݷݹ'~�>�gUSJ��H �^��rK�g�Y}	NXv�� 
f�� ~\�a���f>d�i�Z)���F_�d�0:�#�sF�֣���1����'���g�k��8���xl�A�[�f�{�0�����1�X���2?����/�Tnfs��/������m[3Jn#eX!bz[�i{e"�B��6#^��K7de��yk��Ənc�;��/�
�d��'7�"׷&�d2ɘ�A�f��Y�(iᙙ缙
���1R���U9d���k�"�`��qb�T�*F�?X���i{��8V���<H�~sӕ~f�C�E�2D��gyˤiJ)`�"zÛU'/nM�\��G���o9����W�}�_O|������9�<w\���L^|I�������	����1�Ԫ����1R�o0�P�^�
�@�G����1M86�X�w����J��'}����(�9��)@�T����	jM|�H4#��bS�b��^���Vst݀~��o%�/�v�pI��RT՞.��+`q娧T0�# F��|O&�{e䲺Ɍf�5��X�s��R���.�����ƖOr�0u:���l�p��A��_��.�tL�T���hӐǑ��k������0�����U)$Z���VT�?Vݏ�i�/hr���ʱ̟=v�Rß
��楇\h��	��3MS�b�����	y�����g'%����"=�,Y�*wh�ւ�^��s6##�0'����U��"͚"g��XV�\��ȬF�PSy�R��'�0���@g%� ��]b��x�"p�ٓŐ�����U8��u���OOa�o0��i��ip���k.+}ѹ��G:��Q]�h�
������,&��������l�sVT��W�w�Y���n�s��S
��N&}���Kyq�QL��T°E$�jV8�.)$�Okp_�z
���lόO{C������N�ɏ]t�ɲR��yb����B<�c9~I�r��R�>fmk�G��-2;�60���R?pb��YP��=��B�4�/�Qq��T$�;�IJ�TB���H�O)y�N��L�{Y�U���� ׌���ȋ
J��S,�����Њl����	�E^��.�v�/[����4�a�ۼ���ՖA?��ļ�g݆8������N�Aԕ{:��X9	����r�u�f	�H��dc �}miz�L�+�h��e	�UtakT����"������T�u�G̨�2�T`-~l7�BR�ڙ{|�Dΰ������ro���d�bmu�����e���W��K����/W���"���C���*�`�#�5wsڲ9Z�8h�p����b�׹���e0��wm������'��b� aw�(�W��� �ƪ>��u�-(�x��G�>T��#�pm�~.�'��k�*��q�1VʋG�/S��Lˠt���,cTY
M1�Z���P��c"e�_�ReeЇiˑ�È�D1������~[dDdA�U@���7j��X�R�٪L{��k��Ѯx̕5|���S�S/s�@�(R��`�ΡB�֘���5LL;�����}5��Q�Z�?�*e̲��_ܻ7��e�E��}JyR.��L �d�5�X�����W�.�� pW.1��(���XzmD����B�Y�|��3�A��&�%Ø�����Ҥ_�x�.؍!!N�A0�qg�"���3wm	���x_6��\�4��-�0%Q�Z[e'4&�{�V(��Oݎ���JF�#ez}3��L@��`o󘗅 t0,0͛5)͑]�/p:���е�hՆ�;���ɓ_�W	e����~��3]�?r��q!B�*��N��xo�t�m�_�ts�=�����V�TWPY\C��Ϲ����6zk��n��B��l��P�;x����_<e�ȇ	�qU�C��,r���e�,fE��}����o����$wQ�;x���$����6�拓B���ȗW���m!����p'7%�eE鎮Nk�Ҫ,�w�I!z����	�� ;�h��Q�
/@���V�ZKI�X�<��r1[��yP��^������cB�ն�M��D��y�G�\{����*c�sTc+UeD��٤��!Ǻ#�L�6�!	� �N�s���&	���d�	��K`=:�U{l��k֞�} ���f��"%�w�9%u��m:FK�	q^����+=$�� �w>��9��J������T�\ {F���٤�~aI�tI^k��k�'2�vRz�iX���N�?��R���()o�:��A�hmc_`yo3�2̑��!�;�	q�.�L���q�eK=�2%�(�l_�"r\2�D�\�נu�˝�B�NT}�
�j�_e����;�Cz�'r���b��f���}��d�V6���C!چ��/|��i��~���9@j��f*9���ɰ�4�l�Nr�K�}>6j�93���|Q�69�^+#B݊{㖮����/���zO����f!h�K/C`�4'�N/���l� ��/W�LF��jQ�g���9� M�ݠ�����T�i����^��,H��$���&EL�G���}V�О�A<���#�v�Qp�ﱯ0�kE6!YV�y��k��]�S	Ϧxr� sXm<�T��߄�g���n�>��)86����r'����#A�^@�=οqh�W���V�~�wm�Z�L�ks��Fٚ�r�w�c��#�c�����w����\ȦhO����x}�j%I�&�y�(j�+�)
v��P���d�0��	��<r��� ����gj����U�Ο��Ġ��$Ø�%��Gf���ì:8���,����ɤ5qﹿ���i����n���p�t��0�:��'vp��){����#i�:��̤t�@h�Ć�6�t���M�ٹ��ӴntX�ɨ���M�;@W�f�0L���d�����^'*�г�@��8��Z�g�9-�岺d �|���{��a3P��u� ���o����, _hlY�'/5C{@ڱ)�QT>�F�p1z��rJ�x�y�B� ��p��R�.S6���rO���6P���I���7k��y�����qJ��Z�2���8`�:ڴ��}������
�B/;Q���[H ,�B$����9��ޣvf<r�+~��{"�/��DT��J�Y%L��f{���ҭ������*��ױ��`�;o�0�u�1+1'W� 1c�R-	)��܌�Yj�b�*�v���s^(��j�}��D�}�eԠGt:y�u��O�u_��\���dP-^�@]�O/�QQ׽ʁ#���Z�[Qyw��y����󳣈Ajk�ܰ7JA�NY�2=��ȿ�UE:%��p���v�m��82��|�]�?�^Eb��ReFsC /��:�8&��ī���Gڌ��Gh+�Jմb7<����ܽ�h�ޝ�}Q�6���e��Ʃ�`��h�|R�B����\͞2�Z�������N��㪿�2C}��&�IGu/�;� #�})1�*E1�7
�b{םo~�;�@��`�&�6���4�;1B����x��1*e�y�����̴��&�g�x�B�gX�����B�i �r�[m�GY#
P�u���^�:C����Y�n{b�5<;]��0��fl�5k������H�lHLG�������i�
ޯ���V���-��ڒ���
ʷA4�|�}g9� ���F���FI�E+��@6�x^D^ڄe�_O�:�uȧ�y>��G���q��V.�`u5�(�Д��%T< :����
2,B���_�z>�9����̟5Y�m���U�$P�'_�i�b���4����'���}�������C�Ų��ha��3��~Iٱ�h
�ի��X�z,����ō�e�����rKny����U � �b�x���[{(~�1��S���!U�*Z1DI�z�s,pvH��M�r��	z~����B�6l]b��R��KMU���m7����/�<��N��"�-Rt�MO��A�-��?�R&��G�<���=I\�0ᇀT�����	�������m�I����4"_��!L3�U+��\ج� ���k�4�����D���SH_y����윁�BJ@6�m��甔I���1��VN���]w*�����o0����%5��tB�}e��o~�S��Z�34�܈b�m��wia�����·��?���aX��u�rR ���4��2�D�3+a�p@V�i��@w�ʖQ�ML�AZ{�h����e��������o��¬榲X�x�7o��l#�ґ���b}s�Ǐ�&/�"03r��䍗w,�o-m��B���Û�����_<�v�<h��8�O(M��'���ɱ��{�K"�dD�E�k�r��6ZВTz.� ��1��-�{�e���uH�Ƨ��޳ H�t��Su ȕ�K�'��.8�|��6T`B'�x>�ҕz|�;C��%"0B_.G�l3���P�BlW��X�	B�i^^X.��=�re��B4{ !�y�r\E��h�}8:s���4^{����D���4Z"��׹#��c!���ԥ�Û�j��6�>1��=����%��AF�u2ބ߯�����ض}�v��(�P^k>�`u�nsUnY֘i+S5�$n�ȥ4�*���h�����њ�2`��o�_���