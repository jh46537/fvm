��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI���!qp�6ht����B;dv
�[�܈
�/���t�!HO;���;��.$?�'�-#ܨ��q�X `*Ƈ'�e,��Sg�Bno~����1���V�0HA�=/�c�����)7!/2�����&��������N��Қ	Z�G�i؈�7ХP��^��S�T���4a��I����Zp^�B���,��1�W�؂���K�U��=k{�LcF���)��Idᦿ�_�Jy�����d��iN"����#�,^F"��.P�P�����9���})��ւ}�?�T��;_O�@0�|&���7cgKD��PD��댜2�.��%`:N���n�@�8�ݘ55{�K�l��߆,��`QJ���ɘV��kF�B��+]�4E�`�8�`�-��a$�$$�.~T������n`-*k���_�il�
�J��j�E�@���tΰ�k�wʅ��Sԏ�ϰͬ���eX�`-]���s��ֺEw�i"���sŏk�zhk$�JY����k�D3�m�F�K����[��<�{)4)K��|���mj����l�~�81|I�&�c"~#ցG1�j�=LnI\�w\����������Dhw��ڀ"�H.��:�܁z/�4q���T!}?z��q����
�  ����aE3���Mj��c�Z�x`C;��xF������"/�����]T���$8i��3âh�x�6HC����[�.�.�C�-5��j�B�/���擅@=������պ�A#[힐>wx���W5�.�Վ:l�Փ�{&گB��WK�ɹD�?�R}��%c4��)��M5���^w��W�r&���v�0�>��\O����C1#=
�!�6ɂ �s��(d=&f���v]�$��G���<�Z�<e0- �bGY�\�����\�C�s�Y�C72�� <�߸���q2�Fjm9�������r��f��Əɒ��$9��Z&�Ű@�_��q�wd��S5N=����\�JV�cL��-�y��O4 ��� �}j�v�72��,�*��+�� ���C��14)O�H�+9nV�.��ȼR,�^�;����C�/@��u���Po�oQ�4�6���d�F����5җON�RJN�ScD�f�:���{-X���	�:&"�AǣT j�ΏXf�x���O����26Yg�� (D��j� ��7�����/��Ry�S���6�p�RY�##��S�G�W�`�_��&ٛ�6K*�׭����Cd�M��.US�p�ĭ��_JI9^(M(K7	��
�����$����#x�5�,Q����!�*�C��0CԹ$I��A8�O�O�Z���[c�%�w0���V�B��u�O�v �l*,І��؈����wLy�w�
$��=r�k����Xx�n��>"�����e8��I�����^�Y��ZS3���D�k|=��oRV�����s�N��V�NЮ��a��T��	��A퀱ź�݋����)��Ea$�k�6��{RƑҸ-����JOCZYx�K���ݶթ�r�g;<���Ӌ�HC�7/166���J��2ԉg�����͢�2���fȬ�$���\Ta��Y!|
�O�4h`���$;m}V���L��$	�k�P��8|
���K��.
P"ϷN��&yYY�������d��
 ���aU/54F�M�֡�5�)�Z`K�{)8�?������<������Es���|1%Z���ԗ-(���[��w8���v\��3�p����fLSۙ���C�B��7{������"��5��{@�v��t8o䧌85	��`S�~�<�� �����p�ꗩ�K�K�Ř@!>P������h���z�/������]pa2׸yG��,����}U��9j=�w�oA�\d�M���X9� k��@N�4Ԛ,v:���J,���*`3��!TJ�	/bq��b��y2���;8�*�2��<�:��vr�����,�����Ytb�ʜ_p���CEg�l��~3�����i<O��>�z�X�6���kW5�\��~�仩J�����H~�h���Gq�Q6wNgك.шϋ��b�xX�I	,>���lys�`���}m�@z�PD�	���by�}�[dI���M7y���!et8'�.�2�e\�S�q{{�<���m~a�o��������Id�ʲ���x�a��\�:dm�����{����<Zߙ�#7��L�س5�mLIx42Z��$~�s�K9	PJ��NqM��Pe��E�8�1�$���!*ɽ�lX�rā ���AF*Ӳ�8��5+��E
f(tP��/Y���#���z��N��x��d�	'����>_�O*��X��G1�j��?ɭ�"