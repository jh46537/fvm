��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V):��5�P���!�gPsfA�Qe���3��˘�?H�Ⲑn͐�R���6.哺6��NJ<�E}�H#�տ�o��A��!�x��T���R�V���������΁���].`R՝o4ߜ�WE���&����Zd��VN�J瞳R�JS���x<L�nW���-�w��q��f���v?fݬ�L��t9�R	�>�Pȭw���N�J�y#�	g��F����ʫ��P�n��C���,,�EH�ùC�b`�K�[Y`'�΋�D��D�S*?dA?��g��)-E���ގo�U��7I�'z"Hϣl�J7�� ��yh�-�7��4�8D��7�� O�(�nP1̺̻vFV�Np-�\*>�\��)�\B�c����"-%��>� h�t��I�n������tB%;^a|���vW����|���*��K�jI����B��p�_?��HJ	�ffe�^��v%cꑹ��SbTL��Iyע؜Ea}Zq݊������Wfj-�p��m(Y0^�;kXD�)��H��u�t� A�{�l8�h�������	\j��l��Ⱥ���q�tU���bW��� 3~�L�]��9�R'ޣ�W7Z�X��&��k��p�{=*4M��R�bys-�ӥ�a�8M|	��f	����tiF�g.���{��ȅ�0���Rj�����Ϭ4ѣN�|�?��� 2���k��	Zź���v������B��m�?Ak�n������˭B��|�!)�V��V	5ڿM��I"pa�Mf���3G�Dg�ٖ��4'xdƄ)��F��.��߈)t ���b�>E~�Q��� \j�Q�	Ƀ���ȥ+��,k$��t��#
�}�M�wG�bZ!�q1�)G��[�N{/�
���nԛQ�1n+��
M�x�8�oQ�3��>rZ1"ϖ�N�;T�0�0'�b]�n�i�暁͛!��Z�[�k|�k��Įwh:����$o�v��ʝ����H�=:e��׃�� �h�A����3��|㊾GBQ��r>�u�3�S~32��m� �SZF=H�"��Dj=;O����Vc'Nh_���������(l��u���0E+{Fϧy}o�29�J<R��B <+�F�5|ΆPz���>��"|�~`��:%ɨ��1�8i�|C�l}	�<�#������~�&H���k�NO?���' E�_�IYGv
�GN�3���t��s���7#�O�:�YE��E�����˸��߷#_BN's�Q{[�G�S����I�#m�8�Ộ� &��	�5h��5.<�YQ�&O�Ƨ�.��u|ņ��;�e