��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�%>��1(-fR�6��Oؽȏ�)���V��L����W�H靠
����������~���o��?+h7���!���s�̟ȴg`�AxeSo�zC���k�T��s��k��|�R���9��6= ]�].�������H^ZW��x�L(` ���$H���bAr}_hh'��+�[`��ڍ����ki�7V@.�%W�4s�|���Q�(��]�H�C��+����u�
1����Zդ3����-9�zw��n����p��Zv
k�`6�61��~�T����[�4u�d���u�I$�n o���r��پT�ʯ�H�� �0��lY��8�D)��>�@s���F�ͳyf�/�l��@d�Ovx�f�@��\�~^[I�nS�Ά��X,Ed-��,���e�@pJ5�T�m0Y�M�(0+*���Q�q_[1I���j�����{��z��o����A%r��l!��"��j�'���4��+��g�d��serO��r�,Ȕ�M�p��`�EߵZm��0/��V�Q�a�/���)BvQ����';M>9�l)'�f���'��������W���k��h8>0�'�ʨw,�*�o�``ɴ�A��v �{<>���sCN��14�Di7��_U�36$\���6�-����BV���;�׋T����/}x�)u��{���;��d������e�ѓ�GȠ��:���k��z�� ��;5�^,5�ל*ȋe�f�x������7�un�ŗ1��57�+���1���^oc�F���������fn�(���A{����U9
˷F���@ ��a�jQK$�\E�9��sr;^��R>a[ud�ԫ������5W,|�(K6l����睼N��#靊�o5�u��]0tռ����o��'���L���GߗK�]2s����V'Y�xݘ-�w�3@Y��=�
��HFR���6�ϼ��
��Ne��(:����C��!a�x)���e��-ރ������q-(4�?�?�cI�g��=��,�h���hsD�k�	�s,��8֙�����O�{`Y�@A[�4�a"l,�ܐ�[�K�VXҤ��	R�C�>�AOMJ��*�y���odGZ�%���g�������vLӝ�]{��i� �h�F[���-����x�?z����1O<��
����0"�]8C�
�C��/Ϯ&��^���RnX�D���OhΕ1\�I���Q�yR���������~\�,��i^�6�5����U=�[@�de�ճ �{m1V�t���X���_�,@����{���RҴ\��q[�7�BP�YU���~����3��:I���S����7�{�t3'�jS��Eѕ�MҾpd_�hhiGW\;	����M��g��k��Y @j�e��I`�v�� ���G{�h�W��,�#�ؗ-xR��6���T��%��I��j"��b�=�Q��!e�Re�����`5/N�����p� �/}sd��im���8뭎�LL��d.�K��|_�0�m2�-�pK�1+p!�n��jP��@Ұ�VZ�v��Ű�����:����}�.(��J]��/ja�N�x�!z�k�|n�8�翮�~����MsĽ�SK;bM�My�H�I*R)"��M3��Ζ]'
��U�K�zIZ�%RuQ��&!~u�cۮ�ؓYt��sH�쵹WTV��m�r�H^R�@t��kރ���s4�X ���Z�uu�:SbK�4���3��`R�CT׽��)��u�{�m\=[��b`i��F��G࿅AT,�	vq)�x������R��/@lzJ>�^P����ZL���y��'��2~���;x�&����<��N0)̛&��IZ=�Dp��,�l������EZ?wjU����� �e�c�4|�����er��Rt}g$()��W=B_�T���<��~M���;��$>�3%������u�q�zb(��n�f�G�I+��ҎU�p>!��2{���g�G������.��pC Sq0-�evz	#ux���[j�%^���Z ����ȏfb~%j�a�`��0��(���K��� ~�5��/W=d���6-Kg�)��.�r��AT�'���?9�k��
�!3Y���3lJ#���SYR���ˇ6S�!���D���H�@�̛Q�PLw���;��4a�g��w��	$X�k@��Z�m�8�n���J����i:�m<�\���dAɐ������軷��s���ψW�i�y�	��'w%�b_Eh��v��h7��<�Q�Q�$L;^,��%P̨�nC�M��`H�e^:�W ��v�{�E6N�r66��^@W���iY�@����?�R5>x"�Ui�-j��(	���$3D�������p<�K��nO,�]1�TFF�G=��h�Cjڒ�Lq�����曆��R���Dy�F�I��㒛�W�bs)�Uh��#B?]���sE�u�Ia��>:�M*�գ��a���N&K�ٛo������-���6��?$\d���,劙�PNĔ��\���>wpJ�qvxD�� ��E��rd�ۼ9M��X��C��|��n��R	N�ڒ���sm�7��tB����1��$h���Jj���e�v�N��NG�s�.�U��D�>�F%D�#�|r��\���8�e�E����'���tJ/��06����u�{G��u]U�F��b��?�������¾�TP�x�v�Шf�����j-ЮDX���!��D#V�Xmu~��~h�8��$��s���<%�b�&�Ү�}���vn;O�6�y+@��u�v��^�D���(�Y|�w_�Cj�{�;E�>�0-Gr�B�����.Fr��f�� �cP�X(A>(������5��K��e�i0W�A�`�G�&���{��q(1ϑӜ0�8 �.9�/��:�X�lF2
C)�[��h��L�_D����p
l������P�����%�ƈ�za�Q�˽�Yv]{p�����4����Lw����m��cz���&] �ZB���)��֕������艨2oR�n�G'�1��C��Æ�n?¼Hc�$>��G?q,t��T*���s�6ᩛ|�v)d�#��T�>�������؇���T�x�6�uc$G.�1�~����
�txNۢ�y�����D�8����ׯ�]4�.|��עہD��$W�d���ଲ�W7�p�A��4�@w����V�p��C%�Q�c��Nﵥ���2�j�m��\D�U䞥G�i�$� ���k�U|�ƁR�y<H����]�\8�f�Q`K){q�n��&`����x��6��ǥF���%�e�H�+�*�,�p=�`q��z������Y�%���T�S~��g�n��J��̈,8ˮ��'Q�@Ms_1�����s�8;C4���s�z����&�u6��="Sc׍�n����H׸��l�Ώ
�(��}���z�6Ť�Ĥs�r��
�8S( ��i���
M��9�D���fH�H�/73G�`3.����1/s�ʆb]q����O��tIM��r���.��:�F"!�/Do=���E	�e�F�4� F8�rє���4.��N��L ���R�I�[����Ъ��.
����[m)�P���2�Jh��"��PUF�|���p�	�ð�_�p2�׊�߾ n��#,/�Y3��6�1�N[$QrJ�ޟ^��N�3����0��_]G�|N'�?�%w�C �uR\��Z{	�Q���3XD���T�vv2�^�=(����0�IV�wQ�
e�~��g�Q�vp��q_<ߊK����&�윆��k�e_hd�l�����J[Ɩm.�eme57]}JR�K0�SW�t�_s�&i~�	<A��#��0F�ܕL1�3Kg�wM3��JfQ��/��c�i������{���g�{Kz�6Q��#bZ��S��[|?"���"9@�f�La�*LWaS��1��
7�)�\3̷�7|1Z���~N8J�Q�~C�)u,u#�:}�;O��R��:'�;=��Jd�sa�j)�Zm]��U�1T�������KA��]B�kU��-ZAʉE[��Π#��Oއ6M|�ẑ�O�+����&�]�)	�U˰�R"T�m��?���KF�9���GM�,O�t:��-��F=�=:Yl읨��ΔD5<z���@D�zf��N���?2`��2S��g
��MR�HzZ���[��k1��1�~�k$�Lb�TJ>_Bv����aif�����:�����t�5B>���y���m�������K����[�.������g��q��a��r��Z����e&�9�7	��C�<�)�!��`Kb��*�a�8���O�s�B���~��Ň�%��|��+`��1�%&�3�g�݄�����,j�d�E�;�d�	���s�7�RJ��<h�� ��e{%�T����οꐇGcJ����.�pVZƉ[��Izeo=�Ugh#}�ҹ��~��42��Z���nX��V>�I�g�����Sd��,��au"�z�~�&�T_�`�_M.�H]���d�"�l�/�*���r�h�x�8����d�#��+n�����R:�����3"��(�w�h�\��4Y�A)/C\��w�.�.F�*��y�O�dI=��K���W��V0��o	鲭���"�S��᪺����������kt�V)��= �m�)�@��|�������L%rR�w:w�$7J�΃&G�bS/���G�0�~�p�@����Ɏ�gGI��`i J�|o����v�iҀ�\��s��B�Z��Z8H��ד_^W+ �4�ߗ��Hy�R�;po���Jx
��k���W��<�[��l����1��)�nRS&�W�T�Y
�,��׺�¨����>�o�š|
>ʙ�&@lY5	���`����$�ZΜ}'tIh:8~Q{�_�����k �.?����B:��g�1�V��\��r��LĞ��� \-�a�ٟ�h���r`q({ߠ������Zh!�R�����\��$���"�A�%�B������