��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[v܎��⾍{m�@ީ�I�F�b�cb�J��`_K���Z��:�>�_n�t�W���cj�z��Z�`�3!�\l�x�|7�����˂!��� �!Th�)+����K�T+>��~D�j��(�C�L��@�|"�L��"�:�|�����.�A�`$c����"��p����',�MN(�f�"�o���|����N�L;k^X���RQv���a)��*XBIqt,���P�yb��+h��8�U��v��U�Fíw����~�!g�s��౾f(h�OÕjE��?+����QHA_��+(�ə�mCW)Cg���~| UH�$��߮6R��*�bWY��i�T��G0|8��b�Y�e*6���ah�/Q�Z��|�Ipy�P%��l�x�5<�c�x�d���
*:��$�0L>�P�G ����X�ۭ:ZD��l�r<٦���>a[2H�r&��|u�?	����`�Y$�gb8KA�
YN�[�B���7.�>tA��-��/!\��C��hپT�[��Q�ux.��e����$n�{4Š6T��#槭�Zw�UF����Pt��lb�DO�)����*^E�לͩ��*�_�����݊<��L���Iɤ} ��6� |����.�A���G��]�����>���욷P�<�7��򼨠:��n�F7	���_"P2}!�NF�����}X2� ������/`�h� zqӛ��'y� ���<��H�@�uL�C@�C�9Bb�Ș1 ��������r��(��v%v�L�7 �) ��F�ګ��Єn=��0+FAa#��Qcjf6QD�g����x����^�Y�hZPA�6�%��`pˋ�?����AW$���ģis�����U8�Vn�phW�h�쬇,��!���H����Ӽ[��l���"-_b���s��_L�M�+���"{Q�L��<D9����ݜ{F���c@��|��̣��H9�3�n��1�C��@E��
T��0C��N;#����
GP� ]���$^��SgG��x�W��9�eӸ��sׄ���dB)�$Jj�?u��vG���g�����yW��j�TJ���U��X��,g�4�Y�_ɾw{<޺�
�F��6��/-��]������PO�w��m~���������d��󏸢3Q��č�S��\�yvh`f [O��R�����_������ˍ%��`��b�m ������_��5�RЮ�q!'�E3����=}�P��Y�0��N4���rr	�2��`�������aX0��C<B���w��������y��b��I���Q�k��ԍ��+��c�����pAxB���SU��ꀡ��6�e1�3� N�Q�`z��M�#����Ґ(N^2ju�-ş�졯?N۬�;�m�i�b�&P�4o}Mʻ��W?-���X�1���4�ϦD�å&�'~�G�1��|]O�	f��Z�k��~��2���Fm������gA�֍��1�Le��"_&�1cE;��M¬,h����,]։�0��wt#tG�f��j���(�2+W?��Z�L6�h+��˽������m;�nX$��%|$�� '*)��A��RQ�i���~캎F�aႰ�t�{;D�z�m��h,ۍ��b�̹h�R�����/��Sm~���v��
���h8߶�L�5���Q��!^P�U���3��NC���s����wk�7��:N.C-�݌'l��W�	�#Ն���⑜�%o�D�N���*�o�
..[��J}~"}GD���a�m����1��F�n݀Uw����t�\iH}�}�T��۽����uS��!�1H�����.:о�e���E��f�4R+lm���k�;���Sqs�eD�K�\��n׊(��*����W��4���[jPWx��:�)����yfdŒ�P�����Y.t��} �9�O��Ǒ�0��PM)��[�t�ыԙ�%]���Y��a�(c�+��4�K*���f/�7}v�ڃ��c`��텋�'q8<���:<�M����.�=Z�u�nf���T��p:mN5�Dn᪷��Ouu�*�� ��Q�j�> j�����p����[�y��y� �j������lL^�b,���k�{M���*��?�߀��t�����'�e��"VL���bO�ca�Qqo�,��j�~�hXӊ	-��+�gh��у�D{���pK?��a�J�6=����ɇ��
�
�2Vwkj[}�9!�ֺg�g�G�to�/L{Q?x9���#AY����sK�Lyц��r��ī	P��~���t\��N�ٚ1v���U�C�e"��t޾�:�HZ��0�!^wz8
!��7�^+Gn��W|���I��'�Z�^����_�O�V�x;~�X��
��i�
_�m
���f��vz��0� �<'��ܐE�]�p-���@.�pߕ�����ՎBt��;md�@ �əf�{��&
������$'��P�:��R��=�,n��b����:��t&� n�n�l~~M��n ����nE�H#B�Jc�P�1�}e"�í�`�"9"ˬ�_趋���s�-U�h)���Vۛ�|��!��A����)��bx�߅�f5D+΃(����y���b:��V�g~_�@G���7�*s���m<;��p��3pX��Ĩ�u��XQ[��+��_e]h����� �U����TAjk�L��O��@���t^�l���;b�A��jt��'��u�E���[��؂d��)��8zǡv�D��`��N�_L��؍�Z�����c���5���Q�w`�������qu�触I���^�ʳ��<�$ �̫kMMj=�N$ZX����D{�\ȶ�R�P�I����!h��uQ1dt�0S1*���> �b��t����ϼО\�n=��k�����-�:a�i�E�A���zk��@�|I��I%�2qe�l��
M���Z��N����
_�1�pL`�ZjO�����&W���)nG�G��Z��h�Q�>�$�k��f�L�g�I2(��J]f�{�������V�u�5?^E�i�>���������\\����VJ@�0_�J\�#�ȌSÑj��:�� ��O���@^�Ph��(�fV;a��&�a~O���d���{�=�沤�U��p��$�`�%����h�5�j� N�I�Y���d������^,D=��[	�Ӫ틹k�ZO.�o����Ĵ>��\��6e��=K	��Q� �P��D�	b��K��hw5羽�`[G�O���ZCJx�$&t��a�}�Li�sw_��%�6�]�[�/�G�&ӭ_}q��Wh��*mCǭU��7�0���%�?)P��D���
8�W!k��<Ц������7��w(��	�o�+��L�z
��	�hmPJ���-�O����΄Y9�c)ęm�]�ۆ��T��XEIPPw���aV���#�&��)����B\�:G��q=Z��6���i��#:�|M�^:���dR����������B������*��T���+ꉱ3��§XH�K���Ѭ�g*���gqi+(ʞG���>^!�ɀ��� 7|!�U��Õ%�6z�z�sW蹋4閊4VK��$� ӂk+w�8x������׈���4�/�eo�JjD*uU<������0�ΙZ��Q'爞S<��x:�O�&�BT�찀�(�h�(�����r��
��̇�t��8�lq��FOvo�o�.�|��S�=��ʘ����s��lg�쥨�	�XZ�� �f���~:��gU��_�GPSz͓�Ԛ;���_"�(S��IČ����s�Aj@J�e��yY��m9���ݽ�mP�ɞY�$�*/����v`j����)�V.X��Kь�㮲�/Q6�$��NO	��O�W|ģ ��i�T^��� �ys^���[�D섎e<�7Y��ny4��c��0 rH�j,�7��kÊo�׏Ժr}�#��g[��.Κ	+��Ȱ�����-�쉙��7I���zQ�|��/��a���c��R.fc�st�P�Q�Y����3� �Ó�A_݈�/��O��M��㝨� ,�U��l;@��7���pEB�ۢ˚�����R��8���,��ۆj���ċ�r�'(΀Q��MV K�,�����:q�Ç&���NK	����9g��Iһ����eMG��3����iS�E�B%-:R���f�z��5X�X����U#B�ڼ5���@[0`8=o�e��������XXu����f���^����?���wu��O���h3����Fߕ�ؒX8<7��rFhp�����s�PL�d�����ޕEU���r�跇�x@����O�D��3�ݠ��4��F�B|�l҂��LY����/� j&��mT2͛�<�{��c~�<�Q���Yi�3�b=L��l�Sr �C�h��/��(�;c����=һR��	Pۉy ~x�WM��CP뗜���O���}+��G!�fbD��������|b���Wlt�
���n���Cs�QL9�:U_����o�3j���"G;��a�I6�Yi_Z�א@Q�딒�QF.��54�����>?�r�u[�����f��pň��aڭ�Y�P�{L��A�6�8���,�_�{7�n� �k��\�y7ngI0��S�|.)/��À�:F��p�����ÿf}mF�x��[��5�I_�����FYΦm����e(�N
�r��֩}������{��`ݨw���Q1�ҧ3	z���{(~���>��E#���	ɤ�(U��LIT��M2K(��,cvː�굋[	Z3�Ab�Nv���OM���H	�<\6��kl��5:x�A�1�lR�bnz���*2��P �!쾍��&��YP�?�������!�9�O�y���@r�`�cH����<�������i�*��d)g�JBx�W�ɰ��B#��d-b]�wNA�Њ;y��`Ƈ�C� �#n�$k�z��q0)��b�[����.n���3_�a�,� +�v�o:nQ���V�����YW�F>��U�?�e��] ��#�v�=�� ?�}��Y����g؉+��f�5r�!�A��Y�J��V_��-�Ѭ(k�j� ����R�(��&�����5b�����(�;0E����z@<�(�_e���A�ƞu��I'%��s���ea"GY�-%���I�M}r��[mN��=uzu���i�����[o��םƥ�'�q��/3r�d���xm�,��;Z^ܜ�{:�a�W��� ��*)ꗼO岑W�?�dx�d�2�AB��{v�}���<��E��&Z�IV��L�,�L�p�)ӛ&�D�d�et��VF��5rت��q>����X'��b���*���)�s��^.ٍg�T!@�L��|*\?��@/�Z�/̃?��#KZ{��݁>�%'il�CŰ�]�w(��;�2�j�q-���7����!�*�^0n����0��y4Q�PB�#�78����n\Dx�]��-A�-.L�8����P�M����QBD��3�B`h�rpq��~�;�Ta�%������P����Bm��K?�=��&��1N}D��_��|�.��=ZU���o}Nb�|/�Z��T�*�9)�J�?�	��S:�b����۲��P<L���bM[���">NDmf�N}T=�)����%M�y8G"�"��-��$���	��:o��1�F;D
�<O�L'��КTc�O:��
����~��K�'r�r1&�F�$�B
��n`7�w��g����\s?r;�d�'��"����<!�A�.0�� �w)�~f�:ɇ{K�a
"Ux^%*pXJl��w��q"���ϴ�b� ch��Tl�G���}�𣕿Z���ѷ )�>	�V, ��»;c3����+���z#�i��5 \A�y�ު
���#
<z4}-#��=:Nk�j�n��F=��8~���q(A�d�->�j�r+����8���ղ��o�Ջ���v��{B ��}��ۇ��`
�[@rt9j� J8���q��9Ӌ 9�8����|"h;�6��,ֆ]����ژ�s��g�h;��a�o�GN�I���za����M/c�i<	Ur�m[u��;)y��L̳T��4�L�ΫV��V%(F����T�A����w����	��Ⲳ8;��ƻ�WyL��@����G��s7bwt��t��e�>W���x�B}��y��!�L���$c&/�od�a���%4k&h���n��S)!� �Eo��`�)iYA�}��>X�\kP�Mo�:�%��=l��W���b�Ռn�����''Dm��F_Q��M��y�e��_ iO��Ch�t��5Y�z.8�iμ�%�Z1+�59�~>�~��i���J���i�r�7�' Om/���:�nc��	d+���%CfH�_��:ޞ�"��*q��ܞ���?k��zT���D�9}殢<��g��Wv�Jn��.7i�y]�<��?ZN�t�`C�8_PN&x6���f���S9_�PόMq��֖#�~(�����r�l�F��Y5f��r�b#���Ң��%��ښ�����b��|����|P9MV��}���>��� �j@a+����ui"�P���y�WAF�3�6�������Z���[��)�^E��bb��a�)ŹFH4 �F
S�͒�h�Tq�c;/VH ��Ok��U�Gl�`j�ی�.������ҭ�|�|�)F�f��_���<j�k�K���繭�ɇ�BAD�&���l�&���p#�
|���8.�A��(�;�3⾾�(�;���8��57��F>�a9���-�2���"o��� �N�Gn �.9ۘ�qut'!�M���Ô<�W��P?J���1Շ\)���A	O|�x7���m�.�����D��?�d�j���#+���%f���\}���.��$�?����#� �ٱ��ψ�ϑ?T�.��؜��u��uTV�H�L�^qm���6�ܥ�-쿈2�x����خ ��\�1r��(8�������a������}%\Τ���T�?NR9�k�
TU��A���ªf$�}�R~�����ٞ�Ӄ^�`�@t��v˔���[��1��M����gT�X�%	���d��h��T�A�#SE�0��9�����sw`e=��lѤ���+RK*�=��c0��ϲ��H����ld�6���}xǛ�[`g&�(h�f(�Wےk�{`������xT��4#��\�-`J�6�J&���V\k��r���2�eg�'�V�� ��ϔu8�7a�2���w�w\�K-��//t����$�d}nZsc� ��J>I"�Ѥ�v�W�Y��2M��-ݱ�C��Q�Ǘq��AQ����>2O`�Y�ԉ�է[��SJ��D�K��9I�����zS�~Y|/��J(��X���I���Yq���!��5�\��D�.�̯�3�5b�B�En;E�w*31��Q�x�ko�o�8?(<�� ��0jpv�:�T�/�u�1G��l�� .�΍C��^xR�qN��!�ct_Yb!�:�u��?WT�jܗ�h��k�JVk)͓�!{vߦLX'�B��)�hX�����
����c4c2��1�H� `��6�*�x��P�d�������ĭe,�v�b��it���e���|�P<�$�f��N����A���]��	�(�D�1X�Z�9>c��g��#�[��4���� Ib�GC#�у�vn
Ǩ�R[�E���;b��P�[M���k>�s��t�����شQ�TⓏ{[>`����^0��y����Q2K�΍8+�B�U���?/2�_Zg�D
�����6�=Q�/���MI!��g�fS4��fb��s'�CPd:g���z"�H���I��X�y'�&�L��Lt�E*��3e��(ޟ:�����K*��kc@9�Z�_h����!�`�ɕ�!em F6Ō����U��߆@�����B���	�m�F��tIP;�
��.��)���MY�|	l���_����k�j�?����)/<,6R��Jj�)�.���L��/�[�)@����Ce��q��ȁx�}$�@�Y��>K�����q�o~���Qs��uG��QV�'�0�0�Xq3DM��ٱ֘�,m�z�DMn��[�3 ��՞Ǣ{���}���d��C�5�C���/�M`�1A���V��;%֡a!s��y�=��1��c������ھ��
�Z'4V��n}�t) ���W��DP�iU�Ml��񌆨�mVA݊���Ȕ,q����U{b��[���G���Z��w5�1ĕ �f���񡚗ۮV'����R�P쥈A�`D&���h6�*�<�G,})�D���ȼ4�+t�R����#�,�trDe�r�d���~���~[&k�uA3p��6�6�U#�Ѧ���Y�D���Yi��C|�C,H+JV�= �؏7N�8 �f#���*2�Q��o��VT�ý���f�, ɏ�r�߰�][��lq�Uj�&� jk��;9�ne)Փ�;��*�����?��8mVm�7-�zJ���Vj��W1�&�Fr%������;W-k΋���D(#Tn���T���e���L������~���%?�nCY��m1X�~<(w���z&\�����Ⱥ�Cb�-�Ⅎ&c�ĸ��)�Y��z���A ������Pd�u�.��PC	e�c��R<Lxt�;���f]槔`Se�:�gS����G�G�NR�kǫ�5s$�03��0��Å�gö�w&���\5�E���H7��ұnoc���`�o�"R���&7-�ے�#��NF���Y��(9���%��@�z2�۽��D�y�5bG�P��3�(]�Ft�g(��ڧ�?�ߔ���T�Z��m�!x]�W�@[ƍw�U2����$����J�!��^� ���ۆ��Y�$�f�	*~�#@��N�T��[�ҿ�X��ɔ��!o�>HB�#x�հR�zld�Rdd��Q���J��:�lڈ1j�����˿�x`�����g���"R��iG%~���=���Y�֝L˵Yãf�W���}�|�A+�)Tn������N<��j������ �"B����H��v�d�����v)T�͏�!�s=Z�*򎦏�5�i�Nn��M���`����|{_�L}���g�	t��\MǑH� �C�3��ET�>�fe?�F[!{x'ж�X�D��yqr�'����bw�2��c�i¢y*C�".&��|8��	�H��짲�8���Z��&�
��Zj�ό�\���Ϡ����v�W�Y�c������?dM�2��K#�����Z��#��v�?�L�q�m��$��]�+�&{{u�gW�ܰcJ�\�2f{6Ȉk�T�`JW<p[O��(�Z-�m��,�Aq&Y��,�p�mY�@I7T��1y�5��^b���_�0X#`{���f{_s�qq�b�x:M�ӝ����y�7�I�")���(g���pO��C�0B^:��S��w?�/��9�n7�t{�fMk���LQ;�!P*IjSw���ߐ"ZQ�u��k
���0��D�u)��D���1��i�e_�^[Ę!m���s���[ƹ�v��/ɜ�����AR������$��,��u{�:�&'�t
a��o���2�X9\���6C���֠��]l�Yԧ����~e����C�Հ�>�n�<Q!�K��rG��S���w��ğ����cC7jX���G�X�N�-q]
�I�J	�-��K�cs�����ؓ����ve�#���X���B�?*jG���p�p-Ӫ(J鋊�h�%�@�� ����{�d ���v@��E'v�A��dG�j�j���k���<����Le�!Ǝ}��`p��`M�b���s��t:��O�|ux46��T�;�g���q�P�b�{�������'��<�ey�Un\�!s���qd�l�r�v�s�z)��k�U`�XVmZ��2:�eT�F�hh�`�e2��&ΜfMyDT�Z:i0ђ���ܞ�l6��=%�����F������B���.�A���Z&��m񻉭��&D>����s�?3�f�L?��S!��U�q��Z�w�J@,���"�2Yp�9��kn,�xK��;VFp2���4�٩����H�?��G3�7���,䭣i�*�V�P9a!k)�����W�(�_=,.F�	?Lj�5XN�nܲ�2�VK�|
)�LJ�~��X��<g��fy�?
N�H��$aG�,mVG��!}	��MQT��#����7�y񑗮H7�%jC�	ĕ�,�`k�=�6���x�`w^�O4�U�֐���ЧE�S�m���0BPV�+4:�U����ʊ"�;�]|����EL�|3�&.3}!2��D}����dɆ�ʱV�9̟C�1�Ux�/û�80'ϒgb)ʼC�|ЍBY���wӒ����+@�q�B���7�Ͳ�dP-ӥ^�G�U��/�(@�ٌ�ک��;��k-k�5�B�Dxm�gaw�q�*��zjxW6R�� �N���;��'� c ��A�~��/�@��JZ���Oz+��b����G^W�GCW�[�b�F&\ȒhDj�-[E+� ��=PKV+�l�IG�EG٥}�"�:�-���PŨ���(�G��U}1�e|��0�h��Z�_n�������*Z!����Jx���YdV~�X����砞W�g�y[�����Z}cZ�Eg�Q"��A<^u叓Y�O%��r�G�~C��G����&�^+�>� "N7�����t~�VN�x
OxT��wl ^�E����<��`:��:�����
�-�a,̫q�S23�C��ɋ�U���(yȌȈj��R��K@/��mo?��})/uJ�&���]���,C�~ �nۈ�sRA��)zw	Y����Rk(v�Ƴ�]�,Mb�݊��<���o>�M�U�C6���>�7����fP��RqcOǀ�vl�k�����a��E)�t�m��g�����[��-v�a圅75j�m�[U�B�40+�b;_�N_�����4��S�902^7zHӦ�Cκ�%Q��'���/b{Z�l7�7�>�B�~����Kաd��En���Tr�%G�$mpS����?�b>/^ɂ�?��h`q�J�<l
+�
��\ c��v���9�b,����c �8_�|^��e���mѽH]2�4������1\8�]V��ɰ���(t7�%�d��hpAy�|>��	|������:>�2p�KR]u��S�t��2��$'O���� �:.w�/�!��� ���5iC�}I��&W��~�VV���&1 �,9E�~�E-M}��zt�Sh��;��}.����z`w1��0n	A^�@n�5��y�s32`6KT4l���i�6��T�"���0fC����czZ�N5Ԙ}pmy��0(�8�}[��y&��/�5��6�:��^� ��<B���UfG�+��燺�dF�9>��Q��E&�m�q �Sr�G��S����Rl�ێy�5�*}_R6�g��="���S��V�?�M�Ȧ���s�~�q��r��n_;�F��(�0������^j���@����۱�x5<Ʃ�E8ũ�m�Z]2P������I��	I���Di��"�&I��YX���:���5?�N�x��(���Y�G	 ��N3�����j&��b�-����/���a.���j��0��j.�=�p*���Ԍկ�����o��)�,�#.�u��n����F�'���ĭC�����VMΡ�I8��Ò���8�\�#��[����b|z�RZfA����:7����LX�baۃ1t��H%q��(�F���U|��3�^i����U\2�,������0*�D�����;e�~-�(2�Pt@�첧�*?�Y�F�S�I�tOfN�f�;����׏��y�>E#�TJ���� ��m�"_��G?�E��!y��<��0>*��ijA��eB���Y�乛�l(��yI�Q0��0�bEM��e�,V����x^�=/����bK�ؑ8B��`&�{��P�N�+�"�b�0�b���bR��|M�^1^5�����9���{�>݁����ٺ=^���/���K~<�HOZH�W�ecZ*io�`������?�e%R�>th&�WE�XVH�Y/��_�0yUQF�p��YM�yd�~�j!ZF�N�R7m�y�p0*ZHb�����0 ��m��/��֐ʬ/��f�R��=�ʬ�ҋO�j� �Ne�����M)['6�3l�,�OE����?E%µ�*bx��7���5�AAF�����3�1�>��ϧmdi��t]�(�M��i+���y9���'�K�Ѣ�[_�#���=�qX��IJ˗$�&U�e�+� M������Y*�.����eH��<�Ձf�V������1���������#?����)�jK˟X(v}�㳟o;ϟ+gv��1{dIK��zP0�<D���D��MG[%�0o,h#G,��?8�*�Z�"���3��N%G�/����~�UNW��&�2Y��M��x����v*e�hly�}.zW
".+N�~Aihol��S��!A��yC����aW�[]9��CQ�G]�9��)�T�c�*��j�l�
)�e����R�G�hn~F�;��	Bǂ#�b�f�D�y���y�RY?��[:u|�Z���&5���[�61���KN��I����xWFs�r�	xQ��MT�\��7v����xs2_3��;��;� ���.���4M�?� ��<�]uD�+��)�����Y�����R��D$3\7cm�9w���X�p"� �X�Nq����&� �k��rܰ85���,� &�E��
#$�B���k�
�;#�3]�6}�b3���K�W�m��&���&J]뜭��H@�H�)">�c�N��Ѳu��B�.ο\O�[)�����&x�].� ��q9�cL���\x��7���n<�^��d�a`k�$Я���gC��KWUI[�����:��8��p"��|�>X������#.�`T:4�A�)�MԾ�[6)�r����О����\>Cm1+U*�ز�ࣿ����ܠ��O�ôѨ�{�#�xjr{�����F1R����W���{K�D4ƆO�]���$o�����&r-�p3���vЃ^ٕ�����o�����j�!5�)B�wMܛ~58�Q��+x� 8�C��%8���M���B;Ϥ|6�ˤd��%����MO�Tɾf{��+�;BK�A�r�,j7	�U}�SE��g
�>���BJF�Q�b��X�Q�
.UP���6������g�L@�.m:&��ػ���o�u���$�1)�Vy������n&��z��N��D�>��%[�{��uA�[c}Xd�t�Jf��v[n�L���~t��?W��M��"2?��jMζ�0m�%�.4���B����
q0iD�W��Ʒ;D
���~��ީ�
���bQy���r�S^�ٍ�$d+;F�����B!���腵td�JA�Ѭ�8W&�0IA��?��Σ�zM��W���,���-�?�/!q�/�=�Z�f>��G�Z���^8P���-��-F��Y�[�>Ԯ����Y	�:G�����ܞj���ZWo%�l=���}��&gh�ځ%
���0a�ҞjCt���bFb��{v\%�����iBF9��ĮQ�H����j]��;	�P[�;�r�2^��<<+��F��J�Cm(���oc��s��PjWG/l��.Nm��
��o�Eyo���V�G��l0�YPJ�`�[��j�KpP�R�%~���x���q��cCI}�ܾ�J�q�J�)7����{ï�:D��mZhio�p%�Қ́�����(��mN�#7D���8��*����k���$AǬ�X�����~b#k�{y�_�A��V����kc�v�v���9>>r1���zx��PTT��ݧ��H㱪�t�Rj�Vp'��q@���AFc	��r2�*s��ˇ'Y��Ze��].���S+3����"�F�~����r�-w �艴�l}8x�@[A�$2
2� �/�\��	�2c<���sC�+��<�B�����#�'	�ՊQ�=�vN�����l��ĳ���\R���P��o!����(U�,��|l�.�,���y�W�&�{Ӡ\/-��i�.)� ��<�] �tf�i$#���z�HN�#�Uxc12On�Ig�|�[�t�`�w��+ׁ��O�V�/x�.�'K�7$��.*`��s��gS�b.�#r�,�6k
']�|���z�σі�q-����r��eZo�4�_���7���>ȯ)ӘvL7����I&{���Pe���sr�R'�N�C?����8�����b�g�j[1l�K}���K��DX�}���h;X����2�[��Z����Z��Y]h��i���~/�w@ ��<� �_��Ȭ��J����ePY_�7�)D�����Z������%'u���d�w��w��4�B뙼��. 3�%� ]3����8��T"����vsZ�s�������µ�^?�e�?��#��8��d)������o?�~*���]�q�POe ��a��+5�~�m���ƍ�m,���7�[��/�IMqcB����EA~A:��y���1�b�7-[7��,]"� �0ŀ_��ji��
��O����� 9;�mN���E���3���nX�a�%sN'4�#W���Q�l������P���3�ܪ�Zu�Zb��K�9 ���s��[�	�\TN�Q�}&��Š�ա?3P�@ �򭳛 F�ß�:���b��R D��q-�z�[3��RT���D�G�W��6'\^5��^>r�ي�VW���b������T�����{#Ұ�;u"6$���/�s��7fu���9`���Jr�,\j]�����Z��ͳ��+��/E�FHR�{K��pe�[.�Kg���f=�;�����5�b��K�OLR^�*�C�h�oK����R/��/2#AX�ycn�<��ޱ,*��:���Q��	�G���;��#:p澪����
(ɞx�8��d8�x��+�(Ww�����>��K�,�V|��'���ж,�-�eK���G�r�h��#y���E��3����Q����t|d�\�m�0�Z��$��&�GK�r�>S%���Q�`T���0C�w��h����9��ʚX6Ď�ȒrK���
JK�d�?���OB�Ep�Pa�q��}�` ��r���k�ߕ�J�H)��G9���L_LV�y';��~�V[��0&?^[/�����2�䴪��;�>�9�/V4Բ��-�����t�7hJf�N3��<B������$o����yU2]פ+����>Vl����=���p�ֱ��pl��4Q^�ǋL�Oc�\���%IB��f
Q.'Mc�*��@�kW6���љ��}������J01�r��nd#s�� ��T���з	vt���դx�*M�,�f�r;qP�k��R�
>Xg�Ҭa!���A�16v�-�v}������ڻ�t�v��u���4�Z�\�~�&��Wm�V_i�,W�ʤ�= v�"��7ߖ�ҠQ�#]�[���7[�c���`&��q���tR��&�Q�~�S?j&y��Ǻ`�(�@��TZ�����1� �=��eE\^䴞���1�? {�L�>0�Q�
��֚�Dx	|W�����]�-Q�F�g��@�r��ݐZ��a�(���λ�|<� l&������2,��A�@ZF�HF�����]e�Ó�.-
��o*�w���5�<��� i�#_�˙��2165�*p��ţ8ݺ���7�����&��J��n&o��ɤj9�^��\�)�*IáV�z�;�xu��W�%��M�2�h��Wo�ǀ�eQ��=��&?��Dt�h<�T����R�&�xv��L	XJ�=��/�90�o���(z9��ZPi�F�����o��k8��.vO�0��,?�Px)؃~1 öOP�/JC�}+�9 ����~gI�r��:[�ow�U鐨�47��������I���ozj<ƻ� "+����w�Q,�n4Ա���
�&��#]Ll�H���)4�V���U��Ű�y��,���YK��������:;�6w��({Nv�mwf�j�w-j�������"�Yf�����O?X��Zn��1�K����6J��7���L�{Ĭ�>��=`�CCnx��,d5V�a���8�iR8@(ݟ�gun�<.J��~��� '<s#�ξ���:�NS��\Rc:=��;2�'`}�������!�N�46�F�f_�0�^J!l���CϿ3p�Q��4m���s�����<r
�ҹa���K��|?�#�O�;Ț��vѲ�W󒆴B
����O��'|�������������z�B�����)/>MBк6��ƨ�Q�9��S���;��!R�"�K�������3Ͳ*�̲cH8Y����s.")��F%Ut��dT�#r���'%��2,]K�3���,8�hv���Qx\!��BpN:Av�a��R��:I�i�ѧ�����f!R[� ⮥e�W��u��/+2"I&��%�����`�e����B.|*����]�M&�]��Hãz.pw<��S
C]�<�r�]hy�Ҧߵ���ˣ(%����-b5m�2o{�ÀYpJg�m�癏"���*m'$8��������Q� ��W7=I���i^���}��R�~s�q��rd��&��&����j�[�Fr��M=2�Z�'=7�dJ �eV���2�_�`Ƣf�'�(����d�5x1����ڈ����%��k�Ɏ�����*�p�������; �|ÉJ�D��<�<�Tn�-��BH5 Ȇ�nO>q���k
qA|�p��>��L�aS$s��Oș	Ӆ�iz�k��[�5H�n�~y�<�6]�����w
�����=<�6j\Yכ2x��eo�R8$�j4��J`a��t&�~�����=j��P��!����w=U�[���
$����:L��^�^����S��PO^{T�E���Q[Y�yr< 4o:��]�W9�+}nz}�F������B���p�BN����j�Ug-Nƽ/S
�MBr��6�oW��c�XQF��@��,�P���3����H�YG揓��8�Pl���ߕ��+RFj�w:\SKj�eU�"6���#��Àn���@�:j��efo/e ����i@��Vx#h����>iv3P�͓�@']�a��n�*q�m�m��z���3������qaC	#��|˚(��h���.�E�}B�PIa�tAOl��N�{���cb�����0ؑƚM�@x�����{�98XL�����8
�jh`d�x�?؃�6��y��~-(��W�4!��{s*#�.�O������������V8e�;����@�U�I1Z� #�}�yQ�$SA�����i(�ȳ����D���=L4L�N�J��/Y�W�2��-��b$����`��9�:�_ 9�5��4�a��e(��S��ŝ�i�j*�Ƣ��y+@|�]��S��t��LB�-��M0�.��a�+*?`z��SDdR�)��A�"f����04E��w��"�)- u��[��Yg#���� �a�_�y��e��M@Ed/dT�eW�iμ�U��8Q[��z�dp;�6�X`������`|��ge5�2��fl3y���mP�L3�#B�}�E�NtWdFW�\	��
��ۍABh��1G���{F>Y�~��v?��ܞځ�K0�!:�ӓ6�Wd��Yp�"YW٨��;g{��Nw�t�XR�h�gل-�'���k�v͜��ı�S���Dr4M��s�~�_�{ݥ(���&�@�� �ET�HƬ1 �0{�-��9���"u2$�Kr����4�Xk˅��ȗj���j�t����@H�?z��ZE�n��˕%qB�acL�b:�{�n�{3�\��� o ��o1���~#�ۿ��5s�'n��ah��ކ(\���n����)��DJp6�nZ���S�W��^�R���'���@��W��<��O ���B���6�1�i��>6�]+�iHV~NMa��u�0ߚ:_dpطÌ��f�B�J�Z=�i�.����k�@UW��L��o�^t;3�ǽ1m7��Gc��왲`�2ĉՠ�V��Rb�ߙ�w�<^����@+-��Ì]x�q�~`	�"+����*���?�q%d6-g���ɵ�8Wj���"�w}����ђeqy�����,�3tI�߇�ql��g?/#��S������:9o"%�FT�
_�Ѿ����@��Es�؃}��G��>t%�2Q����?�چ^1�=d���g_O�$�{u�
-_����C\�?b��Ɛ�%��j���+2RTj���Ha����n�g��s�X�	��t��XBe��kCq��g�Zt2�P��'@��b6�!~�]d5�]%�a:d����(�³$���A�Hc��{�)`2�7�	'�XZ�n��l�]���ĸ�{BqGf����
�^�׷A���nՉ!�|�}`ȿ�8�w������p|e��\N1�``����V���UG�ύP I�pt�%JĿ+wN������H��7�	������L<�{KC�"��\Vf���e)u�� K��x�Q�D��y&�������0�s��562���&��o�2�}#����о�~WXB�5@y�P�/��Y�}/�P����ߴ��5��0{o�n(���btV���#�����¤��݊G� o�(m���%�?3�F��]@"T�h/����kOEhP�cI(�HDG���;Tc�� �9
������B�ȳ�^�X�K���W��.�y�d�r�T�1a3N�FY�+�@��C��p����[��I�����.N�ַ����bV#��WX��I~�@�����9�Z�%���'^=�Y�*P^��h���po�>�yok7���v�5��E^c�٧Ӛ�ޫ��ύ��g⊼<6>�@���2�T|,u��ID��8Փ*�8u9�c4N���x� ��ΥZ���jЙ͊(���g��z~�3�4��Y�mJ`�ȴT4@�{?��&�uƭ�,B*G6an,����._���i�����av�ܐ�w�ۘ<ș�'<�E��p͛�>;bY��-䲽���*���d[i5�8��Fʵe�ճ���7�ӌH�r�=�e����$��z��@�<-��_������l�����0���	�	��=�5�	���ߘg 
؍B�u��I�������ƭ���(���	 x�;�7�8�ɴ�w�Je�9`���R/}\z���5�	Z��˂�]����#�2.cӠ��Έ�p��9#Q��שּׂ��g��(� ��Ѡ��6u�;�5��v��.��P�楇��k���f�