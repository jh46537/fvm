��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��_)��%%�.��D�ֹʮ��������7@��=�y���fA-krT������&)���N)������&���8Ol.4��^�t�9��Ai�����q>��*�sv�_٪����qT������\��=�"�R2
�D��Y�$�c���]�c}��Ă",=�Dm�@ B�Ňm� �o�2����c��o9 c�)B�wy��~&�N"x��#�wE�>�J��$������% �YdT^�#���Ϫ	� � cY���A���Ѐ�w:� ��fg&�7���HE�(��L������7agzI�x�ZU��qo3���z�FĽ��%fy�'g�3�Nuq����R7l�}-P��xv���+n� #D�d��b�p�c%�������C��9^-G�w%��-e9I�G�g���|�9ғ�H_�<	�Q&����C�y�z��2�����(��j���տ��oQ�S����Bm�>�m�"���5{��� �U�^�QϮ��'֟��
g����D-AR�Ə�d8�z<z�X`��a�����8�L��e����=�þ��׍��_� ���8x/�(-!d��;3;1��r���}2/Yx1��4�{v�(��&����Kl���a�� �AV\�� 4�x�4�DT��sj'h/��]��Xc�M��
�l/N��O�wr�d3��)��p��5�CCk4�˵�и�惭�m�tԋ��M���o�JWJ�~R�H�k���`�b�(�o���u&z���]���Ȫ`�Y*��u?hMr��u��@�m_qU.�K�d�-���Km��`ֲ���_.~F�=�䘦��(vP�d[�:�z����NOu4�9�����F�F�W�6҉>cI(ӓ8�+w��ɘ�b���USk��f�����:��vz#�q�����҃e����JN�,MZ	q�
���0r�OG��J�wg��w��B�˱�Zm�T��%RC�J/�.�jY6�Fm��ģ\4↝�k�|G�jm0]5VQۼ�]����}W�!��˯/�4��:{�_		q"5�!�1F늟AH�?��C��Hv�LVI��<�|ʀ�2D���ih̷2�ڼ��"6F.�^��-�k*fu.��!x^7(�T����#��b�<\��[d�s�
s A�+���ԡ�nk��	�xG/��V��ڱ��Օ�X�v�/�jܒ����=��%l�ܨ҉|:C���M����ӻ�Dt�C�e��g��L���#��	l%g��$|�̶<.]=�t�~�V��e\�/f�Y��Rro���a3�S��(JBc<f��nw�i�T�/��NB��S{�*�R�%d��Yo�RҘ�;r/-�:y�#Z�EɣSH"bk�k-k$�\v�e����E
��t��e�L�w�[m!>�ch�I�����*�b�v�*#nP�~iD?�+��[�7��g:��!i[� �5��خ�E�/�z=/�W�4�~���?,��?�2Gϲ��~$y���E��U�n��Ô]�G�h��]ɦ�Wh��Y
���'�ԁ΁�G�nϘ� '�|O"��*����_��6����,�\('ZL�J��4���[��;��0s7�1A-�0���t��э�xd�����?yK����ᵗpF�5��=�e�3�Ɠ�pW�������Ȟ�o��]Zx���*�!6l���ƦW˷�]i�g�^�'��>�P����#㉎�{ۼꖣ)�m[!s�:��!vu+R)W �dݾ{�Pm`�����f��q; �R+�]��~ef��k'[q�P�����w��p���9��tRI�X�X{��x��[�m����k�0�j�e�d�*�|R�}��T�<A�����&�r�.Z1쟋�,je�^w_Ǖf�H�(� ]B�rP�.8e���i>��`�����f`>�+��F��de;��a�ա��@n��s�l�~�02�ܗ����w�X����w��Vm��� ��L��|~`��N� �2T�2�ؐJ^T_�	(��r��J6�����}����4)��g��{z��C�S�����;(�b���ܮL3s&������c�(i�\���u�=ߚ�+�FW������9h^7��n����E�Y����������L(\�=d�Ĵ{s)�����q�Od�X����L�mص��(H�NT4�Ct�M��|ca�r�3�#��",V!��X���5c<f5TS{B�j2�5z+S��yy�Q�?+zf�e�lRF��W���Ih]�p0p�=D4���9����{Dl�Us��(:j9��$�c�krA����Sf�}�sO�� ��񩵇�/������q
F�o��#7�V2��nC=K! ^�R/6�R���hj�.!��/���M�}kșnfO�װ�9��1"*R��80��@̲S4�vеc�NرS	�k��7#�u��"1;����4�9��B灓 �k�(��X���a)j�f��&��2K��p��n%R%�����"G3~�Z�����M�G��f�R+-sH�k#���[�%���q�u�kQ<���% F&�X�g����.i�h�>�J�KVYQ:ԕ��$�d\�|R��|�����.��j {�p�6Upmƙ���O�������c�y��SK�{>�VI�Q�j�H�L�N� ��Qw���z�~���b1WY�!����`w�Ld���ڐ)�0b��]M4t�W7���IP����{~��`y�o� ���ݲ"�R����s3�4w�&]�S]��@�zX�t�h�����\�$�#�!@���L�k�.�IF q(��j
8�L���=Da,��m�H��j���qi(���ٵ3TNڷӣ��z���D��p�?<Q_�&f_�K�9�e���w�N)C�Wh�j��@[;g�B?2�~5��G!ڵ �|��F�N��ZN(�-K�\v�K�`H�6N�z�@O��#���s�=3�P�yq�@].�0�^��S�� Ci�X΃F��.�'�=Y@��B��f.|��oM4�8n� -�f%�O��V2-��:E$���n��iu\q��0<Ͻ6o����:ɸy�RDԍ�K�v�I2����eV<���������=<Y~�:��}r�rc�[���:{���>Nm��\K���d��y?��K��O��NM�%�2?�R����}�r	�f��=��d"v���W�D)SlEj!%� �D�>VAb�ʆ�TY6��Ǜ��l�f�>�O
<��c�/�$��٢#��/٩t]���v �'Q���[Ol�_Pj���2׏6��t3�%�-��W����Y&iM��´ �wO�P�$o�m:ed��+�Ddz�X�b������A�?wW(�
���7A�)r�(Y ��\N�\G�Ꝭg�ʖ����}W���V���o�v�-Ѡl�h�ݣ���R��F�� �d�W����g��H�&���y���[��:���(��	���)�֟��],�h�[u�ɬKo�K�܃P
M��BjMCUU��Wx����50�}�*F,X�m��_<�p�gʉ��Ý|F��7�i����Bm<��ˊh�9�(���#�ls���W΢!� ���O�t��R`R�u���m���F��,R���A�1Y6[fe[���|4җ!�s���.�Q(�Q/�bde�o׈�w�_��j
�(`J��y��{h�a�;�⅊�% ����s"q���YB#���b�z�����_�� ��tծ�5�j��t�Ƅ��]�g�-,~�ܮ�P7=_��Ӧ���-ƃWz<E�J�cB2�!�wd��(��)�ԩy�~F��2ks��g�P�;8�����o�Gb������	B����l�TuF��G����V�|S}��ūe�1��i�Xbo�A�M#޹������s���[�2�Ҙnaq��'22ɪv�楩�򛘁�����u7nq�S���)�4�=w���������^���:RΜ?�����ҵ��NG��i�@����Eah���;L��fV�
�%�`��q�j)�a�U��v�����-=�,B�����e`8n'h��vA�`�M����&$ľ
>RmW���'�㽼T�
���L���t����#)3�WG��K����pz�ȾKc�O��v�Y��<���a��,ܔ��af��Y͸����O��j��m{r���N�l��1�X��e9s?����?@��x)��&-T�����u4�$Y��;tL"���	���ȑ䜮I��^����AuR+`�+��緧?\�	��f�6�`�i�v�l�_��r��U}�&��Ķ��^_��BnF}�X��P�j&�����s2�����]���h���Y/m��S�uh�k��?���}?��P�r�'x�l�[�m$�0�7�v�HoLC/yQ���3�d�@�5�/Ȕ(�<̛G+��p�����gD"?� @�Oz�J�z�gW�L߽4+�P`�KF~,�o�նk��'��O���h�Ph��H���'��:Az�I�H.q�f	��ȠI0D�:�g��(<@���y�^�����Į�N\!p�6�E�)�NiO�2�7��Q��B�PjS�g*�kv)}~@��,��r���$�$l��+�඘5�=�>��W�T����=������$�IM*ƹ$�%Cr��.3j�sƕ��pH��J�<8,d cϮE3/�Z(�f�k7bc�\gu{��	H�]���8��B0|��m]H���6�M�!XA^�>���RDB �w��Y�W�V��_�q�e�2���'�jE}�D��M�o��L�G�7$ד���Ra��`bvs���9j�<4���%��֚52Dg�`�x ����Y�uu���	9���H��Q�?���x�����5�W+

��}U��D[����\`Q�9�)�yR�mScR�(�� ����kB��j&K5<��4�}X�,��N��CF�j��ڔ1��pP� ޓ�������7�0N$�9MP�E��U/��B��"Xp�"b��UC?'g'�c��%��*��V��860|�5� ǚ�¸�¤'��nj�T��U`?F���w��5~�Ж�����V��D��q��7���-���;�F�]&O����g�m�-���uf`賦W�2�l#Cm��h��̽�����hø7o�U2�ώ/�m�X��6�S�#�Md94'T�7����ܤsc$��u�O�ZKP�p��$�#Ci�>�hHC>FȖ�(��F,��6e���B*zd�!}���
�K<�F�7>2S��;��3w�hNw8��Bʙ[�Μ�ߒ����e��l`\��b�*U9ج��3�h#��_�h�8��#�9���vp.)��o����h�K��F*���yA�9�F�7Q�v��3�g!���Jp�(X�G`n�.��E��r���Ie2��Q���8����*~4��L�$p�`�秢^�3�1~WQGEVa��4�+e���S��2��P���~iG�l�n�[�+xâ�:��J�����:VR<Q�pE/�~D�2>���f(J?��~%k�냨+��:�\ձ@)������ת>�\���EuKJǞ�]�3���h��T�9.���{Lj!zr���0Tah�����s��/��dڪ�C�*��	������9�ɵ��I��w��(o_N	�%p�0��/�����i��-�����&��H"w3�[g)j����k��5�qul�Ѩ�^0��n��������F�x�J͹�#�Ї���fdRm�.as��e���c�W����a�~��Ge��.Q{br`�8b�=��c���'L��Z �໵�n���2i��#͖��U�T��r��.SY��J!&�N�?�����7�qJ�wp�.x:#�Ȣ��`bIL���y}]���K��"�F��*h�.���.��D�*�ؗBp�G��:� 2}��B)� -Ϟ�ZܲK��F�Ɗ��k��_=�b�AF?P��0] 9e$Fn�J�lWy��Dt5+1AHߧ�r�lre.C8⡉�ܒ�.���]IP�g:\�4��?��(B$#�S<��D�w?�~�Q�̈�8'��]�6��Pt���W�J�F�<bu�U����'�+P��0��W5�����4%����Q��]����:���S��3U���?5���˧9)���Y�� r�T���Y����Z��ʹ��Q7�Q�160�ƍ�>�@V�#j`�2��N���|ix"��2}��J�ibo��܈m��z�^tcu��!�	F��+Hay�r�j��@����]�y��:\[b�����Ǻ�F�t1,�בMb��pP�aH�.��v
�C�9ӹ�!�k�]iD4���³�^<z��t�o��8'C����(�?)Z��闛�3��!��p�|��כ�2{z�h
�]��o�\�n�ήS?v�����t�i\Ga]��JFT�s��j�R �P)�鸗�a[��e47�4c�Fe;q�'�eE��޴nX3��#�[���y�ߚiZ�>�����/Q��Q܊<�ɞ���j��ّ��h�"�-vƣM����������/�,�Yq�*7_����Y������1Lz�H��j�{]��J�u]*��iXQDهX
�7�9`جkuD��x!�����FT���h4Z����DSW�%yx�Fq�e}CPCU,�cO�ߑG��SQ��ڻה�t`x�|���A.<��1\y&DY90�A���T�������`�Q�r��pv@_�F�w�>F��pq�F��?�3�*�]�(Z�P@�B0�&�V-����39��"��CZd�6��3o�ݒK-�Md���m���*W�$vF��{ۻ��-��m�f��-�F��y%Ѯ�ӋKxiD�a��4QG��t)F0{��������nB�Ĭ�[\�e��	��YC\���NN3��#����j�`����~]��xf�d�	p�vF��'�j
�嚙�KKE��Lg[��uN�D���w֠�v���U�k}p�i�,E�8���JZ%׈/����q��LEb��	�%y<.�$��ŝ��a�rd�y�|��1$>�X�5�5�B_��6n�Q����H�5��H�lq�C�a��u�?J����YN�J�Q]8����D���+��^��d�
m����-5�Z��0��[�g6�*4sݣ M/����zh8�0�{6�K�1�U�&E.��y�,��;#0��"]��sT��E~�[�:��f�U�WT�>#ӹ��v{�P5�}�N�2���n�7M��ck�׳�2�J��x_P\�r�sZݯ�z#L¢�H���-�
�.;�͏naE$�g��ԛ#��*o\����;��2y'Z(MO��Nd�i��Yk��RL=�3�"
%�;u�V&���>:���":�M��Q�P��1<��ᕸ��%�OR{:�\��EQ�L�=/h�H:t���~�����t�:Q<�Ĝ ����	[T����cG2ZW�_�wYv��4#ݷi���o��RX�+�@PYׯLP.��8L�Gj�8�j�+��rr*a
Z2�3uh(�hL�)C���?D.�LύMg��&!�����w�d�=�3�aAX��ٲ\��݅��~��]��H�������_���<��+�x�?ݸ�͏�A!�:��̡t1,��z_s���$g#fsX��TQά��/ �V{F�9X�nX��a�D�m���~�҆q(2�?y�t�U"��Q��8�������*~�����?;��}�1>&�����x�o!9lĆ/=R0^-�������K�;���G��0�:#K��~�cwL�~��=xb��M�'J���d��-�eͨ��(�ע�~�'��E׼S=��̈́(�=�I��1��z�Q[��0�s�3��v:��.�xZf��V�܊m��62��Y\s��W"2��A��iC��"� 3_�Z����3su�8����w�E`g<���3���h�'a0h��@q߄������2�"֜ښ��J�b���KW�ζ׻�} 1˼a�Vbs*k�H��^�l�M(��*���������h�o�����qA���жy��=3a9�Ta���âDM���ZNGvD+b`�;Ko���-�3�R�/P����f��ӧ;7�Һ-a~�=���e���)ݗ!bF|l��"-��u�tP_�'�hԗ�>&��	u+W�gTp�e76�8��b:���[E�T��Wk�����.	�8K86�0��z�2+~(' pv����,�Wȃ�sM��<��+RL`�q���s�2Dq9:�cP�[�O���#�:��h�|>|�͉a�}O�C8�c(��S](�U�E�~�#�����74��N>����)>�&�E�|cT�R�a��p2 ݕ΄����� �?�-*J^�=�72�����۩��BP>:Q�Ԧ����������̂��o�����ى�3��UE>0��I?w�G�,�h�����v����u��奺kb^^3i1�(,s܅�N��))WZ�.x�H��EL;�2?"������]a����A}�2= �ԃ�|���I.��E�`s�w�vM����e���F�q�)��mq��f�okze���'�Hi�+;qV����=D��H?ZУ�<�������~�>GZ!�A}�vC�6� ��Vd��~z�X�f� r�M��I_�[��mۧ$x������
��ɽ�*v �K\��^���>~+�6�8<�6>g��yE!~{%��E�?����loNz��ms7JF�*U������O�1@�̅*���kl�������z��B��C}�OYw��(v��O��W��'Kzr����k����ń� N��%j'#ɩz�Ed�*�,��9$�>�FaZ�	��qO��e�-��P�M���9o��yezM��OMiL��o�	�۾N��X!Ñ=9Tc�����MVI�_��K���Z��']�e�zZq��O���.�������%ɛ���.�����vk09S邚���{�-�*��˙V-�@�qB�;*�~cxI6&@OG�Nwvv���j�b~�H;7�:;�ҀKt��v:R��5_����l��*;ky5C��u5a������b�Ȏ�@��D/��vﯨ��m��w�I#��r�yZ߸Swr�H��s�n������ɦH�����oWL Y2�GDڦ�P�=ԉ�U��F�B0�#1�}cm�R�+��%*o+{&�As��˯�<�}x(�[�Z�r��-ܿP"�?�C�Z�l��j�P ����Y��:K�w�Q�B�����	�%1D��|_�MW�3M�Ku�/R�NCKWv�ޘY�~���Gf��6��P��i6\2��Hw��� z.雔����_"y��o�l��*�O_���Blkcpy�"P�N�Ө�V!B�=�j�*1X(8vq!<�EYJ7��Z�Ӟ:��i�Ro[�
�ⷜ�Y`�
���y�A��!�.�ze�.}����V
1��S���|�^��om���SnZC1���D�2����p��䜎鏳`"�e�,J��-9&<B�Q���*�e3L:��I������`_$qNɫ
�CR4h *Y�hûf�ډ:�����!��:��\��hh�}Fݲg�T��Nm<�����X��U4��5��<����́���6�mU����Yoa(��r���"�1�M��7	ɦB����Uq���l4w����jK �7����"s{� ����2��
-�FE�ip �J���r+/t
u���)����/��������x�8pa����J�`�0�o"�C�=�%~�E2�_+(�N��6���r/����L^7�U*\��;�j�["�,e��6�8ǭ��9vY�&�2E����L:�$�lG����a��CGW���]�4Ź��E$çnQ^O�1ᮛ/��G�~Ӹ+G�RK�x<,�b8XO�/�,��{��˴u��M�Mc-ݽG\�s�?����=҆��E��A�'�<�p�%�'�x�^L���@���d`m$/�9dv�G*W?Dˮ/����j�;��Xf!���1 �jU�K��l��8��aZ�wL�m3ј̫�P=���v��8lx~Sm�{��n��)E"����.n�j��O�
J���'E�D��߯F�#�uH{��fm�@֣e����v�e��j�?=��6����V�$Q5���#�����%Ꝕ�J/��nՂ,A��{2�3=}˪�)~b�J���GV�)�(hh A0�W�_�n0Ɛ]���s��J�F!���Zu����<�hlw���iDZZ��Y���fHb,�¨"a3����x�y��/f��oW(s7�SLh�w&"$kq�84���?MB+-��G3��kf�Ș �\H�]U�Q^@��5�ip`���D���l�Wz_��69��;,[`m��!d;?8e^���HUqX���t]����j�&2A��>}���ܚ�Q�}Koq�,D\ims�˄�~���b8T�Lj�[wZ�L�ż������Rڍ'|d+�~�;�c����ῘZ-݁(0�P~F'�&7�@��Id ��fM��!��+��-%j��('\��}�iW,�<����.�"�U��X�_�oە�iA�����I 4y%�[��"p��*k��0X�x�ь���Պ�v�Z�H�<B\��˾G[F+9 ���] [dMP'��Q|�+N�d�9�Y��f�S=�YE����\��h�W�5`
1���?�h�1����y������d� �8;�~hօ=��T!�}�`� ��'kJ⛬���/2jR�~���N���xF��q�U#J;"��%�1J�g�#a�W~��CH��M;�=~��_䤊��Jœ�U�"��B��sE�4�
���U�j����;��5<q?���Am�ӄ�&O��ᅝ	�/���r�[x���x����a#(����a7��h�=Ĩ+�w��O���*G����O����zb�k�+��j�}M�G�g�{�A?�>:<��w�@x�s���a�U"y�����D{.�p���+%-�q}7uO��^���O��
�s��H�p .e���Q�Lv(�a��<�Q���}V�6�{�#p��u��߾��9a��H��^�-�;�
#s8��;7��%3�^���*wO�=ȩ312A��A��$_)�Q`e-�)0.�=����>&$�y�ֺV7i	)dewL`Ó�'�x��|��鄰�<��*��d����i���ַ'�^��3j�S��"�Vcq��yI9�N�]�j���sM�����̏N#I�E�@ѷ�s�� �__�0���x���w[�գ��,�M����K��WU�#v?��޴�H$,�X�_��7������LO	��l���ufgYF�/$�l�x���ɧvt�S���M�
��Q�a�4c���Ll�m� �+�Cg��u3�2�o���J�V���+%ſ':�с���K��M!rپ";��u���@��Uiti�q����R�
��L�3���jm4�$��S�*�P`Y^"{�����?�eqA|LJ#A����R5���cz��jE�t�p�[����&o� ��F+9T;��� Oƌ���j �p����H�,]7L�6�loF[cZ�`e��l�U�_�NmaTd;�k��g5X��!�p��:�4;�<`u61�I����!���0�1f��3��������u���({̙�������N��k�:o��g�)!rLT�Ǥ2�'�88���E{DT�~ik���1��:�q���9뙇�x6o2V
�sώ3_z}��0��_�kΚ�8�]sie�`���i`�ѹ��U�kz���9�/X޻�)q��'�hR��r!f��g
����AcP,؇/)�㘫�oX娪��{�Z։����ЋO5�f�e]�����  ~�J���T�����34���}�#Y�~E(Hz��𳑟 ��;��e+��;5�:�΂ajG�4o�!��s�ƿx�]b�F"���@�-�ձ�ߓ�Y�����ԇ�O[�E'��}���X�Ǌ����CԒ#Y��6_8 ��8^��{��w��ҫ=��Wii�33<���F�<�Y�	�1�^�1�,�M��L,w�z�?�{���j{~�y��J�y�P�{���v�ĕ[���n�ze����\�(+�{k�0at2U�����X��Y�`w���%�D��l+��� #�8��ܟ�9^ڳȟ��+���C�Y��U��sm|�vU��9��D|P�oDa��p}Ƽ��CR��"��<"߉Sy�ic��0�OQ��q����Sg�'��$C�(����;fsu>n�.zG1�%ғ�@DpCn����>U��l��L�ҟ�7�gF�� N=�8R����ith��3����m��cӗ���$�e.U�q�l�|��=w��e��+�B�%?��C��*�f"T5r�˛H]C�V�:��ϗ�PW���h!UH�����bl��A��!Hl�4�[��#ű�n�J�.N�u�Y��u�snF�'�zb����p�� %�����#�X��j��5{f�=�j\+�$O������f��K ���(�7�eMD���`IZE����(���u�	�Q9)I`<�� ���Z���ڳ�G�/`�tk)5��O��2�2��D���Jm���O@�;����L���=��0Ǹ�rSDx���}�������2�PK�	�6k�J�֩G:�.�%G�$�kLp�V�J7@cw�Z�qkp���$�~�ܧ�f��ƛE Q ����#W{�Dx�v���5�*���9sց��I�)}�;��+�BX��q����6��s�O������d�����`�$C7��:G��E���P1�X�TD-f��=#RL�=[�"AT�����f2��6�K�\�����4��IE9��X���ȉ��
ᐘr�n�Ս/�ӟ��ӎ�"<��ksq�6�c?i���J':q��Ӫ^
?���(6[v�m�����]���%�$80���]K2�����\���ϛ�{r�8�f��ڪkj�l/,��M��$C�
����y��1P5?MA�]�*�|�?���O��BLj���v��$|�d�h&x�f����8c��?�K�$	�8��L�����O�,���C͕_� ���`���iKW���=M�d����$Z�^�e�~n��D�0�\�)ҷ�)�A��B��Z��\,��W�dT��z��%�ض8��ʩ�}cM�� ��	+8OI�W<��@� J�'��4B�􈺒hK�~�� 8I��B���h���&b���z
�y�:��A[77���ze�N��eǔV��5��8�#��q�龽�jOY\櫿��4�d�2�$x�jt3��!�D��)n�4��|��հ���wv	���34� ��Cl��r�˲����^P������:ԕ:���xQ��Riܔ_�B���tȝȜ����ј䊀�撏��A��És3������4M0�J�w����C�t�{�8&]PF�5_ԃj�~4���L%)���xZ�����m�Q;B��x<t�p�s����ʠ�>^��J�2I���՛�M-b�Bщk�q�9Aws#7�t�����'��������_%ͦƉ�m�8���Ֆ=EX�A�>=�~���	{N�8̿4e���u�a���i8�ܵԾ�n�dx�z�p{�{{�tE
�P��)��2����4���(TH,.9�}b&�aZ�� ���'��Qo��6�BO�3]�~Ե&��R��kۍI�h�W/�'hd,rbO0.Z�3�wG;�� �Ւ�4���ҙ�!�j?P�$ҽ�OU��ǹ_�Z`iP ������k�'����&}7��r�ò�Dk]vת&�SjΑ)��iN]!��{�ma�|{/�ͻLEg*�l�?����� [��(� B��=C`�:��1�����%���F��Y�=�`2�f�W��7�P5Ѝ]{V	�f�v��K�>�v���U�j���	��T9jPK�4�g

�&��k��\�8��M2����D��֑4�<ŘΧz�O�Jd�R��զ�c�B�^I
w��gT�!(�ڇḢ���Լ��O߲�S/�>$���m�dCW8�A,���
��.#�kN�=��~<�f�#E�X`ă���iG{�o^��~22Z{&)1��k��2����~�5rt=K���Tld��228H��ܲ�o�x`=��8UC�_Y����id�5���YA��
�b�S�����+k{�Kt��I�������}�4�Ν�r���b��vX��r���S�yYVE���%������X2�Ǒ��}A_�$2W���?�_�����]?��	���V|o`�YT[�}�^Ԡ��g��M��!M=q(�wp�ϧ�_FaQ�}���ηn�MN�a� �f ���H�Ѝ��!�������
���g���[�\��辌*�X��`�xnX�ޱ���-gj08�IRҺ�`�ܜB����c�J����"VH���3�1"������錰MmhI�'��þ\!���ؘ�h�q8�1�HC�-��ѣz��UmɆy@����R���>��b����N�HW,ڵ�/�'���߲s����/q6��.�������(��mm���K�}%�����<o@|�x���٦I�F��.�����{ն�l�%��:<�z5
�����3'@�I&F�D�"_q�2Δqw���t6n��\��:hz���r2��R73�n��2�X>��� v�:J��$;͈;�8���w�{$=����1�&���� ��2��ϫ���m�1:�6��*���;	(K���,?�Q�P�Irs�@<�G��(.ONS�s�v���G�I6��q���5�CjrAG0��n_����w�5��r/4����0��o��;���	o��>�k3��E���������Y,s��E��ǫ��P���o�K�43���z������&�F�:*�RNQ��i.�dȨ�����.�#�wi�D\yݕ��W�؈eU~���͗���s%�f}=v��\лP:�j88q��M9S��8(��f�ֳ�2�:O��^�_oF�/��5��t�(���a+���F��Đ��a%ڔ�|"U\��C5ި/ѓ61uO����
DvH���0��ߒ�%Y}E�B�tSI��έ��F��]�.�����ݦ�Bol���_ �B��RF[~<��櫄�h��N�e�:w�i#
Bz����&Hb��Z���Gy�=��Z��y6\�Q[;.G��38�w�*��5�=�2��4��14{����y�Nﷹ�g��I?Z�̣��aw�m8�ϧFГʿԃڭ���{�_]7J<�P�7�;�ŴU�����妄����RF[�o�c����
�Vc�ǂ��2��U?��.�"��_ =�82=STY�IR7���U�f��bu>����Et.{�>&�v���䱬�(��*�
D$'��.4�cC.�8��È��H}�a�u��T}5�`d��wM^g��x#V��.!���0�mh��="�!��O��L(���v�~�^���c(��tL�v�|!io>5���Ԃqr`�＃�p�bZ�!d�q�	"�Q��@t�J�d-���ZLjt>2(�"	U���g��\ۋ�א��7��S͚����5*����u����9w7eD�Ě!�B�X_�l"�I��z�m��.wa��H�b�*�&��ʽ2Z��+N[��/�*��w��Nd"*1���0��OبXy�4�aǆ8�܅��]������\Y]a��?��Me�<Ŋ�\Q����2 p
�By*1[��1�HX����'���ߌ#Q��7�?}=��@"�v�&���=�#�K�`_C-�f���6E�A��[.!(�w���|�RǗʣ���_4�?d�#C�j�ဂ.d\��-��t�HL���*����(:���i�3/�����Մk �;�g��j.s�/�It�*��Ɇd�m��LO����3z�!��4�ۨԙ�)�3��"�T���GV$z��Ec�=g���\���n�_z��i5�j��.}[Z��FN�X��p#w�!��<^��`�ە�������B)������D��+�0�"
�M�O���d �*���:�f��ಇ��l�}�$�@`�\�(����B�2!j$`v����;z �1������S&1}}�P؋��� L=+�=8��^Vr-���q�wZ���ƣ�(��^�	8�dbr����Bx�+ҥS��)�BR�ƝP;K=��� �4\J�P� ����	���
0�W0���^�E~��v)�MYC^}�[�Cs�����\�ʫ6T:\n�࿑�-�����F��ij�*�R�@�Q�1���?����k��Gz�/���^�'��$�x���s7�TG�%�p��2�D{H�w�ϻ��h���O���,�C�%�TB�*f�*|~G�pvP$�d����I)��q��˭��=����hwM��v�ªYbj�JW���E���>�?+;F�7�~Ա�����_[>dWi�؎":����,RMn�=���������֎JeZ���C��
g(��#.ʟD;M��O}> g���C(�1��|�2�Wm�l��G���A?H/�/���v	5��{���w�������D9Z�?���Frol��Q��ُ`-�4':)��]J�B"�H�{U�M�	'AԄ>S��Z5uՃH��X��,^㟆�
��.g���c��`�zm�Si7�jeW�������@RT�BL�ND���y����|!s�m��O���ޫ7�Y��LV�I'��U���"��N�"fx�@��I"V9��(��{M.��E1�v[���&�g��[�n�{h8�=b��ϋ��><q9�o=��<�Vݡ������dg���f��("����e��g��ť�W����>��i�e�w7�Rհa��E�"c[�� �x�fN�h�hPე
N�d�҅��U����g�!��1�j��Hߘ�cS��5y�2�:w�Ҏ�;���@�{���0<G�T��n����W��z�Q����/�jL�Z� t�^&Z3��u �ۻ��0��KX��B�R~BB�����C2̿��?�	m����N4jW�1�[ΤU�j~Z�L�g��.�����k]���#�6��ّ�/�
�H��.]ZgkϡV�)t\�|x�ЛN�Li�����J~�7�Ϧ_?��Ѱ�J�i�ruz�^�ϕ���' ��g�X��/e��ƶ����#w�[�.ϏԟJO�W^��.�D��Y�9aǶ��^f-�Sf��$�
�h�p^���t޵+Zq���k�	�0��J���8�nE$F��ٜ�7L����v Y�o{d��:6��HQEy�P����Z���>���+���34�W,N��:m���BX��y�ed���\����=�1�%J����J��	 0+�lV�krT%��� 5�t͑3�.�&��ɚjG]�Z�9��r��V�Ń��,$<[�����~Lq�`��jD�~�CI�cV[X�;�˔;��*KM�= ���
S��d��,A�qڡ5j�����ھ}6��C�4u%��C�Ɔ-
z�����W6����s0���&����fYp�Q��'g�� ��K�.� ��J�Kb[�ˑ�����X��*m�7F�)�㦡Z;�e������#C�������鞅w}�P�C�� ��oKg�������L #�얛}"��(
xG��B:���dv|��#������M"�ү���K���C��������t7�����I�[(����|��O����0�PO�n�������
����m�<�Y9�b@���_�g
dv��Z<*��f�uv<v���-+���h��¹y�6��;aNDk��zu	�>hď:�;fh1�� X	�`4}�Rc]3��=�b��☼KB�q1�G���N�"~`"��j��WcY��n�)6��������33���E-,Ӳ�­�|l���|0 �;�U0\�yX�T�.6/�����<=4QZ�`���T�}��9��zD�����j����|V)��Q�N^��|�=|�䆚:[�߽"�*����o��&�Xz�ʠ�������0e�7q5��(��R��l��c��^.`�U�H���FwA`��Xx6��e�,԰�e�BL��Ǽ�����ge�d`�"K��	^���`��,�/�w��)�9=.�?O|=lD��;�|��8�?	�ulY�`��]qr���4Wi��{ژy��%���B�e_�ζ���_����$G�8TX\��-�ƚ�é��Jp���C��(��r��o�uV N�in�̻��Y�
���ċ�fy�c �Y緀7�%ΠVQ(�"��mK>�3�l�����[7����#��J�m#��2�0�qP�7FjJ��DC�<����3��ELƁF�C
�E��-���H��E]�8�pBm�����;���� �.�`������I+��D�a`��c�s��i��/?��#��@޻�eUn*�fnZ^���;L1�y�e�i�x���:�4��I٪ג��Ӂ={����)�b|�=k`�/i~�K���7VK`fqM���~����Z�A�jP�� ��5���^���3h#��2�������^����5c���"�%�}ɩ�@���l�S�$M��=C/&��A\�*�=b-m(����GԟDzh|`��$E�\�<�g���&�ͣ%�e��-�#`l��	�"�<KB�hŎ<��Ɠ�T����O3�9��]��qf��K�@�GU��J<��?������:���b�
�i���M��%�Wa0����QG�����d���E����F+v�:I&��JW���V�� M�4���(c���ĕ��d8�:az�6s!u���Xpۍ��.� 3y�ZT���Ӓh6��0pS�P�u��i�C+�w�(;ven���]��w�3�hW�����Sy�XHޏ���=(P_�jk�V���_�q���,���g�3��WjoTꭎ�Qԧ~�II�>A��G��������k��
�h;�̯b�X܆d%e�g�Y�}�7��&�a�.'����s�n!=m8H�tiIɰ�C~x�wsHQ2�J��˗�h��1�,W��?m�p��`�	����y��i��;�H���� ˿qwV�X���b��������:]�\	X2!5��:W&�L N_�L3{���_t�3�m|FN��A��(��X&���a!�B�%��i�?Cܽx��ި��Wĥ��c!*@�艀������Ѩ4�mK����M����@R�cB��*��ϫ��j�*�5���v�tԻ\&me�1=��?�L�Gt��u@�h�o���4� F�	�J��)���6~IZ��7R�N��Ӳ�g��1L�UT�N?�:W�:K��u(0TM�Oq_vh��S�$��uHI�[,F3j��ʏ�NXR6)��ر�c�*�z^�4˧��<�(я������֓�c�F�����M�V@'�p,@��{wg)�ӶM{<�l�K�\���*��Y��M�����7,�<4�З͒�H�A�2J�J����$��=Cz��$Ox��!+5G|�h��7�K�HB;��s���(�B��DK�$�υ�/~�לjz��f��>�@�����ݽ�U�FD�Z�G��<�+�� 쭜���!]�O��s[��%"Ca�5�6���VxM��d�2"�b�o�-#��Y 5��F�+��u���
V�%��T���������$���)��,��s�@�P��jT}��ߘ����F~��4S*�N<��}��,5tJ����⯐���mZ�H�@5����l�Z^��R���=�Abr�����*��y�[���'W���q��4�[?�ܬ�b�Y��M��ٖ��Ǫ������$��%]�|�k�
��|�_�re�C[::�]�:�����ړa��si�A�w���pQ)�n&Vn� ���VáCH��ֿS;��;+ɏ��󉲃Ċd�WK��Y�#�����:�T]y��3%�F+����~�k=Ϣϰ5Ki��JOXT�j5��1�>E	�ڴ79�A�������s�T�;�{t���-	L�O]�C�q�w�L]��I�� �K����@���ާ?e�U ��{��ٽ#��⓹��-t16��⎖�ys�x���y��A�����SK�a����xb�L��LbD�^BE�KU��L�'�	�r����(Xt�x��=3�$F���nY�NN����\���*|߇� ��������*�n6����A�]���]i>̩U�}�N *�����1�86�)�ڎF����?�bsߚy��lj�g)r�Rqր�
��LFQ*Ј��wo����>�I'%�"�O���A�Ҥ�[V�����..�� `��-�����O���w���.�}�%��4H�T�B�Ί�W���]�t��.��"1Meq=�JdmAm]��մ�x�8��*�X�����?#�6#��.��r4N<h�FQU�yB�u\b��)������b�p�ܲ��P�+dG��;��r��=�>:'w��Î+���k!i�)>�	��#��D���ĿT��'����|�e����R�~��Ɗ�Eɀ�:/���$�l��!U���K[�۾���5K~-]C��BC�D���%��%�`�c��{���k�i�j����68Wvs�RJ��lv��"�5�Ŀ��Y�SV*�n���bbF��Cc�O�q1�
4t��h��*$�V݃'��t�v6��3��F��3�cV�t�R�o���B�-�=��g(Z��=l"R�[h	ߢO�Ұ^ښD���OG[����]��-ߞY�x�Ɯ�}lF )��̨��.���B56!��-�S94+!���P�?fgN:	���f�(0�����թC������W^1H���{��ׄ��t�䥴�]_�[ߵ��}*R�7�F�dC
M{�űH�
�5���H��)�ܱ��V����ٝ�B)�*��-W�!�\"��x�{S/����w�Ro)��+ݖ��^���cK�⊄@�㥞�5�L��~F��=�h��X�����T�^�K���qKEJ�<(���	$��T$j��Z�PA%<h�V�P�cv��{���c��=�Ru�bp��>;[ԙ�)�3ϊZ"���F���?������yfYԺ[|���xd�"���41?��?���:VR'+3�1���$1L�ڒ4'�iw-�~^`�C���N����B<G�ec>�S�5�Lw����~�;��J���y��J7z�*��	��)�1QE*+#�P�A��/�n Y�❵6췙X�Y#��{O�$";���^Ds3mf��&��1� >����)ѯ���nJ���al�QJr<!?����й�@��:�<�m~d�6]	��\W���Qt�c����RMV��w��{K�{��ʕVkK�F|O��o2N�(; �"���u18�̀��gs½)�ߘ���"8f,E�O\�7�q������8�:�-��ęHl�.3-9Q�}�,tWN�̘B���E��L�fp8}<p h���D$O�5�̫�7ٛ��s�+]�"�3E�2ўuϾ�S��Q�n�w��{���^8��/�Hk=���h�AJ�YZt�V��,��*g����B�[n��~"��s���9��y���m���o��l�w��Sϙ����*��=��dB��&�<���I��1:fF���|4��B��S5l!��MX�Ӓ��Ҕ�2�B����]�;�/*��m4:����f,�l�S0�N�o�$������}5���DD����{�(;5�æ���l���-�sͿ���-�"=�S5��dc{#V@A�cՐ�����+W����������x��N7zA�͒�O跄�/e#��4>p,�r\9B1s����=6���Q�����SR���g];��S��,?xa�3�W��O��k�<Є�?���q�!�q\�31�N���S���J�lP�Qj�}���YYz|���!NU/ʁ��������1H����,��0�o9��n	��>jq��8_�o-0��y����Z^<]tF��b�j��wl�a�E��A��cg:����r�-%x3�1����n����Vgn���]X�k$z�{~��
!ڼ�\���sQΰ���u{�? :�y���>H�y�w��쓔D�~���n�h�g�(��j+��%��~{FjoK>�24���e�F�R�4��v�1�a��
�ڇO ��B�/7uv:�:~.�#5?��_�(�$��5�~��~�6��;6��I�0��ʈP������Q���
�{κ^�Xmf
Km9 ]�;����)6�:\;#�OԀ��_x���E1k�a~�P�9N�3>Z١^��X����]#�/<�u+���ke �?}�OY��0��`hb�y��4�;���c���!�孕"������V�M�gPk�փP�3,u��р�����6�_y�e����svǕU��;'Yd����0���=�V�k�} �P^!ݤ�����W3�"��A�*���	���2���۰���
*(]ou��iԫ�MO|�v�����4�i=��J ?�̕����ۄ@y���yL��xt���$beF~�l�)�x_�����'�H�b��Ϋg]�����on���h����}z���2���C��!@ɷߢX3��5�3�Oc��t�6���Z�ľ2���D�N6��6�eJ��c��!�[�JZ	�m��"�w����`�@���J?���ji�ͧU�����KwJ�bBl��E|L	N�t���$N�Sw��LIA�nO���7V��1�f��|�9U��/���|�=��.�y��(���K����~��U	Z�
�1O��`O�.��+��0P�T۾�`[�7���g`�o9���[��/GQGwW�Y;b��Uk�#:@�j�?���g2����7�na�t];G�WX��`R��	�Q�l�(������=��l6�1�P�;����ʸ�<�=�^�����;(���؈��nYc��vPa�ENR�ȻiNu~�f3IY�m����j��]�s +�֎���#��l¦��wf3���E��F�5y�͎�Af���3��+�''��;�˪���|�
�/?�hixKB�c) ��<H8;q��*|Ҷ��ԁ��I�)�a�b|�å���p�����?�2 e#
YG��#�h+�*%g!`i���W����Ґl��m�_�+ј��K��\ek�9a)�hA�	�yh"�3��U3����^�G�E�ZS�BsE�g�}��re.�\�nӑ�Jw>/)��OF�Iy�:U|,�h����E����(�|�%� E7S�����*��\\ӒO��/�5����m���N�?�	������,k���iJ����㿧+�1��!���2���B<k�{2��<eI��ǭ����9��9�P���9(�9 �=PBX��������ᖆ�^�nX-�$8�d�̣��Ah� ����0�O6�p&`5*O&�;����e�| �\c#x�6�����&�9y'�b블�wًt��τ���ū��^Q-�a������pQ�}�k<�k�K����P�*��V9g��X����ݑ@���Вh5��)>��P���ޔY�1���|"�Ta���7ʙ*��(c�ɟ�ut(�Fd`TJ̃�i	j^,J�)���@$��{B\g��5�Ϧ߁IzA�O�8eg���=��$��d��
Z��Q��K'Z�K��H,���m��8E�w3;-�ڤ��v��j�Am0iSW���7dB�ۦ�EB�D��K��o���Q#�t�O{��@�jR�Sv�� �9��.3�:d`@�Ѯa���;~���Y���}�ֳ��/�	lw��TJrۚ�*�E.�;@�x��8Ȳ6�X5���̵o�x�F=�o32�n�Q̨/~�ū�~��R�I�F������C�cu���~Ub,�nZDG^y���M�o����Y�'�c�� �\ԕ���&�������y�o�BaƁ<1t���׷��g|Dw�|sH�D`?��Jj���a�"NH����qy��h�o�ah]p�;���Taaݽ��?�nH2��Ǫ2�}����$*[8<Ё��8JȂV�������e�~aY-�zp��2�Ι(L�G4Ǚ���"!j�J���$�X����!9|��.h<���s%����˻Be^k�#�N�iZ���#&����by�y�AY� ���5��NB",�4zTA��H,u�!�9��\-B��^Q��
R��mV���i��CK�#Ô�N�"	H��4q_�h�D5 t�LK�g)�[yj�~�f���R"�綠�y�:�> �zx?K�i���s%X5���q�F�2�Q�;�ה�
�L`|s�-!������K��,�ߔ&3G��� ��&�78��[I/�h�}]�C Ɵ��K��
dRr���FZ��s�م���R�!~]�@x��y��v�_xPV�Cb4M�q������I|/��j�P����3tr�1#��,uf�Y7�Ja	yBOx{��|-^�^{���!�~�������h������W�K������a�'�';�+�37�Iq���,TB�-�J��%-���)�F?l��{�I�<��t��j*X���	l�����{1i�ăKk���ŷH����]$��0twy�}�p+�[Y�)�ͮ��b#"�g��P,pb������tѐ�Bᰲ�.�������.��"�?Ŋd�P�,���t�Wfh��R#_�hۄ%��ͮ�cX8���<%�6ԨR]-�W�9U���z*49�m'P����j�b?�2/x(j�9�|�d)k]�t�}8��G[�j�VzYݚ��Z���:Bצ�Әړ�K>G�l������yS�_�]��/�9ظ�;Q�t)B\k��w��o��&��Lf�����k�ȟh���K0Z�j�+R��ͼFl#F��	�S���h0�n�+�.�a��<�㾕���D���;E������G�Im���2��o��}������W���F��[U"�u��Lr��y:����b���������� ���O
5��1c�`�|��N&0�t:�s�{f��15/���=^ʧ��_T�����[Sm���.��<���X[H�k/o���l�Q5�[L�Β�M��e7z����!�wz5�E���BQ<E�aŋ�/��.fCvU�r���(�h�V�0��yF�9x�q��U���\��'�||���V�W&�4�T%\7����V1I;r\��T���5%��=�{An�gn.�:��z��pp�[@��έ�7� n	�F�=���LDJk��1����R6Oj-��>iW?O�(���ѭ���69��ens�F{`�[!/��!8������o�<����ִ���]�j���w?�@��/Dȇ��S�z٩�e֒̆���$�I�?פ�?�&۝�1 0+,m�A-y�u�������$�b�\U��,�+1VЖo�������Nl�~�}�����-f�����M��Ó@nXb�R=\�Bɻ?�?�B�������_�r�n�L�b��h���,�Y�'�y3������Pb8(��«~�_�b7+��r4 �c�g�2���S�>�s�ع	����HP&��%�e%��ުXe-.�>+��$����0����G��"�����/�y�j��O;_�C���k���&8
�cH<��c@R�%��5�&������_"�����nY8s#��FA��7����p\-����X:9馰���m\Ց�i�
q�y[s�Zv5\Z�K>�qѕ�<k�P[,+����ި��g� �gj-gw���1ǉv���j���{�Eb����*]����ƍ��0*��8��=��\�c�n+l��)3>��ڌ��;�2s���1E���y0Mk��9�|\��q�mg�.f�?;AOHo�k I�k����4$2hC+�� m����D�p�Ҧ>�Ψ�)^��n�K��OA�;���] S��ĕ��@�S�D�����>A=�\��zi��
}�ys��ۘ���^�&�����>�7��2zWBv6ォ�?��/v]e��.��+r]kk��%�n�p+�����@��.�2A��RH�'����ga��b��R3�)@5j��/���]�<J��M�r����U'���(*oP,�\�6�}��߮< ��c �����Z}���YY�4֔d��NTغ�oUCm&�t摦�E ��Ul�͂?	�d��� ����� -/��ȱv(�����Q�V�B��n��֘�tz�qV�9q
�'�<�Һ��;��/�z"��ep}������ةK��ڕ6R��P�Y��S��A%`����WPׁd�&x��O�y`y����ɠi�����I�,.�i��1z�0���f�snq7s��Э��ƕpߠ��B�#W�,�Bs�j)tV�q���A�!9�t3\;�� �v�}���#�qrv�ڸ"}B�z嗣�s.k ��.U�땨H_�ܸކ����dU<im�|N���lhl��Tld ����G�2c-��[e9r3o�����,R�b��yQ\���6
t�Ѝ����'3�$�r��v礑�[�]3�]�)s3>{����g����s�p�m��t�Aq����l8�MVo>��U���=��ӷ�i�U�R ��&����*-P��;$#y�'���Ȥ�
%�&a�ƃ�`�/%��v�Go5��zƅ@�ϋ���QX��W�#�_R���a�T����:�̆���jk�O�&��1ޙ *�;�����$���c��T������m�k6�����F _�������*�}ot�w>B,�K�5�a��OQ��ɞ�9_wMC�3rsc�#��!��Sw�o�\�V��ђ#_�6�?B���.���;}����r�{83p�q'�ڂ�Y����\a����T�䷫��8hL�>B��o,Yc-���:X�@&�gu*�䀡Ԩ���*8ՙ_5��m�8�}�d@Ʈ?{N�!W���9��������к~�_��۴��"�K�|�>cC<�ԫs��lˑ
������
؆z�ق��IU�c���p�������*�e��Uo}��E��><r�J�����]�(5:�e8)��O�	��#��J���9�5[�/���n]؋�����?M�'�$Y��l��DU�$_���,�Tү[��3���K�;�"Ò	���aĘ��.+�>��=:�yq��0��XP3��D݉r��|杰 �]8�����2O@�{NY��ckN�1G#�� �۱e�39����^��9s�PE@���������s<�
u���2G�s���6���n�( u��<ݎ�1ᤩ��.�H�T���-@�A�E��f!�0^��`Ĝ!�Ð��T�֛��꠩:���w��x��yqI�$e�~D��a^�}5l�X�ZR����g5��K�kWl}lr�ԃ��2���?�V??�ȵ�{}��M�p煂�'s �{��e��z�ߺ�b�`����q�P������~p�Q8�}�SK �-��ƞU�$��r�F��;t#�m��V��D�y��ʻ�_����7=�E>��.��R^�ZG��bbk��-{A�����Ե۵�h<z�SpȀ,g7�q#�R���&���� G�����FL]��
i��v�E6���90!�˂��ѫ�r�ʛ���B�5�3���L���>.��t	��{��9�ȏ6�\�q��X�ҭ�`��M�Q�i<��K9�wE�������(^�Z}�x�;=P�|nٰ�~ٲ�A:Lv��S����q�ckm�,��E^
(1��L��k�%���h�Ď�q'�k1���L2T�? ��H�%n"l*���I�b')ӧ��ز�L�f5�Hԛ��}w���ߪ�X�cj�L����+6l)���7����ӤV���JM��DX�1��x�5=�Y]���ϒ8q�e����q���H��}�!��ʁ�d=��cg�{!���'�R�w���r��u �x��{�b� ���ʋ�����g��u���������ݔνί�݁ۮtPߩ8a��[��7T��j6c�������G����CgA�=������u��-��^��g�