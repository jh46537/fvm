��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9M!@eW:�Po��+?A��ʢ�{�&{��JN�����]�V|ӪY��Q2��zU.S��f�AO�+�����9?T�>-�o�,Ƹa3[��VwB�gqZ���z�EC"�@p`Se\���� �3f,u�!|bG����K�Oi��Y��%������e�;�`�
{��g�<��`�7Wbo@��٤��Y,ZT�*t����g[�� ��g�w�!��Fp�b��=4F��'��~?n�H�Ͼ�?|�H�����K�/��`���0{��}�2�+����+NaC��Zg�L�l��C@K&���$)f^@.q	�wi�o�䪯����90�QiEo���~/[�mZN.�ޜ�ʨ:��w�Vʦ#�*�|�1�7��a�V"�j�$��I�j!������j�&AtAUa���s�}�}J���	�
 BiE���	��)LϿ:���٥����� ܮ�b��94�8�^Qnھ]N!�i˕ލ��pt�d�t��Y�a���9E�ܫ����9a�w��́n���ؓշB��@� 7]�r-U���Ph�PD��"�+="��/�� �Ȧ��L܂˰6+GX��=������U��g��#�J���|���K�e���^b{҂�#���#�����ܭ����2���������N����(�$X��_3����)��"�u~Ǘ�����j�dUb}8�H��T��c����X4h���>�=�'a����v�Ky�|�z��#�kh��ыsJ����(\��ez@��f6�vk�8��^��\Y[P3� ����ECNZ�)�5�?��P`(���P��D,��Hp~�=�b�,H�,^܇�Qn�����Z�̄����S1-��;��]����Ӂ�>��hK��H�t�l�6>y5�=>�w_"�7N+&�א=��[�i�okR�����%�x��a
�[R�O�+C4��M�_�X�V��q�F�������4m�����	�͒�h��5������i��RڂU�&�Ǽ0��ǽ�9[-+r|�$��ͨm�U͌i(���偧 ���a�Nt@C\a�ӮO��{��0w�W�� Q�*ܞ>�\c��ݦ^r��t�y���;�����aT�.�"�bR��4h @��A�]��K~�������2��'�����&�]/8��P]���u���Z ���R�]�.K��"�{S��I��`ƭB>`/Qp�dAK�jԨL	\�Q*R��~���R��5��|�;�uw�m�@��:�a-]��MH���g��$��HM�0r�A��C__�8���feˤ���y[�z7J%4���2Z
O��@GԀ���)�l��"n���:>,�a������d.Z]g~?���È�4IΑ�5��X�_��&�,����c�����˷A�,����!�=�cb�B��G�n٭�ݣԍ���$7c5��Ohu,���`@��0�Wm���I��,�8^p$๫��+/�4P�?�3i��X�P~��4�AO�*a�l����p�/�Y/�:\�:_��nw �%h�_�]�t� Ht�hB�/:ٚ���+i�Uʖ��
Θ�p�F�c�Q�[s�����g��9 �c�.8��u�P��F51��~���h�{N���������nۑ�+4_�ʑܕ���sJ�H����i`���&3����ߖCKg��s�����ḙn�;`�/�Ht��K�g�L��z7l��/���O�*ɰ�W� �7���a�C\�f�Y�S�F�R}�wL�$Bx�	�J�c��TJ`�e����H!�dHt�I�~����"�����wppe��Ppcv�]��M;S�q>�s�)����*�?���</A�i?��V>Np�?�+��E�� ���G�#�|ʄk��~���_�[S��<�3��s�&�,9��1�T��U���&���wL�&���>)�b�8��$~B���o\�a1�p�pB�z�B�x:��cPM�z�n��2tٟ�5Et���!��I���O]oV��E(0n>2P(U�'�����V��c�5�(|�b�)��d�X	C��|�U���"�}ھϫS#��ͤ�'ɬ��}3 �!!�:�~t���+(=�G�q<�O���>��:�Ѕ��hK��a�,�y�\��{O�Ӡ#WZ`C][�=A�8Pب���]�הly�	p1��!��:?�v~�i[W^}uI+��GG=�ػ֩�"[k'r,�'T��fn��^\ +M��M�t��ڐ�N��Q_�rM%�{�Z(���s�M���=�~<�BL<�L�0:����_�Ƽ>���lKwz�=굁G�J_��\´s9�nh��ā5M�"v�s��6�c�q.>�S��h����,�+���e��L,��R&ib?+)/�'D���U���`k�ޒ"�����M �ނIQ6/�k�8^���y���%B��J�S�5c?��E�� u�(A�E��O���,uw�32.�y���.��-��-���fX�Lc�:���.�w�*M"L�V9lm�WD�����J���@diM�]	�vn��m�Bg�2>��a�R��:]9�=��4�;�䭰*Ӵ�y�W@���5��a��±u���`o��$֙i�D��N��VQ���p�����>P�XLB�+���=~M���_7��^Y�'Rsoq���7�44A��v�5Er��NS��8I	r~����_�C�w���P�w�"�m[��� Q�=����a S��.`@����|�����x�m�\�n`�#�m��3ޥW̘���.�ok���M�͢�G����.�H@-�Ĕ&N���X�7T����/d��%��jY���,�O$b��4Z��Ji�{]�����sP��1����ۼx�#m���ҭ%�R�Y��>vge����1�%�v3lz0`�c���������U]Q9�6�rCi}��S��9��w䱪������r�X��3��� @L������:�x��z�ol�~�$P��3U�c�bL"���E����Ǉ�a����&��1���y�T��t���8�Y�F�5�ֶ�O��i��½'1�%>�'��|��quaw��a�Q�m��A����tz��	J؏�k��;zkB�TK7��Í�ˮ�I�ڭ��h/��i��:� �K7/eR��Z&"�/C�yj�خ\Z���P��Gi����)�d9�h�vC wJ�Xe�G@�8�H%�^�&W��ͨ.Q���p�Lk��̍$!F.9.y��*�����Npb.ե�����W��m�Ʀ �y����a5��Bmu��6��R>���'�6	�-���E�bR�$�5��
VQϮ�"�Li�R�1{>_�$%6Z%ѫ��%��L0�6c�6�����5�,.�(��m��#��љ�me9�_��-��ѡG��l�f|�2܋�S����_u�u���G��Dw�k�U�*2?[�u]�hg^p�"���Ä��9�|򍘫�$��K�G����2~S)�n�0���so�?B���c�����<6�S�j�x�S}�~�XG��R�%��9H��+2v�� t��d<ۘ"��@��(��?H;Jsuzҡ1DK�_!h�1ң�,>�n�������w��ލ�rȆ%�ݯi���d��Oڃޑ-d�W1nKsj�v�A�	����*T�poW�>~��
�e�UW�ŀ�l��7���}7��qk�̀{����͒�O�q0���������p����*=E��?ͅ��jq�"�
`��Y�GD�A��)����=������>q�q�2ب���{Wb�p�i&����Du��f~����|�>H�$>�$�#�$8��yi.�W[Lmhe�ݣ�
��0�ZwM/g���(U�?X��{a�}��Ġ*�<�,	�qٶ����[T��W��ВU�Y
B��e�Hp�;��dn�+�i7`W���]��J�W1���	���%�=}m�#���̈́P�r��{(�^�s��k�o����=�-(��{y��gk[������4M���s�fxuq3�c�����G�����v�����rL�{i:#65��Hq��i�bp�m B�5�2��}d�(Yx�a�T�:loLm�N�Ee��1M��F/�#L��מ�Du�8z@-�I�s3K�uO�r ]AB��k:����4�W������U<9[���71Oa��3>�� ���� 9+]����T�"�z
Ԗ8YT˅""�/cZl���cqz&\���R�+����LP��/�g�a���Җ�.\p8������4��}8@��`^Z�Mu��*���Zk�O�(�:�c�O�� ���;AL��އ=�B�i�Mk0����:��;��ӿdOP�eɗP<j\CgV��R%,�ڄ	5��A��Ԝ��G0�RY��Z�G�b�ؔ���x�3�ﳣ�͢Y����R��2r��;ToѢ�A�s
�����2���t�����Ͱ��P�/��}���A; �6�^���N�*��P��T�2�?7<�Ta����2�\�$�
��v�x��&���jV�G�-�x#c�A�74�xI�Z_�D�RN:�1��:���Z���=������7��ζ��>q��������/�6`t�44P�3�IwSf8�J���Ν(�V���5oۅ��f�?xy�9��I[\D��������hMa���+�}ɂ7��6w��<�v7�"D�L��Ŧ�vdÆ�N��Y:|��Ytj���[
Z,�����ڨ���ռ��e��0q��2-��P̎�t�9^��Ưi�q�8F�WCT��T�AN�S7X(4�(�3���hz�$��D��R�."�=��;�2��R�d�3�d�'$<@��&8n��uƣV� ��=�1hQg��Y�M�r�L�r�B����������HZ��������<����N'B|�� ��v�3�W�����<3Bei��C�l's+�SeO�"���`K��O/oHd.S��K��x����c@ә�r�ɤ�Kj�xJ|��W�	wf���P��0r�MZUO�>�o��֐R'��|�~l��\7�k���k���A}"�\�R ��0�5���J��L�鰴���<-s��Z�`���\/���� 0�ڕ%;��y�����a�I\�ېH5h]vɠ�Xl[��A�3��M�7TڷK���&zH���~]�	h���3����'AW�?^�Q+�)8 =e���O�a�N5���3n����[#&�@�I���.���"�z��e	�8�c���_�� ݆"m �*�B�Y���b3��������y'12�MV�X`��}`�*Q�b�-�۷��v��r�5j���D1�@�J�����<�!�m�Ï6gt�j��4i�տ���*,5�M\ʞ�a�]W�]Mю����m� -7�Ո�L$h�� "^G]���ѧw�o���p_ǜ\b�iuM0I�#��T�Q��J�r�qT�4=]��f�[�E���ivVy q�Q�"�C3:��L���k�^�r�Li��E���ܣ�;k�ڙz��(c፫f�5�����'ׂ`��g�Y��sJ�K���+�b'�υB��u0l7�u+�Ó�.X�+:Wv�G��	\w�Vb+~��\X�l�Dy-�m���%Ky�KЁ�ءo+��|��&�����K�b�'�ɣ2\��9��dW�􄐤>ʝ]\�1��i��9{�����y�����2�>��T;� sU�w E�H>�8;��a"J� �(^J�y���^�-7�k%z�A�.J�(!NRK��E�2&>��X����-��K%���n�1�I�n�������pW�_�b����9���@�VB3.��@��(�{Ũ�G���g<��^�/�����9�����.%��J+&7H�71]��.|	W��=Pi�|��k��,NZ0A���%A�:��`������͓��w<���m�$9J��]�N�"�5	>��HA��u04���&@�ls��'D^�_Z��A�;�j�Rc��dǰ�}fTðO��9�gYKL �#���?q]z#}��[��K�ϼzȀ����3���:��|I�]��N\!�Pp=7��(���p6w�m�'�>n(���~��F�LC:��|� G8�eu����gvM��C}*�Y������X�˄���9(�W��W�y� ?�)��R��(n�M���v���M/ȋm�W�V�H���A)kW�^i^�����D�ԇ����N�vTd苒���֓=�}��L�F��� ?�EI�� ���Z���ļ:KF]&f���׽m>�ͭ4&� �j�A��޶�o�CuFS�n�U-�$�_��&�u��{b�ߢUd�������"�5�7H�Y���3�Ac��%�mG��Ѩ �hҎZ��v~����1��0)�y�}hTm�"ۚݧ�s�>*�7`A�Or|�a��F��c��8�AK�3;Ey��W+�?�������^� ���V�Ivm���?��j�9�