��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&L�g_���w�����ʼ�ρ.�c���}w�3�������F�0�e�$�}�ΩFV�ld_�Sp�}58h��
�[e�Z,"��������v@Kv"�E�t �8��ޥ:��j��3q+GȾ^����~����;���q-N�ٕ�����r5���7�@�?3[eZ?��Y�w�R8��QH��d� v�n���r��.�|7=��B�J'{�=�pV�"ZTS�C�jq%S�RItuK!�mHlg�O�dB�7�W�C�\������h��T]tڊ�0�$vl���#��譤�|f�*�-�$9���r
~��p�[ ң��EL$fR�t��	�F�U� E�`��C�͐�'B�wAhC>Z�/B޵�Ȉ��G�X e��2��/�e�fL7��hԐJ��,1�~B��N���?b0��R�tu��gu�;��4���} ��n��D���sP�g�83�p&\VDV�*�f �mC��sk�ASE�w�&}Kԍ�5��nv�Vr^���Q�>9�����j��ʴml�y����k��'�=��>� ��ԸF�D�<ǅ3� ��+�2R�V�Ү~��\:�d���O��50\X�Ar��YX���?�ˆ��C���k��VX�޼�Z�۔�%�Q2�u�̓�|;�ˬ)�҇p�t	���a�	��F�)��5R��
vj9�.�࿄��Eڕa������4;�!��w+[{6K��������uљ�nОDP{����z�h�p���4��LoA1;���[��i瘬7i��q6�D�īC����5Q' �C����AyGo�G]cTj���E�N;�	�M:e�N��n!�g˔/<â�`�\�(���ꞅ����J���7��#_���3���{Q��(O2>�!s��i8��E@I/8x�t���8�����`07<&?�e��p�Q0���\6�ë��m$}X��3z��ʘ�|�*ww
��rL�����<E���F�c��=ٴ�j�B���� j�>fge��>�s%D� �i2ߛ�ؘ�.�i^��x�O�F�3�3��	�&3����q��5���,ǨC�}WE;�Ѥ_p9n��!\������Ζ��k�@0y��yV�t�k�/VK���d��
)�W��]
2���a���(�f)�|zX�q����R��6�=(���J��:��&�m��ik_��
F�9�۹�`����_f�_9�Yb�>D��̨`�^L��5<��	��j�q\�Hg.�:��P�ʺ^
����.
ZQD˼<B7��,0y|�����o�{W�}�G#���\)�ͽ���j*h9t��ʡS.�{D�6�!��Or6��m���=�i��0��]����jg��ܗ���$�!��`F���Y)Z�\��S�-h����@X3܌ǉ,�m����)`w���W��+0>�Ín��n�γ"0��8�/w�s�e[��G���ٛ�C�v�̥��ԅn��Wg��o�"Fd�������v�,����pC�?���͸p���Cw�m 1c眆H]s7]����Ig�R!q��k�j!So�����c�p\���w��(�_,TC�`�|��kh��i�+��PC�&{|�s���l��:LB�de{J��_�G��o,s�ϊcI�/�9�� T>��[�Hq�fї���;���JfGW��?�(�z�>�֝t�'��^1�2ȩǷ�?���o�����v�k{.��h��>X��ײ>�� q�F:����t͞�@a�ΞC�_>��t�]��Q�3�(7�q��y��48����&��R�K�#�J��w"e���4ҋO��!�a�) �{9#��uu3%�;��>�VF���� ���B�#����u ������@�P(��٨r�oMV�����������'�1��'�Q8����o<�i|E `-0�M��G^��9YCπ���1S�)O��q<�A��ɽ%�kZ�:��*�mE���T�)?��S��u�0����$����e�"K8�T�]�����b�����.|w[�<��# WJ���f2�|��M�t���wL��SC��l����~)�� �o����Y�n��C U�!�l�zd������v�Pׂ������\��ť������vɈ��(�^���x?���gDy�6;����[Zg����e���!E��7�M�Ptj��G�4E��'#t�vD5pp��kH@8N�Ks�������x#{/�8S�W���1��K*t��K���3%�-�]�O��8J�0��s�� �J�u��'6���wU`�z~�a{sԀ#b�Mw�}���Lj��vj%�jtc�;8�E+����B6;�~#���Gc�ԓZТ��,�
�R��=�մt��Ak�2�n}����X%5��|ˠM/»�ݙoI5����v��o<UV(y�a5A>�#���;3v�1U��5bw��i����,t�{��A��G���q����]�k�(w7K�j���*&��'n/��N(���$n��s(5d��y�����X���