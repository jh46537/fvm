��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)��k:�ث�*e�(AOg�X5����!��1��-Y���	�H����T�s��w�=���ٹf���aC��0�VO�JZ�ж��N{ɣqĐҡ���
 ���
.iT�4h�,e���b+t$�d����Q� W�^��b4����nI\g3��pE(�;�L𣐐����|��x-0}�ZE[�Q�v�]O��a���`k���,��_���e��3��;7��� �M�}�:RG���=,��G��ж��-�j��<D����H4�(t�!&��Џ�@WD�cJ+�g�7/U�HDLG�9�k�b��<tu��6k��1�!�*��P~�K ���l��)�J��A�^/T|?O��C���.����g��Yf�x7^�+�>x�P��F�-���w~�L���wЏy�'�f'�:�לW��,Ҿؙ3/��D��ߗ�����~���jڍC�79k�y��4�1��7��ϗ��1��J4X�����e�m^J4\�X#ƺvn6��&��X��g����[# ���ϯ�A|||�,pE���U�1��?���i��K���QS�R�!��Q�A`$ �.�=F �%j1XVc$�����
ގ�	 z֑���]�T9
��y�;���B�B(��\�*q�{��*�*�j�w/����vy��E**?ef7:	+�֪It��h��|ôΜ{~Q+��b�e��g��Qa�P�����=7�)�9B�'����%��0�ȵm���1t[����KlI��P7t	��b��w���yGٟR�Y�z�ʧ�=�i|7ί*x�y!�@=ӱ����xP�I�y/��$~wQ.S�K������{i-]����_�&T]�*���C��`�%vW�����4��@�=3����_A�!W��B͔��`�	�y� CT��D���)�$�>��6@��f�h���;�`96�$�B��UPm��C���˦��q�Z�*�#8nr�ٙ��p���~j�� lάa���ۺxG�$	�/��:����U�1"�k��`0�?=�^�j�q<�![��p��kC[
C^���K���>�ץ�k���`m%��,�>��&)��"�!�IW�_�x�x�sȶ0�̪mn4��_����+d���4�����=.}��	G#��8�"l���H]�j6�:�IHl�|��������fs�����t�mܔ1h�c_�P:��`/�
�j����7L�	Y�7�#��jȑ��_'���f6V~�{��	c�6�C}!'��mz^�s/�c���b3��ֺ�Z����,��G�&9�/��dU��y��S�զ�:��_����5��m!yq���q�2t�$̮ �qr�������ix��2>����<�>��q�}�7��K���a'[��3;pvq��:�p��l�ĕM�]ް�Z1H��~��C ��q�D��=r��j�֒�.��D�+(y�X���V�������l]Aq���_���2��I/�>�J�*�����fgA�Iݾc�UG����%�;:��<�_�����T)�H
��n}q�&{����ŝ�
�z�'2-�=�Վ��6=y�1e�ځ�v���t�p�h`Ȱ��.*�?4 ������sw��wLu���6���r��l� �4��c� B�je?�N�v���ޡ+'[��\����l��-	�N���A�(�NA9_��L���x�Y7k4�/�TwQ�(�ޗ3ɒ%��n�lE>�'�i[��O b�z���G4 ��`Z�E��=�q�C����;�6�h�Z$��N�Z�t��K��\�.>HP�W�[f�[��:�,-�tC��%)!MS����w�:4N�4�#V�/����>A8v�Y ���s�I	��4"ج?�șXA@^��B�{U��0
3�;��k�ȴ@	P�z$����F�Vә���Kd gpD�P�
Կ��I0��єI<(��4>M&��;tmn��u4il��w�&��F(�(ޞ�o��A���nX~�8�� n����l��=��o��Y��SOf�>���J���T(s槻=��s$3��8�}�o�̱~�xO1R0<�F��c��u�ok�X2Ն�������UYu7�;@���x\�';�,����Od�Ah� ��b�\���N/��5�!ļ�}>O�Rtn|!�"���B�֨P{r޸93K���T�t� 2Ⱥ:5U��)��sP���Q����׹z[:�J�_5����e<.F��D]�������q�f*{��DG���;�
}�R��-L;S�05 �р��$>?R�kק�P������U\�������'l���^������Y��dLP�i�$�XT��A����z9��sF�����r��:�P��;�0�C�POQ����Mٯ7�J�T,��4��5e�H�M�!��_E�[ B����\�I�j-�}5��X8��,�^f�gڷ�zbF�˴`��97~\����NRuH<c�n�s�%_.<s��j��?�Z�i���(ޯ�qc���q�t`7���+.�j��������#�|���V��b>�<���ͪ��~H��4Mz����3�~;�^[��o��|�?}mhY��^��oO]��!F϶k!���;j�}�W���V��!��e��,�Gå8\2v ϝ�^���H���f��o
�g��Ϧ��<�+���r�`*�S��dF3�č�g;��qKF�Y;ZJ���]�;���������{��X�C�8�&*��3��|H������\/c���f��v�{�{��SR�3��:k�#��(r���=nrka���Jkr�]~� >��sR���En�2�h�PIBKB���U#�s�cu�W�d����t�5,W�#/c?C�5Z�5�iL�95��|D�e}�U���>�e��KO(TG��#����_������P��ϐ0C���c��#�!3���î��
g�>׍EndC6�TS1�m˕ 8�'�|�(r�ef��V�?�2�P�-���ƞ}*zG�t #�-1e޽��FC,<�^yh��U�'Ԅ�"`?�bJ\Tںʅ�0ò�F�}�	�� ?0f������r��Q՞�͔�xG ��J���!)65�0v�/I�7<䷱�#��vga<,�c/����!���0�"�Y�`.�;%�^*t�?}�%�>< %�s�)Z�M�2Zr6Zj��u�,m�}{C�1�v:��_�`M��[o���/���5(Ϝm�Q��hu�`\� 鰄�Y��c����1|hB�厥ٳ�u�HL��^�81��^=�rAӮ�L{N��|Rm��F�.�~�\���� ���CQ#���-�74)x�7�j��!	���bT(�~�hqG��mVtQ�iy����U�`$O�t�M(w~��",ݫ2��N[|�~�/��Z�ՙ�`P�6�0_<yMJh�^A���D�0J�� G� �_ϥ��l/̎A8��-�+�#e�tK�V;DP
JA����73����6Ų�8:^���X
���h�ޘ����̶�,t9��a�?x��Q�Ѽ�&�~�t$-���g����Nc���Y�/�r�(X!�X�&'�t���a��/{��Sak�Zb��o&b�v[urӍ?�����&7t6Z1�4����ES����)����_ 6`�SnJHm�gѕ)\y�OHM�k�*�)��Ms;o�NH��z�g2�4,}�9�˘�7UWt_T)۞��?�y&��ʘ�����U6-��v�xO��;\ec�5	��W���w0�B��g�v�0��������u��b!O�޳ 7���P�����//s��w�l�	/4�s��Yv��Բ5���!��TU�A�:�{eg	�V�W��aD~hŋ~X���/�Lū�>V;&T"b��������'����#�J�9�pb+���a��;8ۇ�r��g���!g@��sp�)����*vc͖�e�h0��^+��dZ� ��O����3VT�b�5��a�K�������Digb��i�mP�#���
Y������|�8YD���"k�,��8�xJ���S�Y�@,��ul�]٢����U	�����%_��y8��ʯ�o�~�|x�u# �$m@Pb�� ������7�ֻwiںL��W##�ȁ��x�
�0��|�=��+ݙ�6��8#�hf�9̧O��e ����!���߭�'���jCv=���b���`� 9!�<+͎�W��!��/���Q#�dL� ^FM��%#m�����@�w�á� f��6~jy'R��8�k�	m�CF�VR�D�F=�7/��:�M5�����[G��#Z!Dbk�Ì_�I��`"�:	:�6$U\:j��P@iSċ������g��KJS����FG:;��)ի�J�q�A6Dh"�z?��8� j�I�|��I�b�a�����6f��O�ɴ��@� �i���u=M��q����U��x��C2\A]<�@a�ޢa�"�F�e�xG(�P��c�o��>#i1M�
�W1���[�u|��N*�����=��=8�mY�H���K�%r҉���]P,��1&����ai{m]g����;7>�lk�lT<X��֮�)�AW x�,��Я�ѵ�K����޹���ε ���^��q�����{��i����R-9>o�я,me<iu]��$��|?"H�J+N/f�&��<���q�E�e��`i"�'Vf*�Ș?K�~�HDosP�ֵD9f4dz��H1�H�>��Q��v��/t��Z�_�h��#�!�F�,2*VfZ�H�	r��O�f���w/t��cX�@���bH���6�r��b5�!��|-9u��� @�si�]� �`@��m/���6EW>H�\i=��48i�j�[�M�CҾJ7(ى��IXd�հ�� d����l��X�!����ds?Wޱ ~n�(Ҏܽ/��!d *~|�}�)�`����XZ�#���o� �Z0�]�暆}�n�~�Ǝ2���қxk�A�^���wht��.�Sx��'��'�a�@,����g~o��  �X���6%t��I�H���ԗF>�hPؐ��&|�zlc�8�x��'���:���T����׎Y����V{�+�Զ�/�OA��dƋ�Xǘ�%�F�
FȻ�W�E{G� ��,r?��