��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2IayAMY��{K�(#F=��U.Ā��[qp�Xv�:X��~X8h��#����j�mo w�G�ʃ��{����%��1�E1�(v�b��ߵo�Y�A;t]����Y�~�'���dQ���^N���|ڄ�����zԭ}����~<2,xҭ��7:�}�ؠ��9��ڱ3������û�X*9���z����6vF��7(����(��s�M�N�P:�M��;]w!м��y=;D2�ܺ�����ʊ �EJv�����d��J�Q���%�<�]9����r�^/�&[V��B�wl�	�>Y7}�E-.��)zf�-�cK�ˀa���6$:C����n?b1=�[�����_��O��p�/������]��	�X�����Pjh.���
iO꣇v�CB��M�(�GKx�i��RQ�t��֌4��a6���s/��U�SE�z�[<��F�5�&}���+�O������9��`)��0�cR�o���Y�����x�0h.����a����]x9�V`�怟�6g���i<R-�}}-�i�l�a'��+���l����T�~��0f�>W�ؿ�msM�5�j ~	�\��I�(����:��'����2�S��Rwq��s�U}��m�K���&-���-����*�'6�j ��>�9��b��;�Ǿ��@_�aa�����/�6d���Q���<�rU.e <M��<�j�d�X��)aы1�	�6�M5y^g�;Ivbm�n�]J�Z��k�=^�DΪ���֬��B����x1�y��a���VTl#R���s���Aբ�¬�A����S����>�o#���IZȸb_����G?{׏p_]�fJ�0�g�$|O�V�L�"�y�{R(9Ը���pGa���$ %3��RH�,螺�U��wl�	�����x!ɝ�m��DC��tI��.�r�K��^�z2�U���[����+=F0�����Fj�%hX���L�f�����������T�GK�p��.�liZ@wQ��� P07��ʱ1�2F룒P�v	���x��|�2|8
��kꃉ�h����N��S��= ��gDĶ�ZHB��N��cn�S�&#�
E��M�P�̜;�th��Ѿ卬����(fW����~aIhL�P�Q/�{���a�Ղ6���{42����07.�Y��2����b�/�F>:`���M��=ޖ��d囓���Ƅ:���1������3���ZDU$�͙9|Uu�_~^+0b.?V��N��Y2{���	�΍�h���a�����>e�k�t����x�R���|_:־��V����I�� ���&O�v�	^��⒵���~&U��("v
6+�Y"�ls/V��0��7�3��0Ti��Kẅ��*�E�"S���A��xOL,���q�8���fu��k8S���Դ�����yױ��
"H	��b��#�Ə���)�q<�j��T���_��-<%�+y�?��3��=oW-�J�(�p���i:1E��Q��;>��M'^�1�(������X�&��a���2�����oa^�PEؘg�[�G�O�ղr����P&��O�4p�k��Q����>oK7�}X�i�N�ݲ���9�pZ7��hZS4�`.�	��6�4Z�l��\Z��Y�����G0ʶg4nl���0�0�AK�i_X�����Ҹ޺�@O��?+ضKb_W����J;D0阐���GIg�z�����"`�^I�M����ޘYqj���kn{}���q���M>��)��f�X�
��]�۲{O�tT���N�ǫB�SO��mK|��ò�w�j�.x6$��]�g��I����V��C�g�"҆��@�z돶FKiQ�g�jI"_k��
�!�:E�6�5�>�|�UM�	_� V�y��QL��D{��� |��H���p��>�Vv�_���k-7Œ2O��8���@\ ����ߵjT�'�-��.����Z{�;�	7�'ƂJ��(E��zEk��R���z1��$!9�:����?��V�N]&����G�"\8��|���4I�lő{<h�5��sN KL6���D��W��]Ź�Mh��1)�y��u��'٬���qb]) xO<��&��jf>D����e��e�ǛbM@Z>�=�5Z`k}���.?F��P��(���v�`} 
r��;zj��~��YKպ�wD�9P�p�	�i�)���Q7�<�#�c�UX$1��������.�����Zl)�J-�m�*Ɠ�\�^_)F�Z�Д0V��R�~�܇-5�ѥ9U��:&e!����K�i�q�볚JB�Z��}�Cf�0C���������F�Yk������{އ���Z�O�&VɌ|as�J�(Խ=��,�T�J��r�׼`_z���*G�o��ǆ����%�d��B:J����EIח�����OQʆ�WҖƼ?#D����#��v�� �f�k���������8���.�Y���FA�������j�f�҉fTF]>1Οh��u�	>�7~�Ϲω�a��^7��?��X�E�j��yUo]�}W�|*�~����O�����i5��S^UF���|�"������H����ι����ح�D����Iz��=f�ԒF/����I (	�>���I@C�j��H3�n���蚶��+ �)h�iE��J��N���߲�8z�(�1���K9ጁ\�Q��r�Xx{r����7�@��^�<��1�8�%�����e�3E.���N��H_'+�9Fx�I��&�80b�5� 3h�"`�.�q�*�{��'��C$��KJʤ�]c��9/o=34���lf�*��$���%�����~䝚z��k�kM�aL��W�Fy'��'�C\�MΙ�vܴ��4���k3��H8�x�Cҿ�P`�(���T5��_}G��*������Uj��T���?�9��c�(++��l���U�f�i�u�wK	G���.Pl��s| ���j"В�l7[nr�*j��7edL�05�`p�"�Y�QVT���n�˼��J��!'���&{�~?�]2��r/ B���C�qÌSX��<Sj����M��F�[��4�-�|��8`׏Һ�
P���3y�Y q,#�}����6��X�� /wP���Ѐ�g�����Q���"��o$qBك^v��ٍI|�D����`Y
g�R� [�^��^R�1��WpK����l%��կzچgY������;�'dZ]؎���X�io ��T�^TL����1��Ʋ�O�e?�{�nIA�3��*�9=ek�Cc�c�nl�F��Gj��u�f�g�O��V��
�r9X �jB,�V	�
�R���"�!ҏ��2�SO���LN�������ݚؖv}�04+%�ܲ����V�Fh`M��	����d��A��蕡ϖ�@��k~�/6��kZ��/73�j����wN���rb���C�vjS�Vp��K�:y3��D� �F��ܣy�;a+uB��$�k�|����d"�)�Or���O�B@41�BC�YCT�k�.^��tF��g[��Zkۜ������ۙ%x�}H��n+���r$�_�5��AJU����,ԏ�F����]��G
|�ۋR��ml`�@��G��ߺ�0��ۛ�M��	����U��?8vs(ow��?��gA�a�y���k�:��^lY�R��9f��oӷzI㹑@�������b�im�:m�UV`n�`�P�9�T���"�8�b4�wRI� Eeſ3)qA�+�tO�������M�����S�����B'l�;�d�M_�(0`��K&?q^�P�k�"�\� �`m.�Bu�jMo����� �r�{���_����T_GN�s�X�o����A (��CTꭻ��1b<�^�����N,`�T+Ό[����w-.��^�< ��'c�^t�8��9#.��p)'���a5[��\-Z߼e��9>��t<�`�E@����T;�MG��U��\���:S�gʹ�Їn��{U�#3K�02�c��7$��P�'�Hl���+��Z�$�ftGqN"(�(�pXT�
���ђO��p�YC�sc�ѩ��1�t)����-0�gZ�\@@�_��Y�;��%@S��̮�醋4'�;�6���A��:�r ��g�aI�Inq$P����b����h�#6tM��3;>Yخ8!S	I���)a��ȞT��hKr�n2��ޣ*�|��9�	s���s���� θ�!��̙T+
,:I����l8{}h5�hbb�ii�J�JP{�z���.�[p_��=�����N⽮颮jv�V=��#��E�&Q%�װ���h �u��[���f+��6-�o�?v:�0��ΰ����Xyk��{���k��6�\ɨ��F<�U�7B��W��BuX���ܼ���Ŋ~} �E�Fq�-]�W��|? �`�l��Z���}��k�Q_������џX�I@_�c>b�[oZ%�ny6�#�7ůZ�V�7ۦaV�^,��&ym�Ц����Iϱ��Y�v���	��v_H�p�6�-�B&
~qM�{�ͺ��k^X����g�bK��w"����%�.X<��t'd[���$�B��Ԧ`�%~ćڗ{�t�V��}Ξ�I��N�#}gJ���Mt���Y(���͹�whIj(M���/����Ɩ���l�6{�a�ǌ�"�=�fJ��z�3F
���p�#VL��]�)�~���۹�������B�[Tư:��E0�|s����7(��~�ձ��A eR�{Z������Nv���^��ى@�Z'�c�T�u9�y�R� �����'���N�W���cmYSN�. 
t�xvЁ-�Dr�7[�Hh�U)�ٷ2`g�
رU����Lm���v>�����2q}Կ<j���ؽzf�F��ɑ,��E�Sb�H�O�J����O
�R�-;D�dT��;��[3�|mQ��|�^i��lW��dm'ߕK�-C�_5� �l���[�����rh�G+_�R���v��]a�t���.[��k����`���:,\��5��5*|�I�_�L��)�@�W}��v0�N$둙�}�Z�Fɹ2��`�͚����҆��dF���*��EbN�\��x�g�|+i�J�z����Hƅ�b	]!�e~��=P��P:߃�R?������B�aV�_J�Âl	�GE�h^	�+�Aud���"F-�"Q��!O��vGֲo�A�S`�_\5{< �	 �#�$�K�� a6��-�B��Bw���$>b��Vo��.c��z�g4B^�9[�{�<��N��O�u�4YW��f�8�1e����@ϿF��hrWL�M,T3��2ݼ�	��ä��Lz�(ű�rgW7.ѽ���w��#���K G�%/]NFV���Q���[A��rY�'��