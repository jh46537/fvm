��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�=WM�Q؅T޺HݱCV.�+
^~%|'�A��`�B��ZF�7�lgL0�YC[^"Y̬@��Dbz#�x��)�$?�x.ϵ������4��n&�0�X�\�j*\Ѳ��fO�j��D��g���T�SfbJ�����抵�w���_��C��P,�2�j��{>���?]Rof�,�ŭ7�9�I!��_����׽@�>��]75f�I7�j"�ƕrϴ�ۂ��%����6�:�Hɶ�y�z��Ͼ�h��Y.�uIJ���OpR��RjL��/Sz�s����-Pڜ��v���ʅ��wJ��.�WQ ��j�K�4PH��� 6����4�IjGS,$^�n�V�`��P+�{��2����o�BP���S?9X�Z����t�P��	�;>�����x�P�j�	���Q�a��s'T���/���g�ň�g��W{�`�9��j�r��t�(l4�8�↉3�R�$�e�Z��e�7��ܺ�ܸ/ʪ�l"���R����i�^+�by�b?Y���Û��s��/�ɋ'8����5n�T[R��lYx��rG$��:XQ�i�6Qe�6��F𯭆�����;�2g���Z#(}['�R����)J|j���F[^v{��/������ʕ�+��]���tH�+��r�* 'J���r���!u3����I�Η�%>;z-V"V�'m�)��O�n��r�G���"�*n`�a����2���'n3{X��݋6^l?���F��z��XO��H㔶����[ٰ.fVڏ�m7�f %���m�|�5�(�\�c�1��&	AOͷ�\X}�[��n���t�ak񻸭�@=���>c4a	wL�,uV�
�����C�h���l�zH�1�z����^�����J��4R�q;/s�b,ii-g�O�F���� ���ij]�!��8��v,�|�fen@R�@L�l,F˸a��UO���;��,���IRN��F܉���΀�y#MpT�F��4VՕ��~��a2�D0�D� ��nC�5�g=�(��(��>� �"�b淪��b|^"hi�gx�R�}�Yy�����VM�A�R#	ʂiV���f��So����_��ى�!O��x�s`�m�I2-8][r�J��T��wͬ�A�����ʻ�4�]ˠ'3���uyի�|��ա�8�@�{����yΰ��a�{���ݛy��
!1l�o�������{r��G.�8�@��!S��ľ���t5͓b]榟:��!:�mc.{5�a��
���|X��� �w f�{�:��Z.R��k�1L��+6 ���|;��:aM��X� D�K�=-'+�0�~U�����d��; 5���xr�Z�����>D#NBz���r����H��<�!�����k����pj���@�:X�X�YKڊ�fH�\7�Uyo��ֵJ�,)���o�@��:�|�yܯY��Y�� FiYF����&�Q:�oO��T1�?,�X�{�̮��Κ��L�;ģzƕ�:m�D����N�)W]0��=�����|�d�LS�Aƥ�)�Ĳw�pl��x�SKFq-G� R?�k�����EE�ޘ��)K%
�yb������ϗKr�9Fr,590!r%�h�*7(ɽ�RB�1�B�X�Ĕ���������*�~�A�Ve^�
���}�U,+ɴ�v���\"��и͜ħY� �DRD�ɬ`�N�ᑧ��K�ՠ7:̙��/�-v���BјY ��I� $�Ь�����?Bj��i7=��Ua�_�q�4x�C �4��W��r����"&�k�W�����\�Yz�N�m{�N���%�+��z#T�!�^�� �1��(K��"�*#���g���2H���s�r��w�N��[�ڔ��?bA�.��a@�'�� ����a�.p
eH��oW�]�J�U}Ml^[��x�^��S�6�6k!ß�̈����
�����I��֭)��P)d}mC:wg�!��������˼PRky�؄�������ߠ�~���#�3���}TKmu:����1�q�ȸ�f�>��mg;��.2iTi��(�tA�ܟZe���3Y2_�z��NѴ��ꪟb�BL�-R<�}��;F
M��;my�e�N�U�&�*�Z������X��NMz�����2ԟ�i��R�4�_ň�Z�~�`$ $+"O���Y���(�]��3F�c��CV���B���t	4�N-g�θ=B����9���+�����o�/64�*�G���[����R�N��Up�(G=3t�&J���E��wV�v�3�H1���_"J��D�ф�j#t���A� #�1d}�DńT���.I0_x��A2���M�C�
 �����W�f��B,�2���x��b���;���
0"�i܇�� @��4����D�m>��V��?��5�N¸��N��:�j��Q3Q�v���dr�Y/-&3�2Q�����<� $�B����_�7��t�X�%��؁.Ҳ�Qd�9w���w? �C%���>�L��V��n������F.�:x�Ǎ��@�iN�]I�SP2�k<�(�C�q����2�b��i����@$��% �V(���e�z8ƽ���%�j�Hn��$�uG�@c�!�1��06а����[T��=���2�l�	m��>�@k�Xgʅ.g�鳇c��h1�b�b����6��!}P�pa%�$5�e������������	n��-l�����#�=�Q�B&�.�J?Ds�(�����Bj���j��