��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^TC#�yM�g,�%kڅHе6��&E��1^�"K"o19o͹/��m����ts_8����^$�#�3�ow��T_q�4��B��%rZ�a2�����0X�5�s�У�M�[P+�IC���{���,��_-Z�YZ�S�L����v
��K�xI��Oߑ��q�������K������:��$�'AEO�7��k?�TD�Ѿm-(#������f_6а��$N��O�Z�-rQ��0��7�wC�j�tF�e	�|����CF?Y �H��b�A$|�3��,�"�M2-���Rk������_����)��]2�W���0�ީ�����yBFb=e�c����:�`�_��l}�� ��vƏٚSd�V��:�*"L�@J��jj{{ϻa'O]�m)f�=dD�@��?���n�ۥ����[�[k�	�6ಋ��\��A����4Lb�bu����l1���?!Y�0��Zv�p���Zޒ��}p��(��i��?+ ��gD~t����+"���W�)�?^�/	��2������Ϗ�o�V�J�	��@a��0�/p�Q�)߆	æ<L0b<�J�,�#hh8��f�k�41�I����S�%
�� #�F|�Az|BR��ь���`�=^�.0�g��v��ɾͷ���e�T�=q.V4U`�7@t��	�JS����I���I"�, s�a��9<��f�;j;�+��>��8L��km�p\���K��O����/�醋��W����x�Y9m� s�����ň���xgk�l���!��er[{�ʁ�Z�o��{CqtC
���:�u��z`�z*C��G�$T��F��P��0:@cs}�g���K�o�;Tb
��x���E�8iRp�)�..���/~F%WO��{w0|h==�-��V��pf���MK�t�t����Ja���}�!���l����Y�����;��áO<zj��`5��Q��ƕ��/9����ۻ����C-E����<���d=�.�� 1�hl�8eBE�{���Q�7{w�D�J"S	R�(@��J����p����&A�A�Q u��n#7JU���>z�������	�^ѐ�vxkJ��)�6u53�_�e|a����w-+�۰���ὲ�,W��EY(^��D�\=�ƥg��L|�UYn �g�%��c%E����Νͫ<� $s~s�2$�H]�)�s2ڡ�j9�!ȧ���@�)M��	���so�������d��;[�Z_L亂`��2��n��
<<��O��꣖��Z�cz���%�,%y&#��	rA �0���^���0P���T�%�G�YJ(Jȋ7���â� �����@8�=�O�y8�O���������=4R��k�A .0��U�EI*�r_���N%��[[��xcY�9Y�6W�ĩ]�I�hU�+��jK�jY��_��e��{��%��a����*��F�\��~�7��?p���("���A"��0�$g�:���!{Q�����)������Q���޵�y��;�HU��Q1]���qן��UQ��v��o��"�&��V���ɽ���l�mz;�GT�25bfV},ۦnP��#'n�4?��||�5�ꎵ��(�m6cq����[up�>R��?�>B�����F�:�?LI�L��v9�r;���ǭ�S˰P{�~��J����u��9��t�6tlzͩMAG"Z%Q���!p+$+,��r�3CPI��*���r'���˔�k`Lū����arO��^����ٹw	�W�K�D(h���"����@�2Z�śdy�Xg�Z���Pv���*���U�ٿ��ʚ2�k��Uw��� D����Lg	.!9#di3����������k�[�ʩy���:#ύ��T ݝL;r�L�Dm���<��3��g6�)�g��9�\x*X���_���;���9����hX��S����^S5��G�� Z��%W��!��_#��Ս"-���Rn]����r�yB2���S�9M���5;��U@!0B��ooƺ�K+��̂Х-T�O�"�R=L[�R����!��v.E���B˺��h#'R�;X�F���sM�ca+w,��ݧF��w��y�rݙ�=�����"��j��������},����� �0��i�O��	����ý�?(Y�W�^
����֙ff-/a�#E��kBr�S��chP��B�ڊ>[�PlӯL��ks��B�B��0��Z�"�4�����97h��)6��qfo���cQ6�G�0κ\|����X����S?SD���|%����Ҹ�w�#��Q��(M��W��F��`S�@�G.9"��Xl��_t�!�����ۥa�����I^�'��y�h�)(r���O1b�
b��R�~X����D��7��&�I/����;��XKP��N���+��F}r�Z�`~���u���5�a�pb���b?�*gCO	���T8ᨑ�����H�qB�����PL��1�,o�ׄ�q#VV&��=^�|�Z΂�u
Lc��"v|�B2|ݽ���y�#�>p*#��ul�M5`�p���r���_y�V}`���1�
�9ZVM��@0�h�^%P�ޟ��ŷ�W~�,�wԎ{�-�6&%��<�.���유���iQ �����Оո_���>��7�/$Bv��u}A�U�v@P<�SG�2nU��'�\?W�����u���;�kgw��
��i�ʥ=
@J�i��E*u�R=|���F�����2�s:�Q��{Zq)O4T�O܎q�L�"�x��+ ���T3$��74�F�M�_`�:j
ݸ�H��i-,�l27wC8�34c���6�`�&���9vT:mü�A.�۪��Iw��K��z��=�����\�$��(�@� ��V��4�JS��|��n��J���h�Zg��粷��X��(OOb��ƈ��ق$��.O�{�GH ����oۈ5�Ŗ���\�{"��=J����CÒ���O��#3-��y)ԧ��p��k�U�*%��GCY]��lm���jM�� V]N�jep�_�r� �cVT�싳	>��6�i�����sE��ؽf�����3�}9��V�7[��v�������'��f785,�և��i��Ϡ��+�����+��Rpg�t{',x�"bwG�i3a��J�E���0M�`ʲ��$�8�wd���:f�������&�Q�{�Ԁ~�N������45� �萻x�<�"��gh:!�bz���T���yJƦ=bo
�녔�XE�Z�N�Ĝ�响B�#�Q���MeC�Ϋ+�IЎ�fk���w�U�0
;���w��}<�#�چ"����Y��ʇEo��ٍ���n�:,B�k��ޅU���:�lvI�����犷�M�i�-=�ɱ��xx�,9��m�gL)�oX��v���j2�*e.�0`�ĭMa�����ڮ�,`��z��!׎�Ʒ�}	3j~ҩ�-���`!��c�)�/�X��>�Ʌ>;�¼�[���.hb����d���,���Á*�(����o%�QA��x~*p#�%�evC�ǣ����s9��\��0�:]Y�$*�!׺$ Pޥ�3#>��O��"�@i��],B��v�M�A��ғ�eq/��͵��L1�����;�(��,�
��/:� ��Ke�����d_f�R�2�w�V� �9���ÿGt�v��W���6�%x��O#(p��m�yDѳ���f�e�lxHS��6. ѽ�H�L> F=�n�d�8	tbU����a���Q��h̹�u�?#!����5l[.�i��P,��NM�o�d4��#��x�s�Q��eF-���昛��Uz��5�> �rRe
.6��_1:�=0�������d1�j�C�lئ ��b�
F�t�ǪI'f�j;��s�R�^o)Y���Y�2��-�V9#�NRZ;���p��S�ݰ" �'��V^�~�7��Ʒ�R�K��K?# �N�W��Pq�oE��e�p-�4�Π��G��=��EuT~R��^l�ʵ�;�F�-��~z�:��a��祖,�����
9�߆���}u��bLD�>8��f���i@�F���\x��vI4~˴��hN�����6�ɇY��d��FL$�hc� ��{ �U��)�8�$�;u�,��4�����*=ƶ�6���S�OU��&����|c'6fǲ�x!wm�9�xs �cğf��,��i�}�NRε8�e��kp���~���K�ϵY(�w�A1��������jr��ń���iBt�'���׍D�S)>�'��M���i��*y&���d�z�1L��x��_AM@y����|7��>���}нdʛ�D��{�W�v��s��C$¥������;H�ڦ
O�u�){7=U�99�f�	�a�8j@^av9���J�=�H�&�*���j��AJ(��D�R�}���uң�!3x0���Y5�qiۧ���X='�ɡ� �G�:fK���E���<pƛY����N���;��s�Q��S�jAV����gt
�f}'� f�p�4~Mգ��2;�u��N�k�n'��w����I�e�F�o�x�q��i�X
 ��CP�622�%�����Dl:l�$p<������p65�"��#@�:nM��7�� h�Y+F���?�ԺѼ4�/i7n�����yYk�t=���K��ЄR_<�*���T�<� JC���f��D.�[A�'�����pn	c�%I����`�98����B��[k.��*�j�����ovQX3-E�Y��И��(��ٛ"����=O���"�a�S�F�o�g�,���ᨫ�wZ?��k��+/O�@�*�s]�Y����i�MO0*{ey1=��.�WKЧ�Bs��x4u��B���:�ĳ�=n�68E3X���0þ�	�}������E����G��FѓR
US�R����G�or��%�e�o\���L�6IO�'>�/��a���':2m$�>ao��[�ѽk��ɫ��BPG]k�BH�4anMuևS�`�I���N�Bb��ܨ<�m�a�p�����5F����4�$]I��.t�*U'��y��L�\z�~�W�Z	���
	�:z��JS�
������=�+0�����|��<𰬖9���D��ְ Yu�bG�x�����]�q0j��<�m$�'>M ~�N���(�
�/@�r�#;{��8�/�$<yB����֍謦��5.�i�a1�oW�ֲ�\������*�s��c3������:�PS#�ɹ5��n��D\VA��)[N�211h�͝������y,gs�F��l��3)�.w#Tq�d�ÿ�tt[A�h�� O�럓��!�94MST�
��a�&��ck@��G�����v�������=5�Z�b``y�������a�@���<Z�s�.�_�ݑ�ψg�4�Y}�buT5y��R}�Fۼ)�<�U�@�qi�