��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbyj9�ݢ�J�i.��M�.rGm8.�{�r[���JǳV��TSA���`�� Dy��Y��F�,Zi�<���S��z߆7QTY�uYuE�rrd׆����Hλ?qr�&�.ebyj �k��u6W�+�/�>aD�w��cWWQޞ�ߗ�D��dy�g��[(�}��[�"A&��B����ƽSD�z?/m%�0�c��5��*�AG+@��pU=���������A���S�֔z4�������-DQ̨InfW=#��#2�U}G�2�T���Ţ�Sy��Tї3�WD�����: ����D�^N?���G���mO6o��JX���l9t��N':F
��^��0,k�7ቺ U����B�d�W0��жLC��Qv�ۗ����]'��d8�� ��V@()�8�fE�	�{���,�{\m��mp$[ �cT�rh9 �����}�'��cI<�T��Km����܊��WS�.���6I��i�Tض.������?4�՚L3b$�W&�P������t6T�Ġ�h33��h��U�U��b+����X��M����t�љc����3�G�>�5�ί�<u[,ܡ9{N�K+ 89��E�F�N��T��҂"W�"��'�5`A���)&��N���׶Z��r��0.�sY;��:҄��%V���E͐Q����2�3c��^�3"�fӶ(>ĩ�2#�.;�r`1���{
�m��2_����R�'�#�[�ot��u��[��_�|w������x�'���gxxHa�|)]B��H3��y�+���}�^�{�gaB�A�c�U�c�神V��o&�l����������`M�z�n��'�� �ټ���W�'�c;4���2�C,15{l�Ŕ7c�'C�����ڶ`G��u�+߻]�!wE��b4z���5��e��z�b��05��<����'��ѷ���1��̆�"�Ѡ�즣����W���G��*q6xT!�V�L��t ��Z�E��/5�D��g&o�8#ϥ-
�}_��;p�e�3@▿X�!`�Ԗ��O�6C-p�]5����)eX�R�d>` /���-M����"���1��3T��BP�h����'����N��v9D&]Z�?O�/'�1��.�p:2&7kA�
�����b�����	N{UZ!GH�&
����\�˩�%�H�B�Ԍ0�SG"�] Ù�-��bEܙm�����D�ɴ�͋_��M�F��U#_i@��6йߕ�����R/.��rG�mTdm4To�n���Xp�����s�A�F���޲��������{X�4��T�5�,Bv�N�v��4W�-�{�{��B��.�("�3�zs-�1w��Sn�@��'v�{h75<y<C]�ּ��F�l��I��u�����P���H����jY���B�nV��/�=��
Q�/�$����}��6@8��F��𽷥�8(��Q�w�d���4 @�����]-��N�����H�R����V$���<<�8��xSlt
\�-�	���s��ZlW��Y`u�42��P��* yܒ�/~۰�*=�X����W+v|�h��9��K�8Md����:+�����Crࣹ�n&�,�U�&AF�@e�q�b�[s� &'s�O�a����]Wl�����ăy�bz��D��^G���t���z�����K9J<�O$�3�;o8f���0]<����������B$���c�7�Uh[{l�b��i#Qw�;/KKkoa}QK�5'&�ߺ�
	�@��f��u�DɜG�qo��� �S�Z�K�u &�A�Qx�NL�y)n�y�u�ufQ6�cTn�'7m�������vjb�{�Fw��-�������{��(Ւ�Y�!D<�me:%ʅ߉��'��wi���q�t�(�Z�Q4�+<>���ڕ���%ތդ�c/9ڿ��#`�!�*��,xK��x�7��x? {�Α��-vs}���W�*�ͫpxhN	H@F�+ V���7�����g-�����5����(X���r���0���Ͱ$��=L�X�F����z�Bp�S�/)�����Q����:ctB��y�Bs�����7��$%"o�`��7��P�yVMi��Q�
�M�/������P��k��'��nSّ�[6�6& �6�fA$� �b����KƲ�����C+��d��2O�'��9=r���/����B�m��ܔyO�$����Wʵ����i���ÊpF#R�=�r�	eK���ʙ///�	��'���U,R�L�	]�G	�:WݩL?�*�"�����%+���șV�r$B�%�9<�&"���-y���S�e\���{Z����Uūt��.��Q�E_�~Y��ʑ� VF�}��x��I׍�@6��q�0H%@���e��%V�I�������h:]&�Dv���*V�7��R��B�k��@���0\'�^�q�K6�*!�M��_BO�љ!^�#�g��΄�z�ǚ�Q���H�FQq�{I���e�c��
�������F�>�=��mE+Ȟ�Kd_a�����7;����DB��� ��p��,|��BU\��{EU���aG"=ŀ﷋��W���b�H�QM��z�H(�A$\h���R{�%�C\��H8"Ҫ�����[��X��r+�܀zw�i��h��8�w屴��{x�����Ǥ�9���=Nx��O���;P-�2�IǦP냥bQz��iN���'��s!\��p���j����w���K��G �x����j���,b<=3��iAά�U�D��N���
��E��2���%ac/Z��M�N���F�Cw��7���r=��c�4�&��$t�F�{�9���I�핀�3�}?�#օ���r�\�׉���$3�,�Dg�����)��q���5~��W-�rǓ?�$�-�
���l,)�=�s3Vɥ�I�Es�����FS�D]F�}�PG�e@s�@#2�+�A�?�
:Z7��$i��iF:�LY�-�<��춷�q�����N�6%����f���Y�p�U�D?Y�?�Ės��\�!���ex�v�'o\�G�����J 
��((��a,���U��/*�֦�z����R~D+����C=C�5TG�~5�X��$v�� 4�Fg��� -}��&�"#
��xfW�W.��ӱ�U�~h3:]�u�4F�F�D��}�F���1�����&"-4WD�E	��/�)o�R+Y�e�ݠ�E�#��H�
��
Jfπ=�	'���Ay5��ʖ�*f ��WT������F��
��/|�C�7
�\�L#%m�#Ĕ0i�>f�|W��p�D(����ǷRF�|�?��hf&>��۬ş���`�ڃ�6:��� \�+V����Ǽ�ؿ �o%��u� �Lλ��������s#9WgIr�Mֹ���:j>i��0Jg���@�ߢ(����|�@d�7�S�S+�.L�$�-^1���~h�{�6�v���TZX��Z��{H磑볂�;űkL�Ƈ0�C���;�͘��@�@	O�L踒;9���CB�c<<���y%����R�&/�07��nK&���H#Z�l[ߨ��c���Yg]�r��؇t&�'�U,u��F�z�Yv�]P�&�_�����20�o���yUIM>�|iiǄm[ ��m!���%�*�Sl_,�c?rKM7��lk!*X�h�c���>w��o�z.��׶	�H)��~߹�K#��n��-]�N�F��5I
~��>��B�����v�*+��^���@$��й�W�&0��p�5>>�{�����zc�����:1���y%L��>ihݙw(;>�$b�S�?�>�J8>[���hr���-��ƇL�7��WU&U~�M1�D#�Ub�u����ǃ�5�����[��?M��A�Q1�� �>���8zi��އJ Y�R�J���A�ԡN*�k7��S��09��Ȝ�4�S�Y�^��s��F���Wt������-�"��9��j��-8���eu�}�����0a��9U�*���(�
�o]�<�D�`�R-�*A8ը&E5�]�$����^H���C ���-�?������OIoh�k�0W�ߊ~Ppd���p"��?\�'�����l>�r�(� ���+_�Nm/�ls~��C��q4���$�(�M���=���5���ԊF3�gy��G�J�=Rzگ�Q�!��ݲ���;��N�Dg��o~��"`Lf�:��ցL����č�}�$f�$�h����7`��m�ƙTC��R��^C����w����.c-�9-�g'3�����.j��+�]�^2�V�K�d�G��;@�@	-��c�|���o��a�]'���ɥ����%+	��\�'��"f��;�	n�R��eN�]��KB�m�4,��:U73����,�p��x�	��Z<���%��t~5�K�	/Y�:�˝��+�s.Y;�C�����M�/B��wy��s��^ E=�-R����ci���B���?�ٍ��O@�S	̹�T 	,ZEh�EC$�3�9��1X:?�^�<H���y�Ѷ=f��[1]e�g�/hቫJJU�D�7�0�<Eڇ��iv�"cɋ1���C� �M�X���/�7��!:�g��~��(��Ɔ��rB��/L-4/�^>��޺���ț��f����,���;`�Qz�u3o1K��������S�� O�F����L����O>Wk��7�sp̟��ئqB방D������R]��{��hq9���Hq'�8�}�q������j�<�͎B�I�j��H�I�������ޢN$Xf[�sQ�~��d���(% �^�) /����DX��_���W��U����Q��n����7��$���JO&�Z��MҏO󨤃���E|��2^�8 �q]���8|-��l���R�(F?�b��[�nJ�Pi��dT_��Ad��9F����;�3@��/a(���� �PA�B?���4��>�0�`���;]��/�r�-�G.߬�ተ�al/�ǎ!��i�&�ə��fI�9�n��h�	��z3E�H�)H�������}�Q��FQY
G(�}a3��};��b���꟟σ)������ʬ~ͩ�c�/��JY��+ol��&�]gI�b� 9]�m⡘a&ґ���A&s�K�XK�	���Ħ��S�R�^q{ֆ;��F���\�?R���ԙ��gDf/����vP8�V^���٘�d%�'�u(b���bs�U3�%�Q���/�X�"뽝��f��G����u��ُ� #��|������S��5�kb��*�X�(�1F$%Wa�8�,�]�
ۚ7�d^di�.�P8_����˃���::�$�u=vt���:Vh����R>o���@#��%Ef뭃q7]� ��2��<�{�94X+�4��Vm��ϥ���o'Hp���a}�Fd��n��D�b����8���NPl#�5� �w<㷌��������.�&h
h�3I��%f���E���Ԡ�LѲO��
T�t�;�pcE��W�9Ӹ%e�m7:�C�ǫݪ��	��d������ S
�8:s�A
�n�ƣ����ⶀ���U�����'Bܮ_8�/�i��;���Q��;�G���:d���(����D�`�����ިg����VH*tͫqEWS�y���z�Ϲ��j|0��4�ȡu��V��9u�G.������vG�xQ�7�4����5� ���4�+|�$�k�Wн���fT���:"���ڱ>�2�cw퇐L��/|�P�!�J�A��2��
���{�u5��W$l��/?���&��膐�I��c^�pD���;�io�I*���5���P�`�J����~�� ?!3l�/T/ �%3��ی���`��ŮU�
�x�*�I�q1K���k1�@Du�LJ��S?y��R�ڮ�M-�Ww��u�2�Zn�s��Γ<,��cy���E��z���_�����.Qp��Y�;Z,�