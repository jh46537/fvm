��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O!) ���Y�Q΄�O��*Ȣy�dsuQ���`�Q}SA[�.���(��<
vɼ��;4���͋s1D[
�f�T�[��h�K�"HO�¤�TwƜ|�J�tR:����p�#��;������A&�K��HȮ�!!@<Ȍ��VV ��k��ko窿ae����ZS(�F�FO��2�;Z=��t�)W�{yo��r��(�K�StcN.�����s{P�8��AN�C�/��~Y����[#�z�bEB97�'���?�$'�����ِ��ǰ[�'�d�X�������%��`r��`���8D�]�At���w	V�򴴌���R����F8[4Nj7�-���ιFUEp�]c��$W��9P�|�Ԝ��L�?�9�8	^rA�Ƿ���.�He���n0�u�+}@I�2��P%p���-���6��f�8Џb̝h����喥e n/&ρ�1��ue��Fw�����s���Sܿq󀷀�	�~��ݒ�-i�Ȳ�G���S1	�g��<�ד��f�t0-I���:oۼQ gD1M隬it�;y����4_���TB�چ���thh�bL0���]q~�����4�Pw��Du,��8n�,�045��u�3`G��볮��"�W����`�hR�u��yI&n��xc���&����7���W>=���Ű��T��+�ς7
�73�ȥP#�lm��"8:�K4�j��c��<��d�eA����
���&c.�nP�	�hy�Q� ��l54ꓭ��ٶ���j'bz~�������,��������&l$� �+��D}�4j̢�0��)z���#ef �2)AuO�3�ۉ��p���s�l,��p�J\W?��sk\���k��}�a�.�.i]�q��W���o��9�����^+@���T�ӷ1m�$�X��<�j更�UGk�y��b��}���8uw�h�R�b"㕑I`}�0B���B��v��u0ۇ���A@��D����N�Zۊ5&] ����I��-�K���_å��HҚlL#��^�p�wo�O!�`'����^6y1^��m��7���s�5���"����BM�&+��#��_����'k.�A�$ʎ����ąI�4Nj�^��Ⱦ��4�e�zg�J �Ty�hL�%� �@x*Y�B��2��a�0J.�v�P=�|H�"*���J����6ttee@�`��v��A�`�
����:�]k�5ߋ�#1�m)���✶��j����^�n��p�`�������C���_t���Ḫ��f���S(���R.���26ƌ��/�[?��O�y2��A:+ζ4����61q�o��������	�'U߯K)�k����f�貊޴,-�i�@��?#Ɉ�����=X���)����'����^�05!�L{*껑h�!M� �$.K�wg!z��|a�K7S��������ސ�~=
�@9N�2hO�N+��S̖y=�X�W��i]/B�1QE;�EI���e���.s	ӭ���a���|��Ky`q�� �}�|����2Ŷ.h a�/V�'�jm�:-�n<
'��Ls���P����f!Ν`�D'i�#��硽`�0�k"�s��g�����K[��N9��D�����QGMT����(������*, ��܄�A"�v7�S;�R��zX(��؋Xpw\�j�W��o�D�YWguZ�B9�g����G���с�z�I[خGx,���G�C��I���qo��F!ױ65U�����R<��RԪG+�o������u����(�O┷'�{���Θ���?���b���p�����Q,$�H8�m�A�^Pj���{=M���>B���3ڎ5v0��d/i�s�=�?5z�؁%�+����>!�0�X���[=�j�֠�`YJvY��H��EP�m�ے�y�(;���:����Q)��g�x|1~%	��:�0}��K8���e�}��A� �&�Y4JWBQ��Qő˪E�E&���W�Y�`�����xA#x��te� �2�|��͐�tC.���׶��F�N���P��܁1���U�;L�(�q�E�Vy��d''nm�n�$�&�vH�U�A������Ɗ[Ja�F�4 �|VR������<�ϤI`�<��F+�U;�e����^�ix���V��!@po�v�"�I��|C�uǨOI�jI]��Y-�q����;�)��%C�[�^'���c��U��^=ظ�uD�സ�9���N�i�Ƽ��'�*��c"��U�a��� ��)*��Dm�t����t/|>�멳�S����K%����\���V,��}�?'u�R|:�M���t�rFG����$�c�\DH��8�̕��ǝ�y?D�W��!w�U��°<��� mb?g��n1\�ݾ�9�����m��O_��'�Bq�U8���U�s��g�`\��m���0�hC����I��b+���D&i�Zd�c�/�K�-e�濼�
h�����Rt�x3�EQ ����ԮT3n	� �(�jVH-��u;�]��Y��hN�T����F������[����VU�Z��Ɩ\��qOS~5�{�����$6�y�w3��lڄv���v$�
tCU���lF�h�X!Y�G.�p�Sp��m'Ȫ��>�:�ڙ�|$�Q�.&KK���מBH}7B2OD�H��泪�l_ v��F�  �8Ҧv�1���e2����ಡ���}l	�E���1���GY\�}�iz��_��x�6�}����j8�*�e�fUiT��O	7��= ���GA��#R���%���w�XJ�4sH��lH�E#�lƘ�`
�\C������Pf�
�]��&����Ў;��Y�W���b������ف]��;}�W�\!�<��,V f�"�g�7���#���YVEI�	�M|������okx{�w��_�[�nKZ'+Ӎ�[�4����A{-����U�b�ӘH�i-��5��N�U���R�d��[S��/����z�?��n�&������C�����F�����㛾�+�gQ'�L��]��LW6`b���Q{��$A���|V������ ���n����32����xX��� e�O8�hPx<�$�n��889Gi����T����!=��W��D��l�i��l�^Gv"���g����u�K��j�K��_r�-��}Q���@S�W��l�����&����� ]Z��U�C���{>��D��V ��$Km��jR��/L��C�_5�nW�@������)�D8D=,Q�}�~\o���!�b��qOw�:ZV;���.|sM�A�Q�X^(���TOԓ�n�e�*�z�5�����,��HbW�)�b�4D'VT1��6�Q뻁ǈ6�uL�z�qǱ�+�mf�9��af��:�f�(�ԏH��6��g�=�����Zې�%#W����Y#�r���9ƫr�1�8��8�s��"o �G~�Q�"O���K��f�FƯ�he|M ��M��Lֵ�$camGܶҖ�k�B�m�A$)����R>$PZ�^�3|܋g�N��K����d�RqL�!�1
�1����3��#MfMa)O�u7Ԅ2��ޢ30��c}���`̬A�VAه��2����K�8�����1P�b_+kV����R��嘽Gޜ૵����]:笉P�g4w�'y�?A���������X<�Xo4�Z?x����p��*����O�f�8ȅ�f�V���¸o����Z�N���UsV�����ң��o{/�=�� ���n��0����~� �A�zs��J},<�J�J��E�Xkˋ��`X+ Ϗx���R~���|�zo������k�غ�0�9�X�#޽��&m�o�}Z��N�APC.���3*�/�L��u-F�4~`�����)�yw\@ߡ���FG�G3FѠν���&��s���	���i6�@����_Iø�+����A$��Y`��7��>��=�r�Z<�IBmȽq\�V�Tր�V���D�@ ����=���ZO���������-$z%D�;�>{_x���+Wi�~/v����3>A88�M��J�al^m�dH�M!�	�gC�Cc[QdV��8�(�$���TX�D�P9ҩ\Q�|�.��Ƀ��RT�dЪ�G�L��aO�s�u��>��N�{hj�Cצ�iS�L�u��&�I���ꟹn@�g�{]�F_'5�K�w�� ��1g6��'~~�\�ո P<뺜J�� �v���}��ba���+%��R>N=`�sO����|�E�=pQ�5��o�l�������!}�ϲ��Nb
����Z��x6\�T:R�Ƃ��p�-��P�$9If��c[G�c��S�zMe;-y|����-�v��2�32��r<�w�'eኁ^��5���J��V�+/��HP���^3<~H�M�U�i��R��
m��VC���5a�9Qܗ�+�wmٌ�C��p��Qj��I��&�+ ��>AY�`��[���u':=���Zv3����/��~�d\GL����}���=pn��lI����'�wP��W�o��[����%gL0�� ffA(�7]|jq�h�Æ4�3�Sx�؊���>�[��Uẅ́�f6x�$aw{Q�2>#�U�q���\BN���d@'�u�(��	�#���+�m�
�^�4��Mv��T~��h(_�l&�z�{T���ڪ�e�'����|���5�r`�syr�/<�p�w��+�p�J~������ȝ��$�b���߃*|�kd��TdK�\u�e��%���r���{鹅K���2��#��	�l�ʢ���y~J�t@��B:d��Pcy#T/>J=)P���m���і���L+C�| T�n���D�k~3���[����!��t��{�ٓμ��a��lNb���)>Q�d?W��W5�Jdd�i��'�F�U�����g���#$�Dŉ��Tq����e��
����1;��m��aJp-�d.�s�ќ��<�������K��'�psU��[LW��	vG�]���>t&�7���lکD�J,�Mbٱ��k@�Na;��ቻM��Tp�b����T��'N# �x��o�4�L[��q
e�D�Ax�z��� QIV�g�ÅxPQC��a[[��d"��W hy��꼄.��8A�+ȍ�W8���e�k!�B��
�T�0Ό���PdxL�j =%��FYr�P���R�f"�<gÊ>B0.+@'(�ڻ�/�5���f����D q�સm�N2��<��������88P�E2���`��y2 SP��q�{��@sw�2N���%�X5��E�qn�+WQWx@��U�/�5��qg��)�D� D�3KQ|��ZP���А��R�r����]�|�=�e!�<����o�S+U�)emk�B��y��S��镻D���쁏�Y?huA���ʲ5��/z�iUkU&a��.�Y"�Ӣ���햣�7��"�+Ci�9�{v�\{ǭDt���o9U�ʮ>���(�!
ëDލ6�؆Nž<���{�S.��m�,���º���x&e?e[�b��<�E"���m��:��ȋg��0�O��q�V�5�ՙ_�{��0�{?�K�Hz`9����,yB��מ_��\f�َ�<5�o)���U��?ϭ~��cP_��nCo5�4�~�@�+?�F��f	� Z���s&���77k;���s�5eβ�ˆ�����P������sӲ�1{n�s,X����PRg1�f�2�DX,��ʦ�{븓���<|6�J�-�E��%�V~m�@�Dm�~�q����址�%��? P�Ob�Y�J���^tf��ۡ�o֊&�����Lx�¦��=��T�(;y��o�)հ��p��R;D��wc�~ZӐ{����Ӗ�l��W*�!=�~	H���x���������Q�A�eH��;�پ���F[T���o���x�`G���1C���w���eaΣ kE���e�+�U���7W�y�x�qB�;�?��&�F��c9=<ł]t��0��� ���'�<�CvZ]\�&�x���P��q=UܤWJ��ړ���QG���� �w0Ŝ�#P#�%u�d_ޜZ!2+C�Ĳ�b>aVr-uB���i��Y��6�,y70^��!��J*��G)������6s��圌���B~�Q*�X
�ڊ>��N�[��H]�W���VL1�nܴ��̴�Bj�`��Iܚ�S�7�c��\)��� ��q�9XeXt��$�������X�����RK�Q(g�0^�S��U~���~�ZO�+!�q�I���ړ�K���ܒus?H0@wA������<7�����A��29V'�^���c> �U��)$PE�f�P�c_��'w�D�v=u���HX��C-�x�S~�v��^��x�%c��/����l3��_��8H+�����G^{˨7���FjѢg��"0�_>�b�B
����������n�fm��� ֘I��n��@���X�E���`�*����VK�ߝ�1n�:+�ں�g��9j˯qE���4�7����� BB1�kJ���#��������ܔq��G��'�I$E�|=條��b��:��Jm��'#*�f�i�8_[��5��I��X���1P* h����y�!�^�$�!�����.�%W�-3�Q#�;(��𡵹�P���&of�#&��@����m�����r{b\^�"�@��)ȿ�=�K&�.�}FFpʇ�߫��O�?���*
x� �;�Vk�Pt����D��:��{��� �ޯ�QO̥Uh�q�{Y ��E��M'���L7��%O�i����r@�0,G�Et�o����]z5!�6��.���ۘ��G/���S�|��|cٖi��=P�F`�ĬiӠ�����̙����S���"~j}�8�����K ���ׅ�1�����e����<��4�X�顅
*��n��i[���JR���/�c�"#c��������=����-�Z ,��x�x>�N�eƎ����7���HUz�6OG�CJE)�ὦ��uҜlDE�=4"��;��?$���{�_�V�����+�!��ĕ֣3��kj��8J���v��[�����u�2H�	9b"�����.�V\;�{�Tc�j��ҥ��\iޚ�C����:�k�W�ׅI���˵jJ����9*�E.o!rJ�����˚��;���+1Jz���z�mh	�2
�3;<��S7�&Р����U�tUuO�m�@��HN���:��	ld�&��l��� �g��%���`2���~�n��gK���n"��.�H�yK�v��GO���f46���_K9��\�Α!����yp����l�1{1�Z��'a�r�E��{&�>�GCz'���Ԇ����E^�f>%�îZ��D:{�����4�a�e�����@��0�
�٬^t�q[8�ۂ)P�?��pa�hW��i������Bdo��);������=�oy��zуY9ߝ����$KYqB%K:�}pZ(DL��ݐ����~�l4�_�U$�5�/�(Ϣ.Y7�\���>�YQʖ�b����w�#������{�l���>���>U�ɢ��S7�'�)��	̂�v�G������/����6/��G���KV4�?��Ϣ3C���=����E�0�����L��F0��W�yp�܄D�5OH��٘Si��i�,ع�s:��C�9,��`o�pP� �Gr$\��_2�d��@�����+̩�]VS;�5frOu59���:$s���Z�/��[(x72!���y*��IE��:��fz3bŤ[�Pi��
3M��F�;)���6:`�Q���W�U,X�����&w�}65�zU���u��\Z�8��5�~$�d���NUg�s��Q8q15U]WQ�wvzd'o��G>6A����U��Nw2#3��1BO�|�A�# ��+�T��z�vI}.��!���ξ, �d��}���wͭa��߫2ņv?S���5�s�dW���0�a6���T��CY�I��
F�c�/���/�t�7��ǳm����rCc�"�J/|�@�z��(���e(���/F��������엸���\�����a[:h�]�fAM���uXւ�<!tf�����ǀO!Ԯ�C����,��=�����;djq�u��B\���sB�8���BC���`���Z���BpD��3�b�)�94)qn�S��q0����g<�W���ؙd����k��+�����w��=H�*3��9���d���į_f���7D�fW�m�o8i����61���V�D�H�`���g�������pY1��p���v�DФ�L(���먋�O}c~��3jv�g��rdp�X����ďe�~R��4伅�bzXQ�1 ��G�ś-;ɺe�7a$�}�"��{_�>ۿ�W�*��8(ձ�>z&t�MD%%B@�䃗�p�`���[�Eɹ�x�0�L֙��̾?��S!g�+�7��=��=��Jn/Fj���eRS�b���v5\=�(NH��-��.�'BwG�<X3z}W�l~��t���±��9��3
]s����W�� �E6u4�fK��(?L>�k����L9}Tnm�x��u�'�X:����B矗Z	�gs;o���rw����������)ԃ���K��W���eԃ�k߻��q�!�6�Y���������U����#�sF�
�y�=c�,Õ��)LK�}�P�.���]aF.�6�ˠ�O���w��4nL�<0���R	�!lמ����x�	���~�\ ��Z~��l�Q�}�0@W<�]G	Ds��@h�ޭ^�>�}��o8��&b�~��̃��!կ���q�>:xD?x�h���i���mB�I+�B����oB�>�Or��سb<D,z���*1�O�I���M�꒰H�qީmB���!�сS�b5��à�����y����u޵������2g�@��^� �����mМVѾF��}��$�8K��N~�vO%�|���bq
�?�+�kҶ���#0F.������So�9��Οvٍ��͸��<�I2�N%aE�>�,�ɂ���H�}[<x��a��t
���52��U��V�[sE��U92jN����i�S�����=v�	��0���'�����uH1��yY*���]��+D@xh-�G�?=�IV���JAL
��U��61�b+p�M����&L�����������Ǻ࢙2��&���K^XL	�ù�I�H�C/����K����_��9�'I�G��0c3��<^E��j��s�������)�;�ِ���H��E�x��x�OsL�0���ʲx]��-��������(^���O�����g|�T ��#*|��e�|��؁6	!�b���y����U�u��zW�9$��cVA�&�%K���kD�@W"��I�7��w5�'���F�[K;�~x�3�3�0�S�$�x���R��B��5�'A������@6UZ�vwWVVxl�s����%>BI�i�)�*��o����fA�v�� ��O�-i�H���hl��~�IJ{�[�x��?�<���7��_��
�?��ལ�i.����P�N�x'��y�����H��H|9y�w���K��9iː>��_�/{���,�/��K��C;�g�u{�� VG>M;�!�Ue����G�rjp�L���.Z~5�540�&�S#��Ո|�e�6$�v�W��NC���٣pŮ\k��~Þ0�umx5�k��x̲��OFWL.P��K��F��7���������TE���on&�|�z�P����2fdR�gT/:� G��UU���C|U��"����@_ndj2�A"�!���9��@��ֿ�ǖG�h/9ۮ3=��K0y�H��)ɽE�8˓D
7�e�/��_�mF��бS��:Z�	�0W�ew�U��8���c,I��W�y2J�qحz*��͒!{�Dp��q,�H�*S�C�»�}�y����ӗ�sDl�TCu�LnF��q�N�{�ԑ�M=�ݴ��9�-1VY�����x���g2���Y���Zb�=���{��f��/�I��|.���O�C� Z�˜'��֓�/�����&�DI�/#���0T~e��(ƺ3�Giex�p�5�W�-[	�{���D��?aa]�K}� 3�� zMtW�c�n}`��C�� 	��4�ޣQ}%p��1s��`n:�r�� ����{Ț�$KW_�D���J�-�n��a�Kx(�/2#c8��ކ��k���%p�m�/,����t�w�e�!+T�UQ��{�n��LR���/�n��PU�ڃ�!L�����2�%���uo�0�jU۳����L��2�m �+o�.~^����]4��xy��X=b���@�}�r���2����<6"�
n�@��F���Ȣ���U>tƇ��B[gwi�r8S+������I=¶�\�$x���BJ[=ٝ�ǽ�a�nO��
�������P�Eܛk?�����(�i�"�cD�B�\8{�[�,�C��@��)�̓3?��9���f��շ�����R���z/0=�buQ<M9�ɩ��O���)��P՟.A���9>i=�vt{�*��˂��;Ͱ�76��N��ܡUݷ��恑�a�4@�5��E;2ˊQ�h�6�Z���m�7q��7˱���F_�b�,E�s#<d��+FlJ�x�Z)����"���C|S��D��Ƕ��B�p�C�'���&
cn1��X���)l;FH�j��MuĲ��SccĹMtۏ�L���8�	��gHYO<���Z���CA�7Jy�x���X%�9	�͙�]����XBv�I��_��Lac��|2���!D�h���#o�zCb�a�Y��E��ӭ(�z��FT��8ғ��.�r��W��2����V����/|�Eh�3���~E��X�dT�����7n�`Q��?�{G���|킏�ҩ�U�M��*Hy=���0ݥ���[v�#(�>��A�����E�����aZۺ���d�[nVAi��KƲ���6�.��V-��xr/t��'r�Q˒o,��e�p-�� F����x5�C�3KRf��ܮn�;�8��jVW��v3�ȵ�oLe.�BG�M�LN1��]?��'��L
j4���E	">��wE�@���9��)pČ��mϐ'uM���-٠[��)�e{҆���Nk����jI���= ȷ�q���npH/	�8��[M�*/��S.��l�Yj�"���vJv���X�S��/s;���yQX	Ad�rD*B