��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ7�V�>sx��������������
�?�]���yQw,�.�����3*�?H�bY��w�\A%
YK�#��Z���E�{8ENuM��#VU���vS��60�Л���啁0S@VUv�ȲC�r�d�wh��J}��t�^�qt�/g��7/�3:�?�n���3��O��:ά������w ����˹=|���~�C����3��I�Ty��NR�M$^��f�wR�m�X(:Qpc\�S�7#�`��)e"��S�ޡ 2--� ���D6�@���!���d�-�����\Qi������4/q�;^n]+xOۃ�t� U����j��G���Y8	�/6���KJ�£
]����,	|�;,���)� ����$�'v�Џ�ҍ\ms�k��8�o�a�V�Q�f<3k��|
�Ā�Z-Ժ�/.�)>0��j��\�����Lg�P��#c��?N1����:|�ۥ]�m��_MQ�����e� H÷��y����b�*۾q��0��Mʄm�Lh��dJ���ldg�wnݘ�72o���/+��'H�ͮ��}C�n�rW+G�c��,�w�,{�zQ����Z�n��1d��a���U)����:�bxyN���	u��k�Tp�Թ0�0�����W�Z2�\7E����r�%ұK���{>^[��ETB S��P�G"�n:��$��o
O����[�hh�Q����փ��t$F�n�Cպ��7�f���A.7��<
jͫNF"���o��Ù@�7UXӵr��Z����;�K"dwPz�$kJ[��r���+���JB��Y���.�<M=N�����c	�?��W6o�uj8�k��F��R�T3�Q�e�_��Cue5.Q��\�E��|pC�Ʈu㧰�#�?V�d����-\�{�JXH_��F�Ý�"U�k��TZpb*�$Y�
������厭j����!ү_�Ǔ4L7Q��[���i��j�/a%���T09��\��ufD=�P�����)5>&�$�ǭ߬�Q-�)j���& F���GE�H��"��䅏8�FN� |V7ͮ¡л�
�ElD�x ��/|8�� �<�=ĺ��ވ�o@Ӑy���*����T5etY�n0��C������kfԒ����`;�⠙:m�A��N���V�0�����7��;���3��#���<����$0.���\
^�*��E�^��qi�`��H���%���=�)�p�^-�a�A��~�0*:��0)���D�
�#,�j�+WZ��Č@D��{��)��R��4�V\��7����ɛȐ_*��O<�N�8�+��;Q$R�F����1G?��������C�:����v��_ȂM�w�5��y,|��(��
��V��ÁNI,uϖZ$H�j�yU�AVn�¹}��R5}=��y0ݹc����s�� U��E*յS̸��gc.�%H?E���$h�yԺ�[�����C���S��!XC�W�9g�䑯/�M�8�e[2⑏���t�Cf6�/\g9zi�p ����u'�\��K��2ն��u:�)�g�sX0�ޮQy�PJ!�t�ÇZ�h���j��	\%�+�3���yN��>��w�L�\�h'c체����[�mO���׼������҂P$g��J>�M�Zx7���m��=��{��� �>{�1���6���o�3�K� �)nҥ�p֑.��Ѳ9�!���]ʈ�-F�a�����f�jK�q�!���;��p��x�չ��&�c��$A`��Ĝ�jj�R��~��2@䐕[ҽ`��ɝ6���6��9����\`�}�ۇ����p�;`^�m��A9�'K�:�*��~X�� +`��1:m<�2�����3�|#N�+��5�~�0i��|��Xs�j)~&e"��Ѷ�I�f�z�A(E ��t3J�_��=���Hz��"IC��ז
u���\�cCFx4�林E���.��T���WD��9�S��'�.#Q:��' ��Ǡ�F����1b�b�4�bE@��� �
e������S�Jb�%�p$c� A�����ժ�ˀ�nYع�׽�$ь���)�N�����.2n���%h�f]���Z6�� ����j؀�m��A��?�q�os}��B�@��΁��Ռ(+��C8��@.Ey��U�X�D����0�bk��l����75��Ԣ���I�۬�\�#?U���qюǸ�	��ظ��*�ř���KE��,w�%��{���m�f@��>UqE��y�,��d�\K�&Կ"M�ëMw�x�� �cq��s��t���ǰ%
�L�=�r�q�56��<N^���_�ܺ�^�R�!���q&)�E�<���i���o	)��Z�7�^�g�kѰI�&�������0�?�੡�,����H�,�B(�Fʛ��\Ympߙ��"'�����M��6o!�]7������|%�+�?t�qM`���\	FOK��&�u��-{�5�@<Z�b�-o_Q��b)��0�b�����M�T�R�0Ϫe�1�/��{�o���|�"����m��hRof�|�=GlK>��^n~������1U^O��m�qi�As�W:�`�"�z�m��b@N���䳺D�@�t}��UJ�fik���g)S�E�y$��m�gsΜx��M�l}�Ҟ)
iC��җs�$��L��L������z���@��g�;|?"������� ����|�o�j�}5=N{Ah�:�\�T@b,5$��~�8�v�,5���?�RjF�:��'ޟET�~'�zg��X|�%Z�2��\�G�6�He<�J�v1�,��;bA#(T�w��GxVĚ�n�cġ�t�K�%�j���w��b9�'��P�����z�	JI��wN���ಐZ����P��/��g�D�E��R����=b�Fiv���F�4 	e��`i��k�I$���.J���:^	o�E��@�E��S��Q��F�֘�l�NqL0�j�p����T����SԺ{�ޏ��Tb
 ��g�8�W�T�T�lF�P� �Aw�Iz/�����~��7�p�4�8�T�g���L$^L��UP뎑߉2t]��Q��lO���ď7�ί? ,��
Y���� ,�zeG��]3G��
�c��J _�E�����ҙ��BjmZp\2W��s�
��O_���-�4\f��߉���#��4�^>��R(r�rV��FИ�B`���@ %����ө�բ��,�@EG�K�z{�$�<+�p�c���o^_�����������
���(��v�t��������6V�8&r�\-�m{�%�����=UR�i�t��a���!�dK��D���\jL�tۇNQ��K�A�x����8S��Is��\��~$�*�m��7	���C�B-���A��m�ῲ�2H8�\�3�(�* ���#��07���q�KT{����N�2��gR���%A	ƚ
o�õ�7������l��馇D�v��^pRL���r'�E2��1f ��>L��x����7"�K+S����6���f���x����y��og~ ��`��F?��F�YF��<|�T�׼�݄�L��빡�x�/���\ �%O��$��B	F��C��F�Zq e�����Ò��ZC�ց�bF�d�e�|�u��7`2����/��aQ�,���\<�À{�����D{G��ȉ>��W�}B��,�ǁ�X�ؒ+�eiU���T5��x����t����S��� 8qt�ۢ��X�ӥ�Ap��t�Y��C��do�!'�PE���	~�x�Ԩ��J)���n��{Z�*FCC�����=s^D�U�#j!�b�dK���s����`����Vgd��nL��=QC��fk8C0mJ��D���n$�#E �#���J�	��x�CV���1�e'�<�G��\p ceT�ޘ$Z��rf�w��)�ł𤋮›�����Au�z+�oϊ�EW��B��WV�1o�d�L�V>�ʦ<q# M�'Q�spY���7�G��-ZM�d�I��&�6mh~p�R�����B�F���;�̔�ꘊk�����Y��_B��݌��{��.�Kw'��K�hz�6
���fx��%�]�0w��%\���x��/Kf��s�@fJ�}�F»�H6����7O=G�t)�<�4~��2�Z���&W�?O���16��%���q�N���a_;���J��kA�*�{� �Bs��9�����h� �q����8Z�`�Id ��p�{7�#���=��qB�����S��u��x���5[@\Jq"���	�󲔸0k4��e��o��%[���-��=�|���S-�����a 7�u�������^y�K�-0E\���k���~a�c�VE�_��4_�S��C��ȿl���Ĳ;Y�p���\	�܆%����^�\
���@2$ln6�KFْ��7!�;\��5Q��C�F�\���.�E�a�{K;�^�7,���Z次e"+ ��y����P�Ҧ�F~���Ur{�@\���Why�ބ���n��c�E!Khݲg���@���e�Q�rkS�(��^j��nvPd�d������b]�a��~�$`�',�h���k�Eb�U{$du��"9K�g�(>Kk���U}	�`!li͛>	IU�|��-�2�:{��U�4ͅT��}��W~�Q�`��d|�bBv1s1!>�4<dE��ˠ����E.F	{BUoo��D�%
֕"�$�}EI�M�M�]��g�r��P����?"Xq�X<�$2,�Ċ��i�	��6�(����c�fs���o�P<#0����ٝ�lI�q|0}Mv� �)'y��������m
?==��Ίt���b�^���Ow���!����Cz������2��G�k���x�<4\ݛ3Jʣ5H�,��*�I� qZ:31�S*:��~��cT���&&�]��o�Ѐ�5����|K���/�"�41\O)k��C�6��]��ng��);��%��PYd��u4�]E��Ǿ~r9�t�I�s8���Q����s���`�"�3������� �����#�^����Pe��`Ah�}$��°�Q�LT`�'���H�f�"��!��>�9�W<�8���Wj���hi��{\4o'��͋i�(��f��vI��ceuN~�����+s�8��K��*N�u,@,�b�"
u�g���j.���Z3�ݎ����*�$<H���3* is�熉5
3x��EM���eiT9�	��jx�8��JzE�E*8�W x���9���!qU���*�.
4���m
�� W��[�\63D��I9D�t	��SP^�9�Wu���f���y�Ȉt�"%A|�����uP	�S7�v�� x-4 A��X�A{��N0�����$�����޵?{W��� p��3g09n�tRoJ�}��8����4�����1K�s'���/G�A�J��:�@��Ͽ��b�騬�tX��DQ����q9���r$�����zk�����uA�_����R�����*�׫��j斢`����šʆ&�|��o�cZȡ_
���}@���f�5
�>{'K��J�x�� |�K6V�-~�8��X�7
��2��s� Ƭa,�'9\�%jd^0?���N�g�G��q��un�o3� ��3"6B26�1�;�B���-yU���z5�ı0�G�Ǒ�Qr�Ÿ�?�ТL�0hD��e�y��-`�5�xBg��M\�+R|� �����R����댦�$��:6]�%'�6wU����f�5-�e��|���̪�=�>���s��d{�Ag |�� d��c���?D�1�-9'4�� ~i'kӸ�8%�P�s�+Ks&qu*�|YGu��R�/��$%���w�֌h<�jF��G���==s*���Ļ��4�2C���F�|Ԃ�װ^dq�;�T	�e�:�nyl�[�	*���!_w����>#�����]�8�,u�k�NiZ
\�9	���~T������H���*%0m�����	��|�C`��A�[�"g[��u�����ҿ�B��ZSʔ}�=�i[�t"��N��d�a��`���.C�ܒPH�6�E�����`C�9���*�h��qME�{!�:����-�X���;�Z�{���]j�b4�~�Vh���g��������;���]�o#0Pܙbs�`�r���0��STw�����8���Xh�����	4�ᐽEF�̼(a���<n�E�j�;]3r!��N!��<��d佞����@��q��KB��	W�i�/�qB�Z'%�����լms�g{0�9�pf�>F
ծ�nC`{ 5Q�U,��"!BR6n}�tu��|{�׮`���̅ɳLM��'��������񆲈��~��R��f��7�q�	���؄�H3!1��pE׆�@l�����1�O�a;�;nŏ ����{.��@�w٥�#'�vʿ�k�m����\{U��|{���v�K�m0*����!���o�t���"I�!*w,(G�q�w�����T�a^�^�I�H��u��TX�v��X�r7���ȴ�G�-��ndo�����xJg�l�K\��H*8Q�����#R��k����[���*�"���Nks�Іz�G�A��Yv�/�K�>�#��Y��\��}j#.s�d���)�]�������`Z�Y����PK��c~��4h̩ᷠƒ>y��������/�hA���}�q�@������XtWd5��Ȓ�&]k�-����/���L{;�d<vN���{��Ib�w������K�j����p�͇JzB�W��}��L�~m�#�ִmP�?W�H�y%���>�(@�j=<ϟ}�v�h�N��/u����U"bx��ևOB��G���O�GO|�In�������F�+���5�H�e�u�^���b��ΥX_Nq�k����8������$Ս��w�T���9�pV��uO�+����l���VG����w1�� ��M���W�0��:z`^O��m�p��6�� ��ك����H��ʻ��N!; Iiz�5�$��i�y��~l ݪЩr�3M]����j'�	So����Zn�*�Ā���������� ^D�!��٨:Y	����N�:q��4�0W�p��	���_bC���V:a�Ȭ�|n�T}����^��[8�]cH���G����[�q%s�}N��>z1�І1ކ������/�g�?7�]"$��қ8E�&�;M���ۆEh�;��$���&��Um�8��^"����zS���L���̇�=L��<��.��QČ�&�;m�f�Ϻ�1@H�x�e`�7��Nۨ��U^g�e#��Y`�S5�l{�K����+
�rT�V�6�N~���bm"^L��$J��Gr6��E�ӝb��dO�s�����US;��$
z��|#����M��b��K(�xi��F����3�ܙ�������J�(0���%]i��W�K�կ�h��A���-dvw�CWX��L+��Q�17L!
��R��)]b��+�����ns�A��/��2礆��/6���y�q�zX��-
<y@,� ���u�����.kw@�~l�bЌ�E~ʙ�}|�2���mK"d@���o^�O��+с0MFX_��:��j�?��a�S /9�fL��Q� ��F������D�d���KΕj*st�\a�~O�Yr�@�3�m~�w��O^������7�J����Ғ���^����|�Q�����kd�s%*��L��
�ݧx�U�r@���w�K+V.uW�㉲^S�����C�1'C��q�ʒoG���.���T?���[]��_��XOB-�Tc+X Ѱ+]�È/���bE�m���6�j��҇�D��i��<_���3s������LC��;�I����\���Nߢ���I���O5혐.�5&�]����h�`�	�Nǫ����o�u?���Yi����D�I �~�^g(&����u��g��J���	*�Y5�e�{�j4����|�f�eHu^l(��nMt0�=��h�v|�d�q���\��cg=�wR]Z�ϪE�qIrǡ�gp���6cMMZ�z5)����*�o�k?���*��/�,׾�?=�%2I�]I�ҙL�y�IA�}=��k�"�bD���ФmR����p	�?���7!�e�_1�Q�����)y}@��%�h��.��I��A0���q���2H?͵g��������cf�>�a0F�5����pa}u�|��$�����ف	�pI��7�!����-�[��H�g��!����ȝx<�N�v�X�� �E����!o���߷���<?�"��l/VRd�O�"����	�[�t�(Q�m�g@I}�[kȽ�<�<S�{���)R-�X'�uX�]�Bܺ#P�!I�e
B#%�����g�y��І�A��8�0����nW<o\M(��*t�$ @}��Sl�#A��~���F��4��!Q�s ��E!�Q�2pP���w��VS��-F��ͷ �t�s��h�؋��Lӡ�0���̠�xL�� ���v�^Go�W��d�oU��@�8�z���=�������;�ERo.�N���B�%���1J
�s�Vxs���޹qB�>ʢш:c���ۄ$�=�\cr�bi�Rxn�!��L��\��(�J�?��K� ��� -�.��՘5d�2���!2^uu����n}K,8��o�L�ή1�d�*�Ǜ�Qb��n��$j��Z�H�)fW#�υ9��J"��{	'�c�8$� !�݀==xY?�մ,��<Ε�m�J���}fG[`,�T�K_,:�#N�y)r�I�@A���w�h�R�zGis�M�-�7S�I�)�v¼F�Zi������^���6�Z�}
_�� y!&υAx/T
+�n���X�Xٖ���s��j��h#��8m��P�\�]0�3��.���ĭ�����x��:`k�Zq\���cw`������b����,�f�@D��l��y$mw��F!i����WCD�`�F�?�Zb��b����Z$B�VC�ہ"�m�b���y^[��t�}��Ǎ�K�64eMs%ʓ���<qڞ��)���H��^�Ƀ�A�y����jf��eS�(�7����=��D�����5p�9D���c��⏬wã�I�=�F'�����G���~S�8S=��=�N(ղth#DN�\G9�
�Y��=�#i���W�భ6��Ea��0�GC��!��r���u��,~]��C�bM�ݥ�ϕhT��� 6F�����)�;>��2(������#����ny��p��FR�-��p�KOc�a;��w8�)ںؒ>�PJ&��l ��%�[Ewzd����n{�х�|��l�&�������?����ZIr,�K~#����i�4gh���nK��U�c�%��
W�4����b1���u㘕n����R�Al�$+x���#��9�$��88Zp~|i�m&h���c5pX7����$z�9Yl+̪�jp��,�jv�̝8V�snUQe/[՘��w�ڡ,i�����idX"���ڴ���t�OS��d� �O�3�WJa�^�j��^8�X�%XEFG������h2HŴ�.��>\h,A�� ���g�|t����m��})49a���˟��OE�Y�EC�j٩�k�%����ܒ !���kb-�M�{;�Na�Q����I�5��mx�JX�V���?F:��G�����]�����S�q+�_MnD���t��x�R6z3sY����K���m�Vu��%j���t�Ee&b�9~%r���2;;��еth�h���q�r���I93դ"����*\�J�]�,�?Ԙf�����c�r���p#��9ްz��S6����H�'��y�F޺�
��kj�@�����V���"�j��=��d�a�O�Ҕ�T6\��Y�F�S�h�*�R4Q�To��l3�`]&�2�a
��,G���G�]��g��5�T�\R�!.L�\�Fh.��y���*�ty�h���"�&v^?j�^>9Q����Y�hE����Oǜ��O��e�׬��]U^T�qaQ�#�,Q��^�w��ɑ��EQ4�Oy��qa�)(��9�_0���?�<p4B�<��6R>�d��넞���8���\��Rs��F8\����$н�P[�bj �u ���Ӗ����і��s�oaӱX��-=��q��=��Z����a��=��x�e�JWIX� �g�;BO�=^4���K�A�祋�H��qԗ�=
ٴ�ь^�?�8�p��IZ��aK&�z��a����ű�,v/�﫿P��!0{3�D��l{���oH��P��pu�}]�����	M�eh�V�Na��)w�ǱZ3B��RW&ͫ�T�J���A\\�X�J$�,�2ԶD�����2�nqK����c=O�<�RB4�7B�t���!���,{�z��.����=�:�����WU�G�ZV��y\I��od�1Ʋ�Y��Q+�f_S���D���>,'t,+�] f����=�Բʿ1IV#k��	vιQ�-�#y���*6����7N8S]a~*�L����4W-'��R�'좓���(���]�X�KCa�5�WB�wڪB�*a-�f�����|��"�Ǵ��{-	j��eTv��.�5O̶q7��M�+/�{J�UD�s��L��β�Q���}���z�j������%�7��a�D�c�zx�>�Lq,/��#����.<��pi���<i�'y��F��q�J�i!�������P��i���ӑg�Uj��ϹH���BM�Ax}~e�MLr5���LI4\��O͒I��0Ρ |�~�'�+�Z�>����ҍ���'�M��U�Ѕ�ܼŊ?��}���Ƥ��)	����W��k������"�j�.�q����0| $̑Rq���y��d�f�?���O�B�E�����@#��~��B��HK�F��976|Z�5�V�砧��c��.���8[sh�Jh0�"tV׏tt���<;J�B�uP�|u2�<.��<��|�i�a$�(���i�*��/�
���]�֟�$��2P���q09�}�i��r�6P�@ �J�EE��������.��B���Y��N]Q�$�U��R����r����F�A2��s�=P������Z� ��)h�e~�"��"�F����RSh�����[�Va�z�JZm=z%���^�hZv��cc��3?T��١�.�f�0q	s�kO��� �m�'�\\��A�X���1�+��y�� �Q��Z[1�Mu��z�O"������B�>m4%^��9��v�0�ӣc<�������ϲ)�P���JG;qԫ��˗U�
%��B��s�\~g!�MB$^({��2@N3C�=6��=/�`�-ƥ�A�m�L�p�Ih����%�M��mB��V�n`gI������5Kh`�"v7�rm[#���ل�MQa�(��>u�
$3���ͭ׮���G8n2�S���sY�l�Z~��L�$RM��~�3��{/�\�ѯ��;X->7b�e���Z_]�d(iڐ�M�G�1���+C�+4�b�6�N��?�Q�wI��"��ނ��2�{z���"S>(d�ع�hZn;�9�������o�� [�!�E�^�눺��pB�R:�Kb�2 ��u�(֫�}�e�"�Q�[����0���Z�#�HEaG���>A6W�Z�pm޻_�j�XJXR�)�"����N,��'&�7�����Q��sy��q�F�6�$�e��I헗���g��8�^���Şx�d�_4�Q����]��4њ��-_N¡#���K^��z`�Ft��L���ѢX�	�9q�@�h�$�q\b�a����D"���#d��B��u�.�PZ�Z�8$լkj�=��8�������_���ܤ�!�d9���K��z^����?J�,U�̋T���g�U���f�����I�[1r^ ����8�V! �8��E��E���9�/Yǔ�����s��7>"G)�r�Ǣ����@�Z�%L��R9/���G�ͼ�e���D�HH `:��0�e��Lv�c�f��ֿ�>�*a��C�D�͵W3ܐV�x�&��+BMc�k4��H�]:��ٹ� �v����o޵t͓Rq)�uҵZ�wab�����X��i�(f~�'ճmf��x#+~��5��<w��_R��R[��kޔ�]r@M�������66$�������b�	ZdN����~�������t�j; ."-���ҭ�IH]:����L���t5���+ ���o
�Q�Vn�
n�� ��n+.=~�U�� ���qk��_�iK�e]v�B�����-	n�����b~�8rˋ�����;�l&Q��/0�`3+*�����n�0�^a= q�$�z�H�[��}���R��<2+�C�{辣���&�!�e7�q�n���S��k��>(_�]��?�=���Ք�y��9��
S�sA��Q4J�c�Q����r��Dg2���ؖ��zU����`�f�}��qp�D2'vօ[����]��v��7E�G��ߐ��p���8�a���i�@�Yi�NM���a���30���>�*׽�G�\�!��b��rZxA�쫠J�++���ν��b��$�2
�����gwV4�yvH�]>���F���-+�s4����C������(J3�j��IT���F,�`�*#�Zg�����8F7+�mkg�v��Ti�>��yE��'O��q
�Ạ:^�����Y�!89���s7a�S9��cSޡ�c6����:ˠe"}�91.i߫���������/�T���Nb�K�Z)&=�<[xJ��d�Y}��E�>�H�}��Aa���0�,L{�X����JI��6*6N�5�YL�0%���rͥ�d8+S_���}��!�(l��?Ʒ�p�	�,��x�<��X8���ef�eo3���s���N}�w��	W�G��Y�t�)�iȇd��NB�>��xv.��5��L@*��U��"CLܷQӫѬD�@k�lJ�|=vi�cf�݋R��pǗ��N�,/�h���x�vė�+��q�$6=������?�_�%���dr�#��:<·���J�T+� =l��_9��>���t��6�@�Ѱ�oP�g����U��;�7O|�������R�)A����W��>3	�7��*�����Kޣ��G>G<���
���s��ocT�m��zX��Q%C�,��0@��^J�Hk���h��������ST�j��x��)�>>Յ��i���E�"4^���߁��NS�KR��q����Q�`:^?��+d��N#���(M�Q� JHc�^n�_;K�u�P/bD�P��X
�+g�ҷ�^x͟�`��b@.������I�60�^,܇��dV<@N���ϾhI�V�_�S�!>]�͛��o��HG���������<4�;@��3���W|zN�e��e�9nNz��.X~�A+����7�#��23i�h�0�8%rZ�.�?����Eb�JT_���;��ɱ�(���d�5��4��evG���9e#n�u�����u�έm״6A?b���>Ğ��;�	M�[�OwL\[�Y�'�G���_�!~O
�j�n�LFk[D�����	m����LU��)�E�(`j"b
N}�.��v�Ef�_�/j;м�p?=���=��<�:dN�+i�=�!.�0)۵vݯ����bj�.��u@��ÚN�%�O�|�Y���V��G1UM��Z��~�#��R:f7�3u��jK��c�h�Y:o��B�굓nH}4uh��,v���x&��뇪�w��"q��Z]q�~�'�$X��%X��(���ʁV�R��Ĉ:?�hnq�e�M. VM����k��Hc�s���Z�F_�ΨyTšX��ս��tۊB�С��Ah� �W�3N�n�*N�o��vߟ�^�XGSV��|�s[�����������i&��e�[��$������(o7PҺ#�0�]�ifڸDjD��D�r�h{�E,��z�x���}l��T6�η�9;�=U0{������5�&�:jNG��q;�5���秖�۵n�^�� ���X�i�X"�����z�.1�YFC�)�g��|���$���X��^�;@��#��l��|��D0�)���0�
�ԩ�<�m>�JU1��;Dw�J.[ �9����p��.D(Oy~��kR��O�(F����L)����=��?�6�������&5�����|ڛ�ImN��Q�YP�u\���g���њV���aא�� ��!��{1��!A�_�C�jY3f��lW���,=>��F�gFJa|�jч������]ٷ]���x�7�*�L��I��%�S������ ��A�o5Q��.��n��(eѽ�����L�T�'J�<._��M���mJ&f�m�!����G�:Q o�K�Q1G�<}i&ą��ŀ���ĲY|��qpW��7�v�o�)��c'r3$kc�]��a�ԉ��j���v�! ���i���r�)�۫GJ3��(Q�Ҳb��I�� �>͔�2�n�5SQ�IGw�pO%ց�$Ut��[]N��3L ���s��	\n���x ��z۳c�yE���⦛�,�$�*lJ������Ket*O���՗C&\���(�?24'教�o�yÝ4�"]�X)F28�"wۚ�P�28�_��3[@�$�i�萝M�;�bxG��$&Q��}S�&E֡چ��L��ۥ�*W�)T`��$�;��zh�2,Qe�pÈf�fܭ�#y�_V��T�+;ė�v{���gN��?k~j��)ވ�1++�^"�\u�s4ҥ%`�z�2^Z�	ڤ�-��vn���A���&9aW_ɾ7��)�����e6�� ʯgb��G�ܤ�5��n���[�����YP'}��.��II�[���[�m+���<�C4o��!�m�zC�{9����c<|�:��kǪi 겴�C���[#a�Z�M=�"�>F�·���atɑ5���1������̣���%������*��M���e'���E"*;����3�濄;=�E�mx�G{SF��ϭ�����X��QJΤݕ�J�e��D�T�x�[�XV�1m[�	�*.����s1�7�롺�V�D�<%47�po��r��ع��{G�oT0�
��k���x�^���],��&���|����V?�MC��
��dd*NOT�D뾩��{���T��<}�LF�Cw���4�t�77���;�"so��ߊiI��
I�њp}V��e�Fr��XCO\�$�n�ur��������.���r�¯Վ�ٰs���$�t\%�x��{y�G'X:Qҿzq��)�W��x4�)X38��d����0���y%P����뗛�,po��{-��-����A�T^�;[rs�L�-�ޒ��廉"�pXx~�O	]�� �e�AW-3� џJ��@x^��>x�6����l�<2{Q���r����R��_��)�c���������cr��V$#t0���P|�3���=-J���r��]�HhN^і`F}I��~ju��񴴽[�gO
��&-s��l5z޽��knd��v?���<�8�w�,���b��d4)`iT�u���K�k��'�r�NZ��+`��i!M(�9D�ݠzY��jD�GC5j����n�\���[Ε���Σj���D��o�ߒ��oU+�x��\���0��2�l>�w�Ftv���0�S���*���Ro��q��x��˾S���!o�H���C�R�JG̦��O�%i��X��W�R$v�>��YI����7x`���{zRPc{�D�Cɼ$n���$�i�
\[�Z�A�����g
�@�ӕ�T�#�*���.���D���T���M���҇�)�w
��0����,�Y�=}�~�^l�`�qہ7^��깠<��I�����g�=�?ø��܎,�-��r���w��w#'���p�Xt�12T+��_��<Q�dR��xD��9}BD
�h����j/;*Ao���C�k0����}Q*BS�WI?���M�����&m
�ʻ�Q�0n�\j̿Go�*�C&��/�y:�A"j�ٮO�{d�8�Ŭ#�����$�vF3��w2�}/Wk�_�ol�[C�C2�+��k+�]$�@�FJ��
L�Y�����9p��K@�~��L��-�Ry8Fz>H�D<ȭ�46��7 ��׼�M����x���Y_��q�Oo�1˞��t0*?2��N�JE|��䣊 >b xW��5+�\��
GZ���(m���jިˏ	
Y6�O�$�cj�:<�NP%�29Y��->�<�����(��fg�.H��p�
�uR�jd�Uv��\*����n�t�����O�n#�����$��gJ�|��6�x�}$&~�ɳ�vI�U�kCS)t)�fKѿ0�L=�S�֍�z�H�;������$d�������>,���*n������Hb��ϯ$�]��r�?F�$&�SK�b _i��Ե 
�%�*.V.:� �@�A6�eO��0A".\s5��h��9W��S1�F�Q+$l�+�E�`n@c8�}�W���7�(�]{�o�(����X�T�p���^���AMA���6o�x� TV��L����D*:�o�?4HX"iQ�O����;S�붧�JG���i吡Um�xO'�m�Z7d(a���n��(p��̜�Ǻ](��e%�u.�TD�����y,����M����{rf�����@�iiCܐ�j&�ׅZ��3g�~�i���3�y� z���jq�^���@��U�U	���x:Aöh������+�"v)��O2Y�/�!׀�l�ߝW�ښ�El�˥87ʊ4�G�<��GE�ݾ"|;��+��Y�?-E
����X�O8#�9y�$��e'�-z�l"�ŤxC���fx���r� "���6>���}�=:��}�h�9;��+&����X��H���@���#�c(��AHy�}�B�T
Xԇ������S~g�;�N
����S��*��ѩ��c�@�`it����uر�)Ȅ��`&a���K��yv2/�[)��`��/Q���} N�\�u���9�8�ň[�E�]Kb���~|����^����E��,k�/���8h�,�w)��a^�
�}��_㞮��RMb簵>-(��ZG6y�����^qY������	t�'>�l��&���P9�R.U���0�x'��Q��aW�?^9�g&2*9��T6��fDL�~>�]�'kf���GB�(�S����dW����xőС�+��m�2�##7"���u������u����S���L�"���9�q�N��"�#<��]��L)��V?�l�-�r;����P?5ǭ
/�C�l���r����ζ�i��U��	)y�:D��i�6ݚ|�m[�C̯l�A�Y�fcf0=�|zzZ�J�߇�?��V
�U�u9e&Ԇ� 3O������E��)a�.l�X`�����Hy� ��U,Xs�O���Y���t"�e뇪ݝ�z�~O.Z�:���=A������L�u�����b�\l�u=���� ���tS27$�'�B �52�2��!��m�$�֠b���i-�)S��w}�ɤ��� ��R��P�8��޶�X��U�AX��kF��ɻTf~�V��u�a<��	K�������T�ݧ �r%�)@�����怯S㹧����S�U[�B>T׀3xW:x���xn)4#����+z�Ǟ��������(��(��0.3`��/�ֻ�

	&��hu������|ԭ�e�a;`3�T��P��c�ef� ��q��Z�8!���,l��F�����<,��Y�D�H��^�����KV�U��%���-*���W�WHP��V��*�L=|��7.Y�ߵ�9�b<<>�䄓�0/צ�CFv�:�J��T.&�%܌�&J7���51-�e�""~ˀ�:��%bX�>�L�/͓�uʅ�9���w��B�*�����!�\dA|,f#}������)�8�="]�}z�YZ��~��c�i"T��%AfUYIn��e��n���Ĳr�^�a>�V�<�$\L6~On4d� P~!��!���*Gu�)bPP�<�ޢy�B�T������M5I�L�T׻�8�A�f����lA��+��Jn
'r4��ڹ��,M6-	�IF~Y��
#��]��ꛭ
_:侐ؤK�9�M�����"���1m4v��!�u5!�~"T-�n��7�H:O�O`�ZD�)���P�aX�L��h����O��uV)]���,�j�� G�\�^x�i�T�!"�LBt|(��9 qe��;?�Ѧ���85����PW��>"�H����l)����^�1m��g�g/�s?J���?@1�J���)��J��o9.~��BYU��گ�gj��P6��`x��e�lKU����6U���
��f��`��t����1�T������
 �5�_���]�G0���+����+� =0�/�)���7I��s �O��j,����Ul��{��n�1��j��ِĴ����(�e�=�_f����� ��t'�J+8`��}��������ƴ3�]�B��2^�W�ooϼ�l�m�=vLóP��\Ұ�&w���J���	�LA����; j�璷�v9�*Mw�r�gڑN�6�UA����Γ���е=ň�P�ki�UQ��bjr��o�Н&I�Ŀ����=ss̩�X���]t�pU���bWV�D��0��Tc�kSI�߳��J�].~�W�����Q"+n,�TWϦP�o'^h��yU�}7"��+��r�O�K,�-����cꚙC��_/����9���N� �$��4��tNv��ҭ�]��j��Q�\��Oo!�E#��I51�H��K���g�c��A��e�َ�˻5�sh��������}�Z�k1�c����DR�������O׬
���Y:��H^ډ�\�n���#������kGy��[�L�;�V��}�W��'���^?�F�ܔЌ7�,�QH��Z-w޸j#�W@?ʺ�ٽ��]�K�&�w�� ӈD��U��<H�SID�&�ü��*��.8����[�ÿ��9a^��ȫ/z�&�&���ػ_VK|�?�~~��B�E/8���O����˭t_i���{���"�j#�7!��]l���h����<:+6�5��'�0I��w�wG�G����l����F��� �Q�6��X,Y\�0�\A���`�"� 
�o���� 㳦mP����lI�y�{�<D|T��L�p�z�KA�=�A���
��֢[V����������=�Au[]:KU��>7<Q�����j�0�/�^�y�ek�ztr���Ԯ��Tn������Cb��Q����;�E,}R�	ɾ�z�����#-㿷Z5��k�9KD�,�F�_s�P���(u~|\;�} �RO������wS����`n�$<`s!��(O8e�;�$+'R��	�H�7��d^�2�$��f ʳ>���&�傪��\"��z%�a����
������p$i���m��b���X�@"?�����=ś�lu����F�M5R�k<Z^F3��Q*�l��3_���T�Z���!�*�m{/w*���Ae���_6���F�[��EVfq��Q��A����^A
tl�)I�����a��<��!�\G�\np����̙`��z�?���U�m�6q�4	"������*h%��v��"������,���b��f��׏�A�+q*���(���x���kL7d�NYX�LM���r#&vM���6'�HD�G 	_�;.岾[\۰�����X��$6/$�KD}+��~�M�C`�;E��$��G�+/����R�R ?�!��['+u&�_�d.Ň�9C�2RAց�'E�y1.��o��~�[7�˭A��	��2��{$�~�E������.Vw�B�v�y��Ők6��pMۦ�;mL�Y�S��b&�Y���g��������:�A�re��~�?+G!8�37S�kR����R�,b|�D�+qeKa�[����K���#�?d��T#�D�zy����\�!a-��������¶���?��թPxJ�z�Mئ���=eI�p��Y�v�,�@����H�\j�77�@�:P���i��yI�����Y���J�X	���9q��mJc��r�G�	�����&T]��p�҃���<�[A�nSs6��U<��2W8��|�@E�u�T���,��)(Z-��"z8;o�y�1����q�6ȷhJL�d��ML�&�A.������Җ#l�y֍= X���꽧�ޚS\q��{�_>0�S��銟&2�(8	4h;'��O����f��`��4�⸱_�*%��ֻ�E^PqbJ$����Ţ���Q	�,��-,vB3�7�(�p�	�l.�d�<�-�R/�Y���fM)	@��3O7�G�^�/2�;���_ӥ{����a�F�k��I�u�<�@fcÖ�����+�[1�l�ޕ(p!+��p��K��M�-X2��J�jr�>������ք�ո|L��3�h��\��E<e׺������܉�	�J��� �Q�+)ԍq
f4_]�@�w����i�Q<82üY]=ʨ:+�b��e�� �����,t;谉Mo��	��af*�LV ��Ow<��{�0=p�"�ƹ\<�_����6�3Q�
��'?���v`��~h�4!���iKNY�!��)�'�13v��)��)��7�8Z���yM�������%�c[ւăplTQ8�*��,�-"��.��lۇ�����{f��C�����k�@�JT����j���}�HQ��G��.zYc�����C����8�$�Vݬ����nzY�s�9�����Q��:�Ԣ2���#)H�����1PIR��^���X�1b;��+B"_0�S�L�	��j��~�hSE�宽Z��CXv��H���o,�	�����T�}w�>Z�^�ʙ��-8����6��`�bv�~�E2�����Q+�9��L�g��K��z�`sK���6>�uF��4]����]R�څW_7*2A��5���_��Д߶z��ב��~	�*I%� )��F�����!Ds�p`���S/OM�/�M��m�t����q����	��>0�v;��W{1y�b]6�/�r�������9�_��/�I]�΃W�J<�,��N����oMb��ۦ��1���kϰ��p�];:���Α;9��4������d��#�	��C�)�]�q��3�rt�����ފh@�0$j-�'��+�fF�wW�'�����24aR�	����2��'+�G&���;xd(�zE��r�ؓ\8�+�]��Y�t���,4����1_Կ7׺<��Z[Nu��	�ѥ�]5֜2	os�8ԝ�k�x���9���-����l��|�ňIa��`�D͹����9[uE= ³w�Oy�����h)��n�x��f���UfJM�5tK������eU*�~`�2�^ji����3�
p�����OqI Ū���'� \��]�0rFn�TGB��<զ��pBl3G�T�:�yl�C;3]jQ�Pc;�_@F�O��B��uUvS�D��:Uƞ���CN��W���o��ʉ?<~$1��Ywy�~���Iqa��;���o��eW��5v��M��tж>��=~9PC
ܶK�����A=���c�가R�}�.�,{>u�v&�����4d-�y���e�c\;_�z�m�	Y�C{�~hEt�S��ס4A�*8`�@�ڍ����?�����5� 1/F%⫎Și�-ԫa*
)��,2Ύ�ï�,c�ć#���=y7(�[�Cj�`��BUb<�+��9� �g�K�D�jlrBE�7+���.Qq���=�r���.��'F��hJ��n�x����g����v(�TV��M�6C��CĞ�t1
ve��H�ʫ���Q�X�'�x���b�4NJ�|�I�e�\�)��3�Q�y�\�(L��8��:ȝ-�h�����4Ƕ(L��1(��E:���A���PNlR���#�NG5�R�]�:.V��^��2�!����J.A#��)܍�1OeU<����>���A�^�)&;��x�`G&�y;ԶLs�9�C�{H��I���O�OyQ��;ҳ,͆8�F`D��h�D��7���Q񥍔`o�;�NeEaj=����Ю�i@��d'�4!���M>E��]^v��!���~��П�Ȧi����x{%#\�#��oMGT:m�lv��rq1�*��ߓ������2o���Id�{¢�^@�m/�#��[��=?�e��d,_+/I�j�m���3èI8���9\-�q��nd�a�L�Q�����_>�T^yL!��H�l�W�ͪܕ�y�?𞪌�"���ӗ22�R��0��u��(z�Ӥ�2�K{�_$��V`,۪�&E�]2.���Q��S����ҝa�^�y��wD�)!y��ƿ��p[6k����w��$'	�_�̪}<�T`,�튁�%��_��ZXѷ%\j��*_��钹l�s{�p#�^:�fH��:��"����ᓡ�68��5F�v����q�ke�`�����3�`�:��P��%1��XyO�1a�k*���|���Z�#vƄ���<B��	=��P�ܴ"�ft���h3H���G��7�Ө��xr��+tA��^@1�C@adg.&6wT+h�8�����o�#y��0��zK��&K���v��݅
�ɚ�V �C��Pل`b�KK&�ճUQ�&�2��8�):�����6T����
w�U���m�ܳ���[�$��I�%��&�l�Vp
�x�5�ǫ���(���8Q�2�cp'G�Ua����9�D�E'�4-8��1?�0D5t�QYbl�������P��`�|̐�7#�Fs=1
��-ݫ�O� >c�#�=��~Y#�yg�r��:���T��R���?�P�����"�1I�e�}j/A��up$������T�P�������[��j��¼��Ӟp�R��bT������ݿ���Y�g��:oc7�3�Bל��^ 7�V+��忐��B���6��ovC���9����GT����I�`���x��f�`��^�~���!�w���$6xc5���(����]	�3;ix�Q_i��e�J�4�������6�@:�Oi��ɳ@r����+*cV��C�$U&�A��1L���=N�5/�ڸ�"%��9��D{4�gZ��F��]�]h�Bt������JX���r%�<vW>���
F��W���w�F�1}~�o)	������}��/��� ؑy­��aBN�� {��T=iO�3�Bz��j����R��ei�7��F��ؑ7��@�����/����Ӟ�W���$�kX,��9�BM��\�#�kf��Х��h�����PjＸ+-���r����^����n��S�"p��i���r���y~�ݮ�0\A0��ȃ�"�1l�b��n�3I5��&gt���1>P:+���Ԅ��Z��.�ai�Lsu��\����rK�+���wa��R:�d��ޯ�D/�d��
�LM�m�c:P��<���=
�k�NЬ��C3W
G/���Gj�@Ă��@ׯ	��=���HE��r����������fϘ=�y]����W�eI�b�����1�:����2Wkܿ��0+2]&e9��?�ttA�e���!�)bA�5�癄)\�w��A[����m����4���Zp�;��M���d�oq���·SHJ}��s��nv����!}eIe����A��
��w��z}U|�V&B��-"���C��]��ϩ^�{�-��t�&�]����7�q%�w�U�܄�0P��Ts���7� vqF�X+���d�� qC�#�pG�\����X���2b'�G
W���FX�~��^�/�c�pn 1h��	kb��}�����R}��ɖd�5�f�xBu�8�&jwQ���c�>n�U�փp	�����.��a]�Ū����e�eQ���gFRO��aE>{{� ��\Urzc+Č���a&���ٕ��o���7���}�����wg�-5�#�T>R(:r,�iӄ��3��1cR��ƶ	G������ j�+z��$s�h`��g�r�=�2}u�����O��g�C΂Ej��ѳZ�i���F�2�BO��/.��ɢAW|/�F^xR�'��7y����vb����q�`�_n[i~��4�� �[�,����E�����4�� ��1!L��T
�sm �X�a ���WD�o]���V�
3��{��!����='���G���`���T������5�]�_sj[�U�F8/��ғ�b;��8�']4�����A�I��quO~��z����=�Y��C��2�nJ4<�����x�m0rT]�5-���e�Yy<�L��)�ӻ��8�P����U7Y���S�a�&݃S���9Fa��*U:u��8��;}�SF�
k/�Yߢ�k�1�g?�Q�Q�ΉŻ{��>�r%��C0��Ğ#ܚ���2]/��li?LP<MakrJt��FD�Y�f�HL�_Uɇd���2�i�Ѯ�^�����+B��R6�ZC�7������(���qF��1�֥l�)]$�s���X�l��6�]�w�@����A��L��h��R~��~O1�,���r�%>knя�;���<�O�됪�y���Hj�C�������#� �/wU��w��@l8N	w7�s�)���΃ݭw�}�3�a�@��x١��}c�1ߗDW+ڃ���תm�
�
z�ǑA�V�ƫ��@�!������W�%�t,��1i����T���Bgh�D��^� ��� J���٤	������t���=�T*��N�[|��u���2�9(��Y8Rn������Wݕp*��m����N2�֢J,]ZK�g�LLb�$;#kT�N�*��۵�n}'N<������z�mT��4=�L�$篹���`�`���a4l��.ȥ�;�c�A>i�	XX�~���uf�C���q�2�/L��=�����(����#��ʫ���z�6��'��َ��C��3��7찹��Ga��MV��\$���j$G�d` ��0$�Etє+q��o�h-�x\i$t�p�i�����'���� ���yt!��P]7}	F��;_o��U�v��7S	��*�V�Λ5��t�uD��EՒ��D���w�b�T����b���A���9��܈�}�t��u2z'C�7�0�Z0*��,��-���GG,s����G q�'+�V-�.��l�Rn���Ok�x?���A���s�=�\^8:�l��Qa2H
739�wm4��%н�� ��]CG�2��y�3��+�mR�'i�Z�� _��A� ��./�؂�{3`V٬��  ����<E�Э�Z����F�T�Q�D?���_Iju��3��M:(����Z1i�^��FF)V���p#c:�*�g�]�Lj�k��r����U��,ĦX�{���"��8�$
53j��`h�)���T���z����;�6u�P�3�v����7Ƙ,��~�u����H%�V~̎�l%���z��W�D+kx�>,w�?l�a�:�� �1]��Fn!�Ցv�p���_GG���V��c���J�����) i��D��9z�QW1�f����z�&� Mt��ck�w�����SE��΍�V�/��=*�� ��m\e���k~�4�d]����_C'v���������.�b7�P��*�o�)J$(��bX�]�܊��<BX�f4���Yϱ?�)GrjW�d�;Pik%v3+M�n�YY��I��#6מ�`P-� Makɻ`���h�X� G���34��{^?�rZ@S_����S-�ف�w�Dp�D�uF�]lw��˟Wn_�#<�����2$T���p��}� B��BGR �
�;-p�
 bk�^T�@	 �(��4��Fs'5�}��)�1
9Z_n�ަ�-�w��E�B��rۜ�Ѿ?+b$��ŧ��y��;�4O��b��`hQ��#�o��_�`�2�W�ٝv- �����qU�����n�<��zIPqKk�%�8�.N���(f���@���o�PW¸�(7=B;a����ї>���A@:�@M�p��e�a&J%�>g�:~��R��v�!sP�oܻ�#��D�wd�M�/#��֬�4��#u���9�����Ĉ:Il�U����������LZ�0*��5:��
h�C�[�"x�'ѓ F�:/e�U�||<�?�|�q�������}f>�ܷ�����̆�G ��h}w�t%%�Dy��7������v�%l$E0�TJl�(UaP���IH�.wj)�J��r(��N�QL;�L����2S*���� C�'�M��h��K8�x=q���4�W��=�F��c34Z��6�B�\&���ܝ�~z���%�/}��Fl�*W*"W�N���F��T�~�mbؐ��sG�2��s
�[�Q=�Qws3�g�E:��b�\/"�/��9�0�'�g#e<���뼢A�`�`T��y�غ�o�I#7�q��N�wbQ�*;l���
��Yo�b�E����8��^�þə��9��|��33mt���ާn�iX� ��Ϳڍ),Ϭ����C�Բ�B�"R6S��[�R�B-��x'�ᣥ�!�|�F��)�,x��	��<o7+A[w)�L]=i��qp����C��9���}kO�H�����K��]�W7����e�����Fև;����y�P��kQ/X}9���Њz�\3	�]G Y6��=�3��slR�Y���R�|9��톳���m�h[�h�Ԅ!V�X�d�i��=�ԫ��L�퇧!|��{$�������� G�6(�6u��;�C@��1h��|%��
����yI=�z������U�X	��x�!�[O�Z_ނ� ��/o �B��7}�����r�8�-@��}�)73i��g��?�3�[�4��}d�*�5/��BL��DL���jt؅,�ֲ�;��:$����V5'��u�D�p��Ւ�����6^r��^)���--y�:�p<��\`��������7I�'d� ̹�PY(��gk!�53`c����%�
��$��6G��50�%� kp�O[�0j��V�����Z�K7J�D��h4uG`�roV&�L���*<��M�>X��/�D�
���YK����2�+�J�.j�|���߿�qM�:�s��@�(̔�6�v�)�d��`�ј+�&��rrjo���1�����!��8�( 'I9�夥���Z������r�0�#a_,gr`�49�n������Ĳ��uk��9u�N��I}�-A\�<��/���}c&@7�7�e������Ɯͽti:�T�`/���u���g����/4�����r�E*T�Z�����Fφ��(��B�)�{�5{����R��a;,�ג�+��j��i�J�0���'c"Ryc8�E~W�E*K�Z�y�q��LF櫻 �4�ֵz;O�[.L�j�-qmĽS	�M*!�+
K������N��?׫�̓�Hi�G��,��xj2@�)���݈��t	�B��MR��HAQ���/
�[&د4�҃U��;{2s�����"J����j0?�_�;�x�q�(?"ӽ"�ߋ硎M�I���mP��G�z#6H�9T?�\#�1�*�J!�*8� �!C�XE�
F���j�]����+L�?,E~A; 2��Zl��ܽ,����\s���Iv�����4���%fr쫶��������+E/AU](���N���r��ƚ�L]qv��Їu��ĈF�o�׻s�q�@)gj��5�|�� >�y��֏��tÿ����@K�g��(�`]����!�Ũpþ
��������ū'W�����B�3nK-h��;����'�&���u���p@�G����TJ��K\����%��|����Z2�)�de��8{�(�h�As��9&8�d�}}��hb�GG��X�%�&0��c��k('!c��������ո�˔&��$y��%]�2��U���J(sX��?qZN���Kd��	��9vx�+hw�O��NA8�ƶ��1R�Z��:R=i��xJ\�����s������o��z3�jd��2�b�_�B�P0+��MR�D-@c�aɿ,��������:�JZV�G{
�����:|n@�J,�y2��$4m?O8x�X����/!&�:_�8���H�5
�C����������Nۘ4'D}e(r���FQt�&��Uc���!C�Rm�9ePn� ��F�ηB�' �w�gW���5ĉ���\m��^�ݐ���������تy���_�p�w1�����,p�7s%xB6��=ǭ����[�1�ǛW�9�|E�ü��G�>��0,`��	D��DAt/h�7��fl<�?'}�,�ȣ�5�;��7�A���o�t�(Da���?pM�5���i8�2���K]���pFvxF[S)������UI�H��[�;�vT��tv~U����lɅ���>���;�UBA��Y���<�ސ^s�''�8	��뵡"2�F�)OW������+�^�XT�`�����pѠ�B2+�1�i��g�/SXDL�D�*?������a���3��xrݟaf�։�Zܗ���(v}ذ��r��l�d��lR�D�[<{�z�!�I~ӭ���8q�DhF�zQ{��H M|�o`榸�_�D<Hg�w�KJ�c�]W�k�c�/<�ͪ8������-��cRJ`�H;{�?�'>P+�쎠�`�ǿ�&~V�+�@�R�b�k��4s��/��s=B��I��Y��T����`B�]�s���1�I<@`� �n\+Cd)<�|׷؞>��M�zo��u�`WiI*;7t|;C+�@eL�9V�D:s�bh>	EST��cC��:[�&<��8H�5�K*��˦W\�:�S�B�����!~��e;қ̋�[
�h*ȇ?�#v,PH��ل�x�]m��>��c�]�����yF�g�#�4l�EW�'��W�k~�w��sad�������mM�!��_�-|����E�p��gH��J^��iQ�9�.���ɀ�`�Q�{��A���F@�З��7�0����}�pHN��ѡ��-c¯~�`�Ơ`"FX��N��]B#�u��b����Ui��?�B��n�WXR�pO������/�6~��5,��õ7R'[X̕�-àB��_��^�G�V���8��$�ݱsL�k/{m�@���v+.��k���%xQ��N(���O��KH�� a5ZZ��Q���g�����:;.M�-�9��k/���#Y���oʥ%�0|W'p[k�u^�X��9�^�"��F! 3_�z��OOr�#�#�j�r�S�X��$#�hJӠ̼<�p~[����&���E�R�9�SE�T��	D�����M\���w��5�L)�5��F�.��d�0��1��e�+ ��S����+�9^�- �5��w���m�X}�u*H�O��1��kI�ubY\Ͽ(q?�n���I�{�������J�	^~��WZ��������겞S�:*f��εI�-��io
"ua���*��C��:�K�������3ޙ-���`�r�h�:=�%/z�7�?�������,�m�x����,'H���q0�#�}���=|(����s����ZIͨG��������x�r�c?�5��������sеlaW�yf��J��>�� l�lv�h��]+3�3έ(���)�wئ�����я4C��*	�I������ёd��W�_dTrξzP��N�S�_����
����9J���*�ל�A���Q� ۶|	J�B���Bo�����8���x�mngr�W{�X�9l�uޞ������� i0|�밟��(� E��`'�����#�zf���xg���W,�k���)t��A�h��e�מʊ��;���ȵ�bcٽ��s��߽LF���c0:Ǘ�ӹM�IΘ��_--0zæ�'k}E�# �vJ���LL3����6x�v�$I���#)������Q���؝�-hUD��-;ο�[�A���>�$�s�g"N��fލ�]�Zn�ih�`^l�� 	�Ģ���'Y��ڗl����b���ݿ��<�F�BŐ����Q���?�R?}��d�}�&4{���A��4G��N��pU���l�]%���!�`nlrn���ۅ`�@~�2��1���%���'���t�&v�#w�U��!^.����t�,E�~Z�
���Q�qn����ꦒy\:���lI��`QڤX�"р�2sO�*>%�����(��9Ĳu�t~f��u����b�VE�i�Q)���@�iӣ�oĤ�����ʔf�dW�a����<�͂�?�CE��X��]�-I����A���qc�͍��ku��1SY��
Q�O2�Z��������>���J�#}A��'�tU&r�)��&(\9�/>��5뚰	Zv�Ҧ��c8~h�0WO���٢"eCY	IN����W��b�j�D=/ϟ.�EJ��9�%�Z�W�p�N.q��D`�Z��t�S�g�g����x������`Mss����.�j���='y��N��u�aw_�����ۮ�ع���v|�5_ـ	xϦ���v*'�N�,E3�ݞ��,FG��~�n�|��=ye�b�8���K9�>�|8B�����5/	� /�M̘ eƠ?X�JQ��~3�9��z��8{����5��?�͝�'h�����iv|���R�N�l�2ѿ��o&?U�*;�}��;�b��Ǳ)��0���}�"Y��^X��S"4+�ʓ�p�.[ݩ$���Jo��W �����[�Qޱ�"hg	�R�&[+1s��0�9�n�C�6ݗ'h{�ZW|-i:�
�4d�� �؆,�8���[��H�t)/�-)>rn﹇�J1-sm�'/$R���P�w	H�}:aX��,���u���J��(@v"4��+*u]�.2q���`�I������#V(^�
4aJ"���N#d��Xظ���������
NE��dmc	��P�>i�~�'}#��t9��c1���ƪ�^ k?H ¿��n_u�u&�}Z�M��xs9�Rj�;�b#T�)Zx|w(J��C��I��ͻ��T)��ǔ�gW��$�&P{�5(O��Ek��PY��/iֽ��,ҡ�O,���̀��zH�;<G)��1�U,(4�#��1�<z�к�7#�x���QG*����s�nf	jo�U� �vƅt�J�ƹ�T���=��A��"��5�_��.��~�E����^���E�s��Я3+Z<\���ku�N:�3G���I�1�5����r�\���1�!K�$���u�_�	}�q�޸_\�I�����4�i�'aX�xtm����4��?�t%��l֙K�6������n�Cz�W�v�#��1,�Bۏ����ο��if��GLFo&�������$��1fF�u|!�69��"@�)</x�VJ�!�'�v�LW�7X��D����P��gi���Zx��󇝡���)�����[ˈ��Wa��]h��Ѕ�3uo�kI4�F~r�����4�FD\�Cv+\r;MI�;�i;y%6�H��/��{	 �y�Y����2o#�q��m@��T!
�f��e�H�������4� ES�ъ^��2��vw�U�3Z�X����(7֧p��ZB�������7ON�_W(:��:�&�05�,��!��)��]�q�b���tF9���ɻ����������q����}e+M[�^(�m�1����\�ް�)�iA{2[>.]ܟ&��B	x�1�Yv���Z�b��m��黇<��ޚ�o�i7n�W��/�'	�]���"�6-Ǹ���B6��4ZL-k�Ϧ�Y
�$�(Z�Y���(*h��ww(^#�4`H�	��|ڷ�2���� ���?YY�����Ò���Ԫ�c�M��D�,�:-�H]:�\]�&��<
�-T��Q�KbHe�K�lp�ޒ���AZ`�1��rk�л��D���.��Dm�z�He=���|4@�c�L����А^�ɇ�]8�'���+x��	\j�[������=��b~C&�(kxO��ˮa+q�����4�712�:��9��>a.7W�D������H��s����D��W&rD���Z�L�#�E��L@�k�e�B�\��l�fC�Z�T�����k���
�)/.xZ�iFK�}0�=�@;���UX���!3A�D�e��/�'�&�K�t���:��0v��w��7k	0�	�h1,^5��.�!��� lA;��NH�j����`�J�g͒Q�`Y~��"*%F� ��F�/ѕ�Q5�2�!�di��dS�߷)�'^VF���j��Z�����E&@̷(0�}&��V}he^��n�п��G�(����,yB���GǗrBK�������Z��q��ʦ�%�����t6�W��z�st���r��+E���5�[��Ȣ�/�9$�7�<�X4Oc�)Rą�l��d�F�}�C�wnn�S�--(Ѝ��6~�x���>�\�����C�U=2����0A/H��`�����1��aRژ�憑i��E��+���e{-����G{��4d���~�̢E6��"��X`#1�5к����;�M'���|�40g�4ѡ���(�Y@�,�hG��z�/��l'	 6
n���B���z,w�~���()�Z��Jd!��&s�B�`��h�	�ϊu}�}�=�j�������͒o���� >?s��Y���3��kW���M�x5REO�ú�Qx-�]�z�b�C��5V�D��D�\Y�8|ŏ�jz��1 ~�n@bu�w�h��ej�1x�P�l���R�t2B��>�cڦ/?]��:��j��.`L���8CC>/<,`�I�p6��
��>���W�.:,�����&�65�d_)+�(�S��Y1K�g�0
�v���f�dS�1ݭǛk����3.��:����ֈ������o!"���V��c\�ӷ��+D��3Ѽ	��q����+�J{-���~��r����B�q"N�]��V�IC/�T.㺞8?�Y#�Jȫ�Y�(��T �E�M!���B�~\��'�w��]�A��Z+� 
;hi�~��3d�m �3�8
A��-��4�h������'��B(����f��Nŉ�&�h�џ���)�G*�����A���BA���T���y���E1A�u��.�IW�
����/	z�d�K�����m�uq���a]bpc�� 2��h��a
q��zΘ�����%�����O��4�j2�A,rڹ�:@� ��%k&�i�N<ruԴ���4���pU�V�:����&�����Yٕ�������~�tv^�=�m$�_��%/* �]���<|��FC�1�i�W�7w9��gʸ-�wz6�X�/]͒Y��4�ћ��{��@a�~Jp,�����F�\.������3ؤm��Mm2�)�k�$&V!��]��$�?�t�c6�<�;}5b���7���~����8���B:����鲊��&A�������rK�)o<�f�����N�8F"A���""��ˤ�@|0��N
��3bGF��%m��F\ߍ,9q�����hIo�Ρ9+F<�@8
��#�\%��L���%��CVON����wZ�dv��)��T�aHA^�䋒�k����1C1�Ԥ�3{�<��3�A"�^�ҵ�?Z�eM��3jz�8ro�i(wo�bz�5
J����8s��V	C��^��h�Ǳe:pw�Azn"���a���'��yV
�Ħ#�N�/τ��ӽ�	���T
e ڻqL�dfw�eڅ�gyws/�&�#_L�'L<���ô�(7)����|��<�uǻ�k� 4f�(6�=����$ �2���'�z轇*2��0��	W=�x�p�5̜����
�VB��k��&@�G�k�	��ro܄���V;�V��Ņv4At=�[��wa���@�N�&�<=�~{�w9���>���AS^<
DXl��f�������;�,+�M��)x�ӥ�O����J�#�;��Ԍ�T�JMT�N��lP�f_m�v���_�`�Т�T'n���5������k�#���u(�
���1��@:��,��l���"zL�p O)���� ���g�ys�A`�Z�����1&�f����g����K����R�[
���cO;)� ?��7�s=�4�\
~��d�[�%К��4SwES{PƯ���8��s{��;䂚p�Mܢ8�"��Q`V���UI}��7;U[V	/y��1��onEs���EmI���M�ND�{�*�xu�W�;���p?�	TI�)��+��i��mƼ�n8����MUy-(!.���BMլ�W�b�c���ג 1�,}���K����%�-�t�	b@��y
�T+��w� �y��b"z�M�F�I�x������N�]?�E���hT�Se\�eQ��\�尦��5*���okT��"~�]�=g99�����?��G��,��Q��e]��Xr���T�/�������bB�(R�1�1��:럐�X�����9�.'�4��>3{����(X@�t��{p�~��Cn�^��\*�R�#?@CC�+��,���i#,"�}m@���`�r���G���%?��G�/�� p0DEx���)I�(dF�Խ6F�a�u�}ɏr$�)�O���&�������N�]���E<iG�T�v�n�譑
Zٻ��"I�K��8�3��N�,]�
��D���]k<���U򱆒1gT� ���+�i� �M�1'��%��ަ�琦���91�m��%���F���fLa'�4{�K���ڌ��'�}/OHN����?����`�0��f?Up�MQkm���d�k�
77����y�!GS
�랿ȴ��K�rMF�G�O�c�� u4��h�A�d�P��^B�?��'��Uz�e�SDi�<��A;���` �c����A�ۓ�^7<�i���y��,ܓ�Q�]y�/�]���a�-�S�h=r��~H��/_���%�j@���&��fo��O=��(� �vzY~�"�V�
�I��rZji)�_�߬6�R'/�q��X��p�.�=D�m�|%���m4Ge����M���&� 
��\w4�*
���RF85G�^�,�l�NI�%�\{��}���,��D枟,v�xTچ>�&�~��w#�{(�������j��É�I ��l7}��c�5k��7����{�x<V�!Sh�Z�n
�iL�q����x4W��-z�(��Yࢷ<��S���8"�\�hscX���u0O	��n�6 |��
|o���b�.'^�S�$�o�_�ɩZ��Ly1��DB�B,��@r�CDz��Unt����%S������J������x�PNN��#�Y	�j����N����#�L�,��=��y�\��P;1�����ӈ���!������1�! ]�|f^o��>��ѫ���߂�ͣ�l}�k���Ͱͣ���X�i�4I�Nxs���5u�%8m�`O�b�Mkl�Ǡ�����_X#�<���n"��d]����<�P&��t��>�aT�?�qO,��Y��k�9R�������CI��t��{��:u���$,
��>	���Q��q�5}�gh�Y��o	$�S�C������ip�֗����˧������O�T�b�vBq4?e;�N�n#�H��/B����=���=An��9 um���<v��!L��|~N��t����Q9�q���(jr�#�E�@��a&��ĵ�=ƕg�:3� ���%��dYh��o�ftLJ���m_��%�O5�@: 5���f]��;��}�Cx��( N%ö� ����
�?i�L5Zr/��s�N�k霔v������p��&�c&� �?���l�U�@#�Bo
s^ש*�#�
m��*!�r�oz�3��A"���0��د�`�ԙ��u�rS27�A�Y��µ�z��CQ+( ����8�b�	̹��,/��
7r��l=�̚ S9�Q��\���lED�Y���ϣS�����I+|J�"y�j�it�))�1����?Zp]�� ��4�F���`����,q�f�
�!�-٪r��H����MkE��F[qɞ����0�11()'(��ĻvN��vwy�]�?�ȸ����I��;��~[@ Fi�� ��N<V��X�OC�ڲ��> h'��~����:-�Er�iQ�j"o��ÚK"\��Ykt������Ѣ�<j8qU`"؟!�1�7a�Z�Vu>85���5%ι���u�qP���x�ˈz��h|�-{��fK�G?�N��uR�c��-�T��{}����+�BJ�D���.S�C�T��T6+��r������i_���eV���x4-�T��y��˦*���%�#������ ���6�UG˯���K�G���B����9yP �%C�2���%��Z�����N*A��0Bҗ�CB@��8I�Z%Z��'.w;�c�1�UN���W-��(�7Uy�J;�B�3��#��(a�j��[/rK���%bj���9�P�T�'1h���4�X����ih���������RnAb�g�(ԉ
��Ͱ��s������0�KUI���L�CW]�g@����r�VrH�3���B�E�p�����e� �B�棢P�q�jKo3���tv��?�J��d�1��:@��������݇��G@,ݯ�w��S����ui�G�ު�<���kh�l-D@U��,��mu���9��ŕ4�g� F%���Y�e��p��ʼ>�A*��~a����|�ᕬMb[F)�U3��N8�3q��[;��H�>4��y�5z;���hW�����Kt�`�G�����x�9mh�Pl�Q8�͋a4���S�(Đ���e� ǿY������{)�"��&���� �͌asE����g�ť����x�|�It�� �:�/N������%)�br-���b��,W��ۭ\�cfTT����/������c�&��M۸�`�b̉f{������7i����gX�)8W����x���r
��ˎ]��k9�� �D�Q�02=n$�o�Y����[p�� c�zH��l �ͤ��������i�u;��"_��)�J�ϑ�6�ʰVs�m�A��)=�r�{�=��B�q`=��r9hh>��;��*�G9�|�۩���G!��}��Z��CA�¥H���R��>�5C pG�;+<U��
nDM���.K�g?��Q���27��p����O:���@$_*ߓ�8 ~��8��5W3`렊@������ du�*�~#�q�V*�����w�f��c���Z�!��g�FY��F�Q��Xj0�0B�]��xs=�x~Y�ͥpd r���g&�R�,���V���aa�O�b�<S�x?ITBƐ�|FOԆ�|؍�x��F�#�T�ʛ��H���hS�iob$��?�iݮ�$�Iҵ u���ߢ@�Q�o��{�,���N��0�J�Ma�q�G���Kc���n�v�i����S�$����(�O��HIk������<�\'/���a��wg�C�¡�g��Ze!k�%����9�s�	+C<l������]P����3MZ�>h�����UYb�	N���j���?��-�wt�X�}h��9i��~l�� VQm�N�7N��xўS��	1)�N89h�W��x	�P��ݎII駫V}!�vU�M�8B��ѽ�s֯�V���N�T~Ģ�-���g��X��;g
/��(�=N��D�u�(E��@=	��&�Å�}�0���kD.��3��i\\����(]6��x'�ے�D8!ĕp�3n�h��1� @y�Fޥy^P^N��K^Ð{dvM�ُS��b5�k-�`d#�ݪ+�.M,o܍���<�s��K��8fL�K�ܨM��<`^$C3��{w��1���x,���fH�,�L�3z��:@0�w�l1�X�V#���#��3\��0?L �ܵ�k��B�'��c��[��2@լ�o��ۗq�F�	�qP�L�w�̙-�7"x�fx��C�x�<�ɽ�k ��*5	���q��N��p�O��7�[Ơ�Z-��GKa��~1���6�RW^&Z�����N%���}^^�W��d��Ϩ6��Y
�6%BK����_�M(�#��S�=0&T?��'d��41��'�@��&F���Q(w��ņ�2������	(Ԛ�ڀ�,��Gh��/`��i�܌� TFl0-����~D�(tf[�<a}s�'r�/�~Ep��Igϴ?�m�t���+��s	�L��ɳ¡ o�x�اm;h3a34I�����(�;�c���sD<v�!���kG�$b��[?ώ���+�I��Kï3��k[�r�ٳ�cE��v��u�+n�D>^$�B8J��ƶ,Y���^3������t�������J"�E���:�?T�F�N!�y�J�ݝ���g���p�!��O�� ;���Sj����3�>�.���f�$�x��b�ş���	�
����%4C��\�I�oǍ���������z,��/�9e��,D�;XIr]�0v#v�&���2Dau9HEǁ=~S��l���� 6Е8T�\��#sc��%�c(D�w����6g��gCt�IwW8@)^U�.�_5�7�$�qH�x�8�ҝY�)��A�O-Ǩ L� ��YQY�Q���?sW% 61�<H dj��+m�!�gb^L�_3�F�2�o��C��.d��'��W�L#��y�<�ME���g=��8T�Mia@�����jb?���4���u4ӂ���t�Is����?d�A��>���u�䳁@�
5�h�aiΏ���~ؐ�1��5AP֓�����!�*8q�I�H�d9ߨt3Z���q�w]��b=*p�+���.���r��Ƿ�{��}D[����1.�*�5F64+k~߸��I��N�j8��0����g�'�nd�������k=5��y�K�C���"/k��(��X<+"��K�l����?��q�{���Q!?+�t����(4�2�ag���RwD8���N �Bw��kkP�4�g�HX�����1�d��{}��d� �$1b�e("���6��)f��ݐ��V�>mw�|��'�ҹ�*#�FH�Ic���*w�6ؚ�r�46�̧�'Yϩ)*�}�	OK��|�� ��0Q4�-�[���=
�2�����R���ɮ	a8��ð;���S{?UY��-o��Ay��2ѰсI��*_����n��YA�<��8^��m�T\f��df����CK���*1�������|F��Y�e�o�b��5E�Cv�<��-�F�7l
�
�j)p0�^ɪ�q7�e�����z�tJGw7â}�C�]r�uRf�̌��`&�|�W� ��x��g�"��WC�'(���7�ru���l���׬�b*&IB?�����LG�W���K� �ëd]L�V�;f���/�:�94�Í��1Y�2��\�:�j>��0��v[3�U煗)�u�ko����؋ tk�;#�'ȩ��2�#����`R�+�W����.�,�����Y<�Zlv�#�!��bأ�ܩ�J��0�f�+p��oc�v�b��L]����b�+Ŷ>9�G�Z����Z�aฮRN��+x�_����ܕ�T�����K�U��c����]��2���U�\+A�B�y�L~7�#9��ÐuZy����3�b��y*MB�<þ  =�.�B����B=~/3����� Q|�VT���AժR\]��e�X��������lZ>�f� 	SV�4���K(��gjȪ�0�X�QiX��s7�f�A&	��+�К��2�YP6�0\ް�<���L짬�I{���0P��t�$|W��N{��w_a�ۊ�u���������ż'6��{i>��F�MM��腖2����	mX���+|��L�b��j���L�2�4�%c�0�s����b�N��a�i���Ud	"G�9h�^p���r ��S�)��<��eJ��	��
i�kqm#�[��!��5���Mx�2U�s :=��i�M���2)�����
w��E6&�W<�}`���e��"7���ٛ�S?o��4���=vB��1'��7M�n�<�?��w���h�1`�
{�ld1l Zn�����Q%|�Vk�K�̲�%8�
������C�~��`��\ͯW�p���1!��}1^FvYY\����b����l���\G�w/v�C𱻇�s�Gg��*;n`[�4�7�L*y�I0לm�l��?� �] .R7>7qpo���3��v7�������;���̐����e������9��i�h�$�xw���8؀��##ƚ�v����4���^Tx�`��S�E��:�ovn���<�ʯڮoݔ4����8�����P��1 0��\�yMY���I���������]�w�R�9�Y�Z�&9Uگ�Q<Z�oleH=�-�ia�3c^g���t��k���?:����?�<$0eF.S�_;�e	\1go���!9q��揅��p{��ã�d�����.AJ�+NF��A5ھ�
���j�F	x_%p�l��4� ��A�DV#�i�2�eQGg�*vc/�̉
��;Ԡ��#�L�:�w�I�do^��<Ls��o�ۤh��d?�?p'�@���=�����?�U�,��]�#3�#�L���gx�Qe%[�0�1&��_꒨c$�g��e��o�G�����'�B2����Lr�#{b*�Ρ�D�����"=�}ONl����;�x��l��_'�э����QF�.�������|���+��[b���A��B���&�Vf�>>S򍶣I>y�!�?茀E�"{WyO�Ȋ�����: