// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:17 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LCzkjWKgeyKIzWtQXz0MqvcgDmw/zplFn21ltXmKQq3tFf0jIR4Nt1qIn5002Ni1
v2xDq7tdKiuO6tTwJL9nkPHOQsjJGsRrt4lRRulvfFvearymsfH53MQSYcs7kAJv
79rdQF8ejV5SncKZzqH3HCEE4rUPl3t4iKB/sTl7Yv4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 46320)
QU5vqFu8boxqDlHu25y686iTjardM612VJlj4SUOkNOMtH4FfVo0PWnw2OKvf30W
PwAFpHXO6pb16XI2otW8sGykw8ysG63Ayyc3aIUN4H1hUrGVVMA7l9fa6fBSXnOv
EoGNeNPTXJSLxAQDF1GcPVvSlNz08gNsYzRBGrD7XonFN1S7RSr4DOCPOO4bnObW
1w2nmkaLnCT88tMXpW6PaSi3V4xE7tLo/Y7V6SNo16Y5tnPhJ8hO/kxig+lZinm8
ENpvx+T63IO6TBLtqCBnYqEmNY0FZ/f553/lTrGc3ivvef3MggmsTZ6FAtTMNaio
1P2V+4P3iiowm1ZNk0U4vUiQanrb9+crOmzeoAdh/pCHq/2gIVvLUKonPWk/i8bd
rfVCxXS7IeLyQoYdrsCYQl4BWjR5XQMeIqkio6fdA0QG+Pc7SCQ4coA/cfjqbpm6
hqOOXHwJPRwC2dzNUqpr0Zbuoeo6eXUfYREXh/c9NbNJlbMlN4Hmor7SZ3i3YAFP
Lelb5VdTkqdBadjbGTRFkn9wksUMKf+2w+uMhHGKYHmVmiXHrlGLxZ4PMPg7D0Kx
lWGnJBBJ42HWgneXz9Hqm6U2BAc1/NLZzYh5J8zx7R9DBiDblnlVNXhTjjFXj1DI
F4uMSOljfFZhYzlpBOYd6F7RMrZLmPdid50pUD5a2Qd7HGo6Xo42Fdra2UR8svrO
jl5Lp4hTFIHYQ6IHuQE6iz+RbOp8ehyeHJZ/n5gpTFLJWDSmKOF6h7w/Jxp4lHPH
rA+ORTHLuL/RoiFUJhKOnhyNBfsT4wnfSIJgtOwOjBXXjnJgGC+Ra1A1Gze8AMpT
nLYlHOq5NxG5pYlJyaPeI1XmQwb2Ew309i8j/dDGDQfxO3jn1X//m3NGCa4MUAjl
d9slApqBneFBKEc5mNNcTihTSzfCvjauO8YOxCfK/hTatTyQQ7pRML5g5UXWBqGL
tgKLZuU0bkjYgmFl+xOC2TUeNlDeZblxpYWkGDXt6QZfOG9vrgNi5x/4AeyGPL0Q
yO4s8raBblyMWdwo5uRZhhGcdTAS3H574WbV6Etg/ugPfGERIJ9UneEKoFnRSByj
henJnPE8OkD+cw/9tDfHOOZzxk+jnBdRdLX0rZhcIGXPXC6Db/hoArRbid61iV7i
ZTInYzNqm7OUp1yU4j+qJAq7fkeGwC2aICp+e50tm7GdN51KyMjhSksr5bOfNlIX
79j55lswwm9RaZozSrsJ24SU1qsc5jyTPSz6wKVsYunOYKZvGKaoGS8botH+jMNs
e82tVGPUeB4wZTjhM+YnMZT9j621OlIjmepjRrCy8cySVPMJNJ9484Pvv92qPyR+
XrakywBqjwYpi/wMOZmBD8/1nponXbGphXgA4m9qK8FVfTWinZ8BcD6sm+UMcDNZ
ubr7umF5AOvZ5A/vMXLvj0e3Tufar2/TOVwJe2AZeegvzODSCqMR3luac/UXEDfH
1sBAZoYKHOxc+opjNIKFCRmAS5NWP+5j+bwfDzxyLBSFq+bCcHvyi6svwsAFvCUO
SghsRlHcg2GFRTDE8Y+cjHFA6zZqb6MWOG7S1XdYK89cSEIbXv1JY27A7RS38qDd
S0BAszmiTBZtLM6DeUUqhAin3iq+TREKuikAoA3QoYeKSwoMNWHpLeatFMtzCMrZ
uJkEXLZoUTJXfLK2FkqxUp/jvHol7Uo/yHNzssIQPD7lLEalwBUwDHB0Oz6FZXDs
ylcJy/hFykY0Wv9iIuEU5BVZVwj3YUaKgvfuff8OJUieJvtfYng/NsJYBib8xgIV
xm554ghUA3vrcPEupW0stLv9xpDKeRLsxP/u0FIRU078onWDIKgWtOWv+T5lL20K
wASyGjFGA5og/VO8z9xfPmvGbYHJxeYV76VnFK8CYxNy02mMnx/jU+A8qSg5Xbu3
rh0wStHDK3e/H8RhkssEIRM5WJ8oDJhJq9HgHfx1CJNUqahKe32J6Eaeubk5OBj/
0fAw8AqHHuipgugntsjeabmRzrcvHjxIx1PwFVjiTyWVUKBbUFrxINOUFFcqEd2N
TWcTBOxphqv57JqfLRezjLkfff9M0cI2ZGORzSQKWkGOYxdWYTAC5s3/0z1eP9RE
Bd1DDEGlHErY4CbGK3nBhNzHZynoHnuaLWH2bQbZb9+ptAv2E8vRYOerhHGDuNjb
e8eC1W5oAbgQ3MhghclOlIzN4n4qOU28oeFHzkytdTTuC6gGvLVC9g2kCUiyYwCT
bY8u3KjSjh+NOb0cnr+ByMgir+H0GA+WKPBNzI3dPsKtHBuvhhYOfCV4TiJISMKL
ilDyaSE7DX6X6vj1XXLS5IuS4n0iECIXEsMfg1qL+Fzs7yAj/jDASj3KPzwNCWEm
ZsRqdld8fOL22TkZEOdu2U7ncTNCm76eyc3eiKIC4Y+gXzjxNaV/sr3DU3srZuTJ
1/RVX7MPuCJSX3vuwNHUMA85mv38hk4sifDtMHQcwls4UVB80bgyelhTd0B/+Ebq
G9wjfYQx3BNvLS/owq4FCGvZm+tjAkXY9b9QbjelGCqjfR2geps7rSMJ5h+2aBgw
mxT3PWmbHJbshgppQ+oDSEWIPN5PRR4FTSeq0HW0YsDhGzP8385mPZyb1ihCEgTe
NF0GBLFpk0FuK2047rucKmMQYUST2tPnSIwFsj+9hZuK/fKQm0AsQ7dKkeJIe/Hy
TIXIk9BCePd6auj7UO2Zvh5KUhwwFXEtZAytcqgAlVIhZ5AKOaQXiiju0Fgmzdh6
JtgnXSarzADJ/X6N014OR4uigW4u3VJqncjtEiuaPoSrlE02CbcjyyXGJnBzYtnc
IMkV8WfyIbD8Z1p2cP0liqsVx8SJhY4Maf7YG5psnZshEsM1Cl1RFgco2Z0/hoHH
ZtoJzLw22DL6Eu4sH/e7GoQlFYwDgwFkuGXRgZV4877Cr7two0OA92YMrVcl8/Ti
B2glLTy7tXz89YVSsxigvBwo+AJq7BXCHF0Po9G20T9qYA/2zayDSX+okIE+uo0c
kKt6EAzq4W0VPlcfi1FnP3qTxqUu4+sUr+Suit7hZM2lT7XxzmK3dT3bEl5yGhVe
t5Ozq9DYmdYUmNcPXYI3tZo3aStQp6r7FIrh4H1issaFrVJ/Q0VaxGDQpNRIC3Ym
VIJRaRFufLqK7vyw/84l8hh388098sIGgPHiPc0sewA8Qr4HGiLJNw8/a4UTIPZJ
zjGQQToKsAPfYuMRZomepLKq0A39qJV70uqa5iXzKcRAyBfnruigXabDNFaphC9c
8KGx/eoe85bQv7qR6Knc6fA/SKuWQ7wJv79KTeLRgmLy4d3jXuEMv27D2sjf9EbE
tupDQFRImwARHWHVOls0fkORRmcpGz3Hyye/m0pZAW2nYEIltaxH4gqhOW9ykqEQ
/9PXLUeVQX3mJWJS76n+3eHCFfZf1qvghhGmMwiiRWJBP3GdhmDYN/fMUw/Wna4H
8NRYLoFGviueZ3R5rOhbzC929vd9V7NClT7Tjsd2jDdDyOgg47TxzZwXO4Ql9j2/
moxQbfxqs0MUocAShAWJRnpKWIRUYrGj2JBf4/+1WmFqY61i4tLx2TZJZhtAqYl1
Jq2+P9aBcT06LdP58Qp9dQRRcjtmheAkXRKdu44TYyVrjIB+Z7waQlrEF6NhYOpK
+nl8gqjWWWMz1nCZ97QdT6A4wDu8YLjj21RBhN46FUluJQy1FEf3YmTB9TJydLAb
B3HiQIQX2GKAo8MY0HRVcc8n48rrpKZs7gXlstRTHHfaUP1egQB6DooCHwAmXS2D
c+L+sbt5NQ9QU/GMv82aOuhPSbRSJ11XAu3fkJp9mXDB2muC4+vHkR0yALVy/Bji
x3ecUjMplQqaa7o66tsOJuxFgwYxGaiWGk6E2PHEOj/zezw/EbuCVZCIYL3jEDHK
tKgQF4G08X1/bgJjCdpuAIL0LFYbp7sHt8Nf4v3r6JsVsMqbc0krbxJrcDmasNBK
K7J9mkHtK3aIQnl/hosC2uLSO5O7GoeDxRh90l4c984Urgxh3cRYCUjTtjOFIjkZ
LfWxvMSJA4Y1H4XfSImb+4vzYeV+FW5l2Lm6TtleH1crfmP4srXWrN8utH899hLt
VKq0lZhJWv+FwNY72z39AzWDo/Zez0KlfX3IOVB7FMvr11MaR4AaoGcNaqO8Wasi
thsX0e+MIVf8VmuVjXLy2Zkz3Rjy90JcfTlxhK137gktebMjk3wlIZ2ZVEb6Q8GG
fmQh9A6QKdeg+SpFQaMJEFQEi7vTN4DpkmrG8H5Qb/vIM0wFnEB09GSk3W/1AKix
nQFrA1c5Rt10bvboJQQwvGatch+2hzKiYgVWo4Gp7Zv7Qnn+stUy9+Kp/cBS2eJO
CwWBxRKc1czu8nXeOUl9YLbc+q05JcEA6Zp092np4L+Yb+Ps+696dIzMDwB8FJ7G
MsvzGeywU27l/odBJVuX0lLFkKThbViOOMGMJflkq3X6uxUW7Fynx7r7vncApSwU
3jEDVGs5r1AhsxVogcfGqiqCt2KArfMDwrNZ2MeAOzrb5ZRp7/s+sRJBkvxEEclN
Z/MoHZ0/O5v7hk+pKUfBn2rGZmFLrOW2h0/D+mK+9uAkRri/HYupUcbQScLfMklg
QvCCCdY5rY8kJ3qMceogNms6jedotgAuLKS+Gy5cDWjzgvHDM6P7wqKIHz9nA+ry
PhaKnpvBgT6qlssJ5Y/D0ThSMrTWzmNZL65yS29dqcFOqVP/p3Clim/uXbUcRgnr
tLE6fSHl3wAN6qENn/STW/goik5De4PHQKDcwh3N2G8XYPMyzpN7YoTivSULB+iQ
IOYXsLCruA2SJTQfkma7hGQictBOobOeFm5uEfAAGfQqanwErNNj5e2dFVxafdOb
KJJo7vu2Hnwm7w7QGJLelFdduwT4HIN+qIqJwfp26NaODDDNi1HfPAWcuQSZAw5O
LaRLa6tbCJAfIiEn1l0fPyj4Tx2kJWzeEgfAJoNudl20JYe701obX6SyerWiKjPd
EuctGtoCAuNWUNCz33Ux1ghSOZGNNQVVX+f1bv+zGcp382OOKMymTk9+0mn4WvOK
R4V79cS2W0dfmXKXDfAxuV3PrKINzYs7JiHL3oBaATHp/XRrsNewzRsTi2ucfloZ
MRuch0W6Hgu+6/V9J7xidMvUA+seWZBn8oWjeEDqzgjVg0F1Lm/OUzxWhDYDBcg/
xirP9UGjeWkVlyeJpo8SE5Lq3F9t6G6EhnAiAqXbVCS3vhYvWXs2PLFchgHrW4o9
W4NIvO3tNVmKzDBtRejLZBQfue41eJZe+Z7/KjOqbkqZRwnC3N7tUNpsi+p8kJ3/
ugAbGjN6iizLQdHK/K1gY4j56OARTpF4a16DBmJyU9ihc8OZXeoLJXdAC0j+56JN
hoFxoGHyN9GTEAtAqsaKIastaRZ909F2SmztgxMD3kMwIffqSvwm4unfuIlL6OMu
e0tUVh6LfJ3cY+ls6eI8X+MGEnv7EbCmJvRQyPx/sfdXLny+OA612ZQlko3KEAPU
ljpffrGCSax1WfOt6vKr/riSSS6a5BTdfzcWKOvnjjVu9SvzaMgbrxbkdykjx+Dg
LyvqvZREJz4HfB6p0TQUiotFvjg00ExlovxGa+smV+E53rUKRZx0BclPTDqAvBpP
52sNE+AhCzPmDBytoYHjvBYrFyaFPmCRbZ4dATkUGlLQDLkAxFpyn3KfnF+2Sou3
9nD6dUrmO3xoT0w5PxA1Gs735DMg5zVjvv2zTlu6SaL02qcZc6CJYNa36aYASTrF
wq8EMWHwL0QiHTwwatzsTGQtG2z0REtMf5SVX5byo/kJo3TqXQvuY2A3/C4JDs4U
hRd23ZrKb03HkUeYOaBTrmQV0TslWjxhhuPD9l9zwZAbgHuYxcHv1n95dbCgy+j6
aVWiCpSmbKt6gqBC2owakbXazmw+wUkLxC01yh++gGgWPgQYmZSQy+YhPMhxhKRY
UAxctN8Glpk42nrEvckoWOkb1hHm+ekYWuJWijZEHYkdmgSwE35xislSSHynFcA3
VQr8rWzny+B9BWkmjM08ye4wTklIaIehAd38qyVuT5v5cUuzunpROVGw08Vo9NxH
QkpZgehGyXUFEjAKvuciExNDMl/pAbL3kx5SDPGWniQRyv4efEge5waiR0Y79yPE
VEsPAU+AKEeLz/x/hihmIxCdPozwNQe/liG4lsyCrJ01Y0nSivcV086RUUmDKRpb
jbBeEAd0evc4DYQEuQrj0ZDhy0VRQw2iKfGEx7VEO5LPWG9NdCSuFGzf40f+oJMa
M7r1jTRNehRiwxstL2Ic5+n9ypOkrFM9oQx/jFBhJdDB5EWdqVc3ZCtoQdpg9RrH
lzgqmvn5q95c05qr6MPqMpu9XRZKQVehO3tC2QQzx1fIbdGr9c/gM5pHMmhzMJhM
6bA+0eK/V8ZMOLuOO6QkBdDq2PR9aeyLUZtgL4uyR5pc/cCZtwh+bcn2tWD8dQXu
mPMjOQ6IjRE9Shx9KNTt5TFWX4TgmhPnCDekx5/Oo4Pk7WnSCw3v1QDjvNOwbEhj
MxvgnPZuYIaw97RvRIjvVA6In+E1zOduSaL/bnhk/l3OV/+SuN6XXqBp/JEIZiqX
nksng9MpXBbXv0fVH111RMnop9Gy6QXzb4z4vr2DHK6gYbLn4dVKTHGs6u34ecXy
JZPwx8gbNnNesBOpXqI8otZrKjJrm7hgB8QwJ2gFdyq1MOHCKbGbED5u7VBG4YKr
b336LoOQ4LYi/LwF8QlFCE5K4lguhFMVuovXnGbmMIaP3CAJAlx6PbTZgj9rCSZl
33nEpurBI+lJ5V/9sbiIE5MPjQcW3pAVGBzuQ7IgWJt+NwYZy4r30jYiZtOX0AuS
zEvManCA9fyy1yZ4G/B6m4yKqnP6pD/6YrhoaEYmvP6v+G2ewbUD1r1EMRCCdVj/
7ZOUMnS8LfzOwvk7jCxs7uS2L2PgspdonBET/IFjk+dST5XMAFqD2A12zskX5LzH
gfujK8y4VesJEPpF2vbLacr6k942UmFtqcVsuYJPepJ9xVRA2NYLwvRWm7+j03J4
GRgdlMashwk7rdYWujEtt2J49oMrV8m9YDmXBXnlTrAxaKy3NfuYAypL6O1WHgy6
ZbY5noy34SdhKXnCrjWgTNbD7JpPlN0K67wyQDDKcyoHh6+gC1YFw8JVqZP0LgS2
yy8ZNlNeLIXIgHGk4vjs1lfZL3YK5DYnkh5j8nsYHrXZI+pFx4yZlz2m6MhjDezh
4HyX73o8lnkE0jRlJ3B8PEFFXCwL24wlV7XSCNjBxihMHMcIg+HYOOIFIBvg0WZp
GymyBi6kxjlFDwhdaFXmrspoSEGdCbibE/g65wY9wwMn55u9L73xGL0bHR33Qx94
3oFu1NK62H8qZC3CeOn9ls1qmR9Rn2FRuGzyQeVtuKah+kDmdSX6RRgCfL0LNIMP
/Yn/1vPSVZ31GWK+XkQZ1C1XryTB+0OcbiHld5wLrnrUFiutKAIa/Ry91XdwCsKP
HCAjswmfQnXdSwgZ+vIBi6WBXy9UBps7GDHnFowf6bnoUesoOMi5fAJdUJG0y/cd
BLf4AsMAB++nDfwhPZYFEdpLcL1pZyh43hOAE3LfuBVyfvf79vu68TjJMPCP6qek
h55m3UQEaTMYZOSSX+/wSLVIkS0JljWwgEdtjsGtgN4rgGuSzE+1VWngkCL0LEeN
aszXtzc5aI82rxOM7cfk/07MdiMcZoPrpni3A4LHpOrl2YMKU6Wm8XvwY1K6p9ty
oouiroN9r429SVoId15Ih+oTH0L6SAjt0iKeC0YxeoJR92iWu+MSHpxUJgRb46uX
2cSAtRiHT9wgkW9IUXcvY9w4hJS4deV+H6fzS2lskshRIqP5ICDN/F6aYPugjee1
YNiUHRcP249V3myXjyrDJV08kiV4RKHCRjIv4LD9hNeRGiLJSDix9GflUS6tfL24
AUlhhGdxpKzcBDUzsiSqw9UiRSvSOZKWRcW4cyEzDmMgi4M5K1UW94InMI/eTiR9
2hmMEuEwoKQsGeRaMxrbKBsgISjeP9E7Bvmawn8ER/gUnXB45e3qOkTdvkxdOK4U
Hm4xsVGg3fNeSREG4asFTJWzGIbIueHYXB1DPJRChaLHQ/7zYesDZ4Kc9aDu8OWZ
AxsI1kx48m8DaYkCt8vRMePETfYU2Nxxx1HHT8aiX2xKAlEWv9mEIc9RJ+Kx3dEu
dHZgpTAUUrB3WbYTXNxbp7rnYlkEp+F4ddBgAtm9vroadMVkrb/EPExYYxxYERmc
yhLWCtgQKoUSRfqIQYjD5TwQvpLmP9RU2qMYrPisCukil0vuYjM7OgU3DY4ioy/L
JHqWb+jg6HZPabgPTOgi9IpbIAZHrHngg9xJRjqBde5xZOiUTGcezjql5teM2l2Q
kawQOhRSvK+PiAvVqxBYJ3HyGmVD0tBFAgaMxAelpD+yZ06P60su/00VnS3W0iDX
HaZF6zn99o0hSud98ToL1AYcwK5HjNvE/wvWsf7E5CDm00e5MNLQLXw1p+akgzx5
6zeLZmspcYcFzWtbtvnlWjkBr9hl+T3pLSRmpRpamL/41kdmVQL0mhB/0jo3F79s
a7dcvN0MYHNSDvQ3tirC/8qmr25Ds8O/8jrROM2Y7dwtOtIDbuNDeqfOR5Kp1C1c
Dz1G4hj5QvIQe0MRwCt78rPil606gGBD/uqDcVgm4s+RRVWqiCGoyu6GqS7qgMq/
DBRfDvFKqRdBfyZuHMY8jxFgflOafRREn9S2wm3PVFW6PQxuG28/aYfBd9z4F/++
r/0end8VMc0cOFQLoIMXM32o92qlCop8SKWKq8DXAH7Ik4yecJ7Xp9VPBdMH0sb0
98nwCmQ8zWEhVd1ZLlKyZukOfxRWJXT1JCnmPM0VfGqF9qQN9X9sfmzOGo3D2pRt
bd/W89TwhcqBY889241IY7bqVxfF8+qP0subG4v83AilFUUNWTLVXcEQwJwdc3KH
lLyTf++TdxhqG02tgVjgKIH1tVAcuWTdqYsHSJHMo0XU2cvFI52CLIr1gM7JmfB5
q2yKwMbMejsjJCS3oR4MsFSeJeTNwmbsdOn37lfrQ6MIWXipdlwv4y5uKeC93my+
YclbCV2IVQKQx6p+vKcgSRLfmZ/0NNlykcnXcc+JbvUp3/hI+8Cja4SArk1rW9VN
oOb7fqwDjajXJpL6HvtG3i3BgCW/4pdfcZMJLg3AeLo+xydtm855c7IC5LLjgAu7
3EQwD9oNwESNVeONywRJGsfjJvyBNyh6PDrjernhJfNbVGkrN3YDRq8uvsTtdr76
zesd087iBL2KtPzxBc4VlPg2s7VIEWaeI2L9bjlM7fhsowUsiI//BeD300M8o4WM
EO31AcqDouWYhUZvOxpyI8ABgl5MZhyoAQEeDByxial40D0aIVJXo7STIETOzrHZ
Pe7fETNTY1xv2Xlk9vqw2bKor93xfA1CzU1HkaCd/wwvm5+6jB1wfxdJN15Ffsea
micA/iB2EgcNCJr7RNehTYSE50edAK4gEA2TFKdRkwsgm4/9QMj8af1wtX1U+DsT
c5hBw7fz26Uu/6lATfqsbKDYCSwfkzIaQItyILsPZ3pM7TixU8+BlGU65XYeO/lh
+AqFkm/nXyubJtc8xZz4fmerFHcaL1g10czuGMPG82J+sP4xR3OTtttUKJPCFmU3
LBZXPgZc6SOZJlVwwgJ8KRYYLUYoZpslqyET5Q2fxCYqputj26W/mZLiZQcN3PuS
SSfzzh2kTOyQr6RE21Qy9jmx+QSWSGV2AbfGGOm4MdcgFOsSEMCyGgiHjG9PedJC
zAe+n/zUn+AnUfb0a6Jk0C6dk4kO0YvbFPF2UBVZCLEj7Z/NfriDwYwx9BYnrtGN
estxB/ewbQ/Y8l8904yt14V89hOKVO7/5grWc64AoKdS3kP3btWPnOn2nPNSPynb
LTFbA+h5Am/qJSNvxto8OZxio2rXTMTbjMfAcuno5VN4i0MO7gbJDk7PR2p311ve
BTXtkv3g+idNfC3wG0kyKE6yaGZorA0s09lJJo9W9o9FBTjGsBXT0WC07Z7lLNIB
9laIOGkpmkXC1BkPUzN4AFx8nfA/5H5WyCjjJfWqcADdn99ekRmEC+Dix6hYQxpv
hod9Z8dX1f3M/zpy7KOtSwM0YU/IcLH41w58ICjBDDKPI2/7GbMlzRi0H/4JtgHz
OCvEplpYyj/D9Q3CtDIdHrA1m4ek1AuuqeItwrk8lSUQfUh9Ok1o4vIsU0k4/8oq
bpOr4jPFLI9v/uL+id4kTT8GYeTFPyUOkajQ2md2XBTxKb/yif2vFYpqFW4mOET6
6NYUMQkryC5loFquCqq7FPGyLX1PqI+c7q908KlVIP4Zf0VifzBOU3A+8P91vHMP
/9ZqbC7oLz/FS7xFZSR2neUabj47sRfR/z2VzSakPc3/+cFSy82l9/JBfQz9vLtD
MNy4TBow01ZuxeFYTt21nQec3mpMTW2SPJBuTZ016XJciGi6XfurX2D2IIoi7eLK
Tsc7HLY6uBJkEWGJvnvaL5gJfFaf1Ba0T8iGYpdo5AbEyg+v2pjPx5tR6EZ+ziYp
/GGvFX24C8+0rTUDRhahPc8zSFNTcSDS29qx9KUno9bI2WZ2U2Z2C/OSK3TW8uNQ
NA2cyTt5KPjdm8hLrqVTHNlNXMNWYJ/BKwdzIA6RoEjRxAfxufwzo7m6nwqTj7FN
HkcLlV+Xg6v++2cndu753JnQKl2rbkESpPLPE5mpKp8cCKfylc+nDWY4w7n5TRBp
MIQmqTlbGzi3mOotkNi5PHw9nfm0CjTYOsrMAlVrY40LlLPHlaiyY5vJksq12eld
UBJTANjCXf/GZ3GDELYqsHGavHahqhU/b+0G4WtyD5NNy4ia8nfXAizcv1eSVVPm
hvCYhCrJeh7j+blhr9KP12++TSe+WR2m8g2nn6TuRFgcMwmiVtMri0Yg+Z3AN+Zr
KxEBwOKj+OXu0T76BrOrqxKf95bbgFuzNvioSTknebVJqygMPWnosT/LZLI/MFqq
OaT8xrTeFppEDNoBAhRE54LTkE/w6urBPfWqSysDhuLuk0rpce0noplyvZPLE3dT
ORPVNSEHIrYqjyz2mzZIfyHYqf8xwxCDvIbZnBO2OkdKMWJBHHSq1jtPSnO+zHQA
iBtgJgZoNekdpFH0rIw6ITRvaA6N1o9PmFWU9JRsN4HgWmiMfXMET6o20YY4nXWr
DiQnMCXS7UoWWwbSURBUw4wSGxwC1cVQAyAFtIDdSezQ7Fnrinr50MwYr0KyUF5M
lyQOgtEFY8sk5ndNV7Mlbu7E+VWRiH4ac4IFI/t4T0pWFAvjHU+vaWtzmYUc0Pdr
Cq/4o8MiXk6CY9IFXMc+NyWjhxtWXIAHstINw4PESqIDOlmtqyOV5MmpH5i4ZnPD
OVsTLvD8YyQqQ56SAciBPfkuklyMOCB98M16ngM1Tbl7k/MwGM7SII/lSjTlh/EB
/nNEIGL+kJBrZMfIQ5v3V05wDQbeEOuC6i3IBZnmobjgOjLhgBpXdEwLRemKqPDr
q7eUTZTk6Jz5iLR0sIscH5bQKgirj779QYAZa40R0jQ+XZ8cd4glT7Li73YvMngT
aqh8hWQhF/RqD/73hf/WzOLo6Xfua3HKvwrU5G74wR2vlT2+tHY+/+vDejaUu3EG
E1WwQmoG67sbLxAdgq8AvDSi2HNKugWiKzqgNxXszEuQutzLyuPrluU+46G4vVh3
G3n60qLOiKgcwf52d51/cZI9k1dvPkEEZxZEnV5CVbshXKRqcGfsIz4rbZbpZyq1
76dpuDfF+58PWJHccg2BIO3fLxqz0RIklE0dPlxRaflinKZ8tH5ww+EnxRZoTlFX
FTb3F5+ES6CaxXHGFgjz/fkpFd7JLEAwYJD9bBqZ957joz8YyU4oLZoVPDLxZUhD
4HXqL/P38XPnNa9CsqX0Q15KEm1ANR//3N/UKp/NPFsRU9sCDWf/KlZ0zlag05TT
s9C4W/eWXv3r5AXqeoqsDUC+nPaHfOoNJ2xnlOgPPK4TDptYPKjP2Ian4u23qCUU
46fsrD6akQMCXhunk0kFSQAfrUQfyqASccJCF0aI4qwKmEPowPtt8IMzgy4zzADR
mTO9+gVr3c66PSmD49Bu9FR5MHhAtTME4KHyR6Pz5W8f738K1GBgIzVyI10ABQZ3
y4c3wd3kBl/Xh5wJm8VeZGi8JjZ+wsgQdPQ7x7waRVAR1vEx6xEeuc2fz3RT4Vf2
u4ToR1tsyltqH4Yb2WBgR9/MVCcEKo4v79IHRCTqX5vtJ0T8upMf+YxZKK/AUirD
McWd9rFofZTfjFGwb+O3yt2ZrVk50Ch+MK8tv36XYFmuPt7TSgD3Vriu3vLNz1uf
L3c4OSUFqGOIgkKCyEHDfUvBYWrwz//3Kw7TQcWVZVyv6ugUVWZTrWlxqUjOU/Bl
3z1DppAPWDqbU06G2eVtmOAa20gYw9ic29I0wUrJcejSMuHw2atVyyzywp/sU62C
S2zsXCXc9OgJr/BoQaa+fKfBc1G0deMgdg6IN4iijhkR70oKDnQIY8Hz/kfIUFCC
cALVmmWMzVe6RCRb/XonvzCZzQUNPeOH+v6Rsd1mhyTTkTG2QbVFR7b6TVI4P/j7
pc0Fa0qnr70jbnl6tB9C2LDZ2N8/7c6L+kY1wBjK1DrP1rN9QU0OCIHu2vEh7w8L
cRgk3XrJR3w7e7/f6gi25YhvfGkPEw8UW1tUJELCgZX6PMPDYDCB211+Hl7yzruM
mL/uyEAOLmX3txbRwjJCqOZGxQw7d36WPBqcxm9hVJvN83amWIL0pEnTopsqiPhc
SAwudMoevx5rJ40xlguW207p8jdgycPr3P/rPEeXV2S+xF1mm7+ZS32McITGUdrL
c949uFbAWjCFGTPdjne9mC1SY6zCInvZM4HJUudZ2I7yzpcMQWK/fw2kXXLOtL8a
UYyh55TMBBuUPjryyu+m/5/qDgQBvjQDm3w9rpZ+de+W64WNs9tOIOYsjPeK05Kp
xLpcg9yjxvtKYbusVQmz8X9F0+Wo4nnQn4Q2TrFsovs9wI+3GSXZBnNebdEj5/Mc
6OyteKJgWvBvZn2y6ez5Dt3NjYwu/u99wyMCzO3PrcftD9WP9CeRZgbMX/CGscqj
w+K1CHAst8J75sK1EcoeBteX3SvZt13mf12kTpeBQwYAos4lgy2BU+URmES9UMV+
7jADCa3BS04QSr2DuAtY8ILgA2Nl49nZwYE6tDWaaFKqyp60ZSH0ww3miVsUDIZm
i5tlBxYD6Os3oesnY9lKvu3sHfNrVDc/thnrp2n1rkL9P3ScQBMuipdfp5Jyr65f
vYtIX258hjwI+QRlEsW2uL5d3WVN33VOkHuELLYJstVmeHjBpvY5qKoSzryAJ+Gd
Bp6Q2Pp77CJN9JB89HDmFru6rVnONjVv179AnNsgcY7aqofNH76D5WSyXck/ELUJ
YJGvCdLCjvYWLoqtfuSvWIVlqau2YWWtPJ5sKY1UH5MJedp2A60UYEafIDuo6Mlg
oiTdb3wsceBYSF0CDf4BHZOrZa3DMb+xUbmYTbw4onkmPyjZgN9Qjycjo52HFx3c
z3T1pG2VUYTrIIlwyqaPYVu27C+/rhGhEhheYcEbaFZ9gwZypR6a2g6KkrUDR4To
WC/vFVrvRsdsz0RNavsVwQ4mtLZ2ZhroSb0IkUSrJ2U6HrYxBnIQDMSRqaOnv4wb
B/VHKkDs2n7eN33jfb+dqsBCcmZdwJvmLKlmu5KboNukRSDK3jbTNieUuAURJAIp
QRW9xsBH2/WdtMA4KJmDFlP2YlHKw3F+F+VRf9pYPPf6DezcwHjnppA8U3CXNKzp
797p5Ddc8YFh8RwzA9iW1FRXYR5eRz7YCm8gD5T/RWbjTGAN4A8RX7kBYVXEa66G
lEpkJg3SlC4Cj3AH39ZfxwC0l+C15JP8kdAbJQ7O4MM/IyOv0O01juEmmB+uf9Df
SHi9CqMmnJpbYK9Vchn3uKEmXPVMlmp4rtoch9ygrBA2GCx+Tsbm6M9jZ2fFKSKs
LWo2IyhS0A7uZhZXDvYzB9gdAzNJsjEu9DdFwB7g9VxXcm5jevGN94TUNlNjGsEc
deUlPVglRGQ28fuwqWtxiZzse0z2tXIPxvSfEjm5sBhaG6LC7eT1zx1Z3RYUlodD
CPzCg7awUeoPgMJtefwUZ3hFh34X3l21F6oopH7Z0lYX1VoDLk5QYKSFyvZfwPqT
favXnEyj9xMXq5CmhEmGzl+1HY52nDBTgZAQBnxFEsO+YqaaTdwt+Kg6qayoZnC0
N2S1eTMw5ijUWmgadju0+Y+QVy1KnrSNAfDCOaNslLmDCtNI4K+4kkIxGAHlIS8W
qCn4sNQ0SV3v1srEDi1EHfpDZZCfuDrEA+Fpeq1b1fcLf9r94fV0Nj8gg6++LxCW
zymEWFIIRtxao3iAOX/RB9qiA0uhzaFIPKCxnRQvA+h0Dea4g7dQuJ+Hn6GQdco9
xFlcVw8Jlbi+Q/+V5affftugCfXWzudrNoxJcQR9RvLGbtVecjf9hDtNGS5UbXvc
RhBs2GYYLGTC7++/4PViVywreL0H+eY39iTrrRXtAKxAt5O3yAU6o/N1BxqIEnio
YokaO9GvtEAjVfAwtHPyOpcz529kwvx2etyKRVDqoIXXG6G2vkceLD+0zw7qlO4W
yZCzzzvlUcQULUEmzVrmQRepl1+iNgR6xJLN4ZLYNQ+4X/+CuFOyx/5TCy63Sa6M
EDHNuZqriHIyl0j/AEmZFhqyjIxRTE+ijVvEPLYFpEBXO5t56Z/BGVnBJ22/WbLA
mplGL9VqPOp2221WZ0mbuDa4RM9/x/RNOr3tZRKJe6PG8+g51QmlhQaTg3xx3Qvc
QGHJ1bIeZUYvEKxCNQfZBFaUzQGx0wG2lnLyzmeUleGTLuf4n7Uh+TxEfIBm2k4/
GQ0D4wPGcwvhp8nLXCpOGWeKLMVwaUYVU7gRQUwiAPp4rrgkrMj2PDd7VuaFglWJ
ifpX5ALw377lYNg7o98ChRzhNzq2s6+TNSDjSnhGMhOxu4Im48tn7BdoLI3aSBxz
q9ELR6tyb3mVMUvlDr3gTj9J0Ut4klSMftoqcKt/RYrgs04NIF/EGkE5aAqEjO+j
DGCr9cGtcX/NDvZvpXOcWggv/0wKv11OVlDplVc8PeJbsIvd1Y/9Hi1zr/s7iXfB
0aqlW/stmeBz7E29h7twPuFqnCRX1Yt0AmESb6tM+I/Jw9Jsf6sQ9Gz8dODkrHBj
BWcleGBxTqk6kD2zZljzAPG14thTRq7W50RFfkhcgv8gb9HrKOUGaJoV8N/q1L24
XlCFRgtp2uOWtsQgnBZJGORqRQldjQrdoTb9NyKfyEuGZq6XK9Ewx4XwktIMf31H
tzEmtVzfjtnhe6OMIZbgZCwMrZ3Ji0abNfuUclNLSHK+zQm7deQ8AjIo9Ejc0XFX
P0lixLcsUMjWzhZW3dqzrcb46Wi7VmfvNxYsUV6s/7nWttB+EhPag2Otf9Cfgtgh
Ma8quG0ezUJu5f3LZJ0nju5+OjXkmJ2M+eUEGLWb00k7S2FRlamQ0aYsq45IswH0
G3fYgd02/keOjDr0UuO8TJCwcTCxiUFGSb52e1EDu5ZamfM4LjmShSJgKPU+HJyU
JpA7KN5/qA2d7BaxKQJQzGY5ZbZBuJlU7B6RW9v3lDsGAJZ25UjZ3SSnCgp+9M5N
EhPpix4NjL8OAun9JUrIf99l0Z1Q/MdIVnucIjG1UMih+WWdZCZf5w+3chwFKG+y
ESG5ayZveYpp6PKfF42FfPewYhTTb4XMa3zYXbW6GSd7xwRt4X97t1KnMIdKFpDy
/zZlELSv/BaU0TwpHn42lm78xrX7r7XvjJPfbeQjbfF4ULZrJpHhEtvSl8rZeXsq
L/3rMtfsRhfiwPxjba/zGUxcxZQs9GyWdZG26sGkfjGDrMRRkKAXRCNebtPiK3RR
zeu99Y1m9Xxhh9eKG/JrGYG2oKbLLZyIGgWwGy5uFMAT8IebkX/DQeZiBUHvL2he
Cr5AoWD5sMoRWDmIIKduLx6T7emQwYVY5fOPC4WfjMr0zOaB5rO4dCrSy2NXXV+N
VUCyoYwTSN6OUkcB4PIEg5tXBePkuK8JyR3Vj8ckPzGCFo5OZcsR3uNPrAln+uXs
Lyzv9wfRbFAQpMyvyjC3eb8oF87ntYzsKVK+jWP6KZhMrmGNYutT9tJiJwZXnjg1
JKk5zqGCbesiQzfOLXRpgw1KQQlTZEpmgsOUZp+tOF5Ru2wV60kUXjj/zj6kgGva
UA2tj1f+nUeywitJgmcIQzToKjydhYIjsqYfm6Pr2X2oUVbTHITyl2B3S/M7joJX
+osKKNhyCi60evthkbJSU7g94mJWYbmjz4H7I2GgA8fRNCscE7eOX4AUhzdiBtmY
wS6sW7Z0ltVoYEipqfJG7/d5nqkVfH7ZJzy+mhYU2bH+tVTNeoPNDhXWio6YmKle
qXhtP4sXfT5cFHzsY6VwHrUnaPtqoKnFR0jTyJbfqOUSZaL37ITy8zt8ToeHCBBB
ARKSCvfDw2lGqIa8MBHIKCU6/hVxiSVkgHE9PZLmRs035OvYTN7dLLUmETEi9p9d
AnQXRm/CDXd4JESbrOpVygTrAVVgrTi8/1hFcABhnjrKkG5mOhqjk0KitR62QNPz
BBbXehWAFDXvsrB0Xjr0PB9dMjcVhKi/tGOCcyphhxFDkS75x7dS6ld+eg8H6+h1
96zqSBBLV+AGqtE8JCDjJRugyWKdGY2SXswwFh9tpDaSmhcW35MQ4TDw6HOa3OoU
m7frIXBiHhbMmBSOPNREF9/hxGy2RrLRN2Z22B8BYeg9WdBEouEtGtnTLGWSJMQH
LBlNeoXfWZDYYB9dMsdgQywclWA/nRGQIkZ/h4+FhY+Yp8SaHsv1KbJTX75UV4V9
PJzePCYlHsyFpBZm978J0xKJ0c1QOQkh1MO068dGj/j4GmceqXcIAuSSdMV51Q6D
xZZk87pNYCHKbAG0Iz9URS3Qsu1i/aO7qSUZPWjFvyfqhWR2rMh8NhMxXWtGvfX4
H0m0mM8sZHtP2ccJW+f5Vhl1ulg7NNo7ygy5BHQ6mE4ZMBwVgoHa9rwkwgm7O0Fu
60O2FE62ivnO2lwUwZKTI+k5Xaz3oLjGXTRWDMAglpr+FPjgUu8TgJdjHMLdBO7o
fqijjF69CEZdn9aFU/VBktsumRONyUbhjOo9lziZCHUuX4w7AEEce2hqggLSD7Wa
ezjJnhOB7ivfBkjA9ZDHvaLPIgUP1GQHTssupdErkZe8aJMxlKjMOHUuLz8fzXzO
KJYhnQKf20PGlqx0sZYlX5Sk1FjFAnOL7UPdTshp+RiOdYdGYYrb2oLio+WK68il
/qykfQ/Qkp41yvaVVYkpKFjBQLuTwmloc7uw1kMZvR+H3PsG/uhNOXIwpQsodSUR
Vr4hFxTizTBze90vHjDb3jv9m5k7X6RGCs6PWy1KmFZuONtIHdcGQ2a5BPQtNorZ
YJ72YL/hQ9RyzriZinpWoGKWIjsungpX0nO6JitfmWj6kup5z29xUWPWCHyRDt+b
LI9N4HmDP7bIQI/22CsGqgB3IYyxWNvEgg7zaKi3fAekFXYQzMjRzIOZlQI7vpex
fumxP58/KgqkedzxGQLt+zXr70clgbV7k43ksQoqx/wmXmMIwArvHUPUPlmGlKFw
Pw5siKiluLLi9Emu5yKWlkBXTYVGgCCBqjDBS08j2MITC96kjEJQnzbdBuhnB8uE
ZrwfMIX+9gwzIgrOae71o30qmLNTIkNSVDpKpMAXFLS/kngohCok03+2oFxZ0AM9
eZ2YcJXLGl6ZN7dnJTVoavFQWDI5SZxgjkkKCOsTZkWU7lRWegD4IsKPwcvbmTcA
CXpR6ROO5OVlRyMc09R7M6Sxb5CQDHciEmchPJOVWZuAXpRM0wlGMoDxqGIzxhO1
yYX5Jk752zS+97vR2SQqyRbI/P+DerGYrhI1s0Em90ueAwH/93uxfPE+hp2hOjWj
H74oAYIsjoyeLbU68xV3cPItyCtPzQNmBiL1nYMU3Y6kst+8A4vcxaNqCdzn63uR
lo6VT/HZ9sfC31COp/Nt9dJ52h8ajn+9LKXHThuSEqFAgo2Kt4nPouWKQ1Nhudc6
ZM6wQU2UPNqEXG0iMyf+osUHyco4OdoiFJhyMXMxdlm6/+KBUvrYzIy3rnCVBPs3
Q7yfurtrJCN1EhWFCNPJAbXvXTkNIvXSx61sXxkOyrYEsBhRXw8+C4Oe0vMhuRdu
7VEz4zHBk0KRGrSVbpNpIrJeXIpEDDM6EgTcosRgfLwdpqkFaK75JY2SixSAmx82
vQy5WufODykghq6qyyOc34w5/iXm3JYo5a77YrwzCQpYJAQ4KvaHhJKew0q1suoQ
9KgBrTtBfy/pBC+IZ4ww4tUXv38JDWy2RNx/8irx/dmV+dbThdXc3rQ/mOttYTAj
B3wYLO5kQIHVYCBeHJKDhI9OP7er5qz3VoUkdsgWOGzNszkXtn2bNpwo/cVyJzQE
KgpObVft59sdBOZtmg6vwbhuMGZhE1jyytrXU2WPO4UIYuLRhMKH/hJtlhC6UepJ
IySBDCsobu1RkNG1medq5lGWA6Bl74jxX06q+UMGfSTgmRQ0hTc7WIq39m4zR33k
peEEjpTWzxnx7h/JX4EmPLpWtr9bqt/va5vNbbG1nYqlsC0d/gXy3Q2YCpFdFwHc
j1rXkzma1/UvTb+EvobK/nj73y4ku0QXxY7+zQIzSMZTnMjtCXo3eIKJ9xR2vfiD
vBMZO57KY1VdWYG+toXumVdcc8bDgY/k0rW7WMsiasGsEbrubojxH/Es5kiPAova
YInzxDgvnjaGyvlkgoEah4/cu48/UxccJwzQ7q2YWBXou3Va/cnpr5B5zRksXBIC
1k2PpPifaiaKkYAiQV21jlDr0ZFcNzvS93ymTBjoL+FKcK/dJ2dJtfdb/dlyya7x
PHBBr+nKylCZCTWw5Idr8+fs3ob4GK4oaewJKKdAmGgWu8wHukq6KyqYy1tTd59k
18MLI/annUoF08EQwXz8PmXT8pJx7+Z7kMAMDceeByWBcbNT+zPmiHnJ1zzADs4O
7TvNPYmczepJ+KWP0Q5OAAzlSon3kOLLJFbyCaTH8dhgjz55J/wvRsMxky4u/c+o
N0yZWte3nUyak2prW2JlLTsV8cytGVI2ehtiy9FWjRHL6ucezLUTAtppts+tRfkm
7xUJt3Kn3bDpmR9oImlKtxcXGw2VLxpY02WxXWFpa18btyjON27yqAqlG+ZGKc0t
+dUFVk7SxgbhlYioxkG6aKoPXv0b1jfQLCJGvmMmYHmGS+WBubZR/HtWTlnoATqg
b1W3671Yh0Z+hSUktzGkrZd6AZtsPAzzreq3KlDlnhHVVZx4ZkqDI3auD9Wu8dvh
toMxEPKVr7ecqLSoaEwOyeocWHTjdBaXRxZX/KSo9rc8DyGM9QMZ9PChzSp5q/Uf
FLaUyh5VXXG/3l9nrzILS+rCso9jGWqYtaXDApzMHBaozSaAkr+2pngP8nRisiYV
ljO8Rtn04jbIV17dm5YOxQpiM7HSm3z5GI/qqwu2dmQMXAWZga6dfWP1DY1AZbw/
C4jYdec4yGgueFEhkBImSXkXUhmszHUG+158uq5G6lkmCjuX5I6W7JtzT6EKTXul
qBhS4BM5gHvXksCVKyVT1UYSeavPzuaLdXh/0bLkKaJt7hnhCjXOTVAG7TtxUiEi
6LIbCBKacdv2LiDHJgojwf2uqo0pmK7e2vHeWyfTQj/uY8y0e8U+ZkgUQbvaLMJF
wVPlFwlOYcguTPmQMDM7JgFkZufq137KFpUmT/AOsMTg8fbqBJ8FVItOEJC5wsAU
FVhD+U6tfC0cIqULJ1pi2L/UAXQiJn9lVHaCP/T3jp7QpP3dKoNhMaUm7zWUFm9K
FryMY7oIAaEChG+jQNAd4RO2h5hKnGzvyVj4NW/LvTqvLsmV8UShJ0L/uGSvuTyA
m7+9XnBo5AJ14e8X7dtfl0LU8oqo/MVROXhTfxUjeyTDSjBX9fakCCD8nhwx/aGJ
fhkZlh+Ubm9tE9fkf1MsX0kkkv0Vp1Hw3tJeAfvQuGvC1ceU3njd/uBDPN2UmE9R
mrefaSABpPZjI+Yr708gwaTyQTQsFsGqvpV67/Blr8KWf0/klTqLtgC2Ib3Bu9/m
W4corTpoeQP8xbMYI5seoYkjjRW7AGmdBdRxoOkFe08IJKCQsbEMFDRazl5p87X6
L7NnuaZAvM8pWuQxjv5c+C0RMJQX3dDIWZ5PNOJ+QagB+Xdro5jX5DtmcS9AQXbx
KrgSNaC9WmMQSF/p2dXvWLTA67kwziWLpi92a9Wgw7vKp5L0ra/IblFymdKwRBwz
AdPyjvETd3bZrNdqYFDJ9y40qnzzd/Y9n2iuRWXknbQBz26JBJM42A1ziuknFJxX
qjzINb3LMoBhpIZxZxQxh1GK+dMc5AWe9QwrAhHPjmdXZDGO7v47h7sZKM72s5dB
e2qeT76b4qpaQYLgUI6li4F3Evgo+seObUbwsqjQ6XCTCvPJiq+lkcIn1UArj8h6
bCYBbQlpweo1dYnyAo1G50QiNfbXRk1MUl0U4ECZF2MUN4q0VoZwzqXsgFHX8toy
wIcaSc+cUXOeyoXdPY/+jpNznTuqwmff6GXD4dzLUZq76VoXcR2LfY3LDUYCl8nd
4BP91v4fXzzwy7QQ29TlMcYlZndpO3xUI0jGBFKWPPztutrnLl49rZTWcDhJwuaU
tvsGunBdVStxw5B8MkR1l7sbtxiJohwJNsAVtdzPopMzEmgqAuztqHkhwz5yxve+
5/qQtCC1FynrIau8/Jea+vxQAnX4m+g2M97tSxnjQwIk5CUbk7UrYn3qTClrTvFo
u2TeVqaFFrtChQmpjVuFQJdYvUz/nZadYIyM9hDuLSATzWZ0+abdBY9zkmldKzvl
+cvzdfAZTn1nvDtaLjfvmfe8JoNzjaYsZeWa5X5tWws/FHo8TpqGeTP1eFtox1Vf
XQyBORCcC7MJAhP3YhW2Ss6R0RfIiffdvB7lEnW5TMuX/O7eDcko6UZ2KlEtagQn
GXRM6nx12fSBwVq47weTEskPCc3nVaUZGpRDxPMjoNO3DB9fSJAPfQyF2hNThf6l
8qPIrIVnXYgZfevyeuyNFv+2wsZs8DEc6Wfm15DWpWbta8Vs9kuscFi0jzfsIiuF
S02NhyPUzKK+SpTEw1LG4AudakHRCXArAMVX9jPRfQi9P1kmaFGYg8ttYBaV7Byo
ozSscT/VHsLWYKTKFs6TadRYBiJPVoHxci08G21HRxV9TOAHYUjzJXn1FP29aIjF
cZd86yjMSlOzTnQpsDR22IlKytbvpBNu3DD0BB3kuGQJRvcB5nYFp/wvkqD4TUnk
weinsg/1C2C4VaA7RfZ9vx1fmcu2xtP6/zeb0AQUu4ftFwKGnf26HxXyiozJEBbK
tl4ZNRDBKfrhk4tb9C3H1rRIaVK5zUqlNdLyTW6yzqWHzC8TejllEMyHkHDrCM1S
fNhQpqEcAe7DXj48ReBIVtBGOLXJU7FpEJdeD6z+6v9y5n8vEj66OWmKBwOtOyng
1ez3ePD7TaiqoYPu/Lw7ncOaHU4EEWd3P8Lq9DCvlNS689+H8nmaJA7rTAtTtIwB
FGG710NUwp9jRONeo3P++QJUetW61X3bULWa07EONW6nnQzH/yptcVqxTET1Cykh
Sr+Eh5iW7PWJjZXZIVl5UVjBHQzyDlIMbhJXW7s7TfxFgNnmVCnwr9WAOk9PSND4
A/CAiIJax58vocbvMPokDwieV+fytOXqdDrBRmSAJYK5Qk9ZTjF7kTDrEsw7QTih
dE5vqyIg2j0HS/AtTb5Xox1BU02eLK4p0Y+I1XVanN4MohgPIS80TzMehGORJfF9
gXAwGTsaET3W4TJSUm6wZmNw6SQavzKe8RSkZCFsq7WuF5vdqvuto2dcQ9+Na0k6
a8W5Y1qlUJmIhmN9jaJsb5HhRVeZttnsF8Sp0CkKOTWWCI5z6TahwPXv1vCHoneo
6Zau+w9MGtoiFVBsFisnITROLT+Y7lcb9mBPRSyybOi2P0XsGkUb9QFPUXgu7D2C
EDfp1Yj1M28ogSKbsneTKNXq9r7mnsz7whoY21hXWB3rnwyduLpZ4COmi7sP1Hr5
ZQRlCEhV38KcG47P22FUGbed4KyvaFHH+CF2jwvcw5r+PCGH7H15L1wwKq9WXqis
2frIlmKq7Itq+ELEYensDDv5iIH5S7l42tUNv3Ety5JVEmM7sstmQ55VwJ+hcDE4
8hYVNw55u4SmC8+Gs9shjgOyQy9LkGoBUsoYmBCpWMytLbhINDNxd06pJxhHmN5V
2bH2FZckQaipv13N0Ry4GZJoHt5CcY3dJdgIO4RMngwVeUq4qfN4kaFyB8nx5nEI
7ElaCB2AUrcSeBUXtDPjZJGQXuPpJDmWKaF/8zAJDZwdVTL7Nx+cw+9UwBVTjVyg
iW/cayy3++i+Lw5l39kFbmY/fDePhleoJmcdAxA4gd0v8WLtqSLBXkokwYZp3/j1
kkM1vcVtFu99hSiRxwLBSNEXhKd4qLZhxCSozcT7ld0zRjxswatoLfM77KrSKtf5
27oK/XxgaQ9uUliiz7aG/JvSehOvEF2MNqCRpITO9sG5eQ46a6FU/mW7+ryEUrmd
7V+A39whwqEZgvL/E1i7bdVDdTvG7CgoUoRrgXv154LDwIQm9qoxsIbSz4H+Liaf
ThISIRHlMErlNciYh2Wysbc65tjjNWqpKKa7zzqG2TfF8R2EIZA9dqjtcm9VHntY
IyYv7CKdKSPXv79lsdTDJUkJL8LBiMbhFUCYid2P9jMkyD74UnL86v6Km34JLQGE
hlp8zjGhzjQHq3TzsUrChiWvn3tbwAHKgX0qcdbpkvmHHoD9lT5PkM6VfMdA4zq6
GoTFlD57SPCzn/VZcmNucJCYyHGXP/cs0J1O9z0xlEKXl4EcUldlX9N+shb/ZQhe
nyqssScwV4sd3QRpOcTy5IFOcE5hlSUvss4JJ+krT/gsZMMeB6Bbvtn7DPXR1C+f
+aPzSCBjFTIRK2Z7Lz4emUR6vd5+QRi8Q27Zghtqmf3DXwErCafhk1Aid/5LohP4
C29WwiCxqSq+wXGk0zpUr08Dg8CZPOFAE+uq9uRT0NsRkVq9J6oEXmur7NcN2Y0E
Msvt19dOTO/RWNxGge6gdS9whI0W8br4RN7QYPBVhOxXRYkn57ooO19f+CReIdUM
bSkvUwGl+x8F0xENGdO1GRM7Zisxvf5jzGslv4/nXB4dBFg8aYnokOYbXAzoEKbr
BCoNtp5ZqMEAei+SnmMR8J2sYrHERisaEWRE8F1TK54lHYBwNhKgPSI/ZhcgmQGv
Pycm+pv8+ziW1Wo5XXTjH7jcheI50xzpXO1Lt0ZVeuy21cdOYSgk9ICpE/VXB0tY
wNuuLrilsCXmyl0/f5R4uyjaB3OEWHMIPp/XwW8whSpn0HYghU1TRUy2VTjmtAIY
ERjsKT/NmlAxfhuYirVep2SI8jyNw5QCzXNV6F+QMhn43lcl2W6d8ybpK72pgMT9
yiP1+bRJqiH5vNtkoxlgRheu+3j8j0IrKhbNImvE0SC+T9T7QFm0pbgRk8sOQ22h
c+ZbQWLQfg/cFZqCqCGy8D4PF3qgHEgSp+ynZhGD/3RsxbyJ9T9kfWOGgjzf7l7j
pZf6iWsuEm3g6pzdb3xP/W0wXocU0C4zaD5hgPdRcvwaQi5kA0lG9ctulqPrml0H
jp0gZ56BoRGsv4PO0WgpbHfYiRLEvIEAy1rTVG6+/t/VdJAvkDRRmmmUkX9pm7ut
WiK3x448lJZCNQxm696GUslCzx+wq6Y613lWj0yP+nULI/f9fBEOi+I2kdwMnZ3t
/8aPdhg/qquAt5nwkwUT8MyZorlkYDtaMOTI9S/+t41R95NvRifITCOwg1WHgkTX
+NdTGeil5Mf90r8ZsHaeB099GlPG1REcB0UfreJN4LE6Pa/UiC88HK3N5uZMmSBA
oDOkk5TgtoMtsqcHGNmbHmvgjQwxVZxqUe6I8w2oYs3heb9KA5kYC4Z4jy9L1tob
RKdJCE4qVjM6wIiLdNEaoKIRwiNwRLAp/+kTfpIK3uke2NMLocWkLV6lUEawKVG5
CLFD7axy2BevMp6/S3NHdLhjL5Q1dmIzOzN7gz5CvDgx9XQAE8ET8NN3WWEhQ+Um
ne9zB9imu8rfDCbtHZ/TUKuYPSJ9sFIkNQAsuEaurOzbL2rFuj4XQveVwQkJXo2x
a6S1fQqeu8+Iz62P8NQ0qBV1eT9uYgbBYABNiQzNvwpaq1tAl7SoJcmtnhTn54nj
XW6+Erc4dEE1RfV/SvQXhY1ocX1HTbGFbqbkVIRDH+LWuFVxoKsMaTtHPR++ZdUw
CZ5YkMDn4KUMncqK/4o1spa/hXXBbiqyPp0IKC77GtgkRL6shq3pAgkVtBAM+4Xp
kiNPlF+p/gO2ZVlgpOXgznz1akXhS6MLSJrxkVmeTcDhngKWgpwksrHL9cBsXm1n
GwUUsyGC3vZtij29l0wAp8inLXkWXywBwU/X5OXO7+2XWj4eFquxaw0n9/eGJMJZ
yRrtN3QSLJtMayPRZNjmhICa5sJjqw8/PNZEw6nUdA9BG5Qmy/GqMUeiCL1c34GF
9SCNhSmGvNvJSbIZwSPpDgm8nVg3mxb8xRN8w4XmnM/5a2YGP2FlFV7xgJMLrjsQ
eAHWINzoGKL3EsWzF/83VhNo+69mjyhRy8+Tu5J2JYU/AcyOJF/M+y9eCevYkAv7
B8XvsXAJH7qI+nskw242bwQDejNFPSmG4A7fMfDg8Eqa+b3K63WdjrmgDjtQXB+M
I/A3uNZ1eTtNncKoppB9FuPvwQ9uHXhg1rZewikqM9gidn5jET8QDtyCs9c14TLV
2VNsXNIOSKG8iL1yTWK00sXG8SNMlsoT/x+n6tkx+c6jlI2I71xgfUwNHFGNkBe7
Y3gzBukUbrU8ne9RRFs30JYIFiKbjjapWuByGCvi0+Tm+rbs5SRMI13fyU6l/sEz
W3sKBig0yNxR7sjUZZJVjKY0kO4EuaCZDU07hB4KR1zL88+037unaxz3x85djrLl
dlZ9eiNc0tAoStK0diMr0CNwXhjw4EZzLQ4Dl7kFrtsxpnMk+cX/HsnvBSMKQdu0
4zN9YYejBHU3Rs602c2hBGUu9yXZM0VTveeCvwoS4fJ8zRNtsY0UjrEKAFOcc17g
pDV1iktj83ubeeF/3dECcSGPXwbxOBi2GHC+sp1yb0Zr+/xom7a0hQK0bOk/fZbb
dSb36L5WFREMtRwqXfhkgQkdsRvEtzUnDnOgwdDlYZcCJjmX4r8SJ4t+Y+VUC5iQ
5pdh/VWDbTLlmcm0NaJKkP4QJfFKsHaoW/EJ1RySHzptXFWz6O6Cttfr+XPxzm2c
bAT27ixvFkAYN0+MQS/ZczEMsF9LIWv2K2LMQN/gNJNJVgg6B5nkEeEB3FmGN7dz
J9szMUz5DAIV+dQ8gFjYAYiyJi1Dewc/cI35OipOWjVUNRkk0VTx/MNlm4qS5TCL
yJx+kyEMW6ZEjxcm2w11JLHYRlaveBfXuHr0+uxdBj0TVquPCWARsBQGP01eUY6Y
jqN7nOURjcyJtZWlKW4n270OSP/ECy3SIL3KMm08pkdtCbQwns8FlpCLnS1/NRMW
XEAWbcwoPsyNEswbQ2eU6PwtMa0vq00CQrE8+vLbr2CK4MkoiEmJro8FdmN0VzW3
eUYoaAve+ckHmFUXKASUQ4g9dmSgfOSpnuAgjOc6m8F3Eg91KwUfP6ZCDBiNB5uu
nI+uTjOe54zLjII9wktM25s4hNl6cXL2Y/yEK+EVmcwyucHtRN7ItTcda5MEB+6W
zjnHaObM8OepcWELfgj06sg+qhiNKIY6HpubT6NpvTIdV2OmlCvUp1OWatDH298t
2GEu/LgwU7Wj2sqxdnyI9oNOc/i+gvM49wbGFl4AkWMNdg/jx7vt+fo7PS+PDTzt
e/Zp0Ivna1SIODl62VBkBLXqHD9ijZj+m9JB40ATu7faao229K/E+oXvSvFUCXFs
s0TEGP7XCHPeBmN+ax4QP2CyKfUDjYLwmZvO3CZJ1Kc7h3Kw1tljJY2zv/kEI12s
Z/TYKCECke5/vhD7+JUSdRfxaKG220bOmzfnSL9TZzB6K8uOZbWUGbN9S9s0jDq3
i6c6UmETIAkO1YIn3BnIpP8hIg7cc933wd1x23SPOUpyzEn9PxlXotjql9mP2Vit
5r29c8vg99wltXqvRqiuz41avR92bkrSMZ4y0o49txsKT0Dx4LI6zK00+80fOlMU
M/mw+3hl/tQptnDxfp9VR0Pl82vfcfo33ULPFPWKHfhE0Qq90X3+3uuSg+zNgddM
JjyOeNtPzH1lyAIKzoMqFpVVF8gOEGa0O6vTJzY0noM5liIAnWDUTgchazYV0wdb
kk0ntYTGw8CGDVWzMxA6wKGwl5KKrn2T6LXyKmQCHfyu5LZgEeRUEchsDrzhnJz4
cBoLN3lThBXmN355QULBviKMx0/TxSK/+550rQpL/CCmZDD/mlMRq6sqrJ+7mSHI
h5ddRe2253G1srnHAeP8rJtAFJA5wJVCyU9XUsg1r4W6fcfRPkpw3skPSQUCq2UZ
ICpF7UWklWtK+vj0xP/xGf36Ioru+WLekcfK+FNtCM54rCh7Owsd2uoVJMzooCMX
WuN5kPie8VglAJZmWAJ9yh949y/tu+m41nuehf5U5STMkDJm2wYwJgPnX7eNlY12
LASj9vqce+uMQfPlMfClBx0deR9gEM2fqMZ/QUpKLl8zVY5LSTukcdZ1Clcrq5ay
Y6Q+7zKAVQOt9INbotFafDC2f5NqQZEkN4gHUV7Fhdf2TagrVwsyNqaNLWmge1yO
ZqPWovCa4OoK7svrt093IlKKdkWKpx0bIRQQsZokPMzbgWcI+QxcwuFtop1Pzn2G
sp8c4A9uPoOGkOKJcnlshqPcYvnfKZn5BhRELhhZSiI5j/np+QtO2ykn4c+Dzwya
o9MfynzyGqVDk1D1JucjLEXqmvlwLq6Yal7cCP4e/9Wb9od8SNM+jFYqeetYDEB9
GiWANmWuCc5yXfSBc7YgFaUjZWLOrfTxs7PuNiiaHPSNGGg3MA1KgBsYfyxU2WMz
eFfufifN91aKDmS4/gq653zCWrwZXrnbg5/joktuQRCIHa7DguL1/vhgPN5gO6cj
AuQzuh65ePjyJ0ehX7UOeIHtFdpIHBQPSVRJ+EgM38Ih6iYLdJT7cU0pNV6sYrT/
QebeCqzcpD5+EuP5o11xs2YmO4PQ8fX5AQRO5Cj8QoygL61vfhnRzLDzUfhkwtDJ
McOweSf9KTjCsXCQTCn3cbClq4jMfXaXxf0YRS/Dxx+EFNOyxIVoA9abPQvOvHOA
QYPvdrl3QUAL94Hg9sb1+386KpFkSA3zg/+vLP4ncFWXazmyiHmV+0kKWtobh06K
z5rDWGxtO0wFmIV9IRIOZc4DBW12y4sSkhn1H/5X8G1FEao+IuY5BW3zkrCeVFyJ
yLUPoWi/T6cPIUPx6NNVKcD4lCHDTC17740Mu9c0kxWtf+L9+NPIewWOTdK0HJIA
BRMiCmCz824TVD0XfbcyZ9QqM7ho6SKYMOQ6r8ivd6TPn8Ug4BJFwIRZd0mNNWM7
5CGogKeXWipTaUq3P3kYuMOdnsa48W1CT2QX1kdukMpS6alZ3qWlNYntsqH7uMua
Z5l2cZMXMFE+sxqkVX3Z2y9lNHj5zvWwbVZ9YCsP60OEjjqSwMZLBzDpSKhdUg1W
gmiJubHjbDy0YG/Mle9U+wfHEBbjLoRjUEl+RFZ4ECc6kzc5BgyfBfrB9MKqCXhI
5gjSpCBMtmJ4XLyQXPgeAGl3+F90H704f0TaxMBbqEIKHZXZpgxGuET7XsOxS6OS
PNlo0KAepsToRgKqLZafotteLnmxfm39HPFvoyjXrP8ESvJUkzT+gI8AmK9u8Uuf
193n+D0C5lIyHnXJZOuzKPq7hpGFURiV9r24JrcUjuOOUfi5CkiUnAaWJtdo26ue
WtJDUy3/MZFBnNkTJMCuPcGp8TCCZC8KZuGct39npQQj7jizOiY3+kOe13niuUGr
TikHQZYEF6zhCXPMftJ23RMHvvbQe96BvEsl9bu9i7sg1tUWin5V8eozuISbNpqN
ADdx15yp3dzkLU63hTxorNOS/nMZOUIZ5vKWcGvbAts4YGAZyxhpEA7z+kUyAWiv
Pcvk0R59sfWDyZ4Zsl1hNjWKuKUr7iq+MUFa/HU6KHtc3bW/czBVbMCCCyiy+Kbd
CmdPeIbPBKi8roC1N4iW45ssoQPldeyx1R/nmrzalS1+OLHm/4IE1+6GYXO7BjrW
U/08UL1yyhSQAERauoyq3ca9ZLXwYjmB+F03+jNQL8sU7oFromGcThW+d9jH+i+O
pTQAYyx1Ih2HuNQ0wUi2/VPdu761rLyOd/JY3wWiSmA9f8UfMgfWyyqZkKBRxSB4
OvDmVU3IozDo2OyIxhLuezO/ewbwNSdmW4fo5mhiFUX0RuYW0e67AxBZ78R4JR9W
0FiMXYh587F0lSWVp0FjKYoAtwHVIsLT4Ll8jr0igTnyAN07QzA9HuEzR/LnLcQn
WdlbucvP0Fit0HGTZW8D8ApYMzH9bOwA7ZgPksnVvNnPaFraIPUbwZOhkDnhF8Mo
ILsFpXuI5fpyd7K1di+8BYK72eZvcZ1Isj5sooGwac9dH16G4Y4WSaGFQDXHp0jF
PWCjiv3qeJq77MOTEuNi/0/JXZ55NMB0OPsaOK7LvSgFEtG5N+DmklEfHOg+k+lL
46O20K5oWU7NZFFeSgY3HqjXj0do7jWZeuTJonH/ZV7QnEQDgExmbIMIF72Djiv1
osDUtDtQ1wA9fTGCJeu7ZyrRbr8T1eGNpZEcE/L4o1/tl9TUKHngdh1gD5VSks1F
+u74eGafjccuY/HNIVrqI/Z/elOwFksOfPQd8VtTbG9UtqZijv6rz/J32mtWHnUl
nc9saY4/b+mwg0OF/4Bdhs9x5k++gbDQlscxvZ2PyYGsbRsQ360WUXx/CanYGa7T
UAhp3l+EQdnpnN11md/gjl5cay8yZOXAHS4CA0m7miUCSg1www6fwX3YD0Sli2H4
hoxsuvkoFhV/3OELVQZWpvXDT8Cgb5ci87Ll4Z16lPFtBklaDbe1askS7hjRSP/9
RpaUU66T+DO7Z/XIgBA0Z0/PX5YjVDMCSHFkXjBDTsle0Yz9ewGhM+az7RVp5e5G
NeHPYtorsVDjaPZSL1fSLzjOba2M1Szd1N9ekhvB0f3KYz7PzN1R36bMAeNYbJTB
M5B6+KZfjMgzY+Ea3FQ3S8Y2O/tFXmve0yczJx9a/TQP4WzndBrNCbFIj4vQ1s35
yBPu9wafmcMUseEXqQjics3Ii2ySNDTngZKiosALJChLuaMRRd9Rh8JpltmtnONq
zLgVAm8qHzfmtAaE0+SlrT/LAf+igRuWneOeaeXDbN0tLoahDJDGH1yxgUf2FiHs
5blhnFkzUifN6Lz5CmiLQtOcZgDYv2eTc199r/C7+c4Gp1W8SHXhJMKQAUnPuvA3
f3OpzsfT/sI4WsZ0hD0Mz4+alHvYvo7c1qbchSg+QQkP1fpYqXcYCyc4DVYrKkBt
0b+CNko9W6/AEROjaUrgtz8VWpTnN+2wCqhMV4vEU5rYb9ZO1AN0wX/ymogkAbE4
vCUWP7P9g8Foiwcc00WrxZjAeStnfd32tXf8AO5dk+wOHM5SIYz6AWE2sS15hQWb
RlVhSIEkd5o0ApUygaVm3uGUKgxRgQ5fy+5aw5W2yH4NxeTSjiZ8is/w1Jg68GEn
43SyoOS2bI3crzg9D1mUTYKRGZ6BNOUNgLzFiKV4EDLBmU+tIE3aRguqa67diyXz
IuJWJZkasHrA0zaRV3HvoFIKZB1tsvt21Okj/xJw0CydMsHNgoO265Gx0obwr7pD
RJ6HEw7GuLjuEd95yXUxPuvSLY0eAdEvX3haSjKl4KjAQ7rYLgia1nnTMbdfMoKT
grpHFBCCwX6RAAlzbRpIb1toWKAhqPNPW4tlKy7bth7Q4XGRZGLD58SEWl/yOcHc
L5P5/x20SzGHhZthSekqtttV+epvM20KUiBTuJBCXvqm0LYwa1GE7et7grjp/3YK
IaNToIJV0x2v9ctejyNcavgzD0YmOGmqCa53SxSOeNGuKEVo8TwysCPdXmcLDe0j
Coeb8vOxCMX8mTRdloiiI3G41liNi50axgYcs4oG3VYsIR5iZnQc/SRrxIDWc4+f
AC33LIorHL06NBUls7pkYE9viMkp5oInyAq2Sd2+CqOb1m7N2ukhFKRfxkS8oSCe
iO9sG/nK+NMdqs6NlODwv1COB07yOq11YBtdtvgSR5agwjyruTbLi+oek6Ew4zo4
f8NYPvCLn7XJMAGUjs892zap2/MIAJWiSUcybQFNoKxQu5AUE+zCuVqbZHX+q4v/
ExABEgQ8I61VD8yaWUD4lKP+HQE/+kCGBnGaTVl3OYgbVGieh2uzSuYMuarczIFs
9TH/H3zULJGP3+y1defTzXfH9voztJPeu5wR7kQfwmewe0YNeG/o9r5X/7cGP7Dx
lUwj3ce82YNfyA5r1kF6L0x0yXdS2dzMlsJK/3lOBxeRzS0RiS0tpXkJTKGxFUt+
ShYeRxBrp3MN+Vb/6YVogZHza1GR53xznnzoI/OEEdYOJATeS4jPOnii6T+izEHQ
jkgZdMmQyE5n95Q4gZi8jpUU0ruEU9rV8p/6YzPpa6WZSwSXWRw5Pn0JeX/UmMIm
rpg7IUonGzzRCljMie04gJd24WNqzuUYeKYlkicHFcxGfq9G2hXsd3KBDN0QWZuy
nMShRXCTK5tsFb417oAiftwO6nNjs3DFWu6rYj+Kk6Mmduz1jiRG7tQvD7PCDL1A
f5l2A1ICJ57zS0XVrQCUo00cTfmP5x9foi8QxtD+c8buuepTqjvJVLq8EOZLAHl5
E54IqbYJ39KREtD8/pzp8EeiKPWft+Wu97VN3v9QfrsIJkLxqsITUjgiJ4RpSZfd
D04aUPYMowd2XZyGKcPP3OhBlVQDRb1kdta6NGn2/5vXi9WP2QBxnxuGg7CAs6hT
vKGizBLWbu1eK4FyXErVqn0M5DpT/VXTbfsr+Q9yZy48A/GemAXnoqScT9twUvP4
4wYNxG++8xV1h7LIntq5kPyFFw8ldfoSQZ4VFIdEw/aUnKqVH4BgIw7ilXU8KklB
PILBkiW1OBaNsbL8f/OxGv+PR0uKlGGsGv9Rbl8gH+QJ+r1U+AS3XIIseoUxE+JG
5xHJ7vnFIADNfVOkcuSfDo4eiyZG+u53yjXUsZlgWqXbV19y6p8Q1+aw0h/LDA0D
MbREx/kPi7e2TVb+t4h8RRkiCHwZyUPwrDH3OhgYld32D0+2qQWfCdAykb8oyUqW
I0gFY0N0gnxzEOfTkPxtq2YR/2f4dpBJ6vWZcLzOKnYqfL6FX5ECOUK+t9Olp1sN
VDEhN1JptoYRtn8+ok09djP9GHaDg8omPc/AYnZP4sZZiXXbFLs5S3Nq6n8GWbHG
Cms6NbkAu/LXDI2yYG1BfBOF0QMV3pv7zRxwlYi8DQV3ZMBXBdQJQYOGOrnB32Td
aufihm9A6KMSFRHNjxH42ijqFsLNDNCLVHX6//+IPt/X48m0fBTVoBAQFXeg1sAp
acGM6x9IOlUce6ZkTpo/qwaXxFJUziiXZ9kepfqJ4G7Q4rDdpv0Y6JKo8aVVO/Jg
HnC2GzrU62GezluLo3s1DPI1uDwT4p5NAW+8AOhI4qbLsA5os32UTIGcmX1p3nZv
3jVXWZ10A1L70MWdrNoB2BflLKxAIl9zJEevf23Bylk6t8ZNYDZM2PUh7oACL+pV
gOakAfuPXAMoGu1PA7IIgkoUZRcaGvLnRaZNyXVbVFSt6BYDMyFg26Tj0IYkPbSq
ujpcve4S077KaAdrzky5UchEf4Up5f+ritgmOlZMhwtWp6BU7VzqOW/WRQ84+NyR
L7/5cjp/l7Zjml16tAD14NBb7yu99SriL30vnwkz4WWWIgNRO7ETCw3XzI041/Fd
BGp1jOpSGRxBDwF6gbcDzURidPNoVw0TdNNRPpoQag88Akyn8SrTzihknu7CTmPS
9qJN8jPkX6tNyOLbiiOqTruWW3Tv1tUqdGI84iFiEGuDKyNwV3bTWrTSDT7WelCx
NvIW0SWgIMke1XY0/0b3TTCtzDY2Gd8XVhOAjKC3s0W7rjTnurSfJQ6hmcS1XmNs
n7tOgWWeLiCkACjA7JRB9kLDqoZ47ZPVbUtGIXpmlIi5RHy7R4BX15xZULD/SSJk
KgNmaPJEfliHFfgxI+Jb7XE1NQNsBDe5FIjeLK+D5ArdSnslbiBv+/cq05YMx+B5
Q3Ts+QAJlhops/6Q+8SNgXEZL5iVC27XQvgUO73U0pfEfQyBsoAX59qjd6QR8/VT
sfUWeE5L15AA92BUDNT2e1uGctmjuyzfr3YfGboUgNfqSwm3MjSPnv3EVkHhV+Qw
n5No4jALz48PGDIlTjk00om5W0ivWCtn+i+NpyS2pSaHeaT6g40uR2OskwCXoyp3
XHupBTbdKKkc3InGi2916jvDl3OP84qzfSLM7bV+PjafFl99yP+5BcA9VzE1eY0h
WZ22JC7qUvS98p2i8CLbFn9fGpHWTZapczUDLGwWok9bGleHooC/n2mVOezdYdYQ
11+00ZRgFlHQU8W+DKs2VSVKLjZD7vPGby1vduYzk0sGI3L5+5ynatsetRp3x3Js
xqNz122fHCIxiI4D9rn1CkWWglbaL4Ke74ZFf2qoKlikrL6Ga+kBz4BuIlofXTUp
+JGKcSqUxa23nPK8aGwfYYOkc4zDA2yW8VfkWfWKxGP6qolAsM6WkcDyLvM28t/Q
kR3J7ZuowTs8gAavbIDqW1gvU+GeadiS5X9r3y6nT6mYmS7VIpxVStOCWkhI5oiy
zxKyvuHp7eFn+HIJd+PzCz5erALYX+LgUbHwK89jLfjb73nvwiSWWonmryJZdRkp
1rVLYT3ZcLsGZzLosX+fMJZzGY3jJZq5k2ODEO3sBjy91YpJQI/LImHQnjlQr92X
oCL1kfvz9BtBbChpRXA8ShCQnEsGi+LRwPzj2bKEmzybhP9qbVhM0TmwHVkb3yNV
CcdKXrWEXxW4daZofaQyAMuuTfCLPkqpvkkCjfdhKj51J9ILthE805F2U2guvp5N
74tVQubc7JsngjPRsnisfCPepHSN36YAn9YAutrDHLpUmf3OWW2dvNd7igrZwjSO
P0DP3DNyaS8oQDCsOqOz7XTX9lDGyf1Gr3VlYPvcOpOR30zgFzyr2alUmtXFPP9t
qGvPPSvdIf7ezPBBsRfZ+xoQuzkg28g5v5mHbsFOsiHBDuzwO+f6nlva17RHAap8
7B6lBAs30Xa+ybV1iwJGOGDnR84HrWQS4AecWd6uqgBjpePL9cI6gEp9X/FmIJWk
Rfv96Uy45VWo5MPLN6GukZ5wGxwUx6IbBcn6TLCigICidHW+14OSeKJ0h4MZtNeV
9y8zitW4vlQ8LEE4CYjjuYLOK6rFiIbJ2/ZGOzKDfix1MLNWmkRFmqmZ6geCN/t5
jB66JWUk9R9E2y2je0ySDsq+H0XeBPAUX5emrBhbFsht8tEgzAYrgrKDthKmks/9
8/XEbBpiZ7CH4+0TlYjff9196fe7Yy0bqPwKXzM2rkKW0r28JN8NVk04TX8eATbW
vjCUjKJo8GpqPl7+g//3SM3MDKad4Qn2+d8ZQtXTVoxXyKM0Iwq4SMZqrgyfRCH4
zl5mTM1dCzrcLOsIqChQItVOwIywjacfIe8kxWJG6AqNNEhDQ4yl/Qpqy6rwKVfb
YfoV8+TGBjVq8aEYP1J8LgZcxcrZLs+xJkixVYalHSW5Qf6Nnn74k4MYcPxssBCf
SvNW1Px/mcamr05V5MtKl0bOgXK2DNOC8yqtqdzXZIuMqCNPEK9AYbQGtiVk0XVC
Z3tefa+OHjf5Uv4MApuIMDsWxCpKrhhV7pkmLiU8cJAK8DIQHF7qQDHTdiRpFXlX
0gu64YhmE+ZtR+sGM2DEfQXuZ6Mu9EigfNX8Gmq+na9YAziCPlE0bhc9/NHnCepP
866psVubFCXM0V+p4upWkh+97zbjRCXoxVcybs+oHqYxqtBQTnsUP+CgmtkWRIH1
p4TfzCAvsOCAQWwNkMOynTfpwuD/zXqf0Jgjp1arnY420uc12jBkYDCH6VL6PUhz
DQkeQePGI6OewkAhGxE1kP+0p6p5YZ0adXzhDrlZ+H8OgFdewJ6jkoa94HnVsGtq
h9Hg11MMohnew+hwwVi4QIJNavDBD93Omz3cG5OXmaKsp/fr51gdXM/2hOUHW824
GPT1DGnaHUm5IQj2GJ3j8rK7xgrsoCm8vLFJKWvjVRkHWhrDroqMZX9L/0lrsITk
3DWFHT/iiz0EB8cWA7SYqoJYM/aTDeGF4nzmf1dgxkDpLNddDwExI8SGEAOnEhVr
3s9tc5J4ALvy9qqgaRpR/xi5tT0CQ7JREPcikepWCC4OA5U4uxYn94tVG+Yq181O
/E2sOBIMFQ1MlvKy2vGCrj202GzB1f7ZZLVysZHK7k3D68FXtuJ3LpDD9ZmI+SDl
33kbTQkawY2zhkSQwBLLNJnopmG9J4aga88WSeiGfKE2Q3Sx1/mJUFOKo8/63XGD
l9+50wQQPpxTyjpRXrlOVu8ZcFYmIDdvHmMZUfBgpyNKKviwjTjpbhSTj15gpio6
+yiCuf5SORtkE9wgrPGaKKo2qFHM/BT8kPO1VdFOZ1z67Xgdk7wq6hQSbZqU/FVc
qR/Dkh5VaXNKe8R2PfVE3S85PlJ/B1/0BRTw7FW/AJfj8eLB18c9zwpyxUd0qY97
CT9r21h1EO069gUoJWj9TzOJKjRP3/mR/PnDtmhWwjB/dmlGpjC/Lm9vIdwiiqPP
fLexWkJTmpFsrZSM3CQKo73WmhlWpG8dNTVeYNs1Y42IjANbD/vdymxqbZpPbR0z
wHR27ucR3rdFnizvnrbzVLVYXbGsJYLx0Nnp9krdQaJ9TioRYN8enrQ3nIWSp7Hl
Fj+YCt0DQ9oSnfkEy/wJInQacmvg+Q5AfUo6bW7TGm/lvOB1M+JPvNARFSzHGLzZ
VcOoHwvdCjgWS6CH1RUFWuJVyeGeUieufI6eUihcaOnIeOMwH2eWi8vhcALmEoJZ
oigOvbhZ+0gOKQmKOPrK6BvWuFL8Pu82VisCDNczJgJF1luKPXS9lr48g5uis+uZ
/fTa5nr6o2ZgIgK+SheEYHq6znle6+IPKu/J3GNSSsfEXwtX5R9mGZ1J4siSeL02
7bXMVeSRqCPJ+IA3uzlG7Vchs/D4a6euHPBt/ygN5bCunAebnzgvMURkabJXm1yC
o1glnmlVCslZaim6V62v+RIjmAMRWKOqe24F6NIxupeCMNOlaIlkreYdY8xosJ0L
pYdPhHVGu0/ZK6BWq6wThjIl30AYs+Zd1ZPs4oYm7zeI68YqWhR3nIULA2Cwa7Wx
4sbHBTpsENRYjsBJ7XS0ZVmo4ObTmw7rUuEAcMy/bhkq3R93LYFqRV4CrhVGQeZd
uO9myk1RfcJF6jbCJsqyYm9uWMl31bhgr2wZ+yju0lpEfMbUw4KihacWDU+l2nh/
eHphiHwCyXjN4gDPK7fnNGx/4txMV8F2s2fPsVLnJQ51CLrv7U5Y6fQ/XvFya2LQ
kJEdMYpcnq+ChsBeKtxVIvF4PIzzKGkKschpe0ZJgOwzGlST75FP+K02Zt5dH0UC
znqRW5bH/Rx1i6bVSPIiCBnEhDk0f/0N+Hk2ytEQquRkS3mzCuqIhww5nkdjkLNw
CFCq1SfcpS9dxrTvD+ohlR8juh4GkKsfwJ90LNwJnP3hgxR5Ed0FivH3GjxN795V
X+vJrGhjtZ6N1lSgEFaV+SP7Qha7oA8dIEhpee6JLFlexJQE/3lwu/eplFxsukSD
9UfXgD+Q3gMYafjyR8JcxJO0tr7ISiszUfbft59bCJFqiis2BUcfuBogqlDHb/8Y
D4FT5NSo9GO/L22c5d70mAlwtzcplYqgewSCYLF5rgj37Fv7ibSrwlxB+5qrDoUu
SlLanZQ0hf4ooP3VZ3cDemQuD/HrJSp6UB8DMKGJPOCbRDg/m2x0a8AKYyFlWSAQ
v6IbTtQm6yWfz+xZHrYMXmNbwFHM11WQ8el54Eh+MRVjVJ8KmV4c8cz8j4hx+vaN
oHv3G4ZDKadLdgM2x4cZHJdedoRANyq1VuI03XFFPikqwHDDwNJChQBcUV6viAED
+H/k4QMVTjsfuMIq2DkQrbJGDKBxG1NRlPmBBUMqjNjXp6vGy4DtQ7ON5GFzhWsZ
bRolyeBF1Bxe6dA4JmFvl/V90Q2Q/Wrak5pUorySjPtDMKSuS+E3dwHN1AHTOejT
X1rZi8UrhVUcdlvc+lzX0sgO2d458W1T0k2aIjj93oa6cVTzR9eZNChGkL2oCIsm
tofvx63gLH9cC7wZtT5lJpi93XxT24e647yw6kneXLgdBykCqlDixefAFB9AfQp+
xmF7uY8xy3UOSzFg6ZVvrbVBzlclkRBDSzbUtU73gy7I9YmhbdMm2q1vX5kxbD76
jR/fgSqaniSzNnPSgLlpxQE8jk+y/Jv5YR5+M3p5se1fZ66qmCNk9TSlg2PO2SBa
+76mpHC/6i5hKDX7FZT/a1oITPMp8umeRnYks2h8xGtLLKclGHlIHXlZXIVadJkK
8tNMlpvtA/noPl+XOiMZvrCGXj8UeS8qpNyA4WZn6h/Gjg7QRZJHtg9CnVrUIqxB
05bf54fLuqYGtgOG+x5rcKmlOgJHcvHg5e6so7Y4yOvOYoG2Kh14ucAEdevAiSmd
wawtlWVaDib4Xd1qYrfmR+5eXA4ngIVoI0xujqb9YUz4tTI3RYqJZGQtm1Kdclqt
uUr/Ghf0XL3xqDMduvLYh2YTpJaS4x5UBgUFGTc6MRl+Q8GxbkHZCalr37LStK9V
mfXj2a1MBcMFUBlo7f21ByWXOXdJqMZiGkqIXg5VrlDF7HXVl1zm+324iZFCLvvo
jRKS3gIXb+JEGnnaeFy5QXDwLNda6HgRmHUfgROxN4d4Q1DbXlLDGFOAemTi0pl4
2Cy1Dj7bHFIL8wZLFm5mzkFKeloJCQ8W6wOKZkSkbTKhesf2kAzgd+I04EwCzgYe
6p+zMU3zzaAm4G5LqB6vm83rq7bUafzggLgd+RD7M4nwo+Y+OxaWVakFK/Bo0ueP
+2lznHlSEubiYnqIZ+uOyUJ1F3PxuEH4NmCXLX+coUneiRaPxLqeVNpbBQjaSKcX
EVLIaTE6CpbKjmKYzABvqjz1rNg/DZCEzVxbLjLjB6/NnWVQ4zqy+/4mWrp5h8Hn
xjrOMox4JiHieD/Af0uUwtleoW9bAkWNpj2fplhCDeB6Oj7Ozfv38EqCVsBLf/CN
HJhrEVEn/k2g4YPPZjGGDTq2Z+dH4xpRfBwXDINk+afmanEm4QXKsjUpT8o5wMkW
XXBXRzE3/Fr3v3cWID2EpPqH1gomnsp2UScR7U1fyBYaf32IcdFBgO/EsrZGTbrw
uys686jLN80orK2NuQO4QzrHFBQN3kLd3tqn1ExCQvieGlMdM+NbN4elQMXk2F8j
0zVFVJgry3jTAlkgTo0YQV41eA9osuK0xowuhednDa+ltMGO4fd7y5FR+1hKg9nZ
KHgRkljSRVpxvF+kW+ZvJaW0LNth03y2NxnrQ+3kLKuJQt57vXiAQab6yNBr9+Ed
xJzDk9F2Y2qsPdUNyF44UiAb6NLDNxG+sw//v+rgOUvEAe+ahASRghga/YE/kdJ7
kXoFvPBVtzEBxk7T9L8fmbSe7DZJKtj1eRfusEFQy/u2gI2xJHuvTUorC9pASyuC
n2Eu/oj/tPqJOBfkE9SzkRV3mBFBSVjkyofiMvC74oyS2LNinr3XamEITiW+pbFZ
WWTHwIS8GtlvFrwC5xZKj4TgvaRS2NqzBxguRb+vj28D7jEmVhy7zDGPTKnjd84V
iKaIk0CDE4hpT+uenB6KnIs3xmhfX3YRsEqOPyBka2hgpuXXSw9+jLxY7T425pp3
9KWoX9GC4LSl6gGyS11XTpEPARKZ1/OaRnzLtTmIMO9YStJxpWDvZx7uQEVuQlCM
H/+xNvp8CKnl8m8BOjIIPoZDHu81zhOnd5jEgzdxHhCepmgW9ZDsCj/pstPIqY4O
vOBRiVN3L/C1mNjczgKEW46YZCMIGUXgbADwrhqYM6ECzP3uiCG/AjtxiEX6EbuE
k9MKunvbiNP3wjAJsTOJ2MVXcloLpeubypBoLh6g5FAtm40CAzA0i0kRyCfZl7Nz
JnZi5Ycc6jZOX4E3xc7AMyuM33niQ6QAO7O646oVWMTntTqWN7IuyaIbgWt+1Pv2
kXH3JsM23dQTVz8XE1mMgEVBhatAPzRc2sHlxSZMdvz9WaGu2GhYPoQXZVsUioP/
K8tkjqmqqLk3ZAU4cki0fsknT0Hwoq8t0A5EUvkPOY2CJH7VLQv3cqux+Qaz99Mo
NdlBLfeNJ0WQhN75NFclzK2Ig1xDsLihujQ2bdeXMhUJOr3ONc8ls2VCrrHb41Qe
zBIqSqZfMzySNGDBmgzzXqFSBA2orjy+eRwgK6JE6YXoKNrq8Tz7rfIbDCzQWY5S
vQrFx65gHLlWWnkim8/o6vEmtPJOBDDrc9jt/uGXeBXidFZtwwbOn40PfbQicWxu
WVHjx6vrbzISfJ9RQ8vhWxIFrGJmwmxtrsSfvKeD+lmxJWl9eF9YT1JpTh6Gazkx
1m1rHh7zrRnXjIJnzqgryFQ6kmHCQwVYDPEMCFF5SQbdkJe4ocgZmsnvOqzA2FJy
LytxZ05cdy0NN8mrqTxeq89IWjOMrrw7Vg0LBpddGwdATFGKsehtS4mBratQ8f3K
XIAYMBVyuoexIRhPBeSzw5sWO4TuYt/2i1vV32nLXrZxg4zSebekuE9UcSJGfubG
l0TO41F1b90cvb4PTBpyZChs0u3ux8eVlTE1LNC//3XzcFiFEeY08GjN6+Ru3AKD
eSJQCdj72JqZpiFsWKy+0kLJlMfM0/JzIV5VcHvDEQ1V7df14wgfuiGtl5EY3SNS
LEUWzJ+39EoQYf/o+chBbMuaEBPWHvaFnnBSBcRMt8655JqlPedsfdLfYebCqjyt
jWbrtmHuZo1vs1E6l3WBuL4PKIyrS2Qt+p27mFXssdfHkhkwkXgWhdfeXBQrcx/3
w1hSP01wEP8Bo8aJe6h6I17U45kFabn6UYdT/PB/Fzj5bO+6aaKlDULC07gRQUIZ
L7iAG37JqXv+pNA4sZ3aaUiKbCq+C7AVb8EpxVIEWYteX8Q5u8pAd7GDFqVpZLPQ
Ne1CoxS/rlfTxv3q2DQ7qdcyrztGK6Aqnbk0XvWaNd1FtU5ZpBwD/hHqFE5AimdA
vdUmsRQzOZUBGpktEj7RlLWNxrJNpVrX4sdaLwtTmOdORZutWRahst3nqQP3/5sa
BINGRBuCTxmlxapPQFGNPubdO86u83Ntd7HCA8Iai6dEn2F4cLC5yUvMZUCXhN8c
fbuVIVu1M8aAOeL+2RKRo+CXWqxJe6OxoTm9ivaFyBsw9IE9kQz0FY+NlsoozEwE
bmHsqr38qLoDIqeMevGfz+2mIf9qJs2hOhI09HRE+qIqhHz/aV2jOPOmctW6ehc1
B3DT/4nGcldggjAc/xNrQT1X5oyPe/ejAxSIKqHCqwp5XS8SsDGiB4hrWfFNDCIs
4KNvMK7dQ2FKtD4kyUuBuICC99lsAUo8R07v3hy903+MKm8jyxuQKW8T60iiKW7W
m50IVgdKuTczW0ydo9T6u6jQrztQND5M8PnjAVa2WecskMKd/oIoj+dizef+f7/I
CnSo1LPWOcKcjM/UiHccLD9TTLA1q0vhS+BOKTqaLVAjqVKDhR8e3Xa5e5br69hk
anqsngEVhOKSCNRNJ9dj6Ifs395IIR+hFGJaraVoQlrmV8SA0ijIamz+JOeO71P1
jmIzHxe/6kQ2NvpHlFVixiqK+4Xom1cUNm11yamd/Ik0daGtJGzkiNEm2qE1QYno
dC0Kyg6JLDO9kLt6hMek+aiKRqDaVCAeuRdRLtUCj0EYGGcUf9FmhOqf13H47UKE
UxPVOdoKZo7ZsB3Um9OfFvwteawKr3ZScVcJozFmUCsyinw/XMU8R3ZOn2iLBq0g
IdQ9IirI8ekGBxrPC3wh9tQyOaOwEZAzWAIrv6NCEf46L94N9GtjvMgfDdqjBx37
bqONFrlYPxPTrZreIvh6MMy3QJH9vMhkVfywseLlWu3/7R9h1/6Nb9GciQ29QfQ3
S3audJV/notzDECITbabxWeq7CkkHxjZsw0Dnvsu9nNTx/jjyTeN2fA+Tl4frq/4
P9xribW8KCsIe8TjIvf34ICe7tKhQSL0v+8lIHBXc64wajfeeuK25biU5nxHJ+Oz
xFZ/6rAWQZadRqZpnZYhTQdWEUjflFTNzDSwrDjivRvR1uCNW75IZCMUQu0q1fhN
Aepz8VjGonBuLq+7lZ+zkCNkor0FEMzkiVsLxT71YzCvW2VHgrIj6NyQFx8+BVqU
t4e7KlC8z5G/FjjfORBZ8FRSEbSC2f7rBuoM+X2ye/L4gFKUV7H9VApGSFassK/O
gTMzp5ZnhtuTLQZ510fC+CfYFzj1stBd70R6Inzb4jdS4jp3LL6MCYJzulTBAVfu
IYjOb75D1S15aAonrgyVJU8ky/SSAs81C+guY6h09RNzhbv/p2Axa8vbRIawWtk8
ft0a3EkiVLc0QN/TKWjoRnQiklMi4UcWolA91A7ZSSX0LDyqrqfpTicj2l90qdnf
lOENMtnvLUG36nD7evI0z22BKabv3Y8Yx/zAs8bxse/6/h+XUS+ytyeNOJ21V0iV
Ql1N31n4EyuViE9b56L6F8+WHEX5a8FyMX9R1CBYbFsZCTSO0gxJbcGrfZ/smleT
QClprpYnmT3OMq1n19hBhQv2yfN9kCYxX4EKjU9FggwI/HscXeP2ntI/WC5PVS47
5wewgJ63fpXPZDpoMDRVHJCEe7roBbZcotDPjBs5Zt9acnWloQv555N/mI4oQQ5u
y8Jdz02XERNNE/Ip8/rc5WT7gOE9Y9OBzP1Eq/SyilVbr25Pk4KRFaoBFZsmHMTW
uflUAxEPOv5ufZJX6krl/VHfUfaUHU3qrLkMrlayVJ1fCP+/8qStGKUxoofBXW0y
XraaVMqGfq3Q4CyXHvYjKHIOzzx1zkiiT1vWEQlC30KOcBvr8a8uDgeHP7lnY9kl
SOJWmrCqoj8sIK4p2v0IhBKSYBFsLsDpX0pr4QCXQbV6shj9sgHLWnpccsB1jC+f
2xKNkRGL/gUSzODgHUzIQY/ZFhcncjiHqlFA2GQpdwcCChcrRhoFgL92TXfSPGhg
Cdg/vM+yosNxeRrtwjGOd/qdZtN+08UOLTrl9DdkUoSHCZSa1H7Kc3xik34Rarxo
xcFEbtmZ1L5vn87H80gl2blAaMnlU9dd5zyQOD3+z31dpvXHVhNwwQo14bAaeoeu
GIQxiOI6ZM3Wlsce5DSYwxuNJq5GRsAFq0eHc7oTVYkw1OXGJTJ/8aSZ9JPtMbHm
jv6muotk3KqsZ8Ue9tIefskZHYDL6AywoDEST+senIuJWTiIBpxojP9oYiiwQ8J7
juYn0TDWtaLn6865g4+UFs13Z/TVLnFk7Q1BuJ2imckuusnbeVm594KVVAwrnPnv
pIue2v2q2kKwTU8VTCnustJr1cx/TqeUGN5EbvNoETPSVh6ll0OezT/lwZFRyFd+
QGmcWYQHeVf6bDsWwrBohgss3ioO6h3d1vuC7lQQOLyBx9g7q2AuuO4ebL2vbBNZ
8x0iPmtBnbgcxeEd1XZflFNYo61XlcFFZZX/+WeKIWdfVl6o8RQ9LR/QOz7vNa+C
pDEam8R2+b1MajLwR6pHl8YjJneFCoo9lXpJCb6y/iKZeS5gFph54/wr2hqUnU6P
myaGgVPzvHZYami2hXCMPnUlJZG5MZiSDjfGQtwTx07BFhqVS6WpjS3TWrZZLjNQ
N0F5Bu7sJBgDWVJahwK2LHZzj7enk6iwKQPxgiILEktRY2Y42Yiirnj0Apu6TR+J
ShB9I3GilTCUHAJIo6FyY2VucCNu4IFr/ZqelBJ2UsTuLu1uv9wNARDTi3KcHME7
YDZdEBBbFRVEudCmY0NZFLkgyfZrCRjlzOgShCHfVM7tFMh4s/Md2aWczsju+XP4
PZN/ekEJJ/47X8DlihTalYuHDOifHnTLe3SsYbMNNhz1tQZ9ZyiI3UdEFg/ten1H
x19I93rtlg9fTfkcPEh92DsX11Po5KfH5a3z6t0P0yVinB/x5cUsZdOtK83R5BvK
N76B395BhSEO8WKz9fzA4G+2Df5lyubHndRRSRX6U+NqYFOpW7Zyn2n4P7UKgr3R
ge9ipZv9fGCLZFnmMXf5QQ9OjvTVgg28V9cDB5pb7lr+QrHSMqQRLDStthUocjwJ
JKydXQMfqYv1+BeKOyn0dURvxZGDrMqDUjSOvwSnaxbUteOe1asR/f7HiEeig/HZ
lf6SuX2mCNn+XdruV8OrLW1f1N3OrnqrshHVbXDcn/Jtah/nADmXLRkYlJfIHjEE
Q8M3imwTc3f6z8YIfMWyKlcnGGaJaptMPlPBnVwoGwXDg+Y9311E2lqqdulGmkm3
SbK2D6OuMG9Ridjrv8ciBNOKCkqBI9uBHiLikD4eFBtfO9OgW7QSc72bOQ/QHO4F
In4SvwAGl5TvM7AuAkZblrF1JAohmzQ6RcfdrIJ56Y81oiQ18i+v+BGnPt6S4loT
vFojTXKOkuY9+YMYfGVEKjG8s+g/jcyToSD6pkTsq/rP7Sx3L+R0HqPSWbSuLFEb
TlZh8xvsokUHdHacsPGIHWhCHj9VAY3rm86GYGbhas3laL6naJSx8hn6Kfirel73
TCrHGRPhnV8pIp8BcTs7xeBvQk/P7HAlOtO6agwVmNb0eE6WhWDzmSYxgC+bJRno
2bA2Dx0eqaryg2ih6rB8Y6V0rdvKt+k5BqRgGlX5v9tsiZuSWmkA5UFPjOSMv/gu
SsPMCDGLXwE4yxwq46MFZP38OviHF/6wRLIO+/rkAir9+X3drpR1YaxAuCRhcdTq
EknN7ET6YjVCxirkcbyNX8F6xK7o0KsMiNfKSA0tjT3cjoufh3MWCb2lN/PfaJ15
amuwMsjd1ei46rFz4UbW+NG1cTwpefBsB219+Xs5P1DkAQO6u/TZ/tPxhygxBW6W
Sekn16Q+xtxiPIIZedI+LgA6ujP1uWFbueqxa/t27o2e8AacUT84uVqySfeZhReF
5DdlrlbiLq21BmabJsvBW8zFSXgCKTGq6QdfX3KG4Q2M2DpxFZFZhepF4LJWaI45
ZLSPAXVxLe9nvv4RY5bMolYHetzwrWnEsdZ+zXs46gYU/6OA31Xff0Z0fkzx9T7M
zDhvegon09Tm9AU2I3Bcw0ynJVxWxG/G5qiX5kExIWQozg74N5XH4en8lXorjOk2
N2CHUNhiGcK3wPNryCWdjlt98mVBLqCEDaiC7/k3xyPDD8Sfrtwr1nsgdj39NrAL
slVbRBOxSlHNC1eoVMIFF/GX98ncOov8zLKIpYXEJ1YR7V4cdaNDxjHJwZS0spOY
R/BGqKpyalR6uH3GQZEai1Ov4A2KgbQeC2xlzr1lQEoGJUahbErNc/KdyUwlrMK3
nv7jKAzfuNDbJcyfriCijmbRQClzycjtb4LOdzBBUiWBaN8y/6l869zdUCfnS7iY
G3OyLGyCkG4qRJBcBqgXP1XPaqQvGHie11Sfft5yz4SJ339ddfzqJ+1hoNV/ZDqF
J8UplF6pzTL8qIcK+aMvyVb0TPndSeAwwaJUyx/CS9vsyaejBQM8r7e6rfkDOx62
59KdTIOJrkYDFxoR6pZW1GC4xSHaVSJcWtJCjyMESffPr4XzbqG+QVDiNOl+1EEL
7qjKVjR8t7esMqmeofWIgysVKhsJrgFkihQrAeD8DZR68emC+LJczdccFfwgzszR
XHZ0PJ7IW0S643m+U0sQEMoF6K7x+tmE/VM0ij4b61BoZbPMLNaUF2WGy2HM1/BM
R+2HqK1Weu1KzRKHebejP4swwTJ7pG6EYOJo6ZOkC9SZKJK2A5JDfFuacTuI75xW
CrSGt9i2nlUNPkl638XoVH3uqio0iQt7BOjIt3b9HT5uPGlobEVciKFOvGk/lbpk
K5NT1FpFoRPSE/UINJpN9ILyLbzC60Yueipj2RHnQ06m1SmRfICSOQdxIB9amXNW
TgRLZ6RXDJqUaDY5BECGAYrMLtaaLBGcUyyAQRbK93Tua1NxGX4F4PRs3pbv4rnd
iE0RxzciI14ZDbwU0nOZ1KTAgJ7Yod4YmFyltwZGQjvCLpY8vhhuc5TSAEEUctQ4
/0UQ/gA9M5hkBBL97PFKX7sjtTzuUc+7nb/6FEcaJlaThDJD/ZzsackPaGck3wDR
GJo8ik/qVKLZ24qYcZlncyzSEZPUW08m10ivDJSW8lyBOu6jYE0Zddx0ME6BrZcz
OccM7+sM08N6AP3zHeJAFANzzYUZocDYMwEWL1xde1NRvG93rRfgTEDKQdSTWbzP
Eyh/Bxq9vT+gHTs/hZNnmJnIIV+d/94WG4KqMqLCuF3nTrrfGwgnN9NcnYigd19k
wfG82/sHKoV3OppRZSTQEwbnRQgyRwZTrIP+PugCVJYl9+CPgL+wnV/TJ4xCjtsh
2cxX3TDWDScjRuMj44p/cO0b94Z0Mm65+gnJLZJSsZAaVUYvtIoFKrGkUkGFxr3+
o4uAdRW3uybEPkcdj5BLuae4l00y6WpKHN/YNQzb+MBsxlWxKJhCWmZNOGlsRQGe
ag0m76IzSPd6mygoxb3zqTDCeuRzecT0LzGGVk8OChy6D8L/NrtMaswRnwWuN4UD
F2IKqB1kLGHkAgaUknjFsF78HjGgyRNfYc/Knc3AHS05QcjfF3zPvORkFA419uQM
gAI31K46iF3gIcgMMtDM50C2En5d9YnuZP/pGPYCdrEyCwxTsq0R1RLuYLGV/EKz
3m7fCPsLiMT5d/pxO5QRirjoZWbufyreQVKGoBiegSqkjCK5KFNMItzh/Q60LM9u
7n1wBq9QXVyHBFtvWeJE4AD3FDKOmHekYiv4ha4wKCtXKlUFAkYQuWEXFCrz5vVs
ATbNRWeG9gFti+HibrHTX+T1c8990ppbeadMXObPZWKVvpXIF52vUw5sS/KE0nQi
+uNgczVjIgEh89PKSLGfliYJLp8NIP/+p1erxD8t/cxBoGQ+t8Qv6zQPp0mIGtYp
6umMtExBZUfvmBc6dCl49Qqh7bRTjI9kBN0RtNTg+MfcN6q9+qXCQ9dx3lK8W/UI
n/aF2lZgHrQGAyznHvemthPryCzvjhZawVSEfczL4aGnt3SKZ+Ep7VC7bDSmfAwK
5O7W+8FWgWIJPdBzpOPwMMpcfgqeUjMYGm4Zps/wRWTqRD5ajavIh0/TMaCdDhW+
kvwbfqJ6kw61aWdFWPbM3m1pg1+luT/l5r0PAiFMMygSt34Ey561OrmT7gIF1ZLW
dlsuMIBznuZtj1OAHYv/RQD0kRJZwk5NyNrMgwu3VBVFAG85DbdwxO1N2wbflJ9o
eJfrTxurv+0RiUsCPyBKWjZehhgPm6Q8fyuxELKNTCb/YErdl84AIL4xWJjkF3Cw
99nzJg2MMd1/YNd2kUIwB+YVW4KJtkp1GzteAOJIIGIuBd4DT3QMGxjMA3mD37NT
w5eiZlNvnywzHgOIL8yumxPQpP02OvgGbQ4GfsRNx8GiPxJWO5LLW0+3FGiuYut9
EuKuI+D9tSS7eBhJ9ZswR156Eaa9xKJa7rJ60pPazjqqqS7Tf0LcfeO4/WS1gBuF
DxyeJzlQvDvkQ4IIJd2rKMYaVai5Ows6h2L/BCX3SYo56xyLgvmUEZrKW6uTfhJG
Jnw6j1GkkkLX180Ll+4JJa6/MNonpUQwmsxT4ep1BLSiAGAxu69cNygcUZv0VOz/
XZOu13c3xHxr7qM7HOi2Vso1PhMXR2wawLBtFVdTz4aOkKBl3kFMs/N/kXYVNzaZ
Kpgrvzu7purysPq/99mhBDRdEWC0CAfa0kM3vGE2zXnM9ynTYn5mRmcCuJiTAJXC
0uUrEC/kHWwDD/bgpBc/d+Ej3WuH7kGYe3XyytCQbjGoQ9C7IS+5Q67nT6xxn1ti
BEXfp1CFm4NBrWca7MM4vuCkfQJd2LnZBpsxFvt/CYzBDXTwhWeP6rl33YZwXj2k
1WfbBUZvBJtfrpFId5BGpUPL2nfGF+JdTTd30RR50llb9sC4/gkdRG9FFuPWNb52
UB9a/+mJ/V4PDnjWPjZMVPkNP5yVNfWMEwWB2MrHCIVnnD9OQIcc2PdpEMhk+7JQ
AN8ZBLZ/QKEPrFUbzG+izmxxt0gL24QfFHMvAcASu9HRcMzVJ8zOiKNSvTZtS7jM
bqwTmPIZLrlc/ISARnUz4q2m3AEyNpDKlCHP9Ss4H2Uu+o/cQyrouYRTI46lko6w
KTC0fOAxOPQdE40xEO930z5eBNiOVbkh4dKKVR24r+GOcTR+Ge/6mXY6YMQ1/o8n
b0rW+nWxWe6P25m3lXTvNw8KQO2siYr+U5Ms9awWsYkUgZMRvIfnxwptMk6TDH+t
r4Ds0MNVaHsqz+ls3xBh1yaNdEAI47t5dk4Uj+gBSZYPa/wjFogZ7gov00fraR+w
XKC4rnb3Cyd/K1pbzgSco6jdxqeL0s3n/HpMYKna/hW8KEhM9GES82wrmDSiGKzD
QfKf7s6t2706630G+phet84xPBt6xU/8bqdgUmj4Peh20ZzMwq+eKuEGiiARkk2O
j9ME6iknc5/XvEmr18vZvpKpMVCE9MXpyRiwhnRZfQE7DDrU7HFyrU46k/pDJv5J
43RLhUNlliwKO5cWmZz160ingPPD/CSNGJbZjIgC/VN51epxvJ4RpJLebU3/fTHa
RlJTcJzEjTz6HBgTXihUkta0Ic3mMgOsG6Kg/ye/c0yLR30Gz5cw3bP6KNX+MTmO
PyIKnIWQyaHknjmvG5CbR2iYwcA88ArXe8EAoHgQrzu9zwJQAF/nLDB/1yZJqmIG
eWJ/nCJHHJtyJvXDhpXH2v7QT62XyAFcCl30s/ySBxgZ0iLxHUQGEbETxXJgQkae
FuS8gHrLWQf00w/TSQPIWdEwBPBgsRcoh2/DNLTIrAd/yKxNqk876x3Lmk0fxr7j
TRFQLzIz9n5IB2TuWK+suKx2W/m08NAlXTDSuhzE+DYl4aBI9VO13Hbt4n/ig0LQ
axwwMRN+XkyppyKLJJe4+qN9EUUrqIeb6wRWw+Fw5ZmVhgNJFWrn7zQfpzFu0odf
ZqThGdnSHrdo/F7jwUK2FV8rZbrTBlmfHSVgT/+xFLoNIJy0o67mdTTOwkzNXm60
I8rBnOY7rzr1xoz5sEKg7M9EOlTLNtrb4UzvhWxiLqZplXbuhGKwXn7u4UNPPZ4t
mSsdmzsY07KUSuaYim4tUMU9d+r9lp/iN055PBL2DkgkhagXHN7R8y6wvjqQGCar
5w6+54nTBJS9vSvRFbFCvOtwrzM2GgXDlIAb6k6U7eNolDLZL1z3YOoyUjpBoJRv
tid2Mu+tx0zk1MhAkIkd2PuO1bnpxf7mAb890v7uM78T7v67naB9qM7xwtRhJZMB
rBhpQ3nVKvujiwShD1SYw/nHbenrY9dCcHAP+cW4DYbmARuJPnS8iMkflxhwjaEy
NdFA5Qzv33oSPUhQG5dRhjI2IUSXm5bSzLP5Kq76pRhXYqsNA6L1DDMz8z9awofv
YiWlOhbwDzUE+q613+ywA/8ZppTngTvhReK/cZ0An66CUmOWbKtV0LIemfsIh4yk
hlGWu/JUVCOoKtnxsJ/K1xR7rVzNQVbxSQeEsIpZxw+Of0/Gpi65ohGcP1uayTl8
cV4WUCdt+XX+dl/aWV0Omedl7lSS+M1kwGIxCux5l2sv+83vVKSPg2J6pWhVCUvC
vfVfl0YQNbHqxu3tGO6A5I9fY/Hy4YvVns1vrPeZSpF21fmjIRdq3w9jfiBKYDpB
SMX0aMIFwYXPQEAQI+WCKPSsZgZmPnIZSTZh9/mG9KJnruP+j+nWgTIjoUCtfy51
Sf3HlY/9NYDqiGGrhu0kw+nCsjNt6i3+Ow+2uofSCdM1QXZ6LVgJ232C7VxkAVa6
GT4Umlv1K27T76Deyv+FrrVocyurCr1IWYQbhQ+nGTAXQ6JNb4htxTKAg0Vieo8s
/ZbMckXjd3dJz3xtntzC88pGRntyBsewMsZ43arGY2nP1pwBtaMVZXDUIT/WIwHd
XI9lz9CsK93IpkBSApjzcMVBOZevXGjTupvRrjBhG0NIxBqHg7Y0kKAEHdbp0JrL
NwhKhoOLlCvvL8TcN1l5xzmnhdFdzj6NTmUu7RckSl2f7QQlTJn+6P6zm3LvJ0Pd
YerQOTPWRVblb2L/8HiucDLjg071GkIA0Lbgc73/4tgoy90jdmn5sahtlgUI5vSx
kNNvlrdkzl6DkN7LVpAJhyAxxPNOuGy2n1uLEF8mEsYY2fR9pboYpLN15tE4RVji
XAy/WSAiCKYHrXpygxBr4+QIfXK8nGLqolR0DSTs//GMDOPQlcRz13MwF3hWTT3Z
Ifb4cb4VbMu/YUORflf034JlC0l7sVVYUhyNStGSNBQ7NHRHbcLmmWZVgXfFzglc
1kNlESBnMiIMjTioJ/o5hIOiq+vqFTbj6SLxciYPZt/6R7PXw9CWjMzMSbY4tqdv
k2XTFQkayfiH1G4xGdTe83SLveC3ekeC6eRl+Wpf+CVYhQGnmPKcMf1B6AGgty7f
1oJmN6Rnn8v+cIJfV4IDVZ3U7tpGmMNfQuQP+Oc/Tvdt/akg3BCihXvSYX00eBgh
MM/nWo94KMRWJB+zbzBuiNwl5MqQGk0l5YLmc7rkOZzueY3UWu2l5pwKNjo2xnPB
q96d9kMtuhDb2VwW58EPWqL4SGL+IRemWICQbvyA0vk7iAeSyiU7kwpO9sNHSYSj
LJFhS3z9JTuFPgjiH+AZdJvoNVcees+zbjXSfT2PFlW3hSaTxnGVxMvgBvE08ypo
no7HvwDpOMI9wNZzq7qYWShoIajCnNHLyvi7T6pIuZGe9GyubtYV7Waa75Aggap/
6EVBynKCElIKQliWP/Oo3sywq7jZbbopT2Qrth/Nl5gy84Nwq+R7O3pQ6zVdUbu4
nmDDKc7fGJMe5dJTah5WqcRDtIRxxF54X4DeRc96+7/uMmejnsA/jxvx3aPAQjbb
c8GUCe3hZi/sdrZ91aig0r8OeUvUsiF/7g+qEm8zfqD7OOmQ12QugBOVwJUmCJEV
t24bIut6UhBJOz+bWb2xcxo80n/8TFGLRArwzpfWzeSCnhwLon8W0zO3JKU6v2nW
m6VrqXvTaHbEfjJV+XjkXkhz28Cte2lcl00IAmfQ3SgevLF0UzYbz4f5R04gqTgc
3FIuwt/lOhshczwT0M31sMGP3IcMLyehhEDOT4LMDJvsXtBZhF19luX+adRoBDC9
yT0BNucJVYrx11/uml4i/Rge6yxcZllyDHlyG3gx5qndMKM3Ih5003vtcgVtmWvB
JGxoLhMRZdd50HMVBBETTJLreUIbOCpM6ZjBMjbRShp9TKtY3Ep0VLZSxiQRFuBf
qGYFlI/1vo5tW3iQcKDfbsHYsil7cTusZMvUxocAaDeosXXh/IcxpIEjR3dzTBWZ
AdJwibDOO5MJHDKepr3eOWtnpgfx+T5p+S4pAiFeke99Taxr2hCptM/JOSnlmlo5
inHxT7YHtJ2j3muO0/knVN7mVPvciz3RXieu6EqrORjRnC2qPBPaOwLjcXi0JLcN
nFOI8QR7s/L/sV3CAygTTapLJxlsemsApDZ2V/fTY5JHNQrG46/IgCmaYzSIHqSA
NwmaT+ML4FEbfXwPmIZMLHu2YbdX7Qexgto57Vp3d1875gtdGozhjqSosEDGk7OA
1Ya56dTKLWHo7ZaOZgex1w2eSjhefAA4XwZzmBSPgpHbTms5s9FrX7fieNtByQtx
uYURflS+jUl10o/3Wkx99OYV5zqcd5HgwFfk5bO204TFJ0RPZqIIAfhF8x/1aXU1
ao910vj60tex64QvXcQpuL7vacvb/NwQ9FPRdXay2YCVz6sEeQeaq5rhCKE0WMA3
iJGXlDGiROuBXthYuBT2AMGY6y6TtGM1sCYnn7LcjEUgXpJO0rYZwQUyPyTbpape
oOH1PRtwq78Ccvv5DeXoUk0RlMKlsu+D/EUz68t/jf17cVdrmDutLCDbm7PqmwLl
+mSG1F3ZBtsDLZq+uVEGDMXoWPUbh3pREl7j5DT6VQHn2HMBKz53tm1A+umMynp8
5xktskB8m4YQqovXsmJ82tjwRSiKh4aIoG/OPPDSrEnO+fC3VZKf5UoBQfx5PL/D
ucqzDMadnqe5blHCO2RT6692IQfUkCkHiaiI62Imi0awYJ23K95c4ctBibJOd3E3
e4abiTpi607NE+JOOAtKJpoMnZqCib1TyEVIj9I/rGMbScOxdVhZaIXRT8UdmnYt
9bO1u8ksTzOf+6HKWzC524WtotNt+rXP0VywrxnZzB3n4hApJ7bOCOh/ybwDYuX3
hg70L8rKSOsIZyuFKYoa1np/jxrhhyHp+5L7Uel9Cml7ZHUo3Kw7DNgw2O/+KC+5
0nsM63bSGBkxdngVon19fhhbIkAJOqpOmH5c3+w//zjwaBZ8e8XvXNh6Z5GVxQ4q
LKsBebmPQegio7V2ElpySnpPeq2Nl5DTjxYpJQ5OkNDxgIRoTaiR6z+grjrpJG9m
er1HyODV6hmj6TYlFEHJF6JCJFltQxu8nLF2vJeKUIHbYwgTE2KcJBZ9eopzs4hu
D3JR1NOmINhXhASSj4Xc9YAxnWifIgItDEl2y4dB8MpFs2fhimib6qqGAqa9sUpn
jS/yMr1OuO00oXagmPgjJ3JUFVPZlGkUkxliUvzCvJ4PZiGPHeMRn/P51n+Bu0wn
cY9jXuLzJhPkCRR4JrnAwmLsdMtSzSNFcFWdxfq60NOzlkljBa2bDxA8EpbHOmhT
BFlZj8Y429OxHJtWJCf+9Y58pA24cT7AukjbjUYArR1hxne2toyc3etD+KSVwvq/
/aBDGuHCYw4K+5MCKVnzATDy9A3Ac3DqLNhcNDDjlJfbZfI0Mr95rEhT60wjSOqa
s0V4CsQ42Ya3Uc8U3Nkux+jQxAlNG/hIyiZKqpNltKGM4GV1P9n6f2p/2/cWQmay
wJNZSUt3tWvZD1bX52C+HPzm0Wqbn+wWLRiwabQz9n+zMz0WjpsNWhJnFL9IcK8W
H6BO/KLKxRTbuAF2nbvXcCk4t+F74PPZ26v/ITgK8cXTQ515fMCgMCY9px6vWvjF
7t9H+VVHntcDG6rOUGV0LhoDuJH568kUJ54f+lp9xXSDBoeZgyFrPSRA+Mp78KXL
bSFfQcgv6giTIsUMRjZFU3R/Awh0YES9ZrVfWJcKnr22MuHV3ns39xf7rQPO3Hfx
jOCqgNM6mRakFTABbQcv+no3Sx0P0Sd4ztWvIBRStE/o10fepx09Z+jlXktwKbDO
OX9QACamfYMBLfdd6FKiQ+i2shsxmkEe8kfgTmR4ENk7GwfgaUHAQztAOwRwo4Ri
18CA0kZ1Mg/AMTJeitXBaQ2cVh+Dbq5M0U5e8A833pU5X2gN0uWRK+LQzo56dkTv
K1buosDDbVFQJH281WpxdBHSmKjQyQEp//SuGznpGdDmNG5wFTeULidVBueV7rqt
PIZMS1SOXzq2vamHM2kEilno7uUt9ULt/f3Kyvu4Fco2rThjrZz2IcS2cBsTEUD4
ln+iLa9iM8zVpXRqIfE/cGu2ooGJSJ05xsTrJcr1q4HCy/F653ABOEoH03FX+tNv
BSwe8ygtFxETol1lSxn3TFAVBaAeu9DSDpPQSqRY2u6Q7WWJpPhq+fxoUyQZVIAx
Mx5jW3vhxIqm8bIoYML2nzMvbZx4Jd28/KR4jYHmIh629C0m2jNpLmliLqftAQPG
8o26X+85M2Phv5xHYzNF9D2jCFrZY6L4gSkEhxtT5nDAmvio67kIf3nKAz6h51fn
Q3si+aRYjdof28gozSMncqr/zO6op5ZydepbfGjWnoLn1CeVcJDKlxrpETfX60mP
+6BO/qhOLMZYIEFIDsmj7U+wYNUFHbGji9gtL7SM8BcNKnMSmNfMOfvzt4KaXvMQ
ijJuk7t4DE+m9gzWWCacYWlF48ocRBEzvU10vXt7RfzrneF0yEzim0/aanB2oV1h
XICXVecDQZTM0GJVIVPv3eh8iSedNwRR7a/uzYCtZRbtcUzQqhQjj6bZe+O4VJhJ
FIZ0k7HnL/CiRLu0nqtx0EVCBnCLccOVbapRZlhMCQ+k/r++ZKTHCRORHv3PVmcV
oSeaJT8qr+wxlE9HpyQqr8sMDCGYsvzVsLjfiUwap8Wq314Mwy1h3Nsq0ogmixNm
mPqLQosLSvewi9Ibuc0Bza3zK+aVE0irbRf2GrZ/ZhaGwMMKvzDTLTjcnpPN5p8J
QDCVIXzLsenooGkzSluvcieVk3WK35K2LtBlqs1Z/CqM5Q5f2W1VBLp4pxvM6Lkp
X+JiZ6S+rrIfc39sVS8JFhTQT1F0a/3DD9P+QbvClX6XoE+DFiEvFSP8PG800i3h
EeeXD1bIpZJ+ta9crEgNaNNILiQTlV2/P+6IiYPi38yJuB3h8f7k1BBa4cjTXeLR
B3gpagrJJEF6DGGJt9p4VBl8tWohZm74pJc2QmNfz/8fwAPU+jJx15V70PvXe1FL
WROjfadgXNFSr2o0fJfMHdJQObTbngKQQZ0y9Ytjl3Gdc3aZKJumDXXQ5JKEmnn5
PVG1eU1TnPh3Cv+C8lqV41+FP/0CHmPz/Rz3X39+46K85/waFL57per1jXV8hPkO
onCnzkGAKTKwmk+b1TrIkzjupsNaSJIHRi0I3TPaAWy68Kr5PJ5By3o6TVkCFHp0
W1PTm9an1z5Ofn1+EDPHKaTinJKIDYQV89UpUAWJMR7+vr6lwa941+y9QVsWNPaB
YM+y2m+xSB/mfaIvBhf2O02vS+WYIryqpFocy2+nTSfFE+IEU0PuSWeZBn+tLqMX
SzW8YCudD7IYeS8OPt+V/E3wrZ3vbCDVtH9ql9BnE0IYfKftD+yN7GHwTs9BG27b
OxDSaUdOKOgxevsxevzGaUYxppIa480kl7ZRfcRmEKozeLTwljIDPSz37Y0qe63O
GCoje1MzpCleZRgbaavd/Ym6olAhgZozB06DxW8IC2qmmYv+tRbZSLBTcX1H/GsV
/hn2lKh4zu/0eJzGrKDa26cXi77IKMvxBNocSulYc6Et6D269iQee5EtgrRPzHAc
7pu0lnwRtiZrYYVUDlDzG3zbdvK4xoKQZ2ij83/vfw9Z4j1qqgu02GEGa5yxS4gV
D1pGfwcMHbe8dfYNXThoT5xGgIk4UMAgtMHmaGCGoQE5466zlUYOMOM6p8bS+Mzg
T5B9rttc4qWXOmZOK1zWoBVKKSS3ScGb1+fMzEgL6hi1y12ZW4JIh16dabavU0Tq
rDJYT1tNE0tw+FVEF3ixqr2tBMjId0uyD85VR8jIK6pvcXVrfKI8K48XJEz6FRSZ
3WFSHWtTGZp+3X5P3gKq9NWVuBUN6ovZS///mHYQJ5E9hhUBEkCdCe6B5hkKhT5E
8z3uUF+g7r/00xG4MDTivkUPPmabDLZmPyb2KbzI6VKZCR1WYOHiw+/5mg9z5lP5
IZxibEz4CcMTpeccKddA9bbyAByWAunfTZbxzg+rg0jjb6/Dc4X8ahBrBBhxI8JX
VaOtNyJvr/fW/X+Us81fCdLlkyPUk8AZ3tDY6P2C4g5BDH4aGSPDdFIkuOqc87K7
JPAvi7HBqFKVn5HMLSBU6E7eqTJesSl7XUO+ioseistX0+s3fdjW2ZAYS4GyecMp
+IsqJ80X65jZ9rnXrVS2/cAT8r65OYmTHmhnOW6bAXjnFzn2S6aTwziXKm7m1fjp
uNU7ckQqQJU4By0zipCCPZ8sihjWMEC0NcABiGFALGPQCnu/YA1aoasusBXCyq7B
lVl/HWqUQPNWXLROnzx21lBB/dpUebiolUAPanr/rcrIBKZU3tg4K3SEUAsi4LJP
FdLtIvOFjJQwtoxLflfQohnYm5o8/uA5XXR11Vbxyte/qyQvdgeYaCquf7XBYMNa
cJyqc89iiqEJe8Pf9Ts0tQe0xCjxhE4JxsaDtdUgk14d19PerS5HAM603XGloyjC
lG50Nu9YP81LvDAv6XFZnOvtKL0X1KOJ0mjlsPRPxlMWjT7vi/ncDz/afp31hMXB
7H9lEqYPYzixyKz8hGQ8e9tQlLWDOrH/DNxZBjADWoCNWvIN/I8LnZdTDBznn8aB
i8GdClKxlbReIrNBS8WFLAXHWjflqOe3lo958sJcpEmXdrgGh40SQWATpumwRAfH
JCcPmvZpglZ5WFEYXY9TKjK+4sQaRixtqddOda3CQh/lex6I9C5stH6OYfBm7SjU
oQFt6tTH1qOuhm7CirFOxqoFL619e1ujB0HMp5V/NQiXtCfVTAogm9JI2eJwSyC3
nVG4z9kcE1P99zMX3pRrU9x+hv90rORPqkUJvxx02JAwyDJJjyHCA/OH1GmOFrhz
eDh0TsBpgADJf8lV4X/GsWOtrXmPzpTeYDw8KnJ8AH/V6Q6qM4x+kWKVEIBAWoH8
yeEIhwJfIKzSPQNi85aXf6/ZZ/1fvI4KPo9jrTGg2KFjjYvgagw2d2+fls0QxLmK
J9RHQSUl+zDW1I/W1Pb7utxnTS7AZuZE6DvxcWIV53x+STL1ReyQt0VC5idepeL2
S3XkYBmMyJve2yCTn/0B8EOQUig6HnXFxzcsGY7eftsJ5S6nLiuHXNZECJS0wRYM
4Ly0O3nRTDdJtRzhar2alFwjO2bLm428K365rDuiBzU9cxtIkBpvO03+t+27VSBW
uZ1tEYwuH3R7C5/AacPB1PnXgO+f0G1rbbIDM1UaMzbh7RoqaRaq7t/59WQn34Gv
Iaan2rfArLQSO6Q89D9zDZP8T2daXlbbXbUOCSMG2ZJkxKBoHWK2PuzMs7Et41bU
M+PQ5A7LIHl3hIOHz8f6kGflg77nrMCudO6D1AsDCTEpm/6s5s+i2+09jejF3AAO
c5AP9j/s6SOGfEG+FR0/FImLj4XgDknBHeZPBFBvNhqQWvtadNpSPBIuieJ7Zs7s
EpFGWsQl80zdxDMvUrHP9nI1aWbsEc1TG8GKY7NsVD83E8qbxhS/dx601LJwAKpy
zmODX8f3AntWc3XUC+m7W7lTPfGHEHYf2hQsJt12MmbuJwcW/+LjSGQqmk/OP3DO
+4s0EiQuHLqvBEt0j1b5T9D9fx16wZKvPHeku8aFlnOA6PHSenRhxetvf66ytTnn
LNtyGsLOMU4N90WWbC/c+Twsgd0DF3XrGtto5pJPfvXDoLILDwQ8NVWt6LCo6TOn
OAqGavpf0Aeou1VrR6AVyZVeU2sW0kGMHL7uV9mbdHvyCQJaUGMABjtTICfH3bgc
GBRir/CLMoEl16QwnGaV4mEus6gUL8Wkja/ZlzcZWoeAxfF0vGaCDwdwaYdb2JmR
NUZFSRgfCUFuidt9rFAAGpRhraE17nZUFkiId/Lo2OEzt/LlyrHXWXKg9tgbnY0K
lHwtBs5IwnC30UGiiD14PtV3l4XcyNKFsH3p6i5W+h8MtE+z/st7r4eZ3IyG+PAy
ktLWnJ81jxSWjzX1jtjHYa59N9vFQjTuZfMzp3zuzRHsDkCgV4pPPqdBlozgo9VY
UuWpqoMKhuaanLgMzhjOShR9DyHzDVqJvcwXT9sWg67RO93oBPvB7BS/D+fMPdqG
C3ur5YiWnYqHXP7M+4Mh1nV2C0Faj29nrOSssQGBQ1LBxcgkydMiAiDuozZCe5ZG
ewYQF5xuV0RZz+ih9BiyJQZYmeCLloK7hModANzTCkWm4D9O8IPnZKpFFO6XLprI
+9R997aZ7U+yr6tPTLBeAEagVQArkGbx8zT5xDsLg1i28FyMZzTTfmkNO5tdMT6j
U2wPCf25GStjrFboJgbo2JzyXLCcTLteGz7fdySFXO4ll29pv640GYk4HtF1MgX3
4ne59TGubgOJBppR+xQkST/6GE9KlfmZWeSX7+HITg8nqKYK4BV32usVzQXwldte
EE0sLknLb0QSXbFozU+QteKIK3cTp/rE2cRCVx0WJlhlGJTrfhnPzqGApRDXTvJ9
0JovoI7NAKRv4JoQm/UtxC+WMI7tKlsesOaTg0xyyPwwjvc9zcP/o0eCnSKD9ewX
AqdbM2DivJrkt5PKABu8yKzvEu1eGHb2sA24ONh0wDUZvFua797i4tiK+44nrsA8
d9KjyhZuyBqKV5oc+ckTaxgZUsAkizXDyv1U+KEytWHM0xHC8DDFdtZ5Wk5ku95L
jFZ+FvmrOgrFHGP3gDIDwt8/ahauKDtxXlgGe4RVsB5v9K9p7J8IUulavj87AOdZ
7fCg4BfIgMjI1TZZoXMBnKaM6KWGdRt5jXrlxQ2kdflWx38Ma0NC3S0um4C8TplF
uTP5FQKC5orBX4i+n0QE2W16WOhezQJUOcB4y9EWUI9sPG6mQFHgCimXNGLNb2k9
noFF+0I1HJ1MvdO4E0K8MdDuDiUWCJFCkKp7pulU85gbP3qjoqWaos4aPPuTlq51
H6h8UFQKrBsOjZTjtKarkvoi4IsC1SP7VReTbjdxyvLCXM9vcw/VUcwy7GCrSInZ
etR0Wk/iPJXXhWT39aI1pEx5XPQgQXCmPF3uUchirgXqqUGPKVwffbewOJuzevKh
1iq+m3WAW0rfXl6GDuTFEr7RXOsUlCXAUtepEHNOZPViBirmk3iZvxDlWtn/a5zS
85WMp3wBUVdlKvCStgqj2/c62gzZJoDzP68yz4sDIhbuL7phkoaRLovpRrGrD+xI
OC6aGjonEt3sKfi9dBhV8ZomUWd1AJqhhgBRRmOjsOi/PXxf1/fEw6gPWZe2ntkr
KUakXPsEqULW0l12gKnhPboZZQFafiry5dwjN8qXscF7tGFW1DrWM0V5DukSIBuj
eYb6nX9MYbQwhy0lnxdVqP17GfnbVA4X7xDnSxW2w23Mf3jSNKsIa5Ho7d18ifq6
rmLLDbvSmHYuX+/7ZiQmnceLnlEFCbrtDTZFMhiopHcC1AglMjM07YkWN5H9cuRo
HBbEcRKoqCft0XkfiJYgsaZoPuJ1SHR0yI0g33y0gOfXXrzfXZKy282cC6VxYUyW
gMH6vYCq792J7f7a+dF3pnKl6D9CXpx5oFLMEyLGlefoC2QBeXVRZL6/Kij48R/r
cA5UnhzOz3xvf+1248KQx7/A1xyhlTcx/HPu+7EFhCx6YCRkDKnJaxzNLb71p+7I
xQcMszZXJ3+kQwX0A+joqn/JKTfl7jbC/FfMKtd0G8vNxK7St2XXgSavLzwS5ghl
DPYg7jn5IVhufoF/rfrAq2TdSy6PbMbbTUW+mvXG34l3IL+RAjIu00LxpH1XykBv
6tK28Ah7I09qGkYEo8l//M9/X6/6k0II8KhAA5pJraUce+B2g99vDpJ0bFDA6SZt
IgIdeQXN2lPF9sFu2IxitB68rntqNFJ3skUm2cqMM2xOgANAITXTfHgmqTbycnTL
HOYZtJCbkS/cC19w1necOFskCorXttHwLbAMO3SQ2EjL7qEKhKOZPDwlmBvKh+3P
iP9l+qa65Fql6t2l531+PP7Yi01B4TT8bTiZfdz/nVNqEfnMRb1QLqAT9RcIa/mT
c66oalvDzU02Kn1OU1bzuxMOXNMFOnnIBIvgl5B9RbHUnW743NHrlIoUZoT7kN0p
rXTMFwVOio9D7CuqNOtPk45kZU9tL8iz/7nAmia/T2QlQ1PTQywXz2TNaEyizbe/
pquPCSzSPOuXnHO7NeCYgo0eCMOYL3/hH771foeVu/cMystvXT/Rcrar9Hj/hsI+
QCbTXltyXFsQ7LNbGJCEUPa+npBZbn6sUK0BKga/1MiiToRaNbnahPbVftk5HN7u
Wk6QasI4HcsbHZ8a/QPIIk8UpUK8IVZiBnzOamry31YFO1QWLnGHet8+GGsu9hwp
qKC+whYKR07AtCiBRp467ESiHJnsN8W+KFD009F36oDmmqzOSGdn5e1BQbE0XgPn
Rwde3BXu0qdX7qlcipAoWHtXQR1Ns8wP8cODFA/n5eC4BE1QL7T8eF9FP9GYQs6A
0JkCRO9cIMJFIq7DSvn3cLxHkkuOUF7yO8Z2oEB9yz2UpF6F7BENt+WjA+4B68ST
tzwXT07Mz2iN0FruUXUOZTkANivsBI1cynLXk51aC0WTCpjPtK94dj5CGnuYrAZa
YMW8rOGZPckVi/6vHhjREDQ1fkpM5mGvsMi18lU9TQUat761DT/6W4llIl2Rvmfy
G7m/gGmpiHoGHYAZbE4yWn/WLciUbFYPO4PL1W5yJGdHr9YIO74eIP6/OciYnGie
68sM6gcB4Rql/YnRRjvM2lQ15NV1OyHSgb3VcyVYtm5MsVcTfwu1yG3dQsB6bv3C
Aua9+d3rdAtnp0ENWX3xbfxXyCXA5Rfd0BcBFo6OtknsVSRiDy51uIo8vE/zbs4f
5ORd3jYbRa7ofkFlEBuIdv4ftuoAK/rmEoxCbQf2m9l6ziIR6fOs/vHyqxcNUTNV
/igcJMwarsY0bVcrmNmiTLKGqtyGNG7aNL7FHYW+J66SdfOQBT3yBr4TPAsxvx7H
XjRp+GoQvPHNLyjFkqyVmSRi7egcvIDoCC9MUa75nbcpPnvjnJ7CM0ortiB7JtxS
0ALY2MEccBNw/JgSB3yVRYebWcwyM5LFM6z56mDUmen8l5BtoOvarVi5a/z4YDa4
YEuueqbWcwiMA5C92ivZh3Q/dq5wntRh3wcyhZGCwbDhsTWy31sWzQ6SheF/W7CK
UvUDRGma7QNjANHyPeRS7ZqHX+0kqeYvJ7EEws9UbD8GLwAkxlWJat+ysDAj4KjG
v9j5jMIus2EepY6OMqJ+cIKtc0A1sOLP6hqC9GR97cig4chYrabp3UsY0k5m/9ph
aLVdKbFzdV4uOWlzFM9CvkysZ0UQ6Ddh0ia0ZHQIAmTRrZ3kiF5M4V8SV1b2wD8a
OiE8CHRNGF5SsKsMozWsjEXHDtkj/lMhNhWjZW767ScqI/fOyaYLO/qbxRN5G0Hw
kruFt7s73clJ0v3IkpH3RHyLGEOZCN7wdYouj/CGxy0gigDUm6VK5z2iKoc/tqWN
5n9++KNmUXtsoj7oPNn3HGSFB9Eg+Jp1wmQl5BQc/p9DLxjf4l/7xfihoBxtbtHi
78CtdD5XvkA7rqiy8rwfT3r/w1nOLQ0DpzB+sIZXLi/4Xs3lqSWqYiY/4va+GJOD
ypuQe6lFJIwqI9jTh18IQt3rl4h6AOeJ3PhLEXkYStGjal318yjnXgGLNOkjO/R2
zuARuzfZbkPCN4rhbocofSWIq/Bjtrw0WTTW84en+QD0YNL7Lzn0BZFsSwNtaem7
1dYy3lMEgKotCJK8x0aT4qYyxs6YHIeCEzFXZF4wQUmKPLqA6Um7WuA8Xv5XIHOc
uYLtdzsiqxG0H+rkX1B/jNPtocQ1Lird7ftl7USh3qqOexSZ6S9pudugaxBs5Ds0
fJNgV0BgDZdgkKq27uZ8dHnH5gmKJQ0Hls7CRpvA2fW95UgEL3AsbQT1K5YtfAFa
cZXAWXPR/U93boRyE8pUDOfoClhZTOoAQfTUELCkArmUYR02tyF2SFBIqLxdHHOp
IMOsJQm8YhRuKj+02p+q9Btd3TnzvgYH7v3NKfh4IZOv4pwyCXJd+eTAEmK7zr04
lEyLBUNZFOwD3pW52ZUd0fve2zo4gNwowFQG0JlT/jHlgMDESk5Yuk6cwDwsB84p
Vez3A6MdQHiY6NdcCZe3GGbWdxn6VIhgs6BFSE1uJt2iMF4Dr7Fd5HfgkI+dtqcI
J44Kv8zY3i2FlAA81fhAmCXMH4iOHVeoskS71Zlk9i2nM0UH0yKb4z7+kPusKnXi
06+ay8ZZWFpUXnokdPNSReLuFpmwygTx/DzGt78glFpf35kNOb+Vi0oL4j4I0opN
VxQ6GaimIAFKb0qqiZWPyDmbCY/os4pES9VtgPQIhbGHLOrxdJ23YxODyx1xg+Mo
ugfG7fbd7GjqsKIOmktUNc9ILnBl5ezZkEFUci0VE94n6hi77aC2b6ex7tC403Fd
j6AvHUQKDE5GjhCDIzjRrw56vVXryYZtC9GhthrBxrobWzW0N5Vp1J73lYbBdrmV
PmRibldQrwKpTiGeg5PbSltnq7/Z/DIjED6EJM/DkPKTm+TLrncu3kVv9T/xjQ8i
htGCti8QVSRDiruwcsNpP/AHAqmvmWKPYK90MsvFudK4G+DzghkaReU1xjD6KNx/
SWpvfCq2s3oSSqEqsS8BKs2IWceXkGlZaAWa7NMPQQXSIPJsvGFtgfF560XirISs
89e9v0dbRPJJsqDWHv7oXv8Evnbcm5s0/O6n5ul+kquCjC/Uboe9VTC4XkIBPaP1
zljrvQsa647ypdJK/Hfa1zfPZeL4WzTv8bW3Fo/ge9mdpTPuprA60dOUeN61JrE3
R+8684Oq8Q3RKn0GxNGZmXHan3d/gIiL3qcpCbmFlck7IY+RYi5v3/29zBis56cd
TIsIgPVhRlMyqztjIvj72QPkaZhUqJ2JdaytEp+AyOi8udrC4nGxQOeGSgjQ5AFb
ZP9xi8f/Y17ZjUwFhb/M6zDf1Sr21hDoB/PwF4IDnEjvnvwizXUvT1ZCy6dqxOlu
RsRyt9l/U9ghsGIeycTbXjF552nuakhdF00qs2s7IkUvhs3s3DD3OGyyz5lRuOfB
du8eLftE2T1XIDR7LPsEpq9LqN0rpuZ24yKSOfGbShvF8A63vTV+AyJ9f/CXe4tT
0jiF1hW9NecdjuVgKgPV87Et9krFtTLGBAmrMErz8FoxsFBczSCwCP7SMiwBsLbz
UCNMqxpzsZAaNMDPlSjVAm//HCsDnB/ooMBnR1tkUjY6Yd+QPI21ngEYE75oKC/v
yJiwFARGmmsKCvFKIFdnX1QEUY+0ofeyKHPa9PgsVlnpRO4QvnYgfnytnM7VjK1Y
m1wCpctXIpXDeZNHrVE8bgpNBx2VWjvzLHkAb2EpWEX2gYF0a8mOs+BucsotiubE
45XKb0hemGjgEdmf1AVKkO2RmFLNm0T5USvmQgZUWzxEUM4jw7oZSEpOWRERZ/zj
VNPev6hJxrWzbgsDAnotyIm9b6fcJlUAYt/FEYKu+Vukq/DBAKftjXPs81OfSqik
+OlVyh9o/3GSTDvPnwN433SQ5AnipD3bBg65wifCbRhqXfSOf0ShfuMvgwoCr+29
dVSWpyMD11hjjYQ+ZI5cn5qpMIDAtREJ1JQ2lYReT98UVJAXRbB5zZ0Dtk6LxRD7
vuowukbXBxS8u+O1qU8cTvggYxuX9XH3JN3hnZVSyZN8qZ+JNp/1BcTdOUhXANP6
ydFJJdHQpKjO3lfVh/WW9ar/O/xldhxME7zFxPbgVA/hGusWc2Kf/6wIMFRW8vL9
9f5lRftsY8uCSjz3nXGBitECt8yXt20538pdG4H3M7cGuCPjUFow0a47/C18Qf1a
L6bjPjaXuElFWzLfsTwPD2sCXM+PWPxE3kKAWcEip4V3sytbCx80C2LUMJoRKDkM
ku+IIW0q32x9iEpRKN8eh9V4bTaFqQuKYsy5/e4ANb6613RMmfMmc0cE+LV9Nu+n
`pragma protect end_protected
