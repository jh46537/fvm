// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:18 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rQt+g6KMU6JYoCG1UUfHM1YohpVOpaNMVcETVx9LOTGXne3BmihdgeoRvR2pnAaF
q21TyvwM6eF3jYyuQ6o4V6/oZZBKB4iPX3SRK5rAJsKWLJ5FCVyQ/M6F1FWmVWVd
M/iGf00CMc1rDsunudMGYcNDC2k/Npo4t/Z8o/1KomE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3296)
rtwzQ/VyFeRLq3WjZlXZQaK5atxIXRX4kE3DkoavsROoWz/W7Xfn4y713/bYSIPa
t/w0fenHNiZJGMA5Yzmw0ho0Sh6Gi0v3CSGXEErsbNgtBSmIvV+72VnsHs3uA9d4
jyFEMT+8KzuueQp7/nWjklK1hBhNDzYPVc7+Pa754fSF6/Ug9pJ+fA0h26CRJDAY
I1B10rxCcD8wknLw6YJ5hqqi09jaRKScEkjXNoIRDtQXuLiHMacPJpHXCqHXagSm
2OnC58tRVagwxbQ49xE3WU166eM6Uu9wuxjA/4wPqELgplVqKQV50H1IlfN3RIsL
/RdzROrL1QDqm+Dkgs0BU6DgyvhzPJWclXYNV9awsAYTwFr0g4DhqSlbeiD39N1O
U5fOsNIZxlcr+3lCo5gmYSnt5zBWjb9Lqt2kyXWVe8TP3ZjyBb3Q95bcPcUfjU4e
Ev8tldvM83U5oTDd/bEXv8XhkX1sZJo96wCaodP3fy7LIP94xZFs0Hq7rLzdfCnT
M1HwVf9ftV4GwnNdGKC0Fs7Ns0cu298V+TT3OUwdYfHXpnO+/7oUp1Er0tBkJmV4
19fBUr+QStkOUnq2aXoGdtJvRRyWwZttt+/OIBoWyZsVHC4uzDZ+tnwEYnCmespc
SQhhQuYZomtvCOfXbDjFlo8LX90bILFHWUSKBMJajfvhsi3QKkmk1sfvYrZlBJZ3
8w5LuDrcf84xDxafuF6ls725JXph8oPWB2G/Zf/QG3aQwKwFEpMcaClBBcNC0TXv
aRnBSHktBJSFC+OOdAPTw+ISfxiFf2/85aQ+Tk7JyP8+bHV02fwD8dmEaOt7txvN
sUGDLnJ4MfV/UfogMqjzRRcvjq2GJTgpHBXbmeryoeceb8YUnw1MmJEjkQya7NNu
TWhiiOIFuYEe7+rImcztfWmTwmq6K7otfjuPEqhCx3E++DWus9IBOBvRE0w9C/mU
22ke1qSgIWM66YD7k2YxvEGwYy3DOtEh4MVp68aaAhQNXhZ0UzoCFgK4t7F/Fopp
3Hi4xSIl4ihH4tNjdig9U85AOw2lkXcpX73EGPTbKPqM71J8NqIdiZV21nzINUIk
ei2zMWXOdLMg5Q+ENBQdtaU+w1aJk3I0aeWBOGQ7DNwnSFDLlI7+kg9pZWldzaOH
F44fnd1ZS2IVWo9k6h6Vj18N1BEjuB+Sztp01dqNtPmEC8EknY9S2sFPx+xWxUkI
e9tBg3xn+aVsLr+E6MGd3xduKBQydd1wSsyEHSEvGrpCbRPCxdaEvAmmRaOy2plV
/23VhDRusKC2Vln75wYFpv2Y6S708z3j2v+q0cW2HgV1/YptAy5x7IpBVGVPozS2
/MVgM33m4zc89t/3uEbirnSUghdxUNchlnOH9Mf5cE2kCLhyMtNVsfdL8MJMFdJS
Pw8nodW6CcO+4AaW3kCN9aDfXNCFBGm96i+anEwc1D1oClDV47jlrf0/E60ZLSel
SGKoaxPzDoGlGPkZWyZfSWBvAnY60kPCLp9KpmC3peioapCNuApkb2ds5wNDyzwv
bgwA4I2MIx2aybG6wsqtBbR0kl+RhtBFgBaKpDmOAbUDaYq+128phsr5XDMQAA6m
s40u+yc5Zt83XXvgpmBrA2k1sszLC275f5u69R+9Sbj50T8XXFGMxou2/gqRn/s+
pku21UoCo9OP/LmoqWUNdvfSWz/DzT1xAMmum4UTWURpBV0C0M+MdUAxFV8b4QiE
I/wFLtW1oYC4fYDFrEln0C8Z1i1fqe5V1U7HPgKc8vbyqKKrelZM7F5pBlayeX1K
WX40YiU/xlWjf6if/rhL0580NMbZi7y6SGU/HyY28MoSpAIqC+1BXHSfWQ5G9KZ5
w2g0vx2WP8L7uerPcIUkuV2FWidb9Cg56TRxYfQ1OCrkThXzmLhM/FUiZQFGskQ5
YrCCeBeHMCeoJXHYDqmfVnHT5dgYLdPiKnub2nI3D1MMmjtMuStfcyjwQHNds21I
Lk1JNSRWetzLbGA7A5WaB4QiX14fF/KhUIybsyGaxFZR56trOzSsXyD7JRAXhW5f
yswLyGeCV0LgtPozXRhSLmPAHNCAkigFPNokuozgv5N6ISGWnre09csOf6CTMshL
fL0hEXJssfdmrJ/VArUaL+jeqTfe8nMjjs1JaDf6mbPPnZqv7uloORRtOHCDDSrE
5qRbEQdhKgbBjsuwuvelq1Fbjm1p9wCF/TGZhL5wlgIg1LuPAuwdgHG3wIqZo2Gk
Bt4ng0OlmmrvY12hDz3TwSB6wxtRITOXS+0u+iQ1/UMTu04U1tYCr1g9ST617YAf
UVoAcylB4xYMzlil0PHApJy8R6ROPkFyiiaeTNo4knqrnzUkqL8pFyXtRLwVUrPu
iTc1LIjzXAhd59qtj0ToIPLOU/X1AcQNDKK6Ep8qlgYfXYdLJ0fB/6I64N3tkPyL
uqoigZquvUIKp/ny49UzHXhtlNgj6phGe7Mp9+hca5/DpRnG5P7923Eux/bZIFIM
xWgxxn8NcVHsZgRTq1YBvkEeytwp/RrJxsZTeJXRNmEyDJA93DClkYd/4uJDNhgm
q8sCZZWDtrNR56jVskThj+aToxjyxKi5I9HYQjL7IaFUGmr8xBSleCbGdJJwTqHo
oiPIcsRx/niOoyb3utdcpwpan7si48HF8AksF7LlTm9bfXPgVEl3LHwac/SLGj+P
oXLj8OMXbXVAHN+d+qr6JdtcKExg5pq860XfYAVqdKWG1oEDiYYEx3CkQvAxNB/2
fFGGnBsnRAs+9LwLUibDVTXHGMEj5E+Ruy/wKtE0GQMSznbAL6PsidiVxFQPCivy
c84oDBgY3VBH4TD/OZwMdY4zoZrGZb8o54B78gTzCKuPT2dZdzKz5Vn3ZxBc4X/J
+FWBlUQUl/vYh63Z7WZejfhHbtaLanklZi5rldIVMK6nfMrXLGrNR2ORXzk6I++L
2prND6yT4Ygjhd0Rm0B8+WZocMo/3a0QG3jwbEQXy7yIcYLAg040WoFrjDdcQkOy
QDGL0QtYcQRizBpe38tc0bRJ1AW1QwS3j51WDDBZCrsKcWBwVvH4iMspjlJXQSo3
0clgpWJBd0CLjnlUZNcy8E2aEAbwQPyDLLSne+8ZILkO7gxg1CF1T2/kIoMZBSH/
52hGO+YNPbF04wv4a+dXdzmpeV5hIJNCG6MvAdL9O+Fff6OVu44Y7JlF4UjhFmSe
doD1Qp0PTX+6YHck5H5toOfnIQWiqpUye4jTXB2Z4h2yUQKLx5Ak0+eTKi1XVaRF
HB4RD/kLfDb+wtQEs1CK6qzRzSyWeWisWAiMwOtiB5nW1Ju9zrTpcGJynEo/xBSU
1qtcgrEkwGYcPj70aR9oUTx3N6sBfI9wqAdaP+ygIGOh6YX+dyhHw8X9oD9v6uNM
Nl526xJ0Gs2Gp9MZqKfjFtXt5eZ+j8v2OFNqV3rPubS9M+tCJBymofexBKDXbteH
Z3CQ7KbsGmpEj8A2mrR53iJKJHefnVqXEXcTlfOFz2y54uRkQfnWT/1h41aJMi5+
3jnWJnuMITTSJXjYbyG6qHOJUY86N/5/wC3ToVH3u+LP+oOZ9QvZUX3Nrle5Y8sY
ZFmVAw6jtTWQNKbatVdO/26D+AQ6Uwa4vk2O/xKcrECaW6hXtMfUbubOxeDQgC9y
z3zxzqSYx7ue527K3nc2SAD83NLob8tKCIaTWO3wxb70NHrmAlvtwgwmzW/yvZFh
GVd/FYVmE6xr4SYBcJnkdd0+x+8jgrgwuBAfmkT3FaHG3kO47JRBCNRu5Zad2qh6
2HW+pxqbWCTftULj+wA0Xee1bpFnbZadyVevkHOB1sz+bWUjWGxFktdy7iXgUsgE
KDw+gQFKaCoXKvDcHtrfmvwadlei0g2F4pHXNlSYJusM3HgvCVoufP6wbaQojp07
IdvxofmVpKSwVMgBhedWd6oZLFPFSMFmUsd8xe8sADHMUQ1s8JN4FWjFux0pEv9Y
tedH8qm+taEtmxMKr20BIRTIR/stPKRoi4NH0qEljTSKGsA8o6crJ5f+9hldAJo4
PEwmoL/dZ28XQ0KMJIGTU7EkWzVY7RJ9NwL4EHefv/Is57lLUUXcjUC7AqqvH7IU
aQA43zSBKvhuzBpjM95nE7ccHNU3a73iZUpOV9s5mPoP7k2+P5aqXFD71KmaGVdi
yXz/BDG10WMWEwxcrj2kLR6LUcVkoxv8yXYkKKIfp7u8E73ygvlp8Ll663/q0lo7
VWhARQTrKqz4ha0Ve6xOefhMkH6ZO040pD7Pn1dEnFGkzPcMZ2vJaaYfLzH0KKoE
K2+YZzxDHIFa5NqlxfgrqZW0oX2Unt+UH5EuHefw5uAXO2VrqNVgtc9E39cWbU4h
pxgcPQ3cY6CkrsHvpWj1q0pHio2NH5ao+t01Zbbty7c=
`pragma protect end_protected
