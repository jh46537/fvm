��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���ጨ��K��q	c���1�hW���B�C8q��O�jT7fp`#�X���&g���lI�G���r�f�;cS�%�p�А���Kp�>�'9��8(,%� �O����	T��8�e��z��u�		0:�(y�� I�h�}�Q��t���B���w,_�����.����� Tg\[9$y�kۡSD;���.�jT6���[��Ʌ�/�?H�/ ae�� *|�=�Y	Y���i�I�5ܾC�	M���DD�v�ǩ��9p��gU�vӠW"�l*07�쉠�a׋g�[�,����x9<6�G��R�<y$�V;I�K.����~�m^'�����վ:��T�gm��d(G ���`��ˍ��]z�t�Z-�K�A���k���D�('P��i���KX�U
���c [�'�ﴣV��T.rTe����bdQ�PS���u��8l�R��Oޫ$d%�/Y�����d1KgntOlV�Ƨ�8��D�X�cޕlx��([L@{���q`pU6E��*J��t�c��3����6<�t_s�g�j�ܰ"������� dh�����i���0�	Zȑ��Bj{6�9k{�~�ra��B�@�J�jKT,��A�S+	
:P?];m'��Tc'��2�F��
%H���f�~��2�z��=j��V-M��ۤ_�֒M>֢xI"ɅI�,�F�Ê�H�9�i��/�K�Ms7#=�
��2O(n&�T��5S��k�DS����;߼x����I4��~cǽ�������8`�� ��d�a>X�e����Jd���[�PO�x+@��[�~�	�׳�ֻ��"�� ��9�+ZE�������Y]Ѱ]朼��O�Uw�Q�(�����{& �t<�a$E�]7��( c-�,���H�7���d����9bs9����R��
B5�#)��M�x7H�]��ʴ�3��������J���W�0�����ep.�����]�E�P�͖��1U��#c��d��͙���v�bU���AE� aӨ��48�I�ºU�;RGxd�٫5iU��0���⟭[g�ݴ�P�T�L*�WM���`�������Q�e~
�i|mQ�JH3{Wl�5�[���$u�8�D�AXB'vxx8���ߓ!�~g3�9W���fv3�,��̍kd/`k33�E��m��U�%պ�{�e�u ��ʞ�$�1h�r�G��W`�#.D��+���B��m[<�>Z�H(��,$�nJ��c�9h��=�������^�unR��������0�ڌ%�����;�/�u'�P�G�	K����ʐ���u:�����s.G$�Z4}��1&ϣ�f�/cp����5-Lʇ�u�|�#z��̷�������ki1���L����;��o\m �cЬ̲�#T���F��#���Æd3�,��V�j�!q��&�'��v���i�*]����	\m̓��+���<��$a(�/{�ʯk�<)(��͔+E���J[bߙ̞��'#�~[#�qsFF�\:3:`�܏8�4��oP]dk
��m*g�'"u
����͆��}W�
���(�~�BO7�sX���QKok@�ګg5�H����"�1n�����uFS�a|��D�y�%�79�#� X����|i��ѩҜ�Ω �i=�"]o��l@�n
�v�1��LW
Ud"����/UPj�R��S���x�J��r���u*4��F=W#�RJT%�W5�0�?�C
t\�VB��p�S�ZΏ�ǿURc�Ȫx�WmG��NPq~Q|/SZ��q5�	_�f�l���nzޱ��>��S�'r> ^~o� ��5E�r-��J�g+���X��k̏���8����<$폢b���[%����#�s����NY����hM�cSI%�����G�rj^�V��A�}��V�qS��H;���s؋ܚ�],��Y���M��+�HGL[q�Z���4���H3��໱���<$
�k�;G��Ͼ:P;�ko���L(��ǽ19̯v��,0�cd��}7��E���e�w2���2v�����6(�u�R	?��Ֆ$[NX�{����+��c`�Dw���.����p���)��2��Q�8�e��3E�	m؝))f5N\Mx�,�ΩE��O_X�<C�ݐ��'�U;s��sZ�M������Ȋ��;:�^���a=�$˕��6��zx�s��0���'�Nb�zk��P�}B{�����������1m�H�fҏ2�?����Z��a�V݂n�zY� ���n0�|�}���Ǿ؝�E@[t2�]�8�!����~km�Ϯ���\�p�V~�#" � �[Af2��%T�0KZZ�V�r�՜��㢕P#�j��v�������"��N�6Fog��7�Q����d�9L�
�i�I`*H|�����}`�ЦK;��� �4l��;P���DGՅ�U��v�xus��"P�xڀiv��A>�wz����6������d�g���`&�WNȝ2��г���]d s�F�G���
��Hc�~�z����j􃢪��s�:��Or#*��­�hb�\7ރA�!�Х�|��hE�^}|`v9�g���,��$�����MWP���
q,J*���p�����3�Q61��P�ʛ<�/P?c���#\���`��%=瀓�2����V������Q��I�8��Ɓ\F�<	��<�����I�%VtF�Z��۶�����1Щ{^��!���{��������Ft8l��^M1d#KA�eE��3�/P�L���fJ!)er�/OO��I+�(;u7>��(Y���0ȃ]	��y���')��I��Vy
�פO�'1������[�}��]J�N ���7�'Q�Hץ��ől�@d���,�c�J��ݤK�K��S:���',��O�;d�H��VMbK��``J�ga~#R��px��\L�圁RY�ߤ	��1��6X�.7���0��c�%%�F��t���rU*�C7�3qu�"�P�7�U�Q��nΈ˧���v�T&� =rM�V{�#����9���,yf�ޱ�s����s��i��u{"�Pl���>{nOo�{48S��]Z��9��+���R���H	~w'�R2����F���2y�0Q}|�_U޴�ni͝	o�5a¢x���K,w��˒�(�n���fp	Q	�ف�6�,�Ѿñ�Ǥ�i�F���r�Y.���J*�<��nR�ג�.�N�u�!&q� 1L'����zLw��^xp��]QtQ�
����C��O�C�8A6�/�*��oL*/[59�M���w|5��}��BQ�Fm��~?R�� �����=~${��g-�)MU_k�>��-.9�	��g+����®u5��#n��&�]���۷�s�X�`��h�CŲ�/[ %(6�C/[b����l�n��Nа�Z癒�8�{�i��ݫ��=�S%��	P���V1���̹�
<!��\��4a!H�'�Ro�|}dE�69"�5V�#��],�Y��B���:��4�z�Ah����.�*Dh��<������a�{&R�$�e�?�hr�fB�(:�O��\����м���P�^P��f;�$�����Qf!�1
	gOݟ���'���cO���;`^őrq����Dֺ���B����&��ޟ&.�Ƣ3^r���`�Y�Ifil$d}Α�E���y�����O����r�s����R;h�L:IK�[�S˕c�ŭ]��v�&s]H�J�)���.����7�VC�� Lې��cU_�Rb�"��*V2�]�t�!M[�M����������EH��a��U
)�u�a�ʭh+iz ���p�:���E�e�&e�欪`�u��8s���t���>Nm
O�a	;�9|�n8n��c\��������5�� ϝ���=��4]s\W�r�������7#�i!�H��L��w@*�������t�8��8��x���ZY�[�������D�,4؞d��J��2p���l����jWz���5��j-�¨�,��L�Z躬�|�|"�����"`lRH�	��r�z���Ow*y&��R�>�� �rF:.G�\�$�;�֞6���J�J�،��[����O���>~`½�ɂ����j��H�
7�"�:yy���e�i>���U�W!��l=q�Vb����c����� �a�4p�_^�Z����`
&<�Mg��O��)0~�EŪ��ک�%�*
��lC<��$��&��
�6�eA>������B3��>�B�X�����"���ƣ}��;=u�*��Xg
D�.�
�e
���_�>c�f��{H��hQ���d����H�07*7��~���!��i�� 6uF/��s�?]���oZw��7l��B�R��m�~����G�jk@w��	\X�#���?&�äx9;�`]����%cr;?t;蹜��ϕ"M���=z6in� �1%=/#���;���.R-캧��V����iF�π}P@�ơ�{~�H�d!>Cu�Rw���~��>��;̒��G��r�3 &7�gw��χ 4��
$>z��I?��X�u�1�Q��J1�[��w���X!�*Yi�)*��f�;ʏ���c��R条[S?�Fzh���=Y�@�ig}3�F�Qv4�,�g�����7 �u�jI��9������M�<]:::�@�M�j\{�Ob��~`�[,"#�����Y�����L�7!(�\��i����_w>��̿_5�c�Nu8�C.᜽�oAR�\x�#Sa��z�Ǥ���l���Κ;����t��b�:1�{�G`eE���O{FF0R$�e�E$R����o@�� ����\�g�Wǯ��j��{܍:ɬ�l�:yZ �e5�၄C��c�[���D��N��Q�Q�+��^�V�I�]�Ҟ.>7/�}K|���]R�Md~ib�*V0'!e%�2���e4��Ww��������㋖>�01e�^\��0��mp{>1���"��m��B>��W�S�-!B�k��-����D��?(c�6gڦGf�$�tI���mQD�"�6{�+�O�����1q�~��K�(�W�I��ě.�ʥ�Y�����4��C���D���#CpUq��)�C�w����gln4�A���&L}U.����'�����8E�5ҡ+?sP��d~;b���Ǭ�����&K/h�7�EU�:��!RA7%j
��]B�7��M��"5m��TjXԦ��8�H���Ǡp�ٞ�&'��<*!�N.��K8��g�7��y]��$�C$���T�4����5�Ӳ����oO?mi���̘�E�I�H��^$�K��	~�+��S"Y�..{dƼ*�02)a��U�u��׿�c��kR�-6a
	$N������_L�&	p��̋���F�������N���7�U>{y-L���d��h�Z,�8����nj��`���FڜXz�߲ԉ���?�.'��i��{2^�{�U����,��C�z��ɹc����c������>Y���{*#t=����&�zY��FĨp&ڠ�/:/��Lj��hn�_7ꦪ�M۪��Z_�=��!����%b-��[��>�k�.�"�{��K#�7��A��
�)W]_�����81� {�jY�70G�������N�^��z* �"#]c>�X?nգ�q\��%���
~9��D�Ќ:��+!`W��sQtoL�,Plo�L[�<K餼��[�Ʊ�X��	dh#�e+�����;��OW�^��T9V�]=9����F�C��
1�EG�����?���^�R�fM��{���ݪa��Y�ʻ��ZÚb������WR��О*��V��GͳL�-
���yî3Ak�:b�%�	H�e�tb�C�P�0it�A���1~&�v��@���Es ,���Y�@5ĜҎ�WOD�6�%ӝ$����	�75�Ȯ��������4��^u�(g�0�xjL2�P%=�5�]�)�� �D��t�}}i���h����	�V7g	,�ﱄ_D�AY�FM	��1Z�'�4�E�Q�B�$,2�;�D���9-�B٦�O=��Yǳ����~i����JOQ7� =�7�g�����y�X*3�ޓ�W,b"mGv�b �kɢЧ���x��'W���oF;a0��-��8�֎R|JG�M���~�+���Gj3�⪜)��L�IbC�V�U��7�\ :�����h��Mv�)���9�{��o �� Z�E�>�n��f�;�ƴ�}�4�8�}F�t���rAԙN�؟Z��j�{��'k�v��d�����(�s�L�D��<"��U�
����������}��I�脬	�����/�'��ܔ��H����9ߔ�F�
�W����B�\3ܩQaS���#�4"�.'Ph�8'۾v��=�H�A|Q�~?*�a�{��36�&/�8�������=��%IҎ�����<!�0�R:o�+)�\i�@&l����C�Y?�̎J	������l�>BD�5z
�r]D]�~����:��	늲�I�~��F��Z�o��`@����N��+b(���Fq���І�Mت^,��=�g�?j�)��嬰�4��"�$
��t��-�����3b�������^�l�W*�;��r�ޅ�kߤ���Fx��;w�dRop�(�&ӆA��Rk��R�w�N#(ca����NA�V`F���/	7_YYB#��A� x���6u!vDO���v�(�'b��v8����G�x���P�	�9!������#�ޢ]og�b��_I�o2���F7�"3YȬ�q�p���ucFX���s� ���m���r����K����ZW������W ��r74%�c����@���f`��}�k���{S.����>�sw؀c��<u^-(2�Q�u�
i�V��{�t��W�a�W�����$������ ������둄��<ݓ(�Gr-�P�����;4np��&�k�����z�*���$-
��u_E,#�'�Nu�"넪pG$�����΀N��a����H2�\=��� `D����GE���'}������U�=i� �2>	ϔqm5�����I���p��ϋ�^��F����-�M.��:CoFQ3Cn�U�Zy�|C�M����팍@0�m[���L$}�&!�U8����p�@Z�y7au �	��aҞ\a�֚���q�Y�#�G*���u+�w��g=D�>	��H0 `N��1ʬ��?�\� h"#Hݫ�
�tjd�� C�bd��w���'�^*��
ե�f�(�ù��9,�8��d����@Ǌ�+�:\�F�W�o��u�Q~!�3�3�p�#Ο�
��y$Yb_�U��q�.����H� ��2^��-q�xX��������v��ཛ�� E_�B���2<�E�M�Q/p]$��\��x ֗�����C��5�:D-�3r㚨!Z��j4T�����9��G<ѯ�X�U\�Q|8u��e��Q}��&.����»����9��(�����@��Z�<H�:U��!ۑ&�"7��=�G%#��`����}Ft(�����x�5�%d昀xq�4mMn؂4��,$��FR-�T���h&�#2頻ܬ�߽����t6h��J�o񠄠hJ� �YM���W0�%!�RK?�����"�ߙp�7�SK�Ԥ/�#�]�����Q?Dd[Ĕ���d�g�S�C�)���F�Si*o\��2��Q�?�a��d]?�P3f��Z �(Z�̕5��!Q�} �.}�@C��i�<���HL��.Q�'��$��>jhZ3<�ѣ7�ENG�v�1�ש;�z�Z%�-�`)o|0[^W#�%͑P�>|V }Rq~XU�X!V����Le�����s�E*�^r�k��nkY�p/%�e��#��m�Bڛ�0��X�?�w�0���ؔ�|*vu=�m��B��C-�l�5����Kf�
��_L��W�k�5���޷'�0֦IwV)/�XPKD�Q�M{� v�ѝ*uRyI�W(p.�e�����?����H���v��p��qxy&�?z���2�{5��;�]+HP�j,��[��S3�diE�k�ZA���%��S<o�x؈���OG���q��Cg������	.��Z���9�cy9��ڦ=��7�����m������m	��	�H�M����&��Z� ��B�)�EC�:4�D���!7��`7�hH�I.oK���/rc7⩅�����0^����� {�,������n������߼��N��i��Dh�WN��
H7�:Gn��6��va8�'���ŋ3��j����lj�%B~�����4���C7��F�����i�h���
��(�p�!<y�5�xa{�}����j%o8Y	/)��q��^�KzC���m�!���:m�~@�k������L�a�Q���Hj��iUg�G�<��p�@�k��w���}�;�C�U�=��H��ZT](��U�B	R�J/�z�m/��n:�O�Nb��6�
R\]&�`�h��=@!��b4)o�T��J9B��ɎV(��*�.�~�\��.�&�.�BP�$�����nb5z
����dfIh�¦f<#/Q��ʾ�AI�(4���f� 
�A�Y[�����WPj���įsFk%�1o5�~vI>��,-
)��cO��m��ĭn�A�/_z���ɟ�.��V���E�&�[kv.y�AUE�>����J�oe���m8J��݉�+e���ʌ~j|�%��>ܢ�r��m	�2$���1�D y{U<�-��i��8�d=F�!(~�Gp+��מm:ܩ�d�-�'���#������S;�(H\��s�����+�����cү�ל(axo��G���Gd�>��C	��>��}�]�Dl�_�m�u/6��-M�'c������$I��3���d�W�G��;nm��-0%�ݍ�C
4��$�Px��م+�@ְ�t�ٵ�w
�ͷ��O�ƨ�>�mLB�9�J���vOT���F�������^�M3�ϧ�n�����G�]v������c���[���L�����Y��}�B�F^���U�/q(����Ώ� �˕lE{H�xaĊx�ʹ?^�����|�n�-8��,?ix�Q㥛�a��׬i*��{d��	�OE��݋0�xF%�^�%#�kѭ����U�Y��'��҈�?�r͑H��[�E�ҟ�:;R��l�H�X�?�h:ŮVڽ|Y��0W��E,R1��2-��rn���uQO ��z:�!۱<S�������ӢQ�H��q<�L��z"@rX[+����؆G��N���喅O�	�e�ЭloA����V}� $�]��l�Cc�X!sX>�J�@��U�9�_`Gm���7�2x�46�z9v���w^1s��� AK����CĮk~��P):�-�I��A��PD�B)�D��TԼiqBㅂ�3D��������*�>3��8U�样(DE	]u0#D�C��x����66��F^�/ގ
�P�$�јx;��nRm���y)�(�~P 7}a�j�U�3�/,e�0	r�E�A��H*k����Q�+�a��J��
�@~gU�~����SL���giCֲ�|cn��`_���D��2��^|�H�ü7�I�L�g,�I ��4C����zP}�Բd��B��l�dHG �դ.��,N�ę_Xn[����D<�^o�!Hh1�{�I?�$�]�Q��L�!�9BU7���_��2f2��.���.���EG��?nb�=�9'S��]m�#�']/�o�.��o������Su%������X��aZ�H�OZ}�=p+[� �����*Q�Z��T�w>�ʤx����{;�����>2�v�.l�c�*�I]��I�S���q?��flrX? R�SU����ɩF�B��]�E����y��ut���Գ~�k7|��+�o����;�����m�i$p�r�X��b2�=��#W@l�m��q�R����KҦS�y6Gq�?���{��<S����u����rz��$��X��"��Lf��j�����P2�f�:���5����TO�C����st`X���>�R� Y8	�VRS�����)�!5Ae��>����vf�m��H�-|C��,�٭�^A6�B�nG����§��j|բC�Wfč�%���Ǘ�u4��w��8�����k�/��Ї�Azp:�%Z���������祃5��{�
u�H�YN��e��M��
��{R�9�x����-�v=ͬ\�C�Xq}�8�o,�HJ2չ�qю/أ|@~��X��	E��&`�����0��RZ�� �k��Y0c�3�V,/��:y�In�hi!��29�3�:�mP�p��bR 5ݍ�/f\p�tM�/��|Aױ�4��M�*P{�q���t+���^)��q���>��`_hbu��Ȣ.Ǭ�!����S%V��`d[�j�"DR����M"MD�H��@�J:":���)P�������]��q'���6ECo�]�����:6ޣЀWX'N�/5����Q�2#��	���к]���@�u��!���I�x�f����ߟ�7��G֭ti��@��K��Z�\��2���Sm�
��_��/{�e!��*�u>/�\��$%&?��Dc��%��ԁ����E|<�c["J�m�Ut;�gÕg�;S�WI�#r*�ty

4L�/�����ON��)�Af�z7k���]ϜgK�����Df� ҅.G漆�ϫX�x��߳ &���+fS�9��O�i{J��i����C�}�BNO!�V�sa��c8�2�y�'>��:�3 	���z5��</�{��Lr 1ڡ.�����?���3��r�vO�t�(s8P'u���ڿ�3�@]��8�S�.O�F���n����4��-M" :~��h
G�u���\�`��{�����2�2��C�M�,����A��0��k���\��۶�$��/zu�D���,����Տ��a�����R�xփ���?��'���i͢5M�1��r��Ґ6�{�ma�;A�9�E<O��@0=1J���M��ϻBU^��_��ĝ��j�`ȉ!���y�	p��ta
2�gi|�`o\+C|=%��`'X;K��1T��ǐ����?A2�Ш�>�@���1d�j��u��U�"�F�e�A�,�h_~>��?r	a@����^�U�ňs�1@��<Ȏ婈zB�mQ�m�_�x_t�~�n2�Y�.��>�@T��C�!���
�?�W������Cjj�04�p�d�DN���Upo=�����c�3��YpF���C�gG�a�����=�O;p���r���h�LȻ�Wg����D|�ٌ�=�P�}�g~/�@(�	��e��Z�kp㴩(V�^h(�Iq1TWsD���nܡU��HQD>�2�Ty�p�4b�lsRp��w�9|�i\RM{����I�7P��6��	�p�O�������Ĉ��5�K�5RȿL,9����G�:��3��M���$��o�?�nV�->� V����
�-¹��O�j��,�ȥ~��Q_P�;� ]�P��`q+�r��Y��U�`����j(�}x�wɳ_� `�uq�I��J?qI��>>��7��GwZ@��V����aV���½�gp5�S����-4p�'r��^����R����c��t+;�݋;.�}�o�P>$A�OAu���E�^C�fQN��	C%d����m�����-���w�o!�`���1���m;�ez;��&\_j�H͐6����J�w.�B���^����v������ ��,��-[��#�:;"�.���@�iJ>H���
����W̛�s-���#�23[�/�8��ʩ��[篖�j�Vt��Eo�$���<���d�E�t�2{l��f��Kԝ=�@o"�l�A�R�	J��]�.7�ъ�V��s�9	$�lSQ�U�gԖ�ǧ㮉��R<a8Q��c��#���X�n�g`�+�fͫ�W�j7]�[ĩ�1��c	e3������*M(��U��ze���
|r��a���_V��xv�j2ue��2�S9P����Hk|M}�{=d��Џ�O�������`��ImN���T�����MI���ʷ��Y�_慪~ˏ�Wv��;M�@2��T	��Z�v��|������h_|؋|��XD-Q����03�^�V:�	��<��<�[��>8��5{ѭ�r#������n��+��!cЅ�q��'/�C���$4m���>�M.�L
�e� �51��3�8��ߡM�Q��5*���@A>eeJ����{��c���|K���o�4y��?g�k{�DP�7�@�b�kV`MÊd}�m�xc2��L?��*��(A/6/0)�)y?�ZH�[rܭ�����˔��� ?mH�ER.3�QGJ����M� 6�I�#�Ž��(�'W�=?#gL$U�o�]Rq�Z43���8�k�9đ^��}~�w���t�����[�|ƸE��$���1��Һ�O�Ny�u�����l����C�fY���!<�3�~��P�$^��� ��"iY��������͐��DP3�W�b#�"�a�b��1-��>��[���^��s��٤���m�0�bdqW�G�ֳ�JAݸ{�۷W���C%�gG�)To^�rG��`����.��1�T3�s���}^��W����8��=��h�Qw /�!0UV@b۹G.�1��1����I�wB���sݞ��Sf���l`�/�0���z9��,�����.^f��ڪ�E*aQ���4}q=�O��ɸ��1p+B���g����PL�D�T�EG!���rC����zecW|]m}�`�`H����x~���f?�Dd���$
���B�#��>=�s�̦���gɿ���x��aɽ�J�@��b(��)}�	��B
@�m<2�7ʘeup5�r�Bu�0�t��ߘ8xH�|G��5�6�T@:��}c�Z�B+����\J�!v�#i$ȑ�^�A�#ry����~�?�ʫ�)�]
���F~������zan@2����r��9#ժ�J��٥��5�
չ[x���{QB��o�S�����L����6���St+IwU:�'��4PLW�
-t�����.����7uJK׎i��e��L-�"<���#����hNU#����(E9b�XO��q��YY!YM)��7����?�ů�f���yBw>�y)�j�~�dL�NA�^%2�N��Rz�%z4�nQ��U����J�����9��2
��t�������6 6�J�+1�g��`5�0�K���I��yC�݊���g� �T�r��L�f���CUK7�c C��
���?�9#ro��"bɹ�Ҡ�;��,�d�y�5�^�0��ˀ1fn�P�T�Ⴄ<y t�l�7���9��?�*������.��pv���q;f�1�}�+��T�c�"�9 1�j��|��B�B��ݲ�WX�>��8�,S��P�m�z>�����0uW/�"?�xYދ�n���S�l�jPFe���#�T�b��ߑ�4]%�M䋑�$0$\�eN�X�O�Y.L�[����st���K���?[�;�QW$PG(;ku͛
�٩X,4(g]ɝ5�#/f�����
�I~ݦ�b��׮y&��FS�2_lI�C����:0C�{: ���>|��e���W�6��#��"��Q���A>#�Z��Dn�g��Kr��b�P��P�,��݉2B�
�`����s�9@D%�b7uQ��b][/B�$'r�v�b4:�-��z��'|gs����.�e�H�� b�"+����X�ţ�zo��D����T�E~/vT,
�ݤ?2�9�9ԹXuf�~ϟpedPI�j{��[���DŢ�����X��x/�2z:)�9jo�th�1Kc%z#J���A��ɛ�:��@N��I�^�O6��136$ι�j,W_\mg��������թ,{�̐��ADg=�n(WqG}O��%>����_YU�m���0�L�W*�	�/��<Ƕ��HK�1$I'�K_a�?����q:��S�k`��K��/�ڑ���[����^�j��>�s��
y�"�-k�#	9�')�
3-�ɮ��s45�52��L#ID����S�.���Y@�h�l�ͩ)��)��¤l�Ԣ�L�`�)b�E%����Yr�J�r��׏K۸s��eQޏ%)�o������?��oو�ٚ}��T�cۦ#��NV�Ͱ��MG���JX��D6�	��Ba���;Z[�}N/��Z�߱��}���,]_M���Ss=JÍT���&���e�[+c3m��E_v�Q�d�P�>�>JN�Ifo�[�C��ѐ����؛�ߏ��-WK�G���AX��jmc�zX/x^����q���t.�2�)އ��uY=(�z�k�ɮ5�+G3�x����#X0�(	��v�;���!s�B�e`�����>$O�#-eo�f�:`���&��Z��	G�UwZ���O.����\=���ߔ�u^Fjey��h�j`=f�fkT��.��ωv�^҈ʧ��%�l%�!�8D��oM� ?h�$(��z0(xC�Y�C��JS�A�����_�A���3i����s���/h"���I���Q�׺�� Q����K{���&��`���$�c�}l�kq8�b�cYU�}���P V��c
�;;x.F�L��Gmtk#s;���$n9K���O0vta|��¿���+i h0��8�_w6�G/��Mn��z!/"r�`{�Ng%��Ye�F�������5Z�m*���	�M.75�tx
�C$��B�Y|Xv==�̱z~d:P�*	����K�����ܨt�vM�/)x'��������er�p�wȅ�pNd�[K����dX�b)�W�_)�T~��a��Mo���$�]��0,�A���}��ǆ0����d���IW�ʥ���f�Z�6�'��G�,� G)�����ɇ�NUwwS,��n5tXPz�'Qn#��Eq�j�ny�
(�Y:��H>�� ^M�b$�Ê����M#��0 G���)_��^�������@ɩ>j����8Q>��|�[����VF�L~\w�P�z�<�!s3���o?�ǗR�N}�Hh���w+2����l��n1%������A��w���Gb돺~���2���S��6�<sr�a���&7�����˧�x}!��th\wZ�W��R5���}���-�z0�,7m����<'��>��S	��^vC��b%8�p���nt�ǹ3~y"7�^�����l�!����C[^�<ec��W���:V�0��i{ONYV��ɯ���{��k�T��w��n��-�P�4LH��PE|�L��a�n����rBz��&��,��A]l)��<�Q��d�dE�m+���&F�:�Wk��eZ���]ؑ��}�I�-듧��TѰ/qmX"{����1>��SvM��j�XI=t0�s�f!�W<���Z����(��,�`]��˜��4b�O7�@,�l>1'�$�%8��Cs%0J&��\��&Km2��B�L~��j	B���Wpq:�)��|9�%+��K�)���A��3��|g����Q��t��l͡����]Ⱦ�ϭP���d��:K�3/�5���5pN*��s��B��$�q3GW]���?�5�6m(ڇ��w�u�.�;G�rK��0HXk$k� A�e!%�Mo��C�,L��NJe�U\��ڏC5�Uy���ĭXR'�@i��~q�p6"�X�p)c�{�հ�D�G�U���'�����Tv�cY�����I�g\D9.�`_e������Z~LY�r���X�߯��dܻ�vJ'��Dˀ(UejZ�\�|y,��(��;hDs�*j��,�uus}��hZj(7�}�|�O����-ݡǳ�c��L�z[���S�H?��%�Dv_�G�k x��/!S�{�1�\���ȹ�)m�ZU�e�	L�<=��)���v��Hm�&��>�ؤT+��9�P���+����A���Ѭ�a۸;%m���9��4*��-ݭ(h3��D�>Z� �~�b�ڿ�u�9IM�~$�-b��$�dTZR쬓����s�ʹzs�����I�w�M���n��?}���qóX+���
�$��_��������1�ag� ����ӲU �<��TnG��3`=?G�z��%��_��.gR��I�*��|�ft�8����T��c���K��~fe��e��OV!w1�*u{M�wH͆�^G���>�2�$�=�az�ט	z��B��6��i(���ƺό���5��n��"bDdA�-���S<M@c�͖����y�6�$�c�~WvEN�Ye F�#��{h1��]�K2�3�5�"e�l	-�Wf�@?X��e�jwŕ� �銟'\�+��|Dсh��Q������!C�If(�����b�Z]�q�5�`�g�9�@���<^�'�V�n�HO�6T&o��hb#��&��b[�;/_I��꾎Q�*��]f�{wh��FM͵l)���ο {H�;����_��E�:L�k|/�٘3���z��}��I>J�S�M��X�EE!I�X�4Ձ0u���.�\�`��G�^yk�#���BUz�C��^�{��+;��z�@�Z��j�մQ*���2�.b�<wm	��Z�BN�D����x�-�xb��yc^Q`m��)���#�N�ד��e�w��Ȃr�	�ʷ�����;��O�gTbI�m�9����s@��:�ۅl`:�����8�.8K��֨��,H�q����-@K�ø�g��}i�KH]�UC�4h���v�%�*��%�&��2���6X��=J;cæ��9��-�<`�S^�S�:3��~�W��>����&e�%����H<+L�A�񁰱���I8�J␺����_����_O@�8���!D���VcR�n=4���,\f���b_4?���A�����t���6a�]$+$�ZZ��O��rd��PW.F��^�\��{NT��\B�C�9$M.W�w��������&�^�7�J�q�W	�}4f9-�=͓���Tx���"�↶{XH�h��d)دO�B&��X�qZI�E�1e���<�d���j^�~��ȣn��hyK.�}�Ѱ� ��~h9=K���z�ο���9B��tB�r�ހ�"T�V!5x�R�N�C��̻HϲM}�'_?ړue{�M��{��{s��-7?�<G��j����ӳ���d��V[�-1��8��7E�h�Vр�%�멗K��ޖ���Ϯ�0j�s�= �R�Z ���$H5��3v��a6'��/��;�D��q�J'5���l�^�!;S�[.M)�Ksb��{��~I�z�>��)��\D3���Sr�[�rP�,:5���H�H���̚�ɪ�7%��fA�����̭� ��+�H� %�5�`�^6�F��M�B��IC=���M�����}D0E����_���g�� �#�����T�,%�&�J��+`/'U���X�Y��ٻf���Z�k��R��/�V�E��}���b����>1$�
��!D�jA�A������d�dy�O��	i4��Na�cz8I>#C�⧳�T2cܦ�v����(j�sW�:���3�p�Ws��O�N&$}�9��^7�_�
��n�
�z˵�ux��TX�ʕ��E:�Q�y�2�IW/l����)�KI�gK�r;i�dl�����1��B@��[OA�����t���F�Q�1�UH�+�e}���)�7vek��j�US�Q�4�j�ԍdV1�F��	e^sv!���W�'vm�Dj�N�li!b#Ib�2N!��V���E�ݐ��� Q�?-'�o�������"~��-����8r%{c0�2�I�%�O�	o��䗨�DW�5��y��n�����>5���J��mP,� [$�4Ŝ��M���"��!6�$��s}�7�]wBP�	�x~��+��?��p���Y=db*Bl��+���'u4h��8��
��:k���4�#,��H�0qa2�SF|�����q�X3_½z��[��ӥ�ֶ,��6@ѩ�u�u��,J�+�t�b��a��"\(�*wPsC�]�Q���0�F��� �X{Ųy�"d�@��	��� Zlȗ�Y}��]+��wsl�o�M��un��
�!A����{mK��ILd�fw�L%6�VQ߹=~���rP�!��Y��� ���A��𳊣ɺ�� ��㦑�<(q�)Mi)i�V�w�V@+��|��jUO.�Z�Ę	�i�/ҫi@%�N�:�P�%�Z���/ �1d��rFL4������?�?eÃ�3:	�z(���j>GdsXf�#��.��q��
�.=��a;�JR: NL���Z=v��R�i1}]~DE�(;��|��'��w�7���Ȯ�?U��&B/��:9^]��]�w�t���ڍ����L�r�ϭS��n�8�Q��'�����-7�����_��_�A�� n�r�9�h�t^���|�ADz�>{e2G�Za��{��d��-GR|fڭ����m-��,]�T3� ��U���D��BRk^�����B�c_��<�yϑ��u-(��h.{�><-��Y�B�eV�;�5vS���eޖmfw	Ii���J�2K_#^A��U�zz�v=˜�2i������;�n��H�3�Re[���_�˳��&6�S��td�
����}JPb�.J�����՘rO+�y�s�t��Vh�=nE&�
��m�h[o�K��CM��Mr3����G ���@>	���cM�Ep�b;LDAm��4�C�X�
c4w�c�_jKa��T�
v�zB�ϗ���>��tY�*�v �љ���R�T��f):��T�y�$��i���C 2G���k%�]X� �wd<ࢩ��x�Ju�2�� S�6�IK3��ʬm�q�,y��u��}�ݜM��js|f2�7 ���>�"-�!�b[k
��
6������M��3,�{�6ӯ��cOd�|-�u���B��Du�ծ�$lC��>#��4'�y�So���Nb��>�����.��Q�����ʽ�kml�P�� ����)Xk8[:S*���J��b�� ���N�eB(`S��<V(w���lop�N��X��=���P�-�9���*�F�J}i�S�/�W�N΂Y"e���x~T��"`��Jt9��h��c��T�d�m��
���!HP�����_7U<"'�40���B�O|��%�9�ȇ�W���<��A��Cj8 ���e���j�߇ExPw���"�\��#J���6b�1��F਷��]o�84�iBdz���:W��Ga�%u[�5�Z�����6�5�:�چ� �����h�Q�	�*����{gX��},�*e�~H�T�
*��/����H�i�k�����x�i�8Y1�Y�as���Pc��H(S�����8QG���?�u�N]~�����Z\?�} Y�'��e��P�=� �aV��K����TY\K�%�@]�ӂ$e�"'�)���G%�Iqo�7���o$(��Ԓ}��q�m�5G����my��@���D�+�$@�f�;��]�wzk�����1��Z�M�P*���Xa���P
�TV�6�����o3"8����|i��V_uh}C�/vH��a�^�`��c"�Sx�=�:G%5K�p��Ε��Tk��!P�C,���l&zM4�Hw����{�~�L��D-�X�!&����w ��e��7b�/d�Y�� ��6�Xq�{a��}��T��+J%p����I4׎M�$�'��]�*~������Un�T�[��v��V�y�%�����`?���k����-dƍ���B-�mĽ-!�M�Z�?ّ���(�0���ܫj��v5�����¬�Ǌ�fA4{��h�~�_�������<�����Ф�;���;�X�68X�#���n���:H�Q�m�ʑ"���IB�������5��0��2��?�*d������k�v�a���=��+?@#T�Bma�����ET����z�uF\�
I޷/J�}ߤ�cEb�7����[��5�~I�`l�|߂��G2�b~eՈ8�n�2��0g�=����ʀ��3��	-�''$'��i�q�%;���j��׳�B�U��!��Y�������u_c�<���hw2G~ҝ?Y&/R��Fq��M^��̍�����'����G�E�Ot���i�2$����� �^����jIR��{���;�T_;ɝ�$aƑ�#~Y��f�^��lVJbX|Nf�i�6�-��+i���s�h9'%�ұhAh��/z�"z���__~�~���Rp�;L�;�[����	�Ť���3f7|pH��<i_,H�X0��!י�Zޚ�b��m��f"��8-���F��@sv��O��W l~���.�xO0�9���;�S�/�8b,u8�]n��1��]G/ �xr��"ZN�O�H��]�t�&�;�Fϛ��_0w:u��֢{�"`�{��)���Ъ�g��'��n�JX��/�.�$V��n����2���h,6�$�Um�/k;��:��AE���!�4�u=}=hL�c���ˆ���@�κ��A� -np}�/e��ҥq�^sK֠��4jZ�~���SS��nP��=�6����[����}�����8��|�l��b�:>��o�����c�S��.�4?wn4� ��R�����Sq�l�総��#����p;Ԙ7�t�8,�gᖈ�w�U��gݸ4Zd��b1wjmP�IF|ρ��i��V8����Rt��PЕ1
�$9�t�]��C�!1c�Hk��fU�r����j�o�=�G�&A>�,�f\{r�U���Ud���C�S�&Y�
9�N:'� �j�cv'���D��'�Y��[٪�g�a�����c���"9���^���JnT���w��&,���F��gY�x����!PN���p��|"�p�|/Q#�I�,Ơ^Q�(c���Xt4�9� Qa�:�B�� ����*۬HRe���_��o)[��o�صQ�3e��u�	iۺ�L}6 ������E��Zew�t��00���T�%�� �4����8�iA?�%� ���8� ��Q]҆g|n�Td��	����R6�vY��s����E<��ƁTK�r=;�C�9�݊\y�g�Nz|*�mg�~C�_Fy��Q����ƴ_1�dE\l�Ă����H��lU����-�1��Z�ҏ��vϕ�[����a����~�Fy@k>v�c�z����Q�NYG��D<ȡ�C�U�0B��7��߃�z�hX�Wb$��"/�vQ��ukX�:�h4���H�m��(���1�g�<p]��i�:͂�}����%�e��R�'�4ꄟ�x��	�)��<p�ҜT��~c�ց'���S�oo�;C�A=(2����0�N]�!���4�$���h�Ԏۜ86	L�Օk4۫6W�.v�FǡG�Q����v�#^�����[�v�!�����,�����B7�d�)��������$,ۂ�)��:�a��J��͂A���C�6��l� U�(��-[�\0����5��ENtpnxm
�N5p�a�.�^�dZ^ ��.h䙦�m����އ�����rQ3��1��Z<8R !V�hZI���?�(�3�����*���$=�4<�k����w�IEpob�_֖�q��WU�Q�ӟϠ����}�L^[��ݞ��+r�������f�0-�ڕ�k�l1~�����x[������قB��M܂�*�ƶ!�bj�&�q��eE�jʳ��S}O8<�&���8�r���z1S�⫿[0�}�E&�xe���,��u[�1D�;86�F����];ˇep�4��_i$���W� H�������k,U�G�t(�}`U6�<�A�B}�q�����.-��+Ԧ��/Sm��s���ǧ��?[=$f�Ŭ�C��FVcK֟�\��S����b�9ۏ{��ӧrl�.�b�bjy0�)m[z��s]<�[�pi����D�r/���j�WR��2�mD{r��@� ����Y��5�Ϣ((*�ٽ�2�=3�U��e.l%|�jTe
���~r�ѱ��,�k�8�AUOQ �*���Mt�/�����q��GnJ-�m�Ga��5�Ml/8��es#Wt�X���pM��D?|8	�M@L�� �L;�m5�����sD��	��ƭ̎3egA�,LL�N#zZnM^����E��ݭuy��ٔ�]KH0w��ʍaِ��St�_�3��n����"�1mY��q+�"̛T��Q�-t����l݅L���j^9E�o�\_�ݣ, 
[�_���A?� YXz�J�KC,��_6C�[K��� `�{�sbE�'y��f�^�$��Q�
4�i�����T����e(s��KA,W
�XO��f��b+�|��]n4c�i��WtR����%��+#69r��@/������"�$3�a!���t�b/͙�x��	��L�5�����/����9�k#�o7R*�;�� "��Di _=3H��I'�,�6(1�`�� J�_&]��iJ��c?�1�U����V���
�6����~�[`dh��jK�[1�㘞[)*�c����@}�⮆UG>�O.� xsE�#�-R��u�=���χ dqN�P��!��D�һ��=�0L�E�N�>,$���F��ܻ��4*K([;ɇ ��G{eG�������Ǫ��]�X]9u�;�|Gfѓ/F�ڎrL�VE�i1w��M�Ĵ��Ҵvg�Ǥ���I��!��)kǁY\�E�u��:���;�Ֆ�$|Y�$��^��ͷb��D���b6"�Y�	���ߺ��B��C��o�����j������T�'m�P1k�L.��u4}tI��#��W�>��mT~\%�@�Bp������Y��'�jt��H؅r$����|�i�"]:��Q^x���<Ձ'��i�����[hNV'3VڬT����F+T?3>�;�P��rBg��$13+Қ�&�G�v�¿��*^-(3�\g����=�(k�DS��a�7( ?hPP��9r���(�1V�8������C�G�x��o�;���eش>~j�Ѯ(<� '����Lu_^fo��-�@�ە�cr�u��vv�ퟢn���{���wg�S��I*�s�	�V��pO�ɶ/U��ʌ���J�y�B.���S�����ic81�R9sǱ��m���"��㸹:��{{���y��S�u��)u�0|>����5����G�E=���;��<�k ��7K�������ZQyh:�n�}w�z�|i�ٱ�݌ף�궗�*ڣl.!����]��a���֋Ot��G6��N8��֜��ٓ�;Ie�w��au�=U�A�5u�oagF�Ltٷ<?QY�'�PԋΛQ�b9|	�$Ȑ�ҍ��ML
��&��
��6�5���� �H��dh��$�6s�F�7f��'I��Gt�t�^�O�m��3�<e���Q&�?�ǈqƾ���j6� ����~��I }/!�eED%��NM����~9ݎ�0�2��^a������@8�||0ϡ�~M�P �]
��G��џr�p�B]�o�C|ِdkP�3�����0	`���V�\@!R�6�1�B"��W��|Îk�x���ҠN�\��� �W)�S��JZ�\V�h�������Р���97���<�Պ��
��;c)��n��x��T�z-�;�ń�7�M%���qTtb:��R������n{�3�t5�q/����	*�g�<~>�%�P�(��9�s�n�`8�ek�J�U?�Q��2zcA�5����ZvV<Α��p >�t���⛆�4"�D0I�?�y3NAvT��z���k0�b��t�:i΅�1 	�kG���K���t�Hg�����:����NKؼx��h0�Z�!R�;WK;�)	�Vur$��d��
�~�m�|'�)G1�Q��p�Y�"��?�[O5���i·�u6��y0��˚�<Aڭ׻�炘[;%&��r��ڃ/irӰ_*�*b�+u�D*�AK�2Di��;�q�Q".=�d�a��� �/CDP>�B�9�}X�;2�1�����۪��o1{��DM�)()}%|b�%�8�$j<3���4:cc�߉Þ����ͦ-~�V4yk��Z��a����5��么.��/�C�7�a5g��!i��C�!R}2��'v�u3`�6���>��W�c�ҕ,+F��*�6Y�������]�g�z�KI����h���4�^3	�&��³�+-�;��)v�������s�@{f6HZ
Q���G���?'�kߩ\2�4�U  W��`�9Ap2�a%�^�TyZ�����B ��X1�[(����LM��s���co�04�|��T�ї�anT����]���s�YW:�J�e�M�zry�,��{�����3���n���܇c���L�����k_���f��`�^q@X���Q�
=��8Vs'ey~�y���S�� ]�mrc�eLnu*=��&���71#U-8>C�3ꝑt��?�s�R��ܿ�);���U��
V1y:ޮ��4pV����y��-FeǺ��"�K	3���03�Sh=Kū!hhu�?��7�z�A�?)�	b��JKy_D6�p77�QwV�������Ӵh2�E2&h�"K�P�q3_�2��;�GO�]�찺�P\Ʈ��4Tl��H`6��ŋ� !vE�f�ã7��2�W���G#Dp~��r2�O�2Yvk�R.J�$�Z�P?y�H�D�t���#�}�*\��Tcw���cgV	Y�
G�gp����p�1-�FUl�v�jֆ�H�\��� �x���8[��N�9O�Jr��@�3�3��!�n�"ۢr20-��Y�!|�Y�],�P'��H�'e���p��L�e��yYhO�
��ל�|@�& �G's`��f����Y���������L���Fe��E��N"���
kphсc�H ���ȧ�HT�E�61|H��㰠���Xp̠�c9}&��*E�����'�<��o=��ȥv������9m3ܒf�z�<]<\�9;�t�t�xF8� D�,X�i���!+��
�Mu�>�f6�L��Ŵ�4`�L�W�
���	0?PX'T�ի>�E�Z��&=k=�p���5uGb����+\�+4�e���1�������(z���f ��܈��>�ʴH-��KzvŻl/�B��oPo����GN��$�2��?�u�U8hxs�W��W˶�{���}R�C���H�`'_,QY
{�S�³]:x������`bN��'�,���Ҷ��������m'u�h�qq��j<�F��	h��H�s	"��la�-Ӧi� �w,ܒd���D�V7Ty��@�=�AM�ǹ��ČMz�����E�[����7���t��+�/xư�rĳ^����q�z[���6G�|���{٩5�ije��=�mA},�I}O8秒A<�ɞ�zM���o�rE)��Y�X+7�b�؛�ZLi��G�O5��7b��;E:���F"��*B��5y;N��VwLpJ�f�Z���~J3�wn�!$83�