��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E��`!��O���i�*wX��&��m2�)j>��X$�Fv�Mfca�e��q��1���:�vσ{��e�b�Μ��f(g^�}���S��x0l��wp��s4���圱�I�����@(rS�wm/�.
R�Q:2�3��>��7.�[e����r5�-�I��N��L!�V*�\�P/�t&���<�A:h��������gS�6Ǯ�w�\�8����}�� `eck6�Ǵ-/Y��-�N>5�^!�GǢJ��,��<;�uӠ�wA�+7i-��s�]�:��5�Qr9b����+6#.�
��̆�	j���R�#�>m7n��ݞ�O��#���+���6��Z$0[��0���*��(��&_μdܷ��<Wx7��?�U�XC���,�x��\H�5�&S�ϕ�4<�����Z����E��t�^=}1t
�� ���g��sx�W������>^�U&�j+a���=����0I���_�ϒ�*ֲ������@ @QGA��g��2��t�L��j�T��"��f�)&}\gf���h�T�,,�㲘N*��<���;�s�4w��D���Z�=�7r)�TS���f�j9���!ک�������$�m�{t�h"�!-�,f�ՋZ�[���D:�yH�\mSd3���|�V.'U2y�2#z�ڱ��O|Fc����T�%�J�_��4T�iI��V�;�d/5�i�=NkY���i�?�^��e��1��ګm����YB�9�1Ng���.�)����&u|s�.�0�ѐ��m(��k�-�tf�vs�0�W��{n��ʚ�yI�c��!1q�^ ������Lo�D���k+W��*�� ��o��E��������`���C$��Uy�'ϰ4�b��`���k�)Jf��� .�
`C�U?�N^��E+3�&F�Pf�QrW8��A�_��40�U�u�]�0Um�1ކ\�����z�|ZY@Z�D1�XGէ	ymrgU�E�$)��a��s0��i�6N-�,��S z��<�Fr�V������}��by��v��Ut��>�'�:����ݯ�El����}�O$~g������~�뫋�o7{��v����ed�WX(]C����4�E��]NAi�oM��d�3\'p4��0Y��\V{z�	;Ԕ�u�hWv�q�4���yB~jű�tFG����&E�}e[�ZO�~ ���3Ri*"7��5�t�8
\��8�rU:����{6��X�k��9��ٓ
��^����3��h���_3/i-ߖ�<��������S�W3t���Wk�U��
����ւh$G����e3G�&��	���e���E�/S\���@�U<�a��$m$K��ֲB���p�ʙ3��a'd�IF�N�S��f�FL3�5���R:�����tD��G
�Il洌+�QX5{q!Æ��z�9��aw����!|y�!
�/��J�M�7J܃gYѸ5��f�#��x�k�;�^v�4��C��U�,�2T@�#����5FV�����ϧt�5]�F7�N[�>��+>7�����kh�����$qR�AoeI���/(���uJ�`f��ָ߹�y��T|��M휔F�������,oĺ��Ͽ2T���������,+�b?A�Z#�W1�B^�4:���O��5I�zi�zxps�_��e�
��N���"�D�&'3��.�W��gY��;(aol$}k��R�-bC-Kښ�*h�Wv9��F��TE:�5�rc9宲�z�?��	��U�L�i=�M&���p
���*Q\+w�	����gM��!�&��, ��q��X8:��Y�m�S� G P�	3���6sÇqs ��l�X�l0�	�/��/J#޻+]Bx���n�?�<W��ф!u�&��DmD��,Ӑe��FI�P^���M���>ȣ���@���[���Q�x��nF�Ž�y��5Ȧ�s����@sg�WHm��j��	P��8\U*��!�q�<��`����/I��b<��$���G�+>:`_��CM��!���K�3�s�w��Mƹ/uM��3!{x�4���"76hv�(���	��F!��ዯ�Pk�qН�hf+�����T��P|_c�CqU��@�� ���sޞ��4Y\)�ƓF6���X�$�ܓ<� o��L(�.X���ϧJVCT�F��^8�p��-���	14�:Pb+�SKg�z.�ȼt%lĔ�Vw'F����K�φL���m7v�y'�[q��/2��i�hq�$=j�"��tʢ&|f���Z#Yp�k�aF�o�E�G#������'U9�8*�)�ې@�`�]'��?��j�p�;�9��`�Ch�;`˿Y�h�N�>�O��Ӌ�J����q�wphxB���&3
��||�:�>�P-���>,S�ii`ݝ2gHn���B�j,�p��p�[���h:a=h�+>K�Z����cs=觚- ��c\:ַTͷ��5U�ӟ]�)J�$<Լ/c�w�"�͍��ƍ�R���á.۪j������9�t���C�9�A�Ѓmj������!$��Q~��i׮�1,��V2?��s]wy��G���Q���z8���u�X_�}����N&�iU&��72�./��8�n.��.�F%�YSX�ޥc�v�`2�L;HQr�!e\�E;(��;��vO�����/dv	q����X�zn���XH�K2���95oY��S�ɇt/��ȣ�mx60ʛ�0�"P4���>]���`�1����[����^�>\yRu�͈��W+�FGU�Q(���W�:���[�`S@I� ��ԣu��P������p��%�ơUtʬ.Z R ��b�k���Hy):�|uAY��hOY8�5�y�����R�@��� ���_��MK�x ��5M�D����y�<�P*L��.O�[ܓ_���@g��&�8=���2�ܑj�_��E��G0CeX��l>J�b�M���x�Q����Z>���"� #�������{&�fl9B�9��d�[��yR���&{��K�G¶���!0��C����`�i
���K�uy�ȣ]����Byh��GH�|��Y<��4�ubg��z���P�����|U���qY'��_~#�����0�@�s�Q^��In�j�i0��	�/��!�M1g�j�E�̊�J�#V۱]�Ҵ�Y�Xy��RGߛ�� ��Ɩ��f�~�/W�ɍ�۩JCCW��;���w��N����kw'��,�ѕ1�>�eH�ݺ�q�g5n�\����AQ���UCTT��B��?`�i��?T�����	��<��ZJ�r��(iwa����e4��CJRz
\R=�z����C���𰟳}��'T��M��eI��Mu�����T~0��hR�p1�/t�X��uS-e7��.��Qmσm�0��=��+�(%��3�Yl�[��+��n���%/<J��Mr\Ua
��w�\<^�k��v
�gƭ��=G��gyzVpW�M���Ciݫ�qN	S�l{a����PZ@?�Z�D�{���eZ�f�G�`��>�0��H۪!�;�6	�4A��"�b�<����e�����9�)\p֊GΧo���	6����"���j���<���J+���ȷ�RV��S�'�R7�]3�5��+Ǿ�l��V�6J�O���Yc����p�&��IV���w�Y=v0?ec+(�i!O����1e�~ɧI�kVfh��������=�I?��d��^:j`�>�Z������8+�iA�(T(<m�X��Fpw��6�#�|h�Q\