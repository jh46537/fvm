��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
�u�,k���L��z.vJ~ 5&�a�+�%�����n��=c�DS��D�K�;��.��]�W)5��4jQ�l��u���ݕ)$���r<��p��f�0���G[�
�!������2�n�c��Bl#�L���(��T��
��$�˳2�������O�Q���$�j���5���4�\l`<$S%as��^��n��=�;4��M�w��	ٝ��İ��T8��y���,��k�ne}�)s4=��x4ő�t,�?�~51c5��`�2��hG���ߏ���0SVo��@�+Ht���g��xV�/�f�51��6��fk
������d͉7�q1&�|y��p�Kʟw]J���{��u�ȓ]O�=���\��!���;L�po5�G�4f(�|�	y
;�lQ�kU��3�3FmTo�pܪ6n��<݅��L���h�滊�3�F �?{��o���7��9�A��fr�_�h(�-h�إ�}Fj��K�)��P#@*LM�:�L'�u@4i�':�I�7,�{3�����\�JkX�5��#p�nvEz5�TD�
[~q�qZ/0	�b)�3��vV�s�`eȢ)��-A6EN���c�; ����/'d˳6��mŦ�K�A��Eʔ�=@�������G'�O��7�\����F\�V�Į��vX��3��[%����j�����x������{�y����P�F������`}�ݗeC����2��s�%b x��^��͔�2?5�C��I���dRtg�+`�?��,_�\6g�]SH�2�׭µ�����ߦ�ǵ�P��u��m�\�n��	�Ũ��}�1�ȗ��B���	GT������x=��
�̃e��N��;�G'�N66��<�&��z
�r�h0�}����_�<�t�}y�ƚ$ڸ�1�L����7W�Wg	���]�ȟ���p�ѽ����:XS-���e"tG�`�~��J��ł�e5Ձ	Z��e�l��@7ӏ9�wQ�� ������õC��A�4�_���U�%�I@/0�恢2#aS�+�[)��|���~$S���uJ_K|I3� ���x���]$���iO�y�9 u>K����]��U��9�p�qȌh]��<So^�Fe�?��`��SOHӲEK�t�6a��ƲJUj!�}MO�ۅ����n8{�{�����Ɯol�8"ټ8���h6�R�ظ�W�v>�vV5�!y��$�|ψ=͡���G�TL\�9�2:
;{eh�³�o��4����|��9#��/�cO������*y�H�@�!�It��ܘh[0�X}�x��k1�֘5��$}�F���嚲�E�3�u^_�
�[,���r ���z�|�J��j)�!X �Kfs�ފ��m=�����$�~G3}R�r�1ۆ�����V�FG��4/?L�y��K�b���F"7���V&�1�M�a�A��q��ÎO��U��ぽlt�$2OӉ����è���3L�y��No.R�p"�Ф�J���X��J��V�.��J��%�Sţ;S`�<9�{�!Bp|���1��XjN$_6�S�R�BN�O3�
X-�T�C4L�n����5�C���^����'b^�la[4��xUayx�_����0t�� g�tax�4�q�lg"�#H���2�dْ�Np(��O�aj�����݈���=�):��r�Vդ�b5�ce�D9�>�*��'�['c��#d�PgF��Xb8N;:t�?S���tg���k�F�T�j6�,���hT6ƫ�b&np|�-$���:)��xD�l6Bo ~�a�"��ݍ����vD��P�z�v�i���nY`(ot�W���-��z0�i3��I]��6YBJ���C��/�J���y�g����w{��ur�z, rE���T]� =�ڳ�&��u`M��L���َ��0>�/x��3t}���Ǌ:5�&Ҁ������%T.�練�5�Ҭ�;u0Np�E�+v�g���|u�]���Qm�����Ă�����PT	��յ8+`a5�c�\7���"�J�*��ց;�S؀����1	u�;�B=a�ܓ�9�I�Iq�ZW#3@dDoM�X`u�M_���ܓK^^w�������ϿS0�Y@vr.3���a5��:#�cb���K�ܻ��Ҁ��@��W�!�*3z��6vn	��*���.��J8an�#�3Td/a�N+�,�r�=̀$�=`k-��� J9Y%]Wa1	�eE3���d�V�-x��_��[
V
Z�E�"���*|69�t˂:�6b=dc3 �qꎕv�bf0b9��w�@�%U`���ERXJ+���	�J�CO��%���a�$���$<��h�s6k%ba#kVG�\	�"��E_�K���ĸ��r���c�V� f�O2`Ṝ�x�t|8��l s�)�'�1�̵%e䧠9;� )%H�oľ9_��)�L_��Z��/t"@�Y�� �Q���}k��Beg��̡՞Qo
������Zy8�,�,h6�|8�B�Ƿr�
82a��j�zG�e���-�󀵱ɛa��e�Z�j�)�i���==xhta󶥃����m���}1��tZn�/7u�,)�Ĕ������}�������݃��p�!�8�Q��xl���d�3F#ZX�occ����h�U(����u�K��^�H#� ��*�<��{�eSa����l1�2��:�jE,-D�M%�))#&mYJ�p�#J��Q� c 4w�$�ƺ49����!ɡ5y�*yW���)U#�	^�-�0�*ELxQ��O.@6�?
l	l���%�Z�M�\W��� �!2���$C�~}�ꢜp����Cy�l�������[�*�tD�0�q�+�ZBQ%Ϝ��`X�q�}P�;R�!I׹0x�yM[�����ޟ���S�ne���v.��j@e�h�b�2Л6� iӕ7BD�z���c#xv�E�Bxs�!�*�H��p�������Gq7	��5"�W�qV�>�c��Á݆Z<�<�֐��ȨL<��6�Url\�dhB�(�|�Q��O0f�`�'Dt33�t�'��R|��㚚��1v<G�K�\/;��ӓe��W.����I)p�^��6�58���e?z1ع1f)�·����9�`Y9m(���ї;)XM{��� :1���i�`�jR�2)�6y��d�@�$A3�%�vun���N��z:�c��v(I7J7��&�vd6����;�!�}��F���q�	�|/a��Ap,ع)1���!M}aw��cu��g�-��ڦMl긵��ؤ1<�uym��j�[$����1ugP� /HB��
��V�&q��t8gX�_�.�Ů/���A�$�nk�<�(h�4� Ւ.��ES��(+����$pJȍ=�~�>�}�4HOW$��%��hy�W��I��mqL��Ʋ(�[q o���DB����s�k��H%����"c��"ӅK9;m��uB$�B ��R%����,`|)ip�~S����{ċ�Y����j��pE��eK�$��0V�:���m�o�����'?�|A���������d�XD/��=����s	@���f!����5 _�G�SS�kBFʁ��N�+�*��4]M�ncӣ<�9�l~�z�{��P���SlP\SOZÍ�)�&16�{���a�([�6)ɝsK����Ь�\�\R���Ϭ@m�Q�W�g�'5F�s�i��8Hq��Im���)�kc}v��$���HI���ߌ����}!�8,���bU4�����Ϭf<��IN"�..��
.�����"���\����"`��Ŀ�  �h�_y��}�$�5T:��n�T?%EL����`��B��\��pr�V䇔�~P��D���Z'[Q��P����[h�%1�W3��<K��U���P����?��%�xLDk�@|',�qbhO������|��%=����Ea���;�!�������&p�tjɒH�F^��D��D�b,u)��Щ��0���3a�.feZ`��y��6�u@������<�/�s�Ϭ�v(����ld�m�^�~ ��(렁cŔk�7��Yp��H�piƫ��� �Ke�
Xm�Q��a�3���P��4"��'�h��A�f��	�T8p�*���?o�ڭ-����8z�ł`��,������@Z�)&`�pE�t䩧�p��&,RUS��8�R�̆3ښ�z�bk��3e��w�)���U�a�ӈ�x�
@T���3N\Mg]8�=���	��s�r�ϕ���,`*��.�V��4gW�nO~�px5�ʪ1�Ǚ3���C�p=g\`�#J�=�g��y3���7�4���;�5����p�]_A�]��C[jm���!<� �*�l-%e�|�L�7�Xo�ͻ�49]~��!�s»8,�
#]��W���NI�u��1"�U�๘��'�ި��8���;�̂�a��&�� ���9�6q�0=[w�R
�I�DkG�)���7���u�};���X�A�x7�Z�2�8�Q�7�e�Q/-h4wK#1�p�)�����Y�=�nm�"������EaBD_{�x�G�=�./���vb���h_!H�v+��'A� �tҁ�v�w_>~ׂ#�kY	]ʔ@5��n�e�#�ڃ(+�]�a:��ï�ru�4[{���n�-'��:�ݲr��ᶍ�-���T8q.QQ���U~�U*3"޾%�'1z!��Jk�K䒖�\�m[��\���C��������aH@��L�{jƧUuhS�>X�̆��҃|8����Me�Hd�珴kȵ�s�0�>e�����}��EnB ����2j���R�!��d�t���*��y
�ɸ��Pk'֪Z��>��������������c��^J.~,�OA�Yn|r4H�q����W�i]#|�X���Qۨ3���-2���	dĮ����8�G%F^[�8UQ�޵E�.}�,9B���y��ت��}L�g�U�'O��|m�4�8f*$���3ˤ�'D<ۤ�['�@H��I�M�rNY�C��U�L~�(��m�Z�%� 5���_<U��aw��tu�;e��Ö]�sa6�<�%U����;�<,s��y��9���~�Spl��h<�|7y0���s2���r�`eo֍ƌpmw[�����N�+a�i݊>�?��&^\>w�9�0����Eb1��$�x$8�Qa�[�2����D҂��E�,ѿ�5����q^��2�v��A���eap��Z��몑�����oe3�_���zq��dwm����I�UG�bCG>n`��CA����=�,!�q��J��V>R�k~�����}������u�j�/k3�r�〝�Tw��p+c���36�7��Э��W A�_0��������zO��SHcf�p#�X�W����η�ЈF))})h=ƭ�x�y�n�7/��+��	B�)�M0�?�t �����]Eh��o���<�ˬ��vXA����R��4J��+�"A"�M]a/ �y�5���^��9��8~ �W� !�z�:�I�F#���x��^��+����'d�_�6Ϟ�����NH����iEY3�J����_����]!��A/CT��s��rO�tH�k�,v�ph�s�=8����G^�g�SG�5����K欰=y50�\�>���������H���7�7_�������e��Jر+�nE^3����{w)�4���G�U�l.����QD�TÆR㓕2���v�9�#\�(�J�v�+P�V�؟�K�����ⓛ�!�C���J�K�c�צ�%�}eCoIDd�%�m�F�R.%�!=�f�,�b�k����T��	���}@`;
9<<� �JA��D���k�hָ��m�4�����i@�x@G���j�#�c�\�t�E@��� ���b�p�7���B'��'�����j�2�� ;̈́�r]�- ��容 ��7�w��w� �,�_�A���J�:VB ����bIYBiX��ivζ*��a9i���&����?�j"��$��I &V���$]�ҟ/���{J�ėkH1�͂�� �Sn2��YM�r&-#��Nr�Õ���B0,g�7`Ru�}�cO]�y���ʧ�⧕��t��ڍ����Q�`�~ը�~G��aɻ`���0��L=��,�Ld|%�_��S:���&��y0}1�#��1TRDu^e6���h���-���b���X
k��ς�|���n&2�N-�C��I��<Hr14�sL3H?Q{vdp���ʣ0�[��#�L%3,4�Xm��aJ��Խ0h�]o	֒]�e?��!jU��=X?�z�/�&�W��e"�;�-b�5�(�N��c�A����̏�	>B�X|�������W%9�g�R�«��q�ޝ0C�Fbr[,D[�@�E�\NS�w�� N�|�K��G@{DIWFW�u�c��F��3��B=�hS+��1[I�#�g�B��d�:��O��YF��F���X�~�4t�>d�@:�����	`%�����\�|0�*d��!r���lS=������c.�,�{�:aS�D;�c���l�>����qV�4��oVcJ��կ�-������y��y������u#���I��>
��au���7��)A�� ��>���}�f�	��{O�}I�	��Cs�G�;{<ń`nq�V��O�"��E��x��	A�o��-������.�I�MBI#5�7��K�^�ўo�l��
�=	�:G�쐡Ty�.�gڑ#�1�{�6Q�&ǫ��)��#lG�����n�p��WP�5H&�	���I���y␫�>��*�F���67���7�����`o?{������0����2(��6�^���#�#�+�;��g���C���I_�)/��ըΟ��{7N�Eó�=�Ս�2�/�+;xy��|���ܥ�����~欻N�p[D^y�]����?��������]�����Y��U0�S�Шp��T+�։�
i�J��i��xz���h��9(5��f��3fE�He�z����+,��җ���Qtr��x�gO/��e,A�v\�x���F�p�ݞ�������Ź.����<�\����6'�sa��yܺaO�H��,�-?��Tc4�@ �p���7p����#I���3�X��3�>Q��UҀ�5BbŹq�sV'�k0�	uy�>�sk;d�F�)���v�\�����u�Q�a�w}�"ԛ�¿%�B7`���З�d9v�L���	�Ř:3����k�9��*B�x�'M�P$|*-)����bO��p*�B:��h��g���X��Β݂�1FULN.��x����Ż�̧��34}E�h;����� O�9�
�0��Rrp��a�D�od�̧����%^�����j��U>���F��Rn�C����9�)��_}��'k!~	2^�.rʼ��׀�BPW#�j*_h�3w
��	8�f@��]/A��������5j�tb�����MuiN4����i�k�
�m4/���qP5�^��̻��I�/U���g���e�o�aH�g�������bK�ke�2���f4�y�;D�B��*�{���2F��LQ���a��	k����p�'���vt�8"���̶��FO!GQ�!7�;W�@��rE�bh#Y�;Z5p�6�0�}9H.�� R�VEx�"�x!Nw�b��t�R��b7[����.=k�C��kc�[���a~��j1�7��ܛ��{_b:����̉|�(�� ~vo���A@-�Qp��B����^9�粺�n�ē�|�F�B)����zQNӆj�C�&��AF���?�n�/VY�Ru׋�6~�Q�17h� 
]�eû]�%��m��1� i���5�o[j���f�ţ��ٴ˱~��X^��f/��$~W�*'��ןBY��IP�qt��ID��%L�.��	�0ۉo���e	]w�������^�z,�O�`�_�J��4��5D7��ܦ�T�9�
��;�<u��#n���k��#�4]+;�Q+h�7�ŋD�4���՜�r�'�w�	笞=�O�3�l��{(v������y��F~
`2�d
���"nS�d h����]r�����~Ĵ��F�t�8�O�����r�4�8��s�b�u�|$���ϕ��$Vt<L�����A����8pf�J��ܸ�P�M1�6�Et�Y^u���>�"��x�e!�b��X��.=�]=~Z�&����'���
�0����I y^�o��B3��9·Y�l>Ec�<y������=u�5f5�kpE��)6�p�z�H/�Uz�"��A��q���"J{|O��j���;z���Q:m].�1���T������@}*cـ���_^%|�d�t.�ZG��ڳJjl����v�^z@��^��,�;���2ݒ[�Vk/gp^���H_E!�{���q�5%=Xa����d �U�\�	
�&E��C�\i/>�ma^I*}���ٮ]��c��6;�c,?����ɍF�6��'�Ґ G�l�2�Vr0F`�p�t5�?̊�Ģlr�kW["�����F��3"�.j�TA����q;R(�
R�[$������a�kK�R��O�o�ɮ�y͇��#gvS^�ux��+��0{$2�M��O&a�.Q"����t*a|ˏ��b����%�dE�{�5�$D5�A��˔��#)�Pp�}��}�Y�M��s�|7L��~y��+U��/��_Y��3{x���/e��ZwOP������qvJ�Y���o��8yhu!)�D���ԅ1���.�I*Ԩzt$K��J��Kt_�Ud��6�ȶ9co��vk��G��RoO�}�:wNHP�B��^df�]�I?�����FG�t��ߢʧxm!���Z�ғ�٥�`��.�U�*��@�Ary�+� ���/��F��;x�ڹ�H(h~���SE�c��ӿ͆^���>Wp���H�է~�n5��njQ!^'��c|���"b��<����	V�&�f�bh�|����u�9�kJ4�ob䒅������!^���� �uf0�'�2A4���_���~̌n��JQ�0������..a���JKn3W|�#0cw���&k��5�*TlB���������O\T�k4����ZY�	}�z>R�y:�]և5)�"��ׄ�y�	ϟE��Y�J��(����|XK�������Fe�u�&H��/�~�m��;��eN:"o:�Ӕ$B�=�S�l(/�,}L�`����� ��
�3�~��(s��k�ʵP<��r�A}2
bHa�v٧�;K-[1F�`ݼ���>�*_F�e�)'�3K�f�'�9� 0y���H��������h��~���!U���ț�

>p��������-�p�]Ⱦ/|Ƨ�����2J�^y������.cuWI���!���^�T�]j��bʂ'\�O�)6��J��R�����F�O5��7�[��n]((��y��db�/���qvV���2Gw�i�����ˣ�j�1�X(0W���8VP93�Š	m�>a]׍!�u=/��9r�K_,����SF��G�Y����d��y��S���-=f��@bH|�f;ޙ�l��C�V}s�<�
���Y��$JO���͇�3.��`0�b��n�i���}�P���sxH�#y��&�T*6���f�F0#V��)Ո�����gfp����}ɲ��C�i�e��ױ�z6�)��$���&��U�*n̚��׆�Hg"�&���=[��	�d��ܾ���bi]�v	i�"K�d����#4���hĽ�/�:�9�����-�r��3�p��
zk���Q�-���M�8#A|'�=`��<*._��!��b��B�H�x7���B(N�1�.t��mQ�29L�1�W.��ض��m�N::+\���sO2�3��9ۨS�4V��S�5΄V���|�������K(���y��d�B���rUm�-D���u�x��G��_�Y�d�{�`!h�ٳ��V��t�dx�E��g��='�W�ٙz��7�4�r3s��>��r��	��%�qC��:f���zfS��� I����p�=��Q�^vʉ��Fx뢸�k�ڍ�V7��Ov݌"ܺG�4r�����1�sY��4��}<�8���m q�c��D9��R�Y������n�-c�L��z���
�o�Prk��
J�-m]d)2Ǝ���ݾ?��i$��6/��l{��~�wj>�����ҼпY&rX�g�ve����]�r��x���V�nVȝ��Z91T�kp��6׭��o|Y+ q�N%ɟˎ��m�l$�Hh6��h�T�zW;���Eʙc:ԬX�"p���X��?�*��<0��>9�5�I�Ts�_[?ƝH�I��z2,����3=�I�<�z�c������
�Cf<�b����5ǫf�+��V�j�07�҉
�%��.��� S�b��~���ܷ��2��3�7�6^Tru���N��/-�#����j� �����Ջ1%A6̔,��9����&�r�U=�/���P>v�VI*u�����y��^k�`v��{��
Y��P4���(�(��#���?��u��Ә�����iӱF�'3X�,avzm�h��۹�~#����*ό���(� o�/3]�[QQ@"��<�w<���'�����G;e�8��vs��dFi@�����������Z-�M�R��+zǩ6����EY��=؀��{����W��`�nLX�w 2������T��rW6`~�@ǧ�ر�i,ή��)3e�('��
�Iy��\�����@%p��'�
t��	�t�ܚ����s4�� ����)��O��r��}	,]lD�Z�cq���}Ģ��8X1+V��1�f�����}��u ��w��]��p��c�+���z���#*�}�v���kE^i�LbH�ߧ1�������������\4�� �o,��wz7&�Vϕ}��*٘�?!
m�M� �ې�|=J9��S߻���cn�a�S�؜'t�Mt�4a��OUDS��Z�$��mY���i��4���y?#��?�u��Z�%sV�Tv�JK��ҕ�R���ظ��٫����eS���-��%�/*�P�F�ְ���1�P�C�~�z`ķ*��6y���Ӷ�������ԯy����ǴD�6R����sV8u0���V6�x�6�_���Ǎ�j��LX���=}�?�3�7�7�-���mb���hQ؝�+���{�Y��[{��L��O���GF^[� )���꩏�B��G���L��qL��W.�:Y?��t�yp�����\�� �[�q�Hd�Ӕ��B���6�~�f��ր4l`�c����@9�j�H*�#�藺]8�}��7��ë��^[���������� ��Pw�f��-Q���І�m�n罚y�"�C���T}E���i��*n��īn�.�o��V�<?��[��#���q�m#��H<QGWQ}�+��M�)%$Z��,ԥG�"��`�ZT�K��ÅA�Hp��.zӕs3T�.P5���/��_5�br���iLJ�Cˮ�G;%�_��E2� �׋��9��^�Ҋvz(i�Z��-�D�El���|?z�ML��_�&T��G��-S�?�-E�tC� (M`��?�?���R���|dvƐ�e�M�]l �K��~l�#.z]�P�!�Nu����2i&J
2FX��.����&GƤ��NJV�����-���viMEXCڱY
��83t3�ԚլQ�X�����<YĀKı�GlϦM���\nn�G&_lQ�݅T;F��/�~�ˋڬ�x��x�ޑ�_�,`���%9�1��� �̀F|�V��O�`����������XKb�����)��Z���@=�1`r�֎�㺄L
�ʈa\�(.<��N�;�[�h�_ՙ�J���Gd �e�b�ԝE$u0n��L�#_�����j�æ4(���-��|X���V.宮���P{�;ܖ�*$�M���Ü2�'A�S��-�v�R��p6��*�;.w�ر�C_	����,���>����ӠC,��>�xT�GX�e�ӭ���yQ>��w�ʉ랄j�;ѵr�x����9������u�I[�o�c,	i�+LϸLRҾ���XZ�@��Fs��I�}F���b��2<���渘��m��CJ�:0	�0GѬB�6%���'Lۀ�!�p[j
<KgE��U�����I4��2x�
DɁ�x������*��%F�Ϻkʜ��W��]6 ���߽�-� *����=Ho� S�b<2^�[lH��#=�hE������fw�k_=�@$YB�g��] q�i���_�fe��899Y�e>��l��Lm��o���fA6A��:���3��*�ZL���~�3�|�3/X�	�بh����3^9��,������0���w�i�xOs�w���?%���YDz�e�,L{^g(kԛs��%��~K��xy��S�+�CEnf�J�n t؅~�*@�;AY�$���[�M���$o2�t�fT ��=$���c�o\��'�*`�DI���Y	�k���{|7Ux�k�P6!��@p��g|G�_ƥ|g���-��*Dƫ����4P�Xr������d�7�b�������nUY&&#�n%�j
��|O*��Ϸ��[_�M�n20d�)|������(�K#p^rtY�8��`��I�����4�
ERCS� /,�h;zc/
�
G���j)%Q�f;tW�c�ߪѭ��vU%��H�U�:�lNv�Pugr9f�(��DK��z靨u$�#~g�����;O?�~]�0��� ����P(4'm �9�zt*��>���iM:��36�r��B�Bԅ��Uͷ���]*�/�-FMm3l(����Ec�q�9�>t��̒7f�@���ߜC�w���R%/�*����Z�U@��@LU�r�b1Q�<��偈ť��E?�K�߅	a	[Q�8��*0�3�����N"k�j]�����T0'ѱx).��?��yl�
�o�ruQ;�%�{�B+�b��eB�T^��|x��e�G��C���뇂����L��n��)~uK��т��`��R�C�F�����=�X�$��Qu��±�7��x�����?�%�%������6��/1��V�W�
�U ʧq8���x�Nd@��f_Q�K�h{�+�:Sa9��/ʣ���M�'%['��O�1���(�?ޑ9t.�n+p{NV�1[ie]�a��(�R��9�ؖ�j�M����Ϲ��WfYd[��>�-گ�S��8ꁆAR>Y/��|����?�-dD/�\����s�*X_E�g��]��n�����,E#4�sY@�oW�}�C7��j��P�Σ�+���E��x���yx�P�TGp��^Lx4O�h��J|�ާ�B�uo�|�sG1z�;8�й?ZD��Ȃ1]A���)��C/,�9\����W�~��x����V{���3A�Կ�@bD��g(3��[��B�<%b��I��,��ѕ� +����Qy��!:Q0�����f�Zlט�"�hKp���������O����p�P������]]t?Ҥ{��">�yo>N�4	5�"�c���E:T��ڒ_��L"�*�-�>�Ι��sߡ��F0]��6����[�Α�.�(�v2����7.���ߡ���$��H���]R��ig�,��aBU�]��83W�T��)�������Y#TS�Mu���ň�2�1�b�C�V��WM6'�r]EJ%g6�ш�0b^�fi�N��'�����1zl�N�Q�ˇk;�.�XZ�.?�4n�p�M�?�FR���q 6�Yn�n2���~�]��[���J���m֛|�u�!i�%7-�n���<�5��nm�4��nn�a*��#~@/�艓�Q��
��A�g��ZN��J-�Y|��#�)�x)lI猯�`�,�E{�)�P\˄RW�P�tI�8���TL���{⢆kFzq��q��.4s{(��Fo����y�xy7��MN�7fbU|�d'����i84�-�L>�������O� � �_��'��;�O+A�б��X��0��r�Q��(͗��L�$sY&%���)�>�����w��ym	�3���f�g�"��aP�,"?���W��֔�[T��7��e�����C004�w�Q��#�����ێ����
	Ii�pޖ,?j���[�p�v��f� ��FD���I֜8
�ũ�kj�3����\���w�x�hpY���̳*���]�P�W����(��_�x��;j����u�>(�S?߽W[�D���� �ǫ��r�rK��c���g.�A��������^����Z�/f
�)7��6����iā�.#t��aքC`� }d"���j�{�����é�^��&׏T1t��C��n�J���&E����?�{C��^�]�<�I-�o�����z����%�,
�9H�D�赪��p�v�-m���0V3t�:{kU�O��	��ي��X�lU��=l����#�gR�-L�	[|�*m`��!�K��9� �T|o�<g*�IԤՊ[g60��� ��=&hN���&�����o�}����%�9.է��	!0/\<��8����]!#8�)����{P8���|�W��hr
���vF�������I���_-3�osڷ2�

G��J�|�
5+c❁��c7����s��P6���\��������@d�RH�?��X�%�|(��Ѕ�B�|!y�p�d7�iD�
u����N7��fx�a�f<#�rSDnүӗ�%㊦(�'�[��X��=h%�BDb�k=����)[�	��A��)��L��oYC�m��dl?��C�Eg���`-�9	_:��V��9^��h�ŏ��y����h���A�I}`$*�0���c�1_����!d���!�l�*`r�O�W�"`���vo��.�	K	Q��㡎��E0~,�����(˻z��@�$4WL}�Vm��d}ay�W89��M�u���;�I[���02��\���ͧ���~E3�v(�3w[Ԍ\��H�)���c|(O*��*�[�͠���N����b] r�K����%i얷$'[���t��)�II[:�"�Gor�_y{*[ ʜp��ylQ�!K��۩�|��Г!\u��LZr��Y�k�"�uII'_�v�"/]-�`�:��=��<,M�F�X�`��]�J�e7�1�\9��������!W����{0��4�ߩj��_�F�rXa�9�?���B����� /?g�x/vد2L��o61�p��c�l�B�v�x�xr���텘�-�T`y,0��L������dW��*ûQ�[,,�u��$����'K8hdMu��>o�C1��j�'
�w��c�>�G��r1����L�"����~#7��&�� ۧd�7���Q���V��.��W����6�q�G��7+��^�'�hT?�h�'t�Q����լR�m���$U�P�9��m�m���h�6d�Y�րzR�|�'��HHm��$��k2G��R�ɷZ�G,�%�HI������������C0�0��!�F�is���)�������h����|�pC�7>�Jl�h�*��A��3���aS<(�Ƣgn��<{�5" "�%��?~�d�f����55-����ӟa�7#O�嘌��C�+f0>çX`K���Ӡ��{�}�ST��cN�S�VaK�^kV�О���{|J�n��{�ґ1�9�U�zKv	��5�i����Y>�C7|f,_����	����.{��)��=uw使]a(��nL�E�"�����u�JU���$qh%�ϕ*����N,�����V*~q��s��twa��b2�� ��f�r..Q�� �7���2t����34�̣]פ�ЪQ�{��}@Br�s	���ܖ%�W^�&��B�Kkl��^M�m�{ܹXJ���ރ�2ȀVS̀��A�n�3	����Q�;��0ݪޯ6U�p�*�@Th|?�����%�k@�)����<p@Ҩ�#��r[�.2-�VP�2�͔}��iA�1�[��b	ƫ���.3����Q����v@�����Р�Ժ~���ή�n���ۡ�m۟�E��է��K4��;?�ᄶ $�g�[~m�>�!�h��^�P����u���Z\�^�`����nxC�ׁۑR�;�^&��tj=k���������J��&RH�D����"�EV�4mQ�K����"�ɥG��.��(W��둪�B �O���~�,׀�d��ﴠ8N񘌉�/ܳ\',_��<�@��~[�?�/jԶbA\:>�F�b�����A+|���7�+� ���c>jPJ�:�|�M���iQh�q�e�h ,]�?8M�Q�d��u�1PO�r���6ņ�|)�ջ��Y~,e�g�U!}�*e��L���`�C�N���˺!�0C��t\9`�ͻ�ʳ��+�w���.�&T���8��1E���^����۩�g�{��b�ΐ��lz�+���ʌ�����l�@)3kF��[�[��e�9��z�H�N�t�ro�\3�0f�7J�p�3�XCg`���������:e�$�h.N���e��͜���w�,����R!�52Q��&x�v;���t#��o�
"��j>�sr�/>��Q}WswlO3���Fg��j���&7&G|��ʪ1>��;����"�
j�C!�EҼ��ˋ����Nز����f�?�ӏ̣�Pfe<�f��-�>�=��V;��]!�;���M�g4� O��+��L:��F���v�M�x�$~�����c\S���uf�ܐ��u`=�.!���DP5���YD	M�蒲Fy78�ױ��L�B�`5�1�&���T?��7P�"����qRحǘ祉���T�yd��q�-⏨���_eu?��}����ߪ�|<���f�����lbkYo�w�Ӑ��CET�8�f �{F<n}��rx-���&����X�1��8��# ��G0k�n�ZY ��;���1,}!	���wfg*�n�xf-Pt�\�k���^�KQ���������߂Ѐ��Й�#"�˞����1��^�π�Jw�'8J%Q����g(Aԗz��^�E�� "ؠ��=�z�)�>h⦙&�{�^����C>/	�|J�ރ�8�B�/�Y[�"
� �Q���m(:{#�|�Ȉy�~ae
�b0P;�hghA\��m��S����t�_&����"*aȧJ��Q�.�0�1Lk
���#KH|���-$�P��ゎ.i�s��k���!�/�{ݜ!ed9gs�9��(�s��k6�f���p���m��By÷�‧��|o����߃��w��\�p��Ʋ�JQ���H�ZLx9n��LH�ݹq�f�x7:?��T� h�Ӹ�8p{!/?�̋8�����A���X���u&�^i3���[u���.�)�R��A0G�y^�4���3����x�69#V��m�g$f�4�!�6��Ν瑿�v��IkWuQA	D~Vq�_�EW�|�RS��7{�ڈ�Y������U��|C�\W�}�A�^8�A7��v"�uBb�"Yd�6���g�D7sϏ�n����@����@�x, ���t��(N�	�Y���y�$(�mV�4�j/[�����S�L�S�$��c45>;�0�(�U��x�3:��Cڸ�_�dQv�|�����9�-\�L������!���Awx�e�	%��� ���u�~�ςz��!~M���0B�h`����QC#F���Տ�a5�������!w�\McQP��^!����!�T���և<�f��xA��42�� ��fG����þ�O�
翜���c��bN=�v��߸XBy�>n5ڒ�E�����=DN�gs��r�Q-<u�ؼ�޼�[3'�D�I�u_����?4�.���~{� ���
��֕u�����zzuypd��A�����8R�(n����7��O�*
&���x.���ٖ"OH��f�?����!|p
��2"Z?J��:�{rѵEI��Q.����kY�Z�)�8�#ofn�h�%d�b��L&�s޿	ٍ�"8k[�~��$�|cl; :ԣc��"N���e���5jJ���Y	�ލo��:o���ӔU���s]��tȗ����at����3(F� ����`��eh�ξ�y��6B���ra� ��EI�v$���e�&���͵�A2��M���?�<%�Ź��Z3m�HM�i8�2�*�
�<�O��vbJ���+�Yd~��������A�r�m,1�����V�x���i�C+��ELx/��{�@]�JvN�
�h*��JU�A�?Kש�V��s'����%ܟ��c��'�X�o��&�'B�`{YU`A�oVs-R�D�a�(c�;Z�[�Bs�� �� ����*E@9��r&�,g��\A���ZIC�e�����>Ǌ�Þb��\zؿOry��(ԇ���qnc�e��5��ե�g=m��i/��i�(��_��-�Cw�G����