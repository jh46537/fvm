��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���ymc����#��בsb]b�i��g5~.�wJ8���A������Z���4}}��gP�v��t� �$>����6��:�D�ʸIG�ڏ��ӗu�\X���l��F����Q�sm��r�����)����&NsGɚ94�	�c��V� TS39���wĸo�W��'�FK���v���T�Ö������|���wE�+ ��Q�_4�[`��ވ�v�t?\���Y��A�Bڋ�L*��a�O�_�#Iޕk��.0{�Κ`�z��W��+D���ծ���!�j	� &�P�IE����h���2�)��\*��Գ�_���)�$K����4��'��:��~���*����w���((�-���^|hʫ�nʒن�y�
��AL�ag�b�b�{��@�XOa?/�n�������UV�}V,��E�.�seo{�H������XjË^�P��V'`�ս�Q|F�0��m����&�94q��%� �&����/3Eq���=�&H�6
�wNc?hR���{�dn
���R$�m�yh��	�ػ����a@Z�<ҠJ{U"8���i������`�L�eu[��Q Kj�7�_�J�g߆�I��W��ghy[�35�P;?�����o��NH���_����i�jө9
^d��-������ګ�2���}�5������XS�O�����ljD/��2�E�� ��Kl=�Q�ӖL����;O�ڀr��)�p;���!\�����B�1�w�F�����舲�fJ�|:e�uѡ �.��_�e-�:�z�x*�	;�����'���@)1���wʫ��%T���Ù@-�j��j�?1]�cʐO��~�����+���ʄ�&n�X�("����5s�m;�$B��<�p(uB��ћ�uh�DZ�T�jݣ�ѻᐉ�u��k����A�d�#2���t��6@�UM&B9z�j��]{�2��f����Uڂ�3K�������ƴ{��1��W�Jd��W%���Ym�DNaR0�G��t�ڇ��ܚ��^��nma���*_M�15%� ��ȔlO��a�	N"`Q�� ;�L�ܛ�"؝�)FI��읁���[����Ξ\��kJ�	pO6�� p|>�pU�s��9e��o���s?��ފV���<Ky1�3PXw�������d	P�U�Ǿp�"t�����hx+6��u���5�� U^�~J��9�"�O2�W�.��i �(f{e6Ǟ�j丒~�*�9�r�q����*�TkZ�'6��28F�t�zM5L��-��n��h��O��415f̸k�-u72ƻcW�0�U��������?��]3'#��1,�%!�&�rz�j��KmDe��XO�~�u��,��G���)yOzұ�~хf�����/��n��
l��.��Y��l�AG����v���_�W�37���=�� O�ߠ�GJ�Vթ!��͋u|E�%J�������	���E�oh�/�i���r�.��l�U<#��i�k�ѐ�v�|y=�y��=�����̙@���<��*�~�t����Zh�@�k���8�%�W�)��;�,�k!��m���L9k�(>W�ߜi�C̕��%IT����!f���oҰ���[Щ:&��?C��v�SA�#���sJ���=��
��6�_a��J�[k�����]�#H�,)���6SFi�/�N�JF��*�	���`�Q�������U��e	({4��u��;���Z4��A�Xf�.��ȁ4aS�_G�^�)7>����I1���W�6}����ZA$��!�P�!�G�^%�#
 Z��̩��0�N���ur?&(���ӟ��j��ӽ�4�4N�X��j5��p�G��PN����ȭ3.q���	iE�YȬ�Zh�U�u�.�|@ϻB��}`<��s?'�>RJ��>\�%\���Q�$���x�z�Xě���;_h6�eb��ͅ�=#��z0��!<{Q���Y�
 rq"�4�bF<��/�E�OչS�wWC1֋RU�g�XĽ]�)39dI��, NĒC<�*��[9+��*c{d���|Ϲ�����&b-�e8�i�T� ��;�����S�9�;~~�M�Yj�~�w� �^������x!�6ڤ�G����6�_h��R��3Rc�Vn}���#&~ ,k�P3P� ��$wp�Q����s|x�L��r�҈U4���эƏG�W}V_� G+��-V��( ubf�X6_g�`@c_�N^�����:)6�5��L���]->Y���?0#��A3��O*�M�r�u��m�O�A{dİ�ũ.	(u�ǐV���d�^�`=��5!x��4�
juɡ�j�!
i���g}���Xu�������3)տm 
Pk��"��Gpk-�s�9��[g�;J"$Ok(Fg�������O������t�*y�\���D�_�<�4�@ ��H�d��]�[���">��Vj�/�����PW�Fr��%�~F��n�eԇ�L���м5Y��Ɣ-�BAˠ���(�|˯�������=@��p:A~n�����~��������o��.��E���)�?�S��4Wj-�,����_���_�a:�^�,�1��l��c�#W����k`S7]yPʙu�0�1ϙYB�gg��M�m�Qn��j�Ρ�O�`N+��S?f�xթR�r��g�Z!�"�;��X�9X�󵦋|�G#�x�&�.�dҫ�`�*�6���M����l��ԯ ��`�=�I�Ip��E��J�68��\녮�Sp��E�b��"U���a�<2�2.i��|���/?�B�k���s���_���i��4m����Q3��нDF�w�3s�3�y�i�\�	P ��O��aež\���^څ��Ye�g8.v ���z�4�*��Ƕs\ou#)���IR�D��I0���O��Z�o\m�V5����R+WI;�a|�G�}����'�֩��LY �o�>��R��"}rn��N�M���)�)�.�O�Ij$	Q�pF����;
{'%�^\?������ ���PɗxD�U"��0� �#�������
LL'I¹k�B��b#n'n:SW�o�Tqk�����eQ�@Mu�Yj�~�6l2���"��d�G��/�BJ�������o�uv��P{	q<���Q5���~���oi"|:{���M�~W�6}�d��<��.{+&�P �P�,��� ^��a%P��2�^tl��%v����B��u8�/�j�V�,��0�xY�!�%H�(�p�0��2(�0?�YX�e��%���_���ho��`��ȳ��R�U,�L���|)�o2z���cM?c�H^�OӢ�$��;���ڤ�����B���?�yj���nM.�& 9�H[��Ki&�E>����Ϗ:z��7�#־QH���q�j���i7�3���Ҕ��+��3<:�F����x��n#�����,T�඲<�KE2Q־\�X��\����rM�!(����D���ѡz�	�}͆��`(�Ne����#��?2�S�^hP�q"�����蒎'>e֔g3Tn��Qv],�d���"\��4@nV�P�&�!�QkC@N���;�� ��#����%��[}u�r��m�n��
P-/���K�L��3�_���@D��X���#ӣ���v&q��t�?V���R�fIJ�{�E&��E�[:1�b�4�p>�f�v�S�'�?$RU
��O�`z�DZ��	�p}������V}�J�e��M7�l[^�[������ 8� %
d>�fK��M�/ҭr8��t���~�߲���57�����.SW���VTd��='Ц��­q�kˉĈI��U��1������㔶�&���_��΢N��/b�7�e׹�^����O��Z:�5)OBv�W�ȱY.�W�8�E��2TY-�^O�@���_��d��)Mf*����%���D�R7�7c
j�y� {$��9	��� �l�E��0��,�ǸC��'���9�{ՀKm�<>py�g���������(R5=
l�f-�#��~��ִ�Z��vX�c�۶YOz�v0:�-e��G^RE;�_T����F�� 1bs�p��r�B&�!�_]%���!+��)���a�a������8��ڹ.`_�f��7��Rj�I�6b�%%����c~��Pds��FɁedn9�hE,D~�LJ�$�XI�U�5��������*�W��'�`��s��|� 'N��-���F��H-�a \��A�:?׭3Na���\��8��!�t[9ת��ʌ�M���.,?Ll%š�hs͠x��l��E\dt	ݭU�E]��*v)c��$��u �@�-Eײ���\I ���Ehw#bƵ%P�������ߪZ�:��\9q��.�|�A�>��H� =�u9��>(�syφ����}�t/�qqACȽ���<����ܱ��5h�'!�rX���"����yhFnw_���}�N��)�hî�C�A85nSR�gVjϣzU��Dg r3$��Z^sm���A����k�&L2�Z(�P�,k��
,
���L���mMf+�ʹ�w
����4n�����W7�F�:u?�RኼZD���S��ȴtߋ/�{����!�{�P�3%�>oԿ1zH��c�3Ě�x�`�HXt|j��h^��k��?j8.�QCNN��R#5��ڀLx�]��0r���� � Q�Q�����B۾��b⎨�p�(��i�ј_R?n+j��t|�&W�����ER�۞ԆU>4m#�9����u��DPMW��À�Q��?m�	�Z%��qu�L� �2��A���}c�,��/�/��ӕz��p��{���\�W�഑W�$�F����64�/\�TjXR��#eX���2�-�0�����7q�x��%�YX"1��c��^�1F��ִ�F�\h�r���*|Q H�Me�����Y��V<:�4$V�XQ��H� �|������mX._$�m�MJ@jV�a��!���V�BJ5��}��w��{F,P����.��"W���R9H�[�H4ԕ������ЊN>���)�����n
�⾰p�J���2R��@jV�u�!����,H��.		�rK�,fP�,3ɺ���T���6�z�l�,߇�JR!X���)]�p@����Ǉ�<�%|��>�)܄��T	���A_j=���,���[�����z�鍐�m�R�GCb^|��r��	�̱R[Q�'"P����`n�x���cK�׋��R�p��hVݤfݱ���'��%�Ą���7���Pj�� K �W��F	�fȮ�ӊ4����Ѡ��u��.�o�􈿈�wSL���9˿�V>(_��*>^o�7��n�^��4]9���0���)s"H8�9Z�Wn����p���x�l;M+׮��=I��s�y�E)�i��Z��=5���Qu˄�r��D�����V���#o4 ��ǨL]V�>&�;�r"�rNILD��h�Uۤ�Y����o����L�{]8�X\�Nݜ������I���nu@�W2��E��YDM$�F�@�Tig��|X�%��8	����+b�K��;����C��؍��}��}�C��a�]�w�񭆐�`��|׃��lma'.k7����"�x��'%�o�"I`�� �=�3������r.����d�Cw��?Tv0ڷ[���v� �Р���1�v}вx�*\���{�*@ac�H��&%ы��������3j�1�"�ũ�`���7���6ak��W|�>��t��;�.ɰ�r����ͨϺ���~R�c/:o!ᱟF�<;a�u���2i�[h�i�MP/�u�[<Kޕ:a������X�$�Vݯ�����D���)Aq�A��q��Cj��?Lb����N��Y4l$ ڊتb{�r�azG��*tQ�P�**4[Ӿ֔��r��oW@~o�/���t�)�_0P�ji#���u)�~0�5q;�ʗ��X:W�nʥό��v��:�!W�P�b���v"3ݗ���M��Z���m�7�R�e)�����N���'P����VS.`rǱ����ED������:$��k�u�{�,\C4��7�q]t��˷r�`�o�N|-��Y=�00DQ;��,�o~�䁚�����k���M����=�xK�e׊����=�����k�������	�����Z9���լ��f�)�^8A;N��9���$	��a�G�.�Q�b����^һw��f��v��_�+��hRQ`X��RL	���c���vm|��մW�m9^z�;�#�u���+S0�zU��Z���"���4H�e��m���*��(NÜ����2�#�C�����Mϴ<����|1	����_d+f�hf~�pS��JeW�l�Q��uA��)����Ú*���+�C�.���E����n"e�N��w޿toxï��o����&�k�\O%\0�9��:_�����s !JވE�XC���3t,\T�;���LȈ9"V�J_���Q���T�$��ݗ�ϋ�I��]��!.�*aX�����҃����q�ɚh��mz�Ӹ h�ٷ8�WO�4@n��B�
�ӳ��c�5XN/�����n8��:ŨKA@��.�($`�ٶ	��v��8�%���x��MZ ��<��j_�uY�3��0�$D�fA� G�b!PJ��b��9�@���?��N��1��
d���"GR]G��O-U<�˛��^���@�Q ��߹_��.sB�Y�ʶg^ ����G^�HX��JCr�3<!2�w��c����[p�+p��u�)ni�8G"�1f���N�L�z�ݥÇ��|�qK����%"RLe��TS~l���yb%|�.��Lz��
P`�d���?uz�]ɶs�M�ƚ>���a=��yx;��
�d*i����n~g��t�h��E�"w&~*�7w���L����Cvޭ]>�)�b؞���v�ṨQ��wn��|'�UR��;�_��1d���������j*z�MN��n[����[�o�\[��+�1}���`�#t!���0��d�'��]�O�-�#�4
��8pO��Y��̱L�߾���x��J'I�DC�o�2���8��u�k�\~v��m,0~�,s���m3`�F�<^�w�]Z���o>( Q�F6��H�B��Mr�P�Z@�����fLqf?2Tկh�G�o*�
�I���3�����C4�Ͷ!�{{�*�qZߣ9tؒi1^��o���V�Cuv���ِ��;b⚖��ZV���$��^�rW���Ha���S��H`z=�[��1Q�'Ę֯���4����O��ND���X��0�ݕ`"��m�m:��1��mq���|��#�3ͤ��-��`���T[��h���$y�q�b�T@�����)��-h�Ok���
s�`���o+Vz�#V(�Z�G�;d}_���K������Bi@��%�H%��ł���`��lz1ר��;G�+�����	��\����z�;�4�?|KA�"a<j16�ٖxKE�̫���O��pƆ��:�8��(R�^�=ha�$`����7�rdt}E���.�"`�o���$�-B�C���d���&6�?h�X���)X������ ����q�q��	�0�Ԅ@��^�����m�3D6��4���r�������]pV���ޥ����]�$�j�����ާ�V:>P�E��Ѫ�m-X��s������7��3p}���\0 �-rp�v����>��7�n��ŏ��&P_$�y"�\y?�h��(��zZ�oC�̞�z����c�}0�H�Eo��:)���t�s�h�gG�#x���+<���(�p��ϴ���������)iS�N��P<0��s4�L�y �d�u�u3{Ɔ� @����&1��0X����[��>!i'�0z����Ո=B�-wf�G��{Lݨ�| V�r]�,��Q����FTC��?�yG��X�k�{�*�k�]Sm4�������D5ME����u�]U��n[V	_�q}pY�:���>��?�����]�#<�r�и���|�v��eX��	�(�� �O��4(�YH�_-rJZ��2��T�)`��,`@A�̆��ڑi4���6�����
.�Y��2#��(����TL�ݥ6��Xs�����$vę��
���To���XML�r�n����a�-7�ަ�$4�m=sZ�	kԦ��g��1�So����Pf�~��oMl�ҪP!bn@�ĸ�pE�Z������!q`��>4�c<[b�J̣�8/�݆	=�v���� h�Ω|]�u��)�zo��&�S�JL!�M�S2���b_�0H8$��6�r P	h �`�����l��9��J;C�9R�F0�����?Mf@'����A�Q��N�8���
���kZ�ɍ�ڄFAzY�}+-�WSЦ��$ռP?�{����K-.�`n9�x�uT8}���U?�Z�7S$Y�"�a��B���)��;��#+RZ�k����Qn��Jw7��C6]�����S�%�S��w)�iV_W�K�ʿ;'�h@�@4ӄ����H�s+�{�!6Tڳ|gǔ�^��9���i��"�EǷ%���ˈ=�7ʉjf�Ja�[>��)�N�/ߪray�>iK��g�bVk����"ē'z�j�w,����pc.	Q,�;Z)���H�	�=�%�3J��b���A�c*''��d��_�U����{�ޚLCKJ�����&^�u-��;�C�X'��|+A� �iM��i^*='�E���lz��a�.��#�|ߗ�R��1��h\)[��Z�4RydUB/���[���Sl\E���X�@�,s$hsc������$��"�!�0�Y
IE)�p�Mj�c�O����J��<V@���[4?[X	5_��69m����@� dP=:D9{O���7ܧ$�6��-Qa��*����j�)̿�g>�r�1c;�_�^��e��v5��ZY��c��F2Pʿ�X�p�w(��<�:�$��9�
��,�׋a���\�lQ��NJ����6ؤ��MjR8u05�L�,ɹH��,���Xk�ŀq����n|KMS���f	M�� �.<q�DA&&1U�G�pa>�bM��p���ͯHz�m�UcThG�<2��`]h�g��u��L��w�JFPdV���FF���z:L6I>��x��t)�9N���)o�
��!=T�� ?#���Ox�8��d�{������bg����"��f���C��֭�D7���w�
8G�,Q�S�5�(�U��ɨUю/�F�m�'#j�s����FGh]]ą񻸉E�����l��{�&!��^���:i�fҜ\�|R�l�(1պ>���*#���Jx�����M�hkC��IO�8\�}IZ~(������)�eѿ3�~DN�!V!�h��(E���3_]��_y�+�:\.�q fä�T)fx�l�֢i��d�5�,f��;X�;~-���LQW��"S2��A�j���c)+?��_/�p�nNF����H?蓲jk��s�W�G�%�ݑ�����{��Z�4p�Z�׆�?�q���
��K+S��f����^�(a�b�[F�˛`�t��k�!�ތ��x8�9@� �^���{����V�7��V$[�!���z�{�ZϡH��H�[�hGpF�]��H��'