��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O!) ���Y�Q΄�O��*Ȣy�dsuQ���`�Q}SA[�.���(��<
vɼ��;4���͋s1D[
�f�T�[��h�K�"HO�¤�TwƜ|�J�tR:����p�#��;������A&�K��HȮ�!!@<Ȍ��VV ��k��ko窿ae����ZS(�F�FO��2�;Z=��t�)W�{yo��r��(�K�StcN.�����s{P�8��AN�C�/��~Y����[#�z�bEB97�'���?�$'�����ِ��ǰ[�'�d�X�������%��`r��`���8D�]�At���w	V�򴴌���R����F8[4Nj7�-���ιFUEp�]c��$W��9P�|�Ԝ��L�?�9�8	^rA�Ƿ���.�He���n0�u�+}@I�2��P%p���-���6��f�8Џb̝h����喥e n/&ρ�1��ue��Fw�����s���Sܿq󀷀�	�~��ݒ�-i�Ȳ�G���S1	�g��<�ד��f�t0-I���:oۼQ gD1M隬it�;y����4_���TB�چ���thh�bL0���]q~�����4�Pw��Du,��8n�,�045��u�3`G��볮��"�W����`�hR�u��yI&n��xc���&����7���W>=���Ű��T��+�ς7
�73�ȥP#�lm��"8:�K4�j��c��<��d�eA����
���&c.�nP�	�hy�Q� ��l54ꓭ��ٶ���j'bz~�������,��������&l$� �+��D}�4j̢�0��)z���#ef �2)AuO�3�ۉ��p���s�l,��p�J\W?��sk\���k��}�a�.�.i]�q��W���o��9�����^+@���T�ӷ1m�$�X��<�j更�UGk�y��b��}���8uw�h�R�b"㕑I`}�0B���B��v��u0ۇ���A@��D����N�Zۊ5&] ����I��-�K���_å��HҚlL#��^�p�wo�O!�`'����^6y1^��m��7���s�5���"����BM�&+��#��_����'k.�A�$ʎ����ąI�4Nj�^��Ⱦ��4�e�zg�J �Ty�hL�%� �@x*Y�B��2��a�0J.�v�P=�|/�2��2��_	{ɮ���!��r�J�Eׅ�*ف!��#iݝ��W����hcmx��!�!�5�(,��t����3��N��7�v�I'a������LR1q颕]QK��l�ɧR���36Μ^�{Lcɬu'UbLp|&X�4v�[#T��d�uPd�6�)�v{�� �Fe2��ͳ쿙�v�B���������=������X��a:-8�3^j$��Խ����W�&�]fg�=�SR��!2X4���i$;��e��=[Vǡ'k4$�W�Z�?�hj������TM-�Щ%	��Gi�~&��ݸ�8k�qJ��]�r�p1-$<"�f���A�{�3��pFz]����N8�!����L"�8ђ�gM��ö���Vϓ�Ӹ�Z����e욦vxZ7�R��g��ʥ~J YU�a-�X������a[��ȸ�D�9$ԬJ��9w�xV�"�}E�@o�(u>D�q���)K���h�y���܍k���ٛ�o�%;O'�1#=�j��(5Ք_񦉢�����x5�;ĳ��|��Ʈq��e�[	����	��O�K���bA5̨��[�Zk�y���>{��$�)m����M,Jy��� ���sP�qi���\17_C���ekOJ�h+�[spA3����ᓼ���ro�7�v+�8�挝V$&���ǵ��v��(y��G��,�t:��ׂʵ�����Q/�7b���]و"=�p����t��o�oxٹ�����b9I��Eڇ��ϐ�*�,fUM�*���-�mF�/,uj֦k�� �E�b,p�}:����7�װ`7��v�U�se_�6�Nm��8��Qư��P+r([J����!.�c.�Fؔݕq�5�I�ۦ��C��I��@�>����B�$�nC��,��$}S$�/����"����>�¶Z���qXQtV$Ug�i�Zp�Z���u�ًLKջ�	;9�ӥЖ#�U�������ɏ�u_�P����bl��$g�1���G9ԅ��Y���
�|���d�"�S#}���$=�U٧�U���81��,D�?��ʘi�Zv��
M�����޿�°�9�K�����m�rcД�Ԓ�X/#ə�dPZ\�l�N�Lt,����aV�����+wH�� ���^����NnW�a�h�aس,�� e��RT������,�BiU��g�顮z��|����I}&+ q+���m#n�ƓD�� � �6�mtf����N`���m8�����^"s�va���}�	N���O�^U�Ŋ^�LH���o��<�bZ��"a�Ƕ��b�Vژ���7�t�/�l��=��7b'ƀ
q�l�����m��{'Ħ~�A1{;��&��J��8���K>~e8t�Ç�k�o/���B�Vfz�l7�U��S9(Κ��*xb �q�II`�`U���Hs�x�E�\�ˇ�<��e�։�� ؉�s���{�Y�lU�������`�����pb�
xx�ف!��)�� �"������_ �'��^ZW��&�����H���v9�ίV0�mǄP+P��A�MM�#_5��m[:w��������t��D\�w��n��v膱�=F�.M~{�����DϪ1hc�1�p����O �#>ڞ��P{v��U$h�%q��j�P��� M����a��Y]��\I�${z�t�����լ���G���L]��W��