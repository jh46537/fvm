��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�q��ʵǟ�07P
�����PQ��b+qm�ݘªX��<�Zwg8 b�4zI��ɽ�~A����*�N{�O\/�@>�0^�5��6�X0���-��S��k�sxm��(7cަ��)CP�����$��c��p�l��% ����':�Z�>��$l�T�B�k@�V6*C�Q�iA��r\��=�sܺ�/�Xnœ�{�DƐĄ�ل�8��0+1�ݎe�3��[��&:�\n��&T/���ˏ3�X���^�E���W����0� dJ.�Ys`J҉�c����gN��/\��S��$�VA���	Ɵ���o�j��Z�U�M�B+l	�捉��5N�\ݛ-�#OY��إ9[�c�KͣhB�|��s-�B��C��n �����%�߇z4����,�"	T�9�A�T��a��U��%�j*4����q ˗��_�R��� ��.,=��	�9���p/	�g��s}��}��U���|��	ؼ����EG��:��7�@�4	=*y:��&��	��	�`�aT<�f� ]�"v�0���e_gB7֖�BԱ��:�gKt[	�V�L���k��� ��J�H0�������hd*Ur���ӥ��*P!�
�@��c�"}�9�B��S��r�&�%k�Ӡ�&�� �/����!�򬁢��R�2}�-��H�z\[��j�#4�o�H��Py�h�䊢k?7�0g��L�V�Q_>�J�58��6�[{�.����>3�ʹ_S���)`+"�*u��Lp,2M黵d�"���?�ڕ3��f񿀯^��s�rr��t�,�0:�@4	9?��!֦J��j��dD��U��h���n8�ʸ�B3����r�?� ^C4�2�*iyK>?p�;��G�y���o!j�����~)���cD1�e�s������'�'��x>y�g}�X}�bcS?�w��;���E���� �.�T*�.4�)��c��/�5�pX���O���������f��d���]QDӶjM�dN.*���)�>z�#���P���fV��D�cA����exH��C�� C��
�o�1۳y��Nֹn_ԉb���bg<V,���T��N��\�L��8"�O)Vd��^P\&F뒟�4й�m�Wq��H�ýr�D�{m��*�!�t,��6��.1��"`R�aLr?��l�\�N�T*+څۈxt$x����Z;���ku�������p���O�Obr`�L���$��82�}V귶���<6����X�&Ju�g���<��>��A��d{�J�:^��&R71g�*��	X��r>5�e�RY=6ZX���A�},L?G2X��Q���c}Tr6�bFA�T�� ��A�O^�yk=�����61��+��oE�}��!jAc0�|?��fý0Ml��1$����p�jE��ֺ�G[�Q���W�iF_2�D;0L�����a�PK"5���O�B�
��F=�*C�n�Yq���GR��.��r��g��ɴ0�>tb����������d