��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{�.Ѱ�!�C�8f���A�uc��vh�V�,*��1z�!����vLE콾{�7�څ����{o/.Қew&����=�S�*�ٳ��;���2O+nw_
U��K�����G���Y�zؕ�Z;�^nd�\إ��Wz��-D�%�9!�@��l���#L�͝�(������H�J6�s>wʱ�/�*�� d��+�����<�m�hiht`C����^���F#�!v9%+S��k��ۙ�����0c�mY�:4�nv�EƧ]��/�s:�"TE@3M�_v������:w���:-�Z�KD(�#��� ���dZϴD^�%�
���(z08�q�wM�bW����5꾤;5@jM�@��R�{�8ɱ0���`CĲ4��ӱU��t��I���� {���{� �*j�d %�� ��utG�{ԟg"4R}�Ҵ� ���kyF~��L�f�݅|�	��x��~)[^J�;��F���n��KѶ�M��yH��/`�+�t�im�!̈́����G���OQt��K��]��ՙA��bñQ#���s��lZ�9� �]�V<�=K<'Ue���uM}�3ć�y5f��S��i/;�@;C��E&q�g�}Cf, T{��}�m@��+We&Si|Ny�|�V��T��gRv���c� �� �76!��)$����ڑ�`�qH}�v�����>��p�Lq��[V�\��D�9i���|��e�y��H3m)��/1���0�T��+Sّ�Q��I���y�/�B�v>��{�* 5<J�Qz�\Q�?~�(�!���5��^��9)|���^~����f�YX!*:z'�|�;�\��+�^Y*��x�C�9q��+x��n6�0w�B/\_$��A�C��c>G^���y�nS��B�,�٧P4��mCi8}-���F��ʵ}s�l���\����KϘ>�����g;���	�^���+21���}�L�{p+�Z�d*F45�:ȿa�|r�~tIi�!��g����hA�X<s6P��྘C�ܫ�^�]���׌\���es�e������kܼD�3I���:c�A�Tgn*XaE�bEI��1^���:2fI3�S{*����O�D�R����j�XSZ�Ȇ�������iX���~��p�S�����5�P�Z���Uw��绤"Vla��o��,����F��uu���#}���m���0K��.@j�u�YV\�F�C}t#����D��P�H�kp��!mw���,���o��I��I���lp�z[��?�n)x;&�՟ራ�`i�&�������/����<e�
Q#�m]���)$"+�	�1]A�#��Wr�"]�X�|�t9� ��fA�M�����Js�jb��ƃB�M���$.�󏨖�� 9 �x�c��դ�������li�e�2��C �&}���
r�.Z�Z5i�f'q9_��E�/�|����"�<�u�^�Cx�d�H�/8ngUԦ,�m��1����ǜ����ߊ�5
@��#��%���y�"�ǕwŤ��0#c4�P�
>v����T�i�Lɋ���,?�����o�,	�`���U�R!j�U�;d��-\-���ٲ��k����48!5&��p�["֛��n�mZ�8�*Ⱥ�M��0t���H��No?
�������lo�&9]X-�4���8�l��U1�S����@��+>)d�C��� 3�'���\���d�"��[s{�T9�K4�\��3�$��� �еHh������U[�'�lC�#��j�'ۓӶ�����~AY�h��A59����in�:�L��C�D��<&c �y I(��x��oM5�+F��.I4����;@,�Pa�H��I��6(���-l�[S�A���{%S�)�.�Y�j�9�Dkժ�6�w��
�S)�a���{�<]|�6�޶D��^�ö��zO4'&�NH�ENCF;}��;o},�)Y��^ܰ��/'c�+�����Gz�x'M֖��M�!'�y��NLxC�~3Az�L{
�E��2����y[49� �/���79��(��,Բx�t�5�b�-���@۝��#2��Es�n�q���>]r�