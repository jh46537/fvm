��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�=WM�Q؅T޺HݱCV.�gk�i�E���l�<��H��n���(��!��{�?�D6��'�]
���,W��vt��a�>(d��j�@[�ȅ�j�U�@˝�c�������W��;���;��=��/с��m�IHN-������#�g���]ו����Z'�����WTc>إ���8��>������z��K���(ޔ�����(���#ى[�ݳʥ�ۣ�&Z��,@�l�J�#ŕOKi,��=�������t��4Br�ٿ "�W$�"f��9��S)�_�Ϧ&�����yn[�.�U�Κ��33!oz�"�`f�_�v��I:j;/�p6`D��Ӵ\uѩ~�5"����~�v�u�ل����I�k�a��enB�>����V'��u�E����KY,�&��^�������'U��P��ѬV�G���1A���`Q�Õ.O5�<������g���s* �=�<�2��h�魱�ǠMy�g��(,J�_W��� H�Y.�T����]ܜ@0#�GD�!�&�-��U���߃�?j#fk�ʓI�n���?g�؊�k��^�z�����$��_�Oj
�:�K.��Ѹ�σ=���A�^��"(��h����w�n���3Q:%���Bs)")Wtb�:�L_f���������p�Eqy�xф`��@sսܹC������n�`�o۪ZS�L6{}�;�r��-n��<�2r��Y�,�vBڇ�/+�����(���?$ �;�{1�F�9����������ghv8�sM��n9ۦP7�4/i/�!���V�GV���yx�{ �$M���e`�����{똃�?����h��X@�7�Eh�6^(gΚ�+�\͏1�"b(�:E��0l�+ݎ����n\���z�?�`t!�p�V2�I�O�hA��؍!ɀD�3��\VY����o4�Fc�rY8�����*�,�Gu��&4TYj��ݕ��E>Y�M��|�ab^�.ڃ����"r�D�uMf3X�|?�b6�o��U��G|سT1խ�gv}i]Z�*���
K�턥A.$]ɒ�f�B��(�q<�N�8��f)��̋ZAKΣ �Ν-x��b�*�ŞC���g4,�e����)�B�=���s���W�!B�G��5
g�����E����֞�R�^�;a̱�Vx�N�Wԍ&ƫX��O�����i�܍w��ҩ�[8+ZVkc�uE�e�6?��1�Z�͔��DT8 M�jռJN�2��\jX��M3r�q�$_#�d�'3qm�N��d#�dDfKB�`�	��V���к��6��-�%�RvY��lӂ�ޡ\J�~���p�q|ӧV���K}7���R��㹼_����x�����Ȧ�����0|Y8��5\�׊d��	VGh��������b�n�Em��:�R]�@(��Ζ��ڙ�B�$�QkbnL~��j������)i������~�y��qa��C�k[FD#��U0[���u!��h7�����w].ٵRo@��sb�;�Ϫ�=z�]��ؼ�F��>Y"ǒ���IHdO����*ݒ��HB��1Y�1�qmt��.�t�͸h��F�{�k6����U1b.�`����g^���*<#��:̋=sA�<&a����&1ƹ�K����l׿�G S��ܟ��XſQ	s�/���;�Ը�8|�J��.b�է�q���_�D~z.���AǪ���,�����k����rz�"x
;�-��P�-�YVG6�6kT9���4�1��8Y1���d� Ys���',�3L�6��r:J�?�3����!2B :��ZnZ&����1���T�[����33���(�Z�,r�P23�F;0O�z�
-8�Z~�Z/Ѝ�A�v����q娗��S�K����؅W�֫�?��b��"'��d/�q��V��ډ��O�ga�a�^��*�h���0�ܹ����zݦ�`����/-k�����N��db(�gT��k�h���O����ol��,���#k�tX8�[GL��H:*�1��ě(Sܸ"q!w�#U&���ZI�~g��ݸ��6�ФO���owB)Z�M�����CO����,�;4�&9��!Fol�RB�p����=���ک)��n���7���i�6'SP��ad�����������'ܘ�����hZ^�[e�U��3�E�_BºG�0����s�_�A�){4
�[ǎ&/w1W����+�w���) �5s�j�R��tA,���ľr��Ea-i7ް�w޸0��1�q�;A�)�f�*�����B(�~��dJ#o&����B�I��~���Ǚ?��~��zW��^u!K��p5�[Sw�+>��Y��&�Ƕ�ڠ�1����Fk-�93�����GK�B�.�;zw��h}�)���eM�7a*�|Ԥ�S�t��+WU2�I�\(r4�}U8�z G���|��������$آk����j^�
C��F�3��i%��xP�L	�����p�f����n:�*�r��v3��r��NF{j|;'�_�L$lY_9\�����,s�h�ua��dX��앯����h��TB|��[w.tip�f7�9�.���_��Uk� �b
�L�=��T����� �n\ZsY5��"��h���Ge�a���;�A�/�
�VH�"�.?5�;?f����V�忖(&:�SB�+�[X��������;���/ c�&�*�;��>����|�����L�h9�hel����]q0�9ގw��^o ��aD�X[p?�]x����h������ R�ϰ�2k� ��)r�~э�\��G�\B�g0�҉g��q D�w���M�W���\��$�Hy MJ;{��TE ��k^t@��w��B<�`A_S�5+{�V_Ԉ	��r/���S�A�t}S%52�a���+�#�T���!C�/���`���5�9�5���THe�t�"gf�^�6���xrҎQ��Әb��*�S4��zm�.RA9��xv.$}�HRB��^���b���ƃj=���Q��ي������� }r����T�yE@�O'������ʠ�ʉ��
hƈQ� �]5��\}�GoڹC�{KZ!�	���M��S�Z��]��-?C�Õg��z�˗ǜ�"b�qqP�ǩ�r�'57a/��~,K�0���"�������#(ψ&+b��uX�~#���u¯���18E�SUC���� ��lgHZ�M/�r�B�ɿ`������5(%�,H�X��\m�ϤQ�	PB�k�QV��h����fp=2���7�Rz����u�a���S�Cת�����D暗�)
Ҝo"��n����8og�wpj,!s�G,��$���܏�}$a���6M���'�c�n�Z̗��W��/~)�HE8�*���"�V
�?���LrW.���E�����\�Hx�'�c�<M��͒ @,�tp`E��������HP�6V�I#���ЗT�ԭ�q�H�:l���FV�z��Yxs`�}���Eٵui�XEӦ.�$y}'�iq�?H�e�5�P���?9�.'��]ߘ��H�/�f�=�4��*�:�5X[��(iQ%L���x[.�q;��7��\L��`խ�����*�_��gx1c��=͠�S�gp=JQ7c�����8g�Ь�(<nⱏ����8��8�='��F!`Zѳ�W5	h��r	<�!޾g�T9&��1)��6[�&�������G��oG�{g�ݠ���̬`R�FE���/}�<�m�`N?��Пɹ���&I͒�tq�=e�b���:t�������9��h�k�:�i�a��I�f�,+�p�e` �W[���y���D�9�dc�5-�nLEx{����`���
c��:��Fha�i�z:~���ģ�����1�؄��`���u��>b:օg���R�v�*҃Dg$/�N6�<~�^�޹�L{	����4#��-�	�C{�6�!��C��r�i��p��^5�&��_S��j`Eߡ�1��8����ԙ$�´�M��;U�z�I��������#m��Hg6#=a�p����7���������f@֛Jp���O��n�k95I��R��M-��Hgq%R�T���s?-��'���H4_��#�~+�!{�����Q�\�8p+�O�*c	X���������%Qr���^��wo[~�40��� ����ƥ��|5/�TB�S64;����p��j������EҪ��v68����κ�`^B�m�#GG�毱�r xMRL��:�����(�sz���c�;�.a��%K��� ��ގ� ��^�i�/rS�Q��*�bY?��[�+��#Z�@D�<*�?�]�D!��:���{΋�_oէ��/��Y��F��-����F�[����=�
-�M a��� ��ʊ3%3�w~CٴUZ���|q�_%�m,P(�P�[[~��\���P���˞0�P�ш���yS�JM���v9c������t���G��NG����+�9w\�F���2��T��6�u���6���(�C�6x�$��u�m�F;ŲOˀ��� D�Dm�h&�C�l���'�L����a?�Ƕȿ��G�[f�Hr_ef�ukB���m|������ܡ�g��Q���#�r���^\P�s�{��vuUs������_� ��	؍��ԋ
,t--�+ʇXR����o����!l{\�
9��^�) J��s��?�����q�d0����^v��{�Ui$�o��
O~�$f���ӧ�Q����)�gk��MO�go����q����ƶ�!>}]����LZ�"��x4�6������\�0u����7���ؙ:�?�J̃:�is�u�F�6B*}�γf�K�a�e_����t�=G(�-o�E�z�������D8�p�����3�,J��K��Șn�f*1U�~.I���u_]��E��$OॢD�'�3���P�'ӱ�0�.^���li�K'ٴf�9������e4j�T�*�#��t����ϰc��$Kek�o�C0�k�ї9�7bewԊ4-�r��~�_;Sme=h>�[�<k�[�0{�v�7-s.���ԯgi�B����
ٵ�״*敩54��x	�#�k�Ezpf)�