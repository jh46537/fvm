// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:53 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ihjx9I2Sz44i2jc0Y0C4LkJPYpAPZmyQIdKmiptvpC09Ghhvu5+lcQwkXFmTiOhA
0JxPFxbtV5Pg5AIaGPUXNe6E4B1ob/6vKAFy1DHgjzskth64gze1BH78pRnlYBxN
MR87vlvHBoRicj3Cu2yzbasbEwRm0iUOfbIf55911nc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
iN4zpnXvrTfdlyr0T4J27SxYWcIVjpJrkex8Em8vK2lPYNkX2ysnp+xvF9f3L9Ol
R3kW4i8bkQm5r1gIpptbT4XB4+chjWNQVY05yDrC4V1uZzqake4TGQbGJiBr5QMP
dKqBe22AG504M4izuRpeXiDqBURnxDFhkUnAo8NSuLlhJTUFIyRab8uYkkEE52xw
TmbbfGMwTzU6jei8WvKbKZu6zht8itUjHySM2Fuju0UCjdHziKqv6OQ5XFoub6gF
1WCIE/Wp1GttMZ1BpDPWSPOSP2lQI5tJBZfXw59ictjt0oiyeClmYGn3WibZfxAN
/ElFDm2AIoNU/Q50nKPvEUfOA05PmGoZkfODee83yiBjATBYMYmrBQLANzNVrRtS
Ej+9LZTJ3uTxmEcNizdRxsLy4PwbQq0mBd4AlBpXpSKlbfYsHKPWwUP/QYPIKNLO
JlYZc3g5k5hKx3gtxknxymFn5MGjz5Oz/7WEHfHXyejI+g9OQcR62JcWgJYdbmkH
VkfIWHtHyYz14E4e4L5DL2zDRu2i3ufz5YADlPLQfJLUdg13lWbNyAq4oV5dtBd+
s7dIJhwgwilPf567fsAOOfh2UV8Cd+uYk42h5/KljR4jEhPDXosIIEO5DSbCDRWK
XQs57OBXl9O5Gkm5wVVSF9ei2YOfC4DS8kVRWYOfqykXXF8bqljFaktx1A19mJb+
NB2iUvoZr+HBPVX8xaXJmGHVqRc4SHX84z1SfMqAsg2+IUoKLwyVmdS4xp06DQG/
c2SwtmJn0SBkzt3f81255D7B0F/iHSdz2dGHIZNXt4VQ/zFu0OxPMkj4uUoY4jv0
5ksDgJXNU9Ot9rUc5u5SgBxxV+NznD7loneDZw25zjGcItxmALDXzRHjE4mnJaNd
MqQFUK6qPJNzhCBSyPsPq6WXSATJRoatBSuOsIAdyYYSy0XVjopqbXHyDZSS8d5T
0++5OhCkEOKRvS9weg01ouJUgtev7VTGkp62ChUqyA9yR01bJrarNqsezeyIXrNV
OMsx61EXMixO98BzEBUxFIvQorAf0TevR4/nK9pMfEjPnwpE9gc3Q5XTBt63C2l8
HiPv/hctI0YQ7sCHgJBZmNJUhHih/1BVPVYwCAlDbhC748TZ7VhBwyMGuw5cevLT
AIejCoLyM6i+mzJixu3/YTjL+pod2u0sunb1w5rZqW+Ncp1NH2EbVvgZUG5NfjMv
7mJd0JJukhQQIUWwaZJdx6J6i9MtJAbxw8AZaRy4SUQgCe8V7cIpIvmoa+P0S3qP
nZuTHhDCeKWZVJ3CU9HPUN1zkHJurqLwp4I92/giBzgLkOjJJKQbW4duiOGrcmZN
LbIEFSb4LYzAyijjlwQE2yoHMOfpPDfeMFte+nhSy/n90+yC1crMtd84ECEKv/Hz
EWLFqlOvc0EnwiCry2r2axnK5Ci6tJQCgzt1fxzUaLvXWcf38eWrxB/ydDNhgwRH
QbwdWWlJ31NMkegrmopiYTLyrvkpVlv+D5vI5lvERpKV26G5mT/aPlCnSvchAXhA
5RcbAXXVKAxrw/eSTU70IXLjHQI6hEXFvhvKM6EFzESjYb9+J+vrLblOTISClI88
ERhTBe2Ux83RLaVWfMm7UcXyyyQ2atB9nq8sO6iT0tMDajjDLtt4cmRN09wal8Yp
6007PI5+Z8CStknFaAWU/HbhE5n+NInvBCiGCwR3LA85gm31zJGWbM3saDQ6oALE
tJIhEG3u8EMkKAVfPNlpMn2vpQAlWp1J2/ssXbkYePDcW5kJjqbLqSzbcBZJJ9wQ
2xsQki9fPLSmoEGxA+SNooFbvvK2SlqAR7bGQjmu/iZiqbu9jNJjmcsju949uOz1
ZCNcx+bCZZk44nsek/wUJf7Gm7Ldh72D2X33rng7V/LQaZei7xSZph0YK8A5nsWF
qxqgQZQ94FLILtev3QHJtvsXiUoW+k05Hv5nEKbdLWIov2Rb4eaPqbk/S8My7kUW
da4NspqvrhWEPaN67x4+JYRDlvNoE4AK2KGGJCTh3ZgyVu91m+Xgy8Y0bccyy+kx
ASO4NHxKZ/eao5sqEtmF6I8kYMc49zTmp1zzWMMZKdGq5YCAydtXNuHXOzx9LIEG
PSeg0XzTEiz2anL3/zkYCRiV4ylJ3aY2y9NI0GavTK5J0JuesrD+WQTBTaHgTUWa
s1LPnaNKIDEnYMwmyk7egwO2A4VvHcuekTGPt6YFc7pJ8jM3rw6ReJ64nLbRPhaz
n9jrOGaK1/JHE9vKMu7A4m6E2jBZi5ugfAuKzben3iYjI+ido1P2nyVGCHzzjAdC
F/5PAZxUrUFNiG/J+HPlc4S/KuilI/6bRjzEHXC94E5A9jAwoG0L/42CXznID48D
DAlKP6WaVWlL4uxiI2cvSpcijoAXsFMz5XkqRS6G9/hq0gtN9G9TpKFa30emvQCd
l4RHEoC8XqGCG4EPXgvnAWQntf6DKcVzDu+9sDqYA9N3sovqbETbByc86+fgEyJB
tzUP2Rw6wj1dxlwHKsX3uoPjvR7OIEVqQPhVRnIP7FT1xmTQGlekNfN7P2YMI9yz
nu2LGJ0KLsnqBnuGSKrjO5msaEwTvhY2yW53vB+ADghY7xJ7PL3dcvRiuGD1WUzt
cOskP7lGwnt6yJMoSClDxMwVPPIPCjmSgkZD1mtWLAolJ5FHNqbKcrCmh8tE09Kv
Y2PjVCDGxU8A28koJ7k+4zsRV3mlwURVQEAtc4+XH5YtFk12dUVhjRvDtGfAT8k5
0KNAGhJ8QcpzYsWw4f05gKvsBm/o0B1tqe07EyaPboPPoRZyi9A10cnzOwGaAgpo
Nbu4sy6NOB/LQvCdK29tgEEK+a9EYQ7cKhQ3qmvjA3BYVnV6uSeod6Qh8/JGwKw2
hZ0QfIlXBiQYEKSk76Y1X2Out7qLDd+7Ii30gdwAERXjumFX2VrNJ/mhNRBQ9yKa
AIqKLVGfv45V8OTH5BHVfIhs23UimyvSpR5yuETjaYdJKClzfbMxDRKKhh08Zfxy
RrghCb9229G5seOW1Q0g9bmzvN28Cw27SS636mmDsd4bQucuhVAQvgM4KihCNwQd
3c3KEV2nJYxsYmy1e+f8PiXT8RhvVC5ml1AfLBmyqMgXsIcvr0/V8NTqiHDYmF3r
SIrsXnMyHWusoeCTb+XB4nOTq7x71/Ls32B90pFovOF0trfjykcDCm3Izxg4UupF
n5PAkS7GLjaIT9xmMOinVKwx3OtbuqtWzTM8e+d/OaSoN5BG9SEJRY0qwaWkiLJ5
FNE/XLXovAKBKLWaGnxg2WRterDwuFbg8Wel60FGeBeTl2WXLHkUMFC+g7pfQBiH
mPTt0iaGRxuUv9nJkYAocUhACIb16A0p4YoC+euFeBy5KXnq3392k6l9FlADy1bp
4qppLAyagZXscoVv+FiGkaIUhUmuirkY76bTqsW2qNaw4ZFMnUwga6Pcz8S9yOF+
nhmMYtfjkMb4TbvCFd9JPzVAAP48Sfnnm46IyARFmP1mbmLqq0gTlKoXD6EREbhT
32S1ibGColvVZ4mGMGlOLMgIVLvdXPXeDrvmnZxKUo2umBW9v59d+/kb5Ijl9NW4
Y0qFfYrfTXRytdZ9yuAgTYGMXX9PWVFfJtj8FavmuW4FIkUkSGuzEQ41iVJ155QB
xMzsF1aIHnbMb7CVyKkym8re1xhvCjZIUxdTv7lCT7I1j17vmSaBmYyF2CqJ/5aR
9aqPe1hg23DqJhyGzIf9DrWC7/R3YXkK2ZXBZSYnbIaCMOihQyQj2Nq8OU/OYx7A
24Qs7kv/HwLQwkXcl3/XJ+FZtqzHkAxWXtjf8Usf+tQ13WDGuoCVxFDf4QP7l0Qc
zHGDfRzvvpZqw2XJtsaod3FnnV0g8tTl1zBLC5ztSxLmA3H2Rwc9OIC1KK3fXuPZ
r525+EWza9P4km3GsoMCiP+VdVUrbPR6dNpPjE2fe/c2TIw2zr0yqlbNVqNjC/OO
c24IeUxhub8fMfYYhOwp0/DaZK+QB8HrUkWxB1BbL1IUzLY2av7+sQu4GaKroWWs
uvq8671Wo9f2t+Jde/eG6K6qA6MGNibAUZt4c0B+S+X9sZnPTi51Tge5iVVLJ76m
NrUmv+AHT6CCxA9jcORNq0VMA8s5BiJ2FzM0573VXan1XhoQ0FmyGKjV0g6726/C
S5/cqYMW70HVqszlGqbH/oORrj3AAO5B1ow8GNaft1128/YHFsRilzUDHfkR+3lb
QhRjFkt5IRJRXwUX7nO9E9HYfY4g2GWss7G9bFToYv/c3f7QRbx9DZg2Q2B6j+6e
qyLUwEypP+xJJt/HgT3lejsgmnFBaRXv2Eh9/R+7dvyQE5Fu5p0bOhZHJqmt1N1A
7K8gQJD1v1t3Sc7ychzpUTcJHdWCWrjudU+CABas8QKmEywIDLF7Hx0VNkivKIEA
RaBxMTnqaX1rM05IBp6lmL5GmasUQghL4bYHU7QBNx7sd6cvdRFmhWf++KIlV7nc
jifS7yl10Si4PgaLhowPAG50CrVWzIK3CzFABNLnMDMwpMHF0MDVv/Xf28I+BqBg
BoaJlRnX/dcWGcKgBLcaxHQ3PfZA3xAYm0uKVVvmeEhwDBPmpJo3g3Lze34swUto
Gy5mUy5EJZzYaw8X81lI9/PslQMsQQbtgsqRaPmRzICYTWanLe7Jp73fta20Rl+t
Ct73t7RzkwWTo80vZOXfU8iMRGRzv1LUiOvppYkXoqsUdqMq8OlGS6IAnX5zbicD
i+F/z1AYDUAK3GERenyVdr4xRRlWIow8jrKgBMDC8LR6hoct+7eI7OmIUgY6QMDZ
+dea1Mooq591GBMTu4waxUdcJQfZhHucT7bbN4BuoSo/AqP519hPsJbe8TPo0L0e
6wisGBryKLPPOzk44pOK5Z2xGE3wwezBxQZF0A/msdtg80+RKx1g0+u33JoBW+r7
pemmbQS6YwAm8y3sQTDHbrIegfeE2HJcAbyjS7De5NhhWdjsf4Tx5wYmkZCNpK/d
cCXkdxrnH9sCDJx1Vd+2xn0PpKWq5DY1dWAwWLI0lVWJUw3VNGylbC0JaOOClJVn
uaDmpyl0FDMCLIVPp617ejyy2x0XEgV7M4m/y85dxS5+X8dp0FzILT9mfvoPPiYi
ILvY8F216RQMIFm4WaknWc/KmekaqTxORgYDs0tonQ3bZt3QZcK9g+PeYv3rcUuG
GdHLvHIRk71WoCGJpKK/aP/YyOz+HQYNJ/+hKzi6dBol6oR+BENVjLz3FWgL38fl
R++DBNsLWv8TyQ7z9af9tfI6JWSYyhrXNc2f48BQtvwyH3Xnb1ShEiLY+gYD55KJ
t3o8DhUohurmBexY0kz+ToF6lWD/w8pFyhXYlHaMHX4f94+q6gPUJwBCANPjXNnl
iPGvHvNQkIiubzV/V7RSwJItj5MC1uwHHmkycRH6Q2W215FbEYj2AGsIE1nH/v5U
OuJ+RoLDnZRKs+Plp003GQQOeEyMKTeNb3pHaG9THvnqY12VEGLIkFFhUaMRd4B+
weGiyX1AHKQP75nvmRZzPjnrvjcq14X8JvzkSZ+XlsNTdmIOA1E13jqJJiw/exDA
JVWIrrgZ1Hvj8Qv0azGMnXFDhH9rPWWwvZabxmlmpIqUZwNs6mtggoIzhSBHQmQj
j4I9h9JaCN5GIAA7UoZIsJ8mW8UmAr0/YOI++KJ0sBXvS1ivrTTZBldeOBjExhfG
iS8qLh3mJ3sOBc+cWhR9L8HSOIxJOr/sBODJ87wXP7zgEw75U8fJrabli0bFM8xs
4yX18vSf5iB1wJ0MHkPdk6b4nxnXg66DTGItGWz0iM5nTivDEykiD+wdRYRgltbS
ujM4E5/AVaFDvLx2+M5dMM278QgeNvx7K4updMWnKrNphi9OUpRpeqTqzB0P95i5
yWnpGoJqI+mm7/O2ydh5vWyIknKZcqS+kB/HsKmUodRXQdRBodnbx5dk+kxx4EiD
QATMHF10PqxzYeIJkkABvMv0a2+sLfIPInCNmgZOXXHH8DXHYww3FS8fTOIBbOy8
IpsYiwRjoBVd5tWhoGgNg/RvWf+eTZMiIlAzGm53kHKo1R6fJvLgR9CVgkV3yScd
ZgvqRho5GwXTp2YqwzLTREH6+9hjc7MlKWZ3eZPe8jKPbFFXbw7XV26TPvvIyECH
A1wMKlEOHMHJMtaBxjx/cPHlSvky2I0umJm7DbCQCdB3fuM+aDfILRgC6G2j4Cfj
cBLmWlUEZgKuayK3e+cClv4EButBzcSo/+/RBTNvu/NcQjtfSb4GLWc8r7CFPfsd
2jzyQyy/AAtRe6IZBnlzH/XD218L5ct5GZFX9CKbFVsSBypdM8TADQ1zTPpmRqbM
kCdq2S/9cF0CX/iV58Db2lg4kIpMBlywTyMGPhrDFSSWjAnQ9IXPSjfVSlRRCKaT
nHf/im5PHQGZH4RD9Pc4aapXHJtIOx1Azd5LID11mjpAvP8jvkviYTXJusWmsAi3
vtLo/QLCgPAV+TGZyWv52+nvlOyQxNp8lvra6JmirtWZod9ZgLyYgWaGrK9ihAXS
YJ7DHoZvVRrXgDvyV3Sk8WQCummAyI5UNI7X4QKjNM7mwzt/vJKPJCbdW4zAQBqv
33hrx5zJG7CNqtTjlQxu1f1jB+cfmTVPPtwwNUJMfEtioivBpzvggJGKgI39YfC4
nWIgGr10rve3LBXXhTG1g3AqwMOLkR+fhCqUTcrjYXvqepwvakBjPHzTquDzvyw9
xsRgXRpHySHT3qPw92Vqfu9Ci+6NRCxgo5XdBo62SNcoppABtk3kpVl+TpJ97H6b
5L5VhPYeS8blyCgkB0KEhJbPx/ueRkuuQVe1rZ7IW7N3/sRY/qwfjUt/Lo7jRx0Y
B5Vs1t4TQ4P5jPVdOKr/8uSylqsVgZ31piiQhtV5u6/Htc8H3p1ZvOvWcCtnuelX
C/yydPP4oJ/4g9Zub6nJKWEvAbCrQ3dtf0fUvY60R7RERJbimGPthhFmKI/axDWQ
fuw3+4MFWwN2HP7a6KKFPGB9cmyEs1Id+DTYY/EDL3Aw3ADtGOKgU+4jot3SNY0d
PBUeNyVlEOXUhJHN7gLLdA+t2efIuOQ9jedWGNIL1QjL8Q/MPZ3X3yytW5Y0GVMM
TRBcArt0FF4tY9FkkcfPCXmdG0Gd9Cceix4A0NAmhdoCTWWc9Ot3kTsHqkhs7e8I
tUZ4wP/hWYmpdRauDUu32ph62X5y9/Qf2ixZFrmozkPJQ4lgTNHA38fHCFhSk1jz
302leqUrPstbZp1N0inB6un7MpBLFQlsosoXNUms9GuveAxMB9D3YeeVuVzW3G0G
xtdBcT+kz9HIq/OF+k12uLdL+J6dEnsn4aK0zBM4Muc/3cl6D3YvT1mMvVOB7o45
nro39joQAOek0A4lUjR+ufvuE2Xati9yebzNgvXJyz2hedkNguH2lICgmhln4dq1
70LyrDYJnUmFETUvhm7QDhEPLTHjMuOiiUocwwnhQc4UP8ln/t2jg+qFQh1Bp22v
cK0EYNneO9+wn9hDe7aZqA==
`pragma protect end_protected
