��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%rҦ?��*3
�cӂJ^��iAO�*�1L���2��uYJ�c�P���H��Z@���즌���qT��B{=��ɦ!���-�0�>��?o�d^��3ݫ���z�`��ţf
6�k�t����d�w}N21�Ԏ5 ���XP%�9 �������W�����ಏ��H��lk�T���ϳ�;���_��8[�����Y%#H�<���jwN҄��-Z���[*c���#��c���n'�Z��$�djZ���1=���?���*��)G��>�bpW����?�|}�����1ֆ�l?��<>n%/)g����E�L(�R��Eo]�J�:���ؑ�>�!&���0c�y|�=SI��{�ǽӉ\�����DB�p�#��a���j�����z�2��s"�jk ��}R�x*�$�#��Y��e ��HOѭ�V�Ю��"h�M��
錤/5-b�曅q�Dd���I���!?���Bcl^��*�ƀnq�	�Luዝ�.hΞZtp�
"nl]#J��_�J����4_���9��!G����!F<��r�w{ƫM���� �'�:	"������t��n���q�^� �����Z��y���u��ڀ�k��[���R�l�c����o�ND�K9�8���%�,�1<Hݿb��D0�d����d��ʣә��vƁ��K|����*p�*��JU��[��/�m�Jkz�t��=<��3�u����	f�����%WyN�����������(]��~R��k�r��u��h.n�L�0پ+��~��G���C����U�w+�Dq],9n��-�o���8���|�%4<�pG� A�U":߲��j&BL�||Q[Y��'��}Sa7h'��B�_�#C%��]2\��%��1-b}$q��kԙ�?A� �xY�y\�ts+�l��g�g��kT*�zEٺȪ��Hrڄ�ZV9^��d���m�K�]���~��ҁ9M�c�Rz�+�l!��	��x�� ji���5UqQ{֥ߓԸ[�&@R�k�b�����b�A⌏�"\��F!2QZ�)����}FXу֮���7l޵�,r��@o��kڒ��%%�$��@�њ�v�W�]�O�4���׫5\�{!S"!xu�onA�.�<��|��C�}���w0��+��\�~+c������'�F�[t�ν��q�N,�;����9�R;��i������Hnl�T���t����cY�����}(�L#�wŷ��K6[����.�ۼݨ~Hp��/��O��>m�4"�zk�յ�e|7;�"�Q���T]^c?^�߯���Ģ��!O)S2�9ٯy�?ٵ������Ky��TP�˸d�x�W��.��3)�E������M��mB���q��C�(���RЉ��J��U��$Ho��� )�*�$a�'V�QM�Y	/�����2ӂyP�591��,��:��lC��b^T�$'ڮ�Vhצ9�s&&`�L�.�m��9S����κ"�?kLQ�(I����`�`����5&F�}��˹Sp���S�Y�֯�'�"Y�)9;�Ehl.B�3b�`�d�-�1P���'��%Ƴry�?]�<Ѳ3vw��`������D�KڴB���(Y����{���[p2kr��|#�KY#c9
q����/�3��ȹ����L�QC��K�,l;�\�Q���A=CB|���y�X������"��^�uxge����o
j���`�R�2��Y�r�)s���%���/�%�~���� ����(Rb�!���7 e����4�Y�]4�!�&}"����d�]d��s����!\oG��-�kS:��$&r�v���_��4v��-�ӵ_U�.B����u�ieҌ�pb{֫FRp��wnpxT&B�l�́s�>�i����,Oȗ��e>����S������gЊ�`�pn�4F�>�X�ÇR��xz]r��zB�ekH'��.�N�YG����W���z�E�c�#���x��	����� 
�J�����F�,�̹��hL^�c*��sS.|[((_0��)/��������ɃU����_u�/�K-�m+���m�w	�"���	��K�w��?i�7PcHߌBQK�X�)b��a�c��%bGv��Y&�w�z��roBn�i��w#�ȯ��>� ��ϖ ?]���k� �=���YAD��=�~�*����H�^a�n+2�-�����iS�:���ݷC�2���ܠ�HYՒ},
7��K���拜k�kLC��!�'���ZQ�gVi�b-u0;���@1X"a$WS�:�a��N�!�V9{�RY9�?O~0��\F'j���u6n�Fw�9
7B�7�H}��S/۟���{��y&�Ac��+&�3����i�O����TQ�_;a���[��U��{� CK!宿�Z��V�ŵ�_g�А�[�Ãh���e��	r�<ƻ�TZ;c���N��+q�����zWA�uf'����`rjS��@`P3�����b���	��c3�T���z��S�6Sn3ũb"�O߶5�Q�FrM�+��p!�@d�dA�����#�y��+�ڻޗ��9<͗�'���z(6�ĸ��^�9�C4�	���\�߾�<�ݴaG�i���
������*	]pr}�RG 21}#*Y��C�n��n#��`2P}h�_$2����X �amrldP�T��R�U��=|Cצ���p# ��S�5�A�ⶑc��v;��"��k>Y�t����>��Pb��ox@����J%��yR+g�Ȃ����0lSiVEf]����~��
�Q^��PA�U����>x0�07���*����ۅeT�E���~e;)�w(�S���,�jη/��-y:�,�2T��W�������V��f�f,�/�"�{1�^�C�n��1��] �i��;�'K�x �l�Q�]rZ�2?���\����Ș�?�ʢp�`��P�<�[N8�����^�G=5���(G��P���%I:�6&����|��$�5Dx33�y	��@X��:��H��|J����T5!s�u�d�N�J�8n�٤%QO�A����4Y�^��^����u�^�g%��7ʜF�g��a]x�A8��2����M٘:t�\�^Bzb��O��hZ=���S$m�1�jq��ۿG���6^�S�嘥E_�Sr��A:� Jy�5���_������R��T?�Ga�4�����"�
P�#x(�.���ϩ�����~�F:���.\�Q(������A�)s�j����
ƕ�����◠�u���h�#�G&b;��njҁu�H���3>a{��@�E������Mp��)�B&W�t�M��I5n�����ӿ���lj��&F}��_���.�0�@6�j�O�x�ޚ�@KV@k�m���Q;�D��ϫ)+k$�s�ʑ]���`v��&6�|��p��|8>
��k�:�jPa��JN�����r��M�3����h,?��=���O1�e�w@	R�dC�V�1g\�N��!(��A J"�|>T�Sp��'��������v8��nEY>^�Ż�9�JE�������;� U/`��g�v�eYsk���.�(qbp�?�t�l��TAk�Յ��8���pi�ēB���v0,n�݊�<�y-�`�ݎ�]�d~�˦������7�b\W�t�vc�ؖ�r�8zRv�j3q�(�=2����GP��5�N���zk����#�4{pj8��t|���|���=ց�d�Bk��FW6d�
�"a��2���Ŗ�<��7��O��&�m=7'd����W�'Ȣ�^4ԴgI��֌��tj-ឯb���D�5����N�ϱ�N72�S�^��n���t�)�ֶLahp�l�����F"�^�F���"��9od��_ ����H�K��'k�~��0$R�Q̯᪐8]}�29(��=�˯�h�C���B!xH&�2OǍߠ7P�Z��]�rp-]Mߍ ��
{/��#�ZѼAg�W��ڨ�����͈���k����,�-Tx�����dD�TL營�n��k����|3�̀>���V���:^��Z�:N����5�i���$$����W��/��B�G�j&{�N	m�A�S%4z;�[���"�#&o��r�rgBa�Ǻ� 5����<�ԟdł°��SA�b��,p/���.A\ָ�v6k�P;���~ܿ��o��M��$�u��@���!��7�z�M0����
)�H��2��{T�s6/~��J�?fK�b�}��0몍� <�X)��_���`1�#��S8����>�rY\i=��t�ĬnF�v�r�Y]��� ^���B����П�0#v��L���?��1b����R2_��R�#��
���WM��ѽ�.G7t�j�ro����e�א�_�����nc��b�:�C�����?��q������{� 	��X]A��ҜD_�f�s��&�,�OpoY����'��-*	^��h�	S(�����=�� �l(���	'n��Jyt�h�{�هd��O�ྞ���0�/h�����o+�����3L�_��I�/��
����.!�MX]��G�u�i+M+B�1�y�~�k?�.�<=�\�Wh�ףv����Q�愞sC3��PƼ(",��P�/���E�] S'=AO������̭�͌���� R��B�֤y{CG���F�rlZ������AF����k��5a[b
����Eg�U[���R�Z|g�ǑOS��2D�Ǻ%�	��Nl|���A��í�.�k��_�a�A�J�6$ �Ѧ�R���)�����4�Ue�i�jڨ���#��F:t#����ϷIwiI(P-��ųw�|�ɎL��f�a9�`�T��=�x�1L݆�|��a%�~�	�e�\qV*9U�v`�g�|�"�F;)�,w�l/Aa���~�1ES����N*5����/)LK�
Ӟ�Z�3T,P~�W��i����.:� �m�u��քF�؋�"?����|��Oq��}z�w5n+ᴘ2��F��lT!��'ga��-�Kx~ϥ�&!�
�a�l�i@�e�uB���3+�����>B#t�Z]�r�3��z9�| ��o�� M����(P�㶋W �7~~^Dm'�tq��y���H�O9�m�C56��rD
s#�Tp�<���q�@������m��Fޠ��-$���	vb��_デ$Sn8SIZY���v3�J���xp0�x&�k�W��� �gt4�;�Y�[���q�*�I�|L�Q��!����<@iǖ�|�'=���,I?{����	}�� � ?��,%g�
�g *?��漋�<Ō�ym'Fr�� ��=��<=�����֪1GX�50�f�������I��4�s�!��Ē)�3���ݕ#�?��u����9�Uʮh�@�n�u�{�鞛��Q���0s��Ϳ��w����JO?�^����� -Z��i��"�<o�E��V�AnI3� X8���2��^��̸�qK��4}����29nwܙ�M�J��_E��"���������\�Enbs�8>P�7�k�~��p�����m�̪>\�kP�k�79�a�'����(�!
�a&0��s���b|�k
hZ�C<:j��LI�Bn�rھX����m�=�D�]�V^��2�}�z���	,� �_]�x��(��-4��Qft}�1�71�M��%���A�/���hsB�O\t�x�$���_���Fq������Q���l��q=d;S��L�Y�D��[��P9�O��>�Q��
2"�#���WZ�!�V��#��f2�\1�Ȍ��2�3?I^�t ���rPO1�8⼛)���|�79�<�r.�z�u+E�U�����)�ʁQ��<��	"+T�;�ݱ�c<֐���Z<6IbE 5-�Q�M1����8��ԩ2??�4��
x]�W��߭���d=
��{��T���30���e<Obt{��3��]NU�.�lD^Џ��J����m5=�z~�~틗��ަ�8��D�i���Y�Ҿ��M�{�djǤ#��Lpoe�	� �P�p�J$�nR� W���%P�ڝ��s�P�hU	'�R
t����c�R̬�ǭ�O]P*�	�d�ķ"�)��Q*���=��'[�ʩX���?F�)x�1t Cuv/R�f��P�Ϫi�E�j�B�v�fb9n$���_Z�&�R�|63�O�Y��1�!P8xʡ�\���Y��uc�)����F��VGR3l�:�	�{�����s��<r�uX`�*B�/������k���6���D�����>�B��Re�BdT�xP���\&<9bU'.`��i�C�[
��5<�y�R�_fn�eܸ�+� �}�31��<�Qo�{��,h�B=��"�j�ǅ2�!��ym���DB�����f'D�}I��M L��6ȗ�p��1'�n��[SU����0o���=G��� �{�KR��Z��rv4l��Ե��ן���Upf�$�����X1r��;k�LϹrU�:�r��T��(eSԲ�.�Z@:F����ݚu��^D$e ��w����X�$O�q'1���b�d�;Gl���둟�:��͜F��+�0�kݱ�P���'H��%�aI�l5���ݠ#Z�M�p�V���<,��.G�w�ȴ����M-���]�uӵ0~}����� ba�K���u�P<s�c?��a Yѽ��vչo��q4�S$O�v�G�B�Jķ�GY�f�$&v�ִ�)��&�Ì��B���8;j5+��<ᴀ��"�v�����W?8���X��d��V+��1�c�����X���HA0��ڢ��+#i��}'��D�s��GN����U�vm�P7(j�';�vt�`�#�T`���8�������/�J����ӯ{��W\�c�e��:,|Ѡ4&��RI;���FT"�j=��'�N���$����N` }�3VP��W��(Ŏ���T7мL��X�\sۦ�:;{H�
�X饤F�ᬼ
������3ݞWi��	oC`���KP��X{��%ӱZ��S�dI۟�ƫ�r���-��P��0�˃��g��cHO�|gB�p?�'���2��砭���}���/�bog8h߯�ĠxIMƐ�&`T�rk֡`�7���(U�\G��4ou=H���� ��
G��f����G	� ����49e���F�[���u�}F;^?�g�f�b)V�ƪ ޘ�W�8<7�J�A�I��8W������&� ��\����)|9E�L�=�Xy����Fl�(;�12"ɉ���O��9V�@��l,��Z�C9F�P����$Z�*y-Reӷ;���S�����/��8D\���}O��P	8��xepr�{Bz����/��!)Ym���_��L=���ȼ��,}�'$!W����!�	N��Z�����m�2���n4�ض��s-�������a�{~=|���P׌�zn'�i�W+3;�]i��$�^+����h�o�+.��@���Z��#���jS��̙! � �(H���u�Yw����p)��I�Z��/1c�)�@�ݢ��%D�Z�2$�����/!d����"����ndH�u��I�߯=�_nM���+��H�Z��aE=�D[0�c��L�9\�o��6\��]T�ʾ-`9PkM�N�β(T8�����KS�����y�k��y]adQ���S�K�D��X���La>n�u��3{�o��nٍ�nh ;��ƺHX��?$8oe3jm�<��q�R�Э�sXJ�������%L/'�7`���L���9u1
꽱��lf8-�p�x1]*G����K��'Cn-|w�ב���[���#{%]g�� Ԉ��[7�E9���f!��tR��ߙM>�rA�@gJαzL��,=�2nsڝ�!wq�G���ZQb�j;��F!w�{*�8�Z~wƟT=A+j�5]A�鴹�`�������K
\����j�l|�g��1K�e���í�#���/6B�*��Q����V�z��T��6J��IB���ÿ�sV2m�~D\��P�}P�h-%
�t��[|�d}����Rc[��BQdB5�3�f\�P#R@k�3�[�vsM݈3��S�dBm���J�S<i��'b�{#`B槇��z,�Ǝ�c�n�����O��)(h��>}[*�j���W��9O��������+G��d��AX��,�Kuf)<9���ԙ(R���s�+*���v���ɉ��JD�4>�܍�6�mY�o�������f��:G�;T{��n>�޽/#H�o����);�� �C�d���A9�Ͱ�\o�"2���6p�"p��~���@.����c�>X�T�wVhf�,�B�V�˙E��.���ʒ+����E"�����d%:�j�C��q�`�������1H��	sHO�e�nlyy�L=�6?p�+p�+�% �If#�1lT��r�hY*�n2۸��[�?f��Vw˒|1	~�k?z���\OP5�c��3�ຳq9��IF��а����O�#���$�˘�t�\�&W��Z��8&�hU��[?<Ƣ~?��7�NR|9�j�D�n�"�%�0�]m6��)\`��S�$Q�*�p�����p��^-�)M�[2�Pr&�o�xh�Yh���y(�os9�vG-�OߪN��M=~��yҥ���tZ0����:�3h:t}�=�#>X�UBI0Rq_���T���|O�Y���YZ���X��c͒F� �%=��U����.��=W��W�c��b4D�=��)=��iM���,o,��)b�j=�YXYw��R}��'T���(o$��fv��L��{6F��2���$c�y��55��M�p�\@�>=92�L�Dq��6ĎEZ}��7���C? ��R:��#*�������L�Ղ@s�k�̨f���!U�ԙ��7�)W(-�Xz�~;��ΦCXuR �>�[�#���:�fb������T�gfxi ��4H� ���������V�
4��u�.|�l���%d�bR�GB��;�!U�J��+�v0T�������Jk(��"r�'yǡ���F%v�4����롿�Fj�Ȯ���J]��X�)oB>�2LL�t>�Fz��;T��OIn��c���+Mշ�®q�Y)�׭���7v)���7�p���TI��J�{�S�_r����d�-w|\eA�C�J�"��%�xwm��/����D-L������FL`��0�=�����Hd�W=B6D|=q=d�sv�>�Ώll$��oةɴ����sE��G��]ͧ�{&0A�D�̒���&l�!~p(�S:�pnsO(S�C?P'�����3��π��Z�>5���ۣ�g�E����P�Tgג]��{v�ڂz���gچ�"L+N��ۣ./�Ɵ�B{��%V��\!/R�W��ur�;6�g�(�!���}̘�� ʿ�1%�.�B���`=yŦ[�\��y��bH]I��`�w��*��g���C��k0�
^�����iV]���||_��ڣ�!'bz��'S �gsP	���q���Ϝ��s���T���ȤK��h=~1�ApN��/籑!4�FloU(��2�>���O
������/(I.B#^\�d�K;����8��xdWe/�CE �OHZV�Y���H��2`%�akF�e��81���;