��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��!N;�?'ǝ�{9�1�\��,�L�B�8��V�R?��[6F+�+�4"p���n�d�#�$؍p�����.�{¯q��ěW�F^��A�S*��|��Ea)��sz�$��O�+�d(�W�n{�|��C�:� O��U荈PjZ�h�'#��}�Z7��-?D����͈#�26���1�o%3}V�9M5@�����s���F��	+�5�������S�/	��;;�~��g��JRyyҩ�M�'������Q����4�1_A�<�����E�s������?�I8��6U�3[����[we'C	�De��m�!L�����;ܜ0��V�~Ջ�r|��˛a�1X�=��
�M<3��(&�<�<���U�p�b��)��+1��+�����=�	�"Eβ�,�������pR�Ry�+f߮2j�۞o

�,>��������wX��2�:D�J ��� ��<���h�S[��h��-(��(�s0�9��5�[t��s�Lm�����S����f�fQ
���3��?�$7I��Vٚq*�T���8�!yxɕ"��f���&���4Y�v����^�re��F��������]���g��D���?��EH���2SM�>ZT�Ӷ����k��ֻ,��9p��3��XoS���,������vtD�S�Z0#���:0��8��Bk��{����7��e�ecQ�6~�|��/��8������y�dgO��4Y���S�`�_�� �8|C����6 �N�.���]�S=W�h��5_ @�WC8��#����d���.'4����'5���@FjL�D6)$2Ctc�,?������	5��f �))�\<~	�*o���>_v�N���ZU��9�`�ly��.l(]2ȴG�
vꑩ�/���E}n����'�ZG��b�U� ���-fɦH����eÁ����&�"w
0R<�{����-.H�b���r��.�6=�{���5�3�?,ۇ��;ր������$�6%j�r�D���|�ֿ�w�3蔀�b�pM�-1�3�vȨ~/��X=�H̹j��.�V��������}_�����4���ѿY6�_0
H����Q�9�֯uFE6>���P��9Ԭo�zD+���s��1��E50=�+�����sG�(��SB���?�a�o�C���q��W��
8.����G���͆lb�٩��2������Q��Y�ߑ�O��f3��Vr�y�?�����N�����wEi�S�ɍ�'��|b�I@��2��CA��e7����ePtx"�����_�CBC�3����4��`�"FWi4��~�u*;��s����!��%a~.տ���Z��G�z�O���Ȕ���q97�G����Ӟ���!zz�?X������j�(����SOݕ̎���i���pP�1ђ���=�X�:F^풵e���1�_���������.��h��~Z4��d���h�o�d�̭y�?��S:O�����'�!8.�F�R�7�aiY��M�ͼ�Ům}����&x�(x��u��b�;��p���)�����:{Be�{H�@��S�3��5�ǲ5QS��`ܺ��K�W
$�1N��م�G�"�I#̰��P���Q�ݶ�*���Ug�ѯ����vJz�XA*�����0 `��w'��Z'!`K��-�!�����T[� ckE�	����F��	h.��&a!¶��ݧ����;Yz��'{�0['N��T�Vi��ͬ.�BDy\Kɪ��u������+�b��<�L�0�|rMu:����td����;�	�I���̫-}WI��y��X�,��[�Y%�"��g���P�>=	�8�8A�by5�q;?�o_4F���|d>(e�c{�M��Ec
k�x�� o�W$����V8��,S-���y	���EX��ɪ�/%�tV'�Ϸ�b��b^Y���p���BBW�oTF�/m�!�k�Z0gD|��J��6y?�P���9;������7������Y��[�گ-�Q��K3����n!G��^����y͛�q��s���DF3A��}�@I�z}�`p��q9Ca7�r0b��gh^n�]o,V6��7�mi��}L�[f�i�ip�	��0{Q�b�Fy:)j��/�B�Y9j&ƚ׆0 g!�`vP�kNk�Ž�sa{;t��}��{;��ޖ��w�d���;� p}����b˧g���S��1�/��Fxzi�?�s�9�B�����(6m�qk�"I���ҍ�|>ߏz/���N��~:�5Q�샽d�ϸ��S���H�����4���%��b�y>vRm��}�f��S��0�O�s�����c�� )Ԁu�i�?�	�PS6�r/I"
#���mc&:î�l&�2w�c�����X8J���Pb�@�Z��b[��m}ɿ���{0�Fڄ���6Ǟ������Z�G��uy6:�_�?��G��=��S��Ë�8���}:7�L$a��f	��a�J�c�_�9�T��r|M�	Ԗ�k�B����I8�s"�*�nl[���Qj-ٹ
%�����4��QL'U��'|���$Wm�O��<�ż�`�0	��2�y�6�u8T��ҝu���mX���Q�x�ߞy�o�[�����YYwy�?H{�����sR�a�s�/�6�s��c����L׵�O�R�����(�����@��zH'x�\��_�S�(8r	�}D�:�Z���%hߢ�!�f��p�a5L-�#Ȫz��G����P�t�|j:��9L݃Sz�l�>=H+.��<ND�o���=���N�i���:N�f'�1�>`�G�#u��lۊhj��of��u��h�Sg����-�\�`��j��UY�ވ���
!���P������Uv 
��� 4�W�+���KvI���У��