��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�`��L�o.�/?�߈��Ubԃ�]"z{�y>JԴ�`�rJ���m�����E�&"čz��<�u)X�V9�p�T�/�nE��~���s��w�����0|�_����#�#a����du.C��)C�ycR�����t���0
7��"c�������ډ
�&pQQ25���n�]�@y�Ņ͛a��lP�_BNnD�S�����;S���7�~�7����_?wPv~�8���,�Y=+}�Z<e�����r�
~��iB��8ˈ�����շ��I��+a�{kPN[ ��J��6O8�hq˛K&@l�J�VW�ĨsC�ƃuA�[�N>Q�i|A�>5]��l
���\���^&3�J��ד������ݔOm櫴���t����=^1��a�M0�#�hT�$=�{z�L/+�e54�F���9�3-�<�u>ԫ�(�w�`N;/���{�/-�N�s�z�#��`�!����6l'���U��� E��v�����gV��y�Ms��*����R5�m��yr`РaH�rߌO��|io��$9�5"�c���ך���!����_vf߫�A� .@��[��� G��z��\Fu��s�Y3��a��	@AlX�ᚯ=�yR M�nU�e�d����3���l�hٷ,q�
�eJ�آV��s��`�Tg(����0�f�c'3���>lu��nl)K �A�#����g���k"�u��5H��j�&τ`�u����W|𩭘�����e8��t��99bU�=M%ʨ�l8��/��eNz�iv�Y^���[c�X �}������C��@%VI�(�_�Y2��1�(\��]�R�|ީ�Rk�����q�	sY�E ��x��g*�;��F~�mof�mȥ0]P���N� ��_��0�k{h@�M�^ ��F��!E��L�)�W�������4�agf(EuQz_2L8��i��WW]��@�Uz��O�I(��4�k����ۅvc���	m'�A�0T%����.�"��"���TI'_G���-pe�A6wm�H3-�r�g�ȍn�m��I��!�x>Vp��-���º��B'l����*�
��t�^6��ՠՇU��e�h���K���:$f�fm,ؾ��P(l%`
&�r0�����7�xƂ���Y!�����������c�ෂ碂�q#J;:�cW��Օ3qDQ�/�O�ی?4��	I:7x���3&bR�s�W��H��"�����@K����^1�F����i��E1A�\�P�֔i,��v�s
9�n�i�&㱲���Gn�����`�W� S�sw��g�H�����ڸ�|%�̷��V:U�W��{&=ʚ�@2l��O%���֧��Iթ	���^e�����KԢ|x�V�r��@�F1a�u��fJ�y*q�h�嗿�F�(*J��oׄ��_����'�rOrZm�^KxʦB��k�o��A����8��+ar��>���w�T���
��J"�]�#7"���Sc�N��U
�묺���#œx��~1��2�R�=�;����S�W��:z���� y(�:����*��R��%m,���/U�s ���3*|`p����{�N���Z�8�3>)v@)H�;�o��v�q֬�1���(�J��$Gzj֣X�)k�cY�V(3����h<Ҙ%䃁e�g��K���a���I�>1�4��z����;����'�(���C�N����1)%��B�Q��yx�C��k7�a��T�q��G�i�Fi_��o����#�?�
M�4��x�ե�C`��)g���ރzV����jHe�;�O-J�J�`GK\S��Z�P{��Ζ�a��C�Q�)�#�[��x�~�+L0�F������e��^DQ[��=�����O�^+_����$���>�o�Z֊E:Y�W���4\�W2�g=�2(�>T@��+���`ub�J����n��Y�2�X�2$��d�_w�\@)�Y}������-�����#$���a� �|wA歵�/���-o/��\T�@!�a���d!� ��^	 I�&4�ċ�����
r�[�j�
du��i�^�����#Л��҈�����2C�����h��=ޯ�jo� Ru$L�B������T#��\[�����f;�A#W�<9fQr��|���ǭ��v���<�Q� �
RS
��%�Tz��z�<l]������5�?E]]�}�"���6jFA�o���OR�Z  T[E:������/�"�y<���Ԭ>a/s���s��1��_�"�k$"����,]rE&L�+\B/����sy���uR]�/�
6.�/�# ��\�̾�邵i9��g�H�Oq�7L_����������Ak�5T\�4:<B�����v4��ϑ�2-�ϞmA�	FC .܄�$	_
^�j��GXK
"Ug�Kq�_=��:���ꟅBI^myn�5;q��B�����E��o$W4|��N�I��1D-/4��z .�wA��Db{�nݜ�}��\޻e;�P�`V�	�2�-�懽e����|�L���ڡ�3b���^���'_x�o[9Y3�y���K
I�$@��b���!�Z@��V�yIR
���ظ�>W���dh��F~��[�~~i`��'�R��� ��0a�Ej��2	︜a,�S~���\k��ė�y�䑝�$��m�����x��� �"��H��6�)sɇ��qwg�Ũc�����P�Q�r90j�Q�'�?��ƌt�7>x1�#���>�I,�	���\Ǉr��˞
."�(�9��x��$�����O2F�Ny�|G9N�x�Ll���B�r'%Q�V����房	m��ݺ���U-(+X�/F��?�LY�,`���  Z����Ѹ�E�dL�����ۗ�"�I��.?x�7���kNS�N��'T���d���`"5��\Nj�v{G��y����ҍ�~��m�o��"zN�{����1d&����T�?�ŻV��9x��!��DrS�*f�:L����a���Sd�w�+w�e�/��Ў��q�c�a�ĔԻ3��.�д׾G<1Sɡ�\�K�r�D.�^{�ը4z������gѣS1����]˗�̣�x*�O�:�����j�Ш's��̣>~���<��������5���Ta���P��eY������l�)ͮZ��<N1[`����$��9�0�Z�܉^(�ծ"�	iM����f_A�)yni�N��z����n1$���59ʼc�V��$��v���n�s��O�)��',�M�j	�z6Yc ���sr��mc���[.�����m����g�%���^�m!ҡL��X�