// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:20 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d84P+xuZUOlLcCzMsKOFu7ZSOk72rblvqOojIX/BwRvLi3SwpRaTA4CIPhv+nh5l
4ar6NZwJic1l3WFDHse+crV3CoOiiQDeeCROOO8uC3kjx9GxbhFHmuc7x2zLuUgM
FlzLb0X/lnBsFF9yBC7RPZaaUh/KuGrFCLlfmgyLPYI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 93152)
jZO9TauPFl6SZZmVRnq6+dQz/trReFf0MldotIHubGK3sVGIwDFF0dHItpuwOIpm
RwM7yfI/xJssbwbIyR+IiBo3q+aB115eKqtpSaJ+1Upksf3GVkjgKYWkOt9ZGsUP
tUdWvPGPS60w1yE/V6PrRXXhcKQSGZGegZEyQby3brh/baAxXPldDduFcdJGrUk+
G89AHiulsNQJrls59P/s3sx/YTyIeel5w0Uj5m6k0UyjQKyQbZ4BTGsyQp2DYqhy
zJftck2ymUlLqOoZ2ASN2dL7iWuF33eIN4JX65+X6te++x8jbVbHuLHB/ISpztvR
jIAVssWRO7AX3JHOUVIcNppI4JsvI9X6gOMOSnJUBsuCqzWCNSMhFPS4xl5GRNcG
Mf1Y2McH5qDcSmuIcXJ30Tlzl+4qaZliBFQIDle0uUHgQ8fNNLYgamXNeZII6lgb
s+gTg37jmRvfswaBTxxuQJQrwmMll3JcOOsPmtYVwuxS4bQDyCPn1k/XasUp2V3q
7gJTDzT3kWAd7RPQkZgCymWjjSi0AwWlBjlynGkFZMCqRznQajNwMf1oQ2jBrRgr
eMoZBSEmuV8hL1I/7uRem3jE4OA9/kAp9y7OA/+MkGtiv+8tMGrl4TZcBHVSXUQY
Ey9W0Qk/nUppG0eZ+IBLhm+a3f8Hq83qhQAuNAxbYq4JhS3qOQDEqeXby1NPZ9C+
g64qjiXUobejK1iZeG7izEgVUFaypifJUVvEmIBqSSPts6DHyKRYwTK24h2Ms8oa
1s4I2IQqkR0IOTbr19d9KkT8VzzZW3WbH52JpFvPzUg3s7hk0cOLyCumV6gOrtg1
xrr7+UhLr/bMxa5UWkyOVtVS73dCpOn+iC5ZFNTz1eVLb59rS0WsIICr0bpWR4Cd
9xQmRx6j263Gnch5IutvzHuM87CasnklZainQIR0vf4v4eUbzX8G6CDFL4Q26YQn
UVgWeJyTIje7nE9tmHWnwBAWXTMqWGoP4vPaVx9gTfU1AHVTymkDaW30n73aiqbX
f+sb861fZ4KX+TpspoZDSUQ/K4qTwZaeeb8KTMexJ6iOJXlNIYFKndfcyWcM+S7N
1wNQkMBxzmC4s68fxY8PRx5ZTkfbtvhrVqvUgp9zmNUCKtHCWb68b2cIdBoTVAiS
lRyAf+wWTMuR0QL5Z7AwzmDB/nkKFw7Myihx/dq8wbkDBBJ2BmdujX9VHuGbY0g3
q+f5ZmEKlzIuAkrFMT1f1WfQY20jy1pmEBuYDW40KhYG7WQAyOE5oaXHMrXidVP4
9QPwcboa9b4G7yOqmEu5CAPuYA7XOca6I/xcoTRQlTE6L453ftrqayPWKW8p+dDH
Id8HOaDTHZsl0q9DUuuszrQfRKeQ8l+vEzDyE1yd8o1nmAnSqG7XYA++AY3mak68
FYETu6Myz2ptQMBVcsXRN+Hl6JkBEyjvkBXDppgijyhSUGcPH5LWvatKXPWYArCX
TZeZwjU9DSERx4a8S5BjfnofP4NylIks8iJuqYEqxYmqkAPEwmhdO1nP8mkvCndl
px2avLltn2Ve3h3EHuHaY/dnA4/30xBWVb9JkbcvaD8dR7PzXuc4tJxWvqrzfkUH
ZQlfcOZEkfmkge1/47ihqLCMaUhnMzOGrH/LSYiwRqvho3UiKbj4MvmdQHwhZwrW
L2J8NKLVtwsxUrswnzKMDveaM3vXcQKdj/dQTmDL0UqviNzIEGIZr1pw3O93M0OF
ETCTJUHR9+br8Y+MD9W59CAhbzjhTF7QwQoWU64zt6/T2apFmQz1PaHZBXpKVdc+
YUfcEBkiW5aHNy4/ksfMcLavw+7KEIjM2Y5Me3LzPdJvmkfExhK8QfA3bKATWbs6
DON2scbA4Kab/+9PPPcUtCVU2wTZdNG5BK06axLKSktfJs/CrX6pBKhYOiruMcu+
wgaJX3Y8/BNUObo8ogkaU5YrUjPHuU1v35WJPgMPNOhcOAqYSyQtNQZ2ipeq70Z5
vhmCUnIuKW8yeSz1mOyDGon1m9rjp4hKOdmP5ldFyrvtsNfLZu/6YG8SesI5YMvv
7jT6MrW0NG7RLWEiZBQBxkDfcVSWOeQcqNE85T27MDJqm0kThwNFKHFdsp0avyP6
UID8HejuQKg5F8oy4VDuvqNPCr+VLI1GguiaCoM5cXiWdK3+NYgFNud3VgSts8/m
HyM6wB58PHfSrb1gEzy8CYGipFCRUc6/o0MATfph4TSoqdSufFmyUjlVPzD+llXD
sMe8/u/+KnLM4oH74DUM2JzJwq556IDHUkt3MRHJUO0FlB2S3J8iHdqftqsbpNEJ
BeUFqZZa5rRQSgHZGVUjlr7SOL6bhNi4esv/cg11OrHNCx774ZTJpbkgeSizC3SI
8cKgpdXLUuohQwjxAjEIXXTJgGhP1ecx+t3e/00qaHnrEc7bE2EF8nHiACLbAxZE
+6yEdWLTFO2ZuO9M3MhOq6ZVYIbuUgARIc899jqIekbZV10oU9VMrusUj5T8gVY4
60FHHvadYgT01QxFu/hVCCfu4vNrBuvcojL4qdeTIOzC46S8587c1RGuCoDXPpEk
eGnfAak0TovTxw+o30ureTnklxnbkESCQb6WMSoRFg46QSdDTyMqX109Jqd1b2Lq
AxC0INb0SoHXmdjKUM4Bgki/3bZC9kDF4Lwey9uE9dEA6f0/93YeIq4rTkeZDSU9
cgC+PwbCHTZnXYMfQXXITpb08Thf94grni82OI5wlTkp/+DAux35Z8/K/w5ezErP
4a1Bkm5HegdcjhhaXlZ9uuUqFRQJ3QwePIQrFED43KnfE6nQo4wGcRvqVwqlnFAa
vm8VIHmwJOlt1DHLIZ59tTMs8L4f49mt4pO8dnOTRfYjjjDdyaUvT1FAU4wevG7C
7uvTURus1q0vkWEX/M84T8ETxkSoXLkIEYUORNXTCGD+f07T5zy0IUWiPF8X8Cyq
SQLGSR4kakB/eF68YXUhoHnV8QJOSQNh099aunfzxqcpJOnTqfFUnjrQKbQWSaIz
YZ8SI9oryn8LZabS74B9uZ5lTRnz/eOfECb/Llgk+I4a01k8Tv4frTqZKjTCVVE9
1US75oaAy2HsamuoJb0+hcFFjxuMmbEEfKaaMTpm2OZsoDKu3oVZQ1YFRxePLepJ
bYTAAtkqyUqyyMJgrxX4feh0Yu7j7ogC5AFGwnwMgd2iCfEIFmOAYcEp5l74vFWq
Ydx/4owqrrLa176Q5GZ4OA1a0C0oU+LU+g2V9crwpM+sWthkIdR4z7rqelDOWVsA
Wstf0OQILk4mUI5nUlkFZgV++O1NHQJ1Q/gS1b2gk2lCOQEMbTumXd2PPIVSTeve
C9qXRvUwuNAqpnvfhjAJcKbq2tl4b1Q4Y5Q4ignmgUZXegLgyiqI9ynyaWQjNcQI
D0R3fkOfsw1XGkBhdB66wtXBJdTySLDLhVZcmGV1ERC//uiKm4acZE+M9+A5Uclg
jD0RRdiZSL/4W6i1Z92Ui3C1M/Fox0NKkoGP3eGfFAkcoWCf3jjjc5NrP9B2py8N
Zk7gaqzPR9hWLIyxfzW1eZjQrT2Nu2tblnkMAIfrSH3gw6b03h/2ku72kEk+84B4
8OZBEFlHX8tozQCRZjEZdPTA2IfC+z+FqFZed93vIvKeKVdGWlmC1A5+BGA676pZ
oWEV+AUEyYwvYSaO1EUAFWqvqXCZQs5mE1GM/4cDKp548ccyqi/8zTl0CmyKgUg7
easoaIKf8xdbQbfL/ZHgdVz5yJKXjexNfPFE54XjhwMDCLkcVtokHg0Eds5jdPNf
rOIa1Xn5ApLYMlSkeSGZjFuh69MuPG3w3NO20wRmQ3Mg2T83S+1qTZV43rRZqPAt
zzRCNCR5yiVpgyCiG2/pbnl4OXH8p9di+eFKVM0Pyt+vKXg8i/nWn2im3dVI2JDW
WmEqblCOCGKtxMTsTPaWmPDgu56TcpLB3E3aABgOPOitlhQg9uKMNhxXqdrzfsN1
bGmqkAgbvQwE5uYEwGb9ruhcHitnyEyAyKro0YaFCJ3JZktjx5O7edtWyH8EWLxN
OW7UKfkqt+rsgQPHiC/vYHRWmuu6qbv7l6PmYx7UaydKgbGVO2FEUSfqHs3lzq9M
dvzuJGrN+tsR/Ezo0G6JEEaIwP9cEa1ufCeyJXtDlljMvmY40yD7E10BXDpctnyT
SHQDOpe7tHSGFS6xcUIUYogH5M0UBxyZOnFAimosOfZlJoHly3cOy1exnwkq72Io
7bGqMDPU1cCzghexdMdA1qkg27b8TyDeUYfX2gAPTzphveoVZJBRXSGeUn82ECDk
cdu47VFIc4Dfduui5Qhehqyf/Fk4bUOL+oVeLnGOpt/AfbhxcYdBGGlo2gi7Uldg
qAZZVvJBctWThpBF4mAkjW9W39qYDk1XY6rn1VCw+hATRIb8n/yCe830qBf6T/j6
5krV+q+Nvd4Li6vvaTW4AtPKHtdDalq5kGKoLI3xIYbHni/UO1kVHvrgJhHTylG8
kLsPwyMIhOh4+rcLX5GKujNBrOrsPEIlQbiJnPRKFr/nZs9XxsplDd+/ZXpgfue0
JejB8XugkkoGfNrXDp1GkhxOsfZoH4bRUxksUoId69IMIYbrcG3YxzZOGCnsBm1k
YPahxrcggYlnCNZ9uzZ8YKXgHDESbCCBKRdwtAuHL38RZ+6u9lEFwu3yAwmVLi3N
OCJZoWVHFnxsOumDEwz9uxQ+2E09+mIEDIJmpi7uo07SvZHo1TtAVs7B4ufj2qNn
0XI3T2MPDzx8B2fpFCiSCzo9hkqWdApEaFrZILPf0r1Bw/SaIAgbdASBtHNQB9tQ
JAQqYd85VlldzYwrnMjyTDgRwik0sjp1mwZvyhaa/zzUYPT/PdbYBX2ljk/0z65Q
jFcyhnFcr3lTWL1dOb9Co0A4sOseS+eoeKe9vt/A1bh5dKhXGtkTSpKM629a9N0U
0ACXwu4oMEIbZp4fT+uQmjt7YffmpeGqTTaNMd8U7MqZA2bir4ZmiypaOvrlZbKw
+bedhweQuTPfaZUAXci+PwfkkIru1MOMvWSc23NRPofU1Q26+rsGONumrtJg8Gx3
gLK3lhm7oY1CJdmrYOVpuhofggnfzlVuoltbqVRY0xbsRL3WkjgAEdsoojwEZUFK
jwdJ/BTuWB2zllI3+4fqp3zFQk+1UP7Gym1qF3UKXW5NmiDu5TljnaAH7DoKnY/F
rmMe+FfBlDYGzIf25tgP7z1rx2WKQAvUP8aiVTaOy024u86QEkSteoC5xLScy8Ar
YB1fVBqvS2zk/RgeF+QOty9Vt1AHJnNy4EYbgkwpOOIVX7aB4MzEdHPzud7AQUe+
Bh1ean36Fkxj4o2Mi73VdC+8tkeoMd5qOahhGQChTl7nA2H7JThcHgs7BnYTlPQI
J9uFhP2RR9rxPMsrIzBGqmMFYG/RvET8bfpXFijll5cSlW8BfZgUnz0SxCF6NlFb
gtKC3JjrIWzEEpjTDkX8qE3y7HRfx+Wq6+Y252zaGRkDH4tW5XKdmIfPxWFWNvBL
xxeMc5q6ukIi6Eab3aREp4Vc2pstSVXrYcvTaRn6+WDSWj1zGqNEPVGsboSjo7zb
Ze7zXzZ4FI8jFcTKcEor3nFxtJ52O1wL1M/qQyGzC20eGegTKaAtl89f/a69zxrn
MAgqt2k7Em/b8UPAoJqYLEEDeM9wBWu6BwFgOG4uwGiSzGO7ToxOmO05aQEnfbIN
jJx9VrNTvV86BwoknqZNTpBkmOC6yQeG5WMUEW0fivubtvPFgrjb0qtrK3Px/OWR
J19I+0jUhBfbWyTzVmbY3F2ZZxxHifrWqSvjowZRpZPinNjoNUpbaYY/iCiMDRS8
FuUj3EA+EzuzuSTb4LkT+teEGscvZuxAb73b0X0gU2pXxJ2Uns1Xec2Oa2bWtrgj
20bJmpjElPFooO+cGy+mWwcEx2T48ZQDJFEr68lHU/Y2akzMmDDkX9682zM4EuBK
JVZ2U8mgDGSF7KZZu6RRGd+vwQA2eueeLZBRrbtGo9eanduSvyJgWTVO8Atprm5U
1EiqK6Uc4+ATKXsz7yketzAaxkSzOk/M46uw7jbpQZYtnWN1dXiOteu9gwAjAVwk
1JfS0uI57KKpPZRVGxOzfD3ZVWqxyex04fnWhzknO1JNyHYrfWuDwvLRR5bXpXUn
hwWTUCdJpVUItoU1hhSe4Cwp2tQ503NZzwTmZmsjd6lVDKSZN38osebLDwE7WUyK
5FZ/jSLfciZDuF71v5k8r0oXclGL0SXIxPa/lW6jEqXP30aqlpzL4GTxKtYeRDpw
hAjzcEDzxznctDYJwt/3El38rSzCtrHTuD8vdKm0n5rrLRE/Eujo1BhNoDLye0y5
rn73G+7+Xz/Dw6ErZEmUUSHIWAH/yJckWy9tPspQlo3d3WU6wi5MvMpeGZyj/B/s
/hYbH6PLYTeiQrV7dE9E4C/zda2fcF8kH4yeATWmJmKQoz4Mlq6sewG9BvckiyVv
XRZQ5+s9kujeadeirRUJv5K1S55z6gdihGRtwXMtiPsFtAoGNJALU7uZWPPE7Iqe
busZttox9maPq/6ApsjaxsVhq/CrVdi5AdVNfrkA44GhtwV1s2bQLuGky64KThKA
fzzk668dmdf3slNYPM7ipf3yeFCTeSGI3eFhQ5Wz/QQrJr/m1TkCUHXJYhN1ZUGe
aFcGTxNsZCRaZONNwu4TQIvwYtzMJlVLVWoF6LZShELaV0pzE29prlX/DVrCdkKb
Bti2bIgGEzr+zdDqtvxKfPkMPjQ+ZYnbjlYA3VTBQZAEeS2L0oAxbbxb85qGylJE
E+PcdJZzbpsFsGzPo11yk5olGnVwpt/qcPd5EX+eWHfKCiX2ckHgb+3SfXvDYKWf
iD+dPy1QNTGOUWcyNTWFlJNvDOguD3oIbkpU3WHF/XxShA0MyIHgCXBedy/WjHrv
+MnxhIy0Ej1dcU07RqwB3zNByl9D4dODdFAT76UdJh4ajgWlQyEfmeMxJd1nOKRv
NlaIsuT4131Aqvysv2CMo1GCUD2Uh3xDmGMOOhoJHa3yQXzOGVISJXbV7XvN+Lym
5mG8Yh0/MxlSlRvYperh/kScDH7hkm/sHMSn0Z4xba/jNqpmOV6aXMza5+7oaEJt
BKAsezfO6eBEUtsHo3ouohTB/cylUckOGic34XTOEHFAnXXn3EryHrDDMC3NXk8f
dA8vEoBPD7xtDEOBmP2Zh6/vRgVXsmtWdHoATrK6rWWD1DbU6KpimQwlOiyFCR2z
O1zPfKKeoe46bKS0Z7BFqaP/CgY87eLD3EN/FhMry/Ufez7d0IYotlNgHxtxuEW3
at+Ev8Aqsp2jDWxE5EDtz9bVq0RN0+XFlZskfhauRx1K0qegwvXScuLcGAbs36+q
xzhNEW6uadkJYlrywkVL4nHkiTFoU+aFAXFU/tRk+vTdj1MB1P8SGSeMkt2wiCud
wg8YJxN/vBfRAV8Wzyul+d4VuRdgbNJnHfUogU1YUJD8DzT8uFtN6u8vwkMpGCKr
U6YmuOZ9dVwcfRXBMDQE06IY2Qg1U9IJ3hCfLbf7pb6lpHQw5SeN1qIE5w6FLWj/
vKv7PkzcDwbpvwHMECB79lVPS8mBGYhtvLsr3Kok27GzgdPZUCBQCkxIjJuSD90L
9NSye73bj3AiaWfulaFjFfbxlGFih3bvkW1ne4fHWe0ssFSDecxxx214rWu/D+Jq
3I1ADpbnjvJWEpY5BPQf1QLkDN2GaxSah+extvbGH5nPi/S6ZzlM/yOWL5KjYWLs
np3WuQKscrPA2iF+kYeYvpUdkp0B/ZyVZq+ibJavYMD2CW16GABUkwm/qBnsSkJ3
Dhd4IDqo9KNMDYl3RVJJpH4ep6iuka7v8UEyUaKaJKOhff5V5t4rcbh64K+3F2HV
irmk/HJZJmsGHl1mYckuSNfqmePNg34tLa5irrk9k0zgu5CE3uhDVhv5IN/jai7m
dN9wk+pT+NZmLgLLpXMoV7LpxVL5RIww/VwrlUMfVzDLs57uHqtxNcvOlheAw7tN
w12+scKO81aDUhl7oEX4a5R1/TyoqcIpU+OPaZuyN6L0d+3sh1MgYqIhnrQhUUY7
WwnGuPm08Mgqy74w/Wy9QAhsnPvp41dIbRY4HK8zpVMRDnQvqu68q3n+AQ4Tb3kk
xd/zugJYcFhs2d03hYlaEIZYrrkebELvmfmhqYkAI71gPwjF3HhmPC1djmszdGgS
HV3yChozZNFU65PSYYp5gcRVGlU4ygdM93g+/82233QMGCFiX/O5r2rnU+stsSKZ
jeGGzK8pFySvcfRd7GHPpku5zvs+i0OT4sTTtP+N+IYolPpYTPdXKwo+NZ76smds
9N402pYe4/i4BfQAPM8EICggkMJNiQz6cnYzFICUf/2MpqmTyoUyGUDzvWvqy2oP
d9Zt6LxCdVAoDrhP9e+yZIDRevsnfbKdB/RXu/jbWrdUDJ8TnGFy5LAuUPGvFxjC
63L7YHbfYWFxujYsSPzbqA2jm6iybnbD1hGnDHScRHHp8IQhxpPWT5vnnZrDsuRv
DLii2dOtTjuXYDw9pd1r2NtwxMgO1IaWqm0Pq5ug3PA0NOV7nHr0HLA+KuJkrclE
4EQfy7mhvzwdt5OfO7ikZllEW5R+7Nimi11yleD++zWQOaf50mqoWE2kGfXkFQDz
2ydHRCYOo1lsu/VuN/L8SB4erfSvPVM3/B/3EVZsN6d3CZOkQl8Two2iC89+WCh+
kYVEbXHYOpWCnbL0sU0JAvB2FlodGiZGvKZVBei2Tj72hy3XLq6vUQJZL89yANXL
d8tLknN68BT2Oza5DjPl/AorB7WN5B4fktCVcB3ReC1en2chedi4Ckd4i6cf9Tzr
nwgYCS/fCUqpanmPT7O+envT+oMH7FQTL6tU4ePquDavdMhNlY+5nKti+v5kot2t
a4CjTNuX543+ZtyNBhsDtd1j8VfmngZZQGNU10hEgmVqcdGQrmbDn62de1wefQqx
iwQYYbogm8GxtPINqEU+07Fs/wYu13w1MhYUW2vmwsjaGW6jGNIg5yxY+avmD0uC
j0PwiuSs0sP95JKODWf9gCmjdErwKka3hPhGqPmhe0XQheGaTgX2Os4ENkBjf0qd
RHOZuDSS0cGzempt9IWiqqdnCd3A3RGOCfCr1O1HHxrt/e+CPRUAfiycU1mYPUDo
+RO/Kq2QhvxSr+3yvOqxt3f/Lq2sI9iDlDrV6dkQ1ZCKdgCAETNVjytQ40u3Fc8Z
d+Cijz9S6imSqgNnKvhIUrkGtK5dIoj3PVIX9muq7fuctL8CRP8OEH9LjnRdG3Pn
NxodqioofNIcrKsTBWgvSU0EHsv4vrO30MpJkXt5xqyZeVlwhMf5ftdqneA+FHFc
3sVvV0b2mJR8JmA8nM4J4B6NlDXJBqSm0gnU5L9bjQ7+e4OUeflH/dBnznB6FrGX
uzseErK0Ovus6cG1C4P0u21jTuEXYUiwT7cMckGheozMur8jKOWt1scOCQHP/Osb
iaQCdpNW8GZrysOMNpImNPJI1NSQfZ4zcCfRhasAzz37LczDZzIU9eusP470gQMk
OPncRHFk8nkCMnGmC+gJfzZiv2svl60BUQ75/4/G2IvnkLOBgHUKxjEE6zA7JgKJ
Y59EJ5cI55qBBa4sIQ+A/BEdgqz59rl7+/a2GEmP2LzJvgbim40BB7E1lupI2CM4
2FYpjNUQq74MonKNwFrpo3vmqPGEhFPb5cnfeTgwePYijHw+EK8btZ/3PlDxsmJW
/tGCtWZgI0acUP3y5rK1/yrSp/MFWjYs1Rm/UwVIWgmT4ocdpvD7gITe8z9KBjsx
fO7rLpBVQTNJQZhXEZGwIF4lNaS65WWzPtjFlb6y9A/30XF6dGYPPdlHEHjLDc3f
x2RLHfO2LZx36nfwJljdAc+mOkTKL3WQu1zJIxtxqgr8gLfGHiWYmyk3u+qQJe5H
oBsVWpzhbbBzVXCcVdMnykhrpXnXqaEQOhNoIrVybr46mUFS48KdhbPnAtFuEY0r
m9h9lj4B52tInYsTnxOYtwBy8BMOJjTZpFnXUWWiomeUAzleMaMixWUsNKTJpVbJ
mdRVrMOk5O9zaiAjw/AY0/0MFqpSgLtVdUhWU0cjyHTUXQbU6tkqwFG8brczbxBY
+oqaGTqqv1RSort5hPG8jPYF12dGhS8MVwxjEwR0+CXJSqaARaBseQBpe3L8SWn6
Tsrr8rwCX5pEJTriPc7uM6CcvimMasnHPhOiVJ6CHtbnjil1vBIDmHFhh2YIIGtp
+/tn6KTyDajSwenL2bEHlUKN8IQRHabifLDkDXEqmB+7qvq9hODgT5hxwC+xxAtu
CIkFZVXCAWDQKOwv3pfoCoR4GIMbjo+ANMn3ahXw2A8elvMIz8MvyZy1OI0MzgiX
G/g4lBpzkK3cOSZQ5V7JC8d8JH9+5RIoX+EmBe6qcaHdU/+YGDgmbGPf/77MzN90
2NHy16PedSrznckdfQ3x2EYZMnf63PJKUDZrc5Qkh+jshGhcglA5n8RdOf9D2PSp
IQOUmd24tKFs9SCL7BPOQfV4nyqYvkO8PwB6ghsm2T1zOam/aFl1wE4EKVJgylSi
EUKBq9F7vmqnew3/6KuNLs/MgHNW25MmxdkMqKf0WKGaM1D4ogcSUEjpi/bpaqcH
V1WEm30fu/1isU2I88uCmoy+nomjfnlyK41YwTmn/8ulSp9qSrp9efoA9j+v0Aa8
o5YtZ2/35ABk5335tZZjFucJBHgF+ESRXlUh1xeyJepvcRnUdJCsmtQnAh14oy7y
6z4uI5iH5N6bVzLiD/ZXy6eO+3bsltxzzV/WcQXYmsnQ94ZkJA+I6vEePfLvHvsE
73Qhl0Ym3Dgjl949WcXquC06X9L9wGYhkfVkLG7vbBTmvVCZThgRu/sw3H3Gsmi2
YfhLNPdQClWxqYkpTyPpUZ3zWoK4rNsDnzuYm8ObxdhDBejSS32+L6SH5waFCLjq
jeMP4Bl3UpQQSkbQLjbAgbHxA6alQx2rzSBrLoInH7TrmHeo44heFpXhaMJGA/TS
JTl21vMtJ21is1qsD4IUP/YOYPZZvhneqvAfqiIwiiN4XiWSvgS5dy+LKY5TYi91
9Bfmk9SE1+GzEufzN6Vww0lzECyY2UhIohFBptzXGRrQZr9dCvYcNli4mzeLIX+2
OyqZpXQzgBFRhIb2e826a6jDS1lmRKpuFWEib1MywRSgmnmlUdTPAtxdUnHxwX17
8siE4uySOxBedjfCeaQaDzdNpX18IfwSrccsWLYCKlAj79wu54d/1Zdp2+iJ8SU2
uaKXr1hYf8bz3l2mlH9/hWp+bcVqyMRdiBiLex8ots4N0YftqkB0rLODnWen5A0p
Ok9GzqlRoaSAVnuFO6btYkGGfVo9cMf6F2VCfpNJaJYSFlcgy3pr8I3AjKyVjIp8
wNb5xgMxEvRQLXsXFKuaLK4EwwwFyarYSxBs+d0zmhowp5HWf9DrrFYm7pR65t4M
vjYPRSpyc6M6t7fjlE8WUSKwWex4PS6jMtodtSvV6nathPCYTKxg2D3YzguJwy31
kZLw+8A0udr0Htw4Z7LyUH+Uf99p4+v8qI6tKzPJKje3JxYmBIce+NWarc6x5mQf
vho9rPXFOpVUY9gR9Kp3u/4Db2xsLeRDBi/RKJFsWtnwi5YaE5uiOZ3gyowfnA2v
Umewflvg6avXELNBc/k1bNKBUpUg2F0TApfWkF7RHpkQmiof194hLPAWj4NWPyNu
S1qX51FCD6J9IAijnbqGQUInxek4l+54QDWEFalF+sxmacG7np7sqp6zs1GcUyQe
4vqyu+v11/qF5/HdYU+uX1OpxSi7oc9Xq2pOh6cmqF5r8skvvXrZ7wsIQ59Yk0SC
3FltU/HFfWW4FoHoI25MX2OqQ46eVL6ld+/XL0y8zUA3UjrapinaXUOuq/R6eumH
gM739bGKVLUPCbjLsFuOYQxyH+cP5BLJ8er0lS41svZe3N1UYhKSSPjy5Ob7jd8T
uPwnaFmw0oQw0d42cLoQso7KeiaODuEYFrI3vFyD+Ekvi/0H8NvrG8bwxIPTryXs
uX0evCevP5GcMOvLOnhNaFF2aLeOhrUN59e8IVatCxpMNnXvtc5Zg7C1tx2hAJ29
E5PyNrAYX/ujwOAuk3gvwum7ZO2WnUmOiEofK2cUsQ5sxKJgMx+AaY70fVm7hAri
r9Ks1Gk1PUdEJRqtuksYmSoNKjTG9t5LuITWKTwclg6UrCrN8ZA1B66ZX13+4VYl
KPOiJyxokL2LHtuEtwRSSNb5JHw6cSbOYFK52Ef+iVACA4whEzQvtkFzOm6EXqCR
hzXGHw1+aFkgTFsmwzrhJTF5gL0Veogik0mskc1TMK6gboELArqHl85mK7ANdF8b
QSC8NgsFvlIGhXStoeI7fAyEdwRcGMk38Bd+POElXMHw2dmbtNVKZK8GTe2a/wXw
xvLgWqahHWW5y4aInPPUkCE7PrIBaHLV7ZIVTkn4mTL+aYscycw+fcAWzFvGaYBp
G2b8cdgfeVFc8dJIhjBynxYzureBDzjUmEQmliRkMDkB5BabuuRWsamYp79BS8uo
DSpGexECRs3mlNvfDS9kP4YIeRpKUbhrG/a3+HElYZwKaHla1/+x917fzls8ot5U
8LWOiGpKr3ruQTkW0GrMcYUQ8dSSJ2cZBVHVGeNJzP+mujWbFxchV0r0ayFfKpuZ
HIQaITdwTjKYvIW5POqM1RwC7vtN7eIgp8T0wlhkviaRgEl0+3TBtkTq1dt6E6Mq
FCGE6yA1LJFJJsRoNSG7wX1kVZ5rpQ1bI7YsVXhq1YIplvak29TGq24OQYlU8nNT
XoqQRkW1stU0m2dYzb4PTWyEpSpot5cFKQw58PmyrpMATpE+5y+imgts0cV0uODq
/hEnGTddWY5ofKX69d7ch/4XU63KX1iWUhxeu8Y3o+57k+fdjCVqAqZCo2JnMtgY
6b7ExTkScfJxC1sSC6IIHQdSWMvo6E/PHAeZ5I/JCXGPXPg7UNOmPpQnOKUwSHz6
+FKKPAWl5f80b6hZgAhMo95DafwfrYGlLby96OKgHohBStoo0KzPFC1R9pF8yPZe
NqiccUPeNyzIaltZXn/6tErbAryIV+ve6UfWF0ckHkvbssWVTbyvpiMJ9yRbKXBE
7CjP2EQOgtxMZMYjQ0tgDZhvGy32nSAiJrV2LVUAie84esXgKUPO4tpuCPBLNumw
j2xPg7FRoaU0NU5X1d5WJvE2PghjitqRnj3WLOADQRDP6csoCQ5WcnNVnnxEQcBn
g8zFULqHuj74xA4x+icEv4mZnV6whw9JhUV3w2+Mr4XWkw80sveyDXQT9gXflnaW
juSPyLkAjeL090Kn2BJS00WaOiMn3MMMP7pXeELnfZP4tPNoD7z/o6RZOoHwdES7
mHuv7wHAq2nYSMipxcM0vnYILcGDKhHLrmzfq1j8yYpBLEnpNvAXhV0RZXtNiQ/x
ds5RbdQR+3FEJOp4opIfQtQmFcfcrFuSl/qQKoGI745vzkXposn+AwOIEy6BJQ+X
cxzGTuTe3O9qLp0thmVJ0VOxqEMfZKoXGV8txxmbN7Akxe157KfrI1mlt7fztR5V
FSQn/dW8D4bnoTR+zhOdcQMt42YS99q62o2TbwD1SMxtrDn9wUu4lpN0IlMhAJce
peEpK8KtNs4JI/8vFr6zUCkbEUOnF/idyqXq0EgqWBqWJ78D8T0W6A765Z2Pq1AC
bb7a/FHje9fm3mdhHlyrNqSCAURRSdVH5+NQlvLzdHWF+7FuHDfEag4Pl3epwAmA
ij3sSPF1nZe9pARcURo12IKczxY3Qlqgw5lC0i8aYwC9tmbhKQUjl5I3jvFs63X9
fXarWLxLrkEItTWJv1TMbBa46BENOk0+4BrEizk0VOcphpFc1tC/urSqpZLV03lK
1AP8j3qvnytYKs+x6Phzh1Mjxl8ovLnVPMfifEN5b9VO67oUQsZUOyKr/sSgqmPr
Us4vVW8J4/Mv65spvbxkZMczuAqZzB/JYjniIYQjWGdIWAcLJRCw6v0TqH4DzPk+
ua9niAIpYu1tSt1yeF7Wjp7VBEOaDOKrrGlQWpa3P7GC1pDbmqVw6TvzPkd8RV1g
uIe1BCqP8wC1lSIHUOnwdlHEhVnRRD69hpOJkJ0wOcZ0IzIzzxvN5rXA7SofPv8h
PRMgBID8T+OEgsMmakU24zf807ecv7zn+E0M2wVS+zA/bF0tQPpMC/0r6C5t6PHK
6/0iynIf4R3xJxjqx5JVlP/OXGExBatxU9Re0DR7LzR47pm3HjNI4iJLc+bX6cdu
C+CNpM8yA36QzjiovATJBPJkIuRi9tKb9Njrjh0psVKdIlTjSRxpE40V36lyH0rm
p9lYKdeH1luxuBe/yvuoUGe7eKYY+ZUG/aCKLmd5FbKqxlOBC6Ljvp9rTeS6HhXR
k4cJ0tsD/OFZXTC3Y7voCIEnGsk/Lxjz4nygat5X0Pflcx6sVeBiHIJ2RgQIdZPf
aVntpFYlZf5s9zSEZ2DHu551iBaWzcb7iziZoG0LzuxcwH2t2bnndHD4raAEXkPx
lLWWX6nuvsMwDH2Hjf7xN+syNG3QyMRyi3YH1HhOPtKSX9RjYw7b5OBlip2sF62r
aSCeGS4B4xOSleYUidXyNybpUonngkXkhR84/B3j7FIElv9a0YKo6KWJmlGCXDf0
vfSV/XzYul7LT4fJAASKlMB5+3QnsTLw5E2Po7U/f9xioADb8wG1rDIgOfbEPqrw
owR+ewJ6a7UV/GxQSWhGTclAYGI7LDto1/Qu+O2HJOIBEVn11m4opoJg/SfKDdNy
/9P/3ZpEYMQbGw6otPk3JXYp1O7QLSZwcUZ/LT3ZJF93UppGorRRC0YZydcv73L4
tMxDfqDHBFKmwYfpw+2IAP2vkXQ8OrpPTFUVaFTv0P8tSnap4ftbz80IG5d6eVGn
ye0eE9YWhuA6fEr3FJc+fKNJ1sczNXJRKywJhAz/FUFB8ZnYyNzaLw/YBXGr1pPA
c2G7m4G2OS6orKUCe4jNQZvUXb/Ob94lPYDX+O7B8CaGvlRxlJzw73EhYzLJ1GMt
VPfEdUi4Jki2p5LFxYI2PQHkYgIigAMEqljQz4zPq2WRQkkF5JtaIteiVSRuWTjn
is3VyOQwtR2C1IpixvVcBdbI4oanudnyUxIvJjtIfhWfVNC3qkPhMiA3ewh9Vv+h
hzvH1Ehn833JNuelOk7b/mr2WROGagIxQOSUJOJ/BZiOuwNJqtVSXth+jzEEjqoI
nYuxjHL9sxcE5xX/RxdZBgQy+c+YlrC7N4ZDDJUKyrXxsKbcjAmz1LULIHDSZtB5
xL8Ge50QBeAgkVgtc4TWkMkXmZpjcY+RdeJqzgkXaUsHngwIQNu8bQjPcs9NjOP+
AqPUzL5IolX4V9K7/RwZoSsbXSbWaz9+kiwd65MBTgTLzUdqmYqdfiEVyMbOdChN
fMeeGPFozzkh5cutfICZPH2frg5pHawo4o8FEfXY1vRSxlxZ3hiclQAMheECY8Ma
dcvtanEe3AH4F3Loo+7JSDYqIyBnEW1EGLpme2jH7AfT4aLM6GwI9M6OZ2ccUZTZ
M7uBl/luoyDXPWZ4ZJieKcwFPQAlLBBmdxLEPpLLjbTpJVyb0/TIuRR9js65NksI
SdwpwpPmGDi/zHHvmzev2fs5Mi19pVVpZyLHfbFsi8qhImj+UJguI11GvuhmW839
ysz/Ib0/tWtkOUan0WHoAzFDj9x0BXNvH9gdewGSgbMho3c5H1JnNBkMKlv0Wv0B
3wtlwoux1exXknFOYRLikHvMPg3hXmR5NKJiywgawNM07FuiIoa2bR5lnXsYdNKD
wiyxlxZyt3n4dX/8H7xd3jLjByvVEXQVpkI2XYcASDOcSh4G6EcV6+4YTWZ5eCQU
9R+WWJBrgs+0cni7JQYFErSnLWPaJE0AfZnji7it+zcvSJOz3QZBNUu6/8rjbIHN
2kL8W00L3hxHLenpyjtytzHkljxaI1R1Kn20Qmplg9io6mFgOUdXJAipWBKxOpNy
Cn3sLG3nqvAlS5AXtHJhW4iYWdmPaK7hIerL7UmJV3RdGYm7+oWuPrStmG7RrD87
/fzlq5c0/0lQPxLyLnzaWuu2LQFtI9jY+hXDIyVdEzttvyMAnJ2IHW06Q4H37ely
3nIpnM+N+ebkH+I/lIrlQ3rG1K3MfEUqVMc/kVPb8FOj/T8/3oC8dYIzai/p05rL
7mW5jXN8+QmKcWedFiqGbIujw6ktQicbklpgSLF4FAnKGcRDYBOMsUi4Z+S6EkfC
uYlO9BCJiOo9hRg9XYAgBX45NfubsUCwJGJK7TF8vfwsYhcjdkH3dXnSqfSpYxOH
r9/8DHFk/dBkCrHSPoca/ljJqcaCzKtGKJhZvqmfk6/k4knjjlBlBXBcHNf7jTvB
9Dz4x/YLmjzUXbVeT5yIQfwAZe/PV2znEq6FiYdYsxyZuG8Drfw/aRUaPRkjxz/Z
qNpvaxgx1d+CbQ8wEM0dx/n1SMVxu4/8i6NzJlnBZ3mCGZfOoAOVo+uXtGbCA+e0
/jtlWyJJxrC4BtkFOn2Tj+3lPplmzr3i9ob+y7jQ/NRIcVMGvbW0SMxhie5unbWE
8hym7BbtAEq3MIXQ6eV8Ar3YS0Bh1JrJS/B1/4cwZYmNMo0xx7nRw8QakFHPD0yO
eS3flVIuLGWO43+1RmKHwRVO5/5pt00qsyBfqkYsRvLjqatFSkqrYy/3JpDx86Hh
Lii7gKk7ycfWMxEjGlBM+pQP37L0Cf3r8iHniHb3cQ1PeneECHiMuXJfL8z1E821
BDWg1Ccorp0FNV1vSKWzJnPH1bs4Ls5K85GxiJfClj3nX8q3DIUIpuqrEA8t/Pxv
rq9mi84HHPxvozfhwbI5ciMAjjPL3nkll+p71nzmkiyvQNY6uNyBU5zLCt4i1O3b
Ny+nbC7sCygqcfNHJ6vpGG9kKp5CoWA8mW//GFYyX7t0duH3dXp3XarRDgxgW6vd
OXQtcFUcLU9d9BRM9GlyWdsXCK+iQPcyYzaJ3rZ3VZ8NirDuNSw35PbN4UCFcGAO
VEsF70Ju/kKS5La2AwDG4Sn2pQ5cLn18m/6PElNjs/wE08MsJXPJCF8Z8oBaGhri
p7anBNqvq858Y36jzKy/zK0V4Fmi3sFcDZxM5ZYmyLeXgwa0Nqpku66ydGlgQVo4
ubY0OB65pbbZCxNQIcIMsFMAUC23QAFIeMpwcv9OWSjfqZ/ZuCJAqPjbUfNBYgfG
aiF+CqMiolTpWxVsMhHJlrZqrywfklU9yP6mebR0V1yTsYmYLIsa6t7zciMEk8mP
kxIiY0C4mN3fZM5mUnIa5XJTvs2uA0ALFOEb1c0fhyI6oezetjOPILz5Yln4+hxG
Pxt9dU/bHrlTseQ3G3QwS5EOv9KJgzkCmp0sENtBSQ7pYB23YCYVEEr+ZN20Mbl9
dc7C+GEqIyJ+FFfy09iWLBdD482ldi0cUCGUPZ/4y8p9s2HL/uO/DH/6OdlsuCOc
F40FXIJB9U+Yg/mnNMFMlxHJN4HEwtVYIieq0Kx5frH8oWBSBvibKKx4nmw8T2Ee
gbvfL6gT8f+e789VmKMCjk41FT3Ow4kzJgUtMoonH1+nviDs1Ms2yTJWGtFnos1t
d+Ra1rJDwxoHYMf54AHPaIAncgMG4nf+NCSfUQ2wOfahuyBGoQS1KSHmdYi9CD/v
MmGYfZW9VfIzuaDUQTDVUNgr6w7hZUS+I7/GEwZXONx1YGl21CA31A2nCuMLwYhP
8+PHo5z8ug/uY9hEa3eiIKc9B1irxnWmClXrqSsvknS9jr7uc+SVE1Ur34/iOk/8
IIauYtxGws4UBwAni/AuYZqKQwRZDZRrMtLbKQTvpJOK5TKwfeR8gTJAv8AQdDRR
GYDbMzQfIl1Y3fPupVk1Jp3zRZtmv6A7TxoKgndMkSkeFYtMjgHTMDNutVIvOs9D
jSGQkV1S6ugxSDb5ZSyUYKCP5Layt+tnIOB8R9pHH9P893ileVUT+vk64VazaDVW
zhcYPLXU/B/nivzTNEvApp+ng6NxDqnHS7vm1IXq0DLD1jtOAfYXyRXlnd85PIs1
itDhuLm7krYLc1tXqgF168ALr3LfGaTem724+4NwFQYrhNarF7r1U/E7zATm66XT
ZoZj2Ze/4RTMmuPTJLhne+uFzmE5pnJTy/QSukCPdXJe2QEY6Bzy0+vJHf0zvor8
1IzVAN+aPE9Vjll1r/mv5n0DmAsvatdE+SLtWsFe83B642BsGsQtwKIUNDNywwMk
1gJUZCQ0xHjX7sCCrdBG/ZLrpUopdcx6NJaOldYS1E2Wv9S03oPGO+gNCKV4aBbY
knClN4LyMp8dPpuiP/t2prU0eATcOZH+FFqKXVTUrz7JaxDNleDBIQC5GPewCMVF
SFfI/PAgNVR3Pkc6TkGqK4UcGT1ZcTkNiCGbNVfZihTpQejpBrNEimXySenTlIgM
FLH6WoOLPAzzHHI2EEHaKdDhOwbkEqt8WpTIykDnJgvsYGM8L5OJBkyv1S+paVMQ
G4wRBoIDVw5Rp3iGqkcIgHjcr6wIk85VIicz9/yZR42abfez5xRmMEcF2YDbkODz
S+uf5HtOKjZQAzMvPNp6BLlMVf74QUFbvSrVRSt7QjI4Ljv55HCbqo7/e00vLCwE
VaTB9DaBnfHft0sKi4hfURDKjnLgrQ09vhBSwiDhLKOOLC89jWKWNyaZyJb1hyoB
Sif9S64xY/5ok/MbT4mP1j7VdqI1WE6EykNI/x2U2Dglqf4/Dm5oD/KT/RGnRj/7
fpihOvWCfE1DHTKsPVqdwUC+/jdZppYEs+KulOcpMLoMRzWb+mALfdJtzjlJ9iz6
Yv681JXQzsSchhcwL7hP1AZqvgdN9fXIDJhs6npFlqoRvGDi6Yd4h5a3B9B7bmTD
B6on/4NE6KVElsGp7BS0/Dh8Kv8HqDdM7Utfi93t4vdWNtxJJERn9hNvH/k3d5vy
m6zX0LencVY9pyjoz8WdM2t9lc+djvhEm2rqtKmYmgmYwitKQqC0l7ntLNbu0Lcy
4nRaa8uqMLG38k2kezNfmF5nTjxqIoDcQ2P1/IuJFZZX3P11TQXJCTC+P71vhM+Q
jOiESoOMfJ7MKUibZvAPlZOx8kzpWxcaEVDlVsOrFh3CZRd6ojGi19yK1J2OeT3g
0XXaHyNVVTPMvL9l3m4NVihc4J4DLrbjTtIIE8xgNVRv0HO818WA4q3i7cVsziNh
zB9Aw6iRmPuwIPHyxBZALAAKD5/OT8iupqWx0lhfIa8YSxD4vH826ThOpYY8duoS
VjTJQ6w7/TzCoZfumkCeZ+CztRUyAxoZF9Q5MGSd1j8B8WjA8jZkaHW3M3Vg/2rX
NlSb93wtzYFzujbEiu3K9dGaVn2qzUNSlMcIa/Q5WYHwwQ8gSadHZasCP1fSHieM
5IVR/sZvM30amBgNKzvlewSK4TrVq1f22YvQjVZVxiPz7iFwzaVmacqM7cC2YZfk
hd1W7cCdhoc/PUP37Z0z9Dy+jmpG6Tkc+3AhEsklTVqvB98FH/czMzQNwtNzifyF
OHfv1BSefTLZQ6KqniTg4/40sQf9YS84PWuhmtEM0LSuOE39+Drh5SMXI729G7QE
61RVtxx12zM1FAiPtaRNZXgqOmTsUbmrwMPuSW/53965DZEgOo9ur9755LGU8eql
rNJ0IpoWWl6/xrIn2xOS7iyTUtoW4FssI1hmBwzo9kQnU2ic/mF09C9vPmo3cSCK
fiFvXjWYVBsv65DZ5lz7fPk6tIRtmWzuI0YigJZijxd2G4uu97aQ0M/ZMXzkVJXv
8YtYc2hpIysxvALIAQlbRt353p+elnfUrkwbCBFOCTftKYrZDwQ2cbpwzTVZ7L50
VRqWiTz/K8fcNrFRZ0MdxcQufViIES1twd8QPFpHVZBORL0RYHW+gT20CSAzLd4T
s23z7iu+X4mfGnSakE/vAEBGt1mSeYVEJE+efByhOPxh1dj8fT+QEevDcNpIkw5o
JGaojerMHd4E+qWRTZ6CqtLAYJNVQyS/1uikixPFqsEyOj9od5o5LsCp35c5cqTp
IkkpM6J2b0jqSMmN1IEVWfqFcz75k/NoPQEGy8smWcYexYrmgEELtAysl4/J1T13
4kUNtgDTg1o53Cy+t73tzCRUSS9gna0DzM0Foz4NAz5UtN0bjYkH7KvbTp92dEIK
nzXuT+9STzamrTfowxX4nSqhcEurCgq916/zLdrSIAF9MgXzueNTEvEW43B4GQgm
lhf+W3jdtvvlCmdDmqu/4zu4qkDmF+e9vp6h9huHJub62tOUG6k65abQH1WkfnPg
adUu+3/jJw8a3Awl/VAK9a2XyZHfwis6A/ELrpS7swnYqKyGpM071OMb8RD/JVBg
9mA8Twdj8In7iopeLVLeXqNQIMzfT2ScSUhWvdFGLXpe5fBb1BDHa8dWrp192Bvt
+s7UMefQpZSYmQHgj1J4cjuUx47yajRHIrzqSXfPV6XQ69QHBqurLCM7VQfeRiYp
MUiBsxEPDOkx8eLUbOI9bp3UgZoMvwdBJxqMcMhSi9cWo5tUAbeW6CrX7N2jMj4a
7MLoKafFbQGw/Wuq15wLwIWs8tpMOOQX5SlUuVXWjBgR0AhdUuCrQou4SnJamF6k
09XL0gCsuPt9fMOJknB3iTvMZ7eA35bm1iUaSWa9jaMzweffgZgRSS0emA/pHqob
TD9qHXNLiYUPVbzX3WRuKADU2WGKk0DELCDw2RoVNiJtLS02tD9CUBf3EpObTq1T
uR2OtDHECsgXiD4TxJSn/ep58zmz7TfkwddhsPO/7+6Ud9Fhj3rn/l/zRQFCKxKg
J6K8794nRV3zawMarJazpU/IxZ+3MnNixNbouhubqyMZUl5BKoappw2ayHl9Yan3
JhuKJEnDq567zJ8BX4O3LZGpZ/76rpckE3fFsQWREtDcZWdmIr2JEjODvt0ckPxJ
rz1v6CYQ/nIfnWuJZnouyheeAQxtm4sNG0L76XcchCy4w2KVCM3NtW1hrJ5GyGmG
AzeMZwqIckX1S6OW9ol7+KWkRyd3oq5xFx1vsSfd+/oUPkvBeA1ZZwpYykbVpEPS
dTW5vCgXsTthhc+agq0XNLOrSPbsypuLpKrc5rH1CfP0PXvjFWSO3RQbL95iOROB
Fmn2OR3NiwVvo8ORlgMWidTlqDtTsgp1euQb+zIoRdp4D9zmR2LeEMMeCUfs3hNp
UimngnY5xyRHYURk9LJoHeLiYOJiORrW2DBF2Ztav6ITUm42tqZAIGVJalwWj8I7
4lM9z0UslJhtAmsYeC+DC9U5nlP0lkNgkQFyMjqulh3URErH/dXlVG9Duz7xQros
FOMZnndCwi98FbUGC+ek4TvZ1/+r3QTpEy7bdFRiyaVx0OdcJzQNxUJQ5PZYK0SA
GXEE2HE4qQVPYjpAML+ClMknrbUiywMwbqhlzX4Z0NUziTeSL1G6ZKOHQTr3jXc/
wOndC2OR6jy6Ust6gEbG3zkTZURDtBqc+EYo8z8Yq7D5AG531GfTyIUiMG6pAyKX
Fgd4BEtNQuzW0mmJ+w/WKRdEUt5oragtIQZOXMSHtYWuBB5ARgC16e+Ewbf2Nuw1
VoIRmQDavCsm4zWnsih76JbhRMOYvPQCpA+hhQFuYN1V4ijSCFo1Z1vywbfgAQ2h
E7VcwAI7jsjXvCqinNWZbN0OcwUbu3TsLsLBOq0OVdT8sHMSk7LaDwHudwSMZplv
GzNE+x9PeKF9lq2uO7dVPx6kUY6Hdqzj+/CLzbljN2kYV/agyjWjmfbm93pa/HfD
4i67T1oM2ZflNlJJiQJXdo5qftUZygRiOlpzc1OOce0I3aYKtt+pkRslH27rp2B/
9X6HITiR3IrkVIMp1K1eCSiHDUH0hJQysuYBK/5B9youEY6H1KAi241w4gotqL5J
9jjYcKzo+KG1x5X6RUlZXqePzktm1gzad32UeZkfFhDcaPZ31VIo2o01htXGSjca
l+ieDlcdDH4wnNV4Y1h6IMhfq3ggxpkvAMXae5Sl9hInb5bDklstZ7pzB4ZJMFG8
iRk1tBLlLaPbb1Hf8zYxIu5tgTblATiMH1zRiyV1iPv+FQLIDPWocRVjPYzojhmv
LVeB7B8xhyEGIK1+YlGvW7zM3XaZ5uYPLB6A8uBDB19MzerVM9+i+AUCTnuBY5DJ
kvfRt6jPBVLQ54MznNcERO1CvoUnrzl4gp29PZclQmcO35CTJxWhSw3sbtSEj3iX
8zdoBz+e04sel0jA2qqTg2V95ALhdvKM8KFX87BK8rHtH9eXKpfmHNS81aZpYt/a
mzQkjviy5P5kXvfeYaAp2g77IMl73oqdJeIogk5qQnHdsOcVx4zB4w85uLe+NGtD
r2/cG+mMmTplYkqShWERDtfqXJBCv6StNcYiULzjGEkxMA2nzxRgth6JrVbdM9vj
jXM0WJBENUd3F5KGzatsAy9jDjCy24OfukwIV8t0TGzOxoTvOhgqC9IlZ4vkn5Ft
gRn3GFRyDF8iNS6UOrjPieLM7txDZEka6DVGttFefoUyGhifIZ+2I4HFTbuuDDx9
GQ3R5h2G18VCLkE0dkUp/01BzAMonmVsPKrrF09Y43shX7nJPUJOktN6Vhck2a0w
+/zTlvAzacDo9MDb2NXvNo5QYlb9I+aU6eEfpgRAskPOoov8RjQrIfjXGWsobTGV
R0SQattMEkTpOZnWiRB9HN41d/R7M4Bq1B81/wHydCPcBxh6T/akSA1G47hbaGj4
T7FIEXAj6W2u8i6l5Ao4RgJAKOEoH8zVTgwDhR2nHId3yOqWYPyxN/oiNyiyL+8S
I7hYH3nTWLoG50eEiEklmEUUZ4fYEE36lIB/KXXkWf3tGguHnxfjCWA9F3awQJ22
p2pb3GsC4IKnSPT9Rcxlh3Qs55Jz8h9c0yeIFJGTP2so75D4ZkN9JX/iYJJb1AHl
7glMhdAGpKU4XpCdX745OckLYpgVv28TdslJCS3kLXE5SOyrIINFZtf5w5KVr1cR
CTtWozsyPtrMclhlDK4wA1x9iCKBPfXuTFUXm+ZtwZ6+IhXgIOxkdl0vvNKZ0+gZ
xhZLrL544BwgFi+lPTw4+8oJsk7+fuLbnlu4GZr9J3PxdXLTx7OBM9GMNSDeO78O
udRSy78c9NpcXCUeGbfM9zyaGlAsdKPPgsW0iJKgW+AiULTwDnSfJPqOrRFR5ixk
hMtS6cH3A5B9Tpq4YF1SDGb8B7gCaLvTMFA89Dhb2OWBqSod5AWsE6488etb0hfe
eFOY/a0yapOmRGetX6/0JvtPa9sBYSrws2Lv6fVc5pMXaODsuCEe65+7g6DYq1yi
FrzCrK23B2t4Rt5Y2hra8yh6qmXPb3DEat+dEJRvB2uqCt1ZUQMaFH+R5j23olPv
KbOq4/JnKbaHUp+69YG1jlzAE1Id93cGg6a+Pa5re99fIyuz2A+is7Hvefhb0WZD
3ht/MzRcc91OTQKHFZLUEbJe5U6unJmfWuxSF+/21LrXcik2x+5lGL/NG/K1R1em
fYT02kNoZr1uuAXeIglQqowfVJGfDwSHky2luoOqt/7oWtZRaOQl8k+dJs0Ztb5W
F99Cbpu+jUdq0BMCcIBZgVIOVVVeeySe9V+9UV5bnEDPIRh4K9SAaZUJM1klOwH7
8wYW+UXiBdyZj8AVJkJWYh1ycf8L4j2SvOLpYL5zgefbwybweago69QVbd93qXJx
bVHPerRlJOlXyRuRJelvwSDob+02Q+HX9DyMcwIZBqu0uFmYly7Qtl5E6rsuiYov
VkNiUKFiUZbX1txhjX7x88/gdQtyciPGOcDC5ARikDQRy349x2SCJi2fJaQZfQc4
IBEmUprE++l+YR0+n4SGFpP9DBleCp1Ga3eDPYtrJaDjyAB85JlAKMZ4p2z34DFM
9YfJum/2eNuCsOg4d2GPslGYHhH5i/RaiCaGOemf28s0YwE8DblGj3E5w026OYjF
sn9jQuaf45ygGWNXuHKCzoAoF5rFnaKsD1b/huwHkXYYia0GZjiBGO2KLBo65WBP
/uZ3O98c95YPsfyd1n5Q6Ul/O5AYO7IGtVPoyRLrMf5hsyR5dOzdXIZGDfcZzPpf
xLJdQeQEt54dkOsh0JMZgXEEDkVisYSZRWci9uARkAEoC52qrzCS5qLTz4LgL6Op
yVqF0MZqX/V1lRTNsoyYaU9bWfCn4bBu/alLb8jyok8J14FcTXnnTZzaiUiRy/HY
paM0XkooqyCVijY5w3EKB01va2DPm6PwbXHKHI1pKE851mDOiG4XWUior/H4HGSt
6hbBPHjJ6SPenqXX36DlRynwv+2JCUZ98zoIrAKjc37xzlm0xaNOLkd+yl7tsdx0
Kke009Ith+3ii5UhrV6Nrp5HyYRZSZRhSRuqERueLhZfbJRBGbQTwMHqjkkIfpon
eRD5LJDKY86f1ZY6c1VNkpb17C8g0OChJIiGpG0LNxkre5QUAZGJR2ngBlKjBOhu
1hoGN8RCcwfdblYk2K/eZaugJ7P0b3Y+9rkUzami/SUsy9PB2gFYjPOpILXVd644
M54+K9rUPXbmHM43QqDaHQ9SGt8fa9nBuCaYbRRX8so24pTlqfNkDYhbS3eFqmp6
tYOjUC3Gydg2X3X5N4WDxTYdRqZQlD1unbA0zEtRGen1SEGTwBq1H4kH2LXw8SGb
jgNaBwBolzf1O9BLr+vfdUMwmjri8YX17kyli7s7jDVUUn58EUIQktxrnx2m+nNS
UlpnM49Sel642Cjwn+888tL4Dj/5a/hMX5eCrD9mt2AijIplcfZmrGslHlsW3VkD
u20B3NpAgxPKZ4RrOZ3DXzT6AX9ztTGgJie9MPgHT9yqBm0jm81YhQ+gbQqMGMfP
wq9JqoqkwIWsYyOzS/oVwpQEWMyufYGIqc2Qh2aH1sMLajPq4Ah9JKhRTYQJcI+I
RYPR3fl2gbv6/YzyRPWqcqYkn3vqyu87PeVGzAQ7AHpXX2GWDDnotXVJsTVrn6f/
p52t4dgZHyqVRQxwcgiC/UbHC10Hvpk3zT1tawRtBWKdP5B4FkkRp84bgfAqDrZe
lOBvX4T+GOIxw0kegXbR5XdGDHg+7+zhdxi6yNjaTPMTATfW/mR/KO7avoHA2uwh
K4plXlZSn4owAfPyhdmcTIHozBxAZ7CWwW+HR73or+AUYqPPDvD45zDFG/fILa6H
jngnpuQySK7Q2+UG+f0liM6KKlamn8uOXEhTySG9HubyTRR2zU7vFe70gROji2SI
qpRIH2bzgs6Os3L6txBaXgjSe94DO7ISyuDyc1chBqi+81K7HZxedzExUrn/XyM0
msEg0+xqGBd2J36Mxv8jNghqDAUixcb/2+cOCQH1DvIWybympfDyVCNDoG/+pjDy
qApTgxV8MCEDBwWwBmAhUAgWgXzYMnvnuVSSOCdWYKJRCLiFOJd1p2pzSrvzbLl9
lrCGL75wjtI0hQCToGmF+HsaBgVgDTkuzO0qlRbYqAKIZfU92rc5vSxnT69LdBQ3
FgMqxJe5nI+ZmnoZO4UpkGlrzplMgY0E+F65AkdYdGnYv+BmyrXqBqYL8zHyt5cH
hsVi79V2D50hK3umDQekg3ihxtgO3BqjJrgLbwiVzxs3IYajHiHXo4XyeAuex9BI
AoDCcxuFArsIK66Pt4pcNCInYRfhJEGlbmdJeQQGH4FzNVxdTabLVaSP8buo1OoE
CBcmv8h1KMIYPTBOdt34W2beN/Torc8WpjTRkrls6nme+J0YmA1ZOQXuPMEzwTgE
mCwJa+I6A5KYY0CZNNHx24zumJhisHW8K576ezyikEyYd/dXUBz1H9LHn643D4C8
2hhgmgSEgtOsqgUbfw6nqG9FuNXHBl+xgZbvp+vwtkvQgmHzNMo6J1BkVMB66Y68
i8FYBmSQO/fbvrgPEqywh86DQsdSO4iFKcVy0UH/b5n1teOCghbbg2MNbpFD14Wp
4yeCNzNyuBMaN+GRBM49Kt1dZ/OG1YGZvla9rHWCckoFnhfFTqdi7R+yCtZZlf4b
kiYWk81RRxJmub+hHSm1FuBg1/978CnuDziNIzTI4VWINyxYVrJng8DxKVgMVk5I
cFxl5/6Jv/XBoUlHI24Wc+nMMEDN8FG3ZdNKNTuei5RqwQWlwn0hfdSEaADm3XKI
wiSppTkrpty+h2keUJ9QZ+FZqQIDxYJx9zp7nEhkhX5lZlBKDLxVuTJug7hrd+Qi
RPJNYiAeCY1uV+++Cglr3MRMQf08E9rFSosaXue5cJNCO7XNeOgrDqCRJnP6TJ9R
xWwlzroAJ8+byUoHtQcDvZJ87RJVQuXbw1FHncsuAZjYdtz+m2vzaOMvkB0SAeF/
ZpZbagwa/6LCQTmo2C5Yw7gK/wtCZ2v7HIecxGNFZlYizkJ3Vzr1n0t+fJtXBKY5
1Y16N5+HM5hT0xXY5cXY2rE7krLyfGYalhvl/A0u9i0rXzBTo9+CYXBqhtcvX9sz
J+fZ1FkEFRliUbDLDd9l0u2tXxP0hGe0u4tR4l4ePcYHfBXCjY4KwfimR/Cgfnlx
zXDsuVt69YTQIl7J+Y+Fq+AG3c7gx9ifokhtM2HMCnO5Le9Rd6avd0PhYRMpWgzL
58n7CLFtffdhRit6xgXcqt3NJMqpVc+aqq1Gq5WYAKvih/tvoVG0yP3IbP7TTVbg
th8aX9/dvgf0zFbEp0d9o9BYcXIkTT75qJ2oFynlocnYZmP8y07WChPKUxEWnypQ
hadm+GWR+DBu3TQ+s95bhEF8elClm0vADcJNxI/RbOccAEfzdcW79S5oKo/o6Kpm
k5KiF2aBqdrhmuKzL4NUKK8xJDlLC5J5uGGdIyBR5WLUyz9n8jPqwSmndzxgTw/7
hrDPvOv1///KxdXjBvOgEZ488tUZcwVBSbs2a5Op7UevzNSsrZ38F7cvPbUbhoPF
s/nwCfl55z2GxrHpuOsBLQ4QX6F6W0lteYRTr/RBraahyiw07gXbxt7Z5Ymo3NFr
p/LGINfInbpIZCz3NAVW9ARUF80tt1XsHQQpo9as8Re3GQlrOuEpgeS+MDwZ4MCt
o/Cjm/dmRqR6YvpWcBsr17NZOsddNV+HZaA+oOtVlQ5Rb2DEoqcWxoHKsIw3+8ZB
E+7vU9da/QGob+UJ6fUIXCWuYxqUFuAyD+nxU60PV+WgIVu++E3nAZeFYiv5d7gR
wYqExNgYnPw/x6h5h5wQ/WZbuuzakitclMhc7/7sGLi6148qyLLnSjXHV961zota
FMzkrpxh4m2SqNzcGsBOJEwBjWT062W3XEEI7zG2PZv+AIitsHDe1NiQWVZ0jR6W
HR5GOVkqsHC9dX2zdKN9kMiQ0+8wfs3Ij5shJDmCF0u0nDTCKMxKn1aqAqDQIqZZ
7uq8148TkQt+ToQhi5SGxVTiKDatlOeT8Xy3NwFjv7deA9sbKYk6lklRzTFi7MsJ
5NfrkNSA6o5ckhIfgxFhZFLPR9ytGoKc0aysnKI4G/nusAg8cvwH57HhDTzQOXx3
Anjx8zaChJd//AqoXy/BSxw1Bsx0FXI4qvpQpYca8xJsAwaQ82oG5QMJbmlDyjPZ
gY3WIk9Ym/qcMPWydPbdDxMyXqLfyP59Ko6QFJRA8gsNdg/0FmpM/LNH9d0S8CEv
zidLBJFH5OqcXHc2B/Ec7tKLFNGnFgAeYP+g5yGv1L8pEDJzlYzB288pNHPCuMzZ
iFkvgRC8Mo/ZFw3fdf49LwwfDmcIXils0RARrj5D0M60Q7L19lxY5RhaZ51NedT+
DCha5Ih4xx9E/41n/ixkHWHvKkmMWnBy/6KbE8a8ReUUl22r0MitbISA/D+VV401
bq5NqfMsLcOQjBtTFtONytP8yqXnmsx3SywFQPMvejLcx7MZ7elRxmkMnrGr2amK
MI2w8gj0r6wD+YQTWYi3gfxMKjcijQl5CDdZIR/XSDG31qeWyk8sCqagq49B6/DQ
h4lettLFCsfLjxD0cegQGBu23apsxVBMeqOjMPgYE0ck91Zfy3sLORg7TbWNbgfJ
fS8gwSLG3p0Tvoh6Rc5QdTHmF2ui/JHeaiy+1Hb1CJGnX8L+8Yd77Beko3Sf7Jx4
MfKP/z+LwN8v9A7u2tlnj6c1bDDRgq9mLtZB8+CqFZOuLrsl9CjavSQKg/f8Dmo6
Z1n+YMdWU0Kxaq1sxBYZMPQxzhYOQqa5JltFCuTuFZk44Pv4Po5fqTG1OQJvjm41
X18EECIpbx0SPUS1N16OUlsBZYEqdAJMQzlbx/K5hMw8MEuwBSgzFLFGlRWmo+v+
oDl0kcB1iwOsc5CyC2l3S47TSxYfTXhSHhfE8kizT2Q7Cxn2sNreg46UQbBHFlq5
evVqVqmxFHJ/C7X5TIxGEYGICBa6+lej+oJcoDn8QypBZUIf3dwH9BoDSqs5Qizp
eYHQysRyfUIWf7mKT/3uXV4mYqAFanGN/eLNqAKHBRKjJkB+7rbhCIlPyA95o95D
oYxbdn/DNDKuc/mUMNQNRfMmXXOUXLPpxgWnJ9otOQOIsYD42SdXdVJuSrEJDhmj
7HQT98cfTvpmS2GtKHtxIE6nkpA2Qx7P5CijGsF6qzBTIvLgFY0h3QmyLnGugkeq
gJilA9hZDH3YVfKQw6bZX9L+2AtOjVkNC9F+n+J4RkMtyOuSY2wzt8T6lnQnaCTC
QGMgbM1UfBVp7i2KUluf+k+7fIpRsqv/RZGg7pMyhARQ/l6thTTPnoLj+nRj4aw0
pQlUCBa+p35vzFAsQ9ioGiVv8vcPhIPTplSUaJV5E/Nq/JOvkgOwRbJ4rRItts/a
EJu/1qrzi16DEJKjkDupTTawsDg4tXSxL7CWTA/47LfpLngWE0gAi7AF81MXn+R0
+mzfNFE/c7lUjJcJOz2DF9wXd8zVybfeEmnI3+QW4WJrefsqXTsG/OqSsLlYOOcZ
p+uwLzm5pxe4TEmPyHJYqPz8HA9yeYWJwWH4xCGcRSW6hI4ba4djDvxUIciX1Gfh
5uZT3lFX+HCvJYon9WbshlkCmqySbQdzvPmj+lq2PbL+4rVLhr9V05D9+kVQnkNK
SB6gOTADEjTdiTgaZ9dbHuTqtryHawFQ90yUkjYWPqd8InODvXY226gUOkWvMvkA
3zxl2/X3ZKv4MJt/dfHXaMsSGzvvcvpRGRBQftD8kK1BVKv+NGPabQjx9762uAGk
ZJpLrFLCxqC5CJDaliY17eszOb25XGFLRsuz0Gq0VoqQCP1v/dwSCcbc2aUejJHC
bmJJzelhZP8IbBogAq3LxCzQYjQxGi9CWIW1GvRpv4TKSgnmMQE12AXnVp10G0MU
iM2x5l5dtNax+A854hR9cRnsRPhosAxocQyAsMADc3dvHXu4JLxekAkKKMNyHdJc
2Wu1dhfpCenb7q5RpOV9KZjglI8a0OucZjqYoz/I1oOudpxqcR8+LywUi599Q6Yg
rOQmTYnAweYykvSwh9Qz9/Oou7yY2WWKZz2lar5/zXlVi09cMCBJC5GmD00OdF3j
+NiVdO87l/tH/IMaDodT/4n9BojO8l8TCt28HWwD7XRA9j+Ky6gnINwP9EhN9x6y
cPaBDOZqSymwoIgbvZHZPQYG3EcFWFEyG8eCp+x4MMfxlLFjNHXhyquF+hyJI8Am
mKfWqmaKzkBqsJ7+ljA5AvIhQrVHOczm6nT1w6jmOkzTCQXh55EAoPWTOLTMzsZr
R7JHwFybML6PsKrw7eXQ+lBlBjjaXOHhlsIUpa9Cuznez1Klpqorroz1U1Z9G49E
ZafUUVNANtLsqOE39778iBs6D2Q5rCYyuG0EFozyI66d3ZSTwQ6aKbdBvzUlmefQ
z+PNOh9xbOQP3cgviHPDclQdGIvGNqjcvCImoXF+nxgKWW5OMBdUiK1XbkavdklG
Gai2fYwoPlpMWx6tR1mHcpEYWfTrd5zXeLLnw+zS/qHGRgHiYHLF4rutfdHW63Ax
Faa/ugaKHsXae02Tg3ZQX2JpzgUVGhrNVNHvOu7/iU7w9NoA5wRhGJhcAqz+SiLt
efdOPf7idZg2C4AwhOWvRDWBtnOBGh0Xwrznei9FTHagqeDOwXCiMMxA73QlVW20
cok2jMKhJR0b2OUI6HTeIzUaFgj6bU7xr0HbwdmGxxvkZKMsG1PKScUy9I3WpUoW
Jl9kXP16HN/zcyWBf8AIj1XCwmWyCbw/pB2rkZ3kAJZis35mfvvhWqJ9Yrvvl/f4
DDu2HMnoAyQSXimQSeL1MhEuajl1E9T2ouvRaDc11vzwCNi4zs2471APqvbM4JHQ
NTn9cjhi4zONqGU0vGdA6L/DpLdnwhvxtoo3BCgKpV0dNvXb93bSPkdm+kPSXYFv
muQtZislZjdw6kcW2/tpKahBWvqU/6AF2tId1917xfpyWWyzSkBwtmIgXJARa4mw
ZgWV2WhjhHnJeRThM/Mcok3GtaIGCLQO6QhX0n3Z+L0rnRXMJ1CYE7hBAPbK6tFD
2bxTqmTmauOsqzZsBoTeBt1kr/Jyd+n09BS+qssLN8SVON+QvLAVFBHa1TwVf5H5
qELGbY5C5M2KFEXPk/7r+XMd9QxUS0YGY9VLDHLVGZetNZng4TqWgTHz+g/56eE6
Is2my3E3voRGenegwmIXGGQFTi5wChlZ1lj0SIS+pgHOwBHI1A7RP80uLb/V+vep
XJMCXgxqzYWzveSLEaPQ5HggcY3AM6fH6cOaM7vF5t2GpUPIoXBrWxjv12wgoGeX
J1y0N/ZBKJDLew9WoNbD+S+ojj5l49/pVBbwJS5OLWYNBH2rormLc2AnmN8tRliD
RCHwPEejytjuUQegPi1L2f1exTvgqHS+/c8zzgY5+inzsCx2BL1MrqGxHnA2nD7m
Dw6O3o6Z/a7WwnP0Sh5K6V1F2USEOibZvf/qCDPdjlyu4t+zwxC7uZrBfnpQBXEv
q0pE1983VFqaX64j340ZTEnElfuhxDhzCnBICp7YINXonuGncfgk+hbvKgNkK2Kt
+dugon5XPoU6UiieR3Tq1FNCEuQNcuaZ6yXbqvkMfiWkGT3zIqx1ZAPODCun6nDu
OImQbxStlnbLmh6SvRwlw6U/khSJ9weGTJ1lmULlkV3xOxTdYq2tXcykvOF7X+uZ
I4O5mFhjb5VWK1p+eZCTRecqbagdKM+ZUxtaZ5b0SMNYHEW0PuS0MeBtLmVgyQi2
+W4iu2Vkb5zOyF83RH1mWxH2kCPirqd3OnuuyhGeExOcHF8nC8GL4KoUWXGo7nB6
fCU1VSltuNGy/G0qFQLUi4j2qz2VOXyDchh5aCdhE2M9JXzIzGMch4FIs+ffORA6
3VeO+rVq1bft/zzVG1Ky7bIq+B9mjyT6/hDIkfoKUTZrsEk/QtlOMTIn2am6LkMH
NFDzu1fNvUGZbMjourpQMvhC/ADbp9+3ACpcGXGdfxBBgXu779v70F/S6PEtaZGB
GJZI7s6v1y4KkZ8PxYsJDudK2uluhrHbEyfDwkV7roBeP5fx/mdq4JsbpnCvnIdU
DJfaKLJLwJx57jHNTgUZ5E1FPqd+GsyNyL45RJM0iEDHpjF1a5A7Nu2YsqnVdSWV
j9Np5iyelBqflaCrNFLDVY4iLD11cq1NcNFpXFKLs+EFtUa9HxoQ8s1iiQZUkM9b
Fdy2a4x5V+ChPo4wivXmUy2qeqMfv4Y8Vkh/qjAo49M7b5jjqir0ochRnM10HLkg
DFdJa1GfR5SQxG9BPRSMEBfiry30t+5Rv6DHzEtcKpxhBlAiIDg9iGbATaVH7fmm
E68HCGa61NiY1lWkkqL3+WeIxgclw5eP05A/1wZJIzOF551eR+xv8rHRXKVB29Y2
PFa/B0gTxvEcXN/ZNz0W4uIxMnjc8mhICDjDCs2ns9/FjuxveNIOejpHmwqb68nK
C3H+6yYp3v9gir0o4GoSsZ+81H2cwxnfjUZD+ii4jxj0eCECFYlIdO0LKHLiJzvQ
dk5SrT4K5DMZ13u/9B1mzU9eeIb3y9pJiOr9l/kh3HPyW3vIJJcPqTHD9w6f4AdQ
1uOQbMprwt1eWFJc47e1gZs1H9kn7C4ZWeAi1T57KNCZO4B/V1IBKfNNfkDXOkkv
17Oo9A0EcL8CIUJsadRo7hN0Hm/xHbVt8tHUONI2iJy2LYOzT5Q0kMamiXxoYLLN
u65vuXdLn4P+iW7D6mWDorWiD5vRhBHuj62yFdvtladXWOrZCjZglsU9wE3C4te9
p0ET8WgRBvdB2VRniwC+LAHLD57s2X6uhvfJizNG4zPj/bCSQlJfe0zs7wbdbORD
fGDkeqLYeNokkbVm+QfAXDob1u6cZexfTen1AeBnFLKzNrOl5yA14cvu8NxCpGai
R4eqztUqaM6zP1nYelX0UOlSEsTFyHZYgovQGWsfvouEYDEdsWYAjf2tgtM3qxKd
0TgQKQeRLqSFGQcN3yA3RXf7BBr6xQGEgj2iklMAq9zDm/xJ2i0TaGWYInTtmAkW
h//JDgyG48FwA2u84yX5EWSKUo4ZY6rVq/YPozTZJLmUQsu6UiKmnSIuxwKBJDB4
joBcK1/kIYFCWTdyActTbKHNC48eDMu2uI8zPu9IjEcnYGcmZMdWkC1WgJP3WaVL
QdTFmOe9Pe1UFg+UOYLAAiQZSZLQV1bMKGI50ohfkbnLJGpD8CfKKUpk6bMlGcIt
X1bCPH/ZVEM6pJPREzwYIpRtL5bzpX4WrxF8c5umFsP8EFan7Fu1CLEtW/PadK6C
0Zs7LXR/IGpeei1pSzu6dkrNx+Blazb8yqDXXvw3/QSqaRio+0aMj+3XiJikvGRm
+k24vPLjEG7s5ZSBMbSmB/cUncdvHd4jKWJXd6Z25Pm71ZLRvaKneg0yv/q3VRKq
vj6F7CFr0CRpMr7NtukT5XNPOuy2SmXBSECGK5XAvXX+CqOx4e2+lAkBF0eYqxbh
ipXuPgqWkGuAmNtj7rbLZtE1a0h2cCq0/DGsE9go9Or1g8o+51s75tnILX1crAUr
mzQJGo71ehJrbGN9dTI8VSLtWVYHJ+5W5UgifBmeLcIs7kTAYBChqLpJTyLEvCtH
2U1lowKauwO+4r1C2iQR6LcUd3lYXgkHZTZZmEF64qsP08jJ4ymKK70ay4FMGdNI
fM8nRbJqf5OdWHxw2pubJj5zyQfH6+CXjOygqhnNrTycnB49wEP2Rai9fKNzI43j
f+IAL9QlqdNnlHoJ+FiuWduJkt2CvrYRfhSWyxQiSHLGcHGivZs/MWnoLzECADW9
8XSe65gW+H1nHaskFflS6rKTYNIXFrIu2WolJYm/kwynceYExL0KXuWX6RPO2f6X
l8qRGltjx7LBgiurTttKBI3VfQGNu4UhpGbYh7hzGyxZMzcsHabCF5JO/7g98aNW
CH5VBOjwvMGB38w89wMPFnL4vZXHM88HnGET6VDt73t+hdiH/kKlVP9o8RXxzQbE
6C/6OdhJ5ZmAsEF/6L5nnORIkzA5EHEoPoGRmZAm7lD4VPiD40MA+QAXySWr2+R0
zuxcC5msUfULhtkI34jhXK5pjT5Bn+tCEJR40rXSU7rm5fvka8uNmsaJWzyzibTC
Dsnu9X79ezGII2Qnqic+uLZIW2t6usQJCA65qxkRspATfXVGcBLS7aZcZPkfeaKI
Q63cQ/Da1h7P3lvw7wWkUIZpSkJ/8Vu5a1wFbnQZNiZU8Y6Bejgag+sO/FxYSJW+
yw/ufvZYh90hama5XF97IuiucDMK8gvZ5jaQafMMk/aYBbTT2IPkAVCJCPpEE+Qa
f9Jp9oIEDxBEVa4L6fZH5Ce6NyRiJb+gmTL9R+sTXXOJnQsVCaMKlDDRk74xLA8s
lTsav0u6LRfR942Q5p5i+yQcDiZXRmJBaWUSHXyaGqzIdgOcyiR3FK8YkrnPx2ae
PUWth15OGeCtFMvMUu4gLsuv2g83vjFLtKm/zZfdrMGaA8/Tj039OV+/MwNYU1dB
oATzyco5Zfn18sEcmnF0IXwSH4M8NYNqcMTIV33P5NW/miCECov3QYJVHF7ZPd7J
bXElLMcs5MF+gufCyEdSgOuSvTfEBn0MpmYf9bCZsgtllEAXfmoPpb8woHSS3Njp
ljUgWjQUe2jcFWMLJ1h+Tw9agpggOs6AzybWAy4rOPt9kAKxNpmRVrU8m1SbTb1/
Sta5oN3cKyCyg13zKb9L/uu354O4l4ZwKtZcsL+6f4eOu96aBxq5e/l+9fB2OOPC
dN18wPPlMclXBp8NdioRI121dFUPXs3CrlIhDNPhWtf3qT5CGuzCh7TEeiybGoxS
HXsIR1CqrcwVziegarrsvapBdKR5CMiALH8c73Ijnnd/penwaqJ0bWWCIg4C28RM
xpzsaLtWYlSDONqV4IKE+NTjQqNDrQifGZtxzBPVTWjvZjdIlu3QvxKTajR+Izdz
qtYGYlK2kf5lD4ujIT5g/z8dMM1ITLw+IotyGQQu8ZpjWPOjpBD23k2Mx0qAdOuq
PMv0sGLvsUzNBk3IQ/aw+eby0ebEdWdEolM7KuMdhuqphPRVFNRdNC2WszCl+Sg7
LkIKcMr5D3u7R+buwWuKJ0/avCPyWeC1gxqVIkk9mHSX45396Vpryc5VrS0/Ffle
jbOiahfg1YPJkUxX0XVpR4XEAP1+Mrw/FqyZiTsG1ZPomIrEFBQiHnZMqPqwu8BM
Enub39CWaKzyvnjidyuqwKXmGx/C2d6UQzZ+HirMnqPZTCTtwwNbMqCp9mzyVSGS
ZL+09BMpy2gXDb+E00Pz48NT83saQieS8cnWoB0xDNrRwacRdFbz+2SpxfOsl6h2
rFr7tk9P8e9l/XRhW2H2QINXXcHlgx8kkgsOOrluvGsrIljNYwpJt5b5WFyoBkRD
dhaG2lGCYxOTiYGe7NC6DPoD11aOhITeVgJlmTMW5mZvetjuOdIYQG/D14MNj9Uy
S0SoTO8Esc/zMd4fYpYObqApYz3g7CvDyVddHiXgQq1+DpNLkBh9d9pcWyj6dbK9
sTD5WGO2w7y0vsdvn1njXFlYPgnClacGfykS1B5M+2CrIhDP8W7wY93EXTwLhV9s
je8Vj+1ZW2tz7Tchk6y1Kqn8T0WIBidVMDyFWtnY/grVRVRutGJmN+S9Xv8bzKSt
AN+LOlehDlah22mgxaIb3XWHjAM1OkrM66AKh4SUSb+stXXs4urfs2+e4svO5j5d
qY5ej/VsbwI9htuevYzZDk0R4cKPQBkGV8PSTukAD0g96jfuB3c0GAYYzyyQsIKJ
jkhMZ5zTjiSGeNLmPIRIyoazUdNYfQ5fl7o2ISIEPX4+na764W3t+w/E4BcqFrJ4
4XkhLAtZ1CUiYelhCh+ic8i2NHfflz9/3oJxprRYEmG7S0N/I0We2bRMBIJ+fnzE
UeZgKtiJ3swSQ2OlJ3VbmjfjQnmIZ4Vkf7vutrkUIWcm9W7fp48lzbRaOKGMdIHS
qcXu6OkKtLYZH8LCGgdbK9gEIPVON0Ok6dHxwcVNu+vdJqtpaig/5QCLvbFnhuFw
65NvuvDPaCIcUQndCp3IuTPNOiEFCsLqxOsUy12mXan+VLaJpIdGrehsgYE1qXx0
L3YXcspaxCV+e80Z8TYhS0HsG4AH6dif301RPLP+3slkd85aWSIl9WrbewDaZCXu
KLvtCC7WeDj5DdA5hwuVec8snbZNNmeHc4Nt+xmpDcP6ze9BJN9dgB18sjG6mXW+
w0YfeHpm1c5rA/G8v/+2HAYhABlUYcbm+9wEgYgrx8uP1HIzQTa8YU1HZq8c1UzE
T/lX4x+FdMcLv4LChBmxa5Xe+77bzP1C1XU8c0mERYNVquYKKpyiybgXeepG0qNE
r10uCMD+62M6Q44Gc0mtMKnWO28yTHQoTnAZ2b35ZFBgJy/c/xyvbU6NDbhN8Xmh
NQQt13KsMxN2A7nmeyQhuGQTRWvBSZP3vrGf5/4uPYVtq2TiZYUlWO4DWAnxkeFL
6CSVIoPKCUQiTtO+tl3Igh0bb7Mub0OQKIN9vEweF3Bl8UI2p1eR23l+duaPplzB
N3fC+Cg/V45tX38ImVD5TQanWMFJIY5z7orgA5lKfQdpkz0OD2pOekyZtlv+z0zP
HNMPG7Dm8Grl2hGGSJTrfVEL4OYOuG/xGxbQmBuvm0TU0rftHgeDsoYcf12/wLQM
7XEm5WYpmBniW2M5camra54k1Yf/lQ0sDE2thyybkMs1AxU8Bpr3usO/0ahv1BSQ
sqah75kfzOV6/dTFGqn+1cNVLWdVmFLpEAbX+IW9q323MiOd9sBTZw8gYBAdCU3G
ENiU6R4BXkSaeZNg8IpZL4UQtaQMbYVoE5JWJ4qpzggouaFndhZn5hi1wY3LJXi2
v3zIC6eCf9SKbo6tvwdJiuV5v9o+DoKixPBduv7HTyCNr3vxM1YKwXdBOzj92dyP
566la6bG3bvl+Pz5qk5jnRe6Wq9UqyaItOLAxtnnUHu9o23q41eWftRp0FUULySq
RD5j6D2UMcLKLAJ/3TxYIyPOJrljyJ+uNkvKuYLYGT/80JUwoLlR/rCeDAUlK+Rh
G+5t8ExjS9TiSr5+fkBhXZJapmm5AIcjG3GqsO9sc1HHqK0+rBRMK6NOGYnZJb/m
KvuymvFGOQP1P1fYioYzG+XmkcdgdzAC98RwMJD7h3J6KkCAPiImTbQTMQzUksfN
gE3r+56w46pXr8rXmXSupNZnu0LwP8SIC+9f/qZruS9I0Zv2YfzqTDrPhjPigTms
3y6u06XxQVIJCEYmpzNh/qEw8Nyrm9ATK1BNaUm8/pucNdFvejUahe3zLwQ9A5J9
ELgpkQSE2r6Jz2SpStb+/0mOcC3h6E2h0Y/qa9SZB4Ouz+OgQPTVFJhcc23KFxKb
epk/oUjqR17+XzFjuR8sRtOJwqgHW2/wmU6d5AYOWOxASS5nUi6YCQxwrcS+Jj5G
tWgfKN/oMLhnjH/1v0i6B0fPasCSloff5eMnAiKDUh6WMhLDYsLV0c2MC+NvziaW
6EznxMndj7xqVR/VoB+ui3OjZ7QJSArmUn2+M6sOg30ZUBr+gq8x6f4sPFYIjKJY
zM2FTZSRoUzbIhXCKiBZ/KGwD6Yl3DUYpRCJs5628JEuNhtwwdy0K6Pmu8HA8QSP
zAEBFgzoS9T3QU61BDoOgkinyV3gYtdlq8cfueyJittsBeA+lGKe1EIyFv3vLLxS
swdapySFN+OQIoLZM54sgx1GEb0Ai7A/o1mebesrYZKGSEdgRhGmapYkIv6I2CyH
lLGwxVWXYlZ4H+U9J8EbTTONGUXB1y7eUez3zB61vTnklYYkhNaoxmBdiR2A1gO4
FyE17RVK3Ls15GTwNdMGs+J6Xo/qFz1yNYzKZPgxHHDECBJHT5xXQl5gVjbkktCf
+4+bvdwluyrb0NcUxt/LftL0+To6zqFWoCKLJmLRmdZHfrq5oZk/LlLqDy3KLWLr
fCOWfiMdLv8UtYb8Rjaw+Dbty3Nlwrh+Rcfilwf1xpdZer4oKSp1lftlwSJKW11W
6YRUg2dXOr44gugKnYEdhpCZ9vjTmZ8JQaYhpryny5ykaZUr8VYReh7r8XZHyU4J
7by0MIOq6dlxn4OFYI1dfMXWZKeTHnVl5e16KJrvo5yY9jHK0ri5UIgMC52Q20PH
UWnBSk5jx1x15AQCe8R2/3hZLJaIPJEkJGxOejPSNO2G+ZsaCPP/dKvdyaqYcp5e
MpBnzAEQ5ICT3YTmjEUQvsk7Xusxd1fHXC+gpwuSWNZievSf24vTI/8sX/zutESF
Inlds8ANSyihyIQf7mYQakhKcjb9RKXWJUzffjb+b9s+GAmyeObWCyfwQxS1X3En
aXS0Ynje2m8qasbFvlLq2R1srM7H1B7XT2OgeOWvCgIeTm1Fn8i3IJCbKTC8kG4x
LbG6OGvT+LdscYEWIMv18jn75U10VY8kVk+w+ELXVQ3pQZ2Unns/vBO+N0CZeNwc
Z+VjLUf/dVqZCBbwJJ3MykgWIEEil+VM7ellxkgSXpTqiEwm0aTMV4V/jVEsdHLW
Th/CXfTJQ1QZYiXo0ZJxaAb/tDdu/qoE7i+cca1UdQ95aWxaGY9eoEkv0eq7Wi19
elVPspLhlwsRiXQw1wmP7BM7C3ycS7cDerV0CYpLn9Dg4IWCBLhn1Z56UhuRTL8K
atnYfHCMj2Jxs45FmAfcK3bZixZjMbFbhyIRu+L12wVSkGxRKIYLl8dXYpghdDE8
2etrSR6x/GHHzlPnUZPUkZBOBDEwP2sZ/Q63VstP8IioJz37DcrtluLl+4nuUqad
/ueCwmcOOtmL8A0c+WfbcOEIyRlrdOXCeF5ePkbN+8OhI+pFTo3YKyQdIsQG7792
lqHCnlT1GvbLuxI9ImuC+avyPZ451sZWWpZQXV7kr0kudiqteskQcdK1QCEhp85R
eStq7w31jFaIpQ439ey/tsGikIKKCIEXK3WrCSnn+FiZtoUtr7tD1uSLuTZecBFG
JKEsChgBTy7Cbd4CTcuDA1kON1UCvN9rtriMuu8hVzZrc5XojVMIXjTWYEkWPEBD
1IVGAaWd/SnB0snVypE3XVztB46JPqLHlCurocE/UGx3JmO1fr5V3ddc+meygR9I
JXzINHVCyjpLBnjvG9IXekPXB5DmJJQU1iCdwIEnQFizrbhRomDfHpT5/kVrnKut
XjSZZgEcCXbOylVF2XvtIx6/x1O+DBYqmvZkU5K9x/eVbcDkcEa6EIKdLtynAIwI
D8RBMFYiTf9qOUT4iDcVcjrpVlv2tZZc7YDL8TbNTsfjvzJAaYfiKd/PjaErHULa
8ZthARYqlPqHJsos6YHtF39kwkA751+bhlIRGhpiZVpNQjWW+Rneui7RaPjmLcdO
NJZEPYnyXWkbooq19BnDVNQu6TCxEt2h/TfP8q+9UPZPGw/DhJFP2ORyveP+8AfP
4cu/AYnZJh7RIex6o5wgQBsvZYOD3g8YxY/0qQsJbJqQAprFXSGHqNDsCaP6O07t
392hFS99JQEvdnHs71xa1P1Uhy5gNrCCRtLAp8wIkandPV72VFq3BSXtPsiWIxgt
C/bo/oDp/dbk5cT3zEzgsns43jnH3DttDHQrzmqQMWBmb4cVsM7Ce0kaK122zyzC
pSVfXdQXaqo2Wg5cOzmg1uYAEMMxG7g0BgOHlsoL1VzjJuN635QiJtVMfz52qw0d
iD5HUoJZzOy8uU1QX8jtQ7Y1+364KU/qfRVilPaFh4IXwDnRCcXsb7pnqGwdR9X2
QC8D9r9WGzP4mX0WbjpxJUjaa4qdHOjjpZYiSv/nAidzFq4PYcEDkOFc/nYKBUNb
hY+hT/u/PphG0atLwR92+PvVCW7GrDM9kM0C+q0x90C9+SOaRRPieXnW5G5OmbjA
IQudAEMZM9aCvenmPkPzoTHYz9fAuyp0TvYVJ7PU29+UyhVfPjNSy6h6DLSuAFo8
dVb/5af7xGPQPdrgwoauvY0UpIxkImprhnfrDxzLK+taLDdRs/O1Z0N+e7hgFNHg
t7qCTupo7av5xhMuhVeGM+o6EY/ZN7KrLKsjyOf3UgoIYQ3YJkASrRNdv+Yg0bwf
Mqh9GEDsCNjtudhw18ozMLOKUqlRm1YwpY55kaRBzR8azXnzGHPdrHIG3/GW9Q9u
vvPa9Zy8sKONlWzRx22d8Q8gzyPjzcVU9EjEK7zhuMQpuBziZyXD7hpdBOxcHvoa
XIT2k8L5og59HKDTfWqVEVaqAOIwM6RJMNQW6WvpP/Tm705LGHD7iyCSRuB4r3P5
nw9+KqhArnnwo9ALDtZiJHmz1eAHdI9IS6qsPp9a1mRPYGGmqjTzw0ZPyt97dSEC
LG6/fZ9JxD9OgBhPlTAUA0Ald5IZ2b3pfh1dacF4spL+N75oyhjq0PXx5t1R4Ra6
PgG4YKxnX6aSnb1VcXIbIrKCZHxlO2eZt9UKogoeJrsx08FsriMoDVmvE9Qp3hxI
3vmtQvo1tZufSGRSM7UPk3wJ/XAeNqLNIFpcMO3QoA9ibfloSM0wYZWVyoFkaXiU
XoZzg54H9nDKJge0k4e58CEu+5k7P/yfDfgNkjztkwTS/cetumeTfN0VJz9uqSke
rSEZz3mRpXtXf9NMRQeHcgFomNSRHFdCw8T9I46EkfOV4eoJQQ+ppK9CTjbwtXJp
XZ+lHCWmjb8my89HFFNYgibTsqc0XCPvGfdQNxMYHWLkSDQxat9saZEPLe+/mKTt
a/alDIyOE0jQPfaplWMM2kWIETBSaXCtNMRKSxrJYXT6rFtqVDMIJDhjIvw5RbD1
Lde2Elc2Iu0IcWwC1/2SaQLH7vS/SDvXv19U6gDPddpsxVha9TbSLN6q4U03RbZz
hJqgFMgNBGV3Q4jrikzjYuzoOJQX9vZQuZIBRpJNnhINgrpjhM2esnWUs5dgJclB
fwMAH4VLnJ+mvSkLBnB5eRIquZvVqcc7i+cQ84I5LtgE5naOv/vZDYm/tHpjyxcO
0m+MQqSdqevWfo01/na329rsZ6pSymE4HIJnzzSzA8ER+n6rJCsqFdUqRDCoqgEI
WJnltdzaSHF/WxYQZ1R7RLYwUlKqO9p4sH3fXstOKo5apUpViI/ORZAJ9slnLW+2
nkZA2vQj41AfC+yV1TFlXAgeLnvNyR2HjACdPSPEQMLPbHowbycSxS4hsCVMXHoW
x53AKjsOoSCeF9be3PgdJf7GBZ33sQkQsouW9V5Cvvftxl1f2Q66LujmAsU9p1by
a4uSVNMRDDGV8gm9w5RD1kPw5cJUU2sTg3CSJU6OtlGk7Xd3ngQqg6LKpFI8faUX
+IGEswNomAwmNxw1r8drwTPtGgU6OT/YWj6REwE8UHbu90gR17gCveALcCmG+oIx
zxddu/ciR2X1p12/vc4nKZkjDSG9zFHXsv4UfMag1/OpsZNSvKwvSlLVt/txd0l3
kkVkky10ia7UCfHgdEyu2d8tZrC5Py6iV0E/Zhqg/JgOas16mSN7kVns9+Livwne
3MezoDSVKtr6upEzytRraXi0RSHP02Y7Vcd2p02PUaqcpuYI7zuqqh8nO5QB/1LM
aAglRXazJxKqQvsWH97+j77BDkkngbI7uGL0S9LhCoj9eyEAux9OytdF25lahWFw
tK4T5OGrzegr5El865qfkdKYUNevBCerTfHkfY+v+vMTq+ruhBpPMiAltEW26tvu
Dc4mNFVfo5Uy86cVrThGkIeJWTdEvCkQggQ9fNSFc2OJPwNxLQKuiS/9mShydo7V
1DL1/yJgYOcaUo1RfJjcLRZ8mfBW4W9KiiYMcBZkVIPMohyiZtAbwfOTXXlYuJ82
z88UeQo0Ech52TY2u0WtkXeRUObOUXsmPOm1il3PqdNnXU7HRvMAlfZ0PJwPPpfb
6VU0lQJCyhdrQ2u1rE3q9CuoHiN8XaFmaf9xI4Z5yBzhMTqP+k+pxk2hPhXbEgLd
EoXz/caYM34OoTm4IZvBJrtyjG2yBM9sstZfDfBo+4SuMJ8aR9QedU0cQF3LAiIQ
cU0dgotx4LDO9PGWni92Jd++QkPp8/H1bFnKc2XOkmI2RRbhcGgkq7omlQUVdiJN
Y6QK0hUK30bIz8T4ZCo3pDaRmH/z0qfssffzbAFRNRLN7YDnCAx4kqY4zWOACk91
6QuanPMYgdTk8KzdkfiGn05KzjGM6bD4ORbNa8jaVg+2rUdTbUV5m9RJbXrMrdXX
8pGSugujj6G0CsKYsPSaVAAZNOOt5i5DioLWwLdh54tWQiTCqgnDEtlnGlQyjBYI
5XlU1ulL3Km28UWeODqYxODBQuhsyMgW2SI1RlJZ8c7eZ1XgltHU14kWsbZtK0+Q
BI92MsBQioNckVNqxKjXPAz1t5Qlh6gXkfSCkHXYxkfdlD+WRpf1svS685GKuumu
kfFuY+svzMCJ5EOKlifk58gWVTz00B1qfxGRtw41Myx1VB/jzH+WfcGtbF5y3D+A
1pulzJ2dVSLKtPe+LlQvuHqng5EjsOL9i27Q6TbKNFRV0iPDspF81MlpJ7ruUD4m
Lyd6NwDlSoOKBv0dBTI7tvizvB3aVkWcvh1ercx5+JtUOYvFbILRxJq7IY9imfqi
XxTjzCJ6y/UltDUt6/S1NyDR9MWDkQaRhMQ4q33PMC8pCs2lrmztXWbXt1X2/DNq
crnT0FDJg84Zf+SssE73YZJG6ejAUSQACVRs0iv0CoK5Z60n+w+2/p1G2eR0+raj
BYsIpsc244/MQmhn7oWZFNGsq2uNPGgres69UIX/w//qKfGrtRdQ+JHNBZxOiu+O
jgFx2igWqtuK/4vuRY5qeMvVA/ACzIMlfqmYNb6dVvXdHGs6/zPnG/1BhJXBnSyu
R4UU29Ln55rJfEmqrvH+jGfgG3gR+kwTzPEiHWHaQySj90x3k4Y5SgSk6d0+/pAE
hsMyqn9q4ubVCdxzJdJ/75xnt2AQUythpmS6Nc3a7IZobXDsi1oohwhdEK2MD2Bq
ppTn0Z3i2I0JcoSKzY1FFp59RQkFgIdluhWJ8Jttpl+tIfroR9xERpQGvm4YbOgs
0uAYKpOlKz8J7f02gDlMSpeGoE6gpS7gcwIOnYLbKwMQYBvCls77fQEqiribtHzr
s8M2tlvvRK6+c0fB0OhSdPrOLHISdy8a8vA2Pf2KSqZL/lidsrBRANRXMBvUj4pC
9yq3cyBVzRdW9VIgc1n+LQNJC4ASKwooXrO4aKeqe6xXuBJNijQO27rdgv8bX4d8
+cNn3UtNTnIn6MdeWXQha7OGc5hgtNmc3tg/GscBMoTWafCHAlGNUne14LFoXWiX
xiwcacnVmatadOHuQSvERIL6eJy6PNTEEeoha4QEzzSOYiR0SCLERTLtF2EmItOg
RamfVD+BDs7Y6VKwNWvswEvoiKSuQYXOHpxhuOq3+aWtjHeLOz95IBG+wEzziyGb
hwkpdhC11+wg/k2yY0Pxcl9IAQzumAfUTNZqk1uB4UMY7PmC17oDCEoUFiOm7dtn
XK1A3b19l73vviB6yi+apdxGc9Llbuo2mG5UQ1NnBGN6H1TQCmTsmopRktL+jjyr
USDJ2q7zcmC3Alx71eGCVaYUwsMeX5u4T472KcUbqQ5VujjlpJ98PFGDR1EOq3an
r5r7hNyM6cyr1H4/nb+5DjcLRgT3teZUlOX2SOcVJ5iWgLIm8NRw0g5rmB+kwKMx
hvvs4KQY91XY3XiptyJf529ZNwGmgyI6XD0EsDZuWDPbXL1fLkB3tc3l+3ApdHMT
oCFdBiZBSOtaM3di/K/C+5nwEnW3EqBv3NbVbQK1xCK2pit3yPOoeTN+hThnqfza
Tv9QOKOVdymzlM3V9kMKmkuK1ES6C4apxAneoO3yT7N9E5qQ57gYx9DRzX0YetOM
l9eDthww93hbXbhseYZJj0ItoPjUvol1qHkIgoko/7KXgQBbkW1M+JbT6uGh+Gt5
SbQrh0pQJXmh23A/3NEs+hw3WlzS5Hw5Gybh3qkYDb6eBVZxYukZhhTw5kx3oRPx
UgH0U+3IqGtGnAx4XjFFIiqyqNEzexUJETKTM+YX7aaVkKny3l+nRvZvB7VJZteK
P2732AfrDOo9s76upKdKhwlBPafDqYzIfJPrDMCBUXOjZWniFCRBCZlH95kiumk0
FbIa+NMbGzq4fGw/g6YLZVVVxEPGyy7xtg7blEz6uFWAZ0y0kpcsrtDwbggMOfIs
NqgS5oGehj8/gBSAMwxZz1vvMV8xSXYteyQia6JN6+PXlZa/pyeHSXwVGWUPLJh7
Aznwf6CElth7chg4brOMzQi4ZTsB/Zdjy1U7kq8n2ECgSW9A3FYtdMnxd8Z+rN/I
8l5mZGQJRr1AKJaEXuIl1ZOAqc6d6xIjn860wbYJaE5p6e4Il2V21TareHU3q9M1
t6k3++vm+j+9FVTHqSsAGVsKvUZ46TW7mSdy7gzBJ0HAeGJTjRM+4l5gP9VBhOc3
s/oN8cJ8EPZn//C8pbwzQiIU/yHE3FCwhkXYkzPusD3MeDGjOEOr8XP7i7AvsBY7
lXL0FQ+PlPaXbEgEPbdAqGLClBsTRWyXPMy/uyi0+o7zG9MSz1iK79c4CBmtM1f2
g9trWGv5gs0/fVzIKB9vJTgiTrMEfsTStnFC5uo+71aU7iL8d/4h06RdjU/E52Xd
GLe0SqD1NQfVbAPeYJ5GkTxsAhX2t2TNlxTdxVU3NK8cEtHa/YQyo5fhIg+p2exe
8Uzqu/SCFjIuJPrOuY/v8wY4Az+mOLj0suzUDB40ZcbCnSfJj6aO2SYl93wqRQ7Q
BkHYE/NMkQ3CWKngJUfb7gokbjM+zFucZtyKE4VnhdrilgxRIo8WBstNco0EFfjc
jo5jexYi8PD9pnDaz5yRbiF9an/l9oYDhuDDhDxraukDpSqDCiD2XkDIgMZM5juO
QGmdG/dmo3Auud0WOZ+eUkRDtaaVj0VovZ9Yoju7bx5/lNT/oKpxB18V1NZU6hLQ
eyTwEd8enhuJ4pTmeQFDwMfOvDo7hg9qtlWHz7Uzeg9wR+WBR0E7NxYinLLCcxyu
MuUwuoXmJEwB4R7i40YJyHDP+K9LMxytp2xAuV0k6R5Xuq7P/LftGolIblXIhuFp
/Rh7VXD+cRDWlisOAAsi4YM4CVA05eedmJg78UV2kTIfyOKdzK+p13HKmB6aLGdK
C9I96EJUBnTBESfNcMTH1dvZzRm5gtTTZZHNTyL0DQNbiPuw5iXm//Kf6PUqio3a
S96UxKrweXl7hfXhMNnf09vxFaaRnYX04GJVTvVotz+JotP/m85mzqUi1pnRZD4N
X3d24slBDkl6hNP/RmWLQxBJ1ZI7OjBtdf4ld7I8xALgh1fYzDyYX8rdvWNZuf1G
sF/fsGZE+5Q2FGb17Btn9HP7etOCGLU9c8E/gsyrfaQuRWrFsmMHAmESHx5/nI3g
9B9SKIXTNnXxLAUA1Pqds8uuywFcLOzbqwES0XdtSxCXnaHOOVHOlp/CrisfsHvT
1y2gHlaQgFK3P+hGFGDI1iQ4bsjOShYFHDzNdz4bFwW2DlaL4KDzzSEoayVFXZ0O
hbpd7nfQzlNxOe2PWhB74XWqNmflyUap5bbCCOICymiUoJAi1+aD089Ew51gftBK
8NUEF6rmBT62KPHWEtHQaipfLlyFO0nkQuU27KXj149zohbPHbSIarH0Bj9V/8EG
yLqNDe6uOtlcyh4UCPf7O1zbof+N7KKS8PYfckpC3WQIw15+hW1fDqL2zI2jGiVt
JZwkc9aWXLYnP1akbvCFuOMGBFNwkFB0QENzqS7mVdwDtDwJemlDhU4oA6eEpuDD
LzxOofagF4XNNem0Aw2j9ROxp0DTQ17Vj5ux/9vQMAE54xSPU6cT/H0UaYqSE9j5
7uMbyCdmJvqBc3GDv414+r/npNYkKAKU2KZ5b6+TE4orVoABg4AKfqPZ99v/GCpH
YJd1FvdPaCkDINnImPhvIDZAnF0x6upBS6ZHBbw0z1u0gPAuCd+8m+Sf/wD7Ads4
o0dN8m7geDCtLJ0e2duDTOATzxvJrH8PqDt57bT0/UsC1kV4ENuBa6U+Gb3Xau2b
MnVYv5QfTuHqGrINdZKBAHH+8h088+zxMbV5m/6ScDy1oU3datysnkFBe0MAgz60
9cRfh0qBeoWY07qshCvHggSofdbbNbweaCuYYWeM50stFpw3lKC9KB4JwmvcXef+
UsoYJsU74+ke7CxCGQD8H1Kwn8nrcH0E4zGOLoYvm/03VB42elfPNby3F59/Uxnf
64uXQlo/79lzTH2dfsV0KsYanOsyN+2X3Z9xkeC9tAXF1rnTXAW3KjAqt4qNuFXY
eMEtbgwUsTQWMfJUMKGPYSvBI7sOsNL6t1voGUEc1KjY8T5++bTibYXIyodJI/hU
XTRXZRyvYIYUHotrLbrQETsjEwfrAq90K0RbvlRA5SznNXSkRKQikOm7REPY102i
m+lk1DieTdl3a+lwTKY4hNYV2dIqobh2WXChWMiiGhIVpLVEJ+zL3/JWUnVavuOg
rchzznKHNxM5WAUhtQ+dWDQOzATwJtEWybycizBmVe4eQPKMJJRG6fG1tzwfOCas
CdL7hj7WXE53mQ5c5HN29vS7a/4Bi6VxzgX2Bu5SRRdxyPMkUtE3kJFXDgcgwmJt
KWoZRmPW5RXMa19S8knElUM2PPsaCzSsfRdoS7Pcs+7Q5ghUaJ+uNaT3aMEbU6Rt
FT8oZ6GBvBYC7z1IHaHQ12qeRUbh5Xxua+UjkF4D2HTkXJgMmpR3OB1w9rZ5V1yW
8Vw0D1HAvAQmhzCJ6RmFuZNHcB/eDYxa5/NbRjE1Y01VnCFIecLWpUPzs6o3bHN6
ijO2bK4/8fHnpDtBaPHEFhWZJTbvsAoD/tOsgGt7k+KObHgArhroHgrTThw82y79
UICfZsRyIqFqk43BQoyD7mK0qsMW6c1VL55Aor5F1124bjIsvk1YRY7F7nKrvedt
9ILNtEkJazeQa7KdrICFjYbNrO9rb718/ceSwTK8sFsaA3/u8IAUwCLYgE7VOfmq
DjdlYSFJW3yrZPGyVMEL2SA0E2MRZq717X4TQb1aWXVkvJ/NNOkCXmxCn0VGOQtw
vMYhWzAQ3Aqocjn/XLIdnGYhtfuUCKrZiP+08KslSW75NT8R77puNb04Sln0xbaO
rYXAmHRxjTVeqXOZovroLFlTxUn7pltMI71OrKQPe4Xd9yO9PTRYyBGHpk9nssbd
9lHe2fFYLzIb/tONC46plNsk3vyrrgLNjdi0peN3H+d1B2Utf/5Rt5aDCNPx6s2U
byzQYld3Nzj/SEgNMKTiMBpa3nsPq6KjLCA/RztSbQ977sjaK9azYcYEh+tA2uAe
10qQEVPekk7+LQQPG5f9ZRkk6Il6LDpx6Rm26h76RlqH6Igd+TwiseI74ZG2NP2E
ZzKkcXLw26jB+qPpdhVz4ORDU7B88sXaulf2Y0gNLSsQGiaNvKwOoBQaZ97xEZV+
/OkpORDV2v5q/otn6/RuhNpYlz32nBCiO4eaouFqYey9FNDnP0nGoNXUkDT0hwEA
R1434Z9+jfTeFPQ7WjBq8Q+GHl3ykKPUVhP18qsqu4oglQKpP/kRoBhbX1XJdbgq
BNdO8Nl+VkG9aWC6MTSMv/EifAKIDeejM4zyRUicISqpt77W2Wfs3sova2Y5u+VE
V3dcSGAl3H518c0eDkOgAvVE5LAZqb6A5B3vMVue2X/AqPrkhn7ZtCI16x/SE4r5
/yPVQNxVY5D0YI3aW5OiB7QAtLgeYsNP7z1Gj/bSUKCCB63yIbme+BiK2nH3tbFQ
Yav+1XzSqCi/scdEBqIkRNFCyqQf39F7nOdH58kKOkZ6tGuW+64nlpQofSEipUDI
SVawEwDyFIe6JgfY8D4jja98DrlYzipi8oFlRNSZNY2RTM0mie6tOl2y+B4ISeDD
zdxCBqFMBBdmgBNZR3sluJh/1F64ATIZXyPKmGSIbbGQpccDwzgocHv2UoojeeR8
ZO/ciY6tKA4BBP7zubWvdtaOEOIZc8ehir1lR+02sDXntFfJV9Hvr+l5q9MErvWt
ZwuMkiWig6ROm1tCtS8utN6MrUiSQ7dEAgBklYkqC5rpJ3PR0dOKOV7Xjq8y9Oy/
GVuwqjTcaerE11m8AhITEk3jazf8Cip0oRNnOJQRxromkrZvaHKZEIgKkp7+ZjlG
8DA9DoLVsnSs80QWAD84tVaS8nt140ki/ETmJD4jrHUhZ/SIysAlviA+HS09Ipp1
DeNb1/aj+iz73hTzH5RGAKuP1TSbeYE+kJ922vo1jJm5fPFdrYq8NBL0JRsKxlcF
K5vs6RucnTlwfFfQKHoQRTouQ1cf9F96+9gSvBoZFjNIeubcWSiS2w+a6xqSccs6
LfPHI8DgXXu6XQ40s9fjlWbiI0fhVZS/BfXZm+KxnM/c2Nij1az1fkveYw8z3RqN
598H1lg+3qtX4HOBqVVLRni8LfSV07Fw4d3l8mBZP2ixoT7uM1i1AK2f0ySSC2ey
juO5BJElb9TUGJoc7OHRoJq9s+QKEXlxTqHXq/4NGeuwSKzKqcOf8GwiDmb1o8/4
26IsysXFB22wRYGcDOY4b8VXo2SfdpkrhQY8i2iqsW6B3RyRlu3s0/2r4kILFILs
Y9aoRc6Xefb44qNWudsHn0vg+IjwQ5p2V57GHDpo6+vJVCaWhGYlWU2Iyh/amBWh
SI33U5ds/OpGWjgK5cQzZaa02w/z6i9dVS13vulvmUDjP/w5qiaMXcOL4zlkMbbq
0pMGUt3CqvJWeSQiCRdNT1LWBKAS4QhheHze3xxyCXEUgdZdTQAaCCkYD6u/eraP
3ddQuP8KaEzJBXrTyEIU+n+0B6E1eBRfrmiJhIMbLtKh0bw0A1qyeghB7VJff7Y8
LFWEeduNGUN1kEVxGXR/ljXSJsorPKBqnEjnwKT6CpE8HRdB8OwPEjkzSUGQcuZ1
yKDnhmSCGtF+X1dMxENSZHfu8LkBtZ4GG14VYTm3vcO1ivPGLwATK1z6Wb/UhNMP
kzDbwR3AVbUL6O3cstsg+eozX2hax/sRmWM1iSjXA/i6T5I8OtQj2Fra8rnAlatW
1MV5niwD+gejm9c1ZUBAuoSg+m94Ggoc2zI/VeRmXShMDOvNO497CZBT6xeMgIBC
+/VO9gYXHJ27c4JqRiYxFe+/sNDitubkCrA4YLAtUiYq12Rd5VyS+VJt/qT08Els
KSlxSqTX9DLQg22jxceMYGaqe0lBjdJqbArWb+8E5k7EOixMcKvw6smrRbNLgeUr
krxOFQgvpj8dxc+JXF2vfsEcbt0A3Uk15rzHYQG/K3crm3qDMZ4PwHSykHfiPOOI
Nssy5u23cG95ayYbzC87GQFSXzMcy2GFlsuqnAsCp/PNQUum097+JlRKNOqHOOiq
SoZigoso4L4atNBq7s4uePsSDEOeQXmgcQjhhcO2+OTY23yFpgW3x6UCLzUorqkv
qJwWDACQ684SSBba2vwfmDu0d6H56FIJuWccV7Un/TsLEXazwbX+znrsGs1LCesz
KeqyVxdnNU/ubx1LRmtUl34+tq2Z0Qq9emWuRG6qxT245wFV2PaeELro7DpdW2dm
0mLMZ3Dm/4BPMskzZp+a/BVnlfvYG4eY1lj/gXr2OrFpXHb+1VNV/SUm83zpih3m
IJlD+/KCqjNKBlPTaAIMhg2R3fm6Q+qHbTf3CWC/7atq5fnv+KWGoUS+t+xz7Sr1
YArAvvpfjhqxtbLKMdL3zkTuE91H1vCkZ+8iywzo6dk83Mz0nycNSlPfT2cizq2S
HAcpPSv/8YRb2MuA0GI1LwcGobRVC8pQStc1134tgUCC/EKECMiV2hXOvj0K+elg
VKVznHjcQ8MlLrc37p2Hf7o2pHPuc0/5dBZ1qCOfLtWPFRJ51zzcc8WwnSDPc1N1
0mJgQYtzESwrTdCP9VuQ9TE3da1cKEolvl/aN+vAe5hig8ZyXLbkVAToFq2i+rIZ
2ZtwEezsmqu8Z6Nw3zzGA8/WD9sIfEfNO76D1QC05zOlEpDv3x7F+MEdzw49M4wE
aCnxeOArPB3EOVwn5IIZUUupaiSk691SRYYqQ8DlM6sd32OCoiiEe7kAbsp0+ctN
4i0uAHJw8HN7ZZgX8dq0OERKPFr6NTUHDHApu/D4tX2xFBnil5+YqP/858Nx8nEV
3MT0UQ8te0AGlY2wu23BEYxIWz3nKL7ZuSR+VemyLA7vnBrUp8Lp3cMhzg7I+X3S
u1ywDCx9DYQAkAZfPNIBQ75KHJXhjt+YXfbvmWg/HR9WmVBExQWAANefETkDhF4h
8Z5CD0WNdOfb0rrLRVueUZFOZfcJcWMrvK8sEEiifNdAGOb0cdtZrjjjp/wK//eI
EokWAbcxByvmqlS36M1RujjCxfuQcrhYPKvZWtd9HX/avHAu6z5uFfLifYNls6RI
y5xiqW4a6ROBZ+HRMXDkb2B0yqu2NqjQ8Vj9lIXkLSIg2pv6p0Wjl9VggLLHo7J2
FGo8n4+fVBo1V9pKsFb/qjT0ZxE5rjwvVDvnj0I2WJj4vCMIu2VfI2X5J6Ld0zlw
jAhutBfu7ZXkNXhVRA+lUqNYpPcnw/h5WYZ82gkZyti0TkQiTKpz7yywTXLz6vIp
AhQoOzaOR3pj2ZdLICbVIdd3Lj6JX8aq0eP0BkyjVqLAEvyDq/c4lIYTLQmXBGzh
gcGR8U4ujT4rsmhBHn4PRo7xFgIpZRagmsPSw6y2NW9IUS6SqXfOxuw74AmaOQRG
7Q+0j9NwnBi+DiOy8G6f/ijvQf0io+yhq9CbGhqZ96OdyIw7iWhTDeK4MkKkG8s2
gezF7VReRjf9k3T04Qp1XCJyBXilo7hYCea79tdRO1DMwyKZxrdt76MFYB20dVxw
zEwpCQ6BzE/w7pEUgs1CqsuRz+nRMmPWw+xpUF2duGPqSjqHTxnJIqwbb3uo9vSb
XT7Llf3mpJXbeB6lWiEqxmXrIl1o5Q70C3wJ1++nUKvb7ghDy/rAFs7Wdhk+5YmK
A7PAP29TaQpvCRgiuEcGANhd2uqAbI2+Se8GkfezxvcbCl0saot97khUIMkQntGz
3l7eJm9OyNEKEPhipwBgFUpfsQlQjjjWIaZSBUXJCz6rlINhS0tU2uHqiJKxOdhQ
6kiydgJJDKa92HFAWSDedU9lsqQfWYAlrMHZwkesutNHw3Zp08FFHtxNoh7lMpYN
3FsAdAHSmY0DVkCfYes8GCE0KMQG9aU6vr9yCyEHjEHxuVLisg0TVoii9TSi4Czz
XPCnkuGeBFuOFUn3fQgxwL+1E2nnDzStFd0Ubm/ByJrPTmElRs6N/mk/DyuLACJh
UQU3qywILzfmMnsFwekr3OtCydDBJZvspqIuQsV5Eim/x/LTtqJbmh1KOqCWAeL6
qd2yCoDxT7BwTTGv0WekaLZ+ksEdg9SSGswA51fatuqXTV+0rfeyhssSs506aJZa
1ZkHACy3571jpKvM16z0udTxnStM9v8wolGGcWwiQ5rSIPV6y53apZoQNLAIDWN5
AhwDKvMrkRuf+AwWR+smmaYK5ebQdsk+67XtwgeWCcOXfV4hogbgfy1jNOxgy+Kh
Ole5L0kZ7VFilwy0pKmhp27L+h/G4RWgdxNjYTSMPo52rRIsD1M0f8O8MU1lkwWc
QpepvR87EafrR0JikcplzI/vtPWXdEoBJVXfjNfo0zlzAvzllk/u/RjAHvaFq3yu
f+4XY8bp3QoyfwO8XX6vcEwtVl0EtIcQ19ZwkQbyuIOYGDejtlp9Y99akD2o01uc
m4o4kxmN1SCyTgGICznja10oty/uR7+3yjFb0rZs5dQxqBZmQR0RS/L7a/lZDKF+
MrL/q97muYqrrUCynyI/YKAgGy/gS1UUEXDk4A3s4Gdds+8UwBajwHaqOq5lcDFH
SwTnOD3LMnsfzUDJkELsXwnDqjZVfEhYf9ILzuWROT4i9+A39h8b/opHDH4TUlBM
rLajs2D2QXirbP/74F8FVdvQWAFJ6o4e868gzwcEA+MivUk2+wyTSa9ysFZsLV46
FX0vO9idbvi16iyQVBXX/4iwvxWtVEH13+X8rp6iHJzxmb9vOeLmd/i1KKFmntqD
SXGNsPd7gfTawONOKyaCJkaffh+ZfYFDT/Pv3Nody7nNLlj6szXH+0gZrK33f4z5
BdJwjiCsL6+bfs8ECU5KvmPpkRoRQNQGyjDhyPtYbNsXRg9jrMrwqC+WA5fT1Emy
btUwNxmh/sCPoGv0y7f2it1oz0eWT6qNpI4aWml5Q7+a8Y4w00am9Wo5lkpE7+VM
YmApyyy6JLQr9jeuAoFa7uRvlrCESHRbaqKTEJYLafccD6I7Vl6ju2zCAlNzZ/f7
SVps0EzWh3eqTFtGnFBiUM6tH4lixF7b23RLsVFdS8XEpQ0f5n6ocyRwWMu9HQlS
kS1u/CPv5axHSXfxySDuvvP0DMK0sMXdVmx9vRq+0Mmb+i/DZ+6VDTIUi9aicDMY
gi+bnanYGMtUT4PrXTDpy5xSzYAnXWi05jzKi58uc37gjYzis5P0jjt/N3dw7qvt
kgG/BhcjlmK2cFJaVpHyoRCKEe1F9RN5nsDasmUI0yT2Iu+DijEgR43T7G6HUkRi
Mj86YltwUvAK2N7C157MOGefe3Qb3F4PtpRtq6eJvG612d5IAnV6+ukTQpM+6cUp
Z0As9sVUK1sJUzGXKJ02NN1plCfc/I7cajejA94BVnVeewsELPKl6JS8fzDhM7Hj
7vkTcC5acs1dryw26zJVv1hFz38cuXA5W3pWwXivCqT0R4bX06SS3XcHlvn0JkGy
DonH/5I5bYR5z651u6baGjhanvGXFXzPy28DM3/AzpjQ3y0U5+b/+qv44xXRMdc/
dv67gPGiQsugsuCBvmcR7cBAJAe+fAYlew48kKUHR7XsbI7nK1u8xQTVbjisyco2
UXszU5I8rQhhmoTViwW7ZXUKJK9pzXuorMnCxPx8yPbu3zZ5QpPybZRDDrLZb6j5
CdqtNYoieVXe2eI/iJ8XRv5YYKsNfkWGBfNTKbIBlUOt5HmKq5N8udwksPu/ejnB
0i2BvstxJ9BQ5zogmq2AzlTJtNqOHPKSUPLieKvay4O7W1so1BcR6GflXq16GJWi
dAdWzeF4i8nJrOjvk3FqfS7gjrsU1AOg/K0150JPG8JnKEAKz9uxp+eXZEaE+/FA
xljjT7Vkv6dsZeUzOOG6AdKUdpH7TrEKXlwqdq8tJei78r6N5f3K53XF9FmZMhAa
qZWOYw5QhBY0+IEhFAsOidmBmxgR6jyE4CfM5eNstDuMRG+Yt/2F0cuAtkmhKmVy
085Q7MSvkubXmmMK8Hmlt/gxa8/t3HRniG7T6crBT2+76lH/j6LyaZrtLMpjQnro
0ullSmNldqGsUCTZ3b5GJFszrFQuNRP3D7lQPGQRm3RYkbVvO+nnOnv1ceYGO2B0
JXYyDGxxMAa9XUwhmraRi+QERVJIL7dN0X/74+Lxe2hOqyf6y0z/UqwtLnKpCQsg
hGmzcQOf2Lxc3sdfsINiaYAFloJJz/IXwz3DVY92NRD2lbuzuQLSN8642AkVu7OT
i1d2oDfeeQAtKA2bV2R34dSi/+oM6WjUOpT2RtEtRD58ztlPvDVIjPNvS7jSLK8D
HRaZnltY72ggE1qTsmaQasZKeZIp4xM+ULCmEmG4nAMzljXbG8rCakqNg8rRzIzT
0gw9HR4QtuUIfUIp9IULSrFhPdPHl3l6FPN35YuQkelAZ+4R+D5dwoKU7pzv1bbf
gMWLGQwQ9/vBR/79vZ4VITrCBGH4kUWeXK5nfN/Zs/f8EThnR6DeGgc50RhJWYHA
U6fBEdP87xhUIzzPmwW2e4Bpztn3DCz4ADzP1yjGEMjNRvredDcI5j5+rmwNO4md
2A+GywLS4UhgCMR6DPtcw+nMKfBrqJEDMtb90mSEV3HdlBpDOayY+i2M3s/m07Rz
cyk/uQIXSlWCVl45e58zBG1nGBq3ut+2255FLt/4D0ifdQJnXD7Ap/sQZTlyJkQj
M29LqO8kvyAjs51MVkW5NV9SeOQzfZt0BnAzIK0AUzaJ0f7xDRU4InvYLUlOUwaT
XgR+yRXaoRYY4BNvEqx9DkxCtm2muTEQPRtw8+X48HwoIpEWToC1UxsOiPb6S+Lr
hS3FJP53dCU4usyduB/U2bKMjwIaoL3CPWWae5XKV0gKbKmDUTsuEIrovcG/cRXj
/KmvKTxUQ4T4+/gWwxus8Gd4yUDi76UnnruHZlkkJ25jJ1ejJGctOrfIzYaHZHpM
pvImqFizFjck5Qzw2UthHn6sBMIMPgarnWHSz2gXUJyB6moLm2zUPfceNNONuB2s
2xtjbtozXPmAVTQg/aNBjn1AKOcRbxADtITpYlyp6ohmITfYKVGSgJalH1Ov0YCW
+yqcrSWrEZwfF70slkc9WjM1hMMgh6irXpiG7Vb91EwE8tvJVPzBsdiuePi+03qY
f9l6nQ7YEezrzXrf2tSKTfoLt4vsZGNlWxJcSKh2E/83tCnOfAwQ7cYMURwsYVUa
SibzXsqUhvbKUaOkFHLptdNONMFunLyuvfHJhPVBZChBlY8wQrATOaBsBdztF1pn
lGxNFXP+VaJ49Ph9Q2XFnDvXLvvxuOhDbm1cfwa2yMVYi3nyNoxn6fIoM/UAV/jI
KCc9pWejLBn/r0kQbYjrIovG9LmMy4VHt3JBtGLrGDPhmJyPIuMlbZm/KzB7f+fU
GHkzq/YoOyxnc9wsZVdhEj2UDqQG0YvFUMq9tqmjgk17avNu/+9lDxYojU3cjBQQ
xx7ETgwzRCFfi+J5ivjIF/wA7QxMowZY3K5kTV0Yz5SeSkpV/R2hUaqSkJhqXvEq
dc7a6mr1lLaqu87ojA2HLD2XGI0nln24XpR51wtt8tgJ6RlClFYgNSwweDTK8BEM
N+gDLy8Xu6+oIYPJwWddjCNNjj01fKLj5sYGlY7MXEkHq/agSev85K4fqKmrxF0X
fdprJA8rnyDc5nFbTDTYJjMPXPwu4CyFWrG2Dgd+VROBPawJDYbiqaucwkohdGWS
XIDCYXADOBm9MjfT/bAXlJubn1AFQmx29SJCzATzp0OGrBkhYwJTW5vMbX0tlo8p
s6cyDgG0GGPXPj+DEsthET0Wvwd0rwgNAjQu4oimosNjXwbE5Pr2YRtVrBx/UyZ5
Kzq1tLtN/XELSbpM8viWYfevT15IN6T8aSSOtL4MMzW8HCYyv7ZTa5c5YuRCfG3s
DTrcBR+SVpkw96/nyuKP6Bjh0uLjciKlQO5Y4g0JTiq1TtcweHJkwrXGMTPjp3UX
t8vzfX4nUeZwO7cxgr7zkHYbyNnfsSIZtgH7VxP44INP2jClQVBMwvNRMXv102c+
rSPfJDncR0FWjfF+76g8/1G19hnesLfJWIp8gazVXNhb/xucvvBsbzGRrv3rGbje
XJHbk4aDSkoKXODBRfk8QTubqfB4eavbopk4HeKFclMb8HDkklSl9oyM+cJGX04X
/mUqj9rIAJ/NILS91mQCEu8hRU6dcUGFcYJ1CFmFoh+MWzzq4CqtxePLAGRuVM5t
qAOREqAH7SSKeipgThXK1W7hppG7jgyfoVj0d0aap3SKq8PR79E1kvp0+r3rzyCH
PPwDint/lv4SSeOtyUK++qBYqpT6BsLhaFsv4YWiqCxe4SyfxFD2PdnLmRA9mkPP
2NgfltOxYgIoa+GKT/yR8CJ9qyw/Fl36Kxf00Z500pMqXE4uLBIM9/oaVfic5SBj
EJk7P8fb8BSMdNaXAv+Nrg0qRPuIdfKkgrDvE6QDoPXcKLWPZrdqDwLJw94sKf8e
E5WpRyoB9DJFWSzh0jv0RocLb0ElU0h/xSbPYtuF0pnNWegoBQCU+MGdhGrNavIb
5ifhQtnzjDHqOQcBnrzYQrU64cR4G0HWmKfI8LKn2bGxhV2OPGVxORBSUP480oHd
wi+xjOfRkZuocpvZlrHae1KH3syrihU4PfbBRNsBFf6dDYquq4+owLMZV1Em5ltK
9ZW1O3v6R1Yi7aIXfM2hIFIHuEEljBdDQKTv9BeXj9WG0NBbfuYHB80Tl1Awogx7
2Ep4iLznNa0J7C4FoeXx7+kedS1OLOiggOVeqFmkL16Z8bQ0AOc5uNadgccSOhEV
CdsyyCIW6ok6Whk6BejBZlfPMYNOSiwlaVJs5386JZ0ERsPTWB6dhU9ZIMpmKPzR
fdA+Bc9JzsNrXOTGqJDc3kOgFEJzvjIC6CR7ZRt4rFJpE3a7ad10M8CFDVcqG9zG
o2aVz3UZKUkLkPLqVuAJlsTIYhpkZtWn9r1UssNGCbMqm0nKMB4E6vwNYwys12NT
x7PEOXr6Sop5cASQ4A8YzfPID1S67IoGbbM5UttOGtk0aON5zl8dKmc+M5gmU/um
4EUYr03WvJPAtrNA/nq+KIJwSS1zxonWzHkBRfgn1ff6qAZ5X/MKCrxRkM36cnOx
Smc1eFkR1g8mKatBL7jRMKpqhSpxl2dVCe64Mn+Zf0Q5oLMl/YZIMqjgNfJd+31k
M5yftD4UlOwuFvq88ZIDZTfQCRmyfCImz3+R8HEUmCSU51raMyfxGXwo7JpfkNs6
spL9lIckaPsa1HTcumzdsVgghx2n9p8+FV6/SBq7iNkgCSUNyo8wvK1FTL4PQE6j
4lVOV8CtTTLInhVjQyg2FZFCw1D5U2ChqY/SI9SOrmGXoUw1+xCVxv6hRnvIFQxd
Ae0ki2nmu/hmAIGcncGQxoXp6/QXF9D64hB2kEdBFpxIJv6PUtfnY97Ee5uErkun
+4TTWQIe6FlmIWS2CvkJBE/VSwjSMQuZVlB64V63BYSKyszO25yWOZ/Xn0VdBXoo
hYo6pglwuG+fRP4/M4KMnvzBY8EJuux5qBbHe8nvTgmaH4w3Bp4+t93kf5stZSa+
fyBR65T0xpIWsG5Q+BeIUqtkRGa0utUulqKD+mrwOIcYBwvyt6Qk042Xa0ixJcSd
bJyt2sZlnceqXMoClJNHlQska8wQCyDXHpGLvXnaqdQ6AREFGnP8/ONyNWBPsBwu
4zqEZduxuObl67U2o6DeG0iv1bAh9sFL/8ZgVUd1zunskBxqssXrm/TuY4+BpDFM
MLNHo1zuL5ubEVcU1rjjiTirbso3Yh91/h85KaGTFA6OdJQUgr/Mt75Ueq+qLiQy
fTs73FwJq8fzm2GbuEvZjrsWbKqAB4o46d9cVrVejVJgnYSgLGPMGlSMNT48EaPi
oYjnNynP0wrQVI+pikD5h28919woijTd3M51HSNbS/dRMkS+n27MbfgYq3/y7UQE
gqcFxANTlpAtVAQVqSCaKzhI2zvSTKoTtkg1zHyjoTCQpnPokGkkS0hbJDCep+a4
ZSyWfJZIxVj3utS0dPoQ1fjKu+7T4w8QgxHnYH8jMLOuLGJ206i4WLQylXqJtPOS
Tb0yRM9QKL226ZRa2oG+LHcJ3r/vp5deeutN/AqSRWj9/pC2+aG53Xv5d100dWsw
kjF+hKbD54oXSqBBQEmm/yJStCYtaRlHlRU3K8IIW58K8Qf1kmTwfnOfrbu9dqa5
oMlM+i4be26Lwdx8A8y0PEgAKLMzzOD3jy6CJ7IPSvPegPj6P5AhE3snEra7dtKs
HH9WLyVP0LlO1Y2Gh5XkigV0cwAtkfqZvP7uMUnj6jBbMdwnHY0YuY2ty3lGUM8+
jVfZdb//UepdODAImptCHjEOwQm3mDqHMb0xzWMpI/8xQjgt79pQVZv7DWndJVk4
9LNlGMkNoO2O9688S2pLLO9scr0LP2rRgfH8XWeVpuWmLOs76neSQV6gRbkstJjr
861z5DesO+7EX4bI0cd8j/U1XTGSKiF8ADyeFzXn8EQcuHMjeVX9VRo8vidzUk1W
SqBfZ+nPUUrd1cIzW4r/jSuSQ7y+RAoZYQDIuMVqWHuBf4o1aK8si4GelW8aQ0FY
9LefIPSdOkilVwtv1/3xlxFmmghsEM897okJov5JlxbqXp1FvAvd3hGrqnT/MdNp
FkHm3LYEqoi4s2Gr8xIC0JbtpjWSCnk10NPQFScH8I6y6G9R1IRIrZ4t6JtHc0P2
n1W0nwTMlDIZyLr4atTa6K91GexppdFffJ/Wd2qnQk3j6Bg4PFtueljT46Z73kCf
s8cl+ksjGR8hIQNhHllo5eeUsYF8rd3mR9z6MaZZDRek1iG5GvarH5j857ujcskb
3Syw62UAQsbNn0JAK9qQnLMKLP1h5peNigdPDYuqukcp7OpOAwdVJKA8xb4NWdX7
nsDo656aOc1X4hLhj/pimLjCl66NxJi4WfhOZLDIBzBRqlWS0l0REBujrhsYvwom
wrAVRWsCJ8luwfEa0Bf8LVyH138hN4JFdyKsbdPVGiFWPhQkBGVvZkYJasMIOEu7
xNlhgU19ujNz0uwQ87SGSJeUf5IkiDBGr4WtoaW8MA1l16Jmpz950AMhPh63MHmz
QoXz5tWIgYlg5YEk/i1jrCMUhja9d2eEv+b/txaZ/jLxVgGvlI2D9llcDbe2UJMR
2UtWs288Fwf079bi62yNw1F/yyB3Oa1hk7o5WmZTnuiv/Mccp6BY6M2zKCKpn/3S
TiUmoWJDnHfqT7w82rquYKGOymVi4irhMKN06Ip/e6E2oYcgHJfhEXbygRe523Py
SnpJp2vsoPMN1rYff/qgc4Ki+2BoUizBUijjoT2nspqnGgTMkKTF6ZPFBo1/yg7o
czn+khWkJK/a1sMRWk8FCGT95/zZtmO/XUkYTbsDIFa336NKOB21FV6mJ8DEpmqR
XFdFq5AViKANRLfif15q5/a7KEIKx/gXy85+OhvAqLo7KVp9oN7Tsj8qeumhF4uX
CqZPGD7BTrOYkbhNakWvpOWNFz7KS3ob06I8LqNhGRTjRn/l8vndtB/Iweut5FJq
TjynlLAP3Rng1/dYDlfJB2lAwQiOGalokkdvk6K9NyGDnX1tGuDbNpaTpV8NoHgk
+Gg4FaQQT3JBTT6TrXpd8J4NT7zcasrE34xgcm7MdjpyveagPYzo2XdYV7FTGvRX
scbkhP8V3DQFmrsLn/wRC/jqbp3GlXRuFS67Z2jQReeBvOri81gSEuPg3+897EUA
GjiCLPI2LUeR8br55VgcbHjlcSbtMRLvExIoeEh4BKvdnYAMf4n9uVe0YLEiAxPN
U/jwL2lOvcvmq6Atz0XqkYARDEA3NZdgDT6EgLaN51q5MhGikk/snihbVkOx+CNq
GLvDoR4cRvUO1bAgjkpIhW485DFgknJdtCfOWc9E9d3AVLOv3uD4cxXbiEA6aJn5
q26deTyIkysF641XeZGswmx9S+1D6nCQ5B7WoPPB+rWJUts/qCcu5cRUVG77FA0O
b5ZwsBGHCDn72W2Pkln1nT+UkiSB1JTZ45mEaESspFb+z+YM1OhaUM9JwUIY9baR
Uoyn4LnZLf+UXA4K18xb7QQnDOmCYECkz1s8Zg6ZE80kH0ktS7lR3r7dRCA4IWfO
Nnckr2WxSy7qpwm5/B9muhhtma2+/RyvcuBV7jfhlDY/ZpHQOBxiD3uoNoVR56cj
rCNutaHmq0Vaco9lyunqDMXtnLCEv5wvB80ytH5/zRZuYKnQCXDmBHynHh45GJL2
OhOewXI+N/Ccn9vMXW5b+nn7Zof8cTSxyHb0fd+nbq+56NgZrlvh4wHdoDa+r/IJ
6k6bscjGpMvFAazkEWdxart2ASWKoexL6LNGVnm3BeJG1/U7msDZ/I1lBQWS+/kb
yb03EsivygxXz5csFeHCrReNZai7PeohhLWH6vFBPI/glC05L5BG0/C8j3hMRG5Y
ILblG+BAFGzKLzOGzQG/i+wt8Lv2+0Bq/GocxU9mw+gD+Afyn5SpEFZsT31BzB2K
2GTR7rLAefqavD9xNUeZ7kSAJlJP4YICzn1DP4ERkRwLmWWthyrp6v4f2oISw3wJ
fHiu/veHvzIYCI2PjXxXl+UNLZ7txbA610V5yK+pIjjTom6AxpQQs5TonzQjXZC2
y+ZN87RTVi903gC8p5pNglioZG3ouSohshB/Po7M1IzEeFODySEWZHjafjXDG7oi
SskqafTyDbYd9RVnVuYoxQ0Pk336lMTRqwihDTMIR96/h+Qa5+cVtKFf2Yll9ILO
RTY2D8zqeIw4k4ZIyrJDHf1no/aR7nobZL6Y1pHnVHzN6htydr+w08P3iOR/q97k
ydXKSV+JXChXN+HV8L0qBmgU5C2tpwE3wQPsEaCbCYcjVd4H2HJpz7hXM+olGocu
sav5kzQ3qK+sBV9O+bBhzlLBrLZXu0comAEURfozzViXvW1RwVPUsszLx7vhpsfy
iPvmnlhDKcQkbu1i7gTlRg3CEjHx6pxAIs3D47jXV4JnJdgOlqkSkNTNoY14diLC
2Xj2snBGEnpenYZY/ZfK7GO0aUs9D2oQZ1oIKrmyOJwoHRD634y0+RjKLgTiW3j+
gqZpiZ7V5lhiRI9Hn9O89i3jhrwozXiXyxQJTqRIM7Sm34oL/5ABiLzYb+bUDtjj
rEqx1FH1uXYkGedu/hBTIT2K4K80fpLEZULgVNBHV45Pj8NVw+uVpN9ksuaYT6Db
v7XiGw7apOrkkj5ELDibpv7guqMQwi6+lMxIy+varc2WeVpx5KY4PqDzM0Mdzupx
4xgBRbaPDdB8hVl9jsCoS5EFm3REhEFi37bdcH81KPxTa9ueVNPFHZ/q0/PDLaSn
xZ2AzyqLH8caRhLeJJa0LZ0HjhOO6Ayd7ViKIGuFfVNEvnlWv38eX0nEaBk1wvha
6Ptq7cUyUjbOXl0heq5lzgPXN4Q19vuZzxaAqNq1j7WXHCfKktTkH6HoJC/ukf7m
+hCVdITHaLyOmDGj6vTVQyXWqvH1BTDrVtF245blfIGPVHo4a5ZI/udPKE1vDpjy
T7hnFchfvyGRTsjK1rqkJ2fuKvZqsyd2L74w4h5lBK4vy1rncdcyFs/CD59SW/k4
u8xBJ3vr0OR7gMqFysBKKK3Exz2k7l3pbnhp5xOsgT2ofU61hTvnK6a3Hgyh5UUW
w462VEulym+RoR6MadgLFdTwdZqZCiQ1mWnYOl6D9RHANCQZWVGz3tVA80NjpOIn
32PU+hf306A6KU1xTYFpndWyZ5zxWcjvyQ9DcXcPjZeJcwxc1v2uzIddIlQKC3W5
x98YC26N9nbRuNyhwE87Spgzf+wGajKz58XQ/CbSNCwQ1OSNTV8KWWTB1d9IzeUt
uy1HYk35EVom5NGltoCir4e6ed16AUiq9nGWJeex9tdG/vC+VYe+rIAVl+fsJf3V
cG1DL0eR8STHudd5xOiI7w9KlGIj28aiB0BVdScvtsuPEzN++LEfgUmPb2IU7NdN
mHJ5ifT/O9AUkIHeuJO4uGTF5XOp82WvnNYYkZXKe+ISW3nRgAR9pUAOWXCbD0T9
SXATEYhuAphmgi2PjtJbYDzh6hQeIHv6eLeIVJjcxE35Pio7mLsef+L20kzUMmBW
hh3vwLjWmeRJzsIsNbDVLJ0ucwZyRvIrs0Uly/LLj7Asf36kf4VQtaQ2mbnpyetB
ZEA7ppU1uhRSL8k1lvfL9j0crlzI/MKij27l+rxfat/9Y4osQecHpekcAiYdT5k8
fQpT4nwx6NHMlkuLkBhX9RJLwH/mk+0MNekhkfmgxZ6CU7PCukAKJC73R+TCkwBA
fpH1LMvy1UFCh7TiitSdNtuez4/xlc0C65yd2imgrAcv4UHeUBVo7U2JImaX4NRG
sck6WDocqORDENzBkK+W/MVE1Uvsp0rNyQ8wyXhQtK7TV/kRWZKSoFQBXyJKjVpz
0E20VMZaqi9eAWnWSwCsSh/zBUvAGJTqiGCgbrvg5BvuPZqgz82FJ7eXcOYGxZAV
XdS9TGoaFHIkzrKmEHQZ87wXl8a/+Ribt4VJ26EVguNEf6GXZt9XID/hIbBZYW5D
MIWsMbUlDbgRhl9q8pCYQJqlLwr7BqzyyMwJvr7Jii04Ruj2s+7CNF3HA8UiheZh
/LoZQgvHXt2E4lA51ROeQ8QQzmFD1Nke99QrsO4FuWM35NAWJLZLdwbiq/cFUQCS
4c9PcmmMca8WB8DEyJ/WGJ3QG000BSmemSfLODc8LT4ShpsRjq268vt4E7mByQAZ
LmUVG5ZjaI86NQFn6OC3m8zkBljwR891hNebVkbijz5vLyh6faPtVpHDhicr+mYC
Kli0DsGqNPwiBKQbawycruR7ytAH6+fEJnDMW7Ic1lpYKulL4NuXKaSqOv1IbS4B
tKckf27KUppyC6X1BZzaG+dJTNybofmkfeeWcrLq4prCjxpmY0BnRFS25Dhww56S
WN6Czbrs+RG7uGao3CaYSWY9xSJT6wJjStyf2+ZxL55/xTQWO71nljaBHXg8gks8
5MUkie34lFUDkznFoQhLUFPOqaDtt1c3suF5YnycB49Z4R5NjJSl6nSpwNoFJkH+
dhJ195Bt3DwXG0FhP3EhiAWbG3d2lWA/hshn8Ve+u4JbhCls0HYl1J9YtR/VlZh9
SZxDSnYbo7p2En8UAlB2XaSZtR07KjkLtvEXLlYYQSlxEbA7eAr8/4D5PNoDWEQ9
9Q9Qw9nxWxu0nyJITcIEbv5mVuPRnS7tnwprOmXcNnvAJ3chUxQZiocaa4J6E7BG
6chU7YwCqTRkF6b3w81Wl9GXmVn+bPvken8IPK9xo9bsYH5dS9PIDe/jLi44xuto
W+qww75UBkmvQOvhsR0yJVkIf/IJGuwyu1NP3H+ZxxpoxIEkIIctQ0Rv0Vi+S2h2
1TFJ4vIjQrtvG/ArHnX57ofJ6FUVGakfD2KWZCgbOx0KQyjf//VzU4Iyciy2nprK
2+fujUwytOrFpMokSnDLvkBUky341TvpGjTbL5JpIpaMF9SnmujMGvzVcfyBHMJl
BCat6+7gKRo9ZqAoYnu7oq+PzGFFqIqYWeGc2YCmHVP39QY1BamJDt6WXM8XAA8q
u0AF9WUgyKXG7TfxWfZnvfCx6KppE56ggdLLGkUHD+xi7me/yy4VtL7x6iFGt55y
RAXWNERXVXb1VyR7yRTp/1ykX+yY+M1kCmOX2uKI0lOc35cs0yY6I/5o+ZLrq7Ng
A6iGBLaQ7eTw8xNKexOTlvl2hPKQmkTbE6CDkLl9TSKXGE/7wlWA35cM5KV9Uyfu
ngD5k24jx2FiiO7TlRdrPg/pcS5RRBtzQ2+v+tK0keI1CF4qd0scXSCgDzkAlNqJ
DisOINad2/E8mOe+ZyVluVII6Oju8f7rmf3QaZ2YO0EmstxIVgeKzWUE5LvPIEM4
lJqnqLvFlQkzzPVdHfMrhwdQOg1ud7PVKUM8rVkUlwvzI2XYBg7jpj6CrgYKoUAY
iQCFudGEzVpqLcHEug9a7vxKHSDtBtEaR4Huat4wNTLE3zV/x+FyWf1ehQaYICS7
vaqMgutQDxSfkoQ8gkSLAOL4pngNWLT53oe0SVUaCDyzGj0Ec+864OIupFjNjk9T
5vwXUdqo5zQcbx+UqBvXKBNDvsUJIfFdhWwNd9q/lv/395fCURouB3bruzigNzyV
h4bQEkJGNfbPBSOU23F8ZlTRYMVNdYdQKLx0kKOsR6n3isioPtM9biy+J/pmVfaR
SnMKQ5aAOxafuCgmS+BbxM8o6JW4sgV32UxERkQ/1DkW10RAir5CRd+TK7lwy5pj
+bWRPKVerHdBjJ+vvJ6QWbjEorFlDGPtLaZb7xbYKnVWUwRr3qEXxKNl9XbrUiLu
2qRPuWtZ4QU570eR85qWARHtS5vXWGzPNWJ7RatqJUxEYDBT7pHtYnBmin6tW1Ey
n6qRFZl6D0zkPJ7Ryh0d7YgYZeAkXcmgaLObZkbUnvlt987nnOk5uWMQsDxn8eda
qvtXWpLNeM/6ZZ2c4zExU3YT+7KL0asD3HPcHHMdN7QP8N9XkliyFI6Lh3DQW8Pn
31yOE6XVOYbtOV24rOwmm+lWsUsph3mxg3qknRNnZqc1cLloQcyC4Jxbr/er7NvI
ZHIe98YwWQwvaxERGjnx1LSEio9j19EbUuOmnav9SyVCzY1ue1mvcUReVU6EzzQX
R/TkvdLU1A1fJmdX7a8EFrzy6l8pej4SKlBlrU/LtGUAE7ZVPQETlTDUuiqDbjw+
8Z93PK6ZdY9AVV4ZQidSXWznxTkhN3oAzzIh9GhzdGaFPiQkDlNKOk0mtGPCHJci
7fLwHinRMIk6eRyF5CktaN2sVe/8wrA2hULoYmHYbvVwQ/iMMMNlv6uEu2DJdx8y
VgFMw/ZymONshcWa4smEMDuSk65qn7+2tzPLhEyBCoKAZqCmmMdyRk1xGmpbG/F5
rwpyYPOtXnd6n1qpurFnkSgwWBlHbmo2qU1OcMnd/rCDrj/LKyC7fWwHnQ3KBa41
med2t9lBX3BfN9PGBrbKPocdMPF+mWs3PNhB6/LKm9JM0a+im6QXwsBYfzuxywEh
6AWP3HtnCCHzQb3C3tJixVFK4GoUaODV7axZJBBTApfUMmIN3FchYoxXZVaDSvmJ
DlMVIDfAwtmHO5IQN9ZbYvVq46/HeLcePWArh1quV0auEZsoxpxAVgtwRt/LMRFM
q2deCSZ4njW/hDQVdlbmHTrFA8xAd2kLVZ5VRvZCuqby4rYan6GLkAg4iYkRjOdI
RQ8IKZOP+eFORx3FEWJ1J1oP2qKhulHm0Cxsq6H2sgbOiR7Du9f5pJCQH59zDSAB
YrwmURnYqvg5bkyhcYw8uuGWH5XsaCgggR5Em07Nnln80rloOjw7yjItCHfBDkNV
SXfK0HvArU5rv3p02As6ox0aVx3ruxk+JoEGbt/QZ/D2ZqxUsA8jDStwAvE8wvDu
FoakSpG9Wk6WMPJO/nYWFU3G+tjvhYUoboj1VALwRbCLSL8t44qA28J3UjuoHN2X
VDeet5ewBN0XBr08iUgZUcvUcZT4PTSGsvM7Tmb1sRluTAsdp0eQJciV0k2ytPhh
rowGEewK4cy1nepOI1a7Q9CJR9fZuM6XNrEd/ST6x6xh/wwOZ84pebFAN9jAETLE
BnQu90oMx9BICzYgRfUGXXoWOkBUk0Bf2k8z24JhP1vtj9U7ZbjEMOU+fRlg7s2m
cvsqEwfU/Eprw9zYdiCUofW+9UoUYvOAv8VpIiUK2BOylrJdAXpSf+3JSzqhglZm
HdSerss0IdroF320SSV+s0ov6awOw20Xtb5/V86b22Br2Bl4RXeqknYAnrCyiYMI
VQd4QaZtQyd+O5SMcvIfhzaaniE+vzLNpOF1gn1XoJFruex+sbTro9c08eVBaH9J
FYm78t+u/7HayOfKrBgWjm4ukFWI7Fc2sqSxxPDoekMqBPEqKCqC5nHYUwH/5gs0
gBNfkW7GnqvLNs9E72vCBSrERlnIBihD09qS3NilUV4pyz5xFE5w0No34B/tit9E
ur2yfr3lLxw33xMZSRsUQtXPD2FJl8qyFUN2NQyvkP4SSM0uUx5mCvW4E1qG/gYc
bECa8pWyfsU3XFGEID4ByC7eIqMSxx0o/WiHLyhheaWA7K3pZqWv8ha4NqHLKV5R
cWmcztpWtxG9Fy+ENQUR6XMZPtapcJlAG27t2US1W2YlJ3smhMtqEWTZFt9/4gRN
C9snJPSdsfzc+Po9T0AoR8vaNLhSGteD7zdBtkiKx/TLaSk89wcYPqveT0Lmf+Ek
y8TUysXhMLX5hXkUSFGYFWfL2ZYxK7JHvoacqFE3C01mLst+Tt3klkgaJ0RkTmWs
GAjw07Xr3s5TDxYSKNAkUqA8m8sTVbQ8PND2T1OFSi78dSasKAM/o1UYGU3935D8
fK1N/Ft4cGPlbXuMAmBhh4ppPcYkBtWxvSR+5n1mMeQV8Xp1iI0I5KixbNLPllBX
kYzTbXSBjFrjecS+0YMSVUin5S4Wz3NdZMvGXC4YgKgWuRQvWgCSqwtbuwk7XhCQ
nz5DdzapvO7Nh2488OpzwU4VCNpTNibqJbgrU/KK67XjJLGkYYZBz2jqajHNOVDh
vpQHV7995frDya1ggqWabCRoIaocA86aZY9/kob5+VKsOOhtINysYrC9KAZ67JAQ
GrgAk4aPRgI58LNle4BeEq3Vl0sINYHWlCNoB0w49Fobdb4BQLUjfZ4oVupjymOz
t4/i+MH3UG5b8xuc0NXpER1MoOeWu/SI+UJ7Z7G0KgBe04juKrUrtQrGJCnaKZrG
P0HLzHOF9wPg9wDfOY3H7fK7CNpi1RdUiFgM8VDsEZO6c/KhIqGDffp6/6QUlSoQ
+HLzBV4G2RR/kRWMWazPYFABMjfphF+mGkNlfd7Fs88ict1mFVas3XzqI50B7oRr
OjJR9kDVn5vP6fqvg1FIUisrHrzfBMBxU1navuZjYMy/fcxUpnLjPX/lRFvx7t/T
umwZNzGUFhDrspoiD19wZbYYFNFbTXINaARffZPVZVgmPMKisNVspocJpuGZ4FyB
MrEviqDVXrGi9uv35pghz06NhffqGEbWRuUR0nRvJsvdCjtvU7r3P7p2HUXU7UsT
pFVxj4h6rEiX2GOwOq3EfwDmOCWzbSrg1Ni2Q/BYWvDenovpa0+PK1Yaz2u6DYiw
1ktS8ZJh6ASVtXZ9ryH0CfUIIyNn4sEbqMhFPRki27BbgeOWG6UtCcG0L7PnE0NW
B4mYDv8ge891YH8ZSstwS1qF0ZlbL/qZF6Az+/yxIoZ5b6L6anyqk0UZNeSboUQn
yQZKShW5GeFWHAz9mSwWH6F3yS7dz0iR/5zdG5g7VmdrEKf1iIOcTzFsz+v6vXAQ
CHyVuq5nFbVrISSt9ruwG2EYORhjE77IeKuPN6Gzo18K0CeN9A8MnDYrG59MRXHL
HyTW6DIH/b12F4WuAe1m1/FkUzKYv3D5OgIcWNed/S5NonEnX1PsQgdZgcZ1yu5j
544o9G+m6XUDDb1h0WCUsnkc1WbLUvIx6WD2Z3kaQwA4+gM6NLqH7f2DwoCBluCl
UBPDxhAXsFreqWI2eU0HM0Lk3wLnoIYVTOsX1L/ia8ys8DE2Cm/mek2Gzdcp05ew
sAr0uzCNQ4NXkrFYciQm+9rHK8ruoOlHZ7TOFTLuI/lHFeG4j0sY106NjrIt0iRM
t3Pmr/Ex3W1g1nfpuo1aT0oIWRo8NnZ7YVV6x00eF3Qb3JSaFuWnuz3Ma/JpE/Ob
lZVLwDA0Vvz75hikYwmk1LkDgDrwRQGqI+2nj1r9IRnCHSzYz/QE/IrIlEa4OSui
3Zo7ik8GZbsfZE2vyCJCXSHfK0ZDtCX2wgtV8SdH2Ub8GwI0RQ2oYntbM3uuTpPe
KHDzN2pE0mH6RcTLj//T8AZ0tG9DvKcrTN4buu6DWQWwFEww/4P3UjxvZKZ6GEe+
2P9mMCtoE9WSMXP53PMUjicl4l/ZO5rrhkLLl18VB/hqrrdvQObv61VxRmoPupWo
Tj1Wm0hIvqpEFRvvO63cxKEs9aXX2SZVwrcauuQ46p/W2CQPlDDzNdbqSQdWxU8r
gIoaTCDbTfXm+JDvkzFqGfx1/JD3WT021NyTetZMqhbjPi5b7OMZwN1w5a6JpEqP
0OgaRgeAS8/dfft0u/FQEydcOJb0jrpA7lw3rAsuk8Fv4M+4Inzig7Nmtqow5u+k
W8T5M154o0Tpxqe2Ycpmvg94gf+VWmmEMf5aWq0yvRQQpkQDGKTy6/Ucccv+kFiB
r5s6j/6htlOq1ddwEWYUHluPDjrf6wNh2Dqcej6xcJ4QFni3GHZ7WjXRHxilPcrM
yffs0Y0FynJmEsdYkt18m77GBtMwId/K3ocVXWrpCEJr6U91FY7lWctS388eQFD7
WE1cKrilc5GvpIxFKo5qSiEPRCQ4Ro/mQW00hOha3K16fDA+c1MK1ZWQmiuxVUo1
F7KRbi7zqmFjGcAcgZkScco0Pua5s5yvFuIxZmHADFABrSw51G1fkqaBh7mjAdTD
tlIz/BQbZq7lPRpP+/a2KH4TijwECerrrDzUaO1q3l3wuHkhY+fXQmrDYBH9cLW8
AK8SGcmaht6wjvlKfeSfdML7MIj47hRIF6jgwD6HR1x5ANFasA01Wqb/y8lLWUxd
eJbOS7cUaU63wA9gjMc52kHZKvG9EgRaW9As4AY9VszGVBpJ5sdfdRkhmCyECrlj
vMOmpmhRtdXgo1be6ekyivBynSUQI+z+BkEho6iqqoQHcrHU6E6tKN+j8pIGRYbt
oBB6hTtUV7rLRlQY3n7FoCQPko7ATVfyikUUntN6mOIaG5NFR16CFqmdoAsIzho9
5ifEby+W6frmvC21NB8JaQGaPF7IBl0E0oDfgZg5ru52ty7ET/T6vXXrd99eXtDn
kS7OuwhllP5bC6XqzywyLvxUcfsAJtvWn0JNXIYmIA9EjpFLWfqcYiCXEhF2pRYm
FDp17KoeeWdKWyD8W7mLMTBRr1jJzM8dzm4kAIXs3/WtIk5JOb70x/gq/Yw9K0xT
dXQvkZLJfgbkpcu4JK+Xk6TV5IyRJ+WhPCUJQoarRceG2wq7Xyl176wQISvHkq4t
M2oI+m59tip1voPom1ecdh+4g43UcDh0aUYU5ueqAvbvJhKwZfGOHOes0iwFLFb8
/7KSzrsO9cdkyDXGROKG53HI+1D/sg3/BN/Kq5VZNefKVAuuupk5TaXd9WEfkDbB
Qp5wmMBYIX5WDRh0YrlvWBw6Ia+SCv5dE3RI+HA38ysJuc9h9yNK5wc766okXAre
TPRggkfBxNrP1o1Lwx3thEosnF7fwJaYeV/uSnn/FzlIqoAyHtXoOoaIMIkp5OZz
rs85D5ZW8XwVpdfrxLx4nmkk/gP/yX/T+G387e81v1eo7Fg/IYRjt2Ip/Ie76Oi0
jL+DwefbmysF9FQw5S1EzoypL/Wh/cYJOCgAQu9euJgcGYC3CvZaXB6r1dWKXRZ1
tCrJyQ0y3vaXKZGBv3h6wGAFvwu/RlejMz1rZikpJpAja2zLVkNBwoQk3YJefB00
niZ2O7bTPXLDmP/puxU68Efwg+KtMpvp8G2395lZvcqaVCTnmAdLpQz0bH86MBwd
5Ym0U8YJRZPHPXN01kUCEywNDqbUxOUSflPn47vPrFtcMvB/tH0CCKnQMSQ9hiaJ
SyDBoEWYuQnIdPcsSCoSQjp7+g6v0+6i3V/BlYX2PO6p7QV8chVKLi+gnOM4nMjk
5uTUGc3ONEEvbUNtDnhD4ZOlDQJu8kXXOfK4xl/YEBv8urYawMkVth5zfMOtCAps
pRAcaOTDaHglxxbcV37+nvx1Z/2N8jl7RMeONWtxX0zLRrl2GrG6vdaD3FgIqRRM
kia2dhX2Ks1tj9prYbxoo/lK6RQBSy29cAXqyEZ49e/K/FzXbakYws1fes2eq7zi
sSxl8jW99NqPLbFiZvihc7sCaefgczlxA+G865CzCyhEiuN8dJEY8Ys8GCSxBtVL
1KHdf13w10pfSQyaUyYBAJfop/6ZDrjVmueLpoEIhr8SNRG0TXfRXN6iTI9KrzdP
YIhI6E/qjV/ynKwz+BBWGMN6DnGrBuFvKZOTSDFNB/tnbgR3fs7OfMtLwJyk+1X/
BvJALFc8anPqhaAK7S6ls3vDwFcpkqUI2l/LclluZmynUzHPWKUwX/pW97cEOQen
WoPDGG3RouKRTFDUrxI44O/K1V1HC44zr1+PM0TRGLUy8H8cQvNJ7LsFRIcuoYUf
sKqqyfSU3sUXEp8Spfrgi7hWL/ecJlnKCjaOfTBies0wGGOHLWYlMFYxR0+4vA2k
t+HlZYYdbT2ODvzPRX8oSTuelKF09cznolt8IjSUk3nmaZiY9PBx7zZ3TfQpKwzc
89j5mGDX/r7Ogya3DrV1Pry5IIbxN7RtofMZma818MioHgSrq1vkhZ1F8yW7fHIj
Gf7+Aj4+kL3J2aEyJExH/Dp99cefFck5vN3HXeRVGJxIURaNNgu21vxOQfrcv9tX
1qGLmwrHnf4ZPeh+1VhNF6AHAnA5e6yJpntdNqC3tBL4p4wObbDtrkRtLta8N1tO
oi7gzf9XZCXeh4dBDf3RE9rp+FMMih0jAHYaAGP2vCCqh3UO2Z8WUdvbNH+SkP+X
I6B3XGGKF6qlEBzkfE7sKSMTbiKKg5pSWGDmFledeeUxcqhxctclIAWBsbESz1c+
6ClcVTl9UugBROoIz2fyfVRZ9ppboeeR81hq43+BQ0O4cy1Z/QP7m+aKbAtTw2Df
aelPjCVq0VEGl5mXJoSaoPB2zXw9OZ3RJOd7CwQJAgjVtgcDBHdDZPzv8jTgXJa1
Hmu4a3XIAlty7fcTnmTHlmIuVf0yhjcjss0A+evEyskSWofk8jKqA9ZyBXns6NUh
NqsdsuJkxAUOX0FasXJJa179NTRDbYgowIkLrZoIrMtzD/3md6kYUu/62O4nyzcD
dSBmdmhq5rZrEi5t03EHDR2ItiXa52mf5Y8Ixdh6AkVGnNPHOB9YjBpaMWBnSQPS
m7pQb8f1ozfGndS0YdSlgdzVP4K5656m7LibaMlzT8OSexNmcxJsIz98WnmaCL5n
KGFmSiWElDvxmHpVjqh6fAnenC2jlK40azpF32TaULuOyEujKqo3SGOYGoODzaxI
OYP0Au8b3n4fcNU7RwuLgmCogpFx6RnkZz6tIYSb+SRvVVESR2iArb1r3g1XhFkE
8nTxbpS/xdLhJe5NuJD3CVcSsDp+Z0UB4hstH1LlainqOq2+U//t6l0yOyFBGxUJ
X7lge7drB+fBwcMPZX9eV+RoIrm2Emi2ml877lm8r3XzozSQnAQwlx4C8VFLSzNU
Etpmqui30AQAdLapq9z+LPF1GCtXdJPxPGyh5aeBBH5Itl2cd5O9qlJc8I5+El8G
TPM+VKbjIMeWVvncizDUjasIFOcKTt5MoW/3fouhoZph31GjcsUR88tSmnqp8mTD
WF/os2igrX7mCJTiS6/pn5sdqJVhVLWcX1FRx+EsDTnJMx7cyR6UcK44k8ERSPl5
bQRB/BhN67PFUKsefCknFFtrELAD6qLTejIdJUoy3Oz3043AcK3f5MRmz/egV0Wd
h7qoRISP4UOkCi5pjm6w8HKawQXpf5OlHejckHIv6BcGUZlVK/peOB+1Xo079CpN
hqdXgs9uTboXbtJCkV5ozW0D+vpPJUpVHfJbcVTAnjiiBagSk6yOsHYIF4ZtYPxT
DhC0WJnYL0A8XTpNrMM8Uu7rAwEtYk5Pm/Xm0TaqyT0TnKyCn0BTge06+JDkMEru
LyxaCNnC6f8WKTDeezZ1iqiUvtLNXPHVVriEuWDDL0jJW9PrHfbyxLSyOEhgjJQH
siBIEpF6TDPUfhRAFH4d99uH5DIyH5lZXni/mYq7U1VUidzzYNDsr2/Z4LE7kf2F
JAOYhhRG5IgJiTORxb3vHTRopcf9+kjMUUtxSYDygf0YlD7i+NTEMCgMvPbDIyKr
JUqmPH/Agn951w5JdTMl4cHMeLXQgT9lSfPFgBGOWClPgQJrWiJ+GmQYYjMGiK+E
MkBXml5Pe5xTXF0Rpte/ACQp3GTNyoC5o1NEz/zSVnx4qA7jYkqqIt3OnPnp4bde
StVvgRfiQa9K0ntihw5JrxReM62XGEoVGjBm0eyvByaAl0uwKwbyVYzz4TA6yaRv
EIq70TW0i9C5y/AUlXXQd5OU+lKlOcFvKWBCdGCCEX0n8bL/O1L5XjOFccu9ecde
bqBrl35hGg0bBX8JJF7PkMTLWbaAwM46zB35/ufAWUNEGr+GJgTDInWgrx16/4f3
bVCfowzncI/rSN/ksnrmvoulDWWIKxQXbR5/xhtugMFRFg1DWn8lsZu0wWqrH2tX
4qA4e1cnBD3Bl1eqvpg53mwml+F31JSuPuuWHX1TLD2K2jAyxmCNIf3rQGqwkaP3
4CgqRh3NR4xLeLBL/A/qhqSSnEP7sLl6ni38AoXQyLOkxxJfcpvsHhXYbxSEWfku
gWjuAcu9bDQ/2t1eKLthaQ6A+FZ5pEaPo4rcpmbCzCsLFhvZzo0psI5ZQKFnvs4f
JYOG53eBsu2HTGCN5xryoMu6zxTV/tLM9nsQBn4nghJ3+jRhNBPFAwd2xr2rjV6l
wnNtFTK0fpPCkhLzARx0dPAc/OY/vdFInz/642hXTBVH5M686FLBYBpvXHzC/U0x
rPJNuF0BU+xZ3oUGw6+UIHVmfsTSd+jox6v1vekMh8heKsfmcNqooXGaft2DO04M
s1zSA6ZEJxT/wguoPbn61sXR4pYHG9qcK2ohmiV1UJauRDwklueJP8dLk8Ic+Y5s
MCChLE3O46zJjVu2aS6sQiFSpm/1U3VqeYBLFr1znGF08jAAz25niyWhJYgXMybv
G7Vb9W4xYvg57pToUhGBTl+jvlYnnc/oycCSNFSth7jW+KrPykdZ0TVF6H3b5dgi
TUfp4t7T+6ZfLetRWTVGB9phmxIkhWbIExfQvk+ZxZ71oinJ5TbBpoD/qYmWc0vh
ugsbod76Ik5jGRQL9ocQFTDeRnJ0UvHE/dvGRu80utv3n3+7bY6fZC6Jy3/SdHUF
HyI7gjLO7Oirll15xBZcUcgn43mRdGEVLYi1+uAf0uUO0NGFH+Vjl+WZZqBy9Jxk
mDedGG9eNowqrtRIHCYtE8fIhZuKyRXhjobvzFp0zkuUZt8has6Fh5T/aHX81EIR
y5LkMHrG+oYbr6nIqIYvFYuRXtyMo2BPbCPN/Niauz98HjvuTu2AreqhhuvyYusm
ESp2JnY8XxbFMHE6JlaYr8MF3TNAisfxfDgpPrCKOLEhjKt572Xgx9FWgRI4NHR8
/j9mCBHJkZNm4YNkgMPufHXy8L2323FktgZZJc/JsZM9953C2QvEyWckNE5xnk52
F0zUMXp1eT7q73VPzrfCE6TIb7o/EmYHOqFw4KytRlw1mLkIIncXFvyCYWdQjtId
3eqwv5WQvSV9uGftL2/Bg/6eMLeF7+NapCASts7izhIlyUrGLO9YTQNMm8uNbeFf
zHIU0mWxBOoqjW3pG8OU7sSdV/WY2pIwT6AWKgDoBhEGqasO4AMIkEZC/zYtBy2x
lKOFmxwijrnpRGtiMFjPLtAZeVIVXPMsDER9LiYMHaLH6oBWmBaPDRh9cn/qQdy0
RDgajDbLngR9u/lPIocxEkg2JMgZ1UzxOuRBBZpOIJsZpSRkxKtpdQaC0KsLbB/n
qtkLSO672V8Zer6pLmd7V9aZmr9M/Y2l+3c/GnbnZJDEVrpstcTIyVuu5iRuwdJD
1LehNjIakJxKXtCtoWgkZYnPA6t6OHgJJau4DZYX6v/9S0dQunDPDU8a9Dsgqjzt
xPj2DCYhMi6gkFzdplRXn9hQ/Fja1+s0/OlIr8X3D2v7zvMslAameZsTiGgzW4lN
wf6ZasLxcjhKPTCMlYS1bQct5KdrFo3+Twy+vm/IQISzqbomiHL6qXtdwNM/N4hI
a/3eF4bTYltv2DlDYruQGqPk+3drTdHVNNEAc9OyPCW9IOR4ETar10AN/NpGRXNB
6VLm9FPQYeZ8ZicNviz22751XAY//TU9BBqR45od/utoFC+a5WjviEa0H699+EoS
kTwmig4s5wKkByJUTT7Tj+bN2XRBTyOurqfOkG5VvECWv8F8dUy6Ps86Q4dOAGOm
hW1RVrqJFQYQrZFObz9qVYB41Rie7MBMku2jQPLDOfIskTP56gB8k9+4big4W+oc
JxL4BSP+vj7MPC/Mi5yTxpeIfzE4LBKpDk++SqD2ItrLE40oNkfZP9OdKZot5X5p
frfv5KOo6ZN2T7s1mrpaYeZH/WLmgQdnOMUoBhNr7jN4o475ed0+Iwd3el9FgHIm
T/SyPmjOFVnNKCdrA2VqmoK/2wRcXb2wMENMSzLp8/0i1Gwjm6yDj3RHNHH16aTV
X5ecE4t9hB0t9TypUtg+uTvtEiSEWrQPtb159AzMuCvC/k0yBH8aXThlA71LmSHF
ArDyJnyPc/PbAWPTLxQGupS+JSZQp3MS0S7m5B3gaTY7daeNSx+lAxuRtnPcToOj
peyCuDsrTIw69E+gpb51SZV3ZPp4WA4KiAofMkY5D4VcaMF7pgCwWNRERACWPYNL
grVqouPc8l2OPdCWokbiRIDg45dEjZIVhmhgWnRnxqGKwPnhfbev0jM/lfBWA0jk
21msLwN+Rd5H1sN0YT3hhs8HtnxZrQrbWKeUZlSV8P18AqDezUaDtAE3EAMxt0Uw
8WMUkVRIi5LpoXgezyZMHnXbkmCc25diHEg6dqayy7b5ssOO12QAKiDFHbtDvJDT
xiLb3Y6WV/jRlE1Gz0G21dQuYXlAsLUAUMMVO1WRARnmT1flQ+61UjPZyLpLJvJn
v5JkpXJ2eWpb4dnVqsS7EwGXvlNZ6UT+KOZ7FpSu+OdjHcR4vapJcmC8NDXXW6d4
NtajW71nZAivWR5/9H0NFLnMOzWHKQGUkw/8PrXmZMzNIsi3q409APQwV1SOdLlg
z1eChnRPJ3J19wCMbJ1tBkCbZsfn36iLAamEfZ+Ybu3ByGMgQ0O2MeXW/lybJ4zE
l3L35sprU9NXCzEd3y9zRryHkcw9GHfcQfPvhqrA1em0d9E4QYdQCOvTOH5Juzyk
OYAgEV4aC+TAU+CnmyyUGkQaR1iaRoacpL708ZH4MM4II6KEPaJwo2lmhDap5YKL
i7vqCFJmXmLqrxrNyquB2d3XMvwLpuPyU+1Le1H/r3a4cQYNWockO9bPGxbxcFc1
JC4w5rM97iqXUBdgI4so4XSw4fxz1AQZJznEJGFgk4NN+LcquzpSXviZv5j0Ry2N
nOzQVJWIcfsVuJJ8+GS9CjFOSSvL/iBGieJJa8AOT5SuevOwwopYoCtYTIsXRfKH
FQ31654Er12r47Tf0kz9Eyf+Lsgs5Zsmvawk9P6gXhW1QKfkNTHujSWvpoUhPmTf
wMlqOEaS+Wz+m3u7X7Eq4XQ2R4KIlZ+9N/ICoHHJJrADq7ZY8V5AueQN3n9/fyYI
WGQaN31KXO2Q2ydZ06ZYp1S4g4m1LFOa3V1NqqpOIpFUzt3EQXKnrSVbJERV3NLy
ijgw45ES5uyrdq5KXlFLGI/vdLVJFtNUDYVDRqsP/t+FA3eJRlg+og98O6oUJX+L
nB3qEhRAb6YY5nkwG/RNS5RIw4QlKwoKXWWjAw1rov8RFvJpzIZvjty3HgAw5DET
DURObUSMMohYbAgn6hNSc2XYwWkEcuCqygSyF3ZnVWszch2J7y/GYmkEDucUyZOb
uXogpfLNq6nfWciLNzdu/913XHyBqw630WYSRjD+ypQpaSicZvLumwkfUoaaRuCx
hIa3l/h6Yyjxp2WrzEyHI5ASSW5ZnLGrytsw6K/jWQMvKoBV8dQGChp7nWCGnWVn
szraAEmMNKRhOkl4FNiV51/CxkL42gcO/3QBptcnJDAV5BMbG5b2qAtUhUhDEssM
7dbYchTZ38RADk9DO3k54+b7EvsDoUIwjDz+eMImHFKd9t6xugkUhSAD8v0Ye4kl
4OdAC03Es/a94g1p4rWgFQdEUJTOkX17VLL7keu/khxaL9VXejMUBGTsF6BHDJXU
pO1zpuqTmxAPB9RWY2xqvXqwEDQ+gtZ5cv54VfOzRQCy5SwUaskSxfeKBGtRy9sQ
RVpLjB1dDbK7wYtXROKPRE2yPOZrE+G98zlaFpctBxsUSfU66EjgTZnB0CPvkvhh
V/5uPqW7X+XKAHBfJ6IpzEER8X0jOgeNJUOPcai8256f0SNzxwP0iSv+1eiVm1uy
+5vF6QgGx8WcxwidEGZ0vh3yiSOq8f2pzKwXb+oMNoqw29JfCXlAXicyn5JAWaRg
mKivQM4IcmZMRYUm8ItGZ3gMYIGZR8LYrpdpwJm+ntVd/pNWsf8yNW5Mwuh0DrqX
iBisjldqAeQAE20BKHBtPjSlNM9NdtsoI2McGrONcuTrLUPMgl3G93PHrnOj3yo9
zTtjttVr7ADKrgmnpwS1ULku8eIz8N5VfgEGkkcAYgFxifdzVWnQ8asdOkFXZClu
WaIglG9Tw6hQ4z+SLaNBpEbZt7MwNDRAxqxadIFmdNOJsqeabvAZKl0Aer9Oglsa
Bf47mmAQyx+Z+PAbb3wkUv3Ea5DzrrhLkP7BhZ1FEpQFkDndwEh1OSVT8ePXBuXF
H57/sGucVDPe9x2dLLr4XIRZRzko3uU+jDkvYfsuETO/O023+PV3N+5fA46TbDDN
2G5XbQFNa7tglDMyAqKP1TvfH/ipIAIUfS8NTV6AxX6xtHlIu/UhymPD6IpEoOhj
x7pFaayeX0fOTDD1pRF3o+Cg/8n6YlRgDpUPXhA5I8ZuV3JJqTczbvCB27MABArS
OXVhgadJgelr/GrZWUqeludr1yowEcxHIAxAKlxhU2GkvHeN6zzIs+s1GWaEMBvB
0vobsSw2iil44evtzL68/SWWetv97SZJEO623B8bdwp30gEHR0HcLddy2VxFxlAq
BxZw+mOYVFkScygb2S14QzRZgNsiy3m2TELUHyWfzVhxiFBcLb9a/S17PD9r02xB
saQo1TMjq7VrFVOA2pEMicb5/bYud/UwZaBLcXiN8vY2mMYjxTHZ+Kb+EgYoVKus
uJQRCdKyQkOy46bjGOPBR+jH+4oUsRD6+b7P3MMXWM542tGYpKUXwlezmMSwSyv3
+Cz7XSfFF9lB+Xhv+SxJiTqMDRb1R0UT8lj1a4N2D0u74yg22ddTq7YmRa8wJAop
KhQOqNOsv8vutfvVxbQ0aLukLF2RThEN+ZurRq8r1QVDOrequZ7dipYGG0NiNT5h
Hnoklq/JXqCt13RyNwW6kegagBGVF2nKL/tAO4TtSpUt7ghfoUAowmztE8cXf5rN
6bQXWhHfrT6YE3OHNH/QOuJKsqBG/IHz4NEykrrkPlDxKlgfpiojMMOFGYUzrf4u
FBTZK1z5J94czzBmDY1r4ov9OpepzOXHjVG9NpjXIThJxy355PbTySJCS6/XRHMx
UST3u3ZE3YlqW8qeBKUG+LYe7PkrJLmbD4sSBPjTLMSCk64cxI7Fkkr5qZ4quotW
np/1OPeLCiCAoWLX9NBU1tYXkaaLok+mBzWUp9JV2KUp4NyY0LprTlI3xzgfwJsS
sIv/vx3Svi7xFP54NbLp20eTCcqjMt4PUyFdM33ZtqqkrxvS2cS7KJxoqT4kAB5H
W+jZQ1ijpf2fE3XRY6qkAYRTTlhMIHxz3czdINju5KQupR644ZmZxRj7EzCxhSFj
ODevv1edBxLx1vPi3RWWthaDatnzRX/toDPAS47Zbjh1qrQtKrbRXBW+WpPYHwBc
tLd5DSlXKY/r8MMc24z8oRpDA3ip+vEsIShpuVGE59UFZJHN+aV0g7yyvSjEtzKW
f816p3pwCeGQhTHZcs9IzoTnHu7CRlQ1blfzS6SrglsblRwirZUK83twsTvhNmgQ
7JwTezFABS5rv/sHPC6uNYrMU5phxW3LcU9MOc9X9i+jVeBa2+QKw1dqnI4ViZW3
B/NlYnhwA7vh1PiFggsCfJknxm/3d8RPUEZR6qdFwv57A2ya0wn2f5qjFjlf7yt2
IlzGhcyuf2HMs+ldkPesdPYB+X4tEAgOK3ABkW0hP8ZGLWOmVJOKjHnLX8L94Xu4
oBFyihEIR5UbzerioBiFxOjDHHk4Y0z3FJdtMDfN1BxwkL7mW5COclu1p4x1+aN8
qynFpSaIXyTa6vq2wf9jbevV4AmA7WdQc+MdoWmFPMSpneTjFuWXB9T9iOI9tt4S
+X/Xe94BOszRhU6iMtmA1wz7Q0JiHXxGeBx8i3e9Js9oy42BKFxiuCTyXT6VOu7p
0xFZbg6Zwu8og5nKtmGgClsSNcdLE/rNYyIoXIb9mlZGQQaKrP257X9jPWfsaLU9
dxv8CBe1ZXTuv8NjYKoQsS6Rmvz+QBYY7UkNfxeo8f7QKc05D3oMLr9uEYSg4mrL
+Hu5OHXFHLDnq68sodYcb6YL5NIuIC2Ui63qiqj2cbLqvnFfB7tfzJQ1gCvbheI6
CjROQ1Upm38Zuqm/vUkdVpha1LA15N5fNqYbizAWwysrNlpYxQIzwlqL8N+ps8oA
2y/E7fEobu2gcWxCRl2K3M0e3DfZw4mEVbtfEaUrI3anHpzidXF8IYn5TpADLenB
BQxa7twwkDSSYHVds7+lgvHZFiHvmMgDNX5URSR94fFSoPA1xL9fj7venzdOfvh3
imccGcdwtRwFxJ+mEShRcKuKQ/2bKoQUjitjDGnZrTpx65NWVSOL7bfnyzZ3Esvi
ief6S+wbuDLWGiTQ+ZinP+pRDOhxjn7Y1pHfjeAdCDBCS8P377wx6155xQ0T5Rjm
lvM4uU6SK/4qvAjx8Ex5ZmnvMEALKhVZITj/nDw6jzjMbWrkx0fxL5Ekonnh8Rrm
vAxdwDHYsSV3RQWCt3kDLHX5nyFPFqRCEbe7YUEagmMQiw/jANGQ5z137MXrREyu
1TOmfHifoq3nIfWOewbejlp13mS83cCDIf7sRxcfrwJ/xDIGtmmDrvs9I+2k88Yc
O31k2TwKeyAAfX4dA9PmveQqTIBVuEwP3dOwiN7Omh1wLSTNjKckOeiuVKAHiGXV
bZLKaz8lXKx+DNG5rlAkc23+jbykfdtFu8AbatXWJXLnj9fscQ02hR1oOmWxIZWP
eDCNMP9cj0rjDMgm7DX78WeIzRqEXxD9kdwyZ8CbarJKXYIK9Cl2TZhwICRIPToO
5ka0FHOh5yuFTz2jCl5JKjD5uxbmdwY6r+oIJU7E+ReFtSfJh9ta0n1CZy8FyMFf
n0jFd0h3kMuglMjUbuRdho62X+fgiqo5fuEeRfjhALsBrPZ+NI4nMJCNwtK1g4Vf
8XeZj50KDUoEdU99iVEeT3sYt5TS7YIuuAjfv7lHqzcTbkiMpE4irtOxzVWKnCdj
9abHPTmnHgzgMcjoQqvOtf21D7jTdavpGKs4JoXhZc4ATXYiB1soEosViZ6JNRho
e7h4jsCjyynS/NJXk7tblTkvbFsm2cZqp+XlMhPt0RY6f6jRTwD16R3tgcAJN+2H
HAcr/nkKvpai8ZMVdOU0Dwlz/6BJyUyr7Ie0mwOS3CVchSt/rjprYxMWV9hAGgcT
WT/ONvjIOR4aZq60I1Q985JIV+iu1iY53aI0th9j+39bKCwQ3qGLS/V4y7czQBDx
Lyl4QH1Zpc1Q5YJ+QcBN9UR0iiPCTnc4oJfdtLSeQuXRncMFELgBoPj94vk1lPAe
cXUonLiEgHZY7EZhF2WuWRABsHi/GaUVv2UWuNmBCqEtbS+wOX+hst8CPgKyjWHK
f6ousBv/MsFhtFEjtZ2wTQuZFxTB8aLXK/xvt+aTl8ruI+BAjjshgr0GDZvCp5dI
213oafvzUYCjUHfrup3N+NQX58J0FzNF7w9Nsq/9QMKT2zf/y8BbMqCZI4ymb6uu
0qcEev1YujuwlqOjlgZ9vRoNPWwcPy/ZdTiGJOZQfsMxfmHjRS1BkrY9/Pn4RcVT
oElUkHbpUT0MGMEJBZlGAMsxgLo4xuyEqkF3ve8w6cHpmidRppq+tLH29oD2paft
+FTYKHYK/+TY3Jtat1YpRTNIMQtDaZuLtl9KbwwmIJ0VLQgK/WduiPp/OgJJaDxR
IHqOugMvMfn+fxopsPfHDwiR6+Hw4Ey+E6ii8IsTXEJh6ofnomuF7PMCzqj7b9oQ
regdCe5VIl3dfrdNhBsem2PgGDPp9yA7rBuQjlT7F3cQr/jSEINjrIArTsaHAkoz
QpNKxudTFpHgJhQcHCOb6zfQdyNWzyax/I7Q+oQ9+uh+iVfgmWQpQsjtE81v0EPK
6Uz8l30SsZLKScj1YQ2lkiw/t9XgL+CUm2uDugZdKatKgtNR2KiamYXvfyNygTKG
HmU1QZO02/dCpsczh1mfaNNfO6MqoyCMLZSZqASjXcunsXVmEvTgcpB7oYWUA2OD
F1bRIoDcJXRarWqAQ32fqUWtL13IlNRVEWSUVSq8MOyCrJL+lZMqfCbInPqbppNp
UXQPzvqcQnuwGjSf7bkF/dWnbBBFQ1aGDL7XXbFZj23/jrqgUIYLghWrS0HJPlT0
K06/Th8kRUr6qwL3HIasIzSLGWYmNGwiwI6g7KV8viiEHNZuSl8eaiowjkIuM1ik
G4R3epHZNHVaW91+tb9cBG+BExz+pgKdQemMXpZo5IprhhD82eRe+tphOmYdu18c
kiLUxPiBTndc3aAwdvxF+tTBS5O1sYw48Cfdm3b7rEoFKblRviEALP8+e5mxaZ0G
seXadTX4cgu4mnoclLGSMUFKRB1c2nM+lW4FjeSF2uKfAIHTUjvYpTHYa9o78iqj
BvG6YHGPIRUkKfeN6D12ZAYmirRuNyB2plTVDn/ptUOC0kvN294eYn9Oljc4anaV
3bE98zaakJ+WFmmsaoeaKBTAH37VCH849LQ7iwtadgmKMnGA/dkSZ0gQdwRZQH4a
gCLvFU5gCBL0KefZuo7eQ9fEMUUaxc8FrQWpW7uqD9gpnr39vWBzdki5ew+4V8Pd
x+PR7JgQJ//YOvJ+vTwyDF+OQKijBmDtPDoPMDng7PkvawSece/n06k2asMidwCk
zOPrQOw6InVI78LT/FPrCLo/JzRNyR2NNJhTS7fQ9EStYP9jYCL18Q7/5UNLQZH+
B7teCX4ex1/CQvo+WqS/XkUC/pklJSI93buEyUhEQ4havKRpN/Epzppw+ZVDYJnf
WUWYQypIhK0i+Bgxq/ja2KmBDa/Ix7Hua0Pa/bIqP8f2os51Gn0sqrpGhzjOX3k3
pix90uGcsNL7RPgz/skmVQq86NJoWy8zhFOSre0TfPvOrm9+XtePZnRq9WHRKkUH
wf08XreOdBimodBCJvIxPe2SqoKUsoGfHdiRLZL4JklfwQwiRa3e6gQAyvyyq9n2
MlUVtoOQESQP4Lmn6Z2Uru1Oa1DDYybtZP13D+I9I0o+CFfC0W6yL/SjikBv7Bwt
a+xNXH/Ez/Co/hFcUC+UtM1Wy9B01zoBy9y3AkpwbROZiMYZtbat3cfCpWKk9LDk
Sab2v/F8glqVujyyNanwcir0s7TKP7megANyt1vOsWoCgaBJN4Eb03ajwkYVgt5b
S+H+GFiU5EqOaqKxCtgxOt2t9FlPp/Bqa2t9p2xxjNdkvV8pwHYWUPKdpYnS4QUT
VrUrpeGFHXE2aCkG9R+L1YSS/Rhsid8jONK5Rz/tVOfkgklitcZ/OYqpGpWAJXH8
NKpBrwelVAhxM4dzDezgX1ocFOxGIG4UK1yJlmI415d83Woti/qkip05Hu7DqbZ3
/9riuAd0f6rMeaLHslzsw51dXjyDNQnq78jtjbRmki2/GW087rFfRCe+AZdGIrKg
nIlv1ZZy81RdJr8YZf+3fT3w4QEfD6/vu124NvObClPuJgFyhEQdub3lZycz2eJK
3RuuqzZltRtAZ0H4wmw4f/UMJjoNOU6f3QKD9D3j+yEbolgakAkCqrJQiLGBH7UT
Mj/RRaf7BcGs+/rY+2+YRp0WmX35aiJsvRV+KlBDmVknUBKHOBxd0tl0vGeodrxo
JNDOJlYsc+76gIMmyQ7fLIJIq2YsXh6aPlNnnfGAlgkkrTayHBVn1DXe+JzL6YVn
V93aq9GzWKkoepeRaXltHvHZEHaXKOH7ZcZL5oP5IiaQVWLzK8VTiPn+ukI4jfQw
Tsk5vjdw4xToWdAbeUPYlhASMIFFKzez6XpeNFiqX8VY3qtbaa7alXV2Xr3W3yPk
Kpau35L/e1QISsK+Z/bk3J5Ub5yY+zZK29AUBAD3eRRgOc1Hq6OfGTlxf0TBJ2EW
vkfIZ8EP5boFDUMTyNciy4N7iZyPQfcsx3JXXfxIcj+QDqLTPfilufS2OQ2+ZWGI
lF+jCjuFCEagd5m8/5n1oOog4bLsfrS+7XMYAkgkHeBIeNQ8eXmC4nqXRXZjl1g6
aIsz2ve5itqQobr2NbOvUENvwebonb09SQqfu6bMf95UYjOZCuX8Ap1QnalCYEH/
bBtbT39MkNi2KFplqiOqYDslkR5CFZpu5liKG4HkdevwSh96vumz+OxkjZIcO1jf
2oUMuZMyV46lQcJHRb3BSaz6t0Atkph30Ntc31RMp8ZAO55OjiHVSxBP5I8V8oRJ
kTg6mYyMxocy7p0oYXCgG3NSIH9D/uaTlM2V+0RdsLwMlkFySZPytD5VD/3Lmbv6
ryKxLQVAaGFOd+Hc7M1058I2H/nUO51HSFaHiZkQd9MaXDPiz/v4OXJPriqWT3vW
uGbRv3kZDEDdGvRBjNN+1lqdlz5lZUQDG9kGXZSv8U8zD9WHiVB0OuLMthjCr8mr
h5HOnKB/IMPc31jgoUu0PBylGaHTsQatXTE9mfb3z2rE9urwIR1+Kym3VoFjUHfJ
OSacOzm8VWtbjVrSGb1D+lB1Jsz4s69rm4sl2KtCFknpIny+vFeq1tGR5F3bfoRg
WUUNVCxPZaMlV69OoM1in0DDHUFh5ftTgnGmnPBhSQGYdmOnKwzHHgiKcP+tti72
9An+U/i1diGIdGRm2Y7V3gsvgdxMpY+DGjxb++fN+JLUvWK5+lbHq5lwD3fcPiD+
m0wOC9tJ4on6/cbS0p79ioykGsE0zJdL3MLQhdoEfDgWOTqqoF3/fHbqrtbvOIes
mbj1npXNNRH5Mse/qDUpezn8b+gEuIiT+iuyQvPtKjkG9uK7lPVD5SEcDoRCRTXt
M9OCjUvkkBLIukDw14B/+HkQlHHGR1hwXnyMNlBQhv7lc2+SqWFLwNV12Bv5W5PE
Qc5dHwC688zOijApzB5LkMTElYcd5hUzK2TK708601HY2xD1KI8LYh+09A/TCmlk
7letmRU463YH++zG3FtnhlV/lxiqKmPLDJljd2ukogzDK8APbJ/35nnf2oqjWS+/
oQr1YXDuIR2ECd/mzOMA7bMuAseiyEw0K502Yv6bu51Xg4s/0c/GiFgR3Jg4L/MY
gX6LzKVDZJfsJiesI52FVG+rFIQXqeZdMfzax5vwmSpmGg12lavujPMmP0r1xxVg
x8rssRm6IJgScpDUXYG8fKKPLkSxYChx71rbUI/3c8unzAONfeA2Ngk9/BH1oePG
Xovg5G6IkRB5Dwf773Dgyrl0SquUnhgIFwETIDU1waL21NDvGaHLiTPJmmH26AHQ
LbjM3SQuePSBY5jFsbkOMd1ScdxpC4T11LbfV0xQq2+AzCcR1w0NM1DKZ1PoLaoh
wcCdqc9nMGBrI55m/AVHdJO4qc91U/Ds0MwriD1Jr1fEN4+LNU2BCji6NNkG3Y6o
ByRRjxjvBILVas23ioKKKEXnr+3w9tjuKaYQ4AFaxU3H4QffBjxjDkDlcxxLj27z
/rHShMDRBATzPjVd1ufI/yVTxrtHPHzGtoJmubqDNHMZ4G0Sp5h0gAnHOnaxbq3D
CJPBJVXFT0H8jgczPsoBhk48b+DfbCHDMvWOUEQmI3nQUnIT2gA4j/gWC7jRawIJ
JNGm4alBfYK4h8xMwkyOVY0febuqqJzPkwKm5lrL3M3Dn1vjjsp49EV8RFX8HfW0
xUHIP/gkh6nSwSxQrzt+gUksjjhtg3d51oKyqJ0OoaaH+QJFwsRXgdlBbrd+b3A5
aAsLrY1lwBwRKk9igkHfx5dEEOtlws+GcNZI8Xvca2yFegsih07wHCAZ/YBMuHK2
S5aihdpkdwJtMW/EO+pLsP1GTopKTLnpWf7/QMmR00fTI9szRFSTnNkt5PKabgTb
VH1GNh+Jy9XDJUF64gFA90dll8CCuMw9ieIYJW/lfF+rzKTpnNvEfA4CfkW5Gw2O
L+O5Ukw2tUb/6lclbtx5i3tR4qkF2SDemRRCCF+FkiHylnC87nRrfmgDHTN0W61D
WMP4Nvlzb7EgfD2/F3G68AzP3MvXdNF2LDiW3vRp/9kHlEOF5j6XgYvUEWIRn62u
3fSteu4wEz4iXUJMJi+AlsGYP7ZRfMONnI+IeXoHbFwWlkQK3K7xtYu68NAxJY0x
7IzLs9pzSvcTyKAJ3CI1gAefecIwsi1P8SeQnD7eF36a+F0TwU+5lCVLlnjkAjBl
i0DGoNNTzUjLMQEG0y88Xi5+8eD4K7mq7g/ca2bTP3B65LAvut5ZNkWPFUArEF73
PG5lz3vMwD8eIlGGDiy4Ay6vJTH3nbDThYNO/Ui0ooq++E4pivpiiso4TFL2gnvt
yAL+R3trdGo/8iHVYB4bKz69ToSl16Yq90KuUaen31W5lkW1GYV477PSNe4HI6CS
FwTjWCzdFMLyajBvad4s3Ia6pk5fpbLVE8PyMWVQp3KRJD5xJ6qokBgvBhH6ArjU
sIel3ZxRo1q0ASY5JcSV5Dl3wQGhuzNqeposXMzR/wtp9mC4Tyjf1YNiJdqHdHPu
32ynwujyYiALxL1vJ2xjNN9/pobH31lkkSLcFeFkWt0yhtHw4Z36LOF/AN71WOQJ
zCzgkoi3FiFDriLdgcv9GDc477nTApYz4QjlcoDT4EgfQ54DPW1jJLTV3CpREh2m
Ynnqk+wLMD9W3Mg80T1ac3aWU5uxuWsd9+tKNgIK5Rz4vKxPFM1BBF5xBf5OYE/J
ggEHunds0eqOyyMSMfLHifpzeIx6hrWb0pnx8g9WkzLWGuUfq5dWEStFRd5UKAco
k0BT6QuBjLBX12PX+4BnbLHBYI04wJh5Kh+SdQJl7lRU4X2F1LxP2+K+KDFAsNlr
FKsmyQdo/+uJ4X30xto47p2rZtSRLTckXIDgAeZ2e4zH/At0t/kpRLuZedhSj3zw
UUg0Ct7AQIcyhIVhmxr10nsb7Qsh/NxKrmlVhvoui8fLtKyTgXORwYXwos1m0xuW
v8XyjQgyhK13TEw1U3hDJ6/J17UtBkxRnMas8GG0w/t9/YqDMUmZDfM8RHClCcVm
850pECXHUAoVvl4Vvc+jUdOKkJ/l3DrAOQcEZwcUv4bdIvL/19vpvhnrAaHony1H
7Tzx0OWRc38cYz/0SFsQMKfTHFhHKiD8PJYSqZnvB9SzhYDEBgod5b+0E7O2eLCO
W2+pYojWEdiAgH6MvHzTYgvGgO0PP0ldTKHudTYFf6hKBpEtfA8BunhHIi8nHjq1
WzSQnhg2ycIrplY9Ojo2dRptVxp7xEFZ3otHhilyAGL6unVxImJ4c65iRDmtU5MH
YLMNmQx3Nop5VerPVHGUZzDgMEr4msXrf8T5pjF3hgX0AMUV1tMg8FbPYZO1HRwv
lh0vZr6I/+/yMQfyZpLXJQ7c1xk93FqR+m+DqeIMmdG76nINjE8DnO6frUvS/miG
rJKC/ELXGTSCW/NtSVDaSmDplezaRXwOdcbOk6hvQIHBKDp9dJn27P2RFlJ3atDB
0uXQLH9n5JfkzCe35xbpH7TlZedAZbmQ/e9pKtCcS6BnztVlzjwaHeRwSEdkB4BL
IIGeZXxHa866KH02M/Z6ACiN0fmSz4+RtIBOqh0/FbB3yggDneihcWW7ckWcEDAL
1rYmfXbfyhMar4Ylt2RS1IUgnljqQ7k6QlWSi9MKLL1py15u/fes3cxcnH1BAJVE
CfeWWpFxzRKSjonK2BlvEoT5jtDg1TaXDY0tVJGqtZ7OO4I6Eqms5JMjIqY9D/Mb
TgdPPRgookrhxiHuoJRZg6dZAKPKkMOqy2botZbqbkhgvE9DHItQTyDR3YhNirSG
51rw3WMf8J4tgiS+duKi/+INVDGYvBS8VtDXZnylXsHLmLCSUf4hv4GD57/AfV06
dgPDqEilOudb8Xg8JnI9B/mcz9DbkkYqQopDJTa6z2iA95hG+t+zkYWO3ElmLiHu
4TfCO1YSB8ddY3K16fEYEj5BBzTMsbnDAZTe2bLv4Xb8SfZ1m8KKhc1oBBEbgRDN
p+wfBWp+fohU9P0V+dlcrAx/tCyajxSOZFn38yDe6nAOeewbr53shmY/aZThNyk4
9pAeC67svp50QAyfvX9Q+kZ5rv6fV/KDDV19pGvZB4YtvUOe2LJc3EFBBlnCwzZ4
8EpbNxtQW8wLaMfKDgp/ES8GKFfP4rUE6CtoDvJQYlPeCzaWK+nvxLlefXObzp9N
nMy7i26kvtR02tlKNvSWuHMMeWi7kIRdxN+uMM8mXBMX2Q3P2b3kgh6oYeFu50sv
SdWvhVTeI1OZG8mZXYjLOTNQeEN1fTf8CL5P9fLvigJnCyzL7ZAU54F/9kueb+cZ
ggVc0QB3y87e+XV9bOgLnHc/fXII2PbhycfMMBulcsU6qMJqF/IPzVEpBZPH3HIf
IwApUFkLaAgPyTm7ck7xZOTOqj+4TyNF4Vdwv8QL26C5Utx5C59ia6o4u4VBJ4wX
cqJZfmsqspA9CbkFF0tOtOMZWoUPeHVtaHN3NeNZixTlDIUVjyR7NG39Y3u8muzi
1UP/evXl0Ha5ubFaJQ/mQRrWgRkofsgojsyGe1lb3L1kIhHS/rOetLIlfa4/dpUl
zq3xSd6UFdZtJXaDNYzB5/A7RY03gN010pN54NxmvfdDUs3aFOU4dAez9rp92mtk
jLugP4rQkVTKjt0xJ4kXSt2R6sK1uhkXnMxjAUQjYi3SCqnN2WpkYTtTTKKv0Stu
nzK3HJK+ARwnn8zV5f0ajFKoiVqwRZeIJPmlG1hbLyZnVpPhNLkCfsE1N+0R8BEp
RUFb06VlTLZ7/x5soZ/8qYUvzmiBiqhNDSNjJ5QmzzXHcszADkAMH9H3HX1RQer8
wKMNqPT0bRmerggywOT1qWCrVzBYD+1uNCVFPuA6j29KxM70AroDNariPaFEqWCV
4RV0Xl6pUzBxi9i5ShOCBmfbeZtHgIopq/FGthn0Rya+a5k3OPUe1zDTw32tVNLo
Xhrqaa89VS7cbxhsWTXU4/SF2Bl/9v6O7tRywStTt4Njj9RQ98OWmi8J16XrKraQ
UmXFXG3eULROXY9EtRAVzsNk/Go0KNcXMinlj99Zh1JD0jnUyl5WR/em1bMFdv37
yebbN+mwrlFY9LS+tKm8COED4C11ajtHMfwQtQYlvQMO21CJ1OBwBVXkzeKb9YvS
IDAX/FgWNH89a+NozO063wktqqe5oA7bD1UzZI86y0jC2k1fLlveaOBBFOFjvpJj
cj3GzShqT35XMCeudoCGy8C+1is1wYwWTV5GtFNzDf6NoHHk/WnXXFKLjkvSd1aT
zYUP8+vT3Kk47leURaURoWgPLztMYcZgewAxjsQGkXovfRb47r4M+nkBE7+RMTOe
XF09kfFW+L7y8rRZ1sRrK9diMeJgirW286brjNwWdug7HRiUcfsI9MD0uUw/kweB
HElsJriYdqebgSY7nwzc9B7V/sPuMIgrABYxeMgvYa+uUQZbRgB83CEiB3kbGy5l
lIhPsakgMJOk95MYhn+DpYtgbyXotzeEfAwr5C2rrXE2JeJst/fabfcB90JZraVj
HhyxodhpsZtI2/Rnk6vGWPC6iDNYiaFPsYDdyvmlzeniCKUxdaWdWulC7xMOvfVz
6r8anEpnymdVkK0tqmzxzMCLSiwWRB4MNqmubw0eAHNvhIlLaJXbNKTSQ9l9XOni
VxbR8KsbyzfFafhp/1A453eUYFGUr2nTU7WRFLxBymNY+57kxC++XdBCnSVcOj7A
nOqIh2dflCcobM/V5lmPYU7iAb4Xd5LIPVCBDUivezx3rKHb1xDjWhIcl3omNmST
lSLxQi8FzpSwAo1mOtKDOv/aUsQVf37CwIpCbC3I3sws+dTYl+0qjf0oko16DeqN
1E401yzVdiu5CAgDzOuPyAI9k1Zp6/shUfyr4JEOzqViQa+GUBEsddWA/9A5N64v
5usMSelEc+f+UGwKYUnbjG2HlfTJuCu/oE3KYT6wOfJoEmkiy3EQT8RySfCmvzm/
OXIhP8ZAEtTx5KGU3fnw1LUfN/TG4cEC79l8xBYOC+Ese2uYXhkGMF90ckaVvohH
EA7uWLNZKQMmjHEWF/LzNJuhcZOfD//8hDAhsrBzhd9L44xEvADOPmwozVz/OSLz
OwUOMB5TeX21XbsDa25UQAt249eIRCARDFeSADRpz4dWW69KFGEb62L0y5hkG2sU
HCyy1ffXVFv2uC+Su8BtDfopIN4pzeAII1ppIwS0ZTZRmE8BWFyIcjQh4JyNnEUM
wdlsK5RCt7ySoh0MlhE09eve7mL9cXT3so81ztmG0iDm4SloRSLom3fGkd18H9nW
Sb/hAhY1zK09uEix1LZ4NfNbDANt924q55vKm8yvZlLTYg5zgvgTPAOhxv8zrrEQ
SxQw+109rQWH/6iarojDyZSDivlXlxHK6iN+rSgJAZbUvwovaOM6vVn5YNz3hr+0
o0zSnUDZHupE9wtGN3DJyQPLIZ+AKswYiKeMhYUc7pm6RsHNUkYHsoDTFMVW3qpL
OiK+xF+ANxKZSNelFHF8yxzkTVZzXpK1/9T2+ctpFAydHjdX+bzC4c6MEmoLSc5l
/uov/wTbB4R5UNWgdJe4Hb6U0Iic/zLYTQs6NDUuwCwLxmWgFzoDNi99Yfrw+OUP
1m/v+ttlpSWAo3XvkO347jCc2KUlP/Nm9UctAzqtUDUwD2N6b2wuKyoFLzaJPoop
hO5etW9OAa/LQa4tpm7SCgeOUn6AMcGLM+hVO1MYSCiEHkCnlT70cGj+4Tq6tkoH
RpZfTBsX5d8fVoU8ztoYQ64ag/vz8JxXppryLyQpuuZNPj5sjTOGq0nCcCYVud6o
Z+l6TlUcnM0R4ulrpK9IzVjHvT3kVGDpaUt6V6PVADKrQHu589O0Nm2oZtiaJgzi
NoTxuEzKBs3J8lUendpnFX5WxXE1O+lsCipSRg02WVl593wU/y3kJ/Vs88PHRxKo
jaSQqOFoWb0DwXdeXrserdaEKn1rcPuCG4CVbzflRxrSQGkHkSt4U51nhm9jAqC/
GVPO0Vi4wI6U7F9c7Z8MnFeqJbpNyQMgU+XNaV6ZbxI8bRpi/niOeZfrgn14E6R+
CrP9qtlUua+wUNAy3K/MAayiA83CKNpJgcoFCUuuG/CGUJ0EfikWSwPnsrQtHYkq
8At+4ZCJ9jph6/Zr5x+aHwRSyUKEqp+8oEZ5dMQpw0W+cJ7MxjmcqzCsFxWE+MM9
TbgExp4HDa3v/OJvoUfW4S/yzAq9hShhd0EpbgwQLdt5NzVbhIZcInU089HU91DY
3DM4K5ns8FzhBMoGh2QAy0d5GcOWWHYLTlpQfGvyNrfPPSyMDg4AWXyWwWvvadDK
b77R08RymSIurRGa6vzNfJegqrX26h6i+cBA+R8xgKlpSG8YWde3gAIB0MKUCvVS
DaS4+xgSqBF4YtBDFKhy4IcH+daW8EoaR3aZ9nJgydOLKHvuvOOYvHd93AbhM8ev
399MTCVQ8RA+hZSJDgjtW5AZkJUT+UEnfRrvDDVTXYs6rqjV4Vmmn+SrBaRW33hf
Gv4bOS4Tt3OVjA5jsKD2QmInSy7Zhv8NGeYblMgpws9x8SycRM3tDBJdqdJHthQc
XVH6n39NYzEBushSLBjuM1aXLn51vYgkoij5ea7k0mMz5J2HA+XOcyiPy/q9TDa9
+a+Xfn6Ra55O7OXR4xnT7HrolswxnGIJ8J9U0oR1P53OIaHRiZK8vmFN+pRLIcmt
qINGooWIt5KwwIGjFi7DzbVOoRpqrDQ9lox7NwLekCl7f1xcMmRwGlfDo292YRA0
pGt0VPr7woN3GatCfDhfCSz5NXDlbeZrQzj1bK/frQ/pscF99YYbbIyCgBuu2TAc
Tm/pVMvbxBT8XrzushPyXkcvhg1eV/4fhxUde8QCpu9BrknYfb1FCO5sMp38V6Ax
79o1ybq647ZVTXtrwAZgv3kRUgyAwBu/UvAOiLOgUC5EsorI2lc0Obp2qJKZBoo2
FuPEgYQvAxOMDyNU2P3vRzhCiaXW8EHEbGsVU8tbnmEJEBzvGYJKcDEbEy3uWX8M
kvID3V7ILlkimc9UEDdIDa1L8311vB6QVhcIRyVeaLPPByGO7iepdElPfns1NTwQ
6coKzZIn59noXQRWYXh+WWDF4oSr8IUV1JAVLFJVKffplEZ0DfUnb/uUlm6FAaxY
fHrqMhSc/BfzUoJlxWs7+ub08jjJ08KWIvI3k9XWSTIhWQ9ZF6hkU4uzq8Oa/DAT
CzU5TgmOs6m3T9376FBsmXVGbOaOXy218oodVSAf/GqHf4Y3YBTCZgoJQjP9FZFr
+fuZTnWDCvSzSpQHsX/isdeflQ5fKHxTd6av8Hs3gn4q3bXe8S4UyV7kpYx+HXJ8
GXO3e/PAu5d/CdC3KnsINDT9J1FVWn6RjPPpw19+NFhnhVIHofpKfrrfeK3GgWhw
iJB3XNGQ1uNkD2EL9savk3xROg1w/WjcJHepY0aF62sRLWmio51nwv9p7g60V1TH
cMAf4LVIRjrC656m0LvyBi8/sIx7S+wf1WQlSc++TqnlCo6c42GajbXJs2XejmD2
rwSrLJIA08ky2Of5KzFn/kfeKvpeyyFL00evAijTSYdZG4zY/Pi2VFrP/SJ/1pgL
l6fEshjEJODhgeQQ/RUR5Qq2RliRrIQeqnz0CuXumwakZ8DsGr8RmlSblyd7CuIL
3+IoicGoD8ctwQz0+CNKcTv8t8XOQlLUZ63U+Ahvvt1hSmq/C6bB0ie3/4vTb7HH
xkj3exnoJyGyYwiQEr9DENdzsy/9lsgD4KG/g+ObjkI1mRATKayzNj6gZpPVwrfA
uQvaTseUEbAdMqgMK1s46sDj3eBnOHXXYwxb7ettDxN1hw96bY3HeVIzmXe8N1Jc
0hjUuaFinz2F1+2l1sxWgCCNH3687rTtf1SMn8+QGOBlNSZkEpwBcvj1ynyiN7nD
WUXziAw3uaUZQjJMfsb1Z4I+YavANDR6rnM5FvM1miVryAeJEt4F9UKoiviVSklR
z/DQyc/GbYoLCV7rEnq8+rA61jA1ENhiPFqsBYAPCqu0URYHla9XsufbVztSd0ei
isasAHavOfnLFR1VDrKVC0NH08s+01BOx8Pq46jCnMyRRDb4kgiIZbYQ0vsmSPzu
CUGsXm4Rjkf6wHlsc2imKPvnoEvpbxbDytasU0GDwaj4GXg2xmux8jZf5JpTtXHC
herwoFJRVS3lELupwKEdaD3PvHdaOhmbem2yl19efLOHVom7tTO8YQYvekYvkCZI
er/cKlQBvonrpmyM36EBuhXdugPFhjuOYq+h2pOpaWWNURuyYN08aW49FMjiGZYg
tSGWnQ+xGOabrVxPNIWGJvWARPvscfJM0Nb/9MiWM0kaDedoGRT/QiFDUBwDQ+Dv
iaNQpwVrs1sZITtNYPT8kxotDyEu7uIhnNFKVxrv4hbnYWi6BLLt9sTJUo3+dkMy
CyhMEi4bKbbq823l0nfCtVzZd7yxzTNXbTjdExdnKBQ8xdR3TMtHgnvzqyVm06//
Li20bugXOtAUiDyP9FStMzJsImPaYOxmuCUpDADiqs8XxiO1EGUt34JAJKpOfHUp
mbDA7FluMuGEuUER9ABtdsMA1R2vYrItzAdNyT54mtcF/U9yXya5faqK5lRbHUci
GKJP0a+kgkVbglB8rfNBN+yQSXb2ZUHH6+QmgutwFHvqu48f6EyULKXrm4gWyDJI
u5JyV/HVuGKlzf0NGtLyIuFJxWtbVI/wo+V8aL7L3/FFEDVnYpven0AKViYBu3Yl
gnaKgThp+kAl3sFnVfU/r5scX1pgXzwRuDOvMAzjj/BsTxwHAjQeZvZTZYbG1vTL
tM8u4k+wGQdHUVRnlelQhvsy4QEb3txB/GTRx12bzZhsqiAhH+XVipRfQVM77zJW
Yv6upmh22nOJoa9uYk4Dm90fKa/5p6apmrI2/YoLSvj5mkJiL8bD4VNRnPHqtJhe
s/anylEqlaU/9bOazSr6rfbAXtTaCIQqIN5CtT2Ftrv8wp1ERjRilCjFI88UvQOK
0Z5kg0dJCQ6hkWBMOP7mSEbllGzq65kqW48mvdRLFVVReXKHRWdmPtXB5IN8pz6P
RmIx9vOXiixBZP/T+efYmEYqa4HIovoSSGLEptvZviBJi63aba048vhCxpNmXXG5
x1KacFUzygYCpML5fmi4b229vLGXszZZTPKVbUEYrF0EvjVobEkbrEDirDGmSp98
N9JPjp5yAoYWbqgu+atxC5VwA/KfQdvumGNUtiunSvib8t2np8vf3So4NlGs6B7O
5gKHWKZ1+a1jASHDgj80qtfDWcPxmSdoiuMKqOi2Qub5jvIK6iui2gUuOkMFX0lV
YD0N4uQowyTZt86IUmkI0WLPAmt8KhEpCRhA5H/GdtU2otRZ98jgSn2xJz+6Z/+G
zvU8+gG6/RwfP8nAi1DgkgcNIRogN4pM0juNYAdtlY/egN38GJZLB7/a9ftRh0+b
nYXSCV53nEdQuUVJp0gq4BtURzQTdSoeS1P0PbHTVahTnZfzWwg5pgUVkVH47ON4
+exhSOZ/+Poc1YHBv3rZ4nrCPr9Njz0mgWw7HivbXXnmw237f4bYq4VxjyyA8jy0
ISCOFyVeMlLH4rRpqYrKZNxBd++mlTboJZRg0WyQMeB0pSX509rtXAvXoNSphKo2
aMpcRpEwUw4c3tCxehHO1iAyKhXVh7x74Lh9yj8aiuQEufOuRhcOFPb0/H0vcQOL
bqzO0/k8HW1zQfomHaL0rIT0RrDW3NZD9WNbJB88PTNmq51n9iFBJD8SnS8e52ic
6J1B9Yz1chR5l5gsD0FCqDFQgMdCo/oS9hNWQVPrE1dLJUTdeZsz30fhEliYqk7g
VuN+Nh3QbJc9wsE74ueBmku2Og54sI1EEhIiW7bU195T5tulu5TFuVq6fKlm9PTd
xstD6WetNl/JT2sjxJ3t0envdxPufYf0p2+n+HAVHCNGakKWllqeqYhZvBPbGbLj
jsggPxXYaDi96gP2yoZB65N7J4YjRdEBl4YMO81KGnexwsipb28xe5nfxt/H9S+x
xFe/qRIPYzDsNXu8PMna/LtO+i1fh3ie2GNdHrh9c7XdDu8bdvJQhvvTYpYW1UDb
KPoBM6ppKr9eTtePsEx6c6E810C3dziq/Hi1XAwaWZf+zDERMWKrdS3TyUi9GCy7
Q3dzQGXt7cEk+B55o+6SRxle3soKbcdlKdk1Tx9uyO9Y6P6QLYb82htEs6jCbxdU
N4j7rxlQhUSTco3SdG3Xd5cJHMITTzn6fN9p5Og8SofuZJ32mbd4cJPti8fFd1Mv
1aGRV0IGHhdqm4OLG0wC2PLOOvCr6OhkGWrS83rJopFsbi0tCMk7KpUCDsqobSaF
1PMGpfIq06+aZk85GacVWtUcH4nJ9WzrSCjKvr40N3m7R1TBB91LgtpL3ehhlTJE
1loDR4q+vgFujsQoGftfZBtSgQh3oUnMFOMiZbfTXTzC13MkU4eqkyGGMmz+0iSz
g7Y6ObbZHfwOy3OXj4Bsogay+BpMDs2sHOES7743UsNhTyJXfGiEukNq41gTWDIq
OygrsFqkZ8WIwW23QcrM+GuwyKtMhgslIAfIHb3t1FOmxwwgxNFQbZhdb/OxkAHt
6aOa1BLdmovuSBPsjhzq9V1Of39J33P8/FhFet9ftQFSpFMTDlkVqj4eRbC83Ris
2AxVy+YeazLHSaTAMh0HXghrpiBPWWSdIQQVe8sHOLew8njm3bD6mdZJ2SIPct85
AfrGKJZrwPjjtgcgjbS/BTYjEkmd0ajLeNhX1nq/+78iGmVFjMxbrGUEZvmD0sNk
+rnu98HHJxRxHgi9L9q1unFwxuv9KJKTAo3f3YUK06VDrnv94WN0MMa5G0VPetgi
X6bOQoQP5zIH6RfyMgH8nnTJxI/C8bkMfbsEfeeNCmRU/8AHio2NM2/swxkDJDA7
EpY6DQJzcv0CyHC1D/g8zPSrUZmGTzibM/iWCujNNvI3MuJGVsRQFBIPq1Fm9kLB
D1jgv+7uZOfncbAWQvvUI4e7nGurLECZGR0eY3QWO4YDjKVCpe5BVrhSxMqOYikb
MJubwYHaLbREh2fTAjGCG4AEKutDUFSpuE8eQcnAxz6Ixy7QDenF5nz3ufC72OFL
oGBqCL1z5xyuz8+GHv2eq4IBWmSdR4V2sSO8Pr+CxBWDsVR2b14pXLHh+zYTQKve
MuDZYmoHkR5ONv90k4FlLh4hHgi9fe7p+YO+9cufiMTaTd091WLH7uowr+ZbXqVe
TxIywD/PMIeECpHuvigWQprpBp5Q/G9sTMxA/83BtTfPoplCOZLKqbywpUzti2ph
uUFYENwoxvXHFbzbI5R5L82mMCfsCAZzsQ9IQ1Ecc41UaXGvZSpUAl4qTbuhXWLf
2Zbx4gVgKRHqXsTGijA7q/j+lCXGIS+iLqImfyFN2ewhKUVlQMHoI2AYHlPZ8tJw
GwLQJXan6bs+DxyLbh1HSAnxsmMu3hhy8/nmSXxV7vo7Jb94gLlkoDRVxwfmlmBa
M1KTC3/TGKqA9aZMLiG143MHI9FEdqvyMZoBlK84Vi8I8WttJ1evvM4M5SZ+4hTq
qTG3BjdDJgGn2gacpQJ1rDo7cD1Su0dKslWK5IHKVyLMu//CyBQSVpWBTMLaa1pY
Iiy2v/6R7CIVdFwuYsj8Lo4gr685Bq/W7zGxZNiGVOErnmAGD7HDsZ67810qvtjB
A321xNticnQlydlKPLY0X4SnrlofcDnszop4j8pNTosfQqCso6Ah2DlbUvwvt42Z
i7n71Q2Vdmnfv2ltdWAiHQ9uOzUgysFjtkL0mOxohbnTpz8U0hMuDwWmCr2slhz4
jc+ye/y3WxO2yqZWxpw4fWrV2d4jWisxO3/kK9/0+35NOD3DLLu6lZNFeGRX+6zR
lMO1cWogWrcpCigyFBLYXXbiyFv8NiANlj+QfCevGqtubusPtbkRcmBMz01+pRQd
TvW6Muw2ZGCLC/Nm1mkzLQpSU5WVltCDksREu6BTPJxj2kW1TR98OGsblnT1Drwb
qUl+fkegi1MIlrmavqF9EsTZ1v+pCVi3FBgHCMlNPqZUY61eJBT8340P6kgLIfzS
SAceZd0QpN1H5WPiKnWykc/N1FDWCvyKxatIrMgWiZUP3r64kqVmhzHmkcaddRig
O2SZmcQT1cKREb/mkV++/oeQk7fhVtoGTfoDqehPwZxPuOJDI0DwLDfqhYzKMikP
kUjQUAkgoX8HqEVlsRz/l/1NkPNZ1sOzUnaenukmmHZOo14gjfYpqSRIzO3x7/2b
yddLATUz0Rjlc5Hn8IXdAamOfmLq97S3R1yjsBm6dM5s9S8c7tfuTOuxbtWlJgLn
4+7saEibFRutPM+rDUZoYwtt8S1mTaF7YVeHrR3ZYaQLPRHK7V4xrQOQhBiM7Hkg
wgc4jJSFogwwa0dwVQq3nqTRF9QILvwT1h/ss75gmeI6nkMBxoKbK0j0NEytuDNB
wnBtfGbAMcNVe9TqlR2HCpVnNZrIVxBlQyQZf9UHD0JR5K48TWtbEri75LzyafcA
ZHKqGyvnZfnhDy91LUZPjKbJDyIemDpNG3pTyffNU6V/vtS9EQXK4eu3rP6h/rFA
+Z2WUarZnmyxnRAM0hk5N04XO1ZI1t6FBDAXS6PgmIvJ3qv+HtZ1N65TT/oTy3dh
6FqEfAKzRVk7nRFYNt32l3bL8W27Nqi3+pUhsBkxZLVIQsrrjFce/vsoahQDLHOy
sHwXLRpl6SEgx6NUt7DzAb2tFtQFYGsv36fljFkcTpgyQc0CxYsapz7lBWJ76/YO
aLQc5WuIB6f5PudGM3WXJzYi4ZuEHA1Xh9Ltio5NVmFZGytS1QZEmcMNkf6vy61b
7xq3Vd2EjG1Mck7EnM19OipIrtSvqKqlINLpHQCvoDVnQ1wSguusNv0ElELn/Dgs
OSo6zgfcB58msYuzCjx4kLKrd4rA4xxtqdGD4ttfEMnScWjMnaoodAWW5Fn6662V
bQ1T8hT+Vgw4hl5hUMW9ySSDScdnxchs4kzktfK7hwIZPLXzYAml/F5zxWVstTFD
M4LvCAXpiZ8bsvPouozZ7x/red1a07M78H4c1aOQaSo18gKeA3R92ffWts4grCyh
2Re6JvdA5q26EJBdAAmw7f69jTEACj3y3ZuOMCPaToHprkZuosx3GDE9cfysbHTm
FpgaOKuWTlg1InLJ+CgpERxB298HqB/6VFsEdHsXz5LzIzYLEtmb1kQ3x1AJuWTk
kmaVJAPgDXeDzVVzyxwucrVjjz1YbBAa3rJ599nL3ixP5aCCfSi4neIeQtjUOYM9
8C5sDjIDpDcxYyiZIyIkjHTvUb/whVmBAVxl85VR2W4XpxY0vfE1YUOYQ8unoG+H
zw8AlqMj5/2P7SmGNpAgi4pDP+/sd4tEa3AbCdFUaXM/TM6ItTYSipD6q7cTQ+pb
v/qAzNJaRZWjRmpDkvXB9OCRPGPQDhMXVQUFJeHGT4yIgO7Z/UX814rMMk1inmel
FJL2jiJAXa3AI2++2jCvGMKq7ozW9hmwokJFfHQ+VPEvltrfapuz4GQCgIfNl29l
ApQFWaxZB9RD+yiZncEpnuhfE/Cb+mqrRQmBY9w+mbrYHKozxi3YdAfWM2z9A3OD
jOcRiCPSdljFfyPw6gEFLD8R9H1TuhjjZJSmQLx7SrVtVdYm6ahVhx8+Zj0o2/ps
o7JWY1vmL8nAhDyOd8XaBYKfcpvTl5T03NEtUij8tZPY6vWCyHJJg28RKSbEWazj
/U2d8UCSR4x1WqP3X3hSAJ2nfAWLBAxC94mKbSfKzcMqrKf1LArjqxXI8S2FRNhj
PmcqkYQj6T6xX0+QG2bpi5kv1qxJISYtX6VYJK+lC5C12z/BytZEowQoaB5FtDow
ZN8Ve0nA323MzkUIa3Dqd6NESSQ0+Ejia2Hux5K7rFAIXElnX5ve3G2fWjNMRIiS
IBWIPcqjALLAoW0bFNSZ+MZ96ko7A04AfUMqZ86nksLBcHi0Ep6cn39gxyMl/AUw
P9OlR6e1MRDTKHRR8S1OKT0/eUpluJYGWrr4Qnxnluh4D4iXi1dqGPTsGRi1DMN9
RNs05y9Blq15gw5/z3QEvSKM1uQH2khyMIj6O4aZxBh5mNaXgvwuABhVnMel0XkY
qwksQ9F2OqMXSNNZ4pev7ozruVmzFHksCXKOYWdLIKXjYp4QuuL1wD3Ig9UtU4e0
gbiAazPFujGdkXKNunc/Qqu8AOckPF6kKVQ5EGOa2gsIPYs0NNPTOAhgbns29wmo
YROuQkWm//UVxJg6ILbPLJwx6iRFaVGBYv6Tx+xS98MIAU7G74eiP9nbwrEeCKYp
xJ/NHH3hgjd6yK1naLYx4MFtGpesOWO14WXfMn2RW9d9P7tSFa1SgEHz8GgdiksN
kvCpAA4ksUqdVvb0+QMjX57wcyZ7EQKzTRwBHlMPRUnHFOkwqh5X5EdTibtd2h/z
QQ6i7T+3KsiYHz98wkveFp4g74bpmnCaUHeYw+AoMkHDdiMMqogXAqIoUz1HmX1e
KIVcVS7wyeepBxLWEcEol+Owgfc+RZ89krW7pQXV09l1U5qb2VI0nds0gvYDn55F
a3VpqPAlYkwneMXtbgr9VNFtFAFprgVjpphyJXZkiuKMXppCkqiEez+yfTmw07as
X+3j9ujyW9s9oJ7daanfZ1hOJabcY4LbJ3cxCzrJ/ance2UotVbuvdELKVzR7Wyd
l4llByeKCqUQxzYM7IAgFqsEZwjwQpQZCjanCSpbUZ3KoCM+5O3TmO81Lct4BxlW
xLhwCHGxsfbTUbueM8b8Z56PuT9UqYfwLBAr4/SS8Tv5ARgp+u+Sk/enOqj2gF/P
2Ll7kBQqz/tgSfHQQqcm35jWTWlUyJ+oY/KKzk44PaX1rzfABLZb7DPXZq5ulPLZ
GPak5FottWciRY30Iq0Byzfbl1C92wzUkvX9t8tXCQM1BAeJYjqwq5It/PL1ltOo
ooHRANpnO3Mbr0VabY4+PtkqVafFuF7Eof95qcQNrb1BBkC+/JPwML67lyM3dFrg
YZOYaxvPF2MMo3BImupdbiPT73ZeuAtYKsjZPv/Qw/6EBfYJYn7dYC4U9tL2A505
mfIc8hfCLL3cU43ueEOxmNlGRhhPPQcwiYE1ZXZfi6x8cyfhqHsO8HS2e6CuGyhC
bhoulMYxsndXVpLBYILwxVrtIhSUpyUTFcs4cVnuMQAkZGtTKMQ/vfsjJ2dh8er7
vdcv9HWoR71ClpNcoC1c4xdNgBkUuZHXBkVNEHJh6Y0vfoQcuJnNKHiNWY++qpTi
efeV3n/9B0o6TSKTjB+gShdOHU6N/nt4tDvuxycJb67oKWYNm/+n4K+kalJrrpNB
8peytQYgxgd0djl6q9UOKVul8lMHaEVzXtXvEN2AnXNAVDzVPyiDIM3An9tV0S1a
rTy7h0+aqWXcS6NXHdlUSYF6xrcXwjfNN3mEufqd/GXW/TgwCvdJY9dNg4KgIyrc
FdJWnrQ5Lc06mPGEBP45yk9DfaIYL0fIa/nrMoh8i/+2Y7bLT7E2bFPyEQDQRrX9
NSoUWlhmQSRexnSdBhi/TJpUwLPTRkZWkK2M1gavkneIK6MhNBwK0+yw7ss1j+Zl
A+ik6ecODMCCdEYZuc1QU7y/PcANMxOdXJ3jTzxkbK89M4+HmZfkvQ+Gf/LS4rdS
H+08hBJh8x/KhIzXJ0drf35la3986vlpyNi8SJK8rXdXPjbYgT8zetpcj3/P41+o
A3ci0lmPkwVp8yapdcgFHup2xK3hc4wRR7oQUCpJVzh0JAsedtauv0/zZ/I5BQuh
47hQbKs+qgYekIohcZexifNFc9WlSZhFsgyV7zDpxjC4fVvbvjoUe1rPP6FS2Xtv
Cz/EuiCBw5GOa9V16jEk8BMHuY+itphlEGCkv8A1+s0xRXxjbu+0bIEiYnmfQydb
JSTka5xgeT8y3CognFf3b2/j9YJX+QKixXfVN6emjFEXYnC2cldasdHXGLuYFRxl
owmyUNIXsucnl836+XiyfGkTOnw0++uVP9L9nAsqYvzN2Mt2F8yM+CMym8rTF+Bp
AuOaJ5aP/AUo7umyoV85PYr1UlT/gls8VU/OLraPhhuAgwoHp8PLOvCP8e5WO0Oz
86HODgabSeXFVdEbc5Jls2kRePs4ZG6FuSaVStd69WubYDy0vuEPX4GifsaWXsix
YB2UDj8mlLiyfKu6y/fmj+mHR+qalAD4eGvUMlo7oFKcpHis+a9NjkkNDKmR3Ae2
0zYh+Wzc28xrYELKDVpkrif1UspYV53C7HqQN3a56rJq28MCtMuAIn2SiGxOru87
eY8ybolHkcHMSlZ0+e2qN8Z/wPa1CP/UMYhfp4J52zZk+9JtnibO14RWW/2PwP1c
llmNfUpS2UnVMXaJX35w9Doujj0zMV6MiGD2+lazSj90mFNa5DevVxAxoN23hLwC
EPohP8PmPeaPA0PYW287sTAxWnAnhksM/4Z0gvLiF7bdpbOGD9zKqZFdYf54hNlj
DWkeudoLJX0zyHYPRhzPoKk3kiCBzQmV7hzRX/Vi67nxaYTEA5nIkJXCxyjsFj4V
0fhf3f4oh4gJh/imPT1InO74ep3aXTvzLg/7pRPDH7EiOGIHx5yaDtp03uxK/3qU
oI1f0ByIQ2xiOEy1zIBmgCKpO7Oz2rxl9trTkgeTIOYT4xb+0O+rakJ6SUZ6c+2L
CMOv9yhSMp4TVUGCh/QBGPwsJgu4yONYndlw2CcaaozoSiJgDX7dGERU0GZxHvrk
hR75W9OHPdcgzDv1DqqmwnYrERcqqeZE6FwfdgtWHmX4RDgr1De69iDW5NrkSgYJ
9X9bUoqLIfC38S1/YKtjCwQXSTn865zzyfKgd4n1Z7DjbZM46e/vOA6YDbwSX+tu
9pKYRkgf0u+7BGotafXBn32c0q0mxo8aMawHz2zQBDnaIstSdrMy6BmA3uAZM67x
6DagfDg9mKPK8+NIk8HuRHJPYOmw0lKoNo5EglCMlUEcN8ZwQDDpl4vcOr/AGQx5
CR8P+UVGo5v0v2Re7QXFIPQbH0axkK9JZ3tLE3bzQPEnlUlydWPb6VQ0Ns6+P5tH
Gxh1ZVg8U7eoAoJLQGzAEPsXX+e2oK49RpvSo7f6GlEXJ2m/d9Z5NBXRrZ8g4Sni
W1UI32XUnSpomDoy5yqEVs8TUkmVmFOmNe8Ynho7kEXS98dyEpI6a7R2dchajMWA
bBNhqdSlAMoRlTl15X5cXBH6AyNo6r+0F9uSUIDIg23hIgPIhZeH1lqzy9AnSPA+
iKnilWkpasBiNubMnatCqsG3rveJu0wDEvpip9SkwaSo+Os70j6RDFFADfPI3OsF
y9nZ5axLBz4i9mitjDvlDGnoL1SDoWGKBgyiXeDt4TSfbgpgleaFEbtv8+Z1xJtv
OgmOskACHoxAABY0drgL1A2V5+5KzyTJEiaT8rnQ48CAgFhIH/OzRSXAw2HbbnOM
s3hSPr0ZpE1RCRWc8yQjZAqk169P5zCs9mWzooEDC0f/QsUq6AkLuurJdHo3OBU9
Db8yC82xKzcBYUHh8nXpBz38eb7mTgNpepMWv11l+E2baiF7Mi5dJjboH7iGI/Vf
l1HPMRk9X8OJ5obMXyKUin2nzaHgRF5liPrVVoIJmwGQxnIUyx/FBDIwdYj8IBqt
+F47NtuD6nHxTB79wv+pwSCH3AGHr+5BHPV/JVp+ygx1Kv8VQbo95yG44n1eOFTO
07w06ikDqKZhskcFwLTGOa28bTUNFnh5/BJEhpuhpALIV+Fma7F6suvRXlmfSwuF
J64YRSpmp92061UkXtu8Layd4soxZFrD4GH7Ko27A/DD9xSNKfl5Ajna1jTAfNR7
B23m+a1uz0eRO5xj3rsPzJ5Wurk8MF0i6h2uGyL8JkvEsQ76Lvvj9TtMtO3e5fwa
MOohqAEVT83SunDzMhOTlviUKbPcjiXTeQF2afVvPqOyc4NmHXXKRq//fdIgQZWG
Ur9Lr820OTkUjRhCgqvtEXefvbOFY4sg3GDT34ivbmk+vF+6LMTO6JGvqAtkuqsU
Ey4olH5Aect/CYTK2sU4QBCrgikjwKWbwJSfDk6yT8INVckqCDnngg1caM/QBHT8
bYLxUtf4cddlRQKA/jaVS3vOYakkA+aPJd/lJLUD5V4X3gVSTL0QxkYeuikkBaWu
VXZPpfMnC0wMeHTuP4ebvfyoMWwuGJXT07B6lG2EdGQM4NbOeoKH3vsDjX1IHveO
KWsVWSFKHhQk1nC5Py97C7RXh1zXFzW0L1pwJPS2u+NJxOnDSSHy4DR5bVLIXwXv
Cslqk+Pln05hnMKDZbuClAgvsgJLQZnbuI774dzYPsJQRfsjYJLAEDo9uWQe/rLg
Xtx9H/Wkc9V4vClV6wg/bJ/VX79KyUxrdKjoOjoN1Ebt0OKxGYYuvoyPakuQP27E
vCMB+x2BNOSdV7yKtoLE4P3nXO2nLx78mK71a7voq0aVy6nGZjusYM3Lr7/QHxEX
hu2SHGlGYy2bUQKX++I6bBDMEpd0ECxvZ9yWyrCTavH8/eNrTrYTzzX2yJZuelR/
P2u+uE2gwECRlMQXtiRXQZHHvUxemoKyeg4El/KvpveHWLJPfVDdjkgtPfYtbGUE
g9uN0dTbN1AGCp5V6KHmHxq9tp63Aluq4RHLZu5O8OsLKXz6hSpikmjujh18JHoB
JHYL+gr7R4Uh28D5gIoOSg9jCbp1AGQJCAmsEp4WxqLFtLu47+t6KdHQ6UWDV5Vv
TqbUTPb76wFXSs3hWHol62fvIVJtc2xPDW707mLohPbuUO06dLaFEn3wZJZu09uE
PfHlvd1XYFzeU9xFDnQ2RAdx1A+LibszHS9Zue1PCynQ+j2iJZ9waYetan/595Xe
CL+rHsL9anwmei+F1vmXrC1FQTtK1KeNv6CVmQTdeMrQrYW6kJLnds7W9t/SuoIm
tGkh29PlYYygPnDK4CXMu1r4cZ96OKudghw0Vwf0ETUaCPXmpoEZ+dQrIH49VHs4
U2+Tjs5IzhmMuWr7rV1cqP/P/Sg3AeYhUsq0IlNAIPionmBGo4NlujwOaEPM8l8d
Lsh6cMv67annzCtH7gjqE/JE3tSBVTbHtuGigwri/qMM32CivB35TvXB//cv/YuK
qEdkTmw8W1c7tJ28ix2+Cso8pJcH5sxKfpI9zpt1lCT7fRquj9OdAGpbaNe9MkFC
OKhOElhhNRQF06EkaX3RNLzwsJJwTEbktENOyCDHBSmtwxhJlqT3iCHb38pDXFXH
z4Mm/EV1W1L+bo6CZnJqNeB642CnL1tCL5+/WSsXVsaVyXWWn6qkTTbkKeCdzOdc
yTQrNV6hle2nMd/ggsLjPGoVKH7Uj/ScgGVHyNVqlGF7CWP6wkkSyKTfpbHYhpNL
7RvVNbTUC1w1ytK+fZy3LHtERQHv/4kv//xG//5Sf5IlSFFBdchiTT9xAunSHJZd
jgqZy0Zg8Ra/Xq/9XUYeoVPjq0oCqvS0eiMgIDkJwJjMpvASACf7ZLM2gyeSvB1l
/IUrvRI9fJyBQquPssqdprZOHBZNUBs2MR+QZfSAONxR59+D8CjL0bmYNRncsE9c
1q1wMFpdMSd4WyXeJZ0w0QNfLjC8cTps5aZRyk45jZRNL680KVdVQkz0M0Cu9WKc
m18Hay9osqSUXlnfkFXVq7rM8+KBme5BQkLl/o+NEN8//XdPDTb8934nScEZwFSf
XiPJZMpouxSRcmvMWSI/l7dMMYtbfkz4L8L9VvbMu1uKpRQ+60neykp1kzOM0k4Q
AX/3xZpsYvh/aSgtLmDfoDovhW79rGqcSG+ClL0oNCPmALZLbmN+hKR4aoxsf+FL
bvtpwH8IKhnOk7y9V6yP7D/BmJgTKT6fMWx0BkOZ/hsU1ydtk8MixX5rBCBVMzJZ
pG+PXLbBZGtBodYndWgPnjUYTAArlY56HubLb6TJiF9V35+T8djPpMgoDoHzop4+
oDXKxICL6nNF0mFn53DxZ6rThDLCQwkmsqexRGvILb14wvkR7c4x6pBNZCL7CLpk
hQIDWmaMsN6AeRNGQ6mIkAkSxvZAc+l6P7ubB/RAa9ylCo9Pgb5XnZIRwS03QUki
D1sxXWZwVCpT2q3RbK1cfwLbOAH4gtxxulCP++BXICmrLoNe5+dLIE7Gq48LxQWS
vxTQJvtqIgvNYu3DDwcpfoWu1xnog4cXAey1mFrqdcm7IBvA6V4930RifNal5MzI
ZkHBC9iGgexkglMb0BPG1pqIENUTvPh2d0qbPiY7uSxdKwrQ7DTjQWGyBfPVMNMf
PUdP2ra112/9JCUKIWui/uL/qWREhxvtCEfJD6EmBl5PL17Uag/9KA2Oz4YlkEQM
esxFiijTjqwaKxtGlFK3EcUGQQwLL9D3s0CDL/dg5UtVS+td+RlTyoYXpZmuJkbg
04GUFsGIDvV9YpKw06UWyjcElcg8WU0njxOFGm2E/kxOt5iuVke1FkW8h1d/XBpw
YOk4tDm+y3kboZ/OzddtUyOTuqYSOptUO32jh4GBhGh9NRryLjqGE8rdD/w204Bz
72fnqKrXza/290VZOubyTlDfWiBGrmJ97ekoRF4wfGs/2JiSXRMcW9ouMSFxlNPJ
mPdAfPUts2YaiqZL9uQjnhKKhNBGAwaM9/hf07JVGWweLSiLNrTm0JJ77CcqUTdG
icDnzhoMFi0jhyACgvFBB4FfpVgrqWyYCJ6GOjxDcG1HpWIVLZQS5vwsDTiUFcz0
A9V/JW6UcEkpWv7ZKmDC3/9XSztXiOKSVgjDX2Hv0m4R/vEem7d5Ix8k/LtRORku
g76xXruKcMHo3eQg7dfOVR/hspWtK6HialsBZjCOy/8Y00WaKixrthsb0429jXSy
3dq32hoBZPLja6T2tGJ9Kaw68ow63xFJ1BsHvVB1NT0Q5gfepVS+xZOtkzLKSet5
sU3solG+Er5ojeCBpEJ7eyAc+5gRAMfCr2HkQ6rDJKuipeCl7gbCAbknTk/BRGJJ
sMRIM6alLZ5BxzEfpECmGNs1HDZv63zr3NzfET7wiKw0O9tawHT/lo7lk/pQLj9h
T66uvQQjqNBM9Hffh69Js4oIV2JSrWx8V3femvSqRtYYMJ3xYJGDRRyLPeXSbUJm
5tFZDMV739LeP1e02krUJPWcN/IxGW4Q6XaRMEyL+3VpgmwHkituziHv+E6cJqPq
Ex7/Qd+qDLKYfO0+DkzhwB0cijJ8I7ZzbvP61djdZkwyHmMJ/c0byWIxwyscypH7
KPopUpzLl3VPLjvEybjctBMN/w8XRZ/YaxsfP8Z8Tzgwao2KO/dphgKkHiJH2yUr
iVqVcKB7uWoZ4MreFs8uTBGe4Fm4FjWC1GnvTUIIRFTZJ/wsp8RekdCMD27ybuDf
h4HNm0Fg28/xsOyM4pcun4hkkq9DykkmliMYAosLj87iiTqbxocQ78kIbSfEkP7m
RjD2e8JGPAd5HroHljqJtkwuQBak219EJFX/ffXZE8MPsejXJg8U3aTd+/MmTNKJ
VhhzeN8bssVFBm1saotb5yHWUHxWS+NwlUHtpGUuoJwU+E+3pCVbXnUJizd4rRr0
JW3aJ+XpXKbN00KOaSbarKssUKcQ/INzrXnQTDmXRR2dBEtxyxA3MArKgF/d2mr5
kaPa7fC+x7MKDrDLc2r3o07z1znezRluNmSmyxzpiY7E/whOr8lcgulfypFfFXue
pq+XfHTfWvxxNEOkXHIiEY998fzxoThbfBQnGm/pFrJ9hvv4fwfscWa+lXz3k2hz
4Tdg4gaDMdh8EelJ5S17kqCSqTpvnOe8h5nfRMKd2Pnkg6m1uw8olio+c6hksS3E
RVEZwNI59tjgSedfXPsI4gtBFP/VAsnbx0tmM8fkCf4qNdmT+U+2s8MBr91a4szX
bvW4ExTmJcV/rH0HVFhy4SMaQT+y7eqOjcGPAWJXO6NP3d8buKLRjl8bG4HKzQWG
T4+bzp9mE3+oAd0aZew5JBzkw9/qPLhchbFmz/J0qi6ZCgeBsHcszOTmMUaaZwsV
YF2ixTlnCg+5AlNl3Sv3S491X0GzvIukZnQYdwQLD1lSZ1VblJecpW1Y3koGLdaG
gKChgmNRHXwbBWt8WYGmdAcqtqe/z58eeQtiU+IMP+Q4vA6/Weev4a+znj0LLW3X
fcyldZuUzPAX2ZATs4F7b9jOStyZuDiivbE46u5hBNcHHxGq6Pz5xxsV2/5QFLbd
i30Bb9UtyssM3REdVOYwP3HIKsn5kIBsUahaMdZLI2QPbu7pNB6FIOCtxbBoZwo2
gtYjZA9z3DEuJSB6oKDRJlU7vtDWXHfTxOGMRIoB7zW6muL3j97wD2RUZ5LpA38D
2NJXlPxhykJjohaoUoUG2SFetBULw8WXnxTL/X5nX9w3DM8GM+wljE283C1VDot9
kcvICqEqQ6Xu/QeJ/+RwLIvCWnhPXWBHZjoVJRg2VDg1k4DQ6IqO8pK+e9Nogf79
nWiQe3F6FRjHuKKDHRE4xcEtbddwUt5djp/eTfAgbHRpxJ8rzvX5/MtN7zu3ICdD
Crl96yOJTa0vcj6XutqMIAHCYhrxUnQGvkMhC9xCDKmvmbX5dGJYNrXTUof7+5GV
kDgYnxroEnmw+VYAXoTvdu/g5pxordrAsqk4wGR6ho4I+M42kCBhFPPNyIPEbII6
UGh8kJOmZL4lc7eOIuRQ9EzC7r+fys/Ijggpp+ZLozj6hmf3TCZxhqJ6PhvK/ijs
++0VI+eQwE6e4xCrFTeMC7hSWIXdq4ly5hTVivi/ZVzNTTfSmS3fvuVOVEn1EbPu
doqrJ2pvpC78icscwvf2s2hDGKMTa9D5ZoAMk4v7kmGRq2Zsk0M9LFOxWu5zpo9V
JtBunW0v33/5U/N4d4joroXumdLQqcrJS3BLDtfEKMaWvIN+j8Ki9zDBT/mJY5/T
hdZly5kXUB42XZtrEXzwXXQLaMFZbUWGQlSR6U+prd8Z9z4aVRULHQQIJv/X6XGg
Vym9vqFaXf1ekrm4qFtQbQgyHgsg0Z91YFEBqWiCPsc+4KIMgwgw7OvgUstnIkVj
oGh6zcZK50eKP0MgoxHQrOhT4oZnkxZHiwY/uGTQTIxpsas4/RZqM383NECxSX5Q
9b9vzGVEV9nRMDNVaH++XXea1ZORHaRZvs5nJtLhWhvoqNySsvNwm8v7laAlvHmM
8ecVy2tDnP6wQFVs3DxBdxzBfdGsSctnKF7aHw38xaQi7OxCzwX6clCY7iyGqqeS
Vy6mdjdNGGgdqWvLS5Q/jY91EKlm1y5P4s/cFq1lL+7I4Uy6jpqZIrmrQai33aFM
L6VUI/HrFYt9rJEr+VlWVbG2tBDYcgwZAsp/vWQvWbTPPhx83NUiAN1V58CmKjd4
MkBzpfTmBEYjo+BLuFVX1Ep4i/iQK98mR6cRhAwHjEvw88XFKbwKuzlRMRxbem8+
ofUdlUDwY5P+7KW077IIdZPXY4BRqpr1KdTWZxmt/wS24YorMpmifrgtSYN1KJwG
UfP7UFPe7maecp7hhJGsphJo8uPh6oD52gW/yd964xiRPrrIN7BrNKjD2dxm7kgq
pZ2ckWHsGVp44cIH1hKuIj+HT6J7Zs51iA9wzc6jPeXD/98/MRQwjdBGOdDiEhlq
vjZCI15RzDG/FQ4Utwdc4DPobSK+0+nF2CArSTs01Iq7M5RlS+m/qPrJfwu51M2a
v9cHiFpeqxVKT9rnUYaQCZpTFOTT3RgF665iJXbX5y4BZF597WEz/Ialy28Ic/qV
ViWF0b4ayYF9EAkIFtqxHXx0AKuuEBB9xlfrKyDX2dnM76KWrm9eWsyR7GMo8nMx
GYb+WiChCJQ3+Hz3iHUfzkQmMiR6PvHtaPNTmV7YcF8gZ8dHYRu227CubYtN9nK+
s0Yx1fvvTrAjaGJqDhBkk3nMRwl+s1APsnoWfz7pdqXEZE2OSf77ekTivAUA7XR3
lQVaSjQ4fz4r4rbdBObMHyukjdW9fGbQX8tYGBYHzzHlM5Zz8N0xJrwUrARRhQ+a
aJCWWLGA4o1VV4mt7eBJv+hRjeaobSeDewQ771aoX7gxTDRtuoHLGxo0/Rbk4KYc
G40zsFdM1pIrRutpwBrUhm+LhuFwaXMxZM5ebHpao7Yo2DqyEqwGHMeCal4Ndz5B
2K1E0Zatr4Wt6Fr2t2PtTO1BlvG+Z010ljhwqhJvEgZtUh3a5SyN9WtgYl/MioIu
IrwzJW1iPE0dgFrpJdKeewi0eeHUC7HCznGzPvd9ivqnwLQyrBE4NBnh2sEHhzRz
4JKHMUjzRTYMWFrpvGcKio4RFC8eNYmNyJJB+soX2ToSEfeEoPYOCL23sPj0lUg2
vcXv81sahLL+ZhlosIYtV4fQiQf7z4fZtSZQX/ki4OKjiQJvJ8xi7n/VtSDtTyBH
PnYVJOeewX4hVGvGW7VTv45cJbnzIR5IxEt+ATAcIVx0MOjGho2XOGONNspSkdPd
eI8q91XZ5tc9XTHH+hQkRK/+hVNc0qPU4f8U51AWaenxJRkFTPPsnDZU+U+SBCo8
ugMasBqGTv/CoJxmieoH/g89oV1OcUm03jinjaefDRyHYIfUb6av8E0D3KmxBkUD
bBmPvefEv191uKDofH8tMhxdEVb8mUd5ducxIwAVQRiSP3oeAHVCYXRAwP3KNlcg
sThopYkSHdFGMJlv/5NisoYrwu1VJXXuqDQrhGmRgAqIzisGpCzHKVSiIMHjIQ4W
/EvswWFv7UI4Prhll/S0HEVLfZt2w/VnHSum74VoGeN2fWQUKHFSiJV7y6xinwCn
/0fnAAZRrwTTpE6OGjz6wX5Q0zNFx9dX8AdhLzw5h3YeropF2oxTmed80urUzQoa
gCGUyYPsArbB+CHhv0sAa7g+jSqYclJiEXSA0Swe0Rc5q2Hc4/QMCxdySOZwQAzu
rCm2rXuSYGF4PwA+InPEjCqxJ8vApnuOmUW81OuHTrzpc2EGX0MwOGGcDA0qPIxd
T+/zrDdzBwPogV814XxJD6TBgKetGQxTawFfDWqIzdfbZwGcMHTSJkVnJnTn5K7m
Z7a8vXWwKJxN8OQBJPvWXYPYg8AOkMb5L/h2wGaucEnW6TCBpLY3cnb0HwUgj901
JU6dEt1M3In7AzsggrHSKhrwJ16Ci0NrjL2K1ZtuCqjN83qYjESAz0n4yumz7Z4f
6B80nVZ3IxZ73ahWHimONugT6AB3HnFPVKuFuLpTOd8JdNEqhUj3mWbGatBfmhBi
qRQ3JPSZlKB5iGkkEn/xvruO3yLW5JtReTgSJDpTcnBl4CLmkBYPkPXZYSzE0FFb
S1MI6EH/T/NR2bLnEmpRPUrOw9I0/tsI6xI6+b0WY9eK6jswrknpStNu0TxQ5ii7
bzo68hvT0gVBwy67MJZkqphWwKNQhvpyuHFIiIW4G9/WRp0+9YyfFykbaZ4B5R0O
wH63T7JAK+PbSts3gT5u/WhqA+Gc37ZH3h0CAZ+QfqW2C9prh+pxGxOJeVNHRCVx
0Tslh8XWCJxXDxPf0xIS0nNCZV4T59lRjA4oNos+zQDsesbTz8UJ4EJPmwvEXBw0
YWkuaKfED4a0o1mvxSGoHUhVnNYRufRrN1LnWn94rjFFqx0brBMNi0gFmPQz2a0r
dtJcyTrYLChGFx1uRxZjlueCizgzRBzUY0lOiJl2/6RTFpTqw+hO19ZMSmh+f2pS
+AVrcnyc3suI/B22WT1cDYpBdTW8bOhCABYoDKMVaSBxV0IclwWBsz4ng6Ah3CGM
dTEQUydmzVzEDT5SNt7C04jQVqiYArrkh/E3Ji+NNLWcvXGMxcRghCOmxjnykbTP
e6ELo8Yelbud1HMctMEY/d5v8lop9loQ17BewXkVdIm0YyYUw65ilTIJC4GH08En
0U/tQar6Gv73uc+OrW4DfbdrkDkM4V7L5C6SruYUJyPEP6sH+b/yFVmdN3Ywtdog
EFR0b9U0KIHf7nF/uFdn+wfGr/NPXRKK4iyDv794Ytm3MOEX8CNVVENRt4ezFP3K
5BY5Hcomk3mebcDXUtY6PyS4Fr48/8rUNkZJAOPBdnwbkgvm4HZ12kvkhQXwRe4c
8gUDVQK+GkcfqaaAVmIG1qWlQlnnYVN6i25IDoVqbZDYZDtzoANW3EmWJYuro/bc
jxSDg38wuhZwD9Dc6+xBKtT6FnIQUi0ARerJiJpXIB7Vg3QYx74v3AiS3Urfmmxs
HQ0fBVSg8/f7pA1GsCphacIScMvebv3gt9efjtdY1gOGN3L+KBxMmQsPmTXbmOob
yTzdtO4oMOFjaEBdPX4yWuhaJb7m/TXACQXTTc/o9/GQsmh+TcZJMkfYKbbUdBZC
qfJpcy21k7OWkznXDTLWUSCr/3gIkZWs0Kd+J5g6ZdbfAsIwiHQGZKeo6gxX13qV
sPO8FlzEERlso4/f9stFcInh37pAOJoyL0fmYAVJiKxyP8GRW9djj/AwSyc6d+IC
hqlgnzuZwDdiraaWqVnQfO9fmH7fd8LgvfOfXc0X/Gcm6Gv1kaU1EQBPzvMMFnms
g7OLGKNJ+CZhciCimzCyQbwYwxUtyAQLM8MDY1CZXlqD18MJYL1xKpha8dT8WSBH
j+wlPxQvoz0lY/OYXIuqA3Jg0t/0SMlcI7o3zHMMKhBNmbf6TQH3pKYk4GDijbTl
YSLlI5WXo1cPp4pV22SilVF0dJyfp5NtIsSPVQJ+gu+E53xq//FzKF5EuzB4+WQZ
nWBqHRR1cchtqsQVO6HNGl0fy4t0a0PM+26E8d6t101jc0YfoypcAerdsQDISg5Q
IXUNvwltH3Rwot99hy0cH3jPZj0LlRTUZwFaWCss6ZhK5wsnwu7PqQWkCLXdymbk
RXIOtEqO+yyjFzy4YxE266vCNlunc1lOg+t8Y0/7nw2aT7BkGrTsLyJP2TdVFWAc
UsjKn+ttAOa9P5KTyj0LlKviaef2uquukRURhDieH2h0FY7aVQsK5FtoBDvDsqtQ
6AX8L6t8Gl1EVUqFhFLaOEAErmFznpUx4P1+eUNgMWpKaxVVoVj53VzsrtU0FwdR
sCv4AY4Q2lzl7vHBR6Jeu/Pl9b7foL2NB3EfWTAwFexzJqmfKFS7cAEz5ztq45us
eh0C/M6ukJtxImP3VccHLfuu9IepQgzGNd+7+wffmb+8siVo0tVVAlduxombyKOL
NE+KACSrAGpTLjRHpD34ohfMUdC8TCg+acKeTq88Mx107yo5pjakm7JKEILjtH2v
oyR53EjbFlbzrmmf4LIAeoDXSDtFmNZI1SJDc/484x1ow/wSUbDYqu9iFvlv0SJ3
KDqENK1fcogsOwNcyp5ghEJ/4+MgzSTxr0uB5T+7MFh92LDcdW0a1hnjLH/sRLD1
hhhxRGLmh0z03/HPxK/JpHRmgvUIJdl1I4v/QB6LbB5BrNo1Acq4Es89GUNYh3fh
zauZAkfzhCJu8akO8E5gEMWAwsAgl/kW0KniSDx/jY8JvmLQvRHFV/iD4E4opSfS
061g5jNpo91auIOOVgEQjbAgGomp6x0y9dHHGTV79K/ihexNL7gG5oAhqEREhZph
B5P2MHIxJk2HXawJU1X/lsBgFfP/90gzCvnIhxF8rY2n3xqRMblVmK1Q+/a7k27Q
ILK77hUIAQU5ZfOHe8nMjQ6ytpcNQeDQgkypoRreW8h3d+yHxak8pkXnArC3CkDC
42ae97a+4oG8Fs/xeA9uJDMaiLUcsHGBlxSEw8aK8KJM3lyUKSM+T2VdQrpgFYmR
ATyta3cIhEFWVA90WvZcaFptLI18tc4irCZ18jf5hw9jRXwJTKQcoPSzBotETg1J
8OZ396iBO5jcPqDZUzqKZDuF1tI9RAFN9yYgTe8bbjDtmTuRofF2aGSLhxVvtVCv
1CUwF9isJjW8ZTHjCR27vbJ3n7KkbXCw23/Of5owpO4rWiatcqSGiKCNCGbIhrG9
3GlIZ6Z0brdIKrOnEykNvJzb9WgbRJ5GVASVfHlQ9zR7CrJ2YBtlSmGV1U+XwG5u
GvA2AHEK+xbTu93hNRHVU/0Q5KSyafBUjbJLWeYYC9dgHTzE3xnDU5pDllNs4mo0
9yfUchoDk0OWU+sl6MFMmrrLZ2HBCV3g8/MzMQR5ct29KpPlPBhYxHONPIvhsy5E
O9lgjrfl0DTLW45Q93FsOYu49pIWelPY/kXXqzJR3HzeQigtBum/YS+ZJNGyuvJ9
cX4KKBpvnJgTA8xrsj4ZKY+u8oQlgCi+7JJF7hJwnPl1K6G3/OzJ7eg1n3zCg8qS
dXcp9m6+rMUnRWj8osg+gG0v9US0Kt6vH/fcLQb4X2QrwM7BjOeGW8/C2tF8zX7U
3fBctkULWb6cp5CCkUH5rvu8mrL5WkaBhYGFdp2sqOY6wca9v1StIeujIMa0HeaK
QQ9CS3R0RpqvfkzsIG0HcGHi01zXRY9iZMcBXNW6d4gKeciKKNTu+kBOXxNip8tx
BYRybOqaAXywQtUhtuI8mrH81O6QlcTlADUl14Tad0FfbMkyOUz5AHEaT/asEwk3
sGKkmATLRTinbd7EL5OeRjVdIksXsxgFLgvQSxDo5Tl3tJiPAYC8RDOOboVctXyO
tNyYQB2jJrX8xidAUZqvN11I+aUGtQqBYiI6YtLPlQ7wKAfcR0I8TKGu8GsjrwP1
uFFnK0uYZzx53J9Q3N3AkrQVDJMZWY1Lz7Etn74H//nXfV4UBFHFgIJ9cmsS83Rs
pZv+2cmtl6+ndLB7Lqv3qdqqFWjV9Xn0au4TkpuevVK7SnjY2jq/sRHa8DUrhvVp
qxOBnLxPeh0IS3+G00fMZWTnB+OsfM2uTLHZh6N8kklTkh/ZDes4xilXiukDG64a
/R1ae8Sr6oQHBedpaaL9auKdjvOdBxT3D69/+D+0moe9BmcUhdyOdqhkzsQXNbi+
wssktB8Qc4mDD0oHw3qqdeAEeZEsmoKZn6MdxBBQLALB8fTpdJ4w017uZs5NG/wz
1349n+AmqaCh/yJAwYns3O8yPVeUlSL88tgAr1GxaoT4vG294VZ5gO3zPqmQi91M
Jaai3bVYsIBaJe1s+TzNbUCXJQ7NcBqXblYa92wcvBJRMdmJcozIvb22iBbgwnMj
3OSi+hkLTpIpg//Pm1Mv987nje5+nP1mD33p3/uCrAxcGSzIw4N83mqvD39ViYlV
qcEaib6H7Vxjb6UBkc04n8QSVNBTI5/eUrZy8zWxHmfKI25g7juadEkTQeQR4XcB
y/ug/L/rBp4QROIeyv2N1HwpvNBkjPYh1BOnT0R5XkM+84nk9rRdtCKgElOUxCWo
8oyNw0fuYSv6bAWFNapPXtI6n4Re/9EMDVD/9xrGCExHWnu6DclLXUjxujcSF2Uw
pawfRyFsCcLrzUqXE5GrBJdXZp34orTbNcfaKHRPl31rDwWP3FztGcRs3h7Fh1te
ce7O0zjNCUqnpuHgH2sTe+SsHpL2FhJPRyn1Rhe8pCxDqpOY8+Yoxk8cYd0Uiu2f
FrPG+1EvOVh4Dp26U+bP5MDoot6DFTzVWGEh55s1DlhkiqbglVQjpJ98oLTIRiaD
42uUQmlrjxCM8snOQMqnrpyaKAhTi2fgaAvSAvmWfvwgvIAwky/tTiZ/mqkTD0bc
FOMzioK0m9jTR+gEuBbWMo9wIZnlOBE5Gb8WecdrUYXJvTWHUyO1I4t6BTLJBLO1
pdW6o4RV1FuSzjaIjFALulMNTrh/EhspmKgGHToXldde32BlL0GMLTMVFPUI/ZCu
l7iN82jSEqMrdsIe0PEtnn1AYDd3oCanBKjPiykGibJ+TSlLyybZ8tjMjX254P8y
CG/7xAhdKAxRR1SF76dterV7W587z23tHlMd3BhQowESy/V41PrSZJj3dq6po86D
p6tL58bLKAQN19qPawHZsd8LshdPLxvpZ9iJWI4BjOjqRTW5OiaCTwHtmpxeIQ9r
VwfI+yUtC45LBIKzTD5aMO8igk1+PyiyLVHJ5AFJYjcLSxmhAodkE/Z8MYP7+XSZ
LP1xmXmfBZe0OG3Ne6HKSjmaKmtlSnDtT9yzQ/90w34/GPHMUSUCV534JJAZF7Od
jGGcCV+/0SP1fNxb9/qU7wcRr9S9OlevM++I7HAabFTrp1cbUyoFlv3Lv9EAmaVZ
xkOeX7+ojleKR2rtIUQZQPMEwZb+heR0jaAfCHEMLSlCUfx0RW6lemgus+FS8hyI
kLFmJi1kkFk5A18GUp46sPzDOSSR+hn5T28YLKkTsbDPpznMJx9ub0L5B/G10JAF
3/VJ18585qkWon2BPEuOVSIrSaUJcbkmkYEiTZqhBIcKqzA8vutg2RsmyoGbNcaI
slzW5CBGZcMSGXYwgiakUnzQIp+oQwKOdTqCXFX47Vx3DeN7R0fNSEgbyWz5anpd
LXvBi+7eHj7qvPI8glwXbzxa6lrhqZZX1QQRgLbosSFzfZlHv6Sc4iEhO4YenKTe
TmPCjlJig4alcGiFzzZ9uQtEhmlTmL7/CbBM3L3QjGGenVa05dqE8efuMR7vO1wK
QZ3DYmj7tCg96JHy0yJJTbnhpoOdMFHz9LrxJJ0gkkCBkXhLBMpTJgbbrZn/MGx3
E9s9tOdhj2sDVOkaiIPGRO+jeA7S0P1lqqmR/aFPcozQ3i0Rwj7Tblj7Um7RwPkw
zsPhvDP1A5OCyyxAAAXR8+mFWXnsqyYImbLWmakVxC0HbjZeBL9VtNFD7Q3IyFgg
Pm7xRUHbst42QGd15Jjx1Tolg1wAaSiDZrhelCc+cp6G0OP2kxfz02pMdmzDTqCB
AIAtrsGmX1gp1DwcXeRJFgLgnz+z8LrKAlNxMflw+h/MEMJEK2aQjk3wvnm+/uNO
PFmr/vc4GOcnXNJUmMdyl3/XASdTYo9oXF/RxPHw3RzOI7MSGyuU0hG+KqXNziDJ
bwHaOSg5Nlgj7/lPqUA1x3Oo4J2H0B+WiEJzEgedClrKW+rHSsLOnfOZmdkNFkjn
nVwnrBBYyQzxg9qyGu8hjkWkmwwhGOD6Ze22b8CVWTAVc3Lv9hrPd6s0a4xQaS9e
tAf6S1QSuW55K0lr1/nZV36C+KjQyuN6pCPEyobRPoCOs2lWKO3f2uqEaUt1qx6x
wCsmRMDE/mLwQVe6VDqe/GgUvQ3+E9GbnfmuUpblb4ZZnelRce3MYmZ851/U+TY1
DVttNiOi9/+CX+2eP+ZY4K9duqCfGvj98UflmCU/sig4moxlM+aZrdNDejq6+vxK
id0as2dOa9eD1nkWiARpVE/Tdtde1nIs9/+0Ym1pJnzixVbJfLYP1HH5OwgfLZ8o
PyT5cYcj8N6ifHX/t9YldlKoO9mOuSNHpvYcFvuzZfg1lVLniQm72ZE2l6hqZpAV
XtjQWlneqbLjoLmFCXPuJfZJPPEFWFFVlTDcBP1hO2abNzPRb2pDaFzWgLeKGmGp
ZoyFYbER3HTJQF6oEnh0OIBlhaZNr8D6Uk4V5dCuJWYU5Q5V1LQB9entCgyiJ1jh
zU4waJEIAjAksIhvxppoKpHs9zEmFCMhQQl/NpCOnab972BN6AG8J/RM+M5VCVb7
/j1B5y4UjvcH6SD7LjnYmIvhSvgYMT+dRJZHEjmRyCgsz7cPwDQwhsQQeAPdy8Om
/y290jgQeDQ+P709fZBmMoYw1Ez59nlngxHnaUxb7Lgq43usF2oCvFyFxmxubTlO
BMRIcgsm15tik44iuxXmJ8lcv351vu1jzov8hvcUi3rIntGDIeOBL8r9yxEonxx5
254Yw5yVj5wJ+S45RgER8GC4pGSYSSlZwMFZjVn3YQjZUpOiQP81hxgkLuN9dpuK
Bj3yfcfSnuHDo6ABlICSPbw0Sr/d4IgHqSvZ0C1/78GT4buOUKWwejHO5bqdvZ8y
dYrj/fQsBXsGHvpd9ZVNq8XYqFPo95tIJUBdhm9G3avnwUWQaddgQWQKIKaPtMdC
UxNllDj6ZiwW+8Vm9LHmYhaBgZtCwpsC1VOm4qx7TQsmnZgLxY7G4ZWHGlxbcH3i
637mO99PAjSyzCexiytCt9eBDSrmbwpkW+ckUIKRAJXAfbG6g26crYq3YORiuNuQ
yDahZb1fqZLBxh8qxwdhzgXGtzp1J9Xkc2J8X1etgRFJ7wqpqnwtTQsOJoeZDz+O
/jJb2idhQNs2nXo3tE+KjA+3UNz4rYQfGI9r6njAGaGQiv9K3aaFsgB4xL55dRyP
Qd6gti7KkMVPbazewAKKU/2+oH9H8jY4lQFF8PFAc3HdUlP1+2FER6TJy8wMLf+8
3/QGaVFEWosroDv2AMslTGvI9N3Q/eCDf5xDRkum2qm8NzcAfOkyxLbv6T7euM3K
f6rnByOjo8MJeFOojdylfM2XzO2YpChe+zOGNeClknQCxia3Okl4uJqMeG3vlWMR
ziH0sltP6uuGw5S/OoN7ogjn1yVhkOhDIbmrDjnihqiUbotaG/x/YM5A7drdLNr0
q6eJ1eIbSJE4BpBeoUWyMxoYebYsI/0FZzA194HeUvWIN8zPpxkjhRXYNqW3hU1N
P/sIlYBpE3fM1QFPtSEmNrfEe+sinzyfrtCu7ksgKe4uN5mbWEhfARAb/1w0antx
sOogq21S6Hqf6LjKXH4au9eq57zy0t/QQ89ozQglSqicsoQo5LDwc37tVqoz+r7v
eYtX0N0siXEOCxjmvWUNsCfJJaBxyqhKYgVSkU67BD2xDnj/vsQBSx7ZixcfMNlR
EJJeaZh0yDUGmZJoaBP+qbWKL6sHhU/khUHPJKnEmWiiVPkd7o1zuZy8chSQwZTp
Hl8jjjNwJKTropxmu5jDzwQHawTODp7PwYLH5NbhWyqV7uIzEQ4rVDWBbdnWmTxM
IdWWEL83fWTCeZlgaNXn5LjFT7+XqSwfWCeXhjbVL5/2+dcdgg6tRPpDqeRjJmS1
IrAjQBNTuiWRlRUNfyAYj9NLKyJTWtrm4Bwl1hb5sGtevP8AbcGtGnIRC4gHV8Gd
cycqDuh910itFHkn2kLEXxXlnTHTKPcHoiR4Mx/ler8kvgO3yn/r9sj/AENvCLVx
ODFITF8K699sf24xuaWTPQ6VhSYHe4ScHZuNNTFFfbIAz/IN/4IrT0o9dMqOyYMT
ghoa/nvJSJE/S0L3XtPM5mmDuCJkyuamLXLvXB0AFtBvPs+flAwwS5t4rFo86zhM
zHGg/UP151cPHUTbZQnAbpH1tAcR5XZARfdZnW10GWI5J1TQcVBNAYRLDlpcB8Wx
zf7e+RJAOEdkLBq6NZbavNJHJU/3r0Si+px3cNaX9j4l2LlJ9HFWTIV7efj7XpBq
yfRRjtpWQYButH1fzdENpC2n11IH/9uAE2ixXDW6dn0kzeg14tb0WFLIqLSX3Khs
Oqro9yvAwe5sL3zR30JoAXq6utlcOn2cf0XByBxNDKHAcrLpO0WIsS4355jfIeSP
t6JXPl7rd6WVfFlBpSmLCrc4X2SB3F6enUt8AA3DWUtLcLH+amiYGVuYgMYAP2m+
hpq979UP6J0j53UC65vj4NzNLm4AfLeb1Phi4vhnBG1uCFxZNQhLMLxCYaw8VgEZ
T/frdZqqzUNXXLgR2vM66gBnn7ihoAmrOOFAdOE209l7qpqL8cb+NmWppxxV/v55
5K1DZwHbcUsaxYhHU33o9hcrsoDORgI7OmmH9umeCZHfQma3SkIUUzhotV7r5+1g
VfRjbWkAtpYViVR1FbQPifN2ATP7asbuHruB64FK0qq8zQceM93ETOr7mkTXldZa
gey9YtKH/s+qqOZ5X9kaciWnQpwkJySFXJD64lBUrzllqz6mvCjpraUNQut02c/b
mu4ypGd9Zyp1NFbB5bze7lxvlGhYw7d2glL5OQ2dnjkFxv9JZ6y5GTZeE1CSneNM
Jcz6B+us2l8D/8AbfMZnD4hNlD1amyW5/9nOobjtZ9/0DtSXc4WLISM3m5sSGqtA
gPKRwwVOSGl0S0ssC+KCcftC4R5Lm3gqKHdoC55vzxZhxJdsu6XPWmzOHft49K4Q
ZzvuxqQdPZVA2552gqjaotbycHcUKVmlUBadnnr+W/ZxK3fUM2lPYOMEZ1bD1EAP
0RYWCHUA0ffnF8dN3jMrNL8IAau8KWfOLRLM3Dtfv2u0ChEnkL9DkqRO+j0YICae
0bNh9v4Zmlg+X4MGk3lUB0gip1BpGPyVBLFRdI6LA4x2+qtCrLJH+ohZ/CJ6F+VV
WcVJUBjnDYSQJTe4AeEIZvpk+eM+ZQaVjqdgsjDGGae6ueIwzx+mnJ4XX2z3qmvx
Hd0c3el1QNH2G3E7ZaZ9sE6VWEzjVZwA+Hxp02nshwYkUkIoSopWjs+o0HiLFA88
OO0VNBKAksDu9iPSwnjaFDDBk3j1olkOPhC0a/WitTPDRiFs4hS3qePAhzOkOmAJ
9OnS5gAduamZlbvYBeZXCfJ57kJsWAl0ZWw9Um29s+aCcMLaIiow4Q/bHMMLIs8u
Ela6oxL3dIX1IdUT3q2MZIHvWEpJyfMV+pzUeFuccN4f8nzTkM0J06KLbTXhr+fe
HtJ/08b0l6xCDX7pp4H5e73XT5+glNoVmxOghwzzd/vHHbTjgYNQXNer1tLf4CJC
xxHP9gLm4nU7LPEuOlcAszM7nH2+EndBmefOpiZQngGWp++Yy9gUUs32lOWVJ3fo
fpHfT2r0SQQ2V8PTEDjZug2dMnhTmnOcIuXsvhKiKZr1MX2rnhx+EgdhsdQ7NG7n
hyAhTjhEmq4tk+WDCGUwLjcgmsv0ZDCjbaRJIRIOX76vD/Kf3AzG/fE4kP8AMdrY
sk4oNaETYxIeMEQ6tXTJYzPW1kN/49u1dc4WRLVFI15ecfMoyDN0v1rfhGP7nUln
5plRHR1uunXAjrRkdKwU3EWquBNlqhP1nFlTKluGjxKFNI52vdhJVsRBwByNe0x0
vX3DuiXL3l/DvN683HpAbI8EH6c9OzJDviWlQ28Pz0r0OefdOjN9UGEXLmumyytG
zWwIqRaFUbuZnuAwXqoDWguc8HrLKymuLpskWxFcitwgnmJZvxhbIeargyQWYz9r
RRPxTdoBAOvw7ih9JXABH/lhcfGaByrqlB9JM1nNuB71ukv36d2vGm9pDsTOL4Fb
B81u5CSfIqzMf4MmNS2fDkB2G8TRbA1cLl4GDVE+yRA1dkzixIhaJK0KB0thwg6g
dw08s+tRW3MM23w02UhrniDIcIxAAbyN4Ew04y9IIWE+NxhhYXzyFzwKaoZIaX0D
LV0M+F+QssguWgvITGo9Fu2MFUVTvvI2o0mOPkFX09h5EN2p6rAnvCzBDDADbiYZ
tv387sFXwka4CuWJlNDssfr2jd3bVlufLdbpnx7TDAwUKqnVJBnW77ctxPYDS1ls
MWMgIiiVDxGxXX+5heToC5MlcEjfB4l/lZwqM6CYu2utJnaISLGVtjj+D1PPcflW
UPiXvXEcIL9cSe1gNCpZheSQT+dSLLaiPvMnyp0qJ4kH91BrKC69WAU39h2GZKVk
krvktKdK70M+L1e1Z83kTl29WZTDb0g45qIaoMhHD11oegG5/5abr11IOSsyQqln
dFU43MvJ59Y13IBgCED5AAXHRkq0yk91x0trLzi4qok8tHCPcrQpjZV8ZECbApPO
YXMAcVOBHsWg48rA562bRU8nKsDXyFiW46XwTK+nzJDLAiZdOEzy9Wl2h/9M+WKU
q87AiqmKplqxL5dcRLIw7d6I/092mf+pD9+z8fnxi/c6EsJA2XsfC6YC74WCwfu/
HLc8FhHQpikk5jgCiNNllh4KdXlVHoR1JR0Lm6W9iLmDm+yL90wxoqnPPW1VaL90
tuLw/ArYtFuLOiMu65nBL0brexlK3z2tImBwyDqaVo5iprUYZnDt5iLGcmiSP003
NErcOakVT+td0WaFdgkDIumJci2UBNwI6guBKFWV8Z4y75nLwnF8NUcPqtdaPrYv
kq1/+La/cfy9lJB3q7tUB0w3DAIPgqEV5AnG1J2VsyfUfVgZeVHgozAjWa9MhKpD
iu9cWkR8niUtKoBNyA9dnfBzr8csL/wCjTEe0EKvCqBkio6m3SowXE/DFjWVvw2X
8KrWwd6txbnOTgD/ZPOsawx/vX4/Q++5PBPhHB/UWrtkEJF28l9GjNbxI4zKcRvY
Y6Jpsp+0cUsTI6xaC2EbIU4/zooVAhmRY4R3vq4S2YjjT1SGOwQA47l7Fqr63eUF
R1Lbggcpdf2p/nUG/65R1I9jNfDlfvSYQb4yEiyKl5IWolYPR7/Ds2HLZw7QkcRN
n0yxxjT3YUt8sQeKoDOFzfhOEbLcYWnO7sl3li02TKtZ8ZuUED7I8NaRrT3vDYly
Nf7DnqR/xUTClEz7pTl1268npFPu1E4kgAo8p2izfuipUPPNXwWc98slWq5ibcrp
c2dFFNZ0Wfgbsa0sDuFf22ktIwaxdLem/MhxYEpVjbEKAKbjja+20NB5SvNc44Ad
NW4+V11GJOQmrjCirjBmPiRp4rc5huUCsuXr+Hy3xjSYZV4phY0WSFx5P7dMzhMV
6nOSE9s6ZrBmdLGWymoiSLWNC/sl+wP4nzTPnWKzNP34iK+adR9nLQZU4IlPj0NX
rLNmFsIHE4dMpFP2j1L5Q9/dy74nTEsEactc/6qnwid0yu5C/AGMY5T+0I0UDDwY
awtlpii+4JwGgO6VaZVD45e6Hal+Pza/lEUJVyFc6PEOjJ+L2XG8VUzXYfVTuv03
x3G8x5/q6W+t9Zxz7fkHklC8mPFBEIlIiasEBIusx7Sk8i925Fe7RiWcqmR2dRPw
C4bIo8KyYrUr2PLzY8ffBjbmBktwX2B6q3rdRkTWL7uRaqcrVbFGAeu1Hz77ebuv
jFZ/n0PLzkXq0Kh/tFBum1JUrzJxY9cHedMAMN03Wo+vmGjFQlEl5r46bgvDjT3H
4J3JT6oT17vs0CJFFKLSHAXeu5vdFi/psRZyXQccNlMZAxmgEQdcnVbI/lRmhM88
nRJ2GlOhwpAGAIlGpjNzKV9OZEA2x3O+6e8K/CRfMSjf/ICoY0Tp5/MGeB5dpKOj
1d6ojgl+cB6LbINZUcxJHssiMEq4THaAQmf0weYXI7xTRH0haMv72v/FdKAq0Jry
6BE7BJiO2smxpHSq4I2aHyODSdTrt8Hd0KauNv/6LvXLp9Y+P9HW+gzXulUUiSzX
KXNTi6j09al8enW+CS/C0pMiMTIZGb78HuJLdrFdwD41D2mwqrL78lowJWbz8TVI
5BqRd9ClgIOBBoQAt7POfA4rI0M9YVISM3ldQNNJUWjGxQc5zgy8Gio3dE/40C0R
PbStJuzAuX1v3ZZ+6WslPYOsme/Ek+14yFFwqtesqmBjeSLVLt2v4/wQhFy0A1d+
A8unBKtEl/GgSFTCxAAC5AMT+D+kaVz/5UmMB9/8uutvB4y1gtc3cdDgeRyBNgwh
d2mrQ783ExyE/+bMB5nEGZ5/Ppj1duAsN9ru7zvQL46S60hnROhMsXxbxhTCMMXU
I3xZ4hfA45OKsaAJ/XKjKHJ/owg4+RgtxX0SJyD3kgegNM55sPyGOFk4PRLrYoZp
KmzBjjmFvugAdfjEkNsKdoXCku2lpav6/G4c6kETK5P7dvol32ULuZP3M95IVaTz
Tc7leq+hb1S6sOouUZJBIWZrv28iqSP8SvFDoo7H1nqfZnyShyQE55UxtX9ReHRf
Nc39GD6vBbnSYMjQHwiPKnyNnR5MOi/Uivdcv5swuTUEShYrBzAIQ4DWoOeVTGIb
P4cWTaATcJzW2FcvVIT03n9AQNncTtZE3MiFPU4n3ZWVQ5j03gQ6assbZWtfwy2K
jB9AFYwXfv9TwZqPmsa8nI9iZnxySYa6AaHlPa/eHYYC/7PLxNVPVrfUWUmLj9ns
tvPWa/K+3tPbXbJFjIPWeF9W5Ku5ozVaFlOBGcstGJC0k4jZJjbX67uofJW37dKI
OPPdVwX7aBt3IibEqtxba2X/KSzpHEwBMTgm/9dkxvkJ3JPIEbtGhnIp+djJ0yqM
LgN4093qa8eaItqHN1Qp6i6X2wzRr5RBjzmmuWZnTbuX6cTusSlY6/fs95RXSNh5
qaT97LhVeMPB5lthjI8yqSdKeIHvsDlsToDtOq1P+GrlAlBc/CxZnQK7y+PBwX/M
V+yJQuEM6mPKgzqcxsvSqwQuu2kg5zDSrnGoOQda6ApgVRrShqjUckKGZehpe2sA
8Pz2dv3x4SNW509TJFwhji9tuXWqu5NM/I6S3b5Wffw+bggMVSNO8pZJsV4UCniX
1hLSViVmIvyBKAINpvFFe4aWKVIzdKka7ZJuiGZPTzaSEYuHUIxqK5nZHj8EMpv/
eNa+6hX/o7FcbGkyvhLu3o2d+Mi10rf7kCt+L5+hFMng+r1hV4G+0AfIHLQZxKb7
7EVFo9CHZug4x0NM01SzFB5yIVbdPxYWOx8YyNJwmHgMKLVdgiGGK/9CuE+LOqXM
VEcMWJy/S0JIJwJYw2d332W0UiWWW+2ivgQm0AV88px1bx8fLO5jbHwMCN6tGCCg
cDfyRMjNsx8ffEH9iTLzWeFn8n9sqDEyaFTUz9OHxvnx4qilLnDkDF6FOU67ThXr
1TmBcYkzfJk5AEym2CdTkAurL9SV5LYPHziHfr4KBRXKTznkcKNohGqi+hQ5tFib
nsVw+DFubA6HJwGXAR9Pp2y2V3K3aoqz33MP+P8l5fV5apHuQhV/9q//69Yt3/lx
5VVCYbwheIs0y8jxv4P/YhARgP75vnRNQ/lFW2L84LiDSZgYZLGHP0yw1dS79i7F
L+/n+5D/lr6B7Ms52lP2QJxIblcxOcxkeYSs4+hiYAAZgblmKs59xMHM6nbYesD6
/GgXrZtEBNkyuZLZv4jCmGdvG053P0psq7aOKwWAPrnYtFiSlpQPUKMpL44TSQzQ
KOmaRCg2MZGCjx8Ugnz+FaD1EbWXYlbhBnzJqB14wPjfD7C6VwemdWH0vKr/3yZd
tmFs9yTlaPIq91L6De20p4vgiGiwpSVYDomaVCs/Z8Jy1Z3PYD0N7ylBMxpBtCWx
GvWF5dAQUjoqaju9OV9lmhURroCG9r/GODyy86W2/sFQvYyDhyhtg3n6zgf7C9MM
tI5j4no3WITeW68VFRjVHUd/f0Th2Dn2ZoofyOfvo9wLlZ4O2JoyXXd0Py/z048P
8XT37KdO76Rqsb+iYlJPbAX7Tqcjx+qRpDObJBodcGQcLxLiIAFXWhDDpEMcoHOq
UyBRmoLcFpGiF90a26+l2TgyL7ZExh3HfJY85JEv9+ioolok6a4sKBjPNgm5CUKr
KuEIE+of0GEwbJ7HFvrL7Tzkl7WeR2ley4q6OvnB78bYo3FdPiJ2EZQr8yxAaQKY
9phVif9gjKVFX0v3zfif3TTuBeFk1JbE8o4M6sJuaoWHn60nlJzPV7capGLus4fG
WloVTig2ju5qMzBCYT1l8IGuyvHaOBukhDEXIYC0h+NIX3ZLFHW5/aMa0JUeWDxh
8pSCrfZUOCSkeWV/0FtP4vES30BnoorUzA0fWB0HkrSA+TIUi4kJ10F2t+lFrJIn
BCD3clSsCX3vEXBIqotDtIs/yRmyeJbx8EgaBn0pbQGeS2Fn9DxxhPs47wSU4oYf
hH/BvJaY41JTMdWGPUTHrklWIBvk99Rac/518FFnXlzlPYqNixLouNTkhByem1Xc
2NJRAMSC3Q//50kgVftJd8Ypy+I04DnG2kUQ3HVgYd6anwnWOBIjnnk76S4Jj1SS
l/POiMENVvKztifhpbbJVZa5V6UezOY4cGArfAFzz+s/PQzV0EkHHFsgvwcFcrP+
rMZzv6ZzZW+khoF4mEb2hWmjtfoHBqZ/J+2ifaJCVhzpUHKbjZyIPRPMCt6xHMt5
VWDpPUImj8GuHmOAiyO8yIHsJb2xdOSgauzREfDSm7EGBDugXnRtT3o2Vbm3UgQA
3SjGV6MjZGgh6SX2f7g02jdc/FugUHfWVcSZ6JuqLw5ahuNYmB5eQ37cdZl6OnU6
ZWbuQwOwxhtSOZobtQw5swE3tVCk+ZCUaYVdOIEBROlKEDcG5qetli57FQQKt9wF
RaQ/lMsyhhkWJPkA1bFELr0DZ3qnbt1sq2lZDdWDwDqc5N57T0Aa47wuBckvSSNL
AU2XRP2+9lG/8AUUrhJenIfbIRj3RHES/ZKA2zPuIdBbLm8blNUaqsC2DJqd7fpR
wO2zEGQlEWOWigTS0n4Qwh6A6qMGBsW7nYgFL8BBLxiRe/oO2Fik5JFCzrFWbXJO
44uqMwrHR/Axs4P57yTiNC6n6BNGgIyTT9oyUvXVkzH5V5hUfgrGsDWno8pObEx3
Gk8r6WIIfQ9zspwqKo5EwhTc0GiIrKkz6X2dTjTyahgJmZrj4Eoi7lcA716FWO3j
Vq0a8V6fiRWZ8BFlBrIUC+y+2Os994ui6YuUlpJdoFViFBbhptLyqg20qWYQdBin
704Kf3MH0T2dc6EReh1uTuPV4PNapxhoQMdAhYd5PYYeFPdL/1cIQqWH4UvmPts+
+Nno8ijvjqRdgNRFi1NbnBvHlQtQoftjj9urJyWgQEJNDzLZu5HgpkUFkOcbl8wn
bPFIBK8Px7d36HLWKXXFrF/sfC6OyThyDxyoZ909j8uxpNY9GkvDAsFwGn8xCSgn
z3gzyVrQrYAddNXhJw7NVIsrMi5jQJ6MjMr9SPiXrXoOvaKuQWwwXUC95vz8M/cM
9WrLn/oQC1x4/6Vc3UdDIxp0lfqvKxPDNCeR4MfYQ6UShuv6AgVa0hO6fFEn/wZW
Fm9gjt2fhAVfpG9JffPvOfoDYPasRMMqfmoYDVWyQGNTHfaJU3OZmO9hCp+wmjPT
TJRLiutaKuMWUeKqmyFDzjIQxwwV9oN1WKQwuWIykZ8+q5ZOyCih/wS44Rp2AGjl
73UrwEbN3PltoL9WVx9g9w9/GV0x+3FrmX8w1di8IrKzI4ilicPEATn4ChrvNwz9
3CJTjwWWzlJ+1+cw3nverEVaIV/JGsHx346qi6aNBkOfPlr/dqnx4CP7mlZX2AkK
OsmI+CVYSA7Q2jgj0A2NLWl/Cxue2ox599eyzOgkCBOAhQfpB5I0a6vj+7K5tkGP
Yie+LNQZEkzGMjf2+c5J2lYG32YB1IoITNODjCNFBIEkFP4WWS02KxFUglsT6+XX
RQFUpDqQjFmzCvxZKI7NjY6/OJkfBmbEda07+DfwinGe2gKe2miPbXTZL3vOMxG2
uHwpY2rxsnklyGggWjhGOkUtICRGV6w06M7f0NdIEUnH/X7JzqWaT7ChSDKVS7pd
QNuv/kI1N79WI3Ih9QhoD32uP3TjaG/dx/Q8WrIsigwduD+rwSNDwf3XzuMkWIrN
XndZc88FbrY2mnphx4F3TSA/2cM3ftvxzODVltomb6uU/hD2vmyGMmiYgELT0zuh
MHCQ5LG2rUtAZQc+1rZtB8AqjjXRj/3L10V/jnxvUpBjkXmwgCzdYlXrDCBrzKfJ
jvEQLV/M0voOTtK61xfQxkwL5p6Lkb8T0DpBo592sniLMeBBeyHYX4J1AHVXE8l6
ylSwwh26TSULfyOnOH25bEkYaPTphPlydU7bTSNdvEMyE3xDx4cTGqoTG58d8JXi
TiOSmDIUY0tJ7OdybxXUZS2Kz8TcAz9sg0EBHERYN56CJEoJpiG1ZuM2R0ao19MO
j4/J2GTEl2TorEWWEF5UBQvQPt3cxtxBS1AT0eTZuM/ST7YapVK1IBHHmP068roH
xT6qPcfITXmry90++Nurx/VN9OMXDMMmiAV9V9Rqz5D0zlN59R52XSqJhQUpZzpb
5OSSeJL0DOiBBg+WaOjFiJCu8h6tmiJoWAHNusS38R39g3hbrez4IPeuHqj+4u0V
fs/foIeVs1bkDd751rc5nZJ2nidps8xz+kCJbvk7eVCPMnMVXZqH4iNEjXKGoRrc
/v5A50zO6BoX50MgbMNLAF9lozpht/f43ML9DPkegqb3WpyO3Vr7ewfwxrhl30ko
6gBoTFUQNp5vECGXVN9y6Oppa0GlmoU5fLNnATgSKSvmQp0fCuLxY9SoqMWVvZM0
7kUhgn1HQVL/p7j+B/eYxUCRRM7JT68A2+e6XEMNBY5GUQCcMOD9kqM/AnxEZSCm
uaKIGTRWrUNH7MqHEP7aUZE5DmzjBM/g8R/heoKWaOia4Bj48mK4BXJs8fvBJ1vc
adfxrCPFj2L+v6VlJ+VKPC2N4pUGjWKpMee61FkYBK/mEq5gsNuqh5yEJRCcXEg2
fIsMgJTCQG15IYkIyyFpa8Ak+sErgHiUnW1o0R6y5y77Q2vJYTaRJjb7JxcrDgE5
i0DEsQuOxJ2vJNnduRmd1ND9qHkKbeL04kPJ6phqdybFULl4eXeVgNF8VmUtZ4Z6
SwPCR4nAbUusVbMg5UhU8vGpTtMCGc+do3O6pP00WpY=
`pragma protect end_protected
