��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�=���,1�jӛXT�d݂���"�(��=k�N��'�
�NX�yW-)l�Yc���ښC�eI��bc���0Y��rl������4�Z<Ί�Yd�?��?�:��1p�g�e�u
�`G�ʩ����}Q�-�-=��=G�E0��F�lE����djn懮D�3V��)�XQ�	�7�}go:��K�]��N�B|8��N�"7�ԮR�7�ۡ����s��TE]�Dϡ�G釳��i\[��)��%d��,˦9]H_���3�֭N�����?����*�=�I"�~욇��YE+S5�Z�
�?ţ�p�Rn��n,�eր���T/���\�L��m�g��_���cr��Z�"�x�J���W�3Ѳ�������$�d[&�x9`r�]�f����y�<4w]�β���Njz�!�H���w���`��?�}��'31��˫�%��m3�˟YB��d�ǰA�k��m|����'54X���!�%�)��p@�W��5S"Bs8z#4tQ�v7���l���,B�l ��Cm���e�Y�n��t�Q�^��ն�B�,0%]��H&����UG�I����zq\̞��c�5��g�G���k�p �*:��/fhLD����TjϞz<4���oV�ZaG�M8O��4kZ�x�󴁲�'pyĿ�Aͱ������޷��*�&�X%K<���Y[`D���A�!ssyV["�EE�ϻ'mDTg>X���!(������#)r���k�����m�}-�ۧh#�`Q7{ /5"����;m�)i�L��V� f�:�%#�Pﲒ�d�Wfu�e�M��l���/���U�&��8�L��M��躗$+;�<<�+e�~�WKz]��K���ʒO,�A"m#�����	������U�U���(�l��ʸ������c�����w@g�r�'�ѵ��>h��&��� ��	!�!�*�G�J��2d�XaI�IBD������c&�����@��p�<3!I5��-wg�HƓf�4y�l'�8�K*.��z�:�D��kۮ�8E�����R��A���)X�qS~�
��7$51�����%{�r`3���vX��NE5��R���E��嗫dZ��9�RhR�Q��>��T݈)���֕�"���7v������,;�J�*;N�䇔;]�5�t/�%1��d��8Sq�r'�sθHt$o8�o������B�G�.�F�%~
��\��}'G({���R56���<��=�՜0z�f�4Y�"`��Իվ�s�ߺ��X�}�;"q�(0�&�x�6
���if^�.7�+�NI�=��{|��E�~s�s���AS�bkmzL�=�b�(����	=�����`u]-�+�{��S"R%E�cq�v���\6?�m@C�z%��=�;`ǽ��wu+�U�6��2���!�.|cU�[\"y&�\�WoZv���:7v��Nٰ���l}5כ��N�H�
d�	�F3N.����kZS.��r~�l.�b�G�]u��ꗷN+�<F��nOTU|_m����̏��Lj��K��g<Z���ؾ8�-�R^�Қ��i��W{��N�[��
.�z�O���Y��CR��������ߎ�d=`�y��qj��mDziw�_�2òyJXGO�X������HDE�"j4:�t'm�� ��v��4i�쌬�ϐc����=б�go�|Ǭ��
����ѣ�a�9��0�����\�B�+�Q�fJex�/��A��@�bXz&�OJ#�����u_7D�R�=dbЍ��}*HslXEE���5��q\�!i>�^����?W��x���k4W�<�<]#/W|����~ED�/��e���{9{�>fU����;k?�h9���:�y�~\>����X�~���J��>�ƿIM�&'��V��=�)��r��Ш����cy�B���f.J��U6��A�W:c����1���	٭
��^�n~":?�7<o$:����Q~*�����e5�Ht%	�0��]��5L��i��u�������n�
!]�|F��;0��-Ҭƾ�0�=��q��6i$+�`0��)J�jQ�B�z�@��i�%�Ex񴸴�j�`J"ܛ����9U �l'U�6�L6��6]��|�����PB���[��6@K|c@�ҙ(ćwa�9|���� �fS��Dbp��6��-���.P'����IA�"��A�2,`�y��3M4�ez�>���'*"dD���L��%��m�qAԋ��XRW��b�h[�ی�!��@�&�Dd.�i� �/H�vi�'�̚��͘8���̋����#�m��ii���$k���#&������eߜV\��^�t��l����ЮN1�q��+�j}zX+�AB�޹Q�ۦ���
�2����͌����H�x�e�E�>�M~�iĚ.,��@�jm]��&Eٝʓ<I���+�倹�K���+�k{�;������= �V,�/Nt���p�+F�9�^*xЫb�v�TR���Dv�(�f�UK�v��y��+] f�s����˰�� ބŵf�����"g� ��wMQ���Ȳ�wX�������V��#Q�L60h4H�sl�Ư�v~��!�4꒖�c9V4=�E-��`�Sm+�G�������G�����E�w屽�P匋*�6�e�)����UO�٫]�[Rf�A����|�O�>L[b����d6c�B��c�	XQ�������旦���A)�$^�� �\7
�_d3���;]tgN0�MQލT�SBЛa��ͫ����V�� �aS���k*��XN�ނ��.���^5��§D�����8b��m�*Ҽ�)�]��E�͠��3Wd��PS��_�'��[����=&,xp'�֣n�{��C�xŖ$Q�S��fj���)����tKt]ݿ݇��e{�bذ���Tk���M�\C�Jb�\�`!Yy:��$��l^sJ�U�EMX�G�ۃ�`�\�;���m�r�X��<Q'�ЋBKOU�I��$&�f�_q��P�� _��k[pE@*$h7�c߭B�{vq�!�K��ѱ\����a>�T�،jT\�]�Fp�Nv�*٧`���с��SA�L�5�0:��5�y-\e=	@H�JZ�Z(m3n� �.K�=J9��$���B�Sd��x�McV7S$4��qp�#[���VC	���e��n��[�8��9L:����wi �ͯ��S`���fW������0�iAD2��tC�����Z�~Lv�����ȇ�p��P�5��.��2����ǋtk�X`��a�^.� P����+�T��.�nW��	�o)�����f�fdb\�ݩ��u&�4fW�`�è�<$�C�PTЕB�4]^3ô�~�*�;,3�y�k���e�.䝸���BU�`x0��;2��3�S�aJVO��߾��MX�z���N'gܜRo�,�[͌b���gq�6IK�4��޽��T�=kb_=�7
�>��Z�Zѡ�]L	d㠲n�e�s���T>����nJ*�&c��.;y0��)p/�OmZ��3�� 1����2�W��A �p����,i�����(�+�[���_�߱�8�Y��Le(�6��I��.���Sf_��q���O���uٝ�b�ˍ����+�L�:� C���
��>���]���h�+mZQ�NH? ��e�x/�鳧c�}8����l��6ay=���zL���5dr�̓��n��̒�k��s�0ltXQu����BG�#��%Q�s3��<e���H,���Q�!�;����	H6W�'&5G��^������pe~�*�w��^d��y�r���i0ol�/z��m��N�e�p��*z��!ش�?��dbu�����jTv ��������}5���>l�`~Y����K�.��Lu���G%{`���6��}�&���0 RKz���|��Y�Qc���vr���g�c�g�i�=���^ �AY;!�A�=P�XGJT��	��ZCieۅ�O��H|�Qxx��Lɰƒ��T�ڃs/Eq$���M�=���*_OZhP�|E� ֻf�Z�J�-:84�WE3=��[���h���OA;|��^���G�d��4˷1*�>�f�Q�˕%����t�j�'�ێ�Lw �;<f,s����\��2(�cn�F�	�0�ǮƇ�G�?/ȲD��l��(�V�6� �����$2�����kU���~״���N6�آ��K}��U�'&݇Y��?̳H��-��>��ݛ��Q��SI��y���~X�ta~�E��s��!
{\���[�� ��ˮd��>�' ���W�mKK޿U%���]������:�������yZ�S��0*9�H���U��}Q����Ub�t�!�a��B�v��s߯́hf�~PF�ޫ�_����E�F�w�3��l0a#��kw����}���(���u��NܧE5�)킜�%�]���3���K{���'[�~ړړ�x���nk�D�ԝo��|ԤV�s�H��u:T�#֗�<��CS��@J���!Z�����I/E���r�ۘۘ���L����2�-���&�+X���N8��X��c�q�1�A�Q�����ˢPT�DnxN�k,Qa��J]��墵��Zx����WIŜ�)p��uEae�r[߽�.>��u��Ѝ�9�,>z����E��ڶm��9�0�N�i-�Fo�a ��%�,�۹�%�Y�뾾�������JsHfD���+�ĪuR0�R$�$�C�ȸ�M�?��2G 抆���UdQ�kZ�� 8��]t(������>Wj�K��]�b�Տ�D�4q�)��h�۫�¤F��ڼr2�6����pz�wINV�j���a�Q��v�6�i�f#��BTgy=�a��!膝{"! xZk����>&m�� ����.��vR�[�3x"����vq�X�Ul�Y��skA81�ٕ,!2?;�맼4w�)Ց�x��ҕ#�[!����P�3^e�0.?�z�]�y�t�[����>��t�ٟ�aafA��61�M���A	k�����)#��C�Ol�-�y㉹� H2�*c�78��2ѓ��:��p�eF���'V3ECT���m�}� ��i}�[�{@|���edA�rp(ל>�'���y�@aI���}��9G�h��e�j�r/����H?|*� ˎuc?��=�W���E;�Kb2�i��{��ZOR��Ǿ2|�����
5
��G��3�I-�L��$A