��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9h��=�4�n��͇��B��0��8�� ��xMzd[|��^]����鎉2�Y�O����c�m��7B����*��Ex}����벶͜��e7h�!.iI����H�W��$����t<D��^pA���\�^KGM��?!��󽷲.$�%�p�1=�.�3�Kwu�Tk@��%M���G��,(�����!>�lݝ�Z��D�m��6����9�zxA�fOM"?�j�W~��Y{S��|�_ˀ<w��\�X� .��N�U�@��c�A+�2�WM�+߃��k�8>�N�V����@`���E�9���xQ�Be(�5�}�6�#ECZE�?rO-̧@]S�W�1�G:������Lf�v��mqb_{�=l�Y�N}3�\�t��y�6�a��d`�.�x����:Ӡ.��̈��p�N�E��]��Q;��;�Li��"�JLhܼ\x�v��p��Oa4ؖ���`k�+/�/�a\���w�+!u�0� ����?2G���: ��y��)�ć��:Cd��PoE�w�5��5o��c��0��D�H(�ya�5T������2�<a��)�o��A
1�8�o&"]������k
L%y|�:�i�W�B�1���v���;�"����EH�P3����8^�xd�ѵ�����st�uL1�H_���<����M�(L]�w������T�Z�k���03����I�po7^�~��;>�qX2gؘ�92�D��?��Z��q#�q��fə�����E~�;�6
��cEhG u�,=��C~���#���G����А ���ܷu�?~z;�5�zsLnZ��ε5pmt"�Yb��N�v�a�A���������6��R������/"5�ҕ�k�D�Ű�C���U���ke^y�E��"`.��%�,�u� 蹷0$��ʕ�si���̽-gP��?�K^��F��Ǝ�n��܂����k�6Q|���������L0��%��ze�8ou�ц�r�gl���;e�i��qyykUe��x���'����#b���J�j8��5æ���T���/q����쎚���������]L���+�YBi!XC�=.��:/����bu��������q�z]G"?�#n��J{h�谣U�������J������� ��p�)����f���[ZP��5�5��f��z�y{��`�O���D�~�"`�;�F���������ȿF�8�]Y�AOP�bJ�GF�5Qj��x�`�[dv@D��d����}�g�4V�i}ęp�&N$@W셪�t��P�	�&���L:)G��@U�W##yԝf6��&�l�W׵ѱa�[Hp^��I��\١a���M�BE�Z`7�O@��"Ӡ���e��a>e���K��R �Y���ѷt���.@�i��Z�o�ݭ@�t��ɗ?W�k~uB���>#O$w���0�W�&�r�+�� C����&��h(�q�>��Z>�?����>G�"E"�{Y�QV���9:���$�[�٨1ϗ�I�̱�0k�r�9��l���R���{��R�@'����w�V"d{)VO�Ǭ�硃�%4:���p�9F>KI���7ad�=��d��L�c���/�Y�OB�\E�9�*�����ɨ�˨�6=Oa�����E�x�ɩ�&�/aC�z�;o��Xw1��H8�+M�45�A�����;ܹ��hT�7��+����y���K���u���%�3�J�#+f�(�� �����^t���9weԻ����&*��ɮV�b��/������&r�<�H��WDO�B�!'�zh`� #{<��-p��?�[8�\~��Se@��:�<�g���7_gʙ��z=8؍�+����<q�Ǆ��tE��.�8�ހ�fM;b5���%@�50!a\Z�W�y�Qx��sR�&���$]��9��R�HIY���ɂ{튕�����|Y k����ʞ���%��gj0�&	���0���8�F��4ZH2�O����C�<�S�1����� �y���o W����+���� �@�ae���z8��3�ڶ��a�oz�0�X���|��d��r��}��y���s�^��\��r)����S�>�����B�X�i;5D4ʿ�\���,/��nY(�;)��G�B��S޶�~N�4=�b�󸏔�\�9�i2f.���>�C��SO�W���##�/�ܩC�..��73��o"��~t| ]Rn����,���D�F���)��L���gh�~Z�h�3�g7z�~A�����`�Y�e��1���)@���v���!�~���0x��/FyBd��a������Jө�v� �U��u=�z4��cOu}�$����%�qz_gY.x�������)?j)�/S�Ԧb�ܐY�Be�<���z<'�Rb�����?\�QU���ˠ��@��c�L�b-���'�:��.Zh�>�6yu��ν`��G����[c=���wʓ=��^7GET7
�K8��a��]�������;4�zT.�~L���N$m�N�*�&R��74�e����X���7|��|3M0B�-PX%�Ǿ���Ӱ �IR�)�T����o5}�P�@l�ʢɡ_ݶ����Ec8R���즀�����Ҡ�����4��s�W�U�@A)>NJw�똣4�f:����N�]���*�ɂ������m_b��m~�zme�_e;\i��HF�n阺�.0Jۣ�(E�>�asΊ��:��Ͱ��?"�SϙD�����[��n�ga6�/��(ὅ�]��pe
���`3k�nt8�QfN���P�-^o�<-S��rF�5�N����L?��?��Ku�l�_x�KGO����53�%*�?�����?�0�tZq��Q@���:hUrXi[{g޸xO�V�۝�ao�x`tN��}�M�}:.�g��&o��S>a�fQy! ���w�yyL]lf����k�D�R2�2�ζmW�.l��ee���O�
K�=�}lf�O��8&��E��gӄ�|�d-���������Rz�+ҽj��Z���E��͙��HQѫd<�y�uq��Ђ�znH�L[/ �h�������˟�x��flF6vҮED�랔C>������hO�xt�'X��80cD	�LnS�*Et���#��1̶��x|�	��k;=�O�������s�s룔� +!h�/�#K&/��P�Q���X�b�ó"������2�zȯWӿLK�0e䞫>ܟ�s��[ȕãu30݈7Q�)*�(}6%@J���%	h�v:�Р�+LX�-]9B���84��yE��S[BF�l��^l]�n�`�%W�d���?���7U���D��(H�ɕ��ˡ��nrF�D̃C�#�8�M�>�Iȸ��T?Ȁ`u�?tљL���Q4a"Lg"���s�̰__;-�8�6ܲ�*d��?(L���KOOm��~F��"OAZ�p\�B^�B�ɐzU��.��!屏o�V̻ZQ�A]k����QLm��~u��R2{�5��KсS����De����_oMOJ� &kc�Ë��ni0�qZ�s�����n��Y��$�$�}�P�0�~=Z�('�!Q�V7`��'v.`��+~6��o�x�qQ��Θ��}x�_��u����\�)���� `@�ғNP�ک"~�j�TJ<��XHgݘ(1/��h���E8;!�#0'�ta��,r����@zY���
�7KU\���Ʀ�r60`���F��.
�߉ov�ץ?�e1�����;��Z:�CP�.�kݐh�69s�h���%0q��R#�U}��-����݁���F��g��A��P�N�Ek̷�Ũz���M���õ��B �S��eBG8~O���.-¢�ˊ�q"f Q�6Wo���� ��by���:�
8Έ�O2;L�y���bǻ��T�
Ks�VSd�%�#�-�.�̔��	\�Q�����a!�cs��ʄc�QC�p�P�w��3�=r�e���<��O��`���@�V!��PۤR9(�'�d�U�=���(}`���\e�'�Gt������{X�$BX�	RX�UH��Q9D�:fοF~Pz�$���~�5�_���������+E�8�&��!֔�,����×�<�*���tC�Q�H��R�]RӪ#��Þ#�,�� ��6*����1�Q����`�9f��L��oȭC%q��(�X\�,-�Q��@�P5;�{�����m4O�f�=aۑb�#��o�b{�<�#YEp�L[ٔ<�׆D5�#�t��-+���V��n�D�&�����N����s+�i��v=�z��BM����x���W�}k��r���*h�5�?���^Й&���2�ף��E�Y��&��J�S9���2�HfvI��O*��$9�j_�7�}����A:�W:]|f&�m8��=LR�ĭ����d�>P%G�A�"_�?�_�t��!&X�۩�����n�Ĉ67`��5����4�uH�q�ޥs�m���^E�߉W�<�T������5�!��w�K���sJt��|�Q�_|t��_���E�o �җ����#2��C���t���?��9�H�+7S��p��Oz�-�PIHY=�8]�k�2��V�(�	gJύm_5z��\�n,���7�\�7���y��{Y쏙�����u-���r��P7�5�ik�B���6ǽr�.���97e[w�aފ���~�⁥`��A�w�Z����V��	l��C�d��O�]�j��h�:��68���9H=�UA��g����uf���d@<�6��mM�t�������>��bg�7]�]�JkA�c$�?d@���Ɲ��~ܗ/F����zX�+x�8 S+>4EI�l�Bם\�l���ǱA��gȏô��G��o���u|/kMUZo_�t	7zC�p/�� ��U�J��I��˘^C�ݕ#w��0��x�lKC��i��?4Ũ�H@�^���B���p�~���|��5��+U~רp�̖��jL�kc4������7a�VK ��  !�f��d�d�(���nJg�[�M9�*T}ģ��ƒn����È����L2Wb��t-���"����Ѳ�2�_H�