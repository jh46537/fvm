��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{�YA�<�~Cv<�%�������>����p��i���t������IV� d��~�P.#�U�d����u�eP�1��Ɨ�o?*���K���?�x��;}�n=4pÒ�<�E��炧����w`��DCp�*=�G�Z��~��JeCu{������a�6^��`9Z1�U�Ϻ�L�c�Y����5Kݞ%�DS'��a�(�e�!깽�L	�p(���8[�UB��c��ʅF�b�M�5&���GJ�ۭ��e6Af�����͗{�w7����m��'��)�l��2h�o��>Fk^��Z�rA�����"Qsz#��⴦�'�^�s�̎�� w�e��-�Y�"r'@5��#B�ӵy�ܠ�w�n��e�GdC��r���!9����ԮVH�7�Uʠ��3y�Y�xY0"��I~5�Sf�7	�����3��^�y�T���'�4h���^�T�Q%Hȶ��ˍ�fKI��TF�	O�X`��h��0n��o�IY	�':l&��� �����a/ՠ�0B��1���N��q�h����{��h��?40&�C�Aw�^�w�$pr^%��,Ch!w��2�y�r�CV�Q}c���H� *[�ʳ*�N1�{�ŵx'0�h��pۄJ��������f(����.�5D�K��or�x�"&�h�Ŋh��1�,�
�����%�~A}�4!�{?�32ޡ��|<J����	�p�z�TP�Wի�K [EV�#ق�=3�#@�Q?<� ��nˮ�qBQ��ſq��mp��<U�}�%���,]M��0��w�\*���o��,��	�{ V�]�#3��Xo��\��.w�zւ�i=M�wj#\*U H�C�+4�����L��ĹHY�u���:TQ�t1�'T���(v�P�F� �#9"d�&�.q]�����O��ߖ�U����G�O��d׎�!	�8��ŤP�~���y?��Oa�����J��X��/yr����2�F�R��T"����Ԭ:-1���� IvV	� 3p���&~�]�?CO���F/���O%~(�i�0&s�$�j>~�M�;?Ԝ��)hM��+��a�����0�M����#w�I��(�E.���
�N�r%��擬(E�{�j�8�!e�ʣL�4	��֠�J��y�p
��L��M��μņ�c���$���#�O�*my��6Hش0 ���Ym!����-G=�Y�L�֓�a��?���ֆJ�=U�^cp^���i%�Ɋ�5'���h}sa���|�	 ~O��3]U%/ۢ�%Az �Q))�X��a�"L����޵]]�H�&v��y�{�7��q��5�S�E��q"�X�\�C��pվ�L+e³Fc���+`P
j%Ӟ�����,r<;kG�g��w��{6���Wҩ&9��:>�A�1W�NQ��p�v!	x���x���h���ny#-C�Ip����+�$E�y��0{m�r��4���O��?�y�o�*wRH�|��<8�5��xg����n2،��~3`CKpC����1�ɗ�_���h����S��ު���� ���k�Х���j���l�Si�6V�#�˻�����'�a�1 �h*w3�xU
����6��YE��=5 s�eO~:���7Px&�i��~����ܲ�/7$��#¼�,�yZ�G�UYN��30nBm�*Z��%SW]��h_k�gѴ8��w=�G l�A���$��j��G�Qm�}�}d'3ц�݈GsF��Z�]Q�E}����,��N����Ap@6OGK}ի8}��X-��ļ��#yq/����4��w�H�.(�W���=6����pur�ܗ�����A�(s���y>{+Vk�1 ���C�,R�8ѓ�	:oU;1�0�%�����Ͻ27�U���!��;'��Թ�f�`�X"S�`�����I���^~x���m��X��<�.܄���ͤ�U*R�.D�8�'���M[�q���!!9�Ȃ+��i���i���>�];��s(ɨ60į��l�w����t�_����y�!�̕uV�H:�Z*�7��6�"� �@�ZD5���5x��	�������޻!X��ϔtK���tG&+̙Cц��N�%�	H^�.��(x2k?��ur~	j��]�N<M0��
+�Daj����|0�x%߅�V� ���؅�����dT߇��E�;�+n(����=W.'��ϯ�+C`2ܱ*'��m��ඏ)~�APwf�JQIz$�~�P�AY�ٻ� �������@k?B�n��������TC'���&[��B��q��fmloE��C>Ʌ�_�a��,�[q�V]���C4�} �6Z $O(i��4O�t����hǾ>2c�������aC��b�+9U'W����ޔ�������|�RmA�v�6⢹:ܺ=�ƹ�Y*4�-�2:�T�h)�)��,h�������B�D	}�.��p����rX$�����֓�e�T����CE�Tv��9%l?��h6Z�e�.(�
Cs_����D�ٳ�H�%�l���O,�G�:���b��E:�H�
̉&�3�\�h���n��r�t���C��<��	�RȘ��9��j�ٔ���
�3_�'JȒ�������TCFǤK��(G���ϰ��#}����ݫh�ǡ���7�K���Y�Iѓ��%��3����(w��Vf\1E��5�9�D��x0�FS�ᗏ�?�'��+Z�%pa�ʂ�'�>���� V�����H!d_̄�;�h6δ���~��/ޮβ/���-ݍ���o%-̐��"Ӛ��,��6�7����S!H9z\��f���<jg��>g��J���U�d�3�:o(u[vQ��[���u��]�_�������1�Hg��:�.J��	�x��Sj%��D�9ӥ�w��6�C��@�������q�2r��]���i��KRO��wq��]����#9��a!�V~\ �%��a�yn��Bz�'�&V���Y�T���z= W*�[-[���x/-���a:Vof�	�����ݟ�};��1�#?T�# }�j#e��hf�ƯGԷ��Ř��q=!�ܪKIB+�q����9��mVCTIh��!_Q�J�����	]�hm�&���c}=���9`I�4��Ӄ� T���e�l�ז�ɭh�S������$��U����c' 
��36��b%;B1VI,� �R�7k�2��^���)��f�wLo�v-Qfqb�}Aɸ
9�VD"Yi�a��WWg���(Ǫa/U�r���pf+����X|�^Ur�{�;����Um�e&�����e%�pa�p�������_ O+�F�~G6U�/x'�1h�"����O��KV�K�?>7��]q'$@[���f���UMYҋ�g��=>�����w�t~�l�*���ǲ����kX�\�?�B��H�Pq��<