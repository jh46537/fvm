��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�;O;�n�Q�_I���Qo]�~5.���X�̍��ǔ�&[0>ۡ���n����r�V� [qNʭ��[�_��r� <��V(�݄�J�K�b��0�
�"�x��zJ�nzz��6V�e~�۵��=գ��g<r{^���$Մ/GV�"�����γ *.�+s�()\E�|ۂ�d����OůYMehe`g��h܇���A�]�!,g׌���@������*�P�>���\B�-Q�PR�^�KE���k��w#�A�۬���ʳi��t<2�o�H2��9~C�_�꒎-���J��<�W]�}�ڍc�-� S��u�ٴ�?H�w�h�Y��-�u;'9s�5OX�Ih��-��~�s�9��]Z8B�3Q�Oʝ嶟�~��_�pV�qs�h�WHa��j'`�S�d���W�I ��5l���Lk
��{ZC�1�k��c~J�9�=E�L����S�MU�⾱A].��?Fv6Pi��;�lf��	��6�B�!�0�y�6B6�/�oQ'9öX8\U�ɠ,�+�~{�-&�:�C��~$��D�j_Τ1K
u���Z�ɪ	��<<��T����L�^��D��Κ���ȯÆ}�6(ה���Q�&��(e���]���}������F�6Qn�ͫá���GkK�YC	�yA�b��N�@��6�`[.7��x7l�hB��)S���e5�r b/��P���M�mN6k+(�&%���_����1��Ĝ	/
�qޛ���QcGSO 1/�Y�.�:e��]�p��U� a�x+���`��K�� P�pZ�'��0H��uc��jl�2C�I��1hw�ǹ^�L|�~�{����
��V��@��@(�D*����-�W���{(�o�/�J~�6�'=i���m��n1�ǲ����W�(H�$a�N��7S)�d��/y���@��W���YSs+�ďJ�7מ�ݷӌI-rN�{�q�9PǾ3��a,�ȇt�yoZ�'R��ǱZf|��g$�3	HA��6�Ƙ��v��o2�榲��jQ|�Gd{��j��8̾���*�^s�S��B���iZ�,mN�c�M�¬dsڌ�V<R�E�6��B摘(�
5%��Ŝs!fq��(#]�Wɴ�T��97C���6A����I�R�f}'^L,Q��)v�7� ���g#�FL��y�����t@�buIǫ��--ayd���
�/}'�>p�aN�7[��
��ArM���Z��d���YR���,�/�rEmq��k��2jXBM�Ӿ�	�H�W(_�.(�u�on���L4>���e�ۅO���G�� �>���,��{;`Y��'(�� o~�%y���45t�×_��1��ɓJ����
g3�X��@31��3k�q�H��$��N	V< pz~�A3ԙ��޲O��	��z���*OښW���[�`;�Fy��}p�vK��K2���U7":S���P���o��m�%U�`օ�����B��Bo�kz9���( �����=�:�$��Q���;��3F���"��cZ	����@Tm:k���o�i��I���}�[��9q�<��e�=0���G�Ľ����D^N<^���yQ��><��L?����uI������Z\M:*�\)]*i�f^Ҷ�~�Ծ��0��3<u�v��T%m(B�Z	��/}^���0�$'��;il#�`�V�2�ά��9]t @�6�{��OX�,��Oen����(Y@��x��;?��j���T��?&�7 ���8��C�/"c×��߃�9�U�CKj�]o�^7���m'��g�mG}��:j�Ji�ʹlh�)�E�=UU�����6-,�b���(51����N�{�ӵ=�8��_}�m��iO� �k �c�E���(��dZ����G5��7�P�@���@l�ip��5�/!h��K�H��F��&u{�����V���X\���X����)Bڃ��/�~'.]�b���M�0,�D�9�@����}.G92���G'�Y�����2� 4"��ipl�pڂz��_���*�ڻ� ���w^i��366�d���]��.��w>�E�D��љ!�~�Lug�)f�2=�/_�0^�C"�~p�D��T�MY@vtP&yA��Lu"���f������t�ŧ.]c�gRT]'�f�1��_�����Lob�����55��������E�UhL@|��z5
g���pe��}��t�Źa�"p�L��Iuҏΰ*��Ku�J�P�H]�[E����g��]��"��԰�Ḓ�\�wew)��4?�O�e�־��B�}}@���=�Q ��Ť�/'t!���zM4�{.�e�@(�O���n;�������Ǟ�8%��+��ȗ1�1�'���#��T�Q-�.�6��TRe�b�9-ܑ�Y�o(w�*��k��XG�&#I�h(�A}^�X�&ʬ�7�OSB��o�(�ɢ,���4K�>J,��ز����e��Z���.hN.��A�A61yf�'	��lkɼ�'�Rb���l��a���ȯS�4$�v����i��W*�MX�k��de���:�*���mI��H��T��8�䷱ڦ���%e��B��K�(�`���fviH*���6��]�R"�;�;A�u	��!�]�U��X�ȣ���zxQ�:l�t��2@�O��C�\o%/4QL�T_��K�u�����q��ZL�6<�\x�zUw�c=[�;���ZM����d\XJ^�#�u�ڪ� �{�'{��<��Ade�+ �iciSl�l�
P& C��p�s��	�x���;���Y'v��*h�I���~���͓����ڷ媞̤�:�(z>X�M�>wDy䯱7�/�FO2Q���s�M�=���8�`C�^(�����,U�8f�=��	�m���X,J������r~���� �J�N������p4�uJ�C�v�SF� �}8<��lS�.Q$�;�+�fE��fN�.�x�A����dh��`� ��bg ����a���H�E"t6??i>�����N�b�b����H��+��jt\�a'���ޔTx|��Ω��w}i���t�7�Z2OG]8FL�OQ��e�(�#���Ɨ�D�S9f?͐�h)��Q�W��zB$�)�H�Ž/N�!��x�!��6��6ۤҝ��[6.(�[�]��Q����C�@5w���`Rg���OCS�#{�k��Pa�7��@��.��_�?E���;5���h�F��7��$���TLdr���w��t5���^�YH�%BZE*�b�m#�`��xG6G��s0���,���%��
u�\n �2^6��ڰ�Q9�H�RK���A�Y�G�{�`z��$*ĳ����_N���C ���kT�rMʯ ���Sz�ռ6�gz�����n���'��:>a~�_er[�p��f�+2SZ[���o��A~"#pAi��^û��_��e�\�g�q�d^o�L��ι��^#�UC2����c��C:�
-�(�vE2���W�~9(���A$W��E|}�V:3��^�_ ����P���3p�����\߉��#gdO������CY�: 1x"��a���x���e��/�|[/w�p$�Cäu�����\N3����s~neZ8
U��7�+I)�g�6�g����؁)���i��$n���f_O¹��:�-��2t�e������3HE�Q|�U��~P�ڮֺ��H���2���d���0�,n�ݜ�\�,��Y3k�^m�i^1͸���-���5�x���k�Y�/
n���3%�����Q��kK��v�Sk���G�#}Q�D�E? 
��8�1lR^�!��kJ+`/n���O�h�B��HVSFqz��� �&�����W!����n�t�a�lr4�}M����D%��{��c�^�N�m"b��\5�fT��C�"��S}H�p��m���Rޘ��t�[鍃6R�p��J���Ά0J0{�
��<��$��|k_,H�s�+�J��d_qA�e5��^J���"0���x�%�BV5��X�Z{�͗�J���y	\k�E��8MP��I����T�ǽ훴zi$��h�ןD�X"F6U���L���*��d.#R�:a���ct��Sܯ׽ksU�,���T;@��u��\� y�)`i**��zK{:J�Is!�B���\F�B�I�7�y J�w ����p�U�G��D;<�jt���:2�3��k퍸y�h"����(H�o��Dv�g-�M<e�C���H�mZ��j������I�i	�zh� �����xX�K��8�̸@O��JRƵtɃۗ�dh���rr�0Gin��Α�w���"��J0ͣ�������E&d_=r������;-����W�Pz�wV��d��R4S�#f�W#��9�u� /:�5�����&�B[��bL���0�;�2苯�s�ry�