// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:18 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A7IgNbCNGYl+y19H5XLpcpUVWBpkI+B0jZH+/nyTmygHr4HJAYm8DVvC4VcgRwSo
rrClLFLwlt83+aY8cm/jzGSTazAHZPiy3BkpZ3IfyANiCZjFVP9/PQCt/F0pEKzS
6Dsn+IbnLrcXcvNhhwNlSGIGMqms5/8+ixglh47BPNg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19760)
oJdnsGbpynqPX0JlA0kUx8+BirNDzlWcbw2uUsRQJGiHyjx5bqDy57s6RAquCH9P
n5/qiI2O+n3OKAoMWSXkv/54C0YgT5ENiJ3jUOdAWgNP/ruRUWHHTgPWnJlPcXtK
7gh3vxAqztLz5GGQoS2mv2jkdzbzXWyVhs+1cB//korp2ZnNH38CoAvkOLm6/GBK
iUiAzHgJ3xV6HgVE6ix/i3+7fFHUEyfN1vnafbNB6rAoBSzAyTlZKXEdcT2XeMxU
GvAtyo9xTnIf1V/8V4aR6afG9BmpIT2X7MYo3fxfRtBxPvkLUFv0xKtqac7PCRJd
zde1Qk4o8+Bfwt6E4735UJTY/vdZr7tBMTFcFetOBT00C5FQEcDLDf20ubCNEbkH
iCxSWJoBBpDC3Dv6MI+QPJf/ME+YQuTPLONGh1FDRUZfdIt6LNw4CEaOfy9hadwv
21LeMCPiuMIg8IKIdosqHPuJffTzoEVTFN6R2MgL0Z8vbVbXUltLUI48wnIZbo9b
j2YqfkO4SZgThwOeJYCpgc+9QWla3p3+9g4pXPmEcdMf/Yy/ozUMoN2SgCiyeWaN
DJI6aEAXD8K92OlQIHnqfjI1VkNNw8wzC5HPr6RaiFdqOnRxKDL2afiV1Ee50XBS
71VJY/1H7OF33l5X5VoxTFnG6DYX5Ydw2Pfn5NVt/TbnRROXZQLlQ+PJqnP4Ld8V
yR5vtc1yHCjT3E7UL9q4uzFEQeFxcFiyXcnrj3KCmy+v9w+fT6VKEW0+s2Mosl0x
4XTspLMNX70vqUS8JAxuFHcTiZNlvJ26P7UzArbLOOMRGw7hs7V4s8eP+Ba17iRX
XDT6NTS3nIyTj3ghhjpRmH4Rulx/3SU3DIwkaklwXD3i9kMyEbIfKXUVWIdHG5JS
Vj3RYTyce84Opp5mqs2D87GlvlmOdEPQiyk88CNOIK+yZyqc6BClNrlAtHWA5LXS
gI8EtSxjnQmHbYQ1N8Md2fLXcs8ChwrRWXWu0luNqUihBUKh8Nys8MMtFJZw9WDx
+Nzbn3yXEiCtwKpkOnh++zMRv0MGvjNjlJZbb9oHm1TrnWChzobG0V0oJJBWS9z2
9Yc3OZCq/jy5OD4+1nFzQYH8xzm/P944+xNB19JybMOlt8yWvrCFroqKgcvMOmCf
b5F9p289rzC0bVanhAlPG4eRJmwKuyrRAK1uBvpcZ2sqOAoyxo1J0KKe45rbAC1i
gNKJAKgUCw2eH9S3L6V/JyGmuRxlPOJG+bKHzNv1f/UXfVCg1JR6FSEc0/mSuJkI
66leGqtGgrCjd4zr165bgvMfKBOsAbYtdQMGHMi7xfBqUOactdSjyPQkFrgBNodH
jtGwb2uOLD+gCNAdXyLu0FpQ/crtNc1n+7KHGVCdUBu8C3Cqb3VpAUAe6G9EinYG
52dcZYZeIIHS+bs5cChE/fhFnMVFGyOARbS8p09KRLtPgRPl4ksRc2HUqOAvFiFm
c2sdXVT1fdsBb5JpNeQWxY+sws63MhwaGDXCcpSeuyXlcAFXp+qYuamsVeMKHa0k
NRQPsadHOjWeOoFWwQ1PwJCRP7m+kbw5rH4R8/e0BrC4K/AyUuXi9P4RcXbkWr2h
EuwLzQQD30zkdD6CvsUMYo7cwVVhfpN7t07pn4Y+qXpSwf4QgjWQjhdwYYvGYpvo
vlMnkN0ri+T1hbC3qaw3CaM6t9LzpFhYqKMkg8iWxHAGQ/48WNKeYsBmgz4tdTFt
L/fWHONm6uzIHhOyvHcXG8sOyiK1F6L4uUSk6BjIdLytnvS8l8GeyRq8JfxiXrG5
JxJ3dPSiOd3y9ATrk3zNRJhU5o5qwvLAQ5/QWPswjRHMZj2j17BGad6zshBeLWeS
onhD7y3WCwS5vG4N8pKzHb/58bym9WnjB95vwRb9iHFSIme7OB6zwp4x0eO5IYDj
K+c2Gp3sJfNLsd8Iw8ikfgP2XLWTTS+AQ5UbDtHO7BPJKUUbZuKXpqe3jz0B9jzW
P+wb0Z/s6PdyNE84h2VI33CeuaVbr0ZV841AE5LOCvSmWu+YRbz3SQ3cZqdIfx8S
5+JEuF1yZGp3SvKm3mr3TZMnZizXN6TPBILztKZuESN0iekwHlxUn25dtqzQ/c3x
JWjaXsLCnzUgSEA/vG9VgwyCuhdCBIw5GPiP5AJU182n9udCetyvcBpp00d/LaFR
//IMdYlyeg7MaISeRx/QH+09nRoWQQxyCBvoekTbRLo2DIF646x2GZBidl4XN+k3
ysjZ4YJi4IK929Ae/Rn4QnnjqPcAtItIzUeAFgUiKD5rvsfnlowqJT+YTErnMSyL
gfyktBArBz4wi0k8BhZfU2JTcrIyc5QJ1P3Vriy3VS/OVqO8/pupZ5jAIluswpXH
GXZqfo7utkuYQZOsyfpjXf/ep9JX/G1hOPfcKvqWeYl+3HE1MOQi8h4AVN0SlMKF
iFM03bV8zmR+M8fLaf0v1JUWJ0DBp/ELzz8Pfnj/k2FC3MEonKKAe9pT4Gi+woIb
SJvc6kyVs4XnQH0V+lzeTjnohJVVbULO5gUxdwdHVYxv+Mck4ooJ/j4V8awLD1EW
wDT7O+eVF22Li/lcWaKhUCISXU/ycFrv2eO4dDvGD7T4UImgCzI3fUKtZhi2CVXB
mtLVexP/o2r0YXzuBEtGbCLmuhEFMU9iwyepwELWsiJWBUnfdq6AovWpIWI0tTQy
qEe7XgsF3zh8yMKYgPXFgpefVdMDIDampDBU4xnSK9CzOnLp7d1F8OOiCPWb5sQb
JO080sszA1VbobQDCvCsX2TuD5JB+410dNGhLDu1PPLOJntzIJtj8ouZh+VPKRsP
YU9YD9pDFuGS71IOfu6WQdtHKcr3L/AwyxW1nkvLn2meWt9Yzk5LCgrDR9/i2PVL
n4MHmmyg94OyKoFxULRMh3l8Llz7ZAH/vLiLQQTI1BYtFUlmEFOEMJHWfP5C5rIm
qF9JpQbCxOHCl1OCek6FF2NezXGhYYn/A1KPws+/cEf++al41xx1YHG5frfB9PxZ
dD0DRK+mcp0uzaDjVgW677xU/NtH/FrQTeASu72YBOTzqKy4jTwDONY51dwuWA0K
yPLin15LMahTiUnWt44UUUMHfRbsWVdc3ogAQhQXH/1eSIa/Bpdb9BXA7aNkKn6K
lMXi3yrei/y/zT8wjuQ93NOTqoujwEf4QaPUoitScPynKYRLodJJOCdgGIJv/CwF
XahkIioP4sfSpoDI3XhwW2h7/phVOz8kTwH+0WHx4+SB8Aw0Qy199bvva92jGnii
LWv5vzqOUF1i38E4za62jK4sz+eGV7juRvLHhHf7x6+39m7LrrbfyJhxN8kSN5iW
Hdlx+gZSL1OmAVmwk7iJ7RDRk/a30sDDziaMa5LADCb4wQVmEhvEQz28Go2YFGkm
BGi5b8vLTeSLR31/ZN6Zyhapnk9emuw1vCVTPvw5LzM1mwlwJe9poFHHSqI16GUK
Kr+7kSfyFB9Ot3qKOAxIigRs057ByUa7B7hQOGkUKR0UMq2bR5PHozLHNoeWDCPV
/3i1VqJN09FCFBfxYsmsagGe1canIrcmi73Bk3xS+T7QHHoZO0ro+Tu+uEysFxqo
x9o19P4LJbUN1nu1ZBbo8TKtez/XcuY2d/fJ+FOm7kBIm8O5yathjhiUyKkzgCk+
3nOJ0TVdr2tZrwselMhM8F9HwWFkLju59DQNDeccACafdCEOduUV3n6FfE4t+7Nk
Y0P9rBtWUICDI/a+pYKLOlun2vUjG6O4fECHX0rFJWMC8y1TvlbY+rcuhydnyEY4
yVDc6jMa2V6uPtrzzqQLuDQByuH1Hsb9vo8wlv+XCM4ntr0/9liKklefKubU0A9m
BI+d/LLHZkkt/u2qs+NvKkguckl3Co9kolB6ynbCSvQpV2RIzp2pLWNC7TSLWL1M
GxuGlmPMoOUDLH2UL4m3dG++BTtpRcS6SFpvJy3psB9yGYlmQ+XPtonJIDMjYcHj
0gTM21fy3Z+lX8OjvwDzB1iTC0IRV0EIoCNxJ8HkP4NP8Ky2agQLbHr84SYwIbno
p8AlWu74MyeV+6rDZrEjyDmouNVQ6gE6abyBenQ/YneARWSA2VflsRJ/U17w+CIR
JDnckPLDVJhlihTK1tvWP5xIZBTF42SjQ3QuMsMEw3z3vK7biqJ5eVqRhdMFYf70
/wiwUDhwzKVQ9Ei13PIzqN54tD0BxxNoQR93p2Cq2awlF8/8nME5zzYjWP/KBLWA
01l7iYlJbTCXqXVLaCJRmzuGmJVAqFJfNqRLvDYuWNkZpGwIx4grinZFiUwvHXGC
VSnquFh8IlE2P7PZ3VoawSiANEHFaitct1WvySjfzKK/rE4yVM2892SFpILwX3vO
kX4WEiTXidRd9LektXwrZXAIPe6A1/EpF7tkKqf/JgMm/AdceFx5Xtfupoqk+/tX
XioNbxNVQlaERW3AO+2u3HP+pcBWoCIBlmDzBm0Wy13Qx6qbsWSaicJ1Ug7KSd7L
YR/AqcF5Gu8hM1t9lordKzAh1rO5mPZ5KDl37LiqkXQBTU+ficU3f8Ee0cY/7ZBb
Ex7BlBzSywcW+hwNFKpNq1A0RJ/u38Zd1j2yhcw1atL+5TyrQ1OeH3Es2RKdYVbn
nf5aQ3zlw4xK7pNeYhBTqJ63HD0kOLVaXfC40I2ZYRpAugI6d8JBPyyd1UIPcUGY
OlQUme/EPlQp+fzo+5JIuNfkXVMYETuyDMvoanijJP3brbELxsBhFViq0fMV65m6
2c4YsZ1YvBLTybBbO+gYhotmzTEeuJ4YBdb1kGt/gYQA1FRGRc3svTl1iYKx+kgR
/ijR/m2cIwo68aTHHkZnzQDOg0jbfJ9yYAAiY9Rys28MtZCpixhO00aaaVe4VKLg
+htfDxZMvVV9iXIc4wXvKX9lv93+Ooyx/cXN6EIUqxerVd105RKhcqOyckTOsn7D
yqC5HjrHApKGmKij6Y5HKLp7chrTRSUsKFrQYTKMidtqY3w6NT2yOK2sVHP99lcE
SqEEpeLZNrZtVgmNOiSsueb+F8nghU1H+tO9BkuHQKHH7OJGP/xKrGgRoEVomw9u
upsICcjWpNadLgYc80o9RIefNVBdeKwK14UethOSTxSd6Cc3cUzpMDlYXlStJj1m
0Sv6oYMGL+CL7JLT/7/IglvHPnqn8mguDtOLDo9mzqfGyfLsKgmhyabpZ5oxV6pZ
JIX+2+6tc47AXu67BNC401HrgemrGyMAeaaqSTfBbJE7m3UqNV48gMDkUzFeqVdv
e7uWf42OiliiuX9EAutzOsAYBZjIEldnINcFaA3+0qJSzcTAEx0JqUNf3aYJIhK+
Yxc8jr8asNSI8HOqpRJzuBzdSKOwg9MeAOtpQrwryC3STgAeVf3DK26d/P/Ct9iJ
mfju8UT55cnRiWY3JXC/eZYm82+Nd/Q/JZjJwWzVBTutfjmbgbrTKOHzqyG2d7DY
hREETA6VfbOTcJC2dUky9DTYqPfOOz42sC4wE8XaFfVAjWQop/JLSbgr3VOLS8gS
7WXezVzu8KvYuY69ipAMLIyIKdKtnr/2IdsjvgFyjCRlL0ZJoZOrIrgwPMEyfG8+
jmDjZXocLj2oDx99SGIahRR48HfmBPjJKEexqLONeNJ1fIbMImd8dzpEYbjnm1HN
7pNl2f8AK5is68NHwykKs9rfPpAiyiRHybFu1eEmauC3KlBNS3Ot4IgIbF9ifKTy
bJhDE+f67n+05FYo1XANHiembMPK0k3cbGqiwTw0tnPevTRYpr79zqz+6kPs1P6K
SMnTPTpylsPczV45SOyNTcOiGFEMRCjx1EbzhwP8hhmHiAqJxjxXVQ/4mqP47shC
I7NfP7V/8DrKgywDIrQDd9GxxL1/6G035MrSfiSxOaaZQieH9gKslQxT8aGi4I0J
OqjNIErb78L7JKE39i4QB6efh9lL7evwrL8B8CfMztYKk7KH61zKBJrZw3T24sZz
TYaYT8M4KkQAdrWIWmrbvLIOKi+3uyz8zKMTU9ptWBRi4fu46vIAevge1Eveonuy
3FgzKA27OEaqR5mGjHAIY6n9BnCFXenTFGkwqqvGW10N03/r9pMg7If8T46shsDm
zh87HxkhrRqKm4Ag1RBDuBfcbNuvAN9WlLMxwq/WlEIfSK79bjpkTv0cDE2ITQ+F
Rl0Ok7jPtEHNbjZJNuEmyCfwuF8i9Rvfb6Qv357ciLSSvx1yxuuEyFHNkhPgwLK+
kAezteMgS5wsVB17gecDeNQ0k4ALj7Ctf6mdsa7W8uElScjG5OcqImQn3+zrT5QN
vocllCr+1O2MbSXldHgzKWVq/9JeEBhi5yAZDSzVNGutqL9alJFdtIQh2kBq1CXj
78AUy+7EEHDF4Fu3Dhxe/d/p6yd/KvAy8RxqbITvqE8u+8Vzl/3gpNG1Gfxg/aYL
Z3TUw1y8y1pB0GbVee4t9fb+mfokP/sOnRl3gxls8fZI1CM+DfzodnoL0em1O7S1
n6VYFWKCTFVmf5ZF24Jjd1JWHt38JnKu0ssDNnSA7bxgWLJsi6FeZUmd7GnFKc5P
WScL8F7ZWmhvb7iSXFfyzb7LxoIFs5nut3fx8f48NEuUwNo7aNKxfLvYZ18XILBz
zsqC2jg3ZkVhvujTD1MONQZl9dMYJXvEgeRIrnh+ddXFsYR7jqdehOE1w/mxG/Dv
0uX2v8tpcESk2Jpkhv5zB3BDJnGA/Aag+8UvK3j0Z1z+eMHfyGSpYNPjsds/cnpF
0oe+Z0GuhH10010BEAe7YtqPqpFOrxzvMF/JKB4kSq/+Hbv/gzE+58FZycpd0DhN
/6+Jupre1LMWqFa7MxsNKEBWXuPL0khfEMcHn2qKGZlhc1AsI2XVGahFYlAYlBPU
GFscspxgyoCDlCi4SGtVd7NNAIKd7JfJ+G4C7BqCZTP66mZholb+YxgezvuQTOkv
0d5DriSTaYLb0s5QptNepTdaYzfRXFJ14QthPcy/MnyOLJ88WMkq6EcEOBjmzJAG
iS3xwc8D3vLMaKou+AmEjn7JJW2lAgfEiJXE3TTopfOzveq6IV5HYyNlO8yExDco
gXYzEC6EUl2fDHgwb+Iu0KLiNcrVBQuNfSHTQwdl+I+FjtwNYbx4OCKhnKpa4S/s
MDFkdhX4JswbDTpCppItqM2hHPg/b81J1aSohejpJy67Sq94q70gKnqa9ieRWTu1
i1kunFRdALvnkui+daMUZt/SQubHJ/Tars1BcXTyjMGMWjeQPjPSKsMWz721Mc3e
7P16FeUgX+RZVrUO6bwMZY/Vn3Vl7md9lr266FlFBnCgUascUcO6U9edmcmWgio5
iYJbr7C3pbQBMPo1SHyevbG7FEcjsIEsHJtxytYWQ7+aLqMyg+CSAgG2RVT/V/md
cLXu9DHel5YsqtZW5l7UYkIgRGZ/E88tmkt6sIz8l/w/rlxa3cQZEHDcktIneL8p
3jkXacBfToKUexocB5kVgwMtvq7imrWgeo7pNHAD555IFv6n5D+DtUQUpLZLoAQw
DT/o0udaDIhqJBcgbeyW5yMQZfArPkOD26vUM+J9CRmSosNvrb+E9cQ0MxEbTY4H
4EdXLidDIIE9jEeDO87AB+s8xVjnZvZ6pMMHzhOSAYygm24OhC6rLjv93LUon120
gbhZHSFaggus1Lotapc4pGFU4YbVpqEGblrWH5uSmwpZI02m5bavMJ13g6ys8MEF
xvy86RteOzrJcoeeY8pvwdPxSbxq+VHC8xLZXOEGMnOvzWFP842E7l2YckXevSCw
loUMtfDftfBEr3PEEzGNoDJSGRPc988JwM/k26EOUTT/wufjBPCjaawbO9lfzU8L
QXGn6/yzF3S1RUStATdqmLAn0mUKjiiSUCNc8e+22bvMqkPXyGzi0kl2JRBM0weO
7a7VvdLN0klnCBNgci6CDtWnyw6oR8YgHxTcJ8FNDhPvAQACpzA4925EZh3ptP+E
dCadN4hsG0dcTq3xKK4NDgwrcO94OzavM25/kTvVNFUdZ1cRuqp0BtLHSWMXk6vj
ncKpZYLyjvDGCduq8fbadSz0Qe78UUJ8FDkf8qxSzYhoZ3zebzghHN1lQmMyRO56
GKYuQJ/Emw+HIABZX+jKI9EUXXn5pOIRvBTrn9Fo8hiC6m+dGwCJpzmdddObdm5F
kNCJ2RK+DXHv+FJJ3DW1EOxCHkr3PwaX1XwftcDCSyUt7baU9GcIcTv2FBJEaNpd
EFx/KslScd3GpDVHk+6syCJUCRoVr0tmE2e0MZt/AUQR8Xm6az8XVpdiSPGlfeau
nhJTMJ2pSvqDpKKuScLVG0oaRTMXqTl8lwtWGElfCzpnJqJI4NbqMML7/ABehMt8
Pr9riYb8ohDobNi/UynI7OUZPHGimf4SmaY5DfQQw76wfdmy9jYtBOEBEh6bXao4
TLdHlGoyBkYDvIkzOgt40fPYXMEL0oJ1OyWejABUQxLuZ7iuYhBDzngSEJTZ7O+t
prYxrDe+TKkrJfLo3Hy+g3WcnGcpv6r+kspMjRJ+fBFpk2Z4igOleVB97/8fzQWw
CdDxGxRD6b+BVByeiCz4OnJJzQWZWzQcV4Q49u83yWvqiEZr8zEFLkJF4OcvBWhn
AO67RvCNl1tL0QeAA0a6Tr9jghqMPGBV/MKoyfVr+d/HDXdi8YhKCfN5GWGbdNfx
W27REGhouBuOQAN3rkI37MMacU3YYseZiQAaUy+Y6kCezHJ/OVJTyZQQEAPcMxwU
gDj9rDr+XTy/Hi2sWr85sG3sgRHMOaHWBcW1qxDshHd/mKTXmyVxSQ5BuLP3EjLp
+y2rt9oUQqqW+hpxxyAOicsTa+4uUxqV6T0jbmOr8Mj5ZNTRzconHwhTssxCJlzE
lzCVT0a7vdl/T5WPvkDDi5EbuJgYxfO45IcQMgc5JB+c/5LM3Q2qqe+vOr3ZlUX/
zbBsG/PYdrwo6RcKIuzV0Bi5Vk7UWDVnUHW84N9sf9hUjCMZ6G/rZAcpSH7mURiL
XxmconY176uxD2CmRI+QM4F4Dwz/9+7tdBz3j2xBd7GFybDuSouwa4TtbSCWs4Sm
K+j5lXpzxAUINfD46dlXWC9nroOTb2bY31rO8HBpHiEkc66VH9HOIeD+t7AeVByf
J149v9vlIyOOqOsDYg/Yekf1CiuFeRITHSQHsU0ETqdyfYzltPceKsp2MEq76Y/l
FZmwa9vuPUNdJ23Odn4lv7m6lU+4qgwqcgOnIhwxhpRsf1emKNkofokBOtmgVv2I
T0JzPT7uLUVtrjFN4USzKphshrh9BKqTylNl7raFzYK7KACSUGcoLFLkHfqH+ve6
RSzNHqw0JH3nuzOc3s6GpDqCJRPZx2ISlV+6ic2vsOhmeIRD1ou2DSfOmX7tlbk6
8sLSsUalnys93SYVHw6lTDQEXN44ijhN7JKOgQGjObBFSu+PHc7hHqsZMtpRQ6Sg
luVMYTyyWWD8ZSYMrXCwgkKVGo0FTKmOIC9CU/Fs64V7I6UsTzi3vHorKYC0AsSl
qZheJRCxt/PfK/1qDD7aFI0vY6ULFRLQbHBabLDFwzoQFtyvPPZhYpIgrtKPzve1
Oiv3+tVGdUsBkpMpbfynpsoXHyDuYiprAEJCtNQRwQu3v2EwN2s4xGZTkVb7o43k
VP1+W/Nx9kFDAqEDyYjhmL/LivDve2aiWNllsNddDCmRNtgtvMfBSlP5tKhvbtf8
dQv8SEJQFRJPvEsTQy3bEjgEWRO2qSnOgE1Pv6uvzgNVoAtSSgRv8GnFmy0sccN3
YuxnaijYd4LZQRLbTLJXYMAfACx0O2WIrwjF6S8SuPB9Uuh83Cbt2krM6D6126lE
0CVgXrCCYonHiDpwjT3CwVoY96NRENvqsKh4FZeefcPQMu3/eBLudQJbsW/Ar7G9
LO7CQRVB9ChEUwRwT48tmQLZTsWjJ97vSGGQzoRK1LH0v/x/sFqNRBH0zbtBA4C6
0sn8fotQVc+jqjsBOMEwECpT7jxLoztU0/DgTPQW4sSq+N0qJcoekDREze+WHIad
TEaWKQi6aBk4PyKqMuVOUusw9X5o6qWwwEydnw0AIExuZO5LIWWSjsVbzodMSuWE
1GB+YAJilvSc8GjcHkOkdmmOoNw8EL7yNFH4yBEK/KE4QgQmQ/6c2Tv/kPVq/FsR
oJET8AvyU3QpJFuVr7K1c2mHLtZOHMb13jr+EYNH7o2j7z7Ui1XufgC/8fPXMk5Z
3pWW5j6BzE/wHvnGJRZf8x53ihselSrfOHGDULTFCtsUK+ax4kGnnGwGjMDhgjz+
N+dMNZkmzuirxD4mHCUXTTno6a4UayJL/3yRvZuKIUgJWUjMJUjIo7CFLu1SY1wx
39t9Gdnh2wjrk6S8PK2p+tYUK+YB3Y/2R6zS0abc+9bb1RGEI8JLU8qzSvGza9+G
b87gFjOwYwxTb3qWfK0Tgj6gPdWZZd8Yu4maYk9azpiaM5eK9c7Gyxbwz9h16riR
ZzjGTulusJnk47f9Sru9sTZ5oEbFEHzTGYRlZxRvpHPwot2Bjafg27TSMLvf0mnK
ss6kJxOk3wifjq/PlHQ8cm33LB2wp/Mrh+EW4uOeDW8dRu5iC3uu2iF0us/64YaV
l03YpdJiWZGgbyvkjOD2beEdrtWKUFZYXg4xYtJ+CWZSgLggy0jBGLOUGkfuGtJK
ereluhUtqQFfLSRbLD96aEJjLWrk8jG7vwCIeSqg4uWEsR3+T/C50zdBwG2nvMuO
NbmjdU7VNRAinWknJ06cIDs5rZRc1NEpr3FeETxw8Xh21ST6vyE9Ubf5j1IjCtoX
S0VFYFjksaxMs2ItcDiny4Y5EOX98UvwVqr7XEQNFc+EZ3mCQwREkG1pUdUxrUmA
cqRiwPYCMMeZLoRlwXqOZUXAwjZ6TkWGxgPyNRDw69P6Jr0CvcDU+QsvJRoQ87fW
EgsSZU3MyWSAXdfszVbve+V6PZkwkc1OUIrRRRggusVV+DKd5yoWYg7vbCCB8Cuf
JGbrd38TmoYzrdi4Bvd3Zd9Ki0fb5gPpswyBE4lD5zkbvcaJNrtktu+l2kdTOcbp
LAwGxgSFbbaU1Va9/K+4kKClxJbx40uewxnV/lb3wNb26ru8gHx97UmSv3WGippI
Q7I/RBOXSJsCyOmVFekpqAJipHVb2x8BcmKqmgXAUgrqHaHmX4SWyDz0qBhsxQes
CVZE2zPfOCuPkVKbr9ZybfE3SeD1SRYJstPUJ+DZ3ROyxz8CDpkKQDgZHehKRVIE
o1RfFTvWeCEG2cNf13rxykNNVlCVln+SlcOdXus+992Tw/sEIwSSNebtS5Kv5Ixo
QbWCdaA43Sut9HU4Q8Q0etbL3PidAe1LQbXLOtTmGR4ieYt7VOzcRw4UykTBrUZF
MkqoUegJuPzO7aS0NXkJ0KjfBS6W9OP7BSfO4rRXRoZJAZvVWuB34729q8UfL9XE
DrNXkOKRk1PFf8cX26XTSicGtGCnZ67siFPk3MnET26aqL+oZSAf0bi9UoQtpTs1
qNYdefzkl+cx3BuFLfYY5LDEDMscWFMPeke1QmdYH1HVOy0m3XOuy+EmB8J/kuoJ
4Bh5UjtY4E8VELLzCQDQszeyS/3au/6no3aaFcqnNg/N48RZ5PHs8iQTjQ80agCQ
VxnVcIKV/KCm85XscqXE34pqhimLqdoRe55FwISr1CacXvN/WIpGOfhM18AceP2b
qEo68lrk5gTeQ9UOXv6Mv19DyaEnLceEBOBJoywIloBBfOouu0houaj3FaEEJHED
1IJ0A8+pCalb//CQXoMPkjbDeeUcqoZn/zu9yPQ8R/bKdDN8cqqJ2rBWIMj6/T9j
jUGvTJqXMFGoGcnf/E2NTU5+vYGW6xODbj7xNNnIfBk5H4l5lHz4VaxU6r8Ek5Ou
FMx+X6jW682eoGHtvt7dp2RFcLN9KnBV4+31odo0SdwzJ2F6c4kAdDbssgxr7B8U
1unm67uSL5rzxI3te7amKJVRNpIwIylEXs4MIVOcorfbP7xrFgpceZVNwLs2/0AC
spSkoa+oq80kYGSpYca2CnKil8buLcCtpLLBY5u9zgm/rPEOt0SyVI/y3KMlZwDx
MqPNq7MLXf9KvD96c0FcWqrPPEd66e4aghMP4CWo6kzwOuaeMRtSaMULQTLqCxin
oIto3GG6tpNKKZRwbrLca/KfnrUs2T9DDthkTb9Ny/dMGtVCU+Q2gt16J5duV/L0
cVCWJMz3W8Zq6T4zRcORf30uKVw7CLKWVp/oT5Z6O/oeOoBIDOaW8EK6akGiMJM2
XExDWr8NE7v/WT4GlAfAVniL8CbXCxCDDUwy8Racs/JwrH6jEfmiTo2+Rn/bMXXt
6tb507/zsRB2Uw4a0GkVmtUNMmvx7Fh1Dz3CyJnNHLqI2G/zf+gL25+zM0d5Cvjw
Q3cfmYliK5XJdttRyKYzPuFy/zV2LVRbBOhsCPbx2Mrgtf0skroF5Tc2aFjD2PYe
JJiimQTyIwCFofoGrAgtmYQWCn7ap9gAkVcR6kcD44Du2u3y4tAMYs+3XdltkGuP
dd8Fyp7KGx8jLVwSlk5nlyzh6aoG7BWh4LDoIi4bSSnCjzIrWfZODxT2d+u43CZt
L9JBLw+K9VoBB8b4j0Bn6ZJVoYWJ5hJjD2lgJemDArNk/MuDZdQLG7NzMg0e0lz4
WuciR1P07ogWRNrpQFv43Bcp743aT+abvwZzu0yU0J8IrOqziGZjfiWURwY/TFnE
D+5aifvUn1GA+uT6Qjvt6WAbDLMZx1u56+cfPIU0+zzpUoFYY9f4Ovrwc4ofMm+X
BB0VAhIZRJq1Xab/W6JpLyUSlSyYgyuDs5cGIFJaU3nzEWjQSFIusmbmHxMarblK
u70nijCgwRslb0p2cGpAaLwpfB92cRGG/6pMp8nb7KAnrnsyzxR6TyXYphAPTu9V
Cbno69PHNfHphwOTJsVuCiMXiuum3IdPUebGfEbSWFgPKF2uZrNFlwiRdue0JnpP
ufRDfQeNN/ebmfPHhKqOYI8xHu2Za8PYgKb7LvlOgOcQKXKPwS+xZ/t3TKVCHK6I
/bfUQEA7wZZRU2XHwZwE1L9bwkCYLQGQvX20o+FbI0RzAspZ0WmApRxtHE3R/7Ca
eG/A+Q4kQyIZQiVUp0lhgIaSvBEVY3cbDuFfzycHlhNlHFTIFQPFspmLx3yo/wzK
WLKCC2d4rEOBHBB7gKMDLUtQ0wj/JLqJmaZzqcLOZT6mQEWUWe3pyOrACvi82adG
l0BXXYxMM9TB3YkmaLxrowwvUvCbeyVlS716aynHNxGWugeTlgeUc8Y4kZC9eVC8
eifMun3ysRLzdmKte9q8/sWppUX1otXeId5wYLNdS4s1k2IslTgvB+8Ul3H/nJAl
X66ofglyyMWwEP69/TEh4i+viyAlhAn+M/c/9TW97UNTpGdXGDqoQj9zENeCB4XX
ymeI+Aeki8jn7G4MyeznZKDVQTTfWc4gxp/T+s+hAW19RiAkCBoTW9tBsAUynqp/
GCdgWsgW/bJLhVcu4UPIzXJK27pA99ZGrDMYf96VkZ2aILq/fSITACwmus4xZN2j
YYZGZDe1bMCnqmU5NTE7eRbhK0+X7e9dlEzlfF34f5Uo/SdtbqpfzxUpCal5LWIV
MYlEAV9s58lE2tvjA0xr5D11h9k/fd4rJoxW5F5HoHOJJhMJtr0PSiUX3t6iLQSm
0ENBtxZUaEDYSJ7vsvvxyKLEwvxsIMLsVj2DWWi0g2AfnL6VW7Jq1DRntxUVLUw5
hKwpNMvGTbZB+adiRXgr86eulX8RZGXImN+S7XBcftlo4redJBmjzdFYg2hFUz65
naQ9emLoq0YqGCOjvSTosA5X+czeItKrWPVK7tFVwmt4VHl3YcC17rP92/AaZYSa
K7iEMQWr7BNV5TkS/IZOkNUFDu1ZxqGibBFEyb6VjgeeSbWV2eQnCelPQ91mxqTs
Qm96Jq/thAFhBS8egB5f63CiY6X5C8ZiabthrSyMhNJWxyPf6ia+MoKlSdDEkYd0
6lH/q34i8xkq37jYYhgH555iH/vhewbjfV+zosSe8ZPQHVW5r/OWJaEr6+lLqAIv
umC6CZPQdZkNs09I61n2FtAVjaqZGZzxzXo7lfC4c5G4Xf44yFH7pCClfZ4dtypV
oYHD/qUy0NQG2VT+Zj2/r2mrkS81qOHoLs5cyQ5cvXgegnawfweS6Im8QkeomFF2
Wgx6MwnV/F3UCAgYzADI6GUXLS/4KiJh+21GkjqqgsISfTNexTNYGMLYpcDhiVx/
flNUNW2rrNk2AWnok8fB1UCTjo9lRHVeM6lnFx6U6VhD0y51lEXZ1xI6ZWQb4kjv
8bMM1sIGqTjHYq6tp0zyoFqVm5M61r5jzS/0Ki4NA76oaYvk9goItz+NV9eV119P
mYTrgMN4LTo9WYuxdj1RnMZ3viFFVUWpYvK/JemWWtLTF0tMLh7UHTLa7WDT9aBy
lQbTn+trTc2CT16MTzcZxl3sWSld5KJzp+vCFnO7sN2aLQ3yy9sq/CPemKaNzqCK
egvgQgwL8/TQOyrPbuaKBNTo/5DDb09VfgdmfXZbA6o0jx8wEnZcRKghktT4cUb1
SW1Uk7O1w2siZqx4en1Rlx/77YyDGwhjSW4//nG1nfk5/tg4olk79Z/6BSF1WqxC
bYbVGk25qlRUqowfUbUyjSXzF9JMWV05oVS/t+rd5EfRB1QkHp30OGrA6quE+W/D
K4mOrQFps2yXeXPsU0gDxbM5QH71o9QcJ0L8ldxqYpHXOHzraM4JTjygvYI0Mm+H
d1VBaoXXTKJJBj2rk9aAgl8gMbWBv/2eRul4iB6vTctPFUt+T0zxCXFzv3hcjnuI
OhzWZHrvD+vHI+dtkUHw63X6dU1hpDrnDP8gAkWVLuHKUGk5dYsqkvFYBeMNnaeS
LWOg8adhNeeQFVrLHPHW+8kPwG5oLD14HbModMwkyTAwqoK+/q1hJFeYRzPV0Wge
SrrTD/dTquaFydaGFBb4Otlhl+m8xAE3KMv0bzkXFsdbAoiTMnMBBatPH26RyWI9
wAtqkblJvOSpQlg994rnA7VhmwJOM6q+KVDeMz3yfvZyPl4tV2fTX8runh16G3DV
UwRg99j2dTFV/NnsLQw9ZsQxxCbzwm8dopMDuk1VoHPjjPnH5N3cfP2hRAygZjlr
euc/dgQmcoicgD9kOnUv1T4mCTcOa/7FdeQhjzSBXOKWuc2MW6v+RZ2tug2UZaYw
cMxP0O/1GxcHdS9/qlFrUiql9/avfUpRwDgy+Ot3O0+1OcuB8XLwdDmlxgcZIJll
0bOoaUzRxNIpjull7nI/SB2C7mwBFh+R4SA/F73SguHMlJz0PcebrEI9Kv1sb/vB
Fj5rNfGmBdyZgJFth7eikzeaqRYuqhFPlzksYF6XtKk6jbTZ5YKiHIqpRwojlxn4
ZigfSzSqKH2bla+V5kzhQmR6DibkePx17y4UtZGG6fLudOZzN6atw3JV08YBpHrD
G66e4pbc9k0GFvW1w3Kxk7M8L+Wfbec0LoRMwwd/pM2jX0UOzqybfyAYzoidjRyP
aVSmz3sPivO7Xp0UL1ehhT8W6BOUCxfqFsiO80NhwLPzWSwCXsFzhhMNk7pUmnma
rJ496EnPm0APzpxSMjgyTwa0Bc2eCv+j3OCGjnG7WdvkQ6/W1HE6T84HxPJ2W+RE
dzirrbMaxs/UsY4ray5iLPgfolVEBAATPKuGeoZfjZ1/yENhKx4kPirpg3URuF+t
4I4sjJ0jKSh7c4xlMXFwsZQxFqy7LguT/S2ccCWs2TUXfMRr7qmse4O8AdT9qKk3
sbSUp3vZLYaLCQugUZaCDT4lynJgtX4S9H33O6kHXfJgq46BQjq1PY1XFk2VHpxX
C85APd2RtdNrHzXdtAf1YXAFr6KFretRJWb3n0A1zb/Z8tgBWgjKqFeobPCHgDDd
BI8Euh0p3MnWzya0rU6zwFUO1N9vm2jrrZ4a1YFyjettpwnigkCSvontvquXlA2G
2SQ+NPEO8WxvR8wVcA9zh/KjRo/frsixdF8Abt5qzk7yw/zTsyQp0Tq2VZUvEx7F
jQseNIE2xTRVUvn4KFEHc/u38D+WND0XzvM9RATAuV+uJsmIq8ozeUf/ZEL41RJL
vb1uVjRMYkBnXqh8q3SwpbHX4ZyLhZ3JQCgbBi1bVysp46M+MienjUq8LslAEpTq
aHIA0Bd2vrg5OulMUQQ6e92rzKLvwFv9rsxXqB6aYd+TbDw/URR+TGRmvgZ0Yvek
0gjo0u9gqcUGHggdVnJtrOvBQXmx1vhs1tFuaULMX1x9g+EYf4Pd8MJzg+hICEVP
z7E674x+aCNdrz2bpAQOaUG/tzm0XbJ0S4Q/57NzSu2rul9sbWIqRgEFnR5KguVB
e3/w1AljLKhSCC/y0D/Px1xdbqQah5ID1SG0DL4wgDJXtLSOvixRpqy2BquwZk/p
sv6AIB6DD8CCL5l+Gg20W5j6MGh7wTHLYV3n28S536K1Q+rfEve9cyNQjw8oxyee
GbLTN0gg/uMZCQO2/E5zfm6KDGkLPA4IqNgvA0BMV6oVtRRzAH7Skzaq/v6RmAXn
PYpHFjuVQ8q8EyR72oGGT5FoyfRHr33qfMg6mC+gaAeSnTFu5bFJts76Hn2tHlRm
1cjYDYLnYVwQPMugyPDeoelXgIh4q2cZAOrZjlO51yX/A+u0cZmfjUnJ1XiNlMYr
wAW77ZoAPfQKSZKM6cj48z5XSgIiBW63vzQJMmSH4Cb0ZSq1HlkyeD+/0gCwo+BL
Nw9+wYWWpJYAYY9c8jBG5ARnighqoEgujj3XH7nwzNM6e9ZV833xnHJVWMrIHymT
zDe0P5Wjq+PJiOIOz2+vm7vihst5Wjv4/5ry1l5IrLVrTnaKbGGxY5RCaAfVTvsc
j3q7sJm2NNMyCVBQFMUAur2AcvCxAAvLyx0e8QlYw3aSj4izwxRIcSW1LFeO/t6K
di0Ze/HYg7it2x0732+YOm92mETmaCH0fxBDwUUsnh3GqpRYaLCJFmNs9qnhCf7x
MhCR9Kt6eOMXZmXQoywMmEjTAd2r3HsXGqC3wf9r//epkTJA8xakyw/8tat5rU/o
a96/apo5HVM2jyROJljCSttxccId++BhHwvXtuW/inNOi9QsyYRh0JfPKh2hi5uZ
mumPkV3rBWI6ERgrqeEbDL8JkFFCtRCgtuj6PtwFhYKS9LC2bvAvWHB6gjUHTkBR
WROn9oUoAXYrFQCVRwcxZec+VxxMWMAn4KCBqBWtg2pIK94YyqDPgYY/vbzuZNpF
QSD2q0ImUhx5rr/4ByTEUvoAcz93GuYwhsQxLSKCaEvaT4jGursUUSW6yY3XkeaW
mshRER+cZ4ElmkcrdVz2ab7xnzLu3CVv8QLlY3Kqk/JPrwqGK7HMR7xWJNNWmo1W
+drmaSJASpY+klL3uSviagyRmVSKXSgeLBXWRpWYNwQGcKEv5nx/mwxR7kYTsSUs
30JOaqmB6k6/1+rSdVZLjAQAFj9NHQ2TOWVX16mTshuod8VxPwDcskyS/6wtIVUl
N5oSUIJwlLs+mKR4tWUQsDsqapqcxKJbr8R3Jmz+givMJYC7PNCNfp7K4D4De1OA
LfMNYX+uTzZM11NxtZ36iFAr6wtvV5s8HSlZhZLGloZNwp7URp1TTSOcMq0uf5CT
AcLnXJfgYYzkYbS/UfZYyl7vQmM7tFmarkuJcFyiqbkXqYZAwqOZ1Eoo3BxrDQ1L
kqYNrhZ5/HmKnYPisHS7yxDlVr5GEsHNDzGqY0BU9oi5OwsvFLDbQ6/nt1MCKu8J
VZCGCwUA5VjeXtVxZR8IkhtHxYwr+e+E8MAI2ohZdj8Qk0K5GLHyy/daPlMt4/FP
XhehCVpt12+GbRyunEytTTbXdTnliSvLMARqZ9JMkK6ZnRRBC9hPGrmGgGvAcnTb
dlnhMxcZDMVPwkk6xfk/WsyVno8oSI59DUy4IhR+6j9dJkdsdA+y1GsOo47jQH1d
zrcvAhjmQ+CNHk+wYYmcTekTwxPYMdtkje35tbVKLc/XeUBgQR3jA/6eGAQhk/m9
0VlnEH8M8QB0iDBV9eEdD8NVmFLSH6zyJqC7Bh600rS9gy65Q2vG/58iloWHdqmb
yWErUmgLsuD6bqeh9/i/UZlrswSEI2qLiau/7+XvAuiV8MTnym2W1WCLP2QXyzew
DKv3CpABFE0ambZaRaSebOVPZG0/Oc2HKTSekcfne3fE9Rd2VN6ZII90GYHNnasB
4jw/3WU43Dvfcfo2HYj6+O1c/iyAqFpknLGW+n8iYBIQ1g+FGX0wHa0GwRD/55AL
MmxrBr7kyo4uSaD/1yxW53dvBhktxI2Y1jXVGD2LMSTYIbJFuX6rSGuuALayyczk
D+lUa2P2VuReO6MA0aWi+I+EJJ9rbg4x59yapgNsRp2dW6FP5PQAJMEPwMsYnFXF
qBeWzhy/57q8V6fI/x/R9hB+lhiRp2SnRGKkZEmQ1f/lXvY8M4+NlglUvWWtvVgW
LU5PuKynYbsbRQXe83xSqyx6j+GG1J6rgmDB2Xd8Tp93UgkV/vRXmxpU/zW8Y6KC
gyAqwDtEHlqPimB18BrLpfxbhrOnyEJCPTiJCUnk2VBwh3MSOLoOkJFGy7sMdZd0
xfVf/PFuJTjvC6K1gsyakpCwD18UOjWRexOtU3RgyuyvajlDFNNzoDUbuP0lQOqk
QrdUIsF7J3cB2mTrWK3biT95fnFjZbRQexzeuzLWzbK84m45OkORSoGWlPcoRg+L
7hNaGoUmBuy98iCFighzzlUkHi7+Ri8sW/P+lu/m4r6+3CBIB3cZe9ya0+EEEisU
EeDKg9Zpyw4j1Uc0DfXSvCWvahsgFa9iJRdONdi499k5TFrn+wnHQn5BUlR2ZIKP
RWWYX3Fqa1lLV7wScT+IZigzRfAuolHRzmvC7Upy7MWVgd566AfkJF32b0S5UrM+
lJnFZHWEpstIuxEUej+PoA/nGmZmFq450vh7ofuYDaZRQ32UPm8FiJWIRNjS0hnn
cbQbS74DN8+bUn6TwM6AxiJmxe4o66fJO43EnafteEZ/vF7XLFPeMYukfvqygGTu
RvQcrs9XCaBbDyXshQ/OS/XwYTnMEaLO2iw6JyYB0a73XNnOVrnXrsFUEWOg/QgI
iX2Ih9uhGDcd4vYPMhmEgDLheJZpy6j0q9miZiJSoadiAIYHO5SvFNKDuKHVKD18
XiAJS1Fcs1s9I9BPzrZIY/d3ezXr0hpgNMKZ6uT319FQ/AP6fWsV6R6aPlTqZePG
95ZGr9ptCas7vAK7+41nHlh0hWR2CdlfxFsn2SUIdiMOr5IB1u4y6+Ejlyq/ZBOq
bkPTFA7epAF5aOA55lUTZhDck0+snVFEY2W1J5PV7qYFKHkWyfXvML4FmEnwUQjj
0VBA0bgALJQYIw+4GnG8PfA/IZlTGlioWIBiFNYHkYUNWfV6o4UTGrqK8mRJbb+W
BTdINJhyctiX8Ecms5bi0EJ/BWK8U7LRRKEVQcn1wr2xRgLRfSb55rOKjmpsNE3e
WiMSeY0BaXKjnNrTUPnmGekp4XU5Y8durXqrOSAujQdEzIROCD186rveV27oIDsG
ntUMZyCgtR4lY8SYp/Nwm6d5chsnyLYNf6nHmLLs9HW+vo4UidMpG7m0T2uANGlJ
5a8uBgONgo8DONipiaq93omLjpc2ehLcSCwZ198AnUYrQwttuLFzUJbJWbzj9Q77
PXDSmYcIWIx2Et9fUQgyRMXwVRIf3mHjWyT4C9lmmIOAvjHSjKndROHd3t0uLx6C
RtPsstbcKz4Ti0Q5xzuoOA0ji09bwui5TDrtgjyUp2PSh29KkcI9LYvy0OCAPQot
aE/KtEiyALqZGji25OpYoKApzCXA8Xjp2ata9EZ/JQqGVKHIK3lKAD4uC7lKRcHR
jorXXZYGKjDFaa/2Ha9crBYtaOQ34jCWKmrf266kKPJesihBz6xvj6iT51S7X4qP
HOqeuE5bWdrm5VFOoPpCRuGxo2qEUiuSwdRQud6dgD6Yzo4f90GYsurrOkol/V17
9fj1gSj/2RtaNPOksTHnLMq2RLKAQHJC3cR0Gm+78EZ3ZfyV3RxihVrHcWYEQX1o
UIvKYF4Dr1eHeqiEyq6q914lXYNDtuSxYGNhI6HRHlgAjtaRuH4ryz1d9hKx2O8w
lbutVfk+a/XLHZiDp9lGJYjenGyAq+Octeh3E8iG0p18mgl/cKgkj3k9hlXjgne/
PxMxaOzmdWzSjhFoNZAQmi1MnRpFChiQyuMgXCI8OyFShI0bSm9u6vHzSL2aBuf/
oNgFNkzfXF+7DPFLz7Ei4lHBYZNEHx5YkGc3Z2/hSJFv3QE2oai3VwzSWoN12O8g
URs6TEV046pgKateAc6+AXMp224u5HxNuX7vHIZCangTqn26fM4YrhceoQwGw5Ai
aGEdaUWmeKgarvYDPn/5G71Cql/77oJJzAznicX6kQGMpTqE6ZkwW++fwZAvlTpz
8zH2bRiE9N964jD3xv/fNZa1C9hG6gdTPAV56kgmX1tqOOoMCFQczItGNSNWMNFh
fUnaIXNai1KoSf1Yv3qFSHSIRsmDndDBU/Us2enMiJNBtOqGCjfX4U5sgJDJboUG
s2mf5BRPoCs5g4lTueQxrvwBu+4wWu8PSBJYWlgos0UNA0ljrt5qwvj7IOLd0NAa
JsF35Cv+F/tim9TIaFrGpDtK0iuj+CiTWW8C4yi/2SpHElncaDCUrU67vlJBnCiT
hud8svprQwPxLIhOSyKdQAgsTdorQDaRC/3g07d7Ap0SPP3f8uHXMRE5YpohQ/Gu
Il6/JWTx0/i/M+ldJHpyIZAfn3sHX6bAmooVHKzCS9OMZpLQNO22MZWLXG0a9UNr
/SppIsa3TsvvZcvL6hC17sKaw5c6As/ln3dIWWAtyr9g64YRlGUk+PQuQrhPovb4
wjRvpP0B32h10fWaRoC3vrn16LPFU28fd+bSex9JMlSBweBWChe4NXz+P/7OyW5C
Aoz+EPAhHWr5WUaf+VloPTDKXSw5m22PlELtzhjRfX9DVwYc5yKL0YOm/eV4W5oU
IIXjJDNWrZlKpRO+LGqdFESZM071Dwpq6aH0791LIqzT89S6JMOyAejZ1jJmtq1p
mPgjbOsc1WITG8wabt1YKzr1B/xMPaCVK6hI1gSme9rjIBptt93UEbR7MeVewLmd
vt6WHGeZS8zmSOw+eL7F8Jkm5vW0CCbg2zPmTBJv6rmn9pwjpPDftRW1FghOet86
Ingb8r9MX78ySNlGKN8l3jIf7OIQ2EU9OmJQ/co1LWhTTp8ggHcb6K5vUfWbEr4d
YDdDFkNP4CU9oJxTdrp2C8yTHBnP6t2Vnv1czHGSCpdAGkrFy0AgVbguEAu27YsP
dzG3PyRQbF4SNwP1X0/eUzK2uf1Tz90aHqCUQauxAVrx+zUg50P33ou966dQnW7N
sOvmcHz78kKTZ9Bm+NkthAeeMH9t+ZlWKm00E6HVLhGpCVGno7nhuXy8V5vo+fBs
8OR/q7snMjfNT6//rHVqP1qTy4vrcZPZQGWNbXYc1xvH8Oi//o4ONY6+EwecmA1K
kmle08xgmgtRNPj7FIv9nfWTqwYpr/o/Ilqx+lrqaW3v3Ho4LsXyBNYLqtkh9a8P
E8JXwmcip4TfE0HtWLqLxRbMfK752LZNPZpGKxAU2bnop8PEBk3lvIJgK8zffZ4U
fbuXxjFEk9OqaJoO2REGbjZG9DL4UTFaPxCuPFUL5qmDcaxC45qBeWIxqAMuMg8p
S5cftsbXVYqMMAw1fwVqfzV2FOI1kSvpWtkqVz3nARq7vHXAD98fw9hUTaXNY5zg
sWTu3Db0skYxP9VRYYv7IpS+ctJrl0E7CkP05OhnKqZo2WO10RWcRQ60+OwQ25cQ
ILXLIAJUB8yfbElWqWe/H1eDG8xF6PxFtycvGBsLh+QUliLEHBnZE0cOOJS+LfKn
pHMhCJQEV00CuIiVBtnu4I0C1uxSCmsu3gYHWVHKayvVHdWx+3ShFpxBgLUnhZ/r
AckARAlUSct27HmyL+DWDWDm0ovOkp5kgdSiYSLy6JyRHkObv5G4wbghXBIWmzVP
fBFwFwVunFRBOKhg7tVDFDuZGR4FBKpKSLJXDPzShfbvMP9Sd6MT/R+103Lc/Ksi
Gt3BFVU0vzXd0+W0Y49s1+T3Qf8VcpE/kfrv0ZbinpWuAqWun9AYU46bK5v5/JXj
7FtyLR4WR/2B+3B94Pe9FkTcp6NbXJl6J905xz3khjLLNvIVdwmOJ5n8J6+86RuL
V/ufgcmsvbcxABxpLxJJ5cmpWe4GR6OVW8jA5zRS3ypXwe2wmF3Rz5GFYHWOnnAq
dtkHlmwcU3Zmf/YzQnyn+8ItVD6TDgkZpzv71eB6BQ+tvLJBhLnp9rLPfZ2fdyiK
RMuMxFwm3Yb+Ws8fJ4DcRXWznTJIADtDIkaAnVfk7RF2fix5lgdrdy/ZKMYV+5ke
QaVCXFpZjwRtAAUNTWYiKx48qzriRdtnKSdIa39JRm8HYC680e3M8kdRw9TRQ8c9
FCmFpfUQ6v6yMMnRJjULg0TonlEKL76s0A/cXFnrO8ibQ5A8x2tPLdiGI6rP9loD
VgMlcjP3oF7NOeuIdKOh2l7yDR5Cr3falPPY9vWsv/nn8noIVYxTmrDAL0/2e6jU
/wtxBU/H+qHm9BFeG+OE70FotlRFhedWHc6/WH6IcGjOmDPnk3x9glwFSX+XG3jT
dHlk15O3Z+skeQluCKNS18TUSZ6NkZjP+66p6qrdIU9sTbw2eVjI5oMgTC5EKzGw
YbCZt1eKboDosWdSmC31LXu4pe4f8erDfEMVAEff29J4at6lJzjyLIu1vJ4bxKEp
iZQUUGzUXc4nJh+NEXmonrT7jtvz1o7S80UIqBYpxfwEOZSvBkTwaDPpoDkJdvSc
hhN9uCdFvEetpd26rwBzcuKmGM5tHmQUzagoj8M7KdAw0ycr3GIre3nVfvaUKPx3
zbyVuvETaVJAdUCvK2qZUaiYQYIBuOWxHDavHoEzTuzmn06UvH08yBbXSWiz3y3I
HIyugvcQKj31dEw1mDO8y3d0/NfnnvIksuXups9BCfBmAZ3GOlJ0WdlkSQ28ka2R
NIem8LXEj/2Ve1vYMJYN9Aw3AKHwQMrbAzjru7OjlOMVQrkyx5/MalGIo/TPGLL9
jbvYiQ/VkMsnMjm6hc3vRmYQT7dekn6U3o16nsw/QsW75T6pM0t/clXpNJ6seeFh
fHic0FhmHO4WOE/LFuP/WD5QEjR13BTGpuNM5axCPp05nIwTl3QB5XOn1q+A06o5
d1amo83/GwcIdWldKeQi7/GG9xb2Wx2fu1YbXfqp4JfRsLheytdjqUAmtfNWphdu
2zyNMkRTGt7IWSbGC8P4nG6SBxX24yojDAOJqXp9oc7G7tSG/NH9uuENbq2uM+4Z
3SR6za2gEMogSOGoZEp++CuNu8G8y4284MIy/0bfRjBRxfU5kFGLuJJRtzkS0S1n
iCw0N7aqY3Y3iM5MVzYT9J4t9zi7QsXLtJJBtVol42sPGNN/3Shs6NkhC0qcFfTI
BwrAzA4mitH402kHFgqCLilit4dayA+z8EcE2S27q7EI7wxGd4B8fgU4Qx7xzuOs
tIrZpNxq8GjBOduVaxcSiosT2nAUUwiSmEbfE91WgScGC/CCJcwmCFyL47R4IgRQ
WqMnx75CoPoEjcQEXVdt9P1NFi6oDyKFoEGOXrY7SYNsO0F6Ihagl5ItOawDUnaF
bRkfXvEMIilTjg5pKWTqgTFQXPuNi3lc+ezK9rzMv9brqJiigpoE+aNsA6lB/rmA
ZHLvxSIgUz5vQ+gEiR+06NWuXPDewABTcnVdehciKZVMXvlZYP8vpxcTgitScbR2
XRyhRt0lKKnadOwtInhGFQGu4VmPGUU8D7fuy10iXprZIy4yiLciTAWVYPYOK7Nb
kl1TXpnntUv+Ia9UaB3C4urjqvBGrtEr6wDWenfNNM9LgNg9WJxgmYG7/08rtA6A
K/chP8PiQJodkNB1HWUSTm+XhZHuc7vd0wsuCIKLSlhlVGdhZTuFTg2fVv/iTje3
F6hDvN2Ni0KW/rPqat4+YDrNRIo5Y1GqunX7u7ajLzwXCA4MtLa+8tG46VlL0I64
z7s7MZW9cPQd0S8joMtTKFiaMLyvlJHFdpI8Gm+jUbzq49pfrVBV+m5wROA20XRC
eea48EZmZHiwguDkX0S1fIDxIPUmfkAR6X2ECJakso9Hi/KfT9Ld+PTV7so2/0tQ
W6ymERKY5X2THuyT4sJtprFIIk5Gwsc6nHLYRF6JRAYp6hgCdqUXE2fZ63jmc875
lykdac3HMBc5yoEfI1HXGzJKPkgSzaBHfek/TolYNjoSKzPtuf6mkJI4tP+zYQfS
Gy2qTLMRckCo7lAEndJPf3R+pzA/KGhrvyG7gAjoMH79dhhFiEvPBSwD69Qckm6w
bTMJz4yzZmxP1R/TNP5BHjnXTlm5kZpGvvlYlJ1IA1eaZsj4TuYkOyRZEmclh7qp
J95NaXVyXrUgoHZvzGZJ65MbIhIKHeYUzR/GMFN5/nKvn27atg3Yw3730bCqIOD1
RzRhkX5znecMMT84hXhG1wg0ce6dW+gRvwY8yg+y8+kAuc4f7YpjNsr0wcxGdjyC
YMi4oVFIokjSe2KqCKu7z/mKoIFIb3RRjJeeQVzuBPYx6DYDyCmbGirrU9omblF/
WdZW0VAaUQl71Keh5h8SIirADc2d+Tsk+ccDe0tg/SOyv+ZMR8OMFbv+MKjNrQxz
Bk9acLmrj/hicaMcHUhyTBpL5ZbR7bv2VH2SdAEMqeEJVLMfUyQOnGkfMkoVd+Vl
6Sk+VDcHMXNMMtwuD7vY20JNlFBDEGHLPAf7PhsHbj4hWqp1N4AW2lFuv6B1+DuN
NZzeOJN+0tj+hwMi4aWRFyf7GbRc7kW8qFfWYKOnC1V2tTxo/Rn+2616hVzriDGQ
RJjySnT8xTTl/7qOtlVYtjnaNUnQ28HNzBSMtOzyCwDEmb5WSmpR83NN74n77ssE
Grzf72D4gDJrZjKmeSP6MiVVzjRRvJf/6pek6liOxg/DCxGsRIvzSpiz2FQMf0Oo
ES4lB9L5I+/F8ZJGu8Ck9TaHjLW8tjRb0pgLqiskurBoWXIhsolAr+07bA5MzmDl
eXs7wMjwDBpsQEbJOOiMtksayPNokzTkJ1Po/yVJAcTNEPc0Ux8eD92kF6m7BSXW
ROBUuoQNC9/NHiVY+SvAIHFWGpGJcfwcay0BClUznDnMOlwKSYwc50YgeoSIbHK7
nHxAMIngEvAfipqvvMDMQXGYQxyBm/9CeeoPzAzIWuCU/xznnb9AeXSKBKUgGlTn
lLubEyfRqT5O37VsLg1bpOKbHmtMmlcs++Opy0G67XMuU24DwhxIchXXuLguTw1p
0SdaJdJp+QIra2I6gMzLjeWmQaekOJZzLjKQxx9mw/fx6svHmuN9Lz7EgAKbfxHX
ZxfbPJxsTeDzhccW7KiO+2raOg7Ws1Km7VL12gieelSE33C/Jt9YjSF0Pr0qvLP5
td6LPgY8tDfvptR67nepW03DCb3g9yz8YMJl9YtLotX2N13YveNx6iE/Mu9UQzRq
FgWr64rJ6+SMPttfz7vr2ywpTOYPpEUtEZB2V+I2tWSgCesF5M7f1qXYn20wUWo2
EvawoKpMztnDCC9VahbJ0vHyQjhlWzEokUtJrc5I21gQ8KlYfvfLHIQaoK0htwAT
MjHsxfHcAnIbGEI7RChp6g8iUny2XtoqsUukcg+wnvFJRawc2pv223BJHm0uu64K
DzOZFtz2dYmK2RsqwrqlZOE2aPnUfIIZOb3FamfPgebVyJiUQlNaKdNDNVl1avy7
1YJ6zUnqjNyh2iOrgJ2SdZ+6y61pNq1PhbRpVbKqJXkXJHADC2MEJrlDsB21BGw+
yFvDU/rP80Ygf7AqyYqHD5mL4+P9ON4Qf5Xo/LPzsLRiSqi38H7SNeal/ImUgUVo
uWDnHLGrHGf4fNzrgm5g8cEfRr1qRucEEXqtZHtyeYmlbhr/Tz8v+x+wwQSRSDOY
8EYuVbMQgEadNGqw3eOCIoD1zAyl9ABTX5n3vc/W/5TIKIcBtD001vYHEr2PwGm1
pEJ1h5G9/dGMp5wiM7zKjZPi9gIykUJ0jM/+w5T6ehzisZHXaTLRjJYvyDopgaHL
6m3VijV+MloHJ+pG8ylughbhuHehJso1jyjY4bQtARyl5VHJ5B5832nv0ZtC3pIC
YJEiN3ew3lasWIZ5A/9TIIbF2UpWpibpqw4D3rDxx+mWH+s0prXzZ0JJlQzcXaB1
Hw5f7ZICBlAdNCsW9PASf0oc6KhBfgUiiyp5QtUja+4tB+r2wngonnfLOi3e707K
Jm9nRrkLEgyKtrRIh/We9eJd26eLcVbve2TLjcpIcyo=
`pragma protect end_protected
