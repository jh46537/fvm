// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
s7/qrSpzOyjfK8ntiIi/QYLCiuauZR2BeNyeBEnVLclGS9kaC6zlF+HI7LSY8tsl
cJ7jK5al0YjpFFe1yas8S3lWzr+/RIM2iTDtFHTUS+ijfxCgHGaPWkRZQ6AprJNs
eFnequuq5eIKECuKSKUURm9JYPkZfbi5v2iXmmufiNk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6848)
QUY5r7WnjqS5R1DNyvfF/qwS0TImyYJlvT7icsYb2N1N8tcAAw9y7EvToG90TR32
Bl+24yafawMvtpvThF+m7cbNhsufqkRY3ZNE7s8ihclzpWgCqCKi82kE5DBXcc5i
qKLApBXeuarN6qb4z4nEIqNywRn1kYjRofYvnuAzafm7xTlJrrWqYhFzPXlcxcIM
y4+TBp8hcMogKQ+Zk21ZgxwhJI6Iv2L7KEDESg3mziio786MEVcnqsbhj9ZRA2l9
fGpZXeqS2M54r63gYeRawH6itJ0adtqB7JMlSbazEvJPXbeSZwkD1xSFIz1XPJtK
DC/3SjVK6WzTp2i4CnS0TqPXgEMbeF5gAccY83xw1DrnVRiDORXP9tD2oSW45DYJ
ttGJJ1ZOrJL5Wrp0g+wcXy+hzmKG+r83dtl+qCyRy254sYovjWyf7Ck0B/40P/Yy
bUVcLwR+4Opl/RqjJ8OH3oRx5Nq9EixyN1OEIFOhP7nofUNzhs2wnTX+0u7X2uTi
tbmHbku0jGWl7syLJPhsRuVUpfnyXM2Shit8u6xJDzhLkxUlvF0ZN43wrRl+Bwz9
gP2m+4Bkg6xnyvJJ7ms18MKP/JwL0zZI4bpW93dFEtc8CekpUdFW3Pj5yt8CGA/f
wDgyTKR/B1wSL7U7l3nbdGLBiiAPHdHl2VFg2HcI7kyKSYASLvcTrVU2gu6VXT6s
3TZeFqX3d4fcjgGX3m/l3EdclZj2gSRUcb+No3M/sDvGKbsNSa+eRaHxORLNFyXx
8KdYA5MykjAms2tsP6hCDSTrGKv7RJiyrjEkX46/ejp8AQLUDRiMi45l098jsq/4
tMT9AKW6CfZtoUGp3rWNIh2loEF2F24FJ7kk0gRKTgCSc1eB0U76Q2DP8K63B7qA
38awFElw5xMvD+yr/XRpeEOvKjPw1MOpddJuLXLS90zz7OXOoveD40Rnx6MvSyFx
zniOCMxRo7rf8F8Fofda/e+9JjHozA+nlZMLy8pmUZpVMSiec8VjtlpXlPFeaoL5
pYqyJ+qTgfW86B3gLbnfOxthhecnXMecXBrhAro8v85SBfDbRiE0wOeyDs8JFp0+
7LdjeAWwkMxWCiUS0BIr6KRY/dTut3gnZjeu63UHuyhUx+uCbjpPT4vAbsrpFK6g
uqaLBWY5q8PG53WEA2yme51023xs88i2AfbwmlbU9RIClqwY7GEEVwlu0RpnT6AW
EcY7Xs59JRrD+2g6u7zejcZRS0JNJYud8DcCiWDZYvBYyQe6iymAAQqPRgAtYU22
2YlnKUaz/iAPvSBeP+utmdtRx/ZpX69PJUm80d1FqKVM+K7hydIuUgHsDRu97cUC
uDuJl/BaT5t0a2ggBT1Z/tTnVxZThEV5Pm10opt7Pp0t1xom0OTQ+49y7SvO03kG
hxkxlVSfSGe4pYi3o7MUs5f5tQ3k784p+NC31wMkg6Ps3Mdj3J5Ph0A/prvc8BLc
ABvZ9sFM4ElSYVlHlQn3qMrP2s/k6F4g5oywD5D5ZgFyztTczaxe+kEdKQFMAWYc
aEPSOWGPWrTJ8soBun75Q02QeHqwgnJ0peeElZsyBCY4N+iKfj3HejT8IAQYfs2h
8N1YPHud1HVz5OoS4U12eDlq7+rnzG9F6+8lPCkuT2AFF8nZMqFToZyD/lt+ic8/
1Nts+D6Cc659RpSCWXvQPys7uetR5dnRtPMXbRc8pR3beaWUOlm0rJvTSghE4HW+
OJ3VGa6aU+4ILos0z0tpkUd9Pgvkfp1HAjF6ZWZ+6G3D6Ep33U1OFtxFXkzv30xj
ark13pjUbBLcYdEF/HCjB7dXRMxWm2CI6ijV34kDRao6J7eCelGHJeoMYFxIaQuT
hQIB3J/Xdnt7o4uymAjEimehEdCWfBWcLLrgdS2zK6hOFIQjHaWb5kRXW2HuStdZ
4z4NoGDqcnwNMkrgHhiOcbq3cWuE6pka8HtqYZAcKHb8+9e3p/LL835oV/6YKWbk
sOsaefsNqqgmAoEt/+f7mnPd1bJH3tafvbEjjugNrVM6U6tlniY9JWrZrkD1ep5e
7GHJIHh1uNch5WGX7d9mtme3UB5BmBJvClHxAsettGVnYcyE6nt7T51gmMBEAXqE
UecTEZiYrlqBHKCqO3yTuEj0vkd1uchHkWitXxpnihkYcdkDIYzfmcBWWR/owr9w
2atjOu9tzcpPU1FmJFo1mIwuPvVwOBT2kRIo4qxjdSlb7gecvP6yQXQpvHGmrVea
iq3zdyO62zNAC9KTQlaOWHX/D0lDGWlJMp/D02Xorc6B6R3qqW0meuufgck1wwij
k3ykoWN2juJnjyoNvRqAoK7F9SIEVWBm4GvUaKXovP8vuIJRH8KdS+0tKR4TePPD
VFgEOoE+KG0COQYgYcCF1L9rhUhHpPm3Q8F+LIl/2N9sFwDBPtaVB0aanAbEjMNA
yNBoS/9kuY9z7DWRQhxZ04FTH1XDWGkadzKF1J8u8mPn8+qVJkZrFwl066g3O41p
mTETn/Y99U9p6CEmxeEh/VgpWD1plZJ7GZw+jiSKyRp6m2SAW4MI7LefVPdQ3PE2
N/tUHSUfT5pHFh7wm9Ip4BJgwWjpJXM5ql4Cn+V1AfpUUQTsiLXT0wfQ9DooGze7
1/YLE7YoCcVbaXpA7M3Ff5TEQ2pxO7ziTKyinIKKvHaaSGb1sjUpkHyeVBHIsb2q
NTiN1Xcwiu7rxbvg1wEZgz4U6xbtvCKsgNfQW7rea8GoT/UT8SJtR+uYKR8ohCKS
hwcqahJFc0G912aeccGCqYhN6nRqvraJ9eA7dLRHCMFokzPpRvlEbhOGNEbOfwW9
aZ5ZFlQLl8RpVaH4P/8BE7UE5LHipywPg1wIP+tVJl48LyaJ3qu/OAlRcsObX4HW
0lid0OBEHTlE2jX802Ba7bO6BvVTsJsUfQmbOGT0p/eGJvnFQ0/j/OU0dDlbXjYO
rKq/l6oLQYjk7ix5/WdmUzms3erH8dbhZY2AasEzmSNIQXLq5c6A+BO3OQswzkq1
ms8VTfqAvNtyyud5+qrwMu0ll6dDRh33zQzgXRhyzx0/Eg8UAYHdLJHTKm/nlyHT
dz04oxSSj/A/oNi5P6X2q2EkxqNWpDGhpZ6b6qXFKjNzWSeQzk5VR5w8FGZxXuJG
E1qRzSmgZgWv9bcHL26fd9v0up9EguBDdiqQqEEgawtVuewujlYbucY/c7AvyhJW
BM+9ddE1gOB4Hxp2W+E7xItSjed+8oNxZENwleJ4OGAl9TYdKwVdIgIgCI+GXX9Z
27AsHkkk/AXogilsdOw1D1iesfqAcUzLUzjRGV1cHAnaMO9zBIMtqUUxc7HOUHdD
S1Z9D43VcfQkyHIiSisa/d6Ojjod3AyS74JIvfljUO3f3tvVA1PuPXBJwm4aVq5v
kIkWbIJQZkZTtTeV/dnNfa5n5JNIEXPtO8rAJ/ObYeTHk2wuOotS3pXyt4V2EPfZ
tTI5FIzfJJAQwGR5qxLiPKrGLh3dzO0dVC2TgtsBT3t7rj4ZbnvpVeGwl9WYeC9u
8geCpbZ6HsQE3JFAntBqbF0XIrtpRS6rG3rttHoxPkIxuLoyS4sgD5PgohQHH/XS
WMtp+1Eo6XMnhBAcs2lKglzPzzhi5WCr9zjNv1IaCsbWliL45YwRQf56Jvk+nKL4
IrL7G5Igu0ROwhmCWX+i4paAUCvQL3ToLJcRdvqYKwEwaX0n7eLOTP0oWVcWiNXR
C9uKMgE8zlZfOGYN7601JM2hY1e1mV5s5a/Qe2eKfx6yUZoua9ySU2T0TSMbgGBr
m2go5fugyIHK+j0IW94bGt02KY6iahJSp1iijl9il1/CSpCNB/oYtW/LysbcjisG
QQpztyq7wbtuttw1oq+sZrdAHMI9Kkpy4NEM7L6dF9q+kO0Ga+BAzGZSWoupwlqW
yQR4ckHfxfeJGN8R2lGffp3Iuj4wkvODqZMI1lx3H8p/JbzF6jS0KyuboPLK76W1
rp5QZiJj/jW7bUprkCZOiV+gtPV8eZoR421hYAu6lYhbdWSX8GgRblaJ+6lv+rIX
GX/A6hkVx6XiXZ2724LFnosVQH1MshV2V0luVwMpysetU0pdFRkGEufdRe8+dhMj
8UgcSBxxr+fFluP1i2AfGKVL6J4VcX9qpkMWxX0Jlo3R0ZcwYpDRaxKbWw/sbQbo
hkX23Pagbe4LHJ3EYbgaMLdW3U/SgXZtwsMFAsEQd6Tj8EqtSaDJj8ewKryqrcWA
3aLnIG3ck7PWoiRCaCyDB2pSO6/1K80UA5KflvEKH4yKMSX646rjjCnwM57yj2n7
AJh+9FAaD5uwlwf0dL/J4tc3MaPmq0rw5vivrpp/yafhfSSezOKrBKns7pdbowAV
nrV751aiHYr2CwFD2umtCtE4/nx4N06oH1aQdwVEuaLzKnqzyzXpWWY1nxBY9TDw
ElHv11GmSz3pnW3sdjUgxwqSuz4SSZXEJfWs7jSAVXOObF0I/oTvTO8ncy1KQ/bm
7T2l8dNm7VLaqokZiQkmk4a2T/La9Tw488kWTFfyYdzG9OnLJms1W+6/DIEOhd1+
XP14jTBCMdgf+dMNR7P1372zQhyMH/6w3C4l4CXcFKktbSXZgwcfjbdcMdKbGACs
3jWe2fiCX0XmMTCeMLXmd/8g6FG4cW/9imw3q88Ksz+WMxaTp5vwTVzQ7p+mjVaQ
41YTLFZIphveuldw/V0KSL8g5WM1g6MkZIJclLI4x+/bzZ7H8+zE0YvAd9ShIcr9
Mwo7G4ToBmmxg9kQp4uYREVyTVIu8AfDBWXzknUxKICKqb+ZtNlbhHWv1pSU/tSH
Z8DEm5m9pnBjmhb8b6kBBmN7m8qZ3DtRQf5K2iE8cSyDsid0tvXvBJERMDf6k+IQ
JglNBfY2DvwrWQzTw1CjTqGiEsPsKQgmK3eqdfqZjl/CX2s8R9n1+NN1e3TlkH6L
plYOYw4+AjRfNMG6QMkhsrfHjza/l31LcFYvesX/yPQzrmK4mbrxZN93eEC3Mv19
AcGbtwU+1gcCrgbCpNjhTDKXpgagLqtsz6Ooww6rcJhzD0scrT4S3xl4fwhZf/CK
LijYdkST5eNJMy1vXiNdJeNhLsLA9FFvCLFTNPcb46QfwfYGg2QoQ+mEI2t+A+Ak
EoApM1BMKOp8e5sV2nZQ6FROi6t+7BV2B08CVVNPlYr1G7JWm7gu6C8qeNoV/vVv
nOw9bGsfCjILLcHAIj2pMWpP964U334ATV6dTFKEaPgAL86cxhYEryaUdGlI78xO
GH8qBh60jKoBk7lS0RdpOxvJs6A3P0pY2utf0JhOHPDSe8yxJNCi8BKZWR3iv/qb
w52DSAXx119JEyjPcFEFABDDDyl2Ei9GUeNJPIaKyTbUK38CP8SsSH40TuVv452z
MUV3lGQfLotUz8bNSlISpH1J94oWj6nXnsmkhF3WLG7sk06Rj1mJmLgwLeCOV/ER
SOQWFYA/K937N8Bt0sqfKpIzuHeAnwtPGHgVHcrUWrnEjAu/h/gSh7UZhzBiiWaK
iHyN2tgtrHT0Pim7MCUlNXletRhaRl5itzEswZRuLIjOMH01Te69PRe1nxKzxoaA
w58DXyovSyIVATtMA0qmMsYn/kETpkaTatNWPRP8bR7LzkLGj7w2BTj/ipv2KDWZ
d511FjqjYZ+u6kWTdvLSOZSz24+dOuynSfMuUiVqiYhQZPBIYqYwuGpKQjVkvrLQ
/Iw9xs44ZhaigQ6fTkc77Mn9/xx4JRtMzJKd1SCeN2briHFVV5mEirfK9kzo12iq
jAXyB3Z1HF3N2qre8Ofy+x5rmbyyp5x3wzMI9v/E6igO3zohEpjcr7ALCSY6QEX+
Bj5IbplKiTX/mCJss+D4d8zR4fyDe0KPFsiPNqD56FwztRZSz6XJGYpQp+qM41Nk
PdeV9TY9NIlH5qySQwFac9qtFyN9ocj51Yh5wU/3ejXj8iia32rSnZ738y9qytMZ
GBRmLy7zYB6CQ0HZn0oL7+a4rfa1UjBUY1eAuyXw+EAsruZ9dmjoYLp5IScoIc+J
Ft4BzCOW/oP3H3eN7E7D6z07ZBYHkJ4gUqpNapFfuGCqQ5qnB9qo3IIOcVieaWRF
LvvKATe6bsDEtdOOehkFxuOddI4Yy7dUehsSwnBu3BSxrYyHrYKnk+VXyxqwjAxV
MIiYCoqGI7PdoKYnPDK+I/e77C66BbEGiPIO8eGkkOA8A+dFKU5G+j41GryV9cVk
QMk0z/JJHUJgeSnckUCBRiJdHTJxwteXopGAAY16GaNK1RB8h7PZqI38L/+vvSNu
HTqtuYdSzI+J8e6x6IVFsSHcKAEcRdCNNfLBeGeS/bxuv/oCd28ntN5QxYYzLqs1
vpRGud1oCm8jnuIIwM32q626PFv+GnTYqqTBFooE2B9LcXqo6GcBbFmrOBmpnxJf
l+8aJIzZDzJlDvRtHPJ8ki8BWHpRKNA8v/rMNuagvku2zFzOFFQskKtE5YxEvXLn
KpG1iRCJguDbWTJbAODVaVY4WzxhzOPOaEkcykH+xjAGD5NZBklJuV34TSCSVgB+
S8uwxrg8Ob5Odc557dbaOlpPnuzT2QwLEMUmFHBbFIqrH2fYn4zMRula0Wadx7Kt
PqJByHuRXQozT9q4r/i7lhixyYs/dnOGI27yQKZuHxLfZVnXUGMOOsP0PeAykzkU
x1hGZSs/9vHggEcDlDy+MigzuISWNx1m/Fkeo3RSCadKP+21DPZzynsL7Dv5QUwH
YNzsUxMGQfALykUW/K5pKe3TN4UP3oak++YvokhtHw2o4EBuFvjYQOd675lWqTuI
T/kDDYXB5CqJs8kmW6/l18Es5IDt6UuJWdJVX4/t6/AxgrLYDRwR/13O7hGLWrze
tpo8+rtMpwwP4NkwMVdBFtxHvwMHYUS9WnGV0beRmu0CQQXDl+YuEySWnmF6EA2y
acFNRQbaqGRuYCXpM5azuudB35Ero3Al/bYil6ev531mbpZp0ycf0pUBIhR1gBV+
236OUCxRvLE1MGpBwnE1gkKkanu3d+9i9Sw3nJBeXhLe7AWMVvyNKZZtB0TzYsvp
uFvZev+ZF7O/9Q9TJQxvt5KmvIhWNTqp5g7wyZr+DP6KMiX0b6RCX1FlcQPhGmM0
orrd3AabjMIg6OvKRMyAgM5Tih9+MENYt9K+WtqzksRm75SLh+4B/LeAPUYQ1ANb
V1gRusjuHMDyJDA7XPcD+Z/uRSOLuMbnmVTJ3Ztr8TPEO75z/ouVOxKyI9qOmzGF
Au0Zffxwfvl0sP/SrN5mM14+yTJXhbhWtQAhv1OiGAb5uF+EQ2efSy5q9jP7nGs4
lXiV+ag6zDsgJc0Mch6vanvF3y2y+A1I4eeuQEQ/tmBrt1ABi9LLyORVX3wXg7zl
yHmCoXeVBmKYcyTiTSYJDvxtIQ+UOXxtBZlI6VTUrzwmgR0K6AXDM4K8+yaWCLag
b1aqRlYGJuNZvQjv0N9rbYrCpCXjnZNZnShiezHB+E+V8BZMkp+fnZ/Rjl12bwXK
bkmkcPWk4UMe+/oUh7+R0JjujM6hWXcTBsj7WAxsgSfpeaFz6phNEBTaRpJxMUPc
2QptLG0cjZeIHD0pDuPHnJd2eUb4+Yq9q2CrVmhbYyjGrw3+JD6QJN64t8M83JZ9
LJmGGbBg8VaT1pbAD4vLA2Fub7j7rmLGpqBS3Dncydi7qcv0jh5ocKiipkiEZ/P3
GOGkZdcwAkT6mw0p8aKkiY3n3FV+w5PnO0hfvXvbgBmYZMlG5rXkSwGYvteLH6B4
+nNh64lRZX9CFsJbwkQIVGvHv091oxaDMlfvthGHWD1QTrrYJ4qcHoSQH6GJvwpq
lpo/pQO4jycN8IQAPwNmcVJZ4Powh3u3ekmI/TCGVvjqXmWoyIGgKxH2Fk7+iVp7
oqyIwKA3RZphstzqdfb9HwwRr93eKP+q2N5GahAF2M1A2TMHi9qj0HMbcis7GuhS
w5NkqUdspm+i7EzV8dRlbjESat4qn+pB+0NDw+rv+mRdb80hE1jdqnnbwXo44JgT
yVJI92MZtTPGvRQ9a2NF76gCrVIfHBCs6ev5gAHKzSS7P4h9+uv/O+1XJaat68NQ
4rZqYHgZlK+9jc3pRdH/MUqefzTJMHwUf2QinuCsJeiJ/d6bYB0OG3J10Pl8XZ3c
l663WHyLavZ7YY06titjH2pZ6jDll+OF/tk5tp7ZOK0Q9nirILjTY/9nv+XkWAD1
/cYkcVIN4K7m87HF4KDu4gaej2k9dpdruOupVRbledyTzxgBxtbCtyyMWp7+D63g
9g2A5viVELC7XPjB2qnfhvjagXNZQ+XqHFthlKD3VWlNN4cD+qqsFopVQAJCHSR9
uZRVZJYkCnd3XQKJy4TbSe+tak5sTfU+cNJ+Cd1+fzEm4wM7g5CfpIsog+qtzEkR
LwbXvPkN4yBjPpBsKbs4d2tKJegiNsbH4Zkg3M0gFGySLjobuCnquNAej0GqzltV
tJNooJRO/GxbIsxB8eDTa2dWfEvQXgGXEK6xa4RuQ6G6GrkSMq+tNYFzqP/i3iV0
G/M+jiYcDG66HS7Ft3PFzEIxchKMXxwe6P9mndLFse88CutGwL0ReY8TRKONEMSX
rO4q+SNSLfTsdvE7hd/Py/YokLywPK2h9+40SQ7Vmg8hxjTiRK5w7+LdL/XL0DQ9
etuHgoGMLIiOXymMsyP1ylGcfgLApZnVWgSwXKnPPw+n6kzfim+rrHTr7QD2rI4q
uGpNq3+5PjKUsFpRexn2yHBhzwNZG53m8g4PGISIOmHmP34vm/AIsv1+lc1u6gLz
lThC0dioRAvOUeTRr7FP2Jkg5qy6jrW/eKiTXoJQ0DgM10s/P0oV/WywXvnXxaqe
0O2dlyGD7Mt3XuXsT8ScdZsLJUorHHH+SxDr7lJ3o34TJlKZLoPaia13rsJ+l72+
MtY96rcg6Xw7xa/NbZyg2d8aIOjmaA8ymaNurktwiwWWbpEnsMlXGwrapDkonNV2
8KVVMqBFPNjTrn700t/GaoIGsO5c+1dENZB2Qp1K4MT1s8fK8QHG940JJeODM8me
uz3pu0MajoT8gmcU2qMauIqHiiELQoftMhVw169kLWRUx7pO/N+B2I34NIH8xl1l
1DzrpKCgXbMgtVPjp0m336bx2UYDQ4/cm6Am2ZI/g8g=
`pragma protect end_protected
