// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
S86ptg4Eypr4VeszXEAj16w6/frcsqw5DzGQ5YSUowED+c8qvg12V5IB9bNaW0kW
aeSLgZXbZfMIf47vZ+sAwtmcC5C752I99IlSW2Dd9grS4WL10ibRzdAArdXrDiHk
16nyaHMH7x8buDWB9bAQrea7JhRGO6mL31/3UGRfxoc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17408)
EJkrF7qn1FtxMHuy0TLF+G81jnGilO8n2So2uMxe6biZ837b9udXes6KZjQRQ9lL
ziv5d1MbUCOQhzWgUkdPmkrHFhwFcXdL4ZKvoPvGXxkeKMQVP/pHFuEaiP3AUsuU
hv1xnSvZJmJAnw8rPzcO5E+YjLA4tXV0Qn8dIrliWsFoAdbNSoT9aC0I4A1cRM59
6zu3099SzU6p+IVztMOWIJMNUjWmEyADlXDXfTK0Mcmr6Rl8FQzsMVX4IwZP+nWj
j+EAkjMtKAhT4lDEmk3ieQFpnr4DmjzScD+WzMCdI+sVx0i2R/Q9BLh4H+X0Msux
qA6AIwV/F2BiLJeBtqCYWTXMSONSWPoISN3PNgxyr/NGIPuyofklAvYOYzDDvPtS
mGtNKlC+zcpw5lVdGFlf8xc7DkY6QJivNr3HOhEcD0douTksvKAHDo4+KJ0ilMlK
CkXe5TAPI8hGBdjNM5YMtJCdPFt2jHY4zn+IH9GTryo6Sm/Bc1EBTR2et/2l6mz4
AAgGswv4s2ungxuxcmMLqB748wXTn1KW6AnntVDs3vckBY6BmVCeHrJC4WbKShzO
kLUH4AGT3sdpdeF6/CvwChzGUkUcacU/DJya5CiPvFDFLvDO9XbMIHjrShK5AtZm
c9dGnfVYxKepMu3DsUMp7mHKJ9BMfyEp3MbHr0hcKLRZIWfGHxuplinuMA/W3d/z
QkOPs+hK+buXHwBG5r5XeoW5t0XWr4R+KPkHzEQim5BwPZ2OriEoH2xcSR5UvLFe
YHepWxX92cuI5aVj77sAzpsm87jOsG/8o6Quxx/xgJn85EmuOgg9qCcHcsrLcqRa
Kn8G4Q56oUD88lruULX/xBeXPLtxOSh1zh9jr9NacS7z8su3w8N6ny+HXFBpAyj/
Am8l3cbP5XXiUw0xdEXaAQu/TCE2bmg4IgWLXK0H2onC5FScHNoBa2j2ld1jspFR
ogIDh7Xp03Gv1MiV7gPqVZ94cyE1d0XUsQXxaxiKrvy+9anTHbNKWFrWJh1PuY8Z
4f9NlCOAUMuLwfUCePtRRrvuWBRbTea2fs9Yc65JMcMbYl/iO/3Dw+5OEzj6l8B8
hiKYkr3hTE5fz9UL1FRouzYRhcxAznkwJOij/KbSAC2Md3vh18jTz7vT7AxmFTZF
8AkC83BYWuZZqGATSFw+9NS/sAV2dQmvjQb1N74l5k4icjoCUpnWMPGQgZ34hp/F
TxrBEUXWj7mW3KFtTikyg5Yt6Rg5oxwoXSvZUmPEGhSO56lejsSp6MO9qT/gbAz8
lCaNfe9Wxq5oHyxVA1NDycwZZASfvhCVV8q7UeIbXyoTisPK1Dll7cNg9t7BrmKj
hMj8UXaNDzjzjf8KaTH/t4gD6a3ieMDTeWstOvm+Iwq3pDewZLgubzcBKQ5+ctIP
uwBnFQ2nqLXfsK1ulZLGmRQaHwN2JF7GpHOYGM+ppa91ankGQ5izhWN+M+c14zsB
hHs+6N6+eeLO2jVYdz5s2t7UXB7rPAlfzfhZQyvRCseRdqJNdBVrQlDwZxayT4zW
rhPEDXV5r87DRmkXzViInz8l/xjc+QX77Yj1JdihCowuzTwScmrxtuGqXLiRW3bI
grvt5Wim0HeRoT6iYq6VarXkrjYEVsVdv+dNC3IZodcIN3/49QXTaVSVVoPrgyVl
p31QcW6RAw97ASFrXQxJifFDRXf2EFuXqjyqGPb/KpGq6qZzPjBSwTIxrT0Uerah
N6XXqgmo0sebjC3aApR7/Ymcf5Qhg/svXuvDVnRvfI/1A0Zowml6KfefogS7Empw
eb5b90bu2NeVUEkh80wX6PT/bUW+QCXEKzPo0Ta5L6wGAVOvO8LJp4vgwdRRjjXW
RH+LE5HPs1mSVscIUN7CRrKg6004j0zo1Co9FJEGn1pGDAP6522ZusUw+XC2CRUl
J53rqMAk0IUYXwkmR04jJqvCqWMfy9cjUvpWZeF/yZ2BHSKySUHw5Y3zaPcTNhe/
d9IoOiZq6tbQizLORYPyKURYKBkeZIopaRi+F0sjGWlImsRGb25lKiLeR5Wc+qeK
2DGeqpjNkLFFayycsh36YKBfsYI6sebzySzQJkCoHwxAIhsiVTE3hGYf+PyX49Yi
Wo2VU5HJVNhJozCb157aXQ1Gb0gSKd4WbJplP6yFYUOxISbNLupGSmUSpSFAG45l
4Uj0VNDZzCNPGT/LboY9Mgz/xB8O6zbRk4ABHt+BFVdnGnlm55LceprnhhH0td0z
KR/r34qrGNLzvs+y281pMBPcHRDKQn9Az1UvO5VIGaxCuFaRdDhmHRmvQ0BBHgHH
EBCktXl7STFabXMYfzMSJajyZbGjKCmigQBN5Y+hu99pSEydd9cDZHFHPWmflxdu
aUUL1HrpTtzjeoRHYaB5BqFoRF01T02FeAk2N27OILjupjLiXsUelg1zE8Zv6998
jndwX2tXcNHlnidYf/+89uYTuEAYFlpSGerMyu8ChfLG3cgr/GKMlTgSe4FElOGH
73YMSJfIZs0v13mVxk8I/XOs6lCjVvORO4raEBWfTsZ9E3KKQZVhP6CetLJglxiv
gtpX7lk1Sd8DYn03ORrxjYouURVbXHJ4WNdFhnHd1p8y0Z9/1DI3iluzpYNlOA+d
/548HLdXd/vsZRRuBC9aBV1vwr1MuJYQ3cBm5hIUOYn4QPZN7++QAgt7w1Eok+Ub
u24zfUMQCkat9MzHt46akPA40B0CmqP/WgWitW2OkkWkkL8JRbemKxYXZLUvQMHf
6T/i55UtTJrY7v2ywjg/nxdLzzgxNJge/E+13WG+ngXEyQtkQ6PqSuPzzSU8egIG
fGO5y9AqZCYiaA3C32/v6JhGwQ3Z2b31T4I3hQNh2VBCodhQah5R8LMmxkrBwPcG
YIutfB0pmbm4p4W+xiu1DGCuk7dlVP0nM0bZ0UdpST11YWOTGAfxObIwQxZaO1YI
18tZj6dO8WWEXijd8HVfBE2mw2FPA25FRbhZZsD7mZaxZxpPyyjhqx1gtSwGR1GF
Gr8H36hJD7MbnatBh9x1QDrgN17VHGPvXudwr4js8k4+Nv61G+pIDJeT/bdztqxY
482d0jM8CwUc3ThkY6RpM1kQYQ826iyLNBprPYmdOPWvw99CWfNr/hk/MgcuURBN
AO9w8/5KvV4WdRGIvYphA68hF3kXvmizztsp5TdHFjwvp9I4qNaw3gftlTEqBcc0
EVplOqHMbUDiLFxNh0Fl4KIjWUiCg0nkdZ6y7Rb0RfGKxn5dlLZPwEF9mxH7rvCC
D9H3IrVhggDhf037wMepBR8VAMu4uSSB8DcyYtRXhdQHUp6aVW1gwGuoLrrs3t7y
j4EoQJ8DSJs/BNQPFxkf5SwMpHQnf7cKYr3iY/aC0mpzy55xJnDKzOXchlH2TsTg
SCxbjiVBo1FyWnsnel6+inHFmQ88Y5EMYO/7xJNGeUjwPhzXmXxiorM0Kx5YIggb
VzGZwZRZGsp4Bix84je0FrLWDg1csWznV2iUXfoFYHy1KpslWA9K/MggucxqRdSz
prTFdDLBfY5nczMIpH01hLMGLpdzGCNb2hZ9gC11Xb13K7LQCaFiws4uuwvd3tJk
/6enYp0p45OnPHVnNyi4io/22S9F9eb/ut527w2eUZo5IDGwfRC3DCT7JsObN+Py
9zOKpdY3GiWtyQpJDvPgXkVCE5jpManQq4YATx4cEj0GOlU6JW+jvqV7jop1nNd7
PGrB5zir09NnrFURj31WPsgLVXlm4LzwrGo1JwhUZCntQ3zA5naGav156H9zbd0k
zSjOAPL45t/u0YTNzerOehozSx/gd8sUW+Zn4bU1oj7tAa2KFRByaOz7w8oKKdME
ZGhM2P1Y7/gN8qh+uJIcfrckmpQWGqhQO0Bxd0BLaUBadCFiYcYJaAszVQo3NGp0
pm2fnJ4bS3CeummN6dq1lO67HGPLzT8X0Kyv4Kb59CxW4ZjiB9tqTgJT9vorofrn
D/2yyo4wO8mPn82ch3Ii26cmfVJg6yStdkrY7qREJhZ4QLugstGwDzdx5+4MRi29
uIW9XBfVUCXNss3BdDZxGNChVnaMlGJ0hfIiwa3Av8ET/Ocf80PK5Xe60tN9NLXi
NBMKAoUqs+aTYCzRj5H/Aom9sdOnsZ85DA1QQurN4zAY/72HU/0/lS4baKdxNTbE
vMbnvA7TI1zYaQwr5KXlb04K1kleH6tJGjCDNYZAsbDFzcx8UgtfR0kjIyQcYGjP
JJyISbI4vnnl0Ws1m+vOlBA4kPWtN62uAzLfeRds5vp1C8R2bNn3fAdCOKTomD4t
zq5D+q0SXYuOcPQ9Pg/uce5LOklSLexOCL6DhsnDK8G1R4mt1IIzxDVcPb6q2Ehm
CMVSo/71hNZeYcAMN1PKc38HYJhz5/LkZoKXZ1ciNjf0VZnl8+c6rfTJO5TX3ezS
vR8JT+B2dfQOrudcW9aFcy5ZiT0P4M6dZWTYaSD8egozstk+aU38PlmdNT7tqFud
DujtVd8qyTOxCL01dsBmS5tCzZlA38vIzVupBlwRepGrOAqKVzfSmdQN0gZOwBR8
9wSgaYoXffLa+MW61mG/kArLniJVpSOZ2J9nwHRxAdYWTHKwJ2Tfshl0HSYVTzIS
t2PJs9cDwVGfzpEN/lrJAbSxE7Oi5OMoEyIGnUJKrKm/T48rR4x4SqdFhyrB1gbe
bhQ3sJMKJMztBNzKu9N/c2QDJNemJvKm/YHqcwRkUj0HSSBZuK7zb3Q1voN/n3Md
8oOk2U/xksE2J9ajWiz9lP0XqhdLqexPAUkzNU0h6AMpXxj1rB+vQdKbsKvbmVj5
crB3S9j9WUWC7grrQhu2QJwemnkGP+yYkpA+cwmP731yO+zRmbYsq0OtkRJhRMdt
XV+mT/xKYjCc61stZrqLGNtrGzxNJ8F2rXwi5mz1zO0x7gLDQzZlxWGEOfDjOtD5
i1XIdYGz0JVPPo6xE5OlbFCNdgt9MMGjoZOu+WqWhOACqzJrU+MQRQ9Ry5K7dHHF
c8tJgaJY0NeBNFcfg3/vc2ywwhVhfKdgmDB7AmmowMLiImF1EGB6X8vSaJB6yPK8
gyyO9QfFd69Jt2AYdbF6TVbVSJoaBk5oTFHlOqfjOfMWJsbp5urdZWc2MjC3JxZ8
/IsDnAgJnxmvPNv9i7ZlqMzHsjxok6LfsiDgQdFTa1u5n+F+vsff05d7VJn/ySdZ
MdIy/T8BiT2NX5XC+1EvxzZsnS0iYY+5mJBvgnDPz+vf6xdM6pOri2XBfA0Ab5ta
oOg+NkCr8sBGu8vdp3BPO2dEcKi5COR/6zp2dJ8cmEBrE9VkzTT2VBXA4CkZajAg
c1yMCvqz6WvNhvxqbrLAyqAvKY0ABHBAC18vUXSA265H22KhCOjtU+WWsZE9AYW8
g8GFjP9O3kblScOkkh6vwEwVPoPZJ1CqfTSeuU6JoeHqlQC0wewQkCdN0W5punp/
j3teWsCLNuiLn7Y5KBgu87UZ1hnqc1wcoAaldPC/O6eLo/SZyGUb575b9IDJcqoM
qLL5+ntUDHGhHnJsVYFZU8Yextp6LMEgDlYkzk06WQCsqouM5pLsKYW0GN9K+1QF
01vhDuD0ChpC0KPpQv8UxRNglP4z3IAm0v0L3oaWYMdihCZmfdoC8MxCh9FffRHI
FEvxZZITKZloLJ206vWTcddmgJBPahUOvweRzWdLDO1c/ksCMKrl70f8szVte7DH
nFJ8cy6/Ocx8U3B85zbEQH2Xv3pB6i4Q8NhGAhsmUnys/q3/RCz2IXdIh7AF5do0
ukByNA9SPMZ9Xvf6/BrpKKLNWz6fXHDK6SGIe13VGCkBjaJgG4XvRQsqeCt+nCvl
X6eQMYP5nBQrIz5zaKLc23Dt1QbOw9EUCJXiG1YIaeyFaFHr8ZKbZEA6cYePXaTr
ZP5N3rWTOQajbwvhtJfEI3hax05OFqDabVQeYs0H9U1VqRq8HdEtd03cf/kiNZa5
CIAG6haz62YVU/qaX3IZKzjkYvshlOWCvXujNpEB1QtjLAV4vRIHlhfgqlSn5I3F
35y0+pbQtlcTss54zWOpmH6O9EWnyMHHlTCD51fkFeMRkYLGgv4VO3GT2y0BHj/n
mey4ulOv1DlQw09pqTobKN0OSHSrD/h686CkMaKblC4xnfRDcvWEOQ4yI0yM0C3p
O2vl4RVj9Kjq6zM1z9XSwFjX2LfRunNdsL18lB5G5A+ZILKjOx/nYbpdJlfsijV5
Tj+PpOJruXGtawWad/lKCuRI3h3i4ZAB+JBFjMICyBT7o+X+OBhtAYJqkDYjK4hT
W2JnyX8LpAJQqzahtrR2TMr/51fwO+iJb1m6wEKrl2jbs491Aq0wd2q6lB3iBMEi
JJU9o2GPim08szR9aZj7vhs+igdQUuevY1wlvNspRRTiA0eM1AJT4ipPaIq10Xjg
GVJKelIJZPRIi5KKEFln4d6KQcchNTmv7h9SIcwLJRhyRVk5pkIvCXkRhOavK8uT
oUzqug01J5d+FY/l5hExSyCdiZMfoGgWw7wRXAuzEs3HJCLvaaxrfUcBZIWO426r
qCuu/VrzdYyrloIHVAL4AwHiEhdkElPlkjB4q5unObU1by5CyHCEaCk6KtZM9Fo/
yQ+kuPwJjjfJ+y5PVHM51hwpxME5hZ1pWvD6iO/gwO18CMtTezSH5EEZ1FuvCzKV
d+ZW4hOi0PgBuXmd40Fg8DN2+0/a+2E3Y4ZEVKB+3zj1WCA81NEucRGsUHNWQsfP
0OnVlGUpwJTvEqG2Tjql8jqy9baV2mCeQsnhOeNaFZrbmu/XkItoNNQSURTmsTWU
hXtZZomNEitH/2GpvDPVMte78fdfKpJiboabkSPnMcZcxiL7BDHhD5t3duNarWoH
5ElXHshAJ6zYQyZyVk51eFzfw2ToM/2K+lPh2/oAN4d/3nnG6knE8HiPovXwqOb6
Hm3i/mDR8KHQoX2EyVvUNDrpPAPutus82M0h5k0t/yLF12S8a1VbWFCOzYXW7Z4r
Hzb9D5I/bv/cI7cacY3OXmlBZm0btKL+8fhko19RcRoTJMmvlxqthOCw6xZc7HeT
rmqCPEWkuNydYpq0Nryf8wSmpVfpjPor3OhKA5scLcsbMF46xr3brIkvO4cPSdcK
nxu/qvmxK3KfmTcryC1ga+iFtprC4FpfHE4sYPWeParb9aKPzS+SxC/mkXp1SEtJ
SmB7HyG9Z5aKaRmjHypSvvP6MCpBfQa+inqxHKyF3S4IoY12nY0KNQCwj/uklJdV
u3Hk27hps8p2AfEACZt8PwUgghCBsuR9Vv7tdRWe3qvVqT7UGLPJDH6g061//CaP
2eKtUOlthfXArPzZADbemvkW/iIuo1yMGOSLrOFq5HTMMI4IlAHbRYXAVRIXA8px
lCem4tkI7BvM/xexLIwRum8ghP8Qh/lcd8PlaoZDzhZMsGo84M1Jb8NVIPOjIL/J
o2/Oj0Gdz2LZFtfRICCbkP0EnH/ABnOcgEjba7Gk2D8y9QdIDvgOC4wrjze4r5Y1
PWQLRLr2PLkhzBb6eqZiuRYIKKoYjEHai8G3Pa3V/jZ493GV4+7BFMepxqTByaU3
eNP6miqwkxO2Ld8oxEqK+Me3HpSTAw7CBr0SLpCZih+wVlm8SqXmvPLl9HSiLKxD
ylY7+Evv/1kEtSmqlrv24kFs43VuSVMfenGD/YgUOqMKe3pqx/O038kV731wpR0P
d0jg2v1Toi+j2M9Va1A2rVAj6p96ZvNHMwOrQKMFYIFraI/WJz9mng+BaslZSCHY
vcx/CFRg3bavnFY5xmc1jJKyHyhVRqFFQwEAfTXtfT3I6Vhi7lgsyicBcuFcy3FX
F/sw5iM1NhuFNDvLELaR3Sqx/J6f9W8qn4GZuIgWHq4xpTZ0di0jiWhYCPgz7837
dSK05gnv/k+8GvuLNOTvXVvElx1PNQ+SYg4OVy6Mw1z2MVEgdl1p34di8vGSIGGg
NlVC+QobtQ6YLOafAk14mvnAxl9kNgXuY8vTyuQiyW6Mw5BsAROBf/Xym7LTZzPR
FPtNUFaF1c+tCYG+P4MXnCuDtYJb3mlFPBc/AVmx4JR3GNX5lvbzZv0XPF8znFgR
AOUoVL7TN55w8ymKOVsVyDiWTlcB2ucV45TcFuRNEJFAAAhT+PeGp4RefoklqNiA
ChkfyJP7N4JCZWtezul4A+xJ5qA4Rqll4IYFOJQ5VrVdVEB4YAIpg9Iq3ZnxQ4KZ
lUb1taBImP4thMZYTtgfXZCB/D+9nvsQsRvTJYXEr73xsolJseUCcUvOWJnU8xaQ
4RH39dwJ5qClx1NuiU7oF9NWQXaeDju5PC/qk0YIlxm8nzaB8M+nd2UD0XkrRAE0
lSHx8NOjoO8sLMdCIE5J0m1I5BLAk7ES8azUvjk4L6B/jVEtTkuysIw82GVc2/eX
cjTZSaOhID5FGlCiTpxSKIezILZBXBFcjMrTony6gWz8kVDvWwErTuFJCdMGe9UG
laNlfknCpDevOXOHnnXS5I5dUv4dYM0/H23NtRmbWxcxGfjeHFOAPIl4KoeXZe5K
oCioeYA+eqM7/T1/nnayBKYCRFYi4PzYBFrHYtTUROI8Biw71nfV5tYuqud4vr35
IvlIL3iJAvZNKOWvVeSLBaC8YqcGORVAb42a7X5kEON029mnmrO27D2FuuE+k6bY
z4C+MwnMjJNA2zZJ2ljn/mcVufMB+JXS/SzIgM3y23FgthtGPO0BTXajE0p+cAkh
J/+hIqtlp1AuBOuGvd0pmPkZpohQpZJBvvCJXgcKCc1zJ0wm/4D/C6GM0PnLOqld
jg7GL2rgK5K5/0qzwAR1uFyupklTYPc1MW31GtuJRWF3z6y1mlsCrO97008xcbb8
aAB8RApiK05bz/AXjFv5uR5LZmaapFZTcKCFh7Sc9wfyISrkIg1jbvk6AS7vqhW/
Er8j1NtqIirrTbkpMZ8WUQmaB4NcL+TW6EE8xNnp2g8LNJICkZcfB0JvIdZagQfR
BdXWbA0QZuFRsqhqFaxI1Q5Q1HXSzA/CKm+uCnmCayERhc7WkRXgwJWV3Mcn3c6H
8kKSKQ4+WVi73QXHbQ/8YtDtx2PX5nRuvddYQ2GpSPi+d+NEB4P1yyjzXYGGYwPK
v/j0qpoXZ0KfB07vcYVLytF+StGp9cxiit3AO9rzegIG1QZ0RCZX3JghMoXflgb/
AufeX6cJxGBRSvFnqfA8DLRDMOIwNtfPFz1LS4BOmGpoQGU2z3PQaDkRFq1dVUC9
G+M+NlMzhvA7ivMau0putGNTDsgV72jy23FIhWPhixb5bdNyvBZdYFQ1/kRFsD8d
JUp4ZRO446jIdbJmHwCZVW7vNQInhdlX5PjkWklOznIX8Cv8MAMTHysVBEbDfFBM
izYjtmBDHXbrkDUTRvA40XjLJJLTMlK/nT6oO5lFcZNO7rEz9miHZScU2fmCtj8t
2Pf2HN0gbbjeJyOJtP88wp2oA3gdrXx4ZhWAQoUi6XL2R3jzf55FW+MgDHGi2oLU
wmcaa6AMz13Q7rSaooGQLXBYQ2byufeu2UJa7VBoFLvjgw1WCqfUfJfWIbeFtV7o
0ZUPz74v2UEVCNjEKeBlkbu9Anrsf+vE7SwdLfu+4HQ3YPNc/kZE7fTd7OfU1Bp0
6Yw5czenJWm3nvKJsgzpjSvM1CBHmgKdzsAKgB4XXmIG2pEyiXYTo/LbiBwmS/Vn
KthMquH68VQWcy9P6S7Kkqd8KVLu7WQqcbObQ4b3Nrd1Ed7w7Cp2jrUwPp34A2P7
HZiyAqUVLw9u0Ur/68Mp8TdQNVxpzjPifVck4DHgAnqK2DhZofNdhc4O71gFoU2V
1wG8T2j6EJ1LbLLq+5Xz7DrgFk5yOnaq0+J993xYSsm1m1YbkrMs7efg5+KgHTko
4a2HBwvK+k+uKERASoEuSuCiGlx96f5ywwnhIVligemfoSncfw8S5c+pJaTx4fmK
acCA9QPnS6Y2qDDl0BLl/qD2ZheB35AvDRY4Ww4ad1sDdArNyRB/g4n4AauUUbWw
ANCy4SL2GGb/CzjcbDSPtIKpIuauLPYo56INzXgPdRn/FMSVBYwj9jStZYPaU5PE
PYXInxFBHGG7E4Z0gKhagevFYY2qbY02Kc/hmlq/lqB2fofdUWB/3yJhnOeDSmnx
uoHdjP0M6Tth09XxJarAkqIsukt8hNqk0Y3GywTgA2wHkqGAdy/UMsmN11nWjRyB
eLh9im8mcWsXfZ8KW4/ZKL/gzSe2GdTYoYKLJFXuG6zZUIGQU66WlZhzFbJMqJwW
J2Ndnte8QWpRIyFH1UhAoNgCyFot6Awq344xcdxhe1UL0ykfvx6QnZDpvMQZooum
X/l1ZMelPyX8NctydjdthsgCo94BT9n0VK3fK6qAcA5JslJhAx/hpmPScd/dvJmN
m6Fw3pqhXDGljiaeYIrFGfgiYdATi029V/UCAIjMDFJAq0NVYv9gWs6bxpHAcN00
BcrE4ThGU/5LT9ctvvoJPxAsUKu5B6dG9ao0h2jKhrh9AO+aEHL4GAFZ3dtmH2aJ
a8vS8PpuBKXRNaZh44DG3eQ+r5hNXcXupwbU+cCOX8ZroL8l65dFLN1J2NN3L1vt
6zt8iJG/ahAOD7+HKJBacVG9ZPowYs/3SNfCNDfo9h1DoH8RHqBf26AQvhr70f+i
DzoFZhDphnYK7l+v/v7eKp5Qk6KmBktBxmwYGnx3I/FNOJKZYTZOGD1vmwJuWFE0
7sACbL5MfXkHhlYjIbEAOc6y9fWVKYccxA6OTkbIGMuUL6MHil7SIyu4rHElMvtW
xvxfiSS+1gaKKIsazFeIjjjM94e9ycjwBSllZbqLb4nUDrWP/32egatR/magHhqP
6QsEOydkT2FlcU4yQOVhdGXG7wXdknc5OG3TigGuJ1NoCivTUnw60CLNltmp+k9d
AgKsKu6srj46UiONliREmc3GUhQHh6h4PWzVT+CTYfTwgoZMlpyANSJ+Ldp9Nw+h
oai93YhssfuuJjRQJZdw/hkHzJO/su11giu0ft6YceYKl4llvY1tgfQc71+9LeKk
d3ty9PytMtmzvj5KfnUmW0dOH1jcRRHrfZwSuBa1n2HmBP/8AD8VDuWzB29SMLY6
V1BP2Lpcn7dpY7Lk8bZ8I0SKi2Uq46Rosef2eSlS2NTMdpA5t6zE8P3zWlsmxCzY
/QrIbGLr0Y8jXsDNWYuZCcp67IFv2EYhjEkAyHSMeW/GsYr1nDMQwxMm6tIhJK5i
NHxwLQQXLIeRiWJ6SSLDK3sHr6z4XFHrbOQCsTQmDhTWyAyBKkrCNLlo+0ypMIqQ
J9o3DY/vVsJz3r1ngUbaGYqdYisM3bIsabvH1fmh4G+LsoRY0KvM26mq9gxc4KEV
CmIfJudwGq8oJ5+dER9vQFMXTyzs6C6HKsL3UgeSUV07sxlZfAgoC2ckNCt0J2sg
caW4G1CG6KVtKzfL6lzGtMRtmyagNzGUHjN3BBzvBtgHmzHVGkuEoR8/7DjGhj4o
EIrxSo6z8Qoaj3Yjhs2YHPqO7dErlDpAH1H9xaWZLH+OQ78WItUWb9BJjjPSG6KN
PC2rGlK049Qm9ludLLXGOndp7UgbHbkBPnNLS8ONPrFKoz2CYVbWZP0bYFF+A+JZ
wNXdYjlS7WjoQILXnZHuu0kfDDFB205RvqrQDeHR+byJkOdxy+QXH6y/bYqBTbIu
ewLACAm3k74qAR438ieg5Ptu1Zzk8fJWDb+yw3CL6u23y8DVIvE1KH/+1AZL1z2F
c3+o5p728xAodw5RvTlr3FvycELwnjHnrMjI+iPap6+AQSa9tvh3K78Dhj613A1B
H2+itfiEAN9QRUa0r+i2UhW20dt6ULgE/bHR2MXL3V/GCvGJXFQSBVJvjucZOSpf
EEKylE2/E7eQIS/8uRCXXrUDOi0lMP5FYUoaOtede7pkbx+FmrLuEU0jH7xh0rC5
EaYxUOykVWfUExK22tzDntWxIk4FZYfY1oEJ5XZJ9ci7KO4HIz4/ogmU5L4woAZ0
efveuChm5GsgeqivdPuZjxmHuLPZxgaCfqI4SHyCgw6D2WOpBeg0Gf7PMHtl0eQh
D95anaJOacdD5TcQt9hlYDjajawcSWMRjt5SiPCyMzaWrp5pxnqpLo+lk0M383y5
eR02hTHRy+9MTK6wqHoiCtDpaA17Z1KaFKM0sjmW0g2oOiN6udCjNEpoucxFmeq4
YDBkKfarLFElN8WVDdcx6G+4//s2Q73qHTwqBp3v5Sk10mDfNedBFEwip396xi6J
YFY3FJDef1JVG3wiDceC1IZIGK8VHMxpIOi5t+ZsFrxieLoOOZaQy5TLrZCPGRQN
d2NpdwV33wqY2+zm3QfRybwCoWBWWLkFSl5ydN7IhIZzM3zqmFAhLi6/SGSZfJXy
8pkNRvhekj0fksOPAhOXTGTS+D4KoD0OBmAYIIWtgUBMEATl5IkG1Nk9s3BQGu/X
cZ2jjb4JLJPn4yX5IwRg3KGu+e/ddzOQ6EnNawSiNsDalucY8A41ox3RnIEThKsk
XCA7GY+Em/lNNxSsSfynPTXB/QXGgjGTzgfwUNCDJj8io9Z+oJ3Pb10Tija3ozEa
smbxrQwlhr7PfeUJZAnR+dr6sj6d88RGnOR0ZjOdS4ptXXeen3NCU7PVhDpRSdD0
LecnVZGpZyc0N6Ew4OSBC6hU7/QQ/JNBBkkXxUJ4H6u4Uy1vd/SnfqPx0XzAr2Ed
Oa1T/+nk3H0li09Gd3BQjYNMxuZCKsu6QrEVXEfMqbLN5PUgbdExF2XApKlWKvQw
UgqDCY1It07Y5ZQ9S99LulgPtsamFXxz1b8IYSm5VdK+IgePwfU5V2iu7GBgCVl7
18fh45MxlBqlz2aCMRpvIAgdD1p9iVnxuQTQoMO7nI9RRAym2r7z1fIXhUuGusLQ
qNgyGyuOPuN94WjU1HaZPc0LhCq/3R9LSD/zCLF7GD6mzrL6Z+JlODVxWZZ2999b
nlJQtGO7+6vQV+O6KVBOZcHWCxtSyEObvANGfV2QTAzlkNBsH8CgaTbFd9XRo2RW
4MA7lhXRexF5NwQihKhFwPvyepP2hjUtU7h9ojEUaBCAO48eYbNuCejgtV6tmcq5
RSGtAhzRzaqLsvbkCQvcGrewapkYg+2vBD9n7FV2RGA+0OUSgZ17FNoXzGzqYaqh
yHsz6nZ1HpoqTDcDfwdWgtvHf2vCHG3HwaswQu02T1xfmlOqjCDEK+RDfuldttnU
4bL9lP8ag0ag/QZHVtXbk2hT88PVo6fXkKQJ8pcMvcPfbdN9HkAdQOO6K2vIxlpq
K7vZ+iSYF80tfqZ82h8nufgIbl/Kr1MMJqG2Q5Y+4g3XmrD9iSys//o3pk0Ta2as
lI94cliSbx14Xu4/rS2LpckvThtaqcrgYqSBegBRyOhaWxjMohfIa+gfoYI69l3+
Evu5WxlyClkQfN6ujA//UxCMb97m6tR9Nkb7Pc6SGzfhYlHk2ZeaQqWbuV5CpvY9
y2MkUujSGMdgfuB+acZTrtleloMdEdnWv2oUlVmSWyf2bAFy0XkV5C7q5soB5oNa
n5NSWD6d68uWzLe52C+HeCFpd0RDIEazcHIqtQ4+NOTS6RL4B0Zm649muzTm/qzt
he+uUkzt8cZIeoJ/axaFtqJEwVFlD6X5V41ISMkk3Huecqscv2qSxpsqBTx4Cpmn
lo5dBRWdLkVdNKpSbH0Q/0iDDBxY+8vThuAWV6tZWq4gw2fTKU0dPhaghjAkWbgh
TIPOquLUalndN9bNzxDPP75NxLUAjE2/2K8T+ukasaoAnF8VYj/13Ah9sJNMYVQq
76CW+gmkfYpR8Kdo9lGpXAKl1C5mlWt6MdTBlZKOsonFzlzhe3Mg72mTUfpCH3wI
vOn4qcRs/94efHLQFc5kAv4C+rqAG04Ct/Thz7izioj7rNqT7up4C62J9VluVrAE
3wkV9Di0UI0Mizd2g0RfQcd2Stl7h1eO+PR32dUZg929qAsToSCrW9EF6U+gGd4w
Bge7CsvGsODl7xXUGFrmeFk47ETI7iNv73w/26W5BtOIPopAGg1xwTX53EpPYNWl
yyotnKUpmXx+eMZ4etGSMZjbSc5j8UdslarpyM1HPaHS48iHsbIVErVDFgR0FKSh
cYh5Um2MgsR8SbcTauik6WHkqRpRTNehV4C/9Ih4sZ6Zgxup47n/z1MMeD07qMw7
rbCh+fZ4bNTRYMrtz0tz6aj4zWv/i+4iakx8oelQXm6cMb3UuTmz+n03JuWMfo94
IboMOST6AodaxzxQ0d/znS5pi36sX+3nx3pUAGeQvIzztMIi6Cmo2Osc3fSdQION
+6mtZDY2mBvqM9JTmnPmnbB6DEq5z34CA/HbWw4DgLRVUUgsszWSieGOIE8Hzo0C
teKy7KuDiY0olq0BufRiGaommRXt3lB0du6xr+w66lqgOHZQcA+ko3iYczJpWx0D
btjQGTzARQqGL3pemcIzTAVppvTxFl76fQ3r9ob5rS8fPUTOjfNQfrxwBqwmdWgR
/g16s/PuchJ/woK/hlLfgbrRHmugxYTPWqgYa2fIJZi+64YraUYA84kM+SVpd4d/
Qp75qRvdAxNV8Lz9lDyiXz9DhGMJU/4P6tZV6/nY4hQLpzkRy0EYtpZgsT+sxXn5
jDeRYdwQC3KA7rnr61q/GFGgYDV/HHubnkZPNNq60DNgTp8rhD5rc56SfpvUJU/i
OiFMZSk8Sq+rI0RfmXg0G3ut4NC03ycWkCG+N7snpGTOU/1HLf0zVyDQNoZTaLAF
65jF/FbJuMaUEyyYr+n18SFkn27FqCkayQswAQZx56xchDkSqHWueNb+40G24kIc
iwcnmiDs5jSicERcXHGQ7eBxBV/ADWfuEjJm4xyrxweovpxOptI7zooLobxU5cHC
zjXOzbOq8PBPgyrFLtWAbM8BoLIinXM+uNP8862Ph807WDbGLDF7WRpPsiGtk8fE
46RfBDlayXypR51RwM0CAoXI0h1UZSbhSzcFxsuC8jOp5/EkDqXfA91lz9J+8rF1
FkD9Rlb0giRV/5OWN1uhANQhNcEPdQ9/JbkZMOVLVKsnhRmKezp9jOB5DlHqZQZ0
3Yr2mu8fiUvxbjb3GN5F1MhXR/6xLp3QSxWLUuO8EOifakAP5559AFrzmOwUySC6
Ojgy8Oukq/HxTfrvJWEld4MJ3dPDx1/b6/nLXUYDAZCqpGxBH8Evtka8/vbrDKiS
VIr7oGmGvclCy4zxAGsq6JirHh2qVSbgMWbL8ifDK2n111MBf8EETI/GDAFGg95W
jbGdymIRXRoa9GYYA/MwG3g+KUEOzzLOXDTfYsU+OTUI7jwKNFvXAWhcLSzwzWYl
FV18QjyIVdgqIp/IYuP7dGXuwu5fSnbLLlgjP2X6XeJx+YEmtsDcRGDUzoR3Il7+
RSaAxh3HO5ZO5C+A26NHXRysufJBnG7p+Ey4JrL0XeDJtLwfCsPw/mPel+1phC/D
F5+dSfp4gJ5+KP4qoTmCbjiv1YgbkydiIIK0RTVyaWFw60h5mbvwRSp+2yMAeUeR
+IBaassWh03/T3BkGnmHaTRemtE2/eNM92bIZvI7kvAeINaB0fKjjGCLnGahDuvs
YQqcHbQVfaDPJoYKEqCbLzl4mHMNK3fwCIPzbSLCdehchM4AAw09sV7x/7gEqpar
XmGG/Q2gSTFb8QOrhFBsFjdydCTqEJzdbg2dEEDcDmGXULXvMvU66XBg9phRdu97
5c7LjQsxq5fzaoQNw+Oj4dXLysgGLdB4mSbCmqob+W90/E6jRvKDU8kEw5voD2XE
n3dfxVUTuP8GHxun07JXegK3jCer9BbmhhyFFaZ0M/OOiNO854Jhjmzn4Z1xlWQU
mSDfReI/ezu0zd1zyv/SBDu0uyF3xIIWKvAkeUtKO7XIl6gCbiLb7Tq/wvcS9itZ
uUKUX3cEarPYt79fedMjt8DefPoMVnlJGOIAu+NQ7jhlhVJoIursEzLSVmdj5Jta
DoMcjDqf/4PMBBY82esX6Y7OwLb9FzkZStex78hZxRr8VuyFXINQMs21Ry8s/+XT
Vg5JnZ9P3l0E44zDHY93EGxsKNdMJ4L22ib2/BvENDy0s6mJXu7LzTmFV8VIFNGT
VTdwOhkeSZ3J3RVCyLTUHDGzXu5O86h5crPuX35nGwOZI7CMJVEcbrZ5Ol2oevRL
HyxKl/Eu8Uk09nv7HqtQwbm+zF/QFl4ruvLX2MWRm9FFtypLSTTGRWLTmAJSB7ey
Rg3sVGbbCW2AuLvolsFTKegXzlT3eAFrcDBphKVnqME4o5tY8vxBaVNqjZSbUFyv
zC/B5nC7ntub9qXDTq+lEDQSVAgynimLehRhdsk7o+ufr0x1TaJaDPMlX8f6hhPl
3DOS1/ablX7OnQxQgDtAH68z2PV06jRn5mRjc+UvV23IiSKXmEkFAyF8FhLs2hHt
93msHHajG8vfsxzV21Vzv33DYjCKnRXgTp5LtY1VYojh+L0I8lbi9R6u6GqA+2ql
lVgmPYUtzuiljiqb44NA2RtoDFAd8iTSlX03kLF2j89Ryt8PiMtjuPY0pZh5ZCc+
UuCIYeyzQluWUivVeEGsk4lAqA6iWKQqg3Ygn/xho3IsstS431oWJNFv4X4B/Jqf
CqF2Z3N5V0DvX1ObyM2F6XyGeNcQ0ZF/0pMvXQdybuJh4OV4YiOi1YmLPWbhFBSm
Ik6Xi8+n7cGyHJSmgiXiNUDL0oksi+hBUE6EFvbPyIiYjv7ZBN15akScBDhWchnT
vk5uO491qaILk35sRzgquSZezTjkmvMnTlcXGu6OxKKernRu5NxWbTjIosrpOLLf
q31KtagjrtU+oyQJ0we5c2EfK11QrhcCQXaioW61vK3WDYkiGy8B8Dxxhg8C8tzp
cV0SKK2/s4OkzAuMvKJzkNeKR4uThtTPTATUpC35E55Z9duuGrcmJ0vJjTHT1+j5
FVf0fl0OKe1otXa2IguojpTDxLbSUvol2PulNr3rYWwIZVwi32qo3TtJ6b7DJIsQ
67I1ngRoceu312t9KZjZk99BmdMP1xs47A8pmbD/oMUL/7oLAiEJB0/PuANvQKD6
8ne4B4EEB6BL331wIjPqnKBqGWTZ/rn6l/RhcJvUU7RC5p6W163xtrnj5q04PNXR
/KEvDMjsUdbMuz3b0K+cZGoFh8s+Di81GB0q5nuvJcz7ON1HkHnhg/6GSO1tz90+
h6o3XV5WNdMOBAQjlA6wlq+Ieii2KL5QI6XmKMnzFeqiScKPX1Alb40C/dH+gm34
dnh7oaZkeeO91O3mreGKYcmZ2VLu7ImmvIXID2jzNGvw6+DeJq8Xxp0NMYUloknV
rTITE2/6pAvHaQXo/FZkdaurYBDiINkVCv6YpQceJYgBxiE7hnk7hSzJAXOuhL7i
zh0+V6hgBos31xr9NSwBLyAfoNjWoh8qkU5tNdAka1en+r7GOM51JTL0w6w/UtK7
A5q3QEpTxvwbs39MLFyV4mS3XenMYhczqg1v1ytzmMYEnVPZCIjT139SAehi7ZkN
iJ60ylljvK7hiT6fdzSn3PJLcZFqmWmeNQ2ESAcwHvfjvaRnZ3Mo9UzZDexlD66T
YhWPWpgAWiG0DXwEcqZ+WzhaDEdNaGoKbIiryHx4wLCxccQJnlvnajOgtYQuHT7g
jwwif7Di7F6eCjFCVSFxknYej2Xccv9Jf/Xe/EtaUCugU5ZkSOUSWJkKhTu68GDj
MVzqK5VrZRtlP+E0hfaQTR+qAGIhgIuc7PktI1dIwwohBLyE8RNzcEJ403U5HC0B
5/isHovcRXkbYnBR1uhwXpVGwtqMYqmYhBUfU59AdtdmFNwyuH/vnfhOlqPSckS8
NF1UsuWfbg8GdAlOyvEla3yoTiDDSPiVx6G4v/8a1yBkIgVRvhUaUwvaoe9jjkPe
yslK3RW4exLw4hx9838Y0B4B6c4DUsWu4KZGJuo7C8x9pgghjXMKZlhRwoNu00Bu
WkcCBgXv301jLxZpz4HLgKXlxBHIx90fIN05sJc+KHXDEZEx9XVZuzWNN7UuMyvy
m9R8B3k8n4RRSQdUbYVec7gB4BviDqfHYj1psH20wvfu7RXuC+7t9tRrLGfzYege
TxJ7i7aTbGM6bP4AYiJ2rXP8nIri7ON3L4bBYR3Zdu1vKTRAV1XVHjfXpXRdnCZi
goiT86tZ96/dcYks01V/nLbvbz6m8ztIr4IQP+lOtQrnoFCKdOPJvt1KmuQcY91h
EpFfZME89kafvYa9e0tU0AYtry1w+9kLJmkN88fHm2VIJWStBWM7rc572pIDJu3W
XuUElOPeIf8AR/31Ua69VKZnU0Mvog0kfeouNEhy2K6134iDJtNXCGtKnjhve7lH
T0GMUd+DtrvQn3I/i6BZ70+lzPUldfEpzCn0rSiEX4BxhZz+RfO6rHrwe5+4UCXH
MGQX1WssZKRqjMODQOo+/XwVrgInkjJdft6czOpIvqHmGxg+8aa101aJMeD9f59C
aX+s5HT74dzkpADvwfVCsI2TrMc364xG+DCVrorW8fx2g1afsbVMSG3yoeqY/9wE
M7dEn8tez8hK8UYdKHJ5Bl9/jvCD3HKiHAToYde1FnGxiUWBNgHNxq+agxahUgSP
xHXev7OvxBYxDDDQf5/qz5oIa8pmlScOHV9+z3pyitPVBRvh1Q0Rx1COS5U5+g5z
zBwMfHfvGCDuHR98QZ6a+IqW8sS7p4WN/G9W1j3CC3W/GdvRL7oWb2zNBrY/t+M5
TAXbR7pc7PXoz/PiPs0M15ZrPrfX+qZhZWbs+NrFNDR1so1efESzGYFmDyCNKIxG
0wkkns1aANRdeTlr/DDIK7uCK2/6e3QVDjmTjcwn+nxy7KkH/dRnMSMGVVo5hiet
ySk+byYAcHlr1hsfYOIfMYFJqIRX2LBqXKpkt/A0iI5SqJgp+iht+RrII8t23pc6
hrkjVdBHUFwTcpx//m3t6wKAzqVU2SO3GQDj/vZ749mrRncyaOfDnlcAY8B6ZWxu
fGvuE/xz93Djuavhh22orV91SjdQPpCmWuOolHT/Yols7xGdn06xD7L4Leo34E2f
lNls6JKKfSz66hC1KwYSGXgKNp+5qbh0nn3o/4TDmZmgMBEtmk6RvLNgwusrDCkx
kj8d0gr/9L47CxBLElROKoiQLYrpwcVIz7qKQKpOwJCCrpQbufgAvyjHYFlpIRVA
YkxEGj7TQEctJcoZGsi6MWsDqVVqLOMJxE9+xYIbYiBhHXIbddLPLf+WNGB/kqW9
LXGz/DYU6flrehAP3tuVPgh8QqimlVdrsP6sBUYrNzcR3JxgHM1PC11PVXSqwNbo
nVe/1oCjlkRZS6B/MEqSaxJsKu9epnxUNxc4nQXjJrwVehJrVe/FLTdhgGvQPxyV
orVH8ManpljsPcFzEfpWutua2VHh/8kY616eBl15WaDkiGM4XBsXsKLbKVTwoDsS
UTG1pbQCjfMfTwXGTSwhvOdNC98un/hlQTAE8jB6WMAxm30G9CcZHBuoJzDpNUsj
8D4byIoSliMXg+E5tcrgLRUK03Z5vFpiImO5r5tXnIBzL2K6Tc1XcDJ+xJ5hbK3P
bnj9cMXz2F72rc+3oBheolNfCBVzb9olLaXPo0dm1G8LsjeyNZneTW8++4nlLnz7
3hTkesM28ZLARcO5g27skHUMtJe8taA/Q1ZfKX6HQcXGdX3RFsgQ+LLlOimuAhl1
z6AU9luEnK1RgFkwlpp0+jpOYCvXkI6I19h551H8vk3kXk5tU+OkMOgkTPKEkLIA
xYJDqN4uX/8tlmbL1XzW+Uc8CsqYlbUVGaj60pyU8BZZD0S5/Nvf718Cj+WY3r6y
p9YkO9OxJf5E0kMqBGKFGBkrWMuP2RCd1rs9Ynp3hajkHDt1zdS4zev6/emWcn0L
VUYo8yOwbEgKV+JHgANaqO6bY91C1sWHknJdqGlQIuvPp1h1BwxZRVmZCmyll1pp
RHEQwjeKayRIeF/oLm2aQiWTIW2xtdxpopxLgJFLiTsQyVN2wMgQxj6erxoOdjMc
ok+PHmNpczhyJAQSge3TSuKHm4RBUyTHmyA9XbRHhYnA/ioQIKOP0BIqW39Q3bWe
JKim2Nb+FvJCbbCd5voaOwYx5XDCkT2rfApwGRjcsa/Dsaw76c7u0KPwhQx7v0Ra
8j1C75Wu0T3MxeY1tzqPHBY6vR/7A86bPedTP+Va+cuOpjge/dTc9ZxJ2V39QZvR
whoMtTee5NJkKkxzFWEmPf8X1OcHuDAJ68Bzx5uk24QZCnkZzkGUfQ+2LhQ73mfL
yeX6fGGozJcGkbyD7jIo7QlJo4Jobajnr2ExDBuPGXnAWSTXSueNxpVz6Sw8+b7W
8d64UHol+OBdpYCBcv6F0esbykixsgqO03zFdxVvFColThGz7ZAhRmCtGELA6pgP
y3n+E+wV4rh6gprUTFzr3obK1zDFxoZhE4HDjPWkVIBs/pfp3qASkjuu0lMidf1u
BjKLQVAepAy7fSu95CVG3gSzNw21Vw67MFDtk7FPxzqYFLiEf1dae+mEX4C7MGdw
IR+yZe6hgxFHdkAtkaI2eRT8ByR83rICcbTI8UnQq6o+jdhGRXT2lZ62NP5fCsgM
Yo8DQmId1czB61KYL6yjEiYb/XzhlFBEd1TnNwaxTQOZkq2MFbhw6teTIl+cQrvG
/wO/DK86Ve3IjW+pbLxuRmZJrjJW17L+jxdppU7ym1U3jvjSONI8hvfE6ymGbPY3
pUQ1aDZqbghwhEDZ23S0XRaiNcQg52bNnOQPr7AJT3yHRRE3ElcEJSTF9HK42v9X
th8AdVg1694eDNW4zNZ3qaAbBdD3bccgZlCq6uL1CSBFyyvdSY3MZTfWFWWcei/1
7fA1A/pQG0sqcnp6meii43W3cNC+zLqg/doAyeVeYjEHK2DrhUr10WQsOcrlb1Jk
xu1u70zi6i8tKKt5paljKp52u46FvlVxOSS2NT44UQxQTjgMzb/ZhwYisuZuNaPF
A2pcRTslsTTvP4x0of07omFzPjHa0xWvwAZwi7kLeTYX3HOqR2aHBGST4JVplolX
tqz5zMITLQK+OLw4ROv04l5nOZIfom/5aai4vwEI344T5nhEQWJy2ZcmxKM1XGTe
MlyGp8IuzqNNdOhEg7ejoyyW7WTmqr/Of8GOoBZ3PuGjeicL+94SSkpCtc4Go5D1
OKriYCc9QmSgFv0IKmesselD+KrcVGbiOI6fn9LE+aiHi0hakGZMPq3aJqxVTsBC
HmrI5CscNdue31OAhUDvVcHSbdJv7qGKOrIyao9u9Vaj/SA6DFEal1OXBBp9cFCf
q5rYewk9pRRWikBghdB2B1UY4KPQi9rkwcc++AZZhJgF0Gw2e6R+XpIVCJzm8vwe
4FkIKabwf4Oobxsbux3055GtKeoCAmhZav7gkrcwbBU9ue2h+OFpSfDP9dtAoqgn
R40mabveZ+b366D7xPRnfPaf66gGke9uDocYfNjOaIkZ9bGqwjK6bPkDgvbOcDL9
/5v4lw0qvgc+B72C8jHBpQPJIFlCYb6YSm61yizR5GDYc54arPS/o9Sn2+l0WiON
ZmFz7MngegVR1liT6pFZ8et+HCdDG9GmtbYLhUkhJvLyPutmgq73jAOMEyi97U7F
jrNL1nBAj3zqUHa6wPMIiOE1Tpbeiv34Xn7RrQkrwbPj6WFIBhZWcgQUWQWQAEd5
AGTdzgLiweye8FSUgTFRA5UPOlfWkYzsJUYgo5LTfmeNgthhQ2dFOK0K5mhKjWBq
+NcnBGgQmhj/RW6EbM7NUWGI4/O24x2bLase9rel1pgXMu7N5lCy7FAZkYNQ/DZS
qPsXJRZxcW376ykFLcheJH8wsAl0MB5BzU+rK59OnCuUn/9X9+n5N83JhuUJeltE
zv8M8Ma1BOc4zdq6I5Hql2N8AnJi5iVU3USGRQYSBFnYsk7Bd2rcudNemGSZDcaw
07yfCXRV3UE3vGqLEMvwuKr9/oBlOrC3THGme1wCa7xpZu/kG57IlXMJDHhTRt75
SkF3YOtaKG36VXi7mMaUERE4JMn0QQM1CUO7phfn0nTX6ZNuLyne0H6QJZjt56gG
rHmB1gZYpHS+GszkWqo6QgRX3dSbkgykYqx8w2y0Xft9D9uywu7KBgQoDbYnz2gF
WD9RDtUwMnhvKigDfJiNKWL94Y7WHRVVJ9SLeNHgpzTfoknLO5gh0a/fUDHCvz3r
lJYm10or8DSEuSOkQccev7rPZbgQQEjiiI5TSWorV7ebhDb5JgLsCeB7UqgCsKXN
cFK1ElWCgmWMw/bFXNno5djAOujydam/b0ljksko+wWHf1y+oX2Mrnc7noTUZDKI
AEZ1MoZQTP3WN0MDbExEyIEzO9lWolX0izGaLwXezToVldDUd1wNxgWKaHAzm1pt
eOM2KXBLTFBozZLemLtEeNtX6LDclIhMTvPMYjBoGQ4gFijxMzJ6OY61uwr9sxNV
Eu/bFB4Z9acP3dph/Hnx4cuNkSUOkAw8yMrHhw+pRCtkQr2IDQB+SLsnYa5KTqDW
4uxna/NJtPsE3G3Y+mtcY7Nch5PKVI9so0A58Kmc3hj5pF9jELGpXiMlLorPRUsl
z4GmquTseKIASgx5uNarZ7b3PTFfZ/oq5Q3AS5TbYQuy3W5cSrUyH7my47jNh48Y
3Fkw+gZyTXYz4JYbYwsbtccXNgLVuJwccFq6I6rFULv2Ll1TD2ZcJz6toERi0r1o
n570yZITwabw3EJm/FcYwSQkcKvExTsUJI4Vue5A7aIdLZp79GqbUWPqagkdjw51
8yqk+jyibdEjS9cfsuGQaDwHA2w9uxdYNKBBIVVojYa9YgjTlpcPykkr0Yujzmey
Ta7J19nl/Wh6nifUZOUane9eskV/KyVtFD73LdmnNfKlavoPKdgcBSV4ASQfKG+e
I7SVjJAEQO5u0rewJJ/isqza459aH6WW8vDLLxD8y3sXzG1oHdCU7yRk8lNLHh3N
b4gABfm5VPOCCnSMUrX540sZIs8p9txRkuiNnCubHf61oUO7WzPdUiq0KfDlkqwg
jlqG8Zz7mOJsw+u+ZxmDqqNE12JSZWBSSNJhevY78n0KegYq34dUreeR2RNcykSv
HTAXDCZ7FjqjrNVnaaE/oaqLOuMKxqoJWwwod4XhFPk7tL7PCrpHgILSHDnD4OBG
WJOeKHtrDAYvjHSn/lo1wMvrbrvPsi/tBOlOMLEvKlhImC6bzZcRE2SCQa5YTIA4
dYWl+pXHQI5h5WxV3NV0qZ2cRcHLBhLOBFInRekubX0=
`pragma protect end_protected
