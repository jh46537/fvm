��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG��%�}~���~�<cZN�X���Ĳ��Y��$_V�(MT��Ĩܠ2��l�9-S������d�����\������ U�̉���E���A�{n�g��r��*�q�@���_�q��X�5��YP k�١�u��|I�Zi&+��c���tʱ�e�R��On���u�pu?RM��2�Xd�P��1\k�R]�8h���~��!7�����U����b��n�z�>[��DIK��WN2�yz� _�0�\�x$���uw~Ozʰ(���ռc s_��һ �n[�\��z
��QC�)��B(����SJ�f�Dv�&�����y��W�}�0�,Tݗ���'U�jcҬ��Ǥע4�n��|sK!��m�`�-��������^%�]h6����e�.�E��~:�z׿o�_[�c5�6Q�M*�J���(���n���L~|E����MZa�m/b4�!y� ����E�_1�����N��@S��y�����J+ �<��
m�=�ϳ%|���m3�<�v��5nT���
A�<5^|z��V��\��I��A�@�akjd��9��%�g��k��Z��g�e^��@�>��!. ����գ�2�F<����"08���A����GQ�x��Ԅ&m���{y��sɶ¾
;�Ӆ�78Ì����	����YF�g��q�����X�?[N�V�u�?�5�Zn�����U��z�N�2O~�x�
�����Y'n@ Pl|�t��Z�\?�ڦ�)���M�Õ��7�O�=ݾ��x0L��7pـē�����ej>z�S��O(%)$�5�5�vUg������Y¿Q杻f������S�A��4t	-F xdϺvި�0�ܮ[�)&���.��	Z4�"]􂈣0r��)�܇��C�Bz=*��O���Ņ�J�b��oP��3��>W�p7h�y)}�/0U�L}l(�єEC5�w�Ζd�R#A��i�Y8�<7��*� ���h��J�
�9�s߄���ݟL�1h�r��pyx����)�7e\�v�B�;�"�(3�ӛS���j	s���FH0����6���#o�l�ys��y�*MP��ܨ
ۺ���X�bF}���.c|`���2�ў�{X,�;u��sp��lrhcf��mdl!sV�츦j�Q�BH{ֽ%F����m�{mjO�.1�)F$�!��`3|J�-Um�"=�\�,��[�ZAF2O�pLȤ�s]��X�K���N�:�m��ۈ9��W��s�lSÚ^����CI����L35�cdP|3�����[��ʃ��{���dE$��;W�
.õr.�1q/.�� ���s�-Ī�S_,��G`�qa��A-0�xQ��d�٧��F�B���%���ʹ�u���d,3� '&��\�U����������,��FH���D �A4.��2~�U����<o1��X2y�Y�u���7��'NOg��8=t�Dt���I#I����x�U�N�z���R�l6��(���?#��?�,���|؂��q��5��8*�:-�oIUB<38	���|W�5�>���G�� қ�׵��wY�����h���-_� ZɇJ����Wȿ�|�F�pT��z���������t�M�LRH��%W�];S�2�h�VmcU7��m���>9�c{a�)"�+��Z����JV���t }!�tG>�ϢwY���p\)Cj0�d��tN��[���@��g���U���9Řj���^�%��y��0Q���,[ �@7@͈>�j7����p��#c���S�c������
�.7��.��:bu�׼;筃�Ļ��z�T�s�.�fCٻ�b'j&�����A�=�c��@j2˸����V�tIɄ&�(��)1��Q�]7��^t 9���ʁ���6�I��
?�'?�#y>��P�����vk���g5����	p��`�~��9pz(ҷ��Vt�d�ǽ�I��Wa�ui.�*�~�#��"�'+*���c܊�vu ��ت/�K���@�* b�53Ȕ�O�u�Xw
� �mZQ�mR���;��b����O�/3�9������-�AYP�&a�[}Ab�#��bz~����� ?}�h�`�
����	q�`��Pk�x�s=X��f*Y�2�M&�q	�]i&j[�Z]:?��# ie5���&a���{ǭ���3T]����T��Y�Ӊ\��\j�j��oq�	Qơ'm n�v`ԟM�FF�_WO\F�J�{p���5�]�L��m���-sa�y�_�UQ����:��`7�Ì�h�k��% C(��W!1{9�O����Q/���:Ο����%yp��웇���0����?b7��a��狥H�3'���{4(�o��N�L+�2���Ji�G1[F�6���I��� @��]7 "�,<�_���Q`�����-���_���e����ױnQ8�A,omAzU.��5J��I,TX����UެcZ�3v�9�Pc������-���ՉX���sM�������л!ikd�r�C��9_�ْ	�dp+����V[�nu���Q'��^��M�C�m�[?0|���T&��L����� `%��@��)����׶k��w���j�ɶN!�J[c��)m�nUC�!ĮU�,!UV�휶1��-^��rk#���_��No[W�3e!
]πc=a 9?��Kc�,i#<��sQ|�)SGu�?��%��������d�����1����l�>C������hsV����z����	����\�9�����-�L�օ��"3s�����׺��\��֥��.����7�v�\�gi��M� �Xa��,!���༇��xk"H��DP�b�S�.���;�8?ǥ������
ld�Q恕w���C~���*��ur|`�"�0x�&�dV�|�ӎ���2%NPh){�.~�;-�]����a�s��lƊ݋ճ��.�wߝ�E[��2�`c��Q!�RezHl�����%O&$vN����2J,�~�)4e)�h���ct�f��r3{�>��z�1f8*_���^
�p6���?����F����[�.�{��Қ��.ꨓđ��3���TejN�� cb&�/������Q�p%�l-�!fl�6���W.#���Ũ�!w:�v� �I5"��=�Հ�)��Kq7_=�,&���9k�r�m�E$j�: ��w����v������D�_s�G����:�31_����8���M5.���.��v�����j���nC�aBSŝ�^U���b����7xĒ�b�>CT\,���Q��NE*D�/�+G�c�g�@�U���gt�7��Eh��P7��NeTW��g�7�?E[AO���8�`��}*�#܄������f�W�}bmyW�ٴV@@fT`�_A�mU1�����'J�����%~h]aj��>��Ω����<u��t�0ށ�䧍�����"�x(Ź��ZX������sFm5D1}b(���_9ĽT����eLf�y6li���ޱ����q-�@O=w�*��/[��wm��c|3	��w���!@,m�EH2F%I-%�%�-�V�?GLJ�**��B��њ7v�ѓg<ܕ�ð���fQ�������+^�=�3��Mw't$����n��f��mIdo	z����}a��L0t��*�;)�O�]�9�@�IV���QA5}_����M��s�K��٥>e�`�c�'�p#*�<����������7%�+u7}{��'g�T�7cޣ"��9J�s�}��{��ۚ?=Ez�@��|��0�9Jp��7{ɡ˨	�]֫���o�N�7�[T7藰��v�_�U��!KMtUȉ���-~NK�IIP)��0�g`S �������3��Y:ϐ���"}���﹯<f�	Llj
�'eˑ'	�2�X�����,��x�Z<��A�I1���N� �Ⱥ����!#���,:b��3%RI �dK/<�{'1��P�'c�oR��$8�nTJc�H�p��v�����GWv`ܘ�u�im6�y�@����%*��^f�V���O.h�heFq���	fv7� �\�ڼo�ʹ�I.��-���}C��F���)�`�ۗy��� ��z0L\�R��_w�U�\<3⛂�y��y��ŧ�"Ӄ�1º1⨬LF�����^|eP	-��Ƹ��sU����cߠf��g
�M��I�7��	���iica�MjqhZ�&��&��<����}J}�9 �ek��1J�:cZ���
�����'ykއ�TM4r���؆?��_��Г��Ѣ=���p�{���[���E%e`�g���~'o����L)�i1%#����ϧ�ɲ5�����%�JS�����6C.n���i�Tw9�-�Xh��p�����q�^7w1ak"N�^�#-ޝ���TYϽThm�aO�TА���DU�=���i��w���i�׏a��=e�tp�^�iMw~���"5����/Ä)#����o L\�LqɫCK�m9�t
D���P]gv������{��l��}��rq����鱙�Pu���8�Z��x���'��z�rrR�㶶��&�+EX��É,�P���6�l "��,���E�r�Q���>�(��:�%+�[����9������-Mk�=��3V\8z;x3j�HaB����(�m�u������롃�?K�X���h\~���DIE������+}�Mz3q�G�H���Qbcg*��\`��
-R3R�������u{h9�fE�1|�j	�Ǯt,���r�Y��M��������&�"q�ħ�n	"��q�ru�%���+ǧQ�sg��.%f�}O�s.�uS�.2���=#(4kR�C1 +η�(�R�*?����F�z,����9�V��X�: �!��}]�Xy=p�~^�2Z��wM�x'�����.f���E�e ��Z�D7 ^�m��ĉ��z:6�
�_��娒�J3�T7A��>J�e�h�b�P���=�kh�L��(s\� O=����sb�l\.�w�ed�������Is�i>�Ŋ�S����&zo�C��su�D�?���(!e'���3���:f\�����Y��5�T�ُ��(�����ϋK�#� єC��N,���ɴ-*