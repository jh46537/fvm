��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C���P~�û��2�pn*cZ��.��
Ґ�L�	�2���f���&3H�Mj q���S"��g�)�?׎��=2r���n�2�����Fhx	gt:�T�12s�gx)#o����BnfRB��׵edA��������`+���2�&��D�k�o��j|
�eƧ�9��5�KԖ#�|�{�ލP�1��<��Š���K�vH�ɹA|m�$O n��p����.�nm|Mz���t{A��tO�(O����=�l���M�4�����YZ�r�T�H_�w�R_@K �Oi�y��W't��D-�kI_���pig�]��;c��5�<te�f�G7�75To�2^��2�I��<#�
��^�ne�v�i�ڤ�"?`�Z+�P��+;��1��qZy-e@β�u�_V�����%�J��pP��W�.�����IAN�E��Z�j<{�AVA�3���W�b�LD2��U�bKjv?�Лw�!/�n=���c��1�����%pX��X^�l={���7nдսj���.�l�gdg�����"6"�����!�� �QE����P�%RJ��y��
�.�2yt��!Fc�	����W�:�����"u�өn����A@�^̡ڪ�@�e���U$rc�����R�������H,`�E^b@^��y3Ts��˛�z�jF�i�|l/�f���Fv��]#}�?�]T�OL��?5&Ry��ZJwՐ�_K�ž^�D�#b��I�#���%pR�;}Bs.''.O]�MStjxى}:w�ջl������|Ǔ�#)?e����x���@W㭄'%��z��
��>E�A����EO)Z<��ܒ��;)?�V��|1kD6��-�ĵ�p��}|�U^$�;]���)�읪� �FTܑʟR���a!ZP)1>�$JZf���o���+1�^�L~�Qj���
Y�tެpA��j�J3��ɪ�۾�+�k��G�`�	ϥ���+�v�s���^��#^��P*b��?曬B�^��-�pV6V�p�EM�Q����x���u�qCu�� (��dM����9�Jb"��Mak>�m�!j%�'ỳ�f��5�x�v�M|�xze����`+��ڝe�u���X��[̈́���?[7x,�M�����*�r)�<��ϲ_�$��Dχay'0�2�"��}���T��2����2�)�`T]i�>���j<�%T�)ZR	h�\� (h���y���XT�h�؇�(6���͜钑BFOs0�<������i��A��r����t%�Ì�'E��m�.��:�nm�]�q-I�0Ŋ��WNۂ��SM�`�@���K���(�i|��z� �Ǚc����!jb}HR�,�]���\�� ��=G�7+�v��9(F^_�t�e;(�}�M�l�"�;�8��lU �C\'Ft�spSƹ�Pv�e����.�@��'��Yo�0�ڑ��S����X���/d!��G2�E�b�'p�o�Y'�2+�3�<��Z�n#b��+JU��l��N�|&��ߔE����-."e=F�jM�˛j]�����7u��8�?�,
�M�U���um�O�3�g,�Z���@C�d�����u۔G�=&�#���9�Rv*ih|�[��?J��	��n	�&˒v{���m�f���i�T(��R