��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C���P~�û��2�pn*�Dؐ���U�t�������ގ6�aGWi;Tr�1�>Ч5Z���yo"En�uE�z��m��,��T N�sS�V��.ۭ�����i���͛��~w6��Jʑ������Y���ȚV��(�-}j�HߪZ�~MT_ۢS)�9k�9mOV!%�K ��8�;_@R���&��P�u�@��n3�<��8�G?�A�.�∝_�3U�):�~�*V�,?�!� �7Eዛ�#АF�'��}��DƄ���^�����{1~M�{�Ӑ�B�{�%	.����~�4�U���A��oDI}�dΟ+�M �QvP��(��G��L���Q3f�/!l ������R��4]�/�,]�/T|q�kg��1�2S��0="+��Ʊ���Oq��g����2�N�h=B(ᦥ��|5���̏��E>���hэ��|�0�M��͡P'K��Eu@�P� �>�2	lP�I���u'�������yp!�3�Qw��N|��i(��@ل�g��+a����-6[��*����RR�<j�[�������?I�I)��X�w�k#)K��W;&#�}B�y�}f�|�c��:�g�O9Qa�Fzl�ɦ�@�?���׎�D5<,�qiD6�	N�-�4c�v�[���=��f5�L���}rTU?���]�T�6sԦt�Q˖Hb�i�xi1����9��9?��3V����������+���g|r�mR����o�K��}s���L���r�9^P��v�G����j�����]1>B�tӪ��/p,Z��7�|r��4��$�Vwi/�EA�\s�6�����9@��^Q��k�Z�-
)�:�[���_z�0���UZj ���`�O/^j�2��W_�D[�-��;��ߏ�1n5{�,I���e{V�I"��)J׏ؘ*�7�Q6?�p
���4>�n--�4ݫk.v^��]��z��ALw~mC�� SC�3­�Zם��C\{��5�C
��8M����dA��V'4�P	^����3/��rB捍���D����(x�@p��]B�W����*Me
1��N�af�Ш�3:�E�`Y~[����'8�%:�Iݣ"�	��r�K�{��P���%_�*�U��+Z{$�|<Q3����'}ܪpDn�h*�Z�~�.�?hcG�N��Z��,�3 �Nu�])���S�L	+n�xD��e�6��*^[�zjiL�b�葓gJ�1m㚶ܷ�y}8
ɠ��s���C� ����
}�Me����j��}5H��x�e��<� ���i�ϗ�oVM�.�.�n������w�ސ�����L��4bY��ҿ��Oۖ�� ��V�m�Z!���{�r���iݐ��
xȽf�H<��3���x�i_X�b�P�W}��@b�S�Ԧ��SyZӤ��}���3����ű�m�P ی@n�eK�Y���`$*~�����i����$%T�=���Ċݸd��'�@��O2�O.���a��9�����]I�-hG��o�e�x�5%r��- �T��j���Ŵ����Ý(ҁU4QJ�E�X�WFp �F���t�{�����~��}��3m²�AC��K4�Y$�>@tpLwi��2!�#�	j	Q@��NyNxj�'���&}�y�y5�SҌ=��2o��2**�rC�7�gєv���]�2�ϧ{@PuE�{m|����u=�&��c�ګ8�V�(w:w��%Y�ͦ/%[QZrƴ���k8�ˉr����;�`$=ܨg�D��V��@����{}�~������(�"D�+�N�=��q�Vŋ��,::-���8dB	#�-�O7u�����{8¤#�S3�7�^Ubf��"�b��lLvf�ɐ8~DWm#�t����v_��T)Y�)v2���5U��V�
K����j�1(���[8�,7Y���uӣp�;� zm8�HjC5��Lx��ƿ����}�i�W,��!ͧe��w��6K��?&&�[����8�^*�L�j�
��C��h�8�+q�w�F�@��oK��J�x���b�0
��S�H�!��X� ��:U\+��m���*%��=���u��d��q����Lm"T~TC ���Ʊ�c����*�r���?g�U[�2��N����F�rV6o5FS�?Wr�v7������v4�˲|��A��_�?91/��d�������G����Z���B���!)�d�b�D�����j�C��þ
)lO:�d%�I�2�P�sѷHؿ���9�e��a: C�,��.�vWl�l��B�Ь��3��PV+e� �dĳ1u���.��N����eu! ʄ��4N��7W@��z�C����(�v9c��K�T�YZ��<,]gع���`�f��c0�v��)�	���tW�AIm�Ȭ�r��6\,%��������h.%
�,a�3\��w�Ke( ��0���y1� I�*��~Y��q�z���/wak��ܠ�����2[^��'��a\�@C!��T0ceB( 6'{���y� �TK˭˜+*�Y�)\������#�dT�R��7t�h�:�D�*�z_gJ���e���G�Z�E�ю��b���@�ɕ�g��j�#�G׷E�y����;Q��G�Ȉ���6�_[@BiH9�kT|&O�C�+>TF�i���^�ԕ�c�R��8��Hlj��1�JE�gC-p�&.Xe�H�K|`�WcK�	�>�0�CL����Ҍ��#΃o<K�wDPk�؊�M8�(E=�r�-L��p�*WR9�9oX^)
>������#��o窞*ء� o����qo���K>���6��O�h�~1�	ʁ@�_�s���w�/���J�D(��RN�kXl�V��Jl@/���Ad�8G������Ǳӯ��������W�Z����rC��к�[�KG���>F+$5}cvh}�/�v�ċ�ȗ�~:B�O���s
6�d߆�B��h=��1 hʌB��{[( 	�ȿf����@��uh�����l^k�归O�� �(��`�M��QNn�,װ�Pt�	�x�U�0����wA�d4�g?�(ָͅG�?�m�	-L����rg���qK�ݙ�I�`I�W?�{�pa�Ռt�JopՒ,�����m�Z����)��rv��4��[�W�_�4t�W�M��'�g��Q���iжo�%��� ���)��{p
ui�b�?���J�-�$��Φ�%��Ɏ��DBJĺ�V��;qk��4$9�) ��z�����?f��BC�
�e�X�F�ZǸ�I¾ҎW�"��ﱨ��&
�f��E�|m�0E��H2�>?�D�ٚ�j���nop�½��)�߽��K��=�2ե��d����_v	��DT~A�m����%`�'�ܮ����|-R��f�I�`9�y(�rA"����:Z&K�(2���s�D�(�!$Z`,�=}WSfPZ�4�̫��/ިe�y�4��ْ�*_�6�iz��H�/��b1T����R8݉FX"l8c��g�>| gbӱ~�3��NM��q�g4��>���cw�:f�(h��I�ײPYb�+��GUr��[nwo�u�M��+?�A�Lw<N��d2L��v
Z�M��e��\�g�,ޡWO�~&ngu��K�&���ᷓ-�5�w�F/���Q������	�C͒t.q.�Pu=K,m���8����_T���-��w�6[C#�F�+��oڬ����i�ښW@�{�c�E�W��//z�$�d��?�)�ů��(�>���ťN���0&Z�9	����l�q��>w�J�4e��
sBӆ)[X�x�qvv���U�ҽ$BM����1DĘ���8�1��w�����@,����� kS�rw� :}'�	!���Ė��*��K���[>�]�����t�Xޝ(������G��j>�ij��B#��c�VA���gh��ab�J6aj��\�X��5n�F��#��C�x�+����y8V��E��1����:u&��p|Z��݊O�3=8#z�l+�\f��܈�}u��ߗ�aH�9��ɸb�M
����_1x�1炏ÞV�_%`�u�٬)�A���#�GVOÝ7~Y�X��W�Byq��΅�X_�l,'$v�# }���W�["6�L3X�U�_ ��x�����0� ��7���y�x`e�Pr�!߰��E�+m@N*`p`<��23ا�auK�N*��B�T����np�N�+��C5k#]��k+hA�{�|���ļ��F�����#x��e@Qo���E�ߢ��D����3K��N����,v��ó�I�!����}Ɉ܂E�z45�o�j<
��4QQ`\��67���̶G�6���JL�}sK�%ʪ�̥HYc��8M�,ѽ���
��F���ܟ�xp�0��H��ߗac�(��F��5/��o�%g��T���phJ�pӻ��6p�V���W'�%��.bɨp�P���4�K�*ќ�
PXw�@���b��b��.M���s��_�b\�`��.�*T��Sj{�&Q̙!-a��ū�Q�p��T��@}���<�tF9��TQ��C��4��.���2�,R^���A�Z�?Ƃ�E�����B��B����ܭL�Q#��+��M�p��Dv4�e>�T7^\:��X��H��훌�ᶿ�b�/%�����ь	�y=I1@���av㻒�"ͤ�Z��o�KT���t���hK���Lk���o˹�r�
|�s�˅�E���N�FD�ԩt#��6f?����J*��bh�[�h�Z��� ���AحY]���}.G�69RE��&Ϫ�J��Ġ�j�iǴ����u�!��{�-���k3p��-.�kE��g7����_71!T�$7�ɷ�h�I��p[&�3��i��~�f�*cK�O��v#��o�$��ŅS#��L���9/��*(1�_)����}`�_��1��@��ݜb��J_������T����ܷ����uK�WA�수	�]�b����tO��t��)ea��t�� Jd��˕�o-(��Z��Whk/eCG�2|�.���ߗp�j�WZ��˹�{0k|��^5j��B\�gq�^�Lm�㔻ԗox�>�������t����]��K��ϲ]��m�.�_Y���4��9�gx'D�f��pl1�-P�o���=�r�oa|�,������̊�	)�m]Q���T%�x4���iPz�~[�_?�/r'� \�r�0t�D��]���X���*�?c$�uH�m�ζ_�r4O�&�Q��~�Yb�աyH*!{�+��Q��,�)��r3�(sM��a���X�J�_�;�$����,�-k����Dw�0N�wQE�5��s�Uh(��mBӁ�����Y���[�5Tv0{S����BC��k@N�$`����G�u�~���N��D�c��bwdVh���I]Z��nbMޥ�@5w��қ���(�V}��l�"9	`,IyM"�,�4rI_׳�W��x���9E����P5�]��˕�)!L�Yk������q�5�M����0�Z�H $�e4���/n>^NB����w�RY1�c+.|�md�4�M��_�8���h"��D�fjJU/,�K�~��AD�I�jy�����D������Ԯ@'�f�;+p\�������I"�_o��H�qnW�`���C�H-�ܞ���0{�����; É��ˡ?8I�
�H�)�8W�7���F�9�j!�-�P���@o�k����'��	H�.���������\rJ�6����]�{U���'�C��3ol�_�p�����Iq9��7�
^�n��ĳZ�'�����j�&딗��_����Q��k-��?'E�_�����K�j�6�W�Sr�Gd'�̴�țB�#����k;j���B�jGA��Nt.f��e�W���H��4oj��R~�.[���!�+���&XVE>���:<C�2A��|H7��!�-Q�p�  ��:�ĉ�/rR��	+B%����?\��R��G��l��/���v^�u�P��P��]���1�Vc^Ѥ����.����XMXt��x�����x\��G����3��!�8�z��\������	�ȑ֞�*�
&�ٕ`��![S�}[�w�7��r�T3��Xa���?�s�XQ��:��nP�ïp.D8\�6��Lr��q<۬u[���z�� �C`���9�ZY����?�����u�H[Wv���)4��t>(�B*��jcD��N��"O�N��jd����R��+U�p/��^���M����_�!�nE��*Tr���"��y�����2R�d8��&��� ��}�������g����&�C�ս喝ec�j�&����$�raowQ�ҋ�جk#�h��ps��/�p�\�\O�;5o�k]��� 5�$����J햓&0 �A��ƕ�`���{,���r#?"_V��w�@�²�T/Wɦc%�m�K��0� r̀iz�U��Y�W���IVD%�c���瓆���@RNx�l�*Q��a�p��2/�|�C���E�Q��5���3ᱠI�)�)�Y�"�Mq1�ڽ�$���G�U�K]�k�w,���M�N(&x�Wr�pw@/��Z�׌���O���c'�_ �)\��(e-�{�c��5��T�d���,.���2��J�*J��]��7����G?�j��HNv�K���A�ܝ�^k|��h����6e<�������:��T�s������:�n�_/`�v����ʎ��̙c��h #k?�,�MG�:7��C��SX����P���8��&�,�R�P����� �s[l[�jF��}\j���8#¬No@NR� ��g�
���^x�+��~���c�q���,�J��ZZ`�W-i�����+X>����I�%��<=w�H�*�d��2ʃh=�Dr�<P��S��<u��l�TErOVJ;{@�|����߅�ڞ����Ԥ<z���������������[z��u-����@�HTJ�/,�,H(S�v�l�ѿ`Z�/���[tp��c�4�Q��uM/�R�	.��x)p�m?���1��򦖴r��&_{�-�V�P�XV#�+Q�+�fQgf?*�0I�m~"��qV�Oc���;i��ɵy+ ܮ�ߚ:���J$�|X�>j�������׸v>��~	�a������p]�k�s��QxdQ�G9$?>}�ǫ�YQD���_�Qi������rVjé�\��:�<�b}�wT֧�ࡒ�E	�����^8:_���/-څ�d���k�-=�Z�'��#^G^��_&1���V`,M)���v+�^v�(��X$Va����Zэޢ��zz剢�l�E�k���{ӴQx۵-\]j��@�o��erw�:�B�o畯�'��Z��n�@���{��!��=&�A@�p��,�~�S�3�d+�6�G�?�R�=�_0U���@ط�p1}���)3��L�|����`�A��P���N'�����Â�R����9V�g~���P�n�5����Y6�| ��:�<�<
U`��@�ȣ�G��%���Nc������>����i�T��qWq,:��S �5�(/|߃�kZ�w���wv���>���W����![� (]��6<�h�R@ �A�U֥�wA̯��O�(�=�T)�d\²b��>�}Kʅ�F-� p��\m���dLܾQRG��	޺%���F3ҥ�X6��&�����oo�6����z�ր]%a����G��k;�O����t.��0�ug�uB|jf
��P�w���
�5��Ĩ쩚=��B�����:��K�ޮkZ��z���8��ɲ @���e�S��uCU�Fn�v�D弸���N��^˨|ntaI	�[l��7�E�a�/H�r���t�v�1KG�0�47�������ԱT�1�>��wd��B21�X[iՂ�l{8j=��D�fs�6���&K�" SNN<qD2��f�;r���RZ���FxF!��ДZW��*yv�j��$S����&0��h��'��+ �e��<@&"*x��g:���|Y�&;����5}��, hgN+�+�m�1�3@�Z78l�`�Q�G�c<�Ejei
yҼ}ˌ��x<1d�A��'�i��O�Xl"x�-�R�T9V}L�2e�ᕑ�[�t˕[i�Jc/ܻ=�8sS(+�{�#��N���嫙ȿ���e��<Ey[ٞ�]G6�,A��k
��&c�U5ƘUl/��&�Ї�S��Ʌ�q�(".���̴l�Pՙ� 	���왥����9S�8�c��R��̝�ġ�ѿ���LN�Z�*�������Y��h���Gn���tf���A�_�Px?�n��ۿ�"��e��k��N	�4^y���#��'_3p�F�X���cC#ƈ)iH��s��O��-�'�^���R� �!>J#�FK���m��*����S��jV9�j���2h�z\�ͪ	|��uT��%�]�٧H�����J��_O_�9}��5�ۏ�]J'���}�VYA�Rk$ܚ9@C�hd.}�����5�5��pު���B��$�)�����u�n�M��Ԇ���خ�t~ԯ���-ڟ�p<CīNp�KWX��.&S��'�<![��7.8oXF�,7�/�ў˂#̆�
\�I�ň��2�Z���$�ndS��Z�2�%_!G��y��� ݈n�nS�iW6J�d�#d/����?&�tgh����ݘI.t�R�2�7����&S�j��rm��ǟ���g}¯�����<jS&��y
�e�Ŝ�<P��xj�UEY�(Q�r-Y�I��,�c/mg���O�_z��ХҢ���9$x�!{6^�����'[o~�}�4g��q����v�."��g�J��$��m�����Z�=�ڝ�K�l��9��_��k@,�U��S�p���.ϡ��@.�|�P�Ǐ[XL��R�r��)�(|��0��;��$�6O�3��ڍ�ǲ%��ĵ��xez4���א�
X����.�4�1vUw�kN� 1�A�:X/>���0i�cux����3�9ɥr��RK���#�w����AhO�Y��ꦒ�'#�3������|���L���?È�Z�z��Y|���Hf�C�-��`������(�͜���U���x���vPO�^���`���@�C�����9z�ރgI�R.���V���-Y���7F�{���H4)�?Jn��$�kW�P�;�T�_�!1���=�vD���"C�B�si�{��g��=�PJ�������Ô�Y�n�d>V;�J ���n��^����{����f�sN>�RHy�y
��XrH�1�Fi����~�S� ��д��d�	�hO���"n2�[�G����f!��]0 ��O�c�یॵ՘�|�?�I|��σTM�R9�Z+�p���4i8�Ϣ���k�`]F��U&��gG�W��:�"���Aך�Ff=�ojDi�)P�!��!�6���Y��k�Z��e�����a?߂�@'�T�9Ɂq*��*
�5��E��c�2�*�?���(˹7�>���z4��ށd���s�OrZ��9w��R�IXyu���y��Đ��(�=&�S���a���n+�M��\�zQE~��G?�,j�Va�xQ�@E���pmh�2#{��S᱁���)躍��=�D��*rO����:H��AP���qFϋ��6
�&oGG����̷{L�v|JsY�45��dJ�����!䔰�a����b��#f/K�"V+G(:�qŌ'�w��R����yN�
U�5�ڽ����>J�U�ɔ_7V��