��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,��&VSA����U�i��en�(覘��ݒ��a��������)�:s`�X�-�B9���CR�I5dI��Wl�"O*ڋV*���@��l��o��ᦂ����J��	f�K�u�;��2�z:2f\=�L�Uz��='���4(x�8���4܅1kV  ���%D�n�g��C�۶��)Ҳ��yx���q�zJ7���H��,�����"d�C!�:v^�����}0L��L�M�F3��3���t���w�k�,煒a�Z��k�Tf�P۾�{rW�JO\2� �]+2�ɑ3/�˵����1qR�!e���ĕʫ7D�*��
�!�T�w�P�VU2byn����)�Kϖ3��C�9�&sF���	�(g���m��������	�}��M廮y��B��h�e8�95d�:����?ሣ[�$3x���r��r��׿͘h�C��%�E�� 	g���"ג)���,�s(�;E��������誃{�:����8A�xA�?b������3D��RW"�gme�n�:���
ı`]+p�NZ��/i�>��'�1҅^�a��� ��&�0u��; �]�R�9��ͅ��Җ�姰#�����v��7-���D���zw��d��Y���'�=�)�6�˪a�:�!	Y�M.SߝZZ�ݸ@˲j��w�8Ĵ�w�/v�ь�zL��3��2�d��{z��4�����/�л��Ǯ�o������&�/�{b�
��C=p��;�;��5[��10���,��{�5��07\����jF�9LB9�mh�gN	�x��]Ν:���w#�v7
:{��c`�4Aok�a���eCJҜ�����z[?	��'c���k`Z���x�����:�W]ؕ��q&7�-�_��F���2U[�9� ��8#s�����x~���G����N�|3��Bqp�/"=�Ka�`��096�A��R˱��X�~�S	g���|ʗ����y�|v|�d�H�e��]���a��n]TT�e}wq�oL�4H!o�j/qL>}���X���@O0���^}J6��5p}= n.����� C2�:!��	p]����,5�O'��;ĭ$�+W�i�Th믤K
��=�������#b�nyk�D�X��6)l�v��'X���P6]��ɢ�L��oː�mu.m�I�t��Π��b���}�o>��sϝ^�9y���9���
Q(�\�S�32��"��$����G�k�p6M��Ӈ�j�|�&�p�>e����$98a��-�~��H���
���񙝕�3�`�)!���i���\�1�LPP�ƅ;W'u�h_�Σu)����ò�[s����8�hc�,v�}��S��Y�"��(����%W^�\ ����-Arzc~�Гϕv�S��-��5e��]��N�ͨ����lJ?�o[�'�D1��`sdpٰY5'ݩ��'�J*?���I�vP���e�]+k0zD��d�S4�q�s)�1!nF+ũ�w
�>��f+n��jS�v�В���(R��>��\�����g��YL�c5��0̘�]:kp�����e�"�c��T��p�0���մ���`��j��gd2�Q�!�&A���۬O?*�*�� Z�����"�7A@��XQ����UPnW��٫�+��
�4���waŁ[��6(�'�U/�^\:.���iY�x�K����c�
�'(D�'ɥ��2��+t� ��\�?�0����z	\j{l����*�4ji���ꅋZZ\"�&ʗ�9i9��)���h�AΙ��Z�U�*�Y�&@X{M:=�HW���[��_{�F%��(wWoG0��&"�0��T�n�YDxث'&a�`H:(-/;sCB@o4}���E Q����ZIZ@2l�ڳ���M�	�	�v�[� �t�[�sx��PS��*ݖ��,�BVի�Y�O;��N�ۿ}TL�z��{�*Y'�+s$#�T�}֌`�C��.�C�$oȵRң�SA�v�;1\x�ɶr[�ʰ�~�"�z�G� f�q`9Έ�2䈛w�g)/�/<���&�/nD7�I77�L׺rm��E��I�7�{��sL��