��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c\�esR&{������o�T�e�Z�/��`%�����1�2��g\D"[ޏ�F�
܌�)�u�lg�h���T�Rfd���pD�e�֠��:yc���?����ߕr�p2�{M��r����u/q�[s��j�x�`�{a�|�����_�Qv�������.SbH�nKU�2��4\�ʿ�PvOl&Ħ�^C��!F�<�SY�} B�V�?I�c欄a͇#��3RQx���	0���''���� Ĵ��s��>����3����J�[qy��V��lG��i	M��������E'ي!��3ã���`*�S!��#��s�T�
�P���zC�$�"���a�l5�6�֖��� �>�<zS��R{ot�ߝ@#��8ٌy���-�S�-][��
�{&�<D�ʠ��%e��d�W��	E�8�3܋�k�?j~>Z!i�]1ɕ�x���h2��Py+��^��R\T�U���b��.�A��@J-P-a:�fl;^����Yykb}�|�&�X� %5��W	���U���4G_��p���T_a�o�
t[߅FKT�n�WL�٬��4߬=���5E�NA�ߎ���DPާq^6i�b�'xV�,�m7�n|ha;��f挥r�Lp�*�YB��T���=p�;-T#{P{��XM��a��0y$0�������k�8ٞ)^ 71�OG�MC���|��G�AI�j����6��6u>�*�O���&�>Ks���3{�U@9)n���o�k�)$�p�����)���څx���hQ^8N��\�OG䟨��5����� �Ǖ������½3��|	�#����]ۓԽE�W!f3c��+���֌��N�$�xe^�;>.��\N�W�̫�h���0N�_����n{ހ�\�w�V�����W��9�����&���H;̵�>$���c�o�;釫���h���D;��0	���ߛ��ȴ"n�B��+>O�-("fSAbI��|�l&�l��3I��V�bκ�o��`JH���CQ 6�T�}d�2��O\�V��9f֭�wɉ�[��W[8��JV1\z�Hڷ�p��i��>A�Uް�qN�w�{�f@����>�9Yw~����)�tm�5�ALՑ[���+�SC�|�2�jaj���
u�+�y��Km�l�����M�W�,�LL�_�]֠t��Aq>ȯ¸h�8ђ�
5��ɨ���J����� zb���;U&Y1�zd�4�&���H�m�k{��e�B�"@��Q��O�Cqj����hˎ��uR���Ꞿn�M�+�����bo�?�2{v��^�1�F��V��RY9�1p��TAf��H�e�B��	�S7O��+��H#3`�95u�YD���2�wA�ׇ�P�-��q��#��1�}#/���pD�B��Q�ܫ�=��3�R#��#��d��/B��D�M���	UQ6�����˦�Q�hi�yy��D��xWF"��3��x��Ǵ�B���B��8<�y��=8a�IDdb��[k?)�kh�fL���]�ӖU]�ц*����\ƒ�KY����$6�V�kc�����0y,��E�-ڗY�#������ι�b?0=�d?�!H۷�ur�a���Y�ᬹ�$KD̠5`4��(�1��J����+ΜK  �
bO����"�iFs򑀊����ڥT�\뒊ǹ��\�jz���F�������	�9r	<�B���䘃@����UDꀵ�	��>�Q��U�IUF���	�˗�b(�y�pqR?thr;�\�Y_�m0��%7���f	�����`b�v�v�Cn�j}��_m�sb{� �d���yǺ�j��߇��*55'��[iS�3��[�[�c���~��b�þ�����=��ĥŅ�6S��J>�CĤyr�%g5�6V��dN�P�TFU-�,�'5����.Q�c�Pp�V�6Ů�`��`�ܚS�?~a 0_$��%�46tW�O��Ű��c\a����?��+Ș����wX)�p�|��_t�KO����\�l��\0$��YJ��@1,ۉY�G�-��,$cOtP[��J�FFp��&���W��P�o�B�?���2�n��=ː�ȳ��=Ŧ���d���wO��f��~f56�!^��m���h�X��=[�P�h��%�4*&-Tm=>!�:�v�r��ZE������<�;�~��S4�8��;g����.:������S�{�F4�(f�c���L������������]�nPt��A�a ���Ӓk_6��Rk�����:���0i�6#(�J�Z	L�v�� J�ĺ9̾*F��Q�J�E���p�=�R@���zvp��qz#�z���>
.�"˰�OkMN$�4�x%��
~��@������ o�`�Z�%��m��O�\��� |
����X��w�7�I�e�ܮ^Zza�B}l���E�f+r�F�ʧ���ɂo�H����"�_l�WP���h�FFR\W��f*�����;u��T�� r s��3'+Q�/D�A��KW�'�%%KH���3���:�j�1�ϛ�L?c��P����Yuxv����?������4�D��^�� =��s��o�MB�Dڣ�*���7a���t�b,>�U���c����i���^IQI�&���׊���W�� ��\�|M��1�Q�m�g-o�RV�.`9{��8]� �ѭ-Q�5���GƛKt*�M>����6`��nSΠG �4z�Y�=�m�!�F=�Q:l�p�T���4�y�.Hbp�Tr ��́����>z��z�m?�*��0���m3�d�.e�o��]�|KmӜ��9����ણW,��Ej!��]�g_�*����wK;��?1^t�j�Eh�@~'����6a]���E�ڌcJ���h��N0hϭ��` �ls��&6-8:$:�b�y����6�DPƫ�8�|do��.�!D��V���s�)�?�1@RfY�Gf:��B�>k���,}-��p{��l��Z�Ur�^+�͠/�x�|���X^
Us�����l��c�k��k�7����:�|���I�	�6$.�)����ȝ�'�g��Ȕ���%]���DmB	�@���P$����D|ƠNZ��_4a�]-g"cBN���a����k��WO�T���$Hv�h���:�d�&��e�vl�cvEpr�ܼ�U�2�l��� m�X�_�'N���P�iaT�w?���`P���fP7^x2-N��XI�����UU�����޾:��.L���	�{(+y����ΙIq�������4�7f�2���f��|�<Ɉ��A��a�g�(o��i��g��*�_��}��#�IvĲ��'����V��O�wZ�o�n �o�5��;�[�[N��h�4�'�~������hAc�W�&�9�g����{S����+t`��B[o�����@���IU����q�؅s�me�
Q���ڌ�G!�QV����]���19"�k$d�D#��ꗈ���5ti�nj:F�4kc��� ئ��G�k�>���f�����	���ؗ4�����L�°#����u+��:9��jg8�k���x�(�T�b�o"'�¢��Eq�
e����w�hs,�C�,}9(�D�dK��B�|C�5rD�zQ����`l~��3��F���������y!�����xC��"�(2���������N����Q��(��+�>�bn�z݉��!C�����\����Ua~��<�<M��,;
�Gr#�,K= "1U�:ᴣ���T8����n��\
xM����!���K�X�>/%~~��<�����^)�uiN�|�4.kb�z =-�s���@���A�@�ت�[w���Q�|�����QZ�%n�|�ѕNF�U�e$�(�R���RD7QC�X�wr;`�ѫxNo�g�a��2��.�) ��A�XZ��� ���%�-ޠ�{���2T:X�a�ekT����sc_��Gz���}&t�&�p$RrF0�K�?�pih$WT*ylY���V�XA޽�|��v`�k�!{AeE�Te^``	Psw�0(E�=�F�RbIy,�j���s[�ߡ��T��Y����7.x�xz�����D�� JhOf����m��>�پj�G1{���o1n�}*?���6RRq��<�:�-���(󋞿��ܯ�O�6ԅ����H� ��1c|��o����� �rP��ߒaSe����P`��C������b�~@%1P�Z�������vY%6�w-�~�!�z0@�Y���8�ch��^֍��C|�`Q�;���w�0��?d��)��`��1�]ȟ�2�!f�N%����b�k3���mwהZ�S:�A��L�\��j�%Dv7���&X�Ë�W�L�6���i��	�LW�b�~"��&��:��K5��D�8~���w��t�����e���!���"���Ň�,����Smr���GG�R��8�8�d�^|�o	?ʻ��V����B=�7a��E��>M�T��wפ�,#(;l�X� O��Mw��������?L�<
�/�<v��RW�Ud����������'�o(Y��_'�[����T�?�Ur���
�v$2�#�����?Fφ��o�H��e�� #�6�\�x���?baF�ӑr�(b�V/0�C����lxq����d�ay_\#��4�����x�ܟQ�I[�_����G��C` ��۟eJo�!Y�����{���M�̼ׯE�QIX�G!C?��Q �(V�"��TF%xl�am~�@�!mzP��Y��8&h�_U�G�ly���-���
����1J(>5��ۇ�N(�$墔�I%m&�h��w'��z|ޒ�1f���!u0�U"+��]M��aČ��L�Q�oV���f*�j@�M	�9X���Ȓ�^KL��k
e�� ��T�^��>ȺR�Q������¸O�ڛ+1v�z��.���܌3\k��M6��<EbU�@�p�qL+����ܽ�y�PI����!�1w���ٓhm1+:<@r���>ș ^��r�w�qY �5W2���j/��z�Cɗ^�U=I���W�\��pf����Ar �/�Df�MB��u]��F�p7�����c��d*¿�y�}7�2�Q�p�G�j����a��Ԏu���%�#	�X:���?Fz�­����xf�H`�K�fB������,wL�z���������d��s��i��;����NO�����^����l���R'����~0����50�����o�O�;����\Q�n��ށ$�X�Gb��`�z��[����J�>RX�zo}�ҋ���������hy���MVM�J�� ���,��T�8�hw���}��������E�]Boe~u�<�ŠM�L]�i#��T�GݣfNL�7������������C�������8�罙v�A���
3P������|(�@�;��'2p�M]��+���,#+c���SR��Pv��d���W�[.P@�w�$v��W^��1�g$�f��X���"F�d�]��0�{r��Rb����>ȱpK�S�f��r;�z�e-3�SM+@ �e�ܯ���v��1��nF1֖_�3��\{�9��;��#�vK�0�E�x�k� ���#*kW-Y���O�z��4�?o�Ɯ�Tb:>�B,��������	�`���ǘ�\���''?
x��W�k����f�s�u*ȈW�lQ�-Ş�)�i;��-�H^9_Q˦EM��I����@�A�����!��k���4�Z��:�T���=m#[�L;�:�����2��
��`1�S�c���l`p��k\�}��z���P��y����}FHws����3��O�+�g_�s�k�nھ2l�0�����9 ����8ހ�m�n_CG]X�&�T����k���!�.��U(+���Ej�U�66Q�
�5�Bv�e��q�V#P����s��	���h	`~6��s������s���jɍkH	HF��s�Yf���0�t��~���l�� "���J��7���i���1'����0�#ӕip��A-Y��J����0+2���υ"��*��{z䤲��;��m�n�,_��o��a�6��	�����nb�<����PlĴ�y��W7����~	L&�%��C*�lC2��q�ū�v~�!�SM(�c���A��C�\�ٔtq6(7�,��Ƭ8�a�\�}`�y�ҸC"7�*�gC��99�k��n�Wvc�U�d{����>�kѲT�d\Y���l1 ��j���nS��yiQв�6p�����%��@p�zgUH��v�U�����u�~0�Н����i��n� �+��,Z���=���Di�����M�j�?��}��,Pc�VȐ!
�+�����펜�%ŵE�d�5�#Hf� !-���-��6&��Ӫ� B�Q�B�XT��Nlc�+�Dn���М������G?Ƨ��[|�����D�S'�b
	E�������M!ȣ��(O�1�`�g�{_���wc��j��iE)���h�T�a��[�1�Z���▗���<�&1M�}���"&��A2&�D�����h@�R��$��8����G���aO�ef�>�����+���1^x�T���	���0���w���[�O~P�u��DmJ)�z�z��/�ʇ�S�ǘ����9C��,z/O�K��UY��o�z]c٭+��������¡K��S��+�w�W(���ݞ=�f��Rz*��%�7Wc�cd�b	�HF	LNuڵ�;i#T�����������;�1�V uVw�#���%铹�6�XDx�p�eKB!_0�w'����Q����c�_���cr���<),�"؋�xB)+˵�q��1kuk���\�%N9G���X�`�{�IK�L���3ѿ�`�W*���v��b&�b�fk��w�w���5���ǌ��1+Y�k�+��ɷ��ԟ�<oԊ��^�W��q;[�oO�7Q�3l�@`w��u،Җ�z�E!C��y�)C�Pq{ ������C���,��w�\�yf����,��|�×�%3����Wl�H�9�xL\R���-�1PX���Z׾
Z�m�P���_VjL��2��BP�*D���e���9��Y�A���n�?���C@��$�@��+@F:��iQp�����Q�y-SR�ǊnA�����n_��0����\���Z
�sB�sl|Ȍ�eJ����J>_�d�y�*��nc��_���������P�H�߇�Ժ8�B����B`n,IlF��;�b������.V7�hvt�$�q�#d-�3|!���w��]=�~��Vgʺҥ	7X�Sd�)�T�!���
1ZVw���XvX~:8�����@��}k��9����q�gv�]4~SԐ%؜4G@|��EM� KaPiФ�^�aF�xeӐ�T<Œ�0>	�}!j�f�p�����'��$v������>���&u��-V�1=L x�"�XaXE5��D��df�W��q?�0!� I��������w�y���ߞ5>G�e���mhѩx\���4��hٴ��������?oJ#G<c&͂��9�|t,EIr�������7P��:-콢>&r���$��NK��nA~��Wi���HH�ՠ�X�2MSL@� ��(��Iq9�9a�JuQh�� �Tj�sz@(�x�y��p?>Vb#�؉�l'�KG����Ǻri�r[rd�mZ!�Mǣ ��ϛ1�U�"���C+�攸&c��}���Į�@��|�3�w4G�i6����L�Cq�ԉ���q�ө��\6����@�a�M	@�	��/-���Ӊuα��ݿK$Tt�]J0Cp����=��J%�L�o�nGIk��	��,�<Q�upw�8C�|dfZ~��ە*�Fϯض��r��4q�A%���↧m�t%�0��[O�L@+��{�ݿS橀��2sƂU�0]5����$�o�a2�r�rv��V �t�T���{�.,N�4�,����[~��6O�# @�[����ߤi��#76�8����j7�k�ж�⪾���B��'�v��r�w����s��B������E�s����3�j1[>m�d{�UC֗��>V�� ���DZQB�5�����uL�	j����Z�c�4��]'���&�{�V�&�IE�#���A�)�	�x8R��ϔ��1���|Ȯ}�J�v��N^E�s�Ci���[��@ƨ;[���!f,jlP�����a�:�Ԅ�� t[8��?a|�!'����k��&�x7s�!�O�\�d�^�V��M=���F�����pL=1^�>�ͦ�{��b��K��x7&���7��/Jf>��M]��v���z�=I���g�{GP��G�����d�?yU��%�}��A�>K�7�ܹ�Tzk�֞�����ڷ�>F^-4b%���ĩeK�ɞt��LryQ�+�6|m��S¥q��zU��.g���c�F� 0��ģ���^(y#L�qf4Ն�_�����S��|��c!�C�f)X�Ҟ���(	� �q��;�Av�w�L)f��rPS�+��m"�R�!�"2-�#�h�aǅ�����t�25UI�yD�m����r��A��Ce���Q���FLx���Y�5�xQ�	
�	g����)Χ؝Fꈇb��x��ù��뛠o��R����#���<ś\5��#� �bi������.
\0�O;�Gwd����tȊ��E`cÀ�n�V��?���*���ȃ{���-�(�Χ��1p��/�Tqrs�?h����Vv�k���L@}�K��w�W�;�g/��!���n�~*-���۞����{��9g_�K�f�2\ �c�/s�
���Q�?FȨ���]�.�0p<.��N� 3�6�z�T�����-��_�x�
2�_��\����$V������lW.'�H��H J�pz*S#�Kܯ]��t5���,��2�~�b��u�OQ�K������.����qex&�T���G[=�tO���k�$���ˋ��x��2M�
������P����':�^LWlFe_�_�c�!������pt���8�Veڜ1�t�3�(q1h;ۋ]��n��;�3��l���8h�����>�F�;�uk+8a��%�Q(�vHg/0�V�/���.�e-=��2���l���ހ��?�qC3ZVg���$k?�����t�9?�(R��u�tG/&��������Nz6�6A���5x<���,w�4L?݀����Rc]񋁵#[��z<�c�c��>����b�u{WӀ��O�<��c|W#������HG����TR*(n�N<9����;mKnT�UH�+JIU#Vw��W�\�\r���2���f�VQ��~�W�����P*<N�Q�&��6j�vp8��U4�(��_�[&.�t[p]~Z�����Kj����@�j��K��گu���<h7��Qɭ�A�o"��q�jSy�g4Xb�S�	O~�GiG���f9"NX&UO�oR#[��)�N�P�| �Z���7E*�.4Rl4R| I�iw-!/�@�*�[��1Ձ�N�h�<�¥�I�'A�(5�n_�mt���;�1��0�f��=�y��H��`�X ��glO?����`�`%�V �J`_P6o��X���}����i���F�-�B-��D�3�U�e~B�F"^㱴��?�7�y�8o��e6T2V?��F��(h v̜��]���v��􂣰���/g�˖�gɯXNѝOY�H`��"(7s�K����$Ԧ̓����J�:������O�"����?���b��w(�)�2��Fr�U��ql}`C@v��v�-�I�}�am\�ל��M���������H���_��Z-5��G �\B|���">��t �"�QR"��?�6aQ,����@��Ssv�G��xd�g�w�p̈�rE���]DȢR���~���`�Ѭ�w���N�w��f�u �2�#ʒ?!Aׄ��XZC��[QqO�t�耂�b"�n7�����.;>6	�X�H"��2x'ꐘ�؉S�U�-Ħ���j���@�E_i!�$�>��x΋p���+�A@�A�`G ���ҁ�x��� j!�@������,�3q��v�$�.p~��4Wf�{#z�o����X&�UQ.���Q��N\1/��݈6K� 9��z@�$�������W��o#
�i�lT=������塅�}5��<gY�3ؾ 7J˯�!]�~z�:s��&��XYB$�$��f
3܌Ɋ�^���$��bla�<�:K���*&+�Ϭ�g�����q��?�`����m�͚���Z8���,����3�m3���2�>��p`O,w
:q`��d�ͤ<_��,���Wk��,'�N�6B^��ӝ�2 � ����l�d(��Сg�W+�⠇<=4~R���]���&_�V�
�+]Db�F	b]8A<�߀�]8T��׳� o��TҠ�oؐ��r?�{�0�(�Z/3@�o�7��񯺺��e��r�OY]�W����9,w�n�	ƍ�����f���'�裭u���,��=�TT�-�Yr��,e�z�Zw�)�s�[T4^�謹��YTĄ2�q��^R��3
-�j��ѡ�Ag=�XH���{t��r{�n��}8ۄ:
@�V��ح����w�JJV��4H���6]l��7wxA�0�V2��Ip� ��J�(pp���7�H��p���;��eR<�O��E��J�R��^ǐ����5I���.j5�St�8f�Sp��M�Ț� �"��<�G��\������n����g�at�ޅ'L���U��5���}�k2Am��pv�of<T3��+6��t��*ω�.`�kA����V����_:`��[qp����>r�]>��ñ����Ye{m�G�د�ː�(��0>�s�(���=�?x6Q��5���@�uK�K�#65#*�r��4����I[�)��J䁉� �=la=M�������Y�<͐���y&%
[�\-�5��'����ͧv$��Pdu��Fzb�Y��K������$dEh5��	����y���
�ha6��D�-�&�5ހ}=ɐ�JUV���K 5���K�hPdK�2��՗�dp��lW�1�S�c��\F=4�T�MthKQ�a@sg&��ϊ�-8z	�Q-�5u%�,�������hX�k.��
�Dg��Nwp�F]�ɴwR��鬢-��64/��I�aH�[��g����������y�L�<�Yir�|%�>P�Пt�M���Z6�4)ҤЎRX�e�ay�$7��N���U�erG����*�1�� [Y�Y?h,.��V�d��i�����B"��W���d��͈��f'�/�EWyÚ8�F�z=l�����1��p��b跔
���T��X>�{ǩ��贗����7J�B�.�I��芅>�����=���b�� '�~���B�u��-a^�U�=Xf�L\���ю1<{�h�}W�z6����'rFo�Gλ�[����!��u�jg��WA����M~�D�*	�F�����"�c��M�R�,�;�6T�3[�(L����P���s�u���=�CXӞ)�����\�^����+d]�釆������\��kg58=�Ϯ�Gc�/Dyc�Oo�"�J��釸V
(׶��a)�=1d�ey�R����טG�_z�9Y�ѿK������{:�>�0ǋ)W;)�*��ƶd����rD� f���/fR�z�,��{D^0�����|��=�op@��y?��4�o��D�`�K��qb�W������s3�^D���;m�=�S��_e#"El�|�Ȝ�k(�n�����YvUj�PD��s�h�x艐�)�K�
UJp)M�xߦ��RNa�a�G��e��e�3і"��j*|���Fv�A�;2�<�zKx[Z����ׇ ����@>���+�H5	��+���C���?j���{���(�F�Ĺ�pX�����WR%�B� �oz]/�ҏ�`�2����q�흶%@��^S{��]t�����!AD���Nygz"��pSq+#�=+k�+w/��O�ٻ��Ʀ9��r�6�38O]��)O����e�oPH�H�������6d�bg�/��;pdl �3��_���wPF�e>�$�3���ޝ�kB�د>�ݭ�m/����x�
��'0��]���?@����ƓcD�g�j�Z��,J藡���I:�V^�|�#dTQ��h��F����w����v������$�����@���ə���Lg�2�lSQf�Z��9z���Ic�|�.�)T맾��q�X�\�M�ʜ��&�WPZ"?���4��JGӞ~�/�&�l�=;�w_E�:E���E�:��E��r���ϐM����9z&_ы��n���Z�z,��рp������+����=�b`u/�Q,��T �0�v<B�r���A�QB��/���|6�r��M*�:�B�bJ��$,?�cs��}���7�Y�_m��T��:�`���ۨ��t��b����b������4���e)O�a���4�����\?Z.���O�:g�a�3:-"f3�_Ȝ�'͗N4��nG�Ǒ6� E	�s.�N�N����9�M4��4�� J�}:�jl{p?MЊ��Cw��ջo����ݬ�h9�:y��t��W�鄃F�ts-=���|*K�haQ��<$`~�m��?�����{h�\�Cy�ӊ(��4=]2\�m0J��0��E��(A��u5�b<����e���x6c�AbC���4�6i(�Z<��Ϥ��e9Y#$�mK�uTU���q��N�-%��O�Qd�u�)a�)�8�ŕ�D�GŁ�5��&v�v�Uk�v��������5>S_�7�h��^��5��G��sf��8uE�^uN-1c���B�ZpN��U�1���v����0��*]阇[��$�n�Y��늮�b��5{AS
�r3�&�O"�!F�Ⱥ�%+YȈW:N�y�)��ĥ)�Ś{�=�F˝�Ai�󮎠�E���aG�vS�� �=e�������aQ�*��2��MT�|�����u*9����\��ζ{7���͑MX�K�S�����W��3N�R����pF;�g��I�=�!f����N����)ekm�w��q�ʮ	e�g��U�m�_(�GY�|YfN_�ؐ�xoUQD7ͼ�Ss!ݿ����������y:��7��+L\`��!����k|��r�Z��{=�����r��rf��L|��Ȕ�Z�Z@U��|���\(�<�$���q�i��"��\�YFZId�_#�R�<亶+��c"p\`�?\1[�/Ş�q"�V7�����mX�H�ťAkJ�/ˬ�
�(!�Z9����}�1۞��X6� �ҾiWa+�������,�v��E0�+��)/mD<�|�����OНB��P[z{'!�dj�G-g��F�X�������QFtYy�W�nlN�����<�QY4��m�b���sR�K���hV}�Rӷ�}�
�APxl��i��@��kt���Ykp�㳰���IN[*6��v'Rެ�)F�ȴ�e�C�@��t��:�m�	��@u^���R\�f�%Qf����?�(����*�ژ�w-��k�����Ĭ��Q���{�q k�W~[,�D	}�4��7�B��-֍& ޥߦsفW�IG?�t�t�s��&��RF���������ة�=�� �Jp��k�L��G�װ;�Ȃ�=(8��P1��D�`� �I�\I��pwZ1m:&�Bo��c�5���6F�D�G���ۘ�E!��K��� ȺXF�7��V���a4z����zA�ʸ9oX��~��~J�E;ٱ�e���.��� ��|��/�&61_r�Ag6��!j�7��,C�s�@Kq��B���,%[L,(���N�!op�����B�y阔�Ϋs)]��?(�KsyV��s��X^�� ?S�G$�l䙆���B������U�{9�!���_�9<sXB�ͧ��/�0*�.������ƫ��]r�b��1��dE��%�.M(�־�k+U�D���[��]���M�a���p.�5�x�F�"̪��w���Y`oe��m�"1�T��']!QcfE�Yy(���� 8�h;��־���(�#��Y;��E��D�eV����VKV VI9N��R��a9[	� p�Zxq��@�A���I9�p_�'��t�jI���P^�F$�_�C*}�� CF�
T�*�<���Q}L�o�H�� �1Uy&�ȩ��ʸ�1ႏ���7�����3��貀2�Z��g���9LE㾫��
�{� F|��3�֫��P ���{�Vd�� � ���3�wHX�)��� C��J�����V�K	��Ev�%�,pP���zU��]	)T��.vet����f�!_>��́L�!�>�ag~t���m�q�!]3S����o=:�*7�e ��ZQ:��
�X0c���ۉKw6(3#W<��b�2̳
:'�n9������7��RϦ�<��:޸���cҕ>`����t�3��Me0��_ѿ^�|�XĪ}r��?�jo����4S_�������T���Ĺ�#���V�$�{`3t��f�
��%a�W�.�[���kY���l�z��Fsf'l�ש�R����'���Ӱ[���d[��*�����̩��i���
d�t"���9?h���MU��:�GΎ��94",�y�<�+\�X2w�@�`W��*�|=`8䧙���CQ�C0PF7}����9����I+l`�����L0��*�X�mt!�M�����Yd�c��|�����Ѫ���K���	����(�,�P�ܲ~��bj]����?��R��c3R�xw��å2������Ϸ�m͘%��@���S��w�W��R�q�V��GV�˱�#1��aerY�v�tG��  5�7�{���^-C�\cI��V�A���f0������m���jC+�P�ɲ.��Q��Di�r�\�;� ;R�R�k;��/���O:t��At�d�����L`��E�Qz�CkE|��yU���-��<D{yg�>�.�J��h�!�Y�0���CfB)8������c��G�z{�0N��š�e�K�o6! Й��✒A������2� {����Y���d���ĕ�-��3sr3fI�d�S��=,d��@������烡�!s���4����u���X0�ƺ��Y�k�'�iɊ�%��t�>���8���=|�>��A��rć����E%���� R�ԁ��F�н}�2��|�9n�}&�q�6�4�����k��E-Yާ��Ǭd�ՙ��OBWۘ��c'�ݏ+ ��L�ە}�W=�Q	����FDS��텎#�3&cσjb�W�&��/��\b�&��`ݟ�'4!f�0���J����f�Ї��Q�OE=fc��
���ӻ����Jj���LǨN�4�z�����8�W�2��Hl�mA+0y�N�=o7M�շU*�	`��Wm׆o.\ܻ��[�%x���r�H�H�DMK�P