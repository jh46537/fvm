��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��ߨ�=�]	7�N�)3�M�Ρ� ��B
�i�k<֐�1(�/h�"�+r��ҏ�X�fИ`��6.[���L����Sg�$|����x���
����v�95|b�fUw��e#���`r�|�QZ3E�*��e$㩥�֢H.���a9��[��}h��P����{7DI�y*��f`�K�>BW�{�����z��<�	&u2��<��q-F�zB��0�t�c\��L��U�Z���T�u�o|^��G�)�=�d�so,�yr���o�L1/�%�o ��)X�A��f�H9=<~�/�f�ԑb��ޝ��X����3�5�_�O��AX��ˡr*`�}�1	��83pPR]�B~ƫ�ug�D����2�9� �����/E=4�pzD�<QCY^��}h[
KV �����{��g$_�_@�6��F��7c��m^�<E�������1x2b>�HW*� ���	k��q��f��˳��9Y_��{ﯧV���f>i�E����uң
5����Ky�$�8���kXE|�$������G�OBE5*�,�Q-�^��L���\ȹ(y�1���Ћ����Av�B�J����奆Y�ѳR?��"��a��/��ae=�@�5)޻ۛ��_��3����Tr���kA��MM:4cx���Eh��JR��P17����,ws��2���A���V9
�l6��� C(�������?l�{޻���'��1o�r:v��� 7�
����㗠�LYTd��~�Q�k���k
���a�eRy�LH�Є,�|$%�nKV�M�\��πAC��Z�F���Z.�уX�~,�n*�%D^*�4�J�tc5}�p�c��ϟC��	�2����%�<m���8�O�b�u9n��SΔ��p�F%9���#t�����cG^ln��U��zR]���A�E��5�ϵ��1;�v��j/�3�����N�ć�� �K�Փ�1�_5`�	K��\U.��F�Y�ǯ]�H��r��T����n��`����(���؎D�v�mҮ� ]-� ��:" �8�Ia�3�����U 7K�(�M�k�f=7���.v�e��`�ԣC�������~}+��[��a� ���L7c<�2޼�xʛ�U�c�v�{aۇ�����O�[ �IP�������#Xr��I�4�Kdf[Z��x�E�X���-�˄�Qe�Q�ϱTi��;# 3����:�<�I�?�X�%���|����3:ŋ˧Ur����ps�y��p� �������ƈ�dY__��;��=��j]q�E��, �J���\*�z�3�o���iN#-���A궙	�0�1�~���I0��?���\zY�?Nt���<�_W�M���^�:��fY��t�J{�/�Co��L�1����'D8$
�ª�xbF�f[������6+}�G��a*�B���	���g��s�k���O���}���綼0v$��l_�Fɏ3D�	�<�e?a��oQFĖ,�`��pkkl��RZ2��Y(�6O�1r��LS�K��3���j��_@� �*K���.�[��^2�3Cu��R"U܈N����|�n2���Q�m	�<�u���*3�������kctk�)+ի�zڛ�K~�w����7d��~_v�a΅�D �������O.㶖�_G{�wz0x�Ϯ� ����gC6��8�f��On��D���-Tg�eOu�U��X�~+�du,��E�Nks������"]��?j��DM<ɶ�a�.�^J�7������WyG-����G��gbD�Ї���Pn����wK�x\��d؆�� U��(�/��C61�p��f�'�<A����×ZGp!���-h<A��W�"ħc>�����q�Dxs��8?��m��;\4"A�W�!�F3i�,���0z��O���=��=�뺶�p�W/�bd���8�s`�-s���Q\�H@J�<�^+c�w�s���=�{/M��a�9�*����}�oW�ҩ����@Fi����(��<�(��79�j�s�ޑM	��6aa/f��:�3��c���;4��c����+(ZK��Y�8y���y�mIzր�����M������e\l�lk���Xa&��MS���EB��nF ����P���/{г�d%�ʤq�H`z��Fp��1���os���9��^��ʢ�Kr��Y^H��)OST�mC�q=ԖE!u�$l��4�pz2�96~�N�^l�����!�z��l �E��]�����Y�0u�Fj�s�"�^��)W�Rԗ���lL������x	�4��ػY��C�N�&��G �3�@@�){/>�˩� oOM~�!�&�����~���t�.�Ӥ�)˛S��s�$�n���� �@���]1���$TT��+W�}��lƕ1B��w�H^�N�i�da�vq�$*ZDb�X�Z�4���[%����v��@
ʾ���;H]�S����,�yh �5���!H���y`R|��I�ʀK�袁��s�#���Lh�4^PX\� �v{�����V�s݈:k�6
;JXJx,>�&��;��XG�
�(��'w����ܐc����@H�����1�����a���$cM�����Rv*��j!�9�l��"��k37��E��#�9+���Q�j��ՙI�ge.��I��xa�^�V����Ǧa���vx�%�7淬J�P���|Q���$�
�4��ƺb�V�ܝ� ��U0w�d;�Õo�G��{���E\^X0��uYur��X��q4Y�QY��"������sbִZ=Qӝ��xF�սy�xEʯ%�nξ.6��Z����萰J9�,*�0�ڏ�&�_<���|����:Gm���h�˅h�Yj�CW%��A�B�BqɃ��KVr��3�Ej�;�='����ʰW�2�����bY�����O�t^�#�IN
Q 5s%�VQ��EOK5[�I ���Dͷ�lR[ 9�+,�nZ��Y�	��!�	�W�BT���x�s#%/m������_t�@��E��NS�uVSZ�`zsn�Ήe�X�5N���mz�� E��͞C�����c/���s�P�+*j&\�$� ܦ��^��u	Z��)ܛ���]H  Iydo�z͚#Z�܀��3�Yt<��+�Z�4�J_�D��G�#W^���<�p<0�	���q�|	cCp%`^���L{��R�L5ⴒ��k~��6-E��3 �1�0l�^ �� ڏ0֛g��n��y9�,y�N����	�O�wd/�q�|�q�A���je[NΚP���3�L ��u�<d�銲���C7>���%s��
�PdE���N\���c��#Z��GȬ��d�"��PlU��,`a�j&�c�=��cE�Z�N��� [���a(�;�\�F<{R��"<��;�[W秥�	�Ef���vً(p���e�,�`�m��]>�8i{O��GF����#��������	�wJ�}ITǵ�'BI/n[��y�H��G����"�0޳�Jk�r�6u!bL���ƄQ�~�/vY��N�����H:�K�ܖ���9hAbYz#���l1�8�7�1M�ѢD�ۅ�SX
�r�m۸��P��ϱ|�`�ץr*��� �bJ_2��9f̈3�Fh5�/@_;>~�忬��|��(���̇�Y��p�4^=����{��][��r�:����`�8�D�ލv��?�\4���6\t��0��CY��^��"sv7#k��0��f�2k�����*!RI�L�e�	mmX9N	L"1�1.���_z�c�D^yAb�ܹDQ��j:M�x�)�Ru�Z��"sK&�Y>�tv�A"��礧�9�! ��ERӎ���r����\1��1�f��j��}��+/6��Y�`�D��$j������t����)��#��&
s�����
7�:v�~�2ǣ�'���	{�\֯˒�g<ģ4{�L���M��En�)G0p�a%�@�>��~\�����E)T(C!�R�B���9U����oaG�߹�z�#��w�X�'��	����Vd��]�
���8�P���{3�pTGĮg�늇�s���(G"��7� ��s%��簻?�7z�ب����̈́~a����U�%�j���6�0�'�}��B	_��3ъ��Z�?ɡ��,{��Ոg������BH}-h���0�,��_��!O��U-��&�U��`����M��=q�
��TW�B�W����������٠������1�փ�t8RENn���mI(IZǦ�A��]Ћ6�Yz���/׼uA������=� Zq*�O�<��	�� �s��$�ȷ�D�Id+��v1!��`���&�Ϳ�N@6�Q��~�Pq֊Vt=�`�������R_l�0Gx������`��Կ+�KՋ����AѢ�EM����>U�S�#Rt����"P��ldY���[��k�u{� �����1>c]���rc-���_a5}�����H�G�{����kwzF��>�B�dl ,���"8���y�|:W�" �lA�\��p} <{�m��;��֡�pd�Yb\�+@�_ ���'A{����{ð!wq	8ŕ��]�%���Ұs�ԕ����'F�x���i�����`��f�[$2얶X����Tf뵟�؝i�K��*�s'U�*���_e�)/m@t��gɵ@K�ǐ���7�P�iT�b�������5��r�u�
k�ֿun�6���-sQ��6������y���I��<���]���.N�c#K����r��IA�#�=KB�3����r��E0�?=(�}���hW�����H$j[���.D����w�V�wO��\"�y�]B�,�r�H�\��Ȃ+-.����O��+������ʻ �����Z��豉��/l8�H�>���C=�zg�!E�wL�=Ői���u��(��2Ns�^lp��Uۈ��b��Jjy�R쯡m$0Q)�����x�y�5�﯎@���4���3�C��f�+�X^
�q3�e]g�W!�$�vC��|�NVд�~�#<��i����+����d��<
m�Fo��?�3T�%�s�<���-����S5}D0;iM��z�3s������P
0�����_i��?1c3���Fx���O��vIP��5�a1��p�e��Pa4X��'h➮�ѵFgI�3�i�O��R����'�w��tZ��W5f�z������Hr�6\�ͬdά���Z{��9�c�� �������@΀8����@u���_�,�M�\�_B���j�� ��\#,�:���E�)���rD���N�ѩ�1��E2��PG\��coh���3\4Ĺ}r�Ϣ����ᙦ?�#���!*��W�{l�;j!��E��O�W�d	�qp�� �D�6;(�.�oV0_�Џ�)5�����`]С���y=P{���vx��H��Qפ�ҏ��nKO�F�S-uv<7qD�ˑI�����wo�?B9��F-l ���Ŵ�xd��#�x��9�ĘMNQmT1mS�4���3~�mPGH�yq �SH�*�y� xÿ�,�eS�a�8G�h��%����Y���B�T"q�vw��`n���䩝�g���m��Ms�7עZ���-V�*G��<aOh��e!^ݱ���wy��̗�B��9R�����:*�_]���"��;W� ,q����i����ަ�-�j�O5�|%tH�(8��v>SE��~&�=/3�}5���/��;,E���S�`t���
IF4��D��,3�D��VE|r�3����b��IfC~���ݹl0':U#hn�3
����Ɲ�&۬��vۅ%�:��0�B�M���	Y��H�*FW���:9�0Ö�����B��0�1��^��_��C�x�^D��UY����)-��c[��ʕV�2"�}<�erj���붐�:�sڙ`�ͤ��7���U��ṁ.t�l��77R�� �
������<����E�~��n�je��kM!E{���Oj�N�?��=`�\���pl�Թ������X'MȘ���O���M��;��y�-�D�:k)�p:���)?���6�\�f�j�1u��w����bN��������f��f;9�����V+(��jxc�e�}��̛�r���P��Gh����{�BɱJr���-����*B�f���߉��a�i,s���T���X��}F�LV���*�r�ʹ���L%|�Y��i';�2�_��\���Q�z�M�t`�����T��:��ݡb�m��<�~��Wb�0D㞾S��Q���n����o��ģp2���#k���Y�N�^�� ~,�`K"�Ң8~a�| �Ǘ[%��sr��wΕ=�$���`ƩK�n����]׻���I� .�@M ���曝��O�h�j���m�3�nh�O�_�_3����� ��'�1�u𔭢�>u�^�Fz�WV���V�# 
�zStj�m}��%�Ƣ��AϢ��l��p5�2�b�~a��ҥ�pW��4��Ӯ�WyF֊Ey�J��yh�~y�q���W�����jMJvu�z]wY�x9_b����eD�1/]�G�a �뉆� (��Q�԰�����[7�X�@�T�'��R%Ϧv;��E�Am�P]�\��f-�'��^�ő9�L�*�O+�3>�����Yyk�0K7��D�Y��A*#H��8F�F�������]���36�V���Rc��;Sy.p�L�g{%�
�>�D,�����d��N��@Ark텓vϾ�
�s,u�U�-!��D�e�.4�;u �BZ��S@n���+�Є�ɇ�G����R�"u��D|��$^�~��,�����o�)��g'�ڌ��z� K�%�0:��-3J��^�.y���*$ ���8a?or�.\�$���T��{�}�X2���|�а��Ph�Qh�cIm�.�J8VʚîV��Ò�汝�k�)��<:�t8m��Q��u��?{`=�&6�����W�P����o��q��c9�t��Ok�=k�s��&��b�;w,�Է��^{pQ��к(��X���0|	|<Q�	%��0��J�K3_�0f�����׭��ћu{�'X�<8�g{���17w햫Q��^�C1j���ާ3Nte��[z�4�/�\@mʉ��E�`rI!c�fzq�uX�8�Nװ�[��@��8���9�vX-@>6U��39(�NL���1��H���x�y+p�����R�Hm�I1�X ��[g�>��BS�(���O�Ԝ�[4J��NO�G�W�"jש�9K����(��\��'5�ڡ�1�v�Am:�z`p�3�<�h���k�ۊ����Kct������
`Zk�����������KB�
˟�|�~ow�l0�]옺|C�Y(Ћ�gX�#ĢIA\�P��|e��ts/�oi�od�P[AQ)��Y[Ӗ�(�L@9 d稦��t/�ﳵ�s�2��t2�q'�#��w�)54"��[y\Ue�Um�$gC���6�-�>o��S��#[o��X�Z�A��l���q��#:>�1�r|6���z��3]<�kur?WJ&��f��(��IAXÿ�M�)����Mn`��`0��;�}Q	:W��#�cA�{\���d�FoB�擥8�����&���S�������Ɂ�w�r�]��O:���Cr�E2{�qQ����z�A�AJ���Ýj��F���z�`r=���2��z��RgR��[V���Q��U)39E�����"���?�cێ�7˽o�L(NL,�ڧ���4�0�XL:��E��UQ�媬aHq�"���yoK��FLÀ t�-����  '���$�L�� �lV�.3�o�)
۵Ә�n�'��/cN.���^�=ƭPoKB�!���}t0����1�+�p*E��y��Wp���4�^� _��;��@0cj�Z�'++B�kyv�;̘�R���m]�^E���,�f�@&��j���V���ĺV�Ǥ�")>��U%�u�]3j?ј'X[� ���;[�}�9�{����#�2���N	���,�4+[u�=��vn}N�{���9Ҝ��Jx����4%?9!��*_������� ��6��-r�O�ju��!�ڼ��|m`��O�"n[F���q�;�4�X+ߩ=�1t*m�H�S�"v��E�h@*(/�`'�M�l4�|/$�ox���g �NH�Eg]�*K�jz=9�#���0����'*4��&)�.'�a6q\��5�?OZ�ʨ��~��*dO �y��Ǿ~*�U���{*
;���ܠ���Ў>� C�|p}D&P;�c��.r�I�Y�����W��we` ���W�
�zV�Ƙ4�n�^�K�-�:i�2K?>÷.��_`�ZA�U�v&�(�|x瓽��J4�D�N/}�L4��e�.(�b�*�,����l�Ur�1�:�,u�?"�������e_����b�D�L�?�knL(�B>N���O�|�Op ��z�<��� ��u���0,Gjue���!�R�����-���q���+.�}�jxGwml�����Vt1��X
�����k�=2G�[F��wu�9����bXr֓��jXJ����"���_��B��A���]�-�w¡�F>-_  $k�O�>����ը{6[��˰g�[�9���o���,�G?�QD[tj�8��T~����b7�Ic������qx��w�_^j�4D�:�5f�2�r9E[�b���eP����ō[�WR:Y6�MuG792�;��=R&��)W��g�	��Ś=��6B�
�3��8맅t�
��_�S/ٟ�ߥ�����I=�j*Ģ��Ov���[m˪�����/\��n��n��p�/�����w��R����8;���e
��ꂈ�<��G�!~�[��U��R�������3��7��0�����4N����w���?Q�����}��^��?�Z����Ȕ�@C�b�.��A�:'��>��V�>-��t�D���q���
v�:�����~Q���P��'�W����+E�`�c@�����w���˗4�t�a	3�����L�MZ�ŝ�n 6��V��Y2!:E�Ω5�c�G@�lx��|�󐼈@�����ԃ/�k?���6p�9�L{�Zok���R������̏-mL���L�h��("XxO�r�T�F��*�O�D�>�,\�z�$T�vm����!5����F��$4F@��}��Qg)!Ok|�~���u���|r��!~0g��Qw��2��{ aX�w4�͵��n�C:v'<wM�[����~/�6������Y�>l��nԽ��Z�i4��х6&��GP�3��Z���ϵg!Y�`�U�Nv�ҽ/_,wP,��༆(F��6d��Sa�3�fe���7�壛r4���R�Ѩ��V�${��������?�Qp�Q�X�w�C7`!+��/����%�n�K>�71�Dg��`-�}Wi�md�ԛ��ӵ
��N�&�yq���B,Y�z=O�,Y��&����9g��FUp)�F�49ӡ*�����
������{���m� �6�Ӻ�'���6��ؒro��o��,�e��ܵM��[%���E�]�z�>����A��Oat�}�k�/^��u�)�ZD;��@�_z�51/񽩨��o09t`�O���*+���H#=r�P�Ш��
q�ޗ��kP"�75�����b���zӱ��'�k�I`L)*�L� ��+6�߰O�2��=��� �H'�BX��#i���&�z���\���A}�Nӽi�����ߎ��9��;J��@�Q�?W�[℗Y�jl�FJ��)Kh -�W���SR�y�O��p�/K��N�2��������F_�,c�		'�{T(KX����,m q^�9�!s5f�W.$�?K`?+�-�/�jc��b^)�	�U�*J��Pv}�ʙ�6��&4,��2�'V�F��wF��+�BuïL�o �q��7��.�׏n	�' �
��{�m�lOp�QH*��|T<���>K5���g��������Y�P�^'F'��z�0@m��ώ��$�*�*��� .a��1mӗ_�kB�
m�NGc)����zR������ͱ�K�O���>�f��%/����Q�R�(�~ɼ���� �be�c�L�%���7�&�1"��	x�i2��K��Ӝ������`m���E��W��WZ'���Jz�g��:j��ǅ�Q�X4ʿ�y&�ǰA���v���B