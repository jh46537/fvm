��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{�.���nQ��:�o]0��^���iY���%��N!�z|�5)-�f0��&l�B�aL?4�i4�g��L�����
#�T�p����û�\��L�(?��y(9�\m\<�ɧ���[]_�x�$h���c�`͝j�a/b�(ȏ��fz5FG�#f��;����":�\�~>:��5����-���-��q�z4ª�S$iG��Uj}�,��ˢp�p�]
ļ:hR�jN����ƶ�7��X�^��m9�(����Ё6N��G�	��h���%����R�9{�Č��%X���^�W�������IwL9NĬ"z��n�e����������f��5׫����x[�JC�`�'ͫQ�ᆳ��"��`C*�5|:)�w��>#1gU~!i���X1�~I:tX�Cfޙ�Hc����@o7����M7����4�h��w-ђc�ԏj0
��`/�SX-zz�V�����>�ii�	 ��i7����qP�S$o��eLot{�4Y��B��L�P��b:i"��ok�k� �䆕G������9��)����ѯ�!�"�Y���$�R�����b�Wi�^.d���aÀ�*#��V(tLP���}�s��*�Yy.K�����o8�o��1E�>#�'ŉ	7�g[�q-�Ϸ>w���v�&d�g��=���A��_�=�b+,��%C��gS=R8!��j�䢗�c]��V��-�-��7s��e�f *��i�yb���'Q�eDeD��|�J�Ws" [�x�]h�: ����ZC��1z6�Q��V��
�gRc����(1F#x~Ü&��BH����3�1�-^�=���`�%&�6��mw\�i�vE��|�W��*|���ھ}��ɇ�㰲L�뽯�T�'K���*܄m
�������cG[g��$$�@.GM��\E����r܀ ���O�b�9�Q)Lb���N�VA�q�P��:��X����GI�t�q(��0�úW�v��>���~.����TM���X��s��+�����c��p|t���Oʗɽ����e�i�4�S�Z�@}��bZ�-��<Zd�u׵G�Sk9�{����6��X�"f1�0�r�s�ql*_�Ϲ	W���;W�N��,u��O;b�'M^��)��,�7������g�w<�q�o�w��j*��F@�b�����1�$�)b�g�PzV<��k�Eq��_��ƮįR�e����a1��2�lHH����5��[��\a�nęv���D}f�D���=�f����{�����7�2�Bq��>���Evp��YF*o����tyc�>��ZP�P���r/Z�R����U���Nk!R6��!��Dȟm�9�1tW`���|"�
���G��,��3���^�XB�f�1O�|qf�7P��B����݌F��|aJ �����X_����0�9�Xyc�9&J�=]��: -S�Hwhin���a˧�)���A�"�Bh��\��¢�L2l�������-��^d�N'�D�Uo�bbs��������t���n���z�.���n�\<�Pd½��{�7/E9�_L��9�e�p�3�@�Z�R�� d�C�_��pP���=˶^�)������z��*~�w���-E�?��E��4�Ŕ4�	1���V	����m��_H��)Z!�"��2f3LbX7�&t0b����I:�U!~g� 9}�C�*�,�^T��]��)-�f�V�0*�l�OUΎE�M�g��1�ɽj�����Cܨ�Q�ŧ���"���ֿ�uɹZs����ʤ)OQod�ui����cN8��G�Pa�4���-i�'�b��\nt��i;C�Y⹽�6�U��	FڌAwXg��\�-{k"WQ��a��>m[N��5�!�اS�hS���^���t���S��hPӸH[|�1���/)[��,�I�0��+�������F���	�$�E���#bo�L.�z���]0�d�PB�ыL_!R#=sl�6[؈�[�|n�a��)�-"VM��C����g�@���ةzs�������8H>IA0�G���'���U�$,<	�	N�B!�#{o�A����&��ʠr��5� ]0���\��@�����@���p��C����x�.���[-�a`��m���`-d�4�L��f�r��Ԍ;B2��F�+��|�|'�k��B��h� h���>�Vah����@
m�#+o�����_����_z��H2��|��֑�ܨq�=���.�{����F~}d�[�Y' i.���f��i
��Y@��$we����������F!u{`�e��:�fm�ͬ �a~�<�j�i��+~�!T2�iĝI�ۡ��P�,��?��!l�R���8��}�[�wx�	�fT�Gl}C�#[�T�;���+��1��%���2�X:����\84���
��$?M2�0��3=�S�.��@7+u��3
��}���cY���1vաY����X��a���!�Ne*������]:�3 ���&����5��������:�E�������;=u���:�ag�v�C�Pm�M׿Y�fz�(E���Rʭ�4���m\�������WL=�s����#|���̱�^��|#�c$�
K%)�q2�-�٥�x�
N�$�v���{��2�	l�ܒ*w�w��}���?^49$9]������v�¨W�摆ɗ�wٷE�X]틡�`Ah��$�C��Eh��M:��QT��F��*����)�%\l�UW����%����o"�v�UIoP�O��;�^y��`�5�#����)� �\Y5 ��&c�1��<L-$�Ӗ�,�cVͳ����t
kd-����W_ ���� 3Lp�4�ڿQ�w<�.�1Ϟ���6��h��Eb|Xuz/�  ��;����q���/I	�t�� γ�f���>V���^p���?-g�T�T!c$�o���fz�d�˛ZXю>k�G�f)�����A��6��⯇f���S���� ��E�.9��۝����ʑ�O�=���%q��o���p2%�Ǳ�8��je��k�5��I#�L�����f4�
�6���@9$w:��CWl�;3?��9i��L?q��kF[X�!�"�UG+9z��cc=k �k�]A�%Ɓʤ�6�>�xO������AE����;���}�/^�ϻ�����	YS����oS3�BvĹ�T�<�#�a�t�������Ǖ�"尣?C{��F%/����@ݮk�?x=u��^���8�e�W�q��{gb�_b�t�R´Nb�<�y��.��	�p��1��ş��\����,O����K!s�acԙ,i�+�Y�Y��%_K��-�����:
`j����ڙ����?/|����ett��mh�]�]��y��	d�,
�^P]U��%���棕+��n��:^�-AА���}/�V����nyɷ�,�qƛ��;�<c[��&�,�
Y��O�u����Ը�6e;��*��0g������xGҞ��a9���]�[tn��"T]�{�<�W��-��<��W��N�M��m�l�
�����2�ܰ&�w����I�A�q"y�iay?'�ӗ�	5������D�>�p'=�D��"dܒY�)Ռ�-��l�Җ����Y��	�z���ܑ1[��PR`�I��m�q�D��$��Z�o ��Q�<�Ǉ�Î�}5�h���*)�����憎4��p=Y�r��5Ū9�}�1 ��&Ϣ*���ԑ�t��c���.�"��'u9k�܌3�m$;�Q�/6N&�������v�32�_���R���Gޣ���� ��u�GD�w|��_����������iC7�����r*}�_�#�a�A��2~�3�v6̖�j�UJ��q�r4j	j���I�l�^��J� �� ���Z����y����O��Q'�(2���xQF�m��a �1���^s�-�Dߟ��6��멑u�w�E.�0E�[���������t;�
r@E�����IPG���a%���&Ϣʯ��_�ՙ�H'|&V�5�v@1;�'T�dp�c�hb�E��������Y˕l�!R���
tS����ٰZ��[��7�zn�͘2���m�6U�����YG_�PfVG'Nz�a����Qk�ܜ�j�q�3��ϼc��ڋhP��������k?���d\���a�I�1�ͧJE+Lvix�h�г���aQ�']��o�
P5���}�p �p�����'��<b� �6�y�G���3��7���md�K&�e�g]:��*��Z�\fU����dI�.Ò�y��<,	rf�.|�1����,��{ٚ�<�t���b�F�������!ý�Hv�)�WL���s��P1臣3B$��sPsH��g$+��>������03E鯲���j���ޱa�,�zTPz�(�F<a����O��]-���x5W�������n}�c#�|���{SD�ܞҞ'��[�؏�M�o�j��H݅�\�ϲ^R�c��z���<3�q�x��^��i*a;��5�d���m/erM��"ᚲ�����&��[k�݃����Mv��ĀE$�u�DO"�x����;�K  J(�G�9��_�X��>�%�Ȃy�ϽXX�o�s�6�N�E�aE�:- H��S�VR���9==@j"�]�� ��7:�×�$R�L����l���`=q�ZI| �^@57YM�v-o�%�F��yqYq�#�,.6�(w�`
��/���u���Wb�u��Î���j6��y-�	A�C}!�I�z��d{d<X�
��7��b��`�� �̔�Q>�'��#G�����|��ӵ�����\ɖ���KIH�M9�c^�Od/΂ƍ=�+H���jY����
��s3�5�qhR�+}��>6S�oBl?�t�OB�Y�~�iYF�Q;�}��1���~���g'u7F�FȀV�B�i�A�Tɡ�64غdAq�8sH�L��רu�of��&zS�������������v&�hb �P�f�Gg�*d�Ls}�t�����*gemwh0��i|���G���g:j;՜�	[��f�d�@D�r4È�/5��\�/������