��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�`��L�o��<�T��u_T2�MA�J���?��P�p��z˦|J�Y&�׈��D����"�d��i޶�8uw���Ί)42<-f��|�*�P9u�a���Nͱ'%�?�8��o��K|A�H`8��G�V�30@
��%�$��i,�
9�y�N
�r<3�x*�x�X�R���Jx��E{�����QAZ�tƉ��;·�ʄ�R�E�#6'�.�g1��\FXҧ�M-�Q����@N ��~������ㄭ�ޓ�/,*�&���5�coȁ�<�s�Ҍ�7>fT�5]�Y�˓|A��^:��S�n�
�Q��D��g��j��/v(�dK�y���Ļ�,���<|2UR��~�a�16�r��j�MZ�w���}�.��f,�Kyx��u�_W2�>�� �=_;�!��]!%w?5�^$��c�"Z�z�{t��Ё5v�ԙ��N��7ёy|m�Xq���k�I��t��%��C�+�\����Jl���Y��W�Y�97xU�Z��V�,��ax+N�P��D�U#B�M�q{5~�+�F���`!Vm�ճ��;Q�_�z�����q�5��M�@� �;�[��l93m�F*��`�y+��?
��U�����}��p�E���Y��1$`��8��m,�ib<-gL?�
a��?r��Y��ǿ|!��H��WSr?�@�c�w�!�o��;85�� &�2h2��&��tWq6D��_���ϑ9U�,���G֡���(��u�]��Z�%J�����m�k��Zs��|ɁB]�K��ɦL�DAlCW�H����2y��c����!q�fM\M�I���(� ��@�KNī�gNh�F���<�;��I��E��	�P�l�T�)��mwz�Q��\�iU&��+��T�k��%�ӛ���]Z�����/��U���0����=�f&1�x�q'��_v�>R���d�}�\� "5�l؜{�7��h��Ҩ�>�)���C���W2��S\�p����b@�	����`W��Ӈ��F:�g��z�T�7GN�O2�e�ƹ#�`W��Ž�r��#��e����j�����&n�`�����![�[�O}���T"����L�
H�����.G2�X�X�N�H��P�f����bz���+c�h3P9����ֶo�
�}{�?D���#�)D-���Fd�x��X��������9~�EH���|1m���lw=����zZ+r�30^U�!�����&�2�c�0bL�\+�|�ThǄI�>�vk�a|�Rr����Ѥ9�� ����䐶cW����TTZ�묏�;�� !*"���fPZ�~'S=���>W]-n.�>�>�����oH/��,���$���Q ���-�۽�IG��*"��j��5t��p�,�H;��i�s夔}�ۀI��\m��1��8x�'�t���s&�Q���hx����Ό�@���m���ƹ�٫�1���_r)�9�):L.���h+��qҦؼ.R�Z��j��d�^������Y���p=JFP	�}N/���N
�`;J�큲�dM�ˆ���_!�t�+�2���_��j^���u5�ehhv j,�B���6���m[�l�Ǆ8O����pbI����hoQ��dxŏ������y�.�[��Y�Y"d%������k�?d�a�O$����դ����`�`��U�f��ܹ
(�/���-�lt��e$A��|���Yq/&ɨ A]�]�f����������!�<�X �3�ד�m7`�xQB pv�F#_���	F�r9�M+�G�O�7X�gJC��#Ivp&A6k��/[ɳ���N�"��¦���4�DTm�D�J��^\�CfhU^>)�t���"V]kw|v�k`\7��f�3�H�!�;�d�V���!K����8����޺�B��Czi���f��Q/��h�����0:�rT�b#��i�-�ɝWgPS��R�@��&���3.I�c��<�/Al�@,r��8��9��[L��"
�;�@��iy��_���>�����8�i\ֵ��}A�w��x�Md�SY!�Wp&6���	@�����w`'��|x��&��h�}������ggFc�$�M��XɟU3)}�n˪g#�$��Q�c$[
�<@�