��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0�����
����'a���en�,�=y��~{��i�#�sS�Z�àx�WW�Bg������𓇴r�b�ex�Wv�c���V[�4+9o]��\�S�������_���]U��J��]2c���L��<e�@�&���jX�3r|~�SrOa�{NR^����y�R�ΏD�|����m�'�m@�q��S��Ƣ,(�jݎ�4��>X���w�j2�)M��&�wU�=�a�;�k����K���b���ʎ�\������E�\��,D�`�������A\]��J�o�A�����^�.�c�mC5�h�9����N�
�.�C�!�V ˘�٬.#�]�	ޔ.�⏩� j4pTMt��U�uW#�����3��ɐAw����/5���C�اDt�����e���#�h�e�W��QyG	��,ct��{6k-���w�Y&=pK]kS�g7�̝WJ� �
�Y�X�K���L �n��ӡoQU�Iy���r���o2k�aYDx���v~WX������+��xe|F\u�R��0?ked�1G���U��'i��Q8{���=X��c�H����Մ�t>����Q*���/̗����*$�
�e��N��@���p�[����J$+b��6W�T\�oq���+ �0��m��6���Ǎ6Z�Ss٦W��*�C�з��W�����n�4�� /�� ?ؓ��9���@K�*._ba;w���NTK�����\�rf�C����]���56A���N?d��_H�CĬI̊[v����~�Gi���IŨ���3c�E(b���K�N�O�rq޴�ɤV� Je"
��_�m¿�tt�M����r�@9*�}�e5�U���Ow����;k���Q�!��]_3�N��L�b��Q:�#�0>�$��Hd��^��'yT4�Cs䘋�r��5�����zg�pX2slִe���(��r�P����o8�b�&ȦX4�:4�0��3S�s�9hb�$S����
ھx�[���DwɄ׻
 ��y�$A30�" �Go}�ά��f&	K#OU��ߗp�@/qkP�Jv����Ǳ������cykb7l�KڈK��/>#:��K���WG��tT*�R���Q�I�r�Ww�byK��j�lW(����"2��Y�p�W�n�|�U�z�կ�$��
A�v�d�;ۇ�,\`�ġ�Bu 士|lz��-��]暦��}>�=�ip�`�7�R[�T�6���AEG�W][�Xې�y�����"D[��q�j����τr,e�6-O�'�F� ��Q��(�Aw�F�Q뫼J(<�aV6���b��1.�R���<*�{�*���J�f��t�!)/1mա����H����U>5d!a8�����;��궖<12*zU��\���y��6�Ʋ�y�V�����*�9Ɏ�HR�z+)��A �;E��ҷ�'雛.x|n�x�\|�����Q�Ws��OA\b��22%(��WF	�r��a|�U5!�c�xN��Fۯ��Y�L�Z΀�?��1R��q|1�9�n���iuC�k��I?K u��}M�Qo�"Z�ˇ����$
�P�����ӵ��=n�fu�{2��	`�l#0�������8�V�=�ʱσ�Jy	�A!�x�1�B�n��1
Lzh�Q�=
@r�#�9�Z�x�n�e���9V�٠:�p�\O�HZ#��n���R�c?P'U�\ݷ?f���c�(�8�� �����U�9�>��0�h�X-}��<�x�<��P���X����A�{OǅVT-	=�����4���B�s��tZD�w���d�(˸��3;�h��0�8��6��eI�����X^U��D]��¯2�jMA6y�@��@�K2�m[C	N9�ڜv]����K=���f/���\!>n\q��4DchI��^¡�ƌZt<�ء�+���	�R��q�\1��~g�z�P�]���m�0P��#�Rp�+9���zn/(��G?�^�vC9��uv\Mc}�;��9	\u���Hr���c��Yo?��s*�k� ф@	z�{Tn�p�f�d6LI��W8�%'S���ӟ�h��`I�@p�v��H���ʀ��`��ʆQ�i����k�F��,9>�9�� �ur<hW�,�J�!�f��E��ӡ�Oռ/��}�'��?U-�a����sԲt�j��A�
��݈r1/�<	�����X>����[��WΙ+\��
�ZDN�f�iwE���{��I�a0���``=#��d!\�V���5M�:�\+(7�j��}�*1P<�^�[�����F3,1d2�N��Y���J�!N7�x���N{!�B�F�]�<�\�2���ӎ[	�Ju)dj��[q"�N��)S�!�f|�:;B����8�ka��0�� �d�	�,�,��L�`~���S�v�����"J"5�@���>�m���2��� �*�l��I��d����g�ߝ(K��l_������Ŝ!���O�GS�p���`>(��S��O��o]lk���>��ԏ�f�(v�����ah1��mJg��5x��#�-]u����+�:��M�\�t�o�ik0+���C� ��!R3+��O8���:Ԧ��~ŏ�tCδ>y,�mm!i"��)���\���V��
��(���-�I��Ep*��~Y>F}���T�$��R3�}=o�ѧ`!�||}���d�����p\�E��]w4�
�A������57!�Ѡ�|5��\�����q������|�n�p��P�+v��Ī�|���5�פPѠt5��o�8� j�=1\Oil��s��L�xlQ��3�v�tew_1
������!s5r�:H���S�v�aj��|�u
r��u,':plK'��d�9қ1�n��U���i3Q��Z�U�%8�S�zO/D�'��%?����yə��?��Ζls`xI�c��_R��X�vnS�A�T2���	�|��<�K��,��}��֞oG���P=]=X�y�=��[�w����a���;J�cR�]c�)�k���o��
�E�m��U�tض��X�`�ݰ����~N�BfN����ֵ%�ďc'[����upۇ�US'�}��V(2ڙ��S�	���E�j{�|��s��
�A�c������k��PV��At\���B�D��Y���#w׬�q�;J#��r�P��ou6 g�V���\�G	�}"��`��*F��A�W;�a��ˠ��;{�B�L����@��V5*�m��Obe�db5�ZNBsa3P_@	7��M�`�d�:{t���&[1l|�������*w }�Ow'��J�"�p��B6�k�Y���fW����{�q���XI�����і�
l'�"�9a�C�M�E�7�V�� �ku��S���Y(w����9��f
�UH�(
���6x������U�d9.��B�u������X�{.G�i�Q�H5�P��D
6i]���y�q�˹l�lA,�mt������ʁFdZ����\ҡk0�y�}[���k/�=|蜌��00�2Zp�4��jeW��4��j+$ ���s=Mkߜ_������}U]>�����J�v���8�C`�"����� ܚJ_�C�:fb=uz�k���[$}��A��u�n-#�'��c/�n.ױF;��:|8����'ˏ�ȋ��c��}ڜ�|�����\�C����)�~���6A�	���Z���HǲcBYt�#I��Ե[gS0�h�<����Xu*��������^�Y�Y3ڼR��ji�����>�U¶!�������zQ{�mn�.���\:�q���3n<�n���Ytُ��d�:�ՇM��4iP/2����\�ؗ��ܼ˴��(�B�� 4�(�^�F�/w��X�)���8�-�j�q�7Q�{��C_0Xu_*.�i��e)��o�`���[1<O!�02��hu��%�)$��ۙ~j�uC?��k��!yo�A�R��D�e�D������9��������@���¶�[��4���F�M���aLeqh3%l��i�\��pT,����@K��RP\}�_�3�bΡ����'�V�{ ����x,��޵��J�A��jU��ߞo�ۿ�jL�=�������N�ß���9V�[ Uq�'ߌk�bt����
c!h�	�U�I����3����RH�gs�Wl*����?�{�L@�ܠ�e��А��yi;{�=z`���(�ҷ�r���!2�i��[X�Y��0����M�ݡ<ӪUlS�ÈG�-T�鹫^����k��Ѱ��j(5Ǝ����~�2M��yjm�7&��J��C���`x��6���u��hUZ;�t�BT����<>��=��;T�F�.��
ql��҅D�s����.�z���Q,7��FXd}k&U���r������3��