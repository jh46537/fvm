��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����,��f9t���3>��Ձ�A�7M ��uj��M�0��{�ơ�Wa=Kg��!洭D�2�&�6����2�����X܋��x� ����G1���w�S��3�C�1�9��1+CH�<3�vwN��F�T�\#[�'I���ҒO*K��V�6�k%���D��Sn�&$Y�au��Q�/���OO .�XS}���9��k,[=0�hj��V���w��:g�!,;�(���1��+�\�dn�����W#�5"T�\>��s�b�֜S��� �5�b�s3�T}�t>��7����\�[e���("0O�2C���qO�l��G?�9<�6���w���X]u���yd�W2~�h��`�7�j���s���vFWc@3:nsS�"�/3��r�.��w|�I�h��{̽���rB<���\3'��e#,�=Kl�۴�[<[o���� ���=ѽu"���g��\T=�{�\ ׭��^ֽ���D)�n�6���������IZ�
K���J�?6ɝ8K�M�"_Wn�����tN]}̀	�Uꤳ �*g��x;�.l�G7+���Dx��
QWQ��d3c��
�H��XO��f����0\v*:c0�m��d#��r}����DQ�Ʃ���s����H�-�$M�X�V�r����=h��f�s�.�����_V�nB7�W��Au%�4���������}���5+��;���Dd��!e�螺��<@X�boxkӰ5�
���z�QGF�ȔnG��:	��,�c�|��Q~l�'��>�{㠉X&�%�������F��B�+��F!Mݧ������Y��7���6��C\/M����`?_k�ƙS4B�˴�>�� ��exq!Rq�.�hj�O5V�yhc��GS%�7�ߘ�ٽu��R-Tf>��\� �ܪ�J�pz'�B'�ۊ��2�r-���č@�iÓjaB*��d���������++���3W�)~;bS��A�6���m���f�����2�& AT�l�lXD���̀EE��<[�0l�	��)��e��O�o��ӵ��~��/
}x}Q\��,f�kb8�	�?I�Jtౕ�������\���%�ҠxT�L�e%}Ǧu�D7���v��kfڅZ���'�����U<�EE���p����lAHO�I�`�+��lj)57�.���x�L��#[�F^P�C����K٨G�K���X!�z���W�+^ܑp>^��x'��DP~���I"�^�*Bt�����C�!�	u@��~�������7��1�k�|��XLl�&�t4<ATiݪ�~>4>5p��2D�[�j����T�V�?�Q�' ��*��~L�����)�����Po��F�Yq_�=#�%ѧ�J��d��W�n�'!��1��[J����ę�v�T��&�Khǈ�� �S�5�띄v���$5���Z��;S;B�s��wg�BЁ�H�G�)��E�s�^U6�i���hh\�>s���<�fG��Y�0�*�;YQ�a���D�/����uM1ܢ�-�{2�pS�In�=�/����0��|P��JRܽ��Ƭ07؀���[0,|���A�s���]��x�|�� <��AY�т�h�ݓDͧn��7��u�ԙ␫�^k� ��V��*����4҅��p��rb�x��=�qC>[u'{�=�Qqn�"�N���"G���S�G��^��~����� )8��zjnk�=����0T6c뷄�#U����OX���US8�yV),�������?�Y΅Mֶh�r#��R�l���h��3����ln���aj{���%M�?\P]LX����-
"�)���<Z�� ��v����T��Z��A�=��K��~���=�� R_���M�C��6q���Q�]*6T'mt'dj���p@�(�B�l�G�4�uڕ���"�ך=�9�N�+Y��_@�O�,K�{oS���G����Iu�O~���Z�`p
b`��[�H��^�{M�4�	��f4y�AK�z.�헾z��o�i�a��85!o�B�L�8K�AD!Ar�I����ٹI̢K`�vcP���2��^0����#��Yyi*�g�����JC�8��6����])xI��9$ɺ���,�9�R�w�}���o.`�0r�~\Y~�9�R��No"ƥZ|iC?����׎���J����Dl1ZV0&��/�[�K�fZEp2�f�k�X�9�lu`�$�a0!e�$���"�r�q��҅�7ʵ�ZG#rS�a6آ��}��� 8$�`]���Id��S�WKcv��ߙYf^����7z�� �P�-��8k���-��QV�8��x?(f�xΈU$b�{�W\c�t8��]`�}��=�|�雰lx̀P{O9E�ZCm�B�($@��$�xv�
�<}��y袆}�W#�����:��.D�Ɯ�[����ԇ5+:U��~c�-���[M��9��-��s��~�����\oן�m���C��ʲ�_5�{_�i,�����oz=Z@F�S#K/I����Ψ%^��⡎;�4��M�S���(�eYA�H����nDm���e�#`�v�
��^���h����Ƴs_��x`�-���؞��)æD_(�<k�E��������v����`j�ʘ��<�WO��&E����q�'u��8|!ZwlK������n�=_��/�5�d��bî�J�R�L�� ��$[Zt�C�(;, '�/���Z�����<���?�ݺ��P_��(�J ��{��ĩŜ��:���k�^�.'�
��+g���ɩ��&���, �\��军��uRL�L��R�5��K;oǩ�(�/4����y�����h!a�)P-Ef��r�\��/�6JXQ_5K�5;X}�	M ���"ne��BS��ژ����+����_�{Q�	���OtG��}:��)���}�偠F|��ES�
o�X6�;hÊ��k!�w|3^�%"���z�ò�`
�������U���m!+��3��R���%�y:=6�O����t��;t��Xq0 �Z�w�x��$�KG��t��n���(�0y���w��ᬚ�#k���xlB�]@O����e�ÃO������BR�ñ�K�r�_G&c3�.�S?�]�ن~�լ���l��40�b3L�6�N�b�9��̓<�'��[�#D�k��ij��eu2/��a�	�K�ȋ������.�{�����N���<LfvJ��W���^U�W ����f�a#̧ 岟_�?�<��o$ě*C�￫����2�1�,�r�~8�3�2ai.��nR`/�'��s��X�4`��=�(&��7f�UЎ�L��{��VKæ�K�J�#�J�I|)�ϝ>����_ؤ�9C~jUx�� ����)�n��d�]�fV��!���d`#<��N�)'�f��&R����ʓ�9���s+��m�&��ʏ�b^�z#�)�7 ?�Zm=�B����o��ƾ����>7����~e� xnƛ�5T̖�D����X��҃)G�N� �bJ����(�<�j쌢C��빰�C5�r�u�J�� �5���j+y/*0,�G1$�(��pl�^M=�c���?5 jxy� +�ྈ�!�}R��%�=����*�.�FjԒ	�nL)�>S9�\�q)HG�7��E���o�GA�s9��}@�!��C�/������Db��e���N�%^r����A���a8_h�<2\3vm���d%�u����d���mꥇ�  �;~����8�ګ�����L*'����gdf-���K�7��)IS��@��i�/+���z��R��s�6zE���I���O± _��%̼_K����E�)��IJ������:d�'iW�����a�l�u��̤[ṅ�j�LD[G��g�H�_������;ﺜ\�(e�D:l�20<iMq=��6�n^w: ;Y`NH�r�g��Q�Ĉ�ӕes?UK��e��D �Д�������(#l��l���|��3���"m��;��o��h�T)��L��G�w�]��5�!ֵk?_'�/ɤV�j���P�a��Xr�НfDEY��Z�^z�|MsF{��
}O�i� T��a2Ì#�Q��8FFVѬW��Y����R�w0b� k���9�����	Y�����Mm�o�����$���=m1������ϴ d=0v{��]c4-�� f+]�F�V�`sj
l�{��?ܟnå�u�W�5O���Qg��kN��|F�����H�N��o�=���?^/h,r�0PJQ[����n*�p+oQj�����1�"��p�g�oBi��� ���%,�hܞp�.ղ��8*�A�gp���M5%({��c�m�0�-ф�>~�FO)M����5�ƸDu��N.��oFc�A�E_4Y��+<�� ���,ۄ�T�0��!�SD�[����-�&��Kz?����y]��_�f�I2+��DġW|=�7�R�Z��l���׺��{��/���bsÞ4l�o����11�	<����.@�a$-���yv��&��O�����3:2;��Zj��4�����Y��
V�܊���m���6�Z9��^G�f"vN�ve:�P�"�h��ɜ{G���Q�g'SP�e|�]�h�Ly��AX9�z�]ez47��1��$ؑ�>�m��Sə�(>��e�m&��H� G��½l��)�YN��?�g*d���Ԕ�%��'���/�v�/���@7qe�qI�+������S��	!¤v�s5K��9:����1�c_|Y�ԟn:^�&>y k�F�[�`�ȣEr�Z�t��CM���x�~�_A�-�*��"�t��߹�MkA�)�Z��m�E�Z��%��ї�R��F4���T�#c�됷R)u�0 t���Y3�i
fPT9�ɗ)�����Y8J]����vI2��ͦ��1�xlw=��ײ&MVa�@;�SXu��]����`���3���~�����Nܜ�Y��\����%����8Hv$1J��ƭ�PgzW�*T�`�9�^�}ۿ�A�	�L��,+ͣf��1���d8����߉��ӓ����ܯ�S�
h[����6yt�c����x��'~~��6*����"?�Wln�c��ă-r��aO�C�����&�>ٻ ΍1B5��;� 8b�,	����o�G;���$?l�a�@S�g[�d%~"s��lދDz���t�<ᄺ!�qřc��)S*��Ne�;�����2�Rnč��	�?�6g@����]c��twԋ�ʓԶΐ�C��j�as;(��@p�� f�X�/P&�t\�1�Bê�1��٢P ��)�ai�j0׳���Y�'��Ĩ��P�Q�n�m0�Q���rT��f���|�j��z)�@�]�W��C��Ąl��T��[�3i�7��~}J�dv�'�|��{�(-G�
�HoKX"�f���Rh_u�,)�D��<т�ǻ^�E]$����Xz��ǉ�)�����KY*��7�����ކH$�$xr �'$C����E�~����૒�F
mݓ�w~"Ԇ(U��C|wc���8��~�`���$*�C�_d�uR���Q�%BH(��e���ud���Ί'�1���*�P
ܓR�M��9B�i���F!�Gih����z��$�Sj�3��q�m�֠���2�:%�ڒb'	�|����;"�7����8}g�]շ��:��A6�vq���y� ��z��3PlcN����Rr�*���S��Y.����o�~�j�o-=/��i�""�ˉL-��u�"�<o��$6��b(P��×�6�}�E:�yg=���*7�j�R|6�Vt��].��XI��2ٷMV�刑�j����t�C���z���}� �Eպ�I?~�����4�E��Պ�m��4�=���Ϡ���u�+e����&>��		4��Xo��hJ&���(^}��9�7�� �LG��n�U�e^�����V���cD��E��ݏ4�X �**P�9Z�Y=����öWG�c�1�ZSWPv�����^���v�l��K
<�a����I+�ضBqǄ߮�`�*�ŵj�Zpd�D�汧^�[�g�4Š�*���^܂���'�l��S4�4��rfR�$bS�RC����cN:�h@�N
4�u��1.�~*�ov�]��>Tv�S�ٓГ�@��T�*��m���:�U��"���D�F��ul<(�Ҩ��sԛm�Gg�D;���\(������o9:�e��IgD9����;Phqz�E�E#}�г���`�Q��*x�,��J6�C�P�6�0좌��Q�0=�����2T�6 >�6����B�܇Uo��E� �h�\�~&f�>o)���У^GJ�uiݵB8����U����Y�ROn�,N���J����Eg_L�p)91q/mA�g�K%h4��O�L׭�����"�������ç\�'��]�.c7�h��p�bLI5���.i��i//2R�`��}�p��v�Gx�8V"ߕ1�H�{L��@��-�:�l�'�^v�9����!�&�N�@�Ҭ��+�@	�Pnz|�%;�h��ޚ�WaٯRhS!�� �{e6oY���nd�l�o�f+'�k�u�(Z� %t�3��V'+���������6���WP��[B�/u�4��ʤ�o�R��o�7�oNm��r�	g9��2]��F�v�Eyl�/	�d�6Y��d���6��M����o�-���z�jG0?j�/�!x��3�q��O �~�N��a�I\⠳�H�w���5�Vu���f��6g��+9�Sȹ9.������6K%�\��O�h���x�"�+�*�`�5	T�ccxK����`l��-�pH߳NTx�ti��o�\~Dt2WMR�d��|�	�ƁC8��K��eu�=҆͐�;a6��߄,zbX�ϐ:���}'���"�*�&�z�c�=���m�$j���ri���-u�{p9ei�ʬ�ӘJ��&3��Zݍ�Z� ?8p�m��g��3%�<�z3�Gs�RQH����������Q��U��������AKp�+��d��ŭ=n�W�RBG���2��P��	S� ��M�b�S��PI���i�#/��#d.#��w�V�;?���ca������hrċs����FC5P.�;�-��襤��9���J0!�?�w��:}��U�3�e�aj���-��]�]U�ʰ��ͻc/�/���.�I����t�<=����C���C���MSa�|�Aޘ(T�����X����~�w��%b��7%s�\���Zq=d���J�$[�`n���C6��(�c3y�7�ʻ��g�훧��i��d'����[}� �;��r2�-�7W���\8)�)7~*��VRߪ�����.�Ԗ�;��W�C�������K��3�k�&�'ːV3�gg�Ǯ�1�q�I�v�(����4� ��-� ��8����E~��&�5�c$K(`��v�\�������0�9�t{����-�rXDl&��̦�?���:�d�w�d�QI1g>�T11s�����d���23�UM�N�I���v!�����f��ҝ��~���p���h*��_��/�ި0ꇲ�KD���6x�$BA����]�4Il*��x�	s�����يՔ��V`
$���AG52ධ#sZ������va���i�'+���ta�F�h��#'���ŏ���j$�,p�&p9$MjR�e�}�x<������*�^�_4���}�ǁ��~A4�՚�Q�/���[Xl�'(��ϊ�C?��������u����{�"ܳ0H@�4����"���]����s�._���U(�l�O�����QO
٠190"�,k�p���J�c�Tī�p��h��F�t�ݗ�&81"ŧ�l�|'��p�Bl�;�j񚺢gȏ�0�+�Y�Up.��_����X�!=e4��s5 �wxt�Л])]��Q���_ɔZz8�N�[���L�>�����T�9Y�'��%I1�l�ez����ŏK��{��y]L�,�7w�Z���R�S�=�9��hQ�|`�B�Ԟ��qw����;nQ>"l'����^'V�'|���/}]�s��5�kz��P����q[p�����%�!�&�3�c�q�89k����Ϡ���	Tŧ$�怲º�d��⇓�:��d �R�A�ZV�Z���jY�"=<�9QHQ4�L�����g�˯}�~%���{�c�O�k6ݖ��Uh����[^r�k����\K;f�����.����Yl���$?&��K�ȼ4w Ez��MLa�Tv� үIǐY:�b�o˽�s�(:�Um�%�8gQ��<��.��q�ttc_9�$JK�2������M��\C���]5�HE�JM��,�÷߬�tM��@���wРq;�pA�c��7�<��n!��:I��?\Pj%�,J�E`��gT��վ=O�^�՗=ʂq,�f[�zI1���SgՋ�[�Z��w�O5�0=<�Ŷ��Һ-���fn��w�R��pr�VMPŬ�N��R�-��ɺ����H8^�$'���e���Ɨb#)�04�|VZ��րN�ʚƲ�f,�d������'b��7�-!�~��?U��	�B��b*���+�y�
�������gTB�瓐���OS����C+�sŴ�z�4]M�Y���mB\9�-���KO*�zIUТm�J���uSPQ\���0$���س6[p��0�r��[8�5|�z��&�T�ٚ.�<���UQ�\-x�	� �� Ţ@��='LiAU�~b���|�w�짶�2)+	�	��~h�u�s(��P� ��@��Qj `y%CA�
�v��1yzT��\�,Pm�W�;�oL�Y�6�	!�mk�P�6Ml�7��Q5�n��M����=��=��9�_������W�]H���'���m�i�� n��i��g�+OSIKW�N���kB�\)Ҝ��h��H=.��a�� �Ч��q|�"��Hi����y��e������e7����m����۞Y��dt@���A+�����%��1��|��ٵp��5ȥ�Y���ŧ�<C@n���5�		��s'�����p�w^�/�Ї���Q;�n������
�X���rs��%�Q1v�驔?�)8���ke����h��I�ʩ�zfJ��bq�>(E�N�8ߒ%�-� r�Ǫ%�|ͷ`�mn�>709P�1*�<�C*�/JTz���Ȭ��S�����1zQG5^��]�YDw�z�.J�TmV��4�"
!a�����4�1V)��f-ɜ]Kk���&W�E�������K8���1qv�6�g�����_	W��V���`�"w��/��t�
��n�� L7�'��������;��цg�	�mkIk���$l�u�eu�׬ȁL3��)�j��.���L�fj�������!m�rXɬH�k2T��
G��m���z�+:���w���b�����-�O�f.�A��8$��fQP{����""�i"Ď2�FW��vy�Kt#<>7��pt����|G�¹�>b�o��%U��۠w&o���w$q�J����KJ�����gRB\]F������$녬6����%��zTx����A�A]Z���r�X�1����D7����?
kb����R�\���Y��)�!��w`�̚S�!1�������)�a�{%���?�%���䎀���:��	K�^5�_C ��p���L�C|= �������Pb-���ϙ?�'u���hO�3b"�x����ϭT_�B����uB�R\�4D�a��0vFE�V���9�j)�����w��\�k)�\z��+lQe����t��eW{�IJ���`Nծb����p���K�70,�$`&�;�Ƣ#��(�.���g�\�KI��P[�|�4>b���x�G���{');�\LC�ի~�`H���f����bT���s�R�������{�F� Z�](�i����(�=�h�S�����qt	�^
���]Vk^ɺ�uv!K&�������j������t?��u��zJ[S�k��w��B����CCy:�$��"_HB��Ck�7�KO�Rw�6��T�� nYյ�X|P����B�j��
�Ȗ�\F�D��V���U���H;�(�!��t�%�/9�����K�x�L�P?�����0{:��ހ�0���pJ1m?;��eDI�	�}�K�hN\�.��$���7<�^5�%�q] 2�_Mܠ�j�+J~-��F��0��2C�NgRY$06�8������%*<!��̴�v��ܸ6\�T�&�k8���_,ۓ��_r:�eu�6�8�p�刬���e�*�}�8�	B1����ѫ�d�S�	�������9Hz`5��i��[ H=k�w��$ѐ�&m�3�^�|��ˈ��NpD� i���R֕�ox�$� ��یRms.���HAj?	�V.hT�E��c3Lo�u�	�E#�3m	�&k:�-G5<��S��\P���½�I{��9�"�Z������ָA�F����
�uw�X��e,:n���Z�p�`�x�2X\�Ө?=���KXB-e�dbH��M2��>�縞���t΋!u���lYO� PV�����Ӄd"3�K�i
U�w�ܺ��H����'K�\ǣ�`��E�1�߽��)��mg�ALs5hXU���I�)s�e2(Ml�>�!�	�=� #-�ά|�{zz�=�-�����@x�i,@��g3�?��
C���*�sbh�l#:Z�R�˧�k�%{e1��r�)(����r�h��@��g��[17���<�͠X^�#r�"�.�yBѲ	GND�k��`b�T�4�:̀�����F�fL��G\�̀�&
i~�X�/8��~���w�5G�En����tA���hϜ������f2~F�7#P7T�h5 N�"�~R�(2_�l���WՂ�"��1�k)�?W4�@��	}I�{�TE�r,�qь���V'^��Q�Ւ�i3P
�҅V���5��.�B�,i8k�E�+mw�1�-��� z�ԧ��07u��"�AJ���{l�Gb�(=NZѼ��B9_#f\T�O@��\7)E��L6�#Rͪ���k*�T�˹�vxν��(�.�	z��[�.0.�9��s�X�8�W	�K����΀�>��s����XS�u=� ��1A=�g�����`�/@�{9�P�@�YV��͹���	@���ѳ���Փյ"��o��Y9���*�`a��kB���A�^�s������)�z���#Ć�ח! Ҿ!��˵L�ӵ�ٞ�E�a�� Xd���n䏱86�!w�"���i����?��Qk�&T'�y�*C^fŬJ���$�{�47�l�ɉ�H���M�x��Y<�YRĖY1�<�L�:UhwH�\�S�gb��\���y˚����z<P��&�F�I$Sk��+�|�� �W��k'6E�� ��h(� �,5KQ���VT1�+V�����5��S���FJ lh�pH=��z���/'A?hMYce���
m� Hc��訽 )�Fp��-rԹF�j���sKE�ȃ�V����?P�rD������v#ۨQ�yb�ƀ0��R?��~�0�:F����6������p��b�w"P%w�O�]���\������h��>�ek�H�.(��5�,��G����i�eR=�q;@X�3��{|K��y��
l73;�z�y�>�ӷN6��)|���&Uڴ��F+��\�y6������M�,��A�>�|��U<����ۉq*k�����F��>�d�W���0Ƚ,ԟG����e��7�`S=�V�|X����FL��1��OL�����fu���S�\���i�����q��Ŀ�X}۠��ܿk�SC�*K�5c=����K�4W���I�͌�'��5ک�KqgN�0��R<��>�B2��*��8������;IAHFF?������W�T�L�R o��W��������߿bIx KH�n�1�=�B����2�W|��*��������͊k�r*X30��G�P��%+;����9���Exn��J\����N��}K+XQF5T|��I�S-���G����m�Z�>�t���ZՍ�:�t��$�v$A�0�v��>��2J���|��O���Yѹ�W�Q���g���h����ƪ��&�s��R.���_�]��@dʁ+6�E��u���ܩ0��͛'� 	Z�^'m��Aہ3�g����8����D���8>��ռM�J��@#�N� ��DJ��X{>ܖ� �V����p=0� �w���r��S�u1EضGD��u�u�S�/�tס�����F�Gn���������V��"�f�6�nq$���_i2\"e�}�D�� W��r�L���&մj�i�(��\�~-���o����*H�=:��x�GQ"�cA�^nGq�c�t���ݸ�a$���X���[<� �;�?Y�+��Y;�*X�ՠ=��Oq
��y@ɥ�Z�CLN���Y0��~P���+�,��Zq�W5��k�t�����Xd�U�-*=�P���y�@�ۀC¹��s��dz)rF�3�x��.y�߇�1� ���$ƿv�d�e���Iv�6#����Ctϩ1Yf�|��H�1�D�G�ɭbd�Z����{x�L�����Ea�����hL��M��v�0����CV�W}�yFJ �i������}��|���?��ʚ�v��Ut��bٍ��d��Cj��0�0D�u{�����>@�C�*=O��4'��	��,�8C7Ӭ�f���}2��y��-<�B���I����U/6hY���BD_��~���[�V=��Z5F��5�*���gJ�[��UQ�@˷�/�p�=�l�~T
}�a ��W�`����_^��&ao�X�8s�����7>��L�k�ek�h���ap������2�~r�E��I�\Q��B����-��4���-)�Ty|>����A��e��2橤�ֹ�"��m�-����Xt\@�/�YĲ�as:����k8�v����D-�����< ��kq
/���-$aa�F�4w���%��_�i�"�&�B2�j����:ף�}s�����,pe�3pܲ��ᆶ2��(��WW����op�s�e��;�r;əu�㳂�^H�#���T���]�+ˑ�?f	�d÷E�����d��	��aR	���q!M����VZJ�)O�5�}�6lm0��L{�~!x�x����y�����we�u�"�S
�5f�f����J�#�%Wʄ �<Y�,�'a��V���H��9m����plMӨ�Ev_qHMd@p��[�Z�BgƟl�^�kC��5�X9���2�?D��V��B��F�*7���Fvܦ�ۡ�1�o�X���gAC����
�J�ؒAF2��Pl�өC�H���M &�R2���6��8����S}�E@`��M)�.��TO9���u��1�
V�/J����EN[v���M��)�E��ҙ��ro��F��,�}�������� ��®���=t{H��W�������ߪd�n�5/%�,~Ɓ�hكO�0���תW��T�E��yM��N@5�n��"�?F��9	�H~0,�IhP74���:�K��͈9����!Ò�j^�g9#)<j�Y;�J�q�u�P[Yȧ�_��-�I��"���� P��f���Z��C�Q��F��q��E��ƪ� ���zۦ�ΦPun	c�b[�/��b�� ��9@wo퐽\c�_�ft��ϥS�)��Y�	��o��≼���8�y�,`o�B��b��5��'�I�����]ED��p��R�t�����ȤXO-XFjEO��ʐ����������ܳ]��Q�N��rz����2��"������@�g�2������꥘�ݫ�)���bڻ�i��Щ��A:�$�690/�:�sm9L�O�@�W��L�
m�R(��]Ђ�|�c��+��ٕ���=şƌ��ǩ�fT�2w��+�����xzgWr���:�M�t�wU>(F� מj~�C���E6�;�E�<�1����6-;G��\n�����$t��s�Y�5�˜GW+�d��ȣ��lo�/��*{
�����L�x����UD)�6+����I���Ю�VS�h���|I�5�J�r/���5��n1�>�Υ�����輦�	 ��{֗���Tws��'��@Zt��v,��"A�+�K��P�4d;C�=��d�r�Jp�
e{��g��a\�Zw���
�D~:�JtG)_0����N��s�K9�7Ԑ�� L��I�Lö*����{p�i�l2������H�:�H��E�8Ċ��n���)�Դ
���c������[�S�[Y�BdHI��-�po{b�W(i�.��V�U����lZ�z}s�G<�D�m܈(6I��ґ��/,ή	��= ���1�	n�ϐq��<���3��A�{H&��%�5y����,��G�|�Cљ~a�
^JW�¹�hy���2��A�����JOص_c����@��>$T	���9�6l�*n:��Zdc�h��x�=N38�a(�eTD�T�"��ȮK��<����.I���.��l
�='f
Z�]k�c�:�=��4
R3U�KF���f��D֭�@'.#n���� \ � �j�Y�kG�vH7h7����$/��Q��({,�˿���@�{W;�\�Y�Q߷eQ�gm���`�QCO���e��-��'�Ψ��Ǡg�ՇB�� ^�BW�4����a��'(��`�VN�[G&ˡߡ��_S/�07w���E�_�����^@�\��p�Q|t��E�W+ॢ��4/�@Ņu�e2 �U�l(Z�G�A�ď*k��3̂�<�*����a7"4��q^X�R� 7z\�qDj��k)��*a���5b���9pb�gcR�^_�po}H�B���a\\��$�ՙ�8�!�����h	��u�#�#8pB2Z� B�Z|qE��!fJ�5��o���u�d�=V�*7"���fNC��d]�k6���L��L�@�q��<���B'�x����G��g�<�6�dIju�˷�3�R�	�tې�VI���D���,�'�N7��_����ƍ4���AR�t�I���.P,��VG�C��0�s��A
)X4g�:7cʦ����A�ԕ�"��@s��1��f�ks@�3%�\ć���V�c�1HC�ݻ��g��P?#���]v����9���#kp5�v�Q���[�9>�VįL6+�\�}`�]7]�\������B��sH��]���!��Q�{\}ᘒHNA�����GA�ki���%�o��@����X.�APEqC�^X{��|��b���)ke����zd�{�bg�@��Fk��+���J��ζ,!\Lm��[��T�-�f�N�M/���ѰFIvi�r/��f�~�-�rխ"{ݶ2٤}s.���$9;������ 0Y�va�N���p���C���v������brs[��H�0���ȣ�N�^����l������;��*�+�b)}�f�f{]�x����.2>����U,69	��Ĉ�>��ߞ���of��-�*I5$7���0�JT�j�E(|x�|1ٱO�nYe��:Ժ�g�(@���0��uu%Fu����v��5�|\;�ʓ��5A�!G+�ԁ��ф�Bɝ�l��@`l��g� ݋��	���Vˍ\%w=_�2�kf6������ Evb�[w�s�r��i6�:-O0G���Q֑�+h䎂nn��ʇt�#ۜ�۹�0M���cݣ6;�7|���Uԃ́0�^QD��3��]	��'���ګBv��=)��ˡ�S:b2�N�,x�e|�x�^��ePĎW-=��O'�(7��v&q�ەT��")�4�!�#�˲�.t�te����Yz����?�E4�(Y��1���nSR<��E�x?ke��-ׅ�=�s��A%���!��)����
�U��>�A�=�Q������/������ʔ+���N�`�B���(��Xr[}/�c�>W�3�	��!����0T���:�P��OF`�k��F�Du\�����QN�ꄆ��j]��=
�ҏLa&$3U:��8���X�̮Cr�@�s�~yק"p�9���
kGda^�Y��Z	�ﰻ���`Q·�p��fU!�"��B���<Qk��Y����_����g� ��wޱ��j��q&CE0]Hp*�m���E�,Nq���3�B�J-d����S�$\�Q6����D��IV�s(O>��O�j�:I� BR�;
���TF,S��ov��6ݲ��
�nl�s=��qG_EbE�::���-y����[g�m�aiM,m;y�z���xjM�L�.yw�[�*S��	�P�pZ����Z[���sm�>������_��(PRf�D�{iZ�ރ�
|륥 a�o�gl̀tQ�_��P�,I0�a�s �M7E�ӈ��Fn��Q��RXF��t̔/O�P�e�bk�d! *�ȥ��5��F�,�l���E��莆\���s�ݨR�[�.�:��i�c"gY�R]{���:�����
��[��Xy%��� @#�gU%���z\�*"f�F�f�$��Cp��>�0M�):����Y7o�qE ���p�%"赉a3��]/���t����/]�j5�<R�5��,�q�3~X!~h�"�\Dz��(�Y�x� ȃ��`�݆v5ҩ��$Iu�
-]��ҽ����5+e��8�mn�i��q��pDt{�gW�|.��q���x�Z�P؞!���
��`?��ږ�w1�<_��}�s�?K��|���-xV�L�����Þ����!ޮ;#KXy��"C�XFK)5�7;�4�+mACl����r��AH��u�Kka��^���0_�t��rD�T����J�<��p'�Eς�e�Io��8`�[`��|�;}�����T_N�/�!ngL"�5d��l�j��1���pFZ�v�����~��O�l>����K��_g��9(�"&�����̂�Ҿ&�zJ
������kg����i\�[���ꀅQ�B��}�w���y1���@x�u���E�ׅt�Ԉ"	t��dmpR+L���:�u���;Z��J��xNN��FKH���$��}rteM07�J�2����Q3�ܧ>�r%X����{�K������X����T���$�	&�N���O���r!!Un����#���̬T��`@�nQ�$?��R&Uj��� V�9Bh�.��Bb �"ڢ����nwf�)�I��W�Pn�o�(f��l��L�=d�c�c��{��
��=�HRִ��_2��^rZ�n{ߎ?\����h1�#�Q�m,�M^�V�o�V���Z������1B}���IN�Yq;=��y���z�h:����H9*M����=�˂�?��!��?��Jd��u���*oQ���p��	�/��G�D"�`�P�R⺾/K|�h���_�'��!.x'����sR�����gy,`փ�c')�FX�S�t�r&�B�6���vTɔ8ZI�"=qXAZ&� ��zc��QGFB�Ǵ5�	eN���I�+��H�_�=k���Л݂*�t��
Z����=�pـt4;{3��`�1?����2G쟤��8�����p({���#�}+ y�E�OR�Dk����zz�PP������v|4�ɾ������1 �=���	6s�+�r�P�?�ṅ��Dee�������q�B͌g�-��O[��pf%�0����zF��L��7�����ˤd]�_0�b4��O�dӂ�ô�g��T��l����O%�)�p���s6��ۉ�h{IШ�:bTudV�����@ף��a��#[��W�3�<(�f�d���s;�N*#]һ��F\ݰ�C���+� ����Ʌ�O�`����s2��^�7߄�i�bxn�icV�D=�J�/�s��\����A4JE �Ѡ� ��ݜ)S�;�N�?��K�w��q<���av���������e�ջX B� B�2��Xn�FA#���A����5d�6�p:c���z��V&j����,{!�-�[�`�#*H&}89-���c��4M��-)�15���|x��륱��J>:���6�D��)��Ꙕ���:ƴ;�	|����������Al?/��Y% ��V��)$pk������Ź��J�q`1�غb���j�;�����͔X
�t;�_�)����=ɒF�:�<��.ؕ/#��6���O�dQ8aXL(�$W��KТ���ɭ����ی&6���F
@7 �';��U/�P*�7�9#c&�N,r���j֨�Z��X�G�Xr���r��.�F-����ȥ�]�E�>�E� )N��+��Y���E��U�*tb��O����L�ｦ��h�����!#{Aʬ�Є�WLU
�$���M"e���;I��l!�T��,������h�ԩ3#�|O��b����[j/�a�6ͫ������m�nd��"v_���vh�.����L����?��'���}pY�.H�G0�3��j j5��o�R^���M�z3j�(��b�&��o/�qDj����D�͓1O"S�#����i:`�i���n����-�x���K�Rsp�"��y�JD1��a(�[�UB:�M��J�����d�߲~�ٵP L��@b%�;��L���K]�JPy�t���^�I����s�i(rB�R�Μ�&�_���>���S�=H)B�L1��3��8L��s�x	�v@��*Ra��Q��ca����F�X[��lݯh���qqų�8f���ɡ�Ԝ���H����x��Br�,�!�x�z�,���c����7m�3�M�B�f�Ñ�]+Yi�p�|�1g����J�J@���iT��j�EYѫ��ú���H��[#1/��o5ˏ�
N'QS؈�",9+��U4X�����F���b�I��P��S��N��l�R���J�}^
��[�]��n���;ȩ���ţMYMV:�1`���z�jf�m��6�s��:�:�KY=%,���⪙�������%��8����d�/s�����'pu�~���׭����%�E�_�k̶r�o���\���q�#��;�ЖpW�kצ%�cyE"Ŵ��j�1�rc	<�\�G��E��1~�%�����{�4՚�k]��R��o�|�c�~&:�����&��ژ�Щ�}��}[k4gJ������r�%ˮ���#Q�VJ�%�`��t��?]�_a�dc�Uǖ
\��㞨�Z������A�9J,�cz� ȡ|��e
.�蜢�����[���:�#U}��Q�Ǩu�CS�6������ܥ�Ӏ�[)��q\��х��#G�1�����9yc��dI�W�9|�_���*��s�;SJ&~�'�w�7�BE�J�+^��C�N}���q�4��ۨt����g�����i�7 Ф(N=�oӼC�L4IH|N�[z��$+ڕ��[ ��T��`��k�_����T�B֝Q�,~8�� �W��^A_<:*l�N�~q�FB�`�r�ta�o��B�˂�h���S��&}WCa/#��C�*.�r��F�i��x�y�aR~���ݟ����.'�&����L���KM��a�ٸl�!�Y@��9h;>V��-���e�3�_U�����΢�4h(ó6���1)�F���_.X�7�WR^��i��"����\�9
�q�R��৔��D8�~�vfY�;�������r��@����K�p���?��|�n�:L��u�������xBE�T�(x2~�7�A���G��	�p��o�%
6` s/��|2U�w>��I���:�ycph�΃��V�歔����k�o��C?�#��Ϝ�*�&�`����qY�I����E���)��)'�Ƹ9�?�f�E�]d����SoZ/���IG��� ��B��ST�s�w�5ڛ������P�]w�mc��gmIV[ia)����\o���I�r��bD����O)�>�kn���L-�"�Ʌ �8>�����V�6�\F��a�H�����1�� �'����#);�3���*y���W�݅H#�� \VKL�+�n�;�f�H�L���H��Pq�Z��C� �����З��F>��KD�7�kWr����Iњ�Դ�3w�bk�u�/=g��N"�Y���H�g^*�-�̪\p��7`��hw�9R/<��^si��9,�[�
��l�������y���O�Z��z�/�<K�ln]��eQ�M��H����z˲�궭�bʿ��WIWˍ��U���\�f����7�w4��⇉H�bQ�w��~�eTFDԮ���;�<�3�ɖ�Vа���Qm�_�t꺕�@p��:|VPnI _h7bq�,J#ȕ��Z��vx,G���������a"����G���+�"����^z>aԘ�V��Jʺ�Z�㵧�����
}��Ws 9K�m�x	UMx;r��%�fށ�b鳣����������rcU�s�O#(0�j���
���CgCMv��E^�l�F,�A-ä�OJF�y.#=%��`)��i�v�G�Sm��i5��u� 촅fu����oD���f�T`=����O�Ұ8���|�$T9uTd��	��LGh��r{B�O�m.�
���R�Q�v��fO'n-����vȶ͂[�E ��t�[,���c��T��ÁP�R���N��'��.jO-YW�2���<��B�~��s���4���Ɩ�bu�3,�+���Iw�d�� ���3Xr��!J�2a2��/�7�T�}G�OUvN�ݗ#h�ŤXH�LNݶ�g��\D�0�YɎ$�:%�C����.�q#���H0�O�l�o�vg�Íb�W��4�<G����M{B�:��;T�Ñ@ܩ��Z%���"�G�-����K��춤���Pݽ�-�HA��H�{�er[���������m|��pp�m�4�ظ�B[ch��&y��]��;��
ܟRJeR�{�� ��� _DrU� ��q�9�Q̠���ipl�Ӂ�&��#qW�5y>6h�F_ŉE���оv�׼�@�fm�`�v�[���<��L<�I*��c����p�V�
����_�H^��ѓc��z�O�,���D��A�ڞ��%��N\-$��)�U��hX���XsF]��42v�WՊ���`2�����є��3w��Ҵ^��D���+w�*��Ӵ���s�Q�5�Fk��?o�Ҡ��!��9 9�"���p�����Ԥ׺�ѷxP7N7����w�Q_�`_�HU�	9+l�#W�4q����ٶ�>86��m���*�"�tFd���48�+nt��3�#�,�d�+e'���s�&��zâ��	}ڜ���%��6�l���x�#��8��w����1n��L�`�k�Fͻ�S]�1��/r.��uG�D��1 z

�8&�x�c�)��FD)�;�_>����o6��Z1�7�w�7 E�G�6 N�F�y��1�i��%<�z����S(�J�K$�(D1S>�M]�9��Q7"�)/%*]���A�4^O�庣�6V�c�Z�
FY\2ѣMI���Η���B��,]'�p �h�A x�2�Ն8�9�����w~"m�|*oU��	,Iɒb��Cn�����G!	@d��y���ܟ�>M�o���>g����GJ�\�Ѩ�K�{UZ�'�&��3[�Q�����|'x�D9*�G+��sa%}]2B�1*T+�k���m|����Sg$ݡ����?CC6�_
Mڒ�8o	��B�����B�V$�O�Ã��B����w>N�]���G���ͦ���E�Gj/$Jer
[�x��$�k�⃄G�U/��3��I{���Nak�=~���A[�v�z�%�
� ;B��z[[��?�ϟ��@]�u7��&5�S��}���(n�r��.�(��=
�-'5J��$�rWX��V��&uP;�rJ�;���Z�ü٬�P�в\ɩ����3Z��f��M
�)Jξ��XF�~ZynY���u�?˱��}��Ҳ�/�^:���iei�'�������o��e(��r�i� ��Y�ȼ�C�$�S)���]�Lp)TV�y�.�y�0:Z�kIHO)g��	��.���'d����KA7885�M��ʊB���R](���*�<��U7�枏W��@���.޼g!���Nq�U��6�A�e�/tQl3������_�NFD�;̠:�$a����G��N����|ɇ�8r?�~�$}@M&�>��:`!��@��3�y �\(i�Wp)[>�:@f�x|x����T�����w��䕒��F���5U�.�eZ#�esA�ZC�*X�{�;7��m�J�p�s�X�xrD�[�ͯ���V5[R'RA���O���y����c���uj�@�l�5�����`!$ʠ
�>�w����(�G�y㩐�����σe�K�⟻'���5,���k�����M��F��pJ��W���n1tO͛�����c�W���s����i��L�+n�RC�l���B͕�R�Q��3#��=f~��_�(�@.̋���H��<�2�;���Z��Vv��������[������ˬ�w�� �Y8��͗�
�k��R��={�\�\���3�}��x<�����9��@����^� ]0���z H����g݉ReXl�3��Xnf��f}��3����)�W !/��~�uU y�l��*��eծ ���p�ᚠ��-���Hч=(
����b[�ݟ��v���.L����@c���<��l�M���h9�"�7�p���5m��݊h{$�x�7��k��I0H�)��$��U�c��%���<�#���~(��h�1���<J��j�^PO���c���>�´ٛ�:�&�%��"GW3E�������c�F���Msw̗o5���X�~fkb r?,\��9��Ӧ
vF��,��\��E�J�qX�A�g��>*��l��e$$�ysoݢ�Ŵ��]#��>h�]�ĸ�K�G4)��>5�.��]�UY�F.�.8��H5T��A�ZC���7_�[?b�.#7�Bx�k���/�Q�Z[PX���K U�8�2^�-J�i���4+ļN!=��.^����Mt(������i�p�`dF�k��f�ד����.�����hʴ~c;u>��_�w���,)�"�S��R��r�m��2ڰ_�y�A���7�``S�k�k���6�86�F�����q�L���j��T1e/j���YC���\�7�n�GP�^�ح}0�5�.�1�j��n�����{R!��v���!�G�׼h��������=��oRW�|�s��1��=�*탭v`[�a�OC	@�@L����f0��s[=LoQz�߮
����\eqkC#n[cO.ف#xV�Z�T�
����@z�P��)�p��?>gm'.���"�����G�1%��!�~�	�q�_d��b/�ɣbK���,��� �!2<�	yαc;̍�M��W�E�&6P�a����X�q&*^�`��.t4���̙��nVT�_R�75�`���:���+Ӊ6��K���:��C|�#��yU���;��a�[���\>w>2Fp�]�y�O��8ш/�!A&җ���Y���S�>������e?���ϱ�)I�J�{o��{>>���dr�

�U|��y.{#I�������Ufj�g��jL�_��t��MR�Y^�3�<,q1��ZV/x^V&0wYb�Xܨ�Z-u�#�<��6.;#^oMyA;k�H���HI"ϼ[xqqV2�t�PI�Q�X�$c��G��N�ݸ�Nޙ�KNII�la�ꦎ�ϵ���ғ&���Ǆ��<{{��sА)=~@K��o\�:l}&e�V,\�[���S�p���UO�1�~#�֗��;�S\ҫ��-3$\i�x�pK_8���:s�T�L���N](��H�r���s=l�����~�!�yQ1ށ��	�Pr�DX]��M��K��l�L�u)\E�5�u��Bx�fG�%�P�������e�F�rU:"
 �\JK��56�J�p0/�d@�}�b�f����(��� ��/2��q	8?z!U<U�﹝$�H����%�J���U�?|��>��w-v� Zd�!
P>+'�����4T�K6q��6��栥��U2���in	��j���k!�)M3��U�}�P~��o�xE���7�D�x(�����r�1��0+<[H�Tt�Y�+G,�H��
*Xi� d�z����k▙��Vm{���6���{K+:����-��A`"U�f(R�W�Ô�az1W:�b�ʂ���wb��G9e���6�����\$�nwÑ3����e��& T��W$��0�C��0}���W�eTI�/^�� �!ǫ��ZQ?���k�� �!�S�g
�úz[?Z��������ٹ�D�8�OG��t����(�ɴf�i�x�}u��E����{%�"C�r<n��";�w�%9էۃ\e�G}�M��B��:�S!尫���'5�+;ߙ���>��}6WeV��~�߿�,�L�(�7-(? P�zI��#u����/^��{�JÇ��SNM���$u�	 |@�\��˨t��׸Qke��q�!�O���Yr�)*�k����=�����뗧����3ǄM%E��!�2̽2K�(z!�{���G��n���ZQy����.�b�7nEmM=2���6�qI�Wi������s\���a�&4�D�Y�Ӯ��Eܕ���D�ԐM��fR�%��ǖ��3�9M�5-j/�4������\U�l���};���1i�c���{�9y�U�(�s#(��:��Ȼ���=��m��h���V��u�ea��Z2�CH�W��q��f������K7�\�F��^H��Fbq6 �VgV���	{p ��G�����`�)lF͋���è�94�2�>�tXFxhQ�#�f,����J�*]ۦ���I b��> x����sS�2����ځyU�jꯗ���(����՚����yA����j�5�,/�{GU�1��������
�1	����l�T��i[�b2�|x�8b9��2-La�$n�����>����!������	=Ϋ���m~��b�����Vz�s搐jD�&	w�V��V��䶦�֙�C���bۯ-3櫈��E�1�J2��;��N&�z�t��b�2�R��w6��^r>�6�����(,Ӣ���1!�-}�q�zk���"���ߐ뭥��mW�e2�$��^�#	�1�C���%����Q���Oޫ�1v����r����B�o�NQ�1ܻS���?����zr���h����\	��ad:V��q��,�� PzP3�%A^��7�Mוm�PtTyz�3�ި_#���QyZ���y���	N
8�i�i|iU�g	�����������N�#l'�=
�u�n�Խ�K���w*ܽIH�L��)�%�j��:_S�>��y����y�?����Vp�?u'`ϳu�+B��0$�e"����g���>!�vW�Ǒ�����f�U~.��*>��{���0��ʹ��i�c��g�&�����0�<�,�������<hQ�N��D��ZV3�M8�&Cc"5��A�hΐ���h��${�]}�Nytfj���ҕ5(>�ȟ�y��4�����������";� dN�3!�s
���gҡ8��)!w(C�f���g�;����<Q�_l��?�*'5TX��e`����1�N;>��A�}��㡜�'��Pr��i��wY8�gWS�̵Z�&�0�FAj�jꆥ��2
=N��'-����!zCOn��n���VF�!�o��u(�rM$�7��O�<�����@l�ί��l$�y�(h�2��U랰eH3�y���.�r�ēCv>��+�Ȅ�� H4H��Qg�#Kd��`ۍ�5�կh`ds�y�
�(�Ji�7�G�j�p���W��.�D-5�����g�p~��ʤ�L��k�6���w88��6J"^8��k�h��/t����l� �q��6�n��S����Y�¶��r�����x����1�'��G�/Õ��Ά��f ��#��1ix����Q2q�Z�	lЭ�R��H�x�������}Z��D��q^J���w��icԅ�햵���k��0�v�d#�k���'�����$�W��/KO�Xa�A���������r�1�v1P+��_V�y������s�U�B��;�>py(�c�5l�`�<�	7��1̘ST�!�\�}��x0���"��;w�s�g+x��&c��{��=ζ/*�WZ<Xnޢ��^�� �Gō��|0������6��m=�X�j;��V���b@YLY�iXMM�B���2�Ph�r�إ�f�٩�b�Ni�7p���l�N<6TM�m$J�������IRM8d𚾗U�$�����W��Q���j��1z8��G��y$i�J�&[�?ߧ���=�M`�x�	��|î�3>�^���Q�YS&PPg��``� ��um[��;�C<o.gA`/#��9�@X��WP2o���~��v�2�e���a����Fj|��p���]�a4v#Y�jT�2�(�Q�Rl�e~�@�
b�d`c*�
ѽ�lG��t��8��Uy�T��ؤ�6��i�����]����^ m�;j�l��-�%F�hR��{�N"�*�T*+��)�ᅔ�I��yE���1�\it�$�SUZ �q��?8\�pח�a����
��닝I�������7w�CPC�y<�£S2��~Ȑ���g׻U|�)T ��<vt��Է5�O<�*��`�=;��7wo_%{�;�P���l@�z�Rf䔠�$ �����1�P���LPkl���&�>YD��S�Eq�d�l�[��rD�)Q� S!���,{�}nJ��@�#G�PI��W;	8�:90Qi:������j"��(�&����ő���.�W��Tm�.�x���m���y�ڵ��l+/����:��銎$�w�x�Mu_Z"�tf���mœ�(�J�ac&��9|�orf��[p�74B
7S�zV����JOL�fr#��i��5���Ӆf{8�:/�~��U���Rp����U7+#_\������~�ݘ����͎�H�������M�Be��p�9>�;���3�aӠ�Cl
4�����&�.B��x߾�#:�H�6��hC@�q?�p(��RgA�t<�N���":���k�d,TKT�S���
�:L�,�B��qWr�L��(-Ihia�*��?���"���s��[r�����u��}����Kn�F�� w<+��=���x�����7`Mr�� �e-7���͐^w�
�:����b�w�B ]��|z�6`!��B��`��F2�q'���_X�<s�����,�Źt��+a�q��7H�,<�r�֜
��nU"\�i��X�m3�����֝,=@��MEMZ�`#�lh5Z�-�"w��Hͬӯ���$ر-�8�T)����u_x:*z��;�6ak�����	"Z���I�}ȷ��F�m�m�#����f;���@��:Q.��9�kDG�3�
;�,�G8j�,N8��D�e�	��Kq0�DǢi�=���\4��H�l��;tI���в^E��y���Eh7W
r^�z�e������'�쾵)9�g�5݇$�����'o�/=��������p^��NA���V�0,+֎X'��y�ڮQw�*�s�2$��5�+��xAa��ޞۆH�i�B=%Ǣ�Y�Ǟ%4,���8��`p�Y��Q��%�G �6�p �S�փ�Y;ݧ�H�"��y�	��'1�O;�(~��q�O�pf���|��1T����B��� �ڌ4c6��3�s�Z'�d��y:{�_��H������	c͋��:G��N��̈́�?eZB2ԧs�bw4�D;�H_%"l_�ux�A:�
e?��ݑ�m"TV��G_�7(���E ��|2�c��60��Q��'�6��ۗK:�t�$����nt�ΐ~5=N����V�{d���7�nwG��ō@l���ЛWhn�����U��r:�?��|l~�1k8�Z<�6� �H
��ՏU�P��B� 1:Z�7p�7=P�
r����#�
f_F���vE����P�ܑЭ;q��(����R�-u%���&֞�G�~q�u��BQ�f�1����ē���V[��b�"zz�Cԉ��J(�)�͐�l�g�m�M�!�|U�ʎB^U=R6ٓ���lTp��Qe,<�3F�v�l
��3_-_�8{���z�6�+��Z��k�v)q�b��wgumv)���i$��%��}��Ϯ[�%�65,���%�2�s�ײ<P����վ�[��F���3���j��f 3J��v���O1��s�'k�f&ׇ��e�8W(�cA�O��u��ތ���zB�m�� Ӈə f^��|$��Ё��F���量��Np�����h���ݨ�V5�A��h��,$-����[�7�g�<���]6�>�ϙ��z�9S4f�O��_Zn��í,�]����mڕ�5��G5QQV2}i��o���n Vw;Sl��f��l�bֿ�d�)&�z�̒O`��-/|5�[C�9�b��{RB�YN#T���hb}�����3>��7�|9
�������2K�7P�ۻ�/��ߵۨ���1�^�(�R����I"�1RGgn�oYI�r^[ŉ�dɺ����J	�A/DL�PH�Jg��	��uJ���0�Y� ��a37;@��e��d1�!����Sx,�����>d=���,ֱ�ٓ��S�`���Sq�$J�A��TU����Q].� #��5���>e4��$pw���& 4%���ަ�k9��,e��f�<��(L_�_�e�a���g����?:C�`���i'M	�ulw2L��c���Wc� ��{��^}{�#��CN��`+�v	�4�U}^S5<���� �!�ǲ�(����� mH����LZ"D����n�����R�%ig����s��ۖTbpM�(jUlL!�*+J��*vF� ���~P!�9���&�����v���8�	�q;��Ub�jn��A~;���}���d�N^t��;�]sk���O?��mN���C�9�ʱ�+�6bV�Vt��j�t��o�!q1A�P[�$l�s��I�e����T�*�,���Qia��%>��M��̠Eܪ����B�����MY���+�����쌐���= K�����a-E�i���r����p ��q�r<��d�[�J08����j�|���o��mNq����]�ZX��	�/(�����F#�!�o^S�}���PG$�P�p�V��H��<�A�e.�GO��Ҹ�6 �T�$��n!`Z��{>���f*�;�2�S��[��G|$6.skK��P_��:���1�y��ز��M�ؓ譄�k��jUS^��Z�A�m}��T[�$pl�[T��Q�u��,@<X,�"��rt�t�������vc��~�=J{��N����iD����B�^��lTs��G��CXWb7�J���m�ia��"���q�V��K���/ud�7�!�e`�� b�cO��5^Џ�>bǣ�����
F�v*J[�[|m9�o�t��� fiϾ`��G����Ū�ڛ܅Ƒ�6�����n�EE�.��a#�C9�d[�.Ӽ0	e`8=<~2X�(J�SS���C�����*-T�2�n��ѕ׈�����D�,e�L�T� �rqz1]�d[�p�wa���D ÌD#�xņɐ��c�O&����{9�,
���A�;	C�*!ai+%�8#}?jC}	F~3g�	'�D�*IfQ #����}P~��:���wa �"?3cPtz��}ɍp�â3��-��o=�>���2�������F%�-5F)����1��f&�/Uv�sTS�|��Z+����%F}m������P�`4����ϕ���8�N%e�h�`�~۠�~�"�_�ۧ�?��2�4@�1���tybx�nR{�^���#c�;��R,�H�?�g�n՟�2�|�s��
H�� l��vBRo�ٿ��zʻ��yCH�̞��ǚ�]v�yWD��{` }��Xk�
6�jk�7U��a�+�̥��n7:�O�9��顝�p�ΎÆ3w��0�'��'�-���8�;J�2RBi��Xy � 9SQ#̖,`KA�s)3;r=�w��{����k!8�mb���C2�Ouk��K�=Q��&,�8q�G�2�V*��k�)�ӎ�dw��'@�u�����Xݰ�B�j�eK$��U)�\�
��ڬ��1�U�u��q� ���� �;>�k,�z�F�����Wōq�j&V5�_ĉ$#���AǷ�uW}D
^���ȝ&@!2��8N����x��z���|4�G�W�S��V��֠�튑Z����%�Y�'\�np�K>⭐����>IXXX����fv���P�e�6�X����o��ͺ��b�㰆U�ѓ4|�1��@���.U`oMH���tQ���/$�ߝc��-�F� m���La��H��PW��q۵o�9�^��ޔ�����B���mlp��<7�k6��bhƙ��Y�3�A:Y�����r�Y>?��+.0�<I^��VԦ��N�i��3��}�/�fW ӁH��oˍ��)������j�;b�Ԧ\NFX���jm�O�Z��ycR��A����^����g�'�K/�xP��D�_'0�CY$����;�jOJ�I�C�4M��v��
Z<*�������rBZ����C_�Mj�C���]��j#u?�eId�^7��'t��˂���
)�\O��-�K۔"��_}�ot�4���e<�z���i��7!|`���K
R]�ץ>a�j��}�'�j�RHɛ�!�@�MRe0���]H�K�^��[p�)D݄';���{J��k�:m-�@r��;5�o�������
mz��s	�-�[�CG��Ve%�I��y�7�?�	U6��;��sX{RQ?]�Hw��B0��$afnxn�e?�ېK����n�>XB�H�BNB��q��D�@wmrs��,�!�T2�[��yD�bR,z�&?-�+=�eE��>��T,}����p�zp�i�휪څ�-]��v�A�U�{~9F�I2V`��ԏ}����n�ў(����u�8������|�?�u��C y˛D����U���z�TiU$H*ͳ�砄�L���{����UD�B(��!(Z�l4 V{�S
�cQ� �,��0�}˿X�V��?�.��92��Nͽi,}�}o�8�<�Fڇt! ��qo3V�{w���
y�^�/�ó��p#�`�xSr↋�\J�D�>-����]��4X�r@yc`P�mLH4x��7�FcB���?���)�!�ϒ0K�����[g��m��ē[j9��3�L�:�5y�cќAe0nN��][�J{�-���`�9KP��%-�yU��p�9����`��)���ѫ��S�`2O抧��C�5i��������sz(�T�>��y��(V��x���\.	�6���4��&W<|�F�{.X7oMI����8Xw	��`�X4��k���=��B����~���m�pX��J��G�`�Ce���H�pc�� ��	s�ǫC���;��}Pq<�����|�-�O9�2��sU��|�(�B%�ʭ�ς� �a���@u������]�m )C�T�x_͆8�hTo�{���N�
 �/��	����&��>V�׊�MM\G�X���k���olCW+����I�R�<h&�u������H���rs�����q�F���d����S�o#��Ml.g1�j9z@�U�2��ϳΉA����]g��
�vb��U��n��,�B����vU�_�^��9f=F��2{�k+ۺ�/_Vt��J6X��ͯ�~�ec�V[z���_�3	`zВZN�W���qƂ�/�f^i������/DX������g����b�\��%>��S��1�Mr��,�)� 0A�ZNm�����ؿ�9A�g��_����ǁ�����ъ�'�����F�f��L��X�k���������ޮ��9�6�m/���E#,4n�c��T57��1�c��˔���i��V�-�\�<�6�$y*�i�
��=>Og=᫸rt��7o^�hz��'�ȌpP�0�m��h�����G�}�9X��^9F)�
�!Y�癰b�IAl,��4zpY�۝��kI,x�ڔĔ�<���?L�[:�r��w��K;x���4u��R�IV"���W|	^nИ�1�W��F�^R��ps��/\8ɛ���C��Ħ�n�-a&�]F�8-�Y���,�gi��k,��3׺�Q�M�E�+m��ӎB� 5�Jq�i���f�T+V�Sߨ�T��1��Gj1��	�z�*D(���v����Jy��,��t8d���-��{B��%�jҔk�p~�)����+��&E����bIрi?�Ӌ]I8M� v��mit�n�,@8��.��j��M��W�	�\���"�ɔ*�-���E���PJ Ӣ�a�oh�g�s>�[�X�-2�wԮY���5���b��PH��t2�y��r��g,.0�P_(rh���k����%.��_������`���p�?�� WP��AlNs����Һ���1T͛�n���Apq�:z�wRڒ����bm�j�Q�M����0G�Qq�F>4�?Fв@q0l5vV.!��;Js�[`ܳ���:��߫Sw���F��a�,��P���� �̰]=3�Y�U�.��\M�&�ʑ%3:��*f[>��_���9���H|eK<��H_����Pq者�Sf9��a��IL�/��^�9(�`�3�6D$��.�,���C*�E��?������̮�C�&��{�8�8/L��k�S�������b�,jw�&A ��1$�$e��N~�Ʒ�������5��@�}�=ӛ��.~]q���9:���_;����ZFmg�������~p�Qr���/��L㌠���a����g�����8�ؓ����4@�A n���-�1��>&8���_P_6��:�1�3Oe�KT�H��I�%J�5�����4�	oFH��,�����n.�� y����9P�0�i�k�0���Y����m��V��X�X��U�F	 �A�nzww�K]�w���XUaDc��$o?�÷�ڏ�*ظh�! S֗�@�S`�W46(�=m����H��-�l#B�ˊR���7�h���RmX�sn����6�U��h��G_g(�٨V�_��'V�]�S��,=�����{!��	ʍ��1�`G�4D�zn7�zu��+������2f�a�'�4fE�ɯHA���M�\��|��|6�S���-���߲�!*o�nHߙ T�LQ��a4��V�C����6%�n���]�j�0�`���fx1���5Q�zG<��"��������g[�`C�o�Tn�5}�8[�3��ף_փ^��>���������Eeف�P6�8j�U�|���������Beg�\��vp�24�������v4��c���J2�=Wz��)s��n��t?\�/(QV#]�@�֪!��0�8SC���/2$)��KٱT��O�c��b'�P&���N�)��J��?�1>�} �� _`���F���{�w���zp7����Iq��}��7�h-�W:.�D��O� )f�p�f��V̢l֦@:�����Y���Bp<]�Zj)�<����TF����u0�	�e�#d��}x|��h���@�z
T�S[9- � �x�'@��<�gL�D�E���.����/xJC�M-� �S�5CWӸhV�m��d~Ċ�6��T76��Rг| E�����MB���CG����w�߈l&�]p@^aS��c�������!ע��tH�hn1�#2��<��v0?ف���X�}���+���Y��n��'}#㕌��w�B�z>?�B�$���"N�<��Z���{p�<�K�
UjBI���d�tx���m{h��^A.f��k�:!��x�\���l沧�?]����nMm-��KU�2
���']Q��e�B����qa����17����LO�����z/�[�Fɖ��1���8Nkl+��-#�lr(����IOj-�zO@5�KEv�kX��NCk����穛�xz�K�wN�s��F�q�L8�e��wo�{T�ن��u�/_Ӫk������D*9��fXؠ� "�@X.#X�Lg�C3M�3U�S|��S��5�%��)PB��U6�����a�+�6q�@�e*��+y�
ݒ�\�u\��R�#���h���Ă�mQg�t_��T��T�Q��P!䂳�N���|��&�ޘ�(
����5[�0i������0ذĝTF�z�� 9�ǡ�8��"I��`o��M����Ч���0�0��[k������cD�m�e��:�{�Q��po㜪K)�Z�w�#H����%]8h�5د�(����է�cm����)�F��.�����H갊�_�>�@;�Fqȯ�6i"���a��HU�l������-�:�=��!��X����ˡ~b�RH\�UR�h�aFCc��)Z�]��n�Tr���t٭`c%0���Bڴ�Y�&��As��m?e+&U��'��91k�>��Ӌ�S< ���؎�gL��U�c�d�������UG��v��b��K�
u�N�G�%ݮ* ��K_PU�Ɍ-�s%�)����؁�ׂ�;�eHvVG�`,�ŧ@��0/��oY�\���Yb�j��8�"l�"e��>���^�5Q��O��.�h�1{���@�~��d!Q�+�%��p/�3��K�0H�&���4{骼z� ̿�ݒ7URSTԈ�3�e�0���Bv�F�/��zN]o�ӭj��@R&�B��L�Q�X.PR��������ݺ�"�o, �!�ԁ����kx�g�G���������6n��ŕ:��h�K�C�5�/:yU������OvK�T��(���xu�|�.Iq��&�&��1j�'C�6v|,�(r%���v|�N|�$�j<�Q��M�J��K��"�j��X��1�=��[��3;@���Z��kqͣCn
R�b?aj���/�=(v�g��'!���+uh
]��fE�����:�u����bkZ��O+�,���ۇ�#<�.@�?8:�X�_lK�'�E�zV����l�E7+���-c]��PdfV��2Ǿ�$�
�+Q��c�=�"�&Ȣ�P6N׮k�v��p�e��qS�֧j��2̀��s�_�e�3Q��es����}��0�F�k
�Κ�;��}��®�\�0�{@�)ڿS�ɮ��P�B�&Ӛ��᎗S]/:k�L�p�|9E`�2,����_�[OW�Sv��z�-��~۞y��"{	�����DTd�A���������w�*M��f����ܱ��-���O=+�w,�'���%S2����7NLXf��j�� ��ƌ"9�f���f�ʥ��;�U�V�$�{k��'����!����'f;���m,�x�����#�� (�J�֣���jt�X)��9�]�H�&)����Ad&_#zCi���9
V���g�Zjb�����T�!G4i��n��M?[q��jC7xn?�������E������b�D�G+|G�1*]�x��1&��c�
�\��q�W�����#���:xx�,��"��j�Bq�\���C�k��(��t����F}��{��U�T>Jv��� F2�?�r�&*%�^��Ő�����ue@c�V�?��R����B�N�Y�A�"񪇓,�ō�g+}��&��UO��KQ��\4�j��-�yJ4B�l�=�B֙�C�*���a)��|�e09S��\:�f�W�x+���������U����'�	T�*/7���/�:!Y�C6_������]��9����������v�7��Ciz}��.v��{�?�N��mI
��[������*�� aJe�|K�/P��P�� �8
;��".�Ő�3�
��{FX�KL=c__~�Q�ci�?�^��+ZM��;|G��:œ*qq�Y&��K�j�8�WD1}�oz���uB���يӬ�n*��CI�}���K�z'݄����Ԣ����n����艵C�3i�Lfz��p<�6��Kɛa�m�zw"��d����7q{�]Y-�V�;�Lx�8V닐?o�>��w�*5��˓�H����n�V6�'�l���CjU?�|@k��"�l����'�$��c��I�
V��8u^�Iw���u�� ,g��#���3�[��%/��JD�N��9����
�N��1�|�ZH]����~zʔӈ�A�]F�C-��:��"W�ܞJ������l� z@1,.T�"��1�*9e^q�T�?�j���9S2p�7�os�z7�C�(�}tձ"
|�j���xj��14��$�