��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#���gXݤ��N��um3v����!NVѠ��2��?<�8��-��≳E� �����/e\W�]�HR�3�WB��_���ʲH�w*qRt�&���列���0�zC.FOz��7�h����D�B.�P�B=����5��w�kyn�Z@���[�4P����xo�F����*�Y��2P ���l_	����`_�7t��W��]!������cΊ9wm�0��+N�OYz���R �08V�}����^B��F3�[h����Ǝc���>%�
Y"bW:f�JL?��BR�0 ���2l�!CMn���R8T�.��-0����:����LeQ���Ć�9� �>�n�<+eD9��"O���CZ*yD�0l��ZK�T8/a7�����M�֚Z�v�B����лw���W|���S� {`ϳؿ�T��Og��j(>r����50���f�D>��~�������,���	��N�͓�l���_[b[!���>�܋��}���f����u ��[�4��{��t�����NjF3�usCS{�{7�W�=_�Hx[>���&m^*;���HkG�;��Ϗb���N��;���E (�xm�r�_�:��h�1\"��0t4w;	�����\!���1����x���E)�n���&�ц�<pN�����T۫-"w�>�87E$�D�.ꃸ[��j�����'"��:�hH��7�ߍ�q�'a�9�bKx��AD�Q^�J�y|��t;�{f�
��!���u��y�^,� ��u�������p5[�eM3������T��R9��o���؉�Ή�Uzy��/�^-5�Ļ��C�]���{C��&��$�dc�6��%����ԗ��Vx�\�[)0��x�#ޥ��c��#����q�����J߉c�C�_ ��|D	��P ]���=�&��ׄ\5Va�F�����a��4׺��`�
r�����h�hw&ݣ�=@�"�T�g��٣��'�.B�	ho��9-Ɨ<t���\%����=�����v��5����f�T�F����s�y���l	�4�c��߃�;L��"�N&)��|[��X�g�
�<9�qɂ��ʾ��<��K,*�&��ʰ(a��t�a�6�B���:o�](e�G�f7��\�� Al��;��O%.���]���n�o��e$2*��0+n�g�:�岿g$���#;+��	-���L���Gݢ]^&�w�=�ξ�dl�F0�PC{U�R�1S��?r�C�g�e"��ǑV�n�4κ±��otn��ɁW��$���1특�[�,��!x�b�2y�!I��o�9��íR�f�Y��E���*�w9]�$����6��=��g���|��K|S� ��"�4�؇�gH�MyT����^�y-}��M���&����Z����@��經ic*քj�&����еo��lJ�[�">�e��1*o��oխFd78��%P��B�_�o\XRקx�q�|t�e�6M2�d%N9��>���4����L���`og�߃�5�A�p����y��Ե	��y��e�]D� h�;���u:Y�{Ġ11ӿ��\0R�V-�{�R���a@`;���&Q��5��?��r]�^�T8�ً�h�<�{{<���
���m�V2u��\��3���A��@�Z�)R��}稱4j`��t&2x0uA���[�,�V-(i�X 1�xlw~p�t/1�.���x��H|��A�֡���.Ś;���bǝU<&.�YdC��8g'd���7`��!�=fp2���5 ��͙��P��5��[4��~�hr<kZ�c.��_#�.nF�qnXRy�ĺֶA�H�hd �E>�~�ڤ��H���Df :�hX�7{���$lj�'a�hE���lL��z%��Ӻ|d%�*+�Y��\T���p�����E'H�G9���7k�m�W�#g����TU���&(z܎��Y�=��C�:��.�Bҽ��gp�S�D�&3�����q��06��}ݻkX"�U�4�o��RH=�q�����Ė�e&����\Ei���TwD�p&N��];��6���cBm��0^A���(�>�Xo���`�C�jȭ���4
қ�����u!�,�ޕZhS���Nwr�� ���� )�m>���!ۍ�.Ҽ��C�F&��ݷ	<K-��z�JC���-�swF޿t�As��e]~�;��-�g�/=^�A�c1�Z`Y�RSkK�L�J����ϝ��*T4i���{�T��i���t��X�ͱ�YI���V�9��3d����]��j@{|�g�*w�;����j;Ԭ!��E!�������g?v宏�I6��s�}��/�1i�?�ed�M�`>s�טo�g7���+=Ny ��U4%z�c1��5x5��<��+���eH'v��9�3@ڗ���VN��Y��/cѓ�d��$��ʝT�q(8�ˍ6�CeޕR�P
Kj�ihf�ʡ=i����F-e��6�ZKy�XƔ�w�W�*�b��1�,'�k�	5��������h)0H��Ӝr}�D�-��������7�����YpI��T���C���D�T���3�oËN��}�,��j��Bʹ����t F���|� c��N�>�W�J�%��7�[Ni�l�q��-"�x���m_#I7���o���p��H_��/�����_�H$R����I��ҭG뙜"^1�hӢ���z�p�(����Q�kx��RN�Z���6��F�f�Ev8ԓ[�#�V�2�L#�ٮR�|��:���A�j��I��"�����H�%"���>\D��ouc�� s����!Um�`���MҜ�㠺�xWY%�:�77�f;�tO��i�ڿwiO�0ˤ�૔z�ZN��M8�b�2�ܨ� ��?&d3�e��#���-����&��u��e�3ֳ�*������-΅i��ߣچ��ņ��\�Bc�̰��'R����P�ml>�F�#<>1�ȱ��4�ٷ-J=��ou{���
c�br���e1�*�p>c8[�'�뙅��m���9��t���p�a�@�Lx��fω�	:�E"K�H��vH��H�m�lƩ_}ѵ���n w�̊�P&d!�5p��W y��\�c����|�ݱQr�>G�JB[��L��:J�w��&�M�;��R��#+	��,Dw'����|�Ye��fx0s`�]
��'��n"��_Vˎ��Q��j5�U;�E���ɍ̀��p̋��[ƾ�]a����]�.f޵�
�--%3�W�7_����kl�ν�%��Ui)�^F���'�z%A��r�k�
�+д�s�zr���y��͒� j��Y��e�cH)�8q���n�s8�[|UݮH�s����)m��}y�xt��+D��[,UE-~/h� Rڋ�ʕ�����O�)��{$�xRm��_�
�%��om�G��}�1*l��y��N
�ۼ3��Bhn��y�<!V�Y���,��폰d��� �	�B�[{��Wh��B�PdpAxHqHݖl����S*�}�A%�0K� ��A�GA5���n���j���1
`�%G\�����A�����L��,<E�Q�5�I��\;/9����k�7%	�jR��D�U�n���_�299����A�����l$��U�l��>�g��IJ�r����~^<C�!zQ��hZé��&'U=�ȁ�u��ٹ��d��l��rS�\���+٧Ol�#�P����:��s���L��!zr���@�������hu+x�9lߺ/,�\��h�������C(6�_��|a2�)�F�Z8(�������`� ��61��&��>�gޣ�x�8�kl&|H��0���x�L2�w���3�<�m���z��}}��[�����^�F����(uAe�UK��]����e�/K�͝�^���0�;P�ͽ� �SZ�׽|�K[��b�g���K;����#����TiВ�2�d�^uS�@g��%�0���Ҏ�U�H���Y^:��0��g�� ��y	����xs�7�Den%W�/�iȠ��Qb�P*����Dz����1�f��������Ɔ�zj71n'eU|k�gx�c(.� !;h?�}�ː�`i�K_!������S�&�@���{�/�'9*��T����+��e�Q�0uT0!�]�<���S�	��9��´�0�h��������lKC^Z���5�$�������Jm��a�\����"���.j�Q����V؆^�~��$�4���F�&�&x�a;LC�%h�`�����o�B�L�la�b��G�W��2���gf@�,�_�*ĥ��2;.�h��;q��Z.HB�O"u"?[ui�9��,�ֹ�j g�����Qb����{&K,RO��@�s8	����h��
f�GA���^��AUc@mܫ%�t��������c��&���u�0IaG� ����Tf�8�;�?�$3L�@���$��J�:t�����iѲ\:TM�?�Oճ��Б��tG69\p�v���<	��G���-����. �����r��|&#9zK08��^ ��g���K"�
�$�8���_�]���ܕ���r��ed�1�'�S��\LM����kmp�S�D�W�&�8�[/,ѵ��<��kNE�����Q�]��G^X�N9�3��$��O�<��� АI:kL�&`luF�������n����D谪��L<T�0H�y��f���������+�v������r�@���,��`�w���P��������<Gë ����Y�����"Ǉ�-&}1���l����F�,��#\"aoE�Y���N�7Ds:l��r�t��n��ȭ��zr�B���:`��&����h�(Z��~��,{$�n]2e�J�)�� ���?.7s��_���30�O�X[N����:�8W�I� �=l� �7�S���e_�<�}8n���=|w{ ,鎻�$ǖ��JQ����1kj������V��ZZ�btpl��H���t�/ӑ�s�X�G�dv?����]�0=M������,�]��=g�*��ov�<�"w2��
��APkB�>鵊ɠ�n�Up�A���)F�f�r������u��y���������>�,�1��K�S
\eހU%�����dHY�J5	Jن�u��`h�`!������_�j|���T�t3��𙻪ҫͨ/�	W+�1��K��m��B�ڷ�A���֯= �����D�V��-/��HH�6h@��sH��ݘ�"m%��	��R�/��� �Y��b]"QVL��kX~�˾%�Q��u`�}K��q��,N�L�1��8�g�� ��Ae�y? 8$���%�" v��ʂ�����⤚S9�S��_�?J>���d<'0��I�%Ud	���@�0����)�c-h�����w�;�L���zU���Fd�!�1�Y��,D2KBQ�ǎ���)�7y�X\ �.~�	:C�,=K�d}�e���	��Yյ��hc�qyde~���.�'�>��<��~��4�����s���@�J�Z�Y@NT���Fnd%W ��TawP����B	�7�.���=��=����m'V�r܈><֊�(�}A͸vB����9�6^u{�P����.jr&��?�t������qI���fW�aѽ6܍���OۉP�-���g�SsK���İe-krG�:���Ҏg�ҡ�zm��6B�|%�	��;�"���2��Ta<�������tn�S�����f�=�FF��NB(G�R���+�aP_Bt+�w�SCo�H���M�"mQ?n8���bƤMZ���_%�C�B0K��3����șԎA�lo{;�0����y�o���Ǻ�n�)�L�Q�Z��h�C'h~��{>��R�rЏƆ$� .JV�}�#��䶐�(�X�9�LW