// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eazSNnXcjAJGWC7e8TxPx9pmLR4ApZ4EDjRmwdaCkoaZtb4yT0gjYsyl4/kelJea
dOn9cxQw4LRImbhPFU2I6QsRybkid8e5jRejsqABxyvSsSIkFi6ifJDxMAjePB2c
febGoyALYX/ag965Mp4wnE4gbmHtQpBis+uRaqUVJ1A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18384)
/tEd3v3CYw862VfrQzvFspklCLPGUvc1aibUd3qhoUslYcd6LDoXvfQ1vA1ouXmY
k4+cVXUbuxxHkKnYtCzioA5NCeOnAP3VW4VNVZ3ZOhY1xEM15YStswutxqsNszKH
Yi2vUGgKNLGkn9mtYii5t8/XBzL5g2BY3UiAbSFKiARv4gl27K0o+qXDO4YMG7Tj
/GBxSz/c2dB8Ez0w84TsvdEaDfWA4Jn+qTJ1dyL5cbz3I/+SOj/Y84DydZ8MdZZR
OB/L/yKoNg2lBxaFeD77hlzuC4rLGNl7OfBVNNk03Mrlfr8L6JNEOKhjizJHmtf9
nyHQ2XENTT+AkbvlOVwO1EijR9XCcmiTv3/tozv46MPQeocYD1Mnl7Vt7c1WSgKd
kQtyuWd7vg9UVIPUrrlSSHKayAXwzgFtzXLmSmUkc5t70rYbZxuwk9CrVPSUGZV7
JxPmqB+nVP7tIIPz3Y+51rcIlqq05DkG7CExunaOo4hxZtR1sk88cMpe3z2e+Ksq
87RF1r+r902u3BHhRy7/xTCjhfWsow+0Oou0QgGBrZO03pUSjJhSESInXZROJ1Er
9j6uXUFE9kJToovaEAjFnp3uyy8n+yx8ZuIzQ6DtT4FJnG8fNhabBqpnFb1huOcU
vOuBAGSJK0BKMbthPSLhtvuLUMWbZU4hfXrnLLrMUIgk3dfGf9Asx0KxF0mdxMtM
5xeyd36fWrc5Cr2dCtfZIAMmTL4co5DI37Q89jh22zgxsxq6wyeeheb2C3mkL5Sm
Hh4KOEgGp50fzndihF8LgdVZSY7dW/Ob5ZFRj1KRzXm1MlOT9gtsiGD6cdSA/GpE
a3txI7U+W6lRGj2r/Rn+aPSqph5UK9vWi6Zi2Clt1F4bhl81U0gTy5B7edpzjuSj
FMefeAgd+87gynPNFJefDNsF98FDJr2iAHIqE5eFX1ehT9M0QeCzV/WqHiq2+AZW
ZpOogvsOF8e8+Esp4rzU1IQEVe8kCRKEoOXTKEqt0wNG6/YvOoWCcmWNTSbp1eKE
eP/WZ/LFgQmwgYcln5VdufAobYjRevTp6rGir5zPSFD20rM0eJfPUuuqz2XoOH8e
zE66N9L2BB09ADtryXHAetWjYk0eDdKQv/NJScbBuJfj9BBcRbuPk9cw2gkesAgg
71Q037ppMTIkdFHY9+7Yu9WR+VQ7bneflALb8VWybGSipy0rmAVudcm4+XJiSeiv
ft7n7517Yn4nC/CkNo9VN8PzAVQqor0VK/mGhRE+V2+nmtVYaAU+Uz9NJrSiQkLj
3KPZnKr/iJbgtMd6VQxBmz59LktKtfOeiXSsxr9cbic4hSzsW7sPyvCJHzQaEh1+
4oYyaPPu/pWTAWZPbw24ZH50kCEIKrDrtcGdWKG7Obi50XfSZ5SSq3F08wuDwVgD
7hjElgmhj5Ydx1in7TPROKzi59joIpvtSq7n6M+e+yzMqJmbFpfrQBvJBm0luNQ/
2gjPJyMVDBPqSqwv5XtWZPqnMJ7NGpzbCLqHj/r28EIRjr1DhctJcQcWjIFSIAot
wSoevre/Gb2JmChR1Qq6HlMkUqQ3joSdHO1FDCvJPnxbrtUC3M1nk+yRy50PyUTR
wL8ZMSDVLPJY99Bi61yUy3xXoRz3VuKuvQY4HEvIQEd7W8uyvpLp5fCYgDHOeUyj
9kDBjmz65pIAZjfzHT9FRf2Bhgda8DvPpHq8gNIYC0NXbgucysyhzSqrx8XBVvuF
oaaiCmguswhwzpRBq2BZ8XSuQUaLP2W9fF1QUAp1m2T5MOaF0YJF3UIMnBdH4ZPS
UVA7rJdHYKvaLSHda9u2RoCoqAwXHsvvkh3k9zK2gYcf/VAKqAxmZ2ARj9nu4Dcm
vk6/5rNMO756tDJHNcyBst/z9UtZq90bEvYMG4RXXDQgIu1Mvadn6wtHZD52OdiU
if9A2TcL1EY95biVzdNyoISGo26K6Au7YFq7eAQgIzSjZhjyqU99LMW7AP6PnegA
A5tpD6FB8HNp1L/UFlw2QWXY+chFcS4TsvUr7PQo+254vaTMtPUr14H9epBNpOTJ
9SyfTxglY7Ofqdd0tt/vUl24M9zmSL3+C66TszK9i4oIyxHWXHn3r46A4gYw+IHD
heBFix+kkLzyycsIhmTLKjKethK69z4Hmuyrxi0M2T5qT+cXFaWqud7Jo3QN278X
/BqmZpFyq01qkhKzxUCW1ci/q/Z2zoz20K1rQKcz1yA9X6dxVn7JD3W2MxpFOnzH
bmJtBukVHDPXkeUQKyNSrfyNeZOawMlQGGEadu7f/uKYw+s2L491+aAKDULxF3+v
y0ylRE7i8ulKnO0QrKiZlu0YjlUY7pwuawGPZ7VQH/f7U+QuWy+A/CgGdfI6nEaY
bqPI/kct+7NfqxDYCRrhvxzITaPa9L66utC29C/QXcpAxOSPZ/0fMLmA1eU2Io4S
gDCUFH5s4KthPmgDUgETeB7VQnFF/7Bl7c6zUYNIGbQPVmH+L1eJ0Fsop79W88Zx
fDHdhIjvJp93RaBPV8VWxs82DOluSnUgq/H/lT2Vvoa8rHtfvvwZoQVv/jAIJzP1
7ppehgIyGlni8H8kkGHVUNdOblivD10l4oec2+rS8iG2eiuIQPLTazMYgtvQnMZT
oJyucE5uZMYq8rHLz+eHE+xIk6WyeKUU0j/imTlh4Df4mGedUDk1vDPoTJFY7wLD
asdaskN99j4y2Y4VIFvlNJ2ypI4jYjYpFSQO0cuXQu3+KxvHue8tG1efjbAFCdyh
+bzG7UBgAriSDa8YsxpWa+WzrjpdOT2gC/STRU4Xv2mApDxZw4+BRv5xC164m0sY
Qka6zy4IBm6MgGl1hJQ19o7klVSvpylkDaDWf/AmXrUdlr5Pv7jBctePjQ4ljfiY
pG3Qn9Er+Kl8xHv6r6afuJsidXWX5jKT11DxUiTR50fRe7ZJ5FWg1ivt191/ulK4
wfs1LWslWchCK0utdA0MLxkmcwpVSirX0FRG0nBjop9QGlPauEul2ATkd7i3pzhg
6KaSggVBJDc0kVimLQZAGkFy0fMqpH5zYPR0gYhX/uHj25VCNOrSD4FkqBvKICzy
YciLRopgY8DmxpC5mlAxkN5KxLw2WGTICIfH8TeUHCAJtWapCXXIGVvHJ42FsnLG
F2MWM+LQon94q1uPTllb2lxnd1x5eirMQyaNwstYXCFh81f1zDDYy8P34WKwz+qr
nIXXq27u1DQ8Dj0mLcm2/wC332Nt7EIoH5KfMzumBEtx+cJkJ8rmjujdsMsRAEqg
Tx9SyaKM70Iqo8wIdUHkjqZQmTzMAY3A4yMmeF+FamV9XcSdxe17hPwXcG5DBnIX
wkSyOL6cTpjPNzFaN9ISTiZiXHPHt1Q+6hUl1SZ6KMZ5j+1jZIplLdYx9VSi56f/
fNhRhETvbLS3tu+mdC7tq02nJKe5OX+7rOBDlFBKid2SBRaIIG7ZllEaf5iPO3gC
OcgEk2iiLt1gGP6ckIApGjRD9hoAVn8VSQEmLHXZght5HGBCVufn65QI7+E2ml9h
Wx7HBFjiNsYrvmYzWwfC8gdVbxMLKij1ckbvoVg1K1qOlAeyta1XDeiyT8EZsYMj
9GN5+VNSLAmHGyHFPTpYwzU1WhqNkR/D5sjmmP5WPrZY09TPoGPfrq4A8dIRAhDt
0VksFsCNqub4GsjHqyuLlm3BQVNTi6ycEkT6urI6RzFuLpihmw15di1GN9wa/1qR
MS+dwEfonK8r4G2/MPscJQsffB2hMuzktXmm/WAwt1zthtppKePVdH9X9TdhGO95
MqSGdeZ0wVKgNZr9phpobmlxnFR5ct6GS849sGiK2Uysa02kBdOBTBXovq3dPSuJ
eSmwgTgRpKUn4Pytjes09zk4bCCBjvzlhtnlojDBkRBczObrb/wvM7OGtlAC0Z15
m5sWhsuU4Y+iqxO3g2u9x34ZdgYp9naoIGljmNQ4Pfv4ECreXzbvyUHY0V0BfjWG
2rzazfkMJjUq86c27t96I3+dGs2gCxtxXd8B7moQ/5KHmO+k5s26u/mqxqjaSBjM
TcKUVLOeKwMIrNS0D9f4XTD1bQDyq/w4e6VOEWwLdDZnORDIt8ETldfkGF1JauZ8
0ncwyjJFi9E1TCsXH1FPSqfKLhSdVi/a/aPSkGm8zeJviQR7umPkNIRsQwEx/r4R
crDiRy9gRRUIOJiIGTQMZugz5kOAzuwXxNyX2TXaN1qvvBd8QaD2XG8b6figZk/z
KslcSZWWMI3/n83WIVIjheW/Sv1lMygFz2VCYnPx/fPnKjuWyMYhnM7+B/1rOQcq
rmFztYbmnjbpvybs1REVdhT7Px2SLwF43iNqvt5qHIUG4MUxtOsgY+HCD+p8ho7h
Zay41gMxI5Ey5guEuVILknpW+pcVyTu8htFJWCPhdVjUI2rAPaGgHH8fSRNhs7il
irnidE+2McYNzlQucNXMeHYBfvFhKqsp+1vgLFhtDe9cqbXZ1zVU7CnWrs8Hi8hC
GB2VXtMDBnugEK6G0IGp/FlX76v3kAcFecheT972d6vqbKE2irTfD85gttXieGyJ
cT/FG+rowkmXsZmxKX8xU16zMtld/DWZm6lsUNiiHoCMJfbUJC/xnJE2V639sb2h
rHNQm1+jbO5Ky499BEfG/US8hsYipBJsDWB1g5M349P5KMmY7XpPK8rx3d/moN6N
XMqhUt1HIYQu8xk0cn2tBdnb7qmL6Uv1yaK9IUY6Vab1yMwsR1mizNh2wQ1SoBYH
DP47V1QLzrXEOccZ9zVSHXsk4xism4A5/Xm0H5AV2z7QQ9zY2I/c0Qi/Ox4E6h3c
lOndKDx1Dpy13qrh7yWEVP/f/F3IKon0BRcaccla8DHrnmsCAIkYCOTK5BQHkviz
G+q0+2odhjTPssupsm55Xa03/kDqzJro4ap0gFbk11/ZK10VSoG1YQpAucagsYoI
7NghOF/Liv9PqHEgmIzWMyJ9EERIQ+ZLceTWOjMbiJt+5/scHEU3HLWPhnns9LbX
oy+bWrKFwfjXIA1CPvOnfWftZHIya7u1IQcoX9Nml43Apbz/1b0PohB47vWAse6b
nb2UMYEwGmLoq/+KM7x0zQRBHdbOiX63QihXB87nQrzqfWmlzY1Uf+4GtmOOu3ug
1ZxU5Xn2WL9spfxmykBd2vppIBc3d0C1ASNVLsiBLMh/M1waQwbSwcy1dLs5jesC
wCqSdANiRyfhy/weDdMKr8AMUJ4AQV+1H8OIwnj+8Zz0TxjQP9BCsGyX9zM/BUgS
mbaHrqpZZ5oC1wT4V5jAbXJDFQ2Ixznre0JZqhhiW6z+cZvb6iUHwAHo75M8TPc3
HHSTamdtLoSeHspmwWRsxfWGU++AHnE1r8QdEMJ29RIdLdcyPJbmfC6pQFm0NKuT
3qRxt5y98UZY7vgAjIKJ9c2IaDnNCD5ZciW+6pf4mQCnWsuVnf36LFNTXTHf3kEq
Mx5CZpkxKiTSWGDxEokJeZ5GHJtoYoZSkRF5WfxX9A5I1AXE53WqXvd9a7VUKDKA
ld3rrjJAOYIkDRopvBDDx8Inw9o8Oxf6GMRTdIJPz7BpY9TC5YtZaWGeWlochNNk
yKsHi67CAbjyvsQR/eLQvL8dVuppPOBBDnLcRZ92b+ZFBChLthzYCcmn9x/WuV/3
hqS/aPYp0rNYMXXelLPKXuIGt29GqcZlQry9/tiMFWFqzGCYnYWbcyoF/HvyKzBH
2DWUTttthniSGLjmd/ZkYXYc4/fi0IW6Uc0sn/5LH17MqZHgOcf070vW5uSlka2v
maAMnRgbRshEA3HuJweVSDh2e6JEaQtr84B7S7fMprrZpaa1LrqIRtBblns4FsKa
GfHAkx5G06U+qWKE1rQZuVobCTdL6lZBrsoZv204wQBpXSIBnq4BPMyT9mJ5UX6z
UnYOIYgHujZyQEt5x/pgLc4DXlTkoVCJT1KsoBWdTlR04+joAPF7J8rPET9fYFvR
BeXrtI37QJ5N2KvhMmhUTAuGNhf6Im4cQtTypgLvF2EMc81uDmcchF3bxCFCcG6Y
uJZYf6mtr2SqsMJuOExccRZ6dtOCKkXmMgVaQtK3p5pOg+csMlsqX0OsRd38vZA9
5Rw5zcExw3KaDAzVh9cIZke2B4dQX3AFtp/aJcWAaimfS+/JYE6FX7exzqaLBzgs
JYv2NfB9xmrEY089w+ZU7SZ57w5Pf8iRs+G2zCdQyio1vBvItqq/Zb45HFbUik3b
UpHuU6f0Kaz0Aaq22AfkcUeVTgP1YqbIsrePgfzGP4N8N6b6eebhYyrJWCt1Usdr
ec8pQ6tVilHQMVoceSInypjIs6ws9mo4ud+2JOkKW6ckQKVfZMGIaH0Y3wWQkyBW
dJ/z22SMHcKNu3BljJIzv7TgZAzCzllV2qFLJswUk4sFbb9q/LgQMxsoZcWSuNC8
pr5GbtOHarKZhD7LvhjqkfTb9PAVucUeovcUB0XqGFKHE1DD7aIoyzxFCt59EejX
Ztdvx5mvML5+HV0ZJszcGVZ4tGVO33b+ksmEK1r4mRlI76FEiN9jGd0TiNMtch9E
+aGAu88yUO5mXkWWIsu7Hrtcuvq3E0chzBl5VCy/oVZnjwl0DLcpPzVWyOssAHlL
pvLSc9uzhJkiiVs5j3Jx5JUyRVVAaRglmUYEIUFAX8kN55+3wK80PZPRO30K2xRw
sTLfwgYKFgganlhmId20xcXXlJPo2tG4O9E4j0fCsvgPJfohD0CbMxmZchUij6fw
/Y92yabX4N11Z87Q6Is6XkumQsmUiV1iomXbj5aEJc4bthBpATOBqi6EEu31SLtw
4wCyA7Vpi24QtegrXIZbsE7VMbc+NEDvX8wiylG5gwUfHc/caYK0QME3gvBU8Nqv
n6f6kQT8AwSjOr5DJnT+wZIMIMb+c7QACbvpJfPJ1BYN1bc/wKCcuD0F+aiuatEU
oBfTTwoCw+gufZmSRqswrjTV5JFNZEGUMBciSFSCubsNVR0gqjOyNs+BKukqPSDN
svaM1TOekKsTd4gPfN41Mphy0xJb1CQ2Ix+KMNgsKLFgJgfl5pWUXmL8TcHRGxE4
g/kO/2rv/GrWeeAX0bF672O5BzYJzDJhdk+NK5nywiRXqf6mZ7HG8TKETy/UCfnl
jOu+czNtGtAOsoHSUKwKuvACD+E3I2QSxAWFoxa7HoqUKaeBLh4xed04TezGVW5e
4v2OmJwgaFzVe6xvpwSmnipl3OSaoVvi+a6yP2e/WmgaSZbKeLi1C4VYh8/NGF6d
EhU2LH+fanZpNgdvqRsTr4bhzoODAX+qiNbmyO22HFZHFX9OnluPH+a4CJ1CqtDR
8/D05I9Wl8mbcfXXc4MzTolakbYyWN/x8g06U0EL8gVfxP+r3OucVMfCbJxfWoMr
SfZFB44qcTw9OdngAdMg0Wpmr0v+MbbfbZOp+llgLtXxkn5ii1WyaLv4OP8n5AR2
KExIIrNUX7SzooZoW7XveJt/CF8UF4QtXDGM+hVKJJidbzruVbumeUslmr2S7tXp
2d4oDRcWTzGiPn/px1g1kcPDq4r/Da9b9rR7R5iVkLh0GbtDmvcza11CZeCYIhqg
ztSU6fBA0ToRm9L1kN02vX2gwMYXVysC5KCxPiU5Vsi5EDC2V0abYlct1Ift3IET
s14ZYvuDNxmSi7fuQSZBXE/rvbd+nFvH0LXtSSYXCruQK1wtzFLvfr/GjrAxiQ15
6SemTjXhlyFTazGRg7mJmvW+wOjblgJpixCycGS5K96LnngaMmR57YlcVhcZgqMC
ZFgZzv2bvWfIHhu5G3z6/G54J7mizvqUHo/dk/PbgAb5X+nJe/OfgvMKBQCkoLvD
XpqdJnSzmGQazg89lISJQ+mOp356lf/zdHAL0hyad/QD8w/myYLzvRz7PM3a4k3F
kZpuu//SxA7McVWx6hCqPO5FKFE/qCwnqx2crbtWsmUdNV4BMxpSUIx6b9kgKGYf
POgUY//6Q5Dtf1tGEdq2mLNCKnrE3b/xN3UpNgNGzvmocdxhw38URPBg+3ePKeLr
O5LNPoEqbN1BtcVartIDRBDLvoYB5SALDJ/NlHwN8+ekSjdVZhWyWFXwS4JK0fXp
Pn9+mGKnyK9mXRQK+F8u/2QbasdspQm4o5dZT6RqIhBbIAl+Ccj60E1sLlQzz/oX
3cUeLSU7CDPm7e/gVL5yRargm4ZItEF+1mNyJyg6met0hkS65KdVT1y9TTWOln2l
EPATdU0bf9T28u8Raj8vCkqSVfsLVU+iyhFJJ+m8v4cjnHopY/9Ahl3pJp8LZkAM
XZCmDpgq/OjwghqRcaawsuCc827k6pGsTK/E5Gh7EEHzchu0JZtxyaal9k+LHbAe
UEl8NVAtV4JEZCATqRTryN7dkSvSCTjwu77V89z6SAAW1Cjs4YTKhdhZdi44DHk+
Q7rcEQb0JTNoy5PiPrRKR0Renk6DzEutI6hvT6U2zQ40WyCIO3Q2GH70w60jx2vD
UW1FYGiokBWWLFILI20tKe+Ah8gKLzVqSi2g16Mxu7wkesrWVdw2HyBhS+ul6xBe
S/7G34Ty3Fe6ejX2wHtWuH3BgodHG09zL0oKoaNMQmVjkY0zvXnBOeUrQSHJIP/G
AlH+H2H2sFASQTosXhrppp3uMKzHY2l7BGcU0XvOJQHCd79/iF0aQKIhrmPkD4Lo
gn8fha1ySaoLhsxoFBTRXSjEJoc2aTtNLXe10F1BES/9bEgVl5VUWnzSdmaavTSt
3+E2ZnMiBXUsp4rqFFv7uspzEdrQ6MWKLxm7dA1WFLLpItvS3lLWKqIGa6uQ5JIx
Q13qSE5Nyj23yDIhW93PzyMCHDMszahOKj1Gog/f72gIgq71FUtKNKRpsy7GAira
fOcjE65cW+3foapAOpaes8g3j4hRzcFvn8cOMndckhmfBTSmKpaVefhZbp9SePtb
bkXV0jgv0LUoKb0t1++5sjzogWwa433McYAzse1cnxwq3hgrF26VEzaL4k8JEbkk
Q8DAIXrKwP+8ol+UH3EqVIwo6PxjhArlKm96k+A36nPa0urSWNZuF39Nopcvct3d
hj0RUvYYdo85YLH6p9u7fZVQCZYaBXqLpM/LJNMwAQZmOK+gcJc9UqVkybdn886K
xF6VhivOd4i09dML++SgRBRZ/iH1Fl1lw3LUhsXu+rIJOQ3PqI3qohJEkzAkrw8r
g2XEki5l+0JOOxPkguenUwaM83MRMDYYjWhsY+X3I05shZIE61NmzrK7A4/T6HOA
lbahS4EwMh0wALnupLB+6rdW5xJYhHbVbUhyhAux687NUb2DA3itpjg7+RwRkBwK
fLcSJFgJeFRti7uFBD8cCb4KT8X7njX1qgzHsJSfQS+yeOYvwje8PNjGXDAbEXgj
/TT/AC/4KjvZh/IgCkrfIhtPbZ2Qxx2aaHiuZPUVGhlMQ89Hc02TT4g46/3RCyeQ
W/07CFDpmyalhjnZ6h69W0MwVbghxuZsiFpDe3YrJflarpZezjqsSV0jsl+gWkrY
DgBrOPKu58xK4qjigeoGdgtzSnrop/mcaG31YwkdTLKE9AcXvhrzNXjy2Y1Cilik
gwOUCGw9vMzp+9OrO5LdCfCHVlZl5UzKwlqb4rC4P5C5ZVVkk6itYgDdkUFzhCmD
Egvtpb2HR0HYeT9W1tAawwnctV6sH4e4dP969P7K6lpnPVaa5VG401smrNNts86h
s3TktYMLrefqMI4sx5XEQ8X4WHdzhmSH/VBMg5l5THnfJVxElmR+gjh/Byu4HSiL
vIA0izZWoQwEAJOt3y0hVGDOIhD3W2IemsW7sPPX0ymixP3fryUJC3oT/QbikJ1e
mRrdzHZ3d1BcitLzeO4HW7NI5+5NfCUcKFQYomeWlS9m8kyA3ZI6e0LhaG23o6Df
rOwsRLNX7mH0KaBNNteIMPbYlunPXMHIiSrOAldfsVSpcSi2Tg8aq45Eq6GA2cvz
dbVigiZUYs6Cj/UEg2qtKHJyNc0OA6YzeDw32Vlie9KE4PzVTXaOr00fa1ANyaUV
911grv4LHtIkNJb/zx8K7SYSFBq+oEAMuviQMt2weH1VzvGXQ7/uSXLxHM/S1jD5
FLvEp+QbpKBL1DGyJhstE4Iz7kMrhDTeFjPb+58w1IiiR9prO1drdQQLdZS8M0/1
vlVYDb4b4VU8xCQZnC/Ghm9Mdgz6br9O7WrdEpi0/QZK+lQmYJLCTkSjr26U8Ow0
9s2sBZT/jneediTRiQ/sH0q68qLvciPMHP/8IrNIAkGdCmGZDswADmiNcwL7Its7
M4Q88vik8c/uwimAY1uWIJ1A8sPCvQ2P7Z1xtFN5js98LwdX8rh84sGYe9QWo114
bERfYe9mQiOaEJOvIz685mMAFLaA2xGNpBNtDlvPV8BQjZ90DEIuoBkcGvguc9RF
DOIe4HqRzpgNLhKLzVk5lvbWptD/CInCPPwIwzqdWwkrztNQIgCDygGH7qNpOYxX
Cc2ehxj9YrrC8q7QWD7HlQtwAXo/9UuIfZaCHorPRwQKSKn7fKb77+aNnL5zMfjN
MAnzBBs81MeDCaQmCVcbBmFx+qQ5VmR9SnKj7oHPsisn5TxlInp+SYPo+4BZWFMS
3NNDie5xx7+DglxtiDWwjUYBa2LoCG0QBkI+ErCaOoIbWGcoHKR8SL+0cTnqvCnk
Qzhduq8ADBykNrLap7uIsysO7I3OU2w5qOYok67ZZLXtjTqZGGLOsu2QcQcalmTA
QVV8x9kVXsDUleFPufxkjoJyirEvDBWxQ4KWV8MZAIqBQB9axwL0W3eE8y2sf4Lj
vfDEuZ9HZuDPdRMoeQKptOYwLbiEBNuC5YRJvRAgnRPq7oFvdFgwaHDEd18gextM
aqmC1xTHR1MYMURYcZRPgj6xqhXItUtCivtGMwI4Cmcej46vY7yOK0ajSqqlX2xd
kDBy1Q52j//+Q4oBes+lvPIue24yJyr2YISK2RVpDHOXTXHAMt6z22iV2CpOpHc5
wNJPH8vypkAMa0qEHyzfePvn8z9G3237M+oUTshcpGhts+Sz+lZ5fkD6oEuc6Tx9
R8MbnWYk17UdVjcbk6oDySpKkajIEIYI1PNhewMe3W2jTYgy5CSWLXCo7TEjGunH
JEZHsB3lAoCvp4n2kU4XeFEmjjbteVVgZ5do796fm9BezgkIKaC6FBOHRqu0pq9g
x0n8Gcrg68R4NMiuY2PoKFP6fN9vQ/9TdKU/wNpJrGKNh7t31ph/6x91DPbeR9cE
02iWcNNATQinnWYbJdmdJCNJR3k+RAi9jUw6l2aIKCotGDeyJKGSBU8uu7CReuTc
BIryZaoamqzd+ycaEc/Sbp92xvdCFDZqNXk604znDCohXRrcP48t5aEBQFjXpqwe
vHFXD7iZ0Ug8MBxi9NC1v7f0yRJOhf3OzV6oM7FvRcTrMzZoZxi1ZPN1AsW6leiS
TU5vJXpZ4I/5fz9x+wSm2fGVF+vJkIHNdoAg0mdDl2WLwCMzDcJmgIYA3Mn4Yv50
ZgCQlbcCzFmSinXBAqj/XFdALzJwfnn5tsBeAfXkakd9BwsPA7pmCcZtxsC8T/r+
GFtH4YDfEmlj9q8WVQkUKyy1DldfjfyVqjvLO2Xeg5EmAGbBupK4qQBPvkNCwsPL
ntce3DEk/1TFAyJrc3WtwNyE6V4mVTD0K8oW9Pd+nOEf5CJHxTafpgm6bG/7f2vU
SaY+447CiqKSuzBWFT7zhj1sBhcrKB1mHusS0qhZMp8LOMRrl3bbR5KndUhFWerT
tUJZagyj3ozxUoIhezmNChMzaKmeMSgTMyWTIRKwQ4fJBzCYmqmuIW0WkJhcuxgj
tT037S4kMpcIT1b/8m9lQtgJSi72WLnl4yB2nHy6Vgb+phIy/3Vy16L+BgAtEuA6
opc/86PEDQjSsC+l6dlFaxY5WFU9eS3LV7tK1h86BSHzL15sndXlraltA6i12Pwd
dDRd30wjdpJa6JIq3+NuIJq8nsYDahhTn5lMTfsUUy36okqgnCOgrdfNKe9xeATd
dyiRyUNR6nCoSuuNDg0l4xe6BG/bP4Fndhy6AjQ6hFYnODZvaq4J15/l+S2/ZigZ
Qpsgz0T1Zqu6SvVEyS3YEyl6g9nPr75ISNQrQWFAPi84toiKrvPTTScRWv2buN3+
pUXtQRuFeQHojaHZboChv+gevef3Enhd2afoxNcqE5IApN/jfIbiOd/niaq25+v+
DpVqIbTfyoGzrQ8IlC99tz8cWMyYWLQtUb7WiNBjjH6VQwCMX3Kw4lape8FgRDUB
1wA6It5fB/gCcwzCOO/f0hIbHRgiTnZl16EN9V5poonZ8M7zCrHDHD/MhnepSHiK
fRADuafVTrsex/FLFmF6t0+95z3leFHfLSs+aGE9eAH1+INVbzlO/D0eqPkBf/nq
vcnYdgmdk34sUbRGIYSSWNdt27K5vU0psPxS/YWrES/Vi21k5LYAujSbqCVNN+KB
5JIOU/Vj8nXj0kNgditekJOpH28pk8xiEqfZ6YbzP0+viMckPcIjOdMtCjEYciHs
BRuMqda9jhEnEZZjOaZCHvpV/7tKbYejqLUSb4qsecL9HKN6YEabeLJ3z3ISn2zX
ldLh8qbqXQoR0C250fb0fuFovboexJzjBQqbqAELN7yx4fyu6MEeTTmE7H0P7SBs
AQNxAuKPlEz+1nmLbaLOcatbg6Z9oqNtmf0+fQFzyLsIW62N7wr4DQJ8KmtO1pfe
81TxRVmaeMvIphAu4QfKaRbsy161Ecnn47tQ7aUYbdDXg1fCt0abKk4NhdHui7Vt
bAVOw17Ct0ycO3YxzeJG+bgv6wnUWl5Mid+BIfIXKrJ4hfuyKDXQVJHCHkGOVViq
ClfkXr76nYg56x/Tlgb04z2laa4jlTZ833nlhUY7miGtI1asfjh4cyurq6oyTI1p
5g8ATMdLZjH2eQZjudcvjAjXuGTdjR4ZCVTciIpoVH+CwrH01jb0TeX5QQePMFXo
7SEd203xGZLbx3VRD55rjQbTr9Nsm5/WEUOdPnWm6QIUzr4dHnqx4gDoSWpNt36C
EVQSZZRfR/9oVOk5AJA5Oav0QCJets//n529A7vZTuIj8HDSyrZBhQnSO0/oNapD
wKLUVUtac6Nql9KsMpIE9yN8VUxYybiFscf2zEF3og+keIxjeQTxad3J8QPc2Hq0
Y7/gTqdAfhO/PnKIPahw50koBQvgEZI1qHp854OSWjrKnfW6QVFfTEtK1dXylSMz
Jixqi3P+Tv2AWZjA+fZuRIQmflv8jFKBq8gU3ctvvtDftgGtoR6JWTZRBysJpEqH
mx6wpJTdtmx4QYoXXsB/Oodkd8RX6qpUdR6ckWsvPAgT02Zz7pkZ0lYG3A/Pw+u+
wWJM2w46DQGGGopjmxeH71y8q+7ZsUK64G/MJac7fpdJhBmmNiiRf7SezWX/wepb
XpDlG0+MkXkMY8oFqnkUFwEnZ2qu2bIYdOxIGAe/ddCMwjK3e31AwWpdXD+6rV1O
QyZYU4/myGGpilXFofmZvWcmfOxeRWwbFTHsw48A7BfM/hsFOGm7nBTmHpn13SbV
8BjweO6c3SeruDzTcL4OzubfCaw+woIbP2en9Re8WYSH784kwX91CS9/cAT4e04u
gz2dEbldAqeLHyE79h/LWUo65rLh6Sr2s/4yMAAhqvPuYMf5tWejJlrMsRcOtY7G
uBb5doysQE9rQj0GpK/tzhed65vruvYc3WJEnHgSDb4kizIpZbMFx7cqsigmRM/A
zWiQlAp9blQ0qbjcMD8UtGkTyznJpPHT0t9rcbsKBB9jW9ynJt77BK+zPFbO64kp
wM+WZV+TjVyJM20hsyXG1YUx7bJY0B8DofBQvE67snae3HlRTA5Zki5reogdQY5R
/AYlyIPpLpurRyj8xKlnDiPewJtyKqBc9VboeCqD59fdjc2EoPCQzuHazTaRg4TW
g7mglNqgd+sygCyvQqmYIIgAQokwDHFpd4rOy5vtzDdgg9o9Bm7dHCuHjwPurDEF
Z7meLX0yejmev98iPKy0fXC3lfA+gECJOwRx7CUaZo+STmCOuubj8H1ZbqThdKQo
HmKzAahw/rtrgGKDl692qisHI/0fnrhTE/2HkE8DBYRLHa7LZXISTvtitG0hDvzH
o+cw2DF74xnceO3JnWDdCUaf4qaKDQcreNLYMG8ZhrTz4ESTUgCoqQu/NmiORQfV
AKpOmFhZ8Kwx+rOEmsGtSyYh2iVEoPvDL/bZWJ2BzJufAwTjyxkruK+e8k/0k1Le
VfxT2TsrGgX2Q3fm6nNdPAMkiCOjoghVHTAGINIHSHIpZhu5NNKKCHkE7e89YPru
FOG2xxF7RepWp3BxYs23IjEQqnOLKUddDADyNPzSiB4dgixQNVIps4nMr2famw1C
s0B/9Rc9cnh0597SoSLhSKkNpxrUJ+MNA9u5tOF17iGOwbpBuoPuIgJZlt83svOJ
luvLmyq08hyjydafDLMartylZNBp3CkRQThsN0u4ugXi48MMx70mITt12KV4aa+V
/Rx6905VqvDTS4dF90GdopHP7AGZdwyLcR94FbUYd0NNbYy/VjjPR6ofIqn+SGx6
2hRQUSPhuKeoGuCD9F7K7+O8s/GbQTK/488dtfiuIxqIRLOrbqNQGegn7KlBlDhM
lNnuwlVtM5Wx6DNn/EskuWS+QZIBP7/E6dPsaWPUjMoaIK8dn8wtsM2w2sLaq4NY
057t/vh0UFDVcKXK+++JPyubH7wSmBR9a/5jHdWY6yUWrg0tN280b+H5EJrcm58+
upemdXb27sINkUUT32z6fw4bpWP5MH40lVZkUSXM4KvdydXPKcKGTcKnK+jGiYJI
096YesqEO5FGOuOhRkykq+ffQCUZsG3ZnfjlacQaIdPwOGS2pgyWBOtCvGuUPFpQ
/XpeSeqTu2lDea2d5SORBDy3i10upO8ojoJlZswKC6hDnAtq0QdYKReJaFLE/jDN
zeywVTJxqOLU80rtFyLBbB/auI2yAbtPBuJUocqc+kHySZHch3xcb3r0OV+5N5eU
9jFEFK0SyoN4mOKkX/RPhm42gVX+8rte7CAWdXpkliqzqhgaJh+92a1wIpvkfWmY
ZXmsuyw9Seymve4gpSttsukb+N25JKeglQ/2Bjgi3coE41HRYtIutjo6+DHIP9ps
V5gF/NXLmBYLauhCe1xnUL+mTgWqPotgcE6hC4rAIf+5Y9i/XAfTY5tCmhOSI5Ny
AtXrWmmiVBey6NHcOdIfYs+3MpYDMQ131WzdKBwRe6uTqBqWa1JA+3FHHn2uPkFP
+0+0aH56nQBqpeydWYHahV+BU7JpjMDYPjNTp7JRtGGH6cGna0COEcFtkM1xp/sk
JQwas0C7Uv6WnkwA1hnvAPw58EAIGzfB13z7EaB3NTZqkjzFCMkTlhtxAUakjxt0
DTR3AE0rc6J5st6Zb3wWeJRzpdgIlHMWr3oAtUaw0uq8xUyB6KPtX9TfTaK2V4im
ert2dyLKc6qftjfPESE8XpZ12QZKNiUPw5tKuvMjZDK9ZFYY5p+333tYeEXwJ2pR
ixq3Xbu7lh+Qj3z/8+pULHDaaWVpxfybWl9Gp3aJliJBxLQC2uJH/5fJtwc/+mKq
GQhluiLg/uDqtjkhkKpBUuf4jXUyuuk5gjiZ3nNhjB4KInDghO0zGNhK/pD66J5C
gyTeTDg2zwqzUuTGO3re0GXeIvbHgbeSa/aPpoyIYBphpqAKIiiY4ZVFgT8UnUIe
jzVE/crwSHL6VxJOtbv5Z5RqIpn/C4T7ye9T1iKX94Ep1qbF6IfjN3E92MuiOT5+
21ZDkRe6/MRWSC0/WLGXLVfxlAObjisN99VGpnyDoOLSIQKGgfFVpfybQTqbMIlU
U+md2DxLaYGEOEyRrZedUbpT8MZf5Do7iQ7QPVSPeCMmLd/kFF3AOqCVx7nYmNpV
8hCSsyAMyM6Mzvohxbhx5YYhN8F4RC/rBQiZYtep15rGvod2HP9BEt9FCmxwprQB
I3azZMl/9WVAkBmCxQHhDm1an9ixycO1Hfer4m7dx50lu0g7KvL0bE6YxHR8MYVl
WPJyj5e9s+VwLmm5ECEtUFK+6VAKDqa65Nk46ZRN5NNZlff8l0oNw+1yeo0ygtw8
6lpW8ejrbq7r0vvLApBkLgICvdHmqftTA4Yiw9waCS1vjJ9h5ErCkID5bI1aAd8b
k3S93fvFZi2gHigQfEJCvqoH0lkof+ujfkUDbw3C5PQb6lzHrCgi7E0iTDQWdmYe
WT7062W+fzqF8ZpTuhS9hIogTcSeAwYQzz5C++MX54yVG5buc5/xSp4+yx0SsxgN
EhsVVJoaRin6rWfrCriszWKO9jT7SErNx24CNcaY7KkRpm/y3HnS8n+8PRw6pFM+
yxaEdWl67S0v0cr1NbLQpFB6i3bzpAEg8M7LxQtYOrDa+66MhR71QAZDKTM/Hyj5
zJ2NwjcnzhT6ViyIfB1zr2A9RA0bdPd0afXZIMSucJLs97sr7EBwwz1CFQPnwTMD
2cIycUF7v+sWQu0VIMu9yXMZ8+2Pg5GDEfR0LkI8qGEHrBW/7SGlO6D6P0W1uVJ4
MEftINM3PQoBDvTHc3Ua2pJBnEmROCftGKFgKSRgAvGy+kzIi8TUdCGhkhYNQd5m
ho8ZyDKhTYh6PVpOM9xcuskhSmvn+Rf+CCs+g+hHNxwzkxdAABsGQwsJXo5IfGuo
9GNUFtXKcYXyF1Ijh0QF2uDYqF653D9XknDGfTt3hUBKFyn7zRjAyGweJ6lCqJ5U
pA5ZLW0C4wv+gyn/7tgDYznXeuBjCNU/eQYiR9rCFZHbYt4lcbmJk0fdTLiMcq/8
+a7tFlT63Wd2zfYkFM/RUesd0nvdBObsYUcQqVNVrp3YF24ll+a59hQkElkYwT/x
nbFj8+rmW72LZUoTTPZ3eGhtvUvM5I53by0Xulk8NMbfMc3iJh6+hehrbHoRycfi
anTBywTD/iSuhKUkzwPZ0AmtEG/GkNHZGIA6StXfZ+PqYSihZmOs9mIjHmZRwrua
aGcevMLAaLY9bwwrvkc3wd61vJZRUb8DMe0huc0yxbS3i4Sc6XMrbOHaEAtWIfnS
Uz1x2Q38gUuOlMEqGKMglvffCpnvyK8rHxxGV/1vk7KlUrWjkaf31pNzm/jxRkU2
7ZB8s7C7vrtJ+jGKClewPT/4DhSg0Y0yN5dPDdec5TNVwGdXfAIOIltsHBY3QVF7
P9416VTkAeyCWy52wo0YAtg0NZBcA9V2MKsJrSuQbDEol5bJgxo2LRbBDaJuStjQ
0GEe5QyWbqUzSUyFhU1rif/X6qttF/uq7s2k1z5nR8btdDewVxEScBfg/MOTUXBV
Vb+f5mbvDhc3A83EIfAYYMRO0g3+MWAr1kKcY7XFsm7442YbB+rFt3Z974s77EjI
m1iIUX5ZSElv/rZ0PEvQ9ZoKs+51vC+8v9GdoAKR0A0NaTU3KSFmHKzE4VKiNJR9
cnXCbGFGT99kJbE59jYE4WiGpIS0QlwMEE5WwTn7G5+BxTlqJ8TKTjkRSrw2Shs3
xwVNd3f04VwTQkycfXz+WT5YNXu+ZNjSl4TL6bhak7eLDf+MyFILQQ9YSBW2cgfd
JKeHi+blVuUoIKA3p212fEW7ari9kd3Sy3e1RnMl1TFuPlCv+DOvzD6ICR8kY+Eq
BgW1UAX/p7VDEVwHZrJmeI6LyNMQDOW87eigUNpy/3d1ExvWB1QMrCOjU/3hUgrf
TrSfDQ6rgkpWQkYFp2bx8dYJR3yiZXlLhOFGjS3CAJ3EvndkzsgvVsM/66lfPc8K
QJaczdhtrsGokiyY+SDFGXCov6aK3syVqb+EBaow0CsQfa14I7AuiEB/EIs6HRP6
hJIXJhXq2KisZPVrY8PscxgHmwB5218EEEgdcSeIeNuITByPGhTtNuL0FB+2YgYH
V+caFa795x9WyKSnhMQRh3m7xBZWVXWntK9BkL1LsTG4fpA1F+hml6GgUQS6bA6P
T5jKiBUTdQQHr0QIu/tcJNaPGTm4RwFq9+P6bCp5YdfX0vJnjioOZSgnDNDBo50D
IFtZXVL+WOhA7aY0wVLH/B5yY234zJv0pfqYwFgqo3u3D4CdWRnoO6TD2QOxIh1/
nKk+4kLaBuXhzEDrfY05H1i1PAOuwspXJSdxoQzKDRW5oPW2GhUiuI8744WqR4Ae
5Co2rR/Dp2Wpr7Q074gSMMxZYsEJInt4tAZcHuhXoifMEA0j36i6ci0dfY4mW4eI
mQgtxcOq2fa8r71wwMEmuYFvRVGcZVbEOKiaC6eUvMAAQ2F3wnzqhZtdVkxb4ekM
JiSHdSH47Dstetz3YwPEdfCQ0MgDhpgg73EARuXl3sExwQeIjWqBEzyYjQi+SlCz
E5z86cEJB8l6PJlnOPf7DrM6AOUFCf+IgYDOvnh7bq8R7RwBfWj7nCiXOklbmXgI
54k69Og2/53wlJBUH1+thEYxqd+42nqTHv2XsNDhI+y49hOaHg5/uLOii/60gznv
I71hZP0fgJQpsWuYSJ5gNHLtKsq6jiDuM9GkGHy/R4YoTQVuyk3eQDarKlNrmX2M
MCLfq7fZ4EJaHsa1kYSo9J5si6Gv+dOReo6PJfSaoUU6eBqf2UbVxhSEYssmng6F
1x1+g+3XIOxS/bFkMfTwwkZ+8WvX9Yk8ph0iXFvx8wB4SPxUPh/likeyVV1KYLBS
0Gp3zjZdl3q/kLokIKcclWcyza2uIdjSVkSkJX6RDjs0YrRFLx0xcyCHTC1g3JMW
+CvYe4lOkSrYE+Q6l2QG3tlINDTaTBlbK1AjyU13ct8T+bR67wj5vz+XXVYfB1gW
oKFkBU/+i5GAtWC43RIp2sCUUJQ0Dtpn3P7gcTUdzp+HpURhMjfrsiXyX10TDUOE
LgeJNQR8YaCY3teUSxsLUcLD/n1lqnHmIpqRdqgNK/pfHfXy+d/WdlQ3j2WCdtR4
e6GFZzI0BlijmRFg40YNIa2MyQgHjwObKQR7k8yTrOC+oSJleCZqatpm2FHWWl0W
5tnNd49G+mRQA+h3uA2o3lh1SJ+MwJ5RiOGRXif8DHwvNj202Pc7x8e+pNW40oFm
Kv14RvuetRfd9NxiRIsupWY+Bo5JyWcGlZRXZn4axKuRUCB/jSHwU7lQvClHrwA9
NV3QZk21rc2CzPuky8ir3BVS+O/M/IVinNeFJgEs/VVddOMtapMghYEVVKkfePTw
nBgGVK1BCu7BSIvAAOtAWNDSaLxrp4OvM0iExXKh2qpYYcjL/yYkIJ6Qy1SvZVMc
k0klPkQCxtTvx4C6lIQJKGmA9QKpNkwMLQC0EV/dTJgEDyoqyipgrNFqL+lpZzjs
DGPilvXTTfWXlqcbzDGhwAysdOkR86EoyMCrhbBeDzsSyplOWmzsk39THqjrNyOD
7NXZ9caw217PAXWzLGuCCC5b4ux8HsSua4OHPkdiV0jbDY/VjPfdAMDE6VMuR3w/
reN+W9hrAUxxOG5EkJh2fIFoI5MkMpg7iQhO9h19rxuHTg7Af71w4eSULopwxA/o
PZr8SRFpHHw/p5vM+fu0Ix3LJSb97irc7wdMTadJOqCY+i00gWTuIh4h+Lb03cn3
zkbWQcxLf8ZwW0wAFdF9xZMRgZemRB6zsj/SlmEoQ7CQvbBgRjhzykt3CESDmq1S
hAgygyibnpepyNnbq+aKHpQjNLOm9TcO2N7Yvvb/cjVx4rqVA1GHsYQ/n4Qp7UtZ
drmhPJPOiM4edVjGa3Ou3acgGMJYN00jv4EFFJN/0l92YBczswT890ZD8jrh9V3B
rZWC4G8gcht47gmXtku51kvKcLpmmRWXFZkxv2L54SvvCB0dSODQqbTxern8c5p1
xUXAQTG5LUa2ulLbXEm+i1aQLmEO76Y8PlNk+WNalNMhQgaR3aPyv74ZMp/QTSrP
8girf1bTyNk5L1EEuqyA8/aZwzN45XcsHH5pU5u06o8FkQrr7LpVGsR1A+qNFgWI
sAMYee/Kw9A2622+2qouV5hGiYSxE5f7xTZeYr1TtyxwezAYlf3/gKFbUgp9BEcb
8fgMnsrIBagxxqY7F97KKgiEKgG8BG9ARw9c406Rc9Ncgs28RZrAIyWT6KFSYN+N
p0Wbb/iqp22WX0my8r7sbZXbiAayZyHj4ufg59E7/tmQFkGDWPbLCKnUK4JskJBw
cT9QpVFxRpgQWSh6GKSlJBlTGEGz9ydtXE7XG6u7pgphfV36tsJd2hER4OQ5OQXi
z9e5GVtTGTnguZQnUefjitsnJz2NJ2IEo4wh9KCIvxmqdqAEP8IAA8oHAyS/h4Uc
8NL1NsWBjunOqmdhTL5dDwHrWWBuAQsX8FJesvmIpkZgOYtc14IwshT9uB7s4he6
ODKLQTL42JhX4WGFW8ej3ez7C8wn0iAo6FFX7CFIFOZSsO9STTpGIgyBIEqr3KTR
3g8p6dlQQUke385X2z2w9fo0golkDeZ5PbmeKcKGf+9OCMLJ1tBA1aOUqlnmLRix
mkhjoC6lmFXAymJqhxPZ3teZd/beORGR7iwnaTLD/DIWwAzIJvWO2CtEUScwlwGG
fW7ThofTvQMqjQkGWL1sJ6pPgt278pkSOfaYBe3wMh5boEzZdxUenu/m0lLXitCc
Hoi4gos7369zht+aRY+uwtQy8taYfEVHL6l8YaWLlSjZIJk5yPRHaIjhmO3XyVq8
/Tt1WZeRtLTzSSlq2ssHVkgf4N9NvvJon4ZpnU0SCHIRuffIx0GvptWaVPbJntKb
GaA4X8atmIuT+cUcWdfFNNMGBYEcelgL9c9dABviYxeMhTR8tjmr1YNdsl3/3SRl
6RfaQ9otRYxTkaMfBqXh8xWJpVFLW3lSUnPDuhR3wFgMz7FBeSKww+0mja2z7API
qcUhrJ+dGbYnMj2062LntLe63HrO+X8+FhDcdH85Oye5OVdD1eHFdk/mHtU7ZqE/
QveyyoRJ1MFKt2wHvmzhiVFObMO8SFBIkpYxETxXh3eEMutvlNzu7r+kE2Kbyc0L
9hAfHbYq63SgHpwO+av4DEPfjfcQitjoM4iU3/1ANNzc6H7lZjGzDZI8ApiHKBFt
dMmrtSe6tjRyjVqZ3R4tftc2K/dbGvdZO3SUYD444eTvRsGz7CHYs9TGylPzfnOQ
OA05MkLdk7mSUmpCBOb7OzqWg3r7EENHX7geEwwe0ySCc53I+64dY/Kps+9csT9D
6IgqiJMLx3fVpUA6FHGRwl2vNf3cY47fdm87KpYJPEqRZvbd1wf7JM7l+6x/7cEm
KLn8rX+v/GIeaR559Q/B77m5LN2grdksQ9AeBVX+SJPB6UEl6O4RHIbn2Q094ZKK
msqf8bFfT7CvYC2xx4eWtg98oTks8TZuqqrI+drJLXeHzEPfh4kNrNvkuK3EijLK
hpQx5FNOF2zzLr3rLsO4I6G1rBcT3IzBSQHvz53iZHWL5F5AHxdTWkQKk/sRn8X+
JTW98/0MEEcKyEiQVEdy7Vggnsx9VmlXXmnhI3JG8SG4Oiss7MqV5yI11Y14G3Zf
SQbbux7dPywl2hBuwmC55xmtnwFbY6pRCB2GECzddOEupE3wZNDeXUA0cFF5oEN+
4XymLradTsOJPK8PPx4DmaOtq66Vfd5J6Hw10R50WyyOLH89ohbTLWVbSrk46ira
M8o3TyZTzZBAPNed239Uv+n7OrSWnfD4d+chi7y/A/W6A88lLXjOs85aJneESlcv
enVCjOU9GN66abX4qZ0/1f+UNTUdCsJCPKoiHlYCCMdXRUwky8QY6EX8QmomH7jY
i/Yaa48FvSoNQ7y59Xh3v4ShqSwWYd5stJNgGBeW3LBUBblQdJU1qjTwnWUbAxoZ
COI95MJjcluZcbIMin55h9bsPfd7VrLsq0TvC72km0KJ4yZTfj+AmBP5JrjUs2D7
e6aqIPliT226gH2stEOtNZJj94McnmdcpyEk8V1oNJkSXut/4td5dPsi2DIJdrlZ
fY90Kpsx42NS/Huo1beLDlrv8fwHUwYQPETFeyU0rhmdJsloNMmdcBeuhFkYDmxN
x1fVg6CTM0nAreA38uUKuXldKJImxhqfhHdGkpCUU+mF0qpUrWKUmOoikescCG8Q
fYQZT94I9W0kC3CsbMxgHH5y/c/BzEuZ1vQSZRw1EAt4kPwUsaV1JPkCRxyibrov
I2FA6OM9MC0Tg+Qouo4VZkT3DO4IIMIbIdWVUpJbBwGztWviY3r61RYB4LIYji9d
IYwTRF1/Kn+3QSHrQP/NqcJk8fTybNOVnOO6hpsLR5dQ0xiYbeA1dY7e/WJTb1jf
OXwBC6BVPUMSRdIue8/wa7uk/EtYRdE+K9TjVUKsI1cVsb6cB/oFVsW1Dx1I/+Pm
wJQei2hc8gCl0hh2Xe1SYZG8PXlpC4GXnCEqZ3xp0tChORDuudIWZSk4bvvGob5Z
FKtYMZoypGN7fyKBsez737rydhtTIWuyk06Cvfo4yGVLAiadkkMSqXGneW18dCOk
HrzaguKwrp45y4CagDhu9CGHwWCJftsSpS0SUwT9dtZtrQT+5zipDTE1SubMvlVk
15scxj0qO7ltvIAgT5oI7FvViMAcis91IwKL8GO4aYmkN9RmQU1KLFMNHPD1zbkv
/WojvKLyTnqOw4wMq3Huo61pCaoX/yleYZdFBl3/l4y05vwfanv8QkXDEEg1OTlv
9mRN3/x/cXFVKEi6oradzTS/FKT1Lhlj6Lb0/CWOrG2B3dmzAdl9s95XfQH0bY7u
Sh/40PIJ9vMxsW+T2qa4VER+DWRLE3vFk22bfmQxM7xltf1cNtklOTwe7E59ulBp
jRrsWTAi/Rt4fQ0UQyWoI+QuA6CIxsVY88zJclh6q0FN7fNAAbi2JEVPN1oRoU8c
MlmgwfCyZGQV+ojve/kRIrL6SUrJMVR5LYaF8HHkIaXzsFS/yfjX7bq9AELSU8Xz
k0OpM1PQMu7bHQi1WPwjj7QvhG26m26iNkjLAYtA1qezwTinnMgK1kxVSD8bk0To
StDpRp28QIGH+9Mx6v3A/6dW9+STGiso8HBboLnogYHP3aXypB1ibFvxHcsWcuZA
lnM4YkIsN6AmZ5tjLpkIsA1t47NnKfRTRPSOumkpFtEE8rC4JENSwKTpH+oxjv4p
vMU767eE6ZRFKUcQNGiHFU1WOttqPIlwpFemIp0FbVy0V6TPTVgOflmYXi4od2RK
15Hkr004zlbP5+EXlS1Aw7ZXO6rnxfX1vGgeoSl5KzjRAIXVjla2ih6bkL7VxorE
OR7wyK8/i6RaWWwCC7yhbuooiSUeRqnvHmGRgUltQEn19c1NORGrrrwYwvFCwgqx
d6eSNnL/FbqeeeisYb/1XOhtSb7I5SiroYLcLfjkmTXgUdhpewDSNS21oy99AqwC
zKtK7dcW7X+FPYfZsbMbm5Augh8U/lLiZ7PD7YIA/X1fAjj06U1LPaMryy5N9wWm
XcUmIbOvp9M7MDL5c48iJbx2gnqpmtqIjn5EO/yc5wnvnH/rYI6fGChP5OVxNROe
OeAD/DYGJum4iN+PLBDLj5webCF96IDZ5TT82CXfaQbW/6rWj+Eqplj3JisZvQST
xyMCSqA6MG1b4kam4VZ4yM4UAkCglrQYh63/vo+sl8Ahc5ll7Bkf11+duIPDMtzJ
TpzGsjUmBZmfIunwebpaV+7dFPkJ0ltPup/Crg0oX3YYw/mj/phjtKxn00aCKurx
Z8JkiYHJfBsxSyialLVSpkATpKewTM/cl7iyt7GbPqCg3B16ENNM/9TOTHpHNX2N
HMNQzXTeIZxMkVznTVGf2KPQtA5/Z3xJktMWcR42CF7bLcObUcw5B7UwTM5mClna
rztVhsUbGdIWIfBwEi3dOYYDF8S4kuFvwvYcAOghhT6IA578CkH1c2ngjw6E8Zi9
kT/jrTSaGlY8LU8J/YSpBR9FI/pScFCio8dpEPKxeHUD2Nd/PahenPWxNYxpst4g
Q8McKuztFeOB3BoqLtZeeBIVCatRZfTPmkhP5NCkBp1Yx4NEiWTtj8CoEJIEOzoX
Q9hGwZInfB4evnfOLqzdV4JA5IgAXGUFrJTMouQ2VuaGfu0hAVnIatouEgWLd6iy
+nox66rNsVvAHMuG5hafZ7m+FeiItCUGco2jn3icAR1Y6DMZtAlrAruZ3JSLaK2s
yiJ9rGHtJoMTz2jhKw4QuRJFgCjPwiPWW3veLzogfBKlGofeCUG1tiJZvkwHhPEx
7H+GnAcPzNjZ99hKaggzbPiqu0glUBzuiC0ljTAN3EKdqjmh85Cb+RUQeWtocEAj
BnqSyJnT/tSDBMY6sGSypt6VIil3Ek02NfMZOWvVeL+Y9mJ5tH/k79ZmSzfJxxAo
0I3NFonyg/u3WtW4rx8ZgoNXwKPTeosIiP0YiroCywfq4qgYYfWxPk2IGF/kR+PD
wTnXLuM6QOhCKK3Py3tCieyK1LuAK/LpPlu8f2ZZFdI9hs/gbjst8P9xYHm4Lh2z
Sk69ZYi1S8YAKyb6swPWc+0h2GJq8UYMOtQic77Y9ujpBtd474QEUOD/XtIWZq1p
+mkpEkS85ucHFcKFUGA7MF8A/jbcHVeqhhXonirNWhKuddxkzuuXNFXRlYOkajLZ
`pragma protect end_protected
