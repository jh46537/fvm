��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm����질�95J{۠�zf���J:d4�d2r�&V������n&��s��N��H��@1�`>�e�dq��kz�s۽���-g~O�-	14���4����D�s��P��y�P��l37�;��s<�>�B/���G�㽥P�%�N�ϙG˟@1hˣ>�]�Ă�K%�j��{�D�"�Ls�s�A�� ҡ�CǼgYI���n�9x���$Ҁ���V�\��f��-�87_]*j	e*`5�Mu��E�GEΈ-�$r[�[H���'ܑ�=��_%~�z�u��֟�Gb�C|n�V�v��W*jm.�%<����9�n ���e
�p��ƍ%�n$-�d����8[g	6�e��;���*�l4�9�{�%k�l�W6��df��c��Ob����--J]�A�:;O_��r�ʂO�T�yl�RhB��d����y���G�9N�0�o�o�}~т�� ��&2T0Br�z�K,z	;A��J!$��<��x��>kkx9tsKTD�릲���ζ~����`���3~K��NQ� �N�d��
ёo��Zs�}�C��84��g��ŖBn0���ɁLy�%<�Ҵ� �S:�]t�<��m�?:�P�f��q������B��6f�c5��s9���"�fa�I���j����ё�;&ө� ��<�S1�n@���sd&�<�;4��R�A���Y�;�y��p�ٴ����g��z~��m8Qj��I��s��7��2)j}M�,`��$j�k�Z��p�������d��/�v� 4��7r��ۡ7]i@��O��V��Z�� z�J$j�2��,>�1� �[���#��uÇj�\0U�9�7n�1�F����=��|L��ƛ"}��޽7�ԏn#d��o�Ǿ+�)$��o��n��,[�8?Js7�p=P�N��4a3�
��<*�Y6�.W�i��n�$���.|�7y�1�T�0�>��\H�5�������?l��S�iH#�AL�ŗ�@μtV^���� <Ҽi��n�D�?bË�uP������0�;�S���(χ�,���6z�
s38b��?�b	���7t�/��㮗���e�݄r����&���I�:vl��ait^2U�����r��N�B���Z���1�<y���H:�rײk�U�M}�_ �ϒP�E4H�`]N�5w}{
+�� St�b&���l_�vV�}�m��Y�9z�k�H��t�ez�Z�e�Q��WD������@k���߷���M�5h��:ΰ#�'@W�\d�n�pU	�r����`���ma�����\���`tB2k($����-�.����՛���9����G�8#����6�y�l6`�25;&��m�	3�������^�i�_�[H�y��k+�JY��&*�[i����)�_�m�
ܿ��ʷM3��xw�v�.׸r�m#�� do�|��N'p���6.�Ei��&z<�/{�a��gn:4M��5+&���`u�"��n m����?���-��('�Ͻ]�� *��`�^���K�m�ӽ���yP�(^F�O�-����~��MϤ�wSF,��'f��!��/���^�P����-�bq��rz]�x�O,]ݼ��)��U�z�O{����\���[-��`�X`�n/$�0|�;3#��L0�~�QU689M|�`���!´.ɘ�4U�֭@�TF�[�Ŧ��q'q;�a��lO���ϭ	{�e@�[��'3�=av���c�܄��Qç^(�z�k�a�^-���N3DE'Ɏ�EA�4 0�J�@0Ƙ⏛��PM�nADx<���-����a���J�������K)�#^��vq�j�W�A]�z1�&��գk4��j��j*�&�;�MF�r�zkUz���4�:?>Gkm�p[�v�ƍI�۫�o8y���OS�5��C�j�����yÇ�9z�����3,	�ۖ9�����ŵju��5'q
U8`ϊ�5j�F�r!&�!�W����{}�R[cU�WL�m4��7�/k�Z��!�͐�z�ūJ46v��U�{�fd�c�ӀJHG���`b�$Aǲ � L���	� C	�):��3�LR�Š��'do����#�]�t����LXŖ�<��Etʮ��b�������"�n��V�������=f2���-]��P��$U�":�
;�G��'���ϸ�wM�R���y�lة��X�{�9
#Nc���</T��R	ۍ��h�%Z��D���v��d�h16lXkR�x��N��:x҂�OӬ�l�]k6a���2x��S�t[yΜ���q�^G��H\4
�G��R��{�.D>=ld9�CP�~8v�^���G�N����w��m(q�?Ή�n`#�m8�.c[��Q>>��ͤ�\�˵��d���2��k����J��T65f1��!b��kMFR���v���B�V�-��G/]�e_���hsr!�Zj�X�;a��"�d@V�#�d�͡�(�!� ���q�+�>�_��SY:缾�G�`)Ve{f?]��`nZ�M�EZtЏ����:p|-X��4��s�z�,ٌd0���ÖG�Ф��e�{�?ꌶ��Iq����.7�(� �U�
)����`<�|��el,z. ���lu�I�;Ȼ�A���R��+v;mG��s���J�Hک��sQG�c��	^��ۚg���ꖼYɩ��&|�%�e ��ޛ���b��i�JPK�b���+J�ao[=�5�{��ҭ\-H^�Q���'�}	�{�v�{s	'�߅��珬���A "`�|̯��|R��N��.I4�`�3�li�2�t\(����L��A�oV�U�:S=�� �����p�eT���Ry�,�ܔ��@�/>"9�~� (،nB0"�rFG���-����J�ѡ���ô�}~I�<��&��Ǎ�Nd���pU(ҟ�4"YϢ?o>�����}���Q��b�BI�4A%���|\�x쐑�3����o!Cƀ撬2ć��w~`��I�4��]��Q�e�A�ir#'i�������E�Ʉ���򾷰trO�u�FgK��fMצk�z
�]�E����pmT�iD(�:sQj�bֱݪ6˰|H���@��a�mEl"��꾆�IX��^��ۧ�\�f�Q��B�bVj��2=�l�O����5.Y'WG�h�n|�r�[�F�s��j��_F�h>���r�0���qNF-+��is�!N�]���/b���W�Ub�ɍ�r��i�%q�d�n���h*t�	��UNB��\��X��ʡpǮ<Q���u��ć�<�ϼ��x�9��^�y�c=rx厭ĕ��;�amP�
B�M� G_95��9@ς1|��E�"ҁ@������Ks$,��s/�R1�7Y��S��g�FA��=$$��A$������ �\����|[��G��K��]���^��N�}�}���,R��]ڬ�>�8�+��ze� ����	����!1z>L����s�t����;���3pS�ì�ۤ��	�S�H��4���Q�as�聐�ۘ�s��������61�PIv`h���yg���G��Y�0�g�ɷ3s�����cv6蕥�7�r���ڸ]<��"������q�ҷ�B��k�Bt�T@��i[ô�M&�+3^��&t�EY�wa^������^��>���`��86�c��E��s����4��&`�HЫR�C5��ֱ`eۗ���!+k%������GHBBWNFx�Q�������'�퓯���t:���)^���v�u�Ni�"��z�6�3#<��W�+��J/�s-�ǔMt���r���'s���xȯ�-̭]7�$��RQ�V�ּ��RE�ݵI�w�L�I�2W5��p���G��]_�(^()�R��q�_���������e�_f�� � `�۷���2��sW��Y�b]4�@��BJ9�R���,q+z��m�V�q�G3 Kr|�G3~��N%�~�I��c��o+�&l_9S��H#!�������{v9W��Y�*����8$3��+��,z��lT�����A�	�9����L�9�hW�@d�Sy�d�i%���>�ǵ�vċ�C�\�3=�ڞ�lʇ���:�~��aH��\�N�!OHgX)O��*t�3E�K䍰ȼ�C���r����XV�gS����P��i�9�ZG��p�x�H+�Nך��gRu��JA��<�������o�`q>�rV�
%:�S?X�tx��>4��I��E��<$G#�J ��!�|1�W;�݀O��8��fN����ٴz=Ͻ�w���n݂�\�����q�{Z�t�_I&0���mn����������r�s__T;�$o�h��~z@Fr�W{�����4�FOM�̗iQ~HL�œ&0����Y�Ee[�Ώ)l��?ÿ��S �еr��Ȥ����?�N=Å�M"�;�B��W�:J>�m�ܚ���R�Q�|����e�d=��(3��L�=��x�(�J�$XlC ����i���)�}#�+9����ki����j=�}'�(�6|���)H\�Pᐷ���Gި�vʹ2��Q��}�dT�u����9�y���pµ "��_�S[u���;LNT,r}Y6XQ�"bs?�-%���.�L?�*�����gۚ���1���-%������OŪ���T#��YG�XO�w�t��OW{�e�Y̓�uU���Wv2ɏ�2�joW����"mR���ʹM��݁��voI�	:���\�����m�������ե�J\m��P"�X?�AB�Nk��:]�h�5و������L�W��/��\�#��rq�o�ˇ6vnI�?�pa	0���|@ ��-��<,3[ݜ<�>�G�9��<$9�M��1�Xě@x=��dI�<�(S�T1����+�$�	�B؏�]��F��-50���s�-�b�n+'�h��֩b0���(�:���w�*���lV�� Ӏ�9,����M����Ȕjb�����j��� M��g�0�g��\G�a&����y=f�(���M1�9����J��+�2N5A�x\w�<!��ioDV�o��0vb�Կ��ُ��rM�_�Wo&ۧ�W���6Hl3}yC���$-kp�i����7��~������ �@���Y�q�A�2�á�;d�ͮ~����dڔz�̦�P����w��ǯ�~&Ւu&����gaNM��f���\#1-�R�/y!�쾦����HNA��	e�m�����VՓH��x���XRM� ��={H��i#��?i�b>��a��ψ��)���J�4*PH1�9��YT��W��na7�/ɟ4�u�a� (ϗZQ(�r�ER�.��	xV�L��	�������I��هH�������ܳ՞���N_�랱� ߆� ���p�����h(@U :y�dH�������wЫ1x�ʜ<S�N'Ƥw�gV8��r�"j {�VRBў�\����Kv�3[*��7xDF$�@:(x�����3=4J�[�.Uiՠ1����	�L@�TI�y�3q���v����h�S�Ye���b�F:�!(E�e$M�6`�x,f�������X)gq�/~6�Hy|�o��yG��.�za%˲�X����ðЋ�k8T\�`4u���'��:Fp���H�
U}��|S"��99���.p�\:a������Zd�g9 �1D������y���,q=���z�Р�a����Ż������:�*jL�-͹Ǜo�(@ ..���>��������?�{h������1��ɜ�0_Mo��6U���%�9ԥ|x��l���f-���s��]HHF� ^�NeB��0��a$�_����o�[~�nc�YᅝM�g�lh� d /��#�}wN���z��*���ef���Ҷk�<�z/�*u�	;��r$J�ΛjZ]�5�}`�"p`(e��0��'_���F�OO����ˈ�3:�F��g�̀nݣv� 0�9;"��S�8��,��:�(����ʒJɂ4#/Դ|�ŷ��l��Q����\ݟ��a�X����p^V���F�kG��]�t�߾�!�E�>&/C��v43�	�S��C�B)*�ߌ����C�d��
T�ADB�]����4-�g9�.M2�O|��C�?�"���Iy��I� {�$�� �5�/��rT�@o'�:�D�d��'�S��ԗ`�~��tHJ�Q8�N���D����s�ArҫH�S�W�Nj��]F���_;]L�JJa�6��p���r�cŭq6�'������?�%�T���$x�>z1>T�L����y�I�ܟBh��b���YsM��?؛Vmo�Q�%�a~w�����I�g�0X[ ZU���l��%�~�)@ݶ���Y�6��Ie�U ���zxf��@0KX� �j�F��~.��������ugfV��P�҈���r� #j}`�^lp:"�wa�í� A����~��+���r�1xǤ��X����D����q����*��|�#o`Wb���8ਝ꾌�;D��\�"R�,�ד�������{nmJ@���Kz*�{�Q�(��}���
rޡ����U(�6��Bx���i��  ܝk"��� Քw�~�{�^
&��Y���:m5ܬ"\�tD.��X���p�j�J�9��dX��L*�㘪C���#/n��C��7��Q
�-��q-��jk/H-Q�����cby�`B�K���Ӈx�>)%���v Z3�?]�5��� ��$T���y�utI�*O��^˾�Udc�O�+W���G��}l%8���2��MX����H��6��p�� %	3s���pb;�E�!(�d�F�Vv\��H�2g��7���(~�^���pȿ�ם�0�N(5�} �b%��������omل=����F�<^��:���&xڽ���;%B-�6r0R�H�4v7Y�d4G_M]`pq9.M�6)�G9�2��J0n�?�D�^K��v�fE4��'D�����a��0b-HHȣ��6�[mg0d���4�w�3ܥ�fܮj X6�l�
_s�!<��֦Q��_�q���Yka�iY��(�?�,�nc���oe2��2ݸ�t���� �Z�����Y#f���+��"\f���~1Kd}S�d��;�~�KX���gΪRU�Ã�6o�#LM��l���!��~�v:шGחM�̈�#�-x��ҠЃ��\�*j�ݙ��w����lm�D�$V�>�ǀ�`���O��^~��&��pQ:��2�Q��J���oVq�Fs��-��-b͆S������$���H�$����_O���C~ta��%�]-�N��?���5I0�(J�v\�����ȧ�gc ��^L?�cbؤ�-��
�z�`���t�v�����I���*�*<F�5��-6->�px*L��d��zs�9�udDa\�����X���8�|�O�:����~�@4c���Q�3-�F�@5�3���C[�<8Ǿ3��,��Z[�SEh�j�p$�6_ŝ<��g~\��dnP���6:�n��/�.!S�� s?�i4��tO��H�P��t���%�q}��>_d	�0� #��}Ѝ��JrݞT�N�	
E�Ir�`���7DD ��Ig�A�r�I�:,T+#��c�RoG�a���n�m��$��mZ�Φ��'L�{�cP�����<�6A��(ε(WL�{i0s��[��#-
�Q���Z��28T��Z��h�*2���t�.��9��aMblx�w�y[��br�3N�����ū�x+b8M��������4��+@u��rJ����	{�1L�5���Q� yJ�H
b� �`���>7%#'F�cX%ζ*�/ns:�:��9 �Ae��K_��Y[��+��z���`g�?��aq�c��n��$��Q�(�]a�t�'�t@�pj˝ԡs�y�bW�V\1߂g(g����Wb��#��a�������r�]:���v��ML���)�)�,1ciZ!�)�IC��=�t�G�7b;uY�&6�.���9�g�s�@\0�^V}Z[��	щj��F�U�T�P{�A~�Ry҃d7И��^ا�l<��UӪTۈuei�s"�[].%zcm�WR#7��:�̏�Ӝ@�?�O}y<b����Em'��=ˁ���8� HYR�ZW���XLVV�LO��͞���Jw_�E+cp/���ۛ;�,�a���\|�7B�ܧ�QtO�|E�*ʭ�ba��
"Sm���G��������]�V�*��7.ַ�_��ީ�OK����*�ݵ��Od*�ٛ��iO�$F8�(����.\[�����韖?'mp�N�����q�����:b�![n�J:E$����6���P�" ��H�Q�U��}z/l܁���N��)��Ɛ$AԽ;\g������X;ڢ�8��������pt����k�_Y�O�V��
q��M���h5�:2�cwQ�d>������[�����%��d���dw���>�E����W��F]
9k?��6��bhU�?�SQ�pV!	/Qg�*�q3kwL�|�*���.G���j:a���W8�;�69M��HG����(�e|joq!;U*��(�,��q|w�h�e����!���!�Sc�4f�B^ �芵��%��\T���-!��#�*<�_}j�AP�
�lᓾ�1�q��!G3c��yZ���g>���5�j�h�!�\���9Ū�M�>��ƫ��#k�N���p��d��&�%��#�Ϡ�E�352�[Դ�2�cn`ۈ����A�B2�a���)	��";:�y]�E��ej�ɂ-�z�`����[�]��5�B D �B���7l�~��Q��b-�]s���2F�;RJ |��YOŕ��bѦ�%vNh�r����g��A��qZS���釟K$�qe���&��c�	���L��Eٚ���@��Yu�D�����	�H_`�*|�APr2w���#� ҟcu0�2��d1�6cOql����s�"��'���}Σ@rao��q�I�\��z�!D)]�3��)��K�����*n��N��@�Ͳn�N���gd̍�P|����8�GWM�ڽ�,/�-4Hp�����JY�Ďַ����Czr��P����%���<b��M.�MQr��i��6�����pF�� $�`�Ba���Hv���^	L���7�b��T/��i\^���q�o�������&OF��3e��u�t<�5���T�w��O���oB��@t=ӚuM���>`�<���Ο�G(�*�+%r!9���j����Bs�y9���dk����5޶��@M^�-X�4�S��1�P���3�u[�'")ۜc$��������`����+�X��*]�*U���p���*C���X38?{�A��@G~p{���	���<d�� ��VX'׺��r�o�,Ƌ��є�SJ��S�w�/:�m됕Mul�ifO5���*�
�K�U=���z�� m�p�[�8�b�$B ��m�x�F����#�IYv$����*��}mU�g����6a����8��#O܊Qq0oŤ��D��@,'B���󯺼je�y>HNR��p�YT��m��[�3&x�\��KڗPE{R�I�o�9�� ��&ѓT$}�V��nG�w}�`�#�6p_����C��ֆm/�1����u��T�.]�2�JÒ#'�o��Ĳ9���iBC�[���[�A�ք�1��8>l��Բ|	�h��5���"FE�Si��E�M����?�w�,�M���n
Y���@5��*id��k��R�Xbd41d괩�5#����ԋgKj���([
,<"����4��.����䁛r��	z�X$4dH�ܩ���;8��.�x��\�r� ���N�G����w��^Im`$)~ߑ�:!f��l�U*���tyy!7c�6�6�Vc�˘~]8��_�?�~|t��b��K*�&�Ӷ�I�H�֕�SO��?F��u�~��`�O�6*r��$5$���^M/j�K�Ė.�M��Y�I��^n�w$��P�u���1�>�Ϧ��o�G�ߡd
<��H�"x{����Ȩ�����-ݻ[��!��޶�-�֍T��x�
��S�,<��nc{�a�ߥ�����#-�(L<���<���s�>Rh���<*���ՎXԮ#w��WIG_㹙��?�"d��j�8�A�92@�*X�ֿ���g��[��{PC��~��QY��u�3�>��~ml�E��۸m��#NO�l�c����Ԗ����ǡ��
hp���M�C3�M"\�I��3���?z���~��O��L%�2�-E����Kr�a�	t=�������S�Hj@������n�E���B�ذ��'!�b�a$8B��@%(f?�w9��� D�S�bV��^{����8�'P�!J��ͦ�,�eF3H�b�U�������BHg�k�ZH�&��>����/���X�	�C7ԁ���R%�ҳ��3x��ҾV��B�����|4��yx�c&��-Lw|i/�\9�Ȥ��� ��@,y%�(����A��8�Z���b�^!S�" �Lbl��������,���_M�Uܜ����:�Q�S7���Qw��	��\�_���%f��C��Rsύ�,[zG����
k�}	�0~b@��[C��΃HJ��K��y7ۖ����k�|�s�tL��L�?J� ��XtLa���s^k˱lTc��3��y��o��[���B�E�G��z�r7���'��s�ڮ6	:2}M	��ٺ28�,!a��qy��Q��x6&�����o�j$L�
���M�R��8�:�u�*��}`��Kn�T�7�6����9<�ڎ�$]&����Ӿ9G�! �n���ƍ�ڶ	�>g@,�r#�f��Ű1�\���߅�ݻt�����ໆ�V��J`o: a�/C�������%�%�[����	��1�(�b�V �Kl8`�2�}�T2�@�n�P?��� M>�k[�	�R"��F %N��9>�����X8>�f��hxѵ�\�y��H�ocÍ�II�O(� I�!\z�fѼ �#�@�ͼѴ�D� �-�\ɂ���wIw�(_3�Y����Ѵ�?�P:�ў���Ɋv�&��a�	�� N>���|���/;�z�=8�X R�Q���K�#a�����Ɔ�_��V��2&.F<��y���X��D$$��yԈ9��6���H���l?A/���$׎��cߔ?o�Yw��t�1�Z~W�؇+�뀣�?3�N^j�{����	��x��������+$�=�t<Ys�Uu�${�oXX��@����D-�?�I�0�.���c�����C�)���t�K�_�6��iE	(�M�ۊS��p��t}gS�C���3#�ݾ��gz�j�%�OH�m�zCa����B,bV2����A�ݓtƨ��A�*�:�*:��w_ǖ(����4�B#Ia,&�������.�F0�k� �Fq��m����dT$%i�hJ�Po>1r�`�
�\��'�D�1�?�
�gy����8�$&��� �ح.��ɯфY�#�vʮ�f:ǙI;C���.r>�B���l	/�jSK1�X��w"m��^=�����"�e�����t ��NkEI��XU ��^`P��yY:t01�aeKV��Ls]Y�_�u;��D��m���s��vb�܄�#��#�IT��-�m"-@�5נ���BΫ7R�.�^A(����>������Nò1��E>�`-Hg�p� �:�q!�l��g�͹/���/ei��Rj�[��׼�^�ޭ{�] *��ȅ��YS'�^��Ic�,��ؘ�����0͢;���:Dȟ)tIC��� H����2踧�{��T�I�"�-]���.�{�b��ҍ�m®#�UֆY��B� �up��]�����7�z���1��c=��s��I��u�4{B{�͗yd��yٰEDxǹ5����!M�m�*��o����4/ a�հʹ��ܗ�$�BZN�Z��|嬈S*�hA�@��}��ޑt�7r�D��dd��5�B	fˬ성C�P����f�D����w�VDc}sD۴'g,��%aA'`��TR��;&�ù�H�3���^�����F��9��U�����w�����qA�Y��v)�'SB���hJ�
3��ݞ���xO����Nn��D{�RUE��o}���`�j���Y��cڔ�M�������"o	X��]�I5Zs��ת�,����6ҊA���:�b�m�����!��<�_Ń�~C���w�L����7_0:Z�w>a{�E�p�Enii�zr�z�h�}N�j�+/3�)��T���!I[�th�+=M)zQ��?V�#oA=hb�T����g��m���ٺ�Mfb�����L�gm�9��$����S�??�A�W#�G�VR5����AQ4"m-���X��AaK@hW�Ԅ�5Y�S��N2�?�;���r,D�1K4�_�1GG"���G�7ɉt�k]&�6-�
�-�������X���%�H��S$�'d�ߴr��2[E\�X��>?f�5�"h_�
�X?m�#D����}A���^J"�]���j��o�5.[��<�UWNXu��T�d][�����{�aU1��_Y�>I�x��(��Sa_�󹍍��7u	�G	>�W�� �FĽ2n!o��ue5�(}B�����Nh��7���x�:)����	.����OT��ͦ�;����:ۆ��+��a�&Ӌ�W����J�
Ș�3�N�����B��+��n:Q0nڀ�N��@,��<��W5$&�G\L���@��.�������������ݣ,�)�f^�W����9Ǒ������q�7���߱!�#j9[D�lU3��t���`��FP� �.�a��Bt
�[�﷓�;h��N8�<>E���2J���q�MR��j^"���L��"iy�O <�����wQc��w��9]׾>�(�ۆ������!M�,L6���Vڏ)-F�k�_��f3q��3�p}�&����AG�:�G�nj�|KkTn--B}����@�A���k����ǠqkG���ٜ���j��'�b�ϓ'��*fb���	FAܯ��2<Z'�v��ڗμ �e����L������*���z�P��$[�t�4���������qDP�h5~O0]U���	S�:f���U�l��Ш�	�U�����.9�]����,�!^���Y����*�\��H/sB���87��f�S�w�_���~�o�),���Ą[ لB�j��,�;��q&G�+��1;�P�:P���� h�D�X2Ųb����36m��LY�_7���E��$+a
��B���I�d[������Ru�T��Z��<��R��{�����V�����	\�']*��3���L2a��9{gb Gë��J9���ob�p� 
�3� ����͝����]R{d35��a$���M���º�.�L2��Y�-��/N�(�b?yK��,J!�2S���T�!�\{>e�kd+�@����Nԭ���㤟۩3@x�>�)X9��QabHUU��F2�R���/�83��yEc��93���}-Y0���M������3�S�	HD)�Q�)0Z��Ʒ�/@�|�#���y�?����+���*�Y��!��q���S�ϋ(7�^h�- �.&|���N?w�&��.�iP.�>�Vs89��[��$��gpД�o�`5��JM-�o��%�3_�d����"D�c~�	�-|�����w<kdh�~�e���d:��Q~�H���Pk��	�>a�wD'	�j���2z޴���r�*I��c�/�l��B�$�I�.f�����g���Eׁ�u��䈓s6>*Յ��+���(��-�_�q�E�z�Z��a��u3CL��4�$$HJ_�ջН0���۝�B����S��qY�F^�)3}Tl?F�U���㰝�����:���d�.'�� QX�#O���w�=lH��6��>�Ԙ��~h�zߚ���e��ٯ�
�Q��%�a��<}؇�K��&��4�Ν���%�w-I�L�>��������/s��t`�׬xw'5ع�]!�-Y%���V����[:���-Y���w����F���-+�W�s��:E__��w
�[��k�OQSR�����~N^�4#L˄��
�ܿ���m�����a�ˡ�Q�\i�~�LC!fd5��Z�^�;�A�L.��TUAo�f��a�t��_���Y?���t���ds)a	 �,(��Qv ~k2t%L���I���P�o|�1s[���.'��S_:�1 B���t�&ob�jM��о�Xc��2�P�Ү�����iZ��#EY�妧���z�C~�5����aW-�l����S�&�8@͂W�R��9��\-�������'2��&�%��l�����`Uok��
��O���$Զ�5�O��k,�O#��O=�]�>�*>&��"BFg/ɵE��hз��J'��}�!s�r�v�Lz����%v���[���y�X�y�MS�����p��ں#���v $UY%���=t��� ����v�J�J/�ry�&X_j��M�;c5�߾P�/�����׃��"�������1	 ��p�x���Gr�%�9���)B��@���y�2�oo��RMNO����ʵ�GȖ�w��Inp�t}!c����@w��eF�ù�l<�rT���,Mk����+vŌ ���GE�M9�޹:Z�,3���û;�c�_����Q�1�k�O�!��&�x��Pˌ6r�h	o�rul��s�c���b������ �U$?���hxJx8�C�:�q+>�Jd,3jet�Iǝ�!�k`�cj�f{)(�Nijͼ�����".��`���o0��I�Fx?����V��P�^	N�g7W���Oߋ� ����⎬e d"��.����t@T04pcL5F	�.0�tψ���r�����u/wN����1���Җ��2�l�Ԏ� ��:^1F�;�&g���l[���1�)\����1y�RcE�ԇn� %��Q��-��`֦6/��"�j-D�V��Q(�Y�&��FU�w_:�X�
��BH(9��"���C[�t!\K��p���n'�s;�~�q?ӟ|@�b�z�i@K�ֳP�2�A�}�8�/ZL�P��ꢊ԰��)��H�(��C��3�M�K*]��j('�i^QĘ��(/�)��e7��r�6(��	Q'C�/���`�g��IAٻ~"���8J9�~-��y��Ҽ��f�έ���O�%Oق�9�t�a�����o��tN���5k��s*����ᵡ7R�%�!}S~1�u�	1�bJ~�A��%�1�E�4�T�v�ٻA�!�"���tqPi���7�lH���q������î��4c6D�X efd�WS���m�I�t%��¶+c��b��g�?Nh�;λy�0����.T���&�� & ��� \dQrO�-�5��f=ם8*H��c���+��/�����윯��BS2-��%�H�H�/�-U_kG�����/��饨NI*�"�����ib!�y�K��^��aB�����)	�t�"�6�d�ȱ��x,r4��p�"=	^����®�(��*�P)�I�9��#{�)��\d������9�Obr޼��9'�)�b�M�SE�ٝ^�o�z���*|��s�R
p�j�Y��.� N#깍_W�.Y����U .����(�Cm_���%�\���i�T��U��ٙ��fZ���aZB ��������y1���~�z8}nU0b�+����=��ʧ��m�ۃ!3�'"-��ua(<�E�A�/G�j�!i��<h��4	 �TiF1/�>�[S��?��M���0N&��4�d���p�V��fѽ`�/}���ꕙ������ބ����R���a�Y�1}�D� ?2����ܥ�x�+5���j��
�PW3����ua��gM� &���z�b�:{P�W����M	�Xm���벏%dv]Q�0�m��jϖ~�" RC!y����S�_��#h�.��nIݙۺX�gQ߀~�O����"��?	�ﯫ���7���?oxT5t�t�г�u�k�5���{(F�N�|;�Ŗ�[���R�Ѓ��V��#>����i|-�u�E���#K��\�cTӺ=��dT��ܧ��>�ꆷt���N��7��羠11��6D�������+�w�d�K���Qs�RY����Y�-u=J����b����A�'v��|�m%�S�����w�sph���MQ�W�ۭ�����o���#2�G&�L�2%4�K�iD:��^,�i���Y �(xS H�:��k�-[�+�K85i�= �/&X�	�>�F�r9�>[p��A0���Ҡ�8���yϊ\��{[�wT�,J� �XZl�8w�����|�����4-�	F�1��̤O����>�+�A�M?�M ?֣�c��B���Aֿt�=�N������Z��F�L���F�Go!k�
c"�V���"G�g��#�X�Y������3h�8�R�S7IP<��l�7��#(���:M@���N_����3_]$��^����oVE��;n�U�m�SF�R���>�>����ݿ���gQi;�ʄ=�'?�/4B�$
��Gh�l������s����2j��ےmZ|]a%����)֕/tL�d�r�J��Gߢ�s8UGs��4�����/��6	�uM���y����5sYP�}�4��B�+0`�КZ|��H �JO!��%R�M&���ٝ"�
c6�ebP�f�d�6�&K���	 �|Ί���`H�����"�'�"o��K/������MB����0� *L�h�<`�zp�i�a�e���4�P{a����`�������3�[BP'$�j�	~{�c�@� ,"���
�^���c�!����b���i[{/j�m��r�PavA�Č�0��`� ��56W�� ]�*+�k�s�B�6�g
&�!K_#����C:T��j�yN�H���8�ў=��P��A-��wR��Ri��V�w{=ĩ�w��W@���
��R�v,]<k0���=��%�E�Py�>�	��3��? o�f�6�C.�xopu�	�l�08VɆp.()z���Էh�獭'�8N�!.��|��ۄ����� (�k�_�)��9,��� ��T,��)���F��0ܼ�8�w��S�U��w�i�Qz����R<���	w�"�)`�4���,l	Q�d�,r�;(d��Y�	vg��~�0����&�D�ƙ��o�HA���������L%X!�#����@wZ �N��I�����(&�����*SD^�e��"'e�8 ڍU ���~=L�x��D[N2z�R�&߶7�W�)�k[OdMs[�Ӱ�l5AgY�M�p�0;���t-[6���5.�3���Y3ޮ6�d�îslsI�w"�ԭ������g�~%N�♶ɭn*
+i�iY��FZ�o�~tI�wB�kX3�o��D+V��*밇��7����N��D'z��e$쌓R���n:��=�3�Y2���˙݊��x�b)��hPD�
!'�c\�~5s�#i��;�cNH�zɫڰ��;�S*�V͹yf��������
-�Z�����w-+���ӻ���|8�:a����m����>	�R�
�z�czze��N�8u%^g��s���
�M�:#�&�	Y��M�[ŔHB�Q�tK	P�������>��ݐtR���"�O�	�����a����0ew�"���4}D�ߜ����Y�M�����\��#R�TE��K�ʑ�Ȁ�z�"�{.�i �j��'�¯B4c�a�k�4�1�y�t<�GBϖSZ���u���(�|!��r��bk���=�e'�P�<�a�9I�ȁ��'at����0-}3���P���.�7�����{=Rn��8��!�Z��yg5���i�!�K9D�M�s8]c�>d�������ۍ��|���T��	/�20�L�J���C��A������E�����v�\e��1�a�ӿ��ܒ���Ǫ�V�ۂ e�E�#�Y�pxuń-��9�}����e�G�]]���-�Gx�T�<�f"��k�!��{�↻�����.�s�<���++�Ka��-�Z.���r���ɴ:I�A}	 �g5��
�Ҷ�VfE1�Ut��Ɩ~�,w��YY�Fk�PM�km�WAn�^R^T��������=tI:�c��d]ie��]*��!lK:�ݵ��mWqY�	T�z�S%(E� �m5�+��x2O˃_��g�i;��y��d���s9��-:=���
�o���d9&*^Z�.QBU^��:�:d�<���9�e=1��w�f.�����Ġ}a���L�g֝ �S����P�E\A�Rݩ=(�P��a���BPUpPj|�E����ښ���J��nn87#O�OF�n�F�jvo���
���9�A�((���Q�G�Z����õ�Iܽ�:'V�*a�c��}����o�[�D^��7WX�/�F�xv#GM��<�.������I�VS@Ӕ#5��'���/��q�mޥ?���b�*�-��B��fXZ����)��A��<��w%�ź��rC5Zގ#�@?���Sw�r�0��/��u呞!4X6�
#t����B� I�x��ֵ���a�w���56�m$��w��R<[Y�u�� x*6�7�3�4�_�A�=l�P��(Ԙ45&ζ�	������u|(6��'��zU��3���3bVO"��g�Vb$��ꮭ�m�2I��#��w_�5�"-{XS�t�Sj$�B�/[��P��=L�l1��#�~�|���t��I�?Ѿ�RmE��A��:fI�m�&�X�CL��S �A������G��\"�n���H����G�'��ŰP�j�y��1c��z�?ms����]��ug�X5���b��m#��86��)�l���I���d�P���YGr�Zv��).�+�
{@��RZb�Ĉ�(]�$��rd
�1U�;̿�'Wl�}�9/�ķ����6r�j��+��#��ؑ�N`�/��p��@x�پ�B3mxCw��4���9��m�j�cT��,�U���[f3�UǏ|�h����sAVu��dfJt钲0HUVu����3�8i<�,ޝ6_l����ᑋ��J�C~L�sM�=n�M��p9���鲢�O��z�v�JЀbM]�� cm<5�'寺� �Ц}�&[�޴�7��Uҍ���m�PT�y����gy�;,��3X�(9���en)�p��(��l0��^)�e��u��p����㹨LpDr�4�%�XcD����E�@��Hr�1V_�,ݺ��L����0�PEr�z�4���\��IE!�7%/�M��E�5w\Ơƨ!А�b�p�q�Gƍ����M����E$��>���Ҋ�ƕH�;�&���%w�ŧ�[�#T��GNr)j!�����܈I���R�.z1��Ñ��ϼudb8�0�d��T�K3.�@j'�}�����!�r��s�E~���i-�9�����L���.$h=�����b�j�ܬ��"������8���m@�a���(�FNá'���(*ҍ]�=� �j_��h���ޟ��@�g|��!Y���9R�ƒ�+�]ʜ.�Vs��}�6$uz�z�����*wHl�Э4�|7�=�T��>�6��o�$*g�"HE#
������_f<�Q�:7��'z��Kmlt}�h�\�.��94��h���c`6�.Wsm@A�n��4����w�����؉�!��9�Q|5������u�/���\��6{�\��N]x�MqFP�W� �>�ӷ�:H8[?��<����&=ʓ���La_	���H��'�+kzT�R���T�mh�V�s*�%�Q�@�
��BP}�u���8÷5���/��6�$��+$eӮK��6@Qa�� }�b�$�Dj�lQ��S�`U�x�&s���]���]����jng�U!^��'YF��\}���AS��Z�z�����=�Y�^{����%(�f��9|��->�k����Y�-�hJ����%�?��M��[w������H�:)����eii^�_8�=��qIR��v�0s^	P�a�w��S�H2#i}�˔B��Vr���!H�Ll@���{oY��z �'jKy�DdئqX������M��@��a+]+$���2F~�n&@��ڵ�y [4��<Q�DG�}6���{?���o\Se�#��:8���|���+eK&���g���m�Ĕ|6�f��y�g��(8G�5�G�J�:��r�"6��P͊�|�mQ�C��65��$�Yv�k�N<<�)C]���R�!8�&�;Nʸf#Z���流�v4���=ϭ�� 	������P-�|�A?���:,��m��3�1
����g�&��K��#��B �+�7���O��V��9H?o�Z��EqU9l�a�� ��i��/��C|�����=�=ó�v[?�6$���;/S��%O���_��#��<fr�� �>ANo,6߸��/÷�T�/�9N#�gݸZhѦ�
TxxزDU����5������SZ1F��h1��A�,��(����Na������1 ���au)@�MH�1%�/IE���o���r9�l64���D���4���2{T�z�)��hN�`�w{A)�BJ�4�,!z�D����;;�����n�
�O(���e���h��'��E��:"~c,:B��D����б�2�ZF^9�v�RYGNWDv2��n���S��+޽�����ܺ�����p�o�r�j��鮫|�S%t�b�Fv"����,ML��Zm�i@w�꒕��gr�b�����Sx�|%
����ۛ��q:��03��~/���U�����(o�`_�bN��n���s�޾�Z���"�C( �p곧ޚ���*ȁ�(�M@4�:O'3�@`�B�Kl�i7�GK���m�c-������πISn�t�)q~��{�{��Nc�d�K�N�ܕ�fУS~���9����:S\���Zu-��zL��`6&>�W����=�/L�$�.t�}�,��odF�x8L��n�R������cz� 5��!?G:��h*0ɦ��1y�|��c�[i�d��)�q=M��*���}��4X�JW��\Q���m]����q/ �}?�GF�k
nK+��g�Fs,�Fp�<L	�JO�Ҡe�G�Ġ��.7ϵq�Y@&�z<�L���toF�*p 2�m���m�|�(a�v��B�Q��8n[0�a|\v�+NGy>Ĥ�J�#784pQ����TM9	�AMa���k��v�v����(�'��D�i�{�+nj��Pqz�s5��x.S�"L�'��m�V�5 s��ɕ��G�F�I��%������^Y�S��j��G�+}*kG�֛�|�mC��./����4
��Fk|�0�88��������݇/����k��}��x�4)��ι{�y������q����d�T��1�0}@�n>Ѭ_�j�KDz��./Lp`(ĸ���6>��J7�TI�����|g�StF�ˎAٛ:���{�w�eW8�$�h� L8Pa���q޴0Pc����5}���G��w�}�\U��=�I�?Nh�x[�:����$5ݍĪ
LF����
q3~^��,��)z.caߝ�4�Z�&b�I��a�b���	��L���S>����짮י�_cw�ěC�{���T�L�[���m�LT�~����1��f���hK���p��
�3��]!fՋ�� ѯ��3�wݴ����&�_�U�n)3�m�߈A8i�D�vT=j0�J��Z|J��C5gYfA?T���"e_��T�"0��Ձ�ut2����aV�v��Q�h�6��*�f.�Sh�����Z�W���[!��*���]B�y�5A��?��o��{��4U'�hy�MJ'h?�=4N�"���wF�1�z2��3�w������dSܛ�+	!�rL�zG(�d�@�{o�M;�Z��0<�,���Lq�� %�sY7���=ݞ!Z�F׉H� ���7J̱�3�U�W�[?�Eӥ�1b��6ϟ�M��E+�# �`�̀�|��JzA6�jH�ӕ`��C~�v�(����0g���,�넌�a��ο ;��Q�X�#I�q����(Ӵ6J	�3�S���P%�>����d��I\t�)#�J��:-����?Z�f�ﹼ��Wu�5�N2�_g�*�t,~�U���I�2��Q�\��5��.:xTP��Z��v=ො4�Xw�p;��u`
��׶�j�ʤZm+�q����c�V��"n
�
n��O�|�gNk�{1���֍� o�$g�pO(���i�a��W���)cu*����n���;On_|Y��:���d���#�C�1������u������N1�Z�S�|�v��e�}崌DAi����������<�&�U	�3I�	,��&X�-8��ڀ��M�Y5u��6W��6}MzJ+��P8�r��z��ېep9������"��n9�gNꙁmjs�/�
�����!�9B�p�*"�;����N1�[�9�4�kŋЩ����%!8����';ߑ����-_۷��˼��7_��g�oA�G��|,Jvc�o��T�����R����e5�т��m��d�?��nۄ�r�� ��V0]Դ!�[xZpd���0��C�P��f���Lf��>��sgdtX�����p�!kI�����$r�рF�=�j��V�z�<_�&�f�[B͞\���W�!��  0��<n.+Ƹ���V�!}3W�w4gϰ�z�F�V.)w.�*N<�����n�C�ߓ��,"�Al�c�G>��H�N���	\�G�!%�9d��Φ��3r�ʖ�d���H�2u�KaM�.��if��Ji�}x:K>�.��<��6m�(Qy�D8������-������Z��(�\��h�����ۉl�_�gh_g������	�ؿPW�[tw�Km�j�����\hm����$�R��*�ÓSl6Ŏ�/m���y�wԪ�@Mi���Iûd��H2�!	����i-Z6��H|l��j�E��o�tX��q��B�_x���hܮ;G
Rx���f�q��C,ol]],���\�|'v,�Y�W��Z������LgKW+Vް���A���%Y����ɲ?K�(�A[��)���,�����j���e��T]��S���MB�Z�*����I>�>�)���R+d�te1W����Ds�DY(_y+.WB�V��?���h� �<��� O�.�@��A���%@�ú+���yiq�،^j^��hYҦb6����D������,l+>A�[rE(p^�w�:��e䯺6��ޓ�S/�ZH�D��{I��j�B��s�S]k}�~���>�}�FŹ!��hS�E��'�Zj�kfG��;�K�j���8�N�R������AB���Љ�|�~.�^~�X��%PD�����|"�������j٣�V�u}&�HW�Y�O��p5���v�ZN~��G��w��>n3@Ff�&]��c�خ����$�3(xz5��y�󆅱��7�s��*R�����b�SG�O�jJ�!\b��>��l)�	7Q�H�V�݂�%��X��.���?,��EAՔ�l:v��1W��S:}	�{F5M9G�#(G�J��u���W�vJ�kVG�l�T�� v�8~_���:�R ��3^'�%S!���ǅG��0Ć�^u���.�����MC,��ݯ�k~L*_K�=*Bq��$Ep���rTda.�o��m�j�����3��<��݋4Ry�z����*ޅvF~V����*(�������3K�T��T2o�+�Zd��L|��b�2��j�߳�7OVź������R�g���Op|vx�fM�V��l|!:�x0/��۠�.�6�.D�Ԏs�&�	�UwZ��Jd2��ow�۬Z�<#�?L�L|_7If�K�ON\|��eH6�Z�	d����(U;�-T�v�I�"0TC��,��^�ܐԒ�3?�"jٰ�
���X�akBE��x㟱SDa�����p}���9�Yy���#k�F:��Uu	NU3�FltԈ[�6w�iC?��k�j��h��<��CK�u�8T.�î
�f�����g�AkP���Ɩ	���q�n'�jO O~K D��^�F���YP�+����yd_Z�������x��ݢy������@O��E��xM��������#�2�{;?y<c�?q�Xo�{f:�����〱E�%/Ͻ�e����J�����=?��c�E=���`O����%tװ�p� ������2M���i6޷c<����/U����)�q�m��������^߃hu�d����m�[��r���k�#�Q�[�%�6J����K6�}�dz�N���u'{DE��gx�{�N�m�n%L$��#��t\��Od �(]�o�pB��@�0��Od*0ȗU���̋Ʌ3th:�p��"��ÝPf���.?	�&GD�)+Wʿ=� Je�~9���z~bS;�L����d�\C& {:���}h_xh�wHPʟ]�'%Ʌ����SΌ�R�X�n.���lXQU��C7�Y�S�|���1f����T��mT�����a���8>R�@����"��X4��Eؤ���m��\�$~Z��yn$<��M�F݊�W a��(m.���X?d�7�E����Tg Zϛ���9F����P�Z���M�L���H�J%��(��٭��2�G��|�{"qO�~�g����C�3 ���0�>e�����6'�2���^w�@rSk��C4C�2�p�/`X���g-Ntl�	t����^9��m����9:��5n��MzvE3��E�P�����:0�O�AB!�j���d^3��N�m	���X�u!�7"S`k�N8��EnJ�\꫶�.�9�?w�1A\�fL�e�+�xo�s�Vī�[R��5�M�Ϭm,<~��i���H"��L}�JT��ao柢�[��A��=d��s�y+?�6���9�
m��������LDoxw�ɢ7�uB<=u\��L
=S��)�^p�P��wZ>���u�����q*n7�V[Ge��+(>�V�0G�*��d���H��T�3
�{<s����W�&����]�v}7qހ!��%�I��$!��5��0�G�d��������ֆKbz�Ci�ͳa��lÆ/�ߨ��*v}r��X^Xč�>��Y�p�=_�:���-��$�)NT9�d���/�%�{�ץ��5߁������77/L��uD�9��)��Q_���W�I��$�R0ܫ�lp����S��1��������~R��ʼ��%�s \NC�!�ȷ�|�C ��'wM���O�r��?u�h�T�?�|ǈ��&��+[rq�E���w�M�NӖ4i���2xE���g���L#ґ�^d�l?g�������)�@ci��aKy��!p�3�p�C�U�Ė� ����C�5�S<��N���j^�����5�;m�V!Ѳ1#X0�v�|�i�/i/$�'c�g��?�/@`2�Wp@^��W��
��%��cH���)H���z+�����]4�gw�a�*Q��[�����]�Fw� nR�rY�
��vP���;�B"^'��`+�4cz�I�i�N��"�%�1
�y���,ů��^�69������rޏ\�e![������uȭć`~�Ƈx���yJO�C,�{o�L�}�X�N�;���J��؈�~6YIsCj�`2�ČIyr+W`z�Y%�($�W�9K ��γC,���U�84tC?U�ڭ����ߺ�\�U�U������#%�D�:�ј7�#�Qj<�D��ೱ xO��`Zd0�K��wt	+Du��2j. 롡~g�����/�ʹ�>�_���(��G)���1/��؁N�uTeG��)k*`�~FS�Vp�H�d�>�R�?������]����jGS���~�����:�|�!�Om��������CT��k���ǡ�&z�#��%ۖP#�a��kF:tn��@ �^�����������f�|}$9;I1U(t5jO���-L�!c�*����(>������� �I�&m�h��D/wƎ�=����n�9i$4���Ib�/��oo��8奩I�F좼#1�<i ]s�~]��關Ϫ4�p��<���npo>���[�HF6ɔb��gO�Pœ��s�Jng�ۋ���t3���*+C��B�<Δ3�r4���M"�\�lx��7�ʥ�m��q'�O�-M,F�&GNT:�Vg$�.7c�*
:��o}\�Z@Uh�k�gH�M��T(ຣ���å2 ���1*E�;	̡~<��	 ��V ~�T/U���_�(�y�B!B���x�j�b��'���d@��X-��A����.G� +v#k^V�v��?�	��S>���}��L�!��;m��Q�vZ���r�d)[�,`5}�Gn��	H�=4@�kc�o����A�M�(�=0��m1��Sq�C�� Zؠ�����nq�j2sGDl_��a�V��3D�)��,�K^ϯ�=�?o�����;!�6=G����M ��8�L§1����Ӊ��e���6�b�R1
�ߕ�3�N��L�<|jz��n�"*Ց�g(> �y�'77~Tդ��]�X��S\FuY�����uY��.��в��s��0a�3AV7���
��J�f� ���(K�i�3ی�Q���6i^U���m�+� ����`���2l��d�G��'�&�D}��.�H��������bҮ7l�M�*��F�������=�e�Ж��36&�i�����܏G��a�|�|h�1�e��3�{��<@�6����p0#��������j��f�3.l�ӡ��j�oH����4%t�5?�̿ߠ��Ӭ=9N@5��qw�&���?W�c�kmwv�*��RL�F¯�
����7AX����������*��8��s+n�Jd;G٪h�P�뱡����Q�W�7^l�	�>�ON��'�lZ���-L8��=�0bq<͜�VjQM��2��wuD^96C���rv���`.'WƄ�CV7oI�!�d��㢁_�'��k�W<�ޣ}��ES�؇}C�����$7PT���Y`"�]p�;��$M@�8>���]S���6h��
�6�t�	�$`{'�Q��4�be�K�� q��Ed��z�ۚ�(do��󣸁
�(�W���?{�䒙:��T�w^�)6��!��|�H��"�6�]�l��p��3%�s��[J�f��
�,��-��D
Ǯ����#��0f��0����q� B=4 4�j�:?g�SwO��i���%*��w�
���4��QJ`�>�_.��
��U��3���Y?������3�]�7^��ׅ�y�)�b%��N9�J��+$I���g��f�[�/b@rr0�3C��Z�ކ����ݑ�)KU�l}�@+V*M������=�,�/!��K�SoMdZ�����!�ߍva6-�J��=�,���;��M���U��Ǭ:���%�(�?������\a�%�ؗB��ڀ�4����Õ��U:4��/���H鸵Z�ӕ?��T�Y8Ӫ�=�D���9����n�T+�Bg������/l'K)>�<�)� _�,� e"SX�Y���zQ���Q;�q���!��bjS�qر����S%HR^J�ϕ�~�����k�0����q#7Dm��A��G���%3d��I�3�q��\����T��d���}� �N��G�pS�b-6��mHc�W��*Ґ��|�N�	Fk�βj�!]�tQX�>�{����l˛��E�����$�/������������� �Ht�|!��fC�V��}@vү�I�g�ap{�N7l�g��!*(����>Y��Q'.KС6K��A�RW���ߠN��?��H���$1\}bN=������;��[��n�$�`�q`A.1������_�L�D0 �(��5�j��cj�|♲ooEڲ[HM�=7�2�jE4uwV��K�C�	�(�n�nݚN��y��h������ek�ƕAyu^aB�DTc?�swǞ���uYrkІ�}/��ˡ�/UU9������L�D�d�5���� )��Rs�{�FR�6�IBPyeG��&U�4!���F!��<�7���l�]��j$1����j�b;�RvY~d��٪��4 �\ӭ�Y�8�8�P��x��r� ��qB�n�|�c_<,Tv�y�q�20��	sJ�����,�ߤ��F�݆�$�
\c��1=R,[��¼1eB �F&������]<>#��;��S9�%l�!�8�ڜa���V��e�ɯ����o��T�L�'�}����/�J"��F�RB'��~^ù��嫾PO=�i�����q�s�*ژ�_ӊ�)$�5m��Ҧ�����Ldֱ{N_P���^�g�ɝJ���D�
͊�,tY��\>hΘ,e{���hƩ�V�rv���Sg=#�b�r�,����<�?C�^�Եs���p�X�T�^~B�yQ꟎�(�~��kހ�!zl�:���p�d��ok����<�F�a_ߤ.{�Z���%����4}�*�x� ���O�T͏����<+yc�*�h~�Q�R ��HH֥.� /���H$Y^g����h8��0_Ư ����=�{��w�S�f�	�y$���O�`�|x-��b�*�a���~I_�Ō�YY3a��!�G�R�'\���֓E������K��M���f�g��z;�+lI�Pc�1ݸ����9��ʧ����_Ƿ�������`�p<.��Ayt��G�!*8d�����*����Ug�}^^|^��P�$Y>���j�	�=I,���O��O����f:���� I��Il�G{$���//k�BX�+�����W��i��fNT��n䝻C
(�1��疅�7�w_"�U�_�W=�ƍ�k�˨��\
X���oM��!�w9��
Zp�Q��iI2�ÁG��݊�PP4�ʞQ��)%^9�c�i��k�t�#()���.�w�Q:�n�����{�=��JS�A%?E*Y�g�?�x��$k2����dac?�
d�����B����R���4�Pͱ�qz![�%�1攓:&0�4�a61�c��C��d58#S�UC�9kx�#g��ԁx-�a�GƠK���K�����TH�rT����X��	�ʯ�����x���l��E%$�O �ƽպ�S�.bT����5̬D ����P58��(��G��֦�b#���/�$+��M�m��r��.��R�68t,�oTT����\�U�ےǎ�_�1�!�iqh+z	DE;�� ���#���eC4�Z-m�O�٩��.�Gő�6:=$���9c�ɻ�D�YO�Ҳ�SN%��Y��{5^6Y¸d����C��KR�-c�@�3���;�DL�	x�Z{��S�(q]���qt[����mVY�:2y��Րv���A�t�r����DP�;<k�|p�7�^ęn��Ӆ@?Ѣv!9�����FF"��#*oĬ�h*a@#Ma4I�Ӈ���|�y9Uu}U_����g��ׇ]��cバ�cn�+�n@4Ivt_w`���cm���[`6��L���O�lWŊ�øMA~�;<i�t��hLy�7�����{'�E��>)���b�h���tǘ�u֚�����׌i_���Y|��*��wI
��t���U�è[N�Ȩu����9�PN0��� �1Eч#F>�S4�D���c�U%��x�[��;�%��}����������=p�m�$���2c���X��"��g����e��c���C�J��9%b���Ż��>���[���CF&@H2�O��Δ�Oq�x�̟ƀ0������
�č�g)��ZBΥ�$���(�'%z�jXe��t?e�����F�W1< �0'�maL&�}[O->��m�]�5���9�Gݳ����&	w�AT��.��r(�wEZ��)h����s$���靫�k���Y�f.L��6�����2���؂��������x1�D��AiQ, IG�i<]�k��(eT�� ��OC=;�(da� l"�h���[���(�V�ZNb����f��&j`�6��M�3QL��:9<2.�ut�˻X�n�(��H���Nngҁ1�"I�:� ���eoV�5mߏkV����"7'�3E�3������E%{�}�V�M���#��3j� 4k�.��l�[�����Vx,�n��6f��m�tS�w0,T�b�a��&������g���{M�L�L����X)0e��4�a��i�PiZ:�0�Jt��um�W�f��>����5�<��}49Ю�JiG���,l%�32�X,�i��4sQذ�x#F���JS��HHg.��K�C=p19��d���Ob<s���M�2�ɥ�O J�%olYD��ڇ���W�����"���p���Lo罶1�3�+�F�Q+���T�������b������S�V�c:�[�z�m��̾�k1�k��g��Ӟ×��՝�Mւ�k<���1�\iO���-�$Z���'v�5�<��)Uh�4�� �B�EȚO*F��v$f�$�5�	�?D�N�/�_��_g��<����:XPa"<�J�^�o*�2�Ձ�	"�+��4�ISVu9�{B���_�/Xۖ{خAv/���^9c$������/'�5�=Vɋ��1�
%�,`�|�D��`��|��$��ۘ�������)� &�s��*3�ZR(���:�Q�W7s�~=O�I,`\��{#��G�V�#�I�����
��.Qt��ڸ?N�U�T(4+$y���jnU-�S&�u���֐Y0�m�@%�)��u7�� I�x�����RL`�Oo6�'a3���J��ߙs�a�3(V\bdq[���s��i��JZ����6A��b��lP𻪝y��	���G�6���u��K��0���j�Xu���)b�w�3By��Twaʒ���>q��!�-Πh۽�
��p��V��t���Qh����։g�c�@G��2�N��FW��!Q|��t��E��ڣA�����^R���e��_YG���W��������l�O!��5���V�������@Z,��I'�������&�ͽ��s��uTdZ3��+���"����Ù,�d���\�q"X�xr4P�6���Ct*�.���5�dI�=@_ وF��g�����$�ܢldUrd�~�k��L�E�킘�q���D�0<3>��BYd����� J8X>硥s��ʂGY>��@�,�]��r8�N:�l�h��0���j�P0`��5�c�k��c5>s�(z��NWa�����n> ����K���������&�N�$:V��Z9��m�C�C.�d�s�E	pESO�rk�g�
�p�"[���1�P}��q�pt��dS|�cm��'� �.0�y%��e�8�rr�&Bw>��z6�]��7�6����_� =�^+���3h���vh@���"��G�|L�9���3!F".�2��5���`�v��쪸�Ds����Q��2�q��c���3 ����r;��ϻ d&��j}�{`���'V/T� �����_S�\1��SA� Q�a�4�tX��V�@f�?`ȇz�>�v��"+�m�ڒ�E2�!��l���%+tޚ�]�D^�S8� �r!Hfu;mc�x{G�Cw
����^s�=�����΅�҄�2OH���!����X�͉i%6�WM�S,Ħ��h�\�t�Wh'�H,���T�u�G�1�=�Î~\�BE咄���\�r����5�_{��+m'�s�kqwjI�"�:4�/K�e�esg^�G�I�[�;��-�u[�����?:,a�Z��s��W�zv_F��L�`����z�
��Ԕ\�Z���h�9�8����8i�S�yO� ؃-ԂZ��s�]!N)eR�G��	i�/�1��#0ˈX�Vz��fĿ?�K��(�Հ�0(����rk]�.���e��	<Nc���؞�����FN�N��:�$q�|�[�j�.**�ܷH�w�b�oJC�i�a~�M6kg�SA�x��w�����d���'���	 jŘ-�"l�����'7M}?�f`�!�GnP�fddImI�"�7J�z����D"�@���k�=�P(�U(C׫'?���ϩڠ�F\�? ����_�����+�ʺ�r4o=.pC��{��Fln;�/�k
���N��a�c/�$P�D�e\��#Sq�}�e��q9�iW-RIC��쵒���T�b �S������(`��(=�%K�Ͽ�j�萺�~;��!mD�6��W�z��p��A��z���[҄�]e͖�V��v��4'nh@�K4Fj��תe�}����7�6BP���,������-A��� �?F3Od��'I��	��R tq?���](�K���靠��c�h8����A��=*�Ⱦ�.\�����ح�\(KKZ�}F�������)���ǰ�,�?kO��e#
��`��M+tx���6�|H��xj���WJn�J8g��gj`CGʄ�jۙ�=ތ��Y�E�g�b��pV�>���7��/�������E,Β��Q�<��(�눡�P��H�a�[f���g���d�*��^L�D�
(F~'�J|L��b�Fo1PS�ؐA�U?aj*�ax˳�����G�2a������3}�}���im���m�9q�����A�IEꈽ�{û��� z�{O)*�^duhz��v!$��^�<�&�kG��]���Jv�e:ү�ؿJ>��xn&�m�Co���~�jÏ��^�rM�£�]�⟆ʀﻬRvyj�ۑ��J��B���A 1=ӱ���e��2U��;�Q��c�3/)z�����c��Q��/M������AUײ*`q��E�L	�Y&�ZX�o�� �#'Eȝ,S$&�F��:�kR9y
�+��@ۤ��~Y������=�#�#��F1�8�gSu��i��v��R����cT�q+h�(P)��k�ղ�
�ny���oMB�[���T�g����	
�J�}̶��Ps�L�;z�dX��`���=�����`�
�9¶8�B�N����`կpL��zZH���e�Yx����6�q���d�aJ������˽�j��V*�m� ��ee���X�mzO����6>�p~+"Ց}f���#ڕMv5p߱�\�� c�4��_�^�|�:W)���ρKӃ�p1NQ;�`�x�����Ƙ�ͨ6�|��?نA����hh[��Y�bOl:�>j�]�1aXF�M��H�#+��2s�=�+U�`g�v����8f�sʕ��d�=r��Ն��������;����Z��EEl�����6w6��� ��f��C
�Xp�E�ό�ʁa.%�Yqu!,?�D$l S��1Q��=�\�G��>qn����^E�Pf���⑴6�'Խ �@5��t�=������^�_�Z5ߒ$���iobV�~ }��$�O*;�����=����_#�SE`.JSd`B<+��|�9G@+鐈	�;�P�zs�i�"FowM0�V��GDY匔���2��6���&.��w*�8��3�."ڴ�X���,�<����|#���0m�i)�� ;}�KA�C�7��#�ZX��7R����<�j���yxR�o��rԠi�o�%B�7�3�΅�C�z�F{��	ȯ���0-s�0$��ȏ��{x���a������n�됔��Gd��mmء�Oz�6"mf�Mނr�n�,�R��7qn�q�&Lи�j��}���d�˞v�m�m�.��J.J�ih7m��1m��1M~4�D�=��»�p���Ƀ�]=!΋@���[��	���W��C���(Ȕ1��x�pQ �qL�)_s�#X�f% �oe���5���XU�s ~���u� ��j�y��� �j��B%��u����$0���9��o�IA<������P]_P�ԋ|©���r$�B ���!o�6�Vt�p�#h��vm�ѷ�6��kp���,�K�;�����iqy��'��w�����*��#�94�R@|Ӫ���Y3}x���Ƴ��V�Y�����2ۚˬ�c�%\Z�����Gv�kk�1lV'������6G4�{B ��?�*�B=0��WB������m��".MeFY�I���L�&���3�6>���S�u�a�S�z���������d�k{~�U�ՆLb�G�����9ļ�N�NK���8o���.\�P1_t�sP�q[e��BU$���Zh&��UMM����J�ZnO� Y��o3��f�m��]�΢����ON�{ۉH�,Ge�#ӏ����G $��4�'�W"���%`�Z���\<�㎸��rDg�E&�j�]pc:��ח��TN�l��������:3D��g1�m��%8,�+C�Z�j�3��L�I�~Jő�>�Vzno�k�½�~ �ȇE�<p�;j�ݩ�71r�#�{��x�7�g���A�������N>��k34bg�	�K��N�З�!�$��ҡ3��x���&>���ᇆ!'�8�M�����g��m�ʜ�*i�aS�#���+� Sy�6��Zδ�g��D���)���Z�7ᳱ2r���.yI4�S ��+�t�Na���V:��r�xGPCl8�C��r��k� �A{��S�����z����x�M��z8��`7��q�P�KZ/�R?�>�w��_��q�\Y��H�:������gJ4�VT��@_��|����	P
��V�{�\P��<^�K�����C~:0m7j�s$���b���<ة�Z~:���n��^�0pć�N[�ff
�����YƮ��a�H�M]A������m�.�d�9}9��i*�Ht���h!��JΜ�%V�����%�a�Ml��6H���ረ�e!͟�9癩��e�!��&�s0u�T�E"#���)�x�z ���g^�N��`��O�FƟ
S{�mH޹�Fm|I�	�*� N]v����9ԉ0��Ħ\��.^�ތW��5��U@�OfG��r�ˋ��|#H�Y�P��@~˽>NA�G�S��/ޤB|ʥd+Y�4�I�d�<��{)|K���5Kɮ��6����*V�ӧ�sg�*�`�vI��w�@�R{~�rn��|3��9'~>�Z�Z\Aߡ��B������} �VPؾ����L� ��+A��R2O��WS�����RB��pP(��s�5U߰����p�'ōP�=�y8���	�U�+��h4l3b>��������r�R�<d���$���):���r�{����Ԓ��{_�D%�:���4�X@!����|���uB||������LA������$��R*����+��@��]�b���x�,˓x����� �������F� ����y ���{�y�d�j���ݣ�D�f�x�5QqY깴�qh�T�#��osNe�.�t����� ���$����=^��-}�h������vm�=���:��R$!�X	�j���A*}R��z8|ᨩ��xeu����)v���<��TgL>�����r_��՞%��^z��fV��h�z�M��%%�SC�-d�j	P,>U8 ��|�n�2���6s�̄��©�MI�)�e��H����b��yrg>����o��p��In����bw��1܇�r>�+'��|�y���~����G����1�?g�ּ�S������/&�szq�mw��@�����&%)	�=��[�+r�j���Tꒌ|��k��v����0	���V~�Y�&��	�?'�]��6cO˱�R�7�:�|�W�7��hFHSyxޯ���f����9Z�_L_o�#��Y���L���!�Kl�d�9a5#��p����Qj�rF�2[)"�P�Q�J��sq�`�>L��}�3:bS6����c�R!���+-�r���]���i����C���� ��DB�xfטG['F}ARŧ�}:�_�B&TKO�@��c��g�@�2�Xu�&g��H���=��&/�+J��h��O�E�8�T�*ʶ�����>Wf��ɬ�[ �"��D7ts^Tز��	�k�\{)?o��E.o"@�K���dY�Yl�죪[$%n$U�LU��Z��z����6ӡ��`�8Y�d�p9�#��E�&J�^e����3k%I3`a"������s�]>Y�`�^��gꌹ��%$���hܢ�b3��~{��4�d��_.:��Fg}�[�L���e�0A1�e�s!ie�EșTCZ�/�\a�!1;�����IM���P=V�*�	oqr3���t�"�19�p�<7���t3|�4c~�/�%K��Ήd�=��&$�$�Y��'JtH��r��X�I��|��{�Y�c�И�X��j[0�x[ I�S���%`�\��'%��C����ӠC͟�L���2�e����AE1i����)���z�(������2���"}����Ғ#�w��/Z�.�*���c�UE9�]��[����+��{:6��۫�/b0K��^�Q�q򢡏��>Z�+�!�s�����e��6���+��K&}�2$[��t����d�	�!5J�Z�s���j�e����z�Ø yIL��7k������8&D�8aO$3��[�o�C���n ��$�w*A2����O*����t'G������e��]��ڋ�57��Xl�k0�z�^��\��b�#�B����,2�CȊ�gu�?~pģD{}Nj�<��y0H�đ�E�T���ʔ�F�<u@jz�M.�\b�@4�?�_ya�6*�f^ˀl�s��'p��uނp"7/��
^�$�	mGneɇ,��V7W������2�|�7xa�h�`�n#��z�1N��G��Em���i�)�O���Ԩ��3��쀇g����Vy�e����U �E��y�7���U��?�_O�L2��-�4�]���#v��&f�oԦ������"$`����32W����Z�/�p�����H���A�0�7z��2�HDq\�<[�� *�v�z���X���M�;E��?�=�}��n}&�9>fFP�dz��6�]�|�������lN�@��A��a�~ڵ��z�瀏,��!��C1\��Nٜ�#�P���~��v��K0��У/��-9�$)c>�	��5G���Ԍ�U��&w�=�aX� Xs�ruR�0��PGxNpSp�5[K3;d�S������zt�jன�`NnY�[��r	U�p.�0"q�O��~�ؤ���N \H�2��4�,��,r�of���S6.�Р�32dfԧ��Ov/��x6 ��5x$���CGt�ZHG��c^0���R����~�)ۼ_��ب�?�9G�oA�z�Ϻ)���(�``�h |9�ӌ�~T���-_u�E���0֟bɮ7+�a<��9��+�e&�
��w�(Z{�c��I_Ϩ���&%�4k��5�"P�x��;%�9��K��-�yz#�g4����e������� Q1��'�'���K�9S&��v�,�[���d!W^<�咠!�u!���~T�WcUw\[n����g6�ҍ��k���J
L���
�2��(�[ �L��2S��$��~�0�����\�t��F��2&P�z���V_��l�y~������^�He���ݷ|C�r����Z=˂��jSb6��N6`h�+0���b`͵�I�DP�*�k�f�W1�q`y�{pE�-�/i��n�e�Y�N�O���$���3��0������a�L�ɡ�*����ܖ��卬0���r�/M��"�ub��+byɏ��`	�|����Kr�:�_^�7����B�����&#fM� <ZB�K��S�F/����4�<SG�Kw�E÷�:&8G��G�xO�-T���.��ؘi���̖C��選���sd�@	oX�ԇ�)~��l�̯lD	�q�
Z_p����&�0^�o�3�ֈ_∔mgQ���^���Dm|K���Cݼ1��d�L=���2�q-�`-�R��ҧAc�K����AM���b b� ���d�d�8� (*�W���C�H߾H�՛��c��nV��E4`�:�$�G�_~A��N�o�x�bl`��غ�� �a����;.U:�>����f�U������R�k��H�,��,��\e�&��V���{��7H�هV�6b*M��w�49��^�uߌn����9ؚ���;�����-�_�D�c���[�:�݅9�~DA�^��<���&,/�������5��Ee�9U>-��%U]��>6@ԌbB2w���_&�ۑ:E	d��q�pE��ˁq��k��gܷ`[��Wԣ���=��#�iRX��aqv(�����)�tY����h�%3�Z�3������M�M�9�e'���6a��^u���gZ��ۻ7+�)q[t0F_K"��9�҄������j=��2��aOcE�FX�����i���L�W�h��$g[;3vC+B�̯��2�SD�O��KAt$��#��'�@3����`u|^���7��!��kU������	\s6�	z� {��l�Q�iy�?����PU�ȅ�枆�Ou���3Bl���p
�vD�{{l�����:��8w/�JMcd�\�0��v0/�����á�[��C�8��f��5�ɬ�&��E�]�c�*T�ʭϿ�=���ϟ�b��tG0�|-�7��gI(¦��rOL�#f�ͽ
4d���
�⧸�����W�e�d��n�a����su� ����ۆRJ]m�y���p�f
qQ�]�Hj�t�x��ȫ(�Wo�җ@�$[�\���� �Tlj�j��^�_f�ȣ�)�?�&H}XxHMI[�Fz�d���%�5�j��ӡɏww�c��ԁ}Gq6�m���V����9k�E5���ǧ��$w��f-	j����ǯ��.ûq�E@X�ܕ�2��ȅ�h���0�����@{���Y�H�)��Ncd&�jd��j��=�KN��ڎđ���#v� G�(.�TYԆC0Z�Y�+
���n)�5xn�3����1�}���y�����"�^�+��n,���j6�+���]�+u��*�@�YYzn�� �L8�=�H�^�ۢ�<t�ǩ���/�\2�?��jA�?����{�)�m���U��w�]2��?�������p`Y���Ζ��L���H�7�5�YL���O؍v��&�xc+��� Б�G��R;뉿���뀰�@�Q�k�u�rRZ͈��o�u@<0�I��D�B �d��b�L�d����Zh�<��AD�T�ų!��+������&�P��,��g4�v��#���yP�t{����7m)Ѿ�8>$e�_ɋYQ�ъU��{iLS�%����_�GK�	 �Ð����״�!�f���,�L�	7�м1Ѳ%�/��qգ~'h(#n�E:�SV-�w�0�#?�˯�;R�ߝr�]��t��	j1��'��9=>K^���y�E��(-�:��k[��Xq"�q�zRA�ྃ�~hʂ��.�B�{�y*�|t�}��W��J�Vg��Uϟ7ŧ��Y��p�Rٰ�mO�љh^���C���޷�z�<o�{���JC̗����)�b��q;Q�����L�}�Qr3R��@}`9���TC'1�,���4��_*��S����a�5�1�LS��m�����%|�M.��C��GQz�YtB�C{K�c-&T'�m��7�������bk�����x��\�U���²�JO��#2�fy�5��~D��rp�懸�Of�I��MKA%�my�'�-�e�\X�xj�j�����j�,���(��s��m=Ae���D;�Ƹ�tI��/3���4�!�vm�|nxJ
��� �q�1gls5$f�~':&?��Ê�MX4�&Y�t���h�
B��7�l�����sf~r��Q�Z���d�d�d>�N޸D*v�!���d�_��4��Q*�t��&ĥ��Vt�@�3�&�z���>�M���?�9��7e�z����ׄ����c��+��UI�w�����Ϙ��OKƝ&�[�S��>�9.;tr�j��zΝH���X�1�� Gf�8�*���_q+)^#V�����WA�)s�n�2�����:�7�0�!5�t=�	H�4]����E��=����d�֣�h����f
�7��V�RO˅��\�������Ԇ�6D���Er|�Qvи��Oˢy�{rC�]��N+O�7�p�4�4}�K����Em��qO����x~O�j�@&��;�� ����t� u{�MbHDS�GMD\�GU�;R�D��&<v���@ �V��؄SdܶY܌�&$/��%�1#�ݪ��	��ar8�yh������D��U�@qC0�tt��ȃ��o�@�f���S�ަ�O��B�����eH�O܇*<V2��v�P�+�������͈��d)zg��������C�+��w��� u���U�'�q:�_ f�3���"	�����[�}�<O��(եCܗր�V�p��L��m�s��kr�����3:[>Ie�,'GM�4�l�F�~ZP���qd�lh�_�a��Tv;�*�q��_�n�J9V@��d�A���(,�������������q@nk�a"64�(V=@q_�g��5;��r���4�?�R���O,�@���?+��E��U]E���f�c ��o�۵ɝ�#w������%Q�-���5�q��i�� ��g��(���,���4�ŧɴ�� 	l�G�;�Y+��c�3�]`�#�v�Z�,_��[鍻RGl����L�U����8����uz;�}E�菗v:�>�[�	�*��|'�Ǚ֥#0Q�ʴu�wR-�\ŋ��ǝ��*��kb>��Dz�t�Ҵ�s�����D�0n�4;�%����� ��~Ƹ��M��P�N�HZ� ��]�*��x���1���1�a;�t
�L��}4@�q�QJw�n|9�T�M6�2�ܧL>��P�����וy���;�s^ @��H��9��9�����`W��o��$�u���B����hP�lp��e��gڑE�� tGfc�	P���R���)6?�h�������h	��<z���~���B�T	�`��#!��{�l��&�a	�	��{X�s�:!ϫ?���i�k��x?��"��J�4���/�(|:����H��k�	�A�!N!��LA�կw;�3���s��0\�q��CLmI��L��>�!�I.�첕��Z�4$�W�l�%��3�9�
n,Ӝ?P_\g�1*Lx�K�qws��e�I[�П��>��vE��VF��a tc��7���V����L�Y$�bA]p��LNӗ�i��5�9@�⻲�6���(7 ��P�q=�G�h���S�s9yK��ƶ�ڟ��-炔�K�O4��3S>��ݛ��i(]%VB-6EV���݄��Z9�{�XF�7�;эpF�����0���Y	�o[3&\�.��;���k�z�7!A����fm�J�|�=_�0�o��%]����A}�Y��ۗ����f0;��E�����I7�+B��p7~m�Յ,���7	9�50��Z6U��o��I����w�y�y�%-f��O:��`$}���� $* �M�:yI(~bp˶'�d����<K��{`W+�U5�U�A����3;�4��I�<\��r�z�G�v�����zhD���G���ѻ�\�\���]�d��5h������3a>����>8�j�7A�nߑ�/n�$���j��}�2A�<{QS6��+m�3 �ҵh��>�{Mh�Ձx!?W ��(��T��Z�Sz���ڽB��DG���m��GX%�����R	TX^�M�l�ɰ<�u}��n��t���	�[�"^蔝9�'�r=8/*��_R-�jKV8� D#H�SH�'5ؓ-|��4��5�\�K3��W�lHFE?��X�G�<���?��,�Yi�T/�i����\�����m֑L'�'(��� )J��@�;rz�����ƣ'����I2<�2��K�H<�.�qP�bDVΝ�5�44��yFY^�h�����TN�ߞ=<y���T2`�=J����~�)<p��وtb����I��r�x$�Q�hR2�ӭ%BM14VS��T
+��O�m~��o�z�q����a�R%��.6�݌�(�����㑏� '�D��#��r��چ����{i.��/���F�m�q�(L��p��s���2>��GE���F1�%�a�S��?M.|�	�ᜂ9������lVU��1����_B�g,7�0��5I�H�8ʯ�U��r9f}���4��R`�9��8Ft��S���ۖ�:��&c���������n|�����K�$�˫ W,�}y�Q�r���[��D:G�*��Jl5_�ͻ6���� ����|��t��#�Y��_@kz�#�y�I��K(����n�/;zc���t Vl~���o�.G��iUq��=��1�g�$Мy���L��E��ǎ44�q}G%);G��K��9�C�9c��[u�O6~�dkLw/���'A.�NGË黳� ��v����+��[���W�܍R ����
���~�.�X|���0r���I�k�%�{��բ`	�>���3[BeZ��O���Յ"N�_)��ƭhkZ�~W���@�������%e���S�NT���ǧ^*ݮ5"Jr&�� �]k�J���SX�� ���0����>�`�i�nQu��܏λ*�.lyNg�,�3��C}RJ�#K*r�A�bܓ|*��iY�����,�NU����h��&MI��+���3çZ�m� ^� �jq��?�\,)Q������"ǆF$T���71�\����\6��+��^�K̥��M�`�#�:v��c���QYb��䈶��EI������#�I���D�����#kJ~Y��K*#@a�<bo)��X
?4�P]wm����t���-N0	#����cW|�"5sa�YH����[Z������ޓ8�`T7���,�t�W�Ԑty38�������";z���
F-�_��$x�4^�Ɯ�]�Y��q8B(��7ຯiر���Q�{ǻ��+�L��"杈��[�n��y��U�ƺOj~������t���P���_�o���=(�Wy��,;�Բ�� ����N����L��7g-����c2�p�4�iCh��#圲����Pf���eä�B�nм�<%T��O��td�Ag.��|>�iHR��%�^-��\- �8��h&��sK��HQ��k�r�?�y;������l>���T��(P���q��ǝ?YF%]��l�����G0g-�}���<�&�Vgb�7��)P%d)2��b��D�gd5B9y�xӻy Vb����~)��xM۟9�ۀ]�����,��B..�sE����x# ���Z�z��Ԇј��� ��E'c�.|D�mq3�n���n����f��vY��.�}�RK���2���(�Ҩ+O8 :��N	d[ ��=�MW�'�.USA܌�?����Vne��ߪMe�Sf;�r7�q��߱���G���h|Oz#Q��UT='���Q�1?�A�Xx �58˲ʒ[�ze^�"�{S�jӽ��e�p���v�/ͭ6�[���}��4�����
���h���C�g$�}�O�Ғ�0K�@�Q�\T�C�]|�O����˛�)��e�AZ�:��4B�Z)C�c`��X^7����o�H��M�m@nfNC�Ri(ĺ��d�'�D䴤��\�b��SُDC�26*J+�0�(�{1;@�d`eq#/v�_X�s�����'Pa��&���M^Ug7�
�.�D��2�,[�l�H܎�ؖ`*|�> B҅jg@����9d����,�z$d����T�a�dԺ��UMF��~Ok������dY���[���4�a���2�u��}3��<+�\ bW]�1�y��/Mvץ �>���[Z]����f�W��2���u)��ȢcaR�=��dY�?t�&��{%mV��� E��o�ގx�~�8���Į���<U!�ι�z���d\Z��l���ʪ��6Zx�R���t[,՝���~ztV��A[pqV���x^�'���!�4
�Uw��VC�R݂K�`&��*
�d@6�B˷\��.�2C=�"���vZ��J U�]�:�J��F��m��2��=��5��D�ٹ��C*W�C��O�HO�p`.��c�L�}���"�T��1�2�R��ScHԮ�U��I9�u�`sܔ�_�1��`�V�=�=t��x�y,W���e"������c*&;C�/c��i]�_�2-z_�+0�E�$=�o�7�mن0�i�{��F����Y�5�8���6&H�u������6z�qUP��*�;ҦB�Dy�ؼm�)l�*���D]��o1P�|6P���aSEN&���ݫ,F�Ü��V|�|�n�p~�In0��̬d�9��
��m�V�m�H��)���!jL�}�v:�P�?�h/�H��./�ew��jV4��_4�7�ky��a�����K�̀
vŞ�|ŧ�#8����0,Y�,Jұ3O�<D��FdcG
�JUW�FpN'�%ԱK���9�@���5E��,���吚CVW���O��]���.�6D�^��R�eh}I�}�����@�^b3ު��ay��2�|�_�B���m��OoB�K��Q
�m���v������+����Q�~h��wI{���-Ru�M2
E��*Q{9_O>��7y�[���iT[���(Un���{EQgH��<
����G_�	�_�w߮�j��=�e���֨l���g��<|�����)q��流#�DbI[�g���>l���Q�F ��wW8����S���h�mY�m����K��\s��	k\����MK���@���1X���>q��B v�)����:$iWe�'�Ye�`���Y�@�Å�V��kI�"�*a�ݬ�ׇ�-�Il:��c�1��P�S��E��"!�rO�Z# w'I�<#���8�2`�pUlګfG9��v�[i����x���i&�+W��3e�jk�,����`}8Yz�z7�1�\D���O�~L(��_u���Iُ�#R��ΟC:Ce�*��i���������N�D<ު@�Ԥ�p��1��EQh���鄷���_R����ԣ�����-��e(9W<��&������fQ�'��^��@{�f0�Shi�;��?٨\Ԁ�8M��/���l�8�l'�ql1C��O.����}�$Ȯ�E�mV�*%:����w��e�3���H\z�u��B�M���{��ǝ�t��&�����-��CX�5C	^���R���~�R�wϫ�4`0p�R@��������V68r��2��nu�
��wrg0Ч�y�8YNR;X�Qx2("��+@���1"��L�+�#TK =���[U`I�lŉ�졵1ǜ�&�[}���h��ڮ%H���*U�!B.�M�s�L�	?w�����9H�"��5���k��Ϧr�2q�n=a��m}8!iҫ�6��ԛR��J��_�;���#�� �'@���}�Q��@���ƍš�[���G.Ձ��D (�"wg������$�;~yF+�gG���@\��al��ϲ�&��E�7�p]����C����Ru��A��a��\	����h�;��r�#Ќ��O��p^Z�t�����b�����q�'4��{]��?o'y��3�aM4�ez}�扳Z��&xK?��v�H]������ߔ�r����+Ah�N@(�!��UQ�R�.��~<��wF�ȗѳ�?�D_ETۙk���:��B9�̹�N����
����<5��<���W����v�)<�u��'�>ص�%��I���r�ыO�߂j��Z��h��8B=h6�̤Km ����b���Hi 9gG4�z55ܳW�m��!;O��m2Kp#�Fn��/U�3k�]�)J�|W�
Rnr��v$�W��Ú�a�\F��C4�h�8����G=y����>roH=�O��zK���]�8S��+d$?}�)�.R`6ʃ׻��r�S��3~�n=���Q���(D�x~��:;�ѶJ, �|��)>>�gsj�*�)I���Ü9��8�Q���.Av�79��8f�6�����.E����ï�� ���)>�L��C�%���d�p�%�~XS�ֲ�uU��k�/R+�1��|��䀹��Xt/T�5?�&e��n������Nk2��2���k����r$�	w��5���IG��[��7�D#a�{��-�`�L�-Kc�T��_�<i�vo�i���֌��^�]H`�X9�	>0��GP�c�tʰ;L�|��	�	�w�� \=��Ϸ�->[�b �h�7���y<��fB�	��(p�o:I�����zY��n*�,�A)b����t�'>ᇻ�K��������-�n�Z��I����3��%��*%a�*��6�����(湥q�W��B`����Ǜ[�_�-a�}�$ą�jrF�D������$�^��(?��-;�o��A@�qd,���q�>p�0���א"��V��OY���~o`u���J�+UE��"7� Ȥ0��`�FS4�mmB�pJ"+�Ƿ����vw2&�}�:� �zi>�ffWJ/��	�y�L[YN���h�b	؏á(�ƙ(GG���ɔ��@SA.0��Svr�
�{�Z�Z�� ���>3}��L�2066�f�*�Ҭ�Dɤ��oKOÿE$i�O�҉��$�4'چg@��>�c�5��Y�W��g�#��]�}�E�Y�0$:�.�R�m#�@���R){t�q��rSo
wu�QGN��'1
���:�.z���WR�/�\#O*��F�bv�c/�t���ԙ�:xOSpt�}Z��Ⱦ�|}sY�̘ ʥfF���<>�&]I*�H�{b^ꏎfr%�6�DR��Xy5iHߴr��a���m���5��&���j�r׭ɜ�"%ɡڋ��mfF�aa�#1�j6!������aĶ��]:tR�oHiQ��;�ٯNj��J��Wɐ����@����)65��Y~�44�F2k9��k,:��;��,���v�]�Dx4�#��%eek_��! �IEU�7�,���
���YGȀ����<�G?��� �����wx9Y��*��z�d���Fd�XN�랶�2����3���7V?�#s�({��\�Ea�Ku徳�p�͓6Ԇ�������%�G/|ߢ�6�s^�'SV�i��\\�Z��$�*�G�h~�����6ٞ9�Mǐhp�	�o��1�CK���P$���e�KR*�h��2+��!����r���y�Z�v�������
���4!^�����f�/2���P̊�Rj\L�B�,���,8�{+�ey���k��^�*k���g�<l����Í��+��D�G�j���%v*�XS��79��w�4Tw]`�%��^�Uh��ȳ!h�\���L����iE�]��cuI��^�C.����f��#Z'�2΅�i�s��ȓC��C,�
wbEs�%�dGag������J�9_Ty�k�0�ғ��[�jsAI���;�p��_�,:�yL�*�������������Rub|bI���:(l��x�)#�y�����o���E��"���Ī:3m���Lˁ�P#���`�|@��0ϲ$��:�$���H}���<
��c��/�XY�~�`�_%`�G��u������f��H[��)�t����?.l=v�W��XGm��0h�4�p�a�-��"�N�|�2��e�����G����ଁ��"{�_h�,\��>�:��e<�k�9'|���t=:m6Dy����