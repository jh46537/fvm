��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2�9� ��,�<H0	>��|�5"�!�n!�����V;5���JNs�y̠�4�S%ǚv��=�h���U/�+�*���C*Ց7Ve�%f�n@�%� c?�8c�Tu���ԃ���Y�j��W:-+2.٥���Z�Z���V�;�������~�u�J3�!\b����o���Bk},�a�8�jt�ѻvg���4L:~Y�1��̏��O��:�d�N��{<�F�2�h�$7(pu��U���L�t�< �Z�xʩ�3���Sw]8���y%��	�Q2�ÃY�Q+ľ1��W��N
\���H�F4q?�z?%�9P4%�}��vĂΎ������,���a��	��t1�Q𲈒U�AjP��%�/LV�c��?�䵾��� 6:*�Gf��6{����	�����N��
�
P� 0�w #�̋$ÅOT��#�3����f*�|`Nt�``4f�I9���NO�g�"��݈���g�����~c�oJ[�iLP�I�G���Лd��'��$п��%:����-2k��>��l��z������d��tt�i-*96�������幮��iu��&�/�Y3��y�:�黡[��&�����5�o�%�
Ki�Xk3]4*gS����b7�����+��h)��޻q�Q�|<�7g�������/��hL^�J�V?��%Gbp���CO��{��fL/M`tj�� �E�D��N?���a�әķ�G��8��qS�ʢXې��}<KO�),�0��H7U]�Tn��u�Fɓx)�� ;�S�z��qpm��15 )06?""��+~���E�ؙ*'�nA�BCe�� �!Ғ��=����X�����T�s�j�4q#�]���]!N-���T���!����a��c�M9������հs�w�����N�YG[Z��u��6���Q��Lp����i��0`������|xK�=Fn�ܱ?�u��fAK�z}uA��B��:8*��/�$
|���X�x4�X8�)y�HI�X�F�I���<��i��GG��hSǣ>�Nt�</i	�|�-�T�vg�?���˶ZZz����V�еt�x_�+�1�0=��[��M"�c-"E�� �fn�xΕq��{%��:3l��VF�3���{���9��*U��c��9������[��z(�C�8��h�Z1c�����)؉Ͷk,A	r�z8q1J�D��=�����5d�4U�����]���(��S��Ķ��U"L�*T*D@p�Jo�.E��u�*M�����Ғ���~�)h��c�0����
��o��K���M i.捃6}0^u���
UY������~�+ʃ���Mj�)Ć�(�DJ�]�o���c�9�6��G�Pa>Ċ���.����W8��Y�:dY�助���1QO����l��B����^,�99�Ѝ�ԝ���������`4��c9��Zop�	�b�X���(i#zWJ��-B��ZS�3`o�63��ӎ^�4�^����}����0y^�"��M/����a{����R��u���wȪ1+�����V�Q
�\~�fủ�����q�X��饒C+��P�oّ�sxg��0��$�=[� �,Eǉϱ�n�A���y`HsApu8�~+H�	�f� E���1zo��ѼP64�*��om�Bm���NRk�0@ۨyX�ʭ��G1��:��r�=�m�ߚ�F�xsF[$�Q�Ā�`���C��Y�����v��p���Bc[
I?[�}̖�M4��J���@��ḧB-h{j0Qo�d�=�rw��bx��%/�b�Z�z���/�''�P�bޤ�JC�������#'
r'��oGo�*���\��ʣ�1��9@iˈ:�EA�l�m���d"W�)Qf�@���n�(�6�����N:�1����6#gH���i?�R���'4x��7��
��.|]Z�MdV�T�^��5����b���!�J���O��txE*%�/>P�f�P#U���U�x׳KKGH�z��m-C���U�<�K�E��3�&���IKŞ��=[�� ���,���_}���Fnq!7��ABs��x��I�4�����*��R���O����,����%��P4_�a|�`�ۏ���R�@�P���9�c~J=d���/���0��jG&@�e	=�!��Wt��moKV�r��8��(��^+��u�8t���Ǥ�@�8�ٻ��<C��`!ĚB�	v��{�PUE��;�����~��{�Mi� #k���(M�BK2U�$Cs��r-��?�Քr����q�ܾ�D������L�V��k����μ9*J~W��s�Pw���|^�� �-lR�dY3����ِ)�y��-u�kM�G����"�~v�c�W�dus�H���m����ZA��AKه�d��H)cgq�)K��HΦ�ͬv���?��FE�D����x�:�	�E^���x�g�\ʨĝ�S>�y���J�X��+�dp�/���z�A�C�� w�V��WV�U%1��a���X���#	�Mc���bg��x�m��P8�$�;T�B���ct7w"��½���q\�z?k�6���l���4�����Y}!I�HBb&M5�u/�2����D�m�|2�J� �i�G��ߗ�IZM�\@�g�e�&�=H�V�֤���ە���5�,����?��}��e>y����% $1�vfw7F�Z0:&���M�V�����'��.{t�nS.{
s�c����e)5�-��fg���,���cČ�.Zc�^����hx�==���,@��OJ��O�K��	+�3�hT�j9=	��T6���91>0��Ք�^�6VQ��_�<��Ǒ	{%Z�{`��L�CƼ�A��5B�I�.$IXO��`p̈+�~��GY�"�W�P���E�WІ�'>�TW+u��?I^~L��\w҈GY���y >��-��
5J���j�6�(�_e[����pC�tK\�����h;A��`8b��^����ON�!��^�.O��m����'ُKD�E�����K�H+�v�AM��w<T���~�v̯u@��h@��e~/ER���J��)�0�i�R]F�|9c����a��>�!B��.�pB=��Y��C�<F.�YA�1�����.v�J���e�í�L����уH�J��s�e���r�jn~���������Y���|��J��7��[��rY`R�̽�ğ�n-�<ψ_���Α�D  ������i�������y��T�xz㷞OY��?�}�����Q1��Ĉ�?c�d��d����s����=�r��4�dٙ	�+*��p+��X%>�� �&ԡ�2l�䬂�h�p���`6�k|ˈxI�>�*)M�)�1DZ��B�[U��?�`+���w�))��_1�����_�4#�f� �-��DRZ�Qj�	Ӻ|���Ɏ���x��[�ZpkV7��Ǣ��1����E���O:�w1�qI%0X���c@
e�1��8��GR�h�i�9*B�G���Չ��J��	�FK�9�r�Pr�NQ���g3�����2<T�k炄MO��c:w�ͥ��b�`(o�����g2s%1@��5W����*���T��7��A��fe�����؆� InC|�n��M�v��R��e�Fp��8�%���a,1�*a�oxrDQIZp\�D1a�(�o���:>4rU˷��^O(�Cr�ď���3�c�A�܈�B� z�n^���A�NK�Ki���;(�H����!���	�����uWH
8u��tZL��i���<Bhnz6�G"�i��e�)��t
L�)��?P��DyJT�%�j�v�a�<!�{�N�a9,�$!�;?S��_��
c��yɡ-���I�0=
�^�ӕ{�_�+�Ft�{1������ ���`���IN',L�ٗC���t��	�����q�鎳��ϱ�@����E���u������ؽ\3�$�M8�$[p���dK&�0�U��N�Lbߝ�ƭ�@L9�Ǔ��z�~g ��a� u��kp��	D�gQ�1U�{wg�x� ��H��y50�/{6;셺޸�*���1�2�l���v�[ri�jx��@|o�Xcl�j�i�y��HM@vG;�s��]
9� ""w����$(�����V��P���WNy[C�3�h-1�ShxفheSUx,+.Y�uoҎ�[ȭT��ZJ��a�k��F0 ��vM��=�j�������@��PX�5O$U�?޽ߡ�rl�Hb��/�NPX��ž��$���\�'�y���~ZDLv�3#'"�ڇ���������� s��9tȨ�%d��ў5skc_?��g���XY�+����=@���h>Po��
ŉ� K@ �a�G郌1_�IX��ĺ���@��[��$�I�v����Ipnl]� 7�"��M���/����1R��b&qi���vb��Nr�wFݳ��G��J_z�������V�	��	��XU(y��lL)H�����p\ ���	� =B ��/{����LAX�G�:t���n�t�q+�z�� ��尔:��kl���U����'Q�[2S���a*��s*�+��fr,"��$�RE̛]�٪}S�o*��������Nx�o��ڄ��5!ͼW��%�O%)N���XO��lk(tGO�(��K��ɽN0�o��MͼͶ��9�����\��g�d&�ӗ�Et�4^9Y�X�܇�=���9kY�lSxY.��=�T�.�C��8��L�֭:^��s������]K�N��,q�R�:e8��'��e";ߠ�p�[!�^�uڛs����o�W��ta)���)}~����ׇ��
��=�u�����r�� ]d�أ��j���*Yۀ��W�g14hQ�~�;�ٍ��~P�_�՞�e��6�#U�7-gE���*V0���G����CmX�i�&�6�X���E���4(�ڲ��F5�a�S!N�S~���`QM�U���ZY7p&��