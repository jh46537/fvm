��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�ӿ�J���I43n�lr4�J�<�8��  �@���|U��5�����y*_��sUe��[�;T��;�/]��<y��#����6A���s=���5��C�_�v����KZ�r�=�Ĝͦ�/��|,��E� �ܢC= 9�D��]; �K�k�X��3�9�Y�:z#ޖ��!�����r�i�����G!���ƞ#�Dw'�����\2"͏+w�h�f����������h?_<���E6ߺ��Ke�),��j4� �:��3}�1���
�H'�C�m�:z��Ǿ����I7Bw��05�zpv�z����u�L{�8aP�-#B��c�\i����y�F��@x�H��z�k�ʔt�#;,n�RE�*uu���R��e]����-����*z�lV�hw𒲙�\�hTom�5z��ϳ:�M��Ȕ�?�>ܡ�����)�a�8�x����32�8y_�S�>ܿ�F�,$��	D���;���8�͙��#ݜ�?�cu[���;�xOJ�o|�(`1!����➈�=��к��
xXFəRZ�NT�m��/q��_$)z#'�p�9
�M�F��`;	�3�>xF���l�u�l0����	�-k}>]����J�t�{߀�i�㕻��w B��	w�s�q���N��ը�I}�6�/Ҙ���:�b���O�L%
��,�̎6�;͟��_�C�;}V}F9ݫ�Xiz,&B��
)���i;������)ɛ匵� ��������ͭ�i��ݰv\5��f����~��'W��Fc���v�{Rќ.����|���{�GXңr�E��6RT?�W�Py�=��0.��U0 ,؅�1S���qWq5q�9W���=�� wd@t�W�n
zF� &a�o��B�-�;�Gj�F�]���oPs1���L}��00���I+x'��+c�PB��bo]�����*�|�8�] ����V��5ʰ./y���{�_���B\�G�HumBU�f�[���/bo����ix�KK���7[*'K�\���x���R[���NpG�u�WY>=�r��LI媝z�zrv�^��֦r�r6�	33|�e�d��8�8kGH��Ie-�#o���(G��d^T�F���	}�'�)V9���<��y�m�#�6�7V�S`іV�_bg�kg��+$%�/f37�=o&2[C��'�d���8\g?ȹKæ!��h����{����@�#pG���\�`>��k�Z��(�7<b�����W�Nvt��k��F>Ľ��uM#�����e��]zz6ahR�ѳ	�듡~A� ���qy	��f)�~�l^�B�o<��穆�}���LZ�s	v(F�b
0M�dU�G��j�S6�!��i:m�k��˂P��܂ʍ�8)����=�?�_Jڄ��x0�VƐ�W��޴:����;��b'�Wl:���\�qa�^L;��p���ЇX�;��AXGh�nF���D�^�2�������m9�D_f\����1
�����&BС&��e���j m��u�Yo��7fĳ�7� �T��[X5�oE ��Y��#�8�j��*��]q&Q�2J�X����蝩�}�KN�z��O2F`�.����/��#���9�_ÌM�&��Cwj~P�L�g�' qۻ�t��8�=��,�&g=��@܀
(x7A%���[��$���/��W��R�3��cx���
9r!'�4]@ûڞ�2{���;�!��Բ5$G}�@�go(~1H&�3jD�E�ʒ�+@��g��F܊98�3V�|z�3 �k����	�mIة5:XrĽ<�K(`��܂y�]�n�Ř6�ݛ��<I�����0��V���>�G��Y.R-biC,ISm��F��$���
ϰ���#�n�l��>�^^+5/	�2r�h�����Bը)��ڷ`��-��UD��;C�̩�.M5��c�QVv1�d;H^�I�Bt?��%������]Nh�Nxt�W��S���[�����sWy���/:RD��\��3�ft��T��p�ͳ!���=�]Bx��}|j_+� ���'��qZ���#��z�&�SA����Oo��~CˢG�^�w�'e`6fh�}Iv��:�)�-TQG�}�ȑ,�˶����}����&t3+l�.u}�i���P3:�ԱI�XX�ƿm�E�JL������^$�*�T\}E	NH�T'��9�y$)�d����:�Y>z�c|����@m�w;���؆Ĺ~��A9H{����X�++���������>
n]�+���P��h(;A{r���AFC�9��F���Gß0�^ڭ��e��gR��� |휐����i�ߌ*n�ٝ1�{��������!�=[�L�J�Т���9~y�>3�R��n��v��\�@�8^��ݔe[��v	�&|h���.T��+��Ο���� �����t�6e��w��Ʉ/Sr�m'[(
`�]�#ea�����:� =�U���E���7��AhV��a�#�h����9-(�	^�˭Y��7N�{�>(U���ک#���#6�"�a��[v�y�4�6\t$S�G���C���Y�%��~��u��~�Rل�*�֟���˞"5G�r�-�<��2��i/�60�JtbY�wjB��=�yR�&jK��˒V��[g��^?���T��|��U��CiǞ���5��S�����j;Ʌ_	{ ����|���,�8�$z���}ꁂ3t4a�In�23G:�3Q��P^����Ϻ"���k��j�S5\yҰt�	:��+��^����Y2���T2DY(N.k��Ȑ!�R����5���>S�Xs,/.���9W#���X:�G�oڢ���xC:�<�޿R<,�ۦ�v4��7��tx6�0^�"x��R�^ǫ�	0Jƞ(|�24x��a�9c�ֽ���&}���Y|kC��r�0��m���iq��,���3{���$j
K�=}`\Jc���Y*���)��w�\� h�Mݔ��9�ͪ�M�Nf��j����{��Ͷ2����e��o���p�j왧�b�9�N����(��1r+�l�}�<e�~'��4DQ6��.��/�=�u���>)�Y��+��䦢��K���D�(����v�2�	��1�8qw$�oz�^\��P\�)$e���Vx J�j[�9���/���<�AX�n�[¥�w�U�d�-cz|\��ԩt�`݀GF�Rk�CI��|��PA�(�sD01e!^�q��g��=���4��28s!��%L)���d�4�E�e*b�D5�5���~�1�$�W�srJ*;�GE`�L[�Up�*9��$W�i��IP֠c����+���i��b�#��1I��}�ئB���������Σ�x�a�Ʋ�$����Ŋ(���[h>\��C��
��˞�֦��o<bĿ&rsDQ�
�:�A-v��$�X��Fr������fg��h�M�L���1na$�����vjp�!%���T~����i_����tv�\���8��f��?�M��:���aҍp�eo��4�[6J)������o��`���H�ܞ-Wb�0���ɼ�Z6pe�봇A� �A?�8K	���;0������خ��T�(X@��1�5�Ii	�+f��>�Q~E��r�.=E�o}T�*�$0r�Ӈ\W����H܌lP�A�L�FmA ©�P塚��a��(i{��{�΁�=(a�(p/VCY?���oS�鶇-L?~壁�p��j)üNA�mA����ZA�)2��m�&9Kv�K�P\�\�5MrG65KX�^S���I�T�vA�#�,��.���Tb�oT�0f�����;���-!�eJ��Ջ�e�.�<���J�
��U��˛��������a
b��E����+V��7���	&4��?]��ch5�g9�/�$�) 94�����JDEq�O�'M��fҭ��s{���ډG�_�� �!0��(�ߴr��!�֞���D���{�k�Z23�a�	]Iۛ��_a�B1ȸ��U�",gV4�QZ�sb8#�P2����{�V=���d��n��t�F���B뉑�H���>,	t+�@
"Vc�W��@��.5Z�tr����h�S'��·��4��צ��͝\�'CA_mq!uu�T>�E�3�u�lY~�4~^�~A1��H+���c�)f<
L�m5,Л�N�N��'��X�~i��Q��Q^ݞd��l�)����J��O�-�xp���m5�9<���� \�-�P0�u,����yy��+�@�n�9����ǌ_���oS�p"�ʱ.��X�L�M�Rb8�+I.�Dk��6��ԡ9�W_�."�.%��:䃄�iE��m�����>�.��b���\���N�κ&o�j���
���K�>�D�tN�������b�1��;-t{��`����3����x��`JzAuJ�b��vuN�xt�5����h�P~� ��Z
�^&Q�_Z��呿����|�Q���k��g���(�I�+)��VPr�.�=���K��N�A�O��Y�}X4�֠}��8Hgh�w����:��iQ�d������]��s#]���I*d���Q*r����@�j���ox�A3��sln�d����#�Z�x{�t�;��6 Q��X��U�%�
A`�����ƶ)0��̦��~�
�N��?�t����o�Z+��'CKNG'ew+�5�A4\�~�Hq���	�J>Zx�����Zn�:,��R�w��XD�OIa��8�p@�FVWj35�xU牳�J��cٟӶ[p_�¡qgB�,G����瓼�b��T������:�5�q���Q,�I�iNyF�� ���R��S���W"M���=ڶ�Ur�mD��_��!��n��N��1�UB�z|b���7xo�U�z.��3e�k8�N*� ��[���	�'���A]�\��p�U�t��9�.�sO��g���T�S���˗`L;��~�y�Te�i�A�惡Iov`=A�Y�}� ֨<(IZ�
G�g�ָ��kw4��ś7��]�q"�-�Ka���r\t�8�8>U��'P���*����I?��/sA��U!ぉy�J:@@���)��?.�]]y�DJ[�FNF���v���g��B��n�^���w����n5����v������z< �ߧG��8�oBcd����$SF�Y:.��Lqk��b�������|��G"%��$p	E�@�ኣba��XZS�Ӛ-��V�광�m���l$��G��Ǧ��l�W&��UB�*�^��}�ȁ�L^�~�b bԉK쥓��J2�.74�������� 8N�ru���<y�Mg���4ɱZ�7�&�9��m�_��h3VQ��G�V+7UL����u�E��Zg�~s���[oۆ���9&���Y�����v�sNlzC,L�Jp�W|���Z���hw�	E�A��D:ٺ�=�!@�ű�$(_��K1z�V�-r(R=we�խ�27b����.�u�'(��L���Dѓ�ۏ��X���z"������8*�+%P�ӛ��r��[C�%��zȨs2S[����u��q�h�]���R�H�&@�{cc�z��ǹ�8x�D#��e�<J�;I�%���'�2�C���d�P�T����Zj�y�WԢ�6�u�&3f"ִ.M�.��G:���	�����4�>ĵݺ�7?={��I�[��V��F�x�.�~��wnq��NJ�o����rJ���:����`�Vr��G��������~wA�v{݇����*�{�Φ��"�>�O�>�ɗ�O��sem.I��}��[���}��L~����0\#��;��e���Q+�ٿ���^o�Zi4�s�8(���-$a�*I^��Ġ���ge \_��W;�H)�l����_�oh^�q�l�����~�=-�t	�t�Y?�{|)�3��8�g�Ki��)��P����Eih��nF�O,`�R��f��x{%9��4�8|�Y�ޙ��wZH�t�q�	��F���/�r��в ����戞2�N�ү�|5��8:�j�>q;��gy� J�ڗ���Y�#�gSr���,U6x������nm�Y{��I����z< �0ﻀ���M����B+j�I�ϊ�'u�a��[��BD����Րq�b�83�W��D:�V���FS�6%|�/M^��H8�"'�:���ʢ��OU@P�Uf�,�b�0ˁ�e���S�u��*�=&�V��^��ӯ?/܇��מ��i�{�S���6VA4��oH4��0�ܙ%V�Qޙ�	u��>@I΃4�,�I=�M�W*H�\b��z�`���y ��Y�?� X�&��s�$"t�KvD�v��������<h�����g7����ӑS�Koݕ���Mճ��Y�CE�g���e8�C_��?�Z����S�\J~�ci���w�=L׋d�q��=~i�)g)&���O��>���Uj���퀈�9���@��haL����"��=c`z̺�`C&�bl/�����w��be�����w�W�g#�����2<l��LJ�W��LHީ^�8������w�<�M7��ܭ��Pg�5�Ɂ���:ϡ��� IZ�f���L+"���+�ģ��N�����!c�m���2�K�^�I�7�8G�~��.;�[؆j���e+�`ɇWm�N�'�q:"�TZ/oZ����(8y����{������xM]6b�%e�6m�H�-�`*����ņ���X�/���Y��T�-,
�p��v�2�I��`��`��O����l�LP�@ސ�w̢�Kp�V��3�g��lQ�kM��𭲘�U�#a#��ߧ
W~�b���0L �L��B��@�&�0 H���l��#��|�^�����۩`C!��[��s�i�W�(��Cm�梒���������y�T�糧�B�ьU�j%��)�aV��(�a�a���>r�!H�y��}��/_����h�8��ۙ#ۉn�)�����a���JI��)X3y�1[}�ε	�����[�'>a�x 6/ĉ�Ck�A�p���s�|��4��!>��0�S;~��b|�{B2Q�`��n	A>N�'�mꋒ�V�o��tp�TNV����Ą��⸪�� E����O�!Ws`�62%ؠ��cz���ψ�#²i��^fK���*�����I���/�tm'X����~<ϧX�	!M�9���+p�8�s�T[q˒�\j@��a܇V�Ȱ*�j_~�rH<w�L��W�ү~���ā1y�8簯ࢡ;�+�n:���t���;�[L}��Wb�6����0���T�l�ء�˕��*����h\�,6���TQ�i
6"�,�'oȡvi�i����;ը��v~���	{Ȥ�Z88����'�U��￣�ލ 5��&�5��|������C���ھ�ЦQ���:�5�N�����E0��Pw��/B<cG�ť9�O#�#>��Vm����	��e�d;��Hn|�ǿ!W�7\rv3>_]A��2�I�Ei�v[�}�N�8`����SSåP��d��$�ĥ���Ys�2n�L�zX�Z�u]�?�L����42�<��u�lw�d)ٍ5*.57������v^�N�F-�'���j�$eF.Bg�b-�)	�Mů,�/'f_�ţa�ޒ_,��n�+涾�:A%/����~� e�X�;���A�o]K�`�X����~ݗ&�!�c4`r��)���/Xr"��cDTx+Ņ��`��KJ'�
O���Z�aU�]M�^Z{�_�ʦ��
R�)�q;�&�/[I�̆�Z
b�g���O9�����Q�m�)d�N˧����0 )��|�܆ȱ~v@1�J}asJaA�~�BϠc�ʱ.�gG^�U�=轰�s��u�Ԕ�r�!X��q>Yol�=&H�"�\�Yq�{"�lX�'����:<Q(�3��ls����a,W�~CED�Kei-"���V�R:�W��|W ��<6�����u�`S}�Ŭџ��Eu&w(D�^���t2��'X&���� �u~�W#���鍻�1$�%T�71�CC0����o���LK��ѹ�(,D��_�
�*}��� <��HGb);�U��G]�u�vǘ	��0�d,E��񡫏��?���K�v�y���
;���["�_2PWA;RL�8���'k�9C�c9�|��v׋�v�T�'��*�-�e��e\A��@/LO��Kc�����A�U4��hwoƩBD>�5�2�s7 �%|��8��v��,���N��h���!B3����S�^��z0<��gݠ@}�~ϧt� Ǭh�'P&�wY����2�Q�H�=ȉ�q�O���p�G�~��p�p�^��7�X�c���Ek;�d�_��-�GOI�0cO�����y�3z���������m�8қx@��+{��Ϋ���|���pQ��`��:ȢƆ3��	��w�<q�cs���T9���$R
,����a*�p^�T~bQXҀ�h37��@�f����|�g��D.X�{�#s3|��7R��v�i{������}�n�5��V�Ά����d`��)�ؚ��&m��N=����H��"�����.c���P$�M�̉����IבH�������S���"��45Ƒ�����[f��.�������Y[1m�"�.q�W���9�lK?l�s�����pp9o�0H��hŨ7��vV�L��N��{�05ڗ�?�O�_mD���?����b!>��N���RÀ�i<t���=r�2Tw���s�k��´+����ҫ�i�ۯ/X����ֽ���$��촙�F��v31��M����������A�o�u�����[[�T��-o`<��\ƨ|]�EOf���{�r�1��mm�,�h X[nD�Q�5��>�EkN���$���� x5�I��0�dur���F�Y�k\z��<��?M�p�kHg	�t���;(&�f����0npb��_Iй}/�W*��<ݓ�a���>;�P�~�]&y�9{Y���C������'�����G?�K<��+�gK7�7���\?:f�����d�ET�V[��鞨�!��������J��Ҩ�r�M�s	'��"�_a�F�N���/�H�FG����'���t�gX��z-87�q���;�a���h��R�f���n�EL�-*ܮ�gq9�W{�t�ѡ����j�5��0p��*8�;۩b%ػ�k�\����#\OR�~�kEM��!c��>7>_���^8j���F��il�T"���GR�OOU�t@��~f�v�e��T�#RjGts�X�!�G�;eLG���zT���߇���?I��V��������J:���۔<h�I^��*����cK�?3qp[��7�U�F�D�����i�#��Ts��E�!��+[���{����6�|�FO.�,ްV����cC�NNM�I��,�/%��Mj��R1��	?�H-��9�����'x)K���4w��c햖��(��e��耗�F�b�c�a������PX��&��k{�t�9^��"6�P�Sq��Z�7«̓M~'�bݽ�ْ&V���I��e0)�\�"|n��Ͱ+�1�̐�#:�%{�q��i
O5�zB�Ky�6a��^�`sCq���|R8�$�U<ܢ6,�{��x��3���. ��I7�Ś<`����S6���������-����u��#�?l�n	���wrt�9���>������4�%�v�Sg(݈�x+�&���s�ߗK�4��j(��Jbq!h�%uPJ�6�}�.�B���w��!;����'����l��<F*��`Aam�oo�X��A�<"W�����).����5̛^>F�K!��(s}�>ū���Tǋ����D�)��a	�蛘'U؅�,f`�4�P��XŖ#ʬ����rb?WH2g���_mB��-Z%����H�Qh� κڰG"���6�sV���w�-����9:�Z]��1&�އ0�Ť�M�@�F&�C��j��7\�;鑤i�ؘ��,�W5ˌI��~����,�p�Mb����š���>�ߩ�@9�"!�״l.��(_�k��M�N5�5��U�F�ág��E�������Z�+z�A��05.YqdG��HEP�����94)G�+{;���`���>T�,9�vT�O�a��~3��d̮)���G��v�	���Z|^iQoUJ$E�xv2G�,�OO��!WG�qR7��폤C��I��Z�����s<���E�5���ɳ���vv�T�%bv]�h�e�KQ��~�2"���m��?�Gw󹚔[Rv�a,���h2��<#��.`#�Ң�,�������t>]�I�_K+%��u$�����F�i�c�_�*��T~��&��Aw\S�6҆�r����b$�\]bt�I���+a�q�j���Z���/�`m��b�L����<a&,dc�_���PaT1?7./a�#Ln��\ش�+݌2���MY������$K Q_�'{������\*���͟���2��)���-�^�T�H����>
7rO`�a�$��mcp�X`�ڲdo�����0���$�27Q)��^��sD�=�D'��p��Y�$r�.�@� X������"Y5E�z����@�C�h��j���0�j�L�&�C��i��*�?+8}y�����U���:��h��xa�\���^R�݉��=$c�}uW	��T��q�5��!BٳX���=,P��q$�pVx�UD�u������X����	��Șx.�EVLb�x��6c��%!+��;�`��b���G�;6�2��Q�G
S�������>�X|R��c���Ol�4����0��4�����o��j��t�@��2�5\x&�%�ߌgv;�hr�'q%���J�b����ԹYE��^�0U�Y����J��h�a�+�}�*��o�N�I�MON �G;��h(�H[7�IN⡋W4F�J��<\)J[!�	����1��T��GʳN��Z+Ӟt3�O����n��QZ��R|�b�!��M�S�O:��Fq�k�YjH�HC�G��L��������.�zJ-�s-�nJ��<����M��G��dW@��q�Fg�V��\|���?N�z�=��y]>#�M�_Ɣ���C�hV��dTg�tg 99Q��e�,��w�ݙ��p���W���zhja.
�Ō`�Q�A�.m�ױ[@S���4�~��q�t]��/��f�	+�Fp�T��E�;h���_��_�-1`4�-��th�!���á|��ů���g�tU��~|^}S���aLrˇ4����v�v��8�s�!+p��i��xf� �hR����(�ӹ�_>N��J�ɜ��� ,Ƕ�;!6 �L�^&�ۉN���<	Gd;[�%�T;�U��!ާ��U�!A�R'(�&w�K��bS�hH��Y��/!(%�2���q�< ʡy.;	�2bZR��ebZ�-��M��~�3��sd��', Z
0�^G��ܮ�<4��+�|X:dF(��/���X�Ǣ1p,ZSO0�%X���A���%�ae�`����t�.��ʼ�>5{��T%��o�z��C�LÊ18����7CA%�V�Az;xL�)�R�\F���e����D����D��I7�&�:���X��=�*a��.�m���!	�Y���66��3��G��`�J뮚�5��-7�)��d���߳C���0�EI������35m�qGW����M����F���w���*Ûh^0��,��T�|� �z�I�˲9�GF�`��;N�R�%i���C7Z@��&-H�8�* �V]����L0��,� �b8����i�Is�+�h�0R��g�qan&\|s�p9��h���rsGD���#��`�ZL���]�� ��O�Ζl^����V��b�	a�;�Mv¢�������j|%f������'��z�W��Gg�&�4ӑX�AxMh.鹡!m��������DЂ8��w�È��y�޳7냭��~��v �,�|n�����ەЋ8V�Vh	JXR+=+.�|nQ�'G��uM�{,�[�!t�>�?�FʖǱȟ|��D�%�Q��p�>���R̛���~II4���䒖N}�cH�c��6��ۙ�6:�Q�!�Vsqz71��*eq6b{썀LC���!��t#��#�/�.3ke���NSu�>���&�\q[l%u�9\�Q�{4.cO�?Ym���k�����e�ܖ@I��Ų�m�Ami�`���G�C�t%�S�*��)���<D������2Y}gb�'Ű��T�Q��er鈅Z����魶lk�6n���x���i���A$��\3B��*�>h��\��!�#oNmQm�>%b'?|���`�ȡ _�h}��Q0�4�9�9�@v�VxbU]�eZ�Z�}-l_��]�-��x�t4�����BH[Pn$���I�4�k��9���'8��s��I�y�%�SL>�dA!�f,g+���������@�dV���s�������j�-�B>�寣9W�?�X�T�=�:���" -��Ks�8s2�|Ԙ�<w��Ɔ`��W	7���<�G�.j';���_@ةM����Ι�X�^�}��0�bba^$Kb� {�j S�5<���r
c�j}{����6k��u!��rL���r
ߑC�YkPȋ�^��[�b�T#J�%�G-��3>On���2���˦%"���ןoSvT��I�dѻ���U�TJPh��@@����O�bh.]�W��ϯW5i0q�9���b
@�5p�M��+s�wX���Yq7{�˟����c�����'O�_�;B�SY��	C�i����~e{7G,� �^��zq��4N��"#B�6 Y�2?���.�e��%#e3H�����L�10���T��]�I���آۉ�l��ƱG0�J���9
�,�t��
ꉦ6C���_U�$?BFc�R�Gz0�b�'�	m<]�jnRX��G�R�mHr��N��oArRDt�,��QlN��[�J=y��S��CLtx���Ɍ��Ӷ�@���H�٣$I�Q���G��#}��������e��-������gֆ���f]F1�9
���ic+ ��n'��z�_A�$��+���8��M�+�,՜�ԏ�D�O�X�s��1>�]��N+���f�_b�\�UБ%r��l�