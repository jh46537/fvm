// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:59 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eFGPZc/ReXlwaeyKusLRDXh43XsETtf7Nc5AbokSKViBaNZiliCeobMYQxCI0cem
MFaeNcwvQ6u0IB9IW07MBb/RHNMelN8QQHy9NvP7VhUKSeio9BhZ9dZd+FFQDo6R
WZe7mTTpflera5X0c0XCNT+ry2OeFA49b3qmdxCiMWw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12080)
MzrMG7uuwgtegUXa9xLJRx/kJDFMknRD7H1N4MbGkfpp1UwUepcaaq69Gv7CnDg5
0kNEz9pxb7bPjUCQBPfctFZL+YpzyvhGJxuCzDZDlQAfPoyoHU52pbQLemrVmpe9
1gTrX8XG5PSdoUswf7tEyALEWqrx2Yj/vaj6KoK5zftKV8ArqLkIcdIc0IximVZ7
T3vHpccTNxArIUFi4843BUWqhoxoqs6UO1njaG1XJd24HD4CRYk9zn3hMDJL4XQ9
D5lEbYniZDcHteOkpdyjZlhxOLDPBdPSGFfW1bwYzst8hBvFHPlVLFzzmZRKWKRB
JlT73C9i267mEAHchLzxJBwe18oYdaXO2UoU5eaEqzo5y+gc2B5H/25KEJ3gTJOm
5nACMM+fYE/ffFjkzYby82rYPia8ZCFOV+hFxPpOc7vKdZFuBhKQ98IBCT8/TBHh
lZ/XQUI4MGf3CjrYdgOQzDfp3Qllve4p7hpDweISrpWa+Y0PkjNABGgSp36hII8K
cPiPxo40agnHA0Lnk/dQOjwiSCZx9d0kKBOxP57EKuZoUFagrkfT4KgmwfwHXJKJ
7QRRLN97nrtsjvGPUqvqFwaNxvkaDMuTYehD/A9o8q0nNvZT9xV1TJihhmr5TM7T
kq2ybwxUJOrepQbVLfvIeiCQy1ivPBv/lj4yb14GNCJ658sXWM+3pHncoJlyFxcQ
FWiYRnV1qI3isTCpNeMAM0jDRLqGJ5nJbtfT+VST2bpfGKu2o2Np26tLJbqKFB3P
rv8oD8mtBo+XIasEEugXgbrTFZz4jcjnl3a9aDXxWhP3kF6cSm4ElCP7YbIacS99
IIgr0++htaTrdgSAk86cisqzKsrewJoKOIGp3f2GfQ2PJjFiMhWAVIO4/53aHNE+
KpmMoCxpq0/eHGjmjlMfFOmDPrmAc/+h0Zm9w93ranUc/OVsxeL3VdFkB+wWwM5p
THamvu7+6YSo4Dvlos8DKGuRBfCSo5zixQez4P7EHhPmI2Pf3U+VGjcW6xBFZvYU
DLnhdVl7NLdn6+K2r/NId5pF/L3I2XsILHi7ovJX3vAE6LI+pcmx581BXSRQpp9N
SJBEFFWHlWg2VtF3kCVrRGc38EvatoS+ASJhtQ80aKBYi0z6EThLjww7H1A7qu8e
VxZvW72SZVLRM8K6mUgfVCbXhjroxlXE530HvBzFsx6fRVvbEvcc1Vw5Y7LKo+aB
Q2sOUjgh0oVZY46prv2zTvYsIDCjXmQkesSxeVJ+FFNiAbsIhIPc3uT/0lJHebIz
mZR0yTfy2pUw7L4/HUAeYPa3x49/udyvNWH8+O42AWILHP2eVKCGGVKM/bkK7O4S
HLEmJAz7vF+yqbdbMm5b3gc7AO+39z8u0mDNcXcDpBHphMEvLNwC4B9Vfo2/+qI1
yNAnMkgjACfPq8VcZYDDJLyHsZgXLmJ+e2C63hWOd64/DswjtcHKKda8qRrmHt8Q
mfMDVnj09mj4JhTRcSoYf2WLKkQ7bliqfLqTRnc5tHABNg4MjAfW/mujsFZrhaw+
DGeajekFs/mxhM/ox7ldbfQeoKMVmSfH7/4yZyFvPamZW50H7Zd9WyisUo3PLhNG
e7fU3CIfIlrbpPm5rgeO9WmpM9FMssmraJmXjRkxCxFwp+ceViTPrHCj9FLLhhNw
hmsoq2ZskI82kUFEvnBQ1XAquasCPtnggP0TAhkm8SYSrnG+Vl9ThnvjtiTx0z++
iNEp3qgU9va3BskhvdqbpD1LiuKioEz72m/9evDp860LTvErl3V72/8lksrxYR34
i5EVvW5sq2+szjCJ134Z+0/PqSX29l6cMK/Y1x4ZrQBZeaiMMlvJ9XX3i34rVxCg
VA/jSpRovCK7BtmWSKRBZEPxP1fHlsZfcyPv6Ebu9okqD4nnqYVRhBIa+xWSD/Ty
Oq+wUu6rFYT/jwJmItkzod0pmOIFRTJ//KtKO+KHSWDaK0RXzAUSxHLIHH9DfCjI
pbf/udvFcYAV3Pip+WtbeevUy/ZJblVmhqMhv4w2hTpOAhyCRu3DO+dt2NsIphlb
Dzlwue31mbMbksQfRntd46hkyNhDezIPSwGhEQLuep7G9AJ8nSRz1av7wT4A771c
zvvEMzVqJeknAyqxtdz21fDkKyW8y/SGbuZz6KcGoTJpgw/WpStGh3rL5kgEC1q8
iWkiVNmq+3juEXvrXFAr+Qr4/H/kZ+s7Rz81U+32ekIDATbYQhQ/TyLs+A4GPp2P
pH7VpmB3fIlzpZ0w309KOp+I81DGq8FNVKwtjjzDgD50aqL0jtQMZwVGsDFpOZ2b
Me5N8h12Yo4Lv4JCWnD0ttU2HtGcOBiZlo8pscZuQUCWKgu8SQ97AZbx/T/kHfdE
CbvD7NmNIHWsl5z5/qGDrKJx/fJ2b2/FJUO62AJEZXWXPKRtqGMdSgO0s5f9cJ6G
dDbOCsZ33hQjDt5xeUjvsoUDkD6j96rvoRCYj5wfVHf7QkKy3SzSe8phUl0R2PaV
EeOZJ0WR5RsGqhJv5dNqNFGRhY69YMT2LKVY+VDQfbOs6wnXW/SUCIIDaWHdKFTX
fFFQ1p2oSHwuylk9h6trZPBsFpoiKEibKkinG4/O+tTlUpJZCZpuLzjWudigjntP
s/LLb+nH4nnuFRn/S+GMISadq78Lu8KxQ0zMpqLQu7Gxu21zwUH343zwyhuc0YsL
PqTPhc+vh+sliGZiJPqPl37omSxvtwWIhrfCWdeFquZXnwNmxB5rTI38D72/tYAl
IdIYQHuk9OVCatcGpf5nVicIkP+H1xisJ6XBSIDeufhc2zcmu3zf6gUFqIbDtzfE
nh/kD3Bk22PCMlK7D6ylzFFMGU61x9KNLwVVQEbKYWClIu3eu0LqUin7/pFR2pev
LlaI0SDlLKfSQ9/k5gUpuAHWr39HN80H7rdsUfVDvDWGltZY73KE4AZzOoWeWasT
zg2r4wqswp9S9+kghDg0V2rbtxRovDvvUsN5C3h19ISjYWsZ9HV3pzKaxLScxlbt
Ev747an5mAtmD4RHBHugEwb8R8lrkVnvsbeff8crStcXzaZ6ohVO/0N8m3g/7ora
EIm5kcegdTGc0FtuwVKZhCAnbB4o84yydw8koQAPvCoDWSC91uN2TOkAiPkOWZt0
Pir1frGqqixFJNinEE+5rOjOR5qJzuqdEow4xJqIBIYhlQat4855zdFMgT9X9j4I
FDEE95VEx1FrZC72jy0o9vxDaRpmNFb8LFkRhWH7VX5iU+pNZjDkl3XL0FX/9G1i
JV9imUZQI02AXyfcoPsr/xw2x/8SwmzprQE23KMSrUPXoKW9houOQck5orMAhvDk
H16XH2S5ckhJUdieUgml+CZyw3C0rciF3dFRe7Pb08CN6vRC16c3QRzPsANkwaOS
xrUrTY3iznS5dEx3jtTT3EjD6cJ9kwlgvMmrZVB2DBlOG8MEZ57UwsZ0hfWmWl+L
i6FLin+AdjqfES6n/4xqriw5Fd9/ew0EMv4AA5DOkUaE+A6MZJs4ElvONesyCG9U
bp/e+qLzYs6gvfxyJ4WaXTEwrv9CSSQAcWfIVO+7h4w/U1A116fQb6t+6vgAGtQx
kwQ06tB7xqAOfSKd6KN7Jjaj6LyVilt04a72eqjDGxNaBgY80mDZmIdijevHPKVn
QLUKzj2n8/0Q1RuhgVDmZHXoMN7hi4C9vqsZUbiPYWeJp8DDvp0nAtM5izOR3NNq
OwXUeepkqNL4Hk2afXh33k4UsnOFIKwU3X9Wu8JsTOxCcAWnZjeBObFb3akeMf9Q
hniyn0UpwTlNq6AOwDqQOhdviX7miLdsk2H+X/WcURp888o+EHSlL/FI/W/xen2M
f1O9OMqD4xqJztwWXwU54Z3nrmnwUhuviSyS6puCjdeNUtoY4HN5eLeBampzvapR
v1AFCZtxjpSOhDe+7AG1QQwqWrFL2+Remp3Yeh+Y3WwW91+yuxVU0PY3erpXGgcQ
RrNLbPU/qD3lwbkAS5AnvxxRnqTAA2Z/XEACQ0MCEfuRb7Ew16sUaJCXXBClq4Js
31d6rpS8e4ZGUOhiQ635vm7jA/5V1MlqnDL6qM1UR14zfLZyZxBRDpX7kSS0jAlR
HfF0jd3L9baVBInlH1+J5KsUBdbzhkR+xOLSNNDjRoR5Shb71KFVx4iy1ykZVY/+
JyQxEe7u8WYOwOjC7SJV507ccedvpCzPebU279QboSR1FaA7RiqsoCJKHAFKNfpu
b4bOZvrjaLGaJQaftrWUprj2vNq47BMTedtFfod3kj2i9Dc0diHjgGnNhlaGtM85
/pEZF7WUI5FnHruKQkWX6HhT4HPzv3Fy9z+fL/ig5On6clAa6HWeAVrewVuGGOaY
kdendnZ46jD/OqCQktutsPXUuu4IGMHW7iTJBigu9tYMve2hKk/ArOiqAVkeBRvw
eso7YzH3PAQyn0zWK6+owpZoOAbOK5XMRVhBp1cau8B5tzIRn1h/RLC5qHqyqpGA
QQW8pVZot1hTQ6lo7hemyEiD30fD2zTQNB+NyVhHYIX4Kil3J9Y2fwIbNeQpPxiC
3iy5PgEd6OrfadVcNC9myUE8yMoYaeWw2w+7BptG8WnI5maSffxN2zVJD9FSQRf7
36dJhPXN18Ds0oFO21tKQU1tXof4bGJNmnTIOMDdgaVzDffrnaLR1/YmR59/qZnc
c64lzkaHA6hyWh4TkNSPp3q6X6rsdaEu8GWQVufpHb0sfWCPTbDny5+xWxzqrXnW
QJjzHXiBXiL1t3ICFQzsTs8IIkFiq9Ud0/LH2cl36gmX5DvhWjgy12Qm8BZrUAjC
WWFky94/lNmoc7dDluFRBqVOO1KrGIl9rOAEzHda2i6/5QD78l6i3bjlOARMWONT
Zt6yBHDResAhr/hhtsK8V4o5TEg6QSJMaNm4Zv8B0DEgoGa6FWec6hbspyJYZOmo
17abqYQCwhfRI+zV6yQzs8NCLVEwaR1BsO4UhO7CppjidbviM9ftTGSXgEcME8/n
mw69yfaM5Z4W83XAeLKJZyIBRiorLU2YBuEvljzjyWhfrnoETI8kZh/g+UoG2tz1
oo/6ARMcDnZ68zvAOPP2/kU7NSo9sw2JSD/yr8y3MFzUKZC2AQMSzu6EHVAUkF1h
9lwIoOM/W7B1AdaSdFMAAvUpiLT8/Q2slHcBrnuB8sboDEoa2v1izos0JK+j5pLj
p8sBRdpuZnMtcniMIXdcYJA285wnNj7KM5ySQGPWlBWoOZJirdxqjx5HgApM7O1W
h6TZACe9cl2W0ssca5F/SN3VOf0kICVxjQLRrnDqSj/SCXUsGJWpvSomXvnJcyT2
uqrIB5NTv1TFQIN0XhOpAcMf9OOjL2oHxE596TZ5PlZSxg6rcEIlyqtu4owWfcI6
5wMWdJp3C1djy6TyvSJskdsr2iQdPoa4tPM/ZVZvwHr30XhEvtevtHWVbkM1GtkC
mzd0dT9zJblGehEaYRRqqynSIztRyaTEPaVM4qvEvmLmpnRmJDCmoupQCay09raV
mhXKmKjuEf8O6tVL93a7FgzX8kQBNUk0zBRGORWdJgHomfC/8YGwmm2Wmc/snh/J
C8TRrKpUeRo38HPxLc47pafTRC/pvy5OvBlIIMVKhoJazRSqEsnUlauM8hqqSgGc
NA2pQYfzYDv98v6U6mNIgo0V10w7STgAclkrEGHjP7GSLotZTCtDOI6dH+sWuhMz
gCn+aCuhbI+daFrpNwkHQuFD7fkk9CLn649Va7/3jvnBsFKsXzzn102NQhhkOifZ
IsG1bh9IhxFk0EzxD9mOE+h/kRgr1jy2m6GJq7TeFd4zIYPRiveb+QYtxJvdlWzW
0aFWGP8el30YhfpYuo4Q77Y1kf/ncP/hp9KVQHtUXSt1Wkv/6zVUeAp5lliAbuw9
STnDS3b6qWtScOw6MD9KdzqPoKVrkA6UZaNB65ZdAyFXXX14S+Ni0oH++RJ7cTOA
Lagiq2qtKgyOj/vlkI9Iz/OVgCMnIANNkJrsLHPYIDqivIZFHjEL50X1ujx8rGpn
9YydAEUyg5P8JPRvrdZb3uC3idNl9anpelgwh9JEzksWDeSEECVPhEMTW2+MAfwE
h7KkDod+JL0jPZEtFccLmaj3IJGe7pWYJ8mK+/5gwACiuBIo0/IIlpMFM5LCiB7X
/g/wHXiBO5Vu0TstO5St/9vqVaC1ODTlVE6cxJdOU9AEfcJNx8eGp1OLngZiBJkl
LGExLrh9cWm0em4M9Sfiv1wl2wdeSDnoUFX2DYfAsgLepdzdgxcSP0tSQJSBxK/2
EvFq9bmjFfo696E19W+M/MbEwPNhgKUBK98hvS48E7oMnrME/ISgIpME73/Wk9sa
CH73lKpWsCcKs+IaeTv5xYPV3m40wC6xD5G3dM5VN4+DG4ukZ0+9JJbg5wyabYYx
8t82VO/v3H5D2vbsO/L0m5v6vAZEc+mk8ZDmhkrHYVlhzZMxOw5UfzsBZFeWGdN2
44Z0eA0XJXkvH4+1mvTW7a4TyOogQrqZQ5gUVSgVbXqim2UKtQnkx8WlzZ3u3g3l
RMJDT2zjc6EOATCoxS9rQVwhmN5ivHb591Pa6i4Z+4Ct5WlSssRDYypPRR3VqRtx
sf4CjPiHVMGbR/lVeq/8Fme5FIn9MaC2twHrTzw/zM4ETAMQzA5QHXG8jV7HOTWs
QdOQFQjR+YBnURkDe71OaCZgvDY0fjjSi9TIfgftIKaEiTsXXHBdko4Ed3Q0xRW1
cLBIxBt7+tj4iMSYhPNZWYRV1WqLKfNQ612nXRF0tqnWfIcUqSpWjjYj+5FMtitH
6QfBZw2ROLuqfbhFtbd7sXXZ+YEQKMmb7xVoyyWtfz/+VXf9sKLOJysGnEALtzvf
8vyEctrvuI1Bk7vgdr1u3bUX4kkn+S7qvlUSCttudVq/CMahn1nBrKu3VhoCPCYq
clTx5jow/efCAJcfPoem5+s4q2qiGFg/z7y+3rVHiW8l28hEdDsI699pvGckQ/9i
fBeD/8QSpSS0Ge2uLtMsWQPm1gcH+avrmDFnoIzJokdaxvir698cDXIbf3DbviV6
twdbX5ffTxlsCn4GSQGkK5lPl6GbnfdId//l+xeBig7YHOO9TpbKhPV7QDn7zNQM
vk/psybkbGUtq5jZYBxveOx6k1J8teGBj4k5pi71F7fViAiNh3X9YCIJS+ikuLPU
Fflw2l1f0Ib/ohjTdMzTiHOKygYxXyFHtN6jMj7FITnb6xstoRehmp74SNDAPgQH
4CdF7H+sKqN+xemlBNT/KQQRf9Kx12I3o4tEQWvZjMakhvXxZcxJRuibkDV81IZR
hgxDNmloQjq6LUX/i1P8VXBwOQSD1wP+yDjYRqiGXM6kjvTfWCcuvHDt7anU7leC
VjOyYE2YEP+GedhbH9fT1k3mT2sJDWFx0Nfc5WCTKswwnJnV63K6/T5vCS1pOwWl
H3J6UT14zPU+GFWThb4j7XAFOg363tkMU09L6rnyOCxWWcSezb5NP8DOI/eU/h5v
VGdDV1OS+Dtu31TEFAQEXtZ9+28m8G5Uclqq0WcLyXbTioQmsceE2dXG26wtRglT
4s5pSpwGtV/p6ryEp+BJ5WfSdvYG9n7ZMjwhgKeKRwlxd/FdAFpF0GR78HrqV7Aj
0/n5yqMLzerVKDoFoLgrSVzMSVmFJabGF4LPGrL5hX4uKBYzboUDGMsqvRFL5PQU
bA7SlhAzbRpzdu1NeiCjV1s1rIK/qWQzsqHqxOVvLcZABXqbeQTMkDRQ/Z51xIDp
RFS2lExsqas56WUPAckzLIHUybrUA/Pqzl9Ogooycdvp2cbkchlZPHvv0jBk8eoV
tZh5qjs7UOL13+9w7nbnTmI1WF41zK/o8qZcAfnWFh3gQEgSnPhpKiQAYq9FqO2O
nb+AEX3J3hognfsur0n83aIo/GXEdsrEgcZnj5txEiMDwJDMJoc+IWv+5WnYyySw
wl4MI/w3fCNUomVOak0WJgZiTgf32hZssMTCeEuzYakQk3GcRZpQqEoKgSegRAtz
tKZ7Vrc4YL/8NAawYtkiODWNWgC6DOG6lB8nNHxVIxedXlgLqvvz2K3ijxBNFuti
yyWj1zrQv95GaJr6yLeJzq4l/xSHMECO8jMImSsgjkSaoj6tHGBCg8b7w8IJ3bZW
jJqYUx5ru0u3GfS4wcriynPH5cZJiESeEgvm59fIiI9lhP+rgLPZ7WAUeHJ0lnEV
+qzYWPM/C+8LtWaAotufv0znaBb0Nx0iccl0Afr948MTgz+JpYHuStmsYEIAcawJ
iPmCwzRXrWjFGLI49z5o25zQp4/2KrHyoJmMcaTzDxRHqwJAQ56SXagTf6Qmj1uO
FRwRHajyF29yjTCM37VJ7JIgLCAV+ZpLgo3xeI2A6BLDSa99unqH8U99K7McVJ7W
GqUZ2QAzXeOgXILD5Kn53xJ4g7oWcB5V4jST8smzktUjyTqQf91N1YQsyWsW06cF
sEB4NeymNpsq4gGdSly4v/mWIVugo1ryL1FH7mk+sYbGr6vqdTb7symAEbJsB6YC
GMkp0B1hvCsoJB9fazO99As0tA5d8y3AozPp1YPhRRUCwLYCF6SPVPKcPAnc8jW2
zR4HCSJbrwRRbJlyz4p2lwfl1GH86TdUo017Tqf+ESlJ8eWw2fDe+sfLi73JUcXO
aPxdrncnGo6GCpp0jxE7nHL1OfO+yyFZPGYCWHByHa4m48hP3gzxhvpHBrOkWRIi
p3fGFOLQ71Jg8kEK0Kvmf5bcpXWOkU22C8uCbX7OOSYxXZTQAiwW/N0jLJHUTGRR
8N1oj+OTAgHwwQ4M8v0AQ7+vOS2oG/rzfPFUvMfrBBLCEj+bgWtKVMPlErXL1lZZ
FNbA8I5rHJw1fukM33GLQ0PKM2GS4XIDzcDYDCSTiDN72h7TPSXUUPE0nUn/2RNY
/YwNdbnm9/utj8FdEZGpJj+6vLpuBECkNNvsIUHYa/E8LOMqtlnvh82gDUDmAnSE
FZs0bBzsj6BvRMY/qnCMb5OPeepWcmJzp7EXgFW/rGwY8abnkRdtmqFRg7Df/ROe
9rg+queX5IKcbImj3AUO1Q5Y/ZzhJoIES017nZEUkm1/uTXMP/DpcIs69BJh8+bl
ApUtZjjfOa5RW7wVfGiFS8NZbc3oa2YG9V8wkJs7j83zLpIN47KQVtMX9dqiReaL
RYmYIXJVWdCsXPibjKcLRgGc84Sy2obI0OokDjvk9wPzMEPfiM+biajAeit2Olip
PsQiULEhA1XThDpN6VqC5njcI3B36opxYQnN3PeGTjKpX1d1FPRi3mwYG1IMnTZZ
rpFV0w0/dahBvCR+Ht45Z/bR0U1wJe2ElLTIAeouLck5uD5dlu843fjEYQXsHS9p
kOXnza64KTSCeoZdlYNWVU75Xgh+zZkdoKfGLCYcQHIfEk6HCV8660r5rQHAEDov
7FCG8J3hO6pw48NIFl6UDyK2hNeMOshHYo4mqIJqbftkqqa+tY04yXRXHHUhVfhc
3tmfTj7RtEyKHBI98rRV/bpY6JtA4MboDcGJ0VCKi02yRrEcq7s/h+QKVaFhxVSd
5PqPVM2qU8KwR3vJHkbMEXwDYJGyqFAXOqndPz9hOyAudXeGctqzIsX04ud4IAHU
/f7THkErtfdD9oBy6KT189OTyN5HgLBFaoBrncLYsk0BBpchWF0NDo/sorih8Mbn
WwkNpgclvYyj2K3V6pi37LKihKx5h1WwAiISndFn3mAj/ZADjJBlSUJFWIupTdqX
36Khmrgdk5Wj2XTkQJBbAZgFGFVST4EZuY8c+wzIkfIbGaFJGZjWSq5DvDrhov9u
ohgn1I6MAootPchbJ/xiRVIgoflrmmcTGPvTDeKBtDmaYTHn4SMEDXk/T5k9tIgq
9uiC6+NTePysZxqjDumsdoRqYoWmVbfXmJOLmonI23fU+tvsWNILSRwsDH6FHriq
THvGSzQutevrHUpbNh4RO/QdZK8kGKLi+WaT/DQY0boKyhXCHAuy1IzXjWeT+J/t
er67RZMZ0QNAlaixrUn2FR7VJwp5c/S8GFmNpPHQa8+7AOxq/7FMJpMVhu01rRMY
RmczxvwEXcPTbblxuvFDv/BWQeRb4BXIKXeiQGYsbFjbm8rZlRSpnzs4n4fzNA9g
QVzyxnrR4QCHIGpndh5Awnfh1nuRdbEoSRthlnmsjVf24L46Q8I6vYPRaphUJElM
OY3g/dOwoppP5jM1U2UU6MFGjCs/Fi6nL66ENixKJL5PgkwS5Fu98WFlQfIZoNiE
HvMwzewm/ToeTiOdtXtsADvI3ekS1AwGj0BKlby3YTwKBgF2VALCNgCHrdyQ6hR9
K9h2mBPYaYTxgt6WiCkd21xCG4hVdEH1S7FPKjHRAsMgfO6MQn2FRwCtoLtKWsG3
VEDdTMwXCF3U6VpXC9olWzJdloknPS+vokAq7V4ICYpDKld46fb2LaMJ03tSfTHG
ShCRMMy05igjFINXvYCeQXunRSV/L/2Uk0WdR2TIt7kJDV+AHLXy1MkHzhGkc7iP
lDmF1JT/UN6bJfj/WW4b99pKbQd8h/lbkY7q2kXQKizEDmTOrFgqmLedjF/c+gDO
N3b4oAUVhx+w6NXDu+SeMwFhjix47V8HN8a/CoHG58IxEbQcWacH21bAw11+SyW7
GzlRKXZubT1ENzpCtkKrdTpiHTfYlkNCZSdLEagYRUvlUFM5H/QRJ7xbo9EbdWd6
FBV27kwBrlmJm8oOkD9OHTJ8rDZu/hV1gx1IZqybgznV3u2FOdonRwhoUXPrhHDS
gSi5oYZ2d7JKWNL5wX+u1CT0UZh7D6Y0TamZMLzc9+mckJC7CoKV/emmpbuiKz2L
sfTLXZ5oV0TJgNTyNOUaZ0lU96uaKP6h2Q+hjMJ1aQ69dUAc5ASHCC3hpp3Njgrz
A09/DaWL/HGDkh2iTFSuD19TYpFfLkMjTA+6hK8t96njWDHWmsAEOO1SuUxVxxbF
QUtbe+rlUMSz2LFoMlaPLE2uH7p64qlAnXAYqRp5bMMaB2obfnv5+bsUC+eu+Fwv
BW+B/bqtzUZPfF8UjwDGXqc/OWWiosqGXO68rzg3+Wfmw16GEaYEbyI6y0EGJt+b
xnJ1KZA9XVAV43A31hkvLiY0nkBcyZy508DZwVQkkA/c7xMvBwvVtQ6wARPgmL+9
GPzDk5j0vQjavrM3kNma2m6SNUh5wKLsEACTKMRoriHiQQIsBdbfpo7BZvn1hUhy
Nkh2ESssK3iHcuBhiTYbBUHPN8ea7ycvhLg7OzpybhM5gDCCj1haBLbU8ZhBXmId
jJeUnWbQg2dfkUvzBO4TqJ4JNfuyK8sATVg9hnKygGvg93VnRDm55EVfvYEVObVt
paH8COPxJYPKXROQ9bmfhOd5LdRhj1ZHHxd3vfB0ldPDfjer61KoBeUGwSRvchpP
jq+Tt8lKsN2xCQuLT9Qi+T7az102cFskkVm1vtGzxEuaVA6L6BSI2uER68wmQE32
OuKt0jDu0KWr6ule/bQV2QhhKA5DfeCPn5AMApayYXc6s/JBs3XZZMpw0ZJsPgw7
plnOJfX+C/htj4HgPU3kMLbC78JiTRL9OeVs2yPrIz6TqtQQaMW1Uwc0I/GC9R1h
Ppcx5DgQp82qTbIUo4CzLwO8+zpvkcGMRhz4leiQZ29AEe00ub7EmUY5yJq4dl6U
c4RVptBIpXzSJ4F/CRqs/SZhM7ziVpa/dG0d+WZWEQ/qvPMbrwy6l5ElS5lyjxBv
LLlTbdUOAsjxt8UBY0E3QLtdDL3I+O4803WnMFsJx63f6FMOUq3qzTqMWpJ+QRlx
k0p4+j52k6o0PfAFcXarMItIkaOAtdwDtTad1O5/rD2HTKKwMHbGxepRIC82G70l
Vq5WVI+Sd2MCvsSNOLHqNx8XkJzAQT3GkP71McM/hghaXpF/nIRIiQVWoxlgWdQW
iKeBCfI7bCD1h2e9TkhwoM+xzcaz7v7j/vBQ/EautP+KgHIWWF0TFyxUU1IEQmQW
0UWsaEaNsXgRODciDy5kK0NIb4zcK5XV/IB+zP+0DD2uAroXKfdwuRspHdf/3Q1L
hMdgSNNweqS5LB2g+JXc2kl439+UxiazUsm81fK777SXRKXYMXD0vwTQZCv/p/rI
armBYxcVxAZF5i9sYR3EkT7uFOlFYQqUKHhoRBjoHt4GZYQP5pHBFDMkQZfO+zv9
p9xN1G729j4pz0Eh0JhyZIWXpSHnD5THLqLq/67K52YRma4FYhIXY1xnNdEy+t26
p9CSwHRjmAAFnDHYanzT35Y2FBhY8HieGVTjeXJUYADdw2WNUNFNN62qRjbK7jNy
TCVvuO4ebHpdp8GxoBe2spgpjAtdKIzP54ooZaRz9hHFFZ9VHjJ+o7JStwgL3mUw
8XVnI6DkUYgUGiF6XlEjv7KOQ/QNTZH8WFT/SDvLO8Y5R51uXbZooOFImdSPLBsA
mM1N61u96hWE/Ic7YC/2/u8mwS1U4G8ApLvCDDaTz4z+6e86zHLjx0EmeO6KYEo2
LtbAF3asn2e5R038T//qEWtSc26r4/ePJthCwVX1OiNA0k+wwXExr4gDJ5Wj+giE
RYNflvCRaGUbzlV0uEip53YmUkbK5ToWvxowQI5nOwwS3VczXlI8CIaOv2wAG/Ec
fGWSkTLU/hP3nKgnF3LPVm3p2G1JwfdV4EiawA3krVh8xCwzIy3eAKGtHa+Kgfet
w9MdzPCRLLQ0VhWpGct0sxS6j4xamEeZez6CRGK9/MBwTyy+R5QcZe2u8ldMF9iB
03BblpCQpht/umlnYBWjHiDyyTyHEOlfbO+HCHxCPW4ffEdGm57dvhfO6R30benK
Jz0WpAM6w/y7xACdy/m6XHUB/wcQiVd26QxNdd5IQRgyJtn38XGOF81XgwH4owD7
CKiy6BaBtDjpmtd3xSCIbqesQlteGz7xjzkNMX6pCpLGYUuF/p9yP5zbXIOztV6t
rD/5p2WqkNUPnqODXxzdPRNfAn1kh3MDXDEOdw+9sn2OGiOmTr+VucDQ1IoRBguO
KyK/D7LXpMzbkWRNf0IU20h6TVadBPUuSb3jjpl4sRUtZwBl1l4b6hUnIwWFq7Sr
pcNFYF57xK1GvS2UzT1OiPsdTkqC/ISYKSBsylB6uoShhVHtEAhp29s1Y4Mf6MGc
Acvf83qNJNH7FBd+buzQtkpw4C5Fy+aTqAH9zZvWQFuLHd66Z/amIlSAQUXwb9ua
k3p7NK9CPzTnblyxLLZcgkoIYt6gbvLSvNOhyojEniu8pWt5APvThQ5fxmoIAtK1
C8zDfwyb8kh0MZbYvBrebSKyJUSA/iOGHeZx1dWSSTJY/A2Dl6nIGaW8XAC5amLn
tKT7kDy6UcU95WRd7VuM2Op7I6Iv8PKoFVAeArUMPtZqZLaZrFohrSBh+2s2P/2q
xqEinSb9xe1LLJmW/D5cEIa1O/ZxbUgbaFU9RdqUVLVI0RmQFi9ex4pGG/XDFxo0
JW+myJfk/BfJz9EMhYI3KxlPWSsWqM1YS5zMMt9OIxNXGSwPv2pxanMIDyU3dNUz
2L+r25hEOwlvlmQ1PSO1x8Hz2tV4zc+6ZMnklr+OpnCUxqcJk/S+FOmKC4d6Io73
aQnf0jM7kR+10uoSD+1Uv/AuGIwijsuxIV3o/I87DDSQs7M2/j04faDvHe8CNGfc
5QqOJ8YiMTMCwurZ6Wnp3YrOW2swx78rFie9yTposQzTaXN68m5o5otDZKwPYIJR
iLQhL0WSLLrolXev8N7auxu+TNE7aeuDh0kZY5NRvsi6ib0XPUxoCkLsOnC+i4GJ
DFv1T7diOrsP82Fykxf4f9M+a6DqjLeK3J4Nu2VQvLeguQIIXOlAzZo35odvXtgN
aPD4dWdJIX/o62QRaF6IipIG/qT5H38/ch5i2GpLKmwpd/dBjOpnL/qt1vHopGfv
oBgDGZWontbmfJLzr3AqQ4GuF9jDOrlHEb3vcbgVC2y4UO74aR1bSHjveB3grJWG
FHAKJll+/Tr578bxC1mJ/qsj3niuoIOAQqW1VV8DqWzuryp29dVayKlBc7bc/1B0
XNW86Hv55Prae+AO2vSKgmIgD/ZhnW12B3TNb4Wr1AAzQPrpr5ahMlf2PryDJzup
cHGrTXxQf2K1vKYTT3VjFZJxUkTNmfswDA6c0vb8QdeH2EFB14iQkEy1TlMWOYu2
hYZMWZYm3obvzafNDXNcLwW5o3KUDe1PD8kE6IFq+jNJZQOHo6KxiGoN6c0t8w6Z
CofoQXedtkFTiAAkpg8w79Sw0lmxPSP6HHQxD3xrjbw4Vp1eLZ1FGliQQicebL5d
6+y8NXIONOc2B/pd8HxaSh1SHHEB4Udmc29+RdY8V2jI3ssjIVjvf7Uatl9KFg07
v4wYTBwtZawrieN2pTVKtQBQk7uH/AXBwfhHcGbrZC6ddKqR9tb3RSI6DPC2DhkB
ljty7PJ3JyaFSTlzH5vMGwF5/FH6RWT4BrRvnSGvChX4SGiLiyp+0RQ6ZMhMeg4L
ecftiwvXVQ6M5XKtYjRFjKi3Xh/fQEnkUZxZCVmuL65TEisfoGmcjOHGCwcT6q6C
oKBJiGp3nKbF0CHdrJ8UxJjh07/pbGKqBibciUxz7O4/HGXy7KzLDfBBB8HtTAZI
GSAflYsYGOkzWxAoMD1nt19AD8fgtR1jEBf/TRYJ90SFpo7eukcN3hbfqHSFMaDS
3/iUD5R8mnuA/wcwQ3tcvjGL/gf6+3vZoE9LL/CO5ZGNj+JDzn5VJ6/KouwHQdYA
wpW37HWT6CN7/f0KhzklEqCPdMSms6gTXREJQ1Omsw+Sn1ogHRGUM5nr+U+hv3Y9
/7QmBgECjV5ZBtMSItlsxgyD7KKAOZpO2HRI4hKv4TSFOETs73zP0SiCXjo/WVVi
AUrU6Pv+TCgQm2C96l1XAs2GhfKwB3SMnopSBkmV5dhJIQRmCjvipXLptyTxR8Uu
CoCrZV7eTJD1/3pNpp7YXjOzu31sXbX9aYKYoVA1p6xM+WMshO9g9MCvXmuivo3O
OyDTtGTf0ZikpxNfEXpaq+gfDI/ZwbYT7SZT4VNhQQRXt6JaVnz9WByLskCVlSH6
y52WJJZpkjH4Ek8pajVsj+pyjfdV8ZR6QLBaDRY/SlbqpOSgsaDejIAIQ75GpHHW
9W/QSzV9L4uhgvvNq19R5M8k+ymjr6FS8b5Nmk14kaQC8F5QHvQ0ErYKWsMS7stS
LhjOKq2SwRaQ3JbVDgZt3QZmpRu+lPQIzhXQcJsJxapzt/7BDAaxp8Kyf+su1IrK
G8EVgZUmoqIRnL/IV+QsBf5ppEMf5QsHXIZttsOLZLpYfkMBTSZ61fboKYkvmINs
kBH6BEMMG+tbM1FcMf/X25WEZAtvKe87lcOpZhDAD0+3jWTZOC3pPtgymYvOQ/4R
gLdxEQogGo7JyJS6787kfyUN0Iy7x/FILlqsMtFA7OURD67+EWdEnHuGhkYri3M4
ip5dQUz0CH1kEOoLjMfniBF62HIP09ouZWreWzQnkHTq1yeESIbyESCE1qlzLQ6M
6Ps/AWj7Lpyk/thfREt4fy4gdMXBt7qbuV9azCKofoNQNyslcEF2VbrxEGONBgAU
PqqoKWw+h8ioP5ORPEMmD6w8EzCnUonn7fZCqaiyPP6aQcifBq46oWj+SKzy+I/J
XtodgWxd6/MaeFvihj23WoukJlFKxoI3R/Uui1O5Mw6kp6vyl/EUtVc/Qq4wVvbf
OArpOT06Ur5kUjF/ZS4GeT0fKUOO2CRkkIrRNqmLNcEHzFf+95/imOIdAhXj38Fj
82OQZAyrjF4YaGMPP74bmdcaupXUwsQzEfS4IY+7n9h9jvkqX7UyOhstARvjriRO
Hy+yLiR6obrxUzRJTe2wxqOVCgXIbQDFWrGeERhwzqL9OLOyDSPOeItrngf5V5UB
BQabMYcY3kPXjqsR69SgB2qhU0Lm3K6kK8Xe5ziNjJBV5zWrBCRQhxKekbcLPY6X
osa6qFePHJT36uT5mG8Ud50UDYqzVjj2J5P3QlFn/XOkK/n7ZVPpInCPkKZGua6N
b1UmGls9akbt9Boc4+6RccNWZNW+nrooIaVW6bDVxUYQKrHXrkRw/QEazY0CtexK
JUWuL5VziQ+kI5n3rCjcm+AasK4cFryLVPjaXnDbs98=
`pragma protect end_protected
