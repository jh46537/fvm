��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_B6Wi�KBKg`C�@	CVfg%��&<jx���P`W��M)��(��:�ִ�7�l2�S�,*J�#���E%��G�?���j�3������������6$K��\�bZM�o�n���9�g���ظi�O~)Q}<Ȯ��e�зK��`6�:�k��V�]+�暄�1P��SIm<�$�>�d�I<��)T�ҕu��<�o�&������!#�Mv�CLI���GE\,��;�b/Mw$���VS#�����+�-���k�����m���%TsG p�]'z�SF�f��v�3�.�����k����6�:�!�T�e�E(���UAx�����J�:�*�%3�(��э�?��+�ɐ�z`9I~<q��A23��OIa?P�˄\�;�ݮX�[���Eh���j�~�jн�7���_�P���iE�࣯�F����*��.�֕z@s>8��=�<��� ���!�{�K6`{�t��~=x�g���G�����q�/�ώ�S+�X*v;�����wר���}��C���LZp7"S��х��0�T`f���?f�ỼÝ�c&�Wb�;�N5\tΧ��%ܺ5��|a�+���6Z+�f�,�)�G�98��"���,?�i��N������z��)���w���r��BزY=�]��Pp��1C!�S��'B6������?�?�t�pL�ݱ�X�"���@˂Gv%`K��"�|���FN�8��e��[G{��.P��ɰ�n�OW��붪������9)'�}_�dqر�Xn�<�a����dCE�F�o]7ٜ ʱ@\�����Xdʐf���Mb �gCg/G�c����<{�Ps����G���!��G�o����l(��fʀf���U���ڠ���z���W���f	�a�9���A舘<(f�B�~om�6�Fi�ؓdf�FI�
�/=�qE����o�	v�Py/��ʾ����Ȥ��V~�	¶d!�b��:��xk������G��iD��p��]b܎�u^*�
���?�A4
�+�H�皠��|x
-�l�I�(���m��hD'z(2��fv�H�ţ8k\�5#�~����.d�I��[%��W�(�t�a	[vB�vd��ea�G����\9v��V�w`�.s(4D�kPȹɓ3�z]FF���XC+{xCy��i� ����/��sk�4�u��@*_�%6Ȗ(����ꋻ��f� X�x��v	*�3=?����6�]-J�����;j,���N1�"Іh��s7n��]��;�b;F����҆e�ϡr����a+�%�Wo�O.J��o�2�roR5ʬܖ=���3؋D%^��i�[��R"8���z�~����@xw��6q��M���R�����<�4�%��J���2E7�#�Y�� ���:7��IJ�c��)(o�5a�Y��#���9�i޿FO�����~F�-I�@
"�=��2;ݻUT�{��hkz��6�l�Ϛ������^r��&�d �C�5#8%�۩�2>)��d$�]F�x�i�M2�$狷��U�J�7�2��y�0Y�����]�����a��X���<1��u�7P���!��#w5��
�@T�u���h��+�ӻb�����Z�W���l�K��cJe�N-5ļ�}�-����ߕf�w�e=+L5gM��S!&Q�u7��֩�9�� 88�����fP�zW	Ě��|�G3懅��'�|���T�fQM��d��@��0�?�� |2�:�k��ȥ硈+y��BC���Ai��g��NU���13�^�Fw���F��"��j�k�g��2���|�ʊ��`{�.Be�U���v�r�#�p|+�S60�E�c��xe[��Hr,"ki���:ş:��F��U[Ye����?s}�*sWH�w�;hf�'�,��z���q��ɇ�:2mc�*����eM5����0��ZG������5���6�⺜��GŅ������s�N�`����?���6#�bd���d�x>tHg~7+[`�>��#LL�!q�M��EB$�޾βyx�rd�Nx6w���q�%�Ї�l\9�nA,�|�m�����h����U:�Pm�
Dh�<��\;�0�(:�^	��9�& ���g6�a����J���=)$P�U�fD�!sCʺ���8��І�������B8r��m�!�n}Fqw����*˞n���78O~S��Yo�IQ�$�Qe�.�U���P�����A��ɪ{�RH��l�c��:/��h����K�b����n@�e�㓭�7��b�/2�g3'ȸ��B�F,���u:/���>�S �B�������u�/o~�(��{80n�r�g�_���l.!;>39bs"x���6	��
�.�n�������~�*��;�|v� $�>�ϺД:+�'��!@#��=�WbF��t������,9C�߳�̻�9�ƾ��%Q�v���Ez�|55��n�Ykg��$~'8r�.�ޞ�`�>�x�[I�đ�r:ڞ�?�G�>�Vօ�d�ٷHķ����+�@��i\k0h�� ^���&̷X}I,H��ԐV��U)����f��O�t}R����k�b��E��#i���W���[��%<-B\�j���10
h,貁y"QT�͗WיGS���rZGT��)=�G���I��h�P�-���<�5{��Z-��;�.��aez�a��:	�1�U_�Ju	l�DLKg,o]���y[�?_���msO��,R2v(4��T�}ќQ������'���Ԧ��U~6;�J̛��C#�,���ظ8~~�_\ԕ��7U�,�:b� �Y�/�wDNu�>�\�ce2�9���d�J��,����3�*�i|�]�P"�ǘw	,��Ƹ��Hҵl�f7Kp����Y�#�����!��w�e����U��x�J��s쨛f��o��
'���4d�P���V!��zƶ�O	
)y��?��CY04��3tW-ڸ�l�Q��r�, ���A~��y�|���0?�0�_�(�A�~=���d����ISÁ�xl�L���p�5.L�
�����S��m�һ���X�7�bZ�v�F�|q~�<�p�E�[�/��rLz��l�������?h5ݔh��O�NU`����G 6�[s1���>5`�V�h����Ľ*(ٴ�%BR�Y�$��n��\� ٹ�,>A�-��
�z�TZa8��yL��얪'�J�S�Y_�Z�͊U[[$��3=�jw�vO�7�!B�3B���LyS�P�{8+��ש��''���
��M��5	�Ҟ&`�f;�I�F(��D:����,5`�!*_@e!�ʤ�����`TW�~]���7����b�Uԧӈ�Z�	�MD�"t>��v�^
��r�]�hKT'��MJX�Ɏ3t��ojG�-��G�������N�
��{W�[���b)�4Ri�.�H���� х�Bq�y���\R#%Vy7-��BS�H��-��b���?��a7��^�����"�F0��\�����Q��*����.	;(r�P�f�^/s���(�W�P��&:,ˀ�Z�ʉ�69���ߜ�@����ŉ~H&���"�*yP�["�?�F3B���;�X����uGHc�JT���G?s�dހ�)��L���׊L���$�P����Z�IN���J�0�Zi��)Yd�;��wI[@V�x4�bŲ7�����[�o�����.�f* �$uR߲���Q/��.�Yw�&%s���(2Y��V�Ӽ�`#��6��6��X�����d,��ȴ!��R��c���d�=똩�`�H��q���X���9@��j�����?�������J�����Y��o�N����j�\�4�X(���"
Cק1��"�D�ߔ�� ����\��^r�fOKRԴ��'��9�z� H5�z�j7&m�aꚺ���(��3h����ǥ�W0�rY-��"��Q4��)o�?sgP�u���O�n�#9���2p��笘�/#7像�o�ER�?�+W��۟����9�˹
�٭�ql�׈` ,:��L��!�6��Y��v�$̞�Y���R�8��`.7L8ƃ	]Js��Lns��I���ntz�������u2a$I��`��Pui����!�v+�~�2���`�����Ԋcx�D�ѕ"�Nh���|.������8��V�	<] l�Ӓ�\D��Q�b��G�|�|�4��Lit��*��{\���W�-7q�مZ7��R�ޝ�	��SȐ|��(��5H�O-|�p͆�1�(��2#=�i��u!��2�d���%��:QG}�
���68y�[󨜑㗴��RSq�6��Pio�ck3#��,|X��O���ȧf_�]��Dd_.����z�j ������8ۢ����_�]N�H�p'�3�w?'���(/C�����`Z���yuɻ��ȁFo�vT%��W���id�|��G�M6ٓ�@eቡ�-5�����q�U�Y ��W�צ<3maN�
��LY��'��~:"_,?�*��_[%�n�����g^S`��߿�&��ov9�U�����q�(�<G�lX��`HHԺrL�@��	�sPP,nVd�c��n�ck[Ɛ��Q�v��}�)�bǑsl�Ы!�n��9�Ȩܶ���m`s�'p�������e#� aX]y�,��x��W�p���M�5�`'�	��>� ��~�^nb�m��NP;J��=�b�q�=���V�̹�
[�H��t��%��ĝD�Y�N����N{�Zt8�2���V�krq׵
Rl�:N���p,��8Ο�.��b�*=���R�߱!Ao0Lg[�a(��Yr��z�x�6���Ul�j���*��A^G��4�>|�qyO����$��Yj�L�k��p���Rr��|��?�UW��'Ri��t�&����2:v�Oh�D"w���D���u"�`����u�� .*���Ǆ�z��ID�B!�j��>�;ox���0��hzQ�Kꚴ�d_eF��z��UgoS��8�u�v��O�^}v9
�.{6�K�n,̆K SX��m��ZY�eH�2>:ֿX���C��tU�wR��MMU�­����Ͽv�|F�K�QW'FN�0N��
�����"W�����X||��H_�����+(�X�k�7>�Yإ�[N�z�o[i�X�g��U Y�x>������h������*�,�����FY�8���j?\l�����xǚ^6��'B;���@��
u_TW���cF��	]���A�������q�(2�Z|�
؏��f��rK=���.�Lg_�W��d"k�Y>G1͡0�"ǌ ;�Y|>�<�c�����XxN�i�.�	)�������*W��,�v�K�,l?o�|�(_S!�o��/J��z��NaD���"nB�;S�0 ߂�~�VY��Oc�8��+>��/�ܙ�3�5]���9�иi�|��!U
cB��q(;$ٱ��5����d��RN�U�Wtx&O���B��K,/��ߤ"�v�I�nM�a����o�]"�9����%�EhP�|�1�=��i�&���ML)٘���O�d^b���y�����BȌ�L�J_�Y��g�(]��U���/��7�Z\���"5��Z��2�� �
��㣋�9ab4�K�ܯ��7��2�Q�~5[���^���u2��k�fQ��O�d�3ѿ�A��p�T`4	�&g�K��n �(`D����[u�0�sZ���o$��;���%4~�E��9i]O�����n%��$`����G	o1����S-j���&�e�f"��~�Za����૤y�]_�dO��,D��O���3n㪡��Z���?~�ԉ�w��U�B�/ǔc*�a�I��U&���>.(Hc]5�1�b���<������k�vC�O��?X��6��Cx��X	r0r�XȪL�'����b�M��&S�N�w�Y�CU��
,��%��1����\L��A�Bt-�ou����"B��zC�?��3鯉UY�d���D>��>����]m��+��L�ކhF�}�����/���L�eKŇ�������>�LJ����04���o�d��t
��s@���h����������ܠ��x<$nf��ټa���8�%P'�v�+���Š�'����Mܭh������`�_�v꾒��9�1���7���D�[yy�(!E�'��'k��uf�B�9�S��y�'���탤
�GpH�>(��Hσ4�v�u�B��I��|�A/ޛ���͈u�Bu%T��L�џ��%�Ӡ�N�;8�*�Иl�C�%Z+�{z���:hT(�!��M�k��["���鷔���)�\�+�Бƨ��`.�*�U`�`%7fY��oD�{��b��;C�tqs����������L}V߻�9�'(�m;U1�q8,�4� �;�>O��M�X��Yע�ܨ��I/u�GF�-����Mn�N�h45���&}K��U-E;-'����Ac[|���Y���7�Ed& �i�I�d:�I���k
~ȁQ�d�Y�Oϟ1|�����i����K=��56�2�����%K�5�}<Bv��4xD��	5���#Ѓӥ�!_��+��\�Aw���or�!�m�wgm�x���}���~�� a)	v�h��Kq���}x�#0�zW-�)� �0����WB��X��S��R.ԲUc�9Q�#y��v�]���4��ɘ}rT��=�F��_'W$E��̤5Q�Q�_��~�>�	����G2���J6�#(h�g�<g�f��<1޹Y��ZF����r����O�-�Wj�N�~G#��N�q��k���٪ieD��X�~�"�����$�T[��xq�\�G�c%N���q�җX�nq�U���l�F� 5��#�$�k��+�����*[��S=D��9�ϳ>'K�Z�M��&Sx�{r#�l�(����x�k)�7��U:�m���R���w�K!��Sn�t{&H�16�8^�fC��ڳ\��hQ/�{M��pE�%\�)x�qWG���-��=n�Q�'�Q�ky����ɹ�J����("�.Q#�7 ����FJJbr�Py����b0�8=�T�b.��q�CsBu��e �B(1���4�r&��癗�y�d���!�w�ه�_�����U�;�s���i�����k�R���}�$���]씍lF𗽶��+(����~cU&���h�)�`�E�;#��Hȃ^W��"���n%bE�6�l��`ȱg���:�}8�8�ݬ��n�:��6Mfc��W�L�f�Z�� ���U/US���Vcn��v�Ǭ�_/����^~�y�Q�����PX
2�����Aܳ�EЂ��g�'J�J��1�tI������Q����SꬂWI��8>�d�W�x�U�p��X7�gdP�?֫�"q�-��wo�`l�%�+���]�	M� �]�?�ϰ� j��LِgS�8����oD(�>���:��B->k�V�KFfW�xb�����GaW8�C$BZpݟ㝏B�,Kf�ꀅ��Qt%�<�d��]z��r�[濌2%*�������ˢi���U�"l��f��Ey&���S~���ߡE鏚o��(�1�i����[̙6:��Mi��&�M&��'���_�ږ����;��}D"�����ŢIi�{?TK�~x�rP3܄p�1���������BLO%�9�v�G7���% 