��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&-n�7o���U�����w>5
�~]#X`Z<�}�
��[�JzlB���-|�dv����BZ%�`������I�W)���,��0Ģ� &��uTFb���L����a�6X���6"�f���D��Nw�j�k h1OR�|jj0����O���fߖL�n�v��v�1Ef��h�
C���x�g�`bB7`������biTG��o/Ns�|����̄��:A"-��m��D����M�Ǫ�������ղ�Z�0N&^?'_�B|Z�uAu�u}���L�mѮ��L}Lظ>|�e��z�уG|������H�0�>�V��^���:���y0���d�*>��a@!���	�����X�M��L/�\\��
i�+�?2H�����<,�:��&E�~�Q��dn]���6_�ny�R�i��G-(D�T�PAA)�Ew�~��T��\9���H���3n_<����:� ���>�,r�o����_��!�d��{�۫��f�������Oek�R�
���DHc�:�+�ގ;���t5`�h[��Z� �1���I��r�����@n/�ϠY���v�����Yt�x�����Abv���Q	3��k����3���i9R)+On�Oo]�H��`��_KW���.d�*M�x�o�_�t$ �����yG|sF_���q	I~�$%��5��x�'�I'��x2o,P�brMz6�.��ΒS�ǜY�C�W =�3�X�b���|~��UϬ��,��td��C.���z�����AL�v�W[���m���
�cL����:Y�Ҳ�}�|Z�CP�\S�HyI�Y����ǈ�I�tA���s�#�:[���E�=�f�.8:~����������la}�<�`.%������W��;�pSj��܀_�o��=�������Σ�6��bY�*E�'���1����E�C�%�N�6��p�F�a"�\H	��.��{6z~�Q����1��?_���w�!�Cw�J���f�������(��8���8�h!���6og3�}������	����ܶ�Z�E��$
u�����L�
�=��vj6�6�.{�����(�F�]s���i�Ưk&;pn��4�������`�u�9**�5Pq�`s�g͔>'?�K$;�x�!i����F�`�ϫ�I���*�+ ����>��2�`9ɜ��N���hz#��p{������ۢEܲ�r�{9ɘ<���F�I�3�2C #~���7�G�@�mXC~��-*v� b�`�O�?洧14��ۧ���e<��+�^rvt[�e%����̽��������pZ��)�w�.�s�9�φ�Sx|��%�Ҍg�~ ���A��$�rm2�����rle�*�\�����|���<"�c�$���L���}xU�����ᏻS�K������DڨמnBw���g6ZA�>��2�Oh|�����D�gF�Lh�"g�D�<�9F~���0�$�'�$1�T�u�q<��S%���d����|�l�=�aR؜�V����R^��܍Qy�,geT�P�ՍJCrp��}.���m���t��w*Mn[p"ݚ _o�vs}�� &0���R�I�W�l�1�C��u��¢���f�Hu[�z��Yp{D�b1N�]I ��h��7��ɹ-<bUPjt�99Ee<�6�Y��\�6nx޾d���>4wЧ��Ҡ)����M�p4��Cv��k��?����z:�V0*Na:��	�Re�6J�)���{�翊�sP9e�3!��^*&
��؍���W��+2��%*��V�7~�#ȉLB� �������yQHO�yl�C1mZ�Q��9vWc}K����npk#|��f/hJ��B@���U[#���u�� q�z�����.��)ĚD�����~��>D��j��p�i�R��3C�� ����*� �)!��%�8�S�W\lʐxрB�.
9�x�l�/�q��V��K���Iv�Ol�{ۉ��f�g�L*]Ǹ /$R��;ʞ��g��sP0K�+�
����-���57��G啘�[ͷ�je�C9� !S/��ʯ#��m	g˦^P�V��sk��)�<0��Z6pz0e|Om�y��5�~9�F�h����S�p�+o� �qg��=�iX}�0/�>*s�W�W��Ȇ��?J�f�-��m��ζ�g�^C
�xvl �2��#vt#I(2��jE]�5<U|IIմ�����ؗ��J~�ʎ��^�:�7㼠�Q��\}?��b�v��4�=��b������'t]�~�5AMY�����,!+�!Cql��L�R�����ɸ�m���k�+�#5w�P�[-�n����&�1�������*�h�}a�f���クYh��z���{e���۸��mm�FxQ��Л+m��2�&�\
����_�eCd���Y\\T���Q]w<���4�/����Q��/D������Ŝ�/����\Pp9��:�I�|�Đ(������`��ه��2�K�)�ˤ��uh�u�(]\�N�"�E�����8����hG��h&��5+807=d���h���_��R		�m� �@��Cw(9G3�e:�ރ@h�����
V�R�P���5x�������䙉0��(�����RzS�%��]�a C����&��&	�` ���n"�0(^�O2>4ՋoK�𾫤�8>����yёB�@�����Q�0�"~�[��O���Q�������v$a���P�.����1��}:j4V�6�8u3]���-�c���E7�^h�S�$�"?�iH �� �Ae���!��g��l�2������f3ًU�)nB�J�-.�B@������U�`+#.P[��}su���u:�o��H�ֆ�G���N� �LQ�d���09v�j�dO$9)od	t�w5�#q;�yY��#�KM?��� �����g#m5��<P/1�ݓ��~��B���R��]�8J'T���l/�~"�,�g�.^ƌ15�F�A1AF�:(������6��]�C�2���z]_xɲ
R�d2v�FQD�#�؟ؔh#���70w�%G��?�Z�����m�EH���倧-���o���-�h6Bn�k���R}����>�iܹ#�N�;�O�d�,@2���/���Rw���8��!�~C�����K0B��5��pYj�����ՂN�[�4-�/ų+C��r��w���Bx���\���(��T-b����h�����bD�ЎԐ�_?�y�j�W�8G�m\�29�*�Ą�W���ְQ���6�cĹ�B˜8�R"gz�`��S�I|���ԄgNw�@��{�����ףN�H]�j���=,�E{\��e�nŻ�~ �ٶAR$9���	�K��\̓�Ԥ:~7� ��×$Ic��:u�[ŋ����2�" >'�0�ūn�,�צzi�i��T�=����(�w)f�LJ�k!����JN�X�@d�R ��A�v4�c'�4�u}��n�6�jA�`���kw�$�
�>�tᡜ3������b������yҀ`U����ՙ!�c�A߈UV2�ʍ_ZY���c�l�-8��ß� Oॿo�'��[��f �6]�F�Ȓ7<�QA�i=9�tX���J�{m�(ŗ�`ӣ��K��H���*yG� ���7qy�D�A�T�dW+sk��,./\�d|n`��~x��Y�U��X���WqsX��h����Z#]�4��'�^}�š� ������Pq��~D�����=��H-�H�ɍ��fin��p����v%V��b���'ER�䣢��k�Q��>͞��
�=H ����s���WzɊJ+mK���z�l��	�~��)ڐ��������/u'�owr�;I�Gy�������&Ik�}��H�~3��"����6���(K}�H��V�J V��k�EM�Y����P[�/��b#�ԃ������TW�C�w�	�3�1��'D����U��/�np
��v�?�4	��P��x�w]q��;�ؙ!��8k7y�h��ﭿ2��2Z�+-1��Z���qjɰA�ʦ>�<8&���Au�D��T ~_�:�XD:U����� �@�1��-ޘ����"�dQ�!�:���ݯ�7�Ky!���a��� ,�(������zƼ��[�a0�Y#�1FZrx��d��w�"I�T���p�}UM��^�[]��F=K�f��6q��\����N�p������ki�LWd �u!y?�y
6?g�L��6������~�N|R��I	NR����xF��*t���`������%����M�YQ���+9AR��kǺ�m�n"2=�t�Y�#�r���,�<s���Ϸ�Ji�$le]6�Uy�Sx����5\G����G��Q��e����m!�	�t"v�
���5���,� �� ���,�U�l�ظ��w%��-���x��e�(#�ؙ���L��_��h_�,��R���t����������SO����Yq �2b�@�5�(���8TZ=w#F�>�t㶽O�RU+$E�DЫoҙd�3)ݣ���'i8��d�����m�sA%��j^��?D��q�窂Ę`�hTl=V�,���g�7
���ܪE܌(?�N�X�sM.��u_=�?y�s�uקX�mj�6��7!]e�pxRgʼ.P���^(3�C���j�2�R^SN�$fnayjM����9���`��<�/�հ��{`��o>�SX� �<�O)r��s�?n�=V��3�r�մ�$�]�����>3ֹ�y-�q���e}� ��U)| �LMf��1��E�z�#�]����S�v{�C�ڟ�M�W����、�Ͷ,�[������c��+*k3���wB��<���\j$,M7r�Aq
q��3�� 4�� D�3��4�=W�2���}x�9��!���7P|Y/���D�R9�i���+z˘��6�A�x��K�Q�������x���229��Ǣp����E����/Ȋ�5����_��8�dh]Yц����ub�>��f
�a<�7N��T�#�I!Q�&�V�l�����(������V��T�#e{�f)+�X��:�"2�í.|����Ký�kyp��{,]��������k���7��{kM�{}٩S���`m'����_W�{���7��%e��ōR�.*U`h}���[*ˆ��:���CE3n��+����GN��������27�%R�q�|��a�F
"��u�� ���4�2���p�O�&����֒/�_;�~���WR�$���kږ5t��A|��n������j�WG��2��k�4�v
b��n�4|���U��N�Fk�G	�����kZ��|� ��$9�`�����7H	���&�2~v��E�ۃ������!~��:�3A�Į���еH��J�e{[B�5=|	�[ia�I`=YU5�����:M����N
BZ.����Mg��,k��j~b�;zUUx$GDwEA\���I�堬�D<B�7=O��OoHX���p>$[ھ�
�.C���p(����z����1�`��@�)7S�=�!���B�A�L@a汽g�Z;e
�u5�WwV�p���կ�	"��,���� \���Z��X��^�s �%}u��9%L5X�=��LV3DT5a��V<)z"�+83��ګ����0b���ӎ'S��)���� � /P�ǫ7Ml��'��V�\N*IО��mkנkS��w�09�*���d,9��K����d3-�r��7F��-3��Y)!���1�{M0�mǉ�:�mq�/V�_���T��S�"{���'�捻V��F}�S�8/��O���Ϝ��I[�:p����$rTBcT������	�~��/r��+D���ˮ� ��uj���^:h�4��e�x3�22�ҳ�lF����6~�?&4�ҝ/g�حˇ
�J�}���}gO����8o�?{�0���-}�1V	������~����ܖ���L�b=�X^��t���-�>t�xn�pLC�FJ��"b!L>�=�����.}�~q�A~�  ���9�-�p/����&��\o���v@�_��D����ۘ�D1:H�=LS��f�+�K%9�^�_���F$��$�S5]�wMq��]f����+0ꭸy"@��Kh~#Z���%��JYQ��o�Z���[d���.Z3�n;c��y� v������JV��qx���\c�Hte\xeӀ{g�?�d����v�Yt$��NhY�NU�!t�B���+��W2����5�$X���I=͜��������xa�$��v܁�;�%��C)� ��l�*ȶ�����Zd�t�b@�0��ؤ��Y��������ר�$K���;;�^<��"Փ�=4F����lI�C�<�53eB�O#��o	������L��q��z��4���Ι����V��u���1t�Țǟ�P��L��&�hi�j���C���+e{�PV���� a��^G{��r>�0��k���t|5�c����[ �k·j��eJ=�G����0�~Yȵrp��(����*�k;����\�i��F������R����A� ��}����LR�_�H~{2�O
.PчSutY�)T�/���
F��> !9��x����Tz\r��qH�{�rr-{d��
���n|2���>���b=3
Ɵ�1�Vv���`��}�!�G�3U6�/�'�����)uG��!J3*�-t�~"7��{��*����6���Аt�}|<��t\3'��:�rK�+	���^��k~��ޢF���+Y�g���S�~�hg��y\߅P�*�Ԍ,%�8��_��Ef8}dj6�X�$}}k��+�V�ct�RB[(FSK��6��&�#���A���#��kP{���:Pi��fK�����<{i2���V��f�-m�L��O�).ه5�h�8�b���ؼ�T)-JM�_s@9h'��{U����{�>p��,�'ݽ�ĬE��y���[���ȕ>k�@l���8KC��D�sh��u�āx���=#��ipƑ�S]��M8k��m<.!Tv/,S)���~�	�:�����sO)���lK<-� k;��c��c���6D�i�L�ls�uR`t�Sk�)&�8N��0��q�Ŝ_V�D�\C��hYQ�3]��C�5R*����r���V�*��"��0�*�V�tC���Ӄ���Ts*I��@�9ωȔ��8`%�[,�
�xD�f��:��$�鬆n�jD�Er<޾�m��C0Y���_�[��ە�&��\c���L��*o�_-�Rפo]����ˈ"{i:/=�Dk�6��{ӄS_�
w�Jr�&����ǑE1��껊��IܑѤ�z�g˙K���J�r�:��E���hdl�Lb�Kmzr�+�G{{Y��$9h�O�(���8"�ޛP��8�j��H	<w�ELۡ��w��?�k�uʹ��5.��_N�(�,#Z���u�T,E�X�g�{�A���l6���/.�7�!�w�m�yg��ˀ1�c����I�r�����Oqת�(��o|���s{ST�t^x�'��ujG�}]��ޙ��
�|���9˓_[���^��z�n|�1HC�"�h܀ح>&���Ԝ�<_��I���=g�?]҈�$�w��%BAQ��W~A\��ë�ˠ�e m�kB�&i;t�/�B==��8�SI�߾�b�:N��%��I6h��s�v�	�mV�y�$5��<Þ�9�w�}\}�Oi�́7�(Tb�tit�|���S*�� �b\�p�R���q�-�:!L�ҵ�Q4O��%>��1B��x�J�D:|�JB_K�	?w�q�����H�Nt�����Ì��:I�y�b���?��{�9\��B�]�<��Dg��[�Mwc߬K�9�$
�"�'?M�^�惧3Vo�R*`c�qqcl�߰�e��^����Ơ�=t�OgK��t��Pz�{:�.)��G��Փg���똄$h����*��Uk6�e����<���$��
��h4-:H���6���E;2�&&i|��<r~b�v��4"�M{A��`���Jv��s��\r|�!�����F�J�N+�>�eam؋��eop��7N��yW>����9�Z?�"E�z[Q�{M�*	@�y+ʶn��+iX�����d�hj5ݧ�Z��z�L��<��٘>�%y���7mh[�$��=I�ND=0B	��s�,r�����?кa�1��6�4�5L~O]���7%��o/�'��` &��n\�ԃ��0�=������b�`_Fr��ǖx����<�~�<m���s��t�#p�p�ZB�L������r��1�?T..�W}�0p�H�+Z���;�0:�Л:#'%S1�)�%z� �jO4Dn��|�}��G���[+�gTm�Y��zs#�ߒ���f��dvh�J5E�9��X���D������ԃ%W�%݄��r`�(c��̓=T�Hu�4V�w���0G^ �����#��E���V7�t_qq�	d#��^1@g��N	��YI��@+�m��_���όK;n� �����%i���4�A.ƈ�������SaY��LX��q� �/����މ����:�K+��sIP�O�W�酾�Q�0�Bq	����J6,���tL�CV)�����n���@�Qw$u�Zq�������H�	�z)�7��}>�/�$#n���J@�3��N@y[fB@�U-��2a�o<���W�4e���R	����ӧ��^7l\$*^_L:�P��|�"v�[�{H�t����Rr����m�mt
j���/�v�+}��m]o��lS�Y�ȕ��`���Ӽ�1����d�t]h~�}�o�����0�3h���o�N�rd�!�����}�J=���Y�5@�l!l�s�5�ӝ+.�|�E�q��A��e=c5�(V�Vxtm�����4+���
�N�0�J��<#���و`��˕������4$o��Q�T�n#���uaj+�&�a��o+���c�K��c]H��Z�KOj��]�3���������]'���L���R�Oz�V����a��ְ���D��-�r���$M��{�ޮ(�HJ,��`lk2�Q�j�Oȉh���v4�L�m�R/FXdnݚ�m���^{� ]�N�$��C_���.�y���+�G��C�����e�5����jF'� ��
��ތ�xo�t:y߮&D˶��g�Y��P�\��X��o��Q2��&��~Rf.e��˔�4Rb�Ȼ�N����Ra����F8 e�Q�B�ph�wI#����"N�4�7b:�#�U8��sċO����h��̈́Q��5���쏲�a�o��>��=;���_�>:�`���7_���\��jn��=�JuV�y�-��OvN�V�4�0u���Ԥڝ�f'���MF�q^ׂ_�^,H0�].	��4�n�W�&""����/�4p�������U���:���⮐���&5EP�M��a�����Մ�;�7b�l�'�ު�������S66� .��3J�1Z��7($�O�4D�]��r#9@��]�2v.n�C�ϼ��y�$�'*^.��Lõ��&�h���߬*�uzv�`�c�ۀ{�g�H=6|�6x����:�����RXKW�}
��M�Pno�Zz�*G#R�e�^G��uC�郈�[�+a/�����G<�b+��b���[���
mN>ʁD�^�J�"(���C���ݲM� ԟJ_8�L+rN�֘��7K�>����n#�ʁ;Dߐ��}ꍐ`)4F���)���.���ެ�#���k��jg�L�b�j�q��)Uh�� �.g��W?�����_R���@� K�S[@�����-�.��7����^��g�w��"'y��~!7΁�A=���H���p��p.���w.��7��L4�G��'�_
����x��&���;��lЕ�u���y:뤡�:66�Ώ蟛� �ƈzA˗-N�օhǬ�&�Z�P@z�w\u�5��l�X��`�J��=��n��n�:!�{j�r�g-�ׁ�� �i�*o�"P�/�8�n�^|�K�t��޺MO����N*�0'�C:�ļdM�x�Mv�v�.
�E爮��u��茩��:���Č�]$se�(�E�m(��m��<�w��t	�8k�l���v5����U"$+;p����h����8�o�t�9�0�i�@��tV��q ���HO��r��D���B���B&�yy����N�Hd~����=��P�c��2��1+yaFF±�,���E&2-��Ayc����#5c�:������G3�Թ5�1��:!䟸l�`���M~�D�� �2Yio�F8SA7 u#��tN��Č-����"�0x-�����f@fma�m��k�a�|��__�C=%W�1.{�� �Դ% ��k�] �a�]�b��tbbC>1y�n���a5�N*S�-���W��b]x��L�u� �ޫ��J� ,Au����~܆�����7�Y�z�&ԃt����s ���]����|��Qf0;"D��m(7�������3�@��|:����t$;<�z��{8�	�:�c�p�I�����R\�$�cp�����D<⋚���S�24�E)�����\�F`��������$n�Ę�qsW>s��͆�u�B�ϭn�Yx�b�M�a�{�B��<��dd]�s+F��Yn�L\�Y��px��0n8\MNGCCr�fl*۫]l��ZN�ãbͳ3'���Aw�z������*��*��t�K� ��j 	�[�I��8t]	���/�幆��`�G�Ph���Nt*F1V�_ɽ�� 7	�q�#\MvUC�Uqq1Ҋ���CŚ;-�Ւ=r�g�y����ӽ����Q��۱��&���(-]q�����V��]xX����;��=�8�I��I
���^�u���3s+���U��-)�a����]��s�q��%o�iD"��u�W��O�8��u~1���'��i��K�װ>���;l�3�u�fj��$��~�z��To�6R����R�����Ј����`B����걲�l�J�Ͼ���kKL���I��Un�����H�5c�5��;�"��my��ej�%�~�͝����v�8=�x�1�s�{�����-F�EL+�4+�}P�����(Y��T�#zgt`<|�Ap���e�8�QI�4s#��U�)�ӍSݺ I�<�J��\⯂dp����F2�5�(���CL۞�����V�W��Ū��=�(��%���_��$���шFf[ya�7ϥWC�4������R+�PF#���7�~�A:���/&����1C2��0=�{�ڕu�+0� S?8<�%�����UN��<��&�[B�����8Z��������s)����1��DƄx���ށ;��Ę�ï��;�$��O��=��������M��:f�|Np��
Ɵ�Ri���<�w,��u�=	\�u�#E+��?	���T�`�|�r����aO�m�*K��;�P2���xJp[�SF��?��ɒ�;�pY:�ޘ�H��v�E#*�KdcܸN�z�
����R׭����*^5[�.k�����!�V4A�ze��\U.�24nZ�̀�����G��1�,�:/����R]<+j�խ����������Fa�gW�A֥�VǄ�1�}E������
��E���]����˯��H�&�E��J*�}���H1
H�*���ܠɓ?��5�%�����5Gh5��
c���à�jב��Qf��`��5��G]�|y5��M+��6�) f�G��"�P��kL����y�54��pc3�eq%�M�G-"o�b�i���T���]��`� C|��t��9�#할`+�R3j�:\1 �G���D��,�1z�Ҙ@�*T�y�o��ל�5���A��'b�qʁ��S��I�TJ�GA>� �+����d|�_��W>�A��`��B�:�}q�+�l�u�{�q(W��F�s�}� #�����wnN���w�N7Ab���	�����㹍�lLЪ��q^��h�j���ڒ?Cb'���Px�jn3fD�迸S�gLCZ	-�k*T�fb����ۆ�&ܢ�L�hS.;=��(J��6��Q.����B�4[]ɐ�M�\+m����GY��!e)!����=�Rw��|Y�L�������!��w�9����	m\8xv��x�6rw��a�}.]��o?3Nﳷ&i���������<P���S�o�꿳��nA���˛Q�C_�Q5ג�N$��Ќ���V�#_v�����Ye$^(�l�s��圌��#�!ڎ�~6�i���I�eh^��]�.E~O�β����'k}	��x]��$h�f-_���᭳P,VG%�&x+�? ���G汆d��RH������}�o!1��;[��5ٴ.�/C��QӅq��,yDw����p�;{6d�;-gΝ�p�˓~��)V^+�azOy�Pk#�[{ȷ�a�S�+ެs�N�^���^;�V�0?ԯ���"h�l�C�ìm?M��F;��
��D%Z��vX@$�$������	�����m�aٽ�I�6�g�|�� �_H�7�		�Z��wݟe�d��E���pV�p1�bKs�0 r��od*/��8l)��� ��/nԈ���m��3���"tY��I�*�#f�R�B�Z� �zܯ�����ؾ4}�����Щ�d��2�� ��7�A2��j�����p�@L*����J`x?�jJ�I�;񆕙�̺v����ݒ��43�O��l)����3,EO���q��r��n8ص����ͭ�� �VVN?�*��P�i�Ir �s���}e��*8DTA��v��$��Ob�3�}v�,�=>���)�����v���|S��*��jo����A����[h,4R*~�����IQL�Ո�ӵ��&���Az�R'�6� :.]R���|a���#���*�̈́x�zq�e���ǿ8�G��=M�ХD�2��QF��XB�A��R�@�h����hKN2�y�H:K~-9�:e�UH��Rۏ!�4��Xk��p�/#�:�����`��~G�be& "���+
B|莠u�}�y���U1�g�m�y �̉�?п㤑7%U?��Ylt���� ���V (k�l��s'۫�QX޼�
�]�b��0�}�ܱ�@��sh�t����9�����J�_���#8��@㆕�tc�5X1��Gi� `{��ߒ=��Xh�.@N�f�BǗx�v���g����g���|��S�?H�Ө��J\�u�M���g��6���Q�+kY�K��t��wnj����-�����}'�\P�^\ģ�6�hT��V�������(�f�É�Sf;ğY`��)#���h���IA"��N vMǌ���FX�l�+{|�@�K?�v�����}.��z����h��`�\rz0;9+���0L��rEi�|����uPW�=9�����w�96�׮%�Dx%�g�1��m\Ǖ��v���4�1^.�2]�{�R����j4�GQ��50�V,S�^��,v�_�խ���Èp�ڬ�?:�A٤�{�c��hxt���G/e�XQ7W�3t�g�5m��C���5��m}��Up�jm��\h�I��)8=��������=S�-������r"��)�F?wv �b�q|3�(�m�>P��̓��]R�/4M�,��+����L�o��V])�fn��S%�c��j�`�#KҤ�FM�(�?�d�'+���ہ.��-�b[��JY0���|����k&�h���@�̸Ѧ��/���,��K��H��;}3�>0JF�?��_B��P>I���+K��M7P�=I?H�ͼv�qP�N�S`�D�f��$�z�9���M�����E�/�a8���q%�D���9� ��]����/z���a �������q�9�� �$z8��l������!*����@t/|I`�i-���h�I���g�M�ھQ��x�Q���#"*8֑%�EV�k/"ൗ��x
�z$� �x�+bIC��fk35���I+��5	G����d� �*o���Bq�)C��ėCD�4%��'zup��RN�l~��A�U�Yv�q�g�#D�Ļ�L�N�<�J��u�YT9�����D_K��R����|B��.�\���R`������r�_}��wb����rJ~"� �Z�?>O,�S�d@������N��a��hAZ�)}�U80W_�Q^�o_`u|��g��o��q���3(ML����;//�
���Q5��+篝��cCϱ�}�:���z�07�5!C�+]#�j6.tj/^���R�3$Z�nʗ�����H=�_q`�J�+�<����yu'*[�c��H��)��]���)�*����iƄd�6��9�rw޹�����@ЫE�m�3���ԓR���R3����0=rp� �{��x$N��*�ģ ��¥�����"��(R�Z��u�4b�6�b�4���������B_����Ӹ�ݦ1��96a\���6�K.u���uW��ʹe/�q�wL�]G��~<P��0���o��C k+�5�����P�!.����wI����G�Iɽ���pH��������R˾V��K�QM��zwZ�`���pbu�	��ע|/.LC�'���)]T)I.��H0Iی�Z��}��R�-��wf�̈́j�tn_xuyO-�5Q˽���|��')$	�͔�?c��G{H5S��S 7v�l��:��<$�5�Vy�2����R/�hM�#�շ���ow[Z÷d�%x�iL��^��zi0�D�輲pW;�Vta��\�M�!QH�S�u:DC�3�ІJX2��A�%J��⹑-V( /���-��
�4�Lm��l�j��ə�߸"�n	H�3��Nc�)=<�z�~���W:i��|o���ې~�F]X ��ѐ_\�p;D:�;?�9�H8��+����`V��W�5�$KcKl�P�h6�mޫ����Us� �W����%T���4��~ԧX=]�ʻ<3�7'D"�ћC��K��d���\��?��?|���zַ|[�^s/��/Nd��v�,��ḙִ�b}�� ��}��L�m5y5�B����l�L���-��t~��,4��q�j}���WQ��f��G�Õ`�=58���9�U�J�ܡ����K���9	\C(�����������WU�iU|Y�ҟ>70^��~�F���%}���Ϗ�D��Nl�8Q�t`w(ۺ=#��;}>ט6"q��B�x}��z�H%��9F @�B�Y��ƒ�7IÀ^�k7P�;��1��7<1ʕ@-b�o�0�ˆ�Qb���DA��͒��ه�%��G07�A�^��n_W����1�`���ӊ Ј�(��gC�TW�g=.�m6�1�����[���!�f>�N��=�����Qk���k�`o�_W��<�{��EZ_b�O��+�Z;q8�*񌃳k���U��mQ���V�]SfV{�Z:�w%�dJ>S�f$#9�/�����9�v�2�(�dj �ZH��	�	�#�\�e��62�jˋ��V�&�������*5���ES������[���0t���V0�}�fo b�5����=K�n~J~
$���VLN�eN<����
`�o��&�Um�+�H��O}j��OM!v����L�#]UyO�횗e�}۸V6�fM�'�KVik��-�i�h{�|�o���/S6���	�V��4h(�vϮ��ם�������~��8l�,*SpCΜ����q�!a-k���zs��2m��~ l厊T�c�v���~62�0��G_;/�8�AU,Ml��N `�;�sd���ٷ��s��/����^Y7����"`����
YL�m��o%����.���șXk���X��'e�GW���H�o���6(���f�Mш�j�X|JDl�l�ab���1?ݑ_V�����5���=��d>+��8���8�ϳ���e@Ѳv�\0h��lt]p�|_+�7s����L�����0�OiKr���L9�|�$��o�7�T&��@qjjj�MM��6�+	<I�t2���ϗc�b27�����Ȱ�y]JK-0����N"=E���@~��_�,�m,�!��T'"��W�I��f�l�9/���x@V�O��T!)�&���!{����CD�"@nH$����ͧq `���(����:�9�!���C}�^���cE�~|��H��~�����l�q�!��㔪R��?6�8Ѭ��!X���6B��l�E���"kj�q^�/�p�����3�����:�E�~a�W9�h=�a�z�/8$[I�� ����,&�1jX��u��XO�μ�M�d#��#���hfӊ M�C�~�9DA��~[��q�0��m�˅�Ȋv�r޼���0���6��iG�1`jh��g��w"$�#N�"<P��[�e��3ިͭ���Sq&��� <"��f�P��4κpb��O5��X�֩���l�f�zƍ
U����9��W�vu.4]&���+�0abBT�G@�V�j�0C�5ʀbvE�E�p��S��=���O�>���hz�7�c;��?�V��'�,j+C	2}gU�՚�oE���5o瀥rS��������g7ҥ�}@sK��y��
��;��P��O(���~��ȾD��:�s?.}B�RRJK4���g���ɿ���iWYV�G�px�V�a��X����JT���cY�Ɗ������18�˅'��i����T�
�˼�G�v�}�Qd(�#��Aؕ��=!�F��O)@�*כ��D >�S9���>ֵ�Z�<h���xί�&�U���i"��NV��U�gz$W����e��n�|��;��?<�Ƙ� �gB��#�y+v˓�D5�Lb�BB��J�a��n�b&	S�\��	�O��v�(���	����*F����/2�boU�S�ms5
&,�y�펡�E}��[^�88�� ��B|&:rL"7D3�u�i� ���	K�%� <����=�'?{
��U��(��N��JK_rYP�����V�F�J$�\�T�]C�S�._�I��_�MU�*��49�O�I���[�7�����0�`4Q<� 6)>!��&�U^�kb�	&���
��ڛU�1[]�K�~���V�s�n��&p���F�W�D`�<��Ք�/R~�<�&%7G[�� �-��4S��n[r�4���s�����]�x5Z{H�Թ��G�QU|3VZ��C2�.%s.���۠���d��x���z��6A��4�"t��O�&nf�Uߒ!A�v��q�tV��(��90�	̓z��Hd����S_p�)�B4<�4f䶼Q�������`�n��&ɞF�Vq��m���\�r�^u���{�A�N�� ���h
�,;�����f�F Oʆ'�
�w���Ir��~}�y��"-�YЛ�)�#�&������k�Ǳ�oM[�9[qּs�RI�Ò7�*��4����	�.�s��,�wL�7��_W��y�	~��QM�$ǴV���}y�t(�Z�����0�KA��\Y���9Y�s�18H>i����'���|��Za� 7W
�����Ό���'�'�KN�N�k���0�"��?o Dk�l�#z���OA����Gƍ��R�隡����jg�N���mԔ-�(�/Q����1f�$�_��Uz����7W���$2�*<1a��m�}�=�����q���輓CS�p����A)�ĭ����w+�6$�#]�����X��uf;�Var$�7FVd��H� ƹK7���f��8l3n	� ��/jH#W�zP�k�j5y�Ԕ��&�G꒓#ɫoKo,H���~
�6DOt��!l����	G{d�O�/�ubx�M�)���ׯrD�Xg쉬(��MN���ξ����z�<;~���W��6��G�H�B�y���g_��P����I�Q�Dy�;lU��0��uۢ����[�-���o����J��o�g� Sh;�	�Imc�6��V����2�V➒�vr�eƽ\8���C�����MX�.J�1~D��&��JgN��6�*�?(&P|0��ɱ�<	�u
�|�p!3)�����6���$�>�63�y1�/?���Z���L�Ok�R�
�a�\���n΁H��̘�C����.���?5���J�!⺰����{�Do������i҃��
�?4
v�[4���r&�����6��ѸR'W��zj�=�������mR��c�f
���0�3-�E@K�m�"�I��o��wis0a�V�=��V��]iZ�!����Vĉ��m�3ՔHt*����枍gR΅�l��W���<-2�)�9��òa�Q��8��d�����ł�Z{/s���1�� i<��oQ�k�)�ƨ��|�%�$�;����Cy�g�a��s6�9��uSe�H�7Zm�jC%���h�d���Qc�%���!��H�����H^�2e�Vk>�����ӭ[!�T��u$ɫ�
�DAy�	��Xn� �o��`sS&d$vT)R�K�_-��y�&?O��'�Y��#k���|�EFrx(ym�|�<��AVM�,�W=_j�Z8��S�|����how��Sڸ�x��� ���sUkS.��|����!�r�����U�ǒC�Y�[�C
Wcͤ�
[8Vi��`Gu��\�|�b۟7lb�*���%���9Q�.bB^Xª�ӆ����n&��a��٧]��a��Ƅe������I�7nW���HL00���D]>��ӕ�s�vƵ�t3Y�X�*u�iq�p������ *��G��Wp�1�������ս�z�7:��t|?�:AH���I2�
d�B�1S;E��b�vcέN^�����$��v9�Z~P����7�{}K*{�wB�e�nL}7��D�O�ve+1������ϷTb���,��� ��ob����*�Q6�[� T�+a;i,\Ǔ���������Y�Ewg�KLI���|:���AtA�]*r�GB�Qi�+����b������X6>��tĐ��<N�.�%�s@ �Vʓ+/�
����K����9���}�����H�B2�?�|��u�<|��ID��b�o.�y�\�W<�v�$���11�>�X��C�-��]��������"n��TW���*xd��!���o��ϏL`���͔�7�G�����Fo|�孽�C�sP��;�p�/.�N^��Y�p�A�9R㥚As��Q��@���.�U+�!���jE�.%����R�=�D�4�[:*+��B��7RL���/��	[����3`x*8ZmHl<�j���͓�S,�����/�)�.����,�o����P�X�;{��ɳ{=�`�b���N���H�����4YJe���&�x)\��Q�9ԗ}�Aq�+I/�s��׸�OiC2�14邛Y��nɫ���'lO�*G��u-�D���#A�Ր��8*����.����7̉�u�*����S�0n�_8+�/��d�e��_�@
�W��G�$�2��y2%|Mv���gH$������
�p�W�<_.����Q�_ /^������T�}��X�n����"՛e�����U����`,�J�|���E��g�ne�y|>q��Ӱ'=�,�i�B*SKoM�7V���l���e)���\ ۋ���v^[?P�C��7��fnN��)w.�fXTz�`��U�Xl���'fՆn냇�2�h�� j_8ێ�e:�xX�b��q�tЀ��s�O�5U�C%���i���a(R�Mm�i�)x��ǹ�I�
"�n����p��B^��ڦ�n�!JG�����/%���0�7԰�wd�T͟��97g
ܸD���m�_Ć�@�n��������gF�J�Dmf2����>�/�a�� -�\��Q]Un�ósO�@�c��"�Jk~<�[�^�B�p�,z�|b�z��!ř���q�KRN�4����V��G]��A�V(�<��ee]�����l����Z0<�2ߧ�a��vJ���U0��a�iq����D��̗D�ρU�	Ϫ?��Փ���tW����Ư���5?���(�C>�)Οȭ��I���H��`K�D��9Z�p�30K;VL�#�����(��+si���d!nt*����;)Ղ���cS�&� �M)V_�c�F��'/7Y|2XS#�h�c��n7~�4�)u�V�k�е$�>���6��������&���bTx��o�qtt��s�(`��1��$P�]��Cj�f�R�ȷˊ�í�X�P�>����6�숒�N����Z?О �
D����\�:_���>~?�q[y��BT�SĽ.Ёg�/��+ǳEr�[!���E5��D2�z�����E/��1)2N�D=`٤�s�gQ�����Q2\�2��S�V6����Y,��5�/)ɔ�.�9����-kt�FΪ5�?�*�6�W��AxOv�Tʷ�lpPRv�r��I���vq�i��#��}�7�Yi�7�ON��Bl�I��Zˁ��I�\.�W�oɔc��M~''$��E=������h����n\ӎM���qܖ~XYw ����"�L�'�+�d��Kr L�g
&��#⭊"$�����b��j���[znX��~l'���Ζ]�b~���k��G����� �d��]��o��s�'�-p�?���� �.��>��D�_�8\�˴)�Q��	
��n_���Q��C��.��1�KK��Jm�T�<�^w7�>|�/j����J2�g��'��J�����tG8;!�Aۧ\[Л��b�7<�:b�A� �%5	5uт3g��H�F&%��J�:�h�N��ҥf!:xU�`=�t�pQe/��Ђs�=ʘ�����z�	ˤ��B�)NLa-��Ӂ�"A���['L幭��-�Ǣ6�2g~BO�0���5�D"�ե��+��a���rEU	�H5!�0�tyՂ������>,�w�4��{��2�����3x���>\G�_x�� ����_\�Ç:P�|*���卾���3@U��s�\�;ڮF�N��)�������<��V�&�K�	�2��p�"!h,�J����-�К;#�)��\�&����t �Q:����FEq+?4|x)���� �r��	+���0�'O6m9-�m�����Xj�0�HSv�`q���9�8��V��
ٝ](���	
��Tb|&�@;j{0�R��<jW�˲J�4vyDd�qmYL�%�A ����HТ��lfd���I���;�f5��V�=�����˕���_w ��S��c8"����Qd��"�L:0!2Pb��[Bg�>��B����=ME��7�V���*TD�A����L�j-c|B�!�	cF��Z���V	���.�Y�W�m�[<��ƌx�c~��H��mx��U*"���׶�r7NQ�Y�^F���T�ǋ#���P�j_(�Ɩ�q���u�ac�o���B���ۻҿ�w�ׂ��[�}��Qh~����`x	��q��f^R�4��`�ۑ�sp���G4,h�;K����`�0M�21 3�:�e����P���_��f�'�l�9��h@�if����@�=����-��(��?���/��7��(�ZU���P�:Wpx�^��IS��>�δ�{Z䂌�&1(�*�s�U3�ăp<�X�yMV�4SO��|}��S���ТEGh����g*��)B}�M��84�]+��rEH�v߳[>����vs
x�r˄��SqKAF���̓�ݬE�M�>��{���qG����M#M��Ӂ�+][��0������H�3��YT:j�q�_H��U�A�����_4��N�-=��uO����Js>�8��<���Cͪ�S5���P���	���(��h
�B#����CtH�Q.���+5����S��rr��{ߴ�
1U�:�I��bIE?��=>�����1%����˝��	���x�B�B�XjlJ���Єs��b;�&Z��0c6S-�� j.�6T���IJ��,�@PZy%�/�w=���r�Ł�d5a���2�5������G]�`�S���� ����ӥ���F56w~0;Y��w��L�'��h���H�vhyz��g�-����Z��f������`)��,���feSL�o���	���>o�D��r����&,�t��A�8��|�r��6Xىz�x.}�g��>��kMؖ��T�c��1�e�V�4)��?x�ދ��Eq�����L-�No�m'6ьL��2�zo��<�֥��I��{c���s)�F�	����Q~yQV��3;��*���d���	#<�^�TG�#�HF�K:`���ҮΠD�}5"�{X��`��j�����{U�.��]p �}ie׭�'L�kG�;�d�� I�	T�,�t���O����6���S�ԁ�u�M����ZQz=��C���>��p�5i�� ��:��T�Uy�`�O��p�x�X�z ��3W�p��@���D:�P��7���s?��5��3���;f~��!leV��g��Ƚ�w!�3p�f�h����E:0��{B�ٳ�* �yJ%�W��y�1��j֍e/|�+ (2V����e�/���1~n��Ė��~����w��7y�_�2�E�K�{��ȱ� ��իp�T"T��0DS�[��)sbD��bb����PG��7b�8�$���L��tA�\��p�63�3P
��cX�p�͚j��m�Rst�y�M����(o����&��L�G�:��y��{vG��Z��\`�s��������Z<��ԉ2\XѶ��rv�gU"��b5}�,�%4~1����.Z�LEf��:�C��
f�Z�ūb���W���f�H �j>v�6�v)7�\����=�F ǿ�.ߒڇmD$`!�q�p_�XBA%�\iĂt�d���;�~�����H~��О����9�"�͘�����8P�v�\�y�����M/��x�l7B5~���5�>���0�Y��EM�}$u��N���C(&�[m������=�F������L�4�O�A��|��P m!�#�iL6���1���Ki���;�a�Z��Y�p�����x����Z��;�^r4�����34i��N�mVa*� 욤@H�s�ej����-���6+�]b<Rd�E��ъ���S78�Q#�4��swS�h�BJ��|��X��׏��\Ϗ�y���3n�}\O"�2�WI���[48H��k�Ϥ�G��gw�n��4��� ����I����S�)W�Z��h��w8"�e�?��Av��T�Ƅ�>!|M
���m���tH}�v���t�>䇌�r"��?�'���7�W8L���c;a��׾.�d[���X,"����Y�J��cCUi���E��)��bmm�B�@EN=|[o�d���<ےp�iz��N�*���W��7f�^���`�Ƶ�o�!�4��(����"�5c��V�ɿ�Rdy\\j�����R>��Q�0�S�gi�&g�"��sǥ���x����x�Bq�ͥ�CA��Z�Ͱ��}۞%PSN����X�1E[:�t�q û�J�� g�)d����CA����)��SV�D��e�EWʚ��� �ԐrsV�m݂��jˌ���+�Hb���,�:>#)k"*����^��C0A�R���F3�rS�j���2�%��
żm��0�rc:Ɠ�<aQH&H��A�n9FRϬ�xc��I���/���6���A�(=ޖ��Ae'EL\4�3s�jL0Ҫe�ګ_��h_��K����P�I��g�k��̢��`e���W�P����	�E�Ey����Y9���(�BG�8�;4ꢫ��o
��nM�ꬋ�}a,����e<)���Q!��@�|�D:�uu�lv��O��@t���:�C�nM�� �-k��������U�g�8ۑ��#�:x>9֌v�,��3�qY�����F�%���x)�c
�ѨydX�f3/�
�|)�Iw�e��dL������E$\d4x�y��j����ʪNPJӼ��o�vFE�����/�%�e-^�8?���Z�Du�6ؓ���0���i?���EZ�����G�G᪣@�s��{-��'���e���X �Y<�1;�4�/>{�gZ0�d��6&�Yy/�H�K�L��40m}�y��&+jqx��D�d	�v�y�š�F�|�
.�H�Jʠ'��I���s{��,v$T���t��OR(������~�%���/�U�C���R��=�	��L���\���é?�
pO�Ӿ�0S��K�*�L����ˌu?�n�N�"�=�5��Q�}�������KP�#��) ��4'�i8ډ;N��OۤA|�t����� w��&����1�[E��10m�N@�uK8�:&#5,؟�3),{�$(�r
����&���?�Ab���/z��m)���t(���(bO������E�cs�C畻U���c��(���:ow���)UyI�����)��(	hF>�t�����8���bb1҂��]�Ǘ h۟S�ل�d3�(&+���aS��^B�1?�|��]4�#�@&A!1���h���3F�;ݾ�don���_Qa�P�B��t`}����#m�n�٘H���!c��į�qō�&8J��5��|p���Xx����:��2t-�Nd����颕����o,���W =^���~�$�}��c���;0="f����ߑr��XV ��K.�1g4�aSP.k����E%��X���N�.)p�����5���X�[���W�B]jZ�d���z4���W)��;"�� mԭ8�{�ӛ��.���8.�S�h��k��)�<V;�~������6|�kZ����+p��]���C�N�e����C�m�U��2�������`�ƒ�SL9�^G��]�x�� �ib�Qg*��i�e+��Z+�D�� x��9�����J����l��b��Q�ۜ#�ڇ ���=B�!Ϧ��
��f��ꎮk��Q��b�U�g{n��Hz<���KW�<���$���q1lq����"��m��HX���?�_E�S�R9r�@X���xOl~��ㅯQ����>t�W&"�+\oI�"���l^V8���&�/A9~�{� 2�N栙�%������`@2~���|�4'�rO��]젯�u��N^�k�D�S�F~ޕg<9��N����e�x2�L,�K~��7�tV�2�6f!��rf���xIfz�}N,(6R�k:��c�c��Wp|`������[��z�:��fD�?u�r������׏�\�/���4=����!R��F0�,�T�:��pK�8����vtn~�?�sDf���Bz������;���������Kd3�mmbb�_�ߚ���緙�\�@G����"=�We���n�h�N+�'��{Y�h��w
n���ZK���;�9q��1�F�[G��˻�3�Cl*��p�y^�jO�ᨕo�k��g	,Qt��e���3��h��%�y�I4��xNB��3^8�\"�R�+�_���uV�,;0P�!�V~F���r{sX7�����.g%�����>��T�>�4�
��������xJ�s�m>��)�L�9��8��|F�K���;�1>�	�U�N.X�	�e1�/z�����B�|1�CW9`x�j[�k��)�����*�by�G�[���%|����1S�7vM2���������g�����{��^-!��P�H#�ג��{\��:�A2��i��k�u؟g��F�[�6E���{{�}l��utǪ��Ѳ��`3�ٌE�O5����n���J��,K�%G����x�C5r���>*T���n~��Q��I[m��'��Mǌ�|���>%�R��G����C�"�o��~<���՛mw��^hF�!u��u�	.C�T>��r�n�N��[���������w��	�b=�����!E�E�o�t�H�Hf����V!�c��=��<�(�Е����q�^O�8�y�9�}�Mϴ-Tp���GK����<@o!C��a����Mvl���,a�=�o7 j؞v�4�%`~�w\�?����6k��Z�1}q�8vB�jID�XUGpX�إ�u�԰�'��~r	"3�DkW��C� ���Rq�O/�Jn�;��O��)o��U��wN;�\����G:y"���xf�������{B��Țm��/y,c0�ѹ��]��|�{�Oif�1.U��<�~��ά#�2hD��7����ز�K�8�^�G�8�5��"������)q��st)({/?7���DO�-�k���������%��EU�ݟ�^n* <�����%7�`��5ߠOhI�����Ѯtq�/+lʡđ��>.�y+��q�<���[?��o�ʚ�zM�I*�'��%�T�{�ֳXl�6�j���>a{���u�����ɑ)m}n|�`G:O���*"J��?Q��i�Gz�;��+=�t,#I_&��J�rIl�eq;U����/� g��(��4�o�(lB��4�q��S�ֹB�3Rb���^� 7�/��n�K���U�����a]�3�ϛ�bqٿ�����8$�}��E��w7Aa��=�몱:�w��O�:_����T���<^��`�#IǺ��_�y��H�T�6�/~��[�.�[s��sn��T��e���ᒈ��j1��k��L+O R��"��Q�*MC,X;TǦ�Z&���|��S�ރ��*UsO�@s�(;�é�}ק�˿�Y(�q� v��@��IK5 ��n��GaVqB���&�F��憤�֋�z�J�!���h\��,0��mq��e9g"[Z4l�)Ķx��#�_�� @�:b��m�U�oD.l)&7P��T4�u���O&�
��� �n���1�Ү�_cD��qj�1�p&�s�R��x�\�=��h��G�^��i��s�Z�&�E�tǽv� �Q�br������o�����B��&�F}O����%^���ט6���K~G�T���ݩ���U֩�~��o"�bׯ�g��!�,�)p�"pN��.��P'a���*0��ޱ�<����j3���k����Fw�̂���P�>~�{�蹭u��5��P��i]�nnO1OJ��  ������1�䡵��b�1o=�s ;����FU:��c:�1��[�\\;�\3P����p�Yj�f�1^�9_ʛBa���Ɖ��V�[�݁���it�T+��E�}_���}D�Q�^���c�8�a
C��i7E�0D{�0t�I��e���ϟj;!�?|�T��� <\�d{�*G5d��dDVi�̼(n���/I�L7������šP|.�t�M"��:1�A�S��.�1����U碉������6&�xٗ���]��WT��y���ܙ�~���{�߅�NS�ǖ1G�Nت��l���A?�x����s6v�]�Ϗ��?��������߸����B��jf�0Nn���>�&��ж�s F f���K�͡���7�M�!��6o&�}®r�������2F޻��h�Xg�����=��߹0
�%1 �Q�tu�]p�����^b��)�S��Ŏ{�{�ߣ���u~�> Z�` 	l��s�X�ѣvl`�:��dH*�y���@�}Q�<@Um,�����)
�D�m��_��8��
�ʋx�s;&@�?b�f�`��u6#�3�Z%U��`>�js�|��� ��᪳o0 �����XjgO���<NN���=_�i��Ga�X6��<U4kND.[k� ���3�����P�&Gxc_���M>�IvMW��8\7��v�͂�[��&t��)J'�F�l�Z���@V���賎��Ti�%���If�|k��W��K���ڞ<B�N�"��q�:^���n0knޑ�#��z�:ʁ��Nd�
�>xkA�RM��p��uj�*J�L�)�X�ڔB��	�`�7�lm(�8)ny�~|��$n<M���$�e�bx�:"R�4����x׉2i��'�>����tC�9�W*?�@5ȑ�R_n[��~<���S
���=��6̤o��|�k�3)���`�xV6�0�@�dY[�SrO�E��x�!@�`���1�z]\j��CgR�� ���>|*�MK��iê�M�׹�}����Wt���v �҆���B�NoM�ț^H���0H�t45�P;O@�Q�k]kty�b nV�P�tZ�O���D7ߺ�o�x'oH͇?~��7��H$H�4mv"�0فK��xN����y�Wtm'���Z/n2���)�f�pGc�p�z-�1�]��?s�8��\؍:H��S��K*3e�₽a�s�V��K�gͽ4m��G��ʒJ�uĿ.|`���_[a�ΰ�mi��xO�0�Ϣ�i&�sRyr,�bz�_5��]�aD�R��'�	Fdvn-I��n��.L�ȤL6��M���z���Sa���d���()�^���+� �gJ _�L錧��<?�'y�e��zҭ��� �Xd��^fH��q���F��<�5�phm_[��%�B�|oj�b嵈U�2�nD�/S�&�?,�E�M��g`+α?�����<b��D*�׈gCצuE{�������ҹ_e_P�)̢^_r0PJҥ�b�rWo3�p%f�
 ]@&Ly�����]���i?4(Oe��>�i�d�	^\��<kͤl��[�m%CSXj�i%QG�.��G�swJ�Nj��Do�Q�.KRd^Q3��u8�`�7)o2�W7�<M��ګ)�,&��3La��������#v���s\���ܘUE~���ן}\��0��.x+�V��iG� +�
�?K��d���-S#�����7�n|4�����9�y�^�˲�ۉY?�A%޸�Gۉx�y��
w?��D���ȃ�������Xwӹ��,�1[�.Uk���?�C"���FXt[v�U���H#�}�$֑C*"FY#׸�\��1��2���O*�B朗��I���@�x6ի��訨����w�8't)s��P�F��h��}-˻�6~��h��j���r��P�4e��~�j�f,�"d�b�qO�U���������*Q��(�GW�ي̔���:�/�O��8�25#���ft��[�|K���ٓ3�C�l\�R��P��:|*!�T5ϸ�U���-���ouED��"�� ٔ��-�QD9m�u�DffqmB�m]q}��Y���T�b�j���1���>��e0�oխ���,���I"[���ܘp X�Ut�<�@���xr �Q�����LHa��	�/V魭��]���Mi琙��I�[6{MS%A���|r����w�(yP���lSߧ�o��sA)�k+*2�>gCu�w����ZU��8�b<>���
����}��;s������Ϣ}��&٘� Z?c�}��*��Ul~�;��*�s���7�c���^���=*ؔ����G
�7Q5q�tc=�u��k�0A&n����U�ԇ�!�}�W��{@w�Wb�7�S��U��?c�1߈�Α��/s����F.�^$��N�gv>��/��%��� l3�hʠ����E���ԝu�O�����0���A��\ˤ����N����s�l/�ׂ�p�_�*��>�BW��W/�D�6�҈��6⾛���y�Bۥ�'Q�,s�7
T�R	�}��Z���0����Q�T��?FR���1�9�j,A#u@��؈��x+o5�>W���R�k�C��y\[�p.����mn�����ZÍY:dD�$�����pĻ�b\p:��k�.��za6�7�9)��@����/���j����,�&b|!�x}��X4l�4��űX�0� B��/��"t�]A����@������Q�i;șD�����������F���-��>�u�ƘGﬀU���x�խOD)4`T�ǀٝ9��Q:nT��=P�h�M���SZ��s'KSu�n��]�@X��\w��R0��b �K��}�{������*z���02J^��VO�(g���~�F����y_%�����X�`sSN6���by�$��{��v��O�k`d�[i�[�5�^*��*�>�	����*7m����8ʩ�/~/!���_8�@�Gpl�e*Bl1��C�pi�C��÷�Bh6lz�P, a.3������H6S�s]�V6\�����E^�����xⱓ�'��R�yg���T��뒡���n�y�ڱ��e�����R	���Y m%��9���4���Ť1	eF1�����Z���ލ�o:߿t�F�ITu&���Ozb�i���Y`D�TBŻ_ �ʍ���{�is�׀�hhLNy�3XB�&���ŞU�C���-��4�|���ӎ�C���)vύ{�2X���5�3�s����툀�C���y����k5�o�2[��f��� D���@(Y�Y�%����`UӪ�4�f�Jg�b�
_q]�>�ø�w`ft=С�y Ȅ)�Mm��<%o���ʐgA6��������ەU��cj��:K.N>�IJ�u)�2]�k�~i8��ȑ�ow? ��7$�v7�".��s< n,}(�����A�_�DWs�=�.��^��k��D7����Ρk��*Y�����*���y��Or���X�`f8���*��gv!n Cһ쬈��k�vT�9�H�4p��#;�·�zL`v�]�ز�ʉ<����!�O�}w���<��GOgP�b��S�u��F��i���3��m(2\�}���7a51�p(�����z3�o�}������H��l׋:���گԌ�<X�"u��p؎��_�����w�[ '*��Qγ)�ԁ�ߋ��ː�
5n�ٻ9�ck�$q�X�< \ ��{�"`M�X���������A�=.�XG���`��q�8��Q�
֥�*ϡ�!�1��*h58�#���.�˭�3�b��I%֩�ec8�]D�͟��t�;y7Q�SGDZ1�P�$�{z�e�)�	�~|:!�����.��i�&}��%#�h�v����x��e���k�^T�/��tyW�a��� p{/��cn@��7�.Fcm����j|.�AV)/qIP������aO����e����]�������Q�g���g❞nHuI r�Bu>~�L���o-| ���KF�D^��Rm,P�U7'��i@Y���Y=���C�|`#t��Pqת��T�_��w��V�O���R1�0� V+����hLi)�@Q����<Hh�TJB��1�|�6�7��gp�)��$q���E삵>�$6p����\{34��:�NNB;��4�*�:���1Kw�>��Z!$���2on$Ӧ2P��1���`��:�j�%�w[ӝn-(��P��p�2��!�;���`�1.�Eҩ~�Q��_�z@�,/Y�����+�!��m@&�u8
?�??9��U(�{i�|Jr��>�Tp�����,�5R�F��20+��B�B;o�e��~3ix!�}]�L|}'��j����86ə�N1ˡ��SA�8�6�h�|Dט3�r�)�F�L����?�Y��M�^i=��B�W��e�0�����LP���h`�� N���2�{�y��5�5��0�]��m��+���:g���U����h�[<��#sm�n����D��|�p���t���,��y����[�xM��`�-~(�����h<�m=^�$p/	A�}�K鯯�5��t�#�x�7�Ļi��|'�bT�U��76D�ͷ��"���g�YU�cCQ,u�G�N��?�\�D�zdw�5.m�L�����b�5���p%����M������~�	?� ��m�ݸ*f�g9�v'���&����I��ң;��|_�[����]�ה�(0r�G���]^C�`�(If��\��d��R�t�t��*�-�|^oVD;�^�D�|2������"M�)�)5[�58���b��|7�6v��ɡ�[�^�sn~Ў����Ev[��hɚ�O'��?Sh
�V3�1�$�Z,:А�X�3Q���)a�{�ք.�4�>K���ġ����]s��1�E�"B�3;�OTk�K/�u�����X�VuJd�?U������sq�����Vu���Q�zzd���F�'���B-jQn>r����-�b
���Dņ��E2H,�������h�$��ǌZ~s�����,Qf�!�o�\�	����\��`�(��tڨ��,e��X�c�`D�d�E<&��W��Q���[�j�ױ��W,�-=���V
�Y*��)C���?��$;��E�P��,��m�5�{��r�����TO�R�0�oB��g���?�^m�7_ˆ��|�bp�+���ۓ<I;*�
 �t5�5�4�Uf�vҳ�l��\���(�9�K	��;�U�ˀ�����W��K#;	����"���ǲ�y�j���:� �CM�-�0�i	�y:})�o�n��'�I.�Z~��٩2�y!9��6G�ǒR����8I��A����^Q�՘6A��n���>�A�x傂W�@:qH>��Jzܾu���QV5�!=l��k <s�O止���ϓ��f��lb�|!
&�Q"�(��i��ۦc��U	}�"Ք-B�k]0<�!U���tm��Z7�A�n.�`���B^QL���=>�o��[�2"i�����̘�Ľ#��C$-Q��ġL%��%�}rH�؝V�Ƭ��~w }v��/rV�w_�z��M�����ț�����1��'���_s��R�V݀�m���q�s���ِ�E�������/�XQ��T�����n!L�۵����C�v9��S�~�R����fh�\�Y�� ɓ�-��ۅU>z ���_�Y�t8�c��R��Ωڸ���*��ۚ�^d@Ȝv�JԠ��M������؂��6 �<�Z�"��"Ǧ������)���d}��9=�і;4����|sɕ�f�a�F�k�
�����&(��G��Q_M��J�BG���gbHT�a�y� ��l�n>ږr���~�f��B7�́E)�¾�Zh��~5�H�h����%���bj�( ��*r�K�{+�Eq@�JZ��]�f�	e�m��|U�F.
��Eƽc����f�$$j�IQEA@��ޚ�ٽ�R�ߝ@�"m觲�G*��EF5\mY��C��zzm��gX�K���v#*u�������r����U�my�b�g���M�=�B�Ա�C˧���&�X�-�����Δ�+�A��x�Y����J�7�4��y��y"Q�ޏJ������
��t���m��l��I�:��R�N
��6C/3/���� ����ܞ<�^_��m7�oȴ�йف����,O�U��AՕ{C�<�u��S�wA܇Y6�]��wL�G��j�/�d'�����[������*w��L��a$Xh��]W���
o*���SS���י��Ϲ(0�d�\�Rt��q #�{T�GN�����A�/W,<����%ߊ>���m�x-�(�h6�(}�#?mL�6$ *��=��O	@Ʋ]�&^�'���:S�6�<�mi%��c�ӡ��c�\��Z�ːc5���ȸ�q�A3;�n�</+�J!�ɊC�ޓt��d�r��dJ��+ �Ĳ_j�!h�s��L0�)~� MR�d'J��_C�I��۽�Oy��.�74�D
��C����D��&�yc�V�Fvqjc���'�ʤ�K���.����.�k����ufW�JՏ Xv	4�p�%�c�4}JN �w�B$�F�">M��{d�߲�@��r�T	��qмk��E�W�����EvBI�m����	Kuqd<G��,��heX1|����gN��3cYM���~��A��#�o��O�Ǵ�m��!\n�l(�׀)�2�9�������s��e�TŨ��3df�M�$Ă����?��!�ܟS^k�2L�d�/B����xs2UJ)M��㾜��\�i�/����ϙ��jX ���+(��%��~:�vFh��\��/�>!פ�ޖ:Δ�j����[ ?���9��O�b�=H���-�̇��Q1�����A��W�S��FƼR�e���s +I�/8R^T]o�?-��5�����o��Cp�����]��"9&Z>W�yi����/�I�b�~�b�n;q���O~�S%F�Qx)	�ve��*��yp����`����������}����¹�Ū�z�<�!�AS���"��F^٣�� �/�������~�&�t,�X5^ze����xB].aE|�SQ�����3��ع@��6�oa�v�sG�n-��؟J�8��0���(����~�3����L�*A!�wb'9���y+���~R?�	���F�P�Jejy$�U�l&=I,�B�(��m4���s�a���c���!�O����2
TO����:���5�͸�&ޭw~XF�et�M����#�/�*^&+�2�m�WE���%'D�o�Q�=��2^��~�%B���ה���f�`�~��kk��s�{C��r�@���*ڵI������!u��	�a-�� ��%�e(��5�F�¨���g�kT�M��00�۫��c����㸻h�����Pt�����1
�v�T΋k�&�Xu�=����s0ټ�\��qD���h��S�N�29��} �j�ð(�e*����9s �5?�&�]m�)�(�)W�/I� ���E�������H�_^5I�3<w�h�nߕ���M?��n�З�J��L�h�κQx�ѧ7&���S"�Y�]��r����0J�c?�#��/c=?�6�#����ɴⰮ����� �au,�Q�E4��=���+�׮�G�J$Ǫ��A��e��˃`/���XBB����>
/�5R�R�s���y[��<π,�K��5=�����v�F�$����c�60���+��N�-3E��BQ�/����L9���7� �{���y����#ɳ'�\h�m��^t��������*��Xv���l���/�D�2�����rV��*8�k�R4;��׎{�8}PbM���JO�ȧp��>�\�\��^��G0��AK ��F�Ï��͂�I�9�8��{��c�@�}�U��_n�|`�8|����D�o�2\��� ����d׬�`ܜNMpe��Q�";?��ʍ�N�d��`*�Ȧ�M|Σ|�6� �f$c�Wf���hr�o���0�
>��F	F��,�tDDftԏ��xj����fqGwdD�ҍj��$���I>mV�Ya���3L�	���SJ�tDZ������B������c�k��L��󦺋�	S�+�F CpĶv�HFܒ��s�	Wa�;7�bB�I�4�U�1�F����
[q����ئ�M{��Ҁ��e��ڃT�"^�ߌ*�	�����]}��Qt���(�t�a"�6qA�h��?0�m��:k�/�u�������X���������gY ��$�q�J$!�KJ�-��|:�E9�j[-���kE��B��HAP�/�0b�S�Η�ˏ&e�8���8.�WKVn,m�v��P�C��O�oa���뢠K>�^���+Eޒ|�v0b>'Ǥ9/\2{��?������q�=��S���Ceܨ,�2H�_���$`���;����T/�����`J�glLvqv��[D�t��)t��C0����Y�pd��)�_Z#�C@,�����;P*�
�$f}����( o���f��ٱ�BR�n�;�E�E�M%k��:[�X1(�����},��%��!^�L/�6��s���&(�󩴛�i�Dg��0�:�'%��r��X5�%�	 q��̓˝w��W�-g,�9ñ������Ye5�AqۗZ�l�Zv��en3�},�)�Y喇騻�"�]�K
2�:�����	��鷵�����b������s+��$�OJ�$r�^��P�kG[���h���L*?\��Sו� ����U�,C�m.�\2�	|�w���=ceH/o�>��nO:/�'�١�}���ۂ=�$3�x�A�\*k�؄P�-m>	� bl��4�xe#�z�$:{���5�������Dxfyk"|w�D׶�I�MW!�bRW`��E��J(�\�]=�G͊�z�U%Ek�X����&of_р�k� ��/M�st߅��[����u����QzqA��ti���ќ��Lk��4���������e��|W)��ݪ*���h}k�s�a�x4����]~�s_�W��Knf�1�7�팯|�꺼��.J�Yf�ɆΎ�z��Z��@�Y���]`� 
�ړ�JPs�i�͌�STE�Mx�:���%h�(�K}���0��-B~2��<���2�+IU���M��*�ݗ)�>�i+��x��h��lT�q�nk]j~e��[?�����RZW}y��F��{5|�ۭuP���t5-�X�&!"JMWl����d]us�nj~�؇D�myOH�~)�#�t��s)v�֠�����Ƨ��ܰڔ ��SG���l���U��A����|@���G;m`�S���[���̃ʝΩ��1����,;�L���4a��oyύ��έ_yt���-�Xҟo���Ӽ��/�tI��s߱ic�m�!VZ7gz�<ړ������u�5
�E�;-�<���_0-�ԧxG:^fΙC�J�
k�iȼU?�N�`�_3����ٛ�FR�^)��(���(�_�����f�V��`�8g�i|���f.�����׌"z�P&���������71���p�a¹&
яu��j��c�L��^.�\R�=��x��D��y��KG�nt�;�1M��7�h_�>�NP�+d{HL��'����Q�����7�~��'[R��C�`C~�#twՇ�������_{�Z�Q�e����=�sU�U�.��Co����Z�J�/�!Ů,M� �� <�Z%� ��Z�2k�Jt����rR�u�(?UHi��CJB��\�3g���.�ї8��9��L �Z!�t�q� �$�hR=a��+��hI���W������4��Y��H�����d6����w�+CS~���������9*`YwMt4�;��������­���sΨ�]vR��$x
�0�����z�!��<�߄��s�#Fo��}:�Ybq�مL�9� �rCU��u�F\4�"��ާ��5��/��1$`��.���^&�4�=y`��GgQ��Z�dײ��������B:=_�ic�ܤc��hx?��3�0=����b��h�C�����_���!�����}�̄Ł����pe&�k�keSw���8��w�2c�����V5�xw�LXN�!��e0���:�"�^7�S��U��}�ê�
5De���{(l��)��=o��!�;J*5��Z��M���������F���U9R|�����5{X-�m�G�t�E��� Jwf�ܥ��qB#zi 1*"��F����" �O]�������Ds�\�xM��yݧD�NE���X����\���7���\B/]Ud��cM�}��p��p��X��v������01����c_^Ab���Lk��h�Vug[����LJ�B�����p��v���F�����d{l܍u���BԲA�2�y��yM[S�x�|%�D?�Q���
%�G�(��'Ш?�u�b�7US��vL�0rC��z'�?�f�Ћ��0�1f=��./q餾���"�7{�C*/!7��{���h��q[�I�b�Ee{�U����Rh:Y�+]�oHx2������־������Cf��8c�a�"E-���K<�Y�}��MI$ʾu�	�4j9}���^�Ki6�!���eA�=���[2�>��Yr�Ƚ���k*�87�澫/ߣ�_��fα�֔>�u��0��U�����b�-�+�}���M{��wsq�0ӐGdȋ�R<}���ﲚG���A�\��� �W;RܲG^t��}�皤�q�ǚ�51d.Cqǘ�!��9J!����8��l����84D�6�w���G0w(��n�<��B~�Ӆ� ��{N�����D�%������+��ˉ�vHE!u��B�����}�C)��Cz�SSM��Zԍ=����H��[H�XN��ϫL�R|�}֪�Wz�n�����3�
�鏆{��VvY^���(԰�,�Y�{Ӭ���]g�%W
��#FnC�{OF��
����a�H*�-��[u�������jǟ�w_��a_�,d*1��v4|GZQ�\,1CU%��zlE�Ƭt�+�/�'(�G�t���!�l�t�$�h6���"�3 9��G<2��}Gu�Ӭ���K��H���7ݒ������C.zx�
����H�Ė��]�n�+n���Q�_�����r�s�n�(� �;�ħ�V��N�)b���Է�����&u�X�4��*$�o"��g���8�ƣ�We��V�):J���OF�n"}��&����t�dޱt�^��%*\�Q=9����N:,iY�j[$�yAk�{�\��GDv�Z������36�0"��A�1�6E`�J��q}���c�sP��i{����� ԏ�,��H�여����Dgr&!#l$�ěp�?���Y�gR�� |��� 4߫ȿIӽ��`�\�jۭR�[E�P�k�,�햻7��?�{~�a3C��N[wYbK�^����SV�ol��>ɱTqO�~Y�[z ]B-� �f���8F	sB��p�D͡��>ݱ�z�Q3�����<���B,�6�|/ �\+t�x�2���M&`�E�5�?G�qF����aE���|�U��hK�~���Y�MI�M$j��1j%���>eՒ��O�D��a$rOK����JɆO#N(<y�~J��x	��QuԎ)I��ע�>��A����t���YeD�>8�M�@?�qE���':�Xn���g'�V�����,��k+;��i{��A/��Yk�`��QD
�᭳�����2t�Ҟr�4��C�aJ��ˊ��LJ��4��F�/�XrK��fIF�L[�7��w�(��pzh��^f>U�uRŝ��Nml�w�h���V�+��^W��2$4��()�e�DE(UzMjñ��+)��с�WQǇ�j�Ӝq2����L[mcʼ����GP�i"��
����H�W�ۊ
"�*D�qÕ��R�o�t�$ݓ���j>�s�a�i��~Sm��K@�Z�)[�FAu�7�h$��Y�Ό��,O
'��� "%�#�i.�SiK^F�e�bd�=(�3�=Ph��<ʧ.)ߧ��2��{�~uF���It�S����&�P����yZ�eV:<R�v��b���ʾ�=	���82�R��\fj�O�����<}��?n���4ץ��\�#L_�C��}���R_��@j�G�Ɠ�k����+nP���!doe����~����i+"�9$V�3���O?��O�)���>K�r(�M�Ʋ�{Ļ�9� �Δ0�@9n�:���_&�+/�g��� �7��t2ZϘH�4��r�i��vc�J��q�B�68A��������ֽ�"��iT(�����T³*6 ����D`y%~J�v���?:���` 7�^�4�_Xf:mSĤ=�ڕq���(*�I:H_ ��Qg7�$���	�#�BE�ؗ�\�����U;q�wmF�Ĭr�x�Mr�ڌ�R�����{�q};�>��J�k��R�.paQ'<q3�q�]C�³��w�p'O�pH�]�W��ve(�Pw��Cg���R->Ř�'Û%H���b��J�Tݠp�����.f�kοdu�õc�Y��(��B)` ������L��C�zc�o�ʋy��ǭ�����E�x��P�I��B�$�
�jJ�����Z�|�����c� /��?e}��?�-xlN2������8�ú�)�Z4F�ٟ����	��x�P�UD��%�>�Ӎ��C���Ny��~_��դ�Y~��	���3�dU)yt�5Uo���+
Od�?|���K��B\�e�����D�¹j��7��F}e�Xp�u���!����"�����\�x"���0a(�nԑDw�[��8<�E����;.ڮQ �gB�Yf����5&o�f�ݷe���n9typﳧ.�I�#���щ�F�=��K\���2s���$�u�F=��N����A�!��J�����g����kB��d�d_�z&��Z�%v��N��'v�z	�ӳ+bF��2DK�y���	�?��`qL��5��.v�l�Q}S��*�je����k���D4A�֣mo�A�t�Ws��kU�;���#ag:8����z�A�,�W1���")��9�]K~���|c�x�L�vQ~��]˥��晖Py$���/��=��3?po�\�G��AS����x1<�����By&���N"BƑ�F���(�� ���sO �.M& ^��G,NS���2o�2��p��xb�����4%�K�p�{]?9i,�B���5f ��Ry�FY$��+NW�B��5�)wx�gB�읉�e`E���>v0T�r�.%ɼ6�I��f�����o�L�L۷�m�w|c\:�X/��]0E���"�Hة�L�t��E$)�8<T�f3{�����.�\4&���&6p�6)-�kB)-�[#�X���h �i|~�e�(���$����4�ZZEfpn�4�k@.=��jJ{^�X�h%�*�����_�"o��x�@�I�����QC%��.�����6��ҳ��'z�}D]��9
Q� $�n�x��@ڏ�۬��.�+��4'��H�s��d���Z�	(R�����F2���w�v��)��id -VM�y�㷰�%v)Z��'Cu����!#P=gĮ	|I4�Ȼ"'s�� ���aJ%g��uy�Y�t�Y�|!�A;�:�"EŨ_�\=�q&��3���/��m��V?��%�%��b?_���)�u~�X�Ӊ�:��VnBw�=;%� ��������LLFo�%[��������f�>G2VX�@ժ�$�m��GǙ⌕3[6�Awߦ��x��+tĈ� �#4�Y7��K&��
%����PMIDi��K�zf<Y,��Y�dZ�m Gv3��x4X��Q Fy�M�[����d:$+�#�tr4������aL�$��<�G/\Ŷ�s�o �!8Q�H�"�4�2���S�tx��R�Z�Z�+PP��@`�X$����\+�5+���N��4��#1
_���D�˗��	�Ø���X �}?tk=��sV#�]�%q9�-�����F�tD���TNM%H�fX��0C��N��(�9:(dd&MH,����-��4/r��o��x+�!0g�>��݇��,f�vDD0j���C������𱏇o�����j%�舼�{ƒ�Ʉ�8 Ju�F�/��f�T� /�V/� �X�&��,���X{�i�SF�A��3���8�L��\�S��RF(~MX�C�9=���(A(.N��3��yb�dl|yBG	�6J�o�'�Le�߾�^�K[#?�V�y�W��R��>L�$���J��TÈzm���s7���ㅖ��V��r�}�0c���.5�2R$��a�_w��<9�V,�M��p9
���5y��Z��\�tk�ԟ��t��"�AL�{��LM�T�������A\�\v���s�l��|8HO�E )�o/��{�ޓ}�zq³e/�K�EӤ=>�1�H#��򍟟	]}��$��6e�r����oF��D(�piо:�vc����'ѕAdB�pڧ��G��`G����d4r���5��;���}��%7{��]�Q�O�Y���s����Ƥ�@�<3yohS=s���RV�OC�6�� ���Y��z�^�0n����VECQ�1������-�󵰦������A���$�xZ��~B�ʁW����:29kt�spڴay�)�_{���|��T�s�[U�רg�e���}��^�|>��c��h�z��Ib���m
�����Ϳ<��^sG,mvU&�E�:���^���+��6 �0{,�ɏR;/r�P*�,·
�ĥ��9�S@Ђ��Q5�RX�������Z�;̛#����ZcFu�М��n��\J>%���I�7�B��P�������fgW�JAߖ��y4�z�%���u��np�����aP1�`7X`L��Ҳ��χ�v���m��]����
I8ϲ �k�R�k�U)�rCZ"���<��Uj��x+���fM&� �'���֐(���[.��<�;��c���3�e��r[G"=PP?馮��yǄ�7�י �G���e|�c�|��#t�h̢�~-QN�Dn��í"�X#`���˨Ӊgj}�H��{� lD����(G{�F��V�����;v��E�7jYX�q$j�n/���x�Ҝ�v�'�4ԡGOV��Rפ�Q_��Fkׁ�&ߴ�ec49b�ߨ ���vG%��0���z}�Ŀ�W����OAa������/����/�rPm,�v�:������_�T���ll��\]͡cD$��5~����J�����*�Oa$�L������s_��E+'D:M�=�B���y'n�����ht�QG�nlpXA�i��XzJ*�&��3xf)g6�"c���xb��<��[r3U���:$K�=�ż��[ɀ��ox�6>�O��?1_g���fy{F�LK�bf�FGaa��h�&?��MO�~�Ԋ	Np�c`�A�A��)�"|�IC=;:�
'_Γ�܏U�������
�"��ಬ ��4SxAb�=�I��aKC-D��;��Ӎ���Ąn��`Кy<�	�͑[ 4"^���]hίm�� yz���$�ҹ��z����%(Q�����aY��D��6*)��ᆩE�$Ut����A�]��Qw�D�ɷ$��8i'���Q �e� �e6_�mƍh�-Ѷ*�D o��e1����b�� ��y�f4L��7��ZX,���+�)y��سsj��3K����I-��M�ъ�D�s3q]�<9��%��ķ�'6�z��c&z*��
RT�/���&�n���^�C�m|z*���q�i����>.�$��7��̨J�no՘�W՗1#)��V���9�LS�t�+u�ؗ�p�:섥��z��_�N��]N7���][)�9�{mx�Z! �$��:8w�*�z���n7
��Ճ�Ϩ�^�@?�I��o�7AIo(��k���&�X��}F�'���&�%g:q��h&n�-γ$c���4�����e���a����xƷ����T*_�V������J�ϣ�c�هq�Xj
Y�<|۴��,%l�����Z�Z�2�}��쒊C�n��y+�S��!��mğ�k�7x�qM�EZ�@�����5K�6o"p�	 ��<��
����URVϑkF�WXs�e�ǖ�am�+�S+eˍĢ>@���#]�C��j����W�%m@�h�\�@6�F�_t���p]H��Ύ
���������W��o��;c�	Ղ)V���j]'z���f������PtdEan&6���/*w��J��Q��6jZ�@���
��CK���u�\\I,���c�+<��ݐ��|2��ؐ��;��7�������%��%B�4pocB��[N�syDb�^DSYXң�{���IB_X�ɝ�|�bs�,]J���ӍNݡ�t�:�«��. �~��r�"��$��a�����0�Yv���B�=�j�6mr�[�{��L~���U�#�(#��o|�t�0��B�=�2�u��:�pX�`Ғ*�*��Ɍ��le���i�	j�����R�'#��C]w�8���!S�A�kX Cm9c��I�d��T��4�c�XSI�ԩT�C��������9}g��=B��n3����f��{KDd)��qv�s�R���$
w\�o�=�*��Za����)S�+��b��r�)W���R5�Z�7(_BI�q���9��<���W�?-�@���J?��	�gL�/��;��
�+�/oҺF�1>�!VM4�F����0��1���@WĖ������a\�?)���K��QV�t0/d�qk�[�=���`���A碠2�U�%l)F�8�(�R7�h&f�ۘ>�V� s�M�I�m)�z��&HfW�/C�2ـ��v�6�"*UдD[�%�
:1h��Y�t>.J.,ղ�7�ch��<2M�����A�I�0�ͩ���47�:��ݠgO��ذ��S�֨د3��djЌ��>]A˿�5��w
9!O{P�`�s�F\h�p�AG�t��|=;�E�]��յ�/;�t�HI�_�dn���0�W3����=+EeW�lQx�24���ZL�J���k��R��V���;���>�"�^� ����V�m;v(�!�9N�Y�J%�f���+�f�D��nz�� ��r�t]0�r7Y+�0��j��J;��hq�g���_Q���%);��8T���Y��b� Cߵ
����xiBE_�����/\_3��-�l�r�@��`����n 2����N{y��2ղ����p�
����eR��M(��ľ�|�M�G���@�������=I����i�,F6�9�h���QO������b��'��C:�l�)[��H�m���� ?y��%��H��������������)�De p�:qnʎ�)���x����_�7i���Yw/�xW��(��"푹j�=j&�\ Lz[�Z�k�ʯI�������!'���r�AHǝ3�u�����*��>ZԸ�(,6�@QCMH1m�H*ްt1e1a7����z(:@�αDV>e�Ъ�$���;��A�U`�m� A3O�y�:��,���}Ha��������5ˡ:n��V	��X4�u��X�k
��[��(�4�^қ'Q�/"(�i�t&�� �;��%���bk�]m��8ˡ{|�^�sԏ�%�1�Z�s[�Q�[�Q��r��,-�t��l�5W�$���}�^qz7�^��Gn�	�-�0���"*�����WuϷ"�[�\��$/H�%n�J1��ai����w
F��L0�8�D��h̟oo��ѾG�
-��g��egF�dŕ�o�ϴ�[;kT��U󙧷�/�Mr�p�ѳ��WTq�����6>G'�&QR��Q��Vo��K��������<Q��Br�I��/�^�4H`ů�������F��SJ�G��9ǭ�|Z�B�k�2kH���I����$.�̞nǕmyJ�����8�O�Db�cX�ȧh�u�؆��� 0��SM������;ֳR��7���g���"N$�g��c��hܚMMK���Iy���l-~PR�o6�ƽ���0N<�c��A��
h�q^,��M�0��_�`j��� !�aƕ$�d#�~��{���XC?�ͨO�-dA~�X!E$�U6�W�`�z����Q�-`N�e��9=�t�g}��#h�B��H\eʐ%��fc؀�4xL	��>�]�_�ua�F̩�x�=�n;
A��18���'�wi��m��v�rk���0|�j�Y�5`d��y��[��77��X������^���6P�(|�D< 8�Ac�.?*�� ]�(��*)�B`k���s�6F�W��QJsƎc-J��eG��2-(�կ��`��z}u��Zư>�%�e��rq�,(�A���~�~2�`��0F*�L��4�-i.�H!��M�ћ�"r@����4F�[�
-0;k�*sД ���?l�n4�F���q��2CK���\=9�q��εj`E���hhB�����l���ʼ�|�����H���~ �X����&*ܗ��㭜��:ةd&����]�]�R����y�Y��� ���nv&��E�;�H]˲]֗�_l`�5a�8�0�o�?�F>S�"(�E�~zU�5��l+e(��k`�J�ߜQ�٥�>wq��.�ض��K�=�c���GqO�����g$�:�PU����AIm�0	�>mr�k�*���lGGu1t�i���f(��|���!8��2d%�ڥ���+Uf|��5�I�P��V��R|��-�w��/���C��gC��XJ	��&NH����T�F-L}��J(����RJAbB�gZ��DL�j��_1��
�Z�Rֹb�Y��\1;�^�`��I��)�}ܤ0���G���/�(�D���S��vy���U�|p����t�5]�c�?���̄�d�x_���#�ە�P7m��faB��;�"���[�7���a���w˂�f�د͝�`*c���_cq�H�.R	���T�hU��u��2�G3�xј��l�$.�+�6��c�k֟��@�6�fY'w�"fؓ��~^�6Q�3�s��D�D�Q���
Lͺ�Ub�3C�!���n�EEND@����\(���D�J�F��v��<��zΎmURQ�0[��7��_��q8���ҿ��L�1)Q�  �uց8xK^���H���H��l�&�]D����)��ӯ̒�Qs�n�l�h�b�cG�/�))Kc���myLQ�Z�Y�9^���T�����Ը���Q�1$u��k�.�S���Dۭ�-zd}��$�����Ž/ �n�L���.{�L� �i ���h�c��Nv���w���x��-uɕ���g�\5zPr<����E�9��/�o�E�����Ċ�*�ӻ� ����|��A@�"��U�L�P�EB��!�K��X�v1��
y�m(]B��pA=��i$�ai��c��
�sX��]�_�� `��je��Z<��?b��CQ��(����2�=|��B�ְ��u� �d5%�L�7�j��}Y�r�ى�.�����?���C����^��6�ޜ���N���@R-j}����
���K�E�`:�8�����8C��3?C�"�"�	X����!���!��.5��:g�z����HbԅvF�P��L!���N	��q��jM'8>�~�W�r0�	R����4�����w�A��t�^���_Ba���F�,	w�az/�� �[��:쪘ܲ�
î�i�`���F]�nS%+!��,֊;��';ca����]���3�o� �0��t�-2w�#��H75.E{��;h0���/�.{�݋z���|���p����y5[ G;�;���-�D��*�>����?[�'MY�v]�p���-�jg��G�:gR�	�p�_��Ů�䲜W]�YZBw/g����<l���*-q��N�DZ�pX�c�&!�Z��rz�B)�F�S�8���/7݋�Ĭpn�;}�ۙ��Z�1,�[��p�-ғ�U��� -���"Ю������Rne M,�t�JHaS.�K�$����2a����)� �~x� 9�> }ĖwM�b=���m4���2{	� �
s޵��i4����D���<�L�D�I��0�[�l�"F��d��o���
%K�\�]��[�����hp���-�b7T��Hq��Nyԁ������=ӢX�%�1Ӻ�m��c[w<k%C^$�1a�	����	acm����u���s�M�n,12��h�v��]��Nq�o`\�P8��i��K�����	�o�R�[r������2CLw��A0��l8%i����Z���~�l�ؘ�O���	�i��X�Y��li�#�s�o��~�G4�C��|�w���PlB�E���\s�~Ҙ��t�Ѿ��?�8������/��&�	M*�,b[�$��4sT-3������!�Cd1���jȭ�!�m� ��.��;|�`�Ǚ+�z}B��f;�%�=�u����'�c��Z���Mh�u�N�!FJ0"��Ȯ����b5�}n��$�H�]��%+7��<M�FD�������6D�~����@u�u��e�/'�5P^+��{%B�S�|%�1M��eo�C�_�j����ӪQ{�
b/����:�����w�;"��h�#�#S��t-.��Y��}Mm0f��z3k�d��S��b��E֒�Q~dޙ��1����O���L��Z� Kc����_���c6*��ip�W�Ŗ:uJsf�m{�Bl�N��m����`�n�ۚE���h�Q���[.[!�#����_�u#�gٿb_�d�]s�?���4�e|��1t&�A����[�;v>X��ͧ���Ǭ�Sɾ��[�� �:������a��S��5�wlE� �:6��D^��m�Y�)-��O�T�È��>T�Cyd��d���ܽ4Xz8uܶj֟u�6;.����r�J��:]�B!P�������a_NU�<�~��1���
�I���A������Bx�j�t�{����IXQ#�0[E���x�6 ��ۘ%w���V��+��ǩTzV�����e�կ��s�X�'��8h�R��
j����b_}H4��e��7{���(��jQ�"!�C�4� P�-�]K��H���a!C�b�x��@r���m�\b�BP����a-��Jg=�Z��ҙ�6H�m�#4⛝A���`z�N��4@��_�T6��5�m�10�۝�?�4%���KO&#y�q���ڦj�K��^�a-�

�2:	��^���실X�p�\�C7}:��kav<�RCm�aC�C��p�78��	�K:f���3�1o�uU� ��o99�-��2�(��H;�uZ<Shyp��<��6��g������qlۆM4���	�����Y����:���'�U<�S;F76'���RW��x)T��5�"��DԞʭPU�Za	�WZ�GW��bzV����nOpN-'I{�w�H�3��Ί�:�3`�ɨ�����?4`(��j��H�,{�
p�M��:��9+z�<U�1!�4�����pg�[mn�c����q��06�ϥ����I�[U{���We�u��и�Q�6Ռ&r5vی�m1gT�^��^Y(T��d��~&�i�3B��f�<C��o��9,�@�Y��g����Ne�� ����[�:p���路��^j�lQ���G�TP��"䕗1M)әF�+QEa����(`�	���ܸ��^����_���kQH���� g�~� ���!�K_!��ܺ��wߧ�%t���̬�r� ��x5��h��#����b����������l��
���0	9m�#�w�w�n1�'ĽE����=v���}���:l���Pˁ�ͥ�
k��Sw�;��̅D6��nn=��]d�cٔ��j�/km-��J@��|��Z�Z����"p��3$'R�2���Fޫ�{%yMn\�û��W�'V��� ����ޖn`�`�&i���/���$��y]�S�t�ڤ�>�?��������t����kj6\�i;E�,�X��6�jz��0`\A���>ӒC1)g?`�ݍ�
�9�A�F�c���j�e��p�3U�������!D�gm��k	I�:�\F����! �59�D�I�8�ȯ�� �����̓��I@[����p1�����-0�4�H	G��@S��T�~��]�G]MMhҡ��^�m�8�*`.o~����HV��G�Z���%�����z��x`騪�eY�yZe�"6�x4)T�Yc�s
Q��74������}��o�CCI ���(��;jg���}�eI����՘oά
�<�|I��w�jq[ʖ�܅'+߱�T1	��;M���n=�/4�T]e,�j3ǫi9~���Oٌ��#�&�c�#�������n^99�2��d�k���u���	�!�㒇v��(A���:�S�r����֐8��Au�@GX�c��(�x�Q۲�/��E�"�x�%7�RGm}bD�	��Et���i$�C��@�-d��B!��W�˄ܥ�Z�ثP�V�V�����^��M�"��G߷�>�Q.u��=�*�0'�.A}c�f�R8��΀���>h���r��a��{��򟼦�Q��r&g����X ��E�2�4F����i�8�/C+f"ZW-�Sƻ��L��㐈jt�~}w�gQ�׋/ȵE"���-5]��Dd���H
>ѩ�PZ�k��4_�Ý���W���M[�U����zyyN�y����1�7����(��Wj8{���`�UW��(0L����`ט�D�\��7[��>�(�Kc����+�W�7�u*ds��ј ��kd��~AE��h�A�W���o�׵@ې&A��q� �ʩ�M����4�����>*�
Q���p#|�Fε�I�Y�̒G���Ѿ�ؖ��;k.��2�=W� N0�
�:�WH���1�L�����������j�����_�ڈ���"}�K/J�D��q���dG3���1�?!�
���
(	738�,)���k�^k��	"�/�_صK�
�ئ���3u���\GUD�l��C]0������v���7z*>tc�Z�`a��2*�Tw|�xrmO��R{3@���������M`��
�x}�D��}FN�J��f�R��2����YK��U���@rN��T�G�|��U�L�?�n��~�'����@���}'
鐕A���)N�Q�^4IzXrUK�{��$����6��"�6k��^�lg�<eR��1��8�o��V3c�>8T'ij:7����Y׭��gQV���v�&.�:d�1j�o~cwۻ�寸����@k�=Ń�=7�	�(��C�c`ʸ�n�-���X���*���0�~"|}Oi�L깜H��y��$>ae��-�z��%�f��7G>|n���.֓�D�0Z��N	�� �R�-h��'������%N�=cT����$���c��9$)(��~k���x0tQw{��q�q2N��k@�q�2�)|~m9���W;RD"����!D2X�9ngmZdOT.���G����*QY�nCƗh�n�6^<��e�s�A��Ɋ*�p��v\Q�H%�K���	�[Ƥ�'<��~�ʀ{{՘F��	��� �e���h��p����P'�ݶ�MW�Y8Y���#Ǣk��Þ7v��v��`����]�b�ʖވ�3���`|K>����������׌|�`��#$�1�E4�)��v\/Ĳ�^x��|ˀ!^ý���]&�r�4L���h3�C�lD
V��
��*���Ɨ}����-��s�_ߵ$�tn����[74��d��$������
߃�[��)?��𫻠�#��4�Ԯ��/��2��L��f@�d_�~�wStj���4��>Y�`6#�]���y(:�B�W>����1*���HY�w�����X���ז���9ޞ�n���iJB�
�� Hhl����g^��W�1��A���m�S,�j�Q]���l}�t�i*	�I��Ϋ���1�x��޵@�?�3�����$:SW��)l6�CR��:/B���ͬ15�o����[� @�`}a��HA&�~�����B��]� s�U~���j�[9>�L0h�d3�~�Jݻ���.�\_{���_#��+�`����_F�ApL��A,�7���d��.�;ԝ8��>������DD�Ni
��ܳP.����4�2�����4z�AuFTx�j�Ї��G(W9�v@�>a[	MHe�&;V\c�ƹ��o��mt�@������X��`�M�-�H�F� 2�QO������JR��5�.{M�֠����bBtQ��z�ľ`��z�Ǘ�b8[���6	���������Iݜ/�O!>��)�#[���>(ah,��U��a�4��*RW�t#~���)e�[��}]�Fs��u��}��F#w��M(�X�d����J���YQ�<�;1��]��}0�ň���c̼�&��.��Z(b��k/���+��8P�zW%J,��7/��7�x(�o�#�M^P��23:I�{�ܭ�]�>��`�����E:��;�D隴�lB�p-���t�34}����}�G��r-��q�SL@G��3Ӗg��B��C�C��~��%/mY�WԬf�wӿ��X̮1O����P���� �}�W~A>Է�E�ր�P�%���=a��s1ؙ�wd"n&�=(�� ���r�7���*�@�s-���y�����>�d'�>��F��@7z�,��,��q{���m~@�I��FJ ��c�yC�����O�mD��Շڥ�'���RC��
h����DW�ضCOk�-�w�Q�O������1�3$�(��O���	�};Qox�Q�&��ef�7*90u��DE�KF2-U�^;��l�J����ܰx��(��I}��v'_�G��[��Þ߽>?ع�]�C�	b��^���C�E^��\�v��V���$A
%H�F�s�y�˓�eŝ$�K���tоU%���Q�
�o��;;Oi���4;���2t����9����2���ܚ<3vmV�e�(ay5�l��T��Nr�A�#�����:qʄO�;Mt�T#v��4c��K(��{�7�g��B��x+�1-a��|ˊm+�6	9���.b����B4��ey:��?��x�a["rY+�Mq~�PNٲl�.B�
/�^])���.b)l�N����:{��+5k��2!͠��������Sg�}������*��1��� ]�:�u��(�N��GyR��|+Dg��o	����.�&4�bC�|n���� ��9������Sg�a���~��#������)Y���S�m/�̒z< ��/Y�u،g�%M�^%6#�H.6����iq7�:�)X.#ܙ��d9��*q�1jS� ��z�`�aeWr%��L]3$����e��C��sC8r`�;#���0�Q-
<��ACB��`tD#$��H~��O��q�����V\����,�qftM5|�qk�,�G��ʹľ�OVU�T�!�'�@�U(���2o���J�����g�B�<�����ZE`����,.��*U6�����ތ@O;��2����D��5����":g2��`,_��HK�%�'��j�.�ȧ����p���JS���L���hH�ͫ��
���W�(my0H=E�Q3s��6<�k5X�˭��c">�x���mX�٤�x�m"z���~���VIjȆ[���i�\���У���j�-�j˭��n[s�P��P�*�_�K3��pW
�*U���?k��� ��q���Y� y�D0�Q�hl���[\O=H8ytfT(z��Zɠd�N��܏{�\��{�z�J�m�Z��)���S}k����c9��5�u'����sFH�G��D����:����:�F�l�%�dHǟl���'�.!���k���{�BhlV�r�^M1�X�&e��_�)�3��)��J��+��[���`�]��T������1�1��qu(Ŋ}GK�閇�W�WN<��a�6�3�鯨e�����zq�s���٪�`)��i+����ō��t��o�";k=�=,m(u���+7¼�E\\�ӲZSs�|�j����v��k�W��Hhv��r^MMVϋ�/|�ev�����dx���s�-A>�j8}���"�X����橐i��ߵ-e��J0���{���/��5��:���ދ�t��*ՍŮ�F~����z͟�
!�H�k8C��]�*�� ��%���
�k kW��eP�cG��(Byl��cJ�78;6�o6T������_o$M�]����i(��N)\�_��)���l�z������}S�f.mGO����F�L|�2����_1��'�(S�@�/�ߍ�BXgЍ��"J;6����%S���^$4�d�n���d�=�A=-c�ô�J,�޾E���$�Q�������W��~]�2B��쫵��Kf?1AHM#U~�,t�Nh~�+�"&��eU�����X�2�!��CR����H:�B�Ȗ�űԊ������z���+#g�� �ˡv+�mv	1�ݝ~0@�hLL����'�Wѩs�dV$����dX�i��Y���U�� �I*G4&���0�>4��ͻr]X�s$��n$N��џ��dx'�&2/���_l�N�:�\����f=��ɚ�c.��̉Y�o1D9����gT�rȌ�����x�0G�6�o�#:��ј���<�5�
?D�f�Ư=��:����P+��SR��]��|	�v��*1��?Zs�GM�^��#�CT�2�ڱ�����5D�ޡ+H�Ph����X�t�/�Hk�Ґi/����VA�8N�=���J��'�vt���ee�����]3��2I3���>�h��q����r`��J{J`i�8��3�)�������ʴ+�+�TDEV�����Ү�2����v$`���5���̪�z"�0��(��R�ճG�\����_g3�F��W�󒯾�Z0��!����'�O����8��Ibm���Ͽ�=��ȱ%\��u�j+aI�	|��^%B��ƥ�ӓShɵ��Ζ��}��Ԯ�1`.q����F�:L�;WD�<��Ϊ��c%�m�9H	�	�%A�-*�w	�[�s��P��<���0� �e	!�:�����R�����
M�
���3��������n���7h���"3L�/6�a���埨ז�dv�<�]3����Gv(��I*~Y��O�n�^֨4�_�R��(���h�s�܏&�� �]��_�z(l.�U�h<�Z�����?C	��BՊ;/�W�8�_U[J�;%�B_�{Ȏ%H�r' �8�y�t�g���}Ҡ�u�Iw-=���q��&{���������fc��z���+��x��&w
X{,;�~-F?����-�T�L,�k� @��������ƒ�gA6H)X��>6�]a��C�[��b���H'���~�����
�%]NH� 6�{�����ͪ>��.9��٭T���a4[D���<#���l�ibQg>���>�*؟��S�sg�հ>I��x�o&�
�.4IN��yDu��e^�Bdm�S; �¨��Os�ǳH�]Qa����h��|`B��T)]h{`��~�b2U\�x��� I�gnU�\==O�������Ç$�4g �U �mX�7���f��h�Z����O8������,O(<vh+4{�O:Qɋ��W7Q����ϣ�D��7��_�/jT.��5'��CG�v@?��jK��$��hL��C mq�� *�<�o������а��|��%�M������?s�ѩ���+��s�f�_�?7�K����?��{��B����%�}ev�k��Wx��U��{������"'5��Iz�����u��yy�خNt���(tݼ��?��o�)G��]Oex����ǃU�J�v�-�h��9���Q�}�%�2�Ⱦn�r�G�;)�;��������P5�P��f�5�j`5��b�6B�����v��l���
���?���o]Ë�ii��� A��yc֑����pI1uF�4��T�u��͘�s`����6?��ͼ��^�X�ø��I�le:x����'�!�4C�Z:+}�)��12�+��n�݆ ���!v����[_ɰ	ȗ�
p䪫��.V�z)D}*~��Q��e��D���s��K��'E�82I���k�'4E��f?� `��i'�/�{X��m�8�{��VW@�'Q�{["��P.x֯*��<ij�
W�
Z�׺x�-�z\�`�����U��ٺ8?fSEo���-�����C9��5?�y�V"�Yq]�'|pr�a
�2�X�X����
�E3����!��3���Uڒ�L��<T�A(~��$��(|q�7���tG� r�H?�*?��=��`�ݶ��RƲ)dR\� ���uR���\�]$	a���Z�\���=�8��a�mc�1���4�<ux@2����Ti[N�}WX��_r��p2��a92Ӱ`��s���K��K�wP	�~��7� ���� �h?�'�bC��܍�萉�:P�\�����A6�׷Y��Z�#b�z=������&�!�^l^U7��m�Z���7��?Z�Om�t+���C���)IƵ�%x��;�=�k�k����[����¡6F�-`J�S��� ��Wl1��%�N}��^q���K���-�ǣ�m���� ��>�s����hH^�	�����&'\l�z�Z�l=.9?����G�R*ͩ�8�z�~6��5B�Xϑ��!���\��d0��9/��;s5� ��(L�
�"�s*R�I��y��	@���'��_HeȽ72�!�Q���L;�:���M�!=~wz��� NHb�"KV,(����zؙh�V�J΁@��%��ko�~7K�����
��C�B#g�+�(��� �$ �,�� j#	�{f
����8Wד
ѐ[�t���,.#z8`ۙ�b}�1!9|�%I͢�[��d�,��Y{������M��_�Ƅ^�� �[�ŗ�7H���{L�{���{�kmvz�
~R�Sp�����$K��8�`��b�<&��D/-X�A!o˰�Z9�*��ԩ��&g6�X�렃���#�$\�!^�]�����L[&0FB+O�"뽄��Ì4+��W\cF$��<�=���$��'HH�`.GUi��~��{u-�5<�*��g0�@����R�7@����1�8Ϲ|��D'����Z㮊Dv�� D���?.�ԑ9M<��N���+� �!��u��R�,�߻�>���8=�}�$�Ė��;f�)�sznm~<���nsՆ=P`��ȫD�fO�uymy,6<�����xH�{�'�ʅ���J/����,�v���cOxi�KN��nj6���y��t�d�Ͻ��"�Xt)}%��E�Z��%��n.�Qi�RF��Y�|D䭶2�2T�z:g��&�SO��n�3,�=�N�	�l<�-��kQP����^3�n��lO���u	���s/BW�w���C$�FF��O�ݍZD���{/�� ���!}C����T/ ��\6)�禳]���U>FWؿ�L����_D*���H.-̄wDt������Y�1���_z�7�aF�5f�{훠"J6�G�v`��a��T*��ȋ���$��:�p[GJ��Ink�Z�A�}�\���/�lo�z
P!dN�8e��7�|�9�	�C��0RLӼa>nt
I{��5\:٦	�GRY�U�dI}w�a�F��Cز&F�Y�R��)��r��s�А�R�֢ �J��Y�h�izN���Q��`�3b"R}'}�%7�-�i�26qT��b<I޿����.��XÖ#X�Q�����T=m[׻	��3FMXcHD�rkrA(� N��f���˰��H��K����s�?`��9+ĕ��t��R~LoH�n���R8q!\ksW�;���P�y������Ihe����_?�:0;���y͓g4\zI�}E	��_6o�Sfj���ҭ٩b�zy�V��f@����x�DI�{�/�*@ǹ�ա�(p����&��� L1�}��2/f	Σ䞐$7//��1��|
�d�ep�nik�r��z���U���b�Yٙ���y��O2�M��<t���2>H���P�*�(�*�e0�4 <2��I�
���� �u�Y%*�i)��g�&�.MJڄ��e�0����Ad�Bn�gNFO�d�R�>;��D�޶����'����x�Ʈ*:X8צCM[G����1�\�������X���lYpL�C���"]�:c��$��I !ˑx�� �KC�+{^�F!JyA���9?w�W�0��4�{��j.(F.��m���T�+�P/�Ʋ����K��|G^�މ��;�2ÛgO_�%	��?H�Oh
��8#�
@�~	�BWPj����F<ci�"��KÌ�g�D���<�=�H?`�>W1#��V3yB���]���k�VGNp#���y�n�.5�9z���~DOx��0� ��`���"ؔ ĊJA��mLA"{�O�9F!Oz�s\y����,n����F�a�P	YGT���
9{����sǣ�Ξ�M���'����y��y�I��BY�iW����i�w�a�BqT��i:7��-\�Uй������C�ǜ�1��|���!hb�F&[bK�J�v���s��)�5��*���m^Z*�{�u�heA"k??��<�zgN��m�q9��r��*���k��E��1m����*�ߢd�ٚ���v�X7���"5��!\ټ՜�	�����O�ܪ���g��9�|���CV�ބ*4���f&Y��� -�Ŷ��N��زp��O��d�uF��W<�1�|F��L��@Wvh�=���ٺX
�'7x�%?~�C����,�/}Z=�Ȳ/|�[��|dA��������)%����WE��y=��p(�����F�I���-i���s~�j\e����$[N�ћ��P-4�}$8W�d�b"b�k">�_z�@�,��`z��7���Y����5�f���%>��K�"�3����~M�� �V$q�p��P�q��)^u:����@��+2��<lO[�Vx�LEX�<�]��-�g���c�D���z�O���gr��b��NXw04Av@)ly�zhr#��gWީ�:�ב�� -��V`�bi���u���(G�������&/����{Ү�sk,r��r�F^����Y[�"v�lρ���R�MOv_��
��v����w���7��0����	����@ګ�^?t.ԗ�������=�A�[�҂$0���m�ʫ��z���L:�/�� ��<��ŉḣ�n�K�)m��7���e�Sɛۘ�}ێ�D �C�`w���:����K�P�)��wH��d@�q,!g��措M�Qu��?�b$Ltܿ^��g�OAz���;��1sۊ٬�K�<��D�a�o���!����б�K�}S\�����?��U(?��O�I>�J���q�Z&^��׺IW��r8�ҮL0�BUm����aW]�� O�$����ڨlV����Z\�m�}�od��f�l����4o�7���f��ƎWz�]�SA��N���Xm��I������k��]`>)o9`��p��5�Q wpL�i�S&��F���D=7���<ym�6
+"��A�6�cv���@౦Ov�d%Ѻ�8iU�I��ac�&����=�i�A�G�u��1�?�8H��� 2����)۬��4���U����	Y@P�����p��R�$��(�>td�h�f����瀑�FQ�t&]�!ћ�e��8��V 亞� ����AlZ@�]Fnǉ,��$�'PǏØ��#��c c��3ti�J��ś�[E>�<<n�P�}��Q�!�/1�:nHsƦ_ŽW���h �M����'��]v>?W����TZN`�tk�Ȍ����6ZA}�+��8_�Hq��a�6~ZBP�Զ��A.&��9�?��;���?��O�{ͩ���  ���ݲ��4���.����$�X[���p��s&(�1j%CY]{�[�/{��S�Y�?y�}j���#��ނ9�g��� ��y�w���zKN>V�<���\M��>w�XG%�(�����z�iv~��]����\�`��P&C�����Yڷkkq�*M;m��W����&+�
�������v�I��	R�� Q%=�����-[X:N]n	��i1.��L<��Z��CYN�[�l�{��F�nSG3]���8�T���ߒ��[�j�����^�C3���ۈڪ�{˥���{�����J�X�`�o���\=���$ak]��3s;y��~���������d�Q�FqD�7��J}�`|b�U�a�au�1�8�F�[�G{��#�^���{��������ߛTu�m_�kp�=oz�d��I����hO>� ���,"�&�t>� ���R7Hc��~㢬�y��e~���է�t�g�:{=i�sFB)����돤H��T��M<@>[?��Ց�	b�[�"%�W�V��/��D������=L͒=`��/!���yY�{G��'�Xq�$R�&�ƿc�������|,����F%gnB�_߆Z�~t�$=#EH�5y�Jmk��aV��O���wO���)���:����k�:�}�����پf�q����;��f�J|�:M��yH�5o��P���6�Ƞ��0T�)!���f���w�H[���M���$XЬ��?����t�;_s�^�� 6���95j���G{�"!���ӓS�n�0��}�R�ȱ��5��]�MI@��~��dD��"��ǿ�P���Y��@�?�T��_,�23��n1R-��"���ȧ���,p����ݫ�NVZů0%H���ِ�-��S+g��]�	����h�h8�y�h~��֋�b�Sk��Y�?B-y��y����pp�-�{􇁆qt�r���)�c�0�b�I����8������t7�]�36��7 �ɷ������r �t7Z���.�z�,�mA�(U4�C.���HP9��\�ٹ�"�����և��G�')�]R
(j��0�X���\�L�DvmDxl�&<j�x7�ŦR�F��M�*���#Q���k"��H)�Ȇ���T��)��.�h�[�Q���5�o�Jjh[ ^�F�O��Gz���%����]@5$3�_q�1vX����_�{$P��`�w�+�~4Kk>&��)�Xn��sl���؈��~W#iV1\��������6�GI�.�_J���Gf~��E^]�n���wb���S��1�|g]8n
L��is+4����@�|T�[<K �N\?QswT��>;o0h���c��8�4�k���,M�n�O��5�(�(4��fV⼍��3�SQ@�� ��̨{
�a_��Wm��n���{�����4nrU�	Qk9lZA���܁$9t���o.[�txtq|�R*u�>�B,B�����ړւ�g����d��Ĥ�����|���l���.�p҉�Y�\B%��w�yO{�kM�*��_@���_�%S�K�V�������]d���<�����?�"�r5��P�����D�t�����w�G|�W,&��qGs���A|��_����
y��ܒ�O[*�x�Er����__�Q�|��1�rP���'d&��X5���M���� ���T�l��mSF����Z�p�p�*EM�ϑ6ߐۇg��u�-���S��vH�T�	2�?9�r-g�!y��_�i|Ҹ��D��5�콘A�1�=��ww��Y��e	L�w�i�T&���l��ѱ�B��z#�`�H!�)	�|5���nWN7�<q���B�Č�a=�� �bb�c��n]f�f��p��CGnQ
m�"�@[��{Uu	2��x�}7�#�NT�.q��6���9E�J�c�'{>����y���v>Q�t|� �����Y*H������|�	���~�g�U����$���.�9]k�m�΂��@f�|�T�YRV��'�F����l�0���#ɣgώ�����5� �|�\����M}�J�����.����?j���Vغ;�&�~,�m/�m� 4@�xh���RgPAZ~
�xhlqћ	͠s ����`��U,�ꔚ��2�9����\Lކ7���P4��=�d�`~C.�"�ؖxUxA,�C��n�b�Q����0vQj�/�-�8��[������!V�֡�(�	>���( -1H����H�ms�1t��S�Ҫ��@,�Vr�/mq�:s�,vh�9��Z���ʜ�on��EQ���ȏ��g�9�=ҹp	7�ęxv�غ?��HQҳ3���<aG�(%���R��1!��b?�Ҍ@�1�R�k.gUM��N��UJ��K�?��Ig�n�~h����̈́��=�;�q��?�=���3�Qm"�m"���n��i����z^�[�đ�O��]Mh�b�����Ry��������!��m��}�)x(B��
b�M���t�ǠW�m���e��������� (Y�G��,�E�d1��#�L��\^�;�(��HX�ȍ�-A>qf�5ZQ�!�#�#����t���~Mc״��)o�#�r�:bHBH.*���C��h''2[a���GO%�*.�S��kG��6��+�}��_^߾�Ĵ��;�	H��O��{�m��:�b�	����Q|�����';.F�C:��~���1���2���i�
O��8��.y ��q�T��Fh�s�#@#��ݓ؂�:�ѻ��ۊ+	�wӍ`��Bz�T,C�2j�~����tQ!�v�j��/�҉
_t���1�4Dd�[��s�H����o5�kFJ�9�O��ҽ�Xl����F���s��e�r
�K�*8'F���[�rD5zĝ��{,\�v�ONv�ȩ^�`���-@°wXьvh�2Ҥ����>�B�jj���L��$&�S�c�8�� ^�1u�I �=��H)	9x�7�b��,8���|�s��i�T���v[�qD�P��/� �A���R!C����� ���^�/����@��!թJ��hV�+oA���B��[�PJ8Y��3_���u����˾�o,}pb�BϨ1���sܗ�����f��"�ѯmir��@��5�F�3�YUs݅������e�	�7y����i~i��b伲J��Ԏ����"o
�t�7Ү7����V��H~����EIQ��X$ZV�P�� GO����o����G㡵�޵�B��P_Cݓ�<$Ԅ8���PZ �+J�_��1 >�� d�$�2��LjM3�)��)ʻS������]�<�;�9"����ոG�&��2�IEW@_�A-�F��ԑ��Ԩ��@f-�Q��x���Gf�~���}	�sPP���1s�Lv����Q(��q���⽇E�V�'EBp��&�?7H?�2v'���d����)y�]������~Cѷ��ˮHl�V�c�5/k�������1Z��)J��VxޚC ���#R#�g�}�!���5oj�\iZ}U<)W=H><8��S V�� �wf$O�U�f�������qq�Jc���&V����r47�F�9�s�8�~[�K�?,�]A@I��;�]#fCӤ;�,X�v3�
Y�O�-"ÝV����8Pt��L�(4���yqW�U�������e�O�F�C���)$�f+�j=�;NJh��k5T���S��AI$�����ݛ.ǰIH���Fţ�@Ϥ�.��`��頾�ϓR�Ky���J�#�IV�M4h,�c>������L��'*��bZ�kJ:���{�;REW�*C���e���%��^�9����ǶQȽw0�ݚ=�|�����G� MO#�� ���/m���*�!�yP'�i�N��$*$�i ��$��T�>^�Y螌ي���>�A%5=8>X�ֳЈ�p�� �ఉ����$�ͮ�F�O����$nmk��!C��$�T�u�Q����/c�Ma�8��Wz��o�56T�v�~�#�0���?����Z������}��x^�^z&��:�*�{S��۹mO��~��f�����g� 5p퍤�Iq����~��J	��j�d�n��߅ʆ��q���Sw�]�HR�tź��<y�y�������)wܧ��&]�25���kW�ɨSn0�
�8��pisp����&�*��]��&f�?�nh��ͧh��8�#R�B���� PZ���b��U�]ë��_��P����i�%�@���Rp~� ��D��ù)��v�����+�5ka�t���u��,��� ��*	�W
�ʄZ�q�4+,9ꝭF�!�����ᥠ��3�Y���(;ߎs}n��2�JB�Ǒ����o�eW;�m-�9��3;�7G���43em۠���3��?װ��[�c4�4�/�&p-%Y�%^mY�����M� B�"�s�'4<�>p㶃�ˍS�}�I�;J[{C�-��&�8k�@�{ѣΌ ��&W�(jf�����Ԛ�T`�R��'F|���լ�+jFF��Œ2)n����?�� cP����8J����@i�	S,�������lxL�pB`�>�j�0&�\�G�������'1��j��陿E�8���N֫��},ⶅ��ǳWH���G���}����A����X�����337lcA9�T"c��d�h*آ��*�Kr%="��mA'͢�~�У�&�I�<����i��A�	���[��5�0�#/>۴P+�X�W�ʢ=���Q�r(��;�4���5h5����?�Y�"����Ţ�_u���"�ڮ�$#So�q�,O�O��虖��;J�Լ����:� Ơz�ʹ�?���@v6��7�3*9�N�8�mYTeT��
�z�(&��v��*ƻ�u0o$��.��F�������,T(�p������m���]��nx=\�/�N�����A��|B��K��&�ƣ��<���H�QD	�EY�s^�=#��.���'��r��O�O�j��w[�_��B��+;��ܲ���wK�;'+nk�a�����R�xs�n��;{����$��Y������i5v�T�$�LB!*��)�6o����{ccc�$` �
�JCsS����l[����$e=�//U@�i�x���SMRiDO��_�J�Yҋ9j�G���K� Aq8��L��� r���Z��.4��#Ɗ/%E�M���u�B'��D�#\z��jI��
�^s�t9*��ʻJ�v�;� �`�p���U�h?��r0�bp�ο䄐������Qd���,��(|�X��F�P�0�5W��F�lHoK�~����h�-��!��~iRx��rp�f���	�:a��U����@�1ro|���:rb(��L�ʸ<*&��10��6�����/�����[ͨ'U�������41,Q��u8t�o����� �>���C��S�r�V;�u��y�~%�\�����F�5��E]ѐ�iĵy��~>Ji��˰o�?Z�mc�=���S����a�g�n|b��7c��#����9T��{.yˡ�.f
%�-��>ɣۊX�.�,���*����6��
�ƪ	UXA�EP3(�/���i?���eM���E 9�m2/�K���+�T���R�| )|�d�ũ���']��9������PC]�;y�rcu��7·oz^��ʰVɗ2ূ��74 Q�,�f'oe٣�i�Z�*�r4M�t��	K;~�:[%3X�cf� �=�ܡ��tK�_Yܔ$[t� ������߀�T^񖹀E>���k#�����R�C�'<�σ]�'P��Ƿq��h&�-a�&��P��}$w��P����x��z~�|\a��=���ɛ�R����bKg���o�T*�x?��K\z3�x����5m8��S�Jwh��+X �'V���Gߚ?f�cϺGw����+p��r0�
�C���s�ı�Y]?�a#�qK���v��]{�xK�2�_��P����I��v���0��W�ב{.��m��C���<i�Яv�/�!;S�I�Q�?><�c���e�؃"�g���yQ�L�ZT��H��^p��9_%E���a���x�Nx�O5v���9�^\;5���>����j���WO���PKM<�F�mB�7�Ў��y�=;�z����#�=o�v��K���_�`����	��j[������ۣ8h��~w��e5��\��j���"7"��C'��L�P�#E�Z�_O�4u��KG {c2g����߰�Q���p&��Ƒ͡"�PC��z�mڎ<���X�Sfԅ�G"��X�q�R�:�.`�f�ͫ(��f�x7oH�ԡ��{ ����!��������{�)}�_�d��?u:�[z���g5�U���?�����&xʠ�g&*|A��/F�5���C���N�\�D2��>�����j|	��\2�֟��)V�7�x6����q��,[p�_����[�}���\�s!@��`��&�@�OJ���G@"cT��s�c�7�n4���l�-'�<���w���I�4��C��G;�#ք���Btk�c�#q��zXNӬ��8��u�����U�t]_~9�~A�z>�
u�=��R�Dj�w$��LT���R����a�z�K�@�*;��n��dP�r��P�Y˵A[�]%���Icʐ�q��]H�B�������ݵRr	�V� �u1d�x]�?�/���h�/�_d=���(3w-"|R��bY�P=����+|�$~X�tA�R~Q�m����U����׿N�����/����Bc����d��<rع$��_�)�?eOu	<�J ������҉]��B*�f�4��YA�Gb�DRӬ�/���+�5��F�$��"�tt�|����Q=d��u��O撄����Y��`$춏P�ϳCtb�5�Dlm��~�A��[���WJF(���Cd�b�	��R*��֚����Ʀ�~���D(�+������l��I�ayh+�T�g�v��������4lЍ����xPD�:���L���~�2���QK+��N^�cJ/u7>R���X^C��V�o�`m���!
h�!{~jna�I����n�<�l��#z��T�6ݧ��d^U��sE��?T��I�!�G@y�'.���@����mOH>LQ?�j��*Ce�3���{ZM�7c�t���W,�"�a:6�}�&g�q�j ������j�/
7����Fi���4��`a<�)Sy���*i��_3����UH���Fz���|��yt���H��z�:?���sK	�6
"���:��<�;5Ǭ�V��l�+����ߟ��z ]�,�8FP�S���D{4⡵����@D�mH�5���0zC
i;�z$�:;��eZ��kסP3y�݄�cY���R���LL
��x��uᐫl�k%��}����Q��C+5#�����$��k�2�����,]Ƹ��GM'�47�(��̛�h=7��uŴE��z���C(Eݽ%���c\f��ľ�,�nk�����ՄW�ۯ߄�\ Nq´:>V��9)���EF㿓�,{k�7fFk�Z
�^�G=�5A����[�?Nޒ�����N=�kද����� q��E�ۿ��jS�����:�c�*]?�/���O���T4�d;@����o��rV,��ҋt$lnW�a�N�����u�e�2��ԓ�*�hQ������7*�]	�W7� ���w�ktK�:Ef���~C�7��GӃ{���/ѧ��Jf,��n�x;6��b��Y�~���,؝�?����\��P��2�*n�6�R��2�Bc�t&`u�-?��(YC����� ck/=Ā����ځV�����i�UH�C�!\��ٮ�R/�?�f~��p{�}�U8͟��MB$ Sݟxj��V�zxK�'0S)��l<AKX9N\�<���9_G����9T�s��
��Tg���I������+�-Z �Zr)"?��ȩ�mE���Z������D��34<q����̓���kZ\�AT��]���Ms��Q��8� ii���BrP��@�FɩT�*C7�rAR�`r�I���U�ќv+W2��_4���/�:]1cյ�|�#���;�O��w�:T������A[ �0��% K�nT���9=��J��Gz���#OL� �1C'�LV�)�r\J�ѓ�l������BBXܼF�r#*l���/6��x O�7�an���$9 v��ŋ"�6X덲L�*|gx�8q7�s-U]-q�<���+O���E�/����rC�J!S��C�e�M�1�1C�5�*��M8���7N;�ԣ㘏DV&��O�G��
3��%�z�V-d+B
!�s:{/��6x�@W�޶v�
�5���E�霣fħR@��S'�Q����?��Y�� ���f�=���W6g4Z�*�\�d�z0��%����<O���n>x�RrY,�r�F'�}�4�����`Q���:��3�z4�z�S�i��9q=��ُH����B�
�y��Z,K*�Y�~�xh�6��3�찢3��v���G�
�m��࣏+6�qT�11u��!n��r`�!��>�
�����㠐%���#���~�͹j�}���Z���%b�`�a*�ico�wάm2"�YJYN�����2kI��uQ�";����6������p:��0�ބ�;��m�7>�!O+!���~x���L�o|�;���,o�*����E�N�G&�DQ����x�3^�Ѣ/I�Լ��@ŀ����le�:=�����Db��N3�h��x�q�0�/���0�|����/�OĨ}��rd5��ŐI4�^,̒�����"��霳'�&��5BS��.� ]��C�������;TD��濚�h�uʯz���~�}�{��iG�w�	�M5����T�Ė��".�>��j�y.��Ǐ-��ݟ��'óe�j����Y~T��ՅI��=
A�'��=��8�Lg�n�k�"���	�K��:��D�9��ؙϼrE���4��J�y6kI��Jj��%fC��H��\
��h�.�|�-�}
�h����U�a��-��s&�靰v�)h�y��~7:�����]����З�9�c�-|�P�Q&��v|�p)��Y�gOck�� �X�����b'���Ġ=ݬ`�B��%�c{�A��#�u��r�>ö�k�On�o��q���R��$��h����R�h8e^�F�
��&���#��k��/�,J%��FE�3�Bbʫ�&�E r4�T^��Fi%���|�#O5g���`�Ky�M�a�пw��L��d�Gyj�-�0�r��u)gSE��2���j+�+?39.?���v �9�����Ju�Z`��-���W�%�|Ne���K�C�ΐ�e&N�oa~F%ZKgq�^����W� }y��ٙDn]���X?�l�Hk)�Ao���p�3��d9���%�NAg� ����*x����	a��Kx.K�0=��p7IY��A=����Q+��BA��\r�?�/��nT�[�#�X5B���޳�`c��B���#P��
�ۻ��v�#�@��t�u!RR�����ɶ����w������qTm������C�|�4�������6��""�*�%^C ���P�z�3]��+ ��Yc�x`�����tU$1F�+%t��A÷��U�D���"��Y�LiD��%ۥf�����j�V��U`��4����Oo�d�Q�N�?⦙��)P��M":�|x�`U�NSצ����3�Υ1=І���Y j��A�6�W���E���E�E��b�ԫ�[�9���}�8d���a�%��H[��������>�i��0,L�����e�wF�	����o��"�{�k��.�3�⿠��u�� <,'Y�Y�ý�ٳ�X�zw�����m����^��D[Q�_,����Xp��!U�^?���=s���w2{������Itvgћ���Or����4u,�����Z���m�f#��.�O^�L�V��|����-�u�q�߲�_b��B�Vt]*`[�:���)2��xS�E#^�Ϥ�&�����p�VKLi.p��{i�ALk�crG Uj.�K+-:k�Q��5�X	uA����\OR�G�&�F�q@���6��L6���!:���.o*�Ї�y?�?�JJ�G�Ufs썂�Vd���H��􉲤r\��g�mF�WV��+QF`������9v9i~x�֥pY4B���o��-гE�J�M�d�i����v�ᗠOA�囤���+�˄��3�lS聥̉t��	$3����AL��W}����1K��^���o+�R�g���r�vLֹ��oC 
ԖwI��B~�ʴ�WI�j.6�)|̴r���T��Rĕc�\Y���b�2��r�&���� @Ii��!BEjex.���Cbb�!�l��ؚ��y�Q�N��{����O��yF1'���&��!����XВ��iy����b	m}��<�}��<Nb�$B4�'$�c��h�{)��fv��Z�@t�";C���k^[_~�r���=�=��W����c�I��J.����J^������hߍHńЛ�a��^�eѮ� ���8���X�ĪĢ���ᐅ��>���P��1��,�.�1EZ{S4�2^��e0+3kd�L�$�"THYNt�ު���݇2�*���������: V��}�U����pc�3.qΤF���Ȧ5K[��g�7kc�e�,)@�_S��+�g�/7��b�T�K�>i�2��O��N~��T����X�O�)��}I-O$-��pڽ��'�4�ozzs�<���M-O,� G��HEV��r�ʨѳ����.�P�̧��U+��Ǜ����)5Tস.��Q�����^L�Rը{�M��Tm\H�Ih��q�O���?�΂�/@�
����孩��5���/j��{���/"skJ���3��S2�l��D+�օ$.g0l�����I�Wlͺꄃ��>��7�ť��\�O�������~!�RȢ]V3�~<�{X��7��Kx���n�����J��"��%�����?e΂&T#�Q�5"태���K�����w�����r3z��^����8i%��}&~%uw�Ԇ��+*�Ԉߏ����E���C��y�6#���0�����7�;<k&���d��h裥d;�ш�D������n�`�rW>���@d�4ߩv�c��Ι/[��Y2�>���g��"�U�߳@���^��UL�_������4��I��Y�E��gl%)ٹ�R�Ze�#��I)�j��1.3~��Y2��A����Ij�=���EP��3�ӭ�-�<��[�1�V���.��hjVU�6���XU����`�ą���L����$�o�<��.+k��L���s0�ɪ�	J�u0������^D ��C�(f0��"@k��6���EՒ�6Y',p�	�>#��Z��T$�T���{�i��bU��12X�۫��i��>f��[���-�^h��K;�Xz�$���0kt3z��V�b$�-7Cň�"��6b!��UH��d�s���o��;��@��L�X�{�����$��ٝ>1Ѧ�\~B��'%�{��]�d���	ȖR��TJ䢑t������7A��߸�<+����n
�3�m�(reU�h��"*'R�-Y�� �/��ۊ��.l�x�	|�%�l�
v��%(+�w_y��y��ЇB���g!ng�7Ͷo�[2�&�m�bm�zf�E���M�S���q?l��P�vu�G�w��@��'d�:T���My�����	Ȗ��韎z��{�!M�{�qk�'<���Yߌ�?�`�oo�N�t��5{��1�����e�y9�41�3%���ʣC ̕I&��	#����ЊlP:�9]U��{`O]�
�(��Ҩ�G��U��A�B��2,�x���8���8^�9G�o�,����>OS��-�rS]2���(o�p<��y�M�:iE��N~mqA1Wc#㳱�Q��7P��ƽ�¦�snF���^��-���1µ��ĩd*���O��ޯB%ڽ�v�.��ϐb��b�~�څ�jLIޘ'T͉���7�$�B����xT���}w��.$/ ���;է� */����UC5�պ��υ�=��a����&�7��qGh��!�Xm)�A%���2e�6="����p���A���7�܀;��;��6�U��&#-%/*�����s����s�E�xB#�HU���$�B�E�$f���Lv�{��qa.sJi�����z�M	�0�%ɹ����"�<+�,�` �jʖ�]��9�/��Sx���
�O��_9�C�9�ƥ%p��0"�a�v%/��9ud@i��/B<���:f|[��Z�Z��ǁ]\b&ߧ	W�؈(iG>n��?���]�s�P������!Hⷬ����¿o7��rh�©�G�n��֘����\ʛ��/P�WٝWZ��fq�rtB�A`�7�_h��ET�q��x��%�{l�����(٢��2`�ͩF�6;`�k����]K��h�����ۣU	�3���׾�V�'�8��W�x��c
=y2� ��k�-F���0a#�A�#�o8��)���~��HDT���ܿ�\2�2�a-Vޔ�~�@	��"��%�@��d�B9��luo�F�������`�p���	t����6AJ��U��U�b^]I+��qB��g>��s��~�1��ɹ��w��l�W��1��` sL��+��5��+�l��!+S�T#�{W��Pch�n׫ ���/�Lt��:��~z}8�� �8�ڭ`f�w:t]B�t�I���2+��������E���Ǔ�X�n#�oMF��Z���+��?�a��;!�>B��]�T��X!��f�,Yxh8?��}he+�Ɵ�o)K;�I��^"�U���9����R���i��k�C�9�U߄��-�'ϟY#�K�s�ɽT�f��z�1�u���'+2g.��Q��;n����{:d= 1�7��;��Rv-",�����������`+��>�U��(&����9݈��|���
9����w���4���no��E�#��z�d�y��!�{I���b\[���'�&r�H���o��7��8�LyB�*��:oB��0��w<�C���A�y[��R!V�{ҫ`��ŨYX�)L�&Yx�Z�pY(GU��;Fн����\���:S�	'a��n�<F!�,Rb�g�@��NK�e�������sВ:8�F̅������:h��MQX^H\�S=�6��<UC�\���P�m:�(�j�eZ���&>ձ-4��z��n�ӕ��ʲ��5�zA�Oe��N�-��nz��QLYw�r��qҊ�N���X�(��Y;zX��q]#rJ�Ct�_0��tp��A���Y������qhǣ�$T�뱛ϴ������N�x.��4��&j�9�J1�V��;>�.''mዝSk��ڼ����Y4۩�Y��O�D(��og1��7�1,�r鸇�z� ��|�&� �#��@��^V��)�RW�Nd�+�_Y������l	����&*���O?׋���A���O�WA���(��*D!�۞�#0B�o�nF��$y�#r�/`��4���Ǖp��bb}xS�	C��ᏸ���1!�j����_|+��D
�;��&��Gp�Phӝwa0zE��f�3Xy�r��i>I�9�"z��JX5z�(����L�����'��%������#�F�_U����4"Ή7���y]\c�(���$e�CsL�䊜����)�݄B̶n�cq�!uvΝb�X�Y=~p�!�K�ʓ���}L�}�/�B�<H(/��� 􀌎�*�i�q0;B��9͌5�@�)ꯒҙ6<h��{�z=[?V����j�ٛ��B�Ŀg����[�!���.���� #����'I[1Syc+�ݷ\��Z~7+�b�֨��օ707�,�(_0�q^�c���6�77��Ʃ������� �l���c�ր;j��)X@^3}&��(��y��Um��C+���du������pa!��6!i!��.�`���׋����_m�O�OZJ?�oР��S�qj~�L�Y	o���q ���Q�8H`�s���o �����AOq�a6��]H+݊�:3�k��,H!�����hq �;��������������4�3^�L�%}$�5��������E��3vâ��r����IA���"��O��g�
�2m�b�ӂﱤr��)]��}S���
)B=�\%5h���Yx4��$��'��"L17�F|k#�mLu��x�Fs2�uq�c������6?���f�e�Y/_��B��ﲘ��`@��&���'a"�doZ� �o�3�@�~�x.���qa�������2�KB��j����|�W,caBm�T�K\6T3���0a�K��(G�-Y��o���

e;��q�L`��~�x	���T���ܛ�{.���y�z���(	��*���V��Y����<{�c����n7�(YU��a�"FS|�Y��d�����n6����K1�Z �9a��W���k��L #���mm�A5����@]w����g��/KwZ-t��gjrj	��j�5ӧ6�OfmPXQiR6.�Y'��B��y��M�=p�eEM� -g��ڧw��(,�� �.�c���D��T=�s�T�F �\M
�qS�IG�
�g���H�� M���l���/���#I!�ؔQ�W�|	�AWY��w���,��j��t�M�S�*?���f~��)�ֈ}{E6O�1�>�b�R
�+���5,��]ʹc��H����%�+�������ȟ�*�q-A�S��{����%��&@�O�����Ƞ��LXGZ��ua㴜&J"8|op�rrыR ���G7��Ґ����z�uY>uZ����ˢ��jl@{*�g�[�EQ������𑵼��.)��Q����4$�?_������äi�5���~��s�����p������D��Ԑ��H�Y�B��'h_�w�����d�eZy��ymX`�Cj��k� ��g�M�jC���A��#�9ǳ��ʴ��5�7��l�ś�7�{��Y,ͦ�- ��G�����A_4��_���硩0�üP\�z�p�Փ`��e������тKW	`�h%p4��zs��{�X6Jޏ=t,�,K��ZS 
ˡ�Ix8�����ûs{zL�J%	LZ��8����ř[$�T�&֊4]c`�G��0PA'�p��%�-a�4�M����kv��K[��,~����r��Ў��?�C;�T~��K�ծC�I	����9v�*I0,h�?�JϚԠ�p+���'� @�n� ��n�4�G� ��^�S�	�C\5�'�����P�¾ݢ㺤�T�^mGg�Y�;�T���M�v��	B���)�a��/L�n4�������'��_GD�1l����fF��@,�@��at��;�#;�Dn�Y�l������el����#���+`�#�%��0��� 6�|ۦF|����p�f�W�w�V-���	��z�(-�=P�����G�&��G]�n���v��#��ڭ�m8������8ݮ!���D�$�����p��xi.�3jV{u�����ġ�;B��ض�vy[�I��H"�楓��=ʙZT�ve����r�a��u��`��>?��$dдr�F��w��ؔ9��h���ɟ�T�j�@�������z;M[�M�H��ꁂz"���ֶo�:l�Q�h�,��J�Ɂ���n�=q#u����Ud���8H�)��-h�;_W�E��.���(�'�I	1{�D�h
�(��A-�|�W��˹3֯��A�6T���߄"���:���!W� D@s]2�W|��8�.:��ᵗ)e��xW�������X�:,��mt4�v�j������C���Uflv�%�� 0����Ƌ��%`�Iy0��`l-��~�^6@�p��k1���K�.Nº�'�f�iC�t2��`v����S@$�C:�)��(=v
S\-`sMA�Q���p^�3��hbee��[� ��U���4� �E_�rq%�t��G3���Wh��v[��mY�_��݉f(!^�@'�֨��ĢI!���˷����l�Z��\f����]0]�� �BT�I�q[�:n��阇d�(�Z�s-�Ғ���<L�9pU��w˦�&��,%�X�zԮ���Ѳ6&�R�~�|`���!��W���-��.3�������.R�����	�����j��<���~��3�< ��T�3Ǭ�Z�{���eZy�.@�+H��X�l��@) 3�3�Hijc�����Y�qH�E6U�u��lK�3q��*�Go<��|�ѯ��E��IsNa����8�V4�k���"?�Ì�4�����0�H�5���2�#z����������G/�,�,� ���af{��Ca�|혶�0Ƹ��j`����*��>�}q��5�C��"�E������r����\3������n�)�N�4���Ec ���-�2�
z�p���>�H1�'�&T�S.�����e����A�"�-0V�/у�6���`u]�U�ȉ����l��ǔ.#�oiT�
�Ӓܑ/�-��2�̚�ݥ5s��$�}s\����7�㥏�j	��Y�m.�I�q�׿��&�b��d�����q��M\��h9PY4����4�+�Z%����Zu�CxE_���Kِ��X����<��9O:7�m�[�Gy�9�d.�$G���/�-'Dx�ڤ���Z-��aX*�w
!Fdo=�J�q�Fo	���u+A��̱҉����#B��HE�W�o��A�K\s�����9��K��L�YPHB;�qj&�. �
wA��� ���O婖b�}�cO�!��9c�OZ�()��o������]Vߑ���b#��~DU*��<��EP���#��ϭ�N��̢�ɄV�mo7��O���l�N�׈���u�^7�HJo��a;��m��w�7�Wx��jP�EN��<i���\i�0z:�dC̛�f�5,ب-DЫ��'��T�R�
E��$��������b���v0P˫UI���|�g���l	" ��47P�`=sRb�f�a+")��4Kb}24�g�l��T}V�,H���%��J�5��V�\�4�͢hrŻ�U�C���/��+�<Vj�U7D۽v��&�{A[��9XYIg�����[����[��(�6��K߿x1T��	���>F���{�m����r�g�]�4�ָ'���n��N"�^��6qo�x?�|���pI����F"|�ߏW�hl�7�D"j>/�c^�y��L�����멄��P$gN�L]r��T�i��R�{�n�5_��ك��&����i��o���ƍ�D7*8�������^؅�T���T��=�f��&]��C �w7.C5��;��8v%�SGp��[f'ЄH@
���;�t�: %�ֽP�������g�%?�-k{���r4.Lj����6�M�g�w�����ú$�&%�L�%y�q��W�(W��r�5���&45���*�l�W<8ۥ-��/�Rbs�������]m�S�c����hG�����0�Lg�'0T�K4��X"��V��3�Ŵ��]Q�t��VFmW��<���kj���L�0]��?,雄{H#�-��ڟ=$08D�F .�f��x�[$r}���r�v�} <�Rnh&K��ؤk����tȥ����RF�8��%��mX��b��	��D��|��E����>ٜ��`�i���Q�w�0V�s(^�]���+	t�߇ܽ̊�5�M���<���Dd]W�"�-��2 ܬ�3�,(a��M(�<���
�q�Ƞ����o�w8�|jO�K� >lߴ_Nq��;(5�1ٓ$����8�N��3n�~}>(Jc�Y�u��!!���B1��u���/u	8H��騣�Z霧v����jQ��'}6A ���H��c�'H[�IA6�����"n/cs}���ם�ٛ�{�wA:hIm�xC!��]�;��oP��k�v3s�6<6���J��q�+4͑#p�9�)�ľ�4Pݕ����z3;���Y8�D��?���znz���%�� �����x�1׋l�9���B��!>�*Zd��%_ ��xyHWڡ5��_����\'*����5g��J�Wp���nD��p`G�DCnO�<1�]�0�m��J�mL�~@�tN3�.s�@)����:���4
��|~~2��?��*H���A�tg�-�v6��Iٿ]�$Tb|����Z�����iϔH�8�v���l�Ճ�0JZ���	�|�٫��X+�j@�s%�	�q�.�Ϡ�����g�J�&>ĉ����imUj�@�����=���{r���{�l@-�E�jd,st5
��'�mr�v� �zF�E ꘄ�:�iq轠Ðpw8ϝ���C]�/o�ș�Dq�.9�/����F�@�C:�I	���~����ޜ}𼹈|7�u�߫���[9�r��/�ۘ^����x�	�N��j
p|�r0)}p�CN�X#@>���w�ҵPWM������I]�[X�Z��"�`d8�vĦ]'% s���Ғ����U�b�M	0��M�a� i�u�!�$���^P�����b�i�x~81���+��g�gE�TC�Meᔙ)�"����$��)�!I���ae���s�d&�ދw�P�un�ʲ.��
��6���l捘����1P� �yyڗ!����'�|>����z�`i��O;ȖGC�T�#��x��ۥ�q�����uG@2In�7��T({������T]�n�y�gO�2���ɽ�XeH�Wv���)W/�A^�(�U�ә�m�d
�g��ѱp]�j9U�9�ܼͰ���|����(�g�5�|i�mb������b�Υ@��"����C ��n�bϞG3~�ey�@]˰l���D�_����4A��}�Oz�$�O��P�غ�Kx�d�6�4Gr����xa시u�C�F7�S���������A$"+��k��n7��3�T�!�6BR��q2�q�h��22�L��jx~`_�?V�L���H[���K�Ș��g�%���$�q8*0Ռ�i���CQEX��Ky����1˸l���Ԩ�?/�#���������kP��#m�<~_P�X�[�꣸¦���K�YD�5R&z!d ��5��:o6�U�ΐ�q�L�<��m�XyR���,��1`Wh����U���ǥv���O�s���[�����t��tf\H^}N�%���D��\@[5H/�F��ru	�q�$��2F�� ��/~�j�a�lk0+%n����9ڇ0����oI���p/��[���3ˬ�,������$"���(!|CP�y��i�$:̌�˹��;~ӝu�[�j"^N��řW�������#�^�r�%�����g��'ji�g�o�iڏґ5y��@�Ӗ{BAk��C)�5��F:�>u`�;)&�B�D�w��/�u�k���j`��Ї�E'�`��*T���G���z�ȳ~ݶ D/md�� � jv��(�;���2H(]t�O��CAz�YS�3c�1n��gD*�h���#��ѴV"U������r�(Û�>�Pbbh�+�$����{��"�4E@y���U��N]|�r/�i{�(�D�g^����hc=�}A�U�b
H��]�-lc ��?Pv�qj.~�߈�̼���@�
�/a����~/�cd����w�˄����TB��My��Ŷ�?)���e��W�����Ga^���X��N���z�l�n}���O��Vi���4����Yӟ�ï��
�$w�~���EB��� �� ڹ8c���ȩ-���J ��\����p�h��#�����7�[;��dD;R~eb��Z`�"�.�{=��l+(�z��ۧ	��s`�J��3��xE�s�q:~*0�1lMq��+,��T�{|vj�����h�X��m�!5���7��7 �1kfn�$t��[�(T�.?=�4���.�A�T[\���(�A6(5�4�Sk@nV��k��&	�u@3�-���kjf"I	�M���_�:|�Ï���h6� �L��Bn��ϵ�?S�+0�
+�����w�kq����r=�raV��d��������Y��Qr[��g#�ڔ?!7�T�JG��O�� �F(	r�#��)�~J�����n���uK:aq��̌	7��c���$��{��[�pDbl��k�a��VE���\��u�v��B��^c��K��7��x�ʥ[�zv̝W�l�	���x���H��jI0�;&�4��w�>�!>�3��y���V9�i� `��a������̏Ђ���A=��)�����O��V�MI�Q���~�+�ₔ�oF/���4n�����nr?Z("d��l�!O�{�=g4����e�H土��=����ο>̷P$=ˤ���F��D���$�A��h�:.�>�,6�&�!F - �t�+�l�/�lnQZT_^j�KM�W�)�~PP��>]�$�ZY'(�
�yfƱ��;�v�I��,�H?LP�gv��a�igmP��'=1Ԑy�Ͻ���Ԋ7��7~����A��BV�>h�v���NP�n�p}M�p��\��`�QMȰ���T�Q܃9QX��@�{�[�e�*&V��˺n�,��"*x��5��Ǌ#JI-�D��F��n�p�`Y:#�G|��-P+�oPi"�׃��p��W��&�Xn�8�>FWUЖ�>A��!C��U2�h;qW<�v������<s�/3��A �E�aj�:(���� q��Dh0l�yԪs����$�D!F~�Y����~/Lxs���6��<
�ɶ	N��牾��;�����kC�f��?P�,O���N�?}A�t���;�)���Sc��Dln���4�NX1�L�J�.�*�\zpp���3I���1��k�֩(����H��L�3̯C����0Zq|oh�B�,1_Q�v�����rsZ� ā�@�!��#���;�`c�XD�#�A;��7��9��Q�gU��EQ\��j!Ťy�+�� �f��b������:\��ZD�`�=�G����)���r�P�U=�n\L2��%�U)�:Y�<]	"S�<�,�,�C��6�pcdg�t�����i�R8s��g��J� {��ԅ���t/ '�&�!߬�>��Ќ�ky�aU���ƕB���{�����#:L���6���yƿ�j��F|?Um�;���p����B�	��w-X!~�6=�زNP���t`��S�fn�I��|M:�(�͙H���bL{>A}iзG�P�]�a�9�X���??�R�|.J������y?��Ű;8�cOα�uju�oju���� t$�}ia"ELԯ�h��ͯ�d�e�C������4���>���-	$��N�"^#�N ,�9�?|�L�j���,�;^glD�>���|ܓЈ�v��+`�����
���;����=�)b�����"L_�&I%�9LR5"��b��{O v1$��2-#&r0o�w�θ�>[6�c�����/��J�%8�5����0G; P���O��k�����;�q�ق���膂v`�H��J��?���5�
̜��H�l7�`���F�c��/x��O���-{��:�d$�5'����?���p:�1:�PTR��tv��R
�j}O���Kc}s`U���Au�!3�Qj�~�I"���(� ME�I�>%����e��KWy���k���i[�e�K�@�J��ʮ��C����@:������Ȣ7�d'pg(�
 ?4�����.�c��U�����)�p�]�?BH�sd"8�}��ˊ�|� �2��w%�՞���'�����+�`t�� ��Xw�����4�b��qc5s}M��n�AG1v+�Q{���\��&g�}��ԬS�&5�T�v!~	��fMύc�X ��fP�36�zW��CVk��a��K3�	�
Q��P�L�>*V!�@�	Z���Y�!,I}��D��5��F����p,~�Db&���le���cSe�X3FeT�vz�l.�1�Y�ru[�[��?D����ܲ��N�6�<��(�H���K�� k����CngJ̈́?�;g���� D��錶w4Y��p%���b��wr1>y����Q��42�ͱ`o��3��2�Or����/���%n"7B����P �q]�rs���~/9�}��;.�DKMN�Vy��l}5:j�Z�j,�]�A�Ă&�8�Zˢۇ��j ell��X�υ��ZɅez��ΌO�e^5mH���2J��,lO�C<��@X���.z�=��4ۮo'����谫^7��?�:�_���fb����C�˜J��: ���.�X��^H����3R\o�0w6��ƪ��6%&� _ZZ�D�֒���I)'1���5�I��n�\Ƶ& O�$�k2(���<97�j<�h��+�=FK!NLG�ۓ�rqh�->hGu��;Ow�G6�@��Ȟ<�.>>��Xf��Ng	����*IFq�;��y�q��8����E�@���7Q;?��A�(��<n��ϑ%�-��P�+�]t$/�����Mlk�x|3�H׆��z	�2��q+���m � �����?bԞ6��Q�W[M�y���3�fRo�pF\��t�%:g�I�o�4�#�sf9Ʉ�x��"vŘ��Į�'�xKB/$|����Z��,�έBII�<��k o\k9��`��vZ/���t����j�j����x�9KR�_h�?�^���>�Bס�k����Z�AQ�����ͦfڋ��7�Y���W��=Y4�r?�/_�ux���̽��b��S&���߭��W�X"��*>�m��ȯM�b{٬�0R6�p�T�I���2&�(Z��L5?�ߞƝ�C�j�I���%�gйo��]�C�q�Y������,��ˇd6�P��$L��Le�,�H;�F�L�"P�{���<A�N���6�fN����[0�aG�ݶ��[L�:F�븥<�=쟘&��(u�<�4M�3/��*�6wN	���7�L���0��w����h�6A���/�q�m�r;z|QI����ނ�����h�nǒp�u��0�W�6f�Q*��͐F�'dYI{��_� �sԸ�z��;�_��Q����uJҠQ0�W�_�"l*S�p
������]�&n�n�[��x]r��g-��2������5~�2?���h)��Y���!52k�E�>Q:[J�!�g8w��>W�s=���g�gYܕ��UBӟ����<�&]gCKԸ�$=~$Gᜋ
�G:9�����w`���L���"		����q<�q�TO��Sb6�0�p��.��3!8Rƛ����^f�6��ܑ��PhTT����&+q6ĩnn7��@0LCsy|�A��q�ϥ?L��ަ����܊�ʟ�-����ysq���{�*a7�&��$B��v3�e�wf��oP4��ݫՙ&O뢩,�磪�,�l�#�r]0�	 K�[i">�U�H�y����R�"��v򹩰!o5
�)�I�<�4�Cǁ]P�uŦݴ��CM&�[7��q��^�5��܉Xs��I(G��f�=GS	�Ծ�}ʼ>fm�:�C��K"�A8���T2��
l�`�5`I�p�\��"��M���KP�f֔fV?�
�u���oU�xU��*�$�ٲ�
ν��ʆmߠ:��/��E�v��b��t����h�����+ª�]q9��?�C��Mh��J�?�������S���wP���&5y��<���#�7R��ҥB�71ۏu�fE�>�{%�F���/�; =���#	�?(�.��� ����Fe����1;d㫔�����H��ȶ2s�\i],�iNͽg���jL�����%/�2
o�pv��ix-�����)�tT��w�:"�	�V�t�V�N����Ϟ����o�� ��� !���y���P���K�S= oB-����P�d���2��"��"�xF(��7�j�߽r����C��L�Lo�o�:����֩\w�����I3V�$�m�!������I�HI�-Z����<(��HJ�EgMG��usviz#�A�=RP5����-:�A���T�	JT�$�V)��:�S`�2�쯸`��R�/{(��e��9
qw�kIg�� ��*V@Y}���T��g4j����PH��9�[���=�qlr�{�&�� )L�#������+�$g��K��;���@*{�࿙X������l��;9�϶�a%�>�,�r>�3�`{<f��ftp�h���,ISK�nN'�NTHO&Z�H��<:�Ӱ���E�ۚ�3N�0�j7��&���0�#�� ��O�B��柊�l)�cXE_�K#LMo ������b�B����O�K�~�0�Hu��c`�g#s�"��-���\�<�!
V��<�#<F����d۳Cܗe�h��͢X�g�6M�� ��?9��C�Ěث��̕��$�^�T_'(�t�5�/����R�
�Q����
��l6�l��z�����&[S�j]�^��o��O�
,2��9�f.Ԡ��^MU��=�b{�С�sj�Ì���b�%�U�w�u�����
��
���2��}	���e�"���4�U��7�G�4�7>4���!N�+���d�MO3�0���6���Gw��y$	��Q3�<؃&�	���G��9�n��4Ϻ��*�UEu��d�6�b�����%ta[\��(ZO�&iH�簻{��>�S�d�5l�GW���|hs�0��)b����_���[k�>�蕘Jt��>�����Ã�:	��}����1��!�H���)�ݭ�x��,!�IVE�Cx�&����G�x9�8����F6���R=����9ᒞ͆�����';�?�2���i=,���X��(�#�o���p@X���5Q�7����sl�n/�{��df�7В���)�+�}�"�Er��/�����#Y.���G�ϧ+�Zw�Q¼4�Kf+�|&���LW*h�tkX����"I�_�Oo��O�rȢ5��&s@D���i�4vH"��Dao�m����]����Ĭ�(#��Yo#9�b̵P��Ү����<=n����F�jN�@~�|3�������mA���O<f8�Q�150�V9/�����#U���K*�1"�-�Ĳ�K�i�2 p�hlJ9������#�|%��<��N�y����C��N����<���LƠ���z�E,輂���r�?�J��ʾ�&ZgZ����/.�Qw;��$+��֗o��R��~���ib��SR,�$�RE�M�c�3��:����m��/�IzK������I�y�Pe3�Iɍ�(\F�n�)��%�_F��⛞
À�	}�eе�1�'gSL�������9ՙ8N�!�.�A�	Vj�,dyF�~9�_�Qr�V�2r>&���*�%����R��$��?�{��{fkm+����e@�V's�-*Ӂ� [��yU+^�lr
�&$�|,�$�a�K}V���d|��i�wGq��͔�/�P�o�q�I��`�D�ɺ��٧�ZT��w��o��B����o����nmS2���*�{*��"o���F�����I4z����	�L� {�4Tk��\7���QO�>��!�-�[aKr���S�p~륒rS��ē!ts�ڟ>�M��:"�?V���ͯ|��ׄh�TF�$$�7"�8��(#���ȁ�-I��jQ�*��1wl����U#��21�Њf����Hz�Ӗ�k���n�%�c����FY
�Ň]Lնw��"T��?"��ʣ�JQ[��H{ڥ���[Wb�C�0Խ����B�i/>:Y��b�=j�}N���c!����_cq���.� B^�Ӕ�,�͔Գ9K�J��y`fo�����VE�=�IW��2����B9V�B�0������9d�֕
��H�k��&pe4K�k�U�>��ڻ'QLg辙oL��%�$�g�d��oK�� �9�T&��Q��'�[�b�m
n����C��~`���9�B��[2Q��Hon�P?��A�z���LZy*&muQN{w��JL�G&�FK������W�"�P횺泚=�#C}�8g�o#��&�L�.l��V���k����$}�`G������0;�!��!�.X�@f��q����h�X/ :��,�?�ܤ��ߔV��P�<ᨢtj]y�6���)�yY�(�[�&y������bq�<�xC��������Kg��TN��p�k�#�|��P���Z�c�#D`��8�M���AO��UH���v~u��O0p0B�`�)b��1ۓ��O�����������|��}^��*u�\��Ƕ�$T1-̚�e��^�4��<�+�-��`��5�`�Ř��D�7YdS!7<��ʿA���O	�?�<���Gp��͠N��HZy�o�K�Jz��V��D�z��RIc�fiˀM4nup�u�1���^A�(�t��q_�&	/&����/�U�#�zE[(i�
�ɷ�Ag�F*%������G��fB34v�`M�w�F9HF�����$;=������aTi�E�)���٩[�6.�_6��)�i�v��uH����E#f��o{{�3��@��3�~=�m6y;P*Ǯm��L���`(N֒����fP������}��j̎�'����#�N��\Z�����1��Ky�p�4{� ƪ❎w�D���T�L��P�Mjn%��&|�H�K@C꘰h�2��$�nW1�Trn�d��LC`|X�W
����^\P��m]S�r�6.C�j� �)_W��	A֌4q�WN��= ��85��8A�u	[�?E�b
H-�}C ���ʵ��n1d�C�������K�z0����@�1�w9S�e����J
/8e�xڥecɿx,�i@WG֖4����V`M�R
�X�}�p���4~���#�y�|�Q�9��>�	HK2�lח�l-�Y��ap:�������y�)��]'��0LSk_�ai��q�"W5�>���VG�@���?,s��Q�97�xX-r�1�0� nƻ�t-�g������Y�����O'���U{��M���V�E��*��#%��{�gc0a�1� ��ɟc(͒���f���=v<�;�r0O�'��?;��;��j:V���\��VNG,g��b�Y��ݖ�1�`��6rj6tb����Y�Ji��|e����T|��)���1u^*�p�Aq��e��f8)1����d�ȕ������"E��-�-���_��$�H��{��p�?%-F��,F�6(�̭�R ��;{�"�tKאreߤ�S��H�**�=A�_�nX�6e� 7��;slT�R5�?]ìb��~����4s��Ȍ�I�@E=�OYR؅8��&��ޱ$��tPiWJ|���*�'�}��$O���GY���g/;l*���";�݊C�e�W#*xz��]�)Rs#Y	�q[�c�%�! :$:�/���O(��ܞ�/�Sɟ�/䫳�!C@�a14��:b���b��NJ�!M�K]:�[�ŏ�&�z2IU�I���k�����Y�k��a�:=��w$�u6��9��:|�+�(s��QB������� �?�EHgs��؞�}<��	�&?�Z�bz�uV�a{��ЌAߎ6��?�<�1b��2���SR��gɔoA�vG{��V,g�\a��,��@�}	� K��Ц߆�E���J�D�P
��Q�Ce���B%�}�t��H*�nT��*��,I��m���D���}��N�d��I��H��˗.KT��z�X.$�� ~�HD� ��{�	K���^�-z��#W����	s�;0��Ԕ��PLÌ���.K,����w<�����"~�@a�є��%9)^�=����p�"5ic�]�(�6T1�n�n�z�k��b��}���5T�4A۲9w�=u���	�|R�J����+��Q�2g��G��:��N��PF�3�>ω�$��J���
1"���L�u)��P���3�F��m�ZD�Ңw��ް��"U�m+��o#��!�/�Q~h[��̡�+D
�G�do_�B^��t�_�/�0'��|0*��J�Ew:C=�Lk_�Z��ŉn�=o�a��'+��Z��8�mZu��A�W��۰<a�(c�5e@��Aۉ���"��@��0E`�V��q���D"��Y*W��؍��hԊj�{X�;!�>R�1<�0�.Z�Gܡ=z��e�<Y/`�&��Ik�*L�Y��db�H��:�](ZaRR2���((�H0�Ȩm�:�` �'_��I�H ��i�?Pݔ�تuB���6�'AX�P��1�$l"�=}sn���3�?
�E�ԛ
�`.���c�ϣ�?Zw����e��We�����!
qL��|��G��Y��	a�p-��ق�~�P9}�m� ��a����8'����i����J��{-�����`���bk�9a�]q�X|P!RFGI�xJ��-7VԌ�^/ق8��Q�N�O!܋��X�.�IMi� C���v��]*��j�PHC}�"���J����E11RB�����S�Y�T����l
�2��`��}[� ��0��T!I���)��Y�����I�o^���EO��tr���C!�5��wFՆJYA:��Dv�/.Ӹ��!��=�0P�o�-�͎j�K��T��(H�L�pt���i᷼O�‚)8�"� ����Tɡ+u�\"����#���k&�{yO��}�J2�b����*p�� �_�ߩ~���a�G����v�g>*j��R��y9�T
ڊڀ,E�?�O�y�7$�Hq�ݴ���v*����������WQ��Q��1e�?/�F�8��{8���ͬ�p��n76�h(�m$t�G�ч!��ӑWT�^qv�*�q���F9
D�N�1�|���P��a��/\�J��(��_��B�4��.���