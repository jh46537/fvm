// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:43:41 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qZiglUi8We+YW+PhGCueu40uXuZs+ZuS6YBgVxGiDUFV2am/hxltjEx8204gKWRv
xkK/eEF2n5Kf6QD0Y2GLHq2/6s4ZT2U1zoAuxQOluFBcFTiqoF61n7AJYYEw3F/K
7BxnigvHiiZ9rtXUnUsJYRSZGqyFqI3G43dgnR3cvj4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26016)
h3H6F/dPycGgy442LqMp43FJ4bv3iqiBdm9Gadg++vormSSoyqJ93veLtgcFKCTY
tP3Bu63uvo2n6rUndKkvQ9lcSQCe8zN7ZOL0rICKpDjPcQYlun3trQcH66gcmrdK
fYkNtZcKDdPjVm/yCNRVAsDkSPfQ1hRAaB98eKM5G+FTXbkwiMoosl60y8N5Aaf5
CHWkyk4CIGOo07gDcsQfndIlakdns/yjqyaRCXKccM14xgjyJCFzcOThUQqjcES3
EF4VpSNdPpOPxiyFHRc2mL1zSrLwOCAX3O0JX6hAQXt25MUHh5eZwOuH+Io4/pUb
lBaa0MqnSqUMtbeGn14aKLakWfg84/JB1IR4U4ZNJdWO4s5N7+aZ5LmCmHAljc9S
PhhFzc9SH2HS6eVdNRowYkKC2UJLGMIHtemg0NNRG4g4bAjSyG3Td79qBRWGkHsD
tq0HQZ6e+eu73m3aQ2gSjbOk1yz2+ILllxqObxQx9TsNfNjhEMwazXAEzMS/Y7qK
kI3hHMheaz56nv86SDnSiREVbNNfIeASDkNfSnbKlOiP8U9jctLl0PIMtwA1k7K1
bcfOi08WHEOdGePaoQOF7cjIScwPyrDmiHjZTSiNLrXh34Jc2wd401szn+2FAFnc
Plef5yF6xIbeCE4e9sVu+2ycwXFMqfS0IgkYaS/WWlQusaHBDfTJBL7L7bDFBwtQ
R8+THRvisK3sZIBS3RMhfmEsuSfr3VRM6rqjDJORQtqKrOheaHM2p8c4d2SIY30E
gXWN8aDESMRIk6DVOAhlp5r4Sdwsgn9B8USl+w7xvPaWCPnB/IVH8HJhj2UhroXt
yuEIPwq3kCo0tkBBcFuow1oundAkZqL+b2xaFkDK4AlOzbLS8LMay+xiZWf3dBS2
n9jJ4bwuyZBXFD3Dfl5C7cGgzBbN4g7C6Fvsprfr2Jns4d4H2Xnxg+hFCW+d2Uwt
CdQPzw1K3+Q+QeE2K0G7JrB+Skqbm6ukv1C6/0DxqnDy+t9oiqhEzmfGIaPzpN77
7H1oAEn/95LYkZLuAYYHF41py6Bb803JvAtLm7Pp7qBpRTZbZPgi9VnFnTM0joLD
yenpey8yd11LfNUGghxxIafCtVSfbO+VRIOeLHpmIcSn/8l/9m4oUlYcg3JH4/5r
Sc6+uXbXgjryWg4kS56cOkPD5MyjUQAYm3PF2Xm7XAJY3+9LkqSK6f892w3nM12K
YmFW8JRFMr6kfRYomCF3s17XxyMt7+7SfXzLuXJIPKD6Rb+uCuHxuQ6nxoMLJRLz
NocPwlyYe1+kHEL2Zgf3FaM8ZJmfbYxWZ6jErvXzLKZQzY8vQPH9DwgQJ6pz5RGp
7GuBJF8x3+SgCkf0ng91Th0fGBeUjJLoIY/CgZ+ToSqqjZAQaqKq6xXiDuHv0Cd3
pjg7EeXBjVZKJPyCskB4CkyNbs0sBvsJPd/+E6NHOZhFes0dSjZrJM22YWWF1y4m
sJFSWn/e3rx15eghnoT4VWGCjuK7Fbn70tKRZMRBdxkibqUnF72S3O3nd4attctO
8QLkuISN0R0dQkrFxiWVAdkrZvfdDAXZcAsW0uOGNlQREfgLSOVmhi8oJCljI4ya
2zrf8cLs0K6CakWASpw6kfeYpMhUN51VV8Q+BC4zdHYDdcguy9ffBEgQ9o2zA+K9
BJ/2+h+0pICyZUqwjvntwzB0zMUfPuETL9zdpYsDgAOiGQ1v6PZJi9BSYQjP+ahN
q/Pg0uZtOCgKpW8w+syEqscVcwxNPF/qZKWNzcd/M3cKvoHpEknOEGZaNSn3N9mR
NNH63jhqOWtzg2daucLspBsa61U+eH5rB1Tg8qydQquC5ws5mCCxi/jgbU7su+mh
jvXkqBqU6h2utlgUiSQ7Rt0TP3XrFrw+NLxIiDrFupYzQgmsR6+W0cSdmsK8Of52
jDqd50TPR/Qg5YvHOciHvxQoQoHvm0G8fHkaWVHkPkwZu6Sy7OFj9GmTXG4D0kFg
+pfqJzK61bNdIhMKsHnp16lYNPzBy1l5WQGswJdE1VUfTq1D8BIrSaqaSUffuIz3
PgvARVA4gFdjf+xE9KO15OxFArxkcO2FNgzQQfWCJiwYSI6ArIroNcfQCK3j/L2O
JdRHs/CZtM7Lzxl81ogI1zDnMfaph7LHrGqLWbmFDugSLCXTxHxx0L2j8mThQCrA
/9MGGjmPoWfQ7hKCL8rZtoG2J0U9t3MdMeuKfUsO0ZAkyZuk1bydhNp28wNKWUbR
bptb4h4Dkpk1v8yegoawVrMEL+T4wsXZL5z6HaBNe+uoLafjtrli9QTse3Jy9vZK
DNLEkAshp7Uvf2l6a1sqQXQhdUdJB26LplBImj07Oc3yco4nNXIUlles/J7SZbZ+
3pij9rhLxbP+ocsraXH3mm/MJjMfkYDZ31apl5ihnSGhX/P5EWBafUHSEZvyP2nq
7zCVY4RNSkMP8a58Gx3Uq6p4M63XhQe/WZFiblRsVXzRO37P7F4rjcmeShSf/Ix6
ItpojbdXxyi9dF+7EEun6YJHOrBVWOO6yAHUGyE+6IBsLsSr5dLAOyEPVCAD/RIW
5erLaHOApczbspnQB2dlwUKgyuNeShYuuyXCOvQmNUtLCMlq+pmQUqo4EOChM91k
Rg2YZ3Ckq4CYrDjDjZIJRpvpS7owPaVfAzCbve9MVlSlgKUnGkc27WdB9EfWVeYb
84LsyX1t1R5jctzSt4ts6iKnj2zSFHpQVqOAo3eRuh214jGLaFB3bX7ontgC+G/h
vDh2DFQfHzvd4Gutq6DyDmqYbHGm+K2VYGXCSDF5OwPjbwn4Pi16NwGOHUTF7MY2
vE5700u6rzZ9P2l5KSU2cfKMzC/LhgLGPy57mzBWlrXfxNqYBPFwgr3lxkDIhNAU
1QQyc4frb5a/Ko9tudJEDnZ3eSugNGxeWaVV5ZkcgpELTo6Yw9OyBht7zGl35Gyg
YCqIeaVYiW+xOljiJUYPPmMSufonQXFc59ohYXteUQ98PoQ4N7pOtL2BNEy7iAxB
0ISF4cIaICzymYfOTdHc6l+PqildFVPvmSZvPsb/ky3s2EChJh7Pw6bJ6kxxoPYN
iQMoKW8qx2gMrpRPqX+DuCO9rRMal5Tncc3eeI9dR4/iByXxIeTmc6ZLl7BL19YR
Y0J422eSSbzZChnzppKhChSsYf9rNvMFs6lnpPB6o5sWN97VIJvdsPAvBQz/lt6C
N6mLMy8EkDvkNRzGiw4PDqpGJll1eMALxMH2vhQZOiRIBkQ4eplMbjGFZk1Ov0FH
i2sPEczB1SUxC0gVaJQN65eJJoGmiatMTn53joNOEdFIM5ZnWfZqxKy70XqmfAfZ
gI9ZSTrhQXIWdRPe8VpBzHvxFG17tiDP87qaMcoyJYVJ7Yn7XuXbWXNaktLpfTux
4KrcI9Hifnme2AZtsVqBg5wPV44pUil+zSGkrNKknJ3tAvsSEz2qdT19+pDyDTRs
AyophHugHcvpV6cW/nWjEMVQGt+4B41pxDgoGtJgJ4fsrbRP187+c5r1Is/UC+/t
30wgFSrg3r+jBYJWXRiZKN/iWvqXIEgbzdC88bfheEuSoS5POlEj0hU2GAOBz//R
PIyQxTzJOXDRYT5ISFo3Pn42zK2H6dp1wCScuISo41ktXaOlUz3l0vhTS6gs0azt
x3CHEO7E9xiTO8kzi5THRo1ANjNgqKS7f5ZQRIEIBUdjIvu2EboVgVq9EoONW8lq
Qj3M63/2+t0tNXyfOIt7cjZbbYLnSwV95W/H7OwZxrFOGsnhsIphP5QwGXK1g68f
Whw0IRVnNn9JOPAqX6ALhXLvfrEXgHbUe5sHQDNwnIQSI5vfJdruq3SyjKe4dyFY
0+8ty1lwpIXdsf65rKjDe/UHUIa6havm4fyTZ626fI6piXpWBT5JZi0EnOiNgjnI
6lj5cVnWgSeU6r3KPNV0mLXGgfaOMDjdbabs9iWftq1XSTET22nChS6OANZExc3f
299DE12Tsz9iPl75vJrRCbWIdUDJXxfDhxsstx+6ME7Z4z6wgFlTLfft+OZNOr71
pB5P53rh/skGGDCZji9HtLCrGgD7bxA3FU7OHp8+/dOfp2EvmNKk0MOx9ghU/bjF
AC3eH4yncdHy6D0aMA8PPKkqh1cqHmE5lvcPqF6bfoJOgdJ5siMMqEsc4MUcjCnJ
9P4fy2HSZuBZzZhyD+1JM6pwYUiUak4g7ctIUurUIfoSpGa16Rr63zZrzih+jmJJ
wlA4vokVGJLJszxj2W4yTbcsNYW6zVGWL6lMaOpowHpG2Yaisj0to1bKoYRRa3PE
TUN8wanvYGsv/EOh/tLnh1++Jo9FQkgqw8ZYD1xxAAuj6Lcefm8xbY0NKDEyjN/j
Xvy7GTeB6J9fQSfnwaAypkycg3ITV4aFNqeMO6U8usB4odxqRHoExXd9xuTHjsIl
M2RGvCprp/0Xnx3RoweQRkad/jBBBOK2Oq9HSuDqXt829MwVHYeSjzA+MIZwfT00
pNYCTusbuTtu0vkltYgdoebOLVxAQJesqV+QepJX7jRbUOogfkC/cU8uWnmlGPkV
/kNukvE82CLvrkzUA9t4QCYKabt/Vf+bpaPM5mmfb+WXf4ZJO7b42IlEZn3WK3xC
W45iUJtjIkuuoK/GUjIC+xKfz1pfQM8Ef1bPQTEQOYjqs2uAM9BtGwy+HBz2RWkY
ZMwMtkccQ+Sk5qmThFKd8fEC8JNw/zkkDN7QI7g70y1s4zw9VIyeJq8fnxezTlIV
oJshXF01IvyhzFADNk1wYos2vLi/KXJuRWStE4mPA0xGa8f1Q98mMJyvdSFA1qUa
GTLl4Tjq7tYPzWz3qoJzfCnbMQ7ecElg7/pu9wkEiZUuwHH9zI2yrUETzJjAFidz
ISbPOT35GlgUMClfkGd84ukNTaJ3u/s9knwUaDzX6LpYiFXcZ5t6a+IWSy7zKE+D
GZOStO9YwQwp2pE1qvMVkVw7jsAsb6zClxnzorRSxcN1AioYqYQLWBKPSwqCIIox
kIC6DCOdhSczMDDBZk5T0XeZqtsF1t1mpY/FTIzvVEJ0eIyYn82msFIoAxyjCeUP
c5pBMulk1Cr8EP+i5VGGCzAKF4R/9WooU+AVOMVrUglWtQ8pJ586u8hRIEED4Sln
6taGab0JKPaHctA5S+UbVgGt49t3vgZ/NTKQ8Hs/pVg90J1zh6KBf+jsAxkmJl+n
J/6iNJE+/EIi6MERFM4UZH8zLt+2/f2GtakhPKsGuuyW+Yh2y8JBcfCIR1oYTG0F
ZbAg+SkOpF3WpiM/g5BwwEb98BNgrvUWictBBeZpUEUztyKW0DhujlD35RSSqK5B
quXjW+TFElmme5VaqXySvqi6aDbuGDzUt00LJD+wubgWSJEZBxgz3Ed6x4kJ8BKS
g0TVzY5XcLHHe3YkfbhA1KlovHmchZmb4l8qOwWr0GeOreLujYmybcqofVpn+8LK
9UnPVeDe5ybUA3uzFQjFEHZ2tgtRb9DE8teHGnWxgJ71km1rd7o9gwABrQmjL1cw
xvNkPEl0ZT4SO0I8lYLA03jaSxOMRCsNCEAqCCWvunMHNgjlN+BgoSbCl4PPKXeF
tJn/YNI+osXt8oehxAQPm5fDzFRQMe9zMfoRcqdc5uFK6u4gDNVL8WUA4YRGvH60
E419NZguzpuNS7E6X2ZDfmIPDShrUPwfx/qHLt0ZxcE266So6wlXaWWnvQDydmdd
1kOMGrWEuCyswD0XGhHqVi1IqbOjPdwgrpldyb6OawgU5rczTFUzsmc8RTYa41d+
y7PaKTHn5oFjveoWHc60bxVYov6MKNLV3pXM2xwTfsE2dt2ac51Hh3pWGpvboJuP
SJJmnqAMA12TDLwD65uVvTW1EW7hOzkdCUOK1BIz0R5H62BIsS7/nLilJHCcAAeq
68evC8zDMbNUdWDaxHON00LYUVpwvfESN5hp5ejNGyuZNAgqpMPypX8Ub0jkjGOI
DtuU4WArhVukVMUdZspddWvX4tIDGLxdS8rUa5SN5G1XGh4hv9zJQXhbBKVrFUBz
Sl1/D47O5BHUXCXeaRyDfQYmEG4myw+YBYq4d+qINpE1z9MEg8vrjHuTJz0R7PkD
mTW3pAczA+jXYpB74LpjdjKkN7xMAe9Kp3R/hhxFauAjEnQUhUpVAEuaN8U6mjD2
JUkkJEHA2/PzBPz4m9rC7OzjcwIwSgyLBPcC3AEjJTBkUaOvAlt6kF0Q+Qu0ZRrM
6/S2kb2kJkUQfiDdFploKjJOPjULaPG9qzejOK36SE6wk2Z7vzkzQMrZ7IdaZail
IkKb4BbFWIfiKZuBuIUHmfkVR88PlMu+tgbFRCOOZCdVK9/+pHvlQCYfQpQo0jEE
Duxk4R5IBPE0NQGNUB2m+As8IokKTzRXXgmfrJVjSAQS4UGczi4/X5+ZjGZV/XfL
OFnKdUA/PfVtVi99JyJucT85gwMBMXtf17fXDnUWdRLZnpT6PZrfaV/kUj1uSfjV
taQdZSRRdh6ZuuWn7omCu8Jrjesan2mPkttl+Oty+tlB1/96FRXNcVEwAa0cbIMB
WNk6NcsFUrH7RyB4dh0noedS/Q8+eOz7EiAgMGAWTYdpTckYcYcLOUYerQxu8rHq
NI1gaBoTwrsDPRTOvVo1dMavGYgLlSk1hiXMSHhQRU9O5vsMgpa6TDhSkcuYdB1d
dumQ+aP0W5jWh9ZB4fdmR2a11Kc9zefq+61ej8XMd04AieDBcv13gIwJnBqllkII
w5xfxqOlu/fQ/JAHLtHjR6l3E/f24vzEAh310tv3KBmxCTON6aE5toawOaLelfKA
yRVY1SWi/teK+wzXkgJcdb3ObXLCgHJmNyhwTbnfglHLjpPMQb7aSgp79gECxv4I
on7J3VKn+OsXRTu31bnmb2L+Uj1Gr7p3IwfHYf59AlzRleK/goVsTEzwS38r2wHL
wUQYVI9Qrf6sMqLhCnct0MJ2KV2I++9ErcDQ3xpwgiTNA3FdDtyFp8dfvyvotCOc
5ZmXTeN2K3vx4UExjBnRNB31ABh71frsQHjSJg/ETZVsx1uTLO3+tVjPQlyir2sX
bRTb9aWb9aQap1jDdVPECmbKnvcDYo6uxNPJn3eLHfAp7+m27x1TeyZePChGyxEc
j/Uj1zN4Ug23eeq4DQoBkiZiEJSsr4qooN0JoCPvRX3tsXS0CxeJAB340ayq3VQU
yMQgEWc3iHgvAw7s//7wAKnQjQ1bV1mNPtpAWYhknOx8ghkaPFnqAx3q4rHkOOSn
/jAMXeun2GsynvsqlNtQEzGHvKAdIa8xKZLqE3mxa6Vvx5qgVGsRfc+ZG0apfzfB
a130JjbBcFq/xbSdl/yvTUNiKKjqND0TPVr9jEiI5Z3BdOuRLKq+WZdf+0VBkNSG
9NWjN6gffW8CG+DBwVs0X6BXQGbw7J8CorXoIg689uAC4xwuYKtkJf36TARQ6aqA
9Gn4HDDqwQeqRIjP9IZMIsGW72/WCyynybHEs2C2ZBFqz5XJFM4Vzm2uurbTdBXO
+AbKgTd+iZfiTQdCViNwKLnz0G+BZAz9nxpRp23KvrLIrIvezbEceSdcFOP8ocmG
MafN9O9uAHGsUFLp9ybcs6gCTUATzLHlWnAML3ERoWrhi90gABRs9Pw8iRBrJ/PT
2K6NVmnHDz6nM7QVxg6Jpa01TUgh8ZdcGKU+J9OacBwtjpezpYIgvSI/j1dFFrAR
HsNR9TN8gxh1bby8rGV9Z+hr2/ORR+xytUIAKWfOpiqJLMq24GLppoR5TMqHYu0v
4Bom4oT/3JmJ6sHrLGvCdivWF+4bDIF97ECc85VV+LI0e4ylPWWd/m2WgNUFXChl
orw52JptjxcesZyG0Bsgqezx1RB+O4+KlI3IYuYkl+v3SQuYFlQqJBIeVoEYf9a6
HXDGLbtLqrFIFcHkksAjqiP5iVLsnrdokLLyvCP6XoKgzs03QVQhbTT0uS/w/0QL
YhWxz0FcwfhXWXDAqy1YS/OFwyVoXlNoYKStd/Wz4v1PcoRdGMmqanH0FZl3JAw7
hQ7LutUoTquS5JVaJrEEKiGV73JgipIiam+S1wgV6HM/Msl5pMsZh/a32zPAuHlO
dNMP+D/gHXmwk74NiB/thmSeRQIKFrCx7ZnUirNUk+EKz12eEwxLmw0DyO69y1UA
i8gE9VYUgglD3vbaRUjswUIiCGKU5Myc4IoP+RXeHBhJ+dzTaVd/40Y3MzyIzm4c
x1Bg4GQJ9JGEREqECYHFD2R1g4aVK7y7JFyRXqKy0XQu1QE3VVa1YKsYecwOf19n
p9Gg1CJxVhyvCXr6R7nisN7OhJOsnP1TFPPlYAuyvbXS5MyAkxi77Xg9SDhEqbtY
UuOSpomnusVt5AU9s+hXP2Ib3GzGxD8IQgrW1fQdG9MFwgUKMkFhdL6UF5W39fvD
1ZFAREtE/WuyTxS0V56/Im2N8+CtCs8ZD1EMI4eV1P2TRAUVhZXP8Yd9hPaeWiMB
eD3bB2D2dExfFdoHa2+Rbe0uMnmcGAYVGfYafVsO8DeZwbovLWiqRcaXATeDGNBZ
rRSTmA/iztKspTMCHDySpcMUj5hqKdfHtqFRN1lFopROtQdo4d8/AuAnTleAojOQ
fE5ypviLMcr1pqIyPvZop2BiCeAxZbB7gP85hNy2Rp5OOXLWXHwf5qPzFIInZOZH
76/bVWF1RTZea9o9y46u/Ygm5AEgCgS9Kt1z8mzeY4Tr0gLeUpcVFAn6YCBpydTu
JNFWwtAgM00ROYklaxHJ66irFnWMKR7haKbUQfiOzAI07JZ9yDSvaukIC1o6cHv+
WNdEvMO6ApgmaklGs0Wfr12xipDaD7xGJdr8hrA7xLdRXtiowalsBQNm4tTVXoZ7
keTchcpQv2LRqL5ebJdblyHqR+IYXpHUB4Z1vME6b3BWuYy3g2nKcye6Cw4nc7kn
4Rx4yy5B5g67/tbvoKCqOc7J+1BYZrf725eQ4sBBQJoM5G9fR1iORvZnoEjbtLq3
XliPBby61PuzYcFdEeP+i9GrTOplqF98FwghCJmvM/WBiIoWGot3BgCwd7F7Xg1e
2HfpMRVmcHvyH1hiV7RibdqRextd4gE0EK7y1HecWuIBT95bzimgb09z2bRXMiqX
0GHNHSEN8oWHixRE1GGwSb41Xvi7Q4V7nutbPe7v2C0NuL2ybc048s3MTB4X+etk
RJ4t/Uoq/3hOUqC2Lmrq+PY/PtCxD8Tmz84E1J9VpM06dqXNFobv6KM077Eb+9Ha
n4aROo0PGIe+25VYG2Kv+dRMOxI5RUzd5OWqzgUAUP1qDlawBNoQ8KDrvefqzIC+
nProCbySy1kF3Ha67FcqaU1RIr18PHeOpLkqO9ndSaW+iuZmHAtmTBh+Q/5pdTBc
tD8QLuYqIc4ATQ7Ik2sBzRiZIaJRu26YTlqlEsvl/yP6bfhpt4+g+pC3q2oPluF0
+9lYbyT1jOt0t1cDCuTHIvPNz+46mNrvEC+nk6amAz+2iSZWdSy9L01UOfhBggpv
DLjE7115TdTsLInR8qWdbhYXWvftI69dF/fSDfCemR8dxdfGzo+ytn0CUzVtMPyw
L1Lfsi+yl7eUHL+0kDDOgO8Y8d8ahDPuYQICfnVH/v5ZdMzqCz4OxeT0zqzx/nnH
uNHx8/un/wgwz3hOHMSs9wrlDzNwP7IvL3Y86miKT/shbUVYL1cOcoGPBY1fONN+
mJoTgmGT7hSwT1ewGrWeJeZOAgZOMaX7+d8b3OT5F2anzo6aXfmbQ0sUdMux5md2
PZv6ikvCOByyK2qL93drQPFXBKNX2YHGus9Una92WDglIqdldCgnuQoOL9GCe1E0
WZA9DvOqbnAmRJYYPiH3CEqC1xLlBbArzkEHXqZ90k/j3rDx4ow8rxQaZUL7E/Mw
ULdSGrZnOAJ6qErQE6OLacH1zlvUXbvhI8z/ay8fJkTXFZpczXqisIsjaFvEIYeS
h7kN163idx5eBkja1G8ImVmuWMdXE24hzDvP9XKe6YHHWUD9W+MijawTr5mLZPJG
SnjqUhVnDaoIBvLkaoIeq3dPB2fVZAhgobNoPaZIarGYT/AAuAgC1PydTwfVuejW
1/sK9DpggfNggtP6nuECDoKSwxvP9l9MZAxuM85g1tSzNarnmrsyLUFov8bEjbQT
6ebqpNJ4HrbFlxUjTTEEdPw0RsLjyzDDoY2yPURu61aL9b74tN/3Aq57/yfKFmvZ
J4yPFFr4LJ1bKHk1p+ux6JAjvQ61a5H+d6eQQtM/xBFi89PI8Z0PL8rl6cPQDPHE
SWdeu3jCZ4OU/C8RLgSD7uatlqdo2iPOtAGkrL0E9afWuuURIgEXsE2WwdnCDUw8
yrP4lvCX1BhyM2yV6hitKa9cJqurwedQNdfG5gxayHiyH6OLI4okcTIGbOVilebC
aSnLSHC8dVTm4HEa6v2Yau4k8SOx5HRo96LKMnjdrTtaus+QWgt1ifyoR4Co7KDP
t04COC06Bvu3SwNdQy/1D+nvavrR1c7jAsbmpFblxmo29NMdtT/pRW6tpg0t6ycy
VIrIU05d2pOii6+h96KtkgOkBLPNXe6RFBt5Dr8NX8fhGIZN9vcUYVTqNvVFvZT6
baFZTMCikSo7EKbEOdnAfwTp8S30x3QVNi8T1zB53tiGYbOJ0BmmqddMKNdOPBdk
KN08C1a6ElmCIUP+3VJrM66sa3wbRtP94tkJLxQQd54ITBuPQU5rVy8wZmko4tkv
AWHSE1AH65F3YS406MEr7kI2fBIuQTSYFxn0roD1iUSh0mUMscxBVl1VMAx8iCer
e4vuWKBK9k25EssHluQjq1vymH2yzCgg68EE9D3Ajx1aFUHp8tZC149eQeMGLzv4
GsdJcqZXg4R/uVfapeCsXb+u/g8i8mNw8wC0dO0yJHghvLAPRTcuaWVi+hGXLqSp
kbGXJoXBOBL4e3yn36t+pdgVUnvc1Yfrf+Yhxwt5PJv45ajA7y6MeJp6YXXNV8O5
MjWnFfgYWG8rItBuZV/ir9PLdfzWKu3O1gZ6QiyQcBMpv4HdtSXX3sYRG7q9uTyW
99eZzfUE7eHsYoVsRuFXt3IhLFYYaQ965ZZpNhbDHTr3phHIg06HE3n1dLGi1CPP
f+URZbMgB1gOL1IPVSv2Ry7vMf/VSz8A4A0SWkYT7TxLOOaWAVNtOIFuvyVQAyL2
F1sxM3/eKRAVJTQqWXa01ppSl/h8aOgsbtYO6lmdLHGiR9yfT5Ug3dnX7r1nw4Zz
Yt0dulEF1w1U2+bcnvNiJ84feHFq9MmiFmIuNspPl7B2SY/+GiRa1+ErW+OiyE26
x+r1zoC82NpNBebWG58FIzivAreeOSGKQ3VPhssLmbEaSYyJMHK1ykq1Gdp1ZcfM
Oqo6xjTcG1qwJzrQ3FKhlXXxzuIz6dFftHXAtBQw5gJR1yEOVeABGO1mOA5SdnAV
mxO7+jJN0CzECkVeQ7Vt4sWAHMe7RrOJS8MQRPR3a43eSQvtQ/qO3vnmlUDS3SkL
pNsTLRlvpURKEaBTjxscReVGOxoPijgCLo2T7ThjwtX5uNwFkLIl3UMov6civTuv
nFQwB45v+n8wnsec9jOt9PYTr/eCqAI0szLgA5eyBvGd+/ORt1Hpj4LWCwel2vno
+PJdP3cYkeLKw+hguiTS0KWmXW7XyUDNc+Ws0hFn9JzOYLBhX3vdk4VuvvYRBMzU
vpuJNncOacm9J108aGxNzfBm7jwLRMtQ3T2ONi/LS6S09Dh+iozO674xKVORz5Qm
VHg3qlOS492NkNiZSrbpvgP7hOf0yOxLWzkAK+S6X7Pkx1Z0C+o3Y2ntfQqWPybm
Rj11yn+EDV0Vw8qvHPdJaqVo5c1lr3qQpDhIkc/2mxMq8E6uo/EKkqo6Wqw0m85k
smoGM8ou3ERq6vkdGw+eHXetjZJWvt5MCnHRgH5hp/DVJdGBrtVSOSPQVhH2ngBA
teM1xvGgw1CLWn0r1qKLuGqCZLJyxxcHiIC6q413Pvh9NjzAQ3KM46Sb4j3pqTBh
+Y8NliKBU9x9RDQRM+rnFzikDFvjPQdS/9/SO7j438v1rUdUjhqbt7GT/qCSiiK/
2dKpieuq8yea8xOESQiMyix4V1s72IqORXgI37n7TWqaKZiajiDFYW7zOV1BVxd0
OBnCahGh2ho1BYOWQY9HBnUBDN0NGzOQkGq1V70EzTLOemwCgjC6b6qlMX8EdeIb
jAQ9cYwGhU/ylzkuOuUawWHJKfyGj5UuBrrDZVHH7jsmvC4USV+5CTcwjMpcAzEw
M5W0I2UrsVyDH1ar4BhBI2CAJDOx9Q7qEnDowfuvVCNTVXhsLbtBGCzp44fl1T7d
lFZFUmlWGGNfHKX3yJ5TNwBB6lbRye7hYQNd7gkaNoT/YRvypp0B2yO2gxo20Qc6
T8ka6xtmzOGkEeBRHRpAiI/XW8rn6LIWL6hFzoN4fvrQ2KgsD9B4PZU9IGqI0muE
q/a4ICSGc+av2GXHOWgw+ZOVZqJKDpXOz01sfS3Mbu0pyHfwxWJYEsJ0Jb1HAz3F
vPmw8sEVnouFRVkRg3TYopDux7GjdjKq5PSMk0HNfZvbOctMR8jZJvyP8aZDvOHT
ECdDvL8UU5quQ9oiBbHUmrZ4mvaVVCVjvVxGde+F0Fzg3JciagVwK6QrzBP6ssrk
naBYR0UPR3Fpi7hckJR9BaFexmilcy7hUGZWR9XS6TSZr5TRDP6d5oBw5tJJdRQy
YXCyBCUoUKXiUXLf1QWKMCupsK6IT3KvEfMrdcq4/kKTO/D7O/H2RCMZUr243o7k
SD2BA9WbnWLcyElpbssSp/ei396ZXOd7lXtcEHUCO+36r4WblRdMTv4BP9tAtvR6
iEjjyormoc/GS4aCvo2PbBQr+VmkRK714AdggOqWn3nuhXcgjnrWTH86j2ezuDE/
LBLbKJN0GUtwwaOklqbBHOunJze7pUM0coqU04WtcHObZ3OPsZwIJo762SK2dLUl
MayBeqjYBogVV9WrOlQk02GrmpiiPmX9VmCavpSLRB0sDIOBF3Zvi6Udvgx5I6zx
2Nx3qEnadWtE872bGl5rdMHegmOhc/KsD1ZRXbCMlTEfqfq61MqKOutozMcj0QUI
g+FCnJcQnhaAOLSK8JZe9G2T9zJPj1qFq2nCPzSlXjn8+RHtGfNzgKfXfuYB4/Fo
/n3Ge0yeqGmndJGImDkxdetQ6l826QhkszCxgo9QxhE8nZporWCwyBr8PMc4chaV
hCPpw44HDenCfI9PvbGmWrAjTtd+dH9KQhguze/U3GNEhcN542aZWBxM4eRVnkGV
mALB7vVSJjX6NinX+8+zgLXEQysVP9U2h32LJKL9PRlOkYaswt+5jVCgwl+bEjly
YGnbU5oiNDbOCXpxjJNDv0ZRXAQoraAdFuKvAEHH1+EGfUPFNuB22T4uzrku/Xhj
Gcy4u470kDZ8Je0DlEREX/vYp3XDbRI7JEJE2nkuG0DUP6ZawDPpRT3LcEwHNvIf
5Kxor6KT8EqDgSiYUlVzMei6fbIPhTiln0CODLj6DCy4HbZ5HzI7RxNbCmYzuaeh
h6bnaA7yKpH0WGgW9neK2emFi2z5TFwUa+Ijh7fYEQPTULARRaof9uhSf9JAzZ2h
SNo186Bkoe07dYnN0K0qIK4xwpCIORBIw0sMsWE4bwkzm/OyucIGQ9KDgvL6qUhE
MTVCIqdBdm/BHd5tYkFByt1+G/LT6uHKrDMdO4n6vYq7zplumF9Dpq0EgMtw9iSl
TZWSDsKDyRXmWPMppWqfsYMtkAFS+OO/3boKGfPclCMCnSP2Gyx9NrwLVJurpVL8
ggZLTx/Al19V/EFIzFIhwugtwlQBq6ectErGKh/u0yeq1vdYtYM3GIPBYwbiq6dH
vahf7RUpr6TSBpSEYUzJa8mgsqP/ptPfy6DHYDgGT9DNmlpnj1+VXs4RGDMBGUqB
01dJudaesmhCTFx9UUSpZD/fnjzPdtrNyIrERpwJ+lwJYJCY3FOgOssRtrgz64xA
Trqy/god6vYfVrQBme1KHNagw9wRNvoi4J5LRb8YyEPJ4KyQv9cAKdKbY1ShtAiM
MAO7YLzssnVw/Gv4XzVszQZBegYw5Y482hS2ozkV9bFgU1FXByuY5GDDBrGU6ppB
lEpwe4ykQ386QTCYMnj2xcWm9lmBH5VtJrq1pcnC/X4Jf4evoYD+D/3ALrGR6Svs
NaZiwHkWjle6+MKcGSp4DQ+29yflj6vGJlONWsGcYTDOr20Qcc0ZzyJMslVD77iL
CQGb08RXhuAFM37kpeCSbx1dp8fYNLg0331hGvdFP0MUsLUuRv0J9Mef+nbpBvCu
Hv7bBdOs/qtu30yNvr4GWyFNc8rURwVrV2xE0SoA3H2UlejW2cY0N0I8j7SwkhBL
jWjaFcx8w9T655UIMJH3wE4hmRrW8vNrDFy+fuNogoxOFubsOlBW2eMSytoQ+SJ5
KEM2b8FIcpUvKBn3caV3aD6xSBpE4wtHR4qur0fBf0tGEhZ935tVOm7a5GlYnsp/
i7kkwrKQZwk6NH9Yn4f7z6hHSYUrw/uwXrodC1OUE5M87BuYG+R8dJsPYk6ItbM4
9+CJSphhcytDf/XEhpqamQU7+8ALEfal7V3pgBpoKPyTyZAt9aNeVW81nZuGa/hA
0ufhNFYnV8AGjwA8PuFY+vlhwrbO+DEbT5TjJ72qwLLivDEC1mLHx+9aWDVSUNlR
k2WV9UZTOJEN3Hy5GMT0QaRNCLmchAQhg1MWI/eV4RDdxtrfxaNhUUGh75NM9Lnd
hEtgneDPllY9PVWC2x62NzZrT2vL0pVQzQfP9Bn2isE9ZdCVN+CXPVmYvVuGYqp0
exMHT5PgKiYMkIdtqKxT4PURy2JerhJFl2nlUi04oSSHbqBdZjUqdT/R4lebId9E
4vAnas2UvIdE9jb3gzAJ1emYMMGqaYYDYWBqrTistuUIx/XFfquGXvHT/g8DFjN+
LK9EkX8w+mc7uA2GOGTjdOsbywl+HdWNV94acRLR04KRM9WHbbo+con1DnyL/Jll
uJzdIzUF8hfhuR+IZ0O/Mrbq3Q0CTcrdixjpQkVBafjJI3o8mn1LA7LjcYtaxFYV
x9GpggQWBWKpOPZUjF178I7pW5OM5OOiIC7ZKspJIO/RZghnulYFZ0ZDUm3d9r5j
AFyjjfuDoA13dt8Jy8ToNY01CCThWq6moUs/YuqZujH99XT7Yyl6N7iLWSoUSe5s
AwmbXdX+NIfAuL1P18Qo1fbLy/zak0XRo8XH4y4NY9niksJe7pNUA3/R4Q/LGEGA
16KWPddYdlvErn1QoSzIvA1wgAvHMHTewvti7dqoaus42kxzQjU5lX4nlfNTnDWH
KmuSQ5A7cJ/Ce7Gp7UlYV776vDiPHpzc+VHHj5vsXS7KQpTOoJJ4qLshF9mp/fhI
CBOiSnsRVUqErcOFPj8HuKRX4UZHXngyvVcsiM5PcMf5hduogQYyC4axSbIc+ehp
5SCDp0oaENc4Q8EosSJOVw9I0ld4B+hdjUJlhQChTF/ix6oQzH4pIHgqHm+oGzhZ
jQpg04T8TyEvYLkE34W9r3vDQLd2m6R1P+6z7K1HeggBU1B8NCTZDgsMNpDPEN9V
WVXXDJmx4d4gjUPfsBWu3O+dJR/VDkYZmLJKDvB3UD1rrD78Y6InMMM8wXQkhCA0
SHyvraaErZkyke9Hk0QaX6E3PHeN7v6GHvPOvlXrJjINy3Chn4tjwZBqHYA09yqZ
cQjTcrIcdBdl6wNiCbwokt+v3TqzYkN3NpwVVwpJBnUBjBusTU3xT1/4j0iplDJR
zpApC43B75UhFSskpDa5ZySBM+SNoCbi02ztz4+dNncveO7oPZK+qJVB4gwrUXC+
M1X7dQezvbHruocZsJ3qQ6dHH6U33V94C2rF/tmLJa+AsNpe4IbUuj8AIAlGhiJf
+X/5ZYds+ZVxad4QzcBQqSH55O40ZuSC4AHovKHtC6Fk0w5xHZSMhghRH6SnoB+U
kQDmj3qcJPklEfYfDZMFdNAd1AI3eIO4FvhBrG1IDPKWBi4sUor8/VEo1k2sC3t6
iTI4JC9JziawLygt52CIyqLyZPOj63o+3MzEUan/CA8iZy7y7YOTJ3IPGIofZ+E1
j+I/c9M+VE4HonugsNkhWwxjiploC4OEsE9cbH81C61qkqcpWq298YiXhmoI/Xou
lw5DIKDbcxEx4D29/Qs8Zvk0pA9Qr9y87nWZ4hXkoOxdIEtNyaaBpXz8HOvq+poz
fuXeIAwnzUCcjB1bL8u2pq+tnLUJinLTmfWopaEUTq2KFOT13wMof+px6P2ztWxq
EmrgGyf1hTwgZ3kuL0ot+aoDuWNiA0sTwT3246H/it7tnpCg+AyBDSytCLPcBhl/
ub8JE3d1fQaU/9H6VJQMotpmL0DsAT0MRN9FtfYhUwO+tW9g24Hxlu2GwONDcIYF
E3egoj8/xrXMgMB/ciF6LT0LB5EzJ05qfdFrbKevly0/hLlKooMI1kk990/RO2e/
6bTcaIUCfFi8jSacTMRJ6FWc3jLOCPcZmJPX3d5SUg8Ij4dCggmCzxF/CRuw5zl6
ZDOAme0XqwKJh17BgMr3yPsNMLUfxsh0cB+5SaWqlMzeS9fOZ5Rdb11tOqnxz5Rm
dDbWKWtBcfVwkCzE6H8thgvNrhHtUNZ/45RB7kmjSe7W9vIMNJ/d5MpLEFBDPzEm
9tGQ2ynSMrS/m4iXuFdsMwO8R+NMjcaBtDO+qGhvKcOtYtfhlnT4tMG1uZqEfDnY
rPCC+bTBK4iIIxTXQ3XYjcV6cECDOs3X76XBIRPSI2jHLVjwPb+aMVLMutoxLpWw
FldhiatemjySDoZqIv3JeCMYor8CAS6nlYEsG2wEzeJkkl1USFgpOyyUkoC7p78l
H3DoE85TZoIzjxloCzwfVl3MKDPtE3F6gYSkzI1khZnLrA9vZGb5ACPnHLRX6JtD
Cx89Jd4qt2RaOawhOaay4duR7tU1Y5CUezrw1kayas27eRPJxPRIa06/jBES8EjK
gGPhLHmW18x7MzMKY+9n76fdqIo1tXIaDvTU8J1wlHfCrxJaPaMWgtAyhdpqvwNV
R2GfFRrFhkqcoB0Ytigg0HshkGj6gH76wcKHs7npsHKmofz2EZpWOKXWng9dIT6S
CjJrC475nRN4Zq3hEq7PacbwoPF8QlzlPggiuDo2QV9aFaWdfrI5eILRIkpKyV8r
eF4UOkwicUZQMQOmw41MxB1abUArH/g4fiwVQVkFg85A8PcCs5pW8LxUK4vf9qav
NNbSKq6lUMjpNhtFco2u+K6QEeCiIenfup1Ldf3bEpd9dIH+blqTISTzmZPcK+aJ
4+oueixfn1eBj6KPW4/1k0hwor55l99VpL9/iSUKMlEwll1CcASxEmIPIwt/B1Vh
1xvcJE3EHewqG4GnlXt7agXhiWqJyGMS/EluGboimVp47oX+KcuhBjAiHP7nUKR0
z6/F4AafU5GlOvtzz0RW2A9LFn29WEHtsK967BGhVKQ1rWjSVjFKwUns99XeW31K
Sz+US+JD3iMusx07+XohK/ntCL8YMXkE+/lByjqSyQGN+Am3wYUgvCfb4QIRdNqZ
GccpAM2gPi2Hy5EP8YM9xbyP/phN5iCAUE41krk7sUn6iHX+aB50cIm2pslc6SQT
+UaaMtTR3qLhaj064SNtp0Mu5Xl2PXkKS9yXYJkbo5AzrZ68OdOfLgoD/mfs65tv
5989Pm7//4j78DQRfHIshyBI3z0/2LBLZnas0slQi7qiqQ5z5imQgY3Qh5uSKbmS
j9JtfaVg0Dzn6ZbT0LwVQxunMRZa+yZfpT2ezbd81fmxw0q1WYMLUhRVKgFTc62v
TW1kweQ5cEXlymrjIHcMApWms/FUvwiWnqyWDma8jUXnJ2sdRF9wTtNMrASrO6De
0k5ndmnqCgq8UlU8Hbg4qwGEKQZ3D6QUwe0675K/agGC91HeqeXbpiY+EGYVxWYJ
J+ZP6RNtYKW9qWlGTKEMFYshrbh9tRvzql6niBj9LGaoK3f9pq7zGlWJDa+crI0T
Wz6MXTQFsFMn8pEzij8Fn66jXiCz4u13+K2sjgHTqPb6LhWp2bTbth++b967M3W7
Mh6L7ke0FR3lHHl5qY+wuWcRKCkD5LR0Me02OceUNNZ0bu+g03z6IHy1nP8kr0uh
qS1EytzNiWSPJXArHEF8LZ3IQb/tlXzKVSPfPpy9XjKd27Grsm2pcUZkHYkpQEXE
cp1qAj0RMAU8/rpcIYx85ORd5s0YqML+5C1giY0m75ou80+wYqdP58+WIqua96Qg
dU/fLe0DR5T1kfns2M057tV3RX6GHJsC2bTlUrOva/M+61WgwFKrP06O6R4+3vHN
eLdw9tmk8FJz6FXygkmbuZS3TuV08WeBp+m1HRI53raBvN25NFqQN6uzg6F43/aW
PBydcAvR97Ll+cDJx3zvKPPxkVaGOQ1V9J8NeX2wsjDA8bK1g+/uAW2rDo2t3gYY
DgiolAlrEM9D7KpVZw1GEzH4UCF6c1zebQAH1THE9S3j3TlRDSRgHLpEFOKlMAio
g4hOgoaDNPtHw0SVjPOPWusgHEw0XhVqqlon42Lpl4cOPobXUBc3382BggOFRRmT
CEcijR81hQ/l5Ug/7KJGjrjXW7Kjf70wLPQd3zXivp/qjog5NLXEOgVdx5fxnT56
40KiiIq8FwCmwFvkMLARHIAEDLL0Cjb4Kfrq4TXw5Kpe2SwJ6UAYMaeKTmkPGGGz
rAlvur5bJgepKlNxUEGXIYuLtqh2iuTD7BLGWgcRS8gE1YXzirFzHX6ZZK7R+1BI
Z4+VB/mr9zZkYh8ogygcVdd1eEQPoxfQIBE3CEKLTHPZAWwQam0YlvGq7dgKjAKo
ZABETPd1ABZ8y5+/gxSNtv2b7BBACDzxVdlVWh4BZ0pdh1TiUauKQh/lYzcKRfHv
KBYMxxJp5SyRUuM+lWQzqw2v71Yl5zPlMA6XOAFjPW3LVLBS0zDbEWt8mxNk3trl
csbByMdHbrPsa59RJKYzfDdA7KN8wQUg+0sKtK1wEmGIPagoEP4to/m8CvphLzNh
ex4Wf0sQ4/6l2F9HlWA7ZkMUCkzt9wg/dmakk++psEeSRkLT4guSr2GXfNqH7AjR
a0CLwAisaYe3HsZ8m1tZqX8jV6vFynfU95QxQLYiB9nTn0tSKKCjjVCXTFg2+NI9
i+2CVhVrXYYKQnsCJKCMCGK8+H3q7zLSmMEYpfypNRhh7zyH2UwDua/P8zy7zJpM
rDeCgmB56qS/jjHg9owwJSiG1V+h2YlAWesOhZ7aAuzyN7KRqnuIGfZ5UA2cF6KR
+RfHRqFAyrEaX4QOPdxO7Il35eb5BZjjAzF5o2qxAcSnHsNOzs8/E3yQQ+k19VUL
FKHMWTOR+ogbGe3uvkjq1/W2S0fTHOe2KkmX+nPt6z07e1qEItS0bljl0o+bfilN
TUA1vO3NuZpar+mwIIDMIkjV+Oau2ut6Dh+QEhATm5+GSOghOZ72TPh4lwBhQNhx
y/a5Bkm0Nj9gSOKoAwPG6IFBRCG6SeydnyuBJ/+cZo4AkBcu+3ifcZBEFnlFn511
6THvIa38lzbHPg6F7wsdXOricqi980Ii0ScM1wsl9NV/h7XyHPNlK5FhjuHunQls
BXDbXUiJEOcG89w46P5yE2oRW+tM+FBiDM7LZFWlOu64nK449kWLm8K3esYflQd8
gGxmPhm/sgELS0ImFzI0Yi+qhMFA2/cQ1UyLRIxts/gY9euQhBU+nGmzUUsExyst
332e3mXz/IhZ/b6i+lTy8xoA9NWSV3XKM+pdsbjfCnc1LXym5GwDw6mK4B7hbvyM
ZwiydUEx4WOTA6LQfd5xoigfgShfwvzESBASxYoAThLD2A8yX9nlD2ZspFSzkx1O
kRQXfbQWLbHseIzMEMeB1/DL9FxcqHnA/GGN594gOMzkZB+J5RBO5HrWkBbMdPXy
UUbxDoNrYlK1Z0xK4GIwIfRTrraoQZG4ChyfDqZuK/xChvgOd1HX2RlH2VYGANNN
vqWYByVQChvYkV4QSURrsTpY78cznv+/GvlAevCRokvCgyRMjnabxSlrAhElHvU5
RGXugRKFUSX2Uqiw0kh4s0PZbIcSPTwLVDr1NksspfwmY1RuUgLcL5gZ2igcTNrV
1pI5ysC6Nec9bKhVfhHI697Sv14FOYeqfIxvm5STJaFJjSCcCQmcPWZzs0lSZo9A
VTgJvsd/7mqM+PN9zLQIar2HeDcRoGx2Y+hcJ2kHSoyc7HGr01V8J1VQJ1c1fpec
aSPrf8dT00Uti6djuOq8p0Sfv240rqyZ8H+X4q0UAEwnng3E8nMG4TunbjOGQ4RB
ODdkARjV5NxqFtlez2+rDb2B3C+jZpMrjNMtxL0GINLkiI0Lf+sqy2nJuDdQ60Jd
SjNTV3XLKy1r1wI5wBHv4yIjNG9cMUkoc20O8rVOXuyoI+xHmPgeS8sQaHNlxhN3
2ay2zpMqfCtx1aWgFCullCcNdVTg5HT77vdu1IMZb1UKPtiLVmlRU49fzS4KAn/l
5AK82WD6jxPhpnKOUXezhT/Hw5yczVep5u9O9agMiTPGCTwQSHoAeDP2vgPOEEl7
PKNgTK+45LqNK0c7k4VLGKWY/s1sBglQrShWYXv9mXb+CuBGLTYuL95i8u/IyGWU
zTVLBjaPrHgTJm95eMHXE/ALjEKuVc223wgpcU7eXn6qpWV3wz8WA71D/TeHRu6b
kg6w9jCZFsB3Tf0nH9qwZ/fLowjcDe3S30TDXjnSWBCGeNQZVxuhjYYYtxH+ThFR
H8Bhhjli3GYc0SNbakKJq5/O1qkoR5NQyBbH/AwL3LWk1IhxcuM/fV8esVyaZDer
/xYSaHdYcl9HYGc04NllXgPlUsl+fTQzUoluiHNDgmkV/fnTie1FCYd5O7QwcQu5
unRNuz/qZo+TUsrAFuoiu4hW+4o3OyC+H13f6DlIYtM8nakRjKnh8K9E8l+7I4OD
DSBPcCF1esLZJDzfZIu8VuJSViOLXkeMmiIOg0xE9PBsUd5UuWwuJOJeLIY5kC8t
ThFhKXH0MjeN4ZTybaIQRHYi3z2g3Qq1QV4Dw2zsuEsNaKIQx65Q4iEOIRvhyIze
UyWVWhcMUVlCpz1c4kiTX88hyABDH3om3rJpSCLuffjpjhGOsL9AESXsF8m45ZTV
mxok8+pu9AVaw0Sq6ALwo24BHcY0wrTh1J2tBxOE1PPPlGEJ/xb8Xa8xeWOrHcRv
mgMlzDU1fCamyhCTxfZCHu2R32H99twWQ9pM2cj1suvVLjJ6nn4PmdSEAJ8TsoUw
7XXfZQk4XhqN3kpOwLHt1lWIzkdxUcG/V4ICxCf93AKvyQ+QCsROphzQzV24cWNi
veQF5nvQGzFGT4PwG24DwC57dOWVYoMxnzG2wwZTF9Q6ItpSdyauRFCpo4AWgLkY
054X8AQ2nlg/13KIWQvtxxATM1rejMpxprCIRua3rvt9i3Ci2FX8ai3c9YYKQ/le
L4MS9qCrJfDIl7IOOjIepc+RdAGa6iCo5ftLQyyCCzlU5wT7ZnIE2kKd/uDFIBAT
2V1sExplfwTJL0v+BZSxvDPvqwbB2U56tfq7mDjVjhwo+RIXjos35I2SKZ9f1IDs
zeRFrG+tsm+Ta8g0vyCuP9+upzyjjtMKWjSLfn5tU2A7zKq+ThUd3mkhHqrBDu8m
h9qDJKkYHugaBqdc/DnYxN7vUcNdS91HdOuMYoDh33GJ8Nb2avAAYf/1mkYs+bid
gTw1v096W/3XBapP3lQ7D3muQR5coPP9cw35cegAOZQnzw354s8SFZBjOfkJf4rf
XI7924ZsqRoXgXZ1qJsqb/icZCjoqxyOPrebqWDHdq30LB1TZ1sVDWJidmQhWBYu
BBRamD1YwJtzNTkm8jpSBNar/vaQSmdCKO6jgnoJvDwUS9PCrRArFTic1DjBQjWJ
l0azXW9Im7OIomo+nvu6g2FggklMPeSGUlBY4nedtiO7BZ/wxjhlubkEoEO1FAmZ
lga+Rqi8X0+KccgHz0eAb0tcVVf+sCBvk9JIBuT78Jvl18Xi+muMFS54+GZhzW3M
B7kyrSuAcViC+6dfJZCIqs3/KPrmj7VlZ3IMroq2TYXEXF5k9Vr3LUxnVbp4FGGF
7XqoVwKICl2gY/BI1bAg2S8bN/KiP+dfU7VuZgZoEAuFFqlZ+HTkrhLw4in1viEX
fGuC3pHn9EapoOlCLueRDO4z2+Q5FqOp7kmM6JCjdLEsLUv722v6sebAmw1BK9fz
U009O4VeHK0/F4514L8/6iGhrNCSxzRbbJFaQ52WHm39ChlfWoTYoUTOpW7emzg9
4ScUv1wSghiOSwDCWQ8xGqcLzKAnW0iWE5Np6jrBUTVmIHy6JO8sAPGq+jnCuVOf
s4gO6AoyWMEBCuL+YzSDFneZx/m2KTIfPl2nqvkaiTSQtiaMedv8UhHYhczH1XeB
xMnb+0EBXmFrUo1l4ooQgXeCg0pLlt7khuS38f4zDfutcSSlOzuuxXyLskY8TC8i
tO0msN/PEyddJPxs+F6oYiYcpmHitcZgcuHH/daNXx14d653xM33fBCs0os9z0xD
uCL8MtBzfY2QdzCnE6FN95TBl8LR4K0hDBHjHqIk2XRvSwG2Qhfu0UEc0umgeL/O
29UKv9yVr2gpzR5/jOupe/jlWbcDFc5iC0Y2neHuHyVju0UUH6dDWGHY/9Myh30e
jYnN4VZSJAKZCHgzHAPda57B2mZ+BC4k21sEbZl++fhwSfyUg6tBMP9NyakP7bC+
JpYXxp4y/euc9MuuUa9vzYq40ou7N/grE+xeApU0PscZZRAPPjPj/eQG+QxAJmqy
alSFfs95E/IhgedLjmOLvb5/U/W/hEZaALhqNEZlF1Q1wdSaDEIZqLkFFZIMsf0N
+Hi0qU3E73JfGcVCsJoi2TajT9XkNsmmsMemGAx7MsjIisRDCOex7bVxcc4wIjuh
1aej2k5bDCBSMO8I/PzJhChHNpOOmPA4IlplbkuMIFPM8tdEJcPaYuLkDvFHMNF4
NUaHkxLAC9Utf+OwRqS2Xlf/SRImE5V5ZZg7Nysr1qcJ5clYjrlXRpXFHsWSBZ6/
B8Q8Jjyo5/AgjBGltYWwwRtXFRr1k13bQmyruYwUM4G8pwpKZKlwjprMrCoGQAhl
MxGq5ugNcWD8I/3630TPorOMPl20mhuk28raUHKkzK6bnTyndANOFvqVYANnfK/f
PGFLK855eDu9T9Bbrc1iAaeqTG9s18ivK2vo9jvjfM9CnwzGEUSxH6XxNN1h0XpV
+82bKJR4gOS5HPcO6QY+vYbKHnF8lUnVNi8Ab71Vp0TVOfx3GUit+yfqM5CGqsic
P0n5vK/Yqq2iwgWlzkk9GXEHK4q+ZitxH0ysj1nuWplJZs21g56+XrdY74FplmFu
Yr0eKI7V2kxCaX3pQ34gLUG97cY/3edvOt2Y54AKX5QJLAy1opcWhx8MVkwQSD61
m7EGFxEF+GTJ4mTmsg4ufJ0wvbhOpLGMvRda/OcUKJ35uWN+C/kqJ42y3CEZP3bX
/oQEEfHWDo6VrqfxZkpjiSUpTDYtP/ABWGAtsrjh0bLlYM3aaOkzx6lnh027XOF0
lj/jlDo2tIY/fGvM51oJzU8Y0VV5nQIM+xBjImwlKFt4JZieLam6KQFVcUHm1dr/
01rc/v81l/V7ugrIMLLUCoGOvANAIn3Y2j07pyoRBtOqOExeJt4FYyExVnlKgUWL
ODUOtq7gL+frrmmZyuc9wre5EjnWAkSzZD5P2H8HjcfapGimPs4AfgT7AGJmsT1F
aUwqxY5ITba1IfvfmdgDkPCijNBHYgm+PdAlaJO4cKqvcOPsSKsXCVPQjkeEqISh
h5bbcD0iAgn5spBgRCrJbBn+Wh97UptSsCrUwBKfbhtRYDm4Lpr58uFTLoG4V4J7
gYtXDjDX2g6LtrRHQUeIxw0pyFznWnqyjypd/vTh8VSd3lzScHsiFx/Ww5F6LAfB
JI3WqZQkX2k4AvWwZNJfEWSo2oJxlf4shJ+o42j1Kq3/Gg+M/qXUkei7/ayExoiX
Owx7fBKh6SRIO1kBAbbztGqlOReiYBZuR0eW68Tfx0k92bFL+uij6ho5IArn0pFt
RpVVhHd9SlwJu5VGiia+pRz8ucZA7n6EhWkt+iJYC6jugq6lN0gljnmy/Ig4iSh9
fi5qoFRxgDeTfK6T2C2ekfbeRZPX6C/APMQSwmirUqf+SL7ctVi/LkLBL1v1l9zb
C5OEN9Sys/RW9bsel2FI/HVMHsGWfzdROuy0MYHwtOn4lan8sZ7X+1eO3V+fxH3e
d7mK9oapI93aWo3vJkK6TNze/8PvpqDI7CVYIE7+54tSkZkD5iUGZ/RKU4PW25Q7
nFuMo/kXoRkOTc2/ROK+kVKyQIERWfipNiHevlGFfNVZqBaaZPNbSStfP2q1FW8A
3zO+RyNI2xX+W5BsjaFsoxzvKNaDEJ0InQxd7fYR0jYUp0ybwXvrA2T5xOMv2NIz
UH+bJkYIUzvbiP7lLW1vfSaST0SmADBWV7cTaTlld6QIADoVbB8ecSv8MU+Qjaz2
uHN5Z08t4D/ZWqhiNnvPjeJZAKWUOsfeqJ/ds+K4Kgt6qO9zeQlcR+sEw5FH/xT6
xQEVNHh2/8M6QvRHBAzDbDToGzlHk9ePM5HNKj0bTCcLEceZWePdebzCPU8t1NLZ
ZX+DI34BqgDw44nWCI+rGCW5jdMq7wriu44XtAnHmSSWRABG0wrd9qpiJw2Itzy5
o5RoSSM/QxDb4fwNImIGEC0OxOBBcgCSfw6U/xCMoper7FpPAL7LtpldX52c9yf1
Vqbj3cPKawlzvQilHagsAMNhjAqiXMQQyszuUQtcpclNKGgWCHGZkGWvRut2JjZH
S4/HcXtgXfYR7nlsMASYmcE+xsP3N8RaeEIPEEMOWFSRlrjcRCkf0pb2lOhFA48E
zfunDJIalMVGfaU27AZz3P6P4zjaOX/qyc8qA3tKQS/LvhWVVPacP60cYGJIWHwl
TOiFMakWwsBEHGoWzUufC/UkrJDeLSfJ4nk55szVYljwfXQqjq/yLrC0b6tnzP4l
HRIXJVEW81quDdZgf73arF9kN/orhefk5+nRGK7pXMLWYsddVoK7SYAD99yyA05u
eiAxHqkWv+GrwSqDQtqaOeqkPf3G2HVlkh90ZrE8bPEg/MinjkwEddI8IX+I+UdE
w+MaELvAzJa1stlO4ROFVSx1karCUJPXusR2KbmAO9zFUOlkIKinJMfABt5wkk2n
/T6lS7M42uuqRynaCR3BNyyx7qBUX9fcDJMo7ZTr8LivuXpT6QEjwza5aYMX/oRd
Cx5r3pxDWaiQcCu6tZmSfhuQK8Ypj1NLDbJyCjCVdouo/mtLGrxVNReUqaUu5PZM
huXXn31Nb6hiIltsed/8IuDzgMof7t3dTRVJ0aJv0AzyCKrms1kjV/cq8LcunQEc
9ZPQUDojfAuACbmH635/dZYIGmMaq+OAX8KYcS6OdkIexA0Ngw8JEV2ZrDlljibV
NBoVQN2dAg3ILZBQuE3e3w1BzH6KAK0S9N13W++dCqdy0d2+DmcEEIJTxmpX0Leg
O76gWumkMENJUjvGbHJD/aitfGPQxQpUvZva8+0PHy7qZcIVzUTTVOkA1dvPc4/c
k1rLVqI221K6uvm5STlA8c23+MNqfSHwdwgu/vGudlRWfHhW6aIRzULvehJ5ynQa
vHZEfb7IJayamehrQfgK7y7G6jjHaNMTeZBmKPYlNgGAant1VABXWY+PCMnPBX2T
Bpvz7iGQKIzOMNt25UkGiF885SOSn1zadqm6J800NZemd1jUPQ8wqgkPVde2s382
jriWCGe3Uf0nb1E5sNANJHLvEKHA+BVVByxpI2AeKlDJ11AhubKA7946hBuPg8aS
g4SvyJsYDfz/77u7I++N//rzKRvReJRFEkUxmnmyj0RvA/AI7MP9zuRJFBznnil9
asnoLktBqSm911RUfL9oFQ26hBj56K4xdRV0sOgm+SsYmiirnHO1Bk0Y1tUvpqV+
eMMWYTqNUh1qgqE+he4YQabJJw6pHFTZuh4d8PswDfZHPnFnCMT6egEklO1PV5Jg
3TlQ9B3H+46XqaWWh/Ws0d9KBWqw7W7kCGTU+fS12Y4Xdw2FfP0IhgMHBCRmwGal
h1JVWei3eKjb5/lAaTR7RGd/MLZ/9UXLwsHE9G2HKmG4NrLzUub8Oo3CYpEkxuRy
gYdzZ1xjGBtmVg53DCnK+BQQAKVtF2+zRuZtQBNJL81cr729kGt6sEumbfMBmgvT
Fl2XInqchNLQqroVdW90NzCxvepx62rmeycm6NlIZSiZvYRzhvUT2wqLkBnU6qSS
stUiWJ/siQf7pAayMvp6SLiuUw7pwsKjKu5phTB6GjgpgmS2bXoleQeuBt6tJH0s
NJP/2fGu3adV5OlBUFK6/SX2NtSPY1S5zmLwnZnhrkY1KNa4oGW8dtWFyElcP9VZ
xdVyi+Ig3kVfpawb3m0ss7AjJHKn011GVN/HoZwuWkrS1Eyn4YWHdu6kcxhsOE2A
yYtcTmB/0LRTgKhx5wKZ2nxgmQ7Qjt4YTz6DGvZcJ1rmYpCFfe1azM/9Iu330oOW
ZSYg/h11YRK0XmUG7T6DsEgoz8dt0F0JigrBsIoPOIbJtmDqP45NL1Ow45jdf7iy
PvltRKDR6vP2zzFGucR2xrD7IGJjoqMsrkUpnxakZmN09d+JX5p84zbgOUc7e7q9
WwUWHHU2VgKQD1q8gYOkjX8n8+lUJiBSLj7kvRV97QDHGuKC+UDhwtJrgwWwi+wB
3a+KrrJ7jaBtzlGKZxioH67QKeTuJ6rRbbRuBN13k6QTcXpn+zCDIoVuhIHJOfMX
xzHPnZTThafdkt4YZwaObvobx6b+T9W20R6+iqw7DnVlHz1PKepL5+wdgrOzZc7C
srQaUMu7IiVdh/J+w2QzqMbMn3CZ7KdnjClPQIiWT12Xz0eLqPAWBIark78y2pX/
ICdurm/ngop+DwAkRNHr9Of2s0cujI1Wgufe75RvJT2QEX3p/5rd3zLc7kBwkrR5
cDaflFwraCKRdPd+4KUKssZF7qPcA4Yaugj8sDySGgOW9rciv8ekL/+twe9PZiiZ
XIvmXmi52hAgbgmZPqH9stFw8YjEWfHynZ9G36WRRB0i00Yz5pdmT6CD1Gw+SONm
YEp6PexEuPYh5WsRl1PNonwbRJKRigOj+rzjm9AO00W2R2/Fpsk5BXsJkgWoIQOx
6GigDu2RNI4ZxgKX9KZlPet8xs774B5tChDl0r9Avmxo5L3pOl8J5VUmu05HoZVg
XgvaUYbd/4ADWw5eb/blHw05n3D/ahf3fSDj3xMHZJejUcYubyhIoo786ND8bsF4
Rpf41LfYpfEiOiK1xygHqePo8+SG9+8H5cKjWsPZb5iGorb8f/nQ+0R16p6m3xBj
z1gWz/dBZbZqzVFhdOK6RH1lsyBb/WGB6TccVNu13RVzMwNDt/UU00CqdtYdKzVm
mLZAbGNYAzFTbW77n0vqOwvPJczpQ/AQ7nAmP7+1kBpbQjgBz2ZEoshy3TxVIOzG
vflWC6loAZbH2I7dVB94GodZXHkTiLiHEe62Vgz/2tfMSIXNxSzzCNN/HBz4B42i
7RYH/QsvfhYFMJMV74K8ck6wOoVOtjk3mbrmFTLssv0gSBIJBG44c6CMjajSzA+E
QslFhFJzxSAYQ3qrwdtKdm7WgP3a1e8T/E2igQvqBQc6WS5JO2O+97ER6GWCaxyH
n5JSpQ382fUJyVaEtqy1OeFcPpXPvcMBPqcfMFunjRKujRadtvqEjiJfUkqfRLd2
7vFMGgQySsU1R8x5kFGR5UX6o0Lqu3HvhosqexYTpxP1I7FUAT2EREsYLojXBBmr
yNrle6GDtFH/VAByELyURxq3jPLfayF1G7Engqg5elh5VPg5SvMwbaVV0QMxCzbP
2dkhIxaTJKztq+KrOzW6rDxdNKRZVcBLURiYUol0kLF+aGbOJxXBjlulNSbjRmYP
SddNdXu9PY8bPEkeABebqebFWYn/laWjMbO3IXdJ7fgWgsYyDQ8r98yzxQkC/Zp+
mWwINDv8sbtIZx8XqQvRekYNEITHFEji/X/liwh7usMc+PYSNitGx1KxAoS3wyqo
5C1lLV3q4euT0ynA4CPjBAo4RcWIXgTHiqhZk9jH5OU4IpjaG3FYGvGWxauBvIJd
LwRti1TCSNxTS9vjW8Go0wZX/5rweiis3ERys6/76iaPci7dP9F8H5dEbC4yEVKm
+FopnIdk4BbxWu5hRVX0QtZokX2wtuh/kiLRlzig6DAzWOfsVscT/6PAu5SsVm3H
9K8xGTAil6zPOqhuOKpjHJXXFaPycQtPAgqvG2XW4jKTHBMxxX8Nn2FdkxYXkbE5
EBxbAU8P7/8vUznSkiIHVFjwugpoRRh15bAOVkxu1iXE1uj7/8PuZ6WgI2MfCnJw
IDrYwx314NDWgBEh6obEHf1ZIRHQ4qbgBPWHcjgIqBKJjhNEMZtc0F5ughp1St2q
orSNVebPJwxqtfG7ivxIXNF8OPASY48QvB7p2Fberd0KdNI9nii9zcxe3oMIWUca
UyYF/qdjR268cYsbvF9raDu3q/op3p8rNdGve2THAW4MRwwW8PtgHOo9TCaYPgzT
MXyM6Le6kiDdSQJJLDPrnOsc/j0Ai6PL1rsyrBUCKYuRjOnGs5+zkbnuT1uiFt4t
Dvt7SBBhXy9w9XSEqJ/n6lHRiro8YZH61dQUw7K/x6pl4QIZFNPk4yDEuPIM5s4N
2lg1jPj5fc5z+yXcysvbZQ3DbTLl8Guj8m78pkIDWwp+/szrIZ/fFmPe+7yMgeGo
gqDF6gYxzCrvNHQ3t6GXX8TT3XIAIk/KG6XZ/uPk6DkjBAgtPkfOKEKC2z83ce5A
zcDQS1L85cgvNTigpluw56r2LbqodAORYzjX2efNQKQ4oB8Wu27nenn/xEkmfCsi
mrfPPahUZmDQmaHz6+y83LNixk+sDzQtz+PjfQ9SZ+RKoPjxw1ZA5+54rtMtzddk
6BPbF1eQRyD42djzWpoa2EAk6z+sRC/RT14cCZCQZGC+9zRHdKF53vgR3nJ4pfpD
dGmHLORpOig8KgsYpwGuQaXv8o8Q/D1RvXVkUz3Y7T0NHphR2BIND41nbZgO8q+V
0jXTpy2UM2q1eWWhlUoEDeepDneogizQh+iLgXXaF28n9kKMt/xXvZfk4mtXxR73
hGqTz5ko0bRKSmaBbaUQb3pomhPlMu1pIQm1M3jEaVTFVTkleJbbWqevQ7sQr0wS
oEel/pnoBiyp6BanWjwiIINQ37iiMEZK5ngugp9nsddOgA3DJRZ+BUuCMwTx0E+k
7VXMZXIhVQCN6MPnyZCX1g6FW4s7opKb5Xw9MCsmLTysYIEvDA3yxvfqAFIEE3p8
sexcpaBSYZ8KRTgpAB6RocA6po1dhDe4y5YkyJSJ5BJKTbqxYHEPNDB4ZjuidLaX
wL7q/62R4s7tygLAtJq6QX4/euXdx80en8oZWl7XKrIQ22SqC3eiC/fWU57KTH4l
8hlUDJH5aeMj5m7PQMiF5fXZtxAmfOmDGeLsIuqO2HDDopfTfJi2CB1hJq9d3rY7
7tH+/QzOQ/P2y+HvKFA1Vy14mb46ywT3kvONxmL6l0TW7Dr44D1MBrlsq3vdaN7R
8bYpsxMMmrYhtOlp2siBAK9YT6KzswFMe2Th+gqa5+o/oUxP56LE0a0H84ZK5YDV
TDpvfFTWrTRW8MEaWIkoWI64rX7WSnJuScxx/neGPyjZRgB7GqVOD2DRFQ0eUoFp
LbGEzreTQbyiyF5AHdTWxJIPIDKj6r6QlC979vQTX+zVjJ1cAOTlt2RD4qutt2Re
LIS38c86HCRRSg0WiyJ378MCCJ83tm7SUP0fAI2EuWLIsh3Fk/QVQmBj+ROS3fSl
LbPb/oEoLBZQ/RdFwR9CQW73TusspowTTypWpFqyCpDhYdJesz7LdlDpCU2s+R3g
PvZDbGLGBF85ILCQjy/ApAwhXjPqUD5ZwbnZNVbRVnVlKDR/XPacjRetR9Zn1uHC
OnRNIF6RgX9eLFeV2u/iBLNCdvTI1iB8cdcmKbtYveJI5OqOFCsIAfO/ZGooHgwm
GRBwgHHo7+YCwxgNoMMUzgAkSXd2dFWyEetFRmqcqe4IJJP+55mP3Y8NzjUFQDKa
l+fGGlwEcLVg4ybKOH8baoYeuS9C2AqfKgfI2PGBV0PsrRVyC2L7ASKnAsHAyW4M
sRDJUWBywSVXPk0rnKVaAhgnmVhUNCAiyyUrPzKZVgssyJ6zyRQnK06ykviDM0Ud
pO79JJVfYQVjmS+DMCZe1zB6pQ5ki12myu3XxdcDB4SYWqeWvcqnpx2wJL6DZ6Br
Mt8Jpyj3RCEKDiTFDkJ/mVbWsHONfEN/AoOBlDuOG3UAVEO27Zwo01Lpi2cBwdKq
7IhOMS24P/aZ40ZQ4bmwiPEnbeubRMCJoqgy3oqdY8vtByla7G+WEOP3dLqcHOWS
YjBblrNqn5dxugPJPSgq2uMu6dIXLH4+LM59GngnqAtFxDumCGe2SDJELMyxUla9
ZsAqYueuJq4mHDqmWRpUokv+iYIjOLTYhyEtfwSavLQdbrhabpDi5uwiPlXTQ4Y1
/9G9ZT+lR9NA8Q6fVNnWaJiUDmIkONZGBu++nzszccUFBhMqw7UsKKH5L+eD6viT
tdD4fCJ9qKBKUUUBN1mHN5/FfeMiym0gU5cnNWmrE2OFe6KCJUPqRJ815x9bvqLj
q11c5icYdXtCy2E63YSAPJUcKxdZuYrGZj9NZOJii1r50+rdWO0ezoHRRrh281Rn
oE1c8PQ96lZFi7E040O8MKWiFqZRY0b9bMjbrUweTKrENzAPKVg7s6EHN/B4CI8y
PsW5DK6w/0ZaTVnprO0gRKehboifXW8x5jUXtT65gNbiBI53admEGT/2GFiWWFVG
BusXfPl7DWYvrZ191SQbpys1IEGi6Npcy5guz+Xyy9UTpKpGj8pG2lUfz8QjCAkj
lwiKsJyzEfOM0zJfDEiEn1j3e8YbnSR1Aw5+JnEBw2PaUeZies1QT5Gt7G6ZXdRu
LqUaO4ttt60v2pxGsfAcxlw9dTRp0EKaoA053SU9r8j6q+MOy8jojKfk2ySxoYT4
/jY2VWeqD2uGHAt84R6XC7ExdAJFE24u+iu6pFllLcs6+MVzpAmH8nPJWR6oEkPE
Xau55XYszWv04mbRQiP6EjMgqjmfTc8Q0GhIeUDXzX65HZUb+Dwrm+vwe4/R5D0/
g73GNGU5mRtMHCkb7RzCuHgAbbanrYzBeO8djA2y9+UcbhJEeUj9zRIGYsRYBbu3
Z8ajAHH+xu0bOjKIan/QLclvbNF/NQ0gYcBbBKBEzyRMmcsYOrZC6MRHuLExk9XA
Ej7pPXuERDQHZYMenVTpEN0ZZZKueN279FLc+Pb77pDR9Da+4dBf+yxpfw7Qptf/
rZ5DZ/xAprutc6JWftE8OhqO8RQI8tSguroYRRz4GBg3WyHQ3gj0ZvcOMw/dmK/B
KRf2QeUFZ9br4ViRK6oC0B/CYw9cR6/NNYBvKyDD4ssCXjrkqtl8vhgBb8llBhP2
BSIWIqTRGDHPOkPzscQ4LgpFXbrUOv4C7pds28eZejAyAHGN3GOZyvDjKDdr980G
6t7K3gDoLomFafSGc1k/2LwM0Jfc3HH1FsrsG40gAtRizQH4q3CbQDsmXjZgX83h
+hP2pYGx46o3MOxxFLrj0fIHH+BSYyASOnPidArfsRZCrhPcAuK3qNIwBDOf0yAN
kndELKPT0q18UbQkIJmXh8KVRi88rwmJXATSSkElgNtHU/saWRtVpJRuc+Eqh7h1
IuDoVk706vmBExBSfe7BWc4f1KHC3/E1Iuw76eW7hMbobeNBPL2Z57q5dJ7iftIj
Tzqo4A0iA210Jk4TnX50Vwra+ZtzdTsipKVDpKeH6ZN6yykQaQWebLHp2E3wfeC5
zOSc+cVnEdlUYftNi3l7Q8POMJEiVBzjIqM5Lskj5kdPZ/dCqB+NagFdSf3nFBKQ
LQwkbYuHlNauzMQLhstcwrv0CjApozGuxeRxP5WAod0kz2DurK19F65inwHJCn0m
liO0HKHZ6J/SBElWtzEs+kf6nbtchL3QmT3PCaYaY0kQLW/iRD7yBffhubJIE2Sc
/vDYrtsPvb10Z/D2VKdqAx2zfUeu3+NMUvKc/Y5PwxWeb7ZBkZMQ6nT3kz4/DMr1
7FJ0bnOwIEndZ8LCDoHO8dySONNBMfK9K3ywVTj+xiLoIf9D8n4Ke9xcFkWTC/Qp
q5AhZed2EqpX1mmgZa31/LwarcE4D2Br7SeeLM4Cn/LtRrn4DA2SGCTVy1a2Y7sk
OAKZi8yX/FirStjj8TEmUkwm4E8pDnMNC57K7F3aJDOtwjYIQQy+KHJKUYbk2E3T
HUPHpgMBjpDuL389JH6w1dvDDAE36QN2CKfYvzPRmeFWeS6ns0lo5fjpbedK+bK1
CvzPz7oNjOVBj47YnGhYbHy/3as81XjswGTUXEo/qkY8Tv7GpRj4bF3Igswt3ISZ
wNrnxDF6crshuSuBz+1g8E7+rflIXhPyX8x+n97HFmYZqac+sFRqzHFRHITVC789
G/wn+N4STPDbSm8Dq7pQNZTZsF1e8h+/hMa3mXbLFIyYG5BCmk03V+pt7zAsaocT
bd0b8sy1wVdLdhUf/nN00BqYs29xIfNqq6pHg/L+QkEGlNXymDCI+TmjdzYGuKUT
Fqf6eK/BnEqOWwQAvTqwyecXHsYiv9pTRqmq+f2xK9xlgbWqD4pAODWMSTRxPduQ
94K+BsZm2QfF/G92qf+pE0XiVxpjV2+UHZt8hgH5ErsGWpzWjfou9JWTxKRlaVh9
hUwY7wWC6DBhWVMfTOCBtfT3gdnxtDknyzr5isv2YcbqnLI4Ql2w+n3CB08B3Fva
5TzKv1ATWB6cRKFgmYNNbsM/UXN1dgEvzRcfCQ+VOcctqWF8JJzAkDnMlHevEYPb
iKodd0BeZeQwS/S8pO6CM/yO0+59oDAuXVZ5+Psdy2VEf04gJxM/3WLeOqmK8CuR
eWY6s58Ts3eiTxk1TX+upFp5pMYQSzCcWEi8s9kdtyP7j5c7K4QDu95fwXr5JRzw
+BZTAvUEyO+/I0wMWCziAbAaGc+sBoWOaRfW3bRhacUSb+ncj2V33Cs315gGcIKU
z+QStON0Yc6o+ZL/cOTFes9Cor4Yi08f3cozJ7IXxb9eGR5hQtlQwysHOlQZjZ7K
RjBAfYn7dAoANFWXnrsVPvlCrTki9lyU+MYt2C9ZdSaEw+Fibdqcv8tRV3yvvyfG
hRIZEuSAGtvMmqtx0iK4I7Bq0FOvYIjszh1qwkOEgbUbNJStMPz/nNiuJvtaVYf0
0l6junOEif+Cc/UY2xvWDrGTMtYusUnPJnVwFJyJxmlhZOK1vldoUqUYNnxofvhj
KflgVcnhQpFhncmUWGF7MjN2WONnADBjkQRPTGyh3yXQCrH1JGo8jGizAM+EtDSX
UDyrQbG4dBg7E1vyywlojwDof+rQQqBZl8MIRCTqNf8ka+ekwvsWNIFdEuilwaov
ScAYdU/LRsq3FOSOJWTvUO4BjwJH72qGhglAPfPCKOtsFXNikZAmCXo25Xg6QZGB
Eh7NbimyYVWvBxCb937ZtIKRf+ihWPYswSOY0ZjuHgp8dMyRfH44MeGetsYfgj01
F2qxbQIgd0kVVztnAQ8BEMzwYVAL6OZk0ogDbBXiGUnlarKWC6NFy0Bz3WIu0NlE
2OyTXhGYvJk7xwf7Z4dYpZpbK4As+4UMI8CSNXQQis1xFTuyCGo7tl3RQY/8+5eE
RHpxnqFsPaBdHyAlcDUuhVqlPLjUoJPtLyUYpD2ts8o0sCNgnKU2vgGbjtRc37US
xoXlxIy46c7JgZ40vYCgwRofOQIHB3j8ED+qN7N2ZRre892yd90+Jqe+lDlM22By
bCU7S9ksOvbhoX9InTnO6RpAtn1PBAKCCRDoLN4InqzOxHS8mkbjjkDc/H7QbOW6
jdQUq9zXwSPsoA+439MWRYVHF+xqvidJgo62frlFsq7/x4xnYoJTzvAHuVbpAYc1
n2EQSFJuNUcDwx8Ln7Ip3nYNS9cSzydSQDoT++r9qgE7iEVwfqCcKgJQ/D/BaK3R
SGDr0pKvK5DXRnn0lYOvfbh3eUUuMMcjL6sYSIVCJK4eQrAUgY1txl8gkb3U2yks
U43K6q3AecbnARfwrAPL7WreX/ReoXq76GH1D5f2cbK2u0IK4V8Gi0ZLRjtXZT26
UsSG/iV3VGKakxRUkIxTvq/uveeKMTXIE8g9zoDs+A+WV1Ce5pRlaOEuvEJjIjwH
v3JrEf5TyWRh/Rr8mtMz+veY249c7T1eEtlQbVU+X/5GzZcNxUiFXVQLfOvZVLCl
j4HAoEMTqCpeaNqR6J5wDJpOWVQaMQo2QpRXzmHlDh0U6EmYZ8DW4gE9R/PsxG60
zj6X9Bj6AMYsxUF5tZaQ8BQqfmEn0pWvTG5k6ZO8Wig5FhqTSVWOzKdnNw5kPMew
8IPzBUX0OxH2F0WD05OieVhsK6cGs4wtr1y5nlHIi0gllQ3fxTrY6EomFNS+bz6Y
e+6Is6PqfoUSwRVWDlst/1A89Z3ZySHlfY8bTsFo92pYgUc4GSK+I4lWqoFpHKmh
5UmPPE0+mgPpDSnSNtgOotS2KHNtsZBZTH5QnaqfRz3VJOV6xv4ccJNUT2sBKkT8
`pragma protect end_protected
