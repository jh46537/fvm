��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,��F�X|�ע��R$�O��I%����n�SỦDūrnnS#';��^�?ēW7���Ahu��:��*4wj����¢K�0L�N�)���Ɖ!���#�xJL^-�I�Lќ�������0Юp1*/0��ɜy��r?)��&P#�&PBC�>Ea�w���I��2��tN3�����l��;0k�y�$��55��R{�iv���{�!�X�B��n�!Ww+�<���E2ɲ��4���K�6��	h�gx5M��ұ﷍e �G��X|�ה���l��O��t��l��)'FзZ���A�3[�>�����ԍE�vUV^�U��{���0ȀjK��N�rX%(-k��̫?� ��'�a׃�s�	�������I���/�x�(�x���h| Q���Ǭ�x��b#J�-sS�;��i.ט�N����I����µ�F�!))�;Ĺ� �2}�Z�H߽�_=��FK�F�t��uSf�^]����V��,Ӥ���R�O�P[_�)Rs�Js��=B�g[�4x�G�0$�>c��/�� ����r�*L-GƮ`��<O����֓�ӾJQl�KP�T�Z����a3��ƊU)w��Yv��._\�	D�y'��Fɉ������xK8���t��D�\ �����Z��`�giN�/��y����yxƜ�9akI�S��k]H�b���f1�ߌw"���̨�c��!NƝ>����
E��uE�ßL#o}�p�ܝ���$/o�-y��Zl����l�Qu���S����p�Gұ��ؔd�`��N��AB��������ߍ�	�u��~�� ?���
G1��wBi1��wiu�Z�a�bp�e�}��f�����w���3�$��8i��;�c���l*3�<a�����p	�](���t�����@Y�"o��go�=�k��%I��h�޼�,~(
A��B
���k��OWx��_�b�G��g*C�;�7E�a��Ry��o�����Y�q�Ӵ�J�Ɋs�q�\�
 �t�t��攟�M� �h(��0���;�>X֋2�?�E�D1��O=4��3�k���6Y�y.�������x���b=^J�U9���+0ml�I�d�������~O#GKK�
����$�#y |aHu�KY3�@MBY���x��v!��K������~�w�<�ϸ{���_��|��5��g���W�z	!���-��Q�ݗ,��8N��s�D'K���ݯ�!��DRpY萶7�J1��5�=��0�!ͤOf���8�b���|�q�9��B��^$��N!: �a�G4{��:��M����S��-R|�~��&o[{#H��~ȫ/Vg@�*�d���H�]��3�'Ůj�(�`Y=~�Z�"3�7̜�.�Ӝ�9��޲|pd��q�$W~KkO&�Џ���zȷO�8�^\����+$ct;��=�SNU@������+��CK ���@J��|l7^�$�U/�#��I�cPг����J�ul��G/z��+���r�!.�f�0���_mP^R������DJ�S�!�P�J3^$40	T��W�G��E�H`U�Q��!A/��[���x�%:��O&��#a�V�m����ח"goڱ��Q"����v�q�A�����C5�$�\~�,z����y�S��S�|Z���4y��z�}�t�E���7H �ԼH�G㗎��8�t�t����9�{�q���qH���>N�[��^��.%|���! LǗWP������$y�	���ڛ�/uD~���������@g���<��^%�b0��m�8���d8���۪g̔%�'��.�G�7�p	�*�8���$�5�#i�Q�6�˹,Y55E��r���Q�T��P���^����D�%jςD��
g��.4�'��HQ��.g���]-W�Φ/����1���'�>���c6и���VM�{�O�y��k�����qq�����g������<��Z�N��C9o�]Q`�����XÀl|�n�;�.��h���N��{�S��G�TF�s2����`��8����B(U�D�U�"K����m�ԔY�h�
�7�5���ˆ����9���nlk���#"� ��.�����W_���Ε��JwQ�����U��,� ���'�m\ ��	J���N��x���5�r	��-5S��X!Top�3Qa�1!M_���8f�fu�X�n/�v���s��t"�0,��?�rZrB&��hԒd���}$�ɩ�a��L@D��T+1,��Jਐ}�2��$6��#��D>�<IuaƄ�.>�o�v��p��O�2e~�t�4|I�������
4d"��i�$���9
���-��i�$&6�3�KM4u���n��rL7��_Eu����}YA��hKE\�'�����g]h��T�S$X�/�)>FF^�+/�m�JI�;Xg6C�ck9op^	1��q�!	���/��R"�tZXc���O�W�����}x�ڼ�~��� ��OC��I������B��"�fy%ԉ+r�}�;^r��q�{�Yz�|��=���l�ye�%�����%��(�����Q ^�u�>.�Gʽ��(�K�9��Fki݉����f?0���8��C�iRaj~�b&�pC S"��@�&��e�\�l��Ԋ@<`9��!lA�������tUl�R; >���o3/m(cTUA'<.@�?�PE���k��Q{��y���J�)e�e��u34�~ب����6�