��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B�6ƨ��J�3��yq�&O��e��jP	����a������Oix�R��k�(V�5��lE>t[[���klFb	�}�W(>6N[w�`�6%x �o�)�N%�QbR��V {�h���y����a��΋�J!vo�y�Z$f�M��7������է�O�����׿lxV�
�B��PČ՟�=Ї��ղ�S�O�x�H���Bf�43�!�+%D�VW,)r���='(�f&��"Ig0V�>h��ae,�q�#�G0�֭~��d���M�/!{q�ѥ��"��7��_RD�����E��lv�`va6-��]�}lALyv�F����G��|'��bdo��~Kk�*�}��d����:����9��0c�Yp�� :��/�E����^l��c\-�E�"z5�f��+/N6Z7!'�?N�)r ��.~��6�?���`��[�^��5��
���Sc5���o����pٚ(kø2�$��5]$L?�R�;{Ι�߉*�vhVZq�o�ܿ���]������7U&S�����<�m�b�Q�ƄV)h;�����G���52,�����㔀�O⣛��u�?N@���4Ϝ/?+LM���@�R<��z˽�$;<B�/��B��R���bI8�A��w�W�J���B�'"r�o.W̡4N1�[�_8\u�a �gs�.�qOP������o{�&L��w�m�~\
�#���� :�m���?S����wb#l�.+�e�M�vX�:Jp��l�M��B$j O#\ĩ����u�p��\ԭ��P�ǘy��|l��n�AJ=��[(�Y�"����D�ީșП���8$� (���[�e?#�G�96��������u��Z�95�5V�R��:<aK���g��?��\a:=B�X��B\U��)��&9�)!�ν������嗥H����1�#�D�8������
^ ̎��\�i��&ft�_�V+�X`�R��>I����7W5�xq��D ����>|� �5�j.��n�s+.��?��,���8}��_�1��?�ܶ������`��C�P1��S3gA4�D�N�����^3Ǣ�|�g�u]��)�����S����0�>�)��_M�f�%��s�����]N�N�m�v�!Ƌ%XgR_M�k��4�/USN>�	�I���:��	�cYQ����X�x6i��/z�S?����A�Wo';�ɑ�ť�k�>i����;p^e���c�i)_)� ��5l,��Z�ah��nr��CZ����L�K�p��e��`f0P2��DNƵz�Q���uR8���?�>��l�m���C(y-d�G�}���$Z�a�����_�
�b�Rlu�ֹ�6ɳ��b���3��g��J${g����g�m��m>c�~����x�a�&<�h��Ww��X�B+�ClC6
KX4D������nʭ�z���t�S�:�;����6 �7|Q�*�j��b3������*V�s#%�p���uK�w9����r�U>f�@*�$��#v��3����-�!�\�9�pv�%K��9}ٰ���Mɶ쁥u���_������k�G-�� n�����rzc��V9�kK�50�|5~̃��F��`AZ��������jb�ጌ$���H �W���A��*�C�ҍܘ�_��N;5�Y�a� �`�*3i"g�������� ��!�(;˂vZ#oX��Ai�zHy�_PN�\��i��M6}�!�MF�JE��Y�@:��� ���^��k���˦~��܌��d��h�����tԿ��AH_&�f[�V�dz��r�敗v�h�mL�y����2���|=�/�CB�b���n���+���
�:c�'�@��{O+�d��yw���h[�·���o�*O3K��S��ҥd���`WH��ӣA2�a�ä!�_{���ݻ}Q͛�,�/F����}ە�*�8��َ��s+Aٟ�j=�<�5Z��=����Ul�r%X)UL��)4Q�k�읨>?Mn].FOfngg�7NW�~��V���=k_G�٥{���D�m@�#���
)Pp���t^��c:�11��X�C��HU%��U��v >�Y)�Q$১%�0� �5#`Ԋu����ڞ%������+�*B��%Ǟ�'����C'9�aW�(��hyq�Mq�#�>��v?q8䥅[$��[��G���z.c�[��ڸ_�2M��t�jJ[}�����#�<I3��.�q2=�UZz�N~:�)��{eT2G�1����Vz͕���c�e��
h���[a��*HP
A5`�+�f6_��u��:-#�A�֛3)�������-c�)p����R�Ӗ�y���;���@cd�jďFy﯋:��)J�B�C:F٭�9 Yә/r��2���% ��\�h�	�|������#�H�R�IiW�G����;����"0z�n(�)0EĪf�:�h�#�b@*�lU�[��Bdҽ���Kӟ��B���#0e4��!� ?�����zn��͢1�cչF��]�9	�(P��!�
čH"(�/��Nc�a%>&Y��:��`3-�mR+*2c9��z��K\Y�z���S�����&�X���ì���=q�l,�@L!P���`�uՖ�CG�5'��Y�[��=;����Be)�,�5g��w��	�o,O�P����+p1��DJ��|���I�7���c�% )5�|���(�%�抋.>��%.#����a��w{_�Oؿ��R@D*���uq���������}�Z��t�@6���좪��;���h���̊�q�dyq >��S�[����Ud���{b��!��G�y;����v��i��6�=���9���+�oh��~�ad@ּ������7�-}��Ԧ!��G=�3�[�C�a,�IϨ<-s�d'�i?N��'�j[�����Ix�X�8B�R�PY�>��u����ӟ�g-9����f_��z���� �����9Z��B(���=�(�K�Sj��(�Α���l�X�^�
!��u�դ����Z,5>!~[{��@��:��IΩ2���y#ϸ�U6�X�D���&�����`��n��)봓��E���j������'<�d0C����]�� �e��s� ��aQ�U���pB0�D*X[,I�Ņ�S�F�����ʴKE�-|���8Bjz���p9���*���}[����k/��<x���N��ޗ�t�K!ߩ7��;��W4}�W���g�l0;Fz�A�`��7 �t����{΁���4�u�
��<�\�ϯ�������2_0���H4���;�uTe�#�����=%n��ó���A��wh۔�K'Fx?�ga�du$�	�����g�[���3�\(F�z��j�װİ� ?������M�<~(�e@)MM&oD߮����hr �<��/F�f*���%�`��p�|��4�NB�Pw��TU�(��_�u����騪h�2G���߾�<�SiB�����S6KW"�p�y}w�O���/@	����]�o���?��my��Ļ�p8�}g�G������fC�k�25B����À���Kڑ9<A�(<��S �X���lB����}��Y����$�b��&���Bs�G�f�H�l��'v��{����yg{�h��{!�g��v��Y�����N������"������!���o]>�Š-%���6n.�����-6(&���֊9��d
ݼ�d��'��IS@*�2���n��x��T+-�o��Ƒ�	}[;l�:J� JkV�zl������X�堾[��IOl�z]Y��qD�^!&�2��*�Q���#Ϋ�М�/Ι���be�j=���c@
gE@_�?w�)JT�/�'\p"��JD�o�ٿ�pn�uY�2�� >F�.N��<Z�^Jr�(�v�1��uk�uv�J��l<`�n��>3Rŝ����+%f�l���:<?�pj4�eY�V��OpS�b��u�^¸^�Y�&��&b��`�:�y�z��e�ͧM�a��Έ~��G���x��)�F����~��9���>��@:���y(��dV׼��Q��J�/��͡�\�2-dZi*U�1��,�D�3�<�r�JL ��@�/t#=��6�+f�_�x4�H��i� r4�d�����r��d�&�蛾]Z0E�{T��Ņ�"L�b���D�e/Zod�������~4��wf��aC)�&ofN�ö�s�C�y��J���@��V2����u��z)�wӊ��t�yR$yz:����O>����C�������>��$ ��ǇW�0�ÂE\�4�V⎴`�#C�=Z�ϡ����2���%&(W�+��֟O�C�?%.��/��{�H�>��Ę��5S*�-W�<L�hm^Ҿ��/����O�Ҕ�9��й��kp�l��Whp6����%��Cа3�V�#vtjFB8��rXea2�ܚ*�4lP?�\�90R���վ��J�K���a�U`E��Ȉݼd��3⨼��{_~C'`�Z�3h��Bt�|�7j���'��[��<��?ћt��0��f�m^T�)~4��	�'0��
ۅ��w�ϬP�amNd��y�g��ɬlS���
��Y�F&:�E�Ꞿ������;�����-b��Ujd�?� v@�.+V�'iC����[CF���(K� '`R��"�}+˭��o���ݯ&�\!y�����ym^-�4�^�'LP���sU���	�O��]!�B+]�QCvW�18>��q��%�M"V��v#f��qGu���e��o5CY�Q����Z��#�H O��v`�^!�6CCt�q^q����o�`шS��U��87s'�&��W�6��M�N+�|��lФ�asg����<	*���!B<ei��ީ>�����T�H�����c���l�������K��8�V1r!�'b�����ɗ'���gJ��?� Yʹ����RBK������}����	��l�g�Z�u@��)���/����k�	2��w�r���F�Z��Z��I�}��K��r�h�<jQL�=p�z*?��<uGt^U�`()0
;l���h���J]X��af{zΕ>���4�	�v RFe`�ћ�ש 巪y]P�&y�a�Du����;����9�T��x�A���wBZ�Z������,�|��t�iXG)���Tq1�?�g�0�c�c|u6`\��Fh�I�9a�C?��x/�)e����vZZ��ӡ����	��|޷u���B�.m9t���7���gr�����&��7Ww1�T����m]��5�����,W�ƒ�9�_ZGf��+򴨘�ˇ��3�cq�����e�[�|D�.�BKR��'Ớe\��<�q������Y"���(ukk�\o)��ӄ"y3R��]���K����ƞzO��$Ҁ���x�>���p��w	���3�^$��G�K�Қ'�+]����<xt�l��TD�K��?Θ$tK��,�+��<@�ȉ�ݞ��pۮm���Q59�^nQ�m�J�)�4����c��s��G�-b8yF�Ebւ�ݔ����/��ci\�~��m�MڗxTࡱK�"�<RH��h�w`�**�7���� m�s�~�f4�E�)�#x���%[� GE"9"�{��;�7�<cu	� ������8���z�Fkr.��6-�]����*S�}?�����z��|�D�����̅���uY�n6,���Dy���׼�x�����钮=�Ca�b����pt�U��\�{���^�/t�h��2����d�0�r�K� ށ�q+�x�,G"�
a�EkХ*�#q�6�I�O��k)����K�D2���ᐖ������ؙ���
�Iē
WFL�t�����X6�����L���I�銅f�Dlg&�3�xӏ�l�V��0�y@�Ż�`���Y/�dC���=��<fHlL,~�N�S�Ԑ��bդqR~Z�� ���G���b�M�'�孓�%��[3�:<`��]Q��D�[J�=�L?��IT��e�,�8T�i��~<[��{�����]����V�)Չ��Īձ!vIh��8�KJ/�N�l4̮�䆠���K�]�K��YR�,��|M4i(MTh�lDd����5ڶ.�STN�?-j��>�mk�Fe�ӕ�v	P��=�
�ゕ�6�J�}��gP�
h��G���w�c3�� 2F�9K-����rg�wC����N�k��L����M��m���͂�V{~�F�v4������s�<F��<"r�'�`���ׯN�x?�u�U��+�2'�B�6���{˽~���h�rS��0!"��<>��5/����Q-/Ş�g>ԏw�+��8RS6猊�#�e���/^ƓA��D$� �A��'��Q�x�|�����юTq�҉�u\ܖ���t�4h�Hc�x�1�lw�V���S��(��n �ä���2hUf���^�}�� �����h �M�_�C�P�J�>��Wq�ڷ�L��;-7��{��ﵤqڵ3��+���W�o��gn7�U(��Ǆ��I��̉fR:�[���|��Ȟ�u$�����;��J[%Bs�s��1O�R&5����qj���Gfp_:�<�wܙB[%�P�V�'�'�NnҝTO؁]ǐK��:9�ڶ�u��(턣�*7+K<�˙���$�n�9ѝ�!+��DՐ:����l���xr��Nj�.-��Z8W�JT�٢׿*yG�mMLS���>�]�ܝ/z�:ZuCѸJ�u�Z����S��n&o�5	��p��Ɉ�6'�l����}n�@�n&���7�<ŧ�O}��ԩ���N����E����VW&����-�"e�7�: ?�Y�C���Q�ۮo
q9o� �b��G8�Z&b���#����:䭟��Ă�@m����� `ȩ�Q�^�?�#�����P��c����z){R6:nB份M"迟���˰�p_P˅�?������j�{u�ܬ��ŧ'ۄ(����^*S���Vv4Ѓ,�~'{����8�F���xQ�/�K)z�3�����0���?W)�'�	�QF�)�נ0�ߊrI��kDh�i(߫���(��2�ύ�S]02�T�3�旚$��-9N%T�I�P��� ��N=�͛%.e���l���kZ�s� 8z�&�5��Q�|`��k�#eG��nqM� �l�}�n��,�e�=v��IY�2�-�D��D��n�Һ�+��?BD����:�/T-�x���IC{*����bZ䖤i��6H#pW��l�X�In�Q{%:�m�I0t�IDN+W�������M��_�~[��Ϫ��Ƶju�S6��va�J �:�tL��ժڙ���=G���A�Dؖ��R_��}m�Y7�em�9/���H�)Pҥ��W¿bS�ǎkP�m_����$U�a��o ���w;�0��@� g�8w��7�y���TY�2N�sy��|A��C�,�֯ېIA&�!�J=���%T8�ߘ�k������?ir"@�k���[K�\XBu����f��9B
'םH�\}��a�w8�_������K�Hx� ?§���#42�p|�'66��Zp.@&W=�]��qn=�����,'���� :|�0���б�Q�]F� Spp?|Ml���Bt~stiԿ�G�ш֯8D���0\�|7�Y�٘��P��֯����t������0d��]2껷ƕbR����sV(�����K}��ĥ*/�����"@7&��o"���	B/�|��`�Z�D��;x!Ū��B
�ci�f���u󣟻���~�j����9u����1���	�����d�#��� wo3���h��������jkS"�h�`#c �5���"����pR0��t��a�s!R� fΡ��κ0�?2�Y�	�"-�N�o���n|�r�H��<W�=Nx�$��BL%���䷑zo��N�Z���?��&ղ�x�k� -��x�m�1ߑO+~�F`m|��Z�Ph���淋H�[F������Jx�?!0�U�qv.����i0쌶s3���k�ױ�}a<e*U#�kn�R6F(l�\���KZ������p�X�����w���4 ��1X{ѣ��"װ��7��3<�T	�o�6��nD/oX�>��W���hZ(vB}�0�೧�4RV�R�~��`$�v�� �r�M죵{���Q�=�<fS�-�M����k�7�WF�*]G�+��t�g_j���U
+j��c��r��"��d'#��ѫP ��T�}	N:�}�bC{<G�����R�B32=�2}8u�1t�U�+G<�(��M��
�x_rׄ�-P���㨼	$�O�g��γ�|��A�U�>���e��'@~��\�� ��El��[��`����ƅ�3�x��������v����@��kpx�1p��x͉lj^���_�z���e���cy�k�[-��hÂ='��H#�FV*K]�޻mG;��x�I��/�o�݉�T,Oz�o�qo��x0��b�� O���2xl�\��l���m�PT��.�x���5��� �t�"�w��F���@j^q}�#R�tH�7� ��W|��"�!��w���K�J�ܖ���Pj�JDMޢCr�8�;���D���E����U_�p�h�!8&�<��q�j��&)f�����~��� �y��`���5�?m����9��P��T}20�Mw��)��Y�K��������5�E�#)'�٘d�}~��-��yo~��[2����.#����Z�Q�pw��uL�����{ٽ������*��Č�dc8��!�v�=�[�n�����^-��N���[�Z�L`���3����:����A��Ƨ2{�����%��H-�t�Rb��Ԉ؂L�ש��Jv�`�����*g=V�T�w�=5��Iޯઠ�[o�¿M!&y>܈c&|��� ^ L)v�)i���/$˹��^��t.ш��6��aN�?:��0Ϯ�Q��>�ݕ�>3�f;�R�{�A8��b��Z��5�s�:��c�b�;�E����4BsSG��Ho}��Co��a��+�&������̑��ICp{�cf�p�U� �焈�n�?�G�q��`2�Yn)���&`g�D^�Kp �U�VC&�ۃ�HG{/y��8sQu6h�D��W�F�0�-)�J�ANzQ��kF�+�#6�ĹN������D�^���y')�(e��%��>�1�R���+�eJ��O�#�����c+�]Au��)�_%\�z��D��������]c䈈��/�dd�n�!���ꥰOw�%Zi����GeQ`3�i-Sш�g�ެ�״o։*T��E=
�x��D�g�vV�c/�����Ϟ�ޅ�W
�ن�@�����~\xAؾ�(�|зA;d��M�β�Qbs��$ ��N�FV�Y��P�jZ�W�9���l�:3k�-܏{�|�l!��==��/D!���jq�Ye�'CG���5<��qb��͗�<�>����$���V�ڦ{�N߂L���c���� b�\�^&�p��_Ȱ�ڌ������I�ƒ��jG@-XV�au{Y��������g��%�}�6��PD��Əy*!�T�A��'���ǆ-�uh��9�%]�W�e�M�U�=X�#3��ڮ`Rp��o����/}u�՜`���!M���e���Gk밦.�~GoVʒ�ʆ��������TF}#�!ngA��2�Ո�xg��E�L�iS!�d;�L_L�rr��q�M�`5�w�����y扐��ᶿ�F�������m�jQ�9�i�9Y�C��{�j#���?�&��}��wzwg�Ś���ι�sG	��Ew9���	"!�E�������� <������
�_>��b����[�-Ϫ���J1����ir���nx��b��9�W���}#�.�Lb�����	aדI�XC��݅�:V^ZL��U8�7+���8�uط\[	�們�#}��&��J/9� ^[�t�sy�*�M&��CN��gӬmx�Я����'�>��,q�$�2�@���m��T���Ɍ�m"��!��n��V���n�#\��Sl�����xq��U������W/ouwK�#�E�B����{f�P���Tk��|!�c�TQ�E��|�2&���^x����=���+�b����R܏�&=O0��n�b�2���hL��o,0���,E�J�T�{�Q������K78sr`�U�K�F���Q�W�t.g�=���y��t�m�\�G`(�)ys��9��x%�é9��!4[:5��]�v�� ���9:�h�fޠ�Ū��Z���ʱ6�8��׷�+O*��h��r�06�h�@/R��|��!G461>�� ��'���iCh{Y�`�$��������әr�D�b؛�-G��������7��uV�P�?�L� "�ʙߓ�*n
��I\�S��1j�y�L��h�n�w��j�j�������i��d;�O�V
uk=����\7�v}������rw�����8nGN����E �[����,KH�иz,9�c,��?:�,���T�z�	%%��~�C�Do2���S�T��K��g����#@�[�h��Rs�2\#~�I��<�r�'��W|��^G�
�7m|�lk�Q����c��;ð�Xv�ܵ�:�$Zc��z↙O�aO�tt>6I����ܐ���9k�d��oC���/B�?��8�Wsd���6����u�#ԋԤg�G�ߝk�H<_|�o���C(�TVJ�E`��@){%�ؘ>l_I'I}<HEA��f	ė���p`T�,�#���d�<
"t`fr�9s(�b����;Pܰ@[����
�N�<5d�I��;	/����:w���ư�c�a�!���k��]/�%�Zg:��d���j%�L��m��m�wG�\`Uc��i�i�pu-<G`�b�nՠ͗=Ȗ����\���	K�	݌5�^���3%����&V�܇*�Dd��Q��θ�S@�o˒0�j�dy8�!�6S:��e\*���a�g����6�S�b����hW�.?9���8>�� 
w����%M^��A�(G(���X&�DY��#���1�< ]�fV8�3�9��I�S_�w�lR���o�����&��R�B����@�Dh̵�d2��e�c&L�ٙ�A�	H����>�.|zBp�P�E���M��Bcx��3��E`II#'ܨ���f���u� �~�������p7��C/�gX9�w�˴�3Sr �ɰB,7�P��!���AٍJx��t��D���82>`��%�8RZ��Q����Tn���8�m�m�A��c�iV�&f.C�L�7�S���:1��s�y����r�"�x?n��\W�� �,�����Md��7�	�=N�j��e8
&��}c�°�x@%/S�jR �q�xLP����bɲ��������"�"kU��I�ן|I	l0@�R��)�"C�?�!ܺb�W{�8��T���׃s<R�sd�����!+h�E����Ц�3�aF`A�	�9Ӊǥ�֤���}�.	� ����'ˉ�M��Ң��þ�2d�_:E>������C�LQJ��\���UwUv��+Y���4 ���*ľ�<ާ;Y��9������T,mĔC�ҷ�2��+�l�o%���V���l0qf�^;�9?�iʸz7Һ~(@H+|3&����A����3ˆ����(�s�}{tlܺ�:�|���1/K�G'�f��!�1�_�3Z3w���Ć�7�� �����%�3�� �n�vg�K��~�!��5�\m]ܓ�0�OsI�����Ri����l`�g�SBX��Sk��4.��]� F�\���{v4����n�4W��a��^/-��p8�^�p�E��v�V�p�.�����t���e(y�z��3��y,L� :k��Ԁd��[��7T��o)f����86BO�r�I����p���̼)�ٖJ)ހ��DlѼ��p�������7��4xg"|d�IG����F =L�i�"/��5X��y]�jDJ�W��|��ʿ>Nps{9��@��
@0׮v�	������3�lqnֱ����B��xO�lMx�zC�
��_�x�DN��W�n�sg,Z��8�����m��c!�7D�w���L^���悛�Ѻ�b~�Q�[�}���3T �ϻ�X�c�!�W��_�N	���Pb<i�`�D��g��@J�����8Kw�kWv��6� �0G}�W86��?���F
�9y��Ԑ�߿|�I��i��0�Se��Ɓ: P�aɴ��Tt���@@��������2�~}=�U*�����X
�A)5�����D�Qp�0XYp$ �����ъ�#E��1l�,l[��lK�E`<A�!Y߷s�&�ނp����g��gg���°ο���;h���0�	E���"
H�<Y6��f���$P4$)N�Co+�g�&���t|���&�.�7��VU%h���%������X��a2¶*��(�����
1J��v��i +% ΢��v�̄B\L)xf3Hw$�c���S��&$/��2��b��C�b�����O�B�=����TO��M,��Ri0� c|���_v������*��� - ��3b�=k�V����H{���<�u!��՞	<
�2H��C��f����CG�"�Uo����aw�0�{_?=�ؐ*JU2Z��"�����t��o��h�r��޻s�)��fi�K㰱S�o�c[����Ӵ(�i|�T��b�ҿ����l`�+�l}5��|3��.9$۲�u�=�F���IǂyD �5���rf�~\�+�����h7"7aEԗ~\!�ν~��]I<��hN 抮{�pe������ޚW��f� (}'jl\tRb�D���
8-{�|}�&}9NV�8�����B���
�Q}����j`�ޓ��{��K4��8܆����qWE ���%� ���,;�)�V.IY#���Y���{�B�9�\K9�)��t}Rp(����ff�|�i|���OI�[��V.zuX(u����j y����+���;"�Nt��L�ƭ8�>�n#4�T���c�F�	� @l)� ���/�BB�
�\;������ R�!u��A��J2��ֳ�W�w���TaPĎ���T�6B_�a;�F�2�Z�ۚ2.Ev�T7��1���>��!�#0��@���yC��d:���5[�X�Ϧ�ۻ���fa�!䆟��}b�A`��C��ʗ,f�M�Mh?&c�L�#��9Y����H�]����D
d�y�P�z&��y�ɼ����F����>]Y}!ili�~ �Ve=��j��������U��M��7HY>�m��
���$(?]<�!�4�����P�����	��ݏ�v~)�[��ʠպOQd��\���^�Z��������mfjQy�;!�[���Ps��P$΅���9&0�iJ��ū}���Ê.�B�ľ�R�r����ꕆw�g�oy#�Y'.��E�Z�A���оT� Y�D.e��_M�ԋtl�
`��	���������k���	W/�z������Yo'��G�t����}�4>-��<��BT:�fmN։Rb}G��uA�B��2
R�N����n1V���D¥P0ɯ��	o�ʨ�|�y�}|���P��Obb��@E��(GRh�<���^�N�U�ÃݒC�"ׁ�g7��LDg�
N�(����Q{��Z�F�����[ǖ�)�y.��H���V�뢣:����m�Ea̛� �ij/;c�����!P:���D��Si��&��G�?<����	Ƞ߀.�ێq�=x���!�D��������	:K���w>>����)����9�n^_���.�.��(v�>$�o�5N�e$+&Vv��17'|��&�uK���羈��� =bz~�#���%k�~˦=[��;�UEk"����$u�an?�ɪ2E���(rࢧ��,>s麡��;a7�]%��km,�W�
{����1����.��U-�V�lZVgo�B4e�2��-M���1�?a.\}~
��ѱ�d�!�':��x �g��3a��n���#8:����u����>�q�%o��N�V�V;��㑉c�r�
,��CNg~_�[_�&�I���\�B�B�aP�b4(�݊��Hgy��%4����z�;y��\\��@Jh��''����M}r{m�4����A"=��h1
�@�12�M�v��|�q�O�\�����4J-�խņ������Anm 7�z�V��~}Dg��ϘV����������"�m$�e�bJ�r��N�
WD��%v~��/�ιmQ��CJg�I��]� �FS����%:{��o�"w�,`��t}#ym΃��0��O���Ԥ:RM��7ؠ��5�	y�)��ͻ	�4�����M��03k��w�Y�K���F{׫�KA�Ȝ�BLK�L<6P��3^��f?pP�%� �;ϛ�R���5ɺSb m�K��C��?�㗛ħu�@��=�ca�H��Z��BS�CBg����I���_H�!Wd@�����R���j��p#��Yu��e���ڡ�(k5m�ß�p�+>���xa�RL�Ny��ۻ������v�v��5gnv"��#й{Ǿ���Q�j>�D
�.�ߝ���1��`^��mW͚�R�Fۇ��%�|���jx�(�:�ժ���#�Մ͝���U��73|�kOc<�u���ٖQ�������\����$mY��o;>���;v5 g�x�e��a��_o%g�|��}X��uQ�;�����N�R�ʻ��ǡujۋ�g3���=� �����=rM^�`1E�ğ�\|���'�%m��W6S[$.��Sl"!<,��UP��D�r�����Q}�D�U�����g�rIc[��8'�����#����Q���,������%`��׾��c��s���	n�ry)�*5��A�z3�"x��߻m�d����xȿU+s��`�LX��0>FƄ�D����d�(���X��+$E��I�X��$v�>�����r<��xi1�DU�E&������.QJ��ސ�^�����v>q8����p�-��#y�v�E����R�����>��Qj��Nߐ}�4�$K�O>t��4�򱕣���D������6����B趄������MmrM��M���7߇U��L��i��a9W���rD�n�,d ��/ �𴁈�P�x��=(�|C6�V��c\jv�_l�9x�΃A��H�f��=�m�"8A�@��M-�c�a.�ɾ��������)�t�8�gVE��n,,�g�j����Gԧ��)O"wB݂Rޟ��)���ݗJ��?ez�?��|�<ƍ+#��s_�Κ�t������H!Gw'�|�ǌ��4��f� 
d�KRG���A��u\� �.'g�EV9��&�'�ӎ���f��z�(u@A���0�����-�;'0&~U��z����;{�D��A4�T�p@��@23:��N��OqEm��=�:��aB_�������j��!�K�)D�I�ai^���>:����.|246��w�%8�I�!�3�- {UPp�ͺduu���ǖA+���'$D��Y-5u_f���DƢw��4)��N���T\�3һ|����6���H��a��xz���g�@�[���M���N�3��EU�@?���+f�?�a��g:A�I`���O��I��e��g���ȡ��m\:�&�j������G������G����v�*��-�e��b���]��x�Ћ���9ͪ*������`�2���}��8�� ��pN� ZR\�EdR��F��H�ȍ=	tH6�H��KKY���,��^��S��ws��������j�.�Fg8��e3����M���&�h�Uv�G�J}kF���cw�9��r7���w�'ʹ�:g
�V¯B��u)\�g�Dsu͉�qbm"�P�� 5�0�@O@{3� �ls�"T1⹚�ĔZM��c��:6<�y�!�#���Wz