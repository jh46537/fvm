��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"��Ia�W�� 2Ch���E��ʡ���U�A���1�%�%<\!<��
��l_�؂��8Nh���-�:��y����E�����!c����-�Ea8�d��]��m�D��#���6����������=��\��]@���0/(l~��&JD�'��I���S�^zϼ?��o�Z���rx�p��Nۇb�k٨�)@c K��4f���� X�W�P}Y��B������_&D=�8P8]%ifXmZK��顄5��ϊ��� r+*kʀ��\�h+-�tG���{�: PCf' s�BϗVFT�U�vS�����p�N��F������D�Li�V�vu���qr��' ^���/��lQ ��ż�f��kW�z�i4 ه�+�Fv+�1�S�1I3��d\� ݜ�Z�� F��	b��jMώ_�uaS�֢��$=O[�*ko���J� EsɌ����^w���fc�A��=��p$ZJ�u�l�;�2��Q"�\��0Z�]��5a�d������j6��$���Bai�ת���x��},�B|7.@����d@k�E�xM7aW��s����?���,��7��u-m�%��"-l�-���(����y�*�0�1X�W������i����t�]�C�5��Ѹ�0�t���*}A{E�W@��H��17a��KDJ��b��{����wU�d�Pk��ښ!:<b��;Y)�}p;�i����Q��t�'V�(D�O�s�|̤IF+�]�n�%L�,�Wl=��Gц�9��M|����{�!�k�`1�,ڱr��*�m�8���ΰ���i����o|V������ VG�BX5|�>�w���P�6�O�����N�dD5�)�Oy�	�K��@o��}�=2@)��x�q�wA.��i��k��N��ůR���j=�D�5>q���b7E0�Mz�Ł�w�(�Ԭ�z�
�S)�����-�z|%���֩.��ʰ�һ�z��hry��������?��Պ���n���:\h�����aY+�3����^Dx�D�g]�D�O��-c�QsԾ6�gg��#cY��ƾD��g�t�K��}n	��.J��X�{e�:���O5�2�1��%�d��.��h3�����9d�y}��
�j~D����`���z
������)y���uI0��TP_�1��J��F�<��T0a��T����= �&�c���k�a�@�5��^g���楉���Aq���B	RL>�<����vv�����8�X0L@�N�q�V�CV�V�P9�r���2u���e0���b�x�d�za�^��L��g��wX�K������-`x~qO�`�|�v�x/�'f<������:�u�n