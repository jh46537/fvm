��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $Wժm�5m�ܚ0�.��C�֯T�u^��k�?e�,�d�<���֡�@�:�G�vR�Q�v�j�Y����*.�T��A�����R�ti�Tf�Y̔��(k�`j>'GW�I��L��2Gj�����rB'��w������E�m���i�)f��������{&���*E�H+bY�����[�8�ڔ-���2�ֻI�ώ��ڜA-k"���6�~�U��YX1.O�*���g���\��=q��t�z��YF^:8\� ��@��Us�_0`}���3ƞ%�3?�3;�	_[���X��R��8n2-��kO�a��m����0FT���y�"gY �Ñ�
�����a�ˈ� ׋o����#8��(����v��*��f��r��*DGDK�	�<�Z�Q���)fۢf/�x�	�f۵�r����bx4�sHl3����
���ۀ��g)�Z 26�-����՟Z�m��/S;=1@���s���7��Gdʔ9jF����hÂKrA��������.���+�� )1������ֈ�1��>;S�Y���?f�\��(Y_�ەq��ٺ�r�o���JǿN�(���^�1E�U����sx"����/�A��{�5��L�|������󱍮���.@��\8Őw h+ۚ�7����^e����iV%�r�*t�Y�*W=�1����5�ߍDi)[>/Zt���h�<7�r���8��=�W]�A��4��(7��w(�*U3��u~*�����4�����֏d9��7��`��z�A�x&�bR�rg	�e=&�����]�0�<Q��^^o�X"!.h"�=a �d��>ν������
�k	r��hF��Kc�Q�fJ­�,|�6��Q]��m}����"����h����+O�L7ka�ZX2����xBN����T��b@�I�>�a��)qyPf\ٹ��a��p�����H�B�U*�˹�>rv�	�Dɲs�h�g	w𳄩mP�{#mZ�BX��=izs���
W*D�;,�(X���)c�{.JU�mw����{D��p�fW����>f�C�?nf�e	�z��*^x��wCM0��Eu��g8q%��]�U�v��C��9�GZ��~��|n�+ h�Ģ^���Mo��(N�׺�`��0En&k$���UL���TME��R��P��p{���\��,4qq���%�����U?U���P����ZsۖR'�=�wP��q�zu���)d��0�e��v��-#D�ߎS|+�03�����̿k�PWj
ɢ��j����!`0�|���&��@�WԖ[P�2�ŦL��6oq=G\�}�1��5n�
�����e�/} õ���AnT/3��I����(