��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�n�~Q��x�vHB>��碎��j�
���
E� ��6���ɾ����,��E]'7��1w�u6jX��	Ox^�f��{:��9�p3lM��e��=W�С�i���dt��|����:���t�������2�a*����Y�.��gw���Ա��ʞ.�!�~6Tmʺ��;���5��!D���.�gA�gm�qέ.Ԯpq�1�PB�[Y�jp��a��M��s�#.��R��`(��#��5����ΥZ@�^���bQd�!%��%b8��0a����8�Ɠj�KwȢ��⣑��3.�!u �"-.�ne �����l9}`vQ�H�%Qs�������G��Fq������6�(�!����kGʦ��ƣ�wl?�<J0Qn��;V��o�f�E(L��ρ=f�F������w)�V�@ڋ���*_ �w2*�x������_�3��H`1�l�=c]z>U�g�PG��d��@�=<�u�.]g���&E)��r�`�`V0�*���$�6j:���I¡�'�߼f�
e�0M
��^A��gt���֛�6�et��IAFJ�#�dT/��u�)�QyWg�h����f]�5��[,O��� f���Dܫ:�dy��iiU�8yث��Co*����X�6��l��e���Ѕ��89K)?+��D[�>�FƮ�6l���*���B!�����C�dN�{Z`��l�>m�^h�O
J��!�n[�7���tK�e_~�Ukq�^ۍ�`V��]!��-�����KEz��EM)]*8���cIR��׭&�����t�_�*ES;�߾�Q~3(�듳":Vm7��l`��������C������k���Zzȑ�cz,L���O�}�"�㰡��ǧ<:l���0��A 0j��/0,��{[����@�~!_Y�/��HHzV�������Fo��7g�`�BC�$(�Z^n{��^,t�H/����=�!Z�m��h��?�����k̂�,	Ǥ7/�o7��4o4���
��Ê9N^;�Г��47���EFG�%l';�©	|Y�Z�6vg��U�J�$V����a��bԫM��Cd�C>�?�y읤���a1Bu�S"�iN�݊ ��)s�E��2^��)(�:0�V�Ŧ�o�f�csaɲ�L�t��%G�֨�M�'+}�NZ�03��v�w� ɉm!�`�Z�܉ᖕ������N�$���e҇@Xx�4�1�����mFS�T]v�rq���XmCv!��T�+_l�C��z�E< �3�����$w��B�w�;�D��|��l��C�,�^G!*�KG�A�b��f�b��1�o�Q��ףT���$�[?HI��j�Yr�5�"�,al}�=:[��������#�_�6�|���P��u��]{*�"��*H4�_����({�	�IPl&u�2��y��^`�&�4D��/���+�[-��o-�����x,[�/]��i�,7�ln�o$��"�f�Hl-�E�_m�>ɪ�y,S�M����H��BL����E&nKDL}T�Ib2v'���w�IIDx��Wq(.�m�.c�V��[.}o����y~8@��*��x
سT�b���$38Ce��v�7�^��#Θ
�����s��wp>�Z��;���3<4��'��2��3�\�,�T�Y6{,3]`���O�� SS7�l���NE�G��{&�[�v_jJN�Z���J3�v������S8a�Z��C>��=h��]�n8b*4�VX���_���[�/-���:M�ѕ��z	͸�H�~��d(xSc�t8�5��egy�u�Գ�Q<gJr��bs�b���3��QR��ڄ�D	�����w��*Y�A��N��q��o�4div���@�2zT;���gY)�\,x�b�)5�b�d�u�����Zr��g_p$����2�[í?�>dA>����H�	���5�~2�U��j�nӝ���uc�k���qqW��~�M���;U���%e�\uU\�������,�(����Q�mJ)�W���<�C#ۡ����Bf�Ĥ���.H1ܑ��vv�͖>�3�q��x���Q�MúX[@X�p7�I�k�g'-��+.w���7N�-�@؄"�.�\uG���Ma��[��n裋�@�5n*�,�}%����w�a�+w>Ԏ�$���8���, �-�8��s����ߚ�K��a\/�pهΦ���C�#͡�ȓ�M, ����u7�>���@��"���Yqz�z�bW��"�����	vu� x�?^0Q����D���i��HB��;mK3/zAy�\8c��L�9��5��s����N<�IϏ�vw^������������.3�aOG,�X	�Mu�\��gP<X�emn�L��)ߗY�~,Y�[������5IM4�l���1�HH}3k]��1]�bd����B7p��ׂ
N�4ô�;��R�ݟQR���z�{�E��1�Jͦ�iKF�CJ�����a|e&K��p?�+�b)-�(Y�w���5C2Eqb"�ܠ�aR�ox�
({������W�]�|/jQ�T>��/���a<�R ��e�7��>o�U�"ȓ�����W���x(3��M��5 ���r�.�F�
������.���v0�0�D����x�vSF��"��'DC��3Fw����3E"ao�5��NZC7�����Q���n�` i�񸨷��]K����xpd�r��1�s\�c���9��2w��d����K����}ʏ�����mE��*}���[��+#��m�������s[���G����w�}�j a0Z�eWM�( P���."�5G�_�Z�HqObJ���<��
�wD��؟:y���tˋ�c�F�w�]��0�|ͦV~]��ĉ��ʨ-��p�:�����/���$�Df�������`�����L�sȀ!c������2zKXM��k|I���v�v��������WH��]�S��+�����vl�îpx(K�:u{��U���{a)�P�B��l1�p�rnxxh##��Y�qW|���F���̗y��F�ޔ�\+��JD�d���r֥pBH���r�����ŕ�z�D���w�dD٢ܴB�L3��
�Û^ә�y��H#�D��f����r�I�@���~�۴[<&�}.,b)=؃}�$+^�F�G�@�bOY;}��eѰY;�9Г1od�p�BC��R����29��u<�ߴ <���1l�pT����X�a-�%p��޵�3�b)9He�/8g�4�;F�f�/hS��z�Q%Im/��^�����z�<Z���7���z�ι!ͪ8�^\���1"-��b`��k�F��q7�m�`]:���>t����Y�/������1�\�&�/�����ڢĉC��)�[\�c Hqs Q��K���d ���
F�4�bߙ�5Ѫ�?AeSD��|5{��KF%}��F�JBr���a>uW���&Zd�X�c޼�ý����4�17��fC�몤Ü8�<ו��h_��#��/Q��1���� 5��l�R�{��'N5+�� ����!����U �fb]�R����Ţ�Ce�ax�w��/ ' p��G��8�z�]]4f�>93�\�C�:�O��s��Gyn��@�.�.��S��'�ɦ�'�����g���d릨�Vu�#��gm)�1�L�/">�wV��tp� ��=Bӗ6xo0��O�7
�z:� ��>�o�g�Yy
u��t#����0�R3��,��v����G?,�z��EEPx���eJ�B���Ė�z��%̖�<�%f��ZER�cYRϥ
��6!��=�z_we�5�Ǣ^L5xV0���:������:��ʯ~şK�jKF�!�u(:�K��F�� ]u�z��2���09���[���Ԝ��3{�
$+�ZkStR)��l��DW�v�44��9<,by�����J���7�ٯ���f�Y���k��"bTR`���đ�x[�m�+�������3�:^�)�a����3�9�a
�i�U�}��ZϨe�v�8�	��	H�.eM���t��4������kJW����-t����?{=y&E��a�^�%����ہcq^��:�qm�� r�I$��|{�����N3�9J�^��q�ӭI�ӈz"u�[�7�`2{{/Қ�F�ϩ�q��4�å@1D���g ~�8��� �E����MD��$�����
,��Z_y�"�<��-]�v�gz6?�n>:y��P�P��=Q��&L^�y�bS�A51��D1���O�����B��%a�]����TJ㯢�5+���]-�cy)�(�q��~���E�|�g�a��e4S
�- hs^�Zl�fy�E".d��[��%���޵�[
�������c�]~�\[	�ij��?қ���c��'^��ʉh3�	�N�%��ƂĪ������d��]SC�`'�N}�E��R`T$؆(�ܨ�q�&.�1��@�bݹI��50P�u�S��= �*T&�f�U����$ç�6Z��5��p��<�X��R�D�wf�����>r1�6��xS�;5&)
��;�ד�v����1H��,As��=
�(ڢ�ՆH΅b�Y8�C����	Di�h���D"�0*W�	[��L:�}�w9�A"]��9�$�6�fv�:�iXj�Un�]�;n1���ϜѪ�ϴ��)d_�Y� !���"��(���ʿ�	L��B���Z,�q��`e�l�C%�GƔ�+��M¿��#�籎{���f��u�v�����s��QT��ۍ`��S�$�y��HY��Ot��/$�=8�uc���~aK��j�*�K��W�K���NC���������%Jׅ|�f��뮢˘��p� �{�ʔY���q�?� 6v2���@Ӭ��e؈�m��3���	N�Ո$,*n���M�?�rr*�cl��#8lwn��H���{x�ibg�!�u\x�@Go����E�E�
�F�Y��9�8+O�O"\�e�U�$���d1�5wF�<`U���9���<�v�b��|��T~w��ģ�WJ���y��a����ݶ"$���#��