��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��)Y� �1�c�{�C�9	��܈Y!����lJF/C$d,�V�<�.
Ւ�-!S�h��n����X��ѢS�R#`�ǗG�ݠE^�^HQ�JDbs��:��y��I����@�1��'�1�Б�4۔�K�s�~�Y.3�L���G��6���<\�.�
�m�܇��Q�o�j�>�o���L0��8_����M5ZN阮(貹��.+z�9�Y�]}"t�(&{?���s3�!�ii�ߎ�u�+��S�,�mI�=G�/I� -�Ez���xp�󴽏�i7s�[��9���?�i���m:eT�!��W�T�Ì%P�Y�M7?(�V��ē7�=�@	��$����ֽD�(S٤�����|>
LmC�r}��?]c���r%����D=�����h֎�	)C��k���ˑ�;�,E8��5�'��竣sC������O�X�Ur���M ������{����_|�"S	M���	wH =S�#h_��c(t4�g�d�Ӛ����N���w��l�o>ʏ���cN<�B^��҈^���ls@Qݓ�lP�א�^�:5��^�>� :�rY�-��*�&3G���*䏷HA%�3CU(�"�繖�
�?K0�}D�i�7o��j�+�j<1१~7.�r��$�|�g�Q(b���u
84�d�	iF���S,m�VjIU%p���X�����V�+�R-�XUW�����(��݌�:j�gO�;�HQ��ƈ��d��m���ʡ��O�m�n��y�$�@�{�~�/(Ƥ�뇲��\ݚ�Afۆ��G���'~���bx�[�/�I���Ʃ����>�q��{@H��6T'�S&���ϋ�A�x������r��X�ȓ:D�!���AZ����ܾ�0�B�ܫ�#�(�>��ݒ��^��9���RF��^�W��|��س�Nh���ñC�P֙�񛑜::sa9�YUu�g�B�ܒ�w{�']3?ZM�Jfz&�HS �@�aß�<%����1�;8V�[���ݴ��N�:X�z�4H��^2+ȉ :����+;ʟ��u�� ,���	�T!z*�ľ?B�]ꐾ�B�Ԙ��H�� ��Q�`��m�y+7/���WYS��&<-�"�lE�U����<0}[�-��E�R�A�&�Ϭ����,�(�7�ַ#p�3
����z�mo�֢&�Z\v��sJ.$@��u��]}���e��K˭��|�������|Eō�Ē���r��Ѳ3����f�����x`Vc{��SH�,;�ؾW��a��idm��@R�M_ј{�%O`�ڞ�-<)�	��zb�V�i��;+�����D.�G]�~���_�|��Ƭ�%�wϤ�)A�_E7@��4%���wY��2~��)�j£/���e�{]u[�����I�j-�afS�������1[�£��ȴy_ûb�1�9l���z6Ӷ�[��%� n�3I��SU1��NHߪb���k����B�7r�4uA�۶X����J�h�Y����5�0�7�8�p�
�2įW�� ;=̯��G/���^+�v>VǙp���X���j�=x�7(��^vG�B֜.��t��5#P	���W`&��_F:��M�����u[-3qn�9�LB3~Z0ܙ�V}S*�?�#�Eg��ZF닇bw��)��|\iuo#��ÓE��\G��[����u�c�%˹��d�?�(%��Ӭ/���^'�|ݢ>����-z���K~0,~���0�X�&�u�W�|�`K��4���uهS�ky����3Rě�6Lʲ��DL=)`	����;e�~�Ό)_�3+\^+0�����0声(���/Q'!Z�-ý$F5��dЈ}�jDZ��&5}����+�s���|�������yAȰB
q]ju1j8,��`��?�{�Q�u`��=��>�������?L��R�p�ȷ˨�|��Z_E[~�r'a��n{x�Q�\�/����)(e�H��Ln�95V�};mߩ�-2��@ ��y^�GS�ά�>sL��e����� �%�E�Xy,(%}�)G�Qc��)�Wxn�����i��te�^Ϡcp�w7P����1А wӁ�HQ������I3��
W�RN
%����E��f�|\�Zzh�����{Ο}3�%�"^�*�YS��?/_E��-G���|�� 0Yna����Q�e��@��<�=U�>�:���'f�f���ݤՀ�U4���XFmz%J�Fiy7��Y&�s�}X�L?�9� ��#o���K� 3��ܟ3��G]fk}�?ű�
4��$2�{���ޏs��zQ��՞�-����̿�V�Tv{��J�=�R�5"��9wx��(N�n�:V`*��}����w�Q�����K�;�d\���dU9щ%тm��y�%�ٰt/#-���m��J'��4l��L<��� �+E�(a���*l���9��?$_J=�1�Ȟ>��X	��鬙�d�[�'���:@�;���rO�4� 8#�oCvi���$�Mҙ5hD5�ݴ4�ވjt)�<�̀n�n��
�]�ߒi��$��샌��L�g4��;���{�B-_��D����=��[��$�L�O�J[���OKpx1�@9� ;c����o�%�>74#"�MOE����h%������O$Uz�˩=�p�>��Cׅ Ĝ��b�=�L��*������QzT��0%?�}tlE!�~﮴Mfws���9$��lqJ<7�^%<rz&'�,K"��6�S���&�!jf
�������d7�+������ԕ\��=c�3���V�������bnק�[I������Ny�sƟ}�'��u�GAG6�	J�4i?�?��14�\.��:}���V�q�2�a�"ߚ+đ���^���J & �B�u�Ȃ�޴y���-���(��`I�X�{������%W��M��B�N\��Sn���������\}���ɿb:���-VDe;n(5���'M��Š�ڸ�[���Bl>>��9]4=�Y�V���<����]B\U:Z��>i��ׇ�x�h��T�4��U-�K�Y��I̊��r��P��^�h*�ߺ�-�mO���EGe�o�y(ڞ���GG%V`��L��b>&�R�d�C��k��K 1�u+��8-H�2��Pr����f�L���?�ܽ|�a�+=�F\�x��'Ň�������X0W�VEU�B�ev���s�'CT��3&�ͻ
�S0��9�����ؖ�k�� ��c�߹Q��R��xN��sZ����m�ֵ,�V�1\[��"R�׻T��Z+4n|��H��]�
�2���~��v��ف�m_8#�A�'�i�F�����D�Q[�L����E������9���<�K�E&L��n0�ր�M���(u��p�R5b���yF�[`�������5�yo'�{��ٸ�<�a���$�Wi���S#;xL6�X,�p����A��;��0�2�@=�m����W��;���0�m�#E~"�DQѯ˄��z�Pyݾc����&�;�@�p&���y�`-�~^z�V@`����,����|d��)~���UW�		���U\����{He�&T�`������P��U�����[)k��:߂�E�g-�G�[m|$H��n����uS�Pr@�	���!��c��"	�<XK�]�~�&�ٻ�̞������-��K���,��yC��4٧-ͦ����#'މ5���(��p���^߾-��X�8���YY\�zo��q�@8�W�=ìE���a�{����Z�%��8���P�5��1����C_�?�<�t&�Oi&n������sї���y1aҗ�li_��Ѫ���}��v�LS�p�pd�����xq���8iÃiu_t4 (��M2Uy�!W%��g��1���fj:*�O��gh�s�U�@���X����f�	5��ƕ�;�I-��I'�Nl���]��B;�]ޢ���z+<
���b>�-��a�I�C5)���J�G�=���Q"��ԏ�}O�bA�����0��^[�@���OA:�4x5��ʁ��>,�I�
�ȹ#u@W��w�$'��{����u��Lsd�S�a��Y�Cv�[Lo\O��V��/���rμ^�}�d3R7�U�L~��A��U�٥�:s3�"ez��xܧ��4�+����"x���a��S-���VRn������AN:��H�!P��cm�y��@�w�af�l�:z0o	�L�ߥ;vke�i�hdXxL�BCω���J��̔��1+'c�U�a���Z"���`B@T������)�|�8S/>��ʫX?����5�����obX�t�U��P5c�5u��6����#�ɮ�|��Ç�Sh`L��1�
�w��*� �9��ݔ�5hԲ6�x�_�@�v�Ƒ~���i���X;ىUL�n�����B�!9�3璏3������"a�3�U����V�UZ����Z;Ж�Y!�Ƞ����u&��\0��`��OE3�k2P�78*]��l�p����ڌ$��F�2��@��B�t���о ܻ�'OC�)O�NS��ʢ���,^֒%/S�3EZc�qO���;�ˎeE�B1XR��7Wg��� ��9Wb�<-ao$�)��< ug�{+{{���31cP�����H�bŞ��o2�،�X�ZuS��#CBFaR�uC~���62H��޹Ъ���q�]�dE9���b�:ʑ����Tp�js�o�װ��*:&��3_S]dUQ�<��ˏCs]�H�'������h<�����.��t6��t)���qF��-�nJPn��{QvF�9����6�ђi�Fh��i]d�����Ggզ^�W�䴔K�/.Q#�-S�l��-�E�U���N�t��pj�i:\��E��8e 3���Dq~T�~��¥�`�0��.�2�ɪ�/�۩��1�bu��I� �|d�;�!�E��c����Q��x�F ��*ae�6�A����0�aϱljw&dQ�C�2x�1����az�y���)u.���دT����fp�H��v�0j���`�+@s���݄�C*�N>m�� ��u�~b�F5:��T���#	Hd����7|s֌�| �w韓o�.V�d�V\��Zh��`f�sn=U�:�,%q����oX�3ߊ��,��$�M`�X�;"Kw��'H��r�!�.;}�'��L�;�C�M 뚹_�x#��]��Ћ95�ݩ7�o�m=��{=�O����Љ�z�糡�����\E��,��vޏx��&Q>��+րcx?"���U�V�~�
v��"�Ϥi� .�3;���e�4*��^w���r�QU�߻���N^\�?����k�Nmt��5[������+��-���#�!���f��.�*c�ɜ�Y�w ���3*�0گ��H�9 ;ݶ��ĵ��b ��5�oQ������3"h�KUMc���Uj �_���ۀ�HsX�����T��c*_W��eH�+jh���8���C�E�60�9�Y�<?;�lH��#k��U�w�T����!Z�1	֕M^��$I�>������%9{��,}�S�;S˃���]k.�IӢ��<`Ȅ+u�67���}�g���Pv��`�����v�#� �����)j=Z$ .��>Τ�_6�H�`��8(��R�T��<�';�`KX��_�k���1�.��RU~��ו|��IQ(�����a��;}48�d�󵼛�d3���;�;}�`7�ѢuV���aH��Vޚ2���\66�$3�|2-t��R?�S�yD,���9]��'�"ͩ��0uab�&���:�'s���~��ly�A�L7i�U�������28>�Ϋy������F̅ޭ�����y�ynwԏ��.M�':Y����^�s]�X1����������ؾ��_��]E)� �pE�n�����<���}@:��>�G�.cDB�[c0��D���CE��)�ο ��� �P��Z���	����T���^�I�gt�C�Oy�H���WJ&0U����I���D{�VKL�����M!�[cR�AȤ_Ɨ�����*�=��b�/�}�&F% .GU7��'Yl�f�f[��@1Gb-�zfKG���T �QKt�5� �8mYL�'����ۤ��&�t,(]-jmg��2�JqT]s��-�c4�d���U��寔��'	y��s`x�����s`ø�l!�P�Bd�lɓ��T���d$Z�u�/�o((c������4����3)݃G,_*��6���T��vI�a? ��H���+�t���ۢ�-N���1tXb���R�2rP��Y���B�O���1�6BT�.	d1Z��&�zc{���e�([�a�p��ac�p�ډ��abn-�ݳ��\R�M?��gO$y���1�mR޶�ui�Ĩh�X����jG6SO(r���A�U�/�[Sbe1���}����J��Pv�����9�=�ꋤP�� LpS����?K�-c�%2����?�hjް~��
�A�p#�l�B�������JS�)4]�7�a+��3����VtIJ�]�ڰ�:M�K?��AY|� ���Mà���Tr�?s��Vn�U�|[��!C��'U��<B;Htz����'����+�����x#�ß���� �̝��wO����zf5�Y=�8Qų{mR��m`��Ơ\����3�ѱ�LZB���"�۱Lm
�?9�fAm�w�#�W6�f��ХW��h�%�2:J8�6������%OB�� ]l�EG������j_j��C� ����b[���W	
<�^7@�d�۞F���K�}U��@�LHW��9P����{Ƽշ�GzJ��>i6>�[dP��}��H�Ѥx�=�=�IU:d��m�_��^����+L�^Kv��3���CGX��t&�w�L�$i��g�%pҪ�+&]�J��[���?:8e1H��:�"Ġ�|���al�?Q�(\}��u���I�A�4���XX+��U/�і���������$��1lO+y&R�s���������d�����=��)�`��]�*��T��E��	{���>��jG-�g�8���EH�Ț�nk.-��ae���꘏>XiZ�|�^���C�#D������
X?%@/i�M|񀘺���.���Xpo�.ú�0�:�6�h�oϢ�.Hſ|��ەpA9��W
���	�wɰ�I	�:�5OT��a]fsZj-�$��e���A=l�F���m�����E����[��!�*�GG��XF���ӣ������^���YH^����Y����Y��]���ܲMW�j�%F�g+����=Ju��QG��9ɝ8���L�L���Y�	͹$��)�U�D��2%��&�tAdqC����}Vl����\�#��&&@�؇�j�R�]�s��Ť#7��稙X�&PN+�+ᬲ5]-ͧ�xO<Oz,Rā�ɬL�w���
ȌR����(��T4yɈ�M�D���O
���@���P
�E���3��:���H��gq��3���q!�9#�=+l�W�ȺI���#4I�׷B�[���,�cQh;���%�^MYSEg�����h��=�cK,6�
v��Ɩ6�>2��c�S�]�z���Q_�MM��~cV���X�����G�wER2/yi�����	���G~!��xώ�t��IB�ʎ��h����>���+�q]N��L�͌�c\J��"a��E�ƙ�VH�Ki*��O�X.������,�Q��ê�m�ɛ�p�M���0�\��z��������O*O��nʂ���d.!��q�^m�]�J��ҫ�M��؜��_B���p�>e��˗B��"Fm_��)���P�䬎��c��(����Ts(�HQ�[Y���)��aE lO��c"�`��ܶ��,�C��t/�1d3ӑ�{�Tc�~�wƚD��ͨ(��Z�f�J��h'�(�Oəzz�
�Ӄ�ݴ����j�8���>`B��G��Ba�w�7ߗ�����ΠKA#6�� ��s_�K�?CY��/@�hG����Ω���� �rݲ�'�9��%ȿ�9�uβ��%f->K��,���`���]�C�����ֳ��A.}�D�Hr?2p����F6@Oxi���SDis{'���K%B&��A@�"�0*`��[����ߩe��e���&j{<W*�['�