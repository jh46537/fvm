��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��e��8_����+K>�XԬ=!Wl����̊+��:̑^|;\,�#$l�b���)�OP��W�&+brgS��gt���&C�_�I}ty��;#6������8��(�α��O��$R.�6��L�|�	s�fCg��3�T���Jq�Ҏ*����wa�A<�"�&7U��Z@LƖYu�u�HS h������aI��D���Id�����{�1�����!у�t�M.@đi�l���i��	�S��_-�|ICu��q p��/|�0H�S��T�ˇ���|?=,	)t���T������T6q���#G%?��9�""�D f \y��6o��X��>��k��J�^���O`#\a��#V�%/P܍g0t�=gB�(i�U����� L)8�����E�dZv���4h�*���]]m�X�������?n�c$N�5M�8����ou�N�#�&D3�*�]�x8�4��i�B��	���z�东\4]��G�d5\L馨���4 }"J�3^��2�`��� �|��ZnV�WO�p��	�3����Tj�k�auYw�8���ŚV4�g�SM��A���bՁ%-Ֆ�~�U���:��D��ؠ�[��׏vċu\�~6C�����W	XS�,��/T�%������fG(C(���.Ծl3-�l�8g=�/h���~��� S�8�/�K�z1r�g�	,���.;q���/Z�ٶ1Y6F�l*j?&���%$[I+�A�z���Nj
�좡����}v�7�k��NѦ�ڒ�v�FF+bQ��u��M��p�n����ufz6������^"�����>	�p'�A���y�'�S}�ה���<�������D(t�Q�GMCM���do��|X��$ �$��U���/f�Z��f���Ȝ�P���P9��F|�0��1u�$�m�ybk�&�O�O(2�K�H�=������'=�����1t�nY7�c><���vi>�>�4`�>h�'��ƷA�:eČU6J��ݹ�h�`�<b ��|��)�b�+�NE���f��z�C7���0v#�uc�Z"�
|�S�3�BQ�����m��3bM�/����� |�6x��|7� ��X�*D%~��H]��Τ8>���2��dCR_�KN
�����߻ve}���U����O�$"�Ō�"�qKc�V��'�E�i�Z�C`^S�gj9;�}^�
�Ұ�g�ˉe>M��:��)>Jr~0db�M���T2��	!��~�.����s�I᠅N�v$9���KD�����0h���,�E�YЪ������~A�"9���Q��˜�؏�>M;�0n�������B�ۡ
O��c�X�@��Pٜ c�:�;�] ��QW#���>�3N��������ێ
&�5�F�r���	K�#��w5��,��Fv���ޏ��~����h��n�g5�+�*���ȩ+�[ϯ;��EH*@q�lEȃO��3�ި��i���fWE<�\��:vQ�]ʣc������m�3�ճ2�{����``�LLf����°Iz�L�|﯑��VP�Ow1E��X��7`m�j�%U_j{�r1����>!Ha�ۈn�'x����z���NY�|I,�|!G�>�4g�|`��v �� ��l$��ao K�_�R=�`]�?xn
�sHѲm�e%_�Q���e�'-�h)����]���@C�`Q�8�+�i��Ż�&r_V7��7��u<��l8g`t�ue4��uK�$Fx�Ct�,[gؤ�v�!
x���%�tx4�����K�.*�uQ�9�5��$]���m�aQ���!�4�J>,~Ҁ��݀�B%R�;�jg��E�2��j!Ͳ'U�C�ʆ���
��f�5���"WӐfz;��w��֘��͟؉E��ȐE�.��a�R!�oX���Q)%=���t
{؋�� <������J���!�-��"�DUQHD_V��O��A�m |�K�hwg<��ws*�EmQa9^���~-jd��cK/ƨ�����8r�k�v��i�	�D}�2\O$M�ͦ"`ŏ��̌�a��z��F}��U�'iد�����>���ڄ��2W���1�f�Hh�=�#�z��)����H�oТEjr�=l/�l��M��WD��K8���i�� ��?�j�6Oi�8;�>�T4�U[��|��U�6�:��*�u�UD�����"W0!���JX%�T���Cܗ	��L3���fȗ���jr��;W�M�p�I���������a�%���q�3��[�JEr6G(���h��JQ��v�d|B"����"FN�%���q�2��҃�9�*�,�O�^�<W�&�5�U��0��+��Ud)� �ă������J��^V����5�K��ǉ� ,� ��'��q�Χݩ�s���S��:_J�x�g*��#o]F�>�nɪ�r���c��9���U�ԓ���@�	�*����+���Va̎�l&*޺���{�ߴ%��,���s���xf@������2%=�������x��Ԋ5�л|���lD�s���OQ�8���kUG1K��+W*�}�	֠@sћ�a�؁?���RB����R	��ˆ���$<��ǥ�((3�^���c� ����{t�z2��8j�:����@�V�r3�9�u��nլ(6��1ճ+篅>�܊�|-$��纯Y�����h��
a+�+�~!Iq���/k׮g���;8�@w��f�@��D$	7����<�.����Hn��ې�0*���F4H�.k�ѩƅ#��*"-!49Ha&�����H��kD���)5H��fKr���Gz�q�j���+�U��@$�'�͛�i�Z��޼^���q���j��#e5T�����m�w�i�P�<	��.3��W`��kb�߀P��C���I���״$s~}8��|��?D��sX�T<���]����Uçn�i$B��~J����H��Vx�ضna�Y/��	��4�����I0�LYS�E����������O+*�YUy ���y1�S*��H�q[��8�HSU�l�%�X����@��da��/b���L�t@ ��Lu��)�+ �c��ȸ�����6�CW��o��V����tRӆ���8�"�$�+yi�܅S��֭�E�?P%s�=F�O5�Vv6'�xV.,���ay���}�m�y� �@���noҞk�ɨ�b�!���hE��Z��P����0?g���(=�d��o��?���xܵ'����	��,��B��Nf�l�+���["yJh]8��2�XU��GH��K��c�<k���Ħ���'!������(����iV��5�px(ڛ-b��:���)P�T������K�O����B���=����Śb���fX��'7�ӳ�{lI5����P�� ��?�%�j_ల�!6��~� ��uo�suo½���H��{��8K�ZH���$��r1�}��}4?�k���r"�'���*����m�K��?(�w���d��)_��F����w���� �$ER���/���3�����w�Tm���N��꽷��/je�Fxcgl�ֳR��H�J��@��iC��l#�Q?�M���-}(���g�������3?-�?˧��0?̉�d�ե��Uw~0��	D���2b"�67f�7+PF�{^��+�3ቔ����a�ߦ��y�}j�z��-B[r�^İ��\]g��χs �9TJ{�:�*�t�#�^Z�G	m��pt1�֣~*�&������MXšvy�`�CZ�аo>�إ�r]�Bu �4AmT܄�Ƙ�d���<���(d�*�r"j�Iiw���D�j`sɜ�m�y�7�QK��ouJ��u��(o�Y�G�Ͼ�5��i�g+�̿kg��Z����8 q��x_��;8`�ұ�P���3���J/^���ho��{�C]��ﬨ��>B��c�O�m�%�'���f�r@ e�@b`������`�\dZ����掠0Sᘤ�g�(\R9\"�>LɇS��ƈ`f7����g��u�Ȓ�v
���yKF���B���L���
�Y��g��J��'p#�j3��~�����P��>��7�� �L���,j��@�fg֭��� �"H�˰ޗ����H��皽,���蚲E�umV�(@V�{�m���^�]��`�T�7� {�Q��4~�<�J=2�p{��:�*&z$�8{�ks��(D����������h=��jM�м�/�FBP�Brkˎ��IGy�@��JX�ZS��t+H���:{�Y�-
D��~=|��=�q�/n��c^CL<���M�n�E�A�7]H���9�_�04:��k6�n���YZ�͉��}5���Qn[�B
9F��sv�=���^��
׊peV�)������ir>Fv�$͎�b�Z���V�˳��֎�a��d�"��a�r��9_��	�'����rq�4d��:���h.�Y��YA`b� ���l���Ҝ��h�v
g�F��	Y�4�i�����α��F[��!Ǘ?J� ��0v�?LG�u�O+&��>����ϧR�T�Z3~T]��I��N��%(t[��P?Q����2�^�4$s-�2�7t����f�1-G���'�B��"�
s`>�?�O�n�
�RJ�G��8R���!gj��TP2{m�n�i����Y���%v;�2jh�A�Q�|Sl7?�؎G��H��~����U3��)�ag��-��`�Aܔ��\vL lm��sLoE6ڶM�m���,��)a�	��� �2,�,XH�F3HkgR�e��Fl�Uh�X�f�"՚�� ���!�}���=�S�l��C��*�����u#Ю����iR���Ѳ1o�P>�ԢCi·�$��C��փ���}��]3k~	����*����7�d�^�U����ۄ��@z���Șx�-�)#ƍQ���O�51��F�*��eYP���򣾛��|�sBy�A�j�y��{l�ݑ�؛հʥ�Y.�!��?�e1�jԙ�5�2� �"V�~��3`�a���X������f�砓4,]��02���"�M�kI�H�����w�c	e�<�{"�hv�i@�.QR��ҎP��$p3�������)|���&�Q�P�����(�}{��{�NI����6�Gv�/4��-)]�?y�C�A�M�+�m��S����}�B���t��2J�~��[n}�?����y���#����=!7��}1��䗤6���<l�%y|���%:��v38+���g��5j���HoI˖ֺ���v=>�?��e:�}s�:K��>���.�nv�Ȧ�5�Zql�|/�{�棗�����S���Z���<OMY����	e��6ʕ-��_�m�n)ˎ��:�S�F��9�Z<j0�ʸK�&'�B	8����m8)�hP4�ZB/�h/�0�
B^2��~֑��e�����<��L�'@��@ɶ�H�����t��xK����,�_�<w:}:�2�d�$���2`�1'f��i%:՚fJ옔��P��/�[2i�$	��+s=~H�S+��"���>5��+�#s�.�eunG��~ؖ�i�J��.��?8�V�pdG�����<�VJ�E�ѧ0#��6�����3�Qh��Euk��������j���;ʹrI��%��s.�^]����>4�_�.�N1l�ZڋP�eơΖ�;���2��iiE�;��#E&*#�����\/b�@蜫a�aj�sG4e�)	b˯,Y�ݦ��B��:b0�6jiF��MZ�	waP~o����lw^-�垆�{�C����s�A�0c^�Z�{��Xn񀜨�O���:�؁/���riH�L{�N�sߠC�یɚ`bS������-F⇇EWKkD���[�i7߃�^9R:�pЦ��AB$�Ƹ������`>Y$�yp�n��d�)��Ks�	_)�~.�vk��p�-.��=޴/�,�m�¤����?���=;��zj�Ͷ��_o$�\ �7���=�*ʏ��(�íM^���\�ɘq�!jFH@�A�Pc���4?�:�HT���)� ���Og�̄�%0��ͦ�8��;�<�7����ٮ}�!Jp�p�~w�q�����v#�n�D�B�L��:{�+*��t���:�j�U��", -���ᇵ,���7��)s����ݕ��g�$ΜL�%_e��@���^����|���%��
��#�@s6����k�=,�f�.�<Q�変�d	m�x��Dκ������~Ŧh0�x��o���2��x2�ǐh%�ŭ��/��r�r����§�:)j��B��Wl���K��ᄂ�0���čSB�����6����r�NVL��;��;��}Ŵd>ρ�-��7/��;�����o��y�'�����'���� H�r��pk^�t^JH�	 �br=ZO�cs�J��2����w���_1ñ\`���u�V6x��d��^�j6F�Ě��V���ӥ����0m�|&�(kD��oKǦ5��۠�!��'1/��m6�O$^� 2i�ȹ��zBL�|*�/��Z|�E�~��H�-����+�D���M�O�PMPiQ���k�X��K&�����C얦���FP�o�����SU�f�h�>��X�֬�������4�»��U�!�)5�r����7��1�KC�tH���^����Y��'� �P��;V��2ُ����$ ❃ҫ�̔�S�`/�^�0-��|�i� �6[P���9=�,�WX