��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"��Ia�W���n*���x�W��s�����+�5�C�A�;4[�CL�"Q~|Ӷp���Zj�z����zdm�y�>��@k��,�P2����C	���V�X�� �?%5�qZ��$�bڳ�&z{��*ݭ��C��6<���S�Nk�n��	�E��6g�����������$w���X�Z�n��7���K��ѓ$"F��j崦�W_�"O.��!%��1�GtE�����m�\lS^��g�ڐ�7�R�?�](elw��[�}��`
Ѷ��!xh�y�54M;�7;3�_�q��� YM؈e�(bAS��F� c]I r�NA��5-�~��̣��$)�#9��"�/S��y/�K����(�Xw�.y�;���(�7Y��,�~lRa�P�zr��ߺ����J2�ʂ5������OQ@m+������*6�#+ㄒ���7�8@�#�px�̉H*R����;>#S�x8�K2�v�[�٠xP���-7�����x�OQ�p��������8��z�P��$@]�j����t�+�lB�x*��9;ԳU�}�j��ZF0�J�B:��w5 ǀ�.�������Q7|w+������ҫ�K�u�e�-��e�D!|��?̓6����p���Q�!w�y�gU@iz[S;�x+�y��~�W^LdF����\aJ����n��qRa`&��ڶ�y�+P���zBȞ�f�8�-��5p�yW� ��O�O"������N���b�'d��]��v@�z�Ҍ:����~/E̺�҆�,;`&�,�U��O���Ы�)�AR���J Jd5��Z�4V����"���l|E+=��7-M�':/	�4D���E}��*k�|��F�?<���!5�+'~tG;1��)�?�7����X\��Jn���^�C˩�<F�E�#e�<K9"	eI���:���jX�%�6����g����Jآ�.ѩ�&k��<���K�š���W	q�b�AOʆ����F"��l���-k:�<��)/����Aso��eq6�ء��3�*�zsW~k��P� ���ǶTj�Qǰ���4Q�:�ټ�f)��G���"�Q^/�i.�W����5��(�ݯ�Ŏ9���Jq@R�gx���;a�V�䰆����@��ڪ�����`]�(�z�h�/Q���6���KiE�9
��"cn���F��
�X�3U
.���B��k����۞��V�C��	�K�aH�v6B0ʳ!_l�ۂ�+������柑`���?�h���?㗱n����CK��N���뚇@Ǫ9?_Y2���?)�>�i��üw�clE���d��y@�'���=�T�D��Ya̢D�4�/0X�)������� �I���