��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK���Z��pu~�������g@�����V�����"y�u����9�Q=d-��	��o�O��^��=����5��R��e��%�E3��?Y;��e~E%YVM'��=7��e�ޙ��w�Ov[����].�\��s�sS��F����|vB�+ŴK���+a�V�6�瓢�t�� ��e��^�0�-�Qy���p���$�CĀ�q�F���.ӊ�����"^,�ZQ�E�#]�L�Z1���9f��U<&��s��ѝ@}���r��I5�$?U��J�sH����8�������w_gK	�&���j�Ǒ���؆-���P�Y�TsN����h��̯������t�������Rf�ӗ�'������������eS$�+�����X	'�V����FSB���U��g�)4�y�֛�� )�y�=�JO���|�#}¬���료�n�;�2дjUC&w*_ӷ��*ѝavqw/4�����D"L�ay!� G�e� "m�ȃq$b�$��
��e�%h��e��NxAq|���W0q�p'�տ��2������RvPP�]	���~�)P¹_}(w] ߫�I�$��|� ��8C��0�aE+ZR]���(n�1^Z���z���&��x��o�a�l��ٽŀby<��I �p�p��������Cp)����u(�le+�k��~	�c���(d����2$������4�BWv.���R!6�u"%��#��G(�A�������7����;'*�=�]��q���~���:���o�A[(������|m�o���E8,���rӾs'�e؛��k��`�>��5���N�"��W��O0���S������IT?I��A/JF��3�?�z���}�eC��,�a��m ���%<��)�u4}�v���nb�k�s5���G*"�a�|�5M��a+���4%�iTd�/�bP[r��ߗ�8���ʆ��ϲ�����G�m<�N�T��e�3���~i��y�6;r�&��k`��2D��*Uj��\Π����]�|��0�}s�F�ؠ�j�΃Dy$�$Sh���`kz�����y7��t�������O�*����Ȥ�i5��kG_Wzi�yD���Z'z"v��M��f��k�o�E�q�������=k���'������� ��3�gqg~�N��G6��W��T
ܬ�-�K���ѹ�'κ���{�&�ĞsuMA�2�c���s��|�#�Zf��B�ӝ3_�V�Q6��=g� T!Yɩ�xxF�խkc�р��أ��x����v1��T�qByA����[S�n�V���QG��'5hz�/��jh�H�$YnO��.�p�9�1�j]5`�f=�Ck�@����W�H1^�������n��N�3�����.9sdmMN0*�s�ϡG��;�J�o��)���MC�;��B�c��:3D���C�Ə���Q�!�NE}�H���hR��n6�}>���f,0q(��(4~?�Ɵݔq&�4�pmR��I��}G���R� �K�â�K4Ī����/0��V���G�b�Q�7k���� >w}���l������$��y�1�˪a��+���5�*�+�~����V-8���	���e��@���N�|�a'G��"�]ۦG?KB��j��eg� Y����C��D�mmK�9K���?�Z�xd�S���n.�ck\�)D]�r���}.���� �1���#����������o8�o�~��O�x�:�P��Y��I$�]o�"$�E��0��Ԗҗ�ٺ��9���.<�82v������A�E�1H��	Q��W��l�k��f���pɨ�^��+�2��^ɳ�Eݛ�IU��Oq�H�|�dv,-`ƀ$��`��[K�TWb􋝣���7�o~�̐�$a�r�a[[�{�j��K�UW��+�Ү7��ZS��ᷖb�-��sP8���ż�FApz��g�%nԂSm��<A�<���*��D�@�20�z��{"<U��^�����[��x���]:C+��Մs+�1j7�1�cKA��W��:Q�����0�����9�D�;��y���|p[$��E�:��!�����Dz��;"|�x{(U� p��Q���2��G'?��`�K�!c3*�]u㔗Q o�qG�$lt�f�k�^��*c͋��ȟ�v��c��Э1D������� +��OJ�˿�e��.�`\�p�1��d& �0�!��eJ��jm��>�����zg1+FW�8�������(��ؾ��W��T����{�A6�{ MHX����վ�����
��ߘ��F����&R�D\�b��a$~3(�-��do��ƈ~������d�A���!�{,H��tE�g8��M8V�(C�v�FW6�����í��ׁI�'rM����0���o�A�� 3g��[������������Q�h�?�Sѱf~߭#������E~H�`J;R�/���=Kܯ1vX��?�(��Xbښ�%PqR
��	x�`�A�(g�?��h�@4W���\��`�p0�緿��|~���+��-y;뼕��߄A�*��8����.���b �Ȫ��xcעpl@"͈��p`s&~aT�]sk�8��,1!y}/p�!^�zcoA�2[Df,X�io[����㕑�qs�\��|��G�[�S��r��Pw,�޽�F�|F�T5Ú<�,?�˧�`�L3g��*/�[l�� ��E˱��R��$���u�p��a��v�����dIDƧ{$������2���?�[��jo諠��7�֮*�a�d\I���6L�&�τ�t{�d����s���A5�q�ٷs����j�ӐU:A�{%�r5��'QN��a=2N@�����=R�Q��5́��]Dr{C-��(��>�k2�O�o��go������������%Rj�q�����l�Ѯ����1,�z��pBm�p��Y�^�ur�W�c^?�����X��ޜb�|�MB��M�t\�^Tj0/@W8@D�DL)���{	5R��� ��Kw|'fz9>�_���ӗB�!�����M-[!����n��x�|�[�sh��O�'#=�ٰ3�(�Z_V_m�%؎��	�I�=D�x�T�H��R?�?i����{=���N�F��b`U��(�<�w-\�~����*�5ߵ��>��H�%�g�l�f+J蕟4s�ByA���ޔ���N���kc��[B�{y�u`���ּ�:v�&�)�>�S���&�T9�=�,��'�Y�D/�H���[u��rU#!Ɔ�ߐ����3m�$O@��Z����dȫ�ЪZ&,ȑ��e9�U���E G�?h�eH5ͲyQ۠�d
n�X��g�L[��-�>�N;��B"nbE����D��V����<4����F=�N�I}��`��  ��`Da�{cJ��5^�;P����"nl_��]������BS+��9��1�7���!��QN=�OU$�Ie��ƭ E�l�S7����[Ab
�jf1ߟ��(�-����'٥85A�
��(��'[�	��ф�-l*\�7|"��:#Мl͋�K�a<���a�������Y���=ʁ�F���g����wZ>^�������[
�ܖY}t�K%���MI��9k��z���[�'�WG�_���#��	kD��q,x�bљ],`�馕�Ĭ'R2�����ii���Q�*����I�C��s4�D�Ł�D��[_�Ş����$��>���t_dS7��01�ΓUt��J���������  7�m�M����1��P"N��n�}�<` �ʹc�,aP���c+e��L��s��9y������m,�D+e��Rُ��4�zd__D=�>d�9��8�0���Z8�%�o�����A�?eK�0��`�&�ۏ�J�_����X��� ����n=�0��0��%N�B�����p�QW�Cʀ��˙R���1F��ꁎ�/�ӫu�����,)kŨU����oQ��АỐ�!�r!��OM&��������a d^K�'����a�x��By+�#��VM��>ui�u��A
��u¦������_S��������ň$6�O�C�������'S=M�🄨���e$3�y.�`���4���e�����z$K�LC�&��s����ްL	c�E�<\B�;	^���R'�h2�U���c�tS��Qi���D1� �E��D���+<�������X�m�0��d*�Ci�B>
��O�'6`�i�!��?�|ƺC��}(M�z�8B_�Wy��RM�c�8!��zG�i�Cީڟq�9p�ɵdu����7�J�zvx2��7BRn|�f?�i�yX`U�b��K�[+���|:V �(����'`)h	�OWZX��M%��Y�xN�MgZ�.}Z�	��+��)�����e�_�?�41V���
`����8��F	F�f�m�{�v��X��գ����\,.����Bn��<+K%����� �C:��ٶT�W3$�5�"N�	��`��%%�������9(�~\]� .�p�˂);���8O3nb�:	�F�Թ�5�@�� �\���y�-UO��p�@�`*���;*����Pɷ@*�Ԋ��ƃP��|��QR�?�������O<�����jc2��t��=<�ԥXHɃ��m�U[���qѰ١Y[�Z	�
L4�'*��;�2LR���G�����y_�k��V$K��x��3q{�v���#<�g�=�md�[lT�<���)t����5ê���.Z�p���ysV���o͜���t����=őK�м����6F��f`����|���|�1��٤F�}$�49�TzT}��H�/��x�~���V�}o�k��4�%����?�i��E�#A�A�N�?����tA��
�V���`����m524����6�p�� �ύ��O��Ik�E���BCP̵�9CcMǊ�\;�˫����퀈F���"��rk}���r&��j�p��;Sb�0_��1n�=�>
�&-���O!>�ZG�5d����o�v��ۘI����ހr{���nz�i�`OT�R�$��4�%�
�0 |/?��/ �`�{�La^0��аeA$���c^�k���R[Žr1���"�Ŷ�
��/�Kq��d�5� �k��ߨ�<�(aH"�ّ}����\���z��P{�9%�]r~|g�M��+R��G��ό"|���: *�]g*�q�X���	�X�ɚ=�,��X�M�4�������(�^d�12�}m;n���*�z~w��5вȃ@��RbO���3F�o/���ͣ﹍�)l�艆���C>яh�z�Y�`�>l(���}E0X��K(!��s!��p���H@������{�s6_�A��xg��a~!���D��ں��sv�a�G�?Y��x�L0�4VZ -�_�14t�3�G��Yz� q��9��:Z����P�O���c3ޒ�k��힢|U�6y�*����(�UL���XKo\�ͮ�⇾<t�4|��^��O��QDm���od]x��Z[���w}sD�wگs�q|����鏌���&��:�e�(�v��.x�ٲ�T���-�����עW�$�_$��(R��š:L��V �dF���ѿ��:�v����	��_�	��VP�i8�嵧�E�n�KQ�s
�9�=�`cY1�Irvv]]���^W�X=pxi-0F}g��S�8}����,��h���0��&~�jId��Ԥoc-�`���~p�/i�f4Iz !��A�"��᫢���T�{L��H�����r�x\��O��^�c�}�@�*�* w��A�^��u�#��^��,�ګy4��lI/"q�Iqf����g���W}ȭ@Y�\y�6�u�L�(��Md���{cs�cP��.1ѭ�^��ޏ�>�>A2'>81yYVW�w��~��r��A��Tf�;�-�i�,�n�5�sg�\���>:���_�z*{��t���d�[9.��Smd#V*�%������"{̱��k[w�r�Aإ_������d%�͆�=h�vܭ�\�����9���4���/����'�?r�&��M7��x�T����o����[��iP��+��|~	�]r�P^��Vs���	���q
t��.�����H5�3é/�	���"F���t�\�������f\0�LĽTL�F[df���M�M3M8�K�=F�� �Go2�ci���J�/O�����A���H�@�S�Ɇy��g��D��k��n�b�1?���SW����[��d>�Ir�,�k�?�J��#	�ە��q��o�	���ؿ�ދ͓fA :R��!9�V=�}
G�F�~�Ŕthc��I
*�Q��}�p _��s �"<6��`�S+��o�O\+!�~fnȂvWp��=6���J�}��R\�n�� �)d�l�ċ�9�`���Z�ޢTú��=���7���ʛ��t.ץa?��Le%6��,�j��4C�w��T�F��]�dǦ�D��gfg�(�0g�bv��qhA�<l��C�גXb-�_�l����������8����Y��󢱥Ԙ�U�:Ѝ��y�:G<�~��D]�]^8�g�hSD����`��dPnX��.�Oۈ��2CnR�)������̸Q�*��ꦮڰ� �^��C����g���u�Q���vf������	��u�,V�a�*.v���o'H�ErR\����W��0�:�)q�E/�L�Q��	���<�vR��S6�Vo�cKn�!�{v�C�<�V�u��Y�Jـ
�;b��.������¦HDjj�d@�r�(�<��ݼ�ߨ���9S㏫�e>��;.uä퐯�3*��Hu�����v	�I�"cOiP��^�<�\��lI0T �W�wU���O�5�����d�%��H?,���>�2��.=,��DB\�^*7�]��ι����Wd^��\5�"�8T�N2@����T��ts�c���"�)�Ok���O#}������� ���v�w�l �F�w�[�!�PvV��o=�9$	<�k2ߕ���>����ﻀS��2�֕1� M������ޡ����2S��p}��SD�v��XJ����yp�!͸SCZ���1�S�py�� �=��C��c�N���o��� �z(���V�O�C��;�&�!�ڬ@QUs���+nD�~y ����"�a6�E��s��a��ρb�s�T�`*���!���o9��-��4E2�֘u�Fj#��Bb'�±�B(\/M}��ʔ��@��׏Le����^~*�v�d�'J͕j��Ә˭��\jX�-�{W9�p<W�H-�o�'��e������-|��2���kƞ������N��!���f���2i%:5MF�'��Ȃr��d�Qֆ	���V�ۢ*�m6Yt��h�U�k?��[a��OK� (+^n\��k���D���&�����ӽT�/;n�o��7��r�^Kf'g.��*?@h�B�G��j[���Ӓ.�U��m�5o�2e��9p�3	[&��,���w� /�=�?�cȤ�Nv�W�賦�q<?���J�M��κaf�B�L%A�l�QB�"�~g�,�v����h��#���ťP{�KWN�q��#$[~� ������Jq�K�0��E=l���$.���9����_��㙧��U�Ma�.�`��b�+���(,R�X������X�w.�ў��2S��HdP]�]�hr���vLgpmϦzU�����%��|�i|����ѫ�u-_�i�ߘ�:79��z��_��`�*�܅����[�*Y5�E�/\?��?}l�,&7���K���]��VX!h�80-H��Ђ�Y�z��5��L�ɬ���0�Nh�$���1M�w��gYPg��<��Vv�<E�M^#������na2�;�Hrf����ĺN��B�w&�8z��Q}�`,4hzr��X��<����~Oe�#�s�&}�/
��L���]��i�r�G�x�B���4i��)͹`�M_ ����Tq	\+��[e\Rm�V�`��Pc6x���#�|����`�IX.�Nl�M�m��FJ���W��`KՄ.n��-�jR�xa/�T�Z��j�������K�Z�]�ǈEh躘���zs�Յ��s�Y9�/�I�2���}���B�|Dm�[+�4�,���iC �Z�!&�-O�WD�^L��D���1�V*,E��8R�\	�GP9��[���h;��W�Q2Rp��?��`6�_��KJ�dy����ђ�����1���:��I��Oͯ�X����(�Pبr������[��{d 	� �*�b;�܆��J3��XC��d�w=R<��Т6��L�uB(/�<�$H�fm���B[r~��5�<�`��>�Ҁ]��,Ho��̼6F�n�K�R� "<D��>�h�H���~@�O}��Unp K�5I)�=�=y�}
4o
'��RL�~w�n;&��lMy�Z�x��Ϊ�p��o��ps�E����I��,�- Z�"�K;��˰F'=(��S!�,@X��ͽ�=V��
V;s���,�v܁�O9kS�B�1p뻷y^�$r����]��Ž{��w�?l�.�y08���و��:a��!�<�k�Y��o9r5��f�9�������^Li�x������g~����}3�;24v޳�4c~*W�!�Bb?�r�����D��2:&�3U�\�e�
�T\���3�Kl��,}:y���J�{LJ���y��<����)�?�h_}�d�u�uC	~P>������!�Wbpɦ�10����~:�qX�H����fꩵ� ����c�s�9�D�<��y͚1֔�u�F2��Z&���y�DZ��{ܵ/���!��e�y��Um�jFs�
c]7p�+*�CT3�m
+$��#�9�I�h���_�*�%�99�k5tY;����A����wI�r��#�&׿	WLO�ʊ�&��ie)Ld�x
-p6�Qh���Ɍ~��y'p�v�gEC�u��c ^J���]2����!��B�An�&|#��Rw�y.=�=`�\��V�Q�v��%�Gۥ�r�,9S`��v�Գf�����
���|φ@؊Z�rخ9��}����i�a�"T,�5�]L���Z����� �!o~�4�T�1�Fl`��ٱ�^ S����q)��T�B�b��T�}c/�;��O�V�E_@k~$%u	!]�WHK��o8D(��k�������r��CL�b��s�RH���BO���Ʉ��'W,7Q���v��7�Xt�k�(�,X��JE9��.,����V�F�S XNF��s!�q=� �4�vHq��4�AqSJT)�T��Ð��M>�V�P��w�U��5Vi7�V�p�;�B ̇;�:�m����)D�6"
�?y�w8�P���_�a|ǻ@�A�d>���6 �~w����Y����4��1���j�ȸ�H��l��[9LT���G�U��,�>��cw�0MDϧ9ʲ�}A�8,y@g��K��
�LY�W��EV�H�G��I�m��
�`��i���w�8TlBM�Py���b��a��^Lu�}��1���Jޅjcl�h��z�UU��Tc���e�0y<�G���C�Xm��f�ٗ��Z�^���*��X̭�R���Q�ӯy�HHo�t�:��N�|��D����u�Z��'���$�|��L�\��t���Gd�^ 5��V�y����j)��,0�r#ۢ4ZXu;�~T"}o7�r����SN�-�Um2���\!ְ�ӌ֫5�����ξ���� K4p8������WB�E8��+n��5��t�ĩ���ߧ�ȯQ���Zw���"
���=>���v��*1��I@J�^�z��[����#��H�̭&��F�Q1��fB�ps5"�o�KވC�L�x�W�
��)9L�d�Z^���:S70`*����`C��G�kO)��k�l�w3͉ba���a(��|��r�&�*<>��;:z����͜-P����F[�[�~yc#���SCK�䛩mw����DċD9;GP��S؅F7F%@�!W-�4_Lt�Q���v1�/�':j�_�4�VK��8�F�UU̻e�* Ǟ�X#T�=p0)��E�ab��.e�i�W����=3=�)4~t�fM�$H�b�3X��k2�q�q��	��ak������@�Z�=�>v^,i]��������|���Gl-������0!
K�ִfm�����gg�y���O�_q�I2�L8�~��̚,�&!�Խ�۞ߵ�?Ə���j|���!��!o50��B�~\m%ՙ52�K��D��֐����cws��\!wǍˬ{	�})r���[��q0[��Mr��p��)�d�M
:�}�����z�F��ϖ�?��:~eⵡ�X���{eg|��D+X%��h4�0KDO���S���Pw.(�Bs[�5 ����Z���^K��ٜZ'��b��_,�8� v|�m�)1��c�J��"�r�+[X�ѓ�c��v7`�*�jQbW��/r�K���c�k�F>���*U��Չg� ��dz�{�`h\p�ا��y��MSYl��ƿ��q�_��a�U�o�:���|��C�ݑ"X��݌8�����DT̜�C�^R��{F/~�EV��:�I����B��i6�b��뢰���\�D��r��Q��Q�YOɪ�#|BݫL�� ��������3+A�HPu��zd"X�.����A;�i< ��\�\F�afʬO9;�I�;ȿHJݝA"�'l,��Y�f��Pκp��Ȭ���Q�ȳ�����e�M�xݴ��
�<�;�L�o�)��h�����jN�qJ�m Jff	���S��<�
���A�0�N�.ό߀n��PʌX���
=?��l��j�3��8�҃+�Y"3&���̑nJ�<��p��x~��j�>�'�ᷪ���꽹�l�o�/�EGcfI����]���D
4�1��7���^�cF&�	]ھ3��҅�r[�[Ӱ��C����|��	�Gt"���-op�'`�	�҅�M��{��4�ظA,��X���ݶ�	<�]?%� �U��t�bbǿ�{�&=�ő;�j�e�n�F24�W���~E��D�x=0X�>��x�����\Q�ҳ52��,���p3BFA�x��FmX��*4~������o�M�	��P��H(�#)�8�Ő��_��|WF-1A�Up��dzv���w*����>���Vb2���P�"8'{��� !�jF��S�K�0�0ǹ-��MV̤�k���{�\5/�wJƃ.#���enx1y�x�rg|����DW�ߡ�g�Om�͍� .�F�.X	�y�<���'�ԫ�r�LYS�N���j���
ؿ.���	ǣ�
7��<�+J�
?�+oS��t�(�.���,���\�5+��C���%� ɸɓ�@��N����K<qt'Yx*�^X���k��/ڶG�v���J�[Ӹ�������T��tRs��`8��f
1g?��V�HU/Ly9=$�F�BjG�i5���v�5j8�F5��	��0{�ز|�;��m�e���	�괠z�����/*�����8}��w��t��!�*��Ds�%WV���5#sM���.mr=���5xOf窐E�$��b^>EIl���H��%m8��^H���X�B����o\d��\��1�W�% �nf�s����^�/l%�·4�h���w�C�w��E�5ڽ:��m��%ĕ-�/��2�r���Xh���|��$�� �%D(����!C#��rM��m?��#G��G��n� 9�LQ9X����{�WL;��G [�h��/�Sg��Ŝ!n�k��xti8�g_��E=��wa���@���^����|��m��&��D8�������e�|�$�GN�n�9z��zIki P���9�G���R�恐�I^1����ĬF��
3���aħl��=y������ ��=����U篅���E���.,.�]� F��XARe�a0����rQ�.֚���ײf�a��j\�R�b���Usu�@T�P~Q�� ��W���C��m�I���G�k�-Vֆȏ%����?��d|��}���� �8�z~U���N!��3xc;屒mӆ��r1�!*���f�!q�y��u��.+4Z>���xsDB���U���K`e��K╌>)#s`A�1�N��{���ɾ��N�Tm�o�G}h��� �1�Y�ݕ��cfH'd)!�p������~i��u��)r��&x<8rA�hQg��F��[+���/��:.�}��j[��,R�zk�5�䖁�n ^�n
Y�fM���=:�Xܷr�x�m���ι�/���AB�{{��i��U���� ����t�kDh%㑽���m�]4�I����~j��E�,u��Hb��蓼l.5^!����9�g˄�>��� ���XH(8aeߢ�r� &�[�&���ϬQ�#�e��A�&3嫅��rx��n�\��U&(���Su�)�v(�!M]���`�gm�6�����(�F;u:_)t������j�S�O��*#E'�9�lA���X�-n�V��=B��}�ի�+N��#�Q�j
���̈́N,�Щ<�%���	wZZ]�z�4i�%����Mމ����,�R&y_0J�n����S���
륧S�Q6UO��Ouș^����x��zG�Ok<�Yx(g�H4=��qK����45������F!�ҝ�����&���JD)����Ϟ�>H�|�#����u�@z��p���]�w]�`{f��|�@Q�H��\�v�_o�k�N~�70���?q�0s.W�/��.����B3Fr+���dIa2�|Q�ʕ����s��p�@_�5�9�L|?H��x]M�.C����<$�w�����5=���0"v��vvd:�������X�q�m����}�����-&Q��W�*�
����ۢ]�ɓ�T�zHB�&��F���;��mr]8�f���?�)H4�>��gX��/6 L���cta���-�]����7���S1�����Ӄ�]�<9pQ��jcD��=�"-���؋��;uI�����C�w��m�6��KC� �&�)+pB�����F�Խ����nT"�o���Sm�NVKs٨��(c��sK��4PZ��T�b��:	�󨯏�C�7����"���9g��p7�.P]�.�c��(�\�}՚�Q���s̎�l+A���ֽ�MTg��*����
�9�񉸛�F*[�m���� ���xO�����K;�e�S0G3��g���˃�m�k���M�W>v��E�Z�t݊
��ǫ��#Z��V.E��������6��x�*ZA~d��wHc��$�*Jtf+.����Ԭ	�����[��}�x�L���*��"��ZDV7"��6�s�̵�2�q��C(pIU���|��L�VAA@"{�>�kI�<�S{=���CO0i[����d�zH�䍲���XH��ʎc-���s��%:n�m ,L49:��x��3r�� �`ٛ�D.̭[�1�H�I Mvb���~�� ��"�"֯t��vui�����2Aܲx�vF�}�A�Ы�3��IZCT�_�l��K���T���B�Xs�E��#���=LT�ބ��ٰ��aU�a�����ĕ>y�Y��+�Y:Ȇ��n'/���;�;Rdtj���G0��ō�YġW�o8FI9-�)@�➊p����S��'ktyjl5��;6$�uv��s`54�A�c6!�AI񛏙�vU�$������O j{��Cv�{_�O�(l��:�|�ڇ��qJ�$�9#ѬU��L���۾���(٦Ҋ��ib�z*�v�&���+-!(���7�ʵ9�l��d$���h�ؓ#����$�<�d�]� ���	��E=~�[�k='+΢��~�ٳ�� ��_�)�_��}�$�V�DB����Kf}��ћ1�qN�Y�W�;r��7��Rb�}Π �k�^�@��A�)��%4,dϯXm��1
:vw!����1�Y��i�gyL�5����:�`�/7�=�t��]�/S�Vw���K06��4:mp�O-�4�t�S�a�Ec�Ax_��������4�i����ڦ���T&qWU��Vk�K��[�.�����F��Ո#���(A,�uA�5�޶��E#����T��eO���Os�2Us�j@��ڮfJ���5�����l���$��[�
�"(��o�R�Re�_��~��R�� �+r��r]�na��G�+D!�F@��&`�&P��0aw�ϗ�}k6d���'"��-�E>y��r�b��ɧA^��D��{s�Z"��2E��P'�S.0�����#x�{W��ME�I=#Ѩn��	Ayib�D���	�
*|1�L�0��&�I��i ����-O�Y���f-&A6Fɺ��ٵ��7h����ws��E����ԟ����T���iT���Ft_�B`��|��B�a�4���3��L�x<BWᢋ�M�pJ�5ٶ�ǯ�d�Z�7���\�8AU������4�w\:p*7�<no����@$D�u��gc��tDM���S����VA6��i	j��y��r�E�a4�_��'���j��q�uщOW^���s!�I�������EqU��sf&��uބ+#����nӸ�F���\�Z�g3�A��lw/������� n�6�b��"7�t�\��=׷�kp���2�^��¸R��黄����|��3T��M8.��WU��)M��dŵ��6?� ���ؚ~��r���2���Vd���exj��do�,��=Ow���b�r�쯀�*8E�����(�*E��kj���)�H���na�W��������8�	�t����4ʾ嚃sŅ��Mg�!���e
�������URӉ��_�俒�X}�wF�=$�|ʄ�Aӊ�.w�˝I�)� 8�o?�
� ����~���G5J�۽�<l0�xN��oɕt�'�5��2V}H����k����{��:��Ե��!�epcU�0�H�>�#��1��j�A�<2�aP0�d��$^
�D)�µ�+��
�l	6GNݽ�W;���r-v���鳼?G� ��gCs��S��l[�8�Z�]�E�o���έ��du;����^����N䌇Ҳ�1��1s�=]{I�xӖ�CV��oD���W<v��.��\h�_q+:��$%�����o�v	T�o;�K-Gԉ2=������s�Tm��c�_$���{�Xz��<1,�vIFX*�9�,�My��f���c�IV��Dzn<�Wә�NG��+\T�:ω
����$b�Q��t�z9�
|��| �>�2���~ �����X�*&�����z`�q�=�>i�HfZ���J��%���Ջ���� �k�ө�m:�+=��d�i���zHD�=�U�3�c��Z�G�)cH��FI#Zf�i�Νp�Ř���/b���_.��M�:��گ����g�W2i'��Z���V��mP���MV�u�cRr˼L�Ȥ�OINkD�]a�V�v��V�8��-���;❚$���Jޱ}�=�����kB�]u��.<��`�l$'�2�����,Գ��֛^;�ߕG<���b �(@DT�I!��PAjS��w����Z8��l.BH��Y��UQ�м1!���z�A�O��]XRL�D����N?�e��!�yI�S�{&�+� zK�+~~?�y�T$u��M���X�#�jG���,��-���R�O l!���N}�F�֜)������6b����CP¢������}�Q/ȳ�hne�C�U�̴H���DsMMPxdԛJ�Mh8���Dx���Q��hu���T��6�&Lv�p�dZ�\Pu���z��{|���g/���V���:".!e��L��m6��V�;����	x0i%a0\ֻ��`�����>��DM-��X�h<Aп�>נ��\���&�#R`�V¹7v��k������E�u�w � (=@?ѐN�#����R���I2$�q�r��/7r(>87�VJ�]�*t�
\tM�%lm����ޥpHQ�-�hugƶ\�B�%5[�?:͋��0{�8|�����@
�rd�d\'�@W�:��h(�������蟓\���"E��H	}��n])C�ڑ}I��B���8#Bd����Q����n�H��������&�]j��c�$����^QҜ?��I�>�b+�97D����u2x��b�����GO��MҀ�h{�E�rDf�p�����wP�4I[�D88Z�u�#�W��d(Ea�e�eV�`��D];eDs( �l�DU���*v��r��#3\�Hd�f��%��8��s.	ќ�UtŢ�u��-yV��;��t���"�@��D�?R�����o�{����������`8��%��M�����5?9�}�(�3&�^#x5錔Q�]�� �l���t��=�?D�ޝnR�1�T$"����x����i_�N+�\Kw��I�ovg�8��fj�,*ͅ�t���Ԏ�Jy�H�WUk,7T5�ITX&�1��]�u�f�Le'#�Nø��ᆱ��ս�L���y͇_jX+�߷K�f�fP�9ۑ�ʶ�I��f�D����M�����X���S8����T;����θ�I5�;A\N���z��&��_>p�F���uˈ=g�|_���|���P>Cw����(�����^lǡB��D�D]���ִǈ0�0�V�$Uz8�h�d��ºn��m�o�9ᵧ�͕��|�i��-�#�N��H�Ъ�lt!��N���K ��[��/[i�q�S���bL�4lvאΕ�kwĔ�É8����hV�kl��F�I6�ᖈn`[��U�Fl�X p�Ζ��T%F	*��������Ⱥ���"�z �e�A���>����Ȉ�ټL�r)��3_2�En���9ߖ+i�ѿ�&�m�GI0��*�-�4h��e�r�	R�Z���D�|�?��K�̮�𯉈 g���n���-#7�e��_���	򓕑��
����B��U�^����{�����f��AM����-A�|�*�d���{pi+oΔ|eB�E���\n6�Hc����7v�H)�.!�x���l�鄏z�� ��n)ϥ*��4v%}C�*�b[���喅L��5QLg��r�e��B��
wg�@10�ϳ\_��%������T�X5C�|���j�	��@�w_�[ީ��}���z�M��k�\�Mp�ګP8�v��f�M�	�9S�EpsZ]Z8�m��G�V��j��:e�Ɠ��Y(��zh:�S%�|�6��Y7s� �x��˫W/�rY�U54�A8�c{�gT�8h�\�����(��2�ح�IC�m�65�C��O�����G�喞l�R;�Q�� �P��8OC�6��OX-��*4�r q�o��a�K=zm�E�땆C��i_������I��8L�w5�]�:[~���}$89�r׶8~�MQ�
Z�4��Fk�$b�V���؆�����}vm-��m�Aӕ#��3z" �q�ra�q���C��LS�����o(�(gl?O��)�ڢ�̷}�z�d���ɗ�S���M(��*��:��m�8�e����;)�S�c:�fsj�Y,u�t^��ΰ5���6�0���Mx؇��.�X~[~TRԝa�Y��v{���ޡg�}�(����\-|t��a��]�����}0v -�(R79�b �ޜ��N�t)�`sM�͹l�
�7��w����g��dk�5���֝d�#�REN��X	�X����~�o7��5|��\��+�o�Vh�� 4jR�9���VQn�`�MW����4R�l��g�:d���9��4��*y\̢X=�	���VoZM����4���CF��7����@�q��-�V��� ca ,���.]��P�{k
���Z`�-ɂZ�����{�ըW�(��b6Gd'�@����W��)C��q�7��4���PMz�K�ӗ�b�q��9�d�~�Q��i��{of��|8O@ʣ��Gy�g8���R�?66�|zX#˃$-�M��0\��eQ}m��&3+���F���?A�̨r��B�v��+��D��->�$��g���o�/^DdZ�W�������u���+�]��NP9�)��oP�跉�ܴ@��
�=~�c{�
/�!���TN�Qm���}u�ᵾ.p$��ʅ$�����"�T!��@�ʰ��κK:���qIc��y�xS)�q�J���[Yr	�TN@ەwP1���˕��4�k���,���@M3�����L�x��g�57\���ް�0�����˞P�ޠB�V%شU��p ��@��	�.�$�!gF#�#�����F����U
}ԐnP�s]d �A�	��!��븩��'�+b��T�~��ܞ��o������4~��[�,uW�O�ws&���L�_�A�l��&��e\thYp�Jm4��f!�J��G�W~ڕ���A��+D�:����S�_R�*����[����2ޯ���l�S��ޔ�J<��>��[�Ca�t\׳�H�L;y!�j��%�b�����,���|���޵�ֻ0��~_�d�r�-�ӎ���\��cL?k(P�d�W��=�i��BQ��.q��}��n�+�K�k\1%[�Lf�bV�`��S��%͋���<}c:�w�'�]��u�Nķ���Ch��۲��}&�[�yQ�c��=���]a����-��}pPG�K�*����U���>^�)����Y.�=|�.�^|6��S��w�|��i�$pYt;a������.`9�Z�=����� �n��7���>���d)ė7X�v�
i/-��H�0Q�>09pa�]����/GI��ϣ#dF�]:�\%��ʹ���0f.G)7̣����렘<�odd�mK9��xl���,_���"%^s�Tgp��*Wx�����Y��Nt����k��\ír;ϡ#8�9V�d:wd�)b����J����Ȱ�٪g*]s�8(����H5�d��I��T?`��')h̎4�9��JJOO�?��p���M�U���g�!�$�,,�sE�V�0ZWh�V�I�~�
=)��ӆo¬/�ԓ��P�в��'���Re���:�.臭�\~�pZܞ�H2�,�����Gh�6Č���J��������[��1�f����G1o��#����Ng��#7�N�%��yxEږ������N�62�}Ѣ`����|��^�����9s$�ib�e�%�Ԥ/|lq9>g��&�F؊����p>��pM��z�@�	�{�]�G�����ϗ)7i��|V�ED���Ϯ]w ��Y�	}E��0��u�0�j:���L������0��(�Z	o��\8-���Ll?l�$�'��T�^9;E��U��2���?�����v�#L�PM��������Љ��qҊEI����5d��p�\̩��}܄�@��4�?e=�1W��4C���*�}P��"$9�����ZsⓗAA�э�aK'C��滏j�0�%���&\��1�.(X��Lsp+��R5�ZK��T=��E8�8R�5`#}h�y�M�&��'�Gt��#�����'��"^X0�o�?�������C<�Li�wß7����Q�Y�-������?��'a�<����C�!�)�:g��)�D'�C����VҒG�����C����/�1+��r���h�Z �m�F�\c�7����ڌ/�N￬��TH�ϩ��d�ߴ�m�f�m9���EU�;Mח�:?�i���ٽ�2q)��N�
��4H@H<����Ä�HT����X< ��Z�r�V2˴>c;�|��uJ�/ �Mt����ig���T�{oҥ� ��ިDW�DfU��Lѭ���mob�>h�E��9���˓Zh|�9�L�rA��O�<E�I��nt%r
��H�ߩ��h�:�E,��"JL�"�҈(�c6� [�_����.�EK����$�����͢|r�6����t�1| �b����E�̪��o�)<���?@�� �5���@=}��:v���i��C*Z»�6���y�(��oE ��~�ⱶ��u��s�#-B���\��m�*�=�ߐ�)!5�B�����{t���̝Ka��P�"7t?���+�$nX� �oW��]��
ɥ�k��ǫ��lh׺I�����bZ
@���8�S�lw��S��%��ծXRfk�9��O@�Lը���7��\w��H�6�^�c�����S���=���gLI.����d@�\$G�Yt �$&��r	+�e&��B s���~�rn�Տ���� (B��wN^�Aa��R>���$yI�K���_XN��.�
����§���*Ǫ?�r@j�	�ʜ���خG>����t� �r�wk[	n�� y� ��1O!>)j	�_$oQ3p�o���� ���E�9<�X�_ţ��3z$_��R)΋��29X-�>w}Q� �QT���Z������ǔ�8�}�&�ǥz�0O!k�u����N�tL�Y�`��oA��>�z�>�#/EM�J$�7�DJ��4m}`|�D\%c���NZ�K��y��D(�'$3��3j'�#!���1��vN3jI�Fs�u��(�?z�E�Ĵ)�q�+m���R&�9�W���q�:y�
�n4.he�>�=K���;�4i��9��4�	�PH���L�����0����=|w.���qB���\'��BY�*�ˏ�8Q�E�<�!,.E�$X|�s�>%ʀn���BU�T���(���}у��ظ���
���!�2�l��;�-]{U�&���1�:��!x�pW�3l:��E�8dV��dK��wy��j�,�e�ILL01��쏻T���F��$dď��������}a��B����ѳ�SZPߟ�E����)����V�A���^��q
9[��I���`����AJxW*����U�8Uj�x��k�PԆG�8"��v���G����ȣ�C=�LRW�ix�F&t�I]@�v$da2p�c�	]�b�ί�x�5���L��9�1�B�#�O���.���P�H��iۆ�kX�����Ӎ0�G�c��F��I85����
l��H)��{���h�����g�s	F��V]���mC�=R�`/u��)wt�]l�怙Z]%@Zj���]!\��P���v3���H�e'6$w�<��������5�a�ڂ��d7x���U̖Ka�p�|0���V�P9{a��N�bo�_q��ɻ=vp���������(�a�k}��[�I����ٺC{Nu�(��a�k���������1������DsB>���\���q;F����3>���'�����\�k�U��0h�z�)���g���l�X'�o>������[�����	�u��wl�/���K�R�����e�|����d���lB�s"�})=�[�(�<�f�_,�/�?����(��&�i?�MƷ3�Ŧ7�_���Y�+��	���Ɲ���lȢ��g]�h�{�7\��c�`A���$8�XY7l��5U����?-ݘJ{V|��9o�x�q��͘Kwo�"�_%�x��Xp�R����ٹ�N���j��\��{a�����KB����lg�F�b�E�$���X����zs����������J���jT��K������y|�7T�^eE�a:jb��x
jX��D,Z0�Oov�T@(��wp#NR��VVZmVZC�S�Z�.�+RJ�? �2f�p4��	nOK��.���p�5��9(<����#�s{R���'�>��h�̿��6_���4�T]�!�=�'z�ȯ�CRV���iLt�
��`�P��YY�f<��p
�e����?;u&�f}�,ɊǓ�Y]|���ě!=�#��5���r��m<�
�����RY���q�7���w��d�?��n��anW�X@��6;g��Y���s�0�fD`CLK�����Z�DIjk)�xI-m�j"7a�詥��Ad�-mo�{2�
:�9V	�Ά�p���![���"�v���RE)��C|����F2X������6k��^N�v
b��ӱm�Ɏ�&�*ovƤc���.����Ǐ���֯�\?$�c:��^|jg`Y��2iwd7"\,��p�c��A�c��^��JP���}�|W���X��D�z?B=%>?�m� �q(1�&7���n�S���5�9��@@ޖ�*h�C�u����O�#�e��fuvR�CH�W�,���{s,�����
FM�5.��	*�}�M�x��5K�My&���?�z��H֜�M*IV��������2d4SyQʓ�l���5�`]���وi󻓒(�������Rٙ��.�=��]ۛ�qENLg���Ih�F��A�,����^R`��!'���?ɣ4� vmY�<��%C�e�DU���<��=�t���$��/t���(�骴z�XH�~"�[\�� (ˡ֖���US�;{���*c��.5�m�~r?��rQ� 9�N�b����A&G��넸�<���Ԇ�R<��fH"͖R�N6>.�o��=%��?�Y��&��k�C�0pR�1R�W|^�ߖբ����FzE�J��t`���0���	b4,e0��f��{�\<S�C��2�k����̱��#z��N��s���4fmF�z�u0�znx��t���+r�Y�C3eEjE�2!�Ϻr�üb�b]�
�(�1ȆG���U��bI��ñ֟Q�L =��yW�-N8?o,���x��P��"Y�|����j=����B���q*hFo�tx�eh?�� �c]�r����q�8G4TV�2�{�b�o�-Hva]j)�I��1�.5 ����Q;c��Τ*�s����I���1��R0���i]^�}=���t���u�5h�B��7�&~������946h U�k�R����"�-��sn4 u�H¨_�͸�@4X�%p�L�m=b`���n�z�G-��.�q����~ʶϪ�-Gt�����3�<�_��$�;�n� sE�eW�����r�V{���c,���� �� n&KD���永J���Ep����n%{v�*�8����#"r'��D����%~��]���JemZ��Լ0�R J���Gi���HK����o����QUsh�8'��Kx�y`�Q�[�[,g�2b�m� ����"1*���npv@�3�k�MO�!��=��X��m�gK��u�}��;;S��o�O�B\��S�h!�ݹק�9Ng=N4����V,K-��;�>R��^�'�Z:2��,&P&!�:�^&]����kT����>������)�N�r������#�a����YC)���,�Nt��k�G�U�wZ�2�����RW�O�'3a_��VI_�r�m'T���t/i��/X��&qC����a7��z���Wh�6��N�;�ڃ%��sG���m�FV�xxk!r�?dD���X�8؄��t~��4R6=������;ښ~{�]m`.�!�Y<��	����:���.��[�����9��|��*�����M�Bo	��9,h����*W�?�$g|U<���c�-�d��\�3�^���S�!��;��֏)�Km�
�O=���7e��R��+�m��+����zK�"÷���
�L+��4�l����K�z�n�l����U��A����LБ§K���&g��.����k�R�i#$�X�uot+��O��(������L c��A)	�1����ZO�ir�� �sXIB��L�뢌\ (^�����9Z}8<̮��M&�Y���u�8�;kݵ���,�yD��O�Z�݇�BL���s�U�/��BڪS�sO�p�mB�xdDFO8Tc��xedz|���0�pE�s�#���?5EY����c����㜣����� �T�������bt�jm���ʶ��������_~�����R��b�N����*;s� �7lu��ID���7r쑎&Vn�l&5�N2�P9�D����V"��
��� �r��+"a���������>�bU���.e�$���w��_���3LCT�E������vT�IC�#���=pc�?2_+N߷�6��}��}:��18���Z����V���0�,Q�`�Ŵ�mĶA�A="~�@;P5 ��TO�@k)+(�ɠ�Nq�U�'7*pd�P鸀��D�I��3� �v<�ıB��u���]8/f]�n��@T)�Q/��iԔ�'j���5pq��{�R��0��� �D��5��qQ�i����������� %|��r;{�g�d�1���H@�*��(��
Z�3����L���H� �	b�P�%� \�1�Yb�1|>j�_+�KJ���%	?)���jD*��+��ڼ�<�~�~��e\��x|W�]!ۃiߊ	���j���� �sH�89AՇo�V�#A���I�]p|��\oeZ���ދ� �Os)���	Gb�l�<�PӋh���2�񈢔���
;A,��8���-��=X�o��Q�G[�}�s����|7 ����1O1�c[!��2ǳ���F�#�F��m_�6Au�=Lf�;�3��&4v���J����q;�v��%��_�Χ�{b\b!���작6Fb%˝t<�/5P_� @�ݍۣ��o��%��-�� F1.b����:�\`�DV7%dW�~	�ᬁx�=��?��s���"T�tG�X#����3�t4�"r��E8j���USG�+	��thn^$x25�T�{:��vQ�J ��mɨ�1
��z��M5�l��Je"��(���dO'
(7'$�lQZ�x���p��m*��&<�@��%4G�J��'�$&Wx$��{�B�ޙa4��I�8A�"�=ʔ�V�q&�Y:vݠ���c�y�6��W�����l>{ʬw��I�^:��z$��b�(>k��ß�53������YC�&�d90����������|1`g�I6G&��A�%�k�CP����Y�WYQK��G >:8W�g�|����O}����GӰ+�(�켲o����f5��e�13�v�7n2\l�!;�%��	zm~�̾��v\mc�
�{N��n��"����h��/[�aU5�nV�C���9.Yǁ�ǂ���0���Wx���|{�-��7*!�g��%��Ԕ���x݅��!ŕM2�%�n�9_�1��*����	8H�":���� &���u-�г��@q��m�'j�)�bl��MW��mq0�BY���;q:��f9������׿��\>�%SU9���X�� /�\ǥ���[��Z��{���=����gSg{6�%b��^5�I����:�b���+4lWjJ.�=�A�i��O�z�$V�d��7�FBj%�2�J[�w��ߤ`������_K�M-ЁC���`�Z�@'�|م�E�����;�ڥ�m�8��_��˷v2��d�!E�r�$�C�:d��|>�;B��(�����*j�[Ƭh@Õ��u��,��=�D�ɞ��ugx����vu	J��1����YޤF�~|F���#9���A90B[�"��.j�\D;S��%U�}<{�h���hB4���U���.�E/���~s<w��}��*C;p�R�|R��hGs����#���5����$S-V��N�$]��f��g8���ڂ���\��Z�Qo����O���u:-'T,o��bAPw�ҧ ,B	��f�3.BKil�p����a{���l�;��;���*������_���0�����m�MU|�tb�y��^���Nf)�^]̦:�0���'���($��B׆#�G��v�����̠ן~!;�aEݪ��=`�o�5/�li' 泛
連@��i>�jH��){�az�g k`/���N;Q�����_�-~�A!�W���r�񮝊���K'�4���rߩ�z>��� #USaP�����U#�=m�1�h��՟X�����d�T�{I��~"�Vm�\�c��V�����lT|G[%�5�����������J�'e�+	"�Yܰ�s�&�R�� ��PO���1����e�k�륀O������K(�k����'Om
��{��8O~P��9���m��G����_�6�������c����S�A<L���9�YVdx8O�>���p�MS��*�7?��n�[�la�F�c�����N�����ל�'fEWQ�5' I	F�o��}�-�^ E��>�3j8�Zi��SNA�7�Mlx�l4� e�(e��Ǌǯq�s^0�"�u|���Eb���6dV����0��� ��{��^2OD*���N��eT�5�	��	�����b��o�1-�U,Η�ѽ�yfO��ɻF% Y�� gɀ��|⥂�R�:��]�;76����g5�ے�g���6��I"��^���yz3�����-JFAIZ��WH��)�n��2�B���̯�3ȏ-c���R�C�,��}|!��o/�r����}��@�p���#��ĵ2_�N.�oX=���%3?K{�ȉ��j�e���t|-���6, �,q򗃻��ז�(�6�PEY*.�����Ub�}Q�����4օ˭�� ��kT+����R��ΖiSʸ���ћ���%y�y/S㗐<$8[��4�ucx�]py�ܰ~��Y��n�@������sf3�
)��Mxxٓ!^�P�UE��d�xԬ1n7�w���!��ۦ�i��_W�-�,�m���E��O~�-�8�7�}bT����e�}tpx�vϑz,���<�`!Q7��
���L��J�͇��fr�L}�Y
���Q�_3o�o�.>%ӯ�ԐE}�}4���(��aG��k�O�x�2 v̳O�LB��>{�Q����x�	�q$#Lh�t��z-?#�Z,�6����Q�s�J�J��FQ ��2�@�#>,�-I��V�.�0v�{�����ɿ@Y���,B7F��u�6@\���2�X8b�f����A�H�t�Y��H�օ�M �݆�;i�t�Z,}��;����jxH�Esx�S�V��$�ڨ��_���L����8�Yfc����8=H����nG�v\�
O�<�7!�x�ω�������wm7�p���a��+�X`]��t��zO/�dyoEV��5�9�WN3�fT�D&��L�����a�=�Y~��)j%�?`�U)3/�ɭ%�	���W�HGH�I���B�7����&���:�E{'!!��Je�S�o�-|;�ehSk���-��ҿ�,�-U�I�2�\x�����;�	ɫh����tr�{��� N\h�l�y��[;~Q�m���H3�q�-/�S���3�>�gr�7�u�M�����י���%VX���	0��1bKn���|h��GwZg��z�������.Ė
���|�@��2�2�D2�KŴ����^�T�26�;� ���.o0��2�hB��fT���\=�����Y�Ui�"����?����2�����ߺ��2R2Uы���B�I8I^<�!�uk�(r�6��d�>��܉�v��{�^�&�K9�!��疠�
�x���v��nI%��o<�I!��螑��Nq�GӁ�ԡٟ�ˠ^p�y} �3L~Da�""���#���Rt�Kd��^�l2�*
�F1V)�(N6ˡ��2l�R�p�,s�w�MtHT�}"I	��f(7��x��}X�U帆C�����u��\䱌�L݄H�W�E��.��X,uq��hgz�2ʥ�{s��и�#f�l�<��?} ����7`���|�W��ؚw)���h��0F���u��J��"�/G�<F�3���Z8b�S��Po �1��-�u���.��og�p����L�ZQ��4E ��6��+�����{��p۞+
4���' lz�T������Ib��R�+[RN��ֲ{��b��T'K�u\���`�w¢�L����� �n�0և�w�i/Uc�A	�J_3&�iG���"^��������a%ˮ@�K$����s{�df�l�Ꝁ�*,ǿVY���
�Ԃ�7����o����� (R=*u�'n�<���H�ʌf�<9ܴ�r0���-c�(���6��xMԋ�X+����-�rq��8�F��)�N��j^r�u�3f2�$���h{:���oT�s_m��F�ej����]��{_�B�����7**|X�fR��)�:�_�eQ����ؔ��m�O��~<���ù��'���*�H6�`udH��Bԕ�|�~'������J$V���w �,��h�!�D�<��!��zM�� r���c�*���U��qE�8�F{�<�e;c�G�?�D6|S4X#���qCLl��r�過my��?���v��X���	�˃�}�S\'�;�G7��O���T��܁�\ab\�~]�ƖO�A����,��	#V�r�K��~�1���W�܌�����'d�+{��YU ̫���K��lma�˲��)�|��~���SO���&�Q	�I&�~��q����q\�Mş����v�w��s
&vs��M5�nN��_L���"f'Mn��ƾg��+��������p���M̴�bRr�S�^7<`9�V�$B~N�xN�k[c�㪮�$���~ ��X܆[sj�ah%�:���9�B]3W�{p �|x+/9�!7p��3��?��,��:��z�*�>�F��<���=	'��Vu��,��$Ы:�^��h�q|����F���Z�����ZWmJ�:�gN1f��5j��f�����*�7�2���� ���xB����Q�a��+SS�ttK ���dȣP��ټ-5�t-�	�R��4KR+v�a��Z��M����Nhq�v��w��4�9�FJJC��Ync�&���g*�LA;N�G�v��f�}3|��濪��"�hB:?m�+l˗��R5(Iw80r_=���=$���\?����*̝Qݔ��qsU��J�'�L�`k<1tgRA�F�y�"���c����L�s�_��f�	�~^�����a�@��	��ޕ&�A#��>c��6]�S��#u���4�'\��t'�@'B����f��s.�+�^	�{gh��W3U��~������ⅰ�L ��	A´���������QN�M�9W����Xt����e`!��Ӆ�C@�BMdŹ�s໯�ԧC�H�Ĥ�3�V�-�:��ϰ%�F\�Tj�٥J�Y�`�Bz@��ww����`�a#����be|����-x��'m��%�>9_�z���i����O��ԋ��h�V�^]~(���RoUk�-FbOt�M�8�l��qj��$��۽�k�7�5���Z?b�a�น�k�������ح>��=��lB��!�lu}���:��1��󉖡lo�]߲ӼA߀.����������E�bS�~�eC�>c���Xi�EJ�l�����gi��|�,*�-�*i�Y�3�1lo.g����8
K9��w%wX�ǲ��nQ�T�q��I!��E9D+��@8C������sĥ�cU1������L ��)\�6�z(
R;'y��Zy*:<P"7��!J1Z��~1�[��M��� ��DO���g��q��A��p(���\���e�jU
�Z�]d+��i`.=a+0�yn��m���3��0��n� %b>/Ú_����M��(���rַq|wUfW�:��.^��β��M'M��+���X�P(���ί7�9\�B�X�X�T�ԓ��
u�#�yӥ���M�~HS���X�p�'���C��$���Bwe_��t���?C�)�x���6La&-m�Lc{��q姨{0w^ĩU:T-��;
���ky��Nq�Ag�JtJ���xw`E�\�8����L�,P���l&�R����|`)�e]o~¹L>hp]/8C����_%q��G*��/�YB.U���F)9Bo��SW��B*�/���@�V�A7ձ�2�cAרּ��S�'2���?����
۳��<�_�"Ja�{����G�;�$�蒔�w�t�����B�=5U��l�2��/x�ox����]t���r�dqU�˔7O$��8�M�zF�2����P�V}1i��,�NfY{�"�>��;w�#�)�Xyt"oe����o"S�"A{��בIh�ћ��h){3���.Q���R�
��Xˇ���
5��Bm3��+u�&�q#8���(%�/���j�vMؒ�|L+�w�����Ǳ�oD��u&.���1��u� }S��Џ�"a?�9����K����W����kZ(�.�L�/�9�u`��$f&�<�7<E��m�=|�+r�.a�NI�fY�i��>4d{�1Q #��#f��'�?M�Qv.�[/a-������ıta�d�T݈ �lWL��s-�E=q�23A��y[��8��FNc똝4�nKjN!]�iu��]5/�W�|���j&��GA�Y�V�,��e�Z�=E6j}=�$����&�:�C�D�����|������Q�*}��R)��p�%v-�4��k2�j-C�l��%�!�(��qC�o<�}(x����},_�sPl�'|�X�v½�&�7�ar>��ъ���h��̔r��;j�ޕ���K����u��C������4Z)���S#���9��y`Gwo��.���egtq	J��Wjd�K��%��ycX�5����`	y�.[��X�M���B9[ż��e���<	W�d��Reޙ�BEG�)q�j�u�H!s1W�G���$Z��ٷv>�rw�N�6��쇳.�E	2���Z.�gؗ��	k�>�"4��#������Q����m��E~9����9꟮t H�HUg�\Wj3%�<���JOF�aߙ� Љ���L!�����s�_��}!�P�ؿs�<L��,���Ý��,�x�St7��le�W��^7iu�����T��6].�`j<!�a�|CH�i��,��H�,����nU[[	*�:Y�M��
�Y�s �u��ɖ����G��D���~q�� �@�^� �9q~�{&y��rhpgg@���
VnU�E�4�t,��i��I Wmf�%Yw�j��m�٘�_/o�mi�4�YM�L%m�~#�>L8m�&b�j�����>K���B5�6�a��N�gx��5�^�f�Ӻ�o���|�$�5��ǳ�.�JY�#Q�T�o�ϳ���9L��$6��#ZM
�R.�״�!qAPF�)	����cW~-|CAa'E�s8}Z���2�h�f�2.�[�V��:�_#��� �O�Z��.�IJӒR�#�����=�T���6M�6�K$ìA۵8V����ʸ�?}Fo���Pk�²���#M=R��/CX��c�J�ԧ,�J��g+�z4c2ޔZTBvm��VV�'�Z �{�C�w����|q؁Y���~}ȡ��:�ђ�{0�L��G�+������z�c��Z���7�������|a��x���=��`�7ۮ�H�e�?��	$�:�����jm\�Wu�����=<<�J�n�0�K�\���\>ɪՕUGV˺Q�mW��V�JO}ז�{!w���W4�C��|D(�?�@Ob��D��B�U	Eu�Ă�@��aģ��@���m]�}����=�#�[H~����a�HK�t�:�g?�j߅��˥,��,y0�d���xI0X�D�u��������Z�tI0Y{�,W+��a��P)ߦ���T�t���Wd'w��7����_Ӗk����u��\�ʟ��l���u�����Dˬ��^T�m��\kE���3Mڇ:�"��B�zW>A }�C�G W�ՇS�u��*�ѹ�w��	���[� �Z([i�_z-@��ղJ��]��a�t��l[���+���� 7���� �(ғz��ԇ��|����!Y>�	��Y�Kꢡ$c�p�\���X=Cc�.WfX��]����p)�R�#�X�=ʢ��n�)�l�7(�D���^ߟcu�
b;�3�'�S~a�{�5�R	��uc��eg`�ʆ��a9��1��^�*0�۲�I�&����T�!,�xU9�&b��5�0��O�^�6Pp�8zq��c����U�Ň:�hD����n�f��(�t�V�fB�mHjG�܂��Z�D���AhI������93$��n�j�t�^��p�Ri�/�s�
��?,�����Rd����n����;v�0X�%$��:��W��[����?��>��`uD�U�I��0��૫"G���d�S��!xs�A����:QY���_�	2��Z�2��/�\j.2(��4�od�tM.3��I#�GX��ą�&���ڹ�A/GRe�2�(�\Ä�8��B�!w���@��T��)�Q�o_�1�|:����. ��Zp��A�#��|h�t�k.Yw���+��'f��
��-_��2��:+�Cҗ3s���Aɡ���&J���r��{�H��L��Ңh`c���YW�q�#,�%�cZ�wQ�;C���]�݌��ˢt����aʵIu�to���U= PI�=�|F��p���ﳿ�tg����S��*�- bh7rqW"RS��eq�@�Ϯ'�H�[bbv�����!Oo�Fh�`;�B���Hj
��,��s�v����n��u޻բԧmѶ�>���M�w�K	?��d�ӑ�?s�'omy��W�+�G��rg��z��������x��v���� .y�ݙg����[3��5�����@%�K�7cg�elo0g�n_���/%HmH<&5�[��s����+�>��h>ϠF��w}B1�k?Qn%���A䈋�h�!#e��X�{���<N~�P<�g��E;s���*A^��8(p��Ox-o0��YS��Xg��3߱�*^(JOi��ZM�HƋ��P�[Ֆ��Y�3��9�$��s��2�>��djP����\��$͎�A�1�H�0���2q���'�N�<���Y�.H�f��B	dq��DSy;�[�K���>T�ل���̎Kj�r  V9:��y���S�;��Ƴ�]���A�YG4sӹ�t�G���?p�v'�#�'P>�:f�D�o�'w�RG�� ΃����sPF.��v����&�әS�YI���#� �rw�g�V$���L�/� vvb,� �:�m�3�{��@�z�Nw��bC�z�hd�l9����c�l�Ur&�|�peKk��>�R��m�?1'��mH�7dM������:��ŭ)1.~��}^�#3Fi��ڊ��2�� �q�[yh���o��k��uV��+]a\��6B��t����p.��@�E�s��z$�W�˵。k��{/jM�׍�{�	���
���#�2\���F���ggrt�1�,pYf�-y�q��� �����ig��2=yHv��8h��h�+%���r�
�97�N�
�XB,O��/h)D����j�?6�Lʨ5�#�S����M��KGI4�Y��@��L\��}�U)�T����]�\ɛ�t�pT�\W��K7�c�s ��p��ZB�L}������?44>K~�؝qtE�z�ws:L�-o0� 8&G� �H�!�KQOxpɖZ��Lq�ɇ�z�F��>j#��Ih`a�+t�}��6�>8.�~Y��냒s��{���*#7n3�P]�-�zn�椶�n{�xa0��v<x����]�SgER�n)�
�Lzvi������E�y��/$>�l�
b��T�8K/����,}}�Q�� ���?z���mh�iW}{� 3�ɠbXx�n���#T��
ؚB"�T�Ij9��)�UT+��܊�cDIW�`1u�(�<u���>1<��'s�Q�����s �O�O�c�*�_�bh�J��������d�P$�Gs�����R���Q<* ���1����'#W�^�1~��Z�����<������LJ֍���CZt���#��y�ܞÐQC3d�[�ts���wv����_}v�6F����������Π�ة�q�y݂��1*�dW)�5�q�4��p���笼3~��kI��䩐kŻɳ6�g��&�}8#��>�u�Q�p�"O�M�=���n�S��Mi_nf;��u��z��{L� �l��X`$ts�2��ĺ�h�죮|`�|	�:��:1���K����4p�B�1(�&��˞����K/�e�[��r����V9 �g�C�Q���>~5��>v���PJ��D� q���N}���<��A��4`�5z/�����f�^���{��_R!Q���z,���^�y�H��+jk$��"�R/��tx;�R�<�x34�Hv��Y�|f�ۇF��Z����S���k�L�rz�ͷ�����N.�D8�.��P{qq�*\�H��K�r�f��2�N�����x�"��'�P�`P�.P�hڇzρ}8Ŏ7��BF���Vb�.7�����
�I�@��d��U�kf5�J#{��Wf�  c�!d�%&��i��á	a�]���I�HS���gz[�(�M�VJ�J���v�)�p쥆������۔�D;{�Vb��U��@J�K���3گ֢G����7�����(�橔/�jp��i{I6�){HP�eb�R��t�L��#�=�$��L��邹���?�o;�db?�?`��[e�y��7�EucbYxu��dw:Um9�Qz臹w��'�I��-���y�׈����@����ư�̩�P�xڃzс�qLl��h�0��=`�k�]�܃�(KF��}����r7V���tu���^İ��
���3��'�ޜctK����h��[���W�z߿�m��o���T��tk��G�1V����Ԟ��m�c���WD�����	�������҄Պ������W!e8���6\鸫�W��vG�'�=F˗�.?s�קh҈ę�ˁ���Π�K=Bs�V�>s_pN8��|7Ak���[a�M���3��#��M7�5f��X���g�f�;��~��#��l����4T�7�J�QjH��l�&'�X�����̨��e��> J#7�E��k��p�諈P�'!�<�TJz����麂�HV��H$�~H��ަ~�E.�bd�2��W���!�.R����g����t.�6�}F����6W���c�'�퐜��0�|Xѽi��b�NA���T�<;H��Z�o����{%�"���<�q*@`j�sͨ�Ȑ��� ]pڠ��������z���B�Х2���˅(��k@3cu�y|�z~Ӭ�=�S��7`pƎ�����N@��w���ִF	��eߤ�F�N"e�%�haA�e�`c&���ǽ��3��~���`r�s���n�`�&����R�z�Ex�>g�!���� 
��[�Ҭ�*}[���Z�"n��~�Hj&�3�1 V ��U�]�m�o��-�a�P�*�'G�Rq�ve��[�r?��|�G���x�a�V��ʇB�$�;K�jcq���[�C�w����Wf+�v7��K���K� TNU~���V�ޞiS��4��Cb�9sH�Vb�h]沑5��t���D��҇Ԯ�ޅ�ѹ�$N	׌F`N�WBW�뢊!���w览
).C�9l����tv�� Q�b[5��-�l�r�PQF��y�BL��)��c{Ct�%�0��E�ta�OP��Φ�WT���r��,�g�`h�2�Hݠ~hm�`�Q�V����9����_"m֑�h)dB��/���2TX�I���\N�C���F��E�$m~Eb\%ې���B�U.z�͔~�Z�l�&�^�TN�/��^̒����p38X#3��sw��V�쑉�\��>8NzR4��u�IZ���j���#)��j���D��@yR�
���z�̠��s��0m��� b��d��TV�������GJ���Q�%r�|CxD���R�f<��:�r���n��~_�J�;�NOf�m%���� �N�q�|C���`Z��%\<bKы+�L���n@���j��o�������-��T@3˟�Z_�����/����]�ңh�};�����pT�B�}�zT4���YG]M4	�W��� q6�F�U[*��֞��!,HB��6uc�e����z5P{�ml�4�O�3�:DjgE�+~ӭ�w|D�mR n�1�j۟���-v8�Tq����mѬ�
|Xr��R�Ԕ�L\����d�$�*�
�ʵ_���	�̴���6��j'%�|�M"M[�L���v%�A=}��Ş� -��?��2e����:ַL�����%P6�����%_�?R�6�����\;�d�np>hÝ��stHC"��߅�e�4���~�`/���U�P����YW-}#��1סsƨR`��������Tj�߲��Imy�&d�x#�� u�Em��T���+��MQ$}���>|�����@`͞9��	�M��~�&�l{x"�CM�62�;Q�TH��NL$OP�k��i?ȇ��:����p�Sɰ����7O�B	B_z��t\�)WZ��y|B��|W&v����NC�)����'�v.�P��αp�7%�}��'�+t_N|*�s��̕�#�/���V��&�X.������E�ߟ���x�Ss^+qi�=�O�{�66��nC�6�u�<B~���V�t�~g~�Ѩ����/�u{8_+e��a��I��G8�͐�瞣�1x�'�"/)��.w�J�qwVko<_�1d$½�p��*)��Z��b�(��L6�)�$�m�}��t�`�$ni��l+�(=`������&� �pLa��J��ny�dTnULώ;�=A:D����'ݞ����w�sBQDdJ�ۣ�T��1.?.2�u ��ڏnL��"�5��ZyfRdZ����]|���+��H*����;pɤ5K��K��@beX+� s��ed$cNÜ�oΣ�zY��?��8 ����c�µ�v*QH�$�~f�	��f���1%��Q���b����hPu���ȑ��m2�/\
���N���x��h�8���]�=�K�)�h܌6��δ ����:	�.�ꑪ#ؘ�u��{he�j�>ʡ��T�H��:�1�0��M՗�(L��G���U:N:1A��Ë2[���C{��D~^�b,��OǞA�K�,�h�Ԅ�]Oɥ�A>�C���gp`�5{��b*l�l��1�/`T�T7c)��2AnaŲ&��t����nt��������"h�IE������><%�$�-�e��Aɴ��ϸd20n@��Vyk���T���T����b�댑Xt:x��RtJ#aiY��ؽe�W���݅+��*	�+j�))U��$b�Q���t��Cs��qW!F�ZW6=�i�&o�䦉0��e������CH]��_�����H��~K�2�y��Otaz�``�g��߰�60-��S�f+�[�B�_VR,�GW����	:��B֢y�U����+���!��Z�4^M�{e߸�5aXM9d��Df��w�h���rOx�Y J��T�h�W�0*�9y��,�8oM$�gD�c��a��,�W78�ׅT��9�mw�"��,��Ľ��J0X�P{T�SU��b*S�w�!���H�EV��'�&�*�2-G#���mP��'	�B��u�%��/⨙z��lw��Ku�#�����7ࠣ'�/�4��(�Xq��u��K��/7&[!r�n]E8�����>��A�*f�4��c+��C�d�Y�<�G�KN�ʌg�F[B�4��+aB�v�����-M ;�+�!ч���}N۝ �oer#$�֦�q#��78���W8���˒Gr����n����ѩ$*'d>���:�:1��,���c�/������Q���������QC���^�6֨��<ĸ �n[��+����ل4��Z/0�͚��dMq�u{�`��3��oeG���}A�@V~�R/R�D��؅Z�da2��}L����jZ�+Ѩ�x8��ۛ�J��]��6�b�ց�[��4KTC�hdG芑��fT��f�(�+C	=#E��Mn�P�X(�_!0��h��	o��hs�(aQ��1�t�K�l�rJ�%óG���L*�V���é��d��P�~b x'��uGrjU�1���,��A��F�DPim��lX}�`� �N�C�W��?���9H���Bk��ғ캟[�}ë�f���V}��2��\!�*Y��}.(9�Ƣ�M��S��܊��[�G ��,T�j>���0���hEMX�pt�I� ���U�fq�����MA���S��	)R��F�z�V;0�����H�k�Fh�EO�<���q]�l�����Lx�8���H>كG�s'��2+�R/D7���>!Э�V�b�[�&��,a~�}��G����X�1h�&.���ȺAWv����$�ܛ3�VG\Ќ
2��%�e{& dƈ�鰳����+|��\�q35~g�0�VN<�|b�����=v���a��/�r�ZL�=���Y@���o�Y�b��[���?z�@��qB�h��n�.HOd���ܵtR	\���mɃ=�����=;ꃧ�0��YqʁF��+�d��#��=Cꝡ-��PJm��j�Y��]��B`w����>wu���G�$��m
��䙄	�@-r}���Y7c�o�����p�djk�8{?6l�>'�(a��h<�K�\|р��v�Ȧ��%@�w~:H�kX�#�#��Y�۱s[���
_�x�oMT�>��7CB��=1���q���쓏f�̱��l�Dc��q��H&hDz��|�BfI��t0���^�_�,]�zE���$���rcX�Q�W@R�ַ��� zu�� {��.���bf��q�F �d���.�c"�)�рP�#VEU��[��������͌�vy��(�kp߬:@4�кE�ÿ��1�!s�E|gɠ��:?��a�U��XG�֗���#���c68�0�g��x.�oK�(��	{�z������<��_`uB�q��%�fv��`��)JX}ڣrk�B}��i"e��jni�#�w��{�	m��ˈ�����m��o%	K����n�%H��^�tw�@B�A�"F�v6ҷԢd�6�_���)mQծQį���fe:(Yհ-+����zv,iiM^��������O)[5�P���[H�_z)��⍡�n�vk�(�6��'+���jhj=��F��4����U�p4f�E�-��rz)�A� �9�ԙ��S�^�TD�!��=��^;ȱ���T$GyYe/'_�WA�?\���#8Ml������F���X� �H�0ײ�Υ��r��������ӁHp���̵���ǥV|��'���4V��8��-A�d�����'��|�� 3ےU�O�x @�x���1	f�2��5V�҆���,&�\P������_~]0ا�O1��T>g���c
v{c�W��P�H��:�M]�����^����,���A�A]H��v\��7ъ�o��k�du�4~�2�(���ƶ`\ [��Z=_Jq�U�J�3����
���'��l�����Tc��K2����E!B���؇���Y|�s"�]��<7恜�9T6Ы�_���.K'��R(<�"�8�ƫ&*�d��<��BL��"լ�ɮס7f2C"�8��Snr���j 햯�y��[B��y��
�ʹ��p�;M�* �4�v2�+>y��o�%D})c���S����]����Q���E'b,ldܕ�:��셚؊��C[sܻ/>eB�OFh�x����YK���V����^bu���ݞ4Y�[:��X�U^�1Q0:�ݒߺ/���v�La䘐�u���s؃�,+ͻxmk࿤�!W�C�q~^)z��ӴGʺ�{K��'۳�
+Ҋ1��ɨ����>���q���s���<z�H�^9�en�^,\i̳�+�C|�4��������)�2���5)�� ���<Smo�n(��%d�h��z���(ۏ��B���*'1������6���-�R��-V}'yY���v�\�
�*aslAR�L��Su��c�eb8�	��u�}[��x� �M��A#�B�k�u��k]�D��g1���NH[� =����pu,���2hH��qC]������w�3-L�wUX���F�i~ ��5��#7G�e;����&Έ�����wm,d�5��_ͽd�y��jcq�y���R�)�(;�>�L�o�Ɗ�O�{���包�m3���(�k,�	��o���D�Hr��d�����A�k1���"Bu!��l"g~�����'<�~���-8-�X߭���c	�H��-뜶y��w+E1���'~aX߅�I�p+�j�Sh�L)c��Q�T�Զ�&�D����.�ZM��?���s��"P:f�ֽ-Q"�ݞf�L���G���4��c�{�Z�����=q1Bp2��o-��/@d�_V���e�u/�2�
�����`��eU��|)n���l�J���<5q�is3p1��+ĝ7�H#��5�<�1���jE���i�Dk�dHO��q��!��a[���!��V~��Z%Z���K]���0��i����,.K;�4\t�}�����S֕n���N�[ۃ+�+���	A�MM����c��+/mWև�B;��)>d�
��oJWu��Y_!��܋431Vq�OQa�nE�{7�x_���L��0C$�}�k,�ű�>f���!��yF&��x���2+6�q�%&�Τ+�v���O ?�~�8e��d��Eh�~?��8]��M�0��d#�NcR�Lk�8���'�庰-�Y���K�{��T�f������*aAw��լ?Y$��gHIv�.���� �dj���a�~�>d��v��lAc���S�9+���-�2���p���3>�"�q���>U|��� �T��;j	E��[������2��,����x�cN�zع.!/5=�[Q�;鼀��p^O���aO6�Cr�D�����jʴ}��$�Q�Y-�����3����o�7���ֻ��!��p���w��ځL���Dv�Gt��F�s+��O�`(�猀?�t�4xb�R�b�u�k��FP�kRp�X�ڐ������(��sP�Tݲ󆿥��B9�` �$4hM�q?�l�?��y�����]a� �d��nrw&c�#�@<�6��^���0���gU���$9
��I�����U���9������HSV�	W?�����\��t@���S`Zً�Za~���:ֆ��(p4��_[�]�d}����c Ge��u�2 �SkJ��{����8�JL���1����J5-GqK)tX�1>�l�F�����Bŷ���]�M-s�=��)a�wHT�FN��w�A�Eqp����d�CN��Um���R&�y~�V�秳2�~W��7�FX��qa0�Ew��t"��S���@�Eee�7I��y�ڿ��40+����ٕ�U��I���X�a-�8dx��r�.+Δ�ҋ�c�86sۆ�бh8�9����!ַ��>iK�ܡ?L�'/��(�u�G漙uW�Җo�k�.[)�)���sW;qj�5��Ť��oO
�����|oz��=Q	�q�d��V��?O���=K�����h+ߗU*̔��;�$��JIQ#��X�W��� rv�:�qє��写�|�#�Β�J4�y���홵�sɾ�cҵᑊj�{-�n`+��ݴ��z�39�s�����4B[N�X�0�=Oh, Ѧ���76Y��$�H�r3n==��^P��+���&�!���k���#%I�6m����e�ٿ<"H*ي��Ei�T�rV�2'��ԉRu>�T� [�c��q?��,��u��@I�RB��'ak�Α��k�
WJ^�e��}�&�ؗ�\���Py�Oa7�"�R��v�g
Ӏ��,Ef�p�X$�||	%<�a1�=zd�,`!kJ�䯜5�D%er�7�oIǇ��j�:)�R+;G���%���_YD�0�������~�Џǡ���@�Wz�t=�3J�렘~-YP�б�ۏ��Ӯ")�����No;�(�kV��B�m@�2lԫ�~CߛO�> l�5����vM�����Z��D�p�L[ê�2PA6�nq��J��ti51��K����=�#���y�K����z�T�7��Y��w��&v�m�y �����c�m�L���pz�E&0#q�sIL	Eu�� �U�����vM=���#�u�8L�j��}�N�L3$��pt�:yT.����M�P��U���t#k��s;`,� 2�2��B�)%:@��+ɷ�f��(��p��o`bᙧ�S;� љ��r�		�@Z��n�1r�_~��VEJT,�H��2'n)^���$�r,�a��/�[�n�	Y$St/Ҍ>�G�����S�&%��b;5����xQK�k��q��l����t�;e���a0���=&9-1"��u1�9��qTtI�<���q�!�
Q��o(�R��{�~]
u�J,%�(;Q�]��̊�!�
�s�]t#��+O�*}�"�Ox+�C��?�'���]�>�EJ����T�`����(URH�b���v���jǡ��߾i�!�k�]�U�ր2�[�e���O쪌��lL�~JE4�H�}o���`2�'����!�a/ }�W�%��d�[��A���$	?>�v�s�F��&x�[�YÁͤ/8�=3�9�7�"y��d��6��s��N�(�m���]W4+��#x�%�_�-`Te�E+ᶁ^����FJ�-��.f�k�M8�O��hs���%!�r�*@��cE�d�-uF��j�	.dQv`VV8HjIo�}�ļ��QѶ�a�����WۘF� r��R{���UC����M=�hk���ܥ��mNp�r^�̤�O{�zo �����C�(�e'7+�Uv�L����N}䊵�$S*�-�}��σ� ���G���0�BL}�?v�j��I6�ؓ_��T����x}�Ԃ=H���h�h2���ɮ�����.�u��N��C��[rӛ�Mc�Q����?�>���DL�X��y�h�π�ǚ�q|ۙ^�e�-q$2$�i��^�&�a%?G/���nc-���a�t��ذ ��޺d��0z���'���a[��h�%(gn�?H�$ۍ�ˡ�lFP�$J�G�o�o>J�L�
7���4�����W�b��Z��'�t#��p�O���9�7��Z]К�x���^��֙���� �"�u��[���� A���<����D�bF�5>����M��O����|�Ku�z��M�+�Q�+�����/t�x܄(���Q��r�eΣ/`ʨ}v5aD@��$P:��$�5��P���������F��Һ������瘽�=����(iM	�0Lؿ:m�v�A-��ĳ�|�>�wM52�����@U�`QL��W_�6�Gz��!���x�P�=H�;.)d�����_'�?��\�]�3d�x�sy��v���,�'�Al`�D,�t��7ۨ&��j%Y64�[�6���ї�R��a��j��76) ��ɜ���w����^X��༁�N��]YYA�L��Dg&���G�J ��nY����R�_�	�� ��[�h��[X�O�I���D����R��K�O��K�ʔ<�Q� .���DQ�{*���v�uQC�Db�J; k���5ļ:�q�Ԟ�IIWc8�K���V#���W55�� �W�]�=��t�;O�jW|>m0�gmSM��C3;� ���Q l���}7��TN���� �6��uj�?`%��|@��e{/fP]�:��K�O��F�Q����i�ؒ���I�'���!	�B*ғ�23\����_��c�c�j��t���ϛ5e D!�A}����,� Щ4�d��]~��-j:O�HR|�q
��9}�:H�"!�N̓���;��^��{3�u{]�ѥ�����b{���m��]e���Z��z�N�B�H]8����٢��ElG�_��#����