��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9��m������G|S7���X� b�=Z�Q��6�;�LXЎ�����,t�U��C�R�=��e%�'�U(^g��W* �Qϐ{L�����*�\'��l���F�PjjYx�r�5a�[jf�u��X�h����$S��pgĒ��#�Ͷ��T]=Ӵh�~�f��T�͍�E���L)*x��~ �N��i����&W��P5��_Ҧˋ��!�����m+zu\���<8S���p� ]�$����d���5$�5��KS�\�w����OE�v��-��o1'gp5��/Ջ��}�)~�  ]H��}�9y��{Q�y�.ȋ12��{�ߛ�.B�"!C�XwȄ����u�㏮v���������1�e��߾bv�&˧�b'ȾS$�'�(^�)%��??�J���Ea�6^7�q��d��5�i:��~X����C�5/?��2r"'/���πσAI��\�9eu�U�_w�� o7V��[V��lv~؎��Rѵ�q6�(�K�R��M{1���39j�3|�!�a�%i�):�C(����L��TFu��ȗ�հ�
[!��J%��e�߭}*T:��aZ��i��E�7WPy��¯e�	����S��c�[r���/5��H�����U�M��
P狥��P��.A�U����kܗk�#�����C%(���5�L8�NF�bg�z�t"���z��;:��p��Q�����8r��� ��O�u핗ՠ�@L�l�NAY|�YX�?�h�*������<#ȃ��NC�)!Cl:����Wz^׃�
O�K��D����S�צ���4%�V� ����؟ؠ��"Q� �mɀ�����O���{PƙP�fR��5�����X�*����#Q!��L���R_��2F#+E*�A�h���OT��\��6]pW�v��I���ۘ�^ˉn��eW�a�e��FR!f�N(����ݎ:��h�Q���M+5�84��r�Q���W���m�K��
G�>�P%gXG�.滆�cs[,�bn� e����p�0Rhv��:i������0�m8m3�+q�M_�/�η��V���g#��ә�Iẙ�;��9J���q\�!�a�����:����*��b�AM������Q���:4����?m5���ű| w�G��]�H�!{�t?�1%��������pۂ����Ĥ z�h,1�}�-�����j��R�[gw!�:����a����[���'���R4'�;x��9��;8���0`_��Ij:v��D+0F�~L	_*� �m��� ?���5���}���"�e��>��?T�Z�XMk����>�Z������n!��>�N��#�d��-�{�:���5U΁��&b��v�d�cH���{����A�{���p-R�L�w��$��^wE�Jΐ�T"����͘��.��r� f�x�l{���Pc6�mlV��	t-�T!E���`[�+�=�}�К�,����V���#�Fޏé`���� '��z�}T����.>%������T���y�p��+����|�6��\�;B���H.��SŽت1�H��嚉���	�HT�!��ݩ�_X;Z��|D�� B���d�+T����WX��8�6�����;���H��bV�9�oGz0��8�V1�]W٨���&���rLQ`�7h@��B��#<���� oJ'��̍�kU4��p�����lm�d�;W�0��~J�%O<������Y������+e����oC��fx�C�N�]�ޢ���b���+SȪ�ށ�U#P�O��)��)Cy�1��jĕ8?sKx�C�3,ƖvzH�!�����4�m.���\�a~�j�7�H�A��1�ǜUc��{�u���v|���	��ŪB|7����gĖ��ĮĄ=!���n�D
,�X($�r��zW�P��6U��4p��&`��x��-��1�GXFLr<1��T�j�>��mp�I�c���z�d����� ��׍�@i���6ػ���ʠ������C�����k�;	9�+f2��4p�=�4�p��!|�� �c'@5�:��x���zl;��&�ŰE��_"��Ă/���m-r��°�g�i�����?s51X�>��AȆ3e�.F�$�+�0�C�pU��s�G��Y���z׃Z�1����,'�?tsc��8����B"��Ҩ\-���C���!���r0��i<R�"�l�/�x��	߳�
"X�?Nɟ� #����3;���3���nW���\Y��Q�i�A��5=��Сo����,�� ���A�<K\����	H�A ��*�,�=N��rp�	/t
�j��:����b�����S��O���\���c������9@K4��<R�}�QRAn����h}~�Z_��=��Y�<3\�m��0����&�X)����ˆ��m�1^g*ή(J��r�;��?�ܶ�����g�+k�O��$�����E&�NO���N����]~Wߋ���r�B1n��������VT����mĴ�L(��[���ݮH{�>��Z[pm`2�̸{���֔��A�J�?lSѲe�rC*Hr�@s�x=��l/��eb ��w0!�Kƽ4����R����~�+�&z<	n!^�w�Vٔ��͡����;^>/ψX��/����np{B�@��ܭ���2~��6$�v����_���^6-V�-��2)r&M�MB�R�Q_�}�Ʊ]��b�!Q�Y��,