// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:37 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aWhWPbst1wLhRKWMMOjHMGOXQMJeIEh5zGPPuUxueTbo6TznnmxH4uXKI0MydQJy
U2nH6BHg+pH+4oWYvJ6tNauBqDf1izySgg7rapqQKPGHcABBli87TlmFPiYvbxpr
Oir/6fGQbFRCt81dNb1bDPPVjd5sMpxLlY7fOxka/Kg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28752)
94fLPT8uUH9kC7svGX173WCOunE88eqHAU+GlZu9nvRHITygcr2WRLecOdmfGZy5
mZpbK7agtcpj1+pv31xrskba9TphavUOsqMDWA6/lABf8XY2X3t3UqyTXJM6vM85
vkKUE0KmwJIMXFQYq5jravbPjOMcqSxxjrVzD+aZd6JdMVCjGcs85SVChRiWzLhg
iOq0HjMe1wQ3+r/v0iVZ0DUboD9xLL5esx7D4ujdDDdDE/iLG/oJo+zJwoRBMGHD
Onzw220yWeP9nU/2LNySl1O3T0JuvgPw0YEfB3ooDkJmdTcJFi5vweZ9sXFRXEhW
Fpu+4Fa2240LzdiYqIKsT+Rc9MsRak6Yp8drdoloxumuPPJRceGi+cJyEX9agY2N
R/iJ5o/PpuCroa4bNv2ttcGSTSbGCKDHbLX6e8jEUXJbKyBPer+qkT3zLp25wPLi
Dc3QqqNPRJW6IOhjZQEt869i7qlPfQsMFSS5unmhytfouDn7dOvOpGRR1wB0lnp4
IGmRjeo6hfwcGrlMifxpVTCzHKvsSd3LMK38LDpWGHFIMNgU1E5MY49lK1y+8Dxl
g4cS6YIhZGTMLX5EoFEZ/3FEWaoSqQ9XD7YYnI3fPU20MOYk1B6aE6REXOHE/7Cc
/xSRt//KHgipSVL/Ne5UXJjx3VaQStdgF6YjEFFpqTtkiAmnWBpwmYXgn4RMlGta
S80F2/2Y81mrtZ0lMekGcOfYXlVXRW39dnwIyMSNwxZjCo8CcuUe2YHRyP1juXVf
uCrt7HdM941DEkNUY8q2txna8qvNwnFK8wNZPQLdbZrZrYB7PmeHmi3EWqEKSXOP
O+x/j2gV7E9FIZffFmX+xQnM5S5KZ8Vw1rnVDk+3v3/PI/COfT5XeaORirUGS4tn
FwCt+HIjBK9fZEVHsMMA62i/0Tg91IOmoXM8elO2iu3DN2REvDUDQqaruxgWcZjL
jaVQ95XKAfAXR2xxApBBGc0TbFSks1t4FYsh5JAxwADi2ZlDyen1XfLL3b9yq+gh
V5LkF9U/mhr9QvAEQ2FP+iFPJmCBZ3E3zJK2sAEGPBHWUbzpRvygupj0/3u1vX0V
f39712M4ujDd5Ah91dN/+ZbIxgG6DaLCfHYRj4OLU41u8IMgRMBwtyFOvBjIhvDi
+m7UsLkt9jHdX2wwgjob3x17H0JslWczXwk/SHUodBhpD3obBBgmWGkmpaccVrAU
LFQf0Gfe3bZ6HigBiC9gtWOOB55LF7C9LkIiMNx3duvbGsNYwF56SHJxbfR5Hxb2
cR6/ylaAdOXhkQLliBU6WxVLaFzenFOrNHxyORz5oTekKHysHHBjfIAD8H9sPrmY
nVr/eSZAVGXyNgD+LrsGr9AenhbElXNb74QkEE2jiSvnRglyI8FTmKRCDlNYV9ND
BB8A5Lk9N5M2JFXTJsYKX7heCgdpHlHTYoczTDa23EgeoajwjzKkFWx9nVwhQhI7
tcdIzts5NYnKZgsEOw5nNoZ7ZQPyWVBq79A+p39DNWLs/rFjqdc2gn8X8Wk4FSO1
1gA86iuJR8KwgW6e9C461RcR6ZZmVOzWbkXGYzCr+XMJdj1i3pUEAPnimia9SPnF
Gm2qbsnLNx9CLjb1w0JhcMhs1JvmuZGQvOvNpYWfnYIwqP/83yel7NDw8TOIz6lt
tMP4Hc/D5YrsmYWDjYOyBOpenECtvUEuX/WKUnJITmjHwIufMppoLE/iBbKuLwvm
mH7w8YF9TfXwgqv1eSDuRBpCH0QBfnqcAftA5oT20M9Mi4q14lnAUcIikU/ESIsa
3v0E4nHAqkt2rnqKNO2g0mRyfeFxhl7FM/foAIbGB2c+o6ITnCKt+w4HCwgKV6zY
kux/eqNT+grpJkEU+6esrNYiNHErqEMoMdAjvrauEBldHBM9vEfhTGQpKdzF4lWb
eXq8sEOIXCXp6dpCEoMy2MM5wNH4FF2xj3QggqryUNt7/n7vX7ZYCcInM+tf+Ztw
v2w5wYMcZxPtQBMw7kssmKAMJVwunOmfQrhmDYv2tj3TaFyYsx3cidM/8y8BHnVO
2M4VTH7AM/twihlIPRHX60JWRCnAaANWm/dIm0tfwOE1C1EUzw546b/kfLi/tsCo
mlv4s6MkAY9AfltL0sF+up698B4n16zyQSuQuh5ghnVbwMGl1Lwrr3AncY6I8kwO
2OhscsW64mDNtopWyaSJqbhmdf1zabaX1wZedPjp+USn7wpmMboRkTVHWVid/Tr9
LUXDJqb0THeJ1vsGl/nHpjMyh4XBJTN2LDRIV5VBBjA2cdxnwq7EOWax6WgCvvKh
vAr3lh9SvO/BbYphn2MlJ6lyEtT/2xcq1PmlDqliFIBeJW1kNaGZZY7k5w7mP6D9
o2NQhiGhJOqupx8FKPh6QXu9drJvFpZ9EtYZrwxo+3RESXolCzqqIjU1rirCVUtf
8ddoiEiMgXfrDiMkMqFspj65TDNenc/8CF7FAdcgeErizOcm7qATH8gk420HfJZt
0UHsphIljmB+9Sn1q3AlF85lN8VV4pWHHaarlkN5N+hulrNe2f+lLRb0DbMjgSag
shieN/M+xsBPtMALWATNu9bjnIqnI1PMzy0mwuXZYTs7vctlmqqf05kkrOBxHBmJ
s2DF4sCY8GUI39rVCjjKEEtL4UXgDEk/8ziN5cj6PDNohjNmt/CPcXfQ96Tv833j
YdRGFusRd0s75Q+H9MW5OfPspHI/4laXQUEPq9FCVr5XldR3QGsySd2dUm/0trs6
wRIdJICT5Hv6ruUDkgyEVR2Ak6vcn+siqzSUPINZQOiunq0Bi/H1g+BwPmM51lIo
u9iBT3kgNeHHHDkY7ESzHCgCLu1poB6Ck5RaZhv87uu7X50lHW40wfWmbXb0tvIV
oLQpbVgKnSOyC/ecoRSRI0FDerNFa6l7ZL7kkUInEov7WGxDVDQVlMjVUHeZ8W4g
sumo3mqTFdYQfBe84Mun4YzygPhAAjY6/9StHn6b6mx8cMCrDVbWdD3rQX4Xohj1
w34z/DKvSW5kVogkwwXAudPaBNSTWXCDcrcjI9iHN0Y3OByd5b13jLLs+PXWo3VX
+pL8/9OSzCMHdnbflro8VRhs/hG68uv3Fj9gyLXfFzV9ud1dwUgF//K1GNjfDo7f
tJyN2bRuztoFoJDsNW4zoXmclUQfg/Ei7DWMtVrc88csoKy3/6ixDDwMj60/B9Wj
FRkepbm8Oc0AQ4b6nEoXWURjKvUTmYGFWSpKIIuU/1bNl/DWT6sWss59JMUrbf4y
3mkeemD15/swL/htREtvEKUHuoqmAC36m3+nVwVHZ4usAdEINk9nH4h12kI6taVy
PCKZBGQQaxk8jpv8bAdGDaJoeC+7YCTqeHLVkJIzisEc3kTogz8+o4c9UIgzYWt2
JRFgq/NmssBeRyr2BOffJnzdi4nPJa7tl7L/ZQnUpnlz/q4LOr834IyOLEnmXkEm
5XVRzUimUO4EPNOA5PfJ5COhVx0wEWq1w3lk/X8XfgUW8QBa0cDGNyLWW5F2LTfZ
Cj6Fj5pF7m/U6Ss2/pGLSNDuIHFNgF5zcXZ7lxwXdesKl46U/GHzpYVVh1RCPyvQ
/ZWdpRaurvxZizLQ0+ScLb92ME6ZBGwiehmtpVCNfyAFUihuQr5CkI7sJi269VeT
iCk7+m6bNWAv9qYqTVxfV46lBCMjENv97VYA3VXrF4Ihgo6WhfXhbj/Q95UYW9HB
V2rI+nB7Q4hovyGZYAzAUK2GaadeMQrQT0P9PStfUdQVztdZxAcLlmsLEs6z7U5T
uUC3M/g7K4YVFrHPD/TTeAgKQu+t/Ju5vCPnXwAOUNgBCgKqWVltR96LeS7mkbWc
gWVU/FRCqD0uES3Xlvxbgy16wnj4fdaVvKIX8Vz846XufMVhHpIgSPbQjpXPbyUX
j5PKipAaIwTU1NYLl1WfLUtf/UM4TbiWqRK1jE0aeb4wmcoACo8plsk3x+TVjNKA
1kAufNQoM7LRBRoYLEhAWjaXxtm1bynWSZqLYMaGltGf8m93CCUGbKo7KrGsNBwg
4UaCyakcp+Rg0BDHg1xvp1DhXM2SiI3WMhMfJAirKSZv/zbRZqyFc3T1fTAJRQj8
TKkrWd9V7T5L2QRSh85QGYO+PYS7CuogqCT1m3dKBhItN5ocNiWJbgHS9r7WBLJ3
J+ipwz+MH1w6miVyTBNv+fTx1a5FiSFGvivKHe2BgVynXgxyYEVwkeyiNWQuqede
ygwo1QhmDULCGMM6qxNQl5QmVsZgM7ZcUBKkHhaxEU3GaakozZOeAZArgLOQJPto
QauXHYUzbSsZkobBB+UtsX++xQ1RYD0qnLFuqOh7HNiBzxXClK0fsWmxL1ub4fAO
Ll0cvmk0J7mkdCRRsp1IPca2pRBOuiN9w9Dar4Xn7KbNvkjKZnm8u4e5vSIybhn4
Wm+wxIVXr4bVaHVf8zVQHJmBsC8H/dL2mjtCbNHFPHmnlCYTUAuhoDQwgr2PMbRQ
wIM3Vi/Ue+3jOTG+V83M6LQ/UnQQMJN7yB5x1aIKEYk1J5QLV2vVF2TMJvfvohrY
Yc40/S1cuxHNcsIR80jWXrUB0a5x/Fm5mn+uoOeOQsnxDdc8GWdH8L9nyNe3sqXk
asOqGxCBoTNfiHUGxZXrP5jE7CnOxDlclNCOUekTaE78fpJA8m6SJ7oBFnhH6h33
djlSe3BgxqjER9Pc1lWAYFXE1PNMrSWWhSEN/RqgJxb4EK11YyzWscF6ABJyWu52
INX5WvZUUPLwwQdVPJcI8hj41gvtiMzz3m8ker0RA06TyIUKpM/Xjn353DC6Khw6
xoOSshxFZDyTpbECPuMQJkgfSuSPeBdzyL9y8B6ZYAODKl7pIfIMJ7IS5ezqjB22
+qut9AGLGDAtSeO8kkXHhHgaaMSPmDz/4TNPnGzRwcoyvnjZIdXFL8yXK5q/XKV4
w8ynoe07mHokgGD426NWay7yV9Q+eZb6fzzli869YLBvSRFwSSCYVAWvrWELisRm
LgGQ6sxvPOFrt/MV5K9gI2WXXnxHDb5q+H64QvpceIVguAzWo8aonMePO7c+rcT0
rX2mHuMMY1iyg08lar5zYPwIhCVXKw7DZy1R7913Icc6/huGlqOdS9DHOvmkj1Dj
9yU7ZjvQjxLKgvjbJBpxR7SlD1A4sxhcM73oCbQNQ7oeN9V0FP6z18bedtEOXOwf
/foPF2LREQAZHkipPxDS/WC8kaeBjfnF9Mt/8Px5Z8hfj8rzeFOJJyDDX7fAsIs7
BB241zUVosOBZ3wFghPKtIQuI2UjJZDj7zEwVTF+Rbez7trIVxuGZNZjRIN8Q6A1
qF9IC1GLQnIUgXdK6i4rk1N07jTPe3Ta92ES962R5qglLDbaHJgKRkDQEJknRLjX
I0x5AL6BnB4NTlhAXm9oAbF5gHaDgbr4FImLw+hHBKJvmpu+XD0hLdKEPewJHWy+
F4jVe9uC08t0UM+lHtSlQSjWA5nebhIjqx8kcDboH0sMXzgK8QuQUIPGBQC8htPu
erky3MAMI7l4zulqt2LU2Q4knexNpIavBstRXvb2Jvv8PMTjIJzv7lAt+3Exk1A7
ZRizbN+o3shH7twideXvEFMAa34utJwWqvUBmsb/GXeLFAU1GKD2jnfy4UuNTEj3
OJV4zQqWUuWC6fQsp8WBjsjUNWoABexO4k2uU7XvRQ81d+7d0XJDzVYVKYoosp4o
vbXIE9z1aUFUGSsMwrOd7Bg1DPQr/ilDtgvD5f61Ut5KOu7BSOQuExYYaTJDiULp
98DogGT/NSc70gjKqukrqTktI+8LfRyYfWn2PFWjYVnPmz11pJDiiRgHJA40dTT9
rkN5ywVTNmB4SssUd6a+LRye66Bj00qQUogz65FpguSaIzUPWp0zZQpzBI5CejUu
wTWt1fHx42GhS+WLJ8uqkyrh9kIxxXbc7GLECgbTXfaBuIclEp3XtSCgWzI1BLWW
3kDHWbOu/mPNQRcoHOInZALtb9QbPfiUQ2xue5ZnUS6FWQw+w5oX8VPclHRrmlRn
OLhekWb+SwJcB0IrskhzWg8FgEkm1P1MElw2+/Q95l1eooqfM/qx7qicazJw8spv
PnTvrFAqU0JV2GLvHdtovrGYHgLvcYcfQppw9hqNsVDaMeOregTUBfbeI8SYpkzR
m+rt3qSSsz2CYIFgkOhDRcBxTfFBPj2NHFhuFeR806p5jtfGSplnH3yuJVhUL7he
8WV7rV5ILvg1hS5CcmihKSwUChtY1LL62isknB1Pwz4o8VV+s1jDDzINVR4wnGJp
HoW35CMdKRyN2a6O9jv4rMqI1KwlW1wEF6RacqC6Lkv6AzCdiUVAJYpXkOXPRSyn
zAcMhZJNgJL1YE6bNKrb/+suXBTTZPoF9aM7j7FNBdX16WrdZpx5BF1KQNY9mHAn
KJ+xPIFYNcXhivJ4BMdySP6+aa/ZBS+FSNe7XLDgJYM4fYwFNXx9Uzlw6RneuUX7
mQSF23zrKZPzZdFOavIUyuMhz7ZfAuiq7ZbOIIaby3bHMAJsNuVwbv+ddr+MjJvZ
1TEKg/utQFHfMeGp5B00eg5YNSM21v+4mHx2VbKCNwb+hrXDv8ncUfNzxwIjiYHx
AY4YmymoGA9hMz4Ponuh46q4mTO56CpOkiT5lFvpCOe4DdBw13+uAB09/TT0FbGo
qX/dLkbHLWRbf52ijaBGnF1H/gPGea4PudstuwNGQgu0SHYeymiPoOINCjAOVDZ/
o4EjdGC3wLXhZzDEzB6624GovEstYADGUfbZEoq+iRmC8vmPoamr+XxKto1JZZ2i
2bJqo77qVwd0o+qXTk4cOLFcRQ2rXLB9ZhTKjZQZTVpWq3FtLeSeahhXqffaqUgR
1r/x7r0a3Ero4i5CmsVTXHfgcmF592oqUK3jf5zq0al7j35WhwbWuqGNQabxXpTx
2CjIoFyAr8//Yem092qUYd+FAFNhioZ6emvVI+6eTGLUdVPTCha1ULYbgoZa1Zam
WVYn6ua2sNL2HyryJ+VHIBCx/X8G94yW9HXFvIUVaOtewjlOnd3/T03KzA53NO/4
7tUrDpmQggUzSEh8U8IG5TOpS4AIoBq3H9pQKGgsLZ3PubF7fAF3T51SsFpBfYio
8C3snBSeoXdL/5o1xr5IIt7e+CqqsCn2TcH72v+xeJV8Mi0F+dmr7+38ksuQIAIL
5iloc7BP58kvT7LSgdvSQHhQtwc/gNgnpTVRGlryOFFBQ9c1QTwbwO5V1+8L6NRq
lMAgwGiwAXJzFs18RzvpQ7BVR8Plnvu6bBBtn0yNaY4gPQlutYIZsAGSgI3OZEDP
XLikA1sc2tkIcmr3X2pq5NvnKDWtuyEgKcPkqPl03twOGY8DhGYf45dG02Gqd83N
hcy8Cobr2NaPTVLaN3oj4DVglFjowiRBjnLByPiCDUdFmQHudnb6+n3RITgVoHR9
7CUaTYEq3/cAtdCwvLZGPQnGmZGD4cTTyPrpLoDC3jPmgVtQ8TCvbUWYugVSNzyV
RqovQVZcs8jsyWpumW2MmcI5i5mmadvG8sQkzkVTHeGelfA8VSeUV7iW9Ypxz4NL
e/sHvg9ZMYajI7rOvOiTT5yjuq9Juum+vhKacKu9sjr5GFspuqgXo0oNQzlbtxrl
CBjPIJaQluhGHdXPHzfnF4baB2eddP4DYZrADcTWAfECx4NXOoSB4IqbDWxwfcMo
61Zw08s6Pxdl53+Yh7c/uKpORddjuvKqItmi6luORe7bx2+cF7TfMfNbD4TjHCyR
S1Bg8UqQ95xHRcazauRgqqW/CPj6Yvyh3lpIMFMkjnwZN2a3XsBBf6id0qp5Obz1
TfQn9LJ4qnppIG1AmPET0JQ2TG1xsKFkPUAOCIsmpQJYCVRnWSrOStOMBtSODPa7
xPtTzSor7xHYs3TI9SJnuK4DJjFCIDMJk4mmDuInKB2re9Xti6SVLY5NnyDKeUYR
TDcMrbNBi9lcriMA2So3MvE1iVfueXZzrQeHELy7JB6PRb3lOSeU5RBdA3UOyq8m
r9663HcNElyDr3fwmGMeZfeksvbGQARAM5fCm+YLBYNbfjOM7N/5sSlnmlrRuem8
FmdanDVQTQCnW3uc5AcyxDd/RmQO5gh1W5ZWzYzfJr0KI+xxGCRwmZFPhtEFvQXJ
EbVEbZoyyJalMFvK6Uen1T/xekLmRo+cJRUSR4uVe3QDHWzjpFGdtwns9HiWKDFR
JK8oTJFytlaCUftzuGS4Yxoy/MRha9Us2Yf1dhzS8vUldqrQiHS6vgoSqbI/j5TW
CZsiiwK1iQpxcVTZl8Tna+V0aKL+GiU7vl5eleQ59VMrL4TVP7hdNqdPFm7vpjtq
YGdwb20PabnaTILkY70RxwrYvok6ZMyLn47zzHxSI6xIfE3ySveQOZak+6iSOHgR
fqiQ2T9AvrBOYcRb5HTrXowO0BluYjYsROdieWs/nAdyi3PT6T8EkOmZAnCuMSmE
YWajsVqf2HYC5RrxybhKtDTvprtX1MUkVE66hGgIOdc07WODXy/kd12AgoL0vDHE
8LE8Nw8/w94BPU7N+PgoTgkglg35xtFkk6Xvhpxlgi9S8Z1twM3x0aNk7iH64O6I
MIm/+Cvwml0RawDpEvWeCsVPbpfFm/dU98iPCLFPZGMxNDP9H+nFW6JnsYBmyV1C
ngh+8lO1OVnIVLwzDtlLP9MbJFhKbH85IFrNHfDtN4UVNPSKDE/L0Wahdust0ID5
dn+YQ4kwM5u+hY1Ec1VBmg+D3/qgemiCLLrL7eGDlmbRxW+/wk+Jl557YW4dWWcS
woPkUuM2Eh3IBAEPKBOXxC+K0oUkWIvxCtVcFxuOex82vD9u3QjTr2iigmSh16Gd
CdemNvfyTsmzHNiu8RvWwnO6qWLkITn6lY1DuPhBplG4Pwj34jtnT0IogHAB0hrS
BAoyGdPEL1DVJT9x7IVN/9TxMLOecepADlncHHZjC31GlPeCEDHeB+x0rEpcy2tc
oc+5h4Ik73eJMUKAXwyon1pj5FVLWcZ0FcZ8WJrjnQn3VnkgiR5MiDse0oNyO07d
4L9Mu+7Zdc8AOrsYEWf7Z8U6rn7bBa3nd+/G1fmtbrsfBiDsJohQT8MqgIIqWMH2
EoqbD0n5uKmPAv6HSTo9pLUrFAte7x1Tm84eNBHOO6QQJUZrMmZgA8xX0DPtJgZY
xKQ8OhQdwhnuUdzjZ9B0xx2lHAbJYP1FjGQcil9FN/YzuXVG9Mvlg4zJmgLG2aCM
f0SYV4guBzgRzwWi2UBzlNmBx1mHVSC3N6rxcjvKKIvgsFhfV9x8LZCIxt1kBLOC
SPwRSO3xZG/oVQd/tbHIXJ+Wbso0nR0a2GGdIxkdljsNWHEHrFOx15ZEm/9nJMyc
HJvf9pK9uXMQcwYdxDa3VJWqIFW9QB31boya5cUTM5qJsU9NNH/gv5q7FcaZgj15
qsJ1jS9Zn/iSSTOQd6Sg9WQYo9bTY0mCNPExmQEzINJm+UzhRzkjmhmuwnPXS8XG
B/OqgQnWjZsxyREIDorpUpd0ihygPWBKj/lXxopxCRzlWH9hTLA6v+7V2XzBk5ly
qyChCR5/nQqifNNh2EcYSqpwKxHYvEAJb0ooz3Q4Xf1LgfM1KjB92vh+7WryFohB
/m4k+KJZQuxBYtba74gN8LSqSkRILWyz1MpGJJ+YfERQvTalWDdxx2T6ckkAyXsI
CTRvb25JnM1ADunxiE01zbBS0MCLqR+aR2znb7z97uePVa6U9tkPIMMq7NJuam1K
yBPzkgxSrRIn+KxckOPVypE6szi1GcxC9YTPaGeIU2BIBH8k3u9hR6tBfEoWfrCv
Ak+TrGXzS5fVBZN+NcBR5ex2hKkx2FHQiXdVLuVZkCWRE2hxUZNUVkLw+Rep+Ybu
c47+23+UwPg/BtsiphOVZXTtlWyV0zaR/kYGkyIElfzFWUadyUa2jLh1AEkmWlX5
Bx74t61NSuVLswg7q0rhXbhfKbgtS1qH6kSyNxF7xdoYxLI2mWArbXAc976Fcd2S
ulKkfsYEDfIIQL3bqlrvieNOhS6fEk4lnTrav+wrqyqIXvlBOA8AW3el0q4rlbXW
M8NErcx3P80zGldqv/et+A0RHEqgyjNDdMm4L7XRM2/ddg4VXkeOj8Vd/GL4mH5Y
m2+ct+mWv78//cyLGyKj+sO59qpkOc69jjxkFZTZyRD6aZYvvloFfWSL8uTLg+wN
AflijM72w3WlxAOCd9/Q0k8FLOyeoEqBb1kNi+XlwwlkeHzqCqaME/g4O/vOhcWx
V5Fc0EUb/puT1+mwiPY/aIRUQc6VXy+UG/vB3tH+XPsxr71ZtvyJQDXIdFUfUST2
URX73CVH8cI5C41nHjtWgVYP0snmvVR4knGUzyCczParSZfcxBLD51PsVSoWushn
seyUpI8W//y0Uvcx2hGfD+byHVQks8Svoqbk4vrOvzJCZF64haeYCZyyB15AqvEA
9rQaKUZJDywGY4Cj86h6MJ1S1svD/XsDMhpEv2/bhG74JuKL31ZGiFP8ZAUuYvoZ
9+8rkHLzqi8o4btHqYH9NpSFMjXLduNs5jrkOfAxq6U7e+FPi1ygKlJfluRPwsFI
mKHcPYvPy0QlTOU+GizBHeL+bE5ZKRQiMhAKZspHhH47iOBz0clpRqxukpXw7JkJ
cRkpdZo68iB+Zj4lVDdppWF5XpEZJ7CYnwYA9SHQIQjWTFg9/WkscB9/yENGpdI5
k9zmh3RnyuxoewXYqW9k78e5qlf3lwR78bybZTZnsm/G/3uYE92udD6Hk2agY+m/
kuCNh8ewI4LwBL5MSBg75sfsRdDSZYrUXgfbZJWHq9kKCpQx1edI3ToPQ+uI0qj4
xYK9LWaUDuAXpZxIKsCicJhaoIuAIZaoAIkr2CLGgvBVaT99SLZ7CSJDgT6Uhl/W
mBknO2P8wovnDmhy7PTAVqHPzbSrNFlwA4Yh043aNeDkrbxQ3+41nF+BWwB1r+xA
sPoe8zLSsbI3e2kbt2MbXwHUI54af7/dAqeAY95he3WCHYNbsxKkl6hhtN69IYTk
8OG0zZPrJJOwIU6lz/m9mFhIEuJ6pafPPJpijLKXxp0ObCCKrVVav5Yq2uVrd72c
QAmOkQXYtYhHK2yL7jrhrwXK4bzeHv+JW4V6jghJUWBldOP4rFYo7rabJlB6aWZ5
SdRWNg/Qq6QlXukctXKq/uCliK61wpBZnlP2+argsfsj3ZFLPwxc7xzVRnNdwg8d
GNLY5iNb7cDuqShVs0MbSmoHU7CC/eamtyDJsb9SsQfOqoKiYZtbY3pdgqv/J/Jr
p50p2sJsLJ0cxZjQ+rBrBjg5MlxXexexMOuhSWeSHIMQuPQay5pJQEUW5EniJxbf
iw9kG2xUd6/rzJQt64ek303J/y8d8qk34Q2iWBF8q476kZVlo8B++q15HT9aDR8K
xdExltr9BOTYEeZj3+4s1wxwiI/mI6r5HNSrhZKxYbf7Nap7ehnQCbK4OBmkTBb3
gEzxtA9Tu54o5mZMNYwf1XFr3e7oTQAYzonQtDCQLohzMN9bRtYRFlx1P2WvGYyI
M01tyCGk9keJLfmV4hrKp5x+2s9x8HcysKfuMpGQC5LFEg/kinaWMt/3KTuuBq8h
JX+h7SR4PqxAujoS/cliNCSw8RRtIdGBFtqNNlsJ6+qSDHn14VNnhjMY149ZABvo
bdlbK0+wNr7eSUq71ZoMw9UdsB+3ESvtOTKevfyUgXQrpOE2LiqFVtJ3hAqc9sUn
cvwR9JdgDyhGG1womSXDNkwhGvIbnk9MHgtEJpHOxhERdgZPnxqq9+WSCggMafrM
mn6uoZdbRjO/6ha3kwa+0QVDeq5t2rhzWJ/Yi1RSDROswCAt/itIgfVTviYt+Bgy
arSiX99/BqziPr7sdnkb3iHaTQEWtTq0n+IifnT99niymFdEa9iFIDLtLoJJDfO5
GnqQLRuj+Z9Fw+Kx2sgDOoYAILHLIPMgjpvcPsoFXfEhqTtdsgqF3bb4YLVz9bZ8
m+KTJkb7+KR5ZdMJHx5+v2M/GUWGooGqM1rijNp8jkfTk0hDMIGMCV/H8z/EvHfJ
pK+J6F5WeWo+k6UBZqd2PjXsl7GxvSVwqHrWbE0naSK3y0Gt5jPc4MR0RNojF6en
HmcReqofIaMUgXORSmOLgDCN9oHDjdUV3TXLKWOvW+dvnXVchiIIcpHPuxavlv1C
c+0bt4p8oFOwstqPp4e24jR22lheB+/Yxq4p+MnyzTlhsHGHD1izdOK79kK14iiM
KSk0JeUqqUr70LCdDt4IFuvq5/VZrRBoaiMBA8+UZlMpCdgWkNTO9kf4tSqOjPqD
jPmWvSWEruURWrQ3lUsbVG3J0xaXWk7GaGmWk8riI+8JzdcpKxQVxaCoxoI+TMPN
qeDrQyFpsXowHN5UYlnY0lhNEg46cKFyGGd9QkUe/xv5ijtHynGp/TXJ9yFsZXHF
jhkeX0IcvaJhxV+yEeWiLQ+w/DeGfW7EfHTtGcLlTpq5fEpNkdlnRkJw6f8+eYUy
QUafO4WOpV75DWdrrYrfErH4xPdkaxeWu2D0t9NyHfkD0JE785PRQqD8IBM7CKF5
M/3EGDu8hg1er/fILPK8rrvhrSoxF+dmsPj/6Q/9GUmWdS/DmtciTLgOteDMg+cm
aAUghBY/2QSlWuDLDzVJptWqV/q2WvW7vv38BFgMeVW0qxFgld3i3zR5PEfHcXj/
By9TOYfT1P5EgFC1B83GsvBRGjd9JKwGYw3P/yZ02XegI9Og7sXRlVmhiAtBi3rp
GIHZBrLcty8yMrQTfgWMbWK3wjecQF786Yk/L0Dyoh9rt6YzRQzkcu3a1zzfO66B
ZrBaDSpqMbqcUO/ThGupO9a77E7rIi5jBmW+A/ujXVqaMoGgnef5JWGmtO4TyPB8
JeUofZ07oTFr2FHyk6Mu3Rifo2E0JNbt911FA7qinSIR4PWpYKZn7LgkbKjE1Oum
RHUolI6I3yqDNKPaXrNxDxbb2D4Hl6kygqkYp7zBxguI8Mp1Q7KnqIYYDRF6eyfx
JXFBzMdvL/y5MIAc7PvoK0IuUbsqSxMIvE3yDyDeNyXMAEqXb4dVS/4aHyqQSIx9
VL2Kmkv7c/9m4QHfRutVbWyImzN1cjzPsm7auVj1aLbhvFqozZUVwnmyYgneZWmi
KTFVOpb2VaNQwfwynLYPsmORBvjhiuh17NCf4sQpRg21cTyIsx7LFGzz2zSfHDQz
2AsqiDjksxIOekj7zkdnBg2+y9oMIMZUyWyHPfXO6w8Z86uDaThnOtIB8Imo4WW/
ZlZkbBO3PGZQNbQNHB0lp8ZzkETUr8J9PVmw8YGPetkeHxOHuzTpbXhYT4l9xq/6
hQjl46DdKDNLLpdPcNy8Oq4xbxs+AWfEpvPDnT0LJ5qHSr1nw9wExOXjsFj+NtuF
4yDUGpwIU7dgG2Qn7I0E60zj6z3x00mHti0xQhdtXDhr/xm5U4/tzRhkkW2nHbZx
/3ae0RzJ6hpFEVtry3D7clvigRzYjKSMfMUaJx0/+V93lGEWPC1w8eORE+mb8/f5
pyDWQDNocgdmJcM/tv6iK3J62STjQkH2SZMZTh76aSzn4I8tvDtwHa8+fGyHm/eK
QQJFlAcpa0M2XL2yXKAB563ImGD9hsXVC21rCYLLblodyzA8M/vzARbNXdgNgy6V
dVlyAzFElAWYmjbdLVKBeC52abbAs19fp65ksGxzBXjL6n/MlaPASJb0pp7VwcUY
Uc0GWt2WpCRjWM3wl5lwiHO5V7/86/cxBOXwaG3t7Y4RBZfeTTO6y72kyFXvyTij
0sVytJuueqiri9d1fzXqmdXc2cFMn+TLV0Krsy6vLpvd7vbsB7t83WI/Eb8Vz50j
XSGosd0raVw2c2Pi08q+qVOWTj3cBxR8XD6waLaTYQ7aFJ04U9/M8n2gkyp4soNd
UoSeBlNodWGeyzcPWCwLLzK+YO4MrLTjaySSx057ac1bt7wZawSfQfqCJ+MjK6WF
OD8YDtWySheEriITIz8vGwhd8p3TczMNThEjohmSD6BrM8dUtpK3g2YNtKHgDN5p
zfn0R6UcZhHE3HxePEXdTakLsu4NnWF/tj+ULegJXX0ZRqeNlrK0Gi7r9APYd5eF
qZp4NgF/HHt3baiHxz3jBMakjbuknJqq1ZL8LHv2MjvYPn1xIKq0+97nyGUTABe4
2t9+tnMGODXsBxQ3GNNwFuQPagcOop6jo0VafQYy63IISM8MCiFwNF695HGsi05X
SK89P6cdTTombZFMhtEaYbOgt5FrdHds5T1lqGvhkFU61I+XuWdMic094akqb43O
ednU6AWeWJxAFaot6/pDkb4JbXyDss81EvbL02yt4uJgKwgyJ8lcQWt6xZQCoRGV
1jCI6FiNN1ZsZK96jLG9bfddd3GRvHmCz/6x3Ifxgt0PXvSwG24begWphpe7VoXL
gajlaUTRqb67tM854yWj98iPN+hApwMsvVrkDpZQjqx5zXPUVz99ncM3JYJbpLRx
du2m0HAmGFexjF42nQsq151ahnrGzmvvXcNeWyEPvyIfIQCgESg0qsoselsaTsnp
8hTPshXDidBvZ82z+GD9mSt5EdheTkGDFwOsfCoLJHsybTZYFbq5scrYCBKyzxhr
W+C/zx9vrhbxPEbVnrmpbZlO0gT3wveFMUHqruads8Dz11XrMf5pgXohEO0k/I19
G2hbggqezypxMwRC8xUgqqtKjv7aqrzQjYJs5l4IxPEB7QC+cEmT5Bb5zjvCjfTu
6/ca7wEU/f/yUdzbqa7nhEgCMGm+5nYF57gW0dd4711TBhheQduMvsot7h4ikt5I
eFFqBUOwt5xeJKGcTo4hxbixRISA2ZU33s5Cn0NcpL2bu62eFzeqzlCpHdHRjBaC
DxAZkiBXcTsahrba9yYNXqelxhHOOBDxk0hHJzym86GJ28k5q7sYtUY3JvdnCkt9
SXnNl5Fg8/75jLBPn98qGeDc2MGPQKYraT2krxMT4ykhnl2cYts2JBz8xQO4tR37
N+UhH2hOK2R3MMmuDuHNcBiq0L+VwWamRe+mJe2CFYsQpmOtjGYILgBHXGs2pUVm
flEU9K9wCjezW7Dy1vZUc+zx8vIBQbYHtTaF0tExE0m4OSTzz/MQaBXvDEiNJwR9
YmDjICKfHp28bXQeCSXuA0/el7vrkUdpCvc/b4wIdMjz7JaGsCPyGOlr6kEovyA0
2KA792HGyPy7zS4QtJk2UYn7heIueMbphu60rUzBffFdZqnKCZTkNch+tstZpioY
BWZTwLtgFcwmwo08PjEaNq6ygH7/V0DT3mkODdzMZOW8wkcNz+VyeNjRFqghgJ7N
0n3AwMgKIrKIpLklRkzcu/5McaUETsqh3d7/4ASN8bcFiALLgcr7zJXbQtm5yVGO
2MaA6TY8ipZ55JOjoyBplWthR5namIEHvFjAhxhk4jPUtr2M7S54J9HiITfQRIqM
i1tZqtEHs4yoBVuWf/900lgTWYlv/9r1CKEzIowID9WxnbxmEIvs7YhtNzcLpfZS
fbcH826Ti/dvqWSFK70JhleQHBG5lwaqFjmW/LKk6vOyTGzCdFrMbzr0zx+5mVcc
crKJISLomtGfLoWoMPNE11MODeMI/YkX4c2fjOW8vxskV+6aBuz/P4KUGAyqDKgS
43Qa8ETG3tg+SeMN6rUeKAW+lPUI4p6JUhXfN50c+pKT+F9fTvZ4SwKygxWkP3Hj
skVyRQiIUEGCwnbivFukYS8vdyhzzZbJR7iKZ9HHyyGYkFaKFn6xuWFEkTvUZOnm
yf25SBHPwqtU9prQH7g66JZVazyE9c9NNtv64Z+sbiMucLqsO6jX3Ljn39kTyj0W
cp6GGDfTsj4lPRAO6MLy5XojHwRV1ausc7VtJXwmGpkSQmiF0VU8o1zSP7QE+L5i
8Lz6Y8OmkDeGnm/N9qVoVXtgP3A33sKGu7JR9woJIyXddzDMp0MOiQVpJ9VPG0La
jykcdyTRYxmlh0b3BWfV74DvIFObpkGkov5+B25+wOkWjsQsOiF4KHeSJK+a5TDv
FX7e+8UgSaKdiVaI8iFg8IKDCxZAnrC/OWNmAgxfJ7tW+T5oCoT26R4DyctIACcV
1tgR9IBXyhHMQnBsISS0hpqAPNdOJ7o0Q5KMrHjUX66mYQmbTRUBxNwNtrbYtmaO
aYa4t3UU5vI9VVKbmY+d4DiDz8oZe3BdCXjJoYDQ4ttwIczX0dbXjZpx4QjRAFfg
93Wb9Z0hrGmGhsaYMVWiaRODpBxJ/BYoR2KJUUvVoG+YVXe/39GY752kS+d5rPq6
SNP6ySIkg45d719fHqaSUXbaLELs9YyQjznG1WECXt0sg26Zo78tFu2wLzAl5KMg
SvjFnYKZRt1BRjdFFzkl2gSW9XCSYAujjJ92hBSp1sHU+yHZC1B37nSHUzkK2Gab
71qz4D95kG+ojzGrivYiEN6cM4cfUrdIbY26Oez/OO3k81SQfu/+QFT3nT6tCAZm
vK1GcL7C/tUrcC0Kj5UR7zpEG8hX+stiN4iOEH/wtpfZbG+XML1b/uEbGDV/o/Bo
251PLWtdBVRJabbtBnXM/+Ca5gTToEFi887/58fM5VwQY88KR0XUa4LZ26lnpDqZ
AAryRmWSwFV0l6r/hc5DaI/nYBuLuLvLuhMRFw5wWFM4mBOI3mozT/VO3m9UeAPL
Q2BemnPpWBATXEGYNMOBv3+Xu0OTTpSuacCb1uhmeGwACnom9eCSNcvls6jYBw2M
oNdnhsZH0MhhPl8KzCLkK0iAq0Kui2CXNFaice3lOT8JKHs5pZZAgM90cfJTkJlP
G5v4Vxc+fmTPmmmVMX/56B6h0Jw5RxHr5Oa76st2eliokbxR5dOYSwJEzzF9C+h5
wnbdSX8rneTvXUDiEiU+aHDdR55NUkvf472cJ74Vp4rbZNOpx7Wc2dFjDBX/0+cv
OcS+gBlyS7d0XsAsXJ1sqcupANeJ7IZBw/Gp3wutCKmLhLqskuj30cKNLLZLVEYj
cxLtzYWZqI0eL7ZdWxghB22PgT1wLWHxE78fwaOcopSe6a4yQqzDWolwHxfVYl/6
3LRb1HaU+Y809gjM9Z/9sQmsADEC9bnbIvc4sjdUhKS574Ptv9y2xxYZZ1qlqEQs
hJqZLoypJXp1mA4FJb0OhLRmyURq+B+zFwVp210QxWjL/V1YaZ4PyY3D1bC+X7RI
l1ryGZFRftAtGmCGWxfZBIDngEqnOMMChobcqy8cRvAHFa7qZzAnlAHwMgS5uuHj
7LycN0/c9V98aHzDAziVhoG4WKwty2wHJXMe54Kg+ejYbXC1RiO6C0ySgCqihJE+
jvoPb4ILf/xTqQbfsnjT2+xwymxdKJvR78H9dBZX2fNXtNgKTajUxYeY1WVB5Uom
iao9WPNwaqg//kFqCrpW4+BXhOJasbwrJovj3SjROfgdpcrUE2NvFQpsb5JLLPVS
IXlnwaCjalWFatu8V680DG3yFomGrkXetH8i+9AbKzZGcRDz6I9hl8Ou38P+nQNC
JVP5As/BxdbsUnje/nF3yUSUpRBmpjdFu/wlPnHMV3/yp898SHm+Scb4PLCBAWAS
22503MRfxKq7mXe/pr5u42BRoj9UgMiE+l+7MNQvSotnpJIcosqrJfRKiflgCcor
fp3w8+wDBW1DGvBGbwv8Elh5LSXykaJy1MBI1Iz+h1WT/FgO7nYMyymdASvgkI4y
gRekluOoinNJzlj8W+PesFxu1/9QECdHCy96XKQgeX982Z+SvyLTm/ow1tR6nPQD
slCgf41tppu7pyKjGhVqNkjOg12Q2u0njvsBXgAPkY77Fym+nVobmAXDap+L5kwC
haSI1Ah7WYkaVmbHIKjCagi0ypIK7/IudsR92Ix5i/HsG7Veik7T/yIy6N8aM2CC
LWmWyLkblEHt9VU9ngIhf4qfvONqZiGf9XKBwOMKtfRTZupVmjJ43p5o4f9XxMov
6CLrd59UQ2BXAlP7xwXSzc28keo0kreFIakspJgeheu1/011cCrTc3OZUf/L5yk2
CJOJyeDR7MgEVrE49tkMjW4meeAoqDzl42Japsk895G+OrsNN/UrxyVNyyydOAFM
+5rPfz6dCHh7zRYwC7cWRgBIzt+Sv4hSA0f2faFG5N0YtFqQgwChYmYsX6v0L0XH
/1onWiLPUGh/mSpLxGKOyM64YfsEkeyF2lISbHNGNYKq1ZUN9OT8n0pb9MWl2gfV
vEQOyOeqBKZUYEwSBl8AIOkBl5DbKAKpWA8VVUIuGmHxVaF2iRNyah55a3hnAEgG
7roHpruf7F+nVw5szU/DxcitUGbnqyG5NWmDvSJKOQ99hVwpr35spUlD3MiYuQJn
UgBhzVKqdBUTX+5T4tpb+ghrtJcM+pi1tR+yJUQq8DDjmad+ATBciWzRFDX9vDp2
WpK2zyn8BqJ2hikIv6qwo5Xs4bLiZy4pVKtKiGYTbGipm0mdQoOsE8LZ6Q+JkyCM
n7nEP5afYy3MjriZMWz2QSOdSPFdKAluKLVpo/C1VyJ93somwhWLC4izRUuX2uDZ
78w2Ss8nqRXgpbnt9WtVGBb2M27h+Ffcsb/ojEqJdT4JBK//kkLFRQxqFhxd0vr2
TE+w8yno2oHpdhPjta7f7SaEryE9UQKuqEkk+pjRbUKT96KxjoQVW5Ynmc0oHjO/
kLj3pLJ5hlCpcvJEWOB3WKBaizlzgNdKm1vbdlH5ZT6l+khqIHVlC3q7YT+Wb708
jRkrsAWOpk40nQxXM5LvdmZmC2hTp/aLT2dkW7NsB9ktiI5qRPcyf2ulRgkpCoOo
drAP3uTkN+34YBgHDG5VJM0CunoKc5kHlxbIqX3HmtVR6Blz1di+HCU5Ze7Id8it
4a/syBXQfsJIDb5P6C2QKX9ulxdZtB2sNiCMO3iFf1npQAkhPcyQ5Hh3J8+Gcqc6
fFlShW3VeyUYkxLq/w4on9mHajrqcH8WjF9H+hgIowHHkREL+5sQeMlK505lwJTa
cvLD5KfWuVJhjwhn8NjPIyVxjBhnr7ScTJxi+Ls4/WGd1V7XxVjV8Nf1Tl0CtTK6
AkMkZ5OxQfrJCxrEh/nJV/y84t1kVj2mcl2DYxukmq74jUf88/o4XuQKUGZJ/Y/D
rFLtX409RnyfWhwC+6W24ZUOAx959C0ysuvJwCiU6oWdJaSlKgBsyzEGIS3KcV8T
N0Kulo6N2lH+Gq2T6EYgvnPIhJzyIi41V4+2AJdHY7bLpHD3CAYLdlakvI0uwmaD
p0R7hR7MU0+7Upr0p+wI/37LPNWW7OcGfKS4Z6HNWT4Kq40cew7npn7ris6p32PZ
jybGQNBXInPbrCUDP3w7NCDbK1/7RpXYuSIR19/zARjXUKH8BGfC1A5ZU7WEEjuF
q9KxBjz4NCB1ACJvJjAXLz81fXw6QDnIWRyyu3Ji5UQNT3m64Dk/X6ifS1M5+Asx
zJuejmltwBumgk3Vg23BR+FXCkjzKxOpViLJbygd+xUYMwtnR+JKNDoLwYyd/XpH
B+s3QpUCm5F7iBP+5ZngYPQwlLC0utRczyRxfU8ZSfQXZQp9v3Ba4elf/8d2vHhZ
25ZH8J8PGOmOqywGn/wy5VRNpApyG4Ne4uhe6PxAcCkg9FP3kvB4d7mnbAWJZJeI
C1tMYReeg1OeD1mzVlvQDezmJ6V/V2YBsunGeoeRbrUSWl5qHvJJ+4jahNCidvIO
ivsvS8B+bRa6Mpa138pMGnNcZe/gJc/pHCvliWdrTgKza0919ft5Sy+OkEqjfgLt
ja6ZNj10cGywqKzISz//J+ha2ikCje9dRXgkr2RI/4qP3FLlE7H8yBoeDOkSOlrz
bFp2f4+paZ8wuy6NeOsiSd96OFm8y5ljJrMBPQs1SKTkdi9tLG7/5RBk4/P3ezm9
cykigzBzJmxZrz7KiUMRtmFRlXL/kuj5NpU14ddTw8wbgl5Yplfe/LGByizvHXcx
SDGjiUfpsPVUUmOMQZPM8YktpyOnIs6nlBQj+xWmxtguIEWposPZpIqQgDFk1YIh
CKt6KwGNXJXdxHwj8U/QqjSwhEB+2NfjKYQH7O7GEFgN+n/fMSA51M6F5l4X4IWU
f2NVcdFjoeAidxwUitHtdWePfuELk5inZZUTgki17R9i8Z+2vU6JFfDBiItwXapL
gmDyOU8depwp/em/Rs4twMYELgqeVfSGBz4LrbTYxZykBC8T+ueFjtmuvd9et/a9
W/GP2Xf6N3F+Euinqii4udSheE64NJjuCNrd3pSnbc9bKR/edbY1t/rJDlNrhu/P
a1zC+hy0embEu0J2WAH+KZ5iHN8JOSsJGHFp74L1BxJrJ+2DQAdPftwf3jbWb+fW
hVPZQ4nlyD1F0E5v1dRdUie8CE1U92POxdAXlvSOBJMNJa7FfwoH4ZGXWCJk7YbD
hSsAUVLccT6VmiKmefOP4W91ooPsHAQNZKIjCpbGxTB7JUSHZwHyr3jsRdEWOkY2
osRhNvSL0AHIhQ0KYI7YV3Js8VRrcH/hMLpHVPqApTMuDqJNAhURkR472iISaRGn
FyqXv/Z2SsP/B9DKP6C8EOCJ1UeCwBjhaXTv/n8iZYCdyVmKPehaYXYXrEfCSRnJ
zQsoEErGaXWFGHiiJyHmcPhK7hrJ/rksD+Orxc+NyFZBfHQJLmHVpNSgCETgxNaG
NWIoqs2Y2DnCX30+5mvQQkSiReyxBKDLTdTYpxDNZKRWyDlUA31zsJCi2IBy7F0c
FZpogk08JDOc6gqCdmPs/nctJA9obIS7080PlgEixaaxR/Er1AcgC9Flp57tfzx1
1dnsE/eMxAToUfJ2WQgfvtqoKdpWFQzqDLFPLM8M8LC8ArLRIO5IF2BqeKtA2kfv
8G/vsXgPi5uFL6IAcap9uC/Gn8IfcPg1lfeVUJty4U9Rn1260Mqn3ElUNLVx61O4
N7saI0/nrcFXYSOo11izNEMnuFVbMDcbCzmz50QZU7C2vA4QxX688r2qqgO/dMpV
uM1lmFty0yZ2wCZndwybWVmWoyfstKUzhdzQ423M44glwKCUus1cYeDxW5yWx2uY
rzMChwgk57QMOEjfLC6somxnTYnW0SOWd7xeeSgD3+BicEt+PVVh16QttCwiCuIT
pkjptdZT/Q49kFQ8KSOoVthOvgJP6BF8LzLZFhami1JuBPv+0Q1dk7WP6tgtjfoV
96sDZIxUHKhdfij9+iGpIHhD8XMjYu68eDiNKJ9O89k+TpJm6kuzB26y+9LL3CyW
Dw/ZXfPNb84nb67Xv6VxKbmaopyS2LigYelzk5v+rkPa0GtQUD6Z0kwdKYkvOYy+
9RfVobqtC94OPcXpIaHWLQwCF8OT3r9U4jiQ77hhwNupQ47ZuI0nLXAm+l/l1gpl
+WBAmqORm/B3vEpan0YJtM/p46cnqvePMXfRMGA+ldrlXqJZtIOS85UivZ+E9POn
2HW1hU3Eqj8fBjjix0mR+y8M9JpSKTy8bnCInCSIi27jKmOtF5G4kqEwQ8qpdNI1
CKotpiBtIMhVtKCBRzh09HabmSi8ZCaqNXfeEg7dnkPatB32OTLDtRaMqQd277jy
MBLKNCwZyhNrgSw/DvQX1sazpbBPLrnSDjVdUnDaOAsUrrmg/nuOHNezF1HB4fSw
9eoIkcr7KEPnwfWxg63/hq47uGR8Qvd4JyTCxkrowdngMFuNxm38sqwNEbsLgyXC
cNLZ6SNqr4ls+5DDLr2XUKIoC7ZUOmF2WtY1wFxdgG/CBqEG5O3DHBWyJKpJHaFp
OEy87utOQ9kpDK58eJ46iHCbeLHdgFlRDgn2KjGQpziwvJUlbTM36fu8IJj1dqdf
QKvhtOL0glHCmBQQxqlpwj0ZGAZSFY0MtNYNVYayPAeGTwThyAJx8eAZ9XjrR4ZS
+yROuJui1Qh6J+j9Pz5lSHSJt8qfn2Pk5rRFND1P442O/U8ix+shH5WScn4j7IZb
uXrUb09VQeIh26bjHQ0Nkz3mA+cQRFSTG7AmOKhihRBv45X/jeVZqjQ1hJT2c35H
Jyo26RFffCFRnuy7OTV6HqQ1An3xYQ4YkF1OwChwdrfjb1XnYS9TRjmk8mbm+ua9
VKDiRC/nuFq0NHbb83lL+XeIs787v8J2S0iSg9tO0BMaYZ7o237c9J+4uZeGdxYO
tq8+eVapcgP/RNgeZAUBkwyOzY5lMifOWHqT0nvG3qY1h6B+IuY1v7jSILSWTi4g
O4v08BA6xRR9a4JCpSA0bNR7AziTn+rMsfApLYcZE64AaC0DRPGAJXL0lpf3sFum
JZPbu6+80mLqhINVxEJ5ID0NlBlh5giuHHn8XtoLwB9eE++KCJpZxBvMRPwG2ngG
sx3Vs28KLAik0sVr9DtHLnq5zpnZCGjuE+RL1D1zRTLN59wPpkJ5dDOqHXNbUPcv
Ov75xYSyaDu3ZX7mDmZjlGLrc8tuOOeQn9iEwK70vzFdaR8he7IiIyB6gnUHSPfE
aj7Vbr6XN8KcbP83r4RlLiMa1yfTGwPRNAOVfb9aUPZU7e8Jc8o1ursNdMGvtnAH
6ITsmozXcuNaM1hD5RU4Wq3zs0d/n8wSK8AdkfwmewGgWRaKgsVyEs0EyYQylu7J
tGbLoFMkNXxuV8GyyVSQlKTA4xrLH7ISPe6Zs+NCinvgf8A9Lb945k2OLdWVnPXU
GqXiWQGpkUMGb0+i7u3//HOHzZ43urwaenWBH2b7yoZ15ncf99qVWzdutHXlWNhX
cWoDBPTOsN5V8czqIdCTj3Vz++B8nZBrojgh/92yjn1bp/JM1XNLWWRy3DQ38+k+
aMz29HJQYrHU/I7H72/up6RG0CYuiDU6+QB2IkJHnH5vQyd1EPa+yQ6gt1jbRCNd
pr/VZEAkXwAPyMHDMe96Hzyus+xeQdyAIqcyyIzgRT49Fi7KIol4tKAYvsqk5anf
j39w+upOQNbFgDNTGjpD3f4IT9f/XP0drHqbn+gQNVvuN40a0g3Om3M5/kaWG9XG
dap5rgdUycNbqcpAWkISD15nj494B0NrjyFlN7CgtF5QIQFhNnVwNXwW2/slmamU
jQqNzsbGznZ7VVMpAqOsoMRXHGtNZg86OPVBXa1+6JNQDuz7YmMiVq/GX+IVXI8g
vTpXAkU1HVh0cwa7eojJAmlcHWbDkblNAgtU5xiQ0/ZTuT7LDD7YQLq6MP/uwHDJ
kWoOuTuVcuYV0ZeXsmYGiIiXG2Q/DhZldQGx8/BTvIiHecy/68XIjZR9T9IixyvY
NpCv9K14exsb8D5gmg1oBhwTqsYoLn7m6wuPa6lO4ZSN61hJYFYHAlJHqrey0PBi
NnJnPQw46wi8t2uVt/lKxDMvMLk2BaTusBBfsfO7O27o5niwzcPuGyhfYmod8V0M
ECWDytfNFBHVzWeG5WEv40YBqnmLlpDU5C4uCQvxuafKUF5of7uiQRlrUt2SwPEw
g7p5Y1yqtt0onjxcRuCMSsmndC3eJ5Tke6ZV3j2ZNKGtJesXDY3OCN4BM+EFVTLO
2Bwc6cC126CGwMaoYJMXNaaaD93IGOZ8NlBe/EnnXUCEL+Z42yPqXk37WJdEXgfj
syWRHcGcJw5yMT3EkzSaoXJTNwMLzsj2rMKzOa5eGYd0eAmRuDx+7Iyhnc9ukZNp
GNxqynOj0Nh6y8kVEGE55PF2vcX7/pcgAN0+OAB7Ye5nulqwT3x8fxxjXI9Ckuew
ZJi7jHODYPNdt/J0GbEJ24GzbHya/7A3+wtipnIPjN5lzvvHVoAGbqzvXMBjk/K9
2pJrko5kk+uQb2+ELTXcL//vilfdH38gJ9Pw6vHTnYES2M8M2gtlQEtb9KXdV/7D
JiuAdhXGkUTvxVD/sgeA5uI7E7Vhj6dON2JKAp6gaiGtyLjSGZuaC6hS4MUGR6Bx
X1VGVEJAEAr1rmIfFadIZm0Ces7BsGBz25pBgsxMUoUP5Tddrk2lhqM5F1pLN/DA
RuDJ2WKcFR7ZPPMZ9/udUDtq80Bj94AYxhr09EgXW+bMTkovO/KNqordXgl+VYmR
KqNIj7qEQ/Q9tvgD4uOAKD6qMJfaXWIc3kuC9IXUmBakKRpGmtgeZpnMEQGLgeM2
SGf0Dp2IDsn+yCESJkBXoyq5DdQgob0FPXIzNBUUiKQxHMOGm/rA66Uc6vtAuhjA
qrNg6Jkh0PEEy9jFHwxX9cb39ND7/K1jjtZNdGT0ieqJNw+OX8ykhn3kWgkYPN9I
pN4Rootfn/iH8XIIUa9Pd3kkoOj43okcuY3CWzrAd8CkVx5rRg0dJUXrYCzNCcyO
WZoDxVRJtSm26HvNOdvypz2J1079DhXv2zFiGxuwmucMYjqlyx2At5Qm3BIb7GMY
aYQ8+daIx0XgiVIUcQRt7sW5DbK0C8VEJIpuyoutQoD15LxaD+w8JGOnfkr0JXBX
Wuh4Y4YCvOS0WktMyikoyD6RBDTxoB7d1dOnrCXAzAdEsrYSLWttyZYLWy+ib+GV
cCHfEVLotTIxsRpawbMx5m22SxBea9Hz9w1aRb/Y59gGlhif+Lb2Faok4bpAErzC
oatnxg2zI9erMHGtR/E42Bclhr7+Ba0NZVlMXOKSRbroUEdHYqkf/5guFXngGo6R
EQQC7VSgpv7KJYHLTT7gBho05c3kO9mrvcpSd3YQdQSsU0bJXcsGJV6/65LeUUfd
gvCGlLEaEede0r6Qgt60+xXwQ6x7lhJXorBCQ4/VqDZArmZqEmHugc1Cf226XRAb
30USOZLReN+J6iWgO48Ku0lcXBSbELhexcENvIgHlumd7cAdum5RGmNqkANrd9fc
8ilOYiH6FMrYPwvClCqnj4zDFMvovRkUK7MmO1muxZZDy+wIaauFyaEjF4o1tg8x
fOZUbefU6iifEjg05jFsjlsyxbhUIjZzcFS0khXlPNTu8QT4h+i1gcKrD7oLhrxb
9IG/YHxFK8DUca3szNz6FBEyvL/7egT5IEYeYKGbWrAGes9hG0uhHYoQlIswbaR5
azoWe4cwF9hPjzWZUV4Rt53ofben8SrRnkjNam5fZrqsJhxNs4Mr9+Qrsfz2xERW
9QjKLebFTBCcJvzNhoviQ5TQl1c6Rl+SOxppejSYAa3Beqq+CW+YlBXgQIfdq1gT
BP1IIswywKWzmGbfOq+LElyaR05B667Z2TKC8ZNSVsaImIRohJv0GV5oPmINhlZZ
Cgvd0LHztfYnxi2zG4pFyRdaCm8al801GHu7tS+czkcvhgNrtQL7KnsKtm7A+srh
r2ox8eltwA/98tBdH1E5j5oDByL52nIiQ2n7nD/Kp+bi0O5RmbWcCXwkJIYDh6BX
yt8nKpdqe6dAkpduxkTPxTx2nt2sE3loM8PDfXoN0pkq6ruot2u1rEeoU2hlL/z6
96KE6/RgieyW+ucQu5nP7egFeiWINgMHvlSWbv+P4/T7WkWQeP+iZujSfVOrxPhS
mykcoY15pdLzboXhg0EIKCBy+y3jvhS0jqEmwufkFeIg6caLPQta8vC2mCFctd+5
OgcuUMKzBGDYPEo/gJ4i5c3uEKbeclGYYvyTNzqL9JGMygUNk2eNUhZZTN3Uq3Pf
i27zAxndzXvfisJgbzHvWbkVEpSeKrnZYC2ONfsZ2DngewIW+BBNhZDB1QWfx7W4
lcYMqhqRku4JgvEcLBYQsMxY7CLrqGYvdwafv7fLZ3Xv/FjUUL/A3PBs7VoQkfV+
Lg2xsAy+nJE8anVXjYx7RT4XPrP5UZBprYawyppM2Hf6JGTXWPGd+glMPY3o5B/Y
ssV6r8qKZFxsLSNsXuM2+RplpNeej62rqlvNh0M+5GEoFxu1qhqSFRIS1jIWCTJe
H+A44kTmkgFC4vOtibqU8y9uTM4XRmaf28f7iafMQM2DZpCeZ+JjYrBU/4GscyWT
eWS1c2LrWdm3GxFp9mdAxJaRJhYL9ybxJEHNO4Xa7FStLMX6VbZljQi0PWihjCrR
SA/OMyeaod2bKyjVkw/wJHGnjyhoeQ3ndcdkx+x15B4D4bYa3F5viReMnK2EeGS0
ByZHr5J47gE/o5CrFsOMp8gcgLIr8dIcxCU6zf8FGNK/H+9UwXYjp97tLNn6UR7u
mbTn5wSqHIJuy0uHzWbZjFLsboPG+hX2vWeF3+MuxIUM4OquGp7o46rbtAb/NEDw
Pa4KcaLmNxQSAzqbqgEsoFiGHHRuDymmtq0P9tQuCji+cQTzVvJYhoi7dH1x449W
Qbz3qTsopDuYFWa1wNzAECAR7QWfgEy3+XHgvYEQ8g9pv5Y5aSuoP0lNznbVq26F
Oqgp8TsLt2CTSMA+jGB1tEFeuA0b/MyULePQ0WRpn7pLceCiD9yFmK4XTofBSt4O
qdgNbwGOfpEUTw1dh9Bjk5ZNQvZRJXMKt02av2wzRbc58UpIrkFOIaEqPnD/T9fM
vid/MUKlvi6sXM2SCei37vszI0NW8ghgKldQbYCT3/Z1TCi9WBn6ePqSa3j/rba/
AKRJW+P7szuHzlvovoIedObyHpksVie4cDGsJ/GIx3uDtaRtb3YkDTgr9sJCfqtI
+R0hRVK3JtAQexBCwuCc7TzUNVAP8f7/tKkd4GgM64HHlhKvzKEGPIPZW2xl/0tM
gIgwbSWJ09PJIWf5rrUjMDNurti5k8j6EmOvMG6EBKOS6RpJ2jHOEJVxbMeHbsSf
X6Xgn+AjUsW7XzRKG/getrNC20rPj6nlRxWCnA9goNfxaTXHcqcHePiyW5THjcrV
5vHVuBTbbmE1hZqmy+Vk9o2EXTHOkzDjd27L2Iu0EKB0l5EdJaKtuuVyUYV2TB5e
+rJFxjyxsXErwkOSm3c52uJtQCqgNucGCYgWrfmycrrpMFh1/KlMCTNERplmNglI
qf5cdn3WGWG8yp2q0iivmlhQTMRzHGwzU6GHeej2gB5xb8p0AgZ3KmUWtitaKuj+
PQan7s42T8adqRlxo4Fue60rqpoxGbgvV+eM7lJzEdPP6kZ1xaPbbt3ZAdRtkot4
w++IqXxYgGgeBSxp9zvE7qpXDVALvOBGv9/RMCfSSBYQDbL6SmiSkRx8By9GCytj
sXEq/VRx/a2xX0XnixkmmVFaVO8XBYqcYW72vO8BTtZVi4IaLOV5oihohe4Y4zhU
UrY4V6C+jgFenTUJ/7S4WA9mCMxleQSWDVhi46tixEee4ZYalT9UJTTbuba8JStm
kbrQ5/y9KKAK2CMVlHG0ehwM7TTfDD+M4PAq97ett8HD7wKt20ItvoCqkr3sx1Ib
FADFGevlkAJL2I38stuttlRrhzGVNrZ1JarEy2BJizihZwOejNMknh0VazBqe6Wd
/0bVFBvEWx5i6TmxfNfcWB4JTCB4T7df5zxTh+GuZHwSC3xi+UgNJdqOrNFjYzS1
5spdoYHKQ84KmCTHITtj9uuNGqycH0YtCHx1pzfgoh+cukOSmwPan9ZB5Oe8F89k
8395iEPobSLfjDCjUB/iLzt9SQMWWZKf3cbLUvGxv+ywDOx0CXC0zsIlj5mp/ag/
cQAKfCZs3h+tnyiWzdCz44SOLnnLgYFdUL9v7XybBgeig1ytU+msh6bE/PEIq8TQ
AyAxF5QaA56d8OJVFotZ2W8KMehYeZcKa4yQfZlE0tR4sH+NSnolpLfgWs9RzJEu
aZCM14cbBnf0/BSb6OqYtBlwOSf3v0oJUbvYtjNHs2jud4labRiphlQSUTqCESa6
AxVhqIXpIKnpHq7vdi2okVrp6jPrAQT6WsDNfF87k5Ca9jfMRvtz+/4fCPzBloZa
TCW5P0vnx/gmYvUymq+9rdXicT28uE+f61Ds/uT6OAA/tQwK/EWw4oyKyKqT6F1S
Get24lTXPJAg5N1vXjJ7l4839bMx90g9+R0Ts32BwyZnPwl+va4dpdv4TZWjHRS4
TxPLqDixavwXdyhB/IfVbXWLzkwkcET93TBY8zM8PZHLWKV5Po0biAdpDa2CCukC
RRCkRuIY2iL2WzjJf/i6z2+NfPT+8zVGDQTRsryrnTMg92CcOjf1gnwUOw1dHZBR
0Dn1K4Laous7YaafpnLtUBq7pCNVa34G4cVncSqqmQZnfPP4KG2H5/FKE9LzrzNx
Qhn7sX2SDrlxHa6YVKHYOrLH+OVDhI65gCpEFZ3ORPjFh6tpOUniiS2JXoC9Rvkw
Bj1VYK2hskL6VuKWeoB2xPtVnUsxXrZsur2cVf6s329DZq2Nl1rMvGOD+asYyWUW
DQdpSprlYmJqYSAupUkDhmA54DaS4yubCK+XO5QY8q7mx0wsgHB89CPUtoiAeAYg
c7py3YCCij1kkf6mPGljK70gM6dskLMq48KYMZHMqpPY2RcRKYIVXVkQDVerROd6
6nPPA3ByM4duTgIqEQiu+MNhXsopWymkjLOrPmCgxJH+smuwnBNIc7xPI3ZQ0u/v
NEoX6/WeMJppitflnNE1zGuPcRxqtP+p5D/hucKKjKItANN1r8qhPzzZgajBJJze
CDOb8I/NHH1K20iqgyL+mJo4qTa1Zrj9va0GzA9hfxFem5+kcZ1skXUO9+3i4SH8
l/+rtc8I9VQDkwL37HC2Xb9d1apsoKtxANv5HfsMzVdJjNwvpIKbcKVUZ9+HZ7OS
iIANlj3Iiu73NwHcoGUBo1LCXPzNzoiNcejfdVzTOJ/VpUdqft33oR03G+/LAYNB
UNcCIAAfOpRTjQy80ER09oed9t5J1JEdhy9YdwvZOcySG6XQsaPwto+0kuVe9q4h
i6MpvX5FB+jwCm3eLpqU3yFcBk7MEvRm9v1pyivqzpeTaA9HFGGNLkP0RVAp0QEm
PiZ/LTvhn2XSx94jb+Crrr/9ZxHUwgmyqN4fKRUZBxvijFyllUz5B/k8CioNsB5D
jmMNFHSeE3xnIG0bz5cuor4gfizx1WVDTsTkoysNP5MVjNZqHpMHlie8oYhJQMJp
UQlUgc5beGYDQcJwPSmB7k1XBBcdrdrrYObMh5aQT85YvxdtYNKF1REAdqFurXka
cplFH22hlshZaakeGmGhKDS+Pkke5GRXu8E4/tQ4Gg6JoE+ESusNtScS/g2vD4HD
03viPNqHtEDS1td8mtrhWvKJbduwPrBtknlyaLoLEsdFCyFUwYCn3gz/MGdMHnAX
vaG9znAjBPnXPW0Ip3706e2TdM7k4h8lA2iaGScItjokr7kWAEWHTTS42QWD3DdH
axmOda6PEvQ6w8SjO71HtypcdpMdL15jD7MASwaHT+p9vGWorv6yNfLafdpU/1vj
d4/8ZagHo1LZI+YImJPGDOgp+t/iuFyo+cwIETEsfhsv1X/47lYIWoHFmzvl3TBc
fJ1pdBqIrYCISJBbrMa7MOUfPxHr2sFtX1wHiyIdfn1wg1RH3sesb08z4F/b8Y+i
8EEyWmmNplz6T/cHYzt959D8O2KGO77DYW3QqV/5sda9Pj26c1DTmlp5kE/FrR9z
PMIT8wP2RvPNhkPrYrdjP/KLhx4UKs0wBJbxdGkcrQPOREJfbVqprVzGOFjfjFDB
MV75WQLI1S4ob6vYmcd0cjiEH6qeC4BbwuCoqsNLxn19dbfJg3XkxSEReNQdTezv
mDWaq+P8PlLV1ITZwEKgiWB40tFK5n3jIeXg7h5SQ/oaKByh+W/UXd4ZjhCTzLLG
u1r4zJHscdIE57Oz+dCDkosCoJTECRVIJ64/VplVBrSF3PBV4MtpPWYU7si0O9Pg
qMu/AZ0zHKxZGfN0Vh2YIVOVKkkoE2twL4nhNrHoZx2ALelB5wT5zxGaD/0xwl9P
4zOjEr0MnbNM7nUpMA/crsyUhqVJpS1881/ZyVyDpoM/3MSm6T76JG+acsQC9uOo
BhSM02QgggVTPv+eZWfAz5ZU0Z30Qn3VG14S62XeE1DTokWxVxDIViiHzgfthP6l
wa0JKQSidVBEEyx36v/29yDIJ1tTNZ27Z3o4Tqe/P/ezSHIKrjubze1SrZBXvD8p
HloLOeyPQ3Df982U1Wytw6DnSZlUyb1/PIWFxYldXdtXOu1AWcMBUIR/LTzrybFd
px5t5FvAPCpYEb505uJp7I2m9Xorn+dEvH2Fx9CdemW2uDcrE6QPtFfGYrPjxC6+
BnmZ4PWx6yMU5Ga1MlLPX/quXMvN0B1Nfx7aRlvfM7su6GB8/Pak+olz9tH9bxHh
BxvAtGLl0/0ennWDwb898l1rZB6tpHVZ5lVFi5DICq4L4Ko1Q+k9uhw3GVFCZs1c
Y4sU849FYT/Umx6CuUTP+xyWrEwNmTnQR12GjZJJL6M2KLen+4uMoqUdAfdIhp7O
07cJiXHc0BkyqORoZKpYHQGNjDfYRg4GMHmNf5hpWLDmPx++DE1zt1eX1FQyZEwk
0fApwHfVLOaw8h3AAUyTaPeLai3kOcoMMHjU7+QgjHcyCZf4oAv/QkuK/yrBniZo
5KkPZgT2qSCyOVoTHBQFAmf0U+oSyvMbY4ajo8rnjOE8KJQ0iGhqIQDFWlRJHL2z
OWc9z/iqa3pszacSVaFEDw0qDI9YdB8Dj1cx/8fkQhm7+ED+IlCKrtFLYNmC8c1j
1gATb2BzNwT6z/Ji8sxE+zmAyAFrDAD1uIvgp8RuQSESJdFgYwGDuSgq1jy2Z++z
0LKFaE/zP0KS+DW0/v5EXyfzocF1yB68XZCsMZ8U7ACkeSVcoROHmPeylnvUC5rh
IhQsMVoAl1vsPaX4GniE2b/kM3DbMX1mYjtSQMdZUuDPbETRJZ2S0fB6n8ZrZL+p
dflgfm7osE+JZtBZ9pQFRosQTMlIgk7xVwxJktk9rixWMIq/A5p8+xAqdPjBGqmn
qvj95Oau57SPXDpuMEDDJMgY6NOLRx6zhLRYq8gkwSlMtb1xO02UaYnGUrXzcSvE
DY7nlPDHEE2m4N9fetisXBmJLuqbj7hHJI4Y1IB9aAnDKgk7AZ00T/bft7uh1oH9
3Xs0TXd5lzQG4ikPjMAqUp4DO+/IYota/uoRZx6ES0FMvrLXmLdCxr7RJw87DuYK
0A5P8WWFNbaxVzkCM1zNhM3IuiAO5yb4A0cGB+8wSEjEFX9X92OB3VRvBjo0jcWF
CkuIegL8Ao19Hv1fH6bEYJHz50p6Zb31ygoUGuznS8lSvQhcCJ12c/FCEA1Ij5+S
vek4GUAQewMKFtUUtvwYlC88IY2Y9owasG/4fdWYkwR28XgLmEL1i6vnToHwQOEg
EpEtKEEgLRIUMxGfDXT4UFFKX1HQJH2Ok8uJBXo/DnqQiheaWkB6WBLkruzaiLdi
AdS+be+oujWerAW2t/j3nB0DXG1D1SvPBJBbTJhQW9v4nyHokgd0htdSRovtPaVz
Vaq6yN7Nw2k9T+o1eTEqEch8QU0627gHa6VjED+zPmybLtxk9v+88JgM0NjJEdo9
EXyYJk97irslvPCiDLzoDRAxwWXBhv7plFPagNpEx6VmfGEFvh2KV6OIF7VoV+g8
9jgCPmdt9RkEPx+2R/g7YcpxCEOpxIlYyALDb5ZZLWtifbfGICyFLSGx7Swcdei5
FZD01kD42aVbeqFWUvMWy45G8ONGeDT+E5MXayOnX9MZv096xnJ1kR8lREt5XfMp
4s6v+03ZsrNPbxFbFry4rrnt9od0lnwigR298jD/PCWRTCylBpze3AvujJytlQxz
RKX0Qwd6bUGkd9qhcf8Nf95vqRYSMGJWFT4L7Vx+5vyYird0HZlnaxHMaKL9BDWh
n9W7dNhCtE2XtdyqVqzSszvLamTXE1SwZ4wV93AayXs12htK4nDOtxFclifGt9Ju
mCrZzY1H/2dN/RloHjx8PDwggOZCtZjAmozkESKYOmvIapyZ33bFal6RGxaXzR0B
ZRdjruJ5/NQJlZ9hK6w6R5dI0lu71N6q+hoi3PmlFf4oxDDi/Rnzm7DlaaWscAoW
ll038QQvEdyCgdVVSlz5zUY5E8TVHMyWYK5/caD78+8xp3ZhGcich+eJtyO/TT2d
aMMtJ2/yJZ+GYp14dKySFuEhSy1INoBFNh9ofJ0IzJ3ltjf5XcvHQ0VGPj+TAPNQ
Hpkzd4kfy8+/6nrb/0eh3/BHyj0lwQjFKlEfc/2Wvdu+Cx92NfO+BknApK8p5+FE
3emOlYbYXEQR5gCzuKPXX5b3RIJnwBHQODXjXlkIqI0sPOd+ekxqtQPpQNUrS/Ia
PWuhp0obysbmp0W6+5Uk3+dCRp5qIz8X4IpyBw2Qfr2mDlZkiwxlgWFK0+l+P+SV
/DxnFqtr/4ADgRy8OPvE48C2ml6CKCq2kaCAdkkRqb7+yhOaJZYdEwW1p3LCD4Bq
ykp6XVHzHrChx0tZT1ZpXTtF9yT/ZQ1AsVgesDfK3scwwLT6SHB+q86x7gNKzXg6
/JOLx742w777CKUSEhpgqie/C1BUgqOtZPzsGCbPAITVTo6iIg5Vszm1vk1T9WJa
+FDAygrc6gU6ZojYb1mQxNCMpOG9chujrOGA7vcDYEJc5I9VysOyWnZevUiqnA4B
nsashx2HFtVujLLSVZhnI+R/Kwb2yxGoJymp7W8f3ODlco73Op0c97dP0ZSesSxy
5AwVanjoNYBiPJj4HTaqmDoUeHTZoeJ/h0Q8nR5n1QWhQEvrxfRBuwNL6tXv8NYQ
CGi4LjQmSzOHdjPCI5FMru6jA+XmHQu1bmsnku3BjOxfns3Z+gS1AhVmMTVR7k7+
DhDxVA79E65oXYV+/0exj3Q82k40lBY275V6SCZQa4DG7WtoE9lebIvBGe7YJtnM
wIZHGi/hLRAWBLAAokBL0ZRB7SHNtU9779FXzP1V87zyuNe5F4wW1yzFwk6ZXM3C
gkDoQdYtL3iuopnhSqkSxTKqXtpp3oBd33GzzTiod9HpzsTHOZM0mtRAZ1STF/ng
A8NGL2BtKQNM4nchUnUtbrKYR8PWkbG3zt3W7GBP2mxTvWOGaowB5DG/Y4KHRDH4
RwkQsNbLulTX29VmqsY/9j+FYC/RO4WR044jILN6RMS1/+nnrJu1C+6B+prGsc6G
pJufX6LP6sE9W3xFRlWGpc/dV5C24xQqwW3HpKY66NMD/CKFyv68sI6km1QU90pF
Ud0eQ1/upH9giH8LLkOPd1i/5TESEPOsPjvDO2llXVtsZb8L80q5ZCg0MACRrscj
G2uJ4rQJOL3L+vgwrploihgGespGDeqfZD5pPpFxlmtmBRi4a5ieZ+C5PdAC4ZIF
gbtigwnLLJ6ct+zmFtNDq54rlbNj2648QCkEqurMfXlxP/eqvdZwmFoHprB8lanI
Fz5/ZiYMSs04rFPuZ42DdWWKiE2FXy9c0LEHi2OLlwWkroizU31v6a9aK0/tJMLt
M7smfChNUcg9EoT7mZAOBboYOaNSRhxFpTSf/U05DBW1EZW3Ba4C9gaKRgXMd8/Q
OuU8OfCNL80aE9vc5XNTgu5vjyMSbCjXaDR2658eZ1r5hnuDHEtEE5wBoLTv/xcj
maOQx5frrE/NMIcTCRJatGsiInuabtHRMiM8Z4AFCuGuwgMxHdbesj7d0HdSYP5+
RrlhWfQRQBzIB+j/cuerb3UM1/E8jy+uqHN/sRcy7kEUVtD9VvgKYksIXQknhPUI
tr7MojCsCDkmDnLZ8hikU6znyhxAZ26huSgpQl4Hqo5f84YSyMwFiB2LWw7K6Q6v
mVCZLYcfN6uwGI8d+oVKMl+7MPzw1Ro3Uj/eS/AKx8xsBEXU0Uma9NHWFTWAitv5
fkaRjMHaT4mEZYU5Am7y+keSjPXIB1kZLDK+E+nLMssXRpm7Jg/vAbYKd+Ps+1Ot
ntb1u5vYBqzq92BXQxqRhBO3/NjigJpSqG+dRfi5TFNVFE8rIS/e0jHIsfJgAPy2
K8YyJKIqhEOFlnxWj5TdsSagcGlG7+MNbQHFLkqu2Kp4hHPxYw8Wc/BNiistgye2
k9n/raLarVqXXaE35PfRMu8u9S2Nx3npMSNEWVUyRAGpyY+kS/61NY3j6VrZwKnB
9XA40F9V5BvECT4lZYPOkzrvl4I8GstPA74wcpUhjzxy0ZEWJb7Zl6Eu/O8Ode5d
LjYDztm+mK1MqVyTzJorX25CR7zlqNTSQ6m+EttsUs8rDc7tFY+TKUS+RoemoCyC
IeyMQ30MjFsM+XFJM1ettg7++a0eS2x0b6xZSoKQKK53OZC/Ps89FpUmo2B1SZgo
w08Nnn+tplWoZ1vGPlaAGTL9ERwU+rmdzVdrgP7DGYSt25SYhL+z6Pa3XTxecTbQ
FyRqua/Diz1PIv3t4ri0Sf3Fr8vRENes4g84Pd27hOR0475UkW7NSAEPQhConDDF
YxKL596QnCGb6P/TeCcHJWUjToaeLoinhbjHcc1LVBEytJqricl9GFPCJ48xHSfX
Dluay++8ELC9iMoSFKE/w/nxQ45lVQO10Ap/uSiGWJoOhJMDrMbcKUNaGHruHe+Y
sitxJXI5hHpERqu/TEcD8lzPQV+oJe6jkqVgVB28txUerTKlLHBwWNoYPt4P+mDn
VOQFQo7nN0yUl+OcjMvijEjSS/eMZ4/4uWlpAOsVrJp8t/qQiZ4l/tYRWxQIxjez
bKHzwu0Iq1BDPAiEr3rmJUaTkLH3276RvXKiadwtLsgBUM2xsKmKr9amMKw90c93
f3bHaHS9Qiyn71L6XfowqwYO7n8xJXJW86G4Sl8RnKR15AnOzR6TGADmB+L9BQ6z
12yw7s1P4aomeP/nDvsHcioTytbSBxw3F5FAR9t1wQE7qMNl2moJbcD3/xrysgiS
YMMpMukwWdhk+5vQXt/tSYaNoHdRvamReXSH7gSQQLBVvvIaQ70HTsz8KJmdE13g
EQGaL9AihVXfnpO7/y+yxQtP0wHpf85LbPiYzt2mQC8r0ewOo6OZnTBYOPkZGewo
KQ5GfK2ZY3DZp8B8fjrPayaIqnSVqEi1gI27pRwFlzeFcIg3SGorJfdjBkYqMIBM
t8Ke2Atv4cRJKxOijlMPXnXERGpYZPBPaOB+SlIJakf5D/horaEd1L4CTx8Rmv2Z
JdsN8yTLiGTzqP4N6NsBbBPNiHHo/7udq1t2eOoeNA1wkIrWIK26CAMUByREg4lw
fFN5zgJ/1Dmykpgk5lFjtKSScEYXsbfV2ZExRbhox+iAahp+xDpiJXxTfi99/dPJ
B1Pm/4ent4lpK5okJVlo8Q+xu871i2U/AdYIP9DZkV3xAbzacyY6egEHdZ6S3QHP
8ayx4T63H4SSB/8qrICEJut3RU25UGp8ZOIhpM4NEGVs4q9XXJRiz9SXhjoxJLya
tEc6cB3XUfv8sgTYo1a+E5UWiQh/zsFV6YSc5Korpt5QRmpAtcch85TAYPxnwrJP
oa91IolbrzKFMMEGxDMH9kPDk+806QLnQcMoIS8+vsBwUzjuzW5nPAPnJZjBWB8J
ba8Cisgmfhf9LWoCFmcmontEjaDvNEhYpx8qoTbxrqsXxvqsdrYWFTJ3Vkl3AmSZ
vetODXfm5jUWV4hbgNKdt2L5RdgRKoAgc0TTX2Av8LUDkdfbe8PxKDHxc89J0yVO
mjFA2zXoYaNmBJ0ZgMnwNVQSOKryUE1FrimvYrn56CXik3FKFxjFbXDow45XirPw
6vGx8ImOUi8rqyyUzC8wL2HYZevVWGNPYNFrq3yJfBabEklXFRU+4h6Qfq4UVaj3
3m0alLWFNc6YvoCsVjNTMhHiq4ICSySK27I3/l3hTe3dE0arS4dAUxeNbJi3rH7H
RtxzpbZFKgrhLC7jW6O6fRLd3lab7mCupYM828R/gSxKbSfdPc+gtYnFuQYunN9o
YBmOSRtVkpEPTTdqKuWoeydCZBijkrb88EphLUeoZA4wPzShuG8feDg1GOQErMeb
RN2ONy6GcOTS0GHo0b3G27Fl/vYzGBhmxlvkzdQ7XpdKPfuWeE2q+N+Bokcr8k1V
O5gb650tX3z6mKuGyIU8Zg3tz/eQmwUF/M7fgVdiTJxx6Eool1KHfGdgFNahwTrO
ON4LOu1FJz79m0aKXnSgf5qJD9CrmhenHsSsOOOZfps4QzHAxw9tfv/3Fb73zGY/
JE+Ofi3LDFZaNaHyQh2Xdh46svFBhFJN7tebaQNnL9uXvHq04+LfvYnaD2x/zuqu
6rgF6915KDAzk4EC+AR1YgTmvgmX9UeiEaUyLtc/hXado0ARE7/EBybdWC3lLm1m
n32VrzLJm0InJ8io5COrOr3w1yhl7j9yQkcP8W4TNxAsyNmR30zKAXUsLd+NcykP
UwRp9ofb5WIFKnS80foTfjhVEtyz0UbmfKvgpgLm+OwSz1wAVnFNPHWTF0POdmr5
mpgdv9yWJgJ0iODsmTGYx2y5x7bclBsD2/bRtZEgHgxVdpzubN0wniBwJm5mtV00
Lorbpkj0ydPUwayqJ/Kt+BSES93pnhkbNKshxHmebrq3eD2RTg8la3uc8lqqfNl7
udmISRnBObXnJhxB5LQ9VWINmU3u6vkrxOXZs9zfkXztT4L7ptabFCjTyKZaz9Pe
flF4iKNjuBl9G7RZNXvjJ0kcQN7nAesF4SI7/qK/6sbVxLb7TRZIb/8ilUQdg97D
VPS1jRTqvrhboSxRZH6toPJIo77SY1qnqRSBu787L4Nso0rSz91gN8JxzH9eChrO
UvkbLrJDS4vqJIaF6sxLPkNBQgUqBmMs/DRGVCb+4dnmjoSHd/uuJ2v3eCGY1l04
pxHAyTD4pxViCPScnULoNT6X0a7bFC4FgsMvQ4PAjN1z/9SyIpWZ/T6aFCqWPT0O
Z3z2hNB7vkl0y3m1w336TrvLja1mHG5JB01EimGc3OTfVilHOiWuP46cpxeMBvit
m27CDI8U5kJuACCOoC7XF4bTpuT/meApkC6l7chhj8oSM4ApTFIFvPvjxINV/+ev
QzV9AxSWB1sGxBDIlcAoHejqTsbnCVmDAMbslwcgvdv9uZFDgooPk9ndlOsiMQCF
ehTKM+ytqmIFUMkis12d33JLGdPulePjOvxCnAtYbUYVtZhr2X6f6AicXWxymMvj
ixIA2BCQskiyUaf2h4RC23TNVr/R+Sai67StyWoxDyQwZB3xRcyOPzY/RCgkfNxa
awJRbBFK52/nrrF27+sZHBF1SUgqufelYFrgSqq6WBkG0M4VX+1aK31HPiwuFyvE
TsqF+vYGHmVeZHDkgwrCCTAdAJCoksJpHzZqvu0WkQ2uZFYgjyyqQF3mcR3rPhZF
HUrf4mMl7U/90z1IIDOFgQwPySN+fHZPfvbEIK/PZbAYFgtQW4qRE7Ufu3HhU6x2
6+/6Mmvsne1FwDDc0yaysLepAceOjZUA9j/Lnw97iCJMsJUz95z76MSimnkMhhbN
9hzewz+mNwyunbWrix1/oMV8MoLcYi5K9eWohK5n+opZIStYX+GQM59JMbKKKtBY
5Yap2Hk75sf2xKG2aSfkEyqBDWRil+qxH04lP/W8bR8v3o8Rhg17kOjQKZFG4+tI
An2CEeZPtTAv+1C/uyCBEhps52CdZXwKlzQ6UQDcmwEuiwQWMCMEMWmq0Bd8+mWo
Iy0ADT4IvuqEx3AWIXrX2I5pabP2vplPh/EzyzdDK8OcGN5EOEgHpq6nD9MgAXX0
IQ77rf+nU+XjJDiENtFrIhUKUsk/qKLhR9OruEucpTeKBLq1tw4OC8fXO90+RNf1
v4c40V8Y5AwD1RaOqRcZQpUhqqH4IweQXEN9qXttk/ktkdZzQs3kb/EQwE4gLr+Q
4aFW/pTjQCTUHob6+22ngssG1rojdxBE1GjcFT0Tzf68ecLJSGKFw+/+LBKvcrx7
joRAo2I/iBZWA7Mh/tyqjDyYx1PUzHsO15alaReGiazkAliJzVaXLoUStdcfC/F5
KpT5ClbfLoLE+5LahPj5nMe2+gNgOLQLbgtLTLU+yonEHMyOYj5+6QigUcMiDHtG
30wO4TFFVvHNbGG2NQDJJ+dxEyWMBl6+TpuTqQNqRT8o+eW4QkD8hBoycf46qWMK
mIuu2eVzCRypZVGPU49gB5mPgwlPAMLGOsbrIYI/FhbZLfPiYj3G+2Xz8xeH2PJP
5dv+d0kwn9HJzjy6Pogv/L+6iPZMSP3eTlhmNk3NuYdUdK6XmmkA5xWSzqi4kiMs
VrhorPbDQSqv4ZFmIHk6MbuoSuSPQ1lKEaQw7VbOIPiagpmBRMbI8ABLROO4oV7y
HgtsSUy8LePtxwmNyX6QEOM+DQrUqB+P/STLev7g572lyAYTlGLDezfyDZeuynsy
R/zSvBNu+8CubUeIEwumhj0D7LKs59w4Zsk0MtnXnWJDTE1ygDiFKozSJA6NLOyh
N38mhejlNiTZX6FbKsqsQVnmhHRdCv7JhrVV+BdHp9eZVd1OuUIk/EhT8ojfe6S+
2w98p7cW2cY58OQUhe7J5VVZUjVACZ9iI4VIwsPCHt7vlU2s1lWR8ugUCrzbMahw
081/oMnn3SwuAmfmjsJ9DFNQ/pchQhGblRhO9Zv9cWtIV58bgFCxq6v7IaPLOssn
KwhJyGKPUHiQeKG98pwq4d72CbiJvbiZH8TqzpHJ6ilUcyAzrf2hqqnTctMYoznp
`pragma protect end_protected
