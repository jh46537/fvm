��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�%��bh���p}Î�C#u4����M�	N,,#
���BuSb]:�w� :�5�(c��w��
,0��)R�S�H�nk=L���N��a����"B1�ImW	k-�?߮�0�=ݝL^P�
�U/�2D�R�?؅�H�������-��C>-?�7�0�+���]0�Ͻ�@� ���e3Mԡ��V���bB�l'�@-6KoMR Z:��hc�F��p ԃLͪP��}a9N��	�/�;���n�PJ�K�X4f)�-�yi���~�i	 s����|�J���/єy�i�c��ڠJJ*��(�u ⣯]��mr1_�gx���qL�*�W�����6��S���� �C΁��OY��/0Y裟�/�z@���"�W�k��2)�ԀJ�U�"C}D�qgv{�gތg\�>}._�>����`E�������#3�"��V�0��O�<m�v.��M����_��ۂk����Cr�o�.�q��3��o�;�����a��h�$u7`�)���ضՕ�a�0}v�H��"ּ��3����D�X�	��gvx��"��w�~�m}��2\�h��:Z
�i�F!-�"*[��	�5����3��z�x�e�T3�,f��T��1���b������]�o�"Ir���R�?�������BD����T��pu�d
C��Vˁ��@�M�32��{qRa�w(����pӢ�o5�M~4N1��x�z�-+Ʃ��3a��x�O-f�3�1Q�P��@�I=��n}��2K��O^���8d1o3�V��j���1���ھ��"�����_O�ˮ9�s�@6+�+i%�j�ʕBf�"��v-ٙۺ�U��#�ѣ�)`������=/|W�Y4��N�ƚ�C��q|�lgr<41�����`�Bڴc3�XJ�6���E#��Q)fF�����n8�	�F_b��|��HE���h"k�=�(��m|(�����az��NX���8�bC��}2��b�h����f��w�3������Q��ֵS�ܷv͑s�����O��F�kXK��:��L�0�qql���ʙv��z� }A���V�
�Ŵc���Q�Z��w>k��\���j��v	��++��YL'5Ӌ�����vi�kq�e5to�x��H�Y߇Ö�&�F� �4@QɎ�3`��gw��Z@��g�>s���ƉW +�.e�'�j{"#y��C����A�"�y�9��٦�	���~k��i��H����/�`V�`�ڿ�B'�DPpC�@�;�5����0Z.�=ׅB$���w�a#B˗n��Ұe��#�|����]���%$��Dƈ?&�K��p�ug��;�к��.{���&�CR\�2��q��v�w=LL��f���u;sA�C���$p��%�R������ƫ�ȩWq)�	x���b��ܼ��}�Yc��b�'5�����^��!
�!οr��'O��QЌ�}�n�����st�*����4�rGJ��%��D �.�I��Qxwvq&?���fU���Vy1����Ku,�1���3�����J�R tBIK��^��#W��*ւAT_����&� \�/��F�i��$��5�\I�S���q�k���q�Au��!\;�kl�����ﭏ+�vW�	�XdV���9�5x�	��S%ꮋ�	m-{I�[����2"K��`!�!��ֈ��h~urf��/ϱ͝M�7��_��⮧��΀~�T����A]OYƷ�x�] ���r��@y��1�먕T"e�.�X�F%���We[���v1w�����>�";=�z���&>��ܧ�-�k��1ʣ��|��5H���]XC�Ԥ}e}v,bU�C��ӷ�3g! V��(Nɼ��¦wb���qPH��G�HK�y�3-�pU�e�{���|�#�m�2	-%ϟK[��RS]Q�Q��Za���0��yX<Μ�#�*��Y1�c�!S|��c���p��j��AN4�u��ڵ.5���Ck�r3q��f#Yx���<J��@bEP�&$�D9�E-(f�� b_yN�U��}��:�je�OE�J!({,'�!���_!��g'�5�W�@�� E�lY�&�b�L��� "�w�~��y�h97ԓ�ݾ��=�& ;��]#Lƕp��c{��f�wTt'�G�[x=p�����GB���M��t�e�=<��xd��7�H�.� ,��`QE�Ç�.�S�9��N���,��C�NZ|It)��hn�Ɔ�iD��܈��,��`�_X�M�ᶝ-Eሟ�;O�7Vң��(3r*��k	�[��p������xz�uLq�v�{8g( �Cm@Tk�5��������O�$�ޤ�6ѱ�Mo�O�6���!�:��������PRZ��r$���ּ��4�J������l����
B��;v�/l]`}���Vܝ�+�.�8�揲ʘ0z��h��1��z�-��N�?�"���l�z*����x� ]iR���T��r�ٜ<	0j�%�m��I�A1J��f^�*j��&�)�t7��r$�o<%X"iW������0�g��cP؏��ܱ��Dn����| �46����6��ܐb]&8kB�4�+��N�W5F§6�K�j�c0�UnII'T�2ɖKp��<��ȮX�;C:� �r<����ԛ��|�e�4�ҕ�ޔ��@��V���9^5��<~�=�����c���Y�[W�L��w�5�p��s���p1�=���	A����QKNb�/͋�>y^�*�'���%���x~1[�7����4T9C--M�k\�}�qfsf�]���HW�LRlp�U��#-��I��d����J>��}b�X�����-/�&% �+�s�_�[P �*��&���Ġw���K�1K3�㓠d�g����1H��b_��[Wĕ+�@{\u�F�/dq��48�r���C���6�"�kl��e�-y|x?~�̏K�<����&�������0��Y��h	�`���q�>��e��[eʚ|��G�@g�1*n�KB{}]����(#O���������n+�7gT",h�QSQv��q'#���N������������h0�RA$�Q0�)�!?{+oj{���.&��|��՛����d2G���i��ߛ=�GA<�?����%����C�ݱ˾oյ�V�舗�=���ڝ{�����̉*55`Enh~ <a~��QR1S�v��p��i�=�6���K�lӑ~8rI��,Cb(�o����A"���W��Lh��'���g~��n��{D��P	�:���s��w�7<xQ���-�W��?y��������v':f��歂���8��+��<7,�� w���06��U+�mp7�F���-Ջ�E���[�� �:���k����'9�?���؀��-�`%���Qt)����)S~*b�z�s�>��(@?ܶ��]	4�G�O�jG�i��	�a5`�"!�{��S�1�2',��p�,�/i%���EF�'��r�>NI���8`���4����.A(���x�� Q<��ޒK#���C��M��>��*
��ɿ�/�q&���]�e�pv��I�Ə& �4D�F��K���T����d�rd�P��ۢ+�;{g�O2���0O��iZ����Z�P�LX}�H=��i�Ob�,Z�#�\�sD��404hWXXĀڢ�����r�Q�HS�JuǠ�n�	�'��%�m�<��`>E|L��&K�/�ݡ���c䅑�"c�[%CP�j��ϊ��h]�������A�D�I���ǘ��M��lj�]�l�(�C+gZ$�l$��!�7��^a��%����;�~���p�r���M?b J��������cR.�#l"J�Ա���M]�(=`C4�*��9�6�}/-7�h�v|�Wĺ�ʝ�r� ��\?
B󦎾%ַ�'�v��fE�0��h��Z|ޖ�`��*��xZ���­fQx�td㞳n�+���¥�&L�&� ��&��,����&E��ޘ}�u|��Ƌ}T�Z����v���`lLC����Vʤ�0R��W�ʽ_z�����S�\7M�܀Ę�(�|L{v�h��\J���Y3G�$����⦫*4wlt��,�M�G�֨/>+֊��y�J��[(��d̚�b�)9C*۪)��d�?�pJ�ɟ߅����C�/�针��<��
Y�%'ՠ`���J���B����y�����v横��R�!�ߺ�Y��MN6>J�\Żpb���tU�P8@�ʋs5G�I�3Bh�|�0��0P؋�"�P����ܣkvz�d����	��[W��r��O���J5PҜ	��c�t�sm�����\���s���;Ɔ�:=9k��5 f���蓑4'�A�������>�,[�M��~�m|�Xq0���5��v�+T+�G%���h��_����i�ȰI�ŔW#��͍�-ҹ�H��}^�fѪ�Y�6��B41��raq��˨B׷��$>���D`�rƴ�<u��`2l]�?��׃"��֬�"r�R�P���	��]2o�ɹ���ZDco� � ΙvQ�q�������&�|Þ1�3�@��T���G� O� be�R����N�(�x��F�9\OO��Qd���>�����*��e��7�*⎲׾j�JF��LQN�|3��NQ�����+ ����Z���fL#�S~����&"� ��"���{A�*m�;�=o�N�2�5Ne�F�LM�~n��k���#c_w|$s��w�gSβ����0r/��U���8�ј�=K��Z�P�{⦨�-�ܘ��3����[]��y>��`�[v�	t��ϟtRtlN2�a�������`�"Rq�C7j
\֙g��L^s�OK,�9F��h���^n |�l9��Z>��s�-�qe:�ڒ�#�k[K�W�0�J�K�1�{�+�W'9��0�v��Saw�d�DWȪ�^˺�f�F^e��@l���2�O�Ql�!g����G$=��Q��z�>9���n{�����d؜���_��
#:���-t4'0���H3`�/���k�,�3�h�jr�e�2��Y"mF ��T��Ĝ���(�-E6y1-(�Tm����YX%V.�{�b^ֿ�wZ<�fk��T!U�}�K��!K�e�?0$P�M��\mp/�N��%�2���w�_��.AEh�d���y�5e/�,`H&��"�t<$]��w��G�&�g9��he<F&��g�]7}�.�����c�rx7��:�/��Ϝ	~��L�����[�;i�NW���'!`9�,ԣ9=������#�!�tR��~�-�����<6��s�o3�/?9����A_~����R��IG�C�[����[�tx��	�~iR6�L�eq��5����e��Ŭ��J
?<)�~"��n�X�ل�c��Ƿ�8\���x��(f��{t��UE�&V|�GJ���� 4���[m��]���ER�V�\gQ��aS�����E�bgq8Gs/��걷��yXT�׌���U�؊ѸW�`��k��i��l����N��y7%.�/���D��
���W�q�qL��)��g�aE���\K��<��bJ2h{�R��&k[L�����(��y�!&	-Τה�YxH/�w/�f��}C���$��۞��,A�^:�+4�����Ԗ}t#�%�MS	����ɀ�7"��`�Ɂ�s ��Ed��ݷ��u�w���:�(�-}-)�K�2��C�������.���i�+i�=@F~�nd�TZ=Q��'���nP����sD�۱�N�o],g�*��Ǝ��k�	՝s&��,�]�(_�������9X&(h]��N�ٴ.�L/�1.��i�@��:�ot���C�s�<]	�/+�$�sU(�+Ȁ����s_Lk������O��-��t�����A�ƞ�D�����a*ndj��!W�A��ω	��fG��<�-�Ջ+�d��pt����y�"�����RC:Y�M<�l��u�û�}F!��������b�ڮ��wl��