��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� ��
�˿F!����i�xL���G)35�У0�Y6ɓL7ɶ�4[�Z��K!�Rʶ�������*�r��ug��51��ڬ�v@H�f����yp�1r��^#�����6euo���\��AMR(��=�"�Ms��HY#镐�r�)o1iQ|��]�L��|X�@T`���W!����As�MŊ[�6���%�|Df��2�v=�4����i�9K��Y@�Ի��25}�)vWv���{���"C~[Qt6'�Ftf�h}yҫ��/�c�ʍ����~^5�5���L\1) ��f���S�d�J�W]*B���L����F%���{�`y�UfS7�ms=���&f�sB��Cp]c��G�k6o����ƒ�=>�gI@�g �gWg��-�o�W�5h�ڣ��Σ,B����U�����3!�a��#t<< �
��o��iE�#lPZ���q�A?�]��z;����Pe��P�o��3O��	Dƃ/9v|����$��A��߷V'+����|����&�}KWw�W!ɻԔ��s=�p��Y����}y�v^��P�s�TR��P�m��R�%�a�{��\���^Ҿ��q�Q��9ݞ�.��e5��hti�S�������AnU'�y�Mދ?"��ĚEE����`�f��BQ�<��@�3W�C�O)��.�m+��o����c�T��-��uU��4�.ǒ����%$J{�ô-�KrJ�GU�E@X,����!��Qr�?��:ao��T��P��*�Ʊ��R���o�)��R�b7�2ƹ��]�.��%���󡣒�����c�n&�݃7��D���wy�2y�\�-G!؉��Y�W �_2��ЇLa���/��֭w84�kbm��a/�C������y��_�Y͛�Ç�c
I����(�e��\���L�BS,ح����Ω��Wj�A;�=�\Z#�$W@�|5��ٞ�O�D����sM;�"�@B'�I�$�L�����M�"5�o��ad��s��I�3͠�u�}\��c�ɐ��3F�'��&j��H(�2CiP�p٪��.���NH��C@LI X�ٖ�o��� >���fH�<Blxcr=�p�X���E�����@�3y8�	>�+�UY���p���f{Y�8m�[��+J��q�r��'����<�U"a+�+���y(�N8>z�ɘ#1]����j�ږ�@�5F2&��q�	�U�Z#Bsj�B�p�޴������<���M�J9���=�fP�xz�=� D�Q�V妞�Z�]o�kiin�t�샲=v�5/q�59@�
���5(�������Yo�m�O���� ���pOd�l��w!	�Q2	���ibF�J3#�JZ�z��w�L�,v�/�h$���ц��H0���k#^���U����8�L��l��V�HbG5q�.IK�p�9����ё�$���"���>!86��B�7?J�������h⋻k��W���e�WV��%�t�2VZ5ŗf�r$uq*���-�#-�V(�k�y�K&�my��7~�P��o(zS�QS�����'%e��F�J�|�Ea2��x?�k9>��ԛ�}�.���3��˩ǃ���$ٖ� ��sd�+�����0�.֌�m���O!���<�z�XB�=�CK��Ro/a��n����w7_�1ᷲt��/u����w;���5��V�\<3���h�)"xd�ϙ~�Jq��ə�z�wY�ȇ�,�X3�]���ˀ�͉G��+Lgcx�F��&�s�A���'ҝŒ�-�FZ�4Ί�Y7���'�W��0#�k��Q4�?��ط�ʎ5�^;	y�=(�6d�#6q*� u��씱�����/��w��E���'q����@5�omf'G~\��W�4q�}ۘs��=&�1���(W���7�C�Q���4��Pe>�����|��M��b�O���x��2���{}N#��D��\���k��zP�l`d�~	�_(�b���	�g�=����JM
k�׿bݦ휖<+l78�K��ǓU��`��gY�ҍ�s�ϵ�;�=7p��YTrC�})��3�(�ge��'|<M)�qǍ�(�6���Y��r[V=��)(�3)= �����3���>�OA	r��ΘGz��vX�M�)l�S��P=����H�@��C�=��]t�n)�		�)N�UwUE��/��C;�V!��^,����� �5�1@����Mj�lǁG^�hو6���a�Q��Y�N�ǂ�*�_B�|�sX���a��>��a4���ה	����G*2L)�0|�Eϳ28��0�D����G҄��PDD��ĬhJׅE��VW�VH��4�6�4L$�7�o�Q%d���5W9{�� Z�1��u�r	X�Fn:�+��t��g5�t��+LX�3r�H?�+G`�J���:��<���)���5L�n�-|
����׸#�����`�--���7�	\�����x0U�0���������	x���,�A�]:x���N��A#��nř��!����l�9V�s�d_V�����b�+Ni	]�ej*ܠ�Y����C�����k�*�cf��JfTb���f"�q���T�ۭ�`Xr�y��&+��0�ʖ�(�>�p��=��Я�+u�n�\Yfo��R��c���!�����ʓjW4�~�:����`��f�r`�F-����TҜL���کk]O�\'l|�[�vV �깛��v�+S:98����һ�qBD��\�k�R��=P���b-�VYG"z��ɜ���6b��k�f��*��M�\Ϊ�+�Dy8g
�+�cu���h�M��x�>��N�W�+�&�w���}O"#<��CK��?��K���o��(i%��w�Dv�Ɲ�X��E�"��;�7g�ρ����}��RVI��-�p�<��jz(�y��.K[�8lY�J��ۗ����^�1f Xp�%���"�S��\=�JB������Sx^{il�;;j�+))���2��4j����Z����A^�1W��/ޣ<�ʞf�_I�6�Cx?�xh�@�D��P��Ć�Ų�h�q��6�֋���vg�P+�6vXr��	�G��&�����on�����l��(sf���Y����|� �,�$�]0�ӽ����C-��f滲&�g]gߊa�{�����ʽ@ �R#Iw���� �)��#���[��.�d�[���b55�}M�z�LT�R9�\�q>����z�e�eo���nuVFr5y��'ፙr��]�o��s�P8T���Îpo��u�ύn�D��NX���nP��c6W(8í': +Ԭ��I�N��5� u���6$��18l`Mh�Ȑb<4�D�x�#9D	U`�3UC�U���ܔ��n8���Tm|����(�Zw����4����iU�#ŉ��-'�0Vq��~С{��W����$����1î����n�<�99
7��	}��᭘y
$Ǘ�w�_�d�����X����Y��	;���xL� X��)t�$���@��*{O`����+A�ў�n�z��)<YB+
��d,�J�5i�B'�Nap�Չ0�&P�A�
����Lڵ��U���<�m�S>���܂��V���5��GE�X�E+�$l_=�Rε.���/�R6:��{IJ�w=U��$@OK����ez�耼�Fz��jJ�.����)��v@k0h�?�ymiW�ͪuo��}�	�/����Q�K� �v)r����	��n ��9;�X�j�Ĝ5݃xt��EM�O[^E����+�*P�gtj}D	��@s��D���-�
��Q�W��KW���An���MJ�b����_+1B��NY�� g�am��_��f]�B����ȟr��x������G6ua4�M]$8mhg��(C�Ց��nd