��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��x� �u J䇰`#����������T�jCQ������p&b\��r��q�O@'ɨ)�doi�����L�q�_�U����G�#=��$)
r�ݥ1"G֯9���3�5�4�`�Ɗ��pֻ���<���A���R�J���>?��}Ѯ���KI$�o���U��
��.D���ٻ�ɶ^�u®H�(;�R�*R�ϰ��M��4���E@$��Vpº��d�{��f�J���:�t�bl"l ���))`�ȝ9�0d��5�Ge�U}s��V�G�����I�u⹲���uJZ�ܢM*\�C\/yZ��G�|��l~�k� ؂�[�3
Þ~^x^��C�);�j�}�1�z�zEF5e(����F- � [p^�Bɍ�-��K�9�����a���Y��>��9�3��~IB6޳����Ą��t�0�����hys�h���@Jf��o*� �s[�B�z̸gp�\�ǝ�L��Ǩ��VJ��ˠ$;�=-=>H �o��n|6�z��_�m�L ۓ�Et �J��Y�\G�}�v+��>���n�G�+.,����d ���{9�l�����-äl�n@�U�g��Y��&��Hvō2�+Y�<�.J����i彙��g%co�'6��c�����F�Gd/��.DT�8��*^-eI�+!�$$�vsV#���~1�,t,ew;Ѿ ��Hye|Li1t=��.���h�7"� ����<�0��N�7��9Ė��<Є.K��E"�&m�h���2pyLd��.ف�ŋ_oߦQ��Vh0�	�M��t����m|�q�����5NB��_�]E(�^�r���'�`Vd<� cP��"ȟjs2O`ZD(�SQ� +�*t�+�G/)�I]􆰁��7���J��LӰ>ѿ7�F�� {�B��s���nIƔ�~�FS�Պ�%~�������e��̊4���:T�-�Za�.rU�A5��r+��$c�Ĳӽ�����T������L 0��N�%�7X�&����8�]�ؖ��
��Я]�Q���0'����kڜڜ
hK5%fW��]C��(CH��5ه����Ԓ���rO���ߞ��v��v;!�ȴU�O!\��H߯���~xs*�J;#J@�r��1�'�0�F0Y�}�Qm�ʹ��jQ�9��ݳ��P�vk>"G�}x|�!�k)c�aLE�I�-�O0��2x����B�'G�(�~P�Q*�X��P}>^�)t,X�����I8���%�ژ�ڲNPЉΘ�����5�|{�g�e�V6���i+�_�6���A,���,�89��	b�?�,��D�5���p��?���i���Z9&�k�,�N� ��7r�<��;c���'fBJ��������2��3փ��|���(�����c���pE��}(��\�/U=�ȑ[�KŔ}���c�{.s���UG]������O("$Y ���0'��&C',!~P��?��Y㥒TC匐t0����\	6k��"H�w'�ex@;}9���a�֙ܪ�h�>�(V�I�r����Ŕm���u�?<>.����0�����㻀�T?%��O����ɩ,Ln+���xѨ�����W�"3��/��c����>)Ǳu��s�ZY�a3r����R�З��ef�AJ���I�� �:W�n�	k���t`V#[Crj9�d�*H���-�wX3z��L���(�.æW���{<�������e3ܺ~�
)�9��-�?�����7��o���X7�X��|1aC�óZL@@��|��'��-��Y��04"�т�OԚ.X��V�h�-WUWEvI�>g8�=�&��,	���+ `||�(��V[J�q[��*+�t;\�m��gj���dӐ\(#oEqx5�.E{�d9�x��5Mu���f�X�)�pS�����E��^`rp ��1�9����5&�OJ�~�j�i�Zx��vA%(��>_b��B5�4w%�z�X�#(�k�4��cW�}���[�L���V�cppk���8�3@#����<��h-��'bt��7w0��M0o� ��U���^S�q6/Σ|>����Uqa� t��Y ��oCmf>z�\	G<
�Ȫ)�K�YBj��ry�o"�$[����� B�Z��v~�a�'p<D�rQ��� ѶYf�� "�ac��p|�9t�	��.��R�V�������PA�b����Ի�/Ƞe�)6�P�$$ۥ����KY$5����q�]4�o�}����h�ed�E�����������;<��&�@�?��hP�� �y��) �-,x�Fi��ߜ�r,{��&6�m(K}�'�Έ�7�%	�h[]t�S�ޏ�Ғ��F!���a��K.}�V�5�!�Hr��aX��z���GNo?ۮ���6v�
�؊��8�!Mӄ�4����ݠGZ��O��[7*Y�@ɍS����.�z1�<�V�>W�>lS�]YW
��,;5�9w�,���ɺy��,'�A�p�jl���TR]��U�μD#pK6o����նN�'M7�/�c%������wX��P򲃹�\��'f!/����!����x��[Q��@o��18>#��L��<�,l3]� �gQ �J;Q�\a.�
�c����M�� ��	�W�M�xJX�󞄙�|�]NG`ѝ]��!�DV�����b��Ў\D�6��x��\���Wg�<0��"��X�m	�IrY���3�sO!�/z�и�0�ʡ��!�����Ә/�x��F���w�^hY:+.D��a=�a�){!kwF�w%Xa��n@Q?�Q12k�s0Ph���щ���$��X����ƞC$?BY|C<G=�s�xC6M�^�&7�P[?4~+��
 u� ������f5ZMH0ŔVf���ס�=5�f~�+�嘟��l�6�Q`]�t��
�����4C���4Z{�Ș�[�4(lVV1pR�CLpB�����Sk���uh���p����-z(U��/���W�c�?�W��uJ�b@Ƨ�Q$��v��ލ�D����m�Ń�����Q��m����i��s!y�:�b�M�bn��:��{��ۚ`y���|a9�7��+d����5?0F�/we���C��wo��Z]l�T��O��ؘu:>�~���Ԇ:q�yWW��3���?�V�Ni(�Ռ�X��Ȉ��W�f{k<��Ub`����P������۩TL:R��ԪW-�����M%!�7�V�a�5�K)25�j|"SX�>&�l�//��|,�����D�=�v.��B��:��'Q�ġgԟ�F�#���\������+��X�Wn��=%��Fr��c'F���������rF4W���5-	/\�}�R�[#�?1���#ƙWǽ��G����;WMf�g&�^�	4��s�M*��o	){]+�D��
�|R壿�dqWbbN8��y���3~��R)�����AcL���6/s&,m���)ަ�ur��(]����ڞ��9 ��t0��Z�e��D"d��.]`o���l�^4�ڟN�-${�ϼ��2��G�̩b���'�r��)���_������n�aZ�W�s|FI<���*#��V��d<��\��*Cdz���y,>0�b��҄{�w5���S���O�I�W@\�
�I���4RxRy�oR;yy�,�
z�ͣ���ໂ
��EC*��@L�z�:��
�tԯ�o������lJ�txfȾ���s�:*�W�����W��!���+�Ӫ�2xh��a]zƔU��a��n۪w�92_��/�3�<J������VW�;m�,E+R�qoT �'�pd�$�Ơ���J���]��L�G+���1�H>���"����m��9��.}x��AC��[1&͇'����,�U'jyR>�l�3��O�pxI�C�Me}v�S�������1�� �S����\�)TjQ,�"�&t����|H.����I��ê',�@��~S�j�6��H�~z���o�'��'� 	��a���\�a6&`�:��^�O��I\Ps���m �{`���gH��(����Ck���5TSWx8j��)@���c|IU+Ӡ�d��B/��w�h�U��E����ﷹϠ��N{�&�	��
��W�}�k9�T��l00xАL���jڳ2�?�=��Ϊ{�$d��4�UԪӛ.�y�e'��*2�@�Z�v�i	�W���]�%��2-au�f�9�&8�Z��c�ey5��h���n���0�E9�m�f}� �r'�S���Qa�@����+d���[�ć�qmp�n����/pz~�M+H<p=�V)����0��s�#,؃�:����uV�o����M�8mF�csdk6��:�7`^��1�[�x���$@�~L��"��ݖ'�O�K�ܾ^��Y#r�s�ೞ�n_b��c�(Fh��%=���5Kzh���+Z�gf'+�
�]:���[�j���k6 �_���̰C���v+�VJ?`��=t~"� k���F�- ��;�kifJ�HN+ar�z�g�&�o$Z��_m�p�xN�LgB�<�x�E���}�+}|�%��W���do�'/��6�
����}��k��j��~�n_���|?�k�ɞ7�N�H���X�z�a�gQ���L�A�j�4#Z{�1\~�Q�ޠNJ3D%
͡��ɒx���k��%ؠ��~7��T�����@V�ٵ�a�W�ކ�y���)���J?���Q΁4��Mjc��r��(̑��|�S�)"۴�51�D:Z�	bt8��*?�`C����L�d�@�.�3��~��$����{_ �:��f���� *�9�Wt��k,�S��L��C֞�ֹQ4����,�����x����^�=�z�y��B<�'�s}��faи��V�_��.T�
��{��v�}t�"�z�h�� �L�C��F��m����;}�.�o�N6���l��o�eIflD�>;��,0{��ƆZsQK��hk�J��,����p8ߗ�����۟wU��R��/ۄ��sV�T�}]��.�doʻ+w�z�i,;��ڈ����t�+�ʘ��s �������C�X����|������RK�s~���8��k�Ϣ�V� %���6\���)=�$l��&<�l�!�q���S27�����J��Jn���dpg��T��7�b{^t�t�[W����<�mv.�i�gG��<G�-٬vuߵ�+<��̵rT ��0R�θ�&�{���u�c��y����[�<z�v���u��
�%�s�������Y�e	���1=g86i��.��u�)�����3$~�O�75R�p�~?�������뵀,k��Zn1��/��_j�e;+3xRn��`��k�!q�"S���D����Л
�wl�>�V������3]~\ʘ�kG�֖�/�������i�<h�.QfI@�<G�3dNЮ3'��v7S�����W���8(�����ٺ+pI�L�A��'�C4ߴ���|�K�F�����S��^�l�͢���wia�t�r"���ٌ�6V�ڀ1�$d��	m���K���#(�}�6��	x��,�����Q�t�ƈ?:p�k�-V)w}2�����Vt�z_a蒡���km��5�s݋9��'�1?b��j�YC]1`˞��>�:�:|��2R�:~;��s5��2MB=q�,k��*Y��z(�|A��������p��M]��T����zXV�l�}�y�����+av�ea5�P�i��\s*������	c�M�s�/��X���Fw�.����{���]]Ut4���nz;���S#���`r~3硾]#u��1��c+�t���n1�����&&��>.孔T��#��q���t.V֜��GA�<R��:�e��]|���@��3�8�+���v�!J0��1�[K�	k2�ش�elk�_��G}c1�۩�Є��0�v>'�t�@��y�2MX��)L���,Cp^�;�I�r�#������Zs���$����q̟�rI�9�!����7J��ک�����2M�n�/�2)�,+{?���O�G�6��m�G�,U_��4h�>�a*Bd��uH��6�U��s�=$�ܮ�Vw�h�bla����+;�*�cݠ��i�K����na�u>�U���?K�qq����o�k���e^�w!T1o+Z6R"
��{�}.��ڟ��xP�G��z�ӷ7&�.DL��3�{"i��?fa#� �����֕]�r�kО�G���X���;i���F��@g����5��� (��_�w�u@��'��E�8����*�ȧ�3�4�V�(J�X�]�U�"��r�W�%Խ��bz�=�b:z����0�<��.�(�K�ѩ>����G��ƏƖ�R���65e���t]ThUA�\ں*u�iG�G���f� �b7X$�J���)��� ��F�b�K�-\��>�{I��W0�\���	@56��ť5p�.ܝq�Ϯ�����X��6����°�úJ5Up��Ï�T@N�=M/��#=";m�������j[5�2X
L¾q:§�BV�#�2 �D��{����l܌����P�fQ��@������ڰ]�;`����UdS�ا�S��	��@=}������,;��� �"�ܓzA�j3$=�xPb���	�:&ճ��sv��?�!�t��Ԩ������ϣ��E�^K1�΄}�b�I�M��1.����#.�y��&� 113��0��!��QB�y�dL�s�@� R�1�Hs�4�"N��t_{ߋ�׭D�6;
	3�'x�}n�}�F$�₎�ߧ��a�^�<���j�M�\��^�����a�j{�Q�"��O�q�\��B����h�ƅ�ԗ%BF/L*"�^��6ˢ����r�6I���|�\�L�L�i�-jԗM�.]#�FX����T0�f	"����\�����D�/̜�Xk䃗��{߽棄Y͝�NBn.���.�W|�gs�@����P��4�0#?�0�V����������2���(���g���D�#/m��lk�>�+&Z�4���U�����q�>٨~��=I�o^�73ԋ�}�f#�+k���򳏮�U�ye���J��C��������B(`��̗���y�>�&*��,���G
 I�~���)�.I�C9!��C��7�&�'���J�K@��l�2�ե���4gi���������Fcؽ�L-VD��"�;����Y=�Ցf��ntL��p:�w5���s(��Ɇ8���c�:.����O|'gRŃ��`5��G2����0G'P���?�ź�bAW'�կ���fd�&��`��ۯM�Vt��g%��x���/���E�c*pV0�W�G*���_pD�azleY

�4�U�Si��k�S����Ӹ1E�x_����B����Þ|���Ea槚���	4�����)�"Bz�k;싧�hz��[Z�A�����I(�ߵ�R��x·)���|)Q�:z�Ж�5z�� ��CMv��������z���������K�F:*�t6� �lw12n�W���y.��0� �2BIu<�iNu��؁���3e��M�ӨW\�]�3B���dG�8M�d#-_8��s��c��rlmJf��rB|8��HDĬ�c�X�/�Ϋ,��Gi�2wI�Òų��©�pu���&��Dv�,����E6��/ŕ���FY]��X�m� �MȠ?��H�?�������O���V.)/	�H���_1��B��a�	���@M�jZz~P�ث��#�q#��8xI�c�/fq����um�H�<���ޠ^�sOʓ����H�������B��$�����Z6C���9����Op��!i�Ƈ`����[��m��O;s�;t}�ISz5C��e�W�n���EGy�\�9PP�?g}��h?Ք���a5�vG��$�9��N�x�ֲO������ޏ{,$�2h/\ļG%ƭ��d��hr�N\��h+���U�����;������̴���4?��NGǨr��a��w�[���O��yH��z�Pa��a;|�^i�w�B���-pre"v����%����Z1��5ϟ૛S0���֗�������ӂ][�g������/BE��#�xO�=LO�Cd��ꮕ�U�n�,�)sW��4C~#��4�Uq
�D��}*�0�r>��?�H��E�
P4n���r��x#V�܉�6�'���LP��D�}�c�������\got�M{�o����>݊�.V١��U��@	ם�/
X���sA��n�;�8��`�XH��&h�ߟ��'c�2��kz4����8�T�yQhs�zI.Z�FXW�@�89�	��M$ψV�J���C��j����UX��,FK
�sF��^�4!شkA�o8���Y�n��e<�HҦa,gm�$�H�屮jg��)�*�B��	D�`DPo�K��F�ft�;/+9?��ϭ]EOK����R>ɹ�P�襣?;�N�vS�2U`�
n���F�\�%瀬�n�q�|�\�ﳹ�K^��
6� �ٝ���_��Y���n����5����v@Ix5l4se��C�QtR)��8�Dt�v�V�m�Vɒz���K��?.!�Q8%�7zD�n�����6�H�r���o�?B���cf���YH8�v�\ǲ�>��������܄x�ǡ�
��;�r��d;!���rP�RD�˵���WR9|ߣ�W��K��ub˼�%��P~��5"}�H��=�k����8~v��yC�2F߻��|D�M�
|�ʚe��f�u�|��"7�F�.ak�RH�5񼬺pL`3�v�gx�z2�������>&;kpH�3�뤧d��3�����.���>!��)I�=�'N5s�u�?o�u�"`M��+���\��Ti�V�+�k�G{|���|��3���K�����hsch�D$F[�w�d@hV	�"�_�@T�)��E�U6�-�e �����r嫩S�m҈���j�8��d3�O㲋jp�X���9��T"Sh��x��y���0�oCZ�
Ϣ����c��P�6�l��gRQ,OU�����������}��@�i��x̖�,�5*f8x2v��Yƾ��F�z^��`T�cDl���7�>i�4Ry _����[(�Y�]���pB��`ts��k�Kx�q��QS�:���K�}]TB"�sJ���0�_۪?*�-�(ƕ�����/�A��LGOk2U|�h�Q\hs$�w������Δ|����Q��
7U	� ��sp ���ܡ�U�B��Ը퀺,�� ��O��=[��0N�B�P��[q�������"�se�B�N����;mq�5z���"�?a)�o��I��(G�ppy�+��o���|����V�ǔ��ERI�Y+^��V��U�]7�*$��Nz���ey��!����nU�$��y<9���$ސ������Zp$�c�,���4V��)��HL���	�@�����kP��F��m�ݴ$s{Ҫ�f�3e�d#��4TF�̾����j�&w���΀��-|��jix
<W(7Y`���Ά�p�Л�Q�CVD�&��-Jo`y��N���S���6��[�E"��{�x<���%7�֤�yM&��2r/n��e}�~Ġ38:�'����C[���!=F�Z�W
�㵄�l����N����O�Թ���?�����҄�a�y�f�h���Y����9J�_�4M>S�E{TD�k��`�i���Y{i����2xc;P!��r/(�����D���D�?p�[q,����"dE��.���VQ�r��n2�!d��vJ�D�}��sZ?�CI۵P<1��@[�d�N%!ϒ�?e��'���x	�1��N�ypWV�C:J���.�6`W(�)`�:$</m��=���e�h�5F���L��d���hh���\�n��W�s�/a������M����,�u�����MJ������f�B��E,F���ݼ���g�r����S�o)p%m�:w�MX&OX��`@���bO��p�@�Qp�y�V�3[�"Y%9},t�W�[l��]�}�:D��)�G����ѓ�M�l.7L�X����:\�C{k���k+�Üː.�)��LU�_��֒Q��YP�����aϮ�l�z��Ct���/�I3A�w�*OY��2���E���Ʃ��L�נ$�}r\:_0���KG���0}���xA5��:y=��_���B��g���\��� 4����P��ԁ�s�J�G"��
��[þ�t�:i����ͺ1����
*�S3U���ʩfu�_�� �%�I3[܈�|��>\�L�5����?�̈́���'KC�PL��Ͼ$�<d���6wC����_f���5պ�?�IE.��^�6.T5�P���R�5+�dP��i�����%[����DޡҲ:&(��vQ�������@�4�k6k�H00	�[��̳͆=�o��r���ozH;Y�z��)y�{����|H�~�{���g��$�@�d&
<~�Sa�U8
>
;��4
�C�ҫ�pg]MZ5z����>�ߧ��O�A�<�
142b�k5�aE�a�xD����T��p0��c�T�K �9�:P�K�u�ԥ
�o]Nnsߣ� u�۰�Uh��M6��+��bۑ+|A�,�*��9�'yrN��9�m��V�'��`�T�x� ���Y��
���Ct8I�j@'{���jƀ#�K7@�|�NB�^���&�f9�9�������Y��B|���V�M~����/c���j��D!x.X�5	�t8�d����.@+�M]�ݐ�.��ТOO�ER�02�	�/��Ց�zo65�x����Ԇ��F׭�gD��h�����5��C�V*�2J�G�-͍8]���YC�9���;Φ�V,4��!�_w3��"�6v�C��y��U�2L��e�6�i�ٵ�c����R���$\_�0Z۴��|%��pBY%�Q`_5��I"d�&vλɼ�4F�����U��3�#�a���v�o&Y+ı_k!�%���� �������b�Z�}7�QWo_���3ݕ>6Fw���=����k&__9��;g����.#�z%*P�w.�{x���_R�����>˸�V�~�>a�����X�C=s��L�"��Ⱥ�u$�������(�8�Ee!�[�B1_{�-�4��'z�tZ}`!��?����M_�9�d��{��e�q9�,*����yP�g�+
�Z���!�L%}p� dP�̞הن��x�o�L��\EV%HQM�ב��v[qf��>,�h���ɍ���x�U"hë�$�'�0�RJ7JjF��m$?������F ���4��qqz|�S2�b�!�K���~ڂ�u��Ͻ�ĝ�~�	h��#�x��L�=���
��|��c^��,��"8�D�>�m��|�a��*���2�����B����%g,������4����[�fe�Ey/Y)X�&\��;μ~�Ŷ(�|U>�!E��9�&�y�,<�8�0Y�7�/R(�4.O���=a���'!��>Cwk�<���V@�@�FԌ���=����`e���%��_�ݻk���P���r�QNj��ֵ8�2�B�ii��ZGm���{��l�%q`C�<���AƺJM �����/�i��k� 6C} m>����9�Қ@$� �k��?�yɣE���ڂ���]��>�ɿ���=��b��M����f��lc�T;j���� Zi�Hk�r����ay䨔$X���r�����Z�>��u��Su��Q`��>���V��[��I.k�)�-�#��y�����v��iߔI;Ϟp. ɣ?z-��յ�_f=v�����5<�L	|iȧ`�l��) J��+y�9�� n�iv��K���l�T���Ě�?��2荩��\�e/G��`����'�lY�m�J�v��w��YEGbR�2�����=Y����w7{"��g}V��h����r�%�O:�Y�P^~2�n8�J���r�X�c0���, �?��
\L$F̊k��;�b�ޚ�R�X�xߊ����ol�*�m�I��S��b�ӝ,:�G�ca��م�r�Fn��}����OA�*m�*��I-���m��i���>zcE�=��i}��7)�Ѕ:��ko��@��2+mT��~��c�R5P`ֵeM��po��l����/�w��MT_s �C�OI§��ৡ4�6�cF�k"�W�=�9�ţ�����e�"lɺ�+��p�ό�`��v�#E凑}��ܢ�J�_��+P㌘Q��૆����$
8E�߫�qa4v��.�J9����Pb�K���{*­�" �3��)Ur�6��֭wÊ�H�dh�r�l��m�.�kە��5r^)JD�I�k6nY"集�(��u�/��z�i+2H'a�4��	�D��A�Ρ��TQHY�l���z~�j�cԝ�������"�i�}l�Þ_���������*���g^'o�p�e"�ut1�ܭ���T��mY�zڥM-Yi������=/��fc��'�٭���+���.�U����`�;�!��N�r��젞��i��Q:��>�L�֤��g�W��������{��x.�rZ�#�jL�f���b��M��兪����f���Z�h�s����QD���i�c;b��Q����iEVŹ�͋�.XX|(�Yw�h�t(�H� �����]�f(�k��BA��8���9�&�ӣ5��w|�^[M�D���F�=�D����3I��^:
n]=��h,��j����`��"��sBS]�rSc���U���U�]Z�,g��z"�CM@]YIQ�ᜆm�i�j?[����uVٍѨ�Ӫ e��|�@|�ph4�xt��v ���n��"�j{'!CV���uv�ΦQU,&[�M+�e�
� 8��N�
d�J��X�쟷k�ʿՀ�����6~�mu�����B��C�&h�l��緮�F��3�:�ZXr+&�/���q`jS����`��hH�?��OR�|�*�Z�&�T�ǧT�!E�a_|��������舱��r/A`,�:��F��qS�+���hMl�O��(V�z<�FY�9]�k��6/gڮ�������y�i ���x�* +���٤$b?N{&��N��p=�K��Y) xa(�ţ.����z����z$=�����!�N���a�̖�W�` ��7'f�50�(��{t�-+.*?��\�A�,J"͔���h�\(bxFIPO*��%rz��Z�L�ʚ}X��.P6!�OR���@���]������՝�DGݮ������6�MƳf�~�I.t+k�����%��2fg�h����oiv����nSL��ݗu�}x{yE�+F�*T��X�,H�"y�&Pӷ��g2�R��D@����K�!5�h�x����
&��4,<~�ckp�v��lnZ�,R��5m�$�s�����zof8����@S�G�)�}���j�U�7�둇/*���7.�
)0���_������x,���g,i���B{�-e�ڡ�B���_�@���@$�o�@�%�BEr(h�S�{�A*h��U*�K]��v��!�@�2K�g�5(i[�֑vc
ˢ2f�/������Aԧ����_n� �$�c&��K qs�L��������d�e{�/V��eq�ai�4�)d!>D����1dM�"���A}�_[J�:?�#x"ِs����`-�{\N"!���|�T4��_Rf?J�����Q�"4��~��3!�2��h@x��"����Y\����a��䢺����Z<L�N��	H��۔3�-��*��jCw_���M���N�裲�yY�s���D`�/����I�±n_� �q��O�9˙�!+_������r��[�
#>���W0�a�2��f�}=i������˫z��W��E���sMa���6
��P�kW��%7Pk��eO���L����gm���le����^ �q��<��F�r�:���Z"j۴�<��Q�
MhWW��.R��t�-=!є��c-*O!q�D$#a�����+jǈ9!B�tC}c���I���=���G׎B����{R�'{�h��HE�;ʗau2���Wk�*Z��ƒ�;�F�T�\��@it,2�M�����D	x*Ϗ���`9�j�ӝ�Rࠣ��K�dJά�G��L>�>hw�;T�*l))���!-�7��^��e�� 5�bP$셒�dq�GGP73��4[$S�����>vHW��a�2����0�����^[��ˮ�L ���5r��PŜj'u���X?�ڇ�A�P����<��w�g��9��5�^�&��GlL��]:]�В���AQ�K��̯>���tI���_��T��h�y� �Γ8�ߤ�0�pU���yz|Pcr?�D�u�;q�v��D��،J�{��ۍBӧ��E7�����z^��N��-�@(N�R��0v{&'w�t�J�T�Z�jZ��_��<Q�!��9��ą�e���5��!�f��XH�4RX$8��40��ڽbz�%�]�I|�7Gd3�X��=���G�f�0i�M��*��.Kâ*$�Vk�d�KG�[��(�Ԯ�}W����R�Ǟa�7@�*��7���*������B����q��:�D' $?��r�-ɥ��t��YcD�uCM�|�D}d(=K�u�Z�%��!>�o����j�8[K>�{ڪ_�RO�:cĔs�F*Z��z�-��3��8Rn\����~�5!������%�;G^ ������<��I��xsCW��ːg�x*�TZ���;��d�C�p��5���upӜ4�\����0e͸�$��J�-�b��E.Vws�	���4��U��bqzג3�}[C�)Mڸ��?�\&@f��&|�ա��8����[���s��?G��O��A6�}�D�̑�rq�a��^5ᨿ:�'d�>Kdd4���S+�&!��*W�1�n���!�[����>�mʨ�u�6=��N[ٵ0��2�^��=����~�;��<��M�8��W�/�f45 ���S��"�%�w�C�W+$q>��3	�l2mh�ʥ��C�M�6U��;!�Q��g,�R�����c.����ݎdK9��_��HW��gg�D/���B�AN2� ���.}#\$���ГW�L����ո=��t��iS[1e�̀Q�"+���y*-E�1���� (8emQ��3��7}���g��A.� 9���n��"�ݵғ� �G�S �p����u(=.uv��	�a�*`�L�Dk��W�����ac��k,�f��V�o�@1eocq����'�[�o�"�$��t�n�T��g)�`�V�?�ҕ:;/ =�W��	�vZ��e��|��ӦD���ES��!D���2��i������|!$���{�=��b',F�uߛ��p��)�ISp��J�Z�*هRQ�\t�(؉,2�ܭ�,���R��dE!���;�^{�z��֣�q�7�֖��Ԡ�y|����;�$�'0�f/c�����d (�B�"�əG���7��l������a�:�d���N�Q�ÙH���Ô9��j��TD{+O��h�I�k��]�·�W��ƽZ�)�|����|���~򳇶!8���I,�!�Iс-�/]LK�6�M!I��o\Lc��Q��6�V�q2x6��P2���J�7�F�_�H���K�� M/5L���f;*��oa��Ԟݚ<���암�)��%��1 � W��'r���T��&E�@���aqTeq'#���YHl�g+vQ'u#�^��d�<Bʛ�I���6�}������WZ��z���O~Mv�"'�]�.(�6�;@U�xܬ,���y�3��WC�5�ds�SO:J�{I+u^�Tf��'���p���Sm��2J�/��xhD$ ��_��(@_[i�ba�k�����o��-N�<��ON�߷t����^�c@2 3ڷ�.�.����!�=�p�aj�
��zә�� �� �D
.�z	����6��<:8��!��j�k�ɝ*�2��H��aN�6�5�96�"=JT�� �1�.p}�6 D5�=�Tg0*�m�AD&��k�����,n�i��S�ĥ�E�.���V��@=��3�Lˎ �����bhΡ���U4)���S+#etE3��F���O�{�K���:ߖA�	�x�J��pg������+	�F#��U/^��)�G]Y�Gio���U������.(j��sTa�J�����Q�BT9QL!�"Vm�EO*E�|���k���[�]�H4<Z���,�q(��M��vo�{�W����O푅;�Q��#�M��(XxbE��j}�Z�](Z�FeRٲL~K*Q�g�ėR���o0�iK[W{�%�ɧ�۲a�b_��C�Q�
�8��U�6�^�ƒ=�=�a�MQoU�		Ns5�ؓ��z�SH1�
�8=��N�D�`�����l8L�>7��r��{I]xF�klر�44����7��ES��r�p�(=_BE��|i�[M=��Ml(-b�c�m�NףZF�~���N ڿ�A\��C���������E(Ҫ(��2��u�ϒ�U�0#q�i���7ڮ���i�`L���'~�Z� [1���B�^<@�p|R��\�Hm2Z O�,���au4��70�7���EO������1��6��B�T��;>65�b��ƅ�U91�6i?��R� >������s�ql44��2	��R����JfC���:�i_�G=��*��W�c�b����Ui�t�ݠ̋��!U)���I#6Ot��/Zo�'�
p��d�)��'p@�q�z0fp���y�K���I�݆)���z�ꪜ�")a�%��%��8�k��$D���l�M|q���t�� ��6�q狸������Z�����?dN�r��םcX�ѻ:�U
�y+��@�9X��0��0޽��)���l��z�0���A��&�<$CvAGǤW�p"I�z�ICj��b���
W�T���z:�m��6�!��m���� �bS�#�Š�̏�jq��`������iB��o;"\��w��������`Q�>	U�hC�9Ks=���!�qb�ᓨd��*",3�Ed� T�`Yc�5Wt�4aR��T4a5b.W��%INJV��������엊Y�5H�A�i�����n�'�m,C��&j�K�^�˗x.l]E(7{9�o�z�vz�e./|-(�:�Lu5W9=�X.�﶐�pIx���~�]@>���G����E+m��{����Mt
K���9u)�f�*��3:x���'�N���d:������8C�H�`:�
s�+��222$J%:�]x�V���oRp��e$�]]a,�b�ѽSBI�
�-%�oV1�įY7�!:��2��r�FW���nL$�#�����%�	�~��
���5�wM��um����d����4�IXR��0�Eb�.�����i,�V�͠�Gz��ck��h����WO���1�z�p�a\�_�V�
�z�Lb�Of����B�����빡j2��[G3����/B�-��S�`���(��Z�5VE-��2m�ي�5���,�D�Pe��٠��7&�{$��	-1�~�O��!��W%�b2\�N�#h���K�x���,�^ �H5�6Me���]iX�}4���u�$�jSh�{��"�b;/
W�I�"�>kcrGQ��jeYK'�QRӄ�x�)���>����W%w#x8�5�$NA�t,u�0^�.O���J���m���4�3���v	�N`i�/���ݢ�Uq�q�H·������p��ڀ5����2
�P����AZ�"�M��*��s�����sy�<Cv&��c�>�i�&��nˮ-!���v)�
������+<i2�7!�,�<�:]L+��8	����J��(g_A�v��h?��������|�}$2Z�m�t�U?��qE��%ձ��~?;T7�yK󓔱e�Ȍr�z]�Sp}r�����L��sS�<pW?��Zg����T����c�0�:�joơ@.n�iЉ�FԘ@��Os������󬱩l��Z�Y�26�+�����
d��}B,�@[���t��"��t:��9�td� �Դ�VsV����Vh��я\����x�Ѝ�7�4saY�13`����fu�
�~���x���ˌ~��?�5�fJ�y������7�6��z�6P�S*���y}
7گ�����63�8Ph!���T�XX0��f
s%n�L�K�! <} ���H�8��o1��-���X�v� C8o>��&��2����X�Q� :#4u�$�w����
CG��z(��`(0^�Y�$��L�G�vuf���FR tb7q;\�uC�>9:�c�.N��T�O`�Do�N�9��3Vn�W�%���g���c�����BF'�.l1����ͨ}l� �̥7X�+#�xW1T��85�U;����E0�J����ҒA~����,)=BJ�b[9��<�_�+=V�MUԦy������LY�)�O%���N�r�w��K�ao�T��6�fS������pa��9�ɗ,��m��Q�ȣ�3���rm=�~AiG��s~T�O{�^,��:��G��p3l���(7T�y0PP�c�B��+�F������}m�E��������@�~"n����A�r0]I�s.촏źZS*�P;��n Z���*6���[]����R��D/nX3�e��~j��;(���h>{K+���6� 
F��$���\�:O�ɟ���S���k���s�����Ӆ-u���Ex~�  ǔ��>0js�DÂ�}@����sSU'�T	�I=)��6��KH��o�����G��O�[�uB�0<�z��P~��u���ŝ[r����U���d �M�����J��m|��P�W��NfsTΫa�[��	l��}KH�<WI�.n���d�n��g;K�_����ֆ����/�|>��ZlT�7C��qG�d<���4u�$>O^A�y�)������ly�$�Lt�&[�
�T���ͩ�6W�j�q�W��]29�T�֝s��Q�5�V�Ȳ��(�=��5�_�"2����+Z!�;�b�Q���R���"4�Z��7��4-r)Mq&�d�q ��<�ￓ-{����y8EcJ��j������@(�������4�}��aA��%r_���*[�2[��lR�]�c/�,�4g/ ��x�Id�U�Bc���7,�� �x2A~��S����CW��Q�6���Q+�NՇ����cXH��Zz��4��ǫ9�HH��7�f�X��ā�z5��l��{��#g�HD�z|X�L<qB�+6�fmc���,�̐��1]x��Me�~�I�j�%#姚��R��V� ��73x���Ǣ2��w]�5{�z_a,�ND���ݕ�L2�y�|ȼI��'B+�x�p���t�5��ԲZ�G�.Rr�\����[���w��Ո�5����0��"��U�A/�k�ҫ=���fo����2��@�u��3f�&�h~�B�->��s��v�t���,eyޒ�d�̗��R�@���)������������`�H�А�
��C(��.��@���@�]��#�����g,�+	ޯW�`�n6Yg�k�F1���d�	N��T��#q����Xx\yw��!��s��Du���֔��`>��������xK1��N"���D�r�Th�'���[=�x8�3UFN"*�g��Mt���Bx��ȪZ�<�K�_9\Sa�T����5V�Q��p�0�X���vb{�>C�fCe�O�����S)�,����f�9��w~�0E�~���6 �F�X�#���U�)A\s��ny����j�?(���U�7�M�3Þ^�����߇1zV���+qZ\�����sZų|՞\���%+5 ��<dB��kba�P��5���^�����HJĢ�2��C�G�J���L[9��YiTxW�H&��>�@	P�����C�ܚ�:9ԂB
3¼ ��\xS������M��m�������,��q�1�4�@�_^��9��YN��2XZ�ӻ���H/>i�)����&]���dVv��,���)�4;��L"��C<yt�='D>K�����	+�=��z�]TW�[�[)��"֯��ǯX[*!���f+@')	����j���jO�%�۳j�0]^"�U�Ad�N�$xtV݂�CAG��w���0����x�E
K۲��J����
)���ߨ�s��:_�p�+i��/R*kc���3������٪��"£��A�"NH~/�,��Hw��E:~28sj�;�א]��aO��d8�&�ł��D@$��k�u6�O���,�pd�$�������L��O���lu��%��Y��̃�\^ؤ|�s<�X�EPW�-1��ѷ��d�%E��K!�_�;�'h��YH!�;jE��kQ��@Ԯ[��������J��jaaSQ���O�`�z�`���CoTn	�"�`���S.�2��V�<�K;�B�ar���{<��0�C/�[ҭ4�H{��BK �^��W�I��hٻ�|&K��a>wY �M$����F,��j��W7�J�fF�m�Q���)�T��aj5fl�EA�M��#���ǭsa�wz1W_��Ik��"G-��Z,���h0�*Ֆ�ϔCq)̑	B�`3��l�����`ɸ��Z����sd��`kGd�E@�؁�V�G�d�E���4�S)��Y:�y�mÁ��O'��N�BU����f CV�9�̀��k����oR��<�w��zc�ÒRV1[0�T���� B����CY�1\���pn��'$Qk���M�
~`��c���}�7�蠙r~�vl=/[���歄h	��63�u�|��&{~��<��R��	�CO���6�����E��Ed��G�uI6��v^�R���%��S@P#��$=;O`�G���l��s�e��.�`E��Ҩ�	���yhܬ$Qqe���і\�4>Wz�/���h*N��R3E��\c�@o��fG���$S]Q��[y�����v�('ǐT5ۻX�q_G���Z��;�.?��J��	8���Z5��>�X�2��vB�n�����WEq�}���k0a�Ndt1
ThO0\�%��&�ﱻ�Aiû�� �{�A�ۡ��rsq_S�Z�zv}�4bN:��t}��ׅ��ϫ0��q� ����&�r4[��;�Q+:�G�,a���u͈q�WjZW9`����@��vJ?sO>�rP�cS|�%���/7g`@ޠԟ�Ƅmz�q�k�t�>~2c�I�4��+��x�M�=�s}����sݜ�c�P��W�fcL��큟�˨0�ľkC��{UcH������H�_�C��1i祢oC�ߴJ��t^�T�U��
Th����M^�u��gnr��Nd��<�ײ��!Hf+�M9���W}��!�Z�Iȁ��K�C��Cc��&���YC��-Z�L&��t�MV@(�t�Q��y�Z! Km���I��5�Z��څN{��m��e�p�W��u��������&��hmu���Ѧ|8�����9#�7O���mi�H֮HxX�.�>���q�
��Ě��+��������O�U��
}�#�q��]\��G�A�_��!_Q����*|�o���b��+G6���bX�'�ǫ�N��q�K�� ;�����c&ju-97��^ DJbus9��|��|
n�h3t�3ZK��acĀe�i;��YH�����gF[i��/9�i+��C�KG�΀�)�'�YD�/(���]������%m}�Zc��7����P��W�����I�I�d���i�ޭ�����@�;g_/���!Vz��%ᔰ�_ӧ�P���	��R�9Q������r��;��� ��D?jq!����s��r+��{Gd�=�����+�T�E����L���;]0���Y.4�d����*&�Nd�r@����,5���yj��иX�nI5���QYS4@A+�2؉�Hp��s�(b|HF�}���7hݞwz�`c�,�y�	B�
C�
Å����TL<��"�y�f�V@Q2��X��դ|�ƣ�
x��a���Ra>�������t;?�~"�����{�Ѭ���~�Ѥ���7P18��{��k�}F�zS�<S����|���P��4Ԑ���k�b�_��a��=G�$2��,�uT��z�h�-��lDu�o@�S��3�=qڞ������^�ž��ɐ3ơ��g?�J��)���#!����Oo�(��f���q,C2N��, smA1�7�^����ava�g&CKtm9���ŵtiz�8�%��8q]4G6z����Z���O���A�����cX�+��ƥ�a{��搏��ta3v��zj�w���x���|�T(�0v��S)"��*�����1�_���B%u.'k������a�!�3���t�)��џ��	��U��h)�>��L]�j ���ca�)p���G)w"�f;|L&��L)�:�j6��%�+�ț?�{��vʡ����k"'����.c��m��
@z�s�-�=�r5��?+���䟒Wb�p�zdTu�;u�(���o�*#��W���G��ٳɥ�2v�X����A�����2u������n�ť�tpxi�oU��J��H�pko�b��������b٭Z�ؓ�h�Yd�럄���9��>}^�;**������1�L��֞�O��_��a�E�s����qgas^I�X�ޢ-��r�b�ƃ���$4OSQ�awW\)�:|�1�<��Y���G����
Lf�oD8�4���r�AT��ـܳ�X�;��`�!(�e	��]K �����VM�[U�������+	��+�yT����%]xulh����g;���E8t,�:���l�;�8���%�}�V�_��bKIF�*����x�0��Y�voH=��Dhq�v�)�*��t��M��M��w�)�`˭b�l���?�.��j�[o�.�ψZz�.~���4+S�$�}0���d$Ue�q|p+K���/��!,�?G4�jW�A͌3Ȅ:�p����-���z���"m#m� ���?�0㽿P�M֢���z����C8��[�O����d�c��#�q�<*�q��A��g��%��՚6c���K܁���{ʤ�����]C��R-�.|*�C�]Mwl�����=�"��%���2C"��2+j�fk���1&����7
�n�ijHў�q�2\?t��ۢ��t�By��HN��h�}P%��f<����)خ0�P���8P��
N���H�4��#E-<��n2����Rd\�'O�\P{w� �d'F�q�A֬�QW@Z52V#�Q&8�g�<��c�ܱ=�I�Y3���2��#����R��x���Z>B��~�,�i��2]�q�@S1&�r�U�^]O
~�D�Dq�cE�"OU�h����$���3A�sV�
r�}9:��j.�D\~�S�ʊ��^��K%��+7M����)��I9sͬy�2���p�R�?ھ�{�M�֝n��%%�h��\	�A�~K�Ib&�P\#��vI�l�5��z�.\$.�q��e���$u	Թ,䝾ȍY����ڱv��
�3��JL�C�rZ���3�����8�����d��w�侮��3�(���n�ĵ���6�ہ<����'����'���S4c�i��J)�4Em�1�.��!7�ξ!4yn���"�!mZKT :�g�I�Nn$f�t��8�����)g�%a/�jm �	��z��GU:r��Ӫ�Q��^�@�Q��Q��nI�c��5��ሦ"�՘{�� �WDtמ��Lc���o�]���Q�~���Y:��*��vl����F�ͮ�ASA�/Mo��g4�۬�!VS�lF���%/c�ą����j���`��Y���8ʯwz(ƲJ�\q܄�q�����f&��O֝gu�`Sgw�/*��j�^��ɳ��h�g�@��6�J�.�B+��r'�<�'�����5�����\������u�ɏ휕���VtK�#>av4���wGa�w/�"b���PF&xZ~*�v��+h+Ua�U3@���%�����u�?���%�SWUc%�AUD�
s���T��i���ˋ	TSY�Aqy�Q�P �fۀ���G�1B�}YwY�M����NѰD�h���c�CG�N$��w�Ý��%�28>�ep�Cb�S��:۰�P5��@�ɉ��R��m�,;Y�&|���$�f�HbH��[g
���ߴ�Dyqs«�mK�O���&���K������8h2���m��Y�+�l[�u5L�<��i������Hʣ�6�����O
z�����f�˕�ҝ�K'k�HY�Vw9Ǿ���� S^���_B��Y����W�G�\�A�J�����?�Y~p���)�`e�Bw�����z~�rK���b�s)�67+<��r���J-�3[�AH��8�&O2;f��g���b�zLF)�9%��/
1�_Q
�ݟ��f@9�a�uG̸[/��y�����!+F��^�k3��=�k~gK�֎bQ�[��T
)��\�m���_�gE�E��U��-PJ,!�?��q�A� 	�l2�F�{H���G
�(�!�?��ZuR���"��kCmZ���@>w!���08y���W����Lh�!L<��RJb ��w���2��l�:7�@"hO���|�4V�OFiv�E�u�y� ��l�������<�����Fu�c��$�8N�'���:�c����&�֏�����G"�0�*TZ�]�Fw�w�6��Ɂ�H@��F����,J�ú��DI�B�D=n�6�ָX�����)].�t��G�]�m��bi�WEWC�j�Y����ُ�裳�e�|O�v�kE!u��[�L8�����)MX�������aټK��T;'Z����O�]%�Zcvoo���"��[]9���<�oJ,�m,�P����L� �^�t:���el�Ǖ�'�`c�Mz �雸��$�)M��<Ra�t[� �����E�8U{�ϰ��Dx�r�9x��6��um1=���(p9��߉ی�ny�.o�dT	�?�<���K��/�s)�9n��k�Z���ؕ����h�0DE��4۠��:J����+D�aE���.�5]�^ᱯG�D��hQݛ.��J���|�>��Wf����\�za����-���#�P_={>��U��S�Np��p@H+��91�n���/������.Տ|�YNdN�n� O��*TH��������#���:[^[�U���k
F�p����X
�J�w���Ct��14G1�æ7��ЮVð�C$m�Urv\���1S���,�2Q��U&�~kGp~"&�{?k�vL�@�Jn[#K
�i����;;�y/R��4���_�Y՟�D�B{w��%/��\����D��K dk����@�3���l�r� ���c��6��|p�?7ݔ�L�6����MYv������VG���+��WG�x5&R�Z�x��w����ue@��R�=��R'�}��CQ��W=2fc\����)�2�?����D���:̚R��D�AR�^�=����\;@����s�V����}�AJh9/f1�)�G��_垞y��yl�9CK�S���z��e��G W��4I|raAK��L�4�[�I/���h�3/yr���%���ڇ=�Ea	��{\��e��<�#u��~����I�.`��O�bn^����J��"-��!�Ș��$έDD�ķ@6�����8���@L~]����Jÿ�bv�f��L���z��~�Z�2 N�b�l0�!'%��^���#�)�~��QP`&�݃ �+�"�3@�M����\P*j�N�L�ى���po�D�Ew�B����y�@[�PRɱJإ&��ޘ��5Ⱦ�����Ӯ=Ϫf�Ч���:.�ߋ�W�)�la��o����ޙ{�ծ��7݊�����=��[d)�\���38k��okƛ�=�)�����OΟT�н��L�%��@�X�	Ga��־&�I�J�������S���� p��]����^m ��u�N[3S3���+F� #�PzV���0��X�bq �RF��g\ܮ���=�3���L���?�`F�8� �e���(�<9T����M|=Ǚ]��}�2I��w�B~�A�4ϲ4�g�ca3�w6�R��b�L��v�RT�6� ��TvZ2�Y��|2���;��ȄL2eW��{�j�K�WYʃif�� ���>���#|�S�B�:�J�xh33U�hm�E9������Y�1a6�ݐ>�L�û�j�|�����,lBc7(���_�-!kѻ�U�n<V+�VTg��|
��!KhX�+�	퟽Oѕ�H����Ϥ�iB�B�An�=�0�ٓ�G>��%B%�k4�<�r�:�B� �x`������T�h���Q�I	�tjF�g�xp�	<�xک}����i���4=����`DM|��"��;�;����nl��H�!}AU!��j�n���4�O�t�����?�K720l�>��v���]u��N3_n��2�፷Z���Ev>�M��HpR����d&W:4_ө7�ޒ�={�CvyW���͋ ��V���Ɇ�S��^�*��aֲqݘS�?] |<�v����eҼ�OK?2)�J:bv���IFE�<�Z�{?V�ֵ(:@���Ա�I�?���=B�Q�S2M�6!{��>�O� �^u?d7��>3T8-��$�̷��ԅYz���uj�3�aI;I����B���'�S��'��M�O?l;�����'���C"A�YW�q-N�����(~g~��� �����ؾzA̏��G�3m�d@�h`�݃<<,��{Kxxԙ��%��G��<�Eۜl��쭿�lK��S��� T������'w9�Њ3��Q�`L���R��.QY�X�m}�|�fbҺ:}T6��n��p����~��0b^Aq���0��n�~-���J�,*��J���z��Թ���9ѠqW�R�$y� "�U�@��K�9V�ܩ�F��7��߭QB�n
�D=I�w��!�˟�p�(c=U�=���/3)E��.ETP�(����ΌLic�;��6Q�J(�/�gNՐʝ\ �+�{6bc��
��	W/S!s���-�`�@���Z�p�
��� 4�6�{N�mL˔�mk��q:W!/���c\H�g�z[xe�c��c!�z�6��,G����Ÿ��e��:����p��Y霌ȇ����ow@�]�v>.�@��݀,E�Fߛ]��6c�q�� ���&��Yl7�s):�휕$��Dq]�%<H\��� �]�cG�&��7���!��nX����W��$���t.��ʙ\p5��|G/U]�F�r�F����ʡ�/yb`��C� KE���lت i<��M���B�igiz��'�����~:��B��0Z>��~�飫tQ_YY=�����8�"AtcacfX��U������L��(��C?�tr��\a����n�0���m���$ܱ�Lh��:K�06?�.�їC#c��J�h��n�X�U��퟇:�Y�0Z��x%���z�����T��:�g��ZB��R�?����]MLs0R�K�<$#�ތ�H`�;w��vk_c�2�aXRLP��Y9��̦?;����z�+	�;�����BV\50Io�uud����J��P�����>�	�k��Tz�ש͐^N�hFi(�\�P�����V&���DM������՚g�Z�wޅ��u�#��g/����Su��uO�j�Zy�
ohs�捘]�R�R�ZOԇ�������������)��'��/���z�+�KIW)^3v�t5[����&Z��0¶����a����j��������]K�D�`�A���%+8�Z�4n��{�WY�KZ�H�Y����L�����mm^hcr"ݸ���~[U����` ��q��;,O�GD��ֆ^�Ga܈�։y�9<*5�g�%�����B�kM�,.���O�#u�ksz�h��՗t9y���%���]��3���xg(t�q#��T�TA��VGV2]����Ǚ�TQ�+u��G�!f
�m<g�M��6�@�Z����N�ˮi�	W�J�#ؚ����]xO��5IG�D]beF����8I45�x��(W�~����}b�q����K�i[���H�m[򖺱����w6�d�#N=2/���XA *�%;M rI;MB�PC��#`NnG#�V{���6Z�xcoo4(s�J�y�P�����H$�A��×2�Dς�Vy-�:(�Ђ�*�Q�Q����jXrB�`��Z��r�W�,��#ﯠ>!�E�z�	ͷဧ��k*���ՁiE��0�3��bT��&h�B�RI�{:x\����M.i�zQ�x��
o���Hm�`���)������]�Pq�06����&�q��F�'(7P��f��7k� �A���[��il
n�����ܔ>qJT�?O�s68y��U��9�����+0�}2ӳ��#���=��?/b���u��74����E\���?�:�˚r;L%}r���Oh��\@%j
yn�~e瓅G�������2Z�cU�_ݴ�*�|�nX��az]p)�+��^�sD�k�#�Q%��	-�g���`4��J��p����Q�K��15���P[�p�}=<_0,2�tض �S�*�QƋ��a����=�
����&Us�EKX�(��j��'��I:��w��r"X��#ȣ�>�cx��z2B\���|鿒�+�s,oW�M}��̂
A�|���
E 4@�C�<]��oL 4�4�ki�@��^(5�h��*��k���GA�QU!u�$B�I�#����n>q< �=�ڠ@z�!�
�W�w��C���_	�fj'�S$�<e��Hm�h
�b\�y��s��R&�M��>�y}Zy�Tonr�(�"�(U��g��Ew����T�}���E�=�	�
��~�"�������Z*z��yA.hį`�������Dƪ���0�*�
�n��>������B�cP�h ����G+e��������f���':}�UTLU"�y|/��F'j�ԚN\�)�O��*];���"��$z����Q��9�ԩG��``Rg�?"��a���"��^����z� ���
�����[�N�iJ����l�}o�,�5`�x7Ui#��!�-�1�d�.�fjBAT�Q��9f)��]~�����vN}�������ō"d6��C�>w���=�p�I�,��_����"y	~`H�97������y�Ǐ�r����o�����p더���K�w;�Z�Q��5��TJ��s{����;��}���^6r��u��e��kGT���[��k�hM�7���%�Ņ@G^#��=e%�����d�
�u [GdI����'?�v��k��>g���L'z�����ɿ����àw���.KaT&NR�V�kdF��;p]�,�+��_���r̂�\y ���y#zB���ʓs쀂��K���%�����\2Z2`[��wB��A ȕ��4�%�Ə�[�L�\R�{�t|ۡ|y@
�E@T.��9�hMy|��M0�K�ù
���b�����B��]��w���p�5�(��Oݞ�p�����)EPh�+M{X��6�/t|���P1�t��k��Q9!�ld��ꓘ
�HX���y�ߤk	�N���0L&X�"��jA�Kܿ���[A��A�^�'i�!X�Mٜ�Ŏ掕fwJֱhR��K��>��&���������@}+=���Zq�2H@�&�q2��;�hK(1��8��=$�1���,
��D#	�������ʔ�+3o~\x�ՃC��]E�ee��'����~S\tY`J��U��ӊ�[��zo}5��P�x7���7�u���'b��i�Q��^8���>��Ȏ�N<z�@FI�qJ|VW�����;�{�^�&
a0�z�b��g��٠�)Fb�&���wQ�1���&�<�- Zq-IWoO��-���<�����d#���8�K��	�Mxfg,�0�[I�֒�1�2&��kf��+f�D��'��o��^�Z�b���Z�2�[��N_���~��\�S�Y���)x*c��*q����s��OZ���V��B��u~������K��ʘ�CAiUB����pE�e�$���|��Aת�.;-��pTq2��i��o��h�����5��GU�E�ܕ�!�ȏ<hq�M4��q��i��pMWE����E�m2�Ꝗ*�M����A=�{�C:Q��y6�Kx��yC;�`��#���� 2��oe�ލ��$�����9t�g'`�1��vWg�f>�&XE������HUwN7�'g�>�Z��J�rD�������Ën�`p>�([���5��٦�M��|�Oa.��!�\C�R���T��B����uh��ҁ�޽�5������{5�L��@�4>�7�p��RN<)����`��tO��|����F����;�����J1������9"25r9��Y�b�.�kA@�_��h��L���8������b G�_�`�� �d�{�h��%��in�"��,]F�Þd(.�7�-TB�(��i�
��[�.����~2�n�����b_�����f
�Nj���>,첖/�J;	�i�Hb���a�]���A��p8��JO� a�_���xIQ&1�ϒ�[{)��gџm3G��Bz�"�.�_U�ɂ[�i&L#�ǪKY���8�����1̵,��<��LHk�CS�4�`"+뾃G��� �m�Q^�6{4RW&m��^g1��t �x���D0�����Kecv%+�ؠb�[3��)�ÎC��69H2��ٴW�낔�}?ge���ؾ8c W��:O�?S����
X�6,�ko@�M�s7SII#���Y.k�2�O2�Գ����T�jJ0Q���ZX�h�����I V�5O+l�vK ���)�3�U������1�f_��7@�FC��:�E̔�F�0o�MwP�*޲��߾@NBEp�.7�t��˫Z���y ��N�փ
��`(�)�IdF�el	-W*<:((1�N�]k�����$���������}� (rJf<�$+}��Y#�5�g8F��3�����K�My>�9p7��N�
��XLx�ϯ<%V��|"&XiLT�i��V>�B�?�P�C��݊|�b����7�^��!����(�8Z�_l�������N7_kkXE4p:����U�XD��%�����z$�Rt Œq�â=�%r���*5m���M�غ�ӣ:�����,����1��� ڟ��Qs���5g.�(ḽ����D��0��
)����XFD��C(�M���F�&>uN���mo5���uor!���{�7j��	�u��lB豎FH0�)�*�a�`����hX ף����,��K�O�8��ޗ��Y/v
s�oy�,h���k��$}qjdI���L� �|b7cҟ��q�K��y��P�m�+��蔪;;B3N��*��pk�H�>KB�"�@�)�-�R`D�����U)����&���˘��j3ǟ�����eJT3�t�n�>�6�7Ϯ�	5�mc�VBIw��
-#S5��R�eA9Jy���.i(}̱�'���{���d���Th'�](���2����\k΅�zp_�I
�?����rf�xD7�0Fcw���,�jJ��֪W�����t�|���թ�x#�����ƨ%�7�ak�Z�;)M���fv4�y50'Z䑁�W�T�I �X` 6J&r�i���@ʾdZI�2������� ��A��ΪȜ�_����������������}�4J��=�����^�Ib�l3B���Ξ4�(tm9���򊩆����[�����E+"V<�d�z#�O�~����� �^N��!,8�׻�H�Hr�T�Jo���I�Y�g�_ti\�/b:��_�60��W�r�掟��k���/�i�l{u�Ū�Os�3�+g���T=�3�� H����N[+�u1X�5R�`���i�����s���X	�0�>�A/ʔ��l�*��?��ǎ���+���A	���5�D��	�k�j���~���B+'�S�����l ?�F9����B+o㔈:d��b(�I��*F�V͔��_%�D{g�/�ZeI#%�/0�˄��S�WQI�)� �x�1��G���:P�����:�5r][]��$P��R~�P�������u�ʑ;�4A'ݶ^I%�I������Pe�^��j�	6��3œ��������E��9�d���;4V���a�d���"7|��zZw�һu҈��Uh��OA�?k+�(����ϊ�z��a��f$>��ua�A�R���Vn�����lN�����e����K�RgCp����M������X�f��=)�����j�Sn4� �+��:Nz!�;S@~IW��6����
O03�=9����)d`%���C��3��Z�~XCp���/X���h����'��à�v�#���@�1-Vr�t�X(���TTƙR�՞�⤩��g+��O�-����^��`"�K��v�	���������BM���28C�	
7L�m*�y��u�5�0���r��=��C��h}�c�[� ��\�-r��-(�D+h���	U�B��Ņ��d�v-Ba��������C��2�9Z1�ٯ�<�&��_ϗ�S��Cg��O������o��o�K��� ��mio/1�%q[����e!�gr���7{��yy�(`=��ƨ?�h}����I!�2�.A���య຾�'Mc<F1J*_ȱ�5��k�5	����=-9�l݃�*��F_�|�ڎ��1lDML��TJj[D�N ���cW{�B[�Χz;���2c�X��E=ez1}�@��j���5� z�!�W��P�KWm>;����q3U=(F���'�
��w�|�6\�a�re/�$��X�.���̞Y�z�ח��BhU�hR��w�X��1�G[˨��kKB `Zl��Y;���Ns��>pq\<MY[�ی�.���0�������F밝=�w�\���u.����!��օS��c�� nE��G4�K����dQ�ac�l�G5-��mjoS��q��@LP�� �&n�W%4F�kI���Xq�c��
�4�|p~;��G��ŃHt��i���}t�w\�p������I%R���J]�`�\���0�]@�1'}�j�k���x�4�Wz#ߔ��9��o���34�T�+/����/ifd���`�J��+6���s{��	6y���
-G�I���|�\���mB�#�܈~��P�yH��pr���h{�:�\~�-E*��&q����z`E�YiǆH.��b���~&S����Y}\T�Tl�Jc2%
��O�8����'\���y\A����®�-Vibcb����0�XP%b}�SJOO6��o�CFW��xfq 
މ+�#�K��3�P�~�LVԕ|������|#��*�#j<��JRh�id4,[��1N�9�iE�*O�Hl��|�h�8�)���<��(@.roO�n�3X�tn��6���C&了V&xuc�Ţ!X�J���8�GK��lM�K\I����*b�p��r��H�� KMP:v�k���Ε_���Ga��I��r�;����aq!���o��(hO">�^���A�P�V$��X`4u��ٺY5#mI�<����0�-K���Y�|�0���Z��دn�T�qY�М2��9�ģ>\b`�A�
�̈́ɒ�B"���, *��O���J�w����_���}J�TV3�ӌ�ɧXn^i*���j�����![a�,��s9�"�3��4p�dk�NEopT��/Nj�kX��A���y�ԍe�Ax^g��
��n�*� G˰� �W��A���NJ����U���']V*X&��ʘ��A��Z��6cd���g�|�;�Jf�e`9���%�U�o��6�gd:T*3����sD�v�Ҏ�	��H�m=˩�mݥG@�I}^�0-q�,�'x0�C>�»�Y���kT�~���)u�:W)H6��nՍ���������F�j�`�y-"!�W�]�R�]vbP��=:�
QY�}ˆ{�Y�_la�$��U�"�H�nI;!�}�}3,�F�nz��v��I�V��X{,�ve#)5��1�w���fD��Ic=5+ן�L�P�IH���#׎O��=��-�O�Mo��z.����-��z���4:�䂠Ys�# 	����Z���Ҍ��2ԗ!g���@:�ٕ9S��2���}���o�C��G�Ͻ����Kw�ރ��������쉫�~�4�Vӆ��.��X����8����Cc�N���2����uh���}L�=���e8� ��v7�K�!O�K�C���g���^1�K�V�@�-I^m	�7��P0�/���]",��L�9�E5���mW.�����[�%-�䞈���; b��/n��`8�A��	J��ZY��No�afq9K��|空��� W���HgQ�b�ԀQW4r���Ҿ@8*�t���\u�jw�<n@?=ת�G#`̢5�����N�����ހV��H'mT@�*G����1�G<\��4����k�Dmt8S&<VBn}�@�r[M[߃�H?�b��a�w���7��C��bVգ�.�@.;��a`Cw��HNn_������n����Z� ��U��_ڮFyv�Եj�C���~V�
%��0�����S'J�R�%p��ӡ�lHn�r�;[���`W�֡{��%���n��h�'�{���
��-*��=���tީ=7�@$A�WN`�MO��Ovϓ��8p�FG��S�Q�!����_L;�?�<�Y��B�A�1 C·�#��F� W�gk�7cC~G��f
)��V�	9iY�g�I��gL�~$��@�Ƭ�q-	�����knj����k!�5����U�<�R����hN]%�����4}�,<����	MW�.Ս,�=��O�3]�=n�굩�dW=��ۑ�mo��8o�`�)��	8o��НD#�S�R���N�-Mx�T��u���3������Sx���
��� ���'�3Y�E}��VV^I ����Z���E^wo�s�.��YԹ�9k�Cɒ=F�i���������LE�'���j�\vC!ӎ�g���/�n?Ç�l���Էp
͏u=
�ɻ�IԔ~*֘�B�&gj�XL�g��B�l�
������߳�w�Y��>x4�yM&�F��=ozk���Ex�>����`r%.J7�'�����]��s�0N"e ?9��0�	�4���=�������i�����<��N"�8��O	N��1��n�DmY�욍Q�������K����sߛ9z�H4^�Y氲�*e���,�;��b��C1<"ݐ�ke1�
�^wnߞH�d��jۡ����
D��ϫW�4��D�lv���&S�k���հB��"�)���%���|a�ӝ�J3���k��H��h������J���.�rhosF;��G���j:b�b�@���Z *�i��1AfTUL���bfb�JoA�)���a���cǊ��~�� �Ʊ_W�Q�p���s����	��Ff��xƃ������q�AN(oDʅ8�j��E � KOF��Fm��/۞)�	fvpe���ZT->֐_$:��5 �A㫊~g���y�è��NU�	˶f/��4�6g�( ��q��b�@�xh���"�/q�1�o%�b�f��5I�6�����'��pC
��6�Q_��*��嶺�v�X�ܵ%��B!���Nu�B��'������G8�ˉ�I�~���(K�b4!{�&�h�j����R�ۍ�n`�l�E(���h�� /KWT��jw�_{8F��kWv�[=$=�e��bӎ3��|`0]+��
���؟�t��,=��X��B�&��g�f�?�U�
\~S�z�+�x��LON���t���l�'�k�^g�{Ta�:t�✾�Fl���6C�X:�c_�6����}����`) b�����i|�(3����;z������Zyn,Ɠ2�P����L<�QJ��[OݾT�%��J���KE���*������u��|�8�ӨX[�D�]�; #��y�S��@*`=n���8.�ȣ�Jpm��ZNC�M�����0S����3���'�����%�4݂z��z����[�_<|�C��QQ����w/w�/�j����y������MP���9(��E	����ؽ/de�-���0����z9oT�����愨ň�s��06g�؈=<���޶�]<����x���=��e���t�,�D�?��hSa¸+�������3�cZ\���v!�i掗�^�Ռ5�³��� �7#���n�x�Vċ#>7D�<�1!emRG8O4&2�9�y\�C�mf6I�;��g��)� �j��Z���?��|�\>P	7]E�B���1M5MqՓ&8����7G��2/�;�/`C|_�MR+��Y��9�x���K>1�j_���1��c�)���?0��QįI� ���16;&��usN *6�\dyg�̻�F!�UjS�s�g�����x�*]@����z�|�����xp(���\>Ϛ!t��Q"�aC�?ŦQ��w"\��"�o�8=S��0�{!c���o
�A�yI�Τ1$a�G���r$v��wд��H�x!��6?�rzwI�I�Z��}�S�d*���^jI}s�]!��[7h�b�'�����':^6���4ᡬ�����r���2z����60=iY�ݸ1	��{G\��o����j����،/�䀖�z�f,�V�:�xc�c���O�n||���1&ZP)V���7:C;T�[�!�+�V�W���,��!����lP,���b��T����������l�`�=�<�g�t�]�ʋR+\3N�4jY���i����G��Z��p�: a ��=�#�����NJ�uj�]����* I򩧕�70V��)� ���W����f�~���NTylԃ֖�����/X�\!t��82u�#c�F�K��|�ɟn^$�������z��]���v�	K���I�:x��o�9���L�X	 l�ܫ���0����+}�jr���@�|� A���kH��.�/�|���;�����m5��@Oު%кO�9=NMX�"К;��ht�|�g����5��W�k�2�/�[���P���
;$4�v�Mi����ᥑ��x@��^�PD3�Nv��r��5S;?4�l} ��@Cի|���:�VO~�"�����+�V��(�k�L����:1���l��DLG�Ol���S�p)���h!��>Ä6s\�tY�����:��wQ*���#��)�/7c����p:-k����k"��6�͕ �S�y����y���Ցed9�iF�N(��7\�S��v���k{/��B�ʯ�m����c����ؠ�ȥ)�:#����O�r[u�AR`���X���y���Ƥ�SL|o�V�?��Rqk)��{����7l�(��9�<�S��0��$k���"25�s�9�^iH������ò�m9�������k1
!�� ������t�Ш���p�&����L��k� �
�~A�	��������6,���U�' f�D��F7��õfZ�aGW���+B��H�9re���;�c+:���ŷj筶���u
ˑQ�����I�M6�3t4f��ڹ_��^��j����NS��Qx��sњ���TS�����YcL��aF1�����蒟��f�{�	�z4�u8�[�%p��k3u|�C.�!���?E[�p����(:P�����`/�n�d-���d��L��7O��Mv(J:�]�I�i#!X�7��|�$p��%��2�EB��NH��-zD�����2�����*�����h�R��gp	�����Jn�h�B�e����Y-B%{FR�_�l˒��`��HnO��cY��_�L0�+�f�mT�%^Ѻ㞆̕�Q�Ԁ�!�I��l�(J.͚~ƨ��������2n<���O!�Sʹ�۱�%'�X&�/w��Ѕa4H��)Hǭ�#^5�=~*{l�!W����>[z�Ұ��w^qcu��ݭ�0��ϙ��Wk^H�S��AY]̞<��ʪ'�|nV�����R��U��]O�2n����C3�Z/.�ب�#5�jb!�V�V�[�``=ʶ�d����U=r���n. &�/HQ+�lg��K�,�� ���X�9i(�C��#��a+;���2�|���g��P4�h�֨
��:6ޜD�6O�+R�OTW���2�N w���4
�y!�(h�s�'B(�U��{j=X�kZ]�mC�ɶ�B{z���� T�u��7.�~�
����&�@
����V�֓_��}�[��,f��C��ZZ���D-&}��!�4{�5�M����(@-c6d�9P�<���y�4��-�⩱F/�-�D���>GۤYha��{�k# d���l"#d�I'ocO>ʤZ��),�A��L&1�XBx��,!�@)F���	�����-�pO���	��1�s�*8�bV!�s�ͭA���%��J��_A-N�9ɯۨ��h�U0x!���� �Ǣ&�g�ín�� �l957;�v%�>5�W_�:a4q��AS�S�a�O1�zG��� Lw�P�Y8S/6'%1M�.��O^����]�2g��(B~3��~}s��hF&�s�.�F��#k
+2��������r�]��w�Q�Y�����T��ֈ������Rq+�Dn=��В7pC�Gn���%�5B@�.�����]졾.�YA6}^m�r��* 'D6�&�n�lb ��������u���3S�� ����KY"́ވ]��i�+��>� Λ�Qy���9�8� ��?�oA�D��Ȃ ������4���Db��a�<��9��:���=j���q��]lSBC%��9+G8�M�ܟE����3�&�89��\�7���/oMH��A���0� 4եD&�����`�QK+����k�v��1�8ؘ(1J�����*�۾��&���7]V���b.�B>G`|Rcd0���"k�mU������	�/�\N�a�� E-ȜQb�љ����t���,ɢ���a�_"%3f���d(�I\�B�c��D�Mt0���� ��/n��s4�QV��M�E�KM ��d��׹|���BHu ��Fy��3���j<�U^0��u-@,�m�MN�����*�L��M�s2�g���iѯ?�~K�;�t�XRSn,�Ր��ܵl�C��ì��+4aĳ�8��!��'�"}H.K!�2+i���d >�r*�=U+�x�_�S����*i�&��#�~,�͂Bn�$8����	ը�_��G��,�l_��n ����ee�:�5��BH|H��4�)�Ӧ�9��&�W�r6������	���񁺅n�ۂ2�y������H�&���5�.J�l2�0���=�ئ����zd�]��Mx���ԑI9���#��ͤ:SG_���OR��.��%s理���^����x�hmd�}������tno��v��c�<s|=��m���i�*PL�U��N���]���t�����4���5S>���7�A��VI�*� �+�����&r�+�n=iփ�P1A�¥J9%������N�s^~B�јI
{M�NP|m>��-���V��V��or��",�Gt�ͣ���!SՋaŅ)��t��jƞ�I�G�:�)]�Ŗ"Lbqr��נ*��<%���(���y�I֒{kZ����N�>��� �x&�ћ?5V�4�w=`񏼝���C>�'�6R��a�1b{��9�ʅ��D��Y:Oi��v�I|�WK͍�p! �R����o��BU��#:��憎yR��J3s�͏,Բ�b;
��wR�J�$�{�������%:�<�����Ku��1�\��W2�ʷfX��Y�2�qU���uA��jր�����HTh�LuZ���*��'�}�j����3�۸I]=�v�}���a�m�:����#�\J�E�pT{�x�e�[��YE�`h��ގ�Dm����h�Jt�|�!;0��Mw����~�L�šj�-䓌��D���-�{|ֻ
��&�q7�[j�I�����)n�t]�z������HI�[@�'PN���$�RgzO�Qߜ�����X�'�$���h���%�o�Jx	�P��g
���5f v��U��IE�� �P��\q�YUv?7lh�Y�]t��k�/(��K�L;K��^�;����d�\�?�Ќ߮AJ��%��+Q6���Qv�؟'/��f�(��\���W��g��ȱ�o��Ҡ��P�!]�{0�>L���^��v�y��Վ)G�0�40Ձ]@x�Z;4�t�xm}�y�W0���r�ʩeL	FܖK����$C��	���aH��cv@��T�펥�v���E���`��b�I^�m�%����a�ee� �1w8E�4P���%���q	%�O%�[B���D���%B��&#3~q��Pc$���ӏ�S���������hPz4�n�!��wX>K3�>&x[��fD�x�眄�E<��[js��N��$A�����7o~0�%iB�7b�����KLz�j���)E21���*�P�寖o�Z�$� % ʑ�a�!C�I�d�f�3N��TQ ��0z���w����u;�l���7J����^I?�==,��yV�}g]Y���8;
���c����:@��G!u�Lȝ�����zת�c\�C>�J�t��\)� ��a��8������Ķ�0�3�ߡm�#햊;�&�w�N\P'r\���\����v(��4�,�.��x�d�/k��H����D�>�2-�-.M�u�h#m[�����*� 6)8O�ӆunH��f��'U,�r�er	6|��l��~���4�2�vj��+\�ڇ�qK1}w�
��y�8Φ�w�O�F������*^����ё&����Ax�T5��4���#��:��@����QǓъN0hP`4�/1����O#� �j1���:�ǃQD?L����W�[*'���sg���Ay	�����ܩ�Z�P1o����?#]�P}��q�˩Tp/�9���b���(д��� ���� ��3����I��k̏Œ����p��2��z��^���3c����|N��a�A�����57;�~��ޕ�L�$e�-�sR�p�����>�
9n
��V�T�h��{G��>``jRa:��57�#��+�566��uX*زH(I7l��6� ;wު�F�9��3�멚l���L�ﬂ��'>�(��'�s&u3j��	[�2��I�d͍��O���mϜ	��(k�/�j��./��G��KE��l�9��u�IY��P1cҾB �5mxV6&zi;H}��j�Zg8�H�R�z��*�`L�},{Ñ�x���l�DP�S~�7iAp��hr듄`[0w��4a��H��T��2����4���mj�!�Y�����*�̿U�j��c���qVcL¤>y��f!�y�[ضC�R9�[p��o���ٌ+�t]J�	�etgO�1��wqN4�G�F.�HqY�س����J�u��}�L)�I���"��� S@�:M��&�u���an�&M3���]�b- �$+c>�>����gHf�<Z�2wV�@�6�:)�{g�SD���3*�޷f�Mgnđx�+i U~zl6���7�	Q����D˒��O>�b������EW	�������E ������-D��Gu�Q�GfƇ�)�V����x��^����謘��6vK��Py�$�ū	��f���Uy�>ڛb��o��Q~K޹��CC-��dԞ_�¦��e���R�3��u����@Wx���S�H�ӕB�f�7V�~������K�E6D߼�����m�*U9����T�<RC���Σ
���c���� �7^?z��m��E���}*�����K�;*���J~��?�+ۊ��I���| �;R\�蟲�m|�v�~����[�.�i�P�b "�(�plx�����_;��b��}���#���J�����u�
s�D�	c#H�K�ԟ6HD�3`��v;��D�A>�!p��f�䵆��i�G3V	�;�z�giLp%H���v����<��a�Qߒ�UፍX���
y�E$��'�Uό�xJ�L��&�J>���s�ȝ���;����Xy����QW^�uzKV�͋�r �U���r� ~P��K��?���
��Q��`@3Ek���
��&e����c@�-+��NB�P�UE��F�̃e�E	��E�$�\�N6�>�L����*�xp�./�3�8C����P����3l�s�T�o|}o��y�6�h
�G�&۟�_�Q�tTe�Fg&�>��,>�ſ���<���V��ڰU�G�.�v�S%�~&�
ZJ19��_�өa7Ï�i�5+r�^����֤���7���9��o� ]�df�#���O\�,B��e+���I��}̍m/�Y���DX��߆��T��X-N����GV%eߟoF��h^���HL{�uH�����]I_���d�~�cq����C2�L2W�֣t������VM@�#�9�C�Kx���2�\��V�*��gsY�Aze��c���^�ܣWIe�`���m��ؽ�5Y׫�t��i���Ȃ�c�,������L7g���s���2����d�݀�� ��A���:�=_nݝ��[49�%���(H�Vi�$��������Dl�8˸�bǿN`�=g��(�uj.��	��Πo�b@���4����PT";}P��nI�:�1���l����U��ı�]�t:��F�r2i.mO��[�|\l��>����ݩ��S5��%%�N f.�C��� ����K>G3u��r�z9RE�=�'
i�V�z���Z�@Et7�Wc:��7F�w
�@���V]��6?�خG�%-iF�9[���,���Hj��a�Q^A��XA�q���{.����[--]#���[e�1���n��no����d=S�7H��;���J" ���z�|ű�&W�t߉l�Z�3��%|�& �@��
"Rc�y�>�Xf6y	�)�KD�ʴ�^�~E�$�}m��0�C*�(]F����k.9zJ