��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2�(�*�!n|}�,+d��黯�"z(�Q�����fhb�M����B���Wb��*;��C-�q���5��6Lf%U�	�����[&r�;1<T�M�����G��8$���}F��G���0,G���:_k�����S�s&�!X��tڬ��VH?����A�ZTd�.�&���:^�&�H�V���wc,7�r)� ��������G�ʥ�VB{�lG���e�^hn�?��r7�6���Y��
���bU��x�����琝$I:D��(́����'י�Q����O�=��(�xT;j=wO��^�6���ef[�bA�[
��׾?�cl�˳8.U�� �b#	!R�o��̿��M�K۽d��ơ/�՗Kw7lY�>b��jq�e������H��̎��ZfE��T��DC �D�Csq�a|k���2#��}=,��������1A	����6J�'�7DĄ��$7�`P=�J!��ճCV�4�)�c�z��א�]-i�O)��7�p'j�'�A֌��a�߽ā]��'�o�P���]�o�|!\M��gY��+�@
B��>��AmV���
��EO��~^��
{�{��Eu�9m��5�����6xK��v*%��$�+$�����C���x�<����y�kX�䞁g�@_=�E�'�5�&ʆ���xk��2�g8��� 4�ɰ}�eg۴��Ԝ�e��Vbȗ�wTܷ�X�ȫm��d���.��Z�tgךT%���_R�{8���
i�ý:��5�H���)�G7����D��!�^@L���@R���f/�]}�h���)Y��Q�S�+5��R����]�
8+����g�:1aL�ͤ�٭6Iq���KyK�3sX�4/����/�Q ��v���i�M��������IGc��f�n��O��^N~s�M�d��e,��?�Z�6�7���ZaE���y����<ܧ�F"�w�淭KN�X%rZk�BCSШ����6#h�g��M�_T}8�������h����W��f��k����"������+B�r=8��Y3�T�T��Kʼb�`�q�D�x'�7=��BFg�:�ȡ6�Q)�qN4Dd��� W�9��O��E�n�'�5B<1S�ZH��a�z�,����,�1��~*��x�����مĵصj^+x �.�f,��5�<��&��x��	^�$I�.�x$�B0���vS#f����r������떂�y{�,��S��|��y���|�ǗW^:��lRq�73�{,�� ���}V-�D�� zO.Jo�s��9B�����T�� ��j��):��� �����]�4����55w���i����J��l�LW�l��b/E�6X�J.�[�>�F`�m�?�������@����.��U � rU���f5�m���;�+A��@�t� q^<v���Cߎ�K<���H�[�x/�o66)T���KK4J<�W�$���JMw���`E��:�2[�;�s�i� ����o��%�0>G�Dؽ���)���D�4�L;uj�3=��)��6���~5��D�|���>Ҳc��_<�G���.��^l�O/6^���A�Yk��/X;�yLNXh�gB�ui<�9���,��,	�'����U�\X�6�\�ߑ�Е�AJ���.\^�Tд�F���h��0{�����*��v�$r�"a��x��M����@"�PݵC\ƨ>�ϹS$(}qH�X*�~�m��5A�Eė�U	m���M�~pa�J�7W���-�c˒Vb@�+\y ��K�������j���>�1{	e��%#��]씩�xo�W�=ss��U�ɷMJpC/gU��>hx|�T��yQ��43W;tϽӎ���4�=��_����"{5��d�G��ƞq���/�s�v��:O��%=���%�&~Jј�,�ܦ+�0��f��Â�K�~Ӏѣvm��M�n�S���_�Rܮ`-YOv�3�.�����yT�,��~�Җ�ԵX��f�R>�2��x��z��"��7��3�9�5�.���N�������%�7���4�%�t=�����n�����Phds�/S�������Oh��{A���]�Y9#��풣�B+j�hk��kO��hJ����T1�wEm�IP14i�F��LQ�tj�@�[1��v.��9��t*#<:��j�3���u{9I?�[R��f�Z
�l�=���9����~�|��Aӎ���Iy����)�,�)�Y��Fe����:J�n�W!��
����k:;����D'���^�#x>Җ�̦ �z�������������qa�3��M��?�E�~�o�k`\Z �����&�/��V��Z�kųW1/��&,{SzD��̮���e�Ѝ���/���A3�P�D�V��#��ANT7p�p������o��UhD?�,�w+�D����K�%}wh��;ʤ�	���pm�w]bm���>ŷ�q�6�'>rm\�S?áV|j[���f^\�[ZI��Ȉ���y�v��o�>�ߓL����ʖב�d�>�g�;e�]�����q�tH-�#��	��ڏ�by��U�~(����V��f�M�ρqq"��Y�Ǟ��.^-��-&C���w6�f�㮙ve��_'� ^�!���}�w������.�Y�v�_<���s$G�ux���28d��ƞ��K2�����<m�ӭ��"�H�)��d��/��P�;Dﴩ�LXK5��+m%92�.`C��I�@l��fE��$a7<hDR������Z�=[Yu����;oDY�!�io�_wL_3}Oo~3WU#ûE�0��#}����t�_�4�5J+=�}�͋�gpd���XqQ��a�pZ/���q�"�H�;&Z�X������Z����C�2��%s%$���<��E&�>E�G&䩠�n��py�C�e�r<
X��!��h�'�U-ʩdN�/>A9�dk���"�A[ˍs`�v��F�t��)w��&"'y�X�v.�z߽b Q��t�j���<B�d��|2���&��_��xg���lBej�������_ۤ$�7S��,��+���_7?=���(~���
��*2��`�<��� jy�@���]z��&���/������Y�C�Xt+(���WL嵗���YH{OV�i
��������f�ik�m@,K����T�4��K��<.��ҍ��S[D^����G��-��k������P���$�)�I=�gR�i��}���w�좄���{�B�f�E[��|�YɎ�ċ�C,�Qr,gv�<um
Q{k��Z�s�o "f���g^���?7���c���W��-6��^�o`5ɧ�"�>���ZJ�T��,�-�UTA�e��C�'>�GJ�a�u?w�J�Y�PmRv9�gF(�g�R=���;d����|��nr�\,��AqU�����V\g���:�	\�����D�� �v��.�^S}���L�XA�*x'� 5��@�E��)�*r����Kf�kY	Ů}�ܴ��8#Q���*C$I$^\�=����@R��-�g�<�A���S���s�)����ȑ*p��܊ �����;���=R\��G����35y�ι��Dy淇�%��O�k#$��[Rգa0����%	?�� im�n�8:�����gS@P����$���H_��c:��wa���蜁}�2󭁨�=�MM��	�7q�(���EOD���o�c����Rv �g�0~8�Yؽb��Ѡ4����=��p�Jzt�.8�v
�&3���Z�!,��}+`td?���sj�E�A�J.?��[��$���j�� �-_�2qw�q;�ol����6����&����2�j�h�#՞�I^."��9��y���ӞF�5|�R�Ж�/E3�����hZV�m��!���%1�n������[�h��'ɐ��֠��GιX*H�R�w���]m<52Px��ސ6p��^������6���`h}h��!fA����V;�{��ǹ�f4[:)6lS��ê��w��\j&�9CT��:��6��*���0�$5��M�؉��0�yF)��B�Vn���I�!��"'�vS�d�?��]��ܤ�Π�h� ���.Ns�����}��eN'�S瑋HǶ�K���@3�MR�"���3�H���`Ox
��)�$۶����Ms&��+L��z���E��Q�C޾�ut���?.�6��I�d�F0�\�fs1���4��:l�7��rA�ՊHC�J?A�roJ�25��&�5s�/���)�����������q�}A��q�l�5�܉�+5��T��\2ι3���!������^(��N���Á�hƚ�l82�F���V�2��oĤr��Bp�c~y�r�دU<���7��������s{ϑn\���ɛj�O�rb���Bl{�;Z3�zl������z��^I�:*а�Xjן�^�Ex���lr���X�IZ�����"R��莮>�P
1�6[���[jA����p*����j��˒.$�n�q �%��	�[���7��֣o֫���]\�1����������p����,�[3�c�ϻQ��	�k�+hc=e�z��0J�����Rp9����oj��:��ժgH�ni�{�ל��G�����Hƺ�hˁ�!����з��ᐾ}��a&P!�\)E�\
��R�):	��[����ܪW]h	����_�Dɨ��-YR'���G�nk�u����enp�ϝD���/k"ڰ��K�ٖW�7L,�+��)'�NH\>����TQ�dH䆹D�w�7R&�:@��H�/j�_�h	��4Z JICZ�ћ�8u��[y���Ez�z�����8"2v�yj��/eВ��ch�q�x�-�.I���Θ�E�Y���栻�?�խV<�.WdD�J�`�Ө�j#$����em�.l&���[	n�Kkp�^�S�ڃ�����W[eSt�5	��lu�q�J��v챲Ђ������Kc������Ͳ:���5�iO�J�X3E��8� :�m�}krl