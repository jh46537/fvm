��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�-No�?�j:C�]�;���cu���uw��^&��YſYߥP�膜��9|��C|b�h&�i|�bF�L�O��_JĲ����+}	"��s�h�SuW�Œ�I5+F�N���{LK�ɔw=М�XR��GO�>
Ʃ@		�W�K��|ƀ9hq�(Uj��DXW9��)����=yag�+D�79Sp���.�!@0;��U�������ġ�J�B~��A^����~Z��a�W]��Sh�+�!������Ja ���O��rm�����u�/��#U�s��*�P�a�>��d��$���%�,��jc�u,sH<�J; �pˌ���ٮ?AB�rxƺ�(��#t�dE���X�	Aĭ%�lW�U(���WQ��B���э&`��J���h�[I#�˶Qf�س�#�I���ΔU;���2��k)[��e��sC����Bk�Е�٪oC�3�Ц� 0��z^���'M����{f)����Yg��^��������ȹl�I�i����@��07���u�y��m����]��O���.�'н���+����b��Cc<�pXW���8�2��[�ڡ?Ye�E]����tے���(���z��o���p��V�sn��,rbL��(�hG�5�#�tٞ|���R�`I�ݓ���M>�.�9}���T�Fg�^�'�U�LT����"��덏��5#.�u^�����fF����/-��( ��R)z��9���vQ�x�t-`��ک��k�y?4g_���&�_g����SҺ��#�_����_йY�5,�Lg��`���P��C3��c�����閊�&��l[udZ̥m���'樀 ��-�'Zb�μN	+�ɼd���ǡv��V�GRP�\磕���C;��]~9sQ�f�r�ك�{���F<E�cA[p&��/�l)�9f����e��ƒ+���Q��@�= �j�w�L��i���<��6�@�����\���6�H��R�}E��xq��\W�	A gН��sXn"I�¼���Lk�H�-帨�(�Տu!��+ '7)��x#+�g�N���F�y���:r����(��c�W��@�����s�r׵aC�2ܺ�>V-'��
A��۬��4ab�S�rkw��� OP�Fd�ꚸ'}���Gr�u#��~e�(��#L�hA6���yR�O=E�,�}�S$�w�o�o�z ʖh��Td���q�V�G�ؽ�d�L\2�@`�m��	M$��w�1�n�c���ڵPV#m�� 0J� 0l^�j4�a����9̶��Jc�
v�5���D*]
#-���Kj��p3�	HmFÍ�����l� 4��i9, ��sE�D�0�L&#�[^���;���B��0U[�����)���Tֳ
F��m^hu�Y(8�G1[�Zi��x�1p.mJ�����0�^j?�Ų�rm��Ń.�����۶=��	_���3U!����^�	HUN;U��՟�W���!�O�\���>����|Q4��D}�(���W�*ǝ�ޑ)��x�����t�T�4y>�f q��0�Z�<��4�L#9���T��+ =�b}���:�t��7�1����� ���P3r&c�EB�b�rzU�����X-n��1{\�CW�?�<��m�u�'�^n�я�`�c��#��p��e��=�
�zwG���ؖ�ab�BJK�]�>^�rX�%�BQtC��hA_ƗȖ�l�4J<6,��Yl{����!�%	=�E����yh ?��R2�VO7��i5�v��Ӷc���8P?�"L�uǿ:�uU�y��N�/�����{��MLd�ul��{�	���_U��j�=ZA쨶�+�"R���D	��	�jG$��d���x/͒fHI� �f�w:!uQ�����)���k9���3
�ٓ�V���m�;�hҵ[M�%?��_8*�1O�K�Ñ����D���ztOo�`҆)X L���t������8�ϲ�D��D�GP��PNN6�P�(x~k��q�O�$8�4��ҩ�Hi�H��hE<ʣ~��N�W���Χ\rȏ�g�'&��^�n�|kD�Y����)�,��z���wʄ;��@AQ��Z*�/~|@&ܨ�{�|�ݳ��I��b��tК}'��,b�����