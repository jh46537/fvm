// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:26 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fn9hepHoXdlMQP2pZf69R5O/Ty5A8TxW17CnUD3LfwVGVsQaHdB85KiO9AVlvHf6
/jRF0dOQwvYh1em6HA9h21fMGCxCOT6jqWDSJWwWfmbZpEJGTl4rkTk16U0hls3y
wrc8eLuNZowjZtJQlIIJhx+QvmdNpKUP+SR928R4OlE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2320)
zkWOa4VRExqade8EwQJxEUcj446Sa5yNHjEhoR0m9e1tnIWWAl6pvnsVFjVR1nYd
h1Q3IwpL1qvbIEM53rZlH/z70Lns5nT/rfLESLvWTc+a9aIER7Ar4O1q12LbgsRA
GO9FXC0Zcyi2YyAi0GR+VAsTJ3B9FrfcxPkBEbjuUh07EDQz9GYCXV4QtVyHLiA/
BHhplSADgtPMhheku5eKnydlSaYSR9ckXkF/Ro7WDzR9zios5v8s1qlwznSrsQwM
x6qo0BVLAHAhdxCudUZR+cCakW/8KtfiKwwMKKa/pt3ZSQwxVzIMDTQll1HX6Dit
kV54Cjkqb101Jgh9OJseALNnAPQejP1XxUTJVBB4n0G9gMa8owTRqKw/TnSr9LKn
sQP4y75sy9lNs6DWpS00n1ZyPIwoxnFj3509Zv9T8omIwya5Hci7ej5bHMxE7Wvr
hCC9+lv7cBNp3hz0YPF3xtqy/mOv7v4EY2H/bVr6UB2LYVCSM/sTtol8p69d7/rZ
RtggU21LRt4Da76apBATNU3NXL/+EsvkOCpTOyEnnl5mBgbX3hrFFkFMuC583Nmu
x4nYKf2cM7FM8ZrNGIkfuUDlsAVthQDIcIXPK/Y96cnJRV8hvB0lbIaUXwAj3cnR
NbcdPRlszSIhWzOzjYxz1gRP6DW76O3thKNwJoUywLj/Qbh3Acux5MIFgKr66FU/
l22wwPIka2QWNtezBkJaHkC2uKPGQ7yNT43b8bZxkincPQ+6cJXWNuVCkF6IHHma
OMPL3KM+85nCXdjGMplC5saiPz9uZ2TMuQRGP0+rCm9FCSGMLOckUwGDCoH0XuRw
YeaDmF9tCWIUZu/zMESg2uzBjCVlVEv3p+1CExLAY7bh1zWleztgV2fiD1NoWHn9
IyXJ/gbPpc0NI/ZxY6kExaDim8eVXZTphOT/w6BIQtXwRHVtckeK2HgsynOHe7m9
FjsBkQ042ITo8k51R4CzJtlTjb6HktNHrezs+OAxyD0L1cd7qWIZvGtQk9Iq2Vig
YX68ju182wCcblilBcilsKtjtEPTjL6uC8Y6gT1dGx8jFB8CZCouDH7nxhFhh69F
kkU5mgVzhgMRUVJs/28GGWdF/i4LiLBgYEfSgONJgoMv/+6/73N45uuA9yaWhgdD
3m6jAk0/T2KzURyF6APDrQroB0JcFjtjAYNVMgI2WXmoSpTi8Mk3chZCzDRE/0eq
K72iUdYFghNFVPoijBkzpUYspn4sNQhjm9KkyxVamAtpytovvOmIYQmyCgTS/elO
28/aAvXta2v+zSG4yO6XLEh8zbQSVqTnalS1WaQM18Zx12BYpAmm6URI1cXfeDYN
pp65Me8PT+xsc3QhswHAgsWpQ8yradkrycPZ0Pzx54w0qdUB9KyrmJitYGV0OayO
RHzuoJNEenRKJN9peaKIKbBkmqUKbtnVGlxCwMx4ocDYchI9/wGBQo5B+9lv2Ge7
0DQrWis/r2suGAtW2Z4vXNVmq57LxDdrM/tXp1wktmvly9hjRnu5l6hxi5TCIrly
NknsW6Iy1DljprdTU8Q8NEL14UqrgleT2Ojfoqz9YF7XvNtTBzO5es5TYPY8gmJw
aq5tDE9oxdLayGm2DS37Zkm+glH8z9m9YKEO4X5/Si9At/xldtMYGPl+4lq7yYqx
cfqOMbzQUMmMEz4O1DNhUcfujcWcDdS6bvjvRp3qkpwu7AhxB3+ZIDPHRipaj+Iv
NA3+6uMSzsJEW/y9RYMnyuvUJayJlQs2lDItjDpSj2h4CQK/l6y6fa0bKxuBhMaR
WZIqnmh9Raxy2kOhnb1sHJZI3AluT9KiSsM+JtrJB+ZjSSbo0VhBtvoTi3lIZxoH
HCnlM1jCZCEyqqVrR86fQ+g1DxD3SXelwkM/vnm7YrxaUT77O+OkUKF0qf1BRSMg
D6XRYCUxaxEhFj4WxbpZamTiZz8/lJaFs2aQ8ry1khXm+wOGhmRRhUH2g/QVgEnC
ennZ5CyU6chrd1qNYT+p0gYix56HEDbt4cyjBcWgtS46blSrbdL5jT/3ovUUgxNt
RuqgmOnIqvojwK5ArrORP0AFK7lQVXe40uo11UwnnfBDLlPgw168MRv3SOxEcblK
CiH5DP/j0hGVMoS9Z3RrWIry9Y8sKiFg3XACXV3qwrjOcV+zdnb8Soc6rwI9nrPl
+ePFWnTOSKdLSG2QIB/8P2pFj8L7u4XVZoP8nruA9zkL+VNakCkcgKLtr9EbZc4j
d+DCKzef/nPAdQWG95LCnwM+l8AmIogLH6NwbYavtLPKlSTwLSfnSOhhfLNeEbvK
3ykA0AxZdpcypO3nwFHg6XoksfmvYRBXhwidJM1Ih3Q8ezoohTZEQN+kr5/HUiJn
eixZSn2kb3IMTNos8qMjZ41es+R1xO74y/iEJ7wAUG2eWJSe+76sAkDNlRSlRwAi
GFQKSeA8dIg7GH4v/DrNTDyB37zC2kEp8wptmMK28J9tiai9Wl5dVKBPIXZvuegL
+wBaskN7GtdPzfbwsJnHReFhhCxYJ86Hujz8f4LRE5d8uCiAkgTaxdyGNzpiIKR4
8Z59e74QSexCU9LWu50awWDLdiJqDF+1sE6s+RweT3GbPnSnCRfmG6ZwoxArCYrL
qwMM61ATpREjHvuOZLiuYehS6+11hbUaM7Hef8FUskb2NUAqDqJO/nAq9HyfbCgr
ILQaZXnB0bXHQhtU6L5SZQ+hM3v/AsASI1ncBtDWBZXxyICuWQxfd0iS8kVLe8u4
4fPlNJrxZOTJwPppTLpHi/hH9xdT3VRJXUxq8QNU+yDYssnYp4WXEBhAUK+X6Eis
2WTKLEpr1QdT7QW4UXwLAKSplXW7vEWBUKXZalV2ryWDyB5PzHx7y/YXgq1ajTKf
d8YohCLtX0YHvneFOLSPcKKsCrd0ljImfs4Zb1KQXPaOcsT53QRV9QsFGDwCrVjt
WdAT1FPbE09qipvyuHJU8hF6IkZoDS5Tkd8ScV6DfHY3eN0yOuX5nEDeWlw3NW/V
+D+OxP8ky9SJPj9nxo6mNxHDc+PV/0Y6hiTMWV3sHMDGFCng+khcxME5gUOlvRRm
re4+7A5hv1/xSUr8jijqaA==
`pragma protect end_protected
