��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��<���A�_\�����F��ߍ��l��Z ��%�����
�֑�wj��}1f(�t\z�3K~`B��ł�$/E_���򴁛�����J �7�����o��%&�1w��Q�	���U95�`ru=5�8|��a�m�X']�N}pKb@��"�:�.�x��g|Eo@@��t2��T!'�O,&6���Ց�,%B�G�S�ҥ-�(����1/f��f4�p#�C�rlrd�#�hv�u]�ьR)OI�n��-��07��^��#�B���r(My�#_S%�HZ!~t����{��6��]�~�x>��|���n��"��m�~�������i��4�_���$o�d9KnO�&�_�m�\�����IK�@���^�]C3������`k�3��0pF�z�h���J���r�!���Ue����!���m#��WJ�!��Pѥ��Lh7�^��#\�<���� ��0�u���Ng���c<u��1 ޵ ��+�i��,��_�����z\���!��(n۰�H�7���9�v\P:#����q�1&|�
v@������'��� ���������«����3�+��ݧ�Mm6_[�P�#��1c8Q�T0(��z�@���R��'n~����%^��J�,�$�K]d\M��9����~^�w �RI�A�LSp� �	,��AD��j	��ޛ�PIq�O@'��"�*��j�jP2�p���<��x�� /�zy�I�2�᪜@�]�mڻ.P�)����Z�|��#�$g*�H�]��6�kU~<��l�ŕ��`�9���b��p�zǫF���A$��+♆y���2����n=SS~�l��=�>d4e����P��OИ������z��Z�#]�9����ՅZ^IU\OGgxu��-�{�� 7�$oIIJ�|Y2U)P�����4�./��j���g`�u�t{c�%B��پ�[+8�\�^QG�V��Ft��D'UNA������b���H
R������Yv.\�W������я;[�ڰ,� s��A�|1�/Eh�	�D�e�F�Ϲ��uy�r�����M3��tc5�����uUf@y/S�'�h�� P��O�V<���ŏr�xRJ-܄e�X;@A����)�<�<�Uœ�%�V��ܻ/cF:>*���%#���A[KR�(�qj�Vd�n��#��H9xs��p���9��ϓ�"��,�l�ج�O�9I>q�4��	�A)�G7�d�֞���Q9�|p�yQ�u�J73Si�6X�dQ�~����0!����j��5�J�t�`��N�^c<:8g�Hờ�aX,���>t<����\w�#b~�F�����̰^�#�x!�w'^R&LT0[bSE��*8���%�q��ϕ/����\�-w>�f6&����n)�^�U�(E��%����Y������c�5dkV�L̜���/	���D����[��3�p�L�tH|u��n���H6���"d*R�ӱ�)���/�"CК�	�tbPv(�L<�t(Q���a�ޓ�Qt�Pg濋8���  �>����hVd����s���r/O�/��Ȱ<���j:sN�G't����T��&̡|+�gC�_�8��tpz.0���������f�Fq�#xo��5�P{w��_�����ּ����b�1��`�E��wB�5M�2����d��y +�Z���,MLB+������'YJ!?C�[
��#���ڵ���	�ў�ܳk�	!}�%�t�Q�7��mw�u��٤�,{A�`<��剧?��҉�k��}h��sK,y��?캇�-�Ռ!�=I�d�>��̝
�3�{�j���c	������%�������hw�J(&�POI�R�/ߍp5�y����wmW��&��Ű��L��y���'�k]9���L��@u�NN�`ޝ�����I1cҷ��!��]Y��Bg��O����_;�,g���y�ojG�2]d��Uy��k�PIR�o�/`GZZ=�_�
-��Q�
�N���d�w�;373�~n�2=��V�㘃�a�����=R�Z�##��U��������/����Y�z R�=��.��x����+0�^�_g�'��&'��}���道m�A.�\ӓՆp[��$'z���K3œ��ˁOD}E<ܾ����I�����^���wj"���H���K�Z��%'�֯s�ܙ�s[�䷻&(kX�Tmc� �4�U����@%u�e9	�};��VinC`���+�@u�8��������щ�[C��k�]��%�ʇxs�R=���V�_��Kf�Mv����&�Z^��l������;LK����8-ȯ�n ��Buj�[bl�}�[_��.粰�_Ml��5�^Y[�	�t��(��td+��Ƹa�*��W)�ٮ�T��r�9$$Y;Pc9��y=q��O��)8������"�-	E�\�n��TN�8_Y��G�z>��m��,��'�"��O��Z+�A�T��R���@�y�V�;�y��j�b��P����B��q�`�!z���l�m��X��\�#OT6W��Wť���ѐ���#F �'x�a�&�s��q�7�g6*Gegm�����ֈ;Ԁ9�	.�M�x���0A5]D��L�o.cLN�e��Ŵ�bL�߿�!}�w�I A�/+D�ɯq�](G6g?VF��'��J�;�C��/q�\��r��VY2��rK����Tñ���݉�r<�VǼr��3��YY�NT�K�i?3���)G�F�^�`���@v�;���6,�|g�/�����.�\�4��γQ��_g��"J���P<6�� ;��j���i��&��F2]u�v���]e�t��Z��ڭ��}�~����a2��l�xW��Q�A�f��>��(�z���2 �}@�˨�3T"C��;Ͳ�B�-I�X'�2z��ˡV������qcA���kz�I�a���1�ք���c�Boc�M[�� ��~��{�.j�5��db��=����s���.���_�~��	��bVk5�e@�(y��T���Sn��lN�ސ�&gM�s���4�8l���[W��]ƾ���z{Ov&W���O�+�Z-��	�sZ��&E�V~��뉏�O7��;�Oi���D�{C���B���J�2E ����KǙ\:,yߙN��������
�H�e*vFy��o@��x^ Af���J(�w��2V�@��1�~�9K%( /x�ᶏ�Rz��Au��ɣ:
���h�i�\��s4�]�S~ul4�N�t]\��n%�����7dTϲ�M*��Ή��D7uN�u��'������cAZ:�{h�r�d���\��\��L��3�=:�9�����R�2�rN~k�f���*�7S�[p6��A%��E�2ۈ��cf��F���#�ܾ����ã�^]_B���Ć�W��$i�}��*�j�~ �c����Kuxc������'���pE�\�ϮoS� �[�@׻�S3�Ba�ӼC7�#�c�LX�ȣͨ
�#��l����ʚrT�>���O��I���5�S�MF�5y�׻߆�/R�#^��q�@�H�!�tx�7�OR'k�����'��,	S��Z~w;�b�m%���ZPk1�}�`H�a���D�����u����Mz��C��^��p�;�.<���\�U�_�X^�gl2,��wQ)���w}�'
�s1��l5��us��zw�\-�����:0Z��@�����"et��Vp�g�����0�ۻEb�o���e(��h؍k�;�B�\F>4�;�� �F�j@	J$z	Q�<����VLRTASO�9�G�X
���j�U�W
�;g��7?�sݘ�o!'�\0E�fm
��J���L!��_*Ȟ�t��!��t~��{0��a��ߑ_n�c���S�此����nD����d���py�_����|i��{���s��3$���Z���[A���]��PY�u�2_��<����s�@�jh��^.��<i�n��l�x��S��n�%t�����-y��s;;��͵�C���	g=�� !�p�PZP�~�cБs�KB|�	���d����`�@����x�XS;��!U����H`�����.���j��Lu��n*��*��ɤ�*�ej�_���S�q�YLQ>;���J�+P�mD
T��x��6{�,�|��2@1!�C]�),x�ڋ����b�|{�SR$g�)ūf����?��b1�=�$�E�����9,�(�����IV
��'��6����OU.P��4OvF��!X�;\*x���a�*^J����7���ѻ>��0��hC�����!�M���������Zq6�y�s�z��J��y�r���۳��g�h��R�F\�"�@-
V�LX��Fʵ���o8>j;��� 
WI�4�,ly���4���n�F�@�<�Q�ָ��1�pfh��f�c�e��0k�W"H^|^��!v�Ţх{��߀�C��V*ڄ�ϛpcéD��5��I��˳4�Dm��PKk$6����$�nr�(���Y��J"C*��,PD�pO�C$>�1h���0C׎:����;�2ۿި,=Ht��z��6�hL
SZ�dl�����ʿz}Wt�V�z��;p���4�l}}b���}���<���Ƴ�9 ���1E����3�@d�_�1:<.L���x��f���4X�?(�� �����T�P/�����l�7�l�c�K}b�B�᪭#bv�����ɫ�,��@���.��aq�5�q�a�������M <����b���7J#���o<��B���i�\�NeKo�S_�
K�a���q�������Q�&�D��I2�ϔTm�❲N��KQ�
���.��SP��
F+7�ͭs�k�8��GcKsPwz{٤�h�y<U�G�]��%p���<��_%k�>>K��(����c�gF$^�qE�My�&}A�7�LR��EjkW��r��D��k����D,ʑHD����䩰Z�&�}��x���N���
2-�ˆX��.~�U��+��_"�	�QL R��oh���0X�/6�6��C�ө���j�2- �ߍG����ȫ|S��c�(i���y�FuA�/��	]SiW���(���Qs��sʾ9����5�Y�+�1���NlM��vR`�3�A�`u���wΒ��M�c�4��!+s�}���EyF�T�g�h9�h]�?铰��(+����:�T��B�O�5�A�d��&��1^����6ۭ-�5��!�I���T��V�������01ڳ5������j��@���؋��zd��`p��a��R_`�@& :�]}?{˽G����|+І7��K�g��N�YA�Lw�v\�� m�<� �o��k�����bQ-���X��SrƖ8*�2X7@�Ϟ���{7��J	?䝂����3�S�o�*����~�θ)y�v/�^�����[#�V�n�UE���x"Шyl���O��S�с������~��TH�M�å��;z~*��L���y��N�X��wN&nB~�N���oT�dMd��W�9���)k�7�Dߌ����>U����YI�WCDIV��9zPy��9F#��>tcP�CSJT4���}�m�KZ�xw�ҋa,xx�OGοC�@�ە��!b���!H��	8��d�Ύ�z�{���#�tp�Q��e/�q��q�q!�6F�8�č쒕��T4E�3�K�n�L�v8�ۀ���oN����)��R}��|x�*��>�1������@��L�BT^nT{�t.l�ĶyA�������G�8��K�E�C`g�T"����Hg!3S^��z| 0_�.��M�.�^��M��_��ȯ���O�=kF|�1�a�I�^m��Gk�W�)���!JO�I�[f�r;ۼ��ң6�Y�2Y+�ϊe�,m���LgH�I��ݫ�� f�"�l�r�_�<���B{����[�0�c�k����;��!&�M��h �#�-�-�I� ��YY���"�7K}G��1?��>��%�_c�����Z��FH�7�L��^?�}�/�>�a���#0�4|,�ƃo��u�]Ԁݘ����ofzFv?�S��染���(�lIL翰�j�U `Y��́��]��1�%J6$!����W�������=8�l}H���-�G,a��uϸ�#F�j�W,�1�H4���yP�&d-SZzѵo��#l�t��H/keD�L��uk��A��+E�	�y���C���0U�qu�G��@�
�P=�yw�ڷ�Po�~2����5F2��S����OU}�z��'��f}��a/��ם)K�G�]�m�Qټ}A���ۼ�[X=2)"]E��Y��L�a��"�����QA�My���z�oާ���NT���R��������vF�����Ǝ�^!���G�¼�w�xR��u_[��26�O�U�AFh�-���Ք4�y�z�$���xd$,��������,@��R�\����(P���<g�c��b�����H)���ELe��(��u�.��<E�ř,G�$��W3N~��^���d��ZuP�s�N?� �EK��×���K���q>S	ŖhJ���x��Ǣk������^��:�G֩#`4B�Z�=�!�n)mx?{����es�����m�	���ѵ}x�D�\��[����t%���xk�W�ժ��Q%����4�����6�m)<2�8<�u���ǳ�G�iH�_m�z��y�a�1pxFO|+;�<[�/Y���ֆ�7�tվ��� �G�d1��삻��D4L&���x)|sNک���ŋ���m��@�xS�V@c�g�V�wy��5_9��?s�u�e8{�\�m���Ĥ��k�U@�#2��K���_�YK<�Ӧ��Sj�����-�[�����>�}ݳ��k�$�am��h�Z*�v�0�3����2B�~e"_��+�F�Ѓ�E�����;����.e��I~> �s\)��{�����*�TY�p����oF����+����"ԝ�5���K��.?_o�w���;n���nL�*�N0���0�n�����/9So�v�=p�o^���ͳ�>�}���_qs͂�&�0��{'��9��0�N��҉�J[�ȩ�i!Y������12�с->R.}F8uƭ7| �@4-`l5�艸F��r��/�3$Z�yGp�I�v�� ����,����9�~�!����;p��C8��eC�� ��T���];z�D��0@��;��K~!��	a��� ��,��[	���<�M��,��#}�߶4��?aZX�_�/�/�~R�l�hG5܈���ƙg%*��D��ým���Ͻ�H �Q#���9��A<�s���\��߽����7�S���/GH��>�g��&Zw[hUw7��Ez��\���VT_]E���#T�r}x��P�2�'�I4 ������[���f��I��KE"$��[���G��z�i���.h2GnoL��Ֆ O;�����v��u����%k���l�^���7���U���h3�.�j�ϫd��cz�V�஢��`��0���&8����{O�=ݱA���nّ/�u\z,��o��Z�����h[h��֊�d�+Z�����u�]Ճ�_�������]~#�B�����f�~wTU��ۧ���E��\(�YMC-B��sO1��z��"R2��N�tj��IJ��l�j�^R_��,W�����[��Jxڮv�<�g���W���7sI{��j�:^�Z�������f2��fƄ���ԉ)���5��e��Q��:h_d����;���G�>��w_~g�R���O�dF��2U-={���V)���S,g��w!ڼ�3��z���t�SE�h�V0��򃣹��3\Ԏ&���wpQg�$�\j���0t3X<���俛؄5iB��B��eU���
rK�V��$�m��]�:�L�2Yٱ��/���E5�5g��c��r'������1��y���$�?S��h��?��aVC5���=��=F��vE�8��9R ����_�&%�n,�MYK�K����e���E�[:�њs�����C,9�m�KH���]�r�\�����/��A��