// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:26 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gJuoznfF0oRsYI9mho9QbBF+F29yq18E9sKY1t/CqTvu12WSktsDj/M0ALOOxdPJ
0QEQ/auCJthOv5KfmHSKOu/q38DLGJGaRXfTIbTuyb4Ddi4aIxT7mNqVt2q+RGSH
Z0ekKyrFsTlKLLTcmiK0xujOjFSvSaDHgAC8qhu1aNY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13312)
UoWhrm6Blh1txiIdvioV2+oNjroiDaxzx1oYanK7uzBcuFHtuwtidTktYtVhPAbx
v+TWbBBScSFpdpuoE94nnL77z0KgzReKS+9gJdTrSz4iwxtE2i+KOoQ0ZC1HxJ2D
gqogrmQlqHMuLcx1XPkc0ffxgV+f6JNN6OwDUHS/EqEDFrygw5D1+r/gejOmWwBm
rihG9Tkb9kj/+OOmwS2qvji5A2jIxzy2mJOA/wwTaBbNsyYfzLZPGBQVzhxJg3Sl
Assx9/lwba0+F7Oz0yhA3uVaZxo0PqBFJ0fFUEp/hT4Pu8pM/LW31m5GAUwOW/Vc
QMnOjWT2sQuBhTqVz4WYW5eBziwSPvuEgGgWgVCiN4vO2m5/oHwsLAUmvoo7FvjE
2OatH3503cw24bcz815f1z6H5o8dkze8QnTOvxvY4GbTTOFs2ufNwS7T87nSdutQ
5GBIvSkCqLUeyGtCCStoVexWHpXF8pXzdWn9yzJpJh4+3lclN6dKu14FHzE5vwN0
NzGvWWZZ9yj7rlaEN7Qd1G2CNpAPzWIzTGtS6PDHzBqrpAxGWe6Jk9vwpyOnwTlm
1Ow44r5+Sxk9sSdnbBvhg5rmhgVJm/mj8zkfW9ZmQsZ1dcn6vfLqS80T7K5d1leN
5xk8KWhsujRj9bQhtju5NCKf6TahS/KDosGqRhuwTwz9Vb8G3MfbT44zbqkNHl96
094n5R70wmRv6X0fAgWReGs3GdqJeh+WUvvGWN4JYlvxt5hxIMXqSedOHv5cmMew
DU4Ywc6Rh9o8amI/Pe8oQ+mk+DbUg4+gKreAQ5wz+CyWBS8kYxtJo2Sot1FTuPpb
OUKx9zdQZxXcH/BASBgi+elSPaaZyydck5UfHHb0Lu0e97MITY5emB1nUkD4+pku
ly5UWEqwgxP/zNdnf4jpwamOgThsmGyNh155veDNWhQxkUN82vguHCU5I22sucfS
WHMw3EAXfJPiGHHiqjUGwNVYdICXeDAwKXOjo7riNa/FW/nlDmdMyboJwjv38Vnm
qg3OhXBZR8j46KjFgvYre1TD+/U65M0lycW0uSLRucjIe46jB6/eFdvq5TSoTOQU
IX+ZOkr31Y214NEN3jgO6JDtJVJrUH0ebIf4+K74qc12Y/GcPyjaH5Ji/3p3vOzQ
RzG5oQS4FgBLH3rbp6ewMbiyEZi1HMC0BOVvPTmwE/O6tDyBeo2z54lV309CSQFw
EzhLtrZjsDbAAH4acqleOCPYUpSwiB3HahXaIWToSs7W/HmwkKYfGZNCQ1v6sE/4
O3GGI/CaxzKU/SH7+NpsiMCD/fIXeij6v1cAca6DUBTTxKic6345SCcogVEOY1mN
fVTwHkrXmDp5eG05N2q4WZ3EdiDemcrlIrpqJwzRA6sBNKfM7Coxas2/CPuk9TcK
oqP/CxsdRAWBLxVVMMmBzncVubggxIK7gjwMQHp1j9XU0JtIXHg3VtzDFT+qPndY
6Dcka8AfKD8ClZ3j9h65z7E3K6IKGZVGiFOrp0va/V81o2uU/cUO4HuqDtdGT6ko
r4+laITjlZXCngtnV98JnK0BE1wT7i4vuytMK4RokklwizDjMvFt+SKEp3n7Hdvf
KA8Q0azW0wfMRm9RQJ/Ripab4mbqKBXlf6fZ7PlBntM1AWHzuyoKNcnQCM0GqVqC
Kfp7UHSLlNKscEDEoLYXRSjkQlCs71M8sdWRE/iRU4c9/VcH01bisuppxw24JHIQ
lJ8v3WW6IbJCSdsNxx85CaF7I69ERry0A1RkRLcwwVoZl6RavPBVcol27YdigxVP
ezfpExT9chxfxlUcH6ByH/hbz8Rb0nvPShcF43MWmGksOeFUCJYgxhT2F+c8Hxbr
lUJ5PkuMZybZgetsMB8gydLXeFuhiiCi7kugayueO4SrrX6Ri4JpNYEnYeYA/yGW
BIb2VjmdiMpJ22tKAtpB4e8XzpDsII3/ZEY7DpaBLLqPvmfnWH9Vp0L9uyej0v/k
EhfnsdSI4t0E+NsnceFJtV1GWGTvZIEiIgWV0uR6PU3pQD7cZQsQ0jlMwA/YR7Sh
dMHLDVOLP4Di8eXaFCfcNuHpWuQs6Fm8QLhKbIbUwvded5Ycltg3TqVAj1M4jb7E
hfZq93vEKax3uCZkdlT1jQvsPgB3uwhztD6FiUvFragFHO8wX982hj10ByE1Hczs
V5W9n2G2gEMPWEwRqKoA9AYH7EFmn2r6QJMGukkcMQ/6U1evc5+FKiu90QKDNNjC
XQUGgxCA2hLfE9SL8wdnjYMjOFaOP5sQQVlyvk4EZBfGD2q0zvZFO9xwxIjh/vuB
THWZf91GhXdrp756PiWH9vQy0kWmSQWPLMkmhKPMaW4h4EGZrvPiaKKfVhwUrk+M
5ZLqTa86uo8gdi8Ju5tXl7W710qMnwDVdM6wgFYtaC6PbYqUDtJIniTAwEgqozfB
HFLVsktIKlTW4+YZrXMeNLdsU8NvqgaBcj8hlLgjnviOD5OdJBao6KnNQg9xMO9Q
iM5xRbdl7iKA3kVNg2VJkV+THvVdC+BxzFo+BnC1aDBJi3RIfg6voIRor4ilJdrE
mMky4ntgiyszj30MjQuJqCwPnPJ1aqmx9O8Qw956P92xZJT6n3Ur8o/apvBLW/Cv
MmHuLwcMGBbkwd+qo9Jf/XfTIuo6rfwdm9TiS1C8H/sDKv4LeRNDCM1oJrSr9u2S
4zYcgIFrfNXGspBBdZrC6ezil3A1LCGAkRxkPs3NXOr7eDCljD64QURDZygnF9p6
35TtAXC5GWT3+JVhx5b5KaFeZzNhi/WjojB9wnebaszF2BL7WmZFXfzqjKIj+RK7
ULUHZaEfPlrmSHU1cMyh57/mvq+MhFjitamlEBqT6iC86ZVbwVani4XihCY/2btn
1MQbOx58+FQ17AW2qPCExGVXJU4mYY8sLX1Kjxli0T9cNdOsqjQaeighi8YBGUCr
XHpSrFQSIabGLVUOguFO5lj67DRmXCaKSvOUwi0eUv8XsDt9z8VfwQk4Yt72Qr7H
P2opl/qHw5B8pkP4Ac6dXXsYVKa4iaGRmFeQgaLYNoiFTULLpHWau2TjyfOCM2DR
k6Bv9I3gnvQnXN1sscuP629m0XE9pRiS7lkFtJ/oPi/Dm5rLpULzpzftx5gSMla5
xIGAkf+YNWG9j2kXJl2e7pcukSiXKLl7zYAKKQ68uk/L9LYJtqCxas/PgikRYAF4
41M2IB3HBOMvzubr0kpW8huEWCkX1So7KksQ7lCYW78YCBcf/DvE2SqrUuZbdvmC
0tq+bpsmwggtzlbqe6I81+2X6UxQOWZSN8H34AduZGixK7wz6aOJ3qWeOvAtmCKy
+/1iA6L/c0LbEljnVOk9pgbsgvKlzteDy+kcwrJN/bMS29E64PneNnr+up+Yh4B/
MaXM+UIoGZnvALhf5VqXug4j5RqeI3XuXAcL+AZTjshKVMwKQmGnDKaqy4uW6L/P
6lPiBTfMtwGSYXTqsEHXyJSLigECE9EOmDfAH72oUc96WIk2NKmB80jsGDjK3lI+
RpugVnp7AVcgyDqFwxKypqD6qpU2FQLZaSDzSiK4llM91XhwfEh+m7IS6roYZZvV
NmDwZRAtMa1Di8V/TDShtjRsNEeyB9YJQ/h7FjnYuJG2/RSjiit+16SVsPzChCM5
pIknqeqdGBiJsyK5XHkwfAHho7MdhA8WlAm7Mw1bBlj+jG0TW0c1d8sFAu5W+8Ry
CtdWdJ0fsl3LyXeB4SnMC7zpR2GsflGhPdUXjrFoeTaH9VLCtgGBHsENeUgPcq7O
MfDj7US4FhhLgWY7bariNM3/MW0KDHNExfl2Gixc+CzhKrLLQsg+2CYBQ77cnKHT
BBmKtT0FRYEf9v4/jGtxbNFfpZonY6+F8jv79Ab3r157ObALoo9iEBdulr5Eoybd
v3PH52QNc1cCdkh1F1RnOK5P9V9ZxQRcxgeZY7LxLySERxuUkY9BswpM231IIOt/
u9VjA2bsusTuQ7mHGXWmUTICY/qg6cAQx3pEZkSebFDNwloXOG4CiXEeXD5brf3I
DGH15NiCjdDBCKRkCqF5254FK1JTQGAfDxDUaOJ6TXXEVzsZZGadokN2DS2/VWHc
+7W1HGFABGCu1RfDcQCXzZwUR5HUqx8NIhLUPZq265/yJAmqv4YgGvV/+G8aAa/Q
DHXSpnh8pIBZmPW5CjP3oIVfno9PIZDGHrA32xSMLbrn0mhXG476FRdO6EMdBRJx
JYw8yaVEcHs87hBL/rMoI1RP92w9dJcOJqAgrkLpy+iAvHtcaSZiGNZG5dm1LieI
UzzPGkmneGULY2EhZv7hHbtxanSouT6DRP3BBw0UWiZ2aSmtfwxkCRdD2UOrfsel
6rbTh9R0fedOOGXoVHFq0fK8Ij4qcgaxUz4JU2tFe2qAqKtSE1+4cvF0eWSI4Y8n
M8+8PG3KQHjUdPS6MuIWvT/m0i3Uh4x/IC0swmexY/k2o7hf1ev21obSTkbMRhVK
Jno+SliS2T2w39Ks9zNfWjge8BqGjJmX61HWPiORj2lrtYHpaxN1tFtOyHd+WMCj
F7ohAGWcE2w05o4zJ2eETgDbTxcUV0US+P2lu2A6kQsD8vbCSK3hBE1jx2t0m7vD
pVS6IjVtJWglDT2FVTUrOPL1oLi4SvHKHkvQUYpUkiqUgfEUVypsms0E/o/DjQnF
63rqdDEVE+AbnA89MLvVP6XDpoaMPPOos+jBkhpQDEzdYj8XcHI+QFdUEZXMdi2g
eHP5SH2fVSwFn1KGUARLG6DCZ9zJ63XtufsViL1kEfZJc3f/MXou1E/B1u0GVgpY
ZteAR4alQDI8YnCr2Y7o3lcP0a5BFZPxqJDM0qbfoBV1i5vrghCo0uTUzzHJc2OO
LdVrtItMDCyaQKixAN5qtlWVwMloAziMOWkQjGRJMDQkfLnkBA8VYSqUxtdCbyBu
H50xYgfNWN+qAKiQULN925jJ2Fom/CIIqTOyru2ACJSagPXb7i9HJiyF/IFETfVh
EILOCR0Hld/FXJfzuL7aMvfFkzeeOLWFmCRWtz+zWuMxQK/JrUtOCmrEsjs3VNl3
ADcJVDf7Nm1ZyEzJMywrdfbhQw/qkRCi+TJr5TSM9fs0fS0iN7bvu3I3tZg1Eihj
nrp2HdnWYnePy3vOs6K+j4M29eBqDLPeJVFZG56VJiEyvmX/PZf1c6lvAaYcWwsD
eeIecsA/9GqeRy6fbEQw2tu7jMbCOVyVL+bMtfzFSGl0jTm22iZ40LEc0/1Wc7UF
W7FtYvOLVXwjqv7ZKlluZBd/8PelNTy+FPFYVa8feijzEj+rCNYKaZAxnOzbr0Hq
PCN13OnSKtnjdZiFlbSPOy7uTX8tRJLuYhgeKWh3ubjtiMxYwgsBMxNlaWGxLVcA
DzI0/RFQXJfw04Lq1xGIVvp30q7lX6GC8Z3jEhIY42f7Jqb5fULwb6UmvU36nOhD
whS03IkXYU2GU5nJXm1iUHArPqiXeytyFHFIaYy2EIZKq7xfZZ0mitBjCEe2z9uT
X5hF3javDWnq5gepTSqTuGhKMEG6JR7uydNqGlD5NCFexygHHe25W19l2RBZ4Tey
6HjiBaLFROgGHMep4poTz0SHM8jpn79KJogq2sSloSo6FSb8fvXyUqTJyXk/+7C+
ezYS2QI/RSyocSTrBM18/eIaTMdR3XAjXLsTjW3qfvnuXP5xCdqL/3DLJHYSWmF0
h358GNkLqNK1R+Le6iMHrg5FFg1rEgkR34+AUzRsXADO+aylXyFIabL+zuCPZe/W
SAHlaAwsLgkM8Yh/YiDEQHDLzBkZDsNKbgqUCLWzePGfe3d+ZK9VGS+gIHJ5Rirc
+wix5cU2BxiomE9IIPnGR/OeRevXteCEXCmJbWIOSzR82DM+ebK7ER8m343t/Wve
1diGvwHuVk0crrx7Nrbvj3dvG5sZY6T4XGv+N4Z2XSitXlWrrSExhoR+u+Wer6t7
MKynvs6Z46tbKirde8W1Dqoi7gdeLOcp/cFzSdmNdpXq5iMv0K4rTkd6Lz7d5HHN
LwOcAUrCBWU0Dm4GNM9wYm7EdPb6dLHRyIWgO4Dj0DBf1C+cdN263XOBnyunBUJz
LRXjbPk/yieyMD13gsQyx5dXuCrIYKYHZRW/QA+8eNjsQrQGLcd2yOU5lqHI1Ll/
cb7fST0/QhxKpNdsFFzdJzeXmuvzsfhezAG445QDLZvZFZ2aCwTJcYYdg9j1BdHx
Z3jRHAKlc/+oG0m7w23XWg8jyI7l1MH7q3c9XTMRuNeoAJxXgfKPaNOAP8HemMFA
1Bh6lYf9I9Y0o6FWoHwuqW+vAZ1HzgJ4EG8xlF/bVFFWn98IYD9nBLoCzDElRVzL
EONpoi7QrWJ9Hm3eD2TnOC9nDRppUHYpcvluNvPBy9S51Q1LhW1oDcBSDKS4lx1L
Pnwct15Gnp87I/tR7YBiP0fb1alzLmOH1OcE25eIGyLbfWTr2Sebd3aPOzHdCz3o
bJxA8tRorYQz+AeefIciPsRPsQqG8FTLhXosqOzcDxA/79m8SACR4+rtayqIqHTS
+9RMLXOJaQQinAnOoEmGYwrrkw29nyl5mZWQT0KZcafqXLsDnq47lNBm9Z9s51lI
qihj4QmcrZPWotPYLuRinxZYAy9Bla3ptiCSWOA/beUEZ4VhtvwS2G/pWzVUFfpF
5x7/4j49CxGKuyNqKTNA7+JoXwwI2+uKkV7ppfkCiZOqBVeFuLzdt2T72tAsauWJ
Jxmc++NU7DV31/KIG8nmmJZmvNxkYXr0bhX5SaNT1dZtmVkzppeJc5MZzlF0EGqB
IM4Sy1AK7QVHqP+0RvH0FCW3RT4e586MmV9GIL23PfQf4RoYZpvjYFWgur7pPoKv
u9rl/4c5d9ppadlMj2cEN6gaQvFJoAz1pp4DIBuSu8jGzwG90yFeHztC5hVcigjk
1LIJDnA7aSUXYTqSRjT+fYWJOQtR7pFMCZKYgUXdjTIuEkk90SZzvAInYU6jwJiN
BFfir9DE97Dykw9KH7Um5u2XjHv2G7oNKm67Vz4Z3y0EW6QAd9HUIEiVbb+yrVdJ
/+gxqDZ36V9mIrDVJ6Wcofm1saYNf7r3J78BmTJsFWhyKwVgegvat1C+TN7tF9Pw
AeXjuAOZKmgWBhlAf4HsyDBz8k8CEEn+08g67T3Lf3g8uebA5lZBHO5YM7ujYiBx
FiCeFZPRW+eEKuHQKv6gFCt5vxFP30GcLFqm2i0/CS+rBCNIasOFOaIn+PRuqCbs
jPGX65ftfGEZZTH6+qKi/uN4yiLsiBh1T8siY2FmcHO/qVICsyjpxADbBp1skNsq
U2IrguyrgkfaZ9j/DufaQX/MILsKh8g8G9nXQNkkQVIW0kaLKni8vpiK3TgHAiUk
rA+7DsQ++6tZ5S98e5umEaxE6u6odSyUJg0L01rK5AlDZJzvpkJz6QByyYp5FeK8
i6B5d2zWlufBv/pTsmf3qjCopsyPtuZ1fYTqamYJpmoU3pZk2eW3mF6JAl/bzBD4
6zztUAp9Y60o9w7JZtbdkG8wYoe6xBF88rwK5v7rNp5PtQn6RnPaPrUCEeekyctR
k7GNtLmyvGV7vwPAi+pOaxUABQ+M2/NDDEF7DhjWMhZQBfG06By+K0Upf7garUtl
MbgD+fHOj52Zr0OE1IZL8O8Sk3P4nD/nlD+4gFefaJXeN1Gr9N47EJ8XILrhiXaP
NVH9Vt+uyfNHpOJQJPslMJ5VS2WTlsmuJhh1OoCAw52vpwQ3mP80o1Ksh9xqc03i
vh8qfbjSTkrmBObQXJTbaEuUOtsG17wxM4/s6pZIzbTNnbjF988hUarK5hIXtato
SSuLqfGoOQalcCEw4LPzV+5oEs/4Btr4qNUBKEL+4npWZ72/uKHcifAFFTfhtPEz
pmKzS1ZC+yOEhjoFDBGiuqTSQKHjaldYFdFV9gzsl1iHLlVzyYV3eOw66gxCci48
F6RR6CiuwsBv6g4vyCVBhNaAQ/5vV7gogPckuYEFhbovHUWlR9MzAroZF1uzOuAt
rt+LXsrb9A510h6yIPLFdPaIGOyeHgc33pAFVCLk4cIdmPEcv7QK8hEt5nSH+7q2
AR14hLDmd2Lg6E6E7tN4GtMn9tiVgIUCSZCGG/SQJ3DCz1ANuaGSe/oOaGoD2e5h
l0H+zXQ587IpSO9Zf+Lj/rThQ6/vArOVIBgvjbEe3LWmjhcPdi9o2Nc25OtbgNAz
ZNOGVQo17Djl4LtBg5oGY2exn2s33ckv5Ur+bnDBs0wiunhClyiQqBZW2FsawBGZ
oTg6lNA21Mn/+dU29yj8X2YamcsUSNLOWgqgwotY2fDb4Fq4eJBkpuBifNN29DCI
oSBcqaCOFSvkYPHNonL0qgw1TaKoZrLeRmgH+//DtsSU9WD/P3Sgtt2KnQCTwz88
nin64puZnhl2Ya+p+HARfj/MM3fMYIfOQH1sA1hO0sz0j87IOKWz2JB9WCAYwQ4k
nSlDyPqUcN7gemy8PPIJeYy7rQ8ZL9fgJ2XCU8jbp+TSUh7aCfbq+2FvKREIf5ok
O+0cm1ozMtV9PcJb34M3tu5pRmotUpnj4FsruUHQZIOhrSJEUG/JcnncdDVsRjnS
oT5tGSEOi7640b56jZkHJhf/ITxry9SunfrYfeWES7daZCYs78Bc56CyFzI2TdUD
kdwpoT5CipC2J45C264B1QSMHiPbg5B9DukEw3FB6QBri6G4SZrHGgk1W5Mu+1cx
P3IAgGM0NfOnejDtxKbZ34z+qPTyt/pqvG7qAceg6oct3PyFp+oLF3KY1Bq4jsJe
kMAoo83evzjNsNhBASNujQLZdZmS1af4F+XSDFY5876CNE+FKVUE+wUhWpRU45wG
KzOhY5UH/n9RQmKeCIQ4H4K1E6gzV0CNAxBHKJzBdpsO6tDu3yWrjPrbJTAePVuT
3nNkPIEYEeTNRvsPOAdG77eRh4uZ1unt0z3F0bHkM1BO514abuWx83OSOspj7Du8
bzW0Ca1G9Tg3plRMFIDEXTBYTSKDRXkF8nhcNbrX8jMhQS0MdDHaYxiVUNZXP0Dx
Syd8LgU6bGJOmZYUP/9bayvbyKkzql918JdoHZeI9DQePf099FnFmFSrju2Jddp8
hHGs/bK4F2dfyCizvaql3lbHJJYax0ljPM2qqQVBfVkGBIXEpIRytfLtStqeP5AD
tuxlSySuiVoJaPmPMi+qoKptmF+UOmZ//G1j+KEr4jY1f9GE7b541wkWPUUlJmPH
rAkhIf7AsdfQvQSuLGTolPN/pKhgf4JZ8Sif42qMcNSC6yA4dFPxVQ3sGfrRdoQG
C6yReP9CBAOt7uHnIo9q7VV0xbNXnWlbg+De6vX2j7UsSHE/dQ6GZTPmvbTUBZ78
tJqs+dWXrlM+W4mtNv7Q4CBfklkzEYDjTJt3Fkg3Lu1aB93LSHHOozpoObWhe1J+
kvPx7M0BXI7nGkScZVRFyR+7GYI7DbDdARbxKw1zVTDfntQ6nUH79YiHU8zfM1Q3
LQcREG3/78GY7017WnAbIlptveQhzRJhJvqyxzih0K+oaNbCBvKQeI1Y6+H7QeeY
7s3ZhHc78qgvjCOPKVqWeSJvJBX8YgyvVJJ7CMssWdybS/3E6Fc2Id8Rm1CMXbXL
Uqu2AtkB3Mcsge+ZPZBeuFA/tNoGu5/6Irp55R1zK26PvLXTy1BGDK7S/V2GOMsf
vNJzXN2EsT2AOqsM5BE/Q7lNoWfdvC9Q98Xkxcd7eE/sS8elCoaI9knBkrYwtdWE
NvBQ7wg4jIj1jjFa+cZQfNxdo8kDFQVISGibcqBcQuLdCtQ1l9qmrk15Mzj48o6T
gBD6qYibpvX1Ou0PlPE77FQId6g5b+1zya/aZ/8BzW9Z3cunxFHzqvbhmf3VjRE4
mCLxw5TjvbTyf8RC3siccf3a4pWZUi057iqw9rejozkl7o/oC6xgzKLVD6SoW2jz
wvZSXDxHEr2nwTT17x/75poRcKb3oqCaPEW2zneSBErepCsm/t+s7Kf65u69NlKW
HoU/Vrahr7AUsVeDslMsTrD2yNuAjKOZ71yxKTM9hqmJSeObYFMaEvonLMCrHr5n
Vuwn5uSi5ZhAXzSzCceY3gJ3kZeIWGOHy6LGPGqk1JeIH6ehxwfb467iKgqoWGKE
TWlZ7oy45EA6QlDrv7sbfwROHqbz/+fKa7aIF1HRfeS3z/oDQ2KYEjVu4DCYI9aA
RIz/fAZOfg/HiPi/T3FPO7Bs6Tub7ciZ1MWa6N9PCY2iUAyf+C/T75UAqRx9ZYgH
x9zQfqcRth8FAWcdTTtRu0C3l8XdkUQWTuyqcVVGtG48r69tAJVkaKr/7biV3/tw
0veUsBtwtcUM1V+0AEcCNqobXUWnwhgZV87HZ6v9IYakBdL8RrAOaQo41EgBu6gF
aX+RzTrx/q/cXT3GjcOO+Tghpcl6OK6yhB7A3ODSIq1hfo4E6RBoB36sIIDA+0Ei
/9Nj7DCXLM2Ld7v+7xhx8Rz3KZ8V+/aZ66JqYHeMlq9+HUgQC22Dpfk76k/XuEOc
7myhrv0SF6/xKJVO6yyinYKjnWCwuTzmd+tAKD2W3GZ0C8FCktuv/6XsyWD1Morf
DmUwRgjSOmNsUyJmHr/asJy/MlBiVaxEwApN0PrT6nc/ICXxmXD4d2z4nqg7mvN7
IENgP/4LqbMBUgUt3V+lRavjkhNbOuP/LRQaYL/QbUSkP8pHhekCmC/h5wwTvAZq
IanB67U0l0Bv50KgnCF/bF6O4Mloz2AHJCRshLMB+Ilj/MRbIoQYswa6sNf90gGb
fVED7nb5fkvn/de6LgCNCsVGCJhiuyiHDNwS3C1VXbNiPIg0e/I3nR5Z0NogxWLq
4dPxGEdLgFukVCE7+JOHK3XEr6zaxRtZUrhBJLGvfrwA8mMav/9PYjJGCQCbtT8C
ExXqv/CSv/rdRtSjl6jM6M35ynqM6DYSdVcOibRjtY5pEnpjP3pZFKQrweFQCUfw
9AJCctd+SVL1SeZlz6RhX0h9wyZiZXiEcQ4nlwFgDkLlhzJm8XfFBHfeeA69ndZv
VVCViUAEf7kgnGWOeueTMQvnLPBugJpuBefvPOYYRmORp1fjmSYiLVckOxFoV0PZ
qwVnb+idiOjv6GmNm/reRI422kuKZxUVP7nnGqEw7nv6Hk7tBiVMCfUEDZzb+Zxx
DNC+ai0wZpjcBM/xSTLrQx7k8bEMH+t8qZ23cIzk5kB4WTWqFn+0F4Q7v+nMY+DS
IR1oJce6Bw+pMN/Yxjzwqm+0gMdYTlDZy3cD1eBaNgpmQAcWZ7/JGqPWbKocspvV
Pzap1nAnDrqfntp9eCJz9wm4ph/NBHc9hJS6ZI3LmB37gwW8mwt1BM23NtJwtvq5
8jNW6x60l7NrhLgbHmBN27/Y6jTPN1g+sn6MikL7+0P7iNpYB+PP8Kefgh8p/wya
acGTmzelXcRgR5Kpuz+FzylR4pPflID3p3vLjg4P7buoDOrKFBPC3/OvflqqIx4l
p8Mcw6MnaY2GmT/HO3FunBwGQ0VjiCtV+n/k6ajG5A+zoYxc96tdlxUMOy0ZtI8E
RTqb1pmc0Fcw99dZ/AGQTBVJCzUduzbZ1D9xykttlVSyhbEdMvPwffBB55DpBaq3
Q7bM1zeodDdumxEhOnog62c8xK5qsuRVpiHcQWsK5e4dBYo9paVpqjjYrayjTwG+
rH6DdI+lviUqbSqBEKsX6xLuI6sHt6bJHyJ1XbJon83lhjO7ICxDLJBJu6kZsKqG
OukZd5575M18Yc6wOhJTy0qCHwAp25Sw9BBmoczTPOeTQRkV8LunIEoZqDL9QWoX
s1n8n81neGB8Yo+KNdFmGIfpgiYhSiB6XhWSgQsZ6TP/ITECahh/apBRyjyQEaGi
vhd/VCJeqyTbCqnKX6wk9/r1eHp6fRI8DCtuGx+9LPr/+hbtHIDqYirojaRdlHOg
7oL9rl/6UIimAIRclagO/yak2qPKTTX7ZZS2G88kgBvCBS/xiEANFcFOMt1Qqiy9
lWFiay9DrWYIL3jkQHLsKHe0M6bq+Q/j13c6+EeVATPj2Qn1diogXeklXLqwbH1W
nLFPI5zV30b1J1UFqUvKCcnMrLWhdznEQasBekQ70HXoFEoNiX11U4SAZw4+aL+3
P7qBo8n59XNI+H9J3kZfT5BnFyEUjWMWFi+A3kxTxaSWA9DfpgVfr14yTOZ7nBEC
ecqlpgVMiiwJzgWaIqLfcoI0u51wDXkR/elFl55G0NCxki+0ZZCC5ZNr3Cr5MoUe
JFAhTzFRXfuRhE8nxwEmfv14v8RvopglTpQSix6qwKzqWHxV2RFMGnnlln3lMxIj
M4iYmlAWIsTJxJRh074OYH/OiopyCIILDbkbaQLOwpPiGh3f3o1GRaOgyiCi7lSy
8YutPREYJ1jJJcWhM4v0orMoU4dGcO5gziiWiK14qk4WhJnHM1wTsb3BNmooqmfy
NoxHHRIC6UwmYjTMCO3PGsicfz0BneHa+i7PhiWNIBhjJTx6SNgDIYN+ytjhyrwb
k9x3itHZ2ylAQc7/34ZmK+KkrDEa4LZ5Mir96QbU/rpwYlU2ya9/vIP9S1j1otMZ
l1g4i0fpe9kO2dQqV3IZWTRz6CJhCmlziBiGMMxz6mMOfArthzeXfprZJFe7kbpT
pxXEajt05WD0VYWzCoVEmj/bgS+tz2x8Sim+a0Bhe5XzJiU7NbHNPuDrQpNYkShR
BZupolfx40KoZGv68N9trlxwkte3RMBWdIarg+gHsa71lcOBm+ZLSvgzV9DISr/y
rgo24Pp+ewEGv09mrr3GLen+I/x2FrtHF8cdjH55xHj6T930bBaE/ujZTWqD/CDy
BQNFHwa6CJZB5d2IxhRsYumsRkyrrnPZBlVSoXC278Hr+arE9CvBZsaWpjoJ83jJ
J1m7SwHyUgAfHuKdFkJS01ufUMAzNko6cV/98NgMoSCUr6h6gpuFM3JrLxmGoWpM
vA1z7KwkiOE7pKAMeK9RWAK5vLOIlfwY9P/ucVZXJumAyypeaYhF7nwZTYFXT8rS
S324hHkGGZY2SE/Z/fd7c3Oo3olBKtGGus+I3nZdLRZh1OlNRXEM8cktWvrM3FkY
cHkgmPwJtzMuCxI3GcpGP9Whou9CJuaH1zAooUb+lL3qOeLVDpF2hly0gvzQ6Jwe
JiBuBaeYHPyPjsVPT/99RRUweuWT0NikeIbSrLyV1+Qs/PZ5QzaTN/1r2mqMJn+H
uKEw/OhZah6UdQGUyqQGeuWBqaSKAnZKWq1Kl9jJVdfE8qXizWdnubJmVn/5UTBQ
fpS2DxBW3BHfeXHfrUvtF52yS5XCMopcW9wSuOTWUttQM9TfaMwrBQo+/uJVdsJA
9JkVPu3rRgYpgwRt4qqOP4LxdAFiynTqNEPNf3jiM0EiMwo79/nGaC0PWOA0uBg5
+Dkt8/9rvYx3EbrFSb2BWYlv0caJqbfjkcOu1HD0CbK7RsAgJpX4bfdwE/aw3/uP
uGaZ8gHvmkWNovhANHDxPOUA/cJwBLlCtEVEaFjA6slC5NdKqsTSMZm7zUpuINAG
wgT7gYe6BxpjPgpWjQBVQ28WrIVRQxUMJy7DPR7gvIwS62S5kxYgZni0mTneGipu
Uewey2+lcvWZ1v9a/xYMuLK7JAcV5TiSsVgG7qZhXwVHT7YdxYQtmzLclSgzYdn0
LiqkAFrnYwUsblltzg7eHJVwEOhDzDWlWxBJlGdtengAqO8UXTQzzzlB8/I0iemP
7B6YgcfgQzFe+nEtpjA5js6Pnnzfw5HEAS3uTi5eQRXCi86MnqaFotiSpKuynRpJ
7+8GfVD9qKT+xE3HNZvjHk2lWZaA2171aeR9a2vE/Odhib1lh/a1/DP3tFahROlf
ZWePTxy22RD8pd1DwJNh6qUs8fh96lsi7A3AHFa0GP/DrhrPXiwiVa8pDpmvEb4r
jJV0ClKr3CqRhV4ue1ZjZlF1MRU+UpHMkOmZ+95F7wjRuHY/LctrsSnAGyVN4Xks
by8/54taHFdyGbkeXdkYfPHG0d1I6Cd8DjYhEuoB3qpdp8peVBzX1glNwmvLoNgW
h+nAH31HyRj85kw7Erw5WDa40wMx/AcOPgR54xfeHOLE9ailqvMWw/F3s0cE8Hlp
qpdtMCR62mLA8Hu+AGi3eHrThrYlM7gR6IXrd/yxLTA11hvQFt0gN7MV9CWHT9oA
EQLqVq3aCFlvr3FsWsqTATgD3EpZTpGQXdw47MIoE3at3ipgJkuNUk6egeU5K6t/
WuElKir0ARpJUBmapNxWChEpfKkl+/uuhPyIipanhXiApqaH8eeHY5Pd2tpq/6x0
b1mfL3JPSf2hcbD1uys1Xub1GXA1iZPPou9KZEN84IuUY2VQHjwsqjsWmeK6vMjd
Wv1un/QXmpJTpfDuSRyX6aQgz1VZjeled8KQIwIqMf6siXt6cMPrDxfqJQRmsAdo
y8f3ToDjn6tA1iPJO8N7TWtQXRtd+lnw0MVJO6Sw3+ALpS2SFlC9vnjXsAVorszr
eTDkPyMnUcQqP2FArKzTm65t/Y8uZcyMgUZD5ywcnjn3xY1LdLAriXEe4ylECRUu
pzf6rUs6ZgOa61K8hmU/T85xax0EMCk4VNifuzUGgxVQPiWcnDmH+N3Tc+SWs8vO
2SmcriqN/ME0NF43IDbxrFsauiUIZEw2dTq1pvKQLxdoD3dtIpGkOONfIe73Kx0g
o+V0++yTZTj7BwwqDKUuKzo4fZUU9SIZJGLzE8rq2SpdU1pCy7ktmJQP6qIA+fho
JF2eeL4CL8mij/AHT4VMM4wwNZn8y9g9yYlSzwdWkHHoSwEAEilenM0AkzM1BF6j
xHm2N5XRYbEGNBPcDjizEaE8lxYSJmcAVqJxGD9CiNDLbMuNmuI26hRCpVaH589B
4PmNV+QNSyR3y8nc1Ybbvq35zLk54ed4J3D6kbtlA/cIoUsDazV1tScW2QzKOht6
rkheptskCd7845hXWoVjQuPI3XjtLijEbb7UrPOuhQ0x/83STE7+LLKm4NJKqESF
nxY2P/WvVgqFiMJ3dq/x5yxaurAT7mckgq2bu2mI8QklGqG0ysc4mg9bEJyIuycU
U6l5fQcmppvuPC1j0oh08iBfqv18zgvz0pr/QW88Q401p1VqZYJrypHeXjqLE3hM
D6p2RQftzhTj2ShcHylKOeks0UuKskBj1LErrdwSggBaW+oSUdWdKdCRpIlJ6fEM
Uwf752Q7ZTZXaZxXwpjruLlQ8FISJnr+vRv82XM9AQuLtuN9HwY3U12RERZ+4vOf
pQPfBR827+2zFbRCOu/fJnlyldzUQ45MvSKnGwNy09LcI0UtCpYcTN3n5ehH3mrl
3M8hdWCTcdvbe8z92T+jitJMqvUUZ5lWL+oLJ8cmtLBFCW2WfFpfNvk76mT3NRyo
MsVVG3XxM3jXupb4A5zfXxVcOiahqNH6Qi4H6ehT/aubWCallNcWARVdBvWYa2Z4
j1aIhXM4Jd5LU13yp4aDOD8yZG8ROmHDNVeBef3Ks64o342r9hZ1MtBJQJ3sZDP+
iV9bSXYkVLxLqtkW5Abv1/oqfcN3nl8UDGmrRrF90g4p2b2mqS7jQ0TOXzCL7u5m
KSubw2g0DMeSGI+8yYy0MZmlb/4gCQNOA0l+ICkCmvEHcuLWfj8jA86W8dbHuS7R
PZKsnGN6vEFbLDOSdlCH036VRJgZnTh7cbQQ7TccdrnIwdTrnuPbojbI86juDNty
sWnWi+ZBpytf0pE/p3G2yzmIALAi891GvCjCIHendfgdW02SCWa0ZvB1SLO9eS8H
OdfM7Eybd2liMS5xOcHHSIH2WDUQhtvx6PlymYRx85CvLJUvOcEjEqwZuxlriezk
qd2VA9PGB4wM2JKOUMAtpNrRQj9e9OiAsvvqwELVzZ8GqpLI1UHC5NtBcHRx0HcR
47Wrm4kuNEEG7Hv3RqTfJfi2BSb39YtMwYV4SrHLnZ5divzHEbvulEjFHvGB3J44
8m7Z8J9qVBZ87aLO3BA6mv7jaz+Nf009ljNbg4lZ1/SPwNViGPKvRH3QP/wiUkjn
bYPP3VlJWXPvt1RtAf4lY732cW9aYRK7LbBD1dlq9ywFmr8A6Cn/3TWVGhj2JdL+
kQK+8LZZuOv0Vjy5R80AoYtqHF+KKcIqGBl+pMUXo8ViJKjy7SxYUv3dsZ7LPmGR
YVDYumT2If4phS3Vwbe1OPf+wEbUOOoItBZh49aWhj89X4EV3DxcmPSoFihqW2zI
2jKTxsoxYeoZhdlrJsnTW/zAIr4W8MVWdQ7WzPPGXOtsqMwBE4o8isOZy9v99YPe
9bFbuw71F/4UP72U6Q7CBikMYE5nFKU6n+wQHwhhUj++FM26yiUT1ki2hmwGZ7tD
MqY9edzjsqM+mEkf5WnzHaau86YWbTHgnqFT/rVlqL8ESqo1aNsWpNlk/lqP9g8e
RFgEx/00KtqQtlejQHhq+wx5dgz8xABN5PfPBY+0Vn0DIW1IhA+kk62bE9KbFP7w
miNvFNJ1G3AQ56WTB8tKMOYxDexOWlCi3p5PtYUDVG3Idwzw2/3m02T+n6ul14tt
3Q+SLytuNpJAt/v3io9RttEfez2OzM1t2uImVOEsLB3/Tjxksd8nXt6SSeUD3JRw
5eFM2nmcQi65bZ1XJtS2hlyjJ06pzdAA0mH7Jb/G6inS8KHVXcPQu0sULG/6yo9o
/F7yx/CMCFHWcoyvbVlpRJJ9JwC6m1MeriYTSOS9xWZFeEp1aDdMb1lkfsqELqtH
P6AoRrFPALVsci5LbGRAZV7RL+10agdMmMKXqJc8Yk2uVHo+uNkBCCBrnHYQ4BuZ
6L+xYAscx5bZAbxthY6m1ocGtIhK0te15e/n7tVHSbCWzayeFrUv7h7Cb2Vh1sp4
E/c/ov9n4HS8x4uc8MZLVX13ViOCfbbLJZcxk0HZPpMXwM44YRPS5ZYX+AHBmGOn
pZ8dcEFtHnG0TilvxzuBC+NkIutBlvS7NpwMIZ94aQGTpnjPyq4PmqO9ti+XSWQ8
jE5cagDhAvOfu6bL+efrtBptiVyZ6NHdhUJe2E20eStFWwweV0Zun5vXH0GQsDm3
P1o8deyW9I+y2fQcg7o7xGamCaurCZc/w9ZEIlFdTYwPL2kzSYITOnPr8b3lJ5F6
mfkPVQnP2X5/7qZsn0s7dnj4+lFC2pWcg+QZ65MavhfS14SaQHRpDLfXe2jbjY2d
19p3VQKi1bOqY1WgbuHbxXvc79p3iGu+mcVZWa4/cu0FhmqoVt+4YldCT9GW/iuZ
+I5ZwcbqTwzIfYYlRo5sNjllqBhUcupTxctTTy3fIC/Tt2+LVIF0XTuvYFk41gCD
l+cJkZQSzIWij1Uo7Gi1R1T7YnDXqN7Y/i0Pa7oIn4g8MdQwfN8OQ+NQDpSjA06Y
MAi5QhiEZAVqkuJhPeYM7SxO1GD0FpkHRIcDeKV8ilr3tEKi5brkFl9cVm4AGdz8
bcv55kucxyDWQCQik5iaUALGlQ4yIdq4CfTd7pBieI+iCai3IswYgUHTR5E7xi3/
GOzGDyuRbxtRmHq2ayM0wAJPUqN0pXMHMRzcIR1v8JH+z7Pp4pXrOz76B56yIsSv
IyCE7mSm7O8xjZoMOj9D6VHCrxhpFUdCtj3fmFFbvA2XoO6CNjSpd4w2CR19fZJm
nQ7Wm78fZlPlxmQ1V8rEw6Sm5DXc/zDPUv731+j5IVmZluRDouesgVTrLWjlEd0I
MYZPE/aI6o3hxFLCnHy52LefpVRAxu6E8/29SXKWUrZCZsFh1MWnDztA4Uy+5TKP
xB1Zk+waUsdh8PofIkVGRA==
`pragma protect end_protected
