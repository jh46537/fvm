��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�{���dʂ�V(��p���ha'�ټ�y���'��ZB��r�O��O:T�B�j����w���ګ�c��	���7�l���A{0�ǉ��삇��$�N�n_�D8ҹ�	`n�;�U �.��"���7��#۱�&��s�I�+s�\�dvN�uh��I�[�*E:]E��M��� i�Z�H[z�'�ۤ*�#�Լ1��IO\�؉�_�f�M�n���rw;��"V8�;�Bl+"ޮ��-�}��78�ءz#�Wz?o�k�>�  ��:�����%.�).=��'�ښ�^�;f&�������?�C9�3qB�k���3IIu�z<���{�[P�2`����X�[�AK�Z���K�pl �㳵Bz��9�R��b��(L�jw8C� �F���7龀���]�����P�Z�o���V5�h=��,`6�6��/�]3r�0R~���{�uߖ>2��@�_ʮ�ou�IV 9&�_zj���Ɍ��}�ևMfEH%Z���D�UZ܀@i��PmȳĪ�t�����M��8)��c�"j!�%���E�r[�����&�AB�I������G�_�2�J�g�$���i�y��A㡰#��]�囬�XC�]���m��H��,x&f��7��/�L����w� y0tf�rϵ�
Z�7�(��πބ2Z�f��k7K�m��wR�J�b_uQ���3�l��`Ͼ��o�c�xҮ�V�<ǰ�8_�8���7�
��r��!̣�X�Y��X��M�3*Pם��{1�3I�s�J���Wi���<Ϳ��w��� �f��HےZ�+射�I���<*F��)z��(nu�����@�I�e��)��� W��s�X���_�ݤ4�����W��p�G��n�ㄣT�L�ݯŃ
�����h{��s@h��4�xm�-�3{��U��TLB��쨯���4 0��úޟq���3w�2��&���-{�)�=`jf�����cTG]��=2b��c�����-#t�g��j�S����
�3þo�,T�{x��>p�'��^*�}R�_������3����������ZN�G>.�_�伥�|�����p��p�L�ɨ}ͭ����B���H�S�	����KQ˗�Ϩ�DY��]���u]:�*a_O�6�0���-{ȳ���V��S�q}W�[�R`�R�r���K�Si֌Ӭ�{����2)�)��?H�)!5)�[�|����A8k��r�iԈu������MHk4�2�JH�a�-]6�*,�
�`�8A������>f�?��Bp��7s���p4��K��%* ���F��K�	���b`���IC�|��^Z�Q�[(4�����8�ٞ{wl�w��Y��m����Yc�^�^�@c�D��ޭe�>�z�+Է&�%c��t�
��iC�M�/Pۄ��Ȫ�81R�&��V�l!�jGquhO�ވ���m��j�-�(����Ί�Q�"��&?u�G�i�u���f��C޲nK�M�&��>
�P6Ba��{Ɗl#.J
i���V�{�I�u��f�;�����p�B㶲6e�_�:I垝���C�5��M�D�ɚV�%]r�O�Ī����d���c'�ː�ᭅ��N���xSR)i�ƪ��tr!�Y�.��X��h4��Ѫٕx:��~\���F�MF��aB٢n<1VBS��EU6L��D���EϜ��g���4,�)�\!$��Ƌ�M��
�Ö�N1;�]�A=ԺOG�^�,�16�IO-L'�m��F)��������B�S)p���������q5�Q��4�I�$�&�&h�Mj���AZ�T��Д���ͯ��������޾3�@]�I"HfF�l��ǟ*�;{=�2������z�{{(��4�G�^fx�li6�꘹���S[��p�4a}Y���#�TԀ�`m��Ceyt�~v�U��Aƭ���]�u�-�d��Qɽ�_�y�O�e�m�P�(]�
�zp_�Yެv�r\�J2�]���������b ���򷷓t?���
p���T4$jp�����1��#�-P�̶?���4�'��L#�:}�o���^ҞCk�gS�0l�`yj�l�׶y$fnU���ZAN��h|LPf`�͘��.����8J��^U���t���}Ƶ�aٷA��J�[�
��{��߶�7�m~�C$�c)��﵏����J�6�3�7��_��Y�az ú�!%29{PL/^=c�֕�p�0��5!/ޯ���ݡ�����Pw~M]�Ћ��|����q�˵��e&46 nK0vD��EV^����^�c�IW�Q�3Ʉ��nN@%Jqcc��7�~rLZ�=W��gJl����W��O��R�W\�j���U_�O�]	�l�<�m��e|�r'��v5��i-�Ӵ�2�`�G&~�7��q˔�݊�Ќ����㤕g�l�ܥ��4�W~s�/VCM��r1\5{IQq̮,ݭ�h���T4ԙE"r�3�!0�_������w�a�x|t-�|�"����Q3���|��H�!;��Þغ�3�
�'��}C]>�JH� �@���Fl���C�`�Ŧ��
0����lߍ��^�+~ ]KX��r}�1K=��2hk�#��D-n�'� ȋ�����[Ş,e���U�[aOߌ�o�<�G���c���4�ѹd>M�>�����{�pۼ�;'���������H}M�0CN��Q�.#N�=��9ӻ9X̟`��a�#čx+'�-��1��̬#�	b#�kǠt�q_����иƣ9�)�r 2:4�]�ɨ����~Sv�C�U4��I
�pfw��V� ���(6�8�JY0rr��	1fC�u�����45�0 I,�
��!�c߉����98�R2��䮊�@�hG���0�x�"ۅ��[��aB���L�hkpmgq�B��{�Y�Zz?�Һ�t�%�U|g�+)�L�A$u�5=y�����.�$�/q���Y�$���#���.��w_/��[y~�$F��i�6������bd����.�gS��ʖfz��-֪g��
C�ATPp �M �<ܕ����c����^o���e=�=R�)Ξh����j�[}�\�+g�b�[E��X[���W�������;�{Q�_�2����R�z�ę���@b����K�:���	���ޓ�N�=0w1�=Y�&v{�⧶�Dv~u��̉.�v$��Nh�G!1��٩��1��j?ޕ�W�M̠��%b(�r��K�sPDKih��j<��2��q�7�~x_	�|ͧsƶ�b���6��J�πP�Ʉ{1�9�q�n�h3U+Zܹ��!W���KA`����n�u��K'��r��p�Z�;��{G�����n]�:h/��,��]����g���Q	��ڕ��	]vC'SӻO�M��R$ة����!޳�K��֜�֊^"5��̬9��<��W�)gE�Sf�&
�3ܼ��)�!�P����= !@�=��>�=����a�k�t�K��X�U�W����*�R�$B͋ 'КF�J
h��-�#�M��mg�-~��G����PΎb�D�V�����w��U'��F�k�?��!~?W9�*�{�Y3a]�a50��(;诖���7�vŉItz{p�V��M���u��?�Õ��=$�y7�-Bҫ��u�L�Nu6�-�c~�} i'4�Yh��vC��~-�Qg]@��q��/�SBN�Vg�~e3��<w����]V���[~������+Gʷ'J?�&S��!��`T/�W���������"����m^"m����L�X����E���6`�t�bj�m{�k�D�4�� w0���l���D��Nt�:P� ����G���6JW�o˥	k��M�r�>txP�W�\�n`I=�Pȕl�����.�X�,��B(r��q�*�L*�{�Y��D.�)���4��g�2�Μ}��5�%{���Ր��@�o"G��U"��"�0_-0�\U3�Ҝt�$Ig{0q��dYց�dT�Jfq0!���5&�����d�a�����GÄ�M{S,���MYt�4�t^���  ��L(r6����ď���22T���h;Kf��RՋ�b�˻������3<W��iA[9��~�*b�P,(��Wƶ���[nOCk/3�A�,9���U��xF@��z��ݾ�yR�BgY�|L�^+u��bRn%Ҵ�7�I��9��:���Ō��|UÜ�$�W��:�y"�����/�e�i�b�z:x"���3����>	A��-�R"ie����s4씦h�����X����=Q��g� ��1��}Y&iD���z�!�ɪ��s��9l�qݥi�j)m��rS�e�����CJ���tz�c�)K4-��� �*5�:<�ڃ#n���j�*��7`�܉݇�E�_۳C��9�%��VhW����9ElX��WI}.�Qx�q�w����j��
u���� !���AK�$	��<P�Y(�[��ЂP��e�m��b$6���J�ҷG��bE��8��n�v�mV��`���PjS>9\�����[Rk���+L�ya������yF����(��@a6�T��;���������]P������<�o�� rj{������j�Oae�P�� ��6$Ӛ������^S/
RA��	:��d���Ť�҆zID����;�ҫF�9�Z�c��z���-��Vҫ��:���7�o��6��~V!�'���$I[(V+A\�"$ː�vE4�o�<�$eY��YP�e'����ӊ~V������J+m"D�;|4sC���G(�����@-��M�I"�%��Ow�n�����U���G�+?Uׂh4�vhТ��Ĝ��p�A�В~�R>)i���/a�Q�2=%�2�Kh2���� ���8Y+�lU�Iz�_n)�"d��y���-U'A$4{�c�b�X�uC�pƪL���DC�7�������9k��_��x�[�5��������봻w� �ݍ�&�^&�o$�fw��s�M��/E��cg]�v8cR)*FU��������[��>�u�pQ��#����?ܴ��ð�?�J?�Av�e����T!�;�a�7�J�P��5�1��nϮ!��O9�v:�q߆I����������V2�ɒ&�SprO���г9�w0 ��