��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�p3t`�Q�|.@��Y�������i��<b$�����)m��x�2�2g�<���w��c�`rlW�X��p�tG�iY�#�7�@Sϯ�A��Q���AU�9���:2�@�_Y��Z�6h��W�*�D�Y�P�����i����"��Pi��l�2� ﺮ��e�B��f,��+H��$A����I���ӂ�c�jG,��X�jҏ+�t7UC�p��D�KOfź3D���Ei9��A��>>�TE�~�W�����w%U�(�*���mm:����Q�g�o�_.�bR[�������`�+� ���O���\8mR��ZL�� �AL������>�؁'	�h�A��yU=�C��?t���ڮ����1F�{���b�RX�p��'�V�>���ky� \��؋n����իJ�I�I��u�v�+�{Z#x
7RTK
-�6���ι��:�W���9i_wd���e#��g�W�K!r����	������7��=����IZ��zH!#��`Z��T�^�������nh]�,P�s�!%�G�ݓW>HNT�5E����-F{���@�-�yxYOe�ȵ�}8�+���ƶ�B�(���d#~�����3d0ם�̎������#j�$W��ҙ,�(u�R^OU�F��HƄ}\�)�PV�8����vy�<%j3}h��?�.I	�$=(EL�����o�n,8�����y3��ZQ�� ������;_/'<�RI�A�`_��~WEF��hX\�̕�ip��W�6+�����D}��2�/�@�A�L�2e]��V��F��S��jo/3��$��	LzަùL:'���	MÞn^��Q�&�im�L(0�wM^���Lp:`� �I	8Rxmc�>�5]l�7~�F7�� +���c�R��+3������y���N�Q���yB��$T�
�}\�2O��l��w�|���OL������z>.\�Xx_@�Y�<F����6b$�F�mK�M��30!���c��.��x�]�� ��1��VQ��׌��1[̆{�O���+�M9]OO�t?�u�^qB�("`cI��ԲB�r��;<?[+���3Ep�2����/��� �,ͦZ���_�O#��QSk�\�T���^H��f��[:�q�`Fd��m�1^�Q,q�۟I�X{�3e�m��.��Pj��v�48t}��i��ʷ�T��>�E椧��:yw����<$�;1�3�A(�G�񉢤R�[���J�! ��(�H!��� ���
��0�[��\J�$ܯ${�oL ��䕸7�#�"J�T���JW�<H`TԳ���h�����r�j�e�H��Ѝ�s^��x�o��+����I��f��#V��)�5��Q��INT��2A����.�U�� �`R��*|+�*`�M$`�H�=;���f��a��\s���"�1d�}��f����K}7���u �� pp.��:���JͺN��t{oa{h$�OC���U�Ϫ<��bh��Nw>R���Q���\���T������0�gX�hs�U�X����x��U�V���_����Oi�7��}�1��rp�%!�*�@�x�Rj��}�&�f-��ʙ�����.*B�ã��$QH�A��M��� $?�R�h�sDJķ�1�f0~�/�ad9��V���O0:f8����?9	\YB��Z�O�s"O��O�N�gS����\�YSw�#|��;E'� �=�U� ��qq���籬qCM���tsH���tx�[#>l�#�"�=�p��)�+ W�������G8ua�*9 {�Y�0f�L�m���1�^�:��_��~]�B^� ݗ</I���@3����Q��:,��T9$���e�4�zREa�>�Q����S��2�����(�
���D~="	��u�K��݇�D�N_(f���^�8���$�DB����3Jقpl�ϐ�[��ZliS
̧,�G��D���薕%��	�x���F���nװm�I�&�!x�J����)iA��Zn�l�-�)W���S��ϐP�]�1�E鮁�i�B��������Nٗ�G"�Rt��۔QM�ШQN��:�����{$�ʗrȆ� L�[Ǖ"LW�g��׍�oT���c�Zuz�3+_u����d��$2b��NA-��K��6�{��̄��OG�*ȃc�=Ŭq��nd�{���.5!Y��:����I	/4�O>��:�.<`*6�9QրG+u��?�#��>'(U��
��x<��o(�x̸��xVja�-ؤB�7�:�;9`C�ב�~`L��3��eא��]DB	����[�zF�挐�t��}v�.j�=�\]�o9u{w���~{y֢��J���QT��gq  j��O+��x�%��loV}D�O�'c=3�y6��Y�+�ޔy�6��s5t�ZN��o���i^R���Y����q�S�j@�h3��E2=XY��E/��:�|@�!�A2l���Mb�_��0�o��xd�$�
�>W/j0����d4K%#ԡp /���A���L�2���{`���=7:}hjK�Ϣ��m��D�Oԟ#��iH���ZP������m6�Y����6!������9C�豮��.�y�W�_l�A6�.0y��+%Χ��G���,g'V�2/]T������F$n�[鱃z2�v�Z�d�hs�t-��$�6�h�&ሚ>P품�RjP�$���VC�AN�ߘnk�x��8�"RS~<EXx��>�j��v2���(��� �B���sH�ۉ�+�A�6���i#<w�b�y��?|�)�Q�J?'�B�����Gے�deA9;��2���R���*�N#8���%�>��U�eF�~�A�FC:?�s��/w�m�����н�* �/_���w�7��/�o`�����gP
�������6~m�w��YQ=	0�2F��į�g&.c��7�@ݕ��nX^�(��c�;�vg:k�/R�x6��Η��ȕ_;%/$�ĨJ��T��Wr�~]��"���dc���f���\D7�ƣP�a�l�.?�6����qht�M_,�`����	6lc�=G��ԏ�Q�@�I�%��%���UD���}�T���c]�1��Ծ�=2J�֝N��^�f���ww2���l�P�]�����"P�R`��EoBbs��ω�r19�y���X�~1r�i��R�"΋�l_����j�6��CX?Mik�c"Ei���OY4xC�
��Q=f|����L��W�k����q���:��g�)6}P�u����Mzcj^	�+i4z�W�&�"�#�1���甏/�:��,dD8"�xdo��]{H�}3
�h%�!�z��P5/��B��=/�4��	~���A���PɈG��OFµ����~�ڊIBe�a;���Ol�Ë�A����WHu0�&��(3��%Us`0'.��I�~�/�Q���2LU����j���C���� ���.�A��sZ�-������"�jN"�Q�7��$����37����e<�ֲ�v�p��<�4koԙ=ŉ�Zf����!���>J��h�]$���-����{�����L���{�"U}�P��h�K�h��m$
*	(�#H����ҟq��Y�ͺ�����G5x���Ϡ�_P������������+ë�\,��p�`pxd�86�A���^U�*���o�T�&����"ܳ��2��`3#u;H�Z#�Zy�-&~zǿB����>a�q���@?2��;h���j�P�ۗ�c�b5��X4"��	h�'~%̡��]&<��	����s�Q"?��@C�h��j�ݰ�K�`���cR�Q�LK7%@������}���ƕr�n��OQH^7�y�I�8|/�$[ه��j����R��o���T��C�@� ���k�Of�l�;D��NG�R\~r�,{�\�Oc�F4U�ۓ{���N!W�*�����qص��s�����s���V���8Jh�3n��\8�=q��tc�{����B�;-����& 
�����gԷ�5L!�G���dF)Ʃ�l.�_[S�0��V3�P���bLő[��E7Hcc�=�נ�ژ�G1�8�ɴ��\��Y����zY��)	pa5�ΘZ��"K�x���H������N���l��)��Z����T�'��lَѬfa�C2�{�*�]�'�Sr��Mtm"h�**��^F�w��p4�.�^dxa��p)gfy]p��M��T�+�B0�enϟ��|L'0�=x;��I���T��*��?��_[�>�]܇j��"m� �;
������PJ�{Ѩ�]�_r���sm��߷�������J���]�lUh%qp�n��t��W�)C
�D?��
�;���*�L�7��\��
��A��ڪ֒o���z�6h�u�	b�;��	G���aDIe�%;%P����Y�#���=�b�H�4��]���s�u3N-k0���)ss�2Qdu
Q����K�A�|t���?�M���t>�q¤E�x,;j. c����u`\]*�HuˈXu{���h�Q�eW5�@��ъb��g�-1	����)�9^�d�m\Z��Q�V�S A�x�ՒU�c��g�C�(^�`݇Ϡ!��qiy�i�7�їc��d..K�Y:�sΞ7���z��s�+~��~z��3�V�I�2��~�i�K���r�?H����̅4��ٔ�'b�B^��U@aF#9a#�6b�V�Mfh���<�7�8�S�(�{q����ng�w�� \H��dA�sAM�Ry��<ؽr%�)>���� 흝��8=�w��P :��n(_ag����	�2�9#�V�N���s��ڍ�f2O��"ة�3]�zFW�cp^D����N}�_����}Q�[��0�^7mh;}~�3�\�Ő�>��َ������* ��S�/^�y�?��.J:4�/k�U��
�˭� ��h�/�)�P'�d~�K���k�� J�&�c`!�
߯����f5��e�<�`VL��qƂ�Jx��M1B���rRɠ݇o��UC��KXˇ��w׹���	#Y�-�� ��>�����BeNnw17Nξ��9 ��p���ì;�����,���]:��mx�������P��e9~����Ʒ��
[�0��60"4�t�PvU6D#%�,�ѣ��!U=A�,r%��E��ܣWQ��\�ɂMx�Ԣ����H� ��4��Q�-�@Y?4B���n�zǧIa0��E��-��/:���� 
s'a�16"݌y[𛺛~�l����Z�� K��ݞ����A�:�?h�&&�����Õ�/�5�`��Un����u� z���~�cIA�]{
+���8����.ܺ���ʓy���ܧ�$��of�H�z�5��ǔ�G �"���^�f���Z�pޫ�D���J��5ڑ#)UpӦ7��[{��#[��wg0�q��1�5rP���c�8m\�0������!�����(�RF�ml�]��';m2?&��Q��w�ܬ$�X ��l߰A�x����D��;�n޸v0h�I�8U��UV>���ebo�g��!�`:x�l�w21��P"x�ï�>Ⱦ��!��,ս��g�F��;�%Y$��D�9����	;x� �����HOgħ�H��~�q�A)QAl*_��q4�̔f�YX�_�-o���HAB"���W��AX��f\�X���cr������ñ��
���|�䚆���#P���@��d1���"u���"��8��N���Fv�=x�i��Z��u���,AV/�J�����<�Č����s�mO��2���/�#<g������ -�~,�΀
��^��R��n����ɦ�,N��]�2�ኞ�_�ZD�?�:�yl�-4Lj��x Q���ʗ��<`O���nl	��N!z	d@�1�8)��Z���Eq�D�nL�`Cq�VJ04�V�2<�c,��ͅƊe���k�ӑ�_�
�w�������gew��}����5(߷J�@b�5����5����G�����/�B��VK(/{�&����$����b�+M89����=�g߼L��od�����V�-�㫡5�<��n= V����GǸ��M��4%�Sfp�}1S�(�t���H-�R�R�tiPq�r�{���D�bcw�#�/$�D�S+�����E��ܞ�\�������J�O���N1}� ��֌�O4� E�����׿QF�"�>��3Sb�q��S�%���*"Y=0NZ���-8��Wy�Xū�7ڐ�(.�l��T�K=v��n�k�L�L����;S6�@7��&P�Z9&#=��Ih�SGg��y4��3�#	,�e�T�!#1x����e�Y^�)�*�c�4�N#��v���s��<-m�c�L:��йa�ރ�v�޴��֞P(�Oj���:Srے��ş頝R�{Z ��&9�;����L��ꡓx��v��|	�tZ,X϶�8���M����gn���x��+�s�,��^tgwmuY��1��A{� �y��Nxd��FR��`!�Za��V�Ȣ�!�)�����_^��@~/t��,��b����q�ʚ ����):ňD�i'����k����2������[mZ�N.n1<Z`�ѽ'�=54W(�LR%_b6��{z����V�a�!Ɉh?rD���>���[��"���+B��?���3NZ)`dI�@����}�B�n��9V��+$o4_�k����e[Br���K���3�Y�!�oN��.P�@�+�2@,#�#π���jG�w]�d$���B�WZ�0 9�F �&.�=�7�0K2)����J�kC��,7u����l?51��M��Cf�F�@���3c;Z�b���7f"�C����\o���{ǷX��P�&�6���[ͭ&g�%2b��Y(��J�*�a�TQ>��Ώ�F���K�����̪&&��2<��fZrF�)�eS��g�H��\���ǘ<F��g)���Zy��'걬)U��2�ع��Qz{E7��e ��M�+�����Oi�;�Y�o�	�:���E��eLWL������'�_��$J�W��ޢ%��A��<��j��ȩ��]���(^ ��Rƿ�V���5yi'H�&>) +DkR��pT�)�쿞�3�I5�{5���O��\b�@R2]�Tm��*�X�a{y.�#�����q����#e]p7Ζfq��;��F�r�������Vx�k�8�Fm�U~x3�9o����j�ә��h�f�1]�~��tKƻW24��kao�p�B���l�~��&�\d[����OrF��>Z&��h�(y���Pg�0�aK07dLVu��[ʽZ�68��m!��p�L��]���~8��:)��T�sݭ[ڹO��N08^�7��:vN�ӿ�!��QEkK	�j�2[����YԵ��f�^湾�����P�QWe��3Daڿ��@.(U�m��4�M���＊=P���k��[vO\H}�cJ�-ϹB��etJ���5���ܧ��g8X�+�O}t��}�dRlv	�2�}��[�=V
���m	�󝏒__�ཌ>7�����0��bUS�vQH�<L��Uó�,��]��h�e=�<n_�VC��[�[@�2H��	��h���y�Z�Rɥ1���~�Ð�Geլ�/0��^��Z�����.B�r58<�Λ'l�W,�.�j$0К�ę�hw�J��ϴJ��_�ٜ�v
�汵ǆ�y�J�����<��T�=p�2's@ge(Z�:@M����&���s�,�9#D�a
�W�� �����2���荄eWE�h	۷���#z�1g��ya�Є�2#�wݩJ,��?;�R��w�Z�9���.�i��P���+;��e��O ��$�6 ���ӐR丄�����״�R���n��I��uT%t��%$H�����x�[ӃuW>���,_���U�V�T� t](�(w9���@9X�vYxS�n6H11��0�ikr�r�	��<��B{�����'^�p�a�A�B6aT����,�����G3R/}D�K�բf���	~�0��j�-�-M�X���
'n�+�}}|oog"�Z�z:�r����Ұ�9^�X�F�dyλ�[9�����ֳ�vx=R��d/�瑕��](�O�G�>��j ����X����ԭ�}7�ǜ(��ju�廨���ו��Ŏ��H4"rs�u�T��F�]���`��p��q��F[��=��Xu��Q+k����4+ �U	,L����f�w���s�(o��⻪:i���hN���Wl넅������qu�v��Yh w�v6��0��$�,F�C�H�Q���1����l�g�/c*����)G�L*�}��ue�4P�9S�?���'��c�T��[�\�@*�p?˟����l�z�1߇���	:y�z��aX���Pp⺸����M^�߰�I`g�����T.���Q LP�$��qu����">B��14\��DyR��r���Q��qMC��������0�]KO�
P�*��F�(�n��jT�x�*���JuX\�;��u��,cr5���(���{h3��*�a��[�1����[��%!��y�{� ����9�h���<�q����^��X<�V|2u�tA����b��,A{M��1x< M�M�\�����L��oVgo�Q �g�5��îa"ȒD>�� ���G�OW⟍�ҷL�j6W�ӤE�P��N`O��W�E��|��������O�*ޅ��%`�x��'��ϋ���|P9̜��2]�+���~�R)^���A��Y���L#s��E~���]��Z�9*�]>L{nHz�ZS��*�}��Zt��<���NS��%��D�m��`nD9'됙��+u.�����	��~�YB���K�	�4	�F�9*[�N�iQ�kxP|��Uў���F\��
I
��&��7�A���	(�u�l
�M	���b,'�Q8H�r�cHZ���*h'���s�>�s�Mh�ȏ.�	w6qˀe	r���J����m
NӁ�_�4�:Q��� k��6,�NcH^ad�w��x�^Ĉ�!]��=E�t玓D��Ҧd
x�sdN�e/:˫ߔ�+���I2��*����|-}�Zr��v��0ka�nzz�=	9�OQd�����{&����x�LVva�����4s L*��ױv����2�H����U�^�.�,o��.���(�yv�'[��]�frA^�-J�� �̵xA�5[6�����m�ɟ��`M6$Ff�O�d�Y�b�Ѝ��'��Y��
h���=
0aU��jF�x����S�sp�;9�:���üZ1���׵����N���-o��g��A��|g��@���a��fh<+�\���>�f���|���Z�a�f�K�$_D����p{"�-Aab=�gӣ̈���s�����c�p��ٙ�m@��O��&!�o~C�b����^��m�f�H,�������h|n�����*�8`#E��t�QOUC5m^-*v-����=�����]�������4_���M۟5�(fT����w�B'�(�A�#ˁ� �h'������a����6^��Ԝ;�q%�j-g��U�:Bs�(n�[�WF�>4�����}((�	H75�R�X�U`��ዞ|�Z�.B�m�8!���R�d"iI��
C��y�>�%hפ[V���������4;�;]J"�(v���|��[8�"����T�ݯFӫG9ߺ��%*�8Q[=�/u��2����Cͫ�4 �<"�#s ����\l|����s��,��Pǐ�m����^x �j��$ߣ��;�������������0�g��!LW3�L]Ӡ/�|%r�M1�Fb�(%΄��Xs5w��)+/�|�9}�'*�{|���^���ɹ��X�r�ˉZ#s�Y��biD���Yy [_�d^�Xų�V�~�k6��h�����ws�׃]�6�@��5���()��wgf򰧀xN�����v���<��&�}�K}'Ζ�ˠ�o��Atd�R��!�Ǘ�N�5;��{lgX,M������ZR�r��A�1�=���F�\+���V?�4G����K�l_0~�V<��	#K�%���!��\��)L�s��W�#�"k�Ո�u#�ߎZ�\�S��k��˲��K5�=��w��	U}c���k�_���%����2@�SDK�uf׹�3���2}UW(౰/ձ������H�]��e1u}�������JY��|���v/��t����̣˅](�|�W�:MO�g���������í���s�S�4)ԯ�Z�+q'�Cwv����W��ع���e%ɤǓ����3Y�1ն�w����A}���]�1F�2 �h��ܕݤ�߹�x�I��u�"|�+�ʋ;���_�}*1K˵%�q�;��p�{<I��3@-J�:�̏M���''�Z;]��ٕ�'M����T�Ԕ���"0s�<�z�ӡ^~�k4�#�ĕ��.|�b�*�D�������]�d��#�o�3"�J�j���ʵ��?Y7OF~v�|X@����i��ҹào������oH����b�'G���	�e2�В=4 +~�=���q~d�;W�ˌ�q���C2|'l�EW/1}��Vy���e��~yZ�
v���&��O�)��6۽ۊ���X�d|������*����vI1=RX�z�:�
I�?/�4@��շRߌ��+��!���!AWj�t���DNxI�_i�$�����V]��p���+�H7�����D�T]�hsl/I��ـ��F�|`���q��RA/A4V�%)��T��~�d(f>�+�������MZ��+���.����&(�mg�4�B7�tY%}+Vu�[Ϳ��J�v�ݬ��H��[�R��k�ǔ�E�[�PLR��f��mV�<�&Kps_��W#��"���+�n�w�%�p������OL&���v��	����8�T��)���	(O���{����"3���n�:�<��1�?�O�Baߣ���vS�k�o!�1+��m� r,���BEG�s/g���bdb2}|��뼲�>�1����M�X��C�*�⮣#�%�ܸ"��[Q�ĸ�4Dן5�v��2�� �����4����_e�)^�G���
m��6�x ��N
}â�1V�w�n��Տ�A�~U��頻���f����|�y�VR9cηP��DN�*g� 3q�J t�SH�@��=�FB��>��O��0�U�_|]�j�f�D/��t������7ж�
�R�:=��X��G@��^^$� '�;��$�"� �ny�]�e�_@1�������_���K�`7WU���i��*"B�������1p�P��o��`�H����z1P1�\r.�����t����&%N�dY	FKl: r�:����Aq��,.�;B���	���e]b��5�wo>F�Om3���
2)cor�_;p5\��S��0�����]���	����g����7޳��<��Ҡ�����ʠhM|����fjsB8����;2h`�hhşԠbFb�N+�J��(\
��Eִ��i /���Ξ2�՛�<x�D7;A��kw�e
���X\M��y��>f�3(3wDy��O*�F�e�����]a��=�) ii�� @r�N����.<S�ú��?�䟁H-ZL�'��X0��G'	��ʴ��gN��>�9Xx�L��f�"���z������]y@B�?���cBpjR]D} "��V��m��E�?e)��>�tx����뎎��ڝ�����C�@���.���ڝs�<����Zޡs#<��
����;�M�oୗ�c�iq�L�횠���eV�x�Ͱa���C���)�r�����Q��UW�9��T��P7b,����׋3�K�A�-�cYq�ǎ��h�a�i��X /��uc��bEm��P���e�5z�M��ޙ"1��껹Zx-9�4�F���`ä0gp��	zq4���t�Gw��'�B�ۆ1
K�X��Toc�7iY�v�j�+lQ(�˟V��e�I`�R��;�t��q��A)E��T6����f�TP'�+ ���s��w�뉐7�u&����m>Tc���f�C��j.fbb�a���2Y�0c΂�]����ŕ6;~�%�i��^1_q�ѹ�5,��U�M�/��mý��O�(Y���G�������2�H�ܵ���"fq��[P��7� ��`⇙^0f��������`��Z��4=��ꏹ�\9��'Y*s_Oh��K��KwRy����Z���S�&��0�)����cݠ\֟]oL؋�ʢ�XF�`^���3|���4^�=݈�����2`c�$~E��Gd���1�"��eR`��`/��uo�Qx�C ������?1�
��*
��e:8�����6�nS��J���k�0�nv�-�8Eok�%�2/zd��i!ώ'<�DM{���D�d�i����ȸ\�*��B j^w�^��'b�<W��M\���������щ��k8�xu)�K�j�U��}�I	��.6^,���5 ��LeO���k�p��USau�<N�8w�����6�M����"���56Py�"QS�<;:�����L���������I1+剟
Zjx2�-����9�N+��!p{{�w��=}1)�PF,�vn�J�A��t�_zPkQ9��u����;��jl��3��@%�T�������2j"�j�x�lW�1��m����>�MJk�,\H
C��x��Fֱ���G@�����Ƹ���?���yj�Bj��:�⶯J������_x���3��>W"d'�1�~�n�+��8B=#�M��IW�����{4�\yTZͭa �!�|����ί;�-��n{B�y�ys�
�ۆYo	*Yл�1�.��Б�S�3|y�"����P�#FWξ��w���r��ʯDr1 aۑhׁ.�M��|�B���2��9��L��.
��6�2\������7�#��^O��~n��9#���%Eɝ���g�s��K����-�Q�E�?�k��Րػ�?��Tq^�l��h >�5@��<=`dMh����$,��$��%�� 2�.��psD[ŬӪ��2v�R�GG����'5ڛ�U2���p���cW�]u鳝�tZz�`��6�o�Ot����q��bU& �`2�c�����w�y̉���P�V9���@�O����m��&��c�3�-l;5 �!�4�(��k���g:����R�A.*���a��SI�`1=�F
Q��'�kP�mFlR�7����ݚ��|����<;�g��")�,�wWś�c��_�c��7���,:;��b�/���2���0))����#�x���%�h�o�X���4Gr�H��kڏ�5ӂ�'���M�73������9�d
�l�1��hZ0Kq�0�;��,L�-��7W;��$�ncɽ�-��䀬o�@���0�1�wUr9�5��#�3���.͝~����ql���9,���6��,q~^(����hy)�yjWAr��9Nփ�hТ����m�1��6��Z��(�oq�y�r"'�ڕʓcс8�1�8X�/�̄)����9+��4�A#����<�bT�� ��1�M{�"��E�![^�l�dj�]{��^ا��r�e6��
=P����ާZ>�&�z����D��H�W�����v��ְ��Z|Ɇ{[�f�S ؑ�����!���N�z��v�����䊓&݀�:|�@<�y�o��[&	�G/L����QxP�_��-��۔��L�`.�?��SP�յ�-� ����W�)l��y�M�L��c���p�Q��s�g����e��d�x0qHs̵��Jҟ;��~<m��~@v��b�%.n�+��6�9&���/�)Ҕ�"���b��¡���D���&OF-��%�ݩ+y��yڜ��	&�?mQ�/�|���;�&��QA*_ wx��mo���x�}�!]�.J�� ����6���֌�mn��o�p0RĥӸo��p�C��1@�pt7��稕2�מj����#Aοkz}a�K�ڤ����v����]�ݏ-�qQ�m9Jyml3��M������ω�7��H�!�U�����Y�dh����YT�L�1C����;S�89�v��G3�D1ZC�d���m�E+|��ò-K��I�GR�E3d(�
��;Q1
p@>i�*�e�k%L�G(�ll���N�tX:�$O*����o�R��Jh�M�6�T�(�HM���h[z����S؁����be?d�%s�Ё���r
�꧑=��I
F�d�[����&�ȿ�7L�I�V��;ߟܠ��[䇉�!u��a�ux9@
����NY�:&�S��qo�m��c�^���{m�Rmҫ�P4�� �~o���������f&G�n۾���S/��H �4=Y�S���@���	P���0z�����F%�Z��=yo�W�d�ӣЊPMxK�^�H�,û�T�P�7%Fg�2�~4�Q�MN����ݏ_8j��Sު˂z�9{�ԀZe\w~<�hўr�]��(�U�Ϙg�Ծ�į�g�k�E��J@5-��h9���w.����)�u`��v�f� Չ���r@��6���]�r�����(��m��Χ�U�����8o� ���9po��� I�����M��6��3?�l��?D�BF���7�� I�a�?W�P� ��~��jnN�ߍ`[+j�D�o�'S��c�lJ�.l`T�{�O�\슡ڥ��k��mf3��?0y���5d����@�û�a�M�4D��o-9^�����^����:m��g��l@�zk-	���^����<��z�Ai�L�+�g���kU>���VS$	�v��=:<x d=u��6�hr֐1�I�YE]!�b�x���˫u��T������v��B�T�iv��x��őa'VBGq��ơ����&�clP�㚜t��#(�]�@��d
��tK��@���H�7�Ϡ�۟�����h��+���R�z�\��{�/�k5��`�KKc���gWhl¶M�����:��#=S�P�b2\�@�k�=:��J�c]�v{��7�(�F�#��G5A<	?(}!z�����Z��lN^hz�(��2&�����xwF>9�+B��B;-�A�H%�s��3�jR]�cC�Ҁ�.��Qfy˦��m���{�M[�>u���M�S�tn��G��F�)I��le��k�'f�Bޏ�(�J.�h��.�M���*� �--��}�fr�dy9���M"�|l,d'�݈�9�����|�7>�1�*TG����S7��w�#�Aٷ��FKvts,���8�4���"�d_1��$�A��~'�჉
1��I|g�!�#��Įd���pX�0�]9�E�fhN��~W��	|��ZM��3���55I`�����W���1�q>��6+BD�,���|Bqo��d���9mQZ��M�X�tU�Cd��1<�V���ӫ��LLpj���Jk�/I��F�:��xOY����=����Kvʴ.R��F�ת?wT�H&Ǔ��@)O�\W7S��,���nO��4�M7-iǥ��W����%�Yp��Ä~-��C�	��HLE%�{�Jr��il?���y_�����N����oM��qAQN��%87B:���2y�Q3@A�&n�{+DkK�>���+[�!`�9}L
	������^ur�m�50�4d��*�(�f��KM6�C i�E��	9�r�2�'7�W���F��F�Ξ�hF�

b�!�9f.Cֆ�=ǝz�^M��*R�H.֗�%��1��b�tA�Ag�*.Y��]��'�Vnf �/��^PD���K6���/��P�
(�}�%��m���*M :I�G�U��o�x�0���g�c���$;��(���>��0�w�9v�_E����4�>��kkv�S���H�ő�"W%���'�̎i�+�C�m�N���=8ҋ�˶� ������*M�����������D�>Pc�>�����v/e޾�H-��ϫ�v����`�0gג�m�H5ij4~�V�;��w4C�Ő��{�� T���N���Yग�K ж��Sh�o
�v � �b����\��M����[��t���^���b�����[Q��N�����w����)�pu2y�,��[��T�! �3�2#���k��1��~I���s�"�sw��������2���|�8ea%�*B�"M�P�	��4�� �[��"��E܌	���q�ET��LY�6��s*�/�9��W�U{��`�J����q,���?>;�jGE"�m�%�Q�c%�Up`�?D_bj�j�h8���$Q)���B:x����z��0~�x"A���Ge�
Z���GR8kX�.g�CB��+"`7#!�wJ�s�i=-|I�t���v���&Kc�����g�D�J�~Y-V�0�J�Jk=��-t.-�b�rL��⶷�$�g��"d���+:���3a�������Hy\ }�Lp?8�2� �lҤ7�<�$�V�O�o
��!�/�:`���y�щ|���SZ�
�rk���!0j��J[�7���	���C��O]���E&Uy�r绘���U�5�淄)ǚ�n���$���a}�4�?'̄l �EcN���,Z�6�q^��<(�]�kT�~��!��y�e�֤�޷a�1]�O��C͟�$K��O���j9�xi�mw���ma��#���9��!���%������!�3����?� ����;yVӥzX�bYP{�l��w���N�{��N�P��Ax=���X�u����ӀS�~�F�N٦mG����NE#e9��<8`^�*K��TӺ|9�)�2"�%����T0V�i� ��V�8��Ȍ��V	?�u	�(��b�_i�m���)�X-"$�`qM�NS^ ��+Ç0���`S���E?s)N�����߼��%�����h:[�0�����Q�-��G=o�#|I���X7�#)�����gH��1�;���x]�e�YN�J��}��`_����� ws��
3<���-GF�0�2́$��ӽTw�����Wͪ�MT�T���1}�9�-���ַ���a�;�5T��;�dGc�]���!"�S`ݝ_�lT���j:�8ښG���_i�������U���&ظi� �-��
�o���|E>��<'(w����TFtWEL�C2-��҄їܑvb�T�}U�b���� '�E�H�8B�7s�0>I�ߩ�zDa�j�ԙ|��ݾ��l�|,E/��̻���ͱ�<W�P�'"z�/�'Z��p�n#N$��(����B��C�sOJ�����
g�w����5n�����[^`�=���B��Z˸�����~�ѕ!~�W�l��'��\&�r.'h�X��L��q�Op�S�,`9|<z��<���M�.��f &��W$�I�z_��=�lHs���5w��{]�]Tյ�]�+�3�7������}�[�7��@�3݂���i�7`��%i$��-K�#x�Z۴@����B�6k��8x3�x��?���aK�&�@�}��=E�ڇEv�\ѿ��_!����EMzsq�_�|[A*B.����h�M���0 ��Tx���w} ������O!�$�G-�:�٤��F%}���HˆK8J6���"W����ɏɶ{l0+o-�y`�V��뱨oG�=�]�q��W�ay@��W��my��۴*C.@&q((�ʑ�pb���S����S�*�/ �#�У~���gLG�����t���?�|_���1�⤇}i�S9L�D��ТbH��M�=� (�tbS��UM�����xM�O�b�S�7厭���9�{���@b�N��������G��}�����aif��<b�o�G~�M��:��ؽ�Z�̧pQ/�9�	�,���W����o��%1������|DD���d}�D�எAٴKX��(�$�P؈؋�d��d���qIȴ҉�D�{�����-fa�l� �N��֊e�5bڌ��3�Xb�L�[Ċmr��\M@�*Fm�+
)�h��GI�X��Z�4b^鋳����mٳ�km�_���5\�炂�L��A7�M,+5ɦ�M����@�-�Ɯ.��}9��-Fx/���)s��M �Z�hc�J�^%Q$�P�6�g<;�0?�+=e��L�~�_� �qq~ɦHg	2�P�g���TT{�~os���Q��GbƇ�퇹�v��O�������F�7B^ ������Т�k9x��u=ނ '���12�C�T�.Z�}��?����(�S���6m��m��rs*9�'K������K9/vaH�hP�4���to��`��o�r�zŸȜ��u��!�v@������l��fK��=��֓���d��'����x��C�k�<j��?똳>N�q��э܏CI�����%��$����D��a�{BUb |M��6M��_�8��(�Oђ�!=��F�������s���@'^�4���^�~�R��<�]�zTyY�&���k9K`3^�?/�{���~g&Aп^֢�O�;�3�F_cX(��bE��`~4�p(.��C�d�z'3�}�_�w���Eto/�U��[��0�=zr�ȏ:�*�:ek�~(9�jA6k�F�+'���&\g��w��c�����J��f_��*8�Γ%���d��K�6���߻h9����.z���ĳ��$���&S-�J"d]��x�P�8�z�կ�[��L̟��/������:��o�F\�
��#ZQ-�������AZ< 7e-V�#��Su�F�F���>���ۣ!Y)7����,��O����jc姃J�k�*�Ф:���D@���#9��芽q�hd�jTQ�m��xTo�q��i�ZO�Ӌ��auT��6N�h"�za�+A=��$�P�=���55�3�Mɶ�GR)<j��a�g�2��H���9��>p����?mJ@�Ĝ���)�e���j���	WS_M ������T��ؖ�x��ݭK}��j�(�h�v�n:7:-�ނc�&�X�,INX��
�s�>ڧn~�`V������p*Q<2Y�3���FҞ;o������qo�9`ǹwL¢�o$����Ш�sd�}Ϧ�qk���A^A#����~9%y��(G]��7!������	��K\?�F���/���7�,�� �`��u��&8�ڋ���X%YJ�ъ�ٛ�Z?��d����,nq��C4��I��
ڒ��Yn_9����f]}�?f7�ZH�-ǽ*�ճC�h� |��T ���1�B�W�|�C}������X�^5,FO=��ݑ}@�'�p�y�]���D��L�ր���/
,Sqw�v���Y*����3�?	]�*�8��_cc�:;�۷PP�᠚W�U�#�{��v��~��`�3��u��|���Sѳ�ݼ#Л��&�!{Oxݖ���=�Yx_�DB����A5�n{ԋ�A�cb�s�5���Ĩ���K=I���	�# �lSӬԭ��)�'8nU��7�D���W9Y�q���&���q�)�O�/�)*����E�9nZe��Q��G���k1l:�$�eȣd��OZ��-�YV�!��V:�������CSv� �!b���%A���
_��i�-[s����/� 	��}�T�
�4��H�1���v`�zc���#] \��K46D�<,�������L����p=Sv���fA��|Jz'Dw4Z��f�n�2]bN�p�����eء��r��n�F�R�~:|��� �s����/5�����U�bc�+N�����fJ�|�gP�V�-쉪"R��Fd�#��t�o�?D�=}�3�Wߎ��؎H�뎘�$v�x���p����.l�"���z��h,�K�����/��X�8��ے��zM��Uh?bæ��F�ˬs���T|�a�dWH��S��HO���zB{��6k�BD4��t.ɿ�5��
�79���D���O�$ONK�w����K:�Lpɡ���� �U8G{��Ԟζu 7����f�G��l��Rq�b�E�-p?�`0��B�N҆��4�^�ޓ�t��	��G�S�.���äh������?���kc:�IL5��k�)|A�_Nͬ4H�n��{����M�z�7X��j��t�@�aFwY��S�m���%1�4�M[`|o����4�����+����|֨=�ԕ~�z/�jq�Ց��8*䜒Z��bV6&��ūN'�:3�(|��`-�+����Z�:�A�;�8���A3�:>C%��)z�����ڍ�{�+�,��SMψn�Ry��	�xT��8t3�֘��p�|(����?B���/uJl�;��*����l��}v�Ⱥ��cO�=)A�����#��yK�s"�%�ˍ�d�k-L4�F�R�Hx�0��a�ۨ_�4L�e��Q��pU�>�\2��G~����N�wP�������3y{��"�V�HnxH>�����K�0P:�ïSz �grMg�r�	4hs�+��:���@IπD�V�T�6٢X��ry6��1'q_O��,C&�W�lM��(�e;њw�nF��J�zt�YpN5k���� ?F͈�~�:�i�݌^����K\������z4���n#:��(�xrJYm�K0��*��i��K�8'��vXu�Ye22��|a7/s�`�=�Kn�N�Y�J;���� �"�p.�S�"����U��m�s���n�>gJ��-��n+��r^q� {:�Ŝ����J9L�H�bz��P�Cp;�")��_Xqĩ�ޮaA�}�ّE�8[d�
���e��@䗪3�[�1\uoR�گ���JDs��4�?y�������6���~kQ[���������w�p85J*_�Sf5�CK�"�:Ӭ��T���(�
�B��Y�@eə-�k��9��P�t�ߦZ8�L�$-��5�Z& D9[�*�9O*��sҘZO�6���ЀE��J�pZ�$t���x���� nx#dZ�WEޔ�l�>�y�WC8����	_bQo��xޞxxĽ�X��
odlQ�!X�T�c��9�	nV(W�D�m����v��a��xz�O�1O�L��"�x�Ͻ���!e�V!5`V�6���*�-bԯ���HO���^i�ts�G	[�݋�˪K�:h�u �
� *kAK��d�5D��f��G�K	���EȊ�����?�%ʕӌ� ������+��f>��4�;��y�s�4��S����1�����l���V
R���FO����$�$X>��:��������R�T�ë�R~��3�ƴ�+2E���;��K铨OD^(xs�z)a�[��+�͛A׍�����,w94^����Vڂ�M��{���(�%�>Ô�c���#�8޸���C�ӵ?����un�H
:z=���O�鰂��Eȟ���?7�uLC�����CEr<��^�a�8AX F�bŭ�s%@Ș^{����薹Tq����9�p�t!%���p̰H[⎕�$�#0�%�#%�|��֌�����MB��8>i�]��SS���a����>�W<�"Z�00�#>�V���ܬ��6hX�4�hn��x�����zv1�G�ؓ��k����ϱ�ј�� �۽��,#���~��"v��WR��l=ԧh>�#h݁�3�{٘r?�ﲂ&��^Et�h�N��� =M32�x�8�[�h�τ�a�`/LJS�4z����ԍ�^���!�iw��i�|���$�B�g)�'3��⛜��}��Y�o��J5@�A��4IФ��~G�A�ޓl@�x'o�p��.��&h�����OHV�3�/&"�8��;b�|�o��<�$E.C���m���-wQ����5%\�M����t[�:s�d��ܿ�Y�d�2'��ME�U�C�+w���4�^��4��FdT)�����b��qKMr�B@L��j����Է,�AIU�1�w$sݖ)u�,��@^p ��H����?�DU���c
>���}:A��T6������Yo��)h	��*�\cj��&
p-p��{[	�{�r�ۢ�W��llF+�p�$����7�)�s��Ġ��o�~�d}8���Z����'��x��C��$���zږ� f��85P�+�y�ecI��L���Ǉ\�
9��BO}v�R�A;}�1$�}k�	+������K�u���Ӊ���S2ı��%6�Ӕz��sV�b}_[�Y{W��"��&B�*˖,����J?UX������J���#���������zx-��j	lW�3�Cchn+XxDO*[�`~?��ˢ��m���iG�����|ٸ�8Gb"t�|�N��_�L�b����P,�C�$S��O������;ɓ5{2-w;��%��O��$pz�lFE��~Y`��\��f�i@,���i�R��W#����u��x���y��H���{�[��/y���ng��i�X�g@��}d禓*��b�.]���PɴR@1*R���5����v�.%T�$���"���v]� !���Z��"�l�
�{�.6淥�iD��������������)*��G�dgt�Ļ:�0��
��ʕ~�]����!��+S����B)�i�#�+���H��Z��Z4d
db��i$���`�/k ���;�5{�	��P��2,�mq�����G�+n�/�Er_uyC]L��́7��.}���o�y_��(�k��>���Ѐ���bgr[��0�6���(6��l��� $@�����׻��E�iKݣ�R06��ϵ~��{
������z��CF&P��t��
���Q��U��T}��u��A��5�� �7TYFػ<�_��?_�
A<a���؋ʼ8_�+*�+Χ��̦��yѷ�%����ˏ|gj�ĺ��V�&v4���XbW:����b����&��P��Q�`x喩DC�%��o�Z�|������IA�?)�����p��/l�"�Fv��yk�<+�\��J7Y%��k����`��X��L$��T���a}+��D�r]n���D���fz�@x�k+����>dE�fU���������ti���aI3���L%�q�i��W��?�D�)��2r7Hm��P���;/G�ϳ�LAԸ��)V�����M�J8���ӣ	7F��lkO^]��0�5���T�����zL��%��~���&�z�q����r0��lo ����͍]�8�Ny.��PSJa��
�7��"��A ���8�_}\�&ڭ��M&q�{l���a��3�N!�8|���U.�l�b���&�>��ݫXO%:��>u�F�Q�x��*.���1����܇{!LA)vg�<$RyO��Lѹ�8�N[3zW�u�^9�l�3n	�㺱�|��>ũ�ͭ�f�""�H�1�5O�M���Bc�R�������t�G��_Ez��9�C�aYڥw(�O�����7\���:��`�j����sEμ#2�	Y]� �Ӏ<��lh�B��);|&/��~�����G�|Ø�Dx�&�D�%�7��Z� �u�u��v�H  ��GP�����q�QRV��w�G�n�?I���dAU�S����u+��Ʃ)ӻ'�r�S~Q����-ldÑ�J�^?R�cC����̣Wby�M|�M�b]�j"Źđ�����Z@��ۥ:��o��]_I��V;� ��;�c���KY���(w_�Z�B���AO>�H����r��u��f����ڸ��q���aV� KA�`Z(���(8��v`M<��@��(�F{[�������Tz����,���P�a�$��'��i7^?���,��H��?���L���ˌ���:SZ��a���l�J]�x�y.� #}��$�U	�V<��.�K�P׷�./���-j�� �)~����L5Fy^=�����!Y�E�E���O.�#t�k��O������V^[J� �n4�@䥵�������	�/�-.'_$�[�y�cܧN;;���E/"�J4���l"c���wSs��+���x���QH4F0�S�Y��'���}��@�2HP�s�;����ņ�p�p���;�'�1ĶC(Q�,R���U�+��q%=�#$ <�Y�a����@꧱�3�*2W"+* <t�pj6���I��K�$�X(����CK<����=��Tl��%�� �O�wI`3i="�O���PϲA��E�+cAN��;X���E�.K�OsP�L���9^˧�G�踠}@�J����B����kp�	)U�F%[#};A��p$�4�����0�
���0N�<��Nm����L#{����IƇ��3̖��I͚3���Q�x=Nw���Al�q�3޸9I�
�nC��e��`�/� ��8����Ke���R���G{�X�����|2m�V�LN���HT �]��ViғƢ�.s��ݙ>����;|  �:5`�P��H�f~�l�grL�w�s�ҮG����QO����Mz��/)AI���j��r��2_�K|�Yxv���_&$�alm�hS��s��Y� ܋܄Q&
?���2���J��M�v�+Hv*t[�w��AH��k�)n��f}�7�U:res"��L�>Ԁ7��	ޗZo���~F�J�.<\���n]�+\�*�Ҡl[�aa{��gυ
�Γ����ez�_Չ���yr�E�<*mQ�C��k��,��R�*')�7�x��ҋXsJs�W5c�? ��pi&n6y�>�0���)�%�����G��M�4z<G��y�s{���N-,\<4̂�n'����wG4�j������wƲ6�p�𒂌)S�^���fI�7��o��Lᾛ�x$H��̳"Vu��Z#3�je��|� ������c��!_)Q���`��L�����	�#�&n��RCL�d�5@p>��k���\��j0T=�M�g���0�4~��V��f{��>��
�b�M�2hF����qO�I���?�^4��+�?��Δ�����EsU���z�t�$�t]z��V�m��`;!,�>���1�=t/G1�P�(��
YWף�>��)LE9+�Ԯ��Da.B ?�&8Џ6�w9���0G9�F��D�b�xLuY'ߏn��u};�����%�~��X%[��q�t�ҀL}'�ƁKP��xx��pe�A���=Xg�&���g�+j�rk����F�P��n��ޗ���C-�J�*%��v|p���D�wW9�f���pU1�О�"lE._�<�C�Z.�W��9_���T�IbZG��N�4�K�`vH7�[qWE�du�&�e�ו,f�g�{q�CF�]�@�o��sp�U�&nj6��/�H�Je�I'�怐/�gF�
�[œ�0�N&��3~�)��Y�2��,L�ۛ��]�a~�k:h�#I��E����157�0��F���h3�JI[��F��J���`Y]�.X?��Ώ�~Ρ4i��c�cnWg^к�=�gh���$f�q���W0����s��4�.i�]Ա	6a2��g��9��w~�[�Z|nk�a��t�1go/��8Պ���PL���2^�\7`�r�b��U�m�|�	|�as�cQ�Д.[u���٘,�:�j}���(j�Ǌ��M��k�B6V	$]���/���� ۪߯zeb^N0� �a3��y(�'3�9ұ������ ���G,��������C��<�]d������B�  �����2��P��h!,�ʁM�W4�S�RCA�z;�CidVj߻��K��&�������Ǖ�����_�1���t#� &^a��aJf����{C˚4P�v΂�VP�}�W��e�w�˒HN_��c^�f��)ōZ�T�y�=?�]���JQ��^a	?����bC��Gx4U]��p��xT�X{�Ft�}��,�]j-��?���DWV�3�>zmL�&��9H^�U��<-*�+��O���:e�ʻwe qX���`�!���:0���z0��x��)��F�J�B�uU�ԓ]0�*џ�v��^��4����Gu�ς�'D�/�4�6#���Q�y<Ȥ%�G���*T���:Ä�|P��ZȌ�nŜ&������`��#�%�H����_1�^���-ڳ�@����*;>-i�C��(՘P��_:��v�J3��N����؁����x����U��w��/g=�r��>��m��6��)��ʱB���Ŕd��yt�90��CR�!5���7�P����\�?����-�8�
^rn �4�%)\�!Y���S�>�v0av����ȣX���m`ʸ� yͰ�US2�"(	�p�ê�|C-��pu�<��?`V!\��Z5��8������y�*\�Ix� ##�B�h����!i�?a��q�'OB@�� ��	�Ƨܣ�����g]��̖;�SyOZ"40[��l���VsR3�Z:�0�4�ҟ~�����z
2gU1!��$������kT����c9�=R��x����B�D�18�������/)��Ҫ'owI�#@�(���S���G�V/)����%��nBA��D��_�8�OX��K�rQ�����(6��	�زd�L�%Н���5lJn�o��X�#]R���]ڶ��h!R��m�|��b�G���NԻ���� �=FK]��֫E+�%+I��ˆ��T�#6�k��ƪ$k��[Qt?}5�s����a�k\�Y�ġ������t���������fr�����
w��� 
s��ER;�O�'y�M7י@6V
6����R����j���)�R�V��H e]��|U�J)<��#���� ��g1��@����7-��P�����vܶMu�MO�B���B���إ���F��>�2�k�X���zmX�lױ%B�b���8�"�S��M�#f)7d�+w{P����q�jq���	O�J��87�>1�re��Q[��k9lNyh�?�[�����<�"��L��긆�X�Lbb�q1����ى4-ѓ�b��0˜p�5.�3� �/&�b�o������*�:��ت�*��)�Ȭ��� I�U`���'u��НSso�U�%��W�HcB?�*�:��������~�?�dP�9��f������^�_�o��<��($�맅�-<e����O>Q�tً*�c�P= C�r�ϗ�����y�Z6>��[���*[��[���s�O3	��D"T�?�^d�6�Cm� �l*<A��j�O�I�9:�çƏ�������B�	�MNrw/d�/����]��V�v���g2��H��&�H���V'�/,���dB�Fmh���"6�'����0��Ld��]hǉ��g瀩ϸ&�5)��o��P�{��@^�#�ڊA?	+t�k��C�����9��dX����A�v����&���A���i��� ��aj6��b������<�26#�?��<�Q_``
��|�Qk�bpE-E��h�?<�\�
���F�j׍�{�X�I3�8�P�US	oy141␯N�W�[=_>;��kN����q|�!��}��"�C�g6�G�]�h�\aR��~�-#f,J
�����V�� [;V+z2i�1j�ű�\���hy�R��u�B+�S{R�_A��Fꩨ{��ǧ���uS�<b�(�F\�sn,�S��2��o��/�5*�-�����"L64��{��a	_���!���p�FjW'I����9 wz#�Ӫ�*JU���l{�U���vl?�M�HO�d��4��cW�Mu{o��+)���n�8���0
zQ?V���6ԛg��e<�YֶH&B��������_Ȕ��p���q}�h��6��T�9�N�͈��e�[�A������6h� E�9�RqHm��^�n룕��E>0������eGT��r�7���ಂ�I�&��]�'��ل.�b|4b	|����o�'w��͆���jEN�����/��9��bӇel�p
�I�~����5�&[K	0*�T�/��"�0q���=l�]1 .u�,��ˡV-�:�l�J2>fՁ�S�(�|nΑxN�@�4 ���(H�����o?�M�Ċ�j8g��~);ӝ��؉ r�������ϥ�j�ϣ*j�.�3����5��v���g���r�[بfD�-Ӯ��]�������с�n�G�"����_g���Q�$w���fck�`kU�o���C�㬡پ���FA�O�:���ҏؐsc�<���
s��/��6�4�N�\%&eE��ԕ�(!pN�֫��}���R�,�0��s#�p;�A�G
�D�\�����	R)X3�h�H�����d�#�~�]���7G� �`Jro�� wL��R�T+Ż.��5>�]RW��P��d}D���a[��'� h���a5�"�z�>d�L��X�wOqv5�2]��v�n�i�#�H��X�\�M{�J�ɞD���x��o��X���#�a�8E��~�5P�b�E��V���2��NĈ�w�[1�hF��=H��M0>��-~˷��x�f7��\ge	@�]/B���D�|�%jKϡ��_�{uf�ܹϹd�r���!⣸rr�����(:�W�1X�X��{�8��u�8�s���&k�S���[��(�Q�;�ruM�߽Ě�#Zذ�+9�ŏ�����ɓ��VJ�8��4��i� �(��HB\
g����P7Hq��
)�^U����|#�S`�UǏr{���^�3�|#.{����)��R@���4�t���Y比�6�s��%_k���J�QQ��K7.A}w��+e���<���2�#,���
\8�b�'x�Ĩݵ��NLL՞<7�WL� O�qo��RM�M4��&���� �i�)0f�6�Ϫp_�x����y�%I�)�����Д�2�ʟ�R��8m�l^
@1W^������f����Cل,_�WA{�$l�G����Rjp94�]a7��e��Zt���|*	!m,��}�t�I��)C|�SQ�ړ��`Jk�D��$(���	/8b��P[�#��E���ٮF��u���v�>�1����B}�;CF�<�t��Bl������e�ԍ�M΄lhmd�����s��0�D��=�v��L�D#n3"�d=c�eO�46E�*0�ګ�-1�q	��2*?�[ѕ�Ӽ9j̤֔�x���eQ#K�(l��"��'/���TG:���N#y����h��5�4c�ۖ_uhދ�&��?T�G��ʔ�e��bB?i^αX�:)x'ع�,o��|(
n9�=���r��?b%pu�����Y���oL��UA����)��Ѕ�Sڽ�l����K7�Oun��Y��Lv���ɕ�+V�cΔ�5;�{�����p'��QWbaZ�,�-f���N�� �P`#a#b�� 4oG�t�/��'��@�?q�n��5�wD	�<�|8S�����i�:����i�Y.ۻ�>�_HjyiC?�"t��kR�W�.����S����a�4�1���*���ϰ%�m�M'�Z7�.�&����e!.a�'������$�Vā����edAػ�k��o��n��%�5��q�b�����-r[x�.+��h"����nN🤩�Ԅ�*f|;��>>�nK>5}���~��\���S����##EМ��H�\㎃���ѧ�ڍ}��3
�d�o����a6���@��r�Y�-|�VU���9�h9��Z�Zj�Ը�r{���h�a���ҳ5ֺk@r.���w�EƒK�S�oV;�Q�Q���8�T������\QZ^L������0p,���3��g{��t��s7�|��%}��Ɏ��_7���vT�,I���*�؞��uЛ��t���o��U1�P̡��ܰ�k�s���>�5��w����M�޿��LJ�����K_��z�*ۢ��W�A�S%���8A%}M�r\,?�h�����)&b_�=:�Q���ܬv��)�}K�K��QT�����/` �w\�ޑ��vM����m�t��䘄�ɸg��@" U���r��"D��
Ř�(�c�`Y}ʷ�k��m8`��)^訍D;i1{�$ X���C�4����Rr)�t��罹�'����M��F��I#����N���U�������0�_m�i���h)� ��b�c���0��&���tir���L��$���v�]t����:�+`j*
�� AW�[��ڀ��RCbS��A�4	��@��\�UPX�2f����4t�����6�Qzg�$T)|��TCy��n�Qh%�V�OP'��R�zڹN`�1X��ǩ!W6��O>�;�Bd߻9������貥��-�!鋮�h}�~:���4tg��E��,�r��DŶ��&�����dYg!̦�-�iG�n�q��pw�/g�D�A�~U�m�jnlX��[����K��������o;J�Y3�F������T�u����M�S��g�$��|��Vn9^<�ɐ�D])f��=��w�I�w�غ鋉p�	�^%]-aU�FS,�9<`vC[R<�rd�]W9;��]%5�M�E�9�8�S?�r�ga�t�tО��UD����#B�[Q��KeLJ���T�H�V@5{��9���kG&,�����IP�m&9St��2�[�sĀ�� �-�kx�$�RJtD
Ĉ���]R�� ���r`�#���2�8<��DD\���V3�����8RWV6u�`0%���ˬȫ�����WP�ZH1w��.F�/_�-8�dM�E�L�+��6*t~�\U�����3em����	3�f�z���X�b|BlҞ�����(�sN^`�DG����g 4�D�c���	,�~�P{����@څ�m>V��`]Z����F�<���_����O�s�a�#>w���C��eL;"�o��w8�>��q�aK��N#$�^r 1w����4_��H-7S|C��n��q��� ��-�C����_��?�����ٗC�#S��V9=�e׊6)�1�œ3V!w�NL^	�f4-���HLK=cѳ��*w�@G���(�ue���H�nYW�U �
]�vz�=����ڰm�)uU��\X��n2T�0/R��6r��R���K ��3/v1�D[?��0��=�h-:7����Xv��V��w��d�sc�"�^�Z��BO�NzEk�[�F��r�E��@+�!��O�MՊ�ך��Pc�iz�E.뤲~C�瘜 Y�V�(�g�	2��.�FGv���H�F��2.X%� �X���di��R��Cd��7�d�ܻr����_@�P��Q�?;��r�/s����ԭ�����j��?��|}[�ci�	r��(�ѱ�}�W�s�:Ŕ�,��x+'M(2�."Y�ģJҊi�uW��o��U�mg(�8u_��sc����!1.)�W�|��lD!�ވ���U({��v�iuh��2�����vQ<�B���Ӧ�j0Մz�s�{���"w�u�W�om�$��3AlYKc��t��Dɐ��v&�Y$L�c۶]��l/�>�5j	i���/>S^[w!=ug�+�Gr��±��8b�,�T�a�	_o�9�$�8Uԓ�5M>�i�NpH��؜��eoJR!���Q��A~�q�ogR���Q���q�t�OdFfw� ��s,[ˁbji�+x6ԛ���Z�w[%�9r���sU� 5���`ܬj�Mf�K|�^����B���}�lu�����\��S��M�,����h�:�h�6+�zo�hG���7[f1���`f�#ܿ/�oQS��mN��[�����>�z��-�&�-���8���R�#�	�de�W/b�2��Z�����a:��fb�pG�;IfR�"�h���i6c�{q�sa|��B��q�	#�#E�c�p�'G��!�*�
�|D�'������Sd>�eػѸ�K /&�Ss��I*b1�G,NBq8������n����(5�-�DX��xt,w7�XdR���ⓝt/����c>��$�SE���}XP�!��o"�'}=g3��;�=�k�Xf^�o	�E�È�q��N������ЁlZ��H�{.��O1�>~Q��CH�)=�����.�
�)\����QP3rVY语?�M�����X�ÒQH͗ʧŹ�X�u�.��c(g�0�nl%���X��U���'^c�&V+��]>�t�7�'�>M�j��J��M���l�Y��F����
�*n�>�����XW�����شLæ-��4p��)WXg	��s7�etvKV!����,9�U)hT�Jl͆��OZ�rf����_��ڑ.�4�5u���"e�Z�:| �������������q=�g��v=�RZU�3����He�-9ݱ
�q��.^���(Y.|3M�E"-�8�)���4�|���D9F=�3z5���N0A/&X���(���������9�Kg��2��4js�.��.S��x��1�����z�'�O@�jҍ���na.�)�%��8���xɼ\t[�XO�+9F�P3f0K\4jB\O��)*��# �#�̖�YtKbM���f+���0�Le���l\�Ҋ���!��Mظ3�wx��W��[���0�[aFR��m��d=��������ܭ�5�1R�������Z{��.=��c�ѰL�^ ����h֓Z�����;�09'�':_'��K�ۛ�$�4�8I��+Zz�cm8��y�CW7+vF �xl�w�Im�B�$]�7~�������R�� �'�%�)�ď]�I.��[��G�蛛ɷcJ�i	�A�|Q�B� a��)��}SR�c��+��ԣᗝֿv65���?$�\�o�<�>mȾ��!�y�/3����˻H�Fbe�%�$����B�(�+p1Cj�DhM�����$�b�t�IԶh`hJ]XYP�����w
�.ؖ�R�V�Ȉ� 䢩_�Ӂj[t�����Z`�����q�w�M9�g��5d�'��t�n�a� 9�әol�w��P.���[c��ُ�Q�VA�bN
i�r?��%���g����5�޿(O�-�>H]�?��#�;��m_�>1k�V�X� Y��9Òq|�b9S㛷���{L�h���ߺ�{�8�7���ދ�`�k	�@�C�J�*�>��p�@��m<](&~Oِ��J��J�Z$�,l Aܹ�g��,35�U���.]g����o#�6����tNY#��֚� �k�ڹ��&��0����2��j������:0JՒ��v87ύ���c�������]j��T�F�.T��1y��%ArE�NE�V����$F�'Ѝ옂$���3�i�?e�hXM�w�
$�vA�l8�V�2�L>���o�r�`I�#Խ�Z�	U`�GM��\��t(Ru��:�&�-WR6�$M�(}�]�'���8�^�"�����^?�rg� S�`4�D�ܗ���J�GV��'��@�z{��l��K����NS�F���X�(~�<ڔ�A��oĈ߱g�;�_�L�MҘ�P�x6�F�mȶ�a�����m�h�ceMw���YY0�?��ѓ�&n&���R��6��B)��ܮ��j�a]\�O�\�q�4��:��\#D���ٖ����Mv���)�/a��@+�[�ctJ��Q��H0A�X�MM��ʒ�F�9m}�	`/2V�,�6�U��ed���:��:Ga�G9l��qt��c�~���g�;#6v��߯�J	N��n��yB�1 �gɺ�z;������:�5����25��o����[��Q?R蹶V`�qPv�訮J�>��VH"[7���,�������=qoAў6��Nct�1gV3�$���W��>�,������	Y���vmC_m�߽y�tu�002�Ə����2e�2��%bN!����e�Pn���/��V)w��ii��Y�L�:}7�� �V/TՄ:Z��G
6�ĉ�ހ���V�u�9��V�f�p��rug!�V�q�EmZŹ�1R���=�qC#x�x�{~��)D5[eQ�$	���ZP���-(	`j`&�5�0��PZ�ٖp�,��f�B-Ԏ��
��X���
�xG�YM�0Q���^���#N�lS�a�n/1ot$-�s�]���l�X�P�$T��0�:F���@�|Dx�+JVE�&�2=Q�\�i�����]	���1@��¢�x�8����@��EZ�\�G�
M� �rOކ�a^]?g%3����.ғT��g�qa��s��O���� ���M)�O��z�q
��3$n�^%V�sxȮ8%�mR�c�"]|�B�����*2����m���m3	g�*И����j��1�3I�IiIj����I�S�5��tY������q�U����[#S�p� �BAQq�ĭq0�;(� �VUX����a�xO=���?���n�ܤ� ��Ov���-�����!�o�$@*�9K���\�20�+��
	�C���O,o����ݿ��.q>���=O����������{�@K:$G��Qn�kw��7İ-�^�tf���f��&���:Ra�~�}�����m��|�M�Jd5��:2�+�92��x|@{b�,�I�̻�yt��1λ��/���(�!r�*&���N�{���e��4`΋����dA�_��1�6`m�_,�In�sFP7�|w����Ik�$�_s�nb��T��d��ixcء�AU*B[Vڴ!i��J�>1��wy@ae�z�hwIֺ�X�����J%����DU��&�#HFf&Ֆ�������4ձ�O��e��+�
Կ�Z�
�NZ�+u+{��;�{�������F(��R��;��޼��������o���B��\!�q�9�9=����i�Sb��#�L����ϱ{��!޸kH���I�&5���\�8yk:�!�}R
�I�J���'�xmf���f���v�D�1�]������]�l#��Y�2Ҷ���O�rV.����{���.�o�p��L��a�
�	��P��([Ԕ��A /��&+x:�夾��0���jY�"c]	���8�/�8�O�~��Ć%��dF� ��?���ZԴ��@��sا�6֮%VhiMūo�mfp �;�4sh��|Y���"�sȄ�"�\Z�Y������$'��g����O,�h<1T���ԟ}���s�|!�������邮7ڡ=���q:v����U����F Ц�`|��V��~i�����������2͠g��JF�����\��ow{�QeSNJ�٧�kW�*AC��my�Om1���������ʂ3�(�9�ؖ]?D(��ں�K��e]|7>f�#�Q�K\��b�P�HK��6�@[��U�w��5MX������Ȧ6����
n�y�9��t;sIn�N3�=USؽ�׮*-�Î^����;�׸�`�~
��	�N�M�7E��N�w3�X`3J�R�O�d�=�C8l.��b�K������d���30o�4�"�&B�O$z�!H(1