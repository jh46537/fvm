��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG�`Q�v�E���?ph�Z���x���\� umG]�&�E�	�ڀ𔒃B��]�B�Vh	��'�$��N�$�ů�+��"p��B%��0�KG�-��=�E ���ʠAF���x	x��9��q���s��|%*���AkY�C$�'v����T����;b�^c#�1~	%�%��*�8_�Lc�s�z_50j*��G
ŉ��s�-�sI���LH||11��f��锂��i�l�0㧑��Z ��D}���n�T(��������U���ᤲ/5h\?<�qq��m+���ҍE�=!�G܄����ʌNX��X�G$x������}DK�k�I��ׄZ�A�J/S.���蝟"5����M9C�T���F�t��$$��W�z=�(�8{HٮKa��!rAy��V�!ui���T\�`r,�)J)"�v>4�
v���+ڿ[��T6w'}��C�R����$��0Y!j �<�qd:!�;�V��+*��l\&��R��~i��2�N�BY��������V�7�F,YS�l�ᠿ��?V*�����{��^��ۖ��,�q���`��^��$�h�2W��0	zF_��]��X�
%l��o���@(���Y+�ĩ����-��p�V?�w�ʗ���JA[|(��������Յ�Y3�C^5�ƺ|m�H�(������w��1X��4���j��R��q��QJ�*0b �x��%ׂ��!�^J�X��HxAJ6�"����b>��kj$��Γ���KB#,l롬X�i86�셆#�u9��,"e�&J�L�g)��_��?#7`�w4-z�"��v��\�e������=]�繦A%��e��@��6�����	E�����F�k���CGځ߄1���6n W�e5���*���Y6)^0��>�� x�鏏��=����_�hU�����04�t�n�.�1W�:��a���:r�<�(ՄY��7���
�=�V��N�`\sL�|V�YT]�Q�=R�tf���R#�s�b����䍠ll���d���'��z��rt���;���I�]��yd��=�TҰv� ���	�}����z%]=!;4�([j6�.Uz)�D����٬����gZc�����vt��}"$�#��L�y�����
�\O>� ����O�%L僂�� /�1�\�\P��>�Ct;	�X�yw&�ɢ=��^R3���!�йңn��.���c�i�vhNks}H�w
�nՑ�������-�nF�o��0�|69Aeh�x�ţ�����
`<�0E�}�`�h���]4�g
���8��'�G���4<����|�!H��������� Լ/1��7��K��{��C�JV���{��b}��Nǻ��ni�e�4��ɻ��n�Dm�Y./p+��I�v�'vq��U4�)�7�����2C|��L�v�ʴM�H�dE{�z�������[�&{v��r=�I
��G-���!�O���e<S *��)�uS�� ח�0W��*�!�Eo��U�e��q3��&g�0�{86v-��?�A�A�����O�����Gj� ZL�p��[��S:�v�/1|56]�6���B�o���m8ޅgi%���r�R2Q��}�}�{�2I�ߩN�D�^d��t<��4�)g	4T!m0���b�7�?��[�>�f�U�'�P1����\V�ѡ
ٮ��ϯ�T(���}<��Sc��"�8��C7,hԣ���H�6V ��G���-^�n�2�'B'y�}��̘�MSN-��Q_d곫Em���2���8{X�.�t3Ė_ه�E+�^�8;�_��":oV$��S�@�.���Ε��!1�<�[l��kWQ	�8<@N�h��>��l�N������[�l`Zew�����{2wg�C�w��>ybFgV/)�.x`��\�d�����F<�]��đ�J�B.och�`D*����%���҆S��u.�v�6̦�3���e� ]�J�
�3KH�`,1}�թ��~3Ʀ�F�>(�#<V:�خ�e�O��U[����:�>o�}�����e���:�I��	-־�\�Ϸ wD/8��?I{��`���@�I}-
*?�x�~ۿ?#�����ƾ�����M�"B6�y?N�p�6^�&�|���D3�T��2���lz�(WS@S�*y�9@���$�e�|��DĔ�A)��M!d^o0-���wpU�
&`�8� f�8KL�Z@�4 ��H�(�b/�Y!��?Ad�7������{�ph��x\�ɴ��P�������Y�1�Ea���::��Ö��춒���Ϲ�$K�[YH���`�s�M��<$M�:b�<1��N�`߿�����PH�-�8�Hlfor(��U�]}�E�0�����;A�|1�[��T�S�ԯ���h4?���?�xޏ�%!�$&������+�X`�'2ǎ&LV;u:��b�K�j�FU�Eϥ�X׃�-���k�8�la���+~ �a��?���T�8���/xԩّ\��������,�·�>�󪰜���^��<����5a�Ѡ��- ��[���?�|Q�I�\���A[��nf������N�m�-�f��T���%fcgؓ�f,"���s|06��:v�ӝ��v!^O������7�uB ����\YZ
�}+W��}�z[��NM��L;Y9Z��Wv.O����2�a[Q�I8AO�P �G�=�T�.��4c���`-@�������A_0��3�T��B\�!R0������7D��bE+:����!j�7��֞�Ӂ�&nR��"���'6 ؋7,E뾊�>�s�-1�qm����>r�^�ɩ.�)̞1FFZh����Dbq��9�q`��J�90r�^����#��Zr~���H)䩓���C��(��c��G�D`o1\�N�����x���#�O��j�'s��𓯽fOZ�J�x�A���F�ݱ��/���4��L�g��W��A��.�t �]My��!$�?�+"Z<���e�?�Y���۰T2ɴȸ'�L#�2\(Zo�t{X�`�Q��*1r  )Z��ǒ��j�6�BY9��#�$k���]|�y�\�J �P�řv����JI!��^=�&�J9�W>�I#3ᮒ�k�i��Q��>�N,C2��I���}�~Ǎ6�W�!1Pgut�1:��6$����Z�Hy�%�
TB��fC�}��^y�ja� �	)^�������HT�2F+zfͲ�;�����S���L\؃��%9�vr�P�]�5������	����E���  4f�ʞ���w�В0��;{
d�P��ߚڳc��f�1*IM����Ʋd�",`�����?���3F��+���K~��8Jz7=UX����-��r�~u�;���^�SG,aĞ/�8m�,h�*�`���X}�OQ{����j�E4�AQ @	@]�}�����V!z{CB.��.�������?ܕC(Z76%�n/�9e�M)R��ƍu�&`~e���b��d�C<\�{��L�}�c%;{���/�i���Q��v��i���;A�އ�O2����p�7�h�L�k��)_�+.GQ���*Zx`2-QS��N��=#|����x�|<h�k���6��S�.L���'� ��k��z�>(y+v���n=E&DĽ�qieLo]a���(:",3�$=��;�(�x3er8���pgU���8l�P���wĵ�	����!^e"9>6�Y��90k	��x��c�����ư�9��U��989�a_��^�O�L�ߌ@5��0��㡳/�ъ$����K�p�u�l=�I}z䩑 �L�x����G��e"�F&-����.S��rS�S�$]��T_�Cv���Z�nmK!Ɛ��{��>bm������X�;"w���o0b�K�Ô0�|�ɞ�K6'RV-ۥM�� ��+�Ȃ��/}T?�+�d�aԾ�7��ߒJ~GB&x�֏���>j��8��RJ� �@hX�� S!�4��אG3��X�?�c�v�u=S�{؄�
�%�k���J(zr웏�|_*	�� �G3Kb-t}H�wwu�:��� "����j�|�-p7��XRJ25g�F%��_�d�G����2+:47�{�'�f �JG�sR�
��+]�ڧ���f��̍�� Z�[�b�R�beƸ���
��}�F$i7�e*U���;NZo|K�u��$i���b�7�0��C�n�ʘR�@�E�]�O/�Й���H�-�C
�I���B�����Ff狦�2���)���񿢓4`d!��+^O�)�ZՑ�Z��l|&�=jjc��y}
͠��E���V��j"�o��_v��\�ea<Pd��#�>�lp-�%��#O%.f�X2�}�3?��D"��@ ��S�>u�C��fPw!�B�����@���\L&���P����;Gy��B@ћۻp��f������3���y�y�b�P�v�&���;ћ����y�zB���I�hB�.B��@P��]�*K��6|S�d���u��K�5�߲]SĎ!�)sH�g�$$/�Z�&�%�Hz��R�H��?�#�l�ަ�)��a������8� 	�H�f;n�y�5i���0�j����+J���/ǎ�C�:a�H��K�	�#��U�Ue���F���e|ﲰEU�&�>�����G�8�0G�mG>9����4lJ��	���o)�w�S/r�ֈ$s82�P�L�S@�H���/D�N�@�[q�Q]�Y=����b��ە�(�������:*�?_����젴�ЖT}��hG�O��,��0N���D��,�M�q��ۻ�+�x�,�kג-
�� 3r�c�X]$V��t>���tP�2�P�n+�_:��%����v���z��=�0�	 EFX3=)S�4���D�ִLf�����L�4�d����)m�bM�h����{�r���{'ny�*A�������|W�ÔUK�4�\s���s� 8FYN��C#�&.����ÿ����өg���L��[G���B��e)ߔ/���-n�#��-�oh����Q���[�>F'`^�Z����{��ǎ�pW�����?��c�3:�Y_���/���HU�������xi+8�*�h�.Ǔڏ��Clkr߽���m���w���x��^4�O��/�+�^_��C-�wd^y� `,[�dZS�}��W&8K̖˼�{�4���x�2p�Q�ޙ���N��aM�%_������d�V;H>�z��%l��?�ߘ������5�m��w���W8G��b�Qو��&x�i-5�,[����ę��/���<�G��{�����'T	|l�T�4��ŋ����|�P=�Ab��t �;�qa#%D��Wނ�m2_c����v9?�g�%�EC���E�����v�8w	�u���T-_w�;��<A�����8{20��xf:g*у)fV��Ņ�V����