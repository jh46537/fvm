// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L/oiGMlwu5VKQeBgKE8czvoY7snt+zIOeqSCwk77LYywUpVI1gvJ9CNGoS0Ucurm
WUqlzNjHh6B3CKcDZtNyQ8n1JzSzWyOv+A6hD223Lhx0fECsj9yS61y0c/x4jzQJ
SIMNB3IzmpbvnA+oXqKhX2RKWElkNeTERikRh+q0PXY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8768)
0a6vI5P/B1s/3XVLQF7kqjS5NzqfWJycE2Sr4PY4VKYzD3wbBClYSUjk13PLQRFv
tasr+eV411TkNHs2ysiZnChUiNbbj3Zv5uOmsN5gVxsZyRb1tjEElbZsipnMrliR
vf8QaZni56+cuaoQAoeFr2JUfFIK0EHAZHACfwUNY+TCURaOVk8TN/DvXGXnQB8q
rfcI0uSsXSx4ItrqGmjC3EEXE0Mkc1leFJeIigVhbodDt0SEcpFa+LiscF8apcJy
ogtZg8JSihVSl4jdLXVBf9mndZB7GdkQCI/szk1M6zBHU/KdgSibO+SEO38ZsaEW
83D5+eGRmJ+cNQ4pm8XJ/qkrDvJxlpraF4+zjNLsElOS/uc03cZT0sUvB1sQZ0/u
ogSEJ6wODbU3E117LAIhLz8Lx5WZFDQKsLeqBF7BG9HUbyqEURsr8eRYrVpGUiS2
/RphXljJQVQPl9R8ex7yd5jMaif9erNzWHgC26oJOQ7mtJf6Gzg/N+VTr27wPL58
7GNHrPCZ+xyHOr5oP8UctSl36fmfrEmstwFS8jBm6QpwfZdG2VuoaqZ+vVGGBB4u
93eRZCRs57xuX70BNGkpSwZpg/e+GB7/e94JPx5P1yMAeqDHqCQsgGetEfPAba8X
f6lvNidpZ3LGcxPY6TuXCYH/crNb5DGN4ry8SCVSl1A1agA7ESyekl+itUXBLjAZ
2WlJ9bqqRzy5JRLFWI9HmGBnRIMQ1AnsTXvgy/CeS6gw8jHcx6fWPiTCdJH0t/Dy
fDSodfIMHUGRsBtQ6w45b8o2Bih+D6/s9Cnltv7mS8EbDUESw23YHmvHvpRHdngD
nf+kpnQbF9ol63GafjGguBwBz49QSL0WRM82Ec2VwcMaU1bJ27KQUdxe36zho6eQ
Mty6HsMSQ6F0jr+pr0e7DxAfiG8rgJOfHlRPrYV0MpSrv/iVMj4GqqZkzvTYn7me
FyxmdiPoP4/MOrxuWvoEQkEyQu5Gj5KpHm4Ckphj9GvMAUA2pPSVIXkl+Qvv+B2U
wHwZSsqKPub9pZze/xm8Ot+2VYoBmekkoeq7cuBHF8LrZ2xdByATGbx4+r+RUu0b
30R2l4l8YBoREsG4xJ8W+YQtmqHhsnxZZJE1SnNDISo51bsOyg/W5QnrTJPgs+D+
Lmw+ahmSkb1dJp2B9X1WsMRXwLyZfKzH0Qd9zi7HhcWBdOnwvlwbcs44XEQG/og9
PKq39Iwn6uORiq77tqyigDUj0nn0jqqNYFopPatbjpiLVgeQXjkenkMhRAY+ntxY
+3FFH0vyOpBGafKyLHRHClrCWNq/W6/sbC2yjp22Sfoo0EELTlsy5sjEA51ig20o
BKyXmjipzj/VGWanMvmU0nyg55pKjSTAye9U/87hJ4ir44vzeKRcirfziLPzS5Np
U9mNqZMC6C9kWvJsuQUOyLWDv7GrlwHkzLyHlwYA76SnBLfGxX+eaDfP4M/roZeY
ou9Q2KLAMfHhFNu5pygGSf/yLxzr43OaEz5VHnroJwvq4j5ljEO6ZCbmOmFWojXU
/gWzOTXIRwtvWPQw3DdM719fnv4Nk6ps4r0ksbZtO834Z3UWdE0F9pVT+QIkcsk8
l1Jb0Tk5YWkyb8JJUD6R6/+mDe6jidh7qEUUwXulQmystKW9g7gunapEjakMaFQk
7vr6jdVYDPTOwfixVcciXMpw0L/RoFtIN2Nboe1Lqo7VkboFM03nppw1wCEotjFX
LLVrH6sLDz+2M/B3eCP+L7mmphsT+0M7q25WDdw398qwxOKM31gZefREBY1CV9/b
oBvHmF83UAfvQZXzd/GUIpw+6zhsnGDrF5GFjmuhorGAvtxhRlA9/yVh4a81KOpD
kU1rszDDRjmZ1objlm44DOXnuyUYF/54NAr5ErjrXJC3Xp61d0kq82iCRtVSIIa8
RlwDROdNaKsNnnpRw1di11cplE5+NSZ4fFd+fXnx9RMJTf7QePVDxwDPdY+J7sth
rAlJ/7kjpPP1X7IEPDAfJZ/zrdKIl/Fnc3mLNzRiPA5fYGvOfs1Vez8jhnRlp05n
VZ2RGFsebMmNDC2OG1QKLDW1ej63QZmq/lBjxKk5Oz3EaDtJHSd6mBnC6JYdgTpp
iHjWsOC93OgdNNtZmqUh3AcrpJ8+BGXvUaLdRyWKjWXQ+By14TeFYliUBfClN8Am
0fisbU9mDTqEyQ/unJUxawGVbUdvDRyZGFpY9vzzgIntjjGt6CxjaClPeEkx9vIZ
YBLBM0f3kg8b5LZZJy2RDLIZ3f/0vBYxE2KTA4702X13mqjRfxSPOpR5SHesqnji
wUEjYy5QoP16kEz9b2lkX7CUFvmY+FAbY1iIyb43yJItrTJEUKmOQNN6Yw0awX4e
zRUMrCrFJu4+IRhdUGK+Kk8djPPAtiXFNlQr9fwXFHzmf7XghwZgUYwftGrPR7Kr
40VebMLsIlIM8joK/qIVXkhlvs+C6yVpWJTJ7pwrsjfxcjfaJlQt14DWr3+kuZU6
SOkiSIjTc6+iQK/xh9s51kkqYIn59i2oz4Kc/U8GFpvm5jCaaPxjwGj/S2mJb4m4
R9v0P/glhIzhhR9TjvqjeW1x0mwAdm7tKGbpPt0+Wnn7bFRiskv2CFYE+dN27YCx
a+PCcgznUC3znSPH+VQaquH2Lx4FM7LNtPL3X48hxUcowsAaEJHI0tbqZd2D7eLH
Vyau2OuthY/I/awvs2YJmvenYRJxu8vP6ZPDqOien3zrwZPOsX0+/tCNp+8gFeeA
iI4msQqWzT4xyQNGeY+1vfqo4Oonq45XuMM7i9xj3VWN83YqJqYz6dx56/6zOTGb
jhVeu1leXkqjoci0HmovNx2Ck05c0byCcDF1q8A1GnjhCOMZq8JfreT3kDel2xEt
/SCGkDYXC30/QDh74Deuhf5cO2qH0QS/77o/Jfa8IKZs7fYUBYKXBeVxUqXsf+Xi
QnyHKaYWP+ZG0oP7hevAcqrS878u+z8esqXwyeRlCEUruAvIG434JEwbkMh3k/0e
KmOE/YTXv78ZAgaa/EEG/r75akZS3lSKIWhOgjBmAALRgQMV73DbrxSrBCem465l
+Adtz3snH2EfRaXAvEJOMtSBINvtxQ1tYM/nACqsajrmtoS7LxDorTHnFsCw/vkB
A7+AftJHdlW10IrZo0KrD+oEYNbeYCzGWCXW0JriPjExm9HmH3pJAXrb6dq3sj5h
+7wqBGHiQNED26qhPRXJN7YQ2YGesAYkYSiF9z1UzMDYI6j53jC9fHMP36hcKa2L
o8wEo4hgw2m7d11UHX6y20fU+xQL5LAC2sNOMSFQraqPHC4/6kjfELfHWer3MvFj
X6m5VA8QslH9n9mR+QYU86hSkd8+d2OXhNdh68YNlhLk3B4vn8TKm6sF3d4WYRBK
N6Z5/Emqa6jcD10JeWniwSqFHx52gp9Pgi/39OI2+Di5A2HJRqEfgImmdQQ84ShD
3vFHOkD832kdXC1NJIf6lBJHsRmjRtoHpil0jGeUvpFc0jmlDvmfmfEi+CCHny6q
pIkqxQnLUDul+3PS/9VuzsB/3zH0L6lcZRfTe3AZw0HoLK4cIBkZiIb98Hugd0vp
vKgL47zc+PpIhIcCZlegU1ABhnf4yBxKyPi26bXexw2GZbmi4L5wiZ/ZIWs6YCBo
J2RBY4zKfpM/7Qeyswul/JCziUTva166HDt+s6sXnbiFWTjDC35IiLveIpx0hosq
PJ5zFrsXpXGkqz3AP7X3/l6mZ13B7ectHP2vTMEoyxLE05q7QIuT5JXl7D7pmD0U
Y48tD/0Z/mu3787xopFk946/Wjmi877nXD3dpPz3diEIhWvHrX+THFt39RXQuEil
vOfdMvjXymmzFz/GmIEGbjb1FUwcwdZXBooj0EJetjePlaRdpAudBFg5zqZD57Us
Bwp4ZI9kbQBmM8vUUOP4Oj4/7J0uRJ8yJKd/gr87ubrArPxqNueidV7HhJP9u6zr
YdFPOtbW6axOKE0V7qX8KmWKegXqcpB+LC5lBYAU5vGVYk8bPe4Vf1B6hbqxU29o
FfGW2Veda2lkUkNG9YT2/J1/TszQpDV+/269bwA+M2Zl5kWi3sChwLxSP5H9soOB
TZCWUM1cvGh5TaBqMx7afTYB+AnyPVMztusnSlT/4T8d5PDvXXi3xuvJS4WQu7Kg
xUwZuGYiphGQPwfCmNnP3HL5Uw0fSNA4meK61UuCKm4xF/xdQno1n/art0/87GM7
D9a++oBJCq3mhklBLoF6ArYQa7opgDsEbhIE5Gw7TfZJsPpQiqxYNPrdV+XmgcqJ
k6bgZqC2eAA7XPLd3FW7RgOaIHJJqtBZZNd9EFcJ8EOrCBrCulMDvMg//3n/C2j8
EGhGttUFgkzXBScT7Hw+TrXBPMLXXzeBYIFxJfCcp6G0BI96k0c5yaazk+wzvQ2a
3IQA6RbYNl2TLLxQPeSo/DBijnIe0TLN2DliSjABkrtdm+sHN1LtU1qvOZzMsm2s
yCFV4n/IOcw4R4sDUZyHYCEouG708SQirzCK5bQkh+rwAGP5NCav29LkRl/0CtRK
qawsWZ3Jio4ZhWlJGzIboQDeMqNd1AMx+L55v+M/LFtg+AWRWL9z6B2kWd6K6nrD
mLsy3WNVo9Ps/Xjjoi/s8BCPEd0ZQwlZNssI6EWr0yasv7U7NpYjDrgCvL0XG4ye
qjcbm2f5CReqzpFmGeMclaCU2Hjt4/lE7grNF2dzhrAji02uh38oUPuVGBEJtUPz
3gkRG0Cz/AIgc3VDaKSpZEracx8Nzpw5SZ9wJ5Wh4qcetvciMugLcicvQx42072e
ZJKVpMNzT/eFG454ybXo3FJZ2c6jvgGigcgpV7C3iV4c6dvmGFWb2mGCRw0AIVPs
LmZ30ozrtfPWAv+5g/k2bZ4QvoXsRzd9nxLMdN0k5nNribhxODS4o8sG7Vbh2Dds
nT3OrPckWtNpL8mdFF+QEcPrveaWoOzqWatOkxAweEbxdFfjXIHguSThsWdDmoKS
Ojtw/u2m6hDKWTM/aPzabZrxbu2+gBlKXjTI2KmWeM64ejfoLZIpAjuhCSQ/AvtG
bW9YNYvG2wW8pRRiKb1Bp3swx6c2PPcLU8ljxBzkBtZncYhfk+vF8jsDYBNGeUpE
lvyi4CgEtrXJtSyDX3hz7wsSnj5cqRFSpEFjfOnPQU0Fb+wBFaCXglk8WiBoHh7W
NLcpis116W0KsqeQL2FyIZ9qGkxvzMHdIB4jIexIWUh9kjYv8ghplfyNOk0jWruw
vXyZm/sT+t1GNYT0n914WBiFLetDPqkbOqDnhqPRmHnCwTSJbhxvnjKqvVDjXh+8
gDVCOMrILYfq40BncQMaEgOIxIFSeKefpKV42b2zUJsg6Cw2KmzCVP9RjOCcTkfD
ZFTYdzqtpIIJEpac7UOSv9WEirWCP+doMoQV3GYTP8X0BPXd/4vfL6toUW7dnpU7
7hpvsNYnWQTmd5ihWLbi61GVqa6O2fMHO0aroGDd+5f9Ju5fTdD7j3UbKyofsOrj
14iVEMmgjnE3PJ4UMqYmEPYwzyX9Xa0Kq5UKs/MbA0JmK62tUn2WUpB7XupTTjXx
z18TYrAZrtNwjFrXuxcgIEAT72Z6uUgms7LwdkVkUA+45YK32A5odJMq/JAYVX+p
c6yf/Ufx829ys1O4MOEOz9hw8ohDFXUcYNUWtaDmw9rObZzrnNA5bn00QgU+HjmJ
nnwuX1LnVPkDLrSDsnHlNjBpoKwm4nc1r6/h4hRvOXK/YeV5+QCu+OKu5xD6Zg8P
yAmouQ27SlfDFQnT4xiIU9t+80RBqQE5aiwlBh5Ws178vcDXc8QxQrwa55HxGrol
Zo+K7dAtY5pw3Bn0Epe/+2+NM/tmWb3eLon1+G5dxg+jEUBqNlk5zgX+hEtk4dIS
iqQvYPC9o6zN6BWi40PDLAEJwS2/+9RgackuHQP0wuosE6sIR+sacRH+DeV3j+1b
XwxjbCzDY3bXQbNX/Ul1cGeKOu0w+GohYSfezoNSQ57i6dP3vg1PjXjTdqgnyyA5
6/Ysh4SJJHzYL57uFEH48bamdnd1yvBnuwpJZkGLX2wlwVhiyQnef6a6AOjE4WxH
g5lq+6w75zS8arBRWd8G4DL+RoRnWn0XIe7SiFc/2fZScgSBkrHYRgptM4YQlblw
USev8Xo64NejKPSphNacjVlHEUHXbjckqtx4S6Tvm3f/XkgTw4hplkQ8+rmJW9rX
TjhtfX6fEm6f8YxCc10pFJmvxSlRneRn14vsm/n55MYI/GdnxehnyhgWQrnIcz2L
wyvcORL/YUrCWt8vPg9sOKVmoOTOQ/5wtW4Y6rcAY8I4d8O9wWLAHTbklplBddm7
/W5m60nySZrfMWcIPvsKXuPC0hqtRC7HMKgnTDRzYKRRnnLQzreBk0Utm2AKyzd7
GdN59Sx+IUtFXATPVwogq9trBo843FSP1C3TQm+ydMJmMXukJbF2kBU5IB/q1yO6
FDL5E5rrxESpUTZOZBtuh8mP59esnQ/QekqZdp83g4VNjUIeMRUGZStk7+vEqxGu
DAzbI8AoVVdZjBPCzzPNU1WQ7j21kxk9M2gFqOZQnA060wI8RucVCrEq4WjKYg2x
EFAc1LVAoxjNNL/h08F67V8gb37V4mpISEo23CwtLG7gQFOTpm7SUIEMtcduY5GE
UHfQCR56Hdc+YIn/rV4FkvNS7f1/mJWIHBxZPh8wy5sve/sCLWzVaxcS2+U5yyXp
LxgMK9ImO7zQC3vMAizLHI8mLh4MDR4CKDivCBKf+/DE1EgeOIvFFgnKIiovQ894
ixSLMIAyJ17vuBnCzkyuZQog297MHfiv/eqGyO7aeQsC5mzri3NSAb3u7OiWqUmP
lqPx2z4+wxsbwMjp4F+ArXiSAxz8FS5OOJzTCJr2rJERb2/IX+4exLfk1GUqLY3y
ksjV3w9Bk0cCq/qkdOUtY9AZkYlSamsfhTuGDqC4P38JPUmjGcOQDO1TYCa7jbmL
Bc9F8f9Y0QGH6U4G5jxsqOSunVj8CecaXNtI1dNnwWmS2eOoK626R0uBfW8ttihd
JorJQzy3fry/iSPZKtLlWl08+14qWFcMRljvEgRCLEIzCZ08oMSkPVrTQnCWhD3F
sz49SgFDbaa7x++yT3O82eahT/K25dhlVaSEMBoA7g0eTakZhbP4LjzzR5MOZ4J/
IOoChGIB4mo6Qg7LI2OnbQE1gpER0adtgqXIW+U1gvYq1lSQ0lQav/yB8D8P7SO+
4ieh6Z7g4BbRjOhGZwvY/vfQ6NpLhFDPy1TUFGOOpYNoqttLEbpsoJ/fJSr4DTGD
APCHTJ8tk9w09U7JSypLPbljf9VdwYDTwjIV2LdCcAxs2FsRwVXcTb53QzkTOI6Z
0ipwJmFKAH356XbjQhw6v+KITPoNnuw5WL3uGWhVh2C5Z2qQflZC1x7N5K+CMC40
ER5Q1yLiPyIeQwdpeg2KGvt31zf/cum0MHeL5kxnveTtNTAIXRAdYgabMEiJdWL1
jIGiqULMPuEiEdpo0FtgbrAgojsadJ9PZRtOsiXU3xpHuYsuinQjddKv+rvAcfHI
7SNPny6VpMt6KLGoM+czsEYDf0XMqYqbtrDefUTcPkhP5DeRpmkapE3//SEYISTv
J3NVUeiK2JiYtqn2fhCBB4F41IGiURF/WTv8qNT8rbbCjwFWTFM7UIE1M7zskMyF
qdSJBVH5FuOxhJiRl3pwD5lzs3i+79iuX+XTpavU+4luteQYUxL77tTxfkdPKo4q
ZQvS7HvhoT/feIb9lGf/J/4RdEwyHhrYP0ti/JQHZ4+8QKBGk76D1cQh9Y4Op2MG
8FK8Y2Zb2+tIHDLdpS709Kv0Yzbo8WNW6+Ggj1kGGREjcLUCkLn2SdHwLHEqJOZo
1rK9fACNxWi/sYT/df9vgBWRw6cKoH1ZY6XfsdPBffNVDnlQUCr3MVJeUPrpPxhz
Fmi2cT0hCoATNiHanB7lJ+Gv6zpeMCmruW7CDG8exOKE5tUBZyibPz9IK9vHZKD9
0VlP4F/8+YI4PtSfgssu2WXiO08u23GrlPL2UsHpYUfsh2zNuKlGUEFSWh9zUMbz
Qf1/t/EKO16ZeyzXTUQ0rW830E2tb1BR8R+25ZnUKVONtfSaQamWx3cKyY1veZz5
1CtiG+PuoqsQrN4hRBixpDNakmJi5Ffy0GNcbBV83Mh0ExHwkv7c6HdFpMv94q/c
XXReR7sp4weHffzuldZlAUaM3BcG5LXz4pbuS5Oj0rHfiruDsR9ZPTQRVk170MDk
gg87kwdHCAzYeDThTwy+qF+xRIyvcjCObLAn1RohrIp9HQqlw+Ho0Xv5b1TL18k6
f6hrgnhRbCxO9u0KtGrNqsh37TzsG8vcpApnZ60DA0IWRN/PtZctompmGSbkzJnJ
Qt6d6ro1a6hFs3zko+lsCgKaTmt15dyp6SQ14tBfjgAfAnxmFHmBy2wNdakkiQAc
S2DDlNwueN2d6k9jKlTPanoSbq765Xk+nU9p/fhPxKBEoFlWQvJ+pjTFSRUoXOT0
Ake4ZKAVkDLQic8QyLfxe0o64k5DZnTqvBkT7JZka+cQZGnE5hwt3PdZv99afDDz
c0yH9QSIlbuQSK7CCs+6Ufm2JuHcWmI3X/2dCtzJJVYThxWUEy3nkT4VC90ZEdks
fAnZNvzjB3RrPUSYX+FGdyQuH3q0Z2Fh79AxWtWxIsqwGSKOF5xvqW3x5QA0WXkc
EF1W/u7uwZbaeTr1ipvGwvXUpzQy1BtL7ADV+/siwEEypRp6Y8RKO3sEnJNPxy8h
atXAoxH/kKbFL3riSr8KI4lJJk6CulRedgv1gPEiU8RO9qi+nIcupq2CCVGDh0GA
Z8RmELA8sljQcH5gyfUcEtcHw/3v4/xVLwE8YxohaY50Umx/yksymeJTgCY+Af9U
JbKkCat3jhr/RI061vuc4H7CmiEK+VnLGa+mjXN2VNeqRndQsn7uEn4h9bUHLt+m
USOdVcvxo1/fCtof/mNGKxJeDsWXP6eKDdQCylG/AMYt64pEZSTLyZkIxzQvQ6jH
PpajuKyLuyAgauiYwsAFMbsE4Ve/d/EmK0s4nRALOgH6ZhLop+FjSY27g0FnWrjd
49ZijXNmjWfE/IxmQof9CZaPt9QSYBtqjk3sDnO9ZA/gAKfDBHvmhai0rpOuAMvD
N6rojAcNph7+xfrTDGPOY+t/LxcMaqzKRtXgPgGgwywWOBOAikl+jct0hDYV6cHi
xPqZSB3AU5X7dQMTz3aR8pzRpgZxkHBfyCY4hPGwgyMDzeSj7KYy56pfQw1Vtoe3
tJuZFrYir4wpDoFJ1f3PCyrtrdZvMevOVhmoyui7+QKK4XaYd74EyxIURB6ZRn3N
GAYBrBtTEBcNT9AAqE6SydMKWt/reFckKa/nHea9XodfASQMMF5WbC0LjPYfEg7Q
yLETGattDuk+x9BddQaiby2eZE2UFocRxLsVkilk3exO8s5NpXg35oCVOTDrmHlM
+qJ1zW9FJ58Yb03EHIrkpNXx5H8iQ4nAWO3T0/RcZtykd9Kvmb5jgvgFNbaq4s/j
c71GUlSCctdbpd1aNAFfuk5QC7v5TF3dqP7V4PkOLwrTHGWjGf8gkaq6xqGZk/GK
3FwxLsQt9RfCee6SIErKl1d+LBkX6WFu2M63CI1fXGtqdjVlxcOI9UWKcviaZlof
P2QFhZiD4/+YbOLXVast3Kk/fsJ4Q1WEXAkVXK6yqq9TH45VYH0wv7GIm7JECpRR
r58tBuinro5s85NnTogCyFeNuskXBgnv+baeLsUA0wycUGQu3jnLF1G797pPgk+M
MxOBjD7VJeJen2WXL9e2hlrZsF17+mftDYis3uzz5jiNpEeDM7uWSGZZtp+/mtjL
gGerxg1V9UdPDk7dB89P7qxkpVMSSKFwdT3S4qYHwwb/4K7EivrGQTWaxRKmuwXP
GvkqdLbBvRjIJGOzML4yfsvXpPp4ywQLbXpIkvd4GAq6cR0YFqtMJWl4MwM+GJ9g
hpi7LHdfgnD0hRi77V/34/5+8lfWgldRZNmDQyWhB+WPhNcQ7UNz8BGM+kDVO1kV
GwG0Qy/ukvWkONJWsD74fugZpMPn8NIYM3tXQjrR1TQqmT8cmQvXDiCyt20/Etra
RUWKd8XmIT+K26RoY2QWtQMbmom8rU0eMDF/TaYKGgas67FFRjkERvJBQEAk56Zv
l7XLlKkXyabgmcUsl9xdBYkAkxiyMbX8pKcTWQkHrBBe3XDyOwPDa/SfWi32UwWf
xuEtHHUUgTWoViPx+hpVfAfaVIlR7fveZU4DEEnZpjHsRyqDUdaLT9VUC/vBczH+
KBiGbLhw0AMuXZtvuAzhp1InPjlXMFI13+YEJoC9n916lpx1B+AWMegRJHw3sHgn
ZtcY4sQbM/wYSvHCBQlk94Sbo3MtAzL81D1WSEuJ/oT92jr7h47QArliE74tqm1M
FVBVIorSDrTyVlXpJDaefpFmce7yyhe1Fforg2+WvhMiZyPGvvGshYprYMYd31Pu
eQx7boThc3Fuh6woYBrYCtWwwpQ+XM0zMMYuy8IkMZGBT9/Rxw3FMEITlyuUKl0Q
LVc6pyYHOZl/lAm0BEmHtjvhwWy1Ird1D9plCRx1MvEOeaYar1goOsOemGJv9Qne
rBeNgypwnqXNwVRjKzMkahT/QbtMDytyUHbvc6xFnmhcq55xOidQHTlmLcifJiFx
179s0aJ7mdyrHjaKGyoKm2J6+Zm/9WlyozA/Y9pf7ZPN6zizisWbwskUq+qxviPQ
rMDrarIeCqMl5ichvkGhIAeyEqM1S08DNslaefayLIJUnNbPFFW+z/zk/IeHVmKr
M4eOH3dNO9bfFwI7i7U7iELynzKSptlfoqbgW41w5p9ZTp5uUeWwFXmEDjpNZOKU
G69+Y/4EJgMM1JYUAvFTwzwc+n44SvYWlOveYg7BJWSOIueQvV2zQhUE+/4bsqdn
IvmvFJBAtr2fuuYd9TLv6GUwUCZd79yZDvNBDJMgImaFhf80R9fbLjjry0sjB+YT
eRgVab/I+Ige9xzVJVcawMp/9DJbzOujbMvt1NspFwbwSPC4Ipa3+unc5UYpryie
MH6mhSGflWGpxoppe4wNhFi7q/dzaWzsGIeEngZG2EOKSWUd4mxLN7mzPfOCcJyo
OGJhWbz6lubhbFGYC8Bxcup5Q/uYbMT6SVKRt2LvzwReAxkydqUI5vktIlggQ7Hl
8Z+LxfR4Iqp3hi3oXMtUjki2R4Db5vTV7Zp/0vWHE0bkOVBFVh7hmMIJa7Cl8sNz
XvvukEc0O+RdF4DYUih3LdzZ1z8zO/Y0B69OUr8Y1EVy/zSiCWnzcW1aqI0rbXo8
d9XVzPwoRHOdAmuAHayQzlhi2baBD5ntdpU9wGUe55AvqlX2AF0EAtjGoFr5s8aD
IbCeREziNrnKRj6+7ciYdW/NbEpbdDI22OdwEsbK4YvdvWW1T6HaZ5pcGoD/Ee2N
WhyjpxiCUvx+2X6BsNHoQalnYAGciQ5aUF10pu4kUQWCBQMMqzfeinplS4yCHyW5
KdTuGPFzZuCS0pvx1BFaFcYjfsE5dEl3ng4ufdldBBdzhLVKGgM8AuT9/7IUboXx
XGTtBAOHThgemRUHJPkMR9rlOrGYggGosaDbcopu97BeZ+4rroRq2eicJf2+RSsc
zlHCq0G071zHDFAcpb6DuKHzaZ4IGdwY7LM7c6+ilR8=
`pragma protect end_protected
