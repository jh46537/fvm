��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(|����	t!����YXRe�������U݈�NׂI��h� cw����X�`��\���� �o�H�RLҹ�%��!��*�}�\���&�!Ԃ�0�K�~�B&�p'�=y�wV<'���PH�y\�^'��Y�����������D�x� :
�$�<�W�%�������=\IX�xTSa�n���3�q���$��H�k�X�������(V(U��L���ٲެQCE�v�6�m�C��7�䬷iW�E_߬Z¸�f��G=��E;��Qc�dg�clE{��#�c�T��DV3[�=� ���w�	��,���̏��i�׷�^�v�/��t�rM#�5{S��pͤZ�66&-�º�E8��GhE��Z ^����V�x�)I(���y�y�*����J]@�r�������n+~]��k�b|6� Ӑٿ*)L�4��cx�/������e"ѝ�1
@��
�M�堣%��J�J��R�)�{Q�'����`9x���1�M{�G���=��ԪA�f�%�����}���C{���҅�ʹ����YT��	�.B�}�
��<�69gq�Xf�� S�r
4{��[��e�KC1�)��Ky�s3e�S����Ϣ�v��{Q$��׹�o��~���9
t�[���3֖+f
�O�� �����`���s��\�>�KK��ٮ�$���0iC������Il�����ݵ��h�R����:W�$Z�w�m#I�����\���2H�7��f6��-^o�)qx�<H�b�ח��:����SH�+��b�l���l�ß���t��P���S� Z�w顶-�I�ϴC]����o����9�o�1��Ϻ�M�o��͊Λ��o�S��Gy
�c���Y�S$S�É���=��[�`�v���h��eٱET�Ư���D���o+��'/�ㆇ*���o�<8ty�s�c�Ch��2'n���ل��qv���З�.c����&�D�:U��[#���5�n��Q����c��[���;yL��Ux�*��lp4kQ�H:��\ZA��,�m�=h)�A����y��� ��H<`���3q�_4�L{r�b��7h^y�٬O`���v#�r���}�Ԋ��M����%�N������[���}�Sަ��FUׅ<]�c��=aʯ�qS4�/"�0�'���w������e�ApK�\G-�2-L���Ilx��	����Za�}Yb�@��"�.)�+E�	B�W=�yQ��OJ@^�Kj����flL�N4��9��H@�zڟ�r~��B���O���c�Hvx��7X�˳��k#����ب𘜠��-l�0�*1��J��_��@(��<U!.Q�^}��r���E�ˣ.BXL�����u�t�s��w�������i�w��@����mzTT�Y�e`�P�p�dʖS��D���t���4�eHE2o�V�wb}���Q6
0,a٤^�c<�Y�8�h]�h3#CX���Qk��H��d�1%�ne�RX˗�*�����*�c��=%�i��͗pg����A
��Ĵ�y4[;�e�_��O�;-G��>�m�%�L!����ŕ#��~���-�L���:~�m�x-��t� ���w?�!D�Z$�S�;��
V�������$'���:��\�+C)�d���2�<�		����)�g4�*�Q��5�eI���id!��t�W�Hi��"����^h�G�L��ᢑw�)BEA����d_�ɣ9_�4��R%B�6�:3���#{���2ó���lgɹv�pQ�t���0p��=��_c��r���TP�}�2Įէ��0���S�=@�^��eЗ�F���=�y��D5V�B�b`Z����GvgC�Hx3A��{�7��j�x�~���l5�M-k}��y5h��,�[/46S���`R�3�Ôr�B�12}>��|�Gl4��ӥ:�h�.�!b\f����w�f����4�f�j��a�,� �� @bD�+W�#J�r9٤��/�-$� ��j��#���):�KFM(z����8\z��IK5�_^���s3���}W<���m�s��j=Ծ�4��&�lLd�����k5D����s�[�xda�TP��zPK���;n�<�M)����')��{KƁ~��I�v���l�翄��iq.�':O�Y�1f��������T�&��Rވ��ނ�'�\$���A޲G=#)e�PP,��)��ds�F?[�C>�!��؋=��+m�@ʵ]����LĘ��_���;�f�ۖ�7���/���C�Q����5�Ū�����@��⢮�
K8�/���]D��=�p���*"�E/�E��,c|� �#�'_#$-7�S��f��l[*����[������C"��$`VeIuR�OƮ+8�?��0[`����~Jm&��\�@���~A�3�R�4h�%$.UI�����m_Z�:�9��e��>A�Kƞ��;���^"#I�R�9�>S�)9�?7��(�a��]L0���X�R�� �K�T*�(����7���Ͻ5?πP�<*�]���by���p�(�Y%��?��[g��`���ʹ)N�g�Eof�k�{��Z�v�9��rdY���	��#�Mc��6�(o�;1P�WOA_�?��_*N�;�])�Z���-�N�g@�;0�e��8˂��.�����674 \#� �\ɏ����V���CO��63����W�ghM�a�mE(��wdTi���'"=l����>�{�dv��q�}o�s��K$�`�d����ap#��ړ�Qr����"B>N��+&���;�˼k$2�ˊq=댅jw�h@Zg`���<9�*�����d罹a_|��������2�+�ؘ��Rہ�Xw>ID5l�!����>P�z4��̆�;���
*Z
v�-�v�{�ZV�����Kv��?���Ky@R耙y����\��l\Sp�x��sspس#V� T�/ew{G���%���~�ʜc-b��c�@94���*q�_�2⯮�U6���G�2I9�z��z8�DؠXb��q%������ `�ڭ�P��Q�P= �g�9���`Ja�R��X��&�A��I���k��KIEk^���vb�$���8-Bp���cf�{��ݮ��O�:^]9*	���)���.�a:��Me�A�.3���UR�Sp��r�+F�sM�2牟�nr�WK��x3'��Dr��Uy���lTqM���یB�����Z����taN����"�*���/�ޑVy��yLS.JH#>�Q��\���ulr���MϪ3���U�Y,L߾{V����=u�f��>���Y��R��TqG�9�Џ�1��u9&L�*��z-�{�\T����ͪ)�����h��L �_̥%�H����h	0��q�{X�J'>�8��5E(��0]@���F��R˙�`��,���Q��~o�2�E�� ��kkЯb���;�D�^�X���������3�l� ��^M�c���
6�j��s^.�Oc�k�& '���.��V���9n��&|�2@��q<B���zR.\r��2A�p��� 6l�0�B�� ���`�H�gxv|]�{&�QJ�I0ʢ9�,�#��5� �/�/��}v	FJ�'[��������`��^�[Ԅ�L&m�z��R���U͆H��tb~��C�d��Ꚇ��׆��K�w��tl�sQ��w���Y������Z��`h_�C�pC��/o��;��e���;c�;���X ��GP�%?#
�B`���ss.��ST(7�Um印b�vT�EM��<��d {�
���`^�5�h�����oFD2��+Ġ��}2�`K-80�A"�fTf�+�N �����4�Mߕ����|6�����5i�Rt%Z�c����B{�Z���Zu��>��{�O1�6 �TzY\�>�~ Kgr�-���3v�L�����C���0�@Z��\�r�-J0x�B�#��r���R1{
݌n�h��
f\@����ϗ%匣����d���6�;��B{�7�$R�D�u��(�WL���fm�|���.�ǣ�w+�َB���/�7$��r��
|�Yo 鼨�%�yآ��M�Ԟ�e�.�iNQ��0f��s��Oh�!{���f
�վ�/����2�Ö�E2�٬��v+C ̄�>Y�;C)��/M�MTQe�W������4y�1xa���d8
ڗ:����HW#�3ku ����g(���F��hi`õ|x�\1��\{Kjt ���㥔%���L�d:-x\$R|@Lњ��qؾ�ض	��9��ݎ[
u�ou�i'6>��n,:*a�M�E�7�+�G���\�~_���9\����	~;������*Qv�T��80%���t�2fv�l�Z-wi���/i���CB�B]�� ���]�b(�������,B���'��e"u<D�����Sxq��)�v*�`&��h�
��N��i�`��2W�����ö0�R��_��SWj��C5�Ӷo庡x�
q_�+��#
bcm�9o�en�P��{�`���Z@3���`:��q�n~�V�Q��!2щ� Q1&��	p�y����Vl�+��J��yoN��uإ�n"T��g������S�,�C����̸c�>{����(�,�T�-�F���!��3z��7�7��ͣ+t��xRIB�`��WE�T�ڧxcw|��b�r�G@J��rK��,�fܰ�9��P�B�,.��g&ZQk��c^h��U�� ��# ��G8�,;Hd��t�Ι2���:_�/aÕ�~Q��i[�H�+.�HJ[����h2]��gc7yRFp6�2��vV{�>�ݭ1.TU�A��9�������}VC�my��KWҌ�_O ��c�!3|PP��Y�u��.@�@[�
�US��>�ڀ��B���R�˺�]g\/�i���FV�mo^/�-<�<�k�2���J�$,�;&����4FB*\�0���ɒ���e(��W���\wa�E��gL���<i��`Ǝ��K�n�^�e��͜=Hͩ����r�T�"R��K(KZ�^S��.���M����7o�7�CǘB��֝F@Y����x_��m.߳��뺧l�C��F���:LX�~�~m`\��K���� �r�u�Kr�mㄘ~h��H-o�6���Į��Uf
3�Ú��N3��.�N�)b�z��4KƗ�{Q�.*�=A���0��GQ�Ă��ٛ���A��'��_�>r���/MF}7#�bs��C,y�uy���&�/�F7���|�v��w�_� �r���͡Elw�'���$��q�"�[� ���@��I$,%k�:l���>��g�^ ڥ���Պ[ ����*�!�(l�^#���g�z���r!���d8�ޤ������X|�x�(<�6 !�7{co֟> O,���܏WY>�a���e&&1[�{����*%ό2D��	��Z��I7;FRO�&��f �������$&�UP�%.����4�NCCgƸM����w5�ǅ늠iN�����@�$��8��u\4_*�T�m�ңD��k�;
ւ�n�L�/朒vի���h3d2�*����Nmѵ
�'d2G�'�������NB��9j^G�vb�3Bq�����P���ҎI`XyoOA�/#�E ��/�p4�_z�:q�Cʄ�~�	`�%|$2S��y��󗠰:[,njA�6[S����ټ��A����&ce��08�	V��T�����2η��D��O-D?eu2H��}2�%��G$�B��R��b£�s����{� 2��-P��-��T'�3	"� ��;���vU���I�cdwax��㷵��6���m��*<F�oC�1�m�	��?��5a��]}��"�O)�O���Gc���F�b: j�`��`<��Lb�����|ʶl&�oÞcO5�/f���z^�RKz=^Y��p4��`���8/Ǚ*��X���ޙC6R�z���9�,MZNE�D|�����rP;��:Ry�/���1twɏ�8ި��9�j��|U�jRA؈coI�`@s!oN��bⵆ�@lʞ� »�HW-�!�2�L/Pk�+�L�6�N��v�}L	q_5�0�ϟ�;j�/�?�5��"M���=�0X\��a�y�;��E5Iӂc^�1�C�촗��t�CL5Aȟ�X]�}�wQz���8�G{�ͧ�@K�����n��sp(·�Sn���	R~�tJwac��Q�*U�T��/T�)c*v�{�ɭ����a��2M�+��w�4�A�ZK �ѳx_06'�m>g��ż�u�6�Q� '�6�o�bC���a�z����k�1�5����E���)?����6M.�+�Fp`�|�p���� '�,<X^7s�y���Ⴟ�=k�� �t�!���i����ܒ�߿~̝N�m�T�Ʒ�'��>����:@�yz3]ɒ%��E>{�Ff���?_���s�%��H��VR�]q���rcF�Ý����l|�G�!�d�N~_����?0�{E�(#�R�����F��k���qByu�_kN8�p؃<*ƛ�1w�|1��`�����p���$}�	��D�����>��e(��Q�zf��0��#���0�P H-��mi#r!��r��q����$]�nhxO羖>���hn,�Tf�(^%��lC��ʉ��S���T�_��EL|K5.�^�c�)����Cܞ����^��徾Y�m��W�ޫQ�N����V�_�����D^F��b��x��B�p#�.}��2E��	e�H�M�j�J2C��Q�Fo�2Qrי��'���>Jl���#A��F�2na$�-�Y�r�qu$"].|9���Q��&��#n�@�fL��d�@����U,�	�"o���5�b�rͲh`Ȑ�Ħ�PN�wAG�M}�֢߽��¶�	��q�"�a%���g�:<�� ��Op̭ܰ5��<�Ow-�I!���P4r (���4����*�_t�Y�W�w�B+�g�+b+�sޟ&E�����&m��؃���	���	>���1ol @��}�SV�Ď��vGl����Kj6�|sc�49�����L���-'�@�X�-�ײ�@T�j��k���A�����3�P<�BBΣG���󰧏m����%��k��Vx�cw���(v:���[v�~l ܖH�B.��lg=��镖��˳����*F���·������J�	�����@��K�=��lls��_��bfF׵|Rw��m"���
��Kv8%�GV!.Q����y�E�B����W�:gT��8�L�,�0ɀB�9M'_h�_s�geC�`�K ��]n�f<�}{�fJ�|I)1�v�W��S�Q�w)�ie\5�v���Цb[��a��Z���<i���ʮm�k�Df@�\XK�v����<B�y�{
����������Y§���}+X4�)�QƠ����b�1�ϸ��[�F�W\#���!��,�8ͅ��j�u��