��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���_���W=1����o �6!�z�O�]E�ŕf+��З�۫�y��Z���q?�M�!�(�lYI�HI�䋽�j��x�T-�ѵf���c���98�N����yɁ����.L�W�Qg�ɥ���%�bdy%�ҲFf���r�� ���K焆�ң9�LR���_:���K�v��q�h[�d$���oP�RGUs���Ҝ���	� և�*U�.@�v��9�K�t��	i$` �sǿș��&����V�W����C@����d�Ӭ�n
w.�<�5=5�/�"<�74�񸳾�D�bm�Lz��b����@�����j�L���z�����ʭ�c��6PJd`�b*U5�1�[���[����>�9��kb�)���쟢��Y������I�y������]�D���������K�oL<����ʽ�g���F�@�7 �%��\���g�a/k�#��Xx��,<C��Y�jg��P6��P���,����5����Mhk~�����|��4,�)�,�����3Y�Y������,L�R�N��ÞEƉ<�%P?6�{�G���BTp��c����_��}9��*;������6��ݡ"��uy�l�g��O|d�)qx|����.O�:Е����?6�p�I��)
�~�<Q�w�R)��0��-�p>�y���c��w���Rxp��[璉��]��������ә��Ƣ�iȳ�I��(�EZ����º�f�t<�I�\�T��^LMM�|���6�k�����m�GP�x�5�!Xx����joj����ǘ�v�R����9X�3��-Ks��J���)��U�q�����	��N
*��}�'��m�UUlĖ+�g��B����)l��O�nS��\c���x*p�`o�G���Up��9ΰ��jj��S'=F1V~'ś��3Z�Il��s�2U�a�h�w�_B.�w}���@
W�ؙ}={k�����Q��tM��W6�0��:�))�g�pJ�Jt�R���1��^"�����6����٭=6ޏF �3�;Y�O���K���0��w���q,
Sn:Cj7W{�x�(*U/�ǆ^����F�iR&0U��hDf)��#�x��}6�[o3���N#���<ikY�Z�C�������ؒ��ݞ�!���K+��$����D���W4 �4p�v@-IkrV�U���p���
?��o5�xT��c��kh�<2��9/2����]���u��&�z�+�Q�^���-���e�;��h��'�e�+r�K]���Q	�y3S��b�^I��h�������{���Ѯ�4>Hэ���S���|Zއ�:�zJl���׹z���8�VY��&��/�bM�K;�WYpn2C�J��_�˃������rX�}��3��c����?�:�'�:H&�
	ď;���%��e�(�i7��D���NM�a}����������.22���_"
�ҫ� �Y+S?�g*��
{��W��;[ݜlY��,Lc�����B��w''��︕h���`�E��]pۏE"7%����zO���jM�e��`��!g�Z��a���/�6*zk���G�����e�Ÿ��e�⢀�7qV����M`��<�$�9�ͅf�ljF���CD���Rt��̓4���6�ˊ�5x����7�SD�ݓ�Q�{������C�++��54�:�N�1����?hN�m���5T}��HQT��
��ы�l�x�\R^���S�7��z�R�6@�&X���ڍ�7���o~3�N��E �'TS:�(vc�Z[�ȹ};`���$鏧�'ܾ�m�-���>�(�������s!?��
��r�[��	�ڬe(����Vwv��ڦ��r�A��+���#�.뢽��ꂇ��,��i9\�Ϲ��Gy��D��x5D�e5��<���	�u�n4'���Z���Iyy'y����rdO��� 5��{�`X����)��}��i<�&�����`�h�
��|9A�Rڗ�l����??g�#e�w�A�Z�ܤ��73rq�g�����:�DF�j?��l�&𷆘���I0�B�1�ya�~`w+��.�uD	�+���'5��m�+�A@�s�mn�
���k�h���r~�G|Ȯ�:�/��E���v��S�*�%v8�y�#o9�˱�o�|�j8�e�mʖS_���K�N��{+�@,b�mO��]�(N�t��E�ʻ�?��A�)Ba����E�����I�~-a%�?/E�
�
�2���)Uj����2!�f��n����Z��p�)򀒭�>+��&�����~�@K���#�z�Y6a	��AaC�ggn$7���;��ήn��;�V3��:Pxm��wn��G�TC�W9��Ra�H���躦��&-�,�r!Z5�AW�L�`�꺒_3~�~�B� A����j�8+~��]��sTV�}�n���	m����-��۪��݄¼��X�MU[�QV%��X}D�[�m�N,Ljz�ΗΌ�Q��$d��w�mqǸT+�>����xL��`͢�h��]EoM	�z4�˯ɔ*�^2kQ뙬�q�~Jҥ(�M� 5:p������v=JoO� ��acaC�{7��Z3HD]��
,U��'�03���{�߈{�#R1M��Cia�8������|��HU�bC�&�ڤ���n�O��#�₽ �i'�� :��v�+L���9?�m�~�A��ެdA�"etٻQ.NHQ�(��nsȚ����Q�I.X��I8�Y���t�C���`!{����Z�Hӕ\�5O�d�1wN}��E}}�{��]���4@��B��3+��h���{�V�?|�Pt<s�q$u`�5F>Ξ��c�� ���@]���n�z��B�!���en�:ÇK%�����[,������K�-j����m�'�HO�TO!��<�%�L�B},���y9��Ji#�(| �YZK�)�d%�AD���t�#X�	%Y��Tw�\Q�%/̅ .<�?��M!�/9������Kz1�`�������[[k�+{Z�u�mP5�o^���>�~�UN�|+�3nb'�ary����m����<:,S��)�:|��i�������kNE��נ�l�z�>���B�Џ�v�@�r�^�9ʠ�<�#�cF8(O�]�@r����e1*�a7�d v�q�(	�������O�`/�\S$ň�%s��B4n��;~wJ2��h >ʟB]\GVL��=R�T��)��ZA��I���X���Otf'�
��[(/-y��@M�M{�o��l��]�wzl��apY��B .�Lԙ�*�]�Y*�Bw�*���b{��E6�s:l��>C����}À�����Fxr����:;6j��<m�b�7�Ί�������:~N:X�ݾ��M�N�LP�'���E����څ{�گu�"�����=*�
;��0���tЦ&�1��}W_�g|����	ޘnm����P@���{�`�@�:�7��8a
H`��0���+'��UB#m�{��ͮ@@ׇ���ęE��)6�����Q�=�b��~������|W��5�T�����>���E���ED7]�}P��7�L�=2���ݒxF��n>E٫��.W�t��7$W�~����moj����4�;c2��B����yf��U�n�\ې����nރjk��澋��IB�8P��� ���_��Q��YM,����_f�Φ�խ�y���؇��D�N_��Q��)�Зx`�x����~#��k�`�18�<���'O ��>�l�'CCg������F��+��t���~xSWW�e�jB��\�$I�5����a@�!�����[oQV\�������$[C*�9G�ٌE*Fw������xf�97��S����n���|�}хFO+�G���V���B��p�>y��N]v����w)�<r`��[��[��e溜��)ΫQ����Q��b�ֽ�v�vy9$�4��3k3�	�j�3� �����#�:I��'ߘ���F�����hQ����-6N5����c#r��7[�ԑ�]G�Z'���J�D�=[\H�U|��kp͆�8�n�D�7Ò9g@�_�5��U=�(8s´��T��hR���[&��|S���&����G֧�;�	�
������mqg��ٿMɃCc���b�Ro�[��s [��1����:��@u�d�SW����k�ǳί�	�����*��6�Qi=�>� �ue2H�]�����f)3Q�J�z�3/���8k/-ݖ.H�C F�]�ԨtO���8G�����o������u�ox����{4�X�,�W�7�{���H:+|ط؞����uOq����x�5~ȼ�l�m�BF��2�޵���d��w۸1�� �&k�q	;y�e�N`�*^��H����!�C�ov��f{3�F[�w���1��;�	A�Hn�%u�ᔵ��Qg����#�����Ѿ'N��eR4n1#GTO`�ZU�H�	hQ׼�r��TT5�hm&"G�*��w��`ٶ��Fa#��Б�t��L�wԇ��H`G�_cEP�*�X�il����b.Z�L���@�7n�!?�[��|ߠ�;�%��b��w�	��|�طľN{���3�J���A�nA�����q�Ѽ"�FH���hw����/+������ٲ$D�CJ�vh�����E�^ָ���H�]XJY�C��K��t�9lu����悹��l�ܬ�z�4��@(8��JĪ��Ry�ae�zdv%M���]���^��G>��=^u����ڕ�R�OQ��J�ҋ\0D��M���T�/���7���8]����������K�7_�����=}���l��{`*�i�pv��fcs�^?o@�^=��m�<S��������Y�]c�\P}�e��#C��R� �G�?���u<�Z�=�u{��Hۛ9�C}BA5y� '�����鵾6ĠY���q�-���<����4�J܎�r�KA�,�@Q��w	��w��z�Gv���l	��E�b��5술c��@DÁ�"<Ol������Drj��4
�5�B��e��?Q-C��������ن*Ҡ�9ᾞ���$���۞��&(�̥���Fn�pH#��M�O��'��s��,���Ay�5XC�=ܿ$/m��2t��X���4�^�|�NZfm�wWZ^�p<���H�g�i�"��R�VB��h�U�9� }��rlx��6ߵU��<���N3���X��K��^Ov�!:VXxiL��d7 �C�0I�s���G(���52���o�`	��GP��*�Cd�<�nuN�<��y��v�L�X�D��}� ��F����+O"r����_F��^7�r��f	CϠ{"l�.�{�����yYu�6�C_��+��6/��y�}^8V,/�p,8Xү��B�m������84�)z�;`��-�u�A|��0f޹��p�
$DD�>�!K��{>����=�|dB>� &xTdUfF;��.`!�%37R�
�35:���DX�yv��:�����ݻh�m5ȃf�G/�	V�:^�I�� �*�{kb����#����/��.���ܯ��.�0�l�4��U�Lz�iqJ��a��j�M�d#d����5�,|y�#��SwGKl�A#���Lo�4�I?�C��?%ݑ]sˏqҠ�l.� ��*�s�����kv�H�pEb�*e��Y�_��u�p�Nꙉ�7{�&iɷ�a�����������%��b��O5Il	 ��,N�1_.�;�^{�eN<�����Zz�K`��刦�<���2�̢TJR��5���l�T>��z˥�HGi��Y��<v�r�ԟ� �TT�uQ&A�|�ԡ 9{V��x��`k��[�h�4"lb��5=&JbUo����`@LV���!Bh�F�_�zl	㛌��i+�d����������n�
G�(��8���Q���֛%B��ڑ[��E[�T������	�Z���`?���v�[��9�폛qQ"�����Y��vy^��xF�Ah�KY�jʺ^���W!��6[]t������ʝ���o����W���'q��!��δ:�֬�'��k�~ϕ�[1FM��I�Ț�rz�K"��`���zN_]�9�r��JN�	H���ZH9�:�fCj"�ju��o�g���WS�FZ��E=�a��G&`-�'1�5��lC���T�	�"�'���<�t�@�	��Hej_jRMQL���K�8h��x��N{<3�mzO>�Z� x���|�#��M�BW.^��p�y�G5�t+���Aܫ=2ٲ���}��jv%b(�Ъ��H�@��g�xȗF��Y�
�YS� W�/���i�ٜde������M.�����;�{oj�$9`CW�1�3/�>� ���#���J�<&~+���T�m�����	1U	�`Ϳ0����G'�Quܫ����窔�P'ϻ���S��:�v1���X�^�A�v�-�Ba]�'w男�M( D���0=��Y,��YJ ���O/�P�u�kMy��J�O �
z�8R�pîa]��<c��Aڪ�y\�0�t�����a�(��0����s��0�!�D�"1`��{�Q;5S�D��
��T֤�$;&�_���K ��
Ĉ�"�s>�(^�j�Mz3v�	hA$��
�I��5b+k"Ǆ�+r�Ќ=:�k��qvg�L0���0yO�V؁�r6}�4?��T��`ױ�5�g��,�S;��ׯ΄���hb-|��S���ඖepO���]+ym��7�v֗�9|�B��Xiؖ11
��j���_����Uu��}ɾi�F� �����qRjR�`K�%k�L���D�|����IU��C1����\?oi,���[�?�	m�/�م���]5ʫ/ �I���V4��D5�����6������&!�������_
��ƿ|�2��ٳ	gL��$n�"�{�:|N��h9���{BCb ""�l��h:��hm;�b#9DK I�R���rJ �53�?I�eѺJO	,�IY������;�#��A��N�"��Mz:�<��s�U|���bi�k+W'Lq��<��� ҙaY��y{��x0E;����z���c�.j�ͫ�ŒQ�i�=F�ɍ��#a��0�����!X��C�p��G�Jk< �Ȩ���NBI��>���}�j�!#��������������BM���t1t��"�-�*dG<�u��.*�	�-��:N� �[�B��Dk�):T-�@���lR.��@Q��]+�g�_"�Ƌ���us٢�zB�w�4���ʖ��^Lհ���7��R ";�,�#IAv/���O;]٭˩��]��j��C%�J6|�Tzm����"y�Y��k;�_���mj(a�.���?�$�5��I�~�k�
ce�������$9��ԃ��D��>p,+���H�:��n\�A�8�*��U��̍.��,6�j���R�<^ݲHƅ�-Ӗ��
}����J��D��hYF�ݥ�a��u�b�dD��ma2K²Fhl(��-l�?������r�h�QԽ�`:���\/��v5����M�}3�v �.�?,pͰ0n"<�@嵲��yR���A�{�")�õ��Y���ҼÇ��2���Ӿ)�_��'�00U�<�����M �{��|E�������oE�]P��^Ql�ǵ����I69
C ��^L����9�f�$��טox�*VC�߀��k�I�
S���&XX����S�ث#�xF�(D �q�K��S�� n�q%%AϒQ!u�Vk�S��=�w|�
&�<�d��~Jb�@���b�-��I�b�}r̹������q�~���� a��䅱J�-�]/ށ�❸��d�T���`��L|?��v�R�Ρו���e8XFW�����{{���/@��A����+YyK��m�i~�aR!Tv"��.��4I�o���{��f��&�HzLz���I��c�l"�LK&�V26SeRq9@�CvѼ�D�(d��%��-�bѿ�W�Z�z��m��r Z���\ӋX�祕�5t��G(?�-���J�{w� ���7��C(o�v%�b���',$GQ�_8βM'EhNILa\*��|K6��נɗBrJ(`�mէ�CY
{z���>*&-�HTŻ��� n�7�~�=&�~
��N�r��5Πkj�����_��(hk�w�/���,�f
QdD�14ym�H��hjkd��gvQ&>�\���J���C3��@D�j5%�|JY���{F)�s��Z��t�1�(FaRa!��p-֬ (/��o��E[��m�T��+��Kw|C>��2co�(�|�n�i
b<=Zh�� nG�����[�#����;r;�d,ހ�^ɐ�+���}�[������ۯ���D��#���!8�^Ee�����99��� W\�W�'L1M��91��q�n܉���;��;�I�N���!4[��!�\U$�50RK��eM�����D�Լ�mFR�g*Ι��% C\4<�����3qǄ��S��YjƢ�7����
�Ȇ"7���T��s�^����>gAȒ��&�"�R�z��3�(�8b2���3�р���Pt����[)R�-
�5"c>Rd1J��H�y@�yZ[+����c_A���/�+�E~�'h�*[��}<�G:#�����������3��.U�x�x4�)�x�<�.��{��l����)^2�'䓛)c׶������������X��џ�|l�^�i����_�v@���n��{��8�tx��p���(�,�����	9&��+\B�5Q��]ܢ��z�Gx�tS�0k��J���}
᝟v�q���>)�����t�Nv��;�_�D����@V��V�F�q'�D�R8/�ɢ�K�n�F���x�/ơ]a{D�w%���ޘ�O�y߰=�-��ȷh�+�=�=u�kڰ]Xp^̂�v6�7�x����˿ʪ�A�_	�]���l�RO�2��6�$`]}�&(
� U5�$(;��+�C)���Ҁ� ^�Rq ,��HE�[����L\�[EL����Ȏ�D
ak��>Q�P^��~T5��[�>������;J�����*�@�B�V��`�Q����R=�� ��;��BQRj �]����'�w���Uw���:8�����m��~I��8��jud1�J�A�;����\&Gjԑ�h���ԈVIC������
�Ka ֒&����;F
9$9�l��!����<Md��2Il>�5��J��-���\|��nJ�d=�;�#�A�B����qK�z'�Z���d�	]�y夒qF��U>�ʹ@���a� �~&�^L�9�[ף[��2ht�9���eG>�dMع_2��"<�8|X��ss�BY$Ң�j��Vݔ-��<���Z������%<�gt5��ݭW��~)�l�(�=�+Up���~�-NY$mz�%���N�k ��gE������	*IOt�8��S��ڀ��C&�jt���f�z�Il��(�Grw�_���<$"˾��hc/T-z՜�'�޿�r�?9���T���>��1��KE���*z�aI�!��R��7w�n��N̠V%��j�Ǝ5�����[�6���ǟ��=j�&�����E�5�"ǯ�Z��րNE�������&�ٳ/*}��=' �w���W?��X�J��׭�8H�3x��:+L�M����gו�,攟�^z����Eڦ������9يאAU=��5�C>I��o�e�U]�)�ߩ�����U[+����!������>�~P����JӒ�>L�	�/��.��:��~���<vGR��e*�<lB$w6u۫(s���y�A�+/n0U�ָ(�ޢ0P�K�l�q��CGB�07��S$kt`�.
6�f���'�q	��Ҝ����9T�%�~�)kv�-Zu�u�}�TI�n�aQ��n!vk�N����̆� dOK���~H������_�&��imP��n�O91����ƈ��}u�bĽK�0�D�#�GV\շx[�К���0*ɏD�IY�q�6|Q�V %UA��[KN��=�('�Ƽ�bVp�2껜���R��`Fv�^�nVn��>�~�
��@��=�M�M��<��I.���Ҕ͈����6d*K�9� nv���f�Lg��Q.XL��ӟ���f��{��N��2���OMi��,m����u��IVh��8RMB�A���[�$��4�yA��<�����pu����fԜ�=.���u��a�ٺ�f���*j10�M^z|�a�D;�Ga})a�����m�:.ZI�_�;T�_��<?�����s��6�	���71xd.�nR����\��Zળ/��зL����v��Ы|�~�Q�`���15F7L�U.��,R�-�r�