��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbI��2��Ձ_N�RL��������lx�^6Y6^J�zY�a�`P�v*�^ԑ�t���e�!�x���I���������k+~8C�S��'x_8=�~���#�GT��� E�C:�H���c�a�@��?��!JxE�ǘ]o��5SB���ո�C
d	�'1h������b����9�{�r��K�t�1�N��3��e��L H;cb�C�q����/ز#Ԍ�9"c38mt�������ix˓�u�ճ?_Q�􋹨QY�K�G�n�р���i%���9������Ҍm 9�w$��
��[��Bv��D�f��W�*�8*�Q괽�8������1 N��Ecx����U)�ci�ܥLl���1䄛�M���$E��F7"dj%7IJ�B��V��-��č�N��D�J?�.�!�0x�T�����f���| z���Dv���]�$J䙪�ڛ�o��c��,��=+O~��0*�^��)�����_��a���_M�������V������cF���2~���h�Lr��e�s��n[
�{q��١6;8�w�=�qǴ�1��ځYggt�Jy���X\Lܶ8T
?��xf���ʲ�H
�x�fʮ�b����v(c�iE��� Z����<=[oԹl!�QͅIt+���{�p�H�Tk��@kw��[w�c�A6�;%9qF�"#� mB>�)
��ŮV��Y~�j�P%�$l�\����t;k6����Қ�+�]/-U��ߙ4�Q�L��±@���Li���)����D�OWZw��n��k-�i�(ԅQ��,�����]%s��-hD�t@�&i1py��_m�ĜK4 h��1���+��<3��ᛉ�m#��3I?���b�b�
�$ �U�e�N�m�T���Y�J�a�R�1�+EΌՒ��.V�=�Js�仭ڜۍ�{jD_��W,�oJ&�W��G9�|��5�!�3��?sc�2EE!S��'Y۪��@/����f�! �U �^k����?@ل�s�/��!�hI��Nl��J�����2�;���!��39�1�&�����u4+>�+L8�s|�M��ڱ%�x�[�v���1/�G�� �h;�)c��+�����y/*��мW�e��X��y�����q��1@BIv��^8�����p%��E��ti��7�G��C����Q8W��*eZ��ˊ��8�1���4	<k^���n��#�?/$L�a�q���|I�M�=�&@���Ʀl�9
!3��~��E�O��t��*���q�i��|��f2'2�&�~KH��⧇�?������V�&s���rBL�x�S��9�5��gg�3�L���@BG9U��m��`St&Mna�F���R;���2g)L�-������8��p�l�d�Zg)P��I�B�}5p��w661����-����ǜC�~��O�>H��h�X3tZsȵ��' ��ww���M��>�x�?�~VE2a(��z�{G�䏞K��`~�3:�+����Q����'G�V>�ɜ�|�(��W�'Ќ.۝�_�9��<�@�E�`�x�Ew�ؿQ�6�X���Y����3�b�;[,D��=i��2��7rh�L8_�֌2Q3N��5��`X=mmXz�j�Ww�+;�=/�&�k�Gr�i��-5Eܴ 5K�[�9}�t��lhF�(�b��'��Z{���36a�N�`c�s�h��֤e�[�?�А���q���}����F�y	ã8��Л�EJc9�q7��<�p�w��}X�\��j��VS!��Z"���]��YO��p�g
�5�/����#W��T]�WhO�:a���q�����R�S���$��40ϔ�����3�)钔^Hd�ޭ�G	qmO��������%�9{G(RE��'8;��)ֈ���cV�oG�׭�%�x�_��8&|l#�:v?J���('c�aB5�)<��V�uIe�!���ܿ�ƈ��AD�P��ͭ��f����Էy���~�EAuR�S��1�6�N�"񦸳pBP��~����NE�$(�`���,�N	YӒ��/�Qe��O��ܭ{�1�>BJ�͢l�?^�K���+�a>|xQND�q����DS­����rY�[�[^̸��p����M���GT�}�^���Y�����3FR���n���%N��~��gN��:����	$W�����[�7y����-*k��-s�7�;���:̨h?���U��nT\\��<���~l`.��Iq����i