��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2)��Tق[�	��5�Fy�
������~�}�Y����%�$Z����!�:�O���<�K�G�PVP"�H��TV��W��e��x��Da�	�����V�BK�*��s"C[v%�����Y�����N�ϑ�m2(ѲQ�q��kY\�籾q8_�IagSPvY�a�έ��7�IR�N�50�[�U��+�Uݥ]&�K�ٻگ��`�9/�Fp�cl��{,�?�ILʮ�B]��j�Ը��+��EFN�G��T��\��h�r�C�b��|�p�4r?�P_W���NY��Nm��K����_����5��i�I^���sC��y�&��Kڭ2�0�����}R$��X�NWF%�"fuD]��FJ�I�"K\��~�.B�f<���<���c�D�9�Q�Y	7J����͙��Z��uRX� M��94��sŤ�egE�x��_���C�OYu�)���ST</�@gTٲ^�a�w^	��1��{"�H�5��q�V�r�W�~&�>(��_W2\^?p��<)��RG��LsL8���XH��wr8K��2�JJ�Y�OE����f�t�ek�\�h.����'���Ȯ�1MAU�wGV�%td���2�Ӿ���.��n���	��?�ә'�M˪�G�aJ��"�� g]'�	�2����J�Ǭ�-��+Kwͅ]_'.)T'��~�8`��gs���&쌇��6!D���]i>Ow��?���Ba@�KPk[��ԋ�6��{xB��O��$�W#�ʨ�T�f_���x�3Y]�ޟ�a���/�^�6�rhn0C�^�h��_��J��F�4�'R�{�Y�h��KCc=`7��c��a��$���A�J�k�b�kL�$S��>����X���(��	��u2�q�?��l��~A->�v�AS�{1��o� BE���ak{+�U�\Vx��Xm�J{�B�yt�
��bO�=�١r���<���,Ȩ�8ڵa��j�w+�alz���Ze���r,���a�0?��X1k�T����O�Q���e��& W���vx]l��C���� 䘀HF:̞k{��灗}��)N�����c��SAj��&�Q��p��oN�P%Oz�V����Ym�8d�ۙ��#�!�X&s�g�t��y��׌�CV�Yu�̘`�G���G��3X��!���������~������b� ����⎮�6�� ����@�Ȯ��	>�,0	�}V�o��@��Pl�:�9?:��`c]��=!>!E�D��:���|o<���~�9���,��~U��I�ė��$2��I'kl��H��,"�T��-��d�f��I���Y������M�9�f[�U����kA�D�����I��㮦���KP���ܫ`����P�P���vb=�rr��L������
q)flM�S�w4a<�J�
�ѱ�ɂo�Bցޢ��I����u2��ތƚ�r�j�òU���p�YL3��Ѣ��93W�Y��eS��mx�1LgX쀍|�s��H0�sǘ\N����)2q����d2w}Q����'�ɖ�F�H���T�BPe�mU�dt��P J���f�mz��VyN��b��^�<ˉR�r�u8P�����cq?�T�� 8��F��m­D�6�K�\��5��?H���u�EKF�w֙���ԁ��'C�Xl��ƞ����-U����d��O��ޥk9C����55BwA.�e��q�U+���hS����sH�|��C��W��%Zpꔗe�Ū�������[�q��l$�QoHR�3|��E�Ʉ�v��qq��NU�}�#�42��i�mp��U*�Y�N��tx�8<��&�a�͠�m���/��9-�T���/)�L��� �f�~V�s��tb����dHC`�3��}%r�Ѱ{lAWx>
I���!$�G
'�u\��C���I�r�Z�P�h����F��:;�b�,h�A��־�Z4���h�zL���{U��|Kvl�Ӱ�.��O!�+^�O-#�r�})ݷ���6����Uq:�H��T����f��>l���r��Iv�����]�ϩ^���^߯�R�CjK��9�\1�>M�ϛ	O�iX����$��F�#�7R���>���W���pQ�(2Ԟ��&<ŭ�U��1����Z#w��Ȇ�,0� �LqD�����e�����t�C˭n�ӮV9o����A����Z��b�N;��^��V����QQ$��oH&�HLE0�T{���þ5g)�!'�F��1S��1��3�ɄO�O�U7��,k�j���w�=�=ߥVgBI�2��K�@�K���7�1A�(w�e�/<�:�={lQ�%��	*쓂
8�'��4;�J�	�EUL����OhFa�����7���\�Lk�ˉ�˥�q3`��e�1���
��Ԣ�I
�c���&�J07]6O	>*�*�X���S�>�v+�Y3z� y�JDO����FZ�"���ګ4}H����<V	��"Ծ�+��5��L����"�Uanh�R0<xrv��^5������{�-Pe�.3�+�u�Ys_g{�u�?q:Ry9|�W�\�/���� �׶�-%^EX���Gߓ�4��}]Dq�%�2��e�D�<h��'�G./�»֕���A���[��P�^��7���d��k�����G�HU%M�? ��=7�|�<t�����Tjv������C%���>8�ј�^̕���}M/��
|YU+�-9���A���^i�/��> �C#=?����k@��6!_�]�0Tvw���rY+�b����;�e���8T-��:<u1`��אY��ǯp�w*"ג-`SRD����Ͼ�9�9��:���5��[q[�X.�N�w6��pݐ�+B!"�R�����q@�b���L��U��GT�a�</|�����l`s�;��C��y�p�\v��,͒�s�ˣ��pn��2Y�z�p������	�ĦD����a�����5�Ș�` ǁ7߄��&�j��åY�-rHK�as��͕C��.t��4�$��@W
H�����%D���S�'���8;8U?��g��hVU-Cg�*���!9�3߇��~��B��ۇ�:��JyI���E���'Yx*
�"�
#y��6�a��)��D�Ǝ�V�n�L��ί�z��18Na�/ԅ��AF�CG�m]�������1#�.��b��Ω���G���X:C�WZiP�������B��V&�I��	�E�e��3��r�3�������;14DJ�B�#�r����I�\/����Rr9�؟�2��t}}F��L(�-9���}*�;�I��k�*6�G������T���{\i�pu��N-�b��!l"��jK�%�Ĺ��xB-B�e�\�3S����If,�vt�-4wH�����d����=���XvI�fn��&�x��x���!��$��G�k�K5~��!owǴ�߳pjuZ*�
H���7T ��z�pg�~��-�>�_�jRu_�@�P���Z���ȓ=f /�m	|��K�����Eà��ev¶���#����Q�Ma:L2��I�JplLP�Ű$�'�U�|^r�P����ěcqƪB��b,y�j�x��Q䰂j$J�T}ͨЗG�:P�u�K�!���0�e�u��bW.�k�Q�L�����|AJ_��O�9v�R{�W���ʒ�]�~S�vQ�kt�Þu��u���B���ܼQ���S�UF��b�u�3,�%y������e���=����Q�߶K�6�_�w;L��Q	��]\�l4a�d5�ʹoH�\!(^qQ�7A��IYܘ�9dL'��A+�:�幪(�k;�ƑD�ҹ�z��4�_5܏ r�O���}�F�/?{8測>0�����������̓�Cv��a�nTV�|�!�y��-�ʍ��;L�Q�(�`RZ�I������x"���V�[�^Mi7����1%"���S�]{f��rp��#&Z��.'!:����r�^���؛��h(���rm`���>�=أ�(�lA//_钡�d�D�޿tF��Roa�=���7ˑ�?���{�7Ƭ�;�y=�$#
-��QL�y?�z�*Gɦ�����=Ӧ�q�!�	Fj��Ă9�Q-�(�v}I�$Se�h���:��'����~;o��d��J��H�u�T
�,��~�8���V�A(�*����P���!��p= ��u~3��e�:A�5�
p
)��c�ކ8,�cn
�9W��Ei>)�p�g���������B.B�-Jۡg�:���)�K����|F�yjlaN+�֐������ߒ����﩯�EnbS,�֪����g�� )�o�5>0*>N�f�>���e�jh�v�������;��.�l����U~?���{.�E�yP�ˊ�z�O��j��|�J����TJ NkZQbp�4�v��!f1�p����k|z꤆*�'��� ʆ�̝����(ޣ��� `gރ$�-��y��	@��$-�^�y�2�=���<Knտ��_���"�!	�ק�,�E��I��Mn�i��q�%�[ƽ
���u7�,i"���"1+�!h�m)]�Hgվ��`�}�:+��-m�u�	�,�0#�ۛ�wڄ��3徱t�6����)��B ����P�����qjNЍ�����G%C�� �y��f	�XE�%"c�**gc+;!�n���<y��±�Z�i#U�0`��.�v�ӊ�5�w�;�u�+g�\�W���@2�����z������EW���$�}C~��Q��|`��өh
�,,8(�~��=�n�H���gʀ��R
z��k�V����Dw�` ���t"!�U�#Q��w��Z�}�"����o��8''�!7�(і����9����.���~P#g�}�E���ˤ��2��lͽ�w�&: FJ�q&N�'{�R���EI�k\�İ�kձ�"����Ő�7�*J�%���A��U�.����p-Q��e�qe_Y�I� �c��˚:S�f@��D�;ᦵ">���Y#�<p�̱���uG���֐��C*�쩈c;G�����E�O0�ĝ!���@5$�ef�*��f�~��	��>\��@����s ��|.5C�=�_����d��7ڐ_eԀz �I�۔��f�
u�v�vE�� *�V*�׳q�1R��O���D'-�j�