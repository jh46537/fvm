��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�=���,1�jӛXT�d݂���uL�ퟣ?���6�FZ�;�o�I��ě������ߝ&;��5TAq8ץ�?+ܲ�#W����utF���E��	�[D�N��:�F���K��T�o�����c5i��y<�--qA�~$��,�����}T)����5O{�D!&]��7N	��j�ySe����n~�Cy1Zb:�^��x�,�I��a��k�l�G�z�59uf���穨�Tp��ͤ��m��y6��AA{���E��N���3RK}<�F�{��p����Ď����j �x(��9�B��r�����}���j��P�i�aW�⅝l?���c���N1��P	tfc�E�=&!�#2�&��2~���S��գ¦KI���鋔Q�<�26)�ni;f�"m	�]����ܡ����U��UȤ���"�s.�� �C)�U���������9i\�i*�EƋ�|�YMwl�^�c�ҕ ���N&���	KX�BO1�.̵�ގ���_0���lE��:���)�Zl �-��dE��T���Maж۰�p
�v�p���P�X�b�2:���ݣ�-=}�Ex���x��@���a�D�KRH`iN0�:��mv�wiq���W���_WC�Q] �/�dbu�"���M9��&i�M��z�x3�B���r�`�8|l��?9[��#'�m`�������9�i��'L�6��6���PM��/�\�D��t��3�V��>��z�������cʉo�V�MI�HU������	��JܟZ���Ex+WM�a)�� 4�9�La��Z�۝y�e>!մ���\9r��y�.���]3�=�q�cX<z�r0s�%j�$��~U���Ķ�i��	#3��=͉�"Y��_^��g@`��@���~°¿�k(cB�_'�$5~(�J�0�⛦�l��({Pҕ'���3������yP��?���� �Z�D{F�ߨ�۽N�:Mۤw[=�}���S!������4ǆ�R�1R<埣���u�U1��!t��)��U4�ٺ/KjY�6���cKM te��
�E|Etp���p�ΰABڠӮ���D��3;�7�5����Li���^�!I������\�X4��rD�����e�<8 \9p �(R\(���3a�Zf�������n i}	}�
��|��r�+��g�8ޕ&�hr��G�f6{�g#���R#�2A��Hp	8i�������:��o='�V��Ό\`�}��YAg����V�m�s��̣bW3b� �{z��l���6�ഔ�-�����%B����	����W\Ct�|Sa�:����O�Q����Vs=�MF���A��p�eSdnD֎���WST�BڻfKԀř�Ʋ�1W�F�4�
�@����
\����q�o�c,�]�9HO|0;p�����ԟe�]�!�E�@kr�7�ZG��gJ��cf�ǍRf�U�H������*��mJ�Q��͵���Y!��z�3K�J�gN�� ��G53��Ɉ�ScL�E�]S��I���j��*\�>���0��I��F�˳�K4�Q�E��EWQ+����.|47g���ɆJ�����Z�A.k��p���ڦ�gZ����&x�u�uT�A���NF�ʚU󩋰e2��
�l=��{����i�ŀ���s�����-�Y�x� Mg&y�Igh+�6��y<�9���4?���,>8C�q��G�k��彋���nSG �~�ğB�!QS��d�����$�
ų�D<�����C����SV�M
ɻ���_1t�/߉6?KR��dT۸���π��g����R��2��-(.W%L/:�h�4�b�ʺ��D�Kp#���5S=����W�}~��78������XXCo�'�!���_��S/c��9�����"*^Ÿ��T�/.מ�B��$����!�h�6���b������h8��<v�rb��Ƥ+)I.e�y�H5mr�N=�	�3�rF��k����2@��B��a ��z���e"�,,p�m�����w��|V��S�V�4���Y��0����u���v�\�r#���?o�b�n�Vo���\�&M)H9/m�!PJ���9�]�G�S�av/�矨�I��0�f��.�:	��.�j�yK���x�Z*[x�E	�vU�ָ	Z�0ä��a
��h��r���O�ͳ i fƘ��� ��N�ܙ�$�x��b�\�f8��N4	�*�{﷬��rA���}�{�w��Lx�P�m�Bed��<4�|!F���8i�M��"��*�r�]�,_����ЧWx�?�AK��0�K{��Ls/G��ݹ�����$�6����캁�٭�������KX�Cj�?>��X�x�
�V'�Տ_�Q�[�p}fJnZ���]b\^��c0�zne^)0����"&��D���Z����h��.�urہ!^�V�����6��a��-�+� PJ��h.D�/�í.|H�t��T$�2W|��6��4`~���_ yH�,;l=Dy�蠔��`�Dɴ��;��5����6��x��A�F@��YW�w\,�7��C�:��T���2w������b�H�O���g;H��[JN@v��r�$n�tk�7g�� �I���N����� ܑ��U���D�r��뮚�v-� ��	w�҈�]jo�v+c8�s�x�י�U�TIH(��W�멠��0z|e>����f̐��1�bn���YNJ����HT�͵ґC�\*��X;���2a�|.�L�3�x`��B��@�(�Ú�{dr�#�L� X���)3JW��;o� ;�����y����`ޟC
у�F�KWl�X��HHB�������.����>�Q:�/��ȧ2=���>��D3�]�K�)��*�<�订k,�e�����D���Cם+���x���|y�� t�P���S��!��m4C���:R=�ɹz����)���C�9t�|l}����\߼�Ye�r�U�a4����E��׀³}�� JL�U:~g�؂�%��h�{��ufF�{ő0z#��?h�܌����S=��%��Y�kg
A1���{�_C���ge����(g(L�������<���[7�����K- ����4�)-*�A�ܖ�� �y�F���N�L���w�P�����EE&�Ѵ̻w����Q�t.�=������J-���d�C��%�vYʩ���m('�u����9�3*�}����"�I�Z 5~Cl e��Y+gI���� `��p�{���� ���BՋ���v^���cWF���%��G�x�VuL"�y�3Q�A���L&�+a��wi����*��	���rzj�N�e�ʮ��0s�ߡ�C����^�$HE]5�$�������5~�K+½k�MA�]��&OJ:���[((!D�BF����-~�}�r���3o/W��"�������F�[�z�[g� {��X�4���\T�M��!����l;P�������S���kL@�,t�_)g0f��l%�'O�l�֚^�;P��.�x)��b���)��q~Al�%!?���T�Z,r�ϝJ�M���e^f;��X�-)G>����v5��-��q�Ix�x	�i/"�����D5!21��%����ǌ��O�f��K%�.�uY�k�����h��*4�(;wJiU	���e~ɚT:}�j�7�s���#3����􂥃&�t��w�[�$��o'}Eb!#}�2�|��� ��d�:bh�����yk,�����UP���ٷ�ɸ/��D���"\x��R\  �|� ��٪��e�]`A�#��Yo�mv&
���Ւ�>��o��4�k6��(��ˠ]䌗����o�/�W8��Q#,�C��b�b�-���3[�]��wLXbﱌ�a����Z;bd,�]aG��p����VL��.ͳMLf˘9'�n�|A Ӱ%�ax@}��w)�NK0_��Kp�N����k0��5�[����m���v�ь��]�~=��b#��3��\��|@�X^��
��Zѣ�v33��I��7hl��&ҥT�z�ŷ����%3���M1�Z6E��.�s��9��χBAn;�0��;*���wJ8=IJ.��|���R��/, ���x�S){u�'�cI�c��mA6�����&m���O��C��r\�T�Z�}�䜗'CR�%o��:��d�ۈ������ۧ��V�p�S�M������_<�X~]̸�*�6��%�	N���<; (�l���A��_p�K0A��_�e��1�_���8J�0`�Jٹ�S���[?I���7�"_I�K�Q9^;j�l�-P��u���@�M|��Т�P �]6�#XW�W�	��C��7�����*�S�攬�"�� ��$,+��DJux
j�GN�te��d�j�Uy��|kX����+�d�N[&D����l�C�n\�i*:��vUQK�]���|Ζ��-<�/b+ΞF ��6�F�S�/x����箴�~��`�a��R���k;\�mӨM�z�����O���M��r񜽪����h�DiSM�Us[�8aP�Ef�+sQ�
�ςp��v�Q�<~!M���Q\2qh<�?j�ΓRo��o��t:DՒC}�����0���A�vU}K �N*D��*��%%�9� �"8YP�T��*�
_�3qH� �������T6F��y��ه&G<�;_�~/p�F������ �Q�>�n�5%�hf���Z`� ʰoQEL���u�R��b�#3sH�yy����P�b�y�yX�����ǀ����ӱwqa���S�[G��~���]�TM��߄4�� ��s��p��׸�Q�����]�����<�sR]e�k�R�U�n[���&bu�1�J�lA4/&Ρr��;�{���`���d�F�NaJ������,�Rn\��k���y�(���1@w��KaM`��R��!���[RX��jеH�e��v�֥�⍮~�R�>�^9Y@�H~ZA��
p�e��O+��1���z��)���#霏m�K�-��e@���tC��LP�=_�K��sP�r��u��q�qI[��ݯ�p�&��LH ��K�<Θ\Ax��`���������J���4_j"���!3>G�bSx��i+1����r!⫎�xV�j���ׯ��R�4�Ф�V�E0���@��;�2��ԣ�=G�e��>�
�/����g�$�HKbyfS0k����S�'Đ�����t[�C%Ɲ]��
��Qi�(w&Ur���ڎը��Ȑ�u�<��67Xt��"���� ��.�S�s2[�����5*�vj���^�v@����l3t�yτ||)�Q�X���΍��l�2X�-9လ�$���U�]�