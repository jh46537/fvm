��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*�ũR��KE�q0f�5c���{�싚|p?9�+\.�Y�=aj�h�*�c���k�{�h���"�A����;G�2���e����,jF^+�D"D]'��t�hi�����n��w��LU��C�fZt���	�,/ ~+V��`�X���\X|7jm&�`.5	K�<ש��d�/�;;���=����o�7�m�t�I���M)J!9����F
 �M@ڕ:t[ʾL��-=o"�p��W���g�@X\��qm62�h�/��s�r;eN7N�ݱ���Y:&΅$��T�Y!�v.$J�uyj0m]�h��VT�޴��%)&;;��Rz�����¬��B��rf���N�պ��*��k��~��#M�������l��+*�L���vc��*nإ����l��̓�tA�bg�j��4xW:�XW�+�Â�x�<��86PP�ܓ½$�Kׇ� �{V��_(9�~4�}��5�y�J�T� ��̟��.���&[k�H�es^^D���[��Q*O�1	�(����V��<<SVi]�!'���Oឞ,,�rA��|qs]*�2�ԅ�����������we�[�>��9@h�w{Ne�RA\����s���6:�q.p$��f�����:�z�]=2a0�6��.�09hS� �3�?�b~ɟ�r���F����3���A-�k[?�,hXD��-}m�R�6�҃���n-��l�p<#�����B%"�l�.�&�.��#7����n��B~���|v������-�kG_,�)��y�L/0=�q�;�*���jx���q&F�5��ُ���[�O���J�*^����T�z����=�&A� �}�jIf��T��J���&�&� rcP׺�;[ZD~���t�񹫙���5��d�Je�_C��Y�v0�_�Ok�칬��U��* �1�o�>Y�4]4�RRG�% ��|Խ�X�����ܙ%s�|��ϰ��i�=��  ��ں�KV&����P7�O�Ju,`�'ȍ��-�&��ZRML���U�'6c�E�;��y��ѕ ̱�<��1��ޯ�K_�<k�5=f0�{q��������ڸgX���ba,��o�C�����u�v^zq��$G2��w�<�K����<Ds���&ʹM���]\�^���z�9?(�ѱ�}���]��?|ƃP9���W�|/Τ	x)-�PP�pG턭�`���:��=f%$L����p\�ϼ���$�����/CR)v9Ic�G�D��y��_�w/�u��4+���n�ֺ:�Z���^�l�G.b�pV�au�1&x�����1�őv-�:�`U�8�!����2j{��8����Y��9vz� [$Lht��ֺ��X&3�-Jq� >5�Q(/ ����on�(L��,�UzE��v-��!'�e�³����k�H�ב�v�ވz}D��X����`�p}+�>F�0���^��a��^�2�7e�𼏣b�_,o�(�ѩ0
��S^�%Q�*��� �e��*G��zHY�M�/B?A�2f���z�
�a����5�F ���;�'�����'sf�1g���9;�Ƽ��Yz��0�s�2?4�O�@'J�-��H�"�j���L�Z��_� �$Nn�2��N��.��݋[+IaYU���/_�I��X���ɧa?�e1��S�����%աu6�s2Ruz� �5�i$A��Q
�8w�����������;l���W}�c���Rm��IHp9��Tj�l�S6�q.��շѼ�~�I>L�E熂�A��X������;��<30��;X��AU�s����|ޫf(P��yg%�����Qȥ`*63YYe�z)��3rOV��y���'����JݲR��jR�m��� ڭ b8��O���f���Dg��%Ⱥzz��U��n�i�j��"km�[?�%.��Ҥ|Ǝě�j�����?w�]w���]H��\c��mg�_��0��)����9�K���ī�h:ޠp%�4�m���G�Kv�G�D�W����A�DW���Z���� L�Rܐ�,���3%+�pHoC|�� ���
D^�;�{zΊ:�_��\�[t�p�g¤kz�g��Y�B�w�	Cd�Kxs��9^Na���n�N�9[��������)���0<�ö�1���~����r^�_�&>�w(�xY�����v��%\�@z���4�^�#��.0M��J�%�A
�Q�p������/즹T�B	�T�����NQ���B
��'Ч+������)y�G:�������zO��\\yȢ�]
c�h-�Y��֮1�%5���	{G}A�l�����A�@ܝ�@��l��
�<��h��<�h8`����y̽��%ȗ���g��fEO�g;�2��P6�!C޹m��喯��ѕ���f�����x�^	�	���K���4��8������9��\�v\#R IX���_����BЂґ���߷�>����k<�OE+�=�Y*8,Gc���A;����	| �g�G{>#�pԽD��2R��J[r�=^q�N��[G����_�YH�@���U,w@Ka9Ia@��������D-AQ�~����~��-�Ū�>匴z(�K��k����tҶw�\uT7Zw�E�c�篬��ӄ��J�>�XF�5.�q�.B��A��GZ ��w_8���π�b]�N��aVc�ݙ_��������R�!�JS�C�=�תc<���U����G��l"�u�t��@qt�"q�yK0��{#j�v����.E�4��=;h|W)K;�J��+���)q�kl3��5Ze}�
�6��-����!����(��T�S��1h����� �b���`L/AA�N�p�́LҌ\����K!_wQ����R����M��>M�&�9Ko	X��?�xeK� t��f�����9b��?;c�oֱcS4/$I�T2�M|lƅ�D����IVxv"��$!ʓ�K��S!����\���S3���_��>�e�%�[������{�v! ��bs�x���Vh>8�ec��q0�oG�,?ݿu�O �A��3>�z���*T����9���Rap��L'*�ʑ
@EG�0��hA��~3�O����A'��#+lE^�?��M�`ę��W����D���2ɏ�%RN>� `�y��J!�DC;ڿz����<�#�(m2�k�����u" B�]��Q�85�d�A��W�u�����@��b�ư��`����\Lh@���;T�Qu3Cw�+�Qo�'��T����"�/�pj��/���%�7�Ld<��C�1l�@�����O��u�͂>�JׁF|U�u�?J��˼`k��y����� ��������?-����Ǆ��>%��#��;�d�y��pm�Hlܣ������S]��iт���3.���ÿ��M(�Y7Eo�\���f�{�9�չ����I���GT���{��RD��g�K�eIC���n<�]�E)%��	CƻZv!	p!tJ8At���ԣ�'�XE�7z^�Q,K�_��S�z~q�7���BP$7�:��S󮪑>�|�DF����E����b���_'��!��@'���W3񏠎�m �l`}��i��{�/*�v�R<Y�m]�Ѧ�X%9�F^���P_�&7�.[��Xڅ�/az���m�!H�q�<�t�q��8RG����^o&��WQ�;e�"M־�i�Ü?K�Sy��32���a��y�F����f�̎�|o�+^�3&����j��__��j�mS�b�쉚x�yp�uE"z�[�em*:�՛���ӈ��s�wq��ѽт��1�UP��ڭ�t.��{k��
��a�����+Ix:΍���ŵ����$���
:"�Nf��邆Vy�K {@��+3����6F!uT�j:wGjiPI*L�	����ic��I�⨴;��-���s a����y�x��q�_�uzAU�#COV���B������O�㼋�r#q�[��A�5�%�L��@S��)4D�c�k���SǗX'c;��E��*a���Ko&7,w��ێ�����2D��.v����d���YC��
Oo٠Ņ�_z5���.U������=���/�$ez����&=����"w��M�T	����),'G&���
����El��[��B��ճ��L����'��.w�rMW�@6�#�c�?V4"�l����Z��⽟�85�T�\=�|��<rf�xI��*N"re��l	�*�6M:ל����Ӿj���p�7�S�o�P���j~�5_��d'1?-4��nl`F��>��&�W�.��08�o���i��S��ar�K�~�Ч�E%�;�����Eߑ�H~.%�m�ibX��mEݞ>O$�4�/��j��8��|�-����jm/�4��ٻ��#�!��Á�OF�N�@��L��ĩ8�Yx��l�,Xq�7�k=��c������*�� ���/�{����q�6=���1�W�.�`@��Ų�xq#d�q�$d�#�5+w���1\tNn���u��ОZl;�=H=������"�;S\����a�i/��xH�'��B�l�]j�r�sޜ�@�&J�� ~SUpLx	��0�?�[�v�E�r�H,����X�Ce�	�4N��%'A�r�X^
�$���x��{�.Qt4(8�	<��!����k^a�&����`��6k'�I8�k\?P��/$VS���;*��
"�p�u��0���.�4A�׊(�Y���?�ظힶ�|uuh��0�b:�y��̕��
p�̨�b(�a1����;��Y��l��vE�{)XW��6�z��ڕ� �����#4��y'ak1�� �'�m�5�(#��eN�~�' �k���suu�EO[�����"ؼsZ�����x�
pϑ�N���mp\P
��^��� �~)���$��[��E�n�cs.����?��+�_*�H���1B�L�$o1���'��Q|��L�1+��UMl[:?��K��4����3�Q�N9����j��W7ٲ�����|�O�9�;�A�q.���A{~�!�S�! ������ �v�����G����'��R(kg�?���LR�/YΘ���2��Ɗٷ�u�!��e���R]����c��t!�bU)��ݯ�RsY�E�z\��y�*�/���X�Yn����L�q���Y5�d����n0\���˧�Vz��zYI���?'~�]�	f�`]D���̍��*@@E�F��7(�.�/β�oC<RA8�8������ed +D3���?���xJ���A�O}߃e��◻��>a�s0���s5+ݓ�b8JK.��ϑ��,/
��*y(�B�Ӎ�YC�����|��h�#G�j��}�H�<`�8 ��8"��A��&>u�q�ăxd��a	#��gt\J�<�^��<~�~�Ƒ�#,�e��+#�.~���`�Y�oNу