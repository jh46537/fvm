��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�On��Y��A5���Rw�k��{�,�#y+=�!����0#��l�C8����}�1��zk��n�Y���l��Rm@�����V�7�/����5�����$I;'2��4M�5
+�s��<0A�E�U���gUf�Ŕ#��;`�m��f'�	��Dx�5��W�uhoY�{y�'�n�͊�Z8��a��@!��~6E�G.>�ډ�����̒ ޠ�^r��y��.�n����4�c�D��H��ƾ�����ٍ��I���]->�C:/6����&lo6�9VI������w���� yx��ɏG��/�\���1��*�jA�d�cn�P2f@~��p�T٥"x�׏5�T��`��MӋ���O����gv>s�{�A8k0�w�׮G���b�X"	������J�֭��*��n�m�����1�r��E�\��Si���Aa��}V�H}�/� �h*�Mbͷ��!̥�|8�[)=f��Y}�Q�]:�o��������U�ߑ��"��"-�]bePn��.�f�*>M4����Z�9���D�	<��Q���T��Q)�/�U�]&cښ�B��bx���ѣgJ\b<�"@G��=��D�������販�o>�y7e�L�������4�7�R]k�E'���������ylGP��8�e*J2<���qG�#�8��A6|�,�	�]g��^(���٤nvN7�}z7�N���ˬ
z��s蜘��a�����4`�{[�$��������+�He��)9��W��S��D舏x�s��_L�/��ǘ)y�
1N<��$x��;m���v�b8�b�$�7�^������z5��j�#Z}ℒ�y��_<�(*�'�\!�7-�6���M�l��ʡ��(�9Q�cT�I/����sc���h���g���Pm�q����,T0S<�8���u��p2y��E�Ӿ�f�#az:��R���;�j�?�X�W���eV_�p���v]J��
��2,��Q{\���w����V�l}>􇢂�<Q��#S�fv��^b��x�:������'al���QSA�ҳt�B�>�ҊΓӿT�bn&�=�R�H�k��7�g�#��a&���ݛ��.0�L̋iΪ,(L��=��mәқ���1��B�+5��V�P��q�J���X�0�d��i_�]�S�W����X�3��ˋ�D뚪���=C�n�ս~��LIP�-��Τ����91YG�Εaᚡz���ߪg���z�P1��u�~c׺Y��R��3��@������%�Q�h���&�1��?��A
Y_ M��x!���Br,A��|Ic�}�`pnB���E�D���!n����X�<������,��<�9ܡ��H����p0a7q�u?(9n�y���3������=.�LC�M�O�'ɩ�?O}�'K�!�7���4���E`������mϜ2���Ĳ���`59:�[B9kI~;ռ�~��<���r�PE�uQ�Iu�8���7.7��"e&���,S���=�{_�?��z�W,�K��( I�!,�Z�h�o\^��r��x|W�-"_����/�V��*�G�F��=���s9p ����@۽_,�'G/!z�GΚ����.�<�%A�R�W��A����'ql�}6G��
��O')L�@z
�d�7��I�be�����J2��?<�ӹXrP���iH�UQ �(�e
A����ŹF���	����F?<]VU������5��2ZN��f�%�	��:	�2��z!.�4d!Wl�<�2&o�n���&��ƌ�	�'j�IF�D{M���ҏ���>3�£���1�4��=(��^�����c�&a��aƮ��*-�F��+'K���$�N�W�|��Z(��/�}��6�[S�tG�!�0�e܌�5�ґ�XD� ,J�8��1�������Pl�H���C�mq�C8�<d�����Ev���v���ca��Qq�Ћ��j��5\�gVU�^�#�*L0�{;�|��r�ťA>���H��ud���3�2҄��5Nؿ��ni���I�����-$U'V�`{"(�%� =�DD���Kr�R�T�\6�a��!S2�����dLd:5��X�.6O��4X{xF0��8,��%�_5�~��BN�0��-щ�Gl�~=I��Q��he4��9kN6ڂu�5��"^Ox�HbږrY��#{h_w8��tcC���G�����BE�#����RK��i��0�3ZO�c� ���I6�x�r7��zE��y!Ӡ�-z�������B��MS��=T�4C�b��xҝp�7q�/�8����gq�.�����Zw���<���*�L�g�fQPa^U�U�+,5IA~j��J��2S
^i^/�+��v��:E^L,ݙ�`��v����zi�j��&�RaHal1�1��$D�Sq�@�ȋt�veaoN��b�Ϣ��� �� ��9p��)ލ�J�b�g@�U�եI{5�*6���!�q�$�M;��+��b��O}	17���qBuZ]���7�խ�Ө]ǖq��c ��C/P,�׀bA�W��Ɵ�W�B8�ܮ^m��dW���dq�h��	�ła��{n���1Y�;bka���0gh�A�rG3ct�N��W]]�tbҁ�܉ltw��
�i���}��� ��!���
cX"��H��>�`��du�t�f͉dXd5G��2�e˔M���>�Z���O��-a�|X��N@�u>&{EN�T���˟��v��9&�5u��'��9���Z��lw^YZ�i�b��A���11��D�	�.c� どkZ
g�S�rŀ�[�[�CB��D�)-H�7ǝ�>���CH�������fAR�I���W����ks�����1o�^jv��@(}�l{$��93��W��eo�M�$����d�fO)A��]�*svrD��+�b-Zw�8��<Ұ��2���.������F�X�ҥ�Ƃ����d���jT�9�x.���	�U.�?������)���hYn",}���)�� �, ���&�zj�%q� ��L7��p��-|r'�)�%[o.�f[Bp溭�Z�	��K��W��s �v�W���t�	_�q�}�&q	�cZ�	'�oVȨ�*d�Eɉa�8Ϡ�YD�"��w�=J;���Ϋㆀ}�+�S���:<n+�!~ϛwj[��aD�~������������Ӓ���
���:�n�L�iM�Xa�4����Ģ���B���B�qR��	�O
��'�L|�:w�b�с�l�O�*u�җ�]5߳�`���r�H�y�T�O����@)��5J��<���q��	�(�576]�GXXR�N�1zd�D Z#�-�~s7)��`������v�Xp����=b����(ɗՌ�w��ۯ����x� ��@Q�����|���lKx"Wu	��;�E���>>���.��+8Y���n��?(�.��zn#P:�n�%j ,�ւϳ�YB>p|U�ȋ��e[�������E��H�+� Y�%�'��P#�c��� ,�L�����?K��h$"�r��?I%Za��z����	h�C�L ��NzRov��-:e��(�<���l��"�X�}�w�J�Z�����=��vk�;������� }$���b��YCW�V��s�,� ޶��+8���gf��	��5��:�P� KͶ#!u�\!��oo[9x85,6�K�I�=�h���\к�+�[�:����7o^d�yQ��1n�b���:��+����`��nh/퀩�3+:X!�/
2�v�p�K��x>��s�oHi�ϟ�H%���o�6¢]\=����0c-����d��eb@cS a��B�ۂ��E�\1��[��.�KX�ҧv��Lc�T^�`��x���y�>lȓ�r��*�W�:�-V�T޼ua�z*����,��h�
Y�Ɗ�#H�=��,���f-�̪�z(]��.o！�? ����}cVeF�:�._:�c�|�,�Ά�J"g�",����fæ�:����"U�;� 6�f�M����� n���FUqt�YW�A�֓�W@A+��|��8�����?=c�}��c�TW�E׃�o�k}��N�S�o�/��5���I���1��q�E�]~���'��jsnbd���d�����KI�{]}�w�BI��m�iGi�����1{�N@��e #��Q��;�� az��6�����Zg�i$$�_��9$������ނr����|J���+���ă񊿁*�fV��C�_8或$�����3�e�C��;������q�P���Ɛ���@��6�:7Z��a�{èNXCt1t5x�� �)��rj#P:������"'����x^�}X���u� �$�a�*��u��.��U��sy��A�y|"K�A�\��kx�{�P,����ރ�k�c��L�m8e���y�H˺��I�e��?�8��h�$c<����f<�6w�ו �4����)#L������W
,���B�"e"4'㱪�r�������[�^Xmđ� \�d�ދ���dWNΛ޺�D_x^#����KT�4��I��$�>�Gc��o����!��c0�@��Uv���\��/i��mL�2ѹ
��r�|��?�U���n\���3�X��)���m
b��
�E{l�^�e	��YIn����-��m�9�^5:I����7;08�>tfb��@���^��9ޝWv�:������j�I�df�0U�"_�Vs�9�IG)�T�����Z3��D�!B�� v�c�#@Ջ͕7�x�o����A�Yt7�����IGd��ճ=B�E�N�ߍ(\����f�z G9�{z@�Ҿ�.�v��䎯��	bL:)m�s�� o
����m������j����!�	����F J���)Y1�o����tOi��`���4��^^��,�������,�UR����d0vq�JKV�u{� Sx�T~H�H��w 1�,�G����I	hA0Y1�(�a�e~�K G���S��~��F�,���%/�v8I�q���r��^�XT���;1x�����Y�0}K����N�/�*�'R�O&]a��V��`��>����a��ەV�����c�T�}� ���sc��3��g����9��f{�-�X�H^��>��W�{�fW�e{YЩ�&���p/v�t��!9(�ɚ[l��\*�?����*�`��D��\�Ǽ> g�_�:^=�n]�.���2�3\4o��Ӟ��Y���&�<�
ض\U�^t.+���t,M��r'&��W�����obu7��Vۄn�0'R�<�\Ȱ)Q��M˒�@J�̙x��G3�4�cm�X���J�r�d�[�;�
�[wq�����:>����:�q��,-i�`/��䙱�p~������t�V�ϖ�X��;�f�*>-p1�0���f@z�4�	Ic�E�ˏ�_Y4[U.W�YF
V1��J���H�GL�$���^��z����R�;�M2;4�׹=��x�ͯ��c��(�"=g�L:�s�R��2�}�g���(���P.^ :�ػ����	�#�(�	�O������4ETO�Ry�"/����d33����ニ��nI�n�xd��І�ut�g��k2��@F8U@�Aw�j�p�ٓy:`�KǑ�G!}7�'.���Q��>���"��o ƭ�0[��D$���Qf�	����"9gSgً~#c@��O��w�!��-KF�p�Xj�E$�\��q�cj+��Ā�e3Q��p��v����N{��VdV�����}DE�(������1�Yv��98�<V�pͩ��2x`�O~�A�"d���Sv��B���o}��+����Jri����ޒ  b���94�+��%yO_���A��i�/��ͷR�_<�c1.�)�&��*'

��u$�Sx�y�N�|����,f��ӄډ��Yeh�Bcٜ)Kyeg�,��O�'�ć��/�
��ؖzκ�Ǝ��M�S�x��B�܆��c6��#ۨ�q-q��i{H�$�.ll�������X'�կ<��}���Q=���M$�	�|I�ᎯF��\��EБ��-f1�������^)�`O&l��QLm��sQ)lN��(��ޔ����b��:�az�z�o�n���Em���S�G9fУ�t:i�nT�AeU���Ã���ؑ���~Hb��I��.^��v%�>e���V<�%΢���[4|��c�/�h�:5��x��ׁ�`�=^� ��<}�9�Dc�6��CU��")V�TZ�`hi��Cl�}����'e��� K���[ٔp�����aZ���}�p0h޶=�\l��K�=m�bc��!�6�f�@�Xަ�ǵjh���@��q���N<��^���\���#:aؑyJe޳R.�8���ݿ�eQ�Y�gN�Hv�m�D��V9�qDej���`�& I�NŘ��ұ�dg�u��X�[ew�*���̴46���
�rC���yN�p�0��P���S(��e����e��$Q��!�&EX30���=#�d��¬�.o/�z-`@ɪU/�C'�4!���A��o�����g�����萊�^�W�"��{�p�8BH��S����0�	g~k뷉�`(�5�/��z/�yh��UJfOhһ���ҩ�D�U�mks_*l������W̯�=���E��q�����3�y*�f-@��~ڀ����8B[�f|�������V'P]MUoJZ���%����N�7t�q��lv��RAO�e8 �I������w��x=�XYPtT8)Q��ը�(�	>�+�+�j� }YF݄��n�a�Z����h�����ag��vS���G	��UpL&��QB�N/�s��\��>g�_��1s@(f��N5��O �B\��x��]�8��p���2M�� QU��"a���Ї�D:L�^g��o>O���p��)C��Ga�:�Ƥ��lpD���~������d�j3�N����u<��a]�V+�˲���n���lx�{>�]e�b �{���ds�R�~i��8�����ػܥ�]Bۇz*]��V�7b�c����T��;���-|�	!�{2�8�d��Ν�ouUI�W�C��n�!���,ن�.ҿ��[�.W��O+�Cj'�mf>ƣG�|�I����Kv=�}��yw�����[�;kw)�.n��ؠ�&]�US$&O��6�;��&Yo2h>�=# �ҕE���(��������-wj��/;yX3x��(� ��j�	��h�U"��:�y�5)���	%"��=�*�A&O1-]�ؙn�]�Y|�-<>+���V<Ɂ@0��k��W�*�X��lѳse�]M�3^.��`{f�_O/Q�Z�OZ�줋�����t�	�j�6Ј�� DX���X
,ec�C#�e7P�*d�wb��b�*܋�U��Qpޓ����f�������ʹf����cF���JA#��$d��@4��)�h�l9Pg�
ߊfo��Ø�+�,i%��o��7Ab��:�	}:�K��.�[R2p�﮷û֡����+,8c�A�M��P}Ԫ�YU�[q�%H��vF45�D(�����ĥ��0����cJ4����1U�o%�?_%-��zron��"�o��{_9n۠�H4�^���n0��A�����7�m��Dךּ2@󆦭���Z/�C�~iO��=bm�VX#�uu��2�Un��V/�r��V9�	ϚA�oĹ��a�N0�;��,X�(U�) [���4!F���_���
�}:O���Nado�y)G.�a�}㎛�����(,�"+����yȜ7١�Qpv�9��]ډ��{͂�א�G�:�N���ow�Y?��#��;Ѹ�A��A�eJ���������u�!��e6N�oN�Gf��eQF��"y
g窞�zo�U�ִ�TF�fb�H��ₜ�4*G@Y@A�b�uں3pb�U1�Zl����o���3C�؇�
�5��UM��gM7v��u�ե��di6ս��`S���ú҄V^@g8?ѱ��<0Wu���Ǭ�I��g�t�IZ+��i�ST�e���A��Ct�^a�a��#�ځ�� A�=]�d����}#�,��IC㌡�S���o�#�]Z��;�ېJ���)��F�JNp�9������:>�;8���C�"U��'���M��7�����H�|Un�G���La]�����i�g먫ɭ4u`F�ƞr�G��߰�OϺÙZ���Nw;�9s��*���d����Fb���:˷��?M	L]�H�����m]�F1����q&���5o��V�0c���
��7<�7FN��i='����՚}�ƮY�~��#g�P#W����d��ޔ>F�ճ&��ʺ�x�J'�Y�%)� =��L���;8� [�V��s�YN��]�m��sW8`\������u@���u��=�J��R�q4�Y��+���w�����$+ �r�{;�L��{���2GC���	�����S@ ;>W��I�՚tq��R���1C�4���[U`��yإP��>���I�6��q%��(��~B���q�v-/W�Z�ғ��3	E)ѷ�D��bv͍�S���H�C?��u	��tA�_�_�y�Rq�.|���<��?��8E|䞐L�8�a����`�д��?,�8F���8��s(d����&�_.h���dre	��I{��佅�T�c�&�n9/*�ݫ6z���0����'�/�]		J����6eǤ�EZ�w�쾺𪵴c;��'��f!�6U��#���F~�V�3�w;yP�yQ����X�����ޤ+�����$]�yX���UW"HE)�C��н7G�ʸt���+�/�=+�|����#��Ӊjq�rtg}C�y�z��֭���Ç�IGM��0< [�0�^`�\Fv��`�z \�z��"V�]��EK�o:/���_���	H������Ί���q���ɨi�~��h��/�uQ���yp���E��%��9!X�����1G��޵�ע��ȧ���;�
�g���(!D�9ͣ�Ł��s�q�d֧��L�$�9�z�"t��k�@��h)�?�Z�A�Fj��>����<�8~駰�ҩ�g� )8���s'{��y-� ^i��`�L~���J����"=e�2����7��wi�;'�tl�:}ʋ>���>=�r/в��B`L�p$��m��s�����o�',$K�J6ݲ]k�N��pHG|it�4���q���=����ф�ϒ��c�S7��o��@���x����qq�#M�U	���[0ۊ��TkA#�Q��
|�Sd�A*�1�����*��4"e����*�d��S^&����}�{`���I�8�v����*4� ��Rv�-wD$�@jFé}��t4�1�{�Z+a��^9C>K�8�Y�Q/:��j�%��͖B)��˅�o)b�Ʒ�K�}9nJ�Ttp�vK&ivvwj��)f�9L�Lux>�b�r$�h��(�[1O��ܽ�.וn�;y�U�\�l�0�jϕ�0�{$���yKM��v��Э`4����w8 �-���d�ވ���v�r5�����rO𗐴+���R��kwU�p�����@;����^��DI��7��2��?�"Cn���LD��غ��������+��K;_�(�~Mnҩ^�� ��Y}kB|�WI��o�c�0�1�e����6���4�������ɝ�vx���	Y��f:��Q2}q��(�o�t����`�*��~j��a���A��F�����cEˈ/17�$�FVbہ�)&�j�[�&/nv�у���D�����Q����>�3돔@�H(36n�dʅ%*s�='�:Ʒ� �(J��L�G��׮�eB%k�b���je��	��q���/���4�Ts���9u����a�-m�ǆ�(<�O�v�W����t>�t�	ڻ5ފ1�Pu����1�\�8~��2�������07��XԖ�x�'{�pġ��z�T[x��.aL�+X��	eX���Xlpu,�VA3vô��?�G-��r��&�ݨE�����0���q!4��{��Wd틂�!M�c?�[Z�s&cv����)$g̻��b�8���`�œ3mT���ˍPu�-�f�љG��q�s���@a�La�;P#�oj�{��9������5��K����}���)M:���s�0��0ç��<_�d\�����?��L�MӔi'��Ի�.�9�1�}�8/�kz�Ku4.+A����a�B_'&*��K7�yua1�%���^�j /|"Dli���u��[^3���tf"ں�����mƆ�n��x�'5�2ŧ�I�럖;�
�+V�f�����j` %��_�f4~ja�0�q<���hy,�R�O��I�e�7��Nh  �*�׃qd��I%%��*?ƛà���‮�s��Q�+5�����@��!���3��˧R(�pZ�5��w�%I��9�N�W�_�)�
�&��'�?�` ����%�!��R�b$v�́h�X�ܚhHH� �]�h�N��������q�6������P7�����l����3��'� l��t+����2,����Q�KJ�K���L��|nT��x26��jvJn\\f���+��Y��M��Bt��ied�: kp��z��97<4�� ��4��7$
U d&�����(e�׏��f͇uj�fʽ�7C�Y.��V�,�S>�D��N3�9Р
���mtj4��P=����[jms�M�/���?&�wZ��T�H�JDd��=���ޖiyJ��ۼ����0�deo�B���}S:7�2Ot��
�:)<)�i�v�ĝS��k�2��M�z/^ըvE�Y�g:��v�����Li{��$�g�|����,� g���*!��͓�*�ၘ|��q�f��-�gZ���N^� �j�C�/�&��m ��u��.7�T(�Z��g��㤦�D1�0�}�&W&Oܕ�bU��.�`�\E�'����}!�G�\��Zn��s�\�;��89���$���u1�|_�h�&s�:�Mk�[At-��z���f�V��[K&a��1�3ג��X��W*W���{k�^�k��6AY�:?m��)Hޫ����?9�í?���BUl����-���uL3�d��8��V��>�R��CbjsC24$���%I���M��c"a�����]<pҨ�4�t�)��d[��86�����fd�]�@��']��O���K�F2'z4�R�s+1���V�aR'9�;L$ȡ0� =��q�_0��tc{��퇾˂{+ �,���	@G+���T����yy�=�����Pf���1���t�8=-����J~��h3�B��T�b�V+hEC�w@��emG��>�P��OaE��g��\]q����e/A.��2/�vH_��[G�Jڲ�2�!�&�ʆ?g|���(�"4�C���~�)���|�G���3�SU�c&�,P)]%����ҜcQ�x�ed+�)���y4�(1[�>�^V쁒���#W7�g��(�4�`�粴7���Q��������*_("��%,$Z�u��*��m�t�i�4T(.@7�v�7}��T����:����Qu;�cÈ&�I���๾P�%
>�Y�Lve�dc���Vq�}qS����U�I��voH�~:���O�8/��e�l��4�ś����%��_Ȥ��8���h1�in6��a�������!�Rظ'�Ĭ��f��`U(�C��u0u�4F���k��qd��WrM/G�zq��@|��[���r}>a֫'֛m�^�=}�f��d��=��3˚S����~�g���߈�j����d �e�H�d{y���d=P�Ğ�禗�I��B���d|`]u���=78�-(�v.�i���TsC��3%a��5[��q�m�a�H�����r@Y�	��gZ1\Ԭ)�gHT'K��)�?@½�Q����B	V��ᝬ2O�� $�"������4�zو@��0ǟC[��zn�N-^��fd�"�9�A9�e����x~Rp�WnKz�Q����s|\��!�n�I!�S��]�5|��<�Q���'��w�P��U����-�hj��^�V�ܷaW�^�����T�q���=ܰp�ƶ1�eNQ��7�H�ǀq4�B�Y��j�7?%����#lE��q��3/�
�ؙQ�a��oBNL��z��Ab�s>����3i�ю�T��Z)�I�T�]����j�P��"*��h����.�s�']_:����+�OR�Π[cp�(�_Y�8��2	t �l�Y��DY��DAf H���3�#�"�b��e����8`էK�fRz_81$���#��c�RI
�"4E6��A�Wv�ҕ�E�e�n������r����Y��g�+0	#�J�y���sV��xJ��>;�W(:�d�������;��i��iv��t��y��u��������kOԶg��2-P�=�l� ��am��i����J�z����Y���K���V�Ax�����4���hz��`�?+EW�D�)c��(	�׳�2{ZVR�:5&H�y-c���� �l&��v����Y �� Z-��(_���J���v��>�I;(�@~ѯi�1�t�wȶ1�=k�>�i�qN��� ���K�%�����S9E�2�NZ����US����f�e�bŞT�'S����BP����|K\��(^�h���L<�s#,>� +sQĴ���~g�w�d�
�[c���0������}Q6� �N��6��n����ud��lB~�U:�^��t�7a��Q|*gFwPXaX����S�9��S;��R�|W�ϟ�gm�n�j��X�&��9j�o�H�����R��u�J�0������t�Qe:߹k��6�]����]oo�i(�٧e�P���.K����d/>̴��O���=�\�g�JRe�v������8\U�,���_�r/�^6�@�[ �Bn$ʌ�H�e��L-S�$��i���涧��c
�"��R�������e@D���"^\ר�� ��8��UV��䫛�J��4\�=��x��yO+(�pK��9M������D���lv����ʂƳ��=h�1DdE�
�e����#��I���P@m��x>�@'���IZ���-Ar.�_޶�yVIWٔ1�G��t�������+NF�����@��>R��nB3�fv������%��0���΅R�ۋQ���.��2G�B=�R��rx�Cq�~�S�'��i�Ա����w���;G��6�����"~�%�����E-�F}�F�g����#�\�y��5Dgw�I�U#�,�h�]e.��B�n]u��b-\�����^�S>f���?�8=5�$�n��g�AR2�!_������ۣ��j,����}����F�;.�Ѽ`�JxO-�3A|`%�Yz��K�ǋy����U����i��wb���6�:�Mc1��[\u,�e?|MblS�)V�Nh���FKT;�<�0C��
2� �&�a���.U��1;�s�w~	=_���fp�*���R���M�ES���8��� �$,�)��J���:rL�z�}<h�V7Zq�?j}��h�Y��ꄩB|L��6}X@7R��sh�t����]�W�w�68&�`9�ZW�I������}���20$?�b��V�9x���tv�Eh;�5p]�A��`���j��P�m�r 4�\	�t�O���6�w�E~����w�q��^�r8n�H�ɼ�v�D�״0ޟ��� ��c��aZ�0c1ڜ>���Z����	�A:N�d�eR���?����t��NQ �����?L+�2A�@1vk�W�D]~�G�Q{�\���ti^�򯔭zT�sH3���Q(��)>�#KEa� �h��şf_��j��fts4q�^���%��g�+�O�B0q�9�~�Ir���%��`5K(�E=�
	�Ġ<##��p����Z�/9���g������!a[6Z�˿!U����D�(�#)&��c��:)�ͻ�c���?��h�$S�k$���G3�<[�`}e�ڮ������"��2�J`X�|�0�\֫a�N�F��~8/���C�c�NtA�����7��v&�[D�|��#v���}}W6ܫToXŘ�DŤ. CQ���k9�m�4�l��etcm�XP̭ G�f�cH:�0��b�&y|�&x^�}�M69���*E�DT��L�Ao�aT�w��8���Neq�W�[v*˓�`6���⃦�ٍp��:�*��uR�w	��r�f��{�etj����#k�����z�]<~A�8"5o�	���� ��?�frH��Cѣn�*A�v�EO����(Y\���#~�ط�0E�!�T���O��]���~[�h�a�=�PRܪ�2]R1Dt�����SCG<U��T����q/���DZ���"n4?	���?#[�5!r^����4W�#�+���xw����;�y�`J�K��`(���6��-1���u��ݠ�{X�4Ɂ�D�ݦ�j/Ǐ�"����R�/���Ą�?PV���J����1.�V;�hn�8J4�P#�ZK�.�O�]���'���D��Y�{(/u"��S��O�
)���/�����᭖E1+���Ctn��Fƒ�Nv�ӳ����L�ˋ�[���9\w��{������BQO���)��Qfzt�Ŀӂ*鼃�hQ� ��lЃ�wo��@L��hh�9�]*X`y���&�"�ȲHQ%S���T���7ID�����J|��ݛ���^`��k�*&+�@�wgw���iۘm""�[Rm��u���N��H�V��͠Fq�U�E����7�LW ��ToF�=b��� ��F%י���Ip#�!4q~��^�9���#*�[BB#헭�}{���,�Wy�F�U������\�(���j����Mj�"h�G�@�x9� [����=�}B./�vAy�E�<�p�Zͅ��W�R�(�u��޲���T���ℓ����ʚ�̚[�,�H�O@.]�k���ՁK�g}�e������$U�;iV�1�||~�4gj�����K�z`�T���G$� �2�^,���U�ɱ`����z����.���SW��K.V�����  /�K����]��ٲ��#�Pg��-�9o�ye
�b��gv��2�T(p�@~0n#ێ+*���%g�KV&�b���&x�iNi]�&-B����'t�;��ڙRZ����Z��=u>�>�Գ�H�S9U
�!aA�T��~�
8�����%)~}YϏ�;�B/�y�'�>8V�Z97�&�Y�	�U�Cb�Pt��;ǿ㵺m�4�ZF��z8�vn�m'gs�F�-U���ݷ%��k��A���ݶ �8jKf_{ƹ�ȋC��������Uȉ��u[��$�ޑ��#,�t5&yLH���*�� �bT��>�� � }�X:?���;Mƺ0
��K���-�����`pO\4npϡ���@0��q���G��W��$�^v��n��\r������J�Q�P�]N_�4�6G+�ͯ9�#^��lOA�%�ߚ�U`K���/M�.��jv#:�1E��_����*�����\$F��m�Õ xd)����U���+E�P.e�z���y��m�J��O�v.}�BFVȾ[E�W�]�\�D�\�#p��X�ԍd�F����t���)_,O�3�/�m�|275��!ǻ5�Wt��?�yQR(�����>�����P�t;Fv�(7`W�QN�����ߜ��/�"c�	B��d ̽5��5Ȧ�N-��A��P�v`iܺ�\�R���M�~��ܦ,����`��҃J ԩ8�ň�t	�Ҿ%�k���G����� �a�f�~��EX_0�6�i�${P��8���ٯ�[�l$�E�Y�q>g�Z�3 ItɢB.��T	xu-����A�R�Y�T�k}�n*3@�t>5�6���)�eWG���
qY_:|�k��i��cQ��t�Y#Y{����w�2�����lނ/��Γ8N_��)	���c��+��k�҃W0�JB�Ԥ�vZ5�ץ�����'������?�����c���9��9�O��k�f�Oz�P$��M�y@DD�k=,	u�w#�ʽ-����(��~���꒽ǜ��t^��&f�	�O�E�S#���[�k9jW�@W��*�@�D�ps� ΔuH-���z
*<�8���@�#jfw!/�����B/�82
�.��ق��
�B�(|o�B��s���s%�o�dr�*)P9n�g�H�����Nm���Mu�͆�#��U���2�B�x�l�
�^��oItVP�
�J��O�	&Iѱ �f��ȝ�\y7�Dn]
��pYD��[z�z4��T�; ��+Od�-�|L�Y+�����A~���L|{�_ɖa�qME�~���b`rG�2%��y��r�m!�}1@��j���
�-�����UBB�Iѐ݆��N�A����i��-����O�p:�ʹ�y�F@鱩�hrԒ�Vf��[�V;���SP�s=�X]�ď�����_����~ �P/�	�U�Pu=3s����6�,;X��kH��e��r�W�@�Z0�����1s�4����@)z�������#CҵL���n�G���='��ŅPM�D��&	G���϶JN�UW	W*lx�����ĈA$�ѵ�B�#7�1IU�*�ۯY���B�� ���78�իh@pV�!!t�'�2v�{h����H@�����*H�*��[Tlk�XG���o�VF}�uӴj�mW���Z]��O����8x������bVvRc��jb�z_ �1vr_3_��Z�sg����t���ϝ�ZJU&-��q��ɮ�9懈�}-f�˵d��>��6֏Z����6���Bn-5��Omi6	#e��	#D����|	�1�E��Ы�
>x9�ҕ��Qw�aV��J�ǉ���s�r�BN�����Zgq�F׊��'6!�y9���	�������Ӥ]���+vA�m�z'�������{�|�_���N|�B�4I��@��;�[Ֆ�0�"�VcM;9A�I�@\����xt�l�$}��$؉�r>�����d]�DS~�HF��(�Q#�H��p;� �݁n���K��T���(�{$�z�pC"swܑ>��r���T ���d�� 1j�ttT��ڦ�����`�V^!3m�Lw�P�<*�$�u�����1�5������9��<r�$�B��N��,��o`�=��vE�Vi��qcyc���$5�s:@����oq��>o��Wx�:�C�C�+��5ePǇ �f<�cl��i_Y��d�v�"��@�r��R�BPpb#)R�c@*��#.[��<t�8"�'�I��aw�n����5����E��ɫ(OW�Q\���i'?���C�{Uެ[zS�BYH���@RK�=Z������k����F�-�����V���Y&��(P9��΃s���EQ@&Y+��s��s#s���/( {9P��9�57	�G�U�D'�V���{M�űk�"������_1���e���b�AP����]
,�ad@.\�Yҗ��X��qT�W@��^I�[�#�� �����l8�c���~8�F��	��E�BMj��sf`�~��Q��I5W��.n�p�4 9n�Џ�^`p��)�Z��wlO�'����-T���0a�h[2Yq�\���R�jX$�A�mE�|t/�a��&gV���@�)����=q��[(���Va�n�
��x(|((˔z&[��SM�,oM�Fﳃ�k"u���+<�8<N�,"[iJoV>!��Rq�ց��^�(<��.v�y$"Uƨx��f�C~��e�D��2?�g��1�p�����'L�z���ʜ5�ںÎ�/G�>�^M�ʞ�v�A� \�jTó�ʊ³�V�8g����:0�T�>e,��kvܴI8��f9��%�K��<��9�2��l(:>�L(�]�n]k��Ҷ۵�mW�f���b�a5�]�k�q���B���Ϫ�׶vF�^`�^*�kA�
MK,$��L�wwo�hwK�W�CMP��E�Y���-y��/TJ���*���>p��#t�m/,�<^������3����k�57�g��o����i[_w��L���3sT��gnS�HO�,� ��b7c@L�ɶjĵȧ�-Jn$u��n�q NDp�\��T!ѿ�Y~��@�� xx�R�ϩA77�U��ܬw��`g��)��4���	~�
���M�GrU8��|�W B�ݑ9�`��E�gH�0���LU��/���c�*���2��O LѶ�n��rY*:y��
�	�s��j����i�Q_��n�d+��p)���8sBu����$�@����V�hg���L5Ck�`$i��ZR�9|�l�Ww�B�+�J�s׎*�N�ǂ~-��F�������M���V�P�����HO��G����a��}q~FCc���^�8��������H�
[��.�G"y������J�?g �V���L�5��yv��.6w�&F�|T���T|���+Cu���.sGX�S�A0���s��OG/������y���)�HLGN�h�6�Z9�[��/I�����ڌ��؝�[E�����$^��gc�a�	���ॖ�1�/A�	8g��G�����w��8Q������G��\4,�4�hQgV�ђ�x�~ �3�ո�VU2�Y��M6�
R���dӀ�, I��<��b1.�ۖY+&;�o�*Z���IU�'"�ϰ�-)��x�2�o���_�S��6���[�.O+eĎa�,��c���d� �D�|Z�Z6�|����]@z;/�ghdO��yB�Xi���;"�\j��|}���S�p.Թ���ڏ��rh�63RIp=���y�T,�fYO�/5���_lFbME��Wn�y��j��L8�h7a C
1M����j(ƙ�H�(#����,|��h$P�0)�.�8�Ĉ�x,p�L}?��wO��ܨΛ��/�n�z�S1�##7���-��aR8�@K���E7 ����8�@�������ӗL�+�j�r#�H��/�q�1�؎�����$$E���&�S3W)��A6{S?����ݝOS��L
���Sb6�@�����5���sf�6�0�^�e9~��ʽ��w_q�Z]��|,��hކ:����l�x�|�L��He'}����,����%�bG�x��Y�g���q``�L��I�l��N"IpG��q�*K�u�H�B��-Z����8����3���0u{��w�i���m�xk�}����a;'���.�ߟ��\���B�N��O�
��-�)��j8 xK
���fj�H��^������J�CU-#sn����G�]�Hn	���U���
>nf�����W7v|1^ǔ3@�"1��e��:ʹ���t�'t{�{'�1ޫuķJ�5��+�&�9�ͫ6y���ln!����(^%��oEB(�f�����#���&;��V�b�ѣ#�&�{3�Ⅳ���ȧ�W��at�-E	l�l���I��Y�vS���i�>Gw�e�y�fxg|�� :fޯLI�6�<��8ZJ��^;�P���n���LkqH����>�W/�^��r+4�vl�B�y�����!�꼥JJ%<�Ў�3�g�Jq<�J0#�n#o,�nJ �[�V�O�|b����S4d�'�,��ʟnx^�m8�3�����	P]�[ZOMϤ�9��>^5�I ,6^��f��{tO���U�"�����_:9Rsu�k�I���
D��$K+o�1an�N��W24�Rb����i,����:jǂn���olj�2��qV��}�Ӊ��Hɴ���!�����/8`��F����L��%�����~�!�#T""��Q�����Έ&%�.�� �\�:	���;�ʰ�"�_�	�v���>V�o���ϐ�"+���e���aV24"�:+�$C���(�7�p�ȅDEd�m��	­v�ц�2��������ѝ�䑺5�����p!�.ƴ�ԿK{��e��..��C����q'�O]We����e:�/�RJ�{�`�r���ӄI�?*N��Q�|mQP���kƺ�)�Wc��.=���RQ�*��2�S���T�8� $�[Ȕ5���s]%��j���Dr�M�{4΁�حj���$����FԠ� e��_P��v���U�u���Ҿ��n���_����V��J��Ѡ��Ѥ�u���W���-�Ŗʷ�p�������|�B�ͫ3�����"���w�
�K &j���;��s��!ݜyz�l�í�䀃pD�LC#����MCIuI�y��nAM����#+����*���ly'$�X\B�2"0��U v̥�̮�����Rd�#��9�٧�����Tx[�q��"�����ؑ��w���{2��>� �tT�Q����jɕa�B�=�+�`V�L���T
Ya��.�ˎ�r�к��,w#U���|�ٶE�����qe��S<ko�E9H�S)��J|? ^!1���F9��8�9��ڊ��o�g����.L�i��p���LU��:4��<	
��P���a���q�#O�	��7_`��~�o��S�lG.h"t0}�W=��"�F�5��� ���d�Lw�C��u�>���i*Y"ut�k�|@H���q�*T�\?�]T|��.$�4/�J�������32D�h�XN{}����Щ5ֽ_V��/�����2�G-ޜ셑�� �v̸�p��*��}�K'��G��x��Z�x�+/9�a�d�����R�����F�
E�>��$]$��-8;�~�z9�HO� !�2#����`6�Ћ�O��D �Jr�g�!��2���}���4J�}o�n��z��a=V'��g���X�ۨ�{��)Z۩��s��u�\=��:f,�D��W6H�H���f�Ig6y �A�v�d8��g'Ο0�p�U��xC�-i��Y�m?�����*Ϟ&{>ٶ�;TW��t
ԟ�^D�諄�B�%LC�B0+�o�&��y)�H95�/M{��,��:z.�Y�O�������ws�ڃ�/�w8+jv��/�Yr"a���}���$���k/��X�S=�U�L�ߘ��;������_gJXK���<÷���'JҖP��K�p
� '�;�$��,R����]4�S��3\�3�z8���=��H�{�V�J�0Ű�?[PpD��)¯u����ܩ5hU�x(����iXUa�RO� ZV�_S�%�hx�\�������e?3�'�_����>�L;o���E��ܔ���گ5���w�5�ol�X�;�?��@{��F�a��B�er]��Y -���0�J�� ^?��f��@@�fܶ~�W���4p�G4�d�ٙB�c��s���\�i�����<��w� �bcIU��>H�Q�s�̃֋|H�FdC�Ε��L��O���@H�_,��� ��]��h�ZD~��	�e�^Iֲ�g'����P�[�W�|y��+��0�&�P�ӥ�����WH�h@�Ŋ8M���CmQz�a���*8O7�đYE�+�G++��m+2(�>x�l��+�ֈ�'LnfR��y�-ι�TB��(�5�_�����\6b��
O�y��Z8�^���i�3z8��i��W�\N����K]����)ej�r�;�/�%�{F��٢�qT����E���
��k���Y�&��%�/߈�(a���Q
��o��_֚? ��Kw 4%�d\��f��!�r���^kM+��.�"6� ���lC5�0q�{rueͅ�d�����{`�^tI)<:\��Rq�L��,�f�v�m7{}U<�f�
�`-<�8&$�]��i��׎llddi�=��˹rI�s���k���ΆЮ>7��N�Q��f�N�2��!%�E܊Q]�*��&�#�愂~ ����%�}�D���3F+H���P �`�X��;1��A?�Jl\��4�E�b�2��!���-��ob���5]�Ρ=y��x>:�������CRг7��X�*����.����E��B���+��������`N�-�B˴����*�% j�Lb��*ҀQ�$���;G6�߅�z�
���B�ݧ�|ϱ:�,�������t��X=5���Q���Q���z/��0��$����_q�xM�+��m���nk@���1�}���R��0>����q����ןۦ����a�~����H�����d:�P<J9�L��ש"�K��y&�����.�cj�XV�g�l�}�L���r����6v���ߚ��mu�_0A8����7]l]�@*��=饅G�#H�
��Sn���H��0=��jp!�6�;Alf�9��~)��Y�:{�J޳ˏ�E�uf�G��2{�*kS�U���=���luט�w�}L��M��,��K�DS�f#X��fp��Ia	�[0��\��@v�h�J�}	��-�[�D���P�-�	:Sm��wW}X��ld���@T����� P������h��~���
a��e�M�l�+I��垕{���b2T�`��$���J���Ń*a�%u� ��^��*��;�B���K3?��B�&�W�M�B�7ˏ�6�,�� 9|'4f�$�����F�}(�Cu��:l!���	.���	��[�ް�լ�T�e�g6�uf�f}�!q,+����`,�������OO�F��:�D�Ze�M%0�5Y��g�m���ʏ5��C�I;����Kj�(�$m�[�-�y�4�]�e9�j�|a3���m�FkڛsJg0s	��5��o�'�*>t�o��x�i^���{J,#r�����R9�D��ҦM�Z�R�:�>���tu2�Y5%t�T$\���_� �+ҏ0�{��s����V_�&ާ��M{��δ����NZ��+Q0�/q�L��Ĵg/�ab&�n�[��}��а�$�#c�(Ǚ,�]�1f��y0^��8X�v��FK�[ "�p����ܷ�	����� w�eQSX��;���_V	�U㚝+4�V���P'�j҉��~�-����%H����3$ ��u+��w~?����ؒn9eN/O��ow���K�Ӣ�l�Xk{ykR�?�Fv�1�#g�	]0�o��#X�h�7)��e���B����OZv�R���3��jڝ��F#"K�ݐ��+�����,i��t�8��A��}�[� 1��Ѧ���hW�$"���:t��R�׈�x1�A��[=dc�m�e�Hm��<�|���O�a6�0���R/o�E7��Y��)+H�W%�K� �o@P� ��D�l�b�
�O��RZC��"e����v�,#�_�Z����,lc��Ip�3#PS���s{�؈T�?ǁ���+ �\c��㋺��y��7��Ǎr	8���]a@|��8���
}��	œ�54EäA4�]$\FG��'ר�ob�P��D�����_��)�QM�g`�W���ӛ����Øs\�cd�Z+�J�M��aA�M�D�\��xI0w'4�>E��/����`R��������?�])�>��L�`���ZK[_��=��@�*}�����Amb�Mw��54�-�%y9�
￯��n���
�\XY.g�6��r><u��ht0S�@39qPW=�]�n���ܡ�� �~Ɔ��0�ÊW���sR����Ԉ׷ޒ��6�<\�mi��O}T͹��h.#n?��dr��;r< <���f��4p�Y� pzcg��T%��Y��7W)�k{���F����o[3���1�ꕇ�;��@9u^���Q����+�C��K��ٟ�H���al���DLc鵟IEKe�^TSC3z�k
�d��o�	 vɖ��7^;Z2�o�_�?z����;jEx�>�fx��O�rYc�2����$�!�J���e-f���}_oS���"�~T�<[pE%�ş����V��h�F�q���;������KQ�����S�i�T�+����/�} ��ےd����u���W��;e�i��A(��)���!�7�*(��}���щ�� ��:!�`��I�PNU�f�6�	uf�
�?��Z�\Mz��~Y[����(�k�/:R6�Þ�*��_�7x���U��S���@\c�}ᄔ~`�e��b���K@b�j����;�]F�"F�j�m�30f!�Ն��i�ܘ{Π��6%���V5�a��	>$H�Ny�R�;��XwI��QW �3��jFB��2w���.2�������Iy5�z_T�.�F���pZ
����;��6�����Ӛ�W4%ءlV������"�{�i�j���E���>(�Z<�p�?"tg�����?G�a$&@@�T�q�̦���#c���?�3�H�C)m�ncirfty�?5������Z�"��>�1�9ֱ+~K�d�D�Ū�_�6��2;�1E��>3��-q�l�l��c���Ȍ�Cj!��<��\u�[��=�^s�%�A���mT�_M��rn���Y�>I��.3I��g�1խ=^0ˣ��p6���~�8Y0�#C��L{�U���V����_ަ�m�by����Ō��&〰"��F=�"1��k;��b��X�F��#�G����m���Y����(�r�57� ��İ�!ɵ�Wr	�A�|�j�Ĉ�?|0rQ7N�d�G� d��`�6�,;�nM}�X���]��*�:�ݼ��r2QJ�.��/|�X1%S=�]��yO��iG8��xG�f`7��P[о���f��� ���^�}���[]�ϛ}3+>Xj�^��or��@���g�.�=2��]�z�����'��v�M�-$54$Xϖm�Y..}qjyB�&� g�����)�O�e����Y䈻9L����K�[β�97�;%2X�A��@hq��(���ϕO
g����[��)���%Ģ=Q�o;HPr 1��V��9�G�8�
�*$P�*`��� d��?�2|���$��R�?�
K���f{���)�* Sg+◿�u^��z�Sr��9�G�aa+��r_�$� �_Wۜ}ad��>^���a!��LP�]��7D�F¾&�k�<ƥ�|���h�����R��Op)��,g��r�`\���̿���UA6�	�^ؚF��xy���c�A��IH
��%0�`vh58���˘y�����E[�;��jk<�ѨH��<�
xr����V�f�v�;ۅ�3o,O�ErT^*�%������h@9
�Lk�$���"�Rm6_�n�t�뉑�E�k�/��[!Ywj�_���}d��ÚU��f�����2�$��}x֚�����(j�����WԐ�'�F�J�Yi��\kX�;��'!�kԒy��n�cI�޺Ӎ��3`�w��|2N���0��y]���M�_x��Ijf!zN�(����h-e��-wU`�O���)ך�jN��ꚾ�.uM����5�����1�f�H��<0�%R�,�PrAO���#8���m{�PO��W�D���q�n�P�7�s�_��i�d����#�,�%Y�)Asz�e������ϣ�)�n��L���J���ד���3K�xSsۤ�9]/ �L�r"y8�J�������޿��Z#�A�3��&6��-�%9�5��A� �T��T�+@����#�D���>yZ��I�P)�M�G.�qo�s��w�4#U�=�:�xQ~�l� ���-�Q�jk�)n|~D�^��0^��f�NiǮ���K����qx�l:��+��T�&6�K��5����rqm�^H6E�& �t����z���i����}�ahd�@U�dC�n�c�̜�Ӕ�Oڒ~��H�" X�M��"m}sÔ���(z�[A��-��2y/�+ ؔZiY�C�`��Vƌd�(�ǵ�g �a�\sU+�v��'�]��
��f~ə>�J�!��q�pO_�x|w&�o�_�I��`X��
s��U�'����@�P�KYV+�u}��Պ�)�kG~U�V�<��r��d_3�v3�Iė�P��[�|h�$9G1�9�'.�D�pZ�U1c��K�c�I(�J"�Ô?wp��:U:���o�-e�Ϸ ��9v,g��Dg�'�5�{Gc���@����	cÎ�E�D��_��nYE ���Oݣ9�qX�E�D��\u�0�w�spR,y��<u�'�B�m��
�IG��jY���u��h]2�:.�_��w}%��#�"�ۺo~N����x�����������`EXZ�x�i������	%m�~sA��TT���L���[WR���%{�&r���
��[(���5��D.^���N�A��I���C"��L�X.������<�8��~�X�OS���~Ѐ��݊)~U��_>�i��r� 3��d��bS	¬0����A�E>8"�Ozun�,F�"�t�t���`�s��)��8��u@l�o0�����L�A��5�<�F�z��F!G�&�( ����:a��-	��:TO\Q���y����J�0���"��oT9�/=>Sgi@���A
���%b�m�!�1c�Џ��(��QY����M��P(ϼ5��XB8=���$�'qR�8�8H��U�J:�1��L��A*����:rg�^��ag�ں,NP�����?_��2�ҧrD􎷞]t���������H��2�Oյ�m�q��2�l��!��/�f?
^o���8�A8�.�@~C���8��hC���p""-��^a���B�Y�M�̊�{�v�1o�d���֝��P�<�TWCU w��~QW����L'"�o�1�͗�������U� �"Է��e�J�K�]HYR��qAcV9n�O����ٛ���N8g>ZvQ�Xc��30�.ӽ��L�%�be���;�����~�J2�o����B���E���b�J��^9M��>�]�Kz��@T�<�B��!!jf<p�s`�YY�}����=�(���/lDFO��������ED�!�Q���N��PYώBg�]�k��J:�ϻ�*s��X8�.���4�[�lr.Ŭ�'����f�Ƈސ�s8��\��TX�	g�<��Wg|Ȗ~J���`r��~n����h�-QΩ�))C��ocv���YQ���e�z���η����]T(�0N�!)�L)�����<��!er{F�$�9�b>э�XJ��t�c~I��B���ӛ�S=� �x�0v6�1��f����&��8���z��:��TG�a��**w�CEx�@V;G���	�<6۶�L�@�O�"��˹y�(Z��{&x��﬩w:�+	�#�wt\3Z�#gb���������ԪT&	�ᓣS�h+əsR��z��Sa��)��Y~��Q���z��VIA�Z��zc5��f�\��\5D��`{퐧;�w��Ma�?#[͍��lV|A� 1?S�� M�|���E����d8ul-uo5Bˡ	i;QGIW���c��\�ӯU��@�H�ȷ��T�r������g�Ձv��ԣ���cT��5#��$��^�?��%ն���HmE���5�:c��XFw��3��NM�z{B��̥Eqz�k�Q��
V̐5��:�Cꍪ�-���L�e�i�	k΋-��b���Z!�V����jڵ}0Oi�5)p�.#X��o���C�
�)���W��P�/�S�Ͱ5���x�7$�?>���l��e*Ʒ�6'�ؗ+��ؗcr�C�ۢ��#�=�OZd)��{r�w�i�W�۴�z�W��@�E���.�|��TV��	@&ɻ>����>e����Ǐ�N�����؅Xq��!���I��p��� �q;X�M!5����>�k]��6�ΐJ��A��z�QT02ha�-t(�k���L�����ݮ���IJ�2�IW�qr����STd\Bɷ����0��R�N��ʽ�_YA�(Wd@�dPe�q�zU��T�Z�� c@��CwmJC}t�>�DC�N8�fyތ��I��UH{��A ����mF�L�ZX��=ܪ�]}�.��d(1�kP�EK��w�\�}n�H/C6�>�{,��7�T������>ʮ�]�U�xP�]ҏ��O��kc�$w������_p61�]���Q�z�(qX��hTK���mMjy<�O1���H+t��ǔ 䐒�˴� +��� � �=���8��a8nKl���{��n�A8:���wq�̍��X����2	bx������9��$A���58��F�~��m���!�k��h"X���	��t�u�������������D���.`��s���Y~�����Լ��N%�S��ԁ�Q�d�eh��B'�jp�X�%���͐�|�2��@xb�֚���� ��#�s�0���v�D���BY ��3��pe��cQ{�j��Ǡ#xb���>���2��ާ�1ҏ�J i �*� �E)^&�t߿l���#?��a���F��	$�����?T�YV0XX�"�:8g*��Xjo��h� ��r�ۈǤc7�E?U�ow]�;U��i���O'C�=�_:�XE�][DK2K}��c"tĴ	{M]O�v\�L�ƨ�`���0��Wۈ��3��Y�a;�j~�'M��?-#��Ү�&<,��mk��ݎzr�!I�4��Gl�M�@P�оn0��%[+�W�Q�Ԍx��ھvA�
I��o���!�5��z�%��P<��SɌ�)3��T�@w���R ����6�x��5�ٙ�sn�cToS��0�j�y�`pѾy���JO�?4�by>��ul��!�>�Ƞ㩌�oP2��O���qwf�(�ҖQhT�n�x=���?�`2*;�,Hz�&�`�������;9��+�9!�BiK+�u�D���=�V�^z�2���;��բ�Ü�~F�:_�B pɬ$D�!g����ۙ���c\�L�DI���SEU�X�#<Vk4�`���AF�>�㺫M� ��L<�Էf��Y�:�&�X�d�Utt��V�`	/c�M�+�豷U�ؼdSO�؁����hC��wRLL<�D��=d���iђ�T���n�7���2��"&F�`?���t@t^�#��f�GKD^`#�J�K�s_��谾��g�"d�]��4��E����$�=�Mul�	�찗5!���~ŧ���`�4�{�!G���"��;��x0�K��vR)q�jT��rl!���&������|���@%d��P �; ���&lw�fU)H��X;�be�˜vah����<�~��	��h��n[RWx�����?�1������w�6d�0A7���
:0t°�h���*��v�ě��*�ѣ�J)5P�]����XϏl!���顪\�+d�M��(Nؽj�� �Z���
	��p�[��Hl��}��|B��{����I�x��q<�D���IZ.�{�Tfn�w��N�H?��@g���kn_�/t��: :���#qґi.я=/��=m����^F�ß��"g,G�.��\;�{b�4��kb����A�.��W&j Z~ _a���:��/߃s�vtAN zU�7$+��^y�D$Vn���U �a�:���O+C����� 4�%����a�T���>2E�`�E�'���𛚩�z�H�T���Ӧ�_.m�'��m�~��eˢ���^��`�H5�"e�ڇ�P���g����U=�⪌ZˡjSp���P�,Y�N w��&����rj�,D�$X�=FO���v"�<Hi|�M�A��p%���G{i8"�c,�a7�\��F��b���a�ay���Xt}KP�b�zM���
���mȍ���C&���W�(���Kkȯ
Irl-��ű�i��f�����B�~"����|L<��k�D�y��B�!i�W~dߛ
0P��m��M�FLڀ��>�X|T1P�S�C������s`�����획��E�=�.�����Y��K�T��\����g∪� 3YU�Wm����i�r�nb�É�Ϟ��mm�t���_-�\��t݅�y�B(ROn;H*��� �ԴD�U��U���D��&1PR��G���%�ji��-	�⚛^z��i��m�x#-�1�UǲF���f�s�(lAf�vA�K������H*�#US���̾ΌX����j�Sn2��8M�)'c��UX��I���-�5����:bϮ�ԑ�n������2���L��8�7\�Yp��$��m�s
��G�#�d������U��7LL��٨�9�k=S�I�K�C�6�x��j?�(��e��P�BET� Z��t�=T��K*�t���g5m�~Q`�"�8�/x�ȹ�]�c�w�R�t`�3���+�|��S�,lG�^'�&����/��l�X�S7yϵ*�8�Dz�@�N��f�!���Jh#���5hJ;��ɶU{�<8z���S�S��:� wk���Q>$9���9���D�=6T$�GQ���H\��f7�����&�'��{��C���DPt��X3rH��5�i�D�� ��i��Ӑ![d~��蒪Q$�Yg(=�Q�[���p��t�Xa!E�J�W��|�����[A��h��o!�b�c.Y��y��d��&���F_~sBRG�n �d6޳�uG"I��Lq�:
�P	�V��l��!��ܬ�VmB��L�6)��
�^5�S?�p�ӏs�)����V��E7�.��Ͷ
M�~��(������$#E	T7��"QN�H#ٝ.��������+t.y�貆[)X�R��P'�4��&4���:���$
y"��3�~Џ'�r	5� DzR,��`�����Wp>�6�2Bf�]�x%��WT�� U�΁1c�5�����}������,q����{/Ȅ3j��t
�E�-S�=�R`�(r�K�Kc;���(tK���m�?��+?t��V���}�MR������?�K�F���B&���7'������aOt�ފ���
�Y�ed5[�1r�p����u�< �+��ȫ��q�/Bh*���h��=oG.���pi˳�6hA�/"����"2�l�\��2�.���P��]eUX�J-v6T4�"A��y�`Z�<N�}�*?j�^��&�N��Ǒe+��=�(u�ðy_=oC�yuRу�[�4������_/��y��t��i��,%�B���� �A��\��� �Q�����(�9�Ѓ�bS�A�8���EK�DLfB����*T��K��g=��hT���'�F��R3����_�iѶ�]`ɼzpL��bm�)jqdCU��yV�y������]�/�㘛ى=�t�F 7Ϻ��8��9{.P��+�[u5��!�S��-qDX#��B���y�<��oXǷ�	$�Q:j�3P*w���f9p����M�"I�JU�#��x.-qM��A�u~�ү������-����g�z�Y����Ʒ�w;u��_���iB��蓡����z^iK���RG�E��}$V�r��ݝ����P(Ć���Ō�w8��	��P3�f��j]g���q�>���v	x`VF�`@��M@�5��i�Ω����l�c�\xe��#`w0.�ɕ�P�a�8°�%7�����f��)��<p����V�*T��h�nϸ�ԻguJ ���(9����[+$}p��$鯒�3|��^����*�
颞BcV��P��I�*�L��"����T|�a��M��ۍL�\ٛ�09Q��i�� ����~<��e��EJ��Vcq�S����)�	�!>�]|mj�R��s*$;�խ�Ӄ7���R�އ���1�e0A��ˍҨ����!��Kϫ��$�?�R�����-t�n��=R��(�L������N���<j�ޒ%�1uYύz�%IH�i4)��]���)��Y�oL�=�u��Mȶ�J� I}{���T�ٻ���X�C��m�ʉ+�`��C��qr)�YW��,�=��56� �J�c3I��VakX�S0��D�<�Bl�c� ��?nۘk��"|@��q��V���Ʃ8-��a�Y��0ŐgM��/�?��-%��&�傌j�j`3w(���Ý#��>�����	�[p��f�����PmNIJ�Q̫O��u[���h�v�Io�)��V�c�ȱ��p�O�� ��xa���cz�nE������UϚ`�"�H�X��w�'_�|�k	�a7�ݾb���P���թ�SS��ˡoVr3P�M1%�B?%%
Z��>�}��}|M�O��֗9�ڔ*�2���HAXd�������t�d�W�F)31fdDƥA�o��±P/��'M����5-Q��q���5����o��2*�ܛTŅt���+�&�]��y�k�A���!��^>�즔��[-�%��
��!̰��X�Cr�<�0���_P\��[t@�;�M��و0?�C]ymN^#ҜjA0�Bq�}��Kr�� Nybi��Vjp����uK��iT�̓��k�����;�!}X�c����5)�6�Շ|3|;��!��c<.��S��dW����~�T�b,���hW:��i�$k�˸�ÿ`�y9�V�u�)Æ��Q�y���������<�6�r�%�35�A,����u�!tX{`�b1��[w��_�3����aH�5kP�Г��L��hѪ?�I�]�1�u�Ӣ��M�|o�a�-.s��.��<T������ye�PJ���0Zژ��<���/���&�}ej�K͵D���
q�UY�}z��A��X���������]Isv�SN�H2�,���dP�$Mj9H!@U)	_�^V��1dU���jSi�[��X�p����:s���j�#q�
��^�q�`�$�j�ٰ�*g����V4���1����ɐ���7����@/E�����ލ��܎�-x��O��U~�![���u���>�a}'|;�fC����BT$D�<=UB�����+Xn�����)��� ��Ʉ��� ���U߫����@�I�WB�|������������?Kf��6l(w{w'3��~�M���C�b�n��OFV�a͸��"�%a:ND��b���b�]��׫�4�v���H��P�	�e�z�� �s2�F����d8��7��ƅ&�v��@J����w�"C�C�rد�N����hT�D���¨� �4�=��B�$tQp�=��˗30ܬ�W����4y�UHL}7�V�x��~|�&�w���*���.Q�)�u]�P_ ��Ǧ���	B�b�CL�2az�k�����u�z<{�'Z��ȏ詣���	}K�8 �,_v����dݕG�t���x�R8a�[ֽ`���pK	Ikq����3@��wA;S�_X�;����b�*5�KVgܡǑ�\9��#,]�`W~�,Q���/l��po�=��3�:���U�&�)���a;��J��]�prE0JR�$��\�i��?��4)o��A�,������v*�vk�܏z,���&?�t�Bw"�dl��#��y�}f��،98~�7�I]�d�����F��QG�E�0Nua?[�0x2��:-"��l��X����h��O��j�H�1$:���K	)��mv&���z_�B�Ar�]g�<����BwR�l>;�x�q�`����L�Ԝ6��
)�"0�V.�ڞi?2�SHntV<���г�z�0�F��7��sP�t�k�����m��o$Y�(I����{�7����n���i�����X�hU�@R��J���uL�r�[{IX���� �i�O���� �bB���C����W�����\7���WBVI5	��0%yV
��� ���x=��'����<\��Z� �ZH�s�n��܃������Ʒ�p7f)�2W�v}0ƈ!/��$��8%���-xJ�H�FB��^�	�U��~9K$]?O�6� E�r�"�v�`�حa
��5A��L�;� 5�s�.gK�_ʻ��E}<�y���
l��,���a$�0g;%}�)���U��Q�2�(h�	�dc�����B(�gN;�&'1�hX"Tn�y�|()A:8��+-�	\�ǭ8H1P�"2HL��b�4m#���=�	Av(L8��-��}�v�k?qPT��k=�U�1���.~yF`���)��IUG������vZ<��ݤ�����C�������4���a��4ρ��Bw�qˮ�4Ǵ�#Z�|����۹�d�ĝ�d�L'�No��U�R9��ab�f�,�Yf�t3S�\R�K4��ptI�>�1��ޔUX���#�Y7jQ��Y	�t�ݸ_��AvBs@��	�zV�b4RK.�`�ro�f/�����Y�%��6NIU��,�D����KO�"X���Ϛ;7Ց"�~���ŕ����A"ݔ����V��Z��~g�#�v�,�Ц���P��~/����E�~�%�������q^���.ii�6]�b�u�|��?��n�o���7]�4l���QB������[Ħ�I[�zm��c\g�f0�ol�����{�zr��l��\𡩡�z�W[_�q\�����7���n�b^Iph'�㿴�1PK����N��	�Oߣ^��l�r$=Ts���h�g���@ck�Z�Sn$|v_~���3���'�z���_�8A'��m�R��n�� ��B���ZZ�xܠz^��t�(,a�]����4�J^���Awoò�#�R�Q㓈�;�Y��i�V�u�3Q=�%������w�h�߃9 ����Y������9�]*��4���!W)�c�SOg77����m�