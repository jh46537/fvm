��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(|����	t!�ۿp:>�"������P��)؉+��}�4+�}�0������� wV�B��R8��$�+�N?$��e���2"���l�0T�(j�^�*��#	3�
�e�r���t� z����2��=n���Z�Q��'y�������s��LZE�,�&����5��m��_���Hd�S��-l�<�	Ze�J���ȟ|	痶��;��$��zl$���|Kj�q�?�y�t�;�%�����`��&M�S ����+��!��$�q�����2)�S�Gc�c&Z�ᮝ�b�ZO�m�N�+ш�Q=�e�.�SO�!�S[·4��X�(u�',��O����潻o8(�jHHl*xG]v:�?$?c�`ظ�:��u���8�1
Zb/��AL{�R����8%Y �jO9���0���"}pm||��b���"�3T�oa�wQo�N�;�S5��i}�n����{|䞜r ��W���w�*jSVK���g3
dG�r���99���r��@QNWk'%B
D<6+������D}�+��a����E��-3d&�Z��^>o�h�3U�5��oQ��-��A�m8�S �Y{㔪�R�/��u&x��;m+Mp�����������٠�ZQ�#�7%����L&ʨ	E��<�+��k���J~��CEm6i��������Y�<�;����CtW1Elx9T�)b{�3��:mNa�ֵ_]��
�fǇ�� 	�jvW��D�����#�u�i ���tۍC�$�����g�g$wM+��Z��ܯp	�L]�qj�f�m)S���%0'�~+WeZ	Es�Dw�^��Ԏ��/��H���x� ����`L#w�Md�>��\�5K�����ݷ�Ny�9&q�4�V��㔚Q�T�ȴ��I���u�?6��F�şcDN�nQ�I��N!���i
��U�ԯ����h�%
�Q����t-��R��AZ��@�"V��"*]d��$󖓟~�5�zRE�&PPՒ�xzX'" �>����I����->6*��Fj�MX�һx�S��	�Ŧ�,�峑�\6��.Oa`� ���;SΟjM>���-�No ����]v�����ܐ�}����A�8t���������r��H��m�.ͧ<���E�=95�&��r9�)�F||���`p��!��ۘԛk&�%Kx�j2-`{!�IU��MR�q�o��(
7b$i�~�ڠh�7�}��p}�����y���m���3ȕ2�'�q��wb�q���oɶ_�n03�{����S��=�k��kO/	P�X�E{���$��Rh���h�Z�ul���*-�Vqzr҄$�]�ly��Ĥ5�;i��)n�5F�2��M�cq���9"�,s�ԭ�ܜ�����Ί����	�:-�<�N0��̷��ͧǏ���g�v�)֙RnA��tҒ	=k}���h3egѷ1/
??�5}���sOU���LR�Q+���f�'��ǹ^q��;m�t��m��\��U�dT,���CՆ$��C�j?L$A4-)��ۆ+��T�zr��?�U D`�ڛb94]����iv�|�Zг�&ri��g;<�L��)�s@1e'���e��'3a��V�� �b��BU��_(�=s}��(�H �8�)'��%P�UwHRp��$����P��D�1%��L��/�\(&��F!�,�aC'��1P�����XR�eQp���x�Y0*�	b!~�w�CR%d%�(�W�B�������[&��ʶ���Sw�S
��6���cӱ]1]���E}41'�����ewwںŕ]�E�8٪��-��ܡ��13
j�R��:CЩ��Z�y����Bd���h/_��D����G�w�I̖���7��FvKSj��x�"��*2otH%�RA Vx��p-�X���`�X��xt3W�ώ�/Oľai"uq����Ҷ=�'8n��;u
X��6�46o�A*s�Y�%�i��HJ�z��=/7�QJ�%�+X���mh{������rP���HSC�/��E�-8�p��<	NO!O
�J�+�9Ω�ho�ll�t��������Q�4h{R�������m����8wKȁ��գ��P�JL��G7��L��VɾG�apo�s�A�B�\��nw��������[k�����k��
P�*4������������yIc�z����qN�8�oB�6����{��U
\a ���g�����t"�T�-m�A/�#d��;E�f?�9n��m����q�񻪅��pR��̮Wv|H��8���R:�B����ԓ8��=��
�C�i��z��{�[.{�ڑg��\�`���%���66�_�S�K�c��p�5רU{��2�wmQg���I7�kǺ��
�s:jt��b��n{�����}�¶�JlG�m��R� ZcT�[������~y�Λ��.+��J�B������?��<G�@ˆM�@yL���Z8,���=�kd�a�E$��~��_习Z���7�
O�O������&#�_=�܉�{j��y�m���3�J�Uo���l�G�\�-�O�Ù��e��"+��闡�_(�S�%��8��K���y�ȷ�w+��m'4��*��r��v���)m�]�t/�9ܿ8��4'���� ���˦j�HK�$R�K��n���8Y2+҂�"(��ٵbD�e���h�F~uN��w`j�ze�8.�-%���o�T��-P���
Πk1�+2z�_D��o�K�8��,ƕy�+�_���H�P��}}5��{�c�9*o���Gݛ M����)j����4��?8��4����A���(�g�����ǹ$@�+�^y |���i���؍��mP�e��SR��>1Jz9��i(�3-��G�3���;-��:�g_G�4��Ȝ8�)>��`ݜ��`p�u�/XHq���3�sV�Ȉy�*ۋ�0m��"��#��tF͕�O9�2y���ݼ�"��>0��`��O��0����̈�{�eg'��̹�8'mEE�޳��O$�5���3%��y6�E��w��o5��Oe]��rU�Z�RPb�0��T.u9��5�.mB��S�P��N�ͥ�Y ���g�⸃����
�ce��M 43�Q)-�T m&��Ĕ5N/�$�оXx�&�����yp�|�)t�6Ku�(�/,�MM
`���HŌ�=%[Qh[�?�"L�BT7���O�N&��l&��! �pA�wE���h�.�o�qt�Kg��<������~.�3Ҡ�Z������hk���l�9���pE3��7x:LPm��ԄB7�=8�)�x������f��8Oe3����ӷZ�!���Ot%4�����쯭0�u:�Ug�5�"�J�L��6��;#T�]٬eϰ�����R1]��"# �@��uj�
��?�pE�_�>H��)��w�m�R�?�Ɂb8*��zq�����eN10Y?�+��b���G��sh7���D{���Y;����L����%YCEh� U���
���o�l�mZ5<�LLq��w���)�S;	�}��4]�U(ٞ�͈	���L�u۹<�k�\p�!�*YI��Ȣr)���ߏ9��D��������(A_���-qYP>(LjP�`l�ݷ��s��T��?�d}��c'bF����!�ɧ��t&J*#��5;��2/A`}�vRWFO���i-f��p���w4�����+�+[�����F(�k�)@��$��g����#s2���q	*(.�n-x���͐��;|���k5}󧢽���`���6�K���%;!5��~�KU,�jp��%w�H�V����� sMC��\�f�q�C�p����ҝr�F��d�e�1[����?��CyP�E�B�-:�ڷ�(f���8t	����k�^R�9���]ED�LM����װ���\�\q@�Jwl&��W!a���&-uD�~��0É+�M�9����mBĺ�6 �O�_Vh����Y9j��E���1��Nn��Mg:B�f�4�$׭�,�N#��c��?�����Bm�}( k��=�/��8;�rO{�5�Ӗ��%PR� ��#�����7^$嚛���&Qc�&H�-���h�d���
kn����J��:Ю�����4���V�goڹE����Q���A�1d�����Ӻ5���P�1��0Iv��֐�>}I��u6����e�i>��O�2V
������P�N�/���� ?~�.�_��������F}����f��);4I`����������c.�O,����S�BP��^:�LA����-��{�i`��gez���)��yo�~��p;�Ȥ%T�Za��+�м���+~e|a�:�t���bk:����H�	���)�C5.�p��߿x8�����W|�q���wq.�Ͱ]Q��-�U��ҝ��y`c�y����+|6U�K�Y�x��*,5�I�|d�_;Ԡ���xd<n�:�P�[�˯_�[��w���;X���hz� �?��O!�}��`�`�.�6^��.�>��­������zq�í��3�xK��G�S�ѵ�Xn�Z���)�H���;_E&�H�p�~>N>�f��@5�!�$��V)O܎�o8��:�K"���T�ʹ u�+�z�襚����C&�^W����<��A�ی�����4XBAKD1L���t�+?�"�H�]�:���)����ygI�'�[���L_@`[����;���(�#3%!?��vH.�������<�5��s�D�p�Qp]������9��H��nPS�f�HP"}�ɅNL��8̂=}8�n��NP$�Wˢ}S04��1�M�r��5��G��������ȋ��K0�2.��"X�%#��s�}t����?�'U�m=��� x�U�0��}?�נ���XU�'y�����?��
����N��h�p���� �.cQ��X�9��X\}��RM��%���d�7�ٯ�r)��8�me�(����s�$����o8��n��� ���sw��[�q� !:��'�'UߢN�ՊJ���b��8"�A��D��H��cI�bʭ�ӑ��2��M��b�ue2`%�,����[�,uSE~5~$(P8�,!��5>�&2�4 ��}\��4$�K�"�#�XC��g�|}�XC�{�)�A#�ϋ�e�lޛ���Զ�|$P�2߾@�+	���f�5�vr�n�����{m�3�gF�n^�(g�Au��c�,�d�ϐ��v���X :ܐٰ�T�s	Kn>�ഫ�c��^�P (剰��]T�Y�ÂY ,�iQ�l�����6_r�y������lh����p�D.؊z-�C���r�z'��C�|\yx9�sq���cx�:J�=��U��_-�""pB�yb�6$$s腕�	�������RB,)��f�l9~�@,\��	F�-ro��p'O�\s�Nq�`������C'�5��zG��X��L1�U�6����m�g���Ɨ�ڑ��ku���h>g�𨆻�4<�`;|,vZ�j�p.0Ic5lc4+&�@��m�
�>���WvP�t�HN�`�1LFϪ���u&(��Q����	:��
ɺ���
�A,��W�F>^�E`���E!K�? u�&$��O���0γ�j/+w���d�{��z�ä�{䨠����;�����t1�ʡ*��6
����~XPp�fe�Xŭ��;}����]w
�����}[�y���������,@��ƫU,3�O���}����>���O��ݿ}TF���81��Dg��DW_m�´*��p�]R�P�������B�J���,�9bХ��T�&�q!H.��9��4V�6��|�[�
�2�����B5K����ȱ��������n}҈���6��;�$ex&�;��nڽH��=����x��_cy��ٓ�U�$�k��a�p����lY]�" <�$���Glb�f�@��<蘛��n[�7����9�y��V/��w]f��T]�7#��%	�Ɏ>yݭ�_a!Dz|�Y��f�u�%�5]�*�j8f��In6*5�Z&Ŵ*QXv$�ղtq����v�u|�4�&՜�*��_���|Ӟ��^�\�Lr��:6J�C;��b�M��K���b�B�a%5ɳ�*M�"�8+�+�k!�~��%�H; -���� R&�l��'[��
� �;'=͐�<��f�'!���q5�5cN@C|��Y���2�%.�a���gך{�2#f�������K�eK��K9k�9�����+)5ᯏ�ː��g�F�Ad������X �hO��9\�\����Z�7��=c��aA�6�
-�������	��M-�3��O��oIFoA���w�~��TkT���ɳN_������/M��}��v&$,�-���N�lf )�
i��y"���s��v��J$�|�R�ø�@m��"���TE�����7�� �>	��(\u�l���A�h�kA{��j �P�ˢ�����3��*EM�}� �Ll�KӽY9��A���,��������{#-l)�,��1USi��Q��e�2�M��,%Ҁ-��Û�ܧ�� էL��Y� �iW�M�w���� X>�ޡ^D�e~M�am�b6��e�MTA�*C:Q�~��/?^gP.=V��Ln��b�B<�!�A��L�[��-�fҐ�Yj�`D�iu?\�E�����ѝq̃ i.jQ�]&���4i��5*�3\�,&[.+r��Ԝ;l��bg�5��}6k/y�i7��pI��!�q�)�8�LpK�z(6T���^�8�l1g��Hp�q��0=�����X3��������E� ����|�Z�K�IX��jf��q�L��_����=�1K݃q��L�y�c�D�pJ&I_uI���A�n#�p.5�n��3�Ħ�eY賨�H�?Ij�ئ�H��^����i;�]�j���Vu�u�5��(��盰P"���a�i��v�j�0����q!L��L(�z�H8!d�U�a[0} �X�eӨ�f?4�k�*��i�������J3���`�o���*���q�zta)?�a2S=d<���t�t�`j-=����:���_����*����J����2料��g�bjTW~�M��;P~~̻`��.�?c�����Q�dp�$	Hc���?#@͟����ph��H$+��9�id]������j�7��0���:H/qː�}�5^���_Wj	��T]H1�<��8��"��g���P$����6JX5��72)	���VMM���z�^����<iJ��<Q��E�� Z9��1E]�;n�Sx�tS��gdiĀwyK^�R�h�O������᛼�΄Ea��Lq`��,V�푰>��DY��X5>X�#�	�I\� 8�H�Ec�'�iĜmK��xf1zEn��v���ce*/MO��t���J���;�z�����t�@�h�|q�E��&����g.~5�l�` N
���،���ج�k�,
��;�� �@'�<��kqH���Q���-_ȞW���_Z:"%"��M�[����ϞG�#�?��N�P>Y��Ǣ炊����֌�h u���7O�-��V����;�U�9$4���U���u�ź��%t(d�4��y	�2�!;[GF��%� }�$�o��gw8�x��}~p�X����%��p?��즪it�RI�=����+�uZF��W��߂@��17Sc�?*=;S�@~��BF��f4~�ل���bT`�D>h�2�]�:��z���Y�w�~�bM��&Wm��'n�Ӆ�ٱ��L��b '�>C�;�tM8��\�e�?��ϒ�v��������e+ދ0(6����焣%E�c�x~痛 |~1���nPa	n�6c!ۍ���`�d=����@�&���T��5��F�9������Q�fNI�!�57T_;��G�!� � ZN5�����@t	4�� ����ӹYțΚq�eL���
E?�"ي��H�2���d��聐�{��}?�4���bg^�d9"lz��b�����<�a��$��9�>�_O��c �	O�i6��2J��o"��f��&|~��:΀t�O��W��1]}SM�yy��f���l�%"5vbkm$�!�~�f����.}]�.�E�� T� 7	w��NR�`�Ds����6��St��}��D*���^��豞����_��uU�RP�^��K�r��r6w"�*�~4��p'��*���jM ��
�q*��SȠ��\!ZM"h��+i��L\�A�$�|�2E�;����̀��5oԭ�`mS��vaw�ƭz�d�xN���z~/<���!����44���)��mN}_(n��-��-�����nyqKK�KS�ͅ�'�F�UM�e��۱wT�1����������a���,	r��]FA^�w;�(hLG�����D�rV�~�vN��P4i��2ٛ+vbx��(	3��iޭ���H|�ȉ�\�"$�n���ȿ�0���Z͎-����D��nʁWҔE�??��m�Z�Z���bЖ�I�N �؆�ߒ�R��0�	ܦNDј����i�>�����R���o��v�NַJ
sr�z�A~�d��%��Ύ��VI4���A�������}�Ϋ��y�&�c?I�:KV\�	n
��q�H�u3�:��4P�lFz�&�o���k���bD�Zb�T�9i�����M�Z�f���q� ��.�d%Ϙ"�9�tN��eZħ�dZ�M�I�23�:O��<�v̹����FxexX?�H��ڑV��&�Ɗ�w��FgX��S�v:0e��zV�5$`��ό�^���Ex��=-��%���,GB攞	G��M15VM�m=��cƽ$J�u�}�C[k��#q�z8�Q���US�-ژ�� <��C��0p
ܕ<���A�;�w`
#[�t�w��������Ce�F9�ӿ.����vЁ8O^��=�����Oo�3�˫&Y�ض�u�uL�H<�f���S:���>|`�[죃N��`�s�iƦw�
K2�f �jx�q�� /X�#>y����̞e�#�[A�U��}_?T�D�e�>�d7�#��Eod
d����-�i`~��z ��K7��W�"��-�b��O�N:�G�P�h���q�#U�ui�s�^Ʀ� -@��ؠ��I���y�t[��ʆ�Y��nvj*�/d���y+^��f��6����hN�����_�ǧ�TI��?e�][$� �b��9�*�����QQ����q2$�H�!m�K?];TUp���m�M�}���p����cz�P7��ӯpCA�C�������Ͳ�h½�P�_���q.G^N���:��Ș꾼��$�Q`dֱz2��F"ᙨ��D�gy.kD���m�c]p�Yqk���R�g�K����WzCT�E��?p^q;4�}�\�H��zg��r�SM���X%�HL�!٤��;4,���*^(1- (Y׺t$S�dI�n��%1 2C|T�B{\�O���F4��!�-�������ݒ�+9�괰'�7c;���^{^��i����~����+)z2L��Ì-�O��iW]O3l�=������܎�7�R�A� C��:�ݔ!�qn�9(;]���Mט��]�X	�,:�V0�[+�)}��ؠ��T�w��X�����t'�#�Zq���P :DgJ�N�[�����k Rj"�u��X�5�(:H0v��+[[o�\��\ɓ-7jI*���8e�ycQ��4�%+2$��m	�W�����֋��\�ZY�}���p0[��3�=���&��͔5M^�i:�۬�j��P����
uS���(�w�����e�1`t��rp�ꨒ5����6a�~oO_�C�-��
��#���g�������e��G��`�F�,2r¸����rj��n�o:�@g�Lj�mˤ\���kK܋C��Qz�:���] �D�~N�+&6�xN�c��73z%�����ePX:�=���]��	X�EϚ<Д��$���JI���;�6�
B
�������*�K:��_j�˱�����1D�Q��&+W�a�i%sZ�g�	O��k51ʎ9"�bf��Ѳ��9������=��_�#6�Z\*�s�N�_C03�(�K���EA�O�/�J*�$3��uDUzI�6:,��ņ~��w,T�Ѽ�9EOtv_2���P�e�"�:���>�x��8,C4�5���E���1���QO{��H������!��8G�[>�gJ�X�!�UEBi��O�*ЀMG�G�Z�e=��/-�^�a�������Sa�� ��Ɯ���s� 헟੪;-�!
��T�� �A���+(�%U�^�� ^p_&5��K�}s���a![
@�"��˄�X=і�$�i(�0;Jp��^$_�)�ĩ��g��ܰ���à��"��@�t�\'����h'�vl����Rs�>���Ҫ��	Ŧ3���#47��Kg���ڪ��O����ӽ{�kT8
��c�P���C�t�㜥P�l�$k<uf��B!�C`�A�e'�0{ޑ��6�����Jh1�RoU	�B�G�D�c����ȉK�of;��D6��W�-�3W��!��-7I�k���5��e��2~�ܷ�'(�JY�F�|'h,���(=ƶ���&��o��h�A��F������,R �|x�^'E��+�?HK�ZD]�����Io�R���\��r��m,|�'M�>�����x�D�ܜ4ϚZe��h���DLf�o���v���a`DcƐ��}|����|â�
���+��(���vn|�f�
�@��q`����9��0B�(�Q���+�+�>���a3Y�&��ƚ���jߴ@���O$��C��q"~�I��cff��9;�i��Jn����Hiq�B�����qN.���ݨD�(W@;�ۧ���Rݶv�3j�0M�����v����^��򽩇��gIu���E �aá���\0i�T ^hy���
K�ؚ�,Y��|��L@�ݻ�-4i�]�����]
��w�!L]��Bd���)�a�<Փ[��C�k�,��%|�L��	}QM#�aв&��@�To\t�΂Fw���F@bc�_�<��o��|\�л��_�n�1�|�*��:)=�����4W�V��v�Rb�B=� �7
x�ݷ�[ɥ��w��4M������g���ލ��:�u�l�M���==�eH���`��n��q CLY��u��9�g�\��al�V�G��Q}��E�>���.��'}.��e�P���)&����?q$2��O5�Yh*�TȾ�jIq|��r;��� ��zN6rV�+�p�#�
�١���Q���2��Ʉz���m���]�\����m��X'))E�g�6a}K�R< ��[���Pis6>�jZ����$0Z�w[��4C�9,���!@�xϱ�*�.k���-^9SL�����<�K�2�ʲ�t����hV�O�)�B�I�b�$��9�O�XG"`@�W`�K<[I`�Z�~�t��l΀{2�S�v�C��	��dt,*V
��F��T�m+e;@��q,K�SC@�R�knY����,�Q�*ڤxޝq�wɐqG�9,����t��G%��?`�@�ڭM��V\��y�ֶ�C�ۗ½�_�L �s������)֭����8�(�lMf[��SWsǾ�Ú��bw��EF��	��d>N���P�+OH?�и+�p��yW}DtzC�ţ
 �0,�Y{<��	�mp��BOg��Aӈ썒x���z���sh��d��-D��R;��,�y�5ó�O��?5�5��M�OR&P$J� ��ns���7�0��o����؅�_.c?>"�ŠVn��'�a7Xy�'����	oЮs__Q�`ͭ�Kޠ������#*�Y!E��K���ܕR"�E�����a�i�i/��!oLx���zW��C����EQ2�l<#�mz�'�xb�n�	���>��q�ha(���R�Q~�L������0�#�Q`�H�]0� ��֎�z�m��B��1uӶ��W43�:��{|Q�,%��Df�����Q�rK�ng�sBv>x�"�6Rjv�'h?B�-ڛ��.�C}�o-U�
&&&����r���|�3M�n���3�=�[������8��1,��7e�ЕT��[�Z�Ô�m&`��,�37f��'��
:a�L��[fZ��%��)`w�:�;�?W��;�֊����lo��炠J��*�z	8G��%o{�v��w5If@/៫ 7�O�S�������D����aM�y]�a���: �������l)���+����0��,��]�N9�9��:	�\���U����ɡ\������ ��]�pYPsP�]sv�g�0�S8k�7L��"W��&��n��;N��$�G\0H�r܃E��K�Dp3P/W� >\�$���� ��$`�����}�f��1T�Xm�.!d��%r�g�]�`�f�,��m5|P�<bH�nIi����4���!��a�Y7`y5�ZlV��y.;gq�6")���E��7\�Z!N��d�2��N8�v�&q�F)~KQ_��:��E��e{}�=D�0��#�M��Eb�Y�G���� ?���!��N�+r5D"�.�S���QՏ����W�<���V9z�ۖ��z��B !C��!W�X]���D��{�����Cz��Ξ�&�,d)4z����e%թt ���u��>Y���b��u]p!-�(c,c�z�A�C/�Ơ�(()֥E�dR�AR�M=�X��&v�����ݐ�C#_�J�k����.���ts��<W���f[킳����ު�����ԯ�X��^�i�鉰kH��=��#��f@ {krڼn�`���No y�!���l�K"��&9�9�^�����c�Y�=��捹&�P�[�k�=ӳ�vB�u�����s���Z@';����w��,�S�/���~"�}v�ݸ?��=L!+�-����V���qz�bB箊G�������B��|I*��Jh��Y�+�d
��84�Mk�M<@xlXdG��a�p~�D��3�c����+dv�K�IaBt�����su�n�x��^�o"���6�[�����؊�Q��͕!v٥L���sg��it{��>B k��6���i,�������U����ɻs ����lU��YŢ�ҼDy@PC5&=4�@�Y��8��=�ެ�Z�\��@As���O�L������o3}˻���VR��@�o3۱E|z�¯�^-mn��<�-]�{�K��dbO�x��Oj8F�ϝ�=��}?Ok�^����4��6�˲]�C�(ׯg�M��#���\�d�m��4�Y���Hݨ]%���\ZY�&R)�l�+�,���Z����]��������>����W7� �B�$�θ��&�<���攏�6���	h%�D6}s"-��� ��v����4��0'�R��w���	�6�����R-���9�3� p���aЎ�+5½V���w'�A���y�Q$�k+�?3Jܴ5_�*�k����</����Q*��w�ב�U��q�*�<T�k�r6���F��7]]_��D��k��;1�p��<���v����nm�c��a�9j�Vzߋ�=�6зZ[*�06vl��UoG:b���Cu�w��Yb��:�!m1�G�;vr66�BFE�=�A�8~�
TJ� ��g���v��ca���ؿS�o	(���4Jx5�5�N�#б��d��SR��+0s�d�s �AL�k�  �d8�Yyf��â^�{�^�d[@�c�`��lDî�6Ջ�|��Yp.�e��{(+�8�r���D)�	���t����t�z�7�̡TB����%F�|?���/z���W,(�'������n�������+�
������bݽ�0ͼ�;��5^��'s��Z��M^e���]A1<��0�ܐye�8��QAa �!V�(`�d(����ZkmD��ӿa�j�x@����2/��X���G��؈`�K��Z�P�%�ʋ�d������&�tL�^�'���*��hh�&s�:����4�}9P݂�]���c�-�,�`�L8�y{����6��·7�2�f�����_�GlK�"�H�� h�:@�� ��7@�Y�+��\>u	����!j������B�L�H�h�rkD����gBd|0/�X���Y����Ӛ��-�$���e6糁���GD��d�B7�KFk�f�iqYT�y8�u����t�z%ي㩤��F�S�5f����Ԇ�èx�c��h����2���[Bτ$F��k���֚@�BI)M0��s2Q��]5n~ϒ���n�[3)H�Hsλ��=�����)�!�"�Y��	�l��_�Vh�,� ��ܐR7{io�£��C6X��? ��%庍�&<���=�ͮ�����J�W��1��'H9;&���&��ɿ?ܾ�B�B	|b��Zu��X�������<Q�XA�H �(��H���&K\F�x�&��b3?T�M]P�������Y�B���Ѻ�:���IE�/N��c�0�/�,X�o�c*~y�|zE�ΐ�ۮ
n��c
�O�Q��6U	{u�A��9-�����kF���9���̽���Za�$�'�BZ:�Z8��/�.��\��"��7��"��҂F܏��a@!U�S~Z�uV�|	U���)���!)��,	�_9��D��6�Á6�Ӫ�<�ar�����,&D��%�*�@�`WY�{[e	�ZY صp��m} �P>�Y��*���lMI�,jb�N�`���z��mxQ��R�e�<�/&W0��Vd6�(Tb��(��Z4��KZ/pŶ���b�mX'����U Q5�:�Z#�K��'D��f�~�)�gj���C�����g*�f��pE�Q��"J�ֈ����'A,���{AD������5z��D�2I�Eak�j����8�1���7��j�]U�����*�ㆊ��@o��� ������$s�*Z e*a�w�+.�+jQZ� E��"3A;@bP<���b
	\�@�Os���Y0��~Ar�WޟMZJ�kG��yrM
��wߙvTMҼ�n��֣���W�l�lH���?��	4˜uǰ�MU+�����.U=z�l�s�'���,MFОj]�̶\���#�����c��=��**o��L����LH��6
�R�����*F���U6���Qx� ¥�o��HM�δajV_�#��|�ٕ�1�F�\s�Ћ
�3kp3VhOѰi!�Բ����u~`K��̅��x%��N��_��m�k��o�t6Cf��:�$���p
0iA5칠��+5��G?F�]8��o��Z���P؍�#�W���A�q����GWI��1�iwq�_��H��?vVz�ZzZ�/�!G�+�^}o����y AVQq.�]�|y��70�Gg,#ևi��C������4�7$6Z\�alJ��.�����/�U�ˍi?���
��-�;�灈X�@u��eC�0g����}��7{�lw�*�=W	a�t�$��Ԋ�Bȩ���?�w��;ʩEpN�5��j�fG 
'Z�v�ZZ��?~��m�ȴk��s�zmS����\_����	����AC�p�u��˓Vv�'�U��Ѱk5��>��7�{![=��uc!,d7��7VJһw�|�4��\� ��Cz�,��+�m{����"6>�ze}=�U��4�I~�t�;�2��_y͞��Q6u%�J�x��-ۮ�*�k���Q���k�E8���pY��r�}�#�P�$W�+���OP����(�h>����b@$7�F:>�W�����ғ:j��$�pI;�a���g���4ٲz~$+�Y�,K��S�W�xE�1,���{#><�{�V#x�Ò�u|�r���(-�g�Q`�:Nmb���5�WG��
X��UC'篩�?�brT mZ��+ �V�MĜ�p�Ii���H=�[w�i��xǴ�%~�g����{[ŗ6��[���'����}N	~���7���xnz
�c<�W���|����G�1���4�&��xV�a�aB
��}ϸ��Y�i�� B
m��9x�h�R~"sb�A��]��~e�+��3)����$Y���c���́*�"/�X^mAْ�A.\��Lr��͆8s���{9���iH$cBC�#}�'le) �
�0��d5�|���}3���*��uP�!aч�ٚ�������D��F�[��{�w����}^H�(���V���	x�K<6}�s��j�1��J���M��g-A�={��-���Qp"�v2z��佬�М�X䁰��BO�C_Wx�k�, �D�8��n2�ZR�����o�d�w��E�|�s4��)|!���X!��(����e����3^@ĭ�ҁ�Q�U5�3�w�2��55+2����y�ֺ��M�q����F���E�(?��P ��=nF(�P���Zb�˯��%q�܌ �S�>��s,��T�?G�~]v!���X��`|��髡�嚏*@$�$V�J�lx��sJ�%�zZ.\QC���ZO�P����۱�0�Tol�V%d����A�V�� ��I�`�&�Mq�ž�^b�IUsd��+!4N��&FPm�h�9���n��N���~вB�d�f���ԁ����KDS)�G�~
 �=	��G]���ͺ7��A��fBdt���fV6[r��ȇ\�lpz���7�����XTw�߈���rI���"%	��$|�_ ��?�� X�زi�p��x5ʆ���֟u	 o�>����i�@���S�P{�?�C���g%�7�d;˒tv��_��8�wn_��ځ��L�V!�
�v�^ �d�Q'-����N<�8,����39
�u��(��;:bԙY��������%f��t����c	��(�K�-y�&FU# qP��g����f� զTT�}���^D�̰�~|c"=?6�oM���Y�')	ǉ���w�*�j!i��?��%̏�T:��6���Ҵ��#�PS3a%�K��:(��']�d���Da�:q<�h����T\����g�h�ɷ��x�צ:z�--�?�c�پ�\�/����R� �@�!oM��Ш�od��:qͧ���8y��Z�!&����Eg����S�OSJ�I]z�����O.^�5kI�,1��&j�Я>�����8N����R<pkSҖ�v=�>�pJ�d
#'�"�	C���x�!�h��u��#}�����C�,!mk� �n7�6��I�O�J��A���܆(_���n ��V�P�q�Ɯ��gŶ_	�e���)f^�`�+d���V�'�q�mn0�|f��"�6HR1�!��92Pl����Z�� ���Us���.O��+g'ew� ��[pk�s�7���*�}qQ���E���o�s��[�ₐ���	�7.�]1��wQR���N�x~��4���>
���D���=Ձ�!Q�+r�&�	r�:��Z+�=}�#/e#��o�nx�E ����`ٔ2��ϵJl�o��P';-ئ���ȧ�}�i����^�k:��g�L~l���q'Y >�T�A������c��{v��ON���=�./Y�2d�hw��g�Ҳz�F7�wE���9��s;��Y��)�m�=�Y�M��=��MI�>�hYUMnfPN���y'��6`��VW&���6�T��0�~�t	�>?G�����<��!qB�Ϧ���]��9��Q|��7B�BR���;K0g�s�u�<��v�����5+|�����# ���n��_��6 �#�|�@uv���|ڊ�V@쁑��*��ܽ��^��kƹtʅ�%��W���nD�$|�`����y]��{��\�&�;:�����K&����q���9�n�	m�����Z��p���nicƉ���%Mu����i�O�0��W�jX6XodZ6�[�Л�gx�<�����#E�l��Eu�*pQ��o�S�������A��J.43R��8�34#fm_'�()0N��Ƿ���
Ťސ5z�_�e�dy�4�.��aMSi�6Q��E-Ň�幒�
�5��_}KQ��8�'nH,�!n�`W�^���s`��c,{�m����(��
�Px�zs�X��ba뻒��:b�'�Y�%�)F�d�r��&���@U��IR�4�S�^-�֮y���3��7�rv�����>C8�Op?���,�dC�T�ŉzLe}S�4��yp��~�6�=uh9e��/�Z����#��
�~?������zm�-&1S6��n��(�IV}�+���6��;ͯ���׉v�;�ݫ��{:�ї?L�a�ha�a��:�K���p~��,�6&�rv��'[ez���z��ṭ��H��b��0�e���Er��<WW�́�_�$A�œ�|��j�P/s@l��ҝFS&c�'n�3Y���0z���.D4Ш#���:N��$Y��dFu��1��X�~�t' �S�q���{I���EL��}Y�:8~��t$g 4]}:�
G&0�p�1�9�}�ӳ0��ԙ��8𛜠D�GgV�z$��qb'�H6ǔu�SN^��!P)�˒�[�C�:�LN�*�΀̾Р�d���5��]���z�B��!ٱƹ�ʥb�\��8'�'�q����3��@��Mۿ1�+a��$bn�#>�,�]�͢Q�@8��q5:KU!p��(��֊EvS��r�8�|]���v����E��|���y/8{a��M����P�$lj����p�u�N`��ߵ�ؑp��i[��U'�g�}G�70�Ji�%�Gհ0{����o�7�1�8{Y���|���,�����kek�<�&��u7r��$���Z���*�׍7ߣ�PD����.]�vn4ce�1�%A�nA��/��/�w���L���!A�}�7�,מ��|N���6c�.��^؝�]�C��N��Ϲ@��) X�DGG�D"�sp��AirF&?,��v;���,��i,�s��{�|{	XaŨ��?N��E�s�h,����*�U�qz���q;�"�����L䀸�4�mu�EX�ߵ�3��J�lڐ�٬h��d�Rm��������:IC�H�ˑ�
lJv�1j��)�nV2���*�ʁL%����S�Q���s'��ַ��G{\�D���P��v�B���,(��TyHe.Z��a(.��e�	���|6���@�gj~�X��X��*�p�ň�zx����D���EOn���&	r���X��ks1y�y�7��@�Z�Ԧ"�f�mQr�S�&��a���Ays(B� Z�t���XQ���μk.�D�(OPw����p�r�:�fG-̷�@v�|��}Bm���ئ��ձx��r��u~�%z��L��u��p��ݽ��=x-��G"BM��-W��C���-ix_$��<&�WJ�5p��
��k���Ä=|��i\�V$m��I���BY�ӭf����VH���9��"avꏐ�M�`�>�Ί���0�U�
�i�lk�{%�5Xh c[�[C�����GȻi's���	�,]��B�ү(����Sq#��S�y�c밌�h ��յ�]�����B}�c*��� UX�?p��ԼN�A�I���:���B�}��.����/�s��%g���p�D8e�zLa	AJ�Byڦ��z��n�\�򑁺�]v�r�5fi{;u�zrޓӧT���7�Lqې	��5tN�����@؊�lxvǊؿ�ge��>4�yH�8���,=+t��ǎ�q��fY�����c ��r!�-H���%�ͼ��c��&�fc��a�#&7�����4����ڵ#�;��Ur#�����	q����l�Y�y���)����@<P��C�$/�C�����9��aSe}�Вk;�jg�2P\��������OÆu!�zb`�4R���&��s��(7"��h����e���D�?`8"�O��<��qnr���ʯ���
���T�Cp�"ې�ٓ�~͑����p�e��,Ey� ہ*����=__�*�p?���&%���@9�%�*e@G|Վ�|7(�3[";E�� ��:�̞������p񏺔
�A�����z�-j]�).��0����Ԣ��8�)�%��`.��Ř�Ɇc!��V�`���ZJ+�0V:���"���@Vh�������y����rU꧔9T 5�%^�9�y�<K���և�U�-��%��2T��z)�9.?�L=&�G{�M5��� 3h?�[\ܗ��)F*�G��}L�
�y���r��S���2;��/�X�j3?Y��}<f 57��1�ü��s�{u���[�A���(��^ϙ�h����թ���h���Oq��Tp��[.��\�ϨTm3����,���v��x2<�0�|,��:m�j��I�����`��'�F���phC��8u�;`��������x��O����AH����w��{Mi6k�p�j��������m��s��'2��^�M%xg٤���#�X1���j�)o��=���YI&)�I�F�q/ľ�9=W��X/�@0�b��>M6"�ڰ�8c�M"��X]�[��J�I4���,�w���/�H��{R]�@]���,�c����m$�Q�Wx�:�~�����K?�ԉ��M�H�.��S�5d$�	:V^a�������{ =de��~ZC��y�ݼ�f��f�ȣ� [�k5}�I�8�G�"hZ�W����C-̛1�Iw���q�3�s���>��W�8䓮���j��ｍX/M���|]�ld4�[�
����5�"��h��,��������sqgj�#��#�3�0q��%�����~�b+}VP#��`/�l����
�C
���3�&�d0�	0!���+��Hr~�}d��VՂ3�M`��L�䭚����ZD��B�}����D�A�y��a�HL�#a䯽����w落*�����mӵ������"���t|��M���s��������M����-�S�nϰ�9�Mnu�J�a��J#����y�� '�"'��+�B\yPyK�u��L=p�`ϲ�n`�L���#�{:�\�RTxQe�47i�zңU�s�.ƩȺ�^/���@�`Q�]�;V\I$��`���1�xl��n��&�u*���﹊�Dy1��U�,X7���S�up_!s�",�ͯ�d�Q _7���Xvٺ@��l\�;@^�)}G�E W!W��+ �`�?��TN����%<��H�mde�䟔�r���
�7�+���������3;���"��N������"���X��F*�j�dfQ��$^�R��u�?!��?�y�44��)F}'%
���@��/0_��-u�RE�(����3�vTv��Px��F
�Jz���ؓ@<˿[aG�HR� �?�?A�	��dZ�Д�¶=4��~�d�V#�?@�t�Z�N�7%oj��qћk��V@�Ne�Lx1pJ%����G,�XS�ڵ��HR�Y>��п�Gk����/�E��O�(	��l'l���L�|T���9���:��ޒ�Q���:��u��ý=A&�ЦZȁ���+
����nlH,��85 �d%⏅L��3	��l�)ꅹY�?����D�{���e�N�Q%�j��S� �EA������`?�k  ò�6"N�粄oy/~3�3/��KF^8A���v�6��qx��iϘ98A}TH����-,�=����2��Z��0�#��S�����GTk8���']��nq��P8K!s��G/��[Oo����qc��\"�!�LI��F��C�B"dBӳ���U?4���_e��h��7{:� d�$n�ߤ��>�t6�X�,D��n���hW�rOH�x�ц��ԥ���0��sO"U)⵻@X��d����XojV���������m� [N��D�j�#0'D[�j_��"�B�%p��CM[�L�`ğ���4�㲱�&�hlq�qQ�ھ����A���
U1��&�G7<
h��s���OCI�iʑ�LòZ����u�DyNF+��2�.���ϯq�s�)�+��ʣ���8N��X(x��m��V<H�j��#}u���Юy4՜��='���	�ϲ:-�ۛ�s�S�/ O4_�1�l�#���1���|���]��3�B�]>J�O���aP���D`���)Җ��U�T+P���nԯIO��FD��Ѷn:��$�c�f������L�'���(u)��>~`�H$L!��F0��j?��JU3�5vgn�8u����h�U$�4��#�(bLo�3����| �^c�,mF��ql^�~�o62qgIkV�V�����Y>ڃVs�&Z�352������T�z��rP�Nf�J�:6Y�	)�RD�(P���A+�;x1$��EBu{,���T� L���-Q�����Լ��9&����
�=��mـ�����H4=�4*<mVL�:{B5����N�Nw�-%)7w"*�����j�u���j�.A+z;��Ѵh�¾j������Վ��"x�z�]p�m�@�z�x0,�^v�vR�k%�ZL���lb��xG� �UtO��mX̫��]!�s߲�g���4�<UN���8���3�]�6�Ll\��O�\$��s�C!�g/���4�%7N���/	�n��C���U�nyi9�����������Q���f��eO&G�K˳��(Q�XO�̅Iܻ�����x�B����YC`��O�$�}S�)�1D��愓��%���TD��Hb�uF�ˡ<?#�HNݚ�o���Wɨ"1�$-����X��_������_w�D>�$��/�I���J�������?!,5V�y�S�?���O�}�p�+p�Zy���X�d���!`G�zKt�-oVh����R*�������'��jMA�6�'0���D*�e����	X c,��k�zbU
=i$�F,�C��d�4�����)�Y7���:����۹�a���]���D����`�l��e���;u�kP�+!pā�`w��FT��`�@(��ۤy����)��ٝ�x�/"�T�PV Bk�}ۏS��%.�3��dԈemA�I�|�uG<��gp�+a��su8?q��t��X��\�-,��*���+��U�eYLv�� z�>]�љ��	�x��=�d���e��%�䉅z�Th@T��e�)�͚?7�m�u;�f�I��oC���"��x ��O/e]������l����m�Ӟ��mY�]9i�sN��~8-��"��m��c��ir�BS�Ee@�C��Pܮu�M�&�����WnO���V�^v��������Q�е
Df`7��ҁp���L��!G�	`\��GÂY��m:�~O�/~��g��������z�L�.���j��c9�9e0QT����k@��k�ʰ�{�`XE��e�9����t��>����7n+�qO��Hڝ�:<c���έcz$�I�K�e�F���P�4/tE�t�1�����PQB�>��R�!|c��G.�,�l6C��#��wg��(Dr���|�~��#xIT�s�o�r���E�v	�E����Vc��V��W*�L[����t�q:��T��@�1�����Ǻ�g'!��˰<$k��i0�(@�`��� �;6��a�C �F|`(�=8�,/!�Z.��ܤ�S��H�]W.#�b6�G�8���4���
�P���.�T�j����Cǿ��o.�)�1�s��7/]�v^�&����o�2�=?Q���viȧ�w�Փ^r?�/�X�E/��(��T�k���!� �z5�E��B*at�)h���R��k�*�T���xE!λ��U���E@���I��ӧ�d�.I������d���l.^un��I�H��W�pw_?��`�p��+���j;�T`�F�]2܇2l#�6}�XS���=i��r��t)�@^�2���Ǘ��u��{��`�}�m��=u���:EOB����yW��׸[/Lf?�˃l�O�������GWp`�ڹq�Tm*��+�#�-�D�p���]U7;����5�0��>��m8��̑����3�AEL����u�����:�2���k��0S��N�`g<�V���@L"C{'S����0_��@JΑJ2����9����� �]���z9�3�@VS[�~�E�ktVve�1FNs�s�(h�ت�>��3T�l�؄��yPL;��D0E���R�=�ј���K�� OC���kGz�Y��y��6L�!73T_$�]�N�麟!����?�� $H�o!} ��=2��Ͽ�7ZA9)։�j��қI;��A< -���-9}��x��@p�٣,�/ވ�'
J+�&�`[=9'jڒ %�C�r�)��kմH�w�}�v���ڋ�5�RL��M�K��MuN�2^�w�����^���5M�l�*~i�mS���"k�y%������1��!!������TR[g7�ځ.۫d�O�Pwn���	`7[3�+�SK݉����������o��!���[����m�c�ٖD��[W�np�X/�m��Jo�f�w�������(<����ErD���o��q��.��+I��=@�x3�)و���#
�ci���+���YH����ܑ�M���G���� ��sY�M��9��{<�q��Z[��dvL����5Χ����?�����2G���(��H�Ա��x|O�`������1S8D6�ݳ(������)��I����}ehI�������}�F�8w��_�T��ѯ:�N}����g5���	��w�)�ء{U���b��nU���,�x����Y�r������>�0���_C�4��u�==1��C��t}�G�eo���~�+��Y�\�Ó�9���*���l���.%H���CP�LV<ߣwם^Ëb�#W�բ�ftЃ������v�Q�@3���h}���H����$n���6K
"������K�Uɹ�A�
�S�$$�ت.��m�-G�G��s��{�����p��Z�B���M�=SzS�7cw� p���،�6e����+/�T"��X�6��f�T	ym�*[�0w�=�Qǘ��>YU�E%�_�Q%E,��D���a4j9r��40S�AukMNoM�)�]1O%kN��2�b�L�j�~��=��FRS �5Ǣ��h��F�WUl��q0�u�9�'G�|"WHU��#6
M��J�]�$�EWZN����"�PV��R�<L_|]6M�b����_�Ǌu�r���F]q��\�u�������+��N�JƆ��4BCZL�A��K���5o/�e��[�:�t�~G۔�#,.~G�9�����%��t*vD��Q���C%W�P�O�Ei3e����+aя�h���KF����ݥY��\G���ЬjD��ߚ�ad>`บDuaN�����L�e���*�_(v�9�٨��	Q*@�e
y���X�G\�.Q��ŭ_Y�z�8Q�����8�O��&��d4�����A�9@ek��7���2�4�o�!�{y�����S�!AGKi�G��]����J��ᯈA}�x���f�Bgz�@�\I@O�4����ga�U�^����w�CtL�ֿ-W�S��$>�7�o�w�7r�'ǥ98��<�p�*QOv�"RR!��8
��z��]=���D��� ��
���3��ϺH�J�*_�J�ㄟM�ij{H�Q�����b�L�l�v���B���	�C�]�q�I6��C������5�+�NH3��X<�ʺ��2�� J�ޣz¯m���Ѿ��-��=8�����*�����D�+�ݕY"��ρ`m2m��,��ϟ�M��)w�c��J��f���n@��l�3��kQĢ�R�zUK�Lm��%�k�~��M�� ����bn��(�#���4�MC�:jJ��/�A�0�$,;J΋�#�F; Wyz����]O�zb/W=Q�40���ޮH�ȑdE���W|L�ж������\�wImj�T�{�}sCf�89�%�0�O�?�YK��`�N����@�:5�3�OT�%���fB�����
�b� �y��o?���u7Tཔaݪ^x͕7����iIR9u��A��\�g��A*T���✨�����S'B��#Ҟ$=�Yz��3���2�1A�:^��.}��7'Y�M��	\��B�ȨR��	���1g� .�tH�Gv=ʗ��"Cd�=�����kC�<���sZH�NV?��u�&�D�Q�'�g�IO�D�a8� ���'Z_H�WQY�aT`�gRc��u��^�����p�|I�7�U~�ak�@+0���m 4b�0��Qx�5�/��xd#���eڝ����=�3//�\�����_�_B��D�B�Uw:h,�u&�v�>a܄XC&���"Wۓ�
3�\_Y a]�r�����%py���@��0Ԟ�{�`3�Z���_7�!�Μ+Q�ᳵmE;Sy�. �q�k�qճ?ZK���D���l�K�L"��[1Nx͘~F%.�����.f�Nbl��,�_:|����r$i�xZ^d$�5�]A�\L�P�����}g���{��%̯�}Ϛ�j����:�|S��X�W*��K�yd��;���d��������Z�D�A�ą��Z��A� GsX���K�:�P�L��vw���m
A?������#��s�cc��ɔ�߁כ����Jw'z�j����+�5���y�=��}x��0I$�PT��!��w�S��F�u����c�!ܰ7�ǋ}���W�T"�� �8;H'��d a�K)�v��G�����q��'<z�T�e+j~�pW� �I����<�gm�m-�&�P�}��>Fi/�x�]/V`�q��|��& ���q�X�Z�j��f�ʪʩ����Q�&>� �Z %�������u(C��:����_�A��v!�o̗�?�;�*(߰���l�a�}���T��U�*��*�Z��sf��wG��#��������jWv������I�(}��~^v�,���W~�g"T�s�	\�}���~�[=𓌰*_�QSsPPR!��L@#JF�A�,H��GL[���&hk�U6�1y�L=��9��G��'��D�����z`wG1=���Nw�U-ypmI��Q-s��N��!�l���me�|�>��.{��;:��>*逄��GE|��X�G8�~5���-2�*���@I�`O]pd8�>���aw;��UaK��}��.����	t��[������F3�>����S����V��z��+R�6���Wn���ظ�m����яR��_<G3<�u�Kfϰ�AB��o;yD=��Ŵӏ��i�XW=6�p5�ݧ��}���4@^�����[�.9��Q�b���x@�;�7�s����CG��8
��m��j�B��Jj�u8��*e�ޒs5(�-5y�%�U�	��\d��T��N+#�ST<1�J��Ô?���qYWV���Ҝ�b�(l�l2R���#�8p'���{������p�e��A*{�X#��C`"���	��
���hR6�_�+P�J��ʝ�R�t|�e1L½:dU/�}vY��،��n�O��n�(7�ߦcRkf�(͡�(�a�Ź�9�UA�51�u���Q�#W!������+\0�!��\�!7K-&��	��Z2X�"O]pf�[������&��Q�vra��֖ �
^�}"B��,@"����L�z�B���H�@]�����+�s�2�����6�"����M�V���z`�}�z��	�W�&T�i�N�N�����V�,�S�������-_S��tEpڸ))�C��/�f�����%fԫ3v&G�P��R @t�40�eC��N��a�JI��w�6�S�r� �<��,�F�/7���rzyB�Ŷ�r�`�Eh��Mr��$���O]?����G��Km)�Y��Od��.p[8fE+��[N��W̲��\޸*�zJ�^�^Bm��i�Z�H�mCo����ﾇ����t��}n,����.���.�X2�W�9��!��6�u�Ga>�Eu��$�cEP��	$L�z{�9����ưM!ԩ|��+$Rݗr��^��)dÏ����ʛ���x���=h��c�+�C���3`px>���@F7���^��\�;��(~�G�'�е�4��鶳��/>HL����iB��[G�c��C�㯛
N.v�9#�} R4���lD:��S�T꧊���D�Ss�
:�X�럲����f�hdM��ڝ���F�LA��q��V-,�[ݻ�"=�+��]�bSŹd��"*U7;��t,t*n�g���&��z�ک���	�rpШVc�F�ЇƹӊS�tldM�i����NY%��neëe77!�N�3#UO��n�`�̽���e�d�E��&����/��X���!�i-;�jn��wy��ڰ$�o�E���SZ�0u��J�i���9��j��{�V��_#��*��l#N�1.�3�R.?Y�'��-���G�ߏ3L�t4��4�!�n��gmϫ����p� EdX�[��y^%�.H�<�s��mW��G�v\l�qA	�f����h����&K�f.}�::	��͒ި�L,�ty�(�-c'����LL�Κ��-�H���>Z�k�$�\Z��6�b��*��zf��.�v3E�k�H.��-���=־|�L ���H��~|�m,��Vx{�U1���j4=��*չ<k�ƌ�ń^5�e�g0�ե�[���#��Z�kYd5���|{1��֮pum�s����6���i8"�3T)�T�Q�#���=�D���Y�*"FC���]F��Q�����,���/�}!G�qM�!Y+�ܕ(T�?��R���3˚/�l)g0���-ٔ��Hn�Qt&�c�Q�Q�K���C�?,ۂDUs!�(���r(Tɧ�s	L���� vy붪vH�):ąf���U
z�!�5+��B��Ҡ����Wzy��Z��R&]C3ﮄ�9��vcp�R�>m[�����F�u����Ρ����b��1����{<��4#�C���g�4�*8��}��S�P������*����m�j	7��
���dysp��h��i�O�6��;�fX&�$#O�n�^u�?.��C[��af�!q9u~~h��y�Š����L6�׏�F�lE�t<f�׋�rL� ��K�0>R+X:���f~{WP���!B���ϘK1z���A �����	1=��"�BmG��,��~_S[k��(h��5���T�tG�q� ���`�|���Oy7��)x�0? ��ٖ��k��RP�s{�e�fyA��"�^������&��ccKqƃ�].9 b~�EV�I�^���B_�}�^܌���� R�@則��a����Y��QTh��U���p?%�`�Z{��n�	���T|I�I��s
_�*�?qj+�dHǤ����c��ڤ��ULm	!R�Nr�6��K��:�<�a��Լ5��z|�
�n�������R�ݣ����!�v �i@�/dt�a��n���L�ee��8zG�gu)������M��e1���4w0�Qgҥ�ݷ�Ql���I ���q��&�[�;�˙ƵLd�~�ߪ#���Y�d�v�v�t�xH@c�M��P�r��2ʺB���2Y�Y^/����L侫���Y���b�Д��i��Rv�S��ы����p7�}TA�	T2�g$8��r�<��ؐ�-�� ���j������T"ϥ�>b�;���f�^2.�W&W�0b�G0k0����#6^��H���A��=����a��
��Ŭ�vN��0I�u0D�ҵ���)z�n�CY�pg�G�BcZ��E6�)���j��e¸@C��Ih��H���D��y���(zU^(�}��^)Mh]�Jged�v�"x1���.H��@��J�p;��䐈+��j�n��j�[H�2L�D���:u��-Dv�\�����S�rP}�;-�y"\��-oI��C������&&m�(�pcPK�Oۭ�t{�`H$�Dު��lvf-�L�!>�-�$��F	w���4;���z������_j ��[��m�^],��ne�ӞA�o����~�d\�T�� �*<�����8���t�n�%�%��%�mE�Ym�:OU�uT�;���%-Q��h�o��X�[��J��E��NO�a{v�V����}�F����A���jg�^�ȅ�?3t<Y$��W���ڠc���~�,�PZ[�p�N�XL��c�B�b��zc���o{��G�I�p�Nn}��S������D 7H0 �0��
K+��D֥}n+.hgہr��[�Ȟ����1m��(^��)����^��Ϳ֯�S>�):�G3�8������d�L�
	ٓ\��S��	.�]N�J��EvA,X��H6e���������i�G=�e�O�˗k+���爢������<�����I�8e݀s�hH�ڔ5��}访�;ϻSE���7���Q.&�*R�V3�]x��nO"o���I�j+�O19�Z�q&�s���<R���g�ڑǤ�WN!�GX����O�l`��e�4f��x�d�b��4?;�� �`�GL��s�0�v<�>ŵ�W���ǴF�.�?��܉!BTZS��&�
��w_ey�"S��/&n��6��r�j���JB?�v���bu��n_�@WW�
o,nL���H-��6w�����+����@f��+��!��i�,�,�@Mlz�)1$vޜ��m��c%�6+�S��y�G�"'mF�����V�~h���j^/���cN���{>l��#��ˍ@y�sEx���{�y>��!�}����~G'c��R�\���v�8$h�(l��t6~;R�v�A��w���� ��Cg�"��&��59��R*'5��.j6`O�a�i�׿��{2�Q��wh���=5W�~�ʨ�y���࢕�����7YlO�Z�x�,4��ƪ�*~�4�Se����0�I�U=z�om���Nݧ2�܍VI����$ɖ�*Γ��F��Li;:�Ϫ�=��Š<7j��R\��P��e@�YL��L�L�����G�쓼j�V�W;� �h��dm��>�3�V��dT��.H��߉(L5��le�,�np�s�<�Y��W��������jt�zؠGus�8��\�(��߬e^�S�Ѓ~�/6N��W�dD3���"};�O�g��O JK@Ęhm�w]������rS�w`��J?�p2wW�a�.C;p$H�ށ��oP�����i��N�
��H�jKÉ��#`��~��E��$�@~��鯀!Ȍ�� ���H%ߧ�H�I V/�W^3��'4�q�Ɓy"6�`_K�K%�Y�A ��_Ľ������(�%�V[�9�@�>PK��X{H���ͷ3���E��p�m����|��/��e/W�_*��B>�lR} &o���ܺ=��A��6&�/5� ��тS=�Z2R�sN���.%���g�&c�P�fZe�BWt:s��M�kZ�Q�;m�W�0f�(��oe�Q�9��뎏 �C)  �j�%{����?J��b6uh�2$tC@xl$?���JHmM@�mX��!d�H��*�e�<��E���ه�H5�<�R�3�����&}����X��l��]�@S[<1��&���?a�/�'����xX���T0Տ�o\	�&�o����>�ݜ='ey���G�*���)լy��~��|!`�,��Y ��j�:zƲ咨r�����B��(-$��H <��Py ۋS1#rH���x���[�R�l�S]�ٗ��r�������ze����߆t�G߳%lZ��F�vC�-2����y�QCe�X�8*�Ϫ���rs��T$�f�;��1&D�$�]�g��3�%n}�ͽ�;3�4�)$P�""���%n�l����ܠy�#�Oۤ�Sx��ȿ���$wZ�	����2,~����E�(����T�Pjw�׆��
�ʨ<�73���_	���#靝���L�@�%�V�0�/�_U���/��ƃ��+�F�Y&p��Y6�0nP�N��$w���(�0]��ȁ+�Q>z���%�$���P���c��i9v�'���V���h(&Om�8�!q8�q%�ݙFy^[��{�f+�����WX�@���8��:A��ۇ�"�=��'����G�����uj�R˪�g։�;��Hf�AA����4* �Ԍ#Qˮ��b	��N���!���*N����#.��Z��c�9�>�In�ub����<� ��i����Bh�Y���t .�
�@$u>�.��qa�p������L!�B*)i���5�'n(BrX�F0As����yA3]Ƅ5�?U�i*ҼA�O�_��f+X2BVO�;�\P%i�EA����q��2k��mk%��$��G��Û���8G�������jBh�`���:�xRoQ���ہ�%�����ÖP��*��~K�n}�٢��2��޲����Q�b�R� �E�_�K�i��Iy E�/�(&�*j�A�ﴺ��c��.3���ʅ�s]��?Mq,ba�9A�*�C
��+%ѺQ�P1�$I�^�2?��v0�Q�a���rk���2֪�}E4p!�`Hh���K�)��Zտ\O�Ib<{A�c�Kb�� ��)T�4W�Ji�	�5
k��dz���z����f�W�2/b�T�%��^��u�/�c�oo�`��G��:;�g����T�g���;����/a�e���IƎ�9<�+��l�P8W>�D�{R�w)��7�h�n�M��BnH�#��S�҂�E�ն!r��"�ФLE1�g���i�n�S�&�{��Ғ���1�u9#�5��S{ 9����ʎ�/|���zR�ZJ���[(�{�}ɿ�X\[4Tb�ǭ3k�g=
��@��#[��H4��r1�H�ȩ#���q�ˈE�M/�%p8��ʩ��+��� ���&�v����^��kӱU��r�+G�m���q��P9�d�#ȍ=i� �U�`5W=��ȗ�{g�)�L��C;���:�'X�{�\B�V�]y$���D��A�a�+����6s�Q\)]�){VXl5v�����Ə�K$�1��eQ.B���x�6!2�sS�/^��V��<+�Ѹ��7V�������1��Mh��
�)5��lԫ ~�����!�K���0�s|
��[nG� �ϴ���|YT7T$*T���<4+���j�.�ԓl�W7�P&ݩ�<"-s0qH^e��0��!@��9_7��A��\df���u~�h�s�`9��lw�牵e�j�Pwс�cY�"t~d�9�j�P�~T���e��H�'�s�S�?�� �q(skQk���u>�W�\�.�5Y+�%��Y`��kM��V�Zx|W��}����T�2�W�rJ��FB�8���m��X5\��ѾB�d._�õK<{+��@�QV�4x�^DȊ��� D��h��q���)�Bs��Ɛ��ݼ�Z~��D��ٽ�7�'>˘�xH(H�u�C���ctf�L��E��J����˦F_��0=+�ţ.���T����Kޞ����f�O;�.��l����]8t0ܹ����3S��G�~,H�$1U(7x�",�	�pU{�l���BH�cǳ�axH�.����}�*��Ҷ����w�~��)؏��=��.h���qU����1��V�Ro�}��H�0h>�����c�R�9 ۅ˝xB����m�c�[G�  �o��B�Ti<�jah���YW���^��\�,D�J��Ѓ�S�Q��o¡s��s/b!���Qi�DTƦ�J���d���gs�cl�F�_٨E./�Z��d�i����HX�x�GH&E�K3$x޽�T�����Q׏��
cm3Pc��@#��
�bi��6��ҙ��� �&��r�*��w����7.��8~�����u�+��_�a]D�YCRTb w5� �?�=^J���_&�_O܌�n����3b�h���/�x(�M�@��vak�?�<�4t`��h3)���犍�~���:��9_;f��N˧��Rxa;ߊ��Bװː�w�b
��\�G1;�4Kɼ�*���D�QR�X/��3��*����T��ʛʾ��B�T�G�d�7~(�)���lW��\y0�w���I���^�/��c7n�W*m���+'S�=غ	w��r\@@A�0֠N���&ソh!�����#�ڳD��:�`���zvq [#��kn8��y����	
�xP��X%��j��6��n�!;�?�Y'c���i��;lc֯z}���P��?�9��L�V�n�	��m�U�"��Q�B%������X]6i=W�}���2O-L��K����8dNhd ��m�j�v?ov�6�d���>U���r3����.R�R��`�@�&	��,�8*��hCe�U��1��8Eu�1��֟��)�Q���{�Ր�'�Ry���t���j�Tyz>ɠχ*�AT7�wb���k72V܍�W`E"��Ky���L��x�.�Ɠ�R/��|�f�����V�r���Ŗ�,��� �Hw���K�)�&�G䬣�O1������Ls��n$�G�g �����;{'�9�c`8J#ܥ�Aͥ��*��r`(�$ڤ�Xc�Y�n@%��+ �r ���s�d�G[�F[?=ƣ�����J���W��zL�-G�U{���j��mH 8)��/E��B��NæfM�����eǅ�y�.7Cx�J<�N@�ԽL��q�(��f�tgMW�j��%�����ƖO$�oz5���0���x+��g�3V�רg˾�u�E��hϪ�{�Wؓ7�ZMTF,Zޞ�k�e��k+璖{T�6�ǔ�YV�ɐ�7/z=���׆]��������=S7�++�����)�B,�I���ͥ��w/	�'��M�M����lT�29�gk��v����i�;)�:��ǩ��HHx�U���,�M-���h��",��p����+��ן��x_��.��H]�J� ș��6]�̫&�K3Ⱥ�?Ơ��xW��h���O�^��A+��0	 ۡ�)-�Q���4�SA���u#��z�)��.�n[��`�����`A%R2�O�]x�;�&%z`Ӑ%���OR:��s���������������X`
���C�N�v,p�t�	m��N�Cj4ZmBK��6VMd�*2n���l����`�d�`B�Ы�dc�dA�jn�9^{�t��5�_H��/w����:Zo�e��Ml�~}�5������Hf�wUܺt���� ?�Q��Y(o��i͓�"Œ5�T���)y��M5�vs ���pcxNN��C�NFꈖA:��� v���Ϟc����_�&UD�*�p����~r�S���%-)z�ȶ���^9_S��%�fo�h���K��l�+q�}>E�̠��*��=%;��dSd��6�67�T�LJP�����+���O7���i�o�5��7�9��zp����Ϲmt͟ޙ&���IBp�x���3�*��?]�O�����}�l�$D��6V]-�A	T�V������� 4�'r`?zt���4�"���o��4c�4�ŝ��25��T���韝4������ǖ�RMK�|�����3�&��0��Y��j��_2S3g��V�!�h<�ՙ��W9�A���|�oI�����J��Dd�:]p?��ߞŤ��"�ӑ&�,|�$'�dS$���K�Pm���g��}���	a,���1U��|s6d	?��5���3|���8Ċ�"�NO�:�ܙ�^}��S�f�4�r��n�b�o�,�V�= �ړ�;r!�7f*u�P���=Q���Y�5엛˜;�$o��'	�p>ў����1��y�<Aj핥7;�������E�'MR[��?H�����[4;��t]YN��1I��|�N{��f��^�|�}4U���m���'���>�@f�������*k��2��[h}E��g��41^����&;�tR6����ci����۟n6�������51��+�� Jj�*���'�N�MK�-l8B��ɟ�G6 ���1��%G���j�+cc �nC�6A�J�޶2�E���DP��Ik�{�5��_UHw�:;����s4i�u��p�RÉQ�KA�&�g��Y�+����?`0<���n&��i ,;P�j�"�C,�
V�+�2U-T/؏eHT7Eᔸ��{Rx)��.9�����H^yf�8�2���O7Od��ܞ�-a]��y)�4��o? L�ѝ)褕f%&S_��T�D�|o��xub�ӻ�:)��(9V�'�ۭ�u���(��,w���>��yʥY��P��Q�D�G$��4��mV�I#�����Wz:o�>���La��=132��.ͳ[�!��-FΔ��,�3�y<	y�鶥�n@����:t,�B\��9����cx�g_���dE�� {���m��:����:x��8����KT�0���f�4�i�W��8�-��Pk �%	��cΪ\���Fp�V�43 ���xG���HQ���)�a��,����3G�Y��.��M{J��M��p>�츞f9�kR�ăR�{(`Z���m�EJ�1��ʢ��m��"�����}�`����h�P�(B��w�m���f�L�
V	�%���02���i���L�a�؇��Ş_�R��2G��#S��ʸ�7zrٿ�D�rQq7�/kO)ֽ#������ø��|ik�H����᯷���Ta�T����S� L�V��f�(c�XIW�����TѠ��?�ωs��c�KQ����v/_�յ����X�i��Wpi�\�$�`P/���>nA3��[���g�G$�l���CŚU��F��Z���R慁e-��ӆ�����E�Sl��%2->��1z�X�y��Fz�ާ�����"ЦmO{49�bm�����<R�]�s�橙p���4k�x
�r��Y�c˭��M�������1�#%��	�7���uC)��?B+�K����0 �SE�q��3Y��Tuӏ\L^����p��ܕF(��˿�kY��M�]Z�Ӆ�!���`��^6���:-��f����ɬ��?�e�J-�i�H��\DGw�����8NDMe\1�M����6��KW���^����+����ٲ������>1�n�g��Zՙ����4�23���g���Eۗ�Ӳ�<%]�+ʵ��֧��G�L<�d]۸b(��մaTv*I�BR�<��s:�O�9��rmz��7<F%�1	��h��CZ�*U~	�>�:gU4� Ý���rNin���(p�(�^{�y�����3����Lk�Y`�ʫ����9ǤE)|�����An��Q}0��rA�a���ckGC���x!�W�������u\��+��c���e����q��6�yLe�����DZK���[&��c���+͇�t�p�������|w�4�穉kt�O�:ߎ�|:aD��}q� પ�)��f�-݉���"N�n�G��mt�jJ�o���e5.�8�8�@�<�%����&2�-��*ǃ�Z}}�T,M���m���w3�M��2 Vh��� (ӑ>�k��^���(uF6D��?�@������Z�b�i�F�~$��a�>�v<��z�̓t:W�� ]������ �-BE�ͨz-�oaa�u�v*��0�U���s���&�=�u��J��g��C�}*��e��H��fO��=�B��b�������Xg��)���`��zQ�dS��F}���k�j~.�ΩQ;���ޅ+Qi��V�bt
<c}�!G��	��0A)m���o��~2Q�W��Z��Do76��m3l�ƿ`�,F��&p��
d�����嘪ʖ�����b-�mv��S�uNq���S�V��g�y�P���?J9���R�?� >>����H%����pL�ㄦվ��gV��#������ł�(wpҲ�����; �e�E�Q> }MC�egcOsj�0�t_�;�)�V�hn�&,�7�Djm!� :l��zk����<��1�ZU7"�Ygݒz��
#+�Z�M�S]��:�M�'n�s*����MO�>h����Y�n�=�TrA�n?I3s�g�ysPE˯���A�<a�{�_�q@��TQ�:��bj�FE��[s�Z��B�� ]p{6ՇUٶ���+�[Z�/�.�_�x�X�GRÒ8�[ߧ����+6(�����}�EɾqtRQN�=�7{�O����m�I��hb�9��Nɩ
�Jϙ�R]�h�ޣ�MR3Q���y�gd-�#U�(����lH��<�*vh��HM��OH����+�W�_K�@��;b�� {Y:�pF�R>�"����r�5�"U9]�u�{a�N�jK��<�0&�Ϲ� �*#J�q�5(�����:�R�>H��cM�vw�z��\�O�������^���	��/z4����8a��=���>��t�3�ܵ�0�P�@�}������d�Y�?�1I���`�����Ք
3k�P�"�/U�~������2m����M��6h�rZn���.�G�K�t�����<&�A
����-s�-a�����M:QOD5˝��8�R$����us��o2����(��#� 'H�AJwF�ؐjR�nQ�x�*� �IK�yN%��t�y�E2SE�\���W��:#�LH�t�@�K6�y�,����Qlk��DCL(�d�Knn�Ь4�a\�gK�Mi.��9�:��4P�.��Ø�P '��l�R�"!݀+�7W�E�ܮ�AH�4/K�D?2Q/�(b���ưFm7!M��s�1p�&}T��fVV���Vj$��Nl�8�)�O��j'�E,�z��, �|�� ��6q�6�?S6ʜ�ve��ҙ��-e$�S���,F7֖m^��"�:� ?!W�����^����*K�K1K���J���]�����R/��SEgB�`�����l����`Ip��?E�M����Uȏ�N�aq{D���������$�Ίp��U�1e��j,��LII��į�g��Q�i�8��駒��K]z��Q����5��(L%/-�GR.@�F�m���`� �y1fЌ����%�����b���R���">|��%��ф�"u��SU,�p_s�}�z?
�*L5����Ox��F$Ä�Q���K("����}��hQn�jg�t�>��/�,����D?G�t��:�M>�>�	�@&����8�E�kjU@��ʪt�����?��hɭ����%���>c�K1y�Y���A0�/�cay(�^����2bg��>H�_{$E���&\�	������_:���O8b�N��8���ϵ�Ʋ�k��zZ�}�[��Vl z�o�T!�k��L+dVIUtn��Eߌ��GyZ7��g�yy�3%|��
)�4Z����c��Dv��}}~����Y�3��;ʭ����6�2��������w���J��&}����3�U8Hr���q(~�CB#"q<���z��҂Az	`��	At�e0H'9]�v�Aw�ތ�P2��_���F�� ���T�!1�����Ŗ&y��h�PMo ����\q��T8�7���m�1Y_7�Ҟ��	�oh��I��g����:��mJ����r�њ�9lO@�i�
UĵL�*�)���mg�P�V�5+p)+�2:x�²������D�x��W�ӳ�EM4��/qc=��,��
e���i1�7g��Ǹ�c��̓��+�=���<������w�_��V�R���R��IQ~��-D�%�C��Zh�h``�h�_%��y�
~�
'��/JD��V#�q�G.屰����)­3�dz'*%c�T�G2�#�Et��k�0ݢ������ľ<?�f.��w����X��|�_A�+5��&�5px�ɏ6I�M߃��T���n�@����u'7��wݚ�/��
'�z>�,2Q���: �l*6_�K$	��D�b;#��w.�oO��/u�U������N�E�4h�d
:��i�%��N�gF�Z�����g�۵�:�5!��/i�⭎�}��DT]���r�#x%UN���$Mz���TN�~ɖ�����	k��Z���E�o�:a���i9*f�;��=.D��n��� :����Bg�p&ö�$����}�ݑl��j��(��>��H��{Z��kRs,nv+��ՙ�d�m���.H��g�SO�������ؓGK� ��%�~���5��P�x��m�!�+�"�ܒ��?���_��m��<ˉ����̊�e)��*�D��21"L�Z��ѾR����k�Co�Ox��Qm�❲�Eo��h+���l���V�
mH���j2�8��o��R ��6��f^8ި��j�{��|��׿˿^������'؍�pb�]x�*Reiv�շ�Z��P���r�w��� ����4;�dz�U}�۰�q jhygJ�	�ܵ��U�꽳�KLu6U��$�Ruh/`�On݉�
�OE�HA��_�
T��ix�';}����"�|�e*�0��P��m��X6��Y%xw|����&͔PW�c\�)J�Uy-��uô�@���m8�f�΋��Jܫx��~���y��xE>ge�x��p����*ʌWz¾(�
IZ��;/R2��U�ٳ�B
�霖��~*��0у,�Q�4�v���0��*��%�T�ㄦ9K)0��MT�1}ګ_n����Lp�t��M5rt��/��[7UE�C��-r�L�l�V���-��W��IV�� S���w��{t֮g:}�:�,���4�ma �>�ʌ"��g�q��c���5�OQU殑{� b%��_���vH��dg���Qǅ�WTR\R'��(¹�'�??�9�$!�$�0z`�N�G��K�L�ѕY���5�%H��C���"p:e�R��c
NȌ4��9��{�]mp3��&`�7^i����jǅY^n`\x�m�j��[[��*�`�#�%`,���wvv�BѣlA]^ܽ�xׇ�|k�H�G�� ��d�C�篤v���AOu&$���bM�nN,�R��a��Q#5��r�T�Q'��S�;���g�#�2>��'���M�Jf��J-B�S��^¥r0oP����@>=r$�3ں*.;�������r,Ϟ=�,�qAz��s_tU�3��#����|���l��BD���l��bZ�`o�S�e/3n���Z�59/m�A zr�"t�xi�pfL�ڟ�q�B��Хw1թەN^<�"L�?�ծ�|Z[LFeaCa6y `�Iu�_=y��= ���6
��.�Z��sR�	�d1teNu�6�~���#d��l/t��"�#���ɇ��m�I���g�H��SJ=�9+�A �t��K�ˉ�H�/������"5ۻ,��gt� �~;������� Wو�y��	_#{��w_�zd��O&��\��@iX։��7>�:3��Gퟙ����kd�\�r�v��OC�k�Cx���!�1�1���0+wa�� 5S�lH��]s~%�@>H����E�8%�'Y�q|�Ǚ�&�?byo�m��ĩl+�LM��v8�nm?�^LL.�31�J��?$d�Aэ�	q�K��ى��Ʋ��sv���w��k��Qϻ��C��B(���zF�j�LW�M�f ��7�u8��o�]��	u���8��tf��;F W�e��>@\R�4	��z(���E+�T���Q����eƢ%�=���`�BPtn�,��B��eMs������C�fI�ДY�F���k	��cn�`0堋���������L����SS�xw3l9>��o�akb���^ A������! �EP]z��幦��(1X9�r�fQ�{�Gk��ϧ
�ɵC���Ď"Ľ�)-��,�Tv��t���vc#p�:}#F�N�诰� q��g����5��|MQ$�
Vǀ<H-�����P]f��'.��V�Ʋٯ���Yp��k}�JY�k��h�ex��?�gk�j)]Y��l�=���Y�+���[s�8�}�2?�=9D,s�hG�>�7F9\V�^�����I�������n��u�oo�����T�-$υ4���0�~�F{h�͵3g���n�M6��F[87Zc� ������'��������qI�ۧAr'T~ע#�C�b�%~I�>�к���ON@���w�S^_�&9�Paa�}�x'�����M��}���+��c�Ssc�G8�S*��O%^=�i+q[��,�Զ=`�p����se5�VHN��a^5<x�hהX�57���3)Is�mTA�,=�X�j����j�1�
ѿ�sY���/�Mn�Dax�,��S�����X��s=� "����m؛�l��[p��կj�H)�2��zj�c���7�|�Ň�%hN�*TNM`����Te����Yv3,�[*0���,�>�bX{�/�W��C�w�︛����v�P��t�����G�Y���E~�T��5�zo�>w�~T� �P̓��wGT��K$ ���lv;sk�"�D%7�(���ӝ�.��rDyI)�oP����L���T������P�@���\(Ƌ�#}�Qw�p*y�wY^�@���m�@(�W�D@{)�H\���r����+%~�>'�8$�Ә	�^��i~�9NBi�J�!{ ߭L�_jÿr�p��T�e	ct ������s��+<�Cx,i�@6�����F����:�����"0y�P��ߙ�\���k�c�h-k��q����'H/pK�H:��t�Q����>�Jv������}�,o�<Q@v�قN(��-dV����#VX:>���{�z��c�D�6hF6#&����T�C��ݡ4�39Oz;T���)�ʉ�m:��!��J�Ȏ��;�]�x��+������%���5�	ҩ����wYט��c1t����q885��X�^'L��w��[5V���KH��7C�(�.^�ɮ�QK���W�۟ܳM����]���9 m�e����(�#&E `t֎#���zS��ʙ�[�lP& ��.!��^ɭ����j(�"nk���5	����|{(��(c���*�rSˡ���=�|� &���K�؏� 2����X1m0���ǽ���im���SOE4������ǘ���	fe0!��"I�59A�X�S��u��R��_��6������-a���Q�<��lm%+&�d�]5'-�D�����k����k���&]uR�tјD�u������g�����GV�[6���9a�B�t�u���I���n���AV���+�z5_΋Qv��K�Y���zF9���Ih�2 {)0[�f��RC���#��Ao�@����x����N�$m�qX��+�������ˆ��!��*�~�E�3fQ���{엒j<�[3٫׽�"G3t~2�]3^�.�6�� ��/:rq�fXڡb?�!�D
f��a�ע�ø��>�����Ax�E�s�0n�_���#�'M��Eτ�QB_� ����"�|Hn��h�R�8$������8]�x��&1����a�mk	j��q��@5��4����;ԩ��]�E��).�K=�W�A�q�<�K��F:
.N֔��r��6��w�!�ǋYظ�D�����L���_�f��-Z��_9��A�\�:rO�
�ʧ%x���ʄ=�n<�b�)b�M${�"ټ���V�����\<�m�Rn�Z�!:�&H`[�`��9���	�HA�C���y 7�2dt3�����.���++�G��"\��=��"ߔK�N�4�HQ����=>�Z2�2
��k�b���U��
�H�c��	�v��Ua�Y+(Yr0Ð	2�lTk�5c�O 7��M����\'2$�K*X��Tj��v2�\�|a�κ澛ox������j�B1ױ�}�s�B��*B�N@�?}�@yֆՠk���b�5<�[yq0�og���1G�����xg��9��>*fG����3�0(8�@���U��Ԧn�LC��	�i���{�~����3�x���po�}f���#�f �=�B�<��d��@8{��9�(��Uܿ�Ց5�����T��f���w��$��������m�$Q���\��a ��o�,1,����s~@��$ ������$�waZyڅ]���6�6@�q���[�}�+��Q���n�8/�5^��M{��\��#݋�j�(>@�6}!���AX�ݧ��_mS���.I�ٝF�'@h�-w+�P.��q�o�m��\�� )�j<į����߅.�~��'����èE�}��� ��I!��P��$�4M�9N�6�C��6Q90J�<���Q�d��s�/��_&�Y�GvlF�����_s�ݠ*4n�MS�oij^�������F#V/��ؓR�E���F!I����ʮ��;ҊB-��S�o��+/���!������U_����@:S��:�m\*|�&�O��s7����u��=gxV���͛� "��V���X�$�RV��`�M�ڟ�ov,{��0O�>��z�-��K�H��"�2d]�,�!L.�u���=߫#"���I�`Q�<�<eVNI!�����=�� �$���Ε0�t�=��Bꉬ�e	����O�{��a�dZf
@9��F0O=��]1̾^t���Q�,�@����;�# K������?�n�'3�㧘���l��(鍗�{7Fԣ�PX�$K�Ph�ɖY�m0gW�j�E���h$"�!�g"���;�i��CI�+�[����=��u�2\k<I�ǻ���\�b���:$�D*9��(�(��B0�D�(�{��i�x��7%D���w�����3�`3���Z�1��n�M��T#WO�@�%�l/���ToIO����b�P��k�UP�8��Э�g��XV�F�ƍ�f�~�r�}�<-�W�������X�w��u�%Vt�w3����)�ج �0Уg{?0x��i�?���_�w��_�#�NT[��J��s�lۣ������0W7=rb�]<rUm�$*_皌�V�q��"��?9j�dؿL`zv�/z�r���``����Mk�vh��W����Hk��a͜��o	+}1 �G��"ە���Q���E�I�˹�A�t��b��K�ٟ%������0�5�,��,,v���7�UP�5h�b6"Ռ�f�^z�f&�Ij�^�&����4́�<tE��ei�7c��^f5K�}i~� ���������K)$��+5ܝ�a�A�h6&)<uZoD	O�R��ò�P���R�c��3-��=�?�(c�^LB��`s�� ��f=�Qk���o&ލ�������}��M_�v�V�po��c�������Zv]��o2�|�!<�OB��R��у(�Caxl@�3�� ��_^ cg�s�#j��m	��d��~��2�	����\�h�>u y*�� ��	)����Jpgȴ X����'��HP�%�!j؊��O�'��e�jA̿�L����yqm'=A��U-��Xi��pϕ�u�yXf�ųž1�,kP�޻w4� h����B�9���銮���@���}w\��F �_�\������~����I"p���[/V�����/�0��NN�>�T��w3�ש�bӴL���n���(������B����0�'�z���La<�IZp���u�q�w����3x�2A'�L�����L<b���⧘d�Ls%<�M�ہ�oQ�����c_)��G�j�����h�����S�ڶp��B���+Y�0�Ix7{�D}�����>�!z�Z��7��xDH è7���n�ڦhZ�+����1J����X�mY'�h������v���ĺ	�f��
 �� ��!�K��t���n��t���������)�����������P\��U.���7e������J�5�M��y�p�.��|�7�I���8!��2)�� ��)1�{Qa�3nB�<?i<rZ\�!�ȗ�����i1c5��D��W�qs�n�e�)6��T�~G� 
X�4{��ǃfM���)��� �*��#�t�r� �"�����R�l�q���6ǮT�xS��0Sn��C�|���|m;Ml�T�����LJ��(y$� p�\����I�8Ժ��Dسm���n�z���B��vcB%�=�m�2��}U�y�K�v���GK�iWpmP�'#Y�Da?`�I��k�=�'a�q tm�\�����p�DA!�d��L��3��/���	r��F�l�eP'A�����*}� ,�ל�Q��[���}�Z��K�5�u�ܾ7��e܂�u_|e�����"��t�JJ�G2^q~�_��P|�c�^�-�4�y�"='v,e��PORչ���R�6�Ðǉҟ�j�_8O����{�~�lwR����~�2�r��G)L�lr�s�]����i������i<���~9��|�,^UZ�hmjqT�*�O �\樬Ë$�H�s2Mφ�@Y6eD���0�1�����F`�g�ߊ��_�0p�I3Z<r�V�i�:�
E7��:��6"L�a�wtpoZ!��Fr,���RA\�U���vUj�#l3i��u,;��dB���+�"�����ZV���6X��b�PR�S���azc0Ckj5U�t5z^�R�����?>�Qi[Q3�p7��|y�:2�Q�5�7m<^�r(��p�lNCwQ[��8Z�4������pɘc|� J�&qڕ��Z+\�ߡ���P�7�1��g\ɤ~׻�/������`%胿2��ض�Ѣ�'(�N;�qa|�[RH=�a0r��xf�T�b	�2�^�����h�ݟ�9w��E���M�1^��܁~��/�MZڸt7���/�|&6-�)gnf��Kk����[/Y׶/`��;�g>qƶ?/LJjG`n��AqO���p�I�M&�%�AG(�F����+ND���~:G �M��K	�Æ�;��"U|I��.�>��՟H)a䷩��C�Y
[W5�a�nPC�י�E'Vas�]Ȅk�(�˔_zx_��FN�`O��o��PesP���`�b��N��͛�����d��(�&��xK���n��Cצ�J�����P`�KŒ�h�HN�l�4xv�L>�<i;��7�z��
c�ҐVU~��Y�\�l@(T�
ƾ�c��8�n9۰+v��#�;�Ev�B�&�����P�޿``G�=&��� ��Q��[μ�j��ȓ��j���
J�o�J�K�>�s����j#F@��@U���hK 2�+Q�m_uR�-�	9�-�;�{��#�V�?
��
���-U��Օ��eG(y�s���-�>��)�P�S���������qd�Թ����+3U򾮾�c��Uc�.751h�}�7v�}�VK-Itg����!�x���C�ی-=�a����-D5d2Mv��E�.�-VP��Ä�?������RMtANh(Z%�����P�g�8r{h���L�\.E�|��6.�	R�B����C�{&���,�r+q7O�$���,OH_��D��	3��V[�&9�̺;\,h#(bS�_ݷ{T���]�Iyd_9+���^R<� 2:�*͒�y���0*Nysy1��c��!;=���qj���O��X.ݏx�1���&���������uv��&�1%�j!rƍ<�'�`�n�{�� ���K�B�GU����t�K�/��6y���si��ڧr2;z�1>�"�FJ�x��Ũ���U�s��Wpr��z.o���r:Dk�6Y�j7�́�q�T@vl�
�4��(;�c#��LT�g ��,�=v