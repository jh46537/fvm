��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7Ɋx�!�g���I'k�c�Jӳ�xz�:�-94Q�߼<p�bj��vC7$=��ȭ�B�z��'4��PNGw]C�����贶���hK�e5^Q�uP��(�ӕ0k����ru��5��]W��!�aI81P��ĝ9�T+�����m����X7��f�y�pK�	#&��t�Pw;�UI`�*�ӻ�����X�͕V�KWn�c���nqMF����n����,�z�ը�Hd �q���T����8S R����Yp!_�y�}�C~��k7��Œn�,d���ݽ޺C���G̛e6�j��l:�ݹ�~����<ƌ��@D0H:���E����I* 8ZBh�_jK�jҦ=�Rl�I*�f�8�O�u�q��B�@�`�����Q�~t�S�#*�ىA��1S�T�e��Ň��Fd1���3d0 �}�f����q-��L?UT����umn͔�+5���BE�~���CC¥��K��u�t�[�@���+_�\�߈O�L�
��G������=�c3>���O��d��� �u(�IJ��-<0�K���Z����C2�gc�җ��G����\ _���|�8�AK�x频�= 4��	�S�ly���ʮ2�y_���Tl#���ʼ4W���+2����W��&�)C�YT@X6��3ןxm�g��>Y��*���f��j|Ū.b����B	��C��YJ4M�~-��e�g�f��
Z���C��:4���V_1%%5�^�y�g�nU�OC_.K!ln�'��&��I����K= ��ʿB�O��毩Î�	�24�A��S���8V��=x;�zO��(�1DI���_�����;��Nz��ܛ���xN�L&�q\������W��%�-�F��>����b�y["&|K��?�T���(�(�$��	��Z�ɒu��4/�U��%̴0�lع�mS��)�:��k��C ���hQ)!�"%b���|7_ _%�!n�Qх�Yy;�i2� ��Lnvw`]oi�䉴�#:G��&>���%t��H>k��8� ��Mj_t�i����yx�Д�f��Vk߯bQ�<�S`�X�RY�Ӳ��2�s$S�����_&cukD�v�P ��K���G����;�S�UM:)�1���m�*|1z�Ede0� ��_F��#z�{�3R4�}I_SAdۃ�7��>-�0�7�>ɤ�r��,A�X?a�b�H^�J�����*cAo�V;�K곭�`�f�3^p���Bz!��z>��O�0S���R�ygS�Ӟ�Y8q`]����VȦŌ�nd=ʡ�;��L&G,���R�8�R6��Ϋ��<D �b8~������sַir��En+�jO�o��x��zE(p%�(��v��
�>:���=��mL�~tC�jL�ګ��Ԇ�A�ɠ�m�A�G�ڬ�>+�?�l�)[���E���q���Epv��l������?��@13�jI/Ԇ�3������C�����`��Y���` AYrCe�g�v���/��3^02��:4������sz�<=�����N~\^��F��v�yW ���Jf��F�����h[Vމ�t��^���,��.�et��������ᰕ=?�+�<����n/�)�+����fp��懞�MZ�_���4�����9��I�m�`��oKF$��bWG�Y���a��G��Y�Y"1�ͣ#��d�!����{�O8�ۗ�cID�r�V�o���#���փxfq%8K�:d�%�O����/r�o}����,9t�� >��JTȱ���6B��J�|��I�&��v�ȳ���������=�k='aݍq�6|�:�ɷ���0d�6"x��r\�z�_4N�a��Ta�:�9��jg�V7�z�m��(T�U[ۃn�2��u�oۘ�Ҹ��R0�w��TS;tƸ~�&4��3���P	qg�(���o��t�D_��4t��<TlvA���t�Č�(��Mً�������vtj�Z#�ܴm�0S���$s�׆'U�O�+
�<k
�ƈ0��8�]���D>���|+i�`K�Dl��N�b�ͦ��j�;��g�f���o�Wbbŝ1�``�"N�x�@�V�2/�Hf�|9�.T��.���9���3���&D��4�A>;U�ܙ�h�B�"��&�:�k�|҆\m֓7�[����ɾrɬm��x�u"��C�2����� #E�*[�q4�1ʌ+Aim���i����6F\.�!�;\���F}�ܾ5lY���P��@�8 t�Z��ʒg�7������fl�vI�,��@s���9�����&@�����_J�,q2���:|۾A;��;v�=x��ȳ<c
m��s���&-O�)bTp�{4�*�K���=��&/.��/�#�1�*H&Z�Y���j_O7V���}3E9���C���ƀ�ZH�܋.G�?F��xLz��Y��Je�(��P�KJ�}+1�����kNֳ%d���n$��ǆ���G|̯Z]�O��@���)<oR�T���OG�xi �qlD�}>ݓ��q�VM%�i�x��qapf&�{�������6fZ�Q��o1�"�h,�ရ�1�Ű
+��>k���D��>cC����F��#�ųb��9Ҿڴ��F�>ck��9ޱx����?,�E�4�*�����"��F`S��?����c�%�����V<���+���n�C�%��uy]�9Xq�:t ?n�<�@�� P3ӷ}��DX�F4R���ciJ�y/eO1ycyS9$�ZיT츭�+�V�ci�Fդ��]�����Kk)��58[<��a#���E�`(�2��`��E�(�e��e���6t�_��/}�	�O؄�:��<�I��%4����#)��eU�p`H����au���(S�h�{C�hΖD���}e�Ѽ�۵�\g"09s�������Q�k��A��Nt�G X�����$�[�և�6��0I����G���;&&ʤdH̑^H}B�~h�[�Qlނ�"4�L|0�cM�:kb��B�=O;i}J!��*B�~�q @́4I�e9�i�n,�_�؞�'�DC
ųp,9AC`�A^�Hl��R�`훬�Q���"����7A�{�+'[5��0-��W���n�nؾ��UoX�
	�&��<�8rQޅЋNl	���d)�����̛Y�x��T�"y~=�vŽ��>7	;�>�jw��'�������GK��qk1�G޶�����D޽�g�4�կ {U��oY98L���^�g~|��Tg�ۘj��qb3��S����N�)�+��:�?�u�7����]b1wD��$o�J��T|��I��U�L�t�.eE�͝��ppu�ùA��ԃ���	o����K��U+�a�崈�ҿb��$5~F[��B����R�)9�14	w&	�)�٦���p�G��'��ϡ�Ě����+A�7	f��9@�H����G
�D�f,��R2�+ה?:Z�L�/���p�����z`�[�#FҶ���(#��V͖ф���U���H��
�~���,O>?�m�Wd��oE�1�OB&�>����XR�ك���4T�l��ڿ��.��.$P�>�_�o[��*u��p���Hh¬�E��G�x�'E,��2�kr{�+n,���}*�	�u� �}����`�]��Y?fxsF�����f����2�ڌ�x��������-��~64�o���X��O��f;5�^j{q�Q�jnhz����̤���V��J�x894���5_=�e�T,�]d�^ �#Cm�#��:;������}�U��'"�R?��(�$�U!Q�Z����X��8M�����?i+;����_h��c�=�l.C[���Ȗ���O���K���>�������������qoW�A�7^����U�ۙ�U%Ք����b�CF�ìL�>���5Cy��¿�`��B2L�u��4b�`(����:7�TB���ͫ��`�9޾ȲM�l��r��J�U��Te��-X�Jcg(��m�O���,8�yY���Dό�_� ŪG��V'kZ�����5Ҽ�A��7�`��i��Ѳ�t�0��R��PF����[�c�A�ҭh�Ö�v�5����ia��t�S	�Q 0i��I)�	��f�Բ�tϭ<��н���3��I[�k�蹗t���gK���=tS,���� x�ւ����&�0����$WNc�?%A�^��9�:(ܞג������7��>�{D����#X���W�i����[���?��D:a���׋�Owy�����"�a�a�́�Q���Q����f���_�j����z��s��� �j��e�T�[�Z�|'E	��^�.�xnպu+�B�����|k!�}�3�%)|o.{6԰	h����lzq�ئH���Y{b7�B(���D��"c&�D�K�i67�!A��T��6v�,�iه��*%/�gmV.�G)Q��}�?;p�K�k�����v���0iA�7���v�c�@}U��?]��¥�'�tk�����`�{Y��1S��<��7��~R���@��B���r\��|��KĎ�
*+b�X���8�M!v] !r���~�U�)dY�]�%���̗8���T�q>�N�i��&���ٵ,M�F�~BU'��yٓy��4�5�+��UfR��7�[�X�(�5��@��{��>;�޻%_5�Fe�R����`|��ɛ�M��IAwE�i>R���Q!�J6A�aIYy���>�Ė��o=[҅t:��� �6Y.O��M3}dSj��vO�k��1��5L\�Jq!��)�	S�֭�
�R�f��,�o�X�s
���LjN�,�@�:���dp Īe�u���a�ӛ���/i�(۲����*O�*|7��eA5+WN5���L.�����4�E���ح�e�~��L8vUv�P�B�#sh��J�Vk��AY圿�Y�s�ɚY���&��OP����/��Ҳ=�s<�����>�'�!Q��㺰[&�Ed^Mh��ܙA� 2��h@�B���Y��l��d���V��!H�� ���2�o�D�!��u�t1�TH��6�a��F�6�3V�BT �ʪ�(L���_�!uO1Xɸס��	� ��������ٕ yH�=ڟ���MM���W��d����E֜]����ҿ�9�[�����ȱ�ۡ�s[�$!�%��������J��\�J���̃�@?�c�$˛��4 �{�B��AP���_6#9p�u���ƣ:|v]ak�K��H"���}�L"�s��Ґ��.�M�٣lq*c�E�`j�lȉ@��ܞ��>���=���Z�#y$���/o�G�u����ȉ5�	�94�O��_���kHۼӎ��<�hb-���Ϯ0��X�P�2�>ۯ'X_�����1����X�o�����x����A��*��v�ۀ��	���~MuJFX��u��6������r-ޠ�	9`�Х9]�Ϡ7��D�~l�-uO�^��gH*�ϮU_6B��[��@8��D��� ���i�"���g��b�^�Oy69y�&�f|�W��u�dP`�4�ȹ�68�0�X'���¦=��[%Ƶ��=�}��i�>(�C�|#�s��s���:�^�X��k����1-D	��sϬ����QՅ���������1R�;�B�\z�̸3��Zi���3���q�����B�8�O`���4�7PB�h��8� ���Vި��y{;���0��i4�=�D6]���/g�1Uz�w;�8�.���{��i����l5��C������sؑ��O� �TVE���y5��<D[3z=�<d [
6�*�ME�e�Ǜ!Pм!�C��_��(%��5�I���0��z�^���e �k�u�6����=)6���iəy(�x���̠�o�����}u�DL��O�e|���#�]��i�~�9�JwH��K�=�CAR��c<�bW���F��a|$��TT�Wy%b
E$*�;6b-/�E8�_^��J_bZ�$jࢨ�$��G��H|{+��Q�����E4�{8q��]�8�R�(7�7w.m>�����uWˋ�D�p5�����8�ɓ,���f�"I�F�A�r�{�I���0Dvsc�SL�(��y����4���/��]��8�P3�-�������¨��B+:v�ѿ�i])z0u��b��=�&twB1Ft���K���C�V�[]}�QY�@�C��t��x��������^�!kp�Sj4����I�`G���q�U�zo&�I��9�}��J92��t"NMn�)����؋�A� 9g��_�[��&}�F�%�V���|��9�ؗ^j���<5�I�� ��X�ͤ��v��5�90��1F`Y�ƣ������}&�˼���:�K�Ǯ���-�"#�Q>7�Ȉj� ��}$nnl�̬��8�������t����5�*��V��H�b��qg>�ćLu{�Zo*25g��	�Q�;�)$�E\C�e�-�E��r��S{jns��J$����{i�� �C��K(��ܷ��<�m�\/	�~�j��؜���o�Q}Q��.�&B�sԊ�>_�K��b�]Rw��y?储������=��t����s	@�T 
Sŀ��[����C���n�
���0�r�����p-�?k�S.6{D.,⚄��](v��BԈp������O�v��>$�x��d�M�9n?��!Zΰt�&���h���boT�s^��{��(�Af�(�#�oZƄ<^v��}���C&��PJpHɄF�)����[���r�����N5udC(��`�������B�N��B�.#��j.�`�'�?&gj03��$�e�|;l=�+ҋ���۴��(���;g���)���(t�|HO��L ^�rs.:Y=�Τ��_��$ �[|�җ5�E� QE��2������`u�zzz����8!D��( �����x*�����D��X̠�� �qW@�^UR�(���p^�y�،�~w@��z�4?��iN�ϻ��]n�@�	w�Lӵ���a�J�uB��&S	�ן�PՃV�:އ�Tl��
�]!��9�R�R���r������`��6��p�b>M��1���]�a�����O��?mU%.q �CE�-��:�1v]�?�̘�+;V���u�@=in��m�j0hʕ�� ��]�|[��Π�mNKHw�[_g���l��F��\HČ���X�G��@���I6F�Ю�:E��ձ�Д����>"6���ӱږ%>D�_�zm-�a�(��5�����m�������,��X;:@(07�c�Z�t杗�����ɽꗣ�C���ҕD�<Y;
噭i��/K�.8n�O��� �!4XI�2&�� &��[�gy�����V���&׆<cC�*��^��=HZ�(�k�+���D���)XRy�<��8$w�#�Y�;��h� �#L������75�6X��iЅ*�Khz��U6�c��iWst���c=��Oͻ|�JIH�WN����ޭr�W�Ј'���Qo����K?�̱����Κ�C[2j����kZ25$9��1��jtjÆ���]�W�g�M��e�|�G���8��:,���dTfL��0L;M�F�Qf�����69������>$��o���<���)qm�&����Qi46Hy��z�΢i���uSm!R���JXj�<��q�v������ڄ�Cn��Y�]9���t���{V�m!�|��0�ܬ~N��!�"����#`9ZQ
N��Ȋ�����r�����M�ys6�\˥0�6���\���4�5����ٔ�������Y��axJ���/�zcm�����S4h>�y(�X��]cyX�ڼvNT8c��(���\9�"]{���S�s�X�Z�bf����+^�3��e��Q�|�͍�b~��ޔM�[!v5PR%��$֙���Q����)�'=�uSs+3*/�4��ښ�A�����}�Λ�aM�n,G��9 �W�Q�۪!�����R��d\~9������ߟ����xi�;0�%�ýԲ��r���=1Duk���BO����-|�f��S�As��wp���~pg�&$��M�m$��EiA��>7*,(d�����N#g2H�P>|�a�����S���X��1fr��c�xf�6.��*~Rr�K�xqm�q>���ܼA��_�$Tl�d��#���E�8�Q��T�i�P���=�񎁭����tC�k����/��m�==����@lW�ޟ�ԢA��e2V.�LL��<>�=���n��/{�� ���UH�8��&�E%�k�N�_���u��@��d�)���q<Z-:Ī��� ��름���E���KC���`�Ҿex���W��߫rwo�}�\*��z�]r y��x9)� �'�s�.�U�w8�p �t����ެ´L*�D�o�ߛ��;�'��B���F�M"��������DVKY�0�[0��^y��ma�c]��3�S��H<�R����}��U���z��H*HLjo�I)fr�0*͗��x3p�lG�g����!��82.I�s)�2K?,
���<L��u�f|��>*���EJ^|����t�c9���ߨ&�A$���Q� ���|L�XF��~ ��-��,�(����m��թ�ny�v�\VER4*|��3i���<�V�9	�*��fm���޴��!�����I�lOh�c�_k�-T����2yJ�JM�S��Q3W��H�Z�#GaҒ���/�
93��]�	�\�އ�<>%u�(�8��{LO��
�O���O��.Z���[���΄�ЯO���l~���KT��m�J��O�^8� �=U�Ր��mW�O�ȷ�G�ۖ�7|����oQ�I�f��g;o���f���W��1����4��6�@{���<۾`�������i;h*}׍E�4��"���S�V����w��U|�[r������Iu�[�k�-��a@qr'[�.�~��Ǭ>���r]U��}�F�U���!����j/w�IӮ��N���}ܻ�PM�5���G4Lh�j�g���l�j�����jY��<�%l�d�w�)d������-0ܺ�|�DfW��O���ɜ������Ȑ���Im�I���R�7�?قk��Z_�W�wZeb%�Ƌ�"I���Z�Nn+#�ͪ�s��p��B�����+�N��k�mA`S�<^r6ݎ���I�]��6��Y0���c&VR{F�ù��Q���Hy�s�y�?~8	#�.�;ʥ�������,�������=5��Ó�B�|��Qk<�1[�8�]��7
�l�\�|�ӗ�/�uc��]���K��q@f �e�{p�e�<YI�-2������-�`���b�a��[�*�~��$Jn���W2ٽf)��2��,�|5!d�5��S�t��٭`��(&�:���M,����g��$���U%��aY��2+��3�"�7�ؓL�0��پ6.��K�pZ�U�ةwfz�Z�w���^
�"��m��Vs����$�21�%6�6���Sŗ/����ӯ/�r2N��`����w������H��M����m��!�m+�7�P2:!���uM�6��D�@��o}cn$G�biJ?�1!�����U�����L����Ѽ]�d��:��0%t�6���{������B�&�d�� i0�%�^=�c�v�,i^?{xv�pv��j�[��}z�I�L?���]!����ɇ?�&�`3qr��c��L�S���k�_�>̇a�j��IT9K!�������>I8��҈�-׈�#\��|'_����Vv�$�-B��)�+��f;���4D��׏b[F�M�-���F!5O�A���d���>Z7�Ra��i��8	�%�8��rP�jY����15�w.��>�Y���O�m�>{]��qN���%� &q�o�Q��x	��p���D�"(S�r��OK�mO&XC/�χ�o�a�E�����'�3V�o�zǥc��1���T=t�XI��}�]�ؽ�-jE0��@�BhMO+���D�_��G���Dr]��qf�8��@
�?L�`FzQj*֕��A?��P/v���q�%�k��2�@YXy�T�_bX��4���^�c��2bK���$]#Z�F��Szw�,�e�,���<֫?�p�=.Xv�9tX%aHN�7y}���1ʱ�2�K@���Ԗ��Z����G�+@d�J1Ԓ��Zك�$�n��*�s�l�G1�"���Z�����x���M6�L�\�D��i�;�����E7��UH�[��>���\c�L"�>;��)��d�pSo��y�>��X�bl�d Q�S��E*�Zl�ۿm3�n*O�#7�Ϧ�x֦� ���
M�I�G+w>���,�5��֎d4�nxKC�/�2/0��g|��N+,rq��Qg�~�$��O�!�]��}���`I���� A/���e$fۙ�c��M�L�\'ե��5�6>�7����"�B�)�C��08y�9\ٰ:H�/�l�$����hU�y��a�yZaպ-}���Ǡ$��:�7xj���BK\,�q�?d��hk�h��قJ+K��v�; 2����-�Ff�D��+�*�oS�!)���_��@ԗhU(L�#���������<���O��4ѝ����Xֲ�m���pD-��lf�ݔL�"�1�u)i��.�B��r��ǜ�l�6UPT���6o;y�|75R�u�@@����>[����RΈ��p(��t�!���¡�>�O���dݜ^���=����F^��`Tެ��Z��B�I�\ݯE�nI޴��	���Ϫi��3��S���	�xO�f��{N����+�k�����'���+���ru��O;V��T���B�P�m�5ͭJ�����������~gcH��S��[��uޚ4��D�������R^�d���zC���_nH6�k�bY�QU&����h�Ң���P��R�DB��-��p�)����u�֝fj�K�x(z��+E�0��9��~x�;���{Ɗ���_B�"6�Xa�^��꠱I��n@2�~b=`P���:xDvs�J&��QX�
:�.u�Jݞ=�%�]�i�+�B�y��$yN��i4�d��6(��O$�RG|�(jq��~�b`���t�>�5�(�g��YlI�"-�����!ז�ZG7�3N����}�iB�����W�.�y%:;�ʵ<7�	7�Rf�1?׳�p��?�(�X�;�D�ƽ\��&��H�I�O�Jf�i�K�{"6��gDT^���"���E��Mhb�J�fJ����Io�s��Mno�D�t��N�R�):�O��x=�\Pl�Θ�s$��Z�^��q�b�uf<"���^�?��~��1��a�����II��)CJKp��ͩ����|0S^�H�hM�u��_k�c!^�u��A���_t��je��w+�y̌�j]s�=5u�����6��������~97C���lhǍ��ob�~Qh�L���9��T4ʵ��Hª��}�������1:33,�vrs��M|]�5g��Ԥ����ٽY}�]R��&���Y�޵������p�f��ďT�\�]��ڞ{9�	�
w6�ίQ�T�m�.�r��8ʉ΀�E�gg����1>�]h}獥����e��V�F�t;,��w!��Z\G~�P�~���#}>���Ap,6@��Z���d�����l�B��b��zxy\��c0N�@����. d�2����ٛ~��hFQ.ġZ�
�^��;a_w\8W���ɶA5n(�K\sY�RF�3���|&AST��6��`���%x����Y*�3��\T�z�a���7C���@�>8{����	&2����O����=�	6��å.��M�
��<���x�M��֍ᤪ�4��.ё�I<Rc,�+O��:�h\�?���M���Nj�yLev��Is�#z�;�J�N�	]k���zAIr��{�����d������F����(��� M���9)6��2i��W��`���T2q@N�Th�R;7!#r�xγ��Gރ�e#i��ZЩ�V�iO~x����b}v��␏f�oJ;�l�\��;J\�o�A;dq�?����= \}Ą���n�fD�qތ��b7俄�K��n,x�u2�R�Je�K�\��/a�Ȇ��J�Y��㟩LyCxT��8R���nD�7�R04b�;w�FG��rw7p��5�?9����-�5�O� ����>�;��_ǖM��׽-r}Z�*�,G��R�jm�<�@�1)<����]�����P͹y�����QEeg/D(S�BkC(!�+C���uA��@��`91�K���M]%���'٫�:q��,�N�_�����2��ɺ��	Bcdw,�f��J�
�} ��a�p(B��� ���2�����)FJ�"ET��I� #����"�bߑE@[e�C����OU�^��m��u�/�Б6�dF�-�n"�BǠ�Gӊ8x���#���X�)��o����;��5��@I�lM�s�Ռׁ�I{�"�kY����m!?���٦�L(<��R�!���^��gÜ�F%��|�jB�3��G0x��F�!�\��P�8z���
��Σ�̨p<-.e�b��1a.��4�D:��0��/E�u�2A~V��H�u|�����|q�\n�t���q�Jqy��n�A����j�)VA�f��BLb����#~rS�C�X���������v)�R��r�����"�t<	�;�"[:ӏ�u�Is�h~���׀k %�3����=bw��,�ؐ��<��SoI���ܢ�j�jogCK:�@�'!���oѥ{��5mo6"�)�����~�'^��H�r���i�R��$dJ�I5{'K.ѕ�=�>g�P2I�DFZ$s���'�[���<��XU��G���YWB�ǥ��٭��O�.S�p��Ib�s��2������.OȌq��)VywVK=?7A�j�����=�����ث'B���l�L�@}�2��;H�y@�r��F�	
0N�ї����u���1�0��Ϙ����%U����v�Z���Ng-s�6�����o#������t3��4N���$�Z�\�9/�)��I��[�"S��kB�-��͠�e�<$
����k7�T����l�!�N���Ki��������t� �#����s���9(V�6�@ WcO�`�ZF�d��9�#TJk�
����儞!<���IU(*�t���#�8�d!N�D��D[^�*5{�)���T����r�	H-��Tj�~*&ƙ$=����ư:�ў��V���$<f�����uj$]���<D g�h�|��]�Qb��i�% ��QJd��� (����#�c�$	�o��b�q��}�#4+"��uqo�]�n �Zro�σ6
#�	�d����{q���2-� "6?ˠ���s�6R25׼�	���_R�C/"y��\-ˣy�����P�*�� ^V@�Z ��}�Ӵ�h5	T-x���8/����[����?>��]`�"����8�3����ͺFo2�$�J���K��:2�N���*���j�e�C��FAF-�;��;9Q֖��O��V��3�f� ��{���l�l.��+79�W�R%'�]3�.��jՀf�ϙ�����տz	���bΙ��P�{�D���{�w"�X��sm��B[��B�{"���	 JFҲ��Pj!#��n[ag)�`�ی�Ǝe����]
G?J?nq�>Ï�{<EI~*���\u]��B_����#L�`�,-tev"-r���Gb�Ԣ��z�����Oч-f�P�f�׸�a�`n�R CG��rng�x���yKThy�n�+�ֲdhz^A	�������c����ۆиp�nhӜJy�"��̍uN��3�]���tJe���gҩ��E!Ok�l�@5��I�߸8	��cX��͛���P'�K~[é�B�(��U��ϙ�����$|�����i�4�d¾���_�A�ӫ������#P�6���tol5}@g��-��	��e��������5�sH�����P��1Ƅ�CS[Z��xX��-�@i��8�p>O4���2e�4ZS���:��g[i��3�,��� �R���-�^��eU�*ul?�)-^��cXWSK=�d|g�k0�>6p�޶.me�c�oW���`Ѵ��R�����e�El�(X�C0�͹��	���m�#t w�Zp�aa�[&c#]���ȝ����$;^�YGU��E"�� �N���s0��2/��	�|kd�|�<0��B<[��°�ā�@�o���L�3� ���.�@M���b����a[����=�X��A�"yj�6�X�+�⧵x���rp$�*�W z�� ʜ��~�3�K���A�~��������q�`"|�FӒ�׌ �$hː�8�4�l��#����X��@��6�͆0_��UcM�(ſ���a{Y��ٜ>��P�kk;�^6�������~�i�G�7;����DuP����q�'�����G/�������@����=���3H�+_B�"	�#�J�p�,HD��_A���j�4؝gXR���� ��������T뷎��A��3����R���A��U�&�0�DTk��F�u�Ȼ��x��������t�r&��)Ve�2�o	w3�����(�D����@������Qĕ�O�x�V��zO!Ű���y<Z��O��=����e ��VTy"��y� ��KiΒ��ҽ�b���<br ��S�E���lO���,Ă8��z���'��p�i��h�>hY�/1]���F�>����iB,R����Oz^Gf��k��K��nT�>���� ��Y��zEc��G ��},74��\�;X��m��g�e
����Q�/.�:G.#�yP&, �FB��K�.ǎ��v�k?��N�v�^��5AϮ�Ш�~O9�VAYr�s�X��*��j�ٗu���ڢ �v�cjxF���x�L椦Φ���wE�;kLg�O�GhI�]E�̍m0���P��a��S{Ӑ{�nbm�Q��R�O�s��Gt�Z�a�^��Gyn#��{���JF#��hS SpG˯���}��h�LK�_W��a�`�&���|��[SV|���m�]�̥11!+mH�;B�,q�z\��M�n�u-ٺ�L�=%O��(��eژq�6�,��	�k��`�G�j/�qY�f�$&�H�xM�M�_d
�o!�ł�����N6��	L�z��R���ux#?�&MY{\s��/�Vu쭒��L-NCpb�׆������6��H,U�@
����.#��u��N�JH�]�8P�b,�v:B*��n0����EEP͘�낷`�M�Iէ�6�X���c�����CP�1vܕs��m��oyp.q049ͼ�d��X%ْj�j`�S">0�Tr��K��#����ӻ()��ۅ@�ͮr?Q�z�E��+��l��P���w�@cfA�<�<E͈�?T@&E�Q쵥z(�8�އ�>���Tӊ��uJ��|kmg���U���sH&sȸ�YY^b�O�#���R'��"»��Z�V8]�Z�#L�+�����B	}Cm�cco���8x����b�Z�c�E%�$a�4��>bnW��h�7&jV���X<�y�繲Nv��!< ��vA�Q�4�(
�����!�h�-B'�:��av��|0���d^�u8��U�$ԁ�f����)¾h�8���Qwa��0��������A5���7�����[��	8��IV���
�|�U.������T{J����"������XɰT�M��@K�f6�P���/�8�M��A��C��Һ��9l2�%����4��d{����R��� ً�{���mW�X���R�A­�q>��\����x�|��!IG\xg�'�F���7�S����a���5i2�	��U�Yp��7%�vȈ���<:KVb��e�7��K!;�Ԋ΀����Mծ���_����T�to�}�⥥��� ìv��cs�ۄ!�J#�_�n�@�b3�0�3ﺳx,�g_C�5�sc���u��.�M_̈h�3�|\}�7���/ra;�YR�Z���w*ۏ.�a��h���Wo�x\Ì�ꌖ�_ �O��9�w���C�M�#hu���=(}?Գ��� �i6�%��$�)wFa�(8RO��*����[�2Ri����<�M��pV���%�I\��>|�-����qҼ�d��y�+�8��",os L��d�<�.U�b���<B@l���YD�0PAa0b�`����w���H�������8M��oȿ��29�6X���~��0�6�;��?n�4`��[J�!n֟ze
3�Z�C�J��UJ�~57~� �dߦqH(����U1r�n�wxٛ~�� �#W��Ʒg:!L{dU *�>)ed��_�IYk��)�j"�;�ܑ���*H�L�?D1�:Ď�-h]���)��[��ZcS�Wd���©j�ϡ^	&�ZQ���8��Ȱ�'F�����B��_]�1�僯�ozvϝ�e޹��49�}�Z���_{��0\_���Pm<Ӽ�����������^l]��W�j�_��246�T�Mp`��x͵��d/��}Zz�-̸W.֋5�S�Zc������C_�W��R9��6
���E���*���9fSb��,��XV�g��7*��A�k�'!�'����)�٦�:o�:��b����YL �B�#�[��N���3$_���g��'�9j`=�y`_]�?&�N�C��Φ|�&i�f��S�gF�oWZ���&4���\���h�.�;[�΢��BUTz.�ur���s ���	pc�khz�̞?��d���Rx˧~�SV?	�V3~?te!����b-�Z��j�,����ʀ C�|��p�8s����g�c�QtJzW*g����EQ�M�UU��v[�]��yLӳ����WV�$[�q,E���+�z��()�?&=�Yf��v	�D���$Lv�%rh��Р<D�K�^��q����
W�zAP�E���
����l�3����}_-l�����s�k|S����R�����O���4̓��h�q,���k�m�!�A1�FAS��_�{�ߛm_�>Yok�6���2uR�t��0��&����,�H��v�۳r�Դ�%1���1��2��5D���� w����a�g�/�H���|�	4��>�"Jx|Á��oy7����
@!�ݒS�qJ����ĭC;t~�������F�(��ߐ��}T��:�ά�np¥�BD������!���:�7E�3��1�Ay�0�Ms ���ɹD{"���(�7.H
Ť�N�sYX��a�L��"x'�n�t$A`�������#���SC��� W�XH�k+�G�&����%�T�<���e�`�$⿷�$�t��ZA?�����o s��#5�q!�uG����>����c{�B�+yi��a3K�Q
CN4-f�(�t*q�"�wTj_.]�[p�5�6s�w��ޖnv��)��`���8���z����qK��}���c�|2b�S{�
^���ySO�N�����w֝G"�e�!���;ط_eS����s�������+���:�:����3�\���-�{�B�����W�!!�@�*��&�!�Ƀ%��(:A�@��r�0ʹ�*�-�]�L�W5]�`�>�AF��/,�Z&��� ���|%�գ��	�����g$�� �5��H��z�ҥe�SҲ� 1���$�
��,�S���1i5�H�A\� �*�>����-�2��Z1b��,I=	�ݧ�Ʈ�-�	���	U �j��l�p^@�l��8`� d��Ꝼ{/�{+ր��� )\ ��
�V>k`{���~���ئ��
N\��A��M:�[	��}G�YVᄿ�K�������+R+9�|0�cs��&��Hi����}჏��_� ؤ�$����K�o��I[����۹)�1v
X��_���R�)��ݼ(E*U{����7�7#N�=��X�T�(��J�U~�ȝB�,���UQ��=Q�}�a��mi(��I���ꀤ��/̰����9:����^�����p-��QhU??R�g
�É/��}A���S���07`�A��7J>e6����ag�V�v���i(5X�a���i��c�$2�����"��v�J��7�./�sQU0j}��h�i�%�̀��x|	v�ݘ�Y����v{�A:¢�"-��U�G���+��}v_����]��Dv�����^4���g,��k��`/��E#�7���c�)b61����f�k
�\�G��ѧ-@M�ͼDW�[k����áV�^�CDbIbα�?CPS�u�Hdyɐ.X��ڍ|�ʑ�����,a�Vzܞe`֒��1�zL|x%����Z�&�q�k�sQŧI��t�H�er�?��b�����a=-A��s��]V~�횢(��!�7��ߩD��)��EPc��"0+�v�Վ�O��"����	�+`���I�L���֮%gj���e��4�?�ZEv�%���m9,�s���GDE������.�*�|���UP	�88�����~ȿ5:�9uy�՞�І	-tj֭m^m����PiR�����*��U�P]T��t���av�g�bǖV�����4b����0��f��~�di�W=�IdwS��,C�ZsL�O��	ѲΖF�P9} �=���w-ćD8�z �2¨��j����6S�]?�u�� >���,�V3�.���?n�����'��:M��b��:K�SMǕڈ�M�>e��ƭhP���������\�$�# Ԍvi��F�U;כ�ڎ�&��:$B�,rd�L�:�!pk<�}紆�r��.���2n*ml&����@�\�����K��ss�?����MY�}� ����[��+�k&��X�¶�(M[�n �UC-��ݙU�/R�7`.�B�w[j���_�����3� ���w�<J`�=|�9K�d�`�f��؂IS���('8}�� ��+s�p	�O,�*�?�o�����{l�/S�HZ�C'�����=W�c�#�f�a�b���5,���⠏��]%���϶7��6CڈK�>�ٌh1+��/��c#�#���Ճ�� �m�4(a�hw�����1hL��$F\��7��փO?���=�Mi��Qu����*j���!sm���q?B�},��
�L�w]�3����2�5�,���FO�ѻ���S�[4�R+�'�������u�ʹoN����2W]�����|Z�%�V� �}��w6 �@p�ff$�$<�Tqm�e�q��X̲��,�o]%��J�n5ռ���u~�Q\�n�^�0�Zi�G�e:3EM牿2�Qһז��+F�f촐�����r�~��J�2y�p�$���F#��ंg��#sl�&�^L$�tR�eæ7w�E�9��T���嬗��y?��/1}��$�E�ʏ��[N�J��޼Ԗ��Q�z�^o�ٶ�0a�ͤ|B[��J_��M��C��=���2�\4#��f��6N�����Nd���Dż�AA������1��.��bVɊA�'��6!�?��3C��B2�^k�x��W��5W�3�T�XѮHf(��8�M��_!&��(B�	�ɠ��jβ��}�����bkn��<��
ê;*'r�����f�̑�*���T)�E�pd�f��K��FsG�F���������Z�P f���eo��"(ҡ�2�7}H_{?�����=��bt?N���T�^8���żm\�t�,�N��
����ԟ=77��>����MQ�SC�\<���k�s���[��fe���m��ke�2�z��U�[" 'ܠ��� nm��F�#�L��3Xw�6vQ�[cmUF�=!��uUY�wO���l-�Q��� �&��B1���q�3�o�R�<�VP��t
2�=u�rB�j�f���[e�x��xϖ+V���O`!8N�!�+k��t��N������9I񮯇�C/M �1E����|	��5�cN��R��^�h~n���&�|��r�n#�%�P�ԶX����B�+�(���ZOY�j��މ�(��Hj�R��S�Jއ>�4��W���a����H�Ϣ�"��n�6���/bD��D=����!��%�̣#�k�GSDWl��)S����:u㇎m7NTCT�u�X�#�������y�<Z���U�ɔg�*˥&N��6_ƅ5ֿ��'�_n�p�D"<VUQ�՝�!~�Fu&N!�G, �η��P��û7e���`�!�� �ݰ�@�a�d9C�´%� L5K�JG����7�r���f��������_SY�Y��1Ɓ\xy��9yg�\�^,����%��^����䔼P�ś��Bx�;&Ju��P�`�G�h�!��͗������,�m�R��u���J
h7�S�<���iJt�[EZ<�'�\����u��������В��N�
4SY�U��<:�Ҭ� ��70^�9�%���b1�6CwP5ξd�Jք:5t�ys���(��l<CY`0"�e�%8MN�D�?{o!CP�m)'�WO�I���Fg"ؾ�S�,Zm�c���]�:�(�����>̲1n�M%�*[wg״NU1K1T`� x�"�:U���\;��I�7է�Rd��lտNn��݈�N�j�H$
|Ʃ����X����W����y��R��BM��ס���x��#�*�����ꥵ�pʞ�`�T�������;�/�\�-� �o�̆��Q��T�����S#�A�uEL\��)������oaj�(&�+��w�
��$�6L�f��<��m03�<�\�����ͣk��Ԅ;�]N���&b�>-M��� �K?Ǽ��G!2R6jew�|�ߛ�SmH�9�����q�������ܗAeW<@jQ�}�`��'y��ɽ�b�P�},�#���[؍��ߛ�Z��/en� ��WDw&y����=c=��}��+x��~���z<�f0н���G�)��M�}��F���q�B��ŏF�jʵ�_�~�1���2v8}�B/"ah�7�ox�(�a7/�~�h"H�*�L�Ⱉ��*Qq�A{��b]Jp*i{Z���H=�Ɉs��@G�@����[_��VVLM���<ԫkX�Ɋ��7Q�3���Rw��Ui�T�/}�||ф��wva�:�/�d��2����Ij�m�+�(���J�$�gH�r�]w��p�b��å��{v�W�G�(��E��.?ٺ�]��=�K�(�Y7��69�����X4N���ɚOtB�� ��Խ��.�x8�O�]�_����P(�����<�W�E촙���L|��~��%��x�X����K�|
2�v2~�2�nB��'�B�� ����H[��������Fj����`>��宅��u���Z(��M�[��{"�B���#����[)8�/' f�Ώ�9�b���b����B�!R��aK�q�³ilَ9���"&���n��"�҅k��:� ���׶!Z-��e�$����4�V�����'�3��W�S�f��\T���`���W�;����T�@���.��A�����T�MV%5�ӆې �� 0Q�V;�K7���"�~h"x^�5(���h�AR��6�D��phj�4$��U�c����tcg�r���z�X5�r��4Z�>D�.�bg�|p�^'=����!�͟��̫qL�����q'5D~ܲ���{�Du��Yf՗,-U˜�.�B͌��c���j��<��H�"�ZTX[rʦ���a�/���o���W���1$�rz�����:P�_��v���m 5��+(�ە�K��|]Y�F�WR�&�G`�5K(�x��̈��n�GE]���E�g˰x�A�o��K�fŵe�9�R�گ
CB��\�O�\o��R��T�ܮ���OA�]�|>]�O�̄/���Em�6s#xd-�7�p^L��2�&r-���xʐ�v`X��.�c�|��j�e��I]Q��ɇlԓ�(���*uh+9��>�aQ��s�蕌ޯԍZ����wBFO
ō�_H�PNf�4�UZ������7����Ms�+��+K��x1`v�|�|@Cv�Sn��|С�I���;z��8�jI'g�ylJ�W�1���y4 ��sč�QT�'����6ر���w-�6�틗.פR��o�&nc65�����5ށt��N8�;"����ނV��@Y��;��N�ɡ�L��m5�HPJEt���o4X�D����oO;	r@j�ʴ��}� �M� �0�r#�������_x��S0�C,@����-N'7A��?<5m��ћq"� �t5�eg�,蚇8"������w��9�8a�,�5���������r�,��\Q�ܗ���!Ű���L���8
���� �<)������rp`�3���#2Ea`�����X �q�os[>�o���#Pb��p�;ŉ�t���M"�\vr�rF�z�O�t���K�8̨�o̘���� I"2�/�9�CɁ��Tf��}���)��uia��:��w���D�O�%$͜�*}�@a�?i��9�I�������^��|BT���PY�k8�Փ��#�XKhyS��3F}�{G�A�a�y�}s}r3~o�N~�S�0�3�e�r��`�*�������� U����5j�s�ZCG�_����ɐ���"G���U�QL��V�l�x%◨ı �38G'W1yu�G[��M�$G�ω�@c�A�ǫ�lJ��cv��:t`�tW--1��%�=�1��t�g��y�z��$�69�=�76��eǰ Ha0�Ư��#z0<-��?����#�)���흱q�G.����'&7�ɍo�']O�Yg�!��cG6�d�]�=
����+�m7A8�a�1+�2gn@����F���dm���t��S
!��4g��!D����<Ҕ��Q�d�TG���f��i�j����#7!�&6!+¤��������J�wGP��3]+&4X]�Ұ����u.)<��Bp���$�ޣ���9S�W����)���n�'��p��E�� �� ���L�%]���ǹ�WH�@����p���b�|�b���E������{�M�-����u8]�h�v��AO�z�5Ь���J�ѧ��v��t+�
�1dA<�ؔ��4�"��!����+qc���(�.��5��y�*�mךB��-��3����$�e���H���~��Xi;s��e�K�׻��6Socc6�;$���Q�ԟQ����[փ�D����YQc��A���C��Ɍy�Aƈ
��H�V��R�O�x�=Gϛ�$�S��#��?��_��&d_�0��*{��r+b.��m�[T�i� B������f�Z�A��"!�yT��������zmC��M�9�.K��Iƶ�@���.��y���D0�݌G�y
HƘ��]c��p}S!�2ӄ� YV�����6�����`r�O��g~�}C���_�,�lTz�����䨖�k����԰�).��֊!�����c����7n.)���r]����� �2ۏ��'�u���(�����b�	E��L\c?�/��ՇXC���V�4� �YF�[��~CH�V�B����g�0�A��d�f�� ��I�U�|�N0�*�>s�/u�O��(b�'QG��
�=�8%|�	�����j�w��ᒿc\6F4:�˭0�1�oo�`(� �s���F<�[�ߪzJRƼI���b�t�o����OOT"���ig �q'8ˮ
)��vC#\��S.4Լ`���������UP�͞���j����i�y��9>wʧ����\-�G~8p/a�i��Ŗ�RV����d��%��1��B�z<��U��u2�Lޙj�}@�7�/؇^��� r]5�L�p��,(<3��1+�2@�^i�	���,v_�3�r�����#@��h���������YEB ��`Vo ��c��TmX�8���I�z\!����hFo�@ui3�x����e�N;�1�{�,�ɉR5ɞ�ّL/kvš�1������� ęu��8z���n�i2T%e��1��
�_b��;.Ji]�Z& �_�Á���s�(U��xP����<�s_�F��Z">��:����Xc��.��Zx|��}A4b��1����G���Б�����;�h�*�x�"���V�KU}FQM�"�vb� im^Ji�F��e���S������E�YQ�Y-<{~�h������sd�QUց(�ES�D�a���}���~�wV�N�-yJH��z�B�%��Y!�W����z�nؠ �ڝ��a�����驋~@,�y��]@S0u��V]�c�@�=�8<���|���$�Ï��-Kg�`Э��	�O�R�-��eh`/���7�f���8�&���R_H��t[�s�5.wZ����fv>��.Jr���kE���ϰi'��,�����
�(���b%�%5x���W��Gn�1��tY�B���VUt�R��o�n��`?���[} ��"�
cB3^$�o�� ��G�O��T���E�?Wȶ���b}���yIӢ[5��)(.I���/�����R�[wi�kB�P��t�w����jm#n�0�?�B�-���	/�H6,�N�كz��O��TGA�X{�i��r�M"���ؘ�i�晗���=w�5���(�l'B����%=��Tt��fD]IO�@>���J�z���Y<�ѹ8��Ý!dC��C�N~��N*���g�A���S{�t���S,o1I�X�J�+Z3�Xy���v9PD��.mۀ]y��ɣ����_8KqV�	֝���c�$I8��$�lFM��7�hY�HBTFd��U�X�ƫ>� ��E����v�r#��`ة��n	q��.l6�": [$�Þ�m;;i��e�������tCX*X��Sv��'.���|��e���i�~�Ba�ղ#�i��9W��T�o�	3��zm�7 ��޺�H�j8��Z���M�'{����_l�'O)�a,�B�<DU;5����AD�6���7�J[�Y�"���O���\ҝv��H���Y�}���ؓ��!#�"���\��d�ك���������˺X<���mA�Vh����9a���';ʓ֯ݦ�Y$Z���5�h`��(��L8D\P�e�kF�Y��ٺi���q���i�p�>���ˢ
�u����ײ����ə>pG>�<�Ͱ7�"e^.W���2�c�7���y&'+;@�~S5�)!��{�}����j�G�A�p^|M�Od���C^E��@��p�8!���w�$iA�;�m:�ܯy`Yh��[�W��,(���{���_�����A�㏅��*��f�N�ӈ�K�2>q����nx���
��K)3�l��/��T���b�g|�y˘ ����L��D.���A����gD��K�����,�F&�\3
�~��[X]���uR?E(��	-�K�G�����eŋ*�CW|�Hlfc���!�z��E�'{-櫶��W6UB�
K������(��(=Y���%�@��u!}P��,m�&�'��c_�Hx��Q �߯C-��5; �qz��,+�i/u��<�ϰ�USݍ.��i�6��\?��v�������I�l�������O�I�t�VOhͧ6^���ҟ7���M?�,�[$����'����R	��}<&��;�\
-G4i�:D��5�����A�x��?�����9O 3@�w�{�ծX�|�;���Y��]�nMJMe�T
���٩ �q��3�aM����/B��'�*�n},ZI���E���V7'I�h	�O��r:��Ȓ!R�!?�  |-��	����/)6H�mvnD��"���͔e�B2|;��H)�����2S��$�1i�^6�H���x6��nfy�r)"#�ٵќ2��O�����g��IT�;�U�<���`���F���561�����ˮ�wwY��Y]j��p,
$����)h��*҅��)j<���M�O�i9��q?t� ^� ~�p�w�?��e\�t��	�Nu�X���<0���3���lZr���,K��vA���r�=������np�U"�D�'Y|$�85��o�e�����%՝Ѹ�����^��2���"�(X�M~�q�?O����o9)%�6������'���<��x�\#�3�\� �]�I^0��f�n�j@�&sͨ����j�Yb��xK{������XR�!��O���-k|��N�k;�<�#g{9:�"�pq�΃4Ғ,S�;����nJɉ��_i������x�e����b�0.z3e�F��$;ߏW8���������v�m`輙����e���Nb8�ݘ\\]F�1gW�X����}1^�c�`�%Z��rt�U ��:���
��Q���o)vP$J [�O~�;��	���
p�4�U�˛�ꍍNU)d�N�C��A�7�x�dIW	�J������]/]0��Z[7ͦ]����������1Xk��q����eq�� @�=vW4�ܴ�Y�|�V�V��"7��ԕE��������&�}�GU��B��G�� �@�g���ִ�������g]�3�瞤xf�*��wD!$���9^�Kf��k�;�y����0��b���V�M�-1�dn�u�K�E�-n8w�O	�}w�o�i�-�i�\��ɺ|0;�U��Ksin�V,؜�V�=�ycn��z�ɚ�CM�,(iG�����j��d��NؓX���
��ѯ�^,��� �܏Tm�b
���;�p��0;rM���2�(�?��RT�i�^���Q�[]{�X+RC�!B���/m\�E*�ߊ�z2���%p5{f|�Q���.`My�I�9f�0j�ۡs�����aێ#ml<���������^D��hY�l�(F�V��o���ƻ��oIh�b�j�g4gc��'�K�ƽ��A�b)�͔^�$i�7e��`�g��W�_����̱�5y[�0�=���k��Y?3�S���D�Ӯ�4d�8K��F�g��V���Шl�C���FL�x\����0Ҭl�"WeR�UqQ�4q�kN����%�[��
��&���{��<�=�-@`�����6��h%�G���^xwn<�q�=W�^��C��J��Ѫp] O��T�����>�v Wr�������r9�L[�1@v���K����k5�h6�0�&@�|O,�I!qX��W�K��%nu���z�y��)3U9b��.t=U����}1E�,Z�@���`�DI�I;�PD� �4�*.Sf}�@P\���)9 É���V[j���)a!>dUG�='u�SQ q��<"��& ��9����R����}�r�(ӈ��ªV�o6�e+AhiF���gE�<@�������<�k�0�-("��3��{%�%Y�%�vV��h"Ibz��̆�F-��'eD�l�HN�Q���y#K�e�;�E6�`���HPP��R�Y2���W����v�=j�j����F���;�ڜ��-pQp;*䆩�2�&��I���'�Z���$n��#hk|Wv&9� ��r,�jf��yD 7�����=���
��3(���ZW ^
O�K�z�r
��J]���w}��h����ހ�T���m���S�ՠЮ����±�˸pj|e�:���`�_��f��ݘz��T�:�9ks�,�Z�p�G�F������!����<�=�Y"�3�jm�gI�f�3�_,Yr��AY�fm��T�2���9����y�Z����k#��.�ٌ��E`��#����_�/P>�a���
�M�8��� �2���=C�"999)g^*+��>ND��}q��f%.�	�W�s�k$�U�	�9�P�{��7Zr�QrC�[��0N�=�6�F��.�Ipkْ�!s2k��p_-�q\�;�����@T�P�y��(��c�E�<�ߋEO��>�衢I�~�c����Y��$ɔJF*A�"�R�u=_-Q?$ٕ��X��J9������!�X��p�"� U����3�����(�B�~�]#��`1�G?�pŚ�2��2����� �ȶs�I�� �����!�-;������>�hb�.�@P��>�.?-%�e��7Ҏ4�-usi�*0��\�G���_��]��ŷ=Շ���#M����$�IF@D}���Z�T^Ř��yȮX�}��
l��B|�Myp���8�Z�0I/)=g� ��t�j�d�up��u����l{�ƣ���48 x��q//ß�T=��3Q����/	��7?|�k��g@��ǋ�Z���H�k��������q̈3�/�4p����x��^jX�#�f�'�EC�����ya��۾C͉�����:]ލ~;��Q�u�8��Y�݊�m�u1�G,�����OM�g�ۖY
hJ�_6�@/�����κ�0�D��U���9����dY^Vq:��VGq� J��a��5�Aa	�g@�33��DWc���ɖ�~�/�/����2�1�Kŗ�d�{FQ<;�(u�%d�ED���*�������p�/tu�? �L%�<��x�A�e|+A�C�h����5�g�Y�K.p���iK�[O�w���oڃ[x�����}_N~�����:��6�d��Z��ԙ�/��n]�bDX t�Z�yB�2��R�t)��H,�.�}�Y31���t�g(W���iޓ��,�6{+� ć�(fGq��64��D��}C�Ʃ�.j�b�lx�� �,�P��c*�0�v�=�����Sk��_���#!Ae���v�A�4>�Q�;�WR,�V�f�3eD=��Q>0��ExZ$��JZ�M�җVHWwv��'B��:��n7t�� S�tG0A���K8�����˼S�¹�D�Nx2�e�Tz� �F +���*/C_"ꗆ��F�\7<-�40ƇEZP�6c�ȵ����"����r��%l�R{3��-oS��jv�e���|SMh���#��Y�dB{�����Bla-�Y�8�K�u�+.A�)X��F�$(��Q�!d���a��x��ʨnE7\s�8�^�azŀK�H)K\jjUv�m�^FX�>�T!bѓj$ش��7��u%���zy������W�?b��z�o	�D-�������:>踊�h��cV���;k<���+^��s6����r�������z�g�X����5�"���a��ӈpg��h}�nE+���.>���q�Lg,��x�R'�T�:���W�K�b[�_���2���M��I�M���$l����0`���*�/՝�Ѵ�M�>{�غ>r>�d��51/v�[|�s�a;w��れ	܄5�LA>j�e���g��	���Xf����C5����9Oy{ǌ=?���3�Q(LP����/�?�j�6��
�uK��;�+�E�Oo�|���	�'�J�߂G�t!�������֍vö��bj��j��V;hvvD�|�*$s�]��5ref*�����F�G�2��
�L|��"���~� �N��z[~I�k�;)�;�~}�*FG�L��h	W�� Y��R��h��F���tG�H�lؑ�~!G��o�T8��L< k4��XOP�a�gЁ�M�3)6	9�Znd��BkOt/j��=<f2�O���f5�?j���}X!N/�����ː�,eY��(e-�~BWI>�@�R������=��Bǧ Ku&>Md�?�����H�+F�t!�$1C`Z��Q�t�:~.�;8D�NԞ�V��O��&?����eD��_��}2�QLY�,�[��љ>���7GM��J�Mɕ! �gKWm������s��ahvKN�h$At��@bD5��o���#O�8�c��!ؐzֵ�9e���o�ْ�Ŏ�p�ڋ1~�e��^�4�WR�p�U�@��L�X]}��\_�|"��zh4���wL��y�R������P0��0�[�(i���©lZ8��k�do����UxJd�m�۞�CP�y�^��cS�S
Q� �^ ��2Z�0MM(\�}�|GU|+5G�kO\8&���[�FB�*��J U�<5��؄�ׄp'$x ��Cz��S��)&��񦦔}yO)��BK5���"eʰ���\���L(����rh��G�[�'u��ݐ(0���Z���3!��z��n�!�Z?���h�m���P&Ggz��0W_������{>�����Y��%(Ry���60��*1��N�\Ҹ}�
k����a�7+�U��l�{��;��Y����׼9&y'W+�/�X�+eF��t�q��:�  ]���#c�d���!K���I=�^��Pt��B���u����V�傮<h��ȃ��o��/��Ur��|%�niF�4�7���j�M@��V����〥K-�5t7�B������+�=�\�Q���������0Bħ�7���.m%9x	3�6ؤvWU�^���j�wЀ�/����`yE��`ۺp������LmP@�R��������rj��BsrLq-��#��qד{I;VA���D���lL{{�����VIv�M�s92�����B�$?��LE�"�3��Y93Քw����e?�s'�l$����*G��T�3��X��O� �D�<=$�'L���p9�+�ʼ��]=�.A�b`jH5y�8h������.�(B3|u� �� ����G�5�I�&c�ō�)���h7a��>xï��.޷�s�� 9�k��-�ۚKP؅��N,���h1�����1�<����F���H#ZU�Ϛ3;�HIV}Fp2 [C}Rq[Z P��ͼ�i���}䆅��2KS�	���\#;��}��D���
;S��u	�1�c�>s�@�F ��,����yv��!Xv�+:e}��g7XC�;A��Ih��B"M7��ĭ4�bA<��>}�bwO�)"�>
WH�x��7۝?;�fj��u�������=������_���k�6PU?�ݳ�h7��%�h �TGYnw�W�~b�C����m�G��2`�:�m��^/=�	T��o�̆�i%�<E��05�FQI��Ò� k��\���v��8-9�RD�!2d=6X;%�B����W���v��`�9��!�3/�8�ůk��5����˻�\�p�7���X�&r�o�� %�V���M����qa�68f�cgV�b�f�=}1��ם
���^M\{B��z>l���v	��j
���0m�X��?��x�8��on17-^z��4ڇ�$�!���[>��T���R��ZK֟�TA�$��Q^�&��=1�!˴l1���b�k^p�@p�U\�P3MG���J|�]RD|JA1�?l�J�9(��lq�u���t_�I:�Vw��x̆�s�8�Ae[�_�~
�C9X�˛c��6�Ԅ�uL�s-�0	y�?/2N��0��ȗ��v�901�Bh�w#h.t��Ċ$K��)zt�M_st�*�]�a���y��7B Ӆ`���Z&k���
�Dt�΁7=��+{��"b$,>2�:�(���hD���Y��v�:��m����i�L���.��=[�D� Hd]E7l
�.�G����H@���/�D�=J��M�,��QB�w��)���Nz9f< ��z�Sy��N� ���è��R���}"�1���������+��ߓ�XEE�ZE�#:Ӱ;W���˞��O.�a�Fh�m�I\\:[{��#������W��*f�,���*��~��9Y\)��"�S�7�$y�$~������a+��k�_[B)	���Kn���Ji ���~Hу�6M%g������Zܰ]���'
��5��!���"㔧�����o���S�Y'���a���E�ļ
MqNa��ӥM�]zh���$ �C��t�B=���<��rE�b���Ȯ(`q��8w�>�ǎcv��B�`:�dOi�^����#ս�UyQ+Zpu��c=57 ��d!j� Jpv�j;U��A�݃Ո36PD��3�й��Ð4�*��uP���zL��|_:IH<k2�t'p��)�[!)�vM�*�N���RqNfQ�|��*��k
����ԓ!��J�����,�O ���P�0tK����:�̛e�V��n�Ӡ�,�K+��4�ΡQ�c�'7sE��'d�z�������\����EE�%�V�U���9U-�i�9Q�=������[����;�&���_�ȑs��6��G�e�M�x{����;Qf)~�?	� LBc|�z��@�V��%�|�DZ"�{��b���W(?�Nu�d��Ui�������\6wZ��-�5�� H���LW���s���s*h���A|��Ǌ����������*N˞�z�����$�0��%5.��t����W7Qqf�2SD����cb6ۏ�����84~qd*���{��[�1^��QX�ob�w�mچC�<F�w�v�Of������5�i�b��6i��������)���%g:~�>�߱&E�ח��+��PJ�uՆ�;�6��ò�_D��CЇ�I����%U?e �2�6"�������Q��K�/Y6��L.���C��i�[�s�-�"�qY�z��"E{���-j���R��_��N$-��8ﴨ��_��L�O�3��~`t!P�L�8^����_��|tT���0���K)�&�Y�tzXV�>\�Sȓ���,r؏�?�= �Ƥ�F��"26}[�g]w�U�)��c�#���r���?^	�JT�2�=��DV�x9�.S�	Xd~VE���.(�*��&FE\͈�aNۈ�
ݩ�|��Jֹc���`��� �Bn���%��D*匄�9�Ť����#!��L�8��M��7�Tg�@h%nb"�g�Dk����E_����/[@���΀xIw�j���,X�^:+GqFػ��\�~���x����ᒟ�|WnɤA�l�L Z�M.&S$+��]�;L�3��c���|�@h���j��ۘ�}��n%�W���p�E�Y�D�����~Z���716N��c�:Q��z��g��������}\�TD��cok��O'���6������d����[���f.�Kʠ�ļiގ�&5��/�����K&�,<��Q���ŵ��r��s۴�,���u�i����+-����m�����h���P��j^�l>�<�Tz�h3���r%Q�	���H��C�NA�Z��2��Ȗ�}|�:И��m��\�O�by텲Ń�t8p.��;V�*I�^�{�.�I��kM�����������O�*"eDOF���Х(�yI�Iq�7ܘ-'lGI��QOD�����u��u-~.���E4�K)�D-��RJ���8�x�y�*}�`�T�1S�
��}|��G��Q�}F����"�H�?��H0S�,������`j��BuH��a����	�@�J'!90
צ�1�I3`��wҐ ���n��-� �q;���e��k6���(G�t�d 䡞���^����	S�Q1��d�8!P.'(D����_�R�[�Lg��� Ź������C�8�o&��2���n�i��)�
�z�ܼӦ^H�P{
���w�Z�����_	[�;��s��L�d�%�:���`� L�G�A%���X�W�-H^���ը���u�>��cTP���y�������W�`��`*JE�M�"��f�\@���d�Wi��8��������8���`�%������Ln��j��o����Ru�\5�}����R��	}��}�^D�a�����L� �h�z,�b��F�4ur�Z-�ҹ榑c��WͬmT�����5�wHA�C�m��Q�s&���{�;�-�a�ⴿ	}��?3�D�g��G��e;���Ŗ�#���,�I�EN��=���6�`�����d�Ң��N�m��^��~v/M�:���y�9�2�C
,��m1���L4 ����!s�����o�b�jY�c��s���7c"+ݴ��.b�q,8�������Î��+Y �3��?��#�lf0�C�n�Q\F�-��n��h9�dfÓ�ݽ����p��i'�Q�c�	3� �N�`�T*u����&Jt�ES��	�.��³|p�5M��<���ӵ.���y��uw�1c<ə�p-��#���'5�f�T�S�y���l�����#��/��.��Dv-&�y��D��U��B�8�t"�`��z�.�8���H����݀�?X&	$�}���#��F�j=��GY�$@�<J(Ĝ�º.j� o��E�P�[ƚ�ڀ.R!k�e$����v��?�3�Q&W�������[Y�@��m8Xr��Plׯ�������Z�vȐ�q5׉��`z�2�b���&�F��E=�����.S�&K 0�mE����5�f�W\zos"����)k3�QTcV�+��n6-�,���G�2���'�����E_hPO��"������<����N�IN���Us޿>���$�.o yF>ݙ�ր��C�ث�ߵQ����f<�٩U		в��ӫ$�6�|�L��"�r�C�/yt�X�\H����E�9�Mh��Ae���xVY�;���/�\_��m�Y�� �e�]\G�k�r
�L+֊�A�����*�;�7CT]�o-tǋ��{5g�e��)"�Q,F᷀8hU"��LxPUoU"2!�r��(�֚M|��B�e�X�	�CttyRI�t��n]+蝛�K'�o��+
:���Û�<�����s�z76�PQ��I�Z�8�[���C�#���3<q�x����o�pdd���͉(q���}� y�5KH��3Կ"�s�5$tU.�K\7��:�6���!��b7����ε�0�rj+:�MI��Tջɳe APw{��hX�i���K?�d�7k����~48#X����2��Z�	ۂ���7�<�����_��m�ƪ�4+w�*��!r�B��W���Ĕׯ��3:�2�\t���|5�k��D��İZ�K�#W�id�(�3Ч��5a�e6P�\pb>lQ?��n��8�X��[Hw��VHv�fX1����T�����f�������w�)����Z��0k*��SM���zu�5l����a��J3�C7��C$
u^	�r�1T�>���$uݷ�� �$&���˳�ᷴ$C�Px���ߣ���:�r*0�CPw��U	rK�ai%,��l<E���j� W=#�_��B���}��4�&�R�(G����6�F�R!9��C1�K�uoәSض�:;���){~�I�8��t�A�s4�7:.'Uyf�hdk�\�/-p�8�|���ιa�qH6X�c��g�l�ڴ|���,�J�u/i�cK��������,d�lM~�Eo�x��Mv��qo|�������aE���W/�h��Z��`�Q�L���󂈟��Ԡo"��DI�ԆVPQ:����t�?ֿ�T����"0���1e���W�ib�Z�A��R[���`�_�"��H�	f��a�e�"��$>)Ǐ��� �6��9�aJ�헰��RЩ�
�.���BĢo�=8�9��&����G6H��8;�;��+YWF�?@{�ʀ;�6��)�5ت�y��%d"��.5[�9�7��V̌IGI�\A�5�c��;�7ЌX�ğ��IL��_����!PZO7�XF+?5�-�
�v���A�>�.�Y��� �
��3�?G��r���ol��,{N!/�����u� {mSt�դGk����L�����&�G��6M���&�(�����W�JyJu�p�s�;��",3@�,�P�����3U�u)A3X�-`�J�q�xGF�k���j�;�A�cQ��Λ��1�v��
��&ݴ�R�r�kB3�Q��3wC�u������޿����s��l|@s{`a*��H��VgJ �8�p�0.*Fڰ[�%#�q��1�QV�YgC@�м�m^��tL�f"�U�:?K����떇Mfz�,p�^ !G"��)��q:`��kѲ,b�\���|3^&�U�q��8߶|ֈ.*!9m&`��);�h)�d���m�.H�O��!`^Hǐ��KɏxV��浭Z`(�'b��ZO.W:ל�A���#�Ӣ�0��y�
�j�ߙ�}��h�r�-��5�/q���wɍƤ �2/Ax<�ն�Q�wv��(�y=��ǟ�4��$e��`a=����нL��$���Q�9ү���`?����4L��k��+t	�m�W� z5���vy���&��2��Z���=$�0��x�3�	���#���l $gCG⿆8>���<2��s>I��z�V7M3o�� ���>�4>Yo����4������*NOTUQ��݉c����������C�*�U=�����a�x� �@�n$o�p� ���9Pl~���[d'n0�FɋK9���&[�=ꠂ�ck��u��=�����-g�x&;�Y��h�H�S��IiY��/��32�œ�}��'��6�@��>� �'���<A��34���{l,ح��������J�0�;���c��r��۞'Һ�[0���[3"��>!�X�������=O�D�R�L��`�q)ӮX��� �������o	�e�͸���?�j�w�:�6�$K�i��E�4	h� 5{��_�ݑ�A*��
-��@��2����nP�{i��Z�%bG��U̿M��|Ka��:���X��a����p��ۜ1UN_2�4yޚEX1E~�WJ�^{
��3NP�>��A8&�����x/�hA�I�H��_�M����{��]=��sLn1�V��*�^vm��g�
����=�A�?�q�(rl���j���?�pg�yz���4�{
���)=�mc��'ڈ]����韹s�E�b�ֺ�W����N�<�~彨
j�&�OCYj�3���W$�s�ߜV��W^W'd!5�gR�e*9��Ә٥>_<e�=����U[l�^��%��z�@*��8���\��Щ�3'p�ı�B�7�i<�xΐ.T�C���X�Ig��,���ؿ���K>��S�)���G�"BNyf`�Mfϲ#��w��1�4�a#Z��Vh�:��*���ʎ*s��p���b�G��f�Y	�[�~�e~ѿ�D+�H���׬p�C@�h*HF`k��QZ٤��h�KSx0��PfE�e	�ױ���H5���� Ò�M�N�8;�M������;&�>:�&,�@*��L�-Q3�#�Zt������18��FJ�J/��IU����H%%\YĮs���ti2K<����h���J7�+@��/s��IS��!=p�ڰ\}D�/�|�k$�_ ��C��Uk_�֮�	�]S��U�j���r1ٌJ��s�i�{1�O�9�}̲N�|<����RaY��
���v�/�L.��>�x��DD D;m��s\)�#�=(Ꚛ�1 `W�O�W���H/�#'��+dU���Z�k�A���@Ts�Z�ғf�8���ʷ��i3o�=�^w���8�#����+�$�{G������M(�f/J��׎��,4S��O�%1�E�F�ss}�d>7�ҽ�Z��D'�ٽD��<m��ʾ��.#�	_�'7m������H����L�Ш؎f�9/@ڷ#�d�-B<a.���5�AΧ+o����RlGTC�-(�:9�ǵ��
/Y����ϵBTg��i%p)�G���Ɇ��~6�����I&.� �_��U�Qꔵ�b��Vz�*����\�d@U{�Wo��2!9��Yg�fɘ��Z�7�V�2~��Bnh����@�V�KS�V:���xm�����#���Q����0�V��
�&�tE	��1pr����r�p<Fx�ޓ�ߔ�U�$��,�G��y�T�$�Q �XF��ٙd:���;L��P�S���~|�Q�j���:Ad`�A�7ɢ�G���C]-[�y}�щ�����Gr	z@
�-$؊<��͏�_����HaM睢�j�n���}�!\���{F6�se�Gwh�H��o���F;���@�>���SF��7���q������3�DZλ��M�>8'�,� Z���A>���;F�L0�sc�-zV�M{���P����~px\���oE��?�!V�સ� wVg*b*a*���2�]��M����nG�.���s������@��x���@I|�Ͱ����3|ت���j�����פT�\�߼�ߓ�lv�-��C2y�	fB�ds^v�<����O��F������x=�g ��W�U����a5�c:�s�L��i��$��bFa�d��O��W���4fp;6�c�`��&�+���Ӧ�3�xi���+�-�˃��j��{֨����#�%���N%u�ǰ%]������O�𪓯[�
�^��f��Syϲ�f�Tr_����X
�D?䒟������C�h���H�$`�	2� <�p�WM�g��$^9���k��m��C����9S�TY$yH
ųy%��T%Jv���XS�{C��N�C_�J]�#:�$�6@m�7х�B�d~�����+�h�I-�5�#���̜i�w��U���߬GdE���d�o��=ρÕz6Q�
ӟ�Q��`4��o'���6�}��R��9�Y0���ZŞ;H�6n��XI�@)|h�hz�B��Rۖ �Zoa֝�j�C�h�g����
�C
���^�T��Hj����.����.�*t��=p׿�25��'�4����~��ɘ�f�mY�=��\�~r�;�df���0;M�l���Ŵ���3��@������aa�C׽g�i�)9c� �m���ڈ��e�)9B� ��ү���;��7j���Qy��-:��X\���a���#������1\+�r*�hR\W�ݛ؎�L3b*H2τ��qF�� %�yn`N]�v�+?WKv̸Ѐ�ztB�aeD+;��W��I�4?u)�KDe��B$�mw�� ݨ#�J1��_�C��u�f,Є�QK��y(�y��wc�c�;��"��{}��P�S���Wʄ�v[���PF���t�>��ѦQB��KN�y����ߎeO��-/��2x+�2�� ~^?�)�v��)�^|f�A��l�ض����U��'���QU�'*xB�¸�x�><@��l%j�W.K��J\f�5X������YR@��N �$ϊ��Հ(ܑ�b�F��e�Lh��0Q++�q��ܠ_��g��!�&Y�OG֌Q�=|[��9ؽ*��e������s�ĵp���˃���O@Di-�B�����Y.~>��c���t���>C<~c�Z�c[%]+׎�����sA�Oo1�+�j�wA�S̽�_Fr��jB+eW"<�wW,iH�g��!�ĲӕO��� G��<�a=�h-5���;�ъ��c� )�׃�&,D�i�W�ű����Q�$6&�8d zJ�zR��C"w�CV��4L�g��o\ �<���_�x�Y�
a|3`@:�1*B��z.i¥��:P�8{��C0�v�	lx<"�6�����vbg%`۱�Ps�!�<e��QH�*L��9�=�-69rZ�N{�xQ1��j��U��tWi�E�`D�|a�/K�Fxv�l	�4�f��ao|k�U����b�&=h0L�wm2����7<}E±[�u��G��{�XɌ�Kd�WVr�� ���6���/غ��d+EW �Y�IU1�|>\�~�m�_�C iP�e󇳔�m�[�*4{ο����ĩ�>�% �q��v]��0jkm�f [����~��K���q,��Ι?���9t^�S�B���@���oaG�RI�$�1�0��qoI��Ԋ2`
5��Z�V6�Uw�;�M�mun���7#ؠ��1(ΐv���lH۽Yk���/R��!}gk���,���F�	GX��,s� �[=6��-�d3;� 5�|�녂��V��q`��Ug���V�F=�D�ڦ��c����KhP`�,"��њ�?��Rj��M� @�ٻ41����-����#�8����k�J0_���X�I���܄va//��greX�S��/�����FTz�7:-�(����oY�lө�-"��u��1fZ��.9�Nef>IIe�@@�	<���l�a�T�%�?Q��i�Ӷ��׬���-8h=�Q��(Ɏ�s���u=����NS&�#���=!��co��Ͳ��yn�dX��B&Y�?Ne�Cc��ui�V~˛rX���	m+���
��xq�oƮ]3Y�u
�ؙ0o��i�X4}X5Ӏk�����g8��9˩BR��/8]A�x*�kÈ ���A4
�jc:jK����M��ttPH?�=�ׇ��HXj��"F�������ӡcjX_��=��l��QOϾ�3�w�PG�M]@�R32����I9�
�p��)#����E}��Y|�0���9ҌF��"j~B��q<F{�����%|��8JO<Gz�j�I{^kb�?�U<|Q���딮֨D��46�r$A%�kzz�d�ؐI�ȊǪ�&���;�[x̓��5�%j�y��wRoq��`����w�U��Ƹ�̌op�7�ri�Ǟ�7��~A��@̣|������MCF/UV�Uե�p���Xh������0�BL\Q�!��@w>�Y}�e��}�o�ޭp/%�L���7L�������Oi�^��6��V�q��t�3"�p�h���g�L��! pf�s�c|�'���`��9�F���O��I��v���ȷY���!���:��^pNRa���^W�Ud8��Q��݅\�x�2gH �Ťwxi9n|���u0�1�|}�A�"m+O�$��E�Y��~̉�.�$����fu�R�>�wع&�;����W-�/�t�֚��6|s���������J��,2)f=���u�u_�9���_��g�)s�9��Bɟ�M>U�6�0�z.	�2X��'����iG�N������aR�C�P�H=1�u��i�w����-�H�9�,���r+)��R'��݀>�� !����K6q��Z�"�Jte �0�l/"��=�!<��=���u���g79u�RJ9�lz�Q�Uy�S�j�h��mW����f��V(�����f)�����/���@��r��ך�%YU�#�<���ݥ"=ڒ��ˀT�fq\�r޿"�ҩX��4���2u#&;RëCW+�� �Y�ɍ��>����wi�hz�����䆭5S<���"W;at2eȀ��V�g�l``l�� �Z�t$ɕ�ۙ㈶��KLr�;�o����^d��+�@*���gI���4&X��?�|�Mb��t�Pґ�(�̢���ު��tIK� �n�A8��IeS���0mn)m��ޯ��MZ�`�k�ͫ�k�<�?1�>��	+"�����n��Q�W�u.�6q�="KG.���`�W��[���Q� SQ�5����~B�:8b�e���j���Em@}ûwdL=�W3i�f� ���}	�����ȟ���2*�	j����d���pw�[���0�2<�Q���!��-���.h� �0��AY�%��oݎ~��u����5)�
��p���~�iJ4m�k�ږss[W�����&��{ʻ���v�K���B�G�9'�lc�vX�)�_��o�(Lr�h ��+�`��KX����$�(Jg�qؕ8�#:ϼD��A��8'q�ߪ�*^-/tȰ���g {�Ж��
`��If9�f������mwo�_~�	ɘ)7�V��f�,��ʋ�`X�̍��4��Zv@�����{��7���e�?���d�	9HF�ʣf��iY��(�
t�E�����G�L$.����u�n��;���Z[S��ue���>�P�ǌ�k�Է
h��S�qDy��M:�$����՜P��;rM�)z�
K���*X��?.�[�K�Q|b�}Y�cbiGo	2�$;t�j��m�� tX��2)���-H���jz=6��!(1�-,������x�4����d�����+�X��u_��Ӡ����{a@{=�ȶoxs\��|�Q�SM� �ij�,��qU��� �ٚ�H��.NF��3��M�4����~�T��
=�TE���	b�<�Uĝc�'�x��Y<��� ���u�r4\�z��V�4�rT7��.�1�h���Uh����|O[�Jp,n.h�QC��.�F��r��	@	P�AT�~`�XrL#g\�g�����v*�K�%;�T��8��#�v�����sK���P>��J$��q�M��Z�i׶$@݌�1l��ȷ���hjn�g\i�Mdڵ�5= !�p�ǆ"ږ�p��ߪ�,��b���b�7�<t'42yK��l�����ҡ$u#���@��3)�:"�>�x1���wg���\�<�65wN5�&��ۜl%K݉e5�4�1��ť�Z��#��Y�� h��x���o,/˦�?���uq'�\�&��V��;GkjL��ShRu{����3����5¹H.�-9��̎��%�(�辇X}RƱ�}�J%�ev�t�V�y��d�U���''�&�P���u� @3[SLj=Bԝ�|�[�M�h�r���S��e�K�&uNC�`	g8pv�!���(��/&µNF"[\�8�1��s����{-BU#-Q�U�0n��Xl�'R�Qk�瀐�p8�z��ԃ>��>{C~�-�wǄ�	�77C�H7�[��:;�a�h,M��<Ĳj�0�F΋Ewd֋�p�l�FlGF��:�3�љ ����к�E��mʁ�h���E�h��\KsA%��&�>�j���O31�{2)�+�3XdW��p�BO��R�GߡǾ!P\���~K�Dv��Rp�o�
#ΊG���s֟mVy�R�<$�86|˻4c�7�M��ġOIKzR�y���'���s5�̰�,fUn����j��%��s�Gd�>�'������
�!�t��y�j���/�	�$���(f�m�.�r�Vǃ�Bq,�X����S�D�g�̡o��5��(dk-YܖO/��+����q,f��NZ�0,"YwP�wt���p=�&�Ƅ���1H%�4� ��d� F�@ _=Wn"l3O���t�����E�t��&������{��D����V�B�e���K�6��qq!/v3yB��ɕ���S^`�]$��t�ԋY��9p�]l�J�LC�g
u�:����鏶E�_AHd7>�����f	�e�1~c����P��oE��J���1	m@˦hT�$;�o��vt,��5΢�GDx1�B���Y��m?�c�a���49<����d��,�Z�F_Vc��%�qr#� ����u�9�Ο�NS!�������Hژ����ۈ���Zv�>6�z.S���۝ln�T>w~��s_�}!�Wt������5�M��,�F��cnC���*�x$�E�8W�%���2��-��#2r��6��nH��[W]d���VD�����|qdF�����^��S�P6�p�W�Dm(9���Yp	����x������9��p��B�����/���<�i;v%1
�l��z�`���b<��u�O�B�[���f`�q��έ�<����� WJ�+A�c�@�_�w)��%��o����32����9~��0FD����uAV: YX����m��N 8�
E8��	y�2Mn<KLL	�>�$9@�Zv��|�`�����N�F-�m���~si[ůh���i�Z���K�OyM�(�]\D��ʠR�Qk��D��9H��Ka�� l�ȹ���.��5��*#]��JmDT�l~���3�JI�2�L$u,'"X5�B�u�Yxy-l����<(+ѻ�Hh��69��V��>�W���=�X3���az���ޔ�u��me��@@��.���u$���<�&]�N�B܏�
L�m��gD�h��@��U��M���b�o_�H�p�=��@���7�x��o��#imf��yō��}>�pL$�w���u1:lQ���yf�5n��A@rk6���}0��*�PG����ZK���<u����W�y���ǥe��ͪ͠7�u�����4\~�C\���Y��(��2ryU�'�|7n3-[��Y�iPYI]K$�VC码~5�joњ���@A��u9A�V�z�<ŷr�q_,w:�T֎��Y'��Qqpɰ�7i�C�����8�#ӝ�w���Yq���?m�8���^�C�b~q
=�tN�g�B �ɝ�B�l����]�CD\�f}�5lwG��[%��Q9���j��ęauo��E�Ns�Y+�}���P� ������A�wnS����Y8�^�9O�ܑ�c#���M�4	I-@MѴ
tg=�����u����4��o[`ֈ}@�,C�������l`�l�\��/'�"ۈ�zIEr��]��m߆�ܺ���1`婘tr��[q5���ͩ���*�SʨG��a�V�-
	иB�a7l+�}A�]/���"'�C�3�׏4��O�,[���Tl�ID2,v�]�>��L��1z���9�j��V�v:D`q-YYO:Zw��4�q�6����ؑ]D͠�'9rOT^X�P�l�x/f�0����1��V+Y�,��Zjdu�t���/U���̱{v�}�e?"q��GXd�Ŕ��E�,Ϳ�1c�d|oi;Vu\���]V�����#��j+�H��1A�{��PO a�:_��3���jn�h@�k�Js��X��P��8���V�1�:���>�%��9��ۓ����$�.�9���s�6�k>(�U5Į>��"
�s�G�=#7��S�lp"@8R�x]�3��I�Np���21/j�}�,MW;&����~�1hIM��N�o���A]*�Xc�DT�:�*��(�˱!p�o~#y����n,�R�~�q�:Q�rK*��e�}y�i9Ҫ���D����Hu8�ʁY`d1��i-�,a��V1o$�SC�W���)0_�i���M�ibN[�{KDN%���c_s�+��U�@���w	���qe�Z���y��M�x�����F#&pMGٍ/����]]a����#82�yt=�ו�8�'��;�x�~) �F���S"!o���xAon�R��0��`�2����E��&[��e�k�m%Ќ��$���-�6;8wxUKJق�]�7�S�.�7�+��T� ��Y>.�$��au�S^̍�M�G=	DDUn����b�Ui��RUo���0<�g�T�&ێ�_,\���RMQñ��庆��s�ZD�R�����`/����TWM�fvLJ1>:�q>b���9q�J�!��,]ɽ�͏��ˡ@�����d�B�����w��h�������ЪK���>�5Ε;`���k_�̃"�ߓ��]ev��1�پ�jF̫<���M:e�Q�)	��0RܼEX]��:�ǭ�I��/��,�J�r�	�c���3c��7&z�H�e{yC5	�RLn{bt)7ZK=_�Ja7LH�������n{�h����D^��$fo*����Ɣ��X���ոJ����!t��la-i-�����x�N���.�L�ǎ/[������j��	�+A_����R�.|��A|�6�#>���6_�s���
\"�Ɵ�g�b��JD��b���&�Z��ӈvr(�](nQ��Q2� 3�)s
|�Y���������
��Flzc����,��"ౌ<[89���N�e+8���~�f�&��5�Ъ�Z��o�����5��:��;&��=�SϹs�7j����%��x��fd� S�2�����JU��o_�<3�¡C��d5rR�r��<��5��n�E����ӾI���:�\��v9\��E��D)g���:�
$wX��"�7̨���5���xw����xQ�Q|��W�m��^�8c��J�0b
�7(�0�u��J��Z<؁�����"R�_��j�E�k5>K1W�?��Dan�Jp�C�u��D3[C� 9J�Y�Ƽ�1|N~w����}^= �5������|�E��������g
������g6=���l�|�{%j��rG�F
�5r/�von�:q9���{%�4(�19�v�e�v�B���d�vm�LZ���߼>D��m��I������H$͓�c�q.��!�F��7G,O���]V���c�Vۥ�|�I\}.�����bfU
��8�iBnpv��8�`p��8�%!�BW��'_-?����U�+����񩦠��L���@=��T��?��=���"�6�s��Byڻc�Ě&�ū��k����JD�)�7uT|���	auM�~P�.? R���8B�\��� K�}�l���xJ��?ntO�^'5��W+�+�f���2[���["K�zE���F=�av���d`�l��_l.���o�w������f�ig��י�2�M� Z`%����R��Sõ:ăwe./?�Ƒ|B�6Nk�d��rH�(v0:C"���2��_u�p1�Y���,�bYnu�lf�SA�B⃅����)��&�����N���Q��F�1��{�m �9yV���������#�(/��# 2/����q���8.��ԓ b�9w���򐀼�I"���a�*x4ݬ��?;�"-C|�1�;k���0ȫ���}�0�| P3�2m�*j�K�kPQ|���;��stg�0�'Nd��w � ʯ�	&�㸽z��a�t���t����	9x�\��ETQ*n�+�r`�j�a}:�ѣ V\Z����j����c�
��#o�v���L<OC�����@�Q�j�8�6�6��&,���Oؤ�-Y��U�~��W��X��a��jY��'"X�%!T��z�]���%L��v������w�*H03�G{���'-��h7�}�W����ײ|�IL@��&�2=�����T�	Z����Jq���#ص�=Yq�j8��1�}�;4U��1�/Z��ޓ������l�x�S�U:�Ї�P�@�}���.*�a��v�	��P3���zL��_�
'�=s�1�d	Tu]�s�l�}��3����%�ZH][�矵<ɟ����%���6�f}��*�3)P�>W�@�^-�����O?�l�O�>���X���z_x�.6ɇ�w�Lrܧ\��;[>L�A�P����dn��׶ҺaQ�=D�"ڹF,�!&A�@9��� Z��F\c�6�is�Ok�g�fW��rF�i���p�K���?N�"씢)#-}=����=�򢶳b舵/��}��jT._����eD�t�P��ʦ7#q�P�Y��\��������\�q���/L�)�(�F�]���?��j]1���$��C+�C�E7���)��hh�s
���`�>��̍��>Ms{�Jx�݀��Lɚ����N ���kƽ��X	�/�e>6�D٪XH7��v�=f�ee]'��%��6�$o+���;5N���.��T=V�C+=�k���T T���玅8}oS"�r�����=G_����=F��_:B1��%
k��}\N"$�\�b��F�{Y.-��O�IS��ļd���H�+m/�1c<_�L,,�Q��͋	�+ť�wb������+�s�l�>�oHL'���=S��D
��})��s�
���\F��q��{7�ɜ�p�p�5���fk0?!����tt>5�zc������?m�{���҆K$�4P���ف�j,RE�ĉ��jiֆ���2K�����u��c���ӌ��*�4��"����������zGw�eYR�sz���U���>s�i/Lm����3�.lL[����V� ��X(�&D�=z.[T���ItnFA�Źι�V�^�+�����]����S�0dc���:l�(_R6�r1L���(�u�'����u�����I͸+P(0|��6�%B#4�Ap-��[�h+�I��
���'�7��WV��kܻ�i�8��6c�O�+���*��M��l{qf߼�-�٣����^���#�DJ˚���t"����2�6��R�k��+4�����iV�1�G��N�Yެq9�TK�)�L��t�}�j4ץ�vX�����h`�1���|��比�F<Lt���m0p|�M@��=o!g� ��%��{������vwŠ�,J�{��_�)�m���8F6��b�8r��E1�pO'��zM����4*��8�^Kk�WO?��B��t��^r�|:�d�"q�Օ�fl\r�F�hG���y�d�d	Vj�] \�I�|e?�sNՃC��%I�]����U�r���+9���v.M��͏<�Dj'�U�W����ݨr$9]��E��h����_��@����U�=d!Iu�R�����t�"qO{�ai�Q5��]8�0�!�ɠ� 5h����M^(�q���z�$��ɸ�Uh���Y�uR�m9-LIe']��Epܲ�N-z�QP�L����v����d�""B�;��m6�V�����K��ͺ>`jխ6W��sGU���e~X�I� =�A�� ��/�0�o�*����O�$&��-����Y�XX�I�'�7b"ۓ���FC�!��Tt1/�=�ƪ.ԾԠ��b�|݋�b_fQ��T���_�U>f��W��P-���y�����z$����Y|!Jz}�����L��!8��K�c���/=�Nlo�R��v����
�O%O�t���d���qqV�#)�Ծ&���7�Z5M6���	�]"j]ͳq~����F�6o�pq�E��+
�����λh���!�V��"�����`;�8�y��`r��/���9ǁ���b;+p~O�b�k�aZ�6L
�����H��7�^�����f��9�M�<���l[)��Q0'��$�oDMl����	�+m"��o� ��n��-h˜�
��K݅�3������u���G�YG�	��U}^��4S�[&�=�NVo�}w�7c�K�k�6���8B+9����T�Ɇ�j��=1$�_�ɾ��AѵW�Z}5����e�7�#�{��@��b�/k��i@�Wj�Pm�Cw���T֨��P�,���mD�~���s����'\9�Y�%E��{��4C3m5�^�4��έXQ*�90�s���ՋKo���έ�p�ݘa�G���ʿ@5:� �qS��M��e� ���a��/_$䗽D�Hq|w`�v�H���,ZTH�k��c>�o9��VCf��y��,�^Ѓ�ST�)�.�E�����0�HY��D���X���� ��I�l��Mo�=hT���#���9K��,p҉F��z���y�I[��eZ�1`Jz��5ܚ6督��aAa@�C�&S��@��$���A���U{I̉!�I���nngcA� �3Ů%�_���n4������h ����EA�M&,q�m
�?OT��n�[���}?�ɪC�SހH���j�f̇�'��+}�U��W���h!㙂�^��=  ����ޗ3;���p/��B��}Aq��F\���p��왽Q7Z�fK�!|�����(�?QQv;@�E�	`�ߨg����:��u)
�,��F�ǳ�Wè�R_�����wUU(k�M���9~�5��J7��ei���i���	 ����$	���� f˟�+;��|i�
1���둃� �$7��Yܓщ�a�򕉃o%Kf�C�KE's.�D Z�� �
���o���2�}'��^���tX8�^��څ?�*LZX�7�>�+ԇ�c���c�����j�/�wP��=0�}`ի1$�LZ@2hB�O�@C�!\�mB���?�:��|U�����cq�1(��!:�j��5�ԡ������5��hᨅ-@��Ѷd-�N6 ����l�kB�D@ZX�m�����%j%���>Ȓ�X^ΕB�9�$�%��X�N�fdU@
�
�Q�e6��謷W%PƎo�N�k���]����7���XA�N*N�(�o��lWf}GveZ�^���I��g���5�S>����J��"�_URf�Y��'���l���nی�A�=�Ě�5!����*�w�"�`!��X4{���+��:�Reo�z�5�c��Ȟ�p�h:T]C��`�XS�[s���BK�ͥ��@N�t:C������0+Dvp��)�]$��`���ex	�������eF��Kì���0��.b.G��Ƶ׌�����k���-�w=�[QX8�أb�""'�39ģ��l�wov%@}N{�<W~<�m�t�k�2_��6b�	�����B�3O�ZnhT�vݠ|���Uo}H�\[@?�*�8�e��yd�j�T6�Q(�����\�wS�|SI.�!�oƊl�����4&�����)�;���l��k3,{�p�=��n�B����;�|�4~x1�,Z�A^�߾�,SO�m�(��C5���Eue�'��(q=���e��$_p6�S,��*�S�E�.������Y�ZѦ�.XG��'�42�6g?�I��%^��VaP�&�/��
u�(�$�Kc��@����"Y�i9�4@�!�38�K��
� I��H�U�D?�};��IּsodᖜF�6�+@]BD��δ���X��\W�YUJC$r���Z�A�sEF������ m��٭��/^`k���WD=kP1�i��߰���0u��>½�ra�m�F�"|p�"֪J� o�۹fe��Y�&g��/(���50�9�Jscs����	��E�+��/���78�MiA�.CAQr�ڃ2����D���cK�L��4���&�"����8nQ����ZL>�;;5������C`�[��tZ� ���3L�]f��dd_o����j�;�h2]�e>G��6b�qAnZk{~���b#o���"���ȒPx1��zk+:}����2O`R�1�u�Fk��Pu�~�F)L�����	l�i�.����Z�)�	!���@��1P�d=� ����ع���=xDUfe#�/&C$�J����q{�rSMDpK���W��M�C�sr�L@B��\�fc2b�6GB
,KF�K8�M�s�|��d'��U9>X�^��0ѕ</L��	�1��n�>H�u�$����?��_���Bǌ=��b��tR�M��g�UX?��,.r��
�&PJ����O��@s�J��߭�(�ڂe�%�۞��T%��_e�@��sR�@�e?�+�)���.�*/�=��1K��z�X�^��99ߥց]@�x���Y��ˈ�I�f��"x'"��rW�n�,"6�!�J�$+��ćm�RB���� ?B��j�9.}�	 �jŘ���i�|#�E��TJ$�����@z\���tE.^�\� {e�t��iM�AFfR��-���=J�C�KˊAe=+����4�������NVm����T� >��N�͆��9(�6$����HlW��^Wyj��rQ�������6�ku�Ϥ�Ϥ��CA�� v���e|:D3F0e��4�F��3Q{�_06Mk�[T�N���<"���w�[���!�o�ڃcp���S�5�2���U�#TG�e����y>E,��8���@U  ^%!��O׆�~l�7u���lX�����:k�Mp�c�i��$,Ha���-���_I�O�Wk#����vH|�������#8S����(ZՍ��L��P��$����QF�|�3�]F�f�)���ፀ+M�-Z���+ذ��@?6������8�5���*U`��q�x�u�)����%�8<%w�:<��l��5�S�'��b�0���S����ᭋ���t��{��Mz'��yu�G��i���I���O���n�jJѦ��2_��hr�W��P���'4�c��5��e+?�[:'��W�r��A�W��
���zڧQW� �y韽0�$
ފ:�\���:�4l�T�ɿJN�C䎷&
�jX��5��1��C��4�Ȝ��07��=��h�p���B�hd@�`��@����,V�-Z��5�%=�K�J�pA�<��0�|��جg�M�Q"~����`-�:Wև�&�];��wEٸ�@x�G���v�C;��r�n4�5�2���ݾxL2A�Ȍ$r��}��1��5���@2,B#�]p�����҄��#��At�YU���'fӝi����樈G0�U%��\���x	,�G�-�Y�#4����Zee2*.y��v��~�|�K����s�%CM��'y�*�2$Γ��K�:��	���ʬn�[T�z����h�C&!�� �!��hP�s�� 1"�VFR.��"y�oo~h���f�q,�����^[��B���t��C9:�q��o��� %$���2����6��ɭ�a-/ ?��~ٍ�i������К�u��5|�42gf�'��V��F�,\bv�Nk�J7	+�u�#[Pj�O0�,�=��NoZ}>X�x�B}e��2��T���4�������+-�A褦k/3����_�a���� �%�έ��S�e�n1/ށaɶe���a��1�{*��B�
�t=ك�b�wF6
�ei5
��y*�w �;�,η���',#Qb�V�x"d�#�u�Z⤃K6�q	=��*h3�ǣ���R��,OxM�a�8RUhI%���2��.�R2$��0��.�AS�bt���ɛ�E�U��,J�:�'�I�G�"��ɾǶ,{_#Ѵ0�=�C���1`�D1w1׼��s�}�8�
��(A���y��m}Ԍt�^tk�f�},�A��?��ɰ3:@�_V&�}��:�e���#�%S�%��L2rL��H��ȇ��z#���4o�/#+
�y�; �n"Is+c�g.E4�!��%,�9��4��}'��[��Uڞ͗پZ��^ѻ&ے������4�-�i"��ڄ<���aXbv9�k1����@�j3�t@���Lΰ�\��o���Hr�L��܃BpP4[Nu�BG���>�I�|����"~��y{h�Ӓ+�q٦��ր����>XI�`k�l/!Q;Ո`��"/!T���C�ݳ�脾����@�Q~�y
��֢�b-��4�<�-�QI�P2OQOЩ�?ޣ�ܳ}�����^�jE?�:[���. �B!9�����ֱ�>6��5�����)�}�+�	B/�ѩ�F3b9:�Ӕ70E@�+�<���8�?>�O F\Pp�.�< Շ�ٸ�f�<̂�U.$r�m_A bg���R�=�3@��oE7��a��R)jiY�"0urs���ͦ 5z
[_������._���H��B��/���G,u��Qhź�|Y|t�����ee��zb�.p��P\�>e���O��ē�*`]h����Z��5�����^��4�1�uٙd���z�:�c�J<�C+'�u嘽��;O=%2@�\�j;�	,�b����A͎b)���no�{l�3����*k>f)������ܣ��+ݏ��v�����e���ғ���$b���cjBA�,bq 7��#�	_q���4*�#s�9B�!�y�0\c��gEE�� ��S,�������^�ݑo\�.�#��K��rV�p�+��(S�Q"�/� O��̀E6C#Ďu�����e�^�r���c�Ƃ.��݆���!$�����),�J�B�4NM�^Gg�A��N��]�d��|�ҭZsѴ1���q�Z���?�B��݁���7�F{�0q�a�qFv �:��X���g�7���������>�S!�0�G?C��@s~���鏠dj1�n��5�m��"+a�޳��	�<��=��J��3G$V�X�u*���鿢:���[���e��Hi��r�k+K�]��f&E=]�Qw.�T������]�'p�hy� �c�z(1��Ę��͉@0@�9��0�L�_�&�v:�0]õNR�h���
�C�8���P�o�%A��V�Z�d�6�k-�lR��qla��bC�Z����S��`A�dU $��7d����Y�����Aԣ!��@���"J`]���! ���FDe$q
x��kxY,��rՅ<[vMO���z�R�0*N� �}TB�+נ��Cl�[w�s���S��6���~.�]�[��u�>o�gN�[h E<��,���X�l����ԕZs��TH�LKV��s�{Z�{j����a&!,>p��ZS#?:�9|��3���x���:�������/��z����J��:'&e..����۾��[���;뵈�5?M���ʧa���ŝ�p�aa�/`>�$�� HC� :�X=�R���yˎэ��݄v0C0{A��PI��G�MxD>E�0X7:�A���=pwZb����{������;��>����*����]v{��@�+,s䎎_�J�<�2x֘G��S�/�O[x.'ĕ-�ʳy�2)��8DBI Oŏ�M��D�������fTU`(o�p�A���񜶪�|E�&_��������4=T;�S(�v�fn���D'��Җ���Eܐ{�ܾ�Բq84:Eg��>D+Ϋ�c� ��]�B����-%9yq��3��xĄ����G���2����{��ww���HW<HDZ��&zk��5| @{���DX�* l�sv1!�K�K�~\�o�w��ė�b��ȷR�
ۻ���%����^�}�����ÉE�8�랊Ǫ&C��l{�"��nYXBI�����md��S#ZOO���>��"��L���0���?���w�)�<ݤd~ԭ���zĶT�nR�t����T>
K�����ߩ6�V��̶��~\��>���B�Ŝ�1��>.�f�2E,��/;��f'�F�Mt�a8�8��9�3
��49���K�B��т�
�T?I�;��۾'g�x�����|qʠDR5�Z�k\?:��}�Ȉ?���X��~&��>ܘ��H�}�3x���r'��%m$R�]`��f6��i:A2v�Ԙ!<h��$ \�l�D&G��x�ilX�@�GZ��A_nNS'i��2��V��Q��6�9+ QK�aŎ"ލ)k���չ�6����(�s��`v�i��P��1��얩��,w�4xD��'����f�<UkƵmmwk�����ϫg�.��!ad����.�Ăg���_W���W�`���=xc����d9p0�z*��O�xk�V�,j
%���O���k���b�(�� {��8}ӄ)�x5HgJ��e0z�2wa&C,���:�
��&��(�d��,�6�MD˾p��؉��;��^ʬ�W������Ӂ֓�9��y`�5�9��ЎC�[M���k=�bʽ�_���j�('R�5�Z��wB�b.��%�9� XJ��죕Vɋ;͓z����Z*9����
��DI�T�ü�����nmo��'Ԯ���`'4������L���� *J9r'<��5��+r��%�C����R��o�7�H[ɞ�,���q;�
�y{��y�i�ԋǘ��֚�V�}^�lJE���Z�q~lÔQv:䕙����c��2��vSrF���S9F�l�7�9�:�_�D�B�����3y OxY�r~OR�GkC��0�ؙg7'�����^���7y|�WX�@sx�L����i�����G���\�1T&i`�iz��9ڸ�s~$s�X�pDeq�̯�E�g����Y��.C�7}f�(���ØRf.�����b\���آ3-��'$��Y`3}��@ĕ7�]na)f=��"V'��hPte�&n�#��Ԯ�W08�L�J�Sn5�=�0��58 �23|4������<�r��V �	��i�.F�����!����������56�7��u;�����%,�z�P�z��^���^�s����XJ��eM2#(M�^zA�D��@N�UI61��e�%���]���D��5���x�\��z,z*�fg0 1Y�U�(�[8�N��1-(�K{z��
K#-�)A��^�Pko.�'Z�\��-��8-���}���oL��K�|���kJ_�,8����	�&�3�g!Zg�ʨ���Xֵ�;7�p��k�Q�'��/FC�ԃ�8Ǭ0����.���+3����ti�O��:���	̾����3���5���EV����nąx0"�X�Aben�T���,%�%<�$W�J��i�]��c��ȴ��M'{�u��an���үZ�<�F� ��#�*&8%�(����Cw?/I\5ijA�.7.aZ027��\kN&��l�X����[��L���֩����3K飵�q��k�%� ��z��\�'P|oV2B�#��w��?\�#O�^�iz�����/��
cɎ겊�ݜ:��7�=3l�Њ++M�����rlg�����-�}�>N�,ƶ�@��?z@�"���B`�=Eξg-�:׾@z�7���#��� �alg�B�va`���_�g0�I��m)��gM��n��W�� �o��k;bdz��h��E:�g�|z�h�蟢+B� 
wc5B\��1�R�4
�G��&/2,�bg��1����~���_�w���2��e5h��~�����AʱUօca����yc&
�*$��<Ƙ����j����o=4`�!Ef&k���m� }Z�u���6�+��t��QQ��/7,ה#}#�5Yg6��gN����T�t�^Q�YF�94[~����`�������U��Ay$��n�@��\����L��D��tG�A��)%����2Z+�V���f�Y�=WZd�={w�{�	���j��2���z�>ML��uN�Hh�\�:��4���[��!+�&sj �8�v�r�S��?��_MI�薂�^�����T������,��s��>�0���\��.��6U�pD��АV������.'	@�o����=��Z��xf�Hv4���n���A�l���Z7��O��X��Q�Q��aBT��xh��zJ�w�����~����'Y�\Z�Pc���v�Qϒ��	�S�|�vTFF$Qܝۚ	�F�?o�����س�K�~���5���RVpX�9��$L������{Zh�ߥg�>6�(�>�R����ua��hJ�s�K]��aVQ׿Ӽ>�adɈ�Ȣ��4�~F!�r~x�����"J���<�l�Y��(�Ю���\���x���y$��c��jsӲg,�T���i������ V1�B��ُ�?c\ը� ���?�vsT1�#S/Pj)ad���|d���S����6ӛ��Ԧ���2�$q��/P�_�I���)
0$�ut;��$4ivpc���Wt�3��c�?�O�������8ש��y�M�[���̈��d��c1�K��a��n����䆊Cŷ}�Oa��$G��Ƌ�Bv��"TՁ9貐���`c�7�B[@�r$����C�㝊'}(BWJ�m�"�5�1��#�:�w��߃�j��p�l�@�gJA�� q��>Qt�b��o�B�`�X���ϖ���F��d���;1�-+�Zt���uF��V�g>"� S��/,�F3���Ԡ$!I'�
����x�|���t\ȹ� H?��$U�ڹΨ��A�?HP����ӻC���<CM���rCi\'%;�.��������,���W�`@V�ˋ�����[�?@;�����$��#��k[p�u�� �!�ߎ��_���m;.��R��&���l�?Ah��O5�1�0n rO��� ����rȚw�ĕqn:^W���?Xma�ƑO���AN�����V,�Q!���� ���'���+�����}W����/�ZPe��w~;Ŭ�E�Nz�O�n^��KN��T+CC��8�K�j$�-ӿ���!̋�6�q�O5A\u�n'ߘ��z��o��@lp�VJc�p���0��i�r�A��F���w\-�A�ыi�4�&����,1���3�����.���8��^r�A;*���*A}�X��6Y�J^O��Ҩ;��~m{y]^¶EF�k�s��:�px�Z��
)�S�'L7с�bW���%�Y�3��[��6���S��$[e݆>5�����j��_	s�Q���Vl�L
֓��S��^=k!)^g��\�V!7\�qxt�fVrŵѹ�A��Ӵ^�����7�����]dbr�g��������Injj���ni�['o
�G�^eЏ}TH���a#
��D"�A����p4N<�bTz�I,�<�{ �܌[��m��T�ah1,���-�?˴���aİ��X&q>/��D~�J�]mL����^-
sdǮ���!"�LM,ARm�ǩPQR<�g�h>gO3 V]�-`�	U�h�&
zh"4!��>)�XR�؈�Z<�!'�)3�����^��j�d�c�N �w�Wt��������2�8i����T�����bPU:��y��D�R���.2��� ���� �"��J �.o1R���Om����c1���������dm4�����%"���=T̜1��Q�o]F�r8�M�fFGL�j�>���?_F�u(��:$O2���`�Yd��� 3�ړ]R������fs�gE���/�����\0�7bμ[K�.���݃AN���R�خ�v�Td"��	2���څ��ކ���J���P#�_�$Ȓ}��U�q�Umt<&�$|f���,����Y�����PJM:�d�o4��Q*��xE���Q�O��%�ݐm����f�)��Vvtu��h ���y�R��z��{7w�sC7\��]1J9� VtX��q.�a���T*ȿ�׉@>Ĥ��9��j ��W:q��-�0�q�%xc��NNK�R����t�eOzb���K#L2	pd�\�{Ɔ�^��PS��eo�@@B�A�L��éȣ�?��A.rY��<�ג�1�Y����`�F4.��v���v��8���؀�Ϟ\�Ş��s�mA�ڏ��	z2KW�d56�3<��G�_;՚#�7�Ml�5B���{��2!���?�d8uN�����~�Ti�$g��|�#+��XKXrq�s�$v�'��E��>��m�5y�>d.ˊ:�W�%d'20K�S����� 	л�����!4�Uf���
��{M� 1����|Q�.�5�8jm���!9j9ݺe�/�V �r� �mR6�nf�]_iJ��uY_}i�Re)�]a����ƅ}�Z�C���Z���­����-[��2��t(V��ה �Y ��/S�<qbTg��y5=�3��:��7_�����Ie*��F���ݾ��k�c��(��]��Ѫ9(mr|�u>w���4���g��w�j_n%��Jh{�D�wS!�Wꐩtx�<P��;0������	a�9d�XѪ����H���嘢ֿ�R�B�T��@�

���jm����9UE��Sq(�+w'}��[Ih�<�t����ǉ���(�F�=�a��e�NOb2�#u�H.���d˻��ێ:Z�U�rͼ���;|�"�ˍɬ�ȩ28�zt���P�,&|��#��Xd�� &�6KC@�5��"=}q��/�\��]�u}��0W�@R�e%���	/6,%Ȋ]���|ޝ��Fz(�c���Qz�ب`��d�"8�]4)��`�Җ��fCs�@?���k3��C���#Yc�f"P	@FA�9�1D��)Ī��,�R'���~��RW��ɔJ}��F�D��HK�	�l�"I���o���OL�� !�)C�7��M�P�M�t�d�f
�?͚���V�Wz�e�+�l�N�'�T5�:,ҽźC��&�u�Z����R�=�P]�i�-�-�ȹ%2��/~�!r��Gn	�N�����+6�6[�{�ح�s�O&�gV9�\��1�+��'�wS-I�=����-RD��G�C�tz� 랗�S�T�O�HF������&1�̑�+����!˜�D����WAY#(��s�����s��[}V �9���@��]6�UZմѩ�x�iEo��r���WN�7�ʯ���`X�;���~�.�#�8�ap��֞�|��C�!��?�ҏ�Ε�y�p?ς�I'�?�*���}6�:��%c@r|w���(�r$l#zT�m��ͱwZz��a�ǹ�P��I�����'&������`BT_X���ui�0��}����fri�u�;gg�򝽹4�?~�Y��Ϣ��bzf�&LH�)���s�쓊���-y|�Ԥ�/�+��yE�V��&cZI�O��1��Ip�=3/.�☊�Į�7��a�M���-�.p?đq�$��_��k�2��=;�1`�b��`_C�4�����|
��a��|�d�?����-B���_9,�o9�ۻ�C��O��(���Q��k+��s��6
h�-=9�`��'��F��#Jr�`�	�$m��c�#E�5M��H�����?�]egP@�<�;D�PI���)�2P�)��6�E�jD���ɓ[\�*"n>�jڂ�b�Ƭ;���)��|*�ͫі� ��ٍ��F��*Sgۙ����^���>�5�u������OT�9.�d����j(gI
o��'������2��/�\1��z��j�JcVW.nn]���հ�9O綊�f!�XG@���J��x��`zo� �����P�����Z� �e��m+�ٱ�`��H��ZY�W���K̄�� ��!m
�Ӓ��l>�H[��(%����pe�B���URa�<ց� �ݾ���+�*]���#@铲�#_��_��Q�#1r�<7+U����3�1m�xM�HkP�*%� �FP���BKw�+�^�Ky:�P�g�ӎ�/��N�� �J�]c��0��q˪V��������*#�T��ǥG�5 S��%Tu
t���r�Q��itOf�qY��kVD��G�P��*,�}��Ix���G��]A���i��ߋ|C�ċ4C�>zľ�<)���s��]o�д�r`~Y6����{{�88��������00O9f1�k4�)<.�Y�j�Q��o�a�1-W��#_K�`!����$+&S�r���Ɗ�z/�88���:����߆�����������Z�o���d�vt�丧\����4Dn�z�X���|p��)�1	�,FQ�\r�������2p�R�]v��i���1��O�2�����<������O�x&	��o2�{��B}���$蘅�/�~�`ԏ�Sײ��\�;/�k!� 5j%���:]�������a�]G��t�+��vTck�LNW0����e|PfsbL��_l�_?ٞ(p��������Aw&�g:i��wD]%u���Sw�i���V��R����I��}���hP��{�_�?;�Ϋ����k��xͬG�����k��l�7��1EJa�xg�	��?��a��0��D��-쥉��l�� )����A̅ ��^"���؜�K9�V�#�L��|i��|���$1�,R�p�x�2	��ΆN�k������a5;�lM>_HL�n�%*j��۲�LD�~��|��g�p����	RF�q�����|�t�݋p������&E@a�ѣ2j��j��|z�/�a3��Ǣ�a��JHP��=�t1j�)�`S�
�ۖa�l�E�v�%�� ~����HAy*:d�,�������^)g�g��Wj����Q�����&A����׃�7]���V^>D`r���<���OJ�W��l����/O�ˎ�~�q�.X\���iO���\`)4�d��o�^=���Y� w���R�/6�s�� ��q<�x����hCa_���TF!�.�E�\v.��bH�.�{��U[h�55h��iɭ��l���V��v�؃P[݃�ޛ:nS`|W������V��4�];*Z�>��f8��ruL�;�~MSg�+�:U�=>�i�����+��+2-�V��Y<�@���8,�����Ai|E�[g�K[#�/Μ���(ݻ;Ӕde�u�>E�Kx�n�|�n���֯�����\F-��*P�4�]�-�T[ѵ^��.u����dC��_kÚ�C�4u�&p̧��������WsXh���j5v%�H��n!�!���gI�J+x
�� �Nb��H{R)-n��L��Jء�xm�P���ˏ��Y6��<TmOA3��&���՞�#���M��aėE�g,�C�q������\��ѷ`,���[b�� �d�xO�"a�+]^9��������o��������I�nv�|i��HƵ5�nP<�t-���^>��6 �!%����|�5�g��S1�1[�������_�B�,�ifT��g9R�z1�f���*+�7��jIj	Wb�����C��� ����1p����%뜕׹LUav��'H�tb<���c��X�6������P���v5���*�&�X[!��t�qF׹��	g�4�Y/�R���������_2�0�/��Ai���[��N���0��ݶ��.o���%=e��Δ��j��4����A�6$�4��
�=K�Z\��M�I�d�[U�v�ԳI	�鮱|�k�3�$)]�To���0�BB��k��crr�����|-�TN�̋:�xJY��&�\�suKa���Z�)�oz���gpˑ���
�-��_cl� oB In�oM�Ԑ�^.V��e�f����N7���iI��\��y��Z��@�����\��ejp�q�A�doC�6��M��i��*
����K�V�c��"���b���h�Y�(�2V2�i���ӶE�nÒV��^���q�OB x�ו�Ie@
��/���.�g��l^e\���n^M��љj�:Ab�&�M5�i
ʭ�G�AJ^����Ů�x��=�cӊk{�N�F�5�x��|��iav �������gb��!�WlP�p�A��،:-���LNէX�ދy��o�ŏX(9?�R@�`%� ��.8�%��Gԍ*k�eS M���#Gaz��b��Z�5J"�z:T��j�m)��Q�$BK�׋0eb@tʮ��g��D�2K�u����X��l�Τ��ϓ�21n�ĥ H���w��H�#Y���7�,��ݳ]#Gް5}��U�P{��5�Vd�qs.5j�6i;�RMnRxX<�Y�g�A��9>��-�WX�a�mTfN@��Y�:�l��뵥E �#�G�W�Ӵ�L�ݙE�×��G�]7��O�ҹڏf"|�bH��C9A�d��/m)���8Y �����d:A�T�s�a:M$-e�/�!j+�Q"��V��#��`���io"�^��Ep��SW��ir�c�CsK�$���,��L��E;V����a�92d��Ǵ,�{�`ǔ	���?����� o��e��(�"M�m=�a�Y:�nS�3�Z�������,QEO�]R Qr���E�"l� #��2yp3�??�n�;c���@zH�S߈ux7���t��LH�|�fY2q-��&-�_z�!��y���˩�R׀m��=С���޺��;HZ�9�M}�݃ݐ.�O��j�	q[cUl<ؼ��"�m���k@�:�L��3�@�b�}:]��	m�.hd|q�YH�r�wr�DT�y�6XH���Z~�9es��k����߄u=����̂�$d�҅�˓���P�dC���^Ej�r�UPR#��ݩ/ 7�{��5�o���^<�.3�iEcp��Z�GoCf#|>� dl��R��:�y��<��փ�������vb�P��q�4�"˶�����ꅓ�Y�#���S[q�B��B�1���p�B|���Pi��=-�g)B1ON#t����k�C��Z��C*p��
�u�S�1�p�2��ȷ��LV>
^��Z1G0|r���D)L-�唽y��BhݗP$�4�.�-{(e����~���yi ������	ͅۅ�����
G8�)����/�v���?u����eAƏ�$�.I�\��:��d��8��s�I�\)] �1��'�.����Wr�sx$l�w��i!߳�.�{�q l��
��J<�[}[��F�"K%�|�����5S���#�"7�Bcz̨20�0W3�R� �=r��;,p�]z�zq�#^��71L͈�6ԏm�4 n��")��ʾ��D�O��x5O��I]Ow  �liQo�t^��0�'�G��!��:Z��s��(f��w�g���l
v'�8W��� k�&�Z�eY��ϱ���]���*m��sI}H�g���=β%�CF�%�:��yl�Q�_�Cs�1Ԋ��
���~@4٠y�>�E����'��[�$vV[Ph�Ź3R���s�M߷�j�I�]��$��w-�LY'I؁��urmP���1��\��w۱=b<	<X>z62����3�CQ���hH;�É���G��Fw��K$�>L�-pF��b��#����GY%7xG8!db#�&D΢Q9���f̈�`X>�.ڗt@e��>L�N�V*�'��	�q�����IK�F��j�\dclԐ�X�&nS��0���e2e��h�>�Y���p�N=l.q�	%���@��I���F��Cp|���!Q���9�.�͏%���G��߱U-��fc��4�Ǔ��Oji㻑��l�K�.�l�ra��X��K�}�#t^5 J�bh^�{�
���6�f���(���8s��8��M������wcIB���%>�_�z4����+���X������n����% ��p_��i�ψs�3Zݫ_B~{�
�[2t�}8t���s��qd����=8)T���\d�|	��e8>�O�8��؜�{�s�Pk� �8/��#��:��
χ���\�^Lpsg�P���hm%-r�	]o����x%���x���4�����"?f���Q���i���>e5>[���,� �9���R���i_�9p�缞�44z$�7*���p��A�r�Y���m�F\W\&�PY�^	8�}�B�up�+K�f�<H�0W�͆,#$��F�Np��ϸ\Y�X��U�B���w��q��rbJs-���{�;��� ��(~\���"�s�B�Z��v��7��y��~,��w`A�[�<����T�WƬ�Idi8��l�H�y���Xm*jB���bm�[t{���	 ��W�#�
،׹@��ͧ,O�dcz�9��c�	k�0����mi�M-���R��%��"B���j��x���r���`_�s:���ۆ_�?b�y'���3����A��5quS��u�LaꞳ��N⼛\t4����3�UJ�?�![����� ���v�1O�h]�'�EG��ม�"��~+P�\�� D�4������䕬5�l}�7"�ei�K���, u��FA��#)�u�~��8�snhG��+���E�~z������+Y�H^���hT��`4e��k�A�B���q'�|���1 Bg�b#�a���>:	.eF�?)���~��ؘ��\���{�|[�]dϰ�ޓ�@�2�dϚ�i8A��Z���So�#8]��K�m�����v�e7�Zy�9��}!ն�UB/J�RA�N&K:��T���O�~���h�=�+ x�zc�ߡ҆���{λB���ڼ�P�w��dﴺ���b�YfmIلߓ8�D�]������[-T=�[�����TTGw��{���>ҍ���}k[GӐ��E\���ns�[���	`��I&*T�f�:1%���j%�%@�ަ�9�`T�iB���\����\�f�I���K�oo��|6Ϣ˯�>ƴ��+F�)1�2/�Y���X��;w�*ˇX�u{^(���7�]�n�!NF��	�AK�@�;�f'�&���a�E�IJ,�f�0�;��ͣ	��,s���s`|[0��c��,R�4�՛�9WD�LY�pK����r�H{}�-P�J��\���%!��ս�ܨp�D	��!���!$c�O���V?����I�s�}=Z�fV�˃�}h������ā
?>�aA��~k-_��0�jJ�o�B�7��w��e����fM�5J��k��[�t�/n���M�AD(��@�!\Id]�'�1Q(���#a�[wi�R�UNve�o�Ň�)ub]R���C��w
�a,�x�Fy�O��?S)��<����5=.)NM�ƋnMWv�x��}��+a$����6��RO���'ݬ.����~����ۄ͌�y��=��&��ϛ$8l�K�+;�9g���ӇR	y&�z���?��X�f�??q�7yH��ఆk9.��gL/:�#�1zM��`1������&D�Y=]�:]���n�v���v����h�P����{���䙴/���x�dr�(��k�N��lt�x���#�BR�z�@;��A�Pů������B�n$u_��ZC$7P3��@�cU��2��>̣U�}ZW��J{�l���O�գ�)���_��5���Bno����Ǒ�U�5��{�7�P�q}=0ӂvJG�����Z\T��؇�f�mѮ�ܙ�������~�UC��oʥ�%��Y�W�h	4�; jD�\˟m�o�hf��G�A��yt��ɷ�#��R%��6�t$7�y���."i�_�E�O���V��\"�]���� �%��T�}#&xBo9��66�/l6�/H�?�� H��0v��7z�[��@ג3 =i�6#�o	ߦ�n�3ٸe��\��2�P)�Z6P�mJǗ]>Z�dHf`�*.�
a+l-���I!���z��p
�&�����C�B�E��8�'Sr��=dS,5,vW�\��"�wG���n�y�&����0�A�G8���d8k�zN3HSq��ٻu�
�P~K,G�TX�u��D���J 
ū��ʑ��{cJ�C�?r�$A�΀!q��n|*�MQTH��/d3�h�/�������a��!N�[��Յ� ,YWB��D���r�򊜐3�)�ߙ')a@�	(������T^&��b&<��u�.Y���fv�Vh�q��l
�;��I�T�f����z�{�[�o���O���%�'o��;ܗs�p�-���vU��n?�9���x>����)�f��m����5"b�^2Yk�zy��"�Ie�[qR�E煈� �dT�)��J������3c�-c�
�����C9>��k�B�=�-~f�,o6b��y��]K�a�_'2u� �6͚V���F3}��ZG����Z�	a�,c��C[���}��5�ц�4�X
Y����Ti�*��C�5�=ܶ����J�� 1��u�_�c�_�PT� \�\�8�;/��XVr�j��q��8�-�3�T7ˆ*fi���,�U�g�N��>;gbI9�����6N<=R�H�BL(3$e�Rs!�퍵��!���^��GP��Q��;͂�vz�!�ݘ�N]�(��s�\&��?��|̇�H�vĢ��%�y?�����<
a�o c�o��t���q���u�!ٴU`V����`�i�2c��|������kېg�\�+<&Nh�]|8��F�7�O�`��	?!"vX��6c0=$�vdq��=�19r8O�s;�p$:ߘ�ܾ���8qR�\�b_ޚ��N�-WI�1�ꡎ��L�'? j.Ղoa��˅��̀=�S�1�F�a[��^l��_�ݠC�p򩈦��0��g��z�
�B�$ȿ&g�D!���v�d��w"1��)ĵ��X���ɺE�B�#�����-�fV��D-9�/�th�K~I8RXr�o��c���8E�%e��3 ���3���Ԁ�5��k�L}��H�is�Մ/�yC�0��y]o�����1�t�lЬ�|��,�1����Ꭻ��S��E@e�I�����W��W�/�7��ي��>Bg�ٸ�Sӂ��y*�rHw��'�L^���7R9�X��<�%S�^4�X�i�$�Q��U0�_�*|{�� �eL��Y<L&�qo�[����C�&�u(I��ǯ�diχ������׋�K�}᠃��z�QSN��=�Ά���ѿ[
dKpV�bLԦD����Y7���~��u��#뭗�mL���C^#�G�T�ڝo��6N��Q和ʬ�԰��~�M�U��z��pr�x沣ջ������}��|��M�P[���I���Ӱ�t�ҬA���ŏY���.�"
���O���`2/��x��+g)��Sc�֙�� Ֆ�ޮ����кO���s�eI�CR�yY�](&���L��'ֱ���Q&=/9����"����N-�|=~��(��w���y������ý����	�0+O�a�^�y�@���:�ݝ���T"�c�/����h�K�v7�4��j�N�<��kD� �^��/wK[Y���Ȇ�ڗeG��.�8s=t���Ş��W�����.��b��N���N�!��/���T�{�C�U����KwP�Op-�\B��X$�F�@?��/zw��� i���
��m�S+�� �LKS���_��։�;T��b�S"V\'�&��Aܞ�
�aL�w)Ӌ�wCI۹����.@0��p�ލ�< �|�E�����H;�R��O}�7m��5%u�����CF���d��_��GX6_�XK�[qG�d;����VH/��p%%������߽<xw�9V�Y�Fm����X���I�C�mX
��Ō�U���1�dn�ـcT=�@�n��,�J��|��賥+֒J	L��*��	b�Lމf�8�)^��ò�s~+k��?^�,�����(�y�]|B��)���* ^v�v%�W5�#�� (��T6"�p��3��*蘡̈��D���u��������s�J´MZ��U�c
0��D�i�.W!5�<�a���r��V����s�T{$��I8�hb��G��L�	4�̅�;���ہ��a�!�w��hK��[`�Y,(�����S��I�{Jp�9��ԋ�D����TD{ߴ�O�$V<��ĵ���,T�N�t#���Ǌ��3o<�o�� aIҡ2%,����V�L��Tm��An��-�Z��B�"�6!��� |��^���z�n�����)�'���M�S��#+Ҏs���
��q�h�R��;�s�����VF6-1�c�v\�sTʁB^��,ع�����T��G�Y�<�u�ξ6R���P��Qzg���R������Wtȡ��9���8�Va��;X+U�]�Uh�v��#���p��9�|�Zw��~��,�ݧ�}�[1���^�t%WB�y�OY
���6ۂ�ԛ׍�$�t��%&
�((����O���h�z	�m��4?�Yi��/7l��y|���Zf��ô���+^ZJ2��far�9!0&:��~l����D����+VZYx#��Q�Eo��.9jh�ٚ��D�y����~� �H�s���"��#�J��9����$�B� ����2�v{#��� ���q��B����p��	�_҉�J�rU�f���	o�Iy�6U�<% �D���K���`�8i����va"F�9$�����y�d�w$��1so+Ď��qk���G�����65��V���*Io7K>T�; _Ђl%az�ȅ�Q824�8g�k���מ�����4��	u�9f$�7Z����;	�3n?�&�E��mA�&���K�HҺT��U�H��WyR���Z�(�ѲJr�%�5餆���
C?:w��f[^�(�,�����V��G	��-��$8m\����CQ��>��InP��Jk����K��a��|^�Q1��7�.���V�>X��.����_�p^U�.��	��q/y�O����V-����)��k�>��L�.A_�$\�����:�,v�Ȕ�%��&�x��}num��9�'F)�K�{RI�r𑤵e�ɾ�Ձ3%�|��F�EC ��߅_z�^E*��Z�\�:LB�_�q�L+���(H��pC��)Ou���Lʡc�*��<�oLd����*a��s;�Z'�Z������CG�T�;������g|@*o���}c�ߗH����k衧�?��ܗ�����kQ"�.��о�9w�s���C{Y�ʎ9D�WZ�zw/��]�E�!��=rc��D(�v��f�Xb�.�^�eb�ȋЃ�B�_�w����p�n����~���N�<O����jz9��R&0J�58����I�W/Y�(�,�!��;����N!fz7�dj�`��+�?L��ꌙ���@�E�*D�֑�@".�KYg��y� ��!�H�&+M�:��G�:T^��JX\+�@���A���C)fVᓂs���<*�QI���c�=���8 ���	A�!�e���89c���
�n����"֢�J���
2��Ƀ�
�i<���ec��>��L۱�D+����h0��C�|Iޮ�7����^���hX�9Z��.D��f��v#f��%<>�ŦTF�5Z�W�l��jt�w�`�<�~%�%�~I�etS>�-���{�|��&�b����3�$�|��"�'�#�2Ĝ�y,=i:��ʤ��V���[�H�&��-�~�>BN��\@:�"�0S4���ٗN:�1��IZ����@������(�:��4TД��i�c�xMV�	]eO��q��qf4>�#��E��Ko|��9e[�����a蟷c-R!�ٍ�o��+�V�P�h��J�[DB��¸�s���Vx��C�r�K�b�9�]����j��~B�m�>��]��[��w�IţA|��_�?�j�k�+��aH%�\�+��q}H��6�Lk}�m���K��a&d}i�;w�Z$���¢�C_
2�zf�nթ4��'}s�F������V���A������Wm��'� S��� }y����˴lВ��\p|дr��v	����'Za�Μyt80|�]�)ү5�+?l��g4�Py���/�}ոV�ld���Z��(�����$��N��lޭx�5�$�7�[�r��J&���yH�Jp��8�N�S�^`nl�����!n�$"0�zd4�aS�Z�Ks�okO�"c�D�b�W�8�7J���L������Y�עKWQ����ee�l�Ҟ9��ꮢ�J�h��m�hÖ_܍�MD�-���W�Pf�ǹ������y�|e��ᤉ�YS|�;�E���?S�Ɵ��VRiAv7�{��N�
#�yY�ϘW�d}����n-0�v��t�~.|d�86���P�����hj�[6���@5�_jŪ��2�1U?�a��e�6��� �>w��@��L�7�����9�����Rޠ�r��bM����5	Y��)�vIP,��tX�U�`���v��^ȷ�9?�c�O�np����ۣ�?皾"�A�)�j�J*QtjE�n~������C��{m�P$!�Ó�7�w��K>li���'����jh`}p������Tyjc���\|x�F�pM���
�uL٪�ъ�I��������8a��|��m6}Z2	ـ�t�BF=\�=/�J6n?�\��:`(��N��Q~�_�M�3�C����j1G1WG�U]p"H�w��c�T�ږ�?���r��E�x(�E����q�Y�DRo���p�^G�-#&�*L	)�Ij	L6��0qKhB/<=[�:�]��䭼�g�����M��1x�F>lA���@>L}~Q,`
C#��d
1���1_*7�#���9l�<F��h��s�r}�%V��2ޯ�j�TJ���@S��>�=�{u�ZU��C����8������r��OҼ4	�!6��8��b)ؾʰ4�4�lڽ��*���D� ��5zNq"z'�3ǔv��J����ѯ�u� t.��I}���y3����\���U<���|��>"f�m�M�cS���r���?�#T�;�r?�q�� �~̆?�<�IQ^#��9E��͑�s�����=-�Mcg�Ί���>o <����_�{k��$�/�����s&[��l�Κ/�=�3�wCq����x ��.�ɤ�%a(a�����#�,�?x�r���#���3#tc�"�P�E��B'Ӽ0�T@��.�֚/�#�q
�\r��aEA�s���LH��<8�q�Tl����r�.�Q��"%�ێ��X���m�Y������'��MT�i�v��=`�?��6��%P7��ͱ{W���(o�8��"���k-±�R:��D��I�WE�Z�26��0|�bs���3pvB�ew5���!������{j��Y'�w������r�QҺ�@��e�lIR�����,�lÆ� ��B�3N���uF��8�X���#�2��B,��]�u��˷���-y�h�h����S�� ��L����G�r��r`x��T���!(Y�1�E���Z�b�)��Gn���+�S�x��#镨ݽYu!�b4�܍�=&D��&�u�{'�� (����+x|F�3a
 "�j�v�� �{�=k ��>���
�/���Zt�r���,D��P��\���zS�����P��J::����LH��:�����^�r�t�b͂Jh��|*���y��@�W��n:�"!��E��[�v�:��6�;��dk���V���o�X�4�t��nV�ޱ��d��
C���^�����V���8(��e��
�+�L�os-�c�z����Z��+�>Zi�l	{��X��8oIX�ƹq���a2~�mv0�:�����u&�g�~$����ߎ@�^�ⶎ��I6�J ���� I�ڀ��������b���6��7_���y�O$�6�V+����$_B|�H :�dͭR=������H��P���LT.�M��c��3֢��$���ߕzȂA���QN����0qJ@�|r.D��K�x+��@V)쒇~w��a����h*��Y]��yԸP��@J?B�L�=���͊Q�x�"��;ϡ=!�/[��/��G� ��Ѹ�TQ�?�N�{�1� �B}�>K�.߭[��������90�G9�u���d���tn۞hp"А<�Xz������MHy��'bѾ���:�z��y�,��Yg4b���"�pX�@����9����7t��p��*�4�\t(#�'^��J���1��
y_vd^�qnwaE����dfQ9'Yѭ_b3�o��=m:uO��j��hmxB���q}O�(�G�y�k֣�lŒ]�N�� ��B����"Μw1�Q���f�~��5�DՀ��SVcsC�h�I�?=M���I����� ����p{jQ�;|9�|؇Gi����{Tt�$��٨�:���"*�|,���eP&��&Ԇ8傡��y�]xL��`3�vLz�5+,?��U���
��HTօ RG:�@xé�����L��0�N���\M.�1��M�>���x_�����I�����DҒ��l��i��|�8Jo�I|<'����S��}"g*C�*V\���b�s����֢����S�,º��E���Í�W`�ʨ�HR�D[i�߂��,��S/��}N����5Z2S�����Y)����k�M��k$��0�g���������Ȑ��3�/�EX����^��}�^��v����s4���;���/�rz��������B��_j1�Y��9�E׍��_��L�\��N��ւ���&K�|1�ƷCY�Ң������П�u���L�r�c�]r�r��0�ҽ\��>m�m�ř[~H�9=ըv����ᗣz��81TJZ�n�e{L�� ��OA�#��]e�Zm�k}��/x=Ee s��k�*�
��k����S�_?�h�
�Y����S�hT}���st���n�"�0˥���c��ݣ��}��j]N�oZJ�����{74��#ה��G#Q�8{>���g�@H:��v�} ���=ZD*�Z4��+�u�Z�L�d���_����a��[�>/0������MDX��v�6
��i�CGL�?ޠ�Z9�o����E�(�#�յ�#@U�)'�VJ��BV:��u\r{����%���h��=�q��s�����gQM�<�f9���w|�,�����4�qnǨ>�㚱���Ű9?���}Uy���~��}�:`{%��f70��F���XAex�׬L�7M�_ll��3�G�[�	�x��Xۂ
Q����l7������		]J�f�$|y�\�>`�I�7���_�-��U������!~����A�KT�=�����9��M+ iɧ|�!u��WBM��[*g�jr�`���lPA��	�խ$�v\�	
_'���َ/��W�ݕ��_�_�E��y�������K5L#�5��~��@��b�'��}���p�\;�w?�,�ώӽg��^�-���?6U�ΒY(Q��_rbr�䋼�����@��NN����T�!�W%�v��|^�]�9����Re����5�~ �%��C֕�L-�Xֈ{�x��7T���)��6��.f��Zp���^�L
-�7�X��z��JY\���\��K��&o�E�8�����4��|�\'%ĵ�I���{�9�A'V���O�0�)Fz8�녈s���r~ޟ�$�^Z�(�eI��z�el��X����]�x��m���c�K̺Q�b"�=��|��;i����������p�p�~YB�=�
�$��7�-��7h���?�B]Z~E@UE��g��̚@9���	aM���plu",O& +�S������� 9��Qp�`2����Wᾥ 遀���u�;�U��3ua�S�y���j�N�05�0�=.��6-��I�0�EN�ߟ>Hu����4�8��%!�A�*D�4�BP� �k����nd8ȫ{����.���|���eX�� +��i;���2sv\�jw�g���4d�e�K8ݕ!"e����L|�`�|6�%���YD�n�O��zb��K���a)��N�)�����Yw�E�:?���TAZ��EY,��m�0��bZ�`MQ=�w�IP�]c%���rZ��C��#|EڦC���,�=M�w*��Q�ӎ��~q����5
�L��HvB��.��~Y_�(}���aY%��,�^"�&�X���|i3���'yb�<�|wpm�G�qW����A�p��l��E���z�75|�j�KA"%�:���r| rS�?�-Gq��(@���V����r~D	�_F^3��	U�z�#�u�{l��;f�wjоI!D� CJ֔����������HXT� �S�HgO�J�]�R#� QA��8�W���*�-2���,���� � :� �+��C��G�\�����)���,r����{�'(LR{���.|��g-2��8&������ņc�K�$�p�|^� Z-�y�kB�������JG��ȥ�ݏo�~'�Ψ�6�}q��=�_�C������v��Ƕ�>�TA�?����toz��p�EVE9r�Gy�m�����DuI�?wa���M=!�n���[���#O��}� ��|���e(l��}�LW�2������e�S�l·_sU-��L#2�r^f J�fW��ƺ�R�릏S4U�|P;�>~�Bp㧖���J?9zz֑����}?���p��a����xz�E�������\`��R�SAbI�����n(�h��.n2��X�;0�\Ƭ��C9�(���Ս'Gi�z�d�U��]%^@��x�,����E��b�>���)	�pYk���Z�=��-����{]
E�EL�0=>|�s�'eUUU�ˊ�w_ѩ6z���_>�;;���y�Hς��,`:�`	��Ŋ:㖁.��y�:8֞9Q�� ܴh��iP�I���n���N�lt ȟ��/"���R� �����v<�3k�&�z��n$͘���j�N�G��Жv���A�FP�0�vt�1�l��<�'���I5׺�����]w�*+غ���Ɲ�Vfr�[��v.�`�p�˲B�y��(�Ag�2w ��*i?V��.��"�j�۟'%̖Z}^��;���6m�d	��ۍU@��
�<0�FBe��t���N0Y��2✘���cNH� ��������f�8ZQH���1�z;޾V��3�x�sTo�O��H����C�O�/�J���'�Ug�1�E��y�t%M��M.���2|����0�\��Bm�wD�s��=�5���\]=�~�S��w����݁�'�|Y{f��)A���� ;�	ޅ�����ք�yR����0�J��놅K������g��'�&����:y'��h�k7?�u�@p,=�$�z�� �$̣}w"��1��f-���/�:�Z�o�����,8�P�8�\��C�<�OV _�~G8��)�q����#���2�!�x2�UÅ���§tdJ����������Yb�����&ڤ��E���3�i!uf�S��-O�|#&���Ka���m�hB�.L�*��*r|] ����Mt�+���l�}���z�@�rU3�zY���iF�ٗz�iQ�(�	MV@�Q�gs2ڍ�!���Љ���>�7��2�l��tU��+zrPP��������A�s��)sP�xLڴHhOv�W� 4(1�9�q�$��s�tC�Z�{&w�`>}N��������P�ඎw�>�m濏esRj��+���!�>H�Ab��(������-D�u�9�C���,�X��\ R�Ov_�!<�|�O�˚�h��m�����%�{��r2�&�8�t��oiŧ��'.�(e�-��kaJ�$z���W�/�?��uvaIt%���l~�h����z@�a5�.�`��<'�5�.B#�I�1�����;�� �Z��:�t���#(;0�i�M�$%����#x$���x�9�Ʌg�n3����.Á��q#�~֪֒�zH&�M��TƊ����HDN��p��_�0/2��Cx�E����� ��v��ֺP�����G���<	��P��X�&��I�~|�/A"w�T��N1����ҡ�V�O�.�g�&*�ܪ�xts�p�Y�L;j\�y<C����y�O��A9wԅ:�՛w�JQ��c�[@�
���J��xӏ��5a��uIEtݦ�5�M/��<I�i���6\`6�c�a����T�K����'�w�)�x�Ź*�+�G��ÛX�*E�剌\:�=�����(%sa>g���@�X�:�[�TW�e���RB���'� 9R����D�ڻ�@�\5&�����m�1�x���?�/�X�F����Dŝ�s��ȟ���_5N���C]��אq o��mw�H��a�v6��p���9�v�b� ���6]�Bc�QM�.�N��H�$b�0����77��9sܰ��y�b�+W.�~y��z���\l�R2k ��x�o܂xw�/��S��ʳN�b!������y�a��=�[���Z�ǽ�WC?�A��:@-������d��	�<��ڶ3Tw:{�X��B�b�4Q���p�" Z�w�=4z�4Q�Â5l[9��!R"O
��kI��V�w�� ��TS�{�ż��_�딨,�%n�@9p�(4�I����B�&�e�{�����/����� ���):�ڝiT�9��I6ԯ�AB�(fKy-�;i���8�O�q�PD�:S�q!���yQ#i�����xN�����G���V�k�+.Fn�!�7U�z�I�
��8F{����U'��v�D�7��%(];jbT]	�CmK��tfJV
8/n��q��6j{�ܼ�$�ZU8��lz]���2�K���V1L�c�/]Ԫ[ٝ�mb"��O��"��X&qfj�$�$9�N��WY�;YM�R�W5 ������L���A0RtvC��� .s����>�� �H��e��D�X��B�G���?RE&�HV�$ӷ5�~��4��&U���I�d&�Wx��JA�����grTՙ����O���L_7w篊SE�#+?���%x�����i��l�H��`����ṭ�R�ӟX�+�Y�G��I�	l5\�l�#�J�us<��&�J�ؠsv��/�ui>�sm�4��{UMը�Wg9������6{δǿ����.#��-h��#�`�����t�t��^�g�G|F*K�j���z@| ��Ï[a�d�z���'Fjk���풵�[���2I�g-FxS�춠�1�z��@74ic_��������w�\r������h�v����8�J��k�P�y��Xc��՛�Tؿ�����
b�\�V �~��ꫭeF)�h��]�2�VH�b�ֿt��e!����Ls�/a{����Y55X���q�,<5���$�-v,�[N�"؂z�ֻˌ&j̈́r ��3AMPb���	��7���~� /���zqc�
?��~�DWYfU���E(��A`�D�V��~�s�2H�c�2�>q/��S�����F��G�W��
Ҵ�&,���~�PJV,�X��w2�p��ш>0
����om��]k/�__�)�e�1D�t�;�֟*�Ln��GW?%�������\}��U�#�E����;@o�=B3Ѽ��/��V�v/�ͅ:�>���� �x�J
#F;��"a�����#��;�L3a�M���C��0��M��Ƥ�	w�bDN����
�L�q�-�0�/(��7����,��?�����-@W�ZOS�6������v�1c���q�����,�
����ֈ�K����Uv]R��y��ug���$��@���ٖ�S���n�����?�I\��1(T�H�U��
|oӚ��Z���S��^����w�����@�@��U���Վ�	����Z����2�RO)�@,�գ���W[FX�w}g��{�x�SIa��eLL���B�f�3�tз���R�/� �`/k�K �rZe=����o-D�w6)2��^c;w깽
�Һ����f`�NB���~�>Z~u $�=�S�Za��g(����)+��<�-�6|�i��@ڟ��F8���Ӟ���9