��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨס�>�6a�
�Ys����'Gc�$��@	[��%���R^�/�
�S`�����r������qT�AGe4|�5��Ёhӷ�c�F�ZNXgvC#R+� @����� �?����:p�%�Hl�-n-�*�:I����j}��<��W�g�����0d��n�i/�BʩK�^Ĥƪ��X���D!#�6kOT"�s���3I�G��e�@����� O��)�_�%e�0���<�}Ar0Nm�@�)��iy�uC|�*{���:g�}3|�J�]z?�d�=��nV��e���
X�������A�Y�D�m�*I������n�F�w�d㇌���RS�T��6wi�F/������O�l:�'�&ۜ|Y���e�r`�HE��Ͱ�������*!v�i��^X�d�Յ�5Ԇ��gJ% �n,y��1Pț,W0�N"��4ba{Rh�]j���ӑ�<��c����@H��,��|�ϱ�SJ���]QMd���
��I��w���Mu�]Q���L7�����W�������kj�;S7u��,x�C�Q����ָz�ָ>hАS�������M���je�n�+�������lk�,_�pJ:@��� �j��J�=;��h���u�l�
�v�����r�ż;Nv���X��(Ȍ(O�FC�x�G�fɥa�*�~԰����^���!�R�,_�cj�;�p����Y��_���u���g�Ц������/8R�hcB��>��1J�C뜂�\N����?�r9n)�(%����ZC��J�i�Ъ�cz:cl=��t$TMB�K�*)��Tg��(g�S�6q28�rG�+��H]q���Vh��kB^+r�m���)�vb
�D2=1j��rz�:S���X/Z5E�G)��=f�SCQN{�~Z�fd��z�,�21���K������W�n�J1�n��?Dֳ#�w`�g��zZ����Y��2E���v������Fb<���E�����C��k�.O.�W�l�w�_(�qnH����S�[�7���ڙ�s����B�U�\�T1�+	�A�ي�X�+1��y"�M���Q�+e�:n2�آw���nѺ�)�൮�Jb#���c"���s�?Aw'��<�?�W-�1��WgIA��'��y\# �� $�v�D��b�(]VCA	�	1�-��)�N#�� 5�Mq&wH����2�o+9z	j	�����_jU^��ޭIL�=��������қx��o�<q��n�!Mi�z����vk~|#@��L��2u�,ui�/'�z��P�Rڤ[�N���Ǵ'�?k��[B<��?�G�I�b�h�w�!�r8 ���m+�3��F���E`▐��M�$<����c�%��)(����L�z�FY�{�����Ac!�v�X'�xX<�����e�~d&���uNJ�*�/��G���:2��ff���x��Rd9��T#�;�*E:Vb�|s�E@�Y�7D��HKl$2��*h�58J��7�ӄ�q�~ڨ쟯�C�(p����#�d�nA�Rh�R��b/,�Jص��[���"����I�j�C����RB�{�ty;�TWz:~A4�`�i�z��7�P̂��sFLS��GuE��/��4S�9.2���1<���;�SL��l�bU�x[�c��Uj�y��J��޳�?Q���YnX �hf�f�]w1��1<�W�r��ĵ�g,�.�(���(��n�-ov��(Q�ԃ��cB�`�ˌ�-V���&�-ѱ�qD�JXh����6��8�r�V!,&�H�d�%�2@����%v�*d�0�`N��l�2Y���]�� )��hE�_� &p���D���$w>�h�X��t��T�컉+�Ћ���m�$"��Hw8�Go,!�c�҇�;'��޽RB畱\L@	!wBmރ�P�t*P?��+f���g,���4;Qi]�-ဝ9(�ZjUMA�ho�g�<連ξ���\^�!O��m
%�Xj�q�t�d�2.����#��}��|4��(_�\�Ւ��5k`�Ґ�QA(^���p�h�	S��!pF�ΪY�?����0���>�Ay��~�I�����s)�x�V��x�A��W/�J&v����zpVg�X�(��#?�"���`x���>p.����ھ@1y=cpG�Ş�lU�����I1_.�/pM��@�)<�ʚ�S�����%�s�I��nؤ�~�7b\�/�{�P��8����/�YM,����+���^!��M���ċv�NŚ��-B���3�`=/��o����2Br�K�.3c��8����]��%W���%��&=3D�}_���� �&EG�� ���/%DQ�3��q�[iOM$���l���q�R *麍vV��b/�[H�v��x�	�p� �����/%C�R���F}�3C�G��*_74X�{O�zwÿ�t�_'Иv#��Z�Y�1�v�'��C
���GLa����aG���a3R����0�̼'t�H�0l���bmy>^�g,GɎ�M¶Z�@M�������.�"e[r�S
�R��v��T2���J�(}�/󊮐��*[/���o�'��	�y/����%����g�G�Jd%[�m]Bўɥә=�NZo4f-��L_i�~�m�����/�R7,^d~*kl�b��:���g�ibm1��T��AW'�����<	���!P'�Y��������M$�W
�?iz�&��,�p�NI7/��)�q`�3���J���$>�tF�K�'O>��5��I��n^9K�&�Τ(2��֡�W��]�Ǿ�QNP-e��A�����l^�d�J/��ˢ�nt�.ӝ���13H��u�ꆚ�3g�CT�A���h�@p(CW��cE��ڔҺ��T�x�>�����Y*>[-A%�$�8�"��<�S� i7in����ٮj��Z@+r{�>>�?��Ѫ�O� 9S�3���|��q�B�(f7�DZM*<?�x��/	�~����9Z:ȣ�[����VD�{%�e!ڰ׊�NF#��˛��1>5 �ȇ�&`��!�֕���5��U�J!rM x��PA4�I1	���/��N�(߃8}��Ӂ����e��{q���k�~ax�L߬e:8O�}���M�;�6ڴ�ߡ4�.F�k1�'4k�5�7{7/6�G��ꙙr���&H.w/�\��}��p��|˓Bd��9�vQ�h�V��@�5�6���Af9��{��,�j�}��'6�z,��
��S6������Gr���)`Ji���Z�û���pzB(��=jyB���ܛo*�>%�)Fpc/�̈)
{�N�8^�a�Dp�
2��|��(�g����	>�S���-Z�b�o�@D��U�=�*-۲�����w�E�*G)"� o���awa��?�We�C��?��oe�)�7E�P��(2��X>�We�Yj�I��Ҝ�I[7��Rh�\�T2���U�>�7��r����&�# IXs_W,%��e���̘�:��t�.�T;���q"�(�o�O�}��^#=�6�p����42������>���@�@�g	֜Z���8k�ܢ�6R _"����8�PG�G�TkZR�˨�5�I�j3'�����9-Y���P�؂�&O��B*�U�p�]�j�oO�437�W�|� ��z�Pg��Z<�F;�/���u�	#�
N�n;���`8'q�-Pӎ�R.��R�c����̝0�ɋf}���(0o0`M$�wk���x� �ÈS��J%grUC�x��42	�I �`Rn7�p�`l�M��_7�z&�`��Äd�//�,)���Xq�OH+U
X��O��ʆQͱ����k��O��:,�����r��y�P�E�&,V��-)g'�Ͳ0y#ב��,Д?~��Ǎh.\G��}ْrk�3͓A���k��oC*cG# ۾�����T�y���T�I���x0m������2���/76τ@l�_F��b�N�>)�����F�5^E����J[0!W��U��$N�a-�<N�}�E<ߜ_y�<H����|~ttPB3��ޓ���p��X���e��8R�b9<��'ڃZ,�k��>�?�ǵ5�4�<5l�p�+,�l��D8�U�R�)��F�f���m�Uʘ���ߘ/xgʠ��j�^�o�i�+��?$CG<��n2����2�+�O��&�/�w��̤�1�(K����45B�����~9k����Su����`�P5͖.�f����_�S[��N?��>���7#u9Q��[�U�g�[��Z
#'Y���֋a{� ;=C���� ��۫�.]0�;��U�ښ0���^����!�EC�n�G�D�4�QI����/�A��I����',���1�-�r�˜�TkO�螮1��e]�i���� Q7ll{�Z,�3��n����Jiם�^�0�tK�C�3=`�¤�*�_#qa�ti� �D���s�M�6푬��Y���̓��c�F����Ld�o�;�5�s��vk�v����CQ~8=�'*m/�)��(+ac2L�:���y9d�;&��{av ϨeAW@IAg�x��B����6����.|u��\Ȋ�	�v�z���71��?��~z3x��̊�ly�;j>������?�('��ɱ60�l�k5��=��f.¨ʒOK��s���k�t�t櫁����'�..�q�;d#��_*�=�\xE���di*��*A`�B�v��ӌ������l?�I�:ӥ��5�zx\��Qq�����t��ݩr��w�)(���0}��F�8�p�b��P��9>U�n؏�(�)B�����]ɦ��rY�����B��BT��Y�D�[ǔ���M�4V_�e�������	e@\;1RFg��՗��:��Z���!tݎ���U/��7L4E�ڣ�Ԫ�$U�pGF��D.��{�e�Z$ ��6>�}�װ�^���a�<��O�7�����q��t�<>�&�����!%p �߱H�qp��PSG��s��Jϟ�04�dz6�]��e�K��v����Lz_d����
��SզrH>�s��`��J�D�@��zaYk�����4���w�tσ�W{�ɗ��g� #���?�7���:���TF�D'�I�Eo��9�l@��
$T�i�ɨ�