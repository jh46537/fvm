��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�	�O���T�7~j�K�e�rd�nWWg�kKs�<X�@�U/�T_K���/c�N:5]6�)D-&ω����t
�\;�E�N]Ym�o��|=��~��=׆��۷�_E�� �%���X���RC�ߤ%\3��1S���m6�]�XN�� ��/�l[�S����,dd4c�]�n L�#Qc^��@�K��3\T)����ny�Q#0g�%\�6��
ņ@�<jG��zJ�8�oA���W[���箢�3�v�#�3 G!��}Y��q�s\�Q�Q��j���!"�v�b+�aF9Q������N@�q�� h��DvZ��f�
��\k�����ec�U�Et�y����)3WRzW�s�����'^ P�D35�y���p!��gN:�`T+n�"l�m�b!%pt��|�ћ��t+uf<���_i��"���7A�i{$�Z�=����� ���켁���:��i��%��ID݁Zz��_J��U���H��9g���0��N��/ΐ��Fη�$�u]1�3+v���y���8�xY��;�5&Џ��)�O�Y��8â��O�aB�dլ��
 �Ju���Hk�k��:�/"@�*�	~��H6���ꋀ_Y��!t-�(6��*��p.0���UmE_�V���|�z�5i��:]F��~���I�g�Xܴ�=!b���>���d#1@2~z�úX����`A=��#,[5ޙW�6[1Ǣ�B��_%5�Cֶ�QY��,���5qk4n�Ӏ�U�<��C�\��P����%��H�,�3�+WV�k@~�<�b�!n4��|��z�����5C�ou;z��>\@SE�k�$ado�P�])Ɏxõ��~$��a��m!*��d�@�;"ɨ,(�0;1��^�VBki��x����{�J%�t0a&�b(��C�T�=��̝h��<����N3���O���G@Y�^<�/[�b�˲2fb'���׾9�C�UD7D8����D�r"��<�i��ljx�]��8��{Z��6��/�M���&M��W�mx�)�X�:g�=?B�7-�i�Y�Ϋ�����/�
�<g�6(�}?/�ˬ|j��H~�]#W�-Y�9���tP���
�Q�?4?k�P�ǵ�4:�:�F����

�M����;R2插�;�L^��Xi�!���s���x���x�����d���Cб��x�Y%�#E�M��m�<��XW�6�3*/����fS�z�lZy IVS5D(�
@�,��C���z�������T$�&	�:��R+���X��z��ɩ�|.T��%^hO͑��x�j�o�|�A�VX�b�:�EeMQh�������l?&���
�P3��2��D���NG˾�j�j�Ln��M?�t>�gu���ͱ�R�w���h�$������@�>�9�G��A2����?0�}+�6c���.��<�
&�W�)����xq�<\��)��Iy0��/n�_r%�d~>1� �����2M=�ɩ�l��#P\q�)���V�n�5?���`T�����~#ߗe�]�Cf<�A�K�A*�HA'���Ea�a�%"�������4�%k%6x�{>
v	�<R� �vN�����AD޶l�ϝ���}e4K̪ޚ �i��Z��I�@t;�KSU�M�WsH6e&T�^��Y�$
�PAJ�5�y�����ږx�}>Ѹ�g�IG0w��v��I�$�r����lں�����/�K��wZ�ahh0wYG��;@�)�1�p������mW�q6��k�j�v�!*
���]���B�e���]~V=w/tr�h��/*9]|�Ķۃq!���sτ
s@�߷\/]c	
�F	�;���>�V>���V��9�埆�Yz�����n�B$}3g�^Kn_5rsS1��{�ӧ=B�"/���ܰ��a���'�U\r�󘖀[lC�;)a��|L���[ϳ�����e�oM�d����'b�RW��a�B>s�m��8��J׏0�C�Ʒ��=�t�98R/�#@�R���0�w,zr��:����K�
Ohu�B��uE�F�P�U!���}���R-���n2aEt>ٗޝD��Y}�dt��0A2�N����s%�Q� �=�,�슜q��E�&��@�a�V��/T���6��āoX�P�g���>�G�c)�V�,��h�x��e�9���:oJϫ��,!�R��r���I���95j��d��=`��#��YJ	L{t�Y���鍷X��'tk��<��H�\̗�E'_��~.��Z�>$vE��@w#k�qꕋ4��Q/t�!�;\���28��-ԣ�2�V��"����P#l^a힎���$�?�����cZ&jO���չ���j�1D[��{�k��q
��oR��1�{:���S�>6��Q1�QY7'�x�eJ::�z��:��@�Q�+�?�G�mT A�%/��ݶG�N��jf�=	�X��-ol�7����Ü�1��bp��g��`W�k�|�æ�c���_X���i�p==ZP���Z�Â=�o�G	b�����ڃ��W���f���D��f2l�㆚�N%���/����^��{=�k~�@��8g��[�Ɇ%s�t�f���'�}2�3,l!����ٔV)Ty�\�7}H�IMƎ�������;��R�N���gRisE�?��H;3u_-h���N{�|��.1��h�b�`jȉ�\¶H.��l��p}���_�4}H���L�� �Q������b�{�1ZXQ��v�s*K����o19l��+s�iU���8%$�M\(@��~�7`����&=�g����^Ic�Y�x��AR���tʩ�(��MFႮ�T���6�J���
��K@m�:�����ⓝ!qp-Q2�Dno#Q`�Et�L��`����~�f�����CH�C��c�~V"{���I8��[
64l����*���7݅w�-��~����:7n�{���
�iܩ~E���o~���d�H�48���������]�P���*$����M��Y�?��:��]jf;njf�Y3�:�n�N�|�(��l��^�f�晆�5b}n5���:��GّZ�?J��e�˳�X�*]k�Hw���z>}��
?�Ec���h;)�z�������J��.Gk%��wgv��O!����_��
�w�3Z!3x�3/cYI���K������a�d�zEh����μ��Dx,U ��$�e�_&��VAhq��s��ڌ������h߸�ZAM#>)pt˦����s��!QE�J4�:�1��E�Cg���U���+$���u��"�����t�������knZ}"�������rm�i�<Wvp�5h�*���7KF�\���"̦�2�z��x'�tֶ�dW�x?o�H����)�㸗��qQ�)�Hf�6̮YTr�+y�-GX��~���5��}���z��q��a>u�ke�A� ���3���!�L��'��$��G�{o��.�U���~&I���1�)F����C����'V�W/X�V�x
�%�&*c�(a���iR�ftѐ����e�(b�4n h��Ozts���	L��R�G�zp����f����&%B�Gխ���Nd��s���h�.4F�j�`���������0cW�1����lYݒ��������@�r������Z'F+URi�p�L�G�dTu�����Ob��Ie= �=T��̔����ӳ�}��{yZY�*�l��v1;���E{�j���G�	E���|�w�Ϫ$��>9��4GbK��x�����n
~��G�o�3sC!kͬ=GG�#����-��Ul",�\T����0�����u��]��E��?�锣s�CZ�$����Yf�C��~��8k�`:l��]�f!pp��i����Kԣ�6AM�KM}�ۯ'^	(����h�b�ƾ;|M��YN�#�3�[���;�����tm:_�zg�H,2LQ-T�9q�b��!���G�A^Rclw>�K�NU	״��j�W��ױ'
\���`�_e�X�\���B��wX�`BUh�!S#� ��@|L�ۤ��4`�\ޙ!7����Ί��	��	 ��B  :��,��%�E8�R`OH�3�5�,1Ҽ����w�����`׽���֜�=�D̡� ^��@��.m�eѠ�^bMúE�/����N��6p�Sԕ00��R��K��K���� �J-8f/�[͢U��_x�o[��g(���\Z�x�������.����K�`��*����ؘ9�M�19fj� N�����}W@Q*��{AU8��#���§9EV�J.I?���<��q�93�"~A�K�w/H�SF� VM����~9�%�Hc_j�W���b�;��(�������
͜	L�^�x���#>@O�ZU�=��v����T� �̅��E��aH�-���)f�-,n�O��~�W��DDf!Oa6�Wg%��)<Z�����F�hf4�%�.["���P���W9�M�=�������<%#��6<���T�ǰIo�̦����iT�� ��W�hd].L���K:�0b9��t�\�v I븡�o�!wD�C���M����^Hqc�/���:']a��q����ӬqP���mC�E���7J�����݋~�d�_uz���uk+���L�S9�m�6P���N�J��91�c)3��,��`k�a�RxK-�/�W.AV*���T�]��5	3L�Ѐ�����c'�E�(J�����@T� P�z�ukz`V����f�@��O֮��ئIj}g��)�8CUw��ÚB;C�ڹ'�3Pgg����T*�H"+ut�J��*=�i'���&������rH��N��Z��Ж-�WV>;�a�Ch�ѕ�L���6���͇�a��QI��܍	��"Lq0�k�#᾿�����]y#C���ַ����̯�1����-��&���ݢy��7ǐ�R�t�_v����BA��,��~���֋�kql�?MG'V��gt1�3�_juJ���3@�H=r�h�g��p�ҤaQ+��Ί�F��Ho��W �+�<�7(-�e@W����zWWK%ܖ��K�|�pޞꝝJ����+r�W����?ᓬ���