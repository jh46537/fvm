��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħP	�(<�%5,i v1`��;[���({�F�G��4�r`�:�*���\"��f�O	������O��Y��(����DV�Lg�w|��cBOb�]�����ЂΕ���!�gy��&�ɀW�0]�R'��d�5�pM �0դL<��}�������4|t<��o��D;�����᭹�^bA|�.NnW&U����?����*�~�:ƃ��o�O`�^����8g)��Ц/� ����2'Ǉ�]�2�9$�Z�6�9��Ve��pu-����=2���7�ޟa����a�i�0��!d��y%W``�\����HG�h%�rq�q2����tq ��g3�#�?n�L�l)�I���-	jYA)Z:�l像��21���5M��E�!8Ĭ�L�3Ed1�`�.�<)�eԼ�f5��_�7���?.��tv-;Mx���>���ؼ�a+����mb٘oRi$�J��<. �jJ�\~��ͮ���?����f �~5���l���|�9�tW�:22���$�	����J�� U���"���q�Kl�5��"�Xܒ�=>�п�'~���9�2��_?��bF/�[�t���e�8�v����U�E�k6Zd�V��]-��s���N�p,"����O�IHg����u7O* ���[}�����w�cי�(��r\�ǣՖ�:[�n�'a5O�����N�'M�f���%���50JYJ	�E%2V�+q`�!�{:x�7[/u�=��&�@��S%��p�z�}�`��F��?.��	�o1v��XD��nmJ5 �w��X���-=��Z��^�����+ ��E�U�\+������e��bN�Q݂�9�x�������*��Qz��좚϶ܐW����֑��&SEP�Ƨ��o���kۙ[a��#�j� �(7C��bg(���.��e��A�������ޅ��T��M�:�[(�S�c{S��Q%A)�[B~9�яZ!��?��|o��prˣi�?J �k�YI����DOVQ<䡍���H�Y��'oOA��ˍ��[m��w�\����,�A��۔{��Z�[�����o��uh�^U ���B\@SF|�S������4p��1,�%+��t�5F%d��8���KyIc
,:�4�6���	ii3�M�����òh�[U�Vq���N�_��&�w��]�^H�vt�/9�!(�+� k�8��Ti �:&?`ڔb=Ĥ�}�NF�>j�z�?0����j+��)H![��;���x�y|���/�='�ŀ��r������Ds�S���!v��w
,��/ò8�Ϛ�����r�)�:�s���t� 0�r[�鞌K|�Ψ��'�_9Fn�-X�&���o,ŷ#����
����x�:TAb4�-T��6��0li���OHm<�8�=K
�9d�@1rt�\���>!�g���I<�:1?lb�� ��W�.]��n���ݧBKmFd�&��azU��1R��p5�~q*�E�(�wU~�xr�i��N�;����\�A�]k���Ǥ�����ّ��R%���4۵��0�u���*�(��/0O���7��ۘ�cۧN&U'vx�d��bJ�`6U��ߋ��`΁���m˧_(g�[_C� �h�['ڇ=��&�yH���Ǎ�ڄ���X�h�9�"�V^s��LK�N�.jBc�^o��d+	��&�S��Ȗ��V u�ZYXS��6\�ݪo5��Ni,�1��׶o&�mH=~:6�S1zF��ɇ?C�L���2���󞀦z	V�Q*���������M�&/~1 ��aƤ�Bj\��&P8�?�+�OH!�O3ϔ=I9�v���dr�ɪt,j��`��1_2��F�����Q�N䞼�
!k�_�^!=����d�̛��	��Ǿ�x�����Tgl� �V��`��f#e>5�#O�-�phy-ލ�������!z��SI2sg�(�?_D��@��zܱY��D�K.�����e�jJ:H9�*��V%a��K\1�F��~Q
*��C�c���zȲlmo��_�}�Y�I�a�Ƣ p����]��ɋ#R�b���aYrD�0��\����bAA_N�#���I+���xA�!u:h�K�CD��i���;|d�gb�W�5�P�=q�M�9Ņ�?�P�1}�~BP�ݏ��x����;wiD���_Vx�ո�$\i�r��ޑ漞C�F*XTJr$�6 �L�}G��w�e�±�vz}�F���NT� JBڟ�E�f�.H`��;���S�G�3��R:Պ�qM��
�0Hl���|CUiBҵ��K�r��2�^�ڈ!���,(�fS��jQj7/�3�M��,���j��4��{W"|�X��@Ff�R�|��̉����cDK����EP�J�g���V��xz�)�vla��6���K�N|4���d�lE�- �o��C�E���Ò`L�E,���8��U��Lre�y�����9�Sz �f!��F�I�ڪNJ�I��y��"��|V�O۪�� )�����n!X�M�1PR?��{�蕠��~����wǆY��?v�>^T�8��=w-���0�����
�&�a�ƘkJ�e�/iLKa���w��R��6.������?ß�mcqG�܊��s�g�jI��b��7�1v��;&II{ho92R�'Ɲ���ק�Ȳ����K��Z�L+�9�%������}�G�n�x�������k
�\�(�����<�>��� ȇ$\P|�o�&E��4�y��T��!W��W$Ę���ۛ�U��id��}���T-I��-���!����&����v);ѧ�L�A��=�(+z����Q�k����;�����h]����?�a� ߍEz�&>�����=�J�
�!I�Z�n�ۯA	�D,۾,3&��9����cY^p1�����xԪ�^P|r����+����T��� (��!:0!j�TPS2�Ә2���YŰ� |�G�.¹�X�8�I��չ�^�9<UC��}_�WH��ȗ(A��.��. �Q��uZf7����$�B/QFᑧ����&��
�I	ꇮS�IV|�ؾ
� ��HZ��9�7���*W(���]��Y73{�S�(n�P�5u�r���[�s�Z.�u�^�X���p$��n�N�?�\0\�lj����Ç��Zaϖ����$d}Z`%�<����g����Ә	��g�T����9�/&ѯ���#93����� *�G�f���j�d�Y�wy-�d}���� ѳ�Ⱦk�[����Mm�ËjN�tp��R�O�G�~��!N�C�X��-ʕ��������ڡ�@�WDj�C��y�`�I
�7����o��R/	�=ro�ހ��д/5�2��{R(�n஝9(9J�6�~�צ�=i��R��S�ȧ�.�VfĭsV�{�$$���H�!&|��[����O�c�v��r��������;f��Uh��ae��X)0�=��D0檨∿��ɛ�� �@������PyȮ��KώaP��&C�oZ�3�]����j�=��@�����F�l�U/�Oz�oG�����e5��0)��������v���M�G�ѽp�ہ��=��?72,�ξ}t>��f���܌�e�p9�x��q�Ț���',�*!��:��rӵ��rc}����
��U�3���Њ�,<���7t�+��n���I@�p��\r���,�*�r���7�{@�5&��'��z{d]�k͟s ����|ɷ���
qt�+����Б,��Vm!���dA��ٿ�x��vC��l��8C�.*����u�+Q�ݳH�
[��z�a&T�?6�-��E�q,d��%*�!Fa���]W��-mz�VLw7)8!E�7f�����D�]5��9��⮋�*-4,������G@��.]��4Y'GF��5r�+	.��E��A�[��:�>�
��E��NP+�I�8M��-�\�DaJBON�.B�p+֐<�K�xusk.�v���ބ�j�r����%.< B�l�
;�hFF��݅W�Me7Q��{'>߿k�W��	�J�'*6��:����v����cuq.v�X<�$���I�efj�utY4B�y��N��[��
�ҡ��Ks!�Ԅ!�Ni��x*�P�,ԛ	�t��)�Fn}��1pb�ٽ�'��!�X�!���y����R�%�dU����V
�8�#O����R�b���ބ�����<��a�����s���x�e&Ӂܜ�H6vD2��?I}J*�/;��)���L�Zus��3�%�y��
�ř�6�m�Q��&�j�Y@��<��UJ�)u��7����öQnC�f��̬�� �ƶ� lL���p��h�J�0Y�����-D
�Fz�)ZH_���g��K2/��PoyE�v�Il?��w�*Rԡ\"�k$�/��
E�a�b[D/͌��;��Z�S/16W��n^�u���]��B�@:3�-����(�4��L�,���z>�#�Ek�}3��6���H��"da��
�+R�(bၰ�x���Q�&���2� %G <F#Ի�U��X�MJЌx�i�L�u�7}e�u%�_7�[�cV��BK3��+[?2�����mO)����ɒf�4�9-�^|�:��{I*!�v��h݊��t�2g�Z�W\3gӒ��:���8;i��q+�ֳgj6y�|��\�V����s�H��.&�;t����Fxz#DR�bv!Z�h7<�H��\�#J�K2�t�s�Vqs���F��ym-/j2�!��.�Ӆ][ٯ,��~��m	���
{��3�y�����!��ca�?�ǅD�t2����k�����{v�����]k_&�ao���N��O���>7��#;�7(���GBqM�R,AM��j��F��D� �����	f1F�3h>���X�n�ϱ<�{QU�6�a�g���E����ۓ�����:F)����[�Kb��;�驞p)mG�f��/tZb�k⳴% "�'i�c����� AͮK�V�̅4�m�N�;���qt������]�,�:����������4B�9E��O�4�/m��̛9i�A�Tw�Ls:�Ԅ�ќ��l}8ύXel�(N���F�W�Ň�UsE4ݶ�	\�ʚ�q*�'Mߙ��m��K4ZA��w�X���V���Wr�	,7���� \�oND�?��x����C�[j9�$q�g����_[�Ic�����F��L/��f^��gV2X=#�y�UV��Z飂1����;�y�V�XI׌�ر4��wyoԟ�����$�t
��}��B��|mB#���W��=Ԫ5y�*U���|dB�q��6���N� �K��a;���
q&�z��A�JHt�����#�/�`~���e1� ��'ƀ�OÍ��s�\Q���n��k��j(*�*hS1pWr��-�_��e�����r �Ls��1/�4b�l��R��K�&����b��X<��Ŝ�F	nN:�@4�!��|L�	'��=���gEL�J�穛��{��;$�O_P~:���w�6�â�3dN�K�yϽ?Gd���Ǎ
�}6J8���ƢV�h��F��u4=�*��*	�Ư���37�4ԑr��&�褝TRkG�7��5�/Ԧ0��rK��9��eZōXE0^����P�Z`���ER���	q�f�����q��A��O)7�*���5�U�������.q9���<d�1�?�s��������1�
�����r���JP�>��ZKD�f�P�Q����:z-lSL��#�!xˊ?�fȜ7��&T¬��$���P��u�Re|���B�M�1EUU��S3J��t�����X�������v"���,������-$�y��1��D�4�6P�PPyV�#�4�h���7c���Dq�
�Q�y��{��dm��;;8.2?1�#��	�&�L�8S���E�nр�a�ã1�I\L��toc}rRh�ק�6է����C=��Q���B�R@�k�ήD�A��Pu
�f=�CV��w����Y1��=�*>пX~�}��6�ch�\�r���s2BE�p)��b<��\� �@2{鈡4g|(chr��aX��^0�A�R69K<���̯�36����}��nܫ��qN��:�g�<[�����Ob,*��v��!<�^
n9�6:G�[�#��*�����$ո��� 	�$��䍤?����O�[	Q�|��C��y �g_@�g��K�Jc�� ;"J����<#-�e�>�鋗1�@�a�j�� ��ˌ1{EL'��SO��҈�'`a`��T��f`�`�\^���O��;-�p�[�� Y��gRm�r��5������0�kɌ	��K���R��Ri�8��}�ZH9f(F���ȥ�Yw�ֻMK�tyd=���y��tPo�_w�nZB|doPg�_�����:g$r\x�2_URy�.F��1d���z��D�Q�QQ�ΎD!$p�l��x�۔0�m2��Ҋ0��+�V�O�q���;@���H��e�X��Ţ�ϧ`��>��d�3M�6�0B��CFˎ�0�����Od���.��l*E��v���Q55�2����7�|y�	��@���Idw���2vc&g��7�-�ͬ���k��bOQR���e�ɿ�o��>(������jA���E��7$j�4�
M�%�i��>�G�-��L��W>r^%�B�̮�Ƶ�A����h�ң���H�ټ���&�RY�i1�hB�3������"_���iP������Z)L��\ (���i�K���A�Y���>����.I(�}AŬV��5���$$_l�u�}���v�rh�M��K��jC�����"ם!������#}�� wY|؅���9ӟı��k�
�����{=�Α 7���+�"3�'����e$ˤ�6�!~�![�������������g ���>���`�â�hڧ,�Z��7qsa��l�`_d�{�b�1�&����w�.�Y$�aaGt	���������Z�x_�^f������`\-s�o�5�T4r^:�a�Q�(TÉ@
w�7\y�0UNs���8/�5��;�P�3(zi+C<>�2��lH����n��M 4L-����R3�HC�n(5W}D�X�+h#
����
���{0�
��=�g�a�؁'Ԉ+�3�D��r����^�4�y�����9��N?{Pύb.�U㺘��*j]�'�+L��&&ƑxÑ�Y�z�{4�s��S�o=���$n����~�_��÷Pt�C�n]#c��6Q &apQvpӀQ���n��o��8`��,�s�J^sbh�f��96��0`c�������8��@��;�t@椫�}'��O݈��V�k�#1���q���?��D�<�����0s��u�����79c%ݠ��]`i�r�jӕ$�gW���BH�h?Ha���>��A��R�sn�Q�S��aĿ$ӏ�=�����k?�~�C��Sl�+tz���Y�],,[�q¼�Nn-��<k͢�=����닠^���
䣐rX=q8jD�7)mἊ�4g��&;��>DaE ��)�}���w�����@�l��ҝɘ3��6��������$�G�2S�ile9��/-oK��I[X�q^	��$j�O~!��l֩�mJiܑ[ �l�T��9X���U�-xAS�*��i��3�l�D,���s4�_�&�!K��L	Du��G� ��4{l_��k^�EO��q�-ѝ��N����:c�4��p��Cb�l��G�/*�.a�&�E)mC_,AjK�����kf���NH8�5�Y&m�+�U��K��$�I���^��:f)�����4z^�cM��x@���k[�+ B���:����Oz�`�q
���5�a���mtQHX
1�󋸎(�%�R�{��d2s��	�K~����/(�#�%4�o�xb�lx|����k�8/���6��D�C��c�u�.�r�r��#K�K�tl-�����-���w��SV�R"t'�_�5w��1	������b���9���3/EM,,@->Y<q	�����E����T���u�� ��U![̎|���L��S��	Y���;�$�{fC��.��FY�6����>~���aF.������':�c�4�yZ=P���ΣXIJײA������G��u�^�����
��I���ջ����'���z��)`�y��2��C #�%�-�(n��/rT���TP��g����[����QO�ܽ�"ʶV����9d�e��1�^q� ^1%���	�Т�j!��u�C���"�Ǳ��c���
4�e�����i(�G��e9���RZ4b"��V̋��<�M4}7m�3��簎S�::Jp�G���X�n�ȓ��������.��}m�zI<�]%����զ+)�������,5�=ؘ`^��+e��-*΍��D��(�������񌳦9#	�[Xw3��*V �vl���Ex��'�\�ه�<�U ����v4X��ʏ�~�=���xG-�=�`U��ՍT4���������p��|�%<ߡ8�<x&��_%�V`Db�^z�d%=V�P�<�<�o�����7� ���̸N�O(��J�ڞ�ܝ3���t}������r�"D�;��0,/��e-Ԥ.J�2���� ��Z^��>ThÇ���h7�L��F}���-���!� ���,:~��؜�m����FӴ��B��͜h��96��MJ��@?��7-S����VʎƑfR)W�Κ�-	��1@��V	�uR�8����5trl�$�kzp�-Ֆ�P�[kL�՘X�oԀ�CK)��5���
��6�%O����-&D�<���03��]��ל�/�5�R��#�>�+��sb�3ǌ�-�GԷ�JX-�i# �m�����_Lu.Q=�K�rE�s
��:����Z���]_��}��C���s��-��ܹW�f���wx!&�0s��q�m�����&���hc /[d�fq��]�=���>W/G��UFDFT�b{ ]��ޫ�4!F)`;��z���R���|��$�M���4�H��V���X�0�~[�U/J�y7:�<���(��~����(%w��8�ioU���f���I$��~�Ʋi��������f\��6�����
V�H�(+$�^�5����WJ�f���E���.�)!���fL��3���c�T<1��4��
MbI��>�0�Xr� Α)���+1#��|���v�g�/Mf๡�Lt]*�tT0�E�H�as�,�����)� #�~�[���j��p�(�/�C��F�S���Xrd�Pn��Ð��M�I�ɰZ��	��#�bJ���.~ճ�)ϴY� 2c#��ڸ�yO�ĸ��$\���'ڇ�6���!ᩒ��)Z��i�O��&<bf��$F���3��?8�*���A��;�� Ȏ�ښ��A�:%]WՇ�g��dΫ�*z�	�,����ݞ�XhQvKSS�A��*v��*�j��� i��^g�N�R����B��0��Z@q���<n8-��4�U�*#C:��
6��
i�Kah����=�җ�����R���i�= B{tn�0�Ҝ,*��3W�q���I�ԑ�e$��b�����%��48�ȦF������}
�	q'���mS���
���V���:��}-���@.��,}]���y�t�|aJ�8Y[���^�>Z�Qz#<�[< @a%��
�lR*�{t����ǹ�]�j�=9+ ��,̝k