��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb$�����k�9��1/��%_}�U�������F"�@-��.�L����bCM�%��ƪ���Dn$��9�.�f1k@�B����L�������淒�����V�����1�ęI�1��#�n	ؐ��A�=f3j�G����t빔�mރ)�TT����[j���bj�D�	Fx @���q��������I,׏q�^�x��;
���C�2��y=��L�L�������k�%�JsV*�{i��.��P�~V�n'�57�mMzS����Q�ֆ��&
�b�@��<��o�.l�t����d+F.���-{�	d�d^��9�ڨ�T�o!�&�)���$��)����UZk�t��J��q,�&��pFn����b��Q3E9��T#�q���`εZu������G�!�F��U�Q5����Ӕv{8�O��|`���s$�����*~�B:�ٰZDO^�p���kb��SQk$W�޽j�����l�=�i�rb;�8�"��և=���_U�-\sZO�
��k��93��w/��Ǯ��m��7޻��n�x�a����j��ƣ��-�Eʰ��Ź#��ȬT$;���{��6�S x\�Μnhb']1��r%��]�!U���I�jRI�nAgdG�¹$�k�p�A�U܃��J���^Ȯ��a5e��O;�\ᾳ�J԰S|���WW�I�N�y�I�٨X�[�]��ą��V�m�t%!�sOy��$`W��G*P���[�vQ�P�2!�vb�~�ĥ>4$C��� �s���U�D�TT�Ϫ�y��,P���a�}�1��+_]��%��9 �	"�-�Fn��_b3G��-N�a�_�~r�{V�
�zc�6�~n�< ^4_=��i�Z�\pg�Z�)�I��6��)!�ʪ��1�s���4��q��N
j^�+����00~a�0�q��*IU��0�7tx�Ȏ��U �'R>�7�w<���%#[��(j��z|��Q��C�����6FDz�'�������[A���^�D��QA���Ǖ�kT�Fz�e���y2x��ޝg����c
�	�'AS0Ƒ\W�Z�+2��	�YA��<Lq%׀�zD��%$�h3�;iV�����]���ϕF���6� ���^���Zl��XN4���,�#[l;�7�|C�h�p��Z���s���ǒ�LX��_���?E���N�>vQt7�CY�������"X�H\���|��$z��Tk����b��k"3Q�%O� �TaY����ڵ0jӲ6U�Ci�l�ԫצ��Jz�T5�����qgN&iU�߆?���\�R�T9��K�"�G�P�6ڎ�	�^������x1�
�+F/�,nK�K���T�S߾��*5�j������p V!�k�
s^�/�8Z�t5�jHRG�����.k���~�L����K�o�q�\��c:��׆ba qJ���80�H����'���+���mQ��yr���cn�p�ބF�E�ﾧ`����<Y�ݮ�߇eg�bb��f���@��w����TI��P_���DE\�K;A^�^�v.Vɕz�45���:��;jY^x
��o��%>���:�N
�s���q��g�Tz�����E��
���&�&bjX���zĀ$�ud#��N�:��\�S�}g�s �k��6Hb5�����`���d�iQ$�%�i\w��^�6",������Pց�ϟ��%6/�k�/>�`����:V�{��cv�;�n���\@��l�8�+&"N�?��nLC`$��?�F/�!ھ��2ʏ�&�D������W@f�l2��4���H5��8'���g����SU)�J���{۷$U	�H��5fBd����G��P���ݿ�~X�c�G�:F�tuA�*(2]��{Eg���eJ�x^�<���$b|�Ԕ��vy*`I�RD[e�.OV��D:�Q
iԃ��Xw#u�vl�IZ�;hC����`x/;�%f��[Ȝ�YN������{��	��Z��i���hH����$��P�r��``{f]���=��ް���S/(��%��s@:ba���v��:܄��E����-�_F��d\���q�.;e��6&�f7����W_��-�ה�����#
����X�N���;f$:IS�B����8���}� ��Dsp82�e5#�]��$�ٸT�=�R�j�&�����njC����<2��\��ȩ��
���G��m �q� ��������VcO(��%�������fI��)-�+G(L±��܇� �m'?
� N��*$A���������#��p45��K�g�!����(4p��<�A��Q!���w5����r��|.�$���������:�
C�������_X���S6�4+�V�ۛ�t�?n��Qi_ �}Y���`���1��b���u�X�{�s<3���a��~��u�8���@���+�\f�M��ޥ�_++�k���;� HS-����8���2{c0���9c� ��:�a�dZ"D!�������'Y�`߇�4�.?
�[S=�'���o_1}�B�Q��mY~1�Z1w2�4@���J�b7N$o��lH����tq���m7�w�r�[�{>5ȇ�f�tH%)^+ʯ\?����鶬��th�9��J	6v�G��che�CW�S=��1ž�m1���� �{��v�{#����]}�G��A���2����[�K��U ��|�곬�G���O����O��X�� ?�k*6���Bٜ�%�:��#u���ƞ+��q������=����wr��z}a��da"�"�b�������	Oi��TuH[k詫�c�(|�Y�q���b�a�Ҍ����!$^����V�JG9��qz�q���zf�����r�)%�ײ�Ư�M��8y?4����gv�D}����#uW��鳍�cMʋ�r:3AY6���r�ݸ�#e��6�� T.�ʓD���!��^l�}tƓ�/���x|*�Y�p�{"�R<L�`�p�$����#DxK�o�bMA�����"!Ub��~<�O�Vw�x4iM�ʯ/�����
��D`�!��5�I�w�ۉU�B��>�ĸ��j,i1�s��f� ��D�C�5���.$������iw�fv���[���d�6g����/�z	��b63ӡ��Q��!I��}Gvˤ	�1?��