// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:40 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pvxaeX2ALSzXI9MypKUk2uBzdxOO46ygi0WPEOs73QfYIDrb1431suAq1jgbIrnH
fXPbUyG10AIbOkDOo1Gz+BnOvF/+2PN5PLbqo8GIjX5a9GrjxoOj/WwY7oAJVDzo
Dt2owCcTmmrMcAf6/3eeINixadWzsLF/3xqVFTv23qY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11792)
9pgf0BHGaY+C7c36pga1s6K0v/XG0gTUREd1zUC10sYy3uukgiWM03KO5ZH/MZrb
Vr0jGWSf+yYF4lXDq6o8Ix0c7L3QHXYOxK3zSqlbnvS+RtdAWjESJvXzf7UkDowm
14MrcZaS4yz3Kf/vuXW1mukiXhqosuc0MvC5NW5hi3Kk25x6CdL91W1G/cgjJhZT
wC2aV17KR/7RYr/BhjZUEupUrS9v6LeWy3Qv/0B0eecit9ZGbzq5TG+FwIT6Vz5b
sVfo6WjNJYMAyRN+ApqJFC36DJMkTyYl8WCSuVCPCJ8gt2whOMVsMticeCKQx19d
ZXooPIdf3IrQ+1zvsAz21aXTGvs3f9Awal+KHR0O+cEOd3wZ7WznMxamSTszxpwF
2+JuXRxCaCRtYJwZpXVunj6OBdkpC40mFfRztzCVWUooG9ylI9Q7XD5f0bNE08GW
gs4eEc+iUoOswFlyFrlSp8OoeHjqcWcbIahPH1aX8dSWqoUybUUUtQyLZKJOR5cs
9lTj3cyeqM+kODGL65Z3tIQtZqBZLix+4nNS0rZ5J94cq023RLsydDn9xfQH/CqJ
97DK28XlJXpAVtMuVJx/OLjIJJ/+GEjbj3WjzPELbk+hXu98Khk0+X97Lo9CsPBU
uYtS9eEOczp8XYr3p8GPR9u/0btznw2ziy1Ev+zgv+yR9WOexw9te7kD9h5Fzahi
o/ZR/M8exctxTIywvplofRbONpGy7M2ehdARl97jgPDGpnAiD92DKXhfogRbeRtj
dxG0dhImODXmq7ykinu4KBSMcoN2e/5tuqeSiWG4Zx2KpZWz41gtIUNWRxuaSY/r
nhjjv3Ucy9Butox4L7SVDGBhCUmqpVuuge9QlqJBmAt6Al7hk+rMGbfeayasAjUm
2dY8531CvFixUaZZ7I76VdtOUPbLDxKJRgmG8w4jhopH6iD2ccAvB2oGG73A/dFB
KMuLJ7YB+w/0QlzD9GVFEzQGs8AuUA7fHzaktpU0KotDJCxX5eVSaxd83enGu5Vs
WWFVE8EE3xVwgspgvhaiJKZeS0MEba/GJcaAo78UfE+L1vnBqcpwUV1ps7pzBmMr
O8uy6xPRjRoz4NxnCBxvQyWoy+uUozv0WOz5BPw8CHxwk/89osaNLg/mdYEwQgRJ
LnX8k+s27T4yKdieuI3nKPOka4MzmE4+uYXQceeU73u9AVFwbY01v8+LaXsOoG6h
bbgZTj+Twz/+RGC7COGKt1nzTGLc/IvneoT1a6wlXehAuKX4vI+FeDIObz9L6au9
YmIxAi9o7CKQhTgaTtteKe42058fdSyxUR3HJeClAU301y/KbMPhilEG9DHZa1bQ
F/1YN8ijRADoBy+s8PeixjEKs9hSwMtC5IrNxAQjLTCVeAo7PtL6M+jmJCFIkmB9
LdlWgp2PPLvrwRWpQXF/tnQGP2ybDQgmn/h0IjDaqQrq7Gv9XDUh7gNmizDS/wvt
WX33I9mYLjKV9izCmp/XTQywXTfKd4eduIXnXbLMM03LQ4x6CPKvgZj5z0hhn5An
jwJ2XnuOa8NJdZLShl+MhJJi06fJNHxG5OsP3yx+A0FADREykv4aKlCKFfXEwWH8
DFuftE3A1QmkBlmWbdS6sTiRe1rDd0gngUdKJG+tY38Z0Izo7FuN52D2fgdl8t74
trU9+84wCZK4+jUkNGwt21nvNeoP7jqSjEU9avOfOEfx+xNPTEQT7Aaz7CJPRYqz
CaHyRuhRrkPdi3+++Y11rv/CLkRYtQ2sdhOYH3Cc2gTV7HcXxpgO8bmPbUvtSHzP
y/chWss+b5FfHUPp4OAMSt9yGxF8EBfIJzalLHH0Gbl2XgamdYYjTCzPwNnVgIae
NooUd7TgpWb1XXBI8c2AXRROef4o+0wykbNGFPZQji9casVAXglpLcyEyaXuisvp
DTfMvsG0mhYukn3ZCQu5Th9V6aSPU3khRbUJ/fKDZVLsqzsCdlxEc0KWkZLzr3zP
iFhhApBxCz1+4PRH5s/bTTrF3c+5H4TRhU4ONUJqABCmJu4O7ayyShmnqulKgL0z
XWP9DKY6xlgAKJnsIz5ItmVuiAyNLZ5TSjP6ymJGjO5TWL76lyVnkrtbxaCpyjuW
uwhldiTTSingJ1iBQ0ZCRgNau4WqgUPbOLINYAns/N2iASY3yEgYKeNo5Abv2yLQ
oaqBP2FEWVDEsgS6cemVQWxkjQodgDX3rnvcGejnd6FzxgoMb45qntWz0Vqjk3wK
3CHxsY4VKGqb/kXeMOMqWMo76jCRVrQtQ/6LLLcWNAyXssHPgPsn2ej8KSuFFsvL
C21eHc4frNnc3FsgOK93bg6HmdVt1rew3S8YsmCoHw5ScUDPijzWa+BfzVGrE053
ElSFEf4twUsroRO3lEkKha2RKhryKxmR+gBsFZbdktfy3LwI65nLRDXQbWcliWcR
RGtKBbM4acC6QIAxVu3IOdnNdiN6zz0P07ZoFIVAd1Vbc8umsNDWJw7SLdFIMO80
ObhTptZlySN5n6ENcTrpyyeblr3haf3BZQre3ggrffZlzpNtaekRYbkYqi3CWPQ7
4tCpGGmVdIDJIKyYjNmalydp6ekgVcpEXrrg/h73kW8W4/184uYgVwG+eVri8qNo
frKbwGvSE12ylUsyVZjL0HcfwNhIpObjHUw04Z78M61BQngUfTPR4UDKF5hoCKKk
8FWh80vHl14K1AKxJzI3JnX8JEU3dgZmnNtp3UT8/JRzYagk/iQaaYbiB0jrC7hS
HcdYEl6SBaGsclRK5bABFoClRrR26CkIxQFAsz8BKT8mGMDCA2VHfnvOvNssT+Gw
aqBwP3A+hS7J4a7x2rYAG2dnkCv92ZhinN5uhzcMFcepVo5yZICqtDJG2H3ldU6M
AZw5E2N0Hu2+QOHOHfS2U3ATwE7qd6sJRhGR+W1vKU98GYHamznbTTyD9Z221hPc
RWpSc+yI3BlwVnsiDAhYPU/9VTB09MWLRJsiJsWdph8j+9r02OmYI9xzz3En+pJQ
r+9J6fhAKFhpEY1coGlXWzRUEmfqX7K/fOFVZ0hGf+Rrf0VJ9xBRl0gCegggKpf5
+aLaKkPPwXGkynRzhsQXCb0VKg2N5RK4Vi6m7hgKzHF8AAGNwZdn2YYmfh6ex0Ux
PiGLQEgbyqzgVVidVJPdDFRX06U3+W0ljgtN5gtKQEXEQ7SmsCgtCPaB6Jy7I/R6
+zZRu6V6uyqY6SxUNG7rCAp044Iy2C0cJgZEw6eFeIlgOk2dLYg5LEUO3gb4jk5O
tqNfx06ywphIJDT1CG4RKgSHGkcfgEEqgSqCJUUBwL1ue0UkAeqPorEc/s+W4FVH
5wgiHvrTKfAF71JWz1jk7mWl57dP3bznUu8uibA/fHGsJDCRMgjGYf/x5FzU61El
PWKqlquQ+Pckd9F6Xx1co2qYQGpstJaod+Bnn+bxJUQnia5kI2H4CkxP5Txqp+Nz
VYWWwqGD5UzskAYTnq/sFNO5FibHudZF74pKNoDN/kYRU786Xnrlc22dOCjgBtwG
yCNDxvhKdJettDp181ybbyZL3wS4OdI+0ZCK6jd+pMA/GaxOnCpZsLMSIvGTU53O
0/jtBPYWOyxdKPC1Trr65Q7oFtp0D3dg8SYWKJ11LBKoC/W3fEYqD7crYkhmCEIV
QAhYPf7zcyoBzJm1iP9ncTP5z+dSqc9yXaT3X6dmWgmFsBQo6ISFaI/r9/+NmhyJ
0vYeSif6EzqrquUb20qLRHXdCnxd4euhxdqbEJ0dmEQYI+tobyOBIKiyqhReLymn
PeOt34HUspXRbFiwSdXN3qhSdNlLYwN9eK4zyKV3mp7afE0rlxqyzDT6WdbDUQGg
l8MyS32VXPhU5nhYLIaomsmIn+sCfSH9be5vyhyf17k+5TfW7syXLAKaARGOQJ4q
S2vIkO1RyZKY3FcCvEBN4k6/M3mMnX5c7eHXC8Ii9YiVbzeIW5G+P7hg7rsGW2E/
CLc96wSzxXDj54xdSd80DDxwALNhms+nMr7QD579+JuuScFx+7yFpP8I9sLkeEUu
PMTpz9HhcZPnBBFqKrShjMFx7n9xIYkAVyhfXAqzrJQIoMUTlue27AbBh9C+Uzm0
m+afI/h1ZAO8N18OQHarPFyKZWXtMhOcWd8rFeKIlN+UGXFEgSbMMBaycqrSgq86
HVYaGgW4d80wH1IH97XyNpgkUHLnIqIHNkd3YBagi8xTjqh9sZ8czliQBKIrnm7W
jUQnfdB0+A82luZdaaUFNCXb7VbESQi4cSL5GG6qbZB2F4ASelyEep/5w0zFcr1Z
Nfky6nCsVPqf4ZYSVk8HSTwhuJshVDP7nc5lzAfyncZwj/p1dHwj87RvrouSxXeC
+8Zh9RymnubOqkEHRLB8e2EjNRQsq8QNh4Kt0Sy7Zx0MHd/gIBXf4aVSUsQ7PVBW
xxwGFNvarMRBIpG5nA1QgaaFmhJN01EQEI5JUyB/LoxHg2E98U4/CYLDf1A7pZqA
k0STYCCPgrOahxkWhLXyNwrcTl6R2CZtDvxfDUv/lqDgzkv09vzF7qKWOKx9qH8a
JIrVVVaLvgK3rU3vxHkFJLDMuMxdk3jh5b+rtgFfTGi1FNvmEYvd0eatNgrv7EHN
MvBI93JcfBGxldBLJcSVzO7NrlkSY02ywn5xaQTRMlGlZGkWJPMdf1YBb79de2Qq
XuDXeqfvvMWgYcc61cgNCypJlCjeKPlhV8esFqgrznEWKn09o3fIDIapkRVkFLD1
oQxJ4AzEFwo+EWGyQg6bmCpSU6RoE21hioDSRY3+Tq2FqMRZ7vz2zsNeVDS5OuuR
mEfcH7mrUXuQ3y2OcpzZE4xXMquDpYo5lHhdUCVX272/iqH5YIbH2cpokWbWPFsE
lYPqts7uiwx4+yBny13vt8I/gzlBs1ESwgeiTbjUEfyEz195sWUR373D1/OWn18f
GJzJJKX7AJfvFKEsdN286zHJgq/r0yRMtNg9L/vJQ6GXsaKL6dLZr0FYCiVZYbWt
O/CXRpBSbsEYygxlnskwdCqFpsmoFue2xuLHp2o9xx8Csm4XjumccnyZblt2Q7JB
N/ud61ScOHyCrt+XwtNELyQc2Jz6YJpGF3GeTlF93PwJG3LIAZmW+AxE2PbMYSlh
TYaE89pfEBWn8EkvcebXA2u8QU/QlfqGiIrND5xW8VX1zj7kfJlk7frCGRMUd/NJ
CHRP0SvEGg7h1PQPcc57jqtLTJJKM3aN/rv1EFYWARcslc/qJmC5DLaB/fGr05SO
sOmpBIPZtZXJyXrffUgYn8WQt18D3WAz5tLAY0qpBss2sCFOmIplcpeTGx/Whgsh
SBgnzi6TQQrALAKZzewjtollKZ7WxRBHW+9ZuJBSj7FywnEZ60/TAwZI6GppDIq6
iORLfYSJlpmtIs16P2eTDmuMojwdGhTALkrGz/ork7rNk/CoIrtWNOm/ZKJP+QO8
JIVe3yjShSKYXKAo1IRPPmNIfcUnvkJv4VMGitZguVgYRymgURdUq4yTdAXWp1Y/
8pz5K9lQ6enUKO3zMDmBsjzlTbbZJe4Iu/z8e4TBFBwIaAC/hJ+6kM7xp3ZOOPBU
0Kmr2grZAjNq7Yt4Im2L9iOLq+ZbOwcSFSI/ceZ4bxZdlhKHLlSZTYLGnmZ0nMU6
0KwGf8ok94hKEhNKE6N+WZ0LkJxP2D2YQsPy/0RjWvD1rjLYb0wc7geX2r7mFOhl
XVfjRHKsDOgtL1jdtUDfjslej2ylbLbvarXdjwUdxdHgJe12xiHZVv8OnlDBtOEs
06zStu1NnT1pUUmq1II6Lg6K9tYlKTp3MAo3XxXyZ9/Kg+1jfDYeDdIJbhgPNUil
tck5JZd9mkfHN+GAChqInLh5uWwt4Gcuwz46KYGPJCZW2wMnL4AY7m/EjPcKTf/e
SMqmTqOizMZUQ6AJaHtWzf+2Q85FONAvmejBAVW2leiOSxHQFBLGE62JjnT9VFID
MBeKSBJ0jOdbm7WvdB2B1XFwDWX21oNxWsQc2aKIlFINQfresD8c5eDtNMsTNv2q
Q/IBDpUeGSewwEs60L12ZR2HPGLeDaEiUcJOQtCp373ROktxNYKHNow3aMlKf+js
Zoss83YVh+VhVTOwudfNqY2NwmItwMEE+HHhLlNEnCZGuHFKUW+YHVE+xVlUjVK3
dmKpvBMw1HVt+7Knw+6+k+jwb6UJXbMiM0BzvEWJAdgvIYbtp0xyEloGli/x6T4G
nqU8I/JE46awDDA34OdtkL+q2DD1RmYZvlegnjTZtILdxqPtuvBDDyPO52iYaQKK
1F6DW3FUI7yD7JNaXSNP4Qit57JRv0fZ2crQRuUY27Efb005dilAi9EQjJNy+KMm
K05Vzwtkmb9pizYw36DWefEcwSPwGCbZ3UWJRqU1UvwAHIluB5x708lNLkEXoBR5
n8vsBNB3zBi17SDpeat7l99hDlL2KxH9KR/3hDl0Rqk5sQdDIcZAcD1WTnjObtny
qRPdURtMH68Zydk/5gdPnmDP+xKT2xtQT9hBMJGBmOJoV7N1tIAWkFfVF0WIKWUu
vu4oAS53mBFlGwlteTLmYQSljyUGgEF4m79Lm1ywf1fD+/zlyVDEPZgyNERbny9d
BXlUUOuMFkWnqmnuZ1eb7ukFHmH09SMgISAK9B8QhB7v8anyZHeT2v+7dfjTDZYB
YtFxpaKoIOK6g1yL0DokjKEgrXE31dr+k4W6npfj0C38rr1F9JsPOcXZ2k1thl2H
JCRbovipbgdfco0xiN+ZbeHAWL5epIPUHgemq/kBuuf5P2HbySjFHYQgfYR1sZLE
EN24ZOH/yQ1Q50ZbjWXDT0Wr3tYx5Qe7KKK0FKRj3POKEpYh5yvOknLSPNX2dBlO
XHxc2LbbaLLU72SFQf99ikmZlP4SSBGV81Lc0trGXRBLb8ZK5Fhz4dn8FRX7qTZn
eccEIYNEzjJf156NaBXNcYcez11oD9PqqwlYcv39vWYXZB7m6Yd3pJdnzqn5J7Wd
JNx+AxdUtUNY9Et8I6C+QcC9DkX5WBJA3LYPfUOv0aYN08ng917pAH/su4peuZgC
zqIzmZeGaZoApclCUAKNcsr5Q6OVgqW9iJ8gwLdHrkRiajlmvOm5oQIHa7Pe7CFp
hQMpj0hyLXVOOV8G+hdnUiVpysNrFrxcV5CrhoziPAX+Jm4REFGroCpVuB3wLP9y
+aM0bNh/rC0HrrylkIIkDs5R73GmNuihHzzHBCcGSP9YStmiE+Nwx+sac76SQQNb
fGgkFBbRVTHG4aE42ZfgLd1USscAXXCTR3x1d5RFseRmDizTF/dCzk+KJgu5JrNO
gJXAJV8RDwe7irn74TiNiLzk67PGQYh549ozMlZUBPI6igLXVrofiVjI+Sln8UHc
PVgD78uE/V7DYr+pVVH/KEIMtvQxcVOQTduTPes1RmCR/MM3FYq7EiA84COdmUr2
9y4B9lG09osmlSZXDlIVgMHwtaBW2hLwAzW9UkrjhSpTS8pQX9pyuyRtKt0c1yGd
CkJTmq4cj8dbnPXbkI7HqhODnUKUHYNgt6GBEQcFZT7vPNhRcMOk4PHuq6IsRLpO
32ukwqj1eKrN8WznvS8vJtoRxQfRxWfc6hf81LN+6FevtxYbLAhWmSN9YPN5iPEX
ML+qh7+2eBRfgD5mvNo065RnYb5/mZv3FhmAHDbicYeRP03YRDOMQgRU8tLF0Hsl
WeGnTUS8U6XdhJN2sAT210bhVQiSwgYsYglHGnQ5OlqyG0ZQrGfu10cuj2zq3Fdf
jj0Q3F7aCrqtdJ+xJyRFa8DO/LD1gaqFjj8WBexnHrk2+LUC1MMy+XTJqzy1biI0
ECWhqn0raJEv5LRdTw/RaUO8NVnJB//oamZmBhoJ+VMSEA/oUkAH0UXKlCiRZEWO
qpox4i4IwaczYDiV20aWSo/Uxk9Nks2DnLFmg59kwWuIp4HAR0rUc9E53sDyZ2LA
fyCNrkW7rVRFYgHuySqFjr1uixwqqbs208+6c7TM63Xu8C+CHr0I237xYoiBX8TG
EX8/zpSQVnSEEJzT9wZedSo+L1nVLi4DLnfXVP3ZGX805Wi2P+CFmws3WrEFMqnm
3mSB2/g5BFxX7IEApGyyhdbUHdswCoKcOfwvIlNVeCpWAiJrkf7S5+PInLn9Jaw8
P5AG+Oz6fJiFa2EP0dY07twxzPJynPdxPBBpFiw09qRAUvE/hPuaGRMVRJlaMX4H
HlXdwE8Pwd2VFs4DpxHtJ3XJlWhhOIbH9q0KQaFUCJQEq5MVcpNDDAWIMJhiRBxk
8enbJBv/AvLpOIfzzZr4xNyH/+3s3GYDmPflGXwZkvONJNPOvx19LV0VwuQLzVVY
nklTgsuNi2q9MSBNFsHk94YP3hGlosZivfBahAIxyJ24F1PWlmYQzr6ndgyzN9hp
w0AZPtPH00rdQ2JX6oCMAux1VQRxf7KKsDq5RAQl8YFifnxsmO3JuufP5xiEgJ8J
n1rnafTT/UBMgFPSetMtSv/TnnEwg4tlNs2Xpda+7lwjdL3/fuKugBekH26VT0ap
BO6qdcpyrpDCsixdG2PtA2gK4FC3k+t/MsZHTO6i0wYkRJZqGaPaMfDjU+haDocy
SSu3eWbPlfwbj/RU+TBXsIJJh1i9Tm0nHylWFKSXsyvsJ4Bx1Qw0SOZZM4UNFyep
HD7v3D0F/wd8J6IEY72YURYy1yR4CH8zIpWG77erBvMo/MVdY0dPQIa3+dfy30CK
NUKOOGSWq/0ame0090bIzMnRdpc0pBzjSDvTXA09ebq839ow7p9MwE4YfWmV6jVX
z9rUIAWoaJfgWTfGaxpng7J5wBVpqrTciUTL/P4zzxpNAsyKsT1DID63BH0hIrcx
BeocrtJC2kOJrucRBg6vy2msp8C00RNu33XiWXZiVsYOt7KEvty9g3gis4oV1rDj
RLk2zk025m5JIbLkQvGBJ/nIeBZZDjUEwgE1DEXEezdtsPuS66pxGoDyoZj/UZxv
4lUFmUE+R3LpKbKz87WIT4TGvHq6gRnjKCqIpGM+b4cELVD5YE+zXDRpwXGVnaKC
cccigX2/kwiZ7sx/saHwAx01fh9ltcT5wq7HKxuBzurTttmYZC6e3Azrh8i732Tj
GKPEQR4u6Cx2E86Ry9477WwNNM+Yir9hrf9FFG/qCsKrLtVjWqDfxC0LjCnqGb6g
JR8pTjhMu0QZHYxuUXwtE7jc0vamImR0GKthSLcFe1NibvGFkH4DJRTl1cLO+QhJ
KNySCafVAwdtkKXbCeiB7i8yi2YnME63FK0+OsGMC8kX3peLfstIGnfZIBNWAkWE
oUxqeQPpRXKWUH98gtfkjXaU8VOjKbR6lVEEUiwTagGXBAtNAOUtsurA0pZY6XQv
qjtNY5UXeYL51BxFZZqEPci5X8TeSxG1ge1aeEtEPHd4aCcYfZAexOW7BYG4R/a6
kZ6tnkb/IbPgBi1K4ZTq0Eh2SNHXzBXw0ZXilGesD0zVo0oZ6TwUZaXEcKoNXS9B
xkoeAfx+c5PpeV/KksthENwOqd/j7JwQBK7Z6XCsTKCIv82ltQYQMyK/hEoldv5E
qbKV5pcqhPg4+VWPQHj+WnDyDzKwJmE1fo0PkUqsm9ojFgrBfjEcDgSxmD2NAfCo
VHO873X5zpTvYaFAKfIKpIplEe+JtKkMQdDbo3iCFGi6kc7QK9yIpoGi82BLBGCz
rhOz0fO1jPiVi+CDbVxEMNbGPyRGWvHHJUQdrcPWAbz0Jl0pdt2eBkaDmUIhCYyd
vaurP36eyhhR1EC+ZksiqxrEJg0A5zAymJ5D8Zp8cKCTxljQHjWXsKLqrJk0YS5n
scqsAJtnqc6nib8DEbeJxKJOSgZA+sy4VFg6flpQP66C83EUOqmSEkMZXUJUYGjh
G8Tl5bqmlgi/iO5PzmIQmANyCtur9OAi/mX1Aa/dnn/MI21t021BbA1PqL7xtUsn
LMYYhZtdHdWByjNyHnkQbxfkI/8YU95RRSq+arGrFICjyQv8kQz4PSqSffurnopv
u1M6+TtMIjadLTnvC+9trYd+qkAeynL8MOvt45+gDyWFLNQHv6gVMKxkJEW8Fu0W
d+TxUCT+GKcnxoJW/D4HC1zEqWFaHL7I7t0APUF1BDgAX9klePT85sxFZRRmSum8
dQWdPGXe7xybWKIvBQL1dzeAV/t5aksj8q5RBYUxNkYTD9+RN6fm0thd5cps4gbl
DTOhX83F2C3lbUul7gwPSLFNvnTkZkmcNurGBFmQAfa253vccwmWjbjrBE9SRxUj
6LTFPX9hQkvh9L3gUh9I+bKq46G0wqbjz8Gg9XFN4+iv6uTIGb4BHo3vynmQEH4i
yuUSScKf188Fav0j8ZZ9IAJrNVIuAL4o7yEpGCvv3pjXBIPYHMuwW5p/+zj9Y+nT
0DBkzD/PlFSk/4ly35ZI93+q4KZHuYYa6rQo4t3nyPqy2JprY16lq190olVaeP0n
nZv1+mKuHezciQfSbEdzXbJp5vojPQk3XNYoP5KIS/yxvON1AYD2/IR+KeKWZgh6
97+KDmBm3Wr1dnKOny3YPstnd+N60ooyxMkn4moi2FYGbGqvXndot3Q1mvCfQASd
xND1tF/z4lpoJxuhCKSLeO+CIjSo0npUStR0rBfDu/T1sTCWtZg4v7moOWe6SdMt
EZKVE6y6jKthFQ3RqkD9ipuGExe64ONbZV25ZtJW/lQEGyEmERr6av7VLOwZqFzd
euHlzknKWM2csqr/BZSMxKA2Xkz1JtqEYd8iMc3jekFOGchiV3CYmRtsi9vglK31
LOJbQYW91fT6rOMBXcpPezgfoiw/ky3Eyqlj1CoxnXMnaULD6QIGnryHeI9eHhlK
KpNntRTuvtZ/p4DHZYAuJ5BOYPltWejhh5g04Mb6XX6v+YAvSSKwRJbdT5FlgsPv
xlcO17kCz2SE5ZVenDpfKwFeMJ6kp0CSVEW6UjGS3kFY6QPkjenlw7cOk+Gi5GYZ
I0rQfRcaECCxjYqEPSq90ARp1cnzbOnddHMnOOph7cbS3eVGNzdoLUHmB73dhUq5
Zg7bXSfK3sQAYjNQfj8S3fpd6SaTF7qwRf+VRvNT8dRp7dl+QkatYpmX2wgC/5Rk
WNNqzs2Ngf/601rnl4Rj5ikpvqfni64wqrvpAH3P2Z+d7CafA4B07njF2dB3/FGn
yZGJSgHsQuMlkGZtlQtkLyc5jL+vhWBXdkBy34JsFlxtQq+449S/fhwS4u22lrHs
fCbmF3sKV8msHUxIABTKcHNtQ74gs9lb+kucDASkBDseUDFwEJ4IwvObS/D5e4Kn
dOn2CA65YEmKjKROcTHMs0UILDMRrBHsmIgPgy2eIFyEyWTHRneYWf7VA8pvDRvu
uOTh0DPMF+xxBsnq6no1rWS1gWUMuoiJTJAUyPmL9sfymck9yVI6r7e5TiPxEqiP
0PvT5tIfPwrlOePJ966f6aH7tee9CYOakTC5LMdwFM5hffZeAf4YAC2Ede2KBcd5
4KPYG0tBdEVMr/1wyW3YXK2k21GG23sCkrbTwPAHWDXwPnZhErHbCLuieYoPu+Z2
phY17p9+/+C9Ugb0q7v9uYU4x7/9rSYbTA4nxe02bNhuiQDTSWsPA2RRtk/H+0dn
UkSNcfhDz1ULgop1wCaQ1vi5valmoSzTjEidWSS/7jMEavcfw7WvlOENRoCjdgwO
DpMXWy3xUalPqdTcBIAAxVeKnoqnNYwzmtlWyhkSGsVqb747JW1Rs2F0+krSgbVf
EM/7jlg3Ev8fEjfNJ0F8o2DskhXvdtPP+EXXDsSLOA2KTY49XIN9LCmVMuj9Urpy
hK5jDu/NLcYyQlqalhcTuHv+8BeUF68YFlLiKlBN7WwDIs5otX5P50Gu9U09ftoW
pCn7Exvz4PP1dkpiSnFxh1KUenEMkt0Xh09wneu2jj6AYUzZTgSnuaPPGJMMizP3
Ah7lDcjVlGDWE2z6q+XCmg9WO2whe3xKAhmeIiUge5gaj+3fJnsRQusPvIMLG5oE
XGP0JIGnx2RnTFARYE40bsBoCm1mOQnQ285QXyl0sUgSO1LasMLbpdsEVjN3VmrC
Gk82fqY03C3bm4431R8syry5GgeBJiU4w3xb4LVSColK+MT5EwKiutMS80hg3ck4
a+psswh6Ov/SpnU8hMeCTzhUauNW8HA0yDuMlyoLyk5EQI+607qkz1GjOZtxEopV
k05Bg0zDGiarcMdmnvzqK4EWKrlKMlskCDwKiC+NbgyQZIwmSkSkiJo1MKRaU2lW
a9XYTDsKjc5OLEJs7paWgxUAgGxcIR2h+4tmgHno3IA+iEtr5mo1SgGhnMNhraKZ
pGEu4zgHAj0KzqtPjRRjWTgPCLBzU35fDfCzg+BI3ZyNkmeA0Q+YzjGPtlRuIpDV
XFwollmhWQV4HOFyIE29rvmPTym4MxnHTgFvvcP2CmCArlEBo20InK3qn+LlT0TY
7NlTDuppos7PaF76O21WijVHqO/VXR9LX6aaOUTDnESmrEex+3XZh165Nx9fmPU1
S66ngMYf3EccIa3LK7d7kaVMyyZtU7gmY5uFxtFtjAa/FVr72scib9666nsmDM9w
KYG0Vt+D1TQtXvv2qjr4rBEDKf0ykeEzK9OoMwZlEtWBgTxZn7JYtklVO+i+IhEV
H33vdgwjuXHc3d5fspD+X3H9R390kXEA1TT/hnJ/KLeYY1dN2AB7ELwltpSad2R+
BEaDAl6kG2Jl8LudvYm3RKYnjuYzw3mDEh32wQWvZk+OxGa1utguWkrln+pFu24h
ZeaK1CJFzjOTZNYMpfVu5cuxkyFA9MF030/NTRw11zMp8Id18b+XWo8fVv1KXJzQ
z+HzTVZURm36KT2Fe17s1aR7AsIajB+mXl+ZCRwPCSOoCUaA+hS1LCC/3hXSnp4h
8KMFwLvZoeP/X8KNJt/m4ezD74bo5YvI0TazVYycHAPWpGL1kaplkqFZF4ZDL/gO
GblgCInFgDAnR7V/onVSiOUcfhAL38Ync/rcjnLQSZ4ZEpYnSo0SObSU5OvcdrEN
qEkkmTpJpTvU04yGbWuTDQvATVwIIGNwsVhwrbpTFYk/uWvLx1ZTrtOhCkGOEjuo
Vdt8VSwwjNl3OoKd8p09isZIAi3+cy8FsARb/yR9unTfTpXQa7UQvLk68EB2Btm3
M79VZiQrUijeVQyN/2EfkW0D62W7y9M+TnUPZ8Fz72PMwewTQFRKXzzH2Vf8Moq2
h4WKEkHivPj77dIyCS+fI9yHG/cg9645wpcWSTAyn2yabD8qJ1nD1uqoC0C9r5cV
EEsRg+TiI9Ob6IThlHgAqxEoPTWjAZwiWxPf1xjV2XQyC3wExJLp5uhH2+/4m3aD
7iGZiLZJwKX7/egx00dD4CSTU7en4cZ4Gwp6ZhJidw8HjpSivL73ty9p9XQLHdmL
pjzis5QdjxkzpFV0aaZBsrniMja149rRfNAybboc3aiJs0ar0GXS6X8MjFao6oWQ
YvCzPyT8cqu4gvC2hOB2W2u9aTV2tYTxxIC1fnZa4bI9V9QNTUn8bUa6BTfMu2GG
jpvQ6Dcp/98eAK258BItH7ItSdOSsGlyc9LoY0HcXqd3xHQuW7AotHUBTvh4tS1c
TvdChlyRJgX9xGaAgv1Cw8qK75yho7bjmPMbj6aXyq17y3pSD6ceu/2KdBOURIji
kRvVBTkBIh/wiY7U93dJNrcJYPS6RwrFOF4sHghUYe0dHs+P7VgM+w8UiKHku4oP
AOj7LngJKP3ZZpffFPNVBOQ+GEMwIFXYsJntyFZx0MHSWaTOjCL2bGlaQjHZBzLo
wDVoAaABiQX1quiRauxKmsYhLwdV7W7hvzSXwPlJZgvdsiJJDqfjsLMvSgcIAyWY
pcwYgteUrS8cBNk1EvA1/soTzNKEbYvt4elYtX5CO1ck88AqlMQ+Ebu7Avbs3eQr
u7M+yNqfluwy1JrVCFL8FsparDlGZBrePrg9Wwa0T0WikTNqGm/58grIYIHyjMvr
OXh2mPE3UWLE9kuGj8BcsKAnKjtbuVfCBETYboGdMMR+NZWZzqnN9blx1BdEOjL9
lx80dD77bBSnF18wmw2bn1irQr0Vz6gJ36nTk+N99BPIdw50CWViMl7M28amNkyc
TgX/NvC1ikSq4vIxVZZvVzGv9xuY3GdaOQclGuvghZ5EyH02uw6KsbMHKUIHgV6n
FEn9SuT/UBXuxrrAzlkNFUeRre2LOZOJzcFYvl8xwgLgzcIVPGlHDQodBNLtPBvc
T5lnhBHuaQLhgXmTlHK0q8KUyFDf7K7rCRXa2QxqcxTnuRvwi+cC6VlAmywl/w58
W2IhjiQITIlX82VMZTynN2NNJeWyt6YvMxKxbjaCRluiA54zi7iT2gK7Y7BEYqvU
tqv0QMTa5TVo8nUDlVknJdSyDh4si39sTytxw+7mcMJtbu8iowFmdMH5N/YdmakN
3ak4GdQcNRcCk/v8+b61zb6IPBZi9fZSqHCiAaJZljIn3wDIEaTFJs1FOyTOu0lw
WvVuzqEUe+TAz4FZCbFCih7YS0/67oNufpHOGYgcdE9cLzsupBlYyINQir5YB4gB
kVc57Z5/7YFxQ+pYoBQgV+7zj/5nnRBegkBT07LgwmhG0g9hwi2JKjdE38qYwsCh
wgM8iIQvoUTWPht8IoZc8eYgAuPxtsEwCQCtgq2vHZFmFxv2gV+XCiNOelyHl0hA
zKDcxWTvsfQ1QmICgWDL+KQZmftKAZq6klKTf+5UVtcfsvLWsNn4qbR+N7LrLafo
YCyK+IhtA8JtsEGnoqZOmngXpbY8fVAtw5KXSDu7zj5B0D9qFO2XF0hOD8TtUU4k
6jA5FTaKm/Pq+4yi0Oc5DmgtvP2vFjD1Dfnp+089lbJ7nbvX/11BEjRXb5Cucv3k
LYN2zzVjgcLmgd7q0OWgm9Xu5WMoGAxQu6uI3l6i+egxHbGCWXUgjrdux8CFQLHH
p+EvIwu9F0PQpH+1JPFPQt464iOXUrTQIu1n112RyQ4AAxb6eUm0d1Ju+qzcoDtf
dS0fvPrffETi1//tTenJykBRHM1WJExBwQWIhLdDXESAR4xeSBiCRwAVt9bljM1/
mar3q+Ihsypj4FLK0tYOr8Fibw+czzIOjg+6kpE8hMMAlHFqbxToyr5AF1YCd6+s
CPjVsH2cxDHgPyfd52zxFIXV8MIbwvLw6RaKf2qtoZzR+/Wbk4/TYeh+g5n/o/Ux
H+XSdYY8QQWHH4X9D4ghGxPm8YCNeKUY2YJ03J/odmKgzdHmKpvbXwSDZvuWOYcO
az3ewOZsDCD5/XtRkILYJ1SVe+K/nrMlHHYu9RTXrwyy2aMZe1Z/IM+XgVdNUwTt
TMoEE3Gc8UvNS0AiRGfygyYzTxaOev2UWTDch9807776uEPGO98aJtOiNDAQyxeQ
tyqNgqc2SI8EfWAcU6ZSxplhMtalqKxtv+8w5m5aJwagS2eZF9jqbCrY5L7jbpH/
jksLjxBEYFcKP9PttMjZmqG6PeKoGOJw/+y51czbbR7XiY+iO8CGCrSkWaT1rcKH
CFAPLuBXI1LBRTGoHjnH0agy8iWgnHqtvFmsmAOfWl6I1QD6bLhKPeZAvTPb4LHb
iDbWmVPgb1rqcLECU441W0yrYX/QD1ZWYh3xIjUHfPJaqTmKD8liMeX8UOmQ4QH5
Fwh3Gi0Y3iiVmt0BzmYkfeOAAA6S6C60yu7x/ItByENrMngHeRbu4No2Vnm94w+5
JoQmK0nvOe81hP6rnH4CiMNGjVOx1UEHAqQ462XMxDY=
`pragma protect end_protected
