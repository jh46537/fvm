��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{�CZ[R���T��|�&�|WR�e�-UE�)�j0o1�`��di�ȋS�~���N�k��:l�t}�m�!�7�A�����fn���pΕ��&�����>����Q�e!�-vՈ >xx����[���pH�j���o1��C�̀/�_NHQ��ǡo��{1�^i��S�4���*�?Uv(����?7X�Q�Y�f0��F�($n��g�a�RV�';4˒�UK���:�֡���^N�;-a(G#�LXK94@�l�Z�i_Al2� �9:�R��lӠ�Lm`6S��Z������mn,�t/R��[<�L >P�Ӱ�z,��-_�����qa�Z�x>5�!�������h«�y%�f{��. �PWx�h�yz>31��ec�d!-�h�lfZ�KԸ>�!Jv��s���N&�i����-���H�M���nw��B��X
�yR�=��¶���T�\(QgU���a�ߦ����s�i8�L/�'�O��拓��Yq� �c������dı���d=Q ��c(~IJ����R�9�8+:�Y���(lW_��׊�76�	��w*c �	�\�����Vc��_Pw8&s�8^�x�c��f��%����S�U_�^."�ū��E}M�d��Q����j<�h�@u� gZ�g����
)�ܞ�ך@���7L�PFn��=��� �8�����I����T$OPnEKF�a���N��1i[��G@C�^�o��q�W}ܝe�Y����|�����-���_��G��h�K����}`��O�4����1�#"�z�)9�{�} �cm_��D=���9���H�_Uʺ�}5;R��7%�K:zDG*�ޡH��F)�7%iS�Hx�ƻ�a���H�0z��5Jw~^�8y�H=SG��&L�y]�a��ez� B�{����9�>񨚤g��Z�z�1Ht��z���yU�j��f`��bUP	v��²���rhݼsM �v�Q;�cKNSe6��E,��ڎ肣.A
�)��A�?�E�jy��T�z�r˟~�dѽ[�g���=1��3��W�x����D�XC� Sɮ�7?
�u�'�U�BX8bS��e�.�����σ�zl���:tw�c1��B1�����<��+r��\�y*�/��xX��A|����_�K��Rt��e���!0fz�EK�N���.[�)���f_�|��aJ:;�G=N𫍊�Y;yi��s�R�̬t.
�ޝ
ɡBo6��wk����ۥ�5[+��yn�E����c�\�	��E�w�������/(�<��O�U����ʻ��J{s�v�w��V=g������bq�:\��{���8�`���� "���z�{���q6������\�Rr�nņ-�}ﺖN�T�	�s?;�,�{m2������E9���+k`[Ne�{L�W ��¹��Ik ��� �e��j�\����~#�jC�/�*�9����[�ws�dz��Py0/��M����i��U�+��K��F
EƬ�L�&����o�V�5��r��d(��Ѷ��Trl���o��7���ˢ�?W��=�i�r,n�&Y6��Y��F/�P�o}��X�e)�r�8�G'�i=�K�ې?��ƍ_U�$���q~w�ꯨ��c�!&��7��� g�ކmX�*��*e��u��2d��n`9�-�&��U̾D�I��үwʴb&[�C���sI�9�Eզ�8��`]0���u��������ܣ���	�	�3F�n�|�x�4�#G�PϞ��;;X�b{��e�̝ÃPf�|tK��0ަ�X���W�퉌�yY8X��W������<j��e��M9��rQ�6��mO����%���A܏�h�y��B�*vYeB�(�F)�֔+���љ3U��j���xD/�q;��J~6����E�N84��4:qߺr��=�N�D�ZJU�w]���|��|�q>��@˄�0td/+�m���e���r�_�7�����{���Y�?��l߆��A�F|������4�����#w7��j�EL�Iu��#G0�bO�k̜��F_�7B�.d{��z����d�_!x+m�����]<�q����r� �����t8��_��Y��[���(/�h���R��*A�q�@�k�衈&���|9��/��<�-ў�v��s�҇�,��|ko*� p{u��� �z@�f���F�-	sH�V�f+�� ��L�kwUhx{1��#�_v��*|�Y�/K�Ʃ�' K[+�)�v�dbbWi�,=��ٮ��x���?aA�'?���\Q<:R���1#ƞưG����_W�1-VC�_��Q�bE���U�&!x?�ݧ-K`t,�?���
�/x�mP��t%<�>6��FeͣՋ�#�6�%�<�b$'��}���x^\-�l��Ŭ��6�*TIo(&�������q�E��<��*�}�<q�������x#�t�	f�P<�lE��U��)M(��uV����՝Je+(R��f�P�T�vv���rz����\B J+������8������t�K��N�	�Q�?��/���}s1����z=i�wN,�V�W��0b��"�[����e���mx�;g@�/r�gg(J8�gA�������>�<�d�l@�~��(U