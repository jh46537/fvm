��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}�����°ȣVhX��M�=?o���.@C|�Z�1��i��g��-�5S*#ƪv��8}�*l�>�	�D��xL�kkg5�K8�*�$����)8��(d�Y��j���	�}�d,뭭�.��0�q�����b演��{���Ѓ˧|:^�h.��pz�+5��$>s�P%�kf�f�f�g�@N��dU���HO�ʫA�:T�(cF���3�D{��k̈��S�~��6LΠo�->�u(2��ivW�b�q�*���,3�����y5��A��5�����Ǒ��$�߾�q8?�j��X�B�当Ɏ=.�a���� ��PU6�UyP�����Ɩ�(2 �F7*J#Ea<5F��� !ƷI�p��UG=��m�\)RF�Ņ֭z��f����H��:"�~_���;<��ѯ��y^���q��<u(?� ���9���\aB\m�#2������3�m�������e��P� ����k�b
i�����gL,�l�ސ���	ۀ�4d�+�ZKpV���S�dg�6T�r��})�3�ӑ���<�>�7Ӵ �I�}{������՞�����?6�) 4�
��=���(yڎ`4�0��URH�}�� ��*5�b�>���/M�	c�O@č5Y�]��W��r�ޤ��͑y3�(Qb�x�`Q!s1����ɽ��`�N�3������ln�r�������v;{ �����
toڶ�^��t���O��">�g����ݛ�lڦm�Jv7�k�_mx�{���c\�5o�)�Ȕ�fٽϮ�B�H7�i�����*��, ��̖�������P�0���Zx��S�UE�1�\�v��;�&���}��~=��UHBX�>&@�ǳ����^�ޘ���B6R(��	�Hj���]�&���b�1��<{�R� 8���^����b ��=�󙠺�m�эs��$�==�D�΋<��%C���jcsw�s��ٓ>w:�uF����C�F<8���h�X��,x{��9��P�"F*��H%A���A�����Rn\o�%Y8W�&se���BR4F��s��*�X^뉚��j9l���
�w�M��$F�5
s*z����
��L�`�*����uo|�f���M5jg8_��%�6�J.! �U�VL3�l7�rC��k��[���V_UȬo��b����5��Ҙa�Cԧ�UW۱{�>��˛Q�#4�H�,�ꀑfiyD
��~T�s	�%3�bN��24[,����T&��Z�g��?�o�2�(�68<�zh��6`���b}��h�����\�t"g�b� �%p"U�e6STJ<�vj#��F���
+�U�;3��Kq(���~���m��R#��zĖ~�14O5���3�p�p.�}��i��j�I��|Ex��zg�}K��|�=����p5a\g���R�\�׹@��V�|�:��Do��y����\��s����7�i��0$�Fr���'Imfb���&��륋q��.ƹ@�9��������"��J�-㟀0Y~GX
��]��.0�+�\|����ԑř������L���R^�M�	�E�����nD2x�����ix ��鶹��ܔ΄f��D)a�K����.ם��$Z�)������V��IQCT�g�����A��K̳_��(��FZyq����(�P䵿��
��eL�mU65�l�6�\���1�V�e�h����c,�;�` Ҫ�GCT&�&$<̝M��)��v~kYw/���Ep��S����
u���#_!jT�Q�����	D����$,�)q2��1�.uC^7x��K7kq"�}{�z��F��+�*J6B�lPn����Įa�15�C��۫xp1?������͔�܃�8�Bʪ�v�+,��]������R�4�j����B�}4}�I�(�-#����v�Tp ���9U���==ڏ靷E�h�C���냋D�S��EkHݍOk��_"{�gJw�������{!����E*?��)�<͕4t�x2w�}`ǻ��a#pKˉR�F��f��/2%�w���4��F��4��[M�P�ĬA����@�[BY�0���|�(�h�^v! ��(�0yu��� �D�+|CU��F��\�,��l��x6���Pgl�F�RxV+�TS�Y&08NZٳ����;;���8�S���;S�!�5�XŹ��.r���K�K�:��]��.*S��?���5��K l��P'�����TW���x�3S��_���M�v��|�LPc��KjC|���!:�č�)�uS�f�H�U���p�!�J���&7&k�^�� b����{� v.� #�꜄����z!�F#�C*�J���G����Wmp���x,̠�g�+w����ڻ��"��4��t12�n�����1���8pa��i�S_taJVȇog�-
���������T{7��_�l�4���_���'4\d�?$n~h@t�|c�ɂ(����ƨsv�c�oH�9�.H�ʐM40�a&ĭ�M��K�RF��w�s�������R�;(�J�r�$���,�qV�to�J�v��_�Ϧ#�9qT%���˩��ϻ@����C����{YI{OF��&/�Z9ȸ"���by�y<$)!�������]�B^/�����cϏ�֝F�f�O�>�'�@�C��~!T�k�i�x��`���9��#V0�7itp�QqRip�D��$��2Y�����A�m`���![~��)������ �N\ �ׄ���!�yH�{x��W��V�%��� s��N�V�<��I^o)�~�׮�����`�*S$l��ռ���&t$��f<�y�'��a���Χ��ׇU�c�q�	����8�G�|�Ժa�]ݝM��L�Q8V�n�����u��Ra�`�s#V ��˄�4���6�����|/�������%v]ѳqvW� ��>&o�!Y}�[��Nx�6ĉD��zS�F��>q�F�7�]�4	#Ħe�᳧s���}.iA�<��E���� vMR=m�3�	��h1���Y����+*ꨵ3�݋%u�6�öv��BC_>g�52��?�R:}���җw�P#�b�Nl!���+j���(���N�e�*7?������'ǯ��tė%Ѩ(�]��,�} ��Zf�o�3��`�a�uj�Z�7
�W��Q�y�˟���@>ܣ΋��k�Kȋ�Y�B���ԗ���j�?�Z�$��Ы��]j��]3����L?�>߽��"��[����5�K/T��H�%�=B�=430�dc.�h��$�Ko<_8�� <X�I��침
eӂ�� ��d�D��%ϡ��'�;�ǴS�
�cV߈l���4^x1>/D�SÏ-�l˄N���i���g����h���FD�!�-��$��T��h�_[A���n+A�Eu�Rq�Dv¢�`������z�~uG0��	�4��=�6!c�u�EiU�[YuE�S��$���1��',%�:�y�)����:��B����7P|�-����@��L�~� ���A�B2h~�RMҁ>��~�D�(*��4��
���?�-q'q��UN~RB���)�B�!�3esr��Ͼ���^�˗I\�~nx��T�$d؀+��*�MAX]Ͻ\d��8#�!�0)MͱP��6`k��9]�z"�ư�$�DW)�O����7�J�S��~�[Z��{���߄������}&�c��c���]ֈ�}a�%y麟�=T	�l߰��(�'%�����ב��N�@ϸH��6�����ȳ�l �	�����]1�!l�Fh��0�qb����Ui�$"�+�w�p��Ɍ����:�h��El�;��/�d�k�����lt�YL��Q����	٤+���i���?����Tس�d�i�KvXl�������S{`a�L�V���}�O����v�:n�J�%di;~x����E��=��T3R�/��:�i�v#L�ץGC�\2
������j��QPm �N�g�����6hr.SGdw*� ��a[˲/�X��$B8 [�It>�h=��<>�?7h��`�MW{�|ex�e��l} C��X�7��R����Tմë-l}=9��kG�Ѕ�8uu�r�
�r)��$5�	�1���}��EP>L��Iŕ���0�Z�~=f����
3E>�Q:aSZM�I�L@s�n#��K�̿M��ʤ����G����TwB��W:�%���c�XU�.�9��揽���%���9?�&��|�I�i�x�`~�)G���F#W`/��e�Nj��q��c��~Qfq�TH�cp9����*Q:�;HJ�I6��2�~fT/ �Z���B�"���MJ�x	�iƸP����MH�G4Iȉ�r�
D�>�tw�V;!c��=*f�
�`� ~Qi���l�)Ρ��e������
����`�W��=���j��;��t�K�@YĦ�G�V��еt��i^�j��7�����:�U�aW��~|{R�`�����y���� $2��@������w�pJ�� �?�	��gv��#ɝB��V�	=ĄX#Ǵ�|gF@�8<LL+0����s�A��o@^FJ/�ߪ�dñ�w�B�(:X���<zVqn�q��������9��A+)ǵ����i�#��z���㟊�a���������[AJ%�+���l������'�D��(�w<&{���b�>�f�fw[�:�WYXB��[**#�����p#��̫�ț��q!����g�2	�y�Ҭ����TY�`'��v�a;�Ө�� ���[�D,�̪�t#�j���o��f��q�w��U,CH����pN��I�O����w�1��c�$�(ʓ���F����Dˢ�|���,֓"��5Z��}XC�T��\�ݕ���h�]e[��7�+o2�ȫ��n`��B�����d��qC���;XMb���!�A����,gP��^[�!_��0/��i��ײr��y�S*���q"�'��AB��i���P^*���<*����D,9j�$nh ϓD ��o!0%߳pT�0���U�2��3Y��~�?���0����>OS���k�w����c1�O��dۜǿ�� Q'd`���U�u'����X�r+=p��g�qA�4����;N�{�I)O4g�jүVy ���gP�g3;<b�R�߇i���8�S�]����/�n�$�O���Y���Z��!|n���l�`��@0�����1^�pǛMv�7�t�wȨ�^�h;�±���>�]��z��=b��i�Aa�̆D���{'޺^-�h_At�2^(�[Hu�	=�NN�h�X�j���V܅W7��8=�,��	A���J������y�,�O��K��~l���nm#�cU�!��0茡z|P]�e�����J�\���]�>.�.����Y��QΌP�V5�#����W�=>�