��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9��m������G|S7���X� bU��5V*dFi�0����Y���*�Lt�e���Q&�m��9�-�ա@��H�v���U�D��ml�&��>h6��G�ҧ1�T�K��?׫3u9"�ғ��KG׿\	�"]��ʚ	P�������������"�T��!�����i�*�n��d`�Ƹ@3�H�*"���d�C*�r2�vb[P�%�_ˆ ��,.�k@h��O�[ݙ������,�t?8��;)��Z���wC�Af��V�~D��騸vD�>C>$��MUP�K�݄�ڙ���Шv���.���>3��o3��������~$ߘZ��}�TN6"�M�DƯ&W�����xgNIH�o��Y+���]�Kt��9��,��=TBFL����,=s�Z�]�,�wD�4Bx�m�T�'�}T3����|�7a@K�_��L';�V�X��%�͗���b����V�;o���/�K�s���H���z�`���cŚ����X�!i3�~_����
�JA:"�N�m��NQb���7H��´՗�$�KO_Ҫ6PM�68�K�#�9�!
�񉡬/u�H� ��s�����E�\ ���?�'��� |Z���:s䉟�[�F�E����M��,���a������f��C�1_��ֳc�EҬvt�������:��G��F>�<�O����\˨uI��<��\W���� t]*K�Bc�ڠ�&�����2~a�Pܜ)�5N���æ�E�����Xl��&
Aw�5��ېVP��H�ax�+BSB���*g��)�D`!yC!`|����� ����ױ��a2�R�؃k���"C@����x��|/
����)�y�._�C�V��0�)JO���u÷�[��.�:�`9�4_�q$�Ð,я���Z���]��^�}r�A�5�o1V1�u�2�@T�G���m��~�x�����uC+z�����jGơq}5)����D/��r"�O��N�:O�$	Es4���WĲ�=*��r��7���顽���S�S���d�,:�>��*C��Qo�]�h�I0n]�.��1ٱ�R�.5��tq:��`y�1w�8�S����Ȕ���_RwK�HTE[ܝ C�2��j�1@�E���̚r8v�~��8��@�@�r��5�m��%�74?= ^�	-a^���)~�R�����D�5��k�'A�&�6˛�፥�9��F��<��	 ��P흒��?���z��6�������p���Q�q�o��`�\+ǵ��<�ߠ	�ɺ����l�l��9��:ʾ��Q��r�Cu+��Z��әǇ��\��8��&~#�
�Z�p��Š�G��kۅO:T��oAy��c���MF6z�^��$�=����G D�i��i��6��H��������y�.�-#�Q^o�0#�e�&
�(9�Hċ��g�){�,��I�5�C�����j[A[��f^b���?����W}Z2)���-=��'g��	/��;�;+�3<2�E�Ӟ��h�B4t�0E8X��Y�*�����.,�(X�	�]��7(�r3Ԟj�sjT.;���pZ�6^s�I����VQ=�n澻7�&�������}���!����_��'�ϖ�$ݬz�pv��'��3��OM����J��)���k��c�`7z���lݩ0(�p(��I��V�!#���t�r��XFs�x[;Lm:6�t6"A]\�h��\����#c�K���7��{���1�K�1�/כe��W���8��P�h#�����o����>0�y�RR��6�/q��b����fI��Wd`��Q��ب|�-��X��K�Rg� ���3u�I}�͉r���HӨ�������D�-��#��Ơ4����Q_�z��@�O2�{��{G���V� �����\j���ɳ�C�(�����ʜB2rH�Ҝ"'��K����'�jܭJ��Sj��9����2N��q��Du(�q�B���H(�l�n�Lћ�h�@��~3[��pu�8�-���~;\qk�5rwǻ�c���,�?�l؁����R�F�����q"&�g@q�X"���(��dq�ǂK��L�jL�����x�z�LHZ�RA;��{-Mj�pc� �0Z5�[��Y#������/g�h�x�*=R����R�������i�y0*�h"|��"	��oI�:�K(�
?;�������F��o�"r�&��_��U�$�H���Q%A,g��7��.WP�渭[W^�;B J������>��:�$F��g1QR�A�^����1�թ���O�K�,wa��21/�,��St�čG����|Ž����wt-�i1]�B�K�?%(T���@
���'ػ�(��EW�e<��B0��gO���h+������Y;�<�����X̡s���#��\ҋJ"�`TD�т��"{	�;n�z`����	��w۫,���t�cȔ���R�����F���V��8� �5z&�d[�4������I�zb��N�H���]O���~4�uv-ל��L��]�F��� ���N��u7�7��<�[W���$�7�x9������q�)}���D	P�g�Ւ�얹
�׼3۬͌!aN��&"�Ch�tF��)
i�=ӯz�`0O�)XD���x�<{&8���T~�~'�Q�Η~x�.�&o%"W� �u�k��]HU�o��S�kD�zܑ�W> I�^���z)\���&��S������{�V׋Ɗ�n2�4�nW�Ov܏����@-��r��mC�{2��V(N4���
BQ��a��m�5�yÛ�F�=�<㦹k���	��~�������?�~���I��t*w����=\Ȧʽ�
`���{��+m��]��������� F�US�f��*��ư��eG�br��z�;��"m�V��< |r����P%�̘l��
W�X��9�J����^���V8}O�ֹ��:Ӛ��h;ݟ�:DJ8���'j����+��P��m� �]�뜀l��fc��c"����xYL@Ƥ��%���(r�U�FS`ЉNV7s:'���ڥ���h���<��)���;R�W()���յJFY52Q�v�-G��|��z4��P��q��RE�n��~�p�[� 5KzF("JM�N=8�g��IC^]<�Rzd\�,j����>f4�A�ױ����|g���\ �` ;.�X�)�K|�y]HېFq���]�L���~��Ugo��h��"*'�:[Ū����1l��>�;�c��X�s���f�G��	����y�E�9�c3_T�y�t�ܝ�G����`1"#�Lk+`�{�!���q׏�D�ƢG�e�����.�e�N{��g#�Sꭟ]: