// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:39 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RI7SgLk8sqaG49ZF4P4I2HnoMD//3FQuubJraB1GJBBTeV5DpnF55qXxw6bOpKKe
/Moc6iWGu/4kDRXeqCoSS78Sy8XEBozF5awz5DmKj5COZDcpQW7ZV6Z8nbH9CRb5
T24xycwcE/+A+/47zft7z9dyX6wySC7x2i91bK841Ik=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8400)
7V8dTn+Z+XRv0js9rcrmafqk/HOIN8mqcDFuQJLqJxUSgSTtm5y92C8XOL5WggQs
ApxcVlOd5jjJnTbP+HRcl3GiWMaYh+U2ssSAr8Ve56arTC+D3zxmmc5/He4umIjA
jwZFzK5jw0OANgOx53VDEGLoBBjjW8DIeYiBdGT/wDZ+hFTagp1mT7YF4BT/+hRO
VSJbfKPMlxFM8Jj2nFIXdZxzwpCJL3Os7q3sPIE1HiRdx+UHVyBWFv+XwAh+3+VF
RP64lVgnZu3jnvlX81tzTH+RrAEyTHa4CtgnKjFSHfcz2zEU1USpLHFlSb1eoDa8
csxf/+jDM5rFGnlNr0YRopwjBPWiiidqNcUE3G7qNGMJcl6nhh2KaWieLyAxVjxi
SA778ruq6JYYZ+roQ95l01/vAkrQeamwz483RGJaWrMuQNJuSBK4tRTRRBif/xnW
OBL++YPwOsyu+CAnuWI7UxSG51yE07BvEQkpiJIvxPFMdEkKqjAaQp0TAcPD/rGD
m9J4lr/wSSxC/8Jd+SxnZKq0ysfG9E6FnBzDV47UID9Ekr4D/qDwM3nipFh5CrjF
z4XjwH9l7u+KQWkL90f+ay2QA58Xxn5yNxMNl4rgBRM8RhC9nI2mL7GrqGgVatKi
fVHgejDCNxr6cDisSWVEPZ21cxoErbR2nsPtFE7ioB6JynUnSy8kOdJ1UKRvD1qw
jH5494yj75N0YG294bZwBl+u3oMu4DOY68Fryvz61Yqo6J4Cl9MIbSKZNTuRsMlK
a64Wisl3YiBSEuOuoM2P39pqxPl3SlrU3OVRbrYSaaWfUmQKckOU+vguziyMjHrd
QOSl4Sysx/Z+3eNFk4/4Nxli/2z/w1D40CkC47C+X8lE/V7iAd+b/skuOR8epPdI
ziQgjyMC1Qx9jwJYVIfwu8nVQn+kVcnKiL4YZ5aYW/+qJa5NCZP9BF5DqUKE8640
G5Hd9oW8Kho99cj1PpXAaXkEzLNeg9pBlDxRYKy5d5JZsrBk0zo20lcqNsEekBzb
1ntgNpdq2LVSWVfAKm74eX4Ia7Ik9ZS5McXtrFB2euap2/hRny/Dc/8SGTZ6n0M0
wkziYNJ0JEwSdztmFk4onwtlWLQfyLjWlnZD/gy4adNqw2CyQTN847ZAINzxvmcM
P6VgGC/Bsv561bGjReeSWLqYQhHjh2y3+kyUlI8TbRs3z2Et/BXomH4NsEJytrtj
n6a4wD6Z2ySFIHIMAMiXf+gIgZl13keCt1r4G9bk0lE0UFdedVFZLxp/6Lb46uCZ
FxtAPxg7mQs6w/+bLoY+sMt3l0dJ5VIuWC77GxEUuK4yvYhExHGLZQVDJ0PDpxoL
tes0pb4aEM9Sr3WsFC5f0rTdwDrWC+JGj1qgsNLh3gdIUHjLmBV8buPaLeaVOA+l
YV4YAL5ffQmLJ5rmmzHpPYpWxRQvREXm9cJaVTbCJYvzYnQXjneqS6qy1ELSz6/I
CEpWov6eWC7G3W1a98MMsxw4lI7An1uHyiLqR6SKSYFY2ou8Zy6j7MNhC2AD/DVn
+9SpVG009Ng+PIDJMeLJ4eyAYyEwifaC7krjeWoT5qqzx12XixPeV+RZ//0NIvEo
aa+MMNoN2W7BRropx52t6oXlmk0+cHZ6gZQsFPLuBfhA5p7pd+0Pr1b1r8PfMet3
aYlMXJ9WOSGl2miIi7iqetxihH8/8uq9Xwu5CxaeYXhqsd3oYhHbUyGR6yRA1wRo
h78D28NXNZ1rZlLPDztz9edZ5snsVQRkjCEaMjvcWnw1ANTPycvChlYt+zoJAKX6
/2joUt3nNAFbinYMqCkkt6ujyObc3O+rJhifmM+zkqB5BFFU7Bg8Y6P0scULuAkd
YLkeYTrvl4EEo5v+PIlqNCcLB4RrfVJhhP10IXmI+6cVhlQCz9DOs4iT597jNfti
JE1K/jQTH59B/L2GXpyjITLlzoUBAmSQ0XDNbEuDdH4Bla41whQTN0PEbjgyq8cs
BnRUUMIeAYo7Yrn6607rXU0xTY7++4X+0LfeP0YUJBKv+4pL9xw+U5HIs4QbYaTf
4XyHHR7LQp2pNzHJH+DTXwOoxkP1xSdqujDBv2Wz+oA5M1cMUkuT8G47YXN98tVJ
3FyNAu7J1pEyfFsQxyfIQkIm86ETiwFCkKJDTjjBfFqTGHz6l0vq87W5PTRlIwMD
1KBHpQHmgbB30NpXYuYhYVR62bBaL5zf0LlAnf2zm6Gh9kgNfRLTR/yJdO35XSqz
3jPmYXb6iXJBG1pOIzEXTs9aiCSXmLQQK8GPbRMhaH//KDc6K+npiDcaX3tKc7+k
qyVy966dnTSV8iNxcvUw2QmRxcRQ0A258wJw7qa1wzUATtJBFFVWbmdPvfAibUYh
+MSrzAKt6l/8cXTLtKwAEu0UGpyhYN1X78/FMbfy/SEAe+aeMLUD4LzsnbBKhPRF
4YFcxeZHh8Od1mXNohEre3LFEFJHZ1fvVRGh89UNAF5CzpjMZcwiVqGzYb3HRJz6
RGrW9xSaAyNl93F1iiMzgyIcDjad1kGV8VtfDfsG5gI6vmeQgowzPDG16DqMkbVs
wVTWl7839JJWSByEOAUdRS96BOVMszys5HLn8BJkKK9Iv05YdmRuSJlHEE7yPc+U
AlOl9Bw2GG9CoDQYL5e1J0da9qbWA+LHpZg1HlXQvnBfOgWYidw/jqwdW3ycU/qC
Sx3MiZH8sOeGhFHtIzSzR8uIvL96e3LXvFxzbX/C+TXdzbUFbXRh9tlAi5Fs7XI9
M2NF3OqFqGumkxIgr9EQ9mnvNX/IVXiE335fdkp6VgFcLuRLukD6nW9Udd6i0gjI
FRQdiGE5irn53QNPmy3x+kxzuRN27O54jVGBw3qq04hIaAv3V1Q+r4wx0vAiUwdx
KdDhZdIxx/ykE4HW61ae+5AH0WcbHT/ya+JeBCqHJB2VHoZMfNBWbvl4CuFgHTO9
Lzdm/N8FGAeMUH6TlOs4BCYp+KWZYUHJ98N/5wA7Wo74WK0Sm41qP2aoaSgat9M3
lmS1gi2qNBpO+WpX9XjX1dezRvEdoVqOBGjRqzfWzkcHFUwUgkr3a7bIJBK1r0Cd
+Indl1iIYM19b/FBd5tibKMBoVHmzR7OREbdDIxqz9stx0utBG8ra1zjwC1uf0eO
t1wXTjJPILxzcvssrd9DFAa5imPZ1g8iysAF3BDgzw1y8ZmOCJweSy46OEK1bOXi
iMhLtpAawlTRIqmNCcs2OqIVUs05D5PZEiDB0Shs4Q3IE8b8A6/1JW+jnWD14sIo
mXIYGHpH4atZ/YjrRcMRmZuXwBQzhHwYaD0es8B4RqjfyT9KWy1Sbg31auR5WFyD
5EdhPYEb11QWfffMkpHv4khLGFRbZTx2Bizpc/wv7iz8geRphUdRjfi+LP04hdhJ
aw8TKcgTR+XtYWWmoEzBUsH7oykijaqJmLtXhwSe6oS51QPmesMvJxJLRkSSFqs6
ioVMgrKi3bo6l0PwgGHxPwFvQjkAABTfthqaPjIExqckyk3hQpoZMAIqaimlUVeL
8mPVa/JOcj3YYi0Bk80AEKB4ywnO/cAXb/jdKqhVe0gP3KkESYCWvuGkMGCr828F
QAfCoKLDYiFSra9F1bC/6wFaA9KUvYDBBzO0+3hLWMyZOTZQ+ALlcMtBXiVsXKqY
buttJ2zU2SphlEcvb2lwRlF6JeqkPNrXeOjnCvfgyUGF0aYF17PFV51yVGG12whj
6hCoFlXQ6xjI7/mnvMExbfSKZJpftTrQISdveht3REzd53TcC1QSJvV3q2qqX5wh
gWjkyPWKD6kipx0SPYAtNO/rkOL35oV/wvEFe4pZFQhVGn94PssdMjK5sxBho8ou
Li7MgPaNtEhSbvBQzFiep+tm1rijMMI5uq+rbd6KlpI30C7xvC4HE2qA2cLR3NGC
wSARxnAzdTIldwDGBcNktLielK5UkBpWNNwdk4vef5eOF9xUsHcaIl209hexenSX
kIPqeAqjImlzNz5rc+G2tGVfwSNsHC3DpNDdj99aQgsxyMaY34GM83sVQ34saNq0
+cd9vtBHr7c+3slEQohAqVcCQngMfLv1SWGuo63Ce3U0P1Nq1z65tbzsn05jrOex
T8NcizQDuiNayIkNG5wgbiVORw7/12trH+zt8KpNv69ls9GKdR4Lm5EjczTFqW6A
UcmG4D7WC0abIRpWbvltPybM0xSo6NBQC/HZcbfV166b6VWmPv9aVQLNVI5KIb8u
pRjA8rUvHwF/M6Iuh5aSvjRYs58Z37BwR6X2Vqun8ShsSQY7mKzXona66U8cIV07
hbDef1lYY6oY+HH4lblr/RP0sUDV6Eq30XWCVhINMwOjjT/fltWBAlT2xvmDWmpV
/E+DgYP5xv2MY+3h5uXpaV7WXwf/sDcvZEt5xuB4gF2YWli1UaHNXM4vWuvwkgII
f0koES8uCWRdT5oL2VmdBA+4JH63khOrC7TUZslnm00go0qY7asKc5wXuP9B/on6
OCL4HRcilyBnkPpNWLja/TuQpFXrxm8uLdZYgpcBumTt4VFMjwyVsTPbIt1uznec
WodOuDscrwVuBI6jdznCABKgiKLS5+yemo3LaHBbnk4Bb028kZohgh5EOz+C8QRd
7w66HQ51ZDRdZhcx7C5ShNyg+q+zJTe9zZ978Rji7n7uvbNTo9NPWp4evRuodlAB
iQJbO3w0lKScVxpL8WGuR9pHcZkwTvgul3PYvgGb657VklCsna7HKrw3L9Ii7aPV
sKy4noDOinkwQKF7Rw7bAvk83Nc2kYROvp/b9WbjxZI8WjrGiLIC5l1J2cwsluPQ
HQ2WrQHMfCu5R2mCRLTwYpzY11HWeJtA+j78mOJ5ESJ08bj19i/hoLOqylzO2eV7
NNYL4bWpzhjEVI/JKdLel11ad7qUnoQA2WQisp1UUSZ+5Q+eB0NrzYLcIYVRmxx9
/wEyHegPgWOxOp80J+mLcZu33WASwv5hzAopbQsKDAQIUDZnjVQRAOYED+8r1FbV
AowdcS7kuBWertvidgwrZtlASJD8eQ8hQuJ315KSkSujk+tsqMSLXEDzHt3d0mNM
Rp4FEwDF3F1C0XIzvHShcaoc9lPMp/H25tKY9yy5FjNj9TfN8cBteufuIXr/AanQ
nJtXNcbFqpYWUP0CT67jOrC88utkUVy2vySNB7EupYhThkEEVT0ePuCraKAfpQCD
9EhxvV3IgJCY086rIJDjWbo0Qg+wGSKeMpgAAZMDn9ixze9pHSazFHvjjMVbmFsy
1QTheZlsDGF96LUp1oG3Lz9E2nq8nWu0AFuXgvulwGvjKAny5xySxkoWoatodKQe
m4Ql0a5fRnpTcnYkeXEOjkNdXtqyuEDIg3Srj+FZM61BCh3wSdlKrShT6vsBZcRo
5thn8VrIdWIoGLQn+pwYQluh03FOSIZ/EcxUyLaXLs+tzYyNopYVmo4ZQFv3d2xo
8lwqhYWdaEjmMRgjgHfj//oY8d/RlYimLHB1Xi+heeSqIM/fb+IO8ZahBSdX3Bn0
pvMLg5+FMBjSmWJ3/PJpb6m8ZLhAKpE/2Iuz8bEfkW9ZdbO7VeofvvMurThl1/CU
J3ehHPwUV0qKBDTz7kkJhLHKJhdtOzBzHJ+k8NR9qRdA/AINzPcsUFMUydX0gVXT
TsaZ9Wuy0apPHD93gRVh1a8ZM0NiUUNhhLKrk1YwjE1UhGJsGgWw65ZoZXRnXOGM
vDMIkJ0AfdT0GCq2/8x910v4VyRcRCV/SWOBEJ2Gzs1XDcojvlZUEW9pl2dTxQua
z6id4pNlCgInjbXV40LEXMUVekXsVwAEOUL7xhYuic/bWWqvjb3XFUm+OIzSL84/
BPMWZaeCbhamHMksDNsuzy77s2UUXR1kqFLw6xCU+vevfClqqTZuHh3G4UR7+r1+
8WIZTghK8fkV53mB9Ikdj/oQ0ujkSm7Ay4ke5+tzfjfv6cw82Rc5hJ5mzqt/IjHW
AGdCQiwM3oTtpFk/XBVjGaDlWNxca8Bm2yO3o9AdUHFabOLeJ129HSI0tHJoH2L9
bJ/EuCV/1VxxbDA6SGmqEpdT9HYweqeI0w9yL3187FcRAQRsrPpVAMdPz+/vd7/G
SuNzj3f29ujuPDvoOjDGs+c4DCwhgymseueFteVd/RJGF88nbmjl2no27pQPhQM9
ihBT8w/Uq/n8TXKFuUkHxStTwSc2pWCWeW8ZmYecIDLwPkDSQRSEv+L6bKSlxMSS
xnGeVFdO5mwRtPv9jgipHYMaooUXgJsgAA1nFO0VPAO37lt+kj/Sll678Msx4N/Y
7rRogqbB6kqmOuG1paxYusX3mYpDZi5JC37SprW3XP3ZAS5Ks2ynIP5iGH82RiCm
Ry0PW/ACNcRhqEru0EWQkENGInVx1/PlSlcu6ANh3jtkmzoIf4JKXyHzPL1oHcYc
xJma3ocePND5qMPOLPYahrImMstjb6BlJjqu5WT1ra9WnWhkKeJ6zCscHFo9st3g
kAijN60y2QQj0k0ckTpKuWw6tV19awwAF+8wR92x9lsMajgO8Cz5qzTMQgvemenR
Ws9wZDdQ9575lJsyWgScBWXNvxu7CuMJ2WaEpeznQ0vy95L8oEf1UToMISBQJN1F
3LFFxheABR1+VMZnQGKZVgxVwMJLYDhnhzkZSyQx14oHD3IHgBtKVpcYECKDOri8
S6CLf5z1vfPWnnAGp6ia64MMeIhsnI+eLvx2+LyYbfUkTbECEA0DM6Z2f2DCHJTL
2+fsP84dTW02RXhQaVSUULtYbqt+JOPteUrMUaLoFJFiOYacRNgXfmH9ZhpmEcpy
8EyQOodKbipsb2jSWJS5cUxdPLBySt+Vi1GAGDMUfU3836uNNxW8DVC2dztdGOQf
fGO2pVfgLT30sT+czFqw+LWwsoSxfXBXFVB4hziSGAD6YJYlc5UdDFnU2J3j4uPX
G7VfKlMkakfKayJJOOyKo1DiPTiXa25H37zJp3O/ZD7HHLgEzvzwPs0iG22NddWh
dIXTmetyGVMtN0kKSv+xaeaB3HqKhbBqTsUSpNA+US0LJZdNkseSsB50I1qv7HTg
BP/KCbSuafu1roXMQ9SvVZtLzRO8JYRO9v7UXEZhmh9jhql0AUJi5b270wAlL65z
0pzap2aSAs6W0qqA2SWnrhkJk+xcIZBpuY/fSq7SeMqYAY5VjuWTwnh6lpUsw1Pi
Bli27BQf3juUcV6Hfi/Qu//1/v6lVQvXA5wTvpBm1YPTmhtW+1CtQX1wfIheIM4M
9aKGK5RrD823nQ68MNhBfVwKbQn34kN6LzvWQRGue3WP1pPxotehmASv+F+H+cpw
Bc2I1TP+ISg69Y0habpL/1dqpC+Q8yWwEPuXmuV3yzC69lyK2eOsF5HOVxPifjDm
m62ZBVpqpydt5b9qakLsBx4ZaRVhpbURYTBMkiSQFu1usPmkkZ94oTBtzw2Mv3mP
t26BJl9vnUlRdXFUa8JJ53cqeiEF8twMUNNPFLeEXNpw9TpshqJGjDhOYPTP1Hpg
7ttMIuz7ACbDK6mE6b0rV+loMR1hwKEPcwTlp0nY8VwyualmPq3JM9fZIoMOmlPl
JvB1b8W3ukYXb9aaqkqVwZAlNghfE4tJQg9JKy1qzzTwLxbxttAEbZrPIhKYQmyT
x2DTxw9IUTrW2m53SKBJODHVnyjnJlkRbM79x24+WCK7/o9W8U8wPSMZL6UzGNoI
8KtcGfk3Ibpmr7BvLoS88qjkP6ARXOLi6Dmbzz972f/sPdykOlB8zyNjsUXb8676
86/Ok+jHlEwgJK5XRMu+WBcB7Rz9VEjdtgzNmCdE/V3xNUs3f02xVJaGipaeDd0M
e1wt3sgz0axOGfmGlyyqdSnDWQ0O3eNRXxXD7ps4kZJu0az0voDxCpEPw5g9CysR
rd9t/Zv/8ZCOr+LtR+vrjY7UGnuX4Q198a/z9o69YZXr2D+4c1L0fcNZOhNnhj1N
nxYeYk5LklGinpBQMkWaVCM3lOEZkoyL3htnMkLUQBkv5xXTZGnziFgtWLiz2SZD
/PDVRWFhVacJVICHAYpoMO8mV+htLZwGu4JdHaU1pFd3jSbuPPczJNMUo9gKSx4Q
oqoQWEoLSsWN1VoBixGKRgo7OGFylxQaiSuen2ozQHwKVI1gOKHC9zib4SQ+sS9u
D+qzkzsjisUIffVk7P37zLt0jgkVVt/i1c2MuOPsiadoGyehcSfpVSjXKMA9Suky
gghzdiML1/VWsvvUwsqYTrM35mKjnQ8AfMZM/rGFJV0abfaKltV3+EA+lVGd/04B
5FNg26TURmxKckFwb8Da/m0FYlvuJSjzTFBLnIMZgLGj2GnVi/N/uoE+c/SqMnmK
8rv+prGXCRwLcpeX9gaNAPyWrV7eOvRH7K8gO+86xjjPwK0VVfa5doRVvfe9vdjl
IZ+Jgdd73YzIZhd0iItoHH5/ULw3NNUg76MtlkHnFwA43X4XQE2/KdxktmyU28df
GbcvrCvjjz4djbS83GSXtObulOFnxRI4XcGUg0h7fAuuJZcm19XcSDVT8xZ9vWcV
oA4EBostXWPIJRSahK9FRknKvSO+wskAE5rFEk7FImFXNt5Y+O8om3g1JAKbuXh5
YpXgFVvA8+XVUdPEcAeWK5nHNu/+schwp7I8OqKMj6Cb0ZWVA6k8RpWycB/jiPtd
1Ce+UYlhvMmMbfVJLBT304ucPcZ1BEY/YEq2MARWHrb03nzgTtF0jWYRwOn8kNNt
Em5oOypxcVBuMDDmIXCa9cC8aeG8i+PR34/Hd0VybfB7/UX7X0TZObP5bMCKutPl
pxWqhrtYcZhXEIJkFRzg2kvObU35jI2TXmuBtZTFI1+6OnuYHHgcgQvD3hhfxj+9
6uzrmYuqpdlfy1A5/l2clJhHEFJfyqPB8FhyRSX3Mk8Xb7gE2+XpOGlJ7CQVxiTC
Ey1H0/fj6K03f7M9UTmX+FFM0ejpV1h4C2956oM0+oi78PFDcfor2uaeZ1h9i5f8
T/w/QyeD+4fu4VyEYt7Dt5jjCacPWdTfbZ75FyE0+VsmZ+MWndUdN+9bNetVwMTD
NieZfp8GDcyObDD4R15w6NApVu8I5MQiyUJEPnWPOuOY7hiMqFRZGqoE7e2m5w6s
2mpwGWYD9F3Pu3okslJJSTNByQ1ONTG1gslI+cGfjBUb32wWQlA766xUtmiVRGaj
Q4IbKDht86Z9o+JMySb/4Salp7meVEj7KXILJeHdT0BF5FL6FrH/zPiy/+Hgr8ke
vLbOI0i/9FdtdzuZoLc4Opa6Y+X+z1tPblJTDC2KYC2vEboEPqLP0SySKacy8hBs
YLBSnQsTsPWWOgCWL9gRNJkmKqUGIL++jQGm+oQvrJifC+iQdUI5PIKQFWBvHQpU
Fhba2ZTe9NsgVsCpkyfltNP6i+ozfZEXh9E/Ir+zHZm1j4Sa6Xvgz/h6ncfLdyOj
aI8+GtWvVZhmXg0vAfpJVpvo4jlU5+tIf/Vw0pSfY7tmUwvQWIV1BK1PgCHWaNfY
uceqdd0IvCRqYOS26GIkzzQ4nmoZCXI/buYor3K2gkWvbu4OF/w1ExoBX7CW62+x
5z9fZmS02lshrwM9n1Ne467WdP2GkrpasC/yUPWI8FCzTXFy3pHEMOwqdnR6NILL
/9YIFir1dMGBcsz0MjfPTQatrD5rMNSfuEoMcROeQyR4lfAiDMN9/v9P/Hn4h1rQ
837e/NgGSTH/IaPVovUF5Tw3FNAKloL6rFzLPKDhY/GaZaKsm3y7L8OIfEStSRUZ
yLHESWUboviChL+T+qKLeRVj/dttVVBqVLp/IHknnXQ3ok6tH4ZrwIlyn4wweJX/
PbEPavT82m2wJRaP+JQb9v0lmRU518PaYkb1C+wIa6g8hNLihQWAcdCd2drwCMo2
BYvgtYpCXV+ETPvPYbJS6DClHIMXF1PodCqdNDWBMQWTDSUizdTAH2RSwbRXKC3o
DlLOV4JAmvRxaHi3KaZ+iKXkX1PqopiFMRw0iFe/P5itIEJgyWXVXZ4BBySEK4jO
RXC6GFzDAp9//kLQt9c4amu/qA7aY6PPwb0Im9mrvnXw8P5Rl+bROdjD2Gtq522a
+4R05LsbQOp2dtaWqy3qSPrizlRxKTbm+tfBRnL0TiottH9jpNu0DxdmIHQFT3OG
NLDO5Ngf6Vb/pQG1S1rNeayKt26Ate6S4cXVKCecb0D83spLn91e0weM9LdmjK6K
zmDqDy8QPAw3b2cEdFAXNvXVhNg27oNNPb+8Vz6StvRn4YTCd4rgqYD/hiDvq9Cc
kGKCNZ3odZBsjU+5Yndls6UCvJrRJOAACquoySVbrqofyItekrGPm+vZre7Lc+Uv
+lwmMqRjzBVxtVHvlSUtY2Xn2wupYQpEg7VSs6YyuizZIHF035X7ZJWyydVGEH+T
aBVdMNBSjV5RRDF0XcvPwNGWUvnHMnXYV8P+Pf3oq1xJDsbVRGF+Cp7jJvyKP/NQ
2FhFYqP/VINJ1ufe4SNl6+QOrjDz0QZIxWc5nZaqalljicxRBNfagUDsXVHG8x/f
pVh+UvtqSVFotQaCeQ1xFO9sXUkVOxyP24UicTUL6+4svAf4y3/tKytteHRlnNNQ
dYg1g8Q1YhOV++XNANUUhqJkf0LvjrOiOPB2EhcA72yXTeXLiDx5/52Y28t5OzVW
JDYsf4pVD1625RdY3Ygp2XqHWZPv86HIgh198fKTVGqERSu8n7dPPyshw89aXcwX
zB5ROjlWfmKnFR7c9P9Y+wmlEI+mvIpG4rw95cUFvdftjWX9+enuAsx7PQjp1ywf
HRNTQ28ex9y69kWAZIx9puiXR8pmvAcioLXHRz95AvizuLpeADlPcZsK66Q8+Iyp
yZ0Sy+mmhXN5vFoV/I4WHxdncrCPJbDE56SAeKkxbh4+Gs2xRirhZuEQs1PdaSYG
oEas+ilhMkjazD3qhU4dhZBXP16lCLyPJdaOUQRfKCqx1pLNGVkN9A4opVORazKV
/rXaw1aZJOmWJUqCHq3AJiW9Qi20S9sb1QOxr3FRCOoyIoqQzvYRmIZmp3jqzETd
vXN+cx0kaOQcaEDrx8eAKhKnzL7N9S/aEN/X4aW5XXlq+m1qsERCyxlYmS5I7Wxl
EWBczr/K4HjYWCh2x8SCTody7V7rG7IkgkBEE/O8zl25S03VYz4HkO7MoRUvk3vJ
3mszmEwzXw5wt7vWIatqGLn30BJIUM79GQwwNZTBhD0DkB+ynzKxsHq5IjO2OVxC
`pragma protect end_protected
