��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}����ٛ�!"!/�NV���slP|�NJ�*�C��H�5�4�h1�W&X2/$1`�Ր���������)V0uI��?/��_^ԺLi�k��{��M\37�� ?nՉ�2��w��KR{�����	^��V�G��1W��9�h+	�-)[�舆o"�_	�8�Q]�1���@�<���б�v#�i�,��9Kl#�@���V����ѩd��}�������@�Q��� �\^����=���M0�%%� ehQD�J6����8�`&�i���M����3��V�|{T�1Nɑs6نC���G�?;���;O "L}�Wܧ�J�%��͙d�h��5EA��J����O�{y�YM��LmR	<�#����u�m<�֧�+� 2��O���|��F\��aL��ֿ�Z��wOl}��7 �
]B��r?)�3G��j��%���y��|��+�W ۩jf��'����%9�+�t�1�˝��������޵�Q�b���:�I�U�0���뼴����I��$�t��W��~,y/��~���hi}c�[6�	`a����E��Yu��j�:�'����6���*��=T�=����`}�2�I��"�x�U5d5lj���Fe��1O8�"(Oi���.щW�(��N�E�`y)�fc��OԒcఱ;/�/i�h���'�T�NJE�UH�Je�;L|�����l��R�E]�e��w>�s���g�Mk�/���������s�@�s﹖4��+�@�x#HS���,�{����<a�qT�8f���q;`�Fw6��Z��Mw��.�a��eߏ
Y�z�k�@sH/.�!����k��^a���j�+%nA+�~[B�!��[kjN�8 D,��J�u$�\�e��%n�h����2�9>$�d�2���G�~B�nd�8�c1����e'fg� ��cM���`c��G��f2��=JV����S��Z;~��A�X��/��>@��FAD �Z�xo֩��^
݃��Qƥ P��ux�v��@8�6��CL0�[:�?u@�'�0���
�����\#�Pc��j�%"���P���޷w�w�����/y&j'���@���&�Z6����]��I�8�Xs�B�V���$.����������������>�*��;�Z�,�%d�g����~���B�Z� f�^������B�rz*n�T-�<SOՔ�O�3�5d�|��K��[d����&.�����i�?�Ufb��ɟ�X�a�D#"k�Q{��I *����"�p�3=�:S�9�7���C%�Al�T{�C�����ZNAR�<rc�6�Ym��A��xu��ז� ������r.x�썽&.�� -|iw����.5�Ϣ	������h�1	�M�y���g�S΀$S������&FbhH���2��;�R�)�ԂY�$��O��{Ҩ�`!�H�3#%~�i!�cʯ�o��Zx��^�/46�e�s]òY�Z�ԁ�2���T������[(!zn�����~tYv�+B"=�q�߆A�P�g*�A���c3��L�i��a�˥A�q�{5E�����Ri��(i��D�I�W��S�.xI�HhJ��z�G_�ڔ�e���M��~��]l����xQ�|�w�t������� GR�yLԇ^�0i5����\q��a�a�����bVȍȴ:�G*�K[�'�u���F�*�}2�HǤo��\��v��=��=e��K!���/ۻ�3`���	p�Y ���?T[��`��gX��	��ϴr�=��� I}V�wUis��G����˽ي�SN��E��ُ�z���#ԉ��΋���h2`�y��n���!L@s��Oh�@����{I$�=5���|������Sd�4!ݨ������)�l�}<�0�w�=��+�c�r2e7gzͶ���Zު������*�� k[���	YV���n���Ku=���%{P4�&4�5C`��}Eܡj�7������{�`��D��܎yֳ�#]ڐ�R�?��B��@���&E�:N�����0�����	�������ʬt���g��؞c��n.���q��CyW6)��>E>ũ�(}h����V;�8�8��6���C�6"��2!(mJA�T�i�����~�Ĺ�Ǉ��
s����l���[t�r�F)��22�z�(wS�`��� 6Q�@��s�X����m7��k{$�$��Y���_�?Y ͹h��y��S�.���n��)��S�K��U��dyOΓ�� &�0���c�k�Ħ{�=�}d�n~n9�w���O�Ն����o��4�Z�����h���"��z� �7:'�3��K�/d�2����J�/n�Ha����
>sa/U��XФ�o���5�nѹ����_x�Y�4���Q1_0f��QS�i���?WQ���a��">58B�U��"�\P����4���6ρh��e�5*'��;��,�<eRލ]t�Pq��]_�?������t�h��B1{�;p�2j2���x�Ɋ����Lby�&���4/�͓�0j�`s�w���M��V���n'vEmsgH/)L���Q��z����;��A��ߚ^�lI�q�0���a��h��a�I?�e����2 L2..m#U̡�Θ_�gr���l�e%����L
�oߚ�ҿ��:�QSH�SbGc[��ΑK�f&J�.����X^::�b��^�;h-�z�E߂u�n�9
V� �?�4N���Ȓ�7Y����&��soͳ�����^',��3�]�;���/5bf[c�#)�d��0���b=���5�P97M��f9r_e�℧|RثW%?�#�YX_b>�d����p�,�v�k�-&V��Fx>=�k��]���s B�<.�5.E)lk�8����:Z��@Q��;��)(n��qi�]]{K9HX�E���҅�卓�qݽJ�P�
(ڹ�5��z��Ɔ�E]o��53i���s}��Y}����8���L�c8�{�m�v�Lz������<�<4Mٗ~��xN�˵�qUPc��iU����J��-��lA�ִ��g����JcB�!�l�a�G��o������%��Z��m�Iɝ�+H%W��婗�2=�(�1�N4zNN�ǁ4����f>7t��ׇ���$�\Es����*{2���͆zA[	�ݬ��D�vw��2`s��P�R���'9�HY,�ω�^B*���o3����s{Y *5C��Y��)���*�6I�;�G>�!��A	J��1�d{�T_d��K�T\�n~��H�pU�c�fIP#GsndQC��A*�O�����S�PS���%
���yVû�~*�^$����-}b���5� �G��3O��R]�I���Y�-��2�t���`}��0dmj�I�,:⃲�c���=�g����ɰ�����`f��fK/-w'��*�@v-�\�ѕ��/� qn	�ڡi�HU�������c��*��a�����@�����z�3`�� �f3�@�!�����h��M���k�N���@(�g�c����`�}9N��<#Qo�T�&�<�w���X�8B׫�ۉ�!Zp;��tٛY�P!.cdP�C�nh�oFY�bm���\�')b}�O�(�5Z�Id��.h�`�_YlWt�U���%�ܮ�3��� D���B�똻���v��l����I����?��J��dU��T�`řd��K#'���B�nq���z{ ]���0�H"_R(*� ��	"?D>��������,�ȝ���&�X��,">�=��H$B�b'U��Q�#X3B�2O����7�����O1j��@�I.����G��1wb־י�`� AcsMѵ�5:��c���SX�x@�k�0f.
�{�9ӏM=�76Li�za#����F��6 ]���{+ێ�g�:�%�����P����z�4�O�L#��A�*;����zJPQ,�A1nDED�lIX�r��Ω�N���7���:!�>����џt�D�cs�!�����88�i����5_�q3�3l� , WP����=P$���� Gv�S8`����>��id�2���e��w<Zy��jD���ޑ�p"l�l�q����`���OXػ��l���#`+g4��5���w"�f��3��)	C��.�Nj�&@/�4�7�[9���F�A�,��t���P�c��R�ȋO2ͨ��$�Yb!����>�ST(��1���4�:D'�����4�~�P�0L���� �9�8�)6 ��W��#Al\�%k�EJ��7�6�V(pv��Kz��c^Խ�'ri��®�U�Ec������_��3/�rs�n.k�Q��8Y��q
�|�y��f�;�Y8����g'�ղ/	�����]�AT�3m7!���]�_���tZya��0&FؐJ��-��!��ʛפ�c109,1����H�w��x�����08+��.�>�t�&H��vpl���MU�@A�;�|����Ck֕ �Px��?����<$��i��C8[�oK����A; G[;��40���y_����haÿ,��FqCtx#C�BƮr����ߐ��9V�Tn8�W�܁ a�8�2�9��n�jϯPK8�dڕ�����'7!g�[�u 8��~R ���]qb��i���ѹ���m���(�^��3!l�
El/���OpM����#�D@_��7��{��]tI8�?���NR�#P���7�]��8�'rbtB>��x2i>+$9ͳw�鮅����d�փ��2/j��E!<�N��}�bUj!�t�o���ѱ�֡ �/qՄ/}V�h%�TfكK˥"�@o��D"kp��w��
g0&O�=���[���=�h�����#Ł��!��D([_�?w�����wՙ�m�����ʔ݃8�V�V�'��%#X%������D��t�X