��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0�����(�_?V~��
�r�-����)�b�K����'�� �yq����@[g��Y���<a�e�S��y���G��O\-̎8��M#@>���{�I�3D�ۣ�q|�O�"IV�D̿?��'��:��3S Ń:����3:v\�.�r�i@2��L�}�">_��!�ji�qdҺ;YR_�8��f��F���w&,�dS��+q+Z�V��4�sE߉��׍�7�=�-�Sη��z2D�(�_l��!�]S��L�Q�B�i�/�sR�3�p�h��a:����0�\\����uq��s���;��܄q��3�K"��z��%)�U*���<�cptL��_�-���!��I�Nb���M6yE)�P�/�Z)*�� p^���X%UIƆ��~W��D���������9��?9�`m��#�C���S��[X�בHfc�u�ه�0����^���
�1I��cdt~�\6�.X�m�A�;\����{�^�n��v�5�-��8q�oL.��5Cd#N��CK���t艇V��w`�������Y~���p����_�3;0�";�
L\26����	�Z�6a𓣱�y,0iN(�4�~���7�D�Ͽ�����w��vI:lż�&,ҐW�ρ_x@b�F�|�Ȟ��7�d]�ړ�r��Y���D��PZ�XP��C@|�.�ʋ
U�R�
3����B-1����\�������7ݟ�"�z��pQHݡ�Z8\�r�3�����>��J�m����Fק��#1���x-��ăr��me�ev���I��e�5����ㅝU�O	DWQ:0[HgR�+m<�~���^�����}IaZ�U+���?6�!t�ź6޻��4�2x\Fz���nՉ@`Y��*�P��� �(�LH������R�s3��nu�%8��\��N�oB3��F�<���a��+_ރX��`g= ��HY�#��Gz
�23
�sI�Z�����AA�1����Y$�ĭ�l�ീm7۔"�p�Jڳ�����\F+XD�{�$1ğ�+p��ۊ<=��d$�S�;>����a΢�굵�6�n��s�1'.�$���8U�
_�>�\W�G ��CHՌ.�u���&�g���A�z�Z��s��	�p��/{����5}y
@�r��8B�~�4��:�w	o"�(�W��H�cc���յ/	b�Wd#��6���͡�e��Z�0�4���?�s,�������_���<��!��V3;2���̘�l�u��d�ۗ����"�����n�����(��>10�K`+'F���jAΐ�Ȼ��2h��`^~�~ץ���3v�08_�#��a�R4�TJ��N�͑���;E\��)�"��Hp���]h���wf��7�������e .˪�(8��6J�?�څ��z]R� :��)oo�B�
绲ݗ�U�Ӱf��?px�T)�J��$������i;���c�2�������M褕����#8%#G&
�N/�܁���4�`��1+�t�lv� ԹF���C��!��|g�m��lA;�G	��*R�鍽�;L5b��9����Lv?�e�&�r쭓�A>��;y�=����p�$��0;�$#�{�| |zm��������n�҆%�ڂ��ȅw�d�pS7�]�A�4+��g��
��L��5��|�i�֕�$������+�B?�*O����H%�(��N���1�=�����#�Lh���ɑ�e��إ�kŒ��m�(Z�yD�`�6���"�h>8�#����g�{k�w�J[�.�,�:���}�u�%\��k��mۆ�]S��q|�qqS6�� �K5�Z�t�V	Ɍ��[��Bu�7���v��:��k�n�% �Js�L����r3�o.��#�I���B�[�$KǗ;6~��ࣱ��m�:x
����ѐ�6��2�ȃ2�@��U�g#N�a�n�ϰ�ژ��Z�e0���UZVU�S0��<�E��`���fr:���%��8�a�
j۸�9.�%�L���Wף1�Zk�pÕz�>,�� �(�ȭ����/��$��h���EJ��y%��]�TP��E~
=�}�DM�����^7[�(�����dP*���b�,n�C��ȍ��S�o�կ? �L��>��