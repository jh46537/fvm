��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� �� R͝���c�	���)es"[��é�#�‍?t���4�5!S�TP��k�$��  ��y�྄ !��>4Y�f�j^�~���X�$s	;v߳��|g��(#���u�N�뿑8��$>��8ѻ <��)�X�R�-�e�;mn]_j����0|4X��)�l�E(��{J?8��_Ѱ�R�}�xEbCج�P�Xс�_@_R��/�����/�9G��6�9���4���2���ƍ�SQ�E��sLۭw�ķ��gM�c�ojr�5��,5�$�
u�q�Px]=O秾
�zza1׸������3�BV�%Ba��,�*�	��e�/ۤF���P�x�f�h�? ��tXkP�h6�/���{g�H���c:kS�q��V�V�LC(Tg�����mڇ����M �w"3�����A�����R��2Y�R�z7 jŐ���-��Ap�C��lp�ta�[���?|o�����4�9�<���f2z'0���^�bxk����r�*����H�HoC�@�	�j\P'� �Pn�'��0���b�
�͏G�}��}!Eu�F�T��j5�Y�����UB�������]V�<��F`�X,[���(�Y$��?ojV_Q�Pf+X�ղ�AA��-���!ٛ�`��ej�繙���.��㥖(���u�)�pi�!Q���3oz4>+/+��1��cb�~E%q��V�&��!��n(iZT��K�g��&x?`l;Yz��5/�E���?�Ƽ*\�������>��e��Z�vC@�쬽�������KEߩ(��	0�)8������uR55EO4�Aw�����{�A_#�θ<�>~d� Ӈ?���J�4k,��\n�d������ �O�bd�δ^��>ݔ��b�ԛ�O!b8�MB'�B����ͱH@E����k�Tt������'C�D诬.[��S������ƃ��&Ӓ��݁��E�0�.�I�z�ǅ#P�V�ӷ��_�ߋNcQE9���m�ѯ�*��_|�Qr�=С��!�������̈�h�OC����d�u/���/2�t���}����0�������.D�X����x�>Q���fcR�&hs�r�A��=�����.�# ���·L.I=�4�=�l��è�
���VZ�(yA;5жL ������ؿ��W������I�� �a�B�t���p��{������g�ŭc��>��%l�w��d#xd>�qib�.̎
}����J��?X0َ#����@�s���v۟�%��2�7$`��F��9�/�Y,[scjE��.�f�s�f� ;���5� ���E����*�!�v�Oo���{!0/��N��b������;h���'�8�Z,g��n�L��\pۙ��u���p�h�$z�#��J�w�z��/h
&�T*oi���g��?��[�+��B�������W�}<��a;o��C�:J��>z<��ų�����w/E�+=��[��1Gq���z�8�_h��8��,'�I��	׬I�Sd�|{w�.�H�(���l�EYq���k�0�.�j� _G����&�?�>e�Z�k!�<���@[�4�Go��mul"Ɖq����X�US�F1|�>�
�1��Z[���/�.�_3�~5�$]��T�$���WZ@�����z<�e��)��n:���f�I[IyX�����^�i��nmL����J��X�!�*��#���\��ɂw9�����o�mU������|�r�Xm؏�=��u��/Jܼ�R�r�T��1M���l�D�>��d@ՀQ�"���1K	{�ˈ�e|{��U/l2�C� ��T2
k���@��SQ ��&ݠ	���5\���d�] �了Ԭ;9i:�cO��Y���%G}yS��43c�@�_�AS��\��E){E��)%pm�5����0��`�Xv�i`�6��>�)3�����Z�`�|�|����_�ֲJ�kԧ|7��S��G:��U�=�-�-���H(e�����}�����T�4�D9���4�-���
ڶ�`�����mp�&�i�"Y�����%L#��C�KdC�����"3�%���Uygׇ��Ô۞L�6��RX�@�%��$@�`�.l�k�KR��y��zP�"���O"ќ
�)ӝ�d�D��k��{�������c�9�e�ሴ N��Fl}@��U��E$w��߼\��k���E�Q�m���s��" /���ݩ
�t{�1[%,Q�|�k��4UBݷ1��ه)���pG��uc ��yJAЄu����P�گ�������3s��^k:Q���3bc�S{0}��#<\�K�(�O,!t���$�R�Dq�c����jS�{����/"{� �m���5�^3�4��)�0,�}3�4��q̱�x�H���tߙx�vO��A:��|3��c�Q����$��
e�����bP�[���l��2�8(rk�N�z �s �2���g��X�����Ɩ����a��bT�ΡL�j��42�/�ѮƏ?�\�jS����򳘲iZ��� �tX����c
ہ��[e@Z�Ev�~���)6���W`D@��XdKt0�`����RZހo�\�n+��g�9�03h��'c�LH��P�U�&���FCNn������o�P3cM{6:P�[̬��ܷ�Qs�Q�<�Q�vM�Ph��H�=����!׿� �ת�P��Z���LnД�S���:`g����;w�#�E��;#�Y�hc��Ax����'Mw։/�Ma��
Wv�n�Ȱ����t�g�Ns̓b#'�vѦ�`�Ĳ�d��?�u#(�HJw��L��!$&�z��R�Z)]}],���#ci��+�ط�H��� �O08W��_�p��nK(�1��A��%5^�3"�^MW*}��w�S�E~�1��f��`�Q��B�-�.�.�>%�R�^��`��Y
F�!������[�l�$��������"ʅ�Zk�ƫ��a��Z�Q����k�x����m��ʻ#H�p�F�?�q�oan��C�˓��r᳡k����,��SS`B�b�et![H�&A�H�g�!rW��W��)�Un�PG���ј���1m���ф��q�)�Q�צy�h�~�:�h0eɰo3�bBwi�z ��rPͺ�,�OR����}׮Ӄ^��)`|rGs[��%�Gl�q�JȠ3nCp&+��L����ف�Ά)@d��ac ǳ��\;�P^�����?@;�A�]��ޞ
 e�U�w�m�@��~E�c�mi�d��������)�V�'�,AtV�\��R�
�K�iz��O�ؤ#��e]J7������E�̿ �_��I��o��z̐˺��_m��2�ZL¼�o�ܕv�,�{�������)�S�Β;�I�FpS�X�!���i�iq��+Xm ���o#z�M�@2Ӄr���Zٸ^���A��m