// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:36 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
paKZllWDYRXmBAtoTLPaYv8s4At+gxy5qnwBB3Os+M9ntG90eyDhiIhpBbWwj3LS
cQIrmQFml0+WeVQMIlVl0mn4MJv0YV1ytel6dv4vAsC8p5uKcdyXF9rUHeeEexca
OQ6isKSJEN+26WyeJMq6iO2EDuVS2qmsGNBuFzk4my4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14928)
TpASaU4A5i3hrG16yXnkCxozrd4reAPN9hXgEOcs3jT+tTexOmCjHjOiZ/H+Ejua
qu2AWZAQ8oaWy/4YAPy1Ijr78kEWtdzQzrjffMp6WrWjtBHVoqWTxFFMxJRcs2Pq
mOK9dIkMrMNcrrWxQI1eoE2Mjmz42nB5ldni6IWHgN/A12wXeWpKAEjN1k+W6Wwv
xBZr/EH2KbjfFcIqs8J/FA87Onfj1u4ZRuaOVIk0goTExlVO0mgqLcD0T1NFTqed
AFx3HEQmVuJqQjC2pj2FUq2SvzBe+qtqDvI+39CqL8RHpZMujVoLsJfD3qCMT41F
4436N3AOkHTu7iM90Kr/VvsM1eQpkawp7KW0yZgAT7Ye+i6zcp4Z34cxgZH3mz4E
wwmjXBXMybGXwnFbDF2YSeyanNxtqY5Gw5bOBFCnilsisVyrgR2k3qJR8YJMpsrn
noJrHasQtalNKACVrQfIpOZbpJwy/KGXlfEwvrPtwm93XGKNh9vx2BTcZFzrgWK9
+vCThQKzrUkJQa0ba9Ykl8GU284++tWiffN+5PRK3C1XH/DfOZbtU2u8GfE4/E9v
gE2OW424Cjq/xgB2qjZH3Z3lAF7mBi70iuzoAGAaOr3c4dcwZCqsjNpS/R+3SHYd
R+N4qgGwJFT5IBnJST7vhPxYf34ZZqFxsU/Ho8QfPidfiiSUmPS+wSHJVvTq71a+
5S0r7TEn2OrNoATcc9K2YmSmRZbZqLe4FpyvCN7c/wtJ7IOUf9gETHKG5lqw4BPO
iFhYP05D8SllT41BDzuplpTJ58fFvsWRKq4j+NsfE9ucGzHdxLk7uvlFsHNMwujO
CMNERENgptShZ9EUYxn+BxJ+eI6D6uDlqKCgVoqetvZ1QTOYMmweudc0FxkUbPFr
zSVNDySkPYQVnPSR9GmwGjefkY84mOGgPd5DLBWIyrmjocja12a7Z6vMIUaZSkrc
2n7n97kNN4m/y9trejvuwolA+iVbo1pxhPfq9sqDzTChFVylfB+Qv7/636+zwMRE
v0rSYC8r8qjknzN2mKZz/w0v+Zy8E+tl4zF9Ckdw8LUG8dENcyVDYgjOR1UJrBkE
ne2LXlVdJeXqSPF1NQ72ql94Z7QR1lCYih92oKluc5mS15cUxwnDW9v13wxjcKJ6
yRvYh9Fx11Fh5T070NWyMfTTfYwEDV+Me9kHsxdicYVPwjlnedNyH2nAT+s9Sx9U
8/ITBrNwm6LKOK4YcuL8Gr9icGig3QCNodJpRfdD2s/ZLdJlZsaNPGiWOVByyawU
CCmI+KGStyilYdme5tz4yj0W4UzEB80KB7IvewaU8WFrs0PAnAP+v258EYUbgQ5n
xcHjFyCHaEvh9YBH0WHZd6VqtMgoZ87UXsYH5BCR7sbQUMnGNYW6DHxwU0Qqr7SW
4ArIzpPXe4oKq532DCMfngm8d2LlJxbvvbYNaL2Rih1e4amrbDzTuv+W2ZQ4Foj6
2n2SHmVSxXl+vdbHM56k3FB+zXhIk8OZqGvqMdFwASP9+D6nWrC1K9/bDz4uhuDT
XnQmmqwjGefGAEQWSwH0nlnKE87KnUD842Ph5Hy9TVlVN2LugsXETwCHOKkEGmqx
GcKASMiVJeu1yvbOfKpDQ7S3W1IJLgihigsJdwIG5mkZ/A3im7yATwcnRzZaJBvE
sLVx1D5XQtVYd07BuQt4CfyaJI1d20VhfCIx3eDB9qztDAnhOF93TVlkZ+fMNNIM
iduWy8TK4nwsolkEg5pivwfNL2t+kNFDimqH//k1POM1RRAE0vZlCh4yQaQBXpBt
b1DU52Q7zW1XWIIw9sceUZn2x66RWkbVduIkuKFOFP/84G2vjSGh1fh71uJR+0ga
AjyAzZRe3/CloJwJKpfwORGvsSCAhA2O2Y0jlfJpSvjLMOLlikv4CDNSOJI+K9Nw
q7vjyYGfqdLAjrUYUjQvI0BrVSCGY4y0WNvDhmUDcxE5euYuQQ5+I/qyFH0rWc5j
z7c7GAJgBMP8d6cMkAbPkBV4+9J0Alvnjxo9PInEDeHXbDHvY8pLAXMiY+WlfwuJ
9s5v5WlAlcG9phvTJDJHUb286d5pafnQIWggK2ChCtV8/geuZW1jxVC9HBFd1AQQ
FIlX3tF/ONOZWd0IBzx3txiDk9SjPKz2XPSTqOzAtraq1/XZfIyhhuSAZZqR8+TY
AN18mzyv/43YkNbz2S6yH3NLJ9GJEg//UawyIOpuic/iLMirmT4C7n7wOlW0S+IU
lnBHw1LBuVMiMoPVfLRLAMd6ETVR6Vn/OswPalB9e1sHMH1sG1lTFIgylbR9pGJO
D6IlI+f0izLba0Nxai9ewxTizzASW5KUvTmGCCKIunLP8qgo0+p9EKL1Pd4J/Kae
OvY+cIPWjC3RE0w//q23IgfkRtFyYMNHilNFDEJx+fnWiIuHlyRNlXAkokEf6axC
z2Rb7BtX5TgTCpEmhUUdu28b5XpaL4HYErg9itYEJaXBmm77DXmHwB3vg2xmHDR6
CpzIC3s1Oi8Npvlr7gHE+Nd5oiY00O0b8XMrfNwZSFSs46Lc5epixLRMcYgqrXuw
A5Uf+JDFzcMRy1I7tGOAF6sM6xqxR5IHOb/20PG7Ha8jlajVmMoFFopsbYvOvGAH
4qUY4D6UiLioU2FM0Q7D6gR/Sh/uYyY1pPPtPkZg2dTJI3yeb0pcycGnsyWNZB0Q
bC2d69Bn/H53EZGNH8fMmS7dBRGlLqKMYH7A5bcVnh8H6QYK2cBxlA19QU35UPf4
awMZlWYNAg3HOcFwaRqyyekYe1H7ZLstY/FqvIfmhAtmR4U+euPottOj8qU1Q853
8rg5Xu9DQXqFhmICy3MiSZryT5GfpEA6JW0kwZG0159MAv9CLm9Ejh5BqCMoyj87
2R7bWPuK/hemtWfe7F4vH71rVgAlUervCboUT34RmGoDTlDeXeF5b0YyxzFNgozp
BiuFTJjaeP7SGE8+8rA9Jvqp8kuR9nguECsXVoL8+/gj4F7Ilo/2vICISi35I2J3
XM1cmiXkzILjXQfhlRR7SV2ZPzpmEnNhPPS+GbXJ3kRKfWUeEcXOj+Krf6pAg+w8
G4j0uTW9gJKFjDlRGEDhb4x5vhkhgxjKgJp/JmxrXlcnzxG8WTJxhfZwjt7z83ln
ruLiAoK/9v1UHmRlJLvYFeJhWC1KArZJsa+3x2pMCDCAZyiI8cojfN0Uhig0vPFL
KKNZf6yyTyLZWKXMO5y1bjcB0qx+G1Me3Cz6BBOGaCLcRQ/dshugsaCyvnpchVrZ
Oasx0qWVfBVo+7BEkBldIYuriaA66EPpuZzAzTcTaUxUw+RBxOdpQUM+YY7ON2zX
SIx2bIwKHqfIy3N4dMvogu/9O9kRP/agEOl+CC/tTVqdiyhPVpQWhsHPqAGCBL3V
pbWRMcegub4q+JvBdGpQ7l4NLiwLM644OBqE5L4kFXZMPmmindg6n0QaIXF7sm+8
SJ1q/RUkguEW+M3QSqO4/gqG7qeUFgyIu0MKIvEmI59QS9jYVm6KBJ2mYtTqlF9v
tQiE+8XUoBxxUpiSJOc+RnY3aj5dwSUTUFU03gas6VOpHu8rhq9PGBWF3aoQ9eyb
FJWz5M3HqBaeaZd0aBtExDtizwnWiHQsuOm3++SKh9UQcBP3qxYGsARINw0BV+/d
VMW2MJycfx0jA51lnxmKbDhWAVkufgLdLGkod7zQaXtdVZZmyxN42g5mUbnnQCHe
1oU3H2rvEnxFXxXcZrCsP7/nd4DiQ3rsXOQ0yNrLtu/9FQLwk24QwDqyZnjPuSqj
DHJWtfQ1YvQ8cpTB6dIIwXkCv0KhRxZfMg5yl91e1hq04bwWHBIwEhiRPD1LfSdx
IojgucBuUwO8e5rnOkM1c3y6R5y3wPvxARSTHX6oOCAdEtxezoUivVrSk0+Ewa/2
GGA/ufhUtG1Tx7Lb/EBzUru6rCASTSG9wXLfmEhxDncd0zzRMO9dh6k5Yak4x7L7
GgXUwwChZyHHr8dIKhvdOuprtt0CsgSBLzK32ZEL8PMScGS40uwIvpxpVqNm5kOO
5rC5lWeiTRC24PWTpTiQqH5dZ/KVp62IDdvhQeTqPm9f4lUUhBbELA70LUziTaNd
B2JUZJ8DECa6+9JhhsInog+d7R5dmHfUOHSA/UiHTT7JyNj81SZzrg5GCCImBHar
QiYn1UwxWo85biWRnVYxHFqAnitp4y/0tNF7XybdhoXxarxvqJv+kw0+nop4ViW5
mb9SWzcyNN1ltjDJrbmyUBWqLeywTL+NApNmzo8RyVtniK8+VHqA8or82plswD3E
gGs+6kkAfPOLjf4/W48fnsney6NZMl5/1x2hCiL6e4mFHMg9xSOgcSLjbkFtjJe7
gf+XzB/Ktzkl0Qr78iB+fc0WNOzrz9WfkZQ7rOIP11MnIRf0jN4Q94l//BRM4o7t
xJ8ygaVZvHaN66zQf+9xur2iL/QcCYlife1Zua4XQUwhMC9becUM8ENOaF9obg5/
lsaSuL8MBs57kN2xRs1t//pPd1wgSxP9NNZLwODiGRd6j+Kwh3Wq1aBgemaMYnuv
YFdd5gpG+0xXDkHDvS3U8i2Bs20Mjeq3T5X1saWw/kt7pPX/ukzve8p+8/oo45jU
7n/zGVO0q5xFd3A7DVlp/SUDaWFYN8JeqE8LUKur2vb7VBn2UwzEnPbF2+4ulzx1
8MfUwnOsXAZ+aW7JuwU+TXvUDJyYMx4QGubEqaHNHZ/6GxBcKRqais3y2KfazO3A
pIqMCidfoCj25A4SeB1AlHyQXBtH/AeFYU2W9k5b/SwwoaZaDP0CHjfU2ogcOK4Z
QcreVs7Vlwi4Z0fXP0gRJyzsVqyBHPRk2pfZeKmPjmAKfVzVvTPX37ERmLzzGZN4
m17dgftfidY+ttAPhxs732jqphxo6pR6uIkShOCZn6XtX5/Xycv5/pLEBw5AI3V4
+R0ox1il4gnen05NXFICwnSjFawZ8DGzmtMGFK5ViDwkgMQNz0TWmP7niKIqQIVz
uRpbVBxNOZUQOkrNHp3pQorTnu13r+p5KPYLb/Y72mv5S7T/qQrHE3ez7BfyGqsI
BdkbgTF3rCUAeRiluYJt9n4j2hr2vKHNFp0wFdqtV7cHPpk3VJ9kITICdcbdkng2
9Wi/E5WOln4RViglJMnNMOew7qEpArFuJpmHN+KiJ2nukGo6780Et5F+f0RCXD2/
JTDEqUccu3ln6PnbRwUwVaGyb/zcRIjtWfZe0Zh/UJID+TRzhkm2pucBq+VKavZK
yRMDZnExQQZbw5r2nokmRUK4vyNh5/w9ROh+TyPw/OhZt/ThIarFaBDbSlgnA31n
s49qM+Gm6BLn6o3J5I4QKHQVm1DxSyjMWRhaj97E9pTo0ces8F1eqAw9dE976N+Y
U6mtxNKqWrhFYxzh4XaqjhJ11EjlVeONkAzOHBmueJ83xM7UwV81t97I3fMI8zeD
Zp4a+MXKupYUhjlLZp09ONsI4yDQoe4QMR9UrWC7QK1rwswJVm2ujJoS/N9lmOoI
aFGqoDekDIjzuJAZjnL/pV30DWrqbw3sMwQOwmKONjgk6Yq4EBlwsLkE6XbjR0+T
hjMo+F+mGrm77qZ7iz+HgumiI/QIyTnWDZByTYjCaTkqmujKq/LGrn3/iOGpUXjb
vRgoWV/6F8bSlHfRnIVi7h9QgxDArSSpUYK9q7tIcveKNWPTpeZcPNV9jhw/CmBY
krNL7ESKS8ezq4rtC0cYy20xRP5yBJQ7WctfqsxFnWw/lD58aNZ9ZC6f6tGrx+KN
BAxkCxkmB+h5U5SmaSmzk6V1KzpPxaDbOmHd5PyU+i3/mqGfGVemDW5H2BBs+JR0
gc3JsixMDWWCx+1QkF+pvEu/k9cevqk80Jb63E0r6+vb6g0Mct1PZLY6kE4j0coN
eqUbB1+A88R2SQANZZHJphuBhByLIYgXFAeaO7T4pY9e6k8NdKvgFNap5JCtqwkv
7MjfYKqkD4xiMC3yBzf99Y4MW8zFER1HVNoZMzpt4RIp+QqdMM3O1gFG2Rf3qNfD
GFZ8j5L3vUlbUA3tIKibJfUgnpXa09p46TVlRqQHQ+W8wbEYQh4dnyxCk9bHHDBr
cHkt8oG0AOR/r0Osczf2tLu0sLNnCUN7Okgy/GBIux1rzreU9P5njkVoLAIY6+gG
94ti73kk09s/iBZ95ND7XfujWai3Hsmwx8OsCgZl1NOAVv3s6cR3pjFhW9c9kEIO
lWhi8Ntkr1mDK5Gblj7X7gGKSkVzw/DoQ8hO9k+WsF2HPQlftYiIHHedveWdSOzc
CFiCTRKKdLU1IChPrP2Jh2c0Dh5X44XX9ZSQcjRkNlXaNTTrKziCkwSW05tT2wGy
OUkysdM8E/nVaC2oaZoTdlYl/kJodAwO1Xzf14bu9zp1ta5+1JXEfJrImwvYTMbG
oYNfNuXE35fpGoTUTCMGvb1YwfSohx7KnytoB4+uR8CDvB55bXW3XMBegpuy05ZH
GViQ/8Dky5NQjue9W2CmIpLWVJ4W2JTK1XKGdySGhsN+zGaR0U+DMDgmWh/M+1LI
Pgo51qh3SOcykQGsbhBg4XGR/yeKgC4rCT4TN6c+c4oqO96jB1SGSPY+7N0XERj0
+WBkoU77Y7pzc7zMQI17gLQenhzZLQI+WijrFagOzBiK65HaL6cxc7iB7u2oHZKH
e5jW9IyzULdDcKWhhPbcf/ypHVfiQ1vpkD9WnXQ1DIX1xfJgOWhwiMmH3YYaby9E
MeSmyWFM4u5VElakm0DxBTYQBtARYgFVI7jB5+6AD0cxrxYIlXJAdwpsplQPNoaV
dpu5e5lK4Cs87gGhBON5iAXak+GuVBaz+rl4lkqPgGNJm5/3aSziyZMQeZko62Cd
dWhgktUEyy2xObIwD1tNaANDQ74kBMMTvf0O3J8WsfFiD8GrjlEdB14sxJYHmTuh
scPLvOkhpfi3BFBuOsBK9pf3gCZKgkKIfFZd9s2wC/vWulJVllNd8nTDk42WI05h
l1qcktXaCPl9MQ5/Kv8maVEVTP+y02WFf5GyfSVFWzN38V0ULBM0QKUuZceqTWug
FVt1lkOCBMdc51WEIcH0haFEouYNdN/WfqyLEyD5lj3sgbyyY5es7eTiAqdIcV8U
VtzOMeQQTB21eQOnsVl4qX1NHbGuWk9QZDvnsO4F0IecadgRC0G5avdUIo96ZsTy
bNi8VbY33SfDGeJEcaXJvzTdDpI4bK9i6zFqiQaTUi+GgJ+tndwQ6w+Hx/229PMH
53rnKpx7Pa7mY9TBXwGC5Wy93nDMAl09Rl6AIM5PxoLFUC3xQlZ2/rC7NU9Uec/9
ndu1MZfE1jmT6sJxviKsZnxIBosOidJM5/qbzIGV+I5qkuP6Mba88udfDszVm/91
zCylQyLcXVLjJLg3G1sPmhxaSAlvj2me889LBXOQq0KlMehdpUUEngt2S4yHOCcW
XjoNFth0Hqa1SX4PYgCxxEYy+jrAiPX8zHEX2VS+JdH0vmT0tsL8hF4w7acjjSs3
bJ1OY6mJSM8IY2RlZZEIiCwD7xJ2uIcc65F94MNzmh2b0j8w7dS298lWWSrDkjmG
il4mLa6zXgsplLbKdS67C3f5x/mXujCeKTDs7lJTTKCHwbURcpSi7/gv0JTyYEJo
2rSeCHigkmHJ2qFOaFRFtls07KDkHvNwYlPGngkgzeQXB5ealLzHiA6bAFhPkuSx
zk++6eDn2fBymU6HjCEg0dSs//zSLR58pGHqTlE72j0+ySkGJpi3AsJG17KOSWME
aIWbHguSXR2IpybVUaG3gRv6v1B9i8MNuOJDI7HPGXK1s/xzxFQNHLJWrrxZlPlQ
GHwL7J5nAiBub+k7/fcKhV3iilfHitiSldNj4DDPx9jLRxoAZwDe1m5+rvsXzPhn
LllQk5+1g6PUSw1wrixOpRtoa9YGUOWkrVf6hDnnW7VdVlpC15KVbDkhxskf48XO
e8tylZ0JcIJAnQi0JPwD+or59561OrhmfwPT3OufJJTbDow9H8GKGtfY8uW0lnIb
nDS5LQmeBKbKxX1RPyHwK3wWo3CZDlkTi9/4s4PPiOSK293v7RPAnU17T/xFxkd7
rDk1WRAUN9qfrzswdgXQMe3151m6cGhTJ2huy8kmgB4FR5lbUuxU8YPVnpQWCBA0
7/B+WSx3ffq3ylmmiYc6LUgxjFPQyoT+MGfC95Tgm/XSePAOviXO886wD/lrIAXp
iPgbj5V/z8UJ/bdnWcOQCF9qv1OlBBSuI5qaLRv78etlJbjU7PWz3BcLnNKw5wzI
xZb6bsJLuFJZTw4z1Ji7mrVfeoS54VxnyhnOoDVhx8HiakaOnwnNO9tm/vay9eAu
51v8XkpFkKjG00m0KY5AP0atEwt/x2igyGmllfTnhigbjYyiPhIEat3s4m96uLtq
2WC8YWkuEXietO+8S84EpB/DgKCYdkg08hTGNnq5ftHxrn6XejdKOulYR8QSkcNg
MdZymQiM9AC2W7Ph+M0D7GmF41EOtYyd8J/91gIqVGA7YPdjuKJ26sCctyIiReJC
ZF5+Djvw54Nt/cwOnSNcgdq5zvpx8rq3eEOWL4xNnowwBB77zT4WNrF/y4I1IN+r
9dRJ42MgBqbCGDwvs4uDa7z236ziWwAjoWyOZBeipJhsRfWe1tRey9T2RiM4EuEl
YgCFx23URalUakEMjLz3JMjY7L/lrpHrcf4XgqMgAiVlcZJTw9BPRFocQAHzxDlZ
kwFNcfT93Mhc+HdN/kKhO6haBnHU1bs+ExQg4Jg+5ZF08LfSYs1uWUI1fZN/i+9f
5dvjB7AqtoaaTUJnT8HBZ0fBROronWdopm/r+YpMqHhbjgZ/oAOUr7uxYSlu7xlv
e7PZ5AZ1qyW029pSMC2T0dz58HU3egrzCd3PMKY7f0EjqxJbuv0uzLULX7smhbmw
5CYYzFluwtFiIlEsXh5gFbzUq5ODggVcZpbu4nXXvq5/TAAOuN0lfsY9XvUXM0sm
oO0MQTIsh4qyo5lOhsY62QGA6FAUlWsIhMzAeZDRzGI0EInIsSwPKj2LuXwsjx/d
6YD/C+lj9SYvR94vyN5p+Mj6azyB20hZ+uDXY8Z07FzhCIBp7HceGOYnaGiSPtJ6
zWU7eEcNPZIy6tJCfQ4eh98hyC16jNWD2AN/1O4iQY/Dte+L7OCogG4xo8mONDMO
NtU9EB2xyfyFGjY/awz+smjg+hTHJHckIEg471a5vMZMuQyG3lX84Wwzrb0pnDvH
AuFOzAoSvBOGtxwcTSpNp2/6si6hpKvhTNdWwWHXNwltDJSVPRPJpu8QE8LVAP1U
CX1N+8ywLWqJR7SCH08OlCqCtvABvb9D3OgQp+xR4SKY+2BQUAsNJ6qAKaxLuDdH
2lteClHKwFeKF+cl68W8f6gRkGBVIKTisNMw6XvMEWYGDZsXsyVYD2Ieb+qDk6IN
bU6G5/KzQ68armOUrIVPEwHso7b8J+RRXfKLporFnQTAuIebdP5GBrqYW99HulBi
vbax18qICLcjQTst7ecmXSfnt1T/ujnB5oBqCyt7s1beFk1Zu5l8ls960SloJIfZ
7FG+CU9XbOmpg8X65hhyag4gT4lGbCTs8mNyit5rV6F0NoUgDveXWw3qNYvMdfWe
L56npPrvOA5T8dxL1/03aRuwj8vUWgc3RIYbfS3WbGSWFhfzEwVSEtIzQruHiQmy
cDASUDGdpLqZ2ZfIELShlBfDu3b9+lTyRBi0a39JPPvi2RfegVsHq7Q8aZHgCQlt
OnuV3vfK8fpO1AVJ688iEhhtUnqQb2ulTidfN+meJ4iu7macK7VgYMVC9K3Ag+C8
T9ySYVarhn0xTU7tE+UK0zMm4C63diEYTMCWZ92p2dYjsvGiWD0J63xRzb9uJSGG
9OT4MVJm1MXu/v3G+SCF8qyZvsEmA7gDGXni0QpYrBZpfyrfr00JveAR856UqZGm
kAWk0hhP4kWVJjPGf6i/W2etwmqtWheOixE++Kmi9DBDPc/0EhlRMRKGWi4Qu1He
IbsyJd0D/eAxieKXJCu0Sbs4BR2DoQP0KErHarJinxZNK9PCMb6egYvxOwpE9gny
XS1qAuPwSWO8XnmfLmNTmqzvuO67pqX/5JsQm0kax8BYCobRFhn2gnwX3C2cM/dt
Zf5VVnmHz2Qb1m3QKwm7c9wD3HUEjI8P78wLl0uJeKVySrVgsMCwxA0JKG0nog9E
x9Hw2HYBTYZuqTmselFhCX8dYJ+EfwoE2dVU+9Ac1pu7LDMfVT2IiHKC6Qo2L2Z/
IZXQ+nvGa2247dbTiSnU67wwUQDei+gM5QYejnw5WScmMf8/Znz3L6HAg7pGHuyq
8JQ3+YdWDlPR8XOnz5WHoaQBr+/1L04F+4RW5rKQBrsRl6fKdOG+XLvkw1rj8PKd
hRERcq74SG2ZMGaq/Vxc8yMIq7WW/aqIJRh3LvoGqVlitu4sg5cPztU3fK7czIHz
UEoV3tDkZe/Og7lPHbiwb7ZYY+TjdK7EjiNIVgnqwgDBJK6SXo1Noa0/wbl/C8cK
cbBscOMcKhfbuZCJDvMwgocJrh7oHzCgYJWcHlWjd9uMWU5bKzgAZuOsl2PCZdlX
gPwLVUvCrKBc9FFdYNHwYIRCL+paiAOm8kCSVZWpdTjkqJpb6J4cWSoNH/+yHn89
L3AAGyW6w25prrSXUlJRY28PJS4+TXgouRvpDJL/tL4ePGl0RI9A/2HrRgvbER8F
87ws+gBH+UiQez4zTT1CPZ1RnF35TRJaAGZH1Zb15EdPuhCm1EY1vlLrjOoXymV8
RX9FzOkG5eD7Q2aYRv1dDCZ3e4B9AlWnKRdLEu2qIn+hafADxWJOvY8b4y+XxDrA
Fl/m4QlaP0lAFFHevlJJTvijQrpX93zVz9GCcXX745B/jxt411pt0eR22oeJo3U3
7Octxqgf6xwXqMBhiC+i2kMtouUattaG208d5JsqTOgj4cR4EldELXtuV9MbYbd1
BK1JF1XEF/NsEJSZ40mdMXts6gLcnqm7kG9VNPiOSkn+rmMyNq8jYwb+0Rk0Y7Az
zbdhSz02AiLm8DkIzEUofFa9TOCsN6xm5E2yRRofP295wi50zTwEcf1TsM6p3SXw
6j+20OybcdnZH4OeeUfYux3kUZIS5FqJtvpQKtgg6Qij1aM6n8JKO5/K4eE6+dtb
ZbVCxLBSM4XdjDuEL2ZkUFVc3JjjUXXvpTQ/kTk8gALfAYy1ddVrL0ThVw5hW/NG
wPPGdB4RvyR1T2G/YJZ+TgyHqMGMkYDSZM1a804WSkCC5w3ChiMFWI7XLLpLaXPY
MEKL10j0j8huIRmURSW2/3nxGeoqsLbjp47F8t9MoGFDZ0lHFol6Cisfy+4xUCOd
62Hy6zqNOzSbeoXSfSalvFpLKQ4kzDiHQWg8fBufU+2XRk1cKAw7qdFEXuPUjQ1n
cGwpar1TVwXOeB/0ujCKo/8OJifZZHSGO9TYjvytLMYhIeP9NPBbu5r6T65Tq0bI
H37JhlgjMBoKPVl77ZWaUtCNiEwp+1GiX3UTUAv9Gh7TVJfxrG9hoKfEhzCp0K+E
Qc7LMd8zOz/SmsxZEKs9QZptMtYIlmUQKzhjNFJnnV6V4pNuHHQWd2TVXf8vfrdY
F2pdcYk12e4HaavQ6NhRmpiozDcsEtpUIoJggp0AyH8zi5JhMVkcngYMjRNszfD1
FZdshinwS74KxUklGjDHjqaFE2WGdEaVA5qYHzB4BIgpZWGZMAZrT5epJIoRdvjF
kwj+QKYrL+hKKxRM023OS+vwN+zRlWj8eo39C9KtVXI8ia0lmAxk7CQSWBgatnpo
ADm0o/l2lFaM3Rm9mR0aNbbajqAAYulS+5mPSMIVL5thBWRbAUmXp5xqaF6uRLtx
cyAksvJz15mkSc+L9Tja76K7QLsssFAjFiqA/2sdKM1oVjCoAcb/AyGNSbbBZA1x
n45UrzQ8YAN2ltDUG/nWYfO06tf8LIhNqXpCyXrwOLQIRWPbK2NizOVhqIe2D8dg
TbloocIQ/e7L4n2JILFaauOJN6wXfKj4nTU1quWMWcuvKMzP+TyctZI4z80MuV/E
XF7HAiNu6Obgc/bJ9UU7VQbDmLM3sgClrRtkDNk8eEluhvI3jMuHsVzxYwp4ADqz
/qG9Hlb+Fe/hZNJRPF7sP5qrvXiXUCAivnm//DtA0Vy41tuzaYq+TBg5TANtKlqv
3MnDpZRMtrGrgR8nAl6izggBEdbdEC2mqsPxuJXP6f7n/OsyVL9UZtyi5wATGyFz
/AQThZIlA/soy+yIZs1u/ipwtbNXasegQ5RkPskkGxCcAbeMqQybLyVi3SVHjWc8
fv2fBd2DFYoAkEtrCV/PXhuhGMQMVl3N8IRZcK7UbPzVi3+D14VpTK7uj1sbPB74
IeVGbVYCkQVVH0/L8tqDdZqnjCLz2j14/dQS/n49oIOVyAm3823FOPtWJ/EPql5F
7oyfQ14hFXRWzLgypd7uvj3NkxNZq0IGFT8UTpHwJLEZpdFRcqQI2p5Vaxg0lY61
RpEqoUhOoxW7PaT3RnrUABp8l577kYBRfE2cAponH8b7mBCRaZXr1Rq9i5qHuVF6
VPjks+R1Cl63SJuG0VqXKKqVciPTfyU1zWl7VncKsGW+T/J+Enktt5q0AzqXbQN7
5mW+hGJ2CILeK59Q+sfqaU3jexAvCGonVzivQh8Qs2GGyu592vGhrb35zA+XmJBP
s1kGojF1U83QwE1fk8mIR9X7wN+JLF2tG/S04UgxIoBrE05TWr3SlW3Ld1Mi0ASz
8fdL6ygxKk+YP2m1Ml90XQiOXShh4xV77EmD705O7HCiNxq06R3msMoF7I8/niC5
3/DLFy1o6qfOXuvUXjWqtgaxwoJX240EtiYA8A++cEDtQxOTrEEILo6aH4tELBiW
bRMcx9eOcz10UZxix+Df/KXy3Doow0VawBqJ7Z1h+4O9Q3NlqfWaSADJ8+7dnZN1
fckEaUnmhZmGs3mK1xjNHxxGjrIa///k/0Nig0Da0WBpvyxBW2VS40x+EpQaTksv
TFq7C1b0up4FNrmP6wVWF3fEf+/+BWgcCIUwXcQ7pw+MDjuWJETxzVKzo+ORr0o5
GmCNeCxkeqsbxttnm9AYXO9OWqwAFhlfsy9TF/pJQoFLMCCQSlt0iQOsfZPxn1XT
aFs6REKeVQ+DUDL07IpCn1+mhnLaswgZ08JqA9EVmUMO541qUEmNHrplGP2W2sd4
jQokRKraGbRhqUAnJws6SgGQzDuwVgSULvlgOIokj2DpdLDFlNwDoa2kIN7GMh5l
1vT0rMlQ1fCEbJ0xYlHOSa+QwKvkXsi9CLSqr7Rt7p2RWNL/8A+/EMk6KyVmfXzT
YbwwQ/GyM/2PVvHYcWxd4S/8X5KyYbHJNBmIYMUyvs8WnCWwPKprKU1/aeuzYLxV
WgSWf+zDZ5w3VW2CMKx2caokbgEsynyt/DYrHbKchyqe9IFkmbmuQr+Iimb6en/2
8NHiZ4XqNkGF98CA0nZDdGRZDsLBTFcrIz+3gFvFKIUyKtIIrbcdLq8zbXJZUea6
sVXFWyS4HfpJmM8X/1mPsXQU08BYVrVKWGGnXChm8ae10GqHoyALckgVgspuOlln
sJGOozSUFhBzQ2daoHi0KExwELTRJmSXFRg1AeKPUsHppxbuinuT7wq6QxVaFSi2
IeynsKeWkmnGq1cTJjPKuYWX2+WojqWa7zfPiP9ckDPnNVIZLyyTTFavvKbnWFfs
kihOBcDt+EvuHLe/EKQf6ZEmSZuR6S793mCrnsFR9xZ0HAICSvhdRTptE953Z0JW
VdkVmrx9LRcY4sX6fTrUn3+VwbQwea+kgcCsZQpAkEnFM+T/iHEj384N0DKXTkws
gC8wQyPDzjE7tZ0osLKEx7HWoUcSt0xanoBDLRiSXYwZeOGpwvAcvEQMjrE7mffL
nepwupUke8sddSNzLwPojC1y6hDU0KK0RIL4jmBn4B5I6uhhFAFHABftNcvS8Ycn
ChKmcLJlsCgHaUri2wJoN2vmDgMeKd4kcxZQlCzxeS0qBi9MPp85UmcR2pvG53FF
AaO8gAmRAEaw4PW7TGRkhmgnkYjreIZo0p1KO2Tn0oJiNXriIcC39qTMEFO/bF3V
CScqLjh7EYtbc8X5OPn9B/pENxa/b1lcOLYwgn3DaVXB9IvpIAIiz3ntsbLfscMu
pOOptLRb6rtd/Mq1+p9mQWSKcC9etFOsa62kZBX34e53PVJQaOfW/Bn+Q93dZ7NM
tulKz7psT4q8OfZrPTFgiFoo++cJQT64yXpECsTrSClyImWkBngVwQZf6piRU+bA
Hlun6fQUyGsRXEXVwGFaD/e24XdgJna7LMfn+Fq+NMfOX3BdbJ2JQG9ibTypwsOf
lxeBiMSIyGzD1WDqlJdsqCR5hDJEM9ShO/EN/UBkq2vf9vUtVnAT0PadB78Pe/yD
QN4bHnIqcTH4j37Dj8jCsJcbitD/Ncf8hHaw90TGHiBwbLwIdPmnndfEJRO4CNxP
sopdXZSINxUtOBFACHcCv+fJ2QcrIs2IOnQuBK/wPUKRSA/tZ1D08LuDoSUkQlk7
C9fDAEWVwrQ4gsxEJOjhHIewspy5bBtZKNJVzZbTQYRkBezqW3tG4bbiFDA6RR+Y
DqOJAU9EX5tYMLn3/zZNW5h3cZ+on2RHFlXL9ST2tGAc78V4oVoFH0cQdaF3uojr
D45ffTHnh2UxRtkWrZwzCRotPvCLf62wqqulicK+tjFt4iiRqU9g70EqOLsd4GKm
S1SRz93Oa5SYj93gdDfiII703FEVCaCB31R+GOiuWcUJFKVOeWDwQ9hL9R2qTi9e
71G/5YteVLrPYzMZbdgzCoIdkQhxf+sTnnpJHlrNb1fpiMFF7knQXqIHC5MwfkJM
p4V4vnJwa03IWrwk0wJlZXmizNILKT6VYKZ8L6gc7JpqrjRxquS6jihiBr+3yUJ3
WB7xfCgYVsd7Zo54m7/RCXfJ+eN7/Y+dK9L37FTSjZ52zpE/pRi34rxTHwOd6eB+
BvuxxLv7YJrhdDcrHtPncOCFkBo/0SHBPeOjSZp00vKgfEffA2mvwiW0rQ03ViLf
fyAnKOar9Eb4ZfEhj/c7aidvz/MEk3yHNowvjRjtOppFlGL/7vzy6tOzUE4GuwUH
kHYFTN4ruKNlxz/tMT0hHx7ktBfpHgq+G/i8lyF9zQxabslp5hzFmjhIxd/q0dPw
2WcjupYOgH84BtqT0Rj0uDH6qtItRwzw1VaU2+CpnnyOKzxg0qaoBJS5bS8tzTpE
xQbPbaK7kJz/vQ4/WFg4YD6PPoKYDbzTtweJB384rRjrItrOtDtgxHnogBiCxzqa
fBLfpfEZn/jQqjPMQ0B86ZGIXTZaFSfX7Tx6moEuwwXFECu8euGguDVnlFDbvdpk
uWU4/ZRTMjxNA6mu5tZVgf57wW0QiWm1VsYMPHJYfWlrznkq2jW6jweFr9KMXhDn
H3SOjI6BUnNPwkroNgqA2ocBHU2XMrAGVfsJMqzVS3Y+m78UqWWJrubVAOGu5ehD
whFak+q6q2rCzqOP3dWRaaY+m2nmXIXpO86MzB3necsgAfge2Z92p5Ehd4HMQyk6
NqLmpYEq8wndApJUY00iuxpWEGOoYklheYPW72xtMmY7yJGmIWKq16UWcW0MpAkM
i+MnLErl7LpMlR9kINYmpjpyHtJwKCkXRXFQrwGms90jVRjGRglpf+HPNNn2YoMJ
pxgjQTO8KZuaLH8AsnwRn4SIUxasOdaClPiNbB0KuXhO2XifNQJQ5gfmyv6wSFiv
UKwaYvNZLBdIDUF/1/5e14b/frJ8ZEdUkmfyenTLEcysE8CsPJRJAEAeNTv8vgoa
KhRkHC6vfuDr4MJe4U5InSB/sbhSV0WdNDuCrETIqqJfXO6Q7qoWKAvTqxWrkO0I
I9gB/TvJRLa5tKvH7hoa2Gf5eRKNoNCr51WXjP9adFzMeya2ZvmYQnsDsgLXMTCm
NSb27pBVy1HvN2RPgHTRYG3dflhTj2wI5/dT49bmzqmDjWqQqMHnclAiH453G8P1
rslk9DhM1Yqlj79dZG9V/pZNGO+gkccVRmv75GnSm6OSX6D00WvHRoNr00i8C+Xi
ok2Pd3Rib3ZwhINFuzV1qV6hUFxyTQyaMT1Be2HJfdtE9YG/xlztb322vVH8xLld
LBo2A5JCMby5WmLe5vpNZlogfBdBBljFSsj9G98aP+dsD5TzRA/rtGytwZw1QAgk
+lsqgpkLJ0z7r57MBMlmPzZi5uv+b5M0zIZthARgcJRLWcZ5gsOlyOSkEnfRotq7
cmsumIyl/Cqi7Dy/kXOGWQTjwgAElN1IaRmd720xZLXK/RIFBXT5nMZEgtjZRlGs
Ca/l26O7yWvklLfqxfTGuceOo81hIt9VrDmc1B1FsuJUwviAJusvvpbgfPkCCxMg
I0LMxASerUgcuaGjR5Cw38yjkclkN348vKX4AcMM9+QVUOhoCmWVIiTxT3XiqXDf
mH8NX0PabstUeQawSPbFkp/NLzMavXT5cxuxgwKDyy5+BvaV0mzTZezIE5VHpWvH
EVL1m4wLyzEfNFdwsN2EAFfaDX+aUgg6+IVxpmX+Zg91hZDLxVWoRQiSYJtSwQuA
C3Y59MVYbR1iE6MwkcjxIvGXcozNEyMbmz3wmzw/cg1LuoSMHfQZZoc0U3DIjJTB
oas/H7tAhgDaciQco1oWZkr0+4WzrTk6WSGDld5/cbUX5bMMmdku7MhNY9mIvCci
HD6tOM646T/mm32F8UKhcRNXkEA6b4BzgUZRfRyTRPcRNNUEGCLoxJGy1KAWWy0h
TjHbdjJqJSRdnSRdnVzfuoZAlgQ7eZZjZdY37fC+C18oRLhjGMPKTrNGitUWugdE
dlxvMLpNMOyjP+NqQJrM6E3SZnR4sOLZUPvgNOLVR1d3EVSwIhs5GcCOaIaLk8vv
s3PhWxdTIXCeZhRo8CzHAHMciLx91u/Yx87SN58O4MfBvB60GJOJ00mwEEStOizJ
zfE0cc0iISdNNCqnatFSr44uOic+m6fJ9WRbAuQmatS2PL/He0rXn6f4XhFCpGde
6nxXtR5v6Z+dp3OLdxBZ11ZH/l29yz6WaF8fzg8O10wARV75tBqlX/GUcOtC43XG
/RQ1SueLVgNj15tbgtsgl3LoOsPLIO8Ws7bE6oj/gVwMkf7CXmm7+Iq+TZuLS5zr
ceuYyOvUsRuFoFPT+wSuBFUITNGRSo0VQLdEAT25yz5wBaulmA9PjOThzIRmhPIm
aVDFZPWqdszURRvV4IMz39zB80TTf8v3DsnBJDxd81elv0YEQfjUwV0wfyzv4rl+
5WJezXGhU50cSLXuPgT4baz0vUZfMImXsJk8cEmKE/FQQjl0mQ1xq12hcOV4IF9h
EmtcpXadxwbIbgruwV5AagadfpkYo2yKMFiGjI4BvOOZ+DWTaailr8te++2QuZMT
P4JW2hDMivExwXE08qORvqeC1QBcmTlz5X/da66g2qWzYySfrfh6bCsRIr8R2Kes
OIDeYM71TJJE1fq+uweGYKzGgCnmdGDZs2Mt2BIpGm7F77cRYM8YZ3sRL1iR/WM+
8r36mbvJxH5BV7gea3GFStRXCe/gjAlUMBsN+jEGmN8mwzg8d9flTWhQFANw/KwN
IUVANIbqK0e8hs1CVUr0XItCskc5nkkuGvynj5OeZjnBeTscCjZ56+1EQ5Va1GYj
EF/naWtycsFty6Y8gH+mhw6w/o9xfJTgC4fAP4lkQRQZYSduGuctTqjuyUhv2gEC
UyCOgX29NfVedvlHzf+Dk+iCw5MqO+5BoTIY9fL9RUnbh1ScUBoQEs+5fBj4lEoK
RPuQo5IaWKVhzOovSo35agr0M6di6C/4ri4v47w9OFtQ+GoSCswLWc3PGe1V7p+x
X5qBpevsXy1THSnoD0rRfghdGx9MPqRG5AzOiwDhYcdpRn/RGtl6nKbBQ5hmW35a
at8/MgbLwO7I8CkokEx96XDnKzKP1wH4v0G1K/7hyuCPLdCsdp7k84j2Dg2mHF6l
JJnjjLrw8x4W/vWss49sMlPuUjKYvEAKuMrR8ohWwxa0In/rSo5q73hP1txnZEid
ed2Mh5AEFlJhJFtmySYQdmjG9imI/xiCq8IKFBh7T0m9xjPZrYYhRg9HX2H7ivqo
/Vi6SOIF5nhFQjF3sCBCdAEwE9sjgJXhzUlTSqq3h1v+ld46wLUM0GbE1f258NbM
AV0QJnjjLRjewbDUe4x8Wqs1U3SwcWJ9yHkJgoP9Q40Uf52MOgB46mzsq0gs4mq/
GETKXTUbLfReyKYNUvM3Hb+Sp04Ly1lVlr4+htWHuTk/xGNLwPLx1GzAPAsYDO36
TbpNAx45PN4DcaNaAOdXxdTiui3vyQ2rFKtPvWms/z1CePXMf0XVUmGwcdyX9Q6v
h9QwLjJBXY81l01f5S161yJxxqh4AWN9IJdVqhu43YREVHe4jgvWvkc2/M8jTcZh
cyVx9MmKGq/w6e3UIUkXscx4S99UOGt84Q7IMLBwOojCl5fvv871hs1wrhnJRyK2
Ss93BehqC0qYFrukqBHkKUs/pImtG3fZlscfQ5zreSczHgy6Jog4oZ3XNnZRJojd
lNJQnJWywchH1ZDWprPL9FhKSPlH9H2t/qAI9YzWfPNnGaB7lSWnP/v5XFtHGMzo
EY9IeJ+s95lYgcW8lfsdFPdnZpBFcZPadlwPbGy3sgjC+8IPzicPcVFpvHMRmtrM
bz2pGjAHOyJe1bnt/sSSsQbNu46m/L7xFmImNdjX84m6EyHdCmH5lFha84mPm2HM
cZKRdcRA2fdsrS5wdeSn6suA+NqpFono7Tb4YvH0OUmN2I8UMUGYhNO+HYKuqh5X
zsQHR7JPhtlRt3sXoy/Jn36Ggf5g+2+UXoiw9onqnSp8+XKzDJMD+/f05OvZOUjq
Vnrl84CWCXkkAmSHOX9fC2bQprIpKw4n+XRPkScPSbwCE+MOKVntXy/0yquQ80cM
tjc59Mn0aFeIbXDMCf+dGdXZ9WZs/UHrFpznL6yAJGsFuoV+hPo7qcYeyUCMSRRh
KNRTfYbT+FEzXDmv7ts1uGiFagnMuf0t9xBFK3oD5M4gOTcNeF+2Qc6NAVmcnZ7d
4yGSr6sBo62rmdjtXxxHua+2YNa5dXwUQCKp1rP7QBIeDynR5uW/FeVF8llcw2dH
g7eMEkZa8VwiHgsNB4xO4UMFmL7s0Qg8aWeq/7Zqz5MCX8CW/3EaYVcF8U8Y3eiA
zOA9abaDaft52Q4cBgqziTRoQGsafzeryQUBBPlfX6vWanjjBnSuaLuwGwEHDgIH
zMcedjWlbheXp92McPa9SfeXQQEgd4KbVf1mC2n3S3dYq+EeCzqiAx8kBpQEAXTU
GJBCMKKWrY0cGn8s4h5G+6gHcKjYtn5YDth1jyjeLa7BqNsrSx7iZwDz4RWplQwV
dfzr+CHRhol0B0RpMDRHUlRD7SkQihuuzXetnES5MEywrLcO1GTZGX+RTS/1+xxd
U8yVVfD4UOZhJ054qir3MWksl4GSofJIKyenP/RBL0qPlmRBo8Vy573Vtq2LD7fr
8LcwZiii4wnf/BjyGCANixERAHNEjyVksbiwcaAmUs1/z9TO0X3iXXhdV6lkwBoX
S4cMp6R0shDrxeXISYSQZ2tAoDB7F6iLln/rpAiKxW/ezO21wmlWPfbVUqGGfpTY
KoQ3AACt1OVKKb1efuUmDIS42JDxPpYCmFtBcI4XSClt27h1QNtqeYHd1TVFfrl2
8/ia8Agp21egD5uDTPe9cqphotvMbxIxTvvTnOm+XnOlaAn1skdNOIPracyBSe2B
Wmux1QxqB3f17SPIUu+HwzMM7qarxwg/LGoGvHosc12MqZFpopS+ENkbIVduP/fe
Lh7wpk+kplMGHL++SzhrTj5nwmXQ4gtR3SbB53VdORub2Fkjs9wsJnlWaUkaEwxE
`pragma protect end_protected
