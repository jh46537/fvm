��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�9zrv��^�t��|솟<���+Wz��ke�q;�"��������U9�:�	L��������27�u�Z>y۾�j �|W~��-܉�L!+�!X�%%�¹%[O��U��UA�^�n�v�)e��c���v��o6ٖFX�E��SN�M�8�SC�}� 8���8,M����{4
K���#�4�k}��#�.Qԟ��Ԧ�"�_6�>uo��2����~ �L3�b�q���g�~�G	�� N�l�<��}�|�XN7|� ��Y:%��(��6S!@~Q�UC��~�6�3�"!��v���,q�|��T���>\����-������@b���\�F jm�
z��?�����5�yBG�_t���h� ����1<��|8��v5��4*D�*͚�L�an?aYԦ��ؚhJq<ݜ|\u����r�6v9'v�����po��r	t�ʣJDU�A�����ȿ�p�D'�x�c�t�l��D'K-�F�[�gǈH`V��x�� Z-��uPu��Î�N�\~�@����y�L�!�|i{ &�+t~�ퟸJu܄�Y������0�WjC��cS�5:;��,�y�i�V��Җ6�i�@��$��>"�={�;��f)}$�r(psl1�w���8��5�x��q}(`���af=;� ��0_ѨڸV��u�N%�Z�^��2��.����Hċ��}��z��ԡ��e���������A]��!5�����D��K���m5��y [E��[�<��Z#y^�Ii����h�]O�S�%PR��"%Tg��K/�l�T&���:���B�8���ڟ��3i����o�o!.Yf�0 G�G4������Ws��wY�f�<�7��55�4R�:wБ�N��١Z�8WS%ɞ��D�~9P��[0>" dsPȗ���P�9hM�9��/I��L�����I��J������៙�8�;/����%j����Ɨ���i|e��UW���+�F>l1{ݷnl���te$޺wt\��A�*dg����y��3���L%+�.k�����3��vT���=,�ȖD�^�`z�_����i���1�dҁ���QU��q�4^U�-�UU�g�8'���oB���⮣Q���b	 ���^�s@��k�W\*�l�C���S[��=��SE��A>R��N�O��NZ�+�W t�0����rP�u�,=`O����T#�*b=���!!CTY�T�F}4�;i�$�z�]������l\i^`g���"z���e��o�DT7&��H�Q�1�V�i��'0�{�G�E'��"�)̞�3��ȃ�ݦ:t��j�njx�R'���)}��|F�打ЧL
�*�z�b�b��"�}a_AT�f�>�pC([?+����h��f �*	�U�7�D������7�f��ǟU�J򨧏7_�P	�"'�/����"��YH�ZP��$�:��|��cR� i���U�/0=���E�ot�/�;N�d�����(�C�K���/ܪOJ����������� Zį�c�A��~������Y]�l`�<��d�!x�����q���]�#a`dy�x�G�M��SSٳ�̡^u�xq#�5T��;j)ͬ����Hqv�蠛�6'Jލ���E�C�6�dc�0��q!#'e7*8߯�4�����G�AV���'_�])YzVt�jEV3"�p�ۼ�o���37���妤�Ni���`%W��峈ZB���$q�7�X�a�j�^)���7�0?���I�Ż��Pe<�lJ�}(�>�3��E��R�}]�9 Ǐ�(�Gz� c�)0���'Șan�9�El"������3����!y���U)���1���wu*+H>�2@I`3[/�@�.K6=�{�v�p�`�G�nX��d�l�T�-־��I�SH�m+�HT���{P@ݹ_���$�ow�����!D@$���k��]-+8�*;���Ysf�$ꇽ��뻇㎶�[ʳl�o����^�0;DR��<�dp���i[�_"�`��8p�����3�=-f�9������b�N�qjpeW@��Fxm����#�@��}��$鋟Z�~,�r��`K�Q��Mq�y�d�b�џSz���B���.)3��S���m��'��ABӮb��so�pS�nEx(��:���p���T��e�)�ຌ,l�&�j�������Yj������X{L�[�_�"#����z�vw �a�N��5զ��J
����b+՟�;�L�D�T����#��raa�x���e�e&�0#��E�h��Q&���*���^��{-/��h���%�(-��2���"nK����
i�j,3U3�t��=$��-�/�U�S���Ӳd��X��Ar���h"�)��M�q*en'HlvU~3�h	FM�1��E�G����h�8乪آ��e�=� ��6E�r�$�M����7'¢?0f?@�.��,� Z��?},i'������#����_���tfң1;q�Q�K�6��N�x�­�r�Xl�C����yX�a9P�(���4t"��5MBG�~c4v]+ط�p�pb
@��v=���=?�^��VL��Hv���tR�Y{.f��*�p>w0t�SPQ@2�� eQ-)`(S��_�A��[�QU}�
<��Ǥ��ajvQ5�ə�!�N��6��D���d9��t#KV���&F�
V\W�ºR��n���IXa�0V2�-�<@�5�g.���L��>Ƒi��.+��W�(���:�z��7<�x�n�����2����?�qP�D���z`��k�{��6�\3}3���[s�1J��E�o
J�YE�c�"]]�0$��<���A�����.�r�˄FI�Z�@��p�@�P��j5�@���u���VeH|'���1��Y9y���'�`�Y��1tF@h����O$؂�����YBO��|�C�Ԃ��oi�6:�#B
c�-�=-v�=o�^��#@�Ѕ�",&�-���kU��åoX�QHR����S����S�<崵(���$� 8n_�-sU�86��ths,�s�f$�;5!p?��4x-�V�Y��О����}�0�u���#�q�cf�,ĂD�(p�i��"�#F�ش�L������\��>�pl �Ax�Ӵz�K�d������T�H!�N������������̠<۴ڷLA��Db	��<]��d~
�b�c����H�煨���1��R�Ya�ۖל�^�
�+�Eqi�	s!�ʔp�Oز�������9�����⼚��	�R���t���\�� D2ABZ���8қUX���iD��M��U>�)�6��*|tg�Jdz��!�@,Ok��7�gt�8o����Q9�yg�K�疰K]��q�h�+��g�K%�+���/�$Ho&�m���$#(w�G�m�s�E�̦�����a��v��1�>��+@�K��0��~ud=�<���?���"�A�
��320���ߪu�y}�����²癞��g�	ʇ�mP���GOq�����=�Q�PQ�e���AjN&҃�	�櫔t��7�Y�u�R��w,1�F/ {[u#Ϋ�~W�?�!G�v���;#��|h�Ck��jk!�7���덀~�%�'l<_�a&�'�f�{g��N�qɭ�)�AF��yl��cw�.'}���9�c8C_��b�`�&����X�Sa�����e�c���kr�E��ܵ	c ������n�c��^�����Zx��z���O&X��6���'���I��c.�Zy�*��kB��u� �>C�Z����Qe����Չ�+I(0C�3����鏩]��L�w��f��0�D��_%���!�Ls���8ei�6-=%���E�����a��T4�Z>�9j�h�G��z"o�j[^W�&�C��^&b�x��⹺�y E�R�c���c�K�L�v �� �ү��;0R�^�9� 0��{xzl
�{K8+f�R�*�$^��8U"�nY��}��𰠄g�T�V�=�"~������E�m*+�a���+ЗGՐ�������Ei����9�2�c?7���m����7Fv�
}B�y�Y��(�n� 	4VyAz��W��ߑ�1��=g!.�ebn	+�{U<��ǚ>'��]�7u��?�אo�3	��.�G_�\�̌��S��/��]�������E��m#׊��5�!*C���4�Ԉ>����#�����Ѭ���P�uq���rR��7i6�p�Sa $�V�MiT��f����E�C%Ua$E�{'bΖR~��l;Ś����fx��O��*e61������e '^ʯ��e��b!X�~�_3��"Kg.�m�PR�Z����s,�V�
�(�@���/@O��T�P�b�f�ʒ�-��1jc��b��4�tE�]�ݩ���L�q^���mf�<��D$O�3*�_�S��m &�|��>uH.�g֧u��Ue,Z���R��=;7@z��>��8��W����zS|;�qG=��= �ߊ�E�O�`T%��T~o����S*�>�5B��@��n�m�z���ԚHm?�Mx�a��ȓv�5$EP���#U
;���{ɉ�[�p�|�U�-�J,VX��OJs�$�kM̪^�$���Gh������:�if��~�� ���9� �z7�	-�o���n1�����5�SWf7�|��mX��� �[k�|���l���c�deƄ������ �̽�̽�#������}�G*c�U�4�w���FR_w��ʼ)����;f��^����jk��˾f���h��J'1Y3mn����	�컴���L�^��37-�^�R}Nȣ��H���amh�aԩx%���^�R�i�~�k�&=���6��-��p��(aX�Xk�L��Ǒ��l��Z�zC��l+[9Xa�H�bqA�X��o!�6۶Om'7=H�ӌ�B��C�f�k0VAV�v �oy�f�߶k�K#t{εW0��9��h���T���H�R?�?����c���hI���s)ܞ�ؘ<���L
o*�c[�� T���%������t��W���=`e57��:�����hw*�P�j{�T!�{���v��`���K����3-�� ?`��p�Էe�"�p��\l�l��Ti�0`��6(w�n�D;*sͬw�2ԧ�b$�`�e�M���4�L�pY�����?/���-�hM9pN���x5�@�@�M3�!o�*ꙸ�6��*�T'bt4l�&��.�M�B��9o���Z�E��$�$�?��/���!��r|>3�h�>l�)9/�M�W���vI[.��5��'�kȱ�c�o�c���.���U�NO.!FZ�9��&���|��hj]��tJǊ�v��r��/��,À:I�E ����BF��~��V�% "wv���g�w���0��=�/)��â~G�~T,Ai���w�,���A[��d��!i{Z;)�������vSO6�w�wPã��G�������mm�kW�r�8�ڟ���L /$(^+�+�)�cs=����#���BMw�X}������Sc��y�ī�y::��^3�|�[�giLrX2��I�kOxЎ���*���}� ��z�w;�����fכ�����d��b�Bu�c�H2�,%����ݒ��fk��)<	�ៈ �p��&���g^Pك5�N�{z��W�u!њ�ז�Bk'��*�4e��/Z��\��eP�B^�8M�h٤8ly��K�ꑘ�x�B��`V�o��Xj�4�Jвq�U���ʞB&�AĶ�)"�;���P�W׹�r�6���s���S�X��}4%8U����n�D��,TH��6O���uÃ�U�ލ�	$Gq�:1@�HX*	k5
���:�2�'aDެ-�Ae��W�|�*.j���^��V�@�P��}���S)cL�U��-���Ց�YV%�6�@����l�\b��|�鼤NA�Ɨ.p�S8����>Z�|h��[J�5l]�:1�BX��[7]�{c ��_�F;lE֍x���y�ٕ.!)Յ)��ѡ�<M`Y)��'�i�E ]D c�p=54	���ß)`/B�7^�6����D^�޴�!�-���N%8��D��Z[٢_%�]�*!7"y��
�j�[��N�Vf�G-y�_Hm�9o�Z�e�{��2��[�z���~Ą�
���*�II��UKG�:�P9 n��#�Q��8��/5u)h�O�}`pW�8=��g�/'mR��-'WdS6=E�\�MP�B��m�l�������䩾��Z�T�@E:s�}�\�7�J	e���,m)Ն-�G �Qz���p���χh�}rd�I�F1A�M W]���M��I�54v�f�G� ���K��s���NAƨ�i6����k�riDF��2�lA;%�{�?X�Pj��d��Q�7�"&NĔ3����xN�Ւ�ٻDx��\�_U��h��HR*�S-U�����ՊG-��'�nw�(�ڱ�M��.�h굇�ʩ��7��E>i�<Q���K�?�ҡh��T�m���A����5Gy=�'7*��]���e3z��!�vѶ�X[�(d��*.R­	�����=�k��x�DPo%�q�*��`XS�z��a�!�ο˽�[��׸KL�nGli}1"���{�z�%�ˊB'R��r��s��hJh���U9f���;��D_�y��`bV9#�����������ڷFJ���E�77�.1��,=�r�˥���d������;�w�o���.�O����)D�Ȣ��+F�����$9�Fk�#� ��KGɱY�k��"j����Sn��p�>�G/h;�Q[7='���^���3!(�@�d�,x$�:��,j[V�)^�B�HI����!Jo擛s`�j|
��}W��ӛw�s�l�82*�x���^O*���@B��^��	�A���2eS"r?�y�1��h1}��S+.斎0ȣF���Q�q0�h>@��mz��I�O��i���8�ӱ�Z,�-P�0�ϓ����ʹ?!ݐp�
VA(VjY�������g��+	ϧ�W���b!�Ke���h��ɐ�Ƅ�0�vmJ�QG��~�"G�ֵ���?���}J�`�t����h�I��8�f�t?���6#pB��YYao:�s�F��i�Nw��zTO=}5
,_���8�^�1�gg��YnCb�ܼ�!j���x�k2q��.�.q7:�`
�(��m��*a�j_/����-(�C�=�Nͮ��b�u_Rd�pc�<_�m|�����d{�u9�����*l�vd�-nRU������� w׳1�"�k���X7�Rb�xrA�>y�c��jش�7
������ōFs�ô���&��t���T�〥��р��yx+�^�6���0@Az�>/�:����j,�
�Bu1<J��h�D�E'�A���m�`;	˷�W¤\w=�y+�{��mQa$��\�Q�ʜ"U����eWe�3���᧻�+WL�Է����dAe�޻/:-I�6zH�r����lt}5�}������H(�,����|68�۸�d�=�0�e���]���Q#�����9�}<6m2�x|��ʈ>z������r��uЄ���Ӳ�/��}��!�N�k�X�%Jy��7Z58��ǋ_g��%��x������DW�?����|�Gg�Aj�O<8$D�|��.
G�����EYfc�� ��|�m�$aigb�2����`Nk�#����;YTe�K,�+�S:����qd�=��)ZWѼ��K�z�W�Q���F���)l��A�Ɓ>�7���Q��=�A��Y��������R��A�e��C���:�7M�"[Dͪ�
�eЪ���>$���\����^����x�1�;+-(�B�6�k��7jz��bC}�>i9W�w޴j���~�3A�h��:-Þ(ĕ�p�Q��-\U���������B�W����_��£����.���|=������uy�ݸ�u�x4�Ll�m����Q��4O=�@��|��"g�E��F�8��W�uzU�os����T�|�<� �s�'n5��2�d4m��k��[��o������iθ��[�8v���Ź6@�q�����5��fI�Z��CPy)@Iw���
��Nº�B���*O���4k,��>f��m�+Ǆ��}p��~�=����9�'��#�a �ŵ�v��E�٦
�n3jf���tӞ���C�������c}����l:T-�tr��k���UL���l����('�����-�|�p���m���1�'���/��8��#����!���ޖe²��#�b���k?�X�5�)&ᙓl�iZ�����z��@�Ht-?ϊ��[�;�1�v���"��[Q��l�k>�@'�S�9@��(XL}��b�h�?���fI����WR���ϻ_�%P��	P d�;b,'�/ɖ:��K��z�y�,�61 2x��%�Ϻ|[��k�K�lDu�w4����lkB�_�6>���0I����/�#$�j���ڢ\���1m�� B�G�j��Ǚ4���<���;�)/(aV��Gr�:���Y���4e�z�i�ᚯ�:
��T9�L	�F�}~�J�	��0Zkt��ɾ[��쉷�ǿ�`���&��ԝSq�W?��s�J�	�$���T/
f9���	+���!M���a�{/f��Ȋ���-�;}�w���c����/��(���Ua��Iap<��5��|��3���0p��PFe�W
6=zB�;W�B���3��: r�1�䙥�����=�y��f�
�^#�rNfb4�2��:�:�<.��K�&���Cu�p	^ոj֯P��y�g��~.�C�X��v�Tdh���m7�����B�Ls��-�x}�n�i2]N�L=�9�s&�����l�qB�&�y��g�����z*9�$����� ��x���}*h��U�&������fа
gN??�1�[(݁��)�<�{ș]��VF:*�(��$�:��8���(��-��a
x7��-[�!�y��!��
����]0҄նA��+����۹�d[rm�V��/�D �!���H7bs0x��mq>������7��m��X�ȉ��O�yMýO[�&�d5 2"@�t\$1{0��߹��0�E"@��	�S7(#�J��	Ms��-G��hČt�`��q)��`��|L+q:�z[߉�q�'�5p�TJ��Ң�*��E��[^��0����<�a�����3�6A���➷hzV2�O0���2�����yP�h�z1�\�N��hT��z���I@Ay}��߀e�K��$ӈ���m#�n���?��']��֢S
^HN^�����D��X�*fV �g%��H��5�O}�^9J��0��[��a,h:V\Rc!��͵�G�\�et��o���9t.f�C�$ �ߠ�((����ř߲��������A��?B���qZ��Sc������Ը��[N��@���ȹ��֠�$A�w��k�ӧ 2w8��k�u>XT�\H 6�W`>Rh#�jED4��[6���ɞ��_T��e�Ñ���/��	�hO1�jO��>�q<(�W��$�M���EJCX�()�Α��F]�&����􏂸�'��/<+�T �g�l�r̘��	�����aC��3�4�����4V	9V�Q�]��q �ǯ�l�ܬܶ&���I��0�� �CW.ؐ��hL�#�����N�W4��n�VQ��B�,�Z̴�|���.#�if���N���Wn����zX<�9T� O��g@���(Z� p� �}�E�J�3��Uϣ�W���q�B�aH@��`@���Kpg�#,�O)���*,!�}+@��y+�i�|:Hm����pl�0�Gw:�^a؃�n��N格o�!���f����i�,,G�<���Շ�xo�4^J㳉1v�3H8+���4�yQ`��m�*�,��6�a׷�r%����\��[Tm�:~��*#޵�遂R*|�h�G*yJxX+m���7J�t�T^����#�Av���h8c�[#�Of2Y,�9��z�=w(�M��{$N����|��cɋ�UJ�rO%�P�Ib�V�ul�5�:ژ�Y����Lu��/�'��C� �N!n*���^2�	�@y�51X��5b�Ts0f`���"Ӎ]7_������;��*���&�[�+{�-���x� �`7V��M�N����֞�ip59��Iy�y�_n�V$��1�_�v�� ������k#���c	�.@�Z�.>�^/��M&���4]�ab�#.�>��>���F�J+(䂬���>E�_��A�RDw�  ��=��S��][I{��!<̤�2̷�Ҧ�Y`;1��y�%���ڳ�V3���L�u�������~�QRC�������ޅS8M&����TE'�C� �ҎC�-��{�9�*8�U����
Xg�Xy���k���Ptl�Y�;i�Y�+a[��J��*�<u��C���A[��%lq�)�WK�#�������^��c��e�Ia���<<
����Vl��ya m���MI!���0���޳Je V���f+DBID*	-�F4��Ó�tI���p�l�x	Y:�)V@�z��������K�����D�N��.Z���RF�~�� �܃ay���8k��@$M�z�'qHa.K�睶�[�t�Pƌ�U���|ܭ_��W��l���'z����Z-�7 �nǶ�Lc&��Sr������9BŮ���3f���n5A~߃��po��{�P��~�N��D��	A�Se�i �6ow��( �&��z{綡���3~'���Lb�v�-���h\u^���
���~���z�V�f�}�K�ݡ�Q�z|��#+�ƤF$h��>z$7rS`x�{z��So+��<��ʹ�~��T�' szZ���Q�%��FR��/�����~�hF=�QL�T�щ��e��e����$�C����*G�y_c&9��\�`��Vz��"�q�׬�Erg䊯r�N��������	�T�c~����b:���5�.�N$O��\Z�N�xnK�G�k�D�ߘm}z(���DDx���v`㢆�����X]��j�^�KE��j����ĵ ��[�R0/t_pP/�e(�i�.�}}��|�)��@%5ޱ#�>a.h4�gFy=I��<�e��8�	��;5Ñ$ ��j���1"ﲹ�������-�~��흝|���2��&</��´~1QҞ�%'I
7Ez�@8�,]8c>�?��Ur�/�
��Z�9�T�^�U��a�ٛ�?Y`c�$=����;U|���33��ʷ�p+䪅�^QH'#\ޭ�?C������%/��j]v��%��aVߘCc�Ŏ^N��1$����/��&�U�5�G�a�4$~JuW��L�'��;V`ܗJk��e^�jnO��Jk����NШ�87[>�#�p��K3e��?���6���!k��#����4��.��龉� !|[吲�2�B�i�����e�6��?�Э�E@	z�N�^ٔZ&���	蘓�5���Iׄ&� h;�D�S�^���b:�$ P�`qe#>j�w�:�r% CGѡn|ʅ4�O����.Mj��5|�q��vyK����*B
����*�l�$7�.����䠓3 ~��q�o�s�_�ร�, �?6�����B��ؐ� �C��ւ�(������EǮOKM�7�aj�4�gVn��ABLd���w���M�O�$s�2���,뗡	��I؞��O<�^�I�>zrr�DCܥa���Y~�p�Lʔ�	����Xr��RH8��%ɵ�*y��B>�&� 	A�w7�9� {w�d��_��i�^���`*TQ�[$�YSp�T�if�9�����8t�>P��[��p }�r#ͯM�G�DN�G�\}�3� CH�Y���*>^C%�4\������,U}�@R�H��w�� ʶ(� |2��t҂�W��J�M�q��{w�-���3�V�*�vj�w.흗X%G�S����6�	V�I����먯�}e� A��9�vX"{Ϡ�8��N>���T��� ��gI}���a>�7���=�	� TF���Q?������s�}Nǐc�p��v�u���.Zp�}����<�bx�����㖘h�6���W�I��z�ѭ5��W���ߟߵ��7U�t	���rx(#�@���|{?�ę���MΙ�����+Y�zC��$[����g7��I��0BA�9�3�ɧ�@Ybfժ_��@:�Kt���z�{F��ʊY%�;X/��?9]1�Kϵe3��,�A��0��u7�%̻H��R���z͐4A��L� }FK��b��:�Z��]#�ق�"3O�	���EV$6�+hu�by�$����sg1d��脧8�5��t<��� ���(&�) �K��n�FN���NA\y�&�E��Ӥ��o�������	S�Uˑ��"X�AޱD=���2�k�Ͽ]J�;�HS>����@R
1:0�\c1�*�i��,���d�)��K�U�����@]�	���6�/ln�7���m�pTVq����W��|�ū4.�j�F6��_Z�0&���.�{�K�5�6���,��Z}�4��,ɿ�CA�"?7��A)~�c~�T���l������J�������������[E ��8!}6!�GW&�HτP���T�؊y�%�>}<��#��-V>�A�� ��㱳�K����pX�⸎�OQp��-�.]�>���@̷��'��1��7��ء�\E����K���*TQ�7��D��>񵂋��@�
�։ZX���j"VϏ2�#�}�[w�M]��|,sq����{�j)����Y��<��ŕPd�k��`\��5�E��5W��9%�������e��+b8��~AOak����y���D�b��`���^�[�́� 'Q
}`LziQ�kUN��]!��hy�.�"�=^!����P{i�r<��* ���q`��`���ѱ/�^���e���[���tF�^0�.���2�S��.1a�Hs�&)'37j�ފ��N�3.�b_�bZ��XB�)j�4��[m�d���Ԍc�?0�A�w#���?����A}��v�R��f���\��Ǳq9�� ;Usϯ����cC;Ţ0�8�^�#�fWP�\"5�nAS��ױQ��?w`"��7�|XΩ�?� ������R�����1νV��
�{Z����M��IQRA��)nN@�8&\���,��#����J�vPa��Y���6�|yU3�Wʎ,e�̑;��ܢ�}!1߿��8G��zf3��ju��zJ�G��SA��8�����1i~{봨;W_��{Fv�P�4�/X�I;��~s�U�	(17��5iS'�������#\"x�<�%�b ��笺-���{�Ӹ��Ů��?ŵ�fr[�C�9���b6Lmf#�'���<.�&�2s��vۅ���@E�q�
J�?��4H@;���$}j����<���mk��գ�j"�wS`�t6�zvi#a�h�Y/�4����#����јk�v��,\�=���Ƴд���x���U���8����Q����y����z	�	���|T�8�-�$�)~��zZ�r��@~@<�Ig���h���c��P��)�`C��e�j����J��݅��.�?*W��c�ٜ%�g�(JS�UYL;7��I"Ⱦ0����k��m�*�f̊��C�5�"̑y�V~08ۈvH
^���1vS����f����;%�b�y����c��Đ��x�/
��E��{n�\w�Be��t�2g �e����t0=��mu�^R�Nx{�qJ�rĈ0 �K2tw"u_\�k榞2�CzX����k���TS���F�²A��@�bU�GP�v\�?=�w���ɻ���c4����G&]O���'�@=~Dr�L�È�Jp$�u�֍"ߨ�<?���׶XFv�o������n��P �Eʘ�����ԑ�F֥��A�Y!��h*��*�^���%�wc���"f�u��ܺ���$d"I�v6�����P�|���2g������mR�:ڮc؍�?����5�K]�7��g��@�]NZ��/l}c "����Ʌ����p�uk�a�!��.9�����E��m���1k����ۧ5x�0G��w�8rh�F-ES�������%�R,����mg��d�0�Pt�hd�5�?�/��H��L�+��z<f8}	G�X�	�p�(���Q�uޚ-�3�K>��4�Ô��Q��Q[�S.x��$InWƬ	�9j�h��E��=�E(����4"e_)��p������C$�-�������"���uݍG@�����g=�ѝD���#�o����D���^�99T�A�?��t���$W�b���>I���Q7b�q����T�		���;>-&�Χ!#2���+���.�$?�<	1�>�hn{5�&���#�=�Ո1�*���Y�r J蝏-dIt=�7�:��6��^I7��2�n��_�!���T:�'�@%��u_@��6��p�M�i�[^�!�*a����d/`���9H�ޑ3�(t&^{vî{���D�~Luj�I?�W��.�4�EI�(���'����ss#A:�Cp*`���Y�WPa)��1�-��m^��,���;����s67���2{'c�|�R�X��FҖxZ~�8j�G�R��췯�>���{�`B�r#<��s7ڍ���lb���[������c��1aTSvX��� h{�Ӈ�I?$6s�y�knc�K�� E̃�s+��L���=I�l��9^����]v�zP�'u�9�4���25t|sc���� |��v)�T������`�R������7�4]�`���d��h}�`"�/��`� |�W9�x碋����1�v��hג���^��#�Aݹ���p�#3L�S^�JwHn�l�IE�L�?_qK�Gʙ$�@��+���/�){�������������t�|W���1��ܼ�UT��}o�������t��V�F"�ɰO�q��֏�g����ߎ�����p�������h����;��eж{�e�"ʔJ�{f�s6ѶK�{v3nxix��Z6�(L��� =J=�w8Ok+��P�VG�nz�K�->:+4j[�B�0ۨ.@���`?���̞�I�]Z�9�ڸ��8j����Bb�Gx��/x(���W��%�a$ˢ��G�\ߧ�n��X!*X�/�E�~��{��Ώf�-;[�3�2���lg�ԯ�bB���`���f�iW��Ws�X̓]/�Ƕ�쪂ۗO�ӔE��O�^G�+��3sDk�1u�w%���旒�1c!�9�nbD�����}YW�5Q�ň��!1V�0���%�u&��Uc&9ȩ_L{Ȫ|#�Hef�
�l���Lv��Gr�LW4PL���ܲt �M֮�D�s-�o��)F��5���}\>p`���*���?�;]=�A��H���ycщ���ЮV���Ofu�%Z|���"��R �=}%TPB2�a?�atM��j��!1*[��1�� n�17�:B�J�K
	vs�X�"����(����m}�~���>�3��	�e�;ME~pc����S�^�?�0ՇW]�c���);�~�	U=�uy���r�=�$�4��4���	��Bn����<����V�Gf�[j9ND�ʢaC��k.�nPQ���"�s��i����PZ������nbF�l;T�t�Bԭ�٫ė\S��H&�����t�^z��%��DAaxR�&������ynr�����B8�^���Kܟ��py���!����gVjf
0Љ��U�"�~������Ɂ�ҳ4B�l��:~��׀
�=0�>%Z�}^h`����Sc��m����q]���g���V�ꗮ{	�TPff,��M��z�E�-u�Fj�s߉�h��Y�SΛ��xk��K8����T�t�"eh�=7%��:�E�~�B����
�3��������ԑM�t����Wkht���r@�I6��n����u�cu+B�ၷi�R����O��(�R���i� 
f\/޴�!g=�8�q�*�U������/gM��#f�7��v]"&ـ��Ӂ��r��� ���C����uZ��X���]#7���x���2�U?KA���Ԗ�Qg.���О�h��������/D޵],��:I�Q�'�l�k�k�ӆ,���1��,k��)�$���z/[�*��;$4���h�=�<�� Z��6o����o��;5�!=�L�f<M�8�2<C�u��\�Bu���ʰ�}�4_ۚ�U�Ƅy�1��I�]���m��3�|�fe⡅����o�9�*��wh��ݗSߨ��K�y�����w�&��/��~[�C���� #�i�Xwz%�������i�5�vf��)���P����)h7ײ�.X�+ �G�d��t�p�o٬�\)��
�D`\s�ی�W�8R|ֿN���P{��i�1F{E��N�⧩-Lg��e��Ӟ��#� (�.����-h�|S����Uo(U�|'�N+�����K_�ˈ��~�MΙ�Z"L%��K�)����ϥ�{�r�%K��&������F9�c£����ȯ���Yp�|[�rNZJ��f���[m$	�V,W`|C 8����Ze.�X���Ͼ4�e��7��گ�lg��n�Ʉ�E�uQB���U�j���)�t<�tA��ל���U�]�*��h�y��CK�L3'zF�X�_�]��K0�v�եV���G�j�¯��7����ud�L�$���hۨb����>�JB�t�_-KU�Q1��u��a�=`r��� �$�� ��fp9Z�<��Yr�4��?���g� !�|�kDoXZW&\O�a
#���2U
��~�'��bz�6T�mj�s ���H$�7n�S&*B;�'�2��p��V�ԯ촛��*hG�-�ҖW	�#�(��Fi�p�qb�PS �;������-�&�X����?�rԷ��Z�"C�>/;�_��A's�o v���|E��ܞ�����VzAվa�ӵC��䉕/�Ԏ]����S��t�����@p�wf��t�<4n/$\�P���aw̝�o�OX�J��/Z�'e�87F2:��#�wb���W���|�^n����8?�FT !���"�~�qK�'��J�7������Au��-�������KɕWqBm��1�P*Tm�
�܉��Aq_&�	�OzphN�,�g�D>l�ٲl�)-�Ւ{��-}��(�6z��<,�@��)�Rh�+���Eө�L��Ͳ�{��le����v͇Q�� $O?����+��N��U���,5�B!&�8�R�/?M���4�8�;�<.0u냺������Θ1�Z�(�����fr� 9��#b:+�A��sC^�t���<޴i�q��H�^��?\�&A�Xw���k� �2�6��y7���4,�[Z[����������&��kgSj-5ь�n�"�¶3����&R�'��7��oҵ�c�ܪyԃrc8L�z�,<��gM�Wh��S�xZJ�au���2���GE{Z9U&���+���+�Mq��(�tw�،�j�1�'��@��Z��|]��*���fs*�'�։�����4���~�*���Z�~�x���|�H1��p,e�4gl�;������~{��8k6�hI��;�ܤQ�wG��UCѳ�Ol�J�;�<O�-0�H���F�3|z�'�e�8d�,Z\���;���Y.3���((1	<����e��5���c]���9����A����"����8����6F>gWZ�μ�%��r��u�����P���ѵ[�Ga��@���F��G� �|���
<��E��y���h���!#u�X��6�e%f dtw��	���<��-ꚃ����P)�jM��K����m�+^K�\�E���5���F���x�0��q���8D�]��w�ޏtNv;��܁v�.У�eC�Ȳp݉�Q�����*:rV ������W�n�iW�S'�R����΍���(r�]k�~$j9�}$Pd��r�ȁq��w#R^V�ӏ�>�.YCN���U�#cY&8��!ڭ�I~�}�-"�r��Hj�#�En�1���	\j�E{R���eg�A�HldZP.�P���p-䱲d*/:H%[��<���-�IomU�����o��k�>%s�6���<fC;��F�[�+�v'���F��$�tm��F:疬���r+Bz���v�N�joF�x)]@A+fH��l%�5�A=H0D��ڋ�ZF����:\�LjRJ�gG����Lq�UO@ؠ5�Y��V��r��:I��A���~c�3����mq��v`k���L:SŎ���g�\��`y|ן(���%fUy�%Hue��
�O��(Y�O [�9*�L�U*�YZY�dp�"S ��䲵kL:u�ƽ4�c����'���T�0�@ч��IS�>6�t���ez(m��D8��W8�(��H �� 	�I�ΗBmR��S��6];��@�,��������%��|Ry�凝��dߨ�{�[rN(�@����Ru��'c'Sg'T"0���:�k_ ����n���c̎�c����#e�����$ A^|e}�ﻰ�#��$�����N�]��^�\߱��e��
�����iN�5���:*L}s��Zp�ׂ6�����ß��.�O^��!Q�͛9�LI*��Ҭ��-���*�2��(;n�	}߱T���#U�b���t�}��C[�-�(%�KD�
�~���M�_�,y�9ۤ�g�!���捎��V(՟ ���wT:��@P>$VFH�Tů˻mϧ`����N�R*�3v���
�F�YPN��lX�Ӏ�Y��t]�Θ��տ��(����܎^��S��O�b(~���t��KR��z�눁k�����Tz
���'ە���J��E�G�mF�Ch6�:ᣛ�x�%�!+�B����r\��j-;��H��替�?�Si��!�C�N� �y�QW��o�Hc��\~��� S�U�f���E�ST�Բ�hٶ�9x�fe |aJ	�گ�a��t���ժ�T���1':��p0�`<����G ��r�;A�r�Z�q���ќ�pYĵZ<�UN[�J<���0����������LC�B�0 `�8_�L��M��m��{�&;�n^9sKy83E<V;��}UJ�y��I-���: )x�8S��v�C��R�xJu0���T+ �b�V�>dH ��?�`�Y���ŋ� �u�T[o���5,�[�h_��5���1%0oO��k�?��䖛.S�.�H��0�ޗy�����6�<Z����xǍ�.g����\j���ʨ%�d���E�XR�ls�FD������a�d7��y\��M���N�j0;��pX�|ftx��)��#�-16�l�:3Wu�?��tD�S�_p�E�r����v�����!����>Jle֙�T�� �^�?f��7`5���q�qZ/��\�j�iA��E;����1�Rӻw�I �@������	���-c@�-)�{���'��7q���޹�4B�Ed�T�:�:3X�u���Z[K$�Ώ�8o?����o�T�L��=�l%h���h^��ހ?�j���	�U�¨r��:��S��f�-	�Re=d�Ұ}T٤k��=5�vK����H�B�����s�?�0A�$�n���g��5X�p���f��_��Y�Z�f��id�}0�QbCw���˳��	E�_Rwv����p@��65M�Ð��D��ͱ3� qv�m6x�%���}Y�F"���_^a1�tbK9�r{���:����lZ�<j�nEb�R|�N��|�.�i~¬��@L���:��kY5����2I_jl�>�@�q0�ި��gO� �o�C�7@?�Q%κ��yݽ "C4څ�I�7�y��9�qM�L>�ŷyp�_а�P)`r��~K	l}��48�]��k�9S��Kh��+����,�>�9r�ݢ�3�Ќ����nս�z�V�u�qGG}V�O�3F��F�-�JM�$���O��B�Bmu���<����B6�T<Q�Y6���)>��t�[lr&��n��<Щ�7"�ꗀ�Rذ;�[�r��Ջ<�M��ci<Hӣ{E�k.��Y��hH��L+�l$�`����@����2�Un�X$6�^��(vx��ky����,�9Pr�=��h5�^�|��/�o��h� ��[(w�'��H�ǹ��q�w�������ޮ-���X)�:N~�./��/$��L�xiqB없{%�#1W�#�;	.kj;�`�DT[7&��ڛ5�A�4�X��Q��