��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����u���y��O?��u���
���XI�����e�����Z|��<��@N�B���dK�s���Y|�0�����H���-���6S����+v>3g?��a�u�8�1k���t՝�5� �8ؾ�T�n�T2�DjD�^扷>,,��?���m�B�fP٤�h�驲o%Hۉ��_-� +S~_�j����m�Rr(@6µž����ƹ]/���Q��)��e2�q���Q}@(sZ��\@6:�̤* m�����Y����U+����0u��QP����x[�����W�^A�OR��O��r�qG����6��s�`�@�qZ�3�����ah�RoѺ�@]��>��H��|���>+O-Y�!����(�������J�ڄ��+�#3�I�@S�)i��j��*��XG�T�emr��
�[��h)�y#A����
����ϩ�>�����n��F���Eo�R�Q���E�/M�ps��\D��>�0�9>秼e��h�"�Pi�B�
h�9U������㛅���ѵLsX��{k���UJl38���
���} 4��iM�.Hf��QU�+�dh�[B!�ώ��w�<�,9ΔoNآ�}c�z�(ޢoD_6|��cv�$[�� ����zIw� �v�,F0��uV�InzĹm֧������*�g
�A#�sr�������ĩQ���峀�KT���Z�`��4+�2��MV���Eh���G
䛫j��9t�^a1�Z�g.�n� �p�x�����i��L�!�L&�۵_�!T�)(���� g6Tƪ�Έ�� ���>�[_�J�ډ)�����wg����cλ�<F��[:&Pgּ�H�$����Ƈ�g��Po;E���ѐ ��_1+dv�|�}��04I霯K`f��������jQ��[����P�[����K��Yr���VVĢii����"�o}՗�ت&�̾����~�{f�N�l��6^�B��@˴�4C1�6�f��A�5C?#��]٥�C��œSm��Z����{5�z��_�&�����g��Ӵ�-:�lG�S��+s��^���n�y���|�7X�H�<5��_���uیaZ��V��N˷0@LL�O<O�f�iD�����.�����Nl2�8�F�� �-��b(q/T���;T��p�9�(�$�d����r-��8����RX!}�E��'�x_z��$ d��Zg�B�g���.� �KMp����Zp�׈�z@(P��ѿ��X�K�;z����K!(���;R�� }�̞�T2��M.[���A�[X]K�i�{�;�'��tB���I_��n.��Q�m�U�!�*�Ýt=��p��i�{6����BQI����?�:�P�T����kc�aM��P�2���ۊ�KMFU�ܺ��@�S���K}P%���v��d~������m����f�~f���J�T!��V=��2�O���T(=�t��N�9V9^k�� �G���E*�1pd�zOH5�������*�ZD2��3��v@K~2��<������0\��=͒�:z�`K�7�x�k����g�����_V��=h��k�$Q^�Td�_ch3}f��L�ز��+��'��8�@��-�zN�qhp¥��Ø���I�?Gx�� q��1�Qy.|�[���4���,��n���dn�{�Q�|�����7X��"���[�l�T��Zޫ��1�ib/���Tj<缟W��$�>@��cٺ��;@���Ӿ�KV���������qz����@��t[�/�Z95���J�B����@X�ζ%�7����ܘS���q��Q�5��j�rE78楁n����}�^��:��	{��D'Vq�����7ݫ�8l�y��m�qWu��S��2��4�k�6M��>�o[�{+��.e״Ls0A�� l'�f]��[�������c���7`5�	,R��\�V_u�Q}�8���#��|�Z����+a�fsب�&g#�9m�����#* �K�3o�њ'�,|u��b,k���4�ɶ��t���I,Gҍ�?�Ā;�7d�f�w��w��ao����+6ܘ�?s|����[���^��Y�q8���.��r�m��B�  ��ˡ�.���k0���7#S��	�S��M)Z��Yf��hgP!�M�ydv�N-cj EW_Q���Z#&��̵O�|�1x�7��� ��a�-%\w�M4v���@�;� e'�s
W����^h���S�7��?��[�0��� ��X�:M��H�atU�?���uN�-����ay융�.T-�pa� �P��/gv+��ڽ�BJ[��K�(!�k����.����'l�K�e���;X�ΐ�S��ƢĖ>��,&Ez����P�h�z��� �Y���Ŏ�J� !�a'Њ��,�٥/Q�J�u�V[ǌ!С�pz�8A�6�����ǱY�J�3>?����E@>g�n^
��R���5n�P�?I\�m���e$n��ĵk�z�0m�,�ĸ�-���O��b~�Y�����N�]�e<���qL(B�i/s�w��J�c�R��8?�d�և��7����(����d�G�&随��E�E��|��j	�jz�7K��g�Br��|��_jw"�Y忖|;\�U��n��"����X|և�ÖQ���P�W���vs���rB��*;��d8��A�P���i'`�OX�;A�����kˆ�=S�~����ݝ&����3������w�aZ���ɲ��~/0n4Z��ɱA�6��J-�F���|�e�tļ�ij3;�k�7�W�{���G<���&�&��QM�iw�����0����sɠ8%�z�/@g�?��7���������y��R ���6T��4�̹�D�.~ݭ?�:~瘉d{�Ԓk</��P�k5���Q!_�q������Դw
@�B3+�opӉ���ݠ��q�����RV�S��TN �D��~~�����|o9�+7�����K��F:�� �`�({0{�Nt;��1��=]�`m��х	����T��%��ƶ�������bq���tO��]Z�=@C����0��w*�{����*�k?�k��Ll�����7ь���B�j�3s��������{@��Ho�&�S@)�e!:E�� �_�KyzO�i�������+J�vj^8�Pa`��_��N{�O�%C���<ӑ���{_�!Pu1/���wX�*"I��0�}���OU�m^�n�{_� rY<�1`+)䁷����l���l_�q�m�1yS3��繌���K�cә�K�`G^'�xY���k���~�<���%i<�;��e*��h�+<�Q����	k/,D��.���k�'�%�n+�!8T^7���"���MK�+��y'��R�MOq.��e�u7$�Y/p� o#
iО�yao(b8�͢�����3�O�Űi���Y��%�J�Z)u�'�#k�i�����2�\{�?J�@9 ޚi����1d㱞�`�K�f�a�L� �W]u�=�8���Q��˦�~ʙ4�g�:��g�ٟd>b�aHi5_�c�$�����焢o\�Y�nM@�
�>�IcN�5���ooQ2�m+�2|5{ɾ�r��*C�Ꙟ��1�� /ɵ���G��T�{�|��Ň'p�m,Ej2<!4�X:6;�9��t�!1���tye��ٱP�Ͳ�~�F.׋xWE(��n�<j�v��'��.�S�����t�L�."R<�Q۸���.ʝz�y��,T�9�(4v��t�*��a�C����ը��(�a��c~�����mv�F�.���>���_�0uM���P�ZQߋr�	(}�mU<��]-ia�����П�S�~�m-dxz:$��S� ���S�u�<��h�� ���1��M��s��d�=L~�Z1+y8VTK35��]���A>�Q�'�r�l��|�ߑ��ү��=����٭�	�CWG]�z�*"�q���$��@���M�1���Zp����Wy>�r�>JQ��o�Fd�`M�_z��2=Ull�PD�7)⛔F���Fu�(������{��Q����0/Y'ߚ3uar�C�
��T�70��KO{�k*�fۿ]�Oᲅ��W�LgYn5,zZF�0'�`��>?��7Œ�@ϗ^��p�����03��,]�!����?�(1�ն��OΔ��M�O �8ng#e�<����SY_+ɴ� �������H<����5�KL=��"13.�N�6)��m��ד�nhw�*�CI�jw�xeֳǬ��O9zb{|���@�i�}��& �'XJȊB��E�J���UH��i�\�SjBo(��H?Ϩ/��\K�qy�\�9�"� �L^�CK%Fa��9��xs��|]�AJ�&O~�wJw V\�N:��&6Q�	8����N���d��Y͕������41��X�}�	�k�-�q��ɲ��1ifY}��e� �X�Q��|��!�voIyr�1���6�f�"�X��L?����ǌ����?C��Я ��a���?����ޢ:�nԌ~F�e�d�L��Tjw�f1�#l�������K�P�b_G.���uN2�S��9CSn֌�c��Mo�a�E�6�n�D���r>�A;M
5�Ї?�9t���H�����ü_%:`�{r�285���T�VD\��)��|�&_cm�>j�BTӟr������{�Dz �}1B�x��*�{�M�ҙ'��2�����Ԫ��-���e�ѩ-��ʌeG�|JO���Q����<�8�ڗ���#�NA��"j	F���Ez^�A��ͷ�κ$�:����x��:KZ]F�1���Ȅ�PC���:�֦�&�hՖ���a�/������2�U0fKN_���i�{�U��6���d��E���hj�?�@�ߠg�Wy%�ϽfM���D�+�������fW�b;h
���$a|��`W{(����q�0��~��)��$�I��� ��u>$����r˩߰�u �PЧ�ise�W�q(�³sW�:�6���@&�J����/�:��%�'`�ob$�X������m�ˆ���m�%)�A�+WU�7���$H���?�IK�Aݓz\a�o��5��5�ψU��*�K{�6�Ԑ�����L!�vT�0�{��CD]���T���C�k�����ͦ>~�T�j�.i`a�&����9�Vw�l}�q?�������P�3�D�	�@ �&R�G]�|]�i3��.����_�	�ѭ��[h���U�ҷS~y���E�������'��'R�&s6"���V�9(��y��ݐӯ��I(�
��cI��@����z�z`7';_MT�k�mA�e�5����I-� �h|ҢGf���6�,���D�[٦:����5k�S֖��O_;�?,A£P��v�d�Xd���ؑ�����fU�?=�g�2�J�B��	n��
�Z�%g�B)�Y9���X���WQ4��@��⋽�	b�=� L4�	y*i�@ҋ�@D1oe������:])3���v���ثj,s'�A4�<F��ޣ�O��$�a}]��P[�Eǧ���H`�i�9V�Q
*p�J���n��z��2k˫!���)��'��6�V\�F���ɝ�賫�^:_��m��A��J=����,5xr�z��Qu�����C@�]���n9 R��H�o��������J�k���r�}R�M��7즼9�Q�b����d\��c��ɣ�z�"��f�cl�(ӹ����t��6{��_��>\��w~�*F*?��V<��$�4�#q�ej��2�����mg��2��Č�N(ÄGa�c�'�냡5�82����(n��%��~)�5��8��^�
irV\k����}��'��V���\�
z��↭E8hBJ�_g�-P��L�5r�Z�r�GV���,��B�բ�:�sPǏ�L�j�����b�b��۬��y�tݯm������	��H��R�a�H��
�|�&�c\�{��`+�l"
�(( c�k)�N�`B?ƼJ-h_D�`�f�c� ��Z�DI0%��E&��7�1U�i���.2$p����;Ep�!ꅽ8�򴹰������ۉ͸���kd	~�$[��)%@���^�H>�$@�e!���8���[r��C���S�
�� �>b-��/��%��_��M1c��.�_���ڌ�d�~�j�.�2al�uL'a��Hw$�]�{�v8�z �:m��ȹ%�ʔ���<x�D�Ŝ�mGy���/O~/��*V�\��/2�R2�蠈m�d��*K�ުK�V%l2�o1�*>����q�f	+=��T���L���@��,�It�O-ؘ``�]a�[K(�rɝ>N��(v}���.���(���]�Aيg��)|p���o���X�%F��N���	tT��N�1f�NϽ�3���%���,���G��w��ck솒���1��+��{�9(y#m[LR�����L	�#��<�e ���NSJ���Y����9-����t��.V�q_!�\h�$6�呓�Wμ��y���ۚ�����3ҙ���j^�d>����)n3��I�5��A(��^���0����l�M��>uV��U��`F��SB�h���LHf��*z4��%�������7�V䅱����Q/aDL��渭-��Q��� �eS���7��g�	!�/_(�
�!��8x3W�ز�Nt�!+�ڃvA�Q&`�Ո��e��w�ht	�Z[XIA�n��gq�"H^*�A���;љ6¶�*�S9p��Kƣz��5�%/P.�<
<�D�Ȍ���Ӵ����_�%�Fk�62\g��IGmRa�M�Y�.��ZXmU�Q���ѱ	���9�9��#���'`���XW+`�S��iF}ƀ����E��!�X�]J���j����ΙȜc0O�]�R�?��`�,u��z�f�P��.k��&z�=CI��±�
pۤo�,n1��2��󫟂���������r�f��8E�NKl�H������3�$	���M�
�
~t��2g"Akɰ��i�Sd��u����4E���V�>�wiƃr��v��:~��u�=���7	�>!���-b��ċ�/A"q�r+�cTn�G�cD�i8/�j�D�ĸ����
2/�q;߫e�'_��y��D�EWo����J��^S]�e_���b��O�}�.�g؉O?��ڄ����te�
��ʉP�&iK����P1L�O5�:bf����!����i~�7��G�[�g��n��0=o화8�8PgBΔW����G���zu�V�&��"��=����x�iu�Ύ+,�h������2�^�����pNI��J��i��:�j��j/\{���\y�Ñv��|l�ҧ	Y�pthy&�Bqba����\�S(�b,E��Z}x8)�nl��B�2Ç�/��M0QP҃=kL�b�{�k�os�ր�ǀ����:%�z9>�y4���V�y����H��D��J���A��߳�咅�$"��vj1���J6zT�Υ	eGeM����2�����$�bE�y���@��e���=OL��w. �CXP3����p�~)���$1I�Tk��/o����_�m.�)����^2[��5��n~�<�!=�Ej9�vi(�y,wp�*L��D�{O��u)R��S�ӹg���=�`m��!hP�c^��C�"<K��_e���o�dZ���\\��@��F���4p�d.	��[���|ߩ�Ӝ���l"U����ܻ�H��ǲT�_H8޹F2e<����J��z>�o�Ѕ$Y�U�u�nL�t̎Լ�6��u��g�nu~;����6��ǋ��%�14���ݡ#a�2�����1"s�J]�w�K�B�o�7���ύRQ_��w���j9_RY���|�A�����:a*���ܧn��<
�K���9:߂H4�F� `�	��p��i@M�`�XV�T��%� ��q�c�j����ݒ��ƶ�3�N��O0㷘�֮�ֿ���)u)��;�N�ͩ<0%p#�c �'0yl�&��#��1
Ʀ�5��<@�	�޾vML��^���p�|Ӡ*��9�(O��{rB�)#]�[͹U�8�'�0a�����<��<� ĘB�9U�y� �K�)ߧ��^��|=Q>��3�:�XV���F2Cp���\3;If��W��V�
��R��!A�;�`E��*��a��6 �����h�������UGm8ͼ�8_z���R�X�'�ÇZ�YY�U�B�m��XqL{�6|��~����Z�}������G8F�u���L��w�B�/�wN�9o3֛��5#0Ѹ��qnv��5p�5�?�ӲV��n��Q�{(g[0�ez�a�C"x%�jp�|u�.�
T���Z�=���]-e��dn�'\Ye+#��a5q	�l�%-�}�f_�9Z*r*lb�lEr1Vib}��P�zV����ʥ��c~�y]C+I�*�_!c�֮y6�C���߳��a�H�j׌��������y���<`#�S}'�p�q�����e��;��tf���-�O`��rE7Cۿ�j�:���?o>��	rJe&9B��P�����~<�ȠK���xk��a+ӁEJe,Z�h�3���Y��{_�t%p�=M�lW>�I ��)�]�E��9�q��p�>�et
e�Ic)
��(��+L��,�W	Aӗ#g6e EA�_ԛ/D� ��C:O�e8
������p��6m�S�$4H�/tt�"S�Eʡ`x6֧���ԆwKa�L�]��TD{wi������5���;dY
]n�:��/L��Y�%�E�O$>ەW�66�R�4�
�g
���a@��"��k�����d#���0�0���z0�\b�K�Bӷ���I�zː���|�����_?�#�2�h���[���B�^!_Jy}�67P�����1��[��G�FQ딝U𾾘��f(��=n۴�Pe�	�flZpolY�^�`�V
=H�����Dy"7�.h�����:����;bz��u�u����?tү}�o�L�+H�[MWC�\���wm{���t���j��E���fr��h�0�on��|�m����R���gjR���<j�P�
��&��5U��1R��O�_�p kF����:�K<�lpt�֊Uk�� 8�H�P��
i���*ќ9V�#��['�I���Q�ёi�C�l����+�@T�����	���7��\L���q"��'�NN��s���31�g\q�/.�׾i���W����51�-�J�����Փǽ���`.���b؛������Y.�O5x~�h2�W�v"G4��VJ����0��Q%�	�3��tZ+�6��d�$�c�����t��­�j0���P�I��Ge�0���)js|��;Ԍ���o�����_c��	�XW���q��졗m¹�9��h���mRL�(.x}��K n0������U�;5_��qn9���T��c-.��OG���
^ҵ7Q�U�~��%���i�31#�Ѭ��M���Z�w"��oc�X���H/~U �+I���qgzXE�[�=��VX����ɓ���41lݛ�C�*]߇�7a���d����E�.�RM[���nD(�ͧO�Q�V�_���-�P�7B�)жj�
�!j˘�>]����M��6�w=U-�o�T�ŶD�<ܚ������<�6�`H X	��ӹ��m��hLVt��. �>��r$@	�B�п�tQP)s�l�#��&"������%�Ļ�&�R�1lC�J�M�����Yy~�L(��Gh���y�lc��(o��p�C���6rk���Ϊ�O��c{��a��=<�;������|;�C�s(Jk&�7�ٰ/�Q��y�q5�Yq����AswH��(<%:Dg�,m6�����+?v�B;�E��@��ݸ�Ք��,ҚpY�����o'��Ve�0����0�~�:!DNd���k /F�fڍ���v9�W���m��_T������t���hh��_[��["�U,7䅧GpO�j��a�-x̳�vH���ͩ��p>w�'��]�GV�g�|!7�_(z,D��%��k �����d�`&ߪnB&�U��siu6|����e6x|t!�6�lҸ�lJ��{�	���q��Zaʡ�ٯ��P@�=���gg�\����t���������ɳ��@[�ST$l��0 ?�F/�b�`h��cqyׅ�&H���f;���J2�i�u]���L���G���#���W�|�G�s��S�R�ը馆� F�"M�R���u��I@n�Ta�RV��4<�,2rρ��k����훍�@�{��s>Fs�*���"��[��S�_���KH0߶��̕�:kdi�Xv,!T�}U��o���@�K1N٪Tu�R�c�Β�q���˨O7�`��cz?�.5'��>/�lG֓46Z���l7�VR<[c�a':���th�6���h��9�]K�����5��V�p�8(*:��bǴ���%���j��"u������-@QV��r�6:e`�T���TK��Ť<����K��)�a�]�$�i�j�K�!{�Q��<!{�8���?�l����qA�Dr;-��!����>/�yA"Ǹ�(��'	\�|�50�+{�
��OX~Y*�S�u���p���XW8fШrx70�J��a����sM�_G���I<r��8�-�Z���)H�]�ـ'�G�0���kz7�ঊ��U-�xU'�*��opN��ˎ�R����5����s?�U���u
S�_��٘�o��	��m(�o��(���S�m�5�<���Q�;�'��a���g�����,h�n���eQ�\Z�\�"BFC��؝��5	�;�5����n�5N�ኮ�TI([�q?�2������?2$�Ђ�U7 �@�V-���_3��!�c�4���n$��M]/���@�Z��s��(��� 8�`���A�aڗ������1��P��G�_/�'"=y���+�j��B�����-��-wS�,���]������='��4o�r�7��Uz� 1�p������S�@�C�� ����'�ؙ���=u��q1�J-�]�R%��.ڳN�Vq!��s���v��Z3�'<��/���0Q��.DM�;�J����1X0A��)���}�u�`��� >Q�Y���6�jIƏk������us�mW�Aڲ=�bG�$�C���8�Z�RY�)�90lz��u�]�C"D�*���i2��5�'B�����K�S�sp�a<�K�v���x>a��Ҫ���|�#&��A<C�@:,%�rRjJă/�2�%:�Gcz�Y[Ȉ�
���ŷw�Se��lXx0)�zx�-{��KF1-�����mP���]}�
/F|�7\��(ER�����N�3�d{ *�z����Jm���F0�����K ���Y�H�K�w���t:r�@�!�sp~ϰ)�j��Ja^v����u�vY6����ő��#TL����n����/�`biD�o|(w�+�qs�p��ߛ�&�:j�,\�yY��a�fU��2g�';3�9�hgU6ҼA�Kݣ*��ރ!X�zu,
�������^&f|91�M�g'�^yҶ�hTm�KN��lYId�g�ZY0�*��x��m�0Z����g1�w:C��tJK��0i	�r�{>����dH�Bl��J��k�j
�����g`1��}d�F�@���;�d�n��5T�E�v���j�rap��@�Ą1�c�]

}s��՛����q���C�����"`k���Z����6�����S�:#��ի��g�����"+���c&�#<3�P��L�P��7җ�J���?	�t=�P]����J�<�"h�id�t4�3�����:�1��w����*�p;�>=�>HM���fms�)�37Z�<�U�@�}���M3�q�� %��{{W�������uZg)�;j�()����4���4����*bL!E�ňz�v�FE��cu�o��w���M����G�q�S�sQ%Ki��[��%�*4�o�D٪��ܺ���A��o��V����y\@�!�_ �p��#c�3;�r�.�>R�����?�8RHo(�ՌG�xE��i���,��&���±B&A���	��,0ډ㭯MĐ+m��z��3���־0r����-P��," 32jv ]��a��L0F�M��ż�
s)��TN��oݗĊ��]��j�U2X��֌�T���(4SFe�P
�J��#zE?���\��?�S�,�P�V)iΌ���_�؜QZ߇Q �gc� L��8��3lx�IEr�#''��
؃�f�����fe�A�s���é���3X�i�L}^q�W��mb��L�Q��_��"a�=`��]��م3�J��OZۨ��6�A�b�߭�C�v���(�¨'l��id��'�Y�{�l��~�fW�4����i���� )��MT=X|{)�@���r3��K�O��rmn�:x�}�yˇz���8P�I�\��/��e�Ȩ���gG��N?�sѬm�Uh�>����ro|3���2�4+ռ@�������3��V��V�+��!_�Gf
V���0�O��H�M��n�[�s�j����C�dz��<���gYꏾnz4��/E��C-Nu~�IaK�>�t/���YZ;���ފ�d��aO�/��sѧ,B�>hj\I9��"d[�󼑍�-�A�ҍ���皧7��[��RV�� �?闈�&��^�C�Q��P�ۚߛ1j}~��Q�O��^ �x�
_K���[<�S�P��V����Ybhj��_���z1�'*r� ����ug���iP-������F�öT�-Qo�Q布��֜Պ_���A��P��·8�<;4�`��0��}v��4�΅��ߓ��:/�8����Ee&Y�WI���d�JW AxC��#r����zHi�}�| ��I�o��-s�B�e���<��e��f�z�gQ��dS]%ץ1�-ވ�9���+�n՚4���<@f)�Q�QX?R���qB!�xk�C;4��P��D�;>����k?�j�Z�Ӝ�߁z��K1��$jKS���z�"�� �%ݷд��6;vݮ�O W2[����Au�t$���<���l�SI��p3+v2�����6[�I
�Ȗ�<([Se��K��NS_�^qz�^�6�CpC!�_�_g�\���S2����T��S�;ݚ��5\S��`%����5�O/�y6k����J~e�KJ]��hz�ԓh0bZ\}��sߤ\Rf��K��^�\�.��,.ޛ�y۪�(6;�^�]��#~���k���4Y��,��ܳ�������5�B�2Ҍ�M,�f�G�N���P�SR�w���W�%�V�=�F����ZS~�l�3����[??�(V#z�3Z��RG��Y�GdW%"���.W"10^� S�5׫�:��8�:��(�>?xfɹ���^G�/��G�a��	a�И�%�_���U�۵A� u��A��jr��g������f��I�x��ۊ�.75xǻB:~
��:�lsv2�p'Z��oA�N�@�`��`'��ɧ+W�;^`���x�G��Z�J�s��b�#,Zf=^�\t0�yb��� �_��ǤDA�{���~=x��5�V
iM�0=P�)�&�z�X�SV Ȗ 4T7�:�)%4H#$��V4	�4C�2(@@��m�d�(_?����E�a��-�׃j�{�r5����<gW��&�m2�B�{{���l�_γ�)w��\�QNE�E�VF̡g�b]�G P���4%�k�ǳ�@�}Z7;�T_�V�/:��2�/���D{��.2)�@S�B�ہH ?�*�i촧8i�$)�An��ö�3��vP����Ѫ� �X`���/���,��ڋ� �Pw⊶S3�jG�ʽ{Ukk᠗�D42w�`�E�B��L��g���fj
ܬ�K�Ӳ��eGw�O��m��#�z�Ʒ������%%�N<�lC�:N�`��%�5�\B��2���DO�,VoΣ���%�����"��1}�!a&��dW�u{8����ߒ���PR���:�`��B�8y(�/{���E���$����q��f��8�w�v�R�# 6Ԥ�h�	�ߛ5���f�Xz�����T�vl��p8p�QC�S��U��195ՠ���Ƨa�]N��!���g�J]�����J/�;i�H^�Wz(���pΓ�Rv�-f~�S��=N6�w���=�j��	#C����r�"�����h�������
��pG�T���u�`;���>����/u�����.T���?���+=.ʲ�Mq��6������}E͌�b?�vCZV�H��Lĩ�]�ײ��M^`^X�<Gb��Ľ>���I`�ȏ񙜙b����t�̥TQP  f.���у���1�O�#sl�+�V�˙�yajۼ�Qop�ZmV.�}Ҽ�ƺ6hq@TX�-N��cī����<�"p���-�z2^H''����ཻ �VK�P�����봡��L;ut3�4j�����(�m�OP(�e�+�p�Q�%4�!UЇJG/x�\���������j�=]Jn�J������hȧ���`r���}�Ȗ�j@��+΍���JO,?���v����F�N|�<�e;��G�����<�2?$����B/��*4�v�w8�)�H�b����R(�\"k"u��U���^����E��d|��͐X���mU	�t�Mfj�B�>ͯCuĢ�-|�5-h���Ď�fX9�W�%�!�v���ÔWK�-��K3�
!�K��)p���6���=@H��ڏ��
�}P�հ=���9����v+�ǎ�_	��j�����ݺ��5_7�hj�/��g�$���	I� t��'WG�Un��-�o��lq-�_4��o���V��'z�??��}��c)�dvd�T��x�r�ק�d�a�a�v۝9���Mw���
BWYK��� ,���|#�
�h�2���+mҼzobo@	��`  :�1��IEv� I[ۂ��Ō�yn��I8���?C��O�Q�	�F�� �!��!�R���?Ǫ ��gLtN}� 4�n/3�#�ϩ�*[��� v8O���ǌÚb��Uۭ@i�*���x+����1d�I��i�k+	���9{�qS�.Y-[�k�n���y����$����' �ҷ�HN�5��%�{[v� q7�kω��*��k��t% բPL.<����O�ǈ��XN.P��R�:�Z� b�K�6��y�m0[~�P|M�m/�yǇ���w����^��Slt	�c)��[9y ���Y��%\�,p���W�g�nAk�������ƹbu��ڥ��];TQڰW�"�Ę�?�[	p:ЍUm��WG��P-Hø�:Q�O���xz����S!�[z��yXH�/�9 "�J��+���z nNĝ�N7��{i����}�[��I�*ڸ����)������jT0��/�i�Dw�o�y��|s��O_�h~`D�z* �5v�}v�Λ2�j�Af�06���U��_�7٫��K�� V�@Ra��fV0�j�Z㲂�ʉ�N
��X��zhH1��G��;�'�Yf�ݫҜ4{��m�Ot�$s���N��l�z<��c?5H��s��72F�p#/"�yЀzW�B�)Ҹ�9�w�{lC⺨���=CP-^��bz������L��+d��v�NDs�$S��V���n��St��}^����P.�eS/˿�Ŕ���2�y���.hQv�0��5e���2�tC�p�9�����\�_ʔ��ΌG7��|��H.J|V�&�4IzH��⃢��*�3��>�>��bR�j9�`��[  f+�Q�a��)���bK���̖��F$Cs��g.ߘ��Í��w���ZY�y8����vb+����(1�*�u��8�?ɟ�ӻ�)��s���f�{"�u>�N�׃���x�ցIģ��sg`�M6m��O,hZ�]�2ؾ$�
�ƴ_R1 ;��.D��q'�ꔗn����Cx;��Ͷ�\��_H���.����r�����7�q�y��Tr.�|"����3�e�	�3M�!.WD�e/%��gk��=�E�.��p��*]��K���tȂ�_�TG|�O�N����$p ��\���A��Q�D��"�W}����l��_�_;��5H���Vh�<zh�n���Z�n_�|�UJb�����Z�bGV�\���ε�B5[��]hL�]���?LX���&nv����K��:T��?X�
���ho���q8��ob^7s�=�U���:�O��E�|k�N'(��d��kSfz�,wQգ#��tX6�odu&����իB;k�&>X����J��q�$m�],�yJ`�I[j��3z˽F��#�+�֦n�������T��gZu<�#���1�{A�6h�`LE�2�0��,��~�d��< g��O]N�L/�ˑ������U4���s���]�c��!���tڿj�p*[7O�@�R8E�NfJ�=Fӟ@���DHF:����j����en�C�����XÛ�o�(��T(+�c�-Jrq�+�0	� �lرlR1���Xc���
�ҫ8/
�z�x�.���/���>�b,M=\�A e����(J�8��ӌ�S�.ae&B�'�^�CB�4d������'y�<��ӑ������,f�ޯ����:""#��Le�'"$ߢ�	C$s$�=�rT�� �إxL��J,:�pT�M�h�"�VB:����us�h������t�����stGC�}����N�/Nx6Zz؏�x��/���t��. �YS�̯�-q�P�W���
�$}�G��RGz���}�ST���/�=�P�ʗz��jH�� ���K�!Ԛ�ƪ�88� O���W����>9ȡ;
3���7�����Ք;VР/D���y��;��{᱘#롆�\l��4���l�Q�zs�9-;;���U�.�@`2뇲kLCcw(��0��Q̬Ȱ���rV��j��^w
�?���E^��w��L���xDhE�b�Eaj�����'U ��԰��&�wd��h���YC4#o��#��xj̏�� =�Y&�=q�$$��R7�����!�3���pI��ɡO�L��?����QxĉU�y�غ�,�n�����s8���eJIy���%򆡠��M��0J��Rc�K���6��{��פ;�#ӚmG}Y5�Ԅb���8���U�	���{�8T,�@��tUsF��j�B�ڛ��,�5b:�����WK��1��޻�����*I�����A��b	v��5a���A-F)�SZ�kؙ�[�o�kG�D�����Ş%5xx�uw���%����O�t�UV+5`G*[�~H�\�u���m�ʺ�S\��{`�+B�|����m�����j�K4�����,%��6�k����E�k�,$�0���I���1�f��ϪS�c\���A$�@j�h���Vd�hɱ���pFl�~X��ˎ��������/\L��k�vW��8�j<��ҿ�@�)m�md�Rrs���?C�վ�aYë:��f�4�� JpE?{�p��u�p:�搚?<�D�|��r9�S`3�O�F�'Φ*��xf^��m��xi�0_���c��J���x7`I�;��_���`^^�O�$����ў� ~��hw-�:���}��*U��J<��@G� ��1aʛ>���<$���wr��hD����\��_�iO��A����̻a~pQ�n<�V���P���}G?���E����]�ɔ��,�5�YNчJB��A�ϰ���r%'�]'\E%dp�,�%��j��Z�7qVZϊ~V�����Q�$
\��иB�,�*5�	�iX:M���J���v~��m�i>J�2y�bo�OjHsUQ��gC�8�
�z]�����`���1��F)ϳ��S�i����#�9nQF%o�����(4*vG���3��.��@P�u��t�9�<Ų9�0mw-���8@a�;�AOE��P��d���A�z_�<ޚ-dr�ZA��d�ɖ4�J�Z;cm�s��X��6Vz�u���VBԆ}ޘ�U[�w�-8f�����8Bg*��p���G�2�W>(���+�{��uL��
��:��&Eyn�r�K�y���\��Db�QVZ��y�-�_�Y���$%vߧ�ʨ���%�E�ȡJ"Uh���e��6��G&)r�Ѫ�`NP3I����錅S(�@�7ڒ�����^LV�d4~gV4�Z���OI����-�bP��=N�iՌ���MWw���� ��s	�(�u�Ha�99�
�mٓ���1X��sǎ'2m5H^�M�~CKt� 1SEH�O�B�k�R�&#�M��s��1��H_����}?�nט��
�MJ���\E�bׁ�z��Q����8��~�j����P�g�J,ad��gO���{!�=�ڏ��͚�D�����m,��q.ia��T�������.Cu�2ܺ�צw�*��29��1λ�-^G�R[˽@���jɽca��<3��:hm��[?�i��� �$8|Ŭ�ؕR#HS5��z�q��e�����(�������\��6_O�����b��!�s����U����k�(�G[H�(P��zb��"��3�l(F����	����9=ڽ�u�@r�쮆f��lY�N�X��mdVRn((,���&�	e�Ѕ1'�T��SE08��9�E,w�-�"������lY<�?��E/?=�����.����d��wM+
ڶ�#��+
I��,>��D�q����f���V��_ʩ#����J��(" [�
Qp�`�	�Dx�N�����	�d���0��gA��;��(��+!���l��G�G�c	G��Z����֟gJf�k�/��H�G#�9#���8�Rr+t��&hfq�:!�ܝF:Vo��\	c��#�M��4]��_����3�CRތ�N�@��}"G�#4��1����*�%ژ�>�Qr���x�hGq��r�
��>8�6�q��AQ��"{psі��9Ml�bh��S�$
��Tnw�
p���^԰y}=��3����ٻd���1�6�����'�� g8�7���2A뽁)�G��a�����f�Xy���G*o���Gy�8��i\*�2e[�w?׎�N�f�u"� ��$�Z���Hń>߫czvT�J����	|��OجU�"�E����\/�d�U�����[�e��/b /������e��k�D��y��S�L?�<����^��[Vt?W�]@��&����2�	"x^;w���B�	ؖ�w(���Rۥj__*ib1�L�=����w3.��1���Q��c������#hr\�;Q���	?m��#�[�J{�D�5i�N�A|�����p�)J_�~>�'�
|��,���b��x��	���QC���ry�pR=�%���E/�SE�"e%��o}B�C^j|���&�����h�6Ԝ=ަP��~�	�����Yno�͜^�#��B{4��B����1h!&���;]�9�/g[���m(נ����&`�^�j��f�)�s.�o��l�p�=�]Z��3	�ڈ �B�]i��aw��PDO�+E"]�Jm�r<�f�"�41�&�8D����9�9��)�`Y�4����wd�Y=�͜���Ds-��u-�3q)�qt�{�억n�u�}���g��O�c�O$�q�M}�n���"	�O�-��_d����e׎�Ǥ�l�>�h~���f1u�{���@]����PZ�*"��
��^]����Nwp�A9��ƹz����j�#�L*�z�S����bs��v�c���9�����1��NV�-.�n� ێM'��� �7�9����u��w8���B��z�A���!|�}�V���c{�E��[l�a��&�n�i���*-{�CSQ���aY�Ɔkr\U'ur��X}q�u���V�9�S(2����s_�L�d�}v� �����F��^��q�A=��6��da�}$ed@)w	�yy,��,ߠͷ)+v���M��L_#B���v��Et����!^���	����٦`� �y�1�>��S�'���L�O�)Q��̶XU�VxT.��Drέ��~0����W��j�x��{�r]v�B�5I)y����L�n)*�ƙշK��f�	'.���b�"E�O���y���t�	��_�2#	��΋�p#���b8���=r6�Q�`�}��C|C=�M���ơ
�trˮv� ���7��.X������u���tﵣ�J/���.`�b�nڀ�r��VnE��i� �����ܺf��֡��kG_ �3�o�k���1KN�E�
� �B9ʞ�V�u_�=�,��X��6�I�����#,Ug����A��@O�2�=�46C3��;F�:��r�S��7g�-�٤p"N1�v#�����	�/�J��˒�2��Y |�*�b��T�����;bx�r>�p��O&�&G4�դw�"E:Cn��KT����~���G!�ߴ�h�M#��S)��*)��X�y/���q虺_��烞�KS����3ܷܚo�n��qUY:�.�_��]�q��%�`�>���G�G|;� ��sR%��z��~�7E�� �A#�cD��_A��U|�����)�^^ʞw#�<m%3����:S!�0�@نs�Ŗ���u}&�pH�~[�o��h��>=�S'_7m��ƍ߮�dS0&7����.��W��������#�&�>�����]p��*���-�񉶆���=�PaᾄK�U'3��Do�?��r�wv�v�9~��r�IQ��[���)7ʨ5R��Ҍ"���^�oT���"���Z~�>��]�)y����%�;~h����j��P�a����d��b���w��+��]��&��G��`�J)QQ4b�|~�rB�O�kӯ�`s���M��D��������U�M5nunP�Bi�D�.�b��~�q�����f��s�w��<]i;�IKQ��(�p~�����l��GS$���I%lt݃�nԴ����!'�K�(X��!.�1��J��{�M>x�MP��+?��C�w�҅�b�|�t�Ly�B�`����R}(�k�:�C����dm���4��,�i���l�m��[�Z��~�p�X��8���y�E>R/�y�jgIW"��kr27�X�����|�r�a|U ����H"�X3=rv�k�D	�)1!�Ѻe��D#f�ק%�-L�E�g�f�7L�;C�,_�����a��"��D��ra*'��j@��\���[�{��.z� y^������p_=� j�)����|���67�R��t� ��`ygE�:���g�\z��-3���r��)������T5���5�q7�?�kpb�
9�Whe=���7��7�=��٭w��Y����92�m��Ϫ�v��F�S����ӝ�>��#4A俲q�y��=J[��/J$���],ţ��Wxc�������?!bu����I@����L޸;�җ�kJ\��^+� �t�m�.k
gݗ��zJ�8�]��L��>���
�ϲ��c���'
\����^����B�(�?�e�]�r*~A�}�u�J����<����2%��į����~�����{�@�LHG��a{�����c���sg��i5����+�����!�Ɨ��*��b-,���0�#�F�� P@{���%d�T�7��)�z��]���:k6���,�K�P�1!A�V�%c,�m��U�>�l��(Ɉr�L2���UOѴ����1��_��L��������1����:�-�wϒ�:�y�'�thɉ��A��$emȜDy5�K�}LY��7�3g�S�
X�.�rv}���r]��H��u�)�5�q�֬'Vǲ���͓��5�>m��6�d4�F= P�Q�z�H��M}牭��Oeu�@�s��n��y�^US���b�z���/����qN���M�gbB9ÅQ۫� �/F����8��oM,R2ؓc��iq��I>�z�#�:���¿)nV׊�]D�5�d(�!?�`CΤ
���I��P黑�db�tà��?�;M��Z[r���³�%m.�~s[�Є|���r���D53�Y67�����W�m�j3��qEB��s���R�vNr-�`��|N�ɡ�p��54��y����g��d'~R9�Ui���p�GȆ���"Qb���f}@YYl&��dCA"x�2���Z��W�̹q�<�ya��f?��T�.ޔ��ƃN���1b����6�3�^__��d2��\��k�2s;[d��s���X��e�l��e���$��E��7�^+5�օ&77V�V�ށ������6�(yT@2=b�dA�(��A�5���3��/���!^���K��:`�� m���5��`c�ԭX"����)N����kp�{� P����]�%p
��IӒ�a��t���p9�>m�6NםB2@����j��g3���h�eOu<�|�Z�)Z��Tڀ���Qo�P�ZZ'tǲ�l̒ޖ�ľg²�)�Q��!��x�����g�����w
D KնlP�&��7)��L��L�D5��;��f��
j��E+`�2D�3����۸
�����l|�]Fd�3ݖ�O��؋�ȹ43�nX�_$${kbW����p����i�ł�w��`T�����������=����k��[��ƕH��7�O)Nm���R��0+n�p�3�5���Ϙy�A���p/��h<C�⪱D��J�=�(�wK�g��.i���f�޷��/�s�)���gsؽm���P���33���	R�+As7���H��O�Q�Bo,w��b����jZ� q��t3�eKp�����AVƁdi}��V+�ᾎ�y5V*������-3|6b��w�8�¡��_�YB��k�{�ؒBs���r�5Ձ9,�ɓ�(�aͲ�7����.�r��4\\������ ��MBz:̓��3���N'���!�Jo�Nc7Ι�����Q%CS+I�Q+m��n��#��'4�V�Rw�yB�d8���v�RԚ2v�����$�׼^��<�i¯Lt*�	�sD�2ĸ�7�Rw��߰�/��;k����:��u���V�*U^֪�������ߓ��R��̸���I=�7� ��'t'�h �]L%N�2�&�6��S��k*wV{iߕ�2���Ŕ�[0��\X���u�)�[�m<^�Qr��ޏ�d�5���hDV`��`�	���dZ��4~к��Oob&P8���O_�͎��1�	2��q�k⌤>�QS�0���6oi�����p{��P-�cN[@v�#Ժc^��Q��9�M�$�h�ʴj�8$�M}fMvSq)nH�[3u�n�&0Z|�v���ʤ�p;8�t���;���A����_�k޶�V^����5������|�*�ߩe ���>���r*����.ȷ���"Ќ��*��@�ݲ�q\x�<gr����?	���ێ^����n�ei	�7_�l�}�b���]5��'�o��� M�2��������d4��p����7��{#��^,2t����W^�DOj�a��Ĵ;]��ݥ��UrX#��6��Pl#���	�ڕ������$?<-綉Kڵ<�84��`A.�T�j��z��AA���ݶ>����oE��U��L���N8���q��ò�#���Xj��# 4��#=3�-��:���j(.�Na��2tg��pJ�3X�}gT:g�z�Gq��#F�Q<^�C�h�R�i|#��~3�O�{@ῧ�0�`�E)��/KN/�+Ԣ��~ޤ:�0!󗍱�@ᚪ���E�ܠ�����ŀ��k���Ĭ�D�Ih/�E�hI�K���y��셽��^�>�qZ���37үy��@Ed��n{�r��c'aS`�G��\��-��c���::H$����:��[y	J?��$
�ۂ���Z���!�wb�� +�O6��[nЮ>�|���)���.j�� D-#�V�%�ʹ����L�|��%�Y�5���bh�_�� A�_{�އ�� ��-�%�n�RB'��b��f<5�.op��C���.m"�4�*����)��y�P?{~M�u��P�$������20�t���	�n��6I��`D+p9��}m��Y���MQ���Z��X����h@cgKg��}�!��a�Ƚ�e��*::�=��u2?����>�N�,=�� �C��^�z�-�Bus߀�����P����40�mCd~�1��ʂ����U x���ޮ5�	4��~�@��	�]�8H����lb����ok�m��(�f��~�71�nPM�@�p���1�n�h�M�^!�	���D������浩 ^��Q(<��6SL��uY(}���V��Ӱ�$��ۮY�ܽ���j94�
m��8tW���v�_D9��'P/ ��uO�{���M���m��1����Vŭ����Dn�
F��W��������O� ^�y>I��������S�<�jM��k��y7����"�U3x#�c����ʥ�7�	2W�<�X2�s�
�4ӹ,���g��9&�
DTE e[�3��"��Oڗ�{���";W�Ԣ4��Yv�_ǁ����=n���d��2��	�� �_7K�D�+�K�$8��6}���8���a��p�0T�D(�lMRB	���kj�mj����*T�0r�;C�>�[����=Bŕs��0�R� T�)	��ő
 (3}t�l�h��,]D�$�5|^�2���3#��Ϭ�����:O ���QF}�<��8��?��c�lm$�(�]@��7�z�C�.�i�S�r�F�hLz��(��ܘ���t2�i%�/1�I� � ǁ��ۻ�<�dߥ�Q��u�a�=enhm~j��Y��2�' i%�xK� �<l;z����n���o���=�$��)�{���r�z�)KnN=�����D�>q._��QSL�m��Ki��l�\7��ɘ�E�rcAD�Dd��n�4;���xq�O���Ο�I�]&�NQrI� a��Ż�l���ɣ�,v�a���6�(�y��B����8D.�.
�D���"�P}ܩIH��m	�sL@�^�9�$�l���(�7�5e�)p�5x�ꆋ�˵��F��8�W��݃k\�}���H�w�|~��J��˼9�t�Ŭ��2L84�d��/�X)�	֣��B�~
Y�*Cm��n6b���Bj�C/��3f�kn�;X���m1x��2k�#�%�5�XP����#��Qn���X�O�\�s��v���(dơ�q$[�H��_�u�[�n���b�Ћ�\ <��$����z�W��Ooܐ� �{sbY̖��:�R��P��#"q'U��V�Wy|�������?~z����s<�@���t|-�4[�bwW��i���`�R'�F�I�7*U�Ub詔�ս�xB����r�#e{�)�,�ΖD���݈˜�7$�m(��3���0�����Pť��:����G�7@���#[��
�{�-�[c������K#W�ekQ��f'5;nnj�-���`qЈHH0ƺ���|�ۤlTLE�E}UP��Wz���U����pe�r��G��uʩ���"�~v�ѡ��� ��QΉ*4IP�155���Y��kW��i�y�;T
�/����x�ǌ8��{ 1��u6e���� 2D�}��%H�S$�Ɠ�ϣ$j����7��9�|�a5���2�R4����A� i�tg�����ӖE��m��u��r�:�K$$�9��!����-�����(�q���n�?B��Sg��qm�HU��
H\�{ �z.n�z��1�B�]3�Z�F�y��^�XA:l��C�\c�X��wDc������#%Y��e��ԈV{�u�*(z$�JaM����mo;,�&]A�|V�,kO����7����l&!��&��%B�$̛+��B �[m�R�-u?O��rE���p�"��l�R����"��xdXz ��������QYQ�1����/����#���`;v�1v�x {����
mz�y��f!��6�K{�+����W V�8���q��n�/m�Ɉ*�ݑ��e�
�9:�u�l�6q�}nU����� ��HA�w̶N��yS'+�1o�)��Y&�}�8��U@^���*�4Jcl���΍�Y$�[�|�<q~	�&���BR����c�
P��vf�����[�O��%r6�f�,N1P��|�' ���<�i�z`[���0�CN�y�0��v=X	�b�dv�(�I�|r�D6�����n���C��uB<3�~�敵�:��l��A;b��8Q��˱-.Fث��K����fǾ�a����m�L��S�2�����P�D���<���߼�ɖ��%E 銥�g���7���TM�x	����Qn!@��2}� �J��c��˒4s¹oOh�A0m��gէ㎒$K���t� ab�P����{��6�~N<>u\�d��WQ]��G�z]�(��V���U�_�c�*�<�.>I�d��V��fwfb�)����Q�3rn��	�"!5����� �3�=��6��ʽٕ�j5�^��9�h��t�;���}����g�So�|Ű�D�Q�A��Mb4h[�����6�u�.��E�����u �ZK�_� 鯨��_�=2��ӽLM0X�xk���!b�7�j�fl�����J��B���1�f-��u	�d�<4�G�@M�H��	"� �}^�#��$�\^S�]`26RA��~�s�~�A_:��2]��.�8��	Ę]������K��W�r����t��w
%m-���p�a��.sĩ�+_���HYJ=S/�B���-5?�8��{-EI#��2�0���*� �+���ǘ\y��c���Zun�>L�u������֫��m������t��<N�=7w�V�4�������E��f�d�1�^���������T�֧�hQ87%6=�)��AЧt�+�>��|�i�(�E��˟Ԥ�|�A!v�v�U��9�P��M�`�i�t^^��{w����27/��,OB����'�0���c+�f�4_����h$�W��ծPh�����n�M���XC�[aѾ��c8aY���5,M�EhMX2�+G�U����LO�v��ǰA"\��Eq�6�����q��\5�
0{�R̷	Z8�f�1������I0$*��K@���ϵ�75�&8���;>�:��@c�����t���`^�u���;Xb������K�_��<�&�����C�F��˙�]0lٺ!���,j����g����@��v�}�C�g��T=M��^/$@���.8z�L#��d;�� wԛ?���\�О��^އޘh�,>i�a��@�|�����a���"rs8R�>3��q~����s2��pc��3ə9w���绀�Xj�?K�$��b�J�҃�Z׈oI9�6W*�r�:I����F�|�ii(�����VDTp�kt+�9bJ9��W
�U˄y;�.<�����M���	�a�(||���/Ub��7�̹�M�F�_צz�n6���5�����1|�wAe1UA�z�&�-y��cB�;YH`�ϓ�@��Q'W��2(3�i��% �� �sG �B �s���HJ�UJU�38� �+�s#��Q�d�|⥿��3������7X�A*��U���^��䣏���JS�c������%6-E�A�#�/�!�7#Am.����'�c���t]�U���JҎ�G���5U)�q�����Ϭi#%�����$]F��|��D%"�M�*Mr�8�b� X3r=tf�4v�V���r��%wBBUIaù�q�b�=��m4�Z�����dO�_��ނ,��J!rI��~�*B�8��	��v��_tP4�
�y�o�a�yUݻ�3���M�j6�bn�]jy�:�E+�&i
��ٹ� h�C�2�8bW{\v�N�1yt����-�:�2�U�> x�������R!G`iWM�5����T����1�\���bp�R!�.����&��5ؠ?Z�4����/���ʺRR���W�2�M���Q�	��
]ֻva�1=����� ��}L�;�8�yeҝ3��k�{b�Պ,2R"3,�9��x~�J��ӬE>���ќFH��b�H
F�9��@,4��`���P�܁,��z�f�q��Rw�jv�{�^���|�ris���dN{Z�����'녮k���w�E��=k�n�o�ă����@1?E�y�b�i��p%y�ݱ}��N��$ĝ��q��b�@nfߑ����5Zݻ��\	�8�&�쭻3}�I06ei>��X���Q�e8�pΩ��91(�g�j��b���W��,��!�%x��G]a��$�L��z r�drRr����^�="`@�ͼ&��D�e8���ޭp�;���;zJxW��O읍Z/1͘!�<�&�:�fz������0�	l-�,p�s�w��2?pu��<R���bz���]�6ms"�<�� �.d�*����rꯃ��R��x��2�Z��#\�AC��m:��Ps*��f|t��t�\���}��I�?����?�X�HL�B�9�d�%�=���^�|Sf��e�p�R� ���V5H�N��������@����-,�E)h@�)�}�r\��{�%9��I�3����?���1�G4�"�t�J��Ϩ=�.[�YR�ͥ�����i������n�&|�2[$�HF��)9jt�e��8�������3�"�y/�c:���.SIq���L�j�ө6g�b6��kxU���!�W,ϯ# ���TQ���f�BKڟ!� �U���u[�sXHh�g]�!��T�Em�n�� +��hVCX�ՕLuv�_��rK@���$9�!��6z���I��ѫU�X�N��S����E[Z:ζ'rxv�?RBI�`P 
h��3�&�B��`�S-�Plw*,���	�'fC���u�g�4ֆ=�\J|�7�2���޺ 2m!@�8����Il������Q.-n
������e����l���a��O�;�h��M����-s5 ��yi��|TU�M����	�����}�Rԭl!H�:.���8�F�z���T��w�����2�s�:�0�U�����2��"�Vk�"q �`˂��A���m#-[��	���k�Y�sAD �B��y�C��EU���a��m7Ɋ�{�������|�)��B�4-ż�&Z[�&�:���A��ͽ����&͒�_!jV�˿�бVc��<�����hI^M7�O��	�r�Fec�A"(�hz w��e�hͺ�����8��n���3b¨���Ο����>ׯ8����,:"�F�Qvm�����88S)�n�p��ټAo��]x@N��q�P�L��+��@�_�جoK��[�J��u��q���+t:�s]bP�ݗ�Q��h��ʛQ� l$c�L�=<;q㲗הG�P[B!�.m�b�.k;���_q�	���v&���줲ޢ?ہ��}�p��zs/���F�q5��5R���5���iNW!2��)Ў}���]�P����B��l�Dc����Q	��!��Q�a�NGG�L�y;i�L{P��+�xN�9}Dwd�$h�f^��aw�y���4��I������D��϶Nh�D.���Z�+5؎u*n�v�T�V$N|Q����9�V�|j#���۝�x�)O��I�+9��+𹿑<s�$NO�،u�1����a����t����-����JY-�YkL�\��Z'��<$�_����<�.���qc�W/rn�]���eH����+>v^���.�L�Aeh?	fd�_6����Ve�F��o����(<(˃�,���h0a�`�B<�t].��I-���9�Tͺ��RBz�R\�6H��D'��f���0z�=�=-Q!�$�V�4���sd�S�$*\r;���@��~���"U���?~0����~�d,���A�D�&��n�������C�mKo�{ �҆I���7���<|"��(�@�i��"�� r\�]���*�Spj�{�Oُ�E�&��yzX��qj����*�V�`G�jY7����^���]��@�"�����bm��T�טu��M�).Uc���.W8�N��.J��/�4�?���w��:���jp_>�L�eM!G����Ͼ������MW��.(��d4�ۛ9��!G���FM\�{_�~���(C�e�x+�Y����qȥ�"�I�k��@������;:�֝��=��D��t����ڄ�FS��aqJA ��5���|B�=����- kt�X��&��
��J�d H�^bm�u9�X��ã�� �`e�z�2�[�æ��~{����;т��_ATq�1qdhU��������� �*K�1as5i� �S�E!�$>&9~9�|$)�������>��K��� �j������ο�Nk*�o�P2�#���S�b<;��&z���쵪��/Yi�3{ޟ}X-+���Y���a��q�v���Ǽ5��@�����Yv��ͺg�jO6�C������Y�	b3�ĸ�M|P�<GH"C��p�eeA7������U��fX��F^���8�f3��T�ǜ�2�ǿJ�$[*�9���z��QymC�Ak�NC.)Q����4ڦ���駽��ḑ��[ݮv��b�"w�R8_5������{��_6���3��/�Rd7�U��#����lE�"?`ܚ�͌��N��Д��'p$��5������BÅ��I�"����_�dP����B�#� �~�w��k�T�E0�~���l���ތ� �;`q�Շr@V�T�v�JB��%{��aӂ]݌m�w�Ҳ�@e���h?�Bp����-����YI����CI4�a4���X�cK>@���}������t�^�P9&��m�����~���5v����ae3�O�츰7 ��u��5'һ��H��|;xѓ7t6��)�Qǌ�ԇJUEl\�Ǯy�A��$��pK��HL����	y )����ĞRP�ْ3��]͖K����W�I���R���Dw�tSߑ��6�"��S�G��Lْս��C�%&����I AUo�ՋD�I8�%��ô���g�Ӫ�r7x�L��FU q/�,�����K�c2�κ!
+���<f�^�)��ͬwΆ�4��~�>(s�!�% ��i^� ��<��B!��� G^��'��C%�=N�l}-$!�"��&28�b%/�ؽINotWߓ�@�� 24혊k8WɁ��Y+���c��	�E%7�h�Ϝ��/���8�X�]7k���>�&�R�����yt�����C�xΜ��,._�>���0��]��\?3ii���E����i=��U���x��ʯ��28l�<W}����n�T�fgl9E3z�4�ԩM�	��8T���]Q<MD�2��:f����x�^ֵ�z�aЛ��"��K�U�1�{go��-�#q�����>�cf�T>Ch�>��+��
~lȳ��k���D�v\��}��8�w��D�	��e�M�D�,x�זR��V/�����-��p�0�v@-$�K};��1�t����p�#1c�?0b(3�<�V0���}D]'=R�f�w���6����1���2�9DW5w�����,|}2Z�ڇ�~sT 2���*���9��v|�$rňB�����4◟�;�e����V,6td]�o��֠�ѐ�.�Abi0��6�f̖����c$%�C��<��&��D��`����~�\���'��bh�7��׊u�@<�/k;�@���1]/�^P���c�>{^��/��+u�^�����佲+�ꏰ/�h�.���o_�¬�@â�>fw��q��N�/��� ��*qP��{�`n`�泜j�]���P�Q��%��f' �X���������C/j��`mb�#k|���ДlcQ�Y�~�Xd_]�1��P�m�IE`v���KD�m�9?�l������p����`�v���h����N��+�nB��M̡�;h�)4j���^nNoa�Nn�P2FS��0�q�nZ ��0�]�ݩ��%e>׏�2*�I���-��cB͋!�lHG���Z��?���q��iy���;\o0#�O&4�m�a��YkE��еA+ ���z�qޭN��ۚ�7�m��� ����F�4 �6���+|F
�/(e]�������7j�V��z�eW�u�Ȭ�P�I�&���T�e˛0��`Y�ԅ�ô�8��ao���ޣ�y�殖kG��:��(�鐌8���X��]w�������_�}1}�W��4g	7���}��G����^��J�K>y�m��e���?>`�|c`()��;�8�.*�W�<�����Ÿx�0	�\ſf�r��ok��aNt����߽U����׉W������Dh��8L��Lb���E״��(�jQ��~�%w��x3A�Xw�:��2��K:|9�r�]�ât)0�ת�Z�;Ufgr����^%{a�\�(S�t<�F?u"�!Q4o@�����k�l0�������������Eõ9t�m�Z7������Ν�[�un�$`�g���OCl��,����-�h���(��PPʆ��
�R_��Lĵ�"�܆�d��+�ً2��^���^}�#�%���U٧�!�R�}v��kt�Ȝ���5�`9	">ۏ�k���h��dk�~@=H"l�n���
�ɿ0G��[S��Y��=Y�>xd�߀�a��##�X�C^�Hn�|�o�:�)�_ԣq�W1Û�K�����C�J���=S�UL��#Mۿ�K��}L{:�璤�����$k�?�@�����A�U#��|��*{ؚ	ׇ�A�f	M3�a�@�e_[@c�VrG�AhC,�\�!�ի�0��G��@t���4ʡ�Z���,�,7�����G�m�湖�F*?9#�����cO����Š���T�(����_"�j3�tӷ��c�_k����gGL����S^�d@Q��4u� <�A&�B�o�N��FŇJ��l������"���$�Đ�./d=�iB�ʗ���i����TX�#���?J��D���D����	��������*����gʁ�4*������AyQt��er��gI�Hr;�D�#݋"����ĉr��c��Nq�ϗ���#��l�?c˫�|�#͖]=���5����^A��3��Gm�Y���[͆��H�kI]:XM�;D�ښP���-y�kx+��̲$0�9(5�;?�V��/P��1l_��(�]�1��z�.'44˂����|IB#��>��8��pH��nM�)u�����_��<N7�-J/���vt�i�8)�F�\��O�/��&gx)EP�K�d�@~Cy�
L!A�T߬�a��wn���N�@���/��|PI���x��� v������3�E�=�R�t�!K��KdU9�3�����'G�ɨ&�.I�`$'�<;n�8,�tK3�c#��= �����pОFL(�j?I���Ռ�]̗�Dv��zT��n��/�sKD�_e?q�CY�4l}7A�/l���:ՆT~-|���Q���$n��4t�c�BUZ~O�߷r�Ǎ��j�>�?���hJ�A䩕����F�3�[��ot<7�D�c�d'`��[�D�>:\�&���|~��Z��.T�yQ���4��]�t�ꈩ��{�`٠�WF[gc�<��	��7I�J,c�/����	gۣR �=�p�`3�jb 8�-��A�[��3�;
�19���Y�ؾ�i��Go���H+�U���Ċw�ˏ��_+J�j���m��豦�D]��}���(Ը?[4耟u���T�`z�������k#��	�TJx��#�V�XC��iD:i�0���oI��XiR��4�4e�(�	�%��e�z,���6`����:�h>����o�O0e�J�Ty���j�5JNt���^��m�P(�|;�My��G���:^�OR+��s,�@�&lsu~�B�K��.7��K�|��	��v�2���[��aS�'k����ᳲy��Ҩ����G�~m-w�0��B^^6��S���-�=��`�%S�4���:�� B�cB�[��oȵ'�ռTLҿh2뵭��1���^���~ �m2,�<ڦ�PiR�ɠ����z����x�]0�v����@�<���-"W�"�w�y8���o`w�Sv,ƘV��:�\cQni�/�͐ު��pA�T]ԑ ����ʾ�{Fs����e���=r��b5��vK{>����C��_ԝQ�H���lw�Gl!͡$�D�qu����x�A�NĲ���؍}@Tm�Ry�g���o��'��Iww�,1K�*hq5��y��v���`���e�9Q7�h����k�&���N���G'� �ʿU���Q�]� ,��,䒜�x(^��$�d�ƽ<�+�(e�_�=1@���8���7�(	���>����ݑ
%�'J7�ݳ�m���k�1=���Q�(6��&0:��9f��|�$H�-��|4�BN��,ER�;�;Į/�t�x�����0�K�w���Q�g��N���.AZ������Ja���$L)�PڗN�����[��+F9�C0A��%y9�cJ��'���;�ios1�|���~��zXN�B<4Z3���"�o�;���S�����]7���O|�Yo|��\��KM���c,9��q����g�1�n��)�*�v���0�]Xm�w^_D�0������Flt�X���g��0.��rȁnAL��jD�_�&"ȭ�I�j ɸG/tfj���׈(�e�+A����Z�ZO:��d/���sb�͝�:�\ԯ��T�H)Kp��~�w�0��hK�Dj��ܹWl(����`���>��@}���0ͤ�51�d��zO�8*�?Hz���6D�\�7u�����
�᠌�������d�mK���v�� �r�l����p}� GY���",��s�oU�np���:(�`Nd-�)���hV���)�����tR��4��B�
���Y�%��N:
��?h���q-���ZB�'�1�v�����yE->K�O��_F+v�N��6�ao�T��Q���_~8q2Հ�����^��4����dl��t.�#	[�V$��{5��Չ��F�ʦZF�g�q�K<$莭&7j2��V�ud�5��s���V{�"�mH��A�z;�C����$�0-�l���miOS�$JPk2G��s��ci�%m��\�;��rq5�y�To���dkP����?sEL�-��;Q�Xཊ_�����e�rR���S�8����z�q��G����7���7�K5�:UreKrn��t�a��Q4R�0�ʰMH[�玵5Ì�"ů]9lBm�!�N�+�p���'����Q^2���T�	��l�7vE�N
fCD�;2�:�����D=ݰ#ٞ��1��,���J�N�ҤU��B��M� Ǚ��t
�9֪4M�e�c�o��U�����j ���M�YG�Y_C+�w����r���l4JF��f{Ň��Bڐ�BN�ݯ:}k?+�f�^�+T��Y2����PG�%�y V�"��D�1�GO�X�,�q�U�E��WT��d��9�I�<��C��S��A=�B��� ���i�}�z�%@"��f�BR�6*�/G����8L8��9�.S��|6�ASӲ9�mܧ��^�nj`���׆,�[� :�(����N�W�8����nU?�c�H'�bm,<쪚��6��$6�p�'�h���(L������D�S�Bv�ώn���2�M����˛�?N�����Q�u�$�K�\�G�N����n1��1�y�UѮ}���;�ʈpNf|4���`������n�
L lQ-ݥ�e�q���gЇ/�o&R\�����u|��P}G�_ݳ\�g~�ip:׎��WǷ��2�?�TØB�{-bچ�4�/��-cIA�mm�9:
&r��=���.�A���\��܉C��ƚ �M�����kص5|�m�2
j�)�؈�W���J>�KW�_
*�����mڶޚ@[�����`/߈�v����b�i�u�H#��+gd�������kR|V�>��[�n�g��[!�e����3�+�X���jԁ���h��JR��⧕��)�ɋ�G�w.���{:'�A��
��<	P���H��Wl*��qK�)L�����Q<�	ZH&ە�OT5�U�swӌnT;-"�w��=���6*"���	Ct�C!%�-U�9qҜ��<5i�mź��q�RӔ�d�B����vo�G��'���7��Cq��o<��	���K�+����"Fg�R�`�&����V8)ye�r k^]u��SW����%��wY�f�X�x�7�Ԃ����.Z��Rع%��%�@����{�-�'���5�& D�(9k˰�v`����1\�Bh��vF�֟�Nw���=XK�Q��k�0��q�w�g�>�a!�jȻ�~?y�̸\��嚊�4"Y���뷖K�>�"rdjX�����0�(ʷdɳހ��t�*��ܺ��`^����E�Q#�vgA9������ַN6B���9��J���X�C ��v��)6��ACCe�2��n�0F����@_�0���0��K�"���;/����XH��ӫVIK�o���#�?��bQ�[
���.1����"�-��;s�5B���w��
�{՞d��xlΊ�ձ�[u����{y�]�u�[l�g����w�Ӌ������+b�U9)Ǟ���4�����X�I	�]O^���p��2��	E����P���B�nyj�.럋(x���~��Ғ\>%�Z��ݼ�8G 5��KV���S~#��<R���R{��8��|�J$cGT�m��b�y�
�N2��p�'ݬ'�rsi�q��0�58h�e�N��;#E}̊��>!c@������f�<�8��y����Q<�o:^���%/)���z��Q��A2�X/���`�F������ɽȸ�"!�r�/R���e�4u�2"���	�WvX�^�Bk0��)�1�K�Y?G��|��WĪ{*y���`9H��t�ţ�����r��u���[}�0А�L���fZg�՚ �P�[�&�C�J��Ae����Rǖu"����V�~����;�� �&F���rc&���a����ㇳL�m���'��Ȕ|/l�I�����=�S���Ta.ׂ�u>�3'u�y�^~�G���#�C��ȉ5th/���BDK���Ѻ��U���e���Ӱ��B������XAG5�8N�H�eg5�����������H-�
�P/��&�]C�	Eۡ��o����{.��^=vt��������! pl_��s��r�Q�-��1h#�o=�X�l1�������/C��A�Rn����r�
w]�k*Q�gZ��K��}6�+:��KJ�`�8��g�N�:��u���H���~y�/Q���{���9'z9:�H��+�����i�m��sk�{���􍅞�����_l�M�sg̳ߵֳ3v��h�#V0S���1���c(�`%�_���v���ŗ��]�~3�@��ꂻ��!�z!�W4=q���v��\��j��\v�3�����+#!Q��}��>Ŭ'y��b��$��ZX�jТ�6�����F.᡼�.]H�:kn�@��W�()!#��@w]G�����
��>�2����dE�E�zE�S�����v��^���segǦ2"��5�C�@�^�G\�I}9�!�1�n��	{a�?qJt�&��ˠi���@���i�N����|8��m0lK8�*�L�udOT-*|q��ƌ����F{������1/l/����`K�[A�j������g\` ��/C36������"��j�%�[��;J��[��u, �A��\���T�G�Mܭ?㐉Ek�@�c����)��쮬�,����p�V-�a�������HP�̥�*>C$#t��Bչ���S��*Y�~�kX� Q3�*	��-i֒�("���X��}�dN�O���y:�F�|1M �V5���hh3FV����,b��兒�>��ye���j���"�$:I�=���zTڇQfCjY���ڊU�S��GZ�.��X�	8n��OK������eϦ'3!�/p�]X�P�D��\�/?[�`�������;��2�kK����s����2IV.e@�T3u� ���f}����Ō�4I/���#IZb�=�``$`2ҁ�q%@/������}�:��'���Ŕ[�MG��m�>e����='���z<	ޖ�b0@��鳦������օ��q�|�r��E�`���,�p�{��޿�q�^��N�:f)�!��dw�"�*�l�vJ��3�Fv�4���%��9H�s�ث(^.��ٻe���]��Q$��p�BG�Fq`WT�zc@�!NƉ%|����;��|,��X<���V�̈Q�L�(Wchg��ֵ>k�?�yKI�S������4fHb�Z�|ψ�#ȾYz?���)zQ8��3�+�)T!��;��%l����h�`I�c�m�b�z9��І\\Eۗ�h�����o�+�W�6�luoۋMvw?h���b�7���-��l (i�5d�+q��e�BW�*�f��ҟ��_ܻ��7xl��m��*U��:�7' Bщ��=\�X�����U416��vw�4�1��	A�A���� �e8�@Q-��E��0Ip^�u��'��M@�f����'<� �/�^�����sFF�+�q�*awCV2��ٛǔwA�Minu+k�
#u!
�Pܟ{���a�>�v �G;肜%I|y$��n	�w�7q§?e�ig7�=3�*PB�&>��G�^���U�s%n���+�W�����ݦ)�WP*��YlW݌�P�<�2��Y�Ö_��Lqy���o\̇����0�U+�=�u�Uk�{��)���H~{:s��s�`Sm��˰� ��5��!�6sЖZ4ɰ��2c�h���<��-�g=S�6����y4RX*)�^�{�b8�6��>��/"�\��CV�|q	n
%-j<�t�XӦ������X�K��N�FU��L)Y��r$f��D�~OQ-�͎�c��S��y]�l��@j��w)}j���x}t8�>U�i`T�2�lI��N����4ws��Վ<Ѩ�M�c�/���7�f�*����8��}`u�T�)s»leUt�F�S�٤�e���hB�HU�v��X��
��$<��O�?��DV��今7s6�ӠP�/@��EL�=y��i47�@�E�e�O�^:w�u�9�΂�2��0�t��ҵv�9C�7�;c����*`y����J��]��V�Oz�,�䅙F���ҋN#�h�<h���ҹG'V���Ь�e���%�ޒ�*ܹ�+3�o�A���n�>3u ����+#�!�AHc��T�O��m�y$ʍTD�S�9s]]Gfp��l���{�.���|d����42�/B>7��;�}�OS�^T"/�H)>����Q��"�#�1��	Q�tK a1>O���z���,�翭Z����{	���W�B��P0�"�f�Zh���#��fX�o�CX�c�?L�VS%t'�H�l�87���IV���D���5�=�+�w�厸�tp�X��o�t[�c����%�S�Squ��:�����.adӑ:��4��w���)���e�!��v��HH����J�T&\!)�%!婎�m�v+�\g-�:�4:�Ȩ>��4�W��ىCs�a��S�*�ь'�i�H~�����ٞ�>�x�Nmӄ��:]z{k�S�e�T�a�A`G�ً]�z��k+��L,β;�H���ן/֝�����/ۃ�<���&v�N�u� 9iԤ�A�������9 �2����ك���'xq�*u�9l+�w�F��3�Bl�	�4T�Ĺ�%�C���L�4���}�K���S�􊀠!�Тs�Ы!��l�6M/�`� ����P���
��թCz�D�y ��A���<JCۥ$�b��D��c�w�z��R$��&��&������.� �t*��x�謩�v� #w�|n=�|� u'� J�X�,����JtmX~;��m�;ui{�]E�*�!;���t	�5���Fa N��)�haR��t.�5��*f��l(�������ɰ�w�'�1e��	�X}����o�%6�x`ꦄC��K�}�'(�Z�l�B6��2-����x>��.	��������|d��gr�HU�邭-�g���
�f��"=:�G@�ȼd&%��ϊ&�"%Nh���$�_��3`�λ��HK"�����HAt~)0薪D]>�,, .�_Ŗ��b�؀{���:�`U%وh��D�����0�[8݂Ǔ�Z�.M�F��b�iD�����q}�5Ҳ��̯4G�f�h>ͧ+)2{hЖ򲔄��nkރ��'w����|1���˱��Mq�	Լa`�zP��s�X��5oNߜ��d�wScc�P��#S���j���j���K:�B�b+��ұ{�)�Z�<j'�R��mU���ppO�-U�I&B�u:\A�Qp r�&:�F2�Z���Ah�]�v�l�3i��>ɮ�E�t����vV�gG�}'��Z/��V��04�p����٭:pV���Z߯�W|*6c���Z`����,>`�ar��uw�l�=a)i�0��PcN��@��BΉ�8kn�T-2���y#���k���׉�\(����M�9