��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E����pbT6o2D�&���6͓ț�W�Ƶ.�=�m�B�Z"��I����	P��sfs���e0��ۺ����u(pp�B�M�}%��,��Y�i��x%Y#g�淎+	a������v���nR�}����cK�.E�&�(v��s]�?��y؋�UiC�M�?o�r����Ȇ�.�:�}��DEf<wI;��h�M����z��GϜ��ˀ��ӎ���г�K�w;1)��{��16}Ѡ�ȃ}p���D�x��x	�B��t�|�����f�4_�F����_ ���40��qYDl��Ճ� �5ލ��GN:ۓ���D�9�j�P�"H�<�郎�dj�kb�@	F:V\z�7r�'��tS�PZOH�M'/9cy&���.�Vu������&����ѣ"�:Z���R .���u�H9z��� E-�-����o6H�⣏�j���ק,e/#*�i8l{�5�yC��8c�e�^��']v�鋶�,-��H~��Yg�8�m���c�=1���j��H����� �����W�3���Uŏ���}�D#\F�����xM�s&$yï)�?��9VfMkn.Wo��<F>
�4���A��������rp����a�tS
'��;�Oʃˉ�W�c)�O�5~g��c�t�pmu��5��J>� �~oz�q:Mj }ں�%�g_���������g�U�\GN��
Uo�)��/T��� -���Q�օr	A���h_ኤ)(�
�� �=P�;���:��MqǮX$�~x��2�4��ːs���=v�\�9|��R�8-IDJ����Y�:�S`��ÑzTeR�U���M&�& ��zF'}��)�=�I�H&�|��W����Gmͪpp8b5���8�͹jVds�����gݥ��
��s\D�ľ�0��y�]�W�F���qM��s�6+�j�M<��4�H���kE=0�#�ǁ!�v�Q�[���1�c�A;�;�K�.(d�Fʐ5��2�K��/)VC�nԽ����o��~�\������r�)y��M�BE�j^w�@���� >ts�K�,��R.�^y,U���Ʊ����2���m�:U���_�s8g=A���D^�p�i��\
������y�D	�V�h4WS����A�֪?n=֥.�(I��`G�å2�V�,�inc���x����Ƥ��=KZ�7k����6C�Ç�ԩн֑N!���4F:p>���c�4c&�]��Vуpe���E���H�`]O�<�����+�X��2e��{�[��ӞT0�J�Pt�Sm��E�c���bBJ9:[�`-��[=�Y�鐞���z�b����� ���\R�,M/ɧ�3�[��Q�����&��P���x�Ia����z:q����ݖJS�ԓ��l}�J�*X�%�y[4/A	a���<0��?z�Ņ��ɮ��R�7-�̶0-�HF��ע��
J�[L��-�!���ɽ��sR1�7O���8x�M�y�3t�d�ļY�T.��Lt��]����^��3����Ty��^��R�
�ئfe�a,"�3|��.��d�q-3�VD���Eq���Ф��Gf7��ux��|�C�D}�E�7?����u�أdX�WTzت���,�wg;N\Ø\��`��x�dћ�4����|������t!D�
g�t��ʝ�[�'�7���q�Q�ё���l���%K�P�B�&\9-�E�G��=(?�ON��o;��]�t�zZ�=8
��9�����a;�v1�$t���bf/Ҙ��h�@�V��N@*p�f�4�9��ćmc���˵e��K�<�`%�d,"���x+�G�ǉb�"�󢗔�!p�1D/�9-q���u��Jא(��-E����)$�CJ�7��咺���'��V���?���FH�����Nį0�T�)��iv�t�� Ka�=��>p�_�ƌ��x��|d~/��sB ��)��JJT�A�\r�n�M��\�OsK7�����Z#G�B��\;OL�"��ee�QV��gӉD����q#��H����ڭ��|7��Z�:Cڔ�dQ)���6(���Y\3������
Z��@�x�E1��֪�ϛ�^D��-��M�2��.TLvd��͔���tiV���������<[�w+hсζs��.P�c5�O$��ɤ�}g��@���؁|W��]T�O��؆L|8�����WD�:#��o������;E�i"�YWm�o�-'Wu�!�(�߼n������^+C��xVV�kUV�"�A��g�6�/��HWlD�=��t�. ��w����/��w�{l�Pk�,:k.t����6 ���A�7y��T�d��8ʏ�*>)�do�}�qvPR�Y�bh��TF�a!�Oi=z��9o�/��0�&�C A��ӏ1W��u��G���2��C��sk��r���.@�@��s >���6�^�Bί̆̉S�Q��ܪ0.�\���櫌�+�����a�+�LzSn�a�Rb�3 ��j�&�Av�}f@
#��F#Q]��:H[Gj;�I�m����O�{[Ь`U'��ݧ��jԯ3F�n����xC�M��ͻ"��.ċ΂�,'%ڮz��%� ����By?s�8	����e�b�&@�3���c㤸����<k�fii���V+��
�>Z�=�kK�u������s�v������ʾ���>~���yM��7���0��t� S�Ʌm��&���,���Q�d��Ʈ���8s*_�bhq]�ǥ}�Y��R
hr�e�z\�`7;��7[p7\k��U�>W�9
7^�v��낸�%�;{�D;���U�w������I�ǂ��[?���p5]���	��ǜ*ў|Ξ��2v\���|Ԯ]�!�-e|�������r�%<���(����qNhk~���ݪ!�<Y��e�{<��б��T��]�$�Ш�&w�a	
���~<ɺ �T���{��uP�;� �0��8���یw���&6p�L��8���'��x�ɯfk�âs��O|G2}�Eh���s�n�N���$I����^fh�@@�zC��,�����T�������]\��Y�HPX/L�HۖH��	�U[K����W��N���G�Ҟ|V�k{fB	aQR�����j}+�l���^ZMo��}XJ-BJ�q���X��K����4� ��\�3kT��y�]����H`C�^F�{W���p�~ì0{]Y:ÿ!_÷�i��?F�޺Թh+������Q�ޤ��lYq1�{z�l��~���|k�c�c���(�KFI�w:�.t�p��p�3d�SG]�g�}���L@dp��,������'�Ö��&���d0�)��r�KX8߬S��Z^�.���Ln��Ų����"7/-fi	�����Gw*��>!��`k�l|
�.������(�vGl�A[Pxs��mʐ�`^����Q���;i�O����|����_���Z6Z?*\��""u1S�QY��8_�'h��YW0T�\bGs��2Od�w�����Ǫ�9d�|\DB�v#�f�3�{K��s����	����tȋ!aYΏ�����x��~
�Zi�}YVC<v�*�-�ؾ(�Έ*/�F�sSkd�Ȓ�R����"Ume�=���$��xa�/b��nOZb�ס\��f(j5#M��~S�Hb�����r�&�����~R�������c�q�ѮK� ��nL�����d{4>��Qσ���G�
F�?Uir���c~��QI��< k渙l���~ܚ,��yQ��A�B����o�)[���}Kc�AiD��9�� M��a����u]$.5s _Q���v��.;dp]�uv}�����
pxqQ�P��,�/��v��U��ʘ���g���l^����)�ҠWYu��mJ��ؙ�p�{4X������v�}�H�W�S�	8a�������!�9So^��r\D� Q��v���J��ʮ��_{xlB��d?�Uܪ aгz������#��M߷�!@0L�D=�.���K<�������/d4���"����&��x�5!
\VO��|��$����g��9�3^Գ�ح�!/��ܑFZf��w2��=A��_�/�r�Wr�@��oh�`mE�i�J�$��v�SG��*��B�����r���0�g	Kͩ�%����L�,�Hu��/�u$�bv������m���\AW�����������
�E`�����K0��9i��j�>�+�H�ɱq����τ\C��F5-�񬚭@����@�1m�eSE��e
�g�'Ϥ���я�z�y�(�<�����M� �)��Y�q��Վ���
a;�,�Nn2OAm���q�'bgH;\����F��I���-�4_�{]1O�m���^��1Q��%ǃR�Y��k���,=��l(������'� gL2%0��y^b��UE"*��W�h�f%��.q���m�Mz��L嶮�(��+s{b�ʉ��z{���w`\�8�j�BUn�!&'7?��^���z�~����F-����yX ަ�,7�ʢT/_�g��7�����L�u|j�"CXZf��t���*�7]��u��T֩�j%�>̇	��(�-½�)vs���E�0V�ٟ���%�����CR{Ŷ��I�رR4�
��
����L����-�T-	9^��i�G��w�GPx��ڶ��y�p$�=�b��&0��jc�����{"�{D��h��C��"���k�ʿ���[��=��Vw����J^5r鴪��U����z�a8�eAsG���ϧ38?���.!�-�Ʃ'�82s̏T�%!r/݁"k��_d�R�b�Z(t�xMM�x��C:,�l�)vY%7.��=���)g:�Q\ś�\��s�zнW�I���L���ޒ�=r���z�F�ίqh���Z�~B��M�f�x\�P�7P���kڇ�j�>�<�0{������G�c�P�ML3_�7@��JUX1�����-�wɲʃRo�U����(��eC7c�﹭�|R��7N^w� �5 �Je��Z|:9�r��vڨ�����0�Q�'V ��qk�6]�B`%}���r������4�e�@�����U(�Pc�tL�J��� CS���jr8�u�0�C�]j���9�yo\�Ǧ�]pB��W�R�7�f�IH��JR7Bv�F�*Ex��sT����ækN���������.V�� W?Ńˎ�D�p����J�����eN�3��R����uq�*���F�p`S��Z���k�2 ��x_���D��KTG�������,C
/R��ө�fV��:���WN�mM�9��a�z�fu��fX�wNIH<��>^�C,9[�q�V�����
����a�vӲ�Ixrb�����,�k��;�~m���1=s�-�i���u�E�A�}�Ho���/(u�!����b��2�b1Z9\5-	��v�!e?�:a�z~c�ndd�x?���pk���6/�4Y���W5fߐ�q?.��X��������q�������Q��h�/�4v.�1�]��v#�׽�}�rG�Q�^����ɽ��1�&�&�Z�z*<�~�2� ���\u	\�y�p�4�r,^���V���da�����P��w��^���P�y�{�f�>��`�-O|I��g���:+w<�'�_^(�&xq�,o,��*�8�!���t�:˙q)��A���e��U;��nqV��v�q[<>3�&��o��o�����g" ���2�Q���Np\��g��5�*5��F�U�����k�z�GYT����K��	�>P��	��Y�//���@3�>]F
��K=��ڼ���y�jf#ʝ�H�3�����|'���(a��G���X0��HB�ۦ��cá���h����e���о�����N�_��	�E'9��L#���=�j���� TͺO��h����|n�����2��	&g�1�l�ǈ�����<��&)���e�X�5��#���I����N��W�Ϸ�&&���n�,C�~�D�w���cdd�y�J���3wv�cS5.�>�r&�RZx*�����>�� �rX8I_;0�O���c���d�y� v�m��T�G�"��b��MM�插؅s�VA}�M��ր��n��c�8'���~5�]��غ��Y���/mj�����	�%���Vp�Y��U5��$]/��0q��[����t��O)ː�S�����L���e�� +���p��� ^��0�-��XT�Y�d��@&�����H����X���I݋��6�d� ��UAs���R��$�%�%��_�$�&Dt��;���U:���s(���,zX��!��wN�������|���waDT��,Y�p��QQl���:k��57]�>ْ����$�HT����͸ŃZ[��V�$�~�A%���9�k��7V��p����,� ��|o2~�}�yC����g7�0Ik�����:I�GGnO�.Ln��k^mD���g'��7�a���T�f��"���~'���}�K *B'�X#����M~d��W�s��."��\:��5����Q$�����T,b�
=8dF�
-�������v��(e�ϰ�W��:f'�>�CT|G|;���5���͹�C �e��ˁ4�
=#�
� �fѹZ�-kZ�9��5�8��� >�GeEܒ��e���/fZ��<�z����3���/�I--��ֳݭ�x4om~'�q�tq#!�5S�67����3(��K�;\������d欕0>�9��o�9��J�ͲQ|��b��b$`�0e	����"mTn+9e��7i�$��mȘЩa~(l�)*�cZ�* �k��;@4C��h�Gt�n^�~,��[%���/���Ӎ	{Z	֤al٭^�<h ����P� �ӫ�"�M�̻do�]��O���g�5U��%����b�=���N��� �ɚ�&?�������Ȕ}�������d��Q��(�9l�X��u}�����E���4i�U#��w#�of�rAUS@�9&8����
M̞�*nU�r���Q(T��;) �J���d*<!'L���tl��w�,�����q�l��φ:U��v�\<�j���\l'�9]p�2p�5� EHC�:��F҇L�U��7:���Vqy�9��U��!}�=e��R|�%��I�߯�
(~�N����F�V�]i��e���5�!��_�ھ2�7<�?d�`�1%M(&�qV�끲!��.�a;7*Z �B�7�|?#�Q@=�$kO���<3!0)���~�5#�י���}��tøuBߪd�뾅�ub������Z�3u� b`�������:�xM�6�O���σ�i~K���񤷼b�?@�k�tڽ�f�2���d�3��^k| ��G�:c����͕���p<��U�w�5�o
�A{a!_�88�GƦ*��$-V2֖Yn���c�$����ځ��
�ة���ܯ��d(����{���O�YG�b�tǱz��r|Pgo�Ǩ�f���uԤ�jN�eJ�Ȉi���WEgI�&MA�k��ɭ·�v�����n��sy$^q����ď����_�)�m�u��L�r�J8+���6N�����*t��ĪR8�^(�k������Li��:�ℱ�����2M�1I$��ƍ��8������Yj�{��F��pZ$�B#��&��]��K���g�؆��^��6.�riU>�ı��E관�r��T�G|ktc�b������]�t% j2��n�{��n�#<�7��l�5�݌����(��K58z�L��ȶkf-�`!�~3Y."����&����Z���π�g��O�|<�z& ��^��M
Ϫ�/B�O�w:��}��9_�W���� :^*/{B�LF��R�p�ߞa��_�"�����V��+!��b�w�}����nGf�>������h�rߕ�N?��s��+xz�����N�-i�w��[;>z ��g��"�&����L�u�Ѵ�e��jE>IAG�a
�W��y��NF���唨P�)ݶ���(�'���gQ���=��_5?[��i�0�;����٫00��y����*h.�����#R,��z�����M�f�r�@A%4�T1����J���y���pZg"���ͼ5U����U��ƍ }�GT���̟o�vi��z6����?Q�S��j���H%6�룒��y,�e�u#
���y��w'0<�ڍ�L��H��5`Rp�V9�l���B��g�j�k�����4���:A���u��#)x`GےR�q����������dA3)���%��ݷc�.����2�7���$#�U���qut��(�R�^=/�@���;�Z�1;����]C��Vo����*	 ^d?��w�5S��ݏ�aڜ��ze�51�|��!�l(Vp����:U�e��>�}�%����kB�a����8u���O������N�a������G6_r��߭��'��>s�ӻ�D�_�K����=������$9h�M�ȵ;�c3K(�b��- ��&�>�v�Ae�ǻ<����'�pY��Mh;��'��V�(}4�D��q\�-��ݢ�|paߎ�ƒ��� �u�f���SS�)q���t�����v�vާ�\Lkmb��*�Px�+K$XHU�Sn��';X5�nާ>2�l'^���X]ݱ���<r!n��,x �����=�>4����c�lgG��/���b��& @����C�\�E'l�W86�15D[�����͠�֡�.W�7Σ���V�~��V��'d� ]�1a�;$F������2�+�-'L�tc����q�q�[њ��F�]��P8���s2���*�m���K��eĦ΋GPr�7V�1���. ����.
y��s�dF;���U4�����-��������1���"dcK��<��}}��U��:�-h�&9~�ȍ�1:��4� "���ٙL�<O�I���\��K-��0��eROǂ�}C�k�"��W�/��k� ��`T��K-R�RW�biGGP�1ŏ�b̅�ni���;S���STғ+���Y��[JC���џI�ѽ$����s�j\��J�Q��G�ь��y_Y�&FЬ�H�<J�ixw�:A㦬�5���_<���w��%��8Նۣ����k��nI�ʈ��'g��/��EB8^��Y�3��}�z�㡤/vG��M^��D�%^���Hr�Pګ�"�胋��;2���$�Ϯ�w�V�QZ�)��6^{Q3���
 |���I)Yg�p��̕~:#	%p�=�1�oni��h��/�Ch�9m?n�ƴ2`��'iݜC�D�$	n�D!I鐂�KX�H��F{���������'����7��0w�d�/���I>����^e��G��	���_I���˚�n���z�Ko�7�������p3��MtlE������� 2����m}�>���`俟�����F�7����,	��d^ǵ���e�	_�ԍ��t�j��D���NW;9�՜��*x '�tpEx�[�*��F�1���.��P��X>M�R��N�r1�#V2�m߰�q�UN03g\��@:Z��c̗�s�.�b�ۇVi|
�ߍ!N��#t��5*?[�n�R���!UU���ŹXW��ym�a:1����Kx���!#�5M�/�����s�Z�7k�T}�Cf�l��W^mq��sSM�w_� &�������O�Mv-1r
��u7��-�:=8��
A>k��yƫm��?���MC�I�
<��k1��彺~�C���� ���$4R��B3�C��>�p��:7xsi'G�S�wޫ��4�^�$���Z	m �R<�����*`�,}��R���M��VY-ס�3�yU�$u�e��7`����pm�ۃ��ŷ!5.Zd�H�����<��ވyKg(����8Gɼ$.d}�V�&�N՜��Ҩw>�Yx�壘�Eq��'E~iY�@3�]w{��-Kwl�\9��b����x� ��@�o���4�X��)F���w��GI�)S;�7[�MqB2|w�Uo���竣P],o�������aH2����V�\�/ʰ<�D�冀���b��gS,�POEmٓK�e1��)���r��O�@�
m�]d��h��(,��n\}�$H�	C�U�!M5VK��_[_�p�1��7�I��昊J>'�m��	R���vı�����`=1h���x��\䂱o���.�U�^�xϽ��!����\�n�sd��2�����A��#�xA˱��l9ğy�D6:���I��ʽ��>B��4�J�x�,ۚ�_�Y��y�����^��X��r�tw����p&YD\ Y�o?l��@Y&��TԈy�LE��vxs�w�ɦ���m`ؙ�nD�㲴�W�w��i�f����	������m�=D���L�B?L���p��y	J�]�b܈��UQ�n��g��qI� �a�^�Ğ��G	����ǔ����k�I=���� qK����rNy4�K)�Q���FoH�22�k�R0�Bƫ�4����{�"��|�r,)��{�/�v^1�m�4� ���b�"��T��)�4+���=U��#�n��g�n�P��lPPS�����K!�ʱ����,�ԗ�x�ͫʦM�Wڨ���w0��0��C]﷥f���X|����\��_F��'�.�@�t�>0���i�W+4�y��o��b��l��NV���=fq�jF�ů�tK�Ӝ$���/�{Y���ڪ��d	��4�X��fwk�u��r?W7�ƻ��n��ht�+6����К/��xK\1j�@��'<b��`���\ԗ�@nTD��;�1���!��t��5�ze�;�9t��A����k�<�w�>{��:�EG���=ǯu���N��]5P�%�m�w�^0D�[��Wi�v4�VHt?(S0!~���O������ɳ���j#P�(q��!Q����K�^��P��K'����X�zΐ�N��o�?�$���,`�v🖿����;�E�{�z�e�@S^cD�h����/�Q��?��?p^T��Æ���o(���2����P�B�i[,�E�[p�-�����uK���sH[
U�h�}9huV��c�j�tZ����w��ũ�[y�l��X��}����ޘ�T�,�[=(+}oo�4�EB�gw���l%[s�ls_ޏ��4�z���1C��B���_xWԒ�0�o��"5�~b���\����e/��ߜ,���5d�-�,ݷ��@�]T���|����rե���E�Ң�ت���uU� ��';��)g���6���z����CWύ_4�C�DV�;�Z�Y.~���\J%N��P���$��|���cc��0�T�?w��AנR���6�6���9ĸ�!�O��ז-J]���,�	䠛��ٳAK{��@��Wc�hԩ��?����:��3۽���L�$�#��i4)�?j�c�ov��c>"�v��G���:���q-b��'7��c#���<:o%��;�S�땺���z��:����p,��#���v�Z$�R0Ib�>���A�s!� ,[�!#��0��.���A-�MՅ�=b�%�A�Ȅ��О�<����@s:�0y%�l������7�b��~�Xs��ШZ85�W��KY���z�Q����� �l2g�fb���_n,���~�W���v�-�˜��%hN{�G9@kC�<ͷ����F�8��g�X�5�x$��a �	t���]-�@�����`E�%�R�����ۘ'
n'OGC�+�I����f��6[?�@R��Z���N:7���P���Zmb�0tͩ�T�v?�B��߆U�q�l5G3$%�{�0��m󱝄�S;>�쟶�j\0�U�h��5ӐYG�׿%�A\\�ɉ@�&e���1������@}0y�a;/�p���>N��T"�f�c��o�waަ����}�j�;���=n����W�~Y������cV\�0`�:y��h���2M	��I7&(�(OЭ6��.������v��D�R
�z=MS����ʤ�z
�*R֊��;�-�,���1��[��$��Ⲯ����ntR�����ڭ���-�G�B&��E�v�
e(k�P�͑<�'7++kJ6Lx�����u�����}��ֻ9~� �*%T��¢w�R�Q��խ�ޑ�u3� -�C�9�E#�h
RW�� ��,�Ӟ�>�'gϢ�����=S��.jÍ�B��a�2��+-��������-e�j��a�LH���+�&Z�t+�/<�F��heb2��z�#��� DlY�N'��$���3��NX��qs])t���Vw�_v`��K�{(�����]O�C�%sRϳ�է@��S���'����g��J��= �c�[c�
�e8���||�6�����1���|���>J���p ���I���E��NU��zH��B��qe�^3ޮ.�ݧ�TWan�� ���5^� ����]-����q��иu�_p����O-��l5����%�o�g0tV�yXb~�2$ۖ�zt����i��Rߴ%3���X�F��NOv�Q ~*��꺮=����0{79ݒߘ�L�7������⸟l�8����<�+aq�L�`3�-3�����|�Gn.�xT_<��I8T8��W�u��FHkωi��xo$���[̡ <�#ڪE�cM���������bX��D9�>�k���
�d��U�~�Oz�V,�w�6W<q-��pe~�t�i��F��/q������A>���kh���l-C3J�9���ȑ\*�C,�)"N������^�84P{
�L��u�x��o4��i�D �Ć���M���t�܏͜�����R-mi���@w���w�s�0o�R�2�@���+���3]
#��5��۩����`eA�WR�h�N� �V���9�����B��:���ۛ2r��}���yH��W��1��6+E�SV+&��;��pkP�q�>c�X#��g@�:"@�%[qs4�����x��Jr�W�a��X�2�聠��VP�zM
�1��V�;잗K�MM�����c��~��ՐQ��)�]Aw��>���AA"Z�e�W��U������2�D�R��~D]��ҖSĩ���b�������	*q@��b1I����b�aC��r��A��O)�����HA�1������L�8�q.6�W��]�6k�0���9��|-�3�� ���j�ju�ʎT�����<w�:�D�wd�|2�:(Ҕ���u��iL��n�g����њ��yTc���l8�7�;m/��1�� q���*6�%�M��V�D���~%j(�Mvē笢�{�M��E�fMpq�7��UCBTf�OU�r���x�>A|��Qm{�B!��'j�)��2#O���i�_Qܚ"����`�[N׵ E
�6���K�@�G���-�� )8LBU��K"���FK�WȠ郍��C���_��&N������'7�g_��_��i}�^j���3j�#�eywt�i�G���/w;k��k­�a��|�R,�p��vUh(�����e4�R�r��M�Ё�+Ą�_�[�_O9c�m���m3'n1��}�,�O^Њ�*��2�Υ^^�\ܼ�/K����nNN���Ln�L�N�1�P6�4oH��Y#%�D��6pn�=�P��:p�A�J|LSH�{��;Hͪ�7zycq�tT3�釵ʟ :@��`���vMC����S��>m%�r�\�u���q���.�]�+���B�lj�5�V`̔��z<1N]8�D��l?�K�_�-�⥌Vg��ow�e���#�'���6jH�T)�M�8CY���ȎU*��֥r4�D��?����4Pp�y�Y�Axi�<r���.3Κ/g(�+zX`_��.���Rױ~��� ��g��Tvq	�r���쒿i���(s5)[���ty!f*��R�.�(~�ggP��)T�e��%A��V��}fiK__s?՚2`h|��I�nB
�pxbX��~��ݑڝ�To���ǀ!<�O���������(#���ʩ�&��+c��I�08׶�;*��{
/�/r��jyO\�o �yj4٭�1�w�fgoZ�2f��'z�2T\ېx�ג�����΅�) f��8_�K7�H����D��-x�D�,[�p�@�j D�I gcN�x��1X�Ы��-����J�7C26]��C�..G]?:f��|�5(��w����]E�<�n�X�Au����yv����8�9��1��D�^�sOn�R<6��1��v0��ב����§|�ltZ!��kR$&���Z�)�Ud����0,T�d��K������~�P����d���U�8�s�7>���gG%��x�l3i���fPb���Vϙ7�z�{�|���\<}Mzs��O`2hpgު��~�/_�%,m��W8�Z�K��P���w+��M�1JC���Q��h:{��@���:�����t�HGl\�j�=u�9�5��=���4��{J���;�c�o���2JSCO�.2j~�[\�M
���Х�.I�0��l���wG��̒,%�]��4����A�!2N��X^3�iJ߄8�o�I��lmTj����ɔ�!��-��5>g����`�I��V��t�N�1��S����v�гnT?%�{�c���^id�E���*c����6���Q,���y�ӷo�@%ݗ-�]l�u�����d�z�H�%�Xz���:Y�Q��6a����mX��`�l����"���6�}a�I+�����:�²x�s�Çǚ��ę�,�O����?��ᩚt�ݙ㹅Rc��aB��Q���}լ��!�5���GIB��kGѕ�41&�\jȣj�O�oˠ������^H����^��	~KI�'�F;O�z��E��%#Βݜ���Dz��KR�z�n���*Ʋ���:��ߑVp�A�kӀ�i�Z��.�'ڟ��Y�g|��oz�$h���^��w֩3�DՊ㳛W;}��+�Z8�B���@����Mmy���ы�K��^pà�yNQ�z���k���ٸ*!<c�3"e��8\r��7
QͲ�5�t���T Y|�F �T(��c��9�tc��T�6��3��<�����[!kr�#x'�0I�0��C��S��mh@�5$��>��9|7��R�R)0��፯j��U�����"�֞W�'=p�h\�m|�:�Ga�Ӿ ��8�+C���3�|J�oz���û�-8���t�T?��[Q��be�Oʔ�����cHx�O~�.S ������>�<����\�(mzW̄�V޳=+o��Ť�JgGx�X����Z[PT�+���y�{��3*$�Gl��aoX������}��wL���H�o�{��Xj	����� �k�ZЄe�bv2ok�{�pV	�6�;� r��3��Ga]#kH�*3��b��2�;2�R�_-ֻ�T�ĸ���?���Y&(|��ah��+꘶7�8�q���8.�c�,ᬄ�ߓ��˦��n6]��OH:��O�3c�#&���rs�� �xs���?y�+<�g���W �9>7n��g�$��C�4+ݧ�\�qI�"�����3� �1�����u 6�k�&R�Q��^���0�pO.Z����r:�S��=��	��pSk;�a����/u�(���Y�>; 1��U5U�T�L3�)u⭟1�n�Ĭ%M��ϟ�#���G��/���� g�:A۶d���ƥg!�ynBV�C݌�B���չ�>��0�x�>)��΃�fI���Q�6_c50(+O!m\��Q'ؾ@| ��pD�'�& ���[Kׯ�2���Rｔ?�
��r���g
�^����U�8p��"�+�Fx����h�\�'�ۭ�t��mM�Q�E^��<�D����`t�����#n�}Z��-�EJmap��-@Ǿт����zS&81f�<��HǠ['�F0���'�c��M�2��\s���*��i|w���!�:* �cbG�*UN/�cUb�[��� �U˞��+q�ؗ�e*AϘ���o�;������r�˾����αhB�VT�P��HR�V����x!4���ȳ��^s�/R?�NT��^�S�~��[Q������ ��o"���ȐF���c�=���8δX%&�����rȑǥᒳm��D��)�g����eJ�n*��9ca�d�L� �W�����ɈN?��7a��q�L$�(�y���������'�����>� ���d7]�Q�O��������jh����mU�	�u�?=B�}�]��Qx�I�W^M���4�ѓ�*�$)�x%a�zt�PQ�XVqN-2��w-?��ZT�@�MF�
[ ��1��C�T�R�5_�5�Q-Z���F��-���52k�)R�����Y��˿���Q��ԜT�	8H�g;��-��1�d��9�Wmn�?��\�h�Dg`\��p�׵�zsF�C'`댤>7���f|@��~�{Ь��j��i�*L}J_g������B!���i����%8�_vL�GeuD�r�i];�����g��%]�ͤ X��