��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B��J��Ǯy{{͂�[��N��������]m�ˈ=g$k�n^v�{.��ʠ,�{������ld|N�u��v$�R�i�f�,Y���v��w@H�o�v�w[OC���UQI���&����RF�-�5_spU8��Ʊ���������k+�(��P�{e݅3�S��0��醆�a�p��ڧ{3�n	��?m*��uuTB���1����r-sG"ة��oE�P�pO����N��;woїc�	����aћ����#��,��O�����Vg��= v�ﴌo�ǭ/���9N�[��Xsr���%(Xy� C:>��o��*�c1x�͠�҈����������x1:���C��ɂ�a��ܱ�\���I���M����A �eNY#|d���������e�j'��k�X{�h�Eʐ��Fmg���b��p߲t5Y-輮�>�����c\Ӓ��=gʡ�Q�w�+q���7�� .[v�����������O������[ň�S��?�lYR����6�je��(��bD$Md^�$�����R�p��c��?]^�՞4�ǅ�2i|f�$��8A'c���wIu�\�'e�%�;���۾��2�h���o�E��LQښ�����OSH�],���`M�i^�GYrhg��~��Eg�Ra�z�����`�&񖹐�,�H��>���4�HQ
�����t��y�R�"�\�c�->C�P1�5���G���HiW��l¥jU�>�f�MJt���W�g��&~��,��7E[4�����#c��-�B�0��M��q3��D@ǅ��yB��5MA���L&�d�ܫ�>�}�k9}�F��53jfi�7�\��sQ�OKZ��F��nN��:�
�(������(w�@-�pN�<J�[;���W�a耽��������Ly3�'+R���Y�2����ZE�b� u�wX��%���[��J��HkA��Yl"a����9._RD~�տ
oҏD�t�y�K�#g��	���Re�N������s���:���	����9m��7��&Dn7��P�y���2��OH\�&�B�񜍼m�p�5U�������� �(���Ҋ�'M�3? �6�b4��)>�G�Y'�h��|�ͫ:��1�W�\Z��{�skQy6�x/;���n� $LmzO[�����d��p���q�6�(�$ʆ�L/|��Hɱ��v�C�Ռ�
�$�.8�ΘgP87f�9��(^���5U�x����ӤF�~�1���<O�{c��s�e���W���4O�B�`i���i�G~Wl�ʬ*�����a%/oϜل֎��
<7 �[�dN�=MNH�Q��HFs<�37�},B{b��LMX�V+�Z��4�\�>= �s���C���� `kWr��VM�?4d�ũ��.�[��!1삮szDK�2�N��=l+�|���&� �Q��a��%M&�犿�ݧ��w<�+R��M#ju+����p���P�Nu���� �({�qsC=�դr�������"1vv��~
^��+=��1O�&�/�h���O�76e��|�
�d�p'�S�GW��)?�G<������McVQG]�����9ƞ6������<����L}i~��5y��Dg�� �q�#<3��?�kT�M���mo�II�8gQB�k%
՟R��di!v+v |�� ~ƽI�Y'���I{���T�J,^���B&!���7�Hsyp���-)��K_��{}o|��Xu�ۖ��YM�j�k)9¾E!��L"�ԬwR$w+0k�^?�ϑ�t�3�<S�����秞�%ؚ��5��H,\�
1�����ȕn��a�A�lu���#��o��+5��� ��L����W��;-=���.�hP���l�^E&$ZӦbɧ����B0vҚE>�o��#oe���)�Lt��Bv�x�$v�-���Ɠ���Mٶ.��:�"cS�*�������g����b���c�ۦ����E��.�"6�'Y,��M!�����y���m 5aw�أ�%�ȢA���)`\	+��}�ѱ?K�^u���k��Zk�C^��{lŔ�L�uդXR�Xh!s� ��k���T����u��  �Cy���R)S����9*����QoM�ڐiu�'j�~f(Ο���yLS�/��ܺg Q�������L\Ҿ��tyDV���-F�S�^Z��9��ku'����[��WoQl
_ƍ٢��(ZI�x�~:�� ܖ͜�Lj��0��������S�)�]]d�vmm<k '��5��_I=L��#��Q�P7Z����Z-0����^8�G��*Q�ę&};3駌7�u'��j� �Jֆ�$�k�8ӽ�c���1;1w$!}�LR����,�ԓWsY��df��.���v"�K��w���4�4o⊽���b�������A���;ޝC�o��"M|F��.�f�dX�e�=T��v5��;��^")��:��&>��p"0-m��7!�$�����B�@���Z�VFa��6D��~*x��~
�a�6�������7���I���<4Ȣ�z�n������ʏ�/���T܋�~���iWG.�?�y#q���1������'���D�\"""X � ��2�q��@�K�$�ݡ�}b�d���F�I�|������IA���w�sK�JYgC.�B�E��j+�i����+NN�@!�$fر�O�����}i��W�aݙ@[���Y��wZB7�Uݑ����Ö7��9ґ�i]p`��yFzA�/����D�|�Ȣ �#:����!�J/������<|��7l��z�V�q��O������ۍ{-$���I�J�����P~vϷk�����_�j��d����a������$��*+�+�v�ڴ�_Ƶ��v�;j�X�%�de�lC��7�58'��+K�V�?�\U���}$�j-����T���o������X}n�uih?�q�d�mR����ѹ���V���`W0<�S�2SJ��������-�+Ĩd�ŗ�&�R�M�����.b�-(Gω�)/~��o8�����@�l�__��NS%�ͽ���0�`��B���/2�ka^��M܏����,3��3x���$u�������0���s�$�*:�{���	/��C?�S��zK�y}$��P= ��_$�bix��a6!��87d��0�V��dB<j1��]*e�n��3@S��֫k�U�`�։�˳���ݢ��`�gH��v� �f��V��7�nABο�w`Stq�H���ۀ��Wl䯲4�{U3�s���m�!�h��H�E-��L�v�eA�1���-�(g�;?-.!盲�MI~<C�B�f�:�9�� '���&��L����Q�P����#������~�P|g���mo�z��(>����������:NϚ��4;Z0��9/$����^�r��:{�_��{���<a͹�K��n}��f���2�H�M8�W������t��wy��B ��}�:ZZZ:�����X!	��\J�a��R��SS�ѿ����8 z_��z%�2�=�6����S�����%�c�̛�_Q�+�̒���?��"t�����n�R�L�2�]�`$Q�Vv�Xg:,ez�f��s#O6�[��VvB[tJs̴%�<�ͼ� nn�2o�o=r���4.����mkW���+�e%J9�F������}šH*����G<Ki�h��$�2��1/�S�,��1l���6�2f�����`�+�H��AIQ�ĊmP������\ùL7t���}M��/rԓbv�Bܛ���������-L.�{ka�4k�V>���zŕ������np�Z(��}i⊸5�3��bFJ�1�\ͥ��5-�>���{S� ���&�!ܼ_��[ xl�����F�4�N2��D�b�K�{c\���{��X���7�f�F��zB���Bmy�6��c�����*@�N�F�����`ڳ ��cGX}�x�I�$��T[�3)&$�3���g��KX(�bm��V՜An,F�&>QTR�D��W;Jͽ���ivݥtsN�#�Ú����î�L�s�r�l�¢䯠|���g���-�ԫ�pL�6�67 f ��L�?"�y���L�o~���s�����:j�.����	���₨f�sp����Z������f�)E�Ԑ����ڄS6K�\ҋ��iA�\Ps�ek�䢖v�w�� H`ҡҝ��he����}/��L�Uc�^Ȅ�� �mpYӮ�R��d֐�a�r�B�}�>4E>6N%2�yH�)���9V�x��׌z��XW��89��6X��K���i�Ə�Yo��=��E�|�I�U@v��C$���&x��H�.�����5
���ڥ
F�
�1���>��y��)Ӈ�务��%M㱤�7�ҋ���[�[
ݫVt�$��D;��I=�%'���1�b5t�����䥫�
�?�[B������� alj�l�ߵp0WZΫ�@�]l��a�5='+E�ѥ��Eq�Ɑ��~kWt�{�98�k��˸�їB`����&膈Zca������S�o���My�}��c\*ev=����0�2'�����lZmb.�H����=�i0 ��[y��d�[1)�d�����Nev�N�[\��8U��NET��1��cS�`XL7-տI|
bO�^��`�_`����q��8+�]9o��Z5�A�=�?�U��	�7�>X�E��׿�&j��*��P�D�p�U}^��O�}y&p��J#z@�� *I)3b���q�����ւ8�*�2��h��3p"�	��،�}OA���N�Mw��
0D�JE
F�|���p/P�|��o�:�4j�֙Z4OP��S�xLU;	��'��::�ֆ�(v-��$�b�Z�o���8��)��3>9��x�����s�:d%�1����<T��� ���L5^*X2��`�1\�=d�oX�T���΀)2<�U"����2/$��g��>c�$�Z3�r4SnT�@��+�r�Y��]�R��(ϣ���\:]%�@��;?2�kEd45�[)�f�&�v��)���X�q3d>ژ�	#�L�{"�s}
]�ϰj]d��ѱ+/�;�]d�S(&��Q�I���;oߟ�R�y�X�?(|�@�[<,�
��ڔ)���)��A��j+g�z���O����8�Q�YpI
����0U!�nR��g�Jd�l@�,ubc�E�af��@f�Z͈7�id;�31~m,�m.zT����
҇�P��M¤�[8Z"��N���P�&R\	���W�i�Cb;��-;�C�"�w�eSW���O�����U��}�sƐ�JMޟ�N�0�v�8
�!E�H�?�m\����L5JN��Psq4�a|\�i$��5
����'�&#Bc'�Qc!W�;F�$^9kAl';��a�Uݎ�ts�	j���������x���mש�֖D6cL1�f97ئf�Yi�g�E`�;܂�@Y�Ii#�'���HkE*a�0�ׂ����љo��ہ�M�D-!��.�89�\!˨U�6����lֵ�X���-`fJ�4�I\�(37��W������S=��/�碅� lK�~�e[A��ek�q��[G =����Z1Q j�s&"]Y�͔�\���R����o!�B`�,��5pd�C�_TI4E�*�5e����q����g@�����Ra
`��A���UcCvy�r:MS�lEuO�Sj���ѩ>�nO'��_VI�9�y#�O���-!}�m�.Ԝ#c�������R3�0�ЬM�&��� c�������M<�LM�9z3��\�C��t��T�.+͹5�ˢMQ��W����l��{��PD��E}M<6j�����r�q�� ��J`XH����s��i)��Ί��nSp}���)C���S�2�;\�: j���?�~�T���H��Pst��^R���^_�s�	wB���r+�aH"�,K4�4CmyF���F�������*�?�I �sf���'rGih���.��to-`34r��	��W������ ����%�ʖ��5�1�-�߬�k~Y�5�Q����j߹���'����Z5bs���r�l�80� ��S����ݶK�G��>DO��t����P�6�`Pi�����E�p4_����ǵ}�-�U�7D� ��Fp�1��Q�/w��)��l�M��TP�z���Z���fe���X��c�l���zQ����$�w���@|�.bb�u%���3�\	JXu��I���/4nf��2��������&����q|�Nƽ�����l�������
^/��"����n1Jп/.e�.�#c�8T���*Il$�G_�H��о�c|���"X3��`�df0-K�c����M)4\m�R1E2��	v��7T��{Fpa�x�~p�ɹ�D"�Lv$�s��FD��LÕ���V�����%U5V�N����q=��t^f��(�x�x�e����V����%(�i �_�-. ��;�X,e���Z�H��Ԛ�>L���O�P�#�����#�%<�Cs�8A��T� Q����bk���R3x�ҵyΫC���9w[3�w��M��J��<D�j���	ޞ��
���mN�P_�.��R�XU��_r�c�i|�������3������®�i)2�a�O`
ղҥ((R�+���"Y��b߶=_����-'����[:w�������.�w�S��U�Z]�ho�܈��$}�Gq�i���n|UG���?v,���#�7���{pSbQ)!��5`&������Am˷)N��
����S���C#�F�M��m�g��޶�ah���!�֑#����ܺ��z ��@{X�3 ���F�ȓ���j�^�#��`+�j隺ٙ>H�e1��Qg�4��.����j=�Mi��v���5��wf`��dJy��n�����.��g�ɯK������*8:Ux<��_5ͧ�^i��^np+�uִ������waQ��uL�c�_��24VW0�`�P�e��u{�`��9�`����LG�)�_��pNK�%��]�+���Y��״?yK�/#qŦ�s�/���̵f'�3��v*�Ϊ�b�"	�?i,%�-���F����@���h�[��6��Ĩ�nᣨ,��Qr���ϧ4Ny�orwtaC-��O��էy����_&�E�M.�	�6�T��U�߅F�Ơy�߾�*w�%Ձ�����t���H$�U�pR�.���e�4��mnƛ�	�j�3Θ)��Ӗ�!�
��$�����N�\��o�u�/��� qVC�v2o�����W��e�����ڕQF�$Cr��4G�})�S��<��O�t�ET�?���|�$�;[D��e�,GH�(X37U���y�V3����DWtI5bJn��������z٤f�
�||H�;�-;�z��q�l؋5�<GБ�U��E+>4��~��J�>LsA�(�?<��<��A�*�B�Y�М�����n,Q+�����~�Y_7��b-X��Ua�U�9?G�&��i�%�	�����5�ビ梙�쥹4�qhk����W���6)�i�ۜ��°��j�[���w�[(�Ì�(T#�����킜l�foT��.�#�B/ ��ƌ�"�����7]��������f��䒹_����"�O2���~'�B�]Ya+�N{�h�e�, �.@Q.ăh��>5����oB�f���H��Z�D��L@��h:/�?mn�C��2}�Y�3k���I���1i�N�9 `���#yV"�k��6�g�:��g'˿�Wh}�t�qo���[�j����\�3w�I/1��"�"t���p(u_:YQ�M��Q��
�g��p�.��+$:@���8��7ݯ��L)��{_�3��c=���-M��Htv4�9��� ݹ���ٚ�4�Wqz��r�W�I�iڋ$�Z�T-A��c���2A�ɑ�~T��$7&��M����܏�I��yB�!�;�8ΧL�wK6m'-ng�vv�Ȇ׬�W����0Q��7Qh�t���AL��r�~��?�{,��~剹��l֪�©2fı\V[m�3r������^#ι�俑qX��t�ݑ�.���ԏ%]\kO�t��9X�u�6�ߟ�^.��6JoyH����%��(��a�����E���]�i���P5"����AF����*�����h���&�c×����+Ɂt��i�FG�4Fli����>�h^��|�H�vɻ�a\�-
lh.؊��TCh��FD��Q�^v����*�qH�� '`�D��>'��~��@p�9y3�|���a�*��i'f��}�6�VK~��^�K8����_t�H��7;����6�ò{¡x�Ni�ܽǼz����v��{�8�8�n