��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7Ɋx�!�g���I{H���f�����&1�+)��ڷ����m�/��(�+u@��K
"��?A���yt�tn��@<n>e�q'J1B$\�xG$Pp��(�n�����k���6��[�ھ���K7>wCHYܨY2�d9����\&���~
��z�0�P�`F�����lȭ����>s�jO�aߐ-��>h�Y�x?�p����m�$��l�|�,��*0�J)��$�PC)͜7Wߦ�K�"��i��j/��
�[���IKT&�B��rN��,��<3�FI��;�
�B��Nj�tO.�һ����s\-����3v�l�����Qc�+Q1r�0eP�Z���O���J��	 �'�={��1 �����9��ל�cod�b#+��Xڂ�ܴ��S����2�l�P�ҍ��:
2~	�*���Gx}�:_!�����t���S�ᤄI5�޺6�E�ȏ��[$%M��� :7a0�#`���J��p"P���8���)o,��$9r��T= �!XtH�-���=��J�q��Z��UX�1�CCo�uI\�:b��e��wK�@��(Q�4d?����<:K�rT��R;r�;��Ml�ȥ��D=���|X[��|Te�'��f\��J�%`�~bh�.�>x���{Q*P���{��D�ϼ���W��_R�������h�]�b�V&�_�)3�V��Bj]X�>_�섈���)Bt΂EC�OOj�ׁ6����S��(Ճf[�����r�h����?T`�^	OӜ��$&jE����!o���ܔ��h0�T�G��o}�vo;{H3wcS��~�J/X6lI� ��1��r��W.۽���V��i�RZo���J/R���[C;�v<��+t� �k���H�S����\T��V�oخMu�Ͽk7�奴�
'��c�-!�4��7DJ2��O����*��fp��7(n2����2���n|j?_�.W�h	g�nn�m����k�_ckW��J)�y�䩿��ʡ�|����ū8�aʉ��xܸ����	8�zm�́2��=���v��MR5��Ȋ�3�g�7��A�W�s#�8í�mh�=���Q��޹���VH�U�skXi�t���q[�\<jȢ��Di�R���[o����+W*�<m-��4t�ԜQ��w!�bXT��r�t]��c���#?��ӟ������g�{�潈=��"��d[��G:Z��důyT���jZ��Ԍ��8�0`Hi&9��El3Zg�&����pU�X��>�b���&��j-��+�'w����m��	�?j �.W�L3�v�֒�~%<\L؝��j,�0�����FA�Dh\��k�2�g��B��|�e���d�̾�Ĭ�}19�oHdf����Y���El~�y�Դe =-�o#f�j'Ud�`�n�C����4X�����x��i5۲@b��ZmG-T=Z)
ܳY<�%	��0�6Y�0Cv�Tg��)�}����u��̯uҷ�a� e�0p��u�h��g���%�pM�+߬��{+K�+2[��rs	V��]��6�U�ӵ�f�ڛ�_��z�p�Ѝ��}�|�hV�c=��Z��,�&��n" �b�$���]ǝ�v(oQ.����#!�X��W�h�̾�Uf�B�O�ܥ�����6�����~Zy�#.�ŚP2���«���O���������5𼀓6�XM���Ǐ6�J�e��DXx���w�^�Lf�<�����y���@K�z�{b�*|��K�/2{�]�sAB&�(�>:[(�b]�0*�Xut�0t��a��a"��S+�h%O ���u���I�[�\�`���S�˴:�.悟s��*'�`��.�78�`�r�F�a���G�� ��4��u��D�W��-�Y�?X���26Y^hoD��F����c�h�Q�h��������VU~���բ�����˔AWMk[��I�9�os����9��D(j��� �%�9-;d�m��y5��:Jj�}H��쩕����
�&~�j�� �¡��ҩ��L� ���9�/���;Yv�� �C�e�,�+�e����竦�	����@	�IDaT���M�f,��#�V��zzKVo�ܒ�zk��P��L�N�����
�����0�պ���&�γ'ȫѸ�;H�C(�_�c���v>9v��pfq�1��:���_Nm�<��4?�"n��wά���ba�|��[�I^c���x^����@FB*���:�«�}�f��:�P:0)U�����Q�i��ʡŭ4d׊	7���ϳ80:�]n+,d��D�����3�l�G6a<�V���xZ[�R��q҅~�}"�C��5����U��Y,^|����t��2y�e������@�X��bA�F��+3E��u%�9_}*���M�4�����V�=x���K�6b��|�������ya�R��+BV�a_���e0J���E%���Tf�gr|��k%��sP[��e��� �&D�p�9�/�|��xrY����I�͹��žA�����c{=�S��s�]_"�(g�v�'$W�N.�;0�z�`�\ ��e��
��j���e�υr�8�Ĺw��"����nZ9ރ������*�ܓp�챙�{�sP��6�n���Z��d�<E�bz��hE^v/z�ݾ�(��t��ST��2���.���KlC�V�9�sI�{�_��a�t�:4h�vد�h��*N�u�DmqLMZ�Jg�G����[��p�!��$����DgE�7���אָ�.�4�~��cC��>�;[z���3j_33��r2���(%Q��^��B��Ƃ�HK�κ���.���}1m��#��w�	g䛹`;+��b6![�C�;(�������י  �gB�(�Ưn6Ő�h\�����o���_j:xC)��TC	�kLO�w��q�_i�L�7n˨���ƜP%
Kz�n��_[f�qe�%��d�
Msde �*L7f�N�T��5F[�!����t�a|+(�@I��N�Þwޤ���6��Ő:�_C�7�ec0X��.���x�T� �[�P���g�|{��;���<����Q]z��)2����W#�8Xt
��uy4*5@�l^
�7Gʣ�Q��B�M�8V��A�e�C�gb�}˔ߤ���}�9�YX�)%�V����v��h�^ TX5��0#��)�ˎ,&���/��M��"�����l��t�	�*��ݻ
o��X�0�@�T0a�N4ٺʉ��Hz���O���~ǁ?w1�U좩8K�!+��`ٓ8���mV��J��餯2��>����̎�=" [rn,Y}8���~�s�=(,�Y���tЉC!w@����v�28�s���:�� K� �}��R�m/�N$?%���J�1�]M.��3UV�����pd���n��]B|��`q��xj$��_[�;�.9G���:��e�L�v�^K4ܩ�+��N�Y��+���!�Qp&�{�QI�Ԁ$�H���\��%�s�!��زF�|�g��0I�Ò�GXꀞa�;,�T�}l�=�$ï�[gG���~���K�}���v��訑{p��r�m2}N,��]�w ��~���X �"Г`Uʫ�#��l����WRR���Y��N}r�wnȍw���!e��`}d�,� ��.��������ܓ�,ؤ�e�D�����-<-���y>�������g����P��i?����
H������&���g/���3FBG^�E���6NF�I�s�-r���=��������fus�&�@��B�~��Ht�\?��"�)̲.g�"^��P�Up\�~18�s'\��	�R2-��D|��Ŕwd�� ! ~w��3�2�-7ač�L*4��|�߰S��^���uþO��#�N(\:ÊDC̫�T�XID����㢕��?6�S4���ͫ����G�٣0��2� :�,�SX]A�j1N�T?�ֳ��v>����߈�
�F��I�C��>����j�u��0�m{\�x�=aq!Y��a4���y쇼��=��#�l�����S8��>����2�<\�Co��b���v���;�YD ���)k��,��
qMΓ���"��M���x��U�f�y��-Z�8/M��{T���� � 5��U!̈́V_�,�xj����kE����o���bO�60^���r�����
	�`�Z�T5@�.Ӊ��o�+̟"!���.qiE�a@ ��%�qK�_Ƚ�a<���;[��9^��XswOi�ЂO�hɼ8"~���F�b�ed%���*�P��Yx;Q�Ϝ~Q�/����s>O�'5�{$���������RC���L��
H�t��kI8�`� ���\3�v���r����P��фA�����*�pXv_�?��&��G���/�n�հ]E��^3ĔK:��{H)��/�٦�e�����m�����kڄ��Aȷ�S�n�Z�#���9ӾO�Ǡ��tH��X4ƾU�д�H8ɐ��b�Ƞc�E��S�N�b���.9I!���V"���p�Q_�f�e\g�����?�8����$��t.\@��Ў���n�ˊ�趄���;��K+�<uj�ꐦ�[�TG���!�����'�F"B�ͯW����_x1��[OVf!��l�Nfq��>�#����P���s���\V��1WF���/$9׌����Hݳ�tw:�vk����]����O� k�T�㞇�\�N�5�:��p��>�Ɠ/�D%?n�j@�q�Q?��Ƴ�����νME������B�9:����>U��{�L�5��ӾNw��6�ތ��=��v}�;٧L���6&mOu��]T0�=��D
xh�>�4�d!}���j�ʼPv@�R-]%�+�Ƙ��vf|��1��-��e_r�-�?b���|4S���a���Zu�ߠ:w=0����nٱ;��^�6z"�/�J�S�~ة9�M�c�=�M���/���ʃn��/��=��ã��l�$���(�*hט��N�n��<U���}�.����W�1��z��?y��.n�"2kJ��N��^��ɀ9d�H���N��<�Ļͮ����?516t?��>S�}-/�R詃([���,:V,#x�0R:���*�gJ�b�J��NW���h�Ɏkw�r��ѻ�>v\�ɃJC�e�\�V�G��-jE��Xo��������OQhR!���7�S[��EWsŭ7��c�A�px��0�P��8������4��^Rh_�O:�V�H*:T7���/���"��%��Q��*Zh�T��+Ċ�63�G����6�y1�<�gN�n}��;I���m��}W���~��ޣ�M _�oj��3�gTѤ�  ѣFx����!� ������5������?󼵮�q�z�kbr���r����h 2m/������4�;^���uGؽ�j�u#��j��f��s�D��s�/eN�haňQ�\a�PG��.�p��qKa���t��vo^0{*�V��q�zo�z��qqMLv�N�ʩhN2b_n��i�Ⅼ�p\�/�iTY��O�2>���g�V,�/u���0�G�j�fƻ���k�h1�E�� �qHSܺ#�ҵ��T������1wG)�xKLu��(���'ŀ��=�i���b[%���R���{���`Q>,��d�r�1R��퐎þ��	U�O}�m�*QSH�۾p�=�I�al��:,|��q��_���I�q�s�����mh`��($�j����-c����-oH����f�<�N2[���hd]��Ґmji2Ȍ�{��7ak�/X��賤bn��y-3LՓu�@$��<̌c����KW7�ʼ�1ĊbUz���Q�Qs���Z�3}��> o�W|��C�B+�H��dT�=�L�9p�_�q������nz,��FL-�/�O`��5�rOS<��g)�l�Bi*~�����^���O�c1�f��?�����K[�	t������4���[(a� �.�Q);g	�R���IF�K��h�1����>V�͓)=�� �GF}+��&�U�f��M0&���k/�yI�.�K@x�5��Øjf;ٕ�>���C�+�C~ҋ���suF&�O,���  �q@ F���#J��)<��Բ۬#��ROJ��A�|�t���^i��F��ìT�vd>!;\��ʏ�/ۭ�z��T�S�ƒrHI����b�>Ӛ�!��Â`�������o�Re[��N���1>r汽ξy��`�Oً7t�^�;�����W-�����q��YAߙ�����I�]�CO����_;$*����.3���$�;��`ukӘo��o3�R��X���ڬ �i�[ń��w��Sd�q��-.��B}j= 	�5�O8��8
Z3��>#X7)�Ô-Kr�N�Ԉȉ�.?D_�AqO���j�8���^���;����M
�E4%͊L,�)p�L
)-�Llqy�RZ/�s'xuP��V�'�.���E����@������uyo�NIߢ�ޚD�Fu�F��Z`��@	!�Q��Ȣ�8_.������ۗ���z��9�={�i>�f�\�<��<C0�}��}�<I���lc��15�ȅ�