��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb$�������N����^ﲇj�m/+n��O}�wO����j$�nz���Ցۺ\S(ӡ��_�[�w2e2�s�B��@���+E���L��t6x�9���Hk�D��?��n4��ۄ��d6Jk���X��`���l?��u�sa���X2ꬑYq�ـ�}�k��	���o����X�y�4���ӕѷ��"�o�jlC����ǀ�
ݣpk/?�ȱ�����	(�	��e&�7!E�p��-/��p��+�=QG�k�(���i�T#�#��z�Ԝ\qQ0�=���la����v����;���i�(١�/���pNm�6��ߤ�w�h���|�D�n�`|�u�����='p{�)5���� ��M/�������i�;��p[Y�vmm�m���ы� �K��&���P�-8[`���v��/Jvt�4`�,�-�w��|��X3�]g[gc�@_c�J����ud��
�SáT����ze�՚�Aa-�8ֿ�C��^�Tf�G'��Z]�
�?��趶��d�g|'WV��l2%*���I	u�k���iQ�<;�_��T��9r���̐;\�
�qi��Vae\4~���fs��X�U�u��@�#�y�b�\6��H�^p�PSU��0�j��nI!iq����0L����Ng<�|q6�SI>5��,\�4�V��>a�T�tQ~ аq�������A4�k5crA�r~w
����W^fQIy���	�`[,R�W]�te�(y�=���[���q�|0�_��{���0Xvl�!�'�`;,���g)����ٽȇ���Ѣ삚�Dv�����o�pM��Q�\���5��q��y~�Ѓ#�ڑ��i��&0���7B����'�NJFf���kR�P�+;G
��^E�[Ed��� G������n�=�D_���Z7�+�Y�(���wRFX�Œ}����T��:�=��14CǍ->�*/�u	yx3Q���>8w����NlE�$��sG����5�=Z�
����r���Y�1�MH`Uߔ��̆㼧�Zb�9������[�$��G����+� A$mP�m����ѕ����/3�  {������h� 8�ԞsD��j�m�Oن7���X�Ͻ��@ �d���[�f�0��i��i�Ci_��V�L"-����Ê�I�D0�2Ѹ4ە�}gDX�H��-� �J��^<�Ǯ��f�U��-�8Z�����h ���9�G�'8����� �6�{V�/(�Vp=�@|@���G,������zOI�S�/|�U���/�wn����
������aoK����g�m�#��s�����<�9�ӛ���|�c�u?�F��z�]��F�OO�����:�?+��hi�,�"���P>�or��Lq[�<��u���LdI�D�7'WT���k�x�wQ�}�����ޒp�9%~	'ߝ�\�*X��'��d&Ǚ$Lo�,]Bs��䲘W�6�8�	�x���m�4ERP?����g/�|W���p� 5c�B3R��iw	�K/F���?�|����G����� #� >9<�my����}����-U`�`n�^�Mêb��:�=�r�-�C��_V��P��5H$т*�'Dّ�+�1J�Vsͮ^���)�평�mw|�I!~�6�s���Ϙ݃���@B.A�J�2A֞�!�]@/Y	�2���ud�?Xu�h�pe�CR��� �xL�xc]l��8kO�S%Z���M� +�w �HW�r��OI8(=���=�K�[Ə[�)��o1�fB^F履� �:��vq�\=M{E�)�h��l>c<N~��hי�D�˗H�L�����֯Ɉu-��M�Su=n�&�%�Ԋn�[KS��ΆT/�!8 B E8�t�[
��u�;��+.���m1g��x �/�B�rP�X�Y��8Y��'ܑp� �Q3L?��۳�m�a׀�[U�P(Vc�iU�$8�x����_P�lS�z-~�`tY�[�i�֝��&hȝ#N��e��i 4i!)E����<C�qr�Ȱ����p�Sci͒������p�ף���_ tѥ��e6����:��H��][��@�/���{UDo�b]ܼ��%�[b�U\���@�KB;�)��	j��E|�D(R�L�N@ �@T��p��~��lc�iY���_}��r�z�'a$d��-�-	C�������kca��f+�[��$ͻAy��#��`�)�7��l}���1dLl����H}�'����sGR�Sb��5rC�!_%�vƼ��O	f9j1���9d,��x��z���1A��,�Bӕ�Q@7������{T��l�c�w>@\bH�;rVI������&rҔ���*�����#J﨤�w�����C	�W��U�/�C��ԏ�$/�q|sr+e�+�/ۯN?7H��*���h��j��<L8���S���o�n�6��O�Ysk<1A�z��Ц@�p��XDM���m��k2��n�� ���i@�5S^���"�PSDj�Oo�kI���H�����)�i�S���Tf&��9�x z�/��l�^x�`L��!f{��|���)�&ɂ��M�:�|2�#}�(�����t�)!�+9����ؕR�i�JK�C��a"X���(�I2U-]��ڍh���������l&�Nk��sS�ֈ�"��6 ��@�Ol+�
뫊���@e��aӏ�F����?5�� b�u�Dv�b�?YvL:����@��\i����7]P��#+�p���|:�K@���p�!��cW��f��Pe�x���Z��@rO�V�ߪ�Q��y�p�Ȼ�Մ�6����y8���0Z����wK(6��)��;������8>���=!V'
^mss;�tj����^9�+��b�X2��Bj�*��7�-G�x?�M�����0��[���8�h<�g��o"��b��c1+|W�3g���%���)�j�9^�z�XPs���j���.� ��b�g-���JL���F��
��޷��vSi7s�^FRӇ>����2�;����v���o�'��^��靛o�|�ـ�\�W6xcĥn̞����M��7)�5����L�O��C�x�����tV�:��h\u ���YS�����F�+2��H"�gP=]�gΰ�(B�?��&��}���O���n��}O��yn�e��+ɰ{I&9�;��E���x�xo@P���B�J8�oʢB|;|���+��# ��e������V���9s��+)���.�2���V����
�F��"��	
��I	��u������S��4b̨��e���x_�!�35��*@�/�?ӮM�+���Z1�x���D��q����I�����Si"m�QG�L$&K�Ñ�~�ao��R�{Pd��Z؂y �fk�6���2�2T��m��5���^�����U��O���������%旲�b�K���[�Ӯ��%�y��ų�!�(^�\*%��9�M����w�s(>aj�GJ��D��]
�PH��cӣ�Zb�3>(p��S�i&dʘ�~3� `E2�%1
"�~�7$C�)�B99��&pm*~<�J{�'���m��|�U��&���L�r=�Dn-���\zM-�
'5��pV�;8o:%�j���J�*Uzwr����2FN�ou�♇��){���F�N>��ga��v��J3�KK�G^�?+�V	��͊kEk�t+-�2��~�,�J?�{��L�Z�xi�Y��s-�Uꃕ�������k��M�o�N�ВU@0/�8�:�G��%�����a������69�ǶI�-Q���ʕ0a�ڑ"��X��:�E�"[+f�
mp�bF|ܙ�(�J>k5������Zթ�JV���7WP� [d�5��Y�u5O�1 ��4���dL�ס��3���f���I��n�i����"So�I��yB�ԕB�#�*`��z��T����]N� � ��0U�4e��:&LO̘��#4u(���g�hܥ��`�o`�;����9�T��W<����9 D��_�����㍐�6��3���M=���J>W���
��F}R��w�q}N�L�|W�%hq�!v�����C�q���b�y�햏!5�R�L���*,��G`��$�`xkX�_@���)���w-0;�hv_��.>��;Q��$��$�,fc��^�# u��6�a�j�'^ #HR�n�چ�>6ݫ�D�@o�p��-��1U/z�Z��`r���"�p��Q*,�^��ى���!	���MV�M�HcSH��&���� �������j��'){l�����6M�}�/�_�p����HZx��
��y�1,�d!#�:��KO/ض�9	'�>�#�/!����gO.��)**~1�L*r����NPb��:َ֞���_ᙺ���l�/@Z�A�3�N�;�����j>Q+��J���\��L����L�B�rcW�s �l�H�����|�p���m'&�{�D奣-ӗ�sz|�J�3�;z�F@J4�i���*����b��8�D�aٛ��F�!��A� �����Y�ܶkkB�����f�9t^C9�����mO[�R�9����Zq�#��U~�e����nXZ��	��7	^X�h�As�y1QިI�)J�����#.ҩ�)�d��8ǅ����K.k���.B3�V��{�3��uc@3��� ^����>�Q
�����hVP�>�P�@! =<���6��0�wha�����rSH@�:I(�m��U?�|�����KU�	u0����7.o�B���E.��7�m�\�G�Z�RSJ�fB�>�s�
�t�H)�r�L�#�֠� ]����A�V����Am���wʳ�ʯ''��+t0e�W����Wh��rs��'l�Y�e0>�1\D/��f��l�w-�,Z�T�[�h�9��H��U�l/_�Z�e�߷2���TWH�i����B����+���<����1����7�C���G�[U�C���Di,�CL������eZ���y$AM�m���e��D��vn�V�:Y<A+d�|��e���g�e;	#�.�Xgvd�`B���1�c&�F�X���镦�2)Ҧ�/�JR��� ��m�$+�lFpQ۝�dn3�r|�5��Y=��B�H
ntH'E�A�O.���
q!d�*A�>�a�(�od+`��7��S�w��m&`Y9��V��9��H��̹d��۷=�@����7�,y:A8�ͨH=M�(�W��oz��D�D"jM��H7G�.�w��|�i~\��h���>�6���1 �"�c[� ���Bv�}?�M�	2���v�z���2�H����0`gL�Ӡ�?���XڧY80
��#i=�m{-#S�����^#*J���A_�G�Sw@|��XG�N=3uz�Z���ǘ¯Ǥ��x�	i�M�8R��}H��c.t�}�Ls��dL�3=�Ć���2G6K����S�S:��)��P蜟��^
=�hni|ͳ�T1�Ӻf��(��{����;��ϒ��Y\)Q>+�gX�n��A�D��Q�T�d�X�`*��;��� ��u�ӽ-ۈׇT6�m©	�3�f��=�@��aX ���kQ�#+�$��[4��
��s5�~�y���*�A�K=.�.؏f�ITxhX7�?�+��u.퍞Y*��kQ�1�q��
�z�c�P�1;XF?]Ο�r�������G@WQu�z�-��L�A��غO`��e)lC�`�̝p���s��a�u�>��}�`�,#���Cq	.��=X�s�gH�v�h$��z���W*���u':ៃ9-$&��U�ih�m���Dv�B�v��'G��H
�.	�<T�ƯS_��XZ�K׏��wk̷��A09:ۓ�Im��X �� f�\�(
@إ���~�����ќ��r�rC��&���a��q��X����� �>bI�O�Yp 7HL�e%]GA?U�&���}�C36
���Mp�0�\�g ^��ܶ!(S�%Q�J�)(q�W(�f�BiiU�/x�zㆎl&�����L�:g>�r��E,�B�x���0�������H7��v���o`��7��qBCcc�`Mq��%_��/�˛ø�i���GR]Բ�N��r��*��J�Ke$p��k|g]y���냻Q��Pg/'���4MDA�ַ����j���(�J*^6��?�i���x�;��������m�G��?�:e6うh�[!��2�lP�Z�F�@�n�����E�1������֥��a��RԠ�gq"-f�E����ݹ?����u˖�!'����;���(����:��Ų.� �-H~t�Ȳ������2���=����3rj
���'�|_�BV{���Y�W�
��W�1c�j0I�3�u��&�k�����3�����Z���0��g)Ҡ %������Ԕ�.~4K���gK�Э�.O	)�B@w�%f넆�����k��=ʴ$��| ���̗����������;���j�߭1�p��f���R7Fr�FƊ-��A���@%�����D뻱�P�ڇz�����q��U�{��GD���vm �V�:0�	ߢut)8h���!G�*��'��trRf'��C����am#L�?�eZ�v���Q|RW����r,�ȋ����Dg�Jn=�Z�l ?�,6��[³WjVd��Ц�+���ʹMw~LH�V[��ca	���~mmF��u�3�UA:�#��~AG�i�e�_�K�����v*Tc�Z�Y����G�W&��J�/�5�v�3p/k����M���n�Ie0����"�g�+������7r27��V�^S?�mY�f>��:.���r��^�x�dм�����.?D����m%���p+�i� ������Te>E�K<.����-��r���Ѡ�^��,��Ά��(���D3������C4��3f`R�Y�����9I�+���) p��s!�(�wy�n��F Bym��la�����B`����}�Ҍq�D� �n��r�%�Vt��jX.Z�O
��;�)��N�O�[x�%?ˢQi۾��*��u��2���;���I}{�R���Ʋ5 �"q8{��剈Q��9��o����g���j�!0ľꕕ|CQ�z�9ݛ��1(� �nB�y�J�;�#�26>�L���-�F����|fQA��q�&E���?�Gb��.��]�@Uݾ�>?�U! �ˎB�����Sgmm��4o�#���^�l��p�A��w�,��7�c��I� �VƸ7яie���[.�!����[Le
R���B�8�°�:6���$�	����V����r��ص���)�;Qʧ�S��D�G�Y�0������U�A�k��(���p# ���{X�ԐeG5uH��3�ɔ��#K����Nmqc� �'�C�_)�Z��e�Na���!=��exܯkE7�b)��jM1!'+�������s��x|�y���n��v�mD&v�����:L���e�bm�V�jqp���t�+��	SB����/[!�(ī��L6�l}M+�6���ݡ�������p��b�^EE��,g�V���=�>uQ�m2{�9�Th����o*W���rv`<	Z 2;��P�K^�,��w��9��1|�#�.���9/�฾��ϙ�
]������Ɔm��l�R�N�}.��?=P[p�
R
{���zq��	�3���|�tT�sVݣ����Sx������0ڼB�]�m|d��v����=h�S�2�G�1g��X�m��&���h˜��a'3�yO�dE�������!�{$���k&�<�l�h����ѹ[���k�V	$���;X��bO����2�]!*�o�t.`�'����e����g�F��A/dO��g�0>[���q�pΎ��K����]��J�]�Ȍm��Ж�o��4�(@n��(P�)����L}���=��Ȍ�^�Ocj��}������|HQ���&0B�瞪�R�}�B�跇a���+�-L��������Q��G�r�W�(i����ɾ)a��+fv���Jm˒�k�"����!M������Z���I�� ��h��@�9g�iz	��%����N>�,����P<M�һ�G���#D�ѯ��vL�2�d
�Yl!Eso�"�G���(��A
~Y�<���<U�Y�C�!��p���#��^��o�Ll.'.>�c�.�#߁��fѧ�,U��Zl�JШ�CX�<��G�*����(��d�o<��%�'l�z���>aEd��$^*�����֐K��'��!,⋩o\$�:�!������ҵ�9C�ʬB^�a�ps������2��sb6#��Z6�;�����`�Ź�c�H �=�H����B5���m�z0cȔȜ�-�E��b�>i�uH��Ki�y�>�벀+>.��T�˝Oe��S*��:N��Lt�%U*1 �?n��=�M��B!s��:����#:�����"���a�p�����A�0کE�PK�߆�{�ѣ�W���1�r�be@���w�f�+�6/�n ���
%��H�yɠ�v�=���4��f�<��+����yR�>Ḵ�J4���M(�5Y�1�b��	�k}��B{�
8,1�� ��`�H�C^P�3k͓���òH�F�˄��o�;�=H�K��Ș�ގ�g�^s����� ��,[\��xI�~��=Z���e��`i��Q��^�Z}�-�uu'�t_�jfgUV��z��e:��6(�/�%��I�6��Δ����	���ZVH�2�-���r0k��[���\n�ˡxѤ��=/yZ_8;V�I��k�ݪ3�P'���g�*�;��>}�Tq���L�x ׬f��d��`2
�~)�yc�C5}���%�#�c\�������g���h.���VR�LU������"���t��t�
j=��隊q2,����}���<E�D�3bոN�?�m�۰D���Ӗ�����:���CU^Y�S��5U��^�!9i���^&��E�`w}��o��!��5��:O�E�%��K��&)u? ��{ �!��$��Z#W��qI����e0;�]թ"˺ɠ��W�V�����D1��F�1�ۦ'|��G�$��TI��'`'��e8m�F���_'�w�V:�Tn�+>L�\v|
5v�!��F����_bpZC��䳧��*=c��3.u<���c�q(����u�����i�Y��a]����$�4b]'L^�,<�c�Y�Blֈ�7R�sH��<���C��T���3�:Nh=�G��j�D��J��G����?t�����.����{b��V��v5"q@U��0��/)j�܊�*�E���,pt8b�
˘���3� �򳆸��6����?� fI��I�l��(�G߸�	~^Gxk�@�{�@��\���X���W�N8{xK9�@����|��(W��-��M�dxk�鳀�b1�v�X�v�ǖ�FxZ�p��q# Nq�^	���}��,5��CJkt���9�����dA@��H��J,	E�Z2����g� x�/f!�i�<��#kԾ��+פoe��g�Ch���	�4"�iN/��vy��H{�^WLH� l�1(�|.�_��4���۰�g}��B�n��k�+�pi��ͷ8tL6��