��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbI��2��Ձ_N�RL��������lx�^6�:nn��~���KJ�#���^S�ߢ���#�����a��=��#�5���ʉK��~��y�n�����\���iB\f���8 �!�)��T1Gjp-V�i���Xg�ڊ�-���]�=I��7�ٸ0�>FK��-G�.�*=�!�Ձƣ`�H�C;G�~�k*�N�@3:Lijݪ��2i��O��J�1�u�O��U�(�M*�S߹2���z�gw�o:�+fb�u�{�1����5;�0�0|�
'���[&c��t�]kg�;����&�}�R|��nß]�:`�]b)*�kE�9�������D�e�k@8��Q�Rß��PUj���Y,�K�>`=�ep^P�����s��o_L0�l��鐃�嗛�û�[fj���A�m�k=b�Ύ���o��Ν�e�/dE����F�vy&d��hj h����Z�w��Di�dך:��`�?K�)��v���3�Sj���_UI^�<t�W��ʛ��*�@y������2�@'T�0�%b���E����gFlo��^��n�����k�ooJ�Y�F��W�����J��Ů{קZ�-^��c��!~�},_g(h����y�Y�S�#i�n�!��ߑRn�H���`�>:�˅Z�������5�T�]������~98�vmu�:�J(�_w;\�#����>��M=	,� ���i�b��c�0c�#���⇻�f�]d��j�_�0�E�G�s�u���s�@ZE���>��h$�2�v����Q�E�A�3t��s�D<U�Ĭ�b
~-�o��Q�J>O��f}�tb�1k�y�cr��\`�,�n��W�����0T4�rk���(�T+p5y���Ͳ��M������!Ԓ�B�D�1��ZjqqM�5�D���0F�]:����1uە3���y���t':*�����B��g��CF�{����QOx�*��ʰmg5�Ǯ���~���}����1��#�9C5��fݒlac��)Cȹ!,�u�K�QIl'���,g���twN��#���muñ���b&���K9F>}t�wG�!H �l�⮊"��ͫ���'!�c��QB���*+��\�TU����:�<��M5��w:�Dab��k6G�c�S��A�u�A2<�C�?N�f)�O4CKQ_�j��A?�u�S�F��U�Yc;m�n]��?w�	}��h����z��k��&���(Z�g� 4@�c(*�#��1&o�Q�	:9�My���Wv��s9���"�F|�C?(v9}ռ�'�Ԋ�L<xӓ![�K2�6��9�3uI��q���<��G�����M$g@��1�\���}�2#l��>;����7���GW�$Kz7�vl>�;��*`�%H�ed�M�B��F�`���e�{GO�Ⱥ_������@r�����[�k��څ4ݽ���.{p���Gh��~a�<�{3�y[�BJb�/X�禵����/[�"��%��K�g�ב�_��#��A��u/�G�z��9B���e�f��:C���^�A	Dq��4�'��s��X�BO�I�nI�i�R]�8Aô@I�[cg�gi�O{	��b�)T���H���tJ���i�
��Y�:̂jՔ�����ZSy��Wu�p�&ѭ��p�4������Ц(l��I!WB\����&L����%�/�Sb�K^:�=����&��ҍC�@���C2_��}	����y?��o�p� �M��R��20U�ܳ�|��:U��<Sk�T�Zy=�;u��N����z���@�<���me�߲g�t1ժBOM��/�昤
�Mc��cqA�\��7P�7؋��3��PQ�Ib�?Z�g�
�7�5�5�2�����{6f���ZF��M�����؍n��4����ջZ�4�
�y������/5̱U>H0�Σ0c4<X��a�Զ�"����9+O��4pM^����1�J�f��E�]m�el�QmVw&+F`�'X|KV���fق����.|`. �Cow@ZYU��cb�@9�@��akoo�͘��^0Cx&�A����>w~��������ۍS	BP�*�5Y��<��{�oq]��,~���Q��(�7E�ߘ��圐���G�:�,�V�~ԽW����z�b���m��	�Fk^��(w{qUG@�1ē ����^�0su�u��=" 6��8�L�$�ǧ��5'�,]����;q?�OUY�lq�)�e$֧�|���`���B�� ��[���[��m�ߗ����,��U$r��GqHfQ.�@��b��ړx�a{|�_J�UK��ǚݰ�<n]��-���5�F#�%�A�aԍ3mMtk̹��2gk`�C�� ]��q?&�!�_vr�C�Ҷ��u����A�^�vWK;�!�;l?�@\K�1�A/t� ��C$��;�o}\�L����a6܃����ح��1;.��Ĳw\3r���<\�5�!��L2�&o�-���t��ÿHd�P�ȴ/#���q��E��
���Lv�3�����D�G߲T�3�N���M׎���)7�&��n3�	S��T��A�!(`���5�K�>�V����D/k�fw�'yvM��q�P�������\�4�&�o~}�8�b��JL;l�2���M~ �PGʤ$>�t6�M7�+]��#��	2n7:�E�:��BȲQ�[��^��&t\���/���-ޫ�"as���J�ȂM��=��z��(�|н'��^4�Kᠿd�́}�F��d����#�)s߾�X��	?Q�i��>R&Ӛ�Yo㢃*��r�S�,��©�k4X��q�E$��榌T0h4)�yH�^�iC}X4�D�ѳq���i�"��z�lqU���kzYK��yD��ˍ�=��ӿ���
vzZS��J�ժeA"#L�Ӄ
wҵ�N�5�=~�_���1�'�(�lk��F)D�-�nW*���a�vi���(�)�9ޣg��I�C�iKԯ���[NN}WC]����&��x�Wk�w~��}%A���3�^E�ե=,ņ^�1d\o3_bxk��-��JXlud���([&?�d$2��^���lJ��u�C|�m�t��RA�F��A(�� �҄q�$ṵ�����L#����с�Tubr����6gq�v%��7���kg��KPQ�JX�{��u���j�m)���gȡp�m��;��c��	e��(��y^݌�z#=���W;�(]d^���[���#�_`D�܊4	�����^iP�*v$�dN|�.���@�VT��n��~,)��������"��`-&������NV��:�y�PZ�Ŏ��U����Q��/�y#"���
j�*��p����4�}�yd$|升sߧ�z��A���C#��'�w	�
jl6rd�6��X� X6Hw���

�o��^�`�4X�6,~k*^$s\O�˥I�@���bb�)Ɠ����N&����P	�"7�ג:�e�8�A���%zq�g���=�F����Z�2ߋ7�U�ř��PJW�b�\���|_=���Ț��ŶAW��_���l��~��8����txҸ�BV���T���o��\	�&$aY�?�eԼ�q����/1f�m�b�$]xc��>�PC���T�Q>�Z�Y�_� ��9V�}yn��.��K@Zn��8S1��
׬��R����>�5��z�䤂�:��-�"*��E� KD�$X.����B� �6�}����[:���w���s��+��t/\X���B�e>���bǂ��f>n�C������ �H��Bp��Y�"�h����w�s~0��ջJ�Øп���/�MM �(�G�+�P�5kڹI�Dwxu�u�4��gA$դg�[�y�!�R��P�٭+�����Ñ\��H�O89e�����3?�����,�n��e��)KB2
l	2�">��/8J�v�9�"��aRv4�2�2R�.��u�)��0B��,Y5�@C2a{�,=[���q�Uì ���џ4l��xS�0ACZ�?�R��� �%��^�ɧ�����3����o�C�N�b�KD}l��Ԙ(d�= ��*Fǀ������L �TR�obޕ��Vj�C�~wYU�#��x8�|��K4y��d['/AP'"�m8���3��Az"[�ZXzD�JrV�����Məb�W#t�����k�u����K�)$�p�GN	���6�^��	�O��e�F�.���������/Z�X�?E�7����,5�BҌ-M�B��՘a�O��)">����!��S�NDB�E�S
��3��{uۓ͜��qt$iA�2�X�d��_[�\9±G�s�6M���&w���K8�F ��MD��R�&u�L~|�'(�OY7����S��h0��4�����
z�3WI$/��}sgO��l)Xa�"$|���pOc��0���ۘ�>!�Y�z�����~�����Z��D��Q�S�ズ���Wb�1�(�g�P�08�q�q����KV�s�����$E�[�`}�{v��nI�TM���}�bd'�<Ǧ11Z��h��P��j�>���TZ�q���Y݁% ٢X���:8�H��T��yQ�>��������xo+��e�1�PR�RطFG{����y��2�W�9K��2��6�ӗj+o��>Ǆ�R\(x�>�+��"��P����у�S��t��`�_	tP�E�����]�����d��yV����bt�!�/��ǉ�+tHj`y��K�1��{[�j�ѕ;�&�̚��Tg"������z#�k	�4��:�.�t<�b;B���'`쏼�x�H�H7Ѻl��>�G~���SF͂(b@��P��V��z*؃icO���j[������Y�^3[3 �	���?2��"�JГ�ʪ��{�ړ3�d���B�7 7�?B|`t2����~��]0�
�D�%oQh��O�^`y�%�Ϳ�\�7�2#6e'�	+����}��mN�}���{�������qAUu�7�����#8��X��v� �,����4hДs�@"k�O��_�����>'� ���Z:��á�_���3((�h��wξbɲ�N�H��a��!sђ�؇z5�	@��~�����k�k���͠�E� ��]N3�p� �J��>��X��ڌ����K��敥�D.��$8��x�����o�J�J�f3}S��+t^k��ݝM�|7��F�!{�?�
h�k�L0��y�3u�G�؛ާl�x�L"^�����y4#�L�ΔM��,�c�c�W���\3=�n޾�?,RbN9��)��fj���b��J�����MQº�%����P���w�l?Ӗ7�q/��1��#���W�~��o �b�	��;�L��M;���˛��Ty��om{%���6|�O��,3�a�N׆T�F[k��w��P3��w��Tn_�םn����"�t �z�����*f's�G�G)��$T�5<�a"E�ӕ��u��t����5��rzs@7O��S���d���a~q�D��S�+�&�����\5^�������]]����7o�,��훢��F�P��m8�%����'��|��
��?��D��K3�/w�2�QE!�����U]~�5��>:���)$c�'�2�*o��x�j-h/�o���"��禃}n�� ���n��l��m��цMW��#֓�pU�u�i�����4�;1����ӑ��?l�҃��lkqo��{W��P�����2���aW�����|ၚ�|�V�����t��U"}�����v�Qޘu���ðF��	�)�M�L�o�H��-�h>+�0�σ���~H��#��JR �&��$�#��xt���"�N?`�K&xW�O6��Y�2�Ԥѝ*��̮��D��8��Up�4_����m����R�Gf�l{�u��}93ƿ �tR*���d:�����4��@&�U$��nf&K��e~�qG��i��`?	�L�f�$�葩�-9W��� 
��庱FT��&�0Z�:�{u�����XΪE�4���ܭ-�@K�G<�`9H	q���HA'z6?��;��;^C�c��E�|)��G�E��u��O;��졩���*3��4#�k%m8`��C<r��
�-�Jќ�C����rܩOh�74�.#$c�Ș��Q|�}m��n�'kJn�EQ=���"h�"en�{x�W̚��+8�8Kk���/����!u�ǯDa�|h�X���ɹ�� Y��|7�y|~�A*j�S��9LO�����B�݄6�	���ma,.6j�dh�ѭ~bZD�%���̈m�
�
x��6a�P	�d��-�uR� ����B�\�~X�&#�Tt����ͧE�=z������=.�v�K��h~���6�,f\��PO:��Nm��"��$��h�'����pn��R����{�3o��N�{��.n�ʍ��e+xap���X�͋@h�+�o����X8	o�<$1��_�+s��,�/����wWR1��6��n�7�#����7+�/��@�wUVIAEX�UC}�1^�{�L�jy�.�	���ː��.v.�$���<��-�FS���&�h+g7�0�^̠#�wv�����\��I�=(^���I��(^��*J2�����v��S�⁧�!Jї�աb߂���)Z���@ާ�������/�m1���jg�y'�������	"���;����
�y��u�݅�%��C>������2�e�÷�v�ߗl*>�<�����s����$,q�!ՙ���sp��%�d������f)}XgcQ��?C�mn�7��HHD#V�}@-��&��&�O7�~�@�	;�aE�R���su�
2`HY�c��) `a8q�^�G�-#n�捞:;���f�����Lp��*Q2���_��xvH�L�c�k�~m��_&�ws 諲�C� �3�Ƀ(�A��������0ONһ��E��G���Aŝ4� |�b �%���~��\$�b:�6\HSl1f��]��1�i��p/ugs�Ɂ���qW����nd�m�`���+��LQ�%0/��)`T����5gK_�����W����o�4��V&�1}���`�����7�ތ�B���o`�vɐ����UZ���-]fH�ˠ��!G��=�>�oG��U�?{��6sYQ�d4���x�]z�5�:���sҏ� n��gc�1w��?1pb�}|��.E��tҼ��lDs��V�y���h`�ӝ��c{o�C�90�5b�A7�r5�+C	�o�-�F́]Y=�fy�����7��!�_4vm^��/+C����-��b���`��������;�<�#���-�i\8��3*�#c�J�P��GԷ���1�)��u!T8;���ô�a�~��n�ޠ�R�^a΅�%m*l5���Q�Յ�UZe`��Q�O9D*,S��H��-��#'lF�\[���:�:���&q�����ESL����u�¿��(F��QxA�ŀ�>��r��������D������5㉟�K�������|u"���_��G��]d��H�#�=*�`��1��7��2498\��@�3�`˛n#r���Lխo����hD�2���_D>�S�Uܷ&?�+�k��t=��!�G��5��6�3n@�!S--):
?������L���%H�R@��Մc�i��a�>���}�)������%��b��xg���g��J��t���2�'��Ւ��8��A\^"p�I���0a}��᮸���F�I����4�Rf;Z���w�#�9����"�^�>�~"���I��`�A�־#��t�I�����^�5TP��?Jg:��K(U�7���9S��	$�B֊�d����>@� |���ap�M;��*t����fKx��;'��.~�˞&M�Pa�I�J
bƓ&uV3!�3��k@���D«�:��������0��/Qx��%���b�¡�uw�@�GRz��yI�֋�q9��2ѧm]p�K�X���bݞ-;�F�z��r�C���18�� p��HAT�5���L�����@?�'�ݥ�~5 Hϟjލ��k�O��/���;�3���7������V�Q.]����3�����VO3� �TK2kͧ�'Ď�ڎ,_��X�p��p3AQ~�A�P��[�yWc�����,tJRj�$i�8���=R��^8
�7���8���HjD�T�m3�6�cw@o�</���g�kƅMd]J���V0���0��<���%K�V�_�_���T!^#_�kg�:�=�����8@b�TZB�¬V8��(2��%�g����~v���4˓��QW�?��f�cx�H���[u*��z� �K[���^+�A����Z�ϼ�jgX��U˩�5U�?G�	ϥ�XK��܎�/@�'͸K��K�nzM:�.���li�k@�K�(���1ĝ�*�_a�ؚ.J13��~I`W�Q��޷�`��#�j���˝�v�q �x�Ĥ��8�=?��e���u�r��ZI���u8O��!�j����U'j�)�i�Rfy��1Fl`�!1�`=�̽S�kdi�祢���F�����`9���ej��%`O��J��*���*|���(IE�Ԋ��E��K�®�8�Ps�/q,Ԫ�K\�?R+��6$�Kt8�K�W�w�ȚON�H=һ�4� Y5��J+dU
�f���}շ��4{O7��Y3x�j�^6m@�<Y�_(��|�+N���nȅr���zv��O�;C��ě�T�j#ސiI��/(�ޗ\7������ˏv�k.6�.�8� 65���%X��y�|Wu������Q����l��3陜w"�> �6B�Sz�پ�?�9�}L_��
��D��w��y�\�"�\�%�O�
ǌL��$5���8 �8�u��`(v�t8����5�%?)!���?>��;,�&%o�svq�t�Ch ���&�Ǝ�izX��a�c0I%=�*��d���eA�qK��sIݵ@�Tn ��"ay���_��P[�l���:tI���[�����n1�I��WǖV��yC-J7��W�,f�~��2������P_L�F]'U6�Z��.�p�E<��K=��˲�h��W�S����r/�b�p���l<s:!Oi��%��5AV��oDaZ}��/r���ӎ哚��#ϖ��w�ֲ#ɥ$L� �J "_x"gGZ	S�Ȣ4f]�� L�߆Qw���Q��V0���m����J2���يyj�q�ԍ��w-�A"]����/<��-�f6B+ѭ�]U���y֎m]谙��W�r�2���+�fw����M��M�����8�N�O��.'�m7jI�v�Ҟ>VřN�uC��o"F���al��!�H-���S?ԥ��п���
�ۍ?n�H�azQ���u>�B��cKuE��Z�j�X7]�W��B�F�Z���)��2-�zBr�6�*0�1PЌ�^L����W7���\��q�vJ��&�Oo�^�(Qƻ9������RH�.�[Bь��:�̺K�%��i�\l_�-΄ܒ�@ۀ[�'��	I��j+CtD"�(���k���p1ԇ��X�=��%�`}be���x�f]���z��J�4��<���:�R��G���n�Ȓ%�X�R��o���Kg4�,ɪ
9�ZRb�FY��h�D����P�B�\�l�N�˜5�'2f�(���ߛ�x��J��s�&E�&���썉?��RNK_@�~��j�����q�]�@
��K�=m�C����x�Rݯg�����l�j��,Z�ЀW4Ƥ{�_��q��M�$8�ԍ��y}$��Bd�WfZ,����
���F���� ����-������ϴZ�;�u�����?.`h�9d����fe��kIr�JVgV_w�#B����_0T�@�hn$W��ů������j�=�U��f<D��U��6�4��I��R�yXi�;�!>��u?�j�wy�\M�1=@ >�U�;�O���@X���-�K<�H�i!M�m�b��1�]}Ԍ��t��{�K�e�؅k������*v������J�48����(X/�7E�*�>WU��7�UQ��e���S"��V�t�[A��Щ_�}Q��n�>9��E�{^���r�Y�pz�=���ym�h����ϒ�	�VMX؈rD�/@�ـev�㏜�N�6
��HD��Ed0bP����I.7�����s��@ Ǭ�8mv `?�*�)�}��W<^|��hҸ����On���)R�Ө��&'~O�RND�%�o;=��O�o.A��6����.ل�-�w	_X����A"��E�oi��h�	^O���N����7R��'�D�9<�ܟ�`�H��S#t|f���@9XdBT�2��!�H^c���@��'�~	Y�p�uHD��km�z�k��8��'/�*[�n������8U�[=�!~��%-Y3h��"�d+[-9?"��w��S�mSr�}�ʷB����8UVӰR�Ή�0ogu�o�URc�mf�_�3,��y��������8�:bou��"�����
������lr���� ��O�\7e��2Q�wEv�l^� \�)�k�s�~��W�k;"�xW���c23(�p��s��I�]	h��)-����+��!7���
���GO��'  ѝ|s���2�����p]�5U���㐝'�0�r4l�d>
B�i��8y�¿%/3� ��V�zR�Ǌ��\��xH�{����c�FhR�b�V��U��$RǠ!E2(|לM�'����$LfC;�d5|�����"��q��Ӎ����Rǔ���
Z�$�#�O��U�$N7��'���J�R𮼺i���`�Q$(�ʶ����^n��@������G�2i2!�*��'�r�?#Y�9Lr�*�b�Jt�O�����D��,��y�T���<ަe�X(��5҉*hB��5���g�&�V�E7�M �RB��Z4�د�b���o�q:욺�1�?<8�{Pd�;�`i���Mv�2|��eS=gН�����Q ����}y�"�~�Swa̶7#CaTT�%$S�z��,��`�[��Hrk��16�Gا�4}�th��11$��c�a`\��E���Ak5#�a�J��;!NS�-����Յ�ɀQK5^�alࢃ� �� `��b<��SnP�:XAA�To�gvt�W��u�鵋�!�u�\��P��_Ĺ�EO���HhO׋\d�������D��b;��7�.��W�PK&��l�B(f�5cִï��<pV"��^z�Wz�4���d6�&C��^tE�0�[�N$��w�ԁ�d��;dT�rYF��i��p??�!T�Mr�j8��_p����_���W�J�Xr���g��Sh�w{N
BU3�H�'Q<�o�q�`��1���]�[\�c
6r�d
�zÅ�$��0L��ʔ���~�Nh�v���Ti[���+�~"T�
�;`���H���6I��Ga���*A���J�(��5i\���k���n�� 
i]��RR��]�6��d!<)��O��5ё�������͋��jr�������*��K�*�T��I�~Di��T�:ǃ	?ԉP��[əE.�6@rq9$aG��J0m}�/����n�����r$��p �ܳ�j�b�j+��*wK�M���\��(A��۶\���������_�qoBC_�.���2�2ʡ����S�9}v�|*���?O�B�����2�E�"�����S�;a �t�XU�7>3o��-���C�U�a[������u�2q'��r�J�����Ʌ�l�2�����+�T��K%ZUة�{F�=)sՇa��_�E�{^��zR7���r�P=𼰽�v22����V�?ʅ�˻��\����������;��Iƛ˜�@��5o�:�C�s�*!v���?��:Z(f��ܯg.W4�GY�c��G�R��ax����p�|�I1�1Q��{����Q����C5����=�t� $�R��^��L�Q�O4���b����ߝ���k�	� n&��K�҃��(�B��\��>��+�//�,��ǋ��������I���Xm��D7�|iPXg֦�D���6V��Nԃ۲yaV'��>�n�� _��D%RB߅�$��c��z8��uڕ�R=q���m��� QDs/m��U9�x��K�N<����8~֜gz]u}Q^� 8�*r����P*��)�˽O�k��'$��.�YWԙ�AJI���,2�Nw��+6o+��Ձ �k�K�8��H��:�hg�~��Ļ�)��L�����g`ֆWɤE��`_;n 	W=�a��=Ք�4:rb`���u/��_f.ɾ��ohM+��b0;.�b�6_H��3L�Y�� ����%�i��W�ϥˋ2~�*ow5߮x�B�2`��?@���2�8��Yg�?i������M�bb�c����iiZ�v�V�;��/4,������|�^�@z�s�v�	�>�v�՘�&$�#�7t����0�`�Srs�~���Lp�Z�r�<�5
+q#��6"I��Q2xٞy�:v�݅�.���*ݷ�9�W�( �N��f�eB��hhʭ	�=L;��@���<
��F��.t��S�G���Y�#%�҄.���C����k3�#�k1���J����$* G��ǢЄ%D�*��BS����WJit�}HZ-�<:3�D��?�@J؊���%�;�T�����z%�?F܉���f6!���r�*ԋo�4#�;Yc��C�r�q�W�I�`4kLG���wM���pRXx�}��ķ��_P��8�5M3���S�q���$u�mW��~#��P���~���έ���Z�W���U�e�G�;�T驛ND�Ρ���hǂ�5�_"�f��	�n����9ڲ��UY�� ��5�02�HyiZ3sZ��@�tg_M�.�C�`����3�@�Q9���p7%�+:�p�~haU\S�6���u:�Oy �ְ{ĕ'���{�&O��� �)��s���6ڌ{Q�)0�H:������`o���c�Mʊ�%A\g��O��E�i�Z�k��X4�,��f[A�V#���f�ߑ-leGU�.����'o��s���@t��֟M��O�-�}~3Y�����ڑ@�X� ��&D�=ؼi� �k����T��_��2��eO�ֺQ)�â76[$d%�����|(̏;y&�����`�}�r�ʺ:��o៽�p�=�af����KŰ��R%�G�%D�d��#ϥso�K��{�G�?���1���Y��/���
d���U� ���O��y��S��X_4�L�`�9�lv�`�)�B^7Rs��r�^�k�H$� �F�q�����Nd=Ǆ��֨Vl���l�Kx�*��<E�j��KQ��I$籠o)m�6m|슪��x��$��3�����.B��P�I�t�~'�<����䰰eFO2��5O���,:a�o�@Rg{��b�/�Tk���P6����X9Gfr�B+xhK�������﵇/Ƭ��I#��Cϛe{�	@��=p�K���]�U\�?�P��/�L�Z�/;#"d��ud��jy���h�� ��g'g)�S[D"v�b���[LQ����s�ƙ�_�����P�^�W�)���S"��į�8����i�����[�����1>ks�p�-K̦��d8��Q��΅��h��_9	��`��eg�2���:����Ab6eIQl��GT�
�!M��?z`�!��}���[���Vj�;5�%ȣ<2���e{)�rǳOB��&���"��=���r[�<ܩr�k;f�Z�5N*�����q8Ǧ��,.sV,-�&� �촡a�Aew?����nZ�N&%�����R��K�'2jM�VVVz1ږ��xdhx���jcb.��ˇv���t9�+���� �����s�^���du���ɡ���Uw�=����PO���:!NCK�t�th���� �Ɖ�#��ezm.�e���"��,�0����B��sZvz�\nm������ؔu��!��в}�H���NŴ�]�F\�W2������ �d�'���\��K���U.�x�V�"A�%��g�(�%D��?������#N<�]/|�PL"���u7#�}l��Q�P�C�!#��Uz��z�h�������1�m�O�1?�JaU`(,~��h�I��C�+��N~@��<>|j��M�i�F�pu21e��W�@TP���aRJ=�<��R�N�Й;��s^�ϥ�ڟ��{�}�Dw����ꏓH���G�k^Wf����a�y�M�l�X��
^�y�6��bo��p����/!�Q�1�Z�n
�k��]rtf��+�%�ݯ��ť�'���̮���h����;�� �	�Il��v��n�7���L�TѶ7�A���ParMM�QJſ�d����ׂ#p�`|,�^��DZ���p����L�������:G:u��^��0�c���2����'U�(?�����0*n�8&�Ξ;W8�r����GG��߲�q���S�9}�SF�:�n���@æ�Q{1u��K2"��@�37��l����%Q���\��)�i���e-'�.]�tĹ�z��_x�F<<���7��W>�oO���Y?���$��r|��� ��z��,^�F�Y�ki��<{����O�r:h5E�
�����:�Sq�p�`�E�*U�أ��f\��i�������Bb�r�2���i�~��Sy��QDԜҵ�JE� ��ݙyW��
j�%@󎉎�.BwVl�l�C���I!�\7�UO�F�Y� ٫��x}�y��zY�~�ʞ����������J3H$�ͺv]l�Dy���xA3����$�>q�03�_�#W�f5�Y�nF���_���XX���\��pg�1L�O
����!4�}�+���b�%��VF��s$�U�!?�Q`#g�Q���l7Kyֆs���a-Y�!��;Q6O&�m�k"Wg�X�ܠ5�,���
��w����*q��8��}��N@�,T�Y�j��
�߮����s�ϿE���{#n���1���pGkF3+�!I�C0��:9�b�ȶ����l�~S^n=0�@¦��e�Pnbi�E��!��G_��۬�D��˛+�3�wy%/�%y��\
uq2�4��r��E^PG��6�K��yl
��zD�.#I��>(wH*P{/�tG9�@om�#L��dg#��{P����rx�mH�Fu8� v��㋴��u��TZ'�$x�N������yg��'��v��?�x>5����iιg�K�����u�y߸Ѿgs������mX����,�t"
�!��t������4=��)��2� `��c�Vt�����\׵-cc�2��>����k��q�Nݟ54)�^-���9<ĸ���w忁�Љa1#E?����qj$sw ^�87�-�]������s�����iX�-�&IN�XR��XӮ��p��}���T�#'�?g�B��@�Q�Wu��2���w�י��L�U���	�J����]�_�$V�"3`�u ��
�0�o��O��� hұ�;`E��.M07�< 6P��0�"�ۿ]?���1%��rV��!��鏎��0�=lG��(�e�7;�u�oU��d�	l�Ѷ��ou6�'fL��s�?�k�Wϔ� 5gT��X#����3�F�@�7A��q��\srٲ���$�-�(��J�(����Y�Ԗ�Gt�܆&y�dH8a��$Z�����!�Li>S��{:�44��"��b��m���/��W�=���4�g�
�"a���sKfn6gҴj=�#��H����w\}���X༺Ȣ۵e6Q���H�_�ۜcs$�' I^p@tz?W����	��L����3�[��%��؆�]� �:���Nq�n��*��+�,���S%�-��i�*���Ҫ8�&oU�V�_�|C������l�#vR�W��%��ZLP�];�'$I岐 �:�@������)8��$1��0g$�/�!k*�m�cE�K_)+P���r�g�㯈i����W�N��j��;�CL��ˋ��Y��!*�y[�hk}/�:���u~�_+�#$Ȋp������f=��s���6@��ԁ����!JL�X�7U��`�4���j�:�#�*�C�|����Ǡ���Ԕ*�pb���V3���JV�Q��O��%v\�%'I;��X�~��𨸅(���|�)��ee��ӟ��Ϯ�V��:)�,�*�e� |z��pNW�U��?��(�Y*�h-v��:�A� ���s_êAs�9=�_͖©����8����*߫�����	�k�=^�d�[�V�?xJ��ȧ��b_Z0>��@��z�B�NxI�m�dTB�����]�v��~��}�SSӱmڷA����R��ԝ?~�(H��J}��)���k�i�84[�ؔ),����
�
>�/���7�jb;q�>��`T��DB�K��������vC�nn��I��.�)n�%-A>�LS/������5��u߀�E1��5!R\�/-��6�i��:��Y<(
�}D�-�o�oM�W+t�O4��\Zx�l�@���
�����$?��F��B� �4���gN��*$��z�Ut�q�D>�� �Ju�c%�${�K ����?/�an����x�VI�����e���a'��}��=9r�@����E����xZ_J���N>�gF�j��Yy�M+��'���cQxj�:?�֟�١�k���6[���G�xO��a�d��y_%+[ē�M�L)&TmP8D����9�#"kL�Ϥ�̿��K��0��}�{�|j�JMD.ԥBɫ�������,{S�HiH8g���6쌚�w��o0�sPǦ��Y��2����X�uc��O���T>Z�i:;@�)���A	�3r� M՚[�Ҿ�����xi^��B�?h�P��m>��&g�5`��3�5U�|�q���D}Ɔ壟�� �v�e���v� GN���;`.��F�Xh�%�*at&i|ͻ��d:��I�c*f��Y����`��u���[Rq���犇��I�ɼZ��?���(�è�m0���Zc����_`x��Kt��Ai3�S`��xEL*��BɴW4"�:U����������s]�	`��0��l ���M�a��} �ҬS���|�wz+��/�t�㢢��[�F��m gc3s�����S��g	bF�j,m��̤Gy��[E�v*�(��Fu�wViE�d��t/B���	o�A��p��t�gT��E2xy\�2��r+�hAJ�ַް��|o\��j�Nޤ�z
vҌ}�;fy��_��9��	������<�1�#5=�HBO��I�x�ı� ��Z'0�\���U�Nw�7��r�Hr���(ys�Q�p�Ȣ0۞9�a vj.��ԦT��LR����Z Ƕ��L@<�z�-6o&�GC��.y)��r��rBǇ��0p#@�펦y�T��S#l��6v!HH	�r�����`$|KH�o.��.Ia�#�6G��^�n� �.5��D�ZmX�:Ĉ�s��-e�����z���!}$����1�pj���xOg5�%����b�o�����_�&����4��ˀ��H���G9X�pn�B=tia��Y8,߄�<�I�4G�p}�sp"���'��l ���:Ql��{p�0	в��v�W�-��z����?iJ�S넦���j�����켵yA0�M�ٗ��]�����$`c���
k�����d�9��Ԓ�kG�,����i���i��+n��Z��>���i	�[5 ����{��d�xy!ΰ�S��v�?��%톡�5\�
�-�4B/}V��W�"��+_SK$���h�w��a��s������nu멯5�i
Ϭ�c�aք����b\r��hp�QM[P4���#��}����t��xs�����bC�����v/�T�tg��:P��1�T�����&qH����-[�}D�|'�C�����*�0]a9LRG��X7�*T���T�&A=h��FC�_�i�h{�B<8�F+:\ o/�EB]ؿ�#��D�ZG��d�vZe$d$�����Z�S��|�IBL�X186B�E&po�8b�h��B�q5v"�\�M_�L}Zp�����|�����a���/����F����`��45��4���2Ӥ2��CU�-3<	�1���{.eM:�IyiZC�� K�K�ɯG��f���o�iu��LB�U�SF���y{������J�Jz@�)�*��&��zX�j<����(�a���ܕ�R�Va����sbꬠ�L����x���;M�|�{�}��}9�Y��}�.+8�|�9c�6kc�J�y��-Z��G������0g0hjh��j3�8���I��>SUѸY����*�i.˝�7�S߮JO���mhex�����t7Ƒ@�fה8^�$X�$�]㣂*z���z"�3"�hk �h�N��.�qe:�O�x�\�v:%c�k�5�YU�ԍH�5 ���i ���-d�hIǳ����X�F��x�:�P�@,��Z@2�Į6��mw3#��(V0%��c�n[��Z�B�|��9M?�^�@1Ơd¬�
Aeb�/�zzI���Ǉ��C���G�C&�K�p{��l��p`��]����{v
^�Җ#�l���,$<�8����'t(����m߸`Pv�[0ů���MYc�ų���[�kx(��D��bU�]��0�M�Q���e
D�ց��D�l����I_�k�Z��#�=ж�*����ߦbp7	��ܮ��>�)�&d2ZA���gb/ҢB�'�e�&}6~<J���xy��v�+�
�/[��Z����Bإ5�0�"�66: ���Z�q�[-�;�1Hc9�&G�B�K�% K�s漢¹��pǃ�證wA�P�ǖ+&s;�������(��ʓ5@PE��6�7�HӅ֙���K-b��vIV񫆚���[_����k�4��++��/	�\	^*�C�(�U��r��vs��Z
��2�����P�KVM�Z��j4O"x�~�+�hj4;Ҵ�a��m�����aM��K�U��;���Z맸$��^Y�H�Q(�� ��\l�n�٩g$޼��U�):�Ww�B����P�W3%���yC�L��<lȜ09���
��H�Q֘"	E_�oN���$�ݳ�����5B�k����;�/����L�F�?O��k�H��M���^���4��6���RE6�UN���'��pL������/(��KЯ�t��Z.A���z��9����A��P���ye߄CXϲ�7�	����1�lxoiw<������54u@lx
����X��r�&�؜Dެ�?9�~�z��Xܜ�� YI�rA��Zh��s/]ց��q���DX��R�P��X���9��;Ǚ!�|}�H2Zψ���W�I�ш�āO�^�i��.��\z3��������L�y���ߔD=ߺ���R��_�K�M�������#�l ��b���������gQ,ۮ懈��T%)�;��s�, �#nv����P(�S��)�n�G�L1�f��T���i��D	R��i�AF��:
e�+��^�-^��q;$�����Fc�h;���~�m��t�5��f2l����1��!t -{��lk?FE
:�c���i�~��Q0�����B�/�� �c8D�40�����涾�?&W������94����x~�'t�r����4��6�c��H�C�+'PK0䗦Ul��8���f'�)*�Z	Y!I�Əb�3l�*lzo���V�T�ד�M��p�Vn��!�gRfYӎ��o�}�F=����+Li3:#	lEBp����~J��oS>m�7� TA3�yzY�CW�=��깘����8�2�g�~���\��m9�n��L|�l[��v�U	�'�d2(�ﴴ� ��'}:�c=[��v+K�[�'1���ے�acU�����"x�1�����_�c�c���~`��d:J��9�{��N��1;:�J�^��)kV���;ey��M&� &��n�끿2<f��F��S�ܵx&�iP��T�V1�V���y'�P!�q-�9��������]/뒑S��P<��j��d��I��ILuX���H��(�d�#�����s�sc�3wEi�z��	p�s&&qq���Ѫ�h�o8X1��>���an�FH5��b}��;<O��jOD���v��ݗr�)�u��ԑ��]1S����4�C��~ȀԶ6�������"P�@?�q�nld�$�oþ��ģ�ų��a�6�����m�%�=����9�<\	�n�ċָr�b�퇾~�����Z�Œ���}�y�P����o�Hp(o\4o] �4s�"Ye�y$�R
�R�0)���5��	�}<M1ԝ&�G�θ�!o�<�3�,N�C,��";�<���RLRG�s�	�E��pu�>߄/@`pɿ��ܟ눉֭{���yFl��)o�d���r�t6�:���
ah+!�m����<J�v%8��]�!�h�&�\�;�d��R�r��0����s+H���jU��W���XR�]����$�)�к��{H*sNiJm�l݀�� ��&�m*�2Cpi�M�<`��<���G��U��P)�O:5\)r��H�I�m�������d%�(�;-g�=��I�c��	�i��cJSw���]�^a?��1���"�*���8��d���k�y��Va$q�Bq�Z��Jn��~�!��:p�ͧ�6{mwId�f��b�眳�6�x,:�d�IJ�qx�o9�\zP,(���+-�Y���k��øp�ӽ�H�Լe�;����Da/���� �
eb˯���2xqAu	0�Q�ʚ��>ű_[�D�����lu��d0�zJ���+��aM�z�й��t���F�g��D-Z�\�V�v!���IF�[�U���c��Lu�U;���°��fL�ފ4]w;.�u_B�d<��v���}�:��I�OmZ��dgm����IFR DE�+��#N���%��T�H�'�(��Aۮn �\ך�z\9�Kx���_ˉ
��D:ܙ�V�Y��(S�͎%���8h����#�<yu;�u��[h;�Q�3���<���@t4���FKa��ڀ�Gv�āR�����H˰e̽6����jq�#�~3}��6$�#j�'3_)�n���E �b�}�~ �����t�<&��Y�C��� �t3|��j�E\ӈP� ����F����ه���s'R˛-��U�#�i�[���+-�}��0a���eeд�㠍)b�`ͦ�W��h�	��N=Z'�旸z�e��~X��_��y��4��� ���~u�Q�m���% ��Oy��x6����)���8&�x��0�kx���/���9�ĭmй��A������2�y�Y|�)�$�d�;燗��5��r�����/���h���4�8���=�R3�*p+ �'��Jeg�	���!��Ēά�Q+0Q�pV.
6�J=�=�����-���,j��%	�9	,z�{w��y-x�5�n ����3d����I��<���1~�_4(,��>�akj�!��}1V׃??�?�hJ(&��S^M(������gU����?�M(㛾��K<r������LHN��҃�V�;S_%�Ƶ�o�N�R�+N; ������$���DX`�f���d�UqI���ǌ�H P�;���7a$�1NO�g(���F�[x;EI;�U��b�9C5���#,:��CG�ԙ#>io���{���G�b5{��� �h.�/�V��hvI���b\�\�E�Q�LX��Me��c~��y� ���*/�֘�H76�L��U>_�i��1~䬼�W��u�]#�&'�%��3ʊe�y��զ)�v���a6�ѸI%��V����b�]ذ
�D<�m���GK�ELclB!TS-������t"e��� ��Bd-���R���[X�(yZ�c_b}tv��2�82
@����ͭ��z���ez�jw���b�_�w�.��5��|���|�����P�",�EU���ϴN��l7/�e�[�.��$�F޿v�)4V�˵��Lz���)�
d�Cp6zj�-�<Ή���N�
�5;f%+������%sxy0�����^#�?Qe��	$�z����S���Be�$[���;_���J���^���֢��=�!�Bke���Չ�]S�H�
���$��}��d=�M${x� ����0�vfL"�G^
c�EqĢY3��(,%t�(�� s�ԕ�*B�]BA���Z��N���/���t�X��L"���*YWx'!Ge�R��<<4�QyM��q@+��u�$/P��9��`��ڒ����/�]��T���M�����,=E�$���q��Iǔ+���
�h����.*�K� �M�F�Y&�Uꑰ�mϢ�6S���
�k+=��Tҙ�KF��ab��BT[�:�Ph�ǔ����ԏ�uWfά�{��������z�B�v|&y�����h�M�j��C�un:j���SM!�1D�~�̍��V���\-,G�@��@/~���b�!L�7jɒ�1"��3�w
�k-H��W���3	H���:g���� ] <(Fd*�$�Ա��ձ�7V���݄j#tH8E�|�"�.�kB1����@�y�kQ�:Hw09�Q����>����#��V�gRm}1{�(!ЁlX�����*�hOp�{�޺!��[q�����>L���� �6:�����\$1��\�+'ag�Id@(�GH��X�OnEo�XZcz��n�:P�MaO�J�.r���ϱ�D ���f��?`אt�sq���vG�Qlx�I�w�����D�B�NNtK[�y��G��)
�eD��Vb�����"C�MeAN��������Z@3�!��^G�B3��0i���_@�	�'��w���G�
!8E/a�qa�@��/;9��/�R>/sx(P���VI|���*3�:� �nv��*�t����vh�{T�7�|10�}-�
Z�^1s�ßp����ˀ�QO�F�9��c݀��p�8�b�g������c7��I����I��N���ږ��!jO��U�`!�g;Im�$j�6IWI	�!����R�65�>4����]��޵fA5L6�Q��Q4��2�"S���+���,%m�;g$�`,�������YU�W�D�Ø"9dpy�MrP��|r%.��zH�A�����A���\�K]��d�'�椖{��y� ��|ٺ΋�EJ����\�f�p^5�T�.��@%g��D+UN�g�ŕW�(�#k9��@���E�(K|8A�~ Π.+���p�G��4"�X�a��In� ���K�Z �
>f�tr �I����b�u�"9#�UD̀���A��
x��W��4����o���-P���J�,M��O��M�W�Þ=t�cGeA��WGVa�P�Zm`h[�ҩ"�vr�aM�Q�]�0��cҦ�,BY6��"�7$M�q:�QZ#s�C�o冮�k
�á�v�z�c�N���\������&�%/�(.y��l,W.���xNM��Z�J��=�������
����H�eF���II����6���Ș�����kav��/���S��@��>\r;偣h8��,��h)_�|4\�U����#���2��o��3-1�N_��u[�� 0	�6��_)׉�Z�u�e~���/KbS��r$�(���7�����l�{u>�u�42H��-�ݍc����52�QW!��r2h��@1�Co����׾N��6w\]�i�=b�x�n�����0�C���v����kv�. ��4����+B9�Ro����9��J�1T�]Ɛ�pt|_π���<�Lx�w�J��m1~V+��ʟ�;ɸ�TȴqL���!�c�
K���S��aL�v��:k���vK0��;��6�lȼ�ٙn����p��A+�i�J�
xB�0U���G��^S��D}�Vq�#F��XgEM���ϥ�4�Vt���2�����&�!�q��7�-F�T� �֤ �ZI%�H�9�V�ԁ�',ӏrx!�D���_yꬥ�|cb1����/b�O[����T�`��|2q�?�D��2�Fl����$[�>S�@�����|@Y�n�����&�Y�i8��m��!�= ���q����g@���_qJ1����,uTښ�84 r%/��[�aZ��y0�%�����W����stA��m#3g�+�*���m0m���:a�))r,���r+��Po��.!g�X��`fw����,p����1w�7��M���w���+��AU���E|3�g�9����YTM3�ק"����^��v��E�U�zx�#+ ^mƚi�8�:�=S�N�C������?D1,DC����l��f5J�Dom{O>��5�w>�6�V)%�^^lV4����؞3V�w�|��GG(�Q	C�K�A�}`��KW�6K�;w��3d�u!� �أ�lc���`p���AIi�
=��wd�K�ħ��wy`�ߵ� �CD6�D���[wK��uw�	�f��(:=��z���f��E��C��# ,9=U*�1���TQ��G�A��8�;<��
DE�?,�^�� CԔ�ِQr+l�'W��F�j[���X;Ñ�45ӻnĭͩ�֊��������F܆o�Cbu���Ը0������%����U@��U&�X����ױ����^�qB=�,G�m`|�X�>O���D��:vQ��J�v��-��7��;�4��hc��f��ī��E:ė:IF�a :\�#���W�\�E'R����(��(�uX	���%Z��Y��b͜�"�T���K��l�b����r�u��2�:�ޣ��m8���<ܥ�K;A�Д�$��h��B���t��UKؽ8dtE<��ۄ=�O��0��l�&X�w�g{�$�ݾ�q��e����� ��h��Ѻa��e��anث-�������`JXez\��L�e�|cՠ�Q��J���S��>��.��@<p���]~�q)����Ω%���	/�/��;֣{��@n�A���eU��&($��_��޺���zRE;�P���Ns���0[�{��UBo��'S�
�i��[�=��r�C��O��D.������:��8Rm��r��4�q;�pR%����9���X�����r[���'�-0�r�ӌ����J�;��X
�Ȭ��-��4!�ŗ�#�~�*UЉA�������-�-�"$O"V�%Tz]|��P���CRrWI�3\�{�o��Ա�&q��\l/�����YJ������LJxGFd�d�Tt�Nm[���r<�7'�7�l.���il�ô5��[`@�A�-����Y�>�@�t�oTi�%Z�J�:���Ӑ��ɵ�����.�܁�PR�%���C�)6F���P��⽼-_"�?����`!�XP�w��{7H�1���4���'�� C�����!e�$�����E��{l5�-�cU_s�^��;��@o�^��UGU7�\���� ��G_���������ʜ8k�?�.�un�SKX�q8��:���p�p���d9J���B�H���o��[s���\WT:b ɏ��bu�Z���|q��5XPs޲`��~c�S�x�R�yK�k�&�5q��T� �J�ĦбP��^�d�}��xN���� �d��N�6V@��-�#��Jf�/�3F��rW����پF
؍�����')�#���d�+��Gq�����x��FȤ��Z�\(0q̊���B��,`�����zot������NU�X71�đr��$�n�H��S+��ȴ��C��!\�P<0?Z��,��5l���Y$(��8Rb+�6��O9���h%,��Mh��O�.�Aё�@O&MK�0�|!��=��x��CS�|R͘.9�:-��R�p��!6�g~�{ȷ�MD0Qs�g����Hp�nͮ]!`��ۦ��RG����}Q���C��=clnZ}��dT$���V�� ��	[����gAx_,�|�;��?h��ݝѽ���_̕�!��	�o���1����~G4�;���fh�P���4Ί��=1
��'�g��tc���f�W���� �p^ �:ތJ38O��rE]����,	\��r&A/��q�[E��U��"������G���	��]"H=�p�����~)a ?���"(��T��n�>wЫDkY��k=�����czw<���2.@��0��Q+˄�*X�����Q�#�����u#��C�(l�o��Gvg�]E�u����8��a[���w*���BA����;_h�����K����������\�V�l��HĶ#�g4���m�h%˝��ZF��(.�FUm��enAcn\�{�g������EZI�>�[4�C��G�U*Â�o�}�Ϗ�?�=@�A}��|i����t>������st'3����h��]���s�sW�reL �0��[����:g�.(q3lʕRv�m��#(�'�(N_y�Z�����O��f�CzJ}�Z�����GlK�^b�B�*��> �zm���z�,K6��	
�w���'��R��䡡b����S��z��Y��g=�>�t�H�y3[j���LX9�]�[�ZѯS�3��2=��Fu�����m�D�F�k�іv�W�-��6_�\4 ������l������&�
�ݤ{��lK�:��f�.�*S�zV������$�� d��g�^�Y� ���@c2�L)�?��T��1&%-�]t8v�q��@ �mˌ��P3�����:���+څ���։ɨ��$%�p[���ܖ��<)��Q��c]l�p��ْo�ȱLK�۩�lX��Xt>��)�"��۔,�6��I�6�_kl6��˾?�@v��L&,%��{'d��)�o@o1�Z�p�7�x$�b���A�(��<�7ĩ2�AG�PiI�l�|�n0���m����e���ufZֻ^� ���W=Z����_w������8�䱤q�:��/�Kמ%�	X��W�Ÿ6&��9i�LD����ƺ}8P�<��m��y��N+Hs(��h>6Q-?S�� j�u�G�;��87�
|�K��k�F�
W>��
�q��q��f�z���E�O����~��u��bu|������q\�5Gk�'4��S|��
X� [p�x�(�N��n�',ǫO�+(hc�)xd�s���m�7���<��(<���ܑ��ǝe�1�5�7������Hd{�4��(p�a�c5Թ@�偅P����w�\ T��[���F�sd�D�sʶ�*��m�Zp��k�\S��<��(BpU ��z��4��u[�eć7�7+��2D�*ͳ+���U{E�Yr�� 0h�E�tٺ
���P3��܍���塦@�-xI�m�{)ah���w#+��0u�3��^M'�hh<�0�5�y�B?:�bvv��'�o㤛3^IK���q�����h"D�ߥNg����_n
�+�t��Ʋ����w7&��M��l�Pf�Y��j���8__L��t�p���Jg��lw��(z6�Y��P�P�`�"��vt����C2��$�sxאַٓ.�5~�:��`��30����T�5�n���z|(��,�m)����6�	|�(�`�?v�E٠�@�����W��p,aq��Y��@��.W=uf.�~�_L;��{U�uO�^z�t�9цR(@,�1�m��!!^��ܶ�p����Z�����Ѥ�N����������Z0�0mc[�"��ªU���Cbv$%%Ō�iv0�>/ SX���iw=��^�����l�ܨY�r[�}/%�G�M�y/����h?�j�Xݰ{���ˣvLÂ�8��O~X�ٸ����O���ݾE�����>�Z��Đ3��7�ޞ�j�;�~�e �R���qc�?b���B�yY71��J�Y!��9�@v��`���Fae��+�C�6h��K�ސ;�A���4�T�8g�@dn�(�ū��X彘�"H{�麐��V�ഖ�:$G��{�A'���x�j���te`oSp�ح�Fui�[i>�q�nU�{P��Q !����+͋�%���*2����G4V�%��J)�a����h�`���E��!Z�S�u/j�t���oO���V�c��b� ���,k%�%wR����T�::)B��5�-�J~8`��aY0�w%�:����L�:��5WUZ��'v��K�rw��f��5�9��qM�2*�V;PH�\�Ի��!r]<-���������%67a���wRV)?��,�~���eۡ(= � ��~����D� �b@�y�~r��H�M�T_���ÖD\����Qޣf�Y�̌I�w}h�v����h������e�`&���������{](-*9�l 	�ɽv!���N�:���8�6��B�eDJ��0���,`�z��u�.ՠ��՛
�6���n�-	�Cw�7C��^|`���_=(� �ֲ��
��wh�E0���"�v�.�d��p�9�T^K[�HC;aG4���1�`�sv<ǈ��po��^+7��ǌv�ojd^p�O��ď�g\Y�v����B�9�Az�A������H�����U�$ѷwL�0P�r�)WoM���CX�Һ'ā���@�7y�}L:�������f�aK)���"W	�K��_<k��	�����Mm	Gϐ��,�X"LC�g�/ �!L��$E�7�@��xhЄ���i7���d�LKm3��`#�R0��c�6�����B�GBJ��\�����؏�RB=b1�	a��~XLO���0�TB8��(�ޤr����h���p��&��-�F�p�n;�l�֜8�յ#�����cҚ\�j�@���8�!��;=��֖�
d�`��m����A��"3B�!N���c�qd�
�� *AY���*�K���б����'9̫(b,���+��	�	w�����2�a2!���a�;w��V�Y�B.LQ�[��˅��,����e�u� �?�~�4���y��5d����^����ɾ���`�j�? ���Sni�I�O��X�g:��.�,`����/�j[����9/5r���6�~���@
4Yqule
g��F0�٣���>A����������Ҿ�g����(���i��,vn���n��h��t�'Z�^�7,����s�A];Vv43�)���Yr�s�A�IRUm�"�&S���A�¡� #MP�K���ѓ����6yq�-��+���{�W��R�E*�r��ّ�m�rN��L����}l��#w��˘+<��N�*/.۩�MlSl�f4�0&$u$Kj/��_�IR�~&`&�BFn�XP5�����|t�����`�/6wz�wD�ʠ0�F8oU�DԘ�yB�f�6k��V=S����4�%�cj����Ѵ��b��P}4O_Ƹ�p�mK��w�!�6��R� ����g<X�K�y�*��Y���� xDtB�����=���9���MK��&;��V��x�>o�s^Q��h�T�D'	�����p{��;����0�|���r8�q�	I=ho����m[H^��PO$<x%P�Q?�"p��,}�ձ��<cXϳ�h��
a,�}������ �h����rP��� i�wi	��|��.2���<��M'^v�.��#����n�sY�"�W�*T �һ-�?e�2�n5�7�=���"�[P��������v$�W�7t������K,J�:�_a�r�%���ʸ�Y������ū]�cT�������˞DhRf
lEYP{�TyƉ�Vx#iHS�ю�������qyOhw
�R�ݰ��7��h�k4���̠�A%D�,�Y�0-��C�$��7XQ��p��D�$�y�>�D��uc=����)��A*RCģ��˪b�aR��rq���L88Z�GI����j�r߶��K{��	w�Ԋ��!�}�y4����9h�W�9K�o��o�8�n�iem=?��vm!�4Jy�@i�a4;���w ��[��_m���Qk�Q�p�s���i ���-�!*�b(Q�@_���4��(�fH���0����-�,��C
p˷]qƇ����YD�!U
s����m�������c���ҥ&ŵ���N���o^���*�i@pD��A�d*��0 .�o���d�Ћ�ݐg �����)l�{]���c��$������C�P��"3fK�^:��S=z�^�q�FqFtV��\x�e�����Tզ��Z��#����_�����#�w��_j;_C�U�O��LT�"\����g�đ$�Iܗ�Fa��iɮ+F�2�DN�C�Jʼ�r��l��1k����C�����[�� L���4J���M��6H�]Sˮm���/qFOԿ=|����N���
sn%�ﵭBE�;8�/ z��Ʋu3`*�S8Pgy�9�~�,W�n7�Wd
%pՈ�P:nSB%7�nGm�e�
�F��`�C}>���3�G(=g��Ax�&�d�( ���^�f�[՟�pzk��;�_�L�}���bM�u���p#�0 3T�����1ǟqPp͒�҆%�<j��F��˶���;���NRQc��ԧ �D6��)T���B���D`����Z�Nm�ך	���Sx�<�>}̌���?�%.�G�ZY�2�0ܲ�PƮ�3�hSKP���<i[2�nn���~�X��[��;:�/�v������Lr�;���$TT����Y,X�X���f���\e�q�a�"R��7��v~x�P����\.N,�@�b�����������.�n�HW �E@�Z�rh0�YXe6#Q��C�"��Nps��8?�D�N�=K�M��	�Rş��Hhfr|��@�'�t���L�}��ޘ��s��H�Y�\����H�*&\�f��{맷�LGmh	:{Ky|���z���}��H��ĶN����	�4�[�uE�&������/� 4C��+=8HH4`��y���b�#��ci�bD�99��Z�߼7�� ����{�	 0�h�4�t.�lJ*՚U�s�d��^�52��۾����ek�'���ȫ!��`�z�.�"�
$D:�Q��ϳ�v���RO��/+z����ÌGm=䚕�Y��
���D����*�u�p�㼷w+�X�6����M��2��N���Lf�K����j���؍���xt�����>��mv�?���9,'��8�[ ��$�+��;y�r��X G3�����2{�Q�d�h��UH=����*�r�{U�	`��&������疻r�Q��>�?셰��o��n����a���10IEH�-��h��a�����|ac�1č�CD��6�!}�����F����~"��/ӃdF/nn�6Hs�y�U� 0��2a�Gx)�s[/�V�V��6@nI�[;)o�"~!J���cT�l�T����6F�ׄ��EX�'G�<L�s<�8��'�>iԸ[�x4Z1S%��cS	�%���l)�6�S���<��L����^^C��������a�j�x׹����Ek�>b~��d�f��#2���z�2Ns���P��S�X4�LV��?�<��r^?y��#Dw��kX�����Ab�C
 q>��(�?�.�`#�S4H��ԛ�(%�mq�ߏPh�Kţ����K�<ͻ�ڐ�&��������=ВV2���G�	�N<�L�(�� �<�x�c���0��dԘ�#���e��ǎ�@t��(�+�4x��fR�'٥5O�
�.NC-�p(r���X�;�\��*^�P���I�)�����Ǯ!�R1��8�������ZX�����}3f�w��At���+j�����? ���@?TZ��0��!��r�(��k?kV�v�|M�Q��k�G%j�=@$�cJu��<@�'�u�O�����%��bș���l�
p�t՟ȓd.5��OJy+�b:�I�\�	�$���߹3��s��kF�Z17��V���/'�X:{��OIq��1+�&�/`+��L>�Y��F��,�����l�	%� X��6��Q��'/�t]�PS�!�/�I���E��߱ �( ���c; ��a5�.9���uz|R�	)�Yͯ���6��fJ�[R���d:��S�r���l������cb�u�R)H.��M� x���E�f��g�n�����d��R�h�X��� fk3r�!����]�@����~�l���Z����F=�a����"Ƙ߁�D����~6W�#W�*��Rʚ^D慠�c�FA����h'���!����ґ��/�§0�+����#�6��Mx�,����ߧx�N�0`e�n&�c�)U��_��F�b����k���Tr�l�H��;A�$q����-�������z����W��C�bT�N_.B,���(�5�4/=��`S����4�q�A[M��Mr�g�X���!�� �h��ڝc,�*�9��
M������$M�&���~I��M��ڊ��:,��
uM�F��"N ��~��g���ҽd1 ,��+,T��j����0�[U�).Bܴ�Rh#�� R�}:��=��j�3,���lK�4.Qzsd��i��X�\�k������w����Z���8H1�Z�C}�E�Y�{���K���6��Z�1~�Fj4i���V��q�t_v=�� ��R�H���eC���(R��%ϔ%/aQSz���=MXTB�14:�܇�,�Ca
Vy���X����.m&\P6�� U\Z�IT+��!��rNk��D�e����聚L��q.���K��Xx���&��E$& ����k��:���7�X��c��F���I]��h�%���Y	&?��	m���A *4T���Ů��d�pZ�j���Qw�W]�2�|�AzP�߭�?�Ğ����];{phÀ�kp�.B�I��J{�ڲ;H_98|%$n�+�l|d��?������p�~��6�=q���w�s)T\B����<8�Eթ�&���$���Wh0���=^<_.*��`�4j>��i��z�V$#��H��Ay�7O�R�]�����w�GԤ�[Z�{r����&;�#���H�~"����D�~��_D��%d�����^ы�|���^�r�?~:��F�V�~�3�
8�,��LD�s�,���S��=t	�(}K��y��g���m��8�ws!�MM�C�������H�m��h�M���_:�D��mW9��1Y��k4� 8�>���˝�r:������Z-C$FՄ�!2��}��Q�r�Ŕ/���#n��"��1KDQ�U臫K�aLV�f�?���.����#9��1v�d�����ksӍ���J��'�0�I4���
����ȥ$��|��Ѝ%y�Ǆ��ǯRb:�{��Lw0{�4ᗧ�.��J#��-ٟ����Q��]J`�]�X��O��x���ӽc�����o�`G�%jY�	�w͙��ߔ[5�8��'B}!�*G�]U��B�lE��d,oc�n�jZ������6���t[�q��no$EpcO=''w�@��"������v��������������k��@d��g��O�/��b�h::�Աam���#9+)�I��D;�򠀭]�wA~ο�w:Z�u�kZ5�{��?�}�gX1�U��<\���:69J������7u߶�1��4O��W�Nz:d����b���3l[Ņ�i׌^A
���{;� Ig�=�&B����|���u*�;�$��>��aٙ$�oU+@�Ujx���NK��pvϱ_���=-wZsZ���xU��&w�� rw�?b6JB�y�^.f���!l�K�gxfZX��'q����b�}��J���w_��=2�rU�@I�CX�T��!�KF�{r%�*�O���Õ�/��RL�e�1�ܡ*`�p�5�+k��?1��zxji��hY��"�T���G��P�5?,�ձ���9_NJo�"/){��� �*d�GME�T��E�1��k;�XB��4N�+	�|�]�H�`0�� �>+���'�<��"�<�ȧp_���i�r�Z��a
	�~��q��uH�*���e(���>/��J�Q7�QD�A����oBL�o1�m���U��o�hY�;���� �ɮW�I�K�e�w�Ci��k�H(�ou��9�(7�/|m��ɑ��#����v�Kc3y�x"S��.�	�lE^l����*��f��h���䵓1 {�ފq�sXs�5$�Hnb��>��0= ��k������,�W���
�I�ш?/y�����?�/�V.�z��ѰX�q-���i���L�&�k���Jx����?��+��t��{��/�߄&j<ݝ�ɞ�n]���֊`@�w��'�,̈E���� 4�;�VԵ�����.7W�d(t����t��PKh;��&��TT����݌���'mLuC1����o�n��**���Y�c"�v1fCkc���a��b�X:,z�'ow���n᝟W���2��^4�^���9M�7q���rs�L��t�d��o�y�;��;?iq�ɤ( �Sg@�:��c
ax�o��ڬ��_�+���B��`qO6�	�y��Ter{���):������]ӽʹ��v�0������X�"���1r�����Y���}XxHc�x�t|c2�fwh;�ڙ� ��3L��+9�U~ncI��~l�هY��/�g'�1`�������) �qW���5J�Ĕ&��[�ʹX�%�Q �_�u I���/Ǎ�Z�a4?���"C����r�r�ri���J2��w�aޡ�#nx�T�%��؇X�&-�����w��X���W��W��3G8�T��qK�v�F3{M�;�ݗ��R�I�B���z�S6z���X]��t���:y��:�J�j*`|Qy}��3=�S�p���M;��쯅++��D�b�4�R�p���A�D�en�t};�f�E��d��e  �Lξ%�4z����?v��������z�᪰���0�@u���au�Ʊ�u�~���ݪ?�}�r޼,�b�H�����s��s5�JXZd+ ��w��z]*�'Me�����E�	�����P����ר��\u73j	�{R�+ˤ2�=������e�?6��m&H,��S��
_>R��QkIk�5�c.��Bf�8~�[��d{�z ��چ��:#���Ѣ�T�7�Ytv���~�Hv;��s�͋��l�X�<:D��\�� ��+��Mv��<�x����h�ЪV���%:��&���ҥ�5��t.t�X�L1_햹�B��B,�����"��Z>�}��~4�iSB7C#�2@ޥ��Т� �]�D�s���I�c�A�gj����g^�"�����1�n\x��b�~��Uo�J���Z�W9��fp$^)o���dT�*���
��7�>�x��}���9lf|��%�O��db�$���DL���d����Qe2U�6���׉�"�,����b���e
�̖G�+��8��.����$�ؖ��S�jǣ=H�ﱒK[���8����F�lU�1m��eѺ~�JE7��@(��� ���b<�����^H���/�G���ʎ����&+��W$?\J��S���b�*��@V���@�0?#E&�b-(�N<�o��c�P�E�8���i���������{����?��@l�.���]R�ʺr���,S�����Y=w>���-��H�5
M�T��~�Xk-Xm"I�t7��Z�o�jv;�8����P�N�I�/]�q�#�ɝՐ�v�IF�m s�q����/��H��+[�S�/)ŏ΢0u�w-���BP[G�~9���6�^�j-坨��#�0�yY���C,�Z5�`����X���"�}�����V�U���s�I��;T	�ONPg�	fyI3� [�k 9-nUP�iS��!p�ϛ�693U��h31����}[��[��\�v��t�t2� "�˫?5$ኰ���E�Y��Q��KQ^�K�i�S��V�,����Z�0�Nct���;���]�Un��?΢�h�K��=�����r�`+Q�';�L�d��q���n�y
�rx�;�"�:k���٧)����|���4�����]�����	}�[���	B'���K݈@��6��J��ܐHV�X��L��߯�r����`6@h�w�x����6��V3s�$���õ��)w��W���ׂ�3��j�s����%]Qu�?���{��*V�:�֠7@<�5�Sqt�?mw�"qҷx������1�	l���幂$�BP��3}�xm���)ӭ��|n�<=��aA��&[�����f=�x�� :��n�X����Gf'�SQ�����C����ȝ
u�N���`�yW�l:/�#~ͤ�y�;���mT�ţ@z(=�1�u���Z:�*��J�J�ˆĢ�ϛ�AZ�~�td^fO��ݳ��QY3�PWb�I�٠ὡUwсqN�m�����:>j��pN�@7��n���D��@�O���2҃�g*yÓ�YkR�{�L��E�/�cT]�+���U��s�a-��8$o��GS2SN�<��}�G�JU�|v��(I��}�	�=�xM������뻈0���^����2���с��8܎����_[ǋ����~ˈ~\�h�i�4~�A��.fg���-A�[�~ڊR&;6v⺨�(e�Ǘ^�OP��1#�Y}9͝a,�O	�S����:�rww.[���aG���J�����U��[�w{H-T�O�θ�R�"�����*y��T���s�5���-S�F`�u�m���i�4шa�i$�V� �UO�F��Cl\\����VL�:Ŧ������!/�l~�b�ؔ�]{n�2�l��(ɣV2z؎+u��D'~&ѓ��@X^S,@7O�<-g��k�Oո�3��g�_�ʲd3Ѵ,zR��u?-CHKI�Y��c���;�n3���tg1"�;����:��.�n���Lvs,�6�痢�\��%Y��gо�����Dj4^�3�6�%��&6O)�m����2�3� �\{t�i��r��E���x4x����'���9{c�\8�����4p���qRx�Rc㸑_�Sq��1��!rޙ�oF9ʰl����󰱶�v��gH�2�YCpA\i�V�B��o�b5n�8�s����]����<�/�{9Ϙ18I��8xC<�w��c**�O���'�ED�<�5�ML:ɼ�d4�ɭ���xP��23>[�J��|΃-���; .�Ѳ
�=�V���h�^RE���Q.�{J\g�}��J���N3;��t��Iz�*9�-a�aG��?���'7cEE��iB8b�D'P/�o�ԗ�C�!�&)EZ)�� dd˪"���ՙRF���,	>S���Lu�9�MC�(mG���MWT�RqC'Ol�y���-��Fc�vH(�L^H��b�v���>���d�Ы�
>���D����_��p�_7G������˙��*��m���������G�ʑR�4��P�w*)�I�3�a\}��H�G��������.܇�ŹmKʌ1�����U`�r�������c��9������h����m7F�]�K��ʤ��#��5>~�$<���l:#\H+(���d`��V�l�@4��Z4OW.�|t3�9lM$��wJ�'�k�M ���e�s�����A�b����D�\�a:�"��)����{1,�Vt�&ʊ���R�Η����U�i@��B���p#����D�� �,d<0��㷀���o�!���E��bT\6m���7���[L��ǉ�ek`ZhjԨ�P2���\5v��l����/��
���JI�B�ol,�TՃ�I]���K��Y������\ ��k�K��yf�d���Q)���Z-�#]pe���KzP6��A+��'t��ZLejc�*y��V�����
禤~ΐ#�7�����q`b=2/`Js<�R�6��T�S���!ҡ��	)z�%lc��D�\5�r@���� ������ƺ�qG]���:�/ԚH�Q7*�����a!��(�v��]?* �ZD�bq�.
�q�c�BW��������p�q��`����KP���a|�0�fbwv���k4:Em��P�>EI��e#=�L̛���T���D&��k{��8�8�Ӹ��e�b�&�ue2UtY-$B:K������}s�e�ݤ�y��a�W�c�,�rQ�Y���s$T�=�V��z��pl������&��br�-.]�	��᧟�+�J��J �'t�N���c�t�$6���H���({�rnΦ�Go�D� �*QW���M7�Ȏc�U!��/rL4�d<���-���铀ŧ�Wv�n�g�U��e۔��j+�=��6�(-��'���Rn!_K�93@,�IدϦ�?�k���e0?��j.��� �!8�\�Mb�W{ES��F����>�n�
g`�������&�*�}�Ѐ/OP�:�"riv*�/ТT��j��mA���r���X*E�F�n��1�F�m��,�5�u�	�L��o.��iԊ�H��n(�4�v8�d ��p���!�cY���G�5[���pq�=��e������-��� ����՚�����Nd�����B6�mFs:z��J���5��;?7W}>���-؟���t���Tl��p˗cXq���3���t��/8�^b���#����y&��むQD���=�i/~e�Y!m�Α��Ec��|��N���S�iFj�f�6�B75l���a�������P�KC�fmB	�}�{�Cm�`�(Spg� �8{{��o�����TQ����o����f��&K�٨~�g��5��z��s�������a�L�0�	,�aY�F.c�]��@m�g!@`�B���|�s��beRЪ~^|a�f��	?��~!jb��{7�B�Z�>���o�(�i���r��|�x��)�ye�L��Х�N�X�y6�>���@�����c�����C\���S�r�C[�������CC�Wu�OE�'�*�i�Z�~#�(�w��� ~����5v���u`��mQSV��#� J/2���E�$>���i�^�I4�?R�z����XG��X�jΘ�T+k�H���V<P�tog}�dCW�;����Z_�]��}n��0�Ẍe2s��:��	�>��ߩ���f�N�m�:��V��Mۗ^�z,��נ[��y-�?x)#��ݘJG�5���<�8�bhp��Ү���v����=��G9�Ԣ
;���'�;5�F@�������2c.�0[q�"tQ��v�F�X�k^��� D�����ѓ	L�G�_�e��W30���h	�}�T�t 6�6��Ϥ7�9HV��Uu��O�6�� ��i�e�8���)��1�fS��T(�:pv��"GSCWjkw-mӄD]Q���y��V8��Ճ��י�����v����n��8�]�Ip�������4����M�^���27K�'{yf&�֋�ީ��bp���4�7;s6 ���Z,��ŉ�<��>��+
D������YjԲƓ�?P�A&��M�?���a`#kB��6$#��E��ǽα`�|�Y�mξ�~��S��m���|�^/���~r<�4�$�-y|��H�O㹊<��sX"�EY�V�ֵC1�.L��g����Vy�	���T�IG.Mv���Z�x���n���8�\#:-wP��ʫ"%KT�tp�W|��0T���)�gz+P�Υڣ�^lAͿ��P#�p�Π�-�7@(� ���M=�"�������-����杯��<nF�� ��^uI�@��5x�AF�"5�Lr���20( ���,��;�2tF�&����:4���@����M�������o_�����ė�����!?����y����]��YG��KP�ﴤ4o]]�+����[a���g��Y���gv�-ԨB�k�z�!RAW7aw���ҙ�1N�j�̞=J*A���/���$�0p�����3WԦH��%�70��)����ea
b�3ྫ:Z.P S폼J�֪��ؘ�mr�����o���������Y �daN`�
��L��$��rM)E���o��I�RE&8}J{;
]�S@<v&���s�$g�K�Z=3PU�E�m��^��Ll�ͳ������\Km ��w�_Z>�ػv��FI������*��?���H��B�� �H��]��܆�L�F���i��<:�P��q�W̙��]��9�]����-\�Rᘳ�y�Z�Ĉ���8��2pPsdǍ5��!�H�![~�]�9m����dJ�A�֙8���W[�5����_���6���О�4 �zv��Q�� ��)���@��P���~�ph/6�ۮ�8"��aR^�kBd_=i!��}H8rWtqc^��t�$�1�%X�ן@ي��#S�鿈>�v!�؁�m�Z���R���s_3YK��<wvX(��}�{:!��f#�lA��i��O����=��Y@�o7#D�5�K8�яs�.�TǶ��[0�_�y�c��-�L{����a�p�5D%m������`"�қ�E��bC�\�j�y{ɗ�~O��C�[���U� �[��w`��[I�w2���Y���R�����������-Ug��6���J��t��+��I��i'h$H9�$``�? Ү���c]HW�ܟ���,��r�EOT��qk�nxI���A"֝��E� ����Z,TD!>KG�����;X �Ԧy�5 ��V��"%喌�����P#��h��	c�9�ɖ�H�0�b��&;��]Q��y�47��4��<��F��`�ή���Dk�0nn)Β`�!�����_̿mc�*���E��F� �+�W�^�s���#�\�3�ɨ�Q�<�/������l�u�[��>�'KCK&����H�ik���ɂ�#��N��<\��Q�Rg?��;���.E-����rw�J�LG��L����0�9�J]�Vɥa�)-D��omǏؕc�`�#�;��?N����
K�J3
��DO�e��ߨ��YQ�aqs��s=oc��LB�aK��K=�H�RE�-�L�� �������|j���sh�9ɱ}��Ds�ל����Q�ɣ���˷�j�+&L8vo�`4���ۧ�ҎB[��w�$rj���|���K�xC���w< �ϥI�N�J������9��Gem>�p
�s)}�sN�F^y��a���]��cx^��"�R���T�c���M�8z��b�i�����E�Z�%I��,���rq[0�PŚnD{������E۞�I�Q-FJ��^o�Y� O�����w�m.�l�O�����"|�f�d/����1��Y��)O�Y0�1�f��l
u�s��h�C�}�kFӧ���J�L�����D$!��=���R���Qt��k��dl*�N�_�i_ @��M2��^Nf=]Eq�o�?��(G����K��{e6��!�Dx�]��z��ϯ⼄M֩�k������܄K�&�E�I��S�4.ߒU��@�h�K�%f!���E�2�'y('�FWrR����RB���T��⣌
@S��P��-Ǧ��ȃ����s���a3y�]��*&�."�����__�T ~�Dҹ����O(Ѯ�9��x�Vn'rA��0'6y|;/�⌯>�G
~����m��.�Jxe�ڱ���������K��Rr�G��c�D>�s]N(��P8�/�K~p��3ɱ��V��l�|������F��G� %���]���[�9����H�
H;��*0+W��u�Pd�Cg�3r��6�,��d�����R��mM�o�>��c�Î�A�c����{�Y�H� D�������}��A��e����ҽ��]�v�k�̭�9gQ��@��$ d�0ъ�!��p���K��:P����k�Y:�ϹG��)���BF_���~&���@H~cv��"Լ�?$�T]G��-ib�]�W����v�_ �
+[��5�R3����LZk�^�I���<m��������0By�nl���*q�tļC���Zc�Y��@�Cf��
�u�pcK���EO�no��]�H��0,2���!Azcr�,�!�g�6]b= Z�g��!�W�	���2
K׆K��d�
S�6E��/��E�EFO4*o��>L��!���'S3�n:���?��G�HqWM��b�"�$VK�EI�GyG�r�Ҥ��<Σ7Gz6����������񲨆�ςykN�&�v���%�ib��������뒊�w�G}��/y�=(s	���ZS�����H�̗���~y�w���#�X��.�L��$U�J��4����n	�R�^�P6|k��j�-S���d��ʩ��7�8Tʒ��;���)!��8o�N1V�����߃��B�hگ�9�G[|.���l��IG��^��ƻ�@�gsXp8�gb�]$/h��4��tLdy���B?\��,!����G'"A�'6��B��AX�Kb�F�@�3�Wd�p���g��M$Ox�U.W�� ��V-��>5}b��S�����=0�D�!�����l��` ��W����LǄF}�̞�*!�x���gFxt�:G� ���Ò�n!ӻ�U6��S�1�GJ��	oT�^"u�Zo�t'1$=Mb��8_* 1j��IBY���l�X��U�)r,�ti�!G���)�=ԧ��e���!
����o�ʑ�@xg2��:f'���V�������{Ye���>����,
H�oEkT�rN6x55&�n[E�
t�.PGY�6������&�+#�U!v�g�$�;��=	hWs�l�:T8V+�b���LW�̓K��t໭��C5��,���M5�Rg[��ri�몡��^� ���_H�[���j�[�"����G�s5H���ry�¨�Xkc=���z��Y\�Â	�{�DNXF+��e髮'��10�߲K�]�v�'+,+���I����`�/�K]��jV����g����ꓥ�̍��������Ra>��{:-z\Le��R��;�f�3R󒼫�\��u雳��ju7��gYI5�~���{��d�=~����h�ӟ�K;�o?��f�N����+�9�M�\���0�zӅ���J���j����ɏ�
�r�w��-��Ј�/�v�	`}w�wJ�=�9�
�fnn�ʒ@�%ǘ��S������,���uژ���8@�7���2�F��.��O3���(N9(�*����Guc�g�,~�c�������jer��\�iyOR�VC���	0Q)t���5hi���U��~Lל�uK+X9���Y�^8%_�5`�N
�����t����LQ�\gYp�ۍ}��I����Rs�Κ��DB��\�gA��Y&�]!*t��za����h$�̬��JM=�����\�9��85��V�Od�OS%���{=