��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���<Nv�wЊxNXT�>����g��az��\�Ҕ��w�N �p������Bh�n\"��{�0� �wrç>�Lb����_���9�R>%L��a�G*�BY��X	�LƩ�J�:YՐ�t7��P�1���2ؗaF[��",�	(Bb��y���4����5L�&H'E�|h�}6��I[�1_��?� �Q_�G(5A��O6nP�U��7M#6�~?�P	_��xE��gf΀�S��dӼ?~��jv�_��e,��n��D�&�#��gU賜Z1{
;~G�)�/�x���o�wG���r:a��;�%�s>r ,��h��þM�دU�7�8m�B�*Lk
C9�H8��sO�	J���J�$��$t)p~��)���v�Y��{��1���N��_��(�����t����ف��dP�1HU�9����ngR\⷟J`�H2	,���������7�(N�5������Qø��P��#U�[�*�Ycܜ
yx�q������Q��s�6�Y8ȃ�p��?���\��34G��Ǆ��E��ar�=��qWy�O�9]h7�O��թ�'�27|�'�F<�9~l��{��9�B��TF5�v:
����`B���F=мP4�����K�1�uyrU����)�P�<�4S����JGN��B�}��ֱ�.9qe����50G�\28H����l~f��I;[N�Xb��PmT���`H�7B#��O��&���q��m�_�cz�|���|G��13rE	{Ğ��8ť�gk�ډmy�Br�s��ې� �2��������9=���9�´-���F���؉��s�d�s��aT��h��~s�Ɇc ��L�O2m��o RfW-�	1w�Ζ���y2��`��v��讋5�ã<�ۏ�#*'7v�:y�=y��lJu�{�.���w&���#���L��]��-K�k8
k���7�kp+)c��H��
5!����6�(�����h ���z2X`��n���R &{�(��qV���Vͮ��`�AC�n�WH��؆׆o��h��W�ߠW���ya���݀�`�p�B��%Ŕ�����n�=9��1���:��t�~������Z�o濟npp�d���]~�*�k|�����w��8�c��gd&Nf��5����Yw|���-��� ����#Ё�om�g�*��`ֻ��	m8O�ɴ�pe�� ?�j�g�оV:7�D��h��栧�s�"&�>)$aq��(��2��_��p[���h�A��L[��:-�S�d�-+�g��5]&��S��3 	J"ި1Q8{����KhC
:��P�z�:����<�7��6�;��nm��l+q��Q(D�G�9��lJ�eϡ٬_�-`�R��u����������w��$s��u%,O�������lՌ���52#�t4���v	���*��_�yN��@�Q���ZAPZŔ�3mٚ��%��K��lr�qi}I���M�~��t�hs���Z���%��LgD&��?�Z���%	!�a�L��X�N�!��᪠#5P�$�zl/������u�H�3�C����J[��c��(l5�'��u��[U�G���a~H�̬\\�����;_z�A����Ǹ����� �=? �҂��7�ŭ�/�[�}s�u%��{�2�����WoJO���^���06O|�Ne����vm�^M��<4�֣N�l�) _�
e��6���C�o		��L>�P�𺬽���G��^v��c&J_;y�s���1Y���V���U�^t��\� ��+T	��o�e[5&����;�Q�>�F)N}�|��t7
���|��1��Ǎ8�� ۑ��#EV5��^�_�B�\鉐�����%E=�ι�07��AG\bz�/����s߾�w��񑂇������ FIB�1(��O����0�=ȫ��G��u@�6BP����8�ۿbvO�}6Kx��d� �ަ-J�}���i� �4K7�A�S/L��OѬܒ�;H@_�;%�PSڸ�G��2Ҿ|]%�A]�|�hIT��>%۸�]�h���{w�\�<ڎ���	�e��a:|J �P�Q�	�=*��ܝ=�J�����{��qm�m���g��y�^HUL�:$�έ�r�����b�8�􅬬��U������T�14�_��>í����b[���0&���y��;��Ԧ�!D�����>�z���=��6H��П�`�2������K�Y��-�E(-"J0[M����'EM`���w������".7�ՈA��N�{��;��6@��C����2~(�uZl;���(�`7T��M"�ewQ�E}[s5])N�yv�����P�V�W E�����CZV�ܕ�罎3�=�A6��i�=^�A!�}*P'�P$�9s�O�:N+�1��.y��o�TUGõ͌���.�ǩtE|�v|B��g7J���H^R�~B�����Y�̽^l��
������$��[?!��n�����)P�D@	�Nqf)����Ht��z�.���O,���H�k�O�U9��4;{�H�B,�W����0j/�sx�:#?�'�P�N��'�L�vqY�H��Xy��z�r���Y���g���U�k�ǎ�EL=���at
5U k�b�bd*�g�S◐�>��%.<�gϑ��=bDX=��R0�l�;�F�@�^������ Y �,>�[o��-�h���^�9�o�����}x������I�X �{؃�1�ցѼ�Ƃxv�s0���3��3�)����ʰ�8�G�����e�MN�h</��C-V��{j������Td�B��a��۲)_Bs����~-�t)F�S�6x��D���J��?�]r@|a�z�7�q���S�:ng���P�����NPo�'8����T(��d��ƚȯ�m4+�qB���V� �3�wѭ���
��1d;�*�',5�p}%�X� �62b(�E���4���+�},����N������i$��A�얫��_����s��W�d `�)W/��gBh��DCPs�d��jv������a����^��0:4dF���!avn���}*k�;>�
�ю
�m_:��y�(g\��SjR�߻	�5���x<�9d��gˇ$l��+U�q����L%~����@�F^��s��%&��Gy� _	u8�soNd��q/�ļ��*b�~� !�8:&��:KW�$[�d�t�g�xx�V�=�W��(��k�#�t}UO+(��el�����R��5HȽЈ6Zqpsoܗp��'Sn�nEO,�+�8�yp�pȊΖ����o���iB�6ߢW"zT���K���� ���>g�:!�L�%�$�;�
�� ��&~����if.�0B8���L-�v��V����G<�pb��,*\��At�`���0�G��T�H��s"@����]�s��T���#��1?�8f��+#��+�Ȳ����<�حKF=�*���l�ݻ�~{��l��!��r���r/*�=�b��vw�'�l5Qv��g�@����n4�G\��Ú�5M�d��8��tD�VU�Ϡ4ͷ���ۣq�u��0~ED�ՠ������:�V�ptOQ�egYڪ����	:�i)}����΁�{:U�� c��{�7Uq��n��=��� �H������
R���LV�Pzz.�.c� �Gn����bC������p�c-EۂQq������ �h
���hD؛n�-W�h�Zd��_Ĥ1,s�$���f"\5��sه��������L�]G�ǁ���ߤ��Lr�ʫu6Z6��rrI�P-ܵcg����1�7�>�]⍳���ODF-�Y��՝7���+���Xm[��eV�%�A\����P��G�i�q3��l�3�s!�O�����	Zi��A�r���OnB�F�<�t�ǈ۸��1���U�%��%^#*}u�Ь 􀐞�vO�_�ц���d��Իx���VÊ�Xr0�n�alAՃ�]�-��)��`�@٭�\�t/�_Z��N��K������^9\�م�[8�T������;��2^Jz0>����*�����K��\^�AN��(����I.k��t��n�0�h������1`9��vXf��C}^յ�rЕ3`᭡�nɒ�Ĝ���J��@%�b�C ��fр�|�e:��'$%ZT|�Ѿ�	F��H>łl%�o��� \,j��$�^6�:N	��i�N�����3�*�4vE�ȃ�����H�Vq��kU��ᚣ���_�EȘA��w`�����B?���C�a������>p��+��?���PeY�����4IzZ&�����.�Esq�io/i���%� �Э(8����L�{R�o/��.���KFV��I
��{g�l������E׏�]l[ee�(���c�Y�T��MTN�^C@,�O��;�q������A$�IE�����)�\��ev�Y�ZQ��L��#TOnj��GRR��f����I)ڗ��2��h��8p5��'�'ܸ���wZ��a�'q�af.��z�E�/����	z��_��p��=	�A-��g]1��^}d�\�`>����	"�R���Ψq��nu�����<T��Hl�7�yv6ْB��8��u��Q����NAzf�����*���V��V�s8�OX(5)f�� ��k�왭�o*:m��9�Xʂ3�vJ ���H�
9X+$�\���e��7%q�m����	��'6Ѧ�X��Ki�v�|W�1�f1��	� �Y�?*���:>~]BR�#�ͱ��x
�'�ܳ�F2wO�'L^D��v�u�N���j��#���ʹ�7(H_Vi�-vg�pΡ��*��$ ���i���$�H0��~�j��h�lt��2	����Β��4�����mp���S�kBHd�޼^�ݭ~�\��-::o�jY��C��O���(���T������ye�c�,"���������uʂ���ߝ��J�%:�>�%�aO ��4��h�n���_�� r9MO�"�z��j�]�	"�L��ŝ�wN&�!��g8������1�����
x���	�u�9�	j�Z+� L`�A?1�$F�򐟆'Zcv�	D��h<�fa�y�,����E�:긻9�h�3%�%Ŝ���dAHE��'�J�x�Ě�E�Y�Z�>]l����Quh|�������T�x�ਙL|3'x{aXV��E+�2Agh�����S3��|Vf��ؽ"R���?�]U���h��[�Bb1G��1�+0�p�֓A�9/�׫�::l�jL[�����I�b�ޒ���R+����Udد�?l��fVb�os�����d��ǫEW3|!f��Wf�/YJ.D��)�٣�}a=�-�����?(�">�W�;Y�@BP���2}��p�����-qV]8ب_m"~d���;e�����O�4<<?^KZ���A�l�)v���$~�#{Fg C�6�RӟM�w5�_o~8���R����4���G-0"E�b��hFn�q̄�9��>F���N�Dr~b��.ߘT݁5��9����|�EPH��9��$�^m.e�'_f7�o�`#NJZ]S�ե�����I2�m��)'�C�� �׭�ǹ��� 
�u9w_6)��OH�͘Ew���)��<�i�`��.U��4�SH�!9ej�
��.vZE�e�1D���� �B�4��C,m��57�V����q�L9#'���ԍ(t����&:�g L�^�䥑Z\�F҇?^R潅���kX@)J&aK�a�v���	WUKO"ۖb�~�2:;7(e�c�3l�)+��^��1a�7�R���GP�ɥ�r��#�%:�Kb��3�zxToi�Zx p��/%1�8��E筈�r���0$.�f^K�1�#	wD���#�ar����}��rE�����]�Jp}�L|~�7Z�5TE+��0L�ה&�1��
�K
{jƏ0������|��A�Z/��3��&j��_*��߄�ψ�$�d�\�?Q�7B���s�ng��=��k�ʒ�;ft���|`�5�/���N���
>Sd_�3�+I�~��'�|�I�܎�u#{A���c�~RP�_�:�wл+ ����d7�;�c�A�F�$��,t�Qw��
i�M����T���G3�3Oo��}A�A���$��W��4%��'���ܚܘ8��@���]�
V�[~hD9��ʠ^F�j������V�h�D+1��%f���`q��Ը�d'�1�+;��)InY���Xx~@ld}G�GЭ��B킲 ��hP�Ҷe�.�EC3�]IԌI\'�+�)Ωm}�� (�${2>�N�<��-�}��f��GB�cq{T`!2�O:��!���/��n!�g�{X�[�OH9�̃��H7��/�1+b�(�n{몜���,����p��تW��MW�sׂpS%�n�ϊ��}B�������Ք-����[���QG!X��7赜�y�f�ymH�o3��s}9W`�nl��Ay)`Ȧ=5wS��T��ā�c��6:Dw!,�po�c��?�!ߛ��`�v�c9�R�OMit��x�R����i=���}��jf�����e(�^ur9a�_��x�'*�)�1'Fm �:���h�lC'7��=�IYT�|�+M�i��W�L�{���y]d�y�-%X2��K>>(��$L$[%�.�$)8�Y����錋�Ż2�������uу�R`*�� �%�\������n�c�:ޢ�#�j_Y�ŵ�H����i�!߶��Q�}d夲 �j�$�g��
�v���i�-JE�����ѐM�C7C.2�R�e�p��`]W1
5PnIY6'3�}Ud��+����SJ0�/w����x�V�o#�tx��PMĦ��=��%p��:�Y�*���&�йd�Ӗp�-��u$xtR� �u�Y,t��R�\�T�/&!D�|Y��'7���[>�����{}(�9�����~x�g1�d����~�?�U$<���S�{��"\H������Ǽ���DYU �	!��e)+�O�6�3�M>�n�y���y|#�UJ)��`�K����L�����/����&B0YBC)Е	�Ї����Ѳ`�'��@v� �[�/�QNR�����Ɖ�×o���G����E7q��"Rۏ���[N�����$�8�� n��GCl ~Au/{9����E�$��*�j�s=�
�moTS�|�9ʄ k�����E�۳"Qh-'��d�;r��k���L���v ��j�8|�!�<�O����D����A����|l�r�w���\�5>�Je©��Ym4l^M~���י3����^H��?o��E�I���i>�3�p�m�ӐE�-���-x���DHP
��mw��*�0���-���C��������&9jmj�=,I� <������;8�/iu�u�{(��⭯�CsO�q��*j-q2H��~$;1�qPU���y��X�$��
ywmg�[ۭv�޿^z+$n`���LxO�|�?�u�N�'�!�d�7;$L��{Y�W�S�ݠ4g��	(2���H�bfg�H�C*��#