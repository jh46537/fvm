// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rHU6+r8Gae8+oo3U7ZPawP4Vto8ITdssgJ5nserk5atGOo0F0b0r2fmlv8MrvxEb
7kJ+fp+ZMBwRhf2kb3a9ERM48cVcEpUz8lGywlO0Vit2U1lOLcogtopHBZglblkH
yzbz8fM7NpnGU4C7CjgLMq2wLMRr2F4WtfiU8Cv4i2A=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15216)
NWJAdYVI7IQq9fgc0QiejlLnKBhEAsfedicH8Atu1wVTDaVBWNwBlXPdfShXFEmG
Wa6Pg3hBJoQLW/F4XcoQ/feK4jPlHWFqwbf59vLCH8eh6luIs2JkvX3xPsgeWeBS
HPKs4kSvCMYvdjI5a2nfTQTFT27ZpbdFnqNfeBzAPdLetiw0qjWzlWT+CJatgnyU
8rmKtB+5JO2IOZcZlWpCRNbA/zUQi/dBxrkPFPrsa5f6feEDBrgZnddzKLzlrumH
9d4pWPCm50Xyar2iYcJeh/95TsgbC0z6WwRIGJ86uHhNadHHzZKC05cCcRtQTSIc
+8A8r75nP1SRIcJOmxFfn+7tNte3ThS/tPajLTtFhzLpLUxHq9O4SX1PysOUtRxq
nTrxjNZ/Y0g9aIe/XtkEpRZaQCKk1/nxlaKUQ008lHY+ZYSKWBdOQRKSWKADAWhU
G3yDgUgrmWCabSN2sSj3a6U0FbKNjVqN6SYXCs9IL+BcoaEVZeEgmQ9Igrl+Z539
+QdRq3f2MFIKrp2s4OS8GT/sA0Xph2RK7t7ZgdbJ3+vohuGNLP3c1ChktZn9EnhL
elQuLOwY68lLMEqnEkghzKjv49q2ZDtgUaHy1FUacWxp9WypD9J2DHPsgA2LFYjo
Dn5ekoIphRxOXi46iFxsHD9Cu4pNVBFSx1SKJNGDFimmc9toaw+DopJ7FUogI6ct
E54+VySNnrb+iRP3HG6nWzKUrKIZYCQqylZ/U8jwkfJlY9qwlE7kHtJw0mDhrXtp
8LqFwnJSAEuXICn7Ja0nYzta7A9yTSAxAAUMCHccZSE88JU4q2lhMugA0KLZpFxs
NCI8hJrnohl83k5mcE86duIkozjn9jcUSK/+DUbFru+EzTmi1nHPSLP5Bq85U0um
gEI/WvuO/TJovFHNq6Vl6SwkyDr0nfTaqGQP4E9n39nnvTKr6MiwgIbJ/IeZEONA
9yUMeiIR7Ri7VgWgCzKS+XZojSi21ENeX/+Ce9sHZodiD3IyOvfUa/c7M7E/wOzK
8QqBs3h9ORDzylyVoXz7dsZkbsOjMdqmy0kMG/aOfSQgDBJG4A+irOm0SdSGerZb
G196Rn98q6gxq1saIzhbEF6QK04DTci21ZbiW2IbUcVI/XyHYDlFexzZAjkQ2vtC
p/W21aMIifo592U8VLIgKojindVQXULD8UrsWWr8j5DU943bWNEelMI9kG9Uv0ra
aTPVWxBvr3Ci1R4dYcFJbLrcES6j7UAiF6CFK1O7VpTJTZirfg1vZcd6GpQXSyOU
yV0aXrgjY9Rls4+KxtjFNqqYsQG8vGmAxFklsvV7vdHpn4QOQeulbeYnGicj247q
EBo0q94AJR/V37ewbXn5z0KIoXXNJ930I5f1+lp91Dvg3XlmMbsN+xGugDlLSHRT
I2BhySTsmPIdlR6cAJCIdjxbg4hJNSbnrFVKJU3cNgAlNxgpx1T+fvwP9qMOL2WI
W7kj+soMqYjKylh2BV52c4YprN9xvZfABSBg9RUGQgmKgOrwM092WRkPVV+4LOHC
WP0RNga0k3a6DPwO2BJ9gq4yTjUNhrnsFDmls3cZUjZzjLYdDtgfqG5DykHFUVVn
HAh6/SWSDsjoLSuRKc4SQGx9Z3MHSnQbxUqpXB6FjOk2qHHlGvxCgIoA1nEj17ZM
RCkcnf48LRkvB1+XdlTEuw1WIyt82RDHdAZIgOv+K12LXFs9Vqm+toFO5DIOwMrl
DO6D5ZXwz40s3VhUgqHyGjx3xlulSPrtEnDZZV03tvxP7Ep0fNRkMSW/kkVTRMoI
7JfyxImsE0stCh6HZESiAACS5FxYWYkYFpjPpLRRHMo90HobVWLvIopT3SRORuTr
2C69/rfvJoB1+61ujmYjXQIYiCyvHjRVytyRRFl9WjTzj8peErNEXcJTrCfOqF0w
uHGcpK06gogO1jSbCSmkVlp1JGvyUSy33L3O66scpt/YaPq6a6mssrSAxgmEqLt4
HPBIrpYus6UbVYwh55TD1qtBTqQcfA38PNWnSDF6GLMEAh90uvnnexOD3ZTKkFy9
f+7ZQgnLnp29jP/IHRpRYz4QRVZ7VVSfLxPm7AjLeXeJXEdfWTYSgSw54Imhfgm3
ILqZN9IJqTfymwfcaYtZGywIetKAplkjzpQWZSylH2Mq+YlX2XSaS8225ZyGBnL7
Av9szdEQFET3GXCK2wCdxy3mkDGi7ArwhGE8Qblja3nAyiug/ZVU+QRqWdTpEMS1
3g+loJC1PmywcwKDOVy3bjoEkJotZeZ1zvjbx6GsCkXsXojhgsy9wDDJKH6WJoa+
RblIQaPLBjoivq7JIOXufpcYntQf9ooZWcdv4Y0zXoFcx5CODx6NZBCUYQo4gF9H
D/Os4WLnXqu8UXrJUEQv2QcfC6wqCSy0pSRFSKIjytQUWqwwxhAlR53B/zKyInVm
HCIMTEBjJev9qppkF308AHYH7AI3/AkU3sR3szI8XSMgCivgnV/ISy5Tdh/g+II/
jHK/6WUCGbfe8VBy/+3Rfgy8D7OcQy5mv4YN+Yrx5q2sSmSw8o2jGveIQJ8mmqL3
PwiAzS0jupLM+X7TNrkdU/eJbciK2JtFX8AUd/4XzOylklEFam9GM3PYEn77rPG3
4siB1MT8frwbpu1xDcic1sIip5PoPhf0aoN0rpPE6ePYf8gLUeTFNNRKRejVmGr0
FyWt1i4onM7rA174tbrvdEgGac6gPM43iIqOcwdYqWr31TJEdqeXHn8CCmZpyg7c
BsJ28C/3JUBpFJuwcwr4w2vhulPbIsxceRfwglu76g/EbuiO7a8Gs++a3SChS3E4
pL2t7HRFb3vuyHxO87gmk5P+2lDzEVifw+Ik/0JHvMa6JDenwZbIrEkHdmU2hqXU
SIYRefx+/I0vZ29YxDo0Zs6Ytvp2X7GKMmYZdvrd07xYBl9pOxsthS8CM4QGVkxK
y8JjUf0zIUUhYmGajgb+aVOl8X1uIPojeiS6+Ewr9ghRL5ua9tcnzLl8ia512F3/
1NaBxwfDbOqFt5XywqGPtQcWDu1bxVtnZSXC9s4kUw1YO7tYoNpIiHSkFADdmq6b
9j2HQaxW5SsyJWeYKdqjbpkoRDYwioQNH4u5z6c8+K2D71JoAobvgkloYM07tMp5
G3U126kD4890QV9nIptUvwv+4eucDRQuvYixrCLuanW977b0dtYUsLItj++q9tR3
EOL6xxm1CDUt7/8oEF2NtI/YGh80TLUOW9bNeZuxioWXlxgzU3Vtrp2DK05LUVZA
/IHU7hUXs0RBszWQzJnf/sEKDEkw4OLEuvbh0FuePlz2BLh0WVydA8Qml4xi/lLt
4g+ud5vN6vUpicF13KSFbGiNHIIJnFfbAhNKCmkR1/D+Jv6CKIwmZalD21dKraVB
UZVevtOJPnQ661qoMmhKnNcdAUjyNUI4pBSCqHO/AsTCYtR3pyIdsp3EqDhjzvQp
TWoKJrLvHtynEiqOZcVxckZMxq+jFMJctnWtqLqxHHil2dWw/jGLufLHZHIxpAgi
LUYZyhUFMlbwuL1bACW5KGwpNUOlbBhVbLUV+xtACDqzlkFztBB2wfR1y7462Rrg
2rt0fCg4XFeT19vhHfbRPEqUrldLBw3wnymp9ycMyliysdUjb9QwtLNA66ht98Ej
wbn63LhhrWZJpa3Ao/J61OvnYSI4vxTIQMY5ns0arodhjCBNEQ0zTIFK+cwcp2rx
n71Ut0JBogMJj23XtOh2lVnDHO/uMe66YCisoK+tcYdF+cBZfrx8z8ZevJUVzsQc
mbSlqCRbAhFm9yu4OLH7zhypGEjkyX2VDAzJE6vLWlwIuh4nRoLcfkvzrNTRHOwc
U5HuQlwy2GXpnLp+0E9CM3eYyCdSBtYvtdZ/FbvqkMECSXWJu4TLY0y8QGqtX0hC
u1qPiYN+6IcnM2+G65+0gfgsx5IQPf4Bh81x1uzBSXfk6xoBX4ZyLV9Sw6tpTcRi
QBJJaiDnaXoSV0APMKdZ0tdcCE4J/+QzomNz+z/Rv2ty8W1N9mbzUCt8mdPawemB
dY0PeYIfeN46Z1iifFJIaot3bdFO4mnnFrk2m6HHU3KrcRH4yfa9TcRFTDXG3h+6
fKUGPf2LZyB4nwBSNZ8sPQaiSyymamXTtkmqPSEu6IlRTKbMb7auxPYmzonaCRHV
nIR8EwQOhkUY+h7RJZABIb7EyMM4GR/7eCazL4XVs7u9H7lPocj2N0A87grRD/MF
iergvcY3mprOh4sBPPnF6WZqMtVW4ngvbfm9ReCDYaKMw1RXyTc91DPFm4Cg8cgM
5bUIom8IWc3rwrHkWe+kyR6T93aG6nHTVVmZT5ovnK7UgcxnMiyohgW20lmQZZGY
J6d3J5USA0yj4gT2jh4YATjxRZcGs33kL7w+mkGgGw0tNfCmO4zURxwjuV0IYTcH
7mhk83RkJfbPvEU2+YQANEq17/xfnY6nL/GdoiXyh93h0BCRXNn0/i4c52Aaej9q
/EQOIq7D+U1+GzSjEYQ88v0RfEdX3SKvA4mW2RVJ5JGnX+GjwwVd6w8wVjJuy/iA
bihvcf/j4boQzKquQ1YaY3p2bXfEoOQAhWyK1h40QKRN90QLdpblrIfhLxchPa71
LHUWed3Ues2rpnopOrpdmUvAVmpJ23j7+xwbULXakKqw7D2A4ui8D/mY3oc+K8tI
HSyoD2WySlw/I8VRBpktlQ0YQy0jOS7Zrm6+WhgW5TJUmW+qRYojzKW9SLU/Y34A
Ke82a5Y+ucjqxbQ52icv3kvTP1QnRqu0RjmC+bSZJuZX3khoSuVTFJmUtxLu894P
o8QOm1uw/Ly+BB+YJi1TZDXwQ5X2k9U0f00ihiIOLoGBuUdcoNH9vYFYM8h1BJ+R
8lKLsbcYz0xSjJak/2zvDo4UktB55CUWhqEeXEslfLKJvhxoLM6Iy/PkRgNbGGzj
zKv6rh/A6/ZWg6qAtX4oVqFK9lQn/RRyzMPkOkBB8i1EsUczkby6UIymB9r7igkz
RKcYp5yz3kAtNqDkZF46cnTe08ijfStP5MlaCQW6dUDshfqJlv1nXqybgidCI0PZ
HqFYsE5KXokttdPlf6rdZ4eH6QIW5JKxhKue6HlTtB0R3mbrw3EOXLqfG0VHRGsX
BU1JAwZ03BWlt5qWU88+j4TBpWYkA0pQNGmwVynGkQii7wK5nSkiDwankR8uV4f+
n1eqn83+iYGyTfEK7oRiwsl5WjfLIDfPilIfMxbQN9YDlDm1gytwUr3DY4LOjTRt
aOSDBwjRZ4w3mEQ/+ANxfO0uH7iIxp6bh42hJCRukcJOzCPIFGoQj7SzQrXk1oAM
u+VFoE1a+vDWPLx4Y+tCaK4i7xe5WGmBMWx+zDnvaUZgbV7eEyVTeC4rzPGKtRWZ
EYcQo1U42chWZ/eVbHJpx5ZPssrvh/E3CZQ9CysH+uASiBRfJUM0f1i9WTekuKFN
pFMhHUCg6QkUIjQWmTDuFl4BmTzhUgmy4/hUzKdJKnuYUK0JqvvBOZRBu4Ipf1eV
u0Wr4hX8tz1ZYR6nEsxPCRDtpfl7nzpJHdORQs+yw94P4//lgN1NEol4URC+5iOe
azWxb/ivgc2Iy7S1reSX6QvYLWJtcROC6yQ1kzOd/IChuXogU2hFiZ2JQTY3D7/4
k0L6b/5hQaDH3vyi3HL9TFdrPi8M6E7+s/g57F1iQvzbJVTzTXYT1+87p2dP8A2k
bXxQlPhe3ijzTXGnyO1rWav9XFTg+5cwzO/BfFkgCXvSpHx/ffHCDtlmjCcrYZBO
5r1nd+s7r35WxsEb/sK0WCsQr8dc/TuAIUNJnooWlRwKKjQfOiNvfn4aubtnPxqY
Cg1tzuP0MATc/DJy0VVqioE4Yq9LKR0yRxEGgJ58zdImJeTpTovSru5kh5B7XA6A
ycFbVXVB7B2LZZJ/AYjEmiScgSBy19ijMG4H56xnmgc6oBcsyUKB7ib/itLwj/n6
wO3EPs6DkmkghzpKjWyDWUoyeSe5/sqe1cJWPJsWXFbjmkEDU4+hgqg/4gUoYXR+
ljKlGcmyy9tzD6qQmaawMIk6GQ/H4ztHNY+KbF/bYYemg3AIr65Fdzb4qorHTufN
OeZQjwWi1tikq+fEVu0jDf7egktIr6NtxvD9CslbES13WqkQaxZBoHbqTjSfVmY7
vpR7DR19owXXwBLJ2rsqE4sMQ5K0Qio2KowKspxDmqU8p5eAqu8sj5LoMkmoM6lU
TKCgFf3e+e8eIs8BGSpSFLAPOeAJuI6NCha8FEV9s10FIBtJfDD1O6cCWeS/Vf7f
3p88NsQbzwnjZm9WZm4mU/PPHl9sZh/D3a1/MJOPzMUEIsFR1P+n46TbwNh9ytLy
7PhF62ChdxWstROl+r2ahzPWzyiSRRcGJFhmynBQM9hMfRi3CDL3UKb7GneQHU7Z
ky/Vh4R28GhfATZM8Z4M21aaQ8sW3Caf+Bn8Qh629t3Xrdwk69k96xKd4L214XSo
nnsUL4tC91EGfm2eu6f6TrPCOLHXr+SOFDAshiMx0VRtvPIBbSmkC8ca4lpK49OE
5leFyBNmNFEwYJoTqyNR0qxecnP3qiDiO4WtNb0JxXE5OLtU4YtI+ajt0IK7nFLJ
1ekxTsQvo5qgmZNz1kP0wRQEgXJHJY4f2igNomP6ZhvW1GCaSObH9wZ/bH1NML9w
Z4rOrATcLOMXddeYTWp6u4aZdYMwV3ny0+j+3zQeuS6rdAsrRFQkeWPOQXLf7vi6
rSf9QZXdd3qocd+XxsRBpKu8vmJPlpr+D2CFfiEkWF1hwxgAGwCSsbG+K9MsVShD
Ron//cVgQ6SuJJOKFi9MnESeF9MwOow1gX6kpvqD7Oxj6/N7Ia3cSLIoDXnWXn1w
zve93Clpsh0dgAhRukTQGOUrA0bpqpjj0L4b1aUgotOj4W8qiN/gC4VL0edlGjpo
d0U/2wca6uDvmwcqIS27uTQCU5DsViu/I6PDxwVnXZ97FrYLIwcAfRlA0vw4sLp0
0JW7ESBdiClZkL2QVhARwEJcVyInPM6M2Hw3E9VV4Odk8jCGa9m5WZgjk3kAOyRi
hetz09mXeAPccf/8Ogo+VfgxQP8ppubutRjWcZbal0gI+I3v04LPaHHDUPDDTMFK
jrFsOlBhHh+Qi0oydxMsRME6IowIfGSdjVZnxKKFsg3Btnf9bWXh/M6mw/mZbrBc
RDnh9N/42WhOr6PUbMqghpQRxxkVuW7+V06L+fGMnyakeVnTwTSm5RfW20JdbyFW
fdMiEk4MUjKfjz6oEuU5WxW+yovJ/2S4unYN+NrOgl6OmAawvhz9deQURReJns6u
tUs8OaaFX4k/P+GR861EaBA/w/YWIW2QsKiayYn0/0c1NYIoJIusoiI/YKyRL11p
r9UyG0Rqs8ZqpBYZ9XGjjpJ7x4kPypf+Bs5zu60psPigwrUtCddUQPP0zzGQgLg/
J8+9HOMvzr8RbhVq27ZoLAwf6iCJiMzFod/nr1709yRzZdRzTVKBcIQ3bGYWMKFr
Ynkp+bwBDF+4NZUtXAPfL2j6QlT2X5YrjrQ9pC1qg0gxfOIn+pfhgi3UGOJSGiRK
KObOLK094tP+buIsuqV6fgv7lJWZeZV3PCJeVTIeQPg3FWu7sVL253C38BYgwtbo
R12bXJeAbPi2p+/SLOCuHKTXUAicr6Yz85E2eV4U27AhxAyn1DlVFwR9bywZsqyr
cWX05/jWQTDHrzpjeJDdgwTTIwuMYniq7WVlVmR9AaTRzLRnoIrj0//ajL2Bw0GR
a29BhFvE3xcTkkiJqpzbxELkQN/Coi7ESZkxZ4o5JII5vKgWvI3wMbk3d+MAk1nd
rwGBKh9spaJLUdYuFyWvodHcc+sFcbgMP25RD0bXCXgdi/MC81+ri+fWKCT9oOSb
iUgq3azl/1oz5f99nN0ykezzgXW1noSxviDoTjCyDEF7VjtB46ytZlxIxqpO+eWf
9NmR8e7d9nOvn/OtBno2VZSihS6dUXYJYBe1LXtD6crFhXYNT5nDEYozyxe1iNzj
FK8uCnNFSMRr3tO7YvzQkjO7sxIVLenNidK/FcF4I2Fmgxyz/c2+2NLtruQ0duv4
TD4FE7b+dQd095045gRVhtuuLKbxDYiub95LbD0xXLLYahc6zZbtEUBtdTzwX63M
pV3RqKwWRF21vNK7HAFIdIXEIsKR7n2L19GIDmPBTqVOt/G8rV8U3SLPRsEKesVj
zoKS3sEBg07TGhMNqMa6x/aj7nyAxKJEy8GuHPbT9ubhlTsTmlfXalTWbkacjlfZ
vgUW9xjC0qZxxrn0IINKKEWodLGG8c4D+zh5GrbYto4BlIos2FKCxPcYnKH4Zo6i
NUfc+7m4fvtEGZp+uYJsk3CYYasvqmMxIazTQK3g3irZM1zqWBpuW7im9HzbzUId
Y/aQGBrwuFPEBXEb0cnZ0HA3Do12uQv1PpdjITzJuoYzegSCF7jQ/Qc1dT8jSqkl
VUWbvZs31glncdEwPGjmJGIKwIpZYQzv7Ft8n2v0b2+EGD2GF6/lpgbNKYVklxzm
FIrB8Lslftx/bds9tqhQyhPdpR5IMEEpPS4QpVY4eR3iRNNEVLn7m47ef3U/i+/q
5Jh8++fev60JKvpgKo2bWVUbt9fmpcctNSMgXefcEk/5x7mTSKu7KezyzAF2dwMN
VeHt+W4B5leiQOTmnf4AZvPmxf/SH4AwXmVERI6tTJaiKRKmb9jJj4zXvX3chCRo
6cHyvZFoGrF6HXP6x4CNV/U3yhjfSSsb2pzQPpUXDUnd1+ZOS2CR6XWdIfeJE5Jr
i14c5jTYWGXORMPJkYu7xxQ681Cxe2J5Tb5CyWdrqzGmseS6uoUi4Ykx62aKfyHS
t/kHpTA5ta2pRmxtC9UMu6/O9hrRhxKd8c4METTWwHA/dCdMMEY/BjdtP5J2Ae4A
b1V3yjHXry+YrinUXwRPjX1ni82oEneJALoGMJ2VVFI3ItkWKgNKbtY2XPPXUshp
S5+YuzndWPKjZ0UR/rrVIqV4cDqIxNkFJDueYS+xFsZ30nCduwzgFMabmG7dZ8+X
eEhOizBXgO6b0FVGGpCLEd4NNtAl4n+EsbbtsLtOlM0CcMnXrvs7qKeoPSU6X7I4
u2mdz8crePfPPZq7OYH6X3Dm6AOHco9eLzQhQKZkkGhAIk5VgVKtn2Wu8o+gumAj
DFS2FaxiaOh9cMKStLP7IypBHuJGWhraTmC+Byv6SVbnhhbQYVLLpAWuvjDggq/o
AElxDYKSTcOMwzomvI21ZCdZn7Uin4N+5bZO34+hms3IVzxNuPUjkJzfN0yK4icB
3u1lYk2FW7YW2ljTW4QwJ5TT5DZXd2K5w5Xs6xSm8qum76n1u7jrFEno+EI2BeyP
HDdAChlI7B0KmfPrPKCTNyizP/6Ylk8u0xFMSztyYsDQUzo5xu3eIxXZGnkGmRWV
vYNtX9z9ytHFLvD2wG3i7oc4Q0XLVUSbhnSqiqgbbtH6CSVZqh2G4d0b0m+gm7Uw
4TSig6R8l+tYIoPEqEFYPy0UFVmG2KdPUh3UgatMmu6Mu4u6M3HHaiD0XAO4FYxr
l9WwvfnxNeatilxQJ5kpe9chSqjVd1c5LccfzDMkctWXnv7zE8HB+p94KAjoJ7aB
xALkfrcbBHplJEc7DsFWhup2LH1dhjAxbI8bq8FJRI2Xp9z/HkTKqyKLdBbWYox5
R24kkFWU5afBWc1TN1PZY6MU0T4ReeoUShwWXf0YvXLjaQt5+25zEZU72KWYKhEv
oTaN6SABcwOfh0buvtjQI1Zsji77wutrBOIU74rtRUmDunfLq8Y6oSjbRrd+pDLB
R9VoY8q70figpy7cRCDjcCTVUp5jj1XiWPvY4plkbdqxG3meq386wQQAa70tu0+e
kM7M2v2ZMrc9ok/rV9FQynYA/PTnL81jC6pEN5+jlmFEpRLl+r6+GkAAjbwhZt0V
bITWsj7C+hbzVro95a+jvofzgNNx7cN2rL54zAXEtlgOJWIdHr8JfCmEWNbNNpi4
P4KmIN74srxknXUNdXYrqiOwUrtlEoFMRkaXz4hJhh/9fIhHsmVDlysfeIW1ecIR
nyLPYMOOkuyv4bIjog1bRy+iKtS+WKA5zpall2CBkIYnRgF2rjN6gAhJASuGGPLF
sPvBjDpfYSYDz5VaDD93H3jKC2pZfr5bo254kD9xKRGc/lAJGdXvH1H9vSDFOO25
nw8an9aDDr15XtSJGvaE9qveIe8GhlpPMdc5B1cDRwCxAYS76hOEBJtsdH5cZ74Z
BFY6H4YHdZJz+V1yQU7c4hSlRbkdDMCeYXMNvQMyk7ewjsHpc3uH/FYnQhD9fTVY
TpMBikYvtKe0WNcuNxYCM5V7KsYCndOh7nhwwrb8LR4Z0a5q/si5rEInDS/h+l3u
2CFGvHUTKuxGUSFtB7++74m6ajiN22/7XlcD74y01eiO8Ny05myLfDKphIL8W/IQ
wo9HZ9voTG38rRotcMK8LV0Xww3OXxMknOlfszXV0wp7Td8kWgaBruRfMF8DuH5w
pcJDd/9GysSMZrwE+Fyi51w/hQjVt3XVXWLxf4PwjRUbitB3t72qrNRZPvDKodAw
n2YPD3UQHEVMJDZZojvhUvCtluzRQ5W5iy4ltZ5qpU0u9S6rjmemxENSJZMGYqlk
YStGoz0RnVuuNbEZ2ZlV4ZT7PdT4+TmQQNtSPS6P+V0dLoCYNk6XSJThSa5d9pdP
RRDi4fx01Wx/3XyI+M+HdDhil/0NLJXok3DetC/0tQ9uuEjs5+Fhr0ilDT/0tbCw
R4yFQkS1ppL5h0qoGbeblRP7NkiNbd7wqXe1wlx/a6oBs9gpwLGIVeWRIDj/alLJ
s2w67yJWvTtIcz3nyOwom2cOeQ4Jl6N1nvIIsyfqGT8Pmc8iKKotCuRQgVvuMkW1
LXMGaLMzg93dcLhPiVJMWDxccW3jbKRu4hW0L82EovQpZfidB1th46LD5o9P1Szt
Nk3o4fNJBGElsSXWNIl0FRpB4Mncsro81b3tGx6+SuvXR9QzOHDx63wgJ+4Noa+J
+4twqDp9wDDx1irjEjYaZA/XUn/w6WGj05IpavXeGVVQqYxf6TvlERc+aAsHDAOf
gFqJTF5WsG4zlVzD+mUg8wvVH+Uy/IVYoJjRX5mkdmoXU6ZoIo4xv/EeZzI9+fV3
LApCqkyNKnMu7kB/V34mdEkyo/mxvJ+TJ2nqS2Ddgjp77sBx88Reos4BCPG8b0wQ
ISuD4gCMoBpDNtk2Qf13W7B6K9qk4+92Xc05HyZYlEXBKjMMUwFIAOi3AGarOsn/
UgBBjVMCv0JSupAC7gGscpwo+SvZGkAsUMQ4LiEaZpFoZUtK+OiFmFtlT8VK6+9i
qfAbA13rKde1xmwlsQEbbecZ1GHQtGCx8pxlypzLHuYmPfoG4gbMP5f7x4b7g1BF
PIP8CFx85COh5z4Opf2yvwvMscrToXvUSZSYxP0Bzr0WBNJ0mnv4UfYV9L+Djyf4
IcPSSA2IJ6LBcwVgsnLQ55I3FWlcVd+oq3IhW6ge/DqmYx4kv6zdZ+qoi2YxZ1On
gU9XdmQc8deoDxwcPtUHHjIlKAf+Wp+wd3erygR0yrjQXdXPY07cuda2CzSscXsK
cA73lu4C8CtT2qW8GWADLyjwSsI6WXh/uLx7GhkolbapCApNnKwGQTLC3Lhuy51/
GEAQz7zvybFHYbW3hqOd35+pQMq9XvXlb5NgWUirRuZMszWlQM6C9QB1XDpsFH+D
t6+PkVq/WJteEbFgIqaBnDpz/LmS6KdO+I8ExAN3OLlfd3sSaN+Z2rgreiaDMzhI
8lDfnERrbXKlidqsFzRp/bAn7t2VQ95wAXMh0phlfu/KldAnaEck+yYuOZoneqX6
j97H0EeQNlVT6mQktkDV4kJR+BpP1Rypopxq/QevyS1+RpcOe+lOO/RMOyoIREA5
sFf/0q34tLFPpl+Nzu/OSgCwIgAfvQbL+JKan0rYY91qH/lDD50zlLCx/lKkCuh7
QnVJ6fzPWCegpiEfnB012uEgAtmwCHxUh6HY5kh2Tkjcweiht/H2WC3geRVWstHP
pYam8AGzWwsSYogOGEmAHuOxdXrIZgKUJxE8bMAKNWge12W0RhZWlNnc3hHpQoaK
K2f5FO1dxXodCYdPh5yVqeoC9ugTvaf/WP5X+SJwo3OU1JgiqChG83IpS7HFiBQm
2l+6/moxf8KL3XAw4MR2zvpfC1ipmEBGE1E3jhnVfsZVYtreyogg9hBpRrg6Yh8V
NlbEPNgNYjYsarD6RgYBknc4Yd5cH8Fl2Qe6p9WVcaLz+NQxhUzqNmnw4vx768FM
5RwlSLDUa7R+pQ6m+l21LsDFujHcvbpHnPn3sX5phaoCtyfC4wahdCAe2HefNEeH
3bj42FYtP1XZ9eOtXOBFQhKn1RZIHVgS0LIA0Xju76r3SE/HnIXfTEKEvWYXUqCT
04YjIg7tcNbTveY5Viiir7ZGB3KUiXOW6UGrRUCNbEY8u/vCVS2WU94uSQpw/ISP
2NlvA+rfTPvjkplIZDhHX3VX2zi2e/sBuv3w1Kz+rWMo95GPvnQDrAzQzN/GxIuB
ywTkuczni2d4ppAz8Uc7tw1xSQxsz9lL09CJ//lhN8VP7yODuKmEY+TjoGWvTfCW
3NGKfXHwm9dDRVc7imX93YPuGRnK+64msE0SepHXjcDGaDWvreQLSZ0KZLYVceHw
e1RlaOqaCMt5GJKDoFOCMv82+T4Ynh9OVdGydzgJW39DOZseA0NmkZ9PfAeJ3DaR
eSke1nx0/tChcDdPrPJgvPKMPIiWcBTnnqu14LbIIkw4rEPlYa5z0TnXNzUTBRr4
Ed3OmmwIq9dQ9Cxl/RLcBe385E4r6KS2cmQRqWv5GO2vLO5ev7vDwgByC2I+DQ5j
xQaSCd2gsU7aDXYCeoboBXm7ilWrWpoqUCLXmm9+FmNWgE0W5Sf67k4hHfdnia6G
ko2Q+uqowkqiBNbgQ9jzUnSAuJaNyVR4XP+m4HJaL3d/meCEf/wFLqXmAGkCizFj
cLNSExPO7AoO8uAF6C1Sjr/ffH/IPwkskCyGWNnSW3wmm1FnzzP4bgI819MhZbzB
Xsni7Co5rnqEcnXXmAiRAL1e/H4bKJFIzdKn8+LO9IMvq93OiAH1CCBVG1mOXaMF
4jjnQYwikMZX4nJvFfiNmdgemP0wqj+nR6XwwHFZW/QT79/7sWQcH+Sk0N6EYED6
nhVZIr5mftYKUPX2kEF7pVVGRZHc0On5kFvV0zDr5HaweUmtu2sw0KwBGQPcRSwA
SQRfHpmKlW5f5QQL4/08g+OnJDf8JYTQQGhym2pkgyA4COtbNR72utJVPbt2+vMY
3Md5Z1MQuxFfg/CzKvp3mSKtAsRAxgnfbVl0nR8r6PGZ4eIDTToCaycviIUVvGMs
cE1aE4P9Zj6yYNeplq0kIHM+N3dBzMReN9t2n9BXtwi1Nbu1Z26V2zJr/0meTcXh
mnnCyTBO/WFuIE3qUSjYjgbfcFz1sTpo9mksm0FRgQWMnI4Iq81rysnLuGaAcuXV
uRucSN566Ul3v9ZPyfAIpbPjhtHm3QoITauUrVzj2RYjIfI+mRhZi3Eq7eACXYFj
EZK1USeOgOyOyDpPKWxZ0TjwNUU5IeNBEtAOAl9TDB8pO7bwEBhU5z9gztGfLpPg
6EnFoqqH+zO2qMrNAZxp3P0corJLqG+a8CE3HaEF/2cd6R/bbfEoZbQT1lBa1iqN
DY1GV9IEY4UtihlN8pIgWnGUa6a9FLJjG9AIcK91FvFZfDYdYbTwCjM1rUCtqPVw
hahK2HlVtOO8g0rzK4GbmySfL0osiWI3u8A2sUh6ybpm8vTph0U6NzDQx0qEUDeI
Woi7iEiNcNDg2yMD69ziiTNo34d9cDxJjE1pdYtPVeT30vIWoqOzZpxKvJdTV0b8
pz7N0Pd8yjMsveCBKXVtX62JiKmueKzcatuJpFXOnTSsl+aGhxHoGHUFjYP/JLjZ
E3UqLoGe5OqHMu8qHOtPWuCdOPxvbCxytZz1sBpee3RlNqVu5IkMK+sk+VuOI3jp
smKIR4cV1Yu98yrY8lBWzN5V96Np0Gs8EtWLKB/StgQK6IYEyL9s3vsejQBkHK1g
8vOTEyuEoOH49enxpEuffmNCXDzPe4MXcZ+IkpPia+3CW/bc69RUIkKWJUy5hn4N
MNRSdD/GzmTgKO+jqglWl734w5A4NE9/Ho7ZkJp1cBjEHxb5IojCw+GfaG5My7lO
IP9e9ysUilyxmkY2N/N1Ks2YplIVTavFoROeZumMhZ1/VtnjaUYeZGNck1Knuk7t
f9A+wFNDKsrPEeeUjKl9Gt/WGhuNh/KBB1HoNSMFEK/YdUu6Od0h/n98TU35q4sM
7Y9bXBQ+XdBZRKPu9LdZgR1E9sORmX2Vj6zB4fzClngJek70tD36hb8pXzZ96clr
nml21R62fqAUA8Tom80liDHEgphN0IsfUN61vOQx5bQ8FwSX3kYMB3WUctijty+6
eDVVqfJadpOfn2acmadnIs4JXKOFHU5w2gDSPkbyshAJUrGwtBQNnxHyxMCum4f+
asLu2GLy//YhAdmfSC4G6tUOCNk3/n4JZpRacbUcASHPXk65QBOLpm3HZJQWy66y
uBb2tcl0d5BdH8+n4M8+zsAaeMLdYr1ZiKiLiQZJ4rr8owkp2VEUrrQq5aEkKeYN
dgY8IBeXT4EZl05XDor5AZyFzXyEc6hHBD0huIchNqh5IM6wjrMCgjjUsa4cPMPA
bVs19iCD07Ud/EKfoeSGhuyliTDTyd4r+aEDX7UaltJPm2UI6IzlLj+4Sr5f/u1h
RcDcAJDFwPYucrEQNYww2h/haSWdpSNxAtM5nO1+pfPkPDSMi9xcnPfwf3gTZ1xY
Fhm/alael1kjiIV841pRHnx1FrNIXcEA1b5HG6gyyMqEnXi77waGBNBr+73v+KNv
tBaCkOBZYq1Fv4O9KM/hIJUZs57NXLEtLi8LbEClMVb8eLaMqz5nAWOUHgGkozVK
HE0ikAaHb2LG0fPAYJiNfg6Ee8sjbCs5ujqt9RFZ6gJG8WvlUuDKCQw9wgavT05r
ITxk3f8KqbpKlVhP8Eq1HxHRuJ6SNXHmWOwbnkTJS+ueRoi7VC2Lq5XQK8aTIj6f
0EJpLk6nP4o3RPLF3PWm6odU3sJc+ZyjoPKbfPdDfDcFYqVTYnTgnNm9mOLNqH0a
BCx9pq/u/1Po51eaASwebW3a3EScWnRnLAU9peDsWuJm6I4HnHou5E4z5nYYsnK6
hAuoMQtjjaG7f2kZACTJM5UrbkokSJH6RbDyXzG2E+hrwxCxm/qc9nf+I/AXecre
q8/ifZ7fSe0OdMh3jk13zzKCxB8DMuKvB7rNpMvBza9TJUN7KTgHTsO0rfBgIzhC
7uKkiJLzMgA5EBv8pL9CYm171VmshgQ/9d+EIcT/7eNBPNr9UOCoiin+ftilICtX
aKmHBmUeXr4eMBvh5Wnufq3ny93eCyF9OBuXj2ZqZ3dfdMytNt/VfIWEsZnJJO9O
SOraE4rs8nttltTITxLh2mS8SmN1BQHlohh02cI96Be3cKRurDkAW2M+eq+/an9e
rJ1b6hzv1jJRTERyfI9MQUux8jKbbweW8WgJq99oV/P8r+SbFVKZnsWwS3+87Fu3
t9rNElGchMKrtZDYApXJeFEVmyxAxQOjLL+tv0AkhAKXtVuhPKDCU24YhsqayB2A
sVCnnwMTK2NMOqpTWQxQpee82910v6YE9JYXWHLWJuwI9U7rDbgfc8H6jvs2pkSg
1o0wEYR4iD1DozFsRiXKypSPHfB2uQbEd77jRAJ0mfUACMWrKP3WbKcFQa88yqeF
oCJ9jB58T+sfClpEFrvMiZ8SpOVWdfZJ1cHjYlyUwdFaqRFsgvRC/rs/zBiBH5du
GlJiq+bdVNBUgamcX3BsT4Ex101WOHPNZIYoOmneDzEkRP9/P1G4pxgYa4sXfP3H
QgFlIokOYN7oNc0Y7cJ/3L4kyaPrd1SuqytHnc1apwgy+4GkRRLxNS8Au5iUVO8L
us1MAO4MZ0q68Wc39oPm2kJHjF5vy2aXbwWVfu+kWbGX5ZodlzDy0JBX5x6XrDQd
X3c9oQ1OW5XWwl9qksh8FZ89xpmret9FGcyXc3kGVSmvdz1/knSDPsp/xJHNgTdR
r4my5MODF6rh+bjCPCaPisKqO5VGxn93PqCm9s326FWfOYg1VjqDeHb/05RIO99Z
SfL5R9an5SBALLEo4gu8Deo/wq+sGMb3MD8/uFIivL/BasobEPqTYgeCYlnzSI0a
WGIVD92QW3c75U+rPl19RP7SACCsVvNF0vf4+6fq5IdudQex6k9hL+Q1LKR0BxNG
FehrljoA66UT7v/dvta0q4TkTLm/m9rEQpQExcXDdgx6rncn0tQakKEsExI7IuNw
jsTCaSwQD5wURnpnZySkuGpzcRwAaDV1ZOS+3U0lhDFpPd1UAJWTycCDU9N+dKKl
BavSaECpMuHg76VzQOVGFJZnaLZ+kAe4rKeHSoAy/iKhm9Xi4UZWTNeNzLMve8Uv
NzxTi08sf6QYT5IeaPwo4hupNLmoN4B2qSMrbk+e7qQXZzQqgh9oQJmgAyfSB4db
y1qma755028w6iOVkecB5HXASeRGlt9CugmHXM90CA2i+9hAh208ES8ju4bzbiWZ
ZEtw9hu4XQ9t4H0mN7GIY21MhlAi10PQIG9KGL85ToJyN7WrIJjLpHXGsuN+tCQa
UmpAyiz4UTjF2j1ASHwDDWeXKBAk1Fe8cvozB0O87Mbf1bemlpO4nTkZLick62pQ
wdmxUPdyZBgkIkWloz1swDtUplWaSeyYHLJRLC+9L/Je4XWu15Gvv9nz0K9UIazW
pafqB7ZQ4JeaVg1vo242lGLORn7VPShUxQB1V7FmJaOVx8TiTgMG91FGThJWJu3O
TsX+pe/avw/7L140rKUxPMUB+LriJ5UhYaSU0gn4T++2iTIMr4nW7E++PHPTS//4
ZKEV10G7fiHg0b2kK1CNZITHVItwdcAycPhkh+2j6Rq4U8OqswUMH/eHRJhw5VK2
xwM7WB8QfXamK3P7uXhCZgDqxa94Rz/VVZ3m+//erAcM7Sk8+ca9PCM46cJTcOp2
uHi25HR223WyTgl6Ccd8NHTkH8w/f0RI0ImCFPX0LZRWeOOQw34LUaK4UTQiYrFf
n0TEjUE+aiSfrUlMkkreJNUjzEcWYPRfACW5fUN94Ht8i9W+VCHwZjoLqTnmViJL
3pyiS0IKQx2aJA2KjQYVyZid95qI3mINU7qJAQ+u63SKajZNFvNgkgwWJQy+bfAT
hjeNG23yfUCjzzPhbmd4c9+l1Rc2Cy4zWcmH3iSUeSQ9HFEy84fMlKEJ7Y2CdmDu
QAtNH3mpUDYvRFPwILRXH4xMIRRe90UsjYQpZ1FAibzWnviaFBjuIPPa1+w1CyWD
5ahSRJmRM2vXOSYCef1z6cvKdM9DK9jcb1Z5DKD9UbXGoLUHR83rGbR0ujIwF2Fh
8vR/ilqOtTtALWMQTRl2kWa4O9eOe1MT3V1EgAIruBMqWDL3XHTrkCr5AGAzFaZ4
EtYzlxbDNNc2C2H64dEE5mTj5vJcNqdcP8hehyDZC03bmK9aRQUhPAdiVjSHkjXP
NXKj57ZL9ZwoFUv8JLkGzTLzLPfvgMrOdbnGBs4u59iKmPEaIwBd169xDYnN+IZx
WtDp7aQJhQ7GDPfRzADa73NqcSHfM8SgC4S/tG7F42DypedZQNaQTPYBIM6F9vIJ
JDx15MrrQ1W9Y0IoYWCHhMCpwa0SzGbd0+3B3m2IzAGDs4i4asMNm2uGOKCxodJd
V+6gyKSW0IhWgRn6B3RPfSp3al+SwYnOzo3QAI3B+XrZ2kbu8pkkF/sXdh26I18X
kTEZlWvfsHH2KxHmTzy8qpYJhZigZ8DQ2PTlc1u0qz8u+Pi1W3U72tFMv9qE4kqO
YsM3++j0dV9jCyWRYX3fLh2e5HTNVwzQtRUCVdzHeDFpv87HTdGi0dv+AC2oeAlo
4liEs7ab6nwFz4QVDmiRbPUaz/urH0iGvVcDfcTsHyzVsqjOsBsDIN+eBvYE/BIO
ykWSYYW1ujxdc37sh/sSqjRGiJGZZo8jeKDj8hZ5qyfivxDFZgF/5zHOt2iwMrds
XzlzE0lTvKREqWJXblbV9v3lwBSSeZOpdUu6xJ1DdklrW/yRQ4++oknclaDMEEm2
kmvqejZctKOtf1w624qt/6ah+LmhRd3Olr818u6DnBAPaiDf8pTOlF6uyyeNk4hm
Dnca/NwCZ6PKLtYrGaKU3ftHyTzY5qZzkUMCbCgRGZJK0wFynRak4TU8q4YYKSDe
DhWcmFuEPt1WsRpQX4zP6jKx28wjdZcECN92K812Lu9w9r4Bvg5A3kDh6aop2w1B
xm40ZzEmqgP7U6AUivrRK8idl17Aq662qPCWy662u736JDN/cd8agWqS1yMRpwN1
tvazxvdw1fTLNfTo4ToePqeKZL7eK6SHw5kZfalVqcIfH27I0uBeQDY1cDfHceUK
0D8P8t5v5dWcJEYLBhEgLyypkA3FwQbovsF75tHw++06YSeJz+Wa1p4kkIuLgOF1
Eean2/WeQuFLZS0gGyFQKR3aBIpHJs8jEdqhYrk6Lp//goa5bqjkNsLqpXSqQahF
r2xXdxIbRbkEhUUYRtlg3SKWhyoA35l9BeQoE74QxZa4jxUascPLBj5QD/8gK9wD
arvUDm/bBGsVCDb4FCLFbvA9aagM2BmCwGQjtcoRvOAMWCm3WAPJr2BZxUgb696R
9FqCvw7ZX+6TRFhlHbUyrnUP9mLIJLPtmCE/oPchzKem/xl3TxIdF7E1s+J52dRD
klV152uxkC5jsC9FqLX4lQFYAYgVp7OM9uYhoZz80MlilguBuFV3ZX5HAJB5rGzd
kLYUywRSc6r9GMfLGQbYoWEayqwqk1eHEnIYAinDhwW+drxjUJQU+f9HaleC5kwV
oQFoXIpYjZNlwFLVtBfiUsAy9YHaQiLSDLEvztjeuX7NBLexn4F2oY42Mfn6xr7d
HbvH87vyptssRv3jtWizsNTEcs4WwGbeEdE2jvbNmnkMJ97td1GHOkkRoLCYZL2F
bz8IquvuG4TwlqNDGXEVMH2vF6BHTM3yQgPfw84yYAW4XVKpZqKB8qHCGJWDM8i3
j6Rnrz39hQxvGbsEBASUfLOFSJ3qYYsfoRPBLHpvurjR72M3TkDOee3ZYtwHaZfn
JXeJhuMQETJGaXv1fFK30EBothlL9gNdHyKtp6PN6ybh9MptCaQNq7c82cPk0ImD
9tMsZlYBIlPEJerGkOdkyWH3hw1GSGZIdTsIGNIhFEdLHR6FL/tOFuloXDooROeR
9dfd+Zq9T59sAlC7X1ud1Y+T1U6OL7iDBMvfU6RKgJ7hPRnDiP+oF29v8chOYL4j
x0gHNisfqLTeaDXOdAT326mEn1NsrRAQwTefZh2PflRv2BDB5a+Ge17BFMGc1JHI
1QXrCioY34vbw30ekr3EkteaBgUkRblEw4KxgDI1jMqxzY1UP4FTCmGXd4+zFk7U
2IXNWVJA208h7TMOnAQPCPK/7XD3oKOAl9Mm6IfN+YW21uVL6TbIygPrW/h/RjbD
fTO6Kd/vOz1yCro/U4N12b8EkOMOleDNEIvpn/cjD+CVtfOnXjeEJ11z7qBUYUS6
nrzKUgzrOWJa7J8T8ix050/Y6EP2yBOMXk7gQr2HudEPhLwc6NdCmLsDo+gm32kp
MZL4QdWgO6/wk8FNmySYytq4W38apkVTvDcQIztmy53/XddjnJZ2K2Jnc0WgPxaY
CldzUc/KS35NYiGaYmbKP7bS5iU+uRqzJAbFBRspOUEr02JLXPWx/xyR4YqsRfVY
T/+FFmdpf2E6X49HCqPnj5RwAIdOixHX3ZMzvVGOLQueb/79AOYOOdHnxPfg1PiV
6ohxoZxC9Gjh1Mbui/+xMzGG8f2ihNGHV/iRG7ESPgVrIIzQEVRaOy998sOxu4Y6
xd8gk2By5Ce8owapW/J6hB8XaXrYoPsnpCZ2kdefqhVgWEWpFJSwqC/0t6npwYA2
vGsB+tL53S5h4ke+0S1IU8Alydta544ksbww2bUFnbRnBpLZqXRDIiyuNy7PpPzZ
sSBQ2UWkanC6pNHAL6s+HIhtH/mUORAwwjOXPoZqw8DS8vQ2tza8lbP5mLEAV7yE
W/9Kj2h+J6gQF3bU6eL87y767HOCTuQq+Y30akG7ThyJRGgx11mr2N/DPy02Zspw
eooKMjMDwqd/xqDII1xw0xEKcANaVnMEFZK4/L9BLPM1dHZWzFQ/1yldqhY3Qo/T
`pragma protect end_protected
