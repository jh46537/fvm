// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:41 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dEwZ7ZfnrfzxPgdfEou60pt5dkwk4k/1AJHa6RL+rzb8QuPoUP4muq33aNTShFDm
pw8P+Ma5iagK7sFLZ6z0tnqmesslzOUHL/OPM5omdORTF0GMKDCxmD2O8CHT8Hsi
22rtfXKZBBzTHipAUbiYp09fyMtf5BN8VEEOkE3U5OI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8448)
8WqpUKHFWN6w7TEJc24lugbXdKwjU7X55nSpC1fti8srK5g33OWm0wHiPp8ysvY1
v8LnT6pjxjxxIkqHY7EEEs5XofrDuwezMF+EOIa4jU7uggipC4vE9c0GhM/qw8mV
R17s0bX0pYccGkdpNRB5VuenrudoRHSgNuXvdGL9S56stliMvKx7xCeq4+NFN82W
1fp6S+vEFCUavPnADJa73Pvo4SAOYi8rmYl9+b1vnRyJfRChscbg8FlLxqMGWRXq
hX2lKh4yO5FMQ+GK5jZSbI+3qfHPysnMaX64C5rDL/m40Q7ksBusNAlJK9FKiHIq
59uSvxWMxIXloxJHOe1BuY7mshzx4GhJHhrDqyhlgiCg9Zr4sxD+HZYsRUEHMU9N
AbuHVIuD258Lqq0JXa817QnOl4DrO0wKtlhcTqHlqMZyBCCI2h1fh3B019aE3NtV
kluAb/TKSQOwjaLco+AoREYHc92MJyNrYqrJqHByHkN06ZUir7v1fcgcQGersmjK
OY/HcOhnoX3lLrsYHzwSIHlot/IxLlxoQCZ2EtTs2hJvaW6tq9a/AabT1Vc6K8L4
Ka7G6ORyRTTQ6En1JN7IidlvGj4xB/P411T0aw4gNiLCFrO2dm84/bripYa3Gt5l
SGuJXuK7d3TDNHl1MQHCarmzTSYNxuxC1tTFbW7tbLBnLz0o6awi5afyZluRUia9
B4CeoDWy+417zdvbvZV5ou281bH1Nw1qs8o8R/+1hCT28s/bYs6zAOsHC3t7aiWE
c4a1nnpXw85EDiprlgybRnNjelPmyEi08Ob9y3XXd7Mg7pudmymI3oSzgR4NSozx
IHBp6HM4ArSi8dWaqkbMnS5+F3NkmZT3Z6gf0pS7ISO9SKET8KCRKvC8aBHS5k+c
8yz7QkOhvhdAKr86I3HrShjx3yk4+s9h/Mu+iHsvBTxYvhLB1eIPYe061atBcgbg
YCzKbw6TAmsNcIh4v3qfYYNEvZNJtnRzqflyQYBAfIPJZCWzPAKQyXUsGVrDhx38
0M54cORofi+hT7u+x74ofYnJB0uAA5q65/+M9COf36hYcGpuEKOejy4dqr5+HyZi
xy1ILJvzrC5Z2gaKcraWYsFXSKVcESSxn5cvXI42xnuM1VgLzy1n5tRCQ1RXI3zs
mP0u1h44S62RR4+fstR+bXWC8hk918/mN6IqwmvjyFFTQ6DwJcvQYdX3AspOBxms
kseediDAA0F9H/R2b3xOCVS+31/eFO6bCbH6Uf9HcYPNh/wScDt4O7E5p1dPjWeD
KGJW5SOFzfgwLvA9UhUvfabP/F3JmCj+dLOGxerD4bG22gqIOC/hWeyoWj+Teaaa
xyw+wy+Ia2pH6EitN2TwImdKTvH7utbnYvYZovuVXgpNtwTEoXsAnkw3K3YvteAQ
gdnLqZcF3srwwUMWGy70udXpMS7TCQ8qrQRv3u4q7csBe+kUmIVrXfYqh9xwB+8y
bSsEz2LkJXtg/EF8q0VFFSAlGesP6Y+ZRIU5VJVwzCGLVK9G4sT0Z1jZSDcTBZjQ
kHnzlDizO8EPD2WJJNY3Xa1Te6C+SLKPBptZTarEn9eL+DhaCgndiM2SFIcwOzMc
74zr8dOgMMJT/C/D3PPFHGeYvVPjmFBf5u8NC/F98NXSh5CbvteauX1AMw+dcI/c
4YLCh/ymU300xjGFpqBjWK1EGNHsh1E1Yiy1xmnVs+GsVobUbpTYfcQL2MAH3Eh9
AmhiIazPn25bQgZSvajH1b7kfHLHdQfO232QZzMhLQHwNDsQuvBbLdNRMP0NZTwN
68/mYcqfzvx2RXAdcvLQ2qDEwRriWJUVbFZDuTKcEfRR80PtVLGBEjd+MWzYvS6e
MjQmdDJsn4ur0aH4/xbKM7cqFWXjDIMMxukv/vzfJ7g/StmlNzHyF2YIiLpGS5g8
CjgGhfP/IyFIi7N0i1j+6rPJpMIkpmjdR2/Z0FEGdmTTOUFfvnav6TiCmshHlS4T
yWvJXJvU0Ja88hDLFB5hWMdckzYYCR/oIpA2pl5nFiYVC/kPMtnpCk365KPvV/ys
bbiNrxsFHSFaL3GE29ELb7caC7YlVyMAk/f5tWIqOtyRhJD2tO41Sn7yKONdf9nt
gdoy2y0Yp1hIPEok6hI+9u2JoyHkKEpEivInLgXWvKgbbF3wbGtQCb/EuwXNd4FL
St1K/THlza9i6B1GCCdjoga2kTi20EzbmPLxxqNWFtMmN9p2PlG5+00TSHM9BhLC
joJfi87nfsaJ0jAo+SZlkN52LD76HWfhzE0WbuBifw7JGux0M06lp9IF7Lg9Fdaz
H1xwNeo+ho3q5vt35tKhhm/preOlsbAsFMcOjTBA4GR+zOlKlKzdIcofxX+kfetz
JHb1z/qvvUG1YXCQn9qVEkFNgSldHvJwl0UcFU35k4FTrNKIx70rrwSv5Md9vaUi
F0fV/4zpt0EYRxDzr/0UDQOkHQwfy484h361jLqd07iG2NvOJUxSD9IoZzB7Jwu3
Z5Rqxf/QphJFEzq/eblcxOynMc6wwdUmUoyMefujubc23+b/638oFkWqgaU4npbQ
LkQkT8FOxosJU+298Ysl0SYMEvbfzMD9/DopKnGh3YhYb1wLqnN3M0XWEFb35Nvg
AC/o+M4Qg7EihqwcPJPG4clNSRQgsUGjXFEnokZA2vNEuA+ZbG/uIdqK2N/nTlUl
cGbitDCIRjxvI4ItrjpSPl5zz9cisVVUFk1SoyiiEUwjM7eDoBF5AA4DHL03jAsx
FsXiNxAFbAZgemleKeyIE0SZoLqaox5j09oDJNxsv8mW3N98hLOiR1cFgWuQhiyV
ItzPLuShnmPblQ5RpBzDgvSFezFy548Wl0i/kdHxhHU2MUVkVNV81rUvzSLTUPAk
wP3PC9+C1Ml3J3IQSrDGz8ThCugA/yitxNOGL473Plc52+j7QlYymPsQgzPBnUzL
qjPDQ/7NsaTo9l/H7zxByfObZrFBLjLbO3Yj2xUy99WuvqphBVdXX/oaCtUG7k9E
L1XhTEG7hSPetcV44q98PSVU5jCsd6Pd08WhxNYDhfkMqdSO9mqyX++DmiFdZHyI
xDj660JzaNnGviVMNpScNPAgpCPZ/YS2SYZAkXOo0ZjLmGGzlSkdZQaUtadQG4hK
CToeiCc8yYDQsVH9JsYL/xzOQ4oUkXCP6wt2X+FxlziOAt6CsdJlfpEwCNaHXfXr
Ma8NSSJ6NXefw4X6mPkEymfPld05FEdcmcbRVDTVMCHLVX25eCX3gW21YRH7QtqF
7maTEk8xUZoiJRMpRonXyTnYvbk9hibfp2aWMdwXm3AjAz/zgcSALm6rVjArqeL7
fBqMe2peLkqk33B+EXAj8sCDEaEH9O6McifqkhigI5AMZ0jFUKgrKZ1deW1G9ynp
u2l0ismn/WMcSOj2Scl1k3IMdeUwyDHum8KwtpM5N/B+v63Rg3IarVD29laN6srd
uycPoPdhWsY2B2JizjkMcLXvHnxm1xAFuDwWUKp1EIfeoQVCtELkTTSULMXv3GYW
V6crV6J9QFL2jElmlXP5yohnQxGkI6anX+o33Qx039SXYxjM0x3yx3Ahbin0Ca9q
yZ9WVOrBKGFHD5L5WsPWltC+nAGACz4ozXfYge//7x5M3ltUDf4OjoPoy6MuXhCc
JPxv9gACCVncQ2UNSbBOCOwfSVPOMM3FTPPjYIjcNwqw55PNrxkP9M5B8eu1DNLc
tbTTAcBXmAIQi9TNY77GD/VvQWMpa/P0iKXDujGONdq3RculhK+OItzbRBysdkA1
x6KouF/1eYWO2zo5yIEc11iRZgxZdGb3PYmtl47bPlfb2CWaq6Bfv4+u1GZqYwMP
Jolx7gfrhD3U9v5kPqCIxOUg6/br3Ouqd9v0PjepyDOXLBjC1zaU24Fc04KlcPjf
lpaq+Xl+m3HNFj9JErtJIR/H6gyl8ivw5dlfFQbCfc+S0ySC5FrPTmntxWKaSgLY
4l9QncU/EyYeC6S0SB3V5Sh4QceAHxGncmzgFYfzu6h7m9q1TWDke7SqjzUR3I5Z
fhjHtMpsi5BoDcWvG5fSgcVGIXnTimC3zNbRvJSCyZCbFMjzsJFK8Am2U44MO6MG
1QmpG6ino72Q+Wk4epTupEyvG2CbNI1nDyxV0/UQ+xmExY4rYsUZ0caSz0HKevWm
Ra+eyL7DxUc0rkwfxnNLpLiJIAdoHNFpl4lD0XMTFGTW07OMkCezmYh7KaUZiqux
eu+bFZnQtEjGxCEjCZu6oH3xJH5+kOQwrL7h4MT96fRtQSxOpw7yMtkO6KnLkPlx
/EsqLGIxZyYGC3yLziTA1KSsECdVD9KYYGRO/3tvsaY38chfpqsS+vlBDS2Awdq+
vcDXNwCS9j4CJpI18wXDd74qLYAgYEQwmuPFIwSjRjjoAxhC2zsyAsnU1dM56T9N
p3d9eUVD2n2sYoGb8/IkS1jArgRR0BCOwomV5YBb5LNOZ3Fqj1oEQcczLE1Q4NUP
YNqWB0l41OTvRuoAx4jAHuLBeoj7GDca2/fzlgAvZ1ALUMsVTlbNtN8TvMDD7Enf
PFKv8x0Q4R9RqgsmZGmgC8MFBx2TYj2I/9EVWMvgCUaZd3yyZ/qvAS8X3WAFLutj
fZj649hSiNexw6AiR3eFOe1ilvn2abbmJ8as6+vO5gjfVPdWzxgApZ7nbB5isJvx
nAvMLHosy8H/Okr+tuI3+E409sjVQGV78l0glk1Yfu1K9TMsqNfnha8AHgrWVqCm
klEkP92cBp+3RaCJGalqMwH6MnFw/VVUxQ1r/PXvLiq0UPxNPe79hdqmGi92fPnS
Nb2W6tfnpD+gLRcPiGBuHv2IMA9s7F6baKF7HnxWBebf4PTy5VN/YtMavBpTFrDL
Am9UAkUntxCd2SjYk7+QoA/wk5Ev8MUGxW48A4nyyKC9hEwPNwqCsNYubbmR2VgW
EUycF7IYfW/8DOw/3LOAdb5qD2+UV7sOkAlaGtNmMe5pF/99L2rpO5BlFTTY7Khi
382sXpY71PHc15iMLMuxzN/kBp0Xi7pzWv3r89JLW0AhzHfUAoNL3p6TS66oBBWC
dwDCy+hIOoQtVBMGefWff6mizyNkCNu+ggG/P3CzBytDcFi6xRlOpFUVweqdPUvY
M9HuKDVnbl1q1MLg31M8NMb9Q/HklyWXao8iS20Kntp2lpcH/7K0GhBiRdz8Evb4
wAVE7HcOZL5K7yU7kmkm+HKk7kGNkDjsJt///jAHpCMfoQbP2EU8BKFo1dHSXxKu
udrLM6UiUZCiIVHjvHFeq7wpv4QLLj1yoojsuXfozmkBP65NAwkVb1jfSEimynNc
tqUVrK5uAy2sVCg7UpBsYeTGEC5DUFIEMBxmjQWhiPrrK9rwKkGUQno8OUcuXHYI
uoG4b/64cNMX3VuVLiLUovknePwOANw6ZaREqsKTCMYpnrEhLjwBkYqOVWD4zssc
bhbSg46bhBMrkCrZq+YV/274VtTE2Vze+EVuZgcs1m4+oVbVybMWSt/bAxcfOPQA
Fykgt85/nQanqty8JkksSlwgHfkojaDz3/x/6nMAlZSVG4EvKyTw4FHZ8Zut3Pzx
9LQf/nAHWIiVFxdGyetrEdkdTQXwCrJi1n9gJ6Gqtyfrn2JRZCCOey0v2NKRCvBs
WJZpbjy/P9ROiYfqngvDdNwTB/IEYFix002XHzpaB5cq8w+HkjxfCZiS8rp6iHZ8
rxhO5SpsxK0tkwmaMQhR2IKRYA6fSYvFmRFV1fQG579E9AHdIAx8eGMMBpUxolfb
HxgJtMbudwuoeC5TxnJV8ywBg+ZC32NFeuQYZzHsSR2G2zv73o1Q2RazyZM1o4TY
KejbgMpCjivNs6cc9PcMjdweGYzVkv//iFO5lMSX+8wXmY2sTCMP/5W3wax09i9B
quZnfhWLfxggVHYFiYRhPhGbwEPYnAoW7bmvaxdEEriH/Qlt+W1NU5ZxjWWM43Eh
d560pstxpme45SBkuAnI3rOCdBRn4xEbh/TfchiiqRPz7UgV3IjZwJmTZc5Cwdf6
UDr9KIPbreT7Al4dfbXdpzT7MtPqOlgZIP2B+Txa6a7uDNWN0uY38IvH9JjXbdKz
pQ8gZheJyICVKam+KOhV2aZ2GnKK0utvfIHO/XeguQyXhgw944wops35EP1C1M0g
ZvCZeebqxApU6Um7N3y8hG188XsWTfslB1a0zvODA6LtsIPeg7Re7JmHzLkKDWsQ
NsINHqkIC5PNfk4UhwRrXOSNGgSE2to27b3m/rQSHMzAW38t453X1Qa3EVQkHqdB
2zYDlJGmwD6ZeVFGIG9Rs3BoBDKbjSOb3ARy9jeF37sOV5q//NHfflhj9d0sfgHG
LMkYCRdOx710+PBuYFe2mzvfo3z92Zrqj9xsh4q3ix7PgI0OfvPU6qAeMh8wdJuO
idMeyxxTpCpNlCX/Rd44f9FV44gpS3oBheEJUwBFHoAXXbTDPpy3/1O9fCgr5+ja
DBR8rYvmoB3Eja6wUKTv73otBY4eCIgWps+31imOF14cxycxrzAZdEZzfnvC6gZ7
ZDgJ7oqCAo29tuPgTOlQnubFSZKZBt9wKHGKGKnYka9JuCiFwX+96ZQnm0ILcNyo
t96gnd4YyKrhmHfnIwhCb7/jwCRDoeZwXQpaiz/sJCvdZ8wDYM1YhTIld6JhnWYt
ZRXtzoiW3Nu2BCdLujgLeCokvO4dSyg+CSvnwaGZ7o30RipvuQJSy42wmt+618E2
PrluHUEepSwoc8vBF37ZfO0uMql0tbMedYABauc8Qk/y/PYJj+a5R237ZXe27jyL
k4MXij6GL/0GkCCLRAj1veWoSsQGhSJcs4l3YJDniqQOJ/YAlCRMXNTb3XmxExJS
wjai9yNzc4n3paP4G5bF9CjeuqIGmjUYT7w4yVvBS8w+FcUTrUQV4B8X/7skuDvw
WxYT/Cl9XzCaVIuetCKKcuyCWVCGUVD0zm3yMrubwt9NgHE7sIJhzrKJtXhpbEo6
7r1/GM+LSTWW8USn7KaR9F8hbIzP99wxq/CsbpjY9U4KYB1tVzaFstsY+g3fMhEt
5w8Jp9tFMIxiHQ6QHaCOIBG08kwoRp/L5bqds8hbkoQD1u4EzzPBjzrn9RXWG2CA
89s+vkciiNeT1JQSHeUH3FjtlTr6lVD6+/jCwC5sxY7kSnuoYP6bYm0u0WkMU5vI
Fx6j30/hgpWyusqAh55HNvqFt/qTUcvVKzpuewAz5Ngm4P1jvYgzQrQ1VcrqH2cA
lRSx5rqPw5yZxPxlSuVk15/O3J/3lrvqxbvqXryY9seQ2XqUi2NySqI1PxwVla+n
Bb/1fEcwY/iBdRUijg9WbreV6sk789lzGs039L2iD2svmpXMw3kOiPRwEtVzYEh2
pr3lkEIDIuVLCTWn2GeVfc9wu5FjpOtTEeFR7OioLBH6kzvKxZk7ID52ce9Zi6uO
Fe7dIIeMRxCJAb+0//a+pxsnvMBsyBMMUB5xkAuIvRwpq8sviv4YqE8m3NbRWnVm
WpWucmKIM4yJHGnzW80++ZdBYiU5XrrY6ZPupkdoHhUiWf/GmhPO6xgEHMs/plAs
xo2qkZBhKnx0hM+gMzsiEKSBANb3SxNSAvr66XoWaj2JDxlF81BzdIJ7qQ7IZw+A
x4u+ITjJ5pTSxsfrdxUAenuAA2STQQFSTHyfKdBk00PqL14Ja0Sin5eqLk/6lYeY
QdDBfchqBHVkIW58ai9yt7FSqLXhsGIbmE2Eswm9pGXw2r7e620K38qz5Ga/MaNq
uE4oMj5LfQ7uSp3ol5wbVTrhbREYoq5YmY+eJYOiAdU9vz4pv7SRhl8ohvJXRKMW
ss+zRnEMHtA2Moe4hlaTzLBMeAnCPKxp/cdZPeIod7K02w/d7ihv1xCEK6+pChUh
xtVWlyGjJpDE1Zjq/LetRbcL1C5xQDY7Lk8e/CXug7yX70/XeufbGGC0heW3tNmx
+VQ0cnEbxTVQirgv9PgQ/NFFIyj7/jvAIKjLCqvPwLVzPRGk45wE3+v1+6Srjf/a
qPlTbTtEh+d+xvbdPsEmCOD1DBSn5DnroCuO3ZCej2KCg0EJlHyDsfpUTdsDJRo2
YuM5gQAh5oJOZ83Y2WzwI3opiFgrCaLGsm8j7yyFLgbHuv23LPKCDPi4CVLcPHph
fCaMhCKq6OLyevzN4CKhWxocTygsdX64x+fZFzuTJYTogefLlncheqq7Krq3Sfkn
GKwR/GEUEpioluzA60co3Mf2J2FR/q0feiu2QfSIG3C34wLZm9KqJr/L2rn7optw
2Zm6zxpFfhTnQSfWaFO9rEUyCO/kyN2672G/MZxbj6r+LGb1YCc+qbdtwScHXbSL
TPdwaHN2lyObYxrEw5j3Aenc7VXtdNyAbwm8gPmmjAVvF2GVcHT5s8gfcgs2vAwM
Tvc4NT8nNXGd87f1wo+WLyG9M/pNovfRIcoQu16PKKgCOOq4mWFNuSVEkXngyx0/
9xa/afTX2tnuTdh/wZE3fT6L8NLXkR83R25/PPQ6PYoe1Lvax+S7B5HHRc5RrDUR
WcPloL7iB6KiRIvEPm0wwa/2TjLilv6AWaRAZ1z2i7ULrO5FhQ9KoJC9bmWCqh/p
j4cj7P3Vu5ucM2LbcSdulD01fbhQg88UPACMBRJ8Xsilbt083bzWJdJ8EoVWNlN6
/Uxyg2uYBJ9SNcnk1qavg9o2Ng163+0/TRTTmD9cGdsdP++L8fJb61hdd88kn3mv
09Ok1PKkB9DNFIK3sv44uPwOHxK7oE0+PWgK0TJPUO5oVBK5ZslL7I6ZqwMLIlzw
mSTIBwMhI5WqFFWTG88pp0hZwMgDpRUWRZdLn37YvOVP5QmNC8qWztx43F+BcWvw
rxbHnMg7z5RIUjROgnuu7kE55Q5kh1A1cR3kETFLCnFRMVfRoC5F1KHKulxUdSYl
WNtkjrP9qDpzB++3TsJXYNEseCblsdd90MpIL7+zqlpM0UOuk0uh4HW8e8AEuZKI
o4nhgSW2BkLddYBjvurvIRZjkmuXsgzE14uU5vWgT0saEFBnIobyWjzUjN91nVdV
fQnA8/PLLz+qd50gfe46gv8NzX2yzl0iKQ9LeWScqFsjnKRSadpipKD0u3dk6v6/
PcpMcavZFYAPQs/hpDygbuBKqi3v67V0iZS1X6LkyWZTjTDL2n18R5GFa3DdpwJc
HljK1k6Xy+4kLSVHhZ+u/tVY3Ma0qTaWvpUATSDSUttMnlh0S/A/vESVCIBEB9FA
hDF5+cLc9swWj/BbbyELiyw3Asn5Z2QEAysnPykpyzhUOHEhRFlhvl1RdkJSsRPd
MbYUJ4wONUea9HyXpVg/L3OBMONDfJKCJ9z5eRORgNNFrFjjltkkeErAiEx0T2Lg
HeCSKyjrxWJtNpQrhgvXQeq2UgXbT2qLVYXqqg9NAN+MGJYVQdHOF5YejVydtA8u
3YsY4nC7RKNaX5jqEVyGLKE5soDLqiXgJyaQ/8xpc2y4TMLKxqn4gvC5N9GiSvU7
C4/shM61CaOHUFQlMNmiywGkIA76nobEFfmQYEFNOaA1SQ/Ke1cYjbpHpUTf9al4
gTvKJlLKrSV909dylC7oBh014dJjjiNPkhSozIP6Jojs/a8Y+/MmIP9T0b2IDw3Y
EQnT1bgbYGELnSPnRbHi//Gme7dTcw1NRfEsQhuyt7nrV8vHuhUti7oaDc3yE9sm
sz76KP5VBcaK24kg+h5vKUqFOUapeb/0PvNN/PJjBJ9SwXoeRNpH6nhGXhG6FFHN
jVx76hrG6ZKvhsjWG0OFcSl0BbXZOU7wuacgvZjv/HGoGkFI+lesf/0D1qCDa38e
zac/61awii5c22U0mNQb22kN912pvxNLAMuOfP009bD4HmpesEPkaIhkOPufBTpl
Uh5j4+SQoV6lSxK0zbcXtwFU4VYWrFjkubijZRtlWMkDrvJdwE0XTB2CZ+Drv6DU
+p1nq8JlEEbfHzsA4rC0HsCT0Qy6os1JuXiJHIQbKcu/lXleCHfy2ilQJwwUi7Tx
DL83MJZFq67BKUkP97CrtNKEbaHr5VMQvlQh3HPaJnx+wwpDOHTX2B7lD7quCIdg
N7nUg8twchYsYG7NayOO4264W8kXbAyw1oq8EPa+fuKN/q58wz+ljZMDUDznATJR
3ShcpOJwSJmqIrQa5AW9AoTSq7Wv8/yDPO1pW/pkAW2uKdzlpKxD57EOq1GtVCRR
yXFECuoupIK1gTWviXuZ/n572V3ZvQC620Oe9nuFU+MneZaN9sat+CfHIOM4yey6
KyOzSVYEbPclwARNL1g+Cu05kdXodh95VQGFGT4r8zORHnSLL8e/M6cw+BIVX2xY
6Hn+SeO10soEuh5+QkEO/sc+MLlRUiKDbUH9jNGbTTiBFcGF5HeAgP/Eiwv7Muxc
+kfkqiPkRNmmaGgHpw2ihlusPwze7hbcAvqckAHg/3w0uGyKdYbM9fVS1+0YbMH5
G/50q86dCppNT1FFiR+BM/a6FE/83+Mt7lFRuk67rqLb2sERDEpXSV69Ka/1h/U0
i6uFG02cKr50dQwG7rk6LIjQnGoTb73+PuC5y/UQUpUl3uu/asPY34jXR679Sbz+
Pzt2iyiThTwPDEJsXeth41cEEysWtKH+ggqskUw7c13L6RWdael65hzqgZq90hOw
YrRKcrIeOgR5S8VJ33nYGlM1YVE6p/lhRl/i3PxYrQqjohq4Y1POh6jPe2TGOzw3
NVz+vFk1nebNE/dMkJwrBaoF9B8sMio2uu7Y+grwX+3TJCKlTRRikTr3R3BRqMBj
zE3ZvPp+2PtPvTTSWb+S3DIuKSbgnjM8d43u3U3s1Aq+Prfy6ELd2X9oiHVAtrNk
Iq3qRGbSt8tlt3qy/V967vm8QB6+sx+8hh2Bl7PtLUCzZSOup930U2vcTHaTyZA7
APCiNCUpICqkJKNb3uAPCGIUB6JmdYDhhg3opRSzlZ/9herJj7aNm4Pn/U7xBirp
Hxv8QMdCn64OujnjzJzo40mabc3ucpfgRNUZwkl+/qzLCO2ohOkLEGGOle9dTXuH
9v6xiNmqy8ElcsZ5gbyxJ0EN2ZlseQqbgI6Prvs4ByvOz6zR6DUrbXCesUwg5ZDF
cc0LhP9hpYlecne+V0lKm/WqlEH+UCl2Hyf8gay4rcOAXVaDBsZHnJHWqFXzJBlz
oTEV0GA7WJsGsmAbO7G128fyVDtqacyLx3JyR4ofRgO9I79A5n6kXQGGNeI5zBPV
J+AZWwDXPuGHMNjtUeRunZoakABf7TPQvzaM0uf/cc0jvzN62r+7X6SYLAJWh838
`pragma protect end_protected
