��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B�6ƨ��J�'��GZU��l+ �p��Da�H�7�&�9ޡ�,ۖ9�Dh�g����Ɩ�����h?�rq�AΥ�(�����1��{���$�ջk�
u%�K��:���O��e��n�����t&a((t��26}rEN��Y�G�՜���Ȍ9��7J�y�;�	���'[f�e����L{vA�zPiO"pS��Z�T3��My�`=tE mQ�u�YnH�F�T�)k�^��Ol]�q�Tt-(X���\�xtܒ�vZ���]�G1���Jzc�]�k���N�n	O)�����t�x�;&�f�6'P\����^�.�P�^i��dsC���R1���=�f��h!��Y�%C�bK:�vQ�9�l*c�E�`�_�|PB��L�������e;���٫����>느��/�p	8�o��_�o��&3��;�6=+��|m-0#&���t0�c��@F��I/s��K���3�����V��}@bdQ9^F��Tu}�C��R�#5���K0ٰ��ԇ$p�0`x����Ay�3���ђ��aiE#[����I�0�����D���`���]�	Gf$l;)`�+��؇��L������Նh��dp��"�N1�`m��X���y����{v70���ΐ��i�gz��p�};_�}��(P�D�� gؐ}��U�˭� ��4��;��i�
Ҡ.��۫��=`�a�	M�GT��)���j�kM�N+�ME�r�՘I�|	���!��4|K-��+��t
����$R�23q�SC׻��7H�)-��½�&ؐ���sJp`�N��5�AFd$�K�F5g��G�P�]���M�|�C�A��`(���
c����0g)�6U=;-q�Ԏ������F��_]�`�j�֮��BY6� �>u�׆z�,��z,�X>�4�3�	f���(y�ts��c�q|�5��_T���:�z<��}C���"nق)���j9��]�6��(!�;����\>��eR��a|b#zh݇]�b��H,��)\?�bD֭O'$zV]�> 2I�{/�qkJ�,.�)_�.�����9!2��ˬߊ1�:�Meл�kq�݂��53v���7"�%z�M�#��'����g��^�g���,�B�}��AɆ}��eց�b��@6s_�{�{�n�G���W�1�X�]���cGH�Q($�[�_^K�	�k��w�����|7���V�
F.E�ΰK���7�/�n�S��w�.��Z.�j�x��-����W��3)C4vP�T�t��9��֓ �SAql܂; }��M	B����yR�<X*xw�'�.j2]�I:"rr,ªj&���<�8�D���vL2��H�A��=��ה�Z��/y˖�ɺ�Q�1v+=M�����"���`�= jS�h�c �v��)����Y��r�Թ.-3�+����o�/�a'�(Y���D�[�R��I�?����������e�p�*N�b������W"T�k���UT^`��D��O"^��1��
pJ�eI:��]Q��9���bB������P�
 -\_g��m�*�1V?%��C�4}B?�!�������(��!#���Ӵ#o�PcZ �t<Ɓb��8��y-o��a��?Co!����p�>�˯���|����v>�Л�VOy�<�b�s/z�p��8;x�؏�X:����O���Þ���J�+�L����ڲ�Xk�|k���ZňR-��Ћy���ϥߣw���J��P�O:*ō�?�rѾ���H���K⺭�$j+{㔾�%�B�[{�����s�SI�>&�;uy���g�1���l)��+U�M�͋yRV(Pc�����b��_� �[vA2ŏ0S*UI�;<�$��v�ldFz��p]{]��W	��J�a(�s��ܭ@��:Z�I?��w��'���B{��Ն����D��U�Ǭ�Hu��my�ԧV;�ߴ[6�����6�y���`�B�,�)��h�"� ������=�b��f����I���N����J�wh��.g�O4�-k{�(��A�L����,�Asv�:U��(�Kx����M�b։zV܎3 ��N a8�G��7��TBz3ׯ+�b�{�<`z���듢��(��ڪiFH~r��~��b7��(� 2s>$��U��K���bf)�� ��k���e*�4���l�ʍV]��П4�����jf6X�R�Z:� "7���6�"Q6�2�5*�O��#V��~�D۴�@2��gu����$�0�110 `wā�a�@+���B�u4G`v�s4������B�n5���&�=Q���P��*��n�9��ZOM��V��4�ꤙ��bb��r�cM�%D�2�LV������ܪ�z�F��1�n.��ω�N2֡E�\���# �n�T��(ۭ�I�F	�H�F#�u.�<X��rIĠޔ��=���t�)N=��j�y2a��S��B#<��+�ٱz�r�p�l��{�By) A{�~<��ٝ�$S~����'&��ӻ`I� ��V���r���se�)�T�_[
��T�T`�$�L`J)Q]��C������4n�dR�����Q�n����H*n/�ɻ���նށ�)�{�v#){�ϖQl|��bP�D���R[��cNP���K�sf:r!O���"��X'v9�n�	
=%#��N��O�8�g�f�#/ὥH7Fݜ�9���	 	&Q?[ڽ��9������z5�<mid�܌|U�w}�w��^�Xx4<\Q�B1�I�|�>k(Y6��|z5����MIgp3{UW?y��������x���� �%��{�i9Ā��sW�~��}�xz�)H��b�""n<�ʹ�킲������^�45�޴��d,[�C�Z�K�C��\C�p@t_�
Je�)�m��jS�����(��ܯ�{��h��v={�����\�<��JF����Ha��E�����)qbF�iw�+������:�╠�7�E9���*T�1���TJ.SaN�(x�S����<y`�Ss-�#�zKKk8%߱���H�恻|�S�(�∼�@�9�� D_�������(�ˋH�L��������'L�&6*��GN� ���dnq��`_�y�YSf�=����; ��ռ��3�c�	1���ÇVI6�&����Iw��Δ���qr�0
��,���㒙���O��r��p�\��1y����#�q���Q ~e99Y�;���Lm����׺	�uh*p��4���>�3Ѷ���_�8*Mp��4w��0b���	!�ڞ�"��г�0�J���-.9���Q��`��Гr��`�~��
����b�
��ל\���h�8G�9��+�r�.0�u��Rt`���]D_����ǟu���B�Vp�<zVY�*o�'�JZ�?�ѧX�S�xܙ��ǆ���D_Dliv�#�:Q5� �}�u�'x��d�D�����D��,l����I��V�[��z'��<^���/�d�*����+���ݧs�KE)_�X���*I����~u�y�5w���@ci&>���AZ~����M\ze���<��D͂�'A�(4��8<�ק�����XN��E�b�Z�ӀB	����G��q��Ε齈gH>����w��l���� ٚ�	bp�]�)��%�V�;aIQ�nhÌ��[�*�Z��r�yUNZ����jhX��$��
���@V��R�':��sU���t\�d$���i��,#�`腧�C�!����-�VwP�X�E���z�"o��)��|栐$B۲
�#�'�\�B�������ic:|{��AV��.^�n�p��K���a�y4���0�V�S�a{/�Z�U`P8�NP�#��>������tP\�|q�8���~��çHES�.�Ԑxr��x�E?2X� �3G�R������KbU��~A:5滪e.��Ƀ�/sF�A�S��<`�0�+?��*�e��X��@,��K��½dR��X�{Eewn5݀�v"�rl��**N���.4`5��
�z�;�a��@��L#+|�ǆ����ּ�c׈L�b��_d!'��o�TO5����