��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{��P��f��Oz��Q�y�0"��v|�c���Tm:�o�~?L������A��!X[X��F�yC�Q)x��D���;О�{i���W�2���O�j"�K��y�銒��cnR��#���#r%C���q�����!�7ճ$���'a.���$��ܲmG�MZ���HŖ���%�������3HE)1���f����(Ȟhk1R��V�g�^�LĴ�n���2�k� %�S­ǳ ǜ�˴��@�):��*�A�'�L�+#�!b�bd�7 �oN�Jk\�Ό8�'��2?����[k�� ��䕕ꦂ
m�^o�v���:�u�DV^3塗ѸiQ_1�b��5?6n��}f�h�.��:K)�7��Ѭ��:(!X�X_�G7�ϥ���t2��l���ṋd��17���ֳ���!��ʢbH���%�y���,Z7������x�G:oy5�/ʔ�n�~��S%��clm=t�X�J��=�)K�&>[��8��W��W8�d��M�ڎ��e�}�1;q����6�
�:x�C�SƽVd"�������R���Z�/0�V�� ]����,"���-a�#[w^��W���\��억����s����po�Z�o�*�k�X�X{n����p�n~��SQ(nUGV�����8�M}����P����P����a2����5�d|R�|D�ɔ��E��n�1	��ivH%�S��>��b��[0���wܸ ���V|��{�n�2�����JT�S��Mx*��Wi����9��䠞W��!M�s>b�!�E���
#�U�Ӣ�i�� �:�*0$���#��b��%;fD���ɻH��4O���b��7Ad�6 \�s��� R�����q	��ӌ�@%bq��O����57?��w�*�y�"�B�T-WLU��@$��r=%p�ɉsᬥI�3����W��m@_+�"c�O`�Mf�P
�(oʇ�i�Hv�6�ž��%<}��;(�Tvwʒr�l�U��6ڝ���]��eb�Wt��;��19��Ni�5ڮ��������^���q<����L�*�cC2G�%G��|]5��N�؀�8��~�Ņ�����8��s%{)�- bI�$$��(�bı�ƹ���gG�Dz���>��;�/"�F��-���5�t����b��i��-� j�gI9DiBճ��o7೧'�K^��<݂��m�V�=��ɺP��J[>1yp�<�����t:咶#��҄|��L,/�n%FU�'�#&yt�J����@%���]�7,�!�C�ʻ��`�N�[YG�6�0��ɭ������3�|Ⱥ"�'u�l��َ��_(�f�9iBx�_�,�b��7&���=���%J�KU
��V�'3q	�J�0��^H)&ďN46E١���_��OՄM��4`��]��b�l$��^�_�qߘ,:�_����m+d�cbF���I�m�85e3�pm��tVWj|���R�Qk1��^S�Z��I�t?'��\f� Ҹ'�]��m;�Ix	��B�&���[i
ȝ&TAf���y��Sy��hR�Ii����;i�pӋfV���s
-��cuG�?���T��4�N���2���3��@��(�%��^�$��֖�k�`a�[�����Մ0B�aV��o�s�׶�f��&�͕rPx�O�:~����aex��;=%`dg�JN ?۽�������l��^=��������1�vv(�(���I�*�R��]F�+��^�v�U��L'-r;��*�.,]�&��S���ۻ�(Db�'��������g�@/�l�}j� ig�7P�`Cg�=��K�������vSc�,�~%`
R�0��G)Wǵ�~���uIh��8q%Me��*b�J������3(��~yIC1�ˇG���n�@
������49��ӓ��Rk�M^��>n3V��:����a��Y��@���B�����lzJ8�:�K��W�������E��[}gN�MHU:&B�!��]�5X�l��P�(͌%��@Nw�}�A�4�D���&g$�ՈF��$�jy��V/�͏����o��`S�ɜ�]���c�z��l^\]�gyQV�$)UK���$:p���-)�c`�t�Io�@?{16G�[0&Ð�p3��3�B��q�ouX
���j?c!s��X��N�UNd&,���S`s������4"�jW�"�b��J��� 9lO���`�L�Q�t�Z\�m��$=���.����T��s�b/i�����D��e]�Ȫ�J���A �8�y�A�BX��ٙ ��q(`	����hmuh�{�Y����F����(��()�l�XVW�kj��'J첨���E�7�`��>���v`ۚ�-IO1�4������SF�1?5�ǭ.2���rh�˶|��w"�C��/d��8S[06��d��kx��j*�I����^$2�:��Tg�̞30�1�m�,�ЬBYjA��Q�m��`Y���:b�����Z��U�\@W��ε�|��ʥ8�70� ��+��ݶ~��ۭ�����6�ŤЫJ����
�����`��PXeB^�˝�w�)��T����0ҍ�Ws{�� iY�����B�@��Mh#<4�����Gn�.	~3,�~уX_�&V^��9eD��C�Q���� �l�3��n]�;K����+L�hx�����r`�^r��~ܦ i���%2oVGu�Y��� #��6�|�@l�S<J���x,�ej�1q��Ǉ��*+���-�c�G�tQb��u�r�l��G;��� +c����@�ԫxŜ���O(��ν�[5.���p�O�,�ڄ�6F�Q���k�i�mS̫V�#�=���e+/r�IB�Ц��^q��������{ں��M�e\Bê�?�--u�c��R�1
����Z36gd���v"�3!��-Nҏ�5��;�h���l�����K�Ea!OV���`�(���/�2D���������>�v�ƺT��TYx��%�Bw�%{�,S��@<���<�Bۉ8ꭾ�"�v�J���%�	��c�i5Sl����X\x��Cw'�,\���暘zm�7�R���*���?�e��oy@tT7���EF�S�MW�vAĢ�}�+X�r*��k���߹]��E��Bv������PX�����SX&W�+����������~��?�=�Q���M�����5�9��>b�6���ȇ��%F�zI�9��q��x��œ���cH���)>��#=�V�q����,�G��ӾeC�0�p#�$�|6s�7:��L�l%\�䶢��\QOV�]�H8�焚l�S�w���c_�q�H��mIc���ϫ�~9����@De�R�����AsTc*¯�gSA��<�p���-��;� +���V<��4��G:x�I��N�:JAg�y:`�Iajb3A_�/���_�F�c�~M���2V@�^Ǌy���6b`�Q�t_��Ю��_I��[�L�Hy�!^�m�֋�V<�2�^��e��S h��[%���������ȅ�>�������{bY���i�m�~��"�K3� p{���'o��S��RvRY� ���Ӥ&�dC����cA��d�5����]Z��N67kfj1,�C�ߒ0�f���+A�d���?��]��XX+���o�a�8N�/x��)]wKn��2���a`\�f��z��ؼ	�y�FZe��#��,x��k4��B)�����B����q�_��D+)���ǘ�@r}�<�1*��la��`x6.��1�:�]İU���̕Y����9��:�mv[T�f����1����.�Z�Y����E5`��0��Q��v�{U5(��{������};�j���L�3(��o�g�4Ϝ�Tg~���7Ъɶ�{F|�od���ڨ�
�- o2��	#(-�2��52�����F�x	�,���g%2�kQ"�P�����c�(��Q�F��|�PM��&rSD(��R��3�A*�=6��;Ը���7�j��e�Qz�&�@�
���(6��Ҵl�Ŕ���b�QI&N.,�E.�m��(+(��+z˞|�f�hm������)[9Y���R�Ɵ�s�d,s��-�wN�Y���3e�,l�)�>�jC��1�T�I��~d<�vB���D](K7�XD��&xu&h�ʳ�9ݦ����w�A������}��3��>0dm�z� #�����o�Dg��E��,R3Zl֥����ɓA�	��"�g,���m'��^�e��Z���o�[�i��Jxz�kŽ�>i�"J��h��cl����j�w�I%����c��i����xO�o��HFA��^��H��q��W��"ק��<F����q����>؅��}�<3�����	��o �s|a\������q��Y�F~a9�)�,a�(�g������������Z�;�0)���/2����;6^��F�0�����;��������I.j�h2��[:�c�d�^�8����8�-��$]RjZ�c2g���|��bz��z��7;��Y�.�8�c� sB�c���It3R�ek,�^w#n�ҖV_3��M�v�3ҙ�QO���m��`8l�Q��H��}1g�������m��鳵L4 {�W��5J�n��nw�:c��3�Ku+R0��7x.^'�g�Q#����.�3��݀�fG-�V�\	w/�ܧ�| ��ۿC1�[�A��\�g��V0��
��=n�W�Q�X�g��c _V]%�|C/<���4^%��}hè������G_0QhXV��OˈL`l��12X���&�\��%K�[������̼�5d�zR�L���+b���0p�w�T�|�"�N��f�\���jL� �4�����>3{{_i��|[Z����;�����3�p���ŻEq�/\l�ѯ`�Q��Fm�P��s�)d��}��R��WL������;�jS:��=B�)���Y6+����sN`�L�wO1x�[�ː���P���JC��uLx��2�WZ{�Z��E�&[;զ��U�1�^���x��q��- 
�<�äP|:<�j��d"����J�#y"�?�Մ�h��4���m7/`I�l۶�W/�4c!�{���хSݱ�V+�*�������A}b�m7�TH$��7VE��*Fx���y�&���r�F��'i,2�4��	E@h:�!�|g�Mu����"-�ԍa���}�O�v�*�咸ۙ�����L��`����!�`����_fNM�����T����RL:��K�"���qa�|&)�7��Q�T�7^ٵƗ��"o�n]�����Y�k����!����<���`0����=�s} Ll#�;���b� �Ia���m[�yd�~��3���F1߇��2g�ɤ�k����0�p0i�c���&Wz��he�Zl�9I	�l	m���[�b���r?�wp�af,e�^��ʜu��V}�W}9J��u�*��Nz��:��p�����w��Kz9E��
~�"�����,�~OoVB��q$ʽ��4���8��%���MfE�>�s3�1�Lu�~��I'_G�A�PZ�l̷��w���P���;[��Ye�čyޚ������G#~�GA�����]:6����r���(9�I�[�~��n��	l'�Z�����%�ڞA��2�'�b<������@d��,utxG]��Z�E�6�|`�4����0�Œ�=e�*�?��9c�Lt_ �
���.��ز���T!�>��\�<[�c�Q�v6ʊD��g�ݷ�����B�8���[�^�(�ͫ�L���J��l%�����-3i���J��FA� �vwz�7�B쩒�ij�^��7��Һf��c�ۗF�ͱ����,�s�U�wYع�Ph����[�[꥟�x������"W.C2�o�i�U�r~$H��x@ܩU�׉�|D�HCζ��fo\
�����Yl����,���<	�F9Q�]���Gi�������{���h���m��E ՜���Ž��%W��ԑ(�4��x��?d�ؠO�a����OECd�x����qz�w9�\��	éK0I�hɯ%hcn���dq�ґk8ǟީ���d��|Y5����T:&	ҧ~��3q,l]rv������"H(���t�
6"[�uT��f��;=r��p�,�+_������	��oK|6��L	hrxe�r�hNKO�]�Ș�C��;Zf�倚�'���kak
�u%���7I�( �;�~�w H��T��,s��Tz����^l�u�|��B~�z���Еh������T��������v�	a��*.40-�瀣�N��wdQ�5�rM��d��~�da�ܰ��}$�VH���TG���{�ՓQ���b���#���2of���S��d���vN�q��;�q���^T�i�7����I�8���ҲV?�Uy�0F�n�N>����8NA�G�
�8�x�u:�7�L�7X<U`���K���?�3�o$��Wd��(��ʂ$\@��=4�M�{�d=�z�c�{�(m����ÝP�D�j����V��}A�V࿁[���ɪ�ZX�ڼJ�!�èU��g�YP�?V!$��B�3�S���qxDR�d�2��~ ~j�"R\�A)�Mh�}፼�����˓F���:��f����"�i��I_���H�M%D���	F�5�0u�cU|�r�Bܨ�K�PlT�n"�fBE��j���������H��l��{7�f��qu�K����
�� ��M�����e8o��	�r@)ǃ����aʢ�4��H��nH���� �(^�|��a-�C�I����FO?�x4{,S���0J��W�
��,�[��Ws�S�����U�n�|קN:����3�ڦc��{I��v4�/~��#�4W	�3� �T"脽�_�����4����QRՅ� u�[�����I����7:����dS�,{�`���ܭ+~mU���hF�nh�PYc]N����(���]V�A���]d��ӯxP����84C�ܛ�c
�af|-gB����ӄ_��BR北�f$MkQ�;Į����i-�I��:�5W�H����U_M�f}�i�D�}�s�d�OK��e�+�'�kY��]ʾ^G���q"44�B�[Ϝ#$���A�-��Ί��e�b�(S-���ρ�h�4Ff��]����r�֟��V}s��7~�s;�5����Bh
J�O+	�����+Lq�!�L�;fH����L"�	�أQ�'�.�i伲��m5��ķ�R%:�1���;5�h�	��۔u��_�$2u�a�=��n��d�>�O���	�V����1�.�]ʩ�Է��4���L����g��CoS�L�f�#����'��E'8�����74�h����XJ���w�A)�M` w��$�^��,����������6isﶃN/B�=岨�*~ѯ�=�(^͔�����8Ts@/��v� �ܛ��\=Z�sd��i(�<�N<<� :�?}����ê!�u/�5Tr�gIP���n���`V_c ��7�G4Eߕ[Q��2���*C�9I�:�d��S�zm�'.Iwb��L���o]�7n9h����ĩ:iTD�-c���B���\�2ˆ-i*x�+��(Hó9�B��E7����:G�6�t�J��77}��fo���ѫX@C˰N�b$��:�_"�U��ęk�-faI�'�����@��G�Yg��a������Z�����C�����}v���OaOHTƏ!~Ƿ�����y�����$��^@~^�4���o���.��ө���Rü�'�i b��M�%����U�-!���%�e�=�Nd�������:P	u�>�6JeF���rΘDD�5�ۈlG�@�ʣu����E���m�r�t2l�`T�;x��8�ǹ8�O�e\͐f;�{}����W˄?�^�I^�#^5�z#�w����Zl��M!� ��D��ZC��ލm]�k��>��HBFW�����N� ����h���Q݄>X P�w:�K�Jdb-��U�p���&(�U��Z�lOɄ��\(wK�_4ܶ�������6��T���0Y�$����Zor�ˢ׈�V���B�P�-��
�Q��[	��/��� ͮ6`��H����2�	&�@���#��[P4���z�t�ok�1����g���q9�R��rr��J*ٛ�޳;
4Z��>���\3uV)�[:Moܪ�A	�dN���'���sp��(gf����綏���D�v�=1݈7Τ��VZ_�%�yvk��B��-l�%�=޲)(Jb��Oq��{�&K�I�C�\CX�l��G�X����>���R*m`�I:���H	���2L�U�H�C�h�H�^�LDv׋�e_3��}�b���y�1[�6a�[��`�)0|�e�V���'�l�B����b�X.�kI��[tDcUbz�l|�<�eR�|K���^�����^��nO�6[�-�դ���J/r�H�޽��P����I��,�i�\6���V�@nL���>�+��Bo�<���� �����;���p��	��&��dTddMH_L��`���F����)�4R)��i����1Բt���X8{�Y/Oыf��z�I�~7A�Ƽ���WP$�p�� FDm
|��|�5�M.	VtD�[s~>�����Ǟ�]���	V�N�E
�t�th��EnT{T/YZ$O��ھ��Շ������Fa�`���UNn �L�y6����VC�m������?x���$���(EVȃ`��ѡV���{����hq��`?<�h��8�5��6�pߓ��[~t�yN25�؅!n1'��VA���g��~.wf�x��`���	x�����B���~��O�t�7�.������.���h�t�\�C����a����fHl|����P=�9ʈ�Z�[��b�M�����L#��~e����b�HG
+Y��<U�"ӊ-D,�%�Yi\���tBMq>r��ӑ	��ǃ�́�=;ș�OX�X�X�{�#-�P���z�Gw"f�m�Ed���lvp]G�&�@,�)���iG�<�����vEme�Hk����0ɶ������峐iw/�5�|�Q���os9Z٪���i��#{R`�����F���$�6�7KY�R	�3-:
P��=�͖X�B��"jF ��!^S���r�����w�o�O���<�h�
�n�:sE����;��U��r8�u'r��L��j�E	�Q�`&��\��ig�'�oY�m�h��5�f/f�@.��A��!���!躃�6��v5�E1�wY=��H�|p���7V��ua`,Ɇ[13c�EeQ*\��._�B����OFm�УQj�E��e�Y�u�jA_vE�0=U Rߛ�#�r&&���^?Z����Tm��Y�'�`�A`�ֻ`�wkۀ�ޘrP;w�Q���.�[@@�7�[��M���H�c�O��a4j(B���
�y�]ivо����������x��"௉���R��W�T�f��x�ഖ�oM!�8}~�X�ՅNpC"��g8=j�����ړ��d�4�yx�a��� Թ�v����B9�0ޒ#{�n�k%�a�9V�b!p�3 �3]��$T���k��0܊�c!��(,��] �̛��i���2E[�?��LV������ɹ���L��3F?2��\J�G����Q_�ܶC�c�9� ��k��E�=w^�:RK����$/�$4,%P�c���37�qV�z5W"�8%�mx(0l�d$���_���h:1���t�W�@���#��0��Y55���d*9T�<����\9hj�=�E�
�径�����dU����qX�Tt
8g�cڂ�\���B�b$�YN���@Ӽs)�&�_���K੘�v������N��w>�������O�P�#`(�s�@��+q�"��l̆��È�8���KJ@G/�E�_��'Vc"�y��>�b�����?����՟�;yS�CFZ"\D}HG����nBt)m�F[r��D�Z�Y��S/.��i�},�������,.V���"�Ç5�,NO0>B�<um9W*n&��q�Y�o�2��kP8�L�F5o�
�VE`�2s��#�
HϾt���1i*,�3�7B�|���ݍ�:��;�}-���SN��b�6������9��	���*e�/��z�6�'���R�|���|�P��Kx$�	N	���PA�t3�Og0�m�P�I ���2��� rby��Iˊ�Z�m)+�
L3�Z����^
�6'K�N�H�z��I�lS}L�y�����Ȃ3LC��N3�P����W�Y��[�����:����P��S�����GX1�E���>�س?<�.̿�vE�mJ�OP�*8�