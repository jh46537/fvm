��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S�VJ���ɾ GK�rA�!��}�x�E}ݨk�fի�u�(���L K߲w�.L}x1F2�#5H�:�'))�6_��\j�S��W��w�.㆔�[NQ�6��iM�@��9��eh��L�@�Fb�%FZ�"e��R���W��@�s3a�����膂Y�:�D���!G��j	�E����}��Ui����kh稯ka�"������e�^��6�ɠ�Ij��-���jW}e�@,��=��\�`�Ǩ��:>_2�)����������t*�� *��%/��X_0�2�KwS9�ڪaԟ�	�踷Q����Z�@Z|�歊�)���ܰ�K���"F�"�;�ŰS�d&>�،4j�o�9���xD��h[JH)���m�tS����\�ɑ� �n�{ƒ;PM�����>"s��R��m(ɠԉؔ�W��6���ߜ=�5�%�_��+*�o/�Wv/�nW�S������50�u#�����=�O�3b�w��Z,L+F=5�'�?y{��yN�2���D2�m� �p)*�CW��F�7�Ye�ȼW�xs	p���-0Gnނ���Q��	��q՜o
����D+�g��!!|VeG*�s�1� y��!��FXV/ao�
Z�#o �xE5�_�=��جƒ�K����#������\?xi`i(d����#���&S����$��a%�o5�H��}\�����?�ՒI�W��+|Vz/:�2�T�K���f?�k��A9���d�̺}���6���K�����T�ʫ�n?�塲������*}�Y�9�{��S���c�{ҩ����H���qn����qh��W�"�&sL'4Z����B��,8��w��BFd�8M�Y�b�oe�Wl� }�$�ՇD�O����r,���1�υ�\\v��<Ɗ��h�L]@�'�Z{�e5��w~��t�qJsP�X�q)��"ˀ�-׍����������@�(� ��bx������O�3�Ӓ[O[	�Q�����c���x������_��˸)��+��hNۚ�-�4�G�[��T ����r�͸���6�GY����G��E<Cn'C@>^=0�DFj_�hEň�
����6Yv��ݚ�n��r�'U�d/"�OS����<�N[�-��������O�oH�Xd�K�qF����mʞ淛�vKBDݽ��F*m��W0��iH*�SM�-s��a�fո�5/?�ز�yw����Ʊ�^3�T�%��ޮ�~�N'kK�u��M;�&8&������0a��B��{B�t����@ֺ?n~`š݀۱�
���
��ާ���2o��E1��*?�X ��1֐��g�0� Z�(ӖrA6��r|�5���"M��� �zrU�Y����A��-���Ӂ�Q����Z/*rl8g���1tFC�c���$	�����K�?������5w�"����xG��i�&�k}�k�*|}Ӣ�#K̉|u�_&�o@&.�
�\��w���ߌ��L�S[ {��3J��2���F�م��%���}~t�:���]�;�q.~��j�+i��L�_|D�s���Qa�!�_l����=->݅�����()�L��̾��94�ċ�2C4�N%�*J��&�+N�,'/0�^,a��]S����;�A�H�Ȍ�6ua�=����F��%T\�4���K�I�2Ӡ��R�D�-nt^4�P��y���ڹ,]�j� <;�f�I���\JY�Y�����Hu���RK�C��p�2k�a�M�Ǭ�uR c�H��(1����" >��[:�
�⬿�(���r<3Ku��K���{�/�6���w �z��݆�����-�u� R��o1O�[~�����?�b��)�9��L�	l�vh�/��?�g]be�*N���)N�W�ZK��x�)`�*R����6@ID`����vFګ7��*�^�ck��/�عx��Q�
>�]I}�b�&D%YD�E=�-������m�c"+�d�'i�,R[��a�p�O�2	6��c���~CÈd�BRAڬk���t]VKĕ[�ρ~o��������1��>�t����c��x�X,�F �h��������ő�s�֓ 
N/�m�y�VC�����B�������e��ѱ�nBx�P˿����H)�������p��W�Ϳw��"���4�Z���?��m���
Z�a�&5�=���Ԩw9�����j�����5mM�׻-�z��EN�C{>�@/�Gd�:%xə:�9,���̀C6t� K�Iγ�.�����d�LX]9B8T�R�����l�^��V�ӆ�i��4��g�s?AtH;?�Lw-U�yg���ủ��k�0� �"����<���o�dƗ�pBg��#��r�a(��ho���V,�b3�u@2dk��'<�t���GcV0�]��,��-������iY	u<��F�{t�^ٿh���ƃ��[{����;& �/5|�\�&�3M�v+@�yNj���-����D��9,��������Щ���J;�<�$qkbf�<#�7�4�ҡ$�ҫr �4�B��j�<��
�`,�a����W�˸o��g8��J)`�U
݋�VϘW�4�E��Z:�g��?��eJ0�mrv�6uH��f5�����7�F��̼p"` �)�Dj�51i����	����vb��A)�W*ƾ[��C �Ж ����<��w�F��^2
�O��b�dPI���B���oWEpc�_��2�"?#-p�S��V��#�� ����?N�ŋ��]��W�"#s��̢i�M��^���<�O[i+�+�0���+8>L*#otEi3�w�XB
]�:=�0/�f���P�k�t����VK5��[��Bc�y(�7]H�D9�8����*�}H�<9���9�+|�}�*<׻f����N)u�=�]hS;P���u��ڒ�:�K�/�ݍi��M艳E|NV���V���虘��]�8E�@u �J���}��/�U��j�S ]�e�~X>�J�=���2\���.<���u�y2CGĞ�*�*I�:װ���J��Q�2@ڜ�'O�i�E^m����A;^�x�s�=BG
������K:1�Fd̛�(��8�� c|(V�*�-�@���u$8;a_�i�AJ�2�
����I��Q�{Þ3˷�Đ?J�w�}2�f����r�?������^�	yŒ������{�\-K����N���j��&6�/�����J���;r�e|����F�bT�+�t�|<�&Sť�sW;Z#��M˲u�DY�:��6=*f'���OA���&��nn�Q���J.~qM�-�9P葝J2B���zEъ����( k�H{o�8�˓>�G�rc�A��ȥùU���S�$|���������������Z�,(ž�u�lE�u�OF7UXxN�慧��q�n� �Y�����/b�Y��Q%)<t�}ᗌi`h�#j��Ξ��6��囏��/���|Z<�Ɣ��������u�J��z��c���m���H�>ѫ63I"R��֛P���^�@t]f����_���tv��23C�)i��Y�d-���E��D3xU��+�E���\���^�ǡ�L�:P�������}NT�N쁁��a����N#�����P]9��4eh	,�횣D�36c褠͛�,��XQ��Y��o�"��9(N�,{��I��nz�3^���P�?aX�2����i�>�Ԏ3��=ݥa95��	p�W����G�j�e.��1�Z�e%��2�u�iRIB�:�^z*��ef�Iy3Ũ�O�t��}���Y$q�wM����a��������G�f���Q_V�e�ш��m�0����
N���	�"Հ�O�N�)�mw���Q�s+?f[l�*��ƫt�W��Jr,A%�D7��K�.v�:}�=��7S�5j͋�
a2�������E>��/��vLR<O9a�Hm@��n���s��HR��P�	���P��٢��F�e��x�)�#�ǩ��.�ډX?�4c7����@.[�UK�ы�{�.��p�P�<���BFu����D�k�B�ڃ�9R�k�u�
���k�U�����EOM9B��s�(�:�.��Yփ�{���:�, Cg�U���6�2lԡ/����Pi�.���M�%��o�3m:����s��܂K��o���!4m���	9����dDT��է~ڏ��6�����d�d�e49�'�a���.M.��yń��ƾ�	�(��O��]�X��,����i� �!�*XX�Sa��0&vR	��6>���-BR-@�>��N-P,�0���&(�U�_2�]PI�Dh7����U�x%�m)-��� t�B|�����T�+y)�bmS&5��~atX�]p��g�N-�N�2A��xZ���:I�汹�EđV�`/�Ũ�`�%g�֛7t��Vs���qL^�\���+A٠`@����.�9Ȑ�W@X5�A�u�����<q�G��x������K���T�c�W .�mKo���"�l="�sO�-�b�#U�[!��HL����H1��Ah� �ǌ@���в�k�	��} ���lN�TW��Z��:G_�FiN|�@� �%� �`����#����7�>��2���f�_C����n����	��Η��ڮ�@����I��7>4�3+��w�q�p��P�Qפ;$3G�(������SG�w������9�V�_z�P��i�-!]/�a�op�>�H�}�����&e���߇\�3C�$nv`G�����b�6�K�a�-}��A�̈���20U`6d��KUs������^n���ȴ�_�l��:���AΔ���C(�j��������@��NU��Vޗ��s��3.I�lK)��;����F�آ1<��{^��#ms��e�tʴ}ɎT��(��?�S����a��̽�4��n!b�m���,
���L�}M�*�TЈ��G�-��FA4����z1�2
(Ž��ק���,�Z|N����*�X3�U�]��&�*����m}&-�ht��I��⿄���u�h��D���� cϺnE_��Ug{ĖCS1�?�{����s�o$3F'}�%m��s�;��?&9X������!C5�S�W9��j北�ML�lٜ	h��Ը��"�g�X#����7_�ֳs��G(7�''#<�>�:п�T��L���9�"k��be
7�do���Lg���xQQs��8�4鴑��l�h���r��S���Y__U]���_�I(�P���gt������RFN|bp��`���������&��!on��n�&³08&�t��l�����
�Ψ7�8���v
2���B"O���%i��\�s�H��'��|��@��eZV=F�Ԕ������"�س��9xH���P�(��Xt���h��;r�^���V��D~��*��{(�����_}2��~U%.'��Z8�	{*2ͺX	91�pL��U;�1A���6#(��=�;��ɋ��4�	u�xD��w���HW[�
�!�x=K��X�K6�-�M�>��c|�M��$��	��{;>6��l�A�\z����ժ<�HX'��)
bR��:x)��Z����|[�E��6�j-�m�i�;�`���q��/�6_J����q��X"#��V�:���4��|���O��,^�7W�:���RYl���	>��+�3J�����ԘrA�2�YmϿ�z��V��R!����J^^P����&��b��F��z7Y�U�uvcձ,�N�ѣe��S�ylLV�K�~���n���y�܁�3�i�OC[����[x�%��d�+a�ª��I��-N8�/��@�"P��WǦ�׎2�;"G�OYn����u��5����/���ï1}�t|9^r?;tSf�?	��[{q����be���E�}@W-��>���e9:�_�=�wb�3��2N�k֊�]�G?/J�b��^�d�>+�#�[�L�W��/��O1�S��(�{?��'��PvY���ݦԃ-�l�?Jf�q��ѷ�eﷹO��u�J��M7@���I��g���bM��#?pK _��^w?1 ��Z��4�W����rg��U�����h0܈�C�W�9L�\*�ƣ��zOH7NfL���K��x�r>3�-3jE�&|k�A�x�+N�-����ݔZ�����?��@�-�nh�S����i<�	���|����Z'��h_m�?6H���W!�����%/|c�ɜ����>�_Iײ�Zc��.�S,�@8!U��+�a5��@{����F��:�v*�_��U<e�i8��L��bmH4.Q^<���28�ZǮ}�q���qp�ʧ�a��s�n'�_�i���Ո�	��ڪX��U
ė^#�Q`.En��a�K�<�<�aL@�t'd���NW�eDY��Vp��U��`�|jX�]�̂{-ְ{����5��_f�!nN���	����N#�t�����{���S�k�v��o{z�Ӿz�^��,
9>*�O#������Z[W'����<�Ԇ�3�-`�E,?	[�hF}5�S��8tȶ@�ç/!�������V7�Nʐsÿi'6j36��_/d��*���+�B1V�a��D���7gnzP��g۫�>���OK�!�I�;���,�cf���Z�Y\�xi���C�P����~��'�� ��_��D�h	l[�l�s�l��]f�XÛ��cil��|]�z�qȊ4;����=�����Z���E��,��6�H-�C5��k��b��wwM��g�3 �x��iD<U�$���J�I��:hXgEb���f�֍Hߌh�z]�f���%D �>l3�OJ0Š�}8!I?M%���z��.=n؋f�,}&�&��ה�@��!<����h������\�<��7*K?G�œBL+>xoU����l�KB2� ��I�w�6�o� �G}̲S�<Wf��N�� /*H�DR��@3����Lt��'��?�jGز�h��� x�}�i��BY6�^y��[�cc�����ͻ��Q�����������4��nrq93J�k/�_I}x����#�Pe\�,������V3I��!��xNs�0��Z#χ�0�`����bG�M-Z��oL�3g�A�U�P��r/i�r=,�y��{�4ږW�Ե�i�G��V�DTyEk?�P� @n�7x�)����������W)�s/�f�ߓ�4E�|s~Ļ�m�%