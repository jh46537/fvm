��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)��ޕ�M��T-@���U�&����pi��3<��T@�ꑭ�n I�F��)����N[N��Qo�����N���)���%L䜇d\j<V���&���u/b�x:LN��ɉ�iT����_������`��.Uwļ=o��Z@pЄ,�����9�����?�eۈ<_�1U*�����^L��\U�t����]1�:���R\�F���j-8�u�����{7δT"³+��˥�
��>zs��U�L���P�i�L�c�-*rr+�4�t�f�����#�!&�����=���"v��A����BgG3��pϿo�".���Jռ���9�<+0�!C\(G�*�|Y��(�Y|G�H�F���L���Ψ��SC��W�/���`��(zt)���EhE�)>�kw%rqB��qN��
~͛��G��z@��)�(�a�w����[�Ʊ��F�NU��Lx�m�Ma�rJ�-:��5���(?�����/.�F��"��Pצz�v���WD��~����j�n�V�J� .S5��%�ӷ�Do�&go�(~��4�<��j���	�?���>f&����$���B����5�0��e�(��ݱt�ˎ:H<༄h�����$8�'�o�Z�8.8��MaQ�2�gQ�
嗡�r�(�_��R�[E�i\�n���4�b\�XV��x6�bW����%�/�H`�yy�os�n��s���hP��l@&��H������-��Oc�v9I:O�L�	�N�q���Ƚ�0�.VR�-ͫ|q�$��	6w{�9E}�����P�K~S}�� �c���a�L��d�$<2�b~�_���&+��AD��?�k�>�{o2���S�	�??[%�C��<Z���_L�/-�)o�ןNH@�vD,+Ҁ�
Z�Y-Ěs��e���,�a0<fZ�f8]�ciBX��'�1qZm)����p��=����؜��2�1�i�A����-@��;�d.���Ԇ1U���YA�;�M��̶�*׈{!��lm�����9}}KvaI*3��Z�rҌ�a�D�sO�}�,G긱>ea��DӴKj��ih���9�6�-����)�t8Rɔ���}*���6*��h�"�0 �ﻖ06j�1=�W0S���8w�0}$�T�ÛF~������ -0�(��Hp@&K%6���z�Ѥa�,<�#����e���b��Ǯa�s���(�0�݉�ҿX�>�d��zߨ�΍�EO)��-�@�j�>ڦ__�i��ś���W�wj����Qt\�Β �.�}w�D�b���ERO���P+���`^ǢA�k�n���k����������W=�ג�;�-螌���|��IIjM�l!2|��eM�S�&�GT�a�O΋�V���'���"�ϼp��q�"V#9G��Y1���\����ղƯ�RD
/L��P3�բ��+=5�������Y��v�D�(����&4+[���ר�2$R�y�*q�%kP@H��?E$3Ee_q=r��P�>h'�}~��[F�8m���mEn�2,�SJ�F��w%m0[FI�W|�u��z��o�a:�	ɳ�;��-~9�R�~U�����n1��#o����~��j�΅��]��٪��B#M�E0�)�)�uz}�	<�B]]��B��z���}��|_�@	��Y�M��`�<4�� ��O]h� �Q��
��j�@
�/��5I�B����te��&ͣh��oְ<�]��[��%�!/����	q9�L��ReU���>��N�*��9�[!�k[Z\<���Y�����
�ȮB1��7��#c�����yI'j�~ԛIH�DdY�����7�@%��V��7�Si�go�f �qY�!UB3S��}��\���th��=:~_���4����l!GCo����HH������]�庠"���[s���z�����(�g1��:�t�&�7J[clS�ɟ�t`T��2i��3�lH���ܟ�s�i�-���g�֭v��h���D�ͺ�]y�W%�KaD��8��ʫ��.TY��m��-�����Lد�d%qb�慎t�оS]?�i�`�gI�%Z&>��@C��dpe�^)�đ�f��,���qQ���
�we�
~(٤��<<H��Yܥ��5�2w.������?'�~���v�!�K��t޾6!Ϊ�x�Ŝg!�Q!S��M;v!���/;�����������=H�ϣ��/3$dl���k'�np9�R�V�����Z�D��r�,�k�B;�2� �]�l�TLq8uQ�
�7O�*Ud�%�I��r/�Y����ǰ%#���D$Kȩ�(�2!�0�+gY�W\C���g�� b����F�l)Unm��� 5����؅Ｅ�*�CYXH�/�fY�e������X���K��!��p�oڄt��mHК���E��x���*����%�^���RB��w$���h�,�,T�����n���{�Y=I"8Rh���� 3iY�l� �F��K��)1G*��[f\�p;-^�Օ����Ɲ]�����z�I��ӊ��x;
����B��L����{͕�n���B_r6&����I~'\P���r���$!a�W����sH�����k�j�,�Ʊ���m��t%M0�嵓�bp�������D�Թ���ĕ�c�!��ᴧy@��x%[�:��*�o��T�q��
�xxd49�ַ����;a�ߞ��c��	�j����fO�\�B��_U�?�Jgk�ݏX�=SU�߻�R�hu!Eq4�u�@�i#����2��m\χ�?3��L�";R}v�!H�3����\�&dhM�tn=kV��F�2�v(I� @�R�y%7�Zq(y���[�=%�1���O^U�8�0,����A��MH*W��\��*	��������a�X���h�Q�Q�a���Eg��i��I���N��2������n�B���	��~��,=M~^B+�<�j(���F��9�N�+W�KS�X�J�T��ɪ�W��gT]W w��%M�������u��m��S7�Y��_��Ȏd��D0.9R�����RO�-�f��2se�8|oa��9��	7o�4s�
d٘�v�0!�l���cG��&��T��қ���D7��� (u�]w�8�*��QD�E��N<�ʆca3ȴ����k!�è��7����{&��ծN��e(e�xu��[3 ����w ��G���������*��(_C�g@�t��4�<^��Њ(��Gu8գ�+��6�_lҕV��y�l�>���f��r�#�9�󲓹Kz
.��[d�2�P�A�ŠjgZ6�!����g�R���ռ��w4G+����y��|�.hs+����4�M��5���۴'ZfN$.�k��i��'O4�M���Y���ۿA/��nT@��-��Dq��@ !��X�~@=���bX`NZD9r��N�#W����ù�+V.hK�]Z���P��� y%�0���혉mpl\̞�V����� Ly���d���9J���u��&���e{FX�<YZd��%C�7ꍈ_ָ� U�A���o�h��x-�sjlJ1��L��7G]�Ey�+�ʱH��uP֐j�N3���f�s&$�Đ��fcv���5 3�Ơb/B=�Wr9�+eZtt�v���8�Έ.�n d�B��0Bylդg�݄�v�Y�q���?8�42���\T�$�F"�S�nJK�����\�s��v����f�z�h%��C�9���\�ZOI��=O>%#�<6��g(�eJ�0�V�%�f�w���z��