// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
htLgl5Ha9qO6u3oCYUFZRp38i77QmQxAbGhZIhqubZ0TlizoJ6ECEdhE/ITEaICc
P2IixI0oMw3McBXXDe5bktiaUZ6UvXU9XE+t3cchXloItJXE+Idt8IOz06M2X0cx
OWjbXYHDHVD6urTgck1MIHX7YKrUD5C1NX5B2n9KZ3I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 43824)
Uz5P/8aP2nHlrQaq33JStijiAB6nGVoiqF3xFCK/f82dF/2Qs1gGaM/k2ZKh/+rr
gqbZX7DF+zrvd8R8xd/cF9dpgtUUlWvPNX8SOM6Ht5kHSckjWv/V2q1vqd4OXwzS
gz48GVIEsLDPXEpEu2veksG85IJLpSpWIK8JoCCUiVbqo7+etUomtf0A9RRseIEc
uMEK+eSXaw9qgCrsk4KlppI91D80t+xZq+sse2CnQbUyM8dtoqX+zf8ILixdo5CZ
OdRUUUCzuyHpYvNZ+IwZTESEZSJgV4Q/ewD7F4SUXvTeTMOY9yXJcmkHEs4i+4Sp
n+PiN/PsXpc0+vp+arIrzDgPclNn96ls1EDyrjPgQECyW3XN4thso57oNRdxRgEr
JVer3TTTFquLllAk6P9JY9p5AZLh1fTGNnxoVixJtQp7OcxbIgKVxO3trGztEPxv
57is+XPHKPVUZCKdXD+I16/O/63aOrRy8K4AaCifl9qCpSPma4VVveCjF4dK2gGI
H4eG9O1rqMw9QmwMw7UPDooTxlTXO8khSvzmNNKdse9JOIoyg10w6q28OfMPOD/0
irxzAY3XWBvr28IyKXA57ZqtUAxIWu9APHUldtehHuoY2b74grNlIHrgpQ3KKa0f
x/ed7k3Sib6o+MQRI+w0sN1fsq1jAXPy2IH9OTsN7lBDkyjLs0clif1Z6AGCCTXM
zAd+pzh9cdWXdErX6LIggKXHkAUoRt/7gVjJMjXZlrT9wJ7kaNl8FhzgXVp2SWOt
MN3kXHvliagO2pf6BhswGXbQt4yTbdRp4HqgPs3yi+FkmPCpv4+O1SHb/Ny7Hk0R
lcDI6TviPpFz3Xf1oDm2qWwrNKd7zsG68NHuow3JOw2NFqu1XYpfCW7ne/ybofu4
MVjxEesyHdCeF7hIlrmsFYvUgBsVXWu3dHBSYoiicHACcyAYgPsrm0gCkkhB6VJZ
vj2xuLOUKKo/7uu6ROopkv4ZoPYFZNtKQpTzwx8qi1xnvsZAV4uOV0PYxG1Jn1QV
zGvJ8SlAraavuX4oi7jgWR4XfP+zTcALAB88OuNubQnIObehsKQyBEtIWLyTw3cS
cH2PwLujvH02NPJJpkLVV22dvgnlyAI7PncPVICngtMzAWzb/pcK7rJJXjg6yV/X
yeK0PM8mWzqkRUp7ViMPmuNk+vaaZBTgiTUJ1eGyunm9u0SXvm0Z95Tx0ejrWBFK
PUwtG9U1PAY/eE5I7DrwLMrT84mTJm6ItthO754c9A1y6Ve3AOEpPQZ/fpG+xpSD
0t8roH+vaP1rxSKVX07frQilO6I7kvnBj6D+h4JlR77rx3W84z9R4G/B73cIdqnF
fCQlsthJV2su/DNxiMvuLaNZWR0T5n2EGULpOfC57w7eCDfYDT52pTWH2c+va4Hp
drJXYrQce/TPil4fxD2MMT8mF2SuX5aJzxQ0A8BaMcZUo+e+Xw8VfuJkXomzpbfx
x7fPEVTahgV/Ga/n7TwvUeAFQk17FOzkzf3P07EzKWQsPtBMbm1+VRfSKOQU2lwW
D4GQXT5WCJJOpyNIQpDyQWInJ9LUT63Mh6BOWTwWgU+vTFkGSeysr9X1Ph99jrvT
Z3yVU9oFuCewiEqGbz7RJCmLJqsUzyO9vehIec1iVudvBFeLlB1BspdlxEuLTdG3
LI+pyPfiVAmBJf0qbbBsKxRACKvGgxbY/M7fEcW5jHHgHKt48OH71jXkj6Mv17Cd
pBWp878HrMoD21g2Lt/jkhjY9k7qij2ZJhU8uISrTAPilWWFAuxMCFEqlU7QkSaF
peJLYU1nJxo6RatMrfbCtfwHpJ8QM6V2gvwLByvBb1WKfMjH16E1MxQCxWnWkFNi
Hlc4ZMbDuKkFKQ30TF39Uz54Q6TNPqZGlmoFEK51nDz0BZ1Nec1OsZ7RRHC9SH9E
X5jvxy9onUpUg0SmCw1mW3Hz5QFuVUqv+sSHog2SI6HuE0aTBj9qTumg55xYV0Kc
v/p6n7UDkUcAG9Mt4AyavFPtzfXrv2dSdVHQSzZqIH1pLfiXbhhDJVpZ7u67CQOw
/rycJk/BtxGNWDLZNDqYDDhBmNt6X9+cW2CJ+eyva4Zz5IzBQmvEG0ktaXcRkAM0
hswkEN7YJ/E8SYVxcD0YkD6rQZm1mhPprn6YD/TGK0qv/bdwyRjB5ek+kAYFCjoe
VFX2B+E9EcUul9S8DJ3caL7/w0MAOtn8lAkN1LBK7qB5UCscQsGx6Spd5f6O9YCn
7vJh9HriA2SD8hc7K2ELaWwaIfTsNUGrsq4K7MY574Aa3MSFoGDg8Wb5hVfLFqxT
wktSvm2u/PsLWti7KkMLKPT6DvCFaPW3JImzHKnsau/vOrmstESduK6VFFNNoPUJ
8Sm3F0JgwTaUtwaWG2H1Cdu/dvDDulSMI7Z2WJ1Yfq3l3BxGDgY2vjmXItVcxUBH
1sp951JTNxhjLkGu4p+gW82thyoifkuAQc8v1YbCBx2DWYtuCLYuuMPpDDtAXPBN
7QjJqCw0LJunrlzB9Awgul/DQtniTgvLKYHmJsThchkc9jJ7AIug5ITIV67mCjkC
+ANH+cwGhgA+3mqm5oIV+jpyEOPWyt4M8Nyl/x0j/PKkCOgSZP4vOU+5X8sDj+/I
rWzsNo8ezK+BL5/1dNLOlXcT0KNn7VAvHqy7AxeJ5kc6icPFzPvxqKTzNGcYG7lJ
GKz8DBtGOB8HFp2aTQE/SsjeBebJUf2HKYHpaQMPZcklxLce8VH3EqmudhhHlkia
6SFuykTMhxLVuotn7HloruCK4vNCri08i2nNCsJQpsYGMrOGLXu4vz7ZdZV6vPdG
98cXd4SfKqv9pJxLlyWTFePhOz1hG3TXLD5CPMILJ2l+nL5ausqO/mBBJYjGfaKw
yHFW5tPigFxc+TB2IksXIor3EfQeysdXBmjlGWStiM8MpgSo6h3CwTH1Q082sc9F
32xqDX3lojBX1JZ9NoRjc12xheYh203x0mMfMj9eKlfLmtS1lfknOJaHYOotCraJ
0bS5YMF4lgzabSGcodd+4R956TiPyGqpoVNRYrfJdISTjNAFsdSr5UPD0wXM4mmh
ZTGVh3w7hWEGyvy/PsBYU2kGVoi6UcRO1I9VdwCCfJOGerTq7bzgDFzrgIBLbP8X
cPpyOcHi9W3qmBrARt/WwqjO/NhG1RL40dp7nocsUOedTtaqyrhQuTin72i7uO6O
v8KZwafgwza/izuZQ0+VkrBRi+qcckAU1RR3BAR56LUP3emJZeAV5LEYHOS0PGrk
S1cEsTpGH/REHS3wz4KXU4Rjhb+ZjZgBk2+39HZUJP5b3JdJLOH9U1e6UZjq75OS
7LyGLt+Zin5KX3dxRNZin170fTUUKu4xMe9KAsr7ApCKLodQxpBtxiBDUgrD0Dlg
Y7O6yA117cY4fiKlD5Stb77LzZiiZQQsjF/LkL5YxS7HP+wi/WYkkz9DAVf1QokM
vfUm+twwD4meDY12NAc/2uCSR6kzfS0jswS6QrJqvkNIdi3rUupM1JztMXNDfeJK
BZQHveQWEu/2+pabo76shA/Y8xL3eRThYXgMD+RaWeHroL5WcjW9S19+dOXoJTa1
hFC88PQp6K0IEha4KuNYYR6+PgWui66aeoiwIHhiDPT9vYf1EdangKqceEOsVByR
1lTnZKxxkWgcojr4pT1id6NhKUGiq5DqWnxIJIMayUWJgBVlnHtA6Yttity1pu0P
ukc0EVoRyMSlKVCMwcmOgdqY3Nu85ywzJg+hyrJW61uVD8jX/2B7X2XkYGYzXis+
7h8d8nWBpLCRiFLm1YyMI/veBjFZ9okPb/0J9YLTLhTXeaFbpA7h+SLVblMJvhAF
rShLqVD5BE5ct+DdALPJMs6/7F4Y96HoNXP+9Z+kKQzXLlVJuTbn7ZmvSCQiEtZk
mHNHhXuATVjUMMUQdL/w6bukoZ/sCCkOossiA8kCy6TNwYkLdLT67IefkZwEuIXl
QF2q2+Be5PvdOCpZ3oBhba4chYt19piNY4phLlmLeYwidfh7cA3WSvPZ6+GP+ZC6
cCEGosjejGxFURpHPy12FXrPVw17gXOnPETAiu+2jAXQCDwhQXp9MUANHcyAevFo
Jq3FsOebVcbU+LxTVDN8k+C3Z77roQW0mgFLLk8jxf0dqSvrZmMLmIEATnCE9cTa
3wKPKFxGa7++q9qQYrH900rprZfndM1SOFfT5LPjLLeMruFrP/TY6PpXqmfc/p8e
erhq+ya80n+KM55DRCMYPyQZ92YfxOWdrkBoBu+jBQXy2rlCXP50wPPRx7Y8J5kp
TXSZ9tRh/CrylkMGtFNMtxSi8/lo6PcRNaaS2/VAfRVVUms1TD+2FWsXCpQVNrnq
KotFJ9aLrQliev53DG+XKMD9ep9LAoymDI+VkFBgQjUkENWlVutrHf7e0LkBS3a+
/f6gQfm5ILiymUDaNWVdYyt+x2E2M2AQQIeF2raRipsA8aATJ0xmLRx10y807WSc
YLu9lXHBRgHCZ8NRAutDYUUphyx5LwtQ2q/aWEmAtFbBVmLXqSUaooo14y5nFxlr
er5aSG7TcM2N7F4gnwjHBfpGaQYMAcfDmwcBnCtwfzmPi9wBwUGzhICoH5/96b/j
13q8q2iZCUwqSCtYHIYNZNfHlO+zLOHzAscQAzFHA0TIeVcMhW5zugyIpE+RJCmG
iUQt4+bhOPIUtpFsa0B9GN6lwzk9E1xCAOeQY1H9NuLEqbYZQ8pufZi1w6IW0u3s
7Nohc9h4UudFq5Fh4/Gh3kbuq33bcZu9Az3POAiKxrkqkvPhb2cnRwN+/fbFAiLh
6TkMD98tQPndI/4oIq+r8wYnqFAYwSq05nA4XnfnBDfWcwd30EWr5HKvpjitQRDD
XX7ZtyTVsvER5kNNITRKsxaHexqNd6LJUmUF8ERTjxIYV7GRuzJi7RhCerMNMP9U
JoW7ra59S8q0g/M5wIULt96GVkKQKeUIDZ0LqVUVSjhMfOn7yq+wv/w6GEdZhwhP
r5VcAeKbh+HyvUTeiVRfGSB6PucN702ES7LIsfEDgJZCDJlBy5rpUcGOOipWzb/q
Rz0+Fw7lTXFfwPDjkJHFlsV+r3XpwKac2Uj3MFr/TIWu5Kyw0RVMqtTYWoTn/l77
OSsL+IEi+B3AsNdgwbU9ZajCHVYiVLFU42lbYDTJOKPKqIGuWpXofC1KaqT4ecRG
uCB37C8py7JaHmtbz065JltU0gCMts3WII2ew/BniTW/fDblPmQGaixjkEAFLvMW
9LZbK30CfHsFIN7OgqZiuJcFp4qqNEsJbC9r5p82XOn3euzhjLkafkayHXqaLWkQ
i/5Fb1skR8x7tCHN59Emhx8Y//4jDvZijS9ZRd1/ff65F2GLBIfsnS8zq0B1fzCH
DECAzseE3GRsj3jFWcunOzF4UcrtHThy7SHAvzhtuOLnUMB4KNGvKmZiVmdKR4se
5+icZ+8bVqPEUAzpBomSkjcobwhBhEVbs3f2WKwf4p0MD2FYK25vLfW366HMZ9xQ
SzUMyPIedLd1PWDDNafUW4pmr+AjwGeoxhTPxdSHPeVf2AUXg0JpwHhHDCOSF/j7
3iIAXhLFhc0stoAIRWzF4D1rix9g9U0AKIMASvOPCu3aTZ0pq8BlSa6lYpc0QfkJ
H/sQmhgCxj52OOdffMIQnIRwfZgVtqY7J/MQNkbENCwZYCZlfazXexr0uqbBayAI
j/3S/Cm6pcwvw8fjofFCzsvjG3wrl1wl7KJwXK/6WisrxvLzwc2BzhlaRSfKfssk
eN8vbAULz8FOGeGHaT5vOWqqNbM1Gd5XARnBq93ze9srlHHz+NBp10hOe7V9DQEB
jG5JPREE2wLdm8tizYRyoBrx6e3iVRhhjA7FsxVVCmH4O976UAvicYWVJm79OKN5
tOomNWbpJ7cUFM+LVnYz2plRc5sfD2jqU54m9IM47aSONhnN+6CtW6FsJjzwZGHJ
G+cWOHF9r2Abx+4JxmHYXukW35p60pm5mesgH6VaR9DHQ6emghkYgz4pTcV4TIIQ
JL/V6HDjeY4Tp1S5SxMrs+qu5TfNrEjgpfUn2GWv8msjWcEKqPrGKeWcYbuI/tIk
g81CnjTBEgeRh8rrlYvj1/vMOoDEEUcIBxRRxAtt2oi7vsGkLo2S6pA4s0XOYp75
Ef8e0JOUo8NXdUapbIBZY4nki8rHcF1CznaZzQnf5l1uWehd6ZXH7zyE12UcxNMj
FD/qmo1izZc92SmizeGwfOEy06umETZpN9Ea4/ypWimsh8xfVBSoSr5tS8UlQVgj
huAjflUW6UIbOkFFY+UFFlSNqZge851DurkiYIblwmqaam9x4ycRQdZa9dXBy6aa
L3KHRcgCD1tF+guxZV9/vQ0/eEdyMRl6e5tS6qBGq3VHOL88nahyblDQa2X76tZx
WUYvCsI/TXbIav+c33E+vgVHQlC3NAKBRXeJAjd4j1l/lJlCnuIn+2fJqhpoTKPd
qtJPICHIWjEJG5mPq+SYIlzh4jTR/ZEeSDpm3UAEPuRTNOpsMDow2nTPacR91TDE
77SDasJZkC/B4NMdws+FtwNjT2Z50kWYde7hHSQT7Eoq7LySuo0Whir65LHpx4fq
FSE4zJRFLpyTtKOvUlBnUG1hzj3KrBwbvI+jME332qPQOkRhhwruwKNvpYjfZuxt
qKodIUtrd4mqO7EPxVTbGBtiMh63anqOM6s1InxOVUtX+22MHbnCnBZA7dOc8iRZ
rH8qbTaXK7BCqtsI5fIzQ0OO3jULz1r1WvPMnkf8ebEhp742b5TEXHJ2IaFEHKJQ
/QvK2SlextETi3+6C18CmE0f1eENTt6/c6MlP+M1c6cWsnU+Uikx2ju8n9JLu1i8
hN+I8GvFDP7EtXgBLTUOHB/8jHFVPfNG9dVoArFaRD4fZE+8gDuyFhodxTIYK9zG
nBMIWFG8ukNSrCqLij2v+vSxm2ov3CVXvF5BHAUKjl9kdrFX+j/X4CEMPf6Qx/lp
lozVm4sIVD+q/VqEaNvfNggmKrFJOBRcoec1p50BbpxTtcCBnQFPSqACLuiOc97d
sDyELACxBfBSw/+p1uxaV52APQN8ySSbLqwGHCDFe8ySiVKBZFY5Ia2RwJ5UR8EU
F6K0U43FYKD/zFkPEGqCrkOi26GHcSaiuHq8U08gSWDKb3sNcWH+Aq3v0PeIBv91
/MNYVfo7O5AgKZwi7RYe6bujoTHR5luXs6WnNhH5ZdZoUaYEFkpXD+aqMjEEuSUU
EJNVBsV/0wR6AFIAtSJwnSqKFtug5562pl8CHKL1yzXEdPnB1xiPV5fQpHa4So26
ZLfZB6bHNo1cd7xy83uJ9c8YZmNEUzcIOLQGJE66dsdCN+apB4Znq2XXIMq6dUbq
P6dSCv1/TGkmc1ja5ms/MkCdeIR1Q1E4zIDDhZqRYNH03XBg8H6+nfjUgcuQ2oNm
eSIFa1ClPARZckvFM/9V0uhZjh2WtnZbMUmtPM5h9uZfK9aAjmP9BUyVcBCMpKxH
y4nGj9V+CNVX+PIyl7QYvZuHhtpQAdHOt+qFKgFS1VQV9E69hEf7s5lIW7jNa+uD
AsO+SBZfWrugcm3i2lPiUECEYj/D/5qd5kgEExzz59YQqdCtKYDe+yfMocZ9NkPH
LPQN5WhgV86Q6lsnAvWtawYmGylu0MGNY7pg9xS4VRnNcQ7bbn+J+j3LOxXMPAI+
Y+UWHPvw8qUHTO14LaB/Xw6UX4qFAA1mh5GL7lL3gO49oZZmku9L1pORFR7KZNoV
jhxvNh21DGbbjBhj8/aeuKdyMfWLHailmrJ24Op6CER05kJaGDyQyHjuZ93iNcd+
JvbaO2Q47wPT7Ntw78EZkg5EMeorVRpxJLtF3/Hp5Hkefv5Kk61OqbPETkmn9Esp
Q4x1C/7A5Nn5yv08lrvD+7/xbEi5VgqbpnxgJaYkP3Tzacn/pIVtfcYIX8+BKNql
uc9b3d7T5K+CLa9i4Cw8vvuTMYCFRLDiKqyG4ZqJASBUqWK7DpXpkG5XuKZijkmm
4WzvuL1aBfw+MpX57MA3un0BxYUG55DA6U3Pra1OwTB7B9l/n3mldHO1sZX48A+z
pQ1sj5hHQumABQHIJdKAhqwwYCDz7tbJnfc1WH8mTZhPi6HBoAlOvEKKto8r61Fl
XWi1n1hzy4hWZVG8+WPJyAkuwydObFNM+G7M0EVPOTZRDFZ0AbX67MzCHDWxWT9q
l9qBnUzWhIe9cz8NRMaq5YBmkydHNKtmvbwF2nsSMpul3pXsIkp4PUDqcp2a6CIa
bMw2iYxn8xJZ1VJuiXb0ophUlQchGa8h+rk8QbCLejEoK4F0eKqCjGD0H2AsmnLA
uyCF4XF5qURauXRaf98fqr109ttgKxgcP3YpZ+nTW3n4G1sdecwkYrE/gb+ujRxz
IPqXW3Awfqda5662rc14oc1PlL4JPnkRzrv44gADjf5BLsv8xu6pxPlTeAov7GIQ
KCujFZIEDi30kKkd6JX6P6xZ8iPcTkO1xgT8Oy2xQgyFJK+02AD8sCtEGCKCBc7k
NqVdmWPoa8XDZ3RwWJLeQgnv0JYQQYZBn3GcG1Gxe1aW9npkO2ylF8Aa7M6EiI7S
hEqog6lXyE4j5Uu4wHqinGr/ORmeIGD3FC2oBf7b8HmAP9DrXmwNGV7m5qBXrTUX
wrkZSxenadkQrZ5RRW6HJZsD18KF7uazXfJ8ANsMEmhUOf4357opzcGzlcltjKQM
Zrn6x8Uvzp/XiMTzmzMnZ9sF+zO0PRVgMjhSya90pJP4/13OKKeIE2+5MNJixldC
KgfHRq96yVjQDfHFwx8lg2UaWdPELg8WevK4Ha85UMuYYHXVQjwlNVTF/OFv/Exz
ZIXjIJVsJjXe1WdbRPfIrI942TTgXmD4nqzp+KgouvGYWkx7+DONJ2HWw8FyVt5U
C0eHfbFa0Zzz3vxUlJtrPImxii9xJPal4+VWmMMBPN6XzfqUpv0+utg4lcvq/mqj
ql5Jww67yM2ybhi91Ss5pxVHKQCecFtM6bvDOydm32KiTmFvh7vfFhvejLI1rk5e
m6U2LyxSi3WKAolYjzgPCMdASk8FsVp45eJZmKr6Q05IQpkMj6jCjAwq+NKmtcgO
A6msflI6uTKYMr/aYMy1x2RuT0QPGk/Snk56VzfeFBDY3dieJUTFA7jHP3h5Vf1E
tz3hdEJAxq2tg4v6nGiTVHfSshpGZ2TpWIu0HEIh/rWIlzsf/8elXPikF++ic6Qc
nSgPmUduwHfi8gReXTH6dn3RiYfdceIO5EsLPqXANd4DnTxQfXptRPjRBqFpOngV
+JnnbcPPyQ/x3HgzT5co/v6uzuBLzu7qZNEPrgoo2yrK5Al5dkaNWEerUHk0kJ8z
dnlrKeDyVCTBQW3ifwNIgj8cqZRB6C5EBMeUYJKTgznwAs9qGH7ciXz4CcSLytKu
aPZ8DG4YryvVCBRfNYHjj0TsZoFLiV/gQfj6Clpt1sWW6Cdj01e2Q5CGouKOiCPm
lYFyx8F1TBh4OuCpn8sBMK8kDWyPAcgG9yhpPRavzwnuhlC3rebnrsu07kKAUhnr
0q9SCoHGCv3JKEvrfc/bQf4zWS/8hm71ZYU/cusRFpk6F+KNr6ISQv0AcSvSygmn
YlHr/ecx0fxyNUMSbyRN9imRLtYvkrr73Zop+MsXLVcbjix2DtzaY+WSLVSGCfFt
zawNaEZnEHteaWw/RuQyr4WXb8RG2qiyWDa0tFtLUs+uHCRqGe7xSjuyBXHv7TG2
oOC05ZGMtVQTR9nxuhRsdtJa5dYAVh0bRQdWjeHOC7PUJmIskQhbCpv3mUmUHn1Z
5/y9SGwN7Avc9AyPb3oRLht6B4CrxSz6Bk2SojM27hehmYbHn54YWvj+3TywLWRp
lcUa6c5MhO/cJYznJIP0bEoERZChJxCVsVME6i4Ky22Vy43r/jKFincJcO1yaAwx
kDxv2EyKuUKurN6gUCY8hrQ8LcrfLQSW/h91KoUEZ11EhtqnhQMqGXBGLtk+K7z5
yFXerzrjkwR2nR/BBh78zXbaHhxWpVRAzCz5QjLKb24xL/R/qSrCRKzJtWTYQh77
Q4a4Ex/GFtBOyg6cSySUySAoDQfWfvkpBy/w8PDJtpXOlymSUDjNXhHnCjSqRc0N
Yely+7Z+tZZjAK+SH3iTo9dpCamXgH4pApuJcSW7QvE7MqEslCMU2JKzXxGzOPeS
PKqVSYGWIRRDvVpwa6L/aItNOafZ3qw5x24JXMKntUZcjC5Pv+63KmHvQkSXzT3+
+OsSkN+zbxYJWVM3inqwjeDKdU9OiZOvgVP/hzTfmVTt2mG2CXE4ljNf8dseB7s9
k8HyGLh25P/efFdTnlKZVcqR95WDCtAyf+yaTDKEZLyYiFWsUqbjy7pv9viFNFSH
wg4/CAml/Fv1n2Iq4/Gx3/quOE360LHswtHm9OC3yOum/xz8rDwHI2txHCirAz1q
xWMlhuEWRqXhEbr1kUqUR0HLhWippremr8GuEtlXEJjyJJQqlwuBRkqskohR93J5
t8tgyBC3iYjtv7kr76PoVr9QT9No7xeMlJQwv0YT3wBKtCpYncwx2Bg5x2bO89nc
6KJ2wKA+Qona0MDgwBw42c7uv2fLqyi8OGbG5xW1fBg54kvySIWT9xWAJOAHWVxg
/j82lN5wrs18shVWeP6m+ihfGUFYKnHyeHL1kDmewelhUIymyhLbH9L6x5NUaJHo
VJkthGc7IT/EWur4RZrHbdJo+dZf9s26t38uF3/TLu3vFaw4+u2lVsEojDz1sPgj
XDjR3aZ5R/O168FNAE6hhqk/Jmfcjh3VSKFwdOnMMZ2zrnvk5OE/tDKCiPcml1PH
wLkGUeKVtrXbf7EvOCYW9hsiz/M/cq0L9loV4HpgfRPVSQsxutiT4xqT+XRuqNmU
US4JqBExbZSeMK/DSujSqOicihGxBWRoeAu9izSrrYhEuMDlcl7XXp0Tq0hlUI+J
0z/uOhx0tXQ9x5X/GWx4MGZDUAtFEtdE54h3i2x9sO7QMaM7zmqOzB+MiesHo6S9
eVPEvFLfmJJVyvZBvtdBgqsvbqkqMnUcGgHJxqfbaCW8DqT7Jm797tlwMARNouvT
xv9ceH/FapvCjopdz0ahsg45oy/DxbJaIfsQ4ucTj5mGt+RfAPW+ADdleUGwOgXA
1B97NFYskPtAXLETu2u9q5UkPneNt40Fha42zbLZGdjLW2gkLOnFX4SvzWwA+hzQ
MsbWa8UEuSDnKt2QAMFmE23vJA3PMe+FgRYYDndPjhueH6mRVSo9dPAasEqo4SLh
FlXJ2rsZSnLCHJRXtdjre79FM0GiirxgyKLPxLXDEheBkKoVdSMVjwuEucDORINc
Y4csOU83Z5dJ8eg9EgrU0Cdxln0XTg6JESv8QyLrqM1QbDQmvjkQ/02Mk8h/IRB6
JZLrnHRoILKoDB/r2FSInqP/A6j2WVWiiaA3es+e5V2YMAeJoJ81una2zgnZ79HJ
CzHrl7t3STDK6v1EdlNuzjRWukDOdMIP5pH3BoQZgygOcv4icm3eaB5Pn3kFer0N
61B3IerQYVXPFl8pdYsGXpAcZqBAxzjV47UDwdnrGHIe1EUKp3Foohpv8ALjqzST
Kkh28+S2uD+Vj5Xq6dOpj4w39YewpK6k/DPXUv+6pEx8g3GCA5u7XNVr1Zg4xHTA
zGZLnwQ38JX6PZLRsqwy0gFnFErbjRBLhslexYi70BFHxT+boBBNrvEBNkcQ4rhw
QFFYYTPiPBrwtSy3c36+RPrLmLvN2WBW0WB6s6NxgcIKBd80jekXEVLzXIyzvprZ
ptbA3yMLTZTvYxZgbvYuOPIRqJ0TKfZMp5oNjUOoj2yymSADBUwsyqZuLXIeNDsL
1ajYvX5GlAYX+kQ/yOUN/DMcfr9wHy8HcHHGlJbnZxjhZ8JJs4FFotqlJjrqAPRc
BnmdM5545hHmIJ5RVvb/GC7eXdG4ee27TfOAhPEQc1NMl5Nk39goGuKYNM8HhiuV
kLr13u4q7uA/iK5JIZHPsd7UJJBeOPIWAAptvysDJnlfhlxU4XYC5BLrY+X/S8rg
vZD8k+JenMrlHtJ/5Cw2K9iDENAXMfSirIL3i2PDLVC6WjRldmdg9107hiegJruu
7tIpJ1UMYf6KuvVuJsLZCZfPP/8Asilfk0yQKQH6kZRejQwJ80jpN+KxKQJUC1Um
US0McNWZdRv7cOckvV86E0LjVmhW/2XME2fKAhA5OJhtiWktReSArestUBcJ8ObE
mR27wsv14yF6l4g11rI94cZjP5/TCRzHeLiK+/hIfKieMdVQxAQeFOtKe7HKc3nG
xNVFf84ZR0z+Pbm+bcY24j9trY3EgkRpqZfYwk28YRJJ98X/FCID5JS6O8LVroEi
oapaZZQW+mjBTU6xC/CQJ8j3pWFjB2hlDcs7CgXmfQb7T2Bw46guY9HsvZ88mSkd
eyc4bHcRS+IFmEg0tdfvSSa8fNgwK7WeH8wLKkt59o4sCN0vMmTXVsxulHKMrP5H
2B9TxVwblXt+O7SkZxKAV6YXhcvZN/LiCkmfxrKpyJ2yyrqP+9MJs/AHebypFXVA
3lmILpOH2axsj0FC9mBCp8TaK8F0DUeKUsR4U+gY6th8pqhJ0P675snBVog8bjc5
1qUYEf3KUhWxzaueq6hn7kAx0bnZzdfWTn3PZg9lOyyla5Xe+aYg3Goy+4QMLkRB
uyFgcl1KJWZOYHgZr+33G4wUjxMG/pNaeFxivMYAt6ehOGvGVkBto4WHD6l6/GDg
fVk2b4cfgZJvsgGtHX/KZHm+/5GRKGDopqm6S9aopv4qVNMgOxIsmNGwDFH2QcjH
vRhMmlKsCxAXlteMQ7tgQ0NS/erSFZAeAF0izMtlTTV1ELTTOcn6gbIMFO2kkJDQ
AZ153ru18do422moJ+Atn1phcQj+ePE5h9zaWW/CPX2Ta8nLr8utez5fFw/NWFGT
/Z+SVGpOMho33kqh5mZfWri2w8agnG6T1hUZE3LSNkDRW0r3FUZsvn8vTO/e0E/j
PShpffnfA/gOM8DCMVBqpgGHJzGzC6UIIVg6syGlOXZFsrL0cwyaYCcxAWW40XrB
9i2PfYt3nNInjxad1dkmq5Sac71N1h+Xz2P6JBWoNb3irJUh/zkGvR/MzvZhMpDZ
DvxoSIIQXrqrX/r0sQQmkrwQsk/xIe/Aw6sxLCsRCg/1n8S6US9/IEBJAkDxG4Yr
x2vhrPkMJtWBikNHfkGj7/FCwdcKjr49ZhFnF8YKtU0WPl45pIh701kpxiT2KscR
/1GMpjbsdwhA49NCUljlwAohwAe/V2NxwQ7/sMsq1RDWcG+insJtSEWG0c9r8i/0
G+KTPZZWWNrT0drgqrqfFu30m5lgCp1CQ0fVJUWZn58C+cA0MflnHVr7BBaag2d6
9LwPREOxtRsVZlZV/mDB9MWln8udkeaLndo71KmZzkajK8lhLegWN98AYaq2FwMv
+Ulb7gYVrz6aNhNnSzwpLHOMs3k9AWq5dCS0vneRvgJ6sFwbZ0Z6wzcCwTSCOU6/
Q4q4z4950U4iYKDTCfp3srlAB4irhxyT2K4NocxlY5X4ZflB7E3/juRc92bm1N23
6cbQRvQK7lo7W3cwZ1C+dEWoj9/u6t5vZCwNSb7CZ5zlJYz7da3dlcN/pVAFh2R4
jDX28Hg4IfVdQNP3eLV0zto01Wn4Ev6trJcLxwFeMPDuDxbMj1I4EidNzOCve3Cn
9IwIqT783uVu66kNDBXml+HyFhyEyXEqAqjI2WqlEj8P94Jc7d46syARoLF53JbD
Vq2zMCAops/zpoqnpdKrVV5wCrsOfaaxt4I8k320/4BBk2blsHRnwrovK+t8ucYG
HmY8dQkRUn/oVCXA2vub5VeMBv9oAfvFg2rHwAfQ1vVWXOKexImEYAvhx1ys5nx6
MTMRDYrG187H+Ljaww5RAtsL439K0a/heUND2LXfBXJKdKlHrKwgb9Ek+F2A3Bb9
dFymKN48eTsH2Mp3z8bLykOiAFrW3tH0TweeN7/lfRgJzlyRbN469+L1UFirETlp
Y13s1XNbySogBJzG2ZOLa5U9SgUGiG3gTeMjJYvwVPFFeP5AMR5BpCARkAXN7nKJ
sd1DSRanaXsuKnZ0/BP7jKN4kq0a82kHBmlBBl9K3IX3cT52ystRqEpRBanSRAW5
dKV+fWZurHJGb8RBFVpyw5a5+QuEtPDu9SPTcVBfqqXLc3sRxlcCO0a2U4RQFy3U
lN7ozxr/v1Fqj3N3FNLG14MxKMkQamfbNGUTcqKLRY8YrV9QSg9JczC3vsQR7cwi
sa35ALo6C89MRCAlfWhig1LLaRlAPoSRNuOcjAaDKR3b/Iu3vV3oDDRSi4Y6oW4P
bViOuemiq4BNdcTqrMz5oI2DXl0k9+SqF75F7sMow+Yq5EqgNieESxx6XCME1vIv
CmWxb3+M98XE9bvwcLWPrEZ0LCs0SSEk36yFfpp3NdGkv1dAeaPCNBb9X7wJ+pAe
1WprA6lv5K/xAjPUxn9N7T7S9YGSvCql6z73dl2UdUeJjkMYnXutbZWnF2eXGytH
MaD+jsAJfVFRTLovPow9PiGzQXTInnnePSr1K4RVyySfpwfVv7bFgtcItvgmZNvN
wjRAqXpjd7Gs9W2frxM9KGNEjLEyCvKa5/53wkE0v0u4qLymxkBe+Aj4Ur2rJpp1
LzJFXluzjRiIu8i7qvsuEY2ankMbTW07wO8qV9SPCOOBIpjNsnqxTWdmyCglnbqm
nfhvuEEviEK3UcfNfHAvQCs1kq/cVJbi5mKKN3gRAfVWvupTTVEfQYmAW8NT1njX
OEycCXBEL4vm/7s6fIT0PgJYYm0Qsik/+DGcYtxFy6S6QHpVwZydK4cSIXuupwiz
kGNTSzi1JTHBt/tzYRkMMcflUZIWcF2UjWmdHcF96Ge9Sz5YaRS/GSqIDcod1CMs
Ss+2coU6HSUUyzrBcWNmj1TUsHyoRqVTLMmXNK6yyhJ8OpZhAg+2jxbFiQ7q9rbY
3RksLlfmu5ofbLOydqSKU3VD5UldbRpH8OaKN/6S4CH0b7zWlXueg9zvLTvLNeAN
lSCphLbI5ttFBUQtpeOjT/9UFVTNct45HTy8yXP/4TYbcb9K/lL3BLPX0maTQntu
J2gh+nFcCs+uRTN+XnYnC9+yaCGldBKoV6Pgc3thNMR1t0+Pspkk8mrU93qqsSxt
MxJz/SLcTEuxUkpDxH5uiIhFM0Opbvf9FMr9MouYtBIjeVp0wwptQ6hGIvTjl2lv
G4mPNG6pw2m8y1Wf6JBCT7WoKLwjwVJAqr9VuS1Q2jyzwC6DwpKIKvUwtfZ4/78L
uc/F//mW5R+rH05IPpCezLRG7Q9hCxQaAbkFnbW9ftgNQV/jnJ0VvN0Fjpr9gaPT
wrKbb411++HikqM/RRAqRdzwSyd6zYe/lFphlbtqb7fDwjtZ1z77g4ioX8O3L9bw
KHqRapvKEBJoLl1gfpqUSeeymo6YBqxLpXmjnZgg0f/LrVLruhGWHGTY8uQ69ZHz
/PdRB8DKUINMnBRW1x0uW6IKRuikqf3/5mGtVS1dw4V0APgxLugxiJI3Uau24Dvb
r3xl2L6QCo+3r/j1qNC9iMdWbMefM9i65ykcdhGQ8MDFfjlLWUtjHWdJ5d8B7QWi
XXsy767rMz8E025gaeJUp9zrHg1Gsm+ldNLAe1xBv4IamzpWOKxt4xJAN+2ZMLcm
6Cl1iqBlWHUBi9I+BOP60NDPbUmBSRMd7hz10vgH/vV9kv12+s0GUZh0OH2mLa8P
jcr0M8O9XSH5mK+lfw8uwFkTl/+yT4Krr55h68rKmukKFqwNwyEqrzQpZZlXt/W0
d7Ga+KP9M181FbBxI1oG22vSJHjim1Z3x/tiTgi42rOmX9USDSL+o5CVb5+NZ3kO
6KdEVQfNeZKJyzub1Ohm9NZnqUP9DdKKVf0v3KRa9Fi1dIGoZVH1dWY+dwV5/O1B
VtGbne4rY37oy6izkM5RF0r9wxrNJwi/0ODjaFmPyCKF4lOu4iCBaQLnMDvDjXCW
Zu2u6SbVkukupmVuGa2NBRmetm6T66yk8vESFHa/C9a/LP8CQgFVoESTWufFpivg
EGD8txqvmVYCeprqXQW0B6v+OXXVat3Y4fKd+yoa0cxNY64b69pfhj7cUDxtzCH+
p24ubosqMIR4In+SEeDsOKaAHrtvXWbxWTA2gBG6Cu85RXOR2iegmSvUbde1W3bY
irQSKQVgk7Gi4I6VWuld2kB89xIGBntsD9/Z4pixrcvNWLZSrPZtG8MDzXoZ+wN+
azCNc1W7jTE9i1HN4TfpXNG+UhnfrG9n6Tx3r4BZeVHyi/voboQ8danCgsLwf2E/
du40uQSqDATrq0oGh2ksDsXtCFhqksAmpUCSTVtqMcYa6EBUJjfgt2k5n5I+K4tn
KF6HXuU7rVnfhkgCUPRhlcTRgylplITXOVis144Ji0SSOjBCk+KPUTY6q/ABNC7Y
0+cYsl/udt3vWvz9lFMyZcwSjrru/6sCG3yhtk29bGC4VD7svIKqpZ3K7VorX6ux
+0TMWhhLqjYZ62i0X3HPPDm3ngI4uKXa/dEVgCSCMiKsa0tsONcV7dhL7HakX3Ii
Ikzx+EIZerLO5eAQrwekBlZFbHJwsjWHFuKsztIZ5eJGgHNIkrdlaKOdvLdYUz/F
PTiXx6DZuOjFnAQEzb5QSmvCZWYtO53gZvIWeTKdM5ZsNqztHurMC38D2veUGvz0
MBIGRA2XeCKHK+6VK3AcFBDfmAYY+9cw8ttRz2j89pjgb4yAgK476mhEIw3xwBtX
KwW+VKVr5AE482ZkahtmIa4Tpavv/g5q91EF9e7XYq7T5vwRAC/3zNUzO4njgWim
thvstF9xUp8SatMtkgtToS2Bs95DdpwakkBIlra5vgLFKTQKqYu+C9fRt++iqn2H
PcNJic5+3UUoL6VHrJQP65Q+FpqWnxVvSPYqONWu9LMc2JIuN4tr3S8wNQwbnmlh
N9uIXP4nKQOXjD4vUrjeLIHYkLsqkTJwpaHaPmut8arqCAR1aHimeg/cR/30ZNr1
TJqLw0R/WbHyG/951Cwnf2GQ3AGlVmYDmVzn9IAgNGJF7tK4qJ4xeRTnt0kzpyUt
rbbluh+ek8NKUJVMnbX5EWosDiqb5NwShk5zN9eUESvj2GU6X7YwwVVu3uiy0xnP
dgr8wqWO5KWoKKIvBRu9ThQc2MUuKgzSq+hyTUbiwecvFPIA1nDJ5OCWNhSCqhqX
87an2DNI21X7SSC7sACKqMouZEm/m7bCsIB+Q8Hh+VpSVOGW1drQLhyJDGDz1b7P
e6UtfUubHQwid1z5s9x0UgHE+is7zSl/S8IaOD1IvvW5s0zSZ7V8Oiol/9PYb8tx
2gOXFra5K/wsvPw1BZe/RlYrv+hEXGIb7yKgesY+q8JFmcQwhY7I1dGuMZSy+3vU
d3N6Rr3YwYlKD4af9nqvYv7QNhRk6j2l3DuhB7DLJOEWZ9zfTGSojHRdUIHawcL6
YbEjDa4j7lj4SCyU412Tm56JQX75etqTGaDz8fs0cVZNkziR0b8wcbyeMwbFxTZs
DyGKEBWJWLN4aiYQvCY77Cyk0nNoXY96AA3yT7/ZpO5Y6I1eHhnjpwbEMCu7HHyJ
Zn68pRpklsI+Got5vBRYTi+0ekxe9DsL1yb3MKCOjwKxqDyP7nC1FNFApZn3rmvs
BqBeYnQxhPQ3otwjFYHBV8OTITrGsWsuKUNzIx94gUpJ/Nz7rAAsbpcLCA8N9gmG
QWuHOsH0AjB5RyS8XsFg4VDEtJ2Z56lUKqUXvGoantqwyef1mF3aSFiNyimX9tVw
FYGjxSigOoUdMqvDU5qUcCEPl2bBaQk4VDqxwnTgT/GimmxN7iCt1Gw3KJ87EpBq
Xqeoh1Rnm9JD87Zw6XTQ3v682aAk/SEPkCC89JJ9YgdMYts4oT83nGq3ibS3h8aN
iS+o/qRI43wfJRJkG2ag0gvPsihyadumW22IDynivmjqJOIFxqTCAWsZ6VSDwMHA
bCO1tef8T9zVfXwitBy8w6+v1MQYGzXFGa4wMmnhhUddeyOQWAsSKUvJJ5+Pv8Ib
bVZloJVskQjqkPDdLb0wq+vcVdmlKoBlLlqbyAaBE54jCNJpkn7Jcr75C7GYz637
CUwq1VNTIK690XV1Y3278NHUmAgNvEWQ3zPEm6EeX7Tw+oThoLh1S5hlaVVFGF5H
YcedXESPnwuXfu76SGfHDuS4Iu+VrQZnJ3180vFHf1FqMT0w23Kivr6Ims3CidRG
Idk8b0AAxbyKJATOQXoWCdU/YhiITGUAuP56fdnnG5uzMFWncTfxK8uIOMa9tun/
eyAuskneLsLi1tY1Nv+DQCOm8xdBc/9FD5bVitYPz3dWYP0s52tDeT7BL9nGTFkr
JmLGnGCFXdEXTCYbNO0uHsijC4kypXl2ma5GvT93i7NT1oz5khJ1x//jAA1ai4QZ
K8F1TLjE5b0xXRWPdUJjLdJ2ro+3b51ydjkSiNe9hY2lSC1ffg2VDFtk86UyQCxn
ZogObVgcpUeScT0HFKe/SspyxL+ssjqCRq7q/YtzLGQgZZ4LwFc48eWp+hnJ/D72
E1jFNFB6dVrOfDnpsuQIsjuWnkVkYNuKazEAO++l2I75MCslW3gTi/ru39WB2Hzx
M9ijNLsUKvTUk5i1AU3T2he3T3PIJ0OPCh3EI84hsHAc0F75PUXbld9cNOKK0gt0
yLeug9W1S+N5lxpjlaqcdtSBj4Hqn9ZN9E2SIuJfOUz7c5JLCfmdQNM9jnPc8OJ0
tBBoid/IFePuLokw0hGXkTf9gAH2wIVHxwCnaH19qHWG/+W4UKe+UewlKyRp81vQ
pWkd0LwnqIinRdoKNytWL4SYfodPeNw41HdRYai6WCoYEwlsMpwx+qIkMyQbmoj5
IT3ZCKw6EVVJiAEutObF1Xei0VkaZRd+LkSn5tliLh6tslpkCIpv8rx7fiVJS5Gd
2Rv9blcdYYqbTMGn6p4Wi1JhAnphOyTlUu9ezsallgiyqYz93MPdbwZhNXtPOzaY
agIW3JJYZJitRl17OjVxBK+e0MMRlwv8PJ8tfmaec180tqU1MxKU1UPrKCInvjE+
SnChBOzbn0G/tZoEqEMnSHGNhGXN2NRt/LaE6jc1XEhkNabN/GoslumlwzoE6rrW
PIlud7a1THSiIihBtT/wEcvsu5uAfARw7xC4vA2xJ/HWhva9F+v3CwRU7MO4YLwQ
B9pVIx4S/PajFquzDHwqgQTZJnWWyK9bZjPgdcDOBx/9VhpxkZA6bHmNUSbd9q0w
kXvKDoQHaTpjPdEbGMD1XFd5EQ5XZnnkJVdjBHdUGQueqi4d9fDm7oRckqgasqlt
g2ojcoGRk9tS5vDXZ0mO2EDCZroTbFOQweXNcjT/fUhffKLoP6J6uITRQcNyaoek
85WVPVBm332NNcweCKEeZd1wU9MVN+4hEPvyShvx3j4Su4JK3VkScEgKApiLJ4ih
5xyP98k8IT9HTnWk0JAWnNb/PpX2UhtpAA8LFn02oCyDIpfLagEfr54XuRTpLPjn
Bs60r92aU2J+sW8seiML5cJlAtJ4Ypz+OKlxIkLaRup0SEP+7ogLON62pcJz3qsa
jJapa95zwy9aPxsFLu15d+CUcYuW9jfwYVn8SRxlnmzfiV/EWcyK/hdP95jhNr4O
mTGk4ZlH/hhp994JXLReBOTKLJJZP6/kk2SSVhvvKCx+5d3N796Bu+QmugQNWc7o
6grfnLdCCvf59u62axZaZBMmjQLTV6+OajCuu8ipD0DnELw2NNQMVDOaNOXrZCzK
RkdPILCYkURbTV0laSiwe4eoGlvmbh2W00VFseo3Puhb74JfIfQcudhDi23f5X2p
8xfJJ639mM1Yk02W5jx0o2T8LP6rSyaLG5sR034bRAaQOej7acW9BiqMoxO97lXF
KFU2Zxq4skkRdPdL9uJWaWb5Nm01fXz86v/w/KhAxZ0lmdlnFIhC1VQZGXpnFVvi
VHU3Usdr9IXBSacjvhHAaC0qCiKz6buxcq9ytkPyO+xX/m1/Olm5J8F7+kXD3cjx
R+ZfoAcj0ysOhibwWyYsXyauP7eEpXvXc8oDn6PScFos8qxwphGWtKD4dC3yeYR6
JeEWjPnLMKE+bDM8thDJxF6y1ofcYwpchKt25NaRvcML4LmljfTapjelew5MweT5
X57odCZPCW/FOGcfiD8mhFhUyCEr7T/pry+1KAOoFO+YM0oTHYrCsp89WSTuOfsj
zFXuNwwlKVH5mATYkyO8CVI+e24dTfXGy8ubyX7kKJO9BgwKR2gFi1WsYAoVjPJ3
oFAdzs/Vpcbi4Ae9NptlCSyoKCMEH30DuC5FkVPYouYdhMaXGMln+tI3Dsd67p40
AIKFyZlo6uybN5k8DhXcOnARDjBgBL2TK0IwSUdirSEWlQupiWnWkG+B+sswBxNz
Yy86LL6rGgZs9p+7d4bGED9eXrYTyMHP2rC0QJUHkN5eBMFbhYHbVOQy4jEUZ+V1
vh3VeQ6VWYmiOuVob50i/JhBdAPzXcFS1hu66ojp5PLiUOgCJaAdenGofZuG7ZSe
2H8ZK2XDvtg6kyKprnW63AqALVnClz+JoM+cKdsG/y+5VQZJGhD8fHu7kUamE3kG
4DDcFJaEwX1iviNKc7euorxK+ra2J0aSgz3jaMGhBM5pLE2I6x6u3EU3b/6xfMVy
sy/WD3Ewwvhzqpw7XjNHlezcHf+L1PEj99WHaXp0h2JnfZmHnVW6jFdObT1ydMVC
JXSg7uIthhsidJ+eeWYahzVKaoFgISZPrlE3XlVcTFZJ6AgU/vk0DdNoJiwJBenS
/eoJkVk/tPHtVs/AAiCjN1MgOlDaGLlBNFkVE7d0VrYmGyR35Adw6JomhcYPiDHd
syQO+iFfsvvqZDUgaRj2tdBydU6y4769uQwqNXhBVqezv9mWZG0/o83dJ5tHlq7Z
MVIJNUH7zN8KX3j2x7wdK9ljvGShvIv2k9Weba9Xtfi96zpoy8YHlUrbWkEu5TJ+
2DUc2j356gGC67RM7wCikTDAcS/rEtslNrU2AYuRDSO9kTfTCAMysCB+2K9sKORQ
iVcT0Ss5ct3LIODmGYyvklvlV1c69CdJBLfsCQxlvixtM2vBAF1+RvsDT89Y0pw7
LlFk+cMxN2+QiYlYMWehtvb3Io9MQVT6kwGMopq9vX8ByPQr22gp/AOZwgddnLzX
Fe+sq2vPlYHsRn1SB7aXLiGoPa29qek9R2AN7oIZUl8702kfs2+kmGjPhZWQ877o
m5EV6BIh5QW+ewmzLV/INO8qujOl2FDv1jUSwV73a7ms/Z6haTEX636MeXSwn1m+
0YomdfHgSpQpuMJcp5J8WyA1t44rS2uTa3qmvUgJlIaaHpmQdNE7/hbKsYLzZZOq
JUjk4U//g1c8ROEL5IbJ3oHXptU7haGN2YwCoHH4GJjB782rLpS1KmLODkX6mi4W
IcxnDAED4byzH8YPl9C2Hv98PzCKq4xHtNnYnxYdInxoeZGeprEAdT0OoVdjvs/6
rAJLg8BuVQSJ9e8s7jn+FEMLCbyTTVzxukJBlpiCMHGMm672DQZDtKXMxfYIdejp
Y6C539RiRT+MgFmvj1nWvYYl/yuOn/h5HyL5VVrTkKVjtrQekKM6K0SozycrgUR2
Y74++soaKBstkH7cCwwk153Fmb5IDU8HywRdvNXkLpIWnA+HJxt8kpnPdo5LHjGU
pF1m9xR8oJOUGM5m61aaHoWHoJChvi3z+KZNH0ljaNkONvRFT15HoDDbgTX0Ra/O
pO2Qat7Qp6fD7zKy2uWwq8+9bvrqu8XtVnq7Fr8dY1VKB1w1OHyWYP1In5KkCF30
HWq498SZHATeztjIT2W0581+VtXX1Qujd8ouPLaS3zhiPBq/gCJ0kVBfSvVneBh3
8FXt6RBSOBtTmwf8Sn698gKL5unUBcmaIsMG3heRVHulLz6pO/c0TCbaAzy0C0gt
81Y261OlO3yaIvGwR1yaK8hEj55ih/Sgai/Z5e/gjOZm85Z1PfljEU3IbXM6kC4/
IUTS++IjsA2GLjCoO5fj02nTLrBRqEtnA/iNvQGaWnDw9YjYrcRGBRTELQWITwC1
UZvX8Hl8VL25pwVy2HG+WcAnNp4HitKPfRZlVjewsscSYUYZlwXOShsqvOwMr0O4
iTvlvBQlxJGERHqReMqmejHTjW6MmKdLp090yX/Axq2FW38Q4SYgQQOBNWzR0LQt
lpRYm2WZOPBC57VWUmiJXW8jKZE5uUi/NQRaAoKQk4489CqGsZUUaJ7HosvA0ggM
1NYEB6sAsULnwRqd+VgzmstU2LEJNxvjJ0xESNpPVZY4to1+KxJTXBEVXE8aVugX
yXrJCBEc2e0BqmBV1VhBIYM65DjiOclXATaTPEtHbskkv3upJvq+ehZxwPVDZjiu
BDHDOetNbPHwBEfcTNsY+VqhX8f+Mx1R5GlaytJh/g3Wa1khdOnZBGlHrkWx4QFC
j+RokcyMdt9eY6t7PWVAiPSdk9FE+k0a9f0JFnJ6yUUcBnZRQBi8qGWHZnudCr7Z
0BA7GwZr2Qt+rHGLcro4uWavuiYeJGcq0sne34FSIN/+lVwVLtUa2YohTSnxZas9
pP0Mw/++/TTdL8XbqGsCbf/S1j592nQ9pKa51IgFdVB/f9VlUznu1GjpER4xTPrD
RolyyJCIadYaR8F8ysIMVTZxb7DRkeTlJES8sOEMI85/Fta/uJmt/EnrFJEu/ZDz
Z1LIVihB1ZHKFoOL/sRqgLtBizMDYYapeC7IMom5P6dNDVIX9Cfyybvkli2PCYrN
JNaZLFYnRTUTBXN+fRoz4mUnmfjsVbAlh9sktf0pEasOoaABNboOC1E52/2tH0Gb
vAK6C43mrN529tne9XP9015urVE7aHs9ENX5l2WbuZdIAZBe2okSJsHu+nYRBjga
Fu9ziQcRruAZ7TuHUSH3ttDuvk2ielh/+gQ0xq677HWe73sMNSFqc0Cpqp64jtpj
OArksK1+jdk5Fw1i1OkDBqOBHOPHWOi4GdelrOJ814i61aLKSlYeF7i0x8izBbWj
zJrZndSuwO+z5HWQFPEQtjYeFsEe8cFYBgxMVze4v8jtJeDWP3WoZBOfXMmCPWTq
Eg3mkA61WTa6hP3T+u+me5E/60bhHtAcHsqBa0yWJd+s6UaaUGTdL3h0I81JRtEK
JzKWffHuSYiS6yB6L+HPibbtsG37ExqMugge52FF4Qs50iT9Po9c/Q+gVbowvzgx
MxvFcPLVrg7UI44TKE12YUGJd8j9Au+0VgrOMTp+Jg5lMN+mL43Sxo8P8aULkVWo
MYKoqbKE3QR12bIG0oxUp4+wLQwOM06ecFfomMbFZJ0odiMHRBM0FZ9xOVzIUG4K
WwrfOsBu0rQNfIoS2UFHqWknf5bHX14HshIym4+mt+if4T0ngJNzKzL1FxPq9CgJ
lYzWJb0LoK98lTuSFdFrp/GLYGRLEyD4Kr7aLS1KQbsodyzsuJwtrYQbUn5Cyms1
HymWYM25odGv5nGZP+flRP1IwEMq8AsJOxLMAzVv8MGTGLz+mWfdZf6QH1gLX1iK
pZNBX2dCGpMk+52NIKqH6Q8LCev3jkKkfT1FVMEuSaxPg3wlOQHVHpFjjvzzF7iR
aV+Yms6WQBpaRL7/yzSvKz3P3mz/+hKhEfWczJibbrRcNqDE+0mGUenuNrBfEwk4
2ssy3+B0lqDPc+NIaf6iCSLEx8q9cCE3M4X74wsNfxEOd94wTPGeHXJ4Oc/zIctJ
tNH24QcSPFyAV3rRZFRkW7AEKFHhwequza1ILx8TMX4maXGy1i1Ff9HpWLkWtnh9
4fDiP6s+Ez4pYNmoqt0Y4QMVuwDdfRDPlFByuFfvmJaVZm+BarhZHE4iTenTa6CA
ombRX7bloDbiy/4hNWqpFc6b8QCtIstgwOxW/Wvfr8N14bf5AZJItagFze3H2mte
rNcCf4MHAxHlyQ8/hmy8PrkYAGA13CZWKndVOcLJgkqKkPxKCRO4jm6ADGq2Sr7h
yjwGp9msw5pUlZTpa1yq83jIjiTxF+oW148NJ4fmthUX47+0kSQJa4ibDVa8GcTn
ntoQunwaRXOjWHf3odkHIEzvCrveYJ+0BYlNGXWzUaGv3cGJucIn2wFN1Vz4W9Oj
PbTsTMjyHeh71l0UsDDWsmtskyyjcx/EDND04O20scoizoX2HE+M+/yW/o2ATp5m
0fNguaGnuP29woDfQlnSCUJqm8LWGF16uR97AAoqxu/OBbGyUJv27YvcWuYz5pUu
+qqriZBP3R2YLcNntfHEqITlakd2ccd0IgBo9ZDmmt7Z6s3ofm0Uf/kXWYZpUb2c
ziGE5xd3HnMRoRwBElmmxEIV5/6lafmg2QgoURQ/VukVph7zuZWxi2O4I+pW84M0
3kLxUTK83BPqgy+ffELrB/fYQV1tzl9SECSMN9vxfQOAq/9GMNaldZDYXL2hxXzV
xRytzRggj3k8qfa3XmnUpf/ZtZ3l1s4Da4gbGXdoIDkjQceRyRtK5HPvZfldn1/o
4dTUGqCwQHvNgdmj7VEdi1iSd52e9+ht1l7GhvAHMrcsl3xMOTYA+g+E9cbG/1MC
RJbGk5xX00juKSR3wYZxpf5Vn2G0MuMqYRKlDGd5iNg7kU6m8H0PZNBfOeOt94BP
lwNF0ouZCn+Ku+tE880uDTBXy0Tu15FvqIgvNCVY/Huj0e66JSfu++o6EJ512rtP
jVi5rkSgBL2aNUeiUQ2d9MejpR4hV7Eq+mBea3U65oMcjzW1dz/20oth/F1kMsCS
0rivkskbe+znEbAH8s/5yUFchhrkncWGMvUIh9R1wgTdXwYQQ6vFDwRVyrQwiwxa
PCawH6mlZrq2r4pAMvsgOShkLeMxu5noes4Q301qyMUAEwbPLmH73Fr/CJJyZN2E
nY2WCTHAO4da/FRwNmYF7fH36zUYFCTo5etz3zGVcZQ3aiT2smZaFsqktQsOzVTf
39bQc6A+pNzOPy5zBQapX3bsIdow8VpCU7p2hc0a8bNyqfrEAGvL3cCdqSCQf8+3
33Nwr/eujQZ6zTlZCDOs2lXkF0zJnVA1XOHXb3xJ/cuk38ZZwbd6FAqHrJTYoIEB
jKgIZ3z43ymvuEQjzz1rf/YwI8GpITtGcDcCLx6J5+HiCothpevphnOCvvc/3uTP
+Ff9Gkh5jwqgAWTzrTRrJbehuBgnqhPtoSPKi+YitORanL4/jQ0dfQGx8B9hyzi6
OOp6v85q5kTZaLVS9Wz1mQhax6xDdzBQlJWPuqDegCcrg04q5/WVpvfk08BalzxD
tfhwlUtaGlQ/oFd4WDA2t3/pZnb32MWuvGMyXtSe4HBuYEZluP6HwnFwCrYQODjU
c0EtW8kivY0AQhKnDMU0bOmPe7tF0btl2Z1DDCXMR2dy9gE7pRuJzICPvee11hO1
CWf81emGen5Z0+YxarZPjhYnFCYm/SICw2smNzZYoq1sWpfK4LlQeXyaj6wlrfDr
C+AT4NArPpIwEm+zS9svjMbZkkIO0Iv7RDguuAIx0Wig3w9jZMVSfEzjoCaJwyUc
LQb/M7oYCZqJG1DZItF/L0QvSowYVxqEdb9PvjcsKzMX3UdPSmMVpcRn+FUbrbep
TCSRZxYuQZjS/OsLH82WMQujLAul10THWIbXi5+kXwsybE3dOpnEjCyVz5bJ+W7q
iWB3wwAN3URwYFt48B1NkseDkbBL2xN2hLxWKTq1XiTRLIW+a/+x60VPbMEdpCaV
GFB20b2SkmQcfmkhf2YsNOUJbxpCY4UcuMVg7e54+JIx3uJTbh/w/8lOwkGVHEjz
mlMvvcSoF+l1yq7GICc9l+Q9VrmV6sEQp2UsLDSkp/MooZ85KWlW3uN995dDFKAr
AX7Bo4WrTt1jLLQNK1wI+40szwIzQf8DSjQ30sE8+YAiPCnf72JnAVwaDIbPXRZC
h7YKwqAEaRgmqE/p3GfgOIsAXyoMr9q2dzZ9i/M4WQjy/cEa9M3XNA+Lcnn3K745
UUTj4Lj5owshsSd6ofKq4oY278/2M5k+ZIwzbtPsYzfzpt24E4XWcuszfH1I9dyc
zzNfXZyoxVXic4u1l4HpFvAGAdedoOUayGDkKgNFKW78q3Hn0T11t3LTP8QbfOlb
+ZjEBUqG8xbwTrFmFDA0PQycx5hNUIknVDLNqVcjQMuVYkCx9lp1PK/RxEZ3HpvC
1n1kdOeNSAIT6kRD8B2zfTU51DoWvpuTUXSvtZaZEPWz3CLYst/Dw8Fhn3jzOO9k
OT1yyXUNmnbbk17z4CS6BbM3wKPA6FIKn/h9Iwr9uvjcbr1AgBY/8OHDOLEhyJcN
tNjAAwXCfzR3YHiTKfRtCB81fTrSUSf478v4ubtX8ORltbXACbHcB64ksN8Dn6Bs
6IU1PFTr64dnRWCInJjHeCtrgXaLXIpaZW5p23Cvm7+9+Jj0mALWlUoqewDV7Cep
lWi3z67F+hTCxgf0MvdcuUd70CZUYrJ0hOlTQZrwpE+tWo5Dft2j0gEKqcIy6gM+
z/gGRrS9r2L8/UkCVElzeqHMHLDw/0rRepQTv0oD9ZumInrnwuhxh0y14LECWQGK
ndigrNBSr3E0pyEAQH4SiL6JGCVuorVRhftScSYzi3EdZnllmBk/Dn8ThRhVmbqE
2KJpC+5DdWF/TpZDyYNuV6UloIGIQR/x1fh26sittHgTu4/k2m99QG1eZSMJLcpM
sUq81nQo//mMkZhfxNCx8tgE8mRZIKB8G1FKmouiK2ZgLiuP0h1bariUjKbfdL3h
TBmwMlfv2c8j14MecmLowN0cIZVSaq7w2gUI4eIBOJK6HvwqvPQ8ZifBrfGkgTmz
P/CQqPlWtkoJ8km/dKhvQe76uAx69U6xdy5kAtptYxo/+pXhezdGMFRlu+Xonzhj
UGy704bUDcND54OGDzfiF6y+IdxniPAuv28O7P0BDgNZlJscmrVBrYCiBmQgZHjo
gaewh1zbXFDfcrf+YcfEtTpKvHgvNHDBt7grGYpzc8zicAcUV54KxbpIvZNpFhiT
bjtthfutOMoHBEUi877jJ1PVVpQG9W/OCUIVA7UmltXw+VbqjCWb1qOqgMFJ3rCF
vWfZQk6KHHjSc3Mu/db4r/kc6lZddpML+i3WlbNWTNL3Qnh2kVeMHIjL16c1eVaB
CFlYdB7MnTtOoLTbCn29xVFOy3v6JgVeB7tBgm7Nv7PsVzXUxH/5gyXMfhPqFuwU
u8PHF3nEee7rscAJStwuSEue2kZlXLNl+cUVUMzo0CPhZ92NEomN1Br/jMJQHar9
wFXBw2jfjVCGNMRbYWXQZaVdYnQmDZN4D3if81/v+W/gSg4LY5WjYvq9trrn7c4B
bGPn7LuM7OfvqZvgSgSIVOhkDo3ForyE86B1tMdI3vL6IyjENZUFrLLwZRHK6Y7+
qUlt24aQTW9iAmgm4vIiznvLH7iwLnRYUM5eCwB2VVhazB1e9IsTBPZHVzcTUx+9
S/sYrDEVcnw7tlvIwYR89NtU4+BGXlKhVrAQP2Ds1780N9tc5nq0FV/+iW/PoZKE
GGZbfrD2JeggiQP3tYdFlraZU9Zvc0jKccjo0AQh7ctR5Xl5L8IAlev5LoULQqlz
pLFt7nJKpR9XnwEBtcgHwbjzisXYxz6ywerMjbRJYK+EeyfsrwdcqtT0SIqnns8S
lhq3cduhYj5Z0r6/0P5WHOA8y4W/C9KY0E5C6P3rYlFtAjwYpw74PGBZy51oVgbT
4CZsHS1xbA/HxlFYmiUOE8yyYOxvc9NELIp8Yg3QH76qvR9GRRACRb5ZHycUTCJp
l5J5DEVvvlLJD6QV00HQQBRcSFuHPSOMUjqIo7aECl9gMp3xZGHrRE1HTwPTBFaJ
FrbaYa3r0lasib65QiRAV7V3r69XO/rk344r3Doz6VhUBnClLMNWw6X8kOz22fXH
3y5xfHdbth1V/No5LOxzkJ0JzKCjaWGNMCsE9cE02h0WGIMoUF8VI22YComquN4a
wR5xU9UTka4ZRWCYG12v1NoM2mJH35olYI5rKeDrVoxg9er6ef7kD0MzcurCMnEZ
s29njegdCUGskdS3WL4xjaGY+L2YCkK+mdqDzVg+shWt4e9jW4ozlafgtgpJ4Mlo
+tTalKbQzum7jpg2qHxeO+4XruLhgkt35loxKJVzv0POTWpx5XJ0KXATBKqxEUeG
KIfJnNj6AEsUeOwy7uktk3Qz5JwFXBav8FcESHvGqejCAorMTlLUniySwuclVEmD
Plj7AJJ7p05Jg3FxHLRcAiztNbu4Rq9Gpglf1BCbrnyXbIlJthv0A0BctlKsnm+P
yebwm7LCt/IbOrIHGN82M9hirDcJQYFAnN15FCaYWa5db0Czvm3uSuPX8oNHoPrp
o+3ZK+HK37PjicmSQiLnDX0/dzRRi/OXKNHZjPuAZGyiESQag8PLitBiQ/cjhOgS
Lqa/4pO4RuXARPH8nNOMbrsZmYGIFXiG+9P+a8/jf987FTe1SMawhF/f2ZpTSThb
6Dt60ap8qmISL9M2zO4kgIvWtOo9V6V43Iqm9hy8+lSYUKMPw3O1A4Vrwd+rPF8c
ksZaxBqezY6L8/uOc221UAHNveVO301HKgv1aEPJPKYsV6jd8Ozk/jvQIwFYwbwZ
cZs6evkiNQjyTVIia0KWWhQOJU5Ekph6b1dfOHjPToI7st08RKgGfO+IQ31U62vs
/ZdAx+jYzf0wTTmhtp9DovhEwHI+KjndW07mbPeV/GrxCNfum2vY8CM4laLnNrec
8Oac9pOM0NH6y5QgC8EYtv24bH7krBAPVGzTI3lP/MhrItmAy/rvdxOctkW/N4KS
soLwJOzKA5aBJasPyHj3Y8cWbPP3JMMS027LE/dACDsQdGsEhWTd95KY0xOh+C4Z
pRiS1X9pEW4Ucebuk9Y8smJK4vUpw53g7oKuOIHYj5QliAmTB7/UY41wB6s3Jnf6
4dgIQf4gTq5Do9LZ9wLfCdsMBODxj2DwzkhcdpteLbjXY7pWXDUSmt1dLqEmTF/G
PIgWTYT/oDAjBxyxKKNgt9zQoxH3fKG7lSSR7wul6Ltz9S9BF38EwjHDHxp5Asoy
BRCThWOXwmmhqEsFGXOi1cEyHejV6GHNouXCpH9tiADamLL7iITVuMPM54i+Kp+f
FuaLeGNbnxCUIYvLjIG1Rv/DhUPZX5vun5bnVWoCiCkIAc4M+4f4LA67ySs58KgV
OXJjIm69MiwD3ri8ugU2CaDjuY7hTobbF90hobnBDP3/JuIAUC4MLDRpULRBHFXD
9SXmLRqKXYMoiKlnprLR8WFcLylWc9ySQftjgOOLYrXgP8jOCOGVfgRJw7d99kRC
gZhaHt/wClauN+2iWLpAejJnniqbK9bH+vL7pjSutPptW5qBUyYObj2U5JTKlXmM
cfaT94cJw1NZeUSmNtSoBiPrT4B3GEwkfzB7yyOq06J/940+ep16DoWhvZT7/nxL
B0NNVv5Tv/dOFq1kNnWnvWcKWMZQJxWNt7TtIr3kkeEW6Sv841PmOMwhcx9bTtJi
XkroIrJUVIC2cxazXCV7DEZWucJbfLnQYditwDBYu+w932y3JSD5AAYMUrUVLQnb
Yw4ZMl8/WrQX4kv2Jq3T2PtYkltIRjNgYCf9TLRgB+Rl/IcHISypgziyLGv0cNPo
Kjlg1TFA4FaoI2X6VOOFnCyVefMrdIUFQcSVuVwwN7WEzZPOH10Jvfdj0KUaTtUx
e8ze8Vn4+lQEZxIWTRLJMMRKL/E+6aG95vsQBkKSxJ7239/HQ03G5cNruuwlruoK
DtUZKNfUgJ5wV5YA/wDK8lF/Dx3/SP/+y0kQF/yGiyG5Cqg4laR0hCfGUDQVnbgm
KdjLNeCODWfte8U8s+WK96AnOMSZn8i35LGdhKjwC62eFSmxAs6vIVlDppJvkVZm
Gq/oNpQXuOnK/RneybeU5+An3Nzaf+WBVll7Gp87m5aGc8pO3fE93gV1kOpy+zq0
nd8QlBREIdHotoyGMi+H8QWmP9xQHv+URrKmivR7Gf12wQUaC0TP3fLuTdADoqvO
u70pS7ErxsGRd10AmPdm0j0zzeC8pt2efX6KQUNOoIGTPeX30f/XHLWypjGMhCZL
m4BINQs+nMZdoNUl75200vKYRChG4mJjZjpSQDCxlphRF90cTQk4SkumngXGI4zI
WEKhXxe/CIUpy3+h1WyVB+m1xDkceu5v7MOEg3JA/lwdB/y11Is0P5FNVZ+TejR4
HSrWrLj5ibNa1/ytMIxGPyrid9QvVbcCgsvZWgnU4+MXyjdeQlnyrn8YgO4e1KDx
7leIxeuCO6D7yariFXH7H/s5sxT/JjuxK6pfABwwP4saXdH4NPsk7fk6JaHPXJyM
IcPAnca9COtPC/9FMcQ3Kp3dciChDW93uGG16mP983/AXgfbnGNFaVAuy+WgCN3o
rmcPU6TmuVRc98dVt/ce2Yoj+BihNfTBHfn6OjNT/Y5PKuofKgtkT0iY3a3wz8Wx
3F0TWMMmJdWn67xv7vP8AEsC5T3iKvZjMeAtZrRHRYkFi5omIbEBvxfFTSegFGQd
sj9WpJFsqdSMkEu5id3ChQFJgVU3zWCkDqz4cUR1v6i/K8i1yS4TL4wAWyARBpdE
RdaxxZqfvhw+e12HWRPorFiSR0h8GaC2IrHl2VjTTvgv2sWBE3whoQOBwwn8pNH2
uAdzirXSHM+QQax3fQy9Za8AgZoxczW7TDmy7clbfTyzTPSk8+B1kbmqkTzhOO0o
D4NQQLcFpZQf6Ek+8thE0gFs/XKhq8elSTMTG6RUAy/V+gOzAK5nCJUp68FuEOU9
Lzi6cNNXjVjj8+fj9hg+qE+Rkkwnx9LaUdBOKUvS05fIRrAeuDi5xs3+We827N4/
XBWIn+7CLISdZJ1JJ8NPrnTZZH5s1ui5CSt3+KtJc1wbeKcDGaqXwvHC4Gh2rgEw
I+Qg53R+QujQd2HmhvDxc6cuS9yZUgkOc3x9gy2aZhV42ousHR3986QCR+TXSDQL
9gFgzhdW+7N2CDMuYwfFenQgsoaNrBVwhb28rpTWcB1qTM3vOn3oF07x0LqFMHAo
2BPTbpPEC2J1R+bDjtArdm23zUQGlNWUeSG9YjMa0KHFUbzZ67lIsLKjVsLY+ztz
sIulNndnV0COCGxMjSKiv1IcGTakB6eCJfJX4DoVoz4PKhFZPKQmUg+4XSog3vxr
Hp+z8eYfxa0U5i+hJxMeF/C7hBK4w/o8LiE4u6YhZvqlFH0IQaWkLisk2TpG5bRg
sbrd2+DLCCdkHV+zO0AVauvRxz/Gc8BfgTgm51wtXWfxtQjlqsutgd16S430akqi
6bO5vjC8t3MJH+IvP8NhpBXh0Qo2RST0OsutuUqht87Hun2bYeEaukBrPtWQaJS+
5wBhhdTo5GLwxG1whJ7CW1PmmvbZM/Wjb2VW7uKdRrS4QY6xU/92tU0LO+k1XYDk
TZ1nMq/gi8eGAQ5PqFGDvxvgWnWTPZ2NtAzpm4YUq2/rTXr3uf0+Y2kUTdKWXA67
KujEbb2jpwsUWN0H3FyJZOzl6jYVj8E6YhesmfhpKZvhNb5mjRYuWoE1GZjGSSc+
V6DZEraKR9ldHt4WTzPq9INRS/Hq2Z8ApFvcudSCZBzG2OPG4tWzCZN2SOk4lIPz
/VVHJrhLIpKxnq/ppH1AWISfeo/qVL/+uNJ2JlfCqjiZTIAg2YhPe8MuqXIMMxsV
JQOvEccl54i+fFBOTmmMnrA7Qc2DZry2gLHKsfJWPTNHtEKXwth2yhxPOceKqi+4
sCrQkeckdFJJfYVxhczeuqALfwkUA95zTPnY+PbFmuVCOk6E9ooZejBOYWVtrQHe
R3kK04aqYMwCUpWB0uV4nZ/WzuKT/RmH+PjQN+CG9taE0P7pu1N7DD7ZTtdekhVY
oID4EwG0uGo6INoBcdeqVljTkuCSrd+GGR0IdVPG6WtpVBg6RSQOLovj2m3Tg6a+
Uu/m9Wmv/rP2TJ0ljFCD/YDJW4L1CU8qVlyAGcf2Sb3krlkuCKpgRx//ldz3ZcDp
TB6ffXMvyRA8uFiibiiY9JVEaob3oTl35zLf7kV/wBTLfKcRcCfl2f5upGHXl6oy
OxJeHxmLpHK7ju41gBxD+As8bmOF1u3rIgBKj1ZjxdTgsYCAvljIxZbdv2afQWcS
OMcch0+D1D1aNyWY/Ek9wIKSOKoJYEFmSichf13h5Q3Ucth3x6ojLtIOnx00fY0Y
fji208eibN7b1flvNNqeVehPf7JvOTPQzUSG6Nz83wx1oTlR1mAldU7UmTCgjAez
Hm4087F7Z55c33/KQmy5Ls/eTcc34chvRBlO7r+kr/HiLa42hzEqDxMbPhltpjHD
wqZSo1RByUa+ehyW4MQYdS0z68+fUV9SjwLupVM6AT/aSOon2q5AeFF0jnHs+uD4
i/f1KathHCBF4CO8Axgfkw4GsQJwwB1PcXZeeIvBILUpL5VqNc4XLdePfikZFbHC
LppOr7uXsXTsJegc4GW+opKts7nw2dCHD9WRPboZ13ikKGIfGxUuguT8JHV/+uqh
bkJC5P7vh+4qN1jZ/tnpc2EgCqgEyCI9RalI2y2hl3TgKXIObEYsaKvMu6RjEa/9
fZejpMrW+5rmFuzPuvZbr7OjkEcY5LrbD1Uuj7OiNwGDSj8HVj3+4SX9Hyo4ykmi
CkC07TABLhH+FDuYNopu5U9gYXSRJv7UC2eFOwf/3dOtMHR8f2SNTUmTiZkkSfap
DtLU4KX/iAru2l0mBwXHoy9q81YJuDTgvbRgcbupIGi64ax9kyJLczPeETCtkjir
M9gq3aeUOTXbvbz2UiBeNxJbneibPcrs1+Qp9vprPar5VAykZ6k94ITxeuENWOEW
msPYQFMbNQMDASjDZmeOj4xG5Z7CoY876UIsRTSVnfKjy1jjO6FQiORZKcjLQ/Gp
xvkqW/5PssUQR5lM19wb9XR6hSDxJ327VrmT2t72ZvhFdDLr4crq31B8ohXPdAgX
kbRi2OVXm3GbYwUiDXLA3vSTHfbIx27WbwNqMgUfzpOYborwgz7LC2/soeK6AWhL
7oUqJEq2iTxS8uPR7a+JqFtJbLQ+azbO1EUTprpIj8C/PiI8lBwbGs1Y83PMg9qz
k2q3ZDls7GJ2A/ee6aZf6E3OtVz0Mi98Ps/L12wz1PKTZE8bz2fpq06hQdXglaqQ
DrjOUsFEf6G40f+mxyswFhc1d+7brBCntSKb72UPX1VM+1C78Tjec1PjyOn459iZ
GBTvJf/7qIehCwG3gMuv+SXwq2KjvVZNIIatH5RXUWNkRHy/Voa9QunCyZzyuG3E
oYxdnlMbU6HENnjUVhQAFd7HgE2wRIz/qWWx1znzXnZu0Tnwo3BaH38YCiEKfogf
WmJM09MG2mXs7E0Vei0cV+jiPVIvv0na3Np2WlqKYp6Y6eP1JQnUvEOGabNdNaIZ
5ZrbPEUwwwKSq3sAnBaLQVgydRc3kaUTCKV1DF7sWc0WkEYJx1nG0mSGkXIVe7oO
ES8jlKJZ2UCQ+7cEMkLY88Vv1Ij2ipdldDnM5Ex6KBijHx0flzUyt4PzCcjxnzj7
hgUCovuLjK/xCz/HhZlrr/ipt405K+LBaXOHxb+p4tjfFMQxRJlSDuPXZT4uGMjG
v8BEtNPpgR97T/sLCA4sbBi/N4NM27y3co/s9E3to/4d09193xjdUlbPXuYN3sbR
qvavjT9jxPPy3Duysc0FxDumfYVqqrcmj8ApXFXYZfA4E/YVHe49JBmn53k00fGS
sexMPYz4LEV5FvqcSlCALaKTC47gLwgAlM8jJV9PzB7PtSluRaHfZa1GglXhJzr9
VQoqc8cE0Q6amA3PQ9IXhOcfeD+YxMiOWvnsBqcrEZE3nUFhaoFkjmNGc3ONEfZ5
ESEg+KH7kT3tlCTVdPkcFOiNnj2t3l2+EgiHM8xmG2EYV8kTbZdMWczeLdjoSw/q
A5G0CoAYc1TWY4VH+Exk1yuc5IB0JQ9HVi2L8F32XrzhAi9hYaW6vWs8ldUzcDrb
oluq+wE++fN0oTaJQ2AW+Ktaz9Uqjwi1XcEr3VymakjTiKLoZecYIthzotIkKHyL
OscViRjICPhVvNKBEpUuSUYOZg3PYQfvolJ1XYkUc5U5jVnK7DvhfI9eozR+NkHJ
nh3iw9bJD6lYSgQr1v2tOvG4EKXUkLgvrPtLnIM8e1QYNpiDxK7D4VvbtUZKkYkm
GH+NFTdmC+bOXdoiR82LN8YCF3zRA1oHRKJlDykUF70W80U75e37gTgS0dCE21Ez
1s9w4JPdlyTf7lXwm174yitD8TDeXfcP1JwiUZT5dHf1Wm0/NthnBDAMVV7O+vpR
PF5TgOtxd1ap6jhBqNR/PmQJYIBUj1/Av+lKEp3CflQ1u8CpFCXgr5Efb2fY9lVW
pDOpVzVaqXtFgA1DM8ZNl0zsyJAuAgPQ3exMiJYV9ZEIEKf7w8oHsA5YIjG7RMFr
ExdFSb1fMS6vkvJySHnQ5Fm+vFXeEFRA33eiKb7uqyVjIk2dkQ7WF/5AGQDf7wlG
7C6HT07smcXUKqqWBvDmaIAQ0Ayqsq55iZNfP7hPn9aN0XJAYDioB9vJDni+IJnW
EZJHolri6Z8uH+LXuJdZEN3Fxw9Nouw4MmqzWCpXEebYRZWdQ9A3b6nvlYxVJe9q
d/9MokBfns7C2zAIzgXBU3aLiFU1v/DyZ13ReAb1bEQqAsLMPHNNUEzP5h/spdZT
ieBjpSSNxna29/Cu0AC0DrkN19BNpqA31UXh9k2snKUterljhIItRpZEATv9NeVG
zvlcrLdWyCbSq6R4X8+XLrcXgvDEh16aFBvWf4gj2Kv6rZuQ6ErOiCEG4xJvnQrd
kfFIZjvx4ZcPoR5SuQHEcU1OIbFDZA6bkM+mGSgWDf7AE7CogKU8l6h3HA99lRjw
+e14F7odyVXKxBIeZbE3jlnooGei6H+YPiWdwz4AADipEaaIWSMMwnsACxMHNGvQ
McUfs+9Y3LZUVJi2qzXmGaElhrXxOLaf8IQbI8Zs5GbYxveN9d7+jjOegPXg8gQT
rYtOmo30z3SLxbh402WhKQ0JC1i6e7Nl+gA2ddCYOSUhJd76JCH+tIMRhh1f3OOJ
sPB7ESWivmT1gbrwG45cnOSy50SwgALH1rxTXRVSfdxwWru0DlmcA47KnmcwHAfs
S+AywfVrYD61jm58qIayxrMmSBKAPY+cJofatKmmnwP5NnJlahjKO4DRXGr07Z0z
Jl5dtERseBSxyVq0k0r1juTBXayuAtISkubu3mNZ33Jb7x1neexEtM24IDLTKTvC
zZwEKu8ZkkFIvOjKaWGjebNRTi5HBxuatLI1huMmSHR9GqRo3WxNQ8YshZAJbwVS
48VJkccwI/Qebx6f6JFpvwH8SBCzgrAibWtj0mZbi8rO4wcAWHlPnrAmGvgubBbI
jYGNzW+24gZ3V0hgjji0K8vZ9ryyKxhLkVdUMLG8pIJzhLuCf/lJRobzNCr+7mNP
pAqMcKf37ckKRWJ3NPJZHty6sRlYxCZuZnpS+w2Z9yGiHX7AkXOZSkd3IUDDIZm9
Nf0g/zUUYqem8cBtny+bPUV3x6VPnXseYDNbHtLukV3iYIg6sZpIlwfNltXeY7nI
jK+1E0y9c+sHI0N0Od8Ieisi/Ye1QGniN7VL3cAvWOagZrNQBtSLEJnTVJTK4g9E
8l1fqNrilDAR8Rvr9VgMFKYTkFwRwo3JgGEipu6cX/jjnhFGb9430wWC09fzgLVs
SUyB7jtZh44Reyh7V1MI9tAvXKJSX/o0VR9EEAS4OSHhmVhTzTXZtodwCcgfMsqo
hKYW7x8B5Pzdtkykn1bI8UH4kDuosc9bblR23XVwgPJBJXjUI6NG8RWQtrsguBhr
767y3A5vm9V64JIBdWYP+C09xeiV/d8FTqWB2shrq3hmOHy6BPj6XcKjK1ODQWR/
MdEm7uW/tQBO1SOdUL8XfBoSqYlQRQywbD1NintSffbkmei80jg48zYj8WDkNMOn
R30FXOsJ56qYarGTr5nuj/ohoKTS6KNYWHI75Iy6d4fgSMo3ZtFI8TP0wufOXTpx
B+ovtkqz9E9xWWjE0tNbA6SrdBKMIvQCv9yBAcpfFpOO0AuVh9efUS0DkJRHUx0x
Rxnuq4N6TVR54eIPS8nua9H9gZGM9CpxD+gNpOGATEaJ9X64ypkr6MTUJBgaWkQn
VPUGVZwGN2zJY2X8qUnH59d8oSTHlUrI8JXykEafLq6FBiOxTou4tCWzym6nTs9g
G1H79Gy82K8TvLh51YQU/0Q8xF3ShQMTISpr0XIE4SalUwq31sqk5qNfH03MCcpc
BQa/3lQyOdMvmqIf7iYp08Byg6R7+B1J23zOr9Ml58uEveZylXjdA/d8mTz6jhfJ
3ysQ3QXrqWaXLKXWW7ZHr1zRcdGj709Kn3LDnXNn0YXYQ7J7y385OT1UZQ1/46MD
lUXGPj9UdLEzehXm7ckjYK20lq6vptw5QWHR0sNXI+HDm3ghvBuFAvqKikZTtuBJ
HRaOybUPTdfHv4+91RYTv4DPZWdyd1sA8hrqi2aYVeLV80AXXGNZi88lzqBK9+J8
2OWFqAK6HI7mHx/qYUNXeVX/tFHl2MzcnIKFku9BJYOmh2apRRJbD4WTCfKTUN3X
B8LjJBV4JGan4TSe2XTas5j1/OT5VN+HR2A2NTCCc6HwMx32y+265AlfVnBTyHkM
WYORQ4PSdrVzeoUiRvrgR7DLBoQ04OwlGqLMi6bsJhxE1zioxuNvUbBIHE8h6BV3
x1jpEIHML2GhsVFqFSU40nsIp64K8QOIVab2S5kQcvn0WcgHdLHxiUG37nycKtWY
ntQBz4JVruKPtaz7c9dHkA0ADod2LSkiRIbNnUxDcManlTgFQcs3S3LHxtLN3S5e
ui201ceocMh4x0lXVdfOTH7J33UOlqq+4et+7TYE2vdYMctXKNC0boOJsXrr/ps/
1L/qEkZSon7KrguwwEUReoyQQ2/huVZDlRoKDOU8AiYU0ZrBrp0med8e9D/UTu1L
FbtKaVI2Ldrv3ygrGz26nrzEFppt4vsPojOT1zqP/npfHkLyGK59Fcy6i6kvSIpz
YD2do4hTpt+zpusfZR7l8qNXw8QjzAosnfUtpKTEq+P1M3jLlRCFAwlO6GrtXskO
eyK/SlNOx5ZbiowoCqXcCLu6Zb0C7Rml2QFowGAG17fiCNNurU/rGEKi9B2T4oG0
MgcKTmxOmhC1dczunyOaAHhbJUSumS7jlxzDDVF4zBU5VKMRASKgLX0qxE2ZTxhb
6ltG/nG4jweA/esoVOPxVNH+BFmVJos3700ffhhkNXyLIltB1kP+VyjVbvXW3S9n
1zFR02pN9BKAcNM4gSyYi/SEd7Ruisucz8UldT1d2iK1/dk5ja2TA3aJGX0DRE6J
BG1h2XKBhCtamhKCcckiAhw+yfeZBSzZoagycHEfQguezrI4q3MMd7fMyqfi24hG
jhPIeDZvPjltFq+9vs2d5nAtZMwzy6xXrJwBQBPszxdVV2HiBuxL5e+/0kmwMNnJ
rFavYs1hx3chxC/PJ8pUtglAeq8aHcGBubae9hvNINNGRUySY0/ianXkBKgXFpOD
e6EeHz2u2Dw/uays9FIdw6Q557WYlTO1YE/Lx7FR+xMg16ytRGj2JXhHDUwQ2bF4
CD3Lx3jwhM/OD7VPBFIcpnXlOsPftezfzAhIgsmT850KB5zFkuIVeLv6Ceo3RSPL
+vFaFBgCepenIFASZ8AVC9iGYFX1/aQlayv8UUADxSNPeTnHD8xYY+ZefhpnXpmg
HF7bLtybxi+L/3RY7C9z53KI+8g0eQ1T1ZdZ18EE9S5gMyLS21X3TS4MpnG76eiM
h6MqhfSMHERZbGfotGFQYh0p3DYNnWJTqaWd17eJUDSdwP/7SDKe7DZk0ffy+GTc
7Vt7NrjKVxMXzaZP19V4g1/1nhXO2a0jb6gV89fUwbJW2lGecVgeoFePDddSNJIk
vHyhBVCLU6IWEv6MRJZ2M4XQJ/J+vldduGB8IJCfQApAd57gfWrdJI/7IjmHnQFB
vhFCvQO3iBUS6Vl5TTnwcPluqo6VOWKknGH5xk5DnQZtvoTmy4Y06JTTl7xKkuhg
EZxxRlpGEEiOsIXUcOYO+RUBsQJqDAO4wkLgfiQQkBekrsdh0J5whFo3li1O1cX0
BDRfi6t99CcfIO+aIPVsMsNpm5gipgb58hckSnmVnYdUz0wJG9QCEOY+9PqZXHGC
ffISNBeBsa5WjpMkvf8P1n+ySJHaeNTMDze2QrS2gb5Jk9n34zx8B38o7j4IamJS
lMvAnWbZ+2rUAnZa9gsaXr1X9Im2+UUwj3BY87YFScaPAdatEKByMPnJnB7ynJoS
I5vKYl5vIAtfsWuWROKZNnxdvBzb0V3BDGXaSy2k4Wp2T0tUtQU6zTzQJQDWQcL3
X6b89PgSP9QY3CKlKlhqyyCDrLsj+iRWHIQ0GDfQ0DuJWNylQ/5LVwtWBtPfzdZ6
nBYA1cu2F038gx5V911fFTM4Ektzbs8wCTAWJqC7vArcBr8dL+8oHIstlLNjaamW
5AncVM6KnXrMjraePszOTmK52ioKkE+z/wXWq6SVlgmvjwRygwrMKAezW2mbpG+t
T+IbOqDTG0PfKf0slMDKmujTdsegn4dtTOShV5BcHswmjOsqshRz4nZI5/42khJv
h79qKrFWlZy6uTG0YRuqzuKhTc44MbdnanNkpwSVMb9whgtQqjfnwsDWyUiMBb1o
QqgCxDfQfaZbUV9EJgrBeTnjCcdhxH1fc3+wXw2XNaCJajxGaawwxkjyVj9PSyp6
pIlKIwk/CVAWOpOpYrNvNnfD2PmltuejW3GZlDtZPLr+wwjEtiYnQRXwu9YDIxSR
578XCYBpQVpTCXlNqisrqKBgrAt/z7hEzASd44DoAQ56nSgvLfGWc3Jvt7wAjHGe
NUF2eFt2WWar2lInp9evqkNhyuVq2FNGZjQzzjgkhdN+pHS/Wb6BvfzIAlkdKUIu
7u42cDriA4zAwBIzWl5dxZn6ACbnIGYaUalwD0yAr8nWxPxJOGyd1fhVlVXB2ex3
HHqKzDuQNfm++alPDNRckI8soENqwe5W/mm3dbIOkDWx81D9mutY9ejLDMXeNSL+
LoSHEfz94nBkjYx+KcQ7X8dqRgXINk/oQcbY7V8BeEozd/8RfKXr6/S7qhRRii/9
hU0IA+u2w7ms9QPgPBV1cVQF9E9qMb7YREsDVzqEgmfoEqRGHfNFbLcRfOu7lnOE
k9E03mnwCHnW5mwkRQ0dpQ1NIW98eLyJ4tj87mK0evmNLKnVedFBFJktLpqqcK7w
PHc9QCKpSRhNBn7nKZr5pKl//8uTCbZJnjvVQp6afHTMsuU3k12It5C2Mt//DlxJ
VpAKh4ZrelrYMSCUxXBtceZBj/goRgtPh02DMkCXCTAovqCzU8NaZ0e6LrUNc3z2
k1+LT7u7nmE7JY0yFXdXv2nveU+Gv9KG5JM9r80Husa968x5nZTPO4pV3+Jb7He+
jZyIyIUWbVOSwyFlcE3qM7smvlbm2J4rhMPt/JgwhImVdKCeSbO08KMA72EQvUOy
3dLPOhVo4t14m0rBRjdzadcIY15X+gtgrVD/KqyMiqPt2chyY/qXQjb9gikpcHAW
/RN89QcElY8FwEFbphWHJjB9d9iwSFuzXK2FlOhWWIZOrRPCizp3ryFeBiizpCHv
dVqiM0N8wcOTzyCns/UZn8Wh7M5XeMshMnCysyUcaRJ8jolNKjlB72WaLyvJCFIU
VRdSX3t5zAP/JrudAx6sRzIBqr1Skpd4fQnTzbKDsB+WniR82EXktwxj0g037AkO
fXnTFAgRDOlS6wvHlCbQ9/6WFEcnqPLspkp9gjMOA+RFo9ROa+iKLHgBfUa3/26a
Dx59d/WsKX8PUPbjNFHGlmozAbH5J3ItoS47dukDkAzxyNWLzyV7wHh54C5TzZ2z
ogsvDtMVwGY8OZwEcEsp3OPt2BjDek/Xtoe1QEPj16G3J9o8XOTwIQb9w467ewse
FrkMhAUSRdmOdjXiYNNbUvlnwU3/VGgpRd4+Mb1ypj9TrAYUZ0B94GjOfEA/V3kj
tFQIAomjLWG+Q6vLzr4WRYXeTs5Yt/TGCsFN9AmQJqECssE3ULInivfL/n7WYclE
84OUb40z3P8G8FoNq9n2p6rxqcqA15H6xPSnDGkXleS92pJCLdBvaDGLFAkZtuWw
bDk2LrSIem8JDn2eJcGpJonKBRFuCDh5cOH+Lq0pY8fY6EZ1dkV8fwFStb7CcvRI
G4WpgNbBRhT4kUP1wc/cqK+1prnCKp75n8xhzhpBc9RyESdNNyOP3mSCbzBULN2Q
1uSvdPbhjmYfrBXm+1LCrRsO5e4tNoWqu3I27FDr1ezKxnamaXZKyzIxeUSVzogj
pOeJEVDOzYGt1n1f/KdKcoaFUSgCgMjT/FtdJiL0JSesqTz0Rt2YmgvPpUYUTYMQ
r6iNdBsc/Xss0ySyMqsheBL2ijTmlAW7/Kc/hvLb89OkBgFr05J5N7fy/rja02N4
SyObb+vCvw5sE2GFMvXPNrZT26pu349GrhrnoCUga4VpR8nacx5Vkj+RBtbLOxKX
CG2s747wGZK/r3YyIi0yu5l54j9Td8WfIeAQWLHqx6IMMoNUFyQoSR8DskLfA/wN
fByJsKuhJHydCD8jIp/YWz1KrfYxJKMFaLCO+rzKT23tRcIzOqnU62DqelTuu01Z
5juIpQcLqQxU+RGfbSUalXpEpjE2cdgwESipIyPocLng4BixgCVP7hNIPTOEET74
suO0jFJ+AZKAh1+TdtcQfwadcvlTw9tau8i9tra4iNQAxFjbffXY3q7o+G7tl0NQ
JPHB8Nqxx3Y0FV0qJNU23XlqhPjJuw+PkZ0QJ/SYqBZhGGP1r9Izuo7Mb+tGj66o
m/SGuTolwl3yJoDli8plv+/F9Pxhzt3xcIxpJcjDGoYvGA/OYF7MnNk9AwoUF2q8
iIrnM6gxG70s1WoetUn7m/K6VqTWYhyzABZSt1HW4RWZM2Ml6BEBsmPBiPDr57PL
0MHqEnk4OgbR6J2FFUcKPG0iQEWo1ZgEDIurcY+Ny+AwWkObAy/6KWg37Em56NTD
F6uAip0lCTMhUON/dry2mUv/exrE47zdONAj67PMrbp1vR8ayAxLG4xwWo5KTmUu
mgFY+250Ca3O8bNwlFnv0gqSd1cBkStBi7KrOTRnhKA2k7B441CTYVC58/AFY/0z
g9hc/S/4khFlpeeoFDibr0HgHl/2fTQhnyuLmC08FAChx+REZGx6BfqskwT5U4O9
JJ5C78tnbKWVG2BWOg14sHgEl/N+zstSnFh1mkG7Vgqpm2ki3Iq3q9g/c+To2mxb
loPH1sh6821zOKelBmnZ3PyrFgFszYJXsYS7Ddels5nYae7qbK4rhX+WcxHxUaDM
tZOcRlfsyJDDnOwo+M3jnAmwzCJERpErNfYybq2Lkj0KDwt+dhqVcJOw9yNwej8/
vPGjk2erR6KXsoWueP6Q88hYRHo4qOVzEB0H8Bht4JTDQyJCFZHcFyAzf+ArSWYl
7oLr9C2KbDQ7G2pGgfulbfkKYOvqJ3LI53E06LONjCxxLV/s1ccJKzF0zKfCG0qW
MvblbVb0Y93J/hitOB6VYqhap0xRkwHWYTvr/tgF4cNhnn2cqGJ2Lpg4SRwx1vkM
S7bKMpXgS0aQFDHJJ8ABFbB0pcJZUEnvAAvJh8UMo7C0ca5DA3IV+JA0M3rAqAge
u7glPj6Bz0mP0eUNguWQNokckZmIEqyJm7y8+QqEscnhzRmzE1XmXgHfnD0z4xTO
mlyjxrOAh1uaf7KTxwXxwzdASgh0EQhUTWGOAQ3iL8yEo/beqGsYhgnCuxl8w6DT
3KcQ09MuETBuFLuumzh6cRK4QVdxcLDvQgI2gKyCCEW80XQg6YbNNevDHHLfQzkk
/KEsxgYYCQ2/s8bkfGITlWkjFncl+GvHzdYRvSP69KVgztu2+wnsLJXG3VyRK6hK
05qDMOfm+C8to6UVSYNlnCNOGI3KwOFcqXzFglgKI3JnMkf4TwNrZwgYG2Dh5PoU
Tk2wcP01F3OOiCiHdjA5SmFz1AoFa24hdhJ43KRgJKiTuWDRbK/11SiHOzVX/FRX
3XkyiXff7mtzm+tnLrV2wrK7hqXI+2QXg4ZkHfSvkafYAx5DbvC9vZAWdvMKDPtw
XRTLmu9dClemQaVYiO+rk3JBGUDqsBpKr4510mpaefj9U2D9xCRUPf91DPOzbEk3
/JyYrHv3HK4LjcFgM4OK0DE1LQE0EG50GJKUwYP65ZQ3o/gS8eAPzY+Yi/heK0oa
m5zis/EdM8Xz2/70XSMfa99CG5oBrL2wzRJsr8AmeVgNXZwTW+oQuGWcvFLi7fWt
I+hGk789j8YRbxoUJK8pcx84JW064Mgt1gG4fySzbacjkP1/eFxzv4wW5o7bXwBk
nlNh/YlzW8rnpq00a8rblCF5EKStzqaj7AhE2etjIkfr7ETnZQdHOpInCdMVK+8r
ENaEf/B0U87eyESnEK1Ipjqm86W6LD1BwjR4CMjdup2pdcVGq80Lomybp1NDRboG
y0Nx959gzs89zHdhPQbsTa5s+VAxBWbVcrawVKhDhUh9luUVN8/Qyi9r8zA0CcqV
58Q2rlZkBJRMO+ssPnrSAMKePLrYMXNP42lLdvP1hVFMtqRahKPDbnYG+kYkbnAn
rbYQAMTrQkGKw5wlMJweDtH/PzITjYl2HUsni8vj+SdsMldVMwFQeA+mG0SA8yAR
Ja7snvOdAfQF7pdhdw5PSK5h9XPUy2yf86KX0zEENiQIRyqSwyj5IXiozjNSN944
Yuwfb54F25KUm3LfdS3wGQzSn2/XgeFayLEH/zLBdNMYTbU+MBqiMcUwoSw5zwkl
KEEeDOjPJbqR7rRDmU5IphLiZZRdgV8atRRG2fPcLmVCgLkcWAC4RG530vCvxehh
sgGRppz0L7uShdkrIslC9MBxEZkltlYYwuv+F9JTyo9UjpCGGD2c7n1Wyj9+A+Kb
LbeLDGtU2LD92rnoFQMddRRL1jyKjopiQSMGbx7GpBeZVpDxIee3m2YCMceehhR+
5AmKbQGTi0D9WL86/z17yw0XHQmui3iAlrjc/XCaiLZoUrar4ktkB4lNt3HWouD6
OS8eo6DRgrQgKNlDSIen9vGqXr85euTa1COhVFWPVa7WgYgkw+vlszYZIT9RmvIS
SYW9qhTIGNliXEgVoABcV0wsLEMP+/j7DaGeSd4qpa/sEKUXL0JikUXJDS0bmbee
zrhVUJbl/B5eG+yXnFnvhgXbGTqXSOrSNzIYP413zUd8C5m9EQ9aNLafzuZfWHkD
YkCqen+ZIt7j7u0EiAZ43xG9MT7jeX3pE/mtm+y3OWXbPk0mbLkLBliZAk+C0wb5
DzWyaaiyrayrf2tAXHVoeG1HdXMURsVN3ZWCuDUmuVkgzWhWKo6bf0HuYV5h4rSj
S/E1e3hERZ2WCbKKoTFhUZEdCOzgLR4tZ8e3h1YebJoNkEz1fXzc+EpkjF2bSbmt
6W2nfFsvriihwRGADpX7ZmBmbuUzeo6LwCOrY/MQ6wR6EWh7AmmzcRwc/9ioeZW6
krq7PGtEKS+fjCVfYRC2o8om9uHpEmiX9Ddzc6on9vdztZvk8pCA72i88NjOivsI
mCI9OGW7bxp5afI/7DBH3kjjo4UPc+5RY8sUXeehc+EFJW/HgVYstmaolcAJZhbD
mf8TqFky5fKuMfiNj5JDMPqgniq6rmK+78tYloZmW5WFHnNdjvJ1bAtIcxR6k2TS
H5LZeS+nIylEVc0qqh7OIeZaVuKVpkxcysga+qAGtk+XG4iuvb9URBi3dSYrROKx
/mE2WfdsdMQfVBSmDQhHb0BmYhN60AcSNZvDIvxWuAOt6Ae0FvW3qNCoH6yCcFsm
OrIH71ygafQZ9FmpaTrQQOsBWTu/uYzLqLgMPIxtNo6yH7slJuYl5ndDCKWzIv6W
KlaAR5DB4yYIr2N89HqwqWxR1VKbvDgBsu6h5kM/AqBZnvjhNJY5CaAD1p/xi94Z
Rw1XC0PZgzzYQg5WIWZo3dFCRm/bG2Fs2tpkN00cWpvxwFejSClFNzZiB0fz0w7c
lEvi3dc3J/dO1fzHq21SkdjJWWnASZdGgRFYNcxvmhBuBkt6KHKbYoTp68lb232y
Bc/+4FBR8wvhqAE0G62nE0pqdzInYB04E6H0Uv0RrrR7k5tPMsx2v5xJoZTcXRoJ
K5gOVbiMzt+Gjo/EuTFVSpF2sGzkcIKdCauiQFVpFnJRel9Mn1fghA1y9kgbo19Y
UYh+afYT8zduvgFbj7jwaH//0EhRYF1BSKmIVcZuUrdpp8aOoex75rHDpgdEp0vj
hHTra22DWrX5qzG5+IZfyGzmx++ql8nchDCnYQfGnL+b4QaAVdckwZXRMXPxFYOF
52Jyy1xFJ/ldHkv/ypR8WVq1KBhOvcc9vMJFqj++ZbAGZLumfjmP3z4qtft4SFqY
sO7LPTFWDtUyANuiay4f5wY38ArKKKG2gKqpj3kRpLbF81+vVGx+au3xeZAK/XsX
6yraYUk0XnRUyLanGOaNuWiHYH1ZpEDI5L+2FDHpDr1a0ZL2J370XVeP4jnvpy9F
ib1LWEmcpPcJtAWQcaWeU0jxOpdp1sJMBooChAWIHEJzOb9yiGHMHXw6ZdFTMhEt
4WM3VXB2Ny2UQYMoggboSbpEmb3rqOKhnfWM+WqvMslNnFEE7oe1jZFOx8fTr+oO
B94bZy0Woe6lDy8a2bIPsi20E2rVhKxDS/zdMP1kP53u6Qgr2gOBMR3Tjv1mQTXP
GM1xko6O8tgT171nbRzfqxdcS4ZLlYxY4I8+QhPVwvW31VuFgQ0pPvmdNNF636Sd
qmal5MkCxGnRkhVPD+bIM8LOOY9G3oj6m0NFANUitbkG9vX8coSeQz7V5diH/DbB
s74kI+FO/JXelFmSaHi38Kt/DbqVnKgCsytui5hZvjv4WM5o3QJ058+J4NxrPhEP
FWh59XwoB8f55OWFjEb0qOxa32r90ZYDcZzkHfu3jozE5Gx4DtF/RU8UY8rG8gx8
IyScP7oc6yngi+AiE9qPmZan/F/9VIQ62aoYG+6rtf7JDa1GyoV3R/3gcOYGfv6D
pKmxMid0h0P+aZ19fp1FkYU4ck88ojx+VMj5S/A3SEarC/Fp1wydFsaTC0HQplt/
b2gpuEQHRRHW085vCpviZCW+fbS7tMZQSWEB9ptQyR1Esro74dhRMWu8JLCoqcpj
inOW664rLVAgjRyUaFNxjrLQpY2Mb0Ozd6clz4+UB219BZiLxsqPnee8PHcpDEAP
WrC+YaLO2I2BWWrMbYG4DSDlK0AoG8OWTag+nUs12oGmBECRxJhzapHy1q3zRRj4
GlxfcYwElrudAQnQ/VXv5Wf/3ob4PFmgtGI4gh2y2ZQ69l9LWL4LWB0ON8bh8FSY
XKNntMZ1ii64xQPcJjAqRtc7fdUl5O3UzDAnvvsTQkHjNVQfhhMlzZtAbjjGwT3X
5qeC90IelManSYj8rbxu4kqvKYhVkFQZkHyykoJ1mdvn2tav+VXnBw6tBY8d5NFo
GXU4Is+Zrvs7EYt0X7wKcJHfc691gseo7gvlJF3MO2ZRmVnYifM6cHJTQ7HWOODF
zEgQsKY2le5Nxz76OxVGLCFEKzRRkkWhUOGVZKwx6lq2Bpc+Pcjn7V27lg5dFBBg
gLLEOWbZw/+JIEX6G11uAM9o4nCkRInZzGANHKJid4ICn7PUTcO+3X7DOKFrnJeu
s0vRiieutjTR4IYnxOHV1NImAD3faRIVHlBZ6Drl7/xlXjRd8QJCuGjAsz+GS++l
oceY4FBEs2+koDuKrRsH8L0rtUCidoNvQdFP5iSY/9En9zTtSgZv9NJm8szYN2Vl
K2jAQJEEkh8mjqbXbh1zKwJayBCSnyvwEp96HStoik7q68/GkHA+SUd2PQrSbTCr
7l0OOGlI15XIlTvaoAaA5lHQqthTIb62gY5gw731VPTXjYj0rgcjuJmfC97TQHDN
+P8sMWqmit0PZRbNpwscfvmElpoAvy2C2EVYUSnxEIRJglO16UtuSRO/EiTZSHVD
sR7x4MqyMjmVPeOsX/siEsD2vV/ZauLhACyh+yGCIXvDIb+tSJStM/G7y/8f2eKn
T8qPrYTtr9pjQcbzw2mblc71yzBglZJ9nB1e6eEbmVbdLAp4SM6cS4qIKLwBF612
aok9DXPj0WkCePnc5QSbsvIldtyEJUOgKE5DD6myLgni4XelFApeuZY0zy6kKRyY
8/2/Jo6F1dSM7iEeywtta+zzS399brkcsYvJAGeqr8+PmNSzsW1/SmaGY/wXWCct
TVoE9WJ5m0pV3LCXmqkpVfYwSz3yYQ09nSEOar8KFVO2nZ2zl1GVRINfXFDcLCyw
9c2ixxPvy/GeVLv/e+36elAVtKE2dA8OrG8oK+UZ6Xznzai+9S2lxuSwt2SJir2x
xfbyjKnIdE06vqgG4hZgPIG0IFXYGmKOppphR++GfyY8FXhGCaUs0S2ZHlc5NT77
VqDJf8wAqT2CSNNOVxsICZhlhGJCaCJBg+kOdztjCzLD99b/wPlQWLW3QvrWYzwh
LLsQUz8rPxH1PuYz6/XCvpLL216JOHaA0YCkCFWo5xj1soBM7Eye154LaepyU9dN
BVEa0XhMd+SPPoEhGOo5edYdUCq+5J+GloSxZNiVDOZ4QDgibme9BPpHTMb/H3Lp
25thKo8E/adW+5fywCnwR/5mTDP+Los729wHn7SE6vzc1QQ9npkNZgh+QmZr1pth
ibFTuG5pw9UxusrNYkhK/19QHORfoj+GVWFKw3G7n6SXFaFtax3pn/iVS0Dr8a/p
jNThnnK+Lk7LYzWV7VSI8IqToKImogxEmi0Ygd/bw1Dj9VGm6rzk3LOlHBvmhU/u
DXClKHyeDi4EbyQf/VNWD+anfHmz9z3KuFslFu7S3d3Ph1zhW1CHFQ8GnJp/meJ4
C4aCTADsqWsxBIX5PQeZzcSmk9S1OZ0Ympv8th0Z8ni3HscHnzggVAN47hNqmNci
giLhMSVpP1n9VpzNH/h+PyJRy7/SvrLQghPKgaYMYRm9xPDthiFs0Rkrb1o9Gp1k
xrFPQN5RsJut/GQX8P7rSrZzLbUEkYAcCIYS6ZC0A937NlM9hYOHKqZk//boGkN0
iGOhbWP557czvf4FGBMYINyq8AwI2n3vu7DvqaKmvDquf1kY5WmLQ6z2EEEoICQ1
pfUn7Gn6XsbCzTeN2YQOC59eBZhuuSBPsa+mp4mTK6QSIWg9WcsoGpnN2CyDukrw
eKmG6rD1RZJXq46GivmWYSFi3o/afKve5OsdNAfLQiEtz4XU1Pg4bk2wPlzIKBlt
WpfQpEPKHCIoXMVAPdVTHpY1tzb9d9bSOuFBXtfMKXf/iy6if1IyyUflBHn2t2WR
1Cyhyx62KJpOtcMqVU6fXkxCl8I/QrIDRRbIfNlaCHKiqar1h06tjc4QCYD1O8N/
6quNyvHu6BevKlin/2Wh28VGK387qA9Cj7Zqx4EngFkoUiB/YC4+9QAdKhFgaVar
gLUajFPCba3iDpqMZ2TI20y8+OYebTRS8hFczKyyZ3sodJNAwZGgf+6L7nfKhauk
6nDJXgg57JzT0HUeVWWfvr5s9je/d0ETJWQiI64KHNVlKcHpIYambdqrBczmtwpK
ih/ZOMSrAI/hoRTZcPhe9Nl0EZWUxjAOSCRHWHX3Q0tkF8OEf4+k+5HHcsVhrAt7
yXhpQV/ujxd7+NHHAXluhsVevSEoKG37N3JR7sc4RP1DjenErN04JIdLmInBr7sE
1dm1B0pl45snRmGAw8Vd8iLNN3hOOVVh792L8m978wunb+okbVCQzBbJ0JTOZNWv
ANXibkat4MRwbO17CN1EDtemSl8+J97k+DBdOxiDYi7ROuznWEk8K3GNA69XUT4Q
s9SYl4QQvLt27wGBNmi+sFgImrpcWKercUb2bsFKx2PfSOSD1oS08PPNoPjEJfRM
WfJyqrCN96jvUHAJYxeV97URHYh4FiPiY4Ro/9KM6FMkwSNHWxFikRLktmBrhg4P
NvgTDZohdYPNCj0vqSt86PB0Wmx5PhApPW8EwHzCwmMeUxdVZKnEO9YrHsd+oQDK
42xmldVfnJNdmxMwsBeADHQoNLqGSTHkyXfMjnv3at2MPUqBq7dem7cAugIMjthp
yfuGixotjsAo4RoXDFXVdA4JtKJ3qFjN1iiZ+Y/VrxB9KKfFM/rbvb4TNBIM+H6H
zlXSKsMLyjLtHaG99ut9Olu8PodqFLe/g1tWCm9519cjEKTGyjjxvkysO8XdIamf
ul6KUKhiygdjo7Gef7IU6g8yCpDeckYsOPsYxkzoxLVEAvYt4drjNV5OA7NJh0tt
NnaB49rTdNyv7jywTWJU31QRGGtfS+vkptfZsMig6cExtK61lr6o69mDrDfLTpjS
ytYyhzxx8mBUmb8TZrSE/izbCVhDeJCdeeuAGUZ0z7wquEYbH9CDShfl0w6ZFWl7
NLcb/yqG9W3xIUrFv2vOyconVaKtHw5N5+mZxwSdGigpmLh9dRDsHDQksxVjGM8i
zMI7vWOmCYYMh4Qkw1FFzqkMC89fTHGG56jf22XZd2PE8LuazshzxvAFU7+xdbfl
QiHvhFDaWkAuyMMyeweEpAKvZagh5fs/kH7L7xDoeOCijExMhW/NcSKZE0S1LSGW
vuq0+rEbEdiXBpoUxoK5TyQK1mfNxtzF+43wNPNhqWbDvK9tQwndKrJuZZAsI1Ex
oYTix020YxSdksgwktozNv0QeEGHrNaQeKeAIC98S6NtEt316ASh1H/fGD6eWgps
u/NbdL0y/srepxq41145F9DGIT4HZdh76nKOwfX2262aNWxRaJHWjtDzVpaW3G4B
KqG8cvh/SIQZmgUHf/VDfANPg3d6Om3qUCUg+eDyZz+TYSGll7tgBNIKlCggBj0h
D5erjK0jGsSzRsJuaZiyv8mBIEE7S1IwdU5g9x5Bh/Ytviu/S0b3WnitQ92dveAU
lwbcUgzUFSM+ZMD0S0vA98cVgyUq/NUrYRpTwbb4vz8Ndf67AxvHvP1OxptEFZP3
hiSGYnH5B+bNq+bY+vY6NiHwSqzvXWbhxAkQ8/q0RXvdGOJC0Hgdwi1RBzw1va0F
zZcqa64QGZqBjHmM9r2QKc07js0A6dmvQBVsOwRyqU06VM5RVXN3RfEjKyXqgziH
PV2hERWrRyFIqcQ/1TwNwlkvHANgx0XKu5Olhy9wlQt3K77RZuWl+Xwn1wcP5uGj
NP3/9SGM37xxVPzrrn4h/k5cNTrWI99iLlaj5vdsFhduLyZlS3Xda+72mz4zJJ/D
X+3R1muY0XdTRwhoAR4YNCWdEyBq90B1sAZADERJliiRTU1ZSUqWwqk2D0W5oj8b
0lEE7v+L+6sAstqFAbRjguq0OgYPY0TOXGsK2pwK/+g5M+kotYfGlD8sK62pLUIL
/hjYSx5kAvyoyK0312gu2T/+RcTBkI6LmkPH7x6LNV0vRVzJPNcTdVEaiU4no2zu
20SomRLFLgrCxrMbBPZzdOCT3IfHPNXjl/HiG8yed7wpuIFa9/4SitBjF1KrtrB0
4aSoV+RFh3aucN40DoKC2X0wVyJDRGezPMifYlwVWy93jz0AtxEvv/oUZyLnEcue
CUInJwiB4DC/jYklBf9b5SZ850zbNtQG2HXfZZ6TihxoRBandqpAWFMM4g8W0VeH
gyu178babnFqcPXp96JaLvuSACCh6N6eqJjVu+ORYUV3goJ1UqnIKRO28Ovn6dAn
V7H0MQR3JI9zKmfcsGu9jvQPnpjKlF3KxtgAD1f0PIs7vrfx5o+qPBNDJau65EgY
7GBV6Hd5Xr1ocy5KqPdeHkvMKYdH7iT3b7fP5CNkwPcifxxNH11gETwvOtXeIB/k
NInEwKEktqrBugy2jwPRnNEymH8azroN44RTs8mXKZ5KCIdTtlvPTDEF6YD0k7dZ
MxVvu9BRpriAwoM9zfE7/orzxGnKGuuD4AguJCjHl0bv2aSH0N8jM1GopdH7qFmH
eyeLHR8nH4I0+euHn1vxni8j7JJtDjFRYvHN8YUuluR2xvsTZnwPRYsWa8BSukbV
mN3FuVJr0rcX+VnYOUN+ULi1iMyNguxRo1GqWhsokjTVBwMjocqSDIr+YdFTOwlq
9kEbIJnLYGQCcgMMiwVqmeAlvOZ6z4UTWKIcZM91tSnPRiXcse7qZJZH91ykvggI
cCDPzV+2CM3UYdzCzcCmpJx6s5lfaciYpEDEDRW+IQLJwlMvK/pSu0dUa2dhijZU
0LuXB0KwrIcchBcEBsGufKH+IJZdpGKa/oUWFofR/vmEXQdO89Dcozj6Tt7zJw1L
Hil6z3nJSfZrt6YuL4P05cI3SAPZRaDDPpYvZ0n4DXEo/Me5H1Taqp7u4ExTtTPZ
LBdPLkH9re/SFae9XgpACG/FwwJFcOdNBe9SqmD1PWSW7ae8KL+SEte+zab7qzzA
TRljG+j99t8mO9NR/rVD8vn/0QzJ4+ihaQzJOq9UP8S/vMbDSllVkhw2fy707zM8
Sl/SzKjdxijdKfMwhfWCIXLkKwSmMDLiZDISflmEqscF0b4k3ZMkndIYEZOj18vE
W4qcJftEJvTiRzSqZJWZDj9O0LVobr2MAn1CzOdlHwa/4Og1CMBA7lRrxWPn/gFx
zo/48iuw9dGXmKhDzPvfWA0nlLTvd5xOVJKgEb1uw0ks/UWatWkmWD/Y04TJ1AR/
YAd3CWvmSVw5EqwVpiit6an0wmImjfauNMkdCJyK4AW+RzSdQBaLqks8UNM14+o3
CBkBw25KOlCEzGMJeXrdFZ2NuRZMo+/VrFzXna1UDxdmu/yMHfQ73fCrwz+prKKO
fjg5ZZV2JGfVjLPOfzLfR5zV3Cz6EEw8j6ce8om5+k91bLT2y9elNGwcORcgbUG2
7z//qS29VFvGeKP3+tZ4VLA+uDNO5gB4OHQ0NRWol4ezQ00tQ3o8xk+ARCfvqhTw
J5lsr/V0VtGy4JhWqvFNQzBz0E0/m6U/POj9a4ZlBqtHbna1FgIXdWqL8jPbYv7t
vn7crbJxw+mECPy8vuMmbB+3X8hkNNvKKtYq88dzQHRrtLiLI5sRMgyB5yxaxLC4
xf0236UIubvKjITua2zFnEm4ODWWFQxYv0fb5zuJXSAjP5FZRgt51JYRvYoXBcZs
A7Zkg9pPRGClptK3MVLCP57mB36sty1KnpqHZ9cQym+yZkFf6u08IUgcC6ZKbG5r
8UQxVWR0wI4bK3P/QutxjpLG5h331nRraCehmOrU9DMDW6J5kz+7QeE741APY7Q1
jWFMZDRKnBzOfEhflBUcN/2idXG5Pt6tVRdx6h90NuiwJbvgJyV+aH6GgSRVeRNb
NecHbm1ymdEvnxk/FImDHYfUrYrkZKmO53oVuDpANrihME4AG7ZFolNGF0YfpENX
wC1tvDeesgaMF5AjINU7RGJzdNuD+z0y67dsd8JDvdAbELbaLQoZsPcj3lk8JPoy
pbfJXZqpDkKNZM77IFLlwHNoZFvashDS8+BIdI2LrpLu90zLIBfvjB0CLgZy/Oj7
JdDdG4axIdZbiO1aKNtvrnhdLuNw2ngvSv4kLM8EUURK+obxtX0/1vXgFg+tRQ7L
6/PQBbWBQB7jVqrdZxjXBZO9aIdacPSH9iJ69S91eJauwzgRYScNZ/Kj+lHxD3ER
L/DBvPV/QxCpcoapRw+kS2TTL7zdkoO314QysPgg72Rhvh3gPbsbzhFcjxak/rGn
XSlPSIR8yqcL7yIaiwWgJDn8IKHIaN7RIIuuwNzknm4ie99ql113UZMS4ui1emqU
qbdTLX0qgyJ0cPpG1KsM00cOZALquxcmHdgilzCPdqEfe3u5J43KZkQWVtlVgQj2
xeVsc7+9saxw7P0Pu71o95AJYgBn+PgQwWOLSxRU+bWo6jDJHdhqtT6dnDrTK6Xh
7m/QM6UPHV/awKns8EtpyfdYYhCw1365oUBDlnIjZLVRlbS/fgF70tTKWyEBlmVT
bHqEA8F9MDKR7zBT+/WFeNTMNQuGSMb3jWs2WrTEbG/vvymj0s4iNxtVjyS7Ftmt
7jgzx5ZYUc6wstdN/bkk/cwnCd4sLF48wmfcuhcVHeh00b30UelL+aXxV/cRo4J4
L4xgwleCSjraCfdzpzUdEs4bxwWL5YLaG3w2W3FwecCHtso3ixZyswYgSWu7XVGu
zLb83QPr89FzfaA4OZTybaat/xJVTTC7rWNRX5oYBf9eZFiRFas1n5a8CPQ2v9Cv
hFQpJnkxXaRk97aYe/2P2HK0cQlRN5N/aymgQmyEVu2BBNdzmJAiKJ1LWJEb58i2
d8Yc3Qyu9OQwVDOxTJSuQRV421No0UNbOd9q5jucQ0AyW/S8OE4qBcvfkZ0lMF4F
EzU9xbfkrP4wbJA2aF3qUPBF7Nmkd+VIiwmtqA8HJbEpvhXrVVtrD5sl9Le8Yith
jBch1mCbLaXXWtL87ZfBB7JAQO7WIy5FcSfAO63ECeBVgr/2Ayo5K7PdY5y/8ZM7
oP4SVemUkTuBd04uPnfEbgpeSCXVPIssDAYexpP0Nw9Fa9M9JlksL98IBArHepML
V96bthmaPtdXwQ5KzXOHqCln6YXaR+aLWMvTq2x5QFbxsM4ch5d+suTj6krHRT6n
yi9S80WAPvxhwRJl35VUtwg2Rn9D2ZNlh0tDM4qqGz1ItfKSKtkfu6JOUWoAEeu4
b8hKk2p26Q4wUuczV/gFCrVWhGuEXiehmeMLyX8MA3ZGmwJtSVkgqLr0R1I+lm3M
3St9gwpWA3zLobY1iTQDLHPJ6xJ24HlQdCU3rYX96y0IbLXcX4z9tK3sfSa2B3Jp
dc2mhZv8wxEYbm5ezHC6nxA3PAANL4WJ5Ygqr6dEV4f+/1QypYujl6CJNs1vxck9
I4o+MQUVFBlD5Xcz5d+LNShqYsdzyntyInNfRA7DUu3nk2xAGPP7Hnz8U2rhpwAj
ZGLhAqSTSltrcOFGCJdaHWQeCoetjl7mAAkCiD4QsXH00e99kggUri0k966Ukyd2
NNXkxfHblyKVeMXaqbGweDrS5vn+ymqIX5uIHUHHCFgQb0stczrj/4Diz6x5YnGG
ZYKMB0iIEjdCVHH9m/dt/6TA8S3iVcKKYkwE4wJLJA5v8zCShnzrjBgOD3q86JrC
XQ208e66R7LuZqgG+7Nnl0qbClUWyncZ5EsdEDbeUaRLMdVH/G+Vwr94U0973o+r
ZmcUvBbVr/7+bhW0TL8naQoADelWzvqP2bsW1mGFNnS8eMvpyZyMJg4AawyXGJ/I
Skhs6nLJTDfZwwQUslfxQ+LjRFgD2orAVjIB+/XEDlrL0jgaPZ7w2l0m3RDy3Diu
nttg/mODKwiI8nm4xQRMoZGnSjgXEDKFFSyc2R6MlmRvXDqRlq3cOYeHffE6kNl0
0yCSfjfzghA0t4Alb5OnBKt3nK0PUocY3jifAM36tVNFegQFkpP9dYiUoL3rUf8J
IFmfzeiTCSw9qbRKecTkdhFUzsbExlN9EIhY8B/hkc2HQGfHsvjvNgQ+hzb3aiA+
zzO2QaoOXlGMXcEb18P1KuIjbu5tJcpIHEvqONdnhHIE13DPs+FxKnUxkSxYu0Nc
6PKOIPMt5nWKina5AIMB/RJfGOSc6NBI7EcXgPRfykiSerTR+N0vpSpKoTF6mfGC
GFaHR2e3kkgtpOHazGaI2VjzwWVRUTOggfOU/7V9WYxxOL/4SPVaEvCjKgvgQN4E
qkno95CZ5Q0m0kG7ZU2Bc5cQ9PIh7yy2UE7x8+8kzJyc6vvt3yOZ1vRmtFJTYIFE
C5bq470zR1RUEBmQEeyQ9dMjTokw2L+S0nVFuenWB+Bq6VVxP4NgZ7w3atAQPoTP
C/5mqPC+WwSQl4M4RYfcmEjVCnqeS4ECWHFPehKXDrAdbvcu06vMQrzXIgYd30Nu
7SdHBlaIw6dwxKlrBgkUI9AUIISbjFMHv9XmQAH7xK+s7IFnBPVR6KLKOrKNYPh9
AzrT8rOgmT65/b45GsIxaT5wWIMcW7jgH7/KXEfaPmMlQRaeU1b/6StMZzJu/L/8
C19dpVQbv1NIxi6JkmXBVIK0y3qJ9bIskiHcJrxFrcyPtQiPIYCK2WVI9WJdOwj6
rIPEYc2Gg/ocvKfZTAtOWlv3+UuJPw903K2WeWwFl8l6aCRrPf8Q1Q8YroIJgNok
9JVD4W+f3JydiGuHuz44NUwhHZXGYXqy3xRJrjalk6QQP1MGTx/CwILkX9YV9wBo
3fIXsa27DDoeWUVPf0HnkQtZ/CzqZxbK2brmalNAt3xTkgjdYCDHAw8LHoIvZu7F
wStiBBwD8iQusFJaQ/jvstMXRXsW49rEyO/Af+hqMKLB4p6Vmh6yRwTVF+a7mOuw
JZcFyB6LBslaNdcml/uoyMAjqN7loggdtGH6yuWcwXfnj6fFK5tJzhtuJMQLMwW9
8uCbc8EjkUreVQqAv10qg3CHwTEwIfhlW3BJK3ix7fNbxgR98jVOtNyhmCkiKTSN
YKpNmlY5oFvSKrRYEmGYFyaksynYoZlKom/b4ilvYx++T4BbHkYi5zx7H1jkw1Fo
VxXHu5z0dHev/R7nwjbh/02Jwy3jopsTRuiqxmNQrvsUWBouDtfqOwzdqfc4wSF6
zdKl1zH4GcDGNo+EfT3R9eCUCCiwAZaOPDbYxY0f2VzIOgzJQh159RCCAgKZmTGh
aAd+dxClw3e/GlSe7u2Rw9E80PYDI/cQh/efKNFlU6Wjey6kPeKtHeAmoKlRAwBB
Y720j1dJSmnewHjzCyHKWhzBtBlVlaPdNQrb7i9bYpZTRQS3FCW3bgeJx6J3xutC
RS9cz1wCOAMvKs+r7+NQBsCssFfjiJlw6xHQcsHBcfQZ1H/hGSt3GgfdgRfIEDEC
tLpYdYCw8l8vxkAaCVj/whvfPCIHAFkTr+IsDHqdBP8LgO5WvK+4JsEj9jgrIk8e
crCPLZnt/LbovDXxzs7aYnn3gm+oeb/hDpHPUTjh3LYBG6Tb+7+xCrlM3hsdarip
aOx8zzN9cxyZapkRbvor6+FVf4RDZ96deBi5SsjyQkCzRBhhm4nx2yduKO4xP1L9
eISeudsmcS0QnCuh5I6UTumVcg5HV5LCKKa9TcKIFN9ygFBj6JfwuyvD8OrZyG66
5v82h95tereCZ0772RE30530j7Bj5KjmOOQ37PYiCLvAtF2jHlXxB2H8ABdJH7zZ
4J+Y67x7eh93IIGCfpLWxmr+ZxZjwcTTCC0Fd0rt4rJncOG5ssGAkguakxW//geE
eey2l78KAZOECW0/9QwjgsW8ZayXZN9/3EtWAbK//Gr9roJmIDvwI4nZA51APK9S
TQFiE5vWMm0TOX2moO3LEeI/qzf/eqCj5q08Q+9DT76Q6OwjvVXYdQnfVzU97TCb
LlnjutFobPQHOlsYsZF2yjZhNbUVIKNpSy0Nhr7jK7TxHabDSKrcfvRhakcJN8Dh
ldWOivYOxpEr4C2/SNvjFolmKlhAdEDfGJQVTboXdyEmybwe1F3VXrtclvttxVbH
NkXrCCH2w7sz/nHMhgsvDBwTC6GuoUMA5azEgp1WH3/KdyFpTB1awnvf6W4okp10
vyxFjR54FU78+CCj8MufO0uIuQVb1xL147Mbtj4aqyGQEkjiUYWOr4FNCEtm09YT
TKqj+6G/uauOS/+Eo2I3VKTmSVfJaeEvlEAeEmYeVSlTWhAxyeAu6al3BBExX8qI
N7p9zZeZNxTNiJBNUMlIUFqsjJCkF46NrOLetuRuuT7PZqDCnS+Rz9Z4EK9IdY+J
a9hu4z62kW14YPp46m1hRBc/E7BFX2Hw91FFK3LdXKSvhUEOnbJNtZFt3OLu7oS5
Y0zwJikZ8SbAwL3ebC3HzpLceXE+j8TzQnb6BS5AMgXUgKs3G8GrV4YELPXqri6A
VnBvruLGpqPgS/6ZhkV06ZDWBE+gQYXm85a6KNe+xceO2fb1Wfo8p6SqGysB4ZI7
+RPIYcEsGkHdPTBEGranmFb0wPx1fAC+3JVN9CdQNZd9HZAdSoin/5ujFLGW+fJ8
9XJD+l1CH8GU8rpQ3fupS75IwrFTI2TfPxEIFLcQDzccHaVYYIXUtVFGuhKVDNgk
ouTSC3tpO7qRBLx0a9xHoEU9iAeJvExub/0KFaVrwwqbBOUrEQ792yV7ZT84gBPB
THtMrUERyn33u9ce8+CKqmKFn4Qu8jnqGPhXSXEazt0yjfPdOvwGQOGWb5NcMIGh
6/Ss3Kk41ntN5f8r9LyZ2YEesNuIxe+R7VUKki1xnILnLTGl5u2gL6Q2okV7x4eX
DFOYbJTFz4I2E/ZmmIjE/pHKxTGViqrZ/5e/RbvVZ14WDN7CcTI76QZ1HLYL3Pr6
jKRZtBNNus4HZ013/w2eU7PwvMXiBS/77/rlvykxWtZalxGi5cYNdp9Q7mJJcvV5
cQA/r1GkmwpJXpkg5b/Tfm1TpEfsAI9MTbxVVLcGkCrK1H3UcCV1lQA6VrwHoGj+
79vsAmxd7fbW/jIlz1rJYakR19N52mJTEBmyPIAbt25d2t4tSF+T68j2uWk7G3G+
lSR5l1srmSjObP6oaa5m1/HuCuYpV4fpqVz+BCT2NsmimaLa+0cYHYkneZlLBjbG
weDyLJhnDbR+ANtVfbKoJ5wtVgjJJx6M1+fgsJAEVZs/KVdsfg0a3XXN69qw9zik
7AEoT0yHBa8+Gt97WA+XYNiZvxPX1vBG3IUh7Dfv5DNiYzHITE7iZIcw9adQSOx1
B+7CGwfHpvRSAYXG9+JquzoNfH+hfLUQf3uhd/I43naPlIMCcby3u0c1k8uU1VjP
pR/ybTCChpyyQ/jENR/5LnpC56zf3eT1tIBujOXxOgoO2wzK+ASXjD/JrwQdQypo
bsVnVEOqVUueLp/Of9slUDF8DC0kj1o8zn9OpqHURLT11UqbBGshvK++uVDNCnfp
FZEPunP1uK9pepGTmBqERB8R9hDcI4Y88dxgUONs5mleNDUsdTbsJArkhB22dcWz
3CVeByeP1TwOxTVH90PY7k2t1UdJfRop93Dc4kr0gB89Q7NNko039s8QIYHlwM7T
DhPjDlbBzYo4jH2jjZvPJ9MUDVi4K7dkMg2WhVA/2mFswAZ5uwxfKU8ukiQwrdXg
CwxYZdt3qgdqK+9X0/bfBLJIuC/ev1RSihVGrp0RGXRjg2Wi8pWt2/Z2YJDJgQLZ
fDzfwAgQAQX1+GwNj6Kv29TDrhh3sC+TlO8usZKhWQI2NBKqUV7sGfXXg2/giRGB
2VzotU7UXwSpTzA1UdQKAxBMK+hZe9QXWno0/RzoyuuXNzFIznJJ/W2H+Vfvcnm7
/9/M7GZmMxCpPYsxpEUE9naajM+jsjQevoKZLMiTGlZCgV/rYMXYP4VVrcjBzb0j
gH+Go107pbio7j9tIMPW9G8lb+H9qrDNv3EYlUpiD1znaP48MIbarEUx4VYZV+H1
A6DKdUj5DkdhncTcGgl/Xnr1pBnIX2xIrppWV71erV3I7xya4IsT4yFaAvL+xdmt
MJW1STHsdcBV8hu4lr3QSlU2g1YgMp4bNJkfsdkYG2pIii/Ing5Y60T51GNSghPW
lSjMqCHDOKdXGWLkYXxDW2lDKTOa5LcBkuj4AwGQrxiMsiIUA5RJR7QVVMtJUh+/
LBhNB5F/XWONlmGKypxPBCaKJ9G2H2uis53L9hNNSiLqampJuTNzBBs0YyotHQPe
SZx3cczSO5aUt/tef5/Vjy6bhZQwfMUHXYWIX+nGxyLZ+m6jhgu/HdENOgcAagyZ
TY4mIbiPH1D0Y3xIWu0bhxpDtxAJfsa3NxOaniD2nykhhb6fCpMHfPHPCy/D2Akm
udql6IWWDP0poIuHkgors6olXDZwx6S3GuSgiqw22EsvSiuWQZaLsWY8vUEdD7Iq
mhnyIE4KTLmNpOXdicIyOOO4aUQbmUF5ji1M41cFQ42vSD2x0t7XgrZ4qtvudas5
V3vJtWhUUNWDV3wp3hZTytC0jj4RLs7en2Byq1Z8VssoxGB8s9xhOj7SDJ4mi8Eo
L5XxohI+q5GXln5orOsHE5ofVycfuZnjWJd/+BVOvl7a0ytsXSdK8sWyZbQwUCL8
FgzhbekZBGX/SAKuFl+pE/msV0hIPcLrCUy+pztmDzqjkdYcriqJtHDfmnD5jvGV
Q1+LlkKGQEiTIDcsCeKM8SYUMo02An3bdQmiwh/eLtxgGzjha7aYoto2IId47okF
JTVtk7qM5Dza2TIjNtAb4FBT5H3BHi7h7FbjZe5rYgAabaEr932ZvUVCCSy76ujN
YsEFXg24OpkoRRbaZ44znvFO5f1eB4xPdZBv9bi0xtDufUzJIaGQMgXn0g4z8/wy
dI0+ReYFeExrum98lReZZShQFEyhx0m8xnm2Eo0WJVxEvtwyDZZBL6tVklYHjIwd
`pragma protect end_protected
