��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�y�Sy�;��>��&�MA�)Cʌtg���e�8~�����=H�9����.k������U��U�Xe���M�b�(	
'�m��_�S,(
>ɢ&T^5�[Kم~�WA��Mb�c#�<˃#:}��6͕��F��O�j�7���'AF�9��'�ƹrq�9�p�
o�'�w=��v��("�|��ӏ�I�\.�V�����)���cB�չ6�t3sꀚ u?�({��_x�W������!�`�e�H�H���|�-�YY�
ꆞ �Ӟ냨��e���S�kFd�v�e����y�*D���G�>����+�ᩜu�f�x�I���*��/1\1����r�2�*M_�4j�t�'{)ȳ:�A��!���ש��6�D`��Js�[�a�O[�G�O.�����}�9�����E���;I҄0"}̙�������@pi?%D;�4৶��q7�D��g�פ*]�cK�eB�Liu��nC<c��&2J�g�����qU�d�Ɓ�/��Ydh ����E@i�{�l�ka������a����b��b�t ���?\��|���1��Q����IrG�:�FeQ� ���Ő~"/9}�\]���x����/-Gĉ��U11��)ㆍD����_��מ-Wn��+����W�3 ׆i$�e�Ch[�/)NG��hAo�iv� @k1R/D��\g�tZ&��7�}sF��#��޼�����m��GJ2�?�6�a��:�p���H�v"�
�nwf9aX��v�d�UU�V�nӁldG۲�!+�l:��u���J�Y�/]j����|��g���c1���vp�O�>��Hu�k� �4#X��mF'n��yy>c��I���'���	�]k���*�L��Z�`�On�m���٤]��:��J�S�2y��O��`)��J�f�&KM4�L���LuxP%�v�gcTx��vLd8Wz��4Dl�ك�m�5�g���Qz�#
����{g��u�q�z��xsぁ:4W��4���3��X���|��\���,��oA�x=��h~���BT`L�_�&z�}U4C����A�A�u[�Ex�K'_��aL!��p%���6������PӚϿ6��V�A'��Pv���>D�0C$��g`Z+ݧoW���wlc@;�b���]���D�wP~;�ٔk��a�z
2��C�g��V��1h��t~nfb����4����Z���#���C6ecn�^wj�k�x��T�}SK5�&��&�W��h� \}���v�ȎĪ��ĨCz��Uc���q�
�g^��ʪ��|D}=����1s�����H��\͟�䶆h	j��<�X�<݈E��s;��C��xw$�R�7�Q���HCX?,�u ���:Y�'��i�U��xx�yf��[˲�xk�q�B)/���c�7U��d&��'D�A�H
�	�QAuu-�:"�?爧;,>��J��<g�wp 7�䟛u�r��
= "pNa�pWAJ����.�fі@�yϘ�a�n�w�sKm{T'
,��ț�~����m�Z#�)a0Q�Jti��fw�<����!5U���}�-�̍cN5�C ���`�EV,~�6�@K�(5��6pF }x�ds��,0
|z�~�fx�8b"�1x��N���Sҕ714��g�zXD��C��o<�^т@��:�Pb�3~�����CA����y�cV�9��wt�ςb��l�X��J���~T@h`�%�-5^v��Q�J'� ��0�v�(�B��9��R�Jm�	�ml,�|	�a��5�p'��H-*��vl3����RߠcXۓ(�M�d/;�)k�4Z[p�mR�a��0�J@�7*i	�%<j�!�k�\YZ���3��l|9��Rj�:s�)zn�kC���Tx����x� ����/�{h�	h�}�D�Sh6�+�nr�\~g�0��K��ɸK'g�����s"7C��aQk�31ԾÞ��b�A�u��D�	5�b�$K��N��1K����f�><f{P�Ru�dMd�-Ě4���`�1�D�W�fM��J�>Á8L�%�-9�9���
B�X��5�F馵�s)����ep�b�$C�e}QT����
�?b�"2Ӹ��0��c�_<o�cV��IZ����?�h����H��<E������燎����sbB���r��p)���%�)��c�ya=��[D�v8v$���	�m���N��^�
^Ris1�D�<I��=���	��Q5�^g�R�S,9���u��FQF|��X�W��B����r`[�d�m&$��Vm�fXR�-�(%����Doc_7d�:�s"[���1*g*�����X\!vF�0���o0r��j���S�xCm�I�ȟ��$/�#����h�H�������Ѓ��.��N=�Zؐ���N"G�5�{*vCAu���ȝ����~���/���#q��OhL�u˞�c��>������dUja}���J���6!|}�����H���6bmF(Y�4�3+�~�[�YC:�B��4C�z�Le֕/�n��P�N8��ե*K�uQ6s:�d'c���
�1���^��q��)�cm��~�4�:[�7�}��n��]���*B>�����n/�Ay�5}]��馤mh������_�]1���2�y��~�M��Z���-���|��{�)�^-%\Ui��g��aa�'ͭ��Ym�0�a�����������x�?�B-��b4d������s"�h�'�4�ŀ&���U^��~"�֐���#�?�C��\�fȊ=�ͱ� �/R�� YV)�]��Jnx[+���Iw��EgB�T���t�b��N��_���C����qEf�h���M���^!Q! ]r�>� M?QF5+(j�K��v��W<&��1�&��ؔS���Un]٭�2$y	ucЙ��@��
�t��I�j|o>0��.�W�]��f/y��<Fϋ:�����M��ޛ�g�DhJF������^�"��i*k�k�F�\�jsd���n��[i��Ҹ����f�9ظ�{e	m]m��tm�n9i$��;�{*��=qrp���t�c���(���h�76�jRz�J��`��F�w��|�s����[A���*��@��U��_���(�x6BaIP����R+J���8���(`Ŗ\+%�3�'B���CJ����@���5D^m�
�g��RfR��t|�Br���Hyj�P��7'�<�1�f��A��V�Q���� (Vm7݋j�{}}Sn[�:���J<�r�	��Tp�?��
���;�:�N�k7C��Dj�}�2�Z��	Aeb8��v�q��S�afp�W]����l&�v-�ɳ�������R>�p�Uq�����o�eQ �gx��FvQk���ʙ��9��j�����8'\[-�g��Z��k�M�;��'��Raе���\\1��+SZQ�}CcĠ7Vܰ���u����7�%�aa,4��+2�����ݍ�?n�1$n���ta���ǈ�C�FN�1ڡ>��yhO�e�{�	�V���:� ���LTR;�ܪV��]�W��k7��x��o43C[��J���Ț0<�C�f�`�M�9��E�c6�_*Žjh�ro3�<�/��I�㖥nZ�� ���
��`�l�KG\�{�g��U�$�p��Y�`c��VX�˛O�7��Q����r�㶺S��נ۸
�(aV�N�Vv��;񦱂<��Kƕ��L��At[���t��!z{>|��S����S�s�����ߌf��O�j��!�E�.�D�-#P�e����2m{#��SD[��kqh�oLx����^�5�Fh MR�#y�`'��Pcg����Gs=���Ծ��|`���SA�ϰRBsea����bzǥ,ljF#~�z�ٱ\�c&Mi���=�%D�E����H�&p%̞{�v7����M1x�����3A��pWܴ����H���u*���R��z��7���lU{ci�W�3��7�.���qJG?#�@ա���=;�^�>V�Cw]q��Us���^�k/���p�KO��;��n��s��ԑ��9H��T������T�
&�-�����iA,^��x{~y v�3s80�O��g�:��Q��^b���w.�ˇ��S�S�)&W~n �A�Zf��0�iu��%)H� �DX��:�Df�����2�ǌ>�z�B$�ܔ��6��D��1ہо}�Nz��T�Y��Yc$�����̂��gO�@�����I��z0۸��K�Z���%|17@�����g�����:�����=8�7U�͜4~��
�Ӄ<�e[�c��dJ{8�"A���Aj�#�q�,8�iwΣF���L<�.D��q���tA_\p�W!6������Pr�72d��N��﫦�6\6�&��Ug]�� :N�(U��J����5�3_)�2��.�m|��{ftI��c.ˊ�K�4����cBic���.&�P<y�o�kY��<���O�Cą��<�Ѿk�ۻ�\�F���Pp�6>튯���N1��Lg[u��Ĕ�;A���SUIr�$	o9�pU!p�9�0����r�/d �RU	�f��i�L���^%�����~�>��ɾ_~���ئS �7C+n 9����s0m�P�d�p^���	�,�,A���S	�(J{֗�^���F�`�������!����o`e_�_g�Q�/�8��2?�����
�:~;�����6�t�oLݯ�1��7s����,�/����ۙ(�
��^�GM"��Y�<��۝<�]�-ꕈ�!lK���nE�]�hђ��6(�
�����S����])n��(9�������Ph ���u�y�k�#������F�5�<���Dc�b�+�*.�gut�[�s�7*$/���E�g�^�j������K�x�w�W1�/	��ۍ|o�m��?�54��Ȅ$��v#8|a`]$���>`T�$hu�+��.-�\��1�kW�"m�v��1�͕86�e9%�(��<5q�2������?,M'tx�zJ�U���}�t� ���xDB�bv��?��{ףB��1�%�m�*��`�7�}~�/� +��	Z��_`r�ꦶ�t��e<���>�����$NEu E� t����Y6g�M�D�O�W`q1V�넢�#J������xĆq/eA�9x�D#^H�����G\�$���<����T�CC
'�D��"��1B�����k"���_�d�3��$��h��nţ~+�� $�������wW�>�)�]?~.�۸�e�X5�1��`�����	��!�n����'N��A��N�����)�TA�hug�&R�b�|�6��[��u�ϣQ-g|hע7֌��2D@Q���T�0	H���.�W�aTP�d�կ���z"k�#wp�u�q^�mǙW�@I+����jX���He�FJ���@��Y�7�������O�J�
j#��/T�#N������Jv�4��s"�����?����V�����C��xf�����(0�~T�#qgY\��q���@A��ĆR{F9׵��Ȳ�s�V��m�Ъ>�TdR?"�}'oAx�7���őg&S���,�m�>�iI>��j�d�\��o�p�{1Z3��C�����"�7�)-S<� ���s��4
h����?�_vD1�Σ�E����$W^/,��i�מp��o�y���&l��m!`nj�7^�)lB��D.i�����9�G�A�7i;�<dy��m�c���Ay����v���vp�Ԋ�W5#A334�������'��!���� �q ��ޛ�i݅ܟ5�ؽy�3blo�@^�9=���J%�Ju��V����i��?�Y;��h>��k����)����׉�n��!ʅ�Ny9P,gD�ׇ�:�^/��m�{E�N�яP%������픋�ޓ݀�gA��J�*d�.c� ��������be+����b[�V�ơ+!��M^`�=[�y5���$�Ȏ�{�O昗��N�F��,��%�g�g���^r��5CW��d�LQ��%��Q��D�H�;�V��{�@8zS���i���jb���|$����B�
�D[O�D/�E��\¨y��rq�5	4�h[O�j��7}��v�xI���.+��h۹L�j��zv�tD���{�@����n�"����ٝ�`�����S�?�$��y4z�WN��I��g�th}������C��V�f�G�~`��ƕT���Դ�L���7�o�n4���*��o�;x���C&�J_Y�5QH"�T�|�>�¤1���H��=�=du�M�~y.�d�I�R�%{���)�To$a�/��)COL�+f\�r���"~w�'G����\�O/D0*�k��ַ�y��S�v���)���_ZS�>��r�B�B�9����������m�X��	t��?W^&F�ڸI���P�.v���>},8;w����	�",2���uN6����b٬�v����m��'k�Q���N��#�Q	HYo˞��;IG`�K���F����w���ƾ��|3R��`1y�Pk���|(�T��C�(pbmӵ��Npk��=k���6���ue�L)�����E6�AO-Dj[����
��;�$�B)�!�9Trq�f-�B�E,�z�Yx�{���۴��*�Ig�� _���0N!�8>��e('�p���>r�� ^��u�=��C4s����� ���ӽ�R.3��K�M*�C�Ԛ7�/�V�C��ZbB��d�U���W�x�Ҏ�R�0��.����^I�=��Xg4Ox��K��q�IH�����	,A#�=g\C�98�Ys�mք�C�V�4�!���������Mܕ�������uQq�`���A���hr�L�6�U�K�1��?��(�j�n�Ƕ�ՠ�2(����t&�\18>�� �$?��Ra}�h�,�ؼh�![/��2i��:��FhZ��#���������1e��P����7���L��|)�c6��/C���8�1^b�!J˾I���/��ՔE��Y�L����0���ā��cFif߳]�2�Y1��!u��a������_�B�*� ���%q�"�.�0i:1'>�t����/�\p_�L_��6�$�b$`o�4����k�)qډm
�Ap��	l*����Ʉ�_kr�}�Bu��%,R���B��o�֧<o0�uNu]H��Sq���
�Rl�7P|sӶ}��n�:so�Q���^�%��/i�n�=�#�rS���M�h�#\�\�y=�7���*^�dvP���ꇚ#O��;4ωL�$�WDM��]�{4�7	vS=&�����#"�9=���#�E��4O1�Ud�����s�K�w�[-�j��!����x��9@�m��^�v;{�{"�EF��:
}&Nɐ%��nay���^�>	l�>26�/1����'�L�`���3�&���J(�ݞ�ҿy���3����ԍC�&Pqm�kYdȝ��xe�Kr�m8p��K���==	�ԡ0�&��l/��Ҵ��^�z]bs�Z���/{�!&�8
@-��h���W<�{[��+F�ި��&�էݎ���y��8G�T`
��3��b��dyӘ�}ڬ��.D�.]S�&��4,.�k:օ2�i����q�H���Na�jF*Q<��z�yz@�+�o�=�ŶR��{�J
�/F�>ǆ*�BT���q�rҜq��N)X��R��8@����S���c�<�hщsPjg̣�ڼ����|�`"+���t�*%A��g�'
���c�|"W{��yЫ�q�{�vC��M��A߸���'�5�����GMP	��#L�9I��8!�l���=)4+��6ð^_��ņ���Pu��9�=��#�7E�
~`ɩ�]\3�_�p���?h󣷐l�L� ���)�J7:����)���)�q��-x���mB᫈���6����r�t`�B��K���̷�����Y����3�v	��O�����fi�SE�CBz�Q%Lޤċj6�%xZe93'��c���Y!���� �I���7�)Jn��_~��Rg0�
�d5����]N/!�KL�O��(:�Ml��YV�t�{(7%�����0���UH�AB�Ae����3����ͤ�	j��rԞ�G�9�F�m�*&$�ψ`��3��Z! ��%��A��w��x`ȩ������/
`wU��;�}�0�1 ;G�Vi����]�P��H�Rr�ު���?�%�)�"��1`'�A�7Ն��U��Q�(���o��F�W�Tne���C��^���U�7��H�w��{h��V��n��̱��_>8�_��0�����+�T
H��u��N�
b�A�Iy��EhK����Z����3x�&��9J{RWm4<⋻U�v��m�����X�5jZGU�U�m��DG�OB��8����Ċ�s#��n6���$PYv`0\(Ch~��kž;����횽�����U�S`��_i�\��������Ӣ);�N? ��k�M3��9�	k����,�SD㈐�3q,ӲP���5��A<�����4a4_.E�R̟�n�� �=-Z�w����+U�K�G��nO��h6�4ۦ�y����U��7�Tq:�?�l�P�E����3X`��;ݮ���&�a�7a]\G�2.te��4qB���a@�j})��h�����n�$q�@�(��*	m�gYE���̈��e:.��m�8#
����h'��6�����_w��ڟk~�@�������'���G,��	~N��]}��e!U`�~�}�8l⼴���t�sd�W��Y�)����Xn�q�!d*Ѹ]��j�Q���c�g�X
�\@Y;JV
	�*�@�FB�8,»��#�aӒ�{d�I��Ĳ��[���D%��.?3N�*z�%+w�ǴP�!o���,�1�t��&�uc#�.��K�� S����)v?`Ϳr�>�I�;�|�t����O����~�!�l�$�^>P�%�G��Q�h���o�`�:��~b�4̓7y
K�|cFgJ��ON�i6����%�������yչn�7��={�dg�����LK|�v���t�J��A���.m{HC�;*���q�:L�$�E���{��OV�ݔ����&&�!�
B��PX��zGq 1�SkM[�z0�������w����=�Sy֤��(��NLֿ��~�X8 ⷊ��fa��θD\�VVSR���1}j�Q?A�
C�J����5K�f�������{u����^߄y\�Y�����gtG����n�v�P*Ĺ�p�)nZ�R�T�ʎz{ �N|�݀퀱�iu�آ���*I(s�b��%_�t��d(�_p\C��j^�_�p��9[�oD����eW�>��;��O:��TQ/�Sm�-a���P{�H�+�J�>U�v+,ri,��a�3J���<�p���J��M�bԚ��ڶt��	�`�H�Uz��ob��p����g|����tY��c�<G��_ ��,��Oя�F%��[*KJ@�77*���6�乳���/�>s~����b��<W3�O�wΎa��K����T��/Y�֥�#��u��C��	���P3p�˥�(2<�k_	�B��m`C���B�D�\�$ٖ6���9�a+�P:[
���1���KPE�54>٤����t2��Ѫ8T�'�@V��)��	L�%>dF٭ňMKs��u��F���/al�����/M5�m�J����A
���UO�c�-T��ECR�v]�X�"&n�?b����?���津c�Qs��>��RȊxN��6�ʧl�3S�NxȔAz�g��"��Huj��z+�d�pU;�lp��4�s �,�u5�j��\j4ߦ�koz��%�fzX$�!~�� ��I�yoI��iъ��fi�mr@��P��જ������*W�����:q�����]I�%�f\�/S�0���˚�[�$�PBp�IJ��r8>o�]�!��R����* ��F@X_]綘o�ri�$�z��
�)r2��W`�@ L�;�h����*DՍ1r��F��B�p�����i�-dlo��ӟ�����p!�S;��cZt���ñ��YJ����RsI��l]��57��u�m�`ڥ�=�H �Ge�
u���iC�1Ć复�Ԓ��<;ГV�N�?��,=��̾�ynTS�`���௿J�$���\_M�5E5T%���4���Krq!背+����Y�����C��*QO�z%7[R����/!	؞�q����_��W[�+�����'�/l*�@�{�e��8��9�|������Fp6R*���'��/W`1@�w��~4.f
^�W�:Kvj�t��F�+�kZ��9d�l㻥z(m	�(
�i�U�f������Lx>��.�%�p[�B��_m���� �c�S�^��\�� ���XE�UT������Q�`W��^�i�P���A�
�3�3�gVS��C?<���7A@
���aXˡu�uc䯱��T��*=�pl��Y9�2)�����A�%;���Ih�'�K�#@�G	�Y��('�zas�䛑��7�Bõ�X�X.��Z�̽ϊ���p��q�V)�j�(J"�B��*�>��_ܧ�Fb��KmV���!:H)�^���(,Yv�/U��4�kϽ��:|FB��G��z�	T�?��3���)�������~���k���&9�� �?PA�gh��Lt*y%�
܁�[��9f�{t�Q�ډ-к}V��K:XKF�aS��^�t�j�n����lR
X��"�-�J�BⳘ?sP�7۰��H�E�g
�.�q2t/����v�c��G����w�Lbջ�����F˞h.i�M��:�}t�t����\6(C�ğ�����d�q��K�f�r��1f�S�ثӨ}4�0�	_ $d�t�����UB��$��"�!��htK-TY�� �=0�)?�e��ᗿ�8c^�+��O���JDhe�Q�~�
K5<�J�Z,��&������ǥ�(jZ6"�/�.�חj�%�UJ޴q�B��Ȍ&7��l<������{���D=O�F+N��mI�e��@j��f���ۼ�����/�<wKko�^��X�Ruy	-��يC��m�\:c�2�C7��~���0��~a��	��dH~���/YF�Z� <J
BI]2`������~�&{�'��}�
_j����r�g�K�aoo ����1֊��}��EM}P�d,I`����� �(۳$�YG���x���5"�0�*��ܗ^���2��A/�>������gh��wchO��Z�i��F�p8�F�{'C����Q=!"�WY�Xk�OT�;l�� ���1S���Î��N���ťkTmD[����	W݂6齆-���i�`d����-��|�O�y@�l�S� �EV\6Q߇��S �,�z�Z�B�$<�3�(�u���߼���������c�E��E���=�w<o��`5��*:������~��*n����2�g�zA2�y�	R� [H��w)XE�JF�,���Ic�NkD�o�9(}č��E���u�e�'�C���#�`E;��s������{i!z���<$����7�~����BY�W=O�$�e� 5wK�{��Rቤ&�+#Ay>[;�e=� U��8�X�HZ�lC�G��b�Q/�Kͥ����.K8���v�:�����)d������Xl��T�-}�+�'�ދ��v�5����
Cv�/��*�)Fn�^�%�.��Ѐ��u�:�����4�8�*���>T�v�n#Yfɂ���7�M�@��"�#��U��)\�+}��{��jҳ�}��`��nn�.5}2b�2y�"���ؓ�G�3 2�ZRHJ��8���g8a��g~	;c�85�/J�)w�)����p�{��Z>�G}Z��i��Z���R͜�c(%�jJW�Nd�6������<��YpB�E��O jZ��ëp;8彽��!Q���)0���8�(@���ʅ�^��B<��Fg��}Ñ�9�ؿ�N��n��%�5� �󟁏a.J�-�%� m��]D�|�$�i�&	�)�;	]�I��*�C�⬾��I(�=�߷}��O}5Ҭ�3�&�]2�<���-^�c�:�%�O1.�j��Fv�.n[3�sZ/�LI�G�p ��T�Z���^���5f�t��L��!.W���af�pg��AB�ɣi<8AUz60Mp���~]X�F�nI!��f���k�%%��+��
��٢�T���D!��^��QTM�y��k�?���'�������]D���5���BjWL? ^�֟�{�ޙ:- !|: ��H3S�Ѡ��E
@ȸ�v!;7��8̮������,q-�Z{�8p�Otg��eAﷱ_�Y�l��p#-�}��7���:����@��/	�<
��I��Pm�J�~�ٹĹ�E�|�PMՔ�e؎���B���7���ǣ�û'�������q��V���8Hɗ�����7�j�����&���b�R�A�_1���=!^1���Wlfx1%S^M���H+J_
�A/�^���ָq� �s@{l��~���YD?G�=yuhݍ��iQt��	�k���D<��e F7�m��Ei%��8�&�j]�%-֬G�@(�i�XF�3Y��fi����'V�Д���O��X���1U�p��W9�y�����f��b���P�)�����n�(ZC�.�&�S�j{�ne�;� O!�>W��!��*Ez/� �!�9���]�v�����]N%����r��U痻���B���N-�8�Kc�U܆8��D�����Ɠޣ9=넒���x�?_͖WP���YI��0�������ϩ�u�MO(�8FEB���ٱ̂JxX�e���\
>�T��]E`����~�C��f�|�k���N�S�-�������ߢg<���V"���X�w��Ŕ@m�p|-�6*V
�ֻ|��^��`P6V�L���Qh���&�� Q�
*h� ��6��Z��g��{�K=��e�>X3de����r�@���㻟�S��+�E���v����j@�8��7�Q�;����~y�L��CH�W5�͉'6�����e/m�N��+f�� 6`�H�k��zg���{CC��S��Ǐ���O����L>sU������)��8'ׅ`���=9%�0���hWtJ�κ$Y�ԪVU+Pb��xp�,�t�w�1��
�Λ��ZKK>[Pس�b��CQ��	I$*��q��2I��{H^4��cM�wLǢ��"`S���{�P2OV{M�c冿��	}��;�Ž��>\�2h9�����jR�^�X���
���C����W'���p������Z�{R�7$�q@C��vT]?�|)�蒛�/M�~���'Q��&�{:56�h��)�fo� ��h7���K��L�ڝE�g(��T-ͦmR�$I/�I�$�پ|w
w8:a��"Zh��41Ғ �{0e�W������B����>�S^�(Y����`8׮�y�3������r��0/7~��~�˶;}n�Km.����gyD�K��4�=�n�u��opt�Sv_���@�2�"�q��T��~\d=q���[xE%5`jy��Vnآw�x���?R��i�uRHs�CV�����`u�+������]�k9��J��ݨ,���m
ܧ��g��d2v�0u��Z�-V{�7�z?.cQ� 0��cfM�sk����'��8A���8��u�[�l(�i��`�򋮞�Ȕ,뺖&��2�-���U΁Y��X)v�ǥ��/�fO"&�8���[�U�Rl�4
�V��c/�O��1���a���6�OVF�`i���i,��<��Ⱥ�ڞ�Q�L!t#|��aE�P��7��r��i�*���� !*��(����%P� �W�rx��H&��P��m�I*H:@�v?RK�G��gYo�x1�@*s�� Z#��mg�>E5GE�q�� ����'�SR��s莨]�l1�v*v�S�4\���yX����e�����[[�_3nc ����bd��ڰ�y���V�KT�
M ��cc4Wȃ������h:M�Fc�K��gt!n�I�v��0�)o�0v���|�����ƥGO���z�'ހs�-xu�$W%� ��z!�h����Ey���f���v�<��!Na���|!xT��Ca�R���윺Ex���}��~�Gd��q�P��J��w�l^�/�!z��}^B$x�L����R(j�{�"�T1p�;���X]pnic@:�c�|.NI�VGP5L��:V9�f������DIE�Ɨ���>6�Uw�ZK�G���¤���[���@��E�zDU������Ƶ7��H�s:bOSdڏ��{_�!����uW����<j+�Ɩ�W{I�i2B_�K�q�|�$�f�s��.�T�ӻN�'���N�o��#b�K��h_��AI�U���}ן��\L�
�,��:e{x��Ro���+K��5��VK������F�5=���hr8\qW���{՟c��`�
�mp��_�f�`���z}������]ɧ���kA�@�����k�L�]I5��R��~q�q�5�$RE�7��F-�ސf	�[��$.c/�	+v�Ͻ��5�ɲ�ei��Ł�BdqN��I���
\������� K`s��L���ܩS��ˀ5�x̤@��ޖ���/��wj�O$e-NI@��J��՟�Sdx��%��x C��~KwMp�SC3W���z��*��P�ː�ը,�,�
�z 0���M�"����3�v}�E�]4���X-� ��xFQ�TҪ��c˕���M����;�:F6�K�nD�Nβ����p���ܒ��h,����:k���r�i��2Vlf�8h��Vd��IS�g�`5�B� ���J�aS܆4�^�q��\nFe�-�R�R=�_N=��T�)I㴜cnT��H1�(	?���VBo���Ǝn5�!�"�b�.�&��^���ZBy���xi	`+ߩt�~pa2�C�l�³�2`��őz��)��?�����R?)6���%�`��"�l�ڎհR0���O�Q����gn�T5�]���ŋ�A���u��E�P������x4�N�ɼ�'{��n���7��wF����>�,��J� ߍ�u�j%��czڗ����|M���S���KW����l�C��H��|*�v��w�;�8$F����i����.� x����;�r�I?)�2<FӦ�~I�)$~*WCX�T^J�]yŠ��Ny���2��
����B#!8׵~.B?X����2f�3{Sf9����F��*<�<�G�$�b�	�(�2s����փ���F�z�&wE��YfTv��I\D���垙 ����+�I�5��-�3��N�_� W�^�P�p��8r�U�>��7+/u� dp/�Ҳǧ?����:0�0�	�z���ØN.��Gs^�W�?��S�VR~
4ҏN^���p��W$�uNh�zV
u� �mk�_"%�Z�Jz�ۇ�j��T�ΟS����D��>-�'n!.
��K� '����RuQ����P����Y�fp��h�k��]|�ck�T~OH2	#��bj(ZÒ2��-T��� �����1B�۷�7�q�Ӭ��+�`zj1
r/�_3�՗\���Z����={��]i��Ӳ ��ޒ���(���b�)I82u3��y
�>�9��gH�Z�Z���IZ���*-G����K኶�	pw2���i�(ti=BH� ��ލ�!�hl�D[�afe�[r��/�f��T���I��u�r���5͞�+M����tY�@�|���[�U���#د�p,�ᬫ"m�/�I��?y�C��$�T�1������C��9w.�iT).�����=##M�#�d`�,����L�W�G�}��!Hb�Z�I��޻BQS�M��4
_�����1��I��^����_�_9o�'�r��2�2��b�КR.p���Khh��]`�bx�w�s��`���F�p�T�dW�.Z��t�����§mP{/}�Z.?M�.}��P*�n�H�LX�j)�4�R%�g�~�O����j.V;<��'Y�&Gʡqn�=ѯ]1ʺ���p���I-��4u/��<Yy`J�G� �f���=	>N��gjj�Y��M���@�籉^�1N�to���B�\�'�����[��zr�h1�WN��	Oӄ��U�s%���{�Q
�zөN����J��B�Y
��Y�5K��`z+���{�9�䙬|����� ����5�+^�Cv��'ʺXa�-�.�S �� �\�U] ���4��c��Rue����Si�/O�EdR�0�P��=�b�aԱ����X�?sQ[���	EL9*�e>X�&r!Q�1g�_ +����mܓ��/���W:Z�ș������n!��,dV���_C04��iv�%w�'��³��6(8K%5��n��{E�ftx�}���7?7{7�7�Lg9��� @���E2�$���#�jTFr�L���=��r��h$L��xBl�6k�Ў{���axC!,jy|g�P�������iۀ�X���D�>��pq�EWZ�\�J�c�c�rM�0].���>��T�9�ߦ��+����#��_3�����:{l4|�EwZp�G;�dM����X��O��H������#�Q����P�Lm�|��%�f�v���}>h
%���ɟ&���|H?������k�S^Fx��B����@������:����竳�#��v ?�4�b;�As�͟Aؠ��u�%����u;_�?)�H%��e���)��a;й���;A�Z۰!圭̅z��w�>nJZ��*�#Q@�݀�%�{e�(z�`�1됯�S��֢0�ͥ9��%��@�����t����O�Hwh��s��RWC{Q�l�bL�.��bj�Ͳ��g��AW������A�"I�b�!ґTB5���d�P�����Z��s�(�l�V�X���_RGGD�}����[t�mr��fPVִ�3)E\�$�n9����j���@g�SzHf��f��(K�w��j���Іj��E#�Co	��z_���7'�����i/�j��G�Wa�<��͚Q,�������Z-�P�K8R-oex�d���À�:U�-��������D{H��\�d���Ǹݬ�̞�S�c�:�%���M�A�M������B��  �m�զm�&. �Z��(#oYw'	m�h�a���;��r�;9vтym��*9�I���O�;�Mi����^t�2�x|�D���#��$'�������\��+��_�k�,�:w_ɛq��ϝ;�|�F��tnb-�[ϕ����!�v�v}�FL��P��������ׄ���q�_��c�jdo�~Ǒr���Sڼ�-�NO_�Fg��,�,���a�m��U-f��{��~��0e�Ͼ��y!9y�y�H^�-�b�N����';�Z�[#]��{71J��Y�c��؉7[M��Sj�-��k���'A�L�ʴߺ��.'�Tv8>���j�.z�VH|�-SSΆ�۱&{t,,,2}Տ��<qTi�]ª�b��2`r4c��:�Zb�K�߳�dT���ڢ���|>"j1ÚD5-6�4ƒ�x���q{���ټ�&��E�4�4��)��fd�O-��h�_،�W?lSf)�eU��(>+�${�	rŷW�q��x��g8ٰ~�$������e����z���s���mX3H�a�>Z�q�=�ّ9m�����CF��ٿ|�{�tS*��C^�0��e�Q��4U�Ej
��L˟��O�e���_n@�,�
*�,�Lq�Q�0���2᫈�,)M�ٵTn���GF�d�h@cN��,���#���Ky����OWV��8$lO�1z��[��.�Q�r���N^$�&����-s�6)����:�yfrA�k�9��n��n�W��T�����QM�:$+jd9j��F3��2�=�":Z
�z��}c]�G�NM+U�C�}�p��=�'�1�ְ���� (5.ʉu,��)�ǿ����&tٹ���D���o��/b�r�>Ca��dX��l3�%�O�C��A���Scߛ[�[�$ފ���"��l��ȃ&/��Uy���Mb��*U�}�U���.�9.����Tٱ� �V�s�>EG�*�PT0*؃�{�X�A��Zwq��+-��P0-	A�*�o0�M�	+cVĿ��C7%~�\�G��L{h$[������Y�t�xh�o�/;��t�ȑ�<Ԭ��=���Z�?W��D�>�)h^��u{&��*(�z�����^������ӗ���#M��e���� �.�@]�������B�
v��y�Cr�yi�v��!���(1�I��}��)���P�~�"���~�|<Ap���L̈́�u`W���
+;�S����2t7����r%l�Է��!���&���̎�G�~�oQr��aj�o��#�\{w�?;R{ �5Ji���6�{�߈��8�x�E��Z@m3	$�3��h�@Р� �!�����yM�����f���ؿv��p�<�(l�s���bǖ�� �"|%�3[�Y�EΟ���%0����n�)vF 6����tw�7z���6|>kge�
ʲ6|�� [M|Rv���fX���.���s/�ѺrB��:������d�V]�U�YI���^��g&��&�q�a�J�\�A�V�t3��k�e!�$a�-����w�ɘ�H�)�p��k�A��Pg��X.�T82ًݝ�d���q��$��o���]4.�%w����k�z���y-���ڹ���O�J�^�`�����L M�w|�X���v�A9a�����Mq��y�e%��M&m��'����@eWH��a��'+������)�./�ƙJt=N7�:i~z}�G�^�,DE*�K�-f��?>	�2| ��\�'{ɘ]M��?`�ŇQ���hԽ����س��c�D�
Pɩ�7P.8�
�Q?��T<�~����g��2���\��3Mu?;v|�X3{��Qf���|N�?O�VJ���vzD��B�`��1� �i?G��.&� E�,����T�Pԧ5��xL�1=�����R��p'���E�����B� �Y��\�i�d�QH��������D�)�\�YE1��X�����|�X�l����I��,:�u�0��1��fJ�/0@`��]���wG�/B��C��l<6lᤝc���W�s<��S����3�㡹�����t(�C<Џժ��i����o,��g�r�һ.TL@�R�~OF�<Gcs1��������@���K���,������_7��?XTK�Nl�&���h:W��m����.�S���E�c��L踐�Ȃ}�jq��D�߱7���nu�Q*���|'qO��iX���P���rUG$3f�qh����˺nO<�hֶ���<��"��J}%㯓2Ù@١�������s�_Up�ȳ6u蕕���C�h(�0� �$��>��f�/l�u���=��o�[N��;i�. ����:���^�y��5�6:7�ks��?��/�>��o� J�g�B�v�]��%7X��O��܋����P�y�)�i�� ;{n����>�
I��L\9����l��&��lܻ^G;XS�p�HȾ-ld}��C����f-[�:PMiը��2LD�����s!Xä"B<���o����\m�4T�����8W�,~����r��@��R���n���tz}�vy��:�����io����*���{3���r+�R�w}��#N����� ��"�;��n0?�﫧�:�J�019�֔��5��?���9��3���8�;_��f�,�-�2�8�1���Q�z�Ӽj�;��fuh�5qu��v���hx�_ �1_=�3&���9i���ᛔQ���m�?\_�k�x$NMS�sRE �����C���	5�7�.��	�,�a�/p!��ýlb�N���>��,8�����r@,3/�$~yt�li<1D�!&I���1�Ed�.��r?�d{X��OI�8�y�)D��H�JDN6���3�c�������;�����׮X�/)[���3�Y������N�џ���Z���X,}s�=��lRdK�a�nmԥ^���g�P��l�kZ��MS��h�ZL^6[P��Zj �) ��u�o�� Yz�)�`m���I����+$+HG0@�A�djA0~���P+�ʺ��vz���}XqS���-���:�N�9����w��������K4����T�t�T�`�\�D�;�DAL��vIYH�M�+RkPF+��;�m3�W!�����!�xO�fY��63�s���"+De���N�:y��a�vDb�׻>����UN�O`VG�f
Բ����=�f*;�Dp��
|cB喹����qSWQW�D���5�'�9�]U,��S%~g��UfH};��kښ�����+����wYfSOB��Pw���,m% �i(ųwЫJ"��-MZ��y& �[/�!�xw-����_�l5�4�>|-��=Z�A��C;�}=t� b8e����;��d4~}+����Wh����Ɛ�]�}iϢ����V����e�֡x�[:�.�0����^�S����j�ژ��p��fx�c���z���D��������U�9�TH>E90,QL�؉�t.c�jG�#yW���4������C=�R2�K�?7�TF�h������_˒9XXd��!�]׿����c"�;HED�VFζ�*������/VW��.$�yU��;W��?v�uTe�HӍ������9���'�� =��2��W#����ez��g�Z3�]���lX&��H��l�����z��`�ŀ�/^��)��qY8l.�KJ���0oݪA;�a-��o�XC�.�sFu��:���� G�M�6�]N}�޿��O���RE��A�K�<�n����Q���j��Uh<�#�v�aN�iO���k�C@�N<.�[⋇��O�{�`X�y��
�^��^�+�
��f����T�2V�7��9�m=�s�	M��5�n@�pQ��n1ڋ�M���l.��g6�
Q�g�M���6���u�Q�-�#x��J<D��2���� �S�//l/X'�j)�Z������<2�m���Z�N~O0��~���Se���Ċ�l!��9|��;��G�+P�G��"m�ĺo��%�
�x�f��&�����:n"��ߩ����L:��Ԇ%��R|�`��v�`�i�����
R��nG��*��s�R���V�TLA���uIN!%�s�<�k%Ხ��аXI<5�e�~�ȕ���)��{i���ʌs�㆞��/eE��jG�x��*?�4_�T��7�}cs�"J�r��2$4�e����-#���!�7�9+��_p9�ޱ�
�C���K̨�bEϫ����W���[�e#a�${@3?�n�i�U�Di&%9jf�H���i��Zя��"1�/sݞn�)멬��xz#���K��f��͜�����qI�|���?�s0��}��)"�������&����m��)xd�0����Q��y�|L�#)�ɡZ�t�o��<���F�L:Q� �g]�,{ڒ.� ��6r��U�seЙ��dyv`�[�9r�7սs.`��gL��ɽ��˪�+����vZ,6k�$4F���L����D���"1oq�U �b���o����n��pn}ah���	�F���~26�������c?شDb3vs⳾���7kdn:�ِV��\��iC�����T#���y�U���8�k���J0m*b~��J�
��W�laC??y�퉡t%"e����N��U�w݀�4�*,�%e;�r�����M3��S�"�����+2ԫ�a΂��.��X�K�{�P�t����vz��"{{P~�,/ o(���Ja���7+%����tdr
�[��qGO�)�?�Z r/֑g�����s��q����[a��ښ�����&$F���B�:�M��Y�?���o���>yoc�e��^�j��"`]o�����}w�|Q��aV�L�3�i0Me�u!���fUT���K�(���7�ھy�Ж�QS�����8"M�w��t��Bi���Y2�TT�ݚ��ië�M ~D3|�G��?���q�z�f�<
�s�4���<��`AS�I ky����w�l&k*�QG_�W�����6C%�2����+f�T�/ԥ����@�t�g�7\qՙ��j��8�4�k�-tm��C��Hn���!��-��c� �`�vo�xI=�b�%�ö�`ߢ�u�m��h��?X<.Q,ڋj~�=���C		�� b�8��ˈ{�7�(�V�߇�������!c�)�1��.��G2�^��/��f�7��\;��ݺشw�Ff���k1�a�����`���1�j�>�tX�����H��IX�&��bFĠ]껙	��em�	�Y:�o�B�TT;+*�z���-�+�dQ8�ug�fL�ϯ }w̴[�Z�:��"U"���ϵhb��l3���]E��3�nyZ�~�v���ow������U��"ϼe�'�?���f��q�P��f�`XP\�ls������z�,ք8���~_im"^�8���X��NK��\}P�k-�7]�߈ ^td�ؤ�Q �×��rYz�`g�ٗPf�9d=[�bC����j��\)��|xR����jj�+�a~�@���d�m>��3��-��.<�>)�N%Ed�6�B�ߝ"N�$^8���?��ȡ�Hx.�E2�i�Nؽ�*��T��l��d�����3�؟D!�lj쮓�ﯤ'ӣI����6o����]_+�����7�B��xE�+ǣ?:C��J�m���-xoΰ뿼/~;���p81�+3=�i]�%QR&h���ֺ͐�.K詝�2ܣ���q��A�'h�Fq���2R��6r5��"$ o*��BVA\�L���)�<�ʱ�Q�((�_b�b��q�5R���}v��j�����S�:2�NL��|W��mm(��^ԬJ��4.��9�u�H-�GJ	.į�Ƌ-2��g���v$�3o�:����ٰ�C����  �&�7f���@�9^e�5XA� �R��!�s�����ҩ�p��~��Z���4�	o�(I��v�d�6�e�1Z�R�����ܓ�M�8Fm�v
�6�N	ݫ�癣'�����lz���1&wEY	fg�V9���<M	sT�䦑X�ۡϜ�f�R������!}T�;հϜ�̄%��2D-���d9�B��K��m>p	xqJJ���~��)��Qg��\6�UЦn�"g���QY�K�UA:��%��Z�UB�˃`Ec�MMSd���B����L5� ��윕ʤToyIsI_��%���;c)K檺Z��z�8^�L�Ѻ������1���#�e<��5xA�d�������)v�`�n-lƲ��T ��R�NgP	�:KǬ,�K�ͺf�S�M���ё�{���9�� ����q��
ͯ=������J}!4���'��;�y��o�ê0Փ6��04$ X�a�(��KPqBy��|�|�@e�'��5'(�r�h��|];Qu�c)�j��N^�?���gm�aW���f�)��,�L���aW��S��0)�#qc�6�
}|�i�:�@K����AΜ�L�7�Ic�
D�>?�|5�PdKʆ��u^�ڡ)��N��� LV���A&3��)�Y-�����!�&߭%��yr��D��5nۍ� �b��o͕�k�g�,P�zc�є�ҥ/,����B���D+8��Ηq�x�Y���P8�/�λP����'7ꛉ�n��#D�}0�C+��}��'�{�4�����P�����෇�Ş�B��D�or
`|��8�_TY��[x;]�G@�G�kE��0�+�p��T�[�օ���a�E[���P�+���*	V��K�J/̀ÞzAl��x�q��D�(+p^�
��ߟi��䪱Ƥ}�LN�g���`�o]��q�9� 	�fz>kN\!��=N�.�7��@�ɣ�g�	���r�f_�hkiaq��9�.�YMr��a�$p�ǁA�,�D��<68+L2[8�m֧\�&A䈝��N�-KA9�%�q�)�!���������8FwF��_����i�Nt���I����(&W�+�FL�%���c�D�a�B�3�/�,pG���qx���K�DR��fp�cDw��-j2���v��ܠ{d�M�g��p��`G��zo'�Uq���F낤65Μ�6�.[C�C�?�Г*�Zi��u�X"�5��s�|Bc���X�z����+X����[>�ro��qQ�_ݠ~]68!�Ū���*e�D��Wr���H=�+��x:�qP�F�*E�e 	JƎ� nd��ľ�x�\܌��%�F<��m(TM��s!�m�`��OVO�hl��K��;в��ڽY�V��1r��v1K�^鋼l�~���0*^�Q3��XT�55�
�����ά��
"L��9��1�6��"eC���'i�"=E*���u8oB
/f�E.B�W�*��f�|�HU���E��:�o�A�C�ߔ~�	J�#��HUr6�$��G�H�A�B�.k�?�z��=C�R@2� ��0mo����h�����&B)���7���Z�.Z����<v���#y��7����������S�S���X�Pά��i�^C)������Ӧ<����\$�3)�?:�J���c���UB<>m*偔y�<T��xR)on��(�����-����hW+6�9�D�s���j�K!���u�	��d��7y�k���#+�OH ���P����& w�Ըx�s�J�%7�8�Œ{���;�8'-�۷?�ٹ���4.�)�3�|2�����'}%,6��_�Fu�'��s��?y�/�gTP�=��bb�B���d�ٓ�.r!֋;����vb���
���7�L��S;Ld�q��6�2Ƒ�� -
�<5UJU�4Yy���T6�(�Ɨi\��`�0%nou��)Ql�È)rqb�|_�\-g�5�ߓͲ�>��:��#�s�5r{2⚰���b�@U2p櫿ܢ0ͅݾ��H����x m\Vƙd<�wi�C�*�.����g��
x��T;HDo�az�Cpz���a-	�r�8��;��"�	�y$��*��{��&{� ����Z���b.�3S,� hx_V�Ge�2�p�:��V����6z��!�?����;�^�Tx��s���ڌ
��@��'ѣ-�2�f�����������N�t��AV/���O\��2�SbM��ͯ{/5[���;�K�YZh�о��o�&ݻLl�u%I�f�����t[�%]��>~$"��-��ϐ����#ֶ�	�y�"2S��������@_�s�T�ؾ�5Z{�?���
��]��
-H���E9�EI�m���'�59�� �S!�r�6�u�떰Ou��<A/	 ��^a��kgv�*�~��M��=�Z���^��� ����L3�Ǹ
�ԢD��Yy��Z�\�/Ͻ_�	0.j�!�[��I}JZ����J��3%�@��. ��df��T;+>���"1�����(�x�_�EiY�V���g��q�b�:t��D��S£�8�q�;{7�sZ�{"�Q��!��YU'�3����m ��v�yS/ة4����b�IL�I�i���ϳ�=?}V8�fᶾ��T�AW,3@�;{tG�f�f���y���ФX���I�%۩�?&���ٛt�'��\�ec�U����hYH�)Y�����G�2$!|�Ft�)�J0 ��o&ϺmoR�G;4����`� 3uq�H�S<)��?`�3%P5�])�f�3��} �n=�y�5����"�Ar��z�ކ`�?s�N�.�.�t^���6�9�uBڭ�؊=��Q�adbp�/�;+[��
��%H��e+����v, j!»8Z`���8%׷��ώ'��pef�d��Wɾ�H�X�
�#���ZM٢e�Tw S��^�<��($��l1���J�8��aPߒ���\�Z[=	͕ U�pP�r�m҂��t�0���c�ku�R�SwU��|��-��{�L?Ϳ �D�����fIzB��w�v�=�)gbT7�I>D�o=��,I`V���hk�#⩴WxXtGm��)��e��MH��! ��➭g�h���9K�8�7�m�f^���9�e�� �v~�O�l�b��w�wZ}�}��9�&��������X��9k�n��P��hY�!9�>u=�3��+�e���}Ms_�_
b݊�]\dk4 �m�� X#�f0�àJ��	���)b�칡/�0�/���"����>,�:$��|���v���4���O%D�_"f�"�>���({��N77�Ζ���&�d!º���z~���<{��^�C����%��q��U � A�z|(�%�m=�!�\��K�#�Zl���	����{�l	ӗY�N6@��w����-�46hڭ�Gyu?�<�n�Aq����Q��t=��k��_��6�����}�CX��h?��-Qҙ��
�j��}��Q/���G����u
>�g#V��EA-X�b��aH��(?�vb��R!��w8T�o}���P)�74����2�i�޽�F�?����<��r�N����@4�^���Vן�;���Z:L��F'�+��,~h�j�ڬ^L��R"�We5�X��:��]�Hrs��p�d	��;�51��u�q[.�su��=X{E�z��2������(uO1SS2ǌSNd9�X��Np_s�.H�v��P֢��2���[�����2�MTX�j1��o}��R!�.�� 4�q�mq+�w3'B����.K)��3O����7kc`>��*�̤�3dD(d�>��!;��T�ڍ�gK�݅�+�6(I4Q#Fo����#�{[<�w������B��h�U��Pٸj%b��(�t�n�7	W�8e���{I���P��' $��7�_:(r&�IB-��]�a���P��ܬ\�炴��"�4�;�����T0OH��,^��%���x_W!�7�������K��!u�w�f�ý�ź�9���A��V���Y#vw�Uj1�z�x&��5BmA`�n��7���w(�Y��c��{&R��<����%���*�Z��<i�Y�����������5���e�C����d�/�s���B�=z!�d��hYy�phn�_t��5�~���s9�[3uKp<��������p�~.p��u8�>$���.4_v��E��>#���آ��?�pt�o� ekfe#�}&�'�u�^
����i-�#W���"����7/19�8�׫)���-KtR,�Θ�$�3��4蠹|���ߔ��p�ΤAT��87���De��d��LTb�����"��E���a��������E$��#=�&L�)�>t����dND��flLX��2�d�KҚL���D �9+u"��񰽥7�m�(J���i�ư����p���k7�j����a;�LN{'u���"���N���(6��P��,���<��=�O4�u������
��Μ���4��]� ���L����B���c���c���=f�Ɖ3�U��t�o�4��ǻ8�Jp���xl&�d��T�O�GR���ڨN���c�&H�t�������Ț�3� ���E0K�e�EO��`db���hݹg�dS(�M�k��]%�9"�d�f½������2Pm�P-h4����Ɲ^S������Ī�a�YĚzl�0$bQ��E/����[ƥ��,�fg�� "y%��ds���g�#�9n��ay�2W�u�#2�����@��QmU2�D#h)���̯�$�G����Yܥ<����S�"D?���-p!�F��UƤ���'g�B4�8�z�1��WyҁF�&��*���a�E��LƁ��W�V>�!�t����
��V�;aU�Oy_{8�
 ��P�rj�l���(H,-G_�B��hJm��&O�ʊ�Љ0N^��/1C#��ҫ1V7c*��@G=�!�袰| m���9v��{�VLQ�K���N�q6����.��\��a��
��Q��n�F���P姶/��M�Ν/7����v�=����[�s����/��M��80ob~�\0\"O�����L'���R�V~o��\��系����#�	�q{}bp���-"�$َo��Ya��̘d�ʃ��,����خ�#�5��j�_x=
)[>�Yk�$��/���ѨƖ~b��1D��O���A�H�{^�鮮ъH��53��{},x����Qq���J�~�y֯<�mưd0aH��!K?$�I�z�7ˣ���-:T�H���y�1�ʜ:�K)z�#GӻSV��&�\ZX#������ꡟ��Һ�幘Ʉۡ2���ۃ�؎eJ��xj�Dcl�v��yՂ�ЉVj>�;B�������}1��jJ��\C��r�{CW�:����H���X/{��=si�O���z���t3G�
�����wݷ�@��C<���f� ��r�ҫ�U���ֺ��C�y�Ӎ*�I2d�n��C�k�;�<� 2�V�������2M�3�%+��K-��
��X�,����5�c�e��0�\2�&iZ��ъ�:��H@�-T)��n9-ay���D������گ���2���X�<��|L�^����-K�V�����6�)�hgoDYR�����o֥���AĔV� �tf�q�e�g�N ��Q��ݠ���[���o�!��5�-�EK���o%?dJ�#$a��ذ�x���,�J�w8ɯ�P����p��K�K�4`M�
 �[ Q�k�%f�jׁ�u�J���}3���
�Ȇ&BXp��Rv���5o���Ӱ5��v��(�#��D%<�QwE���a5�s��O}���,��W&�����m+.l����D�Ч����2W�`�}�	���N؊MZI|@<|t��"�T�=��Ʒ�潮Ƭbv�Y��je�Ȉ���Zn跋���|� -܏�]�KK�x�*A�at�t��X�K��&�d����� kze?���8}s��kK�U����d"|�d��><�����cG-�~s����s`=ļ����(Pz�\�h�쿼W�WT
;N��&S/�X`��{h�r�W�ZF}ym$xg�F��J�M�%r�iL��,ȕ0��W9�l,p�w��H�zζH�f�EEs��k�u >��ޤ�Q��I���8��m�9%�����S���ذXY�^Rs�Y��<L�G<����zzHt�5�IrQbQ~�X��#Ƈ��:"���QM袖�c^-9H
ɧ3����n�<"�=�/!Gx:x�/��ٚZn�e�K_im<#Y�]xE�.)Cپ��ʐ�w��QD�	R�c����oơBbfQ��������8n�@�jY4���{��&M�ᔡ��z�����R�]��X�1��M��q �|s�������1�`��#�a����=ZP�9pRа������M��ڛ7�r$� �Y�fX�(��'��\��3|�zs8��4������/��ؼ�L�d3�1^U]���ۆ�E��<���
�e���hw�rX�������Ս�j������P���*�,x�=G�WU������)�mV"���.�����nY�Ӂ��
���)G��ݩ9,��d�]�!ʲ;��jBU����I2��W��N�|&8��}�{Iн����cIcV@n �3��i�1�P�}%����O��]�J�����e
+�O6]�{�	���8 �Yv���b�Y4���TV�%�%�9��ޞ�C�Ô��9\�^٥�m�;�	f]>Ga����\tq!7�WQ#]p��9/�D'����3bF�E���GvY����i��A�dV��_��H�5i�b�<�!�"�%�w^k�+�QjVҍ�U�	4⧺{sa��n���8��23K�C����}�@;Q�����?C��8�L7���~�^�9	�y�>��i����M	\����/jL���Fw�s�-/}��o�*��^�ۅ]��I�~�+^���6@]���N`�^��Fݍ��rZ���
&�	3u��.��Xs�\-���W��B��Z�i�b`��5r���!�D�0�zMSB�I�ǺUE�e/�k),�Q̟�K7̇_9+:7�n]�o��?�n����|Z��>�4����߉�Y�Ɂ��'l	��>iUf�[9Ҍ~����;>&�d�� |;񻝉�5��o�[�gX�&�P��Mڙ���YmX�+(�YY�_B]��dmS��iU���*�W�e�.c��JP��D�����J����F�Gt���'����]�`���4����Jٷ���/2�<���d�ݰ�]&쑈��������*ŒtV;}<f���i�C����#��BeB��}��p����f|O�)�98@�U�[zs1�x��Rzm�sP�Bs
u�;K�P{+�r�\�W�k�/TA�Q���B����|/�"I�)8��N|z���o�αGۺ��
����C����6�!�Kr-x4?(�%]i���iVú�/��?���t@/��=b���8����q ����o[>�+߾��4.��/�Rѱ��W�}�������G3�K�%��jު�t{B揮ʼ�%����̋n0:�,��("��� ꡗڍB]�K�<�@p���r�!R:CB'Y%�@.e�i��'@�W��SA�
eS�.KK-�3�6�!��z��م� �Y��;��q�SU�@16�� Սh�=%Z�ʵ�w0 !b1���գ#͎�a�*��~�7`)l]T����	�8�V�7m~o�����w%W�����
��2SkhdҞ{a���{햗�ћ�.5��&��Vh��|����q�4
I���� ʋ��!Szɺ��Ǽn�u�/���~:��~��A�K9���y�c�m��kG�_e''�2���!��{�X�PCT�]�3/Z���� �f�HsRi0�A���J+��z1��ľ����W�����X3�8�ߙ�h����l�W�U'���y� v�d�ݵ��)
�F�*)j�-}�~���h�z!�o bW̩�[�o�88U���{�g.�@M�Cy�{5#-����A����(;n���z�~�M_%���ʱg��8� {���������8� ����S����l��$_qC���ـ��ó4���l�����+ڢ�6f5�ļ�0ڭ��F�
P�,Jg�z�������CO�<����9�������{Sv��|���^�t[^�8�?$T\��<�cT3����~#��������᚞��1��U�
(�u"��8�GS����v��Ū�%q�m��|�@\	�R^1��u/͝�zt2u|����!FFcy���u�܍�RѲ���[����5K�">:]>�*�A�ӹ6���	k���<U]�8�T4�S�4;���]��q9o-}^��f� T[����=~*��M��Dlz�[=I�n�w[& k����!�u�� �c����l"R���#����#J��6�;#1��+}`�r��@�ۼ>����wD3�''hԉ#q����{�ٸ[�AQ�%��j�ڈ��Wq[_�y@Y��t��	l!F_����ȇ���I�q����-w}��&��D�d�g�FUL5,�� �9]j'�0�R�v�F<	��[�S�%��Z�Q���H��g'�����TM��t��+�tZ�4{N�4&��P~T���ңi3Rh�9laB�9��O�b4]h�ǩ��� ���d��ĭ��o�B��q����A���z�fL�4ߎ�6,��xj�O�3Nv�wSX�$���	ϳ���Bd{Ϯξ�̙ݘ�����͚����R���˜�̼ �0"���aA��'��ym&LJ8U;M���`�4�~�*����eR2�G�P���?���?L<$���Pf���*v�T�Ǯ�CA�w׺9��<=#/m�s�r�~�����4���7rOk��փl⏟��iM���T+�K���<��c�-v���;��	4f��z��K�y�\�+�T�t��i�n\��i3�2�GM�_�(T��{�H���T�X�?GO��7�n�2�X�����������>pDw�h*B�-��BF�t豨7�~6\MW�
��)4k���2ڌ$����0��2���4���\��F����ƖL<��`xYX�n�pR�x���j]������q����I�iǡU�Y�24x����:{�se�T����Z��0 #���h���"9�^��!�ؾѡUڽ�b��*P��iGg