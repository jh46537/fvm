��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����i��;ݏ+��ↂ0�?�ceR
k�&��;T/�h��HKIw�|��&3.��Ů��p�!Q���i(�+��gX]����\G��/"�TDV
x; ��*���1$���'�os�G́�C2�:>�r��]�#A��]F�~?:6�,Ӱ������4;Y-�����|��U]�Ԝ���6&F,O���*Tkt�Zzڠ6]�ޢ5m�IS��Z䝤����VX��@)���t�I��Ml�k�{F^��-���2#��q릍@�BF(S��:�����jm�â.]"�	�i�,��Z��GU�՗��5�P�N���Lh�����	"���>�֞=]Kd����;�'��D�Yj���I��Kv���R�]���}
�jD�Kh-��W��M�� 	����eD��p���.��8�O���lD�Wa2]8)�b�;p![��5E���I6�����>FN�,5��y��zo�����f�_p)���P�Ey������0~$��^F<)أl�Ϥ��uvLi�9���~�Jh,|FZ�:�f�Q5@��-+��KP���IDu"(uB�LY���� �#�9RyD^oMw1��wS#ښ�p��G��a�u��V�Ρ��q�E��_�0���[[FX<'��ϧR��В� �'n��<�e�����C�J��	>����MX7�8��>ߩ�?���\6;������zb�ǝ��|b�;V��D�͵Kz��ŪO7G�ʕ���,̲W��/��N,z%s�`�?5�1E�tf�BZo�K
�=k��td!Q&X�m�PT�|=���H�?�6f�4�=�w�<Q+�١��F���"��o� i��^P��KǦ�S�es`���J��;��V��5���g�_d;��}��N~���v;NX8��&�2�S�%��o���}o�GXn�0y�Ж�;D�<��@�a�9�O$Ӣ��>$�U�'�/z�,��P�-F��:��l�3lb�APEW��ِ���ΒG�K�A-�3�P �e��+�l��;Y~���&��G�]��~&�L��slL4��t�>�>P��4��R�u��?
�o��1�d�⯅'�@-b����d+��Ǖ�L��m�@�� a�^��Ů��\C���x�J��M.���_�~9[>r�YjI��S���yՁ��H�AԹЬ���"p�X�ۀ�!�8q���M��~wE���::i��0IF�����k_`��������CM�Zv�\iǐV\v��-��U�9F�1X��/B��Q^Zm�6���bk���N�u��O���� .��O�83�M��Ay�Zi�V�0��Fo���	B^��)�����;�U���rx&� 
��d��0�m]aN����u�E�Hw�LY�`��o�.��g����Y��4L����;�ٴ��3q������%�UMf�LH��B���"i�0�	#��6h_V�x1�[Iu3%��p�C�1�c�N�C��T�=��6�ZL�1�_~B��c�Ӡ����ΫfFH�Yv*$;�s!�TB����0�e�@�H�R@~Q�t��ӣ�f^Un��Q���ǥ/��.�O��ɳX��b<���~:.K�f:aE�k��i������m�g���&eV���|�UD�4m��p�N�{��+��T�?hW2�*��6�rpv��P����Io�ʽ���v�q��7���4Qo����A�#�!<a���<��_�if�d�����]�Jf<���v�9/rԥ:��t�\�����p/֡�G��(�|�yu��=fQ�u���R�he%I>�,b}䎳Lgg�0C�mef���^�+u��ȟ���nFK�h����(O�a�fb2A=R�z��C����������$�����tK�Lu;7N{f����˗Wy�B���;�.~���D� �L�sE��[ �5%�ÿ%s�N�-��f�LyG��x;09A~]wN��c��5�!��3#��`�_�iĂ���������Y��KR�����C����&nD��G�My��p
WmbKz���,.W���0�&���E�z��s#ƚ�]+�T2	O�\nD�>��TZD#�ky*�p^�J���t��Ԍb72|�n�'��1��,��=�&b&�%���I����*J��3�;0IuL:R��ث��(�I�?lw�1�����J4����5�m-�?�+Ͷ�L�)1(�?I6=����&�K3B/Xi�h�$��Ȁ�h�3�Y���$��v�������u�(�M�XF8v	+�kJx�]Y�xCf@C[��^��Z~��r*���;�]��M`b��[����٢*��)H�˷T�
�mqV����Xwbȟ�m��f6H��'è~Y�u�����.�����x�p�(qw�KN�2#�	�����d�0���7�(���\���B�rU#O�w��&;6r�!�RRJ�~>yɪ1�i��Úy�})��s�B�,R��B��Љ�9��>�ԓ�{	,�%ÐŤ:�!�
q3r*R�1m=,�?����)��&Z��9�B`���E���E�KG��`�1G��W��p�0��Q_̔4x��ൈ����s�1�n��EV�a��6�u��'�5`�F��q���<D<�L�
����{%�[Uv>��������*�-�N�?.��<Y<�|�OH��J�1�F�7�]�ٖu(ټ	>n豚}x&���{>(�aIs]�5h����Ll��!��yC\��9�_U;ygE5!,a��6��P
4�qp���f1��Pk��-윓,ķ�M�1�~"�GW����lxdW���&�H�����}���$Qj���q/)p��4EPvV�m����mZM-j�:ES�
�-��3mN? o��9�>sr��\r���k��� �5^���/,<Iv�XGp�&m��w NU%lG�ն2<�[t_��d)n�����b������3%��\y�5x3D�R��;��5�����_�[�7m�$��7�Gk;(@2/�������&�w-�\i����/��WP�=���!M�P�	;�u~�6Qg��A�w�.����;�]%A�+��)�Vٝǂ�N�s����,��F�"��`Q�<c��ҥ�kq4%N�W��k�����}��d�����FD����Bt��q�r��4�?�*aʡX������!o������]��J��uӀt]>�S�s]!�z���c�^;j-����b����@���K^��0�4���k����Np��B�J�t��@6z��S��\��O� >����/h��=�����ਢ�t�d\ Ӑ+ƟK���ܸ�7�Z��w�j^+ڕ9��5�ӌ����S�74����6��Jx�h,�[H>���j)�[�"Qh����_�P����<���u�Z�EE?���q
O�Dk5)�ݜ�]�h^�6.jp��<�����W����"����8=�9���C����qD�s��F���nj�O1� �NJ���.��$��fw���鹢����ZUM�S�Nu��:�ܟ��t�H+�n��Z?�X����R���w2W�kU�'j��jU�d�CM�	��f\��k��7K��T�N��?�'f�)���]��s60p��YK��$�L�k�Dd&��*�CH�1�s� �x�>��y������R��.��=I�`����4����J�ن� It˂k��܌V�gt%��Q�@��r���7R�<R��a��*y���6<��C?�30��4�V�y�h�xF޲��d܋f[地���}��� �Uns������{v��!�L�I��KaK�wu)')Y�p|_��_Z�d&�f6#;�X}<�>uS�#C_�;�?����rЕ`j��续��'�q�);8<v|3���t�"�Z���~O��A1�kTc�'1#�UXTN��i��M��Ip�I������F�}�r����[�'���,ᥦF�N�4P�JƖX�C�X��j�w���Ȇ�`��-�mƅ�..0��A�8�i�����:9h��gb�oBꟗ�壖=����.��]ݲ�����X����:�5�c�9�>AA!���qM#AG�r!�����x�g��,Ch�ޚ�p���P��k���uo]D�^�[��#D��r��oW��~o<��1
�D�4~�B+�[�ZIqrz��b���2����l��c���uɚ�4t>�XI�r�t��]���ś��n��]����1v�c���-�N�D������d��I�4z��<��I��V�=�ay��,,�Ya�����z���ȁ"9 cP�: Y�����2��H���s�� p�у��l3IC(dǍq����� Z�:VY3ʥ�ujp�_Ȗ�����d�$9e�J*
0�����+e0#�[|k�f���Q��cn+���<��	���h5Đ�V|�q���K��=��n�,�o �w�5�%�X0Z5�]��bcI��$������(ǰ+cVG���F��}��
���)'�C*ZN	�sV�j��V\g�k'�����X�E ����e�1�f� `�����*5�c�|������G�?�9��J�{�͂�a((
��+0u
���d�p݁#Xe!�`�~��Q �ޟ[�*�Oe������P�l+ �3�������s����]�=�t,��"4�� ݏj���n�*R���j���i�9T2���M�����\b2��#�`#M�O^�A�Iiwl��?K6��+�|ƪ-^q-�u���"d��永s,!�7� ��D�mU�Ŏ$� %%�S�M����J��\���/�)�&v���등��������`�����u)�Em�gb�����ep��;/ߚ���A������}1]�k���w���]�WE]��b��PM��-3�V��8��JCŃxA�d��,}rǚ|e�,t��s��
j��� ��֟��Vm��r�j��3/�ލ�@G4?U�E�^�+�'�(н��q���Q�j�?��oA(�mm�.ً��ز9�*3D $rx��W7���.}/e-��PP/�-�/Q�q��8�R�AD��O���U#������詝6�ߑ{H<<�^�(�̻��#�G-���j�vn���T#��9�
�R�0��3z9U�v��8&"����)�}B��	8h#����ҭ"�,d
�V�Bh�����g�e_���b2������5r��<jC�P
���/b�jmw�F:��*:���6sGg�'�_h�|��+��?�����YO��� 1�{#�eQ�S ��[�e��_!�V�O0�.�祱�-�'����hhܧ!�ǃ��4S���0�n*�#�Ye�(9���ρ�V⏔������*�b� D��Z�S��T�|��	�oir�_�͑f�.ug$,� Ys�2\�vϱg���W����l%T�A��k�S�Y�z�Cڳ�5�4^�-ў�Сf_�ul��oD��P���r�c���S�����@,Ӻ�Z0gMN�{P��W�6�W\�HOF~'S�3���6'Fv�G�i��Y���Z�NC�or��@��~��|�ݸ�����d}��y������-NC���QW��KPݟ��KV?�
�7I�>�<tp!�3�F�X|�e�4��ab~�5�yR9�U��o�0�w�!zҫ����Nε`�z��ޤt3��u����<�v�KWI�0��][�k֊�m@u+�ר�C���=X�.���� ]�\����At|T��~�%��Ӑ`b���Q���LV����F�ʌC/^8�6s6�[<W5����^S��*�y��zj4���K��E�Y%l�$'�ŌA�7�h�Ժ'i7I��D�~}��%�S����t����ڵ^����=�𦌻�b[h{#�|�ē�$�:�c��ȓ+�=w���\�=*^v��ʖ�iqZX��.r^�d��(�$�����4<�SHЎZ^��) 9R-~Y;����?������&�bR1��.R��-_��"�	wrb=�o�@A�F_&PO��sio�EL��./^��y��--ō$߹�n�,Z�`O�L10�@��j�㯫�8�4�JN#����V�
|���T��h,it�c7V}C�+c�=1��G�W�(%��Dz�x[~�����W������].���Q����`1��F.-P|},OI�u�v�ӘB$����}@���ji�`(!�􀩌V�l��nPTߚ{ʌT�a[-<8k�ONɺ�[,���M6#�wi���/�Q5��������(}v��m��㝛a�`���c�c� �|>���%٦����ZY+�}8m�4x��y�8̞�/�'���lX���U}�q�{k����^C��jv6�ʎ��}H��D���a�`KaGD�����G'#�/�b)^z=�PLoa�x�^�9����G_%@��
cg�VQ�+E�bt�x�]0��S>S�.Z�~��3��Q8*ni��4ѡ��(���.� �H�ngT�m��k� �Ux�4��%���w�ާ��icBwX�{H�;!���>������m���9����밸}r�E̞� u�	5WW��m�\�ڿi�^ã�1�C\Q�����콲8��z����0Be�b�B$����N���I�����p:( V���S!��e��0�: ��pǄV��.�N�^>�H���lty��h���}4�'fO���s�J�A^$�����jz���t���� ��$k��s;a���Ae8Z�R�9܅m����*"��\������ _L��F)�Շ�k��k�&�j�Q!{E�ϛ�),����co� ��Fxp��-W�?g�K8��6s�����B�+���M����X���	z�^��Ad����Z�pő�ε�	{-���VNvŒL��&��*b�s9� |��%Z6�<'/��8�����y˦tn��'$�hξ�xn�Ȟ�������Z��As�2xHY( "h�l�����3Ѣ^��냑�v�WVи�[u:}M۴�b�U� ~���;�[��60���8��Igv�c ת�|%���B|,��Q`��χ�c�a�4��cK���FYP<�4���ڞ��@��$�q�/��0&�� �F`���|sY�e��̌WD��$�fq@��Tz�+�!��;�
:[�O�ز�g�*�R��84W�Ě�0��-�E��M�`~�9!p��/0ꮒ�J�A^����٪V�4c�ȕ{7�{��{�S�0���4J��pu�U/_����](�嶔j�a id3:"�(�z��Ciԉ���&�@��!|��z���P�61ǌށۖ�e���m܆����ĥ�������Ä�M\��=�WP��{�&������5a���qP<�,E�M`}�/le����:��ǳ��@�8W#^�#pX�C`�Ͻ\��ZE/�sKu�E�,�T���>mOD�v�:�s?��Ͷr�kDmJGlߚ���5��_ד��ޮ�1�z��8N%�]'�1:�����LP��΄g{� ,���b�%N�IYĲ�űg;����KGHU�:;m��X|��,��O����8�j5l���A�4�\�R�׽� �-���u7�M㑲0�i/�w�	�h$���1)�C�]:���[���0�-��o.�Y�IA]Ʃ�{Bڱ)!"�
rM�B��o�����3�Vh@L�R)���ThѤȽ^���c�������)�wd1�)0GW��?f"�m���{S!I�a�/�k-�ꏏ��j=�r`��+Y�U�3T�ɘ�ţ�90:��Ѯy��0'��`;%.� ^��Wq��x�6����`1�E֮��ݟNA�K?��Ao3E����v� ��������J���:�B-u��!$w��(�E��}z~a�_��;�%��c:'�`�4��R!d2��lS�n����/:)�;�t�tN�>�
{�e����Ϡ8Zj`#[ʪ\���E�A|z�Y%vh�O���ˀUTQ��������jEH6L�v�rj?50��,�>��?��w��d�=i��d!��jk��*��G������M+��H^ m��!�,�|����n�(�(�Ȣ$S#z�-!�܉���y4$P�64$��,~LR�[��T �j���՟���x��,6�lm'�m'��h`�{�}8Duz�:(���p�d�b!��+�+�`��U�06@0���4[V��ep�c��/� �z��Z��M�t�̽5�P�0�rori����n�{�z�#eV��>�W��ي� <���c���T<ٝt7���Gd�o��d'7+��k�1�|�F�O�h���G��l���Og�v�Ӷ�x�t!8j+o�3ʔ6]Ы�~M��I�m��!y4���:X&>�0� �+��k�:,"|d��@d��+�@�\�����|�l�>gJ��p6���0a�LW��8����tJsҵ��Q�B�âLz�JG账��W�TȽ���~1N��;�(~���%ų�W��f�����.���䈟>������(i?�6���zl�;>0���KK�)'���|���~i�湺��ig�_�D���S�H����UE[DXL!<S�>Mx:X��'� O �'P�l��32�E��w�@����O���6�b6���enBq�tx�A�^~Fλ&� ���+�SL��:G�7d�K�췑OCZ�4R_#\r%��֋�i���{�g�������F˒�6�Ӗ�J�w��_��W���{jҩ������GE���<^@��w�:Ϡn� s��~�ćبP�XE���𚂱�O���¾���
���yF���ڶ�ܢ�ڹx/(b�s.� mM��6sf�9���c���y\2�jW}}*?(�#�x�e*�� 4�mh�"�Kl����DƑ�7ݕ��-XAV��}��W�7c�jcx���b=FurK7u�Ԝ���Z+�`��?��$����5���& �^����{,5�>`��������x3���v@Ɣ��*�`yg�� �99�ȍh]��D��?�!K�4��l�_�� P3&m��/�Y|��b�ލLj$gl��w�N��Y[���Δ���s�����݊�����M�A�E��{BK�:fK��^���-ch���,U����y6m���A���A�;Bؚ�AW��	���ݮ4��:���X����t7πe�����vi���c�cdl�GK
<\ŗ5	���|?Oq��.tQke={o�N֬ ���2�\.��]�XW�7�ݠ�<�e��l�*}(�a,˜����76�=�iz�~N�B\C\����TzYjN��7��A�8'�|�c�-]���	�������8!I����;��)�E��=�%W(Q����y�ܹT�Er�2ސ�_v�����-\q��nM9��#V��l-gS��;���T�o�z�j 2�F�ҟ�|ܢF���4�5�'��k��l���T;	��f��M���XnWC<�ma!�7KN�[��d �
��{�)�#.�"�M�K����>bZUL"��3 ��ɃB$CudN���&�U�%���\Z����H��ڸ�����ã���"[�ʈ��=�&�ֺ�e�p��l��
A�N��$/hq�~�w�?�{A;�4�Ǆԝ�7�O�,��Z9�.� �����*!"��@sb�!�]���-�?�� IA0�d[�/#o�IC&�i�V�!j�Zc�؅jZ\�R�B�����������l�+]�{��0h^2�x[��%��Ȣ*c���O* T;-���,�����<�m�{��?��#������\߻	����u��]�<�Eg���rtl�fD���q+~�M�G��ͮ
'����q��������@��~����W��1�z�+r�eBT�fx���
�I�ԯ��?\8�m�����R�L+p8�b4x��~$L�o�qڒ�+���Y��O��3^\n�Mtn�{>��7��2B�����ʄ�H���D[�E���O��Hv{\��@ۍ����xJ9W�G�^}4��F��d�4����M�5�QC�ߋ_-��"�x9w��YG�L��U&C�5�=XH?/�ej?�������Q��U�Gj��&�� �{�T}�Ab�[	��o2q'R_	�˛����@�[3��3�,j����k���n@=7Ȣ��
�(}0�?���Jl��E�"ve��eE�;��q�͉tJ^[z���,��<�*C^x�d.��:��Ed�%;��b�J�^s���8�ZR@8PN=�8�\�'�pH�i� �k�k�^�^�`�1�GF�h�j�{;�p�(�q��/�--[�9D@������LL��Q<�hR-o#z�L�)>ق�+�F�UG�!��[�p���~#o%� J< q���]/� V}	U�U��L�9�<�o��Q������C�D��{�.���j�gwG[�:��lOo66��,l�G�(�T80�>�q-�No�����J�v��$0�m�!.֭mQ;r��W�7��ax���O�ff)��\�^��s����a5c8t^��`���qDf��~�t��e�K��:{�z �n��U�h0�C]G'
T��#�E��
����%j�ySSȘ�ޟ�Bh��'�<v�ͫ�XW�`aV��!�������:ףr�͐h��i�a��y�QVr����Xdy�TQ�}�=<#(�Zr�i��O�ҿ�:�%0�y:����*{��QҸ��L��CH��J���́�*W_�������΁^���jj"��x>�nT��� JӝPd,
Q��
��w�H�į�6��~ 7��t���"��8����|{�/B��={guF~�߾ ٚk`,/�*��	m:�w*��[PSp���	�w+�� X@,��q��aD����!����s�VII������cJ-N[>x[QF���N�����nj��"�w�d)�Px!��>,x�E�K:d����|Y��������9E�g��+ ��60����Z蘹�s#���LJ�ؔ�*��m!Q�?�(ۿ�e��Ư�#�lf�ܹ}X�+����Ȱ]�G���/̱׉}�y%~��
Ri{73��;��t�:�_OEI:�g�`�p�ϔL���s�b?�YF�ZB�X,-|ādTڕY�q�� �3�"���L����Bp�/���]E�S��G��Տi�[���t2,.�e^14L����4`t� ����d���%���,�j�uD�t}�H#NeQ��l��PRl Ȳ!L= ?խ,|t����4G��-Ȑpdݠ�bͽ��=�$����Z���KdX���%U9m���ч�& �bI����>H�PMuj"� P��y�vk��̝�!���M�n���S�ޔ�!��K*�$^�퟾�2g�_�xbS��\tBH,r@H~AB������O�=�ʦm�}��K�����l�O�)3�UiU8�`j�e,���Ds��1ۍ���N;x2��c\閌��,`v-�97PW���Slb�[�@��X��X��8�d�6�']%��.���$a.�60�B���F����}<��͋v�o�t1�V��Ү�Y�1 �h���I�7~����+{�?�3� qT�s FL7(�O.ɏ}�sF�q��e٤j� M�#���>f/fr���\
�[�k��11�wS���RI�5�VF�<^��[Fn�Lj;���iß���T�u椰Q�1���iD�`ǟ�򉴽o��$fN����Kב�oQl��p� �/�:"<�\C����~�+��X��վč��~%p�4���̳�E\U`|D�m����XG#�)���\�y�U�����~����4s3&�Y��]3`�c\+�h'f��>�f�r&�I�������6	R�P%*����Eջ���g-�'�~�m�4��S�J<�q� eb�C��ba}���s���ػr= ;��|qݿrl+K0[�LO�z�S��C�ӟ�|kb�@)��n��h��wR0���l�=��U������l�l˟��J�ͤ���wx46�����H�ϲA����-�3a�1xn��H��|J�!�"RPo��/�,'Y���|�ckh�C6�G����ǟ}�L��'f��������@�)��M���=k�z��V��Ѻ���� yZi��P�R	'ư��th�ŨW�T2��״|N��L۩�sWQt��)>\@Е;�0����/�:e�$�F��'҂��� ؘK�J�f^�H�ble��#���'��c��a$_�[�������$%�'�|"����hh9��lj6��+[�U)PQ��_�.U֡�1�k� .2E�����@.���
��	;i�E���4"��&L/��(EE����1�z"�y�[�h-�����2�\�&��bZ6+�,�WX���5�\�ƚ��'��/��I�){!��b�i<�T _$]ѕ�j��J�Ɠ�[t�ʱ)<�Nf����q�7I�*:j�s&�Q�R}T���(s��ʵ�~��*���Ek�:`�d�	��|h2k����&�a>��g��*VKPs�Y�u��mP��*���ݯ�
�0[�[�4v�z���J:I�縡,͐t'^�UP7����X��^�����HΕ"��od]U0n2S�ץ��|I�ɉ�f�I���ÚC'����_49F��Ao���v�fҧ�L�O�E�B�O��_�6�q�.��M|@�Z	�=N��'�}�TB1��[� ƫ��P>5��z�YqW��TX�����u����L�r�a!�CVT�|���#�.�2���1�5��0���DY�����V�u��QOql�V=��j]��v(�O��`)k*��2�/�K�mu�]W��D�_�.PU�v|%ʖ����D`#*~b薆�'C?{3	ڊ@�@Q_l�/�~O�r�7�,+���VRـq}_�����/��03?��R3�g%�kwѹy��N�q�,��}â�T���j)<�3�$�L"���ʒ�t��^�ח����\��B�Y��q<VG�:{A�����O<[@�+;ؒ��?��:��q��O�<�q�aKc�##�&�ݞ >+�n�i���*�����0�urr�z�D�M����o��:!��xvx��u�`)Qu�,y"khn���iK4���F#m��#,2�D���[<�q�v)���t$C[]��\]��[3Il�rM�f/�ZuQba0�
^��c��f�W�w�z���=X�+��θA���'+��.�|}ʜ��GќS���Wb�(A�8�\Wm{�lf��.P�Hbb�/��1Cj��^�/�2���1�����'��mM`#��U���y_�RkV}�	u�I���v>�+ 1E�*�EPL���拱����!/%��H	Ops���˾"3,�J�s�\���-�p��N=���bY��09�FDk8�!Y�d=����j�I����ۑ�����S(;>�*g���$v�:L�(;ELl�κ��Y�ۣP�r��ei��B�$m�V5��+tL~^e
MQJ��R�s����٘F0�>
"J���]@��������rD��L�[K%
�B[ �Tu����E_�	�J �a}��u�!%p��n��O��0f�����G��t����@�h�}�W#��S��ô�K\��t瑕��x���т	;h q[
]��{;c������E4�P��l&>�
�ă��.��H���0���p� �D���1t����.��8��ϗ^������K%�8�ere��ű+GV���7��]�{o�s�+$}��QgB�N�m& �R�L�rڢ�sm� ����ӫ�8�(|��-k��[����1�>�'���9`�jaÚ�kߦ���a�r�Ȗ!��j�Қ����5|�NX���L� [��^���b�����KJ��+?��IS���Q1{ߔp˴��|� U;�#�\�����Ë������?�Kn�U��IBi�SJ����e���>�C������>"�:��R�@���#vIzs VЁB/�q6�p�3��דq~���N��&���Zj��Q��y���l�)�����p��7��f����]	X<�!��֏\�J;|�l��l;~e4{fd��O���q�a�7R2��F�*;��Y���sS��hvx�Z�3Ea[sJ������3ڬ �>�n�ʫ $j&��DV�S�$��[�ba�*��tl+��s�-�1�?CI�"�I:*��"���z���J���e�a��7G�0x�Z],+,r�%�7�ȿh��Z�
Q/?H��`�s;˥���3���@���-]'N"޶й��j�'��P���s�7C�m���N��W���=19K/�P���� BHA��`�O4_�":qtԯ2�|E`����/&8$,UC��0� 9�&B\H��ܹ�@��Y��=����5g9��� �l:�'�����x����d@�<|`QH�WJ�k�X3@+a]�����B���t�5j�4�K�E���S�_�?�4�iw�K���J,m��;�Z���1����[�KW@�"�!�<1���ZRȻW����t<�A��,�?�U>%�
�̪;b�f�ir?
�3kN�d�����5x;T����(���,"nf�jD�
�@(�خ�n�c%捌 ��O[�f�v��a[�|Pq��Mi7�e�揩q�%j����@$%sGW�	�3v�)��YY����9Jx��J:�kl~l����z�䯔@�<�o�r\X��}�P��R��T�6@e@/�T�ۀ�-!ё�'7�>��'�h�l�ܟ��}�P�s��ܬ=��^��; �?0c>��0�q	��Z0����	v3��QD��@X�q�@iT�I���xD��U���?A�K������1}j���	á�O��yT����I��Y}��?J����������El��� ������4���b>Ew���!+�T� �X	o��s�I�$*�;`g��af�Q�Ò%�|t��Qciu6�T�,���Q0s�2[k����?����r�gc�?%%�ǘ4�D.(c(�Ǉ�����<T�i��A��&��-Z?Ja�d�f�M$��k$���4(�c/Á~��6-��:.N�H�P�����1~����bFUx�?7�iJc�<���_8��(��7���^>�	t�]�O?�|r�(��H.B�����ߧX�,�HtTi��Z��>`��=����*R�xg:��W�@���;ƥB%4)Ǧt城�qH�h�}p���sh�}ѝZZ��� ���ug�y�@����y��`b�q��[m�	���R5_���H8�C�C ��	�2:C͋J����Z"�R��{�wXNK����c�Ƣ�Co�!7ⴻ���"�PB���{�?����17ÐO�EOaM֑�-V��������_X��n�E�}����6 �PXV�4
�|�\-��­Kǫ�����*=0sq�&&�,�@����DZIַ�Oy#���ېI�kY��l�ā��<0ہ	�z۱�y��`��3���?�VTN)��c���S�T,�?�Ý�ǣ�����y	;͖n����ʫ���Gj��G�zSq���Cx��~*�����AY��R���$��~�����N�M=�5��[�A��ı(�ov�q7"��Ƌ�QTC^]�)_��%��
:���^2J�~o�B��S4_�+ܴ���&]�%�u]�7��	���v�,8ʢ��Ǘ<���v�y��V���.�����h��_F��ך�i9
C�]_��Tv���.��= �:��$vK@-��J�Ȗ�@Ȃ
��In=3�k�{̑���
�?8ҡ�Zˏ��!ٮ�F��ݜԪ�)�lb
z��ϟ���>���EH����-p'�@pQ�J�$�R���U�ැ�$W���0�"��i^��݈��O+�j�|5>MWW�Y�Z��K��ʝkF�pւ����d�k��ӳ�T�����b>q�V�X)V������w�C{��>��S��G��1�G/4V��* 6	�g��Y���3�<G��$==8�.�'�����gh��^2��4vJ��n�QV�8ǯnq�^��4�ET?Dc��S��sw��z�����f��>i�H1WL�(�4x�H;��j=��v�ۂ&j'����	���7�v�������vl��փ�v[O=�yl��u�ʕ��Y�N�G��L���]�>b�e"��t*��k���&EȆ������v��<�r��-��c�
��������	l��%[�!�㛅iC�_ۜ�1�[�?��U���2��-��V ���:/hJ:�ԫFJ���L�߿�T�g����s�>����
 $��ח������!�B��C�f�~�j�(cӮX��,�@=RF��C�_�4�	{� �fF�P���i:�ݤ+(�S	��s���0��z��$�v����O�t�f�7b�NiǱ7mӈ$kk-ʍ݀���D�L�B���;uS�9������z/�a^d�T���!?<��5M�1�&��6��'���y�ki�x�5�=*G��Y߻5�푛�}V��0�r>}��ŗ���Z00JH��֜�Yn�/R���x�aM�a�qc�bn����{�3���� *�9V"ּIߟ*] ў�3�N�(Z���<ꀪ�.Z�
ݚ���E��T 6���:<�I�x�� O�)�,��=�+�Щ�b
��
�mA�eUK1V���E�*��1�Mo���xJ���M�_�~����:�M�7
Q�Mm&���b�k��~���M�Η�}�z��1��G4Ȩ��[�R%@��JB`"��T�&�Rx��2����c�@� ~�j�+�w��.��[r� +���.L�sV���=f�"p\�S]S��لW�5i�����l�}s�~�D�"��-題nhH��Pv��Ш��͇�X�HZ���t�ȼ�������'�)�!�V����붹P�<��:X&@0�l�w�0z�[��32����Vf�����6�kGH���?����Ų���\E�k}�J:b)��Fu�Ҥ?�@�d�s� R�$�]�oB�H�eK�q�-?������n�by,���aQ��
@�QsΩ��O��z��P;ɂ�lb&��Z��h�Q�1�tH�^ŉөPo����Ao�I��otX�mZ���nw;� t�1ɪ��m�a����!6杼�EI�^m|s����w���\)S~�Z�=�oZxŰ1�)��{A_^T�T7�@F�K���I�����hac��
b\��nA��>m�uXS��ͮ����	)x@�Μ]�����\���3ԝa�B��C먦
��f&(�pqWp��R<�;�r?XS���I�w`�_B��:�	���`?[��K,�y��k�?D�\��=P��'f��ْk�%g��(��( 
\���%Q��{�g����Y?&��ic���+�T�dGv�Ľ�GyĔx�E�1���8�Liʀ2�R��~T�X:�������JD�>^�M�q/����>?Md���X;�H8�񫩶�}��e(�U�Щ��c���k�g�������2T"��	>��د�W挓�X?i�
�K斲P���m��K�FmΙt��H �]�3�j�)A���po��KK�3k����R`�?��������Tݠ)�>�ڻS�^��YP�
&��8��_5�D�=~JGeH��檱A�4��N�Y��3gv�&`�k�� 1p��aA���D��Rh-�D��l:쌳s�˽Ϟ� ����S� �����o0�o��������Of1;�^���_WO��(�B>���	!6A��x��t����� W_n�Ϋ��\@'|p$� �-�������jkh_h:#�����lg��!"Q�;E{9
JÙ�p�A�������"�+J���.���0��!��C{tR����(��P�aΣ���֌Ǡ�d4I�#c�&	����nA�A��v�Ж�׍�H�B�����\+	���U�!N�%2��=6ﻇ��QrϾ'�hz���%bHl���W�`�D���h�V�
�@��	͆���'hm����K��&��	��j����(��'�-樔�hA�D;�E-�J���t�l;B�
�<IL�;E���4hs�W+����(�s��0����M�q����>3].C10V:�P7v��g��Վ��'�1L�T�Х"T�h�]M�i|Gsa�_�Il�tp>N4�y�x��#d��e���p��	h�ؓ����8�7��L�`ش�e3v�@�t����8��z�������?��bZ�����9���Q����7��n��c$r-�:{(����P-"�y����lG,dԲ�{�*+��79����b}m�f�څ�ʡ��sͦ�`��Cw;���s�rH�[����m]�(�����2�ӢtC(<��5���<d����'�u�=7�f�z�P��,��/���}(�.ݩ��.g�5��z	��K�k�,-�L��dȼ{s~���p(k�拱QsR/��ë��of#�0���~�v�'a���
fHHb�=fzL>NN-���'�Kr�"��觠Ύt�P��6ej������A�3����y�pc�j���&�b�1��d���4�w+@9_��"���D�)�R���Ms�C�8�	��_G�T����ֶR�2��_ӗw��j�D��ܝ�z4���DR��g�`x�4������Hy�,Z*eCԂ�y�v�Ԥ�[ e�~o-�9�5q��?}zwjU�@���E؞�H-��b��ޅ�e�<���;��m�x���i.i֮�~��
I��~����a�ߊh+s\I�[]F���w��D�d�a�t1�������N�*�������%DŃ�?�;��\^�*�[�����Eĉ�)�Y�m9�aΒ�R����IJD���3��J�N�����mN�@�7��D?�S����6�܅�I-�l���4��]�>N[�ql�v^��������U��"�5���:-�`�g��]}�-�Th�B|�p	�����"Cs:q�+YfbP�7\�X��(Ӏb8��^�XR^5E%�j!��M���'�$�=�̓�H���Z͏n7�f�]��2eP��EV�_�MI[T�-2#*���v��#8�`7��ē�P�ni�~��T��\�8]��߅���f� ����3�}�\z 	|��+�7j=,a��[0>󡬣~[4JV��.4���Js����L�"s����ʿ)#[iQ��㬱�㇬�#fʐ\��6>\1�h�l�M�̃�	p�����J�2J~
�8�z4-�;�Rn��!R�{�Y�e3�P��7�nj���E�|b��p�ޥz��M"�̬�I��έ%��頼e��奰S��*���ڸ1	"'�/��=��������#C^}��E-֊!^����~DX�	�(�x��"9e��`s[TS�B$q���,�ļִ?�C�ʱ�w���B���;�9�Y<��|y���fUwA���Z�tC�^��+/�Cѳ��m�M/[�
:K;h�+@w���u�<0T?�~��p�s����`�n~��\�I�"]��Sp���O���?گ���p����r�o�az�ߎ����+�lq� �B����?A����Q>ZY2���_�^��������/�S�Yh�̮z�y�LQe��A2�d�������*n���L�G�{(�}U��Q�S�N��K65�e,�b;uy�(��%�p��;c���xjJJ'�b���j� W��~u��ǩ�px9�搻\�p�R/ě�j���-#�����:��o�`�0f���e��g'Ɨ;Т�,��r�]�&4t�t��<��Q�����|��R]ތ�����q-oK��6m��w�h�>�&�����5���0I�Ҟp ���m���}�U��� �_W��ʙ�2��&$��H{�j�FJ�Z�`>��XKA�U�k�Z �?����k�OgМ��&M�N �4�>u@�&�
N��lUÏ^�P�E���!p ��mԘV�3T�S�:8 ��_�/��ʙ�]�ⷜR��������(�����B@���I:����z����挃�̇��O��WjY��g�	�},C^?�+�U�aPD��A��|�Ğ0.vlG��z�ZX�D4*v�)�p��*W�|2-/�t�az	.����6;I�l4�b{�!;��CF�!�O����H	&p�R)I��?�3?�CY�Z("yn�E��˻!��w峿~x�}�钘I'}�BXP�JdmEZ���wj�W.�t��P�l$<%
�~.���,���mh����0I�n�4Aj���6�I>�*&nM?#�>�
2��Z��U��ֵ�����S�d���n���7��&���[�P�|*H.�����4��k�犃��Ͻ�X�0m�T7��ǥu{�㦆5;z�+�$�V�p��"Γԟ�x��M�S���tq���f�f�z��QRUg2���f�Jp"B�iې�a�I�l����z�QY�$T��Jc�43G�e�(8��Shz��VHKް��@�QC?�'�>9�,�1��E�eB�a��O�����MVX��\dT,�&^쫊��>��=��)ћ��BXR��<�C���R�oAn����4����3�2��uԋ03��
EdM$f�s�U�2+�o�� ���NNꨴ.�&�G�|t����@�۳��H�r���F��@j�`څFU�Q4�� ��;�3�Il��l`I�{�#���$�[m�x�d�G�'�p��2��X����뽜R0fg�t>�^n���0�G&} 3�Ee���XMa�i�xV�tG���z��k��$'hH�d�#�(;��P�7Ȭ	���*Xs�9A�m��D���3���R����Z�X�[��lc���}��W�b8�ɞ;��ڳ�.F���`���;�F�w�Z���Y;�_��ӿ�`��a.�EfTt��$����&e.�o{D��0t�@�^A��+�D_%��ż^N��eH7�M܆�Yk��-����(Lp���G�K)k�|A����NEZ�6 /ޤ�eF��ۊ3�t��b�NG�����*�;��svj��UDBE�	�tm�5f��iHY�#[���'�c�cU3~Chb>�lí��p@ZWU�c�+�fg�Y�c�!7GAX؁U1�*���<��C<�S�S��q����W��*w�VfH�I�����$���'�\GHs�����(�i,�U���bb��Ш���bd�,�Dь��&IY�����\b9�3���a3-�leR�7�q/�l�w����k*�'h	�, �B	�;��v��ӌ��^��n�X@�/���u TI��f�u���3�!�ؘף}@���$�|��b�E��� �dK�ArO+�f��\��I�,��2k�,��.��*L)b�+��5�[�#|�L2x����b�l�]葁�,�bm���^�����΍�r��cV�ֹ?W�6�>�p�pD���?
���CCI��E�5]�#Q��:��Tdc�c�*���o�s x��c�g\f�-u�<� �2������Y�m<7>�)�'���[F��$s�@���sV���7��X?� Iz:ae�B63�0�
�qE�mx��&�%Ch��QU�R��Mn��Ԃ2e���VHkF_����Y�+�V�mC:�B�Z٠��[g��߶7tW�Z��:0�q�����=M�jqN��G��A��9Ξu��+f\~R����}d�)�����9���y��T��Ke�ՌMR�o4�p���.q��O-����u��\%�(��R�������>�2j"Rɹ���9A1�M�q�Wp�ڵ65I��d�`����6c�brN�;���>���	6��X���G�_TҖ��Fl�1��u�C���� �� ӳ��	�@��e7���B@�m�&��hd�V�L��2�2+Xc�{Ĩ��' ��$�B��N��4"d�>"��,��f,^c!���tK�.vF�x�h��dg��s�{k��ku���;x�e	,v�!x��U�D���T�2+ON��v����%<�����Xo�G��.A�%Ji�c�Їߖ��i>D�W~�Y4�<(��!#6|�����@[�
j",C2�Qҝ�'�/�W'��~X����2���EU_�2�~�<,j���u���H���nt�	�����畚�)$�f�ä0�&&٘s��}h�} �,U�g\�����Z��هB��
ruc��P���g)�{�قb�(Q$Ay
�aE��
2��jC16ރ��Ȫ�nww���b�,`�S��Jo�f�jd��5�U���W>�|�P���I���@��I�n��K΁�)�Y��7"V�%9��e��}�2�7�l��0��e����3���f0ǜp3�'Օ@��n��\{��A�5j~r�/V|^�/�ﳊ�8���	f6����^5����=Ȱ�2e�c��V�q��N#��K��F��w�:'�Y�_���T����Z�5�0�+b���B�=�w;=y�&*^��?2�0� �/�h�?ܭ��7���_g������x�C������J��-��H��u�-�f�=F9X�(Ѵ��
�OQ������pj ��tC����k�S秚A4#�����Ti��_�+U����e��븙^�Ty�`U�8]хm��h��\�x�|��[�ۢ�؋u�)���tH�@,�ǉ���������k�K!��X�;�)��%sD�s?�5�Ml3��-|�^�0�klի����d�ͽ�.[��1���+�5�܃�z:�
$�fO��!Z��,�� ��O&�i@�L�T��SX�'.?MD��]]3�H'�а+.�&@k8�U�	M�:�?��Qy�]'��<���y�񒠦;E��P��d���0�{�`ڑ01E�N,d����y���-f��~�F�*e�� �H�T��?�w�	S�8WZ�w`�t�����0u�=����2����b�M��Ͻ���S0Kr�%M��q���M"9�m!<�w�g����7�="���v��3t���e�̉Hd�y�`�QǄ�w!Tl�,[��+�g�,6HHC�<�j-u7���I'�Aκ� Da:�B{���'(�4�g���+�zq~uS��np豬�g([~�u@��ȗ�/�@6Í+�*˥�K�R�˨�{�MkWt��ͳg-�OY
����«Ț����P�q:��(B�ֺ������"5k}&Ȑܛ��o򙒽y����K��e�#�H��*�4k�tp���M���+�~˱zyg�^AS�������vT�E�2�{���d҂�u&(��ZQK���A��\L0y��Why*����u����_��pU!a��	 ����`.�ׁ���?zUm��et�����D�[L���z�U��8��" �;b�u��OA�Prj���n��$3WP������.XL�<�I���n�������2Ľ�O>�>�X	��@l9���L��x�{*y#8���0�"`6���6c�Bi2��{ ��E��1Og��K?�C�T8����n�Fo����h?r�!�q���F&')k�͕1���azQ�6�ЎAY���5ƛ�f��]�L7t�=�4ͽ{)�Glm�λ�����g�О��.��:�>>�W��$ۗ���G��ti�_�'xs,o�s}u���jG��j����!K�� �L�t".�ԭe�����IM�g|r�>a ����<�Y�B������4܊�������0.`.�ʋ]AS��6P	���e��jz�F��G��-Dy����.�O�@3D��ڞ�t�y�P�7��n���>��_L�����ǀ�d{��zI��FI�j�7Z�P�;:ե�����`�xaA�$��$  v�$��h?.��R>���r ��ze��R�ǂ�Bֵ^]d{O�$���I#F8|�A$L�� �^=�uƇ���[���~���~Ϛ%�=]&��v�ۀ���1c�;M����l	�鷬����@.�-����zb�zd���14�֍C� {NZ�i!#�U@[��D����Ou��,�����L$�/��a�k�+D��[��M��TF�[Oy�<*��U�	5��������Ӊ�2�(t��������%��q���D�:D��nG�i��s7�y�Q�☇#G�_�z���߭#ri���=�eF��3�m�BarImt3���<0<���Q�{~E/�S�1�K=.t���#��ir��A �l�ȴ�x3w c�9L~R >H�uZ$�sk�B^�2B� ʹ&�N%�a�������]�k{�
үY�Vq;l�E+�$��^�G�O��ݭ����0Q����-ٿ��K�� �Il*���rT��ג�t��M��	��^�'Mk�!�Uǟ�l�1��~�kd�1�xW�vغ!նb�p#Hޔ2�o���CVeT��/�NV�h�^@�]��&?�ET�4���� ��-B��sF96M�]�s�b&�T䵜�k�!�uߨ�A��gg�
G9nf>g"���Ю�4z�qh't��&Q�Ԧ��v˙T�?\=$�{ EM����T.��!�#�DNI'6b�E�>��yi/��Pu�B$Sc�4���xnYɪ�D�J��|B*J|�C���{��F���j�EX	�,��=0�Ä��'���{0�O'Ho����Th>��4�N/G�Z�ϩ�j#n�")��PJ<�k�}�]'w�#v:m��f�K/Qڄe����(�7��&=�jn��ģh���i'-n�����4m�hu��ç8�GtML�Z��WT��P��M��j��X�t��JOEŔt<]�:������_��N�9�M��=5���q���i�bN	n����%�,����Î�Dؒ"��O��SX���q\�19�&%Oy��$�u�Ws�~�E���-�v�sW���\��i�@��yP���K;LtX*����R~�3L�O�0��✜u(��A���B�FsUo#��΀�����?��"cj��%�L�y�dG��Ծ��������[@����,���c|Ó��&��i��A��r��.ǣ��/pξ�ƮQIC2����m$�Zd䐯栵_e�K����KZ<E�7砷66��B[1�5zϺw7��NB��Fr[���"ZH�л����I�����ag�Eu{i��;�6i�s�z둩%W�Ĝ�	sx��=/���!~kIC��B���t�D
���5m���‸�;���¤�oOׯ>��e)#s�9�2����iwdao<UG=
aP7�	o����YB�
t��9��ma�-#Ie��f۱���Q���������o��,U<:]���*���Hv.ȁ9:�wٚ��9�+W��*l�NiYN@)"�i�P@��f�����|��jJ0B�q�n@��I��n2��*=�x�IR!�c���Q,���t����
�����3�Yw��D������HaIA�KR�N��5�Vg�*o6�c��C< ��G���~�4`�\� ]��MM=��Y��%B�O��)ع�x��l�`�"�#l�a�& 6�5���fo���J�����V͠}M�5p��K�O1��a/�����l�!4���#�WZԇ�<��0�?��p�+S��7C찟d�8<����;5'Rg��j���R,���1OO�닆\*C]�,�����	�S�Wr]3���X"���'4�����7���+�mv�cq���7�Eڀ�@[L2JgH:�1�+�̸���ɍ���G�Z������\n_�Ϗ�7WJ�����+N�=iǃ�$(1��Vo�h)�5x�`tRɒ>�l�_��:����!#�W"P��ea*2Xj5�T}�JA��aͶ �Uݐ�Z���w�i'��	р�Wo��x=
s#k�@��ly�D�>��s`6L��!�t�r���Ðށ-;*�a8SՋ�!�
�=�^�ͭtd���M+��'�����Z�k�4�
�oW���	8�E���ǒ���l�t�+��"��H���\׸���gBQ��a�	/�r��b��
��6����._S� Ō��):���\&~y�	���#g�,8mmk�)%6�[�-b�K4�?�����K$����h�.ɠ���;�Uz�9O8%�;��y�>��vzZ�}b\ܧ�Ub��D�S��jH��x�Si����]s6��.�������'}JP�����gLɠ��RB@��i7Л�4�AbMZ�p�eYFi��O�Wzm��I�����!�&�
m@�dիk�A�S�����H<���C����S��,IZz��B�_�"R�5������|���ȡS���1(���yfD���-��}�=+��г��дv�O��r��K����h��D�t���{��[��
����(�i,�IS(����G	�z����F=x�rn~u6\�s�
a<�`�.i�?yJ�X"�AAJr��������m<��������h�=���R`��F��Vٟb���:#{W�C�S�Ò���;��u)�@7ЍÇ����ᕏ��s
d�5���JcmRY|&���VG�|MY���K����Yؼv5�.�x��.L�B�J��V��	�n��Sj���,W�Yy|����\�D��^^��M�чN,b�����}`�qk�S��A������f7�k�0�1�d7vȥ:��U,�vXeЁvtA�DbI�1���x��P��~�4�) /~Q�|g�tWz��vg���a��YH�h�����%t:�˂����3���i��
r���j��GY��� ��n���`��bQ��⦳��# /Ͱg ��_�#FXO,-�6&�㘠��0%�Co�������U��M?Q�u�>�|4��B��ņ,!����e�ʪ(���j��_�q����x O���ۊ�=�V�8��$�������Y,"�&`S����7|h(�#��ޘ�i雘+��"(�������֚�bz�Y?���:�sd�d|I}�c#Z|7�@��b.���W��Ŀm0Z�;9h|��K��vx�jݳH����Piq1�E$����QAK�m{��N���{��b;���"q}�f.L�͉D�pU�P(Z�ϭ�J��Q�oB
��PS��S��%1[0[��EP���^�>��$KR��Y� ��o��i�����L�u����G.��>P��Y��7�u8�ً�u쐨�ӓ��
��q�{��~��O5(Z'M�q��6�N��S�e��x����ܰۢ���[�u�H��s_W���wa=i��R�#���ĉbK,�tbI_-D�
D\�޻��j��To G@6z��3]~��eC�RP
����JpoG/���F���r�ߵ��������ͽV�\��Ue ?��{|z��9�����V��_�w�UlE��dN*�<��N��
��/���k��S_�r�����P{{A �S��pH�܊ZU�D!���Q�3ي��+	iN�96�A&�h"bm�����QM�\��D���  >4������Z��|��F��C1�ou�׭I���i"� ���))0���<�TYi2A�#~ԍ]#�O���ő�x	�%#��Z�D{�� �A�����\5A"�v���1d�Kz9$�)=>��TK���Os�� �p�%����*��_����$�4�$�}�N�}r�/���th��1z\�4�	p7z#�F�\H�;Vި$�U֥�شЇ���T�����Vc�c�'��~ʃ��[ϋ���S.3E��S9�Wc�߂�����`��e��%�QT�E����Sg��x��
��MV����D��~�����5�qf*G�T��~�@�效�G^owMT���|dm�
�� =Ez�ܶx(���-+��7�f5
cWPc���?9��v��N���?tH��|�t�ey���>��������OК8a��b�д�����o�`�`@Q� 8X%}Ck'ͳ��蟌Tq����"��X5{��]<Z�85\�a\&u*���-��Ö� �d`��mqp��;�mD �&��3��������@��A�Pl�ȳ^�E���Ζ"���q/kH���{�£ˣ8�Á�(E��G�0�c�ekU�ke>�<�Y��*��>�A��Y�7$֠k�4�~��Q�#V��2�qW���{,���1#>��.��h�����g�2H�݋z̹Օ�a�?K�&�U���w`������Rr������͋E�q%O��W���b_��̕���'� ���ܑuΘ����ŏM�j訥Ё�׻��{�Q�cm��`���*+�B1�˨Wlأ�~Gr��z
�$/b�)O�d��n�yű��fXcc�= 	������o6��.)�@"a���'��$p�X!"R��"���]x����I���t�Up�l�-o�j���u�HkyA7��$UI6
�H��T����k�Ӝ���K��%}�fU�\Xˋ��R�Ce�^�k�ӆ�({��(aXEʦ��-�F���U��$(Wq���A-�z?����(\1�UG�Y��8��[wK{�wӆ�y�&C��#����2co�^<5Z��7C�F�3�n��	��B�{�d�g���Fu^2;�_���	 
����:�(%aŊ�R�y��q^Kw��}Gf��R���b�}Y[4����m��"���~��yϧ��i��K�j_%8;���^6�j���aK����q��ZgQP�s�>;#2�^��`L��φ�DSE��XC�6�	������]ׅG�w���9��e���l޴v�pEr�,qK�N�Ѹ��wR���b 5��gcel�ӱ0e���.�)���v���h6!�5�e��U��谄R�����\��5`���7�,C�O
fgU��u\��~Xh�p�
ۦ~
%=ީs^z��a�b"طM[�X؟�����A=�Y��'�y.,�P�o��͝�@L�3
�,���:�|����g�:i�j�#��W�(�\n�gM돔(Gw�΄�)J4dl�;f����w�&���:�6�2��M=����I����* #sw���(����젒6t��ʤ���=@��f���>^:��!��ۭ�<��h�*�������lB�n���T]���+� f+@�Y_��1�<AZ�J#�h�*;|[c���J1��������*���2�xwsd�Ⱥӹ̘>#s����ꉏ��e�2v�N9L}wa��aw�OiFl?G�X�5f�͈��-[,�MAL��$k3�(��+�H
~�l�PzF�,=����*̻9�%6���¿��?q�
 y�ڔ�-�6_%6��P*��j���%��s%��R�5h\b��Q�)js��s�W�ā�G#Ni�:gt+��N6M �)�ЄY6���2���oj��� �a�O)��#��o���/�4isz�8�=�j�t�OcE������ �H|�,/�Z�?�8�d~���#��I���@"M�j�� �=axb�9:I�}�.
��'��t�j��j�b��Y\O��|�ulzIr�g��ֻl�nD]#K���q)H˃�Ll�"��h��T�W�.B���< 趖���]��z9WV����a��:	��7LN�B'��Z���\%G����u�H�#�nB�w�D�}Ϝ�̐5�-�}�L������I^]9|fb�i9l<--Y}D@�׼�n> M���9.ي")���'6j�qvg��ؘŞ�I�3��d~�X��ҭ��(� l���ʍ7Ҡ�++2��@���j:j��Dz�O�g�SD9��=�#����/��$aO+����\����r������jQp�s�p�S�TgTl#��U��n�>$�^�Ŭ���K)�c��:2�h�Z��^�N!�i{���P!ƍ>~t:A�|�G�;TJ��;�ӱ��h�B_p&�Μ9p���PѼ[aͼS#���F���Y)}d]
���?��F���P@O#{3i��F���8=C��T6�`��ͱ�)�	�R&���vt��xÞi� 4���U�͍��p�?���w��� 
V���F�B�����55�	q�;1-r�U���`���r�v�0C�10�]s�P��V���>�Cۜ�5+(����+1�Bv��iZ\� _�Ѝ�:u�U�Lq������3Ru�QT?wO�'t�<p��
��!�[����HC+%��Ij���A2�4��V�5D�R��5i����ks����Rp�H�@�/<)�g�������~��� Ȥ��.��+יJ2[�麎hE/h�w2���;̰%��4�`Ձ8��(��V�1�����v����\(p�q��')�i��������ї�5i ��k�����K���� +�S�iثb��%,uR��E��^�kWz��p��'``7V�gx6ŚNlu;M���xq'�̃D�L�M�ޢ�љ�`D~[G��B���
�����M�+j�;n�����0�L�%^����$'Ԉ����C��l�_cZ>��W8ɟF
�GH�������M�;1O���u���?��ᓗQǿ���@G}(LeJۏ`��<jI`9:)�ۜ�}�!��3��NP�E[~��T�|��� �}�V���,�B�� z�H��Fjd^�*���m7�g���򾙴Q�(�~�ۮ���]y�)*^/D
H�c�]c���P5��=y�}X�&�J.�j�u���TҬ`>�9��e�kE͓����+�dE9^|>�G�jP���QK���.ڈ]��1~��*p���;�E�a:��L}��mϪ���)z~�ɗy/������Ѐdj��|M0e[���[�PW�?e����~�1rG����mi��wf��0wI�p�$ETњ���X���6�t^U��� �P$C/�o��m;��ָ�(�7�����a�A��C���/B�DzVw���#1fnwq>.կ��<<�P�:ְH������=q���p�g��!�>�r�洍 ���BF�!�!��/�5������Y������3r"�B�C.���O��{pj��Lc�t��3iz��b�h&�䓙JX�ɜ��[������'IM߷��Mǚq����bg;���e�n��e
�X �&��2�7�e&7�l�*�mS+(���9�m8f��T�t�(G�eR�w��#J��x�2(��������N:���# V���؇<����ot���Q䅏�ҙh>�I:�E���S��R��I{�y&ЍO{�tƹ��c��(MǭEd@���f0�	t!��?�����	�jJ~�4F.�3���y�'m��_�L�>�k�6�!�}IV��E��sڏF����в=�2W$k����3Ie
9�{��%�p����v����S8�Dp����yd� 2h<�����j���]�?���RctP�r֤^h�������u����xK�F��l���<x
LM`~v�A�rC_��
�*��:身�E�5	�iL���%nt�`.Я���>�x��ޙp���5ۖ��t��Yޚȿ ��<�G�卆��~�p>5���r������� ��K�㈞����Bz���B�YW�Ҡ+w��,Ԟ%����������ٌ�bQ^��Q��Y����Ŗ�ޒuzHm�ױ�T���O0�f ��^��9RP*-���������1KѾ���qR�l�)?�2c� F���g^�,��N�$/>����FU��\��0�Ţf��RlU�\OJp��)���sZ��a�D�\o�A�TX����.ϒH��ə� �D� � jK�~��6����J�ۢv-i�F颶fC�L2x�g@k��y2�2,��	!�4���!F0{'�8}��f:-2b�>/$џju�P���	J`X��sU��Rq.8�