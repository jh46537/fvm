��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�%>��1(-fR�6��Oؽȏ�)���V��L����W�H靠_p�X_ ��6���*��0�V��w9�����������n�j�� ]��}Z��M�������v��mYNZ4wc��W��^Q#��_��ɤCl��x,D�����QN��H�m����w*��nw�n,��lf�'���b�Ն� v�~ƙ��%��FXL#��k�~9�S>К��<�ե���P�ǃ���4�^vʱx�(��}�oW��c+;	�ZJ��$a+)��o2�ˁ��Fn�������L=���E�CO�Go�����J��nB[�eB+p#��NW�����5��f��m�Llg��]G��cMei��I �+WPd����FPcI�tZ�J���;��e��re�Ghtw�ǚv�;��._�v&l6~���o&�ήNh\k�aU<%>N�6�qWU�Wſ�$�p�J'�#GVR�Rs�.pU����a8��Kqշlz�>�.a��N��d���?�yś��,�H��˘	�⮜��r`������	�q��U�ā�Jgi�������5~?&7�0�sGb���g�a����=	����k$���r�/v�1M�����ZF��p;�����*�.�Y/�8����Ӿ`&WX%���C�=Ӂ�d��,،(�S�N�=Q�	/!N3���46���秹���V��%�|��X,QIH@8cka!:"� �c���e�EU��e�'# uY��ǏQm�a�Y�}�JO��A4~�t{J�?��M��@�h݋���Oe.��g�N��RQX���p���u��Z�!H�1ȱ2�§񺞍{C���z\��>�V��Vꖝ�������U���-���ء@@$,5s�.�~*��߾���W�Q��j��g�4)���y�2��$�ёۦmY��T����LU�WJ��]�qꯍ#�����������-S���ľ:�������M�e����F�����N:G�\V���>L~��2g��Se�"7r��A�a�?��7'.G�M�7Yu��g�.XG2\T���U�HdZ�[�	�ϠK?@W���q�k�&]T�	2���d�48&`�oPT3�L�I�����\�l_��C��U����j|�����f�v�]���KČ@$��FT���Z��>����-�k�*��v���+co���a'뮦��ʎg���
�HM�~����Co�;R���;�a�3�$Ӓ��gJ7t�]� �[�ȩVC]�����L�(�����5j_y��� �&'��0� �Z��u
�>@�j�\�Q{�J�ĸe�4.�U���ס
�±�,���M����p��8��!Pz�F �x
̓��=�:�7(�4��R�f��^0���H�@���h�8����֋F�S@��R��=�6��[闫��)0�]�y��r�%A����IPt��ۭRw��Խ����vb-�� �&���.n������N8
x�a��%`K��@c7���u�c v%��Y����K�	Ǩ'9�n(N;Wx��V��F��D�N�t����X�4��N�7ꛚMZ ���U>G�{Y6Y���Nd�����!���`鎛I`5�$���cx<.�
����b��R\U���,"5CeT8��i�P*H>�v׿`���Y�� ���/O�E��$J�O_�I��7��.��^��P#(��J�E��Ν�\��vS��PÌ��K!g)AB?�-�`�Ϻ��gyh�U �5ʱ�����"��� /
�Կ�S�"
�7z��C���O��L���%j�,�4��HOOM��[�D=���['>�"�3�/�L���G���>΄y&�cC���ޯ��Zzž�E�ܧ���on{p��-w񺶎Z}f9�M!���H�Ik��c���:���y �����PsS�tk���;���ar�uY
i,
<�}�X�` v-�HT#i�ˎ�Y��27���'I�U�N�u
�7e��F���V !�VV�Z P�:�Ct����/��5�*SW�� �vi���_��������tu�p>�����O��d#��#]��=��U����ȿY*J�#��MǶ&+��<�W�~fO���_3��I��j�0PA�܄�����KY#�c<��ԙH��B3*��HdJ@�d;ה%4�T2�s�4�����`^
�t��Ç�3e�Kh�ш��1�7�ge}�~
�L&�Ҕ9�E�� �m)rEp�d�:I�=��v\��l��Zx����K(�Xɔ���tMqzt|�y:O�?<f��~tMȖ����j�y��پ��XT#t4E��_Q��I��W�TbDco��A�lXQ{�'V8�3�0�������*��&�� �3���A�2�l�������l.���NT:/�������Ǐ�k��/�w��<�F�]59���<t�.��N���|���E�OA2�#�M�H
�� ��=���8�Y� �3��-)X�;-kN�k[43��$��8<`��_��~\�� iR]$6+i��̦]������i(��rW��{�����_h4�˷�S��_jZ?�
oч��j�XQ6��v��ӛ �uAu���=u���e�����:��+��+x?ª��=} y��󸽘L~��zyz&ECh�I+;�S������o
���f��X^p��)A�a��
�%;S��EL��}g�d�C�Q2r��B?��aM�[��n�d�G���fP�yA*�n�X��=�[�#��eQ-d�F�>��U-��e6���/^���<87K?G�g�2�ls�H�l|C����ћ�z��D��pp��$��� u��η�l����+�n+�����$��(nuV��������!r�IF~wt?*���`�<X|���x//�+ּ7v�Hv���w��S�����f���Ӯ9�D�Q{��eU����(u���{�,�24�B���
�����!k�p0���zJЩ<�%�c}�����Z���k������|c����3��2�v{[1�4��S���$��a�ed1��{ݼ�=*�+w�I_!7Z`��������b�n�S�(b�Lk����镖X�������Z��@BMxZ�:�B��.�-Vo��l�՞��wd[V�DX�	x�pzK�ҽ��s:D$��^�x�x�t6���O[@�"�#rb,;۝��x�wb��� b�]��a�$@�v (cO��¥ʀ<�����n������L�#�9��Ļ����ci���a�6q�9���
�g��n BV�v{�dWu�ٮ:YR��<���r���~�bm��m#��]8����&`��p@ac�-�Ϭ��[e�I?8�(á���`�q(6�ޑ�7T=Sa{QS}�s��(�	?�1�M4�/�nj���N���C(�G7�ah7��o��b(�Q_̋���Αܤˍ�t6(u�pD/a��F���&+i�3�t����k����������Th5�T~ ^|ç�Gk�E`���2;i�do��8%�-k<S�"�=���mY�P�f�>ܺ^���A�I��R��LI�k�:jE�H��3f���`;YY�m�;��|듒�����$1]Hu��ǘ&6���BME\�@Z;OK���,��c��B؆�\oآ>����y��"vY�u4��E0�zy�%���R�Hv�&�l�b"�|�d	Λ���J�j��I�	�ݭ���k�J�CwˡԱ���pm9۳n�� wT�����S�}T��d1��۔-�A���s8^'�Q C}�4�'��ʝ:�͕ؼ�JF��@����~����<�a��h��m�q�� �{�-׵�pU��P��Ah$�4��)R�o|��(Xᘺ��i3��=�������)��<(���F��oXн4�U�^(z^V�'�GQ��)�v�Y������J(��i�%��\rkTٻ��%@��抻���9����Dsd'�$�HFix$� [���;�fO��d*�a�V�_,�U�OP{��n��k7
�:�N��+���jb�V�k4a���i@E�l��kc�0'�P���=g�]�x�o������Un�aMs�
�Ǘ=k���G;Y�����0��9k��M���YP�#Fs��R����"D�(g��%'�Ƙ�mp�ε�����izd{Uq�'�+�ݙ��Ȼ6K�%�G(hlZ�l�M��?Շ�,"EFI�b�a
"��mGƶ��X�2m�ه�A�^���w9I
 �J$o�c�
/A�ޱ4uT��0��W���M	M8i(����t� ͵w5Od�"n�(�B��]��i}{���z�V�taS����z�^;����UdV���n+&�g�,��F���`�� �"���M����z|�i�r���Smzc\�M5AK�ũ�-�z����Tlk�EI��Fx��%����	
���3a�[�Aqֿ���3)�'�焷��ɍ�(�M��S���a���؉)�5�,�5>�@��`U��q)}%Wxh�t{�S�dL�I�m(�um�TN��{���@�������IZ�d9���Pe���끦�$�����ˋ�c����h,�Ԏ�UQ]�f(&^ov;T�,HH�Q�a�"�3fQ�I���5��L�~ł��1R/����H��C��wt�I҅�d�������Ǽ�4g`^:��8u=S���$�7�;�gML\h�ؿ����y�g�o�a�|��zY�)���2T��)m�bn�������A��yv���=	z�r�Cf��������F�a�X�X���d����!{��X��Mї���1�p�:�=-OT�����_E6�<�W� �
Ϟ��o��� $�/�VׁJ��ō���4Vz� �q������$Z����c'�e;�j?�i
�x%��8 �t4ۜ��]P�j-�~�)�I�S-���! :��p����}�3p���޴Y�@�3�c����y��
�^����5�G���>KY���+����I�W�����H\V���E�,>�'�J��ʙ)%G-?� 
~ֽ�_�ϩ(Q.\d>K���,d�@��=7���	BTw��]�2V49U���d�bAt�V�B9�/d�K��S�e��{Q�L5�P(�=����WLsm�V7��R��?�����w�⻡��h�G���߲|�mw= ��