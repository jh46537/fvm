��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�~��"yAfEi�)�����B
��۩C4JA?ϋ���n����g�ҕ8[���!�܅r(�=����UG�O((�K�`�0�t�s��hP�D)�w�xJ�[K_
�ԈYJ���LݷV�2�콷iF���}Kq�I�q��h���H�i���m�����-�bH1�)��Z�ٍ�jӰtr˥V�ڥ��L���|��qѷ�&GDq��ʻ<�����n �Ꝿ��d�T�\j.+�wH^E����C�]��b��`g���[~?Ӷ/�}3�oN��ѭc�2!	�PC������B�+q�z��*����� ��z^˥���ER�J��d �-+T��o�9��h�:V�%|�]�i�E�GJ��4�G�xn�XV�Gü�g�4�a�K����ѥZ5j#��T$3�"��!��K�jt�%�8��2�Rk�h�ﾃ�!����sR�����:i|��*<Y���Q�"���֊�}�e���/2�yaȾJi��	����K���`�kB����R���\�|�F4'<sSBA�E�J�
�`O��/� �<�S-��S����Gǩ.M�F�^Ǉߍ@=t[�TO����K�,�g&1�.<Jb^`X_ȳ����~������g�R�A��cP�i��]t!]݋��2�h�A:�%	~B��YR�?���(�9�z�vЈ�p�/4�

I��4�F�oE[H�;F���,���̕��[���E~+2�]��&������T�֭4"�XuOG���5̱�)W���eZƠ>��y��v���?n��&����gδ˲�7ϧ�K�?��f�H�Ň���d[m87쀨X��.\�.��zNߟ������	��;��zvAn\���&�U6ϷJ���e�- �L{&6�DG��:!�C��U�i���4�T�F��Ҋ�?*���D]�E�Ls�Ӿ]���l�U�� ��j�D�o�2����Љ��$ ?J�``J8�[�h�����e����Ϣ�5&_��s�N��>Cn#5��6�p�iI�O��v�����P@1�m��G���OM�ݟN��%��{rG眎tQs%�&�C��6һ��{tU����\�.	��	v잡"�ֹ����gl��Qh���n�|�����i���5(ݏ�t��|�����1�J@.~�I���NM�1�x�(o�!�Rۿa� a��K�]I"q~�wp���TC&�*V�&�US�3�2M�j�d��-׼?y�� O�fmI}X�?�	�d�R ��A�cUᣐln������D�ч	����nHM�w6��C�Ħ�^����
}S�AM�a� �Y���o��;>�(
1�'�Tp����^W�KWB���3��N���(������ >Y�O ���O(�h;6�x���"Gv�g�WT'!~VK\3�e�����_��"��|Kk��9�K�T��TeP jdS֕����'�Q7�� �iis�'i��rYyD��1BS���m�WB�����`�Rљdo}wTU�E�H�|�N��d�8|�+���D&���k��-,�u�tX��O�<�{F��Oab��a�Ȉ$�ȁ�K��/��X�vM����>����iľ�q��9�a�Η�O"����T��B�����Wm���퇬PV��@E�O�P�c���=�Rt�z��n�-�~X��o�N����}V/e�����o^/�̘�E����&�叄y�2ǟ�]�`O��zao}�w�>���a��mNE?	J�\�+���GACM�#��Ҁ��bIRoz��=�%�
|;���(�9��gl�m����b�x��gl�H:�r����5���:�b��TT'd�f}���2���u�1Z�Z�o�ib�*4�^t�����b2*x�| ����~�*Y
���RO�C10��'��:�$Ë ��K����U�҇m}|��A��0o����#Ċ=V�١�ל�@�	en���d����3\�l�]�&��*`��z�������e�T�A���N���lN�d�\�9_�����4�������K+��$���ɤ��P-�������
K!cv�2d󎓬��vn����a�AGG������q��(|g�4��H�Ƞ�iO�;-�k�i8�D���9O�������Ӣ�D@�-�ߠ�fBs�9���찏 oU��~ߩ��Q��=�B��~�3<~���e�(��z�	>�"l�
�!���H�ʚI���D;L�j���ʷ��:�����g&a�_ؾv�#�Lu]ʋY�pz��A*�,�ˁ.*�g�#�Ӹ�1\T���<&�酀d:�w�d�Cܫ=ؘW�`�K���mo�e�b�:��-� I��*:��R��r@4훼s�]Y����>��%����;���^�����X�|)�J��ю����/����sz�@-`��R'(ו�(�aF^X8|j�j4����	�M|�8_�s����t����0��8˸@���$�`5�T�4=�}�n�1i`�#"=��E>8U�6E��Tqϯ��#ܡ�Ab:-6��w����6�=���j���܌/2}7'���D]	�i �;ǿ��yEH������/�qu��L1`�J��~I�i��lr�5��=��O�Di�)���l񦳽����݊̂������w5lC�F����~�9�q$c�Bu^S\{AҪQ�@��@��8��O�vɔ�%d�&;'��	v��\,Q�b{�y����&e���T�������5�ľ��� |�m~�e����)x�2�+�s�L��7�Ԅ����Z��z;��4�ԃ��8��5���`��畋����6)^�Ί?2+���
��`�c��?�ruv�����K�f�N��[V��ꉂM-�o�.x�Ό$���5U~��8�"��Д�o�H�������4D�J'��T�>>��������<�p��۳BzVB���1�	�3X�Q�L���>�q���=��&�m��$U�d>�T�a:K\9�wF��v�J���#n������c�}��X�$g3��w�A����əGIN+�e�|.Y��#��M�h\����$���t�|LԖ9OFP�<�g��qe�˅�d��"�v�̜CXs+�"��:��Y�w��x64_����Pf��eG]�v/r���-�q��r2˂��A�
V���G8��~�.�|�M��v"X0t2�L�/��p�J��.��I˴���Rn䵔�W<��\a�]x��\aO�������qi�v�Eg+�� �o�f��D�ǛHT՗~���#:��X�lg�)v��3ղl���\�,�`�b� +� e���h3m������غVOY���<�V�}�|A2���|M�ev���aI!���J�ğ��J����\�J�e`�p��M����Yү���G�4N�&��"�	Tg^̖ND�e��x&��W���o���!�����M���L"�V�Ȟn�7�,_kYzvAd�r!v�~ᰦ9��փ����;�vKS�T���r��W��.��xK2K���&v��K���B�V ���&�D;�������*A�{��f���4^���9��|��Z tq�$몑J,%,�N�X�=�_�oE~�5_��<�ǃ-oX �L��:9̲ȳ��Qu�d����l?�yE�̭c~��&�&���6�w�*%R����ba���<��t�IT��2�_�'��.\[��w��������x��ʗ��F(L�=�,�.�c:Ex�����vb�����@�eW��ɞov�)��j(,��kH�{��N�`�����!�oݰ�.ը�"��Zʔ�%����۲<6I&�GT͡�ܩlQR�)��Mp�uK/QN���#6{V�|-�c5��m�����Y����XW@�(�[���3�L��aa�a��er$5l�:���P�ATJ�C�#I�c�'�i����M��p�2n!�m���:��4ҥ���e�mQߝN։l�!#��	�����BP�B�fH_2	�y��}e����B�
U���2\լ���hp�kW����噕q��Q0ѾJr���R�i����P�ܺ�A�I�٨��uQ�;t�[ �5����A��p''s�Nm�e����_����@ث2|3Y\8#� ��x�BL��?�,�sȠ��z�$Vu|�Dm��(r��yT�RdI/���Է�Dnl��gg�tF�Gm����I��#5"*|՟<�Q�%-�7�	����8�-�+���Тs*ʋ��J�H߄�ݞ�F���ӧVLB�#UEKU����û�i�t�� xF�W�|n=-$n(r�J$|��'uEq�j5�7�v�A�� ��D`��#o��@,�I�0h:F��\�RBy��	�躄�������OT���$�s�-��[Y�z�ՎO�fV��1fr�Z��G[�fX��R|�ܭ���1���UKl������SxТ�"`&����GMݹN�%�r�u)�fb�k�q)�m|�J�!t���������H��$��6��K�<��,�qg�S�'�<ϙ�Pbww�b�/q��s��Y�X�y	�˵jõM��Ĩm��b@�y���A�$G���X1��ͥ����a݌8P<b�2q�M��b��P����J�J�iN�%��?������I�W��`�LК
(�1���RZ�lt/�r�i�'=� l�Ĳ2x�� 8)��ե�3L�J���B��N�mO�y�ˇL�"���6��\�e�A���=/0�B�������s����������.�R� ���3���	��竱���xf�����{��ڝFcևq�W-,��C�23w�X���"�]�f*A�is��:1K|!&=�֕���S�0GqS֤(,�_��7��K�!^��I���B���Pր��J��+X�<e-S�K3/J�i���ß�����Ɖ��9A~�c���[��K��W:��,v`��!iB!.��3��t�nhh��� ��7��Ú�?�nwr� F(��_9�քJ[VJ�t��FE�3���iL��-b�⡲6��gnX墪M�oil���o�J�s��%�)Ό�~�{�h5Mva��Wl<��7���o7)�K¸��k^i9�y#^|�na���%�a2HnY໅�<�[�]�A�m�`���Π7����`nd��3U����WG�aAs$G�pX��9LΊ[��W�Usn"z��p&�E�<�I��1;�de/����썪�S�����:�M��y��mb9�+�q��F�LgSql\���ovo���+�۶]�յ�ٰ�aJ��o��y���m�J@ڪ��+!�h�#
O(��#����"sK
J�+
��R�
(.�A�m�T��l������Z��%_(�t��f�f�B9�����ʻp�HR����<�gb��B�UU!��L
�f����s�'6�k�2�@`��D�U#�M�v^-�M�t�РT�`V淸%�A�>���0Ժd�v��=��`J�|�)�`톄��+�$���XU,����QU��eɭ��;�5�����@�h) �'f��qM���'00�'�<�y��~(����K�q�q�V�B��Y�j�����ѹ� =#�V~@�3B����`�\�	�?�D�V>��+�vC"�mS���Y��Y(
G���Yd����C��L�a�X� e���ٞ�F�	���!7r�_3� ��=	k3�}V ��ͻ:�����8Y����d�{��w8�������;[��y�.8��ӝ�_fv�M̐ ���� hy9�2���<{����ݍ�p��yJw���5�MӐ�q��~�h��?&�"C/t�W���׮�粵pa,�y��e�y�{�ߝ+5ǡ�*�!�e�J[�Т?
�X�d����yV�@�g�]�T��ʅ�Kj@Y�� ���q��]3O�W"�hd��E2���ƾ!aI�� ���R�{��
��V���o�jxb�7L��a��{sx��7�Ԍv�����Ͷ�����p
k�4f���\j��
�0�p��&u���!�(��3�$��_1�	
�5l���$�*����%�w�sn99��'����8*	];#�a\Ś���� -u��c%���7G�W"wV.-�]Q*���'�r�&В�J�����,�.�y���{���;�����A�|7I�Lws�ϠJ�D<����s����0?��l����I��?���n�2�=�	�ӗ-DA7Y�^9#�u�X�ox�a\"Ĺ"���8`{�v��捪�p&6�UV���.T�n�� �1��JK�1��BP�u���L���%�1����ʬA��j�m4g��P�Բb�}��w.�T������@���>"N����w�I7�4ܸbc��� %����o~.;�~�\8da�K�蛎!�U�ٻ��'�|��"�G�c�A�sĮ�
ԁ �������8���n���8�&sLD�A̭k5	n�$����<)RZC�&T��+p�tVJ�cu�˦�;a�@Ղ�W�.�Q�+�	�}UF��v{'��J�.�N�~;�3�K6��9��1�@O�6��������p��!������k\'����p�L.�����"{9?f�B���#�Ƽ�ф������� �9��:
�9��?�A\�W�6��CsC���	��x�R6�������_8�+�̕�LH!i���_+A��&V�4eY�.�����K�+������/f�=����ه���'���v�h<i�Y�H8��)DNZ�?�C�o∙��?UJ/��o�2�V�؈�r+��Nq6��,3�au�ݳ(#1�{��0��%����8W)����_t�p�E�G��-=i��\�$D/��nk�~%�?9�+o��ʫn�(�b#����J O������o��"t�b.y�ǭ�U%6u��jpZ��}'�%H�|`��>η���X�������@l�8��8�ﱰp�N��o�X� �G��U��<i�lm�� �������F�)=��ڠB�=R���-zȺ-��r߽�hzEY�߽eM�A�?r�%�ڊB|�]�k�i���5�[�g�Ŗ x�8:D[� ��j �,f,]&� }r3O�Ri7��mf�_4�X��Euz �b��q�
��#�؀�i⸣W"$�����vk�yJ���Y�m��ù`�� ���>'w�-n��a�0��#1����ju��ӌ�x찱P��� �zUc�q�v��DK#�H$2n�q��4'}���ǠoQ>7�1��>���CzU��ˣpرP��4q.3,8�=��(^�A��6o���f�{���;���E���h4ܘ�M_�!���7��OJ
��)�>�ǣ�m�bfjE��hH�ƳA��r!wr��?��+J̙��-�"IS	u����ɭ4:B.�!��%C�z�O6�6��}���f�����>�N��h2�p��"���[P�2p���D�M�%W�T�z���R]��w��N�*/�׍*�O��q��B��g�ڒr��4�,�YN���⢙��E�P��ǠO��/��_��,�8�"��[V��};"��QU�A��	��wɾ>�g�'M��(���Y��߇޲23���P��D5�ǗqQ�˓�T����Jî��J�^o!�RU��n�?r���:3�����m� Q@�Qo�>�Qk�:U�Mj�������1:f$rP���k���U[V�h+8Y���Л�Y�<��Jŋ+�*i�l?�T_H�d�]N|�%H{`��NCd*G��Z�I7/&�#���/���;��u^��P<����A��yͩS�`q���4�P��#]&	�d�zA��9���}H�i�r�
`g}t���+��褑)��П3VM�z����l�r�u6Õ݉���1��|F��?�oq^$9������_��_�ۨ�BN9��4@�`v��{�"W�����о��p�I�|����+��o4G��2B8A�&>�+p��^f�4�:��{��ٳh�љGC�z�Y3'q!o&�����E{ļ��ȩ��M����Tlg
}2�׋�����P��� 8���r�)t��d����?��l�o��%9�)��
%E'[�}�i�c7�OfS�U�֥e�[�N9K�E��o| ��,W�w2<r��k�j�u������sp�S��߮c�58إ�C��j� �_�PZ��jq))�pZ�� �-�g�%Im�d���گ�u`��Q�Q��GaGG(���$�,�m��dc�P�����7r�٬�C[h{�n]C�S��KJ�s�D�L�)�Tǣ观I�8~��Ly���9T�G�`��(٣͠|�Eth�C��b�<��cl U1���)_EҌ���U�j��z�Gɋ��^0喝�S��|��X�a��#s�+�-_�b�V����c��FL`um�R\���'�1��!�*����t@�حd��w�ߜ�R�"���4z�(Ǩ�V"�`\)g�aWu�X��Ғ_��r�ht��=�*�pt܂���������#���|ε�ؚ�_�I���7,���(��,�q물'A�ߜ�k�}�Dlu?[��eG9�R�O]]�waC�#I\n �^�x
���X��˹�����{�D�28%t-�~=�EXniL
�[���&�0��L�T����&r$�]��>��("e%��-�/<~ ��g�Zzi��h�M��n����JAf����-4a�i������d�U��ۋ5 � ���7���S����b`����繑���f�נ&�O
�vA��uvȢ�)ad�Ҝ�C�oJ�Ny�׾Axa���#!�(��Y
a�Q-v��+�*v�\����k� a��+V�"�V!���"3> ��>��J�ξ����Ш)M���4#�$�L��>���������;�YW��)��F���Ȁ0u_L�yNf�)��L��b!μ/�ݜ�R�.�r9��K?�]�c{~V�9�5j������>��|�J4�M ��Ԯ�i�P�E��΋B�2���i>��M�s�4Z��.o���o�F(	�l<:?�!�a��=>`���s-K��k�͒�J���.(�E�x�B�&���0ҎI���
\�Ū ��{y���Ίt�|sJ�3�.�A�z�,Э�p�l��n�\|�p��ˢ�*�a��|{<��:ӽ<�+�V�@
G=��X��w�?R��%�:/:^]⌆昐���2����cQdlr���p�U�;�Q��ʬ�4ԯ�ר�3���郩r3�D�sR�"��١]���`���Q���ea�:�*GF�3y�y�)��T4���ȳF$�-���s��c_(2;��Y�5/u����kV�3Ga�¸��3�4�GB5p(wv���rn��N�5�8�|��'��Ð�䉮�.�bn����Xٿ�y����Kr&�l_��)��Yl��S]a�g�*�M���{�����ٳ	`<iDVb�����0�B��\8BF�i��7ǟ5M��`yu.NJc�1�r�7ֲ�q)+J�f�Yg��Qװ�K@�=p-��fzxH����ӆ	�Y'�'yu��gQ��)|����j��4��2`N��?O���,V�+u����g�S&���tz� ֚��������=��3��HdgKe&9j�����3D+=KM�T�I�\@�E�)�J̟�2[tXث})���|�K*"	R������6�h �T��Ln���h��ض> D�����k��*�؏�����P޶}�t�a �]�x56��A���(��@	@��	��L��՜3O�l<�
'B�$�aY���1m�8=�<S�S�d��4V��r�}�?�����z���-���$,��;��d
̡�eC��O6�&��{�5�[�@��q��\#�E�4~�F�wW�o�b¶���Yy�� ��6�������	�ASUlp��d���ͧ%������̿����逴����W�bh�Qؕ���F\��eP=�R��hүC�<�����ա�=g��r���w�J0�ٙ�-&�{�~�eV�ca�W)
���G��u�xE� ��y�,�m:��[��3Ͽ�6�ow�T��,�Ω�MF�Cr���6P��W��'�X����x���zi�P	L��_݀��b.{4�d�C}�M�E�G��Qa�Z�	�F:?�7��49�̴�
w4��/��}�vMkE?�=9�Y	a��'L'i������.p!��s"4!?���a��� +`�sv�3k�|���B�.+��?��EO�?C����`D/'=h��Z�C���
�V��Aհ��vJ��!ǀ]"�l����1�5Xʢ5�w׮����8�:e�G	��»O	�_�/`�l9�@��n��� L��fo>.lb�{�>H1Z�9z!�>���0���*���Y������L1����_���oy��ڊ-���@�?3��dh��(�
�Ij�5�.�>d̗�OV��氘��&��>[*T�ۑoC�M,��i�1R+�<�]��{�Iv��Cw�+?��w9�u�	�X�H��)�:Qf�ך���wIF��s4��p�$�b�9r#�D�6������
�x$��oU�!�Mb�Yk�����W�	�1��ULn�D���R�-0h8PT�)L3eU�VE� ��̂�����3��K� E�C}�Ǉ��x���eg:��
tw�M����gG3� l�6���Ȕ��w��9�-kzu<9o2����)���X�;�=B��Bh�L�/M�2$�0��i��}�r�L��B[��2e۴��O��� �
�}�6��J�Y�.���N���*NIY]7��Tc���Z{_hp�"g~g+A��H�~�mk2?o�+x!�w�@�ya)%���:b���@��Q�� �K6��P���ȱZ�
v���Ə���f�V4�=s�W�˼nc�_�ض�m��2m� pgG����-�\7�H�&i�Ά�7��u��=@YiK��,�E���V�6����pd���w���b��{n�J���w�D�j��G�b�1�/�L@:��u�@(h�m�DK	A�,��U�����A���_Q�ɯ��=ɘpԤ6�=R��"�ŷ��bDj)�z�y}��Fw��!��S[���1�p���7�=q��݋L>=W��?۾ߴʢ����rj�\Z
���W{��z��V�Q:�#�a�[%��7��<cE8�7��N��|��	�"�$�!�����������˧<�K��#Em��הE�]t�4n�d=��E��ϸ��ƛ;ʍ�І�ig��I�%������ь<E��g���=:�Uh|��	�����ܫ�C�w���>f�{�n���f�ha��V�1\b�b��7���K/�����^���`3"h�i}$��U5��\oX�G2��k�6E@���������'����'���*F�g�߮l]&�mq�㠚��K�*��B��,ZtXձ_!3i F7�TK�*�]{����G��(��m�v�(�ة"�����x#���W�
I$�mÝ��j�@<1-�:K�|��o��K.V	s��5����P����ߋ����Uq����T��=/�3"�$1����c�8���R�+Y�6�%�����W
����]��C�2�(����U��]|��k?e��(��=	�9���9��6;U䜰Υzt~��-,
�)��liS��/��nD����fR�uS��C�h��3Ǔ}I�%c)5W�"�.���g��VIZ�4uЯTY�Q����?����LÜ�#���~�϶B?�哵S��')�@��h��\h�\�l����í�ro�����Z�ԩ@��s�m��0�����|���B��{�&c�$TA������8�0�F��|���ANg����Umm~x\��|���;�B�jSo�;�����f�Z�cc��<G��V?�z��	ʇځ�0�Z�ϭ�C�O(����A��ۂ;*�T]���Q�yؕQ�T�2��T�������R`e#�mbBCp&ٙ�@�j?�EN�z6ڦ� ��=:���K��̟`Y�󐓥����:�����%$x��`5�Qe���.���T��|��"��֣��]?g��L3o8�j��	�n��ZVT0r���_ھ�.�L}O�$U�?*og��]��uG�l�\�ԂcJG*��r�Me\B��0*���bj���tD������k�𫽭�*�s�?����ֻ3u��Ayf���?֚�1ە�{�H����|�XS]>'���<�3ѵ�F��h���LMm3�U� ����uc ���l���r���\���]��3���Ξ�� `m�J�`x"��&~<@�%o:��xq]��yY���Fln^�ă��K�K�>��z^���b��h�ن� ØM�->$P������ǀ�o�HW�d;�Q4:��	�s��%hQ=1Ub�h�((�}{wЮ�b��X)����������D�̝C�]B��U�w>\�S����C.�U����z�I��cH�)fP�a0�R��b��S��pA/N�����d9tV�VQG��m�rVLh05v���Hv��6ި�+@X���i���Ă�l�0�%δ�ݲ^O�,@#.śV���A�����
}�����j�'��}��ר˂!�r�
��`*�P���i�?�HŊ�ВYN��sx����������1�����V4.o��H-r̲u&�����K�.�!N���_�� �I/g�U�?���(Ud�b_
�5=Ն��W�ȂTjS޽��@[BR���d����Q��Y옓����$��}�]P��d�yNEL�E��<ՌN��I�D]���x���M�;N�J(�&V6�,G��Y�-vi�,��w���3�;N�<�H�zB�=vA�p�';
Ep]�������w�.�;p��q&9Yz�c��{�d<���p[�_��Ŋ����9������ ��p��)�l����g��QY�@�T�`8�J'7�����WYS[{�,� ǀ���)�۶�H��~_tW\�~x�vp�P�j�����!�/X�f�o��
R1����i��6ù�+�fY�t�X��Z��F	z_p�	D���0l�0o���7��Rݽ����'C�$���M��}�c�}r`�4t�_��Bx��8��=*��w����Ty<�_
��ٶ�K�������M�7��X*Ή8�agp�֩nA�'k! ���o���Tزۅ&!�0�MkJ��AϹ٧�T�C�G�DzL*���|Fy��G"4f���z�S��1!�)�|��+fu�֢U���UAe�M�j˕q��EFeG A��MCЫ�������bؤ�[��H݇DI��(�g�nN����ʠ��Bi��Tѵ�6%]�vX��`����{<�s�+�LoT2KQ=�Ի��%wY�;��!���БL��:�}���I��7�b>W�{c�k
b���Dc"�/�U��i򨆩���m ���'&��W)�����s=�޲��ρq��_}�J���!�^�/�����i̙:�%2_���Qs�����򟓻��eIj��Y�ދ���iP��9`��<ʨq/�v�w�2�D<"���?���ߖ��A��#dXq�C�q�ܧ�s 3 �w���Y�*�7�1W��*�-	+�Ah��Fx�8�Fkdpk?x�k���N�ņ��r�ů�В��;���܇rȭh�O�KV�R���Z���A,��Q>� ��濸�}�tXk_m���bh㻽�r��UP�k���d�R��_e���U����ZMy��P�d���g�F[�-��<�?J�WB_kB{MR��áK��O�*/Ҟ�B��^�*�p]Sc�-���N��L�ӿL�ą����])+�v�f��μ��v�,�*N��ٓK�[�X������D��S��C�Aa7¢�v;]!_�����Y��Z}�f5vp7��&�B@	_�e����&f�7���2�Af�� ��ܚ&b�PV`0��1,Qgd����0uK�d�����@,N������yR2�r�|�S!��q�/��(��.�F�3�$���fy�4���-�r	�GM�q�^=[5*���¦��BS�%ں�(�^��?���Ho�r���oo/�~wf�eZ���ս����:����,�uˡ��Ô�Ƹ�c���촲WZ/`��H����?��p�7�!��73_.����ܸ�L�y�)�Y�o��٩y�L%��8ϛ�#m?�e!��߃ܱK{�k�$���4�y5�(�Fa�%um�<~rqstRS(���Ꚕcж(�Z��F	Y��2�C�0I
�)��^�9'����O�!�ۉ�E�s�p&@|C��C�e�X�f�?�r�k?l��3��x�2�YEгUg��h�a�k�\Zq�p=4�m]���-��e�_�F�ܖ���x��0�%!�{�8T	���@s}򈄡���Ba}ه�~�g���c����M㚫qe�� �!u�g&��ⴣ<�6�<r&�ۼ���y��9?/K�۹��+�>�"£Ʈ�����������Z���?�,�"YA���*�1�Ȫ
��t(�r��ބ�bsF�=�	2�@��5�;���((�P�O��G �����|����8y�^���m}陭��+Hx�o��ܚ��@��_h�4��S{���:���� \M��X��A+����H+\�iix֒�c��Q