// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:43:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Pl5xwcM/jKHJ7GVwDvtlHyW6PVaCnhaw+0rmW9qxCAhBIXlou81oQB6IaiB5ZX/7
deq2vhgPxwNWD5aMejCbYILZCLmld76jZp7cfjUODz8wlQ5wiO+3Bpxl1ZGQRyGB
Jy33mOYflw9UBxG3QcwUobVTBs53RNyFsHRQcNwp3dc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5120)
dpYOqb2S8XSrXcHT2XyoYChsWUotYoTYLFAv3fPAoeldSMzSnsf5ZlsTKHGpfwMf
C4ZwycvvoYCdLAH3YypH+NruZi4F6ywPrLvCL9IjxH1zsOv33z429p0sRi7fpjqs
jsXo2n33xUwm2VdZ+t13YM48HSWwCxdewAxGTS6LBqS55sI78iffmlNVi/1C/KM0
iWpf8Cbz8wdvk156Z5UkT6kjEeLNRrqaXIE9zGtz8oJDRlyPnLcqv8yPhCwwhw+1
8bB6dXZeyCIN9t44ssNHytnpCz92aDnJQKxr/1aSC/yVSxLqhQIzSZXsna125Ct8
uz77t4GMqnhMqZHUaBjSWTtvZwzpl3M7EH5WnJu52P+L9P88ZlJ6Irl4kW3rbvcn
2B5EYGxdnM2ooSukvOJv5unATpckv+fUB9EiQzVg0tZwEy9sH5GXoAzfwKoJwz6i
9QZlsvDFcAj+pDVBwPvfiZM/+vqJmKtdWMDj2BpsDzib3aWddnEic+8YlMjE7G1+
9jqFpSjobc8T+Lh9aVJRx5a/1+RABIpH94MKkJrQp6I3Y2YoCUEgLdDCRN4vOA9T
pxfn7FBTsmNWl9Uffuu7X+bBW3vbNFOArU2+XNysO9nQvj2gnRx8FDvy/YmNwcHv
kML+Iv3vRGpSEYqpOpM/9ZJ76hl+wVUbtmbrRvGbmOL6T9rbtA8Mwoxtdnqaig/A
6wU6XnWoqx8Sbi60A1AEcxhXrg0ivauOzlbsqIMEqsw6IhpZr7BIxRORjoGnoNQ1
HYD5ahlHm+yA2BkmGXDtVtzYpzj5Ann/bLqudA74yb4JxEztTLh+wKrFr1JPZwO8
nd4T/qlYyKJ38phdLT1Dbs72F3ITxy6GfPMxgpzfgJysBbFoAaBWS/JwLQYXuZfk
n4EzUO/Thlhzdu62/UIFVdqfkXo6dmNcXDIjabA6FxpAo0GfW7uCOKLGbkwUSpBq
NJ1SG1OEvZsF7p9yrrl3koZLV2eb0H9wKlzT76evQZJA010Ukv+lAyJ+aIO6uUx5
9fhC0IGE9qPIW4zowzmbxlU6T+GmQU8MY9xCLSCj+eXG0w4itt7fmQ4THk2jYNxH
fLx1SrnVNVcv0ihHcQfsWX/3Am3P7eKIXvggXUMIYkyUCVFCSP2lPLYPnXmY3iBX
p04Gay+ix1qcyXrLdnxPrY9mCSt5Q1y/bCyTGU5PCgfq+vA30LnPS7f9YU7ou6jh
UAVoHuzlSM4msgYghncIOwhS4omFgThmHkiHqzRffKKfK5queSkwMFYCqd/fB6V0
2O4Huurn1vxw5mUarHlhlZ5HyDm1Sbn7IiRhaPHGCJBw8gm/TsbgaXXEzyXYIFrm
sYXRBhu9yPaLDJXHwwxC41lVKCplMJkPXRC528PYmXmNpVhrljFPoFSlsm4jc7tS
azohEIKyPnD6Gpw3BcohZ0tlNTYkJ9FQwoG2wKbosdloc9bwR1+jQMRay2B9onCG
wlkQK5gUMFI/GgOsM9h/i8ay9NKHx+fCaPr2fBjxEMff9XzXv8KheOuADCfE7ng6
Bg9A3343ciQmv9SwbwCeRwqfwIbzg7NedU4QbaFANYX97dmHMIgqigemdy11U9Ao
F/18pLsOg1JR0j2iHMrASvnhJx9OCn7QgaRqOTWtW7FjqIuYQqbahaLMyML34QiP
3JA/NU4rHrCBKpkijeoYtEcCFsW7diIKyvTscXFySRxsKwREZ528iUOnmmWNiL6y
8tZiqLvl3/g+5p3X1cQYYpYPu6GVC90RGiOQDYQyN39cDleM0ik50pEwt78u+Bzm
17K/rxXj3RSRRW97krrx/MlEQLQeM3zwvlOPXNXysfklHaHoIqAseuNMe++UZ/zf
inuwTC+dGthyyQeJ0f02ai12gsq0Gng+xJ+xDmkqrU4MdjzMDRPCR4p17DIZoWOt
ISPzV0ZGZb9QUY3Lzm5nOjTPj0vEE6c2M5S4vgJkiTbBs1P4DDwyVNB3D6bEGuQM
RHPU+DMSJFK/KQE01b6UWWg5mdpbInPuelvvQtO9Ire6OoK7X9RWihmQkR4pxXsb
xOD3AUFvyLJjYH6tORfPkoILZcSEq1IVicaEEtUm2da8yJ4FS0W/m7J5gxzO7fT9
9b1VHwOudHD0RoVKP8TIwrHj/ByJ4JkYl7ZpQf/VHx7T0PKpzKKkHJ1QMgP2OvFP
HxVPmxs+F7OmxYl6dUTIbhlYDVc0AyWRzB0L+ZKJEoPiyGGgOqe19ARaa3Okojru
7ghfEeOiqH932ZNt5AA7O3xq409EIaGW14ZGhuWNANBpHnk/dTbWPkw72TDsDgwq
tRVvy+ogEBFvt6zMCFcT2QW69iN03vfGDOFYdtLcT9o2tr8wUqpz7s0/NJ1xSkL2
v7BSFkILgW4Elzah6Ii2QEYs8sMhxRhtYUQa74j0flhEcb+YRxzzAP+XAZaxtKor
09lqVb+2G76YUpGVfq1m9Pil0nJkNXfTY/fkGtRJywEBsyFOOlBJnrAAHWdDAgRb
afRl9nHdNQADNud4gw9GWuOArdTwick801iPKDL5K6zkZzKfQerep5e1yuOVO1VL
7IE6QhPwL6ojSHgF8cGDAk0T0sLlSrPLeNsJksHKy9tV58ic4emnjmxl16egrOME
m7FhIIgEKl9mZHIYgqzzA/f6oLnJ0K6G2XjU06LVOnLMiZxYyfBRcjnaozplIts5
KZxpHsG+FWRmB2nJ7228axrRtMwNycIUpy8JQbbaWoVBfvtMCV0aWVvyMBwEH6Jf
PcwJSavgNuVAVVBURbVuokuuINgdFQmVTKlvmenjfT0TgbqdW2IdHwxUtDA/ntWI
48lkXW77dz56of+Iw65gerAMTGOfy/ev99WAPP9PoSK9Oj5BDeUyHMIttD4uJdNJ
ijE0HYsH0BNyKYtMPe2TsMQY+w0m+BglZQRIrkhzloqul5eHAhCB5uFQJWzk4TjA
UjPD02VseK5URG7hAa+Q/Xz7w8avapBU18TBgFK8maARHQeeIQVSGVLxuxC4aXEi
oUDtAoyWB7a9WTvpgqo4Uw1WYF05lgNyrrROhu6QBdRIOZCU4vRF0lIxKqEIvk2j
7CEUf00SJZSy2e+kR5qy5Ohxf7rmwASX22HvozxfzgBEz/6YJitOzmCojbacc6vg
np2n2DLac4ADVuAB6T3Rq8i5U/a+w6ZbghajTEiCqHymPOdL2xzMBTSz4q98pJmV
ImkU+YZkpZGw4Am7pEHDdjaxlRoZeqfTsqSpkAUTym2LBwBt0P0klTKBTl3zFQj/
QZKpSuPZNRbeQleoEX/dUamYXvvU8QM5QgoAJ3KIMsMzKUdrgOe4FHpbOhIgp6nK
CbpPABJEchqmIFDEd3rPNWsFKsh4n0ejAzwPSCfUYVr3eZ8wcoQctV+v8buO9lc4
rDxYMMDwZqqkpfnr9VuzScN1eCakZuJv/7thf8qtLoGosHdvo5gE3Z1jSDwV/Fnl
a2IWQZPPL9TI6EEF+BoiGm7RGXQtZnuymQCRKKGTRamMf3gbaB+lQf9onHM4oaY/
DidrINzjTav1WKxlqQHN2nFtUkeC3k+UGLboSYWjKDNmHq2WYV0rycYNpdrx68/H
3nTlxKiqLi7jvfo/gBWDf5DEd5rqEhpjlKmh/jEztyn2iSHCLPdN/uvlEno+RllC
jhfpQ/4z1FS0bFx+547D7+3UV65PNl17PkuProrOi4zKs3lc7Y4NYl1pUND4Rg0o
2y2GguJ/p75TrUcy1yUb6iO+qQsGvoZeot6biot0gD8GqS6GFKggjBaFk1gQbSkd
+sPf2PZt/s+/CNb4alEKaIDyDxlKv7XLegyWYddvbja4lRSg9yR37ZQ9aAJFjKVB
SkrcUcUWjPl4R+6D5vWZI+8uh214JhJN602CREm3um/mnKvq0gA8yYaLpZmOcE1R
4dw6adVKl8jpsaLl+IrlrmPWmn/RDN/G83IHiyLQywIzkfKUfnuwEH3pWnNECAv5
9oVNOX5VKXbfCv/02sjW8mfCqMQBsq0dkotn0gVwBq4P2UqgnyDoeRSBXpq4dpcs
Y8XuLZC2l2dikI566F4ftaiHJEPwZBgheHIh/1beKSaHYMfbRlkcqWcVEC24/p/f
5nw80hymTvVVLqmIHy8rw6PpIaGFmKak7+SA0xwvZVaG0DaSuMfdiZmJnLnNF2Cv
VNV5A67nfPTjEoQBmxuD1fv0drlrpX4ZVNkCsQ88jLO7gRZT7bY6R8Y+Slzgilf+
kW0AuABsArmfXcFne6/Br/uBo8b0LamPfF02rZ+88H/0WLRfgCPLnPNAU5e2g9Pj
Jpd034/IVL/4xnhxXS7qdhLl085yZ4ERW9qIJEZgRy60w1sI7kxo7b7jEff80gKp
+ML0095kgrFIdXPJi7iUvKLCZG28UXPCH8jJ6lD1yENF3m0xx+6qnwnu/3hx25lL
j+eY+Gg4OUrZI59fWETVfO+zMbhDHy4SNw/qvXBBc4ZDHMSriJcu+OihyI4LNIpm
3utoIlZS7Zr4+nzBUwqex0VtVvPfPC36Ba1FjG6IlWVhWrSCDEmp2ExtdIDuWQcY
Xf2Iyznc2+4KGmhE5w+w3nWaEoA+t0dbyAO0kjO8gk2+Hx72WuQGPLphUefOkq42
ytjV7UpDW+No3hBc5fCvVvED24g/C4/BQ6DVVkK9c0INrch5XN6CoP/pn5AFsI90
VVzrhsqMUNJ4Q8JjKqngM2C5luSrcfm98Z7e2K23FW2wisEdKrky5lx8hU61Tam6
oELdPCjYTv4be8tqJ5A7++Rhxwd4XRKXKQcxoAKFwT5xtQI8B0La69SYVdrTnkto
o9JaRvVfTf3+7oGgEGfCBDyJAjt+lJu3dzB81umFQEOLsawg+RpPJClUZhAEyPBE
l7CvCKaWk9rHIn6hwjQqye0hj3aQmAvCX+Lg/9Uk9xQwllFmPGY2BKTdJlRmhZbY
71RQ+eKb+TzdFbryFQs56Y0HFsrtJXTcByUH+mDxG4KkjEOm64NybYAyn95OgZ+Q
Q3WqRMUQXpsLMpF835/07DzU0sr+aGV/PLUxOJrEOy2dkQRm+yWpxDy5yOJKisR/
c9wqv0NZPwGIjKTfQbE6zqJXzAhYdlaZlwXOfRzI/qkBDYX5KYZ0DwYegpBfxTJ+
K5N6lHFcBfxb4IrxgBb8aBjJ2N4wO9rSJz5g+q7nWOUY62KcWhE3cupax4TGV5bM
g+4YzTVe+7YOtYJdEd1DTx+ktr1Zu5gfTKgfxzruIswtCu4bzXwbeXFWOgsF2KZH
iJswFenYj2BpSNxeOe9LNx5/h0cC4EayJNHO7t8mOz2p3R+cFllNx7rVpsy5LZeK
tAh78MC/7IAL5/o4xUz+XNqLhyUX6T+VpnKiKlbdeWh85wYXIdIitpxZ2FwI+MfK
6O11zvZF15f2g1GJG4Pii2QTm08gF3kXoCLLgdOdksCcKU4nF5BO8Zsj9a819hJ8
HVmMUtIj32YyY0cle89PxUMxzqIztzDPACokKtPeMJ8Ao9pTxuDhGr53p5mMnpTQ
R0choGsMrHkqkZKDRVfgoU0WxdbEpzJehmO6bKz1wzuBd8Giy1LEQmrKi0q8ZtT9
XJXZgvhKw/uMqWTtPSNQlruLhvZNTrEir1IRJcMlr3O4p9OcvLodNr66OSfVAbP9
XQXYzA0m1V46g9FSb5U2SkBcsmazlAO6B1SFRbDmyRINl2UiO7tTrnhCiOHOWJzY
AYUt6IYgN0VG2LZ2+i0NCewQOmcfKR25znybUd+SRmDzJiZotGp5Jzqx5vLNip12
bPdiNwZyoVahuwfAomzaZUgme8xT6DxvYIQT03hwkQLd7s/v3RzT+Z92gUa9RO9W
KgKFuxevvQlJshJB1anSjlIPRhzaPd/dM/2H2ODaBKh93T2NsE6u32ck2Z5lxqcc
zhZ7pwEXmSkFWCXHqQq0PCN3ieE1fe348a2L/VuZLtyDFY2nFbg9jSbBRCk4wlxx
QSH7lrlDqKFgla8BtMbROZ0ZeHt8Fpxbk2J6D+g24iwEEzIbHwBCFtP1yAn4B8AU
TedmEIN75QDRC6vhrudHj4fD38ybXYD7l6L+h+ztwv9EDb9vkyRx973LRSg86ElM
uwOXfe7C8Wcr3g5J16ttsH07NMj/y3jxukQTOQuHefig9hGIkDVvP1X1ykeD55AV
6/kjguZO5FrDeHd9lFEPDK8Q2hPwg9XKoogNM0HsnVWfM2wW1K4JlPkMAJQ4dTqy
3vXo0glDKWHCRa/FM+7NNGXt+6TMUSl7CYz/HXz7Jtrjhf4l5bwaFLOttj+slxoG
Eo5aIOH/Lqp+KsdvmdUUywImnKBWqdTWZjvmRmdrpcX3+MeqUp7ivh7XjCwIFNdJ
OO7TK9d5P9fYE6Q0FLvccT26Ds5PdQq+H0Qt+SY5MPY2s6IlHCxNWj/KYGGZLlg1
pghFIV0dyUZgjWFRxThEvuHwgVHx7wquvdzwXDBukSm/inA3m8rYjXOsNKwWH6YK
F4DUI6Ui0YizGfpLSi5qMmIDRIP5PbZNzOgczYrgh2uXlDkkgexUVcKRJrIUfDPh
st8EnZGDFQw7HfadUrOEaaWcly+IFKXeDe0msLXgPP0vhJhWSns7iI0dBzsoQ3zF
noqijOVq3n3SROwE4MzNfco0Ln5n8y6VfYAp3hZYmPhqC6l1jCnKdFiDtAG0QEB8
/uZqwg21rKOmna/CBs3x89cIQT8D/YhiCDRMmOOnFbP6DPmj7pUEn2yG6+8icdEU
SKtM8vYpU2pEuvtkABUMc1zx+btQUZgmPapnJNV7lzc7KRalNj4AuOMik0Q4syQo
o8XHlq0vPDphxyDcHHp1niflLIo+/Trcf1/wBwjUrP4=
`pragma protect end_protected
