��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	����FP`uΪu2άH$Z�ՀA�l}��}���q�z?�pGdmx���AG�"���R��4����d0#4��,��p����+ �]�`��vR�)���G2-��]9��Ǻ̎�]N�²P��1x?09�w25�*�0�Mk�Jμ.xe��^X���s�1k�7�R"<�- ��.,�@HӺ��RC����(d�}�Y�p"���"/Z+��騜�n'K�2}q�4	Ė�o-o��B�|Y���S8�����M'��w%ܗ}��~��A�,���u&�BU����J��5Yk�4+�]��������*"�rxW���0�4]g�$�b)�b�6�Į�c[2鏒�[��c�NV#1���ds�&.$�����J�Z����1Bc]�^��*��<
x5�m����^��j�u��vc�og-���W����y ���Q���.ہd�#A�R쮊�x�����j	��w+��mzf�!}��q�YQ^F�Fe''�&����ٴa�|!҅v>��v�C�����]���20J-cH�H���� f��<�@{�v����돠�!z��i��&+d�i!3�v,/b���<�����]��؃���� �~�y��|��',l	/m�+�``��*��4(���
39�� �P�H�-���YB����.]��lR�,S�O������z��H����͌o��ue��F�z�+����j���f]�B����^����N� ����I?��Ì,���vPN�L w;|j<�H���a��"h���?&�6^�=���~cٞfPs~ķ'*����-x���u�<�F;�U�	�V�	4ϕ�3��j�Y��N��{���	�.��~VG��)�	Yh���;}�Ժ�h��<�;�.1�8�k.e��A=��Q����3���-�P�9��v�$˺hc"ֻ��외�����;��0#&+*r5؞���Z�1?b��:Z��Q2�m�Ѵ�u� W��:��}=.@/�Uֱ�b���Z���V��7��
8	�����oT�%i��@��0�\`�L�s����|�!�G�܄`y��.�%��
Y�2J��d"�"x��>r��۩��� 6�~��
J�o��0X���'���;F�^�V)q��Ȏ���f9� ~t�m@=�$���SOc�4�B�m2&V.@�e�Ɍ�}f�@ٿX9f�
��	1��g�������GN1A��,���v��B����d��9B������Թ�=��(�	5n(�4S����k��<����/K���(�Љ럮�D�°��0����9��DS��L8��8���qB��,4#g0���]!�B�YO~81C6�xK���#Ȏ�Wr���XX�����K��@?���
3���tR_``���p'�7\F=��F{�1C�-�.�x�w ��8e��_�pOE��z4T��p� ~e�6+'�r��8���I��@D
�4o$�P��Sȼ�V)��EO�0r#<t���۪�"Q���I��2'�=t��-�߉	0�,%��s��A_ITu��)a���X�l�A�C�'��l�_8\J��6K ʠ`�*�&!���3 ����_>�&�ؒr�<��8�a� ����e8^��_Y
��%�mD�Z�*��ߴ��w�е�q1�P��\���Mu����I��Y�uIR��,����*|�;e����:���&>\���̃GR����/�Bl�Q�$��{Z�U���7@��Z����6�28���1�s�z���'k���N�����QΥ
g-��M#q���{յ���d�,�S�0g[����-�^2Mq��Gb�^Ʉ
QmwtQ7=�H��x�6��z�l�K焝�$8��W�<��E@���[Vx�Hd��j2��8I�\��r����sT��9:g�m1�Y]w���f�]��O����~\!�ЎOpb�G�"�+��(�c���J�_U��nR/=�N��]�ø��b�f���,d�Q6s�l�D\�ݐg9��Mҹ*�'�����,CC8�:Fr���L%`2��'�3e����c����� �|KE�q�p�ܶ.`pȘ�H�gyR��H�.�/
zk���Iq�</��z/���\�#�˸��r)C�wl\���gOY	�~��A��3�X���6f�Yd��N����ec�� �����0$k/�y�[���MD�|�z�H)r�U��kލ�}�
���xoT�1�J&���ᮔU�i*�/�:f�ٜ�z��"*Lt��|�����,�g2��|��H�9z�� d�bi�[8��.Rː�A��D�wK�椘��Z5�_�[�&�A_#��G�A[y� $��I��a��x�ܙo,�g�_�
(�(A윲*=ǃ�7��M��a3,�{q-�T[�	��׏�}��f������t=�EYd��_X�c����◻�\��|���ά6��i�"v<KP
f�+w B�3>�wo7��q:��W��W%���_���Ư_���H�b
� 31�ybH�y~A����Ii\�Շ��'������ �R�
�f�NI=��uB�J��9=:�f:����E��N�O�xū��=���Θ~K�Ϻ�Qd���0���:���\�$����'!�c9��:����2���J�����yL�	8c�� �Gph1��&a���Z��K�R[^�T����uj��h�>�-k���&��Q�K>�om�֟*�}z�ǚ;���#>���Â4��n�(�#��&��b%��=���LL��]��՘����z���GKY���{}jA�M]����ԅ^΋_M3@Z�+��;M�v.q���)uz�O�.�{���䄺MK0e�ȕ��zf]�i�݉�=�r������濇2�:�Wj���s�\{b�_*q嵯Po��YHk���ǌt����Ix	S�P�
�p�Rl��%#���v���T��vк&�](�F�YDf͓HO^2�x������!&���{�hI�x���E\��֠�fz2��{������Q��&Xz��"�vid���JՕ4�����im�
�v�8���)bՋ�z��<q2� �	�$��A�A����^�jJ�:�T!!���E\��� �g�}�3��&pt�����W�r�����%����ݎ�>�
@�ƣ�\����+r��R���nM�yʠ>XQ�(�)u/���r֤V?+���22�^��a3�ki�Ϗ�h�Y89Iz���rM{��fhx.E�t*���Z��]�;Tm�j�d�h�6����8iV�$�|�����a���U��{>��X��'��&\H�JZY��!�Q;���v��AL� �������Y����qI���3��^�U�����0D �W6�%�������&�dtMQ$ݭf�i\~�c�18�)Hm�}[���
$_[��L�PR/m��Wo~�;0	�r�Zƃ ԟ | ֳrW��+��:	�V8������qHpv-����Ж��}��r�������N^�?�'b���=*zڷv!!��$D��Q��f�T�vxT;O���{YT}2<)zz����4|!ȡ�H�ˤ>l�4�