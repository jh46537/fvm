// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:35 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
o0QM2oc60dwCNcbGYn0Nt3uM+APua/O6/7grVkQkUy1KM5Eo+TKaCmncZJTIio67
7z5Kda3U5ahu0dSlRjkpUi4IbQQbGB/vIQCFSSBA9RCbfiz/1B1C48tQXhFPneEk
VTD5m3E1KQdhlocTn2SORZ/ZMeBHIwaGl1LXZSLIUcI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7200)
cgkdRzFw2ICiW/7JV/AyJ/o8PO6O0fH5EmDi9wP1EYL74hmuyWBWKidrJLELstJz
4fTe4q2thSCJJ1EhqLQzbkWpPiok6uUiQCEpTgdgBj/vq9iLjm2Y6vzKhIBgQSXx
Fk0iczLtomxsWDd/BSL7dL5VMFmNDUzMr+a4zmPs3v8OCISZ4GO58KKU2rWL4KCR
WOO1AhIaMJd0+HrIYpMeckPPKHmnDdenDbLVRUfUtdJvpvyN3VgiHTQX3le2GzOV
koCqyZwc4L3X3DpvR7XuPbzmSq7Ko1lCd7kNiQfjEs79wNFEDlDMpb/Ykt2L0qYj
wcepo/3tzyFMrklebVs8tVNpb906WaK9pMFCGUPP9a+sYciCwZmnPgx7vrR/LAOt
KqMvRn0ZEyOyg/fl0Hq5rJHrZgygqIZuMiuFwZR2gEz7il/audR2kgLM8+/43gQ7
CCWRoDgFL1zru43heipqVINfoZcJ2/OQmJICxxykesg1kfU13dFvBdPoj5BRukLg
Sy7DRenX3ZRfs7+aX4YHWBEBAGIvEG09OmwxfALrRxplsl8Aem1I1j2Xb02QFXEt
UCdW2ACIbFcjeaV5qFNg5N4bQNvY/GfWAGYKeDyO8F3GPsxEehEND3KsGJ1McOxW
t4m5LbT21MPh7J5umgFJ9f5cW8GnGiJmJEm3wJDDFRdjYmIN94IJ4aLn5OY4NwGN
3Pw8R+CBRGXtNHI2U9+aU+j+mpwOplyB8mtK4zQEWZe1iX26mBuKPznaz1fa2GiH
UWubmQzack3wU/pBFj7WLvF4e3YdNnGazsw4NvTTu5qc+Rkq3aLyQ+aJ2bEDdHP/
vCqUUJg4iY/JcAIu7Ca9UdEEsMrJLRd6LBxbjTTHZ8feLpmghmpYyu6b4tSlVFjI
Qgl5i32po85+MYPd56uyLIe1Gw/2vp7QNkB33Y1ycrBZXJ8XcQDi4vd5Zz6iT6B2
RY6f+WTXeUlIxkRMdQ+Ussap1qpzIG66kpd3XIBkO0juGcQBrSPRRBC5uHyP4p/+
9fjX3OZKz/yDHkFbZcGnGhS4bNhcPyZ1UZn/9aBxFutw1OLNbXdoPatF/lB/GDz3
N0ezQNARf00FrA3OTop+ZESPvwr1f+citYp0j6SgNa23LjN0cKkoCV0rWY+pD8j7
c6IGTTPdpBLYNUfATwr9BMqcnfoMGNuZgI6+rZAV63yw/VleQ09ZtXt9RTECiKvU
xuZKuE6bnItPZLrBJ/T3kbipTGn0oTIeA53F4PDoxyYHjABfsav0sd4HSt/QeRhZ
repGM0S2zNLtlqYoT5jVie7bMHgjR34umoC8F1/LkZclrqZ8nsJAKu2A9Ulxix+I
gVOgH9AdIn9W3rZlz1gDdqdXkZPe9WmZyyhV6je2eA9MXqakAWGOn+Mz+jF3lRF4
HmELfEjYifHrsbDlyET43BecXcPYh4qx07Q/1qPHHIlnHVudRL5ezqp8Yoap/24g
G9PjFQ7rPiTtzJxu6o4bSudGjS9ZcIhpz0gwoxZZGaPAvwj0bfr/YnpWv7C9EkF/
VPrSWgisWPhTBfRHONqZNvFaynMYHq8hZm6XDaTrSG0PPFSkaYfkYfmSm7O1fGtG
9njw62GEqohIKAyA2i54WV6QtABZmXwIqViPqPAdLhjpCOSNW+hRSaqLk1rH++9D
CVhdtJ1OG4Y+ZSnpiHcYf3CGH6ew+vy6G+3lE1lZWU5rttG3vjGDcTKjA2GbiGEy
EtzxNOpgtrva9eJ0CxQhfPuFJcH1hVsCtgakGTLXwVB6kh3TdnAmWLSn1XYZde46
Hi1w25Nmux2SP4yzW3rrQ6rch53kPEX0EUOjUdvO5xmy07uwrE/i146ymgkXR9jP
KCxwVV5UmhXO+0sqXeouuDs8pxNgJGabAcj0WpmhzEdi0QckEWKOGK4s813+dEr7
BtcHZAK+4AEkA06Ice/OpCeQee9wgKOwKuQpKtMuKSiIbQsn+RPWs9vCU0sm3Bhk
poMPyLXfYcipejI0paZeY+zce/ZL0eiJDX/bZxTa2t/5HQlibaL/vTTYekCFVXAF
AUKmr5ZmkJog65KRq0hIUjkcm6FCLxEXW/k2DNgW7J3v7tXU5hunGSgVPTe5ytxx
XI9Vblx6kfhdQpNBOgRVOy3vO78Dkj230IveVMTJ3GY7BzluCH2+1MPcZYpCqkQG
CWEqaXBobgfaTmfzj2VYQEIP2xtUrLTWbUChBzkJYiKiDDi6TchaXW28rgdKTKSh
FLvUehbotvhgTVZoDPQxidSecYjkjQQsTO97KOBUp2GqVhQf90Z4ZIemIVPPQLLK
+zMan574M8+7X/Hlgo0V4ZXCIbrJ/JJhvmmHomwFOnLewwMXZixWptOwZgO2ipzQ
SjtbVGSqDBGXInOsxzDwQmVOkxOTcWen2kUCcEiK5siBZfveKytWThnzw0ASmPb/
7IX9idmNc+mgeSNrT130U6LAlC/jw2A+DCZPrKjHRgL0zIu15c80XTbx8bG84pRK
VKVt+QmfS7OvmZ+NcX0UqCtOJPDh5EtJsFc9IL6qeS6gXw+xCw/G2Tv4xagWPiZR
GRfwLWeGiehvIQeS9zX2S8Wfq+lA6B0PdVymgCNC9dZ1ycB3YzOYd5bcMInLqDPc
dQJd2r3W+hwwZULPV0ZJik+AbwPFsTnKa7O/GLsqHOcsW5iU1mWQA7Bd3wOZsgE6
ZkazLU8oJLvSsf+Q8NAZjzLmEoKGqERk4FFiN7GitYc5KTz+ITaluxrOaAyOrSi7
b7RSlT7QSr78tA1lSHnxxEb2ruxmvI62hT/ziTX3xKfNNwaueu68El8vpQpWIrbn
k1bUuf6IyM7uLFOQk8saTJR3BTx2KQRzGgaLJgQuef8SjX8nDPyeeOvUr080o+PS
Bxk/cpTFuFOVCNulLdH2K7f4M2Qkc/QnxD4tC7hMaMxKaf7Me13Qz5SWvbLD9IHO
X9QdsWtqisLI2vnUfygdtqxTMwUEdmqa+gXb0CBmj8jcjt/wXXwfiHNnzk8rXxQP
H26fiWnNdq6i7aomQwJF00UB0XCUmZleQsoecPibFgl+LOs3jzdtR8xcWg0BQHwB
sVKqSFyouehse9L84uDl2ydD+aaOqCkP/GA4EPiB3aEatOU+hgeUXyM8Mbh57gnn
CWooYQZMoEG4nSwSbkmdmOq87P5Grw2bKRY8HIoyDVxSorYpsAPAeCpqpflmPu6O
izxdsMXgxAVpswYK96MDEUO1r8UDoZQmvVcJOhwKdqD+wDYysLdrMdU6FUtuWN4k
X06/KWP9loOQkD7aSvH/5qVDhlAcy+WFeu8iKvJnVr+sLoxxHDXnbVpg+FUAiaTQ
sF4yvyKILWJZ3WNGwLQ7AYbuFVkLomqp0AvXsuPO8VTI6cJEwek8l3G1LFTDVqDN
pSDeLjKlOBj1kDaf4s7qtA2FOOCuXQ2++ZuojGOESfwSZFAs/UBGXr/snWZSa2sA
zjpIqQRZTQP2Ejafo12AfYoZVcZ4ZTRWqBK9w4H4c2o+maveDO3XaKwUDFH24T8N
ILn4FkbUE1t+DItgNkh33aW7X3mOnrxZiv1DoBwcYBw+P34g3jLfbWoH4y6WLQNV
HCrRH3hnRN6/woFdonRg22I1yfKpfZGtumUW9UPrgCyFp9PIjDQlrkwkYil+r7D3
BnuOeNt3+ILp+Jc7r1i+LVWD4D1wSdJ6VAh40MrRoNuVuv21tFbCl93jmzrrprKp
Iqv83ORST6aKEU9G1CvTHV14yEuw2sm0p2KRzO2lNKoR51UYIe3HqAGgkxRbO5yq
B87SbVxsEZALSOFew6mNWWwAWbZLlz6QFunxz3V7wyXfDF4UNZbDJUn0hcEj22+D
w86dgWdan+nhiwNV76FHT/WlAntLLOuJcLD+yUGUZbd5nkwTuE2/uI0bZVTNB7mf
VWSYl2B+WWlushKR6N1A5AuHW1SYOhHnmJFPdSq11Wai1TkRtQ8l95EEGcCGRU0u
+VQP/wHAWagxeyFuvsEXYCTwV1GQOYozgQI4LJUhwcP+9uNmWCf4M1RfIF4D+Zpy
sG3GJjAwDCQ1yRnMR6JxnlAjkce+Cre9YHm84UkNMST1olwUh6YqSiVealyDzKjg
+S9KRVOT36n0WIf+EgaZql7Q1U9RuAGHeGL1WAXWZ+hkBy5SimU3I+tvXR0nRqx5
dvfx8NWWj7NAP5YU0R2zKRzdf+O1k+z8LT/AmvPjznEo5ujwbmvptYvnR2Jd+Yxs
dBfxGTrlltbelM/S1i607IPFHOFGau/yQ2yRFPTv9JTfH6dyrRHmx+EDaDwHSE6w
ZNuJPFWJTSbXXnFmVbWEJa49Yb0bX4dHH3F1OeueKbKo0zVXzF+LY33B8UfvYSmN
Q1WnW42p8N1tCbfxIOeCHCQS2R8ksD/JQyKqARNN6Yvf8sR6L1VuCa/OFCVn8ccp
m8cIqc7eiIw5MygKmjqg2D0tP64l0XGTJKZEyWSkOJ7QY+iK5UGroeD8ocsS3rk2
dQMlD/xws+Lco5T5KFx5uv13HMkIqIWzgrydP1sSlRCq3KmsYZD1fMkytYx1z6dj
l+8antHRsA0lclu9CJtHdzKrYRx4gHT5X06e2nT98HpKM9aHZNyIxxkTAup3pWax
PvnbEZMb67aapdF+BTPrRhgOo9GK7IzHchsCW+RnIv+6TK7uIYXq3q9AciK7+4K4
LMv9NjVEE9INbHMRdvVVeNz+hTrbWiyC01xzVODaTaDOn47ZGqQkhtc+xagP+SnA
0fZDLogFnyG3AodzZSTdZOWYiTUB5X03P/4JXLVREVWn7iRBCYiVj+8wZRZPh0A7
pw9w747j87VSUTBEIdY5pgWZlzZJP0U1mjPPLNkeMz9HtO46IwbYc4/mCvujcGXZ
ClNpmgYQceYdebAeJO+6sljGrNM2oLf+RZLECjAK3l2rCFLLaIW//oEp9/O5pqeC
s/t4yE7I/QFOplivd2CVc7sMcrX5cbGY3gW88DDLi/BfV9fW39N978ED4i4GJfQr
SylkzfYlmooPgEHSjR8YEpLxKHle+TZWW34CHA+bBGLZV2gTcnfTp4uDJMdiAJIm
tTUs6bSvVuHQcukM2Rwkw00i13Hv7P4ZMNytCdiXEKXMFXzDTh5sqi9JbP9B6Y9B
lXQAyDeWJB3YgB53KMn6ANo4QbjigbBt/Lf7aQDUVqlhVBH0H0XRtPVROwbMey5y
+KYG5zZIUySUNcZ7cCggHU1WIRQXjsjf6xR1DXyJN8zGrEuQ0GBnDJ5258nZUI3c
YAA03VE54xUeUs/ZlFYUSGMsvLYWyGGtD/H4IeoJZwzloTD2JyABqcrb04OXCfaf
omIMTvi/cvLtXL5RHwdKXC1ZzI1UdCZCGp4XnBlam2YXTCWcnvMDPcm+9ajqEzjs
9zwwVF8+wyj8tvUiPGXwKeIxh9IRJM869EiiXo0miCT8w2yMq4BNSVHXze0CxRx0
zvRGbG355g//bRfUwJrzQD9/shM1y0iD2gwE4Yzu4qmHMYHpp46ORGjcozBZGEwJ
pk9HMbs7ex46nWKLMivu1BCuBzAlZVkD/E1qXvUU8HVdMPE63gUHIppKHRL93Ls3
t4msrnSrHrsQGYtFj5XRq1MphSte92lrQKQ6nUqgyoIEHLdkeBnrvNSXqS260pXR
s3IWgkTFNSZ0MUZg3mPw3HfAQEGZ+LTI5QcNBOGZMWsUtnTkh/+CQVlvIGVQ2Nnz
oidB6NvnOk/3G6nZ+iIF96/9ca8QPZaLUFmRmyMyznFbIsYU8gHdZl40GEV5X/3d
gaNBXYk2wrJRqeis6xWvuW3SagSY7V7r7Zeq2m8FDnjAy26S2JjfZFzeYM43P9+9
ICyck+lBzyYAR8nkrosveboXEyws1IxMQn/1q4OAMP/61DEvLWSEvDot1GbIe7B7
lj66VzvAeRZHNjEbLEaBVbOR6xXB288Fznn6SbKo7P8zmQVJ0qq5kSu3orfNuvLu
7bpj/Q9nddDqqG6DEhp+GILp5pXCt7ct0Mug/28Nen81kdAbC6agtIhda89oQt0x
culx6aKy02Zf3lc6zqwtOk9YJWlgALHwS+dvFz4ALznucVZnNO5CCjVq7IupsRaZ
g93XrvS/J/YTjCaayuyuWPEssyMLYkEt5CxBZynVrrDfhqM2xDj0zvydaekTZaLI
uOG/L1Dtp9vHXf5HRgZU3irHHvWYM2omu9VIBJGYWx7OmLzw4HrDIdbcI1G8QkwU
934i+9KJGdCmMHxwYWvUOn5jplmugRE09Rk3KrM9Hdy8rA+7PMRR7W5eR1iuFsr1
C+THhXDBOsNwot314poqwGZhqPV/lQ9jICMFhtHEjQv3POAGr9G03J/3QDDd8rYJ
3P8dN1AhxDDdEHDk8FhDZ1EJPPDbD0jFIAD+2G/U02nSzr5egpwGr7rLsNzn+Uvo
eqk0nA4OMUpg9zh+8CA4MZOBj+z4y516Il1NKrEAy0dCmg8OBNl2VAtLJP9hdeOX
IJgNhyFN5s5zJCZRwle4xxpRrFwJXBQAInEPWBHdpari7JlpW8W9KE1PTj3ogmjQ
cnCRex/ZzF4RNgoLeae1y+6u5LlNycXD6vPZRQBAKpSkSwtmmahxDQ4vdo4UupI1
QUgy3xoejOEwtyhEdiyMXu8r2YKR1ajbOwHWIM1w28BE3bczbCcvStmogvHYnQtW
aKpx+GQZCUTLO+npAnlgdncM952k1k35c3dRu5b2gGuuYBMt8++qzxzMfB8vVTRg
aJVA1ri0BYCNTTNI+texm4f+99DzwngnBGRmj3e4TAQY4VhHMlxgUSD47dM597VZ
9GrituMpzZfriKE6u09DJhwfYkjfTsFw4NiQJCT0DWTQ2u8lQhQRhzz/3kWAEEHA
r7eP863I1qu139T+KJnwoDWub6xzCZvccLoa3fEP3wkvXDsWyygiTcvleRc7mvI4
EEXj7123BR8+lqDTOAclCtnmrN6n0fJS3LS/PXpb1YVADtU+t5aaAFKSFj5ajjPv
ldeA/DR+shMZcOQR7SMgPMQdxOlR2OtTzabewz154xBQaDqii3qeYsuUMY4SY1MK
CfQpTfXSyQm6NHU9fq2fY48DBHk2FnixWV4p+XkIuOdUZfs4gcXfxskUq5M6Wzt4
4qwuAq+egRViAxl6JAuiNncYshNNI0jgtqlpyq5tOewXTPYwTwJKapkMWcAknt0U
QmF7+awZicObqP7Uq6e6ZDxXSbzm9yAt1eU97wmwlZvaboxoptPZrOWc5N900xr1
NZ64yeUqIXCRU8AQpS+HIyrJj2G8l+UbZYJp0Ov3J6T6TesY9SMInCGTYCaXZPua
sbGUwBch+U+jQ1ls3sJd++d5namoGOnHqvCwhLJzUH3pBhHcsWPcjoZ94/Y0bpSX
NXNtXzjzZMWIzOpho+lpw3t6gijB+hUquV38V9lxV5IrtBcP1MPFRR6FYd6hue8T
IrIPFi48LLjf9SoMTAOFtgf8w9TQqAq/PT5l924ohHJreAKzjvHIw7ScH3gMfmPN
T+JndlvgtaasWKexWd2xvjL8Ef55PG3q9nmZ4sJb+knQubWF4QYsfm+J6r3zrKS7
ucG3pSLq61OToTj5xOvHOvthnJAwJW+8wU+F+FAP61RPJ7saDS0abY9X6HHGTRKF
+9Tov+cwfUtOn5fnyxRwEKaVzB/PcYbq5y42Q0V+YN54bRK9n7UXMch7yCUZMvM8
PZTo63yvw7VZBp1QJGz50LJ5J0q9vlLneQ7SAfu+yWTrjOH5oR7lcVYEBMKo4fQE
ph8VIJqQ9z0iChrNHKFIQb9pzwLth1e/6dfZ+NHUKoaqq8d0ors+XtVLSZRrmM8h
FffeDUqAg4qEikSI6Zwf5Ip/AXxBnQotUosQ4ljGmLy7icnwP0thbSK7YjDK/Ihj
LmgIqQ08ttJ9m4ceF8GdZiYPDdZ7cBBj2arWvqgVTNjELprlErg7VXYa1wiVnuMo
+dekO2j7PXtV1gMhfO0xWx0Cq0/6ZzTH8crzqAkRravqoMNOvzV6KfXJDOLXrWlq
LgZtLSbkxoUyqtRd2ETG5ZD5sgKxw3uVXGoUOXGdgrp1pgs4/aANxf/ROQl/uhxW
PjUfTAy/l+V4ZUqk6o/f27in19S09Lxuk3r9S3HLBHImLbHt2O2EVLRL81qTpiM1
AAxPdXc8m1t3c+IWRNhcJloD1MbPVRRb/yH1WKxqS4F25mbWbGcor5ij7JgCgOmv
v06tS5VHJt77v4CcHF4Qt4EoN6r229NgkuE659EE5EyYT49goh68WiiQH38Bx77o
XU2QG4NGUmjPnTLLgCtcnZvDX/XEJ3fOjTpfCaGPtaNkKf8/mm/MwyO1NOhmXIez
CHXwbuEd3RBgwCXzuGSGDQRg6lU7Z8WTmKa2WfJhQae2dUbzSLl8dp1NdxW8Hlc7
z9NtRggu6uPGSojQFhfzC8CME3LHt44cAZRIMt1UIskHx8WEJ2PNjZhVC8VOKz11
qGUzujach6LbHd8mgTv+QRQ+LiPCCc3muK6vq1gRM7rH6QWQE56HiI7m9ZBhJh7u
nbt5kYZPIiNeEFXxWoC0obXPxpZKGQDA8T0/jNdmnsThIm9xOlT7IcMjtklJgc9t
JKUhdNhANfYaL+P3YacFDHKCr308aulSkIriIKw5iUD2P8Sfdv1E+nAQNMp3M9e2
XYPk7is6KCHSLB9bNyZc1ysNsGwvCj0gbXU2BkDfWYinj9XFIsAogGFvTxyoK842
ggqs0x568b9jBLj/6x6JP5Zve/FGR80BddxPxq+X4JXemJD0FkJ/7Tv1B9zVHyBI
/Oc7sbFMdg9sWc22BNkFrs5VS7L2UT5+R42sYGLNna7aq5HpzXkp0CBqo0nf0IIa
S5v/nmIFb054ZrtM4ktpC9Cv/VHMDTncRTqnLy+/yfQPSSuXFZ6w3K3vHLDxwm40
6HG9ndBjBz7k9kTToJyr5hgZ4Avi+BYHd19cG7TPUvzgz11ePqfZb3RhTbsoeYQn
H6Vp95mc9fpeID1JN9xtJPYFdhPb7zwJfK+fxcCwo0DvWCnzk7ntD4iSi9JZ9yad
DvJ/TFowETC6j8rntWQ0dePS95VMz9PtVt5DJ+VmsoWBaKIg+ve4zPI9bjORlABW
mUYpxjG9MbCLCj3dezwhvGidrdOTyOEBaIf/aC1bG7t18dT1h3pBY1uU3vyEM5A4
4Nd//esFoJ3X+l2CBrk4kQ6UwYORTugmp+FinQC6nB2a4NAwTchUhHr56XDjsYkd
DsjFdCPABSAtPC0/NQAlVdWnqnBnRraKAl7SMPtcVMbiRvLkLarPWcVrcF+DXv+N
AYzX1r9CygH3Ei1QF+Rqq1DpODBGgW1Ueq8LUfYbIOoza4ml65mTF8fnNTRZ9W3W
I4g9UNAPiFfSY71iNoSEK4m6KUPU/eBuLx9XEc3L+kGI0+eNxxtTaw3fIO73bvKl
Ud1A6CA94zBWMLG3skUKbihG045s+OoTayEFgp5Il03Lqe0tkVOmH4Nw2QapH/1q
FkTo/CCOo+sEU0xxOH5/SWaJcI9cgNtI6xvUt2XU8DrRTKw/w1B9imSotmzTdp5Q
IBss+bwfbo0Bdo0RwD+ar3LNVrFurEifZWbXuQj9WEbLpCl2IJX4F1xd/ruJE7uw
`pragma protect end_protected
