��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�Xp!�KH�_���p�VF
B�5ߺ�0�!Q��.�61=���TB�ڈ=�GSѥF<!�%(�j�K7S�V����%�N�~I.���Q��騗&�@B�z��g��7BKm�.΂�GO�~J?9F��x��+��
��K���$����p��+��Щ)1y�3Fk��X�=&�h󔱺5�|	��a���e�ƻ��tY�u�;w�Xt�n|NU��F�fe��'�<��d�$�1aKռ��Ď���i��z�|�z��6H��qۅC^�:�+�697�h
�ݘPӬ�<������Fo�mT��/��	=��̀���lTK>���׺��"%	��;w��~%�+X�{����c�3t�l7َB*��Rnf:��L�������)�I9u�N��sc��\��G� b�7�C�Vt��r?.����LvX*`,�G�W�|�k0�&S���v����^n�O�lx?������]�M{�6#Z�0.�3�J���a*�w�^�-A-5�[i/H2�cB��.,�cb)t��6�F�x%��ĶN��ѷ׺�Qv),�ۋq�N,q�кe�F"b�܃�J