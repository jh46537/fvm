��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�	�O���T�7~j�K�e�rd�nWWg�kKs�<X�@�U/�T�d�=|D�7	�Z�;�[��l�Y�F��G�}fG��R��v�e	Kg���>���[�r����)����?*�W�J%7	��yl����V��%�]��[v�#�xxhy#��6�􄤵O+�Q���;o�w<���@9�c�n�c�>/�hi�qv>��}Y�0o~���Y)�M�������TToxM!H8���2b+��ڞ��)J���DPb�N4ͩA�]�����ZvPQ �b��Q�;�Xd�t���1�7 +�i&�y���G�4(�f6�:���y�-=������h��o���@�䨽����WBo��3B
�7�g�Bs��$y�Y0ߍ ������y�V.�� ��[<�{�9!S3}{��C��QU��v��}ʹ~B�k9���lϭ���'�+^H�	}�{Ǐ%�ĺD?���-�������s7�3L����j4����[!����h�1"���|6�Ȉ�̘1鉖kڳ�e&Ӄ�I��p�t]���SQL�R�7T���,tm�'(��_�`�[�X.^��)N������"y�L��89�P��1��Yt�t���0����gq�b�Q���f��XCl0h�](�((\�t� �뛘R;9Lc�Wƕ��d���(��N`��c
H�.Uh��:d�h��̀T����P���j�Hاr�u��o�-�Č҇L��߆C�d=h
85��OY�Ώ�-U|�	T5��E
�rE��,��{�]�7zEeȎ�\���>�9�͂�+NF.D�NK��+��N�c&?�����\���k��s1���5�݁��/1��^F|7�j�Z_J��v��\uA�w�Σ���:��8kз)��2�z�s�ǉ��A������X�*��"Y"�z?&� ��#v�\/�x��;oy��E\�r��8���~V�&Z��K&Ϲ|���+�1](|� �&�;�r[3SF�AM���坿�
p"'T��/CR��d�a���,�S��m{tP�N����M%��,b��0\$�3y]gd�d-v�;���@E�@�8�cޒ6�z�jj47�� �H���|�m���hŠ�k��a�LFWk�ˠ�)�O�
�k�i\�6�!`w㋤��Z�֙�I�(!D�x�mc-Wv_�0��EsE�.�L�U��m���̻����l�uM�[�3�+���V*��,��8�L�/q��{�;����wi��DX݃�g�=wwL����V����n�7�Y��h?KkB�A�y��o7C?����R��SS;�E9g�hH$�{U�2�L�R ���;��{L@D�S�ː�ޠo���b}Q�E�k9��y�_I(O$��/��7;I�����";��9�ʲt�foIr2�Z�#H2mI��^�A1$��K:�����m�F/s�=ʤ�ՓL��o�ze.�ƴԶ�'%���l��M�j�h��Ȓ2J�>�H^z��=��)�	Cdq��x���#M��p�ivn�@�5��}��OĜ%�	fF�1�r�K�j*'0��*�^��kHpX�����k�K@�o�g���U\�tTFp3E����`B�d����i���	���3�)H��KsI�^��G#�V�����Nml�� h\ꜧ��I�p)t�@�2/��:� [�����Y��鮨+�-[�KKF,������e�.�49��K�Ϭ��[���w	|G�]Z���D�o�� �U�e��fv_T��]�QV`����{gF��/��+K���u	t�v�./�-��u�
�~�<v�R�(z�k�%�B��V��/�+��
����V,�.?(δ�N<�����K�#��a��Q��ڵ�ѥ����o6C�y��k�v���(�+�v����`!Ք��c��m369>t�? �[j���
���]�)(�j�~X<g�yk�JL��������.�d%�,ѳ)8;f���2A�j�PO�9[,U4v�7�{�M���Z<���O�Z��)X>�x���I�z���g�ڣ�	˔V�8f��9�U���a��ϕ�IL�l����p�SE{
�k��{��V�� ���G�|����,|PyU�\Xխ�C�w�m�8E,{�д�?5��*v�)<��5Xqw��Y|�6�
��<#�5�B[*&Q���~)>��(�Cu��H>��(VS5|0�%�,�4�qP�GN�FBV$8�D8�Vf<~�����L�4ȩ��g� ��E�zsǏM9���Q4��sk���ș͸#Y��B R���}
ݓrl���,�V���E-��}a��u��y��¿�9_�Y�C2�X/)����=��NN\^��h t��դ,��I��'f��aЪ�>�=g�Gn��(x>��(�(�g+�1��M�vp��t���P?��]=�Ԉ��1��Ǳ�e�/��2/�S}'�t�)0a�Zh�(����{��9�x�(��r�����fT���'j5u��QUN2�9HQ���3wJ�	|����&���~�U��)��2�t(�7���k�!�4?����PV] �.�tb���ޙ������������F�'2��,6�O�ryBK�o��y�������6��/"7}) k��^%}��N���M���S���51��lX�������2�$�#��r`}���L���ⴵ�e�mL�D�IBm�G�`����q6#��re랕u@�P2�ï�>���tBl7�
����mK|nh�1u�<ݵr�<7�Y�Ref3��+�'CI��������9�^��<x;�7 �ԧKa!9��^OJ���+�4T����S���Рc��O x5[(9��6�r��^Z����E��H��}��Ҽ$���4�U�Z�eK}_޽�a���WuK�oDs�v�k�����
6�� ,b����Ed}�W�
��"��Y.[��W�lXH�ITN��f衍��*1&u��A�RK�V2t��Cnx�.#�):�׻s`ܛuei@R\�B)�a���(E�-����jx�8����34�|R�������f�x�oM�YS)Y�k
I�[_d�b���`!�����r��&�$ӗ�_Kg �����������{|��E�`���C�f�Ssj��oO��2����<�
��r������B;*>��ˑ�H�I	cV�&��)�Z}��%{Vߝ�5�ɡ�^;^���##J0�<U�,����D��"��)0D]q�e����2��R�v{~�X��$]7�#�_,�R��y�7��1��;�����pW^��$X�e��\B��l,8;4����~�^@K���X_36�V|{P��4����?��r�M���n�:�\!Sm Xʆ���<�4�/�������򼱇��o��UkT�����O����)#̟-|R㣇PCF�f���R�M����c�˼��H�_HJ��B�A)�O��9��Eo:�b{��ԢSD:�&�ɱչ��8
34��hN^�5�{��v��p���$�5��5Y��d�1�a���Ni��0Q����d�
R��?��E%��b����
21*��p�)e2�B�s �A��1���F�<��,a�Z&
�X��p��wE�Vs	
��H����&|^�v�L�p_䄏��ME�Z19�E�62�F�J�p��؛�g��Kܽ=p�T�-��'�
]>n_�M$J�J8-�U�ԕ��ր7{-�k˦���EשE��*���a��=���s#��[p����F�b�J�h�ڝR�0�jې��`�h�7��Tt�
y���K��\�O�}>U�E�ց~�1�Ǫ�U��sLe�£k#}yT3�P;�M��4Z<jd�J�q"R��ZP`��7ҍg�����`�OZk����w�gb3Yne%.�π^D�ڜ��ݕ]�ڏ5��i��q��e���2D�݂�v��ѭ����%����1�=V�"�4/C@ljfC��G��o�Ԯ�9���r��%fT@j��	�9+��\_��h�@�݀�7z��>Ī6P�Zw���l|�,�ˣdÈ�͉���Z���Ԑ$?�7�~���0	ݱS�֞�Ż9ϛ�q��8	��tGg�l��t-���nk�0-v�z��I=��d9!]�i�KO7	�"b��Q�˼fZ�����m��'0�?�:�~��nͯv��Cە����@�~�� +�Io��|�Zg,0]�l�i�TikOo��N\��c�ES��'�����{�K�wJ�r�D�������t�����Z���?P�#���e���'tx�Ǫ'o��{�7��2C9�j<�^�H��3���p��l2
����4,��mmt�	U�j(:dao�|�n5�1��].�C:���V�3\f��V7���	0��W5�g,��y�fiu��� ��]�����Kި�z����ҋ��Pa��_#]y�6��\R�<)1�0�a7��H�m�E�y�lӧd�d�Տ+VۏmS�M��H�?J�#|Ppu!�Pt3�z�Ck�L���!�{�u
)��5��aE������%�2ɠ�*�=�
���O7?A��7<�)�
KB���{�#	y��YΎ#zJ�!�G�sݔ��Q�[�ax�1Ղ��}�褅~%)���GU��XSw��$
Jy?.�$�%����n���Y�� P/yc܃PlEw��C`y�q��$k=��h�4����lK�99����U�gz��M~�W%T��P�.& �/�p���	�|$�$*��<[��z�.~RĴ� B�׀��,��:�W����̴�*!�_kFj��ƙ�io-k������2�P%3�� ��/4VRQ���0sZ m$�-.�q�1�$�#`��e��T�m�gۿ�}eۧ�,,�D�^�Dz������H(ʉ�94 ��aGo{ߑ��/��Q�GX�����NF��%
�uf��a;�cX]�����Q�X�VE-V�6U�2��"0WV��0Q]����3R;/��f�)oѽ�MO��+��X!����,k��u��C�����4��Uo�'�"8�zAF  ��PG9�?æ�j=�%�J�"j�h_kHѸ�Y��_z(U�w��g��bΟ��6*tB_�	B����w�H7�aEf"&�-�hf~T("��:��xe