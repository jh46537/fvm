��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb� >��6\�4-�J"I#wL?2o��e��f�p1�b����QW�����{��E��/z��3��m{"^q��:�r�<X�z�@,&��F$��e?ƫ����kV���%Jڌ�
����b�P����gq<�%�rP��aSs;ee�G�+����Y�i5���y���#�W��U��0�]w��{�6JC�LϪ��y�)���n<�X�����E�m8Q�'���o�t����BT���A��)d�����{��a�$ז !�����X);�".�)��ϟ����rA5�~u-,wDq�h��i����on��_�_�PPk:z���
|߅�{k!Jƒ]����k��Fg�������N�p��U��tsxSI�9�xm6z�{�U>�jm��y����4q�q�v6��؆�A��xB�����A!�e�w�8�2n�E ��Hq�.ж7kH+�L^PC]��X�����h�����h��op'�vO�>f	�Ͷ��<���AЖ<�`y�=�c�aL�{�	�z���6�X�-kR�Xc�����b7��a{����ʒ+���0i����Dy�T�=hT��;gH��c\ 8��F�nn�M��bc��ķ�C����fZ� 1n΄b��������I��g��8c�L�h)ov(��	9��@�iX����߲������5@�K�<r�7�L�A#H�^�ܡ]�fC����}�@�܎嶊ҷ�e���?�#,����tX
U��|�%�?��u[��m%��uĹFtĪ�tӕ�R����!Z�����E�
(��)w�2�E���y��X���Ͳ8�y (.��-[�p��z/��	��Qᕜ|J��W�r��p�O��o�[W����(��U���@vH��e�C�{�� Q�`�,�8���s!8������m8��ع��N�9lX:�Ԩ=�q�$�M��[�W�����x������ޜ*a˲<{�Y�j ����� �,*Xئ�E��+�=�JW�8/�ǖT����L7�7�3�:�MQ2�8Vw��z��|��+�e��#�+��	�d��Ҭ��ϰ�c��?��︭�1֌�
���DƟ)`F+�&�=�p���fCn��P���ʃݨ�7C������݃�����"Z-}6iŕ�������~��DW����:����0�g����[)�W�=1�<oˌg�)��%���8�tڿ���M�/�C����Z ����D:�M���I�b:���J:?g��G
[=�w;�"{���Sx�Cj��UQ��AR
�΅�9v�K��M�S� *rY`G,M�ǅG�y�m"��p¡�|�� \>�7w��ft�&Gf�JW@���b��e1���H@� t���*n=����G�}���0ds�w��~g�B��"�S����W�`s�Xt�a{�5�A�G[#����	�׵�����g8�4k�HK8�ʡ��R�7b�ڊ�B��~��f+�3�<CJ��RA��9��
�+��U�`�TE�,�c�1t�[>�8h�����Gr	Ae�\�M�rT�Yyv�Ǜ��� ������&t}��Tʜ��$��e��Paat�ޙ3D/φV%J���/h�����Q��^��ۂ
��Z�s�
%m�5��,�3"iI���H����h���_{���w�޲+A.�0U��\q��&7�!:4����̛�հ�tH�d&YH��A�߭�`�>����V�@�c�h@�#����Z�uG��ҵ�&�D��R�'�E0:	����"h���Y��4�N�yZ�q#΁D�b��GѾ/�^��S�nw"�.�a�����,�=ْ�W9c��	�P��@`��_��:��v3 �>v��#	C,2�K&FT(�`,C����k���P���-�x$7�=����Mq'�čJ�gmӗ���_��2\��X�X��D��z^2K�;�x S�!�oS#������6���-���s�d4Ճw�gxP��d�#����M}n�?��@����9��6�%\��5�E�X�x�	S͈�X�y*� �ix8�*Z�Jޡn��u무p�~��WR(�A)��f>w���SQf�5�i
-'d���(�!~��W���|>X�gX��P?�i��NLۂ�)����~@��~@��G&h�S�l��{N\y����$�"Ie�4ŉ�e�P)�-��Y��K%}^mb�T��_�� 8����U�A��I�0�l��6Oq#�c Or
g��[��+
lh�͞����;Լ8�U:f\���8�Qg@.&���;�� �S,a|ʒ�������{)�Qd�4P��8���1f`���/�wע��\j�����f
>4�#��Ue�(�E��()5���+�"�/re�1�	V<ܩ��tu�^��+|�c�������f�:~�Z�0�sn!�^�J!f���ݶ��<�U�T0��D.��C��_.���lbF��P[\H�R:�~��a�RzTF�����а!LP4F�ش�n;P^PR� �%ŋ�m���x������9��N ��T#^REA�8�$,�n�9�jj�9ۓ�	-L�ҿ?���'��e��9R�X�xܱ�ò�O��6gGE[�B�Ҡ�mCYd�+璐��R�����U�8Ę|X��q��o����s��ߨe��B�Y^3����*��* P�},�t��h4f#ܛ�lï&5��Q3�t��9������Yץ�)!�X�$�����"�w��4��x�fn�a�a5�%����;�o3xu�a�/���)ں�3����Vk�z �S�%m|V+�Q3�p4vD;ۏ�L�Q����%قE�`$zЫK���K�9���I�;�"5{��s��!�������
w��v5i�N��c��ss�%)�M�r��(��ߥ������F-��p&�J�y35� b�Mt9sE�[�/px~<���C?��m�eྎ~�9zaW-؅���1�0'�o�խ�;s TI�ReK�Y��uGE�R�YM� ��44�-G�>2�9��K��Xw�����q��p�	�m����mA}�����MP�~=(��"-5C\:�;�nߤ���t�Liyz�b����Ό�i��2��=�B�XsطL{;0a�����m�7�(��W�򇩈x�{|����XJ�OV�r�I#����Ϗ��nsi�|��܃z�5{�eN/�d|�(�����Vt����!���QCܭ�% zU�����g,ȥ��nŅ���@ۺ�$�k�'v�a����;��M�'�
�����F��U��L9b��6��.��[3>�~�]J��=�H*v|rn�C�r ���W���#�?�Uk�'�w�yV�+�W�����]f��f�/��Mm�-g?�@�Ëc��5�;&1`_�,m�y����������o&��1�	t6�I���˯�<n'�s�S����Ja�PUH��݀�P�c����K� ������l�?�� O�S��4_�vȪ߮I�
��ҷ��@��B��3-[^%�禘�k��"k����V�:/W�\��@[��9��b"�h�>7-Ph��h!�*�-Q/&Q1؝#�(��^��T������mz����ߑL��D.�@0L�y�y�0k�i�>`~�!��ŭw��Ga|��6��7={�W��O���^g���8\��rK\�bq�����/%�W��s�P��^t�:����ά�nzz����$Φ�����k�M�<�-����l6{�������F�'xV�
<��t��.����`��!�(�)	�7��Cò�3�)IUU�&׻��sD}�Gz�*,�V�8��X��	�3[������/��PN=�Cp;�eT�]v�"�6GFdGuO��`��`olF?����A�]6{�DB|�|�\�+�b��ƾ�i��1P��kc t��nGpZ�%cl4�ʘF�zw�ʜϰ���)�G7���+�{siX�p���[QbϹ�A\8Gk:��b��3䙇����TF�a���s㋻\�9��ɶ1��D?e��YUǍ���T�kL.8�����p<����ę-���{�n���c�"��%Yǳ*|0�&�*Тдx1�����\����c~���N�r���']#�$Ĳ��I�y�G:wr��G�g�9���JZ�9��Q�o5t	&� �uvs��#�E-.�@G���Y
�7�p��?��'��>��S����8��p�2_���G�2cO)��j�]@!�*7[hgO�on�i�HF���ü}&�X���.�nߤ2C�|�jDI�̫��a*0@��5�:�P���h�s(�w?��L��D��33IB�,i��w�߿�Z�#�r��7���B�Ԓ��-����a�d��قKr��-�Ic5~ 7���Ƌ�� k�H�ca���º��� �Ȧ��e�C!�:\�k'�yqt���F��nH���f�5���|�g�ߣt�Ш⋼𜦉j�Gӂp��?,E>��;��̇z�
G��x擩6+Z/9�6�NS�i�负�7������0�>�w
��a�Ñ�%��ǜU�g9#���&��b�z6f'L7��
5ۏ�2b��OkQ��G)�I��G�X �D�aJ�H�P�9Q�p'�ɑf�d�N��I���g���\��x�г|�C2juBM�Vl�ע�%�M�`?}C�x�(���h���\�#�#���W�O�Yl.����}?]8���]�lzD�`9�%O�2��k@� �͜'d��!�.d�cC!g���2�<5�;JH�o}���<I����C������i��F��u���n�e��	-��a��D8쭝$-�xe"~G�?�sl�跾d&0��U�]����Fr��k�8#\YL�YHW��r�p�1�S��Y�kl�B�b���`�� (�g����G���Aw���ӣ�6�y�b���gV.�^1$������cÉn{.�1y��JZyn��C&�&�R(۾�������I�^	�����j����'��*�Ђ4ڳĵΛd]��5C�v������������{Ʀ>�P3Ѿ��ƬU��� �T��@8P�R"�����[+fիr,n�}���~��ئ�9T��^����B��;�yEH�Ŭ��n�]W�j%�I8����,�v����졙�vӾ
�g,��ؑ���?M�K�v��y�> M�-0�G�}��Ƌ�������Ж���Ʀ����ii{Wj$���r(�^OÆT1�V��L�\��"&7��ʶD5���x��4��b�n��0]a`��-~��ͧ��HS#�+�����wwO�Dȅ;����?-_�ȶjxr���� =�9����L:��B�j���E���iu����:�N(���IB��g���CŤ�jC�~��l�� V#��dgV�H�'��x��e�$��9�[�HՋ�����6l"�&*��jx4�A�&!�4�&Sx�K���Ls"�V�'����BAjf���+��L3����ȶ�ؒ��fV{����T�~�]sOg���A ���=P��t�c�o/����7��܈�X�5��;�X�$:��IO>@G��N��D[�T���
c��*z�5��
�+�&�)e�S��)t�Ӳ�r�BT�����mr�cŘ��ar{���\ٌG�猀��l*�&�u�$���F�G��5rw��jvgٛ�K�_d!.��#'�9��)jD�Z��T��¸��0�5�A�m�kG ���K��">���$��P�͛f��}�� ��Ԣ_=�'�ia�=#�ʎM}f���M"m֭θ}� R�|�yC�A�9+��� �n[6�%I�r���)X�jK�V9v�2^̓�S
<�\�-�o×#�_�Zˑ���j�
u�ˍJЯ�E��5~�b8���o�\<�a�ԯ��*U����{�.gq?�6g���-^x�������s!Y\ R#��Hehj��:�(�n��bQ��ha2�M�~VQ��?0�4�Q��|�f8��	}�Γ�ǘ<��Q�/����6�%C?z/�?��a�Y"�`9n $�jz�d"s�7!�ҸY)����Mb���Jh*��4���
"�(�4���	W��n������Ea%$�+s�te��f�I�eir��j��I�O{� ��"�����>�@�&���%ٕ�6��z�SJ)�Ri��.��^�o�58_ub���8���+̓�C|�k�Yi��S8$}��u�Wd
�K̏���J�~������c�b�0D����XC�q�(���#�컁mf��$�|O�W�?X�5�(u��Q?�\�~����x������؛�ĕ���;R��Ա�.���$����C�]����b����R�E C-�H�@��Hsm z/C~A]c�a_|L][e��kv����A�m�A%��5����T@A�J��qu���sqY��0}l�M�{���y��������}�|Fȅ>N�����i'gQj�|C%~�6�E���Р7'�<�a�� mN��l��v���Ѕ��ho�t.kG!�̶fnnS��-� �d�eU�B��)�3{�#�R`�dv��^x��8�#�~- ��g�NvZ�,���{oXߝbz���(�Άs��# ]?�r���>�L� �4=ŋ=O�c�7��JV�{U� �<6d��@P�V�>>�����r3��7�PX-
�?����Lb}�Y<�Th�jML�b�~�����G÷�h{T�l�6Z]\,�N�a���!�c��8jO0���w|S�|Dw��A��R2�֋�i��b�(����n �!}bdW7v��)�7�z"����w�D�ժ���G2�c*ck-��e*��m���F�5�Ւ��>R_ ��}�n.)������l ���|�US6�ʄ�|ݤ{"��>c��U��w��u�^��	�RW�J:R�D��<����72C�%�6`�%��D饪���AQ�rb_ӗ���'�tK��2�Th�f�����K����l��'�ԣ�����s�cl]��[�_JȆ�`�,J�B�U͑Ǌ���.4��Q}����*��3f��N���΅_���m"`��ӹ�R����L�XsA�Bd����+��p ����&�a�ƺ���3~��U꣖n�[���h������^ �&�eLb';xq1�?M5U�P�k[5p�>]�_���N)R�se�Q7g�@��d�~�s_m^qppb<k26�2��$�,���u�W�{a������9��y�U��nc{ؼ��\�R��}hpG�/L������r?�|�c{O���(��B	�wx��F����/=jπ�ZK�V�ʊ�S����d�4�Z�[��ZQ��8&�����#���P���։�Y�+_^m��ߗȟE���~��N3T���uj�V�?���`:}h	�F	MO���6Sj�WƙiL/1zw��ܥ�9�\�za��wI�<TN'����.�W �����>.6G��,��g3�(����U�r�Li����B�������M8k����"��Ѕ:���U��������G�ʖ���H�ut8z����<���cm�4M�}-|�u�<�HwFN�ּ+�٥��Rms�Є\.�F��7u��c(]�����D}fx���Z�|D����B,_`#ʄ@�r��2�4�~�;pK�vu���V��c솊�m�̎���fJ�2M6��lGZ���$���D\�GuV|�Qbtg;�Z��X~P~��F�R��2Z��n)MW���Ű������ffZ��~�>��,��[2�ELr����%b|�}��ܝe�Ϻ3szM9�$� 𒈦;�%CF �B^�%VY�U����>�傟���J0�1e}v��y�JҺ2>�M���$9�B��E��e���� �8MP<Y��"=ZlE�B�u�,������E1Ga�i'Y�k�'�[��&���b���`u�H�n�Y�W�p�Vɑ��z����3����2
�s�,8"��~��G@���q!?��U����?\؊�}/T~���Wh��[?0-L�⯢��x��
�n��ZDlt��\�+`Ǳ��s�7m�8*����E�<_|mmS��h[�"G�N�xk\�On4Jj�l�R�:|)R�3�$�j���*b��<�+k|V�T�-�\���~q`�5���ܱNcRl�ss��d�Gw�K�z�0dt�9:�6�eP:�B���V$�Ŋ�̱U����z1��<Tp��r�! �ҵn/�.9]�]�w`��5͖lV�9�'CY�?]��q;��9���$~.�ӥ$-��k��/6����Ђ�%:�v\�y�"�񰬠$"�Qv��-l���/|���<�a��\+c1?aw�2����hu=��Ra$�!+̂�~Y@j�[�<�#I�����.�e�ɼ��� �<�%��q��W�nB�KU#��	�f�&\���=�9�/����c}�p�`U�'��n*�(ҫ��8�?���DrA?�݃����~��Cm��l�4:�Ͻq�B�K��"r�C��1Y73�����iEޫ8��n�*�f�3���kPq�� ������Ot�sU����as�J�H�q�M	b�Q�G'�r���3!	�8�����. ?R��Qˀ�9�ĝ_+�x�d�Η��јLP��~�*������O��v�����#&��R�Z<㏶��8��M�|��mWe��!�Kt�����]�cr?���e9~�Fo7}��px/�~i1��b�[xb�}���W%�<��J�Kz�wT�Z�y�<:�T�Y9!� ��T�/��Ҡ�C�Ȣ�����\1�F�b�o';Za�p� KǸ5oW����C�>�מ�؋HD�����yx?׀)D��-�K�����ȹ���8�TX�v�:z��C�}���>�̕cI��z�&���bj���Z_1������{�#�t���cb�?��^;{�7���p�fX@f��Cң�!y.��	�x���)- }��`E{:�;�T��N�kX@�P�k���R����y�::"��� ��_~�(�o>��o5�{*�)��k��߯L��y�����ԥw�w�[�mD)�FV�=��:x�g2�`���.���y��M���%.��j���l��C����CWLU������۩kziz˂�u���ڱ�rR���DB�/���#oofb��~�D��DmW�L2�˰�[�4�¤՘_nQK��Q�-� �>,a�����<�%��ߜgE��~������N_O�U=�n��ˤ+)���G�s��dV�&DE�~����۷���4�M�CU�Z�q@���ը���.����xo�=���)փ8�P̸�����Al�P�yJP���fݗx��$��<1�拘ia	Į����''b���������{����($�<�t �˷J �f���LN�yj��p�-w'�ZWa��~L${� v������n\&��n73���W�s��{�!����ul���e��5;�E���zf�+��K/�FKI�c�'<�Z)�Ru�[KL��j��wnv��9#�o��۹mF�5�̼b�~���$n��%��!��h5��b����5�
3��?,����auq�9I������q�l�EVK��>7}d�'�l���d(���Rh���Mo��;ގ����$ �L��"���0N.b�}G܋���t�k�ݹ���ws��ڻ�����0m�������Ҩᩔ�K�
�=��~Q��LQ�ޚ��Փ��:���]�<�)�k����tP�Z��T��I�&�E\oF�),�D2���������x��^���Yu�1f1�e�~���9��*#F��eZⱻI	���)�{ݮ�r
1|Ꮹ�hF4�9 Z2T+EkR~��+��B�۔�ܥi4+'���y�e� b�R˷�Y�*��Ep�,�}��,|�TWq�y�^���2!��f����E�J$�~G�Y���h��vz
?H0q���gU%t�,iz<�oZ�A�P-·M�{h�&�iY^D�{�k<���⿱eg�s��W��5�I>?�qz� �2rEb
JrR�X'��A�o&`{�F��7���E:>�3X���/����.�<@��3�M1v)�7�?#+SK�l#r\��~�ֿ��I�I�����cF�-��'tt ,-ZW>��sη�^ʤ�a2e��t8��������P��+}ݢjh�2%~��T�#/Λ�s(O�y3������d�Yo�h%�JR��B�L�I>����x:��\o���/��ݪ���ʶ�8����d?���NV�Hg)�+�ycu�홗[�~�䆔�T��+6y��Ŀ�5���]g���^��0`�g�ȊnU�%20��K��bwi8a�XC�Q;L?GѼ��҅ď�ۉJ�'��J�qW����?dq�*U�q.w�z��{�t �M��.f2	�U�MT����~�N
l��
'��=��v[���)�f+a��U�p�R���a�}����\�I�y/���um��fӰ;;������9@�(�L�>~H�\���m�70
�x��n�v�SjI�g>Eu�+mJ���XN���k~��?�*�l�*�|��2m�y�d�w�SM!,>��3�"���F�i�25c+����
���M�9�u��죬UM��>��R���%F�؆Iu����xe]u��	����p�5a�� /�d��r��4D�2/!�,W'���e�eɾg�r_G�LI��0tR^�`@�:h��{�L�yØG,*6�/���ގY>���k咭\f��0���Y�ՌV5�dh���v�ػ͒#��i�XL�ծ z�,�}o��V4��������1W�ίC���-��>�Ə��;ئ�1��I&۟ �� ����S����� �����;�&/���նTհ�_��%����zO �p�вg�$l���������'C�.����'���幜
\�Z�m��>��#}�@�u;�(�M�N�<0��5�}XM'P㇉��f�`�	e�4l  ��p |03��s
�4�f�y
C:�q����/ye���ۇ����üb�j�Y<�K8?��pO����	�tӸzH���F}<W� Ed�9D����<�is�zL_sq�����V��Y�#���ͽ�8�SM�"d�u?�i9���7E��yh�j_NN{i��0e��P����j���w�q�`r�J]�438^K'��	�+��l�W������s�aS%+�e3Q���{��)��!��:q�ﾒ�ҟR=��'u�?u�I�r
�Ï�'�1-�d�"��mD�P����)�D:���3�c�D�%I8Ǥ�&uX���L��E�z�Q�t��6���̹r?7=��q�I�ͬH�'�-���`�]�N������#?�I$�,�vꨗ,��z�!!St�>��pTB�&�%7f>���`�Y-�)�W�昲z/����B��v|�	���a�'K�0�G�B�4n�?jV�K�[Lҍm��<喂��;�3��?�){�$6�B�9����yAn��-iy�|GIJ:{y�
$מ��|�"+��!��9����f�oZ�+w�#~����L����c���!}L^�`�,zP'��wث�������Z���g��k{�ȣ6�fF)�i��UX�T�ђ*��_����>�"�Fg�D6�$���J�\�>]�aySf�΃��{�E�C�
�{�F���F�T]l_�׍�5�?b̸Q�z���%PQDE�1���-�*ĕm*{����j�aI_��%X��	Ww̓�=p&Dڕ�F4�u�xH2Y�gj	��0?KZϙ׼$��Ǿ/�X�:�})x����2!���j� +^�r�d9̆���)s��e��7R��&|�r�K����`��
���d�+�N�@b<�)��_E$��E����V>6:���/U��8��0_d�\Y���'5,F�<y?��)��3��UZ����'sW���	�m��6���'�lb<|S;��k�=/�w�$țEvʺ��D�U��j�Bi���� ]}r�O(��y�o������of�o��[z2�9�J��U�]IΕ�7rhn������Ú'�Hp� :$�R�VÚez��'r��粲���E��ʛ%��\�!h���-���D�*Sy$����/I`"|�y���Rî����n��ŴN��w�������Ϊ���r��A쯅�T0���
E�<=��	��"ó���'n�X�Ӣ)\9�U}�yw��Ք�1S<�b�&'X�\i#?2;W����� �տu�G_�hg�!r0���f��������i�����"���t4�c,�E���S�Ң����r���Vq�UUM"�i���0Aִ�F�r�|�X~D�e
���R��\́)?�]��t���� V�6{������ߔD6lP�_��զ��ޢc>���[�q������u�hk�	�1��c��4z���ȽG����dh��e��!��f����1 {�_3̐X�9�I[�p0P�ʱ�q�� �A�%�x�e���@_�b#9Y�>�~^����FQ�t&�'Ib�~髟���e�z��'q�㪃��Ι���m)�d�����j��U�Ѫ���_G��w��ޞdd��S�� �X���1QG�A�ȕ-8\$��7Ɛf0�����tkZ��vyT�DLj�8c^�lߋ����dx�-X�:9���'��-˝.Y��v,�Q����sf�:O6���˓L42�)�,}�ۡ��f�����i�����6v"ܪ��(��e�TR�����
�iQZo����,v��Y>��>���\tv\[�W�uP��!�\G
�~ʰ�u?�}#�l>�E�V���B[���x`g��df�:
����`H�����������Hh8[,#���t|`��6ߘ�"���e���͓�0�i�%P�>��?�z���U0ٍ�r����y�<:+�f�66�q��%=�ıx��=%���ϋ~�n<��w��,�q��s�����횩�;o�Fh��Ɗ��$�oի�i͸Y�"n���m\�޺C�NN�]4۰jH��V�W�� >�Ⱂ���[�3�o�l4�ؽe�v�c�P��?C���n�n�T�CIǙL:?���˿Ua�!~&o<�*-2�eoX ;�#�c)i��E�}�D��o8�9"���BDy�TH~�cA�(�(F33��k&��uJ�����Y�:s-F��Lr+��M�1^�;uN��v�T���,�o<��!$Ri.�D*�h���D��IB;\�=�%��f���O�!�g{�ط�U��H���[�<V%a��즅3�-�@y͹\^�(c�Wl�����L�[&���`�nd�`�_ܾ�J�����)�k��װ��&pe���a�����Պ�&k�Iϲ;��ɼ+	�)z��I���he�)�Ha�9^/)B�hU�"�$�"A,��ܸ����\�'�Q
Muu95�7q3�8hޛSz���8عuƎ��FS�X��er�g�T%a�{�?y�:� R>�� 1j���p��Z�����-�4n�������h���T��'j���$�����CUT�2��Y`nx5U	h�L��0|F{����h}�>���S���nD�G��ߎK���^��0��^���Z!�m�kuc��5�}�ڳQ�^M�da���6�pBi�&����k�D�*a[@�lwƍ�9���!�"-�K��	"�
rC��z��<"(FQ|��9V��w3�I� �C�/n��w�}s5�dܸ�KR����dOE�IsYǴ��Vȯ��0}����Π��	�k6�G�������y������JU)f��1�5�R�oÊ�	�Dv��v�d(�`����q �%�:���i&B�����SYPM(�i
�7�HmK*$Li�9V>%�,;�A\~m�zo� қ���[�/ś��n$�т����O�u��-���M��M,�MB�`�o��\�g�:��Fc��D+*,²S9ΉB�����:����RDڈ�`ʼ��v̐+�ѓ0��Ic�#��LJ�l�q�s�����}��Sk�=�V]�L�\x�	�7���J�b^\<np�_���"<p��̍⩺��M�L�'éSn;��R�s��_�p�'�#R#	򝂢BC�Zn���O�p���$OS�����p/��$�h���~�[����47�A:�V>�Bk��55�ض�U٩_62�I�T���/��	e�D�{�@��5G����}*�IP��3G4�ځX��W�t׏Î�`5���x�V�vvGr�0�Gs�bH|��YALU)^�Db�-��,�9�$�G�i�l�a�b�d�!�"���P�s����2|O���@�z�'����# ��U���ƚ�k�!��A���DJ��sX�3�;��C���w������9$!�[�C��-"��oM�����K@5����:���e�2�m�SdJ����_Q}�=H����öt+��~�ezC$\T�T��'�`������)0� �����R����vH�����?l<�'�;	1��`�ǽɞ�h#ϱ�3��g� ¾Uf{���u�=�#;�{އ]Ҍ��;P��;��P3�Q�t�.�{̾�
'���Rf�a�3��{ՠ�S+ѡf-_X�z���Q7Y��G�Hh�V��g���J��Jؾ
d���r�]����(3nޛ�Z��U2��a[LCtq��
k��W�����L�4x�ۚ�+��Gf� *��$W�t�]�N�@�pc�36FB�&$��H� =���w��6��xr�R����6�����j�˚�q�{�Ԋ"b%p����9�>��WUԆ��ݺ���,����=�W�iS���ĩP1f�`��iRR���n�D�"b�x�p�!����="v�'kxn�~���Qh|�΀��Rl�8�^7��F�DG_��å*�����Ű�TO�!�
$2P�q���%A�:Z��1�Y6k���v��<����p�`s4\���-�%�_��i8���A�{���M�(se:�E��m�h'U�ʳ]Y����I o�x��K_I������rX��B�!�����p��N��>��5ؾ'��B\�^h��WO�;Y�,�A?8��i�Rz��D�)���t��9Å�Ý ��|M��n���8ј���}H����[��8���K���/���U?�>xh��J~�8�Q
��P�E@��)81O7���N9g3(���f��yL�w�,���?�>�j� r�2����'�D&nX,�SIьC��+�-'�QV��V�RB�~� js�ƫ�-�3�4P�������1w^�ay��s2 �E�T���Q�=7q")Ӕ��y��EB@"\�{���C�g�۹_A�3u�����o�ܛ�*�N�-�ЃX# ?]b��j�톮�W!���������b�b�����!��`0c�9D��/r3z���3�۬o����A>,"$�SI��ĭ�^�	t�L&$����8����i5�������&N~]�%��$��O�cw(�Fy7g4qM�Q�o�bUl�����=����:yF��g��,�2*��hD���o]!��
��.Z�iBvXu�[��q'�H��E�46�{��Sj�@�_R��A�ۘ��A(P+F�;��On�vqE$� �����y�(q.��ǆ
 o�o��M���X5�Q�������8���!��]l���#�ww>*`8�eH�����z���|ܥ#6��ux8���p�LO8>��Y�뫡�������ۂ�� Vbҥ�^h�-����U�3���X���B�L?=�E�#%1�c�)U��|v�?Ǔ±!���V���9`�`}L[�#�y0�46�y�Dv���
k�堣=��m	;���S�'_@JJ+�O��O�����h�8O�z`H)��ˌ2��Mx��~�pQ�SٖƲ��l�d���ک�)��f�e�P�"Jx�^bF1h��ۜ@QŢ����*!X繟�lBlݲ��͆M�jh�r_1˓��=��gv�..�!�F��Q�	�&ܡ��Uz�_T�3�F+GIUȳ^J5���t�A@E�/}��O7�|S��r�=��,?�=�!Q�ߵM�3����� ��F�������g��x��P^ݢ����I�������of���������o��Q�<��<��|��I������1�r�M2��a��N`��^�"�N�W9�sM���!����v��p�O���Ǡ���N�]d��b����T�Y�E�4G�Yƿ���\{��+؃k�"4z��o�?-�>��	c��K�lYp���z��kY���C2�H��L�N`�ث~�+� �{3��4��c�F�i8T@Y7ϲ���39�G��z񖦩�ڶS4�r�}إ���>Tr�I%��Q5�4/Z��԰ݡNq�z�K!�r{�D+s��xG֢A������K� w�]��^e�(���7�;�*f2ߡ�$^q��%�ķ#2���!&@5- xG>21.�[�PƼ@�oYt�D*!�j�E7�Lj�{���ў���dӇNuDBmB��-:�A�~9����5�e_A������Ϯ1Yr�y�W���������2��K�X'!:!�X)��$�c#`~��u��R��@'���9ⴊ�l��:�	l�Q>�ޝ'������y����|���-:3������!J�+Nb���>�ƻ�M~��`{����),2g�I}�m�*(�ʡ���O��#�3��۲!Mϐ�A�N4����R}���}����|F8C!���@j{�YK��=Ը�o�T�����տ��@HA��B_O�}�_&+)_^�&���|���e^��	O�N�p��h�a���=:g���²��2�~~����G�[��>���°��RC��g�����(,í��W���cu�%�����;�籈W�ؒp-Ĳ[N��P�"�~G������c�e���R�Q�B<L]K%񜻄ME��@��G�R�N~Q;���&��״�>���,NY��2�H;�ŧv���B��_8I��pN�%f=F&��pkiH_6�N�,1�=K5��y78�g��%왖����6���j�{�����t�f�X�xR��j�C�t&\��I�"D:P*y4�w���]/u�D|�8�(�W�������Kz���������4�&I��9Q̂� f�����\%��G>�wF���-G�5�(��S9k빳�5����ı$=�Rv�D��eU����/��|�����3.daL��j�T���;�3-��%?�I'��ܡ�P��h��};�2h~�Nf�,����p�Ď#D#pUȍ� M)�Ӂ��+�BZ��2L�����i��X�n� [5�B�Xgܣ�⏌�&��'�,oL�j�8[��x���i0����(nv�jOZ��
s�F@�����1�[s�~��ڋ)�]���$���"��0#���-|<�	X�����}I5���Su{59i}5��6$�m��7�6%7�W]FM5�{pX8�OSM�'������J+��R���1n�_d~2�s�.,PҐT�'q���٩�f�㺬5IKnQƔ�jV��.{E�s�K:���C0�z�¼)Y_�քZD�^ 8����V��[=\4_x�����.����aK�ͨ��$�?
KW����,>��X���Lgn)T*�c��$?�Z����?Թ�'�-W�M��#NA�j�ơX���ƆI�iޅK�з/?8Ğ�4��.�W����2��;�M�b��7ϲR7�l �� [��J�N�-�����52��^�Gs�Ç��K��j��_�pٓK�8�Dx��v�uC��lb�D�!�F2��v�>�g�i���pd#��T�Q�gM����zXѓ ��g��Tp��*A���e���@���B�3Z����DSj	5�voez�����I̞�u�A�$)u�}��M0Y� y��p��u0�P��T���_[���IЃ�6��S�O�O�[���ܷ�b�Ml!f��Kw�T��W�x(w����l�)^5�
�$��x�m���95ׅ3���_8��/8�}j���
?%@abn~\@�/��Ҋ5�_�*x��@!�M6t�|�}BcVr+�B���M�pi�w,��;�9#�d"��q��-��6��%h����ɟ|]ꢞ=6D��ϋw����2b$���a��;R�3�����7�Њ��|��F�0L����=��yU!"���>��O����i�H�[j#��8���ܐ5�a����{��7�4,P�)�>�2Dcb<F��=_D!�~�{����v_E���ݷ)�Ɣ�K�mUF�����7-��N{.�!B�%�0ն�ƌ�G_�}�r�$��U~uC�I����SO8���[�'7�]O
�T���̞+bq7l4�F:]�ڠ�Y�^D x�w��}?C��<���l0�Q�H2@y,���(�)o.�|P7V�v7M 4c�܇������)AEO$l�^��<V��>G���.����+#��
x*�.����&��h���d]�=�E���N����q��O�`���`P�!&zаz�>���:��u\�+�O��V0�e�J�eX�m��+j����3�Ƀ��SV�q��&��|�z��h����}��x��b�'��L v+�c������[�r�`b㱄k\�˂c[2G��1;)Ɗވ$h;���c����3��F2�8lb�hb����C���x�T1�ɚ�T��-pv*G΋�����P�sh�V�8pLI���<b�g=�μ]l��/�*�_`�;v֐���3yJ4݊i�Q��<ɱ�\�јA�SQ�=�2����(�M&].�Oy���2#)8_F&H2f����;�ș���j~g0Ǡ��O]vxewE=�P%{�.}���
2qm�#���M��D	����,f�Qi�*e �X2�ڪK{��!-3�XA2���9)`��@m-f��{r0���N�0��'�&rr���8h�hT����pJqB��Q��?̉���-�\���S��%H�Ku*Q����Mv96hM$g�ԗ*�p���AfP�<-a�{��E��q�Rm#)w��a���� nT˖!/c7x:�ņ,\V�,B��U�	|��p�]Ğ�o���[3 �Dk�)�n��
	�>@���֜�.�ֿ���c�.�q<�Cq���K�)� ��dL���?�
�����?�N�%��Z�D2��g^�9m��_��g��'6��������c��̅#�	�c���m����E
��ةˡ�>�]�nSf媰�r�u��m.��D�B��s��D|Tt��kt�<�R_d�T����������B'={<9�u�T���N<��1+�k��'f��?	����qH��z�$�(ځ���a�u7]��y��e��na��3qC�[�M���$\['����]x|�?���ީոs�6X &~�Uk���̯!���"jd�����PC8�����Po�ٳ��Bcx��'����c�O�꽝x��H5���kCF ���-�ؽ:j�j�q]���R�Y\�q�
au�i@�J�@���'�d (��?���]�sw㬘Ɓ_��C��^�Y���k,9��y?&�š���!��{I�rXt��j Oϊ��2~tS,_*�䯑���q��Ds����!�/��;�H��T�@7l�!C����˞�2o���������#= A�7�����??���S��ϵZ���;6]�]2W��?G���
F�~�����j;��, ���Jp�k�7q-��/�t����Fio��eٖ���nA�P
���rN��I���tٟ��r����CU�f�C�7�?v�'J,�p��h����vfZ�����Q4���zm�y��k��6k�]�8�����=�X�H$¥
�Q�G3���V�M�.k���k8�"�NJ�"/!���kB���:�x��F���7 q6�:�	�QO�BC������0��N��ҟߚ*NX�;�6�؍~�w�Q���u���%D���7erAu����@%��K�6{ ��԰8��������@A'Nt���p:�p��V�\ҾGù�M��{���A�����s*N��j�Z��r�������(�
���iH�y-�J�o��a�~��:O��Uz��P��=�Kl���+��h�$��9`��^�ĳ�JǗP�/�~r�� g�GR�H�������vsÔF&Q��	u�-��
�Z��T��Kf�hG[���`/sئvP��0��.{kNǦ�V�_k��nG��t0'�:T ܖ2��Zس����Q?8��{��Xk��E��e:H�!O6��X�1B�zi��ȗ���������V�7&���T����9ۻ��(ܲ[�W�w���_�>8ݱ?�_���K�@�l+AaGX3�Ԯ����S��җ����)5�d[��N�@�D"k]C�|Lb}j �V�]~�>�k"{��L@R���dX�,�"�)	!TטO���5h�h�yx˖*P�P�TMu+�3f�6��:�19�gbђ�b��[Q�B [<$/��ñ܂cҠ�@gC2�����Y+u��}c�gl�vW�#l �T���lswD�$Q�e3)��zϯbP�¶#0gQ*�t�e�봶�a�x6��ȇ��k�(���e���E>��}���_hs�h�������Ĭ�s�Q���� ��\�X�1\��7`lR��T �kͳa�dh�"��N�@��ѕ�,4���2�;I��U��@���TT���Ӻ�a�_�x}��!́���͢��3|���P:o�	
�c��'��_2B�fL����T���lg�p��2}ZG����뤔�G�;m"y3���_����S�����Qn�Q��&C�r��	��t��}���/��@߈����� ��R�������i�vri����F���G��̑��%	��X,��_^e?�h��C�%�)��$XK��CF�<$N�ĪY�]�̕��@�u�\��N+ <�"�S�g�C���~JӦ�����Oq�1%��[I*b��	a:޳<����M�x�=}0���a$�����oA����p.e���m�ID~N�%S������'7�M�;"�
jn�D-���B�G��)����D�v�gup�')�����m|�����|�J�/�9�բ�xsIN���w�s��4h?܄?h��}�"0?�BWɮt+�{6�����mx�͝����w𸖥��=Fo!κj��r�"@G��w�T�%m�#Q$��ԛj����z$N�:C���=(��GT%(�5wW����
�p|)sw��^Nǒ�ԟF�.�ߵi��W�Bv������ش�3)�B�C�@�I�d��:>��X@��gJ|����:o�tʮ�r�|1� 5�5�193 "�ys� �I�� ���KK�8�p+Q��.��뉺ĩ���޼8���Ӵ��(Ca~�(�_-�r�c�L�_i��ɬB̙\R'�����
��;;)SC��I ���� �ս�V������m;�0�ߗs��o�j~V2c`�F�ܦ���2>�+L��d�B��Z���37	�^���3�/�8=�P��n"����	���7s��8��`�v�O쳡��XYR(É��I	��z-�>_T3[����D0�O����?
&�؂�-�a����,XŢ'�Nf���>.tÁ�1WV6с�N?æ�v ���g������n�m"9z�N_��%�o�$�p7pq���~f�HQ�%z�1��,�6����xn��e���x:�"��9A5a�A�c	r�zQ��L1N��T���B6���Q�ѹ �&�p�Yg�Y!@�K�%�31�9�<T_��ŅT��$<�i����#�S����Q�0�v`5�����Z�L���������7�C�SC�������wɇIRђNzme.%|�R�1Fz���4���� |��C�������-Y�s��˺�2��*r�~~�Zp���������8�_mE