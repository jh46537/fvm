��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\Z�;�j�A�r��'��+�n^7N��C����8����f�Y��T�k�I-]�g޾��s���SoƏgk��U��T����]�i ѣF��1��&��h/I�R�^�k���P��Y "�Ҫnj��-Wi"�����z;����y�i��!��	���QG��[�L�nb�0�p�h���'OvŸ�~����&��XLXB�v��ݘ����@QH����cy�����@|�ք�5�&w�m(���	�>�M�9�Z�F4p\~n�G��ż�:�k�p$���ܤW��d�#���l�Ag24�t_�-��K(3ƽ!�c���lg��A���7F�,4:MH���f�(�_�B��2/3��XCJP��@���#��T�׉�2�NÐC��l��6�@�b���D��X<v�1F���>���f3���K�������ID��<�/�����q��H��`��y��/}�@�
0YQ&���=�W4Ʌ/����P:�/���@�yh��0!�ä��u¸�X)������iF1�|�����/���z�l ��misU$JC����6[=jE^D�'�ʽ.�U��M-���Dd8��b���d&�?��A&{�b����O}"�E�WIB0�鵁�d�>ȉ� �.ۜOi�Z����t��OU��_�I��F{��c=6|X/ӫ!l���'�`��?�1�G�U1�/�e�Κ�(W?m�'�G��h^4&��e��ֱ;�6uN��*�����N�3Y
���� ��|���g�Mo�2 
��(אV�|�P����Kׂ�1���܂��\X�O�fe��y�ը2TT��G�lN�U ��i0�O"E"�q#g%�g"��
?%���)�(���I�ILL�}�	�H���hݏ�(��U�1�]Gw����(Z�ET���� yC8h���́#��Į_(�ެ���/Dz�k*��j"�9Q$M���Q���ٲy1�3��D���H�+�RP���%������&��5�3�hPh�WD�{(��Q|�1Q�^zRU�1���̯��b8�x@9�M��u��%ɌO���7~��c/r������RG���9�Zclz��oYP��*�Q�)U�>{�3��T�ԑ�Eh7z{Y�4%oF3�8�l�Y�P@S�P>)ɀ�E�t��i`��@D���/�'
�u��s�KZ$0���j���Y�����ߝk
��JB.a2WL�aw�mⓉ�I�:pO���CS��$�8�r�{�LF#:�%Q{����<+�ܬ���&R��ʸĵ�����S���n�7�������K����^���'5,.���]�O�F^�~ۍ�?��U(�ϧ�bƞ���A�J��[�D�{����&���vV��lf�O���h~������Y���ch_��1�ݚ"�4�P ��(1���޹�(���]h)�Ɲ�'�h-��A��)��g �z���w�\`�+r�!�[�����;/���tJ�`::��GCM���UXc62�,�6D�.�KAsY@>f:E�έ�٪�!�����6���Uq��{�\B���W)�{�j�ӂD�Jh�%y���H�'dk�j�p��Y�7�*.�9��{ ��t�f�1�1�\�P�~�/�'2�h��r%?��9�b�c*ON��)��}���G[J��J_���Æ=��yt� ����|W_>"��AU��9��S�iЈZ���gH��F�'��Yss���aC$�%���@���N�H�r�V��`�gl$|7��K]�]�NL��Ɠ�Өv�l���O#]�"�g�=�\�?��RG�X5XN*K�]�S}��8�.�	0#�Ͼ_�I �d��b�>Xs��ZD~N��W�1�� e�R��bxU����2���Ž+��,����s��:<�A���{:BQ%\F������]阈��,�����>�y��vZ��I���h��J���Rr�E����p�\N�z):�����4ua��_a��ڥc��,����C�4|����~��������_A�|_t���I�*	rns�\?'�)�OR3b��5��4�_��_"�l��Cc�`w��M��e���>���0��'6��zt�ETA���YK�T���=oTF�/�ƀ�G��\��6T���ctXF�y>K�����7<��R~7LWBw\�?�����,��8G#��\\ z�D8����<��gd�G�x�/L{t����_kt�
��M�,f������������<�R8�����ԟ-���b8�����!X�<�c'`�-k��N�܇l�7q�Q�8(����ɤ��
�a���u�&����-Y0��	�������&�	5r�ǣg�/?�`>��1���N��h���-3fAz���2?ڪ0^�r�8�Go��H�90X����lux��Wf�o���SC9�j���t�� �'��񁕳�ض��:�XcM�
��WI�t��
�Ue�uc�!��m��6G����Џ�K�&��T�{������c��mخ�u�{*Z30J�{�)hr*�.~^�䨡|J8]z�*�]��x����N�,]'��R3��\�-6�AI ��ԦW��A_5rA���O�Ę�����)EU���;�U����u��uv&&B�C�m�n���a���j�g^-��'�
��i2�U�IN\�f ݣdüu�ň�"��\a[�X�X����: (�%�L0z������l0)&A+�Wz^��JA&iI����Ǩ��xq�6����vg�����-�Tp�)�+��u %Zz�9���"�� �H��MŊl��	�Gk��O��f�/Uj#�=����+mgw���W�����ʥ��5�;z�0�G�m~����@����h������%Y�� \]�n�!湩=Tr��\�SfG��ŷ����] ԰��<�#T/��-�6��h��%9�bqY�M���jܮ��V�+�D,:� ����+:2�r�E���ȩ���3j=�ї�A�}�-g	���n��!�qEg�d��F=Zל��O���\�|�}�L��kz+�Rɑ㔺�|�7�DW�
F)K|ڗj���	Y��������֌��K(5��"	Š�oS�R�e��X8Ј��6I�,�.�b���Ӯ���@0�q�#��6�!���S�J M�
Vj �Q�EvN�=b׋��c�.r���r���4?�H�Vf�ˊ���Qɂ��� �p��b��	6��{8���x�5�yS��j?5��晿^v�s�}>#�+�#��6(����f]1��*�O���\,$��UX�o�}�Uie��m�k��e"�ȳS�-ǚ�"�M#��h_X�u�T���jvGR��c�a�HĸK	�Q�oP)�LoL����Cu�
�\1�ޚ��y�M�:%ܨ�DN�$�Gx���`J�X�X������Ƅ�h1�[�k�*���W;S����Ѯ��
	#�W�:=�5�x9�#����QvTg|���R�;�P��O�B�_�8}��hD)��%��9U�|	AI�,t��eH&���Pn:���q����p��s锯.�{�r�p��x��)U���� �L_�h�����/RŬ�0�6��mǞ�>�J)���)����Q����Vw�wl!N� ���"J�VPѮ��Zv�ũe���eҕfn;�2����Z�aN�Z2�����fR2�rɠ`�㦝R9f6������rel0C�0i�6���,��%�`���ٚk��H��7����D�w�� 8&^k.:3�*-��E� 6�8����=ǈh�Gن��Rz�B�mTj�"|�CHT��U���� aƽ���t�9}�����ށv�9���;��qq���-d�ޥx��^a���,�K���v?���F��>x~�?=p^�V��H�G���gx�a�&�M��1������BM����o����q������34��)���1�U9b8���k|��� ��ŕ�0Wgv�P���^@z���Z�����%� ��ĤU6�w���!.����-�S@�<�lꝵL���+@I�.����<{�,��u�̆|�q&�����I h������J0 �kxX	���5}���������Hy���AQ�H%$K��I��Qh��(tUdF��,F����@�����&�;8��WIXj�n9;rT�V�K)П+�c]����DY&�*M<�B���a�^��|�:�������R��{���V��u���x��x�J�cFz*u�W2Rv�Y����]��u,���T[d��Ƒ�G�)���W��[Tv9	\�$��3�恍92�4 ���C���m�o�
z�uYd���R|)��I٤��|P}.w�@
�/o�	{�c�u�;��M��3���9F ��G�v�d�@"�9u�_��xּ������9�,���lgL��jAB�!�W�
�]���U�B�����p��2�������]8���'o��ﾴI��\�V�l�����^��TD�;��������ޓ�H���U#�����t��L�!2�!�������=�u�P� �)2��4J�H�j���Җ�6�I8��`<g����ӎq�<9��A����5���!���R �v:��_ȋ%�,@.J-LG��ݜ���[Ĝ���墘Y!S����=�X| �V.'*���-�Zde��l�p�M<ބ�D-�42G�9C���?p�ԍP{��{'<Ȣ��^fm���B�b�} �-)�v�8z3�\��/  �r���sk�T�����N푩�pٲ&����݈uzYs�d�JZ�<`�e�4�_��#NAĞ�Y;ЋH`�������?��ꆭ��֟�������O�Ɣt����y�p��@;�?����9И#3#r���1G7*���
�����Z�5�ӧ_���Ӡ�_��O�eb'���g9�� ��	�\�h���B2�}p�U��?1b��r�:�'�v�jbթ6��3�|��,O@k2�1Vȡ���`��9)�>�8	�n8n(J��寚�Y�