��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^S��A}�N��G�޺��Mj�;c��� �
:� *b�����L�e��g�I�ӟ�?2-��~A{|4��˸ eu1�f'|E��E�W���lmE���o}v�NX�7G
��5#o^yb
�������KT�q�~'=�FIȵ�>�z�E�P�9��b�U�����?��3y<��r���:�J�0�mf�v��ڧ�1.J��T��V�
'Hy�Z�kN��M?y���S�x1�Ց��,��v��6fezԇ� :6��w\0����u�Zz�W]Y��l�*Y�k�H���Y<͎|�78�W�Ê�4eZ���HڋC�c/��!������R_������.��P��{��@�uc0��I�汰�ϻ��;�G��Xv[��?6���J��6���%�j[�gL����2��T�	�ں�.��zO�f���˭-���ިQ'
�I�8N��x�@�Xxw�����2g@LJ�%hLC<,�	���hΥ�=y����(��zɼ�FzQ(��AB�&m�*��D�Ъ�ȏ�M<�N��G1�#w�](Eg�y[:�%Æ��e�/ �O����/{L�B�v�+Wȴ��+�AqN���Ժ���0�2�]�Ts�@��-c��y��yZ�sG��;�� P\et|ج�i$����B��*�~6��=�x�.���/[�� tC�m����-8_��"��q^���
��V�}�=��tt��2��9!�Ϯ�$��z�8ʓ���BS� 86*t�ܣ�^�Q@(N ���;
2�|�vYW�g� ���4�:F�i?�v�J�vlM�}�O���9M�܋�|[yw��5%�yW� �~��ܝN�E���ׂ�޹sd�V����$��K���h}���R*�T�2��i�9��H����۳���৮M:W�#7��)M���	ռ�"XKa��w.�P����ڡ?�ʵ�?����Z�U�t��-@�i��L��S��pt�4P�FY�!�jѼ�T	#W�r���TS��(]��Y&�q�x�o��w�/�5���6.[3�*s�(����P��-w�b��P^�#���4ß�H�����\��1k��6�����&������P}�<@���.撦x�� �Σ�J��k\�Ͻ�吘I�מ��v��5f�y�l�������*�[����q:E�2ZC{8@N�W�Z�mM{�C'���r��c�[�T�,�m?js�q��tq�͖�#F��9�K�)
%�(k�9%l� ��4���JP�Y��LU$,.�,|�V�V�}G\�&x�J�#u�R'v[��K���\��1ݵ&���౻@0 ����r1R����:勚	���5�L�b��9�:Eq���M=�<]0�৑�jH�nv������A��pRH�y�	��#�CX�a�K(���uC�N��� ���ş4r�P8�SS�U�T�fq�{��e��1B�u'��h�$���*Ʃ���&���UN�m��e��}���_��{pC���԰"��@�8�Ne���gGx����X�9X����C��j#��;{���ۋ�2*kSS����_n|/5��cV�����{�*��хYM\�_����z֛��q�H[��̢*ge[�%�2�N�o�)�B��6l�L��e�x�W��1�ò�1ϝ�
2�'�$���6�e�/�r|�W�8h�h�=((�kiG�����y8vc�/A�ID����6�q@ݼwRc�0�N2H/hp5���<nMƦ�UfV���4�"g�Wj�~���إ]yލ즦��&:;�`^̸K��?��S,P�8Dx�h	�}i��0�bXVTL��(�����=т�ń��W��p�=��!X+ߥ�1����ID%Kkc�>�_