��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&-\X�ǅ�2�.*(VuMl.�$��L���}V�3��۰��A	u�Z(��ч~���yI1�}y-�py��M	Nj�?<$7$OA��ˇ���r;��_+"��g7�U��߽���?)��F_�BAa��ҴA�j(��>k0�pN�L�^tF�[��6��
M�#�΀�ԯ�&Wd��;-]��Z�v���b�S����>�aG�Hi5��2�T�T�?�}���Vʻ*V�0��+O"R(�vx��!�ϐ����q��1Q%(�������@��d�]{*Z�Bo���V�nX�[�O'5������v�����j�3�P#>C��ݝ����'f]�	+�z&�+�)�v�iw<ߑ)���+8<BLf�Wr
a�l.�0	V,pD\�"U���!d�PS|��^���öx0a��%`I���;�D�^FEM�:���[h�-].��?�0A-I�$��T~4h>��̓n��.��`e��`e�Zt�9�Q�[��=Nӭ�tc��(p1�r*2��5�L�&� 5N��`�,�q@�9�)-��E����MP�r���}���$�bǟ�ui:G�~`�y͹9]���'�V���*�����1����p'T�%�u��p�GVՉ��Z�7���� &���%o�9Ь��f�Ī�HZD~U�6��h���K�i��H�@L�kN�ތ�CJ������	�!�ޫ"F~�����̻��D�P{7~k��lv�X��#e)d崂����3:R�;�N=d�ZR(�o�!ld1�(rz�G��`�P�;������f�������ŭ`nvr�UN��T�=�E���/n�dUw�Y��%#h�FC�,!��}<���=pڮBw�'-5z� ߶�r����v.i[���ILK�V�bDi��4���ӵI^�(�H��v��|N\a�x��K�7pBwɨ�V�[#�T}��'� y>�P��!�~4�5�{��6�5�\�X.)������zu!�0�����x�^�=�����O7�w��f�7�9a�����	�a6��@Z8����4%S<�v��Kg��n�6����_��_�s�k�^�PϽo�6�B|`��������KGd$뚰�Am�8��J�u�9��y��Nһ�%��:_��ڐM�̜Z)�e� ��O���5�1jOr?f��O`l�o�$�T��Gisx'�5A��E�jW�J�ng��B�Z���>E:4hs�T�����E�!nR|�+���h�MG�ͳ�4��
�F��PZШ��=87��[[7�0_�3��1B3#>
�
!�90�ᘻ����������4�,�Z+�ؘdר2$y�1(ܐ9����UE��(|��|2�@�aVL��8��I&�Ej�E���ma����z^w��Y�[\
M���p�YD����!��s��5r�{�,Dk4�#�I�����9�pi��t+s�ǑO��ͱ��:8��+����#�.�G��n]so�"b�V���jg^�XS�̈́�U����i�SQ�\�������[��{�T�7��ڠVA��>��N	Mދ�xZ5z����&�,� �&Z�PX¯c}��2�
�Fx`��Kg��q��,s&�[����Aʌ�mƐ�wBkؚzjd�I�:�$6x�ױ���Ag�n�謳����"Zd#4��.���3�>\PU�������b?���G���E�3��Ɇf�,O@���&���|yGk�6�6���G&~z�E���5�$�W&&�\��(�Kr9���M��ǹx �u�HА1��Xs��d����4P>�����RR����@��������|���PI���$l��S�ժjܶ�����0��g=kp�M4��z}G�.�}� �i�{ZX�� �ϪV}� dޝ[�{���n̛��mT�|N����e����O�6[F˅����&f2D��R@F�N�U;�M�U�	����9��L�Ģ�3���E["�bV��w���c�4=M��[�E��}�h�/T�C��qB����R!�׬�V`�́M$�i�e���5��͐V���0f褣�7з �z�o��z2Bv??���)C��vLe7�Y�6%��������!r�zٌ&�^���HW��栍����VU�9����C���q�&ߪ<o��eM��������W�iC����;�S�3�w���l�b���Jʍ.��m΃3��JC�H�0wv�ph���#]���-�X-����L۰�ip50����\�ݭ'�ݠF���	�I9��Q�2jqf߼'�syhڽ)'�9gKҎ�^�:E�d3�ȧS������f�*�9�)�ѽ.�ʬ9<k���VTO �a"�T�b~+�R}��� e�X�,�n����x!~�K�Vd�d���M�w �r�<��L���CR;�Y4�"ւ8Ly�;�4�� ���F�wu���՘ɺ�<����l?�o�V�?����nIeO����I�usT�\�s��R�s�>�eL��b@\v�;� �����<��@�+�pZ��^��5p<3(��z���w�����/���,����(�.bi, ��@��Y��0�c�^~6��C�39��x8�5]�����<���Xo��m_���J�V�ʴb	�|xx�1�7`�R0P�'�h����%�KN�cn���0X^p�����F�?��Λ�<Xަ�q�p-��!vT^�Ti�������b��!몎Bݭi*����Ƞ�� rؔ�/>1V�J4�FF�x��J$�2��8��
1��f鮗#2�*�V&+�����$��CH�X��5������������(�9�H<�ˮ���q!��F{JM�U�g�4�ɵ���� x�~=pw�2�fV��"�����#���3�?�2�ˍ$`�1hU�v?WTX�5$G������e����J��#q�w��
���K��>��(H��YH�Ɂ�ݬi�n�݃�JA�m����/ã��CVČw��������L
ޒ�vFӞ�.���=2ͫ���I҉���b�-{d�(F�x����H(q��?C�����ؕ��)&�:�Hi-Fj��[1��Z�{��|c�>���R��dwj�*#l̛��tcoX��)P�
�q���?�;��v������u� h�($�LḰ��*�U�5�&��"M���WF�9h�9���:a	o����#��a� h~`*��*���T ��'�r���л갪�B<�1ye�q�̳A����Y0���1��M��ۛ���(�/q洵����I�ߘt:���h�� �tz�y�b��_�t���d
� M4A=߾#~s�rw�L�`�Zx�so���y��x�McU#<k�Sd�}q�Kd�2/�%@��>��ͥ�[�#�~R	&VMHԗ�"���,C���[_v���&3@��/Q`-�?M��lo�:��Uo�\�e+�,\��Ra������=���5�IY�C�A�T��7eDEٺ��ܢe���#�p��H�ӡ2�@�{�*VmvL5��dѭM��q���B�3���lV�tM�u5V�&$���5?Ӻ8�e ��*�Z�D�����Cro�D�@V�o3�=���$I�C�)g�<���7���]X��3*�^>탹��¢ �3x���l�Ǚ/Ѯ�$'�k~�%F�Ɖy9P9�&y�T���Չ@��K5j�� ��@7�fu0ˁ؍�^���8��e�$�����-�U����	�D���	��h�,���J�����֎T��/jEb!,�k�&�������?����m���K��̖�}�j�ڱ���h�.j�y�x���[QC������#�������/�4{M�X���=�I���o���4�0�C�.�$̶D�yJj#����%?�<���\2�����οrm�6�!Ċ�Î��D��Ԉ�I~�G-��eu����#�k6mL.f�8˧�4l��d��D�d��h��3�\e/��Z�
q@�I;�TIB��I�Ϊ#֜;�#�b���<#�&#���$��TŒK�5�� ����h�R�M����*��sg�N����=Q-�^�c>�۴4^�5jň��$�
�n�t�:�Q�S2�|aF�>&t�(��x�A�/��[爀
�\��rwt<g]��,s��;VC"V�j��f��3U���,WU���D��S�� l�7&�^ԹvR�a�sib���^�_��� �蒶1!8.���$�|DP������h�dƅ��\)�ĕ?�GR��<��(��q��W�y�U[�{����+b��qMs��]���ڂP>.Q(���)U-p�v}�nO�&C�qT�eV�Y��P�ส)F�l�G͔�C|����Ȧ�Ya�x���%sZXCI�<�ƀ�t����o����;�
�Q�8��>2�����!�r�/�������Mb]J�|���&�*��7��=}��E��q��Իb/��^�AW��W���%$[�lUT�뜱�^��$��	��O�|�4�=(Ȅ�N�e����Ԥ�Jq����%N�=��ٓ��Qq��l=��ȶ����CS��~�?ӏ�5������َJU�P��_�.��"��o�yշ(h��X?W�<{��\K&&�u��7B��c�Ƙ(��8if��@��`��h?��)<ۼ������4K�e�q�+Tߥ.���<ʑ#K�Vs��p��WA9:�!.&<�D���ի[UJ�
���K#ۑ����
nЦ�l�o�@�6%_�Ei%��'��]xҦ)�\�$�@�Ny�v^�x����_�J��+�j6��SG��.�Ÿ?�"?=$j�)�m�9�0wp�
#5U��u��� �HG4)�p]<�r�%��VNB	LGR0��Ԏ�S�|�-����t+�D��N�����j�򋖻 �v����Yo��({n�
��s����(!"ضp�!��H+�v��6Pwr"�����S�r���p����;}!�����(���R�tm�A⭔S][�}D4n<7��K���syi�H�V�r�g��"�l������6*HP��n��7�3B�1v{��aP9�;�We�U�_~c��M��f��
�P<�K5O0k9�3݃�"D�o��4?:}�ԓ��:�E�3�b�&3Ֆ�>�3����z� 1��eCGHJ�Y1\b��w(���j�ǫ���Yadz�Z!����E�=Ԯ[�f�'��&g���ۿ�]>d�KZd�ՠ���J�s�F�x����.��MS�@]+��Ad�d	���r�QʔA3���/�b8��| $�0E���|�(|�a'��e&Z�]�Z,�:���R{���{���y0Ժ�Ьߋ�O�4�Y�J�pA1p	��w'��0mf*�v�1�ݹRQcM���z�ݕ�+�m�5��E�5��۵�V�Km��5|�֌y���;�lON�P��������b��l:m+f�2Od�b��P���и0������Fq|��U��� Ko�H*�UiNN�_�bĜg�i,B[���\�!=�̀ug&�?���U/,��f��$;��zHҿ�إ���Ø��	h�ĕ�#+-��2<��W+Dq�>�c�Lj�2?��"n����#:¬�ٌ!�X�V�n�@0�YH����{~	��`�S�X�i"z	%��%$_�u7�n2-I俚>�Lk�
Y�+�� ؓaȨ�)����iq�Rح�1��,/��"�I��i��Uk,�-��1x���I�w����;:5�e���5�A�] ������v��$u�SB�|B/���^P��OA�􏴭!�>c$���?W����>t�W#�X��>� �7UH�� {*U%��1�,�X�&#��R�Ɓ�X������c��)[���ik�M�ͻ��0�W���Ot3����� ��b�^I�ˋԃ/�<D6&'�[��Y���y�����~Rrϲ��>p"j���y��HnX|�`�	����St�MV��٦D;B��C�����w� S��)��9��uQ��Ec�0�6��� ف���4�,I��=�=; 4��^v�<�x�0��)A��������\�c���:;��YbtS,k9-Cش�=�����Z��|6�v�
�naVia(V�=�T}�D*�"��R��K�,����=��آb�<77��� Am�S��5C��tM��o�� �9�mA���U����n���������;�2���T�T`��W��'���7
���wC�+o͑��.�_.�Gg$)��D�9�ҁ�/3R�J�kA�\��zs���?=��!}'���z �1ù�eYc%T���#� V�h�؅����V�+�Aq�=���`^J �(���ٚ&O��=Tִhm�=�hopi��Kݛ��q'���?8(�|n	P�YY��u�`;x�si!j&U��
ѹJ�������
�����*�W�G��90���\�ݲ ˀ���Τ�<#h��K�X��	|����5�|{Qg��=��u���{��ǚ��-���p�q�[s� �;<n��`˄z{��Yႃ���wC����͑ׯ���6L�\�E?�d ��%�&�!&Ϝ��%�Z�Q��͹d�A.���6��˙��Mx����3��-1#��𶒣|���	ˣ�
5��4yh�3n"]E�[���̜g�o1���A���)*0Y}��R��1<Ϸ M$�uXJ�JyV��q���c9�G�L��(��u緓Â��K����^�/װG�,_���J�D�J �X�&6>P���u��V����0���~a�i\���~3�@y-j= 1pWfƲo}�q����Z�k9�n�	NM�p��F�7J���?3�����Ҋ�Y֓0��P�R���h�y�����Kʡ6(�^���^l���!���lM9�`,<��3�Ss?H�S��p_1)�WH�����ri�)?�����`V쳶�#�uX�ֱθ��X����C�#����F� �W�X�%����6���i�0.���(Rs�[�n�h����nP�F���V�l�J��C�Qk]L�ӈ�̟rK�v��i���@������^�yZ��=m2�Ӗs���K���s�-�,�h("�<��N�0&5�M/��dYKR Η��K))䠑�ǵ�6�}1[�Ծ|p�[��~l\6��U�m��M�Y^7��6)��%�/�Sk&^�\Ze�5�nf4:@�}Qhm��j�:�<��Mn���ѳ��K���ѱ}��Y�'�K��P�M�b�{:^��ِ��a�9U���7�S�I���)Ov�&h�(�f5�_�r���	�|������'lpv�~�ԛl�\������fRx]������ėMV���1ΉHJc�������t��[���8s�з�=�gT*C2O;J�1�sj�)
`�y�RO���6��R;�Tf��<R�*��&�i���+d&A�r.E0uWǽ�ӷ0��������{�Lg2�տx��
����a/sڨ�fW�l369����g�!���=�h(v|���[nz�)��:�2XJu�$��zCG�<�SIP��3��`5)�9_��2na�g��L��F���-:l����4�X��[|eZ❣�0[	����_2Rt�SE���s&$Uָ�;�n��%�
�&�	4�'�Җ�0�˥��<�
�VBΆe�u��E�lɳ�0aN��z�Lk�Z!>�wQ��A�D\(���c�6�}��>M�_.�۴0�1�:{���pTIJ��U>&Ld���NLNs�i���b�Y=���#@u<�]zuX�3����U͋�,z	9*e8���i�/%�Ą+�%+�'rF���ʶ$<�̾{SΠ&`8ڔ�3�*�uB`hz�߼%R>�bq?@C��H�[p �Φ|FD�M��7��Iؔo��ho�'Sy�e*�yg�����|��&�����9���Z��y�U����ܻ4Rl�C��P��ŉ��M�V1�zg��#�E��,������8�܋)Y�i��epC���]\�����8s��Z8�*�0q�K���ǐ�fX