// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:37 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BXAHp35gPACG3qwPvPel5P1Pu2PajhPitlu8u8lQxKhc+o4NM0QXPjHfnzdCKaKY
X+wBws8lX01nuKxJeqmirlN1fz5ODPPyHiQKyqTUu8jMRV0I/rr8CBQ5IxOAwW92
/KQfFnupQGpec85ME1KjUYfOTcHds/idhUCFSDvKZ00=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7440)
HvOqc0+8/dFFgNFG649jYlOYPeqW0D2wDDc+XSKdIOVMbey32fBWzz/MB0Dzc1Rm
SIVP9k1LwMkxLHR7xr52t19X2qTh52qSE/rjed4toWU90GHjtb23FFdQdS0Y6sL/
GYS1EWqgCMz0dAdcXCVMBbRb6ELhLkhCgzFveXTPLfPevzFyZrha4tf7NrNavDAe
LWvoUSILvrOMT2TK35LaR+bdVPDQmzxCKLnlhnMm/KfmSg2/6xvrnjOSr/qN1VLP
TqcrAQVdM46aX/8j2fGlXX53Gy6yWmeP1W8c4UGXSTqQu44OzvggTng967m18KNo
ZO2vxF3a3NgHZvpzQjuEXinnPPrn08FF3TSJNrhMWoRNUGoNRjoh+0NPRrcS/sKR
/mZmOrwmbS9nMxji2k44K/N9r41oX18Fs93Gzf2uJZeFo4WmwBlyVYavgzIy/I6u
BL2TGTVJeymZhMRY+xlkgfSWUUtdv0gE2hDlTb8y4UhP4pmcbe+LhadLUtICYGes
Kje3vfnenQGHel+jBJVCiMTO0YG0FAvzOwmUBasftLvviSxrqfSma7wuWVFntqxC
pzOHe4v+bgOXKzLbjaN2nRpXVpkXpc1pS0RFFtNfrwaouZs9k8v8Xom83zER+va+
W7EbvJ+A0FcfoQe3vQgNR5Z0zJ1kt4KsR7l0vtYozvVOIDMfFrS0g47S/f5UVRsh
RmJ8mHjQOELf4vMRPjqiKTfZw21mY5dvhVeLfS8tsOlkwGFUF8QhwddP29YgwWua
vEy5pqZnz0ruxRCRpVo/fzhm7uAWK58U3xvBV9TaJD6OrGKfZLna/M8Hm9dAdRZd
BAIMO4uxZaF6VCmMRwg0qJZrVjO9rNZG1T1rNh2embBa4u3dfyzag0k/IYSE+Kdo
77ZN4GyGBXEd0XXZSrjXoXWwFgHnQzH8A4+UUy6YpNPknABSSf43FDWmn8l/BYxa
sau1CSQ0ZYDqOzpd6FamgqMppldz5Hd3RVaNb+XnmZDLrAO3CAWbDvDVCMY6Ej0/
K08l3coFqjPfFmC8MsHKzGXzzxwCN8FaxDl3jpjsQjM1qTG5MhmvQomljtsnDHYf
RIdXwCAI5GUrfNBGJnXDouLEgYcZdQYhNbWiJx3Zp16VAdY9EVIIDmRACz0ZPPr0
vgbQomf03eNWP12KIeRytltHE8ZdxrgEOz6/4yUu2JHb+SIo0JNSN5oMq/cBdZ71
QEVfqi7b5pbBAdpJYFqavsTBtmSufo0HEt9wlkTnFtpWc+4FkhB7v4gwsb9M4hi1
nnnkIlZuljFU1BFRpNDHVhrgu1SM4PMywVVJXD3g6kEm7yhDLBibM64uCE+i8Ln5
HOjL2yqUsHUtEIepEnksjpGBViY6Mhi/4OO1VVqmWSVv8MU81M8/R77uGeqjmPvs
KvGNKYwGGzvrkDLtYbx1U14hzBymWcqKevbZLq6O6Cmaelf9hQRFrKguWWhabgfL
VT1MujABBJSnsUPYMK+w2WciVDo1LJtQftaraFCQdSINaX2BSczuWs+QejJCSz8O
pF0q84qlMrlL2s1nHN+VN+rc17mEPi8/omz9ZeE6QJQ1HHV39Leva6KzOt4eZNTi
LJPPAnns4xylt0gTNXiOW67tdEKcl9XVUZDpKaUbUKFJdCCi/P8Lpllx8vWyascO
ucXgWiKkjhzbse6n6aNbXVAdfwhpSr7Q1S8CJeVQxqHekh7ng6RyTjnPUzNytqTW
GNxQnHWXUOQ6Be+hSn5ZslZNKCt68mDA8ezHeqpH82f3gh59Q7Kq5Vn+n4UUwN9X
tX8wtx0EexP6rJlVkEzEtcvXR61wZHzxSHc298Ep+u/nHh0mANkAs5DtOXymfmed
tk2c/5QsQHYV2VEogvmO+JXkfko4IlwZYxb6+/Y1/jJ1CW6OyEQpzEiPbZ2rrvgJ
O1JN3/j6f/+L6NXASYXN6i5FuqPuqNloUyQ2MNkA/OXmBPiaqrbvKs5LYGTJDuOP
J+rFg+FoDuNrtQXbRJDdHPsF3N5NfbB9dGcwz/ddZi3GJwgnPdN2tPo2Cq3BXEzf
kQs3rRVudSgYf4Jc+GIjsRvwlonqDvajlwWNZj4RdbkOYnJcbbkQblpwDSNFUCh0
pNR/D3o1/d0OdlnNreVexKEWdx4EGmVcM2OJAE+HyBePk011FfHzcnCch7c50eHg
kYzQze0/685qB5DAzAqAQWt4fQ2m8328orT65/m+ViZBHqSrLtB5idXneQ53ZTNA
x4ePFct5mn1rXkYhc/gxOiphzbYuZ1KgRGkdDMZr0DcCJmblwqp/gO2BxpvtPY2e
h8mimy3lfkh4XIIJyvHmeVVZR9cndVf9itptnYtCIpRtNZUvynOf8Og1EDoUpjiv
v45z3eNAdXcpdaWOeVi5EkH6RzRuEtv5g7srpCP72L4acqFPY+d6hDbVEa75fkwY
Q/lNCxElZYrhdLz115eO1cdy6qT7RK12lIif42hMqDBbmyV0NGSrzbOarsIpGu1e
p6g77wJkN8QN8SZd2qAQR26EoegPlBVikyqUXFPd0UR3qJgc8iTdtFaqs7fOBEW0
/hbmj/4fzdJ87SanNxeEHuJYbP3jwBF5vSePOoDF8l+QJqC3de3aSykmXZZ4LBll
39E9ryHTWstohSFZwchCePCjFB8YbUpdjFN+Jv1sRTgU0I7CYOCZtFOPxiHW7d+i
olVPToF5ADcahdpGScxA3Rpi45CkIT60VALlg/BFZGfo3onyNDjseoryu5sShPGN
6u6gV+HbNi3bPS2KHlzJB0otEIY5o5JvU4gKcJCbaGfCNTJ+NxWxRVpI//oTqmey
ZHIR6ufALMqRWCV5PsdPQ3lcWk+FCE+jmyrM2ms+fabvQlJ6xrp7f1DBivKjckTx
1Z5H2Zj8+JafDmktFbJzIrQbNUM/rxtss+rSSFPtS4A3lqMexWJMdG/+2G2RIZiz
PRqiUf4pk3bx12Vpo+GFjvwv3oowTxPtvzU0Pinhz92MfcKRb7W2IYV1WQwQqN+k
XrLncu2fEI88LUEm8QyCtjRbDsiKTIxMKzdyjyvatTcuFH4+cGCnzGzMLpRhS4j7
a+F/+PD8Cvp7EHrLZ3+8rtY/izLKlWOTNnoE/UjrlG/9niRD2/yahlChrxLkztYf
n7zdgrHoHxC4InCCx0qZRwIufCtoLtBekXS1fZ5EWE2pudRlYitMMU9DHQsib/HV
r8UgEzMhu2f+OAdN1BiHufdmpvdbBMUqcT5U4+801i2bfyx17xZbNIlWJqRNt6v9
o3yWGg3QEZYaMM5idYpbvHltzQgRFXluOelxRIMhq4CQ2YfVV6FGJJBI4MHuqsqr
cRttivCIN+nCLhFlUqmPsKSowTKu4NEsthtONxPl92q3P7aUvdkhq2KOfp+3ho1w
kwRFBvsPALnCHB6Q/LzaET1yNH9UOtOcJXvP/dw3vZmS0CTetFtk2Tec5KP7A1t0
KdwqHMkp/2yNU5EP0H4/iJYA1wtB1R497PiW5aBd1WvgLxx958bLvVi1s37cjD4E
Cn2J3BnST9Na4UYqaNkoO73Ei4NPxQyqYsBHzO4Wloxd4Dsvda5soZ6KG9KwU/rR
Hke/8I0gTCxCpvAKgAC8YU8d/FyOagQrPRyENE2Bzcwi1/zGDv/NCCo1gHkbIWvI
MiA4ekGm5IuGAqTxz5YsezZ8DIW/zuwKbr2aBtkwrF2kl9L/2cypobfzwrQ5UIU6
ST7vtBF/SKOQQ3xzPog6IpeBZQbZD7wZ3w7q7gcI4gy7hklQNpwL6GPyhdF0Oz8J
I9TBgQ/MIKhuhTV2qOsWdCq3XCLtHefPGDxjdRHsnBwLkr3WxvPxUlM9YjlsoH/A
Ocw9GRQNMGhxdR7PRompi4yp55W+zaFdAlNqTqu3PjTu+sYc/BmiBfk90/Wfv1yH
Xn3dr30VzD4al/FK+2tcCFY22fLygtc0emxCbtdLlbiF6UNzecB5iEQpIHix915z
o9z/iubGzxTgTKVjSreP3/20+1AmQZNCUaT0a2tAUcwExCmZyPq7a/OZRM7cNCaT
4mEXos1xvsGvm3tbSufleZcHbjmaDcMY8lE6CKRgmIIHzlZSc+BPvPcNSn15O22l
86A5pEzjUv4v4TAFims2ZvVRsCJfSAlE/C39dQTTcoSMTn1K2dUGcK5zhFjknmnK
2GAYT37TBQKviUnlvIQiC8XoV5jXDl62Z+kAikibkWSl/5pQEs4AsCI9jX+ST9KG
KkkYm0QPHxokaOFqKugrURKjMULtaRQzWMQG8jIlbBeapn0F81Eb1kUnWlHFDr15
fz2BNQ++PTl3r/2skqu+Tu3HhJBI1nCrnZ+qrSn3ssSl8PZgwAycbCrD8I7cIFEK
B26hQ2t6A+ImbNElgggcGF5AAuld/pXJuL6v9iK/FnDGBphpsnovQWyfjdpJSokx
2vvK/rt9QA52WRkdcLdKJvC382vBrNdA/d7nFslg7BbJlkPih0rbWsByqsZgF31+
StVcJirL5e0DPMaUAWy6wf7DUOQ0vTtvhjTNKDzGddDxj2MltwORqf90SXISQMYv
NEM5370afMDIELYq1rvuL8hN9L8cElsyTW+EdGLRUiBRG3qrlcWmrsDrUGxaWJxe
wAN4Hh3m4DYpFXe0T5zxDmj5pnIFywhwnXWIbaBS6m9Mlhr2mwxrz7+r0yMsrIFr
4KQFQYV5SnnP5nDyizbz6opgEw40Q3wW4D3aCNNgu7DebIelWQ7nGrVxGZT8E2pF
Z4dncOUqEoS3HWqHxanIHXR02CBLfTwoWy50Jo/eVr8zc4CvCoWwcJoic/yicOOu
hsck2QYHXg3IRnymIe/rHudkE21IHstOtpkB968heKogzh0LruraDxeQaHQosjd1
0arlOv5uPDTr1zg9trbMVIjAy9FTEnK1zVJZV4UXHouBheCha7SuFXQCTxPpC0In
UB2P/7ZSu9phDt7QyQZ0P/kA8krtM3aJLQnMuDhjiutBqaipgcoBapdk1A4GnGwj
P9pEmuzQhrAkuUmjQgXT5sSIWrrFOVAPlnZZ/IPAFLIgn/mXJHU/oI/ZxHizxevP
ISROcJ+FW+x2DFIUrFkm9rtIUYC0Kg5Ptao0UYX8fFNK4QQ9ZV/d1lPzq4qNqDSK
McW1UtZiWabHChs2FSehXbiqWHXr8i//XtNAr3C71ixVHE/5D5HD18rsiuQ2rR66
7Z92RAcyqF005AzU87bxBaEbUZAunlC2fhZCbIb1omqbEFMiwCraLIxoh8zXDV/v
bzILuPIJZfdCpnaDc/AMt8aGUB3G4c2oYWQSoi5s0MRrF7/6xS/7bZwJHeT7h9q3
+Bs8CyR/oTQUoqSWntECeMuWvsgHOMZjbAvAH5E0gNsyfSpwv4QBDxLeCU45pwhh
bx58sMh+KKS1+gnl8C09ma+yZtNaixOksRUFVyVJ+LWRvraO1fwipes+SJWuwcib
g5bcHHYi0uETnGgWTl1q2VwjL7/kPdqbM212oIhArfboHRu+z6vTYO0e93rnggDd
6OpFhXM7dGgzR165phqhDGj3uESlIigv9TEOK2byvOmg8J8NQJcv+e8U3ETd56gu
XonQHODN1eHiWnOoyE3CZcpwStnHzshwfeiQGAgMAVfTk5684FeDb8DYF7pxZ465
J/ozwCuB/UBuWIvExfirKX6WEL/NfTtTIdC1VocuUh9/IvIXFr91w00HFM74P4ui
28fWRpZbHXnnuNudzQwquMsh+JtVQxpJKTzHNnw9JF2LdwNizdeDD25pjN5+tG7O
Pw9s5xqXQWig9I62KkYkhoXFfW/U3FHFAJf+6Y+a+kcjZAyZpCJToe4n5uC9BR4R
r2N7p1jcy+ug6KXHL8Z4X/6PTt/v9Q3miWb8JOtz8bcpr4buFhw/MvbVuQcP6PZv
fQisjYouVM5KvlUvWz63NYuIAoPbcm6CN3M/85A71CVTuSuHZSIKNRr2jLgp8bcA
nvf6pZCxTix278mMsSmdYAhyXA9cQbeCb6RqeFFTNW4ZKIYAtIho+RUuJgQLNV54
cWabwNWIpqLs+vdw2FNNNT0hrQsNDOCEeB8PCat26OXsumYZLHX+K1FqaYNjIwxi
Q2CL5PVR73gpD43UhK9SKGyAJEbgtooZLLIdH8oSqvS8Hm5iys13YU5ux717MPGG
IcdN5J56VDO+YBOpGTjbARYvkJIH958qu19lmXo0ouPqJQZJK0jUOwjgm7WHE52/
4USDbfCrAJ1WzJk3hr1zaNv5OhBA3UWHUIv7aPSGPFkG9Fg9hpWuWGx7SXYY+006
Si/CrL0h+frhz6vZ/PS++jKYBKUmxtimduDe2dpyEa1BCtOdXJVyzjTPsAkwNK9s
94/2deZ88gY7/TpS+jDk5IVbFDUTlT01Isv1WO5xq+7MCfmez7YU7Bq5HK/H4/Od
8kcXLDyNWN0QosccsiKLsscu6fNDDhIHO3/9f5GS9sp6LLeppAVB6SqAHsS+vHRP
pEUfnY56+vRlxfGa07/Bqkcx/25b2ME5ABD3odw2ifFdcmi8nIEUNQtSm/rrVyP/
RZKUooRAMQDSfk4WrERu8eT5OkgDJp5eUEmOYkXAfAw8yUlR31HeTyWw4AmEylHO
ETdVogfztErCx5WA1KTX0BJuIquQboomPpeQLhc8p94yDQmXAMy1XAEB1y6/mmM+
RtSlaVGIpMr+7tjL0+xwfKpmKp6abmZc9D11DBOoYRIvXkEpMfJdt/b/WpUXUjyW
gPTalER8pa6WWMQIK5+6wsmmYZRmrWUJLjuHIthhgzlbLXLpuSknqGonLBosF227
76/oF1htkCM7cto49R0IzB5gYACccZKTZq0W4kIIgl5M/27bYA+YX9KdoyEYu0kh
Syh0mFWrIhOixqDJ2Qu3r02Zxq1COcJPxxF/SimZJ2IG3IGXgcGUSHXX3TCQHybr
PFd+TrObNNBdH553jIdelD3nysB44n2a4k28U5PP5pbxNTfE0T99JmIr3lF+IzUV
QaQMtPg+7aIGtnJc4/zQkFdHA5k2jvhy/saEPbCQep9ve7Zcpt5wPsnlB/9e00xB
Kr/y9CXn5Ex5S+MwpZEqh+0Cx5JE02OWRyMI0p8QfhrSvoQAQObC01t4zN2XnSA8
A8f7aYQi2T+OC3kFIrm0Se/eg7+Vq424EosX3laFI2YAy3CRLErPlF7wcCgDuHpD
ByTm1PG86s2mgkjXUL8DaeQYc+PFRvVv3FTxb84qgnMAKcFfMuLaUECXFNSH9sa2
j/cAL1PEn6UtLapgSbuzy7dQXrnmZ4AbEvRqpovnMM/IjU5wZ7HmbNWCxAFr+IRL
rzPe61whfqZprCKDqPmVR+OUqBU/ayCrcSIENZVkxfIHev6SofQTOnvWOvV7trbp
uCqC46fWbqE2T3Gipkdpa4LwuhyaTh/5YjdEeYkOnZX47tDEAwVYpf8F28JvtzBD
MIMhXI2V+FxnBn+nLWnIzFjYRb+6UPxBgnVvGRmzVS+liLv8SvAW08i/ehcXH3uF
ZL9A1xxiRJy/kNHqb+nKAux8WRj8VXzw1JAjG4gKlX8dY+itQ9ke/+pKJSIxhmvL
Gl7IsdwMePcF8qpocMxXL6dm2LgvW7JMlXWLYh3u4nwHJwnfGkXZ5rgsOj0uADsZ
Omy6BOhjFtJENVeJpg3RdQb5SRtUvGMeg8A6FkZSzLLX9tr5ildirdT202kqB6F/
+kV8fGyOi3IiPmD0zwIVlgr6ls+lzpLNQqlZb5kKdaUk5ro8AULKmLDRtuguoF+x
/ZYoNqEfI8hA/DoqkGYwRRG+YoelHk7p9BO7505x+ZZon9tcXwgErSGAGO+R/JtY
cjAOG2/yOp6FefNg4PN4wwFFxTIKU0mZ7xoqyFsFLMmRbiWPu/AIaIPRrL7+yu60
1/jB+yavGGTdYNCQvDY0CBPs8O6VOTWNt4ja1ZLbzvOlPRCdl7b7o49WL7VC5Nr9
7EY5cFft3mYykWm4WQvVZyQspaZAAN0dDSHSMhJpm554EMZ2KZV/eqTuwk9UD8AR
EzCd0OqkRMhoKPYlrAzUFfrr7LgpsgqR4/xe7j5aX0RKUBzXvIhNOW01fwB6bZKz
9So5v/M9TBEQ7X8F5hV9M17UMKpVU8anSc+jgUEaJwSQ+sEYXRxv7aCQAsy1vQgo
MVQFg/V0x0OWb3l/BST0a5ZuaImPcOi6oW/r/xGNT68Ht3lWHmW/8CnMhoV4LDxy
ezPgb4n5FYSXgI1wbl91KL1tkVFigFB2ebk0aMU9d6ob69yO6OObJD4Vyz1ctTP4
MvJds0mprPUvVnC5jS8SQNMU5mpKvRaLl9gUuSU6ZJCWB6Fdz8DO+S89A4hiu31A
B89XGKaoeNYkdPtDapnmnQ846fyyV8j9LqY1IOYAH9zx6z860NVW1/tp+JA578a0
4OEThhyX9e+LvPID6jZuMJGheryqHr8KeahJ+jfI7gvZa1MqGTqnRwiixEZRZMbW
KctKqMWfR4s59inumIZsxnzSX/c+I/qFxQmOmV1JssDpWv980oHsqT6xzMtIlBOz
PZTBeRSRByA11h/h/o7xPsj1fT/dLuFgP+IOey5ELnKI1fFFt0t/oNijtsqKuGHt
apHvGRsvKCuU15Ie0pnBeixaFO33y/zYGDpIEvlSss3TCX8rA4YPb0Sq8NWcTGBb
4PU0NWiWFjOw9AV+QYh91KfVQNuuNF0YWWuUwGA1Cx+l3boWvT5+WLQ4FzbpMh/p
4QFhNWDJyLeeUvZ3HSLA5ckvC5MGZNlimicMjDRh8hBXWishBRW2A+jWTOy7tuc6
ut8yUCKLyT1AznrtVZhQHTRsyS3S1Rm+teYZBttZZ5jpbV8nDPdo3I4i2UYeLgWO
pg0dfYU+DvjHV2Pgo7/5H6WqH4CWq1/4hzQT7pmMCvTYnnwKi30j+nAvVSi5HkSP
fSZ6HUwDGIWJSgeHAvsOwWjbbLbHTJiiiYN2a6GwETLlFlyouWqYPiyZR+1eingU
ctw038wEp2YZgVE+nxfns21OlLJlcfOGu0Z8Csg+zf0T82bpqxqjtI+5rpUH1kHS
lw3Xejwp1e7eZHofm8soA9ry+uZCzwLLfvuLnW3Yv0QCMO1rAQneyVWN2InY/fkD
fKp2LOWnzzCgDjg9YQiQjW7px9kZsbq5FzlhQ7BgOWCUlQmmlBEXhMbYKj+waCOi
ZxRA5Mnx3LrWk9rZVLTS1GkYJ8MZ/vWEmYb65vq7koLK25xrBqj5vYCH/dFbYkwA
/Lg5/MZmxwL3W/xnKmqIt8A3ImxEBqbDST8/PHY5+KocSK/EhX2/TGKk4mNEfI8q
L3Kn7OPvUjgTqL5yY0/emjfqD3W47Qacam9dU7A2W0SnKyxVOzofLCiT5pFS+X9a
tCWSWNWUvb5oe+Uqrp9OEx590LxiF6V1YMiT2BuwRtAzbBGBmUrA/PjXibiincL2
sYHuQlUwZWLLbPJryqmfnOPj+JJQEqYojPFwmceWOgU+SmEmC0uUsoFdnsxJ7YGh
1XTNTGN+jNC0BY066Uhnb6qtmZoO/9JcKb87h3TKKgyUqNa6DTbCdJgidL6FVM0G
eF5FoJj8SjgP7BNRWVTCFn9jRmWW3QL3wEcw5HbaJq5HYQwGCX2w/wS9txjlNf5j
1pVP1rRMcseKJhacu46qDFo/nfdr8TuiUpyJvE19eXJcryVquBkCdqG1qH/Nezmz
X1hJm6vbXTfqn3IJRl0aIYqG/nuqX5JUMemZbQ6fsE2h3Ion2zYpZxvV3liB1hr1
7Dpgi6hSps3DlFii8cmirOzXyobgU469B90I6mmdcj13QO4gTillIYEKXGQPh9xW
+dHIJ3PvrySimM1o0fJhVp6XVyG4hf2+knyM13GnIytRNABzl4c4GOjpicuZ33OY
WDvC6V9qbNWmp5y5Lc7ihzNBXlG9ckFud+Fu63o2SrUZGs7VdhSXjAWWTH3HSJ3o
`pragma protect end_protected
