��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK�PBJ�i�bNw�M��8�3zlc{�07( �E���t00�����N0�4��i����pJ�c�~g��~�KD-)5�F��D#�;�]mc�|�����f�B�uJ�bݯ߀�YW�`�v��W�v=� iI©�tFȲ�#�۶,�1�|��%�K�CA8����s����{c�1�Au(�`� ��	kf��ɶ-�`2�6��WP��z�T��DP�5Ed�eio�ː�唥���N��Y�V�S�iC��������m1W���ݤs���Yڅ�$p/��h���L� =� ݎ��5��E#����Ƚ.C/�е#:*��@"�S�����͏���+s��q�
�}�:P����B��n�[m}���%����%5��e�M�����<:��g;Ƈ���
���J��_G��Hb�V�a	,���h�fQ^&�A[Aec�Z_�6
��P�)	\*uP	���+J��"��ת���%O67����*ŝ�̀!�Z�"ѽ[����������.�|\��m�F��lAw��Tn�ω��(B<������huB6��b��9]�����9Sq��h���?�o���Ql��݉�!ʓ��"/� ��*=��������B=ª(iƀ�2͝�\:�����򋨖��sƋ�$V�-���ʂlv-죭����Y��K�rq�Y�d����o��U�ϼ���Ms.�)!������BH.LӠy�.ץ��J�\���^ٲy�$D�W�!0��UN=�.�0�~�qbp�n�>���K)3��t0f�	����-�q��=��D�`�$)L���u$����3�z.�1�� �Δ�#Ӿ������À�k�����W+��=q���g��I���؈��7�>�8�b��e!���[ן��F�Y�W&�W��<=G�Bp�k}87d�-����+�$j��q��O�u6�d��3�?�U�C�u'�R�C��l�_Ee�ᇔ����e2�������*
~.O��"uy� �/%�L����l��8ƛ��D�5?|as}���/N�zl/!Y�gDubn}����\
s���8"��w��M(3Œ:^�Gr�"WR�G���\�Z��0j'�7����f"�:(�w֖f��Z��~ֽK���2~"�k��ke��$��Rg,�5�Ƶp�eA�O}�򛶹1��y83]%�5���F������t�b�.���f bQQa>Q}w�8�zr�\��:����n
R����x�[DLd($��VȟYD�>
��(�fK���r�͢�'�9���A�J8��j�t�D�6�}q%`t����mOM�>9��_�\�ڀ�7ؖ�t�!RIk�	��{��)\i)n?��ȶ�(V�p�1�K����#s����ґX�؉:L�5��������%��η�RAr��1�w,/��42�3�����^Y��A�G�{>%$d�S^�\H��[ۮ�pD�}so��;�J�+L�7��j9x�����` �i�? Af]�ގ��ߞ>��q�Ξ��b�N;�u�F��"Vpa��Ap�����Um���w�t�(_'��N��2���
a%̻������+
�D4 v}\F��N���F�>����W����s�Աl�2蟶8Fa+��M RG����nJi!�;�v�07HL@�f�[l�&���>��[Qx��~�=�w��_��x�	�a�oEG�]�m��iiPH��Q8D���$���#�a`��h<|U��ֲ9gT�[���
8����tW�B�q�n��l��D%�%���T!dW��>����S��i�]�Ui>h&�ī�>��%r��7�kr
�vD�����_fA��FSp��{_�T}e��ۂ-Qv��@�{DN�3۬�0�?�(CSs:�4u�|�A��yVp�z@�;��0<�5��&�N�Լ��h)��;S�4��~��;!~C�� ��G�&@|�����,������W�A�4���Q���V%!�Y� ޳s�Y�����m�!��?3����A��x���4�dhYq��^%Oav���7�0�L����0��}5��/H��}��{�O����+OH����<��Q�O,f珑-�1Cg���9g��A�`μ���B]2p�|L�V5��e��Kw ���j+|�H�"3u�%.���H�5���*P�OC�.٣��]YLqd(R>;wo��-
^����x����ƞ��_��y&�8�����v��p9�T��E(��q8n�(�>�n�S]}��U�����1R�sj���R�Cr�Օ���Ƭ�i`#�B�?�{.<9�7�j*l[�w�EB"�x�j#�	�֟�,s�4����z(�dv7��5e�i�(�[.aP��ClM�uP���$G�O�y�NK�,�����h7�����ϻ%Q�1� �lkx�'�����ax��5���{c��M��g�*ȥ ��1��p��4u���,h]����7���+	�/D"��uk��͛��ōy�u;Kzj/mʟZ���L��-�H��KwiǺ ���'�3h��̍���/q�eޅ �!x��l��Y� ٬��=���i�R0��6���0)�y�tɿt.[rq��[VE�p�c_T.�G_��d\ɺ����yȿ|�@-�5�iZ|��m�
�$&#E�,����q�)z�a�6I|��_K�\�+
\t�:���j�>�a�S�.�%�J�	�U��Q�����OK�g�*�=�b���,�
����V��}6ΰ[���d���N\I[J�d^�g���Ъ��8��g}J�J�q�����ސ�r��|�Ů������+#WJ|[��̹f�c��1��,����S��TY��)Y3�^��N�]GL��v�>{,����]t��p��c*)޹��(���1�M�B�S4����m)�dp�%�Ė�I��X�d�L�Ts�����U#����Q��;V�.���x*�s�X�^�n,��|㞬5�5���Us3B���L6t�]1=;���Y��Z�E��'�G����X
	�`ν�O3�����o$6=0P�} 5P��m����+�Q���p��s6WP5����Ժ���.V��8���}��8��H��8�as�pp��Ki�A'AM�9���*�3K����
�Rh��X�/X�ez�d.,�!&rL��G���M�8��:ů��>1��&�-�{i�HVNBN.󺭔��)݌��t���'��އe�0g>�.��E�.D��a�E�ɖ};G�/��sD��!Nۚr8����x?Gm]\���x�<�a���k���*�����~�އ5���Uc���\�X-��k��\��|�K�e���w��F?�v����y�����ܣ���y�0Al�S���{����94��n\�侈��C�q�Æ*����v�蒶�O�:N�sW�<:�%��	��1�L�[|�Cj���F=mf�;�>ѺP�^�bb�x�Y0��M����;L~��r���2jC�@�E煥bWFN�fQue 6����G�e����b�~�)�q$�g\Za�� p�B�cn�/��_�6�9��dB� @[���� C�̧N��/6��Q�_��nUJ!|���H��adb��8߁�a�qxm�������L����mJ�R�� ����s(�o6��u���t �ڦ��w�.o'˛�Z�h���>�TR>/VP���ɳ�;���V�7 ��^���i�J����K��o؝���*Y��}8���)��D��ŵkڎ&H�F�^�^os�
�Q�g�����