��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb� >��6\��aJ<���[��?כ�4��n�^�V���Q	�ȶ3f�Y3⎌m��
��3 Za���i/�/��ϕ�0���H�ܽ(��j6�1�)���)8g%�o<e����xH��.�y�0T�(�^���>�:ܚ��5(|Ϙ4��<�p��>���=����5-��$^�Q�H�?���{������11����>�.3#ŃW|��4�S�ы�*߭8�z}j��l��ʕ^j��nC ��3@�H5%5D�r	p,ۘHZ���v�ȑ�pNg�j���_Q�U�U���v7Z�(�'�0�X@���#.��H@Y�"YԶۘG%����;��DK1�
���Ǽt�v���� /j�"r���/����17NJXϗ�����e�ĥ��hO�B���0~�nȫ҉Uu!��%(�]�ɦ�}�Ӈ���h�e:�S#�שR7-c�ƿ���љ�}5�M�mG�)lo=�T�%�Q+W�8��%yT�IOV�=��l��@��rZ�
�-v:ѯ� ��ͳ���kY�H���}�J~�M0cdQG��o�!7Q>�������³�LN&A�dT���cd`r2F�MߊU3@@_P�Iv����e��D���04<����U|K�2�oL5��\�0��eF�뎮��RRL���Z����r���h�0�	�[TO=hwx��#㳅�:u\T5&Y���0�_kY�0��J��",l5�Z�1
	D;���[��i�z��5������Sˮ��w=3�rO����F���`����}�RY���u��z�,*o3Q�lD��m�4�Y﯄��W��W#���w��jg7��.��%H[Z%��4Os���E�II�7�6϶�9��#���/�TAx��Ňp`[��� �ͅ�	[yl��c��b��G�T�7����Θ�e5�o�2��M��0ԯ\�/ �Oל���@oJUF�u��G����G�:�Æh���nm���7bG3uzCOT���O������.�<a�����v+×���+��p=j;�b�>��B����[�ЛZ�W��Ln?�8�a �#q/�6f�ur�s\<����}�wӥ}G�ֵ���5�T����M]nRV��:�{G$�\="_�h��V��DQr��32}I�$Xȋb>�d�{��?�Ͼ�v��F�>[$G:��h~������d)��f��|�xX���eU�(5��'�a�[���4��x?륤�{��D���`�\D艋�,�gjI�/)_yO�8�[�d0��~�<Ô�U�z��=����2`oL�;3���)�K��e#�GC`��q�W��l)z���Q6Gʖf��4�X�}���V�$eH?�]�X��t
��
��� }�?������&���c����dڀ�_[/��cs�ǩ|�iF��v��rݛ8}n���l�2��������ws��4�C����ٽH�G�4���K{[q
f �J��2f&-�c+V0�2~k��f�����KАI��g�Z�y��4��U�PZKzoF�����(�Y:>�:�Y>�A��?EZ�-�6�O\��K��a�@DTB���|	\�Y���QP+m8Ŗ�r��O~"x�=!˥v�k�`�N���_���������C	J'w>�����M�9`cM��}����f���k�F0u*����.¾���"_�Qn`�o���)��pp�,<�ܪm���q�oe�L��z�7�����I�����I� ��t�+gd �bz▉��%��ꟅXͨ�5h^M�>��啨�3�X��Q
�q"qZE]����2�
84�0ᗨ�pc���RF���F�{;�k��� ��ӭ/r�li���e���"瓰�H�p���)d0I�$Vpe�:��*ށ�?>d�+�H~I�8��p���?�҇�E}�lx�M|�]1u��MVF6������'k[�<�X<�Df���eϐs��
24�g^t5�B���;<�����(9�!�Zk���n����₱�̏����d+�,�)� d�]vF?�
B��ŒY�+�_ޏ�r]H����M�Ķ�q�b���W������j}@�y�tJ���Å��y_n�͌A�6�'��)�茮���_j�d��2�<+�>@s:f=��@�_W�_� k�t���5[��kr�J����k0�W���f��}1(�����3r�L��ɞ�&r�o2�t�U�%C�a�2p�4�L�^��{48]O��|���	�׳z���g������߫�x|p?�Nno�/��| �qb^g`�w���@�픾TB�OѤ�ArΫ���pr�HDC,��4�f�	��jm]�9҄~���7�Q� ��y_,�'��Zg91���%)��I�M]�a�C{"~o�Pq�ʤK���Mы������;�B�`��_\�,/'͗��1t�.J�Wv� ��?�Hӷ�*����U���1���G�H�tɯ�;������]�D��:��|�I�n�j��Ly��Hr��P�����`��͛��q4|�+�l�\�Jh� ���(�u���SP�1s����Ht�I���B����m��b�
�s�*1���}�-Z�����);/�K�f�$0Y�>���~}"fWC,�*�������� �trO�������c���s�A�i�{g����ГM�y���5!ً�O���8��_<_�j��w������B��3z�@M�����E~]�$2rxcD*��+��zuח�495BX&��Du0|QT͵n��,(��tB�2��_aL��>}�]\�-�g�����9��K-`S�k�z(��І�����O]٧AAό��a4��_^�g���Ϭ<��W5���&�	U�=t׊E�Cȯ�-w������%sn�QǿE��5�Q�o�aW�t��L�I�\��gO��%ھ c�zi@��7d����1s9(���ޛ�+v��