��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����:��=3�J�r	=�� M@Q �:���!+��?kC6U�T/���&��	�bK����V��D�Db������V��yfʀIG�D�Cs㠆�.�`OI"��\��L'1dA_���%��:��c���'P���G��4BS�_VW�#�6����ZT�v�O�! Q1�fX�<o��3���x4��̢�!i}���IZ���C} ���ӣ��L�l�,��Z���#)GO2��ׁ0 ���_y��7�����m��n��tGo$�=x:�U���������3�YX�"}�ۋF1�0� �-3��{^Yt_-����W1�>_��M�-�����������&9�^�?�ʄ�BϦ�s�V�gW��ĉ�Y@B��9`wg������t�I���Y�<���A�T�L�Z5p�C3Y���D��N<�;�n6��y��S�s�ok�򀄬F�͹���AU\?��\	pe�Ε���o_]<�P���:N��f�&@^'7
:1Ȳ&pۅ��4kD�
-~)�6�oW������nUD�٣a�#ܨR��۳�K)��u��@v�	�`R��`�6���6Ԛ�P�,B��u`�^��Q��>yæظg��!�Ζ_++�Btc=޸���[�����-�����u�p\s	�K4/�y#Q���K�3SC*7ʂ�I8�q��Y��6Q�m��6�q:�,D�L�i��f����a��A���0� *۱c�jD%�z��y+y3S��8a�z���%�&<����O�-yI"�PT���\^�s���:��@�^$�u�V|}��Yq�oH�Sl���@�P*u;�0<��w����u��-TI��"\�,��\��LK���E�[ �� ��Xjge��ֲ���4k
�^�b����┵lum
Zu��|�+*��;�A�O���b0-�gB�b�IW�0�>:��>����-�ø�9�n��Vph�K��E:Dl��e�[5U�c�m��a��V
�NhglO&,O����h�,̛v�a�o�8�D�7	��V�ESi�ZLG��B���t)��9�r����|2�c��T��dT�\hS��D?�)���Xo���4�^�Q;��U��N�T+��l�=��K�\�"Y���|�7�Q�]E @�d�0jЦ}���"%�����c#����7l,#k�`_Zn�nc��[�a��MB���b�1�F$.��]%v��Vm��:���uܪ?�h6%u�l�*iF��I����,�ּ��qʠ%/*������m�,�`����+M��=JïT��mʺok��C�~���)E�ߒ��5����r���?�
��a�ʲ��Ҳ(S�O����YH�0>p��Zh.]�^� �X>�68؏��R��;k��� su,���u��b�{�F,L��_�yH �Z�Yέ��*�Tcv	��zG�� �5�2�G&v�]{�qRE�1ݲW�s�B*ow�4�a� с�7�k�����Z����nK(,W>B�`��Ū��j���.�'���]D�G<�]h�~d��_x�D4~�%�C?�����06�k�����D^����4.-�Bi����f�}2���n���E��!*H(�νqֿ4�h���*���]n�L�G��9����d�p�IP��_���ќ�������k&W/���D,����y�{��4w4�Ǻ�����ҥG]h���WӬ<М�)`H.%;��v���%�U�[��RIq�J�H��L�)>��2	*��U�U�� -�S���p���xܟe�F���ybͮT��_��"�*Y�ްnk.7�5�u�`G�\���қo<���畉��xo�8�}#g����{]��U5A�酉��#��Y�"��^��;0kk��i���(���x2�C�TG֜	֓��N��ӾC����# x�UL3���v���y�‵K�ڔ��B�e�fD�,$ໞ�Sm��h��0���;zk�	Ĕ�����1�Z�!nH�Xi��I5���g6��(^h.�U��-���h*.#ŉ7�+7-NGH�n@�uy��vX�	����C����Kj�a���<Y�x�����A74�� �c��Z��BM9�ikgX��2�&B"���B~�� I_qm�4��t;��m9�����(��� ]�q��V��hV�P=�Z���,d4=�:�\��FC�fH^ٲh����TXpN/���a�������x�BJ�1�Uv�x�F
aTo��yUJ�z�x�Q�̰ߝ�ze��]<��T���AqO���j��\�
B�̅����|��k�����)��#�v ���� �J0�r@V���W�b�#��m|��]n��eH�e{�����>?e��	�PG�F�--��Ap*_�|��~���7iM��s�X���'�r�N�[��ػ�X�+���
��>C���8��4�����P��N]`�+��3��`�Dm.nFX~�hg�ɮ����9!DN�_��)����?	�Wr0DIT6X����Y+ָ,;@���	qu��4y�9ޱ�M�L9g��j4xd�Ӊx�~�����8i4��~��-���0�ṗ��YQ�n��RJn�`Ϭo� �A��:�U�}���ǝP1_O<4oM �j{΅�LO-5B�+�ye��z������1���v�+x�(e�G���$���߸Mg���+"�O��: W.�F�͉m�0��\���Ӆ�^���ȏω5�^���Ж�XTm	l�ʬ���������R�cl6#	�I_$4i�x �G�j���~vӫ�J+�����I�]�j�Lq%�]ff�p�;V}ʚ�GF8bH�%��1׺�u;�Ofw�=7�wU���� ���Zf��'��N��+װ�B96����"#���dNR�h�#� !�r�4US�b�s����o��ZX�a�=��{��{�9
��lyp|�`C�M{� ����M%4hV��ɺ|`=�\:�1��&9M�#�ŭ����&� Fl��,}×I�+lP�0ʾ!��x���`�a�&���D��f�؞q���V^�?���d���H*K �1�Z�)ŒkG�cܤw%1�����ے���b-�^��J83J�g����	��mH�sv1⏃!����[��E�귆��b�>�:	�R7�^��3��P�s@�J�V�%���A�%t�> G��+��36�M1)3�F�S�2^�M�K��������;���G�i~.!�K��7�q�N�^��d܉P�j���(�L~�Fq.�C��g��!��Z
u�\�k6{p���/�;�R��W]�Ig�N�d��6R����#1(W��m�F�)L~����0+"��-Z�x�Ÿ�Bʶ��g�W,$�GB��=��|�`xsh鼱g�$̣��[dt��Qi3bv��XG�����~�@g*�p�4�����D�3��G�G���J�Ea-�d^��-V�-���&�2�2^$���QYc�s�����|����v�Z'TGT��v����Mh�M{����a��o�C�~�)��h����	�h7�("V���T4�7�=x�!ABq���L�����-^`�3��Ѽ�M>p�g���=o,����.�W����C�ⲎNY�U��F�ek0J���o����CtxJT�m�}Q<����-�����&�#�)ʢ����9qQ0\�h���6Q��!Z:� k�Q`�Id���r*�޷8�߿����[0���va.��1.���RӫD�  ��iRPރ*JF|x~ފ�O����uW�?dW�y�`V�Y�:�C.Ջk=m���b����x#�pE���z��ȩ|�<W���H��n����BJ۷��?Q��ǖ���Q3N�]i�R�%��d��8ѡ�Ƞx���`�J��+������:���%��B�2n�9�4?���d��k�����Ov�!��I�V��?���{ٔ��qU��`-�d$&�����6�� �l���?�4["{��B7�C��]�C߯�@es�em�E�ϸ���#P��h��<���[��:���\��	%Φ�;��<3e�L4ψ��r�b�sN�����3%��ї�������[;��p�+v���8�6?(HzS��~�)�MC��27�h���W���n�Fpӊ=���Q�meq�O1��n�`��8Yd�rfd������稐8�� �i��:S�G��
�Ru: %Ӡ^>���ɘg��-�n��B/���TY����v�|HS�ڎ!�y���q�A��uf&T솀��{z���4��|���"���a��5��H�����-�{m���zz�_-\�XL�p���e{I� �ٴU�5������ōo����
��%A�Y����A�kP�X0����
j�.{��F\2F���Fբ�i�� e*<�7Qg�JF���܆-W� �x�]�8sM���і�,���"�����K�P�1�[��.!�|%@�Q6\��xx<����-��51Х�kd���K����?���#u�l�-!�}�6S���/[<���Z�H#��G�O�"��>���oL�KpȆ��R 	��Mx�9u6`#�����$�9��'���yj�'�Q�݉8"�Vu��#��7M��c���1=����o�w=�=9�f'� ����:�{J�SK�jI��4������1�����h�J�5�*�I��m�;���N|�?ð%y��>�zM�Vaf'����)�9(�`Ʊ���$�N<ݴ*�i8#��4�;�-�`��&e�_YM���^��a�e�cҗ?]�BJ�6LB��$$D�����'�'o������%��Q<d�wlOX;k�\�}�b�QQ1�)/���� ���6E�a��&n��p���g m��;����ۆmK���	����c���z�3D��E(^8�\f
b��8Y��s|��]("�<��U�8��ĵs�����?Lvu��Z��7�)�ߤh�0�&1�Sx2��4B����=��Y@; �U��C�`����E�BeL����������l.C_��Q���-�^oZI�&���qˇ8�C��)c3���@Q������r�痼�Cʳ��8��{>>p�丼p�!ʡ g25��#>M �1���Z��o^?0HvgS�셪t�_̌)�L�1�\��a.V.:_[��=�J�!}f���@�'��x�N�)��O�g4Ǿ�����mԇ���r�.C
P����8��M\X��	 P��S[ʥ�XCY��-���~��b��� d���lT�cJwvZ�,t�&�B���x,����5�5h���S�y�Ɔm#?7pўm���[:����ⴊ�_t�������{��+���ܾ(��\�L]`�o;@o��
�7��Bｏ����������U���c�Յ衐�d྄�6���t����J�y�ݤbH8�X�A�������8��l��V�Ơ�	ƴvف�C��j837	�l��[(�}u�i��dy����AB�4�g�COϘGޘ�l���4�����U�2j0J���g�U�����lٰ.�M��J��q�'�\l!������z��E�V9ehJA���8�FOb^}2'�5���[����QO�[cF�9�u���fLn��y{ܕ!w��2���)-\��&��Z�F��D!A`[� y�i�V)��8�mtG�|�J.\ߠ�������^�5�7��G ��dˏU9^�@�w�#GJ*��uӓ�3�Z�{�8��gr��Xa���,��mm�n(+���+J���ӚG�����]_0���j���v���n�����l��)��j� A�gd��t�r�WnF�w�Bmȱ�!j��W�k��T��cK�l���j)�m/�Y
h�KqJ�p��(�.�(7��"�z��-��?��#���y�p�L�?�J�=������d(6ɥ�u �0��ХV�p��;������@�)�Y8ON=8�W*R����y���j��2�9(��^���Yo{J���c�v�̟��A�<k���l��K@̍a��l��I��8�O_�������=�����ͦ�/�)06x���ʜ�/{M�M{�^Bzn�W���1!m@�<k�w���o�gO=J��Y�]#5�q��参��A�D;!$VR�j��䙍t.�!Ƅ�?�v��4���`���&�W1��I��II���[Wo������Y���]�I�b�U���*Et۝?��=�ɨ�Y5������j�>�`dJ��Fբ��/�>��{�S�*�o]y:[cg���R!���F�������_fbM]F[̸%1z��y}U��ozr���e�m�J���б�^�Yp%�%�g�2�W�7!��O��}2�����Ag����oTE��G3[� ��;�:(jИ���n6f�(?<����k��p�B�'T!&���1�����j��睳
�_F]�)��.6X6ev����H#pE��\p�zӃ0��XY]�9u�E��zw�0S��f{s���R�c�$*����/;�ή���Jn$U)�Z�FZ�{C���J��" ��|�p &�Y%��	1jl��u}�cv�5Ȱ"�D}���>]�YDJ:n���qO��}����������$8�B��DA���!���$B���S�T	���ݠ�|�C�N�3;�ks� .',�a�:�6$�R��O��΢�p=�lc,z��J�%�+���S¯=R�ɘ$�%�1��(�9au�W�
j�M5h���T�ybZ��4���k���Y��L�{����M�V�0~t��[z