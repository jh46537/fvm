��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzG&jI�#�a-&�2J�@+uo1�C��ID*�K�������|U���7����d���3H���ct�v�G�;��S u�l���g.B�>�(޳��#�Hώh̩T�CH1~��l�����p� F��|�t�}m�q��[���8Ne̛�z~�W�H�b��0p����
���c��v���������^9G� p� K�w��G��T��SJ
��\�ɿ� #��1��'��K��k�Y{��8VwP�^�e�"�ь#'t�{<cr!�P����ud�R�pT`#:�&j�H�C ���cz#��c���ԋ$�臥VL�&x	:����Ӓ�f�O���	gj��^}sx،��`�i�(�?�r�ĬL�UU<j�A��#�D�#�C%�J�9Q�Y��+��Q��M��� ����a��9��(�������ܪO+&�$q�"�i�4�f�Ss��k���|�s��~HSd��NZ��� (8��J�!��5�{����n��7�:�5��j�<֏�b0n@�6��G2�J �"���tL�C����yCh�6��?
*9b�k�F5�mz��<{�}��x�J�_�+�B��N@F`u�>&�m��}/������U�R�[j3��
ͽ��;ߪhT�[�1�"Y�"����'LҼ�js�D�G{��Ȋ.[׾ʞ�j, ����m^�5G�a}5_��zR3��Ku�����zS%�3���Hm��l��4Oʄ"��M߳4p0{ݖ%q�%%[ȁ���R�6�����H�M���K�2(�
��)�q�w���L�k�V���B;�m!���fF{������C�wZ@V�Z9</�� 
v��p]�$�·�_jg��-]�.u؆�	�x���;r�*z�2�v�K�l� �E�7�<��>�g��.��v~��?�0q�H0��no��~x/-�#��+PO�9��Φ1�~B�S�Gh�����V�%T�H5k�}����Ǖ������'����G�a:��1����U�e kB6r���G%0�r�߇-�0:`�ys�����5�T��K�B�e��;6ν����3J?i]NJU�v`hX��]"{S.l�}[�+l�œu1�kP^x��vL:�ѳ\%��<"���M;,����tWr�)T+˿��1g�v��D(�'t7UBQ�J���k"�s�k��I]P梾P��F��=�;���S��l�Ӛ5���%r����V�Kp���,Aq�dwC5ٞu���B�!����sR�F�A�ŕ3_s���784G抩��iK������""6"������*_KH�&�χ���#�&E���(���`�Ge�{�HTGn�XR�m�Z���o�,Q2��	�~o�`@����