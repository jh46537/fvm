��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@���C�X��?�d{w]��T�-����0D+�Ot0��>pG�Y�����R�Y~xoK�~:Z�CF�7�y�9x�r��SY����12�so�{��Gtn��<�<�9������Bk�BB�?�9Q�l��I�G��B��S�l�j�_i_��;�S9����oQ���xӼ?�� 0�׭G`\\��i�V�.�m����MLi%|�u�D�߁�YWT} ���Ad��={bW>��9��Dx��a�g�9�����?z���{^+?�	tI�Y�S�zk+Ib��D+��S�m���R�>	�U"c�-�b��*��w�ȸ�d79i���K[`�h��.3�mc�H�����u|�q��׶�Jb"��`��pY,,nxhHFh�cႍey@Q�D.�~m��r]D������x��e�-���ui��������}eF�v�_\,��č�n_����;>�Mq�z))����<4��$�: {)f�F��|��h�m���/�,��/���R>/���9��]���a: ksvuu>��: 
��C�f��\O��t%�:a�{���Ūԩ��б��Q�_��t��^LB+���f��2��3�>�#�/� %�� �F0��JPB�$
�a-y��l���ɻ	�B�P��]����&���-s��!���v��^�+%��j��r�Ool5=� �(~��!maЧ�3���g�E�6�{�:�tT��H�8wFSÙ��҈z���	��e��b�x�5T��0q��r?�i5-9�^䃟��7m!`��o :���Ap���~�WW����v��O�:3�`iw�?���/�0<p,��p�g�l֡;/���G�@Gx�
S��Ċ\D�7�\z������(ϛ�v�H�%\2�'A#�Z�:g�����ʳ��u�A�Ivc�n�L�#��J����t�}ۄrTxW�Pa�D����H�Nlj��$A�T�ښ��n%�j�u�+/h���A���^�a9{֍�i�����/v�V���B-`F�d�⶗P
�͍f�Y
�Rq���u��& 2ָ��R�K/�2@cs���e��`Ǵ�f6�z���;��%V{#�Fw:��>�⧋��`�Բ�G�ǒ[):��n��Ay�1�r���r^�p%�D@�K��z�����
�0�#����.;%��$|u�a�G+Wxj��i-��Й.�X�g��!��-�1V�S����4h��c�q�~�2otE`�g�����R^5��cUb#l��K�	u ��!R̖��Mwf�YU7ǹ��nP5U՞��y�����3:to;(��7t�vW�/�]���5�\|)��s	r��o�ZV�')� ������V[C����3�ޅX�S"�{n䚻j��pw;Gf�t3t��ʹ=Ut�\��v���y��;���fP�&T�k%�smP��C3Ku����Bq�n��?硭*W���˶���;�9F��~��$[����z���`
S��eR<%��C��Y���ٴ
����4��kt���74��0J����k]�%>�
�Щ��J��N�{�#���+Q]�dV�7�b$�p��as���� G`VV�j��{;3�n���?ވ��jz�.���2�~;����R8c`V-�S�����ߗ����OV�P̷S�K1sr���x�0�F���Yס��hǹ�3�G���M�1���]թU�)��$�p��55�Fv �
����`���&���� *n�^����Jj���:y�K�qe=-�<�����*]��Sz�!��� �������M)�#U�Z�C�x׺�⻄o�e�;���K��O҆g)�uN۫/)�U��J%	ϯY����f��[+]̉I/"n���j��t�i�(�ɡq��q�2$.[7��?�@اԈe��k�p����p��4*�~#U�K� �^�ڵw�
�>hl�{����/W��if����9�.�[>��`'�q����X�:�e��t�F�7�4������P`��������B�3��mx�����p��
a�e�*��cw�BGB��tu�Ǝgw4��pO�I�i�:\���O��\�|h1�+?}��ѹ�)d��k����qa=)�q,�5���h�����0�DlɗF�����s�mh(�\{��K��