��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbM�'���x�|��2.�*94�0�$_ �<��У���Y��L�ȧ�-�s�x�w����_��<����f�>�P�ZnC'��(��􂣸Ղ�3���rJ%�d����p(�v�Bg7_���Ir=���XQ����m�!m�mi��@eo&m��W��� ��ݟaƼ@f��S����d!\
�G�7�9yx�e��]��'���LM�O!�����0�w*�[a�m�L�,֫*�c��pT�Y�]�dp�����4�Ju)D]�=�~��A$�
>�X1�۵(��#��P��}i�-��a�2Q6�$��N9���nLx��`X���M�G��7�}�Ź=�����1��=J�ݲ���C@�uN1¦q�6�_@<��l5<���G���[��gH���/�Q�m���#
�lmA5�p/�v�����2����/��_�t�7/��R�W�zG� ʄQ���4��-y:�կ���4��3E��W�6 ����Υ�?>�R4�zJ�з"��\�Y(^6׿�) vZG��x#RO &��U͙w��7��IA���-�l��۝�n衽��e�O�8�/�.3���&�-��w�i� �܃iB�N��<��@�O���T�
�X3Z1z�#-�i���DMP�c������%�e�+�����=t��o(�pi������/�KY꽩��z�.����w���s°��d��%�
x�WXB"8��V�#�\�n�j����{層b�7&�h��R���<��߲R%9��U஘ge2LP��"��d�g�M�ft�d� y�w
��c22*����M���o½�,���x�A��SI|ę���95�3�)�6�SV^����V�a��ނ�#���v�h�Y�ūΞ�5r� �a��~ɹo tv��rL��������o����?{�O��> ���q@@��ூ���s�#�+�?��;�c_%���Tt��ƚU�����D�)�mn�;��U�KA�$o�0�����3_.�o�iT�1��ov\�n�H�5{�n�H |vȢJ�����)��NO�&+��,��7��؉�T͐��Tu�T� +���[:��IPP`���L�R�L���6����A�s�C��U4K�Bǧet��%�Pq�#)�Ek�d�Nr�#b.�����ixb�@��D�m�J��'�9�����}+�����x^>�X�.�{�"W��ߎ�O�B11���	�Uf��7rs��urM�ԟU��U�>��H����|�Mm���7i�3]��[��S��V�.�w��^�WE������@7d�Lht^�s8�"�(%��L���	�ƒ�h!�	
��)�_��?�Q5	���WԒ	K	n�侟o���75���n$������g�9��]6����~�;r\�;�v��U���Xs��}v�"�F<�$i=�bOP�X%VaQL��|���\�Y��+}�����#�3�VId���K��$q��7nY�42.<���m��p�]�9�&��L�<�]�����8[+��m�a
�8'�P�ǠE�4��&�+�`�R�Ȍ�U�����-�J��k�
��
�����g9>�3n|�Ti��c�ϙ���gl���`��f>j������ ���g�h��N���ڐ*0�������d��V�1ПD��jы�kؘ񁙈����X/�Ɛ�eet_V��fA� ���- %�A��d���}^�I����D�$���c��'ǽc��k�$	x'��4��i֮���K�BVmj^��f�muM�&W#I%�@�Nw��Qk� �;�+������$���64���S}�i���W������N�6=p�hli�5�N���#(t<���,�9|99�z��Dz�ާ�`'�6�ⲣk�s��u�6R@[n��u{h���h�j������kf�C��;N���L��[�^�di|v�ב鐴4X�t[��L$�ѝ�����!ބi�⬿��	G������J	���� ?X}i>��X�(�Lv�~��' ���`��Iu�mS.��]�<�zUd��m/g,aO)Z�ІT���%i������)+�+�'pG��f�
�`5&�b�:Uu�O���}�(⎰��i&�O1�@e$��u�'��啛8��"k��Jۉ)���2n4�1��f��Te���@S[�yF�
��^��BM|L����M�b6 �s:��m/���*��Np�׹�d�/���D�|Xx(�;�Z��u�:=��,O =�јo�a��}�=G�Zv��&��5:��z<��zM���ɓ�&��w_7B]ԇ����Lz����dVL��X� ��gY_򅜾 \\|!e5pM<	��c�;A?9�`�D�����XE�܇u�_�v"���<���D�� ��Ǡ=޹F茁�����݄s\���h���k�e���N_	�⑇�u�}�ؤǝj#�����u��7���,�\�?_p��km��
��l���펲��q��q���M�����iW��Q �{�%��<h�I��x�;jFC�i�Uj�-�.�S�T7�n�d��&�i�PI�\u��2�~��T�������4����[�s���?!�4��{�Jxk�6w3�����5�"�W����0�z�P)�hR8�\�~��,�MQVɑh�Z�o�Vxј$%��Y
+�9z"�"&V���@�~h��`��s�J�E0WlD�"K ܝn;��Z�����jJel^Ғ�X�o�*��[bJGڤ��5�5���V���~� �b����P���O1F�� bT�t��S�6L�t�IE(,��u�ЋwG�Υ�/�|�99��h!:��o�l��8����[��0������v�ƥ�t������"k�*"��s���J��IA��T}ڵ\C��8�I����r_��ײq��	�g,^n��Aۘ����r��N����a�N����7�t:[&@�b���!�q���ċ�,������/��2::?����H�ݢ+LL�8� ��厜�Z.�(�T�e�b�kx� �F���o��)�
Y6r����D�a�&B�YI�N``|��f�m���=�7�f��m�y����Oq��=�%���u�ד�(R|{Ke#�����	jVlD;�b,@������_v{41����4c��6����n���l���C��޼Mk��jlD�''�̯�g-}��r��*E%��}�xgah��^� �)x�Z�ҕ������@&��iU�}-!�>�}�<P�"�P�&T�d�Fm�렦!�R]$��bh�-���5����ǅ�B%FK � � �3[
Ӹ�!���k�x�~�sO����m�j�pZS��B[>-�����UW�<M�������S �{�]D[�:�%%��|�<:���~ǐ'�6}��?��a�o����1�x^;��M��H�C���lfp�Ѵ��m�y�o���ű0�l�a̴��)���;}�߈����J{�n�'9"o����|-1����YC
���:�Y�@^�6�{��6S���Xn���~D��:�J�D7q o�P�Q����n)�>�H;�oW�p6W��]�N�,��� ]D�Vm�X����.-�t\��o����T��1z�_�k�uD|d�H7é�;��-Sᨊp��>)a�l昏禯v�q���\��E��_���`g����0��!���r�5�4��4L 2�t;��1��~6�-�;G*ڻ�1�Bل�һ^gy�a?�WJ����c�#DD�R�l(<�=[D[u��$b��J�
���HQn5�\;�~�g�Y0!�uP	������I6�;:���<C*<��?�vmg�*���eg�;pvAP�vs����g�!��OIZPL�H!����Zy��E������X<E1���4t���d�~t��w*�l���f$��E��;$S���=@]��TF@Z��#�ej�6׷�},�P͇�z�7��~�I&�k�:�,��sE`���>� �T�v�J��
0�X���[�VBM2��[��?�2��hGT��W>����jE7�ͥ�ƵVv��������o�����<a|tK�*����MX���bD��y'�/m���-4p�SUF୾�F���X9s�寘�'��v��L�o��p}Y�!����\|�[�{!'���T��7��^X���>�Q?%<W"�U������{���s=����l���5��s�-{�Uyv�*>,C���UE�B��)D�y�-�sTN�7����ZU���ԛ��4�!���ë��� ��T��ÂKt����:m-��+��x�:d)��F�4��~XYhV~�,0Bm���U��i�k�[��N�Va?D�Й��O~:-k�
c���-/����ɩv�u͓�,�~�N�~O�$5��3��x�(>F��^�Y@[#��3���Jf ����;29�c$��M�����Q�Ӊ�=����Gb�$�6�*���/�ݢv��0�"@��C��ʩ.���ǆ��q�i��8\�� 5Ti�m�q�Or�E� ��~\�*�O��`����pϡ�KR��P_^�o�8��=�VG�����kQ�^�5�+3Nj=�]O����J���Q�ݳ��w���A�&> ��3L�+^�ͪX+����j�6�F6�@g��h\��P���Ch�]9U��z��-�� f_��Tc�-����_���y_�/���2�ْ�����w�����A̼�Θ.�1������g@���O��rT�j�ċ4?]����7���ܲx�(`����H*"�q1�u���~Y�*�K�:�S�l�H1%�΢��.dw� �~n�i9�/a��o�3d<MΓi�S��-pɫ�W 2�Z�AV Ze�T�7�y��3O<��+|/�Q���KG)���`� 4����3K�^�T\kCr��"nʒ,n�31������:�L���@�.����τ�zK珂]9'�qK�Q{�x�a��h4�v����x���GY���+�R-���&�c��������]s�W��) ��!Y`���9�eH���j#��A�T�IcG�ֱ�6!�"�S��S���^��V�Ul/�]$��~Q���3����q�}���6�Q8K�ٵ7�H'u�v�P�(��O�P��Ӧ�Mxl2��a���󃼏��h��E�Y{�h�޺�t�պ�����3o��WT|T ��������ZA��C[NT}��@�[-�*�
�-���01�2�0Or.����E����pP���&�۬m~~��P�F�3沺��"bb�ݼ��!p�CNl0��͐k�u�O(��F#��F��cx%-C��	�m�2��CKM������+!���a���yv[�n���^I�#K ��n� uMe�S[m�ě���ǰc�a/���^ ��rX�]9�<���d�8'�]� ��;�z�H :�Y:�Q��4��A�8�p������{"DQ�8�}���z) ~�rOPLdR���Vw*�	��HGT�4qK�G�I%y}��]��&)#�t�T��.��[���mV��o���[�Z�����+A��|8j���j"��n�u�l,湑����b`X*��g&������lWbm��j��i�P��o��?�:��m4S�.��o=6-�_�m@��o�4��5��Ik{H�@:�7zto��:>�5�@��7��%�g���c�	 «X��Ou� %��8yL��TatΉ_C�H�����:E������Gn/�Y��^0��bbiG[��0�Sx��f�)������d�ߊ5�L�T������z� �^Ϧ{=90��}���Z�}����'�Q���t���cv�4�J��Mߔ��½`:�y��
�N9p��Zk����e�_:)�}kZ�0�(bj#����!D41�������r�`�hɜ��-e���b�n/⏕��2�����Gkװ��J>?���S{��C��	��0�'s�Z]mrfe��5.I�~�Ի�u���=]lX�fe	<	��Yᰦ<B3�ƥ�� H�����+�Q�m�,t��#�Ts�����p�߭�����閤��Fiد�@���l,�#B1�$r�i&手�1&�2���7H�G�1���!��,�N�o�,��#��e ��q��r�Ƈyj���I}M�\�N>8~� �nt��>\� Ć3}�h�!3�j2A~��>�߇�S�RU�Zvŉ�U�R��K���T��|o�:�P�Բ�J�P��+=61+�N�*���0����ߔ�Y͹���*���W�C1�[p�n;��[@������Ѓ�	���8�����{K�a���-^T�2�+T� sɫ�1��ֿLFY�iYf͈Vt��ts p���k��x���Wh/J�X�TuL��-����9����?]w״�I�����e���k,�OݳcT��Mp�6D �+�as������T:�ɞ誳�-���8�l1%�R�\H\�N_=�sp�p�]<:��Y-����(��S.��=V>7�<��-�b(o���ڬ�]}W�f�n���A�U��܌��7�le�~�]>����V$�����x�Ԥ��8�����V
_������1��(��_���H��ȗ���9-�h[�*;=	^
�=UV]V���=��ոJ��BZݗJ���UI�D
Sj��_55oh�A_����Hc��V�s6�ei9eMcE�K(x�C(�>��������2�c�Sy���sO�@��m�s����Oڋ{kB�� �YZF���7z*��䰳w���i����'�~�t�\�``�2�š@%��J� ���>GD��Ah��h?����6�5�?�axG{�ƣ�j�y�vGbôE.R$���F�������<C���l��Dv�[5��јf1�gǻ�s<3���a���7Q�1ĭ�J'�9�^Y��h��k��0q����]��w��o����AIz��Iǣ��%ixy{�N��I��>��]�ɣ��P�/��1,/n�	U�6U��9Ш}��E�����'6��K9�k�ϣq�`^׼b���OMa��s�#!3NQ�Թ@|�Cy�0������ۗrx[�p\�я���e ���i\�q�A�`�"��~F��
��h����5_�xY� x����]_��\���C�8�&���.
RB�9(��[���8��n<�a`I'rLFy
�]���\ueO]VO�g��L(�`���'Jao�� ��h�=>K�P�ޤcj�c@�[����,V��]'�<>|���j�E�j���Rllݘ�i4n���ޞ}��I�z$�w��:k7�no#&�#>����y;��ݽ ��mM��x��}2]���;:w�?)���w�aeJX�?��#y�&�M��Y9�����\4�(`���ИW��է:�+;�_�av���gF/J^|�!�+�1���i�A�c��Q"ǜS������;����Y�� #�N=��?Y̈́�I�)�ЯP[c�щ����A����-_�Y���|M��X���'�%ܪ�k$(L�I�jJ�tn��T��}����
s�+~��y@{�**S��;[�<�k�>(3�]HN�����SF @��Y��vH��Z������	����Ӱe�iVxE�m���aͅjS׆u����U����C�h�g�������vkd-�_ 2 q��OE8"��kW��("�[�"�T��U����޶?<��2�����U�,P�K�ϩ�5��Ԭ�x }�{� U�~�L�6�F���4�R�+C�N�'�A,!j���d���|I�������K�괈���������ӺW������a@�n�VRE���M�3��x�]����Z*�^��ڪ�)�K	ͽ�L	'�
LCw5�ɿ���P�S�-R���xA|����\R����[�۱>��#�:o Waq7ˎaR�t5)N�{��␀
����/!zG۳oQ���O~9�GJĥp���99�� p��ӢW�����F�kį�Kp��][I��4�go=o��:�Xϻ�=�P��k5���r畟n�\_��n��_S�#��a��ט����>;�m�W8��hu���������J�ɳ��1g�$rs�R'��ȝ}U]re7�g:��ۙ^�q��q���+�Q�l�J7	�	F��w_P�#< �3Б�^�A�mJ�Q���������!�d�
+�sʇ�s�_eŲ_Y T}s2qB�nְ�Ǵ!��S3Ʉ!@.#lq������p���Cp�/��^l�����{�VZ���k1�%Jί� �<�����/鼐��LNXO6ß�=i�\Ar�{���l��e����ڑ�h"�Qq9}ưإ̻�D��NF���\*�)�f�@���(|�"o�Tr+4�;rM�d.���[>8 ]������U��G~v�Y�# QZ���֦I��&���`&��&߿V���
���g�/*�N{�ڼ)Z���ِ����:��\ƆDO�*��|�-dǯo-��^J��J�?i1���g��2��E|�~)��\&ф��Yg�:X��v�-����2��Xx͹Y��%��J$��_����1ne}q�O�̲aNxs ̕ST
l7=�0}���z{&�# y���9�У��!� *{~�M t��I��!8ظTv�����Љ1+���]��3C0AL)f��0�|���'S:�e�V�yA3�����F��W���1�"�d_$���^�H�����,Fp'nvQ��Ʃ��)B�1���k�i?��e�E��b��]�%A�0i����+���}P��|�����S�D�&\�(%�{�n�R餙��{1=B.d����@��������Bq�L���1�D{@O���v���AGx�?���g/;i�i�ք
�g|���p*v���	�E��Q'������^�r�胋	��蠄3#���f7'ִ:���;#M�����xa9� �XNTmR]�s)�v"r=σup���#&�t[d�X�?�H�.�瘹$���rshfҕ��5P�Õ�������/	�MS���b��	3��Ƣ�lm,q=���"u��5C�~���=<�o�N X]]܈��lȘ�c�|W�����O/���gN�(k����)�S���PH��j��#��d:m�S뙼�(�]7%�`G��V�t��~~�]��Y]m����P�Q~�ˤ�g��ؗd/�w0�ŬS����0~���3�`P��!'�emY�?�fl������8<�*Q4܀�ɒ�HLT'�4sXriEVHJ�W�.�T'�C@�=���@B��	��ɐxRs_���^�Ȗֱ��G[��l�(~y䆐�-�t�I��J���Ŋ_�yoO_XY�������c��;��ZQ.ɦ#\��O�92j~��t2��f-u�h�/�J�G�U@v���%��]��O�N�2SZ|�+U���?�"����(``�_�_|�R+���d��K��0�wO�rT��,J�n���"��0)�D9��j<��ޑq�G���ԸS8d�B�X��{��f?Z+���!D�)�Cl�j�Z{𛺒k�#U3I�]55�àd����f+~q~i~Un�0������0�_?ד䲲����`بi�!X��S��IX�SM�Np0���?�%'Nk��<}��"�[9%��u�!�BL;V0��t9N�sO�^*�Y����7Y|��;:i觡�!�NF���S�&S��U���!m��?�����X�'1�����5�\I\�tE^'�!�?�&�c�!�,�a��;�<�;D�x���G���#��p�g��ڸ ��0�RW�>���E�u��8�[֠Bg�A�;�Z��Y�vLw�*(���%����Į<$&���=A�<q ��xksv�����o�~�я��zZD�$v�	�űB�VT{��㉓D�:�u�~�o��ӈv	��0^ȹg�I�p`TюUk��յ.�������9�K�	݆)��❿(�k�j���t���Q8{��#��p� 1�.�莊��������`pD�V���vd�z��ʃx��߃��3��1���+az�A<�W���6�\/p��N�zVWb0U�hX��q	@���#ς�H����!���G����?"�]7Y8���� 6�Q�r8!a[Fl.���A��J�{�"{��2/�q�K��%�ʄn;����'"<X�C�|���C5��� 9��ϭѹ��[!.˸�J�fS�9&��n�I\m{�ږ��-t���Հ�!x8)X�����x��?�a��4�,��.�T�mk��.��]J(�ԣ�TC���#���oD��q�}X��vuXO�2,�`���W�$�ϳ6�օ8�j�JR���qo�� ��mmb:�<����R���s��U����D3����h��A���fZ6{=�KWL�D�+L�O�����r��L՚ֻ�p�,\EJ�6��4i}��c�g�*�2�?��xo��f���9a����72gLz�SqV��$YK'$�[���@�FT+n~>
5�������/���I� 0�G�笶c����I��P��!�I%`avy$� ���6��et�9���\_/9�<�$���UF���;M���=I��_j��+����/ �g��g2�?��2?b������fM9�S�ϻP�>at8��M�0�7�O�ʔ�X��ܘX ��C�T_X�͠ڠ}���(�PŇ�ܓ�� O�<U�%BU�i�A���H�$�݅i+�!�p]J��3���t��>$���C��\u�v� �<X�և�a#��^K�>���h/��1�������KlY�,~��EA[�M�ƕ�X��H@��г�Zu��`�]>�����0�2'k�u7�����fn1T�#�������~9�A�f�����aX��������^�L�� ��y�{>�u�S҄S+A��b�my��Po��F.;4�T���d�>��)B�Z�`�紽
Z�9#�,�ҠZ{N��ϛb��y�����оS[�D��.�Z�w_��\����A؍;��&IP��6���݂��wa.}h�
�p�b$ v�H�11,�M	=����d8G�[�@ɞxb�����	u,�4Y4�y3����L_��#l⥃�U��K��Kow�{p�v�l�۶�Q��{��y�E��������-e�'1*�R�9"�|A��N�`�%#��:�����}w�ņ?~�,8�j@�%�,�N���r���Xn�_���� \~�V� P��~���B� ��%d݄�:ηmJ����[�NNu�.���'F���+$U���p�RGv����E��,z�5����VRj��}�r��)���>��x����LG�3b!u$��w�|�e����^@�O���ʝ'�~LW7Y��a�XYʹ�~M4�x3���7��(�7Fدm`����sL>t��<��>Z�սBۃ�<���,q�̛�m�H��| �_
�qo3����~L0%[�T�	繹��eD��$�j��kI��d� ~d��k
,�!���?��"ڒ�o�޶�\�D7n|�z;4�����7��|>uTy�R�a�	��0����]$M��������B�������=y^U5��L�S�?������&R����,��}��}\�Ɯ�@�g�T�������~돴3�T�kE�����?
���<�dXAr��`=O�Q=aV* �RbvF]`	K�)��y��[O�T��GO�{�g�x��m�����%"q�� ��\0Y}�&��o��o"�Ƒ�<��W�_�º�]*���ߺi��+�2�B{W�sP�V1��Ú:!;g{`���	�oN��rQ�[�X*aE+�wC�����H�<�{�_e��p���G�{�C!��;��3����
&�O��.�0p�>4+x��@Px(>ͳ�M�ɢ ��tr(�*�a�n��4���R�e�ͥW���cl��iY�:��qP�j�T4A<F��Ƶ�f�+��j�j
�p}�c�������|�/����_RvحmD�<d$���\/K���)��`��6	�(��`|���b4nG؝��m��aK��֑ƥ�4��T}w�N��`��Lڃ\cSE����z��P@���9��lR%`q�ΛY������sONk-
��k�pP��#�~�����n�j
®��tS~�y��	������\��ʘ��ȡ��rx�\t�4v�Ȝ�#$Gtછ. ̂��|]jE<�G��-9��6�$}d�T#�G�*�!&3�?�'r5�c�
�R�g�%��X�1b Ν��k>"�-��3�ٻ�K�w3/�=� ZS�{��z��ZT|e��
V�X�̳xEȔ>���l%�ĔB_�����N<;P����#�%��C�����>��iI�ێ�}-j; �f gz��Fk�V�qi�mE�*�;�J�)7HѢ�M�����h����0������:Ö@s�\��u��T��36U�싊����'�)׈�O�Q8-�E�/A�� a�@�+�2�`�=�gq+=�z��^��g�<8��]��f�{�+���d��蠶y"7�,�VMB9��H����,/�%x����7ӺM��~L�� �"c[>����2�']���v`��C%�9��G�\�9�o��D� �-*�����L�\d�{���iێ��E�	*E��v�b/��2���cTx� ă�H�݅2����w�� �_7\����0�P���'O칐!�����z�nr���	h�~~�o"��T�k�@2�ʑk�ZO�g9��*�<�N@�pD�RPTr����W���lH�{�ɢn��g�����T��f����b_oY	QN=��� �Y-�_�����Qt�W�1
Mp�F=:e��:��2�6��ծx�30n�d�"�t*�'.��?Sj�`����z.��!�Д�N��9K��Lr ����^W�C��=���gdU�9�I�u7i���;D!�ɄN@ �m{2
��:"���*Ou1�)��}�Ywamx����>K4�-b ����K���@�O�<f�������vU�u��Q�"O�.V���$�e��a0#�S��،��H�V@_�@ˬ9a�Z.�S���/��0(bŧ4��L�A�E;���"��;y��:����*��H�C�p�+v����CI.l����ǒ��O4]p��fJ�%��ݜ����]I�,Ό;�^��U(�k�"��'��ɚ�&�>@��
�;�i��HT��H��	�lo���x4��=�i(��8�@�I\F�qǪrAɡ#�Nr��e�k�"�Ш��d���	�}jM�/��=˥������r�S�؋W3v���cڋ���E��(�7�2�|��B�&�`Q�,�����*� ���W~(;�?2����rC�3�U��@�[�]S�+|L����V��Ь6Q�7�:��7U�����±���@��GW��C�|�jZ�tF����5�GO����c�� ��?r�R�l�/W�}F���{�D�������u��##BA��F���p2[ڼ^k��aY����љ�wrƥ�m�S��;7�>i3����ո,�5�0�ŝy����g�߸ci���������#/�1�ci��{�/�&�#�� �9��6���27x�D�@���qNC��C� ��j����و����:T�tc2�m�=ٟ
Yj������ɰa#��{R'�@o)J�K�W�l�L���Ӹ$�Eǎ�,~�M�)��_�O��M>PQq��>t�n�D)��w��dE��g�U(����yJJ�Ϛ�ei��W�}lЌٍ����wx`�xyX��G�G�Q�
��@YGj::�sb%�#�SΛ���)��N�QAM���s=�;\8!v��H8iX5Λ% xDY����:���ѯ%bH[���h��L����_FF��)6Y������l��v�6ۂ[dQ�3w�[2|7M��2�J@_���IW�0}����!(
���;��o|����Hp0���w0E�qR�:�X�y���U�@e:������F/{���K��og�@��W<�� Wsx��ԥ%$LN&��$������z����L?ڠb�1�ˣ���-����<Ri��q#�)Z�����͊@�uQ��D8lyia|e�|b�r|%���nH�����h��5[65�������]����Q���Ka�I.<0�����3�"~1�|í��H2㼫
�c�Ds�-x\i�9̾k��<��v�+�	!��}������O�����a�K��ў�����@5�J4�����R�8�I�K���b$�P���6qr��=��@�����4��<�{���1���K&Zߧ���V�7�)3���u�z�O� 5�J���v(7��EZ;��H���eu����@(.e��W/@�I<@�V��X�^����k M��JFW��׾�1�vc,rj3��?wOJJ��0�F�3���r�*|��_���3c���
�G�u��mOb����-U����V�,o�K����SJ͂˧ؿt�U�Sv7vD|���p��l�s��'���z�]�%+���?�b5���?Q�o��{���R�t�*8F�\ރ�꽎�_�td ���A�0�����(h
�����|�K�埤l�҆#�,]�X0s<���$ ��:�x4.����x�BD�c��2����F�P�IHؼޓ�/bso�7B1���|�!��#Z 4�L�E�Y��9
�Ik�d���­��\�Hlf���Ѷ�s�N�����H�e�YDvG��VY��'�_/ �-�cmݱ�,1���/�6$��^��u��pF(�?�h���8�C�Bh�� 
~״G]�/���G�oW�&��7��$f�B��U��?���c�dݣ�-K���qk�J_�t��/��3����w�$ɦ������"%ڧO����偬r�bϟ�A�9@��nK}n��g����ˋ�Uȱ���*����ͦ���v�� }4`���|�&���ГQ��{6�X@�Nv���!�]e��o�N',���Ti��C�S����}�`鬎;.���v