��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cqL �$��)����s��`���O{�N	���ˢK=�% 	'�R�j0�z?kP���N���9XvS�J/|/��6�̫��Hi^��:�#�0$(��U�P,w2F�Kg�?"���:w~A)�>�'r�Rm<;����at� R�Xv���]CqzꙔ�"���\^�����!6:&����u۔���,qI:�kog��m�u�˃� 8�$NN�I4Ы )�0�V:l~=k�H�[Li��ı}�_�R�7щ����s"���B��~������K�~�1�ϖHIy�o�3�fX�>��i#�m�\A��y���^����
�Su��5��^wT몍J�]h�3\�\'�N����c݌G��FQ1��>��|B��m	&@�ޫ�d�J/m�*uQЗϫ<���8�x D/eJ�����X2xϭpq?"u�7+Iy�O}[H��p��k矽5�w7���<O�-EUj����os�5g՗��A�(9��|����-{�՞N�dc��p�����@yF���+7�H�ي�+V���J�d�,V�"x��zs�Ju�`v7PO���aԐb�����l�o��n��~�Ď�0�	x�'0�*S_�he �Ҩo�/�6GQ7V8�h�e�ptm�d�O�6GbŊ-t�t���D�TT�ݸ��a0��#E=KF%}���&ky�`z�eI@4�s��m�|�T ��Y�37�k��K8����Z4���d���¹w>�Y�ܘ��y�i_�f�!N^0K�qA(�%�\יS ��'�Q �q�Z���bq�~�'���Ca���Uq�8���>n���ى��������l~�-<�bgxS�?_�=���z�I�8H.G�6�bD�e4˹_;�^J��)�%��כ��	ad�׭0
dt���YN���졩�hк3�x�bq��߲�����n���|st{$2�'��m�ϙ'���<n������QքQ
��3f�衾����`�\�feY�E�qWt��>Q1�Sue"JԆ?��o��e�njȨd��N/˛!�1P��R����K>R2ckب�]�<E]W��]���;�R��F��L�"0�&�t�Ms�Zi
p��.VN4t����i"[h�C*<��X��G�����w���jo�;M�!5 �?Op(Fw��NOc_�uc[���L 	Vyz)�\5a��;I��m�u�9����\&�Y�B�e�oR �8Rf�������,��l�]�:eKQ�y$����~̸���P�hc΅�=pkeA��O�ӵ�N���c���Y@Y��J ���ɾp�i�����gL� C�t�f�*/�cl�n	��&f���o;i�w�ǈ�J�������5�$�I�r�+��:��{�L"~QA/Q���\��d�&��b�	���}����Y�O}F_�|KE�Wq��?숂�%/|�M���ӗ�
+Y�ec28vj�c�W�{�t�Ynt�K}�B�Q��xM#5�6�J0H�$fa��������oTN��ɼ�/9������3�[�z�ף���s�����.����H��y�fL��L�������Z���-I��z�p����	����8�W(�Ei�	x挶�U�<$:?7v�E� P;��)r��m�c��a.2*\�{�ժɫ����S�Np�A'���H��i��aJ�")W�������D���`���v�r��?����#�Th7Q�\��T��6E-�=}�VsP�[�Pʱw�$��hʕ�������:�a�%��CC��Q���*�_�4o=�[��*π�,3e����ｶIk���o��y����=�M�Io2ik�Â�`5���1���7���/����U �?��q�Hp~���p[�R�؜6����7I��z]�4����l���������܊Rt�>�& ���Q���
,�mS�]�,�����Y�[w�j�i�+�e֬ᓬa���7'P�3��ц�!��>DB�����U-cY��h|w2�.�`�T���a�#�T��*�Uy�1[�h=4���jR��T�8�[	޾�asz�k{���-*o�aK�4F�X+�#7� P�<Z�7�0�0�?�-[[�p��j���HrL-��B�V���H�ՌT���?�(�p��ီn`�LxE}��N��"���7��Ie�;R���5��X����ݪ��)$p�C�����h�Ϲ�����F�~j{z�v^X�>d3Q��2{�X(�Elw�M��y;0l"�lKV�hU�-��������!�,_{�Xk\ʂ�A��I����ʑgڕE�0��
��.x"J\gl+�����q�27�[�yǫ0�z��L����t����[��W=d&Aש���}���c@���*��v~�R��AB����fPs��1�"?t�J��
}3t�
�X�\^Y�8�O���>/�x"�_�璨�B�~%�bcP��r��9�+3?�1Gwm��j����Q[Yc�? ��bS��h��ʪӫ<H��+� �~F�֧�o�5`��`Pq�\��9V%Na�E=�6����#oףS�EfM>PǠ
�ap�GdǼC� �������r�}��l�}�'����K�8�c�b��4�zr���Sf��ؔ /*f*�&���C,��^Mw� �(��-.��ؘ.�h�h6@)��4�>^�w�N��C�/e�)S�\�aJC��ځ:���=_���f�E1t��� ��z�U������mO��ݠ�7��#?S�d˯�4S}U�NAJk'H�"�I&_YR�29�&���P���'��
6]C�sgx�~R������aA��փ�fr�.]��`ۥ�~C���^u�<�Av4���>)pث��f �j�a{a�l	���~���r@�1Nm�7å)��a����ӄ�zԅ�D�|.X�e.�\o�=�h�h��x��׽�bZ��߬T���Q��1�´(�Kn�� �,�=tm!��I���
=')[;���^��ωɯ���M�:�=2-�R��v�r���@��ND
U~qlSE~����v��"�Z�����x��:��`�����d>%p�B"CX>�a��E�u�
V�l�>�@K��J�z��1�kO�H�P�&���/�q�ѝZ翴|_��Ӡf��\�{��7�q��30Y�(I�M$�2�� �����{�w �����5V+(����O�P!k���c!53
Q�e~�߂.��;/��D����Ƌ��Erˏ�d�7�Ѭ_�f���mdԻ1�IzM�:�[��H%&/��r����#GK���5�ղ���-�k�I|�%/ۛJ��855P��Ha&R1��e�!:���}�H��q0�@(լyZG���Z���)��Ѻ���4KS�|ua�+lˇأ���c�.C0�>��������!<�����pO�A�y���96��,��J����f49 hW����&�nK��ċ�q��#�VZ���;�>����F��=tT�DA�I��hy������lF%�X���E4z:˗o��ɋ�̍��<�s���Ҷ���=�"�����ϙW-=��$i!N��,�2��&���Y�L�T�qc?X�`�$R�i��q6�^�����p�=>���s����OaCM�7<V�)�)�+�H��Q�'#�M�i� ����D����dDm�"�,i��ly��p�Ӻ r��o������#����~.�O�������yµ���+��!���������8c��
�O�ѵ/��g�����B�c��
��������Ԋ-C2? �96d�!��1�G��S=,��.���D�uk!}�����ށ�F?i�/�ʏ��9֠������Q�����W)��YRIiɞ���'�l&Y�������g<>p��Zf��ըif�0r��9�R��-6� 7��V�;F6����5䀲�ЇW�p��"�#f��,&�2qN3V��Q��R'4Ǧ��(y�$�Ƶ&Q�{c�$ڳ����G�t]�qQ~��﷼���z���<��^²w��"��zp������;">��1+��
w(��!/�l���A��<���s!�(2f1� �1��d��x�^�e�u������	��O+O�8�]�Cx��0ɮ���M|+Y&`���ÝvŽ�Q[;��._�4�&���b
�,�ꋯ�;�o��z����h��g�c�%�v��,�%6�i5+�Nk�.���I��\D4���dzy%�62�g��T&!�"a�&�/�����Ka*.0������'c�~��H��|�klL����ħ~�� \Y�4#-��	a\f�v�;�=�r��E�[ݒ������.|��Q2<���p=�z)&}C��[I��!�-[�GXk���,& s�D�X3�@�H�Oȴ���H�zwp��[8�c��F���p����F���2�H,q.m		ż���P�7��KK�:�ya�𧼣M��x��o���IK �M8���N{*�~��ܢ���{��s	,
T8��ގc~2e9�m���S�Քf��wEZó�f��=<��+���/��V̽����[Q4tv'�q�d��;���UM�w�oy�'�KsS�u��)���?e+<-�sfן����I�<V�߶R�7ug�\ AL�7F�"���Jj�<�ƽ�_���(43���l6d����cf�b�YBk�kč���`�-,��I� :c��(��!���L��#/�
�Uū��Q#��^n�i7Uv�y�N�(e�R��iK_-�s<s�
� �no�Ġ�d��]����ۚu�`j��.P�R�r�t=.�C2}�0�\�#Va'����~,���r	߅�q��+;M6J��zU�����q
���<å<!�d���h�h	&l�����J�k�u�����$Ru���[P������\Mۦ =�;��p���R_������K�Y4�_�6-��6ڗ������L�2���g"����+���҆����n��}�2QE��z�V�߾��}�