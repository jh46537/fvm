��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8��A��t��
�]W˱�ӆo ĔU�!�!5�S8t�Bu�%����t��������6���%�bK�GR���Kظ ��1G�r����8/�tUvȘE�5�s�;�}J�XQ�0�t�O#^P�����T�)!H�>V�G�����[���ɐcʚ��Y6�1(�	e�aؔ�S�Ǆ�f�42	��Y�q����-��V{�<�vyd�#�NʟQ���v5|��`;��b����`fB�Z�H>�����	�M�a�0E}�>��J.쒯'�v���W��=x?Ra=�A-DG>�|��q6�|l\Y�\�)��h�����CQ:��E��)�f�R:����z�O[��A;�[��6kP�&}���Z�>��:R�U����� y���� Z�J-tl�oQuO8�����;Ẑ�V
������ |4��L7�i'��X6'���?��@}��X�G�Rg�Cw�F߽��e!�_��v1Ne��Q��:j�JmT�:]FB%����{��?@�3�UXi
���D��v�M��I?���@Dn��eʰ�Gn��X�~�ta��R�vBW�npg��{P���^�N��\0�цB:0�w�2줨$3�>�����= �K�a
��,�~���ş�d%Lь�-]�P"=�W�q0�Ѐe۳�l��34]�t��UMWw�~���b���X�k�gm&��`3���^R]�O�_셓�N^���*����jQ=K��-����ڙ^ �A���p��Q�b�����-���&ԅJT@IM��!�ώYr����>Ae1i��M�1���d��yՈ\��x�Z��4 !S��Jl�M,;#�g��/���V����_>��VY�1+���A�*�ڛ7$;�$	�;Z�������{��z��ˍ�R�y�I�Jk$$$��ZӬ���|(T�^
}T���K�Ϳ6W ����߻�������G�P��]Ĳ���6�w�N���H�G.�׉j�;r��c}J{��=*��P1ٵ�Q��ut�%j�2A��s)�G/���Q̾p. ��TYjM���Y��B��_ ��.�5�����Y7����M/Ni���'r�\k�%'q�N��p/a�K�Ҩ��F�O��"��7��7c�n����gy3:�T���Y��w9�]��Q�%�P�ōTa�ӷu�w\����h]f����^�3oFB�U� ��}��,��=���i�%,߲@i�
�� ��YQ�`��_������(�G$����?�ϴ���1hlZy�6�;��I>M��
�3�5ͬ�w��7 �A�+i�*�E�:ѕej��������� �!"�b5���]6���N�i�8��v�L�v-�]���ګ̴-�b^VI���Ϯ,ׯ˞�g)8��(?ꚞ7eR"L;ջz��M��m�v�c�H�ٺ$�SDn�5����7C���$�y��d2�d�e<�5X�H��)���:7݇������(Kެx����z���Hߡ�ݐ�ǦcX�X��J�����d���o,�A��ID�:����	�i���Y�o��� S�vm^B�ǉ�28w�jc�(3�N(�b��a^3����= �M=���o7�$�勡��!X�&�g�(�`'��p&ч,
�K_U6�%����Y�Emg� �F���D�79��`���7{3c__���[P�$̩a6'���܎P�W֥�3ïɬ�1`�Y<{�F+��w˅�M�裬K�G�8�{���#|;͌��7�	YՁz1���Tt8�#�����TR�l+p&?^�+ ��G��.ĩR*�Q�#���`޲s�