��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�;<�T������8�l��s�����X(��R�D�J��`:��e�R�u�~R��u�|�9ڜ����A�t�wS��d
Z~}(�w���S�q��D��/J����6�CCV��'��=����[5���k�
�G�3�O|�HcE�HR��*�9����Z����6�sBP��`Ȫ�����.��네�C���3��i��ju�Dh>�4�QEb쏺H�^��� 1;$�Fƺ:�p�ew+��3�b��QaL�L�}k&l��QDH0Y�/\!�&��P����gd�5>f~ƫ"̛���Ο�0�N(�Y��~D��Ќ̈� 9>@�̡�0�*��3�f̷9�)�9��������K?J�g��d�m�9XT�.�i5��z���]�er�6]�v`O�� o��?Ә�65W:5�D�D
�&�[��Z�X����7{(/��c^�A#X8暻�����8�r��B��sC�"�|3����\R��?Ǧο#�����������s����&�GqQ��t��������	�pn S%6�Ħ�9�U�/�TVa��zF�I�YYj���n�Č�ab�"̅3���7?�X���:,�h��U��4Ǎ�>�7���
q���(�H���C����H�-y�(!_S��`l�_R
*օ�rAA��|�YS�>��>T����蔋Kg�8]��&�K:���l�9k?:/�}d*�dV&!_:�bqu��K�odf���Z�~sF3@}��y�J��?�x ���;c��Ϗ�bя�� _�f�c�$i@sd�^��7��~�GN�
{{W7�ը�-�1��mH�E��T�ɤ�;"�aT{9��LT�@���0���'�	ѳ(�'넕��:4k���2�S'���8���8FU�+�*��E����t�hӒ�dW�xG2�q�� ��:��t%�z�f�	�-6ӵ<��	ו�89S��#)Aʎ=ͪ�L��>��6ا�:��'Y�T�b]�0Σ��04����>W��La{��12�@��Yvq�Q�Sz��٥��n�s�B��x��0+���� �yR��K�|��N]o��/7�w�ū�������l^K�$��)rO��ߥ��8ƭ�\��q�����7�J'a��2:H[5k&6@���ѡbL ~.⼕PU�>��k�xU� ��9����[83 ��z}T'�5�V�>�d�x��"�b̊�9�p-�77LxlG��ߐ�NA�����#:�P�k��KJ���F���(�Oa�[i�&��ev��$L�j+���aG�������.��ň�f���.�72��
�҅}��:�Gz;
�ub��w{�]>�%I����A����=�I|j]����0�h��2
Z���¤H(N&��[�1u :�͗ƀ�L+� �j˞�O��'f�n�$���	XX������'�}+��opJt+�q|��4BHvz���F��7���h?�C�O�6���o����v}��{u�da8����iܘ�>��3Q`\*'0����C�e�L3�ݯ�ը-�`�⥳e�����KFp�B
���Hb؛k��=w�:8�)H��i�iȲ}�����ށ��s��o�*L�e���sy�M�jA��t��Zv��(z��u�\�-H^Wy��xOUnit�W���qrm�����7�䏽#�& jVAO��0)@�*K��*�ӆ�bK�q�@o�u
R�#��T� �d��R�e�un��.jӡ�M�|d&5� ӡ��+�ִ�{�>�M���q�?�F �7��ddɯ]���@���s��DgD� L6����L)A�K���@T<��c�x\��ʊd�T*��_�Zt���uUy�得�ڟ���6�l�\6.h7x�����d\�{k
iݷ�����k.*��77-������q�x���E�ȴw|D�	���KD�;?~���|��vK����A�����N )C�����[>���O�@�t�\ۯ2kx�
D��~��a�ͫǓ����zdJBU��#��n�g�#��`Ŋ��)9�3������ �p��xa�5�yOؚ�ں�IV9Y���С��1���Yߝ���hn�f�CL�R=]|���$�����!�@���?�W�%:����(`�P3�����`sb�e���\������
>Ud\I����#�h=��4z���̌=�D�䑚rg ��k�|�~2J6��!FYPR��(�J�u���N}�1P��� G�A�p�V25�ّ6�j�+�p�������P������$>dbR��	�����\Ws�B-eozhH,:����}\��(�.������@�c�`ݓ���BJ�'��Jb��ƬrN*�J��r���?�����S�����1�K=� w�x5fj�hx��9����N<б�_�jn��@�����m�}�K�˧r��O�K�J�T	$�j�c��f���D����N
��]'�:?XlQ��e����&MOY�v�̈́�,���l��zq�ArE5)�Ɏ�����|���D�k�\W�v��̻�R�ö��r�dQ� |�=��d]�`ff0�=4��ZhY��Ah�-�"�0V��m0�dPϞoO>��Ǎ:�ZM9h`aq�*.oUo,�NE���To���^ۇ?��m}�t�ۃ�s�=�rg9���qvz���$��<�hH4��R�q���Pw��l�:,4s���'M3���BR"s}n׺d�V@~�r��L�AQ��쓼(U)����@�<Z���ڿ�C�V��ݪ�bʭ'ޔ �xkW�n�\��?�2G�#�,Z��@07�B�H|�<���P�r������	!�[|[�sd�����:�wH]
N���u����S�sO��2?�eX,��!|/�v����ACE J�a����}���l 9�/G�g���:=K$��i1��(c�ƝQ�"[Vtp����Q��;E�/́�i���%t�cabEA=R)]����mJ��p%�$��|sD(�V��lL����	�y7q*��db���_/���=�.���h��g_-~�ῐ<�& ����ht[�^�ߐ��(K괉�s�i랍̼�!]��uѰ,P���%)�����`�Df�U<k����|�@�#ֈ���u�?i�_�J5�݂����H�3��������z->g�=��*7;yCeƌ��.]hNA�����~��L�u�j s%nR�6���$1��`nM`GN�RLYL�v�S�"s>J~)��(Qd��Q#���xunoǳ��H�W3`�k�otq;-� ���4{S~o��ث��4f��V��h�p�\�G����4��>K����L##��W3�`[�z?�@/�Yo~3y��؎�##�'���t����7)�<�:�X�<b�g����ݔך�oA�M��5}�Ϣ{��N�_��$N��S�9��
d�9��vw\�4�U��:7����N�y7����o>��U&�uU'��8���\���zz�:VO�ʎ�-�o%���P�* ��d��?��+�*vL(Uȴ[�vq{K;%�W��P\J{4LK�i���K��j�����n�t�������9<�@�M(���L8��.d�����2���Y�JA�JJ���?0(���+��)��2-�o^<$nv�~�KӇ�X�bB��t=N?�u��7c�i�M��=a��SXY���S1t��x��ň]��S�j����m
��@��:�9)������eo]�T��[g�!r��٪�o�ԆJk�hB��I�c��yAXW,Q��0�oK�!���/T��ʴ�k��@�������EL�'W�J夺J��Tf3�4'GA	"���/W�M���'I���+J�w�]�Cyc��*B�6�����v�P�Q0̨���֧�'ЗP����|��44���}�^�U��A�h[��:���/�p���}U����{ �^���u���N%O�и��垾��E������9<e�zJ"�V�݈icƯ
@�Pqd��Q�xW�U��_��H��U�ub�	�T��l����e��(�9O�QE�v�p�%�8E$G����C\��!�xT6ݨ��3%�<�����_�9tӻVyǩ�o��\��`��a&����E-�V�/�
�m�i��68�?�B�c֨B]N x�����s��(� a�n�2@Esm�RD�.�r`����c/̑����L�Iy<&�7x��VŔ�I�Ali[[���pcn�Q��͂bւ����M�lg����3R��w������3لl^�ц�L�ɮI	�DB�R�^�D���0�B�a�O�}�I|f�4����7�y������و�Dv�}�":�,�"�@`�7�z>/`XQ���+�h�b��Z�����_��H�zl� jS h��[���g�-Q���� ��wa�}���ui���X����{v�K�je�$�h�[{x�8�D���L���f��~�<�\�z�V�~#�4xe��H��B�H�/��W������8mI�_�A�3��b&^��K�?'U��ѓ�*K��X݈���;.D֧G �X�ذ��B����$��1:흆�)*]CC\='��h��Z9V4C@�l`��c߲��|y���g����*�L���6�h̔��we��4��K��9�U"̳���u:5�n���Q�k5$��i�Bn]��b�-=�Ʀn��'�@}[�:��4�Aщ�Is�S��ఇ#t �:|��\��I>�/��������`U�d���,P�npyJ6+r�!͢�m&���{qY+|N��j��5�Ze������gʬfd>�\ܞ�oJ�aڃ��be�jh�T2�Ys���~~���2��p������^y4̊�hn�j���L9/3i,���W�	��,ׇ3M̨�6M�:P����WLLU�t������G ��>qm�'���-C�^��(�D�j֗����m)����"L�Ra�0�8o)�(�S����G$�V�sm����|�.�V��%E�iԥ0�f(�Uzx��O�0�m!�}���4!v��O�i�>wY:�k$�h�̡�y�K��rG��j�Y�tL�����z�]�=�r!���e�ӫ_���@@qN�{N�kXnQ���ǁ��� �$�[���P�
�W�ͯ���%]X`>��$v��h�