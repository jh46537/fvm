��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�/�CZ�08Kh�� ry�z�����w1�E�r�߆ݸ>G�$��;� ���k��o���,�#��*�߱sg�E�b.2H��
�q*����*�'g �\Yh�v�8 ]�����ce�;��p���+s��Z���'%�q�:���W�����R��6rǛ��� ,��-Fc�db~����Ԡdr�1j�Y_2m�YJ��A��%�N�D�'1(&Q`�ה��%���}�q'����r�&�'j��������^���2|F�V@�'/O'QH��D��@������QcZ�9�0��r�ΪR5w�D�=3��n&��-J��ː�By
�7��ne�!��.ܴ^?�s����S����/�@|����n)�Q��J����(Lߣ\��[�զy�/.B¶Fvr���u�L�eU����pi�
��j!WV�3��<H̏��q�� /Ѻ`��Y�QCB`0A�g���W9��d�f�|���p5Pr�`��24��,:M7I/�f�{l"�`�#;�
_��(�}}y�Z�j̆>��,qD�>�R�
�j�����*�����%n
�����@$��L��b���r+��sB�1�!�J������T�=���{(����+�X���%�P����ʣl�~����g���;a���xyl����$�I>������Ԫ��%�BXX.��&,&ۀY�H۰K��5�w����<�4��@��f@��U'`4�آM�����B��F]��~�T��{LS�S����?�UL����� �R���u�f����D�'2��U8����yjs���;@m�����BoK֬QpH�N�(|��0?��Y;Rԉ��c�0�Suz	8짱7����hU*K�^7�΅�'Nvnr��2s����sȒ�܄b��$u&E����Z-V�H�jQJW��K F��| �z~����'�^��x��<A�S�Ǥ�AB���s�8�!�,)&^��{�k�&Br�B���ʲj#�D�?�⁩))nW������O��ß%{f"m��R�nq!������}�"#�� ��L�
�%[�
�F������K+e�
��USHO6�\eQm��=���O%�/�*}>!�{Qp��;A?<��Ŗm�a�w�`(�#��:��C2Qj�r�MJx��wN�wq�Vg�D��e�_$�8����W�E�r�<�ewiZ��F�'�$�p>�v�-����Y�/��z�Qz��,����W��yWg�J8c�{��i~����󖦦[n�4����fҐ�מ�ng����n)��=���Ч{t��o_�Ux���-���ث3>�q�I����T�6lӺ�L�FVoe��+aSdm_������ ����M�y��ilб_O,��U`H��{υ)M}�b<�[���2�j��"=˖7�*�SZ�l�_�5,솗Ϗ�*W�!��� �{8��e���K2���d�a,�>��1��ʁۀ� �A�;u��\ֆ���Y�DF���?;��$R�e���_(|�t��0�)��e�s�<�{gc-_��ʠڛ�f:|�7���ͥk;_��6Q[���oO�$���*鑎�.��Z�	Э=�JL������d�Z<��ד�d���x�2�MI����V�?=���¤Zi w��]�Y�:�>�s_j���2�����ÿ n.�Ԭ?�6heU�d��#�i��Z�m����_��J�YYS�	C;3pz<��Iwj�h(��w�wl�i
 b"g�uG
ꥣ��3K��bt{�;�C.x���V��b���P�u���N�5�+m�A������{�$\� ҅L8�gx��_I6�Qzl4��w���a�1�KS{�w��{�����ǆ�?`p�uB�%^��XF)u'��Oc����eˀ'j��/����s����Z�?OE,h_�� ?���	���Z�7\Γ��+�UHE���l���\�|��> PÆ3�PM��rY�2�ѐY��u�M����0����
���W'�e�0�`��y�<�7
�<U��+I�R��3����Q�ғ0�S�C4d�5�m�ս�c�K;΁�ʜ3�pvz�i#�+�Ւ-
P�I,(�A��U�y�#^��k6�5�>�%�Lk�?���
�쳿b[�NY���7���Hޯ���$����uƕ���QA���6�ec��/�iNC�K>��f�@���R�:@��b���.r�:��8���:^8��-�ףl3�����
������3T�����*(���ou���P���{�QQv����F������H�t�\Y$�
��_�y:H�d��cꬼU�W�ir&2dHMN�L*�~ y��;�ƻG	�r���݂`f�)fm�Ǘ���?���#H����jF�hz�Y8l�u9^�����_�I�L�pBUW�N��~SS8H���z�s�W҇t����_���&��X�J�+�r��4�Ų�I� D�1ٚy��d�A;��P�'�W�T���)��a�[O�0A�Ɠ��ղb0U�-z~'���� �`9�O���*�'nK����Ƣ�
�7�����{�Gb�"Z\﷉���=|��H
8��E������W˲)5̔��u>�%(."Ig��_^��5U���c�Ds�GR,ͧ#��7x���g��?�ԑ�,�r��`-q�l$�з�/��=^�̽�J��^��К�!�d�����ꍅ��Ix�}��������к���b��c�#Ֆ���>����`C	)�)h����&�U���L+G �2��'1Q��7��Åp�*?.�B�뙜
S\0	�>�<�L|z��4��He��� IuJP�Qy"[�۳|b_)�[����I���[�`A��,�0IS��
��#��\�͆LLؽ��[�&�m����S�v��S~�	c��
A�i3mf�
K����{�y�ޜ_�E��8�׸�y������?�����*��Z�!�}�R� 1$��I��Ś[�x<�����r�(�e�R��Bb�״m�iJn���1�3�.�c]��)�gJ:��'-�|�����7^�@4!�^9���F	xW��C�z�E&:f�x@t�c7S�08����m�k��ܹ�W����eĝ�������N�M��P=�.���I�Ҍ��2y� �����nl�I���pY7�@j2faV�A�~�ݣEUw=�يZڃ�ó>t��k ��9��E>�^���	���0��*������3��z��BZ�$�Ϭ�\(�~B�4�,8�</h��~{e����tgQ颟�ۍ�� b�ǃ���� Ox��Vd�_.�R�Q��\~,`��XY?<��D0���9�ְ\��*G2s�|��%e�%VO�~��\�J�|�B`���b�� es+	��˛��\�E?)�K������R) �dWS]5��F?��B�3��f̤d侷r�Jv~]���eʩY��^7�7-����n����K")��s��z}�� ��i�I�ށ���E�$���C����,T��bׁ{i�1wx��ٰQL���� ә�w3��_��Exc\v@,�Њ��v�J4����[�:��DGm�F�m�L�ˠS)��]��x��5h�t;˗���w��Y�`�Ic�#�S�]��8a/���Ԗ[4���Q\7�?��1���g߂o#�{����S�&LxJ���."j��4t�&}3��Y��!�s��f���[,w9������c�gRy�R�7-qW9o1�}�,���`Z�$��ӌ/�~(.��&������9�����s	_����B6�B��r�I�8����6�9�v��I��cU1��Yh�2.&����O��&Kw�;�nrc-����L�&_��و�p`�.h���m��\��R���<�c��b�Xo�dk�W�z�Գ���n��f�3/q����+倔�������w¹5�a
u��IkR���|�ά��*���I؇�V5�ڢ�\?�i ���+&����Y
z{z}�ֻ�3��˶�^3AD�������;����b������ɋ�ꈄq��j�y��g�Ju`W��<�y�u��M��:C?�b`,q4[��6@�-��<��U<[Ĥϱ���x��* ��g�#��=�� [�
��!魂�H���s¿p}�_0?}� �LϖL��8�2�6u9.1��E�+i�A��~����'�pZ�1����U2ȣyo��-"	�w<��F���㒬���Hӑ���h�tQ�&���D�@�t��@�~�ɲ�5��5˖�_a�zM#�i� 8t��Ơvo�#�
�m����e�1�-Q_�4�@�V�l��)�[|~fz��m�2N�K�4����T�u���<>M�X��z��2#i����9:�-�;����8�3�D�+���٥"��J��.AqG��Uh՜5�E�ڄy߻�,���᥽�k*�#?��� �#�=/�g�����D�nw�#�ڎ	O���e&=r�kk��y{�G=#o,�\����4�Ѓ��4�CR��ʝ���=V��ʮ���;u�)I�U&�e���d�J�);��-j�E�n�cv�8�L�n�S
�����ӄ �����SAVvI""�Q�Ć:ǨgK�O���}���� �\|ǹ�8�H���	mZ��7��1�S�ڂ�y�W����P�^�ϗ9�F��� 7�	�a����3����^��~�t��v��>f��;�+�<���=U�P-���K���!i�R��̫fE����qݥv �J��.��.���+�yOM�����Ũ���B�P+ ��6l�s��E���u�Ѽ=O����`-�3����4>)_;�V�G��e���h��7���Q9�qN�������d�1�n�BS���I���x�_p���ZSF��.	�k:9[E�V�P@~Rm}��@G�Q�;��?�F�σ�y^�J'}+��՘:�sg�V9	�G2n�Z��h6˫y+�)��A;�g܋-8��u)�}�`�q*��=�~�z3��l�p��"Rhg��2˱����[��RC�Ц�W�.q"��G!�k:�T����7���;�ԡ���>�U|7�R祧R@F��p�2��BCzn7���L������lr�p?���Y-�\��Y�Ԁ;�?FILn�����Ѡ�