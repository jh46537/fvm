��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,�������_^�6�3�@�RU:(�3��j�0��w/��e�p�@�Ô(ޥ�#�Q�|���~�GJ��5�/s�t��N��.Z�Y>z�d�K��?��[�݇,��5L���w6>SJ��ѿ?윪ik���(�3 ����̾�V1!��x�z�tݥ����Xc�����%����d:[���q���ab��.����{l�E��M� \�م��}�ю�t�(�a�{w�}�$�����܌��W�l����M�Zr�8��⾹_~�1��|m'1�FoY��S�y�'{��"iDe�&��O��Urd�C��}�5t��e�ʂ�]���CxX�|�y�3��^{���C���\���o(u?�x�'��+����"����
�Ν�M��
1e������f6	�u�L���d�:��7Ok=���ժ.D}�dH��ʘ�j�kqI��xP�K:X}զ�ah{6�FK錇1}+އ��u ��7G0��#�dӀ���e����K���	�(�2�Ĩ�/Zx��g��tK����\��a����Ų523fUzum���5�Z��3����|ǊeR9�Iɒ)4�m[3��@�9��C�F��N���?�.�A8Us��B��Spesb�{���t��B&g[��3�˱���)C�毓�YO׉�Q~��������&�i鲵2-�����u �ެ�S@JY�{'�N�+F0V���0�>G�r�K�I*"��_�G�OW��1�ѩ�>�������ڽu�.�>�*'R���Sl9�3 
�=��|��
_.��[4`��<n^nJf�д5,�*�\o�'�o��}6ek3�uYǁ(wg˻��铝FO����W��b�Q��,�c�h�NEPb"��8H;�Ѣ���3`��l�%�rY�ٮ��w	%�7uc�l��'|�E�$�~��6t��U�E��P�|���^-�>�`0�*Q�6��v-j���Q��ܽS���>)W���׷�v��t{�����T�����j7Y��O�/����`c�<C�*E���8�)I��J9��� �˛�����7��FZ�p*�	�� ��!��&qy܌�
�_��f�2��ha��ၜ�<��}��UbY=��i%U�0Q��ÊP���7�I�5�L���vئy�{@�8E4���5�"t����]@]�y�ܶG��ǜU@Bb��B���:������� �/)<��8!��f˯3XhE�KE�@z06K��P��0�r\����W�)�p��Nn��|�{�ż��^��F�׹2� ����ٝ�z(�OI�UT�H�ǎ��}y-�5R̇��k��] 8|#'=��"���r��藣T�-R��{- �^��%GK��=I�[H�z��K=���±�89��<	�٢�v�D�+�%��0�"يZ�C ��ɕQ\'d'�B#��a@ih��\�wS�,U�T&M��@?����BdNB3��!�1�1��n�o�@lw�F�İ�`�*��!6]�B�~�l��� �e>����	�f o,��C�;b�Ū�/7! �G,{zY�ik����_s�Z��.M%��
g�b�Ư������+JM��ڼ_�V�Js��<-#?<�t����e9�C�uV�:�G��qO˾����;=����޸t1�0����[��Bkd_pB�q�8��F�����