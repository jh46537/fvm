��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{���b�e��_�@�*��Ht�'�>��j��vm�s���ӯ��@�"�恑z���|`T�iݍ�2�Eg:[&x�
8m������p����#�K]Ϝ	9�gA_0X��66�5��X>"YR�a�b�f!�.�#�c�E��"��5p[v��(xBg�������\�'.ؙ-�S���[�n��2�A�^l��k����d��2ގZs�ѦC���
����d\�����!�G�[>b�<�ŢrqB��.6EL޼:�u�S9͗�UO��D�%/�I�H6S6���J�E<��wՉ���ŉ�+���,�$sr��O���lg *Ǳ%������
~Y����$�g���X��R蕛0%�l�����}D��ȿ�,;�M���xP�#D�h��ꌟew�C���}�-/�	�i��R9��3����ٝ�ղ�=��'�ފۜ8fT�t�4[
�E�g��D*̤�����giff�[��DE�ޅ�Ky+zL���S�^ (�Փ��0:�N��[/U@`]�-��K�=��Y^�Q�Vi)�f=g��vͤ��?�Tl�����:d�Z����]�Q�"<�͎��|E���d��T�!��}Z���7}���c�Q�V ������w�d�>�����"��-㾆�����g\�Ѯ���O]v��o�2N�Y֞���x?��':2�������n�����wW�����M�ζ�<܎�[��v������-?��#���]��k�X�#Y������'W��
hG�.�1�.%�;hJ�) �ډu-��%��2����vEA��F�I�h��"E���:�;hqr��Be�2仆Y;}��#Xֶ3�V×ɫ/�h��e���U��4y�_s|�s15�m7f����5i�_�����x����4q���>*Z�K�����\�PU�7��\�Y�6F������d�Q�sQ<�~��:q������Jd��	��]����جC$ӭŞ� �:�W�{�U?���n�u�4���*�J��N�9�-��(�#ح�F>�\?M���c�=�����8������G�@t__W����u&rω�'�j�c��i)������3�N�)qdT�*��*"�p�w�I�D��1$��е�Uԍ�$�F�C�!�ﻭ��15�ץ3 ��"�����|{����VkS���K>/���T�*����ju��!ݦK�ɹ�E�v^�K��/-'Y.��]k#�)M�#R���J��k9R+G
{�����97U�t9�,`a3�;#r{k6�(<���N�d!7!��JD~�[T��хGUk�(����^�QN ���Y��}��1��L���;+����T8�]�.�WrD����Zn�<,���n��������$܏2���w�E�`�I�/��P��]��W[�/������|YĂ��_CV8�M��(�ԩ�����J���W�P��re���`�@�ȿ�^�	����?v� �
�R��I�X!R�Q7��m0�~J�E�����V'���\��U�l�n<W���)��T���9#?x���]~�?��%d,|�yǄ��t���z�1Q�vZ���x��Ϗ-��؇�iI��I�� ُEv\�r��ӀU��*�e{���QC�v���(�9]����xf�X�|,�v/�Zd9��1K����($��2��zY��yW̪4A:�P�ܷό�&�!Cxv*��N��9�
l}���cB�J*���@���SH��h��~B�y��KJ����?t2F���1�	��k�����f�{MC��XЎ1v�d\�6�n��lWH��\�^F?�c�v��
�� S�(�u�bϦ�S{&���un<�0��Q1��0ꁼ�㟓u�Zgg�J��sP*e�}�w���@d��X$O�߆T�����n��k�4�>q`��Xm2Duޯ���͡1�~+��dȢ?�'�e �P��H�N��8d3�Z�Ntܛ�����z1�aN7�EҮ�S�f���8f�)A�&�S�\Y��v�\"u�Ɉ.H#�m6c����{�Ǹ�y��*���%�d�q�Twj�ꮐYw3)f.Z\�'q�G��[�X@�/��Y�\�  FX���c\���~]
za1m�:_s6۝���~a���,�c�!ْ�Y����MV���6��H�m-�b���kk��n��HCR�C�=�N.��\M�>Vk�v��)n�� Ŏ8�$���!��'G���I2�m��:�cK����M운�+n`�����6z+�b�R�	׳Ϋ=�������AщA3O�,<}����p�ķ1�$�S>�J���Us&�1�����N�#�#ӖU�
ȫ��*��$2&!<g��{�������gO���;�H���fs����^O�������"��}H��73�c�u'���N3��f4mI���ܳ�O �/}����P���c�;�:y�(���y���ȶ׾��\�)���Ur��,����r���o��ĀR߮$X�:#��<k뼇,S�ҡ8�^�0L�W[o��}}}���;����K�����iސ��Ka��xY�kd��=�WPD5=�.��	{�f����@�Y���˵	;vu�z�hVC�5؅�-�R�ȼoq����+t�n��ޟl�x3z#a\��h��4~���&i�Jf���[��O���u�&��������>2�@�}ψ�f��<K�ؕ��M2�S�eO\CG�t �=j��U�z��}��\Y^�B��u��׼,�uG��㜘R)��