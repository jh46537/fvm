��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_R����&�'���La,�)&ȓ��ܥ���H(ކ�qH��t��x�ֽ|zP���ɿ��Y��Xg��VU�2}�<�z��Cƴbc��^T�d�%Ƙ#�C�{4�6��ueT �EpW��^��<=���0��!�-�oG�K�	�)�ܿJ�vK�#N$�PZ�8VS�p�0Fn����#������2�`G����X����֮*�2�;],e���Z��� t߻�7l=��m� ��&Z)���G�Ɠ���n��k������#|��g�����ZZ��5������ݍK@}�l~�B|Ie���w�Nz��)K.u�F�Zyf���*�mvkm���a��q�C���)_*8���'K���ǭo7|D�P�6����h���XF��C�*�q4���Ȇ���$��#�h-܇pA %Un�=�%�[�
w�;l~�DABT@O�vxȾ(�d+��b�<�?"����oG��B�3���B\T�#_�@Ԡ?���k�hQQ�ro�	�;������mx����D�vl��6�:��v��R$;ޠG�#$��ʵ�C-�z�ݍ��[�J�4��$n��3���v ���p�IHD/1�uZZ��]g��S���
<��$B��ӗ�8Y����N�%�L:�1�wK�huZ�����&^��l��'J�X��k�bm�ߐ�J�����K�'e�,蘸��cw(�$Sj�`'C�g�E��E����P�e:���YK�-��h�`���l��0-���S�ש�gB�{d0P(����J�<=�Q�f(�ͭMGȂG��<�A���"����@'��v㻴2�Z*i�'޺�˹�	��0$��m2��=�}L�OOX:��(�m38�()⧇���y�����ɶ�-s�P��j��)_1�)��-�n^���.��ck�G ��uML��R���b�Rn����Mcj��
B�m�T4_�ƅ�y8�u����kt�|�0���~o1��#K7��qS��rƐs{���(��#�T�vO5�۹(5�ex�Tb:x��J=(�����ZK8�_�h�Б��]*��|7�6�.:e����,-y��x0-*��F��P�H�^�ѻ��Y��'k6�� ��N	LϴD�A2@��ҹ���{g�As4Ym�A7CR�ϖ7e�dJC�t�=��{�Go�o��5N�E-iX����	94)�b�Qt�K�ڪV�.N_LAa�:��Ud�,2k!��H*\<<�L�GSE��Đ��|�S�j�ط��������v	�SZ�Î.��w�zc~Oʊ��7�o���K������,S�rZT�U+o7�x��?�̦W�!�».WdC��1�jo4S5�+	/��J믺��:��5Vx�}qK���j�׿��]*O�A,w����a���DQSu�sbI q'� ��kmR�6�������}��e|3�?���b�zW���X���@��ݗ)�����Rk��2�&x!� z��3�c�� ��L_$7�tՑ���L"�k��8|����/�05�B(��F/�a0�m�8VHF|��@L G̼A2�~��u�\� OR$�3���#���|���*�����>�(i\��3��{]^1�;�4�t�����ؑ��[�%`$�wR��j���i{��F��W������>�ɿ�Η�s�Rπ	Q�ā65F^2\��ڤ���g<?�S�&�u��)�o��4p��]�--:a�LHM��6YZp.�$-S]^v%asm�2��-�z��:��r �������"'�;��9z��8e0����-����'?ON�ua�q!����l�ڬ%<�AӄX9
}�|�{m�u!X�,0Nno�&�<�?���nF0j���^v�nv(�ilp��u��a�H�m�a$��$����T"�Pr����#����sU�IZ(�r���X�r|/]�F�fh5�R^�=�d�S@�S9B��(�&?p�vG7.32oϼFmX.RԤ�q�6��3C��k����y���b��$�Y�h�%MEr�]�a�k�o���jK������h�O��or�����B��:u����b���0.��V�u���1���j
+�&#�at(��
e')<0���^�e܃���p7��Nu��^��[?�ܰ��;<7U#�!�����/�g�S�=sr�]W��B�WwXPez�>����W;8��u�
 _�
,^klGw}��&���M�Jol�.ln�����d�.��.�� �!爒#�?�M^��A)��A�����n	����˘�u;s#+��(������~0�4G3t�P���f��X�*ۑ9��F�U�2�%i���x)r,*��2y�.4X-��2�ѴT���A� �_(�w��Wg_�
���Y�Bwn�\����7�U2/���d<)��F����L�V��n�c����K��^>	.�5�u�_`�p��y���nb6r� ]|���+����c|���F�lͺ>�|�0	ͩ$5u�[�	e�{7��o�OW�I�vY�TNZ���@ ��<����ϛ��Z~!����ljp�8��)��6c,]�lyŹ�i�MkS6N�#���u}�g�vri�@7�������'�,�W�6���;�f�q��W1�.�@�Iћ
��C��)��&�wq? jȠ��+j�g�H����?�r㤰���|��w����DY�*d�J`K1a^�����A+��`-���ϬS���߂�2��q)�e��k�j�+.Jo`#�����,s��@��0%u���]Kedk�+	o'��jv�E
�S^:^��,7|��͛Iۓ���>���1�ާ�����
[3�(&�xc����_���	�29�Ճ�}�H�ٜ�Ly�Ԕp����"t�zUNp׭0D#���Lj��]�ڄ���:�nǗ�#"���?����db��M�S���u��f�!��ED 7�M�u!�-�N�y�׉9j*�|����K�|r"������O�p~��auh?±T�81#��Y=���+dgK�N�z8Y�}�׏���^*�cd.�\F�� Tӑ�	�/A�v,X���T�4�5�aG���1ط7T� �t���7UL*�)q.��A0b'�����BW���ל�o2,w�~�7���Ѫ�A�X{7z��L���{��=� ,�x�$�>���A�jze���]CˡӔcpb���Y�����x�HoY)� R'�1�iװp�O���L���'�nq��|��Fy!T�Ф�D�qJy���9p��#�s>��J4��Ì�����G���(�S�p �X>��2J�;gg�]��G�1V��5i's}�����r��������������\P.V��(��"�X��[�PJ�"�$&���J����d���l�@鰓�v`�ng{_�8�p��\J&7`=�Ю��-C�g�18�X3rC�-�C�]�",�һ�;������@�[��ཏ*��4���nrNF�f�Jx�Ώɘ��Ԋ[lΨ����4(y�a�Z�����2�p��x��o�g~oȓph������bz��"3���j]m2kt75Յ��?�-?2�̚�Һ2�j�Xz %��փĦi�?}���2�Z���f	|�(����L��#�qMƪ�fc��9Ę��ݽIT��ѧۀۑ����{\
$LjU=��xӗv�6����t.�4UO�G�����B@P���F�A���l���}���� 8�N֚N�$�n�AQ����g	�[���� ��Fڨn-��8�[��{����^K��~f�D�_qTHi�q�|g q��V ��+�$�B>ե�a�q٧Gfu�$���C֦��;׫��:���
l�^xf�|����T2�������]|"X��z?�!l���V ��d���h�?�ġl����Ժ:���V�QÑ.�5����hX�|0g���}k��ƞ�1�����HYBrV�6O�Ӂk��J��+�m�rϢ�O,�XЯ�I�Q#��Mh��Q|`:�_J䠁��FA��iJ�G0��s������5��f��$Z�,>�q��(�n����O��)��ώ�s�?�>�M$TC���ߣ�g��\�# ~��1u��;�?hH8���<3�twiu��v�X��7�CѶwUC�����]@VŨ���L��=�EI$
Џ�����5�r`�F���R��!�6��5|�hF?s$h�N��?�EZY��v�9� p�t�@�%	>"-��|!���ڕ)��^ה���"���g��֢G.b	e�
r��*�#`=i_����--���?n�O�݀g&�n�i0�ҋ7�3)V5�SBƺ�FD�̤6�.�>j9�����Xwp��$ι�5	���]�O�����G�.Ux�L�[��Q���ڹ�����x��,���5 �v�)��Ͻ4��h,�*2j�>�wH��V��GpVз�'�2�d���Ӗ,��$�0�5L���:��	g�1h:p!��ws�`�0����������Jih�Y���)�[ޑ�nR��8��ER&S��y��� ��S��{��^�-�P�N8WA�$�~oxlL���tN�>�ס�����[o����t��|������7/|*'p]��4k%�\HdZ5
ΘЌ������G��x(z����r^����!�\Rh��ˢ����İ��QsTeD*�ܥ�ː+N
�7�1
��s������Ԝ��Y��Qta�㮁VE�I=�|e��W/u����rhe��Ú�9:��=I=G e>_�R�{��L�8�f��#�j��i��a�Q�y�R��h\LN�(�����Q=]�6RK,fP��h�>�+F��&�&5���<tQ��J����="F�N�M��ma���'1�:�x��8�d�
m��DG�u�O+���� /�5jF0��%_T�*9�[��Wō!�wJ:�?K/y`R����m�<��[ �&�$}���4в��Nd8D ��I�������>l�A��*�<�C׋�rV~�I6�:�����O�,-����R?�8�t����N�5��=���y��a�>��u{�}���;Z r�v��\���j�^6e��b9�yk��x���gv��{L�b�/�4���e�R�n�3�<��:s���Z � a�R�$�.r�6v��O� �L����7�oHY�x� �9��x{ ��n�U�ȥ�{� �
_�əP�:0Ѣb�m~�ۚ@*��.
$WŻT�PD&��A��Y��Ǭ ���6�hN�O���tNv`ai:�*�3��}1�������� 9xQm�zq��7^�h���{
Hߗ��Uh���myc��0�B�A��-�c�Q�*�=C
d��Z��wZBcÌ/c����Hu��e������|��*�z�>,[<��۫�K�l"���)���$1��.��T3�J����ܧP��L%�����!��W��F<<d��κ�C������Ci���uL�Of�設���&F�<Z�^�KC�6���Y\{M��}EL��3&'�ڽ�l��ׁ��bX�6R���4@#��>����C����FD������hӱs!4���ˎ'�@���-%b2?�>����В@�>�u��Y�O�F���-F��7�p	:������6(�\��L�62�Gu��7�L|$H�9}4���v�~I�:���ƢT����]?`��n��$[I��s'�=���j�y��s.Ѭ����d�2+��%��g-��;}_6@�J��A��	�w�XSޙF!��@��&l���a�&�_ ��#�uv_tl)V6�R;/1a����āMߡ��Z�2d�.W���ѥͥ�7�$4�c�Lb�8���\���>��i�#-���!.�v;P�-��GR6	�^0FA"^�3Mؚ�V��N��Ȥ���G+Q�C��;�<el#���rOZr�uP$ mEY!t�r]�g|�*)`�!�\/�/{kW�-�ML��2<L�^Z
5�~� D���*Ң7\Wᥩ�*~k輍��e,�x��=�� V���@d[�P�������;�e��;�5��Z���u(x�5?����ح�$��<�(N^`�#Fd,zJЂ)��Š��ۿ9����@�W�EAT��j9��r+�TYXj�#iDp�.���n���dr2^���nY�"�&)�1ygEL"u��yt��NY���L �V�Go�5�m"�C����,?="�#�������9熶y�����i|J�1�#�-u=K�aiIW'ξ:�B�9�r B�k�Ԧ��8Ã��96�}-^���YV�/sY>��Ĉ�f��hl�J��M�N�6X@�}>~ P��T�}!C-��A��f�	A����<a"�zU>hӳ��q��ܳ��^gj�ʰ=H������c=0�P�u�Z�x�園�)-,�}/����&�P����쵎 � YTYwW�mL��^�8j� {����f��%9D��9��}"(|�uᷲ��o����v�v��q�v�j�� Z��ܥ��ϖ��Ȍ���\�JfZ)�i��Q�-�H�N���(��O��~������m�p��q�`���<�E�4���n�#���#3��+�c��83E�*����3���ʓ�.�Jq�5JĢ�<E�N�����<
RD��+᣼<�r�3h<d����@�_E�1��4Β���o�!ǿzC�y�c�C����}���|vz���Y;KWz�ȸdQrG���98�%��.a��L��7��y�����o��@�u��ާyj��e��`�툴htx�Ż����n��O���_~��dD����#�S@wM܍6���2$X~���#`Q��qcKc�A|��*&".��˟���y����#���҇�6n�N0�Ԁ3�	����:���Q,#�̳��%�0˃�$TTY��	�oҒ�NSKK���xc_�'�k���F�]�'�i�X�:��+i}G�vA��FF���~�s��S���wN���f��;+�2��kx� %,-��5�O��bOl;\��,��ʒ@ZUV7l[����;�VoT�K��s��Ԓ���_���d&x����v8�>�4�=�8 LJ��8����WdH��.�٥���3Ő�ܰ^��q�aVY�{�ǪHS.�ss�Sٜ]��3��貓��=k��@]M��dFC��Br²�@��x�=fc�}Vm#��K*NN�ƺ�3%�� SF�xǗS��c/�q�s���U`M�}~����$���!�]3ﾶΪ��~�������-@�9���W�)8y��������z��k���]��lH�-U �#�Ǣ��َ$@�H���B�}��,q��4d-�P
�����g���{�n��N�^��4�D�p�c9,M�%oJ�U�q�׳����f=e�%0@��9�>X���/�is�i�������!���ֺ�����N�@�wC��"pNJ|��n�e7�0[��H<�s�P?��j"�K��a���9olK-�\���Ǯ8�Sw}=0����n#z"dh [n�w�8�R(�%��OMse��:F���2���A�PC�#|�껉�<P̻�}B<S��r$
�Tl�8��Wl�|*�?eRM^U�M�.u�@���}���W�azZ��pX�����^2����Ѻڮ�~t�%�Lы�+�=���:&ǋr�����b(� {>urd 7] ��=�"�ץb�bK
��4hi%�Q%/��Nh]�%f_x�s0Թ�Pe/ї�4iK�m�v�c���=Mx���37�l�u纩8�����Zy;+)�8���V��(�&-����i��S���.��<^�:0�0#�AKCI�<뾣Ň�z\��+a��c�����0���DZ��&H��f�����`��k�K���z5h}���C9w�~���QF���N�9���Tmy�Cvr�f,��0�4/a�ej>���r��C�~D��zwɪ���5c��s-�c,!<�n�V$����++H�^��,��BI�N ��[�����Є�B���k����t]�J��S�`�uU�Z�B�g[F��d��֦H�.Tt[��%�(�Z��N�S3�W�=�Gͯ�1�Y����-��A�:ɐ.X��'��&;%�~z�JX��t�p�IƘ�Ґ�� ��V���R1B���&+ѳ���8h.��M����/�H�O����9�t0 RR���3�ב]�(���/ݯ�ޥ��<��8\�WnW:T�
��#�܆�C���Z���-5:�Og[EK�D[�Wl�fF��;����}�@^�Q���Sq�|V�Hn�=^W���'���w@Y�4�E����1���/�;��>��~?�"�Ε�g!�����͊ �Ѵ_����t��h6R-8���Q{�n����%I��]I_�ǶE0����_��Z�/Sn5> Ŏ�2���GzK����x�B�A���-������5�A7��ϱ4�<\Ec���J��q:7Q�n��Y� 	��Ӽfg�ӏ-6�a�
J����9wa54]���s}�n�2�Dx�r�����ʦ^��S}����_�x
>��PE����6~K�Y^)��T�}��'-Nĵ��|wz�P���:7P�����mQ-�A�ӑKx��r�������:��»�u#+�� ��U�h�s~��,Y.2���W�Fq̿[\����6r1�v��x@.֘�i/C\�x�oMZd���$j^ y�K�WC9p{��9�/q�Q]ë9[M���X.x�����%ƃL˧<�^��}*�`��+��
�1�,����F�~�Xe
���롤v�k=D�D������i2��Ƕ\�!�>�,.�<1\#i�C�X(���`�e���o "��
�2p.4�䏡NC;6�����@u���-�:�p��>I�0;����yڝ� 8o}:�m��J;]\H�V� �gP�k�wн��Q��/Cm(ː3�ʕ�TǌyM�>:w��c��=��>'t�vy�����K�Wk�U9p��L��J���_��QԳ��h���� K�|ܼ�_(��i�)���+A��f|�S�}��zH����3�q�τڧ������ 	�KT��?�m�5óOY�1&��ˍ ��q�*S�|KE�PR�����d�#Kw�'fZ����s�
��Sb�,<�EyЃ���5�P]�7�'íg�Q@̽k�5}P�(Yr�m�4;lSPK_'O*�S�w��9'E�,6���b،Flw�/{�熖�S�]h�NͅE|X�H�"Ь�zӛ��ȜL����N�z��)�e�F���l�� �<���c��(T�{a�&�$f�J��m��_�襏�m{*��jE�=��I6`������Q�d�g�v�]�!mӨy��E
���֣��'��'ݒCF�1E��T<6nqB��3������GVﰬ�=zej�x��w���b{�=�����U|�(�,m./�ף�B>������"���#_Qʌr˷We��H)U��Lxt�`P+]��.��2i�@��ȉM����`F�Pn��n�ږc(�rB��f�^X��;�"��$��c⒌�����A,(�Q�G"��u�R�9[�s���pk�l\u/��>�$Y'���ډ��ú��4 -��9�}d�:�9�p����qN�9���� f�|��v�٫��X7{�e.����cw�U	�����dVc�?c���u�B�Ú%$�j&��� k���lK0�ܮ�(�p������k�x�%4"*��z� ��!o��B��|Bӭ[���7�O	�\~�.Ƴ� Z]�Эu[mlR�b?9r(��/��{��0���wp�]7p�}4y���v��uT�3LR�~Ӱx�;�N������V�6'�n��q��Z�_㾾���I��1��jC7�+w���'�ЏE�.-�R��"���<�W�_�+U��)�X�)���tn�-���5�X8��&a9�n�K(��u�%�8��CZ�����R>��[��Ưh��<-����
