��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���ymc����#��בsb]bJ���۶�*s����vhl���QE�;�����*�A^�?8L����F�z/+��Ĺ�Y�!�b����k6�A�����B�����E(Gء��������lrWP�G$�H����{��K	>C\0C+@%3��JV6m+�@q4:S�����g-�$ʑs`�*}�6bR���%}P�(>J��,<����}]7�(	Щɴ��u��&9��� u��RK���,��W��|�6���2�x6ۉZ�4'%��AzZHV���詅��܏ͼ7�#�����5�ib��K��~6U�;�w�x�:����Jک�;�u�����=6�}H[<�X ���7{�t��;��'��~�<8�KHӢ��"��NJ�,��ؾO^�B�
n���d��N�Z���[.���@�%��$�ʿ0�1*Ɣ���R�r��������d�-�h�u2L\��ݬFSI�*Xrۘ���TGVX��*�<�Y#f|Y���`�3�UM��]a���<���*���ˍo����H9�������A!��o�)��aE��#�63��Lw���w���G�F)u�Yт���,�J���`=�N"P֏E�"5�I�����Mo�f�w^�@�j��ұya�п莏�j�A��1#�{A�����\��h�%,]���Z�F���G~�9!��ERD��O�[l�a�G�b�(*sR57����=�Rr�l��<�@�:57hۤ+艇���x�}�⊣:&�T�3���.�J$k�
��^7:ٍ,� ��Ą�|!�2T��[�aen����<��=V�I;��%Z��	��[Z`݌��IYn���n�(��u�
��k�z��-޸3��ݸ��h����9s��v!$w+��_����>3?N���o�������-��
���"������^�������T��y���	�w)�"	��:�u星cm�yy>��ݓ��JQ�L���o�3̈��`����\�gŔ��7�0Fy��8=|A���y���6����b�z�XkM/ǳ��;̶
��"��UP� H�nP	�a8��@N�4�})�RZ7�еk���?1	pH�z�뵟�j��K?�y�����f�b�c�gKG�K�P,��vk���>}�� ��e=��T7Q��YQ�m���!6A_�~IP�`�H�{�/���G��l^t�LI�Tޚ_\��-
NO��s�w�
p5Jҕ�j��9g]7��uB��B��Sqn\�,7�e�z�p�;:�!"A����h0�^�ö�� ����&l��׳���k}��tn�lg��Ǔ��"b ��|	��sF6eKܮ�ǆ~����bY��,����%?9���0[o\ԏ��F�u���Գ�D�Yk��<�_^��	�,�]�P�J�Ҹ-eDK�GU�	6�_G��DG�uF��8����YеV����Ȍ�[0s�kE�D�LKÝ��W�c©�[�ñU��,�] �dY�f�p[N�,�����N�XQv`�믻���鄾��w���A95�2��V��tqe�<9��Jp�6������\�$�K�3��oS�obZ&9��,���yI��8�������w9��y�8��T�������]zu�J�`�����Ô�p�O�Vo�������z�ю�=�p��`r��Z~����\�{V�N�]&4���7��ucܔ���N�KC��E�CV��9`�ʹ���f�e�d� *��+�zr4ǩC�JP�G�fwj�W��4�r �����n��ȭ�ќ%bJ�K`�ˮ�H6�F4�9D�����'�p��0a�����ry�g��^�{֎8|���P�����ӆ��|���n�s�M�UA���������3J��sc_'Xn�Do2/�M�]f�Z2�^�8��&>	�=�C5�?��py/" T�.Uy��MD8�~I�4�����o�Վ�@�}�hk�����?�t�L�3F�rT�
t�Z�"/�r�����-���nP���'8���IeO+�&~�p�Do�bb���;�;��}6�+�u���*���B���&e�i�_�b|D~H��xO5��/!P�Zz����2�İ����A2&G���%U8^�h���4]s4��� $�9�,\ɢ�{1��m��݆����8�U3��i���G5���_>Vj�9�h#��e�ܶ���_L��⛞�3Q'N].��S���]������≤����9H�%^�ߧE��ZF���tf�d�95��R[��h�<'��Ĝ%s�'�[��<.愿,IYdk�3�.�A�J���-�ju�ëdES"���Qh��U�M]�����*�nCQ��uF1.TY`'��?���G�K]1E��z��<�/3���7l�JS�F륞�F�H�o��D.����Y��Pw6�/��mx�����P.��Ŕ����݈���A�c����j����9���|f��O���A�TVU��ɸ`��Μ�p�>ڰ/E�����;�g "i	�CHb3,��7��I$ MC���/�cOF�c7ǆ0�`�@
����Ч���@�t_�l����{q����Zz�����#��A�e�����?R,������y�sx���^}�<Ƥ b<1VuT �� 2A0�:�M�"h��lq,*:�:�ùfO�
��z�pn|�F�<��_Tka�ybq+Thl%?B`=�*�}��͸D[Z}���D������V��Ӌ����hB�f�ix�T����<c�z1s�����pSLȣ���&i�n����q;sV%�m�{; �,��l$D;h�����Em��+���[����%�E���,ʼ�@'�2w֕�7zk�a,Mae	L��1ڐ9M���z֊X�ۈ�-C�����c\��r �^�|1��w�9N��".�+�6�
0���1�VRٚ����*e!SAr��k<啥<m^D_����d$��h����ے,�sxD+��@�P�^d�e!�a"�mU�C�3�,����[����J�'��]�H�����9�$1C><_+��^��g��)�&nrU�[5�u�|&|�� f8�a;��	)J�\ r�wę�r����Ћ�ћYt�g_Í����r�]�J���3]"�E�S��(3�.��+,أ{��e
��7��x��'�<���<��@�tlL���yD�����|����3�BmL�t���\r�0cx���9_^I�x�P�]����5(��;{&��?t"�ͪ _�����|��N��0O`*�Ù��3�EX� /�w���ܶ᲎C3�'���]�M��B��Z������C�3�P�)sik�,{�
�����[��Wz����bSLr�>�)*���G����疻.A��ړM�x)���#}z<il��R1���	�g ��(w��)�dt���[�n��z)��~JKQ��h;�6�J�i�b�(�B������?��Q:��-��r��{ʺ
u�ٕ��5��"	D�+	�Y��jC�u�YC5,�xo�3+~AV&̜q��>ˠ	�cF�Q$���֫��11���9p	�p<^;�s���+�=:r�
����P_�a�p�u}!@�Q泐#1�� �<�^���O�o�_�6�ر�����m��IG>s��_�/�Qh������e�H��{��c�
���a�9����+ֶZA(��T����ˊ��AYل��T@o��K�ІbIE��(�ʊD��C�v��	`dGf��!����/����t�"��'D��Z�����=�ډA���s�`�������|��?�ح�Qe�$o}A�?՗'E�"d���&�q�zjB'����)���6��d��5�5�1�kҼn�M*c� �=����TG������F1�hG�7�Yݬp7��0�%��p�h����n��NY������m��!�w��ࣁ�G��	��Ў`��2q��D${�OS2�\�qx��5!4��I�	:�\��U��q�Gr�tʵv���m����-Xj^�+�6YT?�	�}��,33�.�םe����̝��Y�v��Ԣo`[�϶l�U?�l���`И���[M*��;kƏƊ5�q��h �0��r[F�@E����,�ሒq����"=wd���@Q��k�+9k����X]�쏌1�h;�
Om���Z��(��=�l[��z8�l���taP�i�[�M!0/���6r-Om�6���&��-�(Qä^�q	c1��o��qߞA�x37�_uTk%�������.�o�Aұ�Z�H�
��1IV)Ǆ���E ��ڹ�:��P2�6F4I������a͞R�Vs20��Q��f�w��e7�L��J�.�oa���'�U���!�Wt�O@^`�W�u��m����M�21�܀�����B]'�ԣ=u�|��n��;��gI:"��C,�U&)&bO嫛��Bm�Kږ�,�� �\�$�1��XVt�N�a��� ��t��#��� ��o�I�'t�ȼ⧳}�Bhd�)����ٜ&�ߩ�T���f����� �#�y�E��bRp��6rD^~�s���j��KN��hD�X��G�㱫T�x�9԰2�a�����Z��_��H���)�e:���[�d�+���/��DQ<�I�
��
��4k#f�kJ"��ӏ�c -o:�9%�9O��б���/�%skR��r!� �P{��^�Y��v/0�o6vj����W�HB4�9��Maͨ�sl����zK�0~:Pl�f/��Y�F�,EY�J(���W9������rC�;��LQf�;}ژ�! 9i2�7�\'�?=" " +��z"о�N���[{��7 U��zz�����t1�������xQ�%�t��>��P!��9�[�Piޜ�N$�܀Mr�Fқe/�Ԉ���S��Rt��P}����_�߁��
�s�	j;�Ul��E8��-�
�d�Yf��y�lZ����GI�S�X勎HǴ��V9NЕD���H �$3���76�5x��D.Ȋ͚h���k{��A����qӔ���qC˕CHO�y���k�С��Fi�iұ�O�^�M*J���'aaF�k����z%���d���4n_�K'i0�5����ҡ*�I���ݮv�y��������vs���7g"t�]]]�+gz���tЉju��m]��!�]^���Q��<=�W`�b��Z�0��>]^�G��^���V���X/�+�f�:#q�bD���p�=i?�t�	:n�ٮPl�j��r-�`UA��ҿM���\f������!� ���j�5��gšu}�*��ǒi���W�~�S�_��,n5�8�N�m�]�;N=�wf�rh]���]��-��*��r���O���QRH���O��t��Ji�vL�J����$7�m��m�:��;���%�D�̆>�F�.�NE����F\`7���k��+���\���b�D�@F)��.-�D��B^Z_m�г�A�ҫ���H�u]o����\Kh�G�^� s��ґ�Sd��nJ$P��H�P�_�B�x
��8F&v���	�'��hk6��Tc0�!0;oK�/�܀�"/y)?$��%8O5������Ʈ�2;�462� i⡮$���,��P8�~�ZҚo3��D�n���^�V�76��~8�	��p����E^T�5~�R���g�eP�R���
�'Qb��u8=��e�1��{���{T/�)\���t�;��doaS#�pj^����N�Mr�{��Q��d��:�ح�*�ͭ��kw6� wo����驂>7v��׹(X�o��\�g8�)���D����T���^z1��}@���%�B¨����(���'�#N�>��cGr�K�G�/����H&������.�<\�p0��pøG�*������z1�y�P�Y����>J����/Sd�<���1���Л2�:r�XZ]x��R{�/���+o�]৓0o��'B�>���ǁ���9n)��7��b��<_h&�5��L|��$���x�?dV�%������F?�Z
�K˩s�4���Ц�\�5�$Ǔ�Z�cQ���@��Lf�KA�"Ȗ5�����+Fi��T��u�e�:︼���f�*O~Ja�s0W;!��iYqc�h��ƴ����D�pR��I٪�q9��]�|��Ve�������_��KN3⭵�#y��n�>��;�9ET� <Jt�����̦��+k�0&H��8P�.����]��o?��N�[�����"��x�ȵ�U޳��q� �!S7�SCL��I�+P�4ZHh/�E�檀Dv�W�h��L����i�ѩ���<.��\���S4L�|F�礞��d,��K�D+
x�}z?`a��o.���N=����ٝ���5�5��dr�E�8:�O�k��:��c�f��wL��7L%{��K	�J����m���v5��^��h�@�n���Ծ=ƥ��X�
|9�9����{���f`W!�G���C)��Tً��[�x�l*9��|j G����bOTm��$l�UF%�F_��:*
�7`y��፬�FNT9H�WKjh)Z�,8���l��Ob������'���ĕ��t��G_�[Y��f�h���<%�E?L~}� �:c�9>��r�s��~�3些�]�M�=a�����i9����eVZ�'��*�Sȉѫ2������]��A$,1)Mƴ�F��!̦�R�C��8uȌ��m�I��'��F"~R|��H�ㇾf8¼'�_�C��1����U[��w��T[&�p���Q�_��%��\M�Lh&.e��S�eմ���غ�3���J4�cŵ�^�j���xmV԰���1�f��Q�U�Io\�& Hl�P)��6H�Ґ��r[�i%s���T�ӫ���)��φr��e�����Ȫe�'�lm䩱���[��J	�&�U9�o���\F�"�"�UG���˚r��N��:F��!7�a��*�1s]l�s���.o@m�W�m�ϼ�w�Q�����+�S�Y���I��.ct��O|d�A��nO��Q�����Ч<�WE�ZZ�%��7{D�K}�O�`�Y��α�Ե�ڰ�pk��d��:c�kq�w�5l`��8靦����X�Аe�h��lJ,�z����yGH8��ʲ�P�{"�9�iO����&��\_*I�5���V�����R1K�$}�w�� O�(��665(���oB����� �L����or�Їdj.���S5�XgɷI��J R������עH�W-��I��lO2���1�pB�p�fV��	�4!o��ѩo���%�����~ʮ�d~j�����$+vN�lx�v�q6#w8�&�ʎ��R��y������׀�7�x�@�y�q)l(����Gk(�z܃A��z�	"_�"�a�Ӽ��� ~?Ƶ�桪�@A���B(�N��Y	������ϕ��� ����U�Ya�j|�Qʣq$h���C��)�.@���|�X�ݛ�l�uP��蝗��۔\�_7�x�g{��([&d|�[{���=�7j�y��T��L.4����Ӕ�L@Y�ԭru���go�X���/�$�ц�['Q�΢HR��g}Ȩ�#�ý~��X�A��2~LI^��p��8�����t(�D�u�B��H�����e���f�[�D��p�W�)
��_@z����V��g5��G(w]sb��Hr�����ݎ��O��!cN�c�Y���'�p��/�褽��b�S��S�g\;�����'�� � �Iһ���-q���cyu(�QNӦ&��h�|��\Gp��;2�Rˤ���V9�n���#�lo�$�J���ڶ�`^�
1-���xy��m���)cO������,̛��V�����uU��O�J�T&��.�
��0�@,��U��h�a�ǆ%�b"%�q�����	����*�h�k����\̞��Y���q/�<U�%��#1$&1��!�A}�ٛ�u�a�b��3���bd��L����;S��l�8-:2�*r�\�+�v"��Mc�
�.��G'	���v���.�Cδ��Ĩ���Rm�8 s"?�r)w�f�R�´͢CMneqxY7>��i�j�Oz�4u��0�7�$x�.�9��G�}R��f+���;�?�̔�5x�\��oG�(
O��u=�`1J������s�>/3M�8�Tm��O�'q��f��8w���-�<Ec���\a`�*���a@+�=�Nn��.�0RUO2p�\�ҳ�=���և쌏^�[~�?�Ќl�-=U�6�(?e�2{�h�vft�NT��0b�@4���1�R�J0�5��:�/s�b����RJ ���F��!�C_Ps��e�81Fk��t�|R����얏{T3]e��h�*>("��{���O8�R+};��ե({��L߮�F+VY<����]MR�c��MZ�7W2YK��`k���>)\�ܖ�m���M�ә�F܋׷1����ܷ�{6W_[#��F�A��J{<	4��)0n�����3�:K���k���js��˜��c��D�����&�\\q���4�����vB�'���(�2��6����3�3�`(�]d�l���N_�jA�q�{
ƹ�E��*-%_�?�W�>C�g��VLqpí��O���F���6+��+F,��[��ۻ���Z@�<7U��~������}@��N�C��=0���Ҝ{�'�����9R�{��������`�K��x�oK\k�[�Z��*��� 3~���`�4	c��ֹl�C�
�|�r�Q��؈-c[B/N�M�ۼ�` ��ZP�������1�����yڶ[� p�<-[s�TAc#f������4���n�ﾼ�ž{�@c��))EZM_��,�]�mr�7)�^@�U-���0n�;؛F�����H��/dG^�kZm�~���#�	���N3�)=�B����>P6��O �l*�I��:�_k:vMj|�km_z�HZo�
l�$��.�a��𗄣hP�7��G�)��mjB�#,����n(��>�u`����1 �X�������X4~(F-D�]@!��:9Nw*!��jb�s3H̯i2�^;���B��c�X=�[x��mĒ���'=P�ۧS `rGE����Z���s��v��~��Qьx)���ڐU�4�_�9_��<d�	�
��A�*{x#� �%�:��3�����c�N�4�σ���˲Ύ.��h[�͏��%���UW>��p
�j�	t���q<Ru�$Vﺛ����?�1z�-���e��]@��"t{T*��e��M@<�ܣ
)c��:����;�(�}�Z©W���߁�?[Ҡ���4����`:P�ީ߶��I/��}vzk���}Nf�l������R�#��o��#M�@��X}U>���l��0;�j]Xh��)2���A�V�ol�6}5��
�I%�k��d"����	}���Ѫ�ygcXTBLS��(�����`T���`��=�g|6k�ݾ�h��hU��O���X�����w@w^�%�fd:*�]E�:~��G��W4l0��ĮƔ��_��$����!@w�(�*��T��V
�u)��$�ûC��5���Y�C��<�C��(��ST�VV�f�Ow���<�Ծ��@�An���O~=2��S���5�$j�4�ͬ�{-��m�O�H	RF�$��j޴��8xm;k�ja/RY/�-�3(��M�Rء�;�{R�L��Ne��[�L�B����Y|��9Hd��z�h&C�6o�W�U�V�����u�
���ս����-�Ǧ����@=���,��|��1��,PK��<԰�; �aӛ��`Vq*���d�=���#nh��{qe@��e��Jt�T:��3����!��i��I(����WD����I��e��5����t ���_�C�@$M�I��8�la.�cG>��z>	�������܃�n���
m5����� ���[`;������qX�4���x�O�.?*]a �_Q(�;��,D6ޞ�ȘWRV>��'���Ժ���nr_)��֍�7�e�mCdP`Lw&�=�oM�м�5��v���wcT����_�I�����^�jǙ�O2��t+5��3�q	���+�����e��9�WX������gv}�}�� �x�RN��Rޱ�a1}R̄��{⺠	S�̐����as�}[&)r�H��(m��n���H��k&�F�0[����XDT�(�A��w�I�+�5t���4YϢys���<�z��4�)�eR����1U&5��hy��a���6�379^L���?��l@����f�{�^���^��f��2Zb��_Tު��6θ>ߐ��.!�M 3��u��_z"3}h�Fw�̛R��X���b���N�6�:��b��2�[ö��T� I=�pL/}ҁ����9���uMN>N�ǁ�Cs��8��--~ᶱ�M1�?�ǌ�H���˘�0�IG��3���g��cj*rL�Y3�l9�uw���� �U%`
Hi�}N\;gg�@0ၴ:�I�J����.�}�RW��k�9]z�6����h#�ϗ�����yѥZ��< ��n>;'�c+)M+���.�m���;�k�4G��uxљ���Yy+����I���/�����.q;)�� N�00{�����Х�nV�>�b�JWég8 �͖����7�²���5��nZ��8�M�H�*���q*RN�9�e3�<�s�G�"����WC���&q��{�^/HIEǛ/���ד�F�E��d�����Rrgx���QWX"�;狭0�s����Q;/�ep&�k�4( �lR�2������dD�(�j �-��7�I�kzjf`��������.�t�IS/.S����ґ���A?�A�/|^�&  i�R%cq��I��N����j=��d�Q�v��Ε�
���ntQQ�K�f��k}�w�>QC#���o>���U�
�����SCaa����m��#Q�h5'�X��z��������Ł/3��8Oc'R�8�3 a���� �hϬ�h�DVρ.�Q�0��Gq�]^���(LL,���'*&��`#�W�\��B8`�_�T Rd3�Ʀ��ꩉ�q�D6S5c�iajs,'#�Tb<[�p��!��b&;-��v��4w �W�S9^�կ��[Q�I��6k'\��'&�D�`-�E,���