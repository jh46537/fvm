��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK��i�vwrU�j��}ϵ��t"��8�-�x�@��2���t
c5��j�р���������\�"ԩ4k"����u%%Ze������i��p��.�kE|���3��s�Y��yv\Ϋ�"�"�[eJ6�Sx�W3��mZ�v�;(����u]QgK?Uv��[���6��(s:��ii�#.�r����g��K(3�
�;�e@H�0�c�V��,h��m:���f�HR�^$����q���_+}�|��7׷f���a��JS�����`ܟ��o��B�N�c��T�"V���V��yJ��('5�Q������r�E���b��N$���_3͋�WP�Ф��=٪���i�L�Eie~[X����-�梐�3���\Y��4h�M��{o���R�ɇ�=�����/�B�x�yh�+�����[~s,1����C2C $��\�#��(Lq��z<0�pWs�-=�4PH�B�$Vj��s��ٲ-k�<�B���K�,�$ظ`�S+���� �p�`�կh��BÎ��S�MU�2�2��ҕk��j^��)+~������p��à,"}S4#&Ý¸��U\׋�P�N���-"��Qta'ճ������^(#�mf�<��i�%���M��D�����)ua��g�>q����"�C9�Q�@���m�a,~�o���2>:MS�i�-^�U-�T�϶5��A���AjBC�R+Y �%Bj��f�{���.�
��,�#��F�����,�Ǚ;*w:Qm;�k�6�?�(o���.2<���8�<�O�LhMGl�ͯj��d�)��|A�=���۸F��T���T��׼?��x�������)3����{Ӊ>��	$�q������3'�E.�6�#�����z����ib2��l�:DZ�&����m���l}%�"u���V�观���UA�`�zhq^��S�e���5�Y��q�q�8�jA��`���o?�s�=�h׾���A刌��Y[���^���R����G��Y���#��3$�I���$�?ڛr��������P��qoƓ�E�5�r����ފ��}�$Ɖ�1'�
I�%HR͚M�"`��JA��k��(�B�ls��Y�1�m�����;&����)V{����Lyp��/�b�[�]���
47���^�r�_��j��b��g��P�Y��k���7V�gO� 淅��DjF��d�׻�4At�@F��玖n�3�.�<p(S�5(����`�������:j���ʚ�N����+5+�|<LE���D"�C��M�}�>���"f����m/�WS�܀�S�������8��Q Moc��c���ִo�<[��㾳�e�#U�qZ�L�ȿu�� 3�psR����Åg5��K��^�#C�N['f�(J:N\���M#��鯖%�gCȖ�>�� ^��2ʓ�W��!��oŹ�,H��vE���C����lb�>��eu����
���{�bshȬ91�d�!8�B�2I�Tm�?_L�J(���Ms�h|QQ"KN�M�Zس��&s��]�W$��@<�	v�����&=�4B�E^%)S7��0���҃~�}霆���X�YWo�k�Usf�%��3�!��Қ=��(f3w��wW\��x���@nRt
��V6����3�l��e-tk��=��ۊ�\����[�H􏏔��l"v��i2eI/����-Q��!�����sZ��b
������tu2B�0��9(&@�Y����ٌۛ��lY��9�H6�mF�nO`v��������[py]?]>~�3��3XՋ@�fK�^���Cc�LR���
 �^�᮰����r��ov�r�I�mj��V��Ҟ���c�^J��0�(a��4H�0��r�WDm�6E����'����aw�%�*y5\
W}�쉄��� �I&�Y�NGPq"&C����4;s?��2�2sޖwҢ��N����mZ�ws?T��,C�Z��t�̑�_����K�^��
����h�.f��X'�%�SB	zEm
���b�gu�������y�`�������J0�R�Ḫ�N܇���;��Mr�;�P�㵗�ԝ�a�epM��~fh�	�s]E-%�g6؞�s���6��R[�����f�P�oP&��l�~Cг�zu��@l{P!o��(E�>��������zc�U��3v�(Uk�`t�� 턉�����|eF���D�`u�1`�.]y�л�'9qg���V���^b툮̲�mU C1�ن�*mk�kxր�qJ����a�-�>�ݒb��ʶv���J^�]���{��fQ�תڱny��ЯL�s[�Fy�l��7�8�L��l���)�źZ]�~8�R�zF݉�'�n��0��4�(OF�*=}Q�/�ej�R}ڌN���a���`+����/N<�5����M/�5��M%Gq���bK�
t��UԊ:��F𶰹0��d���E��(��(��ܞ�����!=��"�&��bZ�"�saXr�n�&��D��9�]�)�t�w �P�Z��������@P��*�o����Ƞe~k���k��05�p���.O[^I��R���\`���Ы"ɠ���m��� 8��~��l�R+��-eC|��i��H��1K�ּ��ٶ̈��&޹�B�tq���;��<�Gh���ޑ�Q��S��5�;��������"��6m[|W8�K�V�U�g��E�=��8�Q���Q*�x�!��E�$��������"�Q��*��`;�q�n:v&M�W�N�Qw�7.n+B����UlQ�V�nm2�c�>v��:� [ 7��z��	�����MZ��Jf�����W����m���p�a���p�~�3��>��Tp*6��2��ե�Ҕ�Ub�Lш��N }�����@E�a�pc��م�9Vq6x����z\8�V����Ʌ�7Ѥ�氄�9,�l��'<���t�d�f�De���1��EA�p�l\�Z��ѿ-_:}o˺)�=��PUӨK
�	Z*���y
���5*U��y��e/ޫ�D���@�.`Ņ2���]��_DC�w�2�76[�~���Lxl�Q�	��3�4c�^��ƿޯ�rG�I�9̓���C��p����<[(NfH�a���ˌ���88~u��l�C�ff9� 9{��M���Fxu���qjUҭ�7��J�!�MJ�����z2ь�3ߢ����]5)>"�0�:�ߥ�Mcv����6-@�H�0b|&u��ŝ
n�C"���-Sr��'gɚ]û!3g1��6?�0��eߔ�+AÔ��Gzg�(/�aw2���|l.b���Zߏ�H��4���C�K�m��_����H~�z��7��tV_�r�?0���'�ي�F %[�*1k+FU�S�D�XeV�٥��X+�b�B�k��_�d������IT���ƍ.V�#�FG���"��t	�����S��BUZ\9�-�xL�ȞG��7���&x�����>jO,Ż�=�V�b�t�8Zx:���aL�����l�1�6-��?����WK-#=��O?��E$���4���,%�Cq�գ�À/�B
l��}��ө}���2T F�/��0i�i,3k�a�@
0{ �-��;�ɅJ��	R����#D�9E������u�ֈ�M�4X�������E�,1�.�E���
� x�d�ʩE�<s�Zw�o�+�eO�)��8��bc M^*>�dp�@�u*̝mK�`tq�K$��ȳd����>�E6'�������6�:Y���I<��=�lj�y	>����f��7��a�-3����F�O9a���Ǧ���}��Y9���n��6����/&D�k�%��>׳ޠYK:f���بF�I�w���fJ@���W�Z�(#��^�_X����1R�eQ6�=in�'�LO�u��CD���Q��$�RcS̶( �I���<Es���z���V�\@g�C~���Y �11���=�@�]�1�qset���hIr(���@�Q䤛��T��ޅ/��9i�}���F���s�~�lϙ�/gJx/#M���0+�شCǿ}4�l��^�w��`�5���}Bˬ�"�!-�#%���n�}�.����<�Y�JN5ٴy���ӝ��PW�Z�W�A(�`ԅI��]i'���71�iEU�+��9�S�P�i�EՌ�6`\p>z���We_�rs�nǄ��SUST�;V���Aq5x��ͬ���8P���s�Ѷ���3EΞ��f=����5�SvxO���Y���嶮ֽ0$�M��Ԩ ����2�X�2����ԪIE��7}�~��+��*py^)_L^�Of[��'�np{�G��`xЂ�G�S8�s�`cW��H��o�N"��!���y���`T�xa�U�)aE0��R��pe�T�$A)�C������y���@�+:eWz���c�,>h���%��fB)wgT�)p�ݐgr��.�Jk���Y����9�ڇc�o�t�����@��g�t�k?S�_�X'W�Z�m�����Dڍ�]sq����s�xC�X�l���&����rs⚧�G����� �����Cd���#��=]k\G��0+��@�ۨT�x�vP�\�߀ƅ�te��F�{��7�,HVHl�n�uж3ژu�K���>�)9A��Q��)�7Md=���,�,�TF��TG� �� s���y�w��"׆a�L�p9��3�

w����or�6�6�75��i���ø�\��	�&&�G�;��gSBPB��;�#(��HC<u�x.��+m� T�S�rl�M�{��3{�#/A\�߈��B�~���4��}Ki9�ϱd��T���������{9R���$��~�2�o��\̪��Eh�w��Q�F�=���؏�����`+(,���p���&�xNOK����;���Q�kxd��-j����ٙ�<��$����qՆQ�"(m�_���t�F�_��>���Y�H���:�����Ƃc���S{�>�^�!��e]���u���bD�G��{��v��h.x@�,��RqVG����۱��=�QIzSR��Ĩ�oi�|Xn��X��TÎ�h�M�|������L+��V�}�R}:�s��:t~y�w�sPO�\�XJd�g�Yl�6��sJ�C���+2�5�����>�,��2�	�!ӌȂ'"�~�.��2}�$̓h�����L �Ae�3���YR9q��&��I(Q���28>�M�ۢ�����Ԣ��L ?_t�� q� �0$7�a��l_+$|���V��.�z��0�`��F�l4!ѯ���yD�/]*��"挄��ޣ����r�D"�6� cQ�[�1�]�z+_��<[E>��fo:ȑ��)�	�}m���4�8�䧊������E��{gp��Ӳ��"��\�x2�:�9�Vu?��Y/c,렴�/ ���^H}��(K�Pj�Z31�Ɯ�K�J�&J��!�����tSZ��fsg#�D� �n�@"�[p~���`{_�����쬚�8���]LE�}��ŨhV�m��a�q�b!R�l2X�]��t�|c����KH:���D�����	�hN��0r:9��r%l~�F<XV�u�Y��80��2|y���4d.�|rD��!�{�*]χ�� Ex��`4A#(���RG������v�ՇU�F3���Il����<�
`��(�� �؏d��V!rX�����c�m�����ב����Î�iI؄�W��ɩ�8#n���+x�o$����������U^7i4>�G�<�7뤥1|�q]�ϥ�Zu�d^z�u�h�@?�Dc��y��4��]��tJ'0����$ǣz9̪����*��T
 ��-)@]B6AɼU)@
CME6��@A�����cY�1��l^ɤ��F����5rdh�Ƀ�plYf~����j]�
���ͩ���L
0��f��1���spz��(��0櫛Rʥ��k0ާ�²c`�S� �`)�w=�D�@��+h�+
�V�����z���R���z��}�tQey�t���tf0���/D�G�ܹ�P��{�̴�����X��E�6l�|C}UϬ���7�(y3ʍ�NBZIi�{Ddid]_�%�|b*5���2D8P�0�V0�:�2��]�ۺ��W�a�6%2��炳G�{��XĤA��54���L���TO������Z� �7�:��`�?㻿 �hً�ɖ)�������}>�yA��LTn�_���c����*������cr���Ӻ��1�4P�%�y\`��LUm���ɐi,d��9y _�TGZ�M%��.U��	�;A��T��	8i�#�Yf��0-�1���+U��$���:�z a����J���b��t�S�!�7m@*,vg��\�n�܊a���ƶ�j�c	��d��o'e�H���]F9�\z����|���s�+�
�����_.�? ����aH2�`CX&F	�(g�F}��V�ui;�Y��������Q5Be�Jo�>��p���)Lek�8!`�RP)��'!b�߬�l¸z΄:���{�O��&�b��5">�����R����ȓ�DM?i� m�Z���9�~�Ԫ
2Y�'�H(+Q�f~#���gpd�B���0�+�A��i�%�Tƻ�(e���&�¶l�քE=G����A�J��2�#ޭCJ��>���7�WU��=�(���*�ޑ��B۟9�>�����Ŀ�rlc�m�G����"���U�IBn8r9��l���2�.*#��` �!f�b�h��Я�1���$wRJY�Vi�����~��,��f�ύ��*&q�PI�/�%_v0���It�K�ō�z7�(���q0*�z��;����a ϼ3Uv���Q #�����ݙ;!oO��y�׮ަ�c�L�	��^}Ru �a.|�i��.��<���o��c��>gn/�<�4�|Uӌ�3�e6��V�s��B��0_�t��Z��&͌95�"��d���ӿ�����)���
�X!	w����M�`���q�����uη��焦o�����p1��"��ȧ�W��.\�]_;����Ay	���܍��gɚ9�D52E�C��O���<Uݻ!����T3���Пɥ��f��pk`�c�(��߅�+�\y*3�*]�t�Z���-'�hN4:�n,9p�����\�m��^L�������r�%��D;$M��Ӥ)&5ۈ%Z*��?��Ë͟�I��/�H�D�VK̫噎X�l+�7e±������T��vM=��6+6���Q��hЄe��.��WL̆��sfn�ю=m����
��x,+N"t�t���Cv�/��t�Ό �a�O`��������\%�����<��)}�|��]���&�)��~7Hm#?�$j�uE�ݸ���?����')�if �6[/��a{�q���AN���)8�O�(�^58��{�"�k�@�ax,�V�o/Q�ޗk
���>�uF�{������ߍh��'AM6_E��[�ǧ��6?:����H+��3wN�y"��~!��ڿ5�t>��Ɔ�;�JQ5D�=}�օ��p<������~�s��&��Qyc@!�V˾O8�f�w���QkaNm�K�K�ƞ��)H"�`&E��`��m�{�4��Oj��M<���^��E��PzI�}�ߜ4`{[�q�~�����p����d��М�S�����"�^ ��O�|����<��b)�KT��4u�>u��Ǣ�&�!U;hL� �y�&�9�6������A��]a^���-��^�Sn%p����c4����r)��,��.�H�M�-̃��˧�(S(��C�
���l�+!L���B��Hs��͢��r���R&~�׍�K�,�^�-����]�C�����IR��0���pn����FGʌMD��6�R�r�9c\]0��X,�˶�t�a��g�������9{�&? �~�"�R����ѡ�xjx���8v�2_p�Pw9'3�4�?	7rT:�{���b"�MR����n5��C�8�|�
!��
� �E~"��50}�՞�8]h�y��!w0[�
�,oA!��@�船�7���5�y�C�J�j�C�dB��$2R>;$��zX�)��L}��&��H�%����]���g��d�ڷ��o~�)Ɂ�h��3�I�-,�~; j����:�YbZO���K��������ݿ�~j��{b��9���o��D�CM���t��<O�p�F�8�u�2z�����JpA���E������1^��	�[	��8��o�1�tBqz�F0���֠����z�ź"T(FDq'?aؠA���}�yf0w���F}!�~SJC�:w��7�CO�f��]��IS\���ذ^DN� �&_LeF�,�,���1�ЭP�Jj�tPTB�%���|�yu vBb��v-��*�R�ߺ�T�)d

V[�J�ã*�|���gJR���V�c]��,����
�?��F@"FU�M��'y����1��f;b��g��ˁ�6��*#�o\ⴅ\B}�
E+�}Pu�T6!*�(�i`��Tb)�e�F�T���B#''�D����S�h��]���Ʌd����a[:�.�0�^���������b�+|�0a*��_H�}��%��-h�#�zJB|2)eҦ������]�|�ZB���w�k%T��П�A�e�1N�7�X+1�a���-���ir��f�Aۏ��gf���Fꀗ�=7�욉;�h]�sf㰀Bжa�b�H�5m\��'}�G�����3���+8��.NE�#}�O��v�B�OJ͹����wa!r�ka͍�b�z~is߾_߬��'�����kr����jِ"[<�>��(}����+�˱X�F|���l�mʷ8�����P�KTŔL�"U�y0W9�½��rV��j;��#�B��P��NI��O��c'"�,�������iv��R%7m{q�4�jb�mue� ���jzX�M��iTr�H��8���>o���t<y�u�Fk\`�t�?��#��I�h������[kvjE /� ��2,|:ްt�b��8�^OXk�i����[���$��缟.+��A��܍�A���m�V%}�I&F���o���Ř�,�\)��4��͜.��̎�sȶ�  �^�o�X��~뾻�s��&������j����6w��ly�+��R�-��@ŦR}k���"����Þ�#x�׋�!�E���@2 ��=��2�A�.ȹ�������E��Gi�*1�Ad��4�u���)|�e����9wV`���E��w�6iBD��N";F2��ꮒnJQ���[���G7ں|؏����K^�@-T�Q��q���<&��C��|
ӑJ5)
l��ϗCdC�J���30^��e�lWVQ��d�{�����/	v|�����=�B^�܀i�� ��M1���P�$�i4& U�l�ұ���[�R�W�A.Q{�=hȃvfȠ^�=�T%ն��R�x�8�,�n�;N=@v��<�#�G�� �a���=}��#6�#��gn8'j_�Iw�y6�}�+���e�Ρ&�:d���;<(w\�:-���$����UIԛ7�د/�Z���Xw�,;�L- Z�8��d�9e�B�+ [���� l�{�x�~L@n2{J�t��"�]陸�S�&� �ň\:�&�)6�i0�㊘�pa:�l��V����a��F��~�O�K�f&��J��̗`3�W�0��4f��~i�;uζ�
�����ӭ�(\�z�y[2�cr���&���w�_�F�̄.G���R���g�y��;��6�Ks�ydC�q����ך�VU"��?�:�탌Z���}�G���f�a���Jk�q�e޾�!v��W��~ B|���0����F%���\��� ^���M� �t7�C��'��!�܋{����E�:�X��w"U�G������Qis"y��ܫe0m l	3���ue�
?x�ոnH7�LT]���0�(�}����?pA�z�դ�z��IJ��_�S�x�8���h_��a%k�,��F>k��p��+���Y&ȃڬ}n�-���}��i�"��+ራ�VfS��e�E��!��qz�#$,���v(}����<�j�>���]�X-�wx��0��9�8$�2�mO{���T��"u�~��-�[�A���
���Q���#�u��}��`�D{�����B,�q�p��'����Uϯ�[	��t����*�[��c��Y���q�N�,z�1<J��砩�7�P8�5H������&�bi�Db�Qz��D��I��;�Goi�1�,`d,��R��`Y�Y��A�ȜȌC��[z�V�m��ZI�s������6����bI~�X[���P��R�s��	���,
�i]�Ҁ~�!n����v�~�_Xoշj�y�������u^%{��(���A�u�-���x��(�y�k�~v�`�'�n�A��s�6��q�ث��yϛ��C��Q@������P�T���]��<e��2p��b:��(b�����|דF��*�>�j��V��-��f�^���Ӥ�#^� ��1ѯ��u(�/�ByC������'�@�H>� \4F'�H��9�s�J~��m��L����.'��g]�?�R�{����E��3����Tu��
�*N�萛6������TS��z/	���@�h����pYjK��6o��u^��o9����}��.�cyh�'�цx,r��W�pK��˻��7�ex>���!���'RjO�$�Rlg�nI���T��\>��$���������u����9n��禦K^:���Y��m�L�g;$����7�!�l�hm������~�W}��n�hkt�It:I�y�������V�����S��2���W.�~C�5]0�x��t��?�7݄	�+s$>���qZ�Yu|1
��4g	��Y����d��0� 8p���G|�~�������˼)�7�#����Ԑ��\�Lx�I5������"��|���I(��ӫ��ı:�_�4��]!�:j%�^���=��@j�D��+�D�zAгM_e�X ">:P�|Kh�V+nEn��'���vs�/��`+�[�.4��L��gI���~���4�D��|��1ײ��YU�[
p$蘭��EE�]����@���1�xE�E�ܾ���9�5�1�kH��D�:�D����]���}�s6�����R���dE�zhgG��1L��	v����2O��!�u�{|�%CC����?�n�z� �ka/�������#�=��HO�V7s�-���h=�z�R~�b4��xE�ɔQ�5� wx��}X%>ǒ��
8�)�-�1^�^����dZn��UĨ?OA�濌~��ۘ
U��h_�����/��\D����JrU鏇�s��C����B����S�cرǶދ!��Bg��6�!�Y��э��\S�7L {t��������ff`y�i$w���!�6ܩ��ՙ�Ffq��J�h����y�MbdB��(y:��,:҂��	<���T�Z����a����d��,^�VR¶6���]u-&�c�XUTeK9B�I�~�]�B!zh��;7aENB|��`��DV\���iQ	�X�~�� H��SC�[��[�z�����~(�}�zhb��S!ö
my�U�-[�V�28	@I��Ą����L/�W��X����\z����?AX�c"i�'�C@�1/�fB��D��*܎�qu"j�.IM�͑ѐ��p�^-�[�P��0x;��,B�'�tГ9�x��J�0��=ѭ�N�P���T��ꀧ�{��#�sV�o����wP���	V�e��6�rw4��Ԁ��X?Ϲ�}��)�YM§}�	�_���6/�����K��3��y���j��mRR2+�,Hѩ�M�Y�����W,%�Z�U�N��V�ĸ�Z��`�8H�5�8�R̜O�bW(�����9-_�`���_����Z7_�*#Ƈ�K��2�Kޢ�5�Ǒ �k�X\բ�����u`g}�R�du��H��L�����-��?�2qУ�^Xo��F7��W�����,��&o�W������ T�E���(4:QU�E�zA�78�Wк���q�XTd�1���0�]=��xm�x{dN�?~�Ax���D�&}�x����UL��A8_ oJ�B%9��Px%��2��0��`������s�-3��	�!-
<���뢊�Ѽ�X�1L�l%��x�o(b�3@��'_j!,*
:����X��Ԅ�.��&�(�Ri���X�I�ޥ��V*O8m�6�\��\�BS��m?��1@��ru'x��@�Y`M����%���<^�R�\H���mK�J�YL�	TGk�k��g�|��72M�� ������Fx�ŧ��=E�2���ƈ�2L�+xy��z�Z�2�iNJ�H�?v�T��+�7���^���O��Ƭ���1����τأ�V�;`c)�|J� �4 nZ�ӆ::�g�1N�&�/}w�sG��+��&�h��@�2c���mG��f��"�jB��
"Tu z6T�4yGk;�d1�����T�����N�����y�+K��5�� @/�{��Zw���I�er���L��d%�V�Ν�~)��2�^��j`v��EF�Wػ���3S�c�;�J�<�}�qtV����Q�����'�^M������mV|'���	af&���Zf�0}��C��:w�1a4�)�DL�y ���#ڜ��� ��x50q�SqC::n��/�������5�m�\۴ �m��qe�w�+�(�z̲���gy&� �G� 4�c�]�Z�UM�	��i[ڂ��q�����yS���=F��8w�C[H���We{p�I/��a+��y
e����/7��T�m�rvAi[��d��G{����y�Q
�� ��|�w9���K��P����R_������9�w6�416{���@w���g��c��QL+�ʃ���
L�����@wI����L��c��m}������=lnӪӛ�(�����K֦Nأ�|�s��T|�CO.@gd.�6�
�������0���}9�D����4���I׸��>��t, Brx��bs����>�/"_�h&�]���꿹̨I�bK:������7��{�ܱ�T���&��*�3P�%�o�2p��Mv5j��(��t�%�w��)��ADkU~�dz�1���:x�n�� ���&��?E�'�Z'T�oyo�e�۬%-�Y# qU�����Y����<��f�i�Z�[�\�Ŀ'庮����/�5�Z,zѼ5<��	LA��Q�D_�|����/�!��iD)�q$�0���3�TWi�" �՞�����#�wf����#[��P�l��E�:C��\3�y� u|���Mw-�5�D%����~�H%?DJl9�=�3�0M\�ʡ�1��J��(��j"^��^��� ���&/M��8��3�w��Y��>�6��Ʊ�g��TI�i�����s9˟���P�Gk�r��B(�ό��ƴ�q*����k�{. ���z�Z�g���k_�l)V趨kd`�S�s\���dh س��CYΈ��o�PG�r�ƦP��?�K�7Z+R�d�b��b�D)�5?o='d(厨Is�3�t���[}�'ں�	��@�y/���,���Y|fl	���VEZ�\qM3��z��՘�h��EDG�u(�.-�����&�oȒ�]6B�_-8��yQs|�@?�
<��D��bC:���eՐ0jiL�z�TU�!�\�/J=���<��0g8Y�E�0��{w�<��X�4�?�}�N=��E��(�za<�J.�
��z��	�KB[�	���z�?{ ��I�lI06�p���8��;�F�G�Yv�'~�[�j��J���7��:����&�t� �Pd��[�����	9�X�4�����J�d�ƨmfcfm�Y�W1�qQ�b��2Q�q{�Z��N:F������$𮬸L-3���(��V�S�)���sǉ�BU�����)Y�t�M�$��2cM��ŤxJ@ʄ#��.�<�5���]�S����JJ7��m<�p�u��R��^uhT�5澑M�j�.�o�����	����!��e�K����5�8�H�
��O|��b��q�_+�|������9`�X ]�0Z��]w�'�2�1 j��WD�"U���j]EA�|h�/�1j��G}�0��Z멢S��)���3��0g��;�'����!pE>3��GMi�Y� Hy�S˰��V}R]�r���d�����Bn{Cz$T� \��Bo޷z�����b����{����I(!�m��'H��w�D�vdع��6�xPݍr��X�m���'��
����	�qy�c՚`�[��7dv��Nb�@�u�;�5��f�-���O�E�kK��O�������'3�QV��yux��dj��n|�>�e'X������t��m��K@����l'e�f����K��$5���EU�d"i�%�mj�-䝤`��1�Ѫ���w5��ya9��@f��$,y�����fTf���k�V�GՉa@�:drvF���q7��t�V{u��Q��?������s�p��F�A�����G2�5�b�*,yd�����܁L�tW:åb�|`����3U	�J�tN��Z6;h����G2��Rv�dIي�����M��I�#*뭈ls�ē,�g �Ool�Ț�Z8�V�D
�*��2�|
�a�}��*`4tf%,��025F�R�=v�/(��[6��K�'��Nnf&;���6�mMz�
wsiO.�TQ��se@ΒY�0�1���T�� �n2)�;#+�@�t�8)앺�l:z{�$��ӺD[��7�9zL�Å�Cd(��	��[��T"����E�r��$�_�P��8�P�  ����A�Ʉ
h}Sy 6�.����/r�%(�a��S�iQq�	؆��cQr8���qSqE�������!���P͖2�[�b�G`ik����Y��+@���"@G�Tm��r~�ר��л��.���io���O������y}�T�,x��И(�q��k���:K^|���2�6FLa��MR�4���{F�Ѿ�BH���;i#�A��ɳ���3��C���EQ�so�z�@K%U���X����[i]��
T��c� ��e;"z�j>���q��y9(�F�B>�τт-��g�Ka������=yk�GV^T5�j�����}�瘑L��@#���&.F���;�mĤ�*]~U�a$ٗ�5�Kb���	�=�K�����u��O�<F��<* �sÓ���tN~8��N*�똹�i��G��ۇ�(E�ۺ��#������h51D���/"��{.
��@;C�){`ji[60Zڝ�TzJ*4�P�O]��	�G���(B�ݫav����\;�ñ����Ɂ�f��̉�����y@Q)C]솒(?hJ�b�jv��<W����07��c$�r��U�l��@t�=�!}H{������L����g���M�}呱�c7�eǫ�u�*�j��yw�u)˓c㌓������3�U> �V�?v�&Q&�캰�O�Ϟb�W\����W,u���Jt�'�n[��R�pw�*O���V]m#�B99-��1��=������'�C�&~I"���-�U��¼7x�nõ$"$@�(�[�F�5�"��tUT�mT�d>�ҩ���S��L9�sa�@�^�k���/����;���J��
G�ZE\�psꕝs�S��i��BĮ �;籭գ!�[�CF�����{�nr}��J��8$ȵn-���m=����,$���WO��
\iB���hoG��9(Eو��s�Y�IenP����L����j��	�Nf�t8X��m����J�G4"����k[�z���)�:c�^W�|n�=�~+M��Uj{��<��W�NGD���������"g�I뀇eRy8�Kv���
�C��������r?�:�� O'�3�O-M����Be<��mo�=�����7�gUfr� �*,?_�����w�iԣ��nh�����+�%�^�݆���͵��Hq8�>�c;�)hC�8xt��o�,h�gdP<.�Iw��M��~���^�nŻ�.fh2Хc��m����(��Åtc( ��Pv��e�n�a%j;З-�d����Թ��ԍ�|�r��kHL:��}F�rsS7�rdB�U���#���홚)Au�	�)v�5�`���x@4,��FD�5n$�[9eX*�Uk����?;�_0�3���N�����Wt'��d�ث�^+#��$Z��tC��axf$s��P��K���Zvt?'ep��Ȏ�n��T�a�c�o�Q?FTb}�G� ��=� Ȁ�1P�8��p���G~�Z�v!����/�uwf�Q��\%�S^;v���x�Z�{I���h����
z��玸���E�N�L!��d+R�C�P;RO���2T��t��;�cV���sG �}�ǸZ�V�"<F>hB�2�����6@=��SP,3�ч9�~���@�X �����/@���N����m�?�3|�ښ��	 m����aʩʐs���������A��;��_u?26IK���9��D��S�	k;i�BКnS�(mI�W6�q����/ ؎���Co���m`�3��Zl��G!�^	��9~E^�"���C���DA�{��r�:�Tp-Ń/ .��ʕO�]d92���O���t=3���͡��a���=r� 3YU8��ɞrT�Q��	����F̵0�&��27�'cC�N%R뚛�I��<��������-�|�w�����gTwb���\��K� _"N�:�������"�g��JVI~K#��[̞L'�+JǱ�8�׍9������"yS	˖���r�:���0��2�b�@�ދ���k.��G�N@N7��������%�~i#t�M��3��F�m�ob���n;Ar��[;D�e�m�C�$XǞ�I-��$��}a���:VM�"�Qn��M!�@JV>w����qt�'�b�o10J�۔�,�S���X�_
x%��	M�2qj$���Ь��yQcE�ף
l��8��j�lgj��o��Ẩ���?���E��K�d��D�4�Z>�:��<����U� ����R��\M��}b� �Μ[%v|�\>ZLws�Cޙ�s'��!���å��y&��<M�\V#�^ �,hO��a�'���Y��^��T^�6�a��e�0��_���(�<5���u���~���[�p�������e���f��c�%AWe!3���5b�{��$h���pAn[����o�W3{���N
اU���!�{�H7�J!��ɚI���5���?�%�P-�|�<�琤-�J�^,LwK֙Ĵ�g����<oa�E@D,��_���dx�%���JʚUb����繢�7<�
�7@*���dc{K��=��
֔[���|��m�.)[v��3��<��>�*�V{�=�8�H�̦q.�.�1�Ѿ�\6�:��;�}h����=١���;
�������7V��mKز����Ԝ��op����Xq�@4��#�A��NM���p}�<�h8J�H �ؤkbW?��v5]/f�M98Y���:c*`E+��!�̂4i^3��V��D�ۊ���¿׮���a�^����l����3|n+\�o5�>���\��K�p���-0x07ix���FZZv�����
m�������s��8_�A�*��x�˷�?����� ��V��s�ۓ�e	������]�\6 ���,q �+��'��&T�c��=Ә'AsE\nW|w��
�N�}�� ��}� Ť�w)q�3����w�2h�y���^&G�8m��c�bT�w���p��q��λ�a�n�9eɦ���+��O�����aW�s��/*�E��>��9�ѝU\��ҁT?0�V-���T��$��M����Od��byЋ�{���6>Ё˻��] �p��GvA*P�zA
��V}���{,�_��y�u��"B��ȡ�m�2Y(.��&���_�N�2�k"��`>�E�8�/���c*�=�:c0����0���Z9�%���S:(�J
k�à���~(z)ޣa@n��o�CJ/�17#����wdR�n�"�t��V�]�,>zi���L�E�E���͉��F���a�׆3S�K�WX��?,�G+r��]v*����SP�5R�,Z]>*v����K=LYN�9C�<����kn��JKo�_+�դ�b�w�߼�-�-���_H�b�5�6�n�\����u�5�k~+?�o"�O攥�T��E6shq��%�#p_�e/�l�ٮp�w׌9���K5\�{��,�a�j?�LXM������ؐҎ�4Q�sH���� ���Fe����c]\�P��^���~�@Rg�,�>�e��{��4%�`�O���U`
9������l�Yv�y��T"���i=^�]87bx���Zb���� �a����W2_���"ew��,��~I�EX�3x�mYf���׌�^y�M�9�5Պ�[�v~|�%�#L�! ���!I�-��m���e���ďXa�;����D��$��#Z��֪p��Sl9B�(���`�*l�z�F��&Q��쐰t�a���.��
�S�q	��5�8�lpB��I�
,{Ԧ�3�n0e*�/ءO���� $�EK�o��tE�"�&�SS�q�}|\sIY��e��3
v�2T�o=���|�ށ���>�6���g'�<�7��i��6:� ����뢏?Jt���wq��=��q�چ�d�CyV�)I�T�Nn�=�"�D�j[�nt�u2��\a�S���Κ>��� T$�����W�x�lc�I #�	���'4��~���9c;���{��4S����Sb	���;(��4j��W���z��,��������B
�d_�Vif�P.�6\�u5��0sÄ�[~�/ӂ.A(r�����8�-TT>ɝ�8���F3D{t����7����x~�G���=Lxs-����3�v�`� ���� �g��J�
�@(���Ff�����T!]�4��А��蘡G���!��m��[��"�&�[o
��k9��מ��)`��&L!�-=��A���'6{�lƶy�����o�&�p����~����	��1M$m+	=��5g��C���"�A2
�P��F�%V ��ߴm�Ĭ1�� M�j�C
N�#��� ��"����W�%jo���;D1����e3p xu���k4������K���KQ���!2�K6�Z|Z/��(��f (>���S
g�P2m��|���V��y�$��rV���I]/���3nl���k(A�8dQ�/��7�dS�eE�*P�����]����T����}�Zu�Z���P
Ǣ8�jñע��6YF[�2K�P�X�
��t�[իK�i����������b���ǒ ,�7�dqv̙ߡj�ȉ,ש�;E�����1���g��y��䇅$�b��Mvv�3��j�߼G���hP��c%S~��z����='�d��	H�S�t2�8�^�6������/w6���Is��dkl�=����ŤK&�p��Nґ�p$T���a��K��|����[�di���>��������Di�Cwh���jAcq4�U��YS���Ɣ�B�*C� V�0�U������<��1���b��ؒ�n6HJצ��`�yY(����|A��=j�P��
F�3w�r�ْ�P�lU�$U^F�g�j	7]1�K��נ��uGWWw&��GgD$��)Tu�*n=z�0���;]&cs��ֹ���n����i��e�Dە	�,e4N
@+V��H@0Z�%�q-��2>Ʉ�Ҧ�I��0f/F�A�>�4ݫl�Ou~4M�J�j�N��E1m��)ê��k�1�4��lu�ùU��I��Sv�F���6��Y�  EBE���7�KN������F����V�s21	Q�O_�>gu��mc�L��9��[21�N��u)،��K�o��� u�t ��+�Txhꆲ>���jZ�s�AG$�6�T�ڜ�h����9A+D�<�o����蹾
��^���Hc�fr�|�7�7s�T���_�2P�����ݾ���*��s?��P���^"#
dZ[ Rv��q�q��L���U�v�wY�-�W�,���4Ò��K`�,۝p���1���G=V��5(V3U�FG��]��"ҏ�S��)ǩM{G��T��v7�֡� ���
`��qS��I�PVp�`^��&��m�>�U�ٔ��/>�5K�X	�ߋl�|��U�b�du��U�m���=}��Ѵ�id+ӱJ��Un�@�WsgO�L��g�iZ�e��ԛ8W�V�&$>��S]�NV0D<��8W.��������,�e�t��W�����9;�%