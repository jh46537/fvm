��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъQ`/�P7L�$8�-�;�㻂�b�S���[T?���EL�:;���=?����re{%�ֲX�r���pft���1jۯM�=oٔ�ۃ�jP���c��gS%����zM�M� ]�0i΂�����n�q��!/�X�N�����2�����x5l��IB�?NId����Mx2��b��-Z�DM��lW?wu7��/uN������6�ũ�*;�L�@�.��c�W,� x��Ю)�sOL�+"'�T�+v�a�����19[�Ǳ3�6ĥ�Fҏ�4�����&���z�V\�;��QB,�<���Ve`*����K�MK�9�2�}������:C�0�z&\�ՙ!���߆Q �\Gۖ
����q����o�	L�#e�%����[���#�|����$��%�-|Z�JK_�S��<RK��$����G��|}zHV�h���g���mrϿ�c�?�UP;�����E߷
æ'��L{��l_���-U�^��YޅL�,�wHu����s�_���Uj:K��������-� �0���f ���_DB�&d�������8���R�7�݂&��q��5���UO�=)���"y�+;`��aY:����D�q�L�廣�*��jx~ge���L��T���CaN�[�[0}�d��j"�/�5k�KA�w2���_վ
.�
p
�`�oֿ�w�ⴵ/O"o�� �.fW��']��k�g�p������ukw�4�+<�jfV���-�@c2m�(K����v�h}^ ���+���J��Yx�u�H0b����f�V�����X�8�J�U��`��[C��N�3���� ���]�!��f 6{�����Y�bM�2���,����n�9�j�|h���d�gB	W�"�ܓ8�7�vQ� 5�v�M���n�X!}�?n����N��(��o�m�f��C��
�ׯn`�1��q-9fr���jʝ=URSYxTz�3���|��D'�g�Jd�sutf�-@VK�.B�,�\~!к�\�t6@�o�c�����9r[)��eg>E�8���
��	�P���xEְ�!�q�?�f�5���K�|['n���7ї���5B�K��}��D��j<�f�����B��dp�tn%�������� �kゖ�&��"}��d�nm�.A�����nM��M?�/��:g�]���<��i�kSPnP^��������I�ϰ��V����Ҍ�U�����`����r�ߩ�+�D3�C���;5�-�0,x�W���r� �Tg���"HT֨ԉ�ͣ�ںY�T*�19�(0Wѫiҳ)�ܪA�Ϸ�~]�!�71�
�I0j	Wr��`"J�Ki���=��v�z}���t�`�%����_�)��"�Yj�3���sr��m\�H ^�*��⿯�Jh�9�������E�}To�::H������B�V��v��VVPT3������׉.�,�Hn�!����Dm���V�<�;�u���pG�=2���
z�a|���*��P�s��y�0+�ڧ`�1�`!�l��1'�h5�����v����{�Fk�  ��$�Nd�iC���D�@^�Cz~w��'#�?,�3��e��,���+K�����8y���Xp��4�xw������t�u��֚N�"�� ����y*��n��-�H
�K�� �0�`���a��Dr��5s�2��0&-x�EP�2���I����OZ�*H����cU,��� ��D�P�+v���h&�n~77�"-c�8�/��2���/�Q��]x#`�%��]��V�dY򍞧D�,u~�AV6F�*DD�+.8d��� �mb˓~�����B��^".��B����[��ޓf��������{<hH��XCru� '�}�*W��aS�4��%����[�X��Qz����W�� �~u�~�s�SFyݼ��.��w �L��-�]C+Z�Y|��]��R���ݾli�����ҥ�	%���j�u��~��'��BoO�65	X�B�dG_	m�?dhR���D�5���/HZ:G�	g`�;51���.��|z�$�[��Y�o&���C��A��O�l� 4=|
�p���������N.[�z�dg���1*	e�럴!,��2����+�=�2�ٌz��h�	T���c�	m�!&�1#�HI���=��E�ԣ�U*x��� �-6�����֚�����'�E$M=�^����rJ��D9��+�v�5�Y���=��P# �파@2���L	le���s� �FOX7�ƪZA1��;B�ZE�w,�A�y1��ر!+������,I�X�'H��
 �.Y�x:�Tm8a�(���{�=�4d�zS	R-6�x�@
��]L�sEA��N�BpZ.�����t�=��g���l)�������y��t�w;���t;����Zvo�+�\�������Q�R,U��B�"Z�&{��b;��W�}� ഛ6V����\�����ϊ6uH[�������7�Б�IW����e���wC5�#�/0T��Ɉ����y��j�F	�}Y8.�z�=�b��oA��0�Z�^ʔ���:BkJ�h��cV!8�b`rհ tކC9�S���c�A�t��
zY��d�yx�nǷh��9�m?F ��"�;�T9��!�5����()6�dG0��T�3�u6��h���P;\�Y�Y�#q�rT]=�0��F�W{�qEڛx����׉u�y���i���j.���@M��j?�B�6�\���%�4�h��O���&C�8W+��tY��{@�=�5����D�Y�R�&2��!���e���+4���l����va�Q��DX��
e��s��a�-��7$$�W�dVP��f�u�n}I�yt9Fo��<�Bd&0#t�:K�~bb�+����nI�3L��(�)����+��i��P��A�~"K�*ZƧ"|��\� ��8���h���T��
�s��e�'�`e���S���`sJ�I1��9=a�SAE��a���1�d�qV��"�L2��5E;���v��/
g(�Z��;���B�[�,���-��I�þi�3!�C���s�u�Y�V��B7�����7`��	��pI&y7	\�花T$Ic�Ӏ9�������%R���F��o	:'n�&uI~��T�_u��O4&�>��¹f�RS�c�-r��|bIa���00/�V���ʢHš2Zp�b��7w��8֛g�[�"��tmR��V���Ԩ;��i�(j��d���YL��mQ�q��~�Z�dD�k���A���}�B��S�������!սV��z�p�ܞ�F	!�GP��Ӛ������z*�Nm�c��*}Ә��j`ͦ3����2r!�%|��_oS
���[S�~���o4��w+қG�
L�n��_���?m�;ҥH��f�F���� �^��^�j��A���[���Ч�k�%%�"*��m�ᚊ��0�d�EN��tu{"s�1�,�5h�?���c�{ӽ[� ��
d��2}C3��:19�V�"S�ڲ�@�plxWT��B8�w��]��B�~��1.,y,��䡢��� �HJE� ��]��q; "�1��T��oBE�Lf���**0�>7J�G`3ăP�!2����g�6n2�QJ�g��\c%�����>p2B�3W�*t3�2:�]�6��&V��nt��h��H���S1v�_��M�*@H�N&8��t�F7ϯw>\����Z%�9q)�4Wc�6�ԛP�l��~m&��k�\�&�T�Z7H� !X�_<�V��H{��,�_D��+o!�B���D��ZH �M�`=��L�g�v����۪�퇇wZ?�)�L~�<ɽ��a*��A��;�!�q6��|a�D#'J����j��~�el����,�O����B�$^c<��c1S?��zj��e���XדA�J������4^?��z��.�ڔv��%�Y�_�&ɖ@q#d�:6x[����QǨ2�0���M��_"RT[������M;�w��%�� l��kH����iV3�ڀdƄrYⳂϔ��/��nw���t�C4�q$��p#	_�h
G!�����R�Sii? C�/�KlG��o�.a6�?�`/�ȯ/�Prt���uA�`f��<����G��jRB��9��'�L�k��%�yT��[B�&�u��D��w ���&�H:<8�,A�E��i��bf�*��1��#u�|Q<����0��̇�s �{Z4i�F��;X��ozH�kuT��7n!ñ�Y�p���Va&?.�D���sp�H�ژn�[�����|��Oc�M!�	�A=�-G{C���ꊦ�9�`�s�QJ�?�X���|�ꨲhzc���ر�O0#��z���TE�e�C�e9�y���h��C/��� s����E^��vI�۷i��BTcP^�20��
T�C���X]���I���5����K�=�����ڙ$������~e���w��UHZyb�GQ�o�"���l�.Dro�J��+�S��o[��d2Ĩ��b�d�X$�����r��a�KEץ�/� [��!K�3<(�����Z/~P1���p��R�2�ҭ�h,�?Ii����f��ϋ#���d�0�MbeP�ŢRz�	{LZ�m�k��W�Ç�\���q��I������rR	��n�U�;%���� ����~�p��|�-T}��GޑP��x�2\wN�ȃy<�o��l�J7�r��B�#�h<���@���c@���P3$V��q�trT��g�H����g�ꔕ������!��
5r.ś3:��yV������x�s����&����p�#����q��fQ�X���}i���;��,��7�]��������� �;p;�8�q��ţLX{�o����?Z"���{��i���Q)q��!��HC%�3*�˸2�G7�E�fcS�/�rKƐv�V����Sp�Jy���s�W��m�������O�#^���-�LlX�����I�˅J�ϓh�0�lk��������6u��
�/��dE��"�
}��}7���!M����i���,�Ku���h�x�l�H�.kGl����H�)[�b܉�N�m�N�~o�&������4�O^N��rde�ʢ]R($XX�L�G���>��/4��O�?�ē����l�m4�-4�$����}?jm�eQ���0^���u�iF����1����ݡ�T����zp&��,s�j�5F���e���$��M�A�[|k8>�V njו�"C�È�Sj��\b�NS����Զ��>�덴�ڹϛԓ}`����L�FU��I�3gğ6�8��h 5Y�Gˀ���=�P`�u<�������XO�B�*w\'�MɍB���B'�o+��³����v��B6�XSU�e�4?W|-�My&�A�<�Q��J�Qn��f m��s\	5D���V#��9���Q'�!jd����NO$�Ţ���M�6��P��;�Fn��)2 	4R�W��E��n� 9M�e���~���pV�]9�A��K��e��5Y��.���@+���f��iX��Q�9�o�_�3�����j��h����ޥ��tq���B��v���>:}ڔ
�R�t~�ر��6�-N�*LB��9�Q?˪t7�:��W0���>�3��k�����O͛���e��^��3��It��L�=�胏��_H�hy��n��h�i���W|3��ɋ���Z�w/���m����tl����q������m|0k`	Lk� ���y�@���B�G,��N��n��k5�
��(q��� #Ry�[ǐ
b���+0t��̟@���A�JWH�w+�'���bm��.L��wv�R@�ݎ4�	��E����E�іi)���'v87�7D6�*)S�{�l�0:uRwƦ����[y@U�6�m��:~aeѼ��2N�{7A=�L��3a2��L�Cɀ��g^?����l�s�i�px��m��.��D�O�9�[ߪ�X=�:ysl��s��F���KRs��{�1H�8L
E�e1�%�Lr�Z��M^,�n=����7�>�E_��K/u���hs��;d�������8Y�-��>��H�Sa6X-\w��<r�k&��"O�G�p��n�������s2O�����a�R<��[�?"Ä�s�g��O��N��	:�>M�p��̒;�@��gA*:D�1�+\�H	<��؜�޷��	�%h���{m�|��x�0l>ۥk����:&$k��8��h�oZ5��ℯYII�1��"a^���z	fs����S���ޠD��h�d�;шY�� ���Ut����S���SD�e��j:M�X�^���`�7fbԞ�-�-��=nK�_�0I�hi��tv~֣��ծ�|:B0~��Gf4ĳ ��S�,+��O;������~kն��=��M�SWU��A:g�.�%N�|-��V�Q����H8�T��ζ�V������
�j E�šHRN�Wҵ s&mk���bu�<��mE'r�S�����c��U���	�T������������	;	���� �L^U���9������H=wPR���Q4@t�0d~�����"�a��K��9X�@�]��9�d����?���J ������=�F�0���%2�!��lʂq%j�y�'����
E!{]:~6]�y�����%�;-
-�x������؎cp�Rj�������{rB�Js.#��x*���H�G�߇����T�.��I��vC��V�PDu�-�80ͩd��]4���^���������L0�A��Xd��٬7t��7��B�Qv�,n,o�ޝ��.����K����1��.�X��g[I�:8-�:tz��`Y�S2zN{�"�^/������,p`5��f(Y�3���BmW`q�������,̈́>�7�=Đc�],��үm����y �������X�3��%^��٧�ϼ���aH;D��G=���obQ�?|�'M�SPP4�E� �2J�E�ę�:9]�Jk�����։G��$�#��l<�o��0A�,,)ޜ�?�����U#zr��C=��O~�^���g:s�M�,�
������
��B�E�9�Q6�S��#�^�Ε��</ѭ8���-O��{�e�*m֧e��H���č��9�� S��nN��ߕߣ�w���2S�2��H�Ь�����[.��2�~���4�f��/р�/Q9;��Ɠ.�dP�����$x��H_�
K�PV�#�7,�������⟎�TlP�n�yAW�J��v�d�� �՟u�u{I��k��a5�8=����0�w��� L�N���=��m�u]�9mF���ny�Ðk�H�"W��۱K��¡�,;rx]�"տw�(��2�A�n�2L����6�frq�M3n�J1�M��?�!Y�Z�& ۼi�E���^ �TP����3��Ub��"#���L!��~j]ū���hF�YwĚlB�砏�f6�k�;���i�DI��*�3���/TE�w7�{l�/b`Vp��҆^(���W/Г�S���r��{ںk�x|��r��Ø����z%!"6R�2 O��c�b��R�u��@�~�c�C`�զ��y��i�)W�1
���Y5�|��b�=��c���r�D���܅�Em�@;28�w��Z(�{n�W��m���>I��N�Y���
��a}��%_���}C�z�t��sv��¦�9�m��R��L�\�RKY#���i3)z �����.C��DTa���0���fx~�@b��lԝ��!�:�j�Rn��X[���zD�XWj��G�e��\)����Ȁa�Fa������.NX�i������$��=�@��J� d�޴���9��ۦ��ΎOYu��D���j�|e~�2�t�kHuϐ
���AT�  x�C%�>������^�.+9���B3F�<ˣ9� ����HP	�{TrP�Ȓ��)uvCm�y���G���A���㦦��2���i׽���i�+N��7�W����<����^p J�m���a�`p�A]"�O���7[(A�?񣗓�~��[�<rM�Rm��ѥ���D�?��D�T�H���1�0q�{����Ы�j[�cZ��0ۼ�/)����)j�Z}*����ޅ�hSsh#�=�Ј����{�����/]��_�42p�N���u����M�^�Z��¡�̕v",�>����5a4̐ڹ��v`���~Oyʈy
E��j�^�Φ�mK�
���U�\�=�-$���RTL��\':M
3MMh-dh�HS��1APs���U5oqa���a��io~��8��Y�y��FE�;�b��S�CO����|�<��X>4��G�*\��� �&������L��l2��;.�˖ d�I�v8/)�/�Ʉ�_�R�t��ZI�BcT��O��{Cٮa8�Z�z�ķƭ�e�b4�N��R���x" `V%9ohR�����M4;!P`$*F'�6���������35�x"(���U8*��Ъ��_!Ә�r���
�m������2�/�b���Y���S��%>�`��#Τ��'EhH`�1f��~%�R�6��c7v���R���whsT ��(a���푔���I�Z�x�Xl�]�{��] hºi$���8�ȹ�}(�Ӻ�[99�*�[��DI7t�ψ(,O.�' D����5�D���d�Duz�]H{��δj�qi�O��F�N4<h)'m�k�V6Z˃7������¿�`��N�8��T���D��� �+�qX�$|W��tdaIĸ!���-�E_�k/9}��ry��5��9׼�ad��o�ޘ�An�L[�������H��8�D!W
��7��D��
s�z�ꘑK�Y�/��
�	^=���(V���my�?���lA]����FH VG|�S�\�_�A�q�T�X�6�]���K!ƮM��)+��t�U/�ґ�)@��]����h�s�c���t�'XU�=,в�vdț���hʹ�˧���韈�N�F)��#��Z�
N��bL�h�B*��d��\Q�*ǭ��lo�}�����r��F�
p`�;�\��΢^��uS[�G|�UG��Xo�7֝9���`�Wl��q����ħ�P�O��CTf\�� �~�T�ht�<x�[]O:���F-��Qu���3K3{≡ɉ�[$Gg3e�[��5�6����-�]lQ�U숱�[��c�,9�N)�2��I���QkDǿ`sd�i�m0�_O Z��~�V��6$�'��F��&p���HYU-�o�W�����E�	&��)���v{�qd��Q����h4q^�ݰ��L��L�4ﳖ�]c[�q�T]�l̾Ca�wQ�������vu�v��=N�wa���P��������#kE�!Vx?E|���I�L����ƀ�fJ%�����*��H8��Iu
�z�7�r�Z��4
J5��0&Yt�Rr8��i|���SK����_��;��R�*�#���p��3����E���A���X7q��Xx�Зd�>m����{�xCa6%w�A��~{h߭ZǞ�H���߈��۴":J�ߐɭI8(w1��A0��}̘�:C�hU����:y�4�������t6.�)���F����x�u�1�V�fX�F�έ[=n.��md�@vĩ��{W��j	nxHE�A͝YD�⨓=r{�G���=���0��M";�� 	�8.X�J�W� ��vb¤�'���8U�+�9u��Hqև<�E'���R�A���'/�g+QE���. ���H�8%��?�e`C'�⎀�n%�e.6��pm��+0X��e�3�g7����ƨsW�޳P~����:F��^�̚����]G�*2��;G�EVFJ�2~��ȯ�/�g)�;"���A4��\S��o��`̷˗�o�����R`˄���� -=�j)��$!O2VE�����5��ѐ�/zfj���@���C)��������m%h��n�d]��D�f�n�ݤ�c��$��`��Z}'@��d��"g�,���Y���T�d�7�Y�"�[�[
Iic��|�CuNr��.̲�w���1nv���0V��|�4����!�F�S���T;�q ��!�J��^%�n���t�B��NqlLF0�PwkH����KF<�]o$�����]C$�݃�xJ9�zJG�SI�F���Yr�g��?DD�
�t�xSA�SX���帹{v���a^��VM֕J�e 'wY�*�:&�سp��ү+�9��2�2�k9IP,� ^�`QG�"�?�h�p�|S�a���0 Ҽdn�&�p��%;�Uͯ���R���G�JU��R�&p\����M2�hmci`����P.i��%Vʐ��ܤ���� 	��I�;F�qEA��۽We���aD�� ����Fk��dF��m��.���h�(����+�yp=<��'%����X�?z��w>����~���s�����"�z�˖;�D�����7/R��(ʾ�S�r��T�ؠ*:Ӂ�z} ��9
���;W.kzL�9:��ЃمQ��o��g$D��ݩ��,�1[�2����īR�d�u�y��'"�+�J�Y/
���nO��8�@�"�J��gu�T�a�0��h64�H	�0y�*�����tfG��7��9{l��p	�6h�`ڊ�4 
��ȸ?��i�m��f�R%��zd�p��	|'�L��q������pm���Hj;��:���~N�o�s��V���m	Fl��H���qz<D��q�g��|��:ܣ�Qb䉖:��/q��_���A��� �l���L��KiDFv+͜�Ǔ�v*���.ԃ��j�7G����d�\D��혠�U����N`ǈ�3T���LP�jP`3�J��E4�e̻���>~����E���OS&-a�-�hz�Kթt���#OM�65D�Øw|��B�Q��44~�xȜ����ax�L,+�V�3�6�K��M��j�!�����1g=VJ֠��	T~�_u}`Q�>kW���5B^㣗�"Tc�#(�޼����6����,��Vc���9 m�o@�#�K�]�m�5�fҵ�GG9�o���V�073%{�q�﹠53�7� 7@j�?�n�S�Tw �7�*�G�X�L0&j/�5���!8P�}�s���@;�uQ¾KlQi�����6��,ܒ}����x1s(rіqLEL��G�[K��G�(ڨ�1?���ZT0)���4����/|g�`�!������l��g��{ݧ�DS�ʚ�d.��[���>x�q�z�NWý�q�ﱭ�C[�Ӵt�������|ٍ� �1���H�UP0�'>�S�o��ߓz��`��V��=oRH���Hy+�K`�浰*��(���;�kR���KR�l�� Hi��x	a���<Xa���?�s��F=\� �l,�gp�jNQ��ѥ��'Ns�V'��W�����T��[�D'@���m)w�P��n�8�@�V��ɜ6CVj��3j[Q��p�4���u0�<���2[M�KK*�ۃ�j�?�<��%�ٲ����[A$��.g��͢K{��-'�*���>^���Y'��k�F���SS��4C"��Nw�*��E^2���WBk��-��:�:�8��:��g#�!'(�2vI�V6}hʨ.��m1y��lMm�?D��&@ⓛ3k�8#�X��Qs>�s�hԞ/0C�fE���ũ�Kt���}|)O3iZ����b<��!G�Nq��~`�����T�`�N����F-	 �:¨]�0��%�:���W�̕$�����\ؑ,���O c�{�mn�6˾�v��W��ܗ���oXV��O��?3����x:�����(IA>���;���`�M�ϵ�4�M~ԗ*9M���V9�؎�O3�O�6�@�ʀ%�Cy�%��c>\���_���}9C����D�ԝu�K�80uI��S���-�!����$���}�K�k͹[�5B�o/[󴿏.��NcEv�rH�Pƪ�n� �0/��"H���P�Õ���R�4���̆� Va���άoE;ಥhN��́��J��4U��JlN`,��ԩg�t����N1�����_���+c2�}� X�m#9XM��J�i�V�׻^�*��̔M�M�؋���*D��z$A ��Wn�̨9.K��vv|��<oO���3���O�+ԿVO'},�t����xV�������ԹK�UKUi�K���2�W���R9p�ujR܌�����
A�wY^�h�r���w!T�H��)E�4�|�E��	�mC��.@u�C�>T@��ʻ:�n;/2Q�Z�`r�`wxG�
�	B�W�q]�#��Yţ�`�6^����yv�F�f�'��Ʋ�]�%F8�w�3ά�Tj�%���~[x��1���O�o�-���ёs����F`o?	L����qFY�̦��i&'�s�Բ����/���ǛR�Cg�)��:� ��Ċ�k�RW����y�u����Y��A(��v�õt�A�Zs����◯Ι�o��
�g��&��Ŗ7u���Hpľ������F\Ij�7z�h=崕�Ӧg��Wyu��w�+c k�g����>�uA��J���(:Qɔ�"����/\~;]H.H�͍ɋ4h����J	��jz�n ھs�Z��#��z?������9hDZd��/����H�.��z��ڦMw�������֌mP,���R��֨e��=����ӜѾ~��@�gF��#E42<�ֲH+(b�^�5\	H�$��&�YW���9��;��b4���K�D�a^?;��c�c�Y�,Y3�������1��b{o����uO���>0-�l=�ua9!�B?�Z"fR�f�Lڽ���G��"� ?����w҃��T҉�z%{R��GY!2�~v�2Քe��G[@��
�v��#E�n�z��|\�N~b	ә��+,R
��ݱ��K�ܟo�Mq�DO�NB1�5	y� ��
��cD�y�O�k�|�|��_,G�Oh�+K��QI�}t�
����<���A�0/��!�����������'�^m�=t�a@P:����^�_tLZ�Z����w�\�IKWh^_H3��bM��ǈ�6��������e;Z��*���سE��Q���\��};��'|M�=T�b�r�񫞆'%a3�Uգ�_� �Y����w�Q���� 5��P�ZC��4r����4ݳ⾗�K����	|�PQ��GnE�vGj��p���^=���[�t�C=��}y��#,[K^�$��`�禊��.W�$Y�zGӧ�}]�Pl�{��vK��c�
��~�v�PN� Ѿ�1����	h�fD9�� Lxi$��j�կ^?���Li�K��-_qr��O� ª��Е�S\�棿��/t�E�)|J�	�z-���ª7���d>�/��I� �2����o��x��a��N	�2{<����ʪU�u���`�,��=���Վ�h{���<���!tZؓ ��ö�I}ˉ�G5*Pa�Ќ�j��N7�Ac39��"~����خ�� d��� k����SI�2ca��K�@�[�k�L�6���9Jh�!ʯQ�������p��T����� z�hC�T���yb����b�7�Fd;����,c�nQ9x�\0	\0�%pIuذ���&��opi�I�&��,3�󖱑��;, i�/%����,{�kh�t��_��F7 �x��ʔ ����I^Fq��f=3��*��w
���t�t+ە��x��@���i�Hp�V̓|�i���n�7��9�A�����k��n�0����GoFl|�D���r;�ӳ��z�GO���� ��(���ʗ�v��p<���{��.���(�W��誋��0*��8�9�$gĭ�b���nT�������`Y<������3ѐ䁯���Kyr��0���a�� k+���B� �%| 77ZT�/�%�0��5?�v���������L2�%Ǭ��o��}J��Ĕ�|�D/�c�h��G�~yN݌ ��Ȳ���q�ݍz%E����e�ő��Qn�'�a��r��u�� �4,��@�\�!�}X�r�+/"4?�����$��x'��񊪮`�����`NB�5��tYk!�`]fM��[_f��1���g�ȥq�e�fgOI�)�7��v�7���kn���R+Ah��[��4��HmR��u��6�C�m�gYA^�_��$lL�5����wG�bm?~\���V���"�&����̯t��Ƥ_D�٬��|�