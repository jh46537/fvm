��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S�VJ���ɾ GK�rA�!��}�x�E}ݨk�fի�u�(���L K߲w�.L}x1F2�#5H�:�'))�6_��\j�S��W��w�.㆔�[NQ�6��iM�@��9��eh��L�@�Fb�%FZ�"e��R���W��@�s3a�����膂Y�:�D���!G��j	�E����}��Ui����kh稯ka�"������e�^��6�ɠ�Ij��-���jW}e�@,��=��\�`�Ǩ��:>_2�)����������t*�� *��%/��X_0�2�KwS9�ڪaԟ�	�踷Q����Z�@Z|�歊�)���ܰ�K���"F�"�;�ŰS�d&>�،4j�o�9���xD��h[JH)���m�tS����\�ɑ� �n�{ƒ;PM�����>"s��R��m(ɠԉؔ�W��6���ߜ=�5�%�_��+*�o/�Wv/�nW�S������50�u#�����=�O�3b�w��Z,L+F=5�'�?y{��yN�2���D2�m� �p)*�CW��F�7�Ye�ȼW�xs	p���-0Gnނ���Q��	��q՜o
����D+�g��!!|VeG*�s�1� y��!��FXV/ao�
Z�#o �xE5�_�=��جƒ�K����#������\?xi`i(d����#���&S����$��a%�o5�H��}\�����?�ՒI�W��+|Vz/:�2�T�K���f?�k��A9���d�̺}���6���K�����T�ʫ�n?�塲������*}�Y�9�{��S���c�{ҩ����H���qn����qh��W�"�&sL'4Z����B��,8��w��BFd�8M�Y�b�oe�Wl� }�$�ՇD�O����r,���1�υ�\\v��<Ɗ��h�L]@�'�Z{�e5��w~��t�qJsP�X�q)��"ˀ�-׍����������@�(� ��bx������O�3�Ӓ[O[	�Q�����c���x������_��˸)��+��hNۚ�-�4�G�[��T ����r�͸���6�GY����G��E<Cn'C@>^=0�DFj_�hEň�
����6Yv��ݚ�n��r�'U�d/"�OS����<�N[�-��������O�oH�Xd�K�qF����mʞ淛�vKBDݽ��F*m��W0��iH*�SM�-s��a�fո�5/?�ز�yw����Ʊ�^3�T�%��ޮ�~�N'kK�u��M;�&8&������0a��B��{B�t����@ֺ?n~`š݀۱�
���
��ާ���2o��E1��*?�X ��1֐��g�0� Z�(ӖrA6��r|�5���"M��� �zrU�Y����A��-���Ӂ�Q����Z/*rl8g���1tFC�c���$	�����K�?������5w�"����xG��i�&�k}�k�*|}Ӣ�#K̉|u�_&�o@&.�
�\��w���ߌ��L�S[ {��3J��2���F�م��%���}~t�:���]�;�q.~��j�+i��L�_|D�s���Qa�!�_l����=->݅�����()�L��̾��94�ċ�2C4�N%�*J��&�+N�,'/0�^,a��]S����;�A�H�Ȍ�6ua�=����F��%T\�4���K�I�2Ӡ��R�D�-nt^4�P��y���ڹ,]�j� <;�f�I���\JY�Y�����Hu���RK�C��p�2k�a�M�Ǭ�uR c�H��(1����" >��[:�
�⬿�(���r<3Ku��K���{�/�6���w �z��݆�����-�u� R��o1O�[~�����?�b��)�9��L�	l�vh�/��?�g]be�*N���)N�W�ZK��x�)`�*R����6@ID`����vFګ7��*�^�ck��/�عx��Q�
>�]I}�b�&D%YD�E=�-������m�c"+�d�'i�,R[��a�p�O�2	6��c���~CÈd�BRAڬk���t]VKĕ[�ρ~o��������1��>�t����c��x�X,�F �h��������ő�s�֓ 
N/�m�y�VC�����B�������e��ѱ�nBx�P˿����H)�������p��W�Ϳw��"���4�Z���?��m���
Z�a�&5�=���Ԩw9�����j�����5mM�׻-�z��EN�C{>�@/�Gd�:%xə:�9,���̀C6t� K�Iγ�.�����d�LX]9B8T�R�����l�^��V�ӆ�i��4��g�s?AtH;?�Lw-U�yg���ủ��k�0� �"����<���o�dƗ�pBg��#��r�a(��ho���V,�b3�u@2dk��'<�t���GcV0�]��,��-�=�Pػ?��j%�V����r+�gYڅy~<
\�ڷ���m
�\����iwg.� +�	��N��6z�MU19�&�<���9���B.��g?��[��?T��F��c1iR:��,�Ψ8١[�Vy(� �_��d� ����c����bц�pv1j�B��v�q:�w�<_�v $��Q&�
L�C�v��R&���6u�?T��K��0xp�@�Ǿ_ުJ���slS�1Z���ִ��3d��䣌�I�Oل���-�\�����7S��kZg8>�hஊ�;�N�����Dz���-�h}�h�������@Lo�Ӄ���QC�-�2˴��Y6��|~�߂n�;�
�Jǝُ����Z	�����-C��F�b�G��G�,fU�!��,C�6-mj��d��IjۚX�m���H�ҳW�͎�dQF��#�k�m�>⽎�>8�.�m˺K���E��V�����p��N��s�I�]g�
	f�i��`�*����-�A���]Z����
#y� _����q�İ��mR#��x�����z�qLl�S�Z��T[���&_[u���Yg	��k,G[�  �L/���=��pf�nPi���޸�-�u.xw�fPlmh2ݖ1F�Y	��'���.|\`Q�Cz��g��	�DP��H�ĴcOo�=��!TP�l>�$!�[-�s�@��b%f��I�PP��Y�	�j��XƖ],�>w�zO��B�����ye�`&�S�o�vxR7_�:"��&l{�%��xY��Ʌ2,��q�u$�-��(�z�hR�I��m$��Ӗ1��xu-�f���ݘ)-�+�� �
:������l`���	[�����{G "�<YG)���y^c}Bp:�%���j��/	[ؒ���W1�\l�!+e~P������v?�i/�n�ܶ���F���o��L�޵ʢ�p(�F�7��r8�F�Y������C%_ʼ�Cu4 ]�P_�.�p�v�W�p�	�<Fmm�+�+�V;1��YiRV1���Snz1�ἃ,�
���H,�]��7�l�+@��#	����I0�Wk�$��+��㽆����n�&1O0�6�t$o�늙3��ނGx,K��m�0$����C�
ifݖ�	ԭ�^J���ݦ�W �PZ�������đD����r_A����^f��8��;7 �\�l%D�_/��y�&7&^E�˗�N��H�?Vә�q�!{o���(�C��F��^`�H��	l��\�� fv�-�������>q�[o�2>�)3X��"[ȳYp�)3&��E%!G�ܞ4j,vK���0h3:�Z�/\�pī|z)#2G�_�c4�H����C*�>��3\���FЂs}�{0�#�	I=��"]7�y}"[����: �X��*�fWQj�P��bx�`����	%�z*���n�O�P�|���b�J����=Q��b+���; �b6���`�����S��/.-~Z�|۬�Թ���������b��s��.F��n���㿎Æ^� �əO&٬�� ���u�O�.�mI��7�m+�ڰ=�Ж ���7��s�Izqz7KJ\����h�y{�߬�8��0ʼ������/� ��ё��o�]U�\)9��K�WpJ�5�n8�����+�������O�f4h5]Ыgz!d<�X����W�%�W���I���OJ�>_�ގǜ=�NI;�#N�/�د�x*J�*����/��&�N�7��N�?)H4�I-ZFD��[1H�f�q>��F��#Ц�r��{�g���O���+|�;����;���pJk����Y������c;A���?$���A�P��t�g���d�Գgz.�������Kc�d�ɴ�����[�^f�4�/i��t����m���Є�М@�0�)��,���_:¥����xR�ٕ��n�%l?x壃���$&N6*�Hs��X��꣮�wJ-#n7�yf�d�Pŉ���r�G��0oaV
�(Ӝ��͒	C���}#�E�������4��0�O��ߟY:Û����t���,��}�g��H_P`#�Ǒ����|����>�F2�6�ʂ��-q�_C�I&�T�æmD�L�p(_����XP��%N}$˵%�
�6N�!�]��h�K�҅(Is�u��8)�ݛ�}�}S��[�G�M�՝q|Ql�m�U�ro3�|]��� �u+T��,�b�3�_6uqj�E��!�抷�c?���(���d�B��y�-`gp9�k޵;�9K�
�;<b�*e��łc8�F]kȦl%��Z��}����;U�U�)����~Q�)g����~��\������-Z��5����I:QG3t�)�j#���1���亐�8؝�����r�H�5�R{	��ɇk���fx$S�m�%2� �ry���md|N�!t�]h*uyБj �<��%�� q�Hzm�	����8�� ���akM��@�㺋��)�<���]�Ijm�ԙ\R*���`��U�
���<�2�6��ޖ�产�:�_5Yk�J�NS:�/��T)�J�*�!*���z����3|a��/үQb�e!(@�⩫�h��!��	�$f��4�~m��N�o�<��k+W/jL�)���d �\2|��#���r�I��z���[��Wq�>0�69ˣ�!w�H{Z]Kv�ޑ�2ԬZw����mQ�����%���A�V�0���z�Wm/��!��}[46��\���d����O鯌�I���k�dg��5Km
=��JO�ި��=�j�(G��M��g�{
}�!��Lտ�Y]���e@��_��;�:�Y�O��Yۇr����¥j~~�$g�m)�� CB�XYdǤ�/�gK�V�g����?Ziȥ�<����u��á�|� �JBq���J�6_�
P}�r�Ѕt��W	�r�	�З��s��I�u�׋0�u:���9*� �K�׼{AnW(B9�f�+M���-��Ǘ#�,
|�r�y5���[j��@J���t�T�X}*F8F
��K� ����shʚ�W��礼��lX�0����p�v�ypN4��#��6C�t>=g"3ґ]�,��S�Q*�F�ɐ�ϐ�\�J�\�)�}���o��!��f6�x���J`bY�ଉ�k��v"W)�?����J�X�C鷐;�r���gM+q����6b���?��ԋ���|�7�cMD�.\�R4�o��At�ԕC�l#���A�K]��O()}8q䊯v���%խrl��B�(ƽ�`���.C�}?��:XB�6��"[�zo)��U��6^��k�z��V��$I�*+ �(>ȃ|�t������#	�"�z�,`3P�3l�>Y�Ԡ�䂻�et��G�τ��b�x�-h~�$q�h`H��(���_�E��<H����wV��ˤ*+7�r3�3�)?J!Lmt稚\��J��k;?�bg�}xg�a�үU\�'���v=��Q��*G9]$�0�Wb����6#C C`l)<�$�8#;6D�)^x�#�kS�Θvp�i6S���j�$�O� �u}!�E X&a���$li��R�rk�1F�MڄW�,>�a=�'f�����e��N7��z�l+�M����N�D�K�[X
�	�S����������?���7~�w�p�8��\ҽ��㦴�8�'E��3�}:����@I��0o8�2��*�>�b��S(C�s�+��ǝVpCSm��~ؕ�z����ŭطN&!ŷ�cŷ�@`9^\"��h�������`�
��!=3���_�2S7H�#����  +�)D����0\vRa#�G{Bm~��
�f2T�u�[,\��Q��Cc�W��s��1�.˞��V����:�	�٩�W�~���e�-�Tk�k�,zxlҩw������ʿ_�����vL`�/Q��k�5�<\�#��`�&��@i�H+�A�b�L�
�V#R����I�ڑZ�vO�W榾W<�wW;V����B&֛���x��c�93f7�tL�z3�d,c�h3�z,�ن����9��F6���+~��},�P	�i��yq>����i��~�;f�%Q��@��CXF;���J�8���y�@�ϑߣbld�I��\���..o{�_2ˏ]���D�ʲ��wӓB-�+�P�{C���f����~��~�]ǿ�J��Y��l�&�	F|�eB,]IXX��% 2�a{o:�̭��4���}x��Ж��NA��{D�-x%�l��F@�ţ.��̪��E��c`���P��%)$���AR&��Vs��.��yaA5˧k���>Γ�g���7<��ٜ%�/��*,j�	!��z�=Rhf�tԣ�V�zU-e�����lI�Լ��_E � �����yP^���w��օ�טfg�ᔽ�Wc��S�\�"ZC��Pm ��t���'���=�C�H) '�:>:Q��6[��b��^7:�i�.	�t;��#<<�ۅ�i.]��;l�U�lz��~|H=x/�N�kLΤ��x�\���C�՘0�Z�����h�eag����濡^H�L`,��a�]��t)�V S	Zg�-��rc[�b~�����'�2c���`F�|"�q�p�T�$�L��d�pY�J�I����ل#�&��l��U��]��� Gk�%�ǳ-�gl#0�� ����!$�ǂ�D����-aY��i��[Bf�Gߚ =�NQ�+��}P��������ϋ�F���xɼ��-&�$; Tz�Cu�Y�k˞|$?!�C쎍�v��(OyB8���=;��d�
"����i