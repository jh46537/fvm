��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]���Yq�<���Md�3fF�qZ�Iᭈ�q4�\<*��e�ۏR��ܟ��~	V&:��?~��Av>�R�܏��z$]�O�y$��N]rI'�Sͧ�T��}#�o\\�{�gt��;�_4#ϔ�n0���ѧo�[6��Nܟ,��Oۺd����wR��m 7��/����Q�WT�Ns���)�֍�%=�2T�;z�+F98(c�K��o����*�Js��U�Tp�d,��%5U��q_R�ӌ�s��Bv>��iwG���}����}�l�2�$������E�5a���Ј]��_�TM��Ve�=ǫ�f\=-����]�8�*0�r�$D�y
CQ}E����r�ۼ���Ć}^���}�a�oRߓҳ��hp�����!�Y��cD^��⪈��l�;��%8��FQαy���\L���"� �4�Q�G	��#��&�l#�_ڿ�a��n����atU��|P��I���\�r�Y�	y�0�>�F��Iߨ
gWJ>������{�pH�Y�h}�X��n[����%5qf$��F$�OMX��޼W��ؑ��+őg�7�vgڭ�y�b�Az�>a��㮾�p`��� V�A^���|��C�**  2�|�TS�R�5&?�����~?�p;n�)!_��l;@�����@0v�n��e��Q�D/Ц5��&S�:N_����2<��V��H����	X������i�����zD{��]�h��(�S������RO�g��:�| ?\a��[�p���c�\���H�*^O(e��R�Q���;�F�O�J��p�B�UVG�K(��t��ִL�!,=F^e�����^m����|{�7�^�#��ћE�'46�T>ôW���6d�;{oC�Ҧg���|����q��m
�en���t
'2N�Sr�V;be�ږ{�jH���o�X��Q�nM`�	Շ�0��64����7����sjSI�P�X������9���ξ�È�C	[��|�� ��Nˈ�I�|k���ڥ#����2C�u��nZ��z����'�ҋ��侺P̮�'ڮd���7f�V���P
�x���Uc��L�cW�v��fv(M���G̰����2�����f��%Y�s*i8�Oi$��ą��J� �6����L�^�h��b�i���O���p.����|�����\���9O��/-'r���	���/B��ԓc�A*�@����7T��˓Rʁ�z��l��(&0U����Ks�r�¢�� ���J&]��y y9���(�s��w/FDd2��6���7YɈ �j�S���;��)�G�/�?HbE6c�	*ya�y'�{)0s��+����3��,���2}�9?l!����B�pfM���s��*tP�`DdOǏ砇�,/�;�X�Ni�����&��溃� �:X��^xM�Ũuꮖi_	2Z���m�1 5wc�{���ح�k�W6!,*s�z#��=� @3�e��ّZR#��K6'��d��o���D&�3n'^���u���m�^$��^�>0u�~���h�c�4!�y"fd�!�@�a�ڷyG�"�WG#�*�-�y���Η���V7~���s�1�Y�_S��fҤ!�����'b�$��E���/�k�:���Y*�d����9(��g�&�o�FH-�P�Y@k�7�I�.�B{}׀�ng�C!;�u�qr�RO���g�gn膛�������q>�c��j-����K��7�Kj��J��o��T�
��f8ڨM�����j�O�<tr���\��Y� 7�P�#>�f	+ƹG�ё�����g��(��?#C8~,\��b#�����;�o�y�q7��ݧ3������͞r:QM�� >�#X�K�+��:��D 6��>�8+!(���=�qN��P+Q5{!6X��F�V�2�0�IP۱�m�N�F�W!\�����m=�Jx��X���@L�*�&7���P8�c�āo�f�u�)�o�����e��ޕ�~O!<ܶ�x]2�͌�q���i�C�rc!���įL��Y$0�i���"z�cƇj7�Ny��u�6�*��ᦒ�̅A�m�c�%������T'|z�{��wz���=c�Z<6�M'���G�!�:��Q��?�6*�7`�	�l�c�D���`)��������P:�~�����%�кsw��3��q�xL�g��k�"�,��W�����������!��`��V��;���C^XTj���V*�[T�/� v��m��9K��_o�����x�}�U\���29�ID	�L��?@h'�a��ҩq!��0	\X��<h43��S��z�1�pL��G���+`���g��urv�<�2r�D�<�fo#�Zd[��I��䑪��sDU��2�,d86�a�&q`l(��}F��ttB��}�z9>C_����h_��翱;2!�H2�դ�mwǔ7Gp�}���'En�\�c���cV�b��h���^#Um�d%ؒrs��Q�
G
U�ڂ�
䨪�����_�L�SI�K����Z����bRI}7�i��� p2�صe���:����C�����0����뷨��W⓽ϓj
�E�u%x�H���B��������$33���q ��������S�Z�,��>�����sc'Ťw)J����ҊB�z��0����6H�.́0a�Fn�UD�;�������	�X@�4��n�
�	�I\#쇤L��S}1А9�"�p<��2Ae�g�(K�}rl�q�?q	M�@��_S��g.b��ӡ
>o/ި�g�ɐhL�L���l6�h���Q�G�8��عWޜ�������/tT�9y)� ˡ��=f`d�w^�܇�n�|1aw�(�1�q�j�!���r�I��ykY}�F�H��`yK�y7�A�,t�45�f�s�V��2�A �A���3��C(e��q��=��f]���5���Q ����U�#�#Ĉ������CY+�W	�}���H9��Ԉ�2�M$*3��8�OٴӒ���o��5,����6��JN�r]�� v`s�b�
��.�LA5��:!u�DJHf�q���ΰ���^�sWt`{Θ�/�l4���~�8�+S%���'�J�Q]Rq�9���Wv�R���@{�Elm��뵶,��������S���C�\��/ɨ]QԄ��v�TMY[S�$�z^�ʐ��(�v�a�Rfj���cƦ�r k�o+�B0��1{/���uUo5(E��et��S콸������}
$���<(Jj6�Nm����*�Y
R!�2p])�������;y��s�aE��u)��̩��8���9C'�\�l�˗�q��C�����c㡊���/%�"9ЙK{_?��^�k�-*9�ia��f�G�%�l\'ݣw#�r�l�=+	JC��fץ���l1:�<Wb,u)�- �x�}�9��pt����W8F��>TxY4�:P������yҗ�Tk��.��4�{e��c�2Yl�&��0��+X��)"�n!C0�kn~c%�Ӟ'!��u`S�8;Vc\�z�[��X�t����1��:�Gm��G��o��JJ�
�����R��y�@ю�qزl�Tꞗ��"��䱍:\�7��=�� #R�Q6�H�o����Fd���Z �؁,W!n�A�fw��D�H]�V��I�~E�m�<�_9}D=��
��U�q�~��sYl���
T�$AJ%�K[}��(���O�8��	*Y=t�<Yk�!�	to�)j��a�Q�&�VE��m��[1�)l �I��Xy����B��ih�U��Jj�]���N''YLOj�_�G����r��_k`�L�(���?��ـ	�7�l%ֈ��|�2�k&���k8�?�&Ғ��	���DCSB*�2��_A����Uͩ��!"�>@�4�x?��V�Gh����^m%*�Td�����X@|��66_oY�R6Eƫ&3�Q'C8,�:����V���9��A�Tu�..1�2�M�x��^��db[�4�/\Fq�/�I�#���[� z��	���`����w�r��{&�LU��C��^4N��vy����@�5&t
1��]�U���U�<qhZ�9q42����p�#L�����r!�8��pW��hM������tsT���҄8�MK����@8:E;�\Ѥ��������]FoiT/r��Ȧ����`�t�y�����k&��>��4I4���2$p�i�F��X��ٱ25�IB6����e�i�%M��d&������K��%8��d:2�۝-ۈ�(��,�
�g-8�R/��~�(_����}����azh� �Q1<�����5Ay|