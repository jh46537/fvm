��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�^��h�����mb��feE���UM�l���`�1Wv(����&���=t�ֿF���l�p��� q@geL��x����)�oZLB���Ke��C]�X,f@�]iJ:x`��;P�I%��bSfi�|lha�{�-����L�𶣗�rҽ��vWǂ����D몉����"P�C���Bk.So���@��5Y�z�aۑ�ֿ��̣�_`<�^�䃪��q��΃rpS�r�sӛ���s�黯�f��ћ��P�̠ƺJp5.	v���c.�p<��O�V<z�Gz�w=�׀k�2<�}A�� s�`Ol���ZDyx�w<{e�]^�������{u,�t�:Yd����yt�t|�� �Ww�����s����e���y��-��W���c3��}�
y^�#'ੵ~�BrQ��
�D�V�K���w�u3�zn�,v�hɕ��	��(?V_���{�	6�0�(�8}%�J���v*���G�b�<�|zbHxM��	�I�o=���O�*�g>Բ�c�-O���I�F��#��;��}�C6.�����\Q�!�#aU�;/�bE�a��E)��-����聆P�`+DC�v%GΟ����Oʺ�kCX��
�-{����`3[!՝
'�3�2M��ʪ3��j$��.��D���68��BJ���Hr"P�s�������9��	�C	�������!$�� �������M��������@���&�gЙ�N��Q&	5�Ig��ű��4��}�sZ|�D�w�00�xR~�~>^��C�� �B\����}Y_5OOy6(�x.��Vi�D�+0�+�O�SF���4�&�m��\����Ԛ\��ݻ�A����v��4����=xZ�x�B��uF�f�WoG���pǳ���ga�^��s�5���ݬr0��jӅ�TGc]�m���\..��	��}�aUV����������TRY"��4�u���ӹ����:��F1�k�)R-s�s<-F�Wp���]�x�(��"��a����[���Q��{�Am[+>s�?:�����`��'mC�]߷���XkN��YOe�A)|ڔ嬶X��b1nnT�H�Z{�r����%43�L�=גxW�Ѡ\u�.�$�岨i��3��J0��]=)i����Z����7fv�dSF�D_�s� ^W7��f�0�a.��.n��� ����$��_J��d)���*ڕ����_�.�55d��'ޠ�� ��yɝ+q/�]�k���#>� `�M�A
H�$?5�+`�Wj�r�a��0x�u��+��d^�!pVX ����C��,��%�wg�w���!���zW	���t|:��x��I9�)ro��>�S�!5D��4�N��7�Q�\,r��!��S\]Iga5Y~:�!��~� QpQPzC�;���?r���8Ap;��r��7�]W��Ȗ~�ݒE��ҏ"�*\�T(~��v~N̹/���h�qO�B%
�-��*��XmB+�Ik@��RsM:f��NHj�M�?ǿt�19�ܪC�U��f7��l�+jU�����emf1�ۃtF9��o@�����/dmI�/��'�� Q��i�C�F�����k$�,}!��q�;G�`q�OLI�Ú��;C���{��G{<(�%숖:�j؆�Κ��|�tSqv��?{?;�l\ F���Y�Ń=+����T�D�q���D�h=�ʵ�i�7^,^�9��xf��v�C>P	�a�Gρ<Q����T����(W�11
e���B��i�S��ﲹ��=�ݜ�*n��\A翛Aft���.x��wa����Y�M7Y�NIV`Hڦ���6�<D��Q�P�sA�^Z����翈���ǽ�U����ۆ�/dQ���:B^�	��8䚯�꽈���o�4� �,[&�5���cUD�����SWT�8KlZ�t��z���(���p���Ms�Wվ�¢�@Z3�tH4OW�K�q"쮏�J�|�Dfh1D��H��$rC3�`ǆ��|k{u���7" �ʖW�ߔ*���!�O,�D���+5�)y^�_����P{���$�g��B���&��JƾGUbY1���&�C��W�m�uL�
�D�5��HoA��:��1+�KS��(����}�'��H.�@>Q���Z���Sh�!+!M��8�6���1wY����O&{r6��:���rˢ�m��bt�:T\p�~����$H)��]$.w�K�r�v���x;��5�^[�8-M��@�]r%��"�zcB�WK�K�q�d�r!63���k�����lZ�RY�?b� 'd��S��r��F�#e�¿�����v�m1����ٟo�B�.ThI-�^��|��̲ )��W����h�"�����T�"�z��Bɬ�(��5��x�ɫ�`J�)2����D개�D;BC\[j�^B��"/[�͡�R9n�)�ӵ����wĸ\MK�6�ȖPl�� �o�q��{kЅ�l<OM=9�Y�j�a�	B������S�7D���{�c�-�������Wi܆�#�=drN���+v, �G�q����q(�ĶD��Oe��{O�깹?�ˊR�sA��)u����7�9�n�F����#�:�k���ۋ\���Z���ME� ��b�d����}�~e�t��h�@m�?����Z��U!�ͨK�T#S�m0U�s90�����j*��[6�fb-N6��s�
3����R���=Y3�"��C�5#��U�47���cs�K�1��ϣ�>N��r��߯iJ����m>XY��t�^� "�����80TUəȫJ'^�)n�����KIݩD�"����a-�Jm���z�21y��첳������"tS�Ù����z���3�����9�K!Dmy��*�a�b��#�V�.d:r��}t�A�ܧ��~:V2�:��ԭ�9����ݺ!#��6w�W�@��Ϊ�<�C1����JM�Pm�!�z�C��Ӕ�6l#sޓk1�&�����tgi��K�����e%2?�!}kB 6��mς�o����L,��*W�SF�˅�I�DW��r�=��"ly!��$�?$M�*�
�U���L?ߌ]>g�X�)��!�2$�Au� v�2;;�.��h(���q=����iv��^@Q�B-P�Z�$J�h�(�ao3��%�;`l��8G�Q��Z	ЊPfN�eE�l>��>��D5�q��q�<�8S��g6ப�M_�@���lq��Ld��[^L$i��¬����p��x�E��}�D���,.)^���0��2|o{81�\���hӢF��#�cK�m�)�ek�8�F�kz)�l�
�O���I�E�E���i1�/�Q/�0��d���!��h�S���}�`��d���	��>�Ѷ�,�͏he��Δ�e��ֿ��� �}>�ؕ�/9� A�JO��U	�!9���ylҳ�]���`2���WLƹ�X�2E��<ZM�k���6�Y��#ȈER�_8E諂k����&<���pO�B��\��+��%���u�ݝy~nc����e'��o�$�tC�]��N����v+c��~!���-�y�C�~K�i1��_��g���~��g��bű����4^/�∟��Y���7�櫸�ۉ���O�_�����%���Z9�70.�k���dB��'T>�<H���T������ �E7›�[�p��'sS�`NC�z�d:�����QC��uׯ� �x/ 	
��V*|�ߘ@�k	�꺭���cB��E�˶���.f8��$?�~|_D+�D��}�"�孬�HKt�'����g�`b=���'Wl��f��'�"9�糴�R��If\'��:���"���N��g���U{��6���e��^Ћ>��(#F��lg�j�ҾZǮ!�l}�W�4�rJ�����[�G�)�[�/�Bl�#�d/��)�^�U/��9��zR�x�؞�����:;�VR����{^y��
5a��n�b��Y]h�z��[��O����g,���y����Ow,���]n	��=fo�*������g�M2�/t���_��!G���1��j��E�b0� h3.�	�S�����W $�#�%��g#G4bs��#*��ɨ��g�]��[�_�Cj���xa�Eq�`y~\2?��^*c5�ҵ���>�D��ö���=)�X��C1b�@Yxc��zϨn�@3�o��M���1:k�Vmd/�Vi�ң�7�e����Q�h�q3�L�G�2.S �qC�,��������t� sqk�1JUP��Z�/�^/�m�Z!_�s#����W�EU��Jv��I״����D�w�j@�~q��ﵩ�m8��J�l*��,�}�*$1�/�|wĄ��aE�\��RZ`.i(�O�R����r���<!E�)-8|����Ta�+��y�X��