��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�ȧ,ض����'���~c D����G�iR�T^#1��fX8GN1����z��٢�06� ���T�L�Z�:��P��\���(��I���{Q��hp��o�~�t˟��C-�#A��L�L��s�و�RjhKN�3sks�b�m�8�ȧ�q6�H/J�t��K�HW;Ģ7��\J���M`>� yA�\��MeH}\}�ҰF��c��Q���ai���R�]��^կ��a�na:�B*�SS��$VK>�L�N�o|R����2�.�[.�ѩ����,� v�� ��h�6�$������Ѿ�!U��*�ɻ*���c����o\��Z��Fm�_�$|1-_�@G�>9_�E��^��ϻ?G�iw'Ӈ�A�B��i1�6�D�L)�=Gn�8I5[��WLO~)�db�A��y�<��?��"s�R,�:)5/`�x����Jk�D���\�������RQ.��F�~�qvL�W��>c�m�ݖex�.�A� O��uD���1T�����_����{��"�^*!�B�Ԩ%�&���	:/�Զ�~�Y)/�s��s�����6��)��n`�U�~���z���_��W�}yg?k�#�� i�o_�Ch�lɝ>�p�񰺥1h�W�"�姈�J���"�p��G��_�4j�."�V �C/xm1d7F޾.��,�e�S�@ ��PSV6�b_�#�,�+�3�v���m�4E-2�e�V�L�()���ېl6%��^��O�8���q��WӕMWJ�H ˹��P�n��ڙ[��\7t�S�c��!�eL=:6�s^Δ���"��a���_!l�^�d�Ws$E?��Ԁ��|����KG��I4q�hO�Q��Y�y�����Ga��V�:4NV9o)��G�y�r>���БZ�(OM�t�L�ж�z�zk���R=Og/��w�_(���K^��Y;|��g,�6���ׅG�5
=+0����ԍAW�H�E�ur=>3�k���4UWT�:#�%���ܽ2�!������a/��ׁO~W�C�4�fT�J�,d�s � +a����Q�s%'�jm��щ�4n�Õ��\�Y'�:ui�t�sv�i8��@���X>s��FsV��8��J����ƨ^Vo`��0]ۓG`�� �T�]^�ٹp2d�i~�O�*\�݌(��=��[�m2�6P��e��ǹVG�#��� ��D���Jv�~�&=���dm�G�)9�'��-�P��g���:�����
6юh6�S+d<҂?]]	�-�4Z��DGg3�ϥ.b���5��}�U��b7��	�)�&_�A�Y�B� C+��,ٜ�:K�mK�J�ΟLI)�We��gW3�o�
٥��e�/5�>��o��N�$�0	R�����%!�e�&�������}�5C	EƈNWV�"��|��	�� n� ��м��s�/>_���?��0h��mb5�MDnm����X�$.7a�^����[k̓��<�޾&�k��v'�S+Mw�����s�Vx���@����gD{��o���!q�*�PbR�GDSY��T�F:�Fq�	�*%FӅ)��&i�뙂��`���[��v�]�zR�� �$��Z�6����3��LrEd����r=,���8 ��-Y!��"����ڪ������S�K�҂d+S-�����<x����>�Ժ��K9�$v7�_B�ʻ��{DD)�n�Լ�Ix�I�[�G ��[�΢�ш��U��WA(��n�٘�A�{t�xu,zL��z>D���W���d�C�͇D� ����I�w�:*c��J��{�� ��TBŮ���	���^�`���V�HI�����~1���(�X�fa>Gʲ�am =G�"��rGh�D�3�gUs=�4 �xC�2)��N�Q�.-�	š���F;+b(1r��K���LZ�
�?�J�Hm�1��u��?�Cc����M�����9��N�t��U2o�ɢ&Ѫm��SP�Bλu��I�`w�&�����f	���v�%�a.��;8,�(���:��1�^>�.邎���5	!\�L@q嫹�8Q_e��1�`�$��&*=,Gu�^r?��~C���VVV1����u���âa���=��U��S���"Đa�V���qV�Ŗ�bMFi���VG��(<�9���h�ɏ���;���T���F.�('f(I����Gi�hIF4B��$��GCx:��q ?�ߵ�L5GQ���'Ƥ¤��.�����ǆ�^0���'|��+��7P���ub/�q<��U̀�U	�K}������K� ��h�
�|&����=L���B%�k��j�K	Q�y�$��Vq	gy���2V�X���sg��_s���o^M߈vxlD��њ/vk}�f�U�l�*U�K.2t�w�����}�Bɺ� :}-3v�a�r�%��GH��??�6:�d3p�5�8���w�=����A������Z��O�X�}a�-w���-�A3�A �pLl�����ErI�EXt�Sן�awJ����.��]c*.�<ܜUx��ɄE�A'eS��;$���m�p�mvK#��k������|� ��gv��+�EI;N���;��1�	��URE��U	�PU3���\LP+��Mr��<���E%Hc��P�����?�pL�Q��]����uW'UP�ޯ�����_2B��j|"V��
�}�N�� ���Z<�g+�T*�����O��=��- q����T#w΀��.��í2/hdN��_* 6WY!�p�>�W�w��[�٣�-z6HS�Oq��!k�(IR�Tc�R*�Π'd�)�#��V�CE�`�(� ���F�t����ʉ��v��A��C a (I�>��GO����	��evZ��ñZ����h��/�	���m�k](�x+��~�6k��s�/��R�j�}O�xL��"~�ֿ+*6ꏕ��<l��񓭡�/d0��d��l|�0��@����Eo�<{\���
�kD��h���׀��bZ��U���-��o:(��iY�d��;�g�:�����@�"���C�E�� M"_�(��Zq/�*R�l0�N2)�na<�� {��Dy��M<�$Qs�C(g��/|�� p;w'-YH�ϕнa>�GH�f_�j���YONy���Z%���.!�U1X�h(rVˢkic[[<��<U������ۦxHX�����^	QQ������3៻ʑ������m:H`��|�t���8�����q�m5�������&R������i�ͅk�q�x�v��� g���vQ3C����Ǳ��ѳ�-�(�L�'r/�;�VD�G�@r����>��S��L��_s�Yks��N/C��H0f���wn~� L�Λ�Y��||����`��]����Q#� �>U�Sh�-S���s>�t>�ۂ-iv*�+�� s9]鱍�����q7�;d X�_��������'<��-��>���=>������	6h��(�/�'T��/0�*C�@���Raq�ِFJ�ͥ-�0��/�!����Ĝ���-�-����`���HSEX������6�Eş��c {�l���P�|F�q�27[�[H�Vת�܂�SE`ޓ#>3�щ��Y��xr��:P`/�̀�-O��EN%�=f�����Ѣ�儈�I�3��D^�)��s��U�:0�/#�ېȦ4n*1z�!���`����=����{YW�9�I��fLJ[B���ȁ�J<��B~��.s�\��P �7A/먜űy2��2K��%�ò���`�m�~�ݨ��̘���Ʀ�n9�Z:�.�꽉�����^Z���z�&,m;�Pt۱v7LA&�&�Z��ʎH���
��n��v�
;u��z��"Z�W �o�'?A<o쓐��
B�ˠ9QmO�{��;�m��i`Xs���Y�Y;K�C�Θ�̴����N�8M�����d���e���rN������}�?H������3�`\�hj����EUDe���*}�1�Jم��S���J=�,�k%g!�/!�����I0��N�-VS<�2ܜ�3l�s��V͆G9���
z�ҍ�o�F��I���k7�=p?����9�����,L�@��Y�K1��7X+��6\e*Zæ��,�IRhwu*�����j]ە�D��G�k��I�X������U�Z�]�
x
p�t�/z�~�Դ�BtF��Y�Y~}�^B�?F�dW(�y�Gb��Vv|hc�r�Jb';�"Q��kll��k3��*"�����ZE�|����j�[[ �t�+�o�8!��S����V%����N��)�B1�kN�#��@b�^�$Tk�^�z�U6ظ�<b�Vk��԰C?3b�^���?t\�.W�����w�q���2"��~5�Q���i��GY":���W9d^*s�CZ�5�t1�*�9���+�7N Ձ�o�{��5��Ƚ����Ҟ�s/�y�Ћ�rW��Ks}&�/0&���f%]u�hƹ��3Sԇ���fӓe�"�����=���/�h��91�2�8��n��U��2��{�͵�n���ʶP��yy@�\�wTρ��^I�"�@x#��|=����,c@Z���_4o��|#�oj�,�Z�O�+�>'�������k��1���cۻ�:�4�������x 5�hv�㻤"�Kݸ�����$��'�]K��	6jP����7E�]U9�zXn\�E8�Z9�4��m�y��P�c�9�#�ҳ�2M�MǼW�pI)\2�A��z����K��_���0�i�]%�V�$J�U��%���0�����˓�ɞG9a9����
���` 3+|��51�&&�-Zft2.u1���,���vj�.�#V�a������I(ݨX�:>P]P[%�U�_��I.� ���8b�#��0����G^�t=�~l�呋�>�[����{ �e�؄m������W�"��w>0N��#5�(P�~J�ĵ.�B���J��f:&	�l>�D6A����x+��v�W�~��&�<�V	�!�o݆�Q�a�y�`��E\ru�Fט��[h}೜g!�b@�v�V����K�\�*���!��&�e�:����k�?`�/���(e�G����0��6�;�f�7f~�2\&��8������K������%�����7Zj�'M��{#	�Ev7p ��V��g���	��TRJ�Pz�wJo�������]B������ǐ�x�EQ�&�A�v6Bn���h�q�p�d���vO p�E�X�wȽ�C������Wmb����Y�<SISy�Z�uCA�0����.g�&��p��*F��C����\��vR�}/ e����7D�5}f�@d�K�?y���'R�����b�$�J�Mт��f(��s��S�9	���S�f�Vp���̭�.4�1G�{-�+�
t7�n(��t{�-����z�>;�� ��`��;\�A��ᜌ߬����2?Y��u��=߆��He��!��L-jA�F��}4mV 	�N�-V�vY�g��\��b���{��>vhX�gѹ���J)+�h!4[Q-��C���`B��9���5�E�vb��?�=��\5o�_�~�8�w��x*?|lu(Y|�Gp3��P�� =R�l��5�"�O�m�3/K2y�sA��'��}$�*�Rja�D=��#�
r|��U+�^�POW�T���r��F՗��>JjL���Z�aM��&�R[a]ʥT+�a9��߼�K���yf�Fz]5�������S������S�5'R��V�Y�?ju��D�'��|�����d�jpHzP)-i�9�����NL��BHrx��R� E��F�N����F���x�`��Xԥ�s��� ?�I��������M3�|k��v�~��p[��n�!�U���#<�G�wKc_�T{�{�r���VO2E�����o�k	7�7�1��ӻ��P�+�dW��l��8�٧6�`~�Xǲ4Oב�#܉����}0$>od�O��E��� Ŧqqu?sg�J��sHq/+擣�Ɇ���1g�!Bd#X#��]�����ߪ�SHS�uP&�X��GV[����u�B�J�)Z�^�4�$$�-�k�#�0޺}����_���@�{[� ?�:�c�K-��M���S��̮�P��FUyiZ�]�w�h�GZ
��:���y�8���]�ޙ�o���k��(�A�q}SҞ|"�Q��w�û��v���q���3|h���U�]ܝ���,��YI4����tv������U
G�:0�����d���z��*��0�Y��V��)�u�EY�p�H�<���	C���'u�k�  �Q0�[{���=D��}�y��Hx$w��b'�)y���ԗ�'R�%�c=����Ӯ��b�ay�i��-�g�U"�U7�BETh! =�o�a<s���A�8(I� �_We/D��~p+�xk��!迺�Z)�e�m�4��4CF�²�� ��{+:�0�6�_�9��Tӷǜ����=ifҩ	>�O��FEc�������� c����y���o���C��mI6E� ?
�)׼�[0�X默���>������B�LoV�L��۵��E���EW	X����O�op�'��0g>S�c�� ���$J���e�N�P�iH��&��Y���������pZ���T��Vkk�/�����ĝZ��e�Y��Ϋ��,�m�q�?��N4�l&+���+��1l��t�)f��®=���Q{�&;Ă�y�/@�9Mb��#��j.����E�.H��qV���D��M/i�*	9CP�K.�m�7gG��u*��Z���+�~C������WXx�dj�(�73H��������a'�"!��*�rP=�TM�3�t���"��Uc���𝳬cggW�(Pi@�D�&ú[�ib�؃�����	=�U7t"�IX���M�tɍGF��	���C�W6�GB�Ta&�4?���:H2����zo�/��;�!�C��{ľ-��k�~;!�HN��_Á�W��ܢ9	�;�`0�@_�y�q*��M�~A&Ĺ�Jt��.dQ��p�mp9��i\�W�*ܧ�Q&֓�-JwR�/���T�u�l kj���"�W�Ab�O|��ԍ��FUߙ��F�F���[t�~�$��f�Eo��{�ml���]��l��L�P�w8n����,:�
���.�BSdN�8�յ&��e��͉��䁒f1��\�`(W��cމ�Éi�v�za�% xk�WR?�Ǻ/e9<��5�3F�Ԓ��2	ky_��h5{��pڿ&�rmH��ppH���\�R���DY>c�T1��!��pղQ���y/L���gL���QX�z�=�yP�W�`�.f� ��}ۿ��a���4M�.b��M�.V��Q�7����r��\<Jy�c7aR�g��������6d�����5���z#9L�(1�꫸����JK1���A���Fj��Q-�ƌ���+��v�}D�|��P�Z�'�lN�Yc�Y<��Sx��HK��ޛҞV��x�: ���A�� �����3��_�����1[��~�֠L������(^8�]�=�xP�\�7��AL��O���#R��� p��I�Ӛ�ؤ���&�h���!
 �w��9�JZ��z���tW���iW-R�kD��"�Ե.#�)rn�(|��2`����k(�݊�[B�ЕdO1�,��(3J��8���k��~nD#��g���N���؋¨Q 9���-6wR�XF��hΐ�W��x��n
͔_��|�_˦��V�f�Z�b%OE�^T�{(���d��@�4�٧���w�{��w�� ��-|)d���eA_=|t�.�m�mq��F)���!��CjBi�If��1�������M�;F�a2�^�IU�sR�e���*����2V4�CL�щ�O����%9�s�k�ff9N�[G�n��b��oB��T����%���߳:�1-,X�B��n�4r�O�Md�������E���dLVX����*��r9�S=']T ����h�~�-iҞ��!$_��R�3R�'X��̔/cq����� `���lf�d��gK���q�$�6l���mz�D���S�<J
�
1�MO�t���( ��~��`�{H �j��ϡ��~렸Y�IR��1�3Ut�%6ה�nMV��e)d�Dv�i����1c�� ,��x��b��#6�55���c�+_w*=�X3�,�z����] ��B6x6�]���"�"�yך4هV�I��&�}���r,^��I��P|���t�K�|�5��3�z>C����{����Eo�0X7��>���n�hI��v(�Wj�&��Z)��5 q )J���i��$�w�h��۝���b錽[���x�i���u��,T����I1Q�qʹW!����2Y�P���{@sanP��r�iEa���f&=úb=,���6Q"��Hف�K�&��`�URy�(�ģ�6g��C�z�(��up�[}N����*I0$��������Yq{�������p�[�c��o����a���1��,������9���aa}���<ܭ�������U���w�q�$`BR���>�w�	�Im�x̯��F[�z�O���5�
���ՠ�m�+Gy���#�{���V�6���3�½�"�Fy�pnb�m��Q��A �j����*F��m3���Oww������~��d0}#�N���W= h�I	Sٖ��f�$��@T$������\f���7o��o;f���B-�>x��f�]���ԋ��ރbM�hu�DQ���F�ΐ@e�K�����\p�ku���a�b��6ES�h.�|�' ���-H� ����@���Q�\�q�G���63�0�[����>2��Cpp$��R�=���M��KZMD^�mq��Q�N�[pTʾ�ʟJ�w4��Y�[sC�w������7�4}��4����.m%̥��c�p`�;�ZuJ`����\��4R���P��x�ƞ�
!�^��\D�%f$&6��G��5���KD1�.��T��4+E����6��\-Y/F�`sP��a�W0sg�B�G\�U�F>��fm��&'�5�J�l�`a�ֿ��<�|��l�[[DKx'� ���ꉳ��cN?��Fn�C���/��t{'��Iޠ&��3��#� t��!�T��)eL�e��]�˓Xh�k.�[��k~�Y��Fϣf���v`ᑁ�����!�YaI�3ϼ�P���ٷ=����'�j&��чG}�J��`G8鍀@�<���ա<�b1U�h2��4��w��#*�nx�*�R|\�T���/Rj�5���2L2�)�w4�b�n�Bp��-y6���hcA�gW�a[=+ğ_Fi	d�G��#	���[��2I�ݮ��"�LQ��o&7[%�:ʰ��H#&o����i�Y�=��$�|[��^�S�o�~Φ���oP���ޓ���H��)#��L��������T���N���(��R����?d���L�c���%컄�i�#~��
ʋ!b~^��t2m����܍;O�(��UI[�[�U�ؕ�%KuR!�lŗ?>
��3+�sQ T����e�50��,�Zg�)k�XKi�5��b�c�0,�xXbź��]'��J&wU7����c���Y�kn���úSk�����'y\�ْ�H�Y��ы�e\����������8��C(zә���BwPT{���#rIQyO�55�'z�O��5p�P�R9��s~�&��j�.H�����u��.��
Ό���8�;�7�A�1ş�t=x<���gk�Bz�^�T��H!���8����Wg��$��R@Be�����s᭯^Й�ݠ�~�:��L�u\̈́�kI��L&�+)�TXE�V9�v
�2ソL��;���=1��e�)���E��@q��6�����=���j�{&�/��9O�=	�O�y�S�����,���8��a�T��\������Ĺ�F'd���B`�
-�\��^�?���b���]a� �;���ѓmc8�n���-P���ؠe)�x>�uKMP����lv��o8Tfj#��'�SEr'�������0t�[�ܽNDF2�����g�~kM�ho��Y��A�7
~�ZSg��WY�rW� �I۽�NOI�sE"�KuQY6��v��~��5I��ox����_��03��y�P��_��<*�xV��Ў��=�tk~N�ʉ�X;˄�����6�V�5�`�߇�i�ۨ�>Y����a�ة�-���k����
z�����|�f�EĘA����h���g�W��4�o[�
���H��0WF�����!<.�)�Q�a+��|�\q�5:��r�!����<ڸ�h��ƘH��!��ְgz6aN9������_pa���w�����m*�EU]�/J���V����<��>ɤ�|7�x(l�G3����ԍ��j=��S� &CW������"�*��H���E�����{Zm�K8�5NDU��48�K �:r=S��ق�@Cj�u�l����[��T�m;�T���$ǡJ�(���'#F������=���3A��u����xm�xdqd��r�'���(�I�K�-���Y���Y�B��ۅW�O2����l�Rs�Ve��4��ꆓ���V�"�J��â$L��G�"C�è���',��w��m\-��=��T̊H�C:8�oP���B��(`���.�2B��$�p�<v!���t�< �3��D"�˳n���Юz�uJ-���W�R^HU]��Y���}V�Pxq��^��d��O��68!�3*�Gh ���i�d,���J�4��ِj�����{��p8ճ@��$��ʘ�Kؚ��o�{���%V�������U}��[�.э�?1B9�b�#5�)��Hq&����O�q�O�e�E��#�N��G�WKB,9�+��qA�@�ڏ hL/������K��аH�Ǟ��!�|�����<�H ����b���r
����v
�vM!�"\�^��/��d�έ�ho���%��o
���N�N�$icM�.�Rw���W��"�
6�Q�$g+�i&9����dj�ϕ��m#.#�B�|�n��Z��y��G� ˘������y�) ��N�a��ˇ��+���cխ�����vn!T���t�c�93����9g�3"Ty�C�~T`r]��*�kj�������,�-BJ��F�~;�z���8�E��+іuWvX�b*/�_	�� P��ɲ��Wgڈ�'~�9��=V aj4O{12z�~�HΦbi@>%KS�׎*�#!�E[�Ŏ���"ë���+ �Z��)���V���Р��C�u���2��7�V�J!�)��
+�Jx�ϔ°ùj[��g��xo+j4��9�'�^��	d��O�N;��
�h��Q'C��T �rkT�����#�)�,G��;���.���Fx��jqFRah�?��|a��4Z�`�n�׬i���>����fkhO�k*S��I\��옌k�ľ꩷���1HѴ��rV���r����FH�?��s+�P4^,���)n��
z E���q5��E@2�j�C�cM+�W���|&�@5k:����l�݅y'K�4˱�3!��NztV�f#iCܶ$S5.���y�P#�H;�[�_!�)�OҎ�ϸ�0���Kp�W�B/䖞9t��jx:s��f,��`��6|����z�,Ŀ���ȼ�^ߩ�6[3iO��I|ݺ������'�YfrƲ���W�6��-��4���p���6�uy3bGt-a�y[h5�B�	0DU:l��h�m��ل8��w�<+�+tA� Չ� #9��/�x�21%��k�0��]ad��M��q��N]^�O�C��1e��㋮yw�_U�1��e�`�D��M���>��t.0���a\���?=c��5��:�t�t�Nk~��.T5)���C0ѣ�:�t;��|�-3ͫ�58
�+��$t�&W�'�
��tgq?�v}RS0�#!ビY$o��?�c�؋��1lY`�t��԰HiS\� �fu�fOA��u�@�1��|����=d�.�8��3��@@�ö���ZX�����!f�3�b�J�Q��1�0Z��Jz��j�0�Y\gX���oL{Ƴ3�ڙe�S
s ����1|��c���P�Dގ[+��X��� /)�F*��*_K6x�����ۍ;o��!�Awޞ��e���i��h{5.�yein�K��z���m�dU�:�l ���Q�󅸴3H��=]�[��>�	��,�#��1�/xB]<�D��#��
A�H�`����X}�&��8�o������U�[%�xx�b�w���OJX��4lҶY��
�v����*��>L��F�fo��w[�ٴ܅�k5�(��֖�Q�Y�����23_[�;�l��M��i��9��-�����A�����`�=����X>�T6�I�~D�8?N�����㨚��=8�y���c��Y����M�t|���'&�H鄈8��w�g��&R�Q@`��bsB�5!���c"P�l��(�Go�{j�J�E�W��,�������m�#��B@%�G3>���o���7-�������x��)���_WZi��@.7��8�%���UR�S��4��5]:�����;��6�T4�)2#ǀcc��X�;M'z��Qu1�z/�Pm�@��gt@�T9�����B��^�.^�>���J#d6|MGނ���Y}�����6�ށz�l�Ru6n[����+��It��ۺ�}j��.OX�
�._-�'.]k8���ޏI���}�e��Ȥ.'��w��h]���!�g~e��T`�4,��(����������枋Q��ƣ�`�X���J�aG����͈���p��1��Z/�c�cMdЫ"�H�?�����|���Op�nG�x���L��V�-~-�3GP�y�Z@nc�]����y=~��\f���D�+�5a�h�ϸ˪�X8Q�U�S����M�+1��%U���	�~�!»ɋ��.��,H*;��J�tv�@`j�Pӻ��ǀ�]R�$:�f��]u�HRՋ�Y�
Zs
� ��߅��a��0��z��+��)E�%,.��¦`:C���1ѡ�@�,�n���� �O�_��B��)n�����qg��LԮv�_��z�TQ�c6��l��ߎ'j�Ci�\�ꐥ0h��6�U��y E�;� %糲լ:�f��] �;׊^K/�~���φ�4t�t>K�(�\��Z/yJ�ܸ�Sz�n휍
mG(��<m;�v�$�N����x��F��bq�^It��� ���5��XAFn�pU޴���A&�C!*�)�u��dN��lo�����(���@=��}����<���"�����;-I�ݗO[Nkx�K����*LIAm:�*��4��y_v	Rw���������##EJW�r���5 J�M��n�{W7~��|�'/���}&o��&�K/�	8���9�",���ځ������ �q�YH/*�A�d	�}�oB6L�·b�c�!e�0F�!��������9�ٷ��}��2aJi���ҟ|3Hǥv�X���/��pm�1N�%z������̕����b����RU�BE&�NIjV.jfl\��:�]A<����J9g_��NH	짿:f}��Л��	��h�!V� ����غ[��X�������|��bM�>�q��)w̻L�W�=Փ^�\"� y�kw{N3���P0hNP�?���'�{������/>��I>ău*a���؆�ͥV����cwXK�Nmu`�JZy�e�kgw
m�r��>[Exv>9�����&��R�����c��J#NzI4��{��t��Sn�F��\�<��M;$�#�Q��lňb�M�ʥ��>��k�/��ss��Qm���xM�:hj�T���^�>b1�As)*"�zn�� j���q��H_���&W��S�f|���@�ඬ�E�p�1���3ܓ0�V�x|t���k&/�Ѧ�=��-����D�n�ˢ�H6+"l����V!���p�Oy�В̘u�����R����jڰ3��&�u)�7�IX/�E�KKyf�}�ә�b�{�js�����ޖ��w��7**'�����s�ZV�'�; 6H�I]��������dڵ����2�P�����Տ({�����'��[^=�(��<�mt�:�o�-B�,�=w�F�I7�l�+G:��A֫�� � '	�x
�Û��d�E�����V`|T}?c"l�?7���,f��*h�M]F��N���;&#,�7�;��ކ�jx��!:T���7E���'��̳Aҿ�f���Z	�y����u������%bp@c@�
u��0Α4�լ4���m/�(2��6~�#�b��E��؁E�XQ���=K��jIh%�ZF�i�d}�m	a��/b�߮*�ޱ��]��k@���KG�S����O��'Q����bZ)����>ce��6Ч�%���볶Z�۸(�*_f=�d�J����J������F���o�|6��M���P_��2~8��O ���!�߸8�(d���ۨ�2"w��P�N�e`u�BEþ���W�EI��Mt�-V-?���u���TK.�ȥa�3Cg��+d�]R�����@���S,B6���3�̅��[U�
�$�jUi���t�1�;���>?�JXH'�;g��<f��y�BZ����晌�g��s���KE�צ=��/��JO���Рr݃q��ފ����������<?��ݑ���փ�T{9��#n��]ȹ'���n&`�H�ήM��>�{?�C�n�j�ee�� ��L�)�<>�_7��� ���i��)B��O����r���?��+��b�h�_�
��L���NB�A��'��M'hfheH��*��__mY���]~,V
c�æ��L�z>,!05o
����y"�nz��^h�gOIL��`Rqx�B�Ql��IѰ���~4�5O�3�"欷�)���it�ym����`>t�V���[��d&���P-�nZ	ǁy�P�3�1�t��U���6<*��+!7!�25ēM�`Ҕ���Y�MZ��1��b�bi��Γ�l�B�2?���-I_��)l*6�.��/�/|	4�i�_�/Iz[�}L�+V6qi}��d�;=*��@7޿#�u��,$s�8z�-��Ӑ�y8����=m,����A*I�n3������#�ҭx�+S����$}-�8\���4p)��k9�,��$(M���r|��_�����G�v�~l�"Ľ�Zw?��KFz�]�/�-�rk7rp�!	�������:��l
�@��)���U%�q|��b�n����{�^�@'��f��Q�^�#qԴ���7�i�<��������4�p���S,4=J%	u�^jU�ݐ���YO�z�6-k�����O^%�f��nRq�_�#j