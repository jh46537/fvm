��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm����질�95J{۠�`\j��G�!�<�ց���&�l,�y�ʰ��D����&��ejP�4��:�D�BH�v�Y��0�����"J�������W�#0���1�Ay0����+�.��g��z��Peˇ�;.��㝨i`#��3K��o'ͪg4��T>׿?^Ti�j9`��j��#cu�����vJ���J�����|N(�on�@u��w(�������'9����'�(
Lh��*���ù7R!�߹O��l��~J�v�8U{�P�{י�-	�3M�b�s�O����	z\8�L���ĺ9�!y�9�R�$eH��>P���1�?*
2U���W5�҉���<B�vj�dW��j+am �Y�23�]�����;�K��Xl��!��]�(�S��Oe^���%��)=��x��@�@�@�WvF���d�➲��� \���"fK9�'8�}�|C���a��"^�7�pF�y޲�ǝ#D�*�¸����g��GPV��ֻ�ܮ��W�۷Y�=���n�>K��W�8nm=�,�a1��,@�~B�K���Ƀ<���?��g\b���j��O߾���C�%��(����ɕH~�z�8��8�)�����1��U�%���uش�ځ���6-i(j?(bK]�� ps�A��fK��XH���[4&�_�~_?��%�@�bf��?:l��Ig"(8?@Y�UzU;�h&������mܸV�*;�ƒG�ڽ$6߇b��[5�����P��J����m��V]f3Z�=
�v���^��u,!��rm;��f+̣~�R7\�;��[����]�<bf��lS�b�F�RV�7���j
+m���c-�k��-@j4Y��0����2��UHXXb���ISl2�����zIi3�4�|� ��7��ަꂅ�����]�[&�?���S����qyU�����ek��ko��d�g"�;���}.�Ha y��f4�`��{X�1�,Ȱ�¼z:�i�<3l^��Q5�hU��}���d��E鿮���Fڒ���4eO��s��P~p� U9�	w�d)�32U@�h���p?L^��s��3l�<��R���kj�܌f'�t�����S��S��㶓$aqy��K�7yk�Mv����B2f
έ��Ef�#�Kk�*�Fܣ0$��5����S�kp��,k*�tc;�C�-�n�#ۺ��ܠ��𬋒�%3W6�LA�l
y�>t�%6�dz5/�������]����M�z��6��k-3Nr��&Ł�]ϲ��%���
U�jP!�<�r�O�<���#�$�7���KE�����^|"�'��H�X�	�2�Z�����F�����לT�n��])��{C)�1�E>� �IM�|����L�b �H*���ZkB5t�$@ZW�<�{i!�n�h�AĿ�"��ї`�w?��h� -�����	rS� �F
.3h��2�z�֨��k��$���.��|��Ł�P��膇8�t������������S��������S��dZD7�i�W~�p:H݄�_��,H���KD�]~�m���Ԁ����$���y(�f�G��J};׍�)޼'��zK�����U"�f�>�~����z:R���ӂE������g~�Y�V���1���M�D�TbM-,RÔV+o���a]����aIS,�F:�e�^5�Ժ�dY��f�P;��"���VH����xd�f4&�_�8�	i6�����m�rκ�k3��K�H�LFɷ���*'��X�;3��`�}��ִ@Y�Ȅ2�3L�cM���&-���s�Ö=>�V��i��ʥ���J֭�f��@x��m�5�0��&"�h�ӣ�,jCڞHf]�b#+db�^�h
(� �� �(���S��k����a��E:d��I7��=<��	"Ή� �D����sQ���ҹ tz���6!N'QT���i��5Q�B���BtM3�n!����VF�c����a��l�-�ě
�B��X�yO�V�������;|+@��4Ȭ�(�Aj�9= r�D����OW�����Ɇ޲�p��VO�_�a�3#zR7�j}W	k;�	����ß�n4��V���Ϥ�������+�;�o#h��nz/���̅4�TsRN�O[��U��ڳq�h���\1t�N�1ד�fl��o#Lb㟉���^�=DĜ �=��e����S�G�k���b��P��_�����Y�ҝ�u�b��7�uQjN)5ɢ ��a��AdND�pۘ;+��{hf#��A.����ĥ�M۾s6�/�2>y��~Ү�s�~�c�wUwKRp�t���y楘XQ5����o�g%�#}B�,����40�z|wBP����u���Q�ޑ'��2|���j�y�.sj���pG�i.��k���}�w8O�x�Oo����e!�c�:�nJ��+Tl,�^VDQ�YTǠC������N�Ύ��Lq��^�c�T�ӢL�@¼�p����c�����
����D��ӱީ�P'Y���ٔ�ua"ݝ������ЄhO!mN��5�x�[�Ȳ-ٓ2�iU)kj��� �*��<^q�jJ�m��$�I�3w��=���F�ç��uIw ��QA�����i� ��f�F��⩖�= ����L�{k�"������Fq�����ʔ#�j阡<.��TL����v������#�����ݟq���:}��"eQpmR���>&.�ۡ���h�%&`��\��c��A�c�)�����l.��d+�������VV��+�z��r��/`A�1�ۚtQ�n�,b%��:������J�7���Fr��9�wJ#��Z����̺��	P2#��k�2
a�%�F$����܎�~�Ki��f�V,���C]&8���C�� �p�f	���wRǵ����) ���1{X�^:��EF�ħ��<��1��q��V��O�S"���>�W�v��3q�w^�c�ǘ���
= �],`j����8�[� �W��� 2�Hd�+�?�J���~eH��M$~�׍*�g���J�$�U9~Ϣr
������J�h,����[�M�#�D6J�e�d;{��ƪ���+~y�\��#ؕV��C.�$Yh��F�m߻�;�S#ޚ����ߝh�7�Gj�9��8_����p�a�33��.4�K?.�������}q~�`������\� ��-qZ�*f����m�
P�rQ�_sLNPz�������"P��u�i��IثM�u�1Q{�i*6$��	N��a@*���8x�;I���:�cS?�E�҂|4�X�b]�8�7Dp<H\菏�Eg��c��y6�+R�Ӽ/�s�?��Κ	�-�_'%�jd�zG�̙���a�$�0x�r�EѮ�=�_�\=d���R&h�bB}6�ۉJYn ������T7������L��dp�g��#iȠ-Y���A<� �%��7�/�X�EMu2���:��K�R���6}�(R��!�5�v)L�
P�O�N���A@��a5ދdN=��Ԁ��l+&�@��nr��ؑ�Ɔǲ�Ej�$5�Z�e�?�k�g��#�w#�FW����O����y�ϒN:L��Y ~�����(?��5;����r��$>D6h�	��O�Ɓ�#��Ї��֧�e���ѱ��'v��0��dc�K��ˁ�IRݭȆx}?1��CH7�a��a���2�'�������$�����P�7�$:��cy5yHf�����*��5���`7onз,�O- Tn��}�PV��3���e>�oɆ���+Y �WW>#�Q���J9���V�v&R�h)�38y�L��}gzk�`�<lf���?HiP�A�<j�N �~-��'߷��ҿS�������9#Њg6㱗"L9�φ�%(Ռ�g��TԲ��,?kP`}<��|/��5qO"�Dh���m�j�r�CG`If�aI�/�(�@lKveX�e2�_p�℄@D�'�� ^fE`�G��/h��T,�� ��PJ�iS:+�룚$m)
���4,8�|c�Y�<ϸ��
9�'
*JBQ�ǑG[2��� �Ff����� �u��QEm�&r!�2��C*,ޡA͜eo�,��퓠��0��!+� �~��a��*AU	0X� }���'Q�����/��'�K]t�vZ9��*�6��p6��V�"a`�'������r�pd����_ E��{y]ߘs-�v�m�`r���r������#�I��p�#�e7/4���@[�����r]p�L�<l��{�}����/�5�^j�U\�%�g�y�*���z�e����3���_+AQw�S[f��^}��G��N�I��X���F����v0Q�.h�k~0h3	�a"�.RMx����h8k����+��/��_�+����1L	ίֹ�<��n���G�6V
�u>�b�mޕJu�p��0J��xp�V�-(����+G��舐�����H9H����ܪ�w�R+���� O��k؀��amH���Ϣ�p~�jAY�TH?la���r��@�o�J����F��ö�4��)����i`�p��N��,[�6S��nŖW�Z�k~�f�5��#�B��!o��.42.���K)���R�ufߥv��5<C���&5_�3 ��`�<�#V�=����.�=�Q�����Ӥ���.��ڹv+��ѻV���+[e+�������y*&Z�҉�!0��� ��Gõ��oL�� ��N���r����.�免�M��wx�T�id)��r��ψ��7/@0y
��m�5&��^�q�GJQ��+��6֐JMf��~����Ǡ^�����΀�ɜ�OX�+��")'���*o�HI��Ns�|�V��ZH��=�\�K��]f��s[I��m�+Y����X�w2|?H��P�J{�Ly�����(̀:0��I��l��B)bt�/�r�N��j˒79�&�f�rS�2f�(Q��-6j���$Q�	�8L"���t��$�X^�����B��~�"�P:�?M�����}�����SM�B���
��'U�b����f2.Z;E�/c+��(f��FPtb�t�c(�"�-�G��A��~���o�*K��W�jNW�c:�&�����۝8���5M�����[eA�H�~�g���WMW�#��PE��W����;:ןy�}5$�
�(K���ZW+~��/���4��K�rǢC}]}��.<~��T����B����h�
4� `�`	���h�iS�r�)�1bExA�ڬ����EU���ǻE�TD:��X�A%���4��	v��'�aE�_�j:��_�n�֭��3~H���pIfG�@&W;��r�+�|1{�xݾ�pN)Y���Pt�-��,���,�h
B�͌H��~Y�;��~H��c�w��WJ2+�]��z��]��W.��jŃ\� ����U��
�)�,ө@�:��J{�|���x�N/���Q;�=7���,�z��8�_�&�x��5tK<z���Xԋl��FK"~�Z7_�W��w��5+.�7[�ʾK�آl�9��nG���Q<Ϯ?(�3�bt��rsW�R��qtի:m��;��{�D943�c*�?&��T4�_�\h�ܜ]�����ʥY�ߛ8�5휽]9(��a����_u5z�![���t�?�S�P|YRQ@Yɸ�z������Y�m��=Z�;$@���^���1�?	�����+�^�⣴��R�XrM��c�Ҡm님�FTm�&*��V\��)
�:a�|2xn�2Y6d� 2��ڪ!f���p72m�7���j�S�"n�j�J�()e�޻ē�Ǭ����:~	e���M(#�q�h�������w�
N\&-�lx���d��ܼUmI��ĵ'k+@z%� ��_7ZE����٫�2��"p�C�ѩ]enĎ̩M��+���}�{؎BIOoU%@1��1��Lz^�=/�,Q�#�N������n.�̥�M���B ί�6�� |{�T�˫"b�v���Y�*exL�L8�2p�$�y:������[���)��I$N v�|���n�!��Mi��rm��.@�Z�<p�)N�Ak�^/�@��6l|��/Eӝ	yS|%��N�{3�C�?��G! иd�=�� ��X�jxׁ��:{)
B���rQ@�A�]���t�E��Xo��wZ!��G_(��BO�n�r����W��+���H'�ܨE� �#�y���їT�G@�'݄=F[������,Ϙ����OMV������Cr�R:wn\�9��!$_Y�2(+Z<6ˠ�CȰ9G�N�� c���v#�g�ntLo#���ٗ�X���$�x.'.n��p����^V�y���2���j�L�