��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb� >��6\����B{�d�`p����-�'m��)p;�w��#�A�s8�r����D�[�~zIۆ/�����4��>
G�)h%�Ԇ�'����m�`��&-�ٛ�I2��b�����C�&t���K�"hy]A D���Ai�$^r��D���atrߪ�$[Yo�\TW��
��,�5m`�a���6�e��>�М�L�Nσ��ʲ��N�|�}{{xDi�M�6%|l(�΢�g�_���g&��]�[�OGnl�U�le.=��=�dVƔ�t!�����p96����?�b;�d Y�6n��mW�3�;�X��na��ў�R�
&yK��J��V��� ��\5 7@��:Zș@:ſj�W����%2ξ�i�%эչ;��a�0��_j����
�	� �+pV�왗;%V�(����-��,�r����·)��[�ǃ>���#.|�qN���1����tUG�.�#왗@��z��ϫZI1Q�?d�L�+L���d������)��8xfIC8�~�[3+��y)����?|Q����9`�0�6��
���� ����*p��zOR�W0ߍ���^�sD��D�%0]�����a����ԛ�-S�t;������){�vu��1,�N9�G���}�������kT�	6�S�����{@��Ljn٭���m���Gl�YCΥ`�v}��ts%�9���r�&b4+P7Q n�8Jձ���=�46��<6�߻�ҽ����ȫ3wm�$�y��iѰM�O��1�9��,z[�#�؛����3���:|��#��kV*�vҀ���՜2�@(���#78i�� �����Q�7�6���"�`X|���i��@/V����~��k�@�aD��
�:�WM�>N� �Z�GZO�a /a�x��L�����f}�R)��[k�l�*2	H�Ln�z.���?8p��$&��Yi&Q�⅗N�b�7#���lDr��<If1�2���J��h�-��d��]ۑ�%��lW�ʲ�/���`_6�`�FN��L������&�$���w�_-el��3�fi@6��E!K.��b��&=���V���Vy7xj��DzkD�nV�۱����ĉ˒n�;����o�E���=?�n��w�Υ��X.��ڍ�|:��:b-�Q'D�:�ZI� `�x�\���־��k|;7��f(���D�>xc@hg�b�n�ݦ�C�	��,�ڙ���T���}fP8*]�π�{�:��Y=�Ў%N]�'��Z	�N�O�AZ�θ`,��8"-�
q͜0k�XN�}�ȍ�0�{��z��o9x�R��)� z�r �n�!<1��S����~;@��ɚe�w��&��ʸ���V�߆�ϠXR4��Ia�b�5�9F|������ '�
����92�r�ػ&��|��d��¢Q�hs�D
�a����plmE@/F/�r��~P��� �CS{�������F�y8W���yߠ����G�׶����H��F����1~qҤ\�bϲH��}��v��q1-�Yyx����ٓ��a�-e��!N;�!U�����9N�p�T��+�;�59���l���I��T�$L��k��8+G�Ϋ��}UB���Jz�:z�������z�b{��]L��kӒ���u�sY�4�X�����LQ2̺�?�H���<�tb�96Ͻ3[��
�{�����~���12b�'	��:���#�6`-3A��(�3��?���*�F�T�K��B=pe��k���%���k�@�i�|b}�p�%�N�W�J>lMJo2<Au��?��F?�7v������)<*�@�\w�Ya�����&��:��|��!G×�:�'�~���|���qP�T�k���^=�í"������WN"�J�VJ�~G�m蘨�]j�o.���-��Sq0�BܠXmC�%��蕗Kd�MC?������Z��Պ[T���T�Ÿ�i>1�yS$�/i�1��}q�5��
�-Q'�{�����*��e ��a(hė �2�67��3K�j��of>\�l�#�u+ F���"������/�4��|�t�~�ܝ�.mP~#1?�Re8���0bͻ�Xe��/�&gC��|�Tu��'|Y	��S[W���&4��d���=�$�����D'w+��P���0޽��Kq�L�Vu��B����E��W6�&�*zIv~���9x�p�hV�<���|�����:���ʝ�WH|n!C9�C;���`}��0�`~A��y"o�oӾ����"���&��Q�Y��t�`.�n�� A7�=:wNr=E�.��'��>�ao����V�G�eJz�Q��!~��tċ���=��?�ڂ��p����ǹ�������1Gp��RG��H���h�U�AW/	�pg�ІP�4�U
���o|Έ�P��Ɲ�>�`>����e�\��?2����Ȳ�1�Ѯ��Q����f�x�>'9!�v>?h��?v������'�#G�$��B��f�:���j!��Q��,e���@ޞ��̘JÁ|7 ��!s��:�\pq��(����AY�������IZ�#�Mȥ�Z����������(A�ґ��s�8`����!�[8ϼ� �<�Y9��s����p��[ƕC+vp��4�J��L��d	�hG�g�!�5�z�X'���Su��s �m�=�}��0G/�2��W�������#��H���������N�Bu��PA�`GV�?E�jfў�`R��,��nU���{UmGOk�Ү�%$�4�����u��,c�ఞ��[�Z�7
����zx�0/IK�����+{�b9���x���K4�M�ꭻJHX�~v����> x�s�-x�ݛ+?�u����Xd��+1^�[s���*�ś��R����TDQ�l�5����0a@)�Fv&s��M� ����� �n}O�ӄ�P�|!ɝ�������������ѵ���E���K������^�A�9zfS��b�ڸl���C(_6O�.���� ����e�	a�A)�'��m�%�"�G�R��	r�u�,��9!HF
7�����ܩ�G9���߻���'���r�3�4Q�<!*H�G{;�٦��{W���Ο�����6ڽ2�Xpu�-�F2a���ʙ��B�y-�������2M$+�0�E��QL�=�Ȩ�I���z�.? �5c�W?+~����)bK�3�n��ڃM��m��E3fD�@��~��?� �oXe�G_�y�w�N �aD��U� ��T��}:�Rb�Pc�O|~�����d�@:E��I��=j
a�^�m�oY����/���K��ш�Ui���+��:���A��Y��F֗G��`G�0,�
�y7�P}�q�t��_�Gd�mM��z	R��]�ܐ��ߪu��>[�m�x�Z&��]�������j��/��+ßϏ�g�B�Ӎ������?�g;�j��O�Ƿ�4Х7��4խ� ��٭����P����G�)��4�yI�YN�=� |M��0�eB�P�����,4��v6��u(v83!�Z�|@���BA�2�+B�㿬_}����R��<�����~ۛ�X�1=���ϵ�S�O=Q�"�}�o�������6�Jx�]����I"��vS�پ�FT��[^�漖�)��Vhj�p���:!$M�ؼ��"h�@��� ��s��)�������|�`�
p��z��j��aI-��;�9�g���8���zY��Z_Qmѵ?|0��9�)�W�i�HV��aQ����S|B����PlWZ6�~��κ��eh\0��o<AGN�m��~Qĥ��c��tt~�5XU'\]��O�����@	1���۫.�b����M�_�K���$6/y�u�w�*�fj;�A���D���$ge\���bU46|2���#��zҌ�0Z`� =?~<���c�3�����:�i7�{%��V|�!�b@ LMVڿ �ٹ���7�+��/HJ�Y�D�LP�2�p+�c�n���;xL�>
4߭9-f��뭤�T)+ё�P!��L�ο�>�l=T�m'�����_�ձ
�c�����JEj�o��xX�!�7�0�d�O�{��F\C��Q�,��i��ퟜu�����mj�1�E3�x�����?���YQ\w@*E�}6�{�Z�>u������U��BR��0� [���`��T�3�j�A���WCdm�z�����nJ���A����S��0A��j}���v����/�0H�9�@��FU�L��IU�9��Px% �n�O��ɪ=��'}
�#�dj_`�[F��ؠ-&0�¯awT,��*�}�����O���Fj���<zK��f��Z����/;�����o&��k�ѧ^v�	�l� ��A`ڱ
w�}N{ϣ�[��l���V��p �U]�е�ކM(�2NH���>rH6�	����01�˾��l�������3�=�/ާ]+�k*��#�+�DJ
�b�2 ��_[�µ������9�kbJ��rm��Jy<LA�O�<��*H";����1_�E�^`e7�d��I[���n5gɭ�� E+�*�NZ�Rg�ѷ��ɶ��tDZ�9��s�l�e��ž�ٞ�����z���:�g��t� ֑�R�X<�i,��»���4b�R�?ϻ�'I����!��,�c�*�J$:+n��(���Ia\?��m+��9��>���D�7jyǓ6��D�%�b Y��������u�g'�o��7t�c����2-F=Ҏ�;y*��N<�l#��\�P���?|'���"cIw�v�6S=Lbg�L�*��úvEj��ׄ���_Ԉv��y���Y�S@	�36$0���h�X�;��R�i��b���[b�F�����k�*^n����W q���kb�%����:��C%��E�K~Z�
��� D(x�+�M��B������Um8�e�������Х�QOm%�w�b�������N2),{�=0�L����o�P�'�U���<F>B�[Hꆓv��ۥ���+�'87��f9H[�B��l�ǹ_Ry�vJ8Uz&qT��̚=���ȭ&�.T"0��ً����=#)�����>�%œ召 ��D |�}��9V����jV}�|W�om��΁�u�F ��"'�۬���񹮺Xv���R_��i|0vH�w�}�A������E�{�r=��4�d�B��m�\�2G�fk9a���Z��#��t��=�I%�*�B�-�q��	����Ծvh|�����[Y\:X`̣�{+I�&���X"or�%`��g
G�֧}FrM���L���H>$Ex
о�N��^>��M�5b�_�G��p���h�{���N\aX��Inqr�����]���XJe��Cw޶!�`!��j�R��o���˿���R���ȁ� w7�^&�*�M�v���F�-�\ͻiϤd��TsN��R���7�`�k'abdU.?�]��y�3�l�+������$[ޯ8o�-é�D L~D/H�-�d�DyE,�f�"Zp��[`��`n�g"X0�^�Z�W���\s��޵m[���Q'���T�a�ȟ�O1vpx�>wGi��I6Zb+��绗�����,s F��Sƚ֚n(�� X(|2ܮW�3@��d���?PLn���RkRFs(�@1��3���F^��;����/Ҟ��9��)� ;�>uV<3�&y����2<	��Ϯg�����[E��^9c1�f JN�������y�(�x���Z)�v�'�����\��-���	�������ೀ!��� �v�\�䳖r�p�hK�Ռ0s@�h�Z��$S�{�x[n���V
P�>��*�l��o	>8�j�Ё���4}.���JO��