��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V):��5�P���!�gP9o�;�@N�4.�Hcʜ�qb��V�W�@2Y9L+�HѴ:/��f�(9�$uvv��`�G8��_hs��t�5�J���=�W׋4o�0Źh�\�\��R���B~vC�B�b��.��f����U2*Ë�r��z��T_��zY�m�� �8��t����:�ڍp+����MHI�:m�Ne t�<ʒUP;��x���Bs���=�x��]�@�awU�'��v;�"��G� ��j㍤T9'ώ ]�5���>"[�\T��JӍ�(�:X���h�����,A'\-^�&bx�
�\�A��_/m�P�����-�k���G��׭�9U�dX���h@G<4��lȆD<�� ��v��H["�UD��Z�Ldq0�ڀ�R���w��łF�pO��6ԡ#6�1�Đa�����u�	�^0:�EL�'������ ���Z��se4Wy��
\e�8�=.�P4|���T�@1�VU�h9��?��(ߦ���y jm&̣����Wv�����4,�_J�Ba���t�-Nn��m���H햕e���`3V��e�,L��n#��pSȝ��MH���6:�ʶl�&]��
$���U��d�eAA�L ��	�^T>��{�hĝk ��K�n����E
6��<��h0w�<I4`$k�j{HI侥��X`�q��H
�0ہ��y�@.�a�?�]'C%M˖*6'3-�wU`��,=��mm��@�!�UK��c�=)�)�� ]e�>�&O߾�T������H+�Xw�l��6���5U&K}ǬX�л��,����kp�}�G��t����'(�/�Rr���*�����T������G���`H�q�Qu�������*�hd�cT,�9k*gDi~|ݒ�X��YC��}��2����C�`~�|a��)��dJ0|O����p���b"�q�X�!��WIt�_�s_ �������H�,�5�v�`i~X93���k� ����hū�H�'^�9����IP�rp2<��q� 2�U�|?�F�1m,�S?	�\�~�Y��="\!UV~S�(g58]n=�uvfᷛ��8
M���r��g~D��\�aה}������z͊�ե�*�a�7��~&!U	�~_ �\rDEh��d\b�~軎���1ф��sqC{={����rw�2��r"���3\&$D7�E�P�J�6_�h'�N�;�:X�R�]��mᏒ�xi��v<��G6�p�����% ���CU�x6)�bOҌm��<�Y�2�{ ��5�!E~���|,��;/U�qzmzM7bğ��nM���*
 �{��	m9,J.�"]˴ɃǑǲo�NI�ںU�ct:Ԡ;�*������WM��G���'W�#�R�_`ޢ������X�&z�gj�ؕ�=���:�^�y�	�v�;\�je��L�bh�z�g��V�AU��*�!եK��cd��#Lm�q��v�����bJa�N)�Xt%XL00�>��_�TIvtp�>�=VcCs�,��G+̲S<�+s���|����`-����⨱eQqȇ�?\􂐶������;y�{br�T�K^�4��'�M�p��oY*�x]��@RpK�*͌����_���Tm+��jE�f�m&��U_�9���k��Zq��]t�V|Q?+_W]䤤H8���� }�ݴ�5��?x�a1��I���m�k�s�]����b���siqKϠӻ��bF�j�EqL�Ț��}?����+�iȁ����f�l�)O*VY�Z�_�R�=nq@��< �!�H@���ln)c�Z�k��zl�ns\�<s����x^��܏�E��)i�>m�����UI4Mٸ��Y	b��^�~��U��B��T����@�\obA�9�|�\�[&�`��ٲ��i�m�9��r3���⤿�r\�D���0K��f��)걤�M28��D�7���ˏ��C�ˬd���Ĵ$B�Ӭ���c��L���Ao�K��Ą�����NgaPǏkҿ�b�t�z��ΝO&v��"��А;.Zn~��a��Hs��K��J���dbn�6t4
f�	�~�-�A�[�5� ���i�CP/#����x�o,�!̻q��QxD��W�5|2��Zx��/���k�\/�{«1ņvU�0D�>�ḐEC���Dk�U:�JVІ4c�\.d�_^�H
��ΖSW|��mG�ǫT!G�oD�w,���.C���Q*���s�~zh>Lv6@\�����e�����N�r=�)�I�V��.Oଵ#ǻ���q���qm�:�+���K�i,&��	�W�>���w�S��(����d+i��f:�OZRY�k������&Ԁ�Q
��Ɉ������ʐ(�E�0��!��r�@Y}��i�)qg}�$/,%~�R�:�����K��z�/���rq�(͂��|J�v��r�����ft#3ee��l����T]"kj�[c�%��R>;��(!��^t8��
#�D�Z����p�d�!A�j~�ā��O�$=�N��<M����7�Z�0�/���1|S�wI�Z)V�<�7|�1ӌ�0n-�4-��,R�����Z�	(����Y��
P�lv=�K����|dm���l/+����`7��R!��C��tab ��ĝC��}_5v����Y֡�{<K���A؉�w餢މ�ǥn���d��&S1��kh��ү�r@T�0_��P���wR)�}E6��8�8N�;l�w�|���a�d�i���*_:���<�fd��O�Q��q�	%Q���mq��8�T�OQ��i��-G��[����y;h�dE�u��Z	"D3ŕt�SP��y�5�D�L�˺+�Lw���-Oy��� ;�a$�,�O�9ЮY�=e:�����v��7���!MVZl��?8�Q]����Q�<i�Ls�C��Ṇ���&#\�ʎ��e��J����F�������|����PS�0�M�ľ�,��j��i+�WsSI���	�<.�'�kL�DTq���&i)bu�ϫHÊj�	
O^T�HPW7���\�7c!+]]�02����R�jY4 �jo$Wޮ�S_�/��y�X�K<	���-A<=�3��]��9D(�}x<��q�^a��?�[70�X�Ws�ޞG��5X���}�^����o�R�)�HηAe:%�&�g�!,;�w@�`��ݬQ���}d��M�$�������k��ld([�Y�I����B4H�Қ��7�`�-F������C�O�C)}��J�f[/6^G�kG�Y��B�J5�`)��l�ۿ] ��w��i�<&���h�W��8]N_s�+ D�"V\`R�o��թT��z���X�j3&���C�c��;|��[�;������	8(<����lc:!9(O��L+P�L��Ҵ�YۇV��ء�h,�!�H�1�%b=��MԄ�#�ڡFA���{���o�mE�6�2dT��#�:���i,q7a��NC��A�v�-M�/40x��d.|��T+B	�j����d��ݺ$��Ƅ7I�$!���{��������Xc�
S�c���#?���"�6�C=�C��=�8� %%
�6_EV��s,���I�<������*#o�cv�B�4O%{q��=3ʝt���?�ֈAOB��Y�����M@����!+R���Ɗ���;'��\��=�j5A�#I���ՈxeV|\ܱh�$���d �O���j0ϦO��P7�W�s�i�n��$�KU+2�����&��W_����VrsS�����_�*���E�)�PtIVbM�-3~@�xj��{/y��!������ ��+YT��-�ޑPY�jZ��G_�� �����F�\���`�p�$K����;����5%����1�D���=+�2�|Ƅ6�Gsr��Cj5H+*x�lY�ӡ;�B�z�	�VA�0�_6�b���ąd��;��Q�]� ��ih������]
�#�QP�N�I��@�Z�vҋ����S��*����_XL/��:w�