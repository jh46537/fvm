��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&-\X�ǅ�?�;�V�00<���w�̢���8�~s�2�tb��e����d��2?p�ȹV a���"T2���)^�rH����!T�R�(.�/�sg޾۩��FK�i�B���R�р�ee���������o�c����y����z�C��]��F�a3����|D�Q!�M-ꖒ�3�!�olM�1s
�foI��ԀH�Sgohf�%�r�2=B2D9��W��x�`�"��[|`8�_�ӽM;�O��	���]������ԏ��.5s���)��T�P�v�<2ǢΉ$��$�]��#�1Iйiͽ\pZI1I��FM�=�q�-�	�@D�%�u�a�	�nؓLjM�h@����F�Lz��\�1����� ���1��m���Ev�R����B����*�㊈G���I���쬢<2ś���o��a�b�`-�ڙ ��1��q|�-X�ݳrz��T���B��^	��Ø7��3}��.���&O���rv@�N��)Ԁ�^�Vԣ{ZW��@��+۔BD� �MVoH�SL��ay�-S�~��z��TԀ�)5{M��h��(����ռ����u�F��؋e�w\܊�9N\,.��Q7�7�q	N�VR��O��Q��u��FB�Œ�L?,�U1��bi\��K����6��W���pL?��V�Lw���ҩ�d^�@
2A!�U,�ה���g/'�z`�2ͅͲ�׿�n7�(�V$�eQ��0����c�:d��"UE���EA� �k����E�hzY�nP����7_�d�J�(�̨Ҽ�K}��8g'}��,O2m��s����U�2��Ϋ�+a#��.�i��Ts=�ȱ��n�{o�\,Q�o_nZ�c\��Y�>�
�ǛANx��+�$��:��f����W�5�����ؓ?�P|s�h���?�p���@�Id�>oWSW��Hst�*�i\�n�O�\3za:~v��D/��6<��R����T8��$~�P �e�M��H~5��Pczǩ0��ܤM���ׅ�:�)t�c�Gw���ϓP�%��M�e4��v�l�n.4#q�Eu"��g����+P4W�/d�zf1}�3��έ���do��;�G[�FP[
�fh����ظ����|ᢶ�!ٛ��u��%��ݚ���F�%0�?W��)��O,�f�n=f���Gߖ�o�e�~�v�BI���G��K�#	�ԉM�����a{5W6s�l��$��Y#�f]�	�h�⬬����m������|P�u^�Z�P)a�dTZ20a�o����8�4��b�`��O}y���k,Ӌ�:��&�g+ko,�]��Bebr��RR���R8�e 3��)�K�r��I�t*�~�@5��!��;��N�*�Ų�(ZO7O�|�,��'N������p�K���Ot�fS����l(o�ǷEe�0V������;�c+��c.CߤO�T��ְ2�z^{��uNɭ�jZ�7g��f<�%�3w��@�_���?�ۥa��1aJ��J`:�tLK��/���cSo+����ݸݬ���Z�K~կ�n�H��73��bE��L&��n`���G��n�O�r[,.K�.iv,�h��>pr%���!����e�J�K)iꕡz�aB��,@�vⰋ�`�j�i���X��t��Ā$d&�#7x��UX6�ʷAKU��wwHm��Ǿ�W��"�ҏ�٭`f�r�a�o)>�೰
��#��gY��2����/NA�L.�5i�܄�N���f�$���)�X����$���|�����჻�-|��Ԗ�NΡ�h��WV��M�v�����XѨ�8t ����6�\��X���:����v�����5����7Zӭ0��&26{	f�����$c��C�l��X�n��z>0��,B^���f212��u1M2�"c���\b�����2�Wp�t/���J�qEʘ�\����ʏP���<f��(��M�ΩR�ZU%����{8I�?xS�&Y�T��l!���\�Zm�p�@I0�}K�:��#i��M��Ai�y7��;�s�v�8�m^���{cW��ov���k2�	�f��2�kx=v�9�t�Xͽ��5����V4	�'�Y���zM��7���4W�*Y,Q�Ⱥ��\�
r�pY����xT��V	��b&��#ɥ)����|Іd���`�_bh�)�n�w��.�ã����N��2���1���EXCm�Ye��;����?.�eS��.u3{c���ضI�ʅp�(�Hd�n�d�<پ��!�Op�[�3R�� {�mM��������_�$Ȋ�u�l�?��OuC��zA�i2���O�����xn˖I�Z�Dʛ���MZᠪ�0�pأ��P���>Q���).�g�N��Jw�ǎ���j���1vE֣D|X�N���M��R�\����jضP��G��?D(�[�yڶ���L�#C����(JVī@���!`�%M/�>ؐ��g�H�B\i��� I ƑQ��.��u�2�	k�Q�Xm=�9��#ȱ� g6f'���>����3�,`�@����7&u.�����Q�$�s�*sg��s���l����֧���}8j�
�p�%��\����L� �t���Cu��3N97"1���Gp��ȥ�N���PBG_l_�PP��E5��<�Y˗8=׶ �6?;�!���Ț$cMk�$:B$8_����?$�I[\0b:u�m��Dݼa�̔�s�'���Q�t�4YN��y��h���@��X�9oJ6�ڴ�de�%)�֫������F :������%��OQ��JQӀy�`�P
�M �����+�5�c�wS@w���ǋ�qd��N753���n[���Lh����5 �����I���a�����7��_3~���8�K8k��~A��4Q޶w2@�N���Zŋu�qV{�:�gמ1y�6f��M��'�I�{��i�"N��@T��=�zW�j1�z�g�L�ו��]F���,� ���y���Y�?��m}���PK�b����jr*��ȵ�`������~���T⁭8�@竂�q��a���튩��M�hY��b�C(�k�!�ᢕ�9&�Lw����H�`�����r&�ѹ��?E��rup|o�;mʬP�d��K~]�&4�9�?ް� '�}(�ޑGx��Q\�vzxCX�Hh	 5=ZP�P,D�`�m�9�'Ĝ��ߎ0(>����'�eZL�sz��^�>B��3f�f��20܇�����`Gu�u�ʺ�\�
Z�F�va�}7��0MĪ�B|Tl( �_;_�"��v�� I �Z@�sp�W�&܎x;�`ȫ�Bgd�h5#�1A��9y;
C�$&k<Oҫg-q�t������韴�1���~ׇ5��x�mxh����At�XH������eu��q�Ş1��Ԙ���@VW����x�|A0��n%�?n�����u�ľ*��_v4��q�ْ'�d6�'����*���-�T�ף�Q �N$��R�|Bh1��H8�|"M�2��"˱Ĥ��Uŧ���fW�'��tM���(�6���dv���� ��R��6�#�V�8���!P�Q��r4���z��xY���ʑQ�
��q��B�J[��QW���Ae���/_՛��ڐ�W;�����>CD��J�H�`Y3�(��BQ�A�!'�&9.��-�2�E�;\��'=>���?2�����]`B�6�W��{aa
��a�f`�Ɨ���;��P-�d ��P��\=�4�nc��*|��͑
�2���Z��70�������La7�e�X�m��p�?QT�?7�8O�'�	��I���}Wch���R)�J��zJ��� oB��iU�1�b�X�G�����7	l�/��]������m,���R�������Z҃Y)V��\z��IR�������V���) (E=P�"f�;�Q��Kąj+�W�D��O����/u:t/������	E�;,�t����U��m�J��@R����Q�;��]B93����*����n�~L�X^�#��qV���J*a��ÍFn�4^��5�M��O٧��"���+���-�˥1�W~�x�O[&��\6����z��R����D=�P��	H
�ß�7@�20��f��w.F�w�L��aX�T\�ڍH)	(��&�r8q	�B�����R#S�F�Җ����o�5���|���s�˖qҁ�7�WS�Xc`���X��q�¨۳W��m����s��t�~bty�j �G,[�����Ʌ��ɨwǶ�ϋϽ�Ez?�] ������7��#3`��O.bq��������#ܑˑ3��n������:���ٞ���4�]���jE������D�o��H�5jdy� ���X��/���؊ی�o���#��_��\L&ҡ��(�ۮ���g(t�5�f�a&�V�r�C5:�Q�l��Wa�ۢ��+�>���b�-Xe��>kJw�ը�N#���S�q���26TP�xC݇�gX���}o��?|.]R��H9,�\�U���$#�#��=At� ��۸/[���ƃ�4�{��/~�w�Z��7s�"�#����1�\�#�T� �{��Ip�٤�}�C
�%]��e�����: ������v��$Ԍ��Qa4tj�]ܒo�5��;}��c��\����V-Gv��ԇ����oHK!u��� u�9�2m���h�N�Ys!���.D�Q�v��@�����E�.S�Ai�D��Bnbb~�t%#�4�(λ]4Hz�F���aH1��0$�hL@�Ք&����z�c)c
��9��U��X!x�!�$F��#�;)�[C���C�8��n��bv�0�b蔗^�~h������k��>PWT�H���. �I99�y���ǉ`��V8�W?'-��1vpX� *LK�����M)��� ��	H#���g8��=3�.c]eם`���& B1(�%+:��r�K]0H�LX+<�� Z�+-v������Z��a�6�"Q6j���:4j��OC����L�C����ʱ������#�9P���JZԹ H�̖����?��(�'�K�B�A�����o���Cl�o�rx"�	H���܋p��Ʒ�Y�_�N�����2�
��k���>+2�	�ǅ��5b��Ml�zS���6�����D�Lhf�b�&ʤ�R(�B$���BE���0��ih)�L��?�p[�*�U, �a*q��P�E�z��l��caUD��F:B��?���o�w/ �n�:�UO'K���]�c!�B[J�}�4Ŧ�|����.�}x��*��#C�����}�#��������?S/��O*���9M�&kLHFb�)A
��~���Oj�g��{�6Z1d��ɠv�T�#�N�ߠ�	�jh�F4��,�tt�G���m��1P �F��l���ۓ��������G3QX&�TaAc �%�(jn��\z�G��E����)4�ϣj��2,MJ�?b['�k�f}���,�v�u8��u���@n=�Y�Gt�㚒b��|9�w�7�QAQ�z�*��vĲ�jB��&��I���:��2�A�
+`�te<�\ʳ�X.:
Y���.���� ��}Wr���e� �|�N�W��!�F��f�`�MU�TOt�G������[�*��Hno8�F��+��9�NGK��G*��B���:j��:��?Ưn�ϐ<3A:ˤ��\����~�؜�i�ib���z�	�GR�(V��{�g�|k��3"k������:
ˢ��s�z�'1���L����eс����� 1ދ<�������럳��^�.*+�9�R-9@D�7X�	v��������u�E(�C�J?�J��kROl�qt�J)��@C��2O�ؗ������Cc[�/J��J�6��pѸ��|����n���J��,jFѧ�ȳ��d ��,�<9���n�:;��y⁯�z��cvs��)ð���֍�H/�wH [�A`�>��u�Vh�:���h~>`RF4�b�?�G�F�F���p����HD�&��,�Vڅt�J��\���[R�c�"�~f�W�t$E�Z���7��%�gz��3�>���`�τ�g�G x�3��� ���' .;� 5���X����38p؇8�A�K��ȏ�M�S��T�//�7�� �Q=��j[$��g?�kY:g�2��"1P�c�%˾*�@o�d#�bi]��;ImCN$�o�j��=z��;�	�P�:[�/��F�FREһ��� 3T�xQ��B��������'n�K�	{
e��X��ޅt\�<Ŀ�!��n����XgDep��{��F&['_�+��D�m����n.��h�.>]{���x"v�[��竤8):�B��43as���:v�V���i�j��C�,b��z�!8j�{�q1��2K_�VN���Վ�~8~���n�RN��Gd������K����x?�7)RZ4f-�Y�=��{$�Z{�~���A �a����O����r[�"��y�ov$�C�%+c!��*���꾆����`�p0Ͼ���w�b�kk-�[8�nm�]ǜ^�$J _��&,��\�X�+-r@p�t��9���+���<�󨺵�2m�f�U0��rC�$�ա�M`�.��*y�>�L;6����P�L������P�Uk�Νbs :0�+_���߶"� ��A���	FB�qvǃ���:$o�i�G�6��E̐~��ZBA�#ջU@�V��`����;I~���f��m)�=�ޘ�mvB��X �o�u��643�	i�ƊO
���/�-����:!AH^��K�_�w�巁o�>"#�m��fp�yQi�F���i�k� 8�k��_�i]@�x�bO������hL���9�$E������-����4�;�2/i�RX�(s[�'��\���q���R~>�?G��f?���Le����<��#��f���@���"���U۵/���5VI�D���w�Q�?<.��k	~�>Kf�b)�,��;�lX��k��pU��X�,��K��%���3��Ɵ2*��-}�Re�9o+?>jDzp)�9R�&�亞�E]!��I��8@�S��S�.S�͸K�Y�B�݄���3�������MW����II�T�Uhp$6(M�{{�XR�`1��p���.��\t����� ��f��
؝�k�)qaG^��x%e1��[_��r����5���A��~G���,/$4ܨ����sǵ*%*�f���[Ԧ�Ř(ĿSj��DS�q�J�,`x���>T`8�G��>�Cl,>�/�c�
��P E���d��1e���z��xݕj��3�B�/{�53�%� �4��jxh�q����3v��J���ҩ�0��$�ąuio����0Z�����J|_�
� 8�::n�w酦�/�9Y2��R˨E�W�=P��5<����rF��S�v�s
�志��O�=Aҟ��Tp��s��2yXk-��1��_���j���*�r��{[����v� :�;J��;�O�������D}�}q��Fn-���I-5���(�~���;�{,�0������d=?LGp��,`���۳�;�$C�Z�ϸqh�M&�5�K�x��O��?�0�\��Y�<.DDg�g�d�%�	+,�������7�G�3�>@��v�����3�����h���,���kߝ�wLg�t���):N��
�r�J�0���
�m���"��]?:8�;�����!q\�E���١]�c��m���}�$�4L�OK�����'o������g��A�茳Gп��a1�~8i�>N�EP�GE����K����ωI��ѹ��  �k����� ig�mT7��s��Q�9��3�lC����3�o��a��0;�#��1
S'aYя��K�gDi���]���Gó�'�w���q80ٚQ} wJL�'iT)m��C󧣎��u4��E^x�87΀m��k@g�B6,m�h6¤E%J�נ�r�ƀU�:(��,&޾����T�>s�=���w�M�b���W�ŴI���^6~p���(	�N�
VЖ�������Ѡs�]��$��1���!��l(���ba��_ua��dR����kL��=޷��h�&���ze�S���ђ�	���nB��`G?{
U2�s��7������	D�@04G��ѵ����nM8�M��&Z��R�A��Z�p�F��@��#�J�_5٠__#��VK�����%�H�����	��NOg��O��W�ؚ�;H�^,�v�44fK�9ϖV��0F��*�"g]~�Ov=ֶk;��c�Upv�]8zx��:�eO֌:)!�EX�Pb!�2g�F;_E"�d�0ĳ&F�+��D�f�~	:�V���G�I���֯��1!ZcK�ҭ|<ȣۂ1�0Ƕ�|D�\ �&"p�����6э��;+l��E���2��V#$D�&��fQ�<�����4H�*t��)�g͡��Jx�N��d���_f>|�G��s|8�E�X�!���d����;�)ݖ)S���
��Y�����L+~�e#�>�&�;vH2K9����^�V�t�^|_����p��"r�WYmq�m$ �vJ�y�IՊ�'yT��\|-.���idN��Wߩ�@]&�.��PfM/��`$�0�hBy��ŭ���p�9ӼY���w�2&��)�bo6-}��Kgm.8��q��w���� ��z�fE4Y'��BD}V!��as43th��P�ot� 0b�%�V7����ᲘRt_�!��!�O�4�ƜI��D���t�vs�ǿ6�y�`�L�I��A���L+P˲6�l��s&	���c��0+���?�#�����el�G�#�<h*4�[��V&Q��(�����
��t�UT��>G��s9�*xRR`y�U�Bc\��2�d�͍�Ռ��b[b����z��	K���7{G"ʨ��*k�C����7~�J잜&^��u�|ws�l��V�Y�l�k|5紼3��&��?S�L���z()\n~�a)k����3�l��I�����]��#�'� ���6:�}Z��3���A*�m[��S�n�:N=MRG� dc��<�]�l��� h����i����~a��T�����3����� ��ќb] �&�r�^O�R�8���w$�62ģ+�H{0��u��z9�{'�}�p�G��I�)�y��⓾��m�������j��c�<;H"��\�f�����934�ۭ�dfi�����<S�R5h��:4��\��o���w� ��Y�3�=/�k��=Yxˁ���C��?s�qaR��e:p�zT������|��S%�F��d���H�qޢ���%UQ�zz�S�w�ڻ*{���S`Ef�%z�B��"��$O��ݬ'6�Tr�b��P���|tD]���Wg��27)��G,ߕ3��ES;f��3�{�ތ�4M�C �s��
q/�����R%�E�y��c�����6|qw�A���%&�[�������,�͋�ۑ����ID	�eD�67�>�d=/�� �؀/	��\,u� ;*��<5QK|����VХ��,���$����^B��h(��|Ņ苒���Uo���Tbcϝw4�Vt����zxC�h�����������ޜ�q�_�/)^�c�ʿ>-
7������L�|�er{�(^i���(>��ŭ���d�D=�7F�����7��O�Ev�Qb3�Fr���W_�X/?�?2��J�ww	uY'����N�4z��W����+��G�����HӠ9{>˵|�aKTYp��E�ђ��q�:�x���1�gK�4n?�\�3H��
���G嵩 !�W���u�iiy�A}�u��ۋ2U�5f��*�d�xv��� ������!�5�]md��{r�Yϲs�Vb��q�
�i��>֚�-+?���:Y;?��1_������� w�c�
�0�8�O��5��0�x�8f�[�]UX[���^��)�\��?߻����aR�Tu*t>F U�Ӂ�dw,c`%�jz"�{i��W��~i(OB��(�_ xT�[*`��H�7��m���5�y�@��a0쁼������Nl�d]v8b=��7ޓӑ1�v�幥�e I�ـ�+@�D�a��ѿ�i�u��:�%��DEqlS+}+�b�:L��,�.&(�Y� �8�&{Rr�+$�m�Pp�C؂�:��h�=Wg�"D]�`�4Ϟ`il赘��qu����1[C���{�CІG1�ǉ�{��+�i{C��"���rb�j�LςE�?ϳW�Zy�L�;�H���s2XB,��F���V��t��p�U�I�S�	l�㧨Hu����L]2O�đ��>�T���������9�р��L6Ȱ��ˢ1��:�(G��z'U��U9c�ly^��5���'7n������;xs�cmO`�f#_�r�}Ğ)U�OH����	qu����~�v��r��~6+�}�>v)+�f c��%(�,�V ��W'����P�	���a�ͨ����I�l��P+M%KB��=�	����Qb�t���j8��+,s��4�_��)�D#��klD���g!��U��+E���(E�?�q�� _�$	s��̞�(J��vj����r'�AN��@�O.u)���F�����pgC���`zIqn���_yi� ��RduA��b)�S#����g�h<�K��Qp�w��+'��1��gx��:<���Rh5�,ڶ�Zq^<�Q O�HP�#�~t����)cr��7 �`D5&��4���D9��*[�pq�V��b�d7�}p�� %%��=�/�⌔�U��h��;���^7qr,�bp��kz"���Mq�H��L�4?�qg	����j�H�w��C�v'YT�4�Β�(Ǎ���!q�=�{g�;��@x�=%��ʔx>^[�"�R��>���(%���c賶�$��G5`u�`��t[�٘���`�ىe��a����($���� E�om��7��ʞm��8~��XT�v�L��+�
��X� +���y�����G�$~�94Wv�L/EY8A�B8i���T��&���)�׷�z
���TD����9 �f�μ�9ܷ�-)�bد����2�29�)6:�^������͑BN��2V�k����.�).���ɹ�s��X�3yA���%֚ڂ�����������M4ˁ ���#$n<���~x�U�Sy�J�	#��pKnݶ�N0��R���;֡kf㒉s�ć`Eh�"k,{|�&�n����ψ*	�b�3�jS��E��yuh������j����Z���@�(��]査��R.%�ѫ�7�L�}�_ӈa>ـ�C�k�j|�+��"Esl��sY�4C�h[!;��Е�v�*�E9�Gf�U˛2�BFW��ڲyv��@U�󔑜�W�x߅�Y�j�&%~
��BB��o�M���^qg]M�����me�?y�!��zoGi:�o��{	�z�~zFJ��z����cW@�����]�g!㏋��9r5�8� Np����Tc0��j�{���Ut���1���A}���ޱ�.�XjY����b����U��M���w^�8�����Q&e�{����F��/��κ��	�6�c��^|��x��ʝ��w}�$��X��4�㪡w5y1�&�]�ê�g6��QS�db֋[���Z��s�Q��b���.B����b�E��1}�	i�D������膝L�H�V��v����-¾k	��ϣ&�+F�`�<b�G��nV˅N�}�<�����'�N�E1Gq�D�T?�6�߯�yW?u@��������՗��l;Ɓ�<-�G��"�gh�YCF�JRK�j��7F�)I��>Լ:y�CQٴ�%6�[�#.��T�D{��rk��r�$�%�a"��Qi�72�S� �ĔA�6�C���G3�|����\s@Na�6�Z��FJ�c��AE�%�}N�=�K�6��~@@BK�-"��p�
�r֬1��E8�[|'���
��Ԭ�O��b�.P�C}q��ƭJ1kn�"rƵ��ޫƁB���-���(j�6�]����*8�ɛ��f��.��E�=8��9U�{�CA@U��P����_�Ř�+<�*���骷����
5J&���������\;^�Lt�TM��5�:�rK�8qK��P|!��vIzM�U9�g�����*��3,���S���6�bh��=�y�|Ԯ/�z_�����w��!*�ͅ�32XY=�䣹�Z���n�.d�w�=O�`õ���`R�Pd�7��_�SXޤX�<zg����֙��y�i�U>Q�A�-lҖ`��n�\}H�i(��vm��?�u�*�wpk�6���}�#�9]p�8K$�c��.D�����O�K/�'�}k�ł�O{� n�%O�g7��¬B�@�<GO),�Rd�N��шӳͥ)�P�My(��K��laj��`X�ʽS8�v>��4t�� ������ڰ�c��2�ǝm�"{���Kg�#Vk��Ló*ׁ��b�;xa5�7��3vns���y?�2�����s�ڇ�l⮅����/ꅪ��Q�z6�2'qPsն<�p޹����~��uZtB�u�ZVK�m�[䮱~�s��������Cb��( �$	���գU��#(�Cĩ�Jo����:��t�ERZ��`e���[�$��d����DWVN1L��9��3*����w���-��/��n�W��5��?R��c���~_�|�+��c�
@x(@Łzg ǆ�b��M�b@ٱ9������E����=�/�ר�8���1��(��E��rj�VuV�JU�t�,tCb��]�dtA"�F��c���w�@��"s��	�P��fV)5�(t��֓}�KѸ���K����;�.��KsA!����+���oa��;#o�S�tZ����	�{�K�����e�Ve�g?����������}R\5���m�#�������K/-�����"o ^�V���O����o6\�h�}�z�y�����Iџ�\�cp�كQo����s��A1��-%�D{�8�z��6�)��)4K]����s�-@*d+w�w?ڽ���G��	7�����a�����V�}u�'��	@3�5��_F�d���~�}�߲Wz��g!Cjb�_��y��0�`|�lh�='�gbF@;�=�[�o�!��CΑ1���V��W�5�ӖBQ2��.�'�pF���\�JY@	c;��E����~SUwr��4PӹY̦��e���ᷞЍ��׏]*�x&���RuC�pR7_:�v;.
�*�屄�{6s�e�����6��r�`�}@-j��HdS4�Ҩ���,d���-���Z��({4Ԋ�i��/��ؖ
�dK��Q;՘�����I��v����\�ML*�K�ݮ1K����3-K���f�>6�6Z�p��H�TQ�lg-�D��Opb�����J��яq+]��x�4Ҙj��{�A�S�0Eo>��={�كj%i;:]؝4��VJPs��H��SC9w�E��D�4�K��������Ig�l�w��?��[W��X��hNQ���@n�g�,�y�⣗�����7M2de~7�D�)'ʀ���[�8����K��(���	��$F��G)&�2^��g�����R)U���f�a�F\+�<��[Y�At�<�ʝZ b2�n_����M���Q��Dy UU-�ܓ�C�H]I�|�$�9v�8mv�j^w+7����?>ʠ�]*���Hj��m\&��4*�؉m�VYG�_�K�A�Is4����'�GT�6��y�J.���	���ȹ��Ċ��`�C��/��1d.��ꙏ��>�[ӸY.��d�͜��E��o�Qb�F�a���d��	�%\�m���{�"rl��t���6�'�QPO���qL�]�JT�+KVΎ1fc��6]SΘ��I03p�W#�ֳ@�mC��x��H��OG�rW�"�����I)�8�H�:���U��t�2$��+�� �d 8Vz����܌�%�Ol�sBYj�K�YJ�pL��R�M��OE���j�M�x�wY��W��5R�=y�/(�����j�I4]L\-�"m�x�p��4_��C�Z��w0I0��x7����n�2:�Ck"Jl[�o���*s�v���&��U�?u> ��A��m�|���kuIn�"�|g+�q�{���aO�q��r{�BCW���l�(��n���	q-.21� ������Hu��7b�
�fN:e�$i�Ma��v�U���������� � W��r�����+�I������z��DA�&�54
��pJa�0"V��KbS���;���M��7E�07SA>�.�D�o��8����wV�&Y�V��<!	&�K�L>YC��Q�@�|p��㲻M��\Q7����rS��\��Aa�\7��<9ѵ]HҢ2m����ۻW�����!�}ԫ��U;	E]`G3�c�JD���'�{��P�{T�
=aA�`6!$fiZ.���-�ǻ�`�w���u�!Soج-�Hɛ�3Xy���r�����w�~�QL	$�i�)��>�@�����[�f�`�����Mժfk��Е�u�����k�N@ցP^��[�#}�m,
.�53T��~4v�o�YZ�m�k0��߂��n��sTC)���F=B`�G�K�!ӍSL��Vn���ױU�xr\�9E�}#����nC٩��`�jw�bEy�щ�iY�0�L4��� `|�AIf��<K���ZN�CB��`@�8�1~�)~�V>��=(C��>����L�̓�'jn�G<��$HW��9��qݔ�$���?������x��������t�]N���2u	��Qn]���t�����Q���Czh���;oZ3Z�_�?�'�N�7v���e6Մ�J�a�5/6�ռ,�b�E%1Dy��Vg��"OZ�blm�v���0�
ѵѾ�c��v��g`�s�	����FA����t�Z�.�߁�L���o0�"���Ǘ=U���X�N��^��h4]Va�'���R����r���v�����m�Z����ۣ��&��ѵPZ�c�R9�?�Vp7����0�@⣓��{a��R�>څ��ʪ�I��{w������7�K�%� �>7��pJ�16;G��ᕢp�Iv�@��ؑ�U���Ε����(�W��~�+�4*��~�� ��$+���V��̿&-�3�X��º���t�˴�u�a}gYI�����~��l)��'�`��c��ۿ"R��^ގ���&=�_i��(DZ�������kЅ$�1��Xͤv�p�6i��쿸��Åz@)$�q�&>`��k{T R����}�,�o���@�~�/�����u��MQr��$�<!ޜM����ס��'��?3�Qw�Uf���=ftuh�D��E���/�����cJy�
�r�sQ.7�dL� �IGy-+�n��i����(���Ũ����m�m�?� ��\��a`P�aZ��R�e�
�Y���L�[�m��
�N��"���@V���b�ӨU4G���ky��D����S��Zt�k�����ot�)[��+2`I[!$kh��UE�D��x��V�=�/+9��X��U+��7��w��4_Oo��<���j�$��z9ՃHY�0�o��\�_�%V�p�XÒK���^[}�fٸ-��JE5��$�kX[�tN	#䶠���5+j�l-���h�[����?�[d(��m��g`e��L��(��f&�̲X\���� ��M�8i�7
�d��9x�sB�~�K�8X�o���ZSf���(w�+�O�҄��Ӈ�}���Qnu&ᣈ�����6;A���R=�R��	���؁�C	�.ldK罺	��f�&3���,]�`������/?_�-�����6v�F5�Kˆ��4�M�Un���<�����J�@�.�MD����:�Ud��c��X�i^���
��q�+�I�b��6�hT�X���`r�TK�\�;�P������5z��
��,�h.L7�;*Ip@n<�H��,|� Ȩ����n-�����9i��Ʈ�u8���lx����8�YH�����w"��,t�`�7����+�Q�4&���R��Xҗ�����)$�J>�#�e7�8�c�哋�(@(�.�h��[ON�H$� E�\�7&�k%��{g�d���O�+����Q��s���1��J ��x@6(��U3 ���Je�S��B�+Y�2�~�d���־F�h[�/6e����j�\��p��hQ:�ń�8��$@>�ڬ�YW3-:�

ڒH�3
w.�m�q2�@E�]�<i�c�?%�X,E^6A!��$_���~��1Z���Y�����ù�Y�������F��Ж!u>���z���A ���c�O���ZY��Z�ۉ?Յ���c�;��$��0�3|�Ԅ�.�ɁYU�5Y����?�` %Ʌ�dT��Zr���6Ɔ�8�q��i_�L��ij�Z�X�N@���*+��	�mA�[�%e=���͒L6��`���9A���:�J���U��1��/K�K��5X20��a3����?��`�6�ט
�*;ą�
�~<W>Ƥ���Lq�M qo[�:�B�a�AIjX(b���V��^��ǟ�L�����J~�̈́L{1^�����퇳���ҹ@>5��jL�%��M� �3�VzmJ�k��N�������������"JOdH��j̮a�}Xjv:��oS�{�l�'�e;��0���t$oqnZ�9c��inCĊX⚇�8܍��Z�z�4�o�u�*��8Ug��Bj�a���<�^�v�u�H�9|��e�
�D��5�	0tψ��@R���o��G�UQa�M�I���c�)aG��m�i�h@BvЙ5���z]r���AU:���ضzD�~t�Œ!{�`�i'"�#H��70t�`LYC�Y⠕ej�)�Fh�����ь��O��b�_[�b�ƩX�~�y���_^�k�0���i��}�e�)��b��q3w���]��x�t��p��s5L�U��fe�o���4`K�����l���E�zb�'�(��T��'1��&m ��Q��UZGU��=vd��~�J{J�������(�V1�)�N�������F�s����ז!V\<�*l���}������[�}�j�E�/ʱ&������#�e8�3I�A#������x2kP篂tv���'m�\�~�����4(�6/+fpR����߁�1�gbϝ���� ma w���]�_	]�Ʉ���xc�>��q�	�h>|u�z+.���pɹ��[\�G��Pa�V�lB15��!�>�HP,\w=1���y�FN���j	�'(�Tx��L���u��܃��3��=��:���lW,H| ���*-E<o);zB~�2��_朆�&q/:��&l-TO��m@�C �P#M�t��ҹ1���-|�ni�(��AS\��"�ُ�EVO!EZ���x諲F�I��>��7_�T�@��`���$�e��*�)�>x�یx�hG�i҆���9�����^�����̫t����,�OE�q�Rs9C�ņ�<�h`�%����v�	��e��ޣ�ğ�v��m����[-�f�k'�O�1�/�;�2l�,���������6�kV8{|ѵ��iQ��}�}�@�J��K� ����]��1�b `���E�:��l`��&�c�R�'yZ��ٌ��z��O���s����x 4�ÿp�RC8���`m�&VE����p#�ͫ+���e��l������a���.ɋT\��$q�ذ8�QTK���!� 3��/5�I=u��~eY"�Y��eW�웆���?I���� 4g�vnLt�|��H�Y���"�\M�d�9�aX��l�[4#���uЩ֠I����ۀ�#�7�]k��)�T驯2F&l>װ�V}�g�=-7�x�#�*�60Yf��:�t�le"��M������d��?�ϲx�k(m�3�N蓬���fs�;i�n�o�l�9�8�R��<�^�%0mKm˂{)B�Bd`y�'�$A�� F�w��10e��]��5%Qo��g��X���h%�����G��R���u,d�S���X��������Ra�