��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���c\�esR&{������o�T�e�Z�/��`%�����1�2��g\D"[ޏ�F�
܌�)�u�lg�h���T�Rfz��9�x��+�E���6FdS�
��:<'���9o� r���l8*W�V��ÐP���jv�,���9�C�B�"H�`�s�8�:��dg��,��k&~~��{�� ���i�`$�Pt�u��)�`���:��t�9C��:�
&Y/"���MGs�����P3��3�͜���ҢA���r���!"�Z>�:����<�t��aր.b'����H�b<\�NN(7L
Q��ق��1PIo���]�$'q+s泤=tE�]�S�:��r�����=��c��̂���u�0���-?� �����e�J�Ƞg���+�����Q�5O����c*�k�``�K ���(�75+s�d�/�7����oW�4�����`�7μ��L]�MhՇjk3��L���ib��[��{�.�ju�?���R���lk����o��r{��r��=i�x��蓄��y���W�d��0�u�q���y�ޅ��kks��W�*~��L��{^�%�l�I(�b� ��5����ѕ�(5.c?Y�q;O �&�m�����'ꮬ��C`)���DN���y�CQ@:��r���'�o[E�1p�׮���8�K���%?&40���w ����Q@�g_� ��=6� �jL����y�	�|���/E�p���2��lyV>7�C��Q�6�r'�x���d�,�h�Sq�GeـF�}*\��1Z�t刡��se�]]����� �h5�
N��'��D���E�e�~ly���G�C����V1�\5��mݎ��u"�0��%�e�n��ѶA!�=��*�i����bf���qc��SeX��{��� F�W�NV�w 	�+�n���=_�/��ڜQ�J�:(>� �� V�V>a1%;N�.���Jt��I�bib���+�+V.8$S[V�hB#2z�A���8s�z��Ծ���������'9��P�O�p����D߻£��>�������q@�ŝ(Ni�ߒb�Bp�8Ū*d�q=�6�ИC핔��o���	Y�lٛy��^Td�jB�v;9�`ܼ�l&�xA��9�+��8����X������Vu[nH��?�!�֏%HS$�g�\��54�E��h�om%V��}�C��a�U��ny�����	�U&g��f�_������q�k�扺E��NJb+�
IJ��b� {��Cz��.~�lJ�E̵�S6�6����
e�8�)>�в��:P%z���z��Q�Mi�J��:U�A�cgV>����7�f�F�9S*�8 [|[L�����C;�³�?���0��ۗ�Q)��]|Ͷ��|�����khx�r0~��U��Q�|X��5�Q�J���!��|_R�{4�����	����3������9./�'������:�%�_*����y=��	'�%�C6����1�� JNB��؟Z��}J��z�#��1ۨ=�F�+������fmx7(@��P�L���
�".7����*���t.+�i�z����#��=]�*4�%�ui�[���#u��(⽝�ѽ�HQ�IN�D��Шc^��V{���K�����m��h�{�q���%;���;�`�b&���M2���c�U|�֥�Ʒ��Ƨ������M.ٺ�QQ&����tF��G�HqR����b���6�H`�q�����CN�|)�@�Ts+�
�q��|(V���(|U79��A�jd+�Ws|���s�M��i��$/{K�W��HCk�A��x�����`��T��W3�xrϰ�<�m´H���� �>�#t���8`�.�������ߒ�eO{��T������ۤ� ���	6d9�i {���1�����e#5�u
���&R���[,L��W��bڤa)r�h��aќ�����G �@<�8F�w����="��	�ں���ȟ�cv1`���-�\\�����yPq�֦u��Q�|y"kŝ��D=O#Mȱ��Y{`�U�2=��n��hh��a�8��d���%��ӵ����JA��>���H���Y�кl�(ϮUs���)H����Us�Z��z��������V�xZ2cL���l?���G�f���.�<b�@� ��FV,������������Lw��q?���MN��_e���(�$E���WL*��`J����k�ؗ!�]��5�ZI���S��H���n�wk+l�=��xw6JzY^�A�g�s��}=�\W=���9@�0Br�=t%�N��_<����[�`����׃��L������q��|8-��[�D�I���X5��xVҠ��Ң����*�Ք
�i�m�!�7��D�}ؘFr?�V��ѹ��6��f�X��odIIhfu"m<��@R����(Z��
D��(j$�9��>O��H41%��i!KA�d!�(��<k��h�����N�x�\�&K�����5N��ϕ5�k~�e�]Γ.���#�2"3��_����P�&�n%S���9�%`�貗0��ӧ�w|�셊��y�LC��ťG�3&��HVX��(7x�����!�8�c��o{�����=݆�n��θ;S�S���}�I��6Nk4��{:��X�:6��[x�U�������OkY�.nV�4���i������s-7�;, 
ws���SR�ƭ��O"d�Gi�r�B�|&%*�}Œ�8$���yH�����'�Z�$p.�9�e�r����Gu��z�-�� C�+�E@1er�Z��������Jy2�٠O7(w�"P�$��H	�s�g����7�ȦQ��j4�� ������m��K"��i�.��Yя"*J�����q��I�f!��ES����1�iR��8����5,��w�,�[�Tǣ��5s�_��b%L~����4�=U�r�EX%�B��$���⧂,-�t����:�����k�K�LȖ���-���T0��~?���u��%Z�$mg�Q��?\o�2��W�=�v;���<�#6(�e�d(��s4җ��YrQ�N(��������!OC��A	LWݺ��\�ؓ��v�����M�Y��*u��7��a�p7E/�ۏ��� q��:pֱ�+�V!���_������Di��F������GDÐ`��l��������a`��e� ��b�r�0��'&����@�|����vT���i� g�4���D031p��R���~g���<a���-@5�FE���K5�뉦d��:̑}p^�MN��X�mb�r���cKy��kY���w��W��BTT����U�p��K<�%@��F/����I���*q�Mm�'m�L��ej���c��N���2��%�}�[�
[��ZW�y �����d+�k��b��	@]�t_2�Ųbҳ����)C��n�a[ H�w��:��)�/��_�����Y�}�4��)WE�{�B	e�R���]���j�I�_��2�sd�ѹ?і�;�c5��A)�IJ��)��7�ۜu��?�wRW^��,��i�e�\�7�#�C�p�V?ѱP^EZ-��,�/��KV5�1$6M�\�s��䶺�uG�0�`�������Nƚ5�;���Eᑌ�}���W6i@���X�h�k��C~�iz�D{D��C�%�������-�UA&�0�L� �.a	���X�<�=c��Q/��鷕�5r��?tu��%Z�D�l�:"��b���j�`1_9*﬏4_�0T�A��`���MYk&�V�DZ�����n��gXe�e>��k�B��e�zn�3[
�ۼ� ��'�eCD���^8�������xfSط��8ߛ[Y
T�ԏ�+��js�H����tv#ˣoo�u�W�z�*\p�X_�����Ŵ�<�ȗN�z��U>)�|����<
dq�$��_����!4JB&wD���'���N:n0�DN2)����gg8��g��[[ޖjB��jޏ	iq����+�j/��ouɷ������tmfy�Y\�O��i'���� �,�?�@�s0Q-x�M�4��8��)�<`׫����d
p΀���5Aq:R�2t͸?��ΘjED��X��O��Fn�!�Ex���4���퇆�et+���T����;��`��0J�\6��[0�D�ۻ�%�&�p�\�n�I�����Ϫ�ZnK7�i��o���ٷ޵�Ӎ�¹{�������J�p(�as�� ;L�s�ܣ�d;G�����k6��`�mC�
�(Q	����ޯ�ϒ���0.,�D�'xF,#ޫ��eY�3(<1jJ(9
(A-pIK���5VQև	��	4�T�{."V���Ou��?�+�ɓ<� g�e��9�(K8��R�\��D~�^驕�Ό�3%C���j�7����'[t����k.��̽�(��d�^������M܄��J����i��ld-m*A���ƹ�n,���ح��-���
�[Xk��~#8��L�t^	 (�VQ���S� ������=���kǑ�U�$���o�$(Ú����$Gh� Ö^4��Ś�Z����@���VI�+�����*	�0J+�?*q�̭���&Y� ��^Q�;�¿J�nW�Jt1Pc�L���/A�#N�cK4��u�}4�e��mڙ��U���6�BV&@�k`Rm'"� �4�H�z=��H�~�s�{��m ����b��.�>5��~Y��~,����T������$u7�8��Y�hU�%I���@�(s몲3�����}��4��[]�V��rs������8ؓ�,Ȅ���3f��KC�S��
�2k��Ĳ���~�t�w�8S�G�,B_������y[����|Z�(g��M����#X��Z�m�.� ���XG�q�Fr�Ey��4
�|4uۏ�:���@?O��/��ث۠�]��U],�U�n豦��)}I�E	Mm2ŋ�
��춬�1�ɦ(%-i��� �ЖxZ#�һL�x9q眙eR�X��߮�Y�����Ӡb�y%κ��EkoAz����f�rH<��6�x������|BXs�3��>�tsO�����=�� �\-V4e�F���N���F�= ;=��h��(��07!Y�)���6��tY��)z���=U�sAN�0�`�i����mY#jt"_O��p_D�=���-0��q6�4�s�h^h#�)~;��W�Ce�&���n�.�_t�����l LB�p?�V��<���4mBJ��&���-w8� �����6�y���9��ގw��Uc� N���ݍ��;8��k��D�{c��.ש[/��\G�ŋRa�'�&�-U���Um37�@��.��
�x�D�w ��:R4��#T�x��׃�.��C�+�L��H����_�Y����E{��5�J�-u�?`�>z�����"U4u�ΑV-�Ny����jyaJ!42�f���[������K\�H
x�Ʌ�S��؎� �R�T$�E~R@��ֵ���'cEw�:�G���;¡W� 9�r>�=��<���r.j$����RD�#��̣�!��G����W�����wM
��
0A��#�l*�b�-�%�`g��<k�p�g�����XB}ђ�d�Hm� ~w���=�IQ�'���茩4]��$�&;g�a(a.o5�h�
��o�����Ŗ�4�V���\9І�?�,�'J���?^�Z��&�X�,_����ό�L�&KhD^3b��\_�� %\��b���������K��XU����}�	��2��#\'
�8j��~6�H���������z���[1P0BM�i|��w�ݥ-��}�曉�}| *!r���
����nͲ)��(&�v
^�ġ1ϡn�rjNv�6ŊuX����1��B����D:&�\����v�����n�j�<�.xhUe�����)iV=
+�~�Q�NbQ$�F/��WGd%�m��;�?������W�����J��,=�1��f(e�4j���C:i˦����Eـ�`"W�V�J�B���Z�"��ߨz�9z�!�G����_n��Ft1ۃ�?X++���3	���6��]�y�6��ޕ*��$��=7�.��I�Y���dP)�����=�`8s�����&�=�ĵ���TdF����-%'��t��w�2_Ͻ�������2�A��k=�~��Ȕ�R^g@�u�q� �x��_u��g���B��;KꓹJǡ����G��:}�l+s���G��/
����L�;�����0=�B��:��)��M�����:ԺwH�g�Lz�}��������X��n�2<�a�D�˽�ة�t��~�\��a]`&I:��g����aX6�r����QH�K����yT��M���u�����m�9��nl���m��]H~�^�@�{Bl��I�c|1OSݿ6��?)��19^��s�$�ܛs�8�cH	T�qf)`%�5�5�r���e.΀1��F�Kr��#.%�V?�	����d)yz�v;����2� Ԟ�)>��@�Hy�0g�Q����"գ�y�t[���t���6���/K���a�H��g�r+<Bf����<��U��ۆ�vٺ���m��G�/���]1\x���Ǐ��e�	���H����o9f�~,y���Z���@�-C+o��a��?�V��l�T�����%i8�ƒGj�}��[U����@D��S��pH���!�K$;���b|�#(#�<`u}�U9ړ-�Ș��/}Ɇ&�ʙ��B�c�w�Q��j����o}H��#�T�r�p=zS���649��N�?�t")S+�S�_�r�C��I�r��y�I��4/�{nj}���q�w��R"C|��n�b�2�� �x�U���}kwyC�MҴO˷z�
��>	"y���)��l�U0�#��ٛ�h�<�G緳�8���#��X��Y?��误�Hܥc��Y`�n�Uפ�\���U�������U���Eu�&EVPЄ�D��/�ٴMX�Zwʎ�%�;u(J�:כT�}q���R��������-H�떾��,�M9�E�H��̔uaGҬ�p��=� ]ަ:�u?��43��q�2_m�a2��O��2-eb�Vƈ��i��i�vf]����h���/���"A�@����7@�j�-S��d(jv$����qsN!ߑ�7��R���T���t�n�U!��!J�z95G,�񓯳�LضG�c�Ťن�ŀ?8��װqc�#f*���z�L�|\<��z�e9�e���	���E�n�_oo��J� pf�Z@�U/��^-�E|��Sm���qv�+���3����l\pKi5m�������U3{����P������z�[PZ+�)l��8�������@vxF?d�a��)�0=$d/c�È��b�:�Jiݴ�ޮ��p&�$�������6�|�-����a^�k�@���2����R'�H|��2�NV�[���Ů�~��O������Zo�R��k.}�	W�5]�^��=d�i�}�3x<	5��N���jk#ҫ��l�*�B�w)w���#�Q[���/��B'��_Jzj��~�V}kx}�/�Pzi��^Ą������;?S�]����:�f>�ݓb�<�1Z��e(P�'�]�mv����}��x�@1��Sȳ[�4p�t���~�tQ<�ފ*�%���w�(���vDc\�~Q���R��g���[�ߞ�S����U�i�pt2�\>�����{�5�Yr/A��j�Vz����讬�-��mK�S`��Y�Ru�ll��Wm�K�4�m]Տ-[M���g���q���υ�fS=�X���.����!�}ŋj>;C1�N>��p��R��6y������҇V~=4�NR���$R9���%e��IU+/�,S�|�[��k��&���PA�vp���������,7[��d�&Ej��6�|R�����኶��}��E~��Y� ���+�	��~��������Wc�� C�n�[ъ:���a�=wm	Z�TTV�m}a�Ͻ_���O(<�OIN�7�ƈ�����Ӳ���0!�p�L�5�"�!x��fY �w��|B��Ѓ������S��_�ōo��1z�EuX��<U�V~��t�Msq����I��̪�*n�[�#I�P�m�t�5��l�Sqb~���6���/��8��3��Ь}f
�Qy�5�y�W���hG����h�G�C-\)�*T�5�][�nU~���2H�8�գ�c��HMΊ��]w����Q�qJ�^M M����.�G���v�o�g�3huڇ؂a&>�d����o(���/�����j01����[Ƨ���eVe$��r&'�.Xа/�Q�$�P|�:O�ӗ��uŶ����s���gܵ_l�Y�#���Z)=�����q�h�Z�+-�����x��1&�t)�?�	_��F��EF7�]XG�����#��WrU"�N��k���	a΄[��G�"�/|�C���2(3��0by����t��f�{�Y�'����&�|f�	Ty�4��\���N˦��8�=\���a3�e���<9�ĵӷԛb�.��.���##�O���;���zG�U��&DxӚɑ�+t�h�LE��33ʸ��\��^��1���� )q��ݷ��X9�b�tT��
�łZ~�s�/�L�[�J���jmפT���WS���w�A�֓PS�&Ob?�?�[+8�������d�m������`��������Tʇ��&��5�P�r7p���%'J����t&y��slZ��Qp�C8gѺA�E���b�l@������,K$L4^����"��uRe- �KoF$E�5ʈ���$�G�3_ �5�����!5m��#���8t\����N#���)8���|���
r��n�J[oLk&^��L'�,��F�p��4N,ي	Ђ�$$/��OH�K�УwQ ����6B*�p�|�v����K�G1�&f��f*[#N���q�kJ�7rd������� ��n�f(�3��d��!��M1�n��5:�_�da�y����o�I=��5j*^��&K�D��nb�̠nhވ��`�-�"�S��u��r��˲\�`�y�����1��h1����
Z�����m&R\rIA��E�r��_DQ��2j����Q����[H�k���&q;���7�$RϘk��4 �9&_*��便=o5�-ٲ�X��l��o/�\ѽ~��,��,����<�����^��+���>�}0�� �0��V4Ǥ�j�9݋��vP��˳jJ�.K���� �YG��!��*�97B@�o~���:�@���#%��Q������f�v�y������&���ێ�	0f�H{���@�����5u˲ V��?�3�Bu��3�-`����f�l��ѵK���QD��f�8�,w�D�E�	�	���}�Q��ƒ�uD['�2��%�-��[@��{�}5Y���;ǫ�U�L���!{��gT*�NqN�eQ�U�}%S�A�^�yk���~��o��ZEA3�(� �&Ӎo�]9�2�,is鉘�e�QNC�Zn��hu���d�[���1�A ��w�Zh�޼݇��.��
��F�Љ��a��C �d��/UQG�?<��~]]��w�/�{1�0��c�:�=|�\�1(��&^���:��䡃��[F�`N@i_�Х���K�^����1QY}3�c�V��x�]�RQ���R�6s ��9Lݥ) �tM�9�5���.'�}���`�{9�,�����%���VάK�c3��
��-�?մF6���l�o�ϣ���f��A�@�T�|�l�~#��-Χ�݌�s���ꐇ�T�W�Y�4�o#s��Q�p�EG�D��_�5�[Ҭ�AO��х��X�ܿ�
�^�D�%��K��p*z� RQ�NE�UD��3�������VuF������#�G�C��j��+ׂBޡ�Z1�-��u9q�w�8�gI��lؑ�v�Z?� }� 8�+�/ȕ&���{ {����&�;	���0W,�7�A�,�?ͼ�᩼5�G����M�bG>����]	��L+VDЮ�������x�rP�VX�C�l?�,u����,E3�}>�.�e[b����uQ��s=9f���$�6v���~����=s�c�G����T�S�#��e���Z��
�@�T(����sǖ�͏���V��zg6P2"���#��&�܍Qȟ�nrO��wÞ��Q��}A_?�5� ���I�<����ڦ[�sDf\�
+WmU��&r��O����n8�jmV��j��йB=�1����	�� ��y�u�S$ǯ��'p�pɼ7��I�K�,Y|Z�fR24�8��,j�� ı�kw�e�AR����*{ǎ����Pa� %G�a(�_�'�<ڝve��F�Cj>�	O� LON6Kd�Nx�ҳ*Φ�>2�2B�Znh�s��pL�M����PӥԠ��c�W����x�o@v���a��Ὓ^�=�>�	SΓ9�S5�zy��3>�5�-�����������:���Gf�3L��nl
A�wT�:��Z#�}���e~�P�d��8�d���^�0RT�D2s�%���'Y~�1B�P/&!%[��
��6�|n*�C�*j�m��� �5+�(p���#�G���x8��KQZ*,uܲ�Q��9�ߜ���O�vb밙I�17xCLx���Q/:=S'�`5|�0'���B*y��$މ�o"��sZ\-�2`SX�.@m��� =���oA*���w	o��_S�V��U��W�W�Q�>�~�q��?�7ݜ#[������:��J�W��ܯ�HY���6c3<���*�E��ڏ�	 ��`����p�k�)����$.�Dأw��ɇw��a��(�aj��Js��8���\�Q7��. �Y���q�)�m�s	�~(úBJ<C�h�gh�SQSy��`�-y��ת�R�k�.�oG�}�;0M��V������E��q*�y]�t�e�ϸ4�Zܥ���B��xz��9��`s�������:��� ������C$C7�f0�s�8V�yHka1u	z鯃+jc-��#0���v+O<��l�G�� ��!���G]΍mYe��BB\�O~Ƒ^�A�F{GN�OW;�b*ԩ}N�t<��-�R���e�]̙�d>.���<�M���1�������a� �����%��)��t�[���g_���Q�������t��Ū�<xTB'����]HO���Pa�ڔx�8kf�I�o�tR8�i�N��_���u8�Eq�3�g�2}�:Z$ۧG��;�!]�P��3x��<3�BM�vj���0P-i�M���M?�<颵����H(j�S��ȥ�ن�	�^�'��˩J�r��C�H�z��"�&ںTN�?�R�!)薒8��`Qm*��a2<�3g�P�TR�|3<4�g�;B�߻vq�U�"��� �$�Ͻ�ѽ���W$+]�<���0໧=�O�v2�Ci4�
<�,����!�kGr�v�CZ-�H����#Z.�_=�z��߼D�ޱiCH9h���`���h#h�֚�#Y��6
��˟��*��8O����r���T�ȃ���[�5�l+�=��hP�O�J�}~�-�#,��ɯ)*��i���n����������8鳋���o5���aހq�D�UR��C�����q0繸�7m��w�N��$�ꀈv�19�bˉf��숣�X���i�g�>	��W?��ro6�3Jj;�? ��T�B/G�]��e��I���?_4c������� �\6<��|e^u5�~ժzsxm�L����|�\��(���8�O��Z�O��\�h P��vI��4Mь�uo�"�|U'�/����)+3�S
���[n�����]������&�U���	ט��6�����\#����;�X����gָ�녅���[N0"��;�֣pȃ�`|�Syh��nGWb�o�F��q?g���@�m�1�TM"a'��7�;7~=��՛3�)�!��!J���I�>��vK������;Դ�ba41�L���Q&��C3���ea�_�p���J�&i{js폝�� ��\ɕ�6�Ep�d{���W�@j�u�Xp��Y�=�WԎ)i1���ah���Պ
�U���l�˕%��\�<>��&VP��ŝ���&Y�b����!���ʻZ��X�5l�Le7u��:fZ���(5�9.s�_M��o�'_�N�����Pd�.��!Ɯ.+`+��fL�~�����60�{��Ud�6I�5$�I�$G��� j� �����|�Z�9�Yb�+�;��W���������zŰ#��1U{�HZ�;Z~A(4�:rf�lO1a�^(2ۋ_�6+E6�X�ME1ņkM�O�'�{�[��u��Gˈl@;9g�N&��� 7��/�:�`�΅"�7^�y#���Do11�A�����dlf�O�V7����~iQcPeh�N�H�0봦r�)a��~�A����k�zx�����X$��y�3�.;c�@��e�Z�2�.n�y{�7a��d�pN x���0D����%З�K��|4���0ٗ����ڇb(������%��W��o�I�;�H�z�g�ݏb�A�1��[t��}5I����0 賈�:��'�!�0bI�0�i��F�>�K�7�mйG�fz$wxS���M&�W���t`
�u����PSK9]CM�ܠ��~sB�Ce��|���-�I#m������[��PO�EF&�����"��D��m��H��"���5ơ+ac�bG:��&R��L�O�7rS��;���i�O��v��$�,�c��� t����*�'��e{�&������4)�a�܃�r��.�Y�U���~¬�+��K�AA���J	=/�����"���[�aN�ke�>椩.2<��QluY����8��f�����% vKӜ�Q�o8�
���{fD��+,{�	+��۷�>Frj�'5	��Z9B�>��qђUw	󗪃��D�� к��M��!���u��L�������0+R�<(Zִ�$a�h|{ȁթ;���WzU�ȯ��_~^�c�cچM8 h����?.1B�"'gw�)	
��-!�/��65f-^56�:\���R�{���{(��!�I2�dLL����,U�jK4P�ȋ葮1O�����o�����ą{v(������$��lI"�1V��D!�g��R�۰�{����KA�f)����Kh���ڃ�{ΰh8�8�� ZN=��D�rW��E}3�d����,ǰe�}T�x�T���B�l�@8���c¹5���2����1����i��dGl�&�v�4������]�uMŭ#�؈�*y�@N^�ĺcB�anH]�,8-LcԀn8Ƅ�z�[� ���m=5KGеkd_�*��
�?�)p�ɼնkw��,n1��M��}����pW�PY�֯�v��["_�*F)t�Je��ك��~�`hm����!w6I��/��X����I�t�@.n���C'k_��٤��=������v�;RItE�Ѣ;�˜^9�d�b.!���k��3�c
+������2�TS�*�爖��r��?^_��n�q5Y)�xL�x�4X�NθN�MNY g�����=�B�	�E����Թ�;Q���ds�hF��@���c���[� � _}�:��i\R��8�R�p,
D�x>����1�<I���8��g��U`��)-���壀�d���_�ҵ��7^��6�YTV.NyK0a����S��1�_�-�["�j�XY$.�'�C3���J׺K�@k�Խ�el��!W���!�Q<^�b�R#����/�_G}�m�M����j�*9^Z
��XݯzJ�b����܉�5��Cm�T��Q��xL��G$���l4c[���)��}4뷛"�a��d��>�Ά�X����D�Lg2䖱�G'�>l4��FK�f�:t��;�h,E�
�K��[?<�>��1k(M};�� ����7���RQ��O6�m6�P�$�#j��Ŧ���R9� �E����[y^�vi�_Y"�̌�G���:?�+����+��Y�ٺ=C	�����|l�y�(��/:�r�c�������c�PT���˸$j�
�U��=�,K	=h�@T��
���LuF��M���!�%	������)u���z���l� �6\�e2��k|�@�\{IW����u��4���1�Z�� �����c���-����߅恽��3p�8�� ����M!�fS~��EI�a\U �B�S!@Ȕ�b�i��Վx.X�M��!Ak�	�xWp�ч���.��T�C���sS�� Ϊ��(�ss�@%�lr�,���~\i�ʮ2���m��uY�'��Y��P׿�8S�kȉ����ym���paFѪE�c�=7T�<=]s�~Q^�K�ht�V�k�u�"�wVF����������&n8���5��S�~;�PTS�,�F���2LD�Ѓ���>�����Dx����M�k�*S�s��=�/��bX9���������������X˘j+J(�j`�����+��.1��'��'X��(��WS�W�0�IHd�ީu���T��_��kfߑ�����LT��c�aq���O��?���i�@�M�OG
�D�T/,��\b�����Mx��N�4 ��ʍ �SxU��H�O�N���Q�ܖ��AVR�MP#9B\���4���͵�n2�C�K�J(b������3
T �ׅ�%�Pj�k����ҖE��֒�c��j����j���v-0�Pi�('Ү@w�>$H-�y��v�
�Nn7���e�M���컋��w�D^���4�H��e�5x���3�X�����น�����"p�Zq�&i�ަ:W:ܘ�
�[/�@p��m���_�{_֥z������\����b/�/���p*�?z���R�q���㸿��Q���Qd�#c���j��hs^=a[k��������זdk� /��W�pݕƘ������_N�R�'�	j�3��{pF\��5����Wl%�S������R��#�?���'��/h��-�/���E��Z�pָ9�����K[�����T�2e}��.���,�caV����{Q���Hӎ�̅�������x|�a5�8�����}������Y�����(�үq��	��$B�����(�ð`Kt�HS�T�o�:X�����L9_ՌdS�%���Vo��D$2���hm�
q���l_��:���r:���a�!�=�J9+�qjAzm��h���b���'����Cf��M����ָ�ȁn�J����� 	'�����Y��g1�ڮ.�����ML�QYJa!#��X��4)�K/����od�!_�������Y�&x	�kZ��(�D�癧m5����`�n��
��qH����֊������8X������b^�BOƚ(gO���N�D#�M�Vw�?�qUҞ�N�7��O�)�M��T�C�8~,��L���4�fj� &���$3���2��+D��͇-/>S�п�+<�ϰ8{���N�w���X�{gѠ���=�+��d>��㫖�Т���1F�F�@�K�4�2i��ق\#mz�����_�)p~Jg[ݶu��~�����m���*�҂Z�(��1w��(c�������p�L4v�VL�<�Ku��Q�Ȝl���T&�ҟH�8����&��`w��*G�f�6����Z��I�,z�*��nz�{��G�rj�A*�
��:Uj�z]ƣ���� ����OH.����#���%ϱ�0 �#��b���r�M":�ޝ�UL�͔�4Z���Oڌ����)�>`Oﲑ�-:��"��f���`su���U	�13�٨x��1r�)�vtLhCw�e5��cE��5'���75����eC]��(��5�M�m`���|E��#E�
3�����?��=�������~G5�v"�YVE��C�d�j���1!Lr�$]���ѥ�\�S���h{\ŉ�>Bg���=�#Q�m�¿��y�ڱ�����"ol����
z�^b�'C9�yt���ϫRՃ����6�;շǹ���Ꭳ�jA4ƆW��a�!`q��7U8'qߨ"Z���6��#�V>�ɧ�]��{n�&�v
����E ̨�E���M�g�l�䳴U2��x@���� ��]��2�Tػ�~c���1~sx�Գ���nu'y
��t�	;���q�ῂ�-/a��i��^+�e���%�nv�<E'�f�A���Ღ��t�a{RE�`d��a�R̯|�8cv��C�آ���?�s���{Dq�:�s��dQ��_�ߋ��u ��Y���4�=EQ�b(�;��cԚ�	�\O9}1s�����T�«;�$�1Ҩ�:�� �`�+8��<=��7F$���ONoi^��~�.""CC4�!�d�xy݅(��`�׭S1�����:�殴�hw+����ØM�����[�1�r�ֶ�Ǎx88Zyu��(�n��r�Q��x5��y�Q�R���a����5�RI�/r B��)�@4p����1G��ն4��]��	�<y�㨅��L~�0m�i���%���k��=޵F%���-�u��b�%Q��t��%�s�%u0�m c��@��{��[�a'�K$���&
����;�̽]�i ��ݡ1�6,bĘ�����*n�i�xJ�g|�!a���yԗ	L$����ڬ!��^L�v5i��(�x��X�����3W�CV��ŐR[��ǲ�j��T�x�0"�C(�2
u���5��dO��V�v#��b>�3	��V��I=ʹ��m��"�8a�:�a]�'��v>�.�9���%��}P\��ؗ�����.Ĕ�Y�T��N LxKu��� �a���{6�)�v�s�[�T)�J�>���f�!)�ߔ✳A�g=�f=�|�����w�٤7�`���qӷ�/TRY�ھ!��1�i��J�)h�����@N-�0W�WhA��$Hߖ.7���S��茝����i,��9T_��b��ێx3�����s]S�um۹$_���U�x'�(N*x ����˫�A�0-wK��N��h׫}(!��!H0�c���f���CFu�ti|�z��4]�����^�^�����^��!�:_�����L�ƛ��v�/�F��ʨf4g|�ͫh��R�v:�j�<��췮Կ^p��.B^1C��l��P��cwk��A)N���D/�f��hm��w�#E��a�Ei=ȈHo8�.�M&.������E���DU�b���
��cэ|��*Z�a���|eW�������VV�q~^�ta�RH�C��Q�+'!���DGp�wE�D��b����K�#
�Ɏ��b��ׂ?���ԥ5���ػ/ލuǿS���{�'ǝg
]NhmI�i��ۃ��ڍ�~Zg,攈� �<�+�a���?�a��I��h�9��:1�3% {�Ov$L���v���2d��<@l&�)f2�����	_�2ME&���?�@�(����Z��DM��.!V�O�n��(4�v�뻙�ז��	���Ш�A���x㎥ Y�(7����w>L��*�� ���FKITX�ң�(dM��R<�)cr�� �$�����*�[@λ��uY�����G,���o�J!��A�ϫ"���	�������@/x��g�8�_�֥�GY G�����L�i��L��/.���!�YÞ��������Wx�tC�����"�|����ء��Bn��c�q/^��{�r����6��t	�x^��k�5:�����_���d��lxΠ�s,Ni�O����w�ۗ6\�n����?���� ����>vR�	�%O��%,����+&��Ǖٳ�G�Ȥ���X�oe�q�i����`�ܝ�1\��	��4�\����)e�>���b�vN������(���Up�F����hP$D��� ���ȗ�e�����/8��
8�R]��#Ā2ԝ�y.���v��["��l�[��wsh��[�F���;�@tV�ˈ�340� sZ�� �?�J�2�%�FS�=+��ve�X͜�a�u�F��T�T@D�l�Z��32p#��N�B�h�?U����G�G�����,�TN�6�T7�kW(ǉ�#cL[�[�Ko�sz8�p�60�B�v;��PǺو�-f�GC��Z��C��r�{�u�:����ԭ�v��D�sƕ-��2$*��X��n���~P����o$Mp�ƍl�-�-%:�GPwT:�" >�'�s��5�8j�H��^����[��k�(�����$��f�� �
����yF��B\�+~��ॐ�'�I��z���q����� !T x��qԐ�Q��K������q��^���4P�уEF�zw:�!��Y]��u��"$��a�'�=<���b%��[��u�
gv�e,�������)S��䝵Z����p�%�&�-���J/]#����PpZ��S�؃@���X!\��u�8SzZ焈Mf���fYDT�{���%�"1E�P]�o�y�&�^Y��ٹ�}A��t�P�v�C��Y
��w6L�QW� $!�H�Ğ�Ƥ�	bH�eoqz΅C�i��,>����oD�:��<����	x��d�z��8�.�L�5?ӽ�w�!)�(S�U�;�!ǧ�+�I�9��]�Pvq�;R�r-n�����[fdH��q��$�E�����|+��y[�Z�@�0����xk���b�1�{���ӼZ@�/Ke����Fu*�����O�k��{�:e�s�� �� cn�=M�ߵ�S��m�!�(4W��M�,�lJΥ�@��*�&��N���1T�����Z�n5?0m�%p.Э�m��^��4_��S��~ ?�S>�����X���w�O��K�Xh���#;�;f$�9�ȉ�Z�K����;�Bݓ|H�r4�ܨ3P�ʃ��8��>Ղ��FN����Pm����&S�PZVm�HM�N���]�U�4≳����:��,u��OL���W9���ө*q8�!/8�3���Sw^�jH@�1�B��)��]m��L\�10���3!@�_�\�ե�ޕq:��ؙo0�%-|hSY�Ӝ�(Qz�>�<:��s�'��ȸ:ِ2���j I��vt�4�\�y��1���=<[,&CӜ��2h5�*HMQ��>��c1�Z�-Am��j��4���6�$kiSR��B��kg�唍����ås;�rVs����^�/+]����1�YT.�k�h�NS���yj@+�E�U�οVs���i}D��w^�f��R�y�\@���[�YCs�'X�Q������tM����?A��Vj���mV̒;�V0��;�,��"�Aq�^f�ĉz���?��#( ���?�8B�p��C�6kZoJƬ>&-��9�[�qA:#8����'��"��N�QX�E����@�������8!�j=oeH�X�l��F�5���|m�q�T8Pb�5�ƨ
�f3o�:��mi�i�(�+��J�Y05��R�����c8;f��6'�V��jՉ[����U����߀��5�d�=�cw~@B��]���}�vN�#m>�M�T4��w���<�3�,�E>�z����Ձ��3�PX�Y�B���\�荸����Tz�AķǱ�ٖ�nP�K�o�����s�q[%�Fs@��=oV`�{0?����GY���@~��嵴^Bt�a�o�-��X�����\��#2�Vf�v`�G�Nr�LǸ��^EI�����ˀ}�����A׳��(*�X��t~����S��];�OPS���M���c$��c-�Q.� OLk��x��kF��U(ǋ0�T����)�.���k(m{���>��_s�,�i���[��K�h)�ozT���6l˓5C���k�ukr�� 7jr�q�3��I���-�%� *2�ۧM���O��� ��@ �?� �X�%Y�?=��ȚE�?E�6�$Q��Ys��*�[��N�~+�a�l��9��Ȥ�F�.�� L�S���<�\L���緊r?�Su���lk\l��.�9~Č�WL5c�/%U-���c/헼]�h@��sR���X��
�!�P���ظo:S����`�X���3��T�ޜ�rV>��9��AZr�kr�s� �Hi؉aP}��T�jE�:�"5S�&�xL�
v���I��$�s�T�Et�Ħ����%����10m��۠��r۳�P����i�v�#��B+�,�S���1b�D�A �Nbx�luk�1�~s]���SUA�����sR(�M��2@8��}q��b�+3b��+%W��l/(N�m[�P��T;HW��eV��MZ��q!�~m���}�t)N��2����-.�Q� ��*�S��J)6l�n3��"jU����s�T�����pRS�����[�۰eF��M �. �W�$�U��O�<��׏"õDaQ�6�Z��M���s�P��T�ˀ>��4u< �u�#�2��3�����ބ��zP�p�(�em>��њ��i�;l}�Aɀk����M��)�uc�?����D�ܞ��O4�ⷶ��s�,33Ch����g�a�q{n9FO�� �z]dM1��r[��|�H l�����;�<i�H���с�u-�r.Z�0��4M5�� �"T�L�i���)����2�#��V񑤝�ԓ4'ۉ��SA]�3oM�������,����A��h�Jyך�&�UjL4�8M�mi�R�2���n��pD����y�e�8��%s���|��`�FKi�~��p�9��j�>���U+?���{�N�j����8�_��+@��!0�@���+�@���F��2E�S�m��^4,�����EQ�����#l;������|Nè�u������:c��3	z����h��ڤ���ögvM!H ~5�P'țP��БkZ�6ٔ��8Nі�30P��8�Fn�Xf�,�ۚ�l����c��^�G\���RwQ(����X�y��{��X	���}GOb!�B� �g2��uM�`���5�2�d�;>��G��ϔKS��Mrl�BOp�7�ыԪ�@�x`Lzf����2*����Kd�����Wi�q�r�jν��O/X�/��g�A6���kc���������,�˦��dZK[MF�r��!�Yr�)�4rJ�|�zU�W�j&�RMq{0J�� L�AnF0I�×�g�6��S:j%v��̲�
�J�"b45)`Ȳ���%
�;�ZO�nAx���c��f�p"i�Y������ ���6{��t���u_'�_3�2�hV>�����4�\k�
�`-+�eqT�����YLo�P�|?ȶ������X�1|�HP��Z:�){	X�_MrFU�	+�m��3%ϭa�a��hU+��2I�r�f�_P�k?��5.E�@\���R��sd.Ѭ����1����o�&s�O,t�3US�i�,P]���U�#v�e�V�#�[�~X�4ȋmPfV|�R����U1���ށi��^hB��r?�A�!��~j�T�CuΎ��71Dsad��fp���ʤƜ���j�p��;�"sV>�uq�?����;�� Aؗo�F%��u�wJML^�A�^\�ڶ�2�!�s�5h�92dZ⇺Wzy#Bv��2&Z61]�3�^ ��s}N��@�N�#�d.�����e���X�n����=鹋�QZ���
.`�3��ת�sȤd�\U�;��&J�6�C���7h��as����'��g;����䂼�P��b�LD^�qA�P�l����iʂd�&�2$i�b8���v+�����Y�ʌ�I[��9����\緁����d�T����h�8�v���M��Z�"@��H��L�
:,Z��9k[��x�|	p���O*<��3G3��M� ��3 �C��͈x���4&��R��2�&�w���<�
,R$E��3,O�����3}=1��A��7��
X~>�H���+e�'�ޓ�E
9Ēռ8��%��pqd/�"�!h�_��n���T^�Rz��DM=����%T:1q򬄺�����J�@�N%�AS^F�3�$ڛ��N�ު���� ��aJp��b�/�9�����1L� �Z�/�H/E+�~�|�_���7��#L�;���F_z=�)��̪n6�"5�D^xk����}�G��27ʋP&�p#�)z����
SRE�̾�R6�$(�f��@~�t�k��\6W��h@�Q��:�y|�A.��dΉ;ЛV����N���Wy%�1��hr������i���-�g�6�X�(��$�.�bgd����h*�ݶ��SZ�M��\�Χ��Dx��0vp�9��`2�=�~��(̈́+�~_O6r/�;���t���4���Q"GTa=yL�05
.ş��jvj���D�x�&	��Z������4�f��7� X��F�ﰄ�ZT_t�oj8��^�E��z�ȋ[��r�G	�D��&Hv�;�1Xa��uޅu�9g!��]�s�g3waA�q����p}~%�*`��`y��b�\��F"C��_�����ᇠ �ll��\�~��G���O2�|.8\+�#�b٪0Y	e��eR��1#�W��ae��pY�$�!����4!i`���?3�僃��S���/P &�}b�
���
k�����Q�՚Չ��eJ���8\���u����#���d
|\�ǂ����h�-*gחHR+y���Jq��O'�|���w�T.�,����՗�1mz��~�V���/B���/������f���MP�����F�09 5^�_kQ?�u�<�?�8V�%�NcM-�pL
?^�#���k�R�6Ӓ&��H�#�A��jn����i���+2�V*ڮ JY�wY�*�������(�	�o�;/��y^��tCƋX�X�����Mc₶%��5�h�$na~'���m��W�j����K��dhFLX1ד5�d�
�5�x�$�T�kPO��<�l0�;���_��X#�:hc��H�R:��n��,%�gN�Yvm�LCE��s��#\��3Y�}c���KLg"�D_��ֱ�����9uW�W��fDO��S��%/��� ��������Z�a�oPO�H�
�C$aܬ7���?�Ll�ɶ��5�-ݚ�n5�����Js�@ZjmY���<ް|���P��z��D�aV"٢�~r��9�,��d���f%���_�%���$��u��k,�z���s� �y�N�
�L$�&��"�7Z�n�#�/��j.�g��"X.�A��J�*����s�Hֶ�X���.��`�a6���e<ykZ6���JZQ���>������c������O^qQx�h �-�3��p��]?.��ۈ6�w��%.I��t��M�J��"��e�]�_�e��x�pi����}���u����}K���'�ET\Y�C�����_\����}�"UQtW|s���,lK��>+ɬrp=�$�\�.���2E�͢7�%#�����K��ZC��2�3���C^���� �^��qwb�}S
�&:��ƗL��0�ʠH��V'1��E�p>92�J\�sÙ�+��V�^ϱs�X��O4������@���<����q S�y9���@7ʬ�y��8�l}���z�4��寕>6��\p��儣���$g�����G�'-��!��B�-�T�2�zZs�?,�$�%cp�1�5�����3����/,����clJ�%W��F�%D9���� ���/�f] T5����η�5�@%˘w��D�3�4�W8��\��]�����l�H��pKt�*k�{�y8+dZ+ov�Sd߯+D���8؅�V�S�P�߆�}��&O8�n�X����%�V�zO�j��&wM����lZ�fn@����Pt�wÙr�>�e5 �M���Ĭ�~�<_�X��+p���w��P˃�J�߽M�$�5���5�����2�6�\n��~�+���E#T=��6��(�u���g3|h�v�����cF��Egx���9��j��&�l������7��JK�Vp�n*��*����uY���xŊ%�	K�n�/8gW/�>��d#$9Z5 �@��|�p��3p/3�����=|�OD�(wx��u�X�M���v�L�������W�