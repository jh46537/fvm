��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���_���W=1����o �6!�z�O�]E���	Rߗ>���b�C���X�����>�F�P����y*�qGYjkҴ&�f�8��V��lzl�/
�Ĳ��S�L�J��pt�U8��5a�I]ҩ!��/Q��+��	�$�48�<1I����C�oV��\�+�i���y5���M�A�oU=aQ,�ӏj������x$Le׆ַ���ԕ���<%�1$������e��ʄ1�n��RՇ�[���"<D��h����[a>���{���m�i����<�<s���@��܈��#�S{��n�Ȓ��S�Ǧ�oc_i�rPiΗF�YN`�1K���2s�{��բ}��{�G��1���*O���5cU�E��yڎ8�倲��N6L�M/�H�ǹ���_V�#@M��ؗ.~������t��F�!F�#=[FR8x���Mgyv���31��5#ܴX��_����5I�-��r���g�À?
�5� ���2�n6����?}H�+.�r�&ElX���8������ ���D)Ĩ5�^�U���� L��7���fb��!�lt������ok\Fa���L÷�C�?N�A��(����"�ہ7a�Խm�ƻ2�����;RÓ��Cx���m�;�5���~|Hs=��P=w�,��d�M���#QుÆ��>S���ۥ@��G:{A�2�ؒ�n�\=���x0Q����i��~+'���ė��Sl�y&E�4\�o�Uf��2�
�d#E�d�݃�;�v�3�:K�nV��cKl?O�-����'OC��K�9/���ӡ���6 /������ݖհ'���I����jf给�:6V��T�R����'���۰%h�cP���O2y��gI�K�k'.gj?��ư��QC�����Q��K7�� ���Pk��=]r�ɀ� "O=�w�fi[�U��ֶ�X�Q��Z@N�g�\�E��	2�=� I��G�͡l����w5���U�����f5���6 ���&sC°�R8ڽli|��{�}wt�~Wi���`���IE���HHaA���eN�{ �W*��c0,X��{��'_����3���|c7��'���MP�Mj�$5�J3��7��F�'�Tм_�f�p������=�ecA�jq�E��>��e�dW�yn�Z��-�H�=��F��tN��`�(��{VQ��
�͎88-�;�/I�*Bׇ6=W�I��'gA�M�%�~��ㆤ~K�����A�Drt�������YR]��V5$h��>���R�͈�9X�j,�7�?L�-s8�Vrl�����N�g.)Fm<����/��?�+��X�3��u��5�\��c$�a�'��Z)�}*���O�,0�&g�-Mo��A>�\X۞�&3|�"X���<��D���(�s�w�q�Ʀ����`u�ZG,����痲9�M]�d$aNW�Z�E4wx���L��n���@Xwh� �<ٖ�5�n灛�}�8X_�6c�J�;L���Ϻ7#�-De���@�蹈0���������C̨2����Ї�wp�q�N��d{��B�����us�!�+�7�T)��z�D �4c�[d�º��]Hh������b���������'���7������1�à�|�å�>�bl��}��"K�q_�IJ��]�(bDlF��ѭ"t��7[l���h�P�Io���o	�