��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�c���G�J�,=N�{�P.�*�@�&��^[��Ԇ�Ă�#�a��� u!��;*ջ�2��n��:#7��l��8����k�D��"3rd+���]��*�a���7�a�W�Ce�L������ ��5u���#��)�g���=!5�g]4�y��t�/�Y��Kw"������u�J�M&
Rܾ�a=�;�D�.[9>��_2�j)���&��%O���b�R#([��%x�E��8[���i��xh Z�ulN�"m*��5ߡ��!���ʛ(k���=���&�}�n	�i��8�=�(=��>چ�����[��/��#�qĪ�7�������m�훓((IF�YZy�r�z}G,mJ��&���\�}ֲ�n��i���*u#R�c� �zP�Lr�U��]o���� J���Y�\�J��_ա叫�#�/��1��":0jO]�T�F~���?r�c$,����Ti�o^��f���eq�d��U[/���s������h~ߌ�o'�%v�j9���sY����2D� -�'%��Sn��x���}{<
��i���y�+N�i��.�w)B����&�`�ܜ�ۮdA��@���԰g�TF[ņ�Z�W�y��t�3�����jC��� �Ջ����4��S�/s�w�,��b��u�ƶ�>��ґtչ�J���F%��j���`���C�3	��@A�#��|���H�E̚n�s�ワ3.���lrӂ�|Q~�]��]�\!��F0�݁ʃ���Z5�;.Aw�� q���p� V�N#���m�R��6���~���R�t���[�0R�Z�aK&.�>����?f����!?��$:a'�/)�P�~w�@��z�G�g	9a�8�F�!Y����U6�<��#������ş�Y��Gٍ2-F0��eJ���XݓJ�a��dgT������� ��1�!z,�g�
�"��2��1�|�kOEV�TZ��e&S[��n�S��� �d@\�E�3����&w̜E����+^A�9,�)��������.T�^5N��8j��{:/����
�d^��U��N{�{��ҩ��I��Rǀ$Ɯ!�M�b!��~��
��Wy?�g�����[��)���lj]�.f�Q�������(AD"�d�*D5��v��rv��+����B���v��թ��� ��)���9�åCC�!��JfU�%�.1�`����nNf3�Ʉi�=���kH�� ���U��%`
e�R�} v�~Ǐ6��dq��wΤt���.υ���֣���gIM�B�r���I��|��]��0̾F����4r���>�������LS�.��@��NY\��`�Й7�"M��9 �+h�N�搭k2}nj��+�
�g?Ϳ=��mU1��ou����(R1IT����u��Y@)�jU��t$�-R�0��1�8�fv�S�m�4�k���pp�_R�,ܶ6��~JQ�cҭMN�3eL�^ހyHthV��v'��X�7@��M�Q]r5@�5�e�9c@���C������&�/^�	��^��S���`k����ü��{�Dx�z�z�f�y<���x����z7K�i9�Z�������Q"*f�I�^֫�����Ȑ����)0� �w�b�o5j/�b�߱S�9<"�y�1����� �@0E�k��#f~OfK{����&d��#8<�#-�ߘՃV�$�P�
ǵ+R�����X�T�"rY@����A������fN��~{�)t�QTr����M��#�k5��c��;�O˾�_3�	!-Qf*ݷ�	��n��yz����i��S����/ٟ��|�����c,�[��i�>�v����e����DϹ�_<��t�M}>y��*� wa��i �B�!-�ϐ2�h�n��^X�Q�b�frg�rn��扞�>��@yǺ[�$G�gl��srio�wy�x��'
қ6�z@O���Ȱ��}t@������?z�O��|���!b�S�
DM�{�i���=��&���#�#�p_���"��-�"yS��K"�I
ӶhG��R� �cn�3W�������������8������^�$I��rs�5���H��n�yq��oQh�����O^V�|��D��],�Z!�	�͟J�*(�qˡR'��r܎�!�cie�HkԒ�|��[�u�Mת1%m}�����h��gmH�~˟h�7���a5�Oq\��lan��r�WE?���w�r�Igk̇������xy܋�M���s �<�`,� ��S��(�I�/4�F�gbB@�m�q�t��7!
�<���v,j�7ݖ�W��M�0���T9_u۪:���AD��AF�J�_H ������0�At�ߤY<;v�T� �ʘE\�O<�rO�HYnD�
��RIh���Y�.�oa�NF��h'y��X�t�-�_K;��h��4���~y��WF,M�TR�M�P��1�7u	B&uo������Rf4\;��Ưm&���DN?^L�{ŗn�G\s�g�0>8�E"�y����_#�z��)�"���&��1sSh̦u�����"��Y�{�<�~���$��AE���p[,�~�͍��v�sG9L�z*���'�s�nyh�M�7d��h-;��ݧ��$��d~V �<7M�� �]�E�v�p0Θ�;�`������S,0�����V�(��ÇZ��d6��\R,�M�C�r�(#ص�љ<|W�x�3��#�>	�yL�Skd'ٌ�5�@/R���5%�\2�\j�ЄTQt�)��@|]�z����=���A���%[�eU�ĥ���K-m�o�����E�ܰ�_�p};sfRV&���9�;�%�tŰ-<툘�0s�&��p�Î��u����	�
�_���h�K�}��m8��4��K8�>;��b���^�%��'M�xH���CGR�;�D��Ճz w�h�~F����~B�+��4ܳ�V�`�kEm���'�'�=Dl��i/5Pk��$���h�~�y�t8���Cߋ�{!��'�����Ѣ��� Zyc������h:�˃)C�S�gss��-�+��cm侃/0繥K���HQV�p�v>\�~I}m�\`{K�Ա���F'y��.\�/�Ҥ����o湃&a`��(KCŚó�TX5e�)z�� ��$�G��Ɲ�U�����ؙ�m��7�����Smk�u$t�Y�64�~ق�b�9X�O�V�w�Qi��8ǎ5�k.]Év����rL;&��Mg?�*-�,%�6�z���e�1]���	sO�	���Y&@�0�$L�cW�l�5��cb"z�!Ѿƴ�x�rϘ�4ǐz�F��	��P�&�u�
#8�I�U���4�����䮏�(���ܭAU ޏ�ޜf	�oo{�rd ���FM\A�Q`��ÚW~�n�N��NY������w�oV�Jp��w������t��;B3��V�z�ا<�ȆPZj���ꨩ�?)��3Z [f���'я���S��h���e�M����׻ev[���U��O�c��C���t$�A(��-i-�~]!y�>i4��'�,�mCØ�G��2@&%y�q�b����'A�愉�M��'�(� c��M[��xBC��T#�1�q/�*>Z(_<DUy��ف�&eQ3��gx������$IC�٧n�^��Xq,�F��9G$d��o"����#�J�R[�-�*�]'���q�ap���7�)�n"МH�b�^��4:$[ȅ�i����ilc�2wm	�:T���9��S5�Z�?I7��LƗ�)˦���l}�|�;>�A�be����Ʀ�P���3�I1���fV�������N	��<
w�=�-0����2�݊�������:�O��;��&��i�Sd��	C����y�^]I�.=�xU�m�
�8���D���pU�q��LBckS�|9l��uԱ��B�f��ǆ�g�/+ '8��8+vƎ��ᓙg�k�b*`u���F�W���
��Lͩ�2�l8ݿ��ۑ���{z�\���0�(]�d\�192��ej4��j������}�II��^����m"�Q��e��>д��{L��}Al�!�ݸ�Pd��7��&Ea�+�"٧$����+�|��&%~�;;Գ� ~Z��9����d_�'�q�������S�S7גi���Z�h1��}U)c)��	�hn����O!��*
Rb�z�L��z�0}iv]:e)׬�PZ����;�e����hz;t�u�k�� W'�Ĵ��Lbr�$����:�%�*�+x�ݰ���7߲�X�	�x�H�����G�a���
.���U$��u?.�KV�������*�I��y�	F@�Em��XPV��qy�>��p����>�M�7�XK�"4q���nuH�ե�"+�
�Wq��3~+k�������5�a��aS [���b}��iꬖ�\y����@���ڜQ��� F�Ws�.����lI��%L� ����$���3e"e1\(��:b�P�DdM�R0[iT5��N?��`jSƋ�Hm
8U����`����$u�(Aq�����X\GV4>����/�F�5V�b�p�ዘ|�8���� ��s��B�0���7s����ބk|NЇ��g�c�Ė��qό��Ձv;ԠI�>�	On���b�'��#u�i�l  yY���v\)�A��>e#���cA���x�n�̥��%ul~�2�f��J���D�C9ʂ���N�@9	�R�y�+���*0@g��#%ޖ�U	x���j�c�X����"-�vo=u�����o���kN��SRi֯��Y���Ӟ��W��è�z���
p��i��}.�#z6�2�u�c��L9����`�P��&���t�w��;�8;(KIeW�kX��B��19���NYxw�QkLC��\o����4<��[�b���M��;�n�������������}0T�r�u�`.�d "��b`sC7 Ah�̣|~�C.׽�4�SF��{ '��,���f2�dD��Ǯ�O�|�H@�&��`��j���	�txb�劯01X{�t<����� *y�>V(�&?!��S�ub�LΈ��yV��׮Li��!XV��d7��{wMy����r��|��W6�Ն��C��.|~����r9��E�5P����" ��t�bW��]���H{�����x�zZ��rr�6� [��G���;��D��{]g]��s��<k2�Sv6+�2)�'~��1�9~��>��+��x{	��n<��az�u�b1��� n;u�}eA���}V4��'xm���C`bP�����9w��E)ٟ�>��m��Q��_8J򻘳!G��z�����̥��{Z�1�v=�ht��Te
}k��Q|삑k����́=�O�����56]�N	�O�V�k\�o󬶸��Y|�w'�B�٧ڋ�!+﫱1��(��S�����cv$��4��������-EK�HW��Mo5��x'T�k�w��md�Aa��irfL��n+�_��P6T�A�8���eA1�0�D�|� .�	��1��R��"�'p�*X� �Ի(�[K�>�o�ky�O�́lY̮���\��j6"�Dzx�Mq�.��� �pu����;Y����'(���2d1<�b������?��:���X���Ҟ�p_�?�5�m܏�K�;�����A8V�%��A�w���Q�֠���ћYGg����lH&�9�s	v��ԃ���å�똜�bZ�������덺O(�We��Q��屧5 $��U��i��/r��>La~���Ic�ī�ܪ��-�3�p�R=����ϫ0Y���OT��O��1�o	��՗�L�@��I���� ���ؙ�|�EչZ*��Ո�� �e)Ҁ��Q4���&q���������G��U���1��.j-�R���w�1B*U�$��l��
��)�����-iG�n�v�H�}�L](�}�(r�7���+��j�"��_t�� ���䮆�I�j��f��C��Ir���$p49K��o�-aĆg��&i:�
A�W٣��o�	"���nj�Ԓ�[���ȤDV�	��f�J?���j|7ʳk6 �|k��;![�Ůtq�:b�S��g���3a����Yy�&�ܳ�S�B��<f�b��S85UX�8/K?RVS��+�S,(�F(��ݪ\S�*!`��}\]�j�(����X,Mn���[�i{���'v�&RJ����Yn�8��h�p!]��T�"�"��+uzC�Jc$��Z��a��|�d�8?���?�P�K��xF�GX�R��4RCnP�*�;@��z_�DE~�xu���4P7$�l�U��{��f�t�e�2�_дQ��ĻKf��Q�2v�U&�)�����-�Q~<i+����\��qֱ����
p0ᤳ�,>�HS�F�&&���@��%8�e�8fHC�a������<�?�+0�'x����@ꔫn�$ʃ�(����