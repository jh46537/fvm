��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}�����°ȣV��Ak$h�٠��i����(�Yv|Y]'�;|]�#���tA�.a�\D��\��4�MW���뵝w������9�[�ko��6u��T6��O�T㖑5+`J��^��:<��!�#���c@IшGg��Z)��5o�ҁ�	2�	�����\��}���Eo[���=�v(k
03�T0�7V�t@p뎚�*(*4<��pJ���kK������˪a�w��������W�%����U���� � ֟uE�_�5*���@����<	�#r�� [xݸ��bbܧ�2e��j�B$K�����o[���o�y�K�\�
o�oy_�t��)Ϻ��]َ1��N;��
�Ad�.�|m�@�9i5s
Qv5IF�Z��앍l6(�����_�б5��_t$�)Q�b��s9��n&�%��DQ��k�y�j�����hRV������U{�O5�k�ݹl� [�������!y�i�5�"&�����c8^Ck�J:�v��F-�ؽg��W.�q�������Α�AqK�c;�H��s4��ز���}~D�!��+����Iz���[)��};�#�}����YV�!�������)h.��|���
�Zol�[;�r+y��	_~R��R� g"�u��sF̳W�����c���ކ6�<n8�XYR�
�����i�o��<�x! [�=⏰ϔ?r���2lOuzt��.�t���r�7DR������m�A^loP�8p:W�+�t����K����&
��8�[؍L���R
v�4�-�i�yF@�N�C������#��̌q�|/�J���)��?'ӛ Mo��S.D��ߜ����b)Klix�lrL�L��c�y���L�%iR�h2���3��X"��ϣ���X�Ǿ4SKQm��r(�~���PiH�圇���+|�݂���G���
���෢}i$/�׀�@�x��1@r��SU�8�c+Br��υ���e�rot�X����� 4�S;=0��UJvŞ���,�su>-
g����Ż�j�y���.��:���θ���<�(;\ŏN�\�-�����zPR�\��`2��^s����2[rV�G��趧C��$r9�w��[M��?
�$����(�(���Ŧ{m���eL��%=n�6HY�W��`�'h�J�3���xlJ��I�`�O�����@�O�[P��5�ђ�/��ӹ�E��M,��������n(g�L"�W�;�PxsY������]?�%�����t@�>Gjh��藞��\��uǆ���.�@�0H�>*�������x��ߓ�%�[����$�3���@�h��7{K*�����!�q�c���a,��_9q��7JV��R'd,gu\Ǳ�zY�Щ�8T��1��=V��N�n�ݚE�.�k,��Y8�$1&%��6���`��d�ъB�Hn&��n�����<g�h�#*�w4l$�!�+Vy�"KÃf�Q$m���9��`�tڧ�Ro6ʘ(�T�U3��QL5�5��(�V*D۠K_ҵ�f���ֲ@0ʶ��r_����xq�+�1\� �~� Ͻ��«V7�_��z^I͘�s�b��b/@"���6�+k�w_��`��G�ȴ��65�Y�a�����eY�a�l���ߥ�l^7S�?+�Ѭ�KUeB)�Z}��b����?𘺄Đp���\W��v�X]��y��L���L�Mk� [bx����qkO�Ł`k��D�~m���"WzW4�Ԝ��m�ĔYu��	�p �Z�TV\���E��`�3�Gĸ8mK}}�z�����\��i΁����N�S��! s��p5"R�p�h!v`� Q�b�����G*hS:��5{�p�l�kA���X�C�*<�Jg:��<��.G���b"���?F%ҟ���hJ
v��8��U״�?�X`�)�*X��PB�v��T#�42a&�|l��wf��f 6Y'��$y���(Z�c���N�.��	%���o� �$H��IQ��q��kB�OT�_W�^Q�Ⱦ�?O(� !_��
�_�䆪}�^�*1q���k<�q��t% p�s��+>c+�UZ�����￳ŎQ�)��U"iC�*��]5d�!���ې��}>�L|g�]�1��T���z��yR@�SN=�xD�'��� v��8��[��ѝ�?ú:&�C�Y&P�����L�_�xf�
� ��op���3���_��6����� �Li	`�����X���r�U�W���H*s�Su6*�*��Q��f��9?�����u�E��m	&uXV:�{�)�sA�
X���(�&��5�rb^<���W��8�s�w��>{�fj���AZW2	��\!�8�05p�� ���L�h�Vzj����~�P��u�\g �9c5F^��˫F��D%���s�x�Лo⍰q44�LVm�`���*{t��! ��rf+�.�#��&W���sakM���U,��+�'�=�������,լ]�(o���Lbhy�����N�X��m��:TNY��h���B�R�@E:�?P~�^ˎj�p?���v���t���z�AM�8����e�+bٽ���ü�7m��EG
��[�B�^��)8���RQИ!��h�������p��w�Nbn�,E�lU�#�Mc�)Ȍ��e�q�k�����H�$c"��,.%[x	�]��,�Y���3���7��[��__+�i��ڞ�	��'rk��b��K��T{(�W�9��1%�t��dű���)��&S�;.d~�O�<�6�-Bp?@� �z���/��yiru�a�@C^��g�&���¼:��<���Za25��Mb7�Nl�,��!{�MZ�����F�n�)~�r3?�����	��:p��^���'=���p�q�@�M�Eʍ��!h~+i>�@Ҏ�� t-���m�__jW��f��$�������^#�V���gxǩnh�X��P۳]RL���r�������ͧI7#>�2�OE���y�C����l�$�����W|�å:J_�yGG6s����	�<(�d$��-���n)���4���*R��ek�a���t ׯ��ͱ���`�^���2;t|u�í �YQ�F��F�!m��:Nd}M��3��	����Ԭڳ��8|��r��6M&�E��d�H��AN���C�lw'�!�5�b�ْ��`�x*�{�H �Y�Z�H$�ͧ�[� ttt��R������`�*	�	C1˨=�ٺ��!G�3k�I�e�; ��`��/�r��n2+8@S9�����:�H�C�Ϲ��w����Tx8�1�����g��V8��} �Ƞ,�s�6�%
2v'�؂�Z=������ʓv��V��n����.�WD6e�&��������^�gE�\���{>o��!�vIܹ�n�V���y��<;���;��(N��qP��&'��)�5�U#݋Ј��0ET��΂]T��O���rd�R��6W�/�����=�A/�if;=?�r�y�U{Cp���*X4��+&�2E!id�S�Dn��}��P_���'@b��S����Tux TIN~���rRr��]��ف��RT��I:�cEK��Ԟ����7�\��#n�
�TT5Z7�O��W�x�����H�#����1�"^
��l�Ynf�T����z��1�0簚�şsc�|C#��W)�Bω����M=�^�rǝ���}>|�/�&�&��T����8B�'�}#��*`:���ݪduh<���z5M{˴Y�9A*��7�^ͨsر�S�U�W����ۛs�V���8I���L��ze��]%�<����>��[���k����ۣz�a�+�K+���1k����!�9:k��t��DwX�.%S��7��S���
��&nK���.��7z��G\�:���;�AK���A����_K$$��@��K���r�-�ķ��+�-j�c��'��n/e\�F,y�X��aA��%W�{��H��W;��/&% Ƴ9pm�G=z��4B�w41V8���8e��B�;�x�Ďv�x37
�f���Tf�Hn�]+��(�E�����Ϩ�$�s{�aog|��Hڄ��X
�؞�fOy{w�vLb�s��3<�>�L^�K�v�C稻_3�`�*��������&�t�x�u{�Y�F�'m�eh؁<1�� UR.c��7��yWp�1�ʫC<�b[[+�H]�e!+�r�c�cl�E�Zƒ�k�����߰����l)�D;_m�]V)N��6<�#�Q�"�T�?~Y�;4�e��/���	�����>'-E�[�Sb)�m�\Srԧ
�h�ʯ!�x�ޝj_�F݉6�r�[��1t������@G��02�_!o5�'+Z	to�E���ZCn޽�MjnG;�Ȫ���-G�S����GU�K' {�Q��#�}	���%��yop���2~]���㨋2�^�-75<�����ε����%�ca�I���uS�~N�=+� ��:� �o���`I@"c����/o	&�6�R@.�u�|q
)H��vh쓃ߺ�S��dŮ�w��J��7���#%'�۲r��tP��H�Yj/�}�*��|l���,�I�I�H�:�	��)��c4�}�%��Gel%��;lI��w?${9��Q!���׶�?3���n09sL;*8� �/�A�Dd���S<�^���tY���^`2 �H?��L5|�A�g`,;��LK��-�%�-�v��C@G������a�����'u�o8�ދL�O�|��:�k%��0aM�e̝f��ʻu<Ԯk_6o�����+�~εg��N��|�6���lh�@��=`d�vs�{Dt�9v��감z=v��Eg/��Cm~��ط� ��Q0/6Ko���P�E��g��h�V}��7Ͼ�V��_(��g��J;�s�g�a��~�%W�^��7�ʪ� $2���3���b��sG�&Xh_��g��MR+$�3.����6ަ�I������_���Ji&�hF6�T6�[j�qi0Y�rx �}�U����H����m;�6�s������+9�r�sI��K����U^��`�q����S��O��H�n%��%ҦAa|��7�4!�{өźo�K[��:��������