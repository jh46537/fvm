// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:52 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YGrbJeOmYD8+v4M2SqvuONO5BecN6hwUABUpzD5Gy0Yza9Xb5N5QeGSnhx5CeaYT
KZZcGmOe4Ci6t8nno3/9TqW/M/IX+nbiw/0gVqitxU2egJX2lFge1N7wW18XX898
d4WWXe9oX++MrrmjPJ5oZSQDS9L8eyIcdgU3ihLxa5I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5392)
Fu0j+h0ePlvGEoKrICsYtgHp8xs+7cV50m9G2Q4IAnRqt6voB4TwPcbRV91xdBTp
S0n4030RqbpSXtsimE1jXJS+x8cIR5d3ejtPrBwgTDUUoctAxPijM4Nfl0pshXnB
5FpOLhFow7P6dtjIET6KRQ+ztS9zsdoHUMEXRDxhaWKyNbvqWbnfqOydJxIudVrX
W9pcQ9xk8C6tPgHTbCr6i137nd+Ltx2jr84+Jp8cVViCA+txIR/rOHXK0KUcsEqQ
WtWpueMEApFaiJ/O5A1AIYX/3wlGOAx8vYHgoHy+dYaZgntEz9htMcGAdghRKyzM
nOEq4z/XrzCEgAhSqlKeyXtK1WyvsGybX4475hPqURA63lbg+rQcAGYvucECdAB7
rHxN1NPVd2NBdProTEsBgZMWE2dvtnlTdMGv20ALS2jP8phmM0y0lc0u10PzEZSH
WhKqtLgk5HLJvtJec8kl86615tq9rv9P+q3GTg8HjM2iGIihhntja82L6fLAqrJF
dZncKASPVCqPjJ905E7hLJAt7v9/PAH1HCkYZcAVm38MaI13iV95bqS0tH4EP9+5
xgAjth3qYdLQ2xBLzlO0he2p+H9SCx+G7SJXSuNMUiCz5Ip9+s2MSf9x7FWLHDwu
faTVFIYf1qASubAcIttP4kHp39aJBdR0JJudhy0yFyqQHeehXxjtGPOQ1OvUWsRL
51zpyNVK3JByg6DW+TC0YY3XRiTMNiNZwwzAmjJt4/3pPvIQ9AD+jZpiX7uGqVNA
0b+6IbhYROULqh6NKyCNs0t5CGCQ0bVB7Zz9oHpCpU51a98uQ68TEb6roQULBv9K
F7K3cjkkuWOiz5GU6swzmBRhR2sg/FdHJEkh5nLb62/9jNAa3nbhA4GY93Nq2aw/
r27cxCAUr70t0XmV945docG3AZWdaJ/scjC82yNDMoJa8TX3ziuSqzGtYmFtQjkg
+Qe+323b+gP3dpS4kaj5+RzjxkRhb+iunPjWX05HG7p0v+aUfY+fu41WP9Bui9ri
AA6QBihjr86NnMkmKHbjk31Tl+gkUozhgZoBvK2GRkPj5thZDXsVlhC+/ULed8iw
For8VEZhLKEjrsognffE23zXq4j4CKpd2B5Vvb5uIOyFLW63ZPNo1sIxJw9RLC8y
rrCsdXG1PYhUCD6D93yrBCgMVsuQgHnrnPebVWBVbjzSVb0w91UVoqYmJdy9DBUV
G74mrtT6cotDPpqMBPmAeND9hAonwVdRnT9fC6mhZ9fg8M2teMzlxQhDLw0flvyr
hZ+4sF8A6PZrUiiEsQ1wR3csLyma5HDwWMRga26CNryPZlIdg0heQqU/ujmQ67J0
8nX+6W87otXuc0ZeXN0VJiaLWbwuCBWwnbXmvX5RWCO8gVmf3f2bren6b5J/SDex
Ihv2DWwWYWyPIEIs4ZbEZR+2PeXfHXjUC5fjq9NXI2Jq7kfOp8zsiV3mfnvROWVd
gjTx37Lq3MdpS0UNgSJX56OvGNA4IvL3K+msxsbaFHYS0mPuj44LG0i2Mua/mY3p
F3Ks6bCvNhDT5uG16YugWrX8GCY+2EvI0ZFKzybv0rJv0Kfd2lQZBgcHPRx0Z9F2
9hKFRSFPi/WIilCiLu/8/VRjD0xieKkYyS5vGnpCtLAe9Fu7KHiNE+ZQzTMAAGjB
Y4FOks/sGRfPCHo9UT4s1pwxPpgMNMmPEOIYwIy1qs3xLyF92d+to6AZCLybLc9Y
jF5OT40xvNXxgxk7N+ipzWzEnziWcYOJCuLBEOZ9boG4fAL54i+nYGiGTcAMF12V
mCgeAVr3M5QiOyzFtTMyHtgoDjkB9eb179QRx05anTlEt2ol5t0v1zjdcA+GdlRl
H4E9mj9bTZ0gpfYYZ9jFHCjabN/F/S3W1/cn/b32Ft9XrjQhHfiQ27KEWMSv6hjv
EqmLycmz8P+eppMMkFTX6SU9vHf5bljLpoiQFPWEg04NkpuT3zvuN82yQsu+1nFS
6BjKE+23RBEaUWRbFy0F6SKc5tU6Pi0YZYeM6wLCaKzIRAHi4LDtchm24NK3fDlq
ePoCvsSXJp8dM6C4H0bvJeuHl7WTlGm08iawVSHZ57ILcj9xBMlvsWwMmiCwY36g
ILjNjVtJk+MOEGimz2dQSLneFEubE9mavN421c43ztQYIqPeJkMjWyHIUNnUZ4S8
hhWAfXYcRNeWCs3sRkSzTwWWXFmwWOePLxkLAfe6Gakfbf1YWcF3Qwam8xY1khQP
RiK5sCf5C/GMns4MTHLuqeb3TrJncPc+DGDVq4VuOY4VPAzs0i19wjs0gm/NVjzS
zjs2GYH0zdIFM19jtLVkwY9UOzBKoSmoM+HcRHny8bN5oSK8SyxI7ddeKGCu3pPq
zrhrIGXDtxIIZQTHrD8VKZGcpvTGgvj+0VWrFeTMZk8ZvVxCEQX08ffwOUfcCRmX
yrTUZauMzIdLku6eOHQvxFeCmVq8qf9h8GmNXNoVyUQi0+eEEtXV1xCZGfPSx8iu
7UA6TzyTf/ccSQp2yITG3OjSGgp4ICukw9IBNV6rgihFLlHmxxSKmOjlNiMfxKFO
7BgNF0Kc047qe7vxV7tG621u52gocwjxk6rtEkxYdBaTLsDyOJajaz1xte7r0c4H
sJmbHR5QF+dKC7BK8f7cfSAd3JS4k+8HQl9bxvv+F6A7KHw1kmV8CIUzOnzOzKE3
nJe1d9jLOHO2SPDJiS1DyRA8p8O5px6vYSa0EaZAQnwWbRlXAV3GYZOqxsW+99f2
y4r5T/cC4uC2Y3/mat8k7HqaZcSGNLj/ndlQxBEb6xB4QtITM42EJBU+9Y/vseyg
koj9BSu3NRgC7Zcm6kTcBxqhqY0cCp0+W+xbTTgYM1U3NCTET5Q8Ut/AQ47YqmEf
BKkpcztlVhICpUED9VNaW8nreIh7HJmJmosjN0A2HDhIITdupNcJTR5Lz2ljcHkX
O1JfKvJsxbF/4jDERIpkgsjBpkCs0bk5/aANhi4cVCX3vjBrSXgE6rvZhxzQJmQ8
iBVT4wlUQ88bVF0aBGhhgBeOiHF9A//u1XcVji4IbEWm1qoewExvvf+mcKeDpz5a
lL3HZf00w6aY+Dkwlxl/fXf9KwJwaZh3Kckq0FvK06MCRcfutPmZHk3KGMCfWgCL
Al9L9qlcVZEA1Lg6DXFgTHjXkyiBFTqgWMiJD15rvDiHt9424dvIxlV/QhgcTcFF
eA/rVrarxcjNjkSLk3eHXRcF5pFNblBlAb+6M36yUkaZBI48Zxi5Py8FCIY53jT7
IKKJJN15iiKWOnzizlcAONLtmrsEJf0wqaZpxPhbwFLL8IDu1lYCHd6lRqQKE3xV
V9JPhpM1R0+D9ywnBIGihLIizbiqDE4UfrJ8SfCUoVRqIOuxcbVk9jqwNGIIMyf9
B5AQRbUZvFm1bJi4tVAAduiyy5OsuITFyOrX3BjqREyTc21fRvYTL39tZXMpEzvl
ABdrunOxKvNv4fswom0yk5RjPurBKgiGcNyszwmAQVWB0OllCL/IRd5PSg/mKMNe
wDdlNJPXdkde++Uru1JljtdSb2eiwknqh0m6kfwjgSY3JopP3vQjZzRfqg9C439A
sTFWwYrEDp6eP8wzFrI79y9U49HL/DisjLhou8UM0rOdyPJYehMZo0EwcpSHVY8n
OEFCF/7VCNr+WREhCtBovZCnuDXUyOYCLV4oN1voNXJi7NEMv9NWJSwrboAVKRDv
hjrmlHL50hExJ0ZJCt3ry47JGmtP2lmZtYz+EhgWlxaDTuMzPkPy2XLT07iacfHo
inozErcOoHHAlzkqw4kehnp8JtlkKhVa2xGjA3Jf2OZR0gSJuda0yxkCAg+Gikg+
ZqjuO+uKiMjSxrTeha23xXKkghcQMVdTIfBtBj2z43NCcihNDKUtSN0D+nPZcCnX
OWFvkytAzPiH9fLK/GpFRTsIgZCpQlAjznU224bUdq7rjpb01aycDVdOIGrOhQmF
2lAG0ZTLnkSx6T5lcf9obCto7YuTfKMHxsfCjFxR+9n6ilm28f5Hwf8ZZ8vMyzur
kX/b8K9+YZ1u0D866bEI18/x6bOdriTCoLNvpieTD8IIyce+x70Yh87cVmpST3af
9LjOK4AppCNMPYtQ6p+KY2Pu4G0Lvzdz5UT9FBfwrSsd+A3ZKzPH5nAf165dbu8F
xw4IwkYRAfl93JIaApEGmJRy92KNlmA0optM9SqgChwVmslHqIWiNPp8p2zFWqK1
BeebODF2an2gVtVAFlf9z3ptcx/6XeHESZu/UOpW1HX+NmYLFMhgxOJoVWZpvxWb
bzapxrE8H2ztbV3LM1jAnv8kfPijodXBV38e6GnWoo30mqSjxYr5GlKbejDJU0Jz
KtbMiWlTrJBHYyEPL5Ba9OzK+x8y5BIvf2zYLEYTh8cKBLpM9UNwHiatuwJUGP7h
aBS404EYwNGe98pusdi/k3l6rhJFEZ6GC+zyJR8LK3ZRWalYUI4BRZiM7BTAL3BL
S6ayjKNMr2cvJe1t0bbMdmDdUav+DXHTeiX/Q3Bno0OXdDNqFbg9S+qVU3Hh5ibc
QIAvLGhmsK7a9g3cK40nUDrEAkvMFuYhJb1mWGOlz0r/47zWaCqGM80S3e91JVZY
wXLK7QUPGv7CHbzXxE/5ZiP2xIwgs4R8IIadaeCo1yQQneYdWldH3yR2GIOCd+2u
GdKZfyE0k+gkAd8SiHwsGm1JpvKSv2LO6k7AxXaOLCHr2qbY6aL1g6U7zH12Vvjj
K8+hyc+79HKv7CZj6dVCq5OhBga5B/XCwPSuvmydxIl60zlpXk0BKmggGN60iqQ3
nWTrZN8DJtUpM76NUJfpnuxFdBRov4XaUSqClMhjJRVKmL3phyXIVGXyB/Y7LWht
WwGyM+FGsjR2nykq43lTZ/U54+vGYDD+yJWOMcFg5pjnLjLsKbJn4Hx1iE+cWym+
BbMhUaui00Vc6DdbqjguvQX1wZKZ5dXqOEvdegU2Uw2cn15UnLcM97XWUnn6xJEe
noqWgtxGs8MwuwYscqHiFIdpCYk6GqIDsV0RiG+wXX0g3Km5ugIvPDW2BtASy5hk
cpRuq+73ieOiXBZwF2YVyK8XM0IU7swpzpXgmnDl2niNAPrXUrqJpNMnxtsGkV94
2j77AneNk6v3ZX7HXHcPmbqLre8OZj/y/69VYhWjSyw8Zya+SbEh51JbvNG/I32x
XtPLf9RBi5hrUq+ioyjEPdp8MJUKhHAoRJG0AbzinaIjk0WyxwvNHiySI0CvttyN
UkeRIvV75r4LW1sUjORkX4HduE/6eKAigWrbemlrUumzOzYbByA9U4OAN41TlQJu
mrUjOOK7h2Dzfi4c5Vd4v0leffsowll9mBVyKXPq1pdzKaI/8uEauwBcxjR6nX2g
2JdoNWHPOVZT5xB8yUzp1iqOg2LEsiIv1CA1NLyqgen/z3aVeLgCrLJUp1JFDMIS
DOAPXTLtmsLP3PLG2ENfZX8t5oSSCwX9xuToCb807ZFtWoGcFRLMpE0VniHNDLBF
JPPuku/R/Yeyno8HShjyzh/NwHt+7kCBr8irGX6XzYh31ZDUJMHBtDbateIsuIRi
Wg97Q7TzrbmTCpCgWhQh6JccbEdJgqQsFkzMiJ1dZObtm2NeNnva/ZqQsfyVdIjL
VjtwfapT5mrxEsgiv/iQaGDCj5gHg31iepigWUulbnjODmV8TPLQDFpXEEm+xDLT
KR5J4VY7LkEAu/q6NBGlIujxVbzoqpxg/jexkzEdSrKPS8J0jZF+y6o3mNbsnbU+
rUmRfsaVwpdJyWFiWxJ3vu0XfQ/cZVuKvuZ0/tcF9Hyo4AZ7bPTUnqe2ba954uNw
6SNlqZjTPKGcYHB7Q/sDSAKOQ5YNS0WSnJR1ZQvtZlOFxK7vqMfTfz4Y30xg8/Qc
Fg9LNdOway4EYP2qXVdYk60FwjwKhe06CiGKyI7N2NvNbewssRFdwM9Wo5AhSiE4
5kVP6Emht1mqLrDTcw6tIEB1Rxx8i/xAiwege+PiSdIE1+VQkxi2ueT99QzGCB8d
uyAir+TXO39kISZkFV4z0+aQ9tqPtP2dXs9tEA2SV0rWn2QH5fCZJK9LOBqTjK+L
QEWZF+M51OjEYdIm+7XZHGyW2mwTXTduh3IOuSH/5nqiQMHVKZjP8J3TYt8bZSQJ
n89sCtSvpyv63JmPkLW8xh+7PKL3f581tmprr9nM2L2iYoLjIZkBlO0+ob6w4Uqn
bTWpz3yhW/vzDx2oDZt9vwZSVeaK0pDU3DCQgD/ew8sfJ7M2tLM/p3f1ZgHABHS1
fX9rWzzF+lTp31OjV7gRswuyY2cxxCVjRFbGdfw3bsrW7AAsjY7HM5+v9wrlaNOe
2ttK6TBigy1w51sX9u878dR6JBSpOkGkVxlXA+Kb77twGwZFhBz1BDsU9GUlcaWK
uDFbTkQv5DD8Z/mbjYTzhV+JoSAsFZwvLlsGPx3PskhhhNyAdmhidNHREZ7kACEh
NhJq7uHY2ftD97qoxTM+b2M2Z/UxeK4+828m4MTBnUbv7l0w/HTS/Y04RN0L/dp8
rCa59NMVOfPRUfNKw6/OBkNE7xFRRbh91GOwph/dhdaK9abvs4z3kPNx4TEyYtoV
i3Aqyv9wU+VHcgGQ/XzOLBJL8DZaSgVg4EXPIeJcj5pUNSfAEf9XEI5KtPz9+M8A
OybMLaYwGOCC3jGVg2NBqMg5nemVUjimdiamTPaY2g96R2E8F2Kwsnl1ZwWhb/u7
TSaI3M/LbTjjFh73F7y9qGlch8k3QTqeZKXiZrSfizVqeSzOzA71Op/KrN4J0UFc
SYjaSOw+q4r6MjD8dgffTikTJRwrj/LMBXVbfNZIgbSnCJXCoCDr0IRHbqFN+NWk
HS2exLLLEx9U++QgsorixMrBbFY+AjWaB8cVd1F4qipOGIp30WcXyBwxa0x4ObMW
VsV/TRkGDINM0ffNq+ybEJtzOuir94bsTHlWN6i4GqC1wjmTjwRHx226PjuwblLU
89KecHkV9LK+IPN3oc+f/AzPGD66GfWJOIv6tuCBleggchjCW2VCJZAa1HF5auZo
BFgirJ8YZNE8B3pGVicHg8jeY3YL73f+ZrOnjhqxD/mTbHRISlHBzqaiHBGHcjH2
TUREBzVf/QZrEI4SCOmgdVbkLqZVB2fF5EcUqpUe3pwhsaU/WZmAHzUpGETN8X1r
650Xh2O6uJUVN0u/rgWJDg==
`pragma protect end_protected
