��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k{de���ӱ��.�|�2#{��Z�V��Iu~�K7�ޱLC|X���W��mJ&j!�Ӏh�d6�T��5��O-��0U
�R90+����B[A��<q�z��U�3��j�m_9g,�}7%Qc:v�����U�Ug�[	V��ߴ�7��<�.��G9]�Dپ�V�}LD�#T��a��,;:�u#`�r󉛼x�Nw���Bd��.�X��������C�
 nF%��
%^yc:�3�ʌ�C�qt�6J\0
��K�Wqc�ɩ�'���`��u�Q�݂�ԯ��������i\tP�p�A���}��t�1f%�<5;Sn�[B�q/�\ݢ����й��f�L� /Smss��0���.Cd�$ߠj�ToWoPVx���X��ц&D���Ѷ��P� P�	SL��l�z(ɒ�����k�C��R��γ���[�|lCê�,�S��vF�Obp�&�����y�7��-?qB�
q�G�$�>��V!��)�y�0L\.����)wg/%����ZW�7������V;����S���:͹�B$�|���;@��A��^���Nt�IXY�������*���E�ڨ����)P��D"\�"P�M!��a����K9�.EIߴ�(�@�n;�b��hרLbI�C�./
r�aٻn��K��5��N#���S���GO����c��η$�X/j�c�OF��=M�	�� �~?�i���w]f�����+M�Z���r��I�L���򸘁����ҡ�0�2�`O�8h ��~��=>���0�N�[�q��ϙ�|'�Y���pW�~0�9y䥤�t�!�]ք�#�˦4
��˚�~ᏮH��:���hsah&�ʱj0�V�T@��V�D���ifjdX��e��
�����m�'m
�o��d�՗\�¾�����ZsR��l�*nݏ�z�+�������{��P�J�u��J��{۷����Yరu�3`zm�D�=�fC,>�4�#(MW��tͦ�\��hqe��2�Ң�]���ʆ�;��,hb:��WЭN� Ebr�GFD�1�OtE��p� ��!FZRw�<\�D�����5���oP:� G�N����N3�{Ndg��T�1�Tt��ao�^Y��]�mG=#�}���r��P��@d vb9��ɘ8Č�V�j`�F������wSB���@�{}���k��?��}�0�aD[��^1¢��T�q��D���rh!$�;���H4X K	È7��}ӳ�H1���L40�
��*�r7�_�:8_7�l�;�iۯe��F�Q#��9T&c����DN3f�x��]TK�����,ٹ�:�?\x~�@�jB��CY��A�������s\z��uK�+]�W�wU��H��q��wD��V��M7���Z̜�׳SC���0�T&��,�>�h��`D��%6j�믯[�a6��ݑ>813�ݺ�Ϧ��D���T��uЛT�PSx�f�Ky��X�R�!'v\��P��2[A}�^!S<�ԉ� m��.�dP4\��c�j�h=THj�w9�����&����FZ�m}3��R:�$_3��&�C�A��v�h���\������ g���סKR����]FZm�GhLb6�!���7�ں��`t����<��L�+}��"'��'������=��&+��_|D�0�-z�D_%R2>�����h�_�}����z$Շ&k���X�R��-h��Gvj+ɖ���D۝s�#�kY��j�6ז���g��炍��ݪi������xM"޹k��b�[�H����F>���N_�V�N�sm�S����N�$
0;*h��h��3i�R՞�X�~��	�5�\�䀵�r��	��m�R4� W{g��[�YQ��-`����b<�cuhn-Ov .�~)*�!JK�A��K�X_�Z1�������N-#�i{]��HxB����R�A�C��%��t�p�L��$�G�~�V.I}��NmYG�_����-���?��Ǘ4"�2w�-���mrJn�S�v��r�
T�j-T�\�)}sSfZ�1����evYT�}����� Ϻ�w�/yJY�O�f���i}0�l@7���\S�"WL-�,���ߔ����ʐ�Z�\V.�H�6�Q%�{��λ::�