��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъœ��i��C�SY�p����7nCv58��B�f����@��;#w�!�X�h��'!�L� -AK�g��6��B}j�(�@����81��?z�XT4��
+�.(��l��w	|y���4��0�X-'4T�(Dx�~-�<=ϴ��A�g��j��H��$N�A�uud�9bWf������ڦļ�^0���%��|��[���a{<�B�/V�����ǥS����w�$�;�Ꙫ�'-u�t\��-hj�uHÞ:�!���2��v�s�0�]�cb�1ģUd;!É!�K�b_�NI9��4.aԘ�f0Dt8�~��sW���,����Ǜc[� C����Тc\x�Ɗ��vg૟�x�]tx���^<L� ����W�·_�aX��Ѳ��gE�o�!�ᘗv(�	.���=D��y���>�L#��=�8�z���0K�ҙ�T����H��8�[�MF��H�S��>�O�����������dbB]H����Ųnn�a�6t���.��͠�Ra7*���?����U��!������F��������wv u��r��i;�3���0� ���Kܭ������	����hsZeu��Ϙ�¹��XKw�j��#�w��D�y:��X�$� E�N����7'^���&��O�k}�T?��g�o+�nm�0/s/k��*_�dE���,ܗ�A#-q,s���Y �K��#���������Em�b3��Ϡ�v?��AL��E��=���d��F�>����H�g�e"8�NwF'S)�A.�MJ�ލ&��$����b̴��c0pd�Yt�qk�~��!��kq<�d����M�vS���R�Q��31�����b+����^�eDu������AD��ج�׋W����Rz�P,@2R}e�q��µ��OS��X����!��0K��;F��b�To3� ����̨�(��Gq������`1�����4�G,���&���^y�~<�ҦDFϗ�?�UQ�(Ǿm^���%���&���l�/�m�جG�b�t�٫��H���m��*1���9eH|X�K��N�Y,�+�ڝ|�F���8հ��F��o�\��6�b�n�)�z���$����C�I���CH$F�`h]J�����/�=�1�ZT(Ef��&�R��=#�b֍<��n���[���Y��@N����^Z�5�=[{I��n��������a�S��{|/݃h
�F��oO%�N�\�%F���N�
�VD�c/) ����C�[�h��"*�'�ic�^A��L�<��n�l2��v�E���z�S�=h��9=�����OI��־ɫ�͗�K�Yz�km;��ě��ч
ܧ,��F} ��l������cJ��s�iy���9f&Ci��������$�t3��������(J�SP���"�<ޣ��;ΠM�D�W�^��rՓk�ҢN�02��oD��$ݡ.*4��FUyU���+%[�����6y�9��"������f�ʼ'�m�Ŗ�Υ�a&q��2������	�o=�W.*���ULV��  PrSļ�k�H�L�c<�)����_�H �_�}��#�qɪ�	m; `���'�7N�-�u�����o�P/�0�����Ih�
[��3
���?�ގ�n:ۍn�Tx�����oyqL����nQ�B;8[�Q��3��])���h�k�a�����ϛ����A�`��^�Wp��"��v����CmP�Q�Kjp���z�\2$��p�x���\�%��P|��9a�|��*����k�-�'v�$/U�^���D	U'�.\��h)Ҏd���K�������M��®$B�c�;Ԭɥ��z727gE>����解QfdIq>jmX�qT�4EEy���]ԉ		OE��)���9{�Mc��(��/��_�N>��"%;��T��7�]�hm��}
Ʋ�GT�&�}��d�Hh\���sb~�O$�ؿx�n6E����m|Q �x��3M�)�%�NO��r�B�0�\��6D����s6�0�9�4����|��������%.<�Ps�|e/W����_�$�)c��{]�'$J*6(����V���KN��i�W2��d����3��/ql<����r����#ע�0u������� ��Mx�%�>--{�엄�8�V��z	����Y޽�Y��W����`۫��i��qF%յ��B�y�� L��m�
i�2��=h"B�s�*Gi����=�b�Q]��u���:�,�5��R����:�߁��FϜ5q�q6�똟M�=�3�胪�6B���f�e�p���6P�	^d0KtQy:�`�ir�0�n��F.�KtoU��^;���쪫X[�5�`2�f
e}ֆ.�8k��`~�l����z��[�v������0��]f��%��0y�|~�{��&�D��h���o��O�^��1|�f���%�.�٢P�+��uC��S� �"]��/��x��??t��	��b��I���.Ox�}7��*�Q�&�D\b�OIw\ef�:����L�j�f|C����=�\PBd�Xs�`�C���Q\���ǵ�ٶ'F ����w��{�G2~nWk��1���1b_�u�1��u����Z:�V��.��I�O�Ad]e�O�碻��u�?M��p+�O'�"&�Bs����p�+\܅�Gf)z
��亱�Z >l*��E$�QFt26�X�ڬ��� I��LCIAC�\LS3�i�
��&�y��#�j��r�V�:��<���4�`�+Gn�����5�� �����kضH�a񖩅�cɽ
�y��B�H��|e\P�J�q�S�,�bemB/���x�H|R$�8ԝ�k�ŉ�8����7kv;�AS����`���qr|匵��������[\D��a�Jx����Q�:=9�4y&��� dL��3������Ad*��y����t�H�a<�_�.QѺ0�z���#�K��(�O����q�Oԅ��n)�.�C�9ׅ�w�<��W��*��6�a؀�3ߺ��cp?5�,���3�
�g}N�i-X��	P�T2B N����"	շ�3����'Ħw#� ���P/ւ�ج��sRtx�����(���|������ʜJM����t�QeR�z/qD�Τ���0�ޖ��t��iu���&��Iz���D���o�b�]� �w/�"*�h���&0k�ɛ3�+29o��
���O��`5cq*�EYRd�@w�m~d�¨��p��	�"���
p�~%�<��F1�sB��Z=Si���!���q�Y3��X���o��P�;�ѓ���U2���^V^c�+N�5���cw�"NS��޿��ع�gdƥ��[ӻ�Q���gz�t4�6�ZN<����Iۓc'�x�o���ˠ��i�\�稙q�yS�W�,40x'��ӥ�m�:�֊�*i�hIt��A�E=�OC"	z�=X�U���� �O*�+.��u�>����"`=ܢюX�[��g�j�����8�v���Z�����v^>�C���g^ԑ��H�I���Ⱥ��\�DZu��8 *�liH���Ul��]��i���a,*JI"���i����ϴ�_��OX�k͉$4���?�05����A#�3H}%H������]�Q��A6܂�ч_%�-�,�c)�z2#���,}*����C�~���m�m�ɬ�P�;�8^7�Z�!<��2����4�Q�V`�P(�3���5�����=�M�^��2ms�@�إiTD����.}W���#�Gp?F�"�h�3ۛ�Pw/ T���uUo�l����`�bh`c�|6�?����iL�J�F�$�!�V����SŵPk&�W�19��1S��� ¶
���$p:te�]��Ob��&��!FZژO�xߐlq���f��'?2PZ��eI��6���YW��4�ZK������1�v65>�usI�0����{��WP#6K�a*ȵ�BX:D�==P��9*(IT�l̽��Ly�)������ދ�0X_�0��ؔ.RV5, N��ku/VT-E���,5Q@�,(\�f�ϯ}?�7����1F�ZoQ�H�N��:Ay��7[�F�[�G+������zf�u�۔=y�+x~ʭ&$׻l�HC�mO"Ž�#��&{�q� ˍ�J2��)B|[�_u��**b�n�ڝ��y���؆���	*�.>g������O�����ezϺ#y�զ�%��RO�x�'��c�މs���}�  G��C�/e����,o$
(�+��%9H�Q����ķ�u�?4����㾱+$�8n �y-��K���Ths�����{?#�pF�d�h���]l߉�d���pߜ8Զ�@r��nI)~�[�猎PAY����9�]�\x�v�z���aW�W�� �hw����&�y��ڰ��3�ꔛ�f���$'��	�^%��n�{�"3D�=�"���l��;-��&Ċ�����N�賔��l�}W��(}h�<E4�3��҉��m�71%�˃��{�+�k7��M{�.��Zv*x|G�O��-%��c.1V7����sא�4C�*�~�O��|f�����a��*��X~�J�#�f��;ΗPC�g���	;�l����$�1)`���&.G7Az����U�E�ϗ͇��7;����ؗh4c8���x�^�X��ru�������94�KEij���{_j����,Kx�ԏ(�P�9�9��c�шё��'��P���%��G`+�i���M9�8Œ�H�rآ����BD{�~�K3�L)������_3����s�3$�� �~��lK9^_=�3��k�B]�i43y�*�/�S�[&��j���I�=j�m"+ŅF��D����Vwv�bj�W�4���\�cC�`~:5��ݾ�����k������2�R���W��8�[\%�K6��i"I��>[���!�����Ϡ����=)J)�(�pr*�N�T�0�`.��+�!���$=Л�cH��f���SI�.���p��橄�/7�T �U2T�=D�����i5*�d
j�C��K�������?]�0��zB��,��$PT3�ݨ_0�c ��;h�&C�y����$3!��xoz�<����M�@��	�˙��v���(	\�j��ʎ�� �x(��9����?��2~�-���#D���6#�������7A�5|�JC�a�7�VTG��sТԈⲡ�2`��ɳp���|�H��V�
��u�q�Ǚ(eX�M�Ί�0��[T�����~�<ի%� �������w���Sby�y<��(�L	�N�^kS�>��j7�]��/y^�'��T`��d�"����,0���zB�W��7���
a�T~Zrڴ�-V4R�#��}*D�W��f�c�I33:����z:PX�eQ�	:���OT���bf�'�<�g[S4w�*��<&wr�w�ʊ�������f�|�Fb�A�iOT�'%�g����I��b⯆�gq0��-ӥ��38�O	S�}:6���|�.���J��lvu�����f�f�my��KiW�pi��Y&�<	"��-�c��-{�Tc�}�	?ǘLe�e�{��ey�'��ݕ��K>�_9Y��'���%
>�G����Ib�|��ޟE���s��(�apvF�����+w�<!������PGr��DS|ERKcⲾ!�~�u8U��3�^�"��*��+��Y��*�ss�?b�϶��6�;���)X��������;�������g���'��$��&�=��&�M$��@�KLq�lV�~�w�1�2�?ޚЎW�H�i1	>TG2����3(�:a�h��$Ŵ,�)��:��Ӡ�����d�K��c�M�T$�.˰�ދO�u�S���� V ���OU��9���lO��K ȴ2 gj�{�������=ƥ���#IП��qXu�2�$�����78	��Hx��
��tM�J�1��nΓ�"��66b�w�jҐ0$�C�`�@��e����~�.��r�@��8��q�(�\\�P�D*H~K��^F��F�!<�c�.�e�u���'�2��}���k�˺����'�sI� ���=�4��W~�|o��2��VE�`�J��,F[������k�z������i���)NNHiQ�	HRD�?'��v� 5�GG{��B7�=��g�~�&P#E�����3�nwk��5ɻH�ȵ~4~еSf�kd��L�����j�)�]]��Ut�<f@.@�J{�͡˸đ� w���"a�[��֯��
����\ �6�*�N��ː��dW'����m��M�T�w�k}zo���0����X�q���е�>5�4}�N2~�>�;u���5v��kf��N�W��2����y��s�ʙ�G����vض���k�x�Ǥ
0�'��@�:�y�Iz%>k��s�|�oi\;����A'Eo���+�yG�o�{^��	^���oʡ�{�=t�P�WiװJ� ��;Տe wlM�d�)N���W�s��ľ�N��v���r�/���,�˟��]<����.���ӧ�L�1�Y����=����f�v�A^�՟���2��CɁEN�;j�qE�(�m� � :���f�8����]j+���mL���D�X����R����Ш�5>
^�qˁ�k���%W��yi�Z=�M'oG>�]Ƅ�"\�KU۔N�x���K�^�.O4�sN^��Nh&>��H3�f��E~�-�)�#��y�y�+Z��o�9�0�{������Zl�p.:�X��#��,i��"��ܠ��"X�g;nw�������f���k����ݺP��U�7�3(tJ��4���Ԋ.*�W���Q=P���)�NhBv�ajtf2tc�ۖ�)Bϓ��.�ĕ���@���>ֻ���!�m�Lx��'#����&6I��k>^Ys�3��z|b�~�w��f]�#�l�ۓ�}Ɏ���j6�+�<i�	�N.kGE��I�^}󢭆�����ʠ����{�v��)��S�j�E�1���9��&��Ą�M�`;�����q�X~r&���٤���.0�_rs�p��o��y����
�<�@@���"G�6D���.��![j�q�Ӝ�+��1�	��3��[(����]���]\$�N�&��S���iͭ�"���/t�q?�J*}g���8��D�W>��|5�o�#U=��>��Ṟt,������\%��rTԾ\M<�܀
�+e�����2��ɧ�P�B�_�%� ������_B�Q��
,��-���s�x0&����H.k [:���< �)fj����Y��ѡ���<U\%0	�5��bjIw� ���8s}N��ks�Y4��to��~k��E��%x�0�	�|K�$��;J�TރW�l�����b0�4�N�	�[Iٵy�ರ�]8a��� ��k����}�p�g"N������1v��R�wM\ۑ��4���r�:�-	��&��f��oI=U���VE�����Hs�q���VQ��Ԛ����ñ���!]�MD�h�<�H�` M�hO���E2��L�J�І~���M�:U�f��&j������Z��k7��H�����?���\d�J�#����yi7T�t�bڒt�Ӫ9�f����pE�����_?�����T�j�<t>Ӊ������>��z�D9�`Xk8H�І�*Zx�|��k=��X%}WSf	+XS<M����4\���c=�Y%q��+�ץw��g�r%�%	:'l<w�T�od����ދ���F�%p��;�B
�Uy�Yu��1�r��o�y���kIp� ��v2<BЉ%R��.:�VZ-��	�fz� ~����J�$yx���bۮ(Pv�� �=o�/ݵbǴXC,�UnB��,#v��3�`(�1Z&���G#Xw�H��do����^"�X�?��<�\���n�g�!�P1�}�N(u����X��Xi9����{M���r�N�V"% D����BT>:hʨ���x/�3�I�x�����!�_�s��&0ָ`������>Q�����zQ�^���~eW}��V�,~���#%8+��dI+k�b&����"p'�
�#EĞ������8�X<X%Oy	G�F�#J��1��fX��?��Vԕ��%�������
O��ϑ ^4⠋��I[�KRKma~a�Y��FB^0\���	�"y�S�+(�&$'�ó��Cj֗�vQ�!��ɽxRC�~�nW�`�� �ԝ���m�ݪ��I�[���S��{MLy-"��җM�&(�eB�~b�Ӭ��{̏W�Ex�C5*��y|zS�K�.
�4���I�@*�{����D�8=䳾6�ݩ��n��*1{%�%WOo:jQ6�?�*��]���n���^�p�A���%-��9��ߨ�^D�7߯�-�A�`>��
ۋ1�1�<q�uu+����"bD������o�֒�xM��qҚ���9���Ǽ��ҥ?��#������A�2�'��P�R�\L��0���s������Y�@��=������]Awq~`�$=��X����T�lV���B�	\��<�r���F����V �i����}x�'�{Ή�h�aJ�v�Hչ��nPm)�2^�l���Y��~3	���b��{A����ֻ7�O���O���P%��BC$��7s?;�xjv���|3Z��d�����kS�K��C߫�� E%�C�C޹��D��$$~�{���#,f���4�W�{IuJ\�A��| 3�P&Fh�g��[�P|?t�&�IU5M��c#�!��02/�nӷj���uyl��Z���\犰���Y(3���)`>�"��в�Q���N�/�����rO��7����˻�)�#�?�!=��w<4�O�K*���]��^� �ѕ��	���QNۧ���ʈB� �;+G���4���]�ѫ�t� T�O��ui�²ݧM���."g�u4�ӁVI?�d)�"?�+4ۊ*5�S��C2K9&:7�`��Ŕ��FV`A9���3�sC���T/�#s��2ϩ*�˞BS53�f��|� �	�px�l���SsG�qܟf�'r�	��I�Il����d��u�4��l�F�ȏ