��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7`��V�b(�554C�3�o�O��D%�4����}���C4��Է��K7�'����e��֨VF���o�o�#�{���KnT�N
��cO)�m]9|z����X�z:=����^r'X�*T��j.�=fD%�� P�sݻ��BZ�K!����M ��͚\��V�3<��ʡo�Z�6��!�TK5s圢��e��R�c����"�5�9Ĥ�i8�Ҁ��Ð��O�ŀj��I�5��}��H����]���R�+��Y��&:�r�a��?��O����w�Q�0��5|��'6���C܁MD9O.r-6|).��f�@�v�&��]���社�{�}jV�Mi�Fo�vf�O�~R�Ʃ�ŧ���"Z�����}�C��́�54x'Gm�	�I-ϟp�Ƭ��38	�ieύ�
_M�v"�s��XĻ��iI�A:y槧�m	����E&c1�&}�o�})ג�7�*�d�qC*ndot��|�XYӳn����_Y=~�0���ɲ 0��Ⱦ����<y�0y�9f\�΂��;~�,��N�@����4C�\Hb�+��I����1�x��դ�b����B��XUA�X��1T|�h�O�f�*��&��T���Y�s��^�:B�N����Û<����N;ֵc��|�N��@��*&���EC;�ss���S�^`�X��K^(�i�($���#+%���w��ٗD�t-��:^76p�����#��!z�wC?�����{�F$_y)�����o�&BF
�rJ��������.�I>�9AU�}v�V�^�׭l�q��^D��0ד����2��u�+[(�"��A�V������&�֛��o����"W�d_K|G�c��zsI`Z衤@�c��*d$h{,R2m��!�J����s��R[�`��j恦�[K�y���BMm����z6i�(�ΐ�8Z��wUVU�O��V�O�&u�$Q��\�$6!`��q�d�<���EҒ�4M��Ӊ�*�ی$��E����6���� A��qIk�7b�����Ղ�Q�ۚ���~�>Q�EBl�y���,I���� f��/@��ʝD��f�$Q��{A��'�{��yĊ��)z�=��X����p��6���e]+
��zr:Ji��޲��2]�ZȈ�48o
�	GH�Tozk-���Z���_Q���9b3�'G�o��W�@$��g�J܎sUn}���ٺ���*!��n��R�D�k�D*Q6�HW��d�������m��;��E?C!�d�4K����Ȝ�2-�Ug%�.��y�_���V6�����t"7Qsܨ#|�zA\�aFʴ�y���Yu���k���R��!5��3:�H�$�c3!�T���R�P52n��D	����;%���4����a�ϳ�4r�9A��9o�K%� ����9�}^�u�o�ϯ��?��qNM5j3^	��[�6q�ZGr��g���,��U�c��9��A��nd���Û��(�}��EuB��qƮ����|�p�H�m�HJ·��-?�qW�^L�c���u��̽�ʳ��� o�'�G�:ʲ�
����Q��>\c;���`�:����<�����7������\D(|���?@R�B=Qv�����U爀��\�	tF��q�3;Y�	�����C�e[�sX�kՠ�����L(��ʩO�m���9^�%��9�2�IW8�X�rݭ��%���O��f�vՕ��]�3�|���<K���<�������0�n�_��F���V���2,⭽�ؽ��S���Q�+���!=����_�}3d�7]ݜ�*Qg	0`�l{a��G�9쐘H�w�h&���c��<yr��|���v�ߎb��mI�3��$LKq��3rgN�;�4?R���2ғa'���@�$���
�i����9��-��ݽ�	����7��v�4�$Bg�ۢsN��j�N�-)�B"q�m�7s��ץ.q ���	M��V��t/뢃q�e�����pR�c��N����/rF\����^��)Z�|�K�E��V]���*���ze7?�W�h�U�ĦQ_*+������a�.�o]�і6T�Sqy����;���wZF��+��N��<�фd
�y��욣�K�H��{l��,�so�S�*�����H��/C9�f�;��3\�{{p$vU),yJO�i[��V��5�k�[�^Bo�t�4�@vY3 �V����J+t��D1	�Ƒ��SI���
�������K�=w��ٹ����2I�`avCs���q?zN߳n�A��`8PzL=V����'�q���̣�<{������q�E�PS&Я4����r�0��jO���N�j�V��0C=��'jmb*�w��.�L+��u67y��w{��m��;{]]zJ-|����h��o����vH��H�����S�0��:h-'���l�cw4��g6h�ft	�Q����x��د�$0$�_3Ѵ��Le��QR�6I�r�~�8Z<}��~��|��eZ�g�p!�")؂=��X1�2�?&�jR��"�^X��^$�4c����r=9�Y�0�~d'{ojܦw�*�U�j-��t�)yϡ3�0+N@܍^�\�[&�(���b)�g��魧��,�<&8�f�lq��Yֱ��E�$�u�>��l�l@^7)ho�Ig�;�J��T�)�f=�2����&���B�"�Zu�*ed� ��c�``�5_@d�z,�O�������]����<*f>A-*7�G����7V�K�-��y��G��	b��ّj�{|�w�N{�ӶՈ���L
(�E�ᰧ�:&��Tu��*�-F{�3Zg5�(���<��\�ԇ &5ML`�>��ͫ�l��,�T§ߒ�U|���b�O�ʀ~ơ#Ơ�:_�ٞjң�A��^��#U�<7U݃Z����(@�cl�m1��Wr���@��+����������4�S򮕚q�<H�8ϒ�����-z���AX�NOno���E׌$�BY�u�gg8ī?��Y����z�X0	�G�J�����(s�j�Yqd���ܙ�;���U~����P�dR���N�^mN�D�˵�5�O*x��m@����Id����!X�F��^ޠ�:�nm�ڨ6�����:�YHƱ�������E�>[�H{jΟ;.vխ4��P��sܴ��\f]�b$p�����-���6s�!T=�.Ğ���և��I���YsY������Y�1��5�����_{�9��e�m8�xd�����3u�R��v��~隒�5+��辆��B_��S�������Bp1��+r�5�kl�ꑶ>8�7/ŀI�-��r�5 ���@��Dk9U�
7����f)T|pki,�^�:�e�Ʉ:=�u�A�^%��o�9�O�؇��o0ޥzؠ�:�h|�: �ض��@}D(9��U�5�����EQ�#%yY��1Sk��ڑ.�њ�18l�H����,��z����}�qa�r�Qr��?�f���'��i�(��
"�(��j�F�k���y/�����H��H�6OF�:iqh2Q�θ2EK~*j��u�����1�q��v���(؈��<�ϊ�ֻف�!۾e������E7��c��c?]rX�n�R�J& �Ӊ=8�<@�^z�<o�p�&Wj��XyoCY�k&�JWp�\��ڪ�>L�TW@w�٥: �
t�>�I�sݝ������}H0B�
ï����d�	���J��E����Z\��7�U�,|���F�e��sڦ�(Q��x]�ߨ�����-3jUW�1=6�c{�y"pD�.�c�=ό��R1�E*uiI �v��A�Y���ͣ�.2�|�VoK�?��;`d��b'��(�#���җZBV�zj���Y���Ju�-��h�f�4�����-�&�3v�h&�L�'���Ϗʾ�)+[���eV^7��8���8w�jY4g?����*�-=0=�9
.b����r}�hC�;�:�ZչJ9�R���0D�B@g�M�ؓ��g�k��r�'DR��;����e+�����yg��