// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:38 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rSj9vZSmP2Tb5xIyisTj0ye+zyjnS4TiOAIuCBEb9QFDhpA/AaIiLbnl2rB6kn8e
g2MUSL4Uh+CNXgNcJy6856USJ2QkG2ypBxQc6FG+6FL1CeYlio5/S2WJFyw2Di7t
M61bSUWf6bHPtTnO4Bnp3GadIyMeI71TsEL5IbmDHFQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3904)
c3Y9zM1RcCXBAw3dfcrZY73VYj9IFE9i79+OHRqxz4A2X66LI2pF8Ib3vKtRsmB7
EcJy9kMiYBiS2X2U+iUXe7Jt04ImX9xRYrQnRQP/wAAoKViepr5f5RXfbvrYuiTH
utYnXjIYhbV9UgljeoQBZ38cvT8iQIhmDo7pUpVbV4/LB8HDgxM24S8G61YFizYq
xv9nYXvLaLa/vYJHBUig2ZbFuJM/c9U4hezWUsN2RRN2+nmMoqo6gZVuMzACjlc/
BI/JP4X34IxThuUsUSAh9i2qQoBeBYVYwszjzPm3cRSxNn1RUG3TISIMoLaDQ3Xu
XOpACklvYpZJ7fooUWHmWAvgcu4WxTslObRupA1XvPfo3RHYmOuUK9xaZ1UUBsba
vkDiLaFQEPHlBei05gIwDMJKMkEChRvyURbG277OOA2qOWFoH97yYqHDxnUiM1wL
fQWHjAuMFg5rVXJcS93/C719Ckh0gtKno3rlVbxfAkvdhJwwPUkDtMQUJSAPz+Fh
kYdaGLROfJGZ3SFczm09unDCv7N0bZW40wdkLh+hr8t5a+8+D2hXUySmRezeXs2i
qgxk8p+QgzZWettBw+2lXEensBCCG3ZNkHKuHgo0yrLsQgv6bYlMcUSAFSZVsDW1
dwqU6MjxaAkJQMkLEJY1A2rzUih9fcKzWZzoDMkbIrOgsuBEm1E2CTldFKGcCamC
w5Nk4842M98IHKy75Ma2nFHKPuOExhig9w2R2lvnaMy4ZoKltB7esPqdBr+dl+zB
vfm1GUq42i9wkyAB4utboBfsWP+1T7ZKFbx8wWzNMBwKgsoj5MLaujxje87nTJLZ
sNn7dastAAea7UKDNJl040D7ix6c/rdIl7wI8mSbu45zOkpR/REi49GfU3wL5BuT
/cPwebTecpAlGtJlInEiAfpZso1SvXc0XRMu9WM7zIIZNp6VU6BOnUZh2E9jl1/V
P3aXD5nicJ1peQg6m7sztbYLF1k33QvYuvkvEEkmWd8iex/xZHjk9dkS1u2nVfeF
0BliqjHjE8RgzvZrtSrSVB6+rT5WiiTzo97L58K6Fhw8zOZ6Ld0ZiIH3AV2cJIeA
k9EW0ZE3XnwEzlEGZbed4vnfsQL8q9ES1K/GcDc5gSi7PqQPMENvsvRKNPzyYiuu
V78qLo7YO4J+WOQydoWrsQOO+n0lc2MH8lyavtceCdLxWhqMtT1Nl1N+J/oPOhBJ
1qWBTst4cBEDbfbfH0lKbMO/pzF6Hpv9Ey//Oi+N1NlXZSK50zLY0cy/8ECy2Ii+
G20/0D+GBFFtisGoHkVodU16zxC+ad5yJEVk5KeNZykCVlz/YCXzBkFk2neuvFQ2
A2wjJncVsTTc2HfQ2XmqfTe+Wy5+9Uk7xEpy0Ynuic9jg/V/qElltAU/zQRWR3Ng
fYb4v4tBNDeCBNql8OfK20C6glcxDJzHRsOlqaBBGAgj7HmHuWx3id85KK0bZGf3
+Yj/Gwc8m6uwuN6DfntMiivlv5+LHq4cH4JGfnIxWa4l1doL7/ou/odW/cHa1XRb
BitcaGn31CeGjCg3azcK89lXaR/dS1pW35cJvgE6gBfjLKZ0av04Sb3oOVR246YX
zGtG07y7RaM4SAJ58JouH1RDOyoU5/z7FpwQz7L7obyg+hDShi/1JNyyqIn0ugR9
dc/g9au4eheneEi5gkoZgXo+Qy7PpnSDgKF+eks7Ojd0vxQIuYcuFUJduQwl3fhl
O3jlMVXpzJafUeTNjar30phoVVXDp+uk2LVAdEFbAsgexpe0Q1cNgPL5A05nRaDX
n+K+Fq2pKUcXjb/2U0bV34HX/o4R6IIqwWOy/HUQbUViXh2X/fd12ZzyzdEUImfO
e+VZ6L8+tsEuuRt/Dl6WJqMKJ5TEBD66EoMc0qhdRH8P2xBIC7ApGZBPez/WKXeA
zX1oDeveWRFoDztHHLJLUUAkIGdc+e8DKSYCgL7ddlF+rOCbHezcWLUybrUJBX0T
y5QF0Q7DookcW3s3L05gXQFfOQnLL3dbzas4m7vRzBiXXBPBFmbfonWBgnSiT7qK
Xktln6d9VLL6ku/RHwi5eNqpYsu8WTLyyGKYMjbw5wMT7TTszu8RsB++iEcsX1uL
gXVqH4Eu4P0EmNtpJJV2jdOw7Rwx+mRd7pi7lVpp+njBjfDMlJTvK1XtOCjM/4WP
rircFYlR8XJPIESs8oFawF6onfIM3RrnCKUJhyU+PVom4FAH1d6vm7ecSV0sUuib
ijqCPDbXmvNSP2FIf9leIpdIglAyxY8c3i/yoryZKzYvJA3V4uEymensrlLF9h+R
awQDGzZrmH6LrOGP4vHhCx6F6f2cSYBKLyVuckRJyoXjKwVyno9CJjxdOLytwCcU
mflgkBXCMPQBwIR8H7M2bbXCRjFmKSldAqsjnRz+U4jSBW8cTebNhpe/Qo+sndot
3tnOfEuXj4FGQ6GFHELnMyRmtA514/bzLfnkERpuScirRWFiZLx76Y+rwhtOVunK
xAVwAM84osMofwsdo7ffIdypFqknLNFoC8M0QtHgBsnZdPtvHt3RmdUQpWkSxNtq
GR1s81a6DQ5ke7gA54ybP6BxH9N1uEZS+AfkkH+nwprT6dmtADtIzfwELTKZz1xE
wGy2cJBBDijOrJV5+ICg5BTr/2gk11YTLh59ASqRNQaek+piXe145LsGUARKOEUn
GviHCpooYsd9WVkCCbZyMkMtjlbTgJVcZnYO7M6b0sHLbbg3Yiys3/IdSF4CTvrI
EEJQa5DEXWkk8AKsmSxHam0/pdA/fPPnt0B8OstgRoS8zoyj4NffM1h8JY2OTVu/
Aj+D8Zm18oG8LPClszOBgjgpV3WC9L5VRNBVk45Z9krGKJd76sFN7WtWoAMK7DM3
ObuxOQAEpqLgNvBgGH6vHyQ0ZXr+FiBcWKqNBhAkTXlhuZbdQP8Zqsin8BnWzhhH
rtvWi4hyHW2xFXiBPznDow46U0f0P/jOQ+9FH9/BAMN/mt72JfWMecCb0MdN7swq
qn8M/+NzxYFAdrrL2vp8JlyG4nUsrhf4dGKPM2r0fTsFn3Go77UQ5h9fxkfwmkYM
0dm/TUkOeQ7WxwshPahh3ZnIdUI18tE7k9uvSULeA+Tdwsz1uuycFmV0eD1z+lyS
ory8ieOv34RSmobRtXA14qn5SM/msxZkBkzRCOykcdzLxSt3Q/ArQ6O/Cb6VgkS4
UH30pnvw6eKTHO47wyKYl+szhlpUGxflp32274kUJFhWk3nHWpwn9M6V8kyHHReM
u3dnAQqoaqw/LDWGjaG6II03zM6HpctwLTLQhAL7FohQ+IhpL6Cd9Zh3kvQow4AS
8dHooMWwcXl42zKF8g9xp9n7i86gjsTqn9p3Fy+nkqRvxAyXU5hpLx6nV6vYRL7C
8EaxxO/LkHaNExz5VdKv2hRacsnbEhbrLgy6WT52vO8jEM48/TwWYVm+BKP4nPBu
qQtJ2swRjJp/kQujlGESxQ6BTI5UPvuHea2XtmtqpQKqTfHqhKlxmPjbG9gi49jO
Jq+udPkd6L7GSaGJKof24McEKLI2/KIBDCpf/0R86Qh77xvVQcK8L+DeSTrq0mp7
lWceDVjFsrkVeXgKOG1BSMfbyWOJblcsHqofl8KB3YQJh9EtK+D0zTXjDL97k9Iv
Xjz2//wGk3E8aTEg+gswievOG7GWFRrLmeh3yXG9Lem+lj44ki+8vAXpx5A1fSmQ
l9dViBhRIHvLtp/bV5YmfDU0i7g5PjMKHPuxpdf9RfywUX80Ld8TbyJNJIl4PVG+
kcG++0G13JsA975UjiokzZZLkrQD8yqYQBsduWaYRIyZyBVxTKYO+ECv2RQ0mQu4
WyQmEajZhABGasfqK5Xv73pMGqTcu5lfOO9beMsGX0pfZh84/g7MXbhEGNXrFT3c
ekMV81nYPzqC8BfLoG3CcVn1/T/KPoJklLG9xCqmMoe5erUnDiCZuGtSRgdhZZ/i
D8A5SDv7NJKvR37ZFs/rF4K1iL/H8C1UWU7KlL3T/WtA1Nzb0zyPwtTkL3ZqHjB5
j/9yU4biPZeMe1xdP01i7V9L7/aNXbImFbHukpGOSgqwcwRPoEhaCu1z07jQ8wgn
kxppBrZHzNsR7gfh5AqBiKkTaASlf6CmlkxIw7pum0zmVjjf9fg+gkrBCUsMRwav
/+bpS23J30S6VGYb2dUCoFAcplpdms3XFS+Wy/Kux+hbSvVJ5E2JYxVRY0bEJYSc
yd4x9ZH49hU+YfQhGtLdQ5BPk3V5MCWDV/aFPfmJ0AI4iSUxZ5t6hFfZ3TeihawW
OuKX9N9kBjzzSV1LBzBOI00HApr4R0+HzUc+1XoOax9MisCTsZ952aiTtFBOoEfK
w+jm6QmvMgKcgha/8j3XMpemghoveCJQA3GptLZr5mV7NL/kGho5PzJAT022Hru4
yyll+Z4FpKjPBl89ExlOWBK6BYyqmpd1HgleTklki/utQwGTWPsk/gR1J7+rGqfr
kUX2+4h14+/fq+QFyTlWQCHhSj0ZAkZrFS3lXYq92gedBZR2TkY4ImxD6w7ItBcG
xsXh5shkD/WblJo+EMC78pzf021crGBkNLfWcbtNhqtQQ8c3CsbHD1TVrjbcVudQ
bTvR7MK7tWtjEJN2YZUWnkGQ2rIuBxENfrjD89GRBriM82LGPuVh3wfb6/m9NGgq
I6UFNkddoDiFmgwNtTwk/Th/eGE31JUoHi8ZH8Mz/S1QFkndHAEcTTJv0Og92A0I
f0P4xkmAL2qRRIiQYx1BFyBREkk3Y5jOYyTfKEiI0OZE/XB2V4wsoaYgHh6nUr9H
qmZR7jzp5VH8fYNDE06mcjwIxclufSzltZaJtGTt3RHoZFKAOLgQvtWzNnbQ8Aa8
CPeNHlbJabg3ufEqV1tIHe7/G1Xha1F1X9t8Pd1vyUyBqYUBL9NjcQAxA1ztJS9Z
BgMofVlx79kZAtZqJdYHKYwPrXTWUUQINRSbjyXhy5jBbQrMOR84uNM23KBwWPUW
3eUkaPa/9TtLT8Df3YxnQTfrEd23mwddv7WXslpBu29QJp4ZdgXT+MkYYao9a6OJ
38hjD/aNsOV/GEzVFLoVFzmIDSj9nCZXr1s9m+zhAHHvOdpkObmDWEnShPD9P85s
yCw3y3mcOwD/LZIC5Ik3977+dr3ax1YAJUobUdFnAqGf2+c9nmpqHLcXWEZ9J/Xy
JgnXkIARmB7OEk0zhDabQw==
`pragma protect end_protected
