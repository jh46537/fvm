// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:58 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BObe9srPaIP/yVdtYUMUoBl5gjkc5cm5xFMuSniz2JS2DFWaXX2/3urwt51zXyCH
XgcHGV/i3w95WdlhHqe+L6kT6/rJAChTjcYt51JEGPO9rO8y8uOKO1dqZ/0H9Dqf
7zBthFMKRnSVYEXztfbhPNRzuh5b/kmFP1Yb3HauxtU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19936)
X5iKaJ8xG5wMq5jGa7TQ69xvI7E+Ao9TADEQMgr/ZFCYIy0gcmg4l+D/a+X6p4Of
WFENUXZQ68I3svN4Vt8eFOA7GwjWGPl7f4iWlqmh9EGOe93WcFUxfK9sAA4jG/k/
rCrUiKBan+8ofXx/rn86Fd7ITJZbHffSTUxsIWTbRLdqRUt3mviNizuySjUwf2kB
fPd57xZFWLVDUZuDya66NgoI9TYHxlzJX7I/HPWmOtb6oLp3/70jk60ui4Vo8+kL
MUTcS3IAfPS0pVRA+H2VnrmgQRNmRdJFmmnuhQjOc/GLjVdUusjY0XmH9nwzIQwZ
8OjA1dm36zDU1HnuCqqQxj9N8mc9a6+7k3pWSxvQFqZWmVApQPcm/ju/HuMv9+yo
3vICdYj+Ya4f+pRCuK6imjSlN/X0ICOAX2Jm5ILHb1cvwXZ//7jByuFrAc/5sWsW
OK2n73B4uazrtGDG0nZOnsH/H/TQDbqZtHLxgi3IZgiqkzIigudyHHvBkEObhTbP
ELkfmmgAaE0x9S+XKz594s6fUD1OEOFV861EXO4VYWfbdCwTDDfWwTcFbQFiLp9Z
+0UQccGhJbjfASOSVudBGW8y7Uhqfm6C5Oo2zjb7nmxVbzzRXDJtcs1XWmnm2F+L
ItIzZdSADl1kJ2q6kEo4I58Lg8rjzvCLI8iR4v68NysSDvymTwf73hUuonvt9voi
XnpNWqIze7z8M/dBi9XGKHfZ3LtsolZSPQalfnBYtBDlKhkBVnFnMO2pPmWKfrR8
bC7LR6d53OA4c/LvFEywGA3esQU6nNEY6NzF+2q6xcAUa6ep3WnPZQAwljvOoYgc
ycxveEciqHDnGeryAv2wIeF/4cpOfAYgznasoOeMvRHiUFJnC7DXw5nGbJyvuTT9
6CVLc4f0UHRa8TyWwrXAobLjXAl7mbwb1eBGjhJaKW6l/0Q3Qb3+kmC8NZjglTDn
mnO/1gmP8Xcc0HM+LGOuYjXPCWzTwV88EGYilpZoM3Fvvlzd8HJWMFfjBLnMUMGi
SItx0QNMJQjOhvfPHXqRaUAzX2FiRJ5X6UGmhd7vxvjz6kVmC3OK/yp9luAdmSJY
vmwS9mpmhJC/x6pu0lhMZHmZSrRGCTcrYeVTKBmj7QHY8BpxodG7qC1SHxkkbEIX
43FtLTSeAh1ZuUu0xds9BbTfD4XYVRtdtQtiSdONt+U7FkNrVs041kND+yNwtKqd
6WS1AyuE4/iBrPLNVBXvD2FuC9k33rdz7uZx0yxbAujtTVxfb2DOvyXl1c45dsJl
tKEtCx45BLqJ6QEc1lL6SpG7I+6TyJICVDUcLlKqdhapknUOq6cCn+UHdUYI2BQf
2PSp0NberwchVGy9NC8XK5atq5pVEQrzUbiT/rA5jGK50YCgTYx/+VEGB7/xRQKF
tln9YvgfO15TZDl4Geecn4XDxteEF6k0NvQm0wlPo0XrGYr41OG6m1w3dDbLPD8h
tz2TIjGrawb+5IVp6gPPCZEnWPXar3pYcqNp9TvkHBuGVDo7XeEPxCUKJEKltFNq
RPi8OqYpx8E56kCoMU8DBMOO0s57kxNpq6b+ZoJ8qkJu59KwMl0PSvvLEEYMn9EI
iTyM5vYgFpzd9GBvN+ItKc7FnIaCEh4YamuaY+5QhUWwzb6TEFOPoaFBzpZf+Wu0
Ghg4N+I4BO33gl+k3HSWl119NBVKhQqgQ+Nn9G2fma3CIyuO6zAl5jafiH+YG52u
LhHgqJRQPt1KGogZy48KD/P5Owz/blmoLLDg92z/0p6FERhRLKKOzyGdBsLMsB2W
YOKlQoA4ljmbH0rap2wp/yRG1/D2H8bShwKPkK1InjShZiRe0UwIl4xumdkxyax5
zm9oTpCGUF4RBl19MVaxWD40RiRNmunVbnQhSknXd3oBr9kANKalFVpgeUSvNt+2
ZYZQwZZ6pyfn/T2SI6wvLDwRmkrbWYqLfaCKn86GIopPbN0kBPkHlKZ6T+JRvXGG
9mKaae5k5GIjUCxmLiBtIJzX49ON4KB/yIOHwdgNIR8+bmOMLd4kqh+v04XRw3pg
iQffveRm0Nf3v8G6v9MKuT+XEZSmak1X2hBm6CdgYtDlSB3dYpAiWNXgbqhqaQbf
dSeSy9QyuY1N98Gq/jAu7h4em3G7rZLuZaG0ag//mBPjEaSqpQXfy1kHxo/PX4dp
YxhLS55gsGi7WSmqpocyh28ndzatXMwB+mBkdEbkr8CJHeToVd5Lt8Ks7axtw1Xs
wN3XVNlpqL8C1XEmpnX/tVmc5vvZPsDYcrdCm/mEUiodMasfcyt/4OtQ8USsuxyc
612Gy1B72fN7LaN2mhMlT9pmFCycZ1pffLgrx9FmegEpaYs0sdpmpGajj2WkGi1b
70emgzVLG/Gj8/gsUUvb/RHOYCAl8lmuZLMix9six4W7BebUEz4yuef/wu4+urhQ
4Feb+nC7kLLX2rgYdfmSEb30cthkvncNYjqUMZIrtVF9vObcMaEHkqJV0Xek1/jb
6pqv9FpedkG+Y332HiT3cNspyzRUziLmsQmQNx2T4R5VVDMmA5M7Md/4xnYQiqg3
TIKaMXEdlJVk+gvjMv5dG4lhQuCH8t1Bia5v0RwYpgAJZX1lOktg++MzFs3FgfQQ
2p9cY1ts7cHOYTpcsW9AGG0DdP0oIDRAoJMfkw8l616nLgsNrKF2CAckrmnpWPR3
9C9O9fYj3QSpFquI7sQJXvQIMAQJVVw++eb5qG8wlOxV9K8h6B153YsTgQwBXXy+
m0P4m1brIjhJR9shww0N7ydyZ19x18yGYprvPTyEs5n96bfqClh3E++WDd9r1c31
k/1N8Y640j1IAWeWQWvezvJ3SavJuhci7Ch/vHHZFEg/bkt2qtiBWoBBoN32Yi8y
leJRQItjHs4FTg2xGtxyCfi4U/H9PGtKzB0FjnOFSaHTQqU5QfyQd+SmFPu8XV4w
pGcO7hT8BGkKydNXrnuCvJYMw2+FpWtlvaJtYDcxclixnExSJPr60lNVU77WAXFv
/vr9jcTkyw+dWBPJUCF9gzzoKlZt8EnNZN4C7E7O69FeT57/m6UJnsoUgGn75kW/
XcEJWOGG6EVedpzd6TcbbLgY7cA7F2VyomwQ0qGp2dNn2XNQ9UURvkV1wXQXYaIX
dH+enx9hADuj1HtEp5L9HN7cKyuU+4RC4ZB82/uW77OoaMZ6VgqBu4LFIV5TZMoy
2G+0ifFY+MLAyXQYvVDDOtpglr9BQGh6Te1AvhbfJUCvoXY2Nh6qKhBBFex64rYt
RzVYX7BniIR+EUjN66PSx1l56MluBh4typa4k4NL1rmBzhgK6qqKPZHtkI4q7mSc
JGeJCP9YY7I8lZ+RwnDbEK5LknL7imSuVMGRTmvKjfZXEHL6gc7+FsdlPws2RJuG
XOhNa6kFpmbL9CLZyahRULrRe634yE2k1CGEdrNwz1r2F92LDylJEIFDeoG78CxH
5bFZgLOaI4UutZJqVooGV2dA5PvaDl+PBy93kjEZaDNayo6sLf4phmXJ0aRRoOcJ
rs9Z9HLxTREdKa8PsHwD0v4zUav1IZNX7ccU/QWU+BOvjedUGWLsSw4HsKRpX7Q9
0aq5/8XcJ5NVvU/QsxGjwvGrYhQxKO1jCT7d8btll2jT1LCVjuZ/v0IaIoB1xXH3
SqN6Mubz45cHoLXhp9+xLPW+MLzFaHxcbbNioLsT+SAdxpE3awcTbWOi2uU2DVrR
WbjPg3FNJf4nWEKGoeqfYH4cUWwu1tTvvsIrRdV/e9vOQszfhaPnd6z5dnZj/3xt
jUpN7HJV3cWc1mEh0I72Is5Y+UJcxjzUzzd+aqqAp2hXsoCJVpNm8DL8VN9JFt0F
BXdl9R+vkkH4Ztq1br5s5aMF/KZQ/sfrcA3OUvG/m2GyakIB4K4u7akFb2eUfrT1
M4QX25sCleKEfditS8zLybOFebDOunUZ0bH2og9gSHodH7QxCV1wxEninV0nmFPI
scljW91j7TTsLx0KNEyxB9SsZ/GAbiRBWksDBkS2jnREFGx9ixyCYOTsGLK3w/YQ
xoEMycMQLgIhDhHFEBMmcEFmrHOHoTtXlUF10L33giEM8vYZNsS8FwvA7qD214Z4
U7pOeKLW3fR3r+Kzq2JbvrwFbEq0aXhxXs1/i2kZbj8ejQgE5kkp05AvVdgmD0m/
pNhXOz3mYUEPkdlp0V8r4EadPpzY1Awhd7OtevJ2oaAfFLWSfE4g1riINI2tPEkz
y7RrTp+8Dfp+xkVFYTIGSlFPoecqG3ur+J4nuuvfHviKzduIVJRZ25OiWzWrLcqE
d+mwvWRrlTec5ekM9ZqqCUtAU6HXaQ5Erev5Laic2jdnHgmZ/kemSICcLaX7ekou
/36xSZFWFffLUi+A4FsJ9bQuYFrhOvL1niMdFlnLAVoR4rwkjofLv0QqacInBtOT
lBZvHIJnsN5vMynUHq1CzM44C3euTegPI/iRHIAjzMajccUkFAXCgvqqnpx3+OxB
yfOgeUR+1XdzYPpqwR3JJJe83O+Y4xK+FQQJgnnZOxo6n7A29DGB2pRTZZmAJe+D
AXfTLDc5I9cGzmHKMTNOqspoVynTzatxa66f9jCPKIF/QeeoMOpf9dvVwW7c2ZQM
3utC1/8YbWBmLhplkE7nw8LxE9wVFY62FXp2zpXbBD55bmLepJVaBhwLx5ZzDl75
OkvMR3af/c/ion2OUZjngtWmJ+BkJq0yIE4wpMJjWY0mUk8rouiq9g0Y5HEl8SvE
+UXZq3Clc7FtRWXXsGx6JkgvRRP3KJbzoxtQI/69vHqsbQwxTCuCwh0YN5HgqAaY
ri75uC1MuukEt8CEX1dFmp7FasfGXoDrlknpCJyte9iA9KR0wN1rG+PO3CrJmlyA
W1gebNJpJ96roPHuPr42fZ/pkojBLSdalt0D1V4Ex/e5K1QZSbRXQKcWw+BGmdkA
i5wyLF6rxS4H3CWfzOeXK9+mqVMl8mIYm0j6F96b/zRPOyONqK2IdGClTY9TQdMj
NKcJdQ81EKWD3PVZUtlch/KlgCz5gStg6r5c2H5wd6doRTy1VFrNhCKIGNZHvFCC
VTk9ugU7PD7qN5Du8HG8Ox962Qpr6ztCul83mkuXIn08q0AKo7Q1xPNRjrnGRhum
RmEkHfb8SOwbsOi8gm0tG8kwDHukjcVzjvFtK+hEKQhnemKDQPsfSbk4NUoWSnda
PheFI7Sqz5ryjagNgcnsUzvKgehgXWm330mxB3n+1FbzuV8EPkEAi6AWN22bo2Co
rEn4DXmlZ4BQ1cOL/PdofIdAjYUr/gxFRNm9IeygMxYglgGJa8iOuNQVrKyvdCpu
cLa1Z/BVk80ioMOe7Xpjbxjckx/K/jGhyh+ArutVNIa7r0UwGIVT3rGBhMlAVVcL
cmkFZB1iJbVTpbd5x7aWJg1UQYhfhYZAt2cDOW/dS6QYlBrX24pMWfgQfimKpIWk
laoc1VZnXqijMdIPGvW4nV+OpJkmmGz+Pu3va2bwpdvQQ4J5UgB+OxJEtZPeUGxQ
Acahn0UmLcKeGE0zxHPIy5O9xBls9slmObS2KkdoEpKb6oWtupIPyfQOzEoz0yCH
WKYsa3juqV01zwdmZg4noqK9LAJM1nNlbYtWrvQdnH3swK7oxhDRjFcA0k69ERgz
bwZleW+CgeLjVJrYpDFldxS672yyyO8Tw7NFoRcGBpOtvy3kTsFSjUUfJSGdRkvZ
891dV8RWAqdLb3770NfrwUkS9m5mL7FRgtlnIXO8gSSYKxOsL5fAEUrRaPfHTaA7
v3kZdWoYfG4/XKUj0sr/+92FJq0dSzvJCfIhmbjnNFeLD35IQvcf8ZC2Yw0fnaZQ
ty5XMln9VgDxFy21sToJzArom84t05mV8ktpL6k8ooTQ7mILdKHz3LY7mEk/Nd6Z
F+NLUS7rDXODLuEfrA6XCL9aZnEOOVVXG+tUFBruJTrTQMY2NpLMP5b2NnqJuqyh
/9ip5SDu3YMR+AzvcuI0gv+Fhjs1ncxY2sKVlUjHyRadufxCrgLrXcFtGiQh/haz
7GUPw+35TsEXyd2fRLds3J1C1FdFtkmG2UOxUTR1V9uJL8by1oLGVuiQR0smxEv4
RPDWgLAehy432o4gmw4LOGvY9qzjFWdzcyNyTZQlT+bWBxgVtHtltB1EgAZiyj5E
WKmIN4v+3KDS+rR85+oZCZ2XjjoymvGyUtGhX6Fhvv/B7LPo6ChjOf+4psFKzR60
OLrIlg+WuKjGZ8X1ITEw7kBX+soJJm9vqbMKY78LkwSzE4mNqK3zD6P0z9GMRrDx
jAKgSvMCAid9F/DjHcS0IqPnrDw88gw2tUvhttEyueM28x5dmjxljAjzCd4/rUPb
vXF7Q4fmLdJTdyyEL0OP6mMcmyiN968qFoTZL93YfhBDzp5S0g9R/rmJMalsd+Iz
R6sKbStm1wMMxZa5k1eflrSPJT7LYRtGvYsgtGvkparwYJGMQ4cLUHiSH5ves7Wc
3R6A4fRk3+imzCwI7V+47CwoUu1W1VUF0erjIPGkCy4NZeUSMf4aLi1wU6OPshKG
0wqzRICoykibPScsK6q4WD66kAMWp46bDtzMP5Xm3RU9QOIzqXf5i+0GTamYDwXm
Un2sAbJL6L21Bod4Evj2mJDtgfD/t91PJeneM0jUJHua1efskRK7tqjYub5+wFiI
d0bT7WyGq93wN7MaOfu9q6FXmNUxGF9uAVrTUGebtwbYV+6zqhPUoetWb+pSvNbq
B7KAwGP4zIg63KgAlpAhQNU2y4NlshT1oCIcHIBoyWBR8B/gNgWwUPD7ct/raKj6
6ki4t9hU8Jf+QSeFmTkb54fe5QiwkfrHD107Lf8QPgCat7oyb2dljCBR4GR9OJ1A
UWsHhQE4r1byQMpbK8wmJ1qtdm9FmcY4ucmro9IgXFA1CjAsVA8NsGgHqOGs2JD4
JtqovFSfKCOGb+HJYo/9rKyKPW2XkkgIERDQD6PPdaYwJh0N9hftrEqOxSmXDFda
4AWCDQQW44PD59BlSiMe1M9jdPehGSpZipiu1AdaAcml4DnuPmoOZSEkxfxRFRnr
jp1FGBA0vOChlpBm0u+qYtoq/cWcPBIHPzLJUpIoyPBaUzKtAjUAZJDUn4F/V+q4
Vb/JU3Fm4AlMwb9w2+sgukh7mVJzUcm2qug0J8+EzV3gQiZVPh7+Vqkr9pHKxGhx
L8wte4j1UaLkAU/hKB6u/7XsAiD/AM+5J15/MUKt4MhMX79yjJEq2nZi+QOjdYzG
DxAJ7EBFtfgxlc6J8qRMunT0qq5aqMVQ/SlAMzjWcZ2rfZdY4kCaCqTHlQBdnwx7
CcBK61YbCMfsu+UF6dAPdOZoLy0Ia3LKlGxr2KYRSbAvhDXcuKUizRZG1xvKIqRK
7z9bDvp6OJ+WOJER5/AEcyukubaX8JjxpIdznMoD9TKrn5uy5oGmdui5Vfu9hcrP
J1AYhMwSMvLHsfhmQ5bwz+qFD1hKB5dCXcClmj9Do6P97DENeKsJgKGs8YjRlzuU
kgv15HN7dg9tLlyZmOzk5EilQl7JE3+2igxe/VpggMVyxUgu+eH5a0bHZE4f0lhy
09z3ejCg5a6UEOWyg6dAlW+UMbWBTWZ1v9heIb5S8zysdj4wL+UrfSIz2kHM+1xx
c8doXp82vYbF4Nfc1/0git49T/X5AMLW+HRht8v5RFvmAGjCbYaJY5A5qGiw919Z
R4m7tWcu4LUkYWBsw5sGMrjWz8RSxvcTBSqRoT5Vjtym7ljwB3cqbszW6CXNe+yX
lHyk29//yNRkz5eM7jnVNsK4r52RatfabANFIY2u4tJH+5pzKd70NY7F1YL5H+bt
/Buh8Kydg9QYkmr8fVTohDJjXiwMR3CmWx+Hxt1ZCg3nCdOW21VkjCa/XtmF8hvL
O8U+kbgWTV7XRtwx5do+12ARi39aYQr9abuSg+syKaSkWesVaGmQmaOFbOiog7wu
j2gw6oPVSUEj/LUv/WipYWdjaR5Ckt+bC6XBHA/A7sRcHyOqv9ZZNcph5blKIdu/
2LpHkya9NzV4f/Hs13jrm2Ym/nUSuMkuBeY7I7ypNp+c12h6TT7HYKw5wIEv4ZS2
6sZr4o5rRLvluAUGACX9n6gejg0BCt0+2Wc5SPKyjDYbs9T3XAAgzKn4gIjRpoZ0
hsxdU18pTZFlGM5t/R/E5OTfeNSjJrDmMxFPspJN++Gwr1PjO4lBworPmBDysHih
Q2zYlKqpRd1Dv4K8C8knWDC9NsJiWfZQQ8utbaY+R2VYXP4IOHKCyCuLXfZGT+Mh
Ry/lHvohx9XVkETVVRCV5XRk3vTMGskEO/8LJ/iwng/tzE8Bhh/8uPC5zXDW0ZvD
t0YHyjW/VI4cPrZlcOhKXNGKszA7D7gktLGSzMz/CoeKehkOO9lUr8+maovmbbmd
2jvKzpo2XD209Tb0GL2fQ5aGv+nPMGYttarz8kB2wOOUOMj0vME/bn26HDNQK7jC
WSI3gJMqaiDJDytHjkhDvXPg8CT2r6yHEpTViqylj7I9AM6+VnyM4NyAIPgwdWqR
CYi5NepmIStTPK6xwywYQwtAKDtwh1IhT9SPAGqXOWqV5xDLQYGCziVhXs039tsD
M2pjstUorSoBziyH7rOIyuVT/IxjNSpBopOCzf3KIlYVQwPou6sx/wDoJeNSQw+g
DwjTX9xa1AyzERa6M9S3ez2KLnl2kyoSnvyhMI6j1won1LBhz/sQAZsQvh8Amg2o
gmgvxd+gEnJwGPRFOiXPzdJwsUj3/X84xca1YmmfNAWFwKVFhlR+1PiOTmQxmP/f
MfW8GbWxj9Bv7uOjVmiRxva7CvM4HWJ2Dhe3zHIqHMrVMwowWHqLwYAjD3QBjkcl
6dCRnNSuytm4fXdthbAiXrJZ14nZ27bD7gL1OR3HU0jw2V9r0LCqB6VoaMzknjqd
08Rp/lmVFMmpI26wIlrVPlvk40r3qBFW66UPRx7uUo7Qtfj5FHJkSgGMlGYm9SBf
SABLNDiRK7NEt1SV2WRlq8abq3b/P/HBNRLfRgKwLThA18uK8u/e4QpMKewE4ulW
BQIQ/uuh4nPHheCy+GVxlFVTdYBfuumlg7l4pgdS07cdJz9GOymLezZ9+25V48Yt
b70a0UBzYwq63G+DcTKuZ3YlnOeuqk3bQVdBoX4a2AZ7k6OMhKAuD25PdE1mixQe
70P3z2WLxTN90Ul7F/is6sM7hHOKrTstfbyzvfpM/K/sQGi3pbRFf5TMF7OYwlWx
AUONbraBwG7MZv+0v394oqPgQj/j+c119fAc+hR1WaRYifd78zPHgoBZBKA6Vu+E
oYQr84ID+geulAqYOhQBmRK0rRXyZC2GC2rdRzQaS15F7M1ODEKfU4ryaYWaUodl
Prgs9OVzIVtNmSYx//kDMZTPyc5xW/kMVJVXQRbSW6Sl/cTHkTabpu0uEb3pjy9+
3Zuy9cjUUl310a40xUgYRlsxV2PJEVxLDFe7ZgSvb98vWORFGIX0Nynd7ynsRR57
6SaW3YQfQ4hdQHysu0mMBdevWOLPUAa6/JPWZ2zmat8gSmV4pk8iMNb61QKeKH+0
tW0t7GKVlsLvjyjVHug5nlE1NI3He33yta8ie7Iiesv7Xe7z/sZdKGpCQQR22lCH
wxzrkt2zzoqkwk+HX52NaS9prMPhySS4M9ADTR43uiBfFEYxvfL41CgHb/etDkRe
ZtPs3tm3VYLePi4wWjdGR7UrbiZBmSdnH7+2wkP6H0A9IpzONSUMSnh9MtElshdP
QZAnrMPT/xawjx1LGLb7E2qP5L0IR2CuITh3OaNrF6NARdFiSqZ2oETtDwinLKHV
Ayh7dfKNcryh6m8Aa2hc+0gXzmDtKcBvbl8tt3MHHdCHGcImwrX4yzBSsUx4jNnh
/OUM1thZLFLWGKoxeqMfKh9wQLvtgaGnCxJhByBIrkkcnKEe1wdVoE57rTxYvOU3
at7I44TxAYkR1Fjrv2yVcFSR/k96ri9YU3UDGtXQ13ivIQOtfLBI7UYHIndjBw2c
jzYOdFMNgx/cla//AOr/Y1IyzlnnV5CexBRtciwVXqz7BXcCmaS3MvL9Rpwd4W61
SI5dwz6UAVn5fIrU6QdxiJIk6jwZF+vjyXeOizX/9A8p4atLgjc6tsaUnmUt7SgG
sRLQvqFPBzUy51Pyqg1492DOTOFRbb3otieIVZe969F/qKSuX1+rJB/H1vpCPOVP
tSY1fXgBGAx/cC0xHRiI5jJ1NulQtAETUq00r57q0Mi5rOq0Aw4tJLRVL0Cgn8IF
7Os6CoJ19qeHtI2IaKz2DyptDWkweQgEaRT2DGvo7DCplkUobH+53cRvKrh+0rhb
K1Vb4MTlmZeJKqkD0Ugh+mQC41K+w6oFJHq0NyaPFReym4lBKrQF3lbHCgkWLUg/
tzRfAeqIDgsplmth/M0Y9ghz5bTfKXkbmKIT1CgDeVp8IB034VVzcR8xVtZ9rtkM
WpCsegG/yrMr81PIViD8fRgkoapEGfRz1KO68n18FJblBqQFQU/fabIuzs2z3QEe
0n+AO03SmoBBFQvoDOwfwbZArh3m9Wilmc1HHuhANg4mlWPtzg3aGSYUJqeWrXS4
9XZ6jMlTZgymTH5ieOp60p0BIJ4Cyy4xxy8u4ODJy4RbWkvJrKHV2ugEj8/SZodi
/Ksh7Itq9AFtJ099mNmAdhvvLM+vgpWrQNb92orgxq4R+Vryj4VZ3DNsrMVZXSNS
rxATEJIM8dsTfY2BWWzq64I8p9aDTRMaSGP+KlymDxT5SgrP7T7/uCnbn7cYI1ok
kD4U62VdqLpX/CkyFSSK/nWlN0c9PceXYwQsA4fqZTFw4CrUYzx4FtfPBcpV9q6t
4ta9fjAhKwpcI9kkdg2AJDhRbiiuYigIoLkm7sujCOF3Tkb/IfMhhZYWlVYwCVCB
MtF/rbTVhrGjJjgNNGCnlqDeGD3fn25rDe76nDLI4Gg9bZOpsurLKdiRRr7rNtEb
SQACn3wfTKG1nbJI0XE+rcy+fPg1ymhNGGsAxslM7b4jgSbE5R3Kg3nZoKlX26Uf
oU/UHNUARFif83veeNc6jrtyccaLY+Wp8dId61ZckHtkSD0bn4a2IaxkFzqAOytu
aaPMkDX7eAeINmfXmSamb4uXGBOVWBExTrMZQRD7vNC0KCnlqkioamgG3MEFfLu4
WzD8vAKKP5zA5BTtAfwOd9aIRUrQHzklEDzeklblrj3xDHm7+EUQxfpClqOoAvjP
D3ZxBOuYI2+pTfutvvGtEBd86a7BGJTDjHjenLmVyH6UjYs6bNef4sz4rpIWbozG
tYH8D3WQg4hMvVoMDt0Vr2UWpANcx4WqBV7GNWWkI8mA4hQpylW8vzts7BCa5mq+
sDPi3AWxUZHO75alW+yC6Rsny8MkqNIYotSY0Z0vJymvg/jyrrd/C4JmXAxTuekf
/I4GcFmA1JOEi/gj53K3HCGq+VQu1IZWQE6fTE5i8WvHZ3Nv2snIY0DXVK7yoB3T
NxjPcajHkv66NmcjPrructlg/wrVE8kfHMy569g7C8LbkTj3VJhshb9DtOUnjhL8
mPrYcfhMTyAhZXgVG4L+InQxNuLG4KofY49Qchvx/Mygzw/fgeoNzGwjEQm7psGO
hZndQ6H/P5VH50+YLIhfBJo4EtdfkFqzr5AUzEcYMAnaw094Uqsb8CxWAEHzyTHT
HGGOjiDXye/WzFSIfW1LKETW31YUKNoGMVHhXR332kKF4DXg6cbzgC6BhsZENh+z
1bW93MlqNJO0uRt/9ArpX6jV5NUfwJwTQGqSTwJanwuwGMKNNG0YnY91wGPzFPaa
3bLnmG+QOvjHAr6fcCMg4tPoGZW18Jr9kIN6t33VkqWZdAapmLh0lVs5kTfw0MbG
fqXucL0VadHCGtwxSgJr6uw1fGanoYF1RPCs2bzfnWU+8Q80BRI7SeWe/ciyg2TF
hOx+xd8pcmuuJVMf2lB5VSz00SV/U2QU5Ok3hMCA65yL0sa47vjFY5J63id/k2a5
2g8MKGE462FeLDNG/Yr+XVZvmYGFTsiCm5yqGo0esTexNjv5v3MM2yEMdrxpLcqX
D4J4UC4b4dg+iRqsHP0G8AHCnmYzm2mk+VSS1hoNKkgYFQbW2eyXWD4wkzT1db3x
Ur5W8a0hsB0XabM9ysqmvf5AyKJfaOU60H54M1qFOAGU7kLYY817KQvx2+CRe3GL
5uTvRCSGPlqwG5Tf/GzjIksbKqfxjZQ5OHv6mBezzCFzhrNh/2Xu31ZbCVbQoR49
1tNkI74XgiSgsbi8QUYk8nAVUaQkcnyeYxnxZolFanYv9U88QIUIJJkm9ScFtFNE
X3GUVnFJu7N7BTn6AICZDa7zGhJtbd/DtYoRdLAKT9BLGwaw/mLqqFmge0nWDVAT
3y5UfDgPgOLbvX87M0kuoUqnHjJxLIeaVGiY1V67D7kGtoMbSbRAhVzvS3cpBmVQ
x0t4TEph8IMeKE2UhFLGi69qElZR1ng6hHursmKLSNUDpjLd3haVLjHcnwZD5BZ5
rLVD4TI8H9MJV5Hy6tLrbw5RNMJsbpxIDQ1HI9xbwbQfCyh9w5iHoVJRsMeEhs2r
GVVB75IFnJ/Zv5kVwcHUbUYHvlvodrmoqMb5TxmMVJb3r0Kwzzsb5jduE02qv0k7
KNVKCt+fV5avEO5SbEczChvl3kj0oBcf/6IllTvO/MxHmSr3oa6ynjiMHDNqi4Fm
Zd5TYDq+rAjDFhctO0eD1bdCFP/JpI17opn1grV3Ul5OsWULG+/zGoRBkyLYQT/u
nBpqC+F6SaFMTWxQCmehxGopeDyr8ur+kbP4PqvO1kT+X3sx/307hKQAD2HAsc65
1eM4mU683JJLpenAPaAlIfZhc9sWKk04p+IOIvk0gwGPxr/JUieXR7J/2js0XUJ6
dZCCFN2Rl3EV0ilJ47VNg4JRcUKIpCUEpKT3CQtXol8pw9M33iFufJ//ayhlHclv
w20EjLcooo5yw3mIZTtERj+Rc5FSR5qizcA8VrQKZjQ1Am2AFLnDjoXkfVRFdYgG
S144Rg+CQhUiBxoJzOBQvz3ERpKMZSGT9YPiZuCFzFWb2ipZ5+Gn1IrRG1F6Py+S
aRyIcFhl+xg9J++4FJ8diYkmUjvHeCCicT7E2riQ+hvE4IVbIENtuSTeKaoJ6/Ca
m4ekPlC10XHdChS97m1FW5fT0rZHoe0lV1aIbFZrBIrFbbW+vDktXI5YlLTtJMYQ
U3bCYuo9dGCCketQC/BR+HJF1C67WzUR30wHMeEjBIKuNmgdu2ojKa566ySjiM/B
Msc9TKdNcN1oft8128CiTkLbBYquS/13eNT77OmDxzY8FQ6P2hwL4RT13zxnmNY+
RcgqAGzfFJCGX63Ix6PJNwoxnq6VzHvrtvhU5D7OFnaQ0kb9zTONakRzBgm/ZR7v
rOotGMZK17vUDs4dY7flGs24U9Hg06UTEgLe9SGR5MHFI6Lac9x6GzfeYDjOTCir
r1WU+en4paB3/5mvPojXSz+q300oau2cRNO+iCLqP/VohMhNPzpqlrXB3uLm5qVY
EyHK5LyHtDSqiAHRRR58cTM2NEaponUSDla2dukmJHn+ZVIU0e0wAfkD/q9e5YNC
pCn35e6bl8iHDZYruxXa+lCqdIwbRmj75nx2w2Tfp0yFMiXQVqsqM6HCq/FuS+XS
hVDp+u/FbYS8dycY7GvSquXG+qhqZtGtVKFbIIgoYh2kCxrHHnIaHisffoLnsx3x
p3RnEU2MmpbXQMqiNX6jaSWRNkhMaVglSpIQsXLXcELDPysqwYXxlRIq0a9tKhf8
fQ9WPazekXrF1JObMvRNbXglqmMOSsZb7jyzkA+e9kTF8ertjhrTEpUeq0jZmvvs
Rn+rmkUpA9M7JIJr+z1t71Ga8ntgECYCigo99OYl+kfgse24kYbP9yl61oLwYO/M
mN8Jb3tzRBVayvp5v1CVyXQcu27VOI5s5LgqkstBvjBqqbVqjxylwK2vuRcGoTY+
F/c6EK8fN//HbGyjdfSV+XNXQQTK2zvPXzGX2apn8zqXUuZKCjOFILBSdmR6d87i
9AdvUsSq3NYgDob2VKSrMC6rJ8QHjJ6vEis2WQZ5iR2FYRQHmaTzy8JAj7Q159BK
J8ekG/VhHgX06DDkQSPyZxAsr4PjuPDjlrkDh8lO2bFrRZtZPmVGrTYVfhOf44F3
6YxvVdR7YmSAkab2Azt8RWDiD4F9LJn4fl39+5UfOiAkGMz2HECMgS9mBv/MqU53
IH7HXHsO0USJ+jN0wpw/9EDrQtW6BZQlaC5dFvUaoSP/nyTiuDMgEs/L/EsmNSH/
a6HvnV6hyjygJfeOv0oGDoynGyoay+NtySnyJp5NfV1qUFI4AF2afYBRXStJ8jnS
Dj4jIGzKlUP9ZVHl2DHnr20qOvinORJscylclyatL8fJnk0Saow7jFf8R+iuBzJO
MCAed1meqZuuz9xFqJsbnw5VDMQC33M25u+FI5GgKul6KnbyBEz2pbJmnRRy0KKF
Ov0TaXDqq+7Jqj4aTPWnT946aKlJVer7eChHm119jFyn5ElAwkC+HZLYPIcjLwod
RvB3SkTx3KJ5DicbAaiFQoiWgjikcD+/T6gyuy5TfwHgVTjrrH9OmuVrjf8aI1GO
z4piBNJHd4TJ+4JZSQoZpk6mftlrP4Et++q5EhWUt3xABCLwmHIjMFKWREuFKsst
gdXs20qp1pqG7HHKZEbxBOpl10DXjFyVef0h2sADPe3kL1/NLHlfLzE2LImDawWi
xuKKsZS3WgVkgVH3vLumqYGOQhCT+ppEWICVlkCe+Ljwi/76Nwtbysa6b2HsA5eE
fMYv4WgiIUNxS/7LD7N+LZbr5Gykb38HVfMXiEtdAYmd4ZfLGkbmGoZ2dZsyaioH
AHtp042axrk42eCZaAyRbJE5mMKcqE42PGdTveNXaAZA+kjTJkEJoX4BhpJD5urp
0nAXTpmJDRgKUuQ4M4iFqjJWAwHWpzBz8kIcMp+qGaCqWowHCYJVzTC7LEZYxwsk
1Bb0Rzxe1RNSLAUycWu3Gd+vCkyjgnmD1GqMfJjNc1pF2UnWLWMv1voPVMzNhwNk
XZIH9rH+mlIBsT209sQl8iiBdgo6aLn3O4nX7faGTP1pqk04Hfk+hourAAscWxoi
1aLCfGik3kinIu74dzc+v6wSZfBEO6f86044uL9WMcJhnvaCKCfgdrUrkzIS0HHi
KkOr6yQJZoZ9hU2n3I+n3Tx+aDNWNXDfJSwSwzWWhfeO0OISWJtsEjDLCZoOU0Ut
B4Usp8ty4NIKSSdllnEe2/169hb60X6T9dIM69heDB55z1joiisZ7HQo2spq0bnf
d7iPpF/KGD2f2kjzfqVvd9pOMc0WTaDHMNE8pCGb+jsVzb+b9rfPQf95ONbtNNog
xUebPNVxX+KJc7bD7ZqyIHfCZK41avIOoLkZ9vL83bFEo0kqQdTaTiel0+kHQPO4
dKXwpia9F5HNSiLfxCMig3vwY4itVt+XHgLTO+AigAxd8CIDZljGZhZfp9LkCdFx
NtnfPiSc+isq/iepBkdk1WwfzshZ/VjNHHqGmD28EPj2UrUZscfmShfLRVhUzETL
FJ2jKBOim/eYuphxWHW8fp0o9TA7CQa8kSxakLhYgEORxcrOIuFe3ObFD5FKxQHH
iTTrCXJSzbAg8kavg3rvi250yIxgeQ0/9ZeDQ+EdG1qD3FN7slcLKor+xvriL+SO
W2VUcSn2X0cFT3CBCAbTM8JFJvUKyYe23U3t6Ovy99tc955Qe843GMfEO2fYcHYp
4uKphOu/dJSS8LL2i8gj5iEr3hx+I5hSI5rBkhTKABaAQM6VHXyYrPP7rGN+Wh9b
xzkwcbwfpFOcwHzaswk3WMJW7zW1NSW76I+4CFAp/l+2yd0a3pUvbS+suT8yvxW+
bY9HhMTN/N9KGalE93wW3uSwG1ERncKZHT4jQVyePmZn/b/RGEzLVt7mgAfM8gyQ
OfYd2fImUlbuAYN5FjXaR0FYBJ/t1HcrPR/p8B7H/H7tAFjfFuknUkC5a1E1VXpJ
i0HZN99qzaudolzijaPTb+dafvlEOsr06RsW+l7G0rKPzwQWeZ06HxFAi0rElAox
gu3kaqdVR/d/OoRF4J2dw++1bTuju3S7tK84kBMmdOIWmHOn59cRg9fj/0vd+0Q8
gQLDkloXogsL6FY84tosTWE3FI6Rhx4Z2nq1lXxPn+sd+QpQQ0ckiMg77DL86ygK
6pKMhXpf75ga/W5EuVMG/JfVuvDGxwhVHszPcUZaDNa89XJn0QvNypBbMdabhMSj
nGmO7zzNuRzmLLTxCUiKKaMtSRlX0oPtN+kD79DS+o8vZ/EDZl1gj+1YpH437KrM
5O1RCchAsIrqV2rStMzrI+17R+xcotadMiheW6I+TetK9JknmC4FNiKMVH/D4DmO
CcelAYy1N8WBx4fbr2R1Ml5DYT/RTrEGvS8BFjWLTn/qd61+bmGQxXD/Odij+MyP
cJWKVhAiq4FkYogNe1cB/Nbr2j5vAgOMWURjE2YDnzWhXREeMDLLkNFMcoRLaX35
tLyBDEhXqK4sB1uMF2PdORf/iGc4u+M0rgaWpzCrIM3mLul9LmSC2q2TgKi6KdpK
xepvu6GV7bT/fpk9YDv1ob3lbi1BELXUzHJbkW6j5MyS+LZK/6kblivVclA7wSke
2XcXHLRUS6Q173Sfk/RlI0jNnddSDtyxsxqlhEDlCK33zBZ/Xnd1pyi5BK3ugAdI
L6K3a7tOAo7PAzIbdI8oeKXfqen+A6nXEAripn+Wu5ICRvsh5eKQ3/HvX9xr4O2u
AmffqMqVg3mnhPT82yBNWY47yUA0XEL8DUQarYRDjR9/NG2+XsnqPncjQ83XljpK
K44p9+v1fUK39oA2KZf0yAJgaHm9F0bb6eoPcu/MdYNxdw+hyCYhY5L6FVyNHuXG
vVhuQj97t/QI6I/wPRAprR/KHMRoLEhoQl9Hw1bWMHcbRdtqLu0u+Ef5geiuyX4t
gLDJVODGbBtMmcepiKx45dXlSgSaEaXTVmMuUAbHEwtF9C/Mk85uGHCZH8DGSpT3
QRcuAZ6YbGPms3RfmRq9YIzkR/fA7VVzbbCpf2C5XGaIaRjg07zLBZ47vc3R1L+i
0KftfvWpiLcqQ0DYWjrxn3ogBpnPKDmyFCCnQLWoqyhFbXYmdGK+hqgOw3WN5zGW
6qTMjzT8fa1jMPG1dkjODV+sji90u1WpaGh2BI5FhR8LYi5vwML0y++/tE2L6Jq2
TvIfdmayAfsSNxxlUEO8kFxOMrzQYlDZGYMySorZl9Up6Uu7lSJqqkCI29vjEt04
i5OHUzUmDk2d7R8ZojSQHJouZBT8nEBOow7t5UbqTeJ197ToM/Ax+nSU1KnKcu1j
+O90pdnqREil7z6CiegFzET6424Osu3Ml+GnQRkdYFrQQCUe6mpgyc7o8R+HilLV
BjG36u1uVx3Pb96j94/VOGlC31ySrjQ0qnNJUwfS8vRnol6BUvdZ0Qttr7n7zy/R
2HnC19jKiytcl8SRL2KaDb6MOiGq0/2nbVRjTzMw/bYLdNytdnOiNejwyt6zz04g
DCG7BPTFTYvpndmzSfVAREAxfjHMNU9pyb2v3JIZ/ijeJUN2Yhe7DRMC8GJqca14
mQ+BQuWoBbDPAew9zlU3f3Vku87S3W6zHGUOwhRxFEMhoGDWe1pO3ogTAQ7j4sgW
pKcSuNngG0F/RCIeNR4KrUEr5pqsMR3jFD6Iv97N4ilXtEbM8yDKtBzGl4BG7h4z
QW01aJ5YiI8iDYdL7z1ATfi+mB7KBkdH9jStjgKexwMv+9yBLVaFVqMhrc+ptYgV
RezHmBA10u1lC/ZVR7mQji7lEqUGO1YTRVZnrAP8UzZUr7xpdJo7BknkjQXXLXbk
CFcAGZRGy8zPbj9a6sBC1fqnZw0/labhTt6ANAsVWaV3RXGUETVI0ywn6ruo8Hm8
OUpK7OmII4n9R8l+vUuVP11EPl5SRdWmjKpTuL/LHeD1KckCYVxw8S4f41L4lGHP
VxMvULxuDHS6ApMbWo0wTrpqkkaRkKjdNtJfN3AwDHjbwxrwK9tPKkJZMSYrR8RN
vfcW5Nh7cDSTRFUZL30NMztnm9HRXG5/s3ihSWimMCpFycdm8UDEy1F3nJHSFGrv
wvza5N10uB2nu2ptcx6JcxzjvNcTfeL3Qka0KbrPeNGFY3tlcJoWqhsQQeesWScJ
f4BDbcZiftMPsAR85Zb+9zrt0wyOJt7iNVdsuCkG8MqSm2jPHlkISOHwOtAB0A68
JMY2l6Bci5cBTX26/o3ZPpc6WIOhPZrqTFHYjRkjb7NLOeqCq5E4Mz59RPJXvcUH
FwRxirVb/wUZohMUV3nfY2QvIa/ARIqpQ9STboSvdUOErGJixmStqoyMOrgo7w0Y
U6/ezwCgLRmC8Uysv74/TGHvyIN4tZ2yWQuC6DWpffL8SiqXdofqUaFv6qOfckz1
Ib1lf9j5x8ICGWD7rNR1jUvXa0Kj2cy08uEWl3xud5U3idEC/+J2eoMsaarf81G3
iX/lnJiPyYesAq2EX8HY3mAKVionztMjqIFBwI3HxPPrAFyyszeh1JyizeffTxVn
N96LQjWth7ovQuVjKLKuMsopzDTk4gOg8hHq80gd0I0NfVDxtrT8duxsghjvFqCw
JFpgaqm3hC2N1VhfvYrHPiey56aBTiE3j0C6VdNW3S7pV34gqtb+JrY9R2a55VbR
vL7wfcpIHJ+GgB2ApqIO6BrcPoQFAJlwVPvoPbNBS+LDugDSk/Va1l+/0Jv/Pjbx
G7VbJYGlf6AF3+u+d+SlMBIrL0maUwnSsDVf76K4HuGzD6DkqcD7NzQpEGgsbW+k
bBmaGWVrKlDEuT2lyq3CdBpOFxPTYIOfR4L3UoDifrRle5zd8lUVBqP0gh/w1rQe
W7pz1wPyOaEtf37O7aBsa0HMpAdcfFFKC1fI7VwiWmp8SieUU6i3D+2Vmjlev/bq
+MOgePuaeMbgEmaf6P+XuwB0rlYFcHctwnHG0RlH9xv/2Dr2PMdxl7hXZ50QkWhN
bCixDan1y7rmzL3+SsSAtgi3k0ojV201OiVwRZfN6K0EmjQXcsKyxESpJVnfGs0O
FG4HDyM5EncS/c814/DhB02t/Nd32dbKEBymec2YdDgT8I2jtTA7FTEP+OCsZHyX
6+hoH/UCwzjXOVHIcEb10PdOKpw/uc7vjNcfCUT/HgysbPFQ/s3De/Oa0j82Uv9m
9Y9dNCnClg/832+a36Th3FmOhgpwfhUx2sz+Oksu5E+n4DvK24X53n7sc/U8K3zg
jBowll6gMLIXnOMQ2f7fB1tBJ/gLnlp0ikpthIxG5vV+J6BCXJ7ZUIFo1za+OrpB
i6Omi+ofydszbx/IZgavoH0uDa6eFmiBDhfhdaWJa4exkvUL0XN7ffDgBgdSSD7l
DSu43KEpgL3Q7Rn3XV1K3Qi678lPgu5zZHnCXzXY6u7pk72TND0/dQGoog1wzVEN
EbQYSLN+NPp4WX9pHV8hXWjrydUXEIfsnJHb8pJxZJXYv6N+bCFZv3NA5Eu9MAaB
Sbq8tyDlph6fo+lg/uifc4fyDJ5VXBsOotJRv++476TQ6b6TPzP5EBtiW6Oh0t3y
UpzjA0zkkPs/IZsFtb2FFwp0JaIWp/OSvatgU/8lLaBS1nkj46NYuSQ85iiJbOdV
j8QTrmimpLPRs5YeYlDteEs5vT7ygPjvLVFsqvDQ/1Uce5uXQyEx6GMnOxkwJLfG
fbO4o0VBPAnK045NU3Eu4oDiUmv7Wjkgf48fKmEpfY8ahM7VDus1HVodFts/lTBc
b5dhKG/LsOyLlkAdw+8Atl3RrjYM0mOaa964gW1dJlXE8pJqBnk1TmGyuVW+TBVX
j3IOvWHjfEQIIGv410OfH3LNQRO3Wcp7oXEDK8cJwtjQhRKCLCjkxrTar6RPcLUB
l0lBihW+sYYaxDyNRka9FsqA2sD37WIJUEBmKx38YmvxotEf20/4kJAltIc/fWo1
NEWA6KJp3Vv9+s8i6xJQMC3qARFrWQluEM0vORGBjFA0lXSiCFCMx1ytC4ZxngzT
H0eUYUrA2rV6CtTeSjjfbO6Hd/NtVZjrLeofYY+vLPG3ApizcX5KGTaDQqoZn93e
nWezWeI3zFu/d98YC2a1CS8Ks7751s2HNuUxlLNiUV/XjqwMAt8Oz4khrd1C+P/I
6LXtYdyS+wQLRsMzmZ2/AnjGIdZUl2J+52MI+Z1TLBhg6QSL+iuuQMs48f5IzaaQ
+E/8gKwhP40E93qfqhO1Vh5S5LafzjfDV986lTj/5RsnEUQu9n6qRYWzvQ8Pnmo0
FuLQGDHxAeN7tsqTTPIgrmqNm+7oukp0oUHEvxv8v0+PPdmetuSqHgXBpvnKINMB
k0BxG49vqfP+UMKKIa1VpD/nE6QcyLrYwTIbvDwpqUx72UO9TeHfnvy1K74vLHri
HDcbZQbk5o3s0awcJqHbQS1eNNmgeGyeylPaURS/AhDNfil55E3dkV+tArsyUo+a
oM5pY5sPBHcEXjUYVRJt4lzPrMpwLPNor/QMYZGhM1NDSqLlMIlhs48/sdnxlmV6
xRKy/XyTWBUgubL7M1VPKyhAJtrbG+NDtUX4ssDEi+1a/aUNk318a1V2YRa/HfMw
16csVqfxWEXH4POtdoWc5W/QudDn6zrbNppAdZzVf5tY9LRbk3Fqf/hrKYxwH1Xx
6PBIMgcQ/k6hWxq/qkWQHC1Mm4E9O6TUiEsIHMqcBodnX2+60Dn5t6+bB7tmlubC
yYtkntsKE+aOhR3Z/eU8nlzXdtHvfWwD1ITrD+NgWxJirYbImUYnynrWhxFMFfd3
CsG61NAQQ1djxOp7AOerYHmL3e8pxx4Pbu/h38lT/KXvirHFDe8BnFpRdS7bbLli
NVNw5lcX2razrKdMEigxO0fojTx086XjGXDQymrg6K6H1b899u2zeFHL9kj49aEC
I9JI89A/bXUbEfiRT4scwKP/BM6A1tETJVTZHpmKZjgOCKge25DfVbtj23IKS6B9
vT7FW+nMZbsUJ7TfwR7gmaElzHC+p4tqXPOFrA7BWLFF9/Sa5aSIJcFZYLVsY1DY
ig5EWjomtUTdqjUu2T9OtnC07QD+4abryqq1vjc+AYPcHcX9ld6DPP9VAIrjV4tX
vXcxMy5BQyqQOcdpQ+QIarJgBBo8SB4NgVH9/NG53KLBU/PmQNMZRUEhcSGfD/W/
4PhKnvCw/loyUdBWoBQIVEogPRSi52wF40FS3Id82yVNkqJe4Z6LwuJ6DqfOg7jq
amg7gpFPxP31jdggtekjW1AsjEuO46MVM1GQnUX21aLHHLydB75Q61Y9Ut8hvLzG
4cxQXxUNYXacdNxm9lw18suLN4hzhHR2iZ80E0yVFquQD+cvTQU9SDU8dr3c5WbJ
EfOuBPeGHAeXhfNYNVRdBi+yf50pfD21Ok4Rna87Qt2RM+FCHK/ZmGrPqRPNVyHY
tmv7aYtT5GfgiGA1M7+wDdx7wf8WJlBG1ndbkQy9NTmnTuwyVtWsBJutrXUOHO1z
aH3HuScnjONFYXUKhE3Uuy6Rr3MhvAKMBabWfy/R1WjrLsrCkq7RohduDdeaA9eB
X7+BsQ8NEJwNQqIQ5K5vdhqKtXQDrAvbI40pk1JQHQj/CN3I0NO7beGB1uRt/ORY
Y8I6vIM83obbYa4KPZlSlVEOw2JAfmqjFYnRW0BWBb6H1TEk4yPQp/MFlLg05jwz
l1o/99aSMkJFKV546dmB37wOlWE3ivdEXgOP80dQOuQIIJxm26bj03CJYvHzxjp5
FlVuCmakBAWtvZ9tWt2McR3ntE5vRsC65X3IlUkUGUOqrLNZcTEIbCCty3//rH6b
c7PuwWnGU5VS/eQqvIXUge+2zKK15oIsb5ftew5RdztjRkOr8KjZiw8f2NNqeyR9
sWu/W1W7CbF1lSYmWYZRT/5mkZZDyBllj/xT07qs5HkZFn4H5rbF5bhFv+3yIGy+
KWekXFI3ZabdSXzD87ArxlVEEcpLdgwWSPYjRm0WCdymu0vbIx+dRUMTHnfXUAui
yYazo6fabszb6IemoO5Ix1XajiAFISuTre0pjSIvxQ0vEnd6Usqqjtdr2kQTvMrQ
OVFf+ECuj24nNQqrT+VFGNCNegOc3BFTbHO29FDUJ7p2Xs8BXhfvvftY9Q2MV/Qx
jZWTJdDtSBjKaq3jRuAab9VcAOptmakYp+GF6jlYCmqkCLlaDHZx0Fty2Xn4DYP+
8zQJy+HzbyJQRNqw9h3bioj+/0SlY4UsaN+YNdMIXvVlQbgmo1SBuoc8uNSfuUSY
Ejdl3yREv7wOe3sseoZMXwATLdP80T2fClq9HhNC3rf1JfCs+WirDpzviMlBkEeI
nSRCCnEVLTSDYHeuVfL6fO4KK4cmkSoallQc4ZVbBtx3+rnBU1mdxbfMuzNS3i4w
PKebXs/ZW/B3T0Wqs+O2PE+HtjNMucOYO/C5GkXogD5L+vYiSt18pJP4n5iYknDb
0H2jWkgIet/HJdEq76G0lcwiR/IOu1f83rUtIOR2mu7WJlst0aYRnrZy3/Dc7H1B
dfcsCf2N798IUOEyFpbDD5FOrV2K/d2Ju/3T0rNe20vlop6tiKoecXMAbup1iIQa
4L13IDsHwfEA1DkeljK5fHCNKbo/KM/76VuzHe3yMOvD2G2p1xYnNimO4ekBEIKX
EQ9px1YLBgJsiSuiNuyivqBZ7TE1jZvXZ790DqGiIPj6fRh4KdkXfup90frXNI1z
fjcVPo0FDuzfWQEUhPS1Gh2DLM5Voy6OmQ6Pu6Dv01/LXaE7OeyOMnxZaQFWhB01
sGVztETuw3Fm68rWq4VULm6S9O9dRmh0ouYQYcnILzOf09PsxC7zpwOHNKTMThYW
YgTV4fBD0DG8B0aUW0JLfFsl/hYesIyUB24ubrZ7hz5BMpNfHAJqL8n6VbhvMvxY
bZQUbhMIpbcfp47+vqevAmgvKtaYmyqcqgY+XjUoIqXgwAOWlVcmlPkvYbCVMLai
YkEPWT27ekztpoUfv6FKN/RwJgtVa1c0I9roililP0VR8IQJCEiJlLnk5za8QVP8
BpQOKdUPIwzfytITSN7rWSkGtwC6qabYSglAG16NNVPeQKYpQtRDzfuhUBKKXLZ/
JA8zmhMVR2fjLjUmTr6lcNTEHqbJJgygfI1Uu/v7smGoIP++7LLweq2xGRdsjgln
XIEQBnLBNWHzBvE9Cd3vXLecVxN9jUCdXivpBuZn86fJDnJkX7KyJ+x/CetBl1Ux
gPvx1cKWT5Mm3t0ycQ8qIlO0Dyv7MrvR5M66a1nlzE327TUH5cvtel69ZBtmM7A2
jGDvEg3JjNa85RfeSj13+LGdOouT3OShgjSgpb17Y08jS7RroRTU2QI6lIO4ajlS
tKDWPBV8wawMpqjpdoUMMsJn2OXMJlrQUaSJ17SFdQLevIb8/KtBrl4oEYrd7klL
NcwIpr6c032W3vnlkq6GRtVE8rIevazsJYxiksfgxWS1GEDkuJrXZY9qh4nZ+m/q
0+VZnmc+3542CgzSPkb0na0pzodyTPQkJVCmxWd3AYrtzsrKR0FQUXPgGRQCTnL3
g2nD4b0ZPyLS/g88lW6/BysS7XyvKyZ/Kqsp2+v4EsLFI/7X21xDWUKaow2W5eea
2AZGXQcqnWD+bHWi6noAMwFsNCZYaXSOzCLDZ9qJRYScYdmoy0aF8pqwmG4n9Y4r
tnP9mAqpOxhnmngwOVxIa/MNbgIP0Ocr7RvmsHiwC1WJedC8grGjNlYK30FPHJio
E9NY7dQp2MAQqnaV76d1dWB57yLh4+TFy8CKyH76sULjHV1gnsEci9WXo/3b640z
tTFq8i1+WIf4ZGyHWb4r1sWPeHk4nacJr9d1v8KJFLbADQHp15+qCu3C8NLK+ICb
lZo8uxLpQLP6t1PDD3QI5MRAUxqPNnq0QD0nIj0p2pDFcLA2ewipYYo/drfMyxJP
IrLF/4nWDvNdVzi88FxO2XDomGsHuKsFk5GMpudEBZRy7cBX+0qdAc9BVKG7mGuG
dOkv46cLG0LErWsijR/OHFTtW6Ah8JZ4otQ2CpIiSdW0wPzJO3MMicVV9XWW5ukw
kh6JFS1bFBQkJEH4GgD5FqAm6yIHB7r2NRaSCflC2O8M+7VskHre50JwdSmNvSjh
HY6r7TQyKPEwnKSWwXr6iceUiJY1sKNvqmCGs3mP1j21KSX7gY/RT9JdoD4IrP4k
v72/D8SDlwYMsGtoFQArmyTR+xPXQSz2Jc1LHKgoL0inCZj00G/rKOLUNS6r34VX
UolN+AbFWOQpnimulugZ6ZWzYC8YNlG28rIQ/ZVvHa5j9VfBhMWpHVLN/P58oC2s
VgQu3ybQwiwA61V92MmCCHzq5/o95BewGox4rwkLkmgKf9CLMGwNkZ9+3IL4iYrs
A4Xt3YC7k2t8oZekQeXL7apVMr+6IwIHpBRMRR9XldFLh32LIQhBnhZQdcPj4KIZ
qeOL4Q0RWaM4K96XEYRN21oVbd5ZM1ShEb2h0OP1x/rOpR8Vq1cZtU1FBG16Br9A
ehm8LyfoqU8ZSeYt2eM15lZMHo5P23MuzK0ORIsIDP+eKdeyx1vXDUcOx0dYbnVM
ozGIw+RJ/gwt7WDY+juB+mLA+gsDPmVmKksfMxMwau+Ktqqrvnxk+PLgNpv4Okbr
W6d0IhXGOtzMsMoGlwIepYeoiaY8bz7PfgoSV5No/hEVy9U3zl66g4gNqB7810XD
A1ac6iF0kGHHCZRya4R9Jo+mTbEOrlEd5K/uiW6/oyoHrpNylcrc3oC3awl3LumE
qT1QIYq7t/KLoevZz/diRSwUVX8iRWORgUF9IAGjzUa4FC7vO+ngQZHd/0rZT7Iu
O4sf87aBfNRsWBcBXdOEASsRS1kvkzmynMutY3PXyjYZnZ8y34zRD5geSgiluYlL
uGQoYLjNPBvPrtZ33dseBCeT0qEo8DI84pUzZuovNUmxfjt8XyqvVqd7MzN/0i4m
lZME2qxY8TCvDaTIm2E6QYGzWs7qK/iXFi344u51Nj7y0huYNJEGHT+eoAfuHdpZ
i9PtGp5e7chbURdgTZuwUnBWAV6fBnxtk5HpKijiirzi6rFfDZ3ENqgo6cKk857J
wBgcs+zCVDpEi87dmTx5FNmiP2VT1C3XZhV0Kg4Foa1CRmDK+DP7f160SDhzFr+f
h+f8NYDjWefNuDHJLA4N2LqHJVnLmHFDkM8tdHpcmvuRcbld7Z293QJwqkTv1dvp
khBRwf92gSnYNVMR4WAKWJb/gMse+O4IAopMv7x31hEmF4gFk4MgESxnxQTRGHXe
6D7WNicpcL6R38I3lu25azYcfwp8gCXwiv8xTkmYUQzXfyw+q6oafzNzrZtCg2CA
QhqK2eo2Oh2eFK46RMg50WI1ESJJH4x5R7Mj2SHJC9ErVA+2NBIokInk2Zg1tcPK
27quqILBTT7NrBCE4KVQHDp5oz/tYN+m4bEY+l6t0mtkMKWu/sY9ujg5FCdijLQr
PgnCgb/XvqqMjGZZnttOn9P+HSYMxbs1x6K32vzL0XMqJZ8BJx9pTjqCx1mc78X1
2A+l9Pxu5HoXXGdK0874o4yjtqak94vOLnHr6TA+5z6IMrQ+51DHWTKT5CSxDo8p
37ecbaRHjSV2rlBLY8+jqzSIzSsQf2y9VFzr7Cbjd9/U99MxmauXX8guoqN7R3Jz
/x7sKfu3zD4GqRlUILOsv0ZY6CSLziLoytCuosvYOiMXx0xpew1mqPhMRZQuN983
pqL31Tt87XvTqnXRNjQpxbHMQs6rc4UOPUZkQnpzmm9rO2TN0EF2sE/zUzd9zDuZ
15KHhxFVFsHw+BkY1Lz6ZYWKonIN5Z+I2dw9G7zsZXbunPgj1aUZ8Xbqwf1u5TvL
DIXCnlaTato9VELp9Ej+1qhzUWMbpcmKh5iK4QJTn8L82oI1bSCJuBssGjpt6wdP
puHIupRhU4VTPwTu50AO6Hhl6sioDo1dXJ8hTfeRh/1EqLTKzPTsuaveLNGqN473
nhdePJrjGXORsO/tiWhXzZ7MozJxR5ZajEoL7zunCluFQfKEqlKbY/l25g9xMGbK
ZDrRm3ctvSibHHk2s82yyoz+/N55+m+o6gEB22FKmPKDuPjRu0ZCeQS8DXyaSvtj
/nFT1LQmxbPZeTpjrlJJGhC3tOEhzB+FIcdvGiDOUygLvjl4b5D4jfpf/DBSaQ9N
VMN6CCE5oh9h/U9cQxg/aatqtF01CM2ZjQ4Ai/D2/KVeVBT9R3/opShi6fBFYQxs
wXQsWVF19oIaM3qcY9vlBjzGchLBYk0f6UfBzfsoRNU+XLiVhZ5LyfF2f4ugz1SR
n3Y3VHwgMii29nVd2OfIibt3gmDrL3NyNzvrV2Auor5BF1EAleOMEvIuPCPyRFJO
6CEDBTXrM1qOpP23u4CvYiNZXspYyaGDjFlwRDsHqRguc7amn/JSr/eiWShx+ehM
N0VaNB+73ENFTFI6DszS0GtWywwzz1CdYnvJ5ec1t4RyPjg4VIu8gKRUny6CxWu/
pO7PKomVi0u1xvCdlkJXQr14OnVT182Tf2Iux2ncoLkUaIOUZ4Qw6B0aPa85Y7io
4nGjl6CqoBbr9Pq3VTSzVA==
`pragma protect end_protected
