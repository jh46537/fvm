��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\Z�;�j�A�r��'��+�8��A
��[��j�'=X�+V��F���Y�����ɞWV�/���ǚ!IVUA���>�W�ŷ@U�d����aU����Y�|��on�)�b��	I�נ�K���2�P,��M�����ښp���L��PY��㔶��i�,�Y<�YQ\�6B�S%qvc���L�品�ry�?[\|O�r�ߑX�Ċ�n�v�ƉX��,�k��L����(�����xZb�Ur�@�������5P�؊�1$F���Y����hpb�]���"��?ORS�i����M_�c����`�	�1n���Y��+s �^��n7ָ��BR��D����a�ʥW�I��/w/��.�%ќ	wY4��7�@���i����l���q��]��9� xR��ڼ̸��f��'hڡ3	���W<T{�}N��� �i�Ŵ��k5f�wd�Z�re�0s	'���L ٍ0�@�s�P�B8d���K%#�����1���_�U���?��J�WB��tk��5� �j�Л��2R�� ���m�|�lVD��Q�ۇQ;/`,�O��h\����$���m����!�T#�E'h
�H�t0����~ŌoB�M��Z�L�p7��[��ra��V�}�6�rO������n�?�U��W�'�����&8���Ⱦ{\O������A3�No���P]B��F�Ұ
������!z�s�1�kBQE�u�	��(:�p�N���c�e���mvh��Ft
�/��vϘR���0R��;v!R`���~؎kHҹ��.�ʙ���޾UJ)5�ׅs_sX^��7��e�w��9�4~��0��8�mh_d>>��0S��+]sH8�8��珴�|���Dծ|�xleҲ�߰Q�ɝ� ����`�����8���� �q�>$6H�ʘ���
Ԗ��ϦcZ��%~�/ �������|S`����J��J�T�:�xS�lɇ����E�o��N�*R{_`J/��ޟW/$����DTz+�B(i���Y��Վ��&�)C�F��K~�#Äh;�d�Z0�Z̤Ss�N	����N�T��.Ӎgi��9"�YO�Ȭ�-����!oأ1k�&:X=_q&!d3c�\��#�����I�)�I�J��LQ��5�n�M,��3]��< ��>�	^�qr����
���124�-;%�����ڬr륫*�'�y�Uы�����
:R3�q����m��t3{w��p:X�M<��1H�d��-˟佂�����͜�q��4=�iUb"�.�[%J�?e�a�U_���7W��o���[#i��w�B����8�Ұ-c�ʓ���lT�
D�]�М��U��V���fBm�a�1��P��+��1.t�]�
`�3��P8��|I���2KR?��/*@��a�ڗ.�'���9K$uX'�6W��h�ߟǿr��S�}~6��[�`�U�#uaKr�T��xX��4�0�Z0���7΢�i:U(�-�� r�[X��U0'iX��f��*��8|�?M��L01�0qʨ"����4��FP2iH%�#��<����x�d��T�R��֡��q�Ws	[9��S^�$�rz�p����� �$�g@�Lz:����`�@��"�$BN��W?{Yk>8�C+C��<}��bS�yo��E`(
��&��'��Е����`.�u������+┤�^hp���7���;��ݞ^X��HU�k��^���}*6��ςN����k�e6���v[F�j٭%���>ѯ�Oe\�7��c�(�i�Ds�~�z9�a[�Ѡ�i�u�����AQ�-�h����I�}��8����>��u���`�&"��fru<��.EE���U�ހ��vQ'�Y�������D��8�cp=%��\�
Q�0�u���
l��'�]]�i�H�T�4�.�>�}zdBɵ�Og�X]U5��m��
�8@�)�V�;E�Gˈ{�G��}�,�������0*�Ou�Y�K
 �;e�W�h�8��$i4�����.���)�a�e<���d�m��r�O�� �/ôT}+a}��w-�����63VZ��}M��܋��W)|�VHa�]����V��q�b�Ax�7<��`�Ko�"v9����>�/��8���-����!�$.��0�@��!�ڪ+x�}�7:! ���Y7�y��M�ni��0�b2�}�6�)�r߷��a ��#ȓ�:��
����ӻ<��DĢ@R������0�~��7�4 S�f�7�?Ԡ��6~](��e��������.r�ˡX|�4B��e���sqy@��Q��ێ=ٕ�i�.08aB�R�{r%���U$s���2��f?��{(	IDcz㠜�����[<���U�d��o�
f��~�zЬ5ϣG��=����(��s��̀7N���ڟD*\�u�3�K�2�K:j͛�FYD�
������"�e�D���[骽��>e��A�����5Z����'M��� �����xg����8������p6��^�i�g_>��S~���2CSW5lǹ�2cF�XTZ$����-�~���^���b[1�I9��]�k�bE����J����u�����z]`yx��!��0}圏���4�[4�p@����A����5g�^ɋxc'�
�&�����N��#�D�0���"�>�8�0G'�w(IT�6�G�Z/��)5��ػ�ߧ�< 2~��� ��hzb����9�?�9�@c��#5���w�������6Î$ң�輹Id��gP���IT�g�g�hN	;ֳ>%���P3UP�Hs$�P��1��O1�U5)��V��(����"�L��F���O��Y,���+��n��N�f77���<��� �KR|��WM�����//�����2@��t5C��CM�˝�U\R3�v����H����a:��,{=�
Xޝ�� ���yk�A�N��S�L����Pw���{˼x���.<09x�*�Td�?��&��q,Cn��-G~Q����&+�"�ڱ<�p�a)�U�b�Ϡ>��x� �?�9!x�o����#M�3{/�̤�~E{gWX9��8:[�����c~%��n��N�r���y���$�ժŤxy,!��s�P't��p8�t
�����0��L\��'+����а҂�?��5G t��$m/t�=���α9�&��Z�7_V�}Zʺ��vB���q��������̥��p�#�_V��z
���~>!˓��Z�Z�QӋ:�U+�(��oj+�+U���A�)�
	Kj�*��O0;l�<K
?��e̹
�g���M4��7&0�b�����W�����o��6����I�r��##��3z���r��'8""%S�rL�<N`R-����YA�v#�5p�b�(ـA�ac2�_c*N+t~AQx�7�Id�H�K�1wG�>р��,_��x�9�t*#�%H�Kd���p�-�SP��sܝ2�5�����|��Q�N�����$ʅ#�i]C�X��_jj���9ښ/��*�E��	c(K�u(;�L\�,~-�֚[e�!R���JUߐ��*=���*[�gd5�FH�����s�g�s��g�S���o�3O���y���L�V�e���2��haF¾K��&�<�*�^{���L5�����~�1��d��y2���|�����-y�u�j�Sy`N�F�;�Toݖ�8JAH5������Sj��c��p�š��oQF��v���R�-m%Tf�֌M�/G!r�u������9>q8�p�U$���.�3���1�e�+�XzV��N�يT�f��%�/ekE��㸿i��Ks�6e������3D?H- m���lVM�����Uc&®�Zx6�:j��Θ,�M�)�u�.?Վ'?��܌J����\�A˖�F$,�f|nBu=��K�]G���u��Ajr��Q�|k�Xpr���k����%c�+<
����qv^�6X���G�c�4f،K���Ç7B.)�c�����.a%=6:s{��-o6BD�б�(O���V/����iʄ�~���<��<��5,�ex�<OHc�����ˤQSw+������	6�I��{>�ݍ�r��Xx(/bC�'b��k�5�f[mb�4,K���)<�7!�oc�vVD���%�;5��0���}& ?�>�t_�%��<q7�Ҿ+�
y�@i�r��kro!��$��<O�V3ށ��do�IQ���v���QЯ�Vn��o����Ӫ(ՇF����K?����zj�� �N�ɒ`*����.���O	gM%�A�빓F�1R�}�~3r	�v6�����&|mcA��S��O�uFm���F^�����?:-�r+R��4����I�,)�CxT!=?ݾXs���	4,`f5~Sɗ��>m�J��r3�$lyҪʶ��ҭ����=����4�Np��.�vr��K�MY�Y�e�'>xP�~6L{��(N*K)'M
"���fZxIe+�3��Lc5�h�gQ�>���u�Xf˙S�Cu�r�$�G�&����4�hR� 9}U�V�gG����������_��g��|H����ӊ&WX�1�s� �_���Y����.�%m� "[Cx���Q?{BV����fƞ�{^��	d�$u��O4F�J���N�c��=n�L�'�]�Ĳ�([&f�,v�.�k�\�#�֠����.��"��|׮�μi5��,����z��U�yO�z7Ө�MmP*ް��z�� �E��5�PT��IO���%i���P	5i��;%��p�(Su���I��ROR�	������G±\F�xh�G�gh`�s��:8G �LH���%����۔=h�K�1���(W�φY{}�P��w΅�8�L5��!6EO�5c�AR���l�x�ϯ_�	+�����6a{�@�Q�����}�y~��]|̖��Wfe�7R�����E5�a����0��˓G��Z��#�npL��w���}~�m����N�i��x�]R�wf�gM�48Z$��no�;l��u��A�{�jz�>>�E	^�y��Hݍ��Ι�#AC0����t �Z�F��:l��G�3I�#J��³Ψ