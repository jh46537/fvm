��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^�.GJ��-��?f�b��(��ҥ��Y�����!���نϊp��=׈�kS(�?D� Y�S���#��f�����V8?�_���Mg�\��gѵ����s=�B_M�E�B%z1�����U����\�����ZI^C'���d�_ ��-[b�DU�Vյ��*�0��/�^�]ݚ�Z���r �Ї-�l�h� n��ࣁLR�5���e��G\"�JZ�z�!���0�.f ^w ϴ� I�L�J�ȷP>���ө�,5�%%�bK���>�͇_|'xƈ�&8�.�7�ԯ[����!�X��fŷsIE�~O�l�d�O!*�W,��H�����;}"���9��k�CD`Y���r|��# 媑6�x��31�_y����ъMd����<y �߱o��)a˘Q7���{;L��:�:�6�w�K<�&W�u��wK�M���b�[���h��������HC�δ�;ի'�(�����Ӥ�@��$ �V]z	u���#���ځ��2G�#�B	�}x��G��߳~��Yi�y+�����(r��ꕛߥOy?���B���W�uuB�d@�Z�ܩv��x= �ap��X��(O�vNleJӣZy�D�o��/�?t ��0��犢�?�T�*0��Z��}N�YE�1`>�	r�D*�>���NqxVJd� S�3459��]n��H�Dﻅ"��7w�a�t^|�p�v�5U->���^� �}�c��@T2��)6V豓�"S����Uf9�g�$j��j����{?��S�X_�H�_\��ݞ�D��.V�H��BF©�;)B�6ƨ��J�}���h�D��Z�o?�lq���U8Jݏ
sP�ҴŇ���.�~���1��?eE��uy�`e����P�S[mbe��� U�O���'��+�+wA���w{���W�Yٿ0aEU�&��0���Y�9-L��s턨gתp3���״a�A�*/�%��P�&b���5�p	`�o��� �i�ǌ�<�B*N�����`:X�d�~��C���ڲoG�3����`7�|U��_n�e%�PeV��-q$
�iZzƘ�y
�1�_�uT�_�8'��l8i�� h��p�����z�����>	��lj����Cm�.H����^ϫ�D�{J�q4e��4Q�%n1�*:rs!r��	����/�ešs��.]�����td�>�3���өX2��S�$��t.�ό���<i�+f|�s�y�' ��⫗���i��D�FBGKu����]�e�$��6, �C�2�Z�r�p'IE��Fa��4������2� KM�(��=sjfZ��W����w���W���Sc�W�ӏ$l�{2�6��~K8'�m'j����rR�#/����ۣ({�	,�v�P.��v���;0v[��ӧHe��i	˚�N�v���]�Âoz��T��E�3Mu"��W�&(�[�oOc����y��X����i����~�fRK=�%G!Q�v6�x���F�W�"��ٷ|�LF@�*IFƆ`}$~#c	�m���}����?�g�yP}x�*t�۟+,U�/m|(��c���$�ɶ۬#?&x��+2f�J��� .�֨��n�C`�U(/dY���.�=K��|V��i"s쐅�2$��N�E�ZQ�����<Lnbtw�O"6H��{oc�p�P�dܝ��Y� md���E�hDz� ˮ���ɼ���U�,[]���ęV?*7Dw%E6���0+��5k��{�}��r$��Vy���������3��3��-�)�."<�am�o�J�QTR��ϗ2�7��L��☩ښ����fTh�Ow�ݣy<Vz�ft���mT_u��!X�eq���$DY1m���$X+��e�J�����%ܳh����d�n��O��SPT����%�a�/�_��;��͞�~��8}R)�����"">��;��|Q����� @���P`����r>n�tC78��0X2R�2OSL!�9���Y�K��(�ﴋp��Ѹ�r��.
Eʙ��ҫ��k}~Qe[>���7�4x�f�u����95�]�Ш���V��)�ޣ>^B����Kn>g��&��O�o��@x�h�PĜ�J%{-�p>��]��$��l�=���ӯdz�t�Jx�7�?D��ĩ��6IEN�(:f"1/����-�Ѐ��'�X�B���2��ݴ��@?�f����\�#_���� L�͓�W��ʖa�M]��i*Ά#�G��8�{ň� D�}�,�r�iJ�q7A�=v��<��q��������o�W�TV�;�+2��@׀�ţ��*�Y|)�	Č�] %���I�Un��:�{�ŝ>�-�K	�K��rU���[�Le���<ܗ���k���2(���ج�~.�^�7�� �Qz\:JN��G�2�-z����� q�$�d�08�Q��G��ʀg����=�DS�a")::~��g�+^0$Y֫�b�c��*���&pagf�Q� �������Qka�t�#L����+(�TL�0$�#����O<[Gq:?���PN(X��Jn��X��QD���0;���2L�)����a:$�W��jD�6���2qq���t�	��
<7PY�*O��1�5���W��6*�����Ԛ�/+4��M]��X 'o���w��(�Ԅ����ݫ����8��Xv���W���[J�!��E/wїG�z@��{��gT0�qq��i��5��B6�-vh�y�F�>�[=�s��3w	�����µ�aU�J �~$Լm�po�P��B�Ù���6����΍L��x�����[ah�p l5O�z���r��@����/9dy+.�-T���<��x��	I�"MIQ��?�]Z��o�\�¿#�!SҜ����l;!��[��B[����ui�Uܴ��a�������8+��=ۋh��?-e�|X�((1�xO��85,�������+��*%Nj�����aKv�8� � �:�k��E�PPyUx�މ�;���Ȑ'S +'��Ұ5@j���kS迊ξ�3�9����n��L-����bF�KLw��=[qqש`��
2���A�F�xLs��Bez�k��I��������RS:��d�:�G�oǕF�n�|s*�X-d�h�Ie�7_H-L�-��CK\��F�*z"��ifA�ѫm0�]�4f��)�>�Y����̈́\|Ӂ��NN�u�TB@o;[X�B�t���{�]l��D�����Lĥ���x�/F�%��e��d��u�}�s�u��>�*��H�x�s�|�}�����#6=壌�wR?��H�v'[z%��]�zV�~Rҙ��g�@U>ݟ�& ���y�J�I�����ǝ��vXX1O9�s�ʸ!��%��I�s!$��'����v�S�@���5��ኲ��)�A@>tEk=�rQ%�����:N�e"�;�����<�K�6t�ˌxvj��	r 3ib���̆0C�~�'ί�4��Z���8�@H�ua�#K���o�}/�F�c���@/����[V����_O��aǺ�g�$4�<t?)H���㛾��y�.��>�/�m�������;�N�w	u�&Y��`�(�/R.�v_�}�>`�V���� ��>����V�����?���ZZԺ�lXe�a%ZC�S2���0d���k�7�KW5���{��` �G��t��ӧk�na�S��UEc"��b4=������p���l�,�}���j��|$�'.�b�Sk�Ae�r�$ynrL:�����Qy�^� �K2�� �.�x+�g�SeQ���D<v�1��lHZL�p��?2'y�K�	8�w[yi���dm:���!�%d�M�>=x0S����c�%X��&h*3`��atrO�������$�'���ʽ]�=�S����~���� o�0q�	$�(T�L���:��u�!Y��t���2"�g+/#Ƹ� �@l��'HdDW�N���.D�,��G]���h�m��9w�a�������$f^lh�|����8�y���2\IUwy��O��!�~⬱Y�5�@��G8?�/]�.�ΑaU�����]��s�w_�v��tz�d�t����|�[��?�� �&Ժ:I���sU ����ҷ@����������a@���i	�TE�v����~c�ě1{�f�r �7$��%c��LH�\4Vt�X�O��z�k�#��(����페c���7|����=�FM*e}Juw�)<���[��2�Ď���5��>������Y<�Xr���W���WKˆ� a=�<�e�`<AJ�.�?r������^�+ܷ3^B9��!c�!���Y���;y�9�U�c����]4�`|B������(ӽB�:�NO�>ݠ����/��z;cq�:P��i���1�`tU���.��G�8O���͜����Sн������SR�zo�?9�V��Ϝ�{�^~�*^ίjw�$����~}��Di��s��x�΃%���@j�K��/	p �Zc����9��/�_��b�p*���d��W(ͫ^a¿��́�R��Iے���GaF�␸�JT��kɢ)��g�u�{(ҸG�ؖ:R��I�ٍ�i�U��͓�* A ��?�i�逡�t����_���՝�{��uS���S|Y3��3@�H�/jc[vнN���k�ۉ�_����J�;�ʶ{�o�!Q�$��x|�i�5N3�I�;�vh�U���9�?;?''�%2��vy<(�G�.Q_G�;��N5WA��ݵ(a�Bj��s��,ݒ��Wۗµ�C5�9��-v�l} 
H][�������0Ï�#�4���������⸷���t�( ���/�j�f�>da��t�{?��.�+L��	L��%�n�[&�b�18�6�\,}'�� xKr�Y�>���i�^�l`ŀ�R�˄?�Qab�?HA��Pz'&�ü����"�_��(V�:�$���M��i��hN���<�Q��3���y����ѳsi"��e
F����v$����I�q�b���Aw�*�#��>��Aװ���O@N~~���6)�A�1��n
��c�4�m�.#�{�(�Kf|/|�ը��=vEs�(�4��*�s�W�D7Z����v����@�Юݝ�]�<l<�#��W޵"Vo��ܹ8�J
�N�L#BY�$�{�!)8�+(0Q؅����=�D���)l��"S�W��D�=4*5+5�����RTۻ,�'���x�V�K�N��q��$dOF�̈S�CΆ^��K���C�_ʎ�{�_�KO��r���H��tv>5��n>�n�Ԝl-�� ��jC�:w~
y�D���h �w�Ȳ��^��+"Џ����qJ��p��;�IpA=�~�<�F��9���A ��H��H��
D&�'�Jd�	
�k��ґ��ڠD�1���ȥ8�[���4e�+�����d��yh�
�����9t瀉�ऄQ�p���~�[�i�L�@�I� �y�3/�a`V!���S Oa��3}��t�����2C�����K���!�5+n߰�Cb�~���Gv��t��N�`!�s&��s�F �HQ�ЮN�rfݳ����Y;�,�PD"�ӓ��Q�wW�����;��-��
I�'D�����ׅ��X(��}2�����H�иX��C��?�Wpt_��'�J�Ĕ@�C�N?O�����&��P� ���&�.ƣ�@�y����`k������Bɮ�M!=�<� ��w��ܳu��>C"2��B�Iy�1�>>�Ĩ�Y��[$J������ؼ!�:
}A��?��*ت�����pR��م	�Ɣ�d��E��_�&���7�SVzVY��'Ƃ�I���R~��/�u������u�c�\���4g��>�9�8����<=NDᄋ̎�fW��^��x�sS������-��Ŋ��zg� -�fI"ϗ�S&QW�o�)��+H�l^)E����j	
�@�ۖ��4~g���!��S����va�����{�;�|���.�f��(�����^p�gY����������`��17GCO~�N�L��������G'������y�Bg}~�M�=��]�������ȏ��[�+�eKW��X!7V���{/B&��#9�>�`����YsZ!S���!���\��.�z��+p�h�:�^g����^)�[|3X�9|����U�������$X�\�T�/�XI(I��@�˟_m���S�����h����h���� �j};��:ʩ�G�Y�+m��P��ҚDO�"��:���k�uI��U��\Bs�F����j8���������Њ�D�ؒ1��� �D<����Шs׆LWzk�9�1���ş�Ql��:m����k����D��Ϳ�)���2�&�u'��o�<}M#Jv&Ǵג`�W�� �&5�Km�����v���͌ ��oY�g.b �x_!�L����-��uǿa&���3F�v��:fZ�A4�,�޼ҥ�l����G��	��0wג(�g�`�[����x$�����#�Pމ�pW�m��IKT��=��H����|3�����{jh�:���8��K��Q�j��3ټ�F��h`J���ixY�܀J���:���oD�KǶ�����7��Hw�ř���V2mnS��#x*���+Z�(u��_ _1+�R=٪-����{�@bj�m&H&L���)����6G�Ɔp�D1�j۶��33�w��[�d�k��LI ~��L�߼��I��,İ╍�<�W�	��U�����R���� �C0R:����N(�.[���E�������ЋWe �X� &:!s���B0)��Ǿ�ց�p�Wr94�����@5V'�ؗ WF�d������b�W��#���7'D��U�
q�I��݁�!*Ѵ�3�%C=��u�!�-j��l�wie��Swٺ��*�Sc�(������o���r|��Fpk^�F<���.�,M^H���L���/Z�C�q��S�ן4���Ma����b*�"�f���5H=�-�3N�{����2�����v�B�@���>���\tr�D����)Ζ��g���{�[nƈ5�i�e,?�պz���W���U�y�{x�����v-�,�&�0F��uq�N��u�j>OL:%`/�Ø���!���>)@�mH��䤄r�`h�%��Q�pG|�P�=MM�:��?�v��"8�!��U����&�gS]\�]���Ox�`p@�G��t6h�nm�m�k���F�`V�@X�;zE���I�y�y��La1D~ؽw\�!H#8\T�"����jv��an����g:0�o�����١�*n�V�����%-}W<.�Q�Fx���|�+Kh[�
N������ �D﫽n�X�ߑlW�ƻ�e��-ͱ��}��	��1����~��(e|>��El}��٥�A꫟3��'�#Ww�>O?ș6~�R���r%�X�	p�6�'qCv蹿�!N���٣��Lo//#�����ZGo�F�8���QG�j�J���2ʢ鑞2%�~\�G����fy%>>_��Q���(V���Yљ-�T����#�׫�C����r]����S%�,Ϧט:���YV����J���-H�F��
=�p��[�F]��N�#�?�]ų�>v*B`i�O���3JN��R�a?�sp�k�レo�gd� o��Z��i�R8y�^�"���.�S.����V���(|�:�e��%��ɶM����~���c�1#[�x��V5*�`��p�S㍂ �'&��#��Ӡa�?���v��`��y�v����7�~s�-�����e=+N�ŨM�qCE�l������"q(`��mRZ�oI_^�4:�`���$HZ* ��� O�es8��I��R�7�����JA����l'&��gS����%��e�řQ$jP[�ˠ�ҸC��a�ho������d7) ���������u��Ә���\B�n�B�A	4އ^24�oBg���%��Q�-m��6���Q�lٻC�4 ���+%��>����n?��;R�Wq~�su�<@�6@�z/�0da��E��'5��y*Kw9���{�r��GЅ<{>��iBZ��Z����g\k�Uf*FE�n���V�������a��Zv���<�m]�L���?��Ԍ�^�LFҋ���0���A�+��ɷ8� EȜК��-j3H���-:�X/�~,,����vof���Ax����@���VC8ٳJK�
!7�=���-/�0�I�x�j{�ų �W�I�yR�w0�l�����f���5A?�x������"�z�%A#|����L����U�:��0�}��?L��'7��t8�2�H)!�F��}��������<��3=�EdOң~m_q]f�R�_���o�yN�ig�I���|%��=�*������xK��`H��~&ْ%��U���W�bkn��!ݗ_c�5-,�!Y)��R�1T[^#�<�C����:p�S��el��n�vE����ݖ�!+ùt�D.!�8�ZA/��D-��?���@��
��2��h�&���2�w��м����M2���k�lN��ɯ�s�k�� [�W���g�:9���'�b[�o���;�2�%�nsς�f� 6�Xj4����k)3�jyD5�9,�0g]Lc!�sb;8����Q ����+0���dpH�?��p�D����R�:0t����e���V�yZ$q��L0.RI�^�]9Ȉ;�E��@��3����z��>����;�R��CCӎ�ۥ��7f�����W�߉��6F�Gb�	.���[�yyuklQ�`A�9fM�o���Ʋ�K|�iVUd�:��IP�۷���z9����q9� ��]^���ʖ�����1�˵}|��Q����0Oة��wzO�1�>� �O0�z0#ѢhIN�E6�'��1�5�p�3'Y�m=Q ��e��>�Y[.&�`�ja�	�\*���s����g�o{B%l���=����=:s[-�SB7X�kZf ��zq�=m��QD݊�Pǘhw�N�.b���R�� *��}E���v�}�x�NE��|I������ȶ1�N��ԧ[.[J��I����]�<���ܝm0􌵵�LKSy�����;����5���I���z� �3���?ņ�0��6���_�قVR�Ռi��@�X��+�
��I�/g�sa�r���8ˢ�(!B��Z�9�>�g=�%�Ё�lBd'U$��70,)�����6N�MZig��f�6���6�ggE9��mw&0T����q6)�<��wu�B�>���N4�~Gq�-��[H��1Ĉ^�8�.B�~7�\�7�mì�p�>m�eI���cq�+�<�.�?g��Ҭ�3-֘��i�S�G?5�QQ4.HcD�#����X*c�5��Ð���:����77����)ܗ~�Q^U�O���_�:�L���%��K#�z��r�ƿ2�f]��S���$�(�e�LC�q��R4��8z`�.�|����`�@	��v��c�*s�W��=����6	�2^����_�
�ķ�O�w,M��0HV�1Y�l�>���_ c�[o���A���[B*�E�����hp�^�
wT�G?���A����^�������먮_h{�.n>-ć��X;]�$�}=Z�e���F�P��z�OID�j���؃���\Z=-�R����Yo�	2�����g����'b��WwQ�ﯲMD���a��dM�&�[���?G�oJ���-��7�$�hJݸDS�a]L�Z��Yz���� �d��X\sYC:���p�.�9z��EB/�� #�7H���-�R���;�s��\�dK�?}��^��?v�6�}�¿�Q�p�]� GI�]�^y�#v��V ��,.�C��`}�ε7LD��ŉ9�ۮ���җ��ǭ�w6f3�&�$�C�3�|����?5)(z�|Nǃ�E[�Fo�/V�L},��=B���o�Hcl/�J���Ȳ.>e��dN��P]���}���"NHO״[Ƨ/��R��f�o�~���=.��.�I 4\^��	��إ�쭀2�zdɶ����H�Z�7��o�n�� �O��/'�a��:Y'bⲿu[��O����1�f���d���9���%�i���gS�-��S
��-�_�6˿�a�[�����"�*\ƀ��� 5H�7>.������\@0M���M�xW[ڎ��{�y�f�i���$�GhR[ȵ>{$n�g��J=�����^ �����)�֫��a�h`M�����'�,P�^1��a~�y�N�Z�����}���}�5�Ѡ񠸺�i�Ę��}(߹�_��@|��\�&n�DH(�W