��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb&�L�S��O�e�m��R��`�=}M_B4O<�o���6+1QѰ�tT敬�k���K���b<��͏��A4L��Dm	�c��\�:�>���ئc���U%g(�f��2��♃��3<;����@ÕG�C��NCo��&5A����b-��:���Pq��;�q�����6�h	6/�;
���6O}��u�g5��:cA"�}ED�$��>,rPY@��ɮ@�~kF��W��d~��Ki���6�� �-��H{n@�s����ꔻ�^�CRM=9%[�6<N&v�6桚45�
�*����dE�����{������U�̩Z*����kG��щV�W�>�D���)�B����/MYLCE�;���Q~)T�[ws%_S8f��`�#j�cf9g�O�qt/��O�Z�>��2I
�CJ�U�% �t�[�ܻ�����⼦��E�µ덒�[�q���v]�kFT��;�|�9V����d�z��Yw&��p_	S7&�tT��
,>��S��诩<����A���ty��w����;֖�բ��(�[�N����2ff�:�_2.Y�M��1�%EM���=e�n���A��r+XjO0�������۾�c�{k������ԋfkY�ӯ�Mt�ݘ.�dUP]��p����)�抆r��_��x�'��~eh�YȄjS�ո.���+cT�%W+q�j��p`{8���D�����Y��!��L�/�1�ɠ�uW!E�$n�b��ҋ�����qc=��/;M�t��	Խ���)VH��xgY��}��l����sO,n�e$�3Ba��[mo*Z��⪻�@��X���R*)�5�t���X�G.�	����
ԣfC�"iL)a�+T��H⯧�3�>j��o�.1�(}����W���	����;��O�̠2W�*�n�v"}a>a5�F�j�nyaS= ���B�i���t�U��E6�8'�ҶYa1z�d��;9����d�O�U�����X�)�Y`�|��b��C�S�B���y�*?Xp8�;(_`�އu���׌o�ؽ;�oFV���L3�<��N9$��e����i�5�Ȓmc#bv��V��2���hX}�V�+!Jݔ�}�o}Wo*x,阩��J���>=��V�.|h�!{R\������Ɂ,)��������M�P��ñO�=�{|K��L���{���
���?�O��rn��o�;��)�pM�'��G�|�1`0n�|��n
zY��y��2�ӵn)_L�)���7�fs[P���_�����7ǒ\J��`�3�4K�a�z^:D� ^�ңbZ�H����AQ5�U���K���g��,�Iʜ��C�9P��L�L�%��:M�l��o,p����k��L��PN��uvW+�i�5�t'�Z)*)�E��d��kZKԻ��Gx�t���?n���L�G7I�m�z�_��۷��D����\��m��o�)��կ�����.O�𭒈g�1���t_@�mӌ�{mڼx�f|�|�v��ˤz>�`�%���s�<��*k�b[��;���`�[���A=��G7�{H����+u����wY;P�IJ9tC�L�{1���<f�՚�A+��5�.��?�:��1�3���O"��	v����w]���h�~���a��gA?�q:ٻ/�M���@�'=d��tłgzh9�=.��τA]N$�f+�&�t�h�V{ �#��/��"��v��fJ�}B>�Dr�P	�`!������������#�u�9�*��ʑk���:���FD�]�B�lX��lw��8�ltT���*?虮����L�T�:IAQo��{3A�Z𸭔}����C�	��u9k�&��D�����dA�b`�U b��[X�[�u����y{r4c�7y��9��i;�ҷ���s���ӿV���j�ڗ�@!y	�������y�=�JbEv�^�z�؊�_`�3��2�څ��˷��:�]˓x��٭�01G�j���I�p5��@ܕV���X��Ǩ-��\$�Q���N��}ʟ$ r�ܞVń>D^ó��*-�|�:4]�Ն�#s��uЏ���>�����g�|�c�t �Hƥ�0[Y�b3�G��$·@����Ua#�e�W�uL5P/���WTR9��� �Tw��w��VML��V��d�z���m{�g 
���~�v��rJ�E�H"�t:�&
��Ϩd��dQO;gq�e+_O��ap^��Tk��b6�vWN@Jq	��-z���>�q�c��D9�B� Ӏ{���&�����vs�(Hz!\�4F�D�o��}K\�l[CyݷS���Թ���>�*F�tIu�	�R�z���*���P�50�hd-�%HVEғ�pq�������Q%Gi�qɭ';��T�\�驠�~�����d�Qi���B�������r�Z~ ���z*�G�S����:%���F��[p+�+����bʁ�"h�B��
�I\Ӫ9M�0f�@f
� L�䂛���l&G
���T��^H�b�&V����r	mm}�l[�R߄K��"��#��AC�R����	/+�����|Y�[�T�n�X��魞�\Y�����}��>��HͶ����������XT8�!4�7y��6�k(�f�
rF?U����٧�����)b��R��N�g��i� �#��:����mm,�}��r %�1c�lF�m=��q��$�n��a�R����]�R��V�l��R��l����c��a��F16�D�ڽ�e��ҏrX[sJ��~��kg��lL����|��D� �oI���<�5`N˷*F�lw���iڕ^GRot��&��_��1����I*5� ��j����)�]W���oA�tCE�0�@H\K���}����� Etk��P����-uO����������:�ʦ�9��q����]9�2�h�^p^W�Tu������Z@\"ʱ���$��vSj��{f��N�t��mEĄs�!~��}�����\�У1�uCXr�R���~Mw�r��n�I�g��TZ�#k��,T�uy����$˕�X��i�Ggxy$]��K���/��$T�������hP���L��c5�~�43�eq���}]��>�
�I�¦�;�E�����H_/C�#�i2�m�u�����Ͳ+ccY. O��҃��	�6D�δ���X=3m>��yc������ڑI1��p�^RyN����;��c��ܲ�����j�D��������Mq&Ct��w9�EC��#����Ğ�PGZ�z��A㝍�$��`%� �*�
�9�ΤMbF�453t7�P's�����y�%��*��2�J��^�F�����Ie<m���i4�QJ�!-�����d��ԬRhY�S�.�� �]��ҟn��<Qe��B�� 5�i�����H�*!,�#Ǉ�)Ю�X���U[�V��*�L�i�Q����%f3���ǝ��/]m�G�K��=Q7�W|G� V�w�*G�E�8O4��Ƹ6�����\P�9[A+�$�]��;f�>7�����6Q�����k�nE���8�����P�6���o�[��E�\٫(W�y��ˈf"����p�s,��C�i������B�]���@���J����M�>d�H�u<^��c���>Nk���FV}E:9���1�SM��`Lj���ʨ�X���QZ��	ɼ���c�<��~�c?�6E$C���ȡ@�y�G����-�������vV�ܡ�R5��ȝ�`���X����VFVL/*َ�0�18�Vʛג+rɶ���v���?�u�U��Hit-Cd��w�h��b+�`!��R�A��Y?��C/v1Ӵ�t"�0�}�a�>�m���궴4t�d~� R7�uj�@�Ѯx�#F}�]>Sڛ����`�$k��ր�\��1k&�'>���w�m`��?ָ�#�j�U�;}����R�_�/Y `طA���6S��8�k����D��_�m����i���%w��h�97KmX�_jq��O��^ʅ6�
<�9Sm��Ee3��K,�4����nTwd����~�&!�"W������ QĄ�v�+2�҃����:ç���HC�ʄ�����\P��y��E����)�8��Ю�����N��4�5��v�J���ꬊ�@)����b>�^p~��sl]�n%�ؙ,ܚ��8�*~��YV�0\'?VJ�X�k�μ�R7�=0�dmG�1A�\C��C1l��D��>`����`��ӈ+�Z$x�ܱ�de*�<�������8�Ñ��R�0�s<*6�ܰR�oV���f7�-[
�h<Cb�!����Df<�d3�q� s��������:���"
�B�r�~�C�� @mc`�,�T<�O4'�#C�ݯ�1'� d��#f|[�z��!-F�
07�gwh�s��)	���)���A��Vl\���c~.��2��������{_ӅJ�j9 5ˍ���Ɣ��T~*S\�e�zZ̈́3[����1&��t�u�C��NS��%4z���`k���Ao���uH�y;���:�X�� �/D��<� �jYسi:20�a�Ic=�5'"��;4oΩ��!զ\^�6 �h���Nm4+5�����}yx0��-�U�zI�Ȍ�L��P�ٖ�F�hI���K2e�������%�um��j;,�����+��*�d����NY�yo��o��G\J��OO>��{|_D�[L�b�	Y�n[w��'أ���kn��o�8zgeE��ƁF��ŵ����i�L��e�)� �Wk"
��y@?!�G'o�����\4i���K��)Պ`�k�0m�:?i�F�� ��E8�I.�ĽN�[�����Y�u� h�f���ê�Z�D��^���?��X)�?� Ȳ���5Եh���bI�\��Al 6��L^�i�/�����c��&��h��Γ1�k�W<��p��IXvD����
��G�ȰrhN� ���x��=��UV�!�1��ճ��ð',�&�SfB4�2-˫>;nҔq!���'As7b�Tk!7	���Ht�33F�AX�����7}��%(b��{�l�6�.5	�d�����+�T�,��Guy�;SW}
al�#��{Q|�Y�J��߬Ic���j��W��[--S[{j��B|��Zr����=fW��lA���f��\o,��H��#E�
�;�So^��8Ҿn;��{����
�H�	>B�y���@��Ϛ)��۷v�[#J�zrG�l�b����N+��/nUߘ�}>ޫj|x��Jg̫��aOI�ɍ���Z�﫮�f�p�'8�8��.��p�E�Dw9o#wߝy,��|#�.>�O��p銠ռ�2_���V��l�52�Jyմҏ�7�+kg[�l�K6~=]�{Ң����"߰��V�(ԯ�� �V����~A��Y�-\ӛ\��/�:=@ra;��"=��C��b=*�z��������,+H�w���G�GmP�� �����B6���Vv�ۀ���<vz�c�}j��Ɔ��暁1�C�WH~�c��H��ַ)�S��fs�Mz�/F�f[
9�3U��\������8	ě�A�6��8=[�(�œs�������!�j�P��T��ȋ@�{2% /�B��)Q��� �x�V�5Z��}S���dqCy^�'%	�Z� ����",��|UT�3@VI��[�@�u�8�e�{�P[�����n�烌�	�@q�'tk/lL_���i����M޻-c��}��Z��6o3�n>���7��V��e������ĩ
�����`��@ �D�Nf9��|aO+[h����h�s���"���ј��bmb���e���W�����O_��P���>��l�͑��!Ǉ�On��zJ��fVB>Qnڧ��$�w"Z�(�$�(js7猥�l��_3�q�_6+֚�-�^����r�f�f����w,�S�������Q����گ���[�B�*���AT<%��1a��t��9Z�Ig�~�5!����N{��5�?�Z�=�px�I��9ծW�?'ǁ�A�=�������wT&�<���R�f������L��v�d樤w��U��A)��u��':���4ߥ��}n���{�S��Xw���ZZ�w*�\.W���`�M�]bL	c��˱��γH)�9W��T*`̗o$�U&v��j{��@��2�5�hS��\�'�q�*=Xc�I������c�F�cTޢ9`��L���sD��JQ]6j����x��#ӄ��[����RA�;����5�J�f���mX?R�l@)Z�뉂���K�s��H����!�"�=k�-{�7�3M��Y�g�j0�� �9u�����炱�=ʊ�E7lo���t�}�BS�)����eI�~"�h����p�{�)�4����}��?_�� ք��WV�#����$��1X��	K�q!yD9������9��ǳ�|7��=�.�֍���j���Q{щ�g�3���iW|CRH�c3�jE�es����e|E%!(=�r�ު|M"���(���E�);.ƞ.\A�*p��7����Y!�v�)s��Ċ#�(`����5��* ��C�iқ)���R�Y�>գ��	>
3Y��t��3��-�1��WA~�t׭H%4�t_���Px�s�Į�#�0`2˪�pd`�k�є�3g�V�h���qW�y������&M�XE�Z��n}�?��د�8��E?�ﰎ~#������	bZ,�[�/Bw��ا����x���4s臄�j���L��w� � 
sna�H<U��Uk�W U���v��vk����|�@�P����qK��a)�����DHW9I��RJ:JZ���:v%���\���p�)k��|ߣ����0��7vF7��\@��^�߻aOáB��^C�U8�it�|&������u���'0��/���A*��.?k��'��H�6��KpS'�9�Z��9�=4��pA�XB��P
?v�J�K�O{�heU	�[�� ��]f�>=P�e�l[����^P��y=t����I�߹ݿ��9)=Ҟ�c+Q�=I�\���ڌ�\y&�}�]�\��S~V� 4�8ю��S�=�^ct����K6���J.f����(�� rӚ��2�����^ߍ�-9��41@r��#/���
Kk��Y��e�M?��ť�C-��]~��WgظӖ�u �i%X*D �>�8���h�2��q �<'K���"0�����F!���\�e2� �H5�ȼNV�[�J��H� �������R�r�P�~�f��7_�`�Q`e�ίmW�e{c����������(�9��~̻f5As�^&h�	è�wG�5"�o@��Od�Tʟ
7�,4�n��9���ol3�&v[_f�`�&[���������ss�$�V�<�#���Na�})��?�D���C?I94�q�����^Ӿi��k�D/���«�^���`�����W`V�}�S��������߳����S�^_Y�K]���添�R޷4j I������S>����8�0������^D\!û.���k[H���sӄ� ����e���0��XB�Ajn>_SNH׺�N#�����8i+�$�mq�}S>ͨ�B�U���i���5����ZGߘO�ˏ"�s��ݑ}Mc�-!����������%B5�Z��T��l �t0X�tG
T�}F���}�] �`Y�?J*�ˮ��{��}�X��@v��^��$C�DP;	g+�Z`��a�\-��z�$9~���.7����6&l�����w�@�Y�|~̈/��b	�4U��2�:�[�&���4Nrs����K��sIT/�c�(c�%ն/�uP�A矧�\�2lGo6� �x��FE
j4�°����W�.�Y�^��58��cʆ❆��L,�S��[���a�����e�TvN ��"���pJ
�Y���q�;���C���!��x��:�(��������؏0��wvc&L�o!�����0_�4E�Ky�W���q�a��O�CG?J@�l����.�Ԩ�
ڸ-
"���%���T���By�7u�J<�x�Ȩ'���^��(������ʝ�8�-<oXs�z7{F��%�j#���o��>�~�XB��;�lӾ,-QT�G����k|�E$�>�b���X\�iK�?IOF;�Ѭ��7)� �f9Hw��\������ �j)��~���N1���i�٘���1��D��hl�H������CB/�t�R��"q�&�H���	�H3T��Ż`U�@��>����5S��9S!z>���Qo|QD�-_
�J<i�U�o�;%S���8�g�"I�����-�Xj=��[#��_d+�v~GQ�	B�("�}����(d�aG>?w*�\�a�縭�񈈴5K���z�]��/�(��.Q���`S�+;�K����H�ýFz�?���� x��ת�H�qsy�Z�<`V/��p�I@!v0�� �ϦR����7Z^�X�2�2w%�_��\��t~p�T����D�ˑ�h�l���r�pl�4��a��ޖ�_q{Qx�
<o�.��*ۅף�7�v�+�e��_hF=*��&q�a��v= ���q�-F ]�n��ؕ.͙�D�9v���h`�4���#�V�:i�}�]�]X<A�P439����@"lƇzKM�OY���s2sQ��2a}x{��d.����'�����J�g���o����"!{G���5�0�����~���
�~���y2�c�1$W��F�Ve�m��*��ä��AG�`�Ϲ5o�m�z�eF�5�[5�D��f/��l/�6�(��5}�*���E��uכ!�Q�f��2Cs >%�L@����^�t��a7'|ؾo�Sˬ��
 #{���GB��4��n��������7g\�bM.4h/��E�n�S�����$u��5�r�`�T�_���{��i��Z�"^��b�y�߶o���$�	�c��v\ߐ�K��ȁu��c&=*�[ �l@���/|���+���xպ{6U��G�!�YZ�I���p.�AsR��t�ű�ј �"�(O���J��W���E���[Q�.�|�� ֕���а�>+u�y�xO
�s�z�Jx�^�}���o���_�e�($h2��t#z��0��;Y�kT����|D�VH$��ͽw��jW���I��Pɋ+l�>&�UԜJ45����@�!��a��;��w:�᮸w�6R�DЍ�
sT��1�7{�+�������J��w���홡dy�����8����������C���Y�6x��n�������ÈE]I�w�G�ǻG]�K%��A��,:h˄����_>K�к��Y����_���_�-�V���A�̪�kEXm��n�Y�U���^�g6���F*�p�ɡ��=�_��?�k�Xh�QVx��Ŝ��Y�J$֞g?�݆Fn��y�L���9�=���.M��7��!Ԕ��M��V-2���*�Îr��i����|~8r�Ҋ:{E?'���{���B]9
���<�A4��wq*/������0T��D�L�KN����a����'�~���_ܝ��w޺5����-OZ.���Ȁ)�DZ?�Nt� �B��"���	q������U�(�:z�BǌK��/͖�̐qav��4QB[e��L/�q�%@�����|�i�v���6V�G �n��H�^�#G��M߽��ݮ�!M��=�#ǈsw:Ҡ�1�}ƺiZڢ�f�B�_/�@*�JO(��Mu:U�<	R�������V
�������w*�X\�����h�	h�n�:V
u��#u����}�4g4<��｣��B�֖h��DD�PV�Z-��|Z�R���h[��>��4���P^�۲ḡ�����iN���?�E��7�U��?�@}Y Ng��_�mo�W��C��tY�0&�7p�_o&V\,ϒ���Y�c��)��zh@ZS2۟�9�>$)Nc��oS��"BW4�b�`ڢT����I7F]7���~�X��P45���p-3��!��b����U�A��=j�,�{^SrrU�����9[�[=�Tj\�ɲo�Z'R\���ɖ�����