��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]ǂ��O��˰�	JL��Guy6A;��%��:Ԩg�P-fǤwA?����u�n=|cc�j�/���\6[_�����lVw�ĺ>��Vuth�:U+5�N���e��Y_P��M����*�C�Ci�"bNq���ů���Q��6I^�>���S�K?���_1��pzY�'�5�^o���X�����X���֨�����v�Np-��ԅ?�qr��YM��6q����"{n�w�[���%|�όWi�N.��EUf����U %�k��
m�P��� �Q��PO	_�e���ś�
�bh%"������H7�3���7��j��A7לB>���D��$'w)��qP�D���iZ�6i�(G���Y�L���n���|[������02���n�M���>MDԒ�{���tDJbߵT^4N]ۭ����f��i[@c����p���*,��r�F@�G�(