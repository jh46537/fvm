��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħP	�(<�%5,i v1`��;[���({�.�6��^�����*���jIJ�c�W ,_��������܅1H�d�ӱ��v7s9���3�qvi7�yk������g�>�p)�'E|ȟr�h.��(Wp�_��T�
�vL�ݞ�6[��Ș@�[.S�V"CЀ�qK�I �e�$Om%�'�![�&�2�7��`���,�3y=in�����;�5W�(¬�б��������uiJ�����-�L�WNW2�i�!�%��w���HX��&��1���v@!�Y�sdke�3�w.7)�h�.u`��o��N���D���'�"ܺ��C�������� x�9��=� ,\&+��BZm��-8a�����F�~&�c�9.]r�UKxe���	��<��V��è�^t�0�O�l �KF��J	�p玄�c�kmA���K�jN�#���q��g��̓%��?��I	nH{;���	T=g=��������(�Wެ�:��IZ�!�7ˬ�D(LLΫ*qEN�e�R�Gۖh}���_UQ7%;꺹�X2��˳g�6y�X�|�g���*��L�������}3|���\�XЍ�>�G������r�8�]*d~�!)�یf��x�m(��:E�L�bŕ���>�0�L��&�Rqz@��������C��~�UHM�[�Z '8��$�g��1{�3Z�ٙ 
ŧ�#�%dG�D�t�=k���-`����o���:ߝ�1�ߟ�c����O&Ɏv�v`�TA\{驩����� ��H1��¥}���򩱃ڣ4ZM��.���>è��� H(m5��ur,QG4_/`/o#:'��`7l�����J�'lPrC�_�y�#�N����B)!>*��3=��I{p�o�h>��#{�K����v8�- #ӗ��
�2��?���B�[����}F]�y�����,� �L-���!yB�a�ֱ�8N�/���G"L}j?��v��sF�V���55�wt	�Y�v09�t��H��f���0�%�T	e�w�Q�T��9�x��;HwXP���S����?��?��´�!D�7���gC���h�)õ��o]�`7^�Y�}^UEe��K �#�����m�����eU(�>��n�)�5�e���{�Xx �����.^�T�����pR=��7oʟ�� {�����}w@'�&_*a���ꋸ=��;��G�����d���O`���!�%^��]W�b-1��Kɽ���������K����.�����k�\�4��<���iw�N��_��Y���|�u�N{L)���>��Wll��m�Dzm����p(��YƼI���|=ܒ'*<�"E�;N4]�aZ[���,�0�6)�c�,f���Cy6<-+�N^8]a"&�u}���Z�x19�<�� ���Dt#�|�]H���az�\1��t�
��k�
(�Cہ犞��;YtQ���!Q�pݘ
��F���
v�t���*�1*:��k�ݡ�y�pE->��pX
�����IkG�Ā-؏�i�c§�Cc�o�ity_+,��o:�K�$T{��v�⎧dW�$�.�5�����,�%
Hq�������x垴�,�o፛��pxR8�|Ԇ[�\���J6ߙ����n�����!�W]�a�J