��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��!N;�?'ǝ�{9�1�\��,�L�B�8��V�R?��[6F+�+�4"p���n�d�#�$؍p�����.�{¯q��ěW�F^��A�S*��|��Ea)��sz�$��O�+�d(�W�n{�|��C�:� O��U荈PjZ�h�'#��}�Z7��-?D����͈#�26���1�o%3}V�9M5@�����s���F��	+�5�������S�/	��;;�~��g��JRyyҩ�M�'������Q����4�1_A�<�����E�s������?�I8��6U�3[����[we'C	�De��m�!L�����;ܜ0��V�~Ջ�r|��˛a�1X�=��
�M<3��(&�<�<���U�p�b��)��+1��+�����=�	�"Eβ�,�������pR�Ry�+f߮2j�۞o

�,>��������wX��2�:D�J ��� ��<���h�S[��h��-(��(�s0�9��5�[t��s�Lm�����S����f�fQ
���3��?�$7I��Vٚq*�T���8�!yxɕ"��f���&���4Y�v����^�re��F��������]���g��D���?��EH���2SM�>ZT�Ӷ����k��ֻ,��9p��3��XoS���,������vtD�S�Z0#���:0��8��Bk��{����7��e�ecQ�6~�|��/��8������y�dgO��4Y���S�`�_�� �8|C����6 �N�.���]�S=W�h��5_ @�WC8��#����d���.'4����'5C�'�Qw�V�m!DP۸2O��Gv��fr˖~l�2���^+��,H9j���@��W�r���,����+���,|��֘����ǢH;�H�xV��q5�nR�<��îɊ���
��r��P��5V�%�R��4{N5�1w�A�*�lO>��㉲��
� �|�w����k�w�'u��G�|�p�e��x��~�'=2Ҫ�y��<��2�!J?�q�؟ +��_K�2A�}���UM��w�-�w���R����R��g����p�aV?.�V�Y���Z�"�h�������3R{?��D}Jik� ��$��ĳ<!���>5�\�?b�䐴��,���pB�L��W/�q� �\d{��#�s��c(�����+7���.��9��d�w���d�6�;�H��{A��hɟ0���||x0��L���O��8?q�B����m��`K0�L��nI\.�Q?�j.f>��������?�.�m��z�2�+ޅp� 0n�!�0dɣ+�P��@.����`5c�C�AMI�h��r�*�ܨ��J�Z�Fnb�$Vc���i6�̢y�tf]׃��,�����wsk3�����Ql�#BϺ}2Vӹ$���f�X���h�����sh|kY!�x�%� ���~1�P�h���!�kQTY�c2�%��{�`ݭG&�5������ߏ)X+ׇ��ٱ*'Aca�땉ͬ���Դ���1E]�F��]>Ҭͯ�tBl�Y(����%��ƏR@��<�#byJ�%-�3s[�?��JQ��h�6Ӡ&:��^?sB�H��o�4<�ڼp��qݴ��E��@��^����$[�ko?�!B�R���3!����.���Ǒ �mDb8��)yMZ�?�Z��=ne�����w;�f��������s���\��'tɺ�P{����"�ZB�t��7(r��b/���s��3W�$�XrZ�k;,�u���L�9$��I[�����A�O��*��J!<,rB�.�<w�j0�bjI���y�J����x(��tkDc���J��;��X9��2$�mf8	�uox y�~F��ӟ&/�����ɵpHq�$d��R@	�����n��Y=d��2��bTv�ޘ�f�M�~V�d@�2���n�M�[�P�KJA%Y,]��h�Ư��$���;�����v*�:]�,^���
���Y�6c����,
o�Ӗ��\�5�X�X�%Y7��y��U�T�v!:	��ޏtB��9��n�y.���I|r[q�)�Y_6^9�OJ���
�H��w�{�0̚�x:T���a��=�ּj�E�}W�˄jU%X�X*��<!�*a��%��X�'L�X��V���4�8��ROl�0�Дc��Л�������)0�m���{
��+j 7�&B��qy�?�1�ᆧXCe5J\bTJ������y�&	�)��kϫ>C!v[6q����82j���wi����ǩ�0� ؾS���R�1���X=]Iv8I�.;�I`��T�δ��	�!�7<��I��)vR��9AX�F��D�t6��)~�z���17��Qɠ<J�Ţ62����e&�K#�\et��h^�>ѯ4hG��^G�1�d�M�Z"����[�)�N�n
5+SWrr�����[\2���1�G�+�� ��?B�R�4���n���a�Ӵ<��u��sG�T2R���И\8�?�����#�紋MF���t�ޘ�^*Z��R� Z���A^z�oSn�]�:58g��'�D�H��o-3XZ�W{������X�p�pӤ)DpG��jH�3����rg;@P8�&YJ#)ww0#E� ����Ss�I��e:����r�`�5���"��dA�;=ڿ���P֠�n>\��{��{;�Z��ss�F������ę���{�:"X.�=B�:��`�>���[�M��A�Г��+�����0�Yl�������,��S`n��>\I�VwX�+�_:&C�t