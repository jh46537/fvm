��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{MEi$ �:r������]	��2��4�/�֢T�������A��\��K���i̜���P�G�(3z�Ĳ h�r2Ħ�, 6n��(ޖ��1���]���:��kwTVWv��8k�Fvʞ��	�~���4��K�wS�r+�iސ���c��zܥ�Bd.���3��|�L34���%c�4���HO��iE�u.���.���F9�pFʽB�}��7�n������j�D�mb���jC��E ���qwL �)����BJ�g��w!�Mq�����||�u-����I#jb��s7�M�W�m��F���g@�9�s���:pگ��x"������!- V��X�u�`�!��~�}7����������C�w��;k�:nO�hH�ޞ��ʟÈ�p��|��>��o�:YGd�]z[<�	W����]��ͩ��Lq��n.�Ԓ�-O�i�f�T�WCb^�/u�.S���2^TV���-D�0��z�%��, �vǽ�&�_��X�Uͨ��"�O��HG���7k>TQ�mn�s�k� f�_�K�7(��3��ݟ�=�\Wr7����-ۓ�)�8�1�����	���U&N�?-�\��}y�<�����P�Ҋd�B)�m�8	���^ܜ�B.:G~��o�*	���9�K��5Wh��>βJU��׊�E/U�B��5�������E��FkI�<J�Mj�q �H}1���������1�
���d���S�Yߕ���.o��Ǜ��Ӗ�}I���D���5̌Uf�P��KYk4A����h����&EAB�0�ؽ �A�������f�Fl�!İ���.i�"A8�k�����3�l�Ǟ�'����UP�l/�q���X�ݞf��}Uw�{�ዠ�I�r��D}=H�mY��?b�ϣb����J����P���v�0���e(e�'��Q׺0�#�����	�o������ kD[�|�cYPTB���h�r��tۓ�#��|�I��*�@�M�`LCR�l�w�ۓ�h���t5�a�9�6��PuE`�D��O�6<y�#��� +����B��)(d��9�f��9.��!i����@]��,��%�Q6[�e�R<~ple �� ��m��#!^s>�y�W�l���-�UJu���HX�s	���Ml\ޞ�c�Oc�H"o��=�h���YQTn���m������G@�lz�=�w�{� s懀�u��گ�jus-�X�.4���̴��U��:�&O�
�3BOzx��w* �Qy�i-�����h#�;e��.�^��'4��O�=	���;� ��ꥍS��ˡ���.Ss6���1�#K�[�����}�i�\�P��[�aT�l��g���|���ON��L���ɦ��f~9��q�d�s��|��* ���Z���Ӽ�P��MB��B��c �z�A�X�(�&��3��H<ywێ����}��,`�ީ	��[v����룄�Ϩn����"�L�sd�HRb��[��m�� 5X?��%W�P��l�QS�e���i2f��
�(F&�qL}n3܂�bN7\�C��l%"����3�ɻ���٘q�Kv��m�s+�jO]���*C�2Η�W��a�!�j��X�\1+̸�'d�7n��J��^��*�Fi�^�a�W����
^y��k�B�.�@��"Ә��`i�������SZ��F$��%D�0���w%hOF)W����`�4�ݖ)���&+�� 4���2�3W����*m=�\2�!Q�2|��5�"����.ڸ��l�����x���m�����1������mM���rC�m}�d�j��/���e�"�|f�5��̑eG��}v��Od7��<�AO�n� Y�v�8��}�̻���k�'�f��t�
�"��R�w|KG�z�{LTpP�^)U%?\�v�`Y�NU��ӾU��g3jx΋nܥ� ����.Y�&M(�H��n�)m>���v�F��/T��?jR�f|0����Ќ�J�D����vDk�\�zf�ߐ�h~���k�ȣv%��&&���f!T8l�~z"kG�.K��a��ۦ���K�9y���b��x�J��<L�.���+Ύ��'��ܑ�h�>���H9^�Rx{/X*;Q];�Y���v�ͦ�+��8�>�����'������ӵ�fX)��
�1lAS�����}R����.�?�$&b���Io�RBs=l��:@V�:f�^��{ ?�؊�0���'��3R���A�V�x�c~U��\�3���R�F�7�=��?�0|�l��7�@=wʏ̲������&I�����{sz�Ǹe�H/=�=u�4HK"��P�4��deD�N�^W��B�:�D�~�f�R�"(L�,��z����>�6�
rq��AH���&��n�����_�v U�cIV�ٽ\�a�؅}�bM,M�̈́��t)Q|Ka�����Ę�x��iI;�̴�:Ȉ/Ԇ��M([���N���5�ZSo��u���$rM��kV��2��%�������*T�C8Z�#R?Ae�3B����ڪ7�����l���tdVg�-�c\M�ڶ4ۢf�u\W�Nl']~�[�W��T���Q�R]Gs����Z���p�[(�H`P�|� ���8y�Ϝ�E4'SHRT�ħ�����rߴ%Noq��1\�I��C��NQ&H��V�O�O"W�)�[���7�n�!��}l��A�L{�w�-��,��(�$'7eM�?_��g��Y���v�x�_#�pk�j%"0���2����w�Q����3��uͭ7<ǈ�o���Ҫ`�(�E+*�Rp8���rpt1���0��~=]�������$�0����Ww��Q"�QD����l��u}$� ������J�iRk0|�|��n�yL��x͝�Z�$����JΩ#��y��t���2�I��𞿒D�p!#쵆��X��Ҏ�n���N���q,���j��y'f�����}�O�	��/���'��A
P��4\{���a�+��0X�s[�(�s=D��tL����`�tE�72������~1X(O��n 5�hR�mo��s#{�}6��_oI�撱o?�aHb��"'�wU)��=C<�O�/��'Ѹ�
�ڱ�nJ�B����Ȑ[D�G���`��l&,�ؙl�?��(����xϊ�1J�b1[���4��x��CB<����122MB}�P|HC�#�Q�q������"
�:�d�q1^1�\�Y5�ڑ�^��A�%��C��t�h5�AU�q�U�ڍ�����yDL��δ�9n���0t/�A9�9r_~�q;AoR쐿�'�ju┣o�o��	�J&�1��|�/���Xa��7�E]���%����*�>C!�,�'����@��8�\Ӆ��l������$�m������sƦ��e�!���s�՘�\-�zxTf |���S}���|,JJu��|�Fn
AP>���3��w�4�%o&߱�<Ηz�xq�*b�+�j�0��V�.P��T���쎱W��s�9���e�[���-R�i����u/�-]��A�3ݿ:�kqaZ`��^�V�����+8����a�j(oB)���h�9�^{<m_B��4��4�F���.I�tR(�RثN���f�1��qQ^���\�#�U��i��>��1��<����Pa��U�i�)�������Z�#�F+�w�/i{.���O}�M�էɏ�9�X��&��!q�� f*��?r,S�R3��^�S|�1sf=@ʽ�����e�ֆŤ
��k*�J �w�{`f8��4�)&ng-7CJ6Ek���	V��wg{�a�Z�1]M�X����gO���㜣ϔnǿ6��٨�8����� 7¼�C��8��Q΋sת@)Gt���v7���>!-Y`d[�X�����fm!��*�x���n�����>��*���\���{�}�8Y�1�]p9�Q0,�v��\%M��Ś�������1�#i�-��>�M/��$؝���kә�p=�z�	K6Ewն��N
��h�B�W�
9N�H��]�vEj��"/�ɫ�^F°n����B	�ٰQ#�v;B�˹,������jl
�& �+g�Aq��BL]���AY�JO���73�Q��k�dO�͚���x�:|\}��=^<lħ��x"�G��<��£���}�|�nT��PF	�鎠.ݽ�`��J�/�O���ϻ�0vMs�x�1v�<L��ca�h��6,B'�E��vD-�dd��$ɐ�?����I�����v��w���%�ge��P(�-�Z<�����TH�BdꗀA�LxPxW�^)�}t����"�ؘ~Q{�+�g�K��+|C����a�"�@#��īj��j2UdH����U��������O�)'�K ��T��M�n����{7��O�3j��fvܻw�\��mA�Hx���9�8v&�����W��m���v����m��rID���ڼNm0�`��j}ڢ>��!#�@0y\��B�0��u��H1��������:lBsp��мm�)�n܉!4�*���R���dW�	��twm��q3|~2Ȗº,i��o����P���{�:~@mݼh��.���<h�<��rs%��\.D!�T�#JMF�Ŭ�i�W�`z�� h^R+#�#uh�O8�Vܳ�c����4�f�����})e�e�`�8TR<�#�s��Y������r�a�z�<��-�pi�c:k�+���ۂ5W@}Z��hx֭!�ʗ�Kی�-�U��d���+#�qd�&EN�L�^����#z�TӘn �-�q3bek<�N���C�z+�aQ	D�]H�s���x�J��tA^���.w�s�I�� ҷv!�~j��_ 3����6�wK�
+-e���P��Ed��������8rA5� 	yO�2�o�3�Z��}�W�2��B{�Ř2c2Lv����]L�G�.�v4vD¹��6���yEBC�~�S��vubQ-s�b��(
 Գט1}�/��©��[`���a�8��3�C@I5��{j�5�.��������U�`:�O��U��)�9�נ
օ�l�F:ť�t���7��gi����1a{7���1� =竸6�-��~<Oa�9���oif�����ELy0BRL�8`����k8�.����*��