��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7���:�8'��� G���Ck��s
�.��L�4�L�|szWs��Q�ʮ��R>�n�����_�D9iM��7�KV���J�/��*|���Z���e;��q̍%���_��b���z�Y�!�W��S��Xރ3y1{�/���p^C�T�c��NvMV�Y&
-͎����W�p6��I��¹��p�,�_����ux��R��/�ޔlR�o���Ih�d�;�:�#� 1�TX������~��m��;H�')w�����JUw����CM���S�@PG^z$�j,yp�9lR:��3"P�f㗞`yׯ���@��W�W�!5L������fv2 �S��v�`/-���)����5��˳P��!�ڰCQ�,��M�(��5tϙ���h���4i[��>���U������{�yhOًy�4�إ�N�Rj�
�i��O��
V�+V(3�N�gRjj��=��J���u�^	�t����( ��e�\qӊ>��K6�d���M�>�" ���A([s0;�U퉐����$"��'�����&���8A��1R��w����'/� �8����4^R�l��6��=���jb[_݄5��g/6p}�xK���H�w��v +7E�\��/^�+��+9ֆҢ��ٜ��4&��~�k��O�tH1���\[� jFi��w��y��K͔��nVD���ͅzM�3��`%�T����B]֔�eB���C̹xiv���|W���C����DM����>�gjTS�}��2#� ����t����f�tŵL`|<��g�5�_��Kj�:�Y��U<�i�ۥ�t4��KR�C�%Y�N�c P������kS�I�H��q/Ƅ���"�N�-�L������8�e�@$)��g1����.8��_��?�v6.��K�� ]����$��x+H�53�4��%�qKu.y���:Z�Ϳo��s>.��GC.�+�hh�@��h��&*�2���:�.&��gw#4�VRs^��/�1�̴�q��,��B%ȓ��:}�|�����g>�H�b/<WUls[;�_Gm�V�M<�- ��r�ɘ�^�x�;D���?��7r
�HO���jI��:i�&P�t�&�p����G�Oڡ^:6�~t䙡E�2V��ӟ��=��Pw,�
(Oኮ�b��'��̤X��[�$�rt�T��Q�V�7ژ�y엚���V�x����9z���g�=M|�'�_W����㊴�XaL�a5`��7�N/����$[�I�p<i�@$_o,Pr�NG�b5��]�F�7��$�������7�o!����)BKM�K�ѯU쳓� �ۥq�$��[�Ps�.jկ)�����^^�����0UXjYE�	6!}�%XpL�os��HI�~_R�N��C�h�i�[zl�s�U��kU_޺��G�'��A/�p�U�Lq�LN�c �_�fk<��b��*����Ɲ��q��I�G�� 3h�΀:z_�fI頳�Wـ�J��h&�nX՚�d�v�߬�`�dŐ�el���ZaM�̌�k�&ҿu���[������[uѝ�a$�tk���	�3���J��,�FM��i����]�2�I��5M�P�a���DaIn��,Ky��'