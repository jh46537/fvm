��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[��Y�PZJ�O�e-H�E�".�h�Eo��$w���I+6~~ɷ�Œˉ��r�s���o?#�;���G\�iv<3&�罟Qq���%:Q�q$O}m��ط?7��
����(GӦ�0�ɋ���N��V@����� ��(ׂ\�򃛧'�쾌˃��%#��8}��0O����|�S�P��0�������K�'�����3]q���L{V4&����w�AZ�y�0F6+�kD�d�����T�R\S�c
z8��1������l���\�x�'Β�O��5h��\��g��0������֊~�cX��c}�ZK72W���X��*}HhG�js��9��u@���rG���ڌ�:��3p����8��+�`\붱�a���Փ��;ҿ��h�T^kf��+�,)�ac˗�-,N���׾mS#��Y	�׭�H��#>褍��蜫UX�u��e�G��*�4�a��I	qU�yp���_S�Lg�6pk�'��v��C6�9՟�����`�� v������D5��g�0ʝ�Mu��]�G�?#F�	�'�Y3��l6�M��g�ۡ.�m�#(%�k��Ϳ��}x��*A��wX���vB������H�NM��E<�#G+�S~�=�Q/�W�X�+;���q��	K676;��<��,A�W�sR�8��c��딂�7�������ҩ8�;��)��wA�],���6Y��|�g!}\䓧�FW���Q���y���vmp��� n]-�rX#�#22�s���e�x����
��f�I?B�H'E�P���*�HRe(�����+ҽ�H���#)�i�Ê������h| E�s�����hD��h�Y�g\iH	8���7�7³�C~��!��J�"9�a�,�-yr��w�C6�<��\즡�?��X���R�q�<$ ���B/�C�J�0G������ H���/�Ҏţ�]�� w���'�x�{qra�U��lhP���H'��`��L��u_����cYa�L�1��^��H�3�`(�
��������`w{'�����joQ�f�cۋ���β�Ҕ�WRɾF���\�E��{=�����=_cB�LMM}+8Z�T�>q�����BxM!���Ftս�T��jE2�}�|��@���|&?�2�2Wwq��p�/5�88�K�Ϯc�2�q��=�q��  ���7k~���\�W!����-�H_	��]N����i&��C�tvs����q�o+ֶy�F��׈�]�׼�a�d������A����?}Å��r�Trq� ʱ���4��*hq�E�'��hn�	�ݍt�R.J��b�C.1�5��)��~���/ھ\;�kZ� c	���:�Tc���T.� B�<C� A��=sR�@���ܻ����F���x`��z����P�a+C�@�-ҍ��!M����jŷ?ds���Jt���l���&�� ,"���6���g��	$�%"my�z��uR���E��~w0���r�0����3��� ���F˹`�Y�7�X���:�V}:�ΛE�D�y|�mU5z�����ɝ�k������Y46��)zEr��h��
;��W��R-�6o�~��,3��o-��L�Wl���7a��í�n*�p�y�3�������@
��cH��4 
a��7>r��u�]`'�O)n��s���
�������B���%S7oE&/Nx+�5��u@G('x!��`Y�F9l$�Z��Pˡ�`��h�mq�Vh%MmOզ���j�6����,� %=/幥�K7��
��u�P&ݶ �J��[�S�B�3���5�쐥�$�Z
S�صX�:�(�m�kU�-Y%�#ִ��_�!�`��s�H��	���L�eK��>���ȫ�U>+��[�o�b@W:�X��K����R6�(�z8U5?��/�7y��Y��Q%,>8~⧜��iH�c��Ô�;e+����0�"p��Fa�FV��z��*!�n�i�^��;}3�ݺf�i07gg������}�}�@2�}�r���R�,t٥����XQ�>&V�0��Y�]�Kh�ĵ��Qa9LbK��T^�b;���	j���8����(�� �_zh�7&�V��"���L�Ҧ�:47��D:�6^!�T�؎M�[!�2&*!�^�~ ~�ٓ�.f����&�.]��)e�χ� ����WH��Vv�Ӈ./ĦWh��;��_H�]_}��@E�od�We�J�� ڂ��J{J��E�Շ�L�PWK�!-1�#깦m����0�𰣂&¥5A>�[�cq����+��O.�]��k����)fs8����4�󟠝��"c8�	�1����5��v�S,Ūg�!;s ƦR���s��2�AA�,�����7j�M�,� ����q�:C=�Twv�	+ٵ��7'�0�j4s*~�nlwN|Gd��I9C� +KC�_
����t����>���:�/̳�W��lY���r�(�5��e�w��Nf�⦹#�ɬz�C�Z�x}"�A���ڋ2*֬}�`�j���N��a�g��� @Ƽ� V���m�~��g��^b��P��-�lX��0�w�c��o�%0;�7%�rbJ�+�� ���P�z\�r\=�m�/�VC�\�׺����IE��*__hSNY��jJBj��	iWR�p���$ġ�`��Au�����](��/$pk�s���1��X��)�ӍTTC�����0�rN*�*��*�i�|AZ�h��\_R6��ӷ'C���q���<;>�\}��ž�(�: �B�I���Ö�Jh_p�=L��z��R2��	�p? ��<p:����+(�[h�j�p�o�:I�A�#L�h|-Ԯ#�|�zV�&?�&�C?��8��օs����a�(zy�+�|A��4�g���a��XuLO�-���8aG�A�rD��Ͼ��k����VRXi��)$�#A�T���J��fQ|�K�4�4�/�7�"{�P�G���(�ޤ��`��3{�'O�2���M��uNI�{~V�F�-���"� �Y�v'qu��G���gh������~N��Dy�5����w�bJξ�)ST���v*�@�L�3��ٿu��|)4 �_n�/�P�=�ws�S=HU3>�my"�,C��z8����+S�B֛"��n=ĠW�0l�("�}�ހ!.q;12U����k��n�G�Z�ϘP@�m�����C8gڀD�h�����:c{��^@^��۳鑐��K]�`��L�zC��3��V�(m�C?8ٵ��$6��eΉɧ��P�1o�w�W���T��B��n)���|P��'l��"��T���i�IM�����"��������ײ׽J�B؆��B�n�k�H?�y��R�f
2"��5PP��K�h%W4 f��N0���1�Dw/&:>#큔]�-���&c"��`�Ǚ{�+Z.HX�be,�߬������Y�ne7v�w���Rv%w�8Hg�z-B��-(���H��E��iVB�l�j�N�����9>o:����؟�|3U����Չ2���>eC3�B| v��Q�z%�Eyx=���p=��N�}�65ƙưhPy��~����	�ܹ����٥�SY�j�ǂ6͏��-��Bb|�2��;����Gx8JG�D�I����~זx�YY`1P��e:�P��D�����,��8��v��s����l9swd�����>���A2X�{Ju�V����%�#��ߤ[,���Ap��[�p���(rՔܫ(�b�k�����?�R(&�A�$���K���kS�ڑ��	�U��ah�.L��m����T����ފ^*�s�;�`:�	[-�?�
kL�m/�¹�8gy� Oڂ�����G�l7ZQlRb"��@du�7<���٥y&�;�����K�����@j�Q���>��ao׸�$�z�����B��Յ|��D2�@�6��k���p�,]�aʱ�4��`��뇘�M���wqj��%ʉTs3|� }wK2 i��r�^"�RP�aO��+_jF8������Nj	]>��j��0��Ƙ�z�ͲoЕR8�'="�B�p�m&k� ��bB�L1�(D����K���q���e�o�O��I�y�m���nE��䕁�~��Pt�Vw����t�C�!�\�Hj3-��3L��0�����vk�.�դ�ؚ|{�������0Z�� �a�Ab����4�Ϯ7-���t�h��郝m	�{G�} ���Sb�a���<��y@���������ޛ��^��dP�"8�*���&�^i��HMn�cY~lV6@�]��t�Jo�����>�ClQ���*P��x4�&X/����t	l�X�KiX��� �r�����E�J��g0�뮥c[?B\�4�/��J��:y4c�M@���E�,�ZS`����s��A�%%4����[3�
�~v�*\%���ǍGY�U-��p1'�M����K[�Z���DvH�l8�z M�mb�B�YjExn�:��/�n��1�'���tQ�-Lq_���5Jc���ȩjJWFpi$єDy�س`m���1�i�p�20���� K �8I]m�2��)���$/V���wt��ul7+̿��ҟH�vZ��2q� ]3�M3��|�}y��-�����+O��#��߂�<�R,���@!�kf��1�i?;?���71Lzwo~[[����yy��sJP�<�`�uO$���A�ш�^�M'f4v|�� ��7w��lxp0�zg��NTJe\�\m�耲�]���/��Z+V.���-���B��Q\��m�a���]�.�=����^��+0�Y��m0�F�Ǹ��9#,s;�%&�77����EZ�b�&���������V6X�~�;$
fb�4�1uֆ|�7)�ĵ��r��T��BG�}b���a�h���F�?4������wJ�c��,H,�8��Ul^���W��Q�<����h��?�y�1o�J6gu�+s�j�Mh��D�zZV/�����#����p�HG�7�Nv���Յ��J����C">fc�k�͌��]�T��8�}��^�������ǯ���n�U,�`����"@��
c���d R�w{-2Rb�Q*�-F_�<GGU�U�^��
u5���KQ�om`�TQ9�V	 �JF��8�%/��*A�R�P�':�%�1@�癫���8<Qg �hh? ����O9�;�����Ҝp����5]���u����"�Y"4eY���I�?�?~jGD�g:�E����
5��9JO����a�<�a��[/�Q�l�{�a��N����if������ҽ�-�ml�r5	
ʅ�����}e����?�(��]�r�'���M�lt|����È�E�7���~��]�
�G�5_�kc(����{�G-�&!���1���l�O|�fSFcz:#��@��Ϫ��Hʭ���c��ĄAz�Ω�C�M�R��W�%nի�7���s\�5=ͻ���
5�]U�ZO' H��o��Y3��������9�F�&e���C
F�Y��x� z�ݽ�su__L��haX�-Ɇig��_k���A�3������ª%�R}�$
"�z�m'+I�5���؅j��u�o#���ϖ��{��z�W�Mp�F:�9G;�A�৛�z���8���>��8'M�ue"a�:���\Ls�Z�A�5����v�w�R�9#���X+s�%���6�86yHlU�d�+.�G����j�L�S4_��OP���﷤@�{9��mb
 S���0�B"QT H�Hr�Y�(&u&��%ֆ�9�(M�n����L8�du�Ɠ��ƄN��(N4ؐp`K_B����&BAY��C��П��������usx.����5C#'*��QOe��Zh���Q#���Q�A���|7���ɗ\���"��Q�]�����f@^y�Qp�p7��Uc���:殪�h�=l+��ˆE�܄l`-���!��~E_z&t��`h}��3�9K�@>�hA�פ~1��Z�w��<ܚ�`@�_E�z�CZ���}$���������q����xZ_Z���O�Ya~:�F��#�P>�P2<e2}�	d�W�͖<�m.�4:|*���mN�2̯����Rbk>HK*�_p�)��$u�1�s�v����m�q��/����1pX�a����N�� @k��)9�PR�P�3B�~5*����������GuSl����>��W���ύ��/ ��_U`'�P/��`=���[�Y5�1��w�#��j�*�m���n<$�,��ɳŕ�'��S`�UJ���I0�3�F*ǘ!I��*8�`�����1}��70��_�a�܍/��R�D{�@���F��vt�A~sCn!�K3$!��ǰd�]n���n?%�8�pgv�A������8 ��_���B����Y�R
2ܓ�]�>�������5��no��G*����6Z�AV�J�I2��ULN�e�A�&.�,�����V.D?�E����'+�0���j3l��zX�7}�o���2^�B�dH-ҁ�\3���׵��e�����&ØI�X������v�B�C��">X���bl���	�T�*I��I'���	!~����`�P!{��f�-4~�L^������#\GZ�n�xp�P >s���
t^.��k�*��۴a#�֖�U�y��0I�m׵�Ж��+OB��euw�Y"�9���oY�8}���A,=���j�MCS&M�3�\��niZ��{Â�Z|?*� ��|N�����t�e]ˢ�/ӞN��+eiZR��u��.��(�?��4�M�b�O�L���{�4P�@R���g��xmPQWq�i(�-|�x��@������.f������)#;׻h6�#8/�kxy\�YȺ��zr�@D�e���\e~�FI�x���Ћ�ޘ9�"6-�E�d���e�a�U��+��[��A9��1̯i�Yi�?^�gn濷�reu'��N��#B��C؄-�pQ�]�c��@u��S9��ߟ�ʢ-m+H~��0��,v,H��M���P��������P�V��F<ۅ^�9�����M��	Wd2?CѨsOA�ΰ��E*:b�W��L%�G�^���J��(�����~���в�3�br��B$��� $�P@C�������U kQ����	�T�S����D���ʌ���<�z�w�->����.��*���B&Q��a_6f��;p"�(_�����74���������*롦��O��� ����c������&*0�Gi�l8���T�����֑�˧�l�֩J3j)8.�3�Ŷ���T����u0nu�6���vz٘��A��+^7��>#E����6:eNϾ<�w��%j]3�G�����E�E�?���>|p�F�s�~��7Cٲ��"��fJ#M�&��ػ���;�=�}��J��(���|�����%.@|��K\�[ws�`��V ��q��x�`8H�(�J$A��f����pؒΰ�r�����*�bK<���l���*t���Jo�t�(����%������|5֢�/?-�rB~{�eJ��w� d?"�2���ǟ=_&���ȍ���/N�v+}����*-D+���v(��V��39�@E�'�v���҃��1u���I������������o��
�\V_�O��۩�0v����3�q�F�{�4vĳ�Gzn�"7�5�s��0o-_]��R �3��3%�g)�X�>O��mD!�ϟ`������iT3�J��FS+s{S���+_]`I!Q��6��b�ǫ1a����c�~�
]Z9g�#=����)ۯ�؞�����c�q�+kI54EB1�٬ޮ �(vȧx�nI�1����>L��A.�����Ɩ�z[�v�f��o'Н+�����RJ��N��!�+��V�i똂��^Ȝ�tB�0�V�m�t������^�Xx#�mnܛ�t�P�;X�`6�>Wv��*����i3VI|�dmH�RU\���\��#Zx��SŒ�o��"�77 r�&	��Y*L/	���\�<g����Y��f��wb�M�����~�L�9�zٰ|�y�d��Q���X����J=����з�t��{�-��
�!�]~�0�p.�!`�K1��KkY��5���
���
<�0NV�Ʈ��SQ.c���g�H��45rUJ �Ȗ�ļH�E2�6j*�J�ՇhԼ ���1�A]4�B:G��M9�0в��(]Zeb�`L���(VX�?��gs[2]N��{����&B��$:x��W8��x�:�`vF������G��:�$�9�p���=�*V���u���}?r���Q)"lws�DZ����`�[��KX%*P����ZoZ�b"��m��M(zD`����v���fQ���*z���la�8`��^��Cp��L3FH^EOl�P�����J���c�*|�;p�@o?�EB&�,����90��q8e�v�5?� ��!�:t4�`�~V��u��˥i�e�<�/(� ��Oj5�je��s u�y�d_j��R����M \-��M���g�5,�B�����Kz"e�����XX��<ij..�'�T&~�yl��Ϳ�WP"O�V� �QjLݮ��=`���^��ah*| ��w��XL��>�y���e��C@3��y�w^I�:�����'�BY�^�n�@,e�3��I�o�6����6{��#D�v1ώIu)gb/���PX���� ��^�U���l���R�b����S$�*���nTM��L�lIv���[����Z��`c��J��N�.0��־�6�������"��7C�s�i���lw�NT���TЌk��(�����ٲ�>o��S��"hsV�4B�zX>�����p�)Tk�g1,���u��{h�����I�-���0��ql7��J����]9X�$�/f
r�OGEya\�<,���C�֚�N1/pZv���5��.ɻ��<����r����ku���T��+���tn9nq靶p?չ�۱��F���ϹZ���B�1�Ҹ@�)c=5�	�X��AV���s�RG.(z@�\�шgw`�)p*���s��+���p�@HY����R�X2=��Z+�kZ�|;�݃t���t{����gJ}���X�����/���X��^po�A��Ze�����)��&Q�����c_��[h��H�lU�S�u�{��W&�v"n�>�m�e�%	��i���L�Z��t���J��8ψ��)�)S-7[�����m��h���,��c�U�*�l����:�B�P�4}�!ԏ�}(N���Ns���Q=��z�EP2[�{���m��J��%���k���(d�Ulچ|e���'�[_�۟)�Q#e�i7��?1�l�e�%��5�i�@� 
ܕ�Zbl}�ЩͩnDwi��Eh�W �8�l�?@��R�٪/�820k��_%�-�����վ7��2�ܙIvQ�����S;�QD�^��
o��]~d��.�P6�?e�p|H�U��W��()r��yf�JG���C
qX�R�zE�鮘�������v�kV�=Y����>��2+t[z]Гmp��{��0e�9���^�ٯP�o�y\�������G �H�\)�%�^���0^ȕ5w�C���&�A�	��*W�Z\�M� 4�H�u( t�-��T��Eךu�(�Y�/��	V�^�l�x3]qN~9���	��'=�1=�<�g�Rk��0����H��8��Ac]�w�h3)f/c�216��T�����r.�{!��I\-M��}f3.|�$��
�V����Ò��U��g�MG0)��L��:����*#W��~(�c�)6�ly.À��Q|�G�bm��N|�kӛ\��i�j%�W+��
�z`a�����!1��ʛ|��F��p���3F�����֫]&�̈́k`��#�(X
	�ߑ���ُaE��״�QG9`�)Аɣ��y���!��X�B̠:�B`��-�q�uH�{�k gF$&��k^ж�tG8mЋ��w�U����~I&��6�d�u��TC�}�(����"��kzq<W"*�8�S�A�Xң�w��ˏK��%(��lGcN�qD4�g=�na��flCO[>��
�풑��e�&~_��2q���r��pe��Јo�\��g��YWcl�������|�t�!J�2лբ�
��6?���q��Oݫ�-,IAr��V ����^�	�|���ZVkTZ�W9����1�e������������>h	�"�ύ��h�J`~�����A�����fYU��	m��&�K�ww"3b_sЮ����wl��%��<$\E�`3HMc��J��
����W[)�nx��Ms������)�?Gku�!������OS+��w�];~g���}�{��><t���-�	���sa?�����iM�ېm#mH�9If��n�N���K�ԝ����Xq`!j��1k�T��Ԇ��$q�oj��?_�-����'�*̯�a�m��F����!EzMò�PnM'�f	C*����j�M�4�ـ��eҖXl�MI�9}	Tө��~��R�זi�+�mG}6O'GE6'�K�P���*���S���*	���gC��^���0b�%��,�&`AN�I(��m8���c
l�1�r����l:0�;���+�6B�.J���)r�����Β�u�'�#i\�Z�!��?�J妗���V�A��<�a9��x��:Y���b��oIgrJ2�8��X�	���=��ұ���ů@��		D��)��C�#-"�u�Xָ�J٠ޱx� �HT������6C�^j�*f�>@�p5m�7�UqǺ��"}��ׄ�ŖԔ�Hv�*��.�Qv7ղ0<�oh�:�1>i�mj,��uя���?�r���B�"F��u(��*�;��0�X�pT1��}�`�W�$INR�A�L(@�3�Պ��&�xkK����&d�{w���aߙ���2�8���ۭ�Զ&�t�~��J�7�ЌɎ @r�q���zLq�Xs��+�Lg(���O_�F
�}"��x�c�>��P~��wH053�_wDlf@;�./Lj辶`l|�<BO��?��iT�H�ޞ\�\r��3�h�`D��d��̞��?�4�C]$w��(���Rي�\(u�@d�I;5W�f�$�	��+ �C0r��?N�����]�B�=��o�p��ׇ�}�|ϘJ<�h�~vuJX����O��1#K�iTF�,������hD�A�ǳxj*�Y	7=ǪR��bi����F�t���l{T�6�1o��[�@Q׋�>�-�P2꣇�ۙW��J68���wT��}p8
)���	���83Ww�2q��^����<j��L5�zUu�en�=&�V}g6�k
��k]b#9&GF�����
�p�l���0�ka���m. ���_�c����nA���@s��r9Dy��{a�q�ºN�V�F')㳙1SQ��Jd�*�B�OX��E@:E�:ȋGR�J��@4Ň�Ѥ,�<��{6�X?�uN��Ɒ����QYB�������-h]�7��J=��b�7��6�Pqr�E��FH&��RÛk H[����.'�MM[Ab���b�$�2W)�N���,�3\L���>a�:es)l�J��$�q��t��L�T�1I]��bI޶}C'#�Ҙ�4��<�ҩ�
֏!��pk55c\��Y鬬g��b�~��`�H��갠:yP�gҿF�&�"b���v���;Vu���4����<l��Z��p�EV�1�h��4�N��J���P���Y+��H�BӴh�qk˛���a=q�{Ge�44�ft���T��gi96-��/��5��|K��8>�4�e��  �"<��(�/�甃�v��Z�}�OK�u�8�6��dI�:�
fV��(<���'�7�J����`B&u4B�1��M}E� �C�kO((��>�2�M����߈9�*nJ*�9�#a@�菭��v�CܼO4����S����I��E(�������u��NWo����6@o��~�a�!���h����вӧ�������x�����)i��)���N�/�����v��!Th�%@�#7D�1��2�&�b�v\�{��L{��Ur[��_�
�h��h�p�q��P�[�/q���Ҿ�Vu�|�����Ar.�A�.���hu�r�=�R����Н��u�lO�#�2�/��~X�����a����t�m����<0_�.^���ö/�H������݀Qw��zگ��R�:]�x��C��Z����Ad