��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�0�w׍��SΪ]�����E��>��顗���="�Ct�QJW�����j��I�����1��5\W�(��3�D�a=Z=���=�UK��*-Oᚄ6��f9�S|�����Sw-�����R�42��a��ο�&�L�Н>m��%^���8L��ݹ���{���`E�p��-�jq.��>"�H���Դ\/���_�#-0�tX>�K�uT��<6��Țs�U2�H�|���GDN��� �̛�al:�/ ��>yx@����_���tq���,�!�o��j�(����^�K5�򯊠�.W�����hط#��@״�`Xo�ۦ����
Z'���-��'�r�a�&n����"%���#4�{�^�#�δ��tX~*v�/�rLk�� ��MWv!�|�IL�5r>guLjj�Q`K:
�!��=_X]W�]$3xNp����h��a�+F4`'ȑe�5�[��B�!�]���9�&��W�ā\� Y�y�2T�`�B�������x��5<st����, m�yi�E���#ְ`�&K��p���3I���M����D�ш��݈δ����E^�-u&����9V$����@*���ӌ�Q�w�k�
~�oy��˛�Y�R�y<���	w�E�D`�-D=y���qG��2`Z���j��������y���r��+PM�ڐ3�x���� ע���B�,e^@B�Şd�-�a�k���}��M��0�V���ܼHh.�x��Ɂa�*Ե?���nz�HA���y��3[�(�����"
���h=�E���"��&��1KoR_+c Su��V�>^��	���F��:�|ɨ�Sw����u�%`�xF��ܬ�1����ˉ~�+�C�E�zAas����TH�8x9��ť�tp#L٬�-4���i�A�-�%G�U��:9`p��~���'3.�N�q��͉�WJ&���s~���+26�����2����#(J�@���{]�s�U�X��(����ސ�BQ��0ޮ�qQQ�-�L+Y�q�� D��|>��nٹ߿���*�?H/�hAj�� 6��Q�T����O��W��V���#8Q�ԋ}�"���<@*&9���{dV��"�H&���91N�+雽:H����_:�J � �?���<����"6�OC�*���V�3�R���"Sf�aM����Z�(gr�e�*6^��_����	��*I͆> ���M�_r��Q	�߀�(���Y�Ŵ��|�B�C�������>a��}��m�XXr>Hm��8}q�&ǯ�0I_���y>0�S/��g�&���UP�4O�Tˋ	�)�ٳ"�(�E�Y	T���Z�s�l�-bh*'���;���GAGm�6H�z���0�"�X�&�w��gE8b4F7Xb������Dq��$y��Tq���KK�w�X�d��(���Q���|��ϐc�z(S�ՔK7��|r�y�B�,O��-��̙�?'�������7急��ڎ���/��mg�L�6᫐��S��ơ���E����5�������>�u���v����F���x�@��
���7GLp�e�C̦�S͸ꉼsm^�UEHI�QaV9{Yf|`��$���A��pR�V�˫�9����8�w��J
ES�P{6gtk�!ƣQ�Ԧ�6���IJ�ɢB�fU!)m��<��9Уz�8cx�jѬӺ�fu.�=����A�ʲw�X��<m��{�H+�n}���QQr�c�(��5��pkk�0I=�$�Xr�M,?��!yf@�#}���eÄڟ�`�}��<G�[��ۜ�خH���ĕ�^ys��ŀy��NĉF�<�b�S��_�cT�=1���Aq'��$� �%�8��+���/���H�x`�xo^$0ظ�=�&GoZ#�� �(PO~F�i��0�����T5��I�E���Y��b���e[2d��?�Lp��L���h�wm�o�;����e���G ���6Y��.`�xa9���be_��(W�]�DQf�]2�sZ[� QT��jN."�����C�2�ZC�&a����Id[#�J�����f�� ��*|~�ޠ�y�&'��)#g_�ڼ����؇�h��B���g�{��5�Y�\��F	���25�$��f�I����T� hwyO��;���lS!��;��,�>q��Y�	Z�I�'ؼ�ҁ��a�DD��w��[`�\�F��YŇ���A�����ܟ����@AC��a�����w3��`�5��-�;:%z�mŎߤ�����x�II�oKM[�G҆����w��n <>��N����BF�:�\�8��[������&C]�~��V������2f��tp�h��^���KlhK�/A
��zQ�9�N�����Pd��#�q����w��l�3�翭Q�%yw���9N}Ό��mS��+�&Z�ț��?�#g�O�:A=���p�jN#��Gc�S���b�E�	`*�	%�	�}m ��>/bn�T*KFYP�C$E����J�3ȸۏ��m�}�RL?J��I�*h|?�eêS��#sf��� Y��`�����{�,*Rǀ�3n���	#W�:�7��×�;QNi���+AN���X^F})�t�y�_:^���q���H�a���G�K�N�O�]�ϯ�
��4�v`(Z�t!� �غ����iv�0�d�d�{`M�vi4���j�5��3	
^ٗ�
i^�P�HQ� ��Ps�ƃaQ-�4�4�@8��J�*��*S9�;1��`�w®p)�t���ʹ"�r>O�F�(Q����k�W�oz����@��$8e���DU�],��&�u������S��ߐU��`؍������c|��ٔy9G���@�0_6m�ڮ��|8�����`/҂Au:d}����?tq�@����/<@������O��Ӎ�:ji�WT&�)�5����o�Au0�k��-���R4�X���	e�Gx�Sq'�)��4_Q	抴:���<����\��F����}&��U��ɂS�v�Z����<#!��>Ӽ�=���ʹ�i4%h�WANQ�-_�e5<b��0 vL���f֌3=E��J(4u�_��w��Iz>I�vۗs-=�$om��ë�Bu�@P3-������j� �V��䴺�o��@�M>�Wk���ȹVjb�,��C��(µ�sDz&q���_�h���(��8�tç�	1���j-�;4s���~�;�1E'�c�k���X�D�~���N�;��@�����\�p�Ѧ����%2*d�n>%��`!��E�{����V�j��&$�?�{���p7��<��kn�p&ņxӠr�4��O�/r�����uJC��A�²=:?��t���D���G-�W ^��+J^����h�H(lՀ扗S�,���a��\�z��)�#�Leڷ��*֔��-~�LIʩ⫠�8�_�J�7Qf�>B�f
S5���/����F�%..��A���Ȭ9M������*4�B'�8O�Y��Js���#7s v��v���8��Y��x��î���-Z�Օ���n���	�)�4w@�����]�X�<�S��"B���ODEg$I����Ke�r͑�$�=k�Io<I�0��=�JS"�9KɊ���L����O�% 1�H'���]-j��Sm��	Q�i>�K2�O�nch�5���/v��,��SM y@'�or�1���?׌)}ao�昼��l~YD�����@�W0�6`������� ���ѯ#���U3���4�Z��c�e&��fZ���4p�^�W����M�/�%�s^��1U�H�0�ąę��JM;&p��&�������p��O�r�Q�����	>��ީ[Qr��Y˵`��OE�"�y*-��;2��^btI�6�\�`�9�
{��Ftx��� ?�*r�3��+P�"R�Dr��������F���Y@]:vA�ۓ���/��J>���<�8����ӀF]�%�l����x'�ˋ���=Ta\5sC(�q��ڌl�R�"t�/܅0s�\:�V	�~߀6"�Y~��NIF&��4艚� �$K��Ϝ��Q܍�<۝S���7r�kpwz@�R/���!ך���_�)V��Ю3q��~���`<Zw~��ͪ	 YߖcV�b,�;&����;�F��#��cT�ش0^S�^�i9�#r�L	���ݟ�$�1�|{�+�7�2�UE��� ��8�����BYmֈ�V.����a�	7��x�KA~*"H�C
��=�:?Ek������PIr�*����Z��H.ݗ���ְ�����2�^ӹ��8�&�pz<E�$�~��W���Ӗt���b&{."�ͭ�sW�_qڎ�]�G�ޣ���-9P�K-��q�k8s���M�$t���$3�y�K�7�~�肞ӊ�~O�q6{l*�}c��� ��������m�cxs֊t�'�nZ�D��ɖHxm����3��]h��uJ��I� Ż˦WF��e!���҂�wi�!ťoT�_�_'Wr���y�V� 6H ��4�D�x��)�Òֵ�u�	������<Wh��<I�Ppc���+��B�N�6�ۻ���]�2X���2?�&�!��K%sɦ˻��W3^�j�Q��D��q��^`�C�R�$4���E�[&����鵜��6���q"� X���G�G���]\`{[m�N�5��pv��^��K!�zP`���.?���5+���c�Q]���OʬM���O@Ov	�!�e�ĵ�<Ƿ���O�z�����ZBs��FHWʿ�,���85+���|�$��8�#%�X3o���A����T(�3!=\�$ÐՐ�S+8+��{�,�x��n����'4Bb�О\�_n]�V��]�׫(������CCO�q����3���Ȁ�ݰ�u�W �����D/��.ǌV��W6��Ԩ{s2���c��Lي�:8�⻎���4
�r{�[����s�cq�b ��|��s��?�#<w˕��v�՛Ϡ�0���A�i��̆,u��Jw8�?6ǬB��,�{��";��x����M�_���a~@e9���!?�t���l�9ܖ�L�Y��U^,�⬅�v���dNd��S�e�j�}O	?���ԫݟ��7F�*[�X(�(}�1���@�qYb�9�����I[h��dP�ǍR���`��;mqP��ˣ��|4Py��A�& ��f�%�ӏ�x:�q:w�S��>�xřs��å�V�9�@L��w�cwuI
��6Wb�'S���u�#(�L��]��oH!�u��|7$"�����_�BR����e�N��Hj�9�"kE��^�s�0���xQ��-�`:Iw~����8�� Q��{����έ�Ӊ����8���x���u���oD�P��}I���HP��]6�Vk�EVNڴ��2����o�'���T���5{��v�'�̶x��'M��(�xCN�n
Մ�pz������'2� �}��6n$[8T�)&s�^����q��yFw�"_����KH]��j��.F�>�ϰ�ӶJ�,�ЬFe��뱈4^K(<�!'��t����4�k��F/��ox�>#�ZB:`8�5����n<�������F��}%t���Ϣ���`����F�6�M��'�٫����1a�M��������X���U��:����c#�4��q��ށ]��w��a����� e�%�AoM_��&ĐE�nR# ��{CK���D�
����.ۙ/�d鸩r�gx�m�L,��ך{��n�� }8��t%hU�n���l@R\L�w�3�..2>�����z�������]r����(��ҁ�Sc��t>�x��;=jr�w�᠆������F��7�ӚH�Py�����.Y�d�)z����<}ߘF��+9��)#�+gp����}3r]G�����D��ɮ( �4��5���4�qВUw� ���H���O�8v}1�/{���5��W�9�Ԙ`��2�b:����D/��{Q�te�#̱`pUI+���G����[�Q�_\�^��B4R�8<��Bu�U�U��&$��\ ����(��&)�Fb�hgh+RGOѽZ�u��YKE�abcP��,�Q;�޹I˓�zl��b>�u�o;��9�j�`�\��T�&Ԇ�X�M:��ɫ0©!��
�E�y�f.֜H��h�4�4��wk�����=��ؚ�,�ڭ��R�F�uc���G�T~���Z2� 7&��;8j���  ��1�{����
R��n=���!�cL�<2`����*����~Xl�E�0 a����2,a�������1�q��f�|U�"ť�u:9���Bj�AROKiw�]�Ҏ���O���`W���|*�Q��mh��e)R,6<	�-����?}��HQ�4�j��s�L�(�!�j��A�cG�v�՞��`�&�b�����U�g���`�t���=РM̖48��,��K''��p�h��]��ۚF�[{ɻ�z���O�$�F��������MF���3rh�2T����-q�}H��)V���۫m��6%ρH��ʈ�O�Qc�e�;�ǁ̝}�i�*ƣ��{]�m�_���W�䠮'�@]����=���i�\�J���N����kT�C����1+K$r-N�c���'�NK�ڠ��@��J���h%���9E�j�|U%�Jx����+9�N�35���?[�P� &��O���H��:'�_��� v<N���G޲�����E��{��n���	�������d+jg�x���+s���߼�Zv����s��;fT*bϳ��E��~�m��z�V�Yo�V:z%���Ձ �O�<dG ��X��zK~�h��z�?Ʌ����ڳ�p�4<(g?�����t�|p�8���T�J=�+��<1�|�:�#AE}���l6X��B5��5�0f�0�W,�k�����bV햣���������f�$ y=N�(%��<�ij@\uS��9�v���Z��9�/%'� ��_��[1�7Ɨ)X���������>���MQ4���܁����؛'%m���vd���ܥ#�~�-Tr�3<f�%3�z�4h��0L��x}*��C�敀ޛ�\��t��j���$��G%��hȋ�j��L�<��J/f�iK:�n���d��D6��$��Jr�B�tD-��g>զ���˄����塦Z���}���kML��@fq|}-��:�v,�9����$�tI8;O��5/�G�byc��wP�1�1(�^qf���G�][�H������F^��Ztn)�j�"���2^��؆bf�4�8�nK)̕w	�f#�Y_K���)(�9�@���le�u���3VO��`�,�1�������UP��;�1a��Sv��17"�=�$�$���T����#�4�h��ݦ��w������2m�IL�x����b�K4���P�YCA'� !��G�G �MlJ@��=A�;����s��	������ ����M�u�&B����Ό!p�2O�0����oo���&���� �s~��ȾE��d��?���_H�G+H�����ȣ�r�nLU�a-���6�6+��$l8�; �8R��pw����6��A���C�q�J>�7!jF��z�H�?�z��~�9gؐN�fk�T�쑿���k�?p4pQ�Z*9G����W;��b��<��?�j {�y�gG�Gt�j�c�m$l�e�}�7��W��������Ɉe��Գtw㨉W�~dK/Qk�ye�À��I���pI�m�r,��͚�n�y�2�@�&�f�V���\�������ԩ�F!*�0�!/8�jl�<�`�K�
M���;���bIn���:YN'Fl ���4 �EG�B���ö�>gd��;dxtװ�ۡ�p�u}7D>��Wn��[[#W�A�I)�=(E3q�Qy�P�:N�
�a'��U�{��(ѵ�/��u@��x��\�L11��a������0������e�g��5I)�H~�%�g�} �hKVha�nb��u�ڰ����g�3���r�P$ta�(;�y7���#���$�c"/�.5����}���}3��:�j�Y��&�{�Y�W�ʵ���M�d'ǡ��u�L�
n���"U����W�`��!���2~�MYӼV��Z+3P[�Y*�v�u��{M@��M��aɳS�U
�� pi�IK0t{�D�|C���j��d��*e:�{)�=�w���e��R�m�i8u�(�Z��(�v�:��_��{�2m)M��vS����|����RM���K;�����o=L|=ˋ�
d�mv\�}��cMse.�4�U���z�>�L�E��t%\��#�mdz<�iQ��a����!�W2�����`���H}�T���u�d0�7@���Y����`2��fE?]�y�2�%������Ƣ�?���7�ீu֢=�����*�Pe���O�!�u�lE�UJ�y����u�w����!T(G�\@!{��f�$���{����ñR�g5�x������E(),��F��1�(��K���B^�	�9ڋ\�qQ�Aө��/Xv=8�W�?fLf��nu��տ`L�Ȝ	z�r�+��?-x牽����x�/[k�A�5��O�Z%���]�%,G���ɫ?7�����$����w�Z��h���KNb��dxd�TyO���F������1җ���L��1���j%|��ofV�alث����ڿ=�O����"���ya	��&���8`�d�k�@rmg��%d��xY�m�0�R%�zd������Y��s�]r�od�L5���$ơ����U�K�ezp\l��d�'\^;T�й.�M}�F��H��� jLw����A �"�Xj�2������]�=Ą)��5ڹ;���Xy���pH:	�F%�!W�;]�����������#�������DW�Q��Xg֐�FY^;��T�/����V�bց9�	 
E��ԉKf
��D���Y�:!I3�s_6��� ��<Ռ
B���qeI��n�75�5@'
���{��y�p�%Nz'U�(�͂["��hnivH.��0� �5�����`"�S^_U��c��أ3�<e�{k�iP,}�B��ҙ'.���� ��F�k��il�g�&�I+�o���!���v���!TÞN��� �;h~7���:ą�1�b+V3�y�Z`Α����r�f�!�����*tjE�]�<�Όg�ӳx��;��.�N~8����B!�W"bP�<��!�*E7QY�e?��B�W����x�Nzݱ �'�<�`	��#nz�I���c�Uh�Ա��%dq|M�'�|d#�
cAëuBKOke3-�c�Oq2�>G�L!��Gc�N�����fmd=s�� �*�[Xbh
莴��D�	�ž�Z�p@�?@@�8��M_Q�p�Tlg�J�MvE���z?�,E����{���T8�\�z7]u��6�6�`�_u�j]�<h�kur"�P�V%��(A���̧�]7��4j���Dz������㾤�s��`��A��J��2�[�bʄ�!?��AM��@r�
�e�Bs�e}#H��Kݨ}��!ɕ�}�_�q��y��mu�����b���i{���D ��*e��T�Y�����4���]�����A��萇��6������'��7X::��A�AIz�}>��х�䫖=�f�37
��v#�A´q.7 uWv������K�� �xM���Y�D����ψ�ЍT�a� L�W��}IM��w�e��H�(A	�t)T 0��d��x�dؗ�%��K��/�c���E�R��)�۹�Nqx��R����$���˓u�{˺4�Y�i����S���G�)D�����]�!m��<�d ���"�B]�Lߕ�!�G�3`>�cS/afo���D�yp���M�o_-rլ孏\�B:�/Z�p�������*��W��a3��TM &�]S;5[#F����W(*Z�r�{��oE��-�X���i�-Ը�㛡&�	�/Љ) �V��EO�����TͲR�g6TɢQp��a����0r�k4���(jЬ���O9-�о���W�kD��2$�(Z��pA�XTb|!Xp��dI?��u���}������N�ǜxʎ~J�����类�b�������I���ra ��������� ����uɻ���h�(?��s�(�u]XU	��Xo����2�U�T��!>a\�FȰ.2u����TŚ�	QN���?Z#i���sCZbt��X���x�=�u+k��N�6����f"��5��:m��X`~^>+TLcBDս��q��n�"\�Mc e�h��~31 ���^pC�ou�q5��V�Wp/�L�6�?��P����k�anY@`</W
����o��(��e.��¿�uT�(��B��/�4����7�}1NNM���R��R��Q)mʻbE��H�K�?����*	�}�4�аA��}�f@��S�?����6nu-rz	ڣeR.�SBrh�-]?���
�D}�l]��aY}!&hƢ�Lup lS�O����#�$�����D�	�}�j�W�Y���<�u����Ս�����r^ Ų�H�F+��y�D���D��I'u�O��B1�4�k�ΗaX�n�ԙ��Է�f�^I��"T�l3z�S@)�sk	:�rV]g�B�E'�+@�$��W/T���J���+jF�V6zN�c��y�J�SY��H������N$~�_F5�\�G*h��쀫
�J��%�QL��7հ'NnY$`�� Gs���_!��nȈ���:�A��%A"��{2���n�=��Jk�u=N�5=�o�F��Sq����m�;�[��,̎�Ɋ��$��4�T��v�Ԙ�����,��L'�S>�����p���d��ˬU^m��FF�U.��S*�:ϥ�,�ά$Éj���Jd�Gu�8�E��@�#���88�.v���z�}�GmP���mb�D{Arş��!]$�z8�P��d����ԕ�aغ��k{BG~v�!
�o"IZ=���$Y^k�l�
�<��r�J��P<�$����oyk�~	I��HC)��)�Tu~��� P�Z/C����Β�^@���"ۥ(Ƭ��u1_[˪E�0�Y��m;V>F561o�yre��d�y;�j���ם��l�Zʶ�q�=�e��4���9l��3�ʷC��:�l��-�
�j��[�������?��k���?kE� ;���F��{��ED�ڈMI%D�e������ݥ5��m`���
E�_B�'~�q��Nk�Y�9x�Q��S�SuG>M ��6H�.YAB0���/S=g�d��Kt���������v*RH�ݹ��r�zQ��u��t�At<l�u�����1P�l�/+��h������<�y��}��.�r���G4ɡ�LD�J��7=�~�e�;��׮5$�r�u[i�b��_���3�HN�M����͢�p*�`~ǪD���䥄
XrF1�������$]0��0I��Y�X~CҖ�$_4��Ky�J�s2QԼX�ob7ַ8�<;
����2I����ɜ�fK����������ڽ'����%���W�7�q�K3e�پ�|0�jwtׯx�05e�*e""u�*<�I�iLԤ���y�S���f6�j?�o�wm)PpN�"k4��a\�����"}ʺ:�)�}<<���\=��r<��hRc����c��>)꧊����J[���s��$o	R~��ǁ�8�M�uG� �M_0��Wڙu��6�n��UEq]٣�'X��Vl��x������%b�x�z���k�-� B��B��ܬ�Cy���S��f݆[}���2e��ݨ�T�+lc�{a�;:����x�z� �TBM��6�{4��E��v�˜a�A� &<c+�T��݌q�Q�0.cR�^�l�.�~a�*ţ	��6:�1W�?�R�t��ь��H�X�
x�ר�����U�8�x�:��lK��J�u��yT�x��'a��|��#AmTJ�����;TD�d�j�5�*H<�.M����k�ں�i�Wҝ`�;�su�2|�'K7ο�o|<��*��c��8&������eK�`٨�nc4�~0e}o��(���JJ�3��6�49���=���õ2�=�L�A�B��;D�NQ�ާ6ߗn�CƄ�W˚[M7i�q�����mw�����u�fe���p-X�����]9Q�'f�R�դ�E[�<�Sz�{��{eΏ`W;��6Z�ϰ�:��z���:����5�ӈCs�\]rА���5J���|NF�ʖ�k��>�	�ѻa�����ri@!b=��\#���ϖ*��>�[ �}�yvdV�6�<��DЂ���݃�.�q�+�zk�ʜ��`���E��_����m�=��Rz���5���mkQ�:
""[�^pS~��}JG����	s����(y���hv�	��^����!��Kx�ss�xÌ��"�(o=n&�-�e���P´�IP�3 ��\�?����q�~����)�?�D׿f����	iPZ$?���A��A��f�.�y���5jugn�ݛJ��,\���o�ْS��#c[�j��=�[ˍ8/��6���n� ���uy�(*���"Pi;�~��w�S�rFPȕz '��Q <a���Na+�s�6c�3]ȭ�sR3��!!l9+!?_|�r�M}�p$a���ϫ�;�f�$!0�F.\\/����3�j�n`4\׾h�v&�n+�k{��lz!:XILy��t�E#���솶}i��xģ�!�z�*s��n�n�V�%r�Ԓ-��B/3�r��&��V��I��A�}��m!)9�c��dU�nR�CRS�,�7,7͛2�[['p�v�Rp)�c�p�.d�.��ϖ��a��T�������_��Ը��0'=���-�}`l��x�Y��Ѿ��@���1��*�Q<'�eI�B ��g�ʊ�V[R+؞T����郌��x��Z��~ ���T�w>뀕�c��d�X���K����y�{�(m4i�qK�����Xߚq�{G�/�����H����PB��p�GZUXO�I'E8N�A�z�^�2h���-M+�����_�Dib�]��?$���B͆��ᜫs�I	�8�Ӏ��B�Q��c��=�4�G�+Ti	)��bo���^F���'����8 ���?�+ɯ�0؂6�,G��[�̜���r�i N�u�']���Zj��O_&���g����
���O^!W�k��G"	��8вH��9�ؤG�"	ZXk�I��-ʩT����!l5W�P�$w��rl�Ϋ��}R��L�~@%�\���P��g?
	Ah�g��+�w��X 
�"�?{�ۆ����$�a�i\��z�G�c�}�P��y���[�+��B�TOdM;���>��`�'��\I�"@mDw׀?"�{	��M�����Gh=��/f�p���Ac@�\��{���k(#9��x>K!������fcTR+-Q0��7x�Y�z��3(X��{c�*�O��/�a�U	�@�X٫Q;'���� U����_%|���]|�aǵ�������C�R�3%ux�CA��������g����'E�ͺ��>yH��A�V"�Ͽ۲ؗj�N �Xnu,@����͗��~�u���� �t���Gn���c��'�-��Өu�Z�UOT� �q����j~��tʙM��&l�1����n����q�	n�������rћ��k��s!��;�e���[�ڛ�%+J}`������G�<�|���<5��RF������,%lSH��M�z���6�kGe<J�="���@���ҽ�/��
����l�߄�	ӡ�#��4������α_����<5&�/<���YW۝!�?aHv�}�Z���a�ۃ����
a1�񎩈-�(3���
F�32FMh�RN�4��
���F���E:qI�7�!��yV*6?� P(F�P⢇�zl}�3�Qs509f�P��5�$�^wf�;���(�#��d�(���a�v�������T��w-M8���0�f?@��?���g=���*�~�fڒ�-��"G��c)���� m�F��NB�}rʶ���Y��g��n�T�"5lHmWe!���!��"��#lJ�Ï�o���>�#ޙؙ�M�R����p���8K]Z8 4�7^�n�30����I�����N���;�G+�W��-��A��j@A��<��!�.�d/>-<� \o4Tx�iķ+D�1-AȮ����u���9ySF
NP�G���G:�����!���sc �Bn�s.��Qܳ��pf������	����]���w.�� $���,Ty+f�Ffn���0!�+�">_��|�;�I��(Sa?|�h���K����jO���zH��5�l2��>yB �5�E����]�w��,��(�_)�ۻ<��O�:�gaձ܇�w�^bޮ��w>�-n�Q��C�J�T�BFʑ�&����7�f�k�h���|d�8���p������y�-��8*����J�0M�������{{�2�j��y�]������`Zw��Pb$�臁�>�"��h2���"�N���:�'fsxfT<�<�"[��#pc2�?��"MwKρ�n����rQntے7�Q�U1�k����Be1 ��߷�)�I�����n.����w�����
~��t�7���s8���d����!��d��3zyK;"�����=���׏�n��AI����*�Uj�]s��-��h���_-���Ǐ��2��[��t̻��ԏ����?~�lMP��rM`�+����*���~����X+�������l�����?'	�7��/���qܡh��D�6��|�}�x�z�JΚ��h������z�({��5Ţ�v�K��4+�(��5Z��a������j�X'����6+X*��d��e�n��fn�M�֎�`ʜ���#��Hp�ջl�6��d�N=�*P�qU�HB�:[rFIY�ZX����h|h�'�֯4<[�:;`���~k��"C�(�d*�]L���>*�R�c�~�e\�V��
u���6�a܆��.��J�f���n���	���?	��H�L-,� Ai�����{�_@����ݐ�l�S���I0�@36Z���n�Xwe��@��U�!q���������k�9zB��Ԟrtt��X�	����~��g��Y���C��5����2�0Ò�#[q
gЮ������G�|V3)��3�t�Ф�O �s�r�1�ABr/�P�g��n�gw����j�J{ǫF���A8l�J��Y�B�"ꃃ�H�_�kDΪM8g�X���h��E�~�p�fP��U@n�4C[�9�:���<m�Ǉg���X��F�[p�">*����k��V���Z��P����<�ڠ���c�Z�)���j$�Fy���x����%��ʳI޽�".ٌ��d�����%��4KM�$��Z�wB
�-�P��]�־e��m�f{dr��
 &��j8U@z`��'�9cA��R��Z�r�F$r�i�e�mU,��{c`�>�Ü��C����-�aX�[��g4�d})<�����"�k���D��������W�F�d�������J��C��@Z7O6���MUY@�� D�2T��tg/#¥X��6>��x�X��b���`a�G&]a_��*ј���A���;�ZP.P�6�b��%�i�y�y~�tUABN��H��j�x�
(O�P{�7�-={�߉���<.%���
7�\�}�VA�ʞ��Z���es��d1�Q5.>;:������s���W	�畻����_>6#�6��]'�3z�<���+�VÙV]x��q�qǖ�����b�|����u�fT�������~0�� �OⅭV�л@FYh��@��%u���^�20�h�K���+J[����(<Ѡ��qn�Q��p�{Q���'�܀�i��5v�3�)�$�-����s�IO��������Y�b�0�z���+���R��n
�ca,=�W���gy0ɲ~��J���U��U��L^��$�?Zz��U'~k	r�E*D�xN�����e��J]��Qi�@�~f���~+�X;[*B6*�FOב��fwP�t1+Á�$�	�\束��,�8n�sD�k�Q7B���r����*��^�&�S3,����9
�{ى�oDF:?^TY�T��һ����w�,�q�DF�ڛ�����v0bl:Ѭl[`���cU~��rL֠_@R�s����6Pi2>����2�Ilo{#(�`*�:nE����L~J�����^��ө�_J���	�h�6S �;���X�uT�W16��Ƨ[Ęg�l �����E�Ӿ��5J
�̯̦� .pK&H�hG3+�7x�g�d�R_uD+�`�UJ�l9z��(F������E�a������9��[�Hxp3��9ʨn x�	���'û�&�������.hQ;Ð�ҟ��r�LnGr$$I���1�Z}9��n�(8��T�W#|%µ�䗢�
A���m��Ѯ0�#S_C�ն�u������ΰ���������̯�v8�w	�T���e@�!�8G�	=��e��0||��\���N�g�A0$�[�7e��&����=~���chhͯj�ƽGhA�����XK��NW}�)2�R.�Slp�|�GghղeIN��:�\/�LG�X�ŭ\d��.�~��?���,��ֵlX0ğyb`edo�i�
n7���Y���LS�a��U����cA��Þ���/v��}'/�T���Ê��=#�%���g�6��o��3�pN<i�(V��I��P1��0�&��׫��,�=o��~L�cx.yV�)]�&��
��<S9����q\�� ��[�?�F���4�?���]�H�5��4��6(�M6,��Q�1�Q�}������|�fZiN��/wN�
v�U낃L5���v��W���!�x����2�wd��i7�Y�|�uˬYL�i#SE30�5�$Xv��c��9
�'>�wm^H"	��0:�̿�6��F�¥�Ǟ�9�Ԥ�[�8�ϗ,{�y�z�Ź��\W5����z9��-����D��|�D���~&K��t��);"��蕵���[�T�-2�6�EE��)h��X \e�k���ɿ�d��`�-�k�(	YE+q׳�C�`$UW\�oV��$F����;��V����NP (��#%��Z�&� y�o(ڝ�:���{G�� b��cr���p.�&����$���t!\>_@j�ʾ�`,����g��ۻ�� �[eP����VJ�UA|�%���;]-�Q�n�d�p�%Es����fc�쮳�U��:q&vI�z��%�ɂ\�-B��cKʏt�g�#��'A��Q�TXﺐ(��j(��kq���8ʿg��y�*9l0.�9��^r;�����J��
����@r�ɥ�tbJYcc%�d�A����c�Lq�ld��Zh�!�IJ#&f�Z�r�&���ĚGWʢ� �1Sޢ�;U�5�3�K4�b�����d����p�S{��oC:`�䘪sq<���F��6���Ik���Q:
��S��pt����Yz������QT��.+����֞�a�L.8d󏩲��N���M�q.����J��$
q��W��æ��o�* /���[������c~�.3B�+}�Y����PE�JД�o�5=�X�жƠ�8���H!�Na֏_���¿��:���>:����+Hkj}��.Ұh}:�����h���{�OR�]��l������ˁ3�j=y( �N ����o{�K��feb�J㡯I���N��!�\*�߯W^a����ӝ�XM�Ģ�e��s�}�v�{�L`��$W8��H�}�C�W>W
��it��2"$�^1��L}�m�<�[��t�w
,��ǰ�����muR�5א6�g�Ѡ�^#9D�p�Z]߷�W<�[ռ�)h��`���U����=w�ύY����K�	��|9Y5�Z9�5-�c�_���D:��� �G���@�]#��'{w� �f���)��h�U	U���oVi�0g���Ab�ˮ%�8'f7�Ă�!>����֭���y�z�rzEm�;�p/��������v���l�4sy2�?�u�(��<z��@�`)��!��N����0wG8�-��?}�/{����%� �ls���:��,U�:�	�Ll�B9�OX� l<mk���5�[g�z?:�i͆�N=�מ�p򐿲(���y�['���*O�|�AT��p~��B��%c��:M�|�3���. �l�î��MgD������3 �
�����ͭs���3L�QGO�n��ס�5|%��+)�]�*�PA��p�"�"%�IU��}�*L�G�1\7�����3V��o���%���*`�V�äv�R�~؍�T������MW��U�!�ƽPb��s�"fݚVW-�'k�-{�O`;�!RjL���O��:��)6Tz�4��9J]1Ѣ=2hL\+k��{��ÿ�����g��&xk��Rʢ��t�����!�q�>���Z1�u�ZO�`mE[��](���9&�:OX$�!�%-<^�=��{�̏��=��yc��Yp��i��T�(o�Ա!Ά~����4���ɏ��y=:��K�WX��aп� $�G�IR��$e�?�(I�(2t�� ��ƃ{�f+�#�mB_0�_� ��Lm�,�a:iO�ŶR����L|\p$���(l&</�<���B1��T��?��Z���q�np�k3ώ$j	�6aZ���)-b�ز7dCc	rU�/�ӥ��,._�J�vѴ
�c�Q?�����顂���J����_�Er�P���O4��u�{Cjb"�Z������⤯�ⶂjH}���@���V̤R��p�a�zX��5�鮾�gd��E�*����Hr�I�q|%�|���C���+�����̢-�QAy=kb1�qX�'Z�H����Ր����@R.�Z�$���y���	�=�n�Ӱ�n7�xե�!ͪĶ���l�E��*�sr�D�-�k�4U ��>u�]����wq(OF��&0���3�R��8����7��q���_׬�-L�&m,.��n{�T�'%�3���w�Ș���橈d��P��(e�ꑁ5:V�đj71��NW�#%m6��GϿ���mb}���e1�6�U�
!�����%e��.W0���^u
?5�V�P��'�]]�,_�Aj��+VJQ-�����l;�<�BEސJ��kۇ ,T`��'�Ke(��V ����dH>���_�Ȟ���	2�EsP�yr��T^��!�	\\�w��3�cXI{���nV�K%#)Z���������[��;-���|�:/�F����N� nJ_�F�Ɗ���S�졭*�
8�U��8�����r��w8�M�L�s%���A̫�{H��@�`��C?��4�O3�Mt`<?��Ʃ�(���\�T�R�:�d�� "�T֙h�53�����=�������*�yfz�4�A��ꮑIpfF;���J�ª�T�t���ԥ�FQ\1�yA<�+0���0�a��T�,�0��|i�	��}
cklA�a���&Gc�&��ZRTexel�A,ˋ���+��'�h���3��N�r��)�L��(5%���E�>�L�Zb��!S��e�B~�r^�i�#�V��<D��}��~�x��7�6�(���LP���nm��F�|���#��_�CKFę�f4���#O�t]�O4�H�;�isX���@��,���-u
�O\����ztN�͢�a�c{�|O��"\�K�Q��lU�����%de<xfu����b�X5p�'�\��(���,a�30��-�I�d���W��wm���{�XX3�$��YtH*$���Uw�tR%�g2k6`�~�䩅eQ//>�6��L����q*��%�-��џ�X�D���U�-sfp�-]�K<�L�5����G�^L�FB��l�&�Пj�D{�ˎ#e�������J&u^R1ҞM(�R�Q�Z 3YR��2�Z1�0?�|��|k��6X���σ^���i4ٵ��j�8�A6~�ʶI�_�7:�C��`䦛�q��w�B�[���"��9���S���%f�@�W���J�Z�9)�e�:Bh9?Y<�J)�oSV6�¹'cuZ���^����m ��P>�����Ӑ]�@������ <���Gb����m�rb})\�������8�,!�'ap���p�Mʁ(��cs�T�8T�6��o�ʱb���x����Y`��8��dQI�R}1��~��)'ƞ u٢����'	kґ.! ������ 3��$[,�@Cq�7s�'�a�=�v6������:(L5���`K�
��B���=��}���~���#{
�\�£4� �$���I�]C�5_�7�O�%�S,���?�e)�,��Ē®�ڷ�a���$/��Ǿ���ͱ����R��`�����0k��z�?'y��ri���`ҩ��]B9Z��$�p/�z���˓f�dd�q�ۀPo$B �s�p��h���	4��d��\s�)��&XS��d��U�������yh���"�R��b���+�c�g�?��W+d�R��Ř+X���;4[*6�� �����?�mt\�-P�һ��������J�[4��$�c�	���[)�����P�o�l�D����[ȷ�S�V�C#��
����=VGl������}G�Uoc�Ub�����Z�K��p �ue7Kg��{o�%���X��;7D�"�����,���̄�!Z��og&�o ?��
qՇ�����<V��_�e�Լ�-G/:�X������{D�=��ݗH�l�v��I=�,h<zit�������^�P�&���P�\$"u�Ydd|\5��b5^��d�dH�����f��C�[��5�yqm�����p��j㶗�uH*�Z:]Q�[mfP�f�kEQ=�R�h�="S�K���eK�����S��"��&���2:*{��Ø������g\�?U,U'�����se���J��F(Q��;�����?�Mw�J�1r����};7��_�d�l� ��<!��w���Uz�4���Z�2@�=��4{�C���x�WLD��G�6,�lO��`����t[pJ�R�{=Gл�qvb&��Uk�wi��V��igH6���x�)��P~ �>�:�F���8��Y���Z6p��-�9��C��qS��V���;
�'[���8��L�
@�/�����M������I)�Dp~�z@��D炷����S���h�Bl�|���0�ϵfsf�/} p�]�VW|=Ⱥ�������_�u�K��oUua��g��-����PrWH����s/��ě���l��[\��3)7A��TqE4����8��x`�²�V\g͸�g�3	�^ߥ��y���Q����v��p�y�uo�EG�h�-�U,�CjyY=�����l�ɐ�9`sw��Y�a�>�Y�Q���CR�l�o�"
*���握�����PZ2�E��0�~��m��ϰY��J#��Pϥ��]8J����"W�#k�Cݐ�6��-e%q��$�C��舛n����1fڌ�m��{��$��y���x��kD�F>���]��&����a���>ްp�9#��}�zs�4��̌-��ST��0V
j�#lۚ��Gw��q����YI��ا̸ɵ�+:k�|;�o�z2�����*��Uzi�\�Oh������O7�6%�~�#0Y��d���Ҙ��4�)՝.�G<�&���b����̰��&�����X��F7�K�o��ӧTąM���g�װ)�k!8s����0�=Zӣ�G���e��}��5�_"i�0�t�tDD>S�k������~�V�l(ob�ۛ&��)u�%q� !ʆ#U$�ue��ؓN䦾����цQ]E�K�:Uy����v�� ���%R�����&�� n�?�e����!�>���K"r�"��P)����&A��^/ݼ��г� ˤy�s�Q�)v0�Ɋ�,�GW�NN���y�K������BaV�sg��8,�R�{_H*q��o�3,���)Z�!4��|U�ݔ,wh!��/��[����[��,���!7�PA��~�NaTD�*�g3��%!	�TF'5+U��B�t����88��_j��n"��2��{��% �����/���Z}�{˻����V����ۋ�d�_�������n�Հ6��u-�3��	kV��;�j��0d�!R|���;͏Oϝ�b'���^�Ea��� |�X�v��Bc�=8�- *�9�?-�H�D3��)���<��6�ȥ����l�.�g��,w�=>_�ޭ���٬ӟ[�8WoE8X&?�0,���F-n�Y�?u��U�1�f�)���گ?��m�7��m9��ȗ'�%�Ǟ���s�(����d���s���ڲ�=�W}��n�_Y#:�.��9�P��8��u���J��#���%vEL
9 
����������6(�xg*4m�|�dz�Z���~�Z���F�RTKb����� "濇�z6/�J�!Y��%ӄϨ�XdC������I�R\�>��a�>78#�,�7�%
;��d�Xk4����dij�
���V����wL���+��,$RY�D�I&
���K"�(Ϲ�N���(��L����7��W����"�nE�o�6���]�{u�M6(,�/qoGʻ�gX�r�T�ЋϘv�¶�L��!�}�85@�;�>��RZ�������+���e�����M��K���PN�/�i^_��|>;���s��J�c��% ~n`B�ےM*_d��F��Ɗ^XF��t($��1��Q��~g9ʼ�&\��m���_MX���<�H�����_$�����yǐ�
�S���_������>áI�y�M��F6=��өu��>^�=9A����?m�Q,8�b�=8fz�>�~��P%a�6�X��-�r�Tc��F�9������	J4���I�,Ӻ3�I`�HC�����&��<sɗ���U�����Ha��t��f�t~��d�Y����4P��x��oz];+�q��BC�AP�3��p���C��fZz#�"�a�@�24$��}��.�`����i�,M�������Ĩ2c���9�ȗ��6�D	9Gf�*}�Mў�?��]��0q���ev���b����s�b��0���p�er���Of��)�P���QtOױHq�V�H֪ͮv�|����G�"$�l5�-/�-���&x?��^f&�{O8���*��m���ܮG5g�G�J���h��4�=j��|z��3����Ol[�A��։��(3��M,0�o.7[�g;_ܓ3|�����Ε�XTu�!xӖ��+,W�]g���4�:�Ů�_��O	;�F�Ч�O�״|��;.hh�V[!���9
"�D$N?x�+f�5~�~BP����\	��c)Z�l�MvNq���SE	���g�Q��%���U������X�"D9H)��m�%����������v,w�!|���T�J��<�f��.ތ��@`�qBrp]�T��&��41��U �O#_+����dOB�&��j�s[`��^��~	W����.���zWc�q��D��,7扷ڃ�O��i}������gbͼ]��9�p��o�U�E?���	{I��z(_�]�k���^��_��"�L�L`���ۻ�˺�����0����QD���FBU�+T�w��9����!y�G����0)���M�
ٙ�~N#�ۈ���va(�|�@���~���U�j�,Sc���ظ_�Z��Po�n�9��3���0�?��y�t���c�Q�i�chO(����d�t61>d���rc�-t����<$h��d/��j�����Ԟ�Q�G*���O .�%9_��nT�f)�`,�����r�#iț�n�j��ɟ��`Q�V��o��g������;_K"ٖ�YW��Y�J��ޮ�6�I �������!���lO�F�)e�|��k}�E<�GLq�1X˭Duy��G���[+�o��*�}�\2W��<� ����G)+\�}��^�����Q���';���wE�xD�ݘ��&<"Ҫ^�%mV&82P��L^�q�f��a�qz�Y@4��U^1���-�Eʌs6�kF�2�í��[�yok�R�k�׆��?������E)KVt�|l�rF�>���M�y���O��*�2z���d�s���
2�ݤ�Ć��5.�����e����L��ɔ�S�.̟��I|���lӹ��?D|�Nq?<+��iH#�f�'��c�Os�O�o��֓������?="�SK�X佁�;X�uζ�wd]�*���g�o-��֮}�<�}(:�Z�)Ƀ{�'��hWK�5E�g\�l0���遤�3o3 P`��촍,;��oD�����R��j4���E�$Ď��qB��S�1��.�ѯ1qTי�����Jf7�]��պ��c!C��(��߭��\� �.��!�����ؔ����;[�@�Z�����!D��"Jo�z�vwP�?#��mJ
�|�?s��%��_�Y�L�5��缏�ϧۈb-�}���c���Y��#��(�<�_���Au����K�.C��r ��[Qy���=G7�æ�օ\��V�1?s�mT7N�E0J�Q+z� >�o����×�hmZ�\R�0Z���&Хڑ���[bJ�u�v�5:,���!�A-,C����q���I���P�6��̺��d�2D�-.�F<���ˠj<���;�����E�5�E������b��C,���n�vu\f���E�q���l��ȧ:���r^(��*�딒���Ȼ���!!��=������v��yA�Ka�ǋ�5�#P��[ �u��.{4I�����'m`$��k����~)���F��X\[P���rm��N��ǞŅY��� pHō;#*_�]��X�pJ�b8�Qc�DtL]fy��;�E�b�ݏ/��o��Ce�C��|�7-��my�?5Mz�-#pd$��h^F���my���l3ր>VI36)wۛwc�X���.݆ FL�F���F�u]Y=��sx�~R|�J��1'�z�`�ӽJj�k]�)��
�q2�w%��oa�����Jt�{dIQ�������y�<W�)���~�o��C�jY�L���e���6R$���M0���� ��T��S�Ih���ǒ���0H�qe񐘜yW��_�z��� �����j�|J��wXf^N�Nn�o�#�3j���I(�^b��P�)f�أ ЛkwD@މzP:�$^,c��5o���e���ny��Ē׻�y��=&�]�<��?�=�bF.�@Pq �7�C�¼����r�Z�.�N�>L�r��SOL�}k��\����׷�BjB].		�\�ꯌQBV����>S�C˂k��:M�:�v�@�Gm���mS�+i���L�w+}$/-�/���
�3�������_V$�0�:I��R��[����5U*����A
יu}�y�B�}���\�n\��S�gy�A�
�Ff��^�LJ�	D;�n ���{���h��!�3گ�l����]u����p��..�Ǽ��h�I�d�z Udw��*������U�z6�hQ���+Լ��!/w*yq���O�37.�Zj�]�1�"��<�IVӻ'������}.�%�J�p'���DM��q�G���L�wK|��'��)�'gB�[a>Kɾ%C�|��#Nkw�}��k�.kX����A�����*���j�OW��_S��Dϗ�z��G̑�=$E�򍛚X���5��a2�O�/�m���K��U�����	��
�ƥnp*y�1-l���q�c���Z�\~?�ke}W�;����y0��0�"��k�_�A�@Q�/#�p��p����9��7���[ǲFUȧ\{J��^'�i�4k���]����/L��#�e�0fi��y��Q��"W`��ɸ/��
�5Sg��6j6���l\":����cԤ��̍�yXC�5D%wu��8�Z���:��1[+ą-�L,.�ޘ��9~P%a�v�Z��-o�j
.,����k�F���K�Ee����%[bT�z~����mz�<���x�Y�ꤐl(�9�؞��;�йg��RL�9
Z�&	�������.$F�m�������%��9�MTJjE��]�6�_�����y`*�LP�����߿�H�ݑ���b
���|�aT%��B�Ap̽/���3��K��G��.�� -rӍ��!�Y�����I��c �p�}Ռz�W����`������k�����rZo�G�$ �F�b4N�k�Yr�U�D���L��ce��|,�a;U��˚���z1�jVi�GʎA��@�t��4�Żtw^1��0H~��-Z�*9[:U+��4K��r>]q����=1��L�z�L�]��������/�ǥ$��/�������7�$�>ILaǕ��B�	E�O;b��p���Ȧ���L0�ņ6E������y����'R�Tv.�/<�ƄO�ʁ�#H%i.F]��	1����7��[ ��?��׊�~��������d��!bi�Zʔ'S�
 nǑ�?L�,#S�[+�!(��kŠ��Na��ѯ��\FJ/�������E��KrSP5�ܭ\WD���l$:���kns[@ݤ��������ɟ^v�\��Mƭ�fN)�~�l{Y�?M��❳�6q�KEVח�VQH#ӳ 𳩻&_-������hSv�����Wc{��,�A}Z��0���Ң����B>'�á��L��ǀk��+z�3p�[����ǎ��r?JO*�S�5�N��ּ��p=M�e����=�r3�E���Oˊ e+Z_��ц���?k�^�H,���ƝTW�3����J:S���Jʸ��s�\�GG����T������k)�JW�t��v�����|��eU^;�ԛ�l��|�r�z��͘�����K�$�ë��\�۝É2�/$���}�\?�z��
��d{���0��1�� 	o�B_��#��Jp���b��K؊��Pj��َ����rKQ0�-��7�,?ro9RT�)��膯��Μ�lI�c^:q�V�PK��=�"I0�9��6{ui����hX{Ɂ���������vC��CR����/2l%~ǽ^0 �>R%�>����C��pp�ʝ�\ѱ�	�{�L�]�޺��N���w��*#� `amj��9��ݤ�&�����Fy��L�Q>�m��In�C^��,��!���p�̝�B�r>�OD�5��%�� ���"�	{����b��s4s�v�e�郤���ǰ�/=����^���}B4���bb˚�QRāM1��z�q�V0'A�G���E䈨�[j	~�] ��3��>*+g��[U�h�<�x�����J2dғ���l1�X�q?l�8a�U��2MV��k�?y{n<�@����Lw�D4����,9%�Y$�P�.C7Q=�"3�6cH�ω\Ѣ;ݒ�&��cU�\��\����S�ξ8%Ip%7�G��^("BA�I�N_��n��$J�s0��f̐i2���U�W����"#���&��Q����ꑢ��W����O��k�(-��ӎJ"Rۯ�
X�y����^�,�F8c�.� )ʣ��I��wX�طΘ��mD&�rmP��iߘ)�Ks�΀�y��yÖ�P�i�p�
�����4��;��[~=.3�ic��Z���K��$.�U��L5b��G�bB����X�Z8p�ڛVC�[%B���^:L��|Uժ�VNx~�d2?�������w"�ED��a}&K>�pa��J��ɇhw6�'"��:���Z��(����s�k��q�jlE�������xZ$� ��|勇�;�C� s_��(�:�n,J ��A.
{���	�~^ט1# �0\��B�?�B������]1]�뮖>������y���P,����⍽V���E$'ovl`H��Khd���=p���"ӫ����᳔4��j2���	�5b�0SR��4�����ɁDq����n�2�����^�Ϳ$�j��,�("
��c��Bq���;���G���"VfI�o'	U���}p��ݡ�	^4(jy�O�J�?�odR������������ࣗ���Pe��mQ�*I����ci)7v	q`^/|�7�3�s�I�@	]:S���\�h���t3��'́���g�`]uDG[�)���q-6� K��W��6�t��2�-� { )��מE�;���9~2�L�r���wt��,���mj�л��U��[��d�W����!�0���TL��y-F�O�r��G����/��M�aޱ�3�,T��W��
����,��JS�X����͌��Zc%/�0i][��d?h��_�r� �q 3@Bi�v�b��O�m�8�.pM�{h�f%3<_}�0��1�j���#d�+/,��`�"-�S�	�!� �qN��u\�̅����yh��ľpkl����{5�\���d�4ґæ��.����O1½7�@'z�!�5����e�)���(���j����&/�M<:z�-Y1�?��(S��}K�L�qC�mΏPvI��aE/�2��bV��P��?k�BE�w���7T�(pK�p�=��Y����y##0bM��]��?�v[�Ć�̳���a�����x��r���l�#���]���ǆU�"�d��I��7��<��{�����N�q������A�9�5����%�A�H/��I�D�%�0��H�'�8�Tuύ��X�MD��������O-��V%����#��1�U|
f7ۀb�#���SƸ�������4rM_�s/)�-!� =I���M,3����x�n�����g �������&�ŶX�;�����t/O�)yl��a�0�oh촦J����o�Q9�A�"^r�5�?�@����䁭�}��r4L<m=����)�O�  mp�����}��9�olz%i�*��s�o����5v ��'�:�4�XO��
$�*�Ew�M*Z������B��m�Q�_�}��e_:0�{p��������c��3��$B禘�����O��ʥ�yK�%Jb�"d2��Ҳ��f��
��DF",I��S�ˢ>�\4��h�A� w��S���c���@d4=�_�~k�ϰ��V�u���f������H?Ρ���"FI��>Ȃ����_?-r���%�F���?d���-u�P�ݨ7�8@T���&��-�pX�r�A�+�XC��XꍏT�.�@d��]�}L���.����/���y��!���'_�QQE�@TNy��?��bi����U�;��	����^�KӅ�IZƢ��B� ���*��M�R����1����B��:���2�3cC��%WE�����$HU�l�'�[�ރ�`\�GG��>��F�Q?'M>�~�E��fn�Z ���
y3&a˳�ᓧ�����4$W5nʑS�}�V ��N��[#� 
��h;w��'>!�c_nw/���L."��6V�1��Ov�x��Ğ@t#i�͇7C2���Q��[a���]Z����J�K1�����$@o�i'�?�o�[���D1�v����}�D�J���d�z3�TH��$��u�}����;��=��D׈t�k��lm��	?`j�Lt����7,AFO;� �¬#��j�H;4	|3�o	SE��oY�� ��kL֢��\�_�Z*��X��5bV�B�}+f8f�}#���o=�)ۆ7{���jK4}��4�g+�޳*�\�h����xK�N���N�s�R5�L��)ZC�f���(�9p��z�ir����+O�52�O�]PHQ�_��,gQ��x�@�4�XCy��}��ߝBث>H���Ϻԉ���J�-[b�:,fx�s�Z�'��\�x�4��_��ݐ�|��,q6�����:5�+/��9�Qe��#�TAi��'
]�ɸ��ii<�yu�����Y9�/
Mm��f����P����X��ƽ(/q��>C�:���Q��A�j�ܘ�wWg+{� ���i#4�p��l0��u��K�z�O��KYgEE�w�>�ˎcUxn���a�C�`BGټ�5$��|i[��\�oӓj���q��7�h��z�I���I�y;���Me�I-������6	h,��H��I�j���&��&ZU���f��[¡XHXL�*gczI՟K�(.�HU�?T6�sgo��M���)E��n��}`s����.���)ҟ�l�`�Yt��2|F�1�m+Ą�"�$ı�m*�� ��6P������#E
,8�M]�(Hh�3H�5��W�,��[d�E��g��JG���.�t͑����;���,���`p4G��1R>
\��4Z
!}��}o�>��^8��J8�kޤ�dm�d��קA^�n�x���qe5؆�ECoyf\)�a�1�����8�@Au(��1.�(�Ձ�h
�~m�h~MRXBX��\�_����^�e]Mm���Zo��i@�^C�����s��w��Q��(�_������[��8��+�b�	�s1���t�'�s��kWgaS�݀�.�C���1W��)[���-��f�6aa2��3��UG��T����& "/��
�7c��}�T �Z�5�K���V8+Q+��)/��E��=�2�"�"�<�Ģ���i������o�
ɇ�&�N��j�h��6'-ٟ����[&�������8`�#�a�����ܔ�&��<Q��)��PM�Iw�;O�&N;���	��4`�gEf|̃����|�z�̤k�m��s�gQt��0�Q�'R`�U���~�Cg�V
��˴%ą Ȟ�ݸ�أ2y	����$�1���Ʋ�ȇ�r����N7��(9�l��J��l�[xs°M;Q�a U�4f�O,�v�澈L}(rF�s�X����D�A�Ip0=���?�/��K`�e���b���Pf��z��<[�a�2|~��]�谐�_A��4g���7j�e1R|$Ņ���i�@֋�y�	��܄I�h��UO<q�wcj'�`�(d�����"���N��)埾G�ؕN���\�
L�8����Ȯў+E�=\{����<�W��-pVv��>&��w��D$U�bN�� �|?B���z�N�Q��:��CݘS��`�S,���w�!AsP�iZ�.<�ˌK$EmV��}*�.������Q�y�k�=�ܦj#E�W���h,�}�B(��q@�Hg��tyrѠO�@���x�M�+����\�M�����ԹQ��t�V��)��TL&L����g�]<� �ȓ]ڴB�(C�#4�`q�	>����3�rJ��Hi ЪDz�5DL���9em��3	�!;��T�,�K�>w����B�f��7`�]p3jK��{�L��
���Z���b-˦X:�/zMT$Q)K�����/�]{6iΈ�/�2��b����I�סN��7�4�?�� ����!qb�=:sd���ˢ���o�\���'�޺�d�e��B����a�����[	k��qp����s�W����tai%KX�F ���M��2�8�Z�PVA��S��������(�2Wׯ�Jr�AX�SB��/��Y6��2ȋ�L�ڵֵ��kŁQ5��m�����~l�p��V�|)nD��`'���|q��cH��լ��e&����\�����}��=]�\e|��=�&K/��)Eu���4�LN����� �|;�C7�J�qP�!������$U�pF�w2�A������N�����t��"2)�[c�����J�B�ƈs�
����ܯ��+\��qQ,6�͔�#�I����w��t)N�_C��{������z-0�(2�ɗ�A�+���
Z�L[��%�2���m��{����-i֞��*�<�u7c��ȟn��Ap�h3�鼉(�un����oe��G���v_$�d�9�6Z�
������B�jX�_�3�����e�'���^�O���&'�#��t�+�1"]�u�� ����oM��K�V�4�~=�|�P�GU+�@�S�6A�3�P7��t`��
i��
횹�M�`�9z@��U��F8@bS%�~ _�
&M} �$~�+�A��c-�qv�U=C���C��;)	�M���z�wX=��ӛ�Ɣ&�H�8�H��+A�r�+�<߿zV��b�$�~]G�7� `��8�Ф�k%sȱ|I��K�ʸ����^XtO�����	�~���l�v�Ϻ/P�[���.^caL��y.^�������a�S۵�����Fq���#i�!�f��s�cv9)d�7R�Y��]�엑�C#IqgnJJ��I���F�Lr��+�=���D��-��)�bM�'ֱ��8�ڇ�{���[L,6�_���A,���q(�n�d�B�Gم9f�\p*�]a����ٍen@�n�rx�JxT�$�8fj�\	���&�<`:=�'v�5��oJ���(b[�0�|��r'_� U>`�R�� z�H��������ԫD ��-��+/C�>�����@*	�lE�4$|��F�r3�Y�j��ʓ?�`f�W���'.%�#�1TO7��l��hhѵ�m0��/[��1<���
+پ�X�:�uϣ�{mC���iL���|2^7M2p۶U��*2�'�~��py,��"����^w��t
���]ǇU4c=�lL ��+�^��`�I����.�*iu��:�I	ޣ���\�A�3�V�)���kA�&r����}�.�eA�]��B��<'X�uEo�i����t:tʍ������!��q`ƿO��]�?��>�J��b��f�����HMV_H��2�2�X�AF�k�e|\�~�%�O�Ꟊ�WQ�{���K� \���RH���
z�d=����O�b D7w7�!�xVo�N�����Um&M���cj�vw��Lc�(m�"��E>C��A���tԧ�?�G�X���f�Y�c�O�GJEU��3�=f�R�up<��\ĺ7�GF�.�h�l}X3Q#��\IT]'̷��G�+��[-�*]?�E� <z�?鴪̌'��oK{��j>���@������K�2�O�����&�����_8[���M���NZ<�w��?�kD�W���H^���#U�ʹS�J��R9~��K��q�=09�g�|E���%# j`|-���"�1��d֌0��^*�>J�׶�yb����f����� wjb�������4��g�z#H��QqdR�L3j�đ��wu���:���d��_1�F*X�5Z�?\| \y�^EǯP`�_�U����L1�?�:�ѷ�I}~(=u^��?v���Y���lk�DQ=H����4�j����L=�%��6,�Ӯ�:O�Y�Iu�"����@����$�x�"x�;x����W,_Ჴ6Y+�tH�ht8{��XZ��v4�=���Ͷ�3]΃%�|�9��KɐpÍqn�doA��E�����=�)p���~�]?�s��b�*�+�'�2�OV �]����ОbJ4�'��d�7��D���9��?��A�#7@=����J�0����w�$G�c8�5K�ǫ�8=CZ?�s���u��V��>�=/��iY k�l{`�d�����	�� {+v�-c8ൣϩ �-jY+_D�����D�_�㩤�rZx��8j���_9���0.D,���s�jQ^fyE��!�-�8����|�1J;�U�u���餷��Mn���{\�ƨ ��g4�֊�k�l�1�U�;�aaH]��]�M���ݞ�
:���Fu1<�~x���������b��:Uธ��o���������v'�d��9Z ��R���N�_����U�xY������h�ܦIO��2�'i�Ei���`�21Nb_�?�Y��YX���+�VrG"@PV���Zm=�,��a�i�yAA�Z�j�#DCE�!���3ņ��^���G�Ijk����P���.J�i�;k+�k�&��]�C�E3Y�K�s^����r��n9�3��'� g^�o0�����������{%l����T������V�$��0�ӧ:X0�[Wi��H��<_Qk?{^<�!���)e�+�H�����?�ŝ�Y�F�����U$�3$���µ�NDx�#�*f�
�:4P�2Y��Y�d�}��z1-9��{喠1F�D��+0��[i��X"���i���$�q�\_4�U�;pt+aJ�1�1���
���,����>`��Shj��8�����$.�B��Io�2"�G�#�I1g������n��n�uP6pZ���9G�~ټ��K39~���f�4�Bp���܍8�<��dQ���B�#�X�*�zRD��pm Q��[ZX]}5�Am#�e���&��Od*b�n�K @��)4��J�)��yF%Q\S4R$��z���ƾ[Ք�Aa�IH5���޺G-�(��{����uv���BU�Vձ�+x44�jW4�@Q�E�i���w4@�k!c��;!8VX:H1�k���&0��[��E�!��M�hN0S��j��X�yu��S`�3oFd��3Q�c�/�
��.'�������"�����XFù��c�
2� +��[�����6=w~��6d��"�GTp Г��2����I����N{��w0,G�0���|4��L3:��ct�7�CQk�[o�D�� y��CY��vSV�	��i"�M���c����̨�&�LK:�#FZ��.{lQ�:�Մ��*NV��b�Ć�^8�_�wܵ�����4��*�#�\���ňR�d�k�����-�Ԣ�5se��ם7��<�`��Ϝ�,�i�~%��"�?{�����q��f}9��l\�=+��P�
�@���MwI�|���_y��̙��?[� �Rb��7V� ���D�R'v;^��]|�iT��'���W�q��*s��;