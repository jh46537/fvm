��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�-No�?�j:C�]�;���cu�����ҡS	2��)b�}D�f_�1/+B��א��e�(��	����6�s����<�(>���HE�:�o)���,�'��r�����CZ�PA_�=����>���s6������"*�6h�\��� ���P�r)���+2�q� j�})�X�X�h��|�G�M�G����&	��ͼ���o�)����mh�&m��y�`�}��نs�xm4��v=0��m��Ύ��Fr6�Ş�hp���B���:	���Ö��z��xtDn��h�$0�K5�������r�����Ҕ":d/PA���|t9�L&�hg�H!L����	V�OZ�1�/=��ƕ@F$�?Y�1�}�~Z��3�g3Ģ��a�J��j (d��&���Q�4�P~	��,������F��K�j�CD*�ע������f�����h>և�������n ��	�(�ځg�J��yx�)r�շ�'��z"����4��C47�%�&���0� ����M��B?�����d*�T,}����~�=)E���?�AJ��X���4w�F�nj?Ѓ���j���p�~>c���$n��nۧ��v���eFyM�d����d�<�e�gq�!F �cU�E�������Y}��*}�.�S�T��Ċ 
=�<r�"A�h�&�1��n���9�M.�j�����u2� �
�M��;�t��+<�Nɚ���J|�=�̗��k:8R�!��ɥ���{
f���g��a���B��$v{�[�$DQC���yh��!�ǣF�}�o�ǆ{]���x����;wtbދ��#�p$�O@�<��ޗ�r�	z{����P@b��س��ɻ0�~|��8��0�t���2�9,~�I��m��4���S6�r�,n��HԿ�<a��x!�o�Ű*���i��$EgsD����#@�Vq���w�J5��z��i2O?��6QD���uqH����>�Hd P��_U�P7ٕ��/��cz�L c�m��V��r�xV ��Oո��L��	���]��@%^�/)�?�4�HCأ�4Mѓ��$/j��P)��s�o��_ ��c��eֈ�x�cx$���)�)���\Ab-L\gB2@��W���1ɖ/�W��� �o|v�VJ:��z�0V�����J|%��Du�e��;�i�nB�������`����MP��Pj�f�h��Uƍ�d��8��G������nW�$#@_���C-��:<-v�Ѿ�5*�D�< ��Eh�y�2�K\���b�l��ܽ�ʓ�1�M<�c����𮻤C�
�<�7����0��G���U95d5����[A4�U��G�ěЋ�E^E��F�N���O��q�(� �c��WGV��ɖ���u���p�zj�ʨ�e�o���X�D���2���� 4"0<
�HU��W��'�wK~��ƭ�'�@*8��:��Ir��=��q�<���(ٿ��C_���h�u٭��s%���3��P�d�hcfФ�aڞF�4���!H Gv�l[8%��8��@��1���=X�^�`��鬪���Xē�K��	?�9U����Th�SK�)硾*�ӧ�_ӄ����;8���[�w,��p���[��n��I��>~VM���	�qL�b�-6
��U�|3Q{�`&\���g�d�*�Z�@k��[=��.��9W�\�Q5�w�(r�4,��1��(/Hb:-�8���{$j8w���p��ܑ뒴�=�?%r͒9Ʋ]�s��O�\Δ�X'ꁰ�?�=Q�<Lh*�vY����o^8ǜ�TU��������,�	*���E����vhvM:�l@G��ï4�{��P�`�����~"�
����m5W,��0��<g96�~!�D%�	ؾ�߇B�X�C�E�V������@�����2m�p���B"f���ב�sV�{M�v�T��']���$�2Bfy�}c6�0�z�/%��� �Y�&����(��'}�wE��kxښ�	��(���̡�F�w ��Ө�潀]Y�j��S���K
��$��G{,�4<J=;�����#,� ��(m�H��C��͹��_~>AX�>����L�)Q��E#�,����+��gi��^{4y�م &{N�>�έ�ν9
<�t�dkP1���H�g�CI���+?ys�]�i�]Mx����p+�ܬ�|��qu���%��圻�g��g�!���V��k�S���T�$�ό$�3�
�Q`��A]�N�	 ��rʧ����� JLEtB����r�|𾻇i�ZYM]xb����I��.�~�%��a�g?��jxM�w]�Aې�E�L�����hs��@�@�#���~͔p��}j0����n��?�#]
�~����t`����+Hs��l3��p�D�"fK�� �
+��w�䰫0h�mEՏo��Ē����EY����$M$v�.�6M{/Yv2�@��L��E{VH6�޺���Z���C4���j�Y;�gN4j��W�N,��֟|gJ�.ϛ�| Fo��e7�;G���9���IϹ�d��旴��"�8����Vo_� $�7.�-_��̷���O�6KQ_���PMem���V0�*��>���SQI�xC��h��#��z5s�&w��R&�%��^�B��4b���HF1a �M�7h|��_���)���2Q�C�E'0�*3�J�2�\�O���쩼m�7���t�<Ђ#���
�/