��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb��N�9��8�
`J�t�+K}=Y��-��.�1bSA/�\�1��Qr5>ڇ�֑����#J)�^���l�p�(�XiP�q��m*����,\�j�DYk��f�%oxy�ɘӈ/	���4`m����\���_b�s[�Ƌ-~�'���}��d~�� B@��谣������(�$ڵ���� �cZ������|�a<�#�IV��αF���b^�Ks`���S[���xt�vH|�X��Iv�i �G#B�ﷱRM���k�'S��Cw����Oi�z��*:hN�4�f��<���+AA1���´���9� �?^+T���k�Wk([�04�Lt�l�(����V��Y���'� "�I:��8���>���K��	�<���X݃RG��r��v���;�DO����m�u���l70dX�Oƅ�#Y�j��w���L+m�,�ZC`
�nx��I��Y�X ЌBW�J�K�I�I6P1�,�TT�� A>8Od.�@��m&p��u�eEU�;65,!��^6Q�9`��V����5���>tj.��wW�C�<��$?���+�����M���ng�	u��x^��#�3KBt#Y�� ح3q�0������8;��k�V_�f�z���E{"�]E�d�#�sHD��G�j�z2�x�#6ֵj�EN��~�ȯ�f��z�%��_��zL��One;}�<����Ya��c�-�����䘤"�h�?����x4�[���3�n8��t��K6&!x��p6��X��%��e���=�@ɐ� ����K���ָr�6XM��� C�X���o����"]	�s�RN����T!N﻿�K�S��FRՉ���B9���L�y���r��z��h� �K�|k��UTt�NI�1m�X�lF���0¿�kZ|/[DmZ�r9��y�=Ȯ�%I�T>+��FW�z�*w��Qi\��l{�l4B(��١��i���hU��劳K ��Lg�d�����8����8v��$\�%�35�� 1?�S�?G�&{�Ǵ���qI���B��M,�0
vA��dаaYe��$~9F�ރV���@�V(���9�E�t�)�7��K ����=�j�6(:�G�[f�{��<<��$������.!��m�� �> X���'�0yRI�J;kU�>$���X{�V�E(�}1��w����R"��jiQ�_�r�R��l�pۧ��Z�7�����ad�9��f|�n�r��*�.��j�4��@']�Ԗ�u(P���|,T�ơ��g�;a�fD��@dk7�Wv!������$�^QK]i�^4#C�O����]�V�bm\�q�qW�H�t7�{i���Ɓ="kJ��=�l2k��I/����Ln�*�MAH������<��$�y��+��"<^�$���W_ͽsP��@5�A~��#��q��tT�����4��ܤ -;	:z�"J^Oq��CO�4�(9pB�W���N7"@�n�n{Ż���ot��^a8R#���̾ȅ(�gR,Tt"Fj���[��7�_��QyR<醡��R$���i<��SE�Yۯw�B��L���y�fUݺC7���4�m��z)W��fؤ��xF��g�)�(S�b&����L':I]�l����� �*�PC�0d��<@��h��I�~�`���`��Em��D��7.no�`J�NDIx!�Tw�h^�س�2�z�L���7���W�!�#L١�e�b�@ߦ��[����P��ߙ��V�q�[�v�$�}�HJ�*�mL���7�M!bsA\cf[P����7�BTj���ʥ�6'I�QFv��"���Q))��O�|׸��7�#i8�)!�E�l\fl?��J]GlX�Pf�x�>���z��єd���
@Ն ���T���_/.�%����t�s��c$~�z.\�����ౢN���Q�҃&ڨD��ԩ={�]\*~/�&G~�#6�q.K�8V򽒓�}��Oa��pa.�����%\@�z�_[�#թQ󰖍>gW��������(�^��*I��6g�΀OA�O��.A|�As����+���}4;	9 I�-�@���'����%P	S��9��n��0��>�*r�ká���  �;�!�p�B��|������>�or��Ջ��TJ7�X���2)�k�Lܝ�����`m�)ݹ���d:�����	F�(��=�/��YR(�-*�t��>�m/���D�� ���q�DC��!����(ϕ�v��r|��+R2���D_K��>���������;��z���Ӭ��&记�㔊DM��O��U+S�"��/|O�vt����������N�l���\Z����x�Q���$�\E��%��}���KĒ�����<\t�yd)U�U�"���-JO���v��{�HPD��f/lf����1A��oX=��(�g���)��3�p|��|��r���1`�q��i�?e�#+�(yM�;�HbM:���1�'��u@�Δ��2��$ʓ�N|g:��i=��"���'����a��p�[�"Cʫ�
�I�+�>73M���FG����FJ���ur���������a}��H�h����?Lh���8W+\�;OZ����a4*!�ɘ�!�J�cm�B4�â:<�Z�!��?)�ʱ�64��.��i�/��~@�LZ��!���M��^�.���ݶ��>~S�f>a�aYq�8ٮY:㰑<qc'�+ٶ�->�a$j�K^CD�"��D�<2�E��|A�)������;ɟ���#<Q,�/?"{\ȍ�q8���$D� �O�N���������<�27yQ�����ތy�Q
����4�H�L5��섇,=��~ l�B�G"���~����-��ٜ�&ed�r]�:���c�-�4T��=j�<��-�Rn��O5kH�%b��J�/��bti촹�Xמ��$���X���w�k��}��g2tza�<M�)�H �I�k��y���k_﯒���{�)z�K��y'u/uK ����7�}Y�#�D�\�j�k�1��w��ଠ���V�����Yak�m�'���Y?.�HF<�r�A\��N��к�;���Sؔ|�A�}ug->J�4x��[c3�&tm��%
���Ȍ}�k��X��271��'�BPb=sX֙0�Z�`����a]%9z��=R��VȢ���,G�~N��Exw�S:�H(S�w���#��ѝG�apWJ�� Dh&��{(�-���f�^C�~�<!�a�,		�������� V��sS׉a|�:��L���~j���6�6L��ݲmg5q����fiy�ŕ��r���/����*ȵ9�q~B�2���|Fz��P$c b�R�Lͱ�.�U�ߚ�9��������>�`�`F���W���M����$8�%�5;c=+-��j��"�1�ր��~[?�0���)0��m_L1Z��@�!�f7�,
^�);�X�P��>٠��v*?[�km7N�d��I���e�.�nf�M���vL��4���kRC�.�5�ʪ�'�6�QxXG]VG^�:y�ц�� T��|x�r��wE��=]���p�۹���s�
S*�n
�5����6W7E�Q�n����b�y������^�]n^�Q/Sg/wOO���?7�S�U������]�'��׃�0�߿���꥿��|�(랭2Ck�ᙇ��U�e��#Ę8��T#H7��0��W9�/Eʷ{eF0��x��,����rP�-p'.�:�
Rk*	V���J�ͧWB�G�FG����NA��H��s�j(��PZ��DX�є	�e����w48��'�
�(�A����bM����v���Tn�D^|eZ����*�T�!`{�V��	~32���{�
�?� ֣D0\�R��i��)�6}�܂��vZc9#��Ǹ%�����&��v������.38)E��F�}m��څ%��ulSN�C|�i�g�)�i��.�]���{�_���l����pAi�nAd}e6^���L��e+�P�c`:����E��i������%�i�H�#&K�-İ9N�me[���g{��@h}Gg*QU|�߬�V� `&j�_��*?�C���?x�ŗc!_5r�K���X�P�8�}K[=����Y{�K�?���Xм �m0u�ʦ	%��O�SB/�qTR��~}%�S���(X8��~DVF�#�58J"?Nң�Ob��О���QF["A��e#9�����&.�"��2���҇��r�b���~L!��2Ը�W(:�<W�)��4�+h����,I�� Awu�v	Q�ŝ��'f�n�j�,ј����b�^�oT�*��N<��.������T��ⓢ���j���D�uVU-;)L'/�$k.��K���u��^L�2%�w�ց[<��F �D����Yջȧw#&�,�^�((iF���W�R��W!P����U�ؙ&��tt|QQ�J1��`�k��4�N���+��e����+�L�Z�Rj�K��O����Wt��Rي���/�.H�䚑��H5����Aծ��9�}�H)�ؘ]5D�C{:����񰳓��?��z�9p�y_�e_����Yq�{��H�yHj�{��|����|㉠�e_�>>��y$eoÀ6ԩj&!�'������!2p���X^z�� �$N\��	����j!��!C�:�.�.�>(Qֶ��j!2��������VD�*��.8�oz.oƊ��O�r�r-���w�Ѐ�{��2&쪋����g��SJ[X`������ԚRc�TmN�&���ܲ�,\��K%�ux�n�+>vd��K>�ц����!��������@!?%k��'���0�ё�� G�Bi��G.Ê�9RAP�bN;>�q�P��=�k ]y��ǋ��~j*���
Z�*J�ł�Ţ�1i2��T��fp�}�;s�W��(�'}�m:kF���>`Ĳ�`����=Z��c���X�o9�)h��T�+�����[C��2��gE�	`�M̀��$��4��<T�G!��&,�R��p�/M;3�/��t���ks�C*�g��I쑞<���g�:��۩�*X���j�Ra�'=\�(ڂy/�Qd�"|^8��y*R�18�IJZ}�T�k�H魏\�3lHҒ������K*ؤ!�5���U������G�l��Gi#�%�:��Juv� �I/`"{�_b�^��RFM~!���=�x��d����Z�p���nW?����f�/5�P��@ h���4����_Ăڢٍ�Wbó�0u�=�d�gx1����o��B�3mZ��9���a��e�����P��s�i�4)ބ��k�큄��{W�{����n�����|�+�|��m;��#�|m�َC��<��B$K���`d��ͧ��y��������_�n��jR%�+�7��%�剷�f���c:�o���[�M{��Z9x$s[�{�#4<����M|�Ò�^���y
��1z�0�bP��/j�VI]��?��;m�P���$aP*N�laj�E��*��?�z�_��8�����q���=
5 ��܂�O�M'��{��xr/���$De���ʯ�mAԱ3�4'�M ��'��j̆�$����` N��Pn��1�͌P�-~�����\4�H�,!� �z`\S���_4�)�!�ɚ�x�F�J�wC�3����N��&�S+��=죴�rA*z��d�X"Ci��7���f7����\S��M��>U�d���~�,)�a�+Ύ"�V�>PӐ��� 3��d�! �������-�! {�l�I�$�!e�?�����_��뷨�A6��V�����4��L㼫9�E� �����Z��� �Wx�}���/.�a���7;U�n2��p4c;�0N/��;�7���ʕ\Dz�D����������G�7���i�����8���̍����a:���E5H @-S1J>���=V7?���0?��͢�"�Ì�I�h>^xΡ��K��$=�9������V~�6���V�"#V�j�<*>m%��<�
� ta���� ����Y)�i���H�Z��w:W����V�����N�Pv0��&����\����Ҧ��N��M�N��i�?օ$D�駘�i[�~yO�b���,���c�C�oI�0A\������H���.��o����[�]�������ͽO���֦+ErqY�e��m�7�ɭ���Xp��U�J%e��խ*�E�{��y��p�@����)Ua��s�P`6��)�v�(C=�����V�gM��Rb�Rs�NZl堙��B�X�G���[S߸یd4���g�� 7i3�CS�I"�����������7�n�q,$ts��!�s�З�L�ry)yР���J.GќN�:/�C�u�e�W!��	BPlC>i�i��M�x��A	��A�G�M�5��B~���|q9e(b���e�+��e�쵝q|��9#����MP�pV`λ(��ML����E6�RՐ��F����T���LQ��q�"V����	��es��W�ΨB1�AVԊ���I4��Y�Jx�:�M"�/}wX0p&K�YH�5
��ԸI�~?����#>�g�)�}�o��d_�H������a���X�v_<w_�~aJ� A�(�(�����v �
����Ӈ �	�D�V�Ztf��q�Z'�"q�Q�X4�&ܣQ��Ăm|A"C�Nr(�l蘒	m=�������U�����#F�6��n������������ŋ���lfe�X�m�M�w`$�"�L|���([��G�fQ�ջR�	odc$���`RK`�V��?hs#Ow���ǘ�������V%��	�T�~�7'Ғ-��0�I�ԗ ��Y���:?�����[;�V���G�v�]�(���R���h�n��Z�R�S��o�]|��\p��^�I��Y��`�2ɉ;p�{(�]�$��-�_�8R��Au�?�ͫ@�oI3��>��PL3q�4i��>>*�=�`_ �-�Z߀��ɰ���j�b���N7з]�*��*����6)C)ID:�hzѲ'��;�	����R�E㮊��#�7��������X-�'�~��+�#����-4��ߜN��4U�퍼�ӽT\��]s@�&i�um?���rU���.һْ!xm-qM�W,���^r7͖�}O�kH��
���3�ϔ�P�����1�-�4�HA2�/)2ﵦ�P�TQ�UD���`���Ku��o 8㤅��9F��~Sw7��*��n��~ߖ��De�n;霥;��]�杲F�̔�lO<��E��>ӘDĮ�;�Px��qK*�<��ċ�p����d�t�{�|W�������)�7y�*�@ҙ�}H�M*���3jx�6x�~�3C]ۆ���b��@��==e��8���q�͛�0_/M�`�q�J�¢����.�A����	�ѓ���/�2���a��D(^�
�B�� ��<���9q]� �	!@���y������=rS{���B�N����5��A��3g����#8�1���	G�8_��jXi�c��\G���H�*���?5}��R�j?�������~KD��$��~�1�+A�d��h&̱��l���D��(��������~F�e-)`�T�|Pjab���fvu���_��<9�v�T�~��K*yZh��g�:G��������G���hw���ϙ�3�f�E���d��+�(�@4*�5�����¬�7��lD�֑8�[�"��q�Q������)�hھ�"���݈�嚧��2���ݗ3J9�e['���+b���O�Y�D$K�'�6'��
%�%}'p!����OsÍ6�g���Nk��C=�X�_;��d}i�^�6�9l�� ~l+�ӫdI�����t��*p#o9c� ����΃,
�e���3Ÿ7��!ڰQw?�TH�X��%���T>�d�'�z*�>INS��u%K�ֺ��c=��p��H��G̼����^>\�����ϡr��Uހ���LH�y��FK1���F�(�«Ix��]��MF"�����mw��n��1�K�	�!�5>�tG����#��E�4}������z�[��4k�*>�K����S^��q#O� ��6w�I#h�$�v�B�i������#�O�:͞`Q���]���6�=;��z�����)v�:�`��@�ko��~���3u������
k�q�S��C�UR�ḍ���z�_7����H ��R�QG�h��L�b�X�k��^8�Z��;$|4�97} 6g63�viNf%!h�}^,�'�w"��Ɣ%#�G��Zu��¨�������yo��~��ANK�h|�TdJ:Ʃ���<w^eCL~����uL��+�:��6��{K�-�r�Y�5�
�zeR�O�m�yC$8duϪ�hgyI�"�}�#�zC+�GH� �/9��>E�)78����#:�$��u��/b8D-^?��+���Xy�wT#�21z"J�<�^�4g���&���cn�bߝ��P�U&���
�b_�l���Cќ�7�c��f5�����6#gQ\�LgCjie�%��b��`Y4��Ñ0n H�2����ަ��e�\P�W*�Z^!�J�P�����%t����N!��
K�a�cW%���]�?�n[�.�����y�\W>�d$̼:����բG��3|�{I!�'<��hdGO��(����[��2���ˡB�|@Vo}5}�o�E���z-�����q����й����;�	����{���t�aav����s@���T�xާ�u�n�V�
l�l(�+ڢ��z��{��\��5�=��ʿ���m�a� ��Mx���<'0�j{��Y_s���,ߜ�����󇿁�r[V�c�3�����ù�f1����3��P�7��~�i��$�{i������c ���^w�; ��=�V
��
G���	'�)�qQ8�a�0=�L
�� �
=H�[2��t݃�᳂׿�#�wkh!��N��M���K1�C����2��]�E��l�
Q�3���X�q�oI�,Vtr��g�$]/�}<�!c��P�̥�%|������ɐ=ũ����)��*� Ζ]4.~$R��sd�C�Y��jɽr}9��3N�E��ߥ+<4�����[���b�U�P`AY��f��u��$�M��>�A��c�ҧ�G�5��[�Saoȓi+8��2��nJ���k4��*_�����\)��I�,����w ��`����D3=�R� 3n��G�`iA��o�,_g�T�sLCZm(�!+g��>)Ļefu�p�+:3�W����NC#q���O���%���)~�z������ői�s��{��~�~�����ھ8X:Z
�oBԎ�f
��>�9K����� �B	���R����1�7�4ݼZ����3f"ӄo�'�Z� �z3"֝����Dh������ɟ�Ȱ�n�b4k�ljX&,��5�������WF�Z_K�>d����ʹ��!�;�/��i^�m>����Q�* �9�	����|��v�HB%���m�c�rn:�;�$�!+�|H�jf��RʉDB����%��2TB�*� �CԽk�3�)�1�xɇ��/�c
�O�\��V ����g�z#O�J�tx���uI�@��8��u��oA_��!n�!kw*�b�5��l�G�.�15��Z��8��tC,5x4j�KmJ:	����'|�A[� {X\��2��5���P1�WhS���2T3����3 ��~L���Lǣ!���,�Uᦏ��(<�5|3�>Y��se��iA����=�_l1o�&u"�9�@��m��	 `�M�zX���R�Զѥ��Z��<#������WdUE� 0�P������+̉���k������T*���<M���.6��U�Cy�o���[�h��<0�7#��_����&�������tJ)M�+�B�I��8����D��*���l�je��ך������rߓ�Dz�M�ݱwC�v9%!�><ȇ�����,!V�$�A]"�m����7V�U*��N���"����j} Eq$	v0��l�@x�g�6kQ��P}��z��י�������o�f�ɩ�Q�1��պ��_vR�DČ�0�
��ɳǓ2c
*D�@�00���hF����	��wB�M���tW����T�?<sU���
<���:��D�����D��,L]U��,�����_L4���2���B��M;�ϓ�A�O�x��Ϳ���P��R;gDn�ப���u�*�M��?n<��B�Ǉ�j�9{|�oW=���[j���.	rϟ���Y�_��_�cR[�-���~\,�����l��,_N���A'\��������G��E�8٦˽���C�E__<�xF7�����v4"���╧�0�������G�i*�c�40W+P�ٴ�}qa�[�M���a{�42f��� �%!��y�t�{b����pE�i�[Ԑ^�.��7�I�,�Ρ��@��u���aT�#���wI��V�'�b4�����tO�
=�.\������%6��B�D�g�� �c~�(%�8�<4\X�<oTj@ƻ��Z��ͥ":p����H�`�\�o8��x��ϿV4��4�D�k�Ik ݨX�}|�rȂ�1�Z$y�zh�[6�B�����Z��o��=];��̄qL�ʍ���-� \�������_b]�r�Ց�}��u���XۦY䴪�Դ(�z��&z�)`�(F-3s5���Oߏ)���ýh� 0ѷ�~[Y���:g�]�K��}����DR��%��蛳�7q�1��PK��<�?���������PV+��~��%�iMNTYr�aP?r�)U�E�I���²�(5'y+�զ���2|�����8�xx�D:��S��Le��#�ڈ
��k�a���P���<���>��Q,9��ӈd�`	&�a_�
�"���g��)?}�z@xg�J��D���![�LӒ�ƹ�Wik���*C���'��p	���`��_�����C*?DvY�ן}r�	H�;r�<xL7 �B���5�`x/_X���+�0c�1�24������OK�*ײ��R(����je�S|Q��.%�Þ�p��@P��="˙�%mT��͖��6m��=��m���L5࿋�R�jLxÔ4��"*?���N/���'���-�s�n��6�u
�0��(����%f���1J��q,#�H���ٵ���t0��[אs����kf��6,D�_���W�B��&^��-����WP�n��~[�8�U�h�C��Z�}��~��S,*�O�e8�)�'ͩ�ˀ"����[M*��IыJ��;�E��Ϧ�}��My��%��ds�h<��0�#��CX� ?�M�^\��y7_%��4�X�X^�X���Y5�����]J<B����T��f7>�����X�M^� ��ՙ�G(�F5ͯ��}fF��/������� =/��A��+�q�{ZCǀ�}}��_3��N鍡�g-hzXKYKbԸ�ba���<K)�|�یI���b ��~�:@�:s'�b��p���ӌ����>'=�E�4�-XNl~!��Jl�S���7�oXt���.tZ\8�I���m�/���0*�NA]��Α&G�`�sl��[��7��E�s����a�׷�s�J/ɂ��7�'�V��������ر�`�z����x�:�����		=�
%�;B���垀��C���c,��n�2ЙPٕ���~����Y�]-5\�w�<�v}�A�����x����{1R�f
g��&�>i�@{����b�i��\�s���+���E[t'�����+�	���8 �Trp�9 �K���-$C�q��!�
D6�Z����8���7@1�	�n\�l�Uϑ-�����Bt0���.� �`6ШI��e5���[��\����	A���>%jk5�&T;k�$<�
���y��}ƒ|����f)<d���@��/oy�/�vR����ex���^���[�4��,���F�%i_�M�u�'��]bē(�V:˂���/ց�<���*��*#�K�o4��X2:�Я�"�^��(u���u;K�/�[�Y��/&V�<��p"�7�W	�[+9[j�΂֦��&�~ߑc �&Hm�`.��ˀ8���;q^�a�o��\�dF ��ZL�aX��(r�JR��
떻:�>�zL*��z2<m/�wx:�P�S2�*��5\�����v(�P�`�4_[�iA� _�b���P�6e%�1&qQ&O�L�0�I��Д�b-�Ď��=$zh�]^/�<m���������LX�֖ �xV�%��g�����&~�!j�!� �R3��м��,>�+�^���-B~=>��e�8��d1�:� �I�'������HJ�� ���� ����v�����ХH�1��/H�K�#L W���W��qb��X�~��� �d�,Y��L^��L�ڎ�c�����iG�~H��/gub;^Rl���wG���v������J�+�)�\���B���3��ˢ�������cG�͇�sJ�]���P>�cWt�=%4������T����Fne��[7Ȣd�� 5�]��,}���?�n�q���k��砀=ꢅ�M�ڻ����[%��]-.��r�v�V�p�O��:�#�_,�Ot�p@㘺[zF��SZ�>�Oa⒕ڦS%�"�N(�ΈmEn����K\l*�QJ�����j�(Cn��B�K�Eu^Ĥ������s���o�?�}�T9�ǵ�S}]/����EJp-�|�A�DX�f{�ݍs��Q���!�<2Ή�QT�t�Af�Qη!x���$9AR��Ѽ�����{�\qB����"��,�|��=[�L�w�:��T/7=�S*�P�D��W�V�U�&�b�ū��nS8�^.É�	��}�C���O���3��EsX�d3�b����a���%CoB�K��A�$]6kΒ+�i`�rTd>��գ�l�2�����=bl���������� ��-A%�Z;�}{Sl~�h%��4�X7iE��m���~�2+Dy�+I�����9�'�P �^b���h\��MT���6�B{o�1���簇cM�ݳ�D��j?�?�f�g�CY���m���D�L6KѾ��Nɸ��G��
�<Q��J��}�}�*6�Ԋ��݉Г{�H�ە�bp��v�����9%����p�oj��6"�|�z[!c���To�by���m�
"Ɖ�*<Y��V0Pç��!�BQ��4��겣�TD7���9N���6,���X%l���:gV�u�䤾Xe�`#2Z	�E��XY�R�{s��6�,׶WU���IG�$�F�rʝ�DH�L�G���םJ�<V�)�U�?]����"S਽�)�1���3M���J���P�ĝ(+�gf�����\��wQЪ��T�q{�+`8�r�ZT}�sa٫�R��[#���L�mR�[l���7�b��m���]:R9�bJO:eKX��C�� ��w�}(;�ڗ�`=kwg|*��=�����O��'.'��j�N|ֳ�P�B�H	�*��)s�-����>�����k��� E��/$�blZ~���z�va��n����Y)��c��	x��2��s��H�)���Z��! K �/� M1O)�X/1�~	�=p���ܭ2?A���`rӴ�N�w�-����	>́:�����.��xw�K4_8œa�V4;9�-��S�Q��s�=k#��=c�!�� C�09��q��>����
X�>]����tKF}"����5����1�<�s�_���\�o��`|�"��9U��e���UJ��)��d�����-�Y�ge�u�,�����)T�����ìf���,6���˸�ۣ��ڲ�!�-.6wu����7헅O�.(��Y 9ϰWޔ��3�ޕ�&ҷ��Y��"����τ "Z!�PZ��-JPe��Jm�����h��G���r��
�E��59������huc���y���ϱ])��jmcWpU�a+��l���&���Yx�sV�Tm���No�x3�X���E���l(�s7����`�:�z��V�wy�-����?��4� 8~�S������ۻ�6�+�>��8�{@۰��N>��BŎ�aZ����>iҳu���{E�)�vw�ٛC��v	R{�ȟ����=	1Hr�����!�A�;�RlDuw��p�u�H�����%�?L�T�-�A#��K�J�/T����K��M�oS�`��%�1&��Y>˯ؖ����ѯ�Usk��hV�Մ%^�{�*��HyD
zbjxTډ%a�C(�Z�<<��$:���A�J����P鸝���,�Q��?�9bH���F*ܡ���v-P���q͍W�~B� 
p���2��X��y&Eށ��v�l(���4�87�����n������[�	�ە��¿�9�p!u�-£��Td ��l,�51XJ���K�Fڒk��7ʠ�h?��1�E�N�&{�������n"Ұ�ɕٳ�T<K^�+��b6	DY�����G�TVu��E��`�o�aݿ�#��A{*F�p
�z�%�����Wk�e7�iB��B��@�\��KZiq��'�./��L��W��,���dp��� �{���+�.�,z9O`�UԂ�#�\È��Đ���A�-���ҽ+�e���G��=	��J)V3[z��m��4kѣ��!i_��L@�u�n9#w�@ٛ٢@���rG,�J�V��F����K�i���!YqQ,Y� ���F��-���>P�������D�~ԡ��^W��qw-��}-)��tk��]�M�C	-��������b���D[.�����Q��+�h%�9�6�%?E�*IN�yL�h�5���0����"6�	�Ga��V��$5e)����j̍���U�hQT�kZm5��j1���'���O���*
I%L�ܸ����U�Rp�,	����bY'$��o�:������<��_�B��t���C�t`d�|Ch���
i�4���恾-�l<}��sO���T�V6�r�2rZc�:�P�h����ň�8�wl���8F�"g��:?�חκ�OV�Yv�1���]_�W�zeCa�q�8�bw��w~�h��� �� ��:��U' ZVN�h"�Y-0��o��K��2�4N���f��T4e�:P�D�a �)2v+ŋN�s�{�}$V��JC���$�d��y/HC��i����U5��hH��t�N"�9yo�7IϽH�=�T����L����	[.�O�&�0�O�D̀VK)�XE��},�͇���@�"{�Q���<�Ku�V�u�~`h���۞N�C�7�9?[�=�/���P�u�R@n,��˾����
Ɣ�`���\����PN� ��uϪ|����>��}�,���ޣ�q���=�L����'=�%
>e4�T�����z�!C��mio���S��8Z�ྥvj�z9R,�=�~����?f�_���nQ���<X�͓ޒJ��pV\i�T�JH����'��U�t\H	A6+/�dSU{���9Y��*{�#�����6����2�.|ީK��2��DZx��$���tb@3�	�y�/2@5�(�}�£{�����Um��7��*��!;ٮ�D������n�,���v�W���NgJrd���QmA�G�����ZG��q�{$r�=TwE�,�u����cV����g4������bl���\0M$̇��>��M�9����y��켮��<��Z�j`/�#۷�py�Nw	��^s�-w	���&&���$@���?٭�W\�]U�8v����]�����U�l�^�d(ҝ�`�p�6�%v5��d��SW��!3r+�]�=�;��^:���XR/��f��ay�N�>.���1�m��k��X�|�ah��%�ڠ���~� |q�HecU�1�;�Ɓ8�S��h�u���$�9Ý|h]*�Ʉ���\���E������~��+o���$Of� d�;-^kq�њ�6������&�m��������e]O�z��OnJ~_�sG�S�fo���2����n���uP;��QZXP�� �F��h���a�|4�d� P���,G�?
�Pi4��3vx�$5�Y�w���	HC�ia=�&�${'(-Z��pMDC>C�.1*w�,� (�_�Z�u�f�-1���3�-��ѤP�Q��+'���&�l�R\D��]�;,�C�ByHX��'���V��_�M��2���(�g�(2a������#������"AQp�es7b��ߟpk��9n�
�?mO���3%��+L.��C�/Va�2Hr�!�&g�������K�D\�����m�����Ͼ�U��9��K"�ȟ�"*�dϮ�x=y�>��Ԡ�L���TՍS���d � u(��=��Y�5����-#�<��L*���$R�Ǜr�M�&�`�X ��P��7 �dK��^l��±F:��� �'��c(���~w�������Y�
�!��f��F_��]˺O+O��H�D�Ք��e��鮬bX�u��c�Ggצ�w�9�!&k�H(ʨoM�"Q�_ԣ�/�q���y�$�W�����6���dՐ:�+~/a����a��s�o�d���� �ݔt��$�Jŉ[ �e�p��;��\ӴV%�i:ʽ+�W�a�X\�u���i���*���W|؉��i`7\AU�-p�+Z�!���{y%	����ǵ����A�ߢO�%r��E��V�}�ѧI��n��ewM���#h������n�h�����%���c�(��Q��j����ɪm�k�ih���c]͂-)o��,�?��w�QrK��nTHL[��m{ �
K�4���Də/;�$����a;��F�Q׫lf;��6w:�[K_n��U��B��w6�Scj��vV������= ��6EQk;:�>L_�8�p�y�#[�H���/1{QZ��izp�Z�O/�1�{�����g���IA���M\u��#lA[�����xɜHe��v~�WE�h��Ԡ���V_EΔH��[�q���Y��F�VJ�R�׊)a';d݀���Y�'W�6�ج��$��՗rL��P���%��*��o�\/�:&miM�z��;�
��k�d��_Ht|�4��bbF��ybMV�ӊ��;�ʂ�Io,I���cafFʌ�]ăs��6���i-���������	{�����E��d�Z&�A�ۍI�G�a��0�������V��0�T�3���k�a��Y�!�k�[�w��x/��3���Y��H�}޺���7�1@�p����;��^��n��}�y ���A������j�����f�%�O����9Uu=�1�+/ ̲�#YM���L�5������iD�n?��
�<%�j ��]X�to[�?Ic^��1����Ԯ�V+r�_V��W�TQ/��V(���8Ln�<��'�p���R�(�|L|P{��L9YY;��{�2
�/�2Tqf�����4�P
�C�#!lx�a��ɓ�]�7�$�1����˕ϲ�4��Z&_0���7�FaK(ys8�;�U~�K"W�*��wb��T�s�-��\L�)��b1GmՅ�6܃Bu1�Uū��"�	��o����Z�9[T[�i�ERZ����6ttD�Oӿ�sZI�U��]�Ml>���fS����j��b(S�������J�"��\���v�*$$���������BOE��>�M��T��*$�S3qK>�Ӵi\`�q����B�,UD�ct<��n\[|E��+�R�K�l� 7N1�Pq�(��M\�]��
��n���D�m[!(���N|4*�r`�@��}XY�{Κ�4���-��y�s�Fi{�o�_=0������c�5����OYM׼�?�d7<~U�U~rYCdiq���,�s-*Xy(�P�M �w���>�Պ�SIh��z�O��5yhb�g����
$�t��E�=ĕ_���`\^d� �S�RA7?(���t�ȡ��G�F�s��2)8�<�2����0z�����D^���t�E=��Զ[{��4$�L�Պ�D�������H�k���\j>S��ye�mY#�N|(,>�M��zZ���ʐ�������r ��I{J܍?A�����kZ ���݁\���!���J���R�p�]y]J�-��>�L

k�#��7D~/��oC�4��l,I�2 �
��?�I�N�ؙO��@ER�������hR�x8�ԕ�B@�S8���쌃�m`�Q���J����J��ଈ�t�-��y��O�����g#�_E:C~I����$6�}�$8d�g2F%��@jֽ[8�Ɯ��=TF���jtc�����їS׷ǒn}�����7�9�W)ݣ'�6������g���f����bo=l��B�ʿ��&�[*σg�ߙ�{̉$����RٚF�VN�]��*���3���9���"�D~��v��ѝ�V�Za��@��~�/����v��,���*�� ��uN�΍c\K�̳�VM�4%Sb�_0?�����ꉳi�Ev'��J��a�N�-e';�G�ЎjCc�P��P{Q���#� ��Z�rq.(����L���R���Y�~fu*���bW��ymr%�U���c�)���j"l��]5��ٹ;I���p�����=�w�g,~^HOR�V�X��l�Q�N����VAzi3�T�N��f�@�	�ʾ�Er6_A@�0��Q3�2���,�ԯ�����`���o�ð,����5�PT60	eЙ!.��/D=�(�awfF�-��R�������+���{:K]�J�	��e1�*"1آK�ir�n�QK�>�H�X�
���"�o����[�N����q�ۗ����C L7�탥g�8���J�#il� ���9	&N2�6D_d�B�|'�F+����<�U�W`���;z2g�ufl������
7����^���!sC��۩���Ebs�2=�>JGH��h�u��R0,7!iQ0>��6�~b�@@:AV��A�"(8B�!�WÙKej���D�M���l=|�ւE����s*8zW���9x.hC���Zs�8>�E2�sP��8�v5o�v���g�޺-r�4�^8�9��@�/E���лN�x�9*>ƭ��m�SU�e#�������V�ᔹY�	`����G�,��a�L���v^��~�Ҋ.��W���4���\�B���	Rڨ��2�Ҹ�q��~���굪C�8��I~��D�_{��h�"�Gt;�c���d�,��P�CwfQ����Iѻ�����.�����Ȫ��#���#ܑ�
�V%�ۼ���AE-������P�)�����FȞi� �ΐ�N���B��d���:1�����4���j�5X@�u�e���Z'�5��0Ȉ�r9r�ZP�.<u~-@��C:z.�.��Μ��ϕ�P���.�Ԝ�C]}�<տ!�7�"vnY~MM��h�����}Zm8f�����o��pD��h7����p"w,{\�kH�t����G���	@@ٴ:9�s����&SP�d�^s*��u��Ur�
�Wƶ|nd�%�u�ɆC�Ϩ��P��eEN�V}ɀt�)T�Up�I�W�)�2��|��V�|���I�T1�����<�����*l�+��3hq�o��v�;�d�V1���vP���o����F6o9�.�ωm���V�/�r �Ro0Mp�F�-���<X�V>#���(�{�}'�F��z[
���N�� ���L;)�O���l���-Q%/��:�#�j�d� ��'~�M_'T�Oj}6X�V�W������Q�[�2�@A�l���a]p祅��`$�ٛ�4�Q^>ս�ED8V)�:����|\�J�{ۨ��}%�DBNl���~B!#��Uf��Y�:;N�Is��(��C�fE���k��ݥ�x�+Dʟ�ⶦ��z?��Q���+��f��a�k������xx'���^W�6�7%�!|&G�@&�f+'��͉3wrԢ"��b��es	�V�ߖpg%�_	�Q�/�m|LK��y�ݵ2e}�L*e�P�u�+z�D�]�!I>�z��u�o�����'�/L�����9#w��㎙���<T�j�~c�v�&�����!�'�1��E�*�k��7�
�ذL�)�\��^wJ��O�o-tb��ʳ��V+d�M��1�i�"mՒk�=����S1�R�L��ޤ�,����)eB=��s;WTu�n��ј,�����D"��I��Mm�2�Us�&)��#\G�}FA�	��l	�׍v:N��t��n��xBg�<��T�']I�o~>O1� L:$��/�amR���)�f�� ��L��ۇ�O��-([�^{VU�� A|C?AOD`l=����?�هk�/��D�i���<tQ@u�#���_ƌ#�����+�@�bv��U������������U�����E��	Nޕ�>gN�M��^�>�8��ɔK���^�5�,(ߌNp������0d��m��T��W�)��� M��1ثw��xT�������(@zx�t�e��I6�A� ~.��"��8�W��>@�h����Ɂ[#�~P}|E2;���a�	s�]�0H���0��&	�jE��۶���hz�u�7�\	ce�2���>}t͐�"�P���V��W�lk�D�>5�yYZ����a� �ҁ"�6�OT�8N,��)��{Ԡ�u�n���Fڷ��W/R�[yJ���/YǶ����6x��X����9�/#�3U��6�d�
�)(MAP�u X��䡚'�����G�7�c��:��1���)u�{��󏒊倐�ʍ�(8B���Qm�L]�zY04p��0�IY�;�=�m�I��J�ZM���i�����?�-��&��e'5�q8C2A��riTQH�=Y j�LnjMB8��M}��%m� ��ث���`!��+�h�>3cY��� �㫯0<x��@|��B�h��D�$�!���g��ӳ�Nm���,bm��b<�O �6x���?�3�Q5D1>0���ʵ�XHճ��3�м�$�0J�	[d���ޓؑKm꧳�Q�r�JuK��x�r.��
]���	��Y����:�͓@q�NT��s��DI� ��~k�a���ÖUa���2�W�D�}ݱ�o��-��i[��,�Ul��"��4�/��i��4���>�ŐT�L�!�'�rw�Qc4�/a�!r����r�g�y:��pTg�6�e-W�O!noɺ��n g�I�&������O�:qB01̋o�:�)�I�l|ΓB�
LA�Y��<w4G�"Vz�O�|[A}�K���>x5���q$s���[X�(����Wt��B�@�<Pśn����O'�68G��-�F5���H&�2cm��j��[e�U�ޅ�gp3��~���p^: 𽵡��01�Xs��I&�+'Ջ]Z��u��h���9ǈ1��E��[ ��#�g���U��S��i}lTfk��6tinZ��qaf�x��H��8����rk|v����ޤXw�W�zٍ��:�Ѳ�E5�\H'���ꅹCy���C�\��������)��~�p�x�n�4��񉇨�BFƋjU����M�8��-�/����nV�T�W���_���"��`T�-XW����������So�o�3�}�2eϴ����*��P3�>��|#c����u|�6�{��/���ǻm�g���<>~��"�K��(�*݆l�F�UzV�t�l��"��=4`@ң�F �6����'4�|M�9�n�"�g�L�w����ѿ�:���Z��0f�D�fS�"��v��ˤ�f� 0�)u�#	��:y��M��2.q��d�����%�t
ėc]l�t�֋��J\�S��F�^}��ލln�Y��Gn- �޳y sʚb���S��'E��������+X���"��*I�o����f�n�|L��Z;�H1\ъ�;�c��/��LI�d'C�*+w��v�b1~�"��?��gf(�	���^d甩yd��,�9��`k��BKx�P�ήN�]k�;� ��ź�(�n;�U�յ���l�i�o�#{������cM�|8��M[�48�{���΀����~Ӌ��z�q�fO&�w�\�|*-=�Ȅ����A�L�5R�7+�3Є�	:f��6��A = �˰�F����OVu�ϧ��8��9F.��A�����1�T-�5yƏ��P�J���9�.�+��-�r�9���ä�	!n���j���~W���S踎����I
k�r��±��}j��PN�^�?��_yj��_S|�i-�;�z�4��D.��e�䋯�J3L�YqX>�3��dU����U1u�WQ�ُ���IX�8��	?�w�6���h��
+E|���S�JP��A���<P�q������U(VUa��
��uzeKx�����^ a�T%t�r���QB_�J͉�!҈7������{���-Br|���0�)��b/T;���
�,��~0=
��=F�2
�Ibvi��~��Ƈ�^�7(}Ka��^�}Q�D�f���U��U��!�Iƹ!�I��>O�F�m��m`���t�a�s����=��km�!|l"ܶee�c��?���_�pىWd#6YO���p�\����zs�6�	q��{�V��v��s�z��hd��B��R�qf�B}aUY_!p)��B�iHL9�fm@�K�FNH���v}aLW�����w �=Exk"��%��V>SZO�|�OJ�=O�O
^K� ;���[���K`�y�{��"mu'$%\�<{�m��{1�|5�n�o���r��6�X7������w%^�W:�V|-i�Oo�} ՞��'��>6`	�3Y,�d�/����G�2�4�'v����&�"JV�N����?�-B<��2�Ы0�^�j.�U&@+��!���|I>��f�y�x)F���p�+�m�n��h�m*�4���^?./8�_!�d�NѐT��9<W�����Y���>O���݅&�B�6_�Wn�=�9�[y��KJn$��iuC�iI�lv�ye����t�
�
T����"�_�Gl��P�d�2�t[��]���K����qQ�#�b���4{��q�}��L�S��;�d�S���D�i���.�2�Zm�U�a��(Ն	��׀G�Z��1�.ǘ�L��d۱ r6��\�U��^ ���:ϡ��h~ۍ�u�ŵ����1���s��⭒O%��!I �٧@U ۨ�'D�$���^<QԢio$0Ҿd����M���I��Q���cܗn�m�'̘���}�
�A,�Y���:�bR�婯_�M���,��ɞgO� ���蟀q2ɖΩ�y�8���*���Q��ԣ���;$Z���'�`eC�e3�E�*��wE�D)α�՚����aRD�@3�#
����l��/Lw���o=3b�s&��7Q�帬=�ӹ8O�'�ޒe�9�n\"�c��$�&�we�$!��$�x�Lc�I�W�	�(-Z��Z�k8����r���������l`��C�Eи.DD�(TD''��6h��p�LR��}\�DC6<��g��rD@��BO�/��!][1�6�[�-�Hb�ؽC,<�Q9k焲��]�8�u[�3E�K��Д�ظ?�@/b-��@ۥA�C��gh��@}�)��P����k����J��9�d�-s��B����+F��N��Uiڑ�81kEH}.i9��&6���tۧ"�f��Q���N�/G,�a�&hTcG�O���h1GeZz"��)d��g�ց}Z��p#T��/ܩw��0bc��>�V�q��ލن��QrqV[��=&v�ezC� �3�C��,MM:^9|nQGӳ%���5054�Ɔ5x}��	쬹8Z r�"��G�}�F����J�=*�tyU<��ܗ���Z�[FE]ho^��c2D�W�!  p�Hf�^o�%�;�R�i�E�kɨ;�m4�̰z?}����:2�OY�)Q\�@�K>N�-m�����R_Ȗ{�����X�T���Oc8�$���q�h����)�p�	�͕ݟ-��`+��>l�+Ε�-"՝?�z��A�_-8ւ���d`n�-s��Зe#�ԙp��8��k���0�d���cڶ)Dbi$fm����u��s�����i�Y1�4B������D/���Z�,aC'/-��q"-�Q�.F׈�@�i��!E Ru�I
�w�-e�в��¤���Ţ�ˡ��B�3�y5���?Iu�Rbf�hB�<���N���� �'pA����P��_�θ��>r �!���]H'�b��!��E�%��8�2�g���kD8W����w���-���q�-"d7ծ&0@q۠'鄜�,����?���c���mƨD?�R9�������y1�5�S2��6�ҹ��a8K�Y�ҹ�'�"�'��������D*D�`�TU)�a�:�WѹIb��3�(���oF��O=a��a��ue	�6�x��㩤E-�[��$�9&����$�k���cQ{����'/\��!3d[�͢�RSᏏ�ʷ���SNb~?N�?��& �P��I���`6����A�쮵n�r]7Hb��*�Ӯx�b�Ԧ�+L�,{��x��2z�SX!>�C����&��݉ҦI�ǺP�T_@(���&{���; g�S��=^g$��g&�ċ��P��Bi���8�2��Ld����P'��AT��E�c�
gl4�9���\�!��=�%�(.�E��G���~�������[n�I|�C�o"�߃@R&E�R)�[�u����Z����3�����wXLeʗ��?���mj�*q"�����$���ͧ[�T+��^�g�.�%X�Z=A?�g�a�!�i� q�	,����?<�)J�cj�Jw�7��}����[l4��UtJ��^��D׉��|C�/������!,�c�B��C��UvP�In��JV�WI FFфU�7�A��u7߯x��8�	���͚:�/O��� �iŢ�Sb1�_��K�7�|"e>�ɒ2�F���4�A!���P(�y!ɩ��m�	�Pn-;(7�ǂ<��`ޣ��O�>�9�����A�j�<�j*��;���f�o��s�5�1(�7g�9�#�p{��.َpg˧�!d�
�1�[��|3���N=�N�a�͊v�A1���qy���{|i$uM�:F�ؒ�����N�E	���Ub�7x4~�-+r�F��	��׊��ѹ��9�z�Q���K�9.�T�w3d���nA��1�E�d�>�µu��0)�k��9�F�m�d{��: f����a|�P_�t۴�p;�~M�2e˫�:A�w�3ǺS��ޘ>=Du��|E��[֨]�9���;J���jҽ{`�[~�
>l�Xz���3qUS+#ƀ���R��#D;Xo�rOaB���he�ȋ�s%�w�
#�[��'7��!T�`g��$P�ZN}��G[�1�4r�v{4f��G���{b�n= z�>��Q�����W��3&��4H�c~��Y�eU��+&'��������nSaL��������lݰ��~���·����~|�>��%84��\f��(��-�%�3�֍&k-	�2��.j�������:|&�ゴ�k����FF��0_.D<4�;�oՐb\ '��y���!�[4���|���iuvUߎAĹ*|�Z��ø�fѬ�$pY7HL���#N��m#ZM0,ꊯra.����g{f1�*������l'*l/���}��PH�y���=Q����j�~(�b.v׵�I^2]�[�D5��#���O�v'zx-B�_8�q����V�|2':�K�)�}6��|��
�UG�6x�-m�^/�IX������w,3��`�nf��^|��D�ҤyL���%��yD��"T�naB��٢�.��6Ԥ��]��<qy�[�%�,>�75 �#f촆�D������l	�ءUX��p�"� �t�?��T�����L26�(Y+xla��a������Is���m�:0K�,i�Pub���!)ΤTF:�/	��_�v��Y�ŵ��ҤO�dCS�c�[�겸�oP�h�ċ����4�[����_�������RE�Z@c7a����.#Ў�2w����u��/�B(&B� �S @�a�x�C>��r���gk�Cw6T����)b$�w�Dm�O��8 XtI'�2��z6�����v٬�@�a\��������
�֍�����7v�ƘT�;!?-Ǥ;���m�����;#�QF����4�h�� ��PS�Cp���D�u�dko�.�Rˎ�hJ��\D��+r�n��7"^�G{��6��GB���'����xg2�$��{�6D���mv�"xI<�?��Y¢���܏�r�v���ׯ�+��E|��WU<��aa�t�	�&��c'�f{0�" ��"=�s B�c2==][��gp�[��S����s!�M�=DX(���㴣�br�}���e�x}V�cpř����?XX�f��'�����o�C�~���È"���!��gi��߈J�J;k�Z�3
��-6���:�&ޡӘG�&d�1�MI\�,��,G��U��+���^!bn^�nVj�f����C")�0���$���VY�3.��G�N�AQ߳���,*�6�퀼��4���Xb �WN&O*�4���ؑa~��>���oV�	1��c�� iMG����6�d���p��|'v���7��&8M��m<��>o�Ð�(|p&)�����.-B/Z��½��������ꍈࢮ+yE�7�Q�$R5��o�u��MGk<��o~��Q<
�ᯮ94�l��dv;K�=^u,��.���p��|=�1t�GwjTo�{�	p���+h����8���M��y"���V��bw��)��ӍXR&��Xbk���s�\��ؗ�órT�"��0�s�����b��%k-�����^�|> ����y>�x����U!�
����XU�P��y�#Vݴt{��:V�MU�)�%N@[E�΄0�Ņy�P��j��K���p���{�R��
r��h,�V���-&<E��XW0a���A�P���g+�Y`�8��1�Z�+W��5X���<�p�+��V6
�$�j����B�Ԟ��	Y� �ͥ^��o� �*@��Y5��%J�&5����Gvgl� �;[���+�=�+<�e\�/�����5�6�R��`]�!O��8\"N��󧁶�͇�����wP�V�z�K���p�I43�3�M8,�.&�W)G�GE��sj7�j�¾@���.<%����M���yL�Ȥf�J1�)%��� %���B�9�]�C�}��#X1���U6G,�����5kB��q���q�DYS�ּ{ʸK
��_����W�c$4������"d�ԫ��Ǟ��e��8�o&���%0�����:�\�lFF�t ܲ�wjm��V���;��ώsU�q��PsT����K��֑Y�^Q��&������Pdx]d�M �vz��w�A��\�#J����ʹٮ�6	
����<pw�5s��!��j�3�S��O����:�����[M����چ2l�R��R�1wP߃�T�QiWk����D��-n�^�S-@��6�/�=[��Fu,�ҩ�L�W���3��)�P���c�w��������+V_�g�jP� c���v���ƅ���m�g���
��F2�|F`
��ŕ�z=
�OQR�bk�Qe��jn�ǎT�Ut���h���')%O��:%^��߄ѽ��N�r��s��DA�;��Ā�G:�Ě���C��:0 T#^O�������d&�g�`iY��T�%�7e�P�m��W��И����^��D}y���̯�E[En$%椔+��8�	md���Ϟ&~���jڍ������X_�2�^�5���3��$��
QQ�т/�uj�ON(���Wu��1�虝.^L԰9�ry�����cr��J��t�f�)��QM^j�G��>�-EP��B~ވ$I�ے�^�R@~��U��~N=�d�*��>�]��\�%n
Q��z�\0���7���j�`j��È��{���!��> �z�}��^4x�p��<a�)�׳DnPemm� ����.w�!L�1u��{����|-j��B�����v�>&�������v�ʜ$f�~}����Ѐ�Ǝ
�Ln.=�BR)a�:X���D�H���H�a�d[��u�f�}K⩂���cu�x�@#�Y"C��i~튈��r���+�����(E�\�w��8C�H��e|j2n'G"��L�	Ŗ��
���y@�4�W6���"o
�[_@�&���V��|+ǊK^M&,�!k��\T�d���i�,�:R�|e�E&6�s*�����]�"�mv���=�.;�X��T�t�u��|�APǐ��Z�M�,�F�"��hX�#k{`t/�
�lݧ���4�4D��#
%;s�I���G﷓S�ǖ��͖�x��c�ֲ�$��������.^'ȯ����7ܬܔ���"��I@A�Z뛠,�����L��E��]D�gX����HDZ�4�n��Uͬ$��@Z�Х��.4�e�TqK�9=|:����>ؖ
��d��#�̇+���u���HR��G�^	����Ab|�~�0���5���ï=��Gb_��m.Jb���<�g=筡?_t�{G��{���W�B 4U�CE�@W�ǞR�M�ގ���(�<sǣ�^��q�dh	��A�"Xp�
\>�eYa��K�sfɒ2�����Λ�[P7|�AY�uif�sfJ��^=kg��7��ُ�G͹^���-�����4.��&px�I�T+��no{�g���R�N�v�ȇ)̙��)��/so��)��PN�7��d���{�R:�;m�9x"�r%�|U2�Y퓤�}���6<a�2�͓�>�C+�
���K<�7�m�;�y��_�3�Y���%�D0:}� ��͘	QR���}����&���<�ĸ|�j<2d|E��8�:�ZZD����x1�c�İ�[�W_Ug�E���6%�G��X��m�8����mk����5�J�!����Rux1�dC��s��@�3���؝�2#�Qr����?���j�|g�1�T_ދ�P\r&���cĂ��+'M�W2��+Q�m���+v�E�|��[^a���9���K����*޵��u����ز�-5l"Lía'�ҭ�@;��H��8�P���j��:��Zh�/U7pΫӷ	�����UL�!���
h�"����I�� %)�F��´���̫��N�b$����� }�z[��1�0%���e6�AX*����Λ*K-��1"�����@xh$@���h{%c&.`(���2�vVy4��S�ݮ�Vw߸0,>�awE�{�eJ�T���	[j��r"A��4kMt��[�u�|yB0 #�OY3��5����;�F��	�tI'�q�u�T[��+n�x��%�zaY*?����㗂��r�%��j��?)��E�)A֖���u����;j��/�b���,�h�t0����1���<�D��O��)��z�#��b�-��#�V����2��� 	*=�wJ�W��RvE���c��H��DP�Sp���������N��]��.�����J郞��l���';�o\��M���]?gÝ=�ʨ��c*�����m�V�̫�asC�NL-"%:Y�}��@J��i���@�怩��x��N�ǌ��b�sW]Ao1J<�(�S�v�r|N��y�V7Q��fн�8��16W�����S�X�a C�R��EO�](���?�6�.80�
l�#|�!}S�@651���]*1)8
F�@n�@�$Ԋ��g#Z䋏Wˈ�/Ѩ�gc�䈭����J\�P����%<n��z�W�=��JPY�/�}�j�1{��\s�Q�M�nNA5�\�]
t��7н��
��%T��`�v?�/�$��M����� ����Ix�L!dC�Wqp�x`��8���u�@�������:�Y��B>�E���B.LǱ��j�R ����:V� ��f��d����D�x3Hv���ݣ6׼�Z��j��5��>P�X�˄�/�4��H���˸D�nf�E7Ve>�;�Aӳ�O���������E�g
�	 ^`tv�)J�>��O�o���MU�ۓ�Ui(�T&�#������6���/:��n	!;Q�?��Τ�B%���̀��T
6j'��C? �y�$u������{[���o"�щ;Ò�ZN��HG�%}�X I$Z�SQuK�j�$U�2V��n�>�|u��U� �)]�*������C��'q�U��7�C��6�#�݌tvt9��$�B��(���Ȓ|ӵ�b�
�̓I$b�_%(�ACص�"V(y~u�$x0���˙�q����L�F���;��%z�v��<��a!C�.(��i&/�x�����Mn�Nה���,�`n(���Д�̊V&s�X�\8�-�d��w�����\�G�5ޢo�*ŗF�F��9���4^�IAA;�&&A���<��0��6�u��ګ�2����N7]��M�b�i8LUAv�b��Z��Sw�,�*b�]��ԥ�3��ˍO uB�"W��2GsDj�>�-$�='�����zj'�Dh $FMrq}����Ɖ�0��_g��%��3U"���T�Y�g���C�,8ڴ&Y���<���t��>���.;�W�o�֪��[%�z�?5񽤁��-������hsMj=4(�{�Jq:3����+}Acȅ�=�2^t� �Dju��L��0|�r]�յ��=��	��� ~"?^���� ��ƹ K�
Z��}D��AHP&<��W���wQ��/��DD"ˏt�
����E�v�k�~j��#=
p.)���@bz��.a�Om�����[X��9|w�{��N����V�q����Ѹ�?ǀ�����r+_�-�<��$����=x�z��ǻ��,z���Tv�)j(�!oo}�4B�@[���H�lA���V ���"97�8�ᴦ뇫:i�2S��Z��vA��(45n���.��QV5�>���DF5�6`���	�I����fJ�@�T��ַ	�@v���{�;�!�h���p�B\f��Ez2F���o���d���멟>�`�CvRf�i�0���5�葞}<מ��!�{��_���s�]��йbn���D
�Q�ʊ���A^n#�ԝ��0��3�,fMR�!�A$w��k�r?��-��d�-Q*,���,� Jh�r��}�������7��U��-ɫu��ιT'��x�:Aڨ���e�vFU�
�{-��W��D^%�H�L�	�ޥ�#������!꿼0��z ��;^B�(8ݔ��*�g���Hd������9�E�V�`�4ޜ�w��4��~�"�*��l��Rk\���wy7`N)�I3b}�͸��
���Fq\�R�K6�!eX��%�f!*�a|�D�zYj�il��c\\!�m�s@�e�:*���*�tJ�)��#�z���o�n�b�$?u�1��!�K^f	T�@��p]����59nTD��q��x���Y�lۧ��檞�.����e"筩O��qk���a�n%���x��B6!���wR�&j��Z�]�6 �g_�$ǆt��s$��߼�i�}
��KX�:�Wu��8ш�Ӿ6t�:w�b",z6�S'x�6��e���hq-M~�\#���4�xʷ�򭧩�fn#E���Z�g�\�P>n���|X�&J�{}�	�mF�L׃Z.�8����N�Ƥʄ�{��6^�?}�	�ڸ�7<�@^�">��X	��qr'��%�h�,�-/}k���E-8��Q\Y�VK':u� (��b�Gy�Ad�?��S���c�@57�oj6 [{A}p����Eڢ򞊘S���)8J��ܵO�Ŀ�pn�F�-��v�kxX|T�q�١��r��V��ssT�<�kg�dX�$g��p���V�x��6�}�a�3�u����@�����@��d��PIڞK����JꊑS*�@������w����1骑����:��M�K���w�������x-��׵j��?�F>!�v�K�e27Nnz���eŭ��y>�*�*�9s�C։��X�ҭ�.m���e["�s=IH���	wS��;4���f8;}T�1s�=H�%�vnn9�чx^���Y��UB! �+�@�u WbD{@�P೽B5�Zt/x8��HFb�����G���ѷ����fm�+Y}��Z��!�a�X�f��#J!�%��a��\1��L�k�̃���jM��0@�������;I�G�B��#֏����0�����&I?�Uk��N�V���?��!�p�^��j�)����ִ��-Q��H9Z�kzwCQ��I,���Q��P�}}���ٍ�E��)Q{������u�(�s���ZDi�o�}>1Q2�� tn��/V��K��[����w�����e��T�'��A�;5}��+�[�af`��;cg+�f׸�xG -gr�N�Ku�U�ra�&�e��v��gj�+��O���l���>�"ݟ�1���W��EِZl��w�d��܏��f��+$�֦#��*aB�:X��_gQw%PZ�g��F�M���Q5�b��w�9���y��g��hr�:���Dm8W�/u*oߠ鏁�PF�_� d|L��^�@�n6�f�Te� ��N$ϸ3F}��pf|ai9H\�{�(�:��=�'t��eڲ&gy�&�,�q�m2x��:ҝe��!"������a޶~������|�^��|�����Y���0}��N��7Ԛ�\��aQ,�f��ʱ.{�8n:Xʁ$s&�Y��P�4�'��r:K��hw�%1��i�B{-�(��g�װ=�<�ߔj���Ğ��}c'\���l`v�K�.�f�!2&)��	���Hf`��2��M�nQ�N����-${[&�yҢ�!�'��9���m�ӈ�`E���\&��&3U6�d(�(fBV�}�L��������O�����rV� ;�7�H0JF(�DN�H�z�o��}��P899?u�M���SU�5�IXu��CiHA�����Rj��+UGUi��)�wU�C��бygN��x�As�!�l�:! ��&&�2�+���aK�K��)�yD�&7�Et%&��ȳ��ß�Y�JJvx���r�ɪ Ey[�y0k�(��	q3��)/mj���D��l���z��P����-���-%)��><ܷ�Y�r�z���T�ɼO�h_�AG���8D%�,K�;��ґ�@j�D1=xEy��8�?�=j{vԤ�f�Lqu�&R.;]B�d
 t{��G6�G�&�bx--�����z4by�8��#���e�L-�R���B4�{�F�%C��i�,OF��]�zڏVI��DSY��;�-��$��\��14]����d��e_�z��Hu[mɗy����*�� X���Q���!��X6CF�OO�iל���#�K�����nw�p�P�����K�|j=�i�w/���W�)x5a����j�X^��䊨qY}0�d�c����~�D��:O�VԄ����2����126m)OP^4=�8�1H\��
�ݑ�	4VuH���.��!r
,�3�\�x9���6�k7����K�����Ҭq�R�՘@o	S��+.j�+1WM�I'�j�/e�z	����pb!����I~>M��. ��lKL�说�A�#�n�fU��';1Lp��;y�qI�1��R�W�&_���@�L:"�N�����Ot��	"F�}���}�����s�ڕ�L�D%�Y�A%�W��
��:M�I������c��o�B�!e4�8�����G���H=��%a[�8F\ѐ����)N�f�D����=E�uO>v�NT�!����K��~�����|�>��,0�"��M�w�]߆6P�,�l
�Dg��o�����(�p��X�xg5���H~V�~�'d��JI0U��e�g*�V@�7x��>��J����xn\�p�`�L�
���w �OԄ�T�/�[�q���B��ѣ��١_,��qJN4l���ou3,gT3bkȥ^�P>}d+���@�u���u�c����j�������#��0Ŕ�'��<�&E��1ra�y�R� 4E�q@(KK���/�lR,����UKֹ��) ��Y'���r��U�Zcճr��g��}^:p����;jw��+�-MU�xY��p:<���$�A tr�o���!i�B��ǆO�XTN8G\J� ,mrYxC"���M�n�e�)ܹ�oY�K��H,e�!z?���M�柔4��Ż��;��*��(�u�c�ɤS����Ɨ��HX��5�PM@ǁ��Q�?�2���q��r4Z_Qܻ��#���p�Z���5-=���E쒧�q���O��D9�%X6�FWۍ(�"Ֆ�gs��-/�����>�8�L�?��Q�����3ϏC����!���|c������k	l���>5�L�w�(�.ѯ�/�W�t����ZEh�X����*��sO�xR�&���|�P����/:�v�n�وrBd�$,�UE��a�۳J�'�B!�[6�,���V߆��L��������5�MtQ ;�JI�F��VZ�g��;���/Z�d���B�C�o$9%O�in�Ŧx������-dZ�T}�-�]����ؖ2�󬚰D�2� ��!��w��\\����Y�Ɓ$֡�
Q��U�*4��-��K7r�c��e���+w g�T/�݆X%�ɕ�St�T���x�}�Rl�����`�8�w/��gp�>ռ����x��rcǵ�f0�%� `#��Zv�����
n~�l���H؅g�fۍz�>/ze��|b:����*۷N�cؓĭ�R�%i�� ��S�wz���@�B��f7��˨3@�,f�li���	���x���̗t�kPޡ1��6YIJ��w�U�FD_b� {��/ý��o�!��"�'�)���**��	���M!�1��IPx_?)'}N�ߙ<�P��n�(/����4OQ������Xb���$�u�Gx���PY'ް����S1�4����z��۳��M����p����"})�:{��E��ҳh�h�@���G3����Rى`ř2�w����@�t���9���r��?8D<�un>,����Q#6�ܪD72�)��j�,R���&KU@1!���@�Ŝ.����	՜�h��P�내j�)��/rѧxf��q7>��-�y�8�H�C#�$�פ��\eH+�&2ڞ��r��o��v���F��=�>'�g�Mt=n��.k�;xT�)���t��}_�S����'e:��,�q �Z�1���mQO�K�r�~le+��g�}��90�m)x��F4X��#�����Y�~�#.�-�&}�{l��%+��Z���D�%�����y��mH��NA`H� �1w�SZV`�t���q���i��>Y�1�c�2_�nd~7rX�s�S�$��!'#*{�G�I_��&���6��h�6�_*�i�g-����K Ng��	4V���#LOLܔ�Rj�.�n&�0'8�z?��ٜ���	g7r�P|�>���$�W�ǧM�B+s{=9�~&�ڼ2�I���B��@�0Y-��H�,U�8,�G2�����UP��;X�$WT`<��0�,~�.�����j�q��d�O1�I�i�VX���-�-��-���^��|�S�)Dh
�6��J�K&F���g`3φ�M������9�0�@B>=d�|<ɍ��D䨈M�KL��y��1�b�XV#A4X1?��n*	���=EV�eT���2��G�% �C�U��K��!L�=�<,̇"����[�l��m��H~�;P	vI�R��L�h>zgz.h�8]�!��ŵp��j���ܸ}H��j���{�e��y�س"R��.��w�VUݨ�CI��y���u)H��e$�仆5�����d�]�9�^K�K�Ǒ�9�[%r�3/Ob����2��\H6�Qm@lJ65�]�kP�VS�DT̓�� 2�G�5^cF�Q�3���B�i���I�%�!�P��iSF��Ʒ�'���e	�ͮ���Zg�_����l_���M�h�?Jvn=��`�.���H4VF����'R�
��H�M���:?;�����Q�ol$�Fb+p�ka�/��;������F��pR,}کv�X>Mi{�k,O��Rj���7?Y�����2��ܹ}����sG�7��k%ʣ��}���Ígc�C�z���5���b����Y�u�B@={�ʰ�3��f��C(C�|WX*�"V�]�9؃S��APC��G�t&hV_���U8I�̾�-�#�Q:�"���X�i2�Qjކ�CD8����\�w�ɯk%�������2���4�i�%�NV���on�)ߓ��#W��}�^h��c��Z�s�mv_�n\P�5�D��^uE�����- �қ��P� I�����o̈��p�f�X����/��`\Ot!��&Fu���j���>��Ʊ���Ϻ񟿨3�O��Y��B}��e�k�L(E	õ�&��Sh���膦�?6��UY^�P�T �?j\�@�� u�̓�J:ۈ�x����r5E�.J[��e[c���n�2xUt
 |e�,��MK�g�ab�ɊO�2�v�!�-�������n��/۬�;�T���u��R��g��4���#[m���uuƷF�TEU��ܾ>]�`m	��� A��kd�	�G�J�R�����"�
�'.K�!��Rd��$ ��KPp���$,��v�A�e�l��*�v!�Yc�x@�Ϝ�ή���k57�۔���f�g~|�/�3T�^��E�s#���jH,pT�b�!�Т�)�g�Գ���J�Y�w�G���)�M�l%݇�[Ǝ?ĺ&�{>���Ki�q���z�]֟ka��X�r��Ѧ�4��L��n(P��-s4��v����NNt�w�O�.{��}�\�7?NUA�yq��Ɂ|[�7�2趴�e�{B��0a�^?2��p�S�N0h6� �������b@�k���$� /9A����4��Nl(��7�b���h&/n�����w�q6#&��`��Oޯڇn���vI�hQl���sZ(��V���p�MD �C��b����~~�$JE�ϛ��׻�6���P���Z
�S����AZt_�j����'M;7�$�J���DX�~^��w��Y��A-�Nx`z�pM��T]t�u���2���|��Y	�[���-�H7o�Os�\���I����k"���9p{�#��9��y�:�K +�-`�M����c��#D�&����*-��g����V�o�ub^��� ���y[�SC�I�@z�y����9g�9n9��'}Y|����@����ɲ-�Zu�;^�Q�%�f�7"[��:��㱛��xW�u �F$�$$,��d�Z`��m�r2��[��{4�l�dc���C��1��ُ���n���U��8 {��>MT�����f���/���"�0���hK�:i׀>s�� �.�K}��C�ȿHf�r6R'�F�F�+^��a��t景0ڰ�{�2��c�T&6�M˲�p�)���1V�8҅1��>[�I�<�d�I�69K�-iUA���u]�@�{�fĮ)-!/ ������d�B���1@ؑ#�I� ��wϨz�[��}55��="��]Z�Q���>y�9n��w9�S���>_}��R�m�Y<H�V�(!S��_1[E�|���y����;1��ʐ�͸�����кx�W���:.ډ_��o''E������aȒ���s�E�k��I��Z�[(�H�g�~R�B���������Q� :��Uʖ�LA5����{=���!A}�'&���3�6�B=E�(C6,	�BE�zV���Ŷn^$�gZu�m��� ������޶����hWԗ�]����r�?�4ei����4�#}�4��A���N�K�U��.h�qϧ��t���[�$7��`Ѕ��0Lc��0nӺ�� ��z��ugwr}G�K�rٳ�}mB�(���R	�)`q�d�!��n�W^��R�{��λ�RO���aWu��弑��]!���xK����;�򡒬�S/$BP�����ށ�wb����*6�_��YMM��9��b_���}Lp�T*u���]ġ���^��ÚK������B�>^(�]g݋n�	X8�P�X
N������B�ޚy�;t���Ðٜ�|s���.��[Y2G`��W�e�`�a�|�%E���'�e�����'��(��m��4��)y��T;�*�K���e�|H\<ș^^!,�U4B�u����y��4�Xe���{n����`��o�F�W��e�A�0{�F�Кh�W�5*�X�1-d!RqU0a���[��
od�:�D"ڞa~���#�(+/�P�^��\S����yZS6m�0}�֊�W��ܞ}�}�*'�� t%�qב�p�d��G!O>`��7š�<��ڱb2h�ګ�(�-�̡�Q���:(ٌ̟<�YsEӰ�}��l$��}��x�ڑ2WA�33���d��-�Qp���1��<�(��)�g�[�}��e�-7��m23K��.vq�D._�U�nsy����L~Y}��Џ�;p��`�����9:[twx�� R���9F�GVTq\��a<������H��������
P����� iᆀ�i!d4��!r���UМG�ujP�(���C���/���e�6|=�d8�]����-Sy�>�sX���yq:��wԼ���2P;h��a�u7���`�����Y��!��Bոor5�m�'=�W���_R�{VĳM�Yy|{�b�Wz�(qZS+��dڿ��/�ǖ,���?�t�|�M�Yi����Ku��a�u"�M��k�s�(W!�=�h+0
�*��*@T����u^B��gw���'��h�%_����HE��޹D�����ܶ�Xs���Ą8()����P�u����(��MCt�y�bR(]&��Cwr�M>�1����sz����m�s7�O���_%{p�@�����\�bE����YD/Y��"8�Q�N��A��v8�q��;gFkT \����`	O$�B�!84�9�Pګh���ڑs���,���7�IJ��N�Q���yS�-������dK��A�xŢ���L���9E���Y�3�mPs�ڌ86�z<�� /x�8�x��Z��X,Ҩ�|}�hd��Ѱ駂���pP5$�g�XRN�@�m$�~S�S��ת�6kQ�TIX�-��`0�'K�۬#�X�\g��iu �����p��	�|�n�;�K̖��,yD�|�����
���4�	�B.w|����
۽(ޥ���Q�pL\��5�K���ؤ�Fu���>��{q`� 8������D�g8�Ro8�X*�7{�uʁ�~���֧�#8�y¤ݾ�D#v ���=�rʟ;��銼��|�z���cH�v�Q��\"��T�^R�/qT����rN��'s �I��*}��e�b�b�0�F���<y��`�Y�F<�Ms��Iw.O�ɕ�dynq1A�I�S���6h��W�Z���k��e�2A�� .E��?b��ar�����3ȶu�P����=��M#��0����0��,[�����%�Qf���I�i�
�'r�|�X���Y���V�wls&�]��lA�"d� ��RK
>oW ������}�5���DV/��b���e�w�Ũd�����`^�z�)�M���GT?1/ß{��;�0�$����3��#[VH��B� �.�?}�����\�-[�62�Z�AWX��AJ��{��y 9��v�t֫F���:�\V	ρ,�#;�}ӱ�r���^�0�_�!�l���.k�ױphy��_��n/�b+���$����kG�&�4��)��N��D3�Ȧ��sU+��̶��9&�s��X��A1}�+��Q�p�|�w=Q7��B��.J�g��U�l�u�-�9驜�D��`E�L�3h�'�/^���-�
�������v�2�q���I�����ZW�nҢXM	�Ԍ�g	vR���n�aD`k�b�~���06�}�Q���*��dt�� =���Fy�/���V��#�i�8F�#L>8�窳�X���T�o�SV�GCQ���������5���=[�u��Z	���H��p*pֹ)�6�9��>�\����շ, TdX���Ṇ�4M���d�A*6^c�Z�"i���,)͠�6����_:��i���xۿ�۵�ټ�`�����g�,�ã�|�ˊ�Y�ls�׹��G#!�	̝u<g�]�	�(�R�����?j�0�~կ^N<g4��f�:a����	����7k�Ex쀣��y�*%q/� 5�/�4Ot��]����}/@"��I;�Ԩ� !Ye��`$;�f�ϧ(B�����Z5�H�Ws-��c-s�ͮ�9�S���9����x�D7`ܫ�l�kI�yK)����I���M�$�A��!��ӂ�4�{�RbdB�L4�C���t�+�;^	t>w���jc1�!;��+x.�()���n����v��2A���i��a���Y_c�G���"0�)_6w\X"���q����ˆXuzVb��k#��$U]�Uws�жV`d���2�5$s��4��-�zLA$��O3?TN�<a<� &�qG�0�Po�̫C$��UB�f¦uȣ��3w���_u l��l����>����_��Ս[�T@��i��p�O��A�7�h{B%���Gp���b �$;r����F�s�]� p����&e�˜k�tt��3VV]>�ìY�C��ER~�堿>0��/Nf�k�DA=���z1�'�+�F�͛�������`�7jT�~(R
u�qr%���������l���!-n)�RHY3:n���E)�0�y�B�3H"<@�o��#=c.B�F$�:�(�`���IJf@�H����H#���بG�.>Z��M�Jl�-�K����G䦿l�2.��D5K�9���b��L{�G�iVà���C��^�x�X��v)[��Q�
��FDBE�6ʂ�lE籄l�u I��/��,>9�=ֈ��j��n0.\2�sv��Œ%����]>��I� s�_�_x�
��JsY!�R��n�*F����9�m�	�-�$�P�M��Q�9���r0��Y3/u���zKk^q.��Q1�/�-�ΰ�B!��Ҩ�@I�Čuk��i�xm��o��kE��?�L�f�$F��!�
��SgO!입�Z��[����Es�,��k�Zz.���U��<<��Aj��l�7�	�e�2�y�'����WYm�{߰��h@�'Xנ%��3*�q>)������6G�G�,�e���q']t̂���E9��Y2_r��I1��:ů��%��Y#��B�<f�@�C�iOE�-��!���C�	D\K��yp�Ť�#D�$�@0N��C����e���௘ұbQH�V�Z���XP(	ӛ��F�R1����LQ�)�8:NEȃ��`[�+�����i��,(�8�[�,sY\5���EP��~�:j[�m�h��P���-J�M���rͫ���s,!A֏����#G�8@�޹�<���"�?�*nE�D(�x,Q�#�bq*=f-{K�3 ��C�(@�,�
�w;R�_���At��b����Ϯ	z��("tX���֌��R��}�n�m�̧��+���Rv�n�ݖ���E�̏1�f�C#�a��:ۘTBCw����tKT� �����F���?<�cd�W����S�٭���\z?������+ap� W,���p�4�����[ƚ�$� fGC��<����7/��ߖ�<I"��P�;$r.����Ȃ�(c�ȃ�0m�0TԎ�����9m+MY��Y�~(��p��	E�����)ҸmⲨ��{kg��"�MS���B=p5�`v%<7���j_Nݽ#��Z��s�+�I�xܓ\Lc���;Y$1��,���W�y�64)'��\�0s�H־�u��f؀uO���X�Yͣ6	�U���'K
�>}���Je��7�%&;׵��w{7n�ۓʀ�OM8�Ew����bv-7a*�:b�u|�)qr��Z�͜yMyxy�����&{� ��-$�ft�(���s�Nر��s��C3�Q�NE��F#���@ş��{��Ө"��)s�:!;�g��!�9��0Y�$"WO��ض�+��))�һ��(�_&� �V�s���T�l_B)�_C��j��׏��
���b��g3���H���T��2,5[��W<te�r�EREcj]�k.�J�"#y������/s�h�3j�g��@����9ᘁ	�!%ESA���z���T���a����\�9�}���8�]g�G0|�n�������������$b�M��	��|��7��������]��9����:	ȍ���L�q��ۙ���3�>����4���e�s�DdZou���84N�ҬfAlN0)���g�)(ބc u�r��l�o��0H�{�ᬾ��;5q!|���/!�u�{���eɡ��P��ϥ@����x��DH,��.]�O@�����y��:D��2�嶰.fv��� �>5���A�B� ƾ˲{����a*�I�{8YD�S�;��4��Y��C����y��t������E/�L=�P���,[!#��+��o�c�BOHƐh����k��ᡵ-B�p�����ԧs7�n"}�9}	_pv�=�hC�`��2��A�9@�,�^I������i�����,�g�M��~��1C�j��ya�g����kl����N�Tӭ0��&�����\�Xn���a3����sS���~B0�9�v�xW�;���ݔ,M���E^���;3�0\N%���c��)�i�M���j4�bL����Bԉ��3�[��"}���g[���D�	|F���	q` _�=hU����&m-a��Ӡ<�A�pء	%R�4iqݔ��q�5��4��G9#kcX��ȧ�0������W�C�Ͳ�!Ȅ73=��Z72�N�@pkJ���1R��:�e�߷(����G�w��W�)�vPZҊ��!�z 7jNY�*�yկad_ǌ*6 ��W��$��^"N�[�l�_(��pB<�č�����΃��b�����J����O�R��'Cx�"h-������wA���
I�X=ih�4I`d��0�#��EN��{�qA�:VǛ_�+����&ڠ���*{/V�d8�u�f[h%I�d���qCV9�!�1��K��]�TM������I k*��u�ԆF��s��	�WOq?���\������ے���b2.�L�G|�1(��Y����\���u�Wse��i�<%R�R2��'녋���f����O侭n�6[)��`�=�]U\��[�4�A��|��J��6�T��p��|f�qVL�Y
��d��߁�R.Z�[R�܁����W &�8�㿛��#� #�7C˒�$�f=J�	wv��C���*^H	b椁�_��C�KCYQ����+{���O�/��3>kr�t�z���5;6W�3"ܠ�<t�^74��cYy�[��܇K�ޚc>,]��wK�{dƸ/�:��e�;�Z:nZ�G5�5Bd�p��J��-�4��(v���Oc��hv���&R�8y��Q3q�C�>��f��W$o�_fF��ccy�$,������x��L�a���UMgR A��H�SvVK")�u��x)X�Wv�@�� �X���y��y�у����e�m$������Ԕ����X�^>ޕ+�qs(���Lt�z3�y���~6oV!����S�����I��IHϰ��12/ *B�ٗƮB��`�7k�Z��d���Bl������&����u-3<tn�V!���V=��1̹��^�r��r�A>��D���18�VI9��>5�z?T�kse�Z ��6��~YPA��.Z�F����|YB�׼���ϳ�!�#ƌ�{�q�3��tUG�\ b&d�8�s��T��;�;�j�(4h�f��J��b�g<��hy(%��<�&lu��Rf-�0�Ǉ�D�x���37�O.��u�?�J|.�ґc���p�5����;A0��Z��$��� B�'�����q�qBQ���}�3X�Q�f�@����R⩡Vh��բj������OX��IQ���ḳ�r�3�3�$��R|6����}��J��(
X��������&F�4 �W��[[`��:��ex$���X�J]���Os�����:�[�͸t<�kk�w�8i��I(-R�ղ��q#S/c�wl>�"_�+:�.