// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NpYvAn+Tl0pNhK/WPfVAtmGumFFikhlPmdNnAlg7OmiphEdEWuI+89gZhSyocVWr
hGDiR8XYNvW7k4ufktkuMAgZ+SSsOoDyJUeMDK5yddaGz52R1QWiPB50KzlfXOEh
sHd2TgJyX0hUU5cf/uxBBloGedVdhZ5ZzEg1YZpajaI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8512)
STMwfd5H1ZaG3VooIMpO6t5xdMp3/9A6IrxN1039PklpnM23U+owylcSZJc1AweS
OYsiIJQ30nd//a0BGYeKjp/BOcl5njWzyD0q2w37DAAaKGUhK9vmDdPzdlIxQKGO
5DxZaL5/ZzPeT9xsTkNrMABPL4YnFLYD9XKHRhxqHeqYjLA8AxuVz8koLu0SwLaC
RM09trHpz/TKlg98y50zgtptKx0oRT6xvRwEuNg0HeItUep6FLS2Z1/P+LJMo8HM
ab+1UvAbWIV9BoVojgIZIl1iZOKhu9Q0C0gYP8rOBwXUWlZO/l/cIbyX1QxnlFM9
jkZrV1fnj0igpeTM5u/7hxMba7gYLZtYlzqstulVkgE4t0LMe0Wk1Ak17J0cD+Vr
pGecgtuHV6NYDFgkMOuKVt/5Sb1iObZixuGexDYH/NM0LvlxV8VmSYMLDrPrr2sh
gUmWBTyu5dIbiq+GatS6wTkyamMfXDG6WB9wdmxGMP4Cbkpxtax9E8jYxFX7ddHr
kEy3o+byz8Qtc3SwCQ0VA6Z20rOnopt0Ms0CU4kCxAlbfqUd63hou//Qo/uUUqNC
1G9M3StnXcKlHFX6pPJ0vvHdEBjMEnDh2YtaD2yEJdPdTmb3E0r0bcD1W7dadrmA
oMPQxP6v36M+QomcvjkozswsbgUdaE1bLkjH4oHGgmK4PCuCJ7oZI8JzkfVhFrXs
xbHoLhJayeM9RlRQTOlGoSdr0jaTDvBOqJAEgayA++tuvtUfhW8XR9WXYJ2gmsKy
E6O0aTUO5rVsn5sPocb3amRaynrMUkjAaCAUaoZgOalCNMtldAG3mhmvfFaRrg14
eC8ZTGZwPjXKlRnGIzToN5K9Z492Vf7Evqldyz7XjaFX4SQzTMQ+KpppC3qOThon
fSFL21AGGexc8Vvmq6v87cGQUHMUgfByOAIF8xZ52sgubcFUqhH+4qorq9dwMAw1
kX9d0W8zidfbZpZsIfsYIDsoj1Q2SxyqDD8mCUz6PynwuukufYqFfdvp11iEhaA3
Yo/9+0jsBCSZ/lQRVuy1M9OSrDwKB5yla3QFXJQ6Fet47bxR2k1D7VeBRmfZpcFw
u5qN9RUTshie4JE0xNtN079iYop3yhhH+aJIrAAWMcgduBRk0dDvHCceulQFfmdW
Ohy+wi9zh+6S30chckTLD8nOVVamhfJ+heih05q9xblU+eaJx7NI0PVtQqRZh/Ls
TJRzBSOawz9hael5vFdUBElE/FHLFv6a5eNKmRdKh5cDXCHlkCXlLf39uOLZFf7P
sW0hurDWoWcZvpO+v8EzArXSpD2jZlhYM+Xs527SQY5bLguUmgxuZp9HtoQPG7cm
XupEomLj1HBHH8yk0Ilv/Z+z5WIzXU4tuvF0VbrH0v5tviCbzu4LPh8Z4O5SDINq
IqYGr8jMQ+sckOT9lu/OuEP7Wz2fWdj/W7WYYFZiPwpyOJmMU+o2v2LbmJp7OUOk
ozSKoSbwNpbqmtm5BSEZ/nahZ3RHKb81ifCSeQrUf4BeNpctQ99XvIEIoEbeK/HQ
V+TFzCWgmQ3n9pAt7G1H6Pirhg/zHfroqKAs3uF1qrXW6ZbOVERR5kqsMHvYdjQd
+2uPsaZsqpB3JUKVHp27wL8DVttpyBuR0S5tf8ycvKbAPDm6La+TNAKbZ/AdYXGU
1CZOjXn7zIUdwDS1n86WysywgzxvVUq++psN8gY8yG7Zs3kGTwzpmx5Me5ILMgVX
UFcFfPoV7bsSp/ZcPRXEIRCcgFQApzOKe5CQ6zgeezd/s9ZCebvQkk4+MDJRnEoF
Zwg7PF5W3NGbfhHhuXX5RzFNF/ulusRactXODSHxZY31AGYGhxj1bokGGYWgZECS
w7pdG28B/Xde8DuOpmotzf/mlMXRn3A0whMS26kCZBYvCEUCGdNEVHl0hJx1/bg2
X6vOIimcYswGjOOwPr2eg751Qa/d0sgekfFez68gH/epZpJ+HzJfX5YbZ9UM1nun
gNvlucFjp652b79OVtXDF5k9vzEePam/AgZi0bwD6UEWRXMPByoI+FWQu3QLkfz9
iMIDn08+T02byM/YVF+7K4SMY6aYsluBSs9yoRBVQfLSO4dIkSr3vKSW+30uiIHD
lDYfvjDSgWk9omBy82hEyAvncaysAASugMVF65SRDG9zJO4/+wHvSFVtx4aZPhPw
0hOASVCxKq/Q7ihBg0fbYeUdGlof+pId308HqMR2OEDVHLOrdcyoK+i/KXgKNYLS
COL8yqxOezeeMx/3ZYkDLVFBFtxhkpGBOr9gQV8EfXp4LTE5jgXWtv2WPEIVPX6O
OYth5NlFSCm98YEQzn++0WP1p0R/G/wcqJy2DRErZOwOdHxEuNVGFrAOwekC6SqZ
cbJjy2QPuhf6NaP88Dhi/5o2rEuP92pY4ceAT3qZXVdeaPrybDU7atNI3zxs44vI
Aloidu1hXV0k6BfOpfhRZTaj6cf6m39qGBuxcsBTGGUNB0U5ZH0wqya5XY29dGhx
igXIHDxkmbAIGm6O8ilohf4Sl6XG5YYvRzU4zFnwoFBVCeW09CX3h9r6o+wr2r7y
F314iL07/FCWSLM8R9XFOH51u6s0PxFq7rqhUbtQtGbSwcj3RfcqaMbWmDdqSoFN
cfNudx2SYrNjwqugbXlMZCDi0j7yc/DMjKwkt6CC1kGaKpt+nTm7SmsMK1ZfMGji
y/oXy4x9R1Cwm7tXcV7sQiupcd1oHh7cZu6A/9QTxaDAvyS9YzA0dMaxCe8SmZXk
zOX9QD5himAWbTOdCpa5/T+paknontU0QZMv2FXUKCiE7yZdQgUzM8idfGNoz6lL
V2cvTUhz28IwLHUU3zGkxCJV68UdT8V12cBqk7I0PuYctR0ZGLtjZvpt5+FSQiWO
sbxJSn8dycQv3cROALWEZBOjc77yA7K3xI2gW5Jl9i0ZSJgAWGK/92sx/vDOtc8n
wfDl5SIUJpyNHx3qKdHpUklFecD4gQYOG+JlSKq00QlaMmHd39nk/vEq/6dZquiP
+68SbBnB0PNr/EvTfUBGGuwmmM+d2ch3RgEok1vDe/NTP7ZJA3DNKrVkjodeVFrk
qkWvUABdDWQAdRYU+8AecyYkNcgVOe/ZOs8CuZovLjZ+2H3lIr1YHjgkBxezEQhL
+6QprVzxyg4iwDN6lqMs/Pf1CcmuqqbWaA75X5w6wBNudHK+Wxk4k4auCYDiC+y/
/rjCtXyQCkvlcrCWuBFdTk+dYtCblR/QwsuMA2XcBqBMaR9ClG44W22hFCxEYcxc
qLq4aG0yeIk4KbEZTieMrtGbYyrS/0jG81QNJuAmhRUxCB1WhK7EF/i6+7PrXYTe
iHLd1ddYMJr45fhJNX88OQFrbm6OABRx2YCw6JkWguYHS749oVO1wHUpTec+kRbW
xXkf3W4eCd1+WHPvCRPuG+rm2g5Uvce3i2KB8hwsAtGEZhPH0Xmss1Y09Pg/FeHw
sD1oHbwDB6rN2RDJjTBSzT8/k7x9BWBaunaL3W7w9Ws9TiUpBOeHHxzCIIerJ6h6
jYq+r0hGptl7jWNEPXAj4OWZDqSw1FFYL4zudsZobJbtVaMgAaVwtzh3rV5gT/bE
v7gRpGVJih1ZqZoRvulGhtvTeWVwGT4l3UGl4RkW29it/SRoy0bUnJkrHsesH798
cPch32c7AfcouZ4HyllS94YNK8dCl2unMXbKVtc3OWyoBU+VAJ92xFETslEGq2Bt
7KaaOTLHgrLMPY1JEseS/p1RRMQWKe3YEmqCnJnQDEKBA8l0FzjPX2nMov8dXeEL
B78DjxNQ4z0FlNvk6DJNJyRBLAPjlPgUQiguJGFGblQgthA5NfnyhP0UORlLiQrW
tLxKpj/7l0h/3sOxh0FzcQ98aV0vb9+0S3hgN7w8Kag5ZouWutMo+f7u26gzsv0A
9vrfPfKP54PJM5mQFqnk8GBhUhlaI9wTzP1pTl2CTWmhgy7Qsl6EJhlhxOuPZWjg
ZurrSWHPYxTyfNnnkVhq5JD0tILByeT+cRuAjKSry8zvSfEuvLv3lFScH9QkM0Ak
caaIIqiUzUC8IPM5FJJeiWG14mqYFK3IYWRPUi1a6pdW9Vxm3O42vZQ+LXaWAigb
/YtD1sOEXbM3/LGjnl7cQXKuo/SM+JuvKVVJq6dOvq9N8AsSv7hW+J1SBFYgv3Lc
nqTrvT7cdqhBhNiXEwuXm7vImYqp0DWjhhRvK8mZmx7Yl1YRhHIYWns1yGidBT5k
qXdfOS+EnPAGr5sVKcn0PLAIdHSH4aQK96bWqGfn6gwFUa7pAlZ3NbENMUyAjFzG
2jhVWcAyRNV1+An8DX8Jjkb+TYaHg+TPJpZ7h4nT7TDNPKJvc2B70lxzYu4mP9+X
h9lbrF1VxC2uKvytMYF/ymCNrSFIDn3TYZlupvjA496TAnJaeewTtSUuBDoDHks6
MouaJZxgGgNTjRP6/ZnZW+pdMnaaCnVxNsjS5Pmq+An77TbEvBplF/I/lUGJdPaD
d6xUz3MqIpD31zVf3axy0KV35+K+u3VTS/etRUxdq4G4eczS/8xXrOJfrU0b75As
oXUTWhexRHXQ5rcVYcxNX0rAKmxdbpj2dVeHHw4+N34PYdnoOip8NwSgmBHjAGgy
3zwk+iiP5lQBdeKXjNvGRMh/qrsGQOUdzBslXPzP05AV85U4y+yjEPgEGzrRe6og
FuZZeb3YvwAaOJHyJyV9ppT/66mgUUzG0QButR0gW4ZFez2xqgWq4hrSFz55LB0y
8i8nIUcsH3De/bH/tPUk1nRv2n+EBSj0AGKuFbdXtpOJw3ZU055sOXgTQEYu1EAF
UPPENysi9PJyMsq1747fnvWqszWoJe44lZKS8C3v9IRooM/2q4z2mkdBm6t0s2uM
7m5RrovpqUWahxqi9NINV1C2N2P0rQS8bT6kpmKLgPcnk1boUqCBToRR9+IIR9bZ
f+clkDWvf0iPmU9tLKu2BYhuAz4H0WOXlYTx8cDbbhD+95or3n2+a32ys1GppyEU
2/r8FfvBQFe11jUZEZcEqTnk0mKz3Bv00OlUALVtItmVHV6pIa7GN41e6yEIkDpt
5ool71cYws+Pzxu2LfRkIIfDlHyicjShKOjL+IEDqfkYU6AAy6MOJ6v+245MLwZ4
lNuT7rfv6xaVBvyRBo1sK9s4+y5tuPuDdT78CQM9NEAzI53LhRQuhl/4RpW/WBWI
KBqibeXSVEI0s+uV0/Z2T0Ew4a8cnpRiAVr5WkUH5OS6/bBE0gxLvharGp4jzhkJ
PM7W0B+PZufg5poqZoo13cAFYaz9wXgNiiOPg5P1aDrivIn1LusEL77SmDNdq1YM
ulCtIAdjuwo1IN2VUb//aqhKHkW+oTq1fupoHOdZ+J1bUJga8YiLRW7C26iFo23j
NvmJbzaAFlSaKJzxSoe9nxtGqcqJ/YR/PEl9jpCOF5zWLnr9oJiTOQRGZPPKOCVz
p1Qe9clT2lbTF2JcVxURxUjo+8MTpJSA1C+WZLrBe2ZMzDYrj9wpXCXrnhOE8jT9
gp+XfXbXAMBPLw+WskhuEBqiz1WuLkm34XVsUovhWr60jEFBvj00nulI22EEqxJb
VtXUoeFVh2RbMmK2CBqXgLpbjBEFnvc8hy0eLl2t/X7os0d8UvpSiNQw88GPD21D
QInJfbObgc92dMiMxp9ffZ6yfQZ82F6Xm1MjUlIV/eF04DTOSJHt8f30wosgOVec
uQh3dyf7vy6yYAIPqGo6tMGDtAr7d1+yoGh3Ee9ui8gFXcGFs7QDnhAe0nM22OxV
pZ3tm6kX2qgbwgXZ1khHGg73qlsLcIqXZYxbQ0/SqKbhedfkh8nnhoX3hvhjWdLr
YYu97vn2B92HzM5Tuz/pppuGwPTBhpjTEm4cz2ztrVMrkhsNf8/ODMLLA0EBfIbZ
bDPCXgWWSxCmrS75C0bWFHvuElFEa/mraRxjJGDVK+OSjKV2F1CEhqKPyh+kPwj/
zQkwyhFXuLGoq+Y1GOLIlwPeyj6hROAVfdqlFPH8sRzzwtl1f5lyh6ve3LhxGbre
ZIc1sukcKod/7ltEzwN3EsLrFCwIaxAyvtNo2ZvqOdV63jxLuKf22/3qZoO05P+e
BwvhZTx0nHrEpVkaJHEvbM74v+cmGuzio288vhs/SaZS+FGWNmQKGela9tia30B1
tBQX9NEGXuzIPy79pGcyiMRdzrCDR/Jh49hKibwV2dJg65lVSF9claCE23mk26SU
rUkrJd9GRya569RS83CxLzJDm6e7nkU6IwHoH685U5S5AqRAwUj7xnSy0LRHcVTn
++dSIvii0Mbj8LCltlCncDYQYaw5r/nWq/Pds5GtCvKh4QmQbZPfRN90T//t7faL
RkG1e+ShVX14EvHHPQmi5t2fCvR64j+7BnGsokjH7CiO6I/+FzdhCJ4Czwf1h0VP
Kr+At0yjpRlr0rVpG/YlcLlQzc9AEPk4AuRxOc9rmGK7X8GwugCK72u6uwDGLXLZ
nGpB/0mfp3G0iQTDqefUIw7tvj+9K8LnSS0MvSk69x+E9A4SSaTk+ByUdd+t421a
J0+SB9NH8DDiHnCyILH5Edk8A+cSZC+M0HIpBB6+HKMkIaIRHJng0WX/v/8fxU4s
DvrMk0cR1RoeMYgDfW6P1DHVIItED5skSKzDi2hy/j60OMijJKpgd+ooVqQWYEVj
L7Xnbh7qPsEHFqi7942NJOCKCLjSECdd+DFvpj6F3vPJPZ+xoa5PM3fBA7Xvuyx2
bImvGe8ctRD1iMrxYJ5xH71f6rdMy9SyUqR+tEph1etz0s5nwZco0QChh2j3LYBb
j9suiN36t/4xJn6HTcG88Xnb+gZTvvYgDDyPMNVT5ti2ABB5fYL+Vy1VWps5Smfn
Pzx+ux074VctVbnI6z2vPfTn3SDLqwIl6QVdTC9kXDTcS1FTVzQEQUi+yC30vZo5
RS2oWyTZPTWm5Yx1MZyxjSiQe+mLVzigzNZJ5AuQn/OrwwR8eQUqvL7uQyuqrB+s
s0kbPHasvxxz5P/LBfyjyg9fdqqT0LxmyZEDMRH1Zz+iuuGRFSf/1Fz8+CHZ0jVF
tHWm+lgsH3rQBbIlUZQfoy/gNpSlM2ocgRsyNcj2yFtElUXoLs4M4hGjoivsiyb7
VN6WS5D4TmEiY7IoVZh0TCuEPdR0zGpxgIF6Fl4uD4fzkObwFSzDuajg4amg27Wi
FmZOtnHSvTip9ChHtJgb789RE8yqW1UrVyTod9FI6mvMSGlIZgIBmuU3g4Jx5IZA
O406BisJ0j7l5SrrGggPOsgQqE1d5LQJRTIc4/+a4HvrOQ9vEX5UecuP3rsSRZDf
+/0nfhLhXS7yFf4ZdPbg3GqLkMf8RUaWF/rPdz51HdOVVA+DXdFOgUKS0Bq/Fm+I
FeiiapgUXloHKfwIVTIQopRALelVBot0hijB31QtySUrnuoudskSp5SO8clijFC0
A85hdP/HCeGQ1AjxFNtUxHq4UuZKuEWbNisQ9vJ1klO3XGwqXVwNc1ofRzmGAH1A
ZcUj1mIs8cokJaYbHsfPuED/3PbTphYKOoQQfpBZIt6byb4Lv7DcEq+m0SVseEE3
s7XvfAeRY0qCgVD8jE/Ydbh0udVhuI27oaddRCjapszwMIFxosGaDopzoqon6tfX
1h342VvELAA3vz3IjaQaLZRZUrfkBDydiiNyYJakSy7+TvXob4BN3zPE1fPjqQb5
lLH9qcsPhgFf+mutjY74WYW5W6ZaPwyrmS/JDDEFZRBQdTlEiG8EJZXH3YRLHT3O
UauGXXokWqu8u3sZ/MW2UZQa62zn71HOJJVnXLsAPByd5IlWYRpAm8t0s2HLGVlI
RtaGFKr0O6OMrH4Fk6ggAKBajxqVAy37VP+nqq0cxCahRscmOIWL1PMc9GUoey1H
YloUgK/mk4bVzh79snUwzjqEPHgfdklYCa5Ofe9/gAgK7wYcS7NNJVRChcuSwBXH
3s6HPQM0MRrocF3craOEiHwzQteZoO7+2mHfTGCAs6xTTlfs0mGnMqHgW3XhzTfM
pl/CY5HtmJAcT2oJxoww4xZojjqFJR4koRDN3tLHjOZHABIY9m+PIOpTRYbFdDlt
aXN3s1Pm/83XZWWiDTv4CmbJkz832Y7y5SOnbOtdDjSul2/u26wZvlapRk1S4oEo
UYvqIS2VfnZSVE5i1hskkh8zdUuI0Fdg+6wLWo5g8WTofSsOwJfdaSx8W6Hlteld
N57Xa4TQHdxiPWhbUokHxuwnOCZQvah7ZeoiVBFgCZlzwNlyIrs9ax8gBpDHLnT5
RQdIcQeoB9llXlvgnVnR+Zi2q1YpNTXnflsDyUAht5srwvQOkkDnCNKuDjFawxbe
gvIg6RqjekAL2wHLMcllSBgXup/mfL9V5c6IvjL+y2lzahF/6qoQCiSA9qZX6xXr
cHljKNdqwsXjBAEn8f+eA5ts+bxXnYRjnCuMuPeF3UitTZm92ghMVKQSsNwUVmzw
N4ginHY2b6yAQjq+//L+O3NtOFJlMq41K34bA4fE5Rbs4mhX6XyJBn0i35z1O0wc
UQJUbmpH0a5jIkWFcE4hGvXCYKJgdsbNc2GtT6nqTgQAPxVpZVUd0L48XXn9Xrtv
tAEEZlMo6qRyyl1+NoDAQxJ/EAgEEjnpfz7xhcOcxz/tWObKK68s5pFwNpib/9AA
Q86Vs+hk9EZ7FfGkyJG4UaOKjRoaD/alz5aMm2Z3uOOU9eKpJUFZZESvuvGUAXRj
G7pwrBhbAvBWO+ZiIjNInphWKQtUSCwez2pIvPhLGy2Bk/BSZC1C8pMTduXBCD5U
/hggdlhT7pwEG0Ez040TiwcS1wEEEmilhuNwXtSbh7fVNjlUhjXjsp7GhDqWymUw
nj77C0c28KI5LUMvHkDl3P8/s29vKK215qWq27DIR2Bq/xyOly+B8XkEmW6di9IE
6DcOjzoZ771yWJrLj7qO5rndxN2hPlAXfej2VvGiPiQBhExo4Au1G601jO+4eR24
hC8SgwOqLBKXzYNIsEnNG44en4SaPJ/tT7+gAa/qkftVRF3djHCgTtC67x4J0tMD
5qdNzlOKcQjU5ICXb1StfGQHqVUfYF7u7L8iqfQ24MNZ4gFc00X8K+2V7KXOasa5
rR15bwHRZplCwRXctHPAjetwmOLhsZFak/5Gfniy3MbPen7PVgTZx62X1LT34UJ+
Zcr6yeY7HstYRWYnBHq1HYDlqLHZ8elSYaYXwzFniDnJNM/EKLqQVtbCdk0nbknv
DmD2q5VRjBpgtOd+fQ25LLhTuG++u7qMKikspsFIfFp2M4yPcee62D7TDtJODpGS
5lNgRRkakde8ItCNEEIdbjjin6pb5q6vXL3VE/Z5Jmie8QkwQi1KXaFUqLlZuzoa
F+oSoJmrlEU06YUm1cwpShYaL0qrCmM2UdQ6HMM89FgxINgEzIPd1tHu1GfOWi5t
oYCXUrcvahKuKSFh/dfm8moLv51WmJS56LYDl4DBsjC3TeSxgcequpzDqp58RIky
89yPS2jTiBzJNWXHuqgFqLDTKva8eFDGsi8Jv1EZg1Ng6NUVLhnOm9IyewK6gGK9
nQoMBC9WUVnim+EwXe73xEnWRTbFGa8E3+NGHpoLgqggdutPYhuyD0iL4sJSc1hX
qkS/IqEcyKbNT/8FPPfSwA4OD00DyzTKXAoF4pcvMsZkdmYi8Uy244Z5KmUO/elA
mzHgd9BXOOjRiistf6/wFlLjf7ad+o+tIBJArvnU9gmwqxuE2BMpydE/VxkIEyAV
xQpfE6bYUpaHH0gJpZ8AM5zxO2WEiyYwbqnD9dOrRCF3v2CQdxb95I9/Wb0iMW5p
3YBFOSGK/YiDgyq7FKHnhvPQuB9GUK8JTf6cAGqwzm7Kp8S7xh6THtbNGwmh/7aF
0RJnJ7KiXr17gnFX6wnpIo6amgmSu1lZsvTdAWSGqCdMOgD0bRMXehfLNMbkS3jG
wJWzlQmaWwdG2txJw+sVj2THsQm6pBFDR7lurGe2I9NqmqYW6eKtqDQ1yOnmEV4R
FmeAxGzkAogFfbeVMXqcmyYX5u9scotcmPqDHancyZAhQfH23Ofi2bRBtbkaVN6Y
bnt68PU60YrdtyCJLdzXKJrv0hCPPFVB4kdFVXZbHFdGfA+zNPklhsaNj/a5iP84
gPJdfKoeZyo/He21sxVBiTzU5zWg57Y7ak7UW0IPXwkGo6Wf080ycl3AgKJtdcJ/
gtnrT4GH8p5HqqYvgvOBhBEe3v6G6HKPHRkkk1sxzy4b8hlUNWhU6X6Gh3E7UUKR
MVF3/aDFCHFFNKBgfcFjfNWmOqofG9woTWwIf3BFlu0pm4GrggizoqH7lz1gwXOK
ikLjn3n2+GxNz4l2ErfXbS1oBGqqWu0cuBwu7PgCYsh78X2Z29zuu9CcSP7ZQEPm
6Hb7+T5AXwFolFTdLJY4vDgnsxYL75AQJxsoy3kzhKveKr+R6BmjiCCNv1m9TwHA
W9ChiCfb34vzbn9/VOdR+HlHjySHItK134zV0AXTiv5M5TL1vZ1Tgp45pFFze1Pm
8PsLhRXpT248frCnzkOT25ogcYZS0Bb0Ufe2iMvFoeCBojTU/KLApF+XVdfDhqQj
i4x57Zi0lHbqwjX7G3zuYZ7fGEqU/Pk+XfQny19XlgmfjMjptTr6anp2xn+UqEzQ
hc1HRqOj9mdfrnT4gUHmJxp65XklqHaK/eBZXYzKBrLyp12GUJ1XWF+SjtAkhB5+
raKMo+T4liIV5J2/8oADAeVOjo52gmkbPBA7M/Fy+P2iXcqIZ8KBY0Pnjo+lGfyv
WUEidStlgm20W8CTtK1C9A3ahuy/jeLqoH5VE6H2OnkGcqGPd5PUFw5fElrv/+PE
Td4C8UIjFjL2XGxrkseLHEtJiREptu5vSoK93QsdG6Ki8gRGDFmtweiCjBXe2OAD
/KZjcDkkQy+G/yvuyxs/n2KRtUFA3EAIqhwwkeWjQwFQG3Lj1jGbrbUbcaxeopVm
Vgs0SVXbg02I10z+x0jRedUy/vZnKhr+I3Lby8yzRFDIKPhB1k5yFasPsAoPIl8r
s74S6RUBrRZK0TRPLS8cFudNAxNivpk3cLPyvaFsbb7Qh9ALerQdqJSJAmBvJBpf
L/gAOLw9cjkcfIWp1vTBUCbnX4pvs2G+SAJn2tFdTX4zattl039flIf4Xg0+zZwz
O4SkbBer9E5Ty5GVW8PRk+k228OWwUUpdVcSzdNrU75e8IGA3PnhIaQ+Y3dKbAO1
oANfUFbUiTeEpJxwPqu3Awkopv9jTfjqf9gvmzL6GsBjzUSPMeA9yIDohUVGN/ys
Ig2mUCO3+5DNO+8riubJGRaq/jRQVxXa+OQdly6gC//DimNsxfNKIKNECbvsoTED
D5e1s/Sh4V+KVCGcCkUftg==
`pragma protect end_protected
