// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:44 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KGg+e37YogGlBMy0JeoxGfRJaiwgEXkcZ0Y1zXcLZX5pJykHHdgGnAIXeiWPFoTc
J2AewfHII0HHYmE2vuY3uw/WY/qi+H/DJIVADCgt/fp0UlULkQBtJatBOYIbv2Ns
0a+Q8qIgpnCQApCNDlUM/VXfBj9vulJbPBh6xtsjfeM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7952)
0irt8Q7X+blBXaw1IYXldjO4xMsjEeWAqH8vpHAECFaH7+y2epnphirJOWckBgNq
ONIipMelTZ6xx8uG52dfnbhKc6yIDjpzMJZzBTIrZVeDBldQvYvHhXSqTzYEIDSg
cYy1TYbXx8UZlMsfy+R8/LwTWWapVopwMwkmcJQL118RWqmaZegRLW+Rablg95Pa
3Q+FSNbkHEduBcZl+yhwit+nJYKUrkLLZC6q/qpgGMV4aGsaUTTmqfDeBK2x9dRu
PD0S9gZAUWY0riDB2XPC4SPX+nRLVb7s+Vyhs3/JgdpGspNh0MxG9F92xCBP7uQ1
PYGhl/Llgw9KKIFiDUNWcenCaDBmuxYvJAKmLL5HSgJMyOSfMOcdr+9cHZu9ZIOR
g7pIKaJGOOFCZpN4RVxi1CGw1eLMhUyd6vfu19rN0DlP8iheu9cUm5DqyG3XFdG/
CtM5/JOnQs43RKM59+MyW27f5EHAoGKYVHpMNTmXsQkB/UN0NQSaG2pyg0MJdl/h
O3NqEmWk4krwJvZLbpA0jClX/xmMsxSFxb7uvX8jL98vVEOYnNf09tpAEZa5e1Zx
odYacexvmo/qFmBvLR6BVqdn2x5WR6qCQcE5XjfRDMv3MWcu6sk0UqP5/0Dhzqks
ZbwNm++QyV6fw5fuK4Mh24OMJlynn9Zezy6kv7wUnLO4X4VKZSdQc5U4ZUodOcXg
0LlxrY6pywKGB/j46QXaHtMuMiZN0PCPND3qx2/iZuZlWqEDIlYekS1NFkz8Eb6b
O8RVbwGs9a61kpJGvrLQZZokUudnDagFSUHep/hrnkSktMkbdbsMu2SXFfzFLaFZ
3uW4F31SRdeHERu0sAn0Z3dZ5Yc7g0+Hpx8RBUDca+tVEi/W6EeA3pElVUPGKPcO
j1WujZJyUuMMk1lJR8JMUrCIuZV3pzIqiKayKew+vumBLI7DEK7Xcj4zYDrP0kar
IoNRHw3TQcanMwsSQ2ckzIq6rk12LvIgiQOWiWefK2D7Mpe0nVZNO6sVxBCFG9kc
uL7Bx0QyLMUoY7LDiDQdAEAt2QAhPehs3Wk9kt7e5l1Op4q66d3AF38w8E9zc9px
nVLQoxpgpBtQSTrWScO3J90lymtTEiLevfHDRMotZ3bw9R72NLqh/bw2cJrbzle4
CkoG8JWDX+zWuxC7UI+c6ILsZE1zvQpoLdhV9BEKXrYLpfyeeeo0oQbbwh+9i2Qj
8BpUppJn8F5wdw1jSjtN8fidFgz7yX5Pym8NFaRZonXXAoWZa6/ga98zkCToxDRe
EqTou9OKQyok1QtZf5Uq/9HaYW6z8XDP+AoxUXK/l5pPtm3hna8rPeqFu/VPJMYy
U6LRy4B81vBKVaSiLkQ10rD1VXAnR/0DIQDL5CLFL+cZLe83Pjdv/su3uFq2lmCN
crzEy/BSsnhnTqBb2wTMTBlDIqlYvZb0ZZM4Rd7+ZJlD1Fry29eyyPazwWJxk3bV
pzy2x+7V16DRVw1Qno9ohV6FrkHomTkOJCrHjoDIstBR2zdHS+/KnFDqarwiQCDa
Sip4R3JtlTFpTP1T+0l9D1Ipi6z4q120wDaahGhN3I0EBYZ+ZVuAuMvVw9UqKiDu
HNzGGLLOu+Ha2lWBXvTRTqV46jsiwlcLbGazIxHddjS8iPDae020BkhiCKB0/NaR
uqYfp5eDQvWuvFShukeoaseZIMZ22/Bc8GQnT2Pzq/uiTwe2RyowRDhB2H8/bl3P
j1Fiz8di/o8B7OK+Fo+3WHqGnCZKySKO2bO9frSzZLQ2rd2LmtT33i/92Y21MZiN
flt9GqHMCEdNFeVi2bK8NLVY35esiLB/lmc+p7tTvZb31RmYVb+qIJY8yS79bch3
sUWaTeXvNr0FikXdMYWAC48/zi1wUslpZmPO1EufBSvw5jlFwUDTjT/tpPScckr6
RgdSeRUKYuJg/8biOv827kR6C03/JC2z1q4B5jVrmy3D+n1WeYlFg7ctIN/dlhFh
zdxDmuy1bGtWE7aNBPNi2XDMoBbIpqs3nd+P+1pGUpX48GiZmxfoqH3AeO2XVGzU
wr0hxHNNEL01oBKH9UXzA+q5Ni9dDmpyA7YC/phE9hC2ooF66sfB4B2gudw5q+eF
kPq6XaD+dJbBF4anTenTTRX0sXxlBsLIyXytKeHLJjeDNFx9XOYB3TqIlMKXsqqz
vRSTArs+VRlnwUXsnn09J8JM0Vm2Sc486WvlueI16EmzhA/2/mcjxtTM87kSf0G6
1CZ35pc+fOkh+tM59nNBVCzOJ9kQkuCSc6CV+j92CDHkIsK+82HBolw35uMTYIVH
7UcAEcvmS+16N+di3+UJa4liw5O8mkCLyeAgXCsieS9O+Qr2m5oHZIrwFP9xCCT/
hZkC0+GTkl4CyJoSEsgPkPAoh0lubcHAC4qQjnco1cAuV1FSI9k0l1RlARk18VEM
fULebIN4glRRFk9BtwOxHn9EnRRse7CtmyNlu61tZt4ptLpIgwVvHqnxxcEK0ckl
Dkl+sAn1pNBztHou5aI6doiEeqNuwwHhgYE86u2eHbZ8gnwwxPdhf3lxjhfmy9hC
mn3srk+tjJa6aeDquGj5isBFoC9ZpOfeil0HaE9kJ7W9L/GU+0nVIvFDTiambJIC
d8uhyeAJFq1lal0EAZJ1JlBVu1tYM5vfzzS+orPSmzitUpUd6+hw9TSRZlpZfgFX
6M9MWICosKmyoGKjqOXom1bBwi0HmJGVaiTsEopD8d74uGx1O2SSNx1OknNdoi2i
6tDkfj7fqdPIspbdGOSAi2sfo1GdMvmPfTSSqmIwwRz+a4ytnnmBmtbOeSlXz4Wz
xixdSsWA7+h92CvRtOX4KSMoxl3PeSBfN6fSYwvNzsSB8T90tRlbW0cRwCDmHg/K
MUqvFXy14HxVnq1V3TvWriFw8KUJ3IqlJgahrOKTYj739ziIok6cAKb4138lSojX
9dleBiLrhAutzd0e8xtVPZ1DlCsQzbBGjX3zIaL1sybyRH6e80Up1jd/EHvF1taE
BVnSKHxcK9jxi0V1uCwz1Pgfuvyp7/D+Ji7OIhAWcXlognkTDIuRGiK9mRX+6p35
eNey0WD+vBiZeACglTESQtLHTjmRGQ6ygzsuGCwF1K/auAJLghYhoCU14Exg2i4r
lD6nLOXta+FjdFpAk/7FPeS51crq/VuAyaQzggRP+rHyQPUQ5iy627btu1KwDFrw
pOv3Bq67Sp/jZdMQZpucmqzSiEyqNliS4ScsfGeOG3Y83Zi69Rjv1wiITZYfvV6X
elq5VCGMD7v8kIX1b9GEPGGTev5cqRZ1OkFZc2qCuYs445jG4gbH4UnNZKs1rSpx
UYBTdLeVV9nN95nkKbaQouGSgKavnmL7hIs8LgIzzBWfAXPN74kTjccbYw2jXWDI
E+VbfgjC+n/NTVrk4cUK6okRU4+oXt1midaBWOC0gr6lM5BIVZ1VhD+hUgJwyx8B
YljBARiQvnRM/86e5gnolXqVBpdHOI1a+tanu+kqUM1B3h9ma043LXALMo00SMG9
z/eNLFERfURcXad9T9g3jo5Gn6WRX+fXVGTFfwIOOpL1UH424gWqaVFdvvkm/Nfh
iFC0HTDdoRQsppKVYDhr0S1/XRQGXYDLlbBcqyQUy38Sikhm9XS2l/Im8ZsXx5cs
Jhx2HvHRHd2TPOPVIZyHT5tRWMHbTaZKVsQkUwnU/Vi9q9a11T2IzfGkQ10EMkpf
UyYQmcvLEhwPypFvIWG1x2V85nfAMuMwZFYmIjYUQIkiQjgmz7fafzmto+7w2KZK
S7IES7OecYkX5S9i+2Qy3lG6wKWcxBggwRcSxPtgMekoG7Slv8bRe5kY9prfN0FQ
NlcMOaEFGVr2HPOczRFlWEbHdnhn5tvDiJaUWOW51OJdjTxzwJsUWA4QEOYmnBbx
2skKXz7WcUYU7j5ZBznsWVM4J9arMaOW4lun0vDkpAR3e5CKYqdAdXd+SDidW0u/
qNpV4lo7BTCrJ73hKgGfI90l0NI+fAGc6njDv5YGLqIDy8rO/od5nwKDTRT0f7A6
owWQzijCOA565s4e7fdCxdID5qChC/glhmCignUhcqP1Fy/k5MM+J1M6AWPSu20y
zZzzbcBmsC0DMvtt1ua9e+5SS7jamPLX0F+RtNgcXht8nnKQfU8n8vli7oFSSAh7
dlzURoj4azhD5cxMw64W89xhod3FKzqgo8FrLH9pGcE1LSHEgLVR2+NJdXy7Y3bY
WoaIkWnnAqryzkLhRmGR5mILfJZHMB8r2ZcmkVKcDcbTsR9zqUPRxYsw/7f15l2T
f/ezXHRlh7HSxfHUCUBFzN055VHcjabwrea6Uqk9he57cNF2AHUGipl4pKL+xJaE
L3s+3aTDfYY9bu73C3syt1zT/J0gdpxYVhcXzmlAL4Fjn5f771limmW5n+V5HuYf
YXNX/WH/78L3LGblDFnBa/2cIbN7zLuKN6FNpuzLw2klUdU1xzxgks6VLd/FU0Q4
bivh1nqWJHMAULOleEMmDBQaYKCO/htGpS7patJdkiMRCUIE0On5LrIZ+Hwz5TXy
prUlX+VEVFwjwC4moPYYOFl2UVQ1pknRbGIa/rwaJqseX3BQYRNUBnflMngtTpf9
JaSMFcxOiCR+rr7TPD6Cx3VLCeqMofOQhZQddwnogXOpizmEwRRsQRns0QzNmvGe
ZDU7dmaa0JCVRFsYHYg5o1QllOGtv7irQnOKQYN5a9WQ4jWkqyAkeHqt3IfCxuIP
EnOGIgXEBET50EayhE51ZASVJr3rirH5LvxunYHwZOiNuKwT9FtVPjsYCF/gk2jm
mKi6NlXkPRppfFSFKWORJdUtMiInSvgmgkA26xhBJ4rSQ+xyZib5JcSsPaotawBB
wJJIEbNeQsw6Mu+xsjSsBvJTNgNKytmSyK5ZucdaGfK8Owi91afT5OezG2Uzqwp4
Xw+urrehkRCIEJ+tpXvLVCkSS0pXpvd/Qh9lMNxjPtV+r/fe50eCxzGDoZcbjzQu
NBfQDzstyXumD33Xvinskb7ODVuE6v7I/gY9EkQxjAdsPbY96onQUSCKUXmc2eZP
ajlMheCEgm3/MwkioU/dojKOO30DXyjZKulzKkqmD3kwwznOtAoJZvZG29tHuvf1
3OhU2e+YaK5nN/7lW3D4lxhjxOZb78/7p13cI9FkfqpJIWg+Zu2Loxt7RQMlmtZV
LDXyD8lN1rnppUMpQ63CeX5xOhZkTNSsADUckxI37Qb3AWcfDZZI91Ez5Ht1w62c
OBU51jlqOsUH1q6p3oLJC/LYlUtwgFa6PtKfjZyq9DlHD0KwQR310/UfJFZgX3ef
SLLw6bHqvcrGESJl7n2/+sOc3lzBJ7Ah4Num+HpeHTObjeDuNz2BaUStpAEYwEWp
cxy+zKPn1vysCSz3bxK2beHKDTulTNlapc5zUD9LRczqX7bC5jtXbOw5Z8ALPyy5
Xd53J8rEqe0U0d61rwYLvceasXz/ROY4w/TUNZ6n8EqNmgoMdmZhkvWiXaEUak9p
0RPmpGli2SGo/g2l8v3k+c9qsZtYr1s6l3zux9JjVSbaDXgClTIIaspS59JL4H9Y
Iymt6/2mYjDiILfbCTBZha0H+O8El9mcWBi1WZXr/yFF+6lQoSAFoh9Iv9k1TKbi
FeUFIOe0dVsvbxu9GMKg/WvI00vqXAL91TWGmnnQ2aVR1NPtzBI2r3jBBK6TJNfL
oKm/6KlSEIASii+A71udzlcGvh51Ie3wMpU2PEFAswN7Vu9aB37TTLHAePkkHODG
Gz1a4PEAQUJiCjwOOWA33gzAkbIKzcZLEYirHifzlX7mgkT4KZhI4lXt3hM1EBbt
SDYDcLkTRT0Ud2X7M9zd0m2gm1RtOJjxgx4NdfjKhtJ4oU05S8nMu2Ufn5+5Alzl
G29rJoeA8Vi19FDm94P4AbzRMRT4zqSIO5bY81rnnAp1zYxPY9KimB+EYGCN8qa6
oGKJwYCz/M13wJued5kmGyIWUBntCEjLM+P/aDp0ZBqsOLHo9goSN9Z1vDip+rsD
0YknsRNqj5rEYdH/m1WesFg4jcxicQc1wv39yo6qq5HdO7IQFDDwK/3cvO/iMEIi
sL2kWXerhna3dvu5kc+a6wLdM51nMu5pmIxaK/gOI3gsbPOLF6taD8njnbZ42Unb
U6sPPIF5l7OpCQwn5hq/cKRBpcUyTdrVcSoe7j4bkxy2J5XewMRM9m60TQS2dNgd
OXMAwSCzr7eZ8Ak/0zEBDUeud1SGHkdylqGBpDNvTYp19/SfJ0ccJA2FlPrNbyaT
dDOIF6lS4XbBqPTmQ1SCEaknrDxlNQ2QqQuW8eccaN6MvC0yOrIJWw3DvlHXCCiJ
jW4pZcUdTGROuRONPyLcUlZvpBxPYNcpuI/wVg+3uOMixHNYAWRBA6sfHziQrGg9
If7yrkeR9uiOqKEBtA9vu7c7XPNrpySpam8qhR7qMlthW1gCQdXtY4JbYrrrTOfy
d2mceUqIhCNZESdn9QRgZmrMlhaAme6WJ7TlPYmd88CGABTHMFQbOxkyN02Ik24A
UhFNrz2SZ30RrrabrbdFdJEb/+cnZxIRFjQo2Hl0RI4MZjdygP7JY3SVmR5D8B9z
tO2jWYEphRAs6EwchsrHJ3YiaLK0gk94YRLFBY2OddUzy4Jnx1N/JqeKv1YGYsHJ
SnWDZWZOhdQzYvMLz927MGmnKzvyxYY61iFPu0B7bVBQ1Ql2Yz2qFAKuhDh7FL3S
YPMWzncHyWx5yCO2s4PpHiuXki3a5u6kf/3T+bHcqWddjdXKoLBSntgCjgxJ5GsJ
vVzTUP295NdRt+5ZicXsIAJJaxzfTLKcYZGdDIe+3seFWX9RY+erW6nr5oOpYtQt
1if87m5Gu+gXmo+A/o8Xa6B9lD4JkYbFz/9FQHQI6pz8sT2XPs34XE7ptcXB8/Ic
dyJfutb4d9kK+jjhsqlps8LNhGxGievlBNHCnYTP5LC4/LtuW9qly/Iin7pWrX9E
F71d5ZSWaM97X7fkKUS6yvpV14w5ceEbPo+mOVmP4Bh63WeDpOebOQgpKtuc9P3G
Rpkj2k48k7BnJUlnu7iIQqjsbQbp/CRyBydG1pBhnk4613jEX5/7KASreYpVEAxd
5UOXPASMNjPf7klcOa2hnYjIueFoByA95wEWc6CuT1w3HzNw3imz3dojjnCB8ANu
4XQj0mEHvaoCgi4XVZ6Rk9/fGBT+4SstDcCdwDq6q/6WuMQN//fBD+WMw8UrjU0+
lKL6BnUgWr7CqkXs1NAaiq3TC1uGFPLRINws37ojWVfrhKOZH8qk6vmuYCRkHl5I
Q0+Wc9+hfRgC7l9Z/Oz784tHUtf8PPQHQOD6iuttdc1aFZS5Lw0eNo3jLN5w6rj/
TNIEzUE1D37lLBvWpGHkFUu92+TXsmGBFHQBCFMVrFAfUwJUrrgvNk5O9jTpXttH
E6exyfzrNkkYT2N6c2Yfd/Y3kPtFWYZonhur216HK2tTdM1Im/3d8kA5237cgoJg
In9cVMdm3RH5mrHQzVwrhNtWkRk1eWnvcH7dYA/1/2VAUpOeFZ8Iy9XG0m5SQWT2
ljQKB2ZLSrQ+SskssrO8tG6ZGNudDvohUwpF+SGfIwfHNYG1SoTXZrHYBtdQa38W
lNAjdMzB1lQlQkrEzOWsJMZaHjl2pfkyIlcdQ/MVxKkr33itRa/o7ZjzgeAsuDYB
E+R2JspQq9DRFk++XovHoEhbfs5WuLWkpnmWDM1F3AWF6HqhlRXeOnRTWG3IcdV7
kjJzkmuchJZTlAGUqXIELtG5uJuls11G1Lu2mFMyQo0AKCltSvhjLQdtDcxiMFv1
wDMm/H308SntaiJGKDkxClEy1w8xirabdcllkHfZ5aYwer4ERLqsqbT1YvJ24wdA
+DLBJL+7rwGByOALf8JOh4w5i5VBGIaBr4Wk9xq52Hg+SYWFCDtC2ffIEiOuRjKf
NtqWV4TO4QSCHpeyVYw+S00MNf1fFGFMZtbkJ93W3F5nDHUM+o5scGpENpl/GYcV
wx9KcCsQwo9R/h9Mi3OAiijXzgxetoqMeO07zhJsAbvhb6L2KcJtR4VXBZcxacFd
Rq0v3aUleSVgDIsC9t1NJDLjcgw3x+Wz/P/kS9T1VUzBa8rPs9bS95tbx2rZbwWX
L70wKDhCy2Rs9s8/65T+sHvVcBDZyToUTZ5LMXjTp7DCvBJHigk/Rgi6vUPrc2S/
6jW2iBHWKmGJQ1yxTL65+x0ohuzWuGWXOSAL48AnZwvvhFWipMsk3GnAM2uLucti
yeg/Rre4rimSA03NqI+iBYskJ58WaDPeyt56bhcdV7npnYgqZwmUbdGlOP+Hhff/
QEXFSvjF8k7bX1XqTrFkFhE3NuQJraAEd140G95OxoqaO2f+XCxvGEbVwH7UhPrG
UBj/YsnJpjJ3Euf3htLYmrVQlq6HrN4m6JNTPhZaK46rTZyItzrd17ha+gwfczHB
6sZwiYZWHbZMgsduYQ1grv6kCOlbYFtdQbQA7s/UVYSwIPl4B+6zVW4ZBLlFma8a
0Z1Y4mGHAgl9XjjtlNFwxUbT98Eg54HnZ3EiEb86DSdTkEMG7rfmKY5rfTz6pJEd
/Ivi284bWjDwtJa5sNp9cpifZyMjgaI1v2zJ1f9wNHDRsui80x29zY9skAVx4YLp
z2/WyQksRX4CMhh5pZWOf1vL4QCM8kAoJiqXzJJLsVZBW2kZNlDZQXn6xMcN7InZ
NboMCG/rw5BgRn6fbKiZwlpbq56++buM/sMsYiGAHzPFKRiAXIR75txNN2DPOpVZ
NyW4NEfNastC+yO7FWn7le0fgnBq2qWuLaDmSsc8Scn5rMiyrzY3sheX/1S5fCEt
7QRFIO8SvxhFvb/Q241WO960KPiAXL0lfX08NNoiqQYOIWaHrS8Eu0Yz1oyjusS1
YhfiVtLwE98EB+s/G7/DUZPk4k6haMUR2DvVYbjb8w0CtJmY0Lh3VD8l5GINIROK
QomevDhclWQUcXrvClTO5vZlNnszFQHHZ1Ndnu0+qrqyBCmUp9aU5R9HBk/Qkdkj
dYJ9grEaKeU02UeDG+qPfSG7Aa4A22PKvNOs2jYfsI5/Iq1vLMiYEAdde68mPBXj
/Uj+NxItkw/AaJphxsUtwimyWfDcTPQIGzlKvmjuVZMmRlIS2YtjihpsWfc/i39a
ZKlVvDnr0Kvb7FdMA9bkIYw2tr4m5LaHDRrTxCMv5oLcUuyepdyKMk2iLpxEyF7S
BBq0e4rwZYz8HbjHYC1ICKr+00Kg5Eqx8Jepbmt2RiUUkGblNUyo1jG/TX++8x2X
HAVxLP7hjdBzbohP10NEr9iMmTbUEQEf8SDh8mU1ejEzqvQ7TPsc+QBvpGdgj8sw
9f/TqRaDhtOokaGJpqbi6MoLUh5xhiAmEEO2jtWBVaJ4DrJVdWEknyPms7UyHW/y
H9FGoIOxxujOBEj4wCItrtmVt7NtwKOiIgCYVarbJmVW7IEBdHRXqwDGOQVVOnyh
74whUDch/Zc6vL69dAhUvMlcOKSu9zvYHp30rAhqvW6/Cz0QQNl/bm7JYJuzzFFs
NGJez5036sY3BEaav2HTWlhi3zx/rCjYBo6MOu0JN7UTC9WN+H1nR+F8rckBuyfD
EzuGp1kLsfzcZlXw9EYHXKImh9k62ANiNk1GtDkCtJeoYHmeV5tkqv/oRE9vX1JG
w14zpsznOwLfPMSWu718Q5Ee19+bfgNtoMJrMszXMdlGxmz6lWGdtziTlwnaXb5H
yushtsfd/v5zqWLZdD2neSQbJriR9/G/rFQWXw1QFI0USfEWIkagvSQntqD6Utdp
qaldJE1fr35PbN0AMi7FbFlSfaX2KhiOiiNfRXWpC1vX386DOvGZKtwPcp5ZD0gB
jZjyTNxnBHOmpimEyorknHKqJJqaPHRLRi2A+KS+9w/Yl+LwI00anOeZtgvToDak
QWBakOk1e5uQ5iIGkXdwzJh1tVFYnSBm6SnCOWmjiUziAZU9Cpxhw2pdQBe9oNm7
Ab2AQ7WUaxRy7zlgj1kNodfZttGKlo4NkjP0N2rOgitT0znG2nLt+tiQ2zplmA+n
qj07mwce4a8zmjVPJz5Q2LYQLbqJ5pI3YQdPA2inoQGut7HEZqcz/93lr3sNtJPr
Qevyrr47jmtBU3XPvsYQde+jbDyFfmou469GJXt6fpgFJ+jnE0+uMvHkWpIy/DuG
c7j+uTY84pcGk5i8RT/zF5ir02sYx1M3LoeA8RVjaNTU8FCkhazsWGAKPWCJJIv/
5lL8uMSgMBUfmy8Afo0sYogP2DjZHPAAU2e474A1qvjCPith0LMInLEQrwHgiLaw
3Z6MNSVkK70BRXPXatf+PQvtDgYQqx8SXRrrNzOCB3vBerSKFlKJhII04QuDY61D
mtPC8BJ8gAt2O64AkrhU73yIomvjpnQbhqdaeldKcQE8TP/N1wrOBW1IRRysyqYf
7Km3RzNoG19kKJvmb3eIKVKq/eXEY9+oXhsLdJ19luTFH5jYcmHAy/Pa8ivdr29f
qahCqp6Ds4w8YsLjQFW1vSV9z8NYK+Ip1DdDcaN7b62UJocplD6xp3HtHeggujHa
WqdMHA085Zy3fFmjsEfKIhZNz3V5xvhdIiUb3cgxnEc=
`pragma protect end_protected
