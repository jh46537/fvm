// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:38:01 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wn5GDjcvY0rrTm1Co4DdDQWop5INVbI5iNsr93UZsz6+8QYkpyOS8Y4WLvO5L3Zl
nqXUW5hwwwKIKKMHbr9aIDg+y9diHP5GaOpd9dQwvOcarOgTG28TLmh18XxKB6Ly
Fe0ln/pF8mqbcXhJtKUhUSGdv7a5VawS2ttpfm6DXDQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6832)
Pk58M05jhpADJDzy60Nv67fBjIucixvw24cF0zlTsQ4w8eNmFvhwtRJprj9THQUG
4V4dyWr89ZAH4UjrP6guovnhx4LkOSeQnk4ZDJ/B9w4nKaozY6XhsTUi8jy+u3zp
afbllKhFgfMMyt4/XrhXG13xutTpOB/01Zrxn9QhGkqR9if7POYtGMceWy/j14/h
ABjyFtb/gCVaCTt3Vm3HTL6/UKDIr2rw8O6UzN4lfNh3xjbSXjl311tawVEjsizY
vrbqbnPKIizerc+8cvsX8aPeYdr6PIFJbOUzOl+XogXcefpz4WNayBQ5gFtdpLyQ
UDTiSKyqQMGQuudp+9uAUsHR92EIbrkFKe6GvtET5iY/laBnBsChjkiMOr9h2H83
IlpjyAKus6zy8sDh5Mb853/kImgqbhbH14swxTMngxMuSaXzIRxZqlO3qxfcJlqQ
wVLH67Upj27Yt49glowULJhfUtFH+i7dJ6wfTu3gilKroLhX//xF+GvRk+qkd+Nw
0JYPjxJ2ahbsPAkM1a+tdMnLLQJ0H96kDgD9obHbMfYjnTQtllLB/VrFrzntNLn9
x8UgQ9lMb1dCYAYdPNKSoUKPgI8SBvi5+M1k0Mh+/BmIH+eLnaTxPMzcs9Dlnu26
7+7Vwu9zyvTgxYUk59mjmCBoBlJN11JS7egAuzuibhb34J0gGIFHfdshHkszF4mz
8K2r9o0ueALGg01XZ08cTitacCg+QaQbPjL8xmH7k/WGgB9zpL++vlFibGUQQIv7
ch3kSfQaXdC/ECbLm9zLwg6Z1G7ii8vJtVo1DPJSQM2Ddn7PswA6MIyoqDk0HacS
rKZ64k1QQwgpoQ1XsVBNxP9WgqVS4c0xc4xmEjVdCQo27W53sYFS9BDIkjREeOl6
YWneN4dAXfd5X/Iwnwmvpa7/uVicIsmI5J4oRO5hFfgFJBcSIf9nUyvn8xFUkuvg
/7aKpBmeWAG35esHkJWU3AlJ06GgKKZTbPCbw436Pe29wPqQ+J7GEPBnhGeLloIs
2tdAS+Z64nFIx1g+JkHQ9fv2HWeIJ/0yc+Uw+vghDSN3NdU/qEy9OOSIliNSkhCp
yLipsqQrCICfPt5s1HQwABY9Lquah4yz7e4CPuShyK+mbL3pWLMGE5/ufziigmsg
AydIVuVrWaqXldCF0LxKE0rFfMynladImZrEMSBq5SDGUYunzWdbWpeX6fnqjEhN
9ehkDw+GO+ffKFvjVqV5k4KDEpLKpq6cBfeFGMX/ZeDMxN2oNmEqj2KLCrh+Lzh4
sBUeyDCgKYjnQXkovzf87YvAO7KAjc7KY0y06fLpV3Q7KhQzykC+UoPAl3M6fVfR
HUc24r42tkmuQu5zNrRi9aQVTLIsxGKG1FDLwCbrkDnFCbGceBFambGvhkIE1p8R
ewcurDUpCvFEwken2yFBc3/+L+Hnyh+N7k0ugFLSpIe60pant7VvZCb0gYkDZf3f
+WpNQcEpaAiRnl7gQPPVGF1UMNlltV3EhyA7ojNmhtdLJxsac+o2ts879TbllJQ9
y2pYpeYkB5HwG2c0pUwmpdMBOQgXatwnw6LGLVogYYWXwGHKdwGZEX9SOjBd9KtG
SFPFuykJPwzTQ/b7EbIX1fW+w322u4CshIidlZSMqQdVTX0en6hfAQRe6uw/J2fx
GDkvCVKzXpcvs3zDM1+TvZrXTogAsyWywux3Awa1Kn7vpAX+jexH3E8JIRdaO3+G
b72mYVAtoyLti4mG9CWwPk5UPWUYkgx0YZcrvh80gfXq6ZInCwfJUiTDyUHXK+eK
XDA1R8AfwEM7IlFgETPbL84Imn6cfrXtC8iuT8ECL0wGdSxd6k5HXHZxSwqCeK2A
TJsWkDv2WCo8hXhJ3vKr2JS4Y/S0G6i+Z4iODhm1li6p9Tlc7mj1p6SagQTMe9CE
GKtXTYoPRkI3adLrZZRJ4HEOoDrWx6pR3za32tzqjJ5oveIj8+QoZ/fcnTqYMnWM
xrMGBAMz6pwDuwqeh/4mFHZrlvskHzBxZFMa8MSBmQkZ+3RLCIsoPNdUIDOBu+Vc
zEPDvT5jLUQrIerC2vRU+ECt0AKE85xb8lKABLwKEmgn9TBRTgGAcatoPlFiT+Mx
qyNDktzyVgqr8v/c3NRViNJPtjbvy5n4YCahn0yJ/b0z4n4WsVc6h+NuTeKuy0NF
xp+TEUb5f9dSbbhVxCu8tWrkRNcrCPyanua7mb4mRPgMaxQFSV/ZL5hy55aX/sNJ
C5UcBPWgSMZ4tWg3a0t1nxIvQfgm41VQ4a8mgrqMPqbr/KF20CQC7ScGvNzdqzTC
oS9ROqr9dYn533K38V+yDLOzl+O7AC8QAy7KfkK6biEX8/hRs5RuMbkNWVtWbNRf
3CSaphD78KyzK/+MapLirbotOUNyIPlb6wcj2kyPJJwbjIPZOwYbE5zlgn7k5N3O
6+SOK4GTRi35eNXkeULJnXpv93V8addkuMcJFq2ylF1AFI4aOxTUigMmTxO0NoLD
bV9OXKzrTtWwXFk5NKluWKakJ8A9HpoobRZxYavZePFPcq39ZzAjwycE48TQLDnL
tRbD4rH8EDJEEzDhDNcYOJBm/lxwVqRQ+kaODckUVf0h6pMulnAWVRPPEn4knuZG
iID9bMVIG3cVhAjLW3G2cMXmXbk7FZfZWLo2WpSHPPtv8wzu4SGMXEP/27ryAdC4
AzRPv7srdcHhEJ3Zyg1t3qBg3goi5dIyw2FmT6tx3kVeeDkv4fyabWdkKm+8a2an
K28BLiOxTb/wXbnZQQujRNwnlHxg2XSqBCo7vcm/hxOLsZUiivxkpSlU1F5W1UEX
phDHC31G5OwotWJRNK7SseCOBC1SjB4erEoC/Xvpi361s5RpwesB/Oxm3bDUwi+r
uT6ZP8CQ7+8i39hs49ZWvgY58Vv2SPl2diNZNktvAS5m7WfQUp50DvAnTHVhL5F4
qSq64JDEbRzEAPdck+5VUMqPZ12RF/kjV7Pf9VRIW79lPXNqzaJNlyKY1BEwuijD
9HKrLTzyTU38tmA8EAzzPumnRef6YA3/HahBjeu42xIuNdyIuTDJxQ2VFf8FtNWc
B9TiLAz0RAUS66mYX+dPr/bJVQGWoQ2Mo1WcQPqUd6nHy1axLBMz/brHaSuj4KNM
H3tf/dxGjWGBIpYYYyrozfugTVoinjBLLml1ITqcXPSfe4WXWkQlRnfHNnbFzzsz
BXwEfks9950y19pqIxb0LMmOEIhxRxx6vl5GuVbGXnmo3S9zXEd3vstZdcfeVQFv
XJgUapJRZTSJitlxvxGoOyh5RID0SjaAsKjWlH3SaqvfNC/DxsLLEB66zgcWP1p9
ggAbqCqFKLzO+9NqYra3FB4QozOD5CsC1s1nwHL25OvdymDvwF2/BEEdUmxCgt0u
RDY6GNc6Ksj0rtibTndFO5Oe2nEAvGJuCSb+RNz9bw6kH4LfEFna/qhdm/fleGnT
rhYqNGCbZdpPoQHeDdigtdST317as/2291S6+j5axZOX9pJG+CF4RW3Vhnv2dVqe
XPUdd5lhIyBIkJ58JEphFYDKp/MCg9zNqssNOHQJCOdUudIg3jLPjVQyJHA++tt9
bGWUE9CEpsKUWR1SoCKJbTz53jPTQxQAdSWTPSSnobE94AQHvV3Kje4zL2zBijwU
FQ0qdbar9pg0InyfI1iznnRUwYNx6Rb/LAbzV9GGCsC6CG4nm1iuFIxxWtHZjuwL
TehcsCdqtsx5Y3YHkvqvsuM6U/RGHiSc9UOSQ/SxAcDFbp241Q3brqD5oNMxzqxV
C+Mr/9DqqZ/0QgllLN6lli4ILfxYmepyBqJzsGICjimpC3fy+azf1TP8hSksvIxP
VlzVoiYCIUIW9D4zwCB2cSND2Lx905KbghHwyoukbcI0qv1eS3g+AILySba7px2T
P+te3EoQDSnSBS7PY0Uv+39cpDlBXZc6RSVNX4j60mF2kSPJSc53A5/ZekPxHLTT
RWqUAc76vX9tp+BBOQZtrsvYUgLbFpvcVVqzAzGyPc14NkyRohiJ7LlaR6L3t51s
7g7h6xTAtCYoKImxIlWluaLKjywRrG97Iop7apZ9BI2MIc5ydIn5i9QLdxPvz9CV
AZHqyOlRSp4hG6GdUyaHkcTarCnplsduB86dGTr8cD2fLjH6eJVuOrWKMJ0z4Azs
hOoxcG6yfulL2KgyO6zKYUadoInBpKNH/tVgIPXE18BGtUwomZOULw6B/xQNOjJk
sNjeohmqlLChQ5kk39xFSgrqqrcrTn1GZzmsAsEqc1pIB+O5q5vxxC6dqWjmv4qU
S4kShtsZbJqIKrWxyUd1ivSzgWH2RH/QxyA3OK9qCn00zykbi7DlgQKxBxntihWQ
gGoewW9lZImnsTGjpIEhX5Sl1iM9QHkqECTEmsZ/4CKJXh9+MANtnKjSP3vEbgHX
OTLsaErgFeMy9Zyd1uGrDrwkpY3SiQ/ji+iQlE7lnXNiueoOQwhwoVSBL4+DdbFz
AA+j4GKkxoDeh0pJjAovjXH7Vv8B53tvQ2ps+arjQLbr7tJeuPsi+O0JHRrwpXIW
tlto4LLGf+zhwpIjPJzKtTTUVhTAIlzjKblCYRv4OGxoAx+jLz8FmJ4fIR01MMGP
JeRzgeRKR8Q7xQJ4/fyJ8oA2JaFL6scoBLjTKWbFnVVVyJjOA0Yzv6cZ3LwyAkBh
12gUqbdUhRmc90BRMErDCTUgDTojvC3M1ZGgirffyjz2Ab0t8cR57jCmwJyeaF/g
KoCUV/mNsL2g1lg8A5b5WN7l6kHAXUX9NeFJ84+Eh/0skhGtYiaeBQlhvlOHWp4+
xuTiTDyDVOu5h4HhbkYQBjPZ5EyQG7hT0OAnz2JqzylAogV/Hh5hQ1BJ6VN7LcyK
PTKmkjn8TZFGVpAzPiyG83OLGorIQf8XCHT2SM0Dh6o7eEgjHmRsec3Yy9bBl+bc
Ucm19fdbbATCdizmxL/NehrHg74Limwuf0oApxc94s5HDnGMvitBTdMBRAguRHWw
8NGNz/WMXQhYINK0MJ2XIUaJW699TKoLstAvNHRUbjKsfLy7gstNz2onFVIc6Cyt
orSBY8nQsNns3baPzHJs5oY5nBPGDn+XajgZbCrRVIVuyF/K4bnpKih3GeUqhDdp
WOd9elpPCaXyGa9ICfllmvJoMU8RugTGA74p2TC7qw6T8vZtzROxqlkMkPh/MCyf
PppBjPFuMl3uyDOSkOS9phU3la6kcwn7YcAxfxMdmKHqpDubGgGtkEqCv/E0X5Om
HOjKPIMHW5AovX3OyAYMwMzkZH91R5mIhE7d3mN8wl0nQ5+aowfhoQgXDNepqEeB
VAYMNCQtNowIEI62u/n5WP+xlTGl3XzVoLCKge5ICWzVEXIRK+M1vGBSkCX23EWD
1GksO0FK25Mi4PngPXc8az9R2WanU+/GoKll+xVPSYzUFqqRJsG1NGrUea0h3SPD
wNEWx3yHS5ibsBQQe7KkSoasbURxfv6Ziyv3x4rKcUq0Ddpf+NTrcAB8fYU3zuy7
zSgDHdPNxfGxrDsYEjFW0tFJc8T6HLt/567IdmGOplBkI8rhLYmLrNg2CJulfjU5
bwrLZwckDpWx1+4R8VxOcUJg6rBJ3uJ/3JcLynmfLTLYdXjwSyumX8OnYG/DGBa4
+l2SatM28YJjINZoTPHUzERJi8kbf7X7gzFuvXUWXyfZBo2/VAVudsUtXF3U2bXB
iECNtUOHWjByoLenamQhLjTCZL1yDY5jn205BnkkUDTm3Mu9RghfqJUqraDMzR8l
jBIqXKbcDI2aNq0u0Th4fJdzlhbrqgMd92Nn/ZGMgNnh2PpNxjIG7klSjQj2K+jF
gXvCMZ08Yur/g6+i6aUYHHF0reQXkFehiQfqnvjssMWwSp8NpZ8qr3yO7ZeWWpfN
BY6efjLdokXsCwMKSTnG5Fh/7Y7FzKhfZ50r0F9PJz7o+aaWfIrcufsbaMFDdkYB
flAbZ4yRZobMGAFlpmqMUfS2DEq5BiqjOyyumxVqTyWVJJBxNV5TY4uuUYWYyfeH
L/j88rCdN1Nt/WCLfHLHGKtTDwiw9yXepmLfFA58HgjbLX6IjtgqmvWDzTHjglha
IhmjtdkZsQ6IYlS2B+RAS+RwzuFxx4CLiPOubWvooeBehq3MSY+kG1NuBKHwemUd
+6MocGYHnJ1Ep1jncqMa1lA7PRXndXnwPu+s1e9ywUgcmkXx+aXD+rXQIABJhE0a
x3KBALXSByE8UEJDfwLgtazkkWJ6XrBIFxgmgM49MtEA06Oyd+y9XiTfJSsCEVK/
BLr92D2ox7ypJ6ufplWyKdgqjKjgFAUesZEvYeI9Vm/TUuPyXAl5t5R3FxJYbRjf
3aPwNAIG96z5rORVn9AhpOuauwlu/EJkgtsAzkP6tj434lcnpoFT7ISvuosIUv/w
WGruXzXcCXpVbvM0IFtvJEQktun5Bkylh2keA/Iw+bGg49TwD0bTjMJlMLRTZjlF
rPvZYB50rEgMRj40tpWAHojt8DxUNQBBEiAH65TI9FAHjFOenfXyfOWtuN+ctVMo
gbJeb1OrePUUzxPQNoS+CMUlK8uI13unv8yHpDTSAXTHlS9IfeqYffP5uYvpn41s
78d73ArR8TvDhWOMhFTQiVtWPfHH5YJIctbbWMzK53Law2KjG4fZRoZkxfnLvBj+
wKMNTRyPHFaJyReySvJ2CgDncy+uSbjGIIxa1Kw4Kxr+Harf3I7LqHaLhBjYKn8o
fLyl1CxSTXCR0PtKypMF3k46a582W5XKTa2ox3VfZsDrr0LZ2Og/cdQOMv1VetN2
db27f2nunNUwrh2Rpbg5tihLchYhfn1P6As2G2GFIulR+dT3B1NyWO7HgGHemfa9
aJZ1Q+v/wpuAjvgwL9PMr1IlCNmx3oRKBaamFER9GhhSFNqrEwa/vIMqcUMYUQta
GDJHTm5W8lyMBwesZC739a0mkPf3Q1Ydaxk9IQemZOdFNG8woc0HCeZETzIIKfoU
UDrgXyl5Efd/bgjg+zAGt0QGsgxB4OXBBPUcCzmsS94X/zlR7GeYxf7sDH6eoa33
0EL230JjVVHcIGRpB9bjHwAhXJYoXYlFqwHfM2Y6WNTrAcAXbYolJNVCtPCEGweM
KxiXi16nAUBBBa1+39Vw0VbPzVG4SgaTbFyMplxSTd7VnI8jQi0VFCsgrGELjjKR
mvY3rYcQarEhHJtLM//MTv4V5B6+bD8zY9U0UvUdVdQP3UdAX+avOmRGIuz6ZJ8U
h0WYHcNCq4s7xZpEUdVOTlV8C4Du2jKcefQBjgQtvFm2J3zWxO2knlzff6O9rVSB
YXSkJv/lFkA4tlSfUh7mBJ008jc6MevogiVrh+0Tu9mxl8pj71YtOUkp7PZwFzMV
vkGoezTZgxaXLMo9orkyTr/G6D6rkuXgBNC4rdaXPFEGOXuGROXQ5Akvn/KczWBv
9azHdmMxbhluRdkLY7rqgF0uqEKYBfPvN/J/k0k3b3FwBZjf+GkGk6Dy6eMarC3d
hfABOI7rM502hunbsEzsPWDXBhuMKm1P4NVEPlTLL6aAkiU1t/5s3tdanQyK1Xo/
o4P9OzSoAc2KC0H7qjkoOGXou5zMKQ0pNan89Ln4TQWjKOFU30dsqP7OvSfRwzIC
rMVPLEpxtQoXs7gIhHDns/zlkNVDItxr/N9goc+l/JUs9JxShwn9oAahULSw4ak3
r3B4L1ycDH9aIxPotEPFyxp30VM2tyA2dRqAWuJ5yzaK+1fWMT6v01gbTfTENcnh
TBYDAoPuQ6CD2FgiI2ZjXfcYtLmLGqpdWhqTga897wvh9dp78RIGv5ja4nh7tmpk
Fsm21bDMtCUgpC4hn9q2XU3bMZBhtr5yWm3AStUGUxZuNiyLjQi/9sS3NuGITKe6
OYmGM5UfQ0kwzAZZCVNHPsoRlznZjgAV4BpuVLZWAoz9oYWxIQUZPJrdPnnYlUqc
b7fGeL+0c7b4TuE4fUZJB3S5cTI5okAAaGtkOdPQJ+8oZhfHmP1OmrGjIh900xJs
Px2cHMS/RkWJ+10S2xYJmR0Me/0FwLlzzwaYAcFL3SzkCedCmfaZVr1G1mjF/zWL
iRoJByAZ/C0ctOPo7mQR2inOWV/OgFklkcrELoSMU2EkSqkJyNzevLG7xIvD2xsP
edYUPsio8AnFVOZSrzFyB96ND+dSgtyCZ7wdCy6oHMwz6jUfQ29JqS3e5dTGbVRm
bx3UD6BLW5XfgqmIVD+v+8Qx+LvCY1+OoqzDxYBj/Qm32OAemmzsC9ZjwfGfWgl5
dAT7giKbXdnz3jpRrqbnL+GCMxtdsIileXTjsGZUKuZfySKKYHhUxgUmd29a0cbX
92W1SKBwQnB8MXO/yrpqw1g89mI+noefi4eJB+Cb5LvqXqHmm4K5LInVQbowvWdV
mV18RikwyopbNT1DNRg+DoDU3O4tEPbrDcahjeIgR/+INzYb5nTVsV1ZzYYSjHBe
xm/rVdJfqz/imAjc8qBHyS68WDuugHzCRfG1SAZ/bLc5Dn148/paBZT++9xQ0kqF
y+uliyoQmkThFkAE1P/ZSwaac+OmpvbLdnP0NN5ASWTzZOe13eVI9FnxQz5sWDuG
buJVD2wqHRwBjNei1vA4yYzeXIfSOUA82J6z8pgdUaHn6XRdciB/sTtVmlK3kwGy
t0gN15uGuJ76lcTb1Hsuzaq8gqjKTrNxLpAfjMaJ80ykniwyQq+m4nxGWOSax46L
fMbcvrD/fzHPiSN1cHm6qW5qqtavy/l6evr/f7cmX/xEI/pHlz30mVsnhP+/gR5A
9sCkvdSDMRTJXWiKW3eGeTgw+VZrh1vH3BRwVSnbWMVB4Npw91nLpIWWBfECImXe
s5O/RGAjg3z236bxNe0OETCscQ8qVu3+2mW8NNE+MQUDc79CA0IUnUmp2pLm1FW9
gL3lt1j/r2rSayW4WZLwsudO/fIF28b2oXSVp34nE9yNcjKG0kSTUu5DUHx+lCJ3
e+yE48sEHsdcn3Wrtlft+CSEs7VzFdvaDbqZyeffmtTOeJm6HY3vFdgUcD1WpWAc
xzp9WzROhWSKIJvNcVga94xAb3fbIwWMGEbLnG5etmrhAw2apERjLRrm8DFAe1Rc
ZVRT7qUTmZMmRxCdpPYTTQ==
`pragma protect end_protected
