��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)��΄���yN�';�2R�D�Hঊ'->��n2u��#H2\���<�n�� ��x��`Iiou�З���)�-0����V���9O� 0b�+X�6�w5��i�K�E*�=��*�Ƥ5j��*�&/3����۔gv\κ����-��V�+��/_��j���4�62��su;D��A��y�0�vP���e�,�G��/ms�
45Y�Ƒ�P��q
�?8j�H�XQ�e��mb ASi�j�,�u[��%\��r(;�q�R��׎AE]ƾn@��I���:h��a�}�")X�:7��v���\���QPx��.w�g�e���5�M㽹9Ih�R���A��+�$�k9o����߅z
S�`e��f�&�M��'$^F| \�r<0U��y�&�%�^P�_��:׊U5.F�D��C�8q�:zK��w}"���r;h��	lO���/5{:E�{	-q����ڠhP?�}�#׬�ܮ<M��h4�!1����n����T%V9��v�c�T����8&�Z�!�~M��zjI�йl�4�[��oj���j���s�ט�/�����kWm]��/=~��*I9� �4�Z6(ǚ�� 0J�E0�V��yZCs����vd	����ۧ��HsQ��5@�tB�6TA~�^8�P���:� 6��߃���9�́���<�,��aF���6�h_2�0��5)�����K/6A,V��^'�����f��|	�&s叺�6qa,ON���Wu �ш�ʅ��c�x������*�1��E	��<{����튯7������rn��2��xpxnB7�A=������{��O�l�a�~h̿��ޤyq�p�,�'%v�Jl:N6�2v�f��c����f�����-��
1�پ�����ș���,���=%AJ��4�"h�۷��Y��V�:�<9��{O����;��������k�S
��.M?(��z�̴�jh�E�������JN�:N	,]	��V�4CXh�C�.)����M,��.i�����[���#l���&���X�Zn	����&��N&K��Q��^vw��I�#S=?t�2���U��?�k�޴�L@���ڕ�c�M��K��$�1�1�})�#�K;(om�:|�B�ߓ���3���n�>��j���zK�)J�~Jd�9F�c(.	�7f����X�+	E�vy3�T�}cC����v"�eۨu�OE��