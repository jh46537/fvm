// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:54 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
A/1VH2OHbWT7fKbkL272eHaO5CcpjBAbv9yQt2B8lmvJ2e+Dex+EPaWYFqMLabJ3
dvxJo5MPvh5oOej0BkunH2tWWs0nZI0pqrX9Cvsz8AxSzxPbNjFcpNBCz/lDB0RE
v1k+4EtyigmI2BjqUMxrv9NRcST9pYWPW2xeLqcj8AA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 135456)
pbZ2ceRSeplMZ4m4dc6RXNDDE6lU44cK7nI2zc8azdgHdo5rgT/kZ5CBjM9qOFnh
Y/lzfkoMuWmjP3aFXQv1igQxcBI5jAX4fHcmZaz4YgDNJihX7VXtcRzI2GbhGXo1
yXo5OjxLLzxYtsda9V9sYqc0Zmx5NzMjVND7dCEAJMFwazHZ2n96Ijz20mAHqeFq
iWY2z3ijsjchuRoTHy5zQ8/SDUyapuFuvmAaKKeuCvgNKk4bal7w+tMuHk3ZbK/H
QBfZZrK2BExNOFbOfWLgbPDolIx5UcTb5lZcaGeNVAMwNArc7MzxJckyl+ygyhk/
l+DGA0DqwzPYKVcgcb1+/i90idHJtwytrjusAg8FIdXW/3jhkK0j6mdhSuJVkrGG
Edmo/f3RWZtxrsc5fn3B9NYk2OWNip1sUBdOPpJNkevqRzSP0GKzuogDC0lmrDJU
GnBiceeqkwSZWt/kHsIvbG5uBRxccoSD1cOzytphqRGLPPrDxCou4O0jyTxcX30R
x1uDltCYYhyCVVrAH4PU49S+1usSc8j26bAtnEEm0V0fWe/Wz0u/g+hBci0mpcJf
npHL1p6GbiarOATEal6DsvoljFsDPRni+BCg8y7xcL5FSuZnoqY32HS9HiHzeNpN
i4HntRj1Se4PInKUc169fY+Y+eHy3L9992qUsX/WHMbH6fqG5M0v9xFrgZKYH4IP
Ij61voUc3ZeWbChGCIsaZCPBukeSdDTby7W8DTl5rbs17vB1gSUNyrnKzJD92kdC
Io6+vrwWN+RuFTSImlsQgVxODS2qkVnWmJdHTPgDDAQ2GOpdTlgns9IQAYI99to2
aYnylDSlmRSQejzwuoJSPXRiEc96O5GDcq9kqYt1E9hvsjutXIc4Hg9Dx3beiw6i
vDoAVXULwfqaG9/oKzse4jYJ89HRdPdgS43Kkv+KWitQR1TQ9mnYhLUEwuW+MW1C
qCgXR+RC12wlFoL18fryHE7dAGGuxMGdLpQ2ixgrjlxfNFlqJDoxcvxrdwkzVYhC
ZDi/ieMelpM1AaaKfE/f2O7XE7y/M1+s5NlGYpuw/Kw+aYYH9y42Cn87vsJfFrBk
kNi+jW+6aYotHQngCo9VGObp4Sqts4AKc4BDcylTVzi7DyC4ZgpD8Y1ggy9Wy6dg
2MZxvx8JwVnrvUoiF4abinT6ZajIvbbPl8SrhJI8NkdyiIhAFgYWkgNgn1E0VYcO
+/4rVWkvdJXMFArKXBEzWyofxDHRzW7ey79C6BBYxf5qgbRucADnICmXetNZkLjg
D0rxejHuxBKDbtJfS5uMPsjV23A+0u8UdY7CvOxCghmy2Ymgw5X4HisEG0zaaOFx
3iU/acO5+ZN9hMcBeD+uzQk941pcUmEOauddqwt9NQdmevVNNeY8h3Ye97vTTOV7
HXKzl5J29Nx0IsyghyeES1/FYlfvSGSP7dDcppBf7NfoikyIz6xMWIrgV3EibrIv
MLAfNH1fduqno8MSWKY4GVAxcTxrFmIVhv9g/hOHet/yRzncTmfOVMYak2w98z65
Ac1YWR3jCKg4d+D8plwORLu4xazC44o9mj2eQs0CLq5ENinYdyeOSNEFG4mnWdgy
/XAp4utBBbtUmV+Mk5e3FtcxDb3YOJgOaQrL5AyXEzLpsTAbgXVA3VODUIefgJXo
gqsGRRWmQhnFcOUd5rL9+CTlOb3psSF+Da1aB5ILIRvd/lXYW1UU+l/Nb7E9Ng6o
RUkou8X26cDSKl8DK+omRzhkf/uESyZbvdaFzg+ocGicP+sxayPRWPm98rxY+hsz
BGq5ftG2kcY3x2Lx/07NduBlDLtf/jdVrZZju4wyTOSUdE5ghcM6SoMrRYksg2iE
dGGtzhIZ4OlTl3eSbhA+WnOACKtEDP4yBPxPFsOh4tnB3ptYA84lbTFpS0lcvSPc
Hzj+1nDNPlzVO22MHHqMnjz06wdX2vk+5N9gsyJk6h7vvXefzZXU6laqDL4AxkCv
3tk5ELbRsAN+NKKNLk6gXZnMM9/RpNS+7tZKwhH0b2Ue6qjbvBdA226/CibypiIr
OJdh6DYJ8CyOaSpRpExngblUKBJexTfRXs8dWvxcsIvlO/h/QZfkfTGpvFkjwaK1
VDbepIQC8lkP/Q8jm70dEKNIhGDbUOlpuYeh8nOnAWqWDNYHgQon+8w6SjX3+AbO
jPKgdsMM6wfkBWL5GJkcWNCpCuD0I4tG0pwOcwlHc306mz2lM2VLrKxGYPV8/bwc
qRDbG1IqszSTxrBYHEP05esI4aF6zds27BKmY5cPk2KvMXIgR4lRLO6ScP6ofl7Y
jpsVF4wPyoMExRu4yQj6GRjHpGO5ZMBFu075066ziJwWHtERHem9octNIklo+fqR
p+KcTDkedGP4wSQUS/qcHgtYX9+yyM/wJ3KxMiTc+wiPRb1beKmPAv1rkNevcxs+
g/IVGmjb+z0HaQ4F2x38ddQRW6tpjfs0gIbsJofmDPGWc/DhGy6JNFgNbmCFPd3Z
BYZssmuyJqJEhbQE2UuFZ/X80z5n5H7qhbbXSL7WciquSx9BHUZ+u7JqGTZyvLAT
T5KxctO8R6/KksIRNt28Y90R5hecVxbXf6zZmHWUyuJGowho4qnVI/FqVkByTxkW
pX1GMDTKPFT2gey1DVPl4cYa+YLH4AiY7cc1iiCho6VUsr15O8NARA64LalG9Q+g
sZ0DI1O2LNK6lAmFy0eZM6cjdY+O57njz1rqWPYrhI95OSvCqUw2QIVVsXTpqY8r
V8z1CqAUi77pyzupUYyapCzWYREyj3XVcKYudez8YquqIfUI+WTf0FCdCR73N2VG
RQnY6A+7QhOTvnPSaEFjXm+wW1Tqjwk5W5rfuUs/Mkvt3SbF6JU9AqCzFUPobvL7
NP0e+DGLCr0VG6IJRnEI0WLWyHuj1Y9is/MYTy1cioDeh4wtMfGKjSesWMs+lIov
jHaRk/qvbnA6zltf+0CnWZR6EUP8/m2nCDF/8VYAB8O3Hi1CPg+6JueLTTnibznN
Z4bVk90O8e2rB61A+rQtQ3NGDoIuO20w+X4Lslia+K0hG0BkapThHHFNwJtWAQjR
CDS1ECouDfjZOlDNi6A45do8jwUmS3kIhKvzPD+s/QXOjNKPY3oNa2XczNKomtXo
mgjMicAL615DYavIoXTvLlDgleH0OhKllaiIAWELuHc76aVdNbS3EtFQmhye1kU+
Gs7zTKpzTK/O1HqK+Jlz7CvUfvmshnqnm7ChLMjfskUE7+l/ToVRNjf6+pKuZFh6
Y5JJcsyR6dlhJem/DTxrGAa1oaZcxvcyDCR6ENY/Aae7aAmrErNIiahNWzItvWep
kbj0fUp+rnIbY+6waKxgCd8j8Rr8e+CEdsAKQn/StMPlqhpvIPE3FeReJttx3DxQ
scKeKIUyIhEK2ncyoVQJCls10WDLoTk0BIHrpAr/1vfKhW7sLxWiOSyTA/MZ18YK
kSzghrz86U68Q95By8TG54QNPD/C3adtRHIm1Z4nKGY4BJ0swS1uVcyCAyu4ne1J
owyeuNg9MDOFY9KTQU2Mrg5znrCsnr7tKDQABeDIR56yVGHBm2uEiQYOoRD9Qbpu
3Ks0BVnCod8Pxugx5jL6R1Uvsi7oOkdToj1V4GAh/8QhGAa+bUVWmjWP8Gh7CVT0
AFKcELDGZ9YZ056UnNUyApECSajGyYY0cinio0YxiwyIKBbig3UnPYnUNqztTjYW
7v7wYxFDubj2yJp1Bl6yPHWAGcP77L5u8ne+wijcmL4SWmXlfza6JWYw48esC5UX
dsQpIY29Ud9NLZGyXSwT+R2vRXLTXTcCdutM+ktXykDFymlpbm8wg61QEXH3wUq4
wMQEO9twNldNj9ijvZPC7ar1nYZ+HKZc6bLts31zjVMh1BlNHYUX5Ldtvkp7Zhnu
DU4yuUR8mF4RqTR05TUQm4G31YM6x6aKjTEHKjdygw5FJkwJM5JjyjIAWYosdFt9
nBDok7v9FyuNoN7YPQT/xIUB3t4AXR7lFdQFzuNLfNfMkpN3bDrx+b4eMtmcOOmi
Xuxd5d11amSObM0bwlQIgp5khipfEHIqobUYKUf/VhOjq2aAC3wWSqENNX5+UuQ+
m6fQnnJw54UbYV6RPmkFQ3wJPyNZ3oZhsXg5wk9gPq3ggZEThMyM8hUcvhL+ZdwR
bmqhiriuI0eIJ/jk6etEkZE9dkwC7MYUJIMa60T6fOJs+a7siMr8gqwgtaXeCcOR
BBuQ/e8EgtD0y+Nwv76xRk3qSvQ56mHCgttTX6ei2lNfOwKaNftS0hqF0XEkUS/y
U6KWOBQbLy7IJfU36oCfGqRBFbNuay6soorbxsnwXjwWbM2e4sP/yygYM2YeTOxm
3iqj1dMFVRN3nCezIP8rX9VkMkVm7jFR+SQckaS+ejS1RYYaw9I9Q2IU/HIVZ247
w/ib4s5495ZUx7j6D0Wcd3J/A4ne68L0mpyKo49yuVT312atdKahjea54xAN+a8x
ponNYaeBgGI8Ac1pc7K46gTN5ivsaq7uxivWXpTDr68DA9VerGD/Lsa2l2YjjbCj
484CjDJ+5We0ItsYKGHz3Fjp11XkQ+pzfKdcCtC+njOF151cyr90yC9kAPdBOoBz
SgaUkSd3ArS3fSRd8BKf0AR/RlyIsMkg0iYrmUWw9diVXLKosQ557aQ/paxERdt2
k6i5U9w8r9h6oM3GBL5K9QyM47wQNb2QQK4g24qscfendUTIKI2PwOTc8NGO9NXf
g7kUjGfdxtbq071Ye97F4tKx5W7XclrwNYudjzl/SSuofaoUIu98uKOfoFbvf9KX
pTEZGJOah/J2lFrAqcmWlmzyLPv3DR5X4vohg1u0jrLeb5iirD03chRBpB4JOhWo
GlSzeoopve3+qBLGw7y+0d6h6S3BQRdk3acxlcZUHKnh4nQvtc3A7Y0mOqp+t5Wd
zgRwlj3H/lYV5TJ8VUb19wBxQ9fDxadpOeTNfeTczSaMu3jozeVa7ymoAYNbgwqe
FI3TMRT9cm5IhaVF/k84Wdlh+R8tvA4EHYPzG45CpkfzsRrKX91sL0qpyfGfRsZK
Omf0nSl3JnZlA18b+V8osquIpIOsooBJ/a9s4efK6xCF50gt2GtzDmUjlt5ZNvlw
/wcyadf0PwIWrmcZAJgQU384CetRADT1L4QPHZPD4z6n2W7HgUsU/W03qSI1nMzK
R8Oz/pTuuC9N29hRJs4+nHLPbHhBHsGcXiAShYJzh34e+1KZK38M7MqFAlqVoaxJ
lqtDxEe+9tnf/P/91EiQWdC9v91AUYmnLk00RSmc5hBPF6y70dPyT4j929ND9p+1
o+2pUNRzZPMstOfDmJqJ/EjsVKFPoD4WM2zVvkciu0Kncyy6vOX368d+LgH6OP6A
CgbHrehW4WAfRYWbOEmr7Cxz6dhqMHy58MtsGnR6rgg5r1IYcz9ddegQShxcqZCU
FZnhdzb9La9K49n+bgli7Pbg8BlmCrV/X9WhhATWqPdl6wx5Je6J4hhoBiTdgSmG
rWv36Pm3kSNDRteiFLaI6VNvvzyHbSqtxCESM3iXU4FFRfmdQcBsN78g/lyB7CLV
7Zv9XiKX0tF6OExYtwDl76L89fZF7hBg/IG7mJRVjxCocg7OA56mFnypfav+81a7
Tqu4cry/XGyE+mUijTYAarybm4P88CCYRQxLRGCuibXVRBHNSDlWgqeJHoQhQBkx
YSYqPDCOApk1zBrSBnhl7xZl1Md2NBErvRYL1AuNN5ExICUYAMi6PUCdMqMWH236
3rvf6+8vFfWOcCVQxcdIOJ9WlzCzAVPSHO28P3SiHieYpG5n0O1M31nmQWHPJBF5
w8ebB3M98alUBj9fnOyTHlgOnTYEx81Jhd1gfCbGIXe7IhuujT+X4IG6KJeP/c7R
ic2vl7cP7q4VnpG+QPMrvORLF2SOMeVTYfwhN2oVJ1I9z7J2nCYrY5kNwbHvUYVr
PYwp4TxuzxS83VYd7PItbUTFl2S+t4S/X8FcP5mElAyaZ/E90CF+wSyXA187UE+3
9MqxdkPIQS6SzpngQ4Xxt9yv+WK8GzOOYnse7IAV1zwJVvryppQuaWmJMJ2VEBNQ
lQuy4E956xR1J+Ee7qHC1EYdeEnw97KFHhl1bpvLasUYrm3y5d2mCOj/zWAc3623
h/hvzY8rz8xZRbrhIon7YuvbgzHZToMhi4P+2F27ddqWRz9OhTW92uGRLySXgRTh
PnxqFAPQDVLloibhNdWBlsET6wV45e6NxGmNv3IsbIzYCz0v7O2FOJvbFlPGZocx
Ol8PRd79d+sk+ltSTwkoeN4eYSFx894gITJijYOp0K8TBGrpOtAHNdysFRf/kwvD
4rC5zYOzwEV1Ihf2WUFePaIqvA8npqyxZsrMdhxR0PejmzNzJmaGrisFsT7UDO1d
AQqwHw8xI1nQiDn/QAc9xzSkjRo6Q65rXcFTrvDFLHrl406+OtYi1+NwPNEI6VI/
OYsJ9dTG4HMnOzLFhl8azvW7pMC4jJm6CxqITUs1jnQrP+HxPuTMxR4ftp5KKX/K
/4xnSsBALlInmBfZm/BLBgxCiq3/NoJqlWYlfl4CpEuWNM/h20nXmRMo4936uDE/
lmiWic2NpnYTsjwWi0gx/9Z5X2HTfqy9ivkI8Ig0slJXfnN6ArZqH3CCWEJGOLqH
n+IhyyWCtEKARajwgIJbnO7kOLBZuGIvw+XTnkKV3eebwK2ds7JUL1nML8KDE1o3
wAHQsySCx1/lEu7/jRinDov/D5Wj9UToSogJHjIdG905+MkKaxGRHtRJu6+42mk1
LpUyIDcorYbc/EL7xHizU2cHP+fmXW/bd/GcfQOfEbewJPmAvPzyZEaJ29Vl+ozB
DAxx835kpaz6lbzCavYwomW4w71OQ1+cthhfapRCLyXgzus9piXgkucbNTCQE9Es
VvZgXmIxDGe0WfkBZqZ5A+Qvc0UcSPnO1oZaADi1mecNywX5he96wttTci3JetT2
BfadwHUHnzi3Nj3l58HcNy66p7WJkLAFSLmd8wiZGsY7bhbdLT9iIwV0OgKcvaBi
jaesRKbVLhvtcJHEleJT92Ss00gTxM1VcbK09ytoIvR6le1LWFZ2ewntnNszqjc0
873AsePagJetyikFXPGNDVsm18/E/C4e9jJmhHAu0eHZRVnKgfyCBeI/RTJtZ5k2
6/fIpqJs8nAMEI3VusBCZyFodn2RM/HR9CS0umPtvAcdzlforpSrj+HbLJzwPn0c
9TgWFO0R0qOwIV30nxElITox3D6kQLX/fVm/RfRgJj4sQW7HO00/fKfmjtED+fHO
dAkDSQ4dJVRGBkyDRVBVcb3DUBSgSMIUSi6j2wYd4r09zaDwHYb5Ouj+QfAwGbH6
XnNXnE67JvGznCaJ2F9ZCpGM6kzbgddZ+4P7K8pK63tzH1/oINEnEEcZkOJO8rqD
oukpJsYvZpyEfPFLQcFW9QTMQL20e2qXEulbAg0ajxd2PayUAsNK3f5WUOzK0g7H
RjarfHYTOqb1UQNhLZVUkxPfmW4mOoqNEASG2pcTwArZ0V0X7G92xTz43BjvJ0pF
7UryAA9KZPzsnNAUehEHsCjLzVqSlOZe62iIk/+F+T3lYzdOgOtEtRIrUiTpPzOF
spm33eMGTd3UWOexgwB11AF5B0mvG5EgyDjNEvN3zDi93NKX1i7CKgEylBcZmYyO
ekrlL+Z67DJyjiiMUwYiCEFOJD+4vJxQuIgxHzC0myPfNMtPJgB5gcb8LgZy/YWT
8cfZ0oZWNu1BrzsWo2+1FBQm8kDqF2xov3h3Rb8sseQhMH9vMm2Vomfrimaux9Rx
xqNb0GcO0nL5aZllhrh8Y4yIJXi8tUucz4w4XLRrCp17x/0sPl2CY81uo1WStkG0
Fkxlu6pFg83ig01OiHepM7e7MZXcBfFHFwKj79n92TaqRM6YTpQbZNG9mymQIMnJ
hfjnw32Nn2XBUAb47RhW+is9xtz0euZ24YYgY44RuBKk1cSrJWy/IRdIhcrPOVN0
0ohgy1YV5o+rJoq9MxrlW763Ni1UXpA7KGGQVEC4M7d1QA3sULU4C6sLHNZ4ABRT
7TYgSE0q8yjxl+2D5v+b7Ukrqo/d63uy/LJuLAyA3JVxWAH1T/M+MPtwxemOXQZZ
qXjeCuMXFBtkQemHG4HA8VGnxDhzOIEbvxWNFVzzjZobto8zjlNJ+5AtQQM/g+e8
U0fabN71NR/VYLrrjPFRZzOoc3TEMUrgTLKCjvWHw5jsT5DuQBex0H2HQYMNJmI0
pT96pbWgocXrhAX7dX9p2qxWT1rjJqKKTLXkuxvMnluPmEYM1zCOskmS7giMBoT0
xZ01T0dEididyQ1MgX5faHuFfAS8JtZcN+4DQFsODEnF8ZUyEtUXD7fYC6QhZTme
Kc3T9i8n3ayB3Q1UxR/H7OvBkBJAN+H9aK1G6hEcuAtRiTcbZnXCpg59PXAdBYkN
gfqqHvwD0koTDmdgiNT+S2DNvBfWPKfxWP7G++tkpS7xqe40cFi3RBbZ75Xlujgh
QNViGyC7eYuFQTsumZsxwP+SGxFxdkPbnaHkJbOl/92r8DnMvRCjfK37qh5NoUA3
23z3UdwLJGClnfNa7glkQXe80B3h27bVh8p2d1WgDTxZZJxr2AAxBgc6/qW8i9Qe
jgCl55/89DoDdOL6iiL2mEUisFqIGCTJAuGZTyrQjzBAewNIsDRyEINjOIMQZY+J
l5bgAFLPvVh5ehkYWFvDDT4B9rQj84W9O7QEwyIMz9Bt3pm09plCYOml43rE9ydv
pLghOWnRiBvOQ0JMnZfqvat0xrVmkxHf9HNIH8YarepBT0otZIIl48L5NxI5GAhH
SVX+yArnVM9gme0m+katcdkM+YMaEj89gjy4QMVtp34PV1kXw5W6bqNjERW3GSvY
7zxeGIowEazZszsma4MIxzZF4WTPqda55IF23yB+ZR6pJ5GuUTlVnTq7sQDwstkz
x4cotZyq/iypFLSEJHvDpMiYSS7aUfeEKNxWCQbly3AtQSN5gd3Ac6lTh97dLDsf
WEE+QWlcBseW8gL9noy8hUffVR02trdJXHabEc/S+yCLYsS7DOvveoUZ371l/SYR
WLUZYk+W/KcuqCal63KuKANSlm2tLflSPKyO3gu8BL0CXVfVlNWUcjAPyB3Ylw74
QGpLWgsvq7YNdddoWCaJEBsBtCuiOgB3SIs8oG332LhRjlnLYS8Cur0omXgaKFjj
TjnRe6q36MfF0sYUl5I10tlhKTZdzYhFNr34kVUzAqtL9/tJ38YSBCZYrhgVRfjl
gWlDBakifBgydgMUyPhB0qI5wvOV1kjmy+/A2grO6sGvnhDhEUSYqPPaG09EB3T3
UtoPoy1Pn9skuKkR4zZABGliSpzC5QmIcNtzsklxPxtm0FwC0LMf6x+npA5rLhKw
Xci9UMrG0keXgy9R7hzf0ksVTvCXOhUODYRY0gXDpXpeALQcMadDfoKSGJOezMU2
DKr7J7lLMafWtJZWV4WAAHOvS/2Apc74nZ0wxZC+voQiTly0RgYPIGNNNCUauQSH
UUixSpIeedwAmN3CxAUAUjHeD1Nd2ghrVoDTLADQ7jsCScQDas1bE+OxyfRvvqrK
JDsc3B781ns0rrV881cwfq3stDXllxqoiMFsWwjCC7X19mNajQhlvhhJ+LyPffqC
A8u7izrF9b5A6Wlx+c7whPrgGgnutDaxzbfNkMFs1RkVeFZC2z0w8UEtOwvtAL4Z
lHVH3hDpwZxYNDNV1fNNM/iwhL7c0cV/U3WXToeb1eme1+Ys46VzHgzFRwMHdDWE
fqDNCJKTur+x7CuB2O4pOWfnTLGuv1JI7PQczj2ENciVufcT2KwdZjRwiGvoe0rm
Q+ESZyO5e7JfYOq/dn1Y6u4jsTthypBoNZ2GoFbcwL5Y2yL7cwdtf5RdX3XCwNOl
AmB5P25puuCVIBZjhZs4Gce7Nfgq6T8oeY72ZdcM4zxmLzPYpI+eOUgmo2hbtaK1
yZtd2HPEG63DW6AOVfJBu5zN0NO428q22eYkD0rhsX0pat1pqelwvzOfdNEJoxfj
yvcIRiqMzsJ9ro4q2glgQCdBb79iZ3lXPAEU2Gu006/gK7ubG7fZ5oPmG7oS605M
MaN8AJ3SWBWKCyD6WoXKhmaAVTI6bE93x0mM9eB9EIHnLesg+eidqQ53DaHSy5oO
lhBDncLfZcY186MkRRPQqR0FvOHgZHvq0nvOyJ+vL8WRuNVWz5IRFBWWsN7LoVoy
r5e8w4raf7XQL9FIwSDk6jysUJ9XmmeC4xj3avJytWEoODWXAqFtL7l8JR3rLjoY
5GzWFCD2DggAmUWEfxywNuAxr9nehxYsJAskPPZOz374JtIQYmRTCK+btrIMo5Xr
xvRhRF5RPQCKTfrymn6202qM7TaQkf6gR/on8rKO2V9LVH2jwKI1DperKPI/MW2c
HxU7FvvKnTwQ4suSjiTyaLpokbb+B+VEO4o/nSfHNUqKd/OHSyrpRWdJbsUUPEsL
pcg0x9HNVws6+wapLykpam741qcsz50kSHL0o0oMG0VzdZUyDfAjo9P/W9utxB3O
ifYAtl2oUODy9Kxt57lSqAZHwtF7nyrNGSD7mfU3RR7qWL91V4F1ber5ptMekWwB
+XHSvB4AqWLrCzPY0sxLF+9JckRo64+ZMQmhKZdXVZFpCyjyGlaFAbDUQxvbh0HV
jVYAi1u9pZKtu+nm10P3gMfEnJN2ACaTN6n1InCdEBu+NEusPzhk40ge3gUTUewB
QSJkjqBZvTEc5JoR79j0x/Qom5/Tgyl5O8S+onnbV40m0yWHqq0aHQLdvZZG89I3
Z145M/gym982SNwdOhBhBx2g+rRGclxPm2Hgq1FwoVXpyrN2YQfIsFbBkOARXqvV
VTI5iKhoDKVFmmyYqX9eDmT2cZMMIUap4gzmTGH69YUh2BiNJOFXdMaSAep81bh2
BhprHtAfWk6zsGhbup7HbytNbuc3bvhkbMAaWS5oCZBwdFDCD3IrY9WCJEvljIMB
q/qWDfwJq0ASdeWx2WHTX3kZqmI6euL0qeKvkkVMSJlzLt5uQvxAdfe6qoQJmCRq
ZBJY4Pb+z7LVXLrE1G1Ec+o9lCi7d+RUiHriJ0ok3TKfDA0QSMUSamrhPzFQyAHf
jPfzTexIBqhInF7hw9n0FfUqa6t4CDIz3lPg6K//4ZmHtvLMTYktOt2gKrAPVBn9
MiVdmF/k3aHphu3MFln1YdrfO3DPbFYAlNyvKGBnYeevNPzdnFOJNVBG+uGYgoTa
P0WdWrwWQSo5g8rqUqpEqrbt3ue2IPbbjSZweJXoqB/2EOmoJWnyMXE91rXwcx6o
Y4MtwUmojZrTAS5eH/c8A7x4Ff+UuyOqsfMhRkjrI6f8tyElLY6n6VsIfzkdLFQh
mYQz2i2y6iT8Nz/EkEMctJxDVeTUAHfz5b/O8MIRgpvrj2mTlvGFLi8/ewWYm9PO
PFUIEYaZ4R8Cs3vgX5hLU46WO66y5rCtiCmB2v9DGQq9NnQg3S4GfUswDh9OyyQt
QeiSG1kspDotj7ahw3RaT8uNLILrkmXCdvO2GXdRn3PD8eTexOeydKhNvqpwJl0/
MmZPZd+9C4iluhP69h/ZIckGLPcr3UH7H5Iz7elLKUBuKdOQ9Ln02GwLU3IAq+55
lgEDtH1LxkV/vX8bJBmzIJP7d4X0oZKjlHPNwnzzsHeooRijgF7TA4Kmh+HCoL9z
ooo1Pxxavi27p07YMqKgnd0aoE7qqhyiGBzGHyVQUon8MOvF+D9xeKb2nymH43dj
PFAurpci3HAhSSpY5XmbmoZ2y0pXMRp3lQgflQLxviMr9XMNQGKhJDeWbnl5dPO+
qvuBnhpD+2m992VYRP0HQl34YFnjwysHtosZ/0RedtNHSvPJ3PPpFy7zB15ipoPt
WCVK5e1u84uzoUB00BbrZDnqb1uib3BAktxJccjZuByY4MGDykAHjJt5bFKsenE0
kHM8mWW8Qz0r1VEv02U+mETMe5kKcM6XQjDMFZaF+wLjnaYgNLsNE/a4iFK0Wnn7
eXytsn24FyxRi14TrgZJptSmrpR0by65uVKm4IycX4V7oo42ZCoVt5wgT+XDN6nx
GKUb4pKb4OVjtZ6lrQfIiUHA0gMGqAMGfdJHDc4RtjjNH62kzOHDf1/fUCvIfrQz
eM0Vgq47D2xwlgRfPhjAA0C6EVISgaxdFlzNPikmyMhoQi+x8jHKVWsxIZve28Jo
IR8rxq5FtoKo0+2QIbIGWbRwyQmGlEGzpOkWVCyV2Ag3t3TZyl0wYXmE05hLVmj8
lC2PbxjVqmEgK5xS14yMH946Nnq3q47NDjH+xsoe2AhWCdhof1NIthv93h3apvyy
XmZgIgTQKjGQD+KxFy6o9juOCuWm9tmKfxr3b06gTXjFfenS7cTpVrYH0RqXrLi6
xkSmUlKJ4cuk9Is5DxLG2EAPfD4XOkjdTLnBbHHnm7LocOo7EdHBs8C2ATNCP3nY
/l1TSIVB6Dp88VRIKFLQL+oJqRSimQYiQbsgEUTBef4ECYWBr400NvJkxjgrpous
1WNYHaeGxUwHI+7+hwoQYxTgiX/ldffvNPYqcGHoTk7m8D8SKKYa6KQ65CByYxHe
O+DkmYqxMFH6nRUpPaMk2Q1BVBHFxMNml2uv2I9iVsV1tFInH0zJnXKapj2SeyVT
VSqHynW+N67r+l45DorcN03LMD65jTlNSli0QZO5OyVtfI8tcXcZe6ND7ootdmTM
mzOMQRHOQQ3eMjIyU8dn0jaO09cpDXxf1Id2KF+zH7LBK/tRdrrLzlH1HawCaQLV
EykkLR3STOFTtkR0+cvhn1q3trCu1nOWF2jrtwkn4fwtOgKTBwPCNQkSm4DxZpEV
SmJvIjKBgDUQxHGA9NBoM+zR8J2Sq2CNYqlcz3Oqq1dWOFTdz4H2jPmWddP7fY5r
zgxBVaMQnFpCMy9VWCmPemYDIkRX94UkWCqROi+eWVV9o8dzDBoFLYbHh04JVR+t
NH4V2jcy0CLmZz2NRmlN5NUMg/3MEetig6HeAVWV/CiY5HH+xO5EcetkBP+M9sRV
pliqJkHjvxJqIXLhF8zWQ/rDAwUPHDkx6qf2MbT8olW8U85M3VWh0kJ2djHFyduM
icILP2pljFubFOYr5HANz14A8NwhkHkHHaxtRq1gmH6V8tVNp+55KfBL4pSVyRes
DmdTTxIDPqNPpRy4L/zQhhZNAiVBRXlfzpl6B73UoMRaw7C4GOU26ihvaJCNwP/k
mrSVyWanupZKXo1Rkz7OBac4HAy07RTtgQDV0e3NcOBT5Zib5HNAUl/R5rV0Hkp8
fzONNP5m4Lqk3JeiNsm8YRYPST4OnvLk9dYi12ocL2eUluyNcmlyjMGk6uyMdvck
+ovqEHmPuQWkOGxiw7yWqtUVA6aZfllMmgVZ2fUizdkVXODZD4mSFsSipxXZma3I
QBvxPTPPkT4kHtnqtLJUwl79rqp7a1mwa3xzOQNqoEgqIAHPz0O1/kVwpP2nP3Bm
RO30LXUg8KJggDIvcz3ch3A4pFu2N+64182wHesN3LNjbxMKWpnroZxkWHJ2yuXZ
Izy9s6KzRLb9djOrcmFx5U+HPnKXzXYtHDe66e3pzJtVfQFE/cQiF5doOKbstufA
XhuWBVTdc6XH/VeY3TFCorbC5n24/e7cPkq1lEri2U98+gPsnFJAcTX0PUjYJvkj
yzyCRZQylqh64nU9lAwlEgEHdhLVhQJMJTy+nZ479Z+aGMt0HDcX2DeY6JTWd/lh
Zyb18zu+Bg0TIR5flsh9/YxXltMO4ISaYQjkFxZjRD6VpAkrshC86UZOkFqFUgA1
BExwagKl2IPTXB9e1PsMEMXgPGwxGutHtflpjbCOjDOhUVRordZIwMzpASjNKQcw
dXLVnN0OG8UwUSdBKmEvlxIusLnTsWhFOjS0iJg9mLoNioO1QtPDDzrXPernOVMb
dJxEn97gptrsx/HV0zKLb+ejFcVQTxD4p8lhTc0+UJEtvaH//6I50fTO5/j/GhTV
aHTxz7UBksx6L5V2ZEcYlCptPdC7XlGDVw+dhnfLTbLOHiNLiVErtoOJeoK7lD2a
HV/6oJPiNfXRvMoZXNOj6QXt0mcFMjwUP1Stfj4TbjjomaJa4ex2+92w2V95Cx+J
bMGdSS44dln2aDWX8AU+/BplkPtIJmbGEEyXhdJzLhpsNT80r/ptkmelJU1BePNH
y6NZFggaCwODSDq61ieIYP848xahx6vmIOkGrst7wJjrPC7VjtG9gOG/kMdEUz4M
j+O2mzWuXLgPSt2+PhBhpCdvKLrFYviI2sy52fje5l7xBFr3RFtGyo3Eiokx87II
cVwXVtwu9NUaHscQgPaAes6LV2f2fcWGOs/YzAygx4Lcs+VztKgINuYpXUipXAr1
ybj8EsB1MR7fUYIum/3/i1ouarsgAqWmBQAG0Avk3uurIt+Knai/lZf2rqs9xdxB
Bs2w4BBtLtMJ6bQKhAihUSD321UK4fP4DgVrL1pLj+yHOu5xd45niKd3LXxwU3BS
m0LvGCORqz6U+rE3It5IwJFW/9jcj7NcMTETr1kNduakqJJBZqfIue1IMj0ggymH
ncJ9uvReT4KJj8bW/hczUCpYiIMlYsgS16/ljSEvwfPEK9s9DzIVh5+UTZzQYNsr
vY5O4MNOn9J2mdWrSxuYFcy9iK0RiJInf8OLGbfX5179lHeys5BE4T4VlXPBpief
wEclSxrYJucSQRummzGsfyCrv3zy6L5sXqt0qWvumSb4AvJYk90WAddtkjFpNGQR
B9mZiVpL4/u9KySV7mhk8CdmftJvn66BQyOrcqXXstjHvMXM737YtyHbpzoGg3X/
OUZZxupWB6ab3vby4QYHjKHDwsD71E75qplz/dNSl6VY/wrE4c7B+zAMhGbRyG/x
bmSbgVG7Sz4XpQza/eOBxdwIN+XDa4VS2jJDKCRaYm2GlpvtpqeVM7fHtsS7yqKo
FgPH/SrfwcHjCvnCmefB9RFs1tHrq3wxZrfuLH89W+dgpjUzdO5MhtaGk/y94YR1
PRPgCj7LCIe9yGJYagca/bBuev3S71vDYyn4ovdwDuT7iTclB+j4ErTJ/+sXICUK
gn9GbrIETLVlnGcsKhIn+C9pX2dW1PidX2r6p+Gx4wCMUuKm7phk3GfJQZI37Nap
gXc7I1ymvzcvt4vmgzmnIJb9O8ePofF9PdPK7DlZ7JFJ5OUqyHdZhx8v7CriDTUh
PfMtZDzEHvQqs0Q57DdKC2mJlg0oOD1A3zjiwdq0DST0vIjKQ1YwriGvoo732A7H
sTAtPRyusLRR7OgfvuauDkrrNsYzaGBK7Qm92N+Rg2fG9kASxgTXyDfzy7kiLZO9
Jmde4Vpt3FWcomwFCGWNNjzM1Xc0t06q1ps1iIl3bTB/c4CG4QcxkjOjJmvyMlZt
ZQ6kjHlMkTXFqfKiNSBM203r8OfHOi7E56RWv/BVDytxKVPrnE30dbob5+hFnSUk
EmIPxN446MTgbat0G68rOGrrGqQlsJkI2EZX6Iwl9LfQ/qfaOGxML1WwTRZMaqgz
BKnexdpBsPsGiDnlD8sUy2aN2C/8wpw7cPQKxMmMXWNIj9ELp7puqYnEYjg02/oB
e5oTo1xAOEHtNljtprRyZOP+IPl8u9DuAt8KM/x0ZzfcyzM6vsAEyS8C8yv2cwKe
BA+1Hj36X+mGPbXEkhJ07b3ooDhtNxoxOBep8dPjNJ6xCh4DydjE4fGwofjnrjDz
0us54uEOGwqyBk6xZXpo1dXLSTPQFluiWlBSa+l1u3ddo33BM7k7wC1mIiVLrJ8J
QAKdaV6oNKLufuqQHfjblATAvTo0zf+rHjeuj1EPLd+wGaY4Csz2jVtl177MZeJw
NO9B0bC7e7k5Xj4SPd+jbUM8VXcjDg95hsg6B/BXzUzTdUluB2Dt93tN8eAb7F9U
AtSgDjQRig6MC8198h+K94rmVv8i1wmTozClRIRE4MgIgN5L8bZ4aanxz14D/qru
lDfphu7v4pkgb46tnizmbEjLoCle/zKSn7FupY6pgC/TAS0KFchaDA2A9kXzwjNs
XuIttHrZ68khRkyrWMC1Eir4TOAiRxB05cxEcORrzzYM9nM1/MytYzo1vqIdG8+j
mTBTVi+z0dguuuoE7QfXLl0iLmBQK2SqTaf+1NeJtX2KpktwOdXMJGKL3h5iCRVk
oSeTBLmoW7iTMx8LAk6xitWoU359oSn7NITgdWCn/r/c7vGSFtfv5HXRiFoZmA3G
TfvoEQitaVHjyXb51CMkUnLEbbBvab1vUHIMrE3SUsdx0AA48+SkwQBmmA8rhGQc
1vkenZrONF2W9/CbBr91ZixiXNJRq570iAst0vGtYsRe6oZBLT+FirVDDxXSuFUh
evwQz1T94RxaQQ1VYjHJDWFVgOGMKLwTEofMobRP6HTLJUqmxC9+ryU8sMWEFJoi
1FVBZepsZIMPvaesUtKjb40OdP/M2xgMepNbalfB2fBofiuvZWz/xdOBCbrYSNME
C2iKnFZ514mcF4H/2jUi+2up+Mg5oofmM614a5+josqB3ufzxIzLMIUZIyO3mRPl
RYrOpSpcasV1exP8WabL3INS1jbo8GW2urh5B1tt9JZrBZWwsKy9y8BOXwlAB3io
eWA7Kf6bG+6g5bZEJlhXiVvXqz/zuaQfNOXNkeuTrk+i0a5ljYAXo/fZfY5fqydM
rYoXgGOWNV8UPCAoRvc/0es+pNGS1/jUqW5uhi7LePrhSqxxo7HMMm8fWThPLhQG
0PVGDhUHZCfYzW03JdHmyQI/QQhyNjShv4qTwGv3In2847/Jn7Vz5wt7o4guBGVk
J82458ICbYCscgNcVByZ6lvHtu4cR43xaV2tr19irMpKfokI/ZvqRuAU1WRHjIY6
YOcpRdYzq15Y5Pf6BRcqdNywUTCqohAXmyES6RmG1bS2JmtZa35M+3prpXWz1/E/
TdZCX6HTessWi5EtMuv8NUmYk2MeMpXTpf/eMSOHOIQbQEdEtiPfTtTX/ugk99TN
Vsr0kbLXYHl/S9TkRCSiZBNJon4lCGNDo2fKHGBeifSvPdJI6DpFhKeXO3jGPp4S
T0Zx/EmjO7pb6ZwiE25NrXQbfz+bIhIv7ezzdwqQ9sy/Y7AmK4bVcoW4aydfpRUd
uWMMFPeEOpN3vSYwIq7scQEW8/pbIDGHHo/Nc4GVwR9nzs1WgLSY08j5CH2cde0R
BjXuGzwGQiKbfbxffL3uh9UGv0DijAvSROl/jioM3tQB1RsZqniXzcOCgQIOwBcp
0INTHCx8PBH3nYrR5fl1aVp8HN/JrsYpu8n27V2QreArsbmpeQ8vjyxpYiH3LgKN
qxPNkLzJR48liXeXNu+g5jCWpAfM6HTOESHkjGMIiGE0ndtSfE6yFb00uUNYw6EQ
Doyc5JarbWvJWSbPGwdOpD3hIr/KY8RqHhHlKKHFxKmcVsLVLMkuysfy5xOajkP6
XMNQqL1gggp7FEnbtIo5ZvWXfQidRilR10AeUlvTRbOnyFHr8K5gYzBWaTv0vKOH
PBp3o20OmO0kJi1rqwBGicVi8oBDYMgL/Z2GQHwAlgkiTY0AoulHvLPuACPvV/wA
RQytE290fUHRrDWKtb0Kjpk/d489F3meovtebyQ09c+yXnyNWdQfPo/JrsH5lVPF
cOI2pXGk2keexBpUbrJMCAcTJKsR023bvKG+cCuO3isqIwnM/hpk/RWtt56GrwDY
rIqNgfEcw7TJS0KVp8RK9oiZacm8eXSIiZB74q8jn3DBdD67dYUmLssNMeXgkOq0
NFIrBnuDxwfrQptbfK3Vlkphwy+HiFxIIS7Wpy2Ty7VDR26HoxxYpUOhV5bhVQCV
kTgCUaKcRXxN5KaVoHMEy/WkIHnsDhrSmjVoWg9sYEo8j9UIeeGlVnbVReHlC/cm
wzrVyVPEMsO/G3kmpUhsILa25c0vSp/ySQqhjYlqCH0j1LlcgX46RWpOh+6tukJN
Sla4AKug6kD53Tl9wYip6rOAhETPhPAgHjdjK9MxQ1ltgWE2qCTvHbF/q9ET/p12
voQ1ZvzW73i/3z8RZZyF69ezsVzZklk7ryJ3yRE7j7jy0ex79qs4WVA4BVIG1Qtg
v6kpMi7ze4akkZu83QaZU8OjuCXydcs50lFkLadfze3MvewzvD/SBIP04b5jr2HV
StWyLrZKWhfSPawe6YxYFg95bNcaPWSkZTL51bB11zg9tN6eJQHcuA5kSl7+nRwa
Idc3Y003+9IaSEN/dJKonJWAx9/hWL1SKahldHe4eDhlF3AZoivvYC1D/ry9qipT
0fcLVLlvO9EjriLyGKjRbhFfvYLHf/M5n8T5yi75CTRu0vuYM3BDYrV5LqWir7fb
J9jGJGA/JvnVVth9njkn8LD9o26De+/XLLGwvlATGIYnD3DK1zK2+mzZJriZ+HNX
xX1aTbHuLJUJAgiiNO5f6WuLgfla7KbgpBuUx57d+K14ISHA/IXuBvA0I512HXDt
7m0UmKkmfM689AW/ij9FsHS6HDYN05lIMtHyk/lTxwSb8/yKRtDWdvu7DEhuWUnT
BTIMBb02nFI4xGgrcW2FrMA8C0eIaScmD3/+YWwRzk6nZd2xuBBwbOS24Oga0llh
srFPdCP20qgOkcNpQW+UoXa0cQQzhnwldBO35D/zR/xe4bdRPzLkmKAkJaOOd2tC
RclJNYIzF4ah7Uiw1M4b1T1p4TOueugSYchB8HK05yY9W4hVw2jTLruLwjO9d4C9
CyckBJ8mA3yhMU6DCJHjHwHIiFvJeNh05ZNyjgzrHEBSA66T6/Bz417GAo0NOmG4
sj2nMuMTzrSDrqkAZa2OO3AbVGwX6QWBjTZEeQp+JIbS4Bqe0kJF6Qu36wDFz67u
iqjIPPI65BbjikjkmuYTsLoDXqzj5HgF8vFZ4lmezsqGGBFMtNzLSpcAmkvwpaBS
9IkKzqK1/UopWFhzB+btTypL1Rir2sOsj3m2m74gi9e0nBcKwPdIX87kGcm/xtCI
vr3NF6dzm/mdyY9O9QPkRAskgFUInmTrfXt7wH0zH2GCGST26OaZc3hs9KkfdCqg
1JJsqDlhY7d8kKWjqh2ocxKE3CtTRQMfRJm5Xjpji6phhuf4NIB3kHuWOBScTYH3
tTQIXSn4j5mQuJGvxUDOd5Ow7n6HpR6ZKJ4YdGmXueo08PnGMdWsHz9LUXvjyo6n
v985muJ0/2bLCOUHiWLNmSiR5Uoyd6PNdDeDYLmcE1fzZryxDm3C9ZIoDhcHVZS1
HLqxfU+xBh3Pp9kwm5R70pgFiWtZl1c0KdHjjTwMWaNSxdLiJbHPfeZy1SQvsxAQ
M7PVWrK27VCBskYjGRuIWMys7GXF3wWM4J+lp7250cghu0KkHNFfY2w1yTkt3omu
OES6prc8w6FHcdroB5aCcBzR8f5LAarszLDDgrqvZ7hT8be+24ZfAE1xp8BOv5IB
Q4+V/tj7Uo7gK/xEUVFeWKbofilSwh3GwGN2xB7MkZMc0guCt3nxzarlB2Manc3e
FpES1ZYlDsxRtUFGC1qkwuH0VHYDD5umn9+AgbpFAc3cYb9DmPUARE3W69uzPu5O
WODghPB0TNNRCnO+6Xlnh6bxoZQehUPnhw/E3Pf7Tz/gZRcXEdKUNNZ4nkC1rzwB
FXnbMZPxu1WPoSg3pVri13jfLs8610FjXabmxqUFcd/SwqapRJg7LsBSDbuJ2Lpb
QcXg54VBfFv/ROCxDYtwfC+w/1GBKsg6WkBakgLBUrlVNr8GY7yW48chXFiqo2AI
9TXM/TChKC/9ylfJxdka6q/fc3inzH3kJEMeQI/M4nd/US9CiDyM5RzcG+wgweEr
zPOyRvaONlXqR4cQtqGoxALB8R4vzSjemnjnG4XS1+RsDOLQ92RziwiebptmJt0m
4ypf7JHn7GHo7QoVNaz1tbn7H7Z047tuPJdXX89VtASk2xlX+2eaDsoUnnwBLLkx
SUAjpK/t3zeetO9aQzI0SCmTBZdL+f0GJddQLdH7ptQBaWCEk95eNfNLLdlURq0G
RtxpyzkQaj7JYrR6kLb4fHo6HkmHm3BIbo5wY9k/LsOP1H48G/5Sz3CP5SQtwosp
u4xpN+uq+93Fk9lVXixyrTma+qtou0/8jnKhS82+wFbcXqtah7THM/z2ZpN3yb90
2nkGK21cjNRaNe70++31yi+Q1KaFlqcTQd/xnWsr4x0jQGys6XOjKkTG0/0I3ueb
3BFbs2+C//i5KKK4kZcYAxwgQuqTcs4bdr6acUFQPrO30WTrxa8EzPnUsIoKn8mX
d0n2DkkmPZXaj9ZFi2Dk2+p3w5U7th449SPvE/r+8x77rASoV8X5MIcXP2fGE/CJ
DDAmUsmKfWx+W9NET0pB/7iM6VumSShEKnrqRaNQCIrId7sEpVPU6WyULHWBuugY
uViVJvAL1IoGef9lpnf6nqAlzCHF3G/jdK0qnlW/c3TGl5tH7fE7UOMDgiO+vj2M
sxNSiWjb8Zo/wGB+DcVWKGsRcTGSBOJZIuWs3oJI7Yf6K1dQr5i6j0tcxh+yBkzg
r1uEGxgu4HtzpXP/SreBQ9f8VwCLFHqzKfexUhPZCrH0kTxnKJezKVcUrmJ2AL1m
0EyTa9mVBHre6FkgRPcnmC4obroCTrSSx2fikx32LK9uT0HFiTSF/Z0OAk/0vTvX
fQ/hsJ9m5+PzvD10Mr32ygF/pb8Q9JgpgqfG2Oirq5nlMatHrWnV//P0Fu/DikOF
4A/Fo4NwJ1qcR0D2cpvo/j1NMJRrSGrNBRzDRER6v0G8DjbnvFh997R9QPRXNRiv
if6Dycna5wRbmFzgiYlLHmRmk1eo765YzsyoA/t+OIBWDasXmp8iImQilkBXuzpQ
v0eBWWobCtGx54hJReZmteQ0fjjbIWXVGxrMF6ThluTwkS6hilnvvurSLFSEagXm
zdCQSWU6ZTz35eMsexXsjOffugcv9J/1mTMYuAlU2/s3vqRK7zEzJNlJMMqQFlS+
dLlSStRNgIy4LLw6e7rbYmG4DTcsjUGExRRdrpMos7pVMO3ENFTfUgbt+JEYqPQy
bWjrT8X7JAYVBFrK98dLIFKOLi2ZAZctY+eEDfKRWK2iWFk6zgy7P7cCYKXRgnMN
sP8Up0rF+5l2FshMIN6lmRPSrrE+QovjTWQNJ6qWzyWNjAvXFZ5pAPWG7/BCAb0b
pgtYeB1So22Klr5uT1tOUhd6ST9p4GQVb2XXwEbHR9iGRouZR0/imkT3s3bgGhi9
2VqqH4mhC60QZzOmt8bDK4B+6hl+KtoqN+hHHCnUNRflHgGWxJQ9QL14DPWqmxiy
kZ3FMyZXG0UVTQupkqTbFVd3lVLNMvqKZXul3hAbC9nnctkjqpz5LRoTJhT5/KOJ
u/IMstqPROXPn7u2owbLYAkejiZJ+efpIDxmh5GgEu62vOFNvljCEsUiBXgYUkpO
kCnlYCRV+ue2kUPiQuz6kW8sdHBgvshfKgBygYVc/33tEe5xMGhZ/teVEXdCg3LW
3M92mvS5yFHrnHhMe6KCy7M+y1Z2W9asxS056tLhvtf1PiA3gyxFUqBDLmhJ0DTL
FrhPzigB4A8Z6GEsMeoygV8Bskq1WGF4bNtw/CGNai+Y0+BQ/+g0CIhH0kUeWDRx
4thU9wnzOHi156TzJtovtvUJZY6vrcuGhZgrXCbgI+XsD16MnedTjXBfuLV9KsOX
WDNBgQFMHsCYJh+fRz4NS/i2pB22ZFun55X+8Esl0T+WMCYaL8GC+axzGwzO6AmO
Oihhyc9pkvplwZmf//k553GFx5JwTh3m5wYRmRU0OCNRZawvcQcRdX28SX+b4sQx
hHJ1Pn040a8dd2AFjYpQ++VOJHEMLvLc0S6Bjztj4buGC1UoEkVbpb9uTVFUzMeS
TeGSCOAy9vI7QT/aAPHszifoBLlB2PaBK4rrEBPzeyAogjNRnIgdBWenK+D6DLnV
Gvd2oTbOz0FJba8cqsRDYeILOpdK5EsdIYy82cvlZx7ne+Uyke7JlBtEXB/eyYEU
4CSS89DeUsC7svJpJ/7+gT/NILjkIIiLhZ3nfKLLXpOpDDPE61UHCFE9zo+HdyBG
lMABvh3mVKTVPGBAJw4k8g3V9HBDgf2oZJnzIdd3k6CXz4ERXoQFU7hl8ZJqRpom
shqt+LxLXkFtY0wADVArKuoiuONiziJt24OMqrG5iHbFVUx9s3EUD87wA3rKpCQ+
5XRk6p+cAaoelwJ++S3MC5hSi9FaDK79oAXNyvs+r1zADhc80uci9vWXMmuWPouw
Ow6HisJbX/ifF9T7sqTAL2hp5rihwM0c5BDkAUq+n8kjoyf3sW8ZrxpOyK1DyPrl
RIIu+fOoab4+RsQ3kyxseNfE6BwWMqtCzmo90MRCx/mYQ9hU3fvcXPatCFTPT33h
lTKNJ4DpHDHGrH0rgiQLNUTQLdflZgfqCysqCePXk61cGqyEJqt9Pyl/7ywDD5VB
6yw6YpMyEd3S2owtQyS2IXvKzAXkhFGQ9tqhGaMbSqXSm0BRyLrfZz6fnIZUFsi9
eVYvHvA/tPRhtUbVT/6U9FHU/WvZ0TzvRDLFs0PA5XfYjNkU4Iu8Cc6X1ZekveWS
4sRl4x4Rw6aZrrfminjhKRljNKY5q7MOKR56YuOPQGRkvsoS7X8T+CEbHgoHLfUk
bBA8PdMLI27ZtI+xMr4zIQUTwPrfrJsj0vo45e4Q0SvtI6YR7oD8w9ya9NO+MAmk
1hADozT4mkJx8zj4uTT5dmJTR161yXU3gN0+U4zL4byT/22H/mL5z8C0foKa6nF3
d0JR/rJxLoTg6vNOE1dQ9EXVKdQ3MbgSz65owworIXjkwEAVVtwXboF1Mly+E+Ou
Ef5BI85A9zBB0HF8xHk7DMcAsm58AdS/cf8b46L8D1uDtCr11jZnYrCkL0UAHa3U
gpGmK4+3y/a6nqk+AW87MR5EMY6javizR3Lux4p2OsAMpzu+cxoN/qvHkRTit6Pn
OYEbxMbvZyuIM0KiQfDsZejT6oluDytaZy0ZNhDgVrgTpDoYAV9r23HVjHvxCbOr
ewLqXcEuAJk/pvoyHBqM3wY8XY8+gEz+rCKncG7ne8R7QIIZYUOxiM8JSe4wjFj4
l7NUdc2+GC414S6IraGA2P8oXQcabfDKgy0hhI/u6fUkNqT79ef5asDTDE9W8NH8
kAGd/bHYFElskCCABOJnQXAbaIMiEx57lSC8hmZfDLAhHej7GSi4KIoGs/Bf07it
Qs/R8Hk4m41mQe+5nNRh/B4U1ysRTLKEPW4/n/3dPvZ20gBDbPLCAycGxE8QMokT
Sdmcbl+h/oR8s93lfGswxshEae5EgcW09ibfiNzU84THYEuE5Y8x/CKbFSDYuoIT
PYvPjDKfWK4bKlo5vsiTjnvz0xGKs2+aPF40PLj4AP5t2PTnmDGB8vCeptzq5xMZ
Qvsp+QWQ9OlI5YxAPByZX6HMr92Vb+eD+P4QqdpLQ63NHrrxpYaTsCTtVS+xsCVX
8dHccozTwWGB5BSGDaQ7H5g47u7Q1CE3yvLfZEKKwaIh0nIXH3sijmuYf3hGua+k
k9Ehk0qXnOyXq0N6YBbljFJ99pMzLtqDJQeOA/hOxDmBNB9rGnXKYW3ycDWOH/3u
5CNH/AUvMVIY4mrhY0bNfWl+zqkTwJghnbL2++R6XXXJcVioKtsXr1gyb9Bzld11
pg7A2Xoi8rQ3HVgvjxpaAiJwsVNo/pLW6Pnm2QFcofYUJiaKoUotMnhu8morFRf3
6QizHd4IKZge9ve/EhlMAPV/tam9UCjtssN0pPLEOOqDKlJoc3VcW0sxgFBgCknd
PdlF/YPhFvecmuvkedFxLokrzXdw4O0YKIENmBOR1jUSM7cSmVBsC7oV6l2SXk3h
U7Fbn+I27J5DdDK5h3OR0m+DjfZ8eHTRHqM2svfdpZ2+zVrnRFOVkkALxrdEH++w
p1HbJjimcSEhSpVTEGhMXMqj7DhNR6kQDCABQew5j6eMgDa5bi88wXsiYLIHJQtG
7jHWsYE841ze5znHGuLppJaO3kkMdZNAStpy88mKMUS3g7he42UCO67dJs5hkure
O82htjziBUKnSZ44uXVRxyZxPC/UzsvxbAUyWNL3hFpPtPBMvMIozM1k0eehEhcq
UfuZhN0GJXHTqcl769TZKY0dFJUjLZNRtY21JbKRYrNzQcdBsVHmrL7lY94gi/do
z+L2H7/Cu/jUtPX7SgJIybuOWDxEBLJpP431ZihjJI7NZvOElL2LWeizLSt0Y/cJ
wCod0e75+k/La1h2QMBAfAMzbO+IbvwyLaABKkUvRCa5ZZahiKg7CF3RbEIx+k5B
f3GgqJaFdyg5fcmDNW1OWBNB+da6lsPI+WUgzGUAUIlOO6XIbuAMOToWwZ/kSgHp
/VRf6RaIIMiXZcVDwN3qqln584PBElc8/oCs+xmMWziwOLsGdETu4/6RUw9VIKKD
4+vGg/Z9E1LVxdAnWfDO+OH6jKBZFXl8ZbbJSAa5KNwPSU2n7SX3vx5WoSOypsGP
oyYnkDFdYM/UMLekBjusH78d9XL/V81PK5ilD1lGP9Hkm92LLLTc714BAyTSRLUq
oc7t/cLUPwDJJN/ujfKdBE4+d+Xwdcechi2TnXcVxXWAOnB6gMCRJpacSNYn4dmF
xExrOZUJpMyfH65YcP2QUDkxdNkGmLfPLH6JbtqGPmOwnDJewPt54UYe54kNPnAi
wuB+UYBuY612BmE6sHgltjTdr8pmK08mDFeklASwBhNEycb31GG5bCeZG1WAz6Bl
aBmio6siY/9VgCzNMpVsJADGIm7/fMn3q+gLBejQaXkcX7pNZy1zyGD20ZHcvPzi
5stPCSjJax1XTMb9ux+41BVhVyD3Oxc1/kIkFbshN95nIHGGmigEpVSsRmdW51bz
YwU4c4Y3jD60BAYU9P8VLPy+qZSLRzgQLwG3+2KHF902ttGpL0+kyndtbggK58Ce
kpSzRlx/QBog0vMYjzNnM0azBfqrMOf6kVvWyMebBn2KysVkavDCb9nx66wTeZLw
1OZdIwz68l75qaBpVHuVVhh33UZtBPchUWAjGiNJtRfpPFKy/etu7oKWmcrBSndk
SlV+npZBwLyxZD5wQJArKNVPFW59nCtbZU/qQ1XNlwN8N+YJnJq2jdijMa8nfzEt
UT1j/7p2xbB6DgTfJlw+JPcKCdFmpCXpvM8C8dtDH/mFL2K6a19g8Q8BM/uTLZME
OrrT6NGSQ1bkswwaRoV9ioNuQuLs6b13S/PdKYiZJ0AbxLxtUAb+MGp/k4INDKsS
432JQ7+YgTliMingfDJbPSyLNWyJnPWeXjDn+z5I2WKJ8APnJvVEchtvvlnFGnDI
JW7X8CISaWFr4C62TTyYfLy7B4hIqFKctvXkPZM6n4rdj9NsVvgOizokRViUSMF1
b37D3VXNmzJad8atQJrCXpIVMjBC9xng8EhnEg2uA6zuMT1/utOvJ2zBCBruioZm
ZN7gr/SsxU5g0g/ba7ZTkPEDB9LMBL07u7viYmz5gyCvEMMngpqD197sFrX9F3A6
tpyzy9zCl8OSRQVNxsxoaQyoFfNiEQnKzhGojBc7OZukcP9g1h/IKzYO3J/fChFZ
GNmisx2mwis1gn4Q5McDcetr8PyP+97JXBMTwClqU0yXITIqNEggS5pZRxzK0NBg
nEOEHxM4WNAu+MNz0xcQiQtTuaZEbXrGqujCrjM58RchJbX0kUBTJ0epIByRub91
DAGVQES63gxhKwBR5UC8ymwdzjKFSGQccwG9CSdGLnuvn8qFJJRNr3phq6ZU2JSj
b8FuRPs7SsrOyKEzJcsIElvDvZei1TnYv0o7xRw2T8bPw90AJ2YejeXCTHvVWZqe
MDsQXdtmfvuaEE0eYCxGXm3lHfGQCZn6Viy2Mxumn6P31FxC9m+OhKxNC9wafGaV
0rnWSyLUhEgaxYaLLqMa2DLPzawEVTGvWKGzIvXpHUNSli+ctMneidynZv2Csaoe
yeTA4kl/LTo1Q94ScRvL3x86QQEO4tCnHjCc6s6COptKPhTZeFBYupIi1Tg1nRIL
mC1T0sGJG8Dk2iY9lWlK0jPW1D3q4RZoQAdsg4q0EFT++eNQpGdDwlDhISuPJ1xD
Cd0Ug09k6n9fXoctLGiWwJfHmtG/JMPEWJmk8XFQaaJs9YFTskfwc5ySTs2wHbWj
PwzspJCNmMYzkf3wtrYVI8Pk1ZSH0oKKl3yFx9e6Ewrua3MjzO4y9Fjgm49DlzBX
+Zaj1c5Owx5oOXNMoik4JbpzgnhMnv64ZRuAoqQfarz4lS4eU3PiKCl2V4R+Afdd
g/hps+A0kAAFKC+PxFUSuDQIj/r+OT44ctKtrBnQ72nE4JdtWgCJNhkEGif+e5cx
wbM4GXsIdgtAJRPWil4SVMpslnn7EpOIqUE6fq7iKuSKXRk8XgalaGRD7y8G6Yd/
deP7DwKdGkogYpUuMaP8wJwe1jyIQT715WRYUZmiJBBD7zIuUFz2AF2uXrbI3DE/
ExeH9DBGRbuNnuJQx+25g/FgimDVEbFWybp3TZ0B60B8FZqsoHVLK6lkVLZDk45O
mcV+K8QllHbsZP9enfE44CNphLWqVKkYllFmkNqn6MyE2zJvC0+k2kaeL+44DbX6
D+Ab97MRFZfdjYwtCGIfI6mC3FRUjF36c2GHWTIQM33rkPsn5UM57Yhdjh96hLld
oisb188gUlqppSwkn4zVquHnQidn2XKomKPNGCXsu+u6t3RNoJ99pKrn9Hx00Gg2
slFnqIWhJh+2gx2p1xsMhLHRs5NgvOAXN8JkEqxTE6Xh07irPLL1wDAt4T6SuGxD
Gn7M+iPFOEo6gIH7n27E9C86ahvvKOatzrM1pnBpa0lgn0EElWrmlKleKhTyiASM
GF/EGY+wy8kgxV1MfbCM0Z8c2fxtj4yHqntOaKCiN1c+GF5rIdYo3nlFMd5h8F2C
kuiNCSBdYm+hGbK6TG40j268gJVJyzaRWe43s7t4h45lEiVWXDayFjP5S5E/KoiE
O9eMU57OPHVfGfmfqI0vzYmJpkf4L7BiS7H+gofLF9DwPt3Nt7kkd31lMscq0jiQ
OHtoUxFaGwqkydfX21Ap1fcjungKljsa5AHa9klxwrFHXbg8tIOzKY/uiZwqw61W
yFIVXnQPFzx3s4ih7RUsD4tpf5r04UH3w1BRxDoEmgSRGCxbW8eMAyeKXja4Inz1
NufglzfXOkek9whq5Wmzf8vWPy/qQN2CcBnjDQFGumrUJkhWWdXD5PPqux25X/38
GADTzRr1cyljjOCSWQVD/HMhVSCpVFYgRN7iu18G12N8CmSWh5kxT/KYHWF4lpWr
GwH8mHRKeo8y9qZ5txHbvAH0cCYjDl6huo7ao+SRLnjwcubVQsoufv7cen6Fmiqd
oW4QiyGJUQCq3AaxMUuc3y/0T2DyXxM/ILncajNDCOBcfH0IJddjQmJUc6Xvszsa
t5z7KL53oAuZfKoaYeyX1H0r1lOh/vs4CBi4S5JlEU1vOPCwkPoUQp8xZ3tGRNjR
p5pT5VC8+tzdriGRwV+rcZ/S5d5QOhEYIRBNmS6H8JSBKDbzN+EY1w/hTbLUR9oI
Cc+ZjU9YCKHvGXIsd/kyXoKWoxl9GWPm/C9w02NZR7L3ehlwjYLOjBs2oD+BqvZh
xw+cLGnWHTTjkiZsgzETrkzGesytaMQ9/ZN7pgdHojkheoAWtTocW8s6L6wHnXTk
MA6CLFNfa08nADrNUzIT2lNujAriWFe8Xp8EHLkHO3R+xbwUIQIAXsL07PBsdayM
Q0IJpoDtqjBIhUz/iWzfIeLLRgQxnqBQOH8RtYi/RzEAQhvKlboDIF1Ec2yaXR6W
NQegFkOQMGoZb7wte5pq/dg5ij8DwxLSVNEt94W3QAhG9gD+s4TTS83w7pTNlTYW
RLf9p0zWF2dctWkDFG+OyJ7IlGjGsZyCrWko6DkAnk5/4yCAKW3OE/hLDg5NOF2f
MIOQM3UzFrqIw0CQLr3ciTB6casMEqz6xV9J7+y3oja297JBNsby4P9AOduh6JpL
PNKbD90RDEXaeHlG65G4q2o/BqWZzbhberSdYR+tS1XzrSF0nOCUQ3mNJKfUgtSX
Mv1hA0II/4wTPlLqCMHK0QQuVfKpnsLymQXlvIjdgnW8gn13N1I4hpYKGpvmWTB4
nqI6BvGN/R+MrZ1mQb5vY3vfMAnBnInsnJqsVRCmXUNpTauskaAjANSdo6HtiEoJ
DbMbbwUP3uCumL1BzfGLGC+RM7F94H3dpeWQUSJybjTos2HDBOyVV2HsMOCmpqa3
3HN38LRXIfkWWP1lCvVrimu4cvLI3r2jkpmDlm7SecwSxY2nfapm4mun+0an5Lw4
cV+G872kCozCnPnSoTYS4czz9z7q1tDTLzp05CXq5oVkVr++A1DwJwnlpVpiQ7VY
h6L5Cs8P0oU1mAZeT9TJAXJl5VnBCdjwpU00SXCGVnliWrbIFGVC0SA5vYJpZQ1T
lREw2JtUBApSdviOShF2vLLNrBQqIWpJ6gDhINXEt3e60/gP7dup3KjKgxJUy8NP
g70B32EcfzxCiWyB0OTjenNqLXElaJjztR0roCkTQA+J0NDdO1A3DrleEaDj+B6c
4KlFUck7P5LEkGtT07JATw/lmjnmAT+Npf0oJureMJv8Qlns86tB5AJusy0cNM62
7+091e2MhEX5CXJEAj5hGDvR9OwvsU1n7yeXnKqk/Iv8Df4iJ3rp/RQi3pd74RqZ
W/hsszy/xFPiaN/lVhQT+pdxviDc+9C+ixyGZtrbgzpVCAuoVzJRdqo00JENBKrZ
O8AymBjIYs9uGt+9PijCX+7zoG6zSsRbNHQcgUmk9uRGHqAMPqEerF5pG3B+qdju
LDamGpfkWs7eD0FcF+B1tL18jV9pMZXNYkNYRcWl0e3IHnZxFob82hLJaa1WdBc0
NOga7OjRxI+qsqgIo0M9q8Q0/OTIShzB5Vj/DYUOmYkJKk47/ASyOzdoPCoTKWAG
talkpxqLn2try4nhgDmGmDccdxiEdsMpVO1COGJm5cJ08QlC7tPefjw7HgfsnDYc
2ec1uyAaEgvRyg/Y4kdpbN9y195v6CBnoRgdU+78lrRKnKbiskSBeVdIC6gpKPC6
+26jU/fDPHZadepPtFlVzlVlDIQYeVur4ZA6KnrKsgFJptEzWTtbaopgCuS/i7kL
spQvzW7TZrugGN+EPDEXQxgMcToykWP4RZBX1dxIXK91tIFOB9KTSqlPSYVLEzqG
j0JZtWsB6Mpq3HxrVFmlDTh6I8OrDB7k2YxFVZmukckhO4PPrHD3Z+pPifupYQTC
+kmbgShEV0vBuIGLsmD0R/pUnvgpPPzwaVxGq1zS5cHsDRTiH97dQxgcTXCu3NvE
tNGHY2vIbxeRBaFr89iKf119Ww6zrVP0rjsB1apccFPYE82LuDJ3Qqz6QN4zHsJL
37aYDvWk5Xq1J/6pTdshRDFbHJMLDShCE8pfK31UM1BUvL3dYrVYpskoFVt3rqsg
XES2dwiBdy9HAfKvwPDDsCfdE1r86IsBzGO+Ujwx/ld3+rT3YYZl2MMGH9kI5bs0
e3pUQS1YkiRGQXABa6aoIPxnnocV6msSHik2bjDohTHBx3EapQpx9fc0fBSy0Hy8
UP2Z5be9G2LCcZIlEBjHbqXQ3AabIC/Lf0ddb26fJDalq6kp/CCKzUEPZpqkjIyO
EKFdpSX3MEJGV2B55EdEeYIetE/AlXWEInFuXR3duNwL0+xrHIxdY2SmiBjtjW3Y
xWTO0K9g65Cu/4L7V+jBHgIKSUgikzXwt9ma5Vt2yaGnOsBE85PxJTJpce+SrrYN
Pkhblw3GYgmSlI0fIZh/Sy0S1gcRf4e89r6J48+ZYHu1/vy7Y6Dku7jE8VQqlbSl
NtZVWPVvQ4baHxchHoG4FCJ8o3WArw/lVW9CVo5SXLlyozdnk9s2k1mS9m5MfZ07
kSDBinGnO8HjIHtwo82iEgUw3wKIb5q5UHWprcaRqo5vsQwp0SLzLlG8tD8kk4HL
0jSivahUNX5TpO8gOeOrhIBjzeGW01XPyi/u5PRF2g8prdhGhvEshbaUcEMFEL8b
/dw39Ihr+wVaq51YWNYCbk9LH32z7/4GMjB4aNxycX4FpfpIVYyItivEiwGRoOmG
NoF+0aMEVpXq8wsoyycS/+le/DWz9V1SYaNjoyJaf5U+LS8HvuVtf+qipMII5nwa
Fvjsz75lEwgH/6s5zSatBtqehENipCCrAcYs25nD3+XVk3fyPIGixmtqCfF5EJhb
kY2JMEyRynwJ7nWaMoZBH5fZBupDgWPyzitIDGR/mA8EPFhveYhn19+eLSXE0M8j
z0XEvQ2QSTROk6WbwqgVtn/Bou1XFexz92uNwMuAC2Jn4QIhRElpA4EEXxENEl0K
euGLfWOkdxiaHO904pUWqXJ5TTuc6y6Yp/lkn6L4jM+4OKKUXBjrKqJ0HEObP47x
KNT6zw58EukdssfWOaG8NS3zuzfqtjj6m1tnP0tCHCbz/D2ftSQVVPj2DVskckTF
tQ7h3IXCn3A8Mm1Ew5l4UO48RcvZilpIIPmkpwUfUwH5+FU32mDFKInEkGfDaftM
MDfj+ZUISbF4JP54uf2jUbIdlPnvkLkpe/TELRJWu2+rDl2OIL7iNUTJ52MFjZqm
9vB62gQNQPTnhEd8IJHJaABuiqA0RbPv/4IvVZOxTxtQGUwiaEcgogOklwKIz9lL
pHap/kowtaDMrbmxcnr2/XLT/bdNpDlbPlUgnvDCTl98cJbqb3tZcg7sIfufuh32
FgjTZ1FM+GbiY/p/SP1yYHtK0ki9dXFv9j93NVTYxATViTRjjlbKIRTwamergkm8
yL+tUWcmKBBXbUZpDPx8sTWhsl6qn+kiFITJ7SmiNW1ECbvWUBG9Y+UHtFG/i8N9
ZH4hsbtz64TYFmwSefjLJ/+lB4P+55r6OAY1WH9Nctz6y8FSpKMw+WTwm3yI68Sb
rYpuioUAEmkAL9IWoTHV8sMG+zpzqF+us9yZWk6hw7JfluUx7+zPMhRRuCWfY6/A
/QGlipnkY6Su4ooqiR8jmc+cHXGbogtoOTwSHkWujQeXxgJ22X5HwfNVZKRcGJO0
kdWyhTxEh5gViSrlGyuynk0MbT697aKOfCUYAYmwvqdcp/bHaSdglEkEW7ejY1qn
Jq+JPLB3aDk8IUeo8ewyIBLBMKdRud+XfuyZjjQfvIemYHjghplegwfI0Y4on/k0
THZYNulXCUpJTplXOsqg2wGY3I5KaOmuZDmKxhvf1ssWMNICibt1f4qBFnuj7VDb
oIBFvztQXglDhj4v3O/cWLq9xiuIdry6UnvTDXMxsuedslJIjU90idl9ISGN+u4Q
o8E0iSKkZ2fDRJRJ9u9pWJv7AhpaZz3comabQw8tuamEr2dySNmLSNvMImjvznDL
/nnqL8zJj4AaUSccDd2u0y2XpQDYR2JFQoi65gP/4ylbtvwShWh9eMowW0fmMXB+
lDnbPiUEgRcvbsaz+twXTeh7KMxILYcKyEakWl8U4/1zLA99uwlGQCIUvM8aDePO
tduom42ZEHPuGGoC5XnxZzlWf0Tg/bYsVLlhlehpjyvwGu68vksD3ZBaGXtA4CYG
rnh2Kj2+0wLpmLE7zC5DIl/t4coAF8CYFtLBCFlbOG83UJ9gg9qiE9PclWKnHMfp
4DC3nqRdlz/WE22/mGL2TQrJNmywXtdw87IgkrTh7vnVVAdXCKnjPeAdFpw8ubYy
K+WK3LVbDJcvDjXJpXej/1PF2tlDwrjb/yAu1sa3Texmd4RBCxnv9sxrUVKvme9x
zFwu1+53Y0yZSNUtjpre/h0VvEXxg4Xn9jthNBNCXcUWU/QixmAhR4QZ5E1iHJmy
EczNuzQ/kKcppxRtJE6V3R3P6X1oHHaAT0Hn4J2ms9rAN/DJTHOi3puG7lJo92F5
VCo8B/5Okxj+opRN2/xPTJCd2fRxuoclH/aGnkYbXAx5mw+C8fQIuD3WBJiHtqNU
jqKW8gxruXGL2/PaduU/0VxJaOz7Gk3qnkUpFIywMk5blMgnC9STyOaUPeMA0s0l
rM+/E/kbmvFW1u0B37KRpofZIImmV5es/cAjp3KNKJui8BnxYz0dWUqiZpQe1G5Q
QvAwj5z4ySKvuI8SGSl9htiBDhQJ6gfIRZLUCNr/Onu/OPO/oKzFp+W1N2NCN3+q
xl2fxxS3uUAlpNIR5yjVje0xVgq6h0J5opg/hatuVkkt1WwGTiBIdw35E24Ft2Xg
7a+ioz4jrQBC22u8PI77+6nDwMhOFBM1OjAQ44iDIgBJJ2f0Ta9p1/A2WGXHtRbN
cXO688roaBFZ7m5wUC0B8GpJiR9SPWnd3cqTtyVuE2fY0pXYAwxYcjzQjHkhIIa3
hOrv+Rtdbs7gp8kF+6YXqWwZtd8lJjhhElFkzIpJXX5H6r5YByH47FWyOlA5rfOb
ftFjL52i9eYuWYVGMyS4Yu2VMTouftObt8LsNoztU4maRDwCR178844DwwdvHlKy
ad5aN3Gm/BmhPzEgN2wuQ9CdH3AWh8j87/AUK97lEBHi/2RCo4IfG/btsyrIh3Tl
8GnxY/TZNffQ3nOwmbqPBdQx2te/weSzsARouh2YGwgjZto/kj/1Fl632tQ/J4AC
xpeqfzf3zC1VjvySNWcOUCSSfvwajKQ/KpsBol1SZ4/TstUOsTPwKRq02StVboYb
oafafFHiO3UdeIC8/VyOFCBLAKhzXKr+Klc8c/Nxr2xEvhIXLAhALVHpUoeSy3ls
3ljVdA2bzn1dPArUo/W85pPOF84K1vV0u5sSiJ5BSLEN9lVGIJvvvt7i48Wk2or7
ga2JBRYeaNlo3DoEEh2czicr3xHhA+RaGtJcHuL4bCqOzFNdJOdGXrFf10Fnl7g7
MsNkFQ5jBwLPAdmXZFJu/Vl/OjIeLyCUxCBi9gayugh1v8RGpR4I4IoA3hJ1p0SK
Vsg5d4Djl6QGnWfcRz5udX9VqPZkyecwrcwt7v3nqdmdIg7CzPiTkbUH4OJNhDfG
FlvEGfCDJgLdAakKiOgMvYUqAYxbnMXaWq/DE+w7a3ZLNf+C99MdRwCsfC6DcSUb
cIfJQViephu+9wlZ32l1QRiyIDfHYbagsIfKwCy14AyLVNgfCB3gKcJmuIvOiHaK
60JF0kfRg8nSjZa4E6rarw1bCaMgn6m66Y+ccK2oBAH131NbN7f18hM8VVYSTuYi
LBkEcq01U8ySTEPl8Y8HsFw1c3NaVQTJAOS/U1eGBIUCTsSlBlv2IinJfIwl4PVT
OcmWXvfaCA4UGYuiyWHDq8bX3VQkrvj6BcPFfPXbC6zZ1SMIfNUTPeHwKQHyubU9
s6C4e/GmaASxrmgearuLv9xXI3KGKYvovqaz6UHMty0l9ma0dSAnNLJ9JQSn2s/s
D9n8cprE9kzinUqHvKzZH9vr8tk0rk+zk6jxpnVWPrLIbsqCLOuF3Jf+TZqBPN8M
+mNR4DeoMWUFN6teIMjAT/O7jkyG+DOqeyWzBDnUphhvzw0IGa7UMVRgn1Cn22cD
Fvh9VeQezzZ1xEEh2tKNeeCj7kZRrs3rwWj0ebLurO6Hlhu34izDIIXRi6sSkyMJ
nuEuN8J0cVhhRWKLg0mJ9eBBUaIugUjE8Hs7T1+MlUY+ET0RS1huTCPfFSGIPEYu
mQOcgY4lVkVUlxmLhmn77NpwkYYz9uaCNxNwutgrlZmM/P6EM3exC6Mkl/42IfLg
uO0fJlUiEfuox2TFdyy2z6cB6zG38GIBnf4Qug1P+CRgJOwsZq0JFuy0Zovf+bmk
fGZTO6JWFnlyzZtOvyJ/noRP+YkbYxbwKwxjlrE9M2CspUKmd0a6tkqYmMGNHrS8
Pcj5VWqJftqoWxOUQd5taj724GLeOzFMld24A/fAOU6Ng1q2/Vc8k+Hg3o998h8v
8bdPmWOAuTYVCAhZ/o6YW+CPjbdXkFAkuwARhi5HMafmdUDO/SuTs222UYI33tbs
HvwwTvcAjh8U3yVPeXlbpLtN1xXz9QMA9mGSoMaHBuKHUmB5dpfsN3muNwgRWXzT
3wU69bRvzfJWok0ATNBxFM99UtlU2lMilf7JLyI4hS9xJsJxe8JMCYtzVV4SsKyk
2mPfxMa3lww+Qw7pIFX/BiDcf3lI+ijKn2sxt9US6g7TtyW4CgXJNXoJitFuspeQ
1zJGFjlF+YMsM4yc2Y6eSntAzAoRl+nrVJLRJstbB9J4dBYCxCWR39DAMG07mNkJ
KN8FCc5Xr31FK6pdDJSPP/9eWpxuh07JRuDvtJd8JFl1G9cZCm3+jbYbR7C+ZTkY
NhQO4y+lNuFFppGyroeYIhVuC9fQYzyYAcbDj56VTk/Ul8TTjUjX0OB62I9PyODb
l0LygXKnTyrFAln2slUU+U36YF4dBD8E/1BtVbfVuXy0YsU8sBxbUEsm53rPHxbq
YzpU6Iar9+fLU5SqICIHTB2UBckuJGVVh8sgZM9KfJ+T1KPJ3SuVxn8sDKgT8Af4
37x1na8VLpxbPs/NTkgoZ1M7uYtaJ4vGLP+CdHuKZvGnquv3ceRiEqzuZaH1OGuM
bq83rYtKbU8/9vWfozV6rTy5ecGdHecofFqo+VXwuCAP9qIKl/exSZ/oDQ3sEAxI
CQhRpvNu8ejzQuvJu7fMbNXMHJKvRxJNSjW6oLLs33MiPVfuDu66XIWJ69iV03bp
SNLDhij76ZbB/Bw41TBGg6SzV6jo1Q1qbrvhLeEkByA8nez6OZR+QrsaH/3uwL4n
fZfD9lFhIyae5DdtBva7KGxUNo2Cwe2YAVn1OblwpnPm83PQYM6CUmOYf+le/MaH
1T8EjNONNN/fORuQJcZY8GTFq7vb407W9YWH/JhhP1TYJGOexHcysSeSXKECb0Cs
PfA3z3ijm02swXq5JoONMM0aln1TO8YG2C6mMwQhRRz50KLuLtrdzAZC6C9WrzBb
TJfEUx3h8Ox7yTYC7jHsIGueQpbxIHnXPab2DpNz0+7HMo52S1QABH3U2RMqB0Rj
vnV8x4WcuLg2900pNQOhIricCFelvzKwjegYgIf7j9Nunr7KeSRqdBeT6aD4hBn+
4ES49szgJRnjsgxxsuX34LgHRc0Gd0NaU24y1pZsg8EIy58U0p6szElumUmfqHGg
QvKwt/8mXfNx2oiz9HTjD2zAzeevdWLdePPEi5JEAQY1NGQ3m0XvO7QKVtQA7MCF
NPbVPJGELpQctDlKU2VWygfUvVgn8LVu5RRT1gV0v/K8YVHc1hgGCSxfSf6roKTD
Nzaho2qRJtQiyGzI7OYYgzG1pAgVVqvoqUVHVi9X6hnErRKiCoHrotR4j4WnxUbi
wJsNAhaPKiLBZAv9btVzUU2/4a3C0SzkykcwRqZ4dBvgUAPj6wrpO9w3j/u+0rl4
afUMAe29cTm2ZM+T/qY6gYmTeNIA4sesiXGRBl7sKZjjssfMVU1EsNjKm3f0J4Zx
luMXhMXx/FjklcHUGwIYMtqHWfDFzAUzdzEdsBJtM7xDGG7EGDOnlHoMibBDtkOq
M3SCabtN+A59tGf4s+LR3RHQPrxkEv31te8YlFsAQfToG64WLDXWvHJi0ZqD/R8M
CCpQqgdsvjMQbLWJ5CBEf1h9YyE7E5QIDIBVe2GHfbPHJbvnwTItS5avsbvYdwve
B/pRl8/LD2ubBHRTuZ21u04iK1mvz/Cuaqj6QALGGAaRMD9x4eTg2gA3eQybVrLU
LgmfQrF3oGJ3UglnKySfSYAzEpeYavZOSt7GVDGhFjY07mjkoTVXBc87+BGbEuZq
OhTGtOweW2h+xl74+rj/NrC/uU0K1hthPTEBkFUfvthBq55egsL1mUll8LuxWB7A
hWqDYTcgWnNUR3neB4TL+CnSKi7XO7mLM+ZpHhzfal+Z+SxgPMvEYYgH6DHmjb1v
FCkRg0Dtl+uVOdZ2eRbNu4zAIKjMqeLHzzlhQ0kClEWPk9OcVcyvG5hdQlgSI5N+
hKcuyrbz+q9JT7beJZQxNtot1gQqF7Utvls73ZrqJzt5KW+KKsEoe3zMwD4/Yk7M
k9VrPseSwlckxaS7soyKLlz8SrH5v9emvpvqzpJOv8qNOes9VDjp72UL0e0zkCEu
Nl3vI4G86AzVZwlpoFNHYOU2o1Gfsr/DYakoNisW2l3cilNpEV4mX3D8JwtXtc4p
wk+QkJXOqBiPECyIeWHRI+S50w97hKXCWTVVPi4+r2yuP9QoKAdCJ45jGj7VEY9D
2wsYXfTpjy97w7f9inc0f5lB+DrzxN2p4o1Qv+zh+UMa4Mp/pUQWzylmiXc5yPkG
/Gr7U/SrmFhcFsVpnqHLUnXbPWVmUNzJ2vdCurGtbsOr4jNZ/xlLM2ff8cY4Bwq8
8oQtdpaiWH1HvaakjrGO/6lKlw06hZwNiYLz9mdR9q5+YFytVpI4H2uFLjBFDQUA
2WOB4cQsay7RmDNzIso7Ti/24FKtNHZTLpe/XxT6qUmDC/W+Q6J4N1r6cA5jWDoI
SyWEkb8CAY/8Xl75GHWbSYZtxyEHk9HqSBxIX2zl6tUYdmgLXOx2xXithL6/EmO1
ONMV2kM+594IAYc7fBOmYXBkk/59tZPJIO0imiYpGMUbzJtFc8/vHjP4J7P0CBac
ypZKUR2PnIsTQMfzbPzl0iykLCMJituwbd5bVRq9QMFVryAZvKnOLt8YKoFJ73px
PaESiklBn+zr8bor1VzyIrE8CuZ+bqAFTF0OK2VkCHyWJNQPW33lkxYC106plMUD
/5Y3v71qAeYwcQr0AJ5u+LpqAXswnUPV1sSx3crXALm3LYAFEduhxBShm+LbksHI
4A3qTiLo3heSyQ7ofdLNlpTgmRkf8WUqkBm3YQvd+bd4ypucZDELcTPVb1UIVfcs
oLTLKikKHKG/fAtbclQRgemCv34t6i6Z2Jsm1JgFWPvKIXOH/B5KsvqA3+ski+sW
FznKXwtNvFiBghyMm7hZPlCEXQggunJVOCMV8G7kJzFlB7FShhIA1BFSecnLzjpC
uEIJLq7cN4DePuJxhuKYDm35Du3o65DYIf085CP/FMdplk7qjVgELBAe/cNFg2eP
b4nyYn5FkU78I6w0LaT9aVK8LDdZOZl9MuDB8Z67ZOfTfOnYIsD1WicJit8qt4II
cJMpF6gBrgNdfE+8tlvlOVkxfLgdBi7gxHtZnB4ogc+9oiP3lcKpqreA/O+Fc+Ub
0OXHWoLlhxb62ZZ5Ptn3yXuXpHF8VIy4e/CYsGdDNr3I7+xBdNHecF0i1SmpJRHn
QMKNoD0oFX979WrZn8CHbswClFPyFW1yesGPgGPjoHcIKR2hwK7zYaDLcYG1K+vP
FPLpljTfqebkpO65nTRFDP02NM2JI6AOX5j6KJ6zewGuCoZt4m/mIOBPpkxywD8Q
x4T5XXKVDyNxoXmg/MmVwWTKtP3IrmlA4hCh4c0kYzJ9EZEJSR9AWXZtirSQor/p
XPGwxDlwf+z5omiSGm2XGjc7RjPCkgqTi1WHI8B5B/wy6zpSYvkzavFmlUaZB8Wh
/wZABpeb4fzPmP/9p52hpaEOEc6SD7sXA9HgpW2HfvTJr35iuPf5uLWageqGJtGQ
SDbHNDVb43/eZcomhMqRtKkIczF+gTuA5hz+S4njOt5y1BavYF0YwJDAg9R5Cu+O
wmGIuVM/teFdR6+ehe6Ah1pGMSjdGpex10CXoiowwEYJUJN0/qto+tvW6yJc1rPw
m5eTp2mxYPHG+R5m53OPTmwt19Oz5CSxxtOV4d8W4b2wwUPITiyktxn/5l+r6g+6
JPH/hkaC4sh9epTT33W3AwgiV/ovWKk+qfP9TiU9qZhhezwVdjLbRllpksvFcE7o
LTvAOq1uCZJq25HGcipwzMraZ4gsJrRcKsqvbovTgEpEsMzhZQY/GzM+8MtMjNGC
IEkyf8XQbvE1zh6IF72BbnuMYmCqntz7fCO82vOk9S2KjL/dmgur3MLk80RqQBZt
ZtoOfnJvEurS2MtsPRfujNHyvNP71IOMuF47t+y4Sah8WYim2lyckb/gB3NvKL7X
vnXmGS+4gduHwQaV35cjriNLfJttsIBlqT+03+q1jag4ckjRBrAbRXWvhqt5z/VK
QhaLWOSLGM8hQuU/sCiw2gxDf0X/n92x/i5ytANwiGqQPigWd7EyNX/X6yZBc36u
rksk+4Ij+Bv949hlewwkTf7RKCNQ9dOezou5ACcxMVUEy2yEZPOw7nVzX/JR0cL9
yBUClpXhDH1Jm0FlfTMnK1m7+K79ik+hlzmxokIHxwgfuei7N5j/Zw7Zz8ShJNEp
ePYuJH+MfrxxJmJwuAC9m/msZ5cK5LsraChDiBDn8U1TnZKLG43fGXhSDue9FVPF
HWUpu9DsXtbmR82dnDwc0MQcbK85ASOmbLnpW0KDzBBVeLxCGulkJXwJE/U80ty5
zCHghCTHT/WaRCZSbVZ3uOYjObdZl3ouZcUPiYZ9CuqQVqNzDKTtocUVej7bIjPj
zJJ6/nd4e30m4TwfYTexiFu675MgstI4IO8hDcffyc1VVTRgSWW58RqyqbzYE02F
7sOcNBYgMylWxrK6Wnc398kEGs+jhKMFkCvd5kcd+8kqXIe12wxNnrBm/VcpCTKE
67EVFANiEn4DCVfLnGA1foHP1FyfQuSi2Hk+JBq9z2NHgoqb/aVs1pHKpV9mje2H
G1XJx9x8sBM0RIpv9Bw4T6lpXwsjRKjRYeJn2hHXaB+jYdnzb2zs0l+qDK2NQVWn
DpNmg238xCRZ4JKYqJNhEEoiYzwYC8DXG8xGUh/IxBC8A15uezQkh/xiXj2P8Yp6
8dbAKn5eaKtJu8FA2WVHE7Yw3SPM/4hRen2HgSXRebxIpb1Q8qA1U5Wh/4uZBR/y
teEdG4hwEGMzx2pWKxpHXWbjUCmHZ3Sro+XWMSXlmzG4jAQ6BsgesgzB/9jhbtXx
k666ocF2aFRHTsgqd2Si3rpWpa7KKS63BE3T0lQNRjmjAoD0zBJA4UUsojTj/Moh
4XVK3TVhbw8hdFvWeuFKRnrT24NAGzw7hbDf1WUmOIYM8Qf44MVRoxKP3qtdyBim
h7ibWbazvXiiNSn/PfiG1tcEyuF6MbQJNAuQuPPb7O1YJ+R/sCv8056LqFXSj8YL
cW5MvcqhWUYr0CVForgwAnqq2B96egMTwvZRSD+LyD2d1mOSCDlCsVHYZzkvR8+u
czJ7X6kKbMlfns03TOQdX4QKZOJcfzUKMnn2IAbEbm9OIiKI/Ng/d60Aulq/eBx6
iBA2ZtaXwgV8a4feV01PH949/MzBqW/iBXjTeGnrMbGR2yicPNmLJ0AdeyL02LjL
Fv3q6nhWwZnMpoVwYHBAtgXH0k0MZEaEM19t7AHvoNARfQaDipldJnYoPQbMM9kg
YMkYXjRvZHSB67in0WGFSnj7DDScMbR6ZIj2c732GFVl4yG9hIFS96bJ3TV9gsiG
6XogmWQhqhHwimNwyz3ShySQhMrlBun71VoD6t8AGVvBqaoKxhorkCoqVNJGJ7FD
3vRS6zJ9X9+ciivNp8zH85IeqsL+J1Ls5rrN9tv83P8ve6teqX7tlHi11xiQQyuc
a9uOdsFTBZJMIwE6CxcHD8TorSRSjGiBr4o+b+fRz8ECEdjRXZ9sESoFVCDht9gh
pLddLW13okwq//y3Ws2av3GW3bA2/J3OUnnVrgtWbNiN5iRuLJkK77bAKU7PZY1Q
PlppUUFIGCiy+ARcD5mhAkgxl07307CTZ0Be8imPYCu2jzCqh8Pdf29jLXxu+xEv
PPOlcN6HcGxlp33Pp7U1LU8EyzuqZa6Ic+NMVyMXv9BnpXyXGHRUqekbkQjW6Wgs
M2R0tI9BZDnucHF8btootD9JiUUCEWQYVpH68yn/sgp3QO/VMRhFoZ+7tVvDumbK
Xmj7HAePYdWS7b1tllDBKPqVymoxy7r6PZxp5LnKb2Y7H+uAA32rXhlS/YDqFkpy
VzxZvcCs6InvwdpOhoR0nk8RZnVQTIDeyNWzlRvRETdZuYhkrGYFgSlXiZy6ws4L
Gysb6mj8qwfiwsdo/DlgjgECQ3fgubufDP+ouMCkVgOMSOT7mXguO59X+DXt331n
JFGFeA2OlZMfq0ksjndWFADiB0LBLEuHFzN5PFSJtoJFAQsM6BXXH6ZKvmLI7HO6
RqHrELyYX3ExMoMGYWrxsg4Xxx9zMI3FV0QKgD4N0fPlwE87YhYJJfPV8vYTUHP4
4eZP9Oz2dDiLcHnK9q0lUpQP/lcTimnuG1ywoXAT4cEisK3wTkxZr47DrzD66ho3
Lz3JCEF6v/k/S5emaGyYTeGmI8OGAWHM2bsWS+XHAP3gd6/9Vk0USRLRgJ/4Sjsf
PFg3ntcBQVH9itizjNhmhii0r0UMXcOQUgLkOZ/fiGsDKkzy23b5pqSrHbZPjUmk
7Z85BkHYHPrOkD976nn47KFeJImJgFNUvP296D3E7/yhTwr3vipYQxP8b8wTUTd0
07s6XrHkQcdGyWmIU1hVsevgKMI+Kws6N25XZe0zakooiUGTZN/Q7HQPivtvGGbA
hKsdo2ljfvMHfxWUnLEDb2BpxDJWkAANcDhn4vNmZI2e/Povb9BYbwaTJ6hpNp4t
zRRxOHVkujXQoKwRBsR2M4IGxonpYmiSR+zDqPhZWwfo4Hd2vwyAkSH6n/FfwyQq
Mx0FlDb1Lb1D1VzKKSePdkab6JTKVAEiN+f4+i05CwVgRtVqx7quBtSeXiNLp0Rx
HtaGgRNXTShSxfXVzvdosfyCHm4OD//9r+ZZ/MX7Jjtvfl/FbnKhbKLbDWakR1J/
DXuzUIvyY0zTft8wHnLYOWUJDFLkde39dFBGw2myWeBSiVyjJF2Xp4sbi7DehNQZ
G7kyJES/1MtEQSjE7qfLqWngx2zLF8O3UjHsb4hvJ3yK94iAlx41dAc7vyUj+XKi
EKslU3OX0NZKk44gLgwphx53Fk8WCgFNa4Snu6GL3E1W+ZQ3YDeg98EU0wbH8cEf
A42p5bl0HKRGmO0fjDQTR/nF87ndjOntT0kqAdYmD9PL/ttc2hmEr/5EFwrYFUYL
fTbTGtzq8U3s7hxGwZkWTJbS478+8OSGjHFVgmRirQ/Y+coyIBFThN55eaYPH9Pn
vp5uaF2AO6sG6YnANTP7nNKgKeTTj0KpxsC0yH4GCm/kkuZX09QzCVlyghWspS5o
NnTKTx2R9VvQRRhoKrhZv+2NtoE0zuRiVdkIImjq9h4GgoigwEmeanAI4QtTLINd
NzvjAEUvLMtNBvlDZ97gxT4YdB65/dyE/ou4KQBgqttuSx0tZ+mCL8lnslBEfYOv
+4a3Rk/lqPagjbjfeAQA9LJufBGaQ18VgYXQeLmu/Mr9PKDqlIfrIFHWKKZBXdts
n9TO8cIVbs4+pnOxr+OtujyzQJFU7KbI8Ut2SKZEV3e/h4xIaCpBneRpsXPOeJNU
FMQLIPtGvYuchZceK7w7wvhfoiER8eG1WnVf/5cAc6UZI6rQt7sFrXTjHTWP8X20
/ijs48rrG/8ftkXh1v6izU7RbKp+K+/Ek60eIlYH0R3DjPaw/F7P9TG9Mzn343k+
1EbQng2LlRHMZ/qqIyAM+3FL2QRm56S2RYc+VYdVhkPojJsQezHXRh5TUCS4D+zG
lh9BlKkckyQjmdjbcasD0f4CnK3pPcD+mdZDWOFNAeeY/MnqyMuIqxnxLhO5CiHU
4v8JozUvYjmPy5gBSaHiPCZ27eWqHbj3yX9TqyvJm7kOTR2lnhZZPqWsrQz4rUwO
kUCT1fm/bDanbKAdaGez1zmTo4EKsbw0d9qtXOiMwnG2W5F+DQuNLDRDC++nkLc4
2jGx0H1TaYsnxjR4RYPdDyK3RzKdkAhaaUvoGPghpJSK54HV+lLvEFyeyg70yowE
iCNGrUHD8h3IvD4RTkOC9A0ukPkRIBlmowlERZhSGADpQXAyM731MLNeK6v+fPn6
Y+b3vdRGivMYmUb7mZtqLJiVVA5DMWj4amKcTk+d055XSJMRSZRO3ePlvV35yE/+
PUp/00hBJuKNF/vuxQHkRS2B+ntOoVaZNcLe6yglfMy3YQ5wo8P3hAx+lL5WCJi4
6vVK5VGrUE2kAWGcLH73tQcv9C2yVw7yltCBXbc9ZKdNxpKwwJwEKcNGP9d4WA53
ViULgzEALCHy4aMkEdhwdDd+iR8/ESAr6/qVfV+qqmaglM+XRTJkTYY84wGxJQaZ
3Uf6SorWjMkcTHAs/gFBMT8LUqBbvbVMTbFpmSqAsxbF1mfYRDDRMxPo4l+KVTIt
ilw3ONrEjdgTIXgxr0Cg0FMys9zVawktoRpUsklypm1S4tOJq4eLJFVA0ySGFv1S
iAyKr0AtjtrgxAt9mwkWRFoW0SSqQpeiI639dWMzK/K7PgJsMBhciop2RImQlFUT
kDmVwh9/WqSgZunTepbGsj0YKTGV9isoy5rZO2Ux0oiS+H6iVMg4QRyLMr2Xi0Q/
YNsQyL+nKw0x8PHShxMe4EjxWNqxXi6tLayloD7+ymvCg6j5v6QRJkx8hQmxvnyP
JVpdDE6WdDoGZvoGFoNP06rsbXBGgPPwEO0e4hkEEyNDxO9pbl0CeAKZD+RDtttk
lRzGdvFZPSikBvxXR24WmJh5K++pj7qn2MUEff8xklTxKvZoPZ+AS9ERVeBB07HY
T4gqa97SXonImFknajpiy9rjS4A0y+aGbnQyTIO1+XEGLoFjP5cZ4olXBHwiDbQT
yN/SoSwFEeJa8cIhJa+qECpehBtA614JaWLMyaZhGIoJ/bWVkCSY8jfmdKeEVbto
Pu5YziSuejh3wN+A7ku1Bj3rE9EJWp+tskAwT2bPpRv9O9aqYjmlSmKYRtmqKg9k
0cvajxqH7BG6LaBcMA2ozrtxQR2gTek15BmGvtxDRE4jmEVPHGQtPeVs/XzO7XnL
VFwDc2OpcdchmNfz/ZM3dGmYwreiRKxHWKwKvuMmI6pNigIy5Bl1o9evqqYgWou6
dBqJR/GVuYIHSjNNmWlDUY8eY6UYSWKyoYbEuKIwWDaSWhvU9Qzvkn8C7lPmPbth
mmVRgQfZ4u5I2Qmxkr1mweF2P4FElNBLWnQ/eaJbkc+mDC4I9d0WF2NQCpqrfDvL
hDluxnEzq+nzt3Zz/ES1OUM31DGdoXP1h/ko+zxGXU9fXlwXFGkJ1x7rhj+OqEU0
8mnaFS7exMgsCVgFjSaiMB0pPcTtHxcjTYeCBo6ZI3Ql8OeqNKjv8p804SrDItXM
8ZmPrx8rrn2o6TdflU4+oBU06LxHxBJ+CRLPPle+I4JnhWi4PRX0KIyBRgZVbf7O
CGlhK/3hxYNqBWY1+RuMjBB+sRWcNvy70b45zBOl8xNWCc0dVwxJTtzrQnRQkUhn
hSYJva7VIZUNpTmk6YuDXJR6RV56WQuJrqzFrZfjDA+WECcYXVsBAmkmgnFiz4AO
KidGcFLG7X6ia756qF9JI36HWUSs9/9gGOc0LC9usH3tiuKTyQqtp1+4lCteAttx
YrKBi7afBqUPsMQ5XTT4tUFv1guKF5dVhFVnmVGrYb2MwXpDXNCLO/Xkehm/0shw
xXnkEKs1n37+/FZRENcJkqah2eWyOrNdSHAZCrYe5SrIl0wH5BwtXckDLQHteUK0
X43jBkIMWWEv4XmTyV/Ut2KhwSiTEsnE8QILea2xuPYbOmDzeU5rCr6KGsbkxTen
qBjh5A1fk5UXQbOYNHjbZ+DuvswgP0BzGZR4ESxv6LXfrivWOFX3vzFd2vizpShq
aSZ028j9jsjM7vpAycSMhkAYF0ciN0SJBKcKilG7kekp7vGlxMRzZ7ykbgdCEvg4
hY7y+a2o5g8Ol/wSUuWkgLlTmVOu/ZxKPM4jN0+eZjeHcApQ/BB2+Joew0iWsnb2
95SzFMhwfBS2QECb01Tkvrd8MtpA0DMznZtrRQyQ0GgGDKOkXwRXCZpzsCuBowDV
YSf7nBdMzcgMo9tCctyu58eWa7mVVA6k9DgaZPxitZnty6Yt/eVPPnX/qiAGYQ/Y
BT8e+ni4+csuADVnbDDBEpSqV4W/KyxYcMdfZkkQGna1i25PLLYeITYXIgIN/6LH
XYUazdGMob1RiE/YNIpZhFAOFGf4jnHeqAG+b/oM0HBFF4kp4GmICKfS/X6sekSz
K4bkup5gM52l64ADzXMMqer6nhWR2OGWb6Xq/q5PrEiJty06qsl5vRnGdrq2l9jP
0tA8YOSiZkWonZoh34MGkkafhViArwf4sZ3+muXpzKsFlSgTeYZfeFUIa0wWQo6h
MXWO4W3N5wQ1DCTpU1UMpo6qYDbIf/UQMR8eXa27IQKezUWrXCnYMwAkFqm/WnL8
mDamCJY0y3UX8wXB2BUnaR5PPGC14OgiPdsAZVBnZ2WeIq6ldV6zrvh5pOjIVVve
BFj/fBl91IWeX+tFmfVkAlab3eCwKMEQevBLJuOQZfIFPkyRz9QAa9Yo35h8b/wm
idPmCapLFkJGi6IHjVfOnksu4SgzQQSEC9wJ3NBbn198aIvntWwaUY2GpDxEYZ7I
Tbm4Cbp0aqg4hghEgjXV2pdq5ZWDY3IkUBMFIcBjphQFJXNbQPH2lzkVMyIk/h5A
+iRbiFwBthGBq2bkxktF+Ufk2oafzPr6lQRzRAEkH24XdJdAgVGAsCWzmJrQxNSY
vA7HETt+YdKq+BHt0YC1MiIekhFpibukS7OIo9rmfOA3oHV2PH1Y4nDePlefpB83
Og8YrfH6BnqCBBQxB/hSAIIH/H8RPSy9yZq7tJKo9ExEtt+EWjkocqHvqi0bo/Dn
sVWoW5nEhIOJqcp8RrP7zc2JGY42X27i2kKcSr393L4OX+MqC0S7KX+8nM/dtv0N
miV6qI7Njcp0MZ4nIGVTVFk07fwJi6NLWIJJgi9Q3U94ANsAUFfO8hIO3ciLXjC+
rVUYRAGIdDRNOgFITCx75DOZb+ysLjyF4uGXaoW8sL3pJdf+KnOLIZanP6uhiQk4
PaO4ATJV88zgoP70HVJxpsxIiR0g3R8EA4MAbYtzPAxoqq0aRl7ICtMuPVPfWmPq
kNTObfbAhbKWJVDmu8M0sjroH2Wzdk7zadEZZx1gzD9G0ANO+wuMshHIR2CtdMWA
+LmjaD2XlssZ1nWM+RXLuNSTpj5k7dYWJnO4bnMxj/pcxyScoTvxllT0aH73QosI
x9ImvfJVk5v50LG1gQiMMPnokoi3wTwl9wwtpRK/RlLzcecZ9yN9ahDyjQ0ghocM
0z2NpPtLEU48a1yvcr2Rb27DNqUgSztqoiBncc0qXIScK8qtP50W+N0zLc8Fb8UC
IA1bIFUlkOWDH7qE/GPcDFVnNSCHX7uc4PbmCTWrGgqR4WoYh8RhPm0KgpkiVdKg
7C7r8+fvyurNQ2dK1VGnqw3WFRvuz+x4LSDrjwOsXnLD3l3YMlz5pRmz+R5U1veS
5G3uxUqH5IWX6yqdBGZ47P6vjxvmrLpN9c3nboJ6zRvlFG2TWSbdY+e9WA6AEjlJ
os3t4EbmKXR+JapR/J2NzhVUdD03Vnw/lKjiRYBZYyE7fV00nklRgZdPf5WL3SKg
rx4VbPAcWDHty1If5shQxwOi1/cEmwODGjpZokcLWixIkkcnS7N/7rOHlgbOZYaj
Atnu6sg2+9dZxPyo53vHu1ECGZPzADDFpopxt3uMdwpPW/YNFwbJrI10b9KoYbFR
nmRsHIqOtQcGkB27RnQKIobTyKYBe/1E3eHjUlmRU/vbE4/3khDTMhhK+dZLQu7p
LpT5bmV7nVfSuNmmDSb+wv0vewosFrUFgBP505sDsNbVIwpdazbzvqXXd86JiYBy
rzloTwbjuH5aFwUgeL+QLID63O078D3uQhWkyaf5Aa9qcjo70zRQLMUTBMUpJPFY
pl4e5uT6yNbelT2sVDCLRfTQa0eTseRyV+/iiUds3S3dHSiqbXCwm8myVNlCmPvN
XsaaA1GKtUqPmB5QNumh5KUJ7/fME2nlbmDRUrTNmxFeNzypWOXJiJEcrMv+OzYD
4WbFJ+iXGtYO/VPGFUgJ/Q4TofdaFT0C770G4jrP7tcoMtF+xHMBcw9fQ63QeBwL
vk7INOtvyb9x6HaYnVnDkih0l3GRPK7pZ85bhsR2XHU/DH6C0Cv+yhRBFtyNicgO
Hf7zCCLfvRu6boOhyavjrqDC0OX48JTb1cna6iV1q0N4ocn7YI2gfSVJBDc5lciN
v+M26IrRzK8TFaNAAM5Jf0OMnK1FlrmnoYa+tMjFQ0vkkiTY7TMXRPbQjY6Nk7RD
WrDYQj33snn6CZbwW+gmmZiGPtWPEdGwFUMbq6jL2IejPjTQ0bJk/9fUdZ8hJ0rx
G84E93XgJNHYwPAwzEiQdD+tKFc8OtooUZ2EOTa0HlH4/FVeFXc3LxnE4ZxKfX9l
vVGN0SfoXglSX0a403FEotIzOI15W4EvatcOvqtPZ1DHGy6CwPY9GPYB7odehIiy
CK/UVQXo6ZhdMVVC+WV70q7T/6LsWFgAuots+R8EomhWw5alRv7nxWFGZfpBWtuf
2G3oIXCYElqpTju5+QSexW+R7BDRvZveGPdnEtI0JpSk6xVik+rCmKuMnh4pXFNX
CCaGP7pDr/4UO3XWkW9Fn1etaRxQN4+ko9BOu7ewBZdgS8aH0JObEbF7A9nANdBy
Zdtl+oR397U3eu8p6SnD0M9hS2Nv3ixRJnJH+ys/Iq4tJYI1Vdpf+uAiOvtJ/Nuo
emEOvjVkyXM6WVbmvHjBEuhHsFFrhH4CQalbnndUwrhTxVFCGfFwi+tqdQHZFnLa
/dxN16Pgw9tL8prM8To6ZpbDK9q+uwu2lIo02Ft3k0x2FVlfu3wtR0wF2HI52j4d
pbA4RvFH4n9Hl5apGP9oj5FVVkwaTA++iaBdfw0tO9QkiA42iNt2X93PTlmccaop
ZG5IISe+zL6uggnXJ3dA6AbSNPu2/nzJxQ4jIVZd4ewHUovCfVlx3oQPV6cL1OWs
7XFcsoQHoRcL+TRMALRXTX51CEbCbo1yB4sa8r1W44DyK1253sqnLS6q0WZOEP5j
J7/QbFdA1ZB9cRPQPgoo63LxU5I3oz4fhM6RUGpN9IAHPaD73nbBfelZ7kPdnR9b
lorhdJiLt5PyEIyjL659kuF3IVtZwCQZvcE5e/wGuqO8z9BF7M2bMC/7pYbxSJlm
WmxG+6sgV497bNDn6cOOsR1gSks2OPiUa+Qe8S/lqPkxfTzjIqyHgkI7XoJzX0og
trBCBSsD/fKBIBY53TOqLkt0m07TO1Tf5e0MVb1cInpfvaQFK+ILNkq/0wz/2USW
6usPkZ2wC/uxgiYACwQCvb3jkcRzpWrywtUtLV2IcW7ZCujbmKdCRJCsn0D+FCVf
SS/8Nq5J0oIcVOtz8GVRZGSaiATe3ZB2SmnEek8/myLxz6OOXjWGMjFRHNAwsgvC
qKOZ1zrfjH5k1q3BcJtFJYCab5EAXgr1pa1eBrDxNC3L0+lwCPSNgKRu8WZhA/7F
HOc5BE6B69U2eddxuNk7xHaiPEqEUrd2ssIfFy7GLjM1U4xCg75zP+8gDQcHke6w
8GOlGnu6LEs9PEDFB5EYECcsXuqeOr+ZQtCJFOcb8k5PGJ/g7u3BcGwxgXUq/Uw5
VTXDqid6oc/VVakqWBDypUd9Nl10qup78hSqnOMHEh1A268aL2rs31PXDgiVYVCq
qsClDFv3XI/itJQCA80+Oqftw4bcXqCcwWHOIhKpy4PmBsiqeSfFYeSkJ3rYGsE2
QAMgOY7eY2XJ6s1Ug/mFGUBjkzzT1mJO645BBQ112ACOMWqTU+iOZkYBPirTvwTC
i6iWm/reuVp7UbR2cSORmErPdtC5kbt0dUEHUGJBqzv+mpsfY5k0aWeg07ssO8hz
2uIJ6ciDZj5k4xtagzCVnFB8Boz2sWvAsgzGZyVd26XFRAwQ4+dUhHeal11Dliyj
Qv0qeBAMmeshcp8bAwYb3ZjPUawpP5YK1sO2Qes0H95inSxfBu/m9p7t5EOutI0X
Puv855eLELbAiSd8v+euk/LTFT95d9x/xGwUZK0OKX6eyD1aXCI13lij1IBmd/cY
uY8OCO590p+VBIHsu/fuOB5R9D32HpleUXHs7k88aHgS77+OOZwieJlWvLQWbUJs
8ajusiHjTTok7gQaciMb3YbvJMKw5VkevLstiZimMSbXOxWJLCnVHrstNYBOsSD2
g9KIkLG1JhVD/fHvprpjJ4msn1sQQuGJ40F9Fra99h0ruXjrsgmdPGfYzsjI8J0x
ePBr11+ZJ+6HW1gR1DDpxuI1lpvkGPTNjECiuYGfaZ9z4UwwffBNyJTek4/43gSY
y0gZyCM0lg3T6nrp67lkBwl60xtxumS4kvYVNmnUDwHWuQrmIEB2kwyOeHQk84Ri
WygfS2wsSekFzCTJmoLuxSV57zsqyyCSEQl6pv0lKxwEiwZhEX4nwS7rqCHEOM4c
9SXS2IGCs8HEaCUJou7zsb8+wEOU1bVhDti8pp6CsjQ0jy7SU8aogLz9/U04lcPz
7VWcGLViBbvUHr2yRfWE9sE9OnMzs3z1MP4s/L5qKWpfzQdJ585DLiS95Sz2skam
seDDPWm48tYbqee8+Dl1v2eFXlPAgah/oK4pzWUi4yrL0a6IFwiGqAvGVN0nlCQN
EbYBL0aCa4pKy1zr04Ls2x5lRPOv82F0+IGlx/W81iIXF7NozQx3+BGHMXUA1buA
YD3hLur4c0xtasHFU/33IdZtqb4a91STOzTgZJsXQli/rpxqvDY9y+J6Tuhp4WZB
z0gGrWe+UMSCy3ClEuDJ4LWt/1XaW9FU8c8pibggtrX6dWuofeCy6hgV6R6EzsWq
vmVIcGvsx8ahXbHguqIWn30IRmfDjPYDdzDr1+6KqvEO0bHMXfYGyACHOFxKxsGf
Aw0kENgIztdZjwzFoJLwIM5HBUemHKnrr2A4jsiJvaNPLPhFMfniuQIZnhsHgJ/Z
P/GMWXnUth33A2SVNVZT9OMMYHJeehVqCExqtPY2Q+mqZinr3qZ05oIuRpm9kmk6
1qHH5Y6e5moNcdD4lXiaHfffh47X8ktLH9+/FkWXAyPQ4JykeEoyat1nEGWVUzo7
lXew2ljVfMjOYxuXBI2W4aKf2KhnT+DLm/xVl1qaJdU72LJicSGfFeG4DKDGIhr2
n6glyMZhAsBh3vzr5zBzefaMMz5sRrQFqbwryD/OYgzSFV0nZ4CpquYFFMtLgFWH
Qp8Aox7DwwnQ7fNqrEzNzKqT4e/+54VpgePXsMcMFaCBlABqb76xm1GPv+TqhWFX
wHTLEY1L9YpBUBmlvGhZmGg7WaH5Jd5BGMA6MhxJ6fWDJzF6vfvGQ3mDZlRgWlDZ
8Kp8mq/UFA//yVTNUw2P/aDPb1n0RTRCBLMXYR/NNr6KKJDfvrhs3T81kT4iDSkp
Rv7uF+sB2gFCvo7xzDGnVloohVzISLLozO/LwUE4SvHy7EhBHvj5CSJcii66GpQ1
s6+zpkSfV/4u0vOCuIVz1LOiM3JgUbyXetvWW9vLliK1N5aeNBvF2/f5Nj7EQlAO
Wx3d+EgR5EQdY9x5R5N9R51Mt0DFMzUl1sk6C/9gHhip4lzsl0kq8m3JkONVnPLd
s1SOp61bfF5W5e1o4jCMNiyOWfB90SedLL4o3zy7rWFCnPFIRYcOL31gBCtTwtEv
MFBr65NblIk1pNsHSl20W8YxWecNR+ArsLu6B3SVHYmPGKLoYdj84wkdP01gopfb
yVXKxKmNQ8GHokFLKcFH9eNs1f40awMy149E9bd/IUhJn1K7O9m9p1CjLVtLu58k
L6vlXvAXGMqOngvsCE7SbSF4qOAAC3shNTGsBC8IqpggnBmjqoZP4HqGeDzIENG+
v/Sg7Jrvv4diF946eUCkmODDLXaTKBWZ3Qt9Xek6o/HXr4pEhsSHZavK+XKv6lJ6
00hABGR704B1IMW7T9KU9gsDtiOvGUjhSGwWpEPVnf32dZ/vycdnr4scA/VjHmzu
lNpt+o+Qeb64iPWUIIlzrzuPjfCW6o3Ol44gcHBqKfWTKe6IThawN9zW50jtm9nU
lvE2Muj60EiJKxHoc3NZfIEDuJmkW/zP7C+sCg5U1NM8LOwLRKTqQuT+Pdyc+x3v
kLk23vbtwiOSVphKQUJIqDjugJIW4UY4jEbSPZctyLiKubMLWHGM7yUKtJH6I3P8
coPVeBoF6N5zQpxiP/mUmUicPobPyEz3pYNb6eRSh5dhtDGwGm2CbJqLB4/hXc05
nTUH/MZmJ0B9twQYiSBS0cao5NmkPBXSKb0FWT47byPotZFlpc0UoTyM/ui/lOWZ
7wzPmwPFK3XFElo+TnOwFK/Gz/O0vO16+TwZKy4ypn2A7Tdrwsgy3oPedJSOG82z
aBoEr9i65xHTyHIECchCE+pSbVDymCz8X3I8P8zyanO22FuUZ4As9Hc4fi3wMC30
kRF11zOI1BoBQioaTfFfAp2MKEtp+MV0vdDpglhD5T5dJTEVtlD20f/ZXEaJb/RY
1rlKgJelwPI5oheFERCYe+4mJuzLYReAXK0pjZNoX1vfJrODUGGWL+Le4eSVUefH
/Jfxo24LMOk/Hfa5jJlO+dbEdbPz5cCIXX3CKrAEP8OHGfRv5sE4k2bUUO5H9ucf
9vkRf4PqGachU+pXQzwzl5L5wGBRoL4aR2ef8GqFk6IF7up1eyf9pFzL1/PZJDFo
q/eAHc4JiIbtGZRl1Wd23zrSfqcj5+TpvWNxAqsIyqtXXzrRO1kaB4f1vKorbFQo
L8FhgjO4Qbe8t71A1bQF4aR+nGecTBees+M3S+8Wmyvy5ysoIi7VrEmNf1/+MyZk
KfO3+b/DR35i4NaWIQRxpBsTFH1GHnqjwYh2VU9E8fdgOMDpYT/LJWzucpfr0r8r
bAMY2RqYh6SuyyBe+c4AIfuVP1QZkNZdrgZZq91CpErnVOsaruCfMyUaexEa8aPp
/DjuRtZ8LzMS0xnUBVVGiQBbNUJuWW/Eml8y2gAUOO9Oh72uLaRAqFy7DcZzy1nz
6PYq0EzWFo03nzhjfLiQFWWe+Xd4bS0X3p1fBDAxkqfNVCZFUlqch8yOpDw1p1X2
fkUKnXyLY0LHvNswATI+EGQh+fRwTnWuquj2iu4h1BBvlJb/FxBhQobVV3Fniu/K
/ehUQqhobHN8zJgJKaPUJtsEo5jWv0W9XGmxknyOzL4y0B6AYQR5uyoaYfaVTCLc
aElu/6/wm2M394v/vtFG7SbAaCRgOHqL0Bk1yeqS1/Jzca0lpc0sQoxu2q3891Wn
/7j61+MMb5hWgdP0t2SqMnqaFTfppnzyyAiT1lzHidvR/VON18gaHMZkh+SQXT4I
jXrKkhlIwQYrHrZ/ds31MXXwjKG+C6R/bG+PmrkX3ztOb4juavluL+dMicse8mV2
MKPUq7dpXfA1N33xklGEeO5obompVRNkAOHe/3eQwq1A7LSjsS034SiEkienft4i
ieo3lQPUPzjrdaRDAT1BO5Ot3qt3KZsADLS24Gd4wW86BrEsnUOAEZlH3jK4O4lX
C40z0cDwFpRqHGDDZ7aorYEy8fu14pJx8ESpqs/Fu6K5RH/TfmI0MIAMzNGxJa9M
2EODjTJCWpILuxoZCwOkV1pkL7JfTsgApHf7QOAIDJxsMuq70+QLnwTinDgRkT4+
kycPsmQLQvcOgoQZeqpucNjjIjVJmvAiY9miD9qMdqWL/S/+ECEdagJdxsENAObz
8ha/6sMXaZm18r2r/EGa4nfMjn3yktLPgsdoVzT7J33Gk0ec6rGqMOqC5eLtldXy
fTZDjP8nHGqTPZsCxP+Y43sSQREnqDSZPYIHkbCwAYW1KUf3/W2axP4mv6goc0bG
fNphxrFprchjRKHVN2x5UnWuDJ1MnRzko/WRgPdE3GBCS2eJkgKnSEumwZ33jhjO
iql74auoh9GO/OG5J9pCKy7jn8PDMVHP5u/mUZfzmCaolwD+dPaf2Jqjjh8yWIIo
BlEADewQXm+D60sXVUSUKVhivvTLP5kQFM+H5trRnAMX1sJ4eBYHQM1tCbrFhfa+
f4EldH75hVLnhFCPBBPeIJh1qeP0nq/HXvOvzoX4Q9Sbr5UGb7VY7sk7Z5wEsXlT
3evEhuKlDA3NI6BcA5IUwA3HU4Sn1iQoyVHMXf87cJm5kGe9obW8bZWnWUYP6yYy
QtGX38Aoo4l8+vPM7JnmHVj7MT1z0MoJAosqNiwQo6N40H3zbVqQAgxbnn03sE3e
EC3d3emLHNg4JqBfsWFMxy99NCqGo9YkZT6mQ3rpE4F6OyNTi18Is5iMVRrc51Dg
EsPRKOSPFjqQoXHGXPKdx53pcu/VaRliOMS7clyIoQTvLn2Sm+wd2+Htwughw41i
EXr19+d/Yn2OQUstJhz1qw63vCF646kiSRgPK1+wJVITaLFDxukw0w2EYGTLieCT
Oo3fIECN27WfyDbGBIkeMqrEUQFYPLCYKSeCQP0r0fdGq/DcwpeQU6OkpokhZJcs
OmssykiYHYAhHtiHWj0BOJzUX2B5s7/9BM0yjk8THixwzblys4/+d+r+F8VcT86m
fXyYBZMQ3ltnecYr0J7fWaAaAYJ21i8z9yZCVFSUFvxfmSLL6q/cpaK7+2MBekUa
1RVmaEhPoQb5ztGiQZ3rHL7EDneAsDSbmQbJ9TXztJdwUFTkmj8FawsLaCNPngCu
QJ2MchM02j9U5ePGulQsC3eTYtVtn56mey29OcilXglYM3yL9LyOhrDkgVHJisEE
tlFfMFuoKhdFk6gplYhPhw8TOQi07GxwTEfkzJONLlvfxSnczGsh2r3s1sG/5Id8
+LwF80JApoFvZ+ZFgbDj1f4t0ACZZBsZa9DVIHdj1iOxS7cKdisUR7LX+4/aZpAU
vmBnMBg7aBI/mL2tv8s1cju1Mw9/nn02Svi0ZlmkVA5CFF4KDabVAVyjbhiuPBwk
M92zwBne1xOYMAR98O1Xta96rprpeUaNzvmjwehNUKRE1qUmbQmb2+VZRO7aJKV2
/i+o2bQqrv3JxfjIpYaTb3qhOKhEFYGVi+oQU8ABmBY1ticx/RSY+GegxrZm1BXW
gxDFv2kAKsZhRRlOSR1UX6w0YvGK8PsilXrdquBaMqLIVOWtMrplcXzkjX7u1ARf
9zJ6MjJmADQV0moVrK3fR5sx4IdWKxRy0EQONlq1VWvOv4cJ50OwwZoj0k/+kflv
1fMAU0Wn6nXnkwkK/KKjQSrNo6QSOnyHtSty2Ve8OMFNUw7eufBp4dDpXBiZey0G
E5FyTq7uOnrXPivhu48aduy51K6k76OR+SM6dPdiDW+zw1nCi9yVmECxh01Qukv3
zxGIHH/glx9KGlI6z2RrpVL84HY/qTtWd7XwikqVGRe01hH5GQDCub+jd5aNbQAB
Xvgl7kx8NFeaGDLajzwOkvpkLrT90D7VRoi4ToolxUsF0d0iFusVJkV6TwNhosUg
d0qdMz38xsZ9UhLiaIxOdYIpcxCCOW2ivbmozJnThsDy4Z6scOoxF0NtqOKGx0T6
BzZrAtM6tO6O7P4VhIaOTLWPsLu+F1RzykyLQyscqZffp9qDrfLc7Gr+koayXBEm
d2pbbXz+B2Knt4suxJ/ytGJD39TKVJUg78OjO5gykz0WvM7z+JIwS0phDhXnCLJJ
pDwRmQHDadAr6qvLuIFavWuDMcwtc7Lz7+xpPoyPlC7eGw1O4Nk2Yg4BOIHXGKw4
rYw86SPSUZeVvSA8JCWFuq9VUIz3fmIB9osWkV6vbQoVgEx3V/tL2evUUg16bn95
dE/MpZcZ/lK4vvAY2wNuaCJpvfpukTDmg7Vb4AZixQiyIa81iBaL+OwqnvYTagys
A/CORu6wBYUQMky18CEcwdBljPOElctqgbnadyHmga3vsUHKKBItq5tbJZ9e4vwV
kpvMC+fO8QZqElzfTeAeyXTCzFIOS9OCtuv0OQB4sX1EkeqHcMnykeAqzjo3qVV5
rG5elmzkm4wr3JV1Z6Shiz+D6MI+MPwsdaDp0hWpofoxd+2/NeUrLsUn48iyeI5e
9x0aAXriSZfhriIyBsn9l29a9vvoJqXbw1IeVoJo5kI7DLAExpnU1i7G/0WHRYNJ
VYIIcpGs/QdyALOf3fh4JNPnselGhdk55129jUyw79qzTEq9dLXr/77h5zttrM0l
pUy8tx58eBGbxg/RerN2jPKr6sYoyKSCO/pyczrqArECctGiEZyLVNvwVJck/07f
SJk1boa0asF7/sCIjEAtB0FgwzK7eDf9RCRMJ1738hucywIIeXNb7OMr2pBcAsmw
1YvXYUPt0FbRm+B+7MHRRH+4Mlbrnzqaybx/0m3TzE6ww4PgaleLLpSxhT0H72jB
dcHqqxiuNOU7RYvkw0UGRGy6PkHh10SZ4hfS7a82ev3DGEivSnITzMxcSoRM2nKO
M5WaW/DRAaeciv+TdghrfjlsYF6e25ODnAHv8nLF4FglguSXyeYSkOYNKGH84zAX
vRx5VLxctR7oy8N06NMe+EdyT7rNdTFcCO4RzzVrUbmkx8guUMI5921A36AxVCUb
wGv1cxAilr0l1Omi+7vaT5hAJKHkMirMW1PMVDStVobSrs5PXtTEQHPBW3Btx5/o
bXdz+zkapLnf264cJRtHwSZIJnYnG1bt+itTm+CL+xh//zl35g8wwtcEWXcpQXyy
PaW+6QD99o9XhqANEmkNdwz8wy4yhY3jW/aPuggZL/stEdCTc1/4gzBpo9Iz+77J
QEmKEX0/e8KMAnnnaeZE7nvtz2bad0DT0CVZ2p81OC61MLQQJLrW2q4hd3rudiyw
0WD+KkBZapXFa8nEByZSb7rOn5IxWWNf2OaYKCPIQQMkqjEH0WGYXMVEz/+Zn1rL
J/rht+fa3XmUSg6xl70iWF7KtCtCfEGJPOCQyKugTiOLyBct/+66gh2pWPs99R86
Xh0gbGidndFaYX7Mnr+Btv2bZTbXRvnuytLif7VfXX87J7p1Vnxty+KJHb3Yt9FY
9n4AEMCFVRVauTUpdEWpSfQ5I3ht3s/gl27T9ojQkF7GsW+9RfSdXxMe1wJQCNUz
e/3U8ysMQBbvyctrNz2b1dInmA1UXsY12ZjXXbb4GDhEjyEq04PmEvj9+Nm/zy2G
c/Wtmkq6Ywm8ZtBfe8pzEcCmftr1CxanMyv2OYLSrB2apuxHbW3E9StryESqyLrw
UGT5FhtqZdfAeHn+3zg+cBvHzwppN8RDzoR53VGFf9EoMIwmdmiMBBKIGxyUaJSv
WrxGm9D5Ii8tbvOXJMZWpRl2cauhEeNaDT18/4uXWYsF8vI8PhMObmda56O2EPkc
RhKN/zbLPV3nnB9vfMa/r1BvkNg9DBXPfqgOU0znzxa2oT80GfzRQWnTwLIqEVBu
6EmcGmyjgLSM+A7hvHygnZt7QeLIdaXnyby9ea84D1TS2mbha2YzfIBY2gc+hlEn
YlSAEVEcpYgpg/d03n/5/eGQ9jVc0sCMbabJkbh4Q4nVl5boYvSYFflw74kGJyh4
Yp3u2ATqYeS5/LKCVQqn8aDENc48/WvKgcb0SGzr2lwSxJF8vK/16r6UAHJp7JfZ
REQ9Et/YwfGztLyS6+wcx/4NSkbPTnQLUrmnjUq1P5CoorM+GrwsO2cft0dxxnXs
56B9CwuYnY1AsxEpkcnK8BBIGnPdCU5RX9NKzGHU97qRQLqGPmhlhkQUXBQYv93x
gmNIPvtLKhd2ljXIzDwD63yTAdGMDTizRd8BZJ8/vV1Sw2o015kzOslKdxuM+9fP
UwMrN+6bGTHCVTKR8rz9p+ZOiM2Jr4i+M0sXh3lJn1hHE5e3pqfP8xFA9ukIz1qe
OCe2l5FA2cOFn7EwJacWt99mhMO7ZRTRWVoX6B64fY9kQ+350NvJHGZL6vAyOz7q
bvlbPO5yCK9wLmvB7utCJco7J59NWZiLkIl6l5uQpPOavjfy4AnPhTjcgdlQAogr
+l8zoIPnVP0EU23uzxY1MrjIxDCdHOX+GqPnyuB4/AREhHwm7VjnCTdgne6YeTQS
oDzW2bs81wtf9NiiLV2a5ViD1PIQz6gXgJrlX/vTT3kxC3zZeU9AX7VZchV5CENl
8SmultjCCdWLwKovZYpM5BIlU1nPLrQ7dme2jQPDBJDY0vgyh5/T5xVZPcGRxF0z
d2EHwczOEHUdrGpOcJfEleI5IwOoFxuNRkwQ1NPH+NDWwIRwZF3W8pt/VbLT7RnW
vyDesXPO6rwrJyBZ3Um7rIZ2us48g/4huNWU9q76TBIu7lSuYFIvqU7G7aEmeTcX
pWRJBHrp4t9hqKkKc+xR13fkBj0gz60/ueAeayYHgEJ82GWg0Wnri3vUm/UHxXWK
/Kun/CrfLLwrodDgcIPduT8gF34n6ezaJ4FaL6hddjb2HxpVGLink8Ojc+5smYHs
Ak0Ke0jC64d3ToWo8lgnSIB2Ig6IJUORnDIgfwa3i67JNuPEdgj08gsGCDQViwOb
Tw8vu2vuNJ4o+WXdstBJX0W3mYqW5LKXNcd1jSHQ4PXqPuHjd/db92V0KbvT1IMY
LFBK1MJtKRKRiencXBnozWQeT+oijefZqoce9g95Rlort3mSwr33E9dSjEamDKp/
UN2QmbJ3Wt0z9I8MsOFRH9b9rlRfjjYJRjlCRN8aAuuqVoROkMXG6vs+DvVkPUbG
i4SAPBNDUX/d/kuspeyqEedeCQsTAIDk3VVcjUhj5el2hi87XnlWsoZyEu5UTlZo
+30BBzfH+C81FmMKgM1v4VYWJIPLSiYHp/yw9ov/bm/LVwO74A9+j1Z3JaLqqBk1
sckNcoDBwcMIgqaONL7MhO/v3e3ACWcfpoZVOqRkKqEguzxLyBxgUY0aBL2amJsE
vpFMFo8/M9wz0GZmkyjyH0n6sX9AgMyh6dg/uNVFBAURshuMYfELotam1mlfw9c1
1jG5wOLt/OkKJUx9w74Cn66iYsFaGX9L+v16YIVPTKs3Xj/Nnql4utx7cy73QycG
iFnvpzDq3IYtBIyDMNGUnNQXUUxos6MQfH0cWsyIR+g8l1aLZsGrfAc++nUbFVHe
k047INW6j+hi67YtseL6/dQ/i8wf5cfVWpcicr6cEh+h5JWyVMUNjov6YzrFguYL
QLoQf9DBYdCk6w3bZZF460FSpB87US4i1y4d0HCrr03Rf34ciJB6bijC8el94xtz
PjBrm0Z1dtqLuqck1lsbwRtDIQ8yumD58G3OacswyezGS2rjYVwmJ+CqZv+yoIwh
vJKJwR8TkXEIRC2cnVUUHUTRmPGJvBqH9sqLBb/LQqkiJqheodHt3bta5RA+tWRZ
O/fxlehPWQWx1M9qQVsE87YgGt5rdrxPwb3S/Yqt4WUAHZfsb3/mU2ms5cocSWyU
mNt/z6xPq/IsuxVpVgpyijWVRWgvZAtj/8OgrMKxllqQrW6De6caSMv7NUI74slX
3FA0uV5RzuP0HJrTy/MTzHRgEbyC+vz2nK+a94ZOdmyiCbwYZuwULCqR1u9ZASHN
xZrt7RVf5/0FCvTbgEa3wa0cR0xRZTQs7YCSNU+RhFkBsfJnI9Qg/RD7RKIus2/1
CcEuTnulqWrsW7MTHkoo+j8xUUuw8PK2mmwdBgUmL7LrG9K5aS+0XD3NDSPg111X
jqUS+zGQoQJEMtxEqz0/5tRJJNpe+qP/LduWYBD4OBLjReefvtNLu1pC+R/AdAk3
i6szhRQUnXRaNb1DmSt7BSD3Ye/T0d5UXvSYTNDq66kuQjGb+LB2Pb8m+hnSQ565
nPsFxZlnIwL2/Wfy9LvPLC3uc1XKHRn9chj7awJQ63go/yr37rv3RBIgQe1UGc9e
hPDSSIzg8c6A7OxhtKYaVXmDB4YloGPwqYKa0YefBAlKeD8RT43u/2sf/jBF8iNf
6ULcL2nm0Y4n0IvApgbFmLW/KbcZMlhiV5zCRrkyMRcUnMT0Lx36Olyq/xCh9AAe
udQPHRyCk/BupNDH+EZ4Rs9u9+6vc71SCo3yoe5AGS4X02FL4v9QTQIxQZJ7d33e
7PnGgWq66Wc/KwATqDqhuWImFN/b3WWJP5o6y+YLZghHJS+KBJG932ohpkouXGiU
qVCsKp3X5K4o2Te2jZ9VchRutgkOL1+aPy4NkqrMNmKuRjWrl7W/iuOvO6IG2ib8
XryDHSjVsT+1xLxmQcPrd92ZLV/s8+NebCT/KT2ABvZk+lKKgEGT+8ZEjKyaKPAd
NkRJYJcurMQ5aOANkQ2qg7KB70NVP4dnnivEHvl1MR0UChGFxLbDaQRTrM1H6zF/
+Txq55pBKeAd7YbonKHVI9BaxCWJQ7RGC/8DqevyOAawBTZ5Lu+V1pQOQhw+JJbH
Gx0HufHV8ix9+s9yBxNJ9kR98DKRK9QlegohSU9Ux1INPPer4pQ+nrGbGx5M5PbI
g7uuBMV+6OVUa+Q7MV7SQaNGKpV3NSYb3mmLA4IciV6i9WRxlK5QjjIF+Uy76PJD
rqf9nSlpqnRbktkN7YVW96fl6qR4ICxcYe5jCkBm5X5I00tuERwh35rabmfXOLuu
lGHjjVItuF8NHp2zc60KGAlUVDgUKVWz5OEbb/hAZKtmwqmzByN7JCMnewE48iqa
QAPN22zWHLg/I3b0oyghDVVZww2kpv4bAG1k0WF0vyWi06kqb1QgOKKIkIpiJF8H
UdK4m8Sn91Drecj61Blz9c1og0q+f8xPUgvCtiuF676WeL8npyOYgrYWq3aGIhV8
qwkuUq/PVNU6k5Ymxb9bfzhLljHLAk8xIHdbZvfdseoYNV2JLGl3f6E/GSMuyU0A
iANyH55c7RFN52zujP6CWJIM5qs6FxMabRmdIS75WBN2OXjvKop/4rAt4H0xasnn
NtvnDPFdxzsPXc5DZJoGcivOc9sMSFxRvt6tnfiA8A+pAZ/aRparvGFXQSFMXxEU
ijnYxGPa8HyOOVfuKmpSBkIBeAsmfh7vpmm+IzqU6qPH3gezZDWPFxK7bOEGa/c8
K42mPPkcDz++tKimhZvZ9g4Z98XuQ/KcarBh9ZZw+jOS2cgLgGaskHA+xDVwXWMm
hsGR6qLcg8uVk62ud1OgL8vxjtO5fdDdIcvtRVh4QfN8tSsQ2K3p5A0dhXpYuRA5
qTfyKTSaxv0kgmf3714aBrAsP64eZZi4XYyTwekuoRgLEUNQvV4ve30IGv6Iw+Cp
a67BK+egGcLcWD5bEzaKyuJlk497V2fgHPrunnnUHqIFCwlmRS6fNDK9yhKij3dy
jBaoCt2MI0LM/SUDazH77WBXE1HnZsf6lcTkPxhgpedj6JPSyiXQIPPksYiVYpme
g4FR1SefXZW+q1EKAMoa4d6rpcQQjUBbbK05JImbOj7VLUPXOTx7l/m1wVwOTe6M
3fhYsnITWgzfkW1W1TuQmIFywGHs+ixdZyd8pxID6kAhtkf+zaUeiYDfYOvbpgZe
hl/MkVLUPXJWuD+MFmYoyMbPcJGUDr6RF5hWpyS68B6JF3iBOCduRDtKT3WLBGjF
6+lzM2ewJVY3Nrn9Y7CEeqcbaUeLFqCYyLVYXTv6xrXSUWBhs9d+Bt/UETXsUc2Z
epgeRCY05lF0wJIRK4BbIwJvBTSpUBLz2iXvnKo3iGuH5cbnPbNWkTAC+K+17oYk
/J8KFhFiWOZeviZFrAbECjhgimD5fmZocXIeAOCW7MmJlqDoGqvYqJ4/YybKTi40
GLyeMPj1zxSvzHFyYBC+CwAEvrX1T5iXO9fXds1+g3N1qEWNv3V8nLWtI/bkCldH
YdvCVL1Gbb0UTdR6+fkS0N1E3wEytDc1wOGh9QA6dXK2NEI89gOqR9ZKEOutzHZX
NnXbtsngSeCoSIrOhvB6LQ/DcM4rBlZdSgE2xSuQyB8vHFx8wmlQK3W8vCCONdQe
rs49Cq5pmOBnwprqvU9p4kkBiPIMT7078O6NU/0QYMwfnshqxklx3QFuWLXQeQeW
T20dHCbl+uy9ii7J3LaN8eNsVyo7wJ6nzeshGX9uArQJqxC7bTsrxbOih+cb3MWi
BAI+KvqrZnXWd27o7XZbsQy/OuCU8tzxD1mIcngDXgIAjT6q/zLHDxtl2pc04iR8
Q03qZf+Thx0o3xKmkumMCTNop7t6IBIUgbJa5S83jd9XNVJGb1V/otumgIHCOmpj
mNmYrAQHQIPYtebyWRUMzmgOJnSG8aR4KCRVWP3HsmFmDwdSakgw25hfH6fLQ7XV
gQ7cRyL9IFUT5grz2lpqeMOGnbXTs7aiyhPWwbcfaGBZEHyzlSD/q6pjGQ3NaSs/
TTgNxUfQliNM+Ct22k+IvM1bd2UpTyiYhkIngh1L7p+N8ST5cA3g+vS4UBMwM/so
bWpiRkGe/Pfhc4BpDqeZkki5WCUjbaxnv+u9BwJAkI+hkVvTGr/0TXHhp2dGrgJn
ROaIVr9w+fK2O2ypFmjSTW/58W6L9etGrnRW94EMdiFXkhh+N+xRHWkf0OM8jP/M
mjOky0XQEGj03KeCpazJD78XiRBs40YDs08E/e+TNxgUI+SBwLG4ndHYfoEpR97n
+TcWsN+IUvHRchR/kQwJKDGzQJNXlpT6b9EijWc4lNNEsRf/oe5OplLIXtpJ/ITF
0hLi6enPb9IIGTxDmbm62uz19wWxUIkX8s1yP6MsuU7D2UDe/h4UCQDvaK4gjP6b
prBdem4YqEN9xUdSos2M1+/VcC/ds6t142YDvFdn/+sRhKEp5OLyteOz97X3tWNn
eS5N3y8EFsqX9S7QKfmvSDA4yhL9eqKIcDHobC6Tb11dpOGFIgzXqgfsFefbE78J
HO3Sm1qqFbFuqSKOZy7EFnp3TYo9oihBIWqQVNIlb365YRCt/OGWRPEib5pQHMRr
mUItEyPkHBs9WFqGOVDT9lAhpIv4lEwhhpQaGozoi7RypcOsrEJd1mRzzTcL5/j4
nXVgHqHqqN09UTo32iCrU7R7ssJikSJsXrd7irbb5bjDs4XSmBFVh8x8ThJyXkaL
A4ebcIqdS92bk1HCcrOp6Bevyb60yeNIGt1+6x2sD04cHlO6/7UkL43e0wQr/dKm
kcayReVWUoBCNPtsrRokHGZx8aSrSfpRFS/NssvL/zv0dwdQMnv9CQwq25zj2Q59
ZgR4In5cvx3g/asrrKiF9sWGgRjtqQINJk+iR093M/z/HvyZO27aTnL5VmF01eCy
qWwtk7hl6wqXIi/kwHExFM3pI5+haLTOgh+OICWCeTViP0/9sdTdH53A1Bqsvtj7
oJowAhBOPJz84b2Q/knHao4sKzZC3G/7dT4XzoCSGOr9HO9AuHT2nlQ6FfxnklRz
uqAbMvqVty7wJRU4VF9ZMH+XwYx2/l3lqBuylVIT9UBu4UcT8sj0Fp7vuPIRBJmQ
EwgqMxS3yV4wuTtAgWw+MnFJ4VhuZmLUGUVUjAkAHs3zzUMkkyQz8P5Ry84ynuQd
szSr430GX7wzUtpWaNlJmq6C11kJ0CsOJzkADYAZGTCHEF/roquWyBpYPvpVF7nM
FEUYnd+RD6ijGH0TQnkrEZ0QuswVaTkCSB97wQ5cR7y/RNr267ZyCILRLh8sLYaG
q8Y/pRm8ykQpt504EWmtOY7RZbb1CPBkFqLzGC+V8q+/dVmME/ZZvXVjSCe9Qlu6
W1AIPZWaY2KQlcNX2m8mteZySrrq1rIdWIf7HH9ET4lHVJgUFvrp8jKYdk9xOjZN
1wq82glq4sF9R6Ea603+ZYQtKqwGvjDNWV4xDxP4JJjnXReWTmjdO/Pd+tsdBi5V
ArH24CQCozOoFlH1n0KTuof9LglquJiLM2ZAWw/jWDOYZCERbx2eWKGBNC0GXAX/
5nl+hv8guROH/5pY2ySsJu+KzhozAvmjkzRSQKdbzK9vGCrJDYZvZDd2WltldjH7
oGZwvGk6vgpIMBLtIcWJbXhgqcPIkaAeRadTJjzvMfWA1AnR3l47pf9fxqmoN7A5
0rPWqlKGYFudcf6+mmTxpGS8bmAMgl7dKy/SfBAHPrYhzTLjpxWDjISziylXRZba
2PuQVJ8xfWg5vQMZnYYmDIXQ6qtCAfEj4oLrH3i63Td5dr4nDtVDPPPBppFhDOC1
o0n+5OCd46j8iWbSvCSm6z0PreVav3sJIfhsJsHcQRA8cgoxEe8sApNOFDtvL3zT
ffU0A+BoCzOWaGIPcYeGYGqqbPiwFnXJNeiqsQEBDRk+u7/pZ8GQUQ1aqA/NcFiL
w2Y6JLW6YqWuqLqVvRraBo/Btlsj5dA0GEZKBxBj2pQQCHH3SfiXL3fZcl9yAb2v
jLMGXfQMy5277f2HJ9l2lI9/cFcvx2A1/UmbEBRqY5pu9BzugA1zNeDw/hWx5Naq
m2jzRWacBkrJviTEVE2vR57e0Aydh2veruE4rtX5cuNKBqkTSpGwdb36rVj8JX2o
GSIuc2MY0flcoiEJIs4o7DH/P5DEKAVYWG+U6aPOeMQXDlGzxo4+dCDv3NeKviiQ
WFeuZVVsk2KOeFTOafDFV1JVS5F/UCwfk8oO1lt4QyKuceUSctEsECEXfq1E5Bro
6JbMXUmjMY1xp3Sxe/wuOE4SBSqbv3qG8tukoX9SsNCm1oj3eDewyGb5OGyY/QxW
Vsfqwm1XJi580bUVDbYwgUQculpAV2eYQ7r8IMKOIBPwu1Uy2aeAimEVp5/S8rY+
fWoVRnFzZlRXEpp+ajToQs7l/GSxwz7fvF+gQG+uCUfSyID5wpLB4zQZve/Xweny
ZPe+0ESDbzGQ7qq62i6A9i0bL0wIiQMijFXIRT9rsdd94fVNZXf+XQ9Z+yF6+xbD
UCN0COvDCmKVha0al6fKp/Q1/5CiZYgTIjsOzYRh5LeDMtGxDYm1fblWMV22TfKy
zGGfLie+2RI/DtCSysQZH6aFCn3XMfnriwJetIJSu0jgMTgbtysLlCQtCd66ib1C
dKU1Lc2SRCAWNI+MxHYMQqMS3tt8fJJD7+dLKDp+mTLUDdzfmhsU4/ptiO9dM/yS
llaVA1haLrDvgi8MhahmnGjExJVTwQnEea5Uj7LjYcuuXlyVRqs1tx/CetJ7h8V1
xMGLtzsPJtFS72zOVs+78ttdrHHxNhWudmMg6MMeV07H0/OpK9LGi2GFfoU5Zs+q
lTJRHLyim4Ynl9IzlENtR0wg1xUhULK8kiHEWLt/8i9vxYy3kgCuHQR2oNdvz91b
cu1VP1W1cid7VyOJalZoDqzNOy5D+szF25OtZnTOB6oUvx3iLYPuSKMW1p9fe3gi
H0d0EZLFThVVR4UY95YCkPM6BUqANR+fWaZ+vgymCHdrP7lwHjPi0B5bTFNVSi6e
PMx4csZf/ES/MqTQPEvy2Nz5vBjc1/LHT2pUD6+ZFKo0Kso7GDqa+Vk0YKNHBgRo
pquKXr+3Q62dO3k/+6Pap43V4VUA5XcWekjl+eDOhiIB3gasqcribNfKvf14RoDx
ePNJkYVF9h3MF1/xCm+n+fA0MXRiKEcxBVw/KWn4XXALY0ApuPBcmXEJYTjDQuam
IwJZJDk2azBofAeIMDsVgUDF/FbyMOTMbVQNnZw10P/XjWDBnhgo7cDA1uUDyibZ
Xwn4HfNB4uqGBhjqtO5EOvTcK3MTcwgdzDozn3sqsT557Gngg/dygafiJ+IurwiO
H2tDvJjh+7lAUkVG5bNcKYBaomELFxgsMVjKqRMoTd4/8u40Il9/OynU33NbxPNA
joq3+fkNNN4sHkb4bK6wxtunDxlhQK+TqsAXo1Ut2OTEQax1tRVCk0x99V+i2kWo
DJjGJg/VWSQkaCDdqHQDHyz1/tJXP9a4ufuF19eLhPqUDvQe/qd5UNl2ouxzZ+Jx
n1hKCI8UU3Ish2lAeQFmtsuHA5ldv6u7DDkMt4hE1zTJaSflD129vHwcAQxMmM85
NcZeSsotXJuYGOZl86wU6s0Bev3sIKtsIpswdwlK6icM6aovexuKIaQ+VhZSOPh9
CxvUP0ASTLP4t1J1C+jNgvy4q4O9/tyRtIlfnPrzBxxY9sJRvjLsU6oJJlzLTm47
GRAdbSBpxdz4lyOXxDa0gDiJmzCGfhJe8+CrCuE0FbI/wHM0ok2lrsJQZFRqu7o6
PqgkCHNL63iI335DEHpVKb5hjSWafT/8mhaAszmOcWCEpWf7Bj26PTFInrSTJ6gR
l9DsLVdmiuVNh2EFNa2fZP89tUAkYQj6kN9vB/ZeTkjo2RHyfPRRPPRTgE+qZrpt
Kh1DO/LjeQ7cnzmshMuGRK4qu06kbOv9TIB3VeF9OtORTp1nBcDsSQ+geaVo7Duu
V5CGw2zCmfekZWbh9RSn35+ZSZkOQ8JI7dN4JqjcyLBnrpQ0+qoepIi5jYxIagO7
1UtOHQZz0WwTFHN/84okWW3BioWfpL12EqA+h6/HeW5ALbWpFzN0mvSOJbvjSJCy
A5hLBwKF0WDDy3gVHT6oWejv3B08GhlT4Ae3V9eyerh6spZSz8XCflrfzuTAd3GR
KjJuCHtirhEmyfXb/uqgxUDNODocI2+Fw5uxcIekym5hT6atscgqmcr/qeh7dGoM
k5VWvdcxEN49sLeHag5bPk/DAjJbrSBm3k+KwvbQNVQWAUmul9DTFu1M6ShwOArX
1rZqrUgVib4/NQ0NkKFvOTTuacpzZDZsZjA3C8uO1SOeRAuX0QZodE1Difm8wJzX
Oebm1wb4nsFI0CHTvvzMM9VCogXWHPEKNanB2d+JEoxryTkZiCMmT5iMpZHU0xKZ
4g1tnLY6dSMTYsyZ91Z56gO0aUiat3s7z9aNLYGw6k1q09sUw4kRSK8BIBPYV4ZM
9569wdmn0LB9y7of5jTRoxoBGL1OBS+4qFWFTmOFZmw115fUafkzJFKiaHBrNU/k
PhNL52uo6OPLdOMkhDM6GDRrgs6fc55Xq8GSW4fy45A0zmfT4vw/SsuVf7MPGwGt
MwDlmU84GlL4PfEpW8WcOI2zURvL3OXy8G9/cnv8thbZzU/TIqXzrkm8Z8fhz/Sz
u905Yzhp3wYG2VJyskQs8lEQwHlIcL+TMxgvID8wohvyvt0lCvFxar8qEZ9TAX83
fEvd3dwm3H6c52XKYU9Wkv5qgqRYgLqdEvj2PgZShLiuK6zyPlgqY7g2dLYNaxY3
jrKQ/fyVAxamlOz7N6IY6asDIe26uSaH4mKydiR78cmufhRsi6JI1T0KJakPnQgw
ureWXi8aRGdR/CoshEGd4jgQbxuzDGbDOGXXeTbqeEHfJVVwhqI8j8ny+auSYNnH
upNufyxgW09PqfpDpDRapX3fWTpP6HTJDQOBLuBG2Jr5hddhotKwPUALoKKm5jJk
ktIEx/C4Me9l4S7UTy5LltcFWjzI3jCI6ztldczBow42vhBPVHAenQuUczswLtCD
uBA0qWdc5BeK4af5Ss+toQFmCV0oVBqBsgTI/8y01Oq9LwaLu5IqNyqKImAQlszu
ssOMlh9ksUah+Oo2/n2FV6OiLmIzPT9OD0YforWZO1djJrk02Lc9naA08q99i1xA
IEOQprv5dXNpUPcYhY8eB/6Gf1lmBvC7pw16y/otPglwP8UVFR0w4GcCFjWte4xc
rlZe+D0R6XCZ85Ia1dtk4oeC7viZkjP2s/aV0uIFmCSkhuVE8JlgDmhZBXTQsaxF
E1mMLogjQjyc727+g6ShBZS8nvHPOPAI533bnVRRokppFjgMbjP9eSP9/P5GlAIq
4ApTAWRiCDqNF/IUJuoF2/cK09ov+bHNICahCDRMCgNAYWU2ksTfFrALnft7kUJY
kEkdA9QfIcBjRBlTa5v7MRp951aBUKhKR2sfEbOJr8ZewOTjz7zoA4HVpTa65GJ5
7cN3Hb8VEZ0WGWnhhcWJtwLeb0HB0ClWkB+TjM/7L1oxiyid2dWJMy3Fh/zMmuzT
GIPjBhc1L7zLre7pxH90yNUkvUY5twF3YeGYiE91IfaI6OEqSrLu5nQjjJKBfQfV
v6kYBh3E6NGPeyWItHW6vPrfkwVPc7dSceglSHoLwSmk9ul5kwAauQc6RqTnbqbh
6l8mmaqxfSf3e/A2DzUsqakKkewa8aWUehVGP7KDbeUPjJzmmpUnuhIr0sMNA2QU
A2vMafwLX2WTecVhGZ3U3B98bwA8bxI/OUYfOXD1ky4DcUYmPnWwcqK4dfACubPo
pXMazfQoGRRcUn6CspjohLPrYc8/4Osp8YPh7lBfOwHNvWlzneVGXH63Gi9YBNUH
ZVDqEs6L+g/97Jr7NPvWNrvmMw/0AFUT/77Q/sonB2TRjkMG67109VbwUu3VVduq
CV5aRua+hETDdNg0xEcI7MW62VnHHYgZ6JrtA6Jb1kC7H9QszSSStTNhXBPuBd81
NGI8/aBz1mT8hMNUoLyF1JX6HkDNTzCO9S3sAm3H64Vr5DYJklOrAdRRcs/Irikh
jZyDZipUzX51Kxodcc9BWdR5RDuQaKEand98JwoHm90aUkwoFyxBARa3mIea2nu6
jMJSGbUPU5elrb/H+87UWluiUEBR3L7OrzAwaSw6Hn7n/wlA4DbU1+tP7M2x7JZQ
LK2IL6X9fjNH4e+Y9MUfHCUj8oSmQhJ/Qz5A94GpnsyReUSBU/Lqk83gd7tACFSz
iVlirLv1YNWYX8g93vUYY6N3yMVePtdzvptOK9zLdVEUlkdzwyUS+kNAC6RrikIg
uXMsubx9kqrKUoaSytmqx7nIzt0agfWQXi0pVSLlzqNkvPQr6hWTBA66S5TGIz0Y
hh8+++7QMcR9k91nxceoyJwS6VDHEYf/pbKbzkw3nYM6HYnOW+AE4mlxE6Hdn0vb
E3aTdoDifiDMfq0HSclHMp0NNh1NcoTxra5ph+p3HsHHnkydOS7RWRqhW2Tovpwm
QWto2BWcINrsPTIUj7TlBp1aFg/WHQIXvQ5rEOe3pQ2r6rzw6gMPjK/PMllGhyEf
LRvm+lJWNQ5DTucwj3AkygMpmhUr/eUeXgvlnTPdSmCKpQeEKalceMbaAg6/iWPI
2fHJkyzjmWJUuc0IoxtEX6rP1RGYlJVXguP+BeQluO+J4JigrNTU+DvYSilhqKA7
2ReZZF8MpiW4VzJi3cFxROUSkcZlfmHCUtp1wsfb+MGbHt3zpcs266rr1+NieatA
5ZeWi8X65GUXBMmEPwXvOU8Q9pCqIBx1OXYftulidx7kIVk4qi7Hyq+AVuCwUgi2
1JtPUmj6893mxlozburdEqqpLxmCD6sOxCXY+xv5ddPCyGwwh6jHLyp9o5QpzvNj
H3dNU9/V0wH/qaJCCJ34C+LSHNC1UWUeR5DP6hvizFO2qk9B7IyEWJwBrat93StR
Ynp9WhdF/uRSqYQUul0QC65L/38Yony/8x3HTgGtG20iNpEeK10tVLlE0eCZc8wi
Cs3gM1HJOPC04059s6cULH6tUlLgzX3rBNBVw1Sd9WGmuMw8K8iiKXjy3lR9LEyV
Eyrfzl6l2oIcthbb5z42atsnqYNWdsKI9ICkouLsF8wZn28Ex9nxt/93wWzZ4ucc
e+gb4aEW47HujcDzS7OyGUmDefOD02mN9T0Ql43e6B1mZ7W4KOcm4Gl9IJcyyhYC
lBzhlZg8ZzTeEwEq4Q2B+cI2IUAm3mPUTgMX0lSPcRBqylVIYRutKfUxf0Vi5hV3
LefTdHqTcCuSq36J5xGFXQ6Ca273yLxcergI7GUiQeA1fn/zlIaWjlXjUzrQ6E+0
2TTU1l/lHnn1B9WBMdOti/gbkk61NEJPV4/PkCSBoRobzr48hcraf2H+DUfUbhnu
aZ5BLyRSaV0l0G0yzECfE5v2CHN5p99j4uUZkW2e+soes5m+zgtpdOUl66aDwGe7
PADImlNRVyKINx8E8YSUEeV5yfsBrZt/0oVhuySsQ125vANSmZuwL6MywqsIwcvm
R98uft8DhFtFNVY61HpQ8/4mqpOwhpK5Rlim//6y17udAk/Etxmuqjuv6oObTNKl
L5EqCU1A1WKgjs/Xx1y0zeiOs6W47rrR+6Hu6cb85/jQZ69Bt0SwjHCPqbBz0TPr
4hwqNUibdmiz4ZZ6JZLtYzBqo1yRt/BhzaxJVPPX6UhN0hGR4nR5zLJGbg5EKtmU
oCSfF5YFTkn6cWJEhmkAxBue3WvtcQAdJgx6k9q7XSAPG/kIE9lQWnVMAo9uoURo
o1Mca+JPAxTaUdewIHGSUFmWSFkSXTaGM3D1HmlO3FVJppYGX44Z9wgaJXuhShP4
Nrop5x8A1fCCEirHEMBBXj6o2RT19HjblrO+FYCfBx/KekNRclZqMwwsp8ztGaln
sXlLvUGL/h8Vyh7/hkYNuG4X6OgAvDBjVQOwT6skDScKywrOmu2/zrUadbgNn2Dj
ZsL3ZXoCNLN264HTw3HVWHDGFxKDWO+9vm9ky1rZMRmfiM8yG+UMHHhxN3Wb2rja
fOYptQynvQejO2OAoxIE5MjRJVvyJ4vLPf+HoMoT3LvV0aP1oIwkifWxaRrcIk3h
6oA+PmgF5QxJZ/cPvbk4qfI1hE/t8TsdEwko4i0jNaOlkxXNSM0yqdj2lr21+Xm9
NyyQlBg+rrSDePf4YAPdl3QMUJrhG1FdLZaXm/a0mKNibB7CQeRqTlQH95JIZij9
et1R+8PCQXtp/2dIGtH+TR7luq7xhV5/C+10ETAVd0XsgJHTTf3rtYpgnpzm0qPr
0qRih3tuAadZCtfogrSUYrsYNxRJ7aSy31JG6Q/KOpQf4/troo5JYDQqI4IvwQUE
nWA2O3mHwK3h26GsyNUXyReA7lqVk2+oLT+2mbxUr1FaSrgiO51oBsDGLgzxeZlV
cwjNWO1guZoBxduRjA8E8YsCS52nSOZkag65xXB00u/gMwjGq76Ax4PfHMxyOCrJ
OYcMttJsq4ksCb98Nva35JMQ2yHyE9IfZUZhAG6Ag/Y/v+kBQsJfgIBVZxGHsoKS
re/AujLzysvrKWrlsJSwRM3b79b3hngb8x++pMMkSnjmE6qjm3+kJMmpkfXGTZuU
pAvFjDLsrL/dEd91UGemxTf7JdNWcVY2IZSL7zFyHdQxGOh38stZEIsUp2hAyOS0
Rq1omGtT14MfnKyPxW2sJcswUjhIUR34sga6mhDuigVmgAgDr9sGuCMtJS7GjWVk
yBcX32HKi8YXTFCKIvJGOo2oUFcDF18ppUaN7l2fmEQgalSXP/BEPyepI4xLNdPn
IdOGjq3Ry2KTF5DlwLX65Rji/n3RnAZxTxoW1oY+ZV4nKoctqYKWyQc3pQ3EDMgG
IlLg26VMhq4gQuNSctR3/812cKsx3RdYckJbsVqsvizIOs8ra6cqhepcFJLz4PFS
QT118mW9JLM5k4bK9lUrs25p6tpekLlOuRl1ocGcm15iwCbthINjWx2V4a0thG56
6lzROIpqdzHEn7zLwOtdpwfmqvax9S5drusaDQQCOYOPUk+04kvY8yWbqRMb9ZLz
q2USYroW/dMXrM/cKix/5Di1kGnRliVhK4w72mj5g3Wmscswd4JdNg2s5aroPpsC
fJDqjFPQcH4sttbUhIw6mGqRL5MFSRrbc7lsa+GWfAwv88yIs0Vabiq0SPHnnHtR
cnShaZqenjo9ZdGclo7vjjEpoLJvyBWU3hQVedYRYqS8CiJnVVPORAqbeX06N85k
ogi24pJ4PDoQuSksZwHZ/UWgqgoeiZagIlVdGw8ezlN5+MaygN36ZZHFKlNOBVnk
BvB2U34zwNsTswPJHtacd7LZRiCiYn82cBSocla3DDetWQ/y9FP8xFzNAQciBa+G
sq3hRjCzj60S4hFx3G+/eCdS7E7scPoDG3qqdqf7w5grHmHymGMBsvxYvphDc+aa
5vJAEy4o77D/tdHe17UiU3CXCELRHmjiFCZBDYLn3m11p5bedPELdvgyxMHORcAu
/53jvm2pYk357VHU3/PppdfVZQL7DQmBsYxcvR3uIJfy3tiOAUwjkZP+sQaMAjM6
ObBDS2nij7zOBdb97lBBiSu/TUom/WUbJblMzJjElPI10Ai9msSiAk9KiDuRiOBI
2xBX2bJS+cU1JeRyfoLjFuYPmBJUFtCKEer5bf6NvjxnDoniJC0M93UNAWGA0XeQ
QHoTS3K77jHV6Ke3HoYZT2GUDCZk0qmtNwNvTGELeeNifF1EFvp7yP0izQV6LEXn
8X06HyPcHtEwF29DATap5LP9cuMImwYFnLVEBeQpYVbdfTCagiyUfOUn3WRuniwx
t7F/Sk2VByY73WFnWyuLHMxvLzEuKpmEX3100ww3rRhENKK/s2S+oFbA9/44+3J2
lySUM8ichSKTibiOR5GsvvKnK6Dv/aRcZIo9Dzt68Asnvg4vOj3jXvXChlDpl1Ly
vsz/r4Q1EOSxVF9YSgsM0EtrRHN/qvIpKEOCD2S5Pn9F+HHknVInplUNQlm/3qte
k6oyb4LsboeZzou0+SVcCUBVRqPK4x1MWmwSJOHeMbtvLHoSg95vGa/8f9O+OcGn
5g8PYYYpwUSgVvwvTKFroZT1//xhE3R/J8klI6hUSsVnVh1OuUo63vNhs18B/M84
KCL3WBg5LLwNHZtFUtA4IviP+u803kDqgUI15sgkf0Klj8mx0CLqZ77YoeWeE4bu
rqhlR94gDkGZ+kr16WEYY0xm2h1/WCseNCm4gPOUR5DPPwHAob9Ia8J+7PpHtuzF
SnuD1bdRHjnvx3IxbU/ZNciNsjuSMehGEBKvuMo8zf5dqPVuibTRLxnz0oZeaCwk
+KsJxvdfhrVZANluXfV9vGxKqzsBXuNKgTKWETX0RZLf7LzEZOOfe51tJo4VL3H8
ZsQymkSjj7AHbm5hdQ31z72QbSUwKd90i+XxR/O4HY7wmJ815l37dMaFIN+MvS+5
Q/5fMYBy/mO9WYyE1W9fbdGZzPxutQNYnazzRrtjYWhoOQrHSbxpP3anEwrjfiA6
9xHwAKmqAdy6D1xZMhQVXumujGSnO7QUez39x7iH7lCR+ojD+P0sq4v9oKWTe7NW
jQKYCDvUv71EbbSD7z2Hpt9pzLZL1iNe2mGeJhhBx0HBFx79TRq/a2Yh9zTuvz2P
mu5P2LAS+zT9UaSqo0QjWsw4tHVJNjHeANlxvPj8LHiyDKP5JoIiheKVVvI365nE
J8JpSNrhfU0lvJmkBZKRG7TyQI/2NuA43FUSnFjhnd9ugncROTRDq4OA/f3g2YCZ
OXKH6nMV+toONyU0F03giQeNfwZAAjDzNPMqxUjSuoUwk9Vom29LGQi4k9usLz1X
nSmsT5yp8/N5EPY9aS5JnlBarSNPUwN2Zr8aGoNAGfOOGQG99GWtQnFXOpymiMLj
wA5mG9ku6Ep4UDlk1elo0AwXxCu3CegxL/XGF1ZsRyhWcPAxZLSgqGGIZxb2+SR+
XwMkgREm4Gly2CJYpXbsvw85RqC72lVWHFnoyakfYeve6zKEoK5uf6zQ7/bXdrna
/dN8oLYEP4WK5elkTRWJA30ynXlxqbm3HRSBvN/a4jhDQGW/jZDyEP/AUZITaM0k
8bMEEQNYw8dVfvrG5MtERZ+3UnR3Oh7o4opdtLsEV7Sz6Yr/7AnHWUsgfLHCXQjo
pDBu+V71pHzSxLOzpXCH+nKXN3GyOKeRUEcC32LlAWVGrMejEQcZGorjtpd1ehI4
BzMDrtjifQ8ZQRsWvxK8Miaa+IWcPgMX92GrAX+5BugL5jVtCi1nJ94hkHlALZWW
Zq0oz/293ck3906xLqd7Y02SPLdjtVObq1nPr3C4V6BnqHyGwmR+SnI2SRQyc/TQ
68CCf2+y9mSFSsIT071EEiI2EjDbFW1NqISG3kDFv8aqwcjve6fsGj6wneU9GgYQ
00nmnycMe9QnyTNWP6DAN6/SOb0Sxi9+WItKTP04rHHV7+A5EXEkj8tkQ8c1vk7v
lFbwQyT4HKkRKy5lreLWJf2XXArxo3XcbxmhwQ4/aKXC3szDrSAOlD/BrGIgdmV7
spBC/kwfzqikPvCQ10exb3ln+Pk+uv3A9lhiamMoBfcmy8lWqwHsRqp+cbSPyzSY
3EmTmjSakkhj4qyVRYTQJSX+LH7tpDL7AOl4+/UxdofZMc4yfwEVqmuKqZl8L+gj
GAzHEAwf0D/3wDQAtzWDazLI7/E2JGCpTU8AYPGv4G7c6f/1HRbFYWDyZutTCHrb
01Rbh3ycvTjfK3rgNzuqGgJxYjQV2cDjjNXw788tnyC04/+9yWuDEcgwpoCAQPM5
LY04/kU8d0AKEuHDlmm27D1ld9Umxkf+h0nJvQgBb7NFAZ8+SJLtJ7+jZ/7OzOab
nVHvumW2HkOfu5Zqe0arh+E8TnbmnxK+Y9WzzjXRWvazh0lok1tU2kTQJHdTd55v
vq9McIybNO6uWcpqVGpSkCBhJoQtpya738tcrCHryYQZeFCzzvRLBVr1x1DnMax2
hN3xCl+9F1ZjkoBNVsR8oO+hipB6mbLlVLaOf1Du5QHSWVSZZsSKDftH9IQY/wFn
ZsABVD1TXv3X1XC/lly+XRilz72xNul1MdPpf/DxXRhcrnTqVYMtjjQZr0tT6en8
uZj39JecNrKWhQZSpc/UvITpwE/ViXmmONdQ9Ks/vKdUwRrENTpMx/rOHgU36Nx4
kFba3hBLYj0zgxVfkK23MtTT5YbfHG7aKEaethy2kEq1EyVofA3/9c9LOQudNXC6
8ejr5kDHKl0eTEDNZGZoGE7aWaJld6zUHx3Tvl5zuUbW6uR5oXEbqY3Z3u5lWI7B
aRsgZStkQoOovVEd8UHkD+5OihXxs7x2m/3nEt4kWiNSyk82RFr4MEMghkp9wzMr
LVtwGKV6GbadcS7eDOs95IZp2ZRgI0n9w/wYd7bEfnye8MfDI62kpCWlgd1T+TAS
NE3Zv1tCkIlD1mK8dVDvWoTmEGCRvrbQrOurklKFahhh9edhb7yjTWZetYz4obDt
szSej31GSIVYxj7PkINxL4PJfKv5iRzpgpRYIKPG4EQBnk3tT8RkVPBO8/M4Ys13
7MUzDK8GO+2GEgF1dzcpzXaCT/3a1E+zDleKLq0CEJe/CedW8m2mUOC8Nov8LXfE
EgPoEUuM6SWwu3DD8Uimdttio4V80ZhrdDXtTeUip/fTXbUik0nuJSQx6a/qPvZh
r9dZp9x6HTAJ7J3dFGr824BxIYb03/wzNsG9Zw9SFw6Zuq9ud7XjUAY0ZpUSLxA7
DY1bg7LgRumQv+WAY9DECZ4fjgpuoq7Ttu+udAVrbUG03hGIgCKSPGQqxI7DprD1
WTfkm05s3vTNoA9QmkhAZssNiEygIp84qSeuR5cY3HCl2U9G25Iobb2QTyHnJgQ+
Q8epzM/3/tulZ0TXtNoRKOjCEr3WhPOauWPdlYGPEQd8Oh7yKZaL/KBLSHP3Z8gV
0vZva14Mw9tIokhPyifIb5UqZOJkyfy9u/fB7kerwuCf7OnT8ofq5Xwdne/7yv0/
LucvaIH7qo5e35OG72BBPZSgT5M0aA2av3L51IyVzBBCP4yUZV14VSajKBeMa4v1
NDSJjeiZ3duViVI3nQD6LFjEk8nb04Z46ej0On1UlGqkwi5U3jEbsHE7qkqZHnH7
DdOpEnb2FH16ZqYqRP0w06jrY2d5ilyJxK8TLOeIi8IyXnmD8R5+9qRJdEUyQ9SH
6CT2uGTqvyIP+LEoyann8rPeD3l8s2Lc2p0RDZFgH9a4+TIgys6O0oM7k5CVIDCa
vRsFZCMKu79p1ppud3MT/Z4MSlrPsNGFppwtlYdnq0aSRC2zJihnnmn3H2d5u37M
Iwj7IOPaaxDd4skni1oXZ2oS40KnWeLV75iaJ13LrEN0WH2GHOhaCtgjn9WIBMbO
pdHNLG5woe6249U7CYi3i6vretLiBNXfFwmaalOY+w/h8gzM2JVWAzgYoqdwraxt
Flo/c56ZQ0odJaetMtvNM91FdNAjfPR6CCS/LxdFdHI9QpKW1FzSiyLm7S2lhdqT
lMLVfVJl5NHJmdBbfI4v9osAR1BtwyM0Xe5OtobbHXDqDYaHgjx2JJnTppqa6F2y
TKaXcUhdevnp8Maxk9bv8EO8PnokIhDgYapaYu8FshTlje8uS9+E4KLezy65ZLgf
F83udMv7Y+KEj6HWfFH+K2Z0KGulrK31LJJf5iMHGuPy/4tJuaZO3y0KdciwDcCW
Tl1W7h8qV/+SxZmnMIgX/lxCy3aJL1aTkQhGWRTiWODo8NoK45PgiSBFAt3FbTBs
qMF45/kiOtu34oVJ+yYJewRE5H0HFUtKEBpjht2gd1yF+xvuXgm5h+Y28UeLhLaZ
g8fDlNxHhSrzuELU2qQFUb4jDE74lkoT6xWYUftVOTSx/sWvbCHUAlBOSTbY3lRE
F1x5Vx9+tZXMgPAqBvEO3rtr59f8078VasMhHQwGdN2cMPfHq3L9/IY7p0HTXgmX
xs8XDdGcBEEZ+TG6M09tYvm5BXcytkMajZD5QPhfZ95dkyGy+j1TCIOLz/NXbBrs
L2CKJvXRL/jO+XInUbQHmcZ1aQUJc1if2uCjqhePJcJ2TDfSJx30MLu45egc5r/2
PLsuHztfmmyTEJn69Lw7rouXAiWEHFvAdj0iw+CwXxvI14ycluOJwC9Hzj8euo+m
VwSlGRLJIjZoX9A84iOUcX1zqVsrE/D/D1y0bQzICFWKt+WVRG+0r3nZkQcGFX/Z
KhQ8TVMMXYVGqkrVEr0/fuQ0M6J8yxa7IFDr4v0OIB45Kt3lPpoKeP/C/morjqRc
Ls+E2e3pc9xI1W1tcF09ehrYyYZsJC3ubUwOdVCtsVsnj500bvlRC1dy0Z1emVtJ
+bvzLiA8hURPbqWLfD1uh0xG5YtF7OsyXQbuv4i+FJCZs4A/P5th5RYz5rCODbs0
5NAvG4YD1KhBtFSIaNmRi7rlty1X3kucWoSRhO/HhJvK36APqrfn5IdFFuA3deJv
zI+cjOylvYO+WYEVF+3tjWu4CO2oA+WWJ7wCSmcmejFEBqk5EsE4AovHKEHW+Sa9
q8ITZfbRNmWtnifv3gz4mOsB0651AY1UMz+S+btos+e9eZzTYGkKe6qMGdN91GHX
IAkl9h3G9IMfX3hsZEq9MFe7wl28rKF0qowqTjsw19yL93Kzc7U6AdN65waxMTeW
hxQ2Q4CvakeU2hVwmT1PzlmrGUQJqufEd+nkd2Q8WSW3hfC3uy/o2jtr7WCF47rV
r5+6suJ7arfqHb7WV8uQNx5SZWrFQc9acbTV/nad0cLtISHu3OlDrPsi27UgsrcD
cT5JCd6UW92r8UNWmH3PPZ9YxL+l7wPgSMPMoBy/RxKkeK7U+9lluD+k5z6hGok6
hSusz3plCb+LCRshAShi4SswXt1jeGt06BZC/PRBo06WNEeXuvmwnBtw+ASIxAi0
QB7Qau7qCRTMhnPo+vGApV2q9V5Z5Nr4WX7+plakliNhIowXMMoFo2e2vhs2GcaT
jKIAK2WRslLoqNR2WBkaH2uJqDTJly4baCvS7IIADqgU1ZRAORQ97qiTU3gfiDTc
nhD1o4o5kGNL5lUKmCWqfpZSzvZW1l5nvh7Eu584QUr5lz743SXdgalgc1L86/kE
J9qm8bIiRN+UGWDiWyroJEygO5NX1nZo2xog8Xti2lLeFdoCsd8XEeohnObfxUTC
/KCs4w2HHPd2lI/moS843JG5BaojH376clmPw7ppyhnoQ4eWkChqauGIBOEBzjqw
dBA+39CE8kLuO738ybtH0u/yuNUAGzm7C6CuYptmP3ZZ3jNTTLxZ+SJ4OPEYzEHk
RjgmAyvmFJNazwubP0sHDxvhoz7AZuNph6uAIs0SvNxj/DQq8+u3xZ8C5XLPTqJH
M7Y8rkiGxjTEwFq0tkPxk19upRYWShzoMbKDMgl1KaAGnI9XmTdd0NsWNw+/1HWk
mXQMnl/lzqXyizW7U7ziNdo+rwwoKHb+mDHul9SIIiu8unOKQr5QviCdJdweMmKW
fpvkWbE0QgIZQ3HKF33OVc7g/zZCMFf76+UbJeNUw+rhJ2gkSftGTfdrPSHa6LZB
nBSgK99UCxNCV1VnEYYrP7aMkUh89c7chX5mWuKe8hPRbsZw8dyNsexce9luKjUt
VYCmey5e5nP62SjYL9jxYPjc41Hw95s1BjV4GPxuF+KxkADKOxOs/l9zm3lPSAMN
2/WmslLOeYTubkd0pzmyUMw28WgNeY0Z8tWjIR9McwZmtpHuz51n4IhBhpEK0Uo5
o1X03JGw4GbGmqjK67hrzZSt0C/EIZIuv8aw3sS80E5GNjqWKzvaOpS6g7C9WjUZ
ElVsp+fRrteQLQ0D1Jf1OaSvuO+DMERZdZTJzoJuSgmBk3trx5K4iSQjx58KEVpZ
0LhkPihGZQ0FicxfDcXqkzkxJEWqefdFBwTk+9yEU6i0i+iFOy1Wu4vUL5qNDRb+
rd4uodWRADHk756C1I5cIWG7eXQMr9ecJU4VRaap29Yq4He+10c9GamGHRSKpxLj
ebOpArJuhMNkHawf8/3mDA8so9W7hkNPqZg6ZA4Sx4ePSA928/hfptmzD66XBYVZ
zeux3Isw4ZNoGQWFeGtzv1ocb03SLyXhKnFXBeZBzVnn0eC1GuqXHXdwTUPWBwxl
sI/73Hf5D6/X4xIb3u+2VOidsVpzGwsInjhzlui1A/S3rh2EyDscLZBHQQ69EFQP
d4wlGHYA24xlQV6TY1x8BCB1u1DXu7HUU6UC78MC23foPMVCNRULZ8sv/YfrDHiL
6zBxRzdGaB4mb8ReYXuWqEsTvCWH/tL0EcSWR6fURQRDcUzOR5bgDqIf9dMl7D4G
O0WR5ylYZc6IUbr+u2MtTFcAxIYEjt5OAabLSVvm/jEuMz2E0c4Me4KzSLnhZ5ZV
lNJeZyik8vyhnHm6mKOshKmCIWrfW1cYtBOmMzEN7D+zkJbyRB11BBkIbgcpgjsU
wn+pq0beVEF2Mdq3ni18/fn5xMbXudGtlDU9s76lL8GZaV/7UDI3fXbll9JGE4t+
v9f7fMn8wJwYe3keLGEb0h+HbbkRhuAadL9cb9qs7JS6GcP/uRiNqZ2wGlxwUMQ8
QKpVthY1ZynF2LM97NQ5DjNAeccp/BMIfXbSMzLFyEADaoCWgUnzSOnotgCl4KDT
mnMVxyoUSWY62kW0yHXpkpOAhUnEigfg3q07cymLTObY+799c/hdoCtUCERBkzNX
pJb5K+SHZNeVxH56uSJbTzWacjUVcqdG9h4kqx130pBBtpIsfycYG2IDJ0fJZBpe
iItnLlDl1ETld8TnV/CCl6DCrggzEKFrRy48a1ospwt4L5MCNmJQkhRGS7lKepEa
yhVmRAu8Fd0PnETspOIJzpUIYhY66QpST+s4szo/Ti6wGYhAvnE1Q1qCPNMIaDif
G3Qid9EKLNp9B0Av9CfXiZQ3ofkX3H9MxYlXfrksstPnCV0ZK7Vz7wljgnqWwlho
opYoAlt9K3RDECLobL6XE6jrByo5MFCJljNdhF9toXxfO69rAH3A/j9XhGKyUcyF
2lktByF02AnMOitVBP1mZN1wvKdh1lHKPUq4+ZVlZa1EyN8H3i+iIld7zLY+hnNm
smNNkEnFIjco/j/GEX3GhksE3EGppqFW5JWaaigGjPa5E9IrBVHvYCLHd893aCss
T7O2cLS/dQMYS/K8PnEp7ogMfvykqzFXP9ZY+eqnRaECP/9zdu8KiFUu4rwL9W90
R3IEAE3mXST61myljkkLoemmJ5Q7Yv2SHSuVU+Lar38uzTtud9RILvxv7DkyoJ6y
I2hn4b2DwTQRHpsSe/mPEYdCQwKuQcsKdJkraGm+1/z6Q1ESFmKQwufAP6JI8wx/
db+KL+3Co2KL3Hulyeg3HoeU9UvBirYgBOgfcihpCxcRuqdK8VQ+Iy2gRSWNy6P+
vy1DRcAdXlaZ/estd1eEe/+39ZKMcnQFK8rJwTlyCgQbJrCz9FOgCAAfIMwfbCCS
lTBeBxstmyYkD0LiZB7Ue9xzKJt7c9AXp2+ERtTVgvXnP5qg3oD4Q9f4BMwyhPk6
JZTGLCCdCCG/UWM0BLVWpy8nrE6SUS/4dpo3L9aF0jUNByFvwkQLEYqeyqAOqOe4
0pbSvrrWuVE+iXef1F+Bb9tPCXRV6xEhIUAZR/SRx5SrcD3+l2etI4SNtAXKNmN4
AWOPSZFQkuyKMwivPLfuqIBuGgglyCQmw4P00X5y3f0ROe3vZlgGqMl3HEzy5yn1
qBUHNKRobbxT4Ths90Sg8czzblJmt9j5sC7fzdV4SLCqulMRngIFNiDmTvzelLYH
pHGF/B0RrzfI2KpQXJ2OJr4THO0I3YWx3UifuI2g6G0KuALymOoGht0jg1w0KIip
OjVAgchBYwC331uJnYfDjOAL7a5xoDB4tatdgO21DG9TE9jQbLSoWUizwcxQNqgv
/TDO04ObT+62/EB42rQPdoWK8eb0RbVk2GwTX7MNj1ritBcGEeydcEPrxvIjMZIi
f7uRbgJb3i6F5Yh1OMQIOckIWhRVws8RE9ezmHQuoSf1nrsHEJsJCdWp9IXdyCLA
aufA8CjoKmk2JgPtcI+FfJEtW5A8QXNZ4gf/JEppvJEHBPbXidsZj6oKh2WngYj/
WVCUt2mwFjARCHpEBF4P2EgAV1G8bzuiBZ9M9PJAxU4At+dsztXRw6nI74Lhg6Rg
bPmZ664TEVlcHHGO7pb/SjMDdaXcdLqwr/KLUb8lMA7L7mN3TdSBIMh2WeOEom6i
xYrYlr6Xk4yNtaOfHx258dROycv3SJOgj1EYsrblSeHi2M+feHHzNrafSCHIfgGX
aB419Tb84w7WZhkE8fIoGBc2EQK+iDxc6iemVY74++73dpEEn3ZIC/Lx3gT3gH8B
4QJUn+RKfoOXj6uY1PFyaPgpcmClL4xoimwNC1R3WV7h9vh5xiZHWjugacrMAIXr
PiE29j2ZISTnPvt6buoUlipt3r8q9MpB8vlA48VDgWyeMYp46EaLGJfQw7Xm3bgG
z6djohUZgvOGqRWVr5w8o22qk//PAMArTbwOCVo5EdYpCvZW6Dx75CQsscsDbQ5u
GgQsnK/s+dOxq7sH3e0FaTZAm18g7iO3xfo5X74nLR9Cuzn05b34oDV+CzABJILX
+EM4nwZTeipUw1fVQtyVUxhWTMaU7XKx5VaVEGNjInBpGDOJ16aL5CPl1Z05t/mr
0MnvVQq0ITS7sYMuY0/dwr1neh5EiahvXz7Vmn9pUHT2ZFjQR91kDa1+nKpUz6jN
0Vfyg27+FYEcK8YpPiU6wF43fULAIJMSjhrvhJ6HbC4+bGuBT2BRJ0SLljUi6KZS
uw3ZqrK5dxdIWFv45q9S4yuyiE8wy6trg5qd0klnOYzm7Wo9Y161yPlTw3/TNvai
hvmBUFwb4dJXfmydr7U83lRS39grsd+Lc0R6ZOzVML6clCJ8fJ59r/m5zSrMaXVZ
wPjehvTsId8X45/hgBA3e4CbExL1ZAC6IGY/DbJ91c17PXqtlKQ36y/QhCALHKEd
QyENyTwT5k/r/4g4hIrdPfUpiBPsRnSxpEMHZ2721YG7P0IZFTFDxYLUXS8Dt2Me
xs0dX8f/6uLQqKWm83z7V7w7XncRKKLI7x+i4Uio5H60b8IFbF59sxPQyqom4c7N
Qo0LVTJUH4rPr255a54lSeB/XYtryBXXLiA5bZaxTKZjdktibTZxQUHonQzd9HaX
PxJsOJMC7Kjny5bzms6XUEGLg6nK3O2a7rxL4qM/7k8D5vaH6L2cVMN2UWSf5eNs
pKPKhbtS5FC/X6sADsJP5uFyONAkdzSyEWV5X+OlImLm7x+nkF/WbKVXWKusREG3
yGi/BoRdTxP9qpyJTZa9aDYmqUF+Tc9n5uzqyCtovZU8cf2/9yfLM4dLUA/+0GzB
l0f94kVFbukNqF0E7rzb49I9KUZqs2im4fU+EAw3DMq4bRdqVRpWWi57m7Gmrj2w
JNyyhg+RTw0Qd5g1r5mmzzVdGXMJvvdup4AdEgd67AwYeYln6Xop2MU4wRq0t7Yv
uTuIxPcaOxS5+NHKddz8tFtXJIxl28OWksyQ8h4IJ0xNyPCbWarQNsZy0N+b/wgV
OJxXjk+TZ2jYFqayxxaKeiODI0GKnbaJfWhRUys3UivLGa3u/8AzTeeiVskkrcaS
SrkQc4L7RBDR98aQTvFdmROzVDUdRaf8BnKFbxfX4f5e2L2FX9Gf6xcIePFX21KZ
6S1EPa1IStY0jIBHD7l2mp3t8kWEc6DXHNInddojezvzfli9qfilI2bEp5T5XcDQ
Qvo/qwoY5dPDOflSeWMQEQH54JXIktol0ATXe8i99C8uEjVQrJSE18ouwTxe2ERN
8QXpPyPOMeEPsQ6roQQ5jlTw7uesEN6KiIhzgS0a9KgIfGs2K+zPbIm0gqhjJJi8
Kv5ar/2gc+qGW9OGNMQpvPxft4wuCGBm4DkVueY5KNEnVBG4eE3z/NyAXjUdRxPg
oFn+O9dZnPppMaaoeHnVnN/53Mp7sC1MkOa6OnBLSloWeCn34ud13Mr8uwNziTzK
Hgw9WAlFbsXwJHf9mDP6Xe5K47wHsMib454EqNoCp4ZJeULwDy5+5ECI5f9a2gTw
G4bX6YOAfvVpN+461MESLtF9NAWvxaaLMkCixowlZ4x7aNPsuUaQZjqer7CHZGvj
/7Acu5RPhw+tysVvvscX/l446NPUtWVD5ZMVonBHxYkM2EnO+JDR5ceG/ReK0uMR
JQ8wBSaSROzvX1XcvnvbppYzKdNL7fn0vHmtEEKldZrc/LyD/UVhJWXgnMSbJBT1
fV8oDvOLOFgBfQxXReYMQbyrk/bwpejMjJweT5lfwII089RyOnFyxcUK3DmolfGg
MOnvO3Hibu6/Z9CtPjC6bS5Ek0EzPOJqE9kaUGdk89Ytc0dmjWzpCi4bMvk+IpIE
QOSAdd/k6uh7jKJh8ldXERFJ2iY+J7V5L7vtwt6MYzor0Z89EgIUbMtrFVQqQMvJ
Kw/y/9kI3++DaSBdFlGZekUkqHa3NPBdz5iAHQoTn0RWQkZ7MEdHQwCTEBscr8pN
r5WJ/bQR3X1Bt12UskqG3aKtvVQcv0eqWdJDYHPvUY8F1kajAy9foqrF/T9VYG4t
vGomWRYY1H24cGxAe6R2SY5k5gLm0HsXuD2OplGjImSf2yBCRKvJbqUek9l5tOQq
c4Cia+eAcT5uDDtA8FVU5l8kHCk4Uty67coslMq+ceBWg+aiuBin16Xl//gSIm0U
br3WKk0EpoXeZ5D1dZZqCDsYt25kRKTepF4SIXgy6K/p6WSMWvsUKROiWmcZ+F4h
iIzTX5hHfYVw753zwIaPw5W/tVt6+Up7anZYC1dF+/0jB9LuGoatVjesSTwHfcz1
HkQSsfBAq+TUPUR8adF/rHlKUvdFV77xPGMFNzhX5A3u6Nty5NLLBvklNYPbT7ei
1CWeH+n4SG0A4Gx5iyaV0dLpD1jwkKtTBsyMDGjc4jhb5QuaRxG3PWBAsAzNhggx
QD4MI/kGO+xaEXQ6H9T1GSy4qTlKv8vhXnza+Qr+UASUG6YQ/C5P4kOMzz+S2V7/
uakZPhoSH9TyK6jjZSC15PQggDEAWF4uS7ep/fLtyEgTkqqPsla/GIWyLCKXhjXl
NDeIv90MKcIiN3mzYWzIsJUbVZ4DhbGFsCAV+MRz8pZepKY35xqMb/rjaVbXeEZK
0ZfCWnMoB2iFg3OsZAN7N8qTWL3SVPYkjWZsbRGDZC1tVGgpN5mXSQqA9KgxPrLc
KyE6Hp+ICW6i5gvP0k9vszWjgUCErz313ruo9t1VBfAzx8IbLkC22PmrkNYNFL7q
lO2fKk2UGaQPT4/0LHETVJy+4gTRHhDNk+N+9IjbkjdKZ4lFdfFgRA33fxam3C5Q
o4T0Ii66Z+S4PXiqkpiM5V9gyih76jrAZ2bCgevbOBGxdwnET1xwA8pd/Z4Q5wI4
W1frWI5/AoOGMNRF44Y96tE60GqZQqzhWCPG8bBn1W4SwfCet5ldSDOOQ/n95fr9
A+av2ypn8oldXFJespRdQNorIy+i1CEnrFSxd9G/58UMg7AwBNYQzcEn5L7A8Yxm
QVDPw5hPRGBiLan45F8oGsgrAI3dy2EwjtfmSCg685HRijpWJ2wmcoW2MRxbBWk8
Ez+xZDfPp+yFRx4ZThrM4YXC2jhueYOpW06LeQ8saAiPwmrVMLV0O1mS/M6tXRiN
5rcXs6HakrPZ2Ds6N+F3YsfKUXKSBLWTqHM/bmon9QbA6b5jJ0J8uGKRVfhtwJrB
7Fy9mcC4A95v93q1xlOt/G5DnCfBZKtIqOnj3jMKtGDrMvS1M528EABzQDJ98605
r0CW0gGdWfznzIEiyr+C4BCnL1E6IUHur9IoPFPWQc5ArhJ7UIN55PgSFxmQhNZi
o5J8OCfKjPmfyCMLbxj4CcCWI54VJLR5vtP71gfwkFna4gSp5VtcxJR4nlLyPzAf
xoUXWfHnE414+PUmpASiTJTiQVeiSM4k71dEwF+7BxsQrxX5OAzsKwnXuPXXhsAX
5VB0ZoOot+EcfAtJQl17ohw2Ijcbmv6S7/BkVbu2MMUOULvRxS4FSum2qQVq5iQp
JqpznOFKeoB1nXx6QFAku2eDzs7DEP/i3HbJORlATKPkElnjqHli2U9A8xkY4rek
SgnjKuLB5srV+/HOVvbq3FRpF95qUB2HT1lhDvpqL+vQlRmMxsFq2NYUpthrbsOF
MH9P8Sf/yqaLzZ5GgieZiLqjn+UxcAyyOieZQuCSnGYk05MfdVpUQ2D/y6oAk5Ii
a9ywOcuVP6RFLVHbixJ1K/7Yzb9fQGqDXz/1hxPqm0ewSvQiv6dixXB0Yj6/FQPC
CH9ezAKXSHYop8e2LYZHyVmBWyLTYrwPVBL3ZPnjGS2Gb79X1wmVLgzCYK7Wy+bc
2pn4AKqDCojGXkaICex5y6X8u5ab9ms4Vy21ZcKf9TVM0SwYUvcJJNWG4/yaY6/B
3g13jdh4q023QnnJM41+hVt431LDqdHCUC26pBE4SYDKD8jLqSKFi8hnCFowECTm
tv8Ro+QAp2CaIzTtrSu9Ed1BnM2VyMwNwfWSEdChg+fGg1ljLKb+0PeSiabfv+/6
kRmH0n8pmmh0dkmgB5dboabvtkfwWw1Mabh04Y61+3X9vd4lxdC7kFikaUgQbaGv
HTbSGE38PgaXgegcU6hO/G2dpaC9BgfrDasDIgUcaSUpeVhyCDjK8/4o3Dm+W6me
dfqPqrPf120NBQQyZ8RCz8CPy5xz2AxnJW448LOKqFxHwyNVhcWguZGEBa2+UBBG
8bXqqXtu46KArWb/kE4/8r1w77WVhrBUt2ZRYfnoN/o9W1Rhke7RkvmJszi/vCPe
vPPrm7UHuOgCZyM+We6x/i3elN2jurQrMOSImcSY282/FuUg3njLYrQsuKDyy5FD
qsQrqAPxfCndHiGVVGZKJs/3cfgd0zF0n5NJX4ngaJPnsn6xXTP58sd5IU0KnyMK
5QvRiC1inUfI0XnGBLlgqlXMgayQ3jzOnLfeJr2zL7tRjnTtbfwtxX5qys4gem6S
n9ujHcS49CdrrQcBp6n7sRNCNIE1uP/80OVkjZTQ/PhAcb0QiXYfcuEgJ7I9hXg7
RCT2kPU1EAJ6A6ljqM4Cf67LGyyA7B/3Y0d6GMaJzaDlWj599y1I7Yl5Azx3mSjO
AWZcIlQ499f93KnF/CFm+X+rsRYunSfZ81KE3O49lIcn8r+yfogR0CKy6lhW5dUP
xfspOfe7HOVVRbmJUi4hnvtMKKhdl/c2cEpsx8D4zfkXwN0r7b8POl98Y7AZrnh2
cnmmHlV4MyXfEOeM73vCqRRk/RUJBZB89fK1zvg1DiwZ8t8PhOC1FlE46n9kAseq
IrkaErPGYzfOU/8OR3OludYkmHsz2Dqrokmhvuy2q7h3CVwAO3iLe+wMKEeG6s1x
EeiV0tt14Bo0STGgrfPXAPAlPYfhpwxDARxrRwypIn2TyPeBvXlcGkRnl6t93XWw
Pntqh6fkV9zR7OoUNKZ9wWv76exfeC8SM9/B8ElQRHJTNzqSuCon5deL5rdmSuwp
LPw2Y8DS/irRk7a7cM6bz6gFEur7txD9r9yc125brga6fcT6u7bkjN/8ycVKPKVh
TwR+aqNrWqnqW7rDiQCfzJtsG0bum+MykPh9w8RV7lA+RIuhqdJrf7OrZYIiQ1nx
VtpZ1YZZYe4viIOZL0xwe4oE8te1vDrzDnGSuVSI3SVpZu7GKrJGiSRNHR6CxiTZ
w26UPGvCB9X3EMmSXJ2YaM31jT7gk5gX7WnfVCiXrplY54a9ieXpswp710ZtrQYp
nu72CcThSCL10gWUoxBpOawuQKIwCzWJbvz+4mGIiab27lhlluPkBpOhAx7urVVD
1RfwhUDffOoeETfdSgNQnKOJ54BBFqw7vcsj+EKs7n5x305TdjJs4Z7FxcvzWv2b
0U1UwomM2ocWzrepkBCUUj+o8iuSJX4ZT5uhgNukVEQstB3VTYLDmg3OjUYxTQxK
xUO6naR3laqms+8llsSkggjuAe8BW8B74XxUWP5q7KrdN0kypfU1WT3nRFenDCPH
kQKPJK8VlCsztuP6PSqzwgOEeQXQG2YB4x0bEmJT1WlaDg0ipEvileYovXPi5Kyu
JZuIo5h+DME0T3M6uHpZL9+VDdrDpIIPfC3a2hOezVN+lIaH7PmKtrVSN4xF/+oB
YCr5tUH6s7gxFaJRSEOU/hPeURCJyCxXnwq99n+MRbcGv6fZWGMnlIqgxQ5py8Gj
2eZjkGhsdVUqtaq/Qy41MuyOWPedeZUW6fV2tzEd9cv068/N00ilSkr06yIolmjQ
b/JtSZX73Lp/pFLaf5LupXowuJECNjOl1c4XdpgGZp/6kivFKcAn5zvtkbyPjnuP
jHjDodTk1dBEYK/NzlcMoqrS1j3UdxERNoiCdEQizSC36xkHAqelipQ2fp7oe+kU
End7P6FhfEw3YVpBYvwVnz/QnS6YbFb/3xKnYFUzFrvieKSGTQz7+D/pWAHhp+7q
E3BOmcFv9sMGjFj0wUXN7AwnvIepFqLq6KaKwmI9KSYqPJ1we9jnIrlgvFVXFpBg
Jb6mveHor6RM132RdT4XtDd1FNkaYafUZxEtE/gSjo1U5VybfuzldJm40ZJulbuj
StwVMDqbXnjx/pGD53EB1H+wt6S/XBxXIit+nZzkUwqNhMfohQzVBCQ5IcCx8Poi
RGA4y7b+CKy9Kn1lijDuknFdZSd4yPlq9nkPCult45n7eJJ761/1/ScNwCEyPWMr
C0Dvv5hm1HV7XpLP79Q3V9tF8xd22WcatGzNC7YxA6lFjfjR1YnULB8PZ8OlyHaV
dajyGa3hIr36Z6K+fPhgw/dLBOo6JeXq2BGOrXt3r4rj+sE6H03khruEcCD0SfAl
Y6zVGlp1CIHgCBN9QIe9oHTHvOfwvL2x3LKxXYrL9fOf+GY5lSM0hcEs+hLBemLS
nwwziUGRUu2+zQdgjVz0tZ1lKo6cYDmtV3kuRbpSaK4/Fh+M8YwZ7PkH/aCrS49n
bvsy1YwQp5AfpM2Xs0b9x/A9aPtHKzLh0x7GKeysCgBZxhAynR4PWT7LeiE2sy77
Eti08nCUJ65uVzUgzqHPMMT4tKW6mrBVL7dIdESOqIWxjilg1WphOkZHT7NZAq2z
MIo9W2ngCMfbRjjMe+7ubsJvHalpOcCqrpAsADNFaIOUZNLL3lH5rx7Xz17KOEfL
ZETpZpm5sNggMCUs9S6ij0KVfXJmdphPpHpli9S5wvtttYjQ5FqA3BFIWrlELWCG
J9PWjYNfGL4BPG9rkf1HujZpOuvWDGTSuFOWNdALftV7171OeAdp0JOvOtQbRjPE
IQysLMmhCAomMeFI0sYTRCf/n0gVzXMmYk9QrgMOKrFrLm5V3FTnr4rAjH4ulD1j
J2dVJf7xyuEgUF0eL2aDPEaFRZtuiMnlGhuTckQqt0AzOvHNOc8SP+IKvDt9TyYQ
5Aac8wbpG03FWr/jnjteGL6BK/lEM8+9LlO7XwLzZfS+i8Tnhg8rw5l4s/i93R4v
DkCc9wzSBE7T09juKBlaksBpSAYq0ZUzC8I8tBTNknN/obz3AU/WNqbJmvf/w8WO
YBSDc/FRkfAhYWX783nds/3mB6+q3B7CBJyzZQxZaCasYJlNmL/f7j7xll8TVHLA
ut0vMWk6Cts7ZiW73NvsEdYcfhdhjyDEIEhzrdk+oDPYe8XXITBRct/4aYsRMz05
XR/NR5NaqOP6sFrJGdchxZnAY5Vh1iPE5s1tgrhLFarW9Zcj3Cqb2BUXvHSB3vx3
bJxapk1Pd25Y0v5/McTZ9beipkNUzadJlTRsX/69ueyhHYpqdM8/Msilq1FS0Ao0
TnnCwK+de72lnJKBsA4F49QC+dCyuaW1OuVqmFVnf1kz1NuhzjEKK1wyBIqJRFm1
TuOnSuqWOyVi35n2bDnVMWZ4Q5cEzXHBTmtyN75s2re4Bsm7K7TxCJr2MbjkukRN
3oE5f1LvPODlm4a0MRMh8ZnPjYjeqEpC7r4HRu+tWlpasAzmbzBMdtxomx/y49Oj
DOomeNXsbJBE0zowdAi+yyIArnqwC4fh4dCi+FT6Baqj6jPwcBygBjGKzqIdRkYl
oJbOUGEH6JyYDU7GFY56sfwjsucBLYaDGW25bOYb1vOlTA54SFLbjRpEW3Wil5Y3
wMuQZE9Y4U5ua4SouRaUA88x1KgDiZoXlgUxzJ7FdxnuHLBZSIcqBBs/mhZoefyB
MakVoPbjG+tHWLAB15NDYAWx94IwdJReiXRLgwaByNWSgBzQyAm5fVIG5Ft4DdzV
h4iQYLXaHATj24YYNraiPOxj7U1FUt3k5HLom2WidDw093NsitFcazSEcAIrl8SY
VueCwCPolWrTuAxQSqwEDsFl85Cc8WRWlKDMZ+iP5E5jm/YBQQR7MaTIeLbHGx5R
7XtuDs6ic1q83DbD8Q3X1+SXifJlWkrdJFFQJaliYxqyXL0dlRvknjpBP2x81M4z
Gkq+4jrUO0Ak3Ixk1LWWERJYbIeHN8bh6IDDn1NzWB0ekYm1tZAE5ufGjAGoJE7Z
oIFa63wdQahXhGaPGNZH1UgxsJLyzuyvDtxGDYXxvSY2MpOZogJHjid8QLwx27BS
ePqDOVAj9ODVkCgouHzBi2HJwl2vBZdrqV6LxBAdyA7s3LR0ikh/MCSQYv74Q3Ey
slewvaVgAcFRMS2mIfbuq3ai4t/zx4HSO4m7vvFalBUcGkx6yQdFEfkAGURQuNZ1
lcSYJevg4G6+Gld7i/sgWVgRY3v9bgsMYpJzp1I2O21nroGtFBOr/3uELKsOO8iS
8gR6SzCq/CHh9XG+kRI/tO/fN9m8jQW+zsU4+z1Uu+JqoKPkcWK4CISVjeMs/igX
fav+L1Zh8ZsgQWouVJ8d6za/vihNnDq7Y7Noud0Dy3PGQdEzJsmsJ5Lze3xDA2He
4xS3XjoHjZRmeaBZea2+lwTixD6KlFytxX2VYS4V7qWwW8KJO+QGX/z7UHc0SxFV
e5Y7B8cob80vqFCzmKr1riDb5OeqTrX3Q0c5KV1AAk4p9D8PxEKYrM2fI0n1e5SG
l+IslKuS0Dm+7OHN+1rsjVVJfVKfOHrcG8gOhZiFrzBGQHJJycQ5OQ2qBRbzmIOV
XCobkZKrxfnNZNovSpMJWHBNhqVdElAv3V3wtx8KEy8zWtLOc1iPr4IUND0ee+3x
pvu0XDrHZiegYIGDLuGJe/h6LZH4X3BkuXVbEhXvxi+VxYe3ppTncDQjAK97wyAR
bYVGHgiO5u6y1Y2QutbIQRJXVAet3d78CS0Ck33NFc7P3kVcxIsicx2+/ZvUKOAI
5h/Zgoi5oSbAoaXKLkWEt6KMeXuFgVGQxPfPdAAxAG93s7/zcRxCs5RtGMo3w80h
02lGqolVT5MxlswOK08BCXfXrsTOXGYi8b/CoSVIFgxD4Nne14yRqLWFk3P1o4Rl
QPiiMyI3AAHJyalA7fCTHO9WgUlryU3clNSbHlPaiT5Uuk+iIgCap5Vmn8ICXUY2
Cat2E1AGKz+56R/3vd0VZ7ydqnUMAFeDAcVMfLhShonXJNkfOBEazEdWiWaNUYc3
wWxtINiGHCPwsa0m3FaWIgFiQQQV5B41+5GgBWS0AP/FFbD1CuY3jwqpFsV5wQwC
c6V3xgonHAeuCLibaIAgx7lRAhMeC1Z5J8GxfEGMAB4c2t+BRAH0xVFSaKBtKV/4
WEDIIwyemzKdarSLLGtVtH3LGwlbgt26bZW6ktZnBy5SSTR92wwx4TkhB5tHM9Wu
OgJ39VUIPCdevMyhwq8gVqNnEhgvEgg3Ubz66EiCo1m5/4uIngYbSvYGCfHVvjeB
CROaPlgMD3DsKu4Ueh/3jPddmp+tRZt9Snd9PsUJEB3iKvj8TM3fP8cDBuPUAtDo
8Ogc4NTIzJEZk2cHrMhnsvpJDQb1HKGVWDwlyByK/VlO6eGE5iJ5hQV+D7hyvR9W
WUrOPrPenTHg0uCQXEVC6RHx1ef94tiSHbH9tg9B9AskEnItoXmIxqYlPDtRLcaF
66Nm2B7da50Bous84dgDOKcLzXY6MkA0dvOyU8LJaJN9WtuXwyO4HFP222tjsJFC
4Kik4bE3VWX8hw/leFJdT4Jx9sSRewozx5pLqRd2QBUUjr3EXhvs59iBr3VDpGS4
vlod6U1MRBv2VYTMpVyvYH0P40ZTdfQTtiDlCdK5JVw5mTiofrVfD6/zHASbgGcD
n3G6KynvKakWEsJGi3Hztgl6OvFc3utVqKXnxdpIEOUTg93z9oO/kJFOFuKC3R58
ECBJ/wFu6l6Gn5NQ/LgRNvhRxPP+P+OfJ2f8a74WYOGJSZdCW/GmQ9KGM2uyGd0o
CaoLSAzXDtK8wr37b5q7TMeE9qw/zHfEt/EbQpti6yurt82XIftiGMxHFMaNDIyq
kezhNb576rrn13Rl+6AjZ4koBtn1gBrCKF+gyEV5BRbkfhK2W2vvj07WbpCsR+1e
XU83wmHW4Lfcf5n1sJ/dM9XecZ1NacgVVCl6/CRHpDe+bp4qH4N0swm0JKupfCHE
oyzEvncNcOIBF5ehCV5I52opps9DZ841b+iVynfftXcWLwjMlhbUfNMtYnifp5SI
+NSqs0krpsJHhBKtMjycDnZ/+Q9a8hdNx0/V/FY94peuHVby7awyddCA/6nlGA+f
2WCSTfFmH1kdqOmVmn2cyfDUCH61ZDmllqQ1DLFXiDFRKM8ZkNuAc4S4gUMsN/cw
EIWqwLWqr8PcY1eY6697l13pfUj5fbwnd/YOdQ6wVOsHepbDXdCq0JZYZlR6dc2G
Id+83YYvzV+gNmSQzx3mS3GEAd674S+wbH+oR8xqVAJ9kn8xzC9dIDUzfH8iEk1G
+yp3a7NYFQ+XbFDBYguDR5uHibIQWpGmdjq+4l/3V8aifd09qX9SWiMjxkPUKsTb
CC1Tj4Oj1E4jviu5pXgQ7+DpjNPwrgV0cc7g0Y4BQ5NEm2dzkOlSfNkV0txiyxE1
MpEyKlSB6fZ40g9daQZfMnwRhUi5Y03pZFafuH3xG8Q63UeEPeuwMZQn1kS0kvpn
snfcxqfBYdb8KhB2UKdCUziOnzOUw70LtnioK2+zKJ8B36E39iKtjvByGEbEdT2N
MkHXUtzN+0WBpf02V2kIPdfR6ggje7Ih4BqPJHNVjh9BZxnDMAJbE+0O1rBnMDgT
k6E5vKC469iuEex2hp9JWnlUOq3/ZClQ2II9gN79AwgDfh611MtyR50GSl638Lxb
8xx97XJsRop4L8Ot0coTzMXIxZrFUF/LZwhkHvWwKnuGd4hOw3QaeBd9ixZWslHk
32/tU923zPfr5SEujhTiGXDYEz/PSB3cI5gALQi9f2VjSU55SzZS8MwgIcba87Yv
YBa6dRzStNJOcVSaxo0nX9VNH63fLJg0Te0lsMtCCqpPC4qbUlel0c9hPfSQTDfP
VqYOROXc6V//DlLCe3yGptJhiRWtCEdkfSU/kqQGSVi4JB8D6+ZKL71t82UpD8v6
7t0dSgnZEa9QiwiF7j750tHzjkeP83C8P+qcBOHjpuR3dgJGIe4ESgmQNxmBL0ec
ELPhsmGHiiaOGJm3Tep5CpmXQxu6riHELb5Ucl0FoF/YRcnPL/waqYG0vqvExPZz
ob3gfJ3h/hyXEN7MaxG+Yv6BT3h3HW4ljwltxptmKsvOzxc46FHV5BU3bzsL3W3w
yhzL3jaKhqP/NZwKp4g7/16Saogxmup5ZWY7iDBJZVBasD2nd9qsVYekNC0XHAKb
uhBqiNjaVQFWHOdEhjX7yQ2yLYmJCKqOeYP/P5W3zKQl9VeCLRtZrincdP6pe/SA
lNpHGsHHKyHYBWV5n04EqT75r2+rC3i2yuFZr/E+8HTlMTz0Jv4hfO4mNEz+KXxJ
bo/TOGJrjU6p5uZIolFP9Dvfq9vRPBa2uIxFaf9tDtO5udEM5O0acSPVA058abCC
eaw7eWMXROx28mUV6H/qiC8GpYn6WvY0IzkSLKrGc+KCUdDg6O6ndgswQVZhF9ur
TXXhCzIVpu0JC0ENdDHY9kbdO6YCM2RsqgkHvvlFt/gF2MafS7hZkBek4B1C+X+C
4qDfoEIC3c6RUxz03TZjhxT2eDAnCYimzj5PJmVyHkLEnzFO2JUlaMQ76PNTkDsw
5Ey1GfVmKwDV8L8PD5OX3Sb7Sy1UQvAu0MV0iAGKJpdWJec7cN8XDQWeAjsbds3W
Ay8nOoiRokI3SRETiFUY70grTTbMLLwW335gFPb1TesqNHavAP5S2qJHvM1QhbSh
e2g8IITPdR3pDsClsWI8q1ejEC1EsaiXcZpvg6uiMw30kjQ7tP/sjMLpjv1DSR/A
ziRPXRwFsnl7KhcipxaUOkOQAX0CQdN5s4I87HsJp3PsJ0MKdtcYpMZilb0KmmyL
8D59lkEuW0JxaNUYokyS+h5bx3BtmrLtyDsC1lrtXT8RKKZs4JJU29ICCvnxGvhv
aw6EiihmP+sO43nR0jIJeU/MHmYzCUFgVMSo6Msp2ipGAjOo1qNeK95F32KM/dNa
2oRA6BZPay/BhloNO8mPW3cVv82DWwr0J77hjciUi9edy3ou3eEOj2B5Kn3olOuD
lFiGSx2qY1NzAqNMqi5vaV2R1vCMBEBuKuNnTHUmtoUYTNK3XSZWG7o/BFiVVz9J
qHjhPXdSRNpf9IjF3D13gBMCfZhtqI7XKWGOu6Z3sZhjz8XRktv0VhoiaFIJxY8n
0bOA2zc8FYtEQKicLzTit5e31xs/Ri6UP0DaHssTi3K5VI9QYNfD8QKy7kiWDYHO
34wcA68PaRacn2Oo4JsBSuJ/2saBXxxkmecTC1S8a5UCTNyUvwTnWt+8xYvzsz6O
wGACaLflTv1KgmoRDadUwKAlmOR0Zay0VMiyyYuS9gcB3JvZErIfLjHjKG8vSDhL
3sC9beR2+2hBGYu73pbBsBbfimqEsgN/KYQWyi5R3kIO9SaarHm6txMVqehgZadB
CT5a2vFuNXxoS9gBLFSnJo2wTQoab/MGkX1kIDUTzpTt61L+8Kx49ubW34mNqnG4
KoYZ6vDTRZeTTs1cyop+3ucKf6k858/6nz/uJ/fA3+A/8T5LG5aTIHK7dgmf6WiI
QuXgq6yvyA30KkGtZpnsNjs/NH910T4GcPiKbs/zCNonY+bOlYbzPTEpF7vZ/9xb
J9Xbr2pKh4aDzKfUwLOBALrdC2WStTRAhCHwmtRuRei9Ac1ENTPX6T61BPTr50FU
KUNZOPfRhQKz2X/KxzqTAPn7BPIqeqEp+DFBSLx8LD9+b0lFJebHWqf4x9rOiYgR
QqD+/yP8zrkrOmXQBn1ZDqTpAqAXkxR/SF0NUyy2SXwaCXNrQc+wwArheG9fwoNz
npRVjKDaxkHoYyFPws9uYImubnQBD7ts1MokEj2SErPFkYIDbcBwX2Ug28otxSZg
ChmEat+ai5o+KJOs4aIQY8NDLJ73j9G8cPmjoT3NAvm7P8yI8hhVkyeLU8FysZZo
mjp8vOa8GhWKpdZVM6r/edpPNu8KTUGSf1wfZj8jfRcP6Q8Dc5rub1i/cnB+qpgh
9wiKCFMTVEIweQNigoKAg9w4NBHbxKM8yEYUGLLBg8pI2SFCcgcM/Z9ST2NNcLUD
YwZ+9dQ1YRNXJPe5/3N4m1SuWo8k+ht864Wymzb1EHFLZGB6/RgzxJS8OjCV2iWx
oYe71k4uUoN3ZlSuDnnRMF1lIlu8vZVDbAE5SCWge9E0taNUgJw8Mv1VSd6h+sUH
NwgvvqybCKFipIXoj5cwZ99RAvIgUhDngkwobvqu2MrhYhCQ0zin6jeVNJma1kR0
80daPAHlbdr7WSkHQhFRK5xoZlqYN+iPm6B8BYfxNEFkwygpqXbWG685NyOGgX8c
g8FcALna3bPsJWRNHOFKb4iFvq6bXfsOZ8EyabqxOsTpikxuYUdS1lvr7F9BdC91
DiWEPCQzcxY4YJ2vXJ8vHHA550jQzmYx/xLWaoUgBPov2J7Nr8qrRo1V35x95/w7
iJSZXctN6mAYAcMDXo5fMcqu9gW16p+LVQCoRBsLXtiz1SsHJF4S+iOEbt5UROvo
uvOrP5dDXNmceOed12ZAzxivKCn5DCsBSGV//yGvUFX9CLfltyIC4FEwmG1Modu7
UO6xLnqaPpugHsavra6gdSp+RNOnn1hfRdoa3VeEi0a7AxlzQMwnISlUvYELIltA
mOAeGKUnFW5FA0I/d/FYZfh/JdhaqDPIx8qEoSfW6PNfyr9xmNZNP1gwi2JgxshO
5bz9lVe3hPOzTEZy1jY5CYL6NhkyOwOKso689TjUh7iGxve4AtD4Ntl02fCFYakj
WEOfEJLO4X0azAdNKSX3LtShE++6b7WsH2rSekrmLe8cciqAmTLeMCOIC3bvqFan
N35jzChUBWLF/bv/5XrSzinRrFkZDVTrFBPjXIp1+702aR/cTq1LSS2HRbVAdCHN
t3pIRJ1i461nrQGoAwg77BR4vAxHGTmn8I2vsXqdVqxclEG5T1lxa1GHY8couR6B
6N6OOxWYxMcoSNkijiy/KxLwBum3e7s3a1Dp2+hHWXHfmzKAASsft3Nn9sLhNQyI
CbI+cISnqQ1Is3x+wCIWaFbo221V32SLmBZjLjcxbldU084/6GAVmdccJkFZfmeZ
xxWc9KdDn4LIJ/72Lgg/HKKC8EEZL9RHbnL1BQfRIDx4eazJuXmnYxnqNJJYx2dY
OzWTaARWdtKewZNiZJZARyIMTpsMgT/P35YHx4+Uxih8LNxs6wf7ug/DWr3un5UK
HYQQmk1BZShzBVjQwHFvcPpp3Vj9BWHjSoIEmmo84oxJciOSo6yRJ7mPmx8y0vvD
24fwrufujQJOR2zafC3I9NZhlyVnh4JE8xkUM1Vo6d+rZ7MIQM0qdUyMCCFKo+AV
AfvXhDWD+1knnndL6sxCWgMhrLozNgaUQz92azFwK2ugJ3lPJ2WI7hxGCyyJI5BX
7KZ5n+dZC0Uqox+8mX+LqBfQzFsmrXQziJapI9V6ayvl8JHvxY1vFjpeW2S4UmFs
bZ3V9A5SiiSbgOSZabE3IBBBVPoz6A+LZoZqgx5Q8uChFGDQSOLe1zbcjn/wK02W
tL/eNGjl4ImUIAduiNEZoAxSE+FDAQxbhkKAD3it0S1NnQhvnp0ZaUeckWpjidaR
SQm4AUFpjtEBTxqDrnL2MW2SJAeYe5V8Zx+yehyj7jPGfXXJUYu5V4hBG1HZis1Y
NLetT0q+K1Fb2Jgrz1de+2I46Iro61zq6w5dRm234CvOhwkwmJeLTbKZWpn++p28
rcOpNyF13MvsJsCr9SCGvxVq1OmLe93XHTV9bLCZbd9b1JtNbI+hn2oQQ7237ruK
L52iitO8McZ1R/mijhJ8WGa5YkoAXkfVLnAytA/FbapsW9BsmuhgC4ExKTa0/HzU
ny4+OxlvFsLfsEGRUvXb4eq30gRiHr37tu9CIsS6Qo7OcA67rbAcFyjHZpvG+2kH
Jrp9Qk2F18iAKkSjCL7mbJpkc1bpNiqY+MbYkBzfFF25zTn8ZjrUg0P7dJTJMUxu
+ukJR3DJhrLXxXl+4yzqMHi6tkmASiwQUCFwfiokpIQOAEeqpVrXT2LnZ6vM9+t6
0pjHBNYKCfpIcnFGqhzziOZ55eTz6cMPEXRTIRiL0tMfHV/KZZMukIINmOer0WBi
HD7Pj0qsF7svVxR4Y+iJ1xznJ5kfjZJiHW+52/YA/cA45qnaTtvHfmMq78O7XOom
lG4PLVqw57cGZ1FHKCb7mSBo78V4DGCcYJ1FrKlNQedcnVV2KUVUuU2jUX1XpGDn
diy2mT3ExrxdAZXSGzd0eOaU9qmFpFHUU/zUW3u1HbMoMqRqeB/BWJ3FmHuJJWpV
m6QYntczysiqyVxiXwfY7pghRWp7fKeup0PokZWLfgIJEEcdv02Y4fHfajMwmcoM
TuUEdfiBnVXoyqEOK+35owcYm5yvgPUGdU3lmHIQjxaDoe+h4I3C8/k9qE95+hHx
IoHOLc3yqAAlpMJZbLdxRV2yEL7Kz8kLhXMIF+/Yhhrg8Vfaf32RJeBRsdeX9AG9
J4s+rc9ZmV6LfFUlGSnYXOu6K4U7/oga38jHGKWUtua+UGffFdKJ836y49VXxHRs
aN5soOWgZskBCSEKexWtYeVZJi77NpRNkzkxL3i7U6nafnTVTv69Y1R6QEbMOXZN
viUut9fsEyl8NiBrxt9Z3MNCm9Ir2sxxdH5ozPDqRUJkHqEUgRQD9Ymy5tugSlX4
3P2y7H4RtA0NghcKKoU9SUIywE2cVmURDN9WY5yu400XtDX0KDQ50yLeTE1Cn3ev
lHRNXrE8erapeRejKqHlvFaVbbxBJwjli5q2NvZv0o+EEqkJOn+OvNs2wETdKIK3
7SYFPw8YeHIr0I0QHSN45fL4jA0/cAaOI62MKom58EK932fqYZ6gZREKySf5x+ZC
GEiPJsaV++A6mI+496DNdxTspmNReHBCDcSN1YQTZyKWUKLhptuBEOWfexDR5M47
U7B3akhAOVth+852b5J7jFzCoEi06LfW5i8Z8Mn606V+vjvPktOsBCi0yyIdlrhU
G5V5R33Yw3Hxoa/rDPiFgXFcfVId4EeY024+PASz0FJLcSmxlxnilRT0l9RpmmUl
Bbp/Ck02A5aG1EPkxX5bR7B0V1/33k8m7vrOZvfYk69dzMUECS3J5fTdYECCr8uV
BNVIY49nh7k/HiSkNNTjnluF3huhNXhny2m3KZvbmADYCb48+/UNLYEsywSuXD16
2VWa8c6FvsCsSS0F/qK9AtdErYZD1HgIvnE5UKv9W8h85FtYj/Oa9cMu6X6UA3OX
KU9Zl8bZXJGIzpmPTZBYvAToZmO2OpfwL/AoYObmamtYUsW8EQXzT/M9wwAYj1SQ
/XMjdAi/RqhRNB3FawmjmtHrY8M4fIifoB8HdgU8xabAIlZ8xwCkcmRcg23oYpor
Tf3UnMZCk1nRl01s4yCuJ6auNVprG4WGvnUq7hAoXpZdF+y3xoYadcynA1uqVsYt
zrmfsuiM0YggfYn0YjPa3q4yB4Ar2gDtHUKOU/6SHqsCgPNgTqTgkzzKK2UQXQi/
zGkn+QfRaicglBKd/vqcT7JSLl41aO4JcdXME/kkKS/9Xs1Pq/m9U3pp94L2VOsZ
JlZ6L94orEACOl30ILSP+i+TUGxoJ9Aal0Ah/RMNX68TTTZCCIvQ/43umZJbs6U9
bWt+dAyuAmfyYmITQ4GEmcOGUwkIR+rXqw4+wuWnGUyzIPYPzzYknu3qG0baK1Pi
cis84qoPRSLYmwUsCaFH4LdPAwuiefAuXL2J5oyBQKihxHl5XpHaB23Yp9gYVjQU
lnN3+3/cDb7gVaUQSFLoo3SnQ6rfRGJxrGg8yWSu0JwKcMc6pZe9DHK1Hl1p0eBK
WfUGyeW2BCJ0CgPyP71HodXMdFWCnYCx6aYq5yeSnC9APLJwbQ5v3htBrr1YpkCQ
zV88HsSDdM4pyPc6qWj+SgpVH9k8gtoHbQgEUMWB6s5lVDzmQ/vAN4QvV6wCnil2
0wpk/BNkg1AdPC6b9iEepalmE0PVi0kKsxjaXN8pkp1RuBv8yGgvy/mNUbim7335
dBmYjP+AC4YhC2egOdIspsye7V3oUfbjJLDDa4nvxJ5nRvGqW9ZAg0M1k4ncQbSR
FEewsJqlky3198RtzHLoQRZZRF/KOayW2suBcuDbe1UrY+umRMVcXJ7DoRVsUaQL
1XHqfpR0CqiQ24xCw2TUqEoWOqeIDaQxnixA7hbpKh2v85i+ohXmZWp2KdDGquxB
103qJ033CLYF2ZppL8YUE5EAFztP1k+jCjw5npPeO21FU2aFS5B0W4FACC/0h9xx
KFBepYCSrjEFtmfFFv1geimq8u7cEMsZC19AyShiizSCVGPAtJEezqpDvGJJMVXp
FjYFXMwhSFjWkmYuzeFAbzdrdTr0xkP5xaOrV2fh6RWnwbFHMdCBxnPXQgiZ63bJ
Z7fL9U9clXiWUH/YoNz6FM+JZP6NRTOfvV+aruEo/xdJWh6L5FnZS6vjqHyA+Veo
XFU/4gjm0B1j7BEIBOBbzjxI4Der+Z4/1bfEk7B3aL7hp00NHq8TqGyp7+aw2jcr
+CE8NLfIK8hWo7eCKnAlh0p0pcHS1lKCK/I3+TJlyxukB63JhSFwHEO1qSyXsPCH
Z/SJh6FfaP/XxLLST6ZbLcFnVEvWwTIX2p0tGBE/nyByWTRqId6bvDEkLoNk9yN4
BFKNWgrHDOhovU+IO6w6DHi5dueRS0JNWTI03v5rWhfmoudh1NtuvLBAk5PYpW3Z
eHMKfeVTP+C67dFGlnUGv46EAb9hjsoq/sOtQJQ3vjxmzIkfaxzBGo+XjZ7xDUVV
MHTEttsFNetoVVZU5PWKWgg7KaKLlUdbn1TFSiGjzHJfRew9MQb+nRRwuYvlIVlt
hIaw9mEeavBQbs0aX/xDOxXpFTbuqfqUmmSITyDmuw50DDtyMEf5xYtO/24Iv05r
ucHcBumNY2F0HmpHJpYbjlJ4dGOltGfLiM8fxVbdwF0FVX/+3VyVPaskHqWUSRYN
Lt/5debezpidwajhf/aXlZ4agqkL+pJsbqatWo07iTbb+oKH/w2cpIRpd8lRHpej
mWhxNEzsUK1Zq0XrqnDnYUiiWit1R62MdM0AqD2gU4jAkfO+ARmGSwUXaYpZwDE0
r9TuVnorQWfUtc1XklA2I5Q2qy7x66b/oOHUgOdA7VPdJzc0EIbrxBKraOzVPZxH
ED1u2D5r79ndfcR2VoIog1GGNI+/v5Z55cBj3MzjC6hQFn6TvubXzOTxUqdmmIwm
aQ0W8m0uXfyVnjm5oOO6DLQEIeG7ofjynaQnRKhdqSrVzSm88WCsLpdvQU2MnKrf
aPMu343VrWrlWWcOgkyuBXT6z59IQy+GEOGqSXgu4LPJJ4cO+nQiSrjHAcXbpjn+
3jtHp8wyjryGgUvgMMa5YpgZqfC6YBBNfphYnYiTzFrP6QrI7hTxgwSZex4vvbO/
F7d2J8CZNBz2avK6+zHlRA1Puo28hNAWS4SP7g/APKxdqWhwtK/qOMe0Jah+OSgS
m5auIJEuX2eDwFtQA8ilQa3EEWFH1tGSsjtQB3UWMofy5L16pTG1fBKQyCYib4rB
uFzEaAP9nLy4gfqWRRHaHT/2sjf2Pm0bQZltg3Wkh0YDYaIVRipHDZyQDeUfiZMD
OU4BYhkoI0nd9blFIvmfDDcfFx3VvUSxQDfX0KzfcTK42iYlcLnGxf0F5PQOVhik
St5RZyzqAFFUyWikf2aXcOCHTDq1yEqIibr19gMwr8XrE5r1w1tic1wUhG4G5aRl
HUgUM3MR9+tNWcjA+esHqwyP2Dv4Y8XKuwsEHkAT9DzLrzJgr7eNLY7eMIKu7Xp6
zebY8wT49WirD+EjxGCY+EOoOjDmZkTzeARBUvtmZqJB6Xm4R/rybMxR3zIExpSo
Gze38j9xEM6UcxRkoK9z6aJrDVqvviSZ+CSaP6wknaxEF7ePXSmwk0uHnB4ex5fN
h/xFcDkzIfFWF2MvHN7BQPraHycFx1ERgIIoXtQqw0bpWRuuN9HQwMIuxq35R8im
WegxlIC/ztNtIacewi3SsGiLt5gc9cK7OEseKgNsun8FynJM5PqxPKKAZAyvFcpl
y2FW5TmZHK4TRxMlSdg+ZyStESZOMcv/VqI9VSb2IXHvEjQ06bca55G63U8iSH6M
FB/QINYvexJzu1ufPQgT9glAjKbes5nDeyUBtKZ6wf4eRZ/rsqo3WDoXwFQBF5Se
suMsXVSRcH3JpQHXkPAoUyzhN+rBaf/g1+7ctqhNnCfEIE4Q88SraKccC+QsDADA
wy3/D65RcsiNnJfJdA0+9Crt9E0I5wSQXrdegDCR/tVF0+x7yX++wRD9sUPlLLov
V86VV1DHrSzF/ExJCLIsKIRX9R3IfOFUAb3dwI0TsacTLiQR3PPCdx0YaNMUuU3v
LTyOObBKQvNhY5Hw5TKLhnHcY7ecG+GuWSBJcVckxzFJX4sS1024yLPdppyMF3GU
PSNyG7mrJ7415owxKHULAcHqMYJN3KSYFAOWkpmYuH+lQ4vDX2/z0tlg2w+G2RFg
LA5yyGMKHoBdasKP9ggeKcskiFC9Qpx2uB9wqhw7dS8SG7mjox2X5y66+X8eRKIw
hU9aBH5n6l3j4TQtdxdTLt+9vkU9EfvcYo2gCgpGfKVE+Cu8t9ky3zARvWWZTmIu
9dVH/NjmYys+0H0NDTrtBW9gP/D/NVGtVeEryRlMJnoccVfyujHZ+GHzF1tjZ+hv
BNj/rfh6IIqb79rRG8TUYj0d2M9TmBZjMJ29BnaPIGUCmh9enBpySd8WWZGnLjPs
4O2ikjdTJJcHmu7LMABaalV1mpm5yraeGSCc439ChSa81bz1GD55nsnfJDdxttm8
o60vYHhRf98eq4rFDIOqNUwQxdyEPkc9RZGOCerR1QQMNNw7N/3bv/1W1ZuVrAHS
2Uj5/Mou2xbTm/h/eaSMKt5e78pcPjvoC434F+KMA/ZQaIvnRzj7cXOKYEHKvnyB
jukzleoLrioBMLzDJ1ZAy8CU5zVu60/LA6dwZxSbST988ket6oOevo43FWqkrPXc
wibEi4nTJDcSZHYx3OYIblMg6xBWcRx2x28ZftFZg9+yTIlX8MdAYRlHaOyUWm49
JP689MsNETjOvuPtglPZVdhhDW6O3Tdszw/Q/leGQJ7VeA7Vhn9LwdTsBbgMlXx5
zaIJNsQEwYi1nr0KNFNK+6y0rm5OD2lN3g8Iihgnre0nsYVLFQHEhZ2zhfcMuGuW
jKHjDYN974XSAuetCqhNcHTOrO3i0T2IWM6e9qifpd1Q0lw49iUhbUVXTEtBkmGP
wqEn6o8kKR3GS07cw/uLvrthkV9XwWROQ80tU4WuaaHP/jRT7J2cawMtFYwNsgrG
RfSMS3D3IYtdGhUBhu2/K01CrOiacngrBWimNCvxKWHUGkTvRTNT9UmtkNYw1ejk
ouN/BP8R7X3QK7mpsbI8UKjldsrDQ6jp5y04XurngaZuzKZm5vlsoMm4A1UTTZqF
KMOAbrTYQZzbjDQdUPpdmctQzGfdltyml4jA4D1nHiRBFDUuYqMxGZ0zxoCDVdyS
geXoZecIaQ+9X8nDymdxh59TC8PHIvSJECW9oEuSawKJijXFiCOwcpCVxA4e0Gf+
TMK1g/jWQkv3EFa1yR6MRGGdlXqP17jweCO0iTDegPkzyvdSK2Ae0iCgq2lAwm9t
vpkYFpDF25C5r+Bhc/2zVySfo6JVmLazdFGZsrK4dHxKgpB46qZzyXkqwHOXjhJh
tghUTFLMlN14tGKbQFJaAlm3tlztm+g64KEvawp1Zfzwj+a10vJSG9QaVp9TP3vc
qTB3BHdEVwmNOTMMzedg6tAQhgdCO0Hr/5vBG53hwGoeTH5EUiSEBvOQ2Ghr5r2T
KYfnxhg8ul6u/GH5oVcKB5lUpvZdxMPpKRjviDdfWkl6c4wcIkF0oC+OGD4xJDlA
rO0ArdoTETSyPhmi2aQdGXSshAiFIDs1vVxOjEXxD1ZwNldR5XiaAdoVv4cY6TKX
aY0gK9JdR/6v+2mX+XuHVymhn5XLHPK3ZTRlv4f3q4uby2jR+Kj1Vxcy/c+A1C+j
3NefGviuT8V09CqbZYrzQnSkOWnDVAxqXL9MDgPQcWb0gd8/Kk4kScMKIJN9gwlO
X3KiGvT3guQWF9aO0OSffzrPyqMBdaWhN2wd5smkvOw5+wPzLtDWjJvGqRyzLsnf
JjNwBLNr4oWB/0+Tr32CWJCkSXHT3LxZBKA7C04SjXj8AhteZpEKPh+3ZmV8Tu4X
vbo7HHi206vwQplQ0NpXo9cAIbgXFiQ6zXeJQZSNChgbEUduafkOIwOAHgvojOZr
UfciuyunXjUyadSIfTWAjIklzpv9d90QDhiw8RemAzVUlvePiqlu3+fHsSnjhyel
TKjYGBrsfA7P9o2rCvFYF1BmNl+suLdRoUsFOXp7kBHvinocM93iNfuhcr+VjDmj
EUCATk+zKUaXZYGVnpOt4OV8/oRkfoQQaOn9lmqMwhUwefzuV9CPSftpW7bET0zE
Tk669IJzSFFIaqzMuZ6BI+Mzk3NG4W9/6RjDb7MB4EzEzRytV0C0DSvR/BwlUPae
I9RM5NN09AfGL5SoNAMI7ZOgpsQcHMRGbfCwZg93bVfpmZas4tMhT9etV2PKX33c
BJzRiE479o1E+O6luDY+wPs73MacSqIpzOYSFOzo26zwsBqHQ8QfHbgFv1iM6fty
IW6kwwMbWhTQD0sKt/QrpOIeSW6FDJAdPUs6Y5hSeeRAoE9cQD2mtBswrSLZ+Jwy
JeH7i0SssntcIlYNs2YvYfPY8uiX1MegwD2P68aasEdx8EkFkQkzoV+j+b+CcuUV
QlmHOt/oW0+cwpSjkr+hIieVImxd+iYDwPA2pFOMUP5YfF8Nk1asXVHjMpQoSul7
K/UEzo6O6b3YD59yKBtEIeyjMJO8YVeyC7Sp+nZPLLjQmSM0dPD4/o7U/ewcywDi
Y33/LQ1+DcfSdk3k3rXY7kZXrg/tQOyOFbG9FMw7fd7C9paVoeBBiVJgkyFta3II
L298KO96MtserLPem+XvJHbAHoC7cJVs7zc4PxI3oLgOqSLNbCsU33rvPra0cgvS
jagBuqo+ExTeMFHXW/4Kl6BQGWs0fAct9c1ISqLmOanPNj+eelNDXiEPqwts75fU
jYY2FJ05JH/XMTN0kR6+IPoYrgQW5wt1v7XBTKDbevrSSKLqHerl43HfmM5lHOVH
P9fZSl0Ezq7I2GflCFzEEnnU2t0fLHJC1HLw7r+qtqatZfIvArUn7GZo++IPlfw1
Bk/1H1K6Hvdo9qAJPVp+UbtKrBdDa3FlHMMYGKeVRRsuyg2bIXkwz/UuvUbvfsaW
wk56g+Xd8/9XELzv9PGT6uzjpMwphdCYOAExxzw/mhp5gQS4lkch6rTuzbNZC44I
7utFu5Jg7krrKdJA4wVeIGInh+Eb9E0omQPdVM/XSHzZJwJPnqIgkmo9+xzLy7Ga
0j5+hhi+6EGBm9H/Yshtfcnk9bWZBvvZKYVvI77wG+CnCxoQGgTVwW3jDoMNeFQk
LoGxMgPN+4uFPX8q+CVWgDqEDQUHmbwaVE4eNbkKi9BL44LRcpOkVfLoGP8ypmTG
RIR2ez8kU16OcWFw/oYvE79pl4xg6kcjURzLjZMsy2tqORoKvQ6akCmXLXuv4sfI
ymcF7HpuqRB1eo+7lC60IEA9dlOVF8QFSX9I+5FNzvwXKIXFCRZBUrzACNjDPeWY
MLWHOUXe2aqyrVSsVJmKEmDGjYI32llV/Cv5X2H+tGtVcWUiVXnMvHFXPM0ibLdy
rcVnA0Ln/U69nhv/SDrU6HVeMvyRq0KzjWG48wchNo2PCrm450iv1S8gxuMODmSz
ZhF8ssNLJ8qiyigD1ZwjY+iRq03NVzoJZXv0uOeSecpFKj5se3t9YW+5TNRbJ0b4
wQ3r4MiIQyFM1GM/0KGwrBKF86WfkURXGx50SwUB9C7k0lMXUU89b4EfaWedKaX0
xCp2zMaj17agDcrcLF0/A4+yLL7UeKS5fZI+S+7uHDeXs6tCLH5XsBQJD3Xq5pxQ
afGUEXc1DoW4/SZXL9NgdGP4kevrmnS7YDGc+Y7UvKs+TgiETPUTvbBHQQYLDJkF
3TtyWHnfbzJiRhlqlgswOfWldqpTXHwBdfW1OLjmyG2uFlV3VHctogHRlWCPVEjk
iTKyT8xlVFmf1ose1W8h/sLw9C2NxnuG1NqxgEADUWqyQFP+HhyS3xyiuiadSuFS
ckgi5zdW6VqX3gwQLEUaHH0QZegGW6a8+nTelcZSEhpifrz7ZhfruT2Qx3/WkiJJ
N0qILbB/hunZGWdIimhrFnohRZyNOAWIeNOv45SoG8cGBKIMjsUOPvIRjF/0kNFh
+KBpJe2GhmTGi0Geo3yFdOOYfnu+9UvsQXqMMhj4LX+xVlZsU9l/5B9dmyqF5wAK
4ET9iFum1Bmi1YQZgVHAlM48GCus91KlzW0JtqxEpVd53dOs+s0LRr7D3qly9SW/
+yn+CHdXMWgjXm8+stUUJQTVPuu92SxPjAg6zglXtvuT7RZVWx8peU7belBGYNZ/
cAzsaqDBiUlZRPTHD37oyaY6TxeDWRwcVbiohZgwcPh3/QtZEC8kRPQBIRXpqGvz
xm0xUMIkXDljietL82raGoxgTFF/SgZytvyrPQJcD86vYaA5Lc68eHgkxHnnuMg4
mmLILKjamkmLQsGRzsmmR8Xoy/1x1p4qNdS8RKc95R5B6tbmzdN1LZ6FRXz8ZA7o
7/APWmbWiShUAUnmOU66M7YOidk1QXsZ5++0ihS99nnvraYYmVuO1HFApWoZmoTq
X59YfoDQt1xnzrattBKILKQUDfJbJGhPaimLnGQN87juWPEPN2fCbj6g2MgXSSz7
MlVy/95PM3jp+BBXvI6HNVB2/4fhrcG9LRcYCd+XHmeXy4u0o5XqLZY/ffhhpNpd
Jmzj1TpljMduHbaTqozQ6vmZvlT6HeZ4WkpOf8kKsIISOaAFAh72FUAi719oG4OP
3/aJaCK4jqGjYjLQbdZnlwDQast6voomuT4s+01849MCvKQz9kGV+YBpOoypmd3/
WDzeNESD8IjxsAZxbvs/G/DHiI7mJa4uIUeVOcCj/anvzsv+HPLWt46yFUoL2sVv
OFZx0sivWZI0NW+BHna46u9GpGPW2Vt7xoLX4yjJ/sTYFeLi9PdWpkD5ie73rGFC
YsiMaTBbfh/qMFzWBbD59BlKUYJfdbUflvuwudtM2Kwws+QSyv/uStov0IBrY/Xr
CCWiFOxqj/7fnu13CGG1VuO0UL5mIe13XGpwFaYxhN3CVeLL13WaFe7cGzmRpOFq
X7sDTO5M/ZDUXZgZwkUZ9HHxCCSiGqLEAS89fko17WTsvpOkdl8erxJU3VwtQXpb
rIE3TYTNHtgPNjb0LDF9h60sUDAmxDTb35N8SurlTA5fsC4gBDJbP6cnNLMQTaqj
8emlbeZNPIKaVcCpbkbkEvP7/Hxu7IxDZwU1GvXLAV1avDuxsGNi252Cvyxz5eqa
ZL2NviCoJIDhrk1+3Z9n5Nk/UhnGHMbfvYl78dnip5rR6XITKIU+9eWtGuTigf/1
4lCqbGr5ZWxUQ/lj13hEJ4vRlIpUH6W1LMxti3JU4VhiMvn4wXO4NF9O1KTssDgd
jQrZ/DXJiDJreJQQGxl0HdDAGJuQVlkdtCLnuyowAHvWscvO8MRkv7NqC7ZOAUGG
uiPmK46JxpGwDe49w817oKltIsA67oJDQzksIZlBTtshnpdvdrcD8b151KD1xLVy
WiLMko7WsIsoyakUwiNZk/LrzDryC3I8IWahgXapxXM5MIchO5kpf+TwOstncSK8
5YhVK/BbDNBvrzI9Tk0YDwNNZ/zPc4pc8NZYiwUoSwBHXIBltlYjTVx0RoHT42Ep
CW1gqEkO6/mGXeT2h0g73zkcpYvPwwvWUj5DLi6j42ej2Fb4qU4Wu2wC3Xn8PZ0X
SE1/SOh3VwIS9spNswxEXTlSDfPyyrV5SxWXd2pOZPBN0vtzTf1bP4LEBoloDki5
FXMc1mMoucZBaPrezsg/eU+rRlDkZSpKndVW+OYJ9MuyG/e9goe3dpFhofPGZiW0
a3UAs5xXco/aPF4Acxq9qnH30zD+plSnoaukP0hF45P7SEGhEkuZcR+sqlqeAIom
IzPqquZZMSq45oZopKnc6TNhlhD2P5mpYFG09OFlUNG3ZLwOEauV4TBHMNN02S1p
aguWCmb06/tHjA0OFuCyxvOCniZmRMOPOWlzhN2gMFqNEz7qF5TQDAV3NP/hv+MB
K/VyMWBpEdB1Te5Rmjkdlqg5D3Qt7SXpd3B5JKvxQS36OLvjFgJmgCudz0ERLSRl
mlO4h/vvW4yNGTefsqxjqvJOMeBw1zTMaWmwnUrhpIm5ufK4n4/jsk1ZAoyFQsO2
xFSRV7Z56pcFaJV5jCaQVN5Yh/4Ugomdd81d00HjqnX0cYHlvsrPlTL0l5fsg26X
7eDNgNOoQpga1xK8lvE+iuOWCp1iXZAHwaonLDcXPgKlqRc/sbWJrMcjd9tgL+pt
oOzgVOiF3Uercm2rPTvXuxNLj3jAmklgu9BFIXcWR0tAPlr9lsesJIDKhcJIkLyM
adTbMRh0XD9iMtqq9Fbdz3di89WGmQSA9qb/ecBS64LzSvnK4RHCWThmuUTDofUJ
FbpAcYzqVM7kq2VgDpnCMhhzcRknHor7xqfA7Lj4P0f7RZrsRQu0Uzl+5dynM8bS
9WUbiSPl+o30/AyHvOVeBn01NOFkqpmovg2nWbv76yhvAK9NbBwry0CoaXphWrAj
nNXE1WhruRXtje2yopIGjCLnD4gIwX4FyAg9vWqOt6msZQSBcHDkTiWe4Qj0qgfg
Nz6xinW4yyk1S2k6wa9iY0swLWu1aswAFwA+JbfmOl8KN60RHzofAwfCYGJv+9Wc
GG2CjL3yS47TFajodZuzL9cyP6hYZ1uCmvn2hg7Xfq1uL96GcruXnVTaN2g7HtBG
9UCAaiQTLFaHfsVIcWafNLv5gAt0P2qQLFf8vUvStpdoC24+9Lm2Lqyg9pwyEnY5
uTN8tCUoMkWdnUuEIBkuR907yqJ08e7d/Ezm5fVLzw6l2DKq4Kzmu9scbr3B9yVd
EKZ58mYTyLGLR4GagwYWKDVeWLuFrhhbPYC/FFg+AMSmp5xzoYZptSHYN7Lz47Wk
iv4gsh8QntUVQQih+g1rkQP14ccAqZZ3fjWMWp+HwFMko77SIO4WjUunDytsW7Z0
jghUyn3Pq/bt8316qNl6svcCpVitD4MgRJj1nwgswZct/wgJi5fIMvWFMSBHKvtH
2CXJjs9r7Sv0R7uowJAxHhxcDDgNI6o37Tl8HHijSda3V8Sbup9c2qskuy8Hq2p4
GD7brJ0n6NcMrJ9rYWdr0dNwl3rqIhVt4xWZ9aTtPPzoHusO4t5Gxumzk5JAV2UI
BP8fsgVolSzrqnyMfw92VD3v54Dyh3NpQWJKLaTwEGkoCdh7mq+r/8qw6jZ6fjeX
PPPvJxhjJPtEeDUsgae+Rbpsg0Kv6cxLrZ8N3vwrUfVNLKyjlyOKw5+blJsZxLjC
6rAtGAeXKGUwLGLCRTuuvVV2bJG9uffQ3WwjCY25yQ8tZid9eUkH6t/zbsrT3tyt
U1B75l+tUbuRU0quLVByflqcENDJdec0Y78rcpLKC0BYFzovBOSroDO17micFVdn
vLh5N6Pd03POqya8U6ISVzVnYUyRyE4MvdcXGEXmAaWr4nUqgBJkirigaH5cak3p
u+P5dhUd0n9aAx15eY8qCUp3IXzmWmdWTIOtHhVicBZfQxxZZCKLgAsxj9Hd/F0b
qUcz42x/VABoHjyV43ZyAqxqQaHZ6GudbLxhjgndDciZlJABvaT8F4n/5wO5SMOn
hRQiSwa6YvumunBl8Rvoc8B8jp++TMcX65bHfeB+8US7x7tR20ao9DHWZBvMfmzc
qAV77MuQRiOXGr0HE+mq1/rvniMmHDtCCfUvemlesae3xxqrgtOYMjw5TUnzYBAU
vSP+2Q6WBGPcox5P5Gpdt4nIePgYMp8jIE9oqgToc72cyLbFJKXiz+mAnooJzV8s
wuutL08fy9I97y6ZqhR9S0tKNl3HxfqZfg+oODpnuNMDxof/fMluSfzInmTt9Srw
Z9lcyzUx3OnmCE0K7iuDfbqavlr2SSHXbIH6aU5v1T5DoUNV9QnIpsXvD6ghgpmQ
LSrlOeIvfnh3WYshBrCzc5Gwrc0zpLidn56RrYux8pXzeG7Zpd7jiZmGxjU0Rjpx
pqcZg/Y2QtUYsh1siVdw6R0pRU0lE+sCntEAnymg5ZJU5PHMqGBJwid69KSnXk5e
gELlyRc5LiEs/H2VsakiveIwFLV7lT0BlVKHmWqkcq+Fu3v3hhvK6bVSHY/15sHh
Y0i9DWGQ2Xq4T6SeQPGVQFb0zGbntSh3DlTXDOH4YVSIgvSkQrrBrkihWLaTDeyo
WYKF3Az1WbXtAQf72ZxOUoImriXsBfEzJ91eUV4BTa5pqCJrH/05Lg4Zd5Opvf8v
VYTadfxpwPQ73LRJDOvH6X0Je+0rVBAGTdVKCIWv2a5wV/p5jjJ9H7fAhPxPlD3P
9n+9NukbrDRdutTDPMY90SKpe0LmaxB6AYW6ebSBQBzbK0WLrVzqNu8vWVUkrhtz
Hl7Z1jh3VfPPvK84xnLcoqkP58N0l42xq06zOHEjCKpkJsZpWzSXdGuCvUhmt4it
rqz2CSKr19ysDDSt3FjlsODpjSRI2XU1pIObh5XWNyAC/0cClQ7311KS20f2b6pT
ejsxMWO4ejKCeIpJQsDu+cp3NV0g4XhRZ1Uq7qvUyt5kczjQ0B0xWX+YzoiXLMdg
LJ6u820McL7lfsy+6ZYs2kLfmQYgW9l3+3o3MqFv024SsoowWqjbCrwnmbjl7+P1
1r2Vk0m6+R0o4LYueem9Rg1q8XZBZ77BDdwNljUZNH0P24wpcjZlmihA2wLRcD6m
2JOormw7MPrC4bSe8F5iCKipNSF+FL7eSNhRFB60YwnhrELoTn7Y7+A2CoTxfvgO
Fq8QyMV98USGouqhJMqwkcQdtxOdkyrgRqNd7ZbMAbzx6F7j9wn15p9WdHYdbf19
0pyukhb5c5DMGt3LesON1UYGjT25wb+/eOI3Wcl5TklegWSNVCqzWnL/eo1Y6TzR
LSl+IT2m6aeyDbEY3ZKHDq5zWwX3DRXNFUj4wcL8KyTd1cH2H5yI2KkGfZd/J8n0
1EDk6u+UUAqucOXNmDXbYoRIEiGTp/yd/tRrwaqgTC9vBXC3hrRCmgNCfOe4NZ+C
ZdJHpBD/jP/t/74vV85TTmVwSMoc7tLYDux5SA3HyyK6RVTNyzB7XCQ3W299xaaJ
K+mJb9h3aHvm5hS/wR54tJ7Phywh6rDAIKfZzqHDICkgjtheKjY+4PcIdLt000Yi
Ph2nilT+mr4yGFizeW3PurlKhZXocO7nJNnJ3d4EwFs9LRjYc1YUEeCOBIwF69uH
iCgWQcpqtq1rDv/chDH3URz0wfT0eKzX+r5zE8kVh84EMV0ik1sIZ7VaEInlnGQM
jGBm75MHlgnf21g4mjafCn5Meiv+WMIjwBdyIgX+YHXyOeHyhIgWmzojKxH0Xgf+
X9fDSftwbFZAAMyOrUW8jpvXPCvawnSHwZIUBoJPPyUnsu4BZ60tYvRPMdhwyTnj
EbLclwly07S5RZiT0PWTmAA5aOpxqVh8gt3mH3dIOtiwRsn8t5qVaeMAxYvnSDoh
YrFxkB0/4E1ZLZeV/DAWA6ZrB+FpmU7JwwDYRNLPTR5R8tRjgEH4avOrPJay0MxI
hi9ltlsBShZ7GVGn0ZrCdOsLiVhVShWvCO4Q7uUwbW/1kOXKuNUUmfsEJ+g/moUI
4/o9jGz2dcN+YaYnkLlJcGrLZYihUT23LSgz3AETIZZnO7rNaBxgvBJLTHvtlc5e
Wv363B0m50nG9ivo04WU+eAULe4bWAXbbQ/eQF+XW92cu559e2+q88V3kOIK4UqI
2u2lx+PHPsdPjpyakG+hljlyI0b01oxZG5jMXPta3hJ3Y9KLPiZ5MwCyF0sjoHx0
z5lhdjnVrP29ee1JoLQOdPIAAeNxhJDcnu3Rn3PGAdmrVu7WjU5rAnG4L1NwULBM
kPAGmjzn43Tfy0X34EmsjznIikWCgQk821xAXiqF7nJ5HBt7j7IBMzpBmRgHuS11
97rvZdYqgZV2/nwMPrjkOmyigo0dB6OwTFXi89APJw8pSiG91T4LBTl7hZbYpWPz
20+fe/fB7MGYm0vgc75SHuIMIZse3YZ5ifCaGEo58VOkJeyInNzdtn6NPM6C9W9n
IOeZN/g+eTjWe1s3odc2GhSCaop38ub3w7cH8W820EVs1bT2b69DH9H7GNs7VgeM
fPZMLKiz2pNoHF+8z+7XGnlsHilBJ8UoTg7W/zC5baqmtnlU5LeqtshUG1hvXezd
qyQQn0q4hFnc8i4MDHu81KdPGeMwYNfq0XJN/dIkEguyp6chtWDxgOB9PQ5v/SSf
zrz06JStQu2XjRB0UfYgKXXxQk9DZPRnLEoMCegI2vwAV55kD2jTnqFzH5O3DYhP
JMLKXBbOVQAj2sjMahUpYcMAhPBf2l2Rv+gtb5qjnkD5gsMPuWwjmSyQJ9Q+P79i
MFeR87PuuZ3b5cSuDqLMpzvTWR7hXcdr2LxR6GITW4ir0KpPW5KsPzfyphhiqt7X
A2U4l9SFlBi8kOdBmedsunsLe+R8tewxIX9Q24LVFkoitqZAJeBdJ49AXrj16Jw2
7xQiw+hujevfI4H/81v9SBg9Wk6i5ORIwM5A/vWrkNKJy8M1Ft5JtZpIfY7rePxm
fJMCBeqjVSKAB5Gud1tzXcAoDU7rNFy0scll83GIq56Dp0+9+AIDBe36810YQ8ES
sXQ3+AXAP4eAnkN1TCKWt003mN/M7lerXn71i3HTZTbWwHumAxSMP8XsAHWApwuI
suxVIASXAn5q0EIYQRvUSnkUZp1NzhcDyIagfQzLDiuOPe5VnYx3mJv0/q5HIOqv
Z7Tp2el7WMQCMz+WhzjgwcX4IjLiRyTrz5GvTEL7FV62tpMRi5Skwtz4KgNszFLo
M5yI7kYqu2evILnEyw7sJkyg+nqs3+NoY/ewYev2Q2zb+7zcEB8qWi4b8FdhYV11
rxMahOhKPeE1+8JLnygbqS/Wx3aQqdMyPLJqtTTBBGv4BN2HFNVorNDaGKaNt/v6
uQK7JL89wxslfFSscE3LCe215xRyzLvTmemNP8vODdxxgEerYmdweMv0wPbq0llw
FvVGdC7ZNTxdM1lsMPssLj62FGnDHEtbBu55gbaqIE5TBpPxTn+YGpktEiHH+DAl
6MHyAFYM6BYHKNgParJkZcqK8jO3MTp44qRbgnBBgsR8i8babivV3zz6YAMfgp48
H5WfvJbkCu/2JiNpuskvPen/+afrCdHkdbQdFIiSQ8OisbHjYsKHE5xXlrLx086a
/6U/ShPRRmJy9fTrTqyyjAQ270tdbYNpUcEyX633SXZJvkRQvNZ9nwKocEXPdgS/
NVmUnaDJuAzCgDAGMGeB7rgi0f660ykWBG8ZSdR0K/r9xewH6o3UZN3UPWcbng/H
9fWSWvdLplv//HcrrYULsgkFpajdZWT7MltnAGyz6HZRe6Zg9zBIqKqgEnvloL0y
wEDzxaUZAbv9Ns5AcYpuJpfRhH+OInOnv+d4wInBlxdod4R5mQs+q2dn34J41RCa
eAend+PLHBliZw1naH3k3yfSHVBarwoTVMvx/0V4DWCaFCbUL+Tl+w/O+Av/XD01
rDJgi1I3/WfSBemcDJZ77qFljfz36NBCHPJtWh6TvGGr67avqXVSNBPwpsb3gMhD
FGrP/JX7tUnsKvLGTYiIS01D9PKHOcMyjtAucONnIL9viz3XUFSpG126cpsLjGLp
nwDKJLDn7wJJpzFBLsyc/P+rBd/qSVG2Vw9IkWGQJ4DkRueQX2LzGc4JYz9aLi1o
GStYN0kYJXp3okRWWEXgDJ7gBA2t+aMuEQshpa49XBYfaKusmLHYTPLYJpfbUQ34
Lu8gIYVwqYUp6XFrGITQZtt02F9j3sXflywyZHRmEPMdpp1cox1GEkPttptUxlN+
hZNxbnDvXrQvH+RUiEDlnm6+hl1NiteVqhAEhNStOJ2nNYa8ck87QE3g3dtzU5qd
Fk+Uol+PoIwreAXp/ijO2rHwGdD6/D2qxdJrKgH3dJX6md8uwFs66bfnfEusX90Z
FJH8zovwZuRroLPaqVvP7V6Ek1xv5TUOxMNcP21WqPdMLDaObk3vgQ9tQ3kt/gss
N5FSIRjjYDMaoRzftAfwQzRzWGmL2uDBKo/GJqgcyQY9V62gv5BE2+rlVh8zJ7jv
FgsuWBhgeHmUryxcuY8g9DVzJjaO0aDNBh2qz7Ljv/WF6njV75LxLRcHmVq4QiQW
YgyRcIiPfTmk3c3bL57H2yI4UJDhYnMbtogyW3TqzM/b4mm9GQj3xg/wnP+zFsiZ
GpUnQuqUqguuAKPufcBJ+jncdU5SQPaj2Sq3Fn88u7sznFbJpL4i/fEyh1VSEVPC
9h0PrQr3cya+lKteq4Z7S22VsHyYqht/56Yx7YaN5tr7XX/AURHFLZP0WIEQ/gFQ
UHKi//uVlBHNg/X4O5bbUv1I8C3QDDBEf985cYSWeGjlDrcE3JHvOnwqaodXLj/x
sRb8HtZwH4x/JBOPmk01cMrA1p0sSGKR9Xh27pDbwZilUlSOgTcOtfJeTS7IjVvX
TBFur9KX8XwGtQLiy3GdgSo3UJ0qD9FGomQ9Zi/64Pld9/YgxefpTpnjsFHoEpvM
wPKDocPB5m6wmUcc2hv1Ma+TH+YmevALTFKw75KvDadHcwhYyHFehGTol+wUXjDj
zhwReidtHvvCwSu/zj5RFbj+UQ+pNl/fdSBuQhbKp+bDMcz6UkeMFpMI4LXrD3op
/JeidyaZyc+2og2SQqdQj2xdCOJGL/LzKFs69NqQP8FT/2uQ2T/jkMZ6GtENrNu9
NtcuzyiKSqMJ4DWrKi0FBlC1b3jkkLvVRyGHxMDldmwDwZL+hZaXm6CnZ2ovHHFX
nAQfCIwhHlGX+IKgjdAvMnxJQC7PVlQP9Sf6RT/emEJcgMGAXspnPb+FcHwlCO1o
rtCp1etXZsD59GpvhIbn7OZqzemBeE3612Ynod9ok3n/J9CtyBUfe+tTyD0YYnBT
7JDOeC+d7x5plaOo4H1cCRxUzbyB6lMmieJYDvAo+xzdlhpr1FpGmUrK18tAaQ3i
aD0hausoaJ2lEKWF1l0XcVdzABVXKpRpwPxilZhl8OR+DZ7mHmZo7wAZiPqOz6YG
dI/6VBhInYhr5WDBpczbkdwVEX5Q1pdNlISviYV0FQC9eHMR3HcZ8I4XtXyqe9F5
mMv3QcvATBNA4cQiADJ570v81n/8TTymAxma6u7h444yxgoHbNR+p4fOTO3jSGSI
xtcpwF6WP/POAVBAiLqQg8O4t/S/Cr5VWSLO+YkavkB8PTvN4nqbG10vn68U9rPK
BtqslZr6AgP8g+0kEcHvcf2JS1kYoN3gs6QEgl63Z4W9KC6iVLxXc7XgXp9wAkxX
bIs0pdcmU0EvG07ZLHlg+g8wEQ0CtAq5Nf14QJwXvg6f/kAPebZorahwh7cHZOLx
WPZd8sv3PnHWpQVLIpNbr5HY4LvzVDxUWwC3D/qG0Z5OX6NMWtrWJYkynxvl4Oir
azp68jeUfk/Pgn3dSKgMuztCX2KSiF09L3Li3uaRgJWCVAvwk+6FKtWwojtk0bHy
aNcA+q5CYXA9Ul7DW3kXIA/vdHH+eOTpOGNGk3Q2IlY4UeJIi7Cz/550VCoDtbjg
5jz7p9qy5TTtofhq7NnLxEWfLX/H8wZmiEP5sdxsVu3o8WiuyRyD5jfbtBv1Ey6L
eXa+iWI9tWiDNbIE9/CsFezO9ltKcGJx/20Lq1AGWH/Ghaz72NeVLQtUOn73c+Zx
IYkmbtYb1lZ92QrNWyb+IdTLiGoU8OAUwTimy+elIAc+mxi3VD6AX+KCfqm/aYPj
NymsYUeSsvfsISakBK6fsH2+KZ3ol96uoM9qhzr2yscklsKmoiQER9LNkGqCWU5w
6nhJ4aZ2VuHeUoiEYRQ63KHNtaelO7Sug3eun0zycwAT+Z2AbZ7FRQUpATGuFinU
hWS6oxxXIPDkbUKArDMJx4r/d+9QZu14FmiE/krEZiyCVkjoAHz0sbnX05WsTmia
he18D/9HARXNDevcHxik53TOSjk4IiM13lNug4wPMySuENkZnWHi4ZM+Ioh1c9wu
1399OSNqIhy7wsrYT0UnL26QcMMefBgMif8bpWzeqX3yDk3omLhogfmzppi8+N4N
m8kJHuQjnL8YmEho6EVwq6Dcbl9dlZ8hjQKbhdwCBpnjP4SLg0GLr9fePkQ8iwoC
rsusKFdXKwky9CRt2NZVKWerUo+OxzMiOpvUnefclFj2gMcG+QwnFEEams12XtwF
g9WybUhwi85/XRfyzrND58tKGHwCgqNTTFttK0jXN3PdS5lxgAP+Dnt4So1dYPK2
v0HUJf+L5jP27BNVvJqCvT9BD3j5OBOoaf6xzaq6aotcUckcWQXWhuxFtZ1gTSrp
hGaQxnH1+iEUG9L1iKEyzKlKtFVjATD7WPCmg0sWZ5rIoHNdWb1OSzP4blWQcnp2
c2BcdZK7B7WJckQk2gszpGZjLPjsImrYlvMVBbdbYwMU8youQrCQI3FHzbESh2/o
REeyuwzT9PuoSRUN3N9YX/zLf+dTbs1972ScL1tUlwdxziNVAQy+1UvYyUwC5A/D
7w28+Zy3OUeuJkVLU9uv0hT4702hbkS03Caj79twpA+cmZO7pMo08I14+C6EeeND
8iHKt7Md24NGY8Vz4WkNghH1fLldmZ7yW2L5bN9by6C3PcPw13Swb+5PEwt4hbLS
4WfJti6bWuNc6/qFuX8a1JJAusSSXEEZf0OsHPV/YRkKe0Szfwntw77kGDSk25AU
omEhjSJVIQz4cP+tFQRlQ2giJZiiys8U9cKwTGfRmYPwqkrIexIhl4ETKlfooiWr
AEe9vqI9Gfq6n0Jw/U03SwZgnRD3EMza+oRPlGj1QBKp2ikdiguA0ljqpLtZEiDD
W6g2DcTR76xu6a6QNlA4aH1u8SmxAtdnLdyxHw+QyCqXYA6sHra6JieI59f0rUlR
DNm8KktbNW7XFCoJWA3sL6jvHAjMGu+0Ls4gNJioxGRQaUuyppjMGkP/l2OLr9df
5uyrERW9sDUYJ/uJAgUsrTjO5b2nHYascPVvNP2adhKN76K9pVQ9WKCT2tlCyHoS
wZHHOTqF22B/C1TIpe4eTaNiD88hdFfsI4m3NrrYy1LwUFbQEA60UsZpZB9E2x9+
gjuqzNxY0HIzDRiPl1jDzqKRLNK1XPN6dsSlEWPHQl1fNncgAW44Of6fzg5VZwJa
kAcvGrShT7ryBpr67/qIj3UN93rxbilfCQPh+Jr4bvEEKrfYQ7UffO7uFuSbwtA0
Xr+V6+5tdcDt2FvCKqklkXei1yZ9fpBt1uB+/DhibG5U/ibKzdEA4l8vQhqkJbuk
Jhv+FnrXsardkZuEkiZwrPf9LXKFe6JI1Gy3CT40gK9DyWyNJoqO/RvUU+4x6XBu
fnjvUwAeGzG7aqjzfleVamb2HImffZqEmE0BT8w00wEZRsm4jXAboQqQilD2frwe
/tdOtdrhd1UTqACYcKJuAo68oYQ8xpKqrhgJEVDDvtyalOpgM2ELU9H2f1fft0q2
L3i4M/KUD6Y63253phnPCErhzem+5Ihwjq6WWVFY5AmkkN/KZ2PIDv2Vi1oSRY9F
8SarOFbwAVVkISbBGxNXzRi69QIT0iDmJzb0zZZzfBVgoUd4q5ifGrFULTWcsFlE
oatXAmdRgxp2LuPXba0Ep+ua/V1kRnhmnqHDTEUc5hdga2TPQZvuT0uer3oE+/Kq
PwFeMIxdfuhmXVwszVRbGyI8nyh01BWcXHNFqdQfbRF9i9OKTem6Q3eYt5VPPAlx
2MXUyImGvhPYLN7yqsyIl8DSXkruRGgxknPkDuwqfQnmbgh6Odjvzlw4icoPVJ5K
gO41qFfOhFwxN1sDR8v1goAkXYRRnO/DYAnBw72ycibmt4e8Y5nXE2UKffhN1EYU
HPn18LmRLUvigOfr/2A7zJUzIE1ZqhK1QtMs2mfxkyX+FI2QHpz1UZUvDAX8IGxJ
Df/07gdkOOLYbVdwMWfMQgqE5WBBAjhSfu7ducsysZURxzNwn/pgniuXjPQ9KSPE
o223jQsO+vYwm3fbtg7ZkLAe1/zwoIyULT+by1wtx+EQ00A943qwM7l4XLvCvpaE
5Ye4kfkm/KTk1dQjeiypBIY5mMfjpwIEXm05KtXjdRIfkE2mll0Tag/AbK6DmcUs
LMGGdozLv2hmKF32vc5MSXjPDR3/smBUvQFvRi1hgN5Np9Cl1iNoYvGjAoWobptp
kYpaJJq6j/VxQXwCmCeeyaPDuOAp/kVhyXtLU2KTC/5zJnvVN2aqBdAstCwNI7mp
SDH715z3VXEwabfhNuxE3Zqbn2kUeDUEID97rbedoKCzgxlGxleHJcjQfnXIziGj
pHs1bmMZgp4MX8Xa2TJS9J2Uw27cS9aGmY7Q045FJyajhnvzPNhd4f73+blLqlUS
mBp46PrM8AVYlEfiy+DZ84oc0aTqg7hZb7I1vOvbRJp5wbsxVAb4fUQuI2E9NqJ6
zJFTk5nxLwtCZgVwJzbKf0fBQ0rFkwdHADRVT16KKxgX4CqH2yv6BugnHFbT98ir
TkX73R29AWyaQUaRbY39Pmx/crqxYwoDjyvqMEKZZaA8esijfTwxynxDMu7v+yJk
9Una/ssEn2ImDCKj/++U2CLscfd5RGiCgbhI0hHCbvUvmX1sqOKs3pJhvl6s0Cm9
dc616WKqrc4QYwduWqDF7F+P/4VuFB9lwhfVYfSdu7lHQ2P01GIvUXXFpBQH7lPz
nziBnWB2eaaSYA13RVkEV/7x4jx88NBAXUfFUVXVxXIm3IUuajA+xZGm+sAGyqms
oKV89CfXaXue4mzP1jcm4ws8y9RqVZHoJvkMnkclgiCRJ9peqC9caffnSRnvs9gl
YNAfufH6U0p79ufwa95ewTUkdJJowbSQSxThSVjR4q8+jsoHqdXJpH5UnKIyHcB4
zqPt54tzR/Bwd88wF2OKjlLewz7fIniIqw9m0fRQQHPhbfOJ9l+GuNzo3V2yk4bW
i7ter7oVPudnwCsND5p2KHXDKoK0JbvzS4lfseHV7fHKAbJ7+xv+nAKRtLQwc79v
UtQ8k8Xg3ReBYEKccC/uhzfMareN+2hBcc6b+sZ3r7nirAkk7ONSDRm4KqxJ7O/y
pFEeUkAKIx1ULmUKkRslTgt9MTABVnFcIE+u2Sda6CDrflWwvXBIDvi6xvFvMi7I
V9oBRQnOgKDeeLNCZokvh9LnDFp5FLLohrbnV0IPrQzl9OjzwNodjuNShJfl7s+I
hJdWmVM9qNb/uzVWYhgBdiz25fmqgSgsI6HW4znyHJOtwnXZHITOyg0J7TQ3K3FW
fCLiNLvwT9jQIkLTiqM+ZN8ULQ3rSO295qOa8MedCnpRRIaTkO00ziuMs/yb14/S
cYQBYrMT4DCIwlofdbG1p4a8KNAOoIokALtIFkijltM3Eefu2HRRyY+oG7ygyUCe
uD4x3oQM3vb9zyoN+e8Kvt6TcNH9b3YYdewsyWNkc3Rr1lqUFBV4GM1eEqVM/6Ee
NRWaTEyyby6ilfgjkwvZBWClr0n6dUAP50xODIpDIffMsS4ZAAkqZuSpeTswW1X+
SLWL+KVcC3XCeEoslHTKYaYZnAfnTYf2iQCS/E99+UHn4EOOsi8cddW2tF/PuBiN
SqtTzXkycr6Pn3QDnoN3jNfvFwVAKzpM6XZn8/VGoZnxIRDb4iCemBMQR3dBYBQt
jt18eAuj8Xj3HNXnNCwoofapaEeDR/7yA7lYA7FrwZ4PC28xGFLYu59ALa//smUt
6jzZvnNLBvweNrMiZzV5RSzqXf9uMlcpV4dSl+jYhb58ZwN7TYBA2bc/w5YzBcJv
DBC/1aduhuO9awIPe/lcG4TZx9uExq1k5F6iQP4czEo1g8Tfh3Emr5vEdCA+i7ty
2RY9XWuERrDV3SBH/px/teYd7CwwUYf3ONE9rCvBPQfmDygf8E3YkTgMMqVC+mAi
5wPrHSS6apkH0J3qYuQf2Y7vLApsTxkxYALs7a9iAkH33mkcZa7bvevIYpB7oKi0
U8vmQCbHb8TaVIGIDANpe2k56VggI2bcqBK8wzScTZCBH+OLzi7dHS2ZNQ0CHhMJ
ASdaMx6WVuJW7qb+aNAf333+umP6X+NikcBM38yvWgt2R+4X9hV2LkEzap2qfoGa
ScHDKvUTtFwnVCG8JRoNBKmhAMR2MqlvTivLZ8WWHFBTWNhU/oqyXHrdxJRCtVcx
zB2sh3PLPzd3iSGt3yLh5ph3or3iWwvUWxPo2M3ShH2xOypRdwt0uuY1vWA5o0g7
x42nCilLOSA7BMyIJxOhR/wTHKBsj3OsQPG4gdLHBCXGdTMNa5spQqzTwy/fOR/r
yIhjbHGIF5flGkQAvlrOjo0/uHsFceV3rDG5pPCNtTLpeMxA2/smwHwJoqZHxFR3
AneAPlKsmw5smQBVCHAX1ljsRYNLe6LyJFWFVFzuh42gPBb6PW7yNlErsED6azo+
UWEqHUQ3mxL/Pd5IyD8KjnwxhfBVKZto4Rbfe+o75EjRShZnxIMqVHjPRhjWYxVM
LbZ6Cw6pj6DuNvC+gW/PIgVbtXg2O9NNAbL4WjXEDB9HtEGK59JaCpyhDjT7mbuQ
eWseTINx1rBQDZMkv3DQQuLiXYkfBXtS9+pq+yDMq3Zg4TmtJttkEq9hRgz0TUic
PUj885z/tFEp9+4O7dcGWhbiZT43bnv4P55Ck9MXaYXROgezHjENKOFbPyjU32RV
cM/wDh/eBjbJ79qkVmK98fTo8AumbzLUtHMozz98Fjw8RTrRRs4VbqjIifK8AkWO
ptH1agaeKIrKVZwrjamPFN2T5TfAPlkkBCXsZu85lHBiiIm0tuwZKTgad2vklxAZ
7i++bVOryqUtDntwmIixsdceLL1tAQPM3GeMkbjc6zfu0CiOd9gzwt8iVx/voqSv
priGvOwPQMKtiyb7LHeI0kt3CFxfMGnKYNpVDj/jib+nI5ND1fLNSnA3Ek+4tSL4
AaLI4b85dMsBUFVjfA7wtBn5rzrMeXJwZ10c7oKXgTHGYMSDYd980sbVq2GHio5O
W2oqv0lWjbzLvDEX+JbRGfzShh84swQ7ufdH1WfN5m9+lBIBxJg35lX8ZfK2Scxc
KgohuxuH+/z1YdkNvemV85CwdTvYpGX4eKm3Enqh7E1ShCrvJE26PBHBDGPgsPRE
pVSWldM+23EHCzaXR1SjYou9BzYsFOna/Wxz2y2zx/2TMtNDIsW5jDZKfoK4dBHn
9pnF6VZqKna5CF/E1oqsuBR4FZPNL2VFpaJfqktw4ZsbN3/wJvlLjMFIUxcZdDsS
wog8szAlU2BDm3PnA8PLvZcRcmkEv9GixJUxhpYKQwKeyNn5P+20IFX23H9GgrXG
/YXf8yLL8GdCnj9SHGkZ2dI0iBaYtCw5nKRG092MQa+bBSaejYYOfm5Uy9Cnm+Bq
8Dj+omDSHhzgG9yW3GOsndUGAQVsF6nf6dY1BYu7qZ0HEufftjBu48JM+wGUUM7T
NzZXTNs7qC2qQc82bBo/jxsPosqNN8VMOzNctjsRCbFQH18y8B5h/WEj6DzJo7zK
a+3Nkzj8DIEyjKbqNygKI5G4BlomDdI1VmToRtlPXKsbQCYHoYzOZ1MJiuxR/1aX
JuE2G0TaD6ZZL7lmy82HRfo0aHGvd+ZJl3OzvRCp5uL4RxDLkQ+kcBVxKECO/6J6
cMnXpodlL7+98C3wAX5DdJdaOLV57TFN4XHg14Zft08c1IA8QTe7X1mA9JVM5rV4
Jna4H9ZMcE/ULQd1OB8NYm8s4KRlwKoecRkfq97vRoF68cZTt/wDREkXl0cJeq0r
SNiIk5EYV8G7JJSldTJREsj8Y6XgiKTMtzvs+OK7m0EnbNAsf6NnRiywsIXu/xIX
bF+bFqDYDbm/mreC68BNvmpX/RWecIeg5I3oGfm9kTsZWyXKQGyGcVld76Kj8AwE
kfwvgBOEip8lpMzZ/KjyTn8+lLP83VZzarGRKpyJUzufHKVewoAXNu3seG4LaPZG
y1MAVmXb0/vsgzfC9RxjqJNTsJ9oHxtqnQB1AvVJd61VkbZr3gqp6OqeiLOBhPY1
u+09RszZYSa0iZfSWlYruZddyK/pAdAbGCQ12Fm3iPhbrg7nGXKSYIUJOtqwXCRu
/MW2kxO00TUj4aZiKDoElSHImUqZA0TRllt6NMP92Lh/HP261c4iDD/mhiHbjt3T
ZoTqK4BMJkUAltIfPSU6YkUbMP5ettwPACoaV4+8tLnwk0oUArDSE3ErB8l6mPCL
vt0qvyb5V0yTSCckMQy+juNhexk+ZtIYBnA07js4wtAd77/I4dFTXPTAKCOda0EK
PhjIUusVLVls0rV15pwiP3Zs0U824eYf06UTAj/Mgelvq/dt39SE3UtfdJQW2zUN
KECv50WrXQalRvzlHR0cggcyH8dhpj6CjYL8nAPyXege7YOE3gDBZctIaaFojwsn
6fK90XO0jBey0Dffiq2yKzHLERAEasPi7xGIK2O0nRcIElib8PnQlP/tJ77yy7IQ
s5GU398cK0qsf8YK3Mwn1dqEgEez04cIFiWaLW+DzjUtpAFa+hdvJF3CPVnsb5iM
cL1q4RNxNJi/MsMw2E8bddvUC3iA36SHNaY1DCECQ+JBamzyQr7m2Pr6Ti2YEROP
FWgamKdTw033dlctwf9rzeLcvCIODQWMCe6+DRkOQ6cf45MhdVHgIkfVjf7X4jkE
AouL2ALRf18xb5crJJPGiu9Gtni9YPMtI618IO9Ec/K1RylRiiGujBtt1v74qNoD
nkULK/ICDxJ3FMCjBSzCl5w4tAC7IqoZhAIuf9/f3srf0eYCqCKswt08inOzrmcH
Gtf2XDx1AHNGw3PxkZ6DzLrWTmq0k9GCTQHkCERYpOtD8HHavVJTQQfvq6LRM94r
9p/TqohwirULtreW42i/eTpcHHeOaARh623Jw5vlKpvYzq+qQSzuZXEDE78XS0hx
TIVHw3NrsyfBEiAqbkoNRC9n0fv4nBhA7GptozhfXrJ/P7uqbAdAxe4BTphknAw8
aZQed6La/Z3ax0a/9V/1e8abmMCLaljGJlT92f7XnBQlfO0k6bM61lAqqBKPLW6b
wK7TmG7/o4xvO/CG1F9SP9qFAYgUPAeH2DJiGxAgsVGBk+CJRoGtciorseFdvbcU
WqQcYyghMsD9KF63Z2dgyk9xCxRoKzdnofysU7/AjKJ7wYSudw9mgtBU53XTfo4D
8WUQWuBrop4cCstHcUs31cCwZhh24HrxIchF5Dhp0ODMq+fZYnb9QKVDCJO+p55A
ed4EOOmKmK0fRhz7oVEuPqWn5RPaJ+wbIoaGebwGztFUM+wzKzKXqBzm6tuZbbeH
W1FSvBN4H0iTiBnX8z63qe1wnMgC9ZbwVUrW3NEOLoMeB7gLXbRB3/tiU4OHCDbr
jPelGPH1cbBcLPSpDim0/XHQMelQ2vjpijO3QxXipH53kOwI0s0JVWmXHAQPCCUg
bg/GaGdHjAQHJDBi1NwFrlAMsRODykRfzHLXNM6JPvL2Nh808no3B5xbsxKJjv6B
wTXq3tyHRADMrEELC2LCk1VdvxsOarzlXl9XwRopi/QK7N90SFEeH/8YBi0i8ZB6
zDEzTnVD/sI7UqDsmBDIb7K7PiwBtLWDQknso/ItyXgSIQ8nFUBwOXePxzEncI1C
dYD1kPY+mMNhGXDbYO0yl24DpcOaaENJxErcePGwJHxKnCeMKl/jbXrZ9GRvvDjr
G4uScVyBaNfTzkR7aLU4i5A2DHRHxB4EpVLY8R3LJhzeLX1eXW9LnbWHNp5y+6IJ
Nj5ADBzbb8a2xPzsFtX7II38GEmVPIcqDK4Bg8IBqYpeCuHFNSGqBn/pivtwD5IB
zG2wUe00sGZFj/70rKs7A/RzLJQxeP9eQCeWDaDcVW/1B1x4qVCYZFAhxv2ArAXO
WApJuXuQSPsj8hdN+sgvYihHyPoYUXYIca6bF0NB2FlDjg6atrJzaUu5YX4ah3L4
E1FcuvGReksFSyQKMTbrtdV3Q/e9SXakz1gNUJ/GcvDdfXXVkir/Cw/92C5icWAs
1pvgDzA++ENezYJIXT0UpgJvZwPWbid10fUU8H69ek28XKMp1G0OikW6XLZjVuDz
rdqeZbHPcq1mQxVb2NmTXXJNIxYZ7uTYltFubrzEMF2m2xR96Uz3VpTW4fmV2kLG
rL3WxuMQWNDm0eDh5PDits4CegNdKXov8nia3lMjatzBI4XYmxOsZQj8i1f66MVR
F1rzM/KEoRBCH59xC+mfzBmWO8gnfhjQ8oxDgEYiy/50pNK0E8ieUuQgM90EzI8B
UZQmWtDXiDy+KNqhXF4Ca2GykROv0hks/b8dYGxUIv/JIsPCK/UvSLCIUEtEkA2+
ilQ6KutP/Lkcu4HJRGEWe7zCfMQT+0FP6P2832K407MARNsqdZZOCf1bXjjuV03h
7dRMIvAADUm2+a2aNjDTjKCq99MO8J+YMMDnPaZtenHXQgobDvr26sb+0hDHU5jJ
7af3TssaKatT9hS5+aLLk5tT8Jcm/kptTlrzdR3yP6WKN+OzjAJTvARQM/xvxwG/
0E3iRXWG9CDGz3LKIpZGTn/M/hGQXI5eeCxBdCvkhS15X0/7Qg+8Z4nLixbIoGdO
cNnIWbEy+/IOPIQXD5D+6szGFs5LQE3v40vfXuXJj0mHitw7VkdoA0rExd5uXnWF
DCcQwMXDC4H4gAEHamBmXmd9M+d9wQYlnXmp1MK/PvnIx2wPAKs8mFmGfViH+VnF
OGSPVz7yUZD/OgDuIbdVYgISl7lQZ8W+F6qKq9x8fvbA+1g9GmKCgEgVhf8TFXh2
n3Y8Jt5Sq+/ELYYVHDl+DiM91FKHRSGQjJj8M4AwCTUeMh6H4CTA6hEmxQ7VqRTY
jhkNXTn1yZP3wVOa9Ej1oPIFI7nAoow1bSL84SyDYmtzyRdsNDvPe5JNw/kLeR9+
vlJ7LNSe8TjjXbyg5IHJgHM1GV2tU5RhEQWdPdwImMbZUFuL4Bn9oeYCnyUiGRVb
F+5BOvTOCiJFKX+tJFuQ0pQFrznhUPDOYeg1P64jSOTh1HAv1Bab+0PRqNDtv2ut
iocv0D0dsrScKqwD5/7uqwvUrgnZ+6aHt+UyOUeY8RE/7KebWBnQpfq7WAfTWIPu
nXNP2mkwe24MTtVc8+oe3n7/koryHtZaZr+BNCdxmtK50ZHjQaSm3BWuzDs3HG2G
U2ZtgB7bYyJQj2YOmHYWtp8R79tOAcsnQ/Vk0/9pVKdPEcffn8zg/4AYk3GoA7JR
Vp9Jnp8hPQk5n8gCLT+SdCsPq3e2rv/JckGyuEQKbjF/Ok5lixa1v5KjG+sND1xY
+DvhfQ6PJMl7Gzk38optr+E6pt9wsLm/CFfHkv1LtUnqMXCC9WQ3dzJP6Y6+ZZAt
Q4z4XssRqLohjxxKp0NCKMBeP9Sv3j6a4CtsvABZ4wWQG5zRGc9CHdjZ1I3igRED
DLXYr/H2xPrnZxng7HG9uYPIxlBlrtNvkDoavfuGgekGK0QyQWop1FpiSiBjvJ0/
nFxGiRnEWGPmAPoXyRNA3tJ43Txkcwkv+dnts+0kqgxYBz+j9GscI6J5CijL/Mmc
HkJy/+612DvRy6R+8gT51jGUYe1ZcTmgRrsFj2vdbpH75jGtycOdtG0E/tO2NKso
NzD5KLgKPgsCDWSVRvFWxmP3Pf6ewRXHfD+uBE/blmZ/u9U7Vb0diB9XRgzTl/ap
WyrhHEXQFOJtHH5p6eyu6n1Qes5fBsVfPoJQjrd8quG5Cgqy672nc2Yc9WiAeMoQ
DnnNG8FYiYwtBgiwjYV/8EBnY76bSngs+9noUFFbuJ3YCLy92xLsfuFOnv8drlY7
n1vjfjw/fN+whhRwjBVHIR6tIHMyJPuZP4Hg18liX3RDPDsZm0ylA7vCv3UHIYxg
vh4Un6ETWVkCBXC9ikWMn8/nNDCUZ+CV/Q6TFWBgpHy9Qv1z1xPLBKzryx3H7Zu4
UFcfo4J0JJAFZdYsFdEH1fP8KRH9s5ATk5xA9Nrh4zlPAC1B6llqHXjfsK+mu9mK
mhPYTzv7U9bHVKe14gLP8eNUKRXbrPlsGSAEmqrlLA906CQy/I6BzrTs+Vpe/P9L
5httH8aZ4i0j3KEiaAmbe/3Af93UbINlPZCdSISJnCmJMaXUB/atI0zIzyZlBfOi
HWcFjJOMN6nbupCfzDu3R6io99SCIdgM8ifKuw6oiWnVQxrLyZa+OQd5k8NhOdPT
RwFJlz/NYfL+TaXV+ayQ5NztiZxXV79ERiB5LQx786GPQcoh6Qu76F6fs/a2uMws
D6e0x/iuGHnOtL9xsI9jzqSOXZZMsXX+Yawn/6DYRH7qkV4/Uk3dh37hTguzruz2
V9hQ4mAhJ5ZwHCmxUHxc3WTP/ClqCjPbWmQDBAVsKpDSpXmDtFtYLigmPdcwAmhm
FW3Tptv+dbhgVwtlM+Q4Myvrj7JNT215UNOzN4HBTy85XhkOUt73C1+3nAb6txgo
TNZlQ4mOtjxYWrRogl961ybTLwu2Xxv06ZJa2VztcsZiSuhgsqhAwYcv3PJrgqEY
7zQriUlAw5zyyZvgnwc53uchLFzFBVYX45GPhANSs+Kz5nusH8gh4c8hb8++6c6l
vsF7e0HwNVJDrdQdvSV4pcY9PbeA4M0EI/mzhnRwjkFLseZcpOMJNP84wHgUQIJf
inl/nkQN5wbTJUs/Xb4gP9KvAT6B5v+y+CFebJSaLEuNxNIQm2UX2EKL6Fr4K3T2
Ml3VtbB5pDM/ujs7fepjmLyHQJdq9qDtwt8+ftBOXA80SJ3WwFpkTKcsuqx+XNZA
B8wN2oOqOmPosWmkYXEeW4wE60ka1IlfCSPvtDCmKDcnSM159KdLuACQemhQWgIA
cWF4z9333sZr3njg8iuWXZ1/HK6v0a6v1vPkiw/ndqpD/5pNNBHbBBcTCVS4XZSQ
xmWtUsOqYvpulAHwf3pquG+R3wFL26uyxIDendvk0bHng7mXvqtDto9F1bRTNRjj
ERdNdIWewG5T9VLI2PE1W25C599QmV93sbVGaZzq356RTIq7EnmoMRskHZBGATUN
rXyu1Uo4vDlId7wK7O0VJF7SJXaHa+IQvBC+/AIRMML7e74MrxWZBilB+NGnFc1U
g7M9XNieW7KYFU1h1tW4OCbdxqYpMGYR398b1NCjaXSBJu7TMY50fkYZoZvDoYuz
YAhEYtl+nPgEv7OOVg04av3r/qhawYMwP8nBUdosIN8ggeF9TFdGXtgqkpLzaE6i
Sw0ILSkZL1SlmKpWZw0zT94nfVLtIWQigydOWW5QEJFJHNIGkc/yIqARUWOr6ERz
ejshmDTza90srfGwtPwsCLk5S4mfv/QU9JKOH8ZF2HR6fze3WlizsIVdpLcjyLfv
wIqTkHXZvYjF1h+tzeEwti9OO+wgK5k2f5AD7491JS16sEXIPNHG3YOCT3F8EIgp
WqId4e5SsngCG0uV1n6VCfk39VxrYfjuGYPOYtV+Z4+tySIUigeeUrzV1QHOf7h6
XfG9a/KjV35RWvby8UrY76t4eMaQNldBGG+xw2dAko3QM8s7qxbMS2KQTV3QOIzV
Lu+jPCh4klcbhzy8WFxF3ZPpqcKyCk/PULFP/XxuefQZJJh8pUCSaHIUBzJbOs5W
EPLmeqSVfvBxBuz4wt1AtpRejbdKRDxlI5UNkTO+N152yG6Cr0SUtoiIiu1h+OKG
jfkZYlydawY+dt07W5jhDmPp9l+Rgdqsc2E+uCMiIaNj7hhs/naD8zjXrknMG8G5
GkHVE4YUDweBotdEDVxCq7vntJLqfHMOk0RhNoO4CFm3/v1F/RO1TRgBo86DNiTD
zA/NZMd1NdGZ9vj3zI+AQrymxyyLrnfBBAmu+HM1/fe90yZs7ys4xnw6XigMlJ/6
1+FDzF0mBSfyFHsnSLrwcKxmWVBBhE/AUL2SjqK0R3NPiQE2P1JYd4M3X2y7xQdX
THhJzPrmpqsArAFlN7akh6Nc4ZjKFLNSxmIobonhjgotyDBxq4fI74pp1Aqejewf
PcAGMnhO0TU3/s5oumsYCpWIv5dWXu9FLUO4fVdOceoKlOLqv+HqlVxz9lZLNQoX
Ew1+pf6SoDCQ9MXdEgEdwcW1DyLVyob46/oKo0uxBVZZD4Zzu6ooWUQnLecPBXM7
Gz10GF2Qf6gqRVfw+kwKE9paggucgCo0QWR2E8KVy8YLehVbJ3Ey09rtv4HvF5Fc
hsSu0a8XFpjMv/nnVe3z4561FDf+0PFDsr1T3K1ir7jszk80LNIUGk2oFAOQvRgR
YGWsywEUdhZaOeL7rbixkKkCsH2oSm8BU4WR3vzpvQXRzFn/JudxNbSvOedyQ9mZ
E/17B+3uQNI6RCxqViNmltJW1k+vEf0UcXTGOG2WPcdzSF7V5eARlCrMZpGIiFFn
I3yu/fb04BvQFz1bkTCmganarwyHCKdsmaZCRrA0NyqUTo+xgcPtQofKYNSgxJyh
P/sQxN3OQ5u7yxureA0ezofDPge2XNajNn/IcLZT4VZqNosKEx1TbRCPDuDlxHpo
6tXMAi7W8qUGKx0GMVc/9Io6jdJRkpkKQ69go7jeQrtadf+I7JRZmi2+OMuhEvrg
JEjmO4wL0MZpbH+Isy57Y6KjMuJ+JJrzlR6AtwVZgWzSdpGpL6LaozHOqdMAXm2w
61MawXbKdKMjWctxjmNaygNLTSj8q4Zp09dhwGLvooVHevqIgCtstZYjcDmozxfB
05uwQqAKqY1n4rwAU5l1yfHVkj67LhyMJqTRX3DRG0uHedhT9sIR+pK9b7s/rvI0
WyVJADE40yygbhuqOtWbBacHOSUL+IEU/yTuOwO6qREEJCEm0bO9OP2vVrslb9bq
+TKiA69wIg/hkRxvCWJKnRz0jLKLTjnafA3A2JytEm/V+QQRYRvfcXItkzBrE9KB
Q+8F5EYKtK8usp8jmgnwsxAZZthZNanzZhNAsn+bUsftFZmnlXDX07mveJ1zXaZy
z3vXN4Pr90sMzP2BRs+57Gp85I9Tra8obX6lQCB+AHv89HFICLyyGxy8Uezna1k4
BNFDrq/OiucOnVR4gjipxsDJ3kHrU2vJbx8oCZsqWf2e9lszlbN+0f5tVBCTGodE
YKoIP+agi7EklEZjwuz4AFHVb14QuIGPCMG7V6FylXOTrDiELq5IVUBY6QfVE45J
L/P2cWGCvg/a4VrC9POlw0faXccpjjW8YxxF1sHcx3xDFbOuWZmh85gZ3mxGWNNu
2yXHTSupZ7eujMIbrwTTCNXIdeQazdQlsomA6X31C4XQyKDQcRA8z2bJZYo8INxj
QgnyA2K5u0gPRd8++Ac2YEF64Fq0Aluer5G6pcRgwLnXcrOzlCICLbm6tW8ooqID
MjNx21VfZQF8ltfColuIW/ntw+z4SY03KtRNtj4jfFx9I6CMmGLsu6dh5WJcPjVW
izSkYwG5lWqX16EDm82ERjgIlO/c6wzoAFQkhmnC8DUF00/QsNB30F7eJTmedB00
+zgOnqIOTfjx6cwfYL8yiS1uqQ2CZ1XGcpERQESrpwETyclYAOw4vg4q4tLpxazn
h4XQDSxKLNoK27WhCpFFmTxKgep86grM9eUBpKaUj9b2RiP2YSrqQF4HgSIGxjRn
Pgm7bkOj1IyWIigM7xqjMEYRRXjgOzabKhfmSCz+17cfCB6YzZv959gRNtOPxLob
jsB+2uQhmDARdME5tn7pEL8KiFG/leOCl78PxshWMDIu2kkfi1ss3XsGtwSxXR5i
GaKiXWPzFipDOLsFG2qijNq3s7OfuLtyz64EShpT80rhwSXvwzNvQKki88gak/Uj
MhiPJ82Spri3DWbWsY5V5+V90f5J5sbDE4/4bOY9BytxM90IrKnPSVSJV8DT/4ww
EjJtwcI2CBPvKj56CQ0WOSdmna1CDVappOQSY9uKJQnE0tXbWImFc5l3lAJL6ISA
CjpqyHQJCJsk7xq0cc3MHb43DRYHHfKe2yFjNx793onOwwDEyRBrhc4i5ihcOb97
ATXlSIfYLTG6e1otWL996KEgD4t8HUzEimMu2CCiEKHmZq3VUvP5+AQHaJmDLt0+
586ro9EmCsO5nfXgYkevgqwCXdGkfJ9hTn1v/KP+Fj0rjQ75cFHv4aQnAcIa0Z58
Q+DLjnh6jikuTqq3sX0kcwkVVtOS6lKlMG6u55wUl8qjiUeS+S+YkH86I/ZgwKr7
9pMpgax9ESiyExLwcnXi959hBRr6zhbfdhGu0c3l5JZMxYwK/6sHgc1spa396yMS
E5YxIrJhLnBNX1STVAmBX5nAQDolxsenAjkfcp0VdA4s3MRHlmNW7Op3pJJJXgui
fbhBmuGNz8Kg0oQ1Git4hVdZz/7xpuGMSbMYUUDdnWXqc2zEm0Mo611Pzw16PcR8
rFLepIoIDmtmKCpzTGCzB1AEjY955ovdq0YuqQJnjs7nXAuo5jbCAEwyW5dc7bos
p5Gs+EkEyb/3WHxx30EjlPoOQbAN8WHK3M+3NZrogeXQl1UNWz2JcWVi4cXgsD4x
auoYEMLDm1QNaF+Ae4ZhssiycnnOGuuAh9XYDcW3MTK/IceQ+UP1VsLokH8oDt6k
CWXmp3hoohI77v5EW0HbABc3QPKEpgEMweKq5TpMupXVs7yyFYufco9ElLulyOo8
7sZcv/bJod7SIQsqq5phFpojEFTU1HS3NKLUdw6bgRrzRjOLidi772Pc9aFFRcn2
D/h0GrDYJULChUM0VxT5feYLaB+qrRku/tjhB32BMAhjNqNuya3BoClznZzXDBw3
JN2wW/QPxMq7SvB99bvzCvwn5dAIFtifhuHVstdcb96vo+wWPsfq7T5uLHUUrrcW
w/6C1HXOmamFl8fFlQEmJLmpBz9RYa8qmKP3fTXZdHr55Mw0snM1FLl/dWhd45D7
WnObOD3qFL+d2fu06ahz83OEoQmEymQLxBHSDUt6x9PmPE46UdjUfR85wsyjoiwG
zKzBXzLJuXO5oWowDjhCPaHaDAs7ExI8GG+YWUDuFymaPsAPWcnpaPuveb/nVn2k
lT2NJ44orZPmm2L43uf6yA9Q/pxNylf7OXLR6iqL69SEQF70UhchV2oYL4Z11JIi
klQYLizVGdkK2nsbFKKRa5SisKQcIbh4eyjJJoDeojFRRA954Gmlb8k0K1806ykH
013hLBPJgQ/woGRK2xuQdSf+Jz9z3fgCgGlSO1emLtNcjk0C4AT/O2xmN29dHeHt
TJ4j9aoAP3s0YGvw1jKDnDdwDSZLsuM0XAesiji0sXVoUGO30lL1N95WSQcPkEm3
TZaq6sE9p2+Yn2A/PdiPKAlgd0yThHXb8oQuIinz+EOq5mcYMVJFS3ecAjxD2Jkx
Ni86vCBMpRh60O1uDBLWcc211ChIF0F56DTO4PpqZpR0+2KS+e4klA4RfFDjADap
nFMV4st441xX8bsTAsGy00xgVNdu6OBK91CEqLuFS6U0xzjmqokclv9dOZFUowSZ
2uGdNI1/u7oLJmB2VGyc15AmH8hnm84h+yqo27eiDQTiTCbeuBJnHPsTgjWEsUHT
CxSoUwW+GRMKiPyLzHKbc/HbMYOJS091wVpmLjNtu9tRBHqohdIVWtaLVEvsBA93
R3eLqbxuGdeIoc61T+yQjOWxoeaJTgXHeW5jt4q7iPkrtQnErto3/VfplDrMuHXw
8hjbBiKLAtdhTw2R4TOvKtnSbUEk0BkP/Thkfj6Tsa0EOzQF5+mTvLil9jUkvhhS
ca5qeTClbpmAET5rPfCqtaRsgdrMsC0VVODYP/tSMxDGAx5sTkuECnuGOleWVlNK
xdtgPzw1FI9Znr9aZ9hsNaj1fzbAGJuzapH+dhq597zkhuGOyxDckk8KpoJekR3E
dK3Y1kOOWYp5GsasMqD2Kk9qrkSA5JeKDDubawDkYoZCgKR5fOV/sUkT8tQy6flS
AqwFVnU8ITftOhrCfO+K6OM++bYZdzTuNSnnPHJfpAJvpFmdDY1fGKIyDEIP7bTn
qrO5HhkjqkvKWSInk1pKn+aPTcNaCoa1D2gHu9bG2TsUnPvaY2yK33tYNCX/5SFA
OsB40hfHfFzlEIsH8q1Zc6YcydF7r72kPE64i6hFSumIxW+CFgfhPcpOjF4Sq3I/
xWDfWQAdzvS11RKlPlEq1uuRKcW3FHy4lGb96ZUhMtXFx9TShrPccqkbKqjCaa5j
+Opuc6FpHngfh8l2oz/N8dH7UuKYJtdkykQQJnrvKpMItgiB9B7ptZH2wNrF3tmF
WVt/S/SkfpIxN/RhDQq2Ey+jzj+x5TG1iOWW63PP1PTOBonXezz+8SQuyQh9F/GF
ytKhy8lC8UsALIcydVMJ6Vkln6vVonuFqgDSyvvBSSvnQSUs38/kjUFZnXvkf4VC
eOKk9Qt7sfGVoDpdfmdJwuRJxl98e8hpLMfmv8HTEWS2+W2DiHRhWM7jgza/6LVO
3G0oIhvY3VbDJKAM5s+i1jGmkJLlHv0RLsXfuiSrf8Z7NjBuX3m6/3/IeTcDZ6KO
M9JEubjvhNuzX/JKhikQpW1mYcUAw+i/1ZRyk6y5S5OCeqKvym4CHSafpRnhDgo4
ItLzttDb7tDeAzBYAzh3iJd8DPFTCixj+7Me0BJcq8T4XoO5dXupGkYEA31YpGmN
cAgy2UDFnbKpBbMdKX7NgsEKDFE4m+/YM7YCsgZlfubGbxjy5PSSUqi7MVbq6FrG
AxApQFfwCxH2SAJEKuFno8wU09oc502ab57imj4xI22970Dhi2/cPYh+6Obw5a02
akRcd8dtU13NfzUwmr6TR8jwPBYuYTAUT3JadKd3cei6DDe0dolnEPyFyLTAKqja
u+phdLhzVe38Rqu2Ba5YbZwMaBGoMwLaEeOY3l07nrX2VRiGilwWFYOXeG7odn8Q
jAdWUCJ9LpLAcN3Ei1jNMrDMUBjMvrQO0cSIQgyS2pm2efh3jyhK+365Y8AlViUU
ZILcR/CGKYEDSb6zP5SFJ4US4Ib9iDd4Iz+R9kvqBmNhjNTjUMaldRUfRhwe67aE
TmT9PxeQJhELxbGyQLustIjJxhUbV5Mk3DUF1gcG+VVX8kCqo+IplMhBZRI79jDY
Ew/NpIXEL9ea33f4iYPyWTdsmJyxKV6gUNKIelaeVrQm1DcaEYcDmepPh476YSJ6
45/nFMWzjizhCET2f1W4U/qdAW1ntySl46nYw286MTaKIHVbQslts6OLlCzoUO4m
1Lbr11MLFd/0NnI2OP1t1V4QXmzkpRZdrpLjF1r4S9KKbB8wLoUcvtHnH1tG+xVf
NYzRFTlmppJwGNaxFqOv4FjGpkVVp90fgzhMHxV8P/2T480IFcz6tD7fcw+fD1gT
z/WdqwTE89E/UBlI8gj103/or4jo2e2B1NtaFE0GhfSM610QBC27nZTilcOfbya0
uUp/mQteDmLY9O8ouxp78ZJanlDAcmLdqfhld6THZeflfai4S8ZAwhWp36081hvb
Bu/q71zXgUiYdPCgcon1tT4TFvZfEojKpeIifxsR/AZWr53tNehCcqHKTAWWzz+x
wY/jRuZVjQjrXlcWaM/Odhke0heWRFF3hZ8BXK1d89q4+Xr7jRMPm71ZBCFY98E6
2HZHRvM0gDyl6ITe+odogITDatmuJY1MU9ya/yuUKBt+I+K6d20to8KyrxaF4pWN
uFkpSR/idw4xEMCVwgCCG9/bcrM0TrY6okfbms/0lz//YeUJkNp14K0QTArlmflZ
CZL7eW+HpYjFOUBq2tS6eUsSARRv13wznh2SpIc7FlfcC7pT9nfbtCYH4sZsRq7h
d4nYe2/iHwOARJQcwQowcXTQyZD70ZocrDltce01xE6hfN+4rXIwNSuKLWm4rIW8
vbA4Xe23duEE2lRmPimNstDFMFihN5oK/iSuOm3liZELON426g1nr8r8EHVisKKo
tZCzegnCxNyCjonZylAyQOrohCf8cv2u/IF/4TLaSMBbnsENCzyvkhmL5XMVG+s6
hJHSxgJXKM3UdnSByKWV/rsorpV6rUv6UZNOm34zlNgQ432vxwRf5RBbQHejZjl5
z4itZ0h2KgYr/UK2RTqeKsoDTR9rmQsSc/DEDRQbuZgXgrnewsWWsIdfI+dMQnWW
EapYBJLsV/qJWpg5P3EQ7BvJC96I3uCD8pML5yBTFvJmpJ35rPcn933x4C2P6Ev/
mmX3PpVuXHXQSPzBt+/G1hOW9L0y/476uoZhgP+a4crGQ26P6OqQyMOMYN7+MSch
BPybuAnDdzBAUZ+phxAfKf6pJ4TJ1t2uvrZTIqAHysnYDOOwrA2dNtxMd4Khy9tc
r7mNd0k0DigCR115ZWu7g0BoIpfXHxZLim+9NH++JtQHFTs3Q8sPl4Ud9wQvrHWm
BDJECV/79hJQNI2LjROX5Yj43CWtLtCAyahPMCseHyAP+eb0AG3p5SIHlJZ6qvzj
gnvFuiK04n4iRR0bsNUB6ZMNl2gt+f4FWsV1OS60EfbdGMC/2vzvyrdkONXEhoJV
iSDRWWHZacUHpfYrkX+Y4XqSJG6CmYJMR4xNu9cWgc6adLft7S2eSEYRXFO7CKvJ
WGunkq55/pvnSo+w+M0d8Kj1nF5wTI143NiCA9/1yaslsz1V3kOP7ZfTHwNVaj6Y
KfshCpA1hgeme6piKHntpHwbstCeau5h1xDIH8bF+GcmeB3vHEMjFpqiigp+FqJd
zfd6GMlFLWyaTzbgzD4qBe6jl7fs9OWk1Mo/cNnCbts2GLivl0mc9Uai3HJs3mKB
IbdYnE4TVSQtqaN9XcgJP9l9BRjyRf1BROPlobz3MAgpAcNriXwcTwZWFG5OKUx3
MrYhAlK02VmPf9EyBbNVaYZ6tMScerYPZwRJZkk7Ffx2tbq+hthmT1kz3zKRC0Vu
w20/i5FTs5VsnOPi3IZgAPcP5uyrb4mFjeL7yE+7fwRxStD4WeE/HmtGrZY/GRG5
bPBsKE/KPzxBCZNh/le6/alEuXezBd/nJucdHPa0mpmC9j+59rnJ7QXunNvBa8xH
2YbdK/rOcfJ2zVn/va/kuwDR+klFOY2B62jP/0TSv8s+NRzYmniRLzoJ6kSk4uqS
bpA5Smes1x0B3SR6Acxd4PpHaJLkCWEkfl+4nMIeFXAe+yu6gyFQd3XhWc3kwhaq
wxvHKEqQl1j1dSJORW4MZP+3YE1MVoDIs8o+ocq08IIcohfIVNsmvcnWkoadTLin
tKzbSiVsqVBe1MoEplRjhKyFnBi8r56cpZWQII6yvdQeRV6paBgcwutP/CGy7syg
2Ofbfc6QoSqLqP19/f2ttRVnZ1NfDFiht9VeZPhKq42ZTxXMty1x0uB1IE05egAL
ZpVojoMAi6Jf6GIYapxW1Vdyldu6PoveXij53w/YpziWw8MDIHzITaIg4Ugsu7Yb
IJhKxrCzU0XmcpdLAWVBJdtZ0JWtFDGnP9Ys64kCZeBKy9VTUoL00IpikHT4SO0N
X8DarpoCyvnSTLn6cLY5cvuBQNZPuSATiZgURhMAuQaNCDtVJ+TUC1a8xRsBNNdu
JcPKR9r8TAuoKO0VQ0ESm3ngvq9jJjrEKOKjhsL60i9XzEB7qvi/aY1PHcfunVp4
tl3aubRLmhWFKsfNdObtvuIzKSoNGEhgjYnDB/0tNwVYMDXcrTICPTT/ufNL9Lfj
irf1b1tdz02XL1qbHlnf/Yk+DeYK2zdYI0t6kQRpNCb5Ob5cSgG80TJZ52dmY6f6
WosGmgZTFFWhzaeUy7xUZXcv1iGdQP9yFttGoJvJZtXTgmvFC0W8vSy1Yk4++9zz
7v+c/hcvpKJ32fIrMnmUcT3PP+yypEgvjkZI62MUFBkSHrUZODqv3PeHH3dUfFPT
tKZ2dIQH8ipnUT7Uu8vml6VgYSrKb/gX9uLQmPviYNpalbzUSUgudUx7IrMhO6Os
FPiP2SJvYZiaKJx70Ug7goTRceb43J47mmyDtTIpz8id0j4yQ2FtqKJSpW4c16dB
Rd3bOHCEYCGDjr2MRh5qenxCVvwdHWxoMptCvY1aHAuJ6BPxGhECVHrAEmEczH8h
847cIYtUH4ZejUEnFzXXfwFTvBS+Y57JwHCGl+iOXSbkIaV4+x17lYG/tMQlKJrl
F7ltFyB8oDsQuVO51Flo+uxIlIbbnL0nSBJaLglrvLfT0ra2dSYlQ0IrcAnqJfKy
zy94tvKOaXZmKTfeAhYVN7gPJnPFtNzUsyMRJcXN1GYD8OxiC9mShhx9ECz1Vosr
bEFzFumUmtRqz5EX2VprO+Jx4HBmAM74/9M0BK/4IVgSbB6jmrUH0/MbN50SGau0
0VKHFREI+VVejDmYWFe/ms04x4g/mckiVWy2mes71yKDgVnR64PxTynRP9qILIo5
pv+cwcn9chK0f8adaKJImAmtALrvj9/n5Xakscg1mAqVW2cl4qYCO2HNrDoHUTii
t++pszOJBjg4QZQqW3yOj7LF2JkZrCQeZRh/b/6NMu9/KJDHaYQFl/Z1jOZu23Kh
CCAVNsrmj30YyTcYkniqfwU5k5UmXza8kXlGLVS35wy+oFP6Y1mt98qlHdwYCYj2
ZLSyH8947Ghbu6hGEqjgp6bBGr4Lh2dlqhccTqMvIcJuOvmsPjNwUhvJbmrKVPeF
IkPJOwKCmUlg+yKsKrbeNawrOCvDjXoEI7HdfELc9mAH13MGUH33Hmf4H94DtNjq
oYQZ4clM0eVCzUvH5n2HGshD48+bs64pOUnkIsBG7FxnLUiRoK8P0C9Gho2yGRgf
e4c95qfY9C9ZitFWgPyCY9NpPyLMULmsevAQJpj63BCPXW7uI+sA4Q+DT7RzDjEa
y6yOhacnG5JJ4zskMFTubxE9HdukEk1u2ptLXwo2JlktGk3ZdcA22MqUMUqry1fG
KPIAkjBD5OIbm7yDpLPhYa1OmA/4r6Nx4hkphQbafsfBQUMoCsuMuCG6kHyh8wIz
4W3yaxmAtavXeWYiHZJoaYDJqtuyqRhHbVyQvXaD0ai/tZXB1eITknYaYKL9Mv8x
iGKDYS2GOOS0BJiGY7rqo1vXVGMJASqPCEbR2lBbwMoObb7/1IQDbAm6e4OZ+jPN
8DqW6saXYUDMQfGLc0+YLRImOWtQEU07T2gbNIem3OKNlbMdnzXvmqVDHA6IlRj/
+NWtGgjpR/MX2MdyVqZcX+i9iH4GktQ1wFrlzYVQBsceLP7A3eD58rlQGn9BXjAy
4HQXqY0kNDFG92dbsG0z2h6Jut4MG/d+n9iGP4SksZUbI5OoZyTHiPZsYsFzeycy
6VRNrJUTbz6HrBPW3SeDvlPIYQ7tlN90EC8hZgB5iYwYfjqqwZLfTntmzDnn5h4o
usdP9RhQx46aHA8BYAi5KxmNGkxTXCKRwxB5Gcgjp0a8F874Z9q8TUOlVdFUJ7h6
VvmqFQxhVWySYpvGlfxfhyD/O6nqynI0qBGK2ESEDkuy/G3hHZPzDSjeQrGRs8pX
lLWOacy0Tfg/mdjeyIkCMqy4wnP1/TQqireat2jXfTPm8s7YFQZoJzE370qL/dLj
Q9kXp+Qw0ez/NsFvs7Guro3LYXdhV1O69JJCNNKKFw56dBGYxxolaqXUQDQv6CKm
ZzA4Mn7978yMlkgjMaIwjsL++EBNCX2vcO6RVjEIN6+2HQzwm44SludGO1Z8dflP
bybmN5feZ7M118ey/LAbkZruL//fQAOgniL7skdsuCaLqUWTxPdc32TfHAia3it4
Ma3D8gvgr008T0+Xb2rW/bqI3ZrJm/RdlulKcfvaX01lLvZOn9QbQ+afea+4is5L
+gWgJ+892FHJAA2MmmqjogVjNOTx3HeZk/BIuIh/YIv7AiYtiMCzvFX2OW1vgEkN
9gcKsLimTadY/AvRfQ8h05VKeq/XNHjLQO6D+iIc0qce4K06U6IoVxm3/HIBqKJj
mtoX5oxAQOz5j5zLuzB6uqSP4/yvHMnfO9K9EDolrsPiG6YqZCOdLgsXkPV5DLK4
5+9rvoG+6J8NlC2xhcvWh0TeYHsDyvhI818Gz0Xphf030p/w/9iv1+cUtwHEmGcE
FXLyPSJuToUKAUgbtoa3Tdi4cIvYNtsK2DLshYc/s3q6VbbpDL2gY/MbBp0HveZH
NPurzFsgkqkTwjNjFS6Bmxz6X2/RWFmUVkzOoGO8/GWpMmu8IDaBFCjAoqlkkegT
qal5PupvdPyKx9t4N4UsU5XKUCcK1c9l8I1ZboQetdNeMiZg5Ox+P7eoDdv8eZ5f
WPvVM2x9kSDFLnFM8wy2StIDqJp4muzJybdPGkYCLRNQLVYmpJux6l6oCN2qGNBx
lJfoHYHhv/jJuNNAsvrLx5nQpwHW8etr+Vn1ScbY/8MCJjszbDpm3EJVoje/RSb7
V5sAhyaOqnVDntL1/H6kRCLTq8czxymvqV8/qHVtEBcEf7J4WA4DNunCdC+cGsP8
luY0vnaKQZXSZPlmC/HUvv7unzZxuadMQZ60qqYDdu0qJzD+d+cWElxsGp88x8CX
x40T2wBLjHJfQYOY95kCmmu1OG55IuyTRHfksuqaFtIsTDOSatx5Xqh26Sm5wO4y
kfIrCUpL+LBIXIkdy0SbpCfXIgQ6XfZg29vPbAyX9uPPwdoTPTK7L9nXBcR1jPTD
1zNNSz3psYHt4L5OPWUZIh6Deg8LeZ/fUvVgJPrwmHMLLDtH81+RN630ILWpYBYn
MCG3x7DLN7Rg7Wjc7kSJ7mm+j7bFT/Fh0KZd1dZOkFPJdeCTm2G+1fUtJmNrway7
FYILWJec8n2ha1KeomkVJzLVvFT9DIcjlRZOYgdt5ACs+CNimUYp+8u7DgkO0S56
nWUHa5gL8KteeIfEl/mj4eaVf8sMNTTAtfQEAaRzAV3qPOxU/0bpmFWOuOW50uR1
EASLP5oRcrCBZSaIZUr7TRocZOFobh221JzAb41L5cG0PsgMF4WHExYx0PxbxZ7X
HBgkV6gredm1tEdzYIP8KmpTB2ajFyp4DliCPtMgn/jdHDhjssWXPiJkppxKaC4v
sqJhcWWHVKEsIlj93VAJ9/DUhp1VzUr/QIsEO9DgdvbenY6MYb/LxIlvEwzIkL1V
YxJxjLAZJDMc8mOxwb2IjOcI+3xYjzLFddcJ0S6XQm7I6nyc0qu2Si67ZPkB+a5K
Rjm2tzlm88I6UsvzwXvNbox/KgjdLVu5PRdj1oiUHovqY/qqGk/11/voumhmpSxC
Db60UdGmQCQ3cBj8KZ8pkbWlYrH38KPGxMhEOx04nGMRw912hoiC2s5SzvdshE6m
J0ee1aKgPCXYvmpgjGYmevzs0zaL98B7bguaQt4H61ML5Blg+CGb9g9f9YcFjZzC
njSQE+bCBEjw6/0XNwVkoMhbVWFLCaaJZx5zCv4DKfuHytOyF+1RQWJmSNlnPjhw
+/WfrIjr4jOucGuBYTHceRQkhJmLBOe0HHWOB4vpAi92Iow3OxLGExNG+sAwx36w
XK+jwLmex1zddaATmfCTKxn9dVLaSMMwV7BCO1b8vp28i3IvNarpAkoetKeQnt7Q
DWm2RCDfi3HAhq9gtWOXLctJ2peVHBk0jXh/5KYghr31w4kFy9mplCwHfQXbdLJL
mA0vd7hU292tLztlJ9s+sBAepphXpqLsm6X/egfPIHV74j0487pM8/pHihdHMTGT
sD7RijCGqMypn4HATRIT2I7aoTSsDJHB3qlqOMo+4LqDyk9gwFdi/HYoGi6zktMp
ozn1OOscuQsY36vpFcFgfRazoElTEKza51cpPEeK2o6p5A/THOyvVcfOteoN67e6
iQWsyiE4XnPA2JeVWKxP7ij+6e87F2RCTyGLPSDMj9HUaSSWMQm5/FyPcH+1GTub
JNC8s8cOdFga1ocZvznkgVd53RNXjOcJ8dhYUlVg631/IdPm7D0yn9IaLK3Tkc9I
rlyJxFUd7Kw6Xn85hc/gNcXtkFPjsMnbAUAo3M+GkQsOCUIPxrGqI57GoH8+7ReS
fT/DVB06vDXm6r+gwgfQY3EZHsbX9fZM2mbUQIegnMI/O8xqhFyaTtsrYnvnx7iE
vK/gpuC4dS4fQjK87RlQTqCzBq1z3Vu4vB/kHRN3LLHResOMhd7QKTYtqcnfDu44
EJSqqNnvcehRkigmJ3DByxHzzRFndaff8idF2IufucXpu03mXaNP1EiJFsyYYDpk
mf/jbQxlX+RJj7ldyPCjAowcPpfZ27RnKUaJvUVlKGq+v2m3lHvFyclEIdtkfUxL
aPrpIbpsD8XeaCsn/3ZRkwRm8pHMi13u8A80K32Ecjuo4+afJrA9wxAR5o7LVWPE
hY0Ca+dudvxn/0NsfflVKMFTqujy2nReyASh4DiG+xuX94OPOCngJbKXS87D8Is9
3HpggA0Ag931EG+G5dNRXqP/10lhQN8jwQn2i6E4w69VqZ771uAmnsVRXowCDxbe
Ucc9+YvyHFTNo9YVv5FwOYKvV6j4ndawnVf746o+LDlqFxUBSA5CH/f7EL8IUy3K
afX4b4k0Oirnn8idATRtUAeUxVP1pfbHHnAwb3FAk50q+XID1q4mMoPdMi+lTGAt
wS5MLXVv/nG2K6rDtrOymX1NYhyRjVJy6XyU2s9NCoW36GtmuYVtkt66H4l70esJ
kdLD1lvzckvp9U9RqEzKHgTi34UuajgPRvrIExBjXcBXdgWdaEwWogzsk1CDojTo
L4cqMFGFNWEGhud9miXss8xcD2vMS8xyUfmJ2ToE9huQXe4zLr3hYRolKcop3FYZ
yifehYeAy45rwUsFVezxGVRgvjzgKsi6B199wEscQ8QJ9X15NS1ylkBENQCFMTRU
kQ25RbGIjiULymoLNdGmKe9qzdjvlGHW78ILh177FMYuOO55wyMzEUiokblVu0+y
o3tnyeTUjBkV+y0r+a+PZ1Eg2hOi1SHQedB7J4Pm5sR3egMvmQZcVT4vrGLwFzOP
L3uSw0UWxYXB8AHosS6L/L3rDxDzG870uKiBNW6MlhcPMr/Hy2d37BNemXlyboeq
6Aj4w581Kkck8pFIhUPHpmbSYtlPd7Q3B1XSQv8gSFnNNU3e4wPIgeSxejYW0bTn
24Z5zxLNz24l8wq+/bL8BTnnDxWFE7UwLp4a0rqCpdXwl5ztIokedv2Zm5r4+bdy
ipjP8vxMKLPtBiL7o0rVvCQx7KVNsLrAfSnq4ufia9/rVagQmGhuyzweTyhPbOQl
x1ebkE6OQyfh+NBSDeU2+YRjvIas4IyslU8UlFkAPstTqI6KQZuL9B/eiqZ0MSlX
YS75zYE+DEGILvoB1IchnCK48KjKDk0h87XZ+IlvGSOQKjpFpkisOPiajTsvQTjv
2WldN2CE1blZ6YT98H3JJNWCHusfjR8y8p9nDi7Nzk4I8ikx1XdFGDtmT3Cio3ha
Kz2+EFgjwpfmAeKMi51S8IFRJ5djMt/dyxOXGDAuxYqdReIo777Vu9ZAWXZvhjVb
to3zCnuAWnIRa8lFzBKQWI+y1Vb0ULAeJrtg9NrPRpIAZDNFTnekvQFVNjnMDXIo
ALVVbWZ091Csrj5PqrYpu28a7SIk0aLAbHV6TCIdeXb7SKgwxTE2L3F65VNnI35B
DLhOtn3FeDdciFoV6+f/837NZxEhY9eH+ZnRVM2KXUJxisHEJzsC1vJuHIH3XC/a
iMRmym86EFYEeyYPXMTRiqWmBw8gUQI9v0vYJoFF5dUGwQeoa/I/nzblw0CzK0j/
ub1XlQvHwHcCLhtUAWocozMXGFmeye8Q/5uXgBFewCdFugCNfJ8q9YKXs0DKstcO
6ynW8vhGBIgAbBZJjaoxlwFzGcZNl/x9IR9z9dv2RmQ15Q53DUilfSDFr6RGZQkU
3CUjIDTKy6pYwhCh0BZz+c/5CJROFjDisz3Lv13hKkCGVgWH5f0LNYHL5/xy0w2D
//WHfPkW7e5dEuoAMRtwfHIIaSEWgDbTprouXvsN2Xehv9eR6g1JsgZfPe4t4mm9
gEYrI9D0TiBn/e0r5h9ZdU7dOylD57IR2i2PymNofjso2kvjvtac2GPjBuM6R4nU
DcBR+ZnidbnVmcvsLZSSkni57CaAP5P87Er510X2Cb7MLLrJzqDFNFI65BJ8BJ9v
uCeYTKXzdpblJJzu/Hu7tlQCLZpuSqcG9Thb/GUQSkpyMmJGLOBfRy3BGprIigo7
GjG9wK5/SKiuFPwiekUvRAiUhgjtbB09nQOlkAldbZM+++B29RrSburLK2ikscnF
fe7Mr2jAt2WqJ5H35XPsPeXReFuudu2Oqi01RrFpOFfk+QaUogmHeigERyuZBhzT
1nXfwzyspHc9DvEvCjaUi1Y+I+4rkCm49uTAfVYiPKkrvp0TgPAJDhV2//xR/bTD
/NtOuxcWBppMufoGN3fMkEQAr9BALuVqSEkoryHicLcG5z4RcjyZ/5C+8vA3fEI0
rFIgei5FaX1aA2bFLsOKwYWs+PQ93xBQVb2zzauATkLRWXLlxucWdfLFoXCZg1Kz
zynNchJuhRdLXvqibp9F60Zt8YPEZGO/DXWCarzFQAebiLFuNV7w4yQQEx8G1I4K
nOrqWP3bRj6mJYpcQBsQip6rshg8FJ92rApo8s4OX5yc0SE80ZteVhOCG0/lzDjj
QDUQ3KQ0ftORkbCcujXAH7OvjYnKDfPHLOOSaEJQtUAQK5hongP/E/RXR1vAhafL
uNYrKN/HvkXDyNh4uSLlHra1Xf5LPgJgfbdTsgTgfvIfKV5m3QmZQcio2Ii/kaVM
6xe8I4QhDghIAW26Q8yx30LKeWbFkJKZ+qT0FbdvTstkElf/Z/WAq6KUg9zlJ20M
ou5GIlRucQLnWWmng+lu2t9m68oeLZvk4OsCGcJfqgCRJp/t+fMqKI61kSHegZb1
GPFUxgoPNxC2wSLG73w/0Cw5TcF4vfGDsEgSZU96i95iGTzv3N7xSg94hfjcQD1h
txssGOGWaYzGKFFBTrXGmL8nUXDgieZtGpefEB/CvYqRMXnomVey/WvLwZtxcXqd
8WeY1a3MetSrd4gP4mFtpBU1vDWzjA9vUV5AkiTFCMiLLYER6fMNQEVfMShin9hS
TmNd9QkotrMb08+5mhqUdkeEALcxvozZ4g1Cbv5WnFuo50BXc8tz6GSBikpaxl4v
2pdKqtoXHnU5Gt+77JLZacWoEB+wJ/Fc8n/UM3oi9EsyaWySlNbbWWgin7rPy0L7
AjSLBQ9X6HpSXEOBAxN1p7aZYDalaN/g3rCRDB5fgargiH2n+5bLsQXcdqMju6/q
/1wnhLORLw5xvlDg1CO0PPZLJDa7C3Uh+UMWXlw08/RcGA75XVe9iruO3sXDEwoO
5IpTMQmQrSe3PTlfJMLmwu9JksEgIEOcViRZmNtF5h7XdISEwPITOJLIjGWTsSQg
rNzNDd3TKQheZ+IpNIkpAubK2VdSKdGKHCKoI7vsofurGg4HyWzzAtSmzmGR/kuP
yIPAGwIwRvQJ7uP/uSJqajBm+bKJ5gfnUsWh9dLzBj/+Zmp9PpKbkucwH7le69Bc
3xPleLCeWLuHuxzwWIdjEaiogUBG0pvlKtH1Gm7dksN9vsK65fN9Lli4esIeVUtp
TTxYswvGANFbts1n777cphhjmrXyuYDd1KCtnN8wwPo6soQmyYrzjZg7mCuoGjP1
/0sh8eY16NH48BlI3XZsLRzXHyRmw4lbwFZGgBKc1Ci0zocg5NuEYMw4sx6xJplb
7gNl4LWCgsl1326RF21nm+TbSR8zam/R+SWpODn2K2ssZDo/bdYPAcrrx3lmuSFA
QZNeZSQtWaHE/mCs6Z+II+dPb1pWiesah7cR+a6BjcV1iKmvwvAnYlV67ZU2tDtA
Gcjh3OgCZSdqwulxlLEzCCGTar5xDnCXOVVLk3+HYAK1mR1RQKKAq9E8SvJ9rwlW
7A4cYwPk/xSs6BZSg3ebDiO0hgPWH7xC3O8dwyqb3N4UAp2dl3Q/Pawi4W16icLo
gaTxdSPS7M8qTt368+uusF4MJ5+cwXWP3C6/1UED9nAi425iYtdSOKa6R3shZQbF
y9gD1ftDyBocoq+qleTBs48kX1Y6M18wP4/DRxVaFT+wMKpvhE4kAcYKAoR4Veda
Qp8Hz5zkErGbI9bc747AVZW2S1EqZs7XYnqti8mqRHiDYpo1n52OSGcgH9lHuAs9
8UtCNjbeCiqAfK+Jf2flULLhOnvFqZuikHmnKkFCADrso18bHB1fAfGXlcFkHSgi
mGbiHTn4qFer/zo2i/lm9bLtkEF6iCqXE1klTVTt9FxWBaKWllmR/XqVA6p01IQS
AaGG/o2exDPM//Ptjf9hHQPLcK0VvEl/2fZP8Tb4U+n2hmIrR9GUX5rIe40daoq5
RvFyXx16bnI4VwGFLr1jx5j20TyT2v/cI1txkcwy4q+KrwKOi+isRJ3UcB8xVROA
JkGXiPGMPfhdgAMPvcA3EI41E1PUSnsUv9f82gMDTSLMaQXiADiBJNd+S/RXpz/2
/l2TLPnC+jmz/Zg4Ri+cUy5WoIsUY9Hh77tj8Cropu3fG/VsJAmObL9t4fF+eGol
J1UIUgdjV0rGgIjrmgQua8GMAIDHKq97mQd4B+WYbGoA4ylc98YCdMKAJPAN1Ee8
c/N6FwOATVs/KEguxba6XL3WJbArCQrIZo5Ooz7dGDDprVtLAR/dX7KWE816RCOR
4k94JrmAjOIwLfES0dfIxGfYytGFKsP3lkVsTVq9qHdrUyO0JtCrE4ItUNltASwE
mKoUM2QimrfF5pAugtCt+5DrcJc/a3wiCyyJ047g0C03Jpz+0/wnqOsgaG2CWj92
Oh0rarb8JioKpkqHbSMaaFplo5p4NaJTkXMOPYAWNTWBJPseyvUKYBAePB/8DoIJ
cf/x7Q1XeUF+UOyThnomJzoRBYWWcuG9ba4VPTXkoSq7dXjM1HC3SceAOSJ0Bc5h
WICIwV1/Hx2kHL78x82De/XQxyzKQUOcShjBw9hYqmUmMwW5zja83gw8Ng6b33CB
p+em8rlKQNJ2jwxQ2+Cxv2im95wwcVnaqULTmmUWFwnkQuKzmmEkYilAjOWiAMUM
5ICrnLY2vhxFq3INwB/Hqz2vxL0He+4RnbD6s75yYeB0nOkqKaFeRH6KmI6Dnd16
m8ajAfQNPowEDrnXvLh+sCsDh7POhZzOxqGv3MxZAbofGka+uCvgcLFRVR1B/STY
auKCpFNYNwcgM4JzGoUf1HMWn5sobJSr7stfcZdW1F2DqX6fyksTj7sLiZlAZMiX
Xx0RPsLXZvj5ktBhW19SuiQAT5E+Wb8NIR3c8zXSd4ViDg//XyDj88dEYBVqa5ad
JLQfm+/cOL6cu+s/6i9oBixmdqNRLVLokKTOsCQszUktEK7ROJu1gHultibVWTVO
IcEKrocsbeDsTQnw2Qny5SYvMnjnxf4fXaht1askVFYgN708Ly20m+ywDkPeTvhR
Aqcm+vuj9YNoEZG7DhRCKP3162fDZ3UnZypyiSuEWUMbp6VAZJScSin/hVr87Hye
bgrfmORUhDXHOyr95MoC5YZEXD52R0Q7Ek6pprFxUqGIlGgE+LbkxLDMGQ6LfgkY
sINAQfIBbJ5VOTP4At7Zu7NRny+XUOp1gOPHp/4BTM9lHFcGp31MpXdFAImOnGyd
q4UBptofsRig6Im6GiWB+1ESGL5l8gxWLCXXbpM+YjyDtcuS+eBmodfNunQn0pmJ
gkEtMSfTpWOl2td5Xx6gF73tSGaUxZTVqAGN5BXjGIkIiM8L0lXIlFIWTUNCN6wj
pIs8WsU1scoDwLMYezkSz+I6HFnPOrESivnprs2a455Xl10deAwyK8QP+BSi57wN
0EBAwL2NRjWo7ASPPMCb90XS7zl42vgxrZ+/i4BktKz1Rkp1DcNW76iEw7XFnxcF
uL4W7MMXwqsjZFcMcCnF52/e+VmKxqaeFx8mnzfbiIn3fbDx2/Njt9KwH616vRQV
urxrfsgIvxoKS9ou+4l+v6uAwCiwn2tFwZMNCL3h5z6sj8hL0AxvALBKzeRUBxXC
EhnaFlVlawBcw51Dnb6LG8ARKKImN7Sw0pGRG+2CtcQe8JlgHO2qt/s6Nz9Xp5JD
OHsTXzOYtfStEIy3Nt/seAil31C6lVEpQCJA0aff0A+5X9x6f1KAf2MT1bPDJPHS
VDH/kWCORaOPhHEHUnJy/dH3Dvg/YDKhwmwE/rFt6AEE28aWoTnH/D11l0/hoFUb
D70/Wn3+BZInJCKXA++TL+Zf1uBRP2vY5IfdZJuKbsYNh5h1ZL1xwFN81iSpN4YF
zYcapvCNzcPZotHdUB8401YdpbNCSrm4ZBCfiEHtofvxIAijw/ol4euIVYXnJoyr
co3QbnI08dZq2qXNRepl7WwBGCQxY365Bn4IDeDYjxJd0X/9nTGVincwEFex0L3L
/f8ldsLRoccqgCwTw1i2SobccJOq7a5wDy7WuNuKgwNUgzg9oMXWOsajzDQR2Pot
VXtig0JNp15kMQev0UnZ++bKrV2BaQElZ97dNTQdHlFgkOThmpfJ7jHC3mWYRK77
0+N4oEskm+9z+uCYZmy9gNFOCUpthDpRF9LTqQ2P4Gjtbcos+Eu6htaoJ6+GHi2G
a7mi1OOTlWfb6x0iWYkMp0c1+4cQ6U/7hdZTMV8taaSnBKSB94zmoNRLr5XsmWHz
DaFWpP1VMGyzDf3tBkzkbOD5re3Bq3eV3rAWfWgV7HFky8Vg72zjSP7MIcyZtQ0k
D2kA/iPXdDy0wC7mI3FjaRJwiIbFxE0E3cXPXLR+hmxQdtgrsAgjsraFxK48uZQn
NK6OMMDSeLltSY0ukqHMDjWhUngYuMyzJce/U2u0EfhedJ08AKpDX4hA62LFPIXi
0Q3mb76qdf7M109aWiuz3T14/WpgGODVT5KDJiGr6zgf9T5huhYqZ6VXaHCPA20Q
chBC2vW0pCc6GYpv49XgKYTXSvsA4LtO9QVNB0w9toeB1dFH+itg9o3mMa0eL3ld
YZbqJhtPQhWjZyolcbS/5gRGE3FrLTsoQAiq+hRhAO4d++pbLSFMObu+G2gAcLk2
EDxR8AittQoz99QK0cfF5u36tYvsbtoCuEYurDoQgrd1XcQ50Rzd6n0Lu/eMfOtq
uSVCHBhzsLtNkszmmHaMba4EdLtW76WsKshrS3lf7fOFNKrNeIjXZSHr78j9h7cz
hTk4VD4S3cpW6CkTDreXjBupZFRW6BL29x20in3pNU5CuaXvyPQXVYEIB/wI0kPK
VQvBV5VjuH7tgmauZzn1dpXL/4naF1JwKIS3W2O17IdwULvpdVpkkFtPydIBep+I
GhP2zpOE/yGmekIbrTmPdoC0OfuflkuOI1y1NoYerISkaCzjD93qInVp0GfFvy8B
aHGgFU/Qpfca3LyKi2CXJDo6J/y2h/uwzx6OiN7tPceFye1NZAyRhtlPJwl/bXoo
vm8WEVPsasAdPGth/1NHS8iYVwSW/bY22Rwxq6NqBl0DnR4NNVUEh/KRLoaT+TYA
ricAcTIpJA/474KtawtXEAfSivpFy8My4G7JtFT6wzhzWR1C/pcfGtTYGzjmPTrJ
3/d8Osz7HYJXcQTxaImHVjAOuielyMYi13FdY6jqa4z/CYw7TExLc7yrNd8hYl12
ueFornrH49ZZkKUw2ZxwQ7RRfM1boJ4QLPIBzgRZt2SWTlC0BIdS+sOoMneIXvMa
3Jrk9PX4EAGCBouFkHcdgW8glA4l295I951N/XTKOCCcLaNCnMtIXg2h2QfHHU6e
3T52oMrIqZ0eIVrcmyeeOAy8qCfySNdw2GwGM40dZ8s8BYfucYN3MAYKCBHtYd5H
kMfquu3qlnPbwXUi108HzcwQsAA3o1LD29JdCMotdJca6gXmMcUfwc22DZsEv+S4
P92Dxd/uCLTn25gSA8qAfGomQHQ/i7tmdtKP8xHMFsPwp7/yprBYdUHGqwL4KdbN
0xZrSTZPySu1x9QXCQH+OdPaD1aMEMbANF5Fw0QeW3WDPM6WlpieKIQpIQZY7HGl
T+FBd4j/9yUkzxQftFVscVKa8qjNm4UzOHl3hXfO3dl+xtFbefsvJVEo9DXTcZMk
kqCOPrcb1zrqNvp+/+to4RB/iZngjKWvO6J/dhXP+7A3m2dqPBLp0r2f7Cal/9o3
Tq8uGtimq4kaLSvVmL67KXVu8BkUualVHyIXsHqDy9XFpMiKWVlz312VJI2EiLpj
fgfuMZZ8Uyoyza4vyF6RkOVaU8hYnXFduf3jqU8t4ueh6s+WQ9cnwlpH6gCqzgsU
iBtteyrWZfGBLU4SNDxofX7qnP44rr6YP6Fe9l91jxkS+qoZ8yInUa5OO4KObGwd
hanp7wuWAQlajkCzGAgOxyCdQCed+maITigMmRhWgY3RMratkIKcglCrUePFLMyw
gwKwZHOx1P6MmZZWEJCb/7Ipso+OTti7BC0BpEWPx1/bd5005P0gQGEzN6UG65xk
3o1Ky3XKtQuuboyhyb+WzepRE9dteKhZEZ0fpPtlH7gQl288yuEy22q2suSOyAwh
b9rgyOmioK4PD10SRbpnhtLU6NNZI1QdJFL4PhM5WivuS3NF5MyUYktBE1xA0zHa
G8hMuIuT9a4FKh6Xn8fL5zoFDSkBxt3Zs4NLxdFmBzqav/SFQ4uurMROlJeG600p
wiGRAMAabR6kp+jSPpuRQ9NRHU8lQf0JR+K3ReYap90GyaBrkmShG7ZxodkCEKjt
cey1E+dwi10F3MgGPrUOvB2qJuDU854kkv7yQNMoAr9RNzZ4MpYu8HpHVakhd329
hC9XFFvV92bJ/1V3S4vspC86/rKMbjIccrRN41A6/MvNTL7W5PImpIZtoFYcxuZS
UwHzWO7+B42qfspbU6HBLU+/P2q0QvFT7jCz8UnqOyhRw0rX6RAeBksy61TGt3lB
yhyqmK5evIpx1PFqTyhNogPa9Jxg8jiH5m/ZZA7kea1Hsw+kl+uBTvq3iDm0dgxA
NlSwVqt0GUydRNXplZyocV0vGS9bebibPreqm8GuRfLifqdnoBH5Xg4nWusuHyjL
eGTEXsPY3NZ/Vr6ceFTSDEaKOL/P8W6TguD/bfz1g6k5+x6MKkqsbS7OSlF0545/
k6FcR5u2xro6cyIz3ASa64FlP224GHTnTEYvJAAxwtpDP7jsAx+YQ0zIg9gv85Z9
GH6odTwxRvlrD1MHvUiMZtNGsHQc3sCO2BsR7O1Yo6VUdAJN3v8aKms1F5PYARnN
86kJvsmfhOo+aUzappaFIOy26oCdYsZr5xOqfgYTpcvZXR4Q77t1UVHIP+UUMpLD
AcIRxkKeLKXvMQ+b5JO9QXH50xKSSB+QrtKWcp5O994Y6LxKL1KMDm0nRpryMzr3
r4HG1oEtvRyv2WwuXMItRuVEEn+1yHmd644uQt0Ihhn0TP/howUKHBAA/bYpTCCZ
VspgpV8zA6374KMCAXqLbQwcrhaVnIz5XPBJEuOksLvWQLxM3fMApJ/iG2mVOPTR
+Vt0uiWJfkKvxoUiSnKz217SHcn8WONl9FISviKrEXI4HYMsTUCg4eS2pHqnGeLR
3oiCIlTiKp+lnjfg/2sDXz70pmWkFdeLnF5JF1lQ1h0FCZVSotdzG4v2Bflo5/0s
SMJEBF3ep2cD+e48atyG5I+f0tvxekgc0E28UAgVrfx2wnKhwf49/gZdmKykhW/Q
DgVMG2aoNJNRIETRudvyMB7kr5ixX/fJSDcL4ZueZBhpVclbPAW72WGH27tNScGW
Ik+g1kelmZGYi5dgu3hu0uc2uQ9K2liMJ9RE5Pns1ofFLMukzcuJlxaoECWS9vNF
4lV5x7m2eopVn/dlRyB4eBOz2vzT5Zj6Q/MozgqQh9KKDjFm5Nq6v0WSZ9pc+SKk
+cmcm38O48YrC2Qks4ftRXeDWy1Tr596pu/XyaiiiOX5R6qe5M1kDVuecJWTQWq/
j/m1N4SVUy5a/xUHt7RjlLRUsavYQ5zLjFzm5QXlRByGv8WCOO7nAqgyu/gVDMaA
2aZxsN6RPvpzkvlFOmx7M0+O4XTt+Ui6lkuXY69NUCLzUGKFQSmbiyKwIzUrLi2S
l3SB8q65JgeKJZBB5uRa2a5wCyA7UQJ0lQpdQPSl8It1PVwbBFx1klTZ9zXQoONo
PC5iZ2DjYugbnh6VFdO0x4Mpe8tYJH7PrLXQLGRyErCpejurFn2R4DlLkpawTete
sVS78FswmyfJ5QGvAGuElQYi6yfTMFeQL2+YS04hrAGyA4IZTrtZ3bNBwHQGIIr0
b8mxm+OoVNnIvJNHHqrfzN3Koyv+5T03n3ZHbMPmkHwgWDNOrOhTWG0oboxbj0j9
OcBNkEVk/pE+o5IyLXoheranx+Z1ne0YRqeKXH+y8UwAl5D7UXfqrqfq0OqvOHHZ
WKbS6oqF6eZIspVxv3cZvK0mwa7+euHJxxhYgZYRMsdcb/Aoyr47CYi6ng7N82LY
AGFBpzwMjsjCjg1eLPc0byCnGl18MljlmmypLZEe8Ju/qzOmAv9XDpNis5gVfu+F
dQddeNTAxUolcWmhV/Rv6HSAPGt/IQgezzcvx6EpJgN7snS7oSdj9DSp8CjG1289
ZpmjHRjpIie8aqDjJ33VETYvmmH2sJiQnrQUDGDYqNOnGGPXjQHXdMxPlRsyICSX
y/Td9mK6CCIrAQvqHVXSNjSFivuKzMvq9go2NBpgLs+26penGPTRG756y4WRZO96
2DsMqPW1Nzco4yFR2irUaA9wMe8FIpLjIk6hwEJ7GMgyB8VENoeIve2fDyOUke3t
cLi71jbSKVWx8rGLpXEwWgPv9HJIDMeGp843JPvR+EeB0QguO420olWUugk4jL3y
ZR5l/LtTUMe3gtHcI5rwGT37uNqNXQ+H98JHILQ4bUpMm5G1YjvXCjZTVq6htUJ6
EwkwGw5kvKNk0JB19I5dIOV0ES/ifPPsN0QpVsoM8PDG6jn6ZcD/Pjy65TuYmWTV
airKh7H/7weHz/k/A40NgZ/j73zwiVpyrFexHMHDBYYGAEbOPfcS3m7rSECQIwjT
1TkmNDc9akDhxFcV1sZEyrXZutwfyBjZk2Ci7qlQ+ksIK0CDRkA/eqO63Ap3bRln
uqxOJo+62xEMQVx47sOy/ysnKsP+N30DgajqwtjCSiNUNyt1sudgV0T2lrTkzAVq
TBjotljVAJFjAcvgWSgxfHaCX2OdMyFWkM1yhiwekMcqTg7MSdeqU+dGX9tnD1XY
+q9+bCOOpL1DJLDuWD91c5hzit1ILc4xr5P73JAP3SEZAL4IiJOMsKyLaG8s1cwb
COW+YiV7nDN1AL+qMdlkcmeK3lkprH9NF+pdtBJECppbGPs51wng1D1crgoybPWu
VCGnL6uzhtdeDTRdvUtKGWmbfhmOMyVbp7RJQFMcAgH0C619EdF2gwjXt4AuTAIZ
D5FUFUGmhDk7imBq+Lpcs9NrX4502NWSfJma27d4S+D4lFRS82Nl1pQMnnS1vBAn
H172nWsuh53Ox25u5wzYC4nlaSxsqtF7Winmnv+btMh0b8tPEPe+FGKZP5y+F0n6
fSrd2+qfLirdsdjruXfXAYHqZqOgbYdPRUK2KC23GadpMsTMW5qjtROMsGi7XgCl
RqqjlTU9RpJjJ981XFF64qZJw2VQbjzS/c9YC3ENdbFbb6uZPgBG3nrA2em2wmSe
vCVetUIqxF+oZ3wqWX2YpdZzsYYDd0eT2J49tKPI/L8uaxDzRv3YXKJOJXZjWVM/
sOv97DFtXgq8HbJT9OcyVH59j/7kNL5BHwlK0azS3NyEw8Dc276r9RvGsNgPlfdn
p5CDKYIR9ic0JAPNWyi1H80NJtaRwEk34jT8yobnWAUj9TfEFKiMrbVHEzuhH2Pd
EPiCVgehVLCit7/qGLgxiveo0ntgfVpJvcYXSKcoDSE4ouucATKMrlmz0j6q6umV
701TtR5JqQREpZrVlcC5JopHF250GOkAHBTRgjHRrglvee4oqpY+e/N/DxFPyW/Q
rE63OzyMGS0IUcTHksHvBk8Yzuge4jyHOcatTANnkEy8XpQ5Ml1qQUYf8ACVBoan
NevA0EZ+z/Bjsq4Tztd2J9xBT8XleH5vVWtiBPzKxCcfRj+6bNyB5Z//VJRq8S3f
IzlvFLMF2jC3x9F6WgIahMltdBt5MaH9HpXrIfvS8I57voC4JIcThs16TnKXEnb2
lQt4X/QqOZFwfnPXOYFDoJrQnfiEb17jBkKQo7wZXGLjcbQlyPQqQbpAy30XFy9S
pxellORgcPWDU5hyOGFBMuhS9chPAjCE6IkOYo7n2qqsT7/MvEiiseer1uRswQHX
q7YM570+NJrbuYIyA2Pcr5mbPX0pKQhECV2tYWUOJmFB46+vYe6z3oTYYP7Nq89w
rhVxEkDVOlyZ9DxJGKk1k0d7EjajY6iEleJ8z4HrG66Mm4aTOyvnq+IgQA1LWXs7
9nJXOn+VTANLTrsOU9QAizNZ0X0jTjqEZYjWMTZB5HEQkSvPFbfeHDUqiprxm388
dlhOscHsbqQ8xhUKYt4sPfClU1WNMnuaqz6ab5Z/qO7ePdM+5PH4uEkzHbSi1D+m
7vIi4iiBDDfijRu0ksBFN4hOKYKNsx5VvafBwFvVk+epiyRqrShUo/Rtg0iuVqgL
Pa4RhA3j3Ct/Th58iAV6yOXK1ApEA5AlWSsajjSKu0L7Hur9QHqVfK3CBLJ5GAfE
va34RF5Qw1kjuzPWgBM7h7ebrNHZiMwWIz5Evg1ELMqqq0LRwy2Xc2n5GwZcJBOe
dRgJSGPypndPvvCiJZ1+i92S3vfcSgk5DhudRUyKh1mcmdyy1By30vYyOB/fSNV+
e3c6gmudQ3ydH1NHGQOczFS/Bm/KcglZsHIfU/onJLJzqfAzIfcIsjMxrmlLzXiJ
Y65v3DIv6orXVDCz6vLV8ZY5YLXf+oKwo/KhFkHGfeXxhf6I2bpL0xO78Dr8qvJU
+XlyclhD3D6IRSad9R3bnsGjusUpavxAckn0tBwKlmuIhANdleXx3fRYyVuboVFR
8CoEn0DXFz8WQ2iZ546FlbruOpP0GpL9u5SQ9msIWCHCGc0HckO993fkokkndR6d
WPkBxK0uJHhZ8uuMB8vWznFO2w+A7go+ppeixh/BleWrOd5THIES8eCTn+ZwhAHv
MUMUvXPtl+ybYEVpf++lR2KcbzIK/MiNn3kKt6bCsoXquBtjmkydq5n/GUtvJoiJ
CXTndxHpy9+rqGG6ZMHPu5onv5fPY6eRxuLAzjowLt/ePZ43ZZWDi9dTECBAq5ef
NNTLTsrJocZbSc+NrLbsev/uQ1S/xgTCIw18FIQAk2HBvDBI4jMZCiXH517/r2nQ
qafwPMqi2GxImN027TSNY0YwKGAAl5/Blpn+bHfTc0KIZ1aXFXHaiPL4Z93OoOAx
KiKTL8Kx8M4QbRlfTOifWJHxAiJibc59gTynx7cOm6sjLWWFjLa66mm9xFVj6BeP
oOXHGJyiUUTXdsiuaMDdeXO+EGIczjZMTmYgeAgW62kYQeAYD+swT21n2nLH9OFU
Ql2DjewP3lHNEKGNz68y1YB+DG8En4WaqHW/HKOqzba25LooVjo2INCwMzILEVZO
EjQrF8RnyUJXH88MwtQZJ0TNYqxehHKI9OByGG/UWjcAM7riOvz626eSDP1Ufj2c
jyDNJZCyJftq2pOuAAJSVC0BavKoDds9uZSOtoMqiRgPGsYR5agVPbPrwvWD2QMU
Mb47XkbR9CTkxlQTCMJ3BAJbTMoHdsBUQWtK83njdpbuBBg+vnMVW01JPMflJKnC
ljyDhTsV+QcYstE4vbTymuKGmZwljZfR1jNkqbqDVQwPviAibkNBR0DORatV2dx2
3dTQo7R5k6ylRPIKmmPrwS33H+NCbYl3C26P09iWeXZ8Jjp0ZlkEuBDBRTEeMLlP
WKQ64lIIFv5cI7hWkzgGV5Nr9dmnyKUiGQOe4DDwOvgEwooEhEIs8fbDVSkcitEK
457gYMGPIa9oz6eVeSTbGJHCMe/7q+EKspjqUyn+ZAWbucphyAXyV0ThjHnqGn78
oUKqSxISJQY7ADHh4ToqCpp55ZrVJ53tlnL4cmrfnJd57oXu90EwxbczTFcPNvdR
e/YknTPw893qFEy9pcR6MRauJWCI5KHaGdPAZQTIPFqL4XGcBspFM+LO4qsMmtpb
wT7HaiPgjAuVqRLF1oqQwHK1gZq1AsG1KZ5hn019Ca8A7D7wSFlmHm80dkxflmY+
2rzjwVlMLLJLF5/LYXtYf8aBP0jio2JGMnY4hJq1aF7IH+rTcNdpIjTBCdjkgH8M
7tM0EkFI0y5nmXbj6Y6izlxEQ45JmvUtIWoWZoD6qunC232JySaCTZUrUB0rqkKx
kLc+J/6HQEgs6FCFrj2TNSnpEidwMYBwTHRPrWhWesuPfRRgo85WARyBq5j/YoaB
h7Op6RKfTSUbwZ8DI8aIK+yqOAH9MPO7CmDPmrPL/a9KDM62TpOvPxwFBG0WEqyb
H/bCYXRr8yoKCHOGzthwZuT3bGcrvagTr1d/hyGDckw47+q1IHfRIco87uta9BHc
f+YPp+UqPqqOzUZ5ftfbcraMosQ6uep8FPyu5vNE3WL1eIFOy1YJMpta+4TugO9o
DAZM+DF6ZbdxbDKCL5mEXYgF5yVxw6Fqx4Rz9NxmKwx09lGVSoswmgmCuFvAdjB/
0BV0nMqdYgZADUYF/cToCL+FYBdlO3HquJ4myP4sR5pRrLcj7JKDoGcJucJX1L7G
nytM8cC7b4kRUYSe1tEvErc9SYJ/1UQLynX7RBnRo4TI3WrXAMUL2swNX7NdTQ7s
NyByQTyi2FWXkLvMyMZW09tLGl2Ipt5QAbuRwlZIU2LqBCG5jCCY8OrcbZIZU/Dj
HkrvqqdPH84cH/ktoxyGlwAEDnclO/le7ulasvbgcNzd7glEMbhSdsjLLLqMc6IX
JpAi/rpTXjlMHbMPV80SIKWGWoVF3X9HrwsBQjTmkKRrVGZizlYINF3/CmqF8t6W
NtqAgbW1YBIEEGKTkI4lwZ07ZIvkpHiqQ3xr8keQTixpI283i8LUZRlWEMS2jBSI
yR3Grm6hEQm5yA7dsUR5Oh1JqLNvfkIEmG8dpodioPoPxNmVMSRSX4AUHyd4LNGe
LfHT0ABjEVDBZYX9KXZw4tn4T00X9PY2nRC+jYauIe14oHctR/GMaWhK5oUfNC31
VheFL24dSZOjv0NId2GbYE2SVshdc5FBuRoKEk9S7X+H2iLh06c4ca9lOwZP2cCF
jEOwURwAB1cBrEoiODmi3LBNlNmrqG57JCFXdaqq6IzeeIBVQptWDXEhgQnmyRiU
sNr2BP1CQsh+axkp80hjtB7tqZhN3vT6qpq5BhOecNIGKwWN+s+M2oo/s1Brm1Pp
6PTjN7egDm52FO2iqlWM1J8U/h12GBpQjcTL7Ost4AWyTapIrXEh8jN8LITYDnjT
DZ1cJAXqXvKHpDWNJPBFcDHU6bnzDGzzRNzrhCU/Ere2hVehogITuUrfgBIbTcJP
9/czQaYxjkZLnVDyj+1x/fpnKUHRWH/4T8roJv/VgxvL6sc/9n/BR/8Yer3ELZUZ
+VmRXcZHZKTmd2H9EdD/RfKsocRJeWbSW3GhtX/OWyKFo/K1YvZ3GTqSJkL+nhV+
y5K2rIhGDPEpMyoUO+q3EDBltqJm9Rs3Z+5f1HE5TeQLMfimAMADBkCAZcBFM6Vf
WSbqRjYJ6+zYXwEqEFdNjsuffaox1yGZqyO2M0HFfOLCrt4EVRiGLE5iaDFRpaT4
fOEKIiKqMdU8zV9YaG7Bw3pdLnmRIR/zUOkk16flPrtW736f7hBzPOSTWyXDZVRe
/PehK/attT1HZHFeekO65IgjYnhGbfVqFekfeaL5aV2oXrylwZLwNafhZoCXYK6r
NTnKukgtwUN+IWDByUG/5/5ReUhPDloRVoeKG8zTHELQCtm920T/ViaqgWN3riIP
393hvdokf3a6vmNNVQnEPFpQXVZCTQh+dVdFAzEs0kJYrP8gZ9RELerzU1IDhOpI
Vr8PXtBTVkWk5d5hap5oIRFnh5jXWNvFfPNGv3IlYzr5YLQcUdu6Sd8D2+IzZhzm
4xyEndLufvFzLyxpwxpPryoiy0EkErDukB5McPpAaU2wLqRvWuIVmytLc1DP6SuK
R1V+rded5Pzd6sk0PARcrTv0dy4L0Gj9l750/edsxhtHVhkOfR12rBsbMdVfQ1oX
3ufliMsCyukYhJs8VYEtAWaVzsNk6SSd/D6nJ2sa5S8xZTtVEVMmpDlU12/N/azB
zeDJtH9kvnR8mZMYqwj1px0fwa5VQmdE++prNuYwRbKmeBkTMiSDnuwhQ+m6rLdJ
ni9cjkhJ6Qd5e2bHDOExoZpLfWAXx4ThFECV6jJLbYWmX7f0+Y6TfRE/kTk0jfvZ
s6y9KG3lFq2MMaAiPhRY5h+W+sLVSwBo45dzN8B9JM3zZYbwQ0n9u7XpEzaB/0yg
GLs1ntFUD4+Lp9URHtUV21OpKMeOFofqVEhStKjia2zlSv3+r0IcLBbV6s5bfgRt
krRkqdzA1UmbHS16eBSSanSBx41X9gSTVvp83zbJBjPUmZ0x5vP+2lHFY0l6b88m
Dx/lUVtM8NA8JldiZHp6H2QwTki3GILiQ8U7cKIo6+4QYhoRsbiFeqDhtPsZWIV9
tC+gaZV0KtdLuke/d45RlPDXrTThrPw5FuHQWZssQELFCSZr8fOt8/2LV3oTc3rw
j5XNA3cx1Yam7u3PwXD59TyZUNZvFGbe0tuJKZ3e4Z/2wdT3OFHWpP3mo89Yw6Rw
HH1IfevkwblL8xcOEaro2BPJqwvsIDv2rV1OkA0Y1hu7H35boISTl/CJDlMjUl8h
zIF2NKuu4Rjd1vuDKGDZB/uIT/rH2JnqBpcj7AEJmGHPcesc8F8gpZB/8jLahCBK
EAQelOpDEy8G+Qz+8nsKUN85a/J6ccz+/l21ixABSZYjGJvae9dSX3gqSgV9zbWD
DeH/keROASRR2xum+Z43Zx7SIlobosOy5M+skreH644ND6J7X4VKsGlCTSEteUMq
YKre7wVLXawDx6Pa3uuqCOi6K2qezTxHre1Am9S/wxOwSyxbQ9u/LcxPsDxmCRve
YdVO99F+bLBrMXfkzmrc/MTKbMArexK2UbPvXXi+GrZwXVUhIdiakmgl41/eDG3Y
XmtQySyr2aX+on7Q+ILt3m3+sP6Tkwg+xuzKFqzqwhTqQtdTXMIkGVgRPkcGODkN
6A0o4vrqVTOuzwm9k7g9kq3JpLeqDWfdPhop1HV7arH1zKhSRXjhvN3/TgfBXEhf
sso5NkmnDjjvvRm7dVDjXvvIGTmPMo0bX0RuEa1tqvWw+iGJIWDefO/eRmM6o8a3
6tOVCQJQ1ho8X4nGcI4OBu9PtIocw0V4TdZOLH77xKyb2Hd2ptEbPYbb8Dplrb+T
4P+v5ZsIExiNsZQj8KvSdLkruCsAPo/xSaCfUuwzRCfzu+KWShV1C6OJVLag8Vzx
kit4xVydEAomJTr9VXsvzMYR2sClPDI4md2XHvLh9NkJfgKL0pGIJirn+j9cy6rj
QhpQno+qKpnLjRBtM8XnDtpsydoE5FKmxj5WbeuYoYGBQPFVlesWoWaXmDc34PME
/C1rLzJhxnQaaqPvSPGNIL/L/qAMTlhELDKd2x71OMuatqY8eTbCWQmYE0jS2DXV
tyqTPfZnjwh6r45ToNmh/HAPKOyGKRijOv0y5ep0bel/hRsgPrHyUHhRp0VzC/pg
QjwXWAHiM+x22fbnoGx/2x/FoeGU3U1FCjG5uRZ0POwO88RbJkG45HzmLWtDacAT
kMRdUlohxYjnbpzol9AYyxtmDbpvWXOxfj2OeQXxHdGNqlb1fkHNXvCN5dHS5DOn
NtXKKFN+n+Nk7GaaMKWtWHRbav1Bx0dimmz7kXqx6wdDrYN4hXBfKS4yCiJHkwr3
zNetgyvTBNmr1GybJh0lJ2KWu7YTrNORnRHVWiGhNJKR+NdEVuwINM+nkv3vyc3z
e0RRQkO7kiKAdJCMV+FGvUoeuMvCdsQaTvGHhBdznxiG84424yvI0n6yTVWjF4+Y
2Fo1MKWBeoKsU93oqTRda/NlX2fm6veuX4IZS9C4zz1+xB6cTgBErKVzOkwRC+0c
HjZEgfacdCGPdvIo6tITHvUgCM6USmCfdJYMyt9b8DtACH2CipeEIojOSzBhQ6Kz
+x9TRaEleoA+Wi41Mof/SVJMJbE02o0CEOuVk4xJm3Z9sciLoFx9SvAL7hohcXQF
rlfzqGF/BbpFOPkJWdrW3iWwQm1msdytdQwAr5qrIBegyNPc/CmoffmG5wWmeUD9
/MuD2mO8DBGyuh56o+1BP2sP9H2iy/9Lf3T5mrFszNKNFEin/TgQmHxTHv5j7FYA
6CpMy+idDcAdIbUz6vd4nVJuSt2zAItfA71YSavsxPwRA6KtyYBda4Sv3wDIKbAh
lLRkJffXU7iWPp9ZKTkMvmKwzMwrH+gxQlTJFaTE8JgH0muDT2lElWV17hBkOlFE
JW7tDodKN2n6OUVHZ80neL/nJk4LEADACM1AEUSXi6ggOY+1mc0QdXxGzd9NotDF
+qp3dm2TN2NVwBH09kLYYQkGKMQsaBvHOf+jmj2pKwZg/Kj5kZ5VM+FsXSDxCtfe
zLFK2UE7NxLLq9G94i3S5r81lO/6lcYNFtKTziZRumJQ+XvkGG7u2i8UbORZdLUv
Us3ciPum0Vc/bpUEoa3/PF+knPDAfgweymGeHuZnWLj2A35ludTHfEHuggijvrKn
Q/vR9ETw8EwyCrlnlQjd+jboM6UTzMs1g2VJVWg5p9biWjG7usu8gUWJv2Ovgpl9
kToBj7he4EKtu+eTjRxo32VlK6xzOGn3fHAJ90yN6urPt3kToVuhFGviyJu+TOgd
OKeZhWAXpPDMVcXlBD7Nz+advOZnTp6qLlwk8r2P9i1ROJ+arQ+gODA0S0NHneHS
hJiS/j6Fv2PEv3wqPLJkNJRr5C7tZAll9Zq226Af5IRL5Qi/fTznRkqdj5PV3ONK
O/g3fadlXL67Sl/6mITBjXzEziB5zfLXpnbPlOh0XCDMWjzYufORfezan0+NVFBP
wl0RSfrMWP7iNjcrp5C1OJ8PKJW3PIa0lZM6DjZKGRtfUjcq0/SErYh9Edm79WfA
A4wiL1/8Ai14RKWSs6w1P5DvVml7FF7kA3HOIhgyL0Hqpk2CI5vCA7FbVmNdjpJu
loVS0+J+kZzXO1tYUFjA6ZB3JkUogJul+FCDU3UZd+QoCoLJ6/a7lfdHuyCyWC5v
t5Gzl+m7ghakzIXPerPCNRbIX+yhdNLHWw0ZEFdGkLgErw4mrqQPgYiYRd3CBGMv
xFlvHhmNG8HBA/fv4Nl05t8eZ30+EJdaFqs1IbF9aJiAHExHvHe8B6XYcSgxk8Al
FCmvVYisEvPZIbCiLKga2K9LKH6vYLltsTafiqenH5elRt5SJS3a27DYP9aUQlhO
B3bCa9sw9g/Jf+xhAPtGE006nFVmQzYcbIYVvU/EcRuh2p5eEvMbuKfk9ok+YRkX
JwPYkTg0Z5juQeLCDEHMEVx7Q0W43x+GvbqOHR2uEHI3hupMxP3Gmk0HAANZmPdl
FshKXrBHWrMBTGKBmaPJj2HCA75Ref5ZYuZAIMCwR3bDKWPrRT7xi627dKgRYM5u
AHgsz/tuVguYZLHfLb64L6jlgzqTSpN4RJ4cEKok44LhtxCneJDFevQ3A33pnj3q
n23Ya639ivdjg1w9NulF08CQMSrINwgTjAbv4V/2sEZ3o7iQWxDeIw53lOjccKDi
sFcT+QBlUoCiDCZh7q8ydRBV8gXoa7Q2Qu187qLYCjHSF+MK0BwPdwHbRw9bQjXj
eXahDrqpMfLLJJr8y1YZjqxSJpv16rp334b56bGVoXOVeBM7e7btmgEvwpoTsPdx
+EHLftn9MPBaft6gyOKCTutKnnKjTZclbqQv+JispFAyaiGfKT3CC5/SVnnRUMYj
fnlkxnyjxO3Wg3A7kCgQB37w5ACBtmU5OvMIDLawxtBGma7xZJn/8oPUILLIdZCB
/Ck52YWvZtHTsend/eWyHYQAq25I/4WZXeADnQ7CBJvUpQM/km1jVmwZ4/ux6HDZ
f1fSMIDudvsM870YhQQtmYI48a2GsmCmccsaQPJrMWfqhnk5Yxke70uVgZC3ft7g
6UHB0GhJiS28wJCzN7RfgTuLkRcjx6K444K7MMy14eNUMRYS93COePH7bVx6t/bY
09bv6aO9GkRvO7B0d8i37G/SfLPIk0dsKw+iMZp5fCyfOcZKTg2gbHRIWc3Tu3jd
gGuKYWxObyWnb+lvFpmq73EVT/wbPKNQ7eSHN4UFToIK6EeTIry8OgdvzyNsyzIc
hp/e6qIzge3NYVZeV7DL5QUSACwAtqdm97r7ikho42L/vMZbULHDO4KY8cxW9v9K
eGDD5SQm23WDwgDROMvGmCuC2hmBhU48U08CWz0iGScE1ZqjpGL48EfEOlKh6AUC
3mYEtAEnoLNLcb9pT61DOMP/MHwanpx4d7+qAlKyxaE3mpIQyAT/x5LJIg8wDJvh
NpcVkgZS8ac5Fq9PmkaW7SMV4CNpRKSVWMVj09RCFBnZ/DcSVFRUcAStmA6wjmGb
6yLi4tKChbNfza6/YskoD10iyAl0I+vaDsBdoUwZ11AfjlqA0egkGzo6CfNL5PiQ
4Wfa6WMnu/4cJ8LgtLXVnzETP+VAEesYXs/bOOzoFu+BaBPG9kwtX0lUECx66jPB
8TVyJadvJgiuzPkwHHt4L6UDL1oeIAWDJOdAhW+MWj/oYHF287fd4RUnyxraBnAk
dL+HS2+go7RmpLpQHPVMeZR6YAF/GK0SnWBLAT+tftopSQITlnk42BZEeDh/U64L
W1SpmtcVU1EHq1XgnM3qxTmAe7omOSgWgKZSzlwNUheooVizK9dzAfFRVsD+v6/O
vgqSCkV9vJozyucVu0JTYg35LOAc/LI/qf85cs3ETFog8YT4yuVrsW1w6fSpm695
bZtqn+IMFdgieNjwMugfPBhgJXoOY5kJUXQ96TYtiTN3UlVJOkiXO2+jT8odRGKT
bsFWuCjVVVX2ldr0IZsZnbk5QYRvk/u2moyxUkxpo6GPU9WnIA4gjGdjM7NQFROR
HK8IvKF0nBkFZ5p2E1f5sQUZyxu5J3bmY6J1CU5mdupoooIp2t0i+I7FH6xX2yuW
aUA5c8eTPejZA77T3VQMfDvym2ElcbjpYkGuxMRv438fa5iAdYsx2ql+eGChNQNA
rLmYkMqcGS9oSD2ASSdMGIQhmu4UgHqbgyWT+F5heQ2K7eZPGlBmKfMyPqpLuQst
nw3vKnztkhzazVzwdGl86KsS/HSQOL2PzLPT+VSZInuUGncvn5ioOhWk+6f1CJAx
929PxuGU5tKcHTXTjC+f0DMVh4qGgMUi5KOHEMiAqEM47s8ULPilyuo7XHqdbov7
oX2X2YnnsfjqYswj4ZKY6SjJUb2bEVbNozPoGx/yKnRA3B43+HRjbKLtETIyV7hp
SOCvL3BnBDY2GXZu4pQEYvq80NsDcMNRwfE2MJfKU4NPyS/MWGwDXh+Q1fmUuvhS
ewvRpBEXiNt5mtHDpNPQ8JTEsjfy6XQVfF/pV2hVPxVeYFGliqB/XQwGPdNR4xKU
VOaMAC+AxFaUndF71/LpOT8uptMSCjG1OLBktEePQTD2KlsY79WTE5ppiAzXVtP+
sjiC/qQSatIZwGkPWGSPllQHbpcOCKzA2zaljxpXf7iTmNXmk5th+i/fkSelivfb
qW3yBCA4x1U+JaPiZ0MuDvnCQPm+gqZ4OqU2Ke9f5A72lCcIgiRKwesQOXN174wN
2uRzQe1wvM1/NV+mbQpodMRcUW9U8a9Ly9/wMJxtLfJZprsrX9nBdp7tjCTRuKRd
WI/EKlDJ0KZWrNEP1C2NpmVXH+Cx6SNHN10TxNZ/RjoIb01g/2eF8OHeBFfWXNGe
i8Vot/5e36/tnuGM8ykBIr4cw9VcAykrAUXyE16eIjOIV7t4h0EuuSb5mz813//Q
2mjFIRDl/D/7xk/IuaGq5GCx4XXwGZEeNeGfFwAcRqu2/ynvHrogeio7bWA9XoTF
X1D0U7i5W+Qc1Hs/iwjaddCnuwCyfi4MBC+6PPr1IsngTAoFAHa0otMe58QnuJsA
pL4lBMIFTcKT3BqN4y/Fx2AAh7eWAV8SoqNkI2ym37glaJAGoV2MVVhyQc/Yjw3M
qp788YT7TeMu4Z+JRvSqsOcTtK6+R0xvUQxe6N1qB13E06l02itkyvFqqj29oBOR
rBbq9e8dCg1LilBHam02nZ5SlvKIGkM66hZktfl6ahRCOlFUnoBckrbXt1Gbx0dz
cj1yfyczOOhXIADI4SagKuYCBK7G0GJV8WSQY1ssR7WDk2dSb74V2oucUZEgegpx
sGnyHqKbtSkPdorUWZaQlq0q0I3Y/+c4wd9PrqQMOobGKsd1iqEU20caIzB92kTS
NQqKOwPj6CB/9Rmo0PdHZyaIwIn9jaobjCLGrJv7MJHO5cPYyvt42O39A3CcLbdS
9+otZ4kXChNSJp8u5Srf9vntWj2kCjZS9TSm7aLYE3cEJnXqJaLH8ilUBvwjicZU
Wbl8KVOWoGa6Vy1MetjH95RKCQt9BTV59C/hSKjKaftjPvS5KJ3frjtvFD/K9Ppa
C7RReM3X0iRd/u3l3RipoxvUf7WsjDPO9r1OqcvG2frNG4B6x5AhKhgBRgVi32LF
vQPTDL0GzNZ8BhpYXlzMrKMYfKvHOkJ4/0a+KHiKpUMFby8rwnKAce4zBT6IIlbc
QumBquXA2cjWPhmjuYzF7BlaJe1ASodTKnENfTNXZ1x7+6DoMwD6hih9aSFKT3vy
KQFekKF0ReI+YMsx7FtrkyWmMY/Z9bWnp88Bm+Z2aVWG1cy6UBY6Vk20flWrkAff
nNbuehZUUquOLrt2S5dGD+5bizbclewwiszdVGwiXYuU4YqWR77lkEXPcwXQGKoa
vwUbwTsimdJC9JHVZSyAz/M+rSCaZ3pBYk1jqlVSfi0EpVFXfBEzk4BRFYYGBreF
4JMz7nf06n8pEzKurx+/AwG9rzfh4AsPWFZ1nxs2eel839ANiHzaxSXETtf8sVBh
ThA4Mt2cSi58We3c7zUTYUQrRV8Um4/p94CLPxcvpBASRqGScp1lzx9zpDKG7eZ2
FLYdbm5q+pyxpYKB0TQI8o80xhxHGWZw02S6LIVHHfybfixDS8Fzy7QaZj9A6prd
NaYzWBnMTKTK6ITj8Ohx3vZL6kba/v1wykJ0MUi2Ew2nEoPkGe/ooA4Y4/+RDrJG
NOfIp7uw1uFbBYplsyuFljhMsfwn8X23Jvy6SezC/l8d7KHA7BRynYcfhR/qrSUX
olpCE/i8BrJ9fzJ5XDr0fDnm5AZgwydOPyDDAv+y8UJizSr++Z8mOjrWXHYFSRtp
PcYAlUmi87YX2LueIJmWy2NmC5avz2sz0CV6DcCaAZhyIJAPK+HhFE9zk6JOe9Lf
KYhljRMDSvEbcecaqTi9casfashlXBlpVCMy0ZbsNJnVmyVDs6W82cWU0GzCA/DM
HrTAuYBMct/uIGLIIU+P9Ako8KDIVNctUKSXTAr/YtHlVWvFx59te7NFTEHCWqLQ
UOO5Td2GRVm8jdiPR7oU5db0sVARdObNYNuCiiNdKmmXsGXVY7i7wsYZQ2zN7cGl
5fSRCPSVFkdyVuhbO5oaZLLb8zgkOjHlnfdJgEVKlfBxKeQVjUJ6a2doy/Cwh5Zl
65mme62nRntY0jY9Fd/eiZN6YKOpqfkoSiCViPJczzS/1nCqPFFcYH3J2KaQTNDK
306N4BtIWMmX7s8I/9IbdMm3SA1k4aKhjXjHef9JPId8J/BbwB3b2uxDngSdN3Og
AXUvaMSNOMvqzvr5QifHkcndEg7V6OA8TRFdoK/BXkkdRikK/AEV+oOhaJDVDvYV
t67Ka9PRWu8py6t0ZW3wlQm6/BqMxA3aw8n8IGWGt8AT3gtEKcKdjrmVxWAbYZeL
MCdoGsPn7kg5mFseITpKbHUjR3GQUjfU5eGPAyhtweT7380jh7bJnJcZEJkwEXxE
jplVIEEqDrJZca5MepFdLe8brGBZvdPAz2sjsqgfqwnz6CUB8bDCCBZztYQkLM1K
W9owbYPLGE1CrdV60JEABROSnAJBQ/DXYazyNf4oxc+opw6LqPldMikUIhAyeQil
GZCUUL+h/U9JeUYg5Hy4b4bBmKdTRjtbCSFDUp8FTmYNHUX1972iTHbaXYMFRxG6
gOz0Dy/MxhgoDF68aw0Duf8hS9FJprtv+eCcdpn+3Hfqg+dYJ/fc4h0R6tkq0lPf
N1IjZEzU42khfdWlzxYoX/LVj5USlk3/0oZRJ0D2j4OGxpRiWCDyefDVBPTfqld8
lNLLURqBak6ZKQCNsi5SFo2qVo9qEGAm1eX6sL8J2GOPXBhpX9UsUhe0J8qtWD89
tvV1lg5BL/njxj+pqxnARkv/68vJukV3gZVTE7kOivIgcQEx3cZ1LFEplOmh4LoG
PnlBMGZ8/q98tWva3gOLCpp21EciXm4RrnTpL9G7JaysviNse0AAgdfu4d+VUTOp
nwFKB4Jio8jMGbs3/sx0CqCRPeAEkLOhed8tyj0cRlFYpIqGCXGI1AvFhPJrtYat
tuRA0c/a/mdimdoY5BKyuvxwEq+Jt05IilucIaWSR7zQ7njVR+Dw4ZVJdh/F0RK8
P8cQW4kiH0N/r+wFfFk4WZk2wxJgpik8jv6vguXj7hCZAt47/P24u6IclZuV+luS
Nk/pRHugPDA15bd7LN/GGkiZUFpPcEGqNCnZlYm5QHZDnAEV0CYocCg36njQQLzs
qfDvW4uwdyByRS5Y9aVteojWFqu8ivpYeSbTXEaVaL4QyR6gU+lMrA0xss4fIfhk
6S7oMAy18Edf8oF0eJfdlRDNajYEjTXaLXRn05T3mavtaYZXdhUE3yNdqiPnfJa8
9xWGCvsTqnTJjjGhJYQgzYrcIaS4R9JygtVMcIrXuP9eFjHh806xXiwyyVOarxX8
xGIdWcYjJeEMiRsDyf6Q8NpEe5V/m9ZhuzNo9womX+C0b/UNdfPKYXC79mPeaon6
Xqe7pKdJVdgw/kQxMxsWKwF/3v7uo72RftEO+xrlH0zY0FEAwHrFHItYGsOgtSi7
svrZh1w2uzoEL5mOvkCZ/VStQXwHaaCoN8QfHHE776v/33PPDvBEwtudV/z6h5XN
MGK9K58KCAYqDOCkJ3Ev10unexy2scVop8F/0g6e1VbYKi71hb/vbCWzk0LiqTFd
4JyV4++GmX/Ur3c1QVWc5fCenLwnsC14MsYHSeVn0JXvGjodFKZFXkRW9l0bs1Ad
Fo0HILWPNRkzq54EvfFaPeeTrfR6A/FHF1OWU4fH5bO97GZlcc8jyxLPmSHLiiel
xNiFF2UPlVh/3N8z+7cGDXD0h29p18dPkATGkAs2yEbYzWnqkHYVDHz1b6Gn5CMH
tLGJ4ZnzwL88Sj6nYK/kMmC0jPixzCjv1HKBTt9YYcKh5CZURYmthiarSNUoJCUO
6QS1Z5daWOFYqpDUTAk9Asdr5VvXcUjYTnhPDpb2NYe5NywZyr8uAkRIQAVCUiTj
MiN6AI8IUoGuEsmXa+BMu5C8KkjdM9LmeuVTgWX5zRs1QQHx5YTuKmJqlGJMXo9L
hjT9Kdz521fNmYFxhoLEQEhWfkU5KPaWxwnY29TLvQ7250exAFhhxvMv5Hphwjd/
L7LsPNkJsYTM9YLSwBPjwAIqbIIiJ2vkNg4mxM5FgCStfjoF/wN3uK27tCfoygDe
Sx/Wpp6kd6+J+VVIxWL9Ei68PlRGgMJuFSAG37EkVb2lR/nxQ7+3xFT0jpTbFjSs
MabQnBvUkWx2E6Fr63K1nwBozH414euLQlFiNLhJGJsLXuDci5mlC/3W6Y5oDnTj
OOCdVzgstOx1iH4ERRLNmqXED/1IM/AavJqm5hdM4nfwFLIj9GkdYIifY4UjZTSY
/26Vs1lk4HzUHIgGKQ+Ihsq/3jKv7Ix0eU02+g+aBq/V46tl7IfVTzfxrqIqtNeP
jQZNwkxCMuOqXnv/ckHCd66hO5e6PeTbVoZxLBhRYqSY9GArbnyooT6JA4EqtPmH
sgcj8wKVsZTe4fpOLlEAXhGOVIvY6tdXmKrL31W6kbr0Qflufq6013SU5f9vXWtc
EDsDIOONqq46p44FKRtbX2GV+9qftprwSZBCxS8dGO85XHu+fQNP+O9ZFqxJ3HM5
oCpFEGGYVpNkR61D9iEq/L1WZ3kWX1B3+qaU4q/4KQUtczN3Nc/67g/2QnhjG8DE
zv6D7z9Zdst4G+7B27ArvOvmBkTXM34JbZ84HVxkaovxe3Qx4FmN+IfxAl7Mc+WV
6lP0cbLclOxaRM8Pu82lbEOt6PwKXRoa9ujhPOjU8t9HY+liAzq40uKKEjvgzxDG
2yxs7jbW7/QpWA7xDEhgs9M0Va2G4iOB7K+LRjUPabw5KARqX5PMOTIISAHNXAs4
ZXgJ1rKURi08ep6OTKKqdMwKBP3YEenFM0ZIzRC8zbkUIXbZmR3oYQIz8Kb2hKYh
QY3bVVUkfUwzGqqSd5C+x7MWC4KLqE9piDL6dRJ54Z1YsDunZQdBw52k5rA4dZAQ
G3hNGsoIsLPZyugGcMFUa5BFq7/ZhG6SJc2cCFZuMJDhHNpl2TGF1xqeniBW81lU
ivfcH13oLQ7JXaGyliZEu+YSfsLfjsI6X2KruVMNqdonkUACb5TG7Gsaahh+7hUe
ABKp3HZecUvjKjWcxRGxNXOx218sBRJgzQqeScgTUBDoSHhYv26++daMSG+lzt9O
d58YFsglHu7BkbsiKKDCy3XSwopPWGsauHV/jDzA77SnlCbwCM2lbrZdVHni4Eje
+L4r4C58cbNtj/UB0x80VrI7ekabuoqw/ihHe3ElE04b+g2NuMVMp8T+vYbtwH0k
P13qNaB3enccyvDrDKkcr09XZ973mgO+4pd06CpJQ/OyjBqbN0yIlrcStgkMrGvW
n0Tz9DPJ5eSU3H6KLtFHXBB8f1zSPrNdrqh5Ln7hmxuLIEX2g+a/C9ovuTQzNRet
8LJb6PkaqObCqYoC8uuO2k6XtAfhKNIyYnjc+21k6+XkEBIAabyERloVbycq7Oll
DmyBnUNG49VzV02KmbCRB6yPjZSg/bbw6fOlEh7ZgdLkQrSEiaxUmbgGQPKPzYzP
63QQrtSWvih0YF25Fl+VmfQh+UI/Jpk+CXrWYxGLqp11M8s6+QDvAC+Yjlt7NOqt
DnGTYLKxxad2Mmo8x1GXuhA87cLkDEsF+AF8lcQBxVTO+g9SVui2wZyEjwPOe7ck
9djUWbd9qL6EyccTz+k69QRmxVAGixmjwKL/u5qOYgDKkt11PuIrkzCqZozXippw
juvtlhRkTu6RnA3+mt1oe/RCCXbcuNo5ftgTGx77+H38zeSIst+L2gDUaNu38uiT
JrMHlZg9BgKSFlLUnoDgq1OQCFZYTLAv5TBOMcSHV644rcV0uoJfCzHiRT8dN562
mgzOomBTU7ciMkqf5OjJblNxlfh+lRVGcHP1ukQPFfeo/MEzNqZMRAxwF+EjHIx3
EA6AJU72jmbd70tYA8EV19ihSYeWhzjgeTVD5lvVxjwvMzf3ogNadvIiHRpDFqHK
8WYy05gRJwLQ9Np7viYcaRgEej4P0QjXGu2T47kL1TGoMMxzOE0ktJJP3tqxpVIV
l4V4AEop5LMneGAotDdz7N5ORBItz7AFGDo52sdX2PwQjDS2KtgUlXV3f8OHJ7eT
Api35NKfWf9lZP9zlFifDH5PG2HHqyXD0eq3YcNL9Ykta68lQaYist1QVVSdXG6j
tpzsteInQEngepj5z40Qjvjn6zrOFD4mKz348Ylm/qCC+Jzu/pmUYVPGJEFnKsBO
NluKlDV/+bFtLW9XD3IGSPNJSYiSZ+xhYz9H22P7VivXwlJqz3GMPwCPpmgnkYXn
1eQWNqgLDcj8jv9pV9nOfmT41pXes364Ol6hz8947Z4WM1NVOyjCRRJdKkdXLh+w
nwWHDlzIE+gZn7sBMHoSsx1jZhPywgzDkiO/dnxMFUMvvJEdRnGTsDqDc5DIiMq9
aLC5LbFApdNDe/QGEvmsv4+ZDtsFVGjaIeCUqtMEvk7xeaGupNSQDajrk+Lwq26O
Df0BPiv6rpDklHb2N6NXnYXWsdgL6hYTysl6LX40AR+vLhpgJIFlI9c3bLG1CpWI
y5oA/qdxoezh2JGUTL3jNJqPopf/+q5HS6N+KUWumxm+6UirJHHBzKNiB/gbfUGN
oc/pTfzoAgQRS3ImW8c2FJ7sNieLyEn6mSZ3Zm614tv48l2DdVbFSg4UhpB/l6so
NZcoj4L3uLumR9lIIv001Eu9nWZCyAxZ/YxByafINj3Qa2E9/c0aa0akdarXP26z
0+YdBY0t3wRruxQ16l8lQaJSjy8lVcOBZoFXleIbYtGWNT0mLqicMN/b839waogV
7Szo+FTc5baRUxbkWYsTWzCkvQacb7t1Ol4Ks/AiqlmMpjigSXLGMAABeGOU0es6
zGP11YDgZVCxdHEDYQXLEl236fzIYP/ETnmfij+MSgHeEPDYJ7hdcEwNVDVeZDEk
A08FyOOQkm7+qjI4G5Z0IQJgjiegyE9EWNgpXjrOsHX55A3M/SlVPAX30NBxJvg4
BN8VWbtEPiOQB4zO4WiSKWYcsFamr9fu4yHekKjO8QUmRGVuyIZhnqA3d05JlwXy
C/DCFszhhkPomgPNc1C/qCL1We/3lP852WtNiJGNGL9LqF53Tg9GHqLCNuO2cUUl
mj/7/5LrtW0uFFUWmSGZDSfzu344+n8bildQQJiqatESBy8gLgmhHCKLW06ElJX6
oARPAHBVzL9ZPHnO9hgO9x7jQUSlSg4ZnjjzrBusi7vU4NgPfX9Wbcce6MP5plPP
3JZLdOefBzujrcktcFFdrvExVgQWZFShBbr1XOfw8fB0b1DH6zECtGINAm+SKPPU
M+Y0ZU0kVFd12FE7gToIoG9JIMUizI533mHX8upxNWo3J+FB45zjUE3Suc8Ya7CL
pSZEsz+OFDx/0DZhmQvjl1jh0eYvEo5BARkt1tgcLY5hi2+Vq+0kuM313xus82jA
T5zYVS6Sg9CBE/E/R8WdfBUhGUZ4e6fYiR9Cn5k4DWrU/ecS3cuu/RGPLUH669Sx
1gRxYOD/fHZbseVL54OKfTQ8bhB/bFLzdTJHWWGym7kbQEcMptsbpUtBT29TIpY7
itSvAAndZ8SdX8lJTpGPHDHcUxSf4E/LlEbwyll7XXSxQsQcVXfnCIsd1i9sMEzO
iIoggZrb8l42fkjcurRVIv5k3Vw1D9jMjQuOrRs4ElQ2ZlY7UkzfVAz8NT2+RcJO
YmWDY1Aq6VyOCTmc+Jw9OZsocaKlcgI+HXh7sBYxEsm3UnzxtlXWmxrQiQ/8ZZBP
40ryPVUlvaB6Jzjep1xYrIhaHWjd237mNq6Z6RPCT2nkqG3ENazFPW1YVEUd0fRr
rHTcHlJY4CbZUMRNLZ2EQCbpETIDlo9AkzyCM/7M8+8HJ8TS+Uk21fv/Sh+RXJAd
kdVpMrsBc72fpgqJGIJnxS8ZwXi2saV/qaKOR6aYOZpoUHV4m2dp7YxGDm4YK8CF
6zECjGLlB4ipK93WRM/wXREbXxZc4imnnvkxJGWug3kgcLNhXPBTyPSZ/Agfznkg
5jVueQoH1BB5v3NM5k9OJuk2kqXkiQqkr5tJ9nbVhacZw8c1FYmfvKPDZBio99i3
TC5K16UqaHtm4SYxcD6Pl0xrGcsNH02xoDD7/FQDgvQFlpqbwpm073oemVLHL80/
TGO7DQpb8MwE4DkX8Hc4YqRM9fHkblRPOe4jap2meWKXmNEuhWdmtFaCWSzo7B4s
RQNTygljuoYIKbwloRCL7pfso3QvNzYA663e5CZ3TIlxJ4/cKPq65RjgNfUbxGja
G401IEfyJIPV7XLUF3s8zGq6Zzq1jYbqyzi+ajqD+wpu60MbCEY9+w+Rr97K1q0M
MttJsu82tY5aONM7qj1ibCDZM2SYf6RTI/W/Xlu43+BvSmoQFojYFWH5YTkGbq1n
KV/V+SzuvXUbKvNsAoGHgm7JJKwpB3N3lrgd+yMZDdO1vQSL4dwfShxaNXUuvm9c
XYhwufVlqtJmzQ905n8KHd+PtnLVsybyogMWP4LbOBEi7SE96GLP00OIUG7SRINo
Oa9Rq61dtWfCNV29cX6eyYQRlFP88DLmLr3gVgqO+p3Doei4a9DHV/gQ+HvDq9tE
LzQdDL3P1ymB/XZ3shbqi5ntHEbT63ppRMQ2Osx8/lwW8hPs4nvAeM8KDbDENMgD
qmNLd3frtVsdg5kBc6wLR2lY3YLXX8n2JZ+H24ffMVsnbOgJ2xX/3hWsRFbmiUSI
+D/J/m6rDCATPFuhWL4F9ZO+5VSw+6geDGAJ+6gm03W/bp3QszeMFDsCmGY56Ms3
vQqhPS/bNF5m2jw75NKJN8Oe0vlMWwLb7+7fo+o+cb8kaXjfhcBOFj3AO4ymDCx/
cRO/hRcfphH5K6UKPfCnTuvdOKtCx03O+Q4Pzp3OW1dlTPDSHcuTegVHcWDGdx8O
E5juGQ8prCcidxzAFgj4Y3MAMlYuwwQ1js349Ec39Dk19SDJiLywf0UbiWz7KRTs
/Bi089IRHkN5VyqjO1eGkhZLyjF6pxHup9YbFR0EJevNY6VXmH8LAvx7pzzHwRUP
ZkqEgLI2+hbSuRN4p+RO1KtJAH9Oe2O4MWtSQm6VoZX+pea7cqn92dg22XbHWsMy
O1zszGBUuuFQcLi4/ho+jhkEFzMB6DnQfdgGVwYOZOLr9UcPU9eq3zEX6rPvKq7K
hjZnTER0n4TVmiCPV+cwu3mMnbrV9T6dEET29aau8mk43D9KdQlu/Ruytk+pnGkK
IGM94Y4FardyCUuSSFSKVuy1o52I+PuY5kf9oqkL+izt6t69q1H4sBTjgyAgp3e0
RJb3bf3s0Bvlrbk9fqETOl5+1gW/QxaXgZmwCDsK7CCpKKFm7AuxGicD+ajMTEvg
gx4TJHKyoXhKTrz1hepSBKFVziDsYAlsRKDk1mrZr2YDY/2vDLYnBfJNE6xu+ocI
9B4yr3vxCDd1V3hP1DqwBh5SdMmaJQ/BMcdvhdijf2Ad2dNiuHweji5kwYwf84iW
NvFUW7uLTLJ+OBazluNHn+0kp8WGTaDtW5eQodFCS40CzFWN322V+devcR+94DK7
7EZhz3MwJZC0BN550M6Pf3LRZwq1vZj9+p6KcJnJlIpfRO0g3bkG7MAVUoPKj1lW
ADprEwpbF5QiMAQx6QaH7RaEJNBHhm4nYBdIlDEzMknY4rygVkTOr4jwo9R625Nt
uctGm1LECs5qktojqhnaUms0URJ71HmUmpmuJ1Mo/AtJTXHBKcf/DeRgRjr4iBE4
677zhPRW1U++f1JVSWXj8MabpcE4BF6KpXp00kLO4B/WIRlJHcjWCzlijbZqFXxC
NIG+Y3hzBG4XMwjmtSe5iMFSyCbP0IsTCbtBGhmP+TqUwl/qmcB8cyP3QcRHW+j9
cNC/gd42Zm/Kn4UnSJiyHGlQALiqqjI3NDd8E+AvwPgyasppW+EB3wlqyjW/Pvar
1Qm5NyYdmToLcRypFkDuhrHxtCs6u3KTF3PI3quZ3olWgxka52LiTHrCHgGCd9Oe
M5kkIg8nyWwX9JLRXOzyJfdYDyeWVGkb+s/4jUTBTwuctVmmgyseHQf79ydf09V5
ZBCwKy9nU92fV0Bel0if3LKafOAtWMxm8GaAq31T30cSLCXFiI5LvkbFq6DAUg2b
iS3GNTJYyL3HdBcPyJFNf8f2Mam6mAxRJJBnSZ8YiGntpBuLVm4OwsIeMHwM1/LG
xVLlKdcAJAm87MbMPVw/x4WzfzSOzVCwjt2z82meKc8SoRLTHr4ZuSdhfFqy2ziY
0ESW7xVoo1ePi/+2aaHbveQlyaGAvdwT2j8/x16RUX339V3cCVS3TeYTfHnndmQj
O+qWlyS594QYzlQfaeIjAXZqdiS7Guzi31WxRXe49FXjKT0PTO9TrE2n1AnEoCcm
c/4MlK7I41VSLlN0cQVbCWJYHSzykeRwFONPjvW8soj05lZzevIKpRCSqmjCJVLk
b5+TC3rz9EyKzAcE76xaP8MC/pSSrfeNimB104aXHDCkXh8cpvHI7onj1te/Kqnk
hVBzOVpkkiixQcrLfSJs3NUohJXcn+LEkSKyOg68D1kNEX8aWfkDqgi18ZUI7mSn
nwZaYE6SP68bfHCFCrC/+R5No2lf7zr4K1qdKR7GSqCqUk5PP7unY93mqirdwv82
lUX8pYlBhFSGoLL0aT3MWU9ACCBvKd3as09YruTeqqOwOBjHnehsCixl/2HBfZjh
DK7/MXq8JXy9Z1HNAv8jSvBYPdr5IfiMog1SoEaCeTrNq9SMFaIRK4Il0/EpJ+3r
DmW74fLMiPlfKHWIQ8lN/MR6i/+ubfXcx0uaW5BR6aoGRn2R1QVMg9QbpaEA5/EN
er7ZBvi2aTlrPMU4mZKB4dc5n24PaOh1sW8eHSPV8APQ6dkDGDgLjI5aSvKHZf9u
syV/29N1QL6+nIP3Rcc2S0yDOqHz9ryF7UXf18zCHOFp3jUnMc7lYrOXVdNcrW+0
zlmrjCnJJbQ6uVax3IR9pYrinHkMzUlOv8X8834aYN4qtPzf8vPcFMbdm8aEcIRY
v+muI5VCKvcdYzRT/0T71p1QsD+OofYU3+2zKSkkhYlNdwf4kog4ec4bk03uoJ0q
EKuHSbn/w2L6sxlrSWmTUEXGTRcrop1J4el7dAMwTrrCNL/oHpOQ9q2DXW4y31/T
0o5dB6ssI588+4qgMu9eJUZ53Qq3rZb0BQYI2VT42VXwGpyXqnz46koKvlcOTlEB
V1iohJaIGYKnn3SVH/+/96Z0kVSCFCZ35gZPy0BQqKV7urFvAFLor34pb0o5Fj4E
ExZbm2yazc8i9WYwgCn5TOmAmdt4dOCAWJ3L6qG0/3UR8eXJB57nAVu4OIkUDaCU
iMrTnKaIH7D1DZQBjcYgEucCaBgwedhdl9NPa8hJtD+1INl9WhwcJdfKBc5xPYcN
Z+5QDwY7BHshHaJJ1vSpBFYzBQW/gr8xw5w4BAZZvgIb1gxAPmEKjBwj9x79Z1Xy
uKbhphjO8TOlldBRT1bC19Zvyo0cRy9fBRhZFlUD85wWhiXNZXMoYK+8zsZEmxJr
7C3HJSyRwsf1R3U3SDD/dy6ISuq7CKk9Cqbf5dLqtGf0VRdDCTv0WQ2idC3BHW0u
STDTLRnFnFbMUxunT176nIvOrnX5pIffeRFxeWw6Ah0Vw+04AAE7Th5xIYVcS+G4
XD1gpCgcshi5EJdIc5sketC5YAWOpyAKy4qaFRVxHyu1U1r/AcwNRqoUgjBtGOvu
SZKUqQGGipEeatQCAjMra3oOhAkjHmDUiMPzK16F3xuq3WrhChV35zJM7RnxEckF
YIlSoYMLj+bMH4l4TKh1VuJl7rwvACiDoiN4H1/xq6DqY7GG3IPf2gCVCbWTQZdt
m58xupgWLZ9a1RHx73snTahkWzrYUcXqh3LXsy2DLxmP0pAotYxljCShkTckcreH
m2Lz77v+19lShu2lqHxmcopIR6g8Ldy9RQHw1FUKDgXBe7lfZsI3z4WRcATP52Ex
RrYTHgyZYruq4asdbutI2Vx95I45fWmkSxnXX7iF9IF0kIiSLq+IBv0k59VpHmgq
n2XPyrNeq6s0ck+GzxC3qIByRVsYNo3XXw3ERwPQJKkGFLLKFSRq9VMG1SgS617n
A32XRsWiI3k1bY2Mmoea6dZDHGLtyyEN6EMHORiYkEnSManxoUT7PgMJPpzUM6sw
mQQdfujfN00Wp9I7nLuqtAlteqRZnWfw47U3vsxSEvqwjBfve2OAna7Znw7d8CbF
pe1PNxKdwGljUKWshF1sJwy0y6iWrVUpYrdhTymmx4VprCDuCfTMleekUcMDM5ce
8BRD07QGX44230yZFu7rb7V/rOabqKTX3sWJ++MADqWw1x1iRFH6YWDwuRizaJXg
DN8xYYBBrhLzfwqv0JDiWHAfsHtZNzHphdyP8D+/E0EBPuoIoGkVAajt1BZw3rZK
kK0rH50blXVL3zpPNJ9nHjDZ9/ZwlLrgVHelV4xBvWKPoUs3pQoh0PmBndLKLek4
ASyyRPMinl7L3GEcToeCvx37P/AGGxzdMKMmwvqFlkNHWomeh2iTEAeBTF0VgNXa
U6V5QSbcBliVlRLdvJ7k4raH1tzz3+D7ug7YrgQ/h/W4TUcR0KsKW0c0FqFvMyqk
lTe3AlFlwFtOEH9dn13iL9yZlN9GXVhqnYiaV9vp8UXsOsHRysYMWI/ip/ZCy0Xf
fWOiKXlGO2lT4wvxWuNQkL6Ym/tG8D4zDtl3ZiU6mPAzXxoHDvP/s+BN4auFHJJa
alSX1RrWraeChDOVYN0ATAaCW3fn+/2/JgX7pKgvGCxclTSJa1u+BxBLTzlUIl9Q
236uiFwhWPqd1buHJSMq6hJTGrfkvtewMoCt2Wp9jQC/pNOg8tVPj9knOGbYV7tN
SvkyA/8Go8Yl6RG7/NWrk3uDzzjwfyoRCOBxllWMVYcP4lEzUUUyUA/ec14zNHwu
1U9tLhslE7715tf4r2YZ6VdQKvSQlzeX5Nz8FGtydXHtFc7OYja9MWga5DkrVlkF
vkkG1Dy73qkoqAw0czAhGya93pMpkaK28prhfebAkDVHSJxMKiCMj1HtPqeUzKSM
2/txSquL0XZ7mZPV1g00Oj4RPi+m5GqHwS4+ZGECOcG9Op9w9teHbeuBlQZRhSRO
clts+aKnmdwDXmznpi/T5b784uD1x7eao9DsrC102864kUklEp27+32XThMM0itp
zxcKbWlavOtSKAZ6gP6JNrGzGi8ryEkwnpQf+vS+o6ONzddgigX8AUJIn59wSBCu
mbuUk2S+XNrTRL/ZngSuc3iwMaUMlrwaO+br0Os+fZhO7fA4Nv7YPwaF8QF3VXI9
Sy3ZwffoHjkgP7LhLtvOb7mCxShi76aZA50KIJWJPcY5QZEtkGwOaVHLuVgBl9ez
4S+VbDSD7K4+WdksKMbNqZ88385tG4XmLeFKThSuG9RIg+VzuF2cXmUWrMzB/2pP
48IYpqo844HljvyMjmiBMjR/jt4UBlVUWBENM234zue9FCwK+4FUeLtZ411o6Fcy
So3UWG9wjVj+ESg6glR06VgQgaOSSaKQm5LdkgL5tGE0DtX31uK1QO/QqBatvJOY
jUOf/xepu27AZ4IMitV2+Fd3oVxj8cbv2LIljTT9Ejsp7dTvWpxGAZnHu5vx6Rbh
eHtmAoi8EZGPJJSWaCNveCd5imbSFm1DYG/Pnn0vJC0bYIGJi4S3ywtsiPSU5XDD
vaN7Cn+pYAj0MOev/IveI9/DpzSxZQScQeQCE6EezevaiBJgDV7SwVVkOchOR8jh
+6RCNsIZkxhme/a5leB8iMCNGXC9IdPQSdUwSei8jvY4y+SZV4egQu2zQ1jn4BOR
rWVywIg7aCQqMC0d25HJa3fz9l/jGSYcbuggZnOvz8vYH3wx43VmsIl6uRzekt6w
pSitvbOd8NgMgnwUuXgN1mSH0Gafvac7CMOofftDmGYg97cMMtqc4PwayVvl+Lxp
mOoHvNziuMiFllF+/U2/rH8xSddjJ2zjLG7ULgSz9AKisG1eOLpPc/x+a0lOd/PZ
27wmtBhiHKJx89EydpqIoQ6Sa3lEfxQCC/5Oqczli82noNKHni0lp1en/i1ZKKag
pmpVmObfGlTpBgs/is3JBneIkb92zNUenRzT3D9ahRS7YPOjIfq1qPujW0EAZjrn
BBQyr+YpSaICYVwjl8MmaYC7gAwRttmUeKlTZBtvnvkV6EWDQTOFOPLNfPvZKz5Y
x+wmGTeMtwhjLCFh5I6Jo2FXj+kyRaWzh+T2fwGOUImg3BrazdpS5ROKV63SLQyk
6xchwiS9CnJyhoelz8isaMcrM1aVRbKSlURS85vryZL5CoVt9nw/4dnTKKY3T45U
XflV+H654VnQ7gbkIVOc/3H9dWNRi+/GGNtRAW87QfFEop4DQ0KeRC5qBM2v2jkO
Fyf3TOoIzDs4kqSYeOrZy/ZEJBuZVMe+rNWAvw/+xWWh8Wv34eWZ5rPw3wu6KAY/
ADt2gqkZjqfQRq3br0r+v8AcrIMnc8YRoiQn5Y7ufpe2B9keEa33osQkJHKI0mxl
hBeIIFaG1hNUxXpiggY6d69TDj5Q2uNdtu6LBSoimPmyECatAJUdAZvkFreWai+p
CdqZoSHmsBqfXE2Nub2qukOWL4x/KPr2ZK/MPwdTifOSKKHoF013IqmRrUbkeCXT
zbd6KM0Z+g7BIz+4UvJLJZttSTGAZ16JJSJdvTJLAJOJ/3fykI/5w04y5+/tkU7H
oHB9HRFSFnnHcweo7JmNI5p3sTRqpSL0V7u1x58I5YB5Ys5EAFAhovS2tJKHSjdU
gD0r4zTKd1ziOWc1bO6bq+em4ZFU6jh+hGshOao3HxiXfqnUzoonP1BFeDOVMq8M
Sl+yDTwvEk/qzPHO2mGnWjPiL1UrqO1yYuyj1LiveKMX+uEmxgayds+PVH9LETNC
RHI5wVgGtHhlVAF2dvLN3PiBMZ3ZwFvYHBBiu12Y/HAIGh2Z47Sb0OhcBrAnEeUH
WFIhNkbALfm6cy4AVE5wYsyYImOF54eo0qVKoiREdty5TrBBFROvpcng4W1hTysp
0MtrWC3ytFo6YKG5JkkOvC1o3hRBhnEYoLRSmxS+L5Q0+bcdbIJNBynYAagTpKMe
s/cNG6ZOneZPjjJnra7l6Gg7OYIb+0d3Fx5eMpahlDt1t/M+b/H5lG+kycmetnXe
rb9mmWSiNx0gh4uJ0K94UfYIA+Bmy+gnLgGCyMfHbZhsDfF/veQLDC9G5o0o7ahY
sP/9zN/Ym4JWiSJRuihJzzDBe/GL1JVix+QlCCeqdUWqO2YtPYw6otMHiNQ+LC/K
MxhVfn4XoXH2380hwUGx9La0xEL+Wb6/6tGZYquiP2lkZtLxy5aVNoBF3ogEQ1Ir
mLvXWYmaJnRaJvwOcY2M13p8snZBHiQt2QD+yTWFRBPlSKIxolAT2rmvpcEdLwoT
fgiFWFvP+SZ9/DlMEMsoFsBSPcCA/rdCxI6j5Xv92FFYLdPihCVUUALF+xFBgd7q
Aw4PsSB9Q2DMJL+9lnCTOwyZOwQ6jy1zfTi9IEXszCqr7hrleFMzofqTBHYFc7y9
h8OkxxRUl/5nXvF2UwMSOVuwPocccCXnKI7fNhy0PnU6cnSvylR7b+tZQwM8iptQ
wWmG6QiDZooKw2o/uDMCI5YnXNU6W8mPNyEznlA64qx75fmWoQBtiox0aKb9Escg
OrcUyOf0tlb9flsfrjTJU4nBCHi2xHQoZwnDdEZndIsmV16S1R64rs0ClXdpJsXf
x5NQRtknieA0+DS1UI7ngrhDL2B3J0HFqvdLS/Et+7fEhdPBUbGob48jj/Nirz7s
wOOGsWvHSt6N4fZn6lXXHZ3pVernsKgjpjxKkcb5p0y5ZrjIMDB8AerXsA//6r/A
mLtebE/uEMlik24VYH5QFpdB2BngHbm2oiamX4rK8vrdgRA1t1L/Y28ruOXNrQAr
9cqzFombZXQskcAF5kAqQfcyVEBxnv6nZPIwbpfVs/2azfH3e58xuVflFwI0XFzK
Q02zblIOW12qauzhv+AVWW70TDcgbi4R6m3NAIQVOONeWzOKSseVtM4+06QyrH7Z
2KX+OmVoD19mElRu0yXYZ6x+e8CdFvQiOLLyrQpWqZB1bbp0X2Nrz+jcpE8vK2x2
81SmH99lt6LWcubMPyZtfNU+5EMFn/uJEPkJxEzBedU0YlJJET3yaZPkm0V5+0cn
80vg3O0mCtwdk10/c3pFwwDpdC4o3uZ7XNagcA0PleZ/HVAxKRXRjMe6r/2XHu8l
iLYjKagwJkOLuPWTd1q0bSzOgCBY5Tf01Zrj8OhW6fFoLFdSbhjB3uN9owNq7VeX
3Iphg6MQzhFGyY4ruJh10ug0GKkrTP8h5O9j0I7w3EPRVZgSqQ8RrSFZh/P6ttPa
z8uffhA+EqmFrfKm9axbh7LxyqI/DQ15aiB1Kaf21cQo1d7ldIQnImsRY3ojfrTd
5mMTMQlPI37CJ8mjRDy+w8CZHASLVYy5ObgIY8/aurNi+p/3kuHWRFpe+qo/nPFM
1PedCFXUt93JGNGACL4fPQuOe+nTWdY1qD5p0g6wmA5q9U1gefhDm34lU0oK+K1u
2dOQ+a+UrmSToWHK7XJF9COLkWItFk+Dg8XgEOC+qye0WMMLLcmzR9ONr/dnYw9y
10DMI+8uyeoRdTSRlb6iitW1Ex+E/4f6TfH2T4JLcM3oXMojdDNMmGfuyNoMPve5
CwwKqMqvnncbmVlX4W6kQJ+W6Qt4vmqXzDJs7Z9xn0mh0fY/1y5a+1aRBjRQdsXy
gmtgfNY2NFI3mXpuKPm9UHbQkbxMjfbXAbJvePDAFxsPSaFgzLb+quBXGvvsfWYb
tlsvQIdqwuCgtVkLr1KqMncl2rQCYd3pk/z1YtfKWwyLtQiGZ0RDNyyQoHlA+KUO
ziZGUkuS0IYKLk2J6gRZsMxdng1Esrd/hK18hxk4/z+KYds1tN8/NYhe0BXNBB05
NoL7Ib3W1I+BeZpGKVbnMIM7+I1a2vFTM/bwmChM9isJyQYD35ThUnptTRzfvoeq
+5gdfBbP6Ug5o3OuxTXbpRBIfbyV8XG0CCDTNCtzIsgcFnC/4OJvc9WtQm6VDqvG
Z7RPIxlCAgLSzZ2TJVw930lbXxU15Tcb2zDLuDjDDk7PqB2ekTlOm4VLtZWJFCqN
UVlcg1kD4hn8k2o36yAMCB/NHr+OUt0gnjLaSG5xja+OLfPqLAJUMSOvj944xMiF
5oSDWzUaJ8609wYxZyfdIZ0DZ77muwitkvLs0i3iAUGCHhCnQclLgagPiNxK5LNe
Y02znuDe9PUZxlc/sxyHZdpTGuLA/RHcCCmZIiv18VeMj6MsXk2XIJMprbn+a13u
ykkwgwOuCT767Uq2qAxkCvPep32D9uUFe8EVTRdMr1RHRn71jeaAwppXZTcVgNpH
6mkYaEtrZ/b7HSkHtW0o4n9nfXcB59BGUjRgrl+Xu/WCD/mFLg5FB/fCfKMm81NU
agKMpP2LvP4RGD93UQd5barMOEub4a8hPTTXQCpM3CSp0i1GH6bu+dvpRMfVN/j7
KgVE4I3xMljy/1lOCRtJi3bnLqTNzAesyPptPs9ijKXp+0O4apz4kaqsecjKuSeV
l+7tAAzhkfS4uZluebMUWcZU0edSb/JOX8i9kXPvf0zXyeKlgfbjDVqo2scbG393
63OLkEo6rSjrVYtfMT6b6j7TgttM3z9iX8SEWZiQV/bzmFh4bT8ZCPb7US90yKKw
/pz2qbpBpFvvKtR1U26smjxIVuWUDhuz7WWfuxrg4tBKzVEQOnb17pmI8K9w5Tyt
aYK7ZifIAqw9vWtYqW3u+DOBPBIEpNTyRTMMO8zqj0yeDMcnn8T90HslsxgZ8St5
TLL5dqtH1m1TDtKfdHJC4yqp+N6YkC//Apa7YZ2sNwjALGmT7zS2NP+wL8nOJ0bJ
YqKsKAWuyeq8ztT/AsneBvpSDkxus3dIv3mp6PioxAbBoZTvrdNowURHxj1hDGqu
5SoPA1SOFTC5X1ldKC7GJw3uctmN4VYFi5MQ9nhClHT4sF2D2y5dwBuy3VREKEJL
IdjGU8c+NTO/ljQZcPV0nN8tJNMdPKsogZUpXj9vM/TrGJKmBsrp6GgPBTQEhkud
FutJ0Aan+nxoYtFxD480ZWokAPwLm/a28+KVcQ25vHgA0nrMT+rpzNvTbZwdWE4T
+cbK6UilNANht4xAGyggWQt1ACPFnmSbYrx3TwBSAaXW+9uiUza6SjDGZkGXAo3H
R6sgjV65mb9P6YaI4XBynW5oaaqOg91KeZ/KdE+sZinABqw1tRrxdhKkwmLndgk9
q94BFbg0tPrmdnZ9q2PWaZNZ87jcD9LAdmvV8pEbZSxGhVaR8C2oI982ZOPBgsoP
902P+57Z8adbYZuWkyjVdbFVWYH8RnSI2b0TCKfs7F4aevR2fGez5ec4TfUmXYvF
ZTFOHZDMDLIs6AR79mskNxtcTaHXoyLJcT+Xx31ucx1SXF+0cOp/4JBJaqJuBwpL
Q5TojDcNVlSuApj8q0mpgYV0LMRljQxT7x6q1vDHrfvVE197do+BPzbOo4lDOGu4
NsMJaQfZwFxsRD6oz9M7HcuqSrbVFcSvgdN3MwXU/52zYmzfYr+F2RrOqGDeGhh5
3YxYT4ham+6R/ZNyzrt/AYPX7Y3zzRXQrpwuk4VlmYTF8bsM4zijlWzxapISbSLn
XZeQjzsnS5JZsWmbUBu4YikuPCgUQY7wXXIJWVa5uME9fzgupTQ5kNGISQ7fTkWX
5m0VWDk8izSDMM8KT03JCcqOpzBROqP6AglioLV5YOG+aafh5zbr0/z1anBsalNc
MPEBFMiMEdn2ZWMNo3g60lSa0mulsD/nT51KZ+lQ1BIcYs4InbanuEOzO4ZFJB55
WH412SncrE0Rtdi0BmDyW9D6ksm1InYEvfVwDZYcgxYEo2S0Z7u7MrZ7kS2Pqk4F
BuM3E9/3helmJVoRuO/jNsdkwvPkReTOTrE+5cytkru8/qDzbUOi7Q+f7eBG+B3N
lU3busRPvKytgne1kCGMrfzexBCvMHVHQlEJ86uIi5c1g3G0H9r6h8UzUq2K2VJl
n9RdRbR15Gmd5i0ix8QqARU+4GuMZVILjRUuGMeCXxFoJdKP1x58L6D3MqpdZjd6
Pf2f+UQUPfBkfgt1djbk0yn5EFfq/jgHAchgvv/mWaNX0N6bbgsvb11LRhHxML2L
5WdGHWGU+xGeHwsqmfvdtOFsYcAKsfwtNqJUD7wg3BasUP1TsJqhXTYtaC8k9A0U
X+9Jo+syoWgADF4CTEv0Cp/jTte0auvcl3s/gvILEa46jTkrLzqdbsxaKUG9sRGC
GFqK7q7BaiAGbMjeu5PJc4TtNk2v9kNiWVEzlXeyBUechEF83I5hkkzz1gJxUSKm
+yyisTYPbtio5yhMXn3m5OPBkYsLskT7RsZsyg3492BtAjRet6Bvtrw1YyJSKHwv
eidYpHQSFjvUu/8lEWLJZ9fBTxpR4wrLfosYXjUJ5vSZk4s5iHuCsBANaFSQf2jl
Mb2nUtZKqNj1vdmR/ZtUtObECeZB+dSWVaYgXI8FLD6BPVjhlSL6CKtKn+SMwtag
LJyaX2c9dLdkfo906/GM/cE4LiMaVxADu4QOEI85PF5opnxN0jzIvoEQ80ZJaapD
+ARCvsdXgiqQrDgdWsjiwaeb5FGA27/tT8PzUq5OoSqR0XWo0xaguIlWPQCO9yjG
yYra1VPvn0SCfRKYm7Zpxfd/tEeb6qyF4F3z6M2YOZauwiwit2yMninsSq65tx0R
WMY1XZ31s3m84vaJ9b9e+B2zFMRLU0EcEi5McdGxTI1qmIWxYDB7PpCPmsERgLMh
PA3WSAidmpSHoAFIdz587HNtRh9751jSnyeQ/NVZ2Z6fijC3+drUSL1serN540RO
5GtMF6JvecnqCjx2Mtywlux2rMMh112JsY7Z8+hnqzkFwEuzHtISLotYHRrHf6mS
qLsKOm/xnY5EHc7RRy98UrYjXQ9mJjcU3ImJbNif0AbMqpnE1LpHGO1rhDtkQ0+/
OUV0RI5vGht/AqyRp1H2XkYwJW5Tk85fL4wY2dEbqYkBmDSD3Mxmj10iQgjcXlP0
ZnNwLFdfiNFsXv4C2Ww8ttEuqe0VOShWeW5UEUoDj26/ry/PMjV6DoestNPX1yHj
M0KKZ8QFlRXou7nuT+zfboPDgZ5zJM+JLJJrr9OrgLeipQNGAVH1wQelXs/8/mEm
k0ZW/ivUvk8qUiGEoEjugRW+JuXD85n6HCCo3v43HLtjzPMi2MzVKdTdYfAhgzdR
BCLTwCA0PtsZr+V96O5rOiTcg09ZCiLHkEE6bsJhBOvduzD+Ih9EZUU2B031aIsq
B0UQJJT+DpwoQf+2qrM7PO1MPRLoMSU1cugiGvVeRkjb7CxxREV/zVO9NcI8Km2g
106KT1qYr7F1jRedACO1jFB34l2lVNjmxHIfDeK++zxqHVAOJoUR//5/O5ffgUm0
pblWBqzBb/aEo0+MwSz8jt1+sR1m3dpTYWPoTldPmjupVg/VzLlK1z4wwdYnx3kH
GAjHH0GzooMBhuFQUVL+flsCpQioAPZtACxOG9P3ctbk/yTO4iAhazM+NNfA6JaQ
mMLoLwYK8oigxdVFL1ZtZk1hLlkkuWEAJ/wIUjqSzzVTtS6G3vVNQWJCfLznmuXJ
hksns/M6aDuZokbbQPGW7xlEodUp/Q/oLc8CFdTQpBjFZlYMJJ+l+kbaWFggO+QY
0xohsHYeuREgSZOI1T9MQKFxqvhxLSiMLneDckh/5AT8TJdGJifua6pTd6jT1lZl
o0kyMvpqD7mQj3TH3xk6hMPaskCE7BhV9DPg7WeTgE+YPiDEdzvcKJSO+Audj67E
Su51NdDvus0NgTh8s3wxRiiErJfZaWyrEcKKgumrEM9kPY7ctXSJ6nDWGCLgFAh/
9j9T5dqQRa8rTAl47R58N9BirT+1CWJmURPfPv3yfmHox/dipFcAU46SWYkYBsey
0XKCtI5kQN5Zpjl00FbvEkD7mkIv13lk5qXwB40d9yfhbssEyRYbCVYj3hanoDpv
phTcL7GdtuDtQkmYB3HRU61HoudkbzAWHobj4Uc2ktkrxOEijygI5WnmT1daJ9+i
uzkY6+ORGERggBZ0Oujfo5Wq3V0eOpF+X/3TK++KB0lMi6E01Cva6/obBtA6jhqq
38Uq42jlpPzKUNH81Y62nOJNo/s6/CgmyXva+lYR4j2wexZYus758wqubaB5CSGZ
wbCJ5By47F7jp+LUgz7KJkhSgvp0ZseKi7mwzsAANDPsnH0UN3fS8L+tvoAwdo4O
/qRXNSATMX55YnVTV7CXUvvcv8Pizhd68zuodd4VbIKEC1DB0YMTe4hgIFYEfXR6
2Kq2pIKWOvciMKAkohyQqU1q+TPq4JZmJw1H77rKg3Sc6ztj1ZyvIkTfInZhkU1x
4YcHRaHhN8xHQKyHjK/sXn4owBppxN8TyMk+HRMpTwAmg8BwdYGQYGI4F73jfRgJ
kevVeejtFcweNUnhQ2PzRVurbZ750o8zuhWxulWJPKcBFy9SF4kY37Yu9fHhvrwB
Z68ROQWPn4si/uPod0vPQsJGj52VB/kWyvmWXbDnxD8+G14aCzmTsSm/w6ePugLz
jUyg2FvMnQQkfZK9qGTK8XaNPMxIqlWLBI8XD5bS48VyC1vrI2VUiF28rfNl72yO
rfktMwM4oteCyTSFicWnzXRwdOKT1j1Y6pnELWlEEv4m/4VJby6XTTYM8lhLFBeQ
y8ASYZ66NO5zWlJxoFo6xsDTtIhi/ijYJ/VmPosPaEpSIhEc658VRefG5rNN7uqz
CNuvVwkDl98o1w0gmPjdcN1r2ZkjdONtBMC/wJbhmSo9tu3ATKPswmRCCs2wB5ri
HkTe290N9HWMZ1l9yn2BceHCQIb3xCrZJQDb2GHYnJrTbykxx8Oz4J0/bmbsC1CS
PeYtKj8Seqbn9NJd0jiII57YwxxEQ3g5iPE1SDQ2rF1yA4rUXmu9t2ViTjxnJVHa
/EER4e1bSJitAj+XXy4vu5XcJxjdbOhEGd8tSKbn+LQGrM+c5MHPn9+23U/MVQYo
tS8WmQ6LDHB7vSl9za2UedSocTTH5DjTmhvhv2KZs59Bq8OAlrgJBtyntGCz+YW5
rvYYYDU8E0SY0JvuuDB99415KUqmlmsIHr85DVFQ1xpzzRIL8iE9r4e+7ArkC1yD
4vmBm9I6xwu1blCzCr/0PvUtv3vSZLIL2wO4TPWfth6A1ss8ZD7t2GT09YD6y9bO
HrbP4Nf5bnzFvGmJYLzqHm2TqX++rnJDSk0voQI135ho7fPnBYo8rmFITFpES3Jw
ATCHrDsvcSxKALfHhYybrKqVNgQz1b93U9Vcx6zLbXYAEfNbpcviJyvoPxZy+cGB
c/euQQiG4h8DfaEx2elYGdpXc/SQHg0yyUN+s/xJO/dQdAB7Dty12856VbRlNdgo
ZuMqEejTWxSGziLsw/SuCdbDzSGRerniY6NYKVdIxaQQFb4lPJP8r9TGQwSvAi6w
3bci+4Kx8kazTkCr6lj+F8q0vUnZhDeyWVJTpjeBznS0Ko3lCOCHRog7JJxCT3Tb
+9jeM80mW1QTPXb1vYU+9bspdZmNrsQBGUrhnVszJisNEEljtC7dO0ds+Mm+thmx
doAeo60iS3mmEAAOiOjqqoUZs7l0H2U4n2bMyrx6W066HXdZjQ+6m/+XWKo+SpoP
2AXRZAI7FsMeii1OCDxkl4ay5mUwgulVWmvbEl8vpALQjmDhe6l5PCOSUejD42Od
1dRUGxLvfthugh/CyWW5mPvv2/2+4BAvnP3vieWvmY5JSqO8VlnN2ceiJfKB8+gg
Mps9EbmceF89vEViEAVtPm5GVJVOLPY6eIEZod2y4SLxJv0TsFbijfMD0E4cm9Kw
ZiJBaqUrh4QYm233EKocmxG9LW7m/V6ga2c3xIRvrH/zx+WJc+dCk0y/BZvv0V8g
`pragma protect end_protected
