��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}���B�an�gu�e�^ӹ�|d	�^�roD�3�c����.ݦ2nPWn���dU���bj������gr]��i��z��r�9JJe�(:��	�|�:��F�316�b�U���I,�u;�� �JB�#+t�\�	�������&X�*��zI��BDfBE�R�{,��B�}GW'��F(�n;�)�(�����Fq�SmX|�L.����#fІ7�!�P-��b����>�rG�<5d~��$K��!j ������}�W�'ZQ"3u�Mf����M3�8U���*5�*���W���F��_�b���X�~���}Qs�r�
����Bg������
��^P?�'~c_��'�W֌��w�
�z�����X�O�Q������b���/��D�6r20�$�V{cC�Y�u���)���F=�+R�a�m�}Ob�Gw�OX�G�9of�_K�o�e��D�Ln1�חnO_�����G�('�j�HwSfnJ�YhÒ��^������J�yNU`�KS��ܪM���VxM3C�(dE��68��J�x��F/�&��z�	�����;+U�`[D%3~M7��\[��`���� zf��'�T*v�ϒ��s��7�L�]$��1�t�b��7��~Fg[�|��3yD���?3P	m6n�=8y�z=z0�]*7lH��sEЙ�SS�]�3M,9��왜v8C-1
�������H~G9�ʇ~kmmse`4���)����9�I��@R��<B�Ěv�+����L@L��ܑK�)p�T���Y�#�T����F�M���3�2H%����;<��˛�R�K�K�=U��-�}~��w+��{A��#*E|��ִ���Ξ�����r�+��c��C^�ZΚ�@惋U�Q�d�t���y;�0�Խ��)�l}�NTk�P�Ft��--.�7>� �r�rB� �i�k��3�t�	����ꂙ�B^s�f}!��9L���1�b	L��d�qG�y����Ig�M}�:����p��j�W���PK"��5?!3z�Ƒ���V�q�1%!�/��,����(��?s��#�=���8��I)aD�X�S�[�ct1&���ݜ%���L>�c*=5�x�r����7K5ݟ������,�R'V����X+�<:͓�A�t��j�[95JFM�܁2|��>	�����P��rRNG�j��v{�,�bF,O"�Her�v�7��Z����*n�W[��6�d�]�Pw���0i�����gEĦrכ���G��K�
b��|�f��rJ���HE����KjY~��<��:~V��d����F��?c��
"å�JjFPI��Η9���}���w�$�@�bu����u��#�1!*"�� +��HeUu��vK[�q��RΘ�F�����K��yUh���Hk	O�#Ri������/�9c���Bbr�%ܽr�3z����°L{��5pJv�f�<����5��k[uK>�M �jX~�ُD)�Q+�ף~W�95�~,��n��A2G��L��m޳���K����==����XE��/O�4�����>e��Z�dd�;���O�#�D�	&�Zu�x=�8Z�+=сW1(Q�����ή��7Hd>��m���[Z\R�0ߋ�ډp�`)7ށL�*��\��4��2�X�p�I}[z/��Ri�	'@����?�8���$f���"�?w�I��r沛̏G��K���M��;���E��N���I�L�.y��x��ڊ*�d\���o�3�yBf�e~�5�����y���{��/��E�!�}��l�)��a$�m l]�O偨%%{I�.�K��fu9i+�g���������B�4&-Q�P��>�](j'g�7�[��ׂ��m|�Wƨ���ntY�D"�S�f�)�ւZ9W�)��Y	�j���	�eg�X	���n�0`��5W6�ZÁ���ʺ��˃�қ��z�5H�(�-��KU��Ws��6���,4��v�B����c5��KT<KII�}p����kSi7{nO� N�����F�'�m�#���LN�E���Îit5�\�8�z��8�a�m@P�yN���D�`	.�6>kH �lb?N1��#��M����à~c�Mg�죸���O�٫Χ⟘5çJ]�Q"��T�w�*���,Okȹ1���o&Q��ǏH{�ܔ������V[z��?����Oi[���$�VM����s��LB��L�3=�;�wsJ$�^V���1��~��d%�Ю�œX�\���}�s��֣�a��W,�W�<�>��K?�bU�G����i�ˠ��R��+7�IS��"��'WO%��[j��3�*��Ƅ�eJ}$V�c��}�ڈ�c���h�
�qs�����otK������K�e�4@��r#��5�u�7^#5͆b*�����?���b�_��k[���fs�N0;y�D�Clr�>}�+V���-��i�V�i*�Rf�oe��P�A��s�Mda����VQ�* b�3�C�Ę�T��Xrb��5���q-�"�v��Qs�M ȸs�fy�D�/?��
�Œ^p�铬V���i��(SR�7M�a��aG��K������XGT-j5�ހ��R�������{����Β|z�G���� ?6� �t9�ݙ:�zf;-�is�gt�%?+�W*�G��^��i���� l�50�o�P�1�]M�w)���ˈ�@er5>;VA!��d�p�t:ؼ1;�C���Bf����i�E/Hgߑu��-�!�>z��������V��f���%��c��LӅ���|�8����`�����M����L�se�6�����e��n+��
�y�s�;l����k�P�N9�e�]��V)���)4�%����&۬[�X���Wl�ʃ�AX�#uc�RS���O���VQ�s�����.�vԐ�vG��y-k��4�7:��?A�>�)�.D���#/��Vz$p~t�m��A�
XZ8e/R��~Ce������V��2�{��k\R�H��𾣄{��F�-�j�=*k"�0B�x~��d������E&�]�\3�F�~eu�˗pO���W�	bƬﲧI^d- ���{���ρk��	��Q��[���Ծ�����&J��ΠBf�H�hVx>��F"�֞f'��J���XF[���Q08v�����GKI����<�`�U_�P#-���=x�|?9v�z����/`r�� /~�`mܫ��!a���ٙ�>�����)F�8M�mB�,|A
����L���o~t�[�ūOT�kZW@IY����W�}?���q�zq�� t��;à�u�J�
���9jo�ֆ�A��0��_�g����B1���|���ѯt�H��9)bM$����B����.R��'$$#��	��+\��#�tCK�%���>H�8X�Y@��yb ����nS�9��`z���XC#''*!~���*k<M��;0,�^s�m��%��X�xK�׿6y� ��=���}Bښ���`lo�kk)�%9����<��-�Q�sP߭�)c����4[�|t�ᐙ���Xt?����&��=ה�&�lUlG<�5�(j}!%sQY+�1�3��5��GgJ��ynRpb��ڱKE��~�["q�\o�<�a�o�Z�Ip�!\��kVio[A�ɨh��(�.�z��F�'���K��h��zO����od��� OT�ђ)�
� Ы3��<�YY)M�_���O>�ߍ���e0���f �,�(�M�̶�G�Q�wN���ϯ;A�J��	��{E4$u2����$���'��@F�Koz?sc4g��bF���1�K�)W~��`UL���}���_@4Xo� }BY�wSMO��*�ۉ7�����n3Ȁ��"���g8~��y��bT7�H�cY}2* 9�R.�l���{+�I繤�0�_��F5l�;R��^�&!�j)o��Z��Ɂ�v0e ����^-î�"��Ji�<x7N���?[��f�BtEYT>d�)�GT�[ŹCd>�jZ����aA��n�Ԃ��F��n�595�w��'�� B`A�v�Ҹ#z���z�����Oxg�9sٕK�%��j?G��Ð�v훧3/���.�&�ěB��^d^A��$������(2���� |t;�æ{���޲圲�c�
d��B�RT�`�I���!TVa�q�$���F# �k��rBߊcĪ�myꣴ;	���%�Yks�-�g������3N��q�_\i���ַ���fҠ4�/��@��>oT�z��hE�>��L�n=�d��,�~%v�*1��6YȤ��ϣ�|:C��+���ݞ?���_T�%��W)���5DxG��G䡍�X�uow��x�ة��e;n�<q��]:l)�gN�B��6�H I���ȍ���~?j�Ǐ��J��|����~���eW�gH����{�#Kӑ_:����j�;6�x�xҟ@O�¦�YR�̡y&ڒn�� ��p������g�d!ڵˍ|���c<CNl��[Ȗ$�Ԭz��lM- ���9�@�E�F9r��~5ωe�Xٺ�|w�Y�i?Do� �� �?�8��\�A�)�~������Mb���x�6�X�7Y5���	�/(��D�X��hi��	J�@�#nƊ���`�̤'����!����b!D�I���9��)��*�����t\mS�vc�_�k%�.r�.�z�qzXY6ɀ��H<|,LW1����)4����T|��o��b��2�@8੕����R��$q����ϳ�p�`�K�� p^�Y�7d�Q�m=ʱbk˅ۖX�|��5� R�>=p��g�]J6
�Rb]ң�4��g��*㊴��i�OR�ڣ�����D��H6;��Șr���.��A����N�Q��x���Ԉ*K�3}�lbd�M7�+�P��Ƚ��H톑Kp!x�p^l�p�$qe�@z��.��"9�s>��U;��7n#������F�V!��4}	a���ԦOB�r��`S�VĪ |�G�t�yO}͡��H���!YM 5�9&�W��e�V9��O:��6��gHcb8x��PV~�J���s#���xt`gF�Q˗e6�_��,��D�I޷ɮ��l�Ь^*24c���,�������ӷ;��+��
u�WWE;�6��G:Zh�w[��9l���@A�x�'Qy_8��\2;���J��[�+��HO֥0�<��5<���֝�F�0F��X1�B89+ �!3����i���dI���b�p���Yq�6ܶ8U/�'$w�B������m���'7n�[QM+a��y��o�$r��l�vU#�ݾ�4���*3L���sƷ�~�e �2c�d��G�a(� ��TA�Փ�>���M�	�s��_4��������tʎx����aj�0,�+6Pr�����Kٷ���y�*u�����v �ʥ�]	m������N�d����Xa~A���`%i�ihQ��ö��.6u�c<U}}� ��+7�)b��v\i~��Ӆ�y�
��!��[��������`�����i�u1R���L5j��=}T��K��/�\:P�hIR/�=��#�&s���	��&�������|?��㣗ÔNC[���[�Lj$���qn\>�?�ď����y���bC����H��^��T�yH:6E��9/�=�BSC��)#���M�[�=.6kx\Q͔Z����|�s�~Q"�,r���	��o�Y��O�0>������K�'2�KDm�3�7�o�ݍ��?�Zw5}~=E�l�j&������%�B����U_Y����ϭ�P����pV��h�h��+z���I��&��x Yq�Nh�Y䄻�y��䣍H���4꼐�}��!��t��+}V!������ �>p���>�Mۻ��@oWb�"��6��(�d$J���B=$�9rN�S� �ߔ���ͬ35�0:�C29��DEݯ{��8i]W� �M3���iSZ7 (�H�אVT<o"测$ʫ����]!̜j=��ҭ;�Թ�&�Y��:2����'
vƜ��1P�p���K6��ti� �n�J������� ZƗ'��R�����ǝ��"�x��u���
�HK�n��.c��p/�Xanc��ʋ1�������eG)	`�\�Yf����.M`ĩG$7�?�)R�%**����1A�&�{�'J�qL��g]��[/�J�xg=mx��J�,y�$ZrVQ�ލ�� h�ˑ�h�*��ª��a�*=�Xi8�Jo٣j�Dٸ1&��l6_��-���X�燸�fsv�����|M�G�n�G��nD�m�ʲ�5�U�6��H��aVcw;L�z�g�i�J��R��HP�L�zY���AbC����1y(�c<
���aX�޵go�M�R����N��?y���`�X�9�������Ň*Ɍ �����ª�v�T���T\�sf��d�R�xZ�a �"��f��Z�S�&:��g��՘�~��R{[Q�^{�_B���oV�8Ee�Y��7�HU��X6#i��_��7��cu����^H�æ��w�:
�T5�z��'�SO7���/,�� ��b������N�/(4xl�Υ����E!ɷ~�D~ds�.�3Z�ih#-NF<(8����d~^T_1D�>�~�*1���
����A�b���CV�%R�Ff�[��$�ɪ�O2�=s�c��Gs���tB=��Z;g$Je� ��ú6� W�6�n�٤�������Q�m�'����1��֟V�5�j�&
4�u��$���<�F#X�~��_u��Gu�/!�����y������)�J'��H��h6g�Tt5��TR6�$qQ(��hѴ�6���XE��v�u'������\̫DL<�m]��c��-�شNGD�9*���X�T��]�'���9�������FL]��c�������;I���`6��89��B=�8��1ұ�)��f���dT^U��r��FI���|��t�����@H9�K��S���s����1y��q������1�F�������4��A�ꪪ|�FPw	��{��D`��z�y̶hr��fL��4��J�5QG?�po�k(����z�y`,�a��ȼ���Vi��	vY�5@�u7���o_�psG�P.n��&��\$�Y����gV�ڇ� y��^CZ���?Ht	���j��SH[��)1S�j�D8V8������?�.���Q��:Y4���V�;�.К�!���{�L�E�ѠԎ���,�l2�#
�Rsכ�)��כ�M@�`	�L��.+��,��O�Ek���(�懼�0���0�>Î�C���ZR#=�7#�?��)� �xQ��y��5������(�YIL/��^�4qJ!�P�,�G<���WT�(����G蕾�BC��V�gJ�{\L�eP�]��E�QF':�/ �fa�Xю7���d����t*z#h�}C�jm��v	k��K�T�F+��}��:��m��=�ԅ �L�]"���p9�����mI�u�̂��&;!���$� �5���D�i ���:+G8ME����3k�������޻ڼcżzW�p��Q���	)	��g�V��כ��DHc�^鋾���٩�s'f�*���Єg��m҆T���M�"�D��߼sx=�r���3x�+e~|�$�s3"���g��Kт��������[���q��l8��V	�t~Q��|?Z�NJ>\!+��A `>�MB��ذHЦ�%$�ą�����jt�@v=�J����,�M�zdD�ل�Z�z�����_�l	�v�I#[UB�;@pʲb��п�	��p�I5c	�ς�E����"��5<�`����ȧ���6�S�ESȭu Ҿ\	O��;9�m��|�>��5��|�VΜ\_ �������~�&�p���9!Q�� ^!�eͫY��c)�pp�nQ�@���^*��*�B\k��TIG=<gv�yb��ǁ�DZ߆����� �~p�HIܳh�mBG�K�9zb�p�X;�[�_�QnR�K��m��d���<����ū�"�Aqy���?:�x�����=eVw-D�}�6G��yZ<�v��kʌT��D�e� �i>�Ȇ��w+{z5z\@j묨�z<<A����Ȼ�I��h�W�k�׫��1_k�:wB��]ђ���c�,�1�N�Oj���O2c����#�ċB�`m�/7�����t�R{��\��6�Z'}����}�nR���_�!b�*Ӓ����)�C�/��_��4NP�C�6���X�I��"|m�T1�8�G(J�:�oG�+���M�UW�&��-���,.��A;0�-,�^��2�����=�n��O��æw±���:猪��w׮��9�0Ν�U{#�(P6�v8����g��%���:u;�b3/�*���62g�w�с{�n�AP��v{3�U���+����B�.w��t�!á��jۛ��[K6�o�D�c����+Ò�S�������;�\�� 0��,�@�/];�vٮ[1��!����+�����(������k��e�4�;���#k��To��:T:�a�Z/���BsF�	S�~n��f����K�o"ɔf�)0�G��FḳׯJP8��:L�bPH�!$�$F)�1>��B�5���2	[�ek3K�����_�0;��
�׷�r��LT5@L�ݣ�=�W-�$at���,�86�U"y�����Wp���M�#	�e��i�D�変ej�E��hCﲓkF��j=�)tc�����V��%p��X���GU�������J�}w
jun0�^i��M���J�d�[\��ꃡ<�3�e{���n+#.Հ�a ����/K�d'y�w�$J�Ih����<h���:]���,�g�\�r|���ʀ؎�tf�߇ܳ��z&z�o_�7B[���Ȼp�Z~J"�Go�l�#����W�m���$4��,':���]�UM������#��P�	E�%�N�k�CG��MPi�x7К�Ģ$*O9�0��J|���\}����\�L��L��ڻ�o�H6q�m�􇢬��Vj�c�$c5���.�Ƞ�����Y*-�-�.	"�j��G���J�[��#Q�`�/��}�>+��j�4vM��7�1XZ��L�;��7�hy��"�EO׻gRF��JL�`<�N�i<���V�p����E�Z�B�i�O35��2�����#w����m�T������l=�3ڐ��Ԍ�P��)i�[�EtX�B��0&9��*A5$X��������_"�e)����]&賫g�&�#.���R��������F�^m/>`Ix-��M*�b���Q$t�:��2?��j�W�i�������4��Z�m���RY�z��?ָ�+���~�� b'K�j����c���V�l�(�i���.ۻ��٧Kz\��pYߑ!9*��8�8��e����/˵d'/R㨆ĥ���H�Kܿ����b���[��)�LE�܌�)��*��1����#��q3v���%���dX���m�&��[Ὁ낞��@�r��v�Er�לj�[ �R3�ƣ|��^��"Q#A��#+)�ӎ"����3��h/�(��Ѷ�3]�R���'���{YĪ�d��Ch�E�6ߠهa�����QTZ>�{qħm���	QK�P1�ّ]W8I�"���M��]�J�
K�*�����7JM��p
Of�f0����#�Ꟈ*�>� ��^��3.Х�@W�k��5<�Q�^�4�3o[A�N�1��';��:$�n�z��pӻ�	��yc@�4w��� Y�#�.N�4��m���e�����������bH�b��_{��>�ǵ'	?k{GgE)���I6���L7V�v<�ˎD9�������F�6:�w��o�2 |�Cj�s�h��iA���"�i"���E��Q�����6�.uŁY�W?�mخe._ 5�R��9qa�&'����Z^�,�m�KF�ڻm[�l�֩x,��5b�Z�e�l�$q� Q���\��^�� �b�/F>m������-�ٳ�׺V���T	Dw3�-&��K9g�<��.�s%�\�GU�Q���vN�;Tc��:T�2�5q��*�F��QK-.ٲV�ԯ�V�X�KLQ�C�`%�Ek�kO�Ϳ��{ˊ�t����+���:H�@��C��of�.���\�8�n5�RC�!8*M�xiw�D�u��wȳ������p��X����H����� ��1�T�H_4 �G[���+���Xi���{7;��@72�ރ]D�_=�[�"�T��N]#����z��8ǺȐ�����tB�G�I�#�u%�����D)�a����&��u�	7���V�Ot⓬
A�P*�*���:�t���ט�W79]��6�Wl�M���և7p�\rU�\@�^��*�؟�J0gjmhmɺ�Mv���~�������$�B�t�z����%�ةkQ�oL]���<��q��dm-,K<L�y������h6�X�P�1�9+��/��D�ڦu'�j&�	�y0�`Y�%����K�S�����<���S�Yq]�����a�9>���h���*'J�+�� Xj�㩌bp����
O��k��m�Z�ǝf��J���e�ViZ)� }e]^�*��&=��/�@N�mk��e���`K�f�{��'����xx�ڬh�@�45��b���y��v���^gY�Қ�nF�+5��O���~��{�w,�m�9�%���Z������!|`�������f��nRO�A��E配k�Zd���
'[����a�]i�~�L����boT��� 5%@�pf�p�_> �a��m2���0�X����gG���b%P���FQ�p�:�zE�V��y�B֊v0�[�	;zpإ3�pM�k�nN�b��c����9�Z�P�f��FK�"]�r�R	]+f*Α?ɹ���~'kx��I�����CLX7��r�f!�Y1Rq酲���+�t�t B���\$�;B�hm����xR���P(ά-���)�YcҶә�iN�.ɬ����2���}�\';�mp�$�-MG�qP������J��K)p.��I���*���.��z,����9��G��Z�%z���
5��Z֪%#����PA}�e�l &�_S�ӣ�?��C� {��I;��rK?���	�|?���tP1	��� ]5I��B�q3���0X���ײ���EQ_�5��*�t�|On��^{PA�������X���q;1��u� 7p|�B���z�y�9s?*K:隶���;��_̽Ŋ�ܦ'B�k�#�V q]�cb�1���g��%����4*VF�4w=Wϭ�+���7|@``/�g��7�!�;�o�YF�)�	M��?�X������"Z��"D~���`	V�zm��r*��̰����K��D�!��E #|'Y��-���-�CΓ0�T�벑�!�C�%[3i�xgO���I��=OC��6�3IU}��jϸ�~��b\��[7��n	�����¶��I��씄h~��ۧi �.�lP<]b*�RoA��
����zS���A����Y~��im{_�����S��{e���?qĤ�_-د6PDR�a�ܥa�k��{�m�}Ӽ�����Q�yf��M���'���	n��v%�L�7{�y�L���Ҽ����b�ׇ�2_�976���.� ��^}-= ;j2Y���(
�-�����w�b�z��X�Y�stp����Cq�T��0�2�P��K��%@}LT�ߌZSNP�J$�)*��7���2դ�����_��.&S�<g>���3�A0�?py�J����}F�?J�@D.��w-�b�F\z8e� �2uD�f�X�N��+�K�ZI0�BS���&7Ky���bLoH>�a}&A�&�<�o����.�������|t����wC{�&tx� Ȱ���C�����ښ_~>�\���{(�")�͝ɇ�$yi�(�;G�{���_|q�������x��^c�cffȬ�G��<Ą�4��8��]��]���MQ=�������3���x]&{HЍ���4i���\�r�g������R����ėH�N��t,�2�{pe�:�WWc^��!.* l��b�)�I��A�*lTK��\v�^b�����c$1�V�Ѷ1Y���c�Oq)%�?��[�'����I��<0c��n��M�8G�K���ޠ� dr8W�@����Xr��)�6�ð�zt����|R�fhT-�'h����K���ڟ��_+�0�����6,}�
��(�Q�6a^�#�o�2ó��9�x*)�<lL"��ۤJ�����X����7�
�nQҼ)�8ˤ�0���Z�9����K��F�pcT�5Emeժ�x��.�
q[I��AvB��f�� ��ջNk�����J'���rA��W��Ņ��N��
��c�'욆���&?�p�i��)Y��һO��I0�G�N�n�#�O/�.���>F3�� ?ح����*���˄�6��,ߐ��4`G��2�� �eux�A}��$�x�v�����oDRay�`'Ho���M� ��\Wd��'_u4n��qݔ �7cokvBM���C�M�/�Y�v�flxX�x��H�8	<ʏ0�9:�r���G[Z�DN�����a��q�X�iրb�%���3��<@F�S���
θ��|�"콓�$�ȍ��2��L価����P�@�"v�D�A���d�:�+��'�O���o$�w��k��R�fX;H_<<��O�߁���-9��C�v����FT�(�j�:�t[�]�AŪ�O����wc���{�j���kf��>���:�x�KRX"�����AN(��8�ݵ�� a%o�%cRIeؕ)f���9&���Q�*���rU-���%��k��"{�@���~N��=��`E��Wn���0Ѽ�=�k<��`� ��ٟ���g�c��c������p]���P2��$�X �ɟWw�d�0�����ڔ�Evk�����G����Qd�t��'���n|߻�%D���`�Ǫ�u*e�%x�ZAf�\��q�G�r��pt��5�n��g���x4��(�����+3��ZY]<����h��{�j"9OZ7��P�;S�O���$��O�0ﻦD{���2D?�=9)BcҖ�$z�!�?15a]�U 2�EX�Z�ر����9
Y�N��= ����mSh�ֿfA��bP��
5 ��A
^Dbϕ�~�	x��m]�
^�\�
��:����N���H2�r.Q�Q	i����3$�W6V�D�e6�.U,�vR�$�w@d�~'�pGv�u�y�J���SK�T�d�$�[(���b*&����4�w!*��
A��AŌו���m\^4M��N2��#�B���4r�zJ
���u�ʤ��@Ņ<��uaC������P�䢮�9qU���8`�6Ws5h ݽ�=jODMȇ#�r
���q
�Y�{�.� D`���^b�������h�G������=b��/��""c��/U�����:���%�v��)�Q@�LzE#�\!B������S+��f��w�/TnTE��gϹ����hu����A@�_1Q�����5����� �s���n]xʈ�M����k��2��2muT{�q�.�P,��Q,N�7%�#Gi�T�1�\�!%� ����]x��{&���I�qZ��#���2��R�o�(�&v��A�����WrH�>w�����Jb�U��C�ݜ{�MG��vHp0vC������Ŏ�k��ܓ_�UR�#�P{z�P+[?^9�\c�81XqO���:w���Z��I�J�5w�d��]`.H(��8[Wu�\oF�r?׊8*��I����{W둘Q�]j��t��	ɳR
�E�tzI���r@^Xl6�8�w��w���Ih�$�ml��tX�������Z���*�"c�Pâ�[`��B��Q_�8�cЛO��	��ԑL�xw��]��]����H���H�|S��zhN��A�Oţ�)n�hX�i�UVw|%Ut�aȭ�0`�k�DM�U�1�wS-HV�z��Vr/q��`��w;�$�\y��m�^(�T��u�H��B�&e�u�L������(� ���	�_�wN^/�Ƽ8_�막�F�E:`��4�����@M��K@����*��@S|H�sm�����wtNW��}G��_sC-@Ob��G0��ss�t�@}�.�o��:S􌩯�W��A��-h�(!���	(p���2G�|�v�!�y���gG���Its�D3�/ʫ��^vv:jC��m�tZ�^��������8�e�/4~_C]"��е2��� FQ�m����t?pm�Iy�nr��[q8Z���N^�4��E�����"9&׮*E%7��l�x�E�tnq�AF��z6�|��䟃���Jv�-9Ε5;1J9�ƷiO"^ˌ#���L��$r
E*1 v\16�@�fR��M��}p�igW��h����J4Ǣ|08��u���1���*S�!2�����e��|TH�8�V�+�z��N��R���h-=6��{�uV��$�����}�;����;GNpJv̨yB�wzw�����Ky�pQ�K�{/�d m���W���)�k���"�v�	�E���᷺�|���;���d�d���q��^}�D^�>5�P��w���S�%��l?(����X���ǜǆ�H�?��^�`M�Ӌ6O)�bM��|K?����+�R�{�����hrYs��N# �x}n��$d�T�]�4^ 9ui�k�B����q�FxN��9����೾� ������jX�;�x�&�e��Z���k↾R���WЊ�skKiX��0���iS�w8
�T�1�M��\P��,�TB���8A4�o'�,��ٴ;Zy��k�\��h�i��A���\�8���jM��;"N6U	�j7"�CN��V|�'I���H)�:�`�� q#i4�[a�~���̪��C�6@�q��Jq�=N�$�BD�&��g�d�8� ����/مMV�+9e�ڸެa�I�'x�(&�Ѥ�u�VQ�qԎ�Z�dW3w�Sӊ(��1y1~~�z�:�_�=���,�(�h���Y�f��v;�[��J?sw$^�M��a�s���īi7n�9���r�5�H�e��&=,�àADs�G~��ܹ�V�f�yM�a��d'G�A�[{�_�4R+�ٮeg���1E\��gjm�vk�V�:��G�"���;,�+;_���C�)��I=��)��l?��1p-"9��+��b�G����ή�ʡ�TjXD���p��$ػ��^3��c8<��B��#s�rG�0�u�<����i6UK�"����_�� �w"�)��%�mj�3]�'J>������4�S���лJ��d�_68�z��>	����L8�%!����l_x���V�i�����e��;{cOo-��M�t�B{��	�l���+{)`��N�f����M�(2����Z�X0^�%i�e|7Ǭ���f��u+數��җ!�6��I�z宔��
�o������Cf�ao܉
X7c`��s�vh���l�!� ������b��yF8��������_�]�Ӕ*/O]��W���=�}H�Y�66��+D%V��O�n����&V*���D����s�:؊�KI._�����;x��l.,R%��Jw�@+���ߔ V���e*����7�l6l�@���AOV����.��<��ߦJC�ZS5bUZ���(Y�$�x�7L._W?|n$��X1IB�<ߝ+�m�d=V���u���(uxԓ%�����w��?������Dx-1�S�3���I�P�/҇2N� aS$W�������������T�����4svVQ��Hr�[�>��kvo���RY�����y �A�@�1{��/�qY�!����D�b��u�<g�!`~Pp"��M�iM~p�V���sENh0�T�z}g�0���ţb��uLxG-W��k�O�t����Ԏ��7�a6N�Xg;Ht3�p'���Ճ5�N�MM����� %u��� Y_癐����k�gñ��R҇K\>��P/��v�HsYCK��J�֩R��?����y��-�@;��-�������M�HLK�A@��ˣ�`"��P��%j'`[d�&ȇ��6� ��YpA�G��>8<m[Tĵr�ň�2�@� Y��Ep�H��t��䗢�r/1iG�Ug�xԚ���q�ʃȿ6r������Y;p�uN�:Da���dGHE~����!����qZ����Q�K��t7H��H��L=�&^�3�ٴ��]��&�r.Yؗ�M5��GcX1ԕ~�X�:4AsM��w>�v@�B�|����6�����,���r�f��mY�)U�ha��/����K�ne����ib���ܔ܏��J�[����i�c��{�Q���'8�B��E1(NmY�b����VM-�޹d�q	+vf�{��2�H�^{e��bX �2(љY�<�s[N���tN'C"��`5��)�ಃ����ƅ��F�7�^�,z�ʰ�7A��MN�2I���J>��������1�u��8��{~;���l6�C�L����~/1r�?�샚1��K�v��`�#�IW�hJI1���N�W��cV�����ΰ�bt��g35�C����C���[TK���,͇S\(�|�7�WT�a,�O�0f��RE/��[KJ���r��@ap�H{��F[�Ж����=��	��n�#����8 �#g�.Q�	,��~~(���-��pذ�c��S�t�Q%�����-&��	�ޅ>��Y\5\sl#
ܵ\�o`�f	1ƥ�o{�}�SQ�CU)V����*���7�C�]j�(���ѽ)���s]i����s�!�*,��>-�ۻ���g�8�t�kK�/j�~=�Dw�*o4��˂�w9�Q����Nǥ��g�㭞�_D�: 
Kń@?V AY���C���-�L�eM�|�*���R�?5߭�ԡM�zC�7p;c��;]�k5�7�Ѕ�*AӉ��  I}�	(wr_R�4��]�z���)� jpW��x�#�PHw9vCQT~��8b�d��Ő�W@F�;Gh���b�R�����^ڎ�q��,�7�P~��ם,��	�����˦2�3;������|�ک򽃛j���!l��:D̚�A�i*̛hD�3�#���
���9MַRӿ�<�e���B�f4i}tN �V
R���i���T�HI\Ó�	�#|�� l�>BX�R�.!&����$�v?S\��Wjq>��gZLH�noPqĺ��:������(%C!OZD�Т1�<]���>���w1��'� ��DͺWA�7g�휷xY�厐��{#��j�J�Ji˞,�G�gk2����d��+�D�VA B�����T�:~���$�Z6�+�t�����ƟO�B��JW�����T��qt�9�k����Q_�OEu�BAk�$�eX޳���6����M��QɑjA��x�n���~r�8���X�{Z�����	ΠgZS�O��|�^n�E�?��8���v���.���O2� ��4��������Sdr�#���3׃��˯Y_|��w`(XY�