��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&*���α�&֪_�ս$9v�WT�][����N�b2�F���x�+le{��L^���j<=�w#C�.L@�R%������}�.d#=�ʳ���;���C�����<BǛwjLN�S~�&�H��Uʴ��l�t7(#c�{X�v���Q�Y�Xs[����W��9��E�v�d[�'q��h����3������Uyr��i����K$��c2�-�2ٌv��+8�-����׭�a�<�p������M�B~즢�E=
��B�Vd �(8�q�!A�2o:���c1��џw8}���O�l
`GFi�v�6k�O���`�#�B�����;C��ur���6y�0�I�J�w�	����fه~^Z���t�:�����)�Dċ�ڂ����H�|4�90���'���z����1�W�\����u |=���/����l���E���i�RXr�δY�h�F�����rғ��B���O���ē'ұ�:���!�0�k�S
��c����-�x�u�����ns�~�dQx\Ų�d�g 4��{�p�X�H ��aE���F�5_*��l%���vLT���p'Qw��e��|�>��L>(b���'�����v!�靆%����~yz�ul���(0����
��t��j���iL�T�V<�;�&�
��Ϧ��,�R%W�_m���	��	q�m:5rK�+��O�p{�2�bӀM�D)��1�yU���0��ֹ:5V3ߵ)��D�dxl�	W4�Yf!^�E���\+���Q�?CA1�hɈ��3�`����DP��c��\a�p��M/�)�XMŭ�.��9��*�	�J���B6;��c;�&\[9NϪk��O3�F2w� ����;�0ߦ0���ajª��ߙt���;��W9L4�G�\`�|��l/5�@���ǬqR	��|��z���~����-�'*�\Ƥ�R`���9z�t��ܖra9~�~f/O�g�ݨTX�m8xN���d/=�v�LÝ�;G���Ⱥ��IY`�T��al�~�Wr�g�p�)yE�𻛻��͕��S�ξ����r���)�I�ց��ky_��<H�; 9�a�jk4Q'���X��~W��g}��F�?�޶���� ��V��fx"�n9�x+��R/�)-��Ec��e�&#����a�i��s�%"�=��L1&Zg�s/\�4�m��q韭+��8t�5v�7�OV;:yЬt����'S1��.mg���,Q��U���yZԞ-�K�����1������J	����S�xs�[&Aį��A^b��6�
a��ђ�K*<�GӾ�[��:�մ�B������2N*a�aބq�5~Z�.<�rd{��$�R�{12��Z�;x��W_�"-B�k�)��q���oU�jҵn]����eB
�գ6@hi�1����חnZ��tp� c���FXf����,f�ojT�_�~_H	R!�ά��a	ۖ���'��jM�1�O ���ɢ"78��͸x��N{>~)q�p�*T�D��&��HU
Eo��(5M0&�O�L1�M\,� ��������h.mGDcm�BB��n{��ݰ'���7xI��
���ȓ�;O�nWlk������G)�����L	�sc�#ȭ�@X�na�C�)No�>H�۬&`��f��s��;���������,�Kbzg�0��*	֬'~�<=�F��.����?���s�s��?�N6/x/���mD����I�WJ�oW�uY��%d���}o�ھ�ey��I ��&:u��t�OI�D� `�~��j-���	&�d+��4�e�O��`�������~����ش_���}�I��3kk��zj�{~<�(�w��B��\8�*�E5�-A:���v�}�}��`0`rدM�ӌ�D[>Vh�f��X��\�);���m����[�6�ۣu���t����,<~�����p�3͓��R_�s<N�G���ΕL�J�<"ݶ2#��)�W,��熒�����i^�������í^�`�� ��W/S0���>̯���J ](XŗܧA��Z��X���+�M�������ni�ș��V��;[�FB����'S��[�ce�"Z��p�d_z�F����۽��7�rA@��"L%��G����B�E����
���W�f~���N&B��j��,��w�����*����O�"�Av<Obv��r�n�㞄��N5Y����y��� "��W�@����p��\��mP۪����x��t��A!��3��[Tk�w�𸐖��FI�����؉Eɗfb�8��$�Y�P��AN%-��EO�5p�e��	�NdM�i�m�i����{��w����dA�`hG��,�o���o&�>��d�ءa�NZ�MЉгa�
Q�A�%J̊le�v�
�2K݈İ.t�y���%���Ʀ^aN���W��Ŧ0�2����E7�Ո�~�ƼI6M�TH�kc=G��g&�ciq:T��)��Z���� �%�L��4V��^�Ef��3ejp���_GO����.�9+IHV�e<ó.�)X$�O�+@!5��4��M���wꚙ���nbƞ��FW^�j��*�tA��{��TI�[�܈:�5��4�M�:s�S��ʊUƺeo���U�h�˸4j����h�}�':�X.�9&���rd!$����{-��Iz�5R����-!
S:+/���p-����O^���Y����k�|�_�gb~����wf}���["p�n�A��&i�`V�H(���|�לU8�+-����V���w�������Ev�n��S)��B���������f��L�