��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�9zrv��^�t��|솟<���+Wz��ke�q;�"��������U9�:�	L��������27�u�Z>y۾�j �|W~��-܉�L!+�!X�%%�¹%[O��U��UA�^�n�v�)e��c���v��o6ٖFX�E��SN�M�8�SC�}� 8���8,M����{4
K���#�4�k}��#�.Qԟ��Ԧ�"�_6�>uo��2����~ �L3�b�q���g�~�G	�� N�l�<��}�|�XN7|� ��Y:%��(��6S!@~Q�UC��~�6�3�"!��v���,q�|��T���>\����-������@b���\�F jm�
z��?�����5�yBG�_t���h� ����1<��|8��v5��4*D�*͚�L�an?aYԦ��ؚhJq<ݜ|\u����r��
�!E4�b�4�,:��9� y� �l�����g;�D
�@�.qm�2n���.�������u�8.韥eM�|�ܻ��	�1ϟ�%�u�H>yEd]6r����7!��p]�	\��!^U�;�k3[~!�ꞡ�k=�o?�_��i{}`v=�D�J$ETV��f{ﺐ��Oa��6H�C�kY,}=:T���#; �:����������O��-%����D8��uy3b]ڥ�'�k
< ���^�����f�e�Њ^K��9���~�W����*Wj�n�>t�TWN���
�D�<����������c'��4R���"D�\����],�b�)����+�!�� ����I��ƚ�/�^}�oY9���қ����臡��}{�� �{޽a��*C�8=_��G��B�01��\�r��2�|���|^|��(o�ue`D���,D�7��$���/��9'x���|�r�fL�E�7���w-�|m�u ��:\��SK�߲���C%2����iQ���!�2����.�m@�K1)�ij�Z�goMPp�c�w��;��`:t��,�2��5����A�^�>�p��E���Z���+�j��e���-�G/���E�-ͤ����DF���7"O��?��޼��wuxw�B����6��%�]ߓ/=B��b@FbdV�(K����$�1/ +$����3�e���O��@��4��M���2A0����;�
��s?4����m}J�A���ψ��23x|ϖ��%�#�������|�ֽ�@�"�H�d�ڻ@���kYwœ#���R(hG_�lD��{���&��q��x+H�K�)p�(x7*8f��C�2q4)Y��)[�4Y�x�P()bM��kДMC�lhf��x�lۋ���(��sX-?[����>�7�����,4ス����⑋M��R�@��w�$�E`T�|���<�~���fq��Q��? ���:�hKp	mm��w�c�0*�}�0enB+�:�k�[먔c�asǶ�"� .~��V��>!Z�}?��0T�P[������|���-����;�g��9���?�B�l%Ő+@~�뾭�����C��}�v�*�64tϵpT�/%#-?866��^e�s�b�O�����&�9.��!���;��;�u}F�X�=�ֶ:�ؐ�3�Fҗ:`��[Ƽ �s�焂]".�"fP��[@_�U�bzT�iE�Io��x.�)��p��0V����P1�l4�氬1Z�u����p(3�p���0��.b���c���&{��Q���o^l� c�S]ٲ�a?ich�(��&f�V��@3�ll��=@�;���00�L�w`�g�訡�akE�{NڥVK� %��{7���q�V��S=�'^MGL�q6�{������iqRԼ�X��*j	������ț���9�Β_G6b���6�p��x|���w�ڞ䩿���,��b-]������f-"Rlg�Հ�Gw��P��͊@���	�ز��kI��0�Y�_���,����*���|�-7��5���R�&8�w�'M9�J+4��#��l?t���H0�}���E+�1�+)P0V�X�Y��@xXs�h�y�hvf"�߸����Sm�9|�,h�k�����f���^��qH����EwըIJ����4�<qn�@�jf��%�/1���L��FP��4[��H���=����K}.᫗�P�R�hV#����x�hB��/�К�Jwe�����h& �/��i�7�Ef��oF<�`��$�D4M2���=�D��a�h-M����4���XI�AZ�q[c)��j֮mZ�����,j~<����
�%L�=��@y�H�"�����'�tB�<�ko�~d�Ne�C��ݑi6?���V��\X@�!��	�i��W
�&���K�Ff�#S݆�`-V��(�`��;�$!Ґ�� U���4�'��?̒�>���rq�5��JA;�<'2�u�AmCn���_����ҭ
{CfQ�3g�������a:�R����IǅGuH��T��N��m1���ڭH"MK��
����ZX��p��X�	:�}��u�۸�J�0^<2S���ۑ�$��LP:��d�Ys]�Q�D�z��������?�$�P���m�}���V������W0�x�M��$�ȃьg�|A�L����:���f�Ia�\�)oF��t��WBN�������{U'qaΙ~��%1RA�AY�����߷Vw�@:�m9G�PF��K��D2�� �4��)�:_�M�鯍�gn|�|�<1{�y���6�m�P��]v��[�LU���I���'�FR��7�yn�/�#K��ӂ�H%"D}���AA?���30�'"[ؿ$��zط����^C(�ߧ�/o0�X���r̰aZs�-�;���K�)X��Ck��0��$�R��#<�n����r�W`��l5����H �<�ǿD�d�h��jС�ƞ�B�I(�M5�x�)���h*+F���Sܬ_�80L�7������s��V��>�繗:���
�A��E�H)��ї�=q!iG=�2�j�����iM��M�(o���v����T�\��K|]�?�m�Ԃ��"����&d"�xC�йÇ��[�ӎL���	����xy�Y��Q�pԅ�}���c�%s�e(�"h��j���7��JY�䶨,�o�]�[��F��tsM�RK���؞4����  vw�%z��mX�]��'u�8��]ivP��}��\�]�b��蛲�]Z�bn��Q���r�e���H��I
�}��tSF-���DYޜ�	�i��Pҏmapr��M�Rf_bf�"7f�Ix�7�yXg�86�r|������<��)�%��x�X-iS��Q6�sp��e�k<�m_�5�=�v)}�J�d��_��7ԁ�>:��4Q,B�,�d��� {JQ�t-VD�`�Ð��1���"%���ͷ2L%%a�����j4���d	C�ɫ�x.��SеN�SzQ�A���������d�rB�q������(�/�]8[�D;�r�@%�M8}5�5QpL�[v8�*i ����'���d����y��I0�N���iO�Ф���}�����<��/|�3��3�ڮF�< ����ԱZ}����m Ɂ��kT�P|,)�3����!�$��|{�g5�-�1t��,"qw��US��i�Y�EЍ*\��9�3zx���Z�@��ő��sE��2د�.��� (�r����v�(E?�o�ޱ�x�϶�^���� ߯��#rA2���īk����A|��f(��w�A���T�at�B��	{��U�X���"�⓯ Q�QW�ƈ\u�O�5HPo%�W�0]�Q�SW{VR>������*���w���b���S���R���X&}�0���-�&�r^���  �03����~fԗ9y!��ƭ��z�X\)���C����;b�j���.'��x1,��/vr.i�I��+Vm�Z�*d�&1Q�L�Χ�C�뺑�z����t�r"�_oD�]5EBEt�p6+��\��f�3����>�
'�/ӵ!s>)���1L�5��_���k|��* |L�M�>�P&�m֜<xt�4�ޯC���.�F@��lY��<�/�4�x�r~}"arϑb=]~������@��u�))�	5�F���Y�������[X�,�Ο��p�$���1�
�i��g��k�o�h&C\L��.�%/���ݪp��)?r�irѭ�ͅ�0�'��u��-dJ��t�?�+��Oz0Bn��L\����>1-H�L��f�!ٶ����h�=:A�܊�a��7�l�Q|�q?�w����#�I�d��`�K�BP�k��8��Rچ�?�!��}+����Oa�)FA��������:$�4�ZYG�ر�\!��`�5G-�$���G�6*�l��������a�"�'%�L.?�n�d��J���$O���\����F��&��`]� :dr<��V�_�%|HNH�a����"��r/�E_��g��ZJlѕ��ٯ��3v�J�ç&u����Z�tjZ�����s����
^��'��~kF)����ǰ(:�U��N_�u6� A�=
�n=iI1��/��-���b�$�f��	�|����7����,�P�.��É�[<LV�=|��y�Sf���;�V<�͝c���$A�w��?�+JG (�\0��=� ��Sc�����d��i���3����J�)���G75���",u��gSř�j�Q_p�oIKu�W�-9���j��C�uG�R�H��H�-�;7�G���g��t?�F�fj��2Z��������GIP��
�	���Ю�lb�kXV}������X��yQ��_��CyH�ѝ>��S��0Rs������⤂Y�D�7C���Q��З��CU�O�H�Vp��'ڥ_xM'/cA1;���K�|���,��£R�zE��x���F�Ÿ�0�y"7�(e,T(8��>>2�.���s�<Zg�9���� ����p�܉T�ZdaT���d�%��g}i"��/d��������b���O�K���|Q8X�ʁ~
��~7�I�!8ή-ckҞKG]xYr��'a^KH7|*g��FT�ft�Q2/���N=����^XaI�)Qf��eR�6��V2^�y�4M��ح�n�v7��m+@QQ/�����Ə<ϭ '7��ję.��А���x��B�I��lB`P�:-�íj�^H��rh��3��M�3��L���q�oO���ϤH�fQ��[]���J~��eO��5ŀ�^�ב�2ϹYZC���O�??���,N��ѭxzg��4�?�u�z5)"�i���*O�[O��X�����H����c.S��#�i�5�MU�,mE]=��#Չ��|����M4k{N��l����ԧH���KS|ז]*���`�m�C�ق��5EM.j�HS����֣g�y�����?�e��\v��dg{�S��{s �%�<�����;�{�c�يRg��O�;�=�$�ٳ�\�5�/�R<�)c^ʊu��mܵ��<BN��������2{��x��mĚ\p�����1���b=�<�:QL�ʕO��eL�Sy��ʾ�����?�MY��V�+�����%�X}��`��nn
%C����c�Z��~��@[���i�D�#�ͧ���V�x+��N544�|��&����n���O��e.��?B�����l)��6��%����q�)*�-b-�
6�p+��t _�pm�4{��1��t�6ď�Q=�Ɲ�&!ZHd垣�Q)��땵Se��S��f�m�ġH�"ͮ͢����ȧ5�� %��'/-V��9D��.d ��������0���sb�$�'J}��r󾯒a��<���S�S���;���5�/�H��&)�Ϛ�a]����F54暗¶*�Zb.xeG=
wn� 8Ѿ�9��HN�N�#(�_���U�r��/�<F�~�u%�ֽM��ɎoJ6�2�����0���!�f�O�$�`N��C١���O���J��ca�g����x��ߖRp�����Ȇ�1`u��}r:��kA�T��k�k�(퐗�R�_5�W��1��.����V��2;�cӈ����/�9����vt�ˢ�ek�R�S��l����̝�	A����N���j�+�[������x1NKQv�\X@����d�wy:�)����o<���|?�6�MEպ��ȳ��4�#W��#��g���X��n++��W��*�@W�gĞB�3sH�)�'Н�8Y��P�d�;��s>��&g!�5V�+1��[���Pj��g��Hwq�z�=�G-5x'�__42��m�4
\L��ӵS`GP��Ӊ�'��w��H��Lu�1"��s�;p~��h���OJ^�{u%�Ơ�X��l��س"O�g0'x�U�R�O�s4�'.P�h�e�'�~��Էu�,�Lly[WD:$�n��h{*|��hw�m����Hj�w���d}]��\M���p��SҶ��'�<��K���xh_�����I\�
��)��������=�LV��{�̙\���nx�Hoe�R?-'Tv���U�������'�>�����!X˺� ��ƒt�)|���2�O&���xl@(2TT,�t�6gx���vT5Z�L��>�d�R�j�򱓼����=���
��O�f�N��V��]Go��Ŀ�H ,(pX�U,��A�|K<��4	��`ޮ*u�""ce�~���gfM��!x2�v�.�+/Wn![����fbh KY]�	C�~^F"�iEHk���r��C6S=��,c��Ot��'�hݳ�=�.���k5�m�Gى�mF|�_�;�����uK�=m\I ���|�&fp��B��mL�� RՍ+�pW̸�:C~^�_��I ��>+~��y"er�h�_�o����zY�n=�^ܣlD��O5�Mla��X����5��<rX׍١c�-O�3Ψ7��89����gI/��@���,�{cLW'���
��<��M��58�O�z�$�s�$^:����v��~�����;}pր-��+FΣ�?uAC�A����
�dU�~���A�<a�W�eW)�AHJs>��< �����R�&�Q'����"����?��eq;Spb�q�M
;�tk[�DD���ےG~A7�zh؍��4��Lg@@js�2>k �zDf�W}��o�lR[*��5	�\���`J���,�m�
�������]G�:�������٢�f��Z^�7"�.��fx�:�͝A�ল����ϸ�h�U㡞���g������m~n�W;��w����0��K�{��@���<�a+�uy���}�in�������qk�ل��e��`T�� ~���:�0���>��9����.�?�K������+�?�<��5��,�����'�������i�*��������Z�� ��xz�����{D��V˰@��)N�UG���=���T��%1A_�`r��
N(Z�%�7Q�(D�����zD4�4��sg�8;�ԫh�;�eޅ<��I��f�_�u�Ÿ���������ٜ����k��~`
_��g��^���>�E첶"Φ7:K�Sw�x�LҪ��ѹ�E�^� ���{����9VI5)�k�{�����P'L
Soo�b"���͎�L`�s'�H�c���(�yr�\\�{.�?���B���x��`�Sp���A�Q���X���2&U_U���S���
w ����j�[�24/�p���R�M���ڝh�	���b��;�|qfS(�p|<GE+��z�ta4#;#�r��9�56!�}3���! �v��H��g��B�&ǰ��z�{��v֨om#_� �S/�0�1�n����&to�$Y�awITJ� u��'�_ǔCg����z���6{�o�ٟ�2W|�3Wh�TM"J��=�Ӵ*���/�4�%q_G�n��텲E�)���I��1���l���NX���v�:��������%��lk�[�4|~\�����yJ$�k��	z�$6�ϖ ��'�w��U̸��r�Ԓ�m���4I����l��e��G��es�n/C�A�[-����7�����Û��j�6�wF����h�"�&;���0p�e�\��^u�EД�^�_�Z�F�y���o|�����v���\���I���q%o1�Ͷ/O$��E�ٚ��S�3h`�+�
�# ���i���e�ߦ�dE�6��Q22,�u�w�B��T��~:}��2�A�b�4.�t���F���-Pm��������(��igP�L�%�b�簀r�}%T��H$|>��;ӚD��>��G��]��KXn��0Q/L�𸢓�H����b@zY,�ur1�cI��wo3�׌�Ei'j��?	�>����e}�5(�L�(2ӵ���wI�E]c�f�U�b��5�}k[n��YB[l�`d}!v�c�ݤ��_Bm���uu�-xq�(���6u�����G����X��j��8��{��<�uZ�����u��p��+�Yv��tЕ���}*i7��l��f���B$r}�Xu9����y���ae������ov.z*�;\~�Es�J	>��H>iw�4�ve6�B�F��]���h�A�~����(~���]�f�Ko���T�:u���,���ƀ�Uu>��t��M^g�:[�qBBz������'$3a]YU�����S��i��.q�#ުn�6�$ѥ�;i4"�h�@d8��Y`�T�w �ļ�cԺ��(�w���VJ�f����`�a}���������OE��^o��QԽa��i]���U����ԧ�蜏��D���ك�>����S��+t1&ӄ�*���g��`n#�>�n��g4�s��-��@^�Um5uE�G����~��1[�s����@��S��҈{�P�Oo2 S�gh��/��b�C�7���ۯE�l��f7��
��U+5ߕMo�/F*j8i��5Z⢪�p�W 6�W�S��Y���p"��8u���e�����3V�zWPOw�]����G)��#�t�@���_��0BMr�<��;՚ri��%����m���Z�F�W���Ͳr�wc
�~xw�*̬.M��$��O:^�,B���oC-�� �b�0����tw��>=�~�aG��I Q%��j�G����E�]��Qy��PEi��$�2�\�.��]�n�b���<~.������G1%=��f:a�fa
źݫo�}�����R�:��-�g��*'�#��#\����+�r럾p�e,ӌջ���/8 �������M l�7�)�(T;��[&��5y����@�<1PX�V�]��owh��R@�ev��o��D�ٰX��0v ,c�c�׶)�*��Y���q)�z�1�D$�mHip�l�L�ȋ�dM����o˼�q,,�ͅ�3ޘ}����8f7�Mքx���)4�#���T��������$8w��^\|L�PY�ʟ	򥵜Fu{���>�?<@K�k]���wQ��fP��oiB��?Ȗܺ�+���6!�$����� wzBs���,�3Ͽ]h ��G�*z�sSA�#���f�c�L���g���t~ �F:\�m��.�0�gB#jnk���3��b_R6�6*�{�k��!ㆨ�Y�+�[�����PA� 3l|�%��6Ue��^��G"8�=7�`R����W֯������5�Ȱ궸I(8��<�KK�Q�cZ��	�׿��C�M滠j���YIϷ�f�tyI26L�cJ1g!o�\Un�=	$oi��Ņpo;��C��uD�-ŞK&��l���nu�3J6�8�Jo���i6��"T�@�oF\f�6 �K)��X�0�޻\���F��?���|���z^!��֫$�۸ve2�^·:�7���ȯ�P�Z:��{US���M��?�щyQC{�T8����;M^��Ed52\�^K땥�����#����s�Zh���uZt��<7!un_#m���hl�rR��M�@A�tj�k��V��>+�弾����G���g%��~Z��$/p�$,�/_x#W���� ����P�G���YӞr2��	�J��H��iE��;c� ��r;CF���#`�q�1ˡb��f�-�gT�웘�(V>�i��y?��*��"�'죵��R�#���=J�?��>� ���� �yTb�`���0��0ݦn��5YYi����_ؖГV=b)�W�eA�8-�1Nd����o�yr?����܏1B���� DC������QlxsIL ]�e |�r�MI��I �*�LӬfp�ߌsJSNS0���$Nǂ�r �}�1��vM�����n���T��׿�Bmܒ�NV廔��ֺW�D��ŀ���
�D#z�ת�`L�sĔ_&�?ڈh�.G�Ax��C�)!��{`3��Z \ȃ]~`��}N	.��/�ц�����]<� ޺k�b�@���V�,ǃ����sWlc�{�غ�c��`h�����vZ=���ft*�f�WyLH|!xM��j/�w����bΈ�I(RfA��  ��Cu3G��L�١O�d?AZ�5)M��(i\��,�X�@�7���w���D���2l.�Xvi�$� �������)||����V��?���mW�����'dg�{ a5H��h�qr�qwa7��,��/ei���$G��,X�$�<�"��}�fl�>��bu(n�qY�6���7�W7�Z1� �`�]e$����i���a@vȾ�� ;_�c�P�s�]@s:'s��ҹ}�#�R?<=QSϳB�J�L|t/saę�%BN�9��������=2Z\ S��%Y
��V�f�5��V�%�����r/>��n���&ߒ�~u�:$�d����nxn"�Q�J!���4t���j��|v�Z)>��?�&��B���Rl�|b�Y���[o��*͍��_��� ,M��Nf?Yu�5u�&x!5`j'��ŘD<l?fͨ���f��:̑�&+�##n畴���;PypXX):�6M���-�\w5��q����:�t=Q4iI�?Z�q~� ]" 3k��d�x��%øl��|����1<6+NѳmP�t�
��N�W�� ��w�EG^�)KW���qP�j�Ugr@@{�,);���<�y�i|�v��0+>�K�z$�h?l�Y��8;|�� �Lc��H�gS�!ʅ�,����7�+�/ ����4jX�]�E�� ��y��i'���������g!(� �)G
M�;��E�*�8�Xq$5�<���:6�*���&��ͩ������ մ�����u��ǫJµ󃠈7W<z��~9 3TM&k�3��M_?H�A���	� `	�*ʾA�4��M�9x�����
cr,���Oڅ7y]��9�L�AN�2��.p`�ep����TOj,���bP���k�R �Nz���ҌO�`�ӏΛ����R�G�(���o��]��q�DnY���]��5~4x�ҶH0S�b��R���3nh�rC$q�*P���%�C��r���c-�Z�0�.
u��B	Ý�ڢ�Jw�m�D�:mU$�UK|��Nh:@]ˉ��/���#5�Cj.@N�1��*�ܜ����]Q�B��blx�K��_m{�Qh(�΋�^����ʧ�_�*���Ŝ��4���p��$Ӻ�#[�>	�Ɛ��h������]E�`����b�]K�x@ϕb��bё� ��=E���^����ma�s̥�N�>�ǰ�����1�W�m���7�R��<��u<s3����O�d���Y~-"��P�����~ߵ��lo������	k�\'�� 8�Ȯ-ޫ��Ϡ�.�i�LȪ�x�~�<�l�^�+&�i@E������@c}����QɊ������1��2�?�+5�n�۫-,�FR��'���e�C�Z��TN�?"m�U��}G�!�3U\�<�JKiC�H�	?��d����Gx��0�β��ˠ@8�8F�>C�fg�9&fq������;!5\~����4U���������`��<���73S�-Q��f�\���@�g�,�M,�m��ҵ����B�=a�ǁ��6%�z�S֍W�3����7����oc̊�W��s��}6�C���X͋ �k 5�!��_�Ȑ�EXS�����	#���;���	Y�7���;@����]�'.B�d�;*_�I#i�M,d�5òJU0�\�yF��uc_@��[��b��2����`�03ҔeI/�y���!���j���ܗ0ɾM�v#���^�S�w���\����r`́�G��t��v���29Jh�ѡ��3���-�."�8�NQy��i_j�1��]�Џ��"B$�A�rPz��|#���Vj�Vw�v��q��bT��R�hݷ�d�dGڼ�%���}!A�H�X��,,?Pr���J�.����`m�W�$ia��8� U�s�«�m)��\����jѝ@i)~�t���Qn8�D����4G���1d�w\ʩM���Q�}�ئ0S�m7�϶1.fR�wO�0'�|S�5������)�)��}���L ��ZF�$@���ڗ�Kl9�6���t��9j��u�
�d�����쬘�~�[�ᚙo��D���ޑ���d��\݆����{W���T��ѕn����jrUp/̍c��f]�"Y7F���*i5���.�־��Cc���E_�ݜ�l}������-��i[XN.ӆ��-�����X�n�ח�-��}nq�P2� �,���O� ��uiS�O���k���%���s%�>�Tər�Y�Ȉ���k�(�������<r�]є-r��Y�Tg�!�Ʀ
T��1��6�0%~�a�r&۫m��q�2��56�i�Ay%��y�P%[��C;)2p�Hj���L�s�t�z/�ZJ��d�#�hL�r�Ȗ~��f�t�#�����I*�ud]�U�K�xW���/F� ��#���
�:��u%��VM��՗�n�Z;Z��q��O��-�>��T���7a�݃��'sZ;���0[}_�u΅B�,�+5�K@*;�>i�6�#i��������H��IAϋԼħ���t�f�}乻������[��cu�t�
����:;X"_���<��d}}%?Ԭ�Ch�¨K%���M�xM��$	��>�W�c�z�Q�:gz��c:��I��s�GcjS�O2��Q�U' ��&�D���
`l����� ,zʸ���N��"��06+����8i����	�7�D�y
��i�d�����m�.��Sh!�n�#?�	������f��f��V�z��>�&��"*6ˌ��5�n�L�@E�����2�[5��Uኀxv_v�T'Jp���_��9Nj�t�ݘ�~��}�}]��<���+�k$_�M4}'sQ�vƚy��-ᑊ#
x~��*�ӿ7(�i[멵�>{&�3;ױU>�"ľa��B��	�6-�ܩ�^�c�����}��5?�3G�f]��8���݌�u��AW�����@�"�Bt(� B㘞I&X���X�+-v/Δ*j��}%ç�Z�I�qs�To.��E�{b�S��ĺ����J��g���'D 5�L�R|`�f�%�c&�2d��-����ޢ��ۆJ�� �Q�g=F꣤�l���W�gNg�2�Jp��Y�3�6k��6V���������&�R����`���?M����i�d�FIԇ�9�)���K�dW�N�p�P�J�S�8+d�O�>��d��8����b����Ҵ�~|�eC��{¦���ҩ����YV1���.�)�l�X����**AV͑t�;�R���$��:�W9���P��'�$��_PS/�Ew�ig?���͏�,�Q�Nz�oK|�BH�7r�A�Yӄl	�����O�VU*{%���p���T~�TFc�m���
�$lL�~��Do9��c�W�w�� �7AI>Ɲ5�ܣ,��4x��p���2~�דY�1�h��o��jJ׫�X|�)�s�<����٣�c�gmEmb�YU53�N�x��^GUJ{��sk�67!�cafh4����fF����J��E����d�4�`�?meT~#�*��F9�֖!if�~���U�bPM��=�u)�{Z�pq�����7�?%Ϝ��4!���@�r/3a0Ʀ�g���řȥjyT�Cv�k��ˡ1.��v0��^��"1�I}!��	6�5�9vL!���n�'��+A졨���~��i\!��;p���z�0sZB�f2b$z�?|�}}��Իǔ��ri
��ٕ��b���u���0b��m���7F������+�?t���[�������󿘉y���Aè�iC<�VE���By�'��������)g�1��E�rO����E+'����_����IvpF�t~��_�d;1����|URU�Y���TJ�ͣ#O��[�reQWow�̓���u�ݠ0a�1��T�;G��GE��aj��(M~�~�/�uvAh�K��(��O�v�k��8.C�bŦ[,���]���H��]7�{>8^��f؎7R����65�uu���s�\"�ާ�;E��?�x'Lƈ��/���d�	�k+gB����P�c
!ƻn�RQBL�q.�FOW�W���U`�[���jtZa'xATV�bz���N�(L7����B��a\̌�59�#W���*y���N�G��>lүl}��18�d3C�}+�� \�
��U0��C�=n�EG�n:�c��;�9��|����,~լ���jܤ>�jV�EMn��F`�^X�Xd�)w���T�����-�,�Rk}�O�%���~\�}b��W�׈���|U��;�� l/J*dN��>�q�EfX��8^� d���%�&�Ż�9�6����Zt�C�H�	��Y��K=HR��I��[a����&���M��Eַ*K[��qW��"�?u4��]�l���ع0��9�`��L�\���乱Ka�'��;?����4�L_L�zD����ǡ� X�C�ޙ��-x���݄���`e�c���6�ٴص�C�k2��v;:<]g�GJ2H�,_׿
`=�5�����%|P��5��ICՈmܳ�W�D�V�}w�b�$Yo�q��<vl��	�0�C�D\�	���L�N��c�� �y��0�B�����7�Ib�>e��/����Vb���.�l�'oۼ�u+�QU��	�/��5��|�Yf���N�@E��[��s��s���Qϳ�^~H��F�nOr�k!g_��8�L6~:|W4kk�L�6c�P;�	����M�hڗ��@��Qi�B2�F0�6�C}�j��9�l_!�/f��"�@98�L�(���w��js� ��^��������)hc�6x��VtŦ��:�C$�)	��9%*C��0p��J�YblԄu�r�������_zš�7,�)��ݞ<��uz���'�42�u:��V�i��-�*�	��pЭxL��=��}&�x�X��~�a�̊�4�h�u}6�g+������P*����?�`��_=fepԕq�����{?�-t��N/-����xڇ48��,�(m\�5�?�9��uG���FC��S �*�:��/���T��d�I��4�Ctg`u�n��.ޣ�N"Q�
l �/��t���-�Pk��y�����X�W�ko�������-�
��b19���3����c9��yBѹ�&}�G�W$z�aWē�������4����#�v�0���Y4���#�?� q��^4��������a�󦳝�
�[��D�#��ʈ��=�5a;L΍�ޓrj��{��]�
�I\W�"��/M��܌�h
���_��M�A�o+a��5z��ٕE��8�X�t��]�d�fI�����1�d����^ ӏ���Ư��'�]�"�RcR�q�˙b��I��R����$���Yu�F)|#�6��s�j*B���lz"mŶ�Ƙ������t��{�7*ԯ����f����i��5t�����4�Bu��ޖ��,/D�J~�6����j��q����в����y��/�?���%��F`y�v�:��(��{��]!�X샆��HiwG���W����o~�\'1\�l��R6;���-kiO�AP;3p����b�آ�)iB�O�0�3`�D@	'1M2a=�[�K����Cy�u�s�~�[?h���7B=ƚ��tv��h���C}���hF�����E����G�]Y���PO/�0����#������z�d�Kw.ZT���m��ؕa��6�sU<����#;��O'��ǘ�!�*.�I�{�����t~I�7�}�x���p��7&�^�q��G/~a��p������W�-��В�~*K�g�x�ץM���<P�&rmS��gqwv[��N���.1(�[���~�A�N��O?��^��c[kLf�ɒ��p8" sV���Uy��<�x�a��r���)_,�ob����ͳs鯽5�'
8$1�G�l|Ѽ�*�G�탠(���l�{/�Si�J�%g���f1��$�����\��C�^�[_na��+3A���=b)<7T�a7,�>����kF����
n�v��؇�.��Py�QD�<�.LW[�W�WgK��T� Rw��\)lO�D0�F�@9$�4.�!�|L��_�-�ʃ������R˔z��� ��!������+Gc`�_��W��;z�K�mb^�L$Q��QB�c"����/�,/�C�^�L��A�	�z�{�'�S��}
7T w�`S+���F�ޗ�r��>�"���I�I[~��u�p���c�QN4��y���f9*S�P�p����:�Gn����w�]+b:.�i��]Ԛ?����u��b�'����S�סw�d��e�����V�� ��D�����5�Z�
M��2����	���uK0'�@��}t[��,� ��Ը[��4M�qhJŰ�3�8�ѣ	�C�iH�4zpʬ�|���݆\4��7d��qǭ�����%�<"�o�\�%;���">���s��L��b��kk�)��I>	ra�;j�������R_�g�%��T��.��w1��f���Qb�6���[��S/�O���������������$j;���>G��g��,D	�$���=��ƙ��jy��菥�N�?�:%�� �mc�q,�b1�:K�5-�Z�Ǳ�L}��G�-���(��]�X���NR�?q��j���5U�Y��R�ZJ�eAAH���=������|��7w�'&Qx��k.�t���Msm�u��%�|�z��W�/?YNP���Hx���*%AQ�������8���=����\�Sm:�� ���F�g����j\Z�KM��ҭk���:���a@Wtc?�+�Z�[��"a.���"]��ߠW�M���>(%�Ԓ��p�9N�s��N�}��d�=�&@��S,�'�y��E0��q�W5#�<���P4
���񔯛��8�����e��&�!L;�EP~%�x��gR��TuE6笜��9�Y�EA�����a,��A�,�	���FHg���9�G���*�(q�x�U���1�%j3�S���)��\x��g5�-B���%�ރ�Ou�ԛ���%�W(�ѻ�� n���n��z	���I'���
�y��d����[�!�:�V���AM�,�SB��cI�.��)�4�~��������G��}wĝ��H�Z&(J�h�l����0��U�kc?W���M*R��CU?/*;��V.���
Ir��M�H*�,�a��P�e�ߒ�����T���f�1�ժedjo�a?�z4����J��y��F��Y�P�B��i�Aq���������|��&���+�]颮
�6EE�11Z;��^9��Poj>=�kYW�E�V�s��� ##�(Zhڏ]Bo^�>��>7���{�p�=���)`�l;�*�wı�X�H���f8����oZ�e�X	��Tf���o��t�}�ڲHG���,�A�(I���U�H:l�nğ}�
9[�?��x�� �su�I�0�R� ְ7)�s�{��(m���B�Ģ��tk�&�WTO�r���i5?�K�:ԕ�!�S�l��)s����_o��C�G�`�y��XH��}F7)�¦yV{�Z���.�}�����lu�\���N���!p]u6iAwv�4ǽ�͆	��R웶W���ޟNm�^�@���(]GS�<��,B=@���"�f�x��po*%��~ۄ��]�bT�%y���$��jx��V%�
���RYI>�u��ސ���Y��Ӏ�qn���0����.�0k��|�W�CbI$�v+O.��������CH&��s�!�)R�à:Or\�.����cǔC�q��.*Oڄ��ӟ��T��G�c6�&�"Ǟ�ʊ��>V	���������$�Rd*5�L	Ѹ��l,e.S��&�a��er�	��8�y�{�x#�}:������q�W�*YĖ}=�`�r�zh�!9��CC"�����*f�,A���:������+
��t"P,	�>�pm���9я�w�䯚W�G��g��4�Cj�)zi���]���}^VX̡S���CJ�!���?>'��k{�.��Ps:�WS��X*� ��&�BRT�������S��<%)c�;eR$roT;�:�����%*Di�Hq	��1��1�t�1)&29Üp��j�1�lm��<�>�FC~?^9&�N �)��R�Ԥ]�r�=����)���G1m���՟����Y�#��������#^YcK$cV���Wr���0-�y�dx�]�1���H8�g��7�ߙ�C��.<�L�HG�?�������E7�ԅ�G���b��"�bz��v`��#lח�:	}�
��oT �XI��b�h��Lki�T� Sc���(�WK5?Rq3��0ɷ�"e7f8i�ۭ� 6"�羯m�fg͂1�P�Ъ��Ļ
�#��3�1�}�޻tN��>�U���%���A�Ez��GE�H9|�>f���RdnS����H�*��?�utZi��U��=��F�
�z"n�,�W�|4 �U̬��AQ�TĘ��&W̛�w���0In�?4��(�d�ܻ�CE���g�񅟲k�|���;����0^���i���ը�b_�+�Ź��_�.����wq@�9������)����c&�MǠ���!��q)�te���3�2��Yo\�Rf��.��F��P��I���v.|Xj���nr{�4@�h�����|��k �$���/�θ[�-����/"�^��F�h���dpkQ��ʻ(dT1N�л���*f�nz��I;M��<���,A�2�����j�����2O�O8��t	��@W@���jb����/ >�{���pf�B�	�蝿\���.��֓�7'(�XuT��z�}}Ϩ�g�N��U]Ɩ�(oJ*���D�%x��͕�!�'��ǯ}���AUdyp��b�Z4|���A� �	��٪v��JѲ���H�}xڄ��J��Z�R�ǫJsoo���d���<kr{��b$De7��6�����W�&s�k$ε~�?�`6���[H�a.�2Jf���ܻ;�7NF�ԡL���Wt��Te�o	5͇�"4����Ɣ�A��:��uk0����-�(���=(�9tҦ��,	�_�	���F��^�PuG�ح5���7jkpAT2�XGv�"��~��a��eP!T]l���0h�zZ�gr��;;�W��Q!�L����n���_���#;\�� �.O��s]�겚�UǚB���JRT���,������f��Fc�sN�܎yD���w�)��j �����k����Ճ���p��'��A]G���<��0skg�h��a��i5��*9s�6�<��з(��>2�EJij��{q+Eq�y�	J��۽O��,l�� ����cH�*s�ḧ�::e��}��M�O��t��n�@���V�A˿��� ڒ��B���5�Nq2c����7�j����O��ȗ��_GNK$�[�w�1�a�}I�'�E/�?ńܰi��������jS��ܯ��m�� $�G r�B�|�A�'��
�>QFܨ��
���4�����{,)�`UF�S$x��@l��ï�����0>�R�p>@�9�z �t�ů��<�d��Z{��>�B?�Z�I(+�츌��w�wP�P�^�%����fZ��2��dʊv��(�4Mi��
駸�E����l�ɗ-2�s�KrA��\��B*L��x����t7����V�X֜"�~�x�N�Tt�T;���d���|Ѷ ��Y���o�P(%א��c�[u_G���G�GzM��*��œM���xyR|_��Q���RT�g2+90�\:  ��ƺ��
���2�{�#UN�)��A�m.k���ʦH1�D��"V{�����L���$�pJ��[����X�w����O�!�<d ͮ�V��検���^���ῳk��9.�=�H�͘k,iE���_�D�w�[�T���}9���j[����+�%-�+�%�қ��"��NŨ,:Y�ȅ�Z��#��f�pг�Pڤ��e�5xY�V���ܼ��;�~/�;UX��e���t�txI2NJ�|厛.R�Wd�б��f�< b����j0��kf�R�$�m��p��$&B)���	���[�����#0�e'�^�u-�ܶ�H�cuM�}���%�4����s��b`��_�H�[�wb0��v�!��i�/"�*����m�g�����P��)��x�Y+�9��@PwOP� ����q.�~�ܝ����<�R��������hѦ�Nm�ݬ �\��f��_Rlf��i��p�y[���	��-X�O��oT������3�آ�@��4�`!��d�%�NSL)L���'�������3�b�C0x���D
m�L��6�WzP�q���c�%�J�{�����Y?�̺ �I���Ys��>a�h!��S�@�h-	}�_��V=n�v�*�8���l3Mi|���ln������̉dV���[ުڋ�m�F`x��!�}�cc��a`UR[X��������G���[SF�m��$z��5��l����>��D6]�I���e���_1<!���Qr��_?'�s4� ��gb3A s�aƚO>啃��$��Dqz�����aN�����+/Dow�kV�w1ddN����u�5�@�:�\�S�#q?�N<�(u�W��?��D�*+��5���7���7���}��8OP#Aۆm�(�󢫅z�����B%�c���3�yq��a���֬����;r�/:_A'>>ܛ�Du@{���4�\��#wG��W�7qX]��d䡧6�Մ��~�Go�PS��9��<��_�xW�5>��>I�z��`ٔ�G��;6#��]�I�c����ܠ۽o�(�ۄmc4%Iܽ����j0xO|����@!)>��X� �}ϊ�Nu���S�ys�
�?���h�ͅ���p�w��z��`ͷW�G�c=W����N}�E�h��eS漐%�[!C}��xx�cg�)h�� Aܦi��gO��1�ÈX�Xi��]'�:�;��^�ki:�x�Z�W9�ft���4���!�1�'�PβJi�y�u>���4��j����;�B]8 4X'�~f%���k# ;g��TS�%��MW�Y�2N��Ѽq&3� ���K�/7<�E"��~������L��↚����틸��T��!y!x���,�4��8�����S{���>��o����F��� �a��-+w2S��-omޒ?I~�ϰ���R/�q奵�on(#�gd(������i�'s �E�+�����)F�O��l@A��U2�lW(t�*P��6��\���	C��u�'��.���(��6��G����_&�HCX��n�c
c�B3o7gXB/��Yw�)�h��GO©ܭSĈjٷ�����(�Z���\�E��w��Iz������~�6�F����O��1�q)7
�3DxZ=W�2t`V�ub���V�TF˫�sχ���<}9���]��H�l�io
�J���n�ԏ��;
��Ƚ�i�}"���A��Z9+�CK�q9)��^��E4�a4���� �hFz\ X�rm�����|�s�P��v���A��r4H&�L"�L�V�<����S�IJ��h�^�	��O��O�t�]�����2�����@��O����Ѷ:):�4eؖ�jBGU>5D�aې>�)�Y�*C(���O@�w�f�>Al�A��{�]/&tZ�P��uhဇ�;X��!B����3��ޓ��	U�qy3��,O�?�ؑd��z�ArХB9�"�qU�Eɀ�ȵ�Y�ovDG�K �p�o��D���{�ێB4y�i�R���9H�x"�u�����#4L{��ԃ#�V��� �O�S��M֐0(��4z�~h�8Y#ވ|QCM�s*�u�t:x�Ǚ��j���JR�=���n�S6�|��oR@M�_����ش���!�����\p܀�'8ö�J��R@���ˮ�8����G#?���_��S�q�j�J}�tf/G|��
�F�R��0}��	�x��?��(����]w���T�ն5W��7��II����%M����Z��C܀H�s�3,�4C\�����ԑfv߳�+IZ#����^��Ʃ��h��E0u�.7:�羡�W,��]ـ\y9���\g�'�~E*��ġk\r�>h�n����� |�V����N)�����0��_T)�ܫ�k92"WЏMy�J��Υc⢱����럸�nUC��"F�v�}򏷼6V	p�(�`:�_�Rp�a�4���	������{æ|��[�9��!���*�h���Pт�Z/�9؂W�u����7;/z��6��W�f��H49-��Y�v���;�JN���Ȫ0u�����@�x����(I��$H!mh��^.wN�47Н���; ��._%o��,���6)u(yvx?�n���p7��99�$ڝ�<���f�ɫc�|}^�F��oꝮM�$���,m�c�z+���NK�U��ՊF2?�O�c�޼�^���Z&D��˓sKG�}�}����]"��!�N�"�0��1�U/��jl����"k�ZB��o����2\�@ҏ/�N�f��#���f�z�K�9�>)��:���X�M���+�I�_O��ǆ�I�ۅ^�:�r	�^׾�Z��酚��#
�-��L*"h�o4�_�}�Y7lJ�ε��������C�Q'*�����]Α�P��s^#����`@��DH!��m���ӡ��j�`p���x)��x�K����y�&T�U�bm`OC��-��D�ߣ�S���<{(-VЖJ���|�Q3�a�V�}�y'cZ�
^+������\�@�C3�v�++@?9���	c�<�g�-R}&�����E:�
����	D3N�/�,7�_�`t�[ k ���2�S��ch�D^A>���ܚ$���|zN�!�N%��)�D.���Q?�~��0�7%�$�_�QQ���_nP��!�U�ᙠ����9��Y�Ų���G�<�����S����hR�ioȰE����z�6�:����[4��L�_�������&Lt�v��Ӌa��\sc\e�V��1^��b"!��]���A5�E�UT� �:޸�z�[Gg�t�n�2�!���L��|�j�B��z;,I��r*v�{*�q=�s»�}��`���yc_�+������<�T�I}x�bI ذf�lr�`���a���v�[ZCd�A�&�7�"=Y+^]b� 	}g+�{ h��6@������YY�/˟��"��%�c�=GY]?:tA0FrG���O@	k�)�_7��{&�0�EAWC_38�xD����Ջ>���k���ez��2�}4Z�0��yl��;��5��k;��v�K��%�>��>�)����g��E�������gld�)X���H��s6������t�J횋̓�i�g���iX��hM�H����+>1r=3X�~\�M�{Ŗ䔺GH
���ް{�tt%�y��@~��`��c]�F?0��Ѧ�iN��_��]	��u�8�IHbj��1C�$�(���n8�"�sX�Ȅ�u	�&�,x�D�������1�os�z���J[N>u⺽��J"n�`p���x�L�сX|��=�.��K֥BS/6.��/�r��0�}+/��K�����jW����㜔;I���f�Wn%�Y�k'=3q��C 涐��g���!Z��-� �4&ĩ_ʙ>Q�m�}�6:�B����*9��$��0ЧU�A<:�+je�W��p��6�A\{2"����1�~�In�.��-H��`茅�S��=��8�p	q�F1p��u����$_��g�!O2�}N�n�����V�h7ن��ZW:8a�T�g��Y�{x<�Nxې��,��rmb�J}B����Nϰ;�f���j���O��$H#Q���.��.��������Ι�1ˑ�kr����1�J4?M����;�qDژ!c�[�ڙB���KvT"ҿ�	��?fy������7,Ζ�������$ʬ4��*�si@�Lv��=޲N���8$���d�7���\�l*�jE^_�q�iFĉyt�e[N�'� ��:�is\-tc�B��E ��U�u;���ߪɕ�,̈́j�Շ1��1�,�C$��G(�Fي.��CM�2�h��oxj~���Z<a�/�Yx��B69����X.��Vka�ȰUm<�Ü�vp$�k�{�����ޣC�J�Z�b`uޑ�� ��%�8w��!ϓ��x�P\y���\����$����i8����mH��{��Ge=2�(1W�K��''#T�Y��& ��/������c��^Y��	� �1�ܾ�e�5��o��"k�~,���4��S�x��Ug�8
R�]bPFu�_��z �g��)�*���0�9H�rme�%��櫤b���sݮ�(�u���ekd�,�d>OZ�����Έ*a��g�^�,>��W��L�W�L���	��8Dr� �'L�3˭u2�L��E(�%#hv"![8n��u8mJ�H�Rq:z��<�zN�`|U����W$�п�&"���?���>��� �!���k�mr�{9C]ۋ�+7p�i�����&l|7���� ;`�T�d���q��E���녱b����b�L쓥�=��h�R �	A�}����v��QR��3^����O,d�m+��
�����jos�a�	������K�?�E��� �b�{]�Y������x}�6q���Lu�1ؒH����B.���N9���f4��tpȝzc�9	V��u�#GK+��O�VF�D�d]T��4 �3�!��Ф�@ְ?�����=�fΊcY~��`#<�a7��}s�l7��aa�6�.C�*��%{��$#mT�螈k�U�Zq��/��u����J��B�3�2�)i�E�I��Z3��;��"&tܠ�:�\�;s;7ah:���meA��!'�ɏAQ�%r��MO���?���z�u���ƙ�X���̗.4WG���ߍ�IӍVD
y�v]wƥU.�ЪkT�K&s��|���L`"�^�`U%%~OIјz�9&_�==- ��#�/ʅws���0�Q�`�ח|���IƄ����ኧ������gD�f[/���E`5���)T\9�ؒ��&�.��W�bUQ�;�ج��(�͌��98O�	�R���[���=L4v�E��!�CNj5����>ȓk㙸�&yMn���Z��l����t�3��	�[�C�(����m���.@i���9&���s��|��e�H�<jpǱ���GPo�[䨄8jW�	��Xs�"�@�72�Ô�pO�_�0A�ع YT�w_��g�U�Ȳ�� <�ѕt�&E������������G���N������7B`3�C�K{�%��Ug� +d��ȮT�H��<����6�L��`s�v����r"���J.;7�e=�����E񟆮���� Q�t�މcե��3V�������)?�Ql�����;�,�:M�Z���������j~�b_"�E~������4���r�Y�(6����`�[�Q�W-�$�[� �u����B0L�2Jo�oz@b�L~�R�m޼9�G� j)*�b�_�;Z�{|g�F{Ш�2+w����Mw��|��j�P�c9���F�5���E���V �j�b�T�C\r�oX~�;l�z_�?! ��^EXa�}��n՜/����� �(��<Zn]:	CdE)'2Y%&��]��5��:@�����Ӹ����Oۣ�B����Z|(M�**?<�lJ8���
m�(>�9�x�t$7�룱��^�����7y������Hg����g��R>��� ����:<(������r�IIҊ��ğ�k�TOq�u�N��_��<�-6���]�l(�px�L	�we���F��K�d�9�����x��6���:��C���n\rD��F�=V���?y�˙	�m'ۼT�*,d�;�w������)��f5*�KÏn���SP�[pm��O�?��J��u�#�h#����ʘF/X��*Ӿ���.�>���8Z���=CsKJ��v�����[����Yy{��1�[p����U����%����*gsK���@��_;e'�~�����Z�����$��G�q����ь���z�C�4��^��RY��������!y�vt�>���@��ҏ9O)1��h�'맿�QL�B���b.���d�E�9���ƈ�|�-�\������#�U�d�~[�g$��&ۑ5��Y�˷�Y�Y
��
���̂���2�����ל��i�%؛a��PQ��C�G���)���S�T���"��B�/��r��(o`3�R����}��;���Y@Bl�Z�'�~�_��%M�ԗ���J�χ'+�2�B�		�Fm��7��̦�.��[��{(�]�=f��e7s�2�M�3o���S��M����3���c��?I�wU�$�>pW���AO� Ea5c��U����D)v��b��K"�B��w��<� ����U��9��Ǌ�W"!N�q{����x+-�����u�� �7�!����˼hJK1�T�g	p�c��r�<������[��&����
��y�*Q.u�G�i��]����g�b4I��ؓ6�5�L3�qz��Ql�{�P8��vǼ�"�B�� �h�H�=��(G��qe��X��	{)��ı���s��
,�?��ฃ[xc�pi�.����O�y�γ�;��*���L�4�l8E�y93�i�S�blI�>�¼�0DC`�8��c�GN}����i+!)q�	/�p���\���f�P iv}U�gc�{_�ٕ"0�w��աC�b(��ڭ V����S���#��R%����7�-)���:��4��)����Wf�*BW-9����P�Y0lv�6t���篛��8�0�h�����P��R��7��5�C)�pkˑx]����<�I@|\Z�G[e� '3�lٿ��֢3^�ew�x�� �Sms�o$� U���F:����)�a��8��J6`'�\gq���� �jߥ���@f��7��s�����-'vR�o� P�y����Ҵ\�8��RD�ߝ�J"ibmZK\x, za�M���'D�a�(�AyE;��p
@[��0| ��дÙYG���kz�u��X��D"�.(�x�v�(e8S�P�ې3�D�|Z� 5�5,}����;��	Z���ߗ.� <zOz�@���0�*������m�����[�\jE�:���o^�@7��3y��Jt��)e㭓X�%��E�(��_QO�6�a4��:�?��'��3��Nf����O�\��FwP�'$��_x�����)����c�T�U�f��ba�wY�͙\�p�N�m� �LS�� ��E�lİ�ɻ{������8T�b�Wa�ѝt��},��a��hl+�H#O�s�e�}�@L�m��=$�lF�/�8G�p�1�B��`�ĭ�UF��.i�9��+��,��;�Z�:���'Y�x3�)m�$PǑ��R����ф��=�H�@hd\���Wc��I?��><��S�q��g�X�l �7�]�q6L�3��O�xM�]������rQxi���*2��A�}�y��Ʉ8lH���X"�gP�����g��F�w]`%&���B�;vPxwȫ�4*�< P�3�m��up��<����`�`��V�`���x��?�Դ���ˈ?��q
�j=�������(�����U�+�����Is͖���¹�3 Ѧ���x�N��-H4J0�_kd��2�Fe� ݀����s�K��t
���2m��Q��a-�۹-K�B�So�)��D��x�j�#��ڨڋ���)�b�A��M����x�v�=V�4���B�!����/������ǽ�^r���$��Qk�6?�rp� v ���r�Ze8�{�*�`7_�S����˗^�G�M�@8�[��F�ْگ:�%h@�!�5Z�1٤�/��,9֚�Sc��T{ �ug���g�]�4��Jt�*6f@FQ��9�7E���(+ɡ��J��'^�����_r��/�Lݤ�g�hJ�8ۉ�*|	Z]���	�%&���- J"W�+t��������"R��9�%�MN���1�,1>Y4�p)E�q�Cqe�8��􌏸���"ƥh��
�[z=��']��Wa��v�ۉC�-��<���"Rkp��o9Fd)0�"w�m !X�@n��CnɏY^�*"����iQ���mgo�7�y!�1��eŎ��Lt79|��Rh��.��} �|�4�Bl����u=���}���d���D�q&�M��4=�Yf(x��{�����Q��e�)��K��d_'�%���j�����#����D�O�RZ�����@��2׆�x���1+�>C]j��ҏ�z�'.-����th��a��c^ca��Iߊ����a�� ï��񙌗GhrO!�\�l�0��T6����t�/�B-����F��t�F�>h��^N���{�m��M��ʼ\ʆU:M��wܕ�Уr!>vS6���V��$ W�r�4ƹV�V�<���h�^�-�S�����v/:� ��
��3��]�Z�ط���3�ů��M9����ڽ�����!�!0:H���i���� �r�s�T��gH,8�O�����?+�/@�#�ʇBp%��mH�̯c���]�Y�爘���u��*�R��������J\,㵉�n�䔻J$	|F�/$i�����
b��̔�K<>|��V� ��I�#�&f�Y�dZ�����~XC�Z	�=
Ø;V|�Beu]d�C�Q@�W԰�8Z��A�y��V70�ɉ���~������-�E*Q���y.�%��;i�Ԙ{�$��y���&��ֆg	q�1�*�cy_m��wMR�zYt�Lwe\��;=�W���Z87�5�5἟�)�s	��l��ǉԍ�e��UZ�D�s�('�����@�5'
%�*���PE�`Z�^�<�8�T5�BSI�*��yL���`�����2X2ܮ���T����{o���կ�e	$�W��>a>b��ola��.���s�$S�M{����hD��lW�͖QRCCB���&��ǇH��^�t�^j������8���9�4�s8Gpy�"�m�UĿ����!k���5&5�r�x��mk"2s)-�{~��B,Op��_�	!����%��*B�ct��CN<Ť�����e��`�zp{%�x��.��'0��O���(K��cP���C�==��s��:�m�|���D�4ؒ���H+0��R|H�u��$ʬwՑq~���1i�%>e���+K$�-i�D�_qfu�O�kye�P�,�FrTw_�����
nrNzq�"S�@xUa�����O�1�F�i6фG7a�Y�����/΍Y�.ϝr�*��ȩ�*��w��V�~���ߘ�6���v���/�^O .iVG>r�}蕆挨�8#5�
EƜ�
���2��i� 	?�������`2s��q=3	��عv/��*m�is��� ɍ�tGT�B	4SI��O��^���n��8�G�`ŀ7d2�pbߺ�i;�!��E�n�I�F�/`Oz�(t��q���q�A���Brt�͐���������l��Ow%r�`�_N�V��-��}*/ ��7��{��׽/z�*U4��?U�Xɔ	��dQ0���> �c�D
���Q��1+0�s\�m��%T:�y�\ ���-<�J
,[u�JQd�?M/cݟ��v���e��}d�ط=1sQ�� ����{ꮞ�dխ�*T+�~�O��;��=(i����&D��=�E��\�ɱ���������|�U�t�
X'�><e$��!K4}�*#�.�J���\�N��z; �8�fqt^v���cߺ6�Z��4�������߄~�
[}����H�ž7�#YOŗ ��	[A�O�h��j�m�����+�s�4��5���1�&@R 5���;ui�ka�˵$l`�����I�#G�o�'!���C��ۥeM\+���������ֱ��D���4�J���B�b�r��roE-�fR�qߞwiMp�S~�3q��<&r��Ǚg��ͻ<����H*v>��-%��W�*x@�L�R��nx��3^Y���mn��#���yt�R�F��u7���>��y�OVР�袏��3?"�j*V��zv����mQ���,���Db�����=��E�Z�. ORp}KR����:kH#L��V�2+5ȝT�h��P�p��Ϧ���;�|�OMA�D����܍V���xdb裊7y�/�m����F�Jq9�ف�p-)��m��@(��`� ߧ�`;2�!��1�2�'�tb�[uQ*��y����n���U�r�iY����bB��B�3�1�w��hY/@E�%b��D�W����n;^'7�4UJT�X�K�E�~�M�+c��^,�@������֣�@�CL�څN���d�>Z!����Bgoߝ�N}M��Fk���0�&��UQKI���{v��0< A�s]љ�������b�s�	}�|��
�bHdO��:��Յ�8Ň\���%4N��/��h�\=�
g�Է�j3)��t�n�gV���X�3��Z	���ќ-s)Ή�����L�,9������#�[�
�uAW���Fd����W�����ݽ���^6�g���П��#�,Z4�]Q��A�iӈ�RTb����^��7�CNe ��Ћzs�g���k3�I�@-��Ԣ�����PU��7���e�%x�zh;�4��j_rۖ��\��D���bSY��� ��(z���qt�9�wF��{aOi+��Tg���ӱ���=�ܐiF�[�u+���M��]{����2:�x���(��O��͍�L>��*�]�ʷ�2�;���F�-þ�e��-z�g\�v�n������]�7�"|��l����
����]��=���*WOg�}���d�Dn,�f�	IռL�b6����)�΅Ӊ.ݸ:�>��jk�DG��o�����{��)i�h�t&���~t�u�h��o�jwW���LU���-2�%�iOs�h�=�w��L{x�
�]��vqW��e�qj����R)����3�$����(��Σb���g3�r���c6�A2ya�U6��`9�
�(�ڨ �NOl�-FX�yC	kь��CB hz�N�wV�%�a�xׇr�{��r}0�xL�)�Uj�Ug�Y�M�+�oN������u��/��:�7İL���4uV�]����BQ�]�Q���R
��؉�`H'x���:�@�^�D�i�=�I����VPq� ɉ�`dڷ�hB�����qf�O���ի�6nQA��nJ�c�&�y\%p0��}Tͯ�̻
�Vf��\Ѥ�����U�ݢm�_��fJY��T*:�2P��"ӛ���j!K
)��ŦHje=�3�8F�`Q/$�n������2*�l�V
=���^�X���A�E�x�H���H(a�<�,�o`��h�/�����y�ҹ`��є��1+t �����`�u�Vw*�.�TY��`23��m_���g�k����q��̅>����Q��Ч�r���҅t��3�$f�C)�z�5��@��+��g�Y��|�h�r���
��*8�Q6�UPy��
`G/e����)s��U�H��i�ܮ�T@�
��Q��*L��.�J\G����Y���J��/!�)�6~����:�;W�<��_���"~i�֭�ߍ�o$�ؗw��.�a�JO�^���⪎��$�nHa�؛
^��m�~��w)���� \�����ZOɚ@����<aC�O�_��2G�����[!���k�&��F�t��wҧ^l��a��S���{��[9��j�7�)a�9L�e���Ы�k*��[4�� �F��6�!�Bv\���f�������e�7 =|��ҁbu��HS�	%��j��<�2���\e\��V|:_ .�����@�B���6�&�#�]�@p�Қ-�8�`+L�jb���^���N����2���@��΢A�)�`Zn�����ۂ�汯�_���"K��	�`�����|�So���s9�l�'1�nY՛KY�K>����b�U����l,��*_J��9��͑�F1z �+1�k햦Q�`�4i�s'��/`"��P�_>��F}��! ��Dz���2��#뎏�Q���y��L9Y��;0P���+$H�zj�,%7���0(5J(Wÿ|��̲V�%���G��ʜT޼O=�����P����I1�I�Z�5��@�v�E��}�%��;��9��~�J�d��T�
q��8-|A7�K��a�Xl������Φ'9��bI��	-�hi,n��'mpȝ���\Y<f��&��J��
<����/�S)�g�ByRN�փ#|=�b�.��Z�W1�U��J¬^��ɿ�Hpf��=�_���r�u���D�������j����ʴ'VR��!���y��4�����⋺({��rI�-��!�A�B�̍2Πt�HmD%�����1��,ӏ.�+_X�����ڳ�!����鄸bŬ�:��3b��g����S���$M!'���m���EǑ���ϿTnҼ��9��y]Qѫ��u�0YD���L�֓L�ʭ�U81���I�w��['x`�Y*�z���}�[a�(��N2�[�`�
��dW{ ���4�[>s(o)���|�I�������e����,r�|�CݾB� �D�N���(p�9H���f��ϰ_�L��x&fա W�gI{�q�*�8��f�ht��6�����k[�lx��3)3�eob}���AUA��<�����ۓ��7�t��������q��?Q1���� |]�+�Z���E��<� &ڥ. �iP�Ʒ|̱w��J���|�\���+�b����ş����Xܓ^�7mE�u��S���}<$��������bX�4�^~�B�E����{2n�jQR Ҫ��]#$ǐ�]VWG��*m-O�Ȟ�)y��C ��+��"�w_B'̨?�d�I��)H�8���b����FFA�׃�vw���Na��Z\�@�[��Q��N�^��<��<Y���m=\Y���t�2#n���5�C�A�[yuJ�$kGf�~�Rt�����]d���}K}�����+�/�m���y@i:�@j	��lqz��Oq��m\���� ���P�x����ϼ)(%iwo����g��b�o��Ί�M(��7��f&(�| �s(�jB�
<��1P�g���՘��q�N�D+��oY��!H>7d=�� �����}Af�����ӥ�Gk����`|L$�WӘ�?x\x3Ԯ�����Q��Sɤg
)��c�d�tT��B��߂��Lpɞ�vA8�z��Jʮ͝�9��J�x���=����:{���}u��$��-�W5/��.z�
ڛK�J���8�\K+�	���U���v��0�fS�c���q\����� lo!u��.��2��jXӝ���QS�{�꽊���:�pb�k��h�W�`t�[t�͔��1�*P0dl�>m���\�+0ziU��lܴ��nzۡa/>�q�^�3O���N�$
*o8es8����3�u�8�[c���
��#ܙ�1)�re�����!��0�VzKGx���T�_G��Z<@��p���V��T>�eLE�퇲��T5�Z��v�Jn���^�$𤠷�c�sT���4qp�>�]R8�m'$�:��;*�q�¢�dD���$>E���]Ag8�1M�jP�����uMm����^���	�L����Qs�F=��z�y�29�ӥ�ٿh�,aﯽ�����m�v��"� h��&��K(w�>p��Ep[�ϐc� �� W%�J�˻!,��;��k�zw�~Ц�lE#�/�[(�����.A��yr.o�NU<*e1s;b��S`@)U'J����ۻmD�M��5�	j(-��@Q��9��n�좄-�*;��1�Ѕ�]ۍ)P�� 
��+p�|f2�=C�|�)��� �dL���f���i�����>���*��_�r�V��#��Ug�S�b���1=[��5��Ή�4j����,BC�h�8��[]�� �&u!07J�mz7��v�&���{��;� �W@���:�r�(�m��7��Ҟr�+n�	:�4��D}\V��o͍6�JH��K�����^٬�@P�/�)��[���ߕOX�����$d�&�fa���&Lj!�s���s9������AQ��~�HU�s8eF;�	$e�玉2��[�z7��7<�|��A�Z�pɯ�=��gv�����7y ���9���]\�/샅�`�U���튊��wC�6u�����lp�22�;o�EukvJ�엋I�B�o��[� ��o`��/��z�[��j��D��v�2*H�*{*`������b���n��r� ���=-�f�x�Y�I����.�	k3\�+���k�?j����-�fL�D�&|��!C�& �à���Ou g�k� ��R����*pе�\�8@t;�*��m#����@.H	z����L��(�Nu��&�����3���6�J��
fDT"y�p"w7n@{d���¶��6c�È�����2�sq��2�*�j�<%���?N/J�ZI��<\Q���.=PTCk������#�r�S��4Z�Ta)ÿL�3��Q��P��-Ht��R��L�h��N���)�[��HY�2�P�n�0�N.E�z!\��@�|�OG#K��l����4һ��r�� ��t~C����')���Q�O�����AӼ��c=���E����/L�7�K%�A�u��~�}���ld9��C�����{��y��O�)�|�NN�ɇ;�4�'0$����=~��n�qy���ƍi���a� ̇��<vb*�ޜgP��������C�=4����~�sY�Z���.�;�lfK��dr�E0Yt7RY_m���6�����-&�V�<�.a���}[7x��6��~�ԣc#>WR��<J�MYW�t����F�)��+ΡG`zKӷI���O�ܒ�a��T#n�-º�Jg�V����vh�P�!���G�Q�
��q;_��^�F~4�i�a�w�_#q474�9*>o�ׇ���� Kj�6z�D|do{������%l:�v��fGm��t��j�Z;ԯYb�vnB_����
�V7�g�Vr<����'(F$b�A�v��dvY9�=��Y9)�06� ��gu��"�h	lx�v��ĭ��&��y�V�:*by*vs4F������H�?�P�����Rg5Z�.�Q�C�Pg�p359t�YF� }��Q���sK��r}�+e"z��)Z<S���b�[UP]��)Y˅w���a{�D�#X�K�dA�`6&��,4y'�V�h�h#QڂW�䓐�6��ޙD�ʀF/L�`	�R�_�}�o��`T"��6�$���z
�»��۬T8SXҦu�EJ𺥎!B:�ر݋%'��6�Ŝ�d-\�KA��g��L�ؖa���x��e�*�����󻧿@M�X��dX6	�kQ�!��!�"c�i��O�2)D��W�� �%mպ�Ϗ�U�G��iZ%�p�����} �n�Rs3�i�ӝ"�h�=}1V�� ����0���{C�����(�Du���(�SW<^�A�X�i�	6{�&&
�K�R9�P��/���0�y&�_�dO��'c��� �P?�J(����m"S�F<��X�	�9ʠ	��N�(=��7y��S>���_���Ƅǂ�o��h����]��b��{NC�i������M^��(E��Hա�X�n��m�ڒ]�7�D��]��,��J,$����˳&��
�!�,Q$�*�� �@*[s�qBS�4�^#5��ah�����_Κ}��F�*qɁ+?j���&�J���CO�Y�r��, ���O�W���*�{׾�U�y'?�=��������a���Eo��s�X$�'��u���[楼ZA"��R�t�$�$+��Ҷr�[��͟=�Ln(��^eB�(�#}2Ҫ_+g�gig#�p[���z��ҏ3FDMW�:�`��fڋ���.�E��q@;w'��_�T�T��/����K���%U{�_p�|�a:	�nj��U�1����� �"\���_.���6Y�M��{�<{JĲxr���.R�4�D���r�kP�r�$fT��1K1ǊQ/T>``�DM�8\��������W���,U3���j�0���L�2����t����P��^D�������<�.]�jt`Ɲ��ęev�%CU��} _���ȃ��8��� �6V��iL77���|g[C�lX����ǘq��)�����0Y���v� ��9dV^���,i���z�0�Q�IJ�s�nk�O����L$�����/�H� �2����CbE����$A��wPAA.UԚf���O���" �)�����/YD'^͙ʀ�����xr��?����i^�4N #��~;�y�x�P�H.b�QN�Z�X�BT�XV�npJ���,)C��KF��a	1�#r�R����c*�2�u�>��^z�4�q��6���}k59Q�@�̯��i��7p��������/���"%��_=����
��	�x)�����O�*8��>[�`����J��+��\[^\M{_�0����rF,㼠��H1��2[Wsc4&*�ɭ%��x���fhY���>��n�!Q��Z$(A�;C)L��'j~�[��s���W^�m���ut�(N�ϫ�hF��`(�+��{�Zi��e���U^mk݀3�)��X��A�n�2)ru�!le�R�mV�C m��k/-�N���P�t�`�#�]�U������K7[�\.Jwi��� hYD�Y�@���&���� �՜!�
��O����=k�{���)��N۫�5_�<�G9\He=R�_CN��	Aec�8S�:L���]&..�
�m�suG��.&8���y�����5�m3d@̄y�U����g�G�K������7`GΎ({��ɛ��6��q_���⩠�P�����0oQ��(�A�؈NŚ~�m�mÛ<�)��P���v�4�r� +(ݺ�!�/�����s��?��in�t���&֛��Ѹ�3�'���I4�����h��-j�֘$*?bۂ4:I��isՕ�|�>�2�Z%tГ E�EM��	�벨�����̰fK����:�q��2)�8a�\ԉu>����M'(��5N�I�lڟ����$��ۺ�_�ʯ��ha'��߫ŶPI'�R-�4DU
*�a�}�ҕ�R���knIlcf>)p�� *���|�3.�`a�M�����єCmDb�p���N��*K�+l�>�a�(�E���,�M)�:0%W�l�&}�H��K�F�7>�ϫze����I1)�.�򤀁۾�+�Z�Ջi`{�E�uu�r��#�K��R�jL�2����O�W���/��Pod 8�z0�.eδ��Ӕ�C�-F{�M���q}o����ȫ�r�ڸ���Ү1 
!�̒�J��R����"U�u������)�����B��jq�ж*o�V�TU{�7�u�Ò�u~<j-���hZ#<3ޛ�w%���ϖ-�2�r��nS6�����޿�A[p��cBٔ~��mk`'cj?g��A�a��o�:��ssv�B��ϥ�1��u��%���j�k��\��a�9�`i�%~��Ϲ�U�+(?QPbD��wE���n�%���$K�E��=�z�_Ȅ����D�Q�/�ր�]1�9�[��Mɤܝ\�P��ksa�ɦ�!<薬Fc�K�:�2��?�B����'Ew0ɂY�{���ɮ$��1<G-fh�Q�1G�T�G|�#xb�Δp�Q�������]���'ns��:�����_�Y�D������o��U6���hl��qL!���)A��䋬V�҅�䇐G�[`��w�kұ3�ÑinDEs�t�cZ��p�;��i=�"=��V�TR@��	Vm�K�e�|��ܷa������+7< �������:��?���Y���� �D���6~Ny�Nɯ������]�����%6e�E*��Q� #��!z\�i��� �d�߆A0M2�J�m,�3�ǀ�s�ԓ��3�X�hQ]^�k�k [*abp�t�V��#�3X�aʵ<���NN�R�)�h82�'B���� ��6�]'��"��u_�������m�w�_�3Ѿ�ʸ�]wWqK�"�2��>��v���La��?��R����q}I*�o:������P�	g�XV������-,d�T���~�mŅ��m�B�l�T�斧�?+�����D�
M�{�A�m���Ab���Y��kh�@ӗ'�L!D����Ƕ�����0ɸ>���s��Q�}ԃ�Cj�����!"3/�P��Ȳ��*��^�K�	�:QF1%T2U�V:X;�ߨ �|��f"�CIGa)���hă�/3�����6��d6�̑�̱�S�%3D�^0�A|P�x|u{z4��?���Ɨ���u�m*�'�����Ug�PXj	����3f=З&vbߡ���_&��#�_����c��H��0�g�9����k-tŜaCArBbU�M�QY<�-0����1�*N��,�_��3�Wm=2t��N�6���W]�6���Gz��Ўj
`)ZL��spVwY�'���#�;������o65F�� 6�$�ڟ�"z�)@
Z/\�#�?B�`V>�R��-X�$����u]�L��D�Qo�rR��6�3���C��B��P)粧�E���<��`���f��:+S�G8Q�BL^Ί"x�NA���h��"]�������\�jZt�/{�?��tfB��EĲr��n\���_\�*1�vr��wͤq�zv�����m&�k�9��,�.�*��D���N��y�N�-@��#����Z"6��X��`���y�(�#]'�m
%�!��Ԡ������7�%������f;�����֒G���D���l#P�q�����f�m�+|�N���$�z�}��v�>J�<�wi��ߦ�h����[����)��#?z67�
ĵ�״�a�D��g�o���E� �+�3h���P���f�^;���Ym,Fwd���a�ɩ�-����v��˥d�I��Jm��������:����"�kax$!��(�eFN��2���m���<�4ҋƮ�uez�n|>��W$���1�� ;��G�IU�j�!lۧ9>�S�J�����,�	�c��ڡYr�z,^��H�/�L8Z<"�,�A�n�*���������ƿ+�}����Z!��� �: ��i���ٗ<�[�4�䯙��'�hO4�D4�wkͲ1���X���:1(���7����BN�7YrR�c7���f�as����H��|F�~[�hf�v&����,�����qK$����T��1���w"KI{�ش̦����[<��o��V��������+�� �9a`�(�+�~�#)uD�`��� U��-�{{��=�[t�ű�돞�ed�I��m�"��]H'7��d�T@�	�x$g��O�^d��s�3T��f!���W�f����TO9G[q�M�d�uն�����R��VU��D��������\�(jτS�}ߧE#̑M/hC:^h�$��K�x�l�o�t_��=�b���m�	vB_�*��G�^�k�q(�$�����-ҍ!q���Y:r���Vw`}!�F��5m�B�!P�~��p5�Mݛ��e�:z�%�ŀ8k�<������*�{�w5�	�;ť*��ۂ�����o�)�/2��<7>��/C�C������!��O� 
\x�)�-���&i���t�l=�]�#����Ӳn���;�߿��V����,Ҷ����x-H��G����'�#�n�+��.F������X��{�������]Z-%���]Ě��f"���O�z��[�'8��]R�a�04̦��	w-��s�����hA:<��C�(ɸ��#����X��Z S��$��<s�����3���#�W��Х�))�y����9JIÞ�>*�j�3|_2?���\MևTڐ��(��Al y��8�^CFs�W��b���R7�cl��b����-�� ηz����#��h�SP�PڨA~��,�6�N-	�`S�t��{���,MvF_�%����ܗ�P��"�<�� !���ۻ�{�<q�|a �x�/اx��R�{��(��wjm���B!�ɵ�8��Q���85&��<z�(CG7Aj5���>m�&�#��M��F�:�A�<8�
���'��O��S��J�b3�^~���<�d�9�[?�r��xb����A�ޔ�}��l��w����Zv���Tw�y�E%}�!�s��lB�e�mЎ�09Sm1�?��F<�&%I��$��)i�l�:�'�r��{ܻv&���
����������C�e'=�e4e�����7�q��x�3g��s��AQ#I����h^�1*Ќ�Zr%D08$0�C�M׿B#%Or3!HK�h�����^:��"���`��/z᭢,�,z�j��]��_d-�o��M�V�qQ˞�y��X���*����][0��;`�%�-�iMWء�����;cy�v�o'�u��px�1�P������a��H+m:��������6}�1uS���Gl�ŷ�������78Ok��cjI3�`#����]��_��^i��j��u�/<|�����P�If�?�d��6��Y�E��⇨F�