��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{Ns�ȭ��+{do�;��F�0�Sa�K!�f�gԜ��s�\!1��!F�wX{,!��p�V��&a9��*���O �a~0��r����0�kn$�K�%�'��N�,]x	�f?SPfS�~�F��yȗ�4��j*q�w�n˪Kr��|��k��E�a�]gq���YEB���4�����<�G���#z5-T�c���S@C�$��0�x.T[�j]h2Z9
�d��;�2J�"�5W�7�BH��!0g.�{'��O��x�3e\��B��T͈)��L�����pb�'������n�Od��jT:�"��P�;��Oy�_5	�hU��r	+����J�ry�<?�^������;��(f���	�4;�u@Ejph�gb���BZ^��p�d�/\���9w�?����s���X]x@�1�R�q�F�l��ڜc�c�ʨ#���O䥽{zF��Q�bD͗TImƝ1��:ۃI����ӟqµ����v.P�Y������g�g��N��mm�De���CK��H!����ӟ��"�o�l߀5'1���eC6HS��@7ȳ���2�����Be����� B�N��p1��g�������(�	My���0�)ĕ�^|5�KR�����&��L��^蒾ۣ��L�Im���W}V��D2`u�V�D���)I�{����7��C�?�)����8kx�/�"7�~ǟ_��if�Rb��esT�g焅wl�_���U�&Ҷy������G.��"?)^]��'��NE6y�ϱ�Qc7��7��7���q�kF� �-\-i*���u��ђ����F��.�py,9��(��iç2�
db�ܓ0'�@a�l@��AH搻�V�p�(<�����^�1���o���i��ٌ6>W��^��������� �ah�@që�(�bO�)<� �w(�;���m������7�e
"���>}L��@�C�p�?�����6�M,�b��7y^����,�J���:)Z��>m��D��8zcYŉD �V�u�^}5z���L�k4���8Kd ������v���XWIL����F�����e���~�� ��HLT�]��H�̇�e/8���-�޴�1�Ȉ��KoH��pH.�n�����ʥJ,M�i�`�L[t���1sc���t�W�w���݊�.V�d5b��@_V6���j/M(t�M��͓B������L��1č)9��#tݜauTO�Ω���<D��4�|"�MC��B �h~n�P��ۤB�c�fexMK��=W�Iު�O��.K�)T �D��^t�/��+�����sP�����4i̙�j�LX����!QW�:�i�Ũ��� B��bV��!��Z�8'��{k���4��U�7@�t@vѦfj���+6+��E�D�aNN$�YP���dH�r�/���&�.0+c;~�7��ा|����B�����0�5��"��i�P8ޝ���	�]W���w��~��N�
�ǿ n2|N���M�^�.����;����S��睵r<l2l�[OL�Z<��|������N?�#3�c�����܀��X́��9��~kkk�ν�S������pDS_�4NVI�X뻍��J�,�ce��n3�����)lZ�֝�s��h�$�55{8��2?J>�q4c�4f���L.�aڨ�	S\\\�cpƻ�W@,�+M��er5�(sfݼ��;k�wK<�E�fW\/�X^�K�ޫb�h�;bٟ�>h������"���M/
[��,�F�����[�]gB��^9� A���I�k~�{�������S�i�yYc_Q�N�oӬ���4�:��G���^�
�qX�F�[����j R\m�y2\�����>fY9a#�w66t׳>���-�����W�%�����(��T;x/���F���� ���drр����9~��}A4<��SF�t)<��2�;�Յ���� Fg�H����[	��}���!�{Dޮ^���G�[sH��Oj��G<I�+?2W�iX�᫣��{:l��}{T?v�wO�>�F�+��:a���f��M�N$"q���.�3�6e�0_���0+��b����	u�^�*�����X`��o�q�P�TV����ab�R��c�����cf���J�s�ɡ�̳�Ft�����@��p��d����B0�eK�C�.�7�>��.�V�~���l�O�+��\r]���8�n�C���r(��7�=��SD�^I��9�o!�|�/%k��n)�O���+iñ��S��v�p�9�4H�PWu�h����a�����'r?./�ΗӂA��Q��i��9j�6�_��M��E=��8pL}��j°�U���*�������GF*d$@�*ۺ�E� �Ո�A��Xwc�����z��<*�J�9]�!��Ҙ�) ���L��Y��Ed��uVI��?s���ּ8pL4��S��D��#����y��\!��y&P�d���޻`���8}vzb1+�R������gu�C̏N�V �3���Ir�B����<ND!����Ӱ�ӽL�=�O��ҐZ��i��W��<Y$� Ѧ[h��^�a����E ק6/i�1ӶWgt��C�������lcZ{U�F��f�G��Vȯ� ��W/���|I�Q�m��S�����q4�zC�c"$��6�Ka�{�N��Stn�1#����C��1����U�?���|�UY�X�XR��f��_���V��.�{��̥�C�P=u4;��P�:��ߊ��������7I��/��>�-Y.�k.�U4����,�G�d-P�Q5�2U�PlvS�2,;21+e�W��j�1y
�) lS鿀�Xttqp�&TQR�>��GD#���
. �4�a��A�����4S�9w
�H-��H7M(�0>ҩ�"U2��%�9�Jr�,��4��$s(�s}T���,v�࣒�\I@�;��.L"�s�����O�z�~�}Zc��&���@O��bW�V�����=,�X�ܒ�������h�G����)���yB�� �wo8 ���Ҕ�8o*���\Z��~�)�Sc��%e�"����}<�H>�A�&�@������Sn��������X���`��q� 9��X(�f��"��i�"*$��K��7{�%jT<�آ�AE�f��UCN XZ�P���y�\�.�+��[��v��ߟ�*$�2�Z��T.@>��֙n�Y����ŋ��*�� ʭc�]��e����J��L���^NV�d�
F����#�E諷hH<�ú�̽�yG�:��<�����G�S�F���> �M--�����8�.P{�0�s�h�5L���,�	YQ���!�Ey��@�������֘�F��ċD�(�3�oU�Dj�C��D��V�[�Xk��G{��L�O|u��H���N5qG�Z��R��%�,����P�m`�!%;zX����Vx\��W���"��q:-w�D�TZ8��v"7�}ab�'���U����*��.�[WD���@3�ጆ��VO�f���U�=�N/�8�=�>.r���Y�ΠP����s�N(Um�Kd3��E�_�h#7�eZ�+�M�߬��t�D�.Uu�k����3�+T9kZ*�x�'�Ŏr��L�é	&;sm�ǜ�u���<��t£jy+}�Ie81HߌԓGx�?�L�J�pB&޺*�@TΚ[�陫��L^J����➷wԁ�j�vEo�"��&m�q�
1}%2�=}�0�P(#i���u'ƿA0���\����W�:M࿄ی�{��|����sq��v��b؟�n&%�΁>?l�_��J��g��S4��W �]���U��,s�U��*^Ӭ�A�#w���/o�2���:x�N��	��O�V0A˽�k���[#<�GΩ��O�<�8Q���'^"�,)�{H��򛆪J�����Ayy��\�RoT�{�*���t���U�!�iȗ��n��ً~�v˕�-?������^�b.\��ˈ>#�CC�+�+_!_殅T�^�24�uSP�"$D{�￘��(�$��;�Th���eE%ۥ�[n#���+{g8[��%�9�~�t���X.B��[�J�����$� ���Vz�V��u9wN��'�������;Q��i�Z׏�=&/�>C���$�������80#M���`�x��F�^�}*_ԭ*{eL(ʪx?>o�X��L�\�L�~��	|�?�/���Z#���]��ՄN��ۖ�D����3�XS*	�w�����c�y{Y���z��w��AΗ�o�!dw��g��-�o���P��P�%��J2�_/�}���ܡ�H� ��Ɍ�F�<�f��h��;���n�S���<��YY���8^~ʖ�-�+�a���j��.�pc+-A���U=<͕���8pa�]#@"�dg"4| �*�̺:������ 8%��)|[�Tmg΃-+lX��Z�_%�	�b
g�y`I\P��Q{�4���6Zr��!:�7ޤ#�Ѩx��iؒ%�>J\OGd�0ߎ-+@�ވ<��܆�1óļL@��>?s�́��
�d$_�9���C;e͝�h6ۆg�����%�L#c8�C���L��2�^=c�-�\f=��tZ^�ƪ���g��+9����W�W�����i(�����+H��	���_���	s�^!X�	J;+Z�oo��x&�c�ci��F���*Kb��	�����GZ�7�D��/��9��畻��2�9��;+�*�� �E��X���M�<��,�@�������Q	��)} GGd�;M��2n��dZ{/�����;6"?�g�5.	�(̷�Orc(|�DL:r�N击���y����1��
�e��� � �*/��דY��g^:W:��	�^`�2����Ԇb��%���E�=K�*�)����u鵒21{?��)�p1��I���Q�Z���^{R$��j_N���4�`-�[&<��pFN@� @���f��>���zjbC��1[�5-��CN�imB�F�i��[{�K�Ea~��ϯ���t�0O��:Q�S4)��OQ�W��A���0|	�Dd��˻��}�1���ս0�	��*���ysѿeiƲ��a"�fmJqm��6�!�