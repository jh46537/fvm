��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)����\VH7�d��6����]�:	JȾc�ޢG��q�@�(�0E�+���N�)|�~?�|�1E��vv�(K ���'#�X,�ӊ�tJ����weo�����t	A�\����]�*��H�<'���c�k:2�D�¥I��P�����+�;���^�~���A�Ipg%��b��4�$J�Z�,�NɕG}I����S��OO	3�A�K�{�@]�(��-����ː�~����rU.�w>�V��S�����C��C�E�J�7;�!��]�	Sɮ��8�WnI��H �w�3���N&~ ڛu��EX�(����;&����'�]on�L#2���0�G&����c���*�_����o����k���M6Ϳ�`�ʄm^bU�2�����w�g�r��U���*g���BԵ�Q|�~D�wHZ�y �� P�\#8��a!�-��'c��s�݊:J�*>�	iSw!�3e��x���W?H�>Ң�#�O�$3�3J� �m4We1I�k��(�7��� �t�P��p�-k~���67�;����!�3z��(p�KI	���Y�Q�;ȩu�����3�?t��BV��,ꜻR�vAyLC�n��m�s9�.�jXfV�-e��i�P����3�b%<Q���y�ft�>�S!�p�P�PL�SKˈ�uKK�H�܆�E�`�3:�����=���U��ŝ���=Bc5���J�ª�dP҇��^�S?�jd�:��l��;xi]�)d�;�Q4���r�_��zx�7:�"B�!���f�� c�b�_���Y��>�~�2z�ϙ��!���@���'v���:�ڋn��6Ef妵9�@�m���o�xc�ԡ_&�����U@�u�l9�7�0�����O��:>FE��g��^�uA=	N_���J���2�_(��5癑=f)�?�]V%;KV���0Bn)i�'<�G/�U%5,xa <h�M
����Z�~��ƀlg�|!��6A������L9���?�הI��?
�ְ=��f��������p��8�ˆ�{�m���`�1��n �Y�CF��E��z0!���EԳ��������]�4��w5A��n|>�k`�s
A�XX��&����:m�|�]���2��o�ژ���4�nŬn�S%�8Tm��v*ނ�y�s.,n<�
^�
�0'e��JvȬ�N<m�w��Bm�>�/�z%�
I�����axL�w薏hA&eF��/���,��XM6$�͘�'��B귅F�)\R>��P�4��ڡ��`�,.���:��O�:f:�y�R�Y���S;=�M��,u?��σ�j��{$�b�A-S "i�Y̡��Iϡ��3G�I�e>�h� ��!L�Y�_D^	T��A��[s�C��l[�n���F1��_���_�d��|TJ�����c�zM����U�|�}D��Y�AV;,,Ҏ(���':�Ǳ��Ãቻˣ���^�`������M��3}��e��[5�)�N����=B�)Zf�-���eBNƢo�L򀱗 e�Y QX�)-V��6�P�ꝎB���W��{ސQF�����B�\�O��O���b@53	�����v��_{�U<5؅�h�������^��Qu\.R�ѝ���gY�.#��,p�0�|�_��b�'�w]6^�A�C� �.����ҜEKH�|wF[�A2�:?h�9�+R)�x 7�AfR)���P�hߘ�j�y�kWT�47���n앉�����~���Q�s9�������WY�\���G��$~�-��f:��D�b�kK�"�˷,����ͱN����"Mh-ŗ;r�|�}�&���a��0�~��LP3������_f�CS�KO�}�W~:�����f��U%Y$s ���;b��x�ŎQ
W����:�MWr"~*-)��g%�f�JB�6%P��OMH��cȩ�$�봼�D n���?��tĨ��M�C������G="͵��OuǹeP�.ds7�DiwAO/�c:�ؖ�� �4���I�Y���ry�|��0�i|,�H_�'�ʾ�wKΑ��ꯣ9H9�{��ɴϣ-�a�:�C+t6D����g?&�x_�o~���.�|����0r��pV�A���grD0	��-�r�/��2-T)t{�uJ�yd���J^D�w��;ZU�Dq��{&?��%���K-��(ſ���ѓj�E� &����,����:����b+�YL/���خ�(`JX� f�y�<)@�I?k�e|�����d���{�|�ƭ��Tr��gw*ts<VR�d/��_�iO���cM�I)�g�	Ӎl���L!������{�Up�?�z/g�NeB�#��b�-��@9!n
��Yy��O��Iӈ�A�� �Q��$���~�524$���Ln| \����Qt�G<�����ޥ}U�)S�t��᫅=l&j���n�9%+I�W�0�;���/�(V@�6�������o�WR��O��~e����QD��h�Y�#��htg����l��C���)?B��-�P�g�ׄ��z��SW���q�,S�;ϸ���n�T����PN�<U��7�����ó� ��IF�dP�j���	c��E����x�8��qĴvuIN�>�v�R��1r��@Il��b�_,� ~˷�I!�⟍��iV�&�ҳK�WCe0` IĎ1�8�6&�<��� ��z�����3n�xV?�� ��wL����V��w�O=Aoh�Uu%�O��C�%B�a��m_cH�Pt���K*��$�EO���r��B_���Q5e8R�Bc�������|�GQ�a��h�ޭ����@�v�@�����L��Vߨ���h���s<���˕t%�un�cÝf���=s�Y�Vo�i�=�/#w�<��t�g�f�j��k����QQ���a�(�G��.a��u�	��O��M}�>��Pm3��O�fЊ��'�����L���(�\�a��H�)F}ļ���x)�����Y��[�Z�Pw�7���5"s<s�ݖA�����)ٶ�iH"O�
"A��h�&�Z�&�%�!�Pf��b�LS�U�>�L)���~�(*w��ѯW�)��Y�R��pi��ʛ�2����҆ۻ|��}�]C;������N%�2���������'a|.��W��}���&C���ؚ�|���F�c��ʴ�z��B6��};e �G�������O��� �8�D�O0)�¢��ѫv��9AJ�.,����1�y�Lc!�����)$��*���&�,�9����8�F?H���ؖ@�E���}�B5L�����(��m���Xt�����W4�ȹsd��J���Ϩ[~�\dyl��JN��bڣ�;��/{�dhK��B���;
8����
�.��^�\T_W�D������aR{18P���|4��vx�۱l��:��yXD���9Q��p7���qm\�|?ĝ���lT���Y�� <
�t]��֯_�3Ğ,⻒X��z�"Gh�3_ �F<K�F�$��j��MM��j��j��S_�g�P��f�*<��vS"�߅�\����;nz��}�Hѩ�Tܬm)1.�d�J��UP��2�p"��츀hnfZ������A�{(BB���������%�,�&�~\4�^�����~��0S9�P�Vh��~��=�נ_rf["<���'���Y����K�IYl7/\����}2�w�CQ3�9Y�@��b0�-2�1���pP�qO)pO�O,�0����O��OZ�N�2�q��YG�[D?ì�T��+��;�r�2��b;Sa��D���A�/��43��,���%j�@��?��
�#������2��+)w�(�Q },ъ��\�Do2��EU�Z��7��+��&�����t��Y�~��1���:E�i�"��H?;�4��h<�m�)J������ �J���(f<p#�������"tD+B��r�oPk��w������(6Ec��g��[޹&5-���K�Qp^J���I�P�C8�5o�"^!�@O7����:q�0=3b�>��cŅ% �ŭ3$��&G����ෟ�U�jDrY�Bh����M��.�H�h:f��缶�_�/��Н��$�]��y��E�Kj�%�w�p�Q!���l_v$Hc�*d"c�D|c;�h�J+ ȱ[����[�3e��oc��'*6v<����Y�/������&^���t9�ofW�����8(�	2��*�5�.����4��8\k"�ݡ���{-���:>��8��v
r�I�F*\�#����WiM�M)��+B6�H�q��0R^H,�1}�O%�=yZ��Od+�M��Ou��$��� �^��Ifr(*�%�vҨ���p�L�������:6
 �{�2Z5+Ll$g�|�[�(� TB��V¯��%d��Av� 
HOY��:K:���8'k&�(a��4I�(W�mt�- ���6C��)v����$7_���B�v�M���*	��E����+���'>N��؋�z�|-�v]P#������t��J��sLǝ)AA����hH�]��A7(]��^�%�Tep�7Xuӥ45B�y�M����f�D�r
C~���[��B��C�mKB�R�G�DQώ׫�F��mz^]F�����P��n���-��,��c��i�,���Q��x4�s8⭖�Smh���%�D�
Z`���T��o�\�0��3Y	�7��ʍ�eW�>3���&ځP�.�q�~��ʩ�p��5�e����T����(
9�<�jlԒ���t��QL��� ��.'T_�Y��U�~��Mq������+N<�)��DҒ��F�f�^4���s+'�:D�*�׋vґWY�7�};Vd�f���7'y�wǀ�}L�Vp�@z���ݜ���˖���H*��	��X���\�'�~��P\I��Fi�Ţ�~F�EuJ�$�ȫ���#�Z^J�IS�6� E�/��_$�����^ٶт���dB�	�]㵁r��W;]�=��G���6�nNJ�'���`�1��X���g����$l;��.U�H�i,�2NE-|#�cx��m���GF�����vVl���\�����I�i2%��VXXj�KU��y�:|��^���n��"h����l�C2�>֥����z��0!g9LI��%��LB�<���I�/���GIW�����&V�)�W>&�!t�%�ep7�`S��c6�cE��*Y��S�2���P�l�р>S>�Z�r��/����E��1D9A��	�Iqh����:�V���<��$3�ت�2^��~X�(�3�<]Y�$�|��bG�f^?G� 3��ވ`�syXG�F��7cD�F���Ƕ=Va+\�&��Y�b%�J�U��Q��E�@��*�X���8o�{�zɡ�#��O��'�mJ}������F�<�7br�ߴ��'��-`���puU���_�ΤYlQ/f�`6]��E��͒5�;�K�	������Rn���X��W`�Z�*���?h�M|�o��G�}JV�����囁��ƕ�k��S�8��׈�W�p�I� ���t X��낔K�9$��%��W��_ټ2�̷9�8��Y�����~9�XVK�
*��ô�od�6���1--Φ�c������XU�9�sY1Vn �iƷ�R�CV�U���[.��uD�Y��H �BB\�~��L��CBF�\<v��Um�ZM*�\{���XFc�m�$��F�݌ϭ`5g��-��9�6��U��������S�����g�M'�&ַ�K
u
r����j5v� ��%�+Y�T�>��#��5l���F�~w��Ou�g��3��+�g��>�-7 ici�m�q���:����/xD����2��\���
r����/��H���+B$���mdp���Mv��47$��o�Ue1㷑���/P�r C/2b4r��n������7���`G{
����[o��@*?)���ڡy����_�+K���η�[u}�w] X)��ڐFM�-(..�M��B6	w`]�]�\Qz����X!�#5�Fg��5�j���$s�v;ݵ�Rq�x�X
�ì��O����px�]\`��%X�0���HK7MvSͥ7Xu�;rDfN����㽜W��,�����p���!r�o��������!%g��	���R��o՝�?}�-l�ە���Q�1߉/���θ<[J��/�36�&�,֤�3+@K�]n��:R5O�D��KyAb;��օ�"��OS�☖b���]+Զ����3�.���TC�/�7K��R�Q|pW\ր+u�4���^��OӖ�{Ɗ�n�ڴiJ��h
�?p� vP]|�8��(���(��1�kԽ���j�_%j����xZ۠TF�u��F>ag��G��jqS�U��訨�/ܮ��y�$�~�
���ٸ��`���ឨ�>N�=�ǜ�(k���;��ĳ#v�J�\t�\���`��."&U��&�����q�'�Ix		�vhѤ���'s�ܬ�P ��+0�F��nY�'XB}f��\��̞h��nb�����d�1�Ԁ�y��1��zck0@�U������X �zX���5�|�])	Ǌ�#�ho���7u�v,������fX	:�g�Ёg�k����	��!$d"q-���'���U� �X6$:�j�'�<�QZ,�Q,�r-�g�x�֥]1"���<��u��B0x��"5�����x�X��#î-*����}&�Q�c�En��I��K���{��k�d}����{
%I�z�l�� �zO��rPz�����,�)� ��U���_�C'�'O�Da�!�b3�e�;˄��%���*��.�ZɈj��ߍ��+�Pk���p�e`n�T����� D�_ @5�0��SbQ
��I8��]U/��x�J��0�\5%!x�N���y_�$����x]�8�����:�rܾ-�o�':�9��u#���H���4�j��f�	����sNDԷ<"J&�.���z�5��H	4�ޅs���;�(�<O���W�$�����i�"6�[d�>�d�~�������p��������f��>�p��0]�?0����1�+�����)L'�8Z>��]�aoJ�"�r<���OV:�����>�},�4~�Bףt�5���w6�f�N�ڙ`��)���I��$?��[LDz�
�)�O���d��8�/�wx����%-S�k7�pY?#[O]�ED����{rդ�:,A���b�B�q�����!,�y�5�8|R��ڙ�6 :�~����Ϫjg-Cs7c��G�&Jc(���e��ш�_�}W{)9�҄�h���h.�hk�񩫲���tt�K=�+5�j�HA�u(b�\d�$0�_`©�O4CT
��m���M��9��uxJ�C��Y��*o�	��'o|J�y�%%����y���br��&���s�?|l#�N�+�F�V���D�r�e���. [�� �?� C�Ql�%6j�e��e���?4��\���rE�ÚB���T����蚤,۰�� Ym[V~x��_׈�+fG�a�7��L���ZA����+�~2jl��Y賸?ȷ����\�j�@+%��)Oj#X�/�� �P��$���ҳ?_�,K����HEl0?j��G����?ʷ٤l趢C]�6ڈgsQ�^���R��	�����
<z��yt��ZI�����6�8�4��������A:HG����[�Hn�ɭP�A�h|��I��nRK�S��f�|�7X�a F���ZgV;��0r�D1]>!zB�w�%Ėz��l�,�bL��E����� �'��x�j�=R}@��d��_�m1��]����b��Rى�(�7YG����2�������R��e!�{9�����;���K��:M߼��fT���
6���G��T�-�v��&��#bY^bYnæ���%�*�Ϗ��_����[}�i�ڎ�F==Ƚ��i��zp�^`x	��W�Ro�@���91j��L%��9����kb�ٮ�ēы��e�"z�����lV�=���?��9-�7dw�-<�VC��6�c�)�oaʣ&)����|�
��}H�O���+�̦��~Q�����K5��.����>ڄ�S'�]A��1��B�_�&����6מ��G��U7��s�r�����y%�N�Z�������LKД�?������8CkZ��?���]Ԥ����(�ӁH�j���|E+X�a�� )�H���8�T�v��RY��t�#��[;3,|�u7[�g����.��H�9�ҫc@$��zT�����U�6{x"�
�7l���Sw�C��I����|�;ˎ�&��������RC�o�\fdM! �!2�V^�̖�̰���F��.S	�JtLl"�k��������se�$�[)ȸ�b?T����t�&���A*s�^���}��NF`�2�L���S��{��<��S�<}/$D�T����=�޺�''�9��q�D��c��#��=N����Llb�H��������\��u5⍳\�����?�g:<Ϫ%�%�i~���e��3��\[q��q�ɸ,S�9��X�G�t��OKD�&?�l�h�*��R_`�j3c�0Zq~���Shh�X������� 膝zfB���x}����Oߎ���I ��d2���r�qX��b/����$lC$����QY�BݕuB��|ڲT��_�o���`O[1)��m�	��^��-O���L�1�k�L#τL�ku��C�v��2�^ЋnQ�=�Kc�h3�:�����گ�DrOp��Q��l�1�'֦?c���JD�7j3]���7ً�I9R-�sT��/	xl��'�.�������s�t����7���^�.�=QI?i���K��4�3P����[l��.��ά��r�'�K���,c���T��dk�Ԁ)W��05\4AS��{|��<�&��g������?+�`҅��a�p�G
b���D���&?�)O�#苅�;�4��%"��i]������ɟ$�Rs�PMM�'#��ɏ�k�ܰ���N���	�����R�l���fd ̏z߾�,�1���$�FG[Iш`9���'������>��A�S���t���?����<�F��*]�{^{H�h���<���j�M���5�`�|�'��'�Q�L�Q߁m��%��Uu�h�d�t����{�)x��&;?q1[w�m5��G�%@�([�LFf�qy,YXM��Q�u�5[2��6��.l����Ɉ�
���#M��	]��l�����)�J������Q�6X�� �ܵ�&�����Zg�O\���,��^���]]XL���i�%�k	���(Ҩ��@ϳJ��cd�������J�j����e4�`�1����"\�5��hkо�G��y��(�]3'�T����J���H\����e�/���c���~����=Aut�q{m����O����vU�8�ۄ�/�F�"ξ�=#�xdA���~��cSʯyY�""+[�h;1��������0��g�A�G�;ze�W\Q';Dk�\�  J��ѳ!n]8)��!�Y�B"Y�e��>����ш�0<:�0C;��t@�@�aX������\oz�;3����0��kF��'�o�Uzc`��Z��D[D�8�n�ı���g�X	�t�="�t^�����a��^�_�A����:.Kbzp��0|�ڥ�A�X�7�ƥ��]l�%!��-�a)#�|s�Aww1�`��o�	��"���J�}�~Y����&=�]�dK��@Ժ�f�N��7M�d�V3j����g�1����(\���7s*��C,g�[���۴PӚ�7����v���L�N���
�m���j��*�>j�_L=_��< M�Ad���������͞����52�>�M\�m������o�U��Ւ�/�/#�u�����;dזv@﶐����bPv͓��-�Q&EA��~