��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<�Qҽ�������v+u��/�T����i�Y�h>d���7	&��m|�hK�#U�7QA�7�P^��N�џK7d���7sT����A�c�58�8�{r{���@&;Z��̶�HS�#4��ᐔ	���i��nm4YiE���[b�L��!��&�Ei$��ζ��y=�R�Ԅ��[����H��i\h��e�2c1L6V�5^��m3��C��i�Z%f�����F �U�SZ'�ǽ��y���U�w�S�m�ABC���!sQ�o���y��Ss����(Tԡ$���XZqn�q]�Ң:l{g�+�	�i����"��N�s�N��*Q�M�|��l�C!�-a�OM�}X
q����!CY�M�0/�5��u�&�4ɘ1$��@�EK�闧�^v��ѯ8OE� _/㊚[|a��,}���(�l�$4풫�$�U�����)<�;ekN֪W̝�[�Ȩ�T��.Ht ��:�2�~�д�P��>r���e-�j��/7������\��G��L���<��G_k��o�A�����NF�=Kr��n�[�Y:����ŧZt���Ke0PY���[k�����Ѥ� �v�T����s�O`B�Ϟ�|�/)5+ץ��rHNprR�@��:?�%KI�0w� ����"'ǿ�F���;��)D+:ڵD�;�{�3*W���2@�B�|k�.e|0�c��G�D�G.��S����_B<K�L!�	y�I=�?���smՎ��ƝK���9=�D��G��|z_D���ᄅNU(08����k(��O*Ѝ����%������L�\�c@
�K�9/�KC�ZB���`O�����Cdە!j(��Y{���RXYd����������$���hQ*]�&������ �Ć�U٩��g�ܘ]�����jC
k���nS��N�����Յ7�9_,8�b|�H@�ba�e\�?���Ȥ�4��zQ�?�ȕ�����ĢI^sn8�`��=6������:'�'\�	�k�2@���p���rZ7����N�x�*O!P��k�/�
iI�]�\�9�w���Z�$�i��#u���
�H�;� J1��`PB�F���Ks�����<�����V�3u.��r�b���ۖ��
�r�I�^&7�m]��Y�v�����֬���zT#��͆_�%�6,6��ͼ�No�P�E���.����	�0��_�ᩳ��������]�D����|e�����rL-����E0!k�e>	��%�J!R�i�\mv	lL�R���9�N<n�x`B269j�E�����T!fq� 自�\�8S�d�82�9S��Aè��a��2�t���cu�{��|�c��g�����{�����Q2I8sFm�l���z����r-��"�v��C�}�s��9��|�c4���Q{��P3�q2��@�'�����h�y�"�f`4n�����"��8i /�~Cx�k���Q�^�(�*�I�s�qD(6��8��92�꒱|5��eӞ���Hl��$�Xb���[:J�5qTAY��_�K�ҹ/T��?@(����h�g���a?�o�|L:M��h��؞D��>�.i��$!ة-�Ļ��q�os0�7��>���K�@:��d�%I�t��)����+��}�f{-(yx��R��nȆ�ٿ9R ��>��Lf����M����3�^�+O+�0;Ԯ
�U�	�@p�3aJ+�j�gz�)b��m��ʌ���Qd�Ώ%�u\,�PT�p��O�����A
7ӖQ�I�즅cm�0}��@NG7�V��F�h���|�0���;v�g���hFA�矚;b��OJ� �c6׳t��z#���v���˸(�)Z"�{{��/T��U-�Ь�kcxt��\�R �������ܞ=d3�W���7Q��o�4�y�h��3�Pw�|1�IV_^�濵�ǡ8"�^�Ay���w^�_�B��j�L�����?���3E���(su�s�g���4��;�͏���LV�vF�����8S��m��D��øXus�ni����y7�N�*�w`b�]�8C	� �c�"�|`���������T��8�K'�P�G]�b����.�s���T]�T�;>9�VF�{P:u?���F���*ޥ�c�2��0N��)k�7�!��'4S)}V	:`ȳ�d]?�Ⴀ
:M|���T�Z&�[�'LgL���J�;�4v�Y��
B����t� r����#��!i��0�i�?��t�"+��c`ٲ�C�=�u@&�:�S ��f�7,���kc�+�f��ԯ�)?���|�4�m��d�2�n+��j(��(ZE��
d"\r}t�f-Ĩ��1,���I��	��jA+6S�,�W
3c�xH�_�ܼRA����Y��*�J�.ʟ��,����r��L�^4э��sX8�'�7��ǁp�pٕ�4�N�d0$���(a&Zt�1��;	�]� 7����QT���گ�87E��b	�y3��d���<Ac��ɹtoV$��<�;�*қ`���Ξ˩��d�{.r�w���M��k)��j^��K�b�	����s〲:�f��l�(;�X'O� ��JN���hh��J�U�W�u8��-9S\X�s���D���L���*�hC��7�5#���z�n������GX�<e�ܗ�>/%�&���`�I�jcep��.�i���6�x�ǮN���;�X��Mݨ'�� qu�*�k�RA,)خ���;bWN����U޶����}� Iڐ�
�-@-��΀�Aw)~�K���,F}^XA��[��@.^{�n3�pt��_��)@�_%-آ��ijK.���/Q�7 Ʈ�����%%�,'N��n\1��T��-+�b�s�杨�.BdAy�MxSum1�@����u�v#������#�����Jm03iQ|�kQDU�9+��x˨`P���,6��{��pw����|�a�v�T�G��g�וĽ��#0�岑F��l~�1<XJ�Dq��L�UT�V���_�)�y�!����g�^��!��/�Cޱó)�!'� ä��,ۚ���U	Q�.�.��Þ��滃7Q��3W�D54t���:N�'�&�Hʤ�����Ո�7.�Q2r2�Gs�VG4��hw�����Ğ��I�X����!�)�AI5�+i���$=]ͣ��	b�=�0�̔f������]~s ̪l��̊Pu��_��E>��DK �ղ#ܞ�W%?�,�Մ��T�Dm��Su�ޣ�"����?]`zu���Ҋ.#�4��0���f\�,���-����H�'�e����b�@ VB<�t!�m'��Ꟍ~jy0RuފUt���Y�S���iE��9�GEw��{&�:�"��JHY-�1��coNd�G8zu�E�t�!�$>����@.S�E�2l�2�fȦ���F�)3�Ke�f)]��U�f1�ޫ0ӟZ���F� �ӆ<)�y"�����}O:��
�0Łq�,{�y��prF>�FX+.���:̛a'���>������!��C˕���)�$���c�Aj;�4J��A�O��$/i�`,GB�ʚ&nY���jLK�h�Q����7��#�Ư��rE@���[=�p��n��)�Yu�)�R���s�2��P/n;�Xr��:�%?n�O<?F��-Q�R��*[���������.a�`�kר�A���1��<tGsk��Є%J]�\�+]L;� ���x���b<����a�2
'���R��ǵ]UU f��P]i�OX�Q���ܠZq���}a7enM�*��n�5_`����)"�G�ˁfgMe�WꇊJ�[��h�+1��ԩ�c6U2��M^�uh:��q
�@�����ٞ���������R��:lvӗ��6A��ſ�J���nb��
��
��=�a~��+�A�R�����*H�'�W�o�"ڰ��ݡ/�08�*�z��V9&xtD_΍�z ��(/U��̄�d��>%Ň�K"���4�kTn++�:�A�� :�F�=cF�B]@}��n���V���=MȠk�!R����V���.�Ӛ��Xk�k�w�m��O��Cg�A�1��VrǛ�i�=	hhh�l:���&�P�ygۚ2��9 �t�k��̈́�a�7��63as�>?��^sH��:��_�2V1Dn]��i�Y�#ьڋ2�X?=-%�I��s^�BDO;%��X�z��ܪ��I1)�������K��77���1;��M�%<�a������ڻ	p4jv��u_�/�,_���b�E���@��+��;�އ��duJ!��y�I}��$�o��āV'Hv]p ��(��@i�F�C��N�l#��wl0Xb��<����}_�N��ආd�����[���2���4mi��v��G����G>�>W��An᠍���~R���S7d��U���jT7� �誀#`)�_�m�� �Pe�ŶT"��r������_@d�]���#��WF(4É��l�:q����IM�:�/B�c��M@�MFݽ�o�*F�����J��ڥh���%V��.QT}h\��0�B	;����O?���
�V|�-?	'���eZ=�xz����1�<Q����حik�[��٤��\XJ�1�Q��`�b�ӛ�{E��`�]�S��R�.�$�=p��F
1ԯ �#+;��i�مT�N�*T?]"F2uϓ����"5$�fA����?����f�;+�0���mR6"Q�Q}R.��3�%/��$���= F������e}^�	��n�wf��.*���!�s^����P7�%���>�?���ٷbCج�=D�b5�8+����~|���	cφ���Xcp�x�6�I�2�ڋ���ңц��,�ާ±���� ���$TQ;,�%}%��s���\������7����нgY�*��11�8�e�KO�H PTd���U \y'�����>=�RMڔ�w5�,b��k���Ԧ�p^�S9L���|)=C�B��ka������ja���:��[Q ��X�4]�����E�?�]� Y�vX�.��!M����6���p����)��9�r��=��w��!p ��%�a�U&XD���L����şT"�@�4�LS$a`Y���]if�F��X�yP�I�3XZB'���2�	!{�'2��>�VZZ�dS�h#~wgS�+���I1�Xq���9,&��D�x��y�w���L[�o�z}t�ϼ�@�k�8VBA���Ӥ��.X4Z����eV����� ��e�s�����兕��UFyMƔ
�����4�UO�M���dww�'O 6������m?ǧ���/���c�'�g����)4�!�F�|6��-�ev�򐙘
ƟOPfl,y����h�t����%��U��V�������u��2k���9��������st�ז�V���E>����8�!<Y�O��@X�U��x�b��!{?c������݇��-���<3��Q�����]zI��up�U�u͐7�7�=�K�(w��4�(���y����-������d�G����L��aZ{ls�iCT�:�<a'*�E���4~3�&��G���3�a���kG5߆�*�h6������;{�u�p���@���A�_�hu�y�:�Q7�~�����&*�+v�c�צL�0P�V�9C��X��u��G��;"6d�:Q��-�of�CO'tB}"��P~����E2�h���9�9��!a�I=�.�n�Q����]�Js�����"�:HS�n���񴲟�jǯh=���|S�=��G��2h����e�N{(�5�I���C�/�\�s�S����u�U���Q��-Ӏ�>QH��h��U�"��Fk{uCL6�S��\��"�Վ��X����;��p�W�"$�3w���̕��)Q�O���0��W<��
u�UK��0���ֳ>
(X0#���y�?���w~��3?AQ=�SA�!�Ϩ��1�A�0o��5��IDԫ�=��"W���6���&�iҸUCDK1Vb�ja5���2�����q���AV���v�HT�(�����	��gÐ�8�}�s�E�U����W�LA�j�?�� >!�J�o����g%�WǦ�Q�O������8�>��~T�y��,4��ѐǗ>�ux��-xlf�n�/�T?�_�@�[��i]�35��\J�+j���jm�b�T�+��A���wȑv��>%���i.�:j�C�DG2�k����6w�x7�{B�$���N�.����6]C@c���@�+=���}RަS�A�l�+�+�<��mHa�1�=�����N�1��K5�(����$x�*�3p���,���
fnC��a��7�z��o�m�Z�2�GǞ]gS?�D|�[s�2iٗ�D��]��3F_��,�~!�^��l�����`� �LdZ�h�����$Kß'�1��q��("�=ve�D���'���3Ru*�h@������TT��@�K-�����n2�Vh���B�ؾ�0K�zE�4�C�v }��l>�y�ZRb�ﺧ��;�� ������~F�)�:@�
R�w�����8��z6�+t7Y}��#�(v��SL3>ÚG�h��橭�Ժ6#�t�<B�M~9H��=�p�]�[�<�P�B��h�����!����A��@����4dX�e�XX9[(W��T(V¸�:YpSJ���Xu���|l�N&j$*�z������<Ӑ����+��D)cp����N�^���fu�x��W?Db����)(.�}22�?	g��y�k�����w��+PK?dƨ�ʘ�XI����Z�;������BaE��׼�%���uˎ� \��g6�l����_���Ccz��!��G���n����V��������J���Z���ZPM�'��"��׫��E�00R@{˰��lͳ?�_�%K��h�� Ӵ�N�e}B�z3�QVw�m��W��(Q5!P�������\���^ޫ�WLw��&���NbT fK+�f�d2��%�l �;���.Dm2���8&�%�����ԟ,۳�E��cr&�Qr��g0�&�9�)�1��{��p!��IEAMω}ڴ�U�s�P�%ڕ���&�"W�rA��<k���RWx5`z�E
�]k�S����^%!�T� $1d�gvh
z�y�OLa�pAO�ឲ�;�q��5��j�ASd"z�+�s;1��ߒ��'ig�j���0�ʅ_���U�w�X��,wg�J��;�"�0>���(>��aZ����N��1~$�*3�����d�8�</��'-�eE��~!\��֞�t�|�|��}�p�cc�Y���p�r}Z[��Ŝ�zu�}Ӆ�K�F����y�1KY �m��
���� X�'֟�Ġr)�qL����"m����I�}�Љ&Io��k�#P�ٺ�P]�6���$��bb�⟅U6�FT�!�	"2�Jv=m\mڗ{�zh���֢%��xM�j�G��rR}ŧ��σ�E�H	_�_$2��m����P�Ɉ'�'ъ V��g�Dje���ޣb�f^���h�OGN*9J���J	��ػCv��i��7�N�gz���=�M_�{
��j�M���Բe���k������d�'�?�"V}cgcb6&�;�zw�#
(��^d�#�Mv��*�Ow{�!X�K�-�����`��(��;Ȱ���R5 �p:�梮����c墦A�,���z�)�U#�V��ͨ����ڮ?�� ��-P$�K���ZS֑Z��T1y�-oM В"�񶲟z2n��1	�b.�"x�[t=H3j�)��
=���-�p���
�>@�N�E
&n'���՛EBL�˻�������8���o�b�Q�_H�2��s���Q1A��#pR���,�h�\�5?1+嗀����CS�����`��"5�GŜ&�Yį#c�軵jm@��Dy2y;�J�[�H/�qۂ�9ֿ�"���0Ko!�Kdh�p5��3�Zp�*�[�R.T@J��70+��a���[��C�O���NJ����8����O&iwUu6'|6QS+=;u�n��ı@�����x!c2��>�,:�J$�%o��Z&�6�t�~�����qU<��鿋$n5՟5:i�ܱ��kpD�g��d{�
�˓�^����?��q�~@�jZm�m
�|��ɹbL1�S�k�>2Ǐ���13�	���s
@jX��@��?��Fu*��xy�WC�$�������Z!ɡ�s�A�2~=L���G��o<9f&�k֝�a�K�!+��=���"�o0'�i6�u����|�/������|A^ �V�2D)�Df���ѦI�^E��<kş<^�	y��n�1���FrՁ��̒�x���#
G`�*I�M"�ûF8�`"��S ��8.*��C>M�g�A��DG�@��m���G�J"G�I{� �jM.c(�#lAf~ύj�[�a����[S��b��"�ѧI��s�ugwv��Ʒ��Hbux��-OΎ��L�*y��ʡ��lb �-��� �N\\H���#�g]�?O���{�s'�)<��w��骬�F%�҅�6��fa�Of|f�V�gk}�"zUc���b?��".�$L̲���{�0�.g�Ꭻ	��?1�$��Z�B�<4V������Pbf�Kg�'��d�(3���ϴ�E$��ݠ1C�6�Y�Z�%ȶ.��-hN��q��ㅽ��@����%�7_Z�jԨҒ�K���"+38;����.sT��S1�����N�j�S`fC�u���k��
���*(�+c�������T1S���1U4#��/�PƝ���{�θ� �/&�s����b+<�����W�YpK�=Ӊ -���6��/�Q.������6 -������
�m��#�_x��\2>ە��"j�D&�R��e0���U��9H~^խ̡�X�1&2Q��2��7z�`�7Β�+4W�a?�d�BE|RZz�r�!8/��jf�/�f ���yđe����,�[X`�u���zua[1��t�<�T�s9/����r�s����1dj[9�+5PW���E�LO�}+s�ڐ�UB��a��$b���� ��)��C�l�ˋŌ��ܟ���Û�,������>�lJ�8��WL���@���Y��on���hc��Բn��-��:��e@"i����u}��u�����fr�'��yfD�]�6��T�TmC�.gm�C^%]�c��^B<�֛Z�����gd2Bq��ي1Ub�M��g{��K#��G-��X6>��;�@��ƸB�}8���Ju4�:A&�ױ]"=�狻��Fe��4�r�8�����Vvp�;v��U���2^��~M��QM&y��w<�c�|r;�M͗�s& f{.�Y4J���?/���Ȍ�G��ᶂ۠����f�Z=�;{Ԣ�E������)����E�����lsx�#>	{`��xBpuLG ���AP�[N����FHu�:wK�~[��Bao���ud=;3�����ͬ-H� ��u�~�,n�V�]
�2���mK<���U1�x�ˈ۪��a'�-�����Z�B�Ƥl�<��)7���W۷����C��S`��*]!���Y�;l�t?\����<Pm�7+�E�r(8
^��畗k%������|+6,�d��͟Po�ic��1�-t�py
�q�y�=B�?C���_��V�T��K��[��|���I^I�V:���|�/�P�:Qr{ �wDx F�\'YM�!涔i��	v+�.1�Q�:�s���p���p6�Ϟ���I���\_�8��	��h�D��4�5�v�N�\zP.đ�������&5uI�\LV��
zџ�X1��@�h]L�R�&GZsS/UB��,6n�UH_��i,�?C�覀�خ��U�B�"�3S�ߺ<��>t�&Yg��G���ӝ����7��%WF���oV�'���e>����,�/�b�7��:,WlȺ#���C���'�N~ �!s��e��	|��.�9�y��a:@�Z߇X������3�ĩK�4�_�&¢�������'�b����p��"��_r��TGsI���&�ڴ^[>�ypN��Q��r��D�L3S�yw([�/I�b�����@�4����<J|�����nt2UtZ2e�J��4�ES��?����(g��E��%���to#&�J���!݋?o������0.0��7��+io���<�Y���J�]��<T����XpuE6��ۡCY�l3N�*
7�y�
�
���2wKҲQ%K�)���u�vWSW{��q�@�>Po�u��h�4X�{�]���̜O�ᠴhk] y�b
U��҈�a��}EuX'�RM]k�|�I�!'�&�E8�VP`hћkm�vV��9Ը��A����(2���F;"��x^ɯ���������Y%�����Q��ݚ�aEo�� ��uEX��S�`G՗l\��_<��&Y��$���li�K�E�N�3�Ix�_���B=��B�O3�j��a�9K����-KX�	����9�5;�w�96�j
�N��]n��"AYD̺���#/b� ZE���������F�����(�[�V3�G�s�$S�$<!���.���a�����F���d5�mЋ�t5��Tc�
�b-m��#�C�	k{r�4����:�W�A��o���JU\�/ ��;ZN{)��.Y�E[\������}VaY��-���4�Om��kIt��q�X����'Up��[��Y��zR�Լ쎼�C��52#,4D�G��{�jvGj��\�?�lS4�џo9Op�5��⑗^��D�"���-�������_���z���e�f|#-�g)�<�马6�b��` cyIv�*m��?Ph���gm>����W��y��{��� sĦS�N����l1���h�z��x���S9�%B���t����*�S	w.�6�apn����7n���b����W(��tZ��v��a5��G0M�b� r��^��i�ؓ��Kw��Y�ǟc�2Hq�w���m� BU�Q|_}�z�d�R'��)F���ʱII�5���=�[��3�ڕҔ�D'��M���k�8Mj���'�݈�~{�)����U��'��S�@�H�����J�i�Y��[mBK߄%��݄6�;��k߰��(������}"���
�,.�!t�������ܾ���p}qI�`����L	.fu�$��e�Ձb�[<g.X}�QK�c
��I���惪k�����֯Z���fC<7�$p�w��%��{T!�!jW�ܟ7^�Q{�P�0�=�?��\7Dk3��"��08����AS'9�Y����O4����5|v��C��b�!�VbJ�Y��o^��ߓdM(�B<E��8;j����E'9�*���q^����
�A9����7<�R�3>zE�}��\x:�]C�%�?a�+����������'�\�k��뢱nZ�Y
[ޡ�'^�d�E�<�ؐi
�ѥ~k)�Z%���ⵄ�Ԅ�R1|�cq��悃��T*�8��h���_^�H�����/�0��"��c�#	�໥��]��I�'8CSv���(��?`*Y�^��L`'F;��et��A����G��-y������j�����0A��*cpB��������:K�@Sm�\N����h��	M���7��ܝl]�)��j�
�_ݤ���لz&����<Sժ�	�T�e뮌�]J���P�C� ���Z�5���_�xB�������� ��$��=�t4�{�	,]rF&Ƀ�Lϟxt�����l~&���݇��m@�pK�6�SfzI�]Y-���j�*��a�� Z`03L���@�ג���w�=�&J���8��O�ٖ�L�{�mr~�X�#N7�xN������~��#[b���3�0D��?N�������tҥb�\�پ���%��J�|ѧ#�J��Z�#��Az��kɩ��e᧊��"cp�*?�,Fi�"|ΪX��{n S��-j$J�7s�ۜ.��&���6�+�L�6ӟ���C�*���
}`V���+��y�O����y�
��BjC�F߽7�b�	��)+V�z�#*h̒抬��s�`�z�*v�*/{ǟ�4܈L��Y�KN�$�"�������0��.�gM��}�~���ꝦłZQ���$����>4Q�q�A-2��1J�\�k��!��b@����:�� q�+�K��SE�X�J��_�L��g�d�U�!�age�L\r�M]�V8�նz������80�Ҥ51iY�(H�\ɨ�w�|X�o�5��I��*��}Z�dj��VE��#���c�#�^c\�4-��Z<�*�*-�{�9/���@���
�+d7I�CCιODVk�4��<�P[f�����]��W�j�|�īayd�����}��[�O9�����Q�bƠ��]��v����u&�`{xP�4��+��!�6���IO�t�(�a�&�E�/��Q������}�u|v�=U��/�l�ܧ	�e͉��Ĺ�~J�N�����\���q9K�׃+���p��W��W-�$�\��HK��r�[k�1����1[
�됰{��@c���0�Щ�n�����dfԶDl��Gj��o~irOC��\!��zz���ÇR�B ڃC^�q|P����%�v������v�:4VT|]a��f�u��c40}`Y��t�@����Q0����Q)�3�g��SCZ2� /ZV�(9���nn�Q"y�J
[3ˌ�!n��;�Z���aV7��7h�QKM_��3���.�j^����r��5О� PC�l�T�-�C��~�:VGB2ౖ���v��ϸ��y&0�\�j�����7�������c�2�ng���B��1
���g�8n��}�9*�FT#x|�䉶�)��S�Nh����o,�����y:T����z��^�f�������F%���۸��"b^�(�����Յ���"�`f�P�5]���/��E�0����%\p��I��p/X���/J�x��<� ��A����7���I��d�_k�m��	ouS1͒�2bl��µ&����-���_�-��lK���ä�	��[{;�?�gu��(}5[ rը�c�;�+쯶E����w2�]�Z%�|
"�	��Dz�9U}Y�BP��0�X��@&�6��"PnO�2Y��R�Ū�Z#�ُܷ����  A+Z��op���z������������G�	숗M�0I�r5*���θ���U`�vؼ\$�������kf.ݼ�Dkt��,M�ŕ�B�A�h��uӒ��V0];*�9���0�����{:�Ϛ8x�w=nT�K�`�_r��?�znr[7��ڸ1��~���)��,��~��!��j��&]�U�Ea�+�1��O�+�j!��+����rZ�k2�ϫ�uSb�ݶ��D���Sc�P'�ƪu�⏅;z/�-��$�涠���p{�.,������}�e���4���BT��ʯ��g��Y�ɹ���<NH'���-����4�Շn��t�6T�	�U5���w�d���G+p�#�u�]�����-�=�7Ӗ7*:���*}1c����S�Q��-��Z��'a�R�����"j�?�Í��R�UW {A'����Zo�edZ���kޝ����:����Yw�gEM���Y�p�V#4>��[�1�"[��ʽ�&eB����ZǺ�4
 A��ekLI����%����k��e���L�`���l�:Jz���7j&��z���Ɣ*�Cj�t'X4l��A#8���v5�\y��8^��x�X|�EO�R��Us/��9��g��`ޅ�D���A�g�X���Ym�Bo���Q���_��6��B�Y�f�q�5K\�.������l+�c6b�0���-�u��������X���I��;M��ؿ*$�Ix�+NJ���R���
J� �B��+��:x�33��m�"�L�����}��C� � ��-�7"H�U���!�}���>�F i�? �)�al�v0Da W("��K��P.WiE/nKt����kT��{P�>Fe�Q�(3�&�������9o�1<�w�o���O$"_����y,�'yL7�wߧ���]ȭZ�I�p�1{:��}I��6�Xz�Le̹��p4�/�C�BFO����)�����7�%�F>�C�M��h&nv��c�*[!ц^Ǧ��.�"�<���8Z���y�7kj;>�mѮ�}��K�B�9���RŶ��U�+r{�xw���pt��:T����u�����pqjj5}
2�z��Wꈄ�Z*y�J���Y�C�F���E$r�c���R��1@lg���l*.��x�� �ec�(x��
&���ˤ��~��k�o��94��n�1��$��,+b_�.�oP&���"��1��s���$pc<��?�b\n�8���L����gp�\)�5�~����I��ڇ�S�G9�ҍC����7�ET)]�j��/Y��[<������w�=5ȥ�C
ӹ�b;>@�5*�L�� ��d&���"ng�'+��hu��s:�7YM����X�k<!���8Mm��i1�� $���j�=¸9�**�V[������`ǅ|B��� ߴ?����[	|�\�pe�t}�z	kV�5�E�i.��0���y���wr&ia.��+��l�#)�&��\�JD�%7�>m*�FW՝�?�V�`�e.�(M�(o<�9!�&��jBFp�)���k cD��X㞶��Y������[�~�l�ߟ,^ǯ����w���J/��f�h�L"��8�ye��'o�&�3���A�yΜ�E~�χP2NS����y$c�l���ъ���,� j���cPT8~8W�^�Wch5F�F�7B-���=�>�����ʜAu���0������u+ök�~<=_��(��[ryw�55]�c���@@�����N3�ĝ�0���P���	����}
���(��p�_�����Ů8�;���1>{y��5�o���5yNP<��`��*�)9
�9���z}����J�>�fPC�B��?MF��G]��r0&�`�t�Ɣ�����z�~�v2���gf�Z��3G�ӵڙU��ccKJ�x�5��r��V T�K���׈u�b��Y �%���Ֆ��<(!#�L�Ķ�1�ʓ�b��郷�Щ~Ȱ�*S�<W�!&m � Q��(2
���n�r24RRI_z!f��t�?z��v�3Z�T%p�dn�]�ϓ�c�#ˍ�=a
ʠ�e�z�l�u��|�zK��|4�a��Y��XL��� [\Q7�g"yV�w��y`+���2�@�qPj���֤|d9&�����V���+��Y���z�o.'D�7��bԶrw^K=�6o�n�(N�۶�4�HT-f����,�^���&����E��ם�DDhW� �ʫl_����s�d�t�w�]�C��S��	ua���_�3l��K��e��r�
��iJ 3S�F��Ł�+@<��&6�D9��E�ރ���,�!���7�(�k���T��@�<~�}K���y�L_<GE��ыkPd��*Q/=,-~���d�P��KoAm��d�.^6���k�_8�������
�u<ms!h�4�7i�H4F��'��;��pA