��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbg����c�i�?��t^��,�~{�q�E��	YjpA������2o&����ޛ@������g���U���0�2���.�%t6�_Ii,
c��)O�~�`�&0��5���MY�U��.n���-�,�I�K�j�0	N����0D��<�}[�]k��������#�w��4�ް���)ba�@�ʘ�btN�fށ]6��u6+����Q�����F��Iզ�������.��;K����_�GY@A��a���I�`���e�ax��ܙ���٢Φ򑖟�:v�� ~�p�w�+R=m@="se�ӭ�f�>���>>����=V�߰Ys�W���va��"�N�参���6O��S��#E�}G�2i���}.��߮���숺�����b3��x����샅��{qp�(�3�����	j�t,�)��h%ĩd�! [�ƿ�����/�D���$�u��pZ$ԏ���7*�Lr����T�Gd<�u Xȶ/�!����MCAja�K:�����6�n�V���wnS`��&_0�7x��e�hQA�
ٌ��-�Q����Cd�漾.=x�Z�괔T*V��c3�g�[	(��h�9�ѐ�����殆�q�ƍ����܁b��,[(/߃Q]��6�7SN�`��È�X$�	 N5hh�5����r=b�ٷ�ݑ��7����#2Sj�4�m��0~�������I�8�*p�Dia)\ժ�,YDF��w�+_���U�6�\�osk�^�z����R�׷�zkc^����8�\� �����J�<ҫ���֠GV)` �}��,�&3�������w�G>���Ƭҵz;�Z��/">�0[Ŵ$<�L��%>�B�(�z2I軬�2ױ�
Xo4�9��-�!=��쯸�7ņWYhg\�WCqw� 5"�c�G,�A��EE�0yu~}eҡYS�`}���WM��g�(Bv!
:-�p�j8]`1Ri�g�T6�,З������Y���|���z,횳���jo)�U�Ǥ:�q��h����%\���?>������=�%�ل��� G����3�o�H�}��a+�T���ڈ��G0Ұ����(^��gb��Nk='/Xi��W�w��(���:���Yz���_c񳊄Om�uMQ��@k�f-q�80�j/nk��K�I7��f�i�$��+թα=u=_o�v�͑ ��R�1�E�"�g���b*�����°7{�:�S�.��4Zq���*]��3�Wq��\��d{��95�G��X���r��m�-di1�!M�k
�-D��W��Vמ�6�vî'm.���e�Z�uH|���I)j��2JDg"7�?͌n�̹	�§���_�z �~�#��$x���:q@�k}y������*�>�ռ$�ۊ.��ޣ=�O��R�Ji���@W��w/X�"���8M��=�6?����R��c���o,/�uCF��Z[� L!���p|�5 �a
o���#E�$�_ZiV��P��e�В���R4;]i�9Uq��>�Ok~ct��G����O�Wee�B�O�V%j��t�$t<v?M��2��wY)m�_�����|��8�Z2hlx?��Y�ץ�������%%DP8F���2��0�w�xY%��)34~D5�}!'�T�&�{��:��r|� �,�޲��&�����E���D���[q�׸ E�G��B�xفȉm8	}q�VfYL�:���蚯�Vu�l���������L�c˵Z���X�G��K]�b^P ����%ͣ�>�ps���_�=�f��q�aZ��	$_� vg o�5�T��i��!"t�q}���H~��� wӝ,>�,��C�Q�
�B�_���H���X��u���-?^��\���N����L*�b��Z٧6�17���wh�Pʤ�і)����C�(ceOr���0ft���%[]6�9�~�bc��I_Kiʪ��o%*��R��P m�c����6���y�O�>0���*��%������_�<�?��W��B�7���ꓚ�q{���?d�a�j,�r��Ŵ'岸iJ�8���!�O@��i�u��#����G�Fc�	�\��b���3NoeYvH9�R�2�;e`Bi�͢4�xBu��=�wP�ß�V�\����.�5m�'ģ�E��P�\�mvx֟X�Q�u�W22����������筹��h��x�1!�2����L�1�
����i����օb�:RL�a�U�Wr�����y�m�Qt䁊e�A�c�����mV�*e�ڠ���ÿ�>Y�xr��U��d�;n�9�uh�y��,N;T�
��?��L�U��p�_���5����=U���b�Ș$ U��.Wngx'0�x���+1rĳ�9�JZ'�!/�g�8mO�\.�"ʹӬ��h�C�'�?p���sv�G�L��3V���kT�T&|F���mgIL��X���G����@@tBj�<ob6���i}���=��Mz�\	�$��+����v�(��8ơ��Q�[���2���V��"ʌw�W�F���Vb�����S��=��=�����e��ڍ�Ҍ���]�C�9�=�͍����t?4�ut�O��X�����������ۏ�<��)?m�)'x�E�䛯���_P�M���w8��B�����ø����k^�b��l~MO\�ڃx
�@�O0l�]}��CEq(� ۊ��
�c��-*)�{w�~�<�V!��>�{��=�Z��U��퓃]� ����c���҉�1	Fᛷ원�6�2��tm�]&8���u�(��Ũ�N�I�
Ҏh��1�r��\f����+�`F��1�9b]��LP��Em���R�UnH�`��;�gZ:g�Y���5��*v��isl-�J�?�\����t�G�Tr����"�Ԩ\X*�8�g�%�����RpX�dxr�]{�:S��Y����[lS�r�Wa�[%�R�����Z��D���p�K�=tsL��c���e}�v8���hOWr%|�kЍ��XO�����1!B��\��T��la^'�g�J*��]1x�j+�rk�����P🫣���㾊��1,�~�!l�8|)�d�w�Aׇ��އf�����c�&�]p����-�5G�C�r���O[$�n�����?��%?�2H��s�]#n�O�/��st��,Т�)�g�������o-�ix���Fu��?{���:U[���S��ŪEH�:@��W}�Am���qj����;���ؓ��s�Ņyo�zs6+/����9��G3��� �<�Y3<���MŒA���x�c���?�7��|aZ�]�q���9�X�ܔ�!Ÿ���c��#�����3A���3���OY@�� �#�̾�́�2&P>8�#u=8���$�,��Q@���8���:͛u�:L��r�Pu\� }�peۂ��i2 �S}5�Aӱ�ikaVC�:�3��Y���Ȥ=��q*Th�T/��|Z���b��Tб~�Lň����o�u��X�q\�;�H��`pЬ�p'݂��ȿ"&�١Q�2����Z��3�3��5B��T�\�`��\�f͋ȶ' Lo�~�9�:�9�r�."���Y�M�^3��+�7嫓�*�y�����Ny�6��恗s�[����a�i�s	�c�M�C)ⳗ�Sd�ֿ�Ujx�o�7ۚ	�(^��u�/�7�|t�H`M작%娠3tiR(T����LŜ{��ٔ�_H���0j���y0�b����W�j�b�U�}{mX17�$w2uE���(��)��CQR��<���,���YX�4nԌ�P����Z�P C�ӕ��o͗d���8�Xy�CX�x��2�ɹ`gݬ�UOu�&uZc�tF0�]]d��o^�I�X�rA_�H����� �B!g�5l�ΝБ`�;��F�����v������q8�&�j�[iX�e�˙�W�ʱ�
���6tW4�6�1� mP�*�V���L �g�)-yv�X�a�g�U�.WWRQN1�����J�d�/�X�C�`��]�S�,2�|{�ϑ5B���*)���h�z=�����yE����Yeꄇ�D뺮�l�V{?�
�O�0?ԇ�����ݫ�$��c�WX�Q�	N��/^������l'�m� g|�A�b6~����!!Ve�G1R.�jA��`�*RT^�~��xA���v���߀7����;�KxtuY�4���gk���&�YG�~?yA���������1��cQ`��(���w� qT�~�"�䥮�~?�G8A Γ�r7}<^|g1�e�����|���J�/�f׺�ѯ�Z*"5M �/`���֔@��T0����߉r�{"�>cW�9�RdS���x�X�؂�H�#��ط�PS��+��#�WP��_s�;��+�u����|�TfBSV;�5��<���y��c^�Z ��DFV��!p�
���{�㋮�n��kw�ļ�v�k4"#E��$��©F�(���GV�z�:[*JU%P�ꃕ����0�B;|�F�5|�ր��>��Ѥ�e���L�Z��[TW�t:�0�`��qQ�h_Z�w+b��"g7�f,�����6q�z�2�wW8����P�3�⪞�<�R!��"�[`��Y�%݋���<����yM��~]�� �F��Bc��k�/J>�r�dI2Ў��l�����&F���t����JN ���e�+(����ڕD7!�V�V���>�P�bݺ�w&纜X�>s��J8x��'� uǒen�[��"֛�-n$-W��Q����FP@�f(,b��tZ#J_�����"xf8Q@S�����Z�Nc��s��.����K�uL��ȅ����MBړ�
J&Y3���I�ǎ����8�ly��uk�������0V��ɣ���	*֠����5��o�k�K��h�����Ce�)��?�cظ����V�@h�4$�Z-��;XzXf���\�J{����	t�D(�J3��݆���Y�>�$K��e~�p���f4���S��D��	zDK{�iwv��%���[�@+%��嵰�<SḁAV���`�_��G��9��77�H�%�o���]#�J��gf�R�A9���B5��)r�/�:Rn\���G&@9*�s�{¶ �I���
�u��IM�<��u�x
�K�l��������W�*��iԊ�K8 ;��-�/��5�o_te�HG@hhւmw�Q�i.UpZ[�`Xj�L�T���0ZR4Ur��C��"{�˼��\�5#���$["�Gy�<��K#�7�OR���Փ���u�ã�!f������LBS��={�������@Ŗ%�#�����R�0�����B�ӷ�����LL��ͬ����X��X��F/��
[�e����
	��o$�y�$ �`AT!j�C%NmK�������8����˗��
AT�|�0:
�/|�q	�*��yr�}��3�d⍻&	���b���	��|��t�c���袒j�&����(����zt�T�vUh���[c4I���z q����&�uD1��be���ҿ�N`QuW`��[�[����ѕ3N:0���yS�9X�<9}AIL�ʺ;L��׵�8�לV?�x���
C������cZ���a�4ǧ��r��|�)����$]���=G�:6��ʛU�*	4]�_d�C�����S�o�����^i/�4�&��0��^����-$�6���5
%�5`�uw�����xc $�;���L�H�f��c�����R@�(�T��8e�*��I�a-Y�Y���"���m!�'7�Y����j�%�n�Մ�b�1uui���Hg���]J0����`������T
!��6I�t��8�����L)Qݭ�笃�ȓC�ǘ���o�d*�㺔l~�3�j/ ���n~��;{XnږɎ^�X�g#)�Ppr�`�嫓�������:IMq�����=ȿ�� ��RkN��w � D�a,U(�+�����5�4�+������(f߻Q��1�������[ Ug�VSu�u ���8���2l�^�ֱ�n��g�XCӿ�~����R,"����Y�q�|Ò������um�Ħc�]�:�߬�Ȼ&�h̢�lѠu�E$����<Y0�{����ݔ�,N��`My^�3��F�p�%�j7�k�+��/ �W{��B�\ꄽ��'��fI~Y�������6 ��4M��ĺٗW����C\�Y��*��I��L��%�|/�U�RXj��� TVe"h{e��b�I���{�`@&E�]��9�|<I�j`) ��z��$<y��[s.��R���͗du���b6��)M��±2,�|PU�����)�=7}�����(3k�n[�P��k{�Ё�BEĴfPH�2[�p3ٽ��R�[j76���|Kr�;�ݯp��\�6��[��~ld��,񌳺�m�����P� h�A�xB��s����E|z�^��>�!���%^�.��#m���'N3��0��ݴ�Z�7J�|4�%"/}����&Q�W�F�BR�{�N-`4�jj_�9������N�6��1��t��%P���wQ◻���d7%T��(��.��#��r��wh���HT�̙��M�7Y�7�.EM��Ӆb���T�;ō�����T�x�%4T�-�FG�,S;2�^�yDzo��)��9�j��n{�͠��"C�L�[L�4%�>%�5��M^ŷ&}�4e0�@0"��>=��S͑P���g3RWm��I aK��:�۶��rt�|y����4�B�|�;U�*��|g�2���6��"�DAZ�>ng�5C�����p.G����E��7:�GxCikAr�'�*���
ѱ}���P��K���qp�6]�k��qu;Лol��U3�+���q�낗p��%!A�nO���!b�ڵʍ��(0��m	�{��dQ��ll��Ƥ�L��BV7���TI9�u,>�'(�2��bK��s���q�p'�E�`���'l��$�\6���<��~i�S�?u��B�q��$k!)�/7��:�h�9�ϊ��f4�8��Fd��|���8^�kNJs*��7y���/����J1��$�C�8��/��HQ�P�H鈛e�*����$�������6�P^����|nf&�|��-_m;o�� ������h�"���LYw�eح%�!�)�k�z�(�W:ҧT���Ɯ0��rԧ�F�I�|���5�L�^��6�_߈�/d"~s�wK��ȕ5���v��X�yGh�RO:�MϽ�a��dY" ��lǻ�`B�m�1������48�ߧ�u[�*��I3
�Pf�#�:����d�Κ�*���B�>ѹ�/�c���j���+Z�<��vCm�I�)|̈�&,�/�<�H��t<��)�܇�e��ϖ��NO	���4�݈_C/*���r{O� ����]Ė����7���驡{����cT�[�yD�Wk��3&i4�v	�v�λӕ"��?ޅxN�\��=�d̙�����c�&KőH�ړ�(=������t��L������pطO�-u԰��v��H��V탮���G�#��NZBc�Ʈ�cz��*3�rEq���^���!v[�Tz��uN������xT��S�5�0�U��L��d�~��@��X�K'�` �
ExoE�^>�"M�
Q��0� ���8����\�_9�y&=���l�p���9Z{ T�0��[a(\�=�
�,]Z��2n�Mb�W��C6 I���_ #��.}DI����v�-�d��^yH�Ȥ^R�����p-L��3�����ѓHf� Y�����1.L�a�a��`�@�)k���!x�Z/�x�Vp�Njϟ�G)��#��5��/��[�䋲ao%��r/|5���2�#�1N���h�(iX��LE$7��AYVB}�;����:Xl5����I�aQ�xm�Y�]�����%��ev4n��#!�j�wN ��[{,/���Q��l�/�(ǚ$�`��*tU�A勜X,�����X��o���q����HI�W������F��I!i;7Y8�wJn	����>T���ɠ��?$�<�~���&��9Ԍ�u8a�m,�g����쉳���揭l]�6��(	J\�
"z��!��2�]��H�*�d;du`᩟��0:Ix���uY*�J��l�;'լ!�����2'�%�c��`�Ŵ*𚗍�_W}ST��q~fD�l�VG�� t��9�T@�wF�������l�kk�)p*�+<���D2�g�������;9����s�D[�w"(AS�D/��`t��o�)~8Ý����+�ԕ%����D�J:�e�����A�׌��Nv�aP"�Ч��r.������@5��G+@6�i��k�O����M�����@>RN�����3������ro�,�puQ3�0���L��Ь1� �Ǚ��l�v�2{�F)$���B�l���3���Y,�g_��x���`8��:�����4�jw�%��wu�8G�1E<4��P���oLQ�7;�
ښ/(գ�����E���!�:��JjXy̼�u\��wG^C�;�� b�I�9nb��_�1�sڔ-V���w�N��U��"v��@6?�� ��]��(]�܇�I��@TSR֓��rDzT!`�LG�7���As���#e�j
ܜ��]�-T,�����hr��OI�`�oæ=����<̞�A�����P/@�Wj�\�W���)R�9��'��)m ��ja��V����Y���V���#28�1��vpa�\���8*��uн�o��`�n�T�-R&�ޟ[���\��I:�؏��^J�:rʢ{l*Q�֚�)�	Tq�#���:�P��ӛh����1s �$ʭj��g[b�z��gTVs1��f
�NǞc�g&~�QWF82��)���.�W`xy�����u�d,W��m.ϑ�����c�$S2@2���ֆ4$�Q��+I���F:�}/��b�;�������M�.���g�pBe�`� �IֿPs��[d���3���_�k��$�4�"U��z�)w�^�xk�s"�U.���R����� �'�U�B଩��8r;���ҩny+[�r��r�l@�{C�V��vo��P�O/�a?ta�
tu��w��:�a ���>Ó �E�'|�T�fY}��>z�*2�-,cC�C� ��v`���k=`C eKx�ɘ�)?#t�D̡��?O�y�Ǜs��S���D�K�͟"����sf�\�<Q�D��
�7��,Rs/:^�8-c[w��zw ��CEev��	�d)C���'��i��\|2S�c`�3��gƌ��TDd���
o��S�o��i0q�J�:�����#l��h0;,_��X#'&��׷��RiW��;/_7�7��DRD:�W�R�oD����*|"NIC�*,�O��Ӄp�_5�R0�=]3)�fG���F^� &�rW��K��%�>�[�k[]�\g^b�c/�t#��=���0K�zLS� ����������b^�4�p��S��4�?�;k���L@񊄉`N��Af cG���EY���S��7Pt2fa��U�٧?����~ۚ�KC����)-j���7�~A�%B}�ꂘ�g�~�&ζ����X��Z@m���.���3��Rqn��B�
�r�ݴ��gC�ǛBܾɓ{��y�JE�猉4%��$�<,v@���S�ܲoܩ&���]��c&0�`41��/�y���7���eJvTֲm
o] �3�9]���Q$Z��ݔUwD
ʟ�W虻�ȇ Ov�l�n^���=���m���vQ�@�@�kc��i5�Ah>��z�^1y(�+N�{�^݊1�\�U4t" �]h_���OF�>ߕ�J�;:��i�H�2���{�=W�W����^��31�E�Z ��y
{R����h�^u�_O�\�����g�Gҏh���>�T�]�M��EUҲf�S��v��uN v#6;���� O:�^�D�ϋ��\��[?XM떤�.�_�N�֤�����1�ח�5t`