��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK�-߿�@�Am����#���i��q�>��|#��Tx����L��N�I�������f\�g^l�γ���=�Zg���Qm:�cݴ�Ng��`o��e�Cq��6#Q*@�V������T9)��ۓ�!������r�RS�� �SO}g�S$A����a��+J�e;=�e�X
�dm�-J5�3�=�'�J��q�]�p�\Xz#��:e�nV`��c:�ϳ��?�,�+�50����vKy&�H�̃�X�bUw�3�H����ı���#�&B�5��r� ��!��6ʪ��
x�SE��pٜ 2����H�Ti��3׾���"����j�|����%��2�% =�+�q�3!$�|U�V���-+G��U�xєXBk��t�R�6����oƢ�n�ueE-�J.b3�1cM����T�&B���4��m��wu�I�OL-�ݗ�M�*,�c�F��}T�i_m>�v�yQ]���pE�AE��ڦ�����~߇���t�pz���qI����X�ȖEA?�b�Mg3h�d8xga���������J���n��~ۤ���{_��i� >��yH��@U�n��i���]X��a���N�tFE��n�ʤ����!nA��&�����!|wQ,����7��/�؆b�j��Qnf�\�F�pk�N�q��6t���5�Ӏ�M�:o��ݨ����'�ר�{͋m�2n��s���sL(�'EP�]	����0B�҆��{����K ?�k�<�,�G�w�+o(�?�q�6��@�=#����h{xGJ�s�Z-"�+�孞Y�mFk�����������������	���@y���];p���8��i�T�Ӄ��	3�������.d �S$��"��l˄	sbl�\�q�4�}��>Z�%+�9�N!�D��kW���p��р����������!PS����T�kl�R�ց���*p{�!�Dd3"�y�V�J�#J%�l۵�-!��,�,�����O���F%B�6�%K��8B�H ���Z�<
��K�%�u:�Y�`>���۟j-b�cm�а��{�n���$$[: Y��H�oJ�>K�K�����IIX��Ҽ�'��<��}c��]���6�MU.�A���T<I��&�t^��>��0��Er�|��­�Q�M��~��]]�����62��,�Q� �0��WZ�u��u6QkP�sJ�*N