��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,�������_^�6�3�@�RU:(�3�ݵ���_�檀:��;[�M�+����z/~�T�M�@�9��%Mި��fRP���G�G�IS�p5���Pp���.��>��ǕC���+X7��_�3��w�'3St���<P���
S]�������t�/��x�+ޗ�ȡ��S2��b�|<\>p~��e�kb�̸�B���
n�9U���=#oi���s�r+�Q��^]J�PU�b����!�P�����K<�E�r�i2@�B���p_���}�DR��}mSW�g����a�;BEn}���r��B�H~�~��<�|�yQ�*U3�j@�������d���̸"�b��t#��J���e�t_�u��y[[�.�ϺT�^>�u���#����x0ԍ���{��V�ꨤ�|gC�;��S��l62���Ccezzcuu
ɀY�ǤU�RB�B"��7���3 V7�!bO!�/�(�Jq�t,;��n��NV-l��7��]�΁&����@?���L�.�$��)�!�$z5��hҲB���bm80�W ���V.Y/< ��.Qu�W�F KU��"������qP0��������-A�KfE�ǹs��{��a޾��{\����W�C� 7�tsW;�\���M����A%�В���pO(:��^d�_Aj�o������|�|��ÌYS�?<5�c.�>��6�31fS�5��xk-Pb��lO�0Q�X廁�!�
���(�_��P+Up�χ�l�y�\��UU�2X#�e�DEww<�t��ݐ
��U�W_%E��խa3'�o��N<mK�?q���ؾ��O�F�%�> UF�����,\�CQH���n'���B�k뀳�����>�E���>*� ��2D����Ŭ�!ۤH�p�ٰ�z(�%{(���8 ��4������^�4Q<���y��S�p��l"	�)/d��_�	�/+:�|�H�3�z7��_�k�ӆP�p�#Y���_��C>?G
W�A�R��4�P���E���ma���.q�wJ����6l$[��!�Φit�f�����ȷj���Q����,��T��T]�=ݞ�}ıgXviu�Tj��yuv`�H�w������77<�ȟ��~�`�)F]��@Wx'y}���l"��dG�b�{��_�O����@?�<��P������J]�ε��5As�RL!����F�t�!I�x��V���j�B���Wl�n���Bn���^���&/�*����:���z�5tZ7J/UK��9*�Ֆ�jag�;�r�֓�8*����Ea?���}�˯j&�u6���kϜ��ʘ�$�0m��m��0Gi9�a�j�6B
}v��YV��__8ѝ����!�uŧMj1��q��#��{��\;}����^C�3��:�c���4MS����d	{�b�����!֝7��o.�1ۉ�� u��x>��K�^YO���ϥ�/�`G��3����9�:�\�D	
�٫Ͽ�L��]�ܓ<Ll���l��������x���+� �W|(_�ۛ E���R�����(���#\��/�ă9�>д`@9�Ð���w�}���"���)�,���7��4��?��x���VAf5���b�+��b���|gD�aM�E:|�#?�=�r����|���"��P�����$�r(����{j�Mw�av�F�s�)�|�V�7*gǞn9A��r4�=��?����3�43CQc�nÿ� �������d�N�]}���$?ʽi��Ǝ��x��M��<.���]�y�ŗ<'�`\��L���`��O��썑��0��������A�vة��0��'nu�L^^����Y����[��h��)���<)􆾘9�`8h�
�����m��݆M��5Mc-�N�^�Z���ӖqӪMt`���^5#1�2����7,Ď.�cȹ��z�D�.([7c�����]Gx-����~���I`�����l�Pm~W�f�� Z�_�X�y�#<� ֘|�~`mw��<����:8��E�_gez�9�q7�c�ތ� �W�p�� ��4��r���+�=��yG���Φ�����OC���;���>����~��/w�v�����t]Qky�޿�����)R���D®a�i~@�C�9�Ď���G������o[���_��_~���xRg�B�u���Ju#�+<R����l��g�w���4� �z��C�ڒ�/�I0���I�3��M5Hnm���O��e<cMi0
%g�Ii��͐�j{ƯM
(3�����Ӗ$�m�lP	V}��Y:I.���Wg���d]e���Gx��%lT���D�z�3g�U����H��*}�r�y2����{iu,� zVB�u�� @s�뺃��l��-(2�k�_���u��Śӈ�f���d��b2�"v:����3vo�5����.B�^@
�EY��p�.H�f����U��(�	���r�����(�*�J\�!�"��b'T<:�>�.����������!�=��z�8�;cֶMP�4��[����]|%��c:zj�����'��w��&!���;��fg�L
�\ZS�}�I���F�����b�C�Ijc�<���������[��C!^֒!�1�B=_Pp#܃��a|q,�*���u���ѧ�Qu+��O��1L��!3C	�OYU��uj.	y�!�Vm�P��w�"�V�9R{IL��l�����{�Y�*ȥt��a���*�_�/�$�G�Z֚�q�
�G�̊�T����+�S.���t��gY�^S~��EI<��"�Y����H�*�3g<`xo	7Y�={2��N+�M�"��s�/��7�(�\�g��7�pŃ.�h���VA:fU�Cs�KT)���mS�)m��[����%�Z������&�(�S䑖HEG��%g��9�X��9A�`�B�����/���o�P&������$��â�"�pf�'f��2���������.��*�;�y/e�%��/ٝTh�I�p��u8��F�q*>4`$A�����nB�����������[A��ٺKЛa��4r������Y�� ��Ɣ��o���ʌ�-{��\��S��j���#�4��5�����\=i0��6�����V���N���X�>
��7����m�NЃ2qi���G�/���wc_S���@�a���Y�r�d���Wr�T8���H��:�A���b��S�'��S�-����+󿰥��4�(��/X���}�;��fl��y��ޏm(��p1<p��f��1����P�}HX��%Q���*Q!�\�S er��k���p|����e�$��Z��#XW�U
���<A:(��mrw��d>Y�_��(�����6�`[�����ty#�:؟Y���5���%c*��܁�҇�!�-a�	�E8�+�-9��[D�A%�\�2`��-ɮ�^�c�G����҂�3���t�zN�7�EP��דٺ��t�	��s�₾ qPA����M�R�J��R����k��u���4��d�Vk�N� �������,��!�ׄ�Gh�'��%�͠���x�P-�cU�ƴjg��ۜq�ƣ����h,��J=�Ǡ���%Ūg�6�jS�6@�ϭ-����������[�RU=g8���1�t�H`k�*/�\1�n�`�q�S�%0nhپc�.O�\�0 �w���b֎��պ=E<~)�n;��w�j���:x�_��!��Ƀ:G���C�,�UQfI�r0�s������+	��i�gK[�wRGW0�q��7_�n�a�p꘼�VjHƠ�x���&�t '�1���:����z�41��!�ca S�X������@[t["Ňe�)�_'�2�k
˜��<�+��a��KCwO��N���ٵ]qٱ�9�������G4/f�U �*JQ_ʺ��^t�m6)�%��j�}��ZV���� ��g�&r��؆�����[1��G�}����G����B8_������=-�~��v�d�O�7C���%��5�G{4^��0���H�ᚇk�a	ꦺ�zT��!�ˮ`�C1 Lj&�l�h``8h�Jݡ����j��T���W���|����;,��>��l?WlJ�)�`��Wa�X��O�y���{#c�x~�~RdT[��5�ϒ�"�0E��3gU��ew��L~zˈ/bӹ��T/��.+俢up#��u�&�IXk��x�wM�wpD��4A罯�<{��'Ji��ī�����l�j�cxh@�%��kX�s�ݡA��ye!�;A+`��X��T�r4��.u.�����`@�4�)/���jm&RaM_ؿo��W!�j�
�d��.���
KAdC���U��q��Sjn"���	×���RZ�C�)~�;��λ�G�1p��>�]�N9ǤbXυ�.G#/�-7�5"j-�f/�e��z�(�#"���?�(�+�H;h����P�"����#�O��KC�� �M�v.�K�QM�b�FÄ<��*�I9��Gr�bW�v	���rH�C&;�����g?���mT�����l�p�f$�A����%]�Ć 3Ê�^��ϓSEF�i�&�}=8��K�Y\��su!	m�ݽWm<�e�y�]���!g�Zs"����ٽ+;b�ͱ������ ��|A�֫�7���V7�����d�[u�ʔ�����~��^���dCsb~ə�L�����Te@_:��P�nY���9�i5���-J[Y��mǙS2B����	�,y�Í��5D|OZ����R��L]���蛔�=$�"�z\�[L߾���=w�/�v�E�A9{W�kw,�U��	)�{�V'�|�|�յd�yN��[�<q}Pa������;�Af晝af;���9@�˕&��
 �@S�|����{2h�B�.��C�@a�cQo�"ق^�œ,=+��j�L��}�EQIj`����A!�!
���4ǯ�heFS�ז��^YyEz^�C�0~똡��� �cNT�5jq}T�w>���!��A��#��SÞ45��}yE����_��Df6��d�B����+�.�p�*���a�] ����n�_2��X��>�t��*���y(۰���aª��f�I+`ZL��+���c�2� �l7�\��zQ@r��A~��}�ٴC��z����YX��LkC���o�\�0`g=���7����8������K�\Ȃ�'�E�C��@��w�Qt���n@����\�����?���U�\W��`Ӳ�6*J^�@cmb�)��c_.�K
 ��=��;���VM�]C� Q��s	�MB{b��Q��%�k.������ψ>#���Hf'py^]�`��F$�ώ6s_����இ�Q%mZ�KG?��
ld7�˻y)���3Չ���XԐ� �H4����_2> ��4j�
�`�;�b6XXs�RQ��>+*�k3�"U����p�Fjj9v/�J������������z����X�� �ٟ��\�z�}$:�.$��p9H�g0�PMw���PU��E��/�r�;�����lN�-@��P��v,�U��Oj�`�a�k���[=�r�xk�]v`���qrc� g�cC1��^ B���]�tM�"J3}��J����1���)(��f�ۏ�-��vzn��W������cߩ�����Ph��=�ز�0�a�Qv��}��(�hS�v��7R� ����2���R3��'��
��K8�G���T2��߂�d���&���l�U�3��?h�f�9��n$�)�_u��Q��.H�Ne	��`�~�V^Nd�������I�� �s�4���.Y]�m������Y������4��u��:��Śi��<�����3�\��(8�UA��y��?�j9�(�S�d5��(a'64��o�k_ �	g��T�_�&�@s�I���p�O7��c��Ǜ%��e��LKT����O�q��
��(\�L��%�@TsKIGP)��{7��$w���@$"7��&	��B>�B�R̹a�%r<!��3�2�HűUϝ��2��~YPX���F1�7�֚}�I�O.�"m�3�0ǆ�V7�ՠs�"i
��E7yH�
$g	Ohs��f_S1q�U�ov��L@���ikq�.�����KF���0�Z6��Q��x�Ğ�$�3��79�-�>�'v3yF�Q=s�L^����i�}�+�X럓 o��E���A���d��Ͼu�\z�E��T��<&�����߶~}��X��A��2�A2:G�x���QOx��ntJZR�&�k�A���X�T��kt|�� ��ݫp��'�u]&V��!��<ͷ�?���[cnr!�����t�U��C��$ס��k$Յ��#�����Ui��I�����#��F�9ڢ{�=m�L�	�p�-�Ɔ��%l��XH�1�;�o����f�5W�9�(�޾��ܻ,��3YU&�Sj�x�p�)�AbY*���� FJ#s� �'6�Wom'�gc�2ŗ��"ZcXIbj�"̇3��j�Ջ�Tk�q��jal'mvlx �~����o���&�t���V�䢷g�l3m�z|M�����>�_��E�X��5���'�h�S7׶�P��1�{�B7��A
�z���*�kPnK'I6J���<���ܢ�Ź��=V�>����~<J�^�u���hHO�����vE(T0�ī�S�.��B(�A	:�v��
��X��y&�����U��N�D�j��ck+P;�E[���ϧ�TN���u�-��$��\�����B�\Hݔ��H�1�5!�R�:}���'-b)��\CWm@�ɶE�}&��yx	G� �V�%X$Ql ^�pb��2+��]i
������:Ѥ*�����8��yv�)�gޟ*�d�X��L���B]ڭK�
��~���p�����f������dܼ�\�����r��KdH��)��3,�נ��(����i�:v�/FD\��)����ݗN�C\��sy��@�!�q���>m�q�&
T|O�HW���d�y�ډr��gpziN=�?�20�t!��q�S�1 �fj&���ݾ�g�I�;�ao�O�n�4�Z��8��d���I��~����3��E��С����Vm~2AP�r�1��燕Xc_ڭ]���ι�DP\�W�C�ǝ�׽h��Ф�l�490R���hy�/��j}�&�
rޠ���`�K��Cd�Y�V�U�\����S�����Z�ۈ���`x�]���N�t�)�+��@/�㓎�i��H�B�{���H� �<vֽ�eU�6�<�7Q kiidg�ǁ�����+N�L{�J���ׯ�iP�Լ&cf���?�e�ţ�~=[�O�q�.S�\hE�#-{�h��p���|=m��Ο)}��`���:�КWV�:CT�4%�X�B��r���U���V�h �xݻ,�,мPb$��y���t�Q H�1xd����U��*S3ӌʲ]qc�_$��ѽ��h$��#�qC���aN�5D��yh��n�pc�k)��I;g7@~/j�������}
���2e�/�fu� pjɡ���&Ȇ����ӕm5Juq�Az窌�d�K=5}O��J���-�l�Aȋ�i/�)�a�96��s��u7&΀���4�Bק0>�k�CxE��*��3��]?)����{�Bg,�sr�'���]9��N�(�:�|o_JsW��C\��p�]��OS��Q/��1�@r;Nf�����򡲺�`tF�����V������VA۲�
�-�d+��7�1"��P��^���3�ۄD�)���{B�v����p5�d��o�f��;3�jQl��v��y�^���� �E+3J��Y*��n��|��7:�d"�̈�l�i}�/���e]��q��Z�����l�}��ߵ�L51H�~�g�W`�N��K�� d���I�95�!�H�ƧP懑�1!�� � 4�Id&�h!�!��[�Ӕ��s�gx�^IG�����EuT�8����P�Z�v�#��%I��cn�hDD�8��ᢟO�8���5L�F���*�N`��W�h�(���6� TFta��vd{������U�.�;��;܆s2����S8ib_�Х��T�E��Xk��]޺_Η͊�8�v��BH�L��E�V���ZC�K3�-;��n���g&�
o������{������*�KnXӄs"�^!�&�K6qp����\���A���΃og���cƟK�k"zB��!��1��Z�.��> [�BWϹ�����J/y0k���5{o-��8�^��3��s�e��Fy'�E�����0ґ��h��T�P)�}VZP�s�[���Jo�]���T��(�Y˗�	Lf1ݽM�-�K�e"Z��lu�W}�B��I	9�7��_ĬK�N���:sH�W��Y,��UN��'OAaxL$�q a�F���Ʈ8���^�l�]Y6�yer��{�U�z���͸9!ϡ����eQ@㳉�$^A������4	� ݦ���ә�ZT΋��7�gK9�'��P�� (�7;Pcx�x�}�Q�op�� �@� ���_��uc�y,+S�O�P����k�g���*�:�4�X�T���~f�n@On��
��O��]��o)���|d�p+Y�p@ϧ���a��Q09�A#�a�V�R�&�@��r�+�ia��3�'��XRf�������Ou��������SX9���AV+�ѕ�4�+}��O�3n��	u�<��|�%���%��k��h6����"o���ʱw�t�צDy��[�jAX��
���ښ���MIhK�R{E��p0���C(��aO���v��i�UbU�E?4W��JȮ{0�^�ǚ��L?i
�CO�%��R�\���>���eﳀ�3ߣVL�{-X�U��#� �
�_���a1�Dͽ���u<|ߦGܽq��坫� Kpr6���X:���／'W�oZx�������(�<�a�h� ��`�,�B�\�09�	E��}a�"�/��j�2"طS�^�ȕZ����w����I�޴�J!8 �7Mo�2�Sy*1�e|�\��J���z�]��#���n�3�'-	fY�(}����9Йp�t��u>�9Ϝk�_��o5�r����/Ԯ�u���]�x+1u��F�~-�M8Xg(�����V��EA�Ț�2�?�/uKS��B> ��)]g9���e؂r�i�P��k�q��4����Z���z��N/���$'�&���T������ؿ��p�Yk+4�e�D
Õ�m�ɟ�K��y�#JY��\���e��{�vK�o�(����Xij[���B{`8%��Z��RY�a� \_FA���J�_D�߲�'.{�������<��`��=���Aʬ'�LN�P|h��p��NL��pMi�R���|����	K܆^9Ejt�B+�Uп"�܅b{�F�?,J��9���#�蕝QZn*f���h���s��sV�]�Kg����GZ�T��v��-^������	@�i�������(�1�����;S�^����<��V�;ce���ɋ
��i�>�����flp�ۚ"��B��|�����L��<�/�����G�q��cF�u���;&�O8��e�)
ćr��yF��f�����i�[	�\6��)־�5�̆��7̳��v4�Y���(��wjn��D��ة"'ݿ�$��w-"G���@����Yj&�y�C>$��`.!�7d1��F�b���{�ZX�x��y{ݥ�#��	>?�E]+gKQ��w��������EV5^�WtjN�0&gd��3��>s��t�Yy��)�aѝ+�,f81pȲ� �,w�X��*]�߬޿�}t��.�9��ũ��2dmd
�&�l��4�}W�%�'�>$�lgԫ�Y
0B��&�pϏy��N�h�� Ǚ�0$A�x}y������$��r�O��� �
�BC�os橕�����W!�{i�|W
�:�}^�?]�v;_{��\�k�C�K��I��W۪ڿ����+�H�V;�?C#V��	�7��Q�6J��M���s��I��ƫ��I^y�m+L�s�\#�6�s��Ē���&���{I�M?X�8x�Kꃦ7y<�X@�����Gl�Jd�Y/6���U�Ql>H؞Is�^�:��z��0�o�ϲ�:-W?*���������vlx����B��Ho7�u3��h?X �1VPf|\�h�G��+�R�},��_y�%�]����D�䥒q��G8�"+��:=�ɪPԄq�@u�Si}�
F-;��c���I�r~��[��y.�0d\�z���3u>������4U����9_������3*z�~��K,ɏ`�%"��e?x�ءD���l��o��s��<t_Q��$+Y�N���Օ����K��_�n!���Y�;����cw���]�f�!��z��*I�L$*�I����4l-�B�5��3b���I{g��մ���=DTz�[��������<|]EfS�?C�,L���=���|����5�E��{�������A%I*�^�G'
N�%<�Z!8q�1'&����W����$� r��0n��vt�Om��RK��u;�Q oZ�h3�W��r&Ƚ�g��R2$"�vK�B�}��|�<&ѯ'FTu�Ti��&H4<yd4ͻ��Rg�b
��:��������� �W;Q��+�C'��v1�}�+C���������!�3hL���o����D������()4���z����N��,į�G������"�^�]�d�P�+RHj�J��STT|�ɘ��I����e��蹸f�`O!��^��hi1J�b���8�:3�ǝ�n���I+�h[�|¬��
y����ƉeK-p$|'<@�\����,c�dQ�SҎ��T�M��d]Ꟃ�l��'W0�+$1R��~��١u�F@J���獶��/�C����^�s��1��"(�N��Y�ܯsN7���p��𱍚��P��k}�N7k;�����*�3�J=,�L,Ro���ex��%? ��ֆ��QW.?��������$�������d��R@}�9�-�!3�� ��ؚ��(�gk��\ �!�x$����]�M��5��ӡgA"�~��\;e|�Q�Rm��͊n*?5� �1��.��Ln��N�2#8���O뵲װf�I�-C����Th�u2��X�Ú����7�u�c���O���O�|g���(�{�-�|Ws�