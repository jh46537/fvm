// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Am24yLBWdVBKwliLbEboqtICIGuXkfbO1K3v6k3DQikQC+CEV6bF7bWR0CAXMjb9
Nd7rFYnTBYO/hpcAfmeNoj50pfsW4fjkTBXbTW+4hk6/WuoxPpx/fD0yQ/EP7wCA
zSAr/QvWLgaG355e16jzNEYBPYH4Hdr9278GpASgsS8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29232)
d0FF29Mg8iCujXpfGn2+0UzcIBWFkGAikBX+opb+kMIiAMr2ropNpK8l0LlYVwAg
WWEzteY36kyrZv5l47aiEBb700lCdu1KwRGTbuv/xxpxlXbsnQsTudoRpCMV8xdI
bl1Xrwu97T1nh9mnJm6soVuXhJyMJ7araqu1zxzp68WT0oqvICctcaMm7CPi0EEy
jIT75PwX5d5bm54QDdbpgjv+vwSNqySVhjEcMFTQUjgcx6Z5Iv+2gNpFoUsu3dvV
tdNuHJ+pXToUf6ZEWB6teR35D7uAnCr+MqQUQCqyAi6Mvurl570sb1A18XMOWUs/
aQwjS9Z60BHtE/pVUvR3/at7BvKN1EUJyzP9EeS0JY1NVXrzVT2cmqWtK85PmD0k
IEywBlDj8/vTqBUt6gR7F+Wswbldkv4zho0dUiGt2dgHKqWjdTRJDQzp8JnLgPPC
rpdcbGrN3dCvqG55iOTHno5ORzBi1i9o9i3yU90GrPZ5BPHaTRcBuOa+Xj0rLJJS
f2If+xZyGT4avCIoiyqor1G+IWn4/Yk6LqzpEpA3aJ06fJDfCBSkq/KGgRXUsXn0
vSFRus8sF5AYkDxGfNro2Bwutgt7tkKdidR1K5XME/Sg7ciRMo30SQvRYnp0iD5l
Nw14dUKG5n2V4RTs1/sMQRor30JGaSPy3w2aqUScwJQiw6V5q00V1lhycNUgrGU0
WX1gBABLcyYGj9w9ZgLnhjksMWtOa8DiXklgXyZpVnHV2uepU2PTMxXBCOBn1XX5
08/Mu2CRB8ul6QpliVyKZhB8uoN9Nzh6FkOU/dhmP9861I/WkvuLxiZma8Jb4v82
gLZ0T99Q/roxMYhqLNIaIgoYGuLwyIDQi+r/6B+ho1+uT5WnOebUXpKtu8Hv17qT
o16lVDP5VrFA5KoHiM4XMzPBlTL1RJp0JVCZXLZyv3jfVRtV0xB139enUr0amhik
BTbZn0B5x3Yyz6n73q1CsHCe6rLRioGKBN4G3rfsth2VA5Re06VmRoShCFg2jojH
zNRVRVS6crUdkNCUjdLWuKb8v2HUFm9WCuXumX39fpV4kOLw5izBQWEPoKVBP3Lo
6x58O9cdjkbOW3/LdRdEGquzdrnVI/MTSCK4t2Yc9Wt1cAyf8Gb4px8wFpzGyuyV
9LsVfvMvMXHJ385nR18Rx+yIWyLWBcfbWzksKQd6LIYidu5pQ6mMaWeQAhYb1t6Y
fodW669jA1zWx8HUT0n38zIoipPai1MGY7p2mnvT/rFHFOo8LWNTc/2LBlVAdF2W
+hizsjyw3n5Bgj0SnaU/V/7vdvYdMOd4VeVSbK0TX80/ZE9pa3mh8wytJ0a5VcKJ
c4AhDzWU/LDV18164GpQJW22cSJGOi9L35uTO4hDQNiNobdix3ZG6y8VeHrz1uHH
/u8km4G1hhdEgs2UiLawAr5/bLCR6LquXkDTI2XE5D67DB43WA7FQXiFDVEGtwvm
OJJAWCsjvOca6jzoln7W8WfWjXMJyZeAUkkc79m+zz6UYQ/J+jJRkKVFi7uYP8lN
fRB0uGsTSQl0RXKtaARE8P+kjf5aaquuauPMVpIvgtzRrZcWQMGRGpnUrCdc1vb5
/+V8ZefynEPUJFCcguSo8wCKxOW8inqaVzqSUGJojXBJ/C5YUSulzLQWvhfzZAKn
+XBmjt8xdHQkxC4ioGlDyrUUej2YgJx+z1OYYW10DmVGpTSXvtCp9H02L2hmCLvS
KgNbDATFJBxsql3Q43mr2ls6fcOiiYNjgUvM79h2/uqOkgrWQmVUxnv5Y18tYMYo
MNvWNz9Ib0GSkH1a6uQx25MDmCQxCaB/oa+Ct5+iJze1+0hF4XGO2OkzubtZcsBQ
BKbOe4lq8O37OX2KIb3B9T6+AkuUY94YoBbrzzBSxV0mkj8eoARaY9So5wpqLxB8
VPu9nrD4t9hZY8N7J9S92clGRUh0QatUuqXWOCJx/XYQJxDRESZwAnubfx1H79zt
l8KJFoaf/NiPDssWNcwxMk9p1GoMH/jDHLaA6Vp0yoR1yMj0ocuq/MiVxG0ocDcT
rrenTgO4tk7S4hVDllxgU2n6BihMKY6Cide03US8j8bkJEFDMSwz/83x2TaHui7y
zvMAyR/jzlsx1zYW62CA85kA8gtDLdVOvXjiZscoIq3ZI+D6oOWvqouCvKWtMu06
yWpTUp4aFNsmgs1LHgBdlhxorZpJW0D8q2EbFkYmuS735c1Y0BuAr7q5QW2UxnxU
UQtS+4RUTAyK4GozZ6nY+VTLxjy9Soac8K0LlZM55sCZ6007YxB+peYk4Ra1Hw5D
cb5NVxYFXeagwx/ZEtQ5824nVkl7AUUXSP+XP4drIvGbaBs5uw4FL6bjbjjuoBtp
VvHwCqeE9l6uilXjoK/p/5h4IhLReGIFFlaTMnTrGBlwor5OqDilhkpu9609Pbdd
Y5K6irsUbgdp9hPpcksMjLcLCEAxXGu6AL22RkswzU4dnQrN7iQhGqSBAYMbxiOq
lOGV32lJHysC45Nr0tzkaPlI5NdKeELbMlKC55D97MMGrABqm7bLgDVvNavv3sml
QZXA7dRGxDnRgdAfVvo8Xpf3MbftHRU9hWHWPANB9xcl9/GUnbghQhM2snUKiGL+
6BFdHt4v9SBdOQgqGtifTLX2pfPXw/5XxPIYOoOl/TkiFunpMuwLOc9oJ102JY0j
kURpE8RttWlC5Q+H1K64ZqmvKXZP0oZhtbebIh8jmg1lSWGf2nLupgyx8AyGp8zr
xgL+yEg1gjyKJF53Zzqqrhhqvv7MV135gDC83Yn9vqAODRlz4hSq8BkPXWwAebYK
v7xJ//bYgxqT4O/O6R9KiVdRJ/b9jgQYCl8j1/lFhlqhFYWv2Sn2ljNBKnXPa6g7
Zy2FzTofUcaMosvnl/NoAce8XhAQIK3xWxSiRDKqtawQOEpmqd3a2MYs7tKckW8D
kHvaoIzfFt+FLs42sk8fcocbyuSoWAZM+nVJUpBtUQU0LFRDAvmA1UCMoApAK6lI
/jwCZuv0mRQ/qQ/ohI1sbH3RTQzB8Fh5qiW3Mc2Wu65RwQIlSbinzKjhcIQoouz5
DMzzfmrdk2kR85FsUV7//uY/yY9tyNRlqwpwlytJqwRY9QF5vgqy4H6QYLElnkn0
miEo5QVNDVYgPvFO9x/LRVhOYRXyPOYE9TByMuZo3s5N4+KfJSeC6O+2GiR4XdfP
jWZiaiVustFdzYsM0wXpL5Fjd2Nk/0g6qnoZHGF5xun7B22zop+rh/6DRP2oNc2P
3M/8eMfV0+wYRmgWN/uRBwWdvHqciYD/RD9gLH9wfZQZ53ofJdgcaS8gh9DzddO5
i8RVBJ1zkcJhfZkeOyf4pZ/T5INrSCYibM/YACFpuOf5blWCtTl0QROjgBWFuuF5
yh5meF0SLkmaZfhY/xiiM0xtCev9nFECKnUJ0TjbVRq1dNt3UTZQteutiFeS8ljE
f+fhkhDPRii2eAz8GcnW6MuNfPE2PhM6T0kbVZy73cWdQ7L7oK41kgCgBTJCQ/Qa
wBBil7y8N8kJv2GWy3od4qsYQRzj+bRXbIQVGzb0NzlWyZBRwj+DtircjILh9TQ2
wgVF3GBEh/vfCqeZrVn58TTvGJ0aDNC2RE6EKW50fGPUDQIKVX/N1az/dzk/oYO1
lfyFBCU+5/H4E68fhQ7lFgvdhAgxZKYwRTw1T2Ze8RvHZ30uzSiNZ3HSnrvS5+iO
NpJi7PYZ4eB3AeodrNN64nlPMgpgQ230u8+vrA0acvh6LSg4As/1LuZM8Ko9MN9P
tFcieG6320gURo59j+u6mDtDsZlnGs2cE2hPChNkf9V2dM+0D5GggkSPuBD46vKD
tqgdTC+sQTUJWdoIT8Do7gRA9ickVynpK6wwjRjT6t2QHch3TSyHmE5Gk+3IGsI5
dUtHpO+F8lev1EKBLgNrIrDK0LWe0u/1EnnV2gByR8L+iHi3milf8AnDoI3Wcmq9
IKZZhI5bIPTLniGZvKgd0Ta+zAnUSz4xFDDaNqXuDzb+RfIS77vNktz0nW6CzX5M
Wl5yy6QSwfPRGVx4r2WQ6gGM8uxlwRjL3MRKcNw1y17H5TsZLRkVwddIFEwNC+aq
zAaYq762BhZGW0G5rqqk+wn3Oo1SZVG60mFnYGpmX4GjQsl/y8oE6pQTUBJQ4Fts
U5IyS/uU+/Kxwpi4D6xBgTTUStxg1zZ7z/Z+E4SLXFn2fLJS9FnC4OQ0mSI0Oz34
8KuCPFy+gxsfwaSieM9oRCI+uw6HZs0wrar1JBxPCWSxuXfEJ0oUIrx+nYH/d0Ct
I3MPfFpjdakFDDoTLGxC5v3HjoJcsrKsg6ZqyVQsrTVnQZS39BJHsMmT24KU/YFN
PaW4KikxxVR0ybYtmz2bNeLm/Itc76YBkuqCNzSRlFif7hfXQYeaEVIMJ6ey4tF2
saH5NKIM2mvpqfiXUfoaeQUFUAnPtI2wR5UX90ag3UVCYnw58CbvSIOBohEbFbaA
6W4Pvy1wE7vv1wosADwZEscIr5mD9yVkGkLJSsGDgHXGVVaw+n60v/O0RvzR+61E
UG6RhSxjAqahwA5DTtBu3ZvIRqmAn2w8Z4d+5RghFbacXNp4C3nlkgRq99l3wtrN
BCfHUuUw0AjnNkBbSZ1mAHIBcQzol63gF2hG6/dlU1zxU8kC4U6kvmLtNhVgnOG2
XlKd/K84qznEkmLLTjwXuBGpv+9BUZ7ReA6tVp+r4GADFr8liMx2j4sA9GrQmel0
6SOKJD8C5vrj+E+vHz8/ieFPDHK4JkMHkibmkIpeXbc5OUFeOEBNGtxsDa2jbSsT
TRJKo0XIY9GWqvng2sydbfrF4zllAwa2qYffCkKQiO50hZADgbmyKdJCoD06va+I
ASKVscFOn0lBjFjr5Z/foXb2n/NaGbDfY/5x3rsUhVzXTAbKd0g9qiZYMudKj73N
hBKcfbsCXjDGlG1MIuxOCJib9aCUvXDrJ4ZyrKGguHUSmo4BK0EKm5kfGbNeUS0C
/dcnsKum++dLoI2UNqjzx9WqaIICqZLvptm0NM8jNYUMAJedI6l/72vTIQkfjnGt
tCLx65ZlBHRbNkEu+2kBmI3mWXCz9AlkYtPmFueV6oz2NaEMuJnK9qD1b8gTQOTu
Rrzd9unkFBP3PKJ76GBlR7Xda7tzef2AjWd+QQO+84KtJxrsVCmyCiHROj41tJhq
doDW0nVT2tZoNSTxK1BJX1LCblqddw/xlcOAn5IUzRrOk7JciJ5k8Ln4mF+89gEn
HoV9beme3Y1vAOkXA4ReZKei+enK5y7LYMwV5rnGJtikDXxwMxDVyLUpWD6fK6Uh
hgUvgYLcNHOhkg/noH2jv+fXF14VTt7uI7YXS/Jp/kOoCoLRNIrn+ukX0zYTIvQk
YVcucFzYBEpbJSuvGG3bKamt0eTgUKJmhCX2Na0VH/P+6VHJCVYk+DdTS90qkAky
9EleF1rk8pHdVPhUV45m9F6kXHgN8GzbWGoCVhRbdN4q+VeE1EOzuPNEs+Z2bISn
WHIq8jFQm1W2gz0gU1tJ09JRa9c2+Ja+DIEnOrjpHidqyXsh2qcB0UlrJq49q/2s
5tXkHrS/vGcdUqP3ES/vUHlLqqcJF1YWqj7Vq1g62gOroEY2rVdbLyNOSdiyFDv6
uEkn0iO0svNxMki/9xRuVChUYPkDMRj5d8XWS+1Vr010Nz0y4hp1TrJ3yOvTBwy8
tEBoNejVZ1Zo0oVxXrH6AEECaCi2A38A2izuwIZ1hf4aFIjVWLojYgNSJa+z3RtP
qL/qnGuEufFo+mWS4It8sy5Fh1C+Xo5sWunpXS5ouo5mm7B1OBH3rpIBGdOSe3QR
sDy2BIvax28HOneqyvlAqv2adnhy1BFGl4NV5zLdcyzxgxCkNTIgWmcxCR0LX1pR
SfVPIFTrk/epFBBSzINtNCY43h4TqaKM8E5+N/b3XCYnCmJJi7alRCq2iqQHEfP4
r216q1xfRDAMwzUW7IdVs7dTpHZJPyFXNwcIpYnFIj/WAhvFPmeOzrIfmYm+s/qK
ZNWQ0jmADlYGPnQV9VeYTZBquF/uWp3zNpwsyGdbXNfuPl1iQrS4gRD5oV7+fDAP
tCA/TMkQphWqJACLuVMdgXBgnoHYeVYS6e2Xq3bs/XcDnYF6VfK0mk8QJZ1XXjYM
tlj+07L+UmJ30HQFq34pbIj4bc9ya298zwhSDYQdBCGf8qvc1TdDapAFeDe05j76
pfUXHCqEgb+YLtjm8zPhkZGXu4kWJkqIpRWuarP0E1xkdbEFpqr2qscOUqPrfEtA
FPUQrp9rTIarPC0Knthrw7O3Zj3Yf2zw0Sy7ZuRAA3uTZjuHDoKBkXHESDwE+QLX
bohU+QkW47KeI5lBktt87Q5S3+RpYxr8CrDzSmcFF7Oydon3fI4u6m6/ZiuB2N16
UbIyaOrn9tPBW415gDHLE8TweJakW6iSGsM62AD+JjCVFlEhuFv29r1CHH/CMHPY
Ms7HOz0LZZNyUDSI1QDVSyHhBXjD5NGrAHWv5r6CB9iP2XYm7UFh9qC/jLISH37U
DLIUYBXR8NtIwY2sr6aeWCeIgghjAZx0YXRlQPxtBWDYe6Hf9E2OTJsL72BpG73u
51JNILxBuYHBfm3D+dgfxcRspS4NKprY4w90gbAOU46ba18TfXo+HKhD1RxhzW9a
DjKYJnq0xWZytLno5cEsIMfoWowLhWGKV2MaY+lnMFhjhW7k5LfiW8//OHVfUykq
GIaISyDjtlxbTPuGjx2OE/FN2ZbQkzT9z4fjJTpsjMfJrT//PXPUKaNicWRy873j
Gf5a+sgtitXXPBpHJBy2guR3c8WH851pu8oLTlBrSSi6b5ZXv2LH6R2WPDnVdxMG
NqADDLBSGGoQU3KJi8QE6ziDt44TyRDzMKTG0BvPqhdNuuT7AIR64OD2sfjyF1aX
YcuH8f/4yZBDJ0i/pwtABLX8PzSe1roT557a0QEGosP6nz718kBHQYTD5cHTgh8M
hEVi9kb8huKeGZM7lmQHKzEEQpRgiRy/22mGBgwM3KwhwSFxWXAmbp0RSx388ODz
OYDd7SzBADtcTPFOzgv2KDH58G/kiUl+b5UIPHso+9qzmoVRJCi96AjZq9ohbIdN
XxeJx/y2w/3FTCIWw3ooGaev/Tje4xdiPiCU0MabFFsnGio3CdMGJQiO+GqMXOO9
TkoLLYvo7K1CWtmOSud4cqXKAqBHxkxGWUi3p2bxyq7INT+3WS+Cq0EFQvQpRPGz
Cfq1AbOwrx0XTsIKzuZyDxe4fxOVPjnfsPi7Om2HCw7KTwf6gNRI7W4fQYCcxMTO
FygJW9buEjywW6LsjNVvB3dyA6Xia/zTCWY0H/0u+Hv3qarGmr+cB2DoWyzQLaH7
BE7cEzDQq8KetkE3FptqkrMx8AQuG4KlSO2ndEEh7x53AqMUbcT2l6Cfixml0bYr
mtHjKzLLu6U+mLkKHPUDqWU+sKVB65fqugUVR288Krv4nBeSVDqat9/DfxKhcoJE
SUGr23mSWZMJjlRBwHkVuBn88XdI33X3P0il9Mow6XGOLA+pBS5M13CJ+yByQAiM
4sbnlV9Aeemj95j3ASi6V5hg9/dlKgG5coOUakEJZokjT9Xsp0VYCICzmuRliwkL
mDRIN7oGWhIv9DlJyrH/lsOrXY+XjodmsdTmiQflbBrxaikgRJo6J5aMtP2Qv/S3
KkQQfJTAW4DC+Tp3WrVwwtzt0ZRBzPteuzghRgHWn577dBOszql5wv06di+sCoMp
YUx83StRS2OTK0on7nrTukWgfBroPz6C4FVdxASYS65qaUAYUrnkym0d2EzxNcbB
kHWsPQs9AMRCeHFRJEd95EmKOw2od2q9990F1xcvxMxQFBchWfDGWtRfgp5ZJ424
LB1FZyOqPysj/CKr+o/yCq+mXO8CBjmQRpMQGDp68UKgWvV6X8udKVPTInEo30+D
NSX2Q7isouHS7r/xYfB721RyweleStbV768RPAe8qiD8ZE5U89TMHO/qdGaUa5Ai
cN3ClLNo81P72flZhbzSYw1eNhDuAn3R0jq8b6AL/MF1F6XuEZnHSWY05AqdLB6O
3vWkYt/w5O2NXXuotvSxQEGS0M3r6sxMws346S7FvWHaa9haWNrpB0i2AfXjFe6P
n+9BaGkqIf5WktKZK+LHqYTxImsgm2SnV0vsvgTDJOqpST+jrNDXetA8ZeSryzpx
mZtZ+mKqL9kv6FPn15PImarJ8JU/X3KSuj4xpQZ6Jt/kcqcJTszQMJFUSJzYA4Ro
a/VmCbkTqa6PyTEKAovy2SfvHtYqwEbcpKo5BRtMepfTQGTVxfPAMcTNcW0jgpqY
yuViWGIO+G7jhoRCz07H5etYCvwOw6lTer+FLaC5DdCvEQEGvKfrVNM86LujuDQS
zpreiu7LkUsZ1TLYg8dhyKWjBtOGFwSH8Mtnlhl/XniQj5N9ribiTHKz/gL+n2mv
ZpM9JOGsf2qkZRzU+EGpIGisYy9ue49DMp6mNNNqanuEloLparEdkjTzFbteoMZu
ldkMx4TP/d4dppkZNGK9iCYLyGBpBpDcrLTzP4v4eHvS3y/5OaZVLhfACWreYsAh
0KLNcEsVpPaqI4pM8IiHC25VjNABndhvbAjBOxZ3QZmVS7Z2O13ZWnApjiaAMZ/r
X+3kHfjYMvO0lSOXC9ltd5mOX05nUgZdhTe4aFMIppRoBVn46LUxIJ4rSQdElQ6J
afEUV/LzGOxXQb/RTqGZn+JV07IkeAQLjRv5Ht1qc31Rb9WVq5Y+fwFRRNg6gGSq
K1349WwsKuge4Vz5NMqombofc87qd6fnrDmFgT6LNU72fhHEENCrjNknVnNVjn4c
ikSe6j7E01N4wI85l/8XEX7zWrz6OEvlMeHiVvgHiyrBWwB0wMrfWtxJR1942HcK
43ZIY7c+erY9R5vjV9+Kyh43XnhOyRDLPkSoVVf/jl80cTeQRt24SUAreFQMkDwK
dUueEgZAeBrEdL02s5CU+ZnHgYvpSG/2KFDW2u9F/gkP7juhjxMyazQn3wOMkBK8
0RiqOcF/5DBdygQaaga3m+fAekIQ6gXRgLiBL58yIQiE07ra/GjJ7M1BsARiEM2U
bfTb1Zs76tqEOnV42T6GAZw+kQPQXPceA7blMxelxpE815IHM+F9dUl+9QlO/Hze
ddrFczPigKBlyMfyvfTs18oJNhwTiRkTT1Q0hpoeGxs0/MooH2Y+H+g0MI32fQzR
L3LWR4Bxi5NPN3uupAFzMeBV9sAvl0wIxfxlvGhh3QbmI/4jY5jmj6TSGt+tIyAa
owWlDOdIbLvktW3VaVP+k6FuQzqexcivTSUPwAercK3bajLp9szk01XDcVWYv/Zl
ho6VGeXxwvWlK/axfQBDGejd72hCWyZimeZRwZxfe2OAVgK8RRlDyk0G/Mj84yDg
hvy2gmA3a26ieV43HhEru8Ak0Yw0c6KtAhTaCV3BQrGAZEnKCNURdnK7iXp/f/lY
8AZT1HEk1raRAY0RcZvvKAPRXpxSs7NJRLpoPNiB/NA5naim982IuL00teqJ+sdH
Fkr35d60xLAnnrWb+19ED2sfvBMibjNxoZOr5MWh/aAS3h/KMYfWbup6ohDvPfkb
fiPVSX34Cdr3rD4xCflLYnZER2SuVeO0UxyHEbfPuoiHQkCsmgXOEPrWuVvw0ZEU
yIjiJO6eu5aHTJcrGN6Gjr46zfM8qnYSyO/VR8qX5T2f06I4xV09PIujhq7DwLQy
+7A5Ajcc/V67Yy77qLtqyMpnZKmUSG6+voZFMJ+meiXs9IeCxI62afAFQA9tAezD
RKRbTdBX9CGrIfstjKj0Zip+6buUMa6ZUpxGCQXJx6YoSfmJwbc5cp9/IubqI//Q
98CUiHHKaHMN4dfX4tEiLGSW7Va0egAKQFqf37F2AWs3v8YkH4BLLxmw/JZP+MQa
p3AQ1exDkwB2WY1v13asifWV1vk4pPMXn7T2B0cRjjqhAK+g7n7oNk77iUNJ6eHJ
E83IqFuHGg29RsZ9wC8AR0jYWc+x8VD+KGxfY+CuvwYmqjuLoFscvWwvAbRDZGWs
0n6i17wIlxKaVBD9IHTuijnfRweYwv223o3jwNlKqyZyt2LrMo9w/tOucwNpDUME
9nKbd6tOoU13lYGCX+i6UbkUvekuShzTYVhDl2FjPfDR2YKnVf7PCl+y69zaqTQo
GBWeQRvcsfrHIXZfa+hsmzCAAMLdaHinnWdheBeM4R5JzdcIGs5NIU+2CRwNHKbR
Pw/dJYZ5nyXEAET1ePpYIBGuo+IXMcjCAkpUanRFhbjMHnV3/H+E+vvEoKpJ4OrZ
TE9feZHJzZWz0MeW4P0CzOWwCGkFaRDR0+2htJN0TbFrUAZHT//jneShfmlYPf5w
sJ2UTs2M8Go4dPv/na5RlLCWL43EsfkddERiYbzxgzIszfVGt7KA5ptbTku8bRg7
aEme0KjuurvK8d0hM+p5q0zEjPuE26PWzXrDZxvzZk49A3hQc5vXQWQE62u6tMOn
NNO7JZVQEfZOfWJkUnRKjaZl1BlsdpCRkyyPsPMNFQPxxsg+Lw0o12wI5xhmim2u
iJl4fvoE515lj3dErAIoptQ7/wt0VvHLPe9jKMdbWVphJL9E0iSHvhRhYxknD8Vg
cKYaIfGkazch4mD8gGVVmTf7yxyCk7NMQiBgA3uma1oc2oc3b49npOgP554TL2up
+n8vgqZvuPmE9rxRv+QJwXgO+2rFsyBPZ0fxAatSidGigbxQYf4QhH93FqGMFp9l
h3/YtEsR7rzMjgZlAHdD06b9dJn+mBTfOQDV3XH2LIZi33KuqCLbqy2Rn5GtnwpT
GyIz4sC56Cj9QC46UHP1jV+IIE/AXNyQLohZ++qufrt2ufdBhEjrlHsnOXT9wxd9
owjLwdC1RPJT+SkB41Ku+PEiHXOeRptmTgit0FVLVLMzPHAnabPujWIvtknBka9a
yEEOCf6SP80cachYgUVjxoXXI8tPkkpWytsWcd8L42927FkJ6O73AEuDnpeP8E5v
17whzK2eP7gebSWLMrec8D7KWqLSwZinPv9s5wsoD27fc43Lx+y4JX1sfFQaTqWB
DTByyWmUyfHhn4AHtc0DJUfvN/6Zt6l9AXDCs98aJxvM5YS/0W2J35p++hT/aq68
3gxMnkb0b2jnlLALnchodddqdsUg2bYF30+yDNiTiltv5VAHSEjBpBDnt9FFlJM6
y/1pt+ZMmAEBjjhjqg6sTbsHTduI1aXNAorMShG/stpTubOVKCRvnyNIwItt/9AT
7FMO+kF6VbTKEabxUpm6JM+SO0weuhW3c78eWykZY2TdeVTtcBCHyjqNaVyn0xoB
rzGajHxwUi17f17D1shm85+9nWZ1dCr6EwN83MHmH+gcS/OnvzoZTkDYIfgoHUrz
OV9r8X4iGePGi1ovHiwBgbAPSid/bGjQHV2FQY/63ZqSFj1MeFH4Q4cNcUDkfmin
/kig9FWf+rxnJ/mo/PF9HC5L+S2+SAztiuLsJ3cnSoO/k1Ite8o2PQigO6Fn9g1z
WMPkQHuEn027xAkG87EYT4aoN6lHBBRvFyKX4RZGf9hXqe9nLPRJLHZuT35GTXhw
287t6os7ProH96kPpa5Vm/6iy/T6QPh35y56IzB63A4yhlWDY00y61Nhuh3+XimI
kZbeDXqVcrqrFZV2P+GxUs6Pjc6XgtqvO0kMPVneKIShFLUy3W0q8rk+5m18bqd3
L0X7O4npw6Lf0ZdtfonwKUFzTRZ9/H0QaVgJ1PJd9m7XNHJBwobxU3l9jPkqcsov
xrm+NJjNmFQVHRWgDAHXRlTMGnhkJ2N0sCmrMak3X6Gsg0P5cHp/4g4NvzP2TXk2
GKCkkGkKxfqNlCmYROhWQg9a0ltmIBqZRmwEOis+1ZG9cL1X+KU2N4hBZr0IeFVJ
ShkBMJ+JanicgF+sAoVsEVClQlYi8stFa2uNAuxZ2p1dN+EVFS17gBPLuQvYfM7e
4P84TuV2Nu7Eh6hkhZXzEnGcBurTzfoe6h6iAdMe/ulLdbG+WGEUPjAhj5JASG81
FrICuaFivsWPrcnzEKTXPTlh7/o54qDf1/TCqcWqvqKwuu7sswLPTjySVQDo+iZK
Gm3jZIrtcfX7Kx1zmsfwKwE9oGom6pX7GBs5MVuPKbiLqa+UeuP5Q4NSFeeNnOl8
Zprn0pIS2wxfbi9ARypxa8MQ/zE2kiGa7s4gCD8SN7dnTO6ZVaGH6OqZVBi+SsMU
9ftawL0cb9wXoAIWSl1P8HVKwKTW1QVAmESTFwpR3GcDJKfp81oEnUrl/esHgTx7
iWns47YfQttVIFNtky3MtVCWTb8thOMFbM+S9fWd/Ix/FDivuD4K+4FWhAK+3Imx
ztXekOqXUx9MOWL0Bj0sxRKCjZPHMmsO9sGryYCpbDXBLE1b6NJEJ/LRIpMikO0e
7Bm5FkgMaAbepkq0H/aVXninzUCVvN96uUhQ7xWUBdfw6F3dy9eLgGCsRAPRWyOZ
AHC+JcmL2ZVEV7huw3J5HYS7sqCoAz2dwy5cfPxEln/QHD2x1X8XaIkZOXnHlsQi
w1yOonwFupScHQR04VoMVq01dEyEz++bzrK3SvxaUinplCaX3NOoPhD3jgv4BnyQ
yU68VmZ8Kh/Gbt1UYi+9PaK7J2Ye07io1hqLxynOwvYuYO/gOiu9wbmHSBm3E1qW
v8PZj4K0v/JCdCPbDcB9UlwExfyMrvzAXKdv7HMMqYAizkD1qDs+23vr5cozAuhw
d8nyD1B8zsf9I2unhb6IlA8ZkuyI49DdakTPO0DJPj6K5THyR1a7maOgYUSNopJb
7bwCHSIJePsa4uVfcTxPmpYIhu1bqg1mIp5KHh0eGWkuJCBp9GUl0wpD7WBTXytk
7YbbusNw9UOB0Pw9/nh/IJ+yd8jWzOdusrWvdQy2aHtscM0Xnri1IayxoB1LQ8QX
0EeAR8UooJfV9bXExmmFQDcVD80ZkhlOUnWmWf8utGtG2BunprKSKWNJvlxj90fU
JcC5zcNi+wmmEJ98Q3MVZEllS3kt8HDT2AdKse5Ste54mZxAZsXQ8ToREm6/zJMg
lNlz7YCNaesJDJECWYu46u7PH1VUbHH/IVtKj3GQ2hhpJmIesG9TSqG/dgo+kcb/
6P2ray8uAL/UBcaVcFSoQOw7uwYCNdnQVsfk0Nz9IEb+csto5fqHkqTSNURN2dNj
VQpm3dkP/pPZokgxBDAlTAclnRhCBX+uDb0RFH7Gds1HznTlOfRYY7b1rzKSO1Cp
05t4z+C7IUo6rJwUCeD6VjLVTLpKk4CROe2UKZuJOHu02wgxvOV6c5rpf841haOG
otILiKQpGSmnEHT55527uqWHW1ZFU6XLmqhKZY7t50Of92uI5I5Ge2p2HPpInWef
H/ejbqie1jgcMLpgy4U5apK7D4Csw3gBbcKAvJo57mBQWkAHolkgERjMDeosTH0G
SjWJnkzB4B30BNhQkM19mDUU0vQObFOnhS3Xdn8c1oyvKvBn/OE0GtDkF8/Ca3p+
EYBScrBLUZZzrcVp49jQ8NyldH+k8QSVJeMhT+HxulNxb7WdE/YgiqgMgsHMZz1P
1dbegesGH81m3YmTPdgstc/tYSoDiYVw4Y7HwTL5UlMIXV6eSRzBlBezsPT2e60A
CSueEIWWSgFjvZjGSXWFCbAVnsF9ZEIqbog9ZASbNg/K5totdeOzBCJiO78+gxrY
BiKV/Zwpf4YZZED8yhbWn+c6BxFNrduzLnnUpCDfOkj1owCi/Sbcx07BMy4YRpHn
DoqjH0hvrt38dBQFL4wBPqqyS+wdCFmq5nUeAkPgDIO7AEW6j4qnPnwiv3F/EcM8
IhP/gm2GGwO7dhktRqOZepifGz1HedzzLVR6LNtD2yAkJrOqFzCb4+53xdhcyBko
9X4bpCvgawgkeEMmnemsyvEVOKC4fSWCCCywFUokoI8qWCbqNLpoFkc7bn4HMtCr
xa01OmbO8kBPjt7z+xh4pWf3+pVc9iEyw3dBnpaXQhne6Tv3h2D7SbEW8yaAyXIt
VJSMTlIjG7e+Uwjyr0PVeC2cgMq2h9Ek8YpYq+WnJ7hGnqENbHLaB0/WZlO1l88P
4h9TlO8q7oRuZhaY/VPBkfwYIyIiL6HBPjc9UtZ/Aibn6ut+WT7pZoe7Cv+QEyIT
MEIywPTTC2V3yvr6sOlwbp0OhCUYUp53DiJVppV+yT6jVYqBFjxDmBl9FCbwBtie
3K2YWM46T2ZlC9GXaEhYXJZwt8fmK48/Vx97BrkyWHNsUzh6DxhyT/KuTdpR4wRu
sUxDHo5g52qUlEOiZepamnLIzgCS0MXVV9JzZX9tLujEskTdLgN6k41mxhPN2oKX
KaEIP9kE04o02TEtWyt5jsXa4fX9Zq0ntliYRh9AzCQzO0KbUXpjIBW91DQLKCVF
yq+lIHe3gNW4mSkdwJOvaepaM+IwBy2yjDNqaN0Htk6Z0gjgNooJAI6ZRiPm/eHD
0VDvgaQwZX26YwK8il0f3prxIy8Ny6xiFjDXSEv3iMfb3eJb+tvDjSkISyRiUf9M
Kz7vbin3IWTZ+i2fKSpj/o/6T8Y1qeD6LJLpbLM8WHO26GF8BIiqKsihXZHZWQWr
61here5HHtDWrJkD65VghDzNwjb/qyF7atI+BOFCBqK4Fpp8ImEDX1WqMR5ih5T4
pzZTp52jBngmWCPH4/EdDYaXZGwY+boY05xUyoGq3DloWvB8ha+KtSU3+srotaxP
M2raXam4R36FqyPZZ1o3oKrgl9bAMCK2ncHR+ycb/KkQbMtBPFeYZ61cD5Vb4pdB
p+Jm/xxvMrkobzH5mzuqIFfqMNlcUHKgmTtLs5hIvnPfJUJvCSgq8Uap8dkgDnvk
CQiP5kdJG9LRlYWPtgHFez0XAyxnRCdTag+qzykXiU8mVJp8zMkDwtoO3LBcgOIP
NRhTCT0ePt/mvf084yp73PEHlJmES8K+9T1Ux/q2T3lzL3V6YRtUGwr59Ur/qWBI
UxT1LRtLARCWwEBmasV/2eNtIoP90olKVx4P1uKyXTQ47Nja9NQN1EDnNlEKd9id
KjYSk7gh+3p+kNb97QtSKz/pVWRyUXAciRvYt2uUSo2td5rebX0Hx+KsQqHMK12b
YKaP4t1+vTe3t9uoGikh6daCjW2REKpsr1Iif8rQzcupu7XxbBFakAc8xu2XkCzd
ascpHE12pB9WBqmnPO6r9kAnw6eL9FdqOZCsi18xJ+4Btj69QIbBEGZ7jBuYQK7m
yWjajVbr/hHdcLrkR0DE7+G2GSTcwozEM2PIJo9Z+w2RjJUmrGmHvZqT/e+MRkOT
q2M/f7cQy2xIO95+/TfxPAAMVW24tDe7faWOcMovIuSq221GNsgHCG2lv81mpVUf
JyAWV4XmpKut6VW7dEwbK+DReKvJ2ln1FVhUcCERQ7UI4beV7ImKTo+qTAfEm63F
Kv8lEvRb2s6Eg+JZttdIy7AyFfYMiCx3WLjmWQ+6eNCroWGKfZZanNuMZtiy9Y1k
Y2ZDqq+bwsS7anwOFvP2alq/n6EsEiyKCRnpsDaXYfJ0Uf2FZ33cSJNou6HaMQTn
WljBzJtL3IpRl7AU4WaRXtY5dmRnvNlGU9UJhlbuzYCCXZI8nkcLxEGTatpUDAY7
NUMsvvlh8uWBy+hw8W7F28ZrUEQ5RqB2v4l4P36RECthIF+o3wGrBS+cwxbIm61F
sk7Lm4jkfvjsS9G5pUNQApFB0dcWwk2qPMajZxNAnqXcxoScTqo+ScAAI3u7Z1W3
s+Ts597ST5q1RGob37Ey/gxhQD4lHYIpWoDIFXfEzEmai54OF7cDCGWj4c+1My3v
yqvgPGm3qW2FztClN6bHk2y+0DCd0Yz/ktK6mMXc79thtykSQ3cMa8gJ4MjgmSAK
QMoRymr/fnlhgBQGC5OwflCadV3JldBbNafE8OuPtmMFc6nB8B33fRtX7pdKhe6P
zQuL9QCdUnOO0Yr6pMKWzOiEEzYxrt1S8s3sX85/oOSDIYOMUlZmCTAMsXaIcWnC
wS/ZTTQYjj/3rbUv+yBL0uVNWaM0lmHj5Ygqz7Fic4I3Ro3SfMi7CuJg6Ptb7b3Z
p1JbDIXB49hQI8RF5uxBAJGyr5SD+Fhia8xoWhnhOBsq0+nYtsVq5jwc7sgCRwhS
ZupsV43Qe0aPYjfNGhLsNRA/j5hyMlWWHr8tfeKaqo1ztNtMZMiL4zW6pwsvrnVG
5fyHqRsxGu9gfI2QzCZu0BILYABMd1upEe3z7s/4dIGsGBzfAykQqED4xlLU6llR
slIB7UY1flo0nZyGETWtQylQ1B8mVWjnE10pKM0yK99sIXIKg/mNwHrE4hvyz3ix
L9p00z4EwxclyMDU/yjj1n3ulcx3brTKKAQgaz8DJkL1Xpx5gKCs3acdUBfVyIsP
E8DIXErHE8RqUFCfvS/EZIABNbslhtkp/vYwiRUsD6HjlDWz470r/v+N5ccTtNaf
uCaZQ+4oRoC3QKaZMC79E8s/mJO418DcSL+nno+gi2xfk1495a2WP4wCcex78oxW
1Ej6odAFuSv4/gfNqy2BSN87whIZxL7CsETjQUuJ+GFHARZbW7Q6L+90AYRKHaCG
4q7hOakhD1nGgF+t5scMDTM0BwRhZdLk+/aURa7VUA64SqducPoRShtO8ULZ+TCC
G+jAQyylG0nfZSh5qSP02PE+BvXn3b9LhiiNFvebSP+knvDuhQZXnKSMi/VScIha
KGDSUKzsCsHkOTva8iFM5zlgkKY+vuBnIuW1DTMmAmE20zuvXtlVThEULz2GtBP2
6Eou8MwZhEYrx//wJ4/OP7BGfadfnuUVKyL8KhfojAe/rr965gULM5zZ0drbr8ga
p9mKpudsRlxDBcHLpzII3/aS1cvbjfqzNV8VxPAQzpwprsdw6f3mbINh4RN3IJAW
Fa33SH4d/fKZeDpgBF3VX8KFzRaPC5CvM0zkA3KvTN5k2WSGx49EHdv2sbaUBSBg
liu5dE1uKgfwpoixTkfs7qgitvMXd1c1YkNJj92P4xl05szOafsLrDLfA4qVcxMc
ytI5fOeExoLZwMM0RNt0SRHXzlkWPmi97kBejpLQbjx7bLaRx/t3oa08adxOJVtf
7qLqTIlsATtuLt6lF57d5hJWtA1GXNqjo29Ej50MWod5q3Jfh4BS0Kgvw790Yav+
UEu/tuh495LG3yZsWwtpILuF+vVt+t3F50IAW+vrEu4WZjjjDWxypUKf1Uabu/4B
o770CXQSh9qtL0SsNH/iP8SMbUWX+YzD+eu7O1MrrqavwOqOdb5e2YVzY8qJ2xFj
SdHuigkfYN5dwLCf3W7fBsWu1ZO2NQRpXuUop7+XRFBHKmfVsGKuNYzGT1aDsB89
VSqqwOy2FyBsxx4WULAoRHJEkY5fH8+dg56dqKfAlGCpyVHYvNYnp+yLNIyzCF8T
SBnbM0Cntm6gvS23mxHWt5eyMUS6rs6MOff+pKN08pPfYU+5Ujc4frVFQLvMdcUD
zDb2kqtIjmqRknnT58w61oGo8Mb9J6iNUJnvRVEGnKwZBssCpw0GDu18qc4LYyCs
8ehBZ3frdFbWrUGpbGq+Yq5l+9bLU4ZEfkINp4/0NN694huRueBjVKWtiDNoJ+bn
71BkLgGW8BPwxTvR6Y0+aUa0KtJmzEx0FMk0soZ/SMMpC3Opf+rnm2OERIJO455H
x4h9fo4qfffjfH47VMSo+LRB1f//zIvBxTWHsjKKzXoo0Su3oB2PqyGLG5wl4h5e
CLrTYHOpkjro1F9K87+W0AYSJWhcN9c1tyryfuWd6qXmaGH031DlM0VABE4tC9/3
ZWvTRKUVCfZ+F49VZavrVywj1ZUOxJoyxjndPMIVFfgvedAQyq7C/lM7Ts0Srx7p
NFY2dTX6BLKGNSIVGk9JdCGJGrydUj4e35dpChnUIArVCMcp431Ist+aeu5XxpEL
SUmXRcgukl5bnxkqUPpXcUWJFg+VDw1f+iQdyNKZ75qIEQxMm18HnxYufJBQFAHb
m65Vulg4kbA9m16wAwzPAhKie4x2Dto1IWj4Wt+mg2rjmP5A4XLPrYjfi9lC+buC
x1b+iDTjFcAhcpKSb2UhI1MXoDRwjJChfkiHC/NmOll/itmNsScIxk3JPUaUmCwF
nATnl2kAWo5F0sv3UqnLWbxNjoDrLKDzzZ+IJiP8ozhibiHQ+KcBbC9vQZGRxN92
68TtsyMtcCVE0pOaeWhtaRoG2OQ2Bd2W2NVzBas04By8Rw8A2Xq4tkcSC6mdEGj8
MWbHDjlKAbRfR3XtlyhUG24vX+L9slSdKhOgie1GLw6tDz5yjc3BfbMV75DkemsO
Np1Yo/bl57ZuOB3WVYgBuohaKfkeLKBFb0MTzJDKBvemSJysXVyRr5YIlfyLAJhf
jgFcTZsLlfPStoC8S5NfHHRp2jW0mlOIPCz9WRmYt42j9gYZTXF1z0wJOhEORVUv
RoeMH/IJDqI5Kem43ZOXn7pTPZ27KRSXFgiohQ3YDFQlVMpddd5kxJzlyY+Nk5Tr
yZlW5/xshMtBZH06SVupbFimgyXfd4SRXEwyXGsm2PHy6ql4x0EtnMj1w7UDwq2a
c8jEOWapcBA4gffvAu762TODJPnghoK9l4qjr/bni+n2lWvlTLxy8qsF9VAEfM4B
tO5AyvRQ2WkWXBXeSR6902NLEiZk3ORWeEHW4WwgV4Zq1TYeQ2O2dt+7+Ek2ZbzY
p8lNzQaf/lnHEA8Ax5BJiptSPrPLfENNwcBW8O0oFP45TrIRZV32aBsPcNbVofWv
4fa9GZCclWHImFn0g94uUMYMXDE/lDLviC1lQwGXVKCz0adE/HFwilxRsDHrIfV9
sd7RxtqArcR+qYwKY9qi7h7lFwnW401x++/DHptcDim42ew/dqeP8pjWekze72BO
X6V76xguJDnCBptNNc4DXjoklNr/5lJD+YLFsI8sKWEp4RS9ztvYEmxhzzuQo+TN
STSAgyev40eUdLPWySUTHKpTN7ggLtSy2YyGpQLCPAalKEQ2VMA1NBiknXPLvvNz
f6vyPL8JdzXUlvTxB2DYXaj+g3iDnA4jjmFRQzX3zn5B+NT8lpU1fmeUPlgQ/9Lg
w6o7Q96wGExYhzaxm9VQKtSaJ5meZRlXQlWQnruibcCwF/3iLsJLDIKP2E7viTfj
IQDgPDofyRG9vzvN1thWM8l1mpkP1NNATn6f1mKpFy3OZyZSEpf6EWGrI4wplx9k
vIMvyi23KWNIVNIP596z9JyCbBo6SLGGgJe//ZRDPpazvKbWwiOO2kBASXRAmBHI
8cVz132p3jH6r8ajyw48066Fe9x7CQHi/V9SzpuVsR/d5gSkldhMa9YHOU4lzllc
nXNKf1f2VFGu2piDA4R1O8YvnI17Hg4BwPkJBhiV8I3vJZTjxhXUH/zdcl/plDl3
2aW5dR3/aUwCPabzJ0EbP9zUBxzsVmRyJgzj42CAxUl5LOcDVsHTYxGNSxk6GtIA
ehs/MBfxIUK9zBlITLLft0jOTZ7yken2HJKyqjK9u9atmn2Y9EzoTO0XjmBiP4n6
stJq1EO8W0R+2ExvGBjP/9zhcfAq2JlNToR2zstNCtHrNzN2tHVAPC9M63oKv1eX
l1JsVDoLixJkFciV+pwvKP7Z5n/7G3DJH49nJd4fGoF4ECoaCjiEviOvyJ8bruJY
L153eIAA7PGk/H3QjZicTffj4k97kcat9i4jube+8dQg0k/lBZPK5kfBOz0BMhlV
MOKk8wQxzvc0oFj8B247aG/oXhzymDM8JBtV0MtIkQ0B0pCVekNfUPGj0nfhz1ym
uBbfn/hmr+jzAq+82nAJ+PhQBkUckee4jZSvk7TkVkUigvnfccXNZ1f50Jx4KMtD
tUmF4VUr1rLR5OBKUnWAyzjcSEeeL3gCzOUJEV0GvaeLmMv10BdGAEeYCA/nxZs6
QCEowFoW5P/953XAd4uXCkLJq1W9e7yUCZFPjDAnPsA9zJhPC5QcYtbsfIAELPPO
2CTdo8o3GFdgEll1wjubL32d5nHv9wilTjlXhrjveI1TVowwnKNcbNekrVSZ8lji
Y4mVycbJ4QfwdVyJe+QVbTKyYLF6kLe8ITxFk5WctPjD/RqocG7c0KWxPle4VpPY
Uuih7N1eDejyPQ+dr2uJ0L0ZLF34AK5DcYv1VlxIVlZ2A01qeBemU7F3uDYF9X2R
H4q41Zmwe0ZqLqLiFoYM44FVQjU+jPjq9bPaCjmrQGuJN7VBDwVpd7QJxhunpkW+
tzUhMNTUNFtuxwThauhqVhHHly3xKfP+I8TDASlpiQwaT8IAmKY40rXqOInOHhJD
mWRaGFSZ41JK+DVOXpCboThI82qxpoNg6bW2dAghDO7tN7SU4ZbIa4LQq7PfppHP
izUyAyXlepzBcexkhyyrRAKnUQkZS3fgsca/YdZAO7fl2aQZaPq+jdTVVYYwe1qy
5hN5vzaThv/MeR9Q7YehzxrsxTs2aVnq/XEUgxENrabg59xIeTlQZbkJVacDq3TM
BRftc9Qj6CMZ/gHMQN2v5lDPLe+WTW1lzlOFMl26GvYnyWLls1+6+Kohq2CJv0Qc
vcLEYVKBPR/JamBDe1Id+uKfhzPw8nKdu3xHe9TlaM8ewQVUmdSxEyB9PMyVz0Ki
WvUaJF/jw0cKjXzuBVr4x0M+TwwbabNwF9l0bM2nmJlKjB5ijTHMCt7MRQLv+mJ4
mlb1fAuQHEMyzeHW39Ia5eCxFQ5neSeZ57QKtuBHWhg4+4C7sfeAdr6Nu+M43mN7
beSqHFO3Tzh89l05Tv0zsyVlaVhTXagsetYp3KWcICcjjGh+obYyIkRdykras1+K
IpjmTbZvJHs+yqvUmq5VMXgVY39HG3xcfWlhLiqyJEgnomT8mPJ3jkAlsVr9UMMW
+nDmOfLn9RbkAbAhaC+1I46VMgcOfUtwbtzrl6dCAgWOUNKxcBj06ZAsQ2ssZygQ
0c8a1v4m1TQ0S3us8Rk9g+98lswoxWbpwFmog3DQDCY4c8gX9bjgiO1sVMXhJqql
I4hNAnGCZ2m1RD3H/iOUCkfnQrvVMInvyickzowb4/YE65x/Il7IvHFSlKFxFIj7
eQKanxEjZ2Yz5RKYY72WVe33DkyDTJfTGE1KJa0TFTWanTPrJBbYVUOjD8i1TNXw
WZiXFLeIAPpsp3CKEOkjjR/QRaAMaoeD0nb0n/qlSjQakyY92dIBSagwDQzbQ8Xg
BOdaKRKCPt2yrKJF+wnfBaxB5h6ORRuEWDPwqQEhKnS+1rFpMoaXtTPGy0zwjjfp
fP2GDsgIBMh8X7KPQXfYyZLGDkoATTDTSGAtWt2jXiO1X1VRumm/7reHn3DvrI4n
6v8yTHDrLfg1xZoipREKv6x8WOhqktx3skzUnEwprQg8d55YJEpMbgWeRwgH+JFe
0PKDCJptHrwOea6k5cN/P1pf+yEF9xf92E0oyTsOFayiBzc+zgyv9O3F8Jmcgt1H
8CSWqDV6wvTOPSU3gKENWYpPz9vW2nZcGzNSO00oQAy7VCmrvGbgkDuC9Qe+6GyV
rLBmp3a1J7maQVz70UYbE73/HBoaNRi7Y+xzOTlBBLGKTF9aU7K0GRCKKP6f7kwG
7bWnugovjWSmjiXfu8exv9VDjoVSiPj63Cd/dyOVf9DpBa3fiyLJ0SULiaQYCfJA
jaw+ExGQk1r9XdAF5sWMbCN11Z5Lv7e2fVw5cS9ZqgsgMRIjNOazLrIDyxKva7E1
LwtDexe404zO3AkYExb69KVjjZt6O4siLQbYBZNjSrnbhsuOgA16ao8+vniRbM0r
HBYXIvlgHabJdFYUqdcXgk6PGafe5L+o8j+RH6Ev6YJkIul2vrGSq7oq5pFN/pBo
O4kKsQf8TJvasng6xMy2hF866MzC7i8a1fOrMv9yXZsohtYLmthTwuj2J4FacMun
661Ad9XcaxGL7iYDvSY+jRZInvLRaYv6qk9vKYPNNf/U0c9Noof0+L7/pzKC52k9
S8S1nvkrOdF3iWMq2m+KnkFrdlXaoETbn+7WJf/Js/ONZI2KV1oZOGgwxmpVUh86
Svm0AnuLY8DZeTcPgOk8M6LGQuz+B5rOCupttQRHFa2BPc5JQBeGHMM69UGCKlac
27jhY3Gy9rC6b+zFoRs042P1VY42JWD3EIaq2Upsdf1XYdRHi77J03YPEsWVRPO/
vp/fpvJAFfhxJ/7v56rG3/ykT60E4q1/bMP9Jj37mIwkLXooTnbef4wJ8o+lD2zV
qJDJlVgpJ1F2g0jTFD/uYi+vjdDc+Yn+vyAiT+9mT0r1SXYTctLj7J+lqWTiqAqE
gq/SLlTnZbZ0WGVhkEWF98Gq1H3B6M/ZFnhKo38ADc7YPPtiK/J0E4R5MET3S/wm
inbHst/H3ZgDDgw/oOZJYaV9k+lrU1yqbzoNHh++Yb23FjdvzWDPdN9bQ0fgPy21
eftztnAZ6/rev2b0RaQ2SQzU+WWDNl9R8Gri0MYAF+wAfPjuc7JZ2fAyr6dqt3Rv
I8MP5rzDGC2EGBSudu6TuXffJcP9QkQGjB0Z68CIf4JcyLmGLIzgaVhIpHtKmiSb
rL/I2l7rXs975vewRPB70K7kupTtzwpGK0IzfK/mo0cJgufbb9EHzmAtVNx5R+0R
8WhF3lcdHsTAxvYdIZsEwtTxCmDsAIu1ROiwla3SjnzjNMQWaNUnaztqKyNSpsRc
9Rkpa/+k1tmljWK94lJf3CA9sHg4MOmu1GhBzkT9CQlxzyOXbG7NRjWbxFpgzcEq
qvWvjaAZZIlgP+oePEcK3CogdWv4nipDR6XUOXmmlVfoVzBbDrWRdv11rIw44RJA
fk477OcoI7j98BNnV8FdeCpt6UEKsY1cv/kHYHE/5iXXERH28Nk0HHjVzN5vGnkc
jntkqzZ1Cs2WzPF2/B9d9WQNLPQP5kc/uMx182xfLRK7yhvk45slMogy3G8hODGh
bMCSU1Ouf46LUjaOPsYgmzD1dyf3825rBfYl8fz2yEl211v6/jTiwO+v4ln+OTgq
g/+RqIT3U2PWdeyH2wVuSP1zohd8BHD5Vni3ZgiJlm5hfSW9gHCdrQRdzQtH3FvH
D+WwmXSaQoAmrlzbZ88OlrIr3zjYtiPurkviW7lx+CNEEMwXslp5ZHoPQ/113dUl
8GjLsQYImYIrdcbPLoW8Mk3PQ987D4SkQIuP8CwLnciELYmZ9x+OGorIDrrAHXjy
r/IgbqLINPZRaUj9tOYJzm3AlDevhUOxnYFrMOYGSfDw4QLjCeCQzejcVlbG94st
oYERTfr94WC9RDA+KDrLh/kJdbOKz65Asp4o4RSdosR8d50fww5ianZ7P0/U5tST
Mg8SXmNGInnT3K4xNACTyogREpa8GWTt8Acxg1fwdNHBbZiZ58/vyqAxIoiP65S9
2NOd7cIrZfwWadOW+S7E0/GlGixo9DtY2xjtEttuTD5rOylCaQIyA7l+TACJrgCb
0uU8ISGCttSWLRS0PD9J5oELpM4r7AU/ENPEFfG7dAiHg5jLiSz0QGNgs8eH4mff
0KXyC7dvXgXiglb2WAj98xl6Qj3eZbg3sckQL7IA2xMg7V5tKRTorUb3GWARZoKp
iCikKfYDW1IZ5/aokafJV5key5X1X6bJ7llVaVjj6WS2UuZ9TNvAtykMHNBZ66z2
D3ozlDgUmZztTXAEYrF7r6IZZhNq/lUDDjTHMqflV7aLQDmgSzZuU1RvacUkcM6f
/fn+EvXPtzOLzwc94QQEVaKHEzEdb4olSXXkk8mJG+k+epFbCLYZlMQYHKTD95Rj
/tVYjVr9l5bohnGteBpxXx7OduGOQ3A0r5qGcpSbpBiEoc6cjcM9e/P/IvYg/Q1X
E0OArwQ4IDgpN0giVWH2cXe1rc7p2/nuXc7uOoCar9QROQXJw8RJb9IUa25W2gKZ
PqgHWUiLDzClX3FFd/lOAawWSlUyLOSgX/A2ksW39qHj/n3mXcIMskfMK3MAr5DU
PKnYsXA7ege/TJ8Z9BO0+5qeev9GKltq+9rHdOV30o3IkLRZ1vYgu9FuaDHwQtxs
YEGofOwmgJ4y3QQzuo1y/q9wHYQdqz3D80Ys/jeL3JiMF5+PPclyQ7nhWyQUy8bA
/GWPUBx1sni4rTaj+LTOAXWAA6hjdKxdEMbs7pqB9m7JrAugh1rqxXUXry6/X2mk
OxNrUzzIT4GLftRs3tV+bfSAH58T7UirdRIX0yeil7p1ssQpLQOK+JDJp/9KkVK+
Vt5d+os+nRbnc6myMyJXFHpOUHHcECoc2PKgHUfWcXKbOR5CFjyKQkB62qQydBFN
SqcxSuipqksB8sWF5iPGnD/A6E/wLWoWmFKWp+CqexKZHWIai4dX5lLsx8YicARV
XJWgk61pjxfoI52iwlU1p/2F2AN3YWQXtxaQo9j/HRptN/V5xER5GEH4ELtOF0tB
5BUf1lGCgL+WzQFjHgnSVrLu7+HwLAbo8VKDI0kHcUh7uZDbxZC8eIGvJd13gsja
6DbAGQ+aRMjw7DDvdroDGznd8TCh/qdoe2UpLtJu7E/9bcEXCHVQ3M7ANc+PEU7R
rjZ6g44bdkPBlWco9eb5Xc88Jwz3Iz+j9/Ym/yJg+3f4QkpsHg296VyO45niKNlA
w6eGJB5F8X5HMXC/WanxUlA02NXB3ESxOm7oH322c0PZE6+/4xjQZF7FXiocKW52
0+VQ6pfW3Gz9vDuPCpBGzUTF2FrH+5nQx7sAzz92HqzA8CeOzyyWKzWAAAF27guS
m34UvAzXb8jAS8Jes8wHjKxmVEhGo3MG1rEaDl6jAkUKD4je+TsEEGvBIcg6UVrs
DALz+mrZSGIrnY6rCwqgKExhVlUenN7NBbs5cwXfia0AGYGQ0grbhmSNR4vmR8yz
oZVNLHlI6y0uO5S06iMBsE01hi/zbD6bzLjoQxsGE3RsIQsuXVMgYjZDL3TJHbmx
gLTqpVklardmdqZDAcxED0CmkMvlvC2TjgysvjyhkPLDTxCl27U6gyNuTiizTOn4
UAlyHrQGf6YVK1iCJo/PC4PDcX8tXt7LXP3cTmwmMUCgcpJZUYMCNW/qdL0j6fjx
rmMMRU4mASZH878YFCq6YJUDVmrJPPDuMAow2xZMCcl2onjk2fICopaGn55dOJdE
GJqSsW7Rjr7EN1e99dWOPonETMrCuoSGkC2EM0lJ6+7qKZXKDP/LDio81gkoWxbh
8hgJuNljFMpiZaIPI1JFm+K0rCDAl0RlEruGXudQEKMxF2bg4fKbnjgKfsr7RF4k
plSduO/LCUrhacOCapdk/kiyvxXTZDvz5k90sqlK7PFRn/uaLSvMvBYU2e43ro58
3MOAWjd4sIoi+9qya8qr1WajHeIOkJtLmGJmlH6Pj4LfUflRsWmf+s2fyegBHpx7
2huCFP/7guC/YvdtF1/cRi+l4wumRbo47OKkGFSqJzOtDieaF2huMLb8hkGnAmPw
6znXydtG/cMGe7lYYV188TaFcRrBPJnb8p+VH4C/w4paqHNyt108LFrlfkWFCbV4
Y6YDxahdDOKyYc0b6z7CCi1UExbyWjHQ+ut+RrYI2iZ5M68v274EWKDf2N4jrXFv
ZZAYCRxAdl6c5jRGhareQs2lzKnQ7hIjoG87e3mz2W6PrtSkEkTa2BkX+Z6QvqJ3
abRpWebiurFeT8cb3l3x/d0dhis8FDIx4dHbAp5j16Rv9Bv9+BBYsNnMQhTMK47n
UgmPo6B4cArNTYLFyP01pkviMGutfjAFJfNVv/wf1SuepBWotJwm6n4u21szKC5D
naVzPhuzeQQh6OKwuBCbJevWP3r2p9K9eJDhMNL/z/u1H2H9+bvHRgM0Gyw5VFWu
79Xr5ZvsrI37EvUCg9fKfWfk7AIwQVv0/v5ThTKZLulzRapOK2QjFJucnqPO1Sg3
dghXxYdsGisQrpEAcOs/0l+XZnIxdO3hSLCjH9jVszVx6dVh46zdBSXoo5Bdv4+K
dTLjIAzBWvmGR1iBSLHPxiOs7Q2C/XnV5sWjl5PQZ43Vi0un6Vknd9FMPc8nZJ4b
5tYPiypfH4p+ov/FioHdV7m1o8wNUQY3uvI2NxTTprnKIuWma5gxd1O+m+Pocq5y
2+BzWGMNMS+w6F1ya2ffyAkWwCmGDJ2x/5bt5z5q0g+InTf49IrLjRi6FE/EUXSV
FE/fjMKEwbAr/tpiOoqFCWP113vFWfZIRky9t+W8oEg8LdGCEjnOdHCpgRsiCwdi
w9uuxWWezN08aQIOsa+VOzr0LJxtj8vqd8KBbq4zxJr5hUeIA4KdQ7MtKb8Vshva
ZBG7Nu5wzBtZ3FtwMhAHPbwPoDxAQwCa71pdTZr1U0EQ8dDgqvjL3PVOr4cpkEh1
im9I26LN1TCriioAFJKbYzJz8tWWNdgWWJEfFBAHrrweVZOjuR+N2Wg/TX5ZxRKp
zumTKRlDaQymbFyrs1BCYDxJ4xPwiC4pArd5kECKYKiBB0/I1zeV30Gc0NuQYjEW
2bfMHEnDanImkEKlqsDn1W1xOy1tSWxWCDPYyKKQLqVtgf81l7z4eDMF4grAKYPu
5AyQBCoAWDgyiQxrOGWXoaopaB5d/PRLIIYwQ+FpOialVDTWLTOQ4853o+LdvIS6
wKoMX9m4jrs2C5wKXALB6lBuDB7siHmZGZL0j2aG9FHqKpZpqQ23ka1ZYqNZpXu1
SsxnE17g02NIZAdtQLL+nTKl/dzhd3sqTjq41Z831ojfE0NJeBdi33wM6X0WwfgP
yuoeJ9wYOEdf+Z8oJIKGh2kz9T7YKqb7vhHK1JJaLi2Baze0zPcsIE6co/0VrUwl
QEKmk93p1CHaT0Jms4cndjJkZJfjv9dSzDGwaYSmaAJsojyi9MPSWkDsc5Xv5R9H
88KkZcLIvGxh69z9qbE5EAwhTxsHubk9hI0JUuIwKUdhED50g+P1KBOWs3Rv119J
XOgyW10bnRiJ/RBOE3c0cwiLh+jWE3ZElanC5yiFAdPF2S624jUQAWmCDIK1wSty
tATeA63qtXcv9U17pv1U63df+fqCw8moBwi/oyXuo2wwNzsane1AzbZ6RcI3IRMQ
XVNi2QQsv6gD8Z8uzTJTKqC2c61fICebtd9reFZgQu8pSAvxoG95xaMDpis63+v9
6veTc4bcg2n5vB5Tg0vRvzdBuPLkeS0hmTBt6hXc00C/S0v5xYSC8Dy9PolD+rlp
8eoxeKPv22WEjYckAKnxI023hgRhZS+avsV0CvEUfobqYjcIxR64RekBKcdxtAtz
YsqA2+FoouGrwGucLfSzea9cFX34gamecwYQDQ899KFFXEeZOyZlj28KdEaIwIJs
UcY74UYxiRP24pIVis8ZQSQUF1BFFE3AWvBwrUr1s05SY3KVE+NzBDTyQohtmRz1
eV6PunOd/IJTc8HfgpnuJh7e8u1scWLqeMwX02uSNIFXVMDTAbabI3pWmMoYhiQF
JnKQBqOiQPNxnYdsqLM6LkMI9DrX36PbyksPQKfjCpeokcqYmfliUdNa8QjKZ6WE
5Fa3GN56KKfzvQk1HxCXJ9kIxMgiycz4LY1LPL+CYSkVx8RMzHy5w88DI1Gh/T8Q
8hwYp2Kgk9AzkyjR27wANhfPYXS9U7iSrKzjrxJkh8EuwOFuj/icoAbxTB89UWfM
CBjDhnIUzrf8wpVzLdJuwLJpe3VihVaQkxUNIqPmWGzU3xgid/CxYtQEBTHQzqwN
GYUdJfN3b6bSWkbqwt/g48pamC/Kc3jVdOxeM47wp7teoZiBngS2ONOjKbn8KrI+
8ONzm+dwEFSdFU+QCG+4NvoeGjxqn/nMX9kFM+r4c6UdpGgTIqrrXswR2TtF4W/u
FBKaqPDcXJbh5LGDk9nz8igWHjeIp9E1BKS9IEyFdCw7cBW6UMfKMjs1zHDsJhTh
UU0gd6KoWiKzS8mqRmH1a6BlE9E8mgLub3dODjmjFuYC5UkZ06Prg1MlRi7MIxrr
d2LfmWT04FMIrWGC/y6tGwhA7auUame0vmFFJooEb0/4yVOEJHN+4CEEBWcsNJ7A
+zbGqgokNxGo4kKS+Wq0WBvGLH09nSf133f81F0IWgT7sDbdaeGKneXWJkBzSxHU
jqQvdcnpAmF9xuCHb2PYp4K0t3/bliFiNaYO5692cn4XRpNTnbtHX3svLihM8DCd
1iQiMNEOT0MZ00TJE3/0YROFdU6TbgZiOjMXJZGx6mPHNVf4tjavdpzWm1V5K8G/
uDeBYgkiqQS8+H6K57RGGf+vVG0EnQA8YP3HNhD1zFyKDjkkrhzJG7avKiYh/eig
ixZOfzaQQSC1ZQvbUbD3064zeiLwFAhq6CSkHgF1qO3LKUuUaixweSjCsoiBeE8x
GF2qSoVu2t9JwU/hFd97JzfYG91wsucFYFg0/Ht/BAo6iiTYtkaOwoyXOJBMwIjp
HCiHB1uAZbnrS03YvcBetqjRgu07IhBbBM/Dsvf3WwoXaqzrTevqGAQgQUeee/cz
YfFOi4pKouhIwFU2ljHHlgrkAmxQ2ly+FDX2HlQMytb61B+jBtgR4AYRDSRFgRUc
zOccEA8wx5tJ/hvJJauCLlzSQEvPBWP9+XVtJ9gZQDMFn103z4k2scDtscod0c1Y
loQ7bsLLRSZfWHxNZfue37WnQxc/MdXvqNd4fX90M5ap/N3xO9VUTgWzoWyW8wkb
w1+DpeLa4zI6v4zKkdD+ywQUGz/ryoMC/aKQ3pGDEN7j0AM0FVpYdBkT93T8GhVW
SVncaVqikVLBtj6vioNXh8QQARRUY+EFsH0Za7t8A44pd5U3gZ9vTZ3uKJLVDJnt
BcqPPQ6acLZPu+8p6QJSsGTLikSGnuDvmH63h37VbEzR1IItZXw+giwNuJ4DRwp0
Z75PXC7ZcTBj56xZWdTwFeLQX2d9KrTdqP/7Cienf5WQdRcYs0QVJHEzalSTpqK6
zPUYeHNTUAd2JbQBNdOTfOqiUqLzem7ICnb8MCHOL5FRyNNPjQgTDQdCOmS4IxAj
0tfaAX0ZGJZqkuIT5AejsI/bocupGpkwfGI7zpQCpKmVJLl0Ss9vvMYZwPB12qdJ
2rZpZ7LxYmx4IX6iQKO5dfyJ3AXgfdxZ5P0iUInYRrzZ2BHr5NGKAXt00rtHjkRM
zTLFYMgC8yXcqkbgoLgHtZP0swNEbbhwgj5I1JB5TLqey1a9YP0T3aamRsQ7kneT
tiBaFWBGme2ZoZHeWWZYBohxvOdxfkhYxV8zTi+t+CNkqY1MpGzKBVPgMeBrdu4y
43ddsFrvSWVnmTPNo2MzR6y8CfZjkx8Uab39QBmjQf8NmAOorJ0kx/Y8IGPqCC1i
2RU6EzVueaDTXzFyNGv7THob8BvEYaZE49aFZ00NV3bDAkITkDm12ilnDcfy6C8/
QJqVt3J9XQbYylwvjylN0fHZts7W3B4fCqOcM7rKLI2O2vrqxE21UBOz6Kepee8W
LPenmVaWIcMbu0uE4GAfWrQ8w6iKFQYjxIisCGw0BwgF0WmuDI1hCRxwMfL48Vd4
bcBU4UbqvrWndgmrgxAYjnPMMNDtevnGYsJDEdp2k9CWh8fl0nng8zh6IG6WJcvT
8/0Ob/bwI5/e0USdWVREF3m4MyQ9j9H6+u/iBOzhAxV/GpNkfQFAPFY+ismwiXsV
+9QUmeULnkw+smA/k9bebd11z+T1HGStjIgOGrWDdKtRvxKhvfaz7PinoOFVXCEw
qjkC3WVmaufm4bnNleegycfAoySGZsWp6+8gF+ejm6M3Wtjd0KAONNWCsMlqck5m
HC8fo9QztoRtT6g07Nyg9pNbkVahWBtxUI41QLEfX/z+kQDdRPHScpZ9UC/qg9Uc
Ypfc5d7QUwh+XE5vSpJE0ioXC42AJ9FqqBO6QBohEotNs4jhhm+qojVBVd/HN4lk
fLdLsgMP7PZDTzRBn1hW0TXFEHT+VQAHW9CxNlKK7YAe54RrKTVwi1D3NiBMfdRI
YQdHwD/KwfXqYAmJa+J70hx8Fz82djkjVm8VtTjnu/H21+9QyWlfnFu6eIG7OG7I
cnA1tCXR88zPOvIyiGUh+9CR74O74RPudMaJpziuiSrE8f8yLXHdg1Z1VIRTvuvC
WEypu3h1Mg5PllStaokAHWaROboTre/n6Qkh2DOcIm/0sLavNbmdpTHYtVCwTueN
AWBL/ugKU1Uw/+3qbD7UfulPo0PV/FK2jEd+wyfXNEcCWEX/SiOQdZY1f9euV5nl
xt7Gue7sdAinlEQeDnQkCSfmN7ys1NNyj1Gnd8H17aN3SojQXBWiD6s9AOlVV+F5
NzDOduA1wLRxxcqcMTIvSj3ZLfqhy5b0NJoj99+X2NN6JZzclhGbufXqJmlxmGIA
SQ+zSD9BpkZed+1QyEEgTY0hIEXVyZmix+oOnZGgHpuevGwugzvPaQn2y7FB12b4
ztfs+2flBykjDei3aqaissNIcVNJPVGt7KU/H+cDfbCCuDXiaPnNpzdz6gVYnP59
dv/uv3oAf299dH3WcvuOUrg+bFfgsI/wGEYIJWsLRqok+lMz1L3l0a+HrBbScIZV
ZhDDRZzptQnLxI8w+9nQFG0ya7n6mbeZZBWsvRFKNFMAG/Riw4JnAbY29BCMl1MV
qKIJzpvkSLfFi0DB470al7hsC/U226ytUIFW7hnw9CR0NWOejMr1pac9dyKEvFZS
irwChNDkpI2ThUASod9Z9F9ZhmTXrAKCuYscOty/3fGw7o/Rm/vbL0oDH3RJYWgS
bbN6/pskuYCXXo7m2z7gugbmV9K23gaOMcDkBvL06um2+T0Jby5gBmy7PeRMekw4
HwZQtgXuVaRI6EJHvYnSnA/ifWhnrUENVgojbOt7Zjw4qZWeIZ0Jm+dNQakXaPhM
lBmiwgdrAsbOmmGM5N8d+OmvGvvAPMjJfdAH6lscy2GL+59mrOwOEo/aulkIqRM+
BW13hTMPby9ND38xpX19wLE6f5vLDRD3Najqemjrq8rff+e0E26Vi5gl6DBJRe7p
XmmEUawGYmMefJeSRofL4j6LB0Vldi2cW4HE+07k15jNyS/dhkGqueBrfo1jyJs4
S7/+jOWOyogdml+Ant40/SpmkwNy0BPW5ELwI6QUtjsn9WAQg4KqrlLNjuIS7zCr
xcJsBw5T+CO2PxobT8DvUW3agz/aP5M907MeJHz58aIhERCZKMg+kbD8w2HbmzLb
Subl0kBb6CS7H5lpgM3SDTkeNT7Ri/q400S4EutqmCf2CZOPUtNJa0WMlBU9JlGJ
kfmS1NwKFxU9yIkzF02RaO6Tswz818IuZ/xQ3CA15OtBsAuQpHbrQNBomrh7WcCp
0tZeF+20mWVLbRiqtyDmCieOjVcmfzmeD9uPfpbR8Uwu3yMVha5Juyra+tyi9OJi
1pEYSYoSAfqIHj+LWgyp28pphb2Ii/zZMA0UVZ0FJpmNN8Ih2W+/EaVQJP2u3A0E
doDUPDKIzwfa5qO8B2ofhLHyVikBxwex/eOhhHcj/6MACpsHqrLWq1/y7ZDQhmyH
IiNq7sDkA4pjTqrL/QFh3Jp6MZ0Q+EwxgMDq09ZLFOHxKXPayOVfU/yHLHwRw4VV
+BPPUgNFnwEebhQC+XRm4UdFMi0pChpHwLYbT7O7VNm3+Yr7qv13+LPcKXMlRwJF
BEiJyMRzVqFXhwYg80/OyFnSmGmVLDlneIwIXl5S83I0hMpkoJXJ+hovZVqXGgMB
3QC75kjY5i33QX8dxKPyS8UJhcRQhI3r3XfkYcgyZV7JkuHTG8NnoqeHHZI+KSqi
G1FOSznSeW9vlMNqzSHJTSSdQdBebppHbpZVsV5bBwaLp3gFSB+j8r7vA2D9erXb
luF/2DrcwXUTmv9mej9R2u4ZcK4GV24c84NZbJradHbMR7Xrt/U1zBDqlE4WirDr
jR/oSsTnxkOIram1YrL3kuIXiRsKIcXDCHDcTn5/fxPopeY3f3AeG6r2JB2pzf3P
nST20LSePSQUtFKawcmw4noAfEiq8X9/mpuSktJB4RGaPpjLbdUA0oBt8Rbv1mPf
8NxaTGqh4RN/QzCeNyQeTnfga3N+WdG0NY5R2vHem/uDSng4R1gFjSL5t80DZXO7
IyS9QIXs9GW9Lfr3ojizaOfwFf/Nv2iYSheOzmASQouu7aVIvIsiqw0qVqD3krmW
/mvyQiW2GarGlHrRSzX/wMrwEzBH0GBZ9pqe0zzKgkR4OcYUXBSlZEQI1gRZogV6
/yRFwcvHWg827MCNpy2V9b40CypUhPyC3fOYMJFBOwTax6LfxTQcbgy7A8saZOlr
OCxN9Q0I5DEa9Q2ow9qLQgPBrwCvVXLSvbjrzzYyhUVeqd+93BpQurF3lHBjoxM9
/MdnynJ+V/cF4CHabeQy5hw1/7BsYgosMcq490gfMhKGfdabKZ8WCzeRd7b1MGkt
68LJYZ1cdQmdFokYO2mw9RyZcvLq9OLwcGYb96rOtn5eyh+zIpgq7QgBz7ZVdUrx
uvUJdKNlGwTdqOAdRjtqWJNHUoniMFOD2R5SUGCqZ3sKQqkVly+qu1k2lGM6wpR5
heKHveD71ykedP+kk8PqRSasbAe7oc6uksG+LSVVtzg4+WvrtRBiyXc5tqswAc3e
yF44eGuaktu1e4YpX2YTvtpUN3l4rvY7zQ9HkPFwuQq/o8ISR4k4SIXCOdtcifcC
o5MvYaWz/qYGlQ78L6Z5pK43D/mXgmakGk9Po8Mq3sTJbtPmWZw2pmhsg7BXRK1g
BbS69WCPgm6cwcKbMtuJOpASJ/AP7cq4Xn8jo2M8PU7pm1MEGqRu2mxU5U3x8znM
87cyvjJoBDnMrCRZD4pZ+cYsQLS2+vcgzeTBx/jPvTj7C3kP7jS/FDC1yL/eIYeY
vdGc9NqcQrL+lYQQUI1xMlyzMMBj1v9H+ZOZoeN1s76vVoDpUBsy/mAUe6KHISIO
VH0xvqomKiuS2jHoeVKxcGqNCCxqY6cSqu6LtXst5isDFuAvOIdFlDs+rUHitQA8
uV8Nyt4m51IyMiICu3+I7fTOjPruV7tz8VNvf5qR950TZ284GMifJJxfm35+lN35
KAGQ9W79JFsdazhjjd+GBfRKIw9qDmelV4yv1m3QvJoUPhwM0yfmVRElcC7jc4A8
HQnLP8v5abm7Hk18V4+xTt4dlAMSH+Pj9lytoZY9opSzjt+fW6RYvSxkHtI9de+T
hkVj00gcXUudHEmvMlGxtfu5vont3LCwC99rqdZAcXLX8ctl2NEl/le3Qn+QOD2X
6pAGMkpGfnfjM+aCa0SOfqzePMpQpB1nwEmJpzGI8b8mXEP42vZDwjLTle5F0HBi
gSnkFx3nQZ2JnAyf9E98cj7xQfztQ3hK8O0gD7hz0p4svx9lJlrVaJtSnCRMld0g
uEUxnB6qFsEdGDPBKDJAalftNPyAE6zBd9R8YZo1iLPpxQHWUAG21BY1a5zflb9e
dcXkOyNfg1NedGT1Kal7OSj2TMTHLF4JswJ86a9Of3Aws89cF6u9BRP9yYQykJef
dLBNm42YfLY7eW2baDpK/zPWc+cfnkedoh+LGIFEvw99Uu7E+mUwVuxNmgtFXdJL
zhmfRHfKtJHs47Qp0bLVHe/i6R55YPH2g1oV5iPOQPFjs8XW9HSKF0O3ZfFssx7+
VeWzKMceLWITxttTZPx8oSBSEXAIsSZ+piTOxQB/cCzj0PvGT0O/sIWM6J6O5fuw
Pu+87T5QkV/vB8Upfx7b6nS1rgAHmVK7Q4agL25e3x+3MdR/7gVx3QDKBdtwFWwh
adT7hd3yqzjqxpf7VAjSSpaPJUapfvQHxttzqUwpDFRwDzH9b9L5BxkUgDGASXsf
clTDnav3d2Z5UGYQDnWHyLgz/qhFVkkJV8kbjMYfo8T+DaJ/dN1LW4EZqQHZkMGx
a0KIWna+HP0mjNEhpg9hnZFZ4w3eUg1wASNF7QxLL9ucbH1Pro64b9ZeulOdtshZ
6nZV2Y7wl0ucATLIRdJ3h/9LZfsWmvpPNq/0FaCBH3JwxRWgWrVWNxxZy6Z3GcMr
3Jf7XF9Q89Sh1jNoYLfZvmfa1Mw8vqvOgb4JnNtbxcDikbTkoTB2xX9mkvKcaK0F
nJkEU7FD8H69KBsBoIjLc+ZmxmZjSITaJnPBAyV/GK8CrrkIhcrCvoa7YpZE3Y6m
GfxGbwplo1cZoz4Ts9DYWQBlTTmMXKUxnhFMr1FDPsNiFUP4b6So6DIHiAYSYqcz
bWBDJCAHy4ujxDj4H49BKQypKrzBL7ORDLxNRjpb1E3ipr/alMTZlzj3TSv1AzLo
xAK6dIMQOU4mhjdAZyfBg8gaYRzfYVaP2Yet26sgqjxaHJ1YE/L2NTLY8Gp2KTwO
PocTxeVGIEPakG5fuYcle69vMuykG40wLQCixZ8lMJbdXMCJKkbwGEK5ghPeacNv
XCsvwVXzDHtyBKU8rx1xSs578w16K/Yk21THwUasFOUHza8diSZ9bfIikFlUJ6tj
FUSYHX/EUpcMj6CCX7Ub/zJ5ptph0YzTRZSEan4Q6Zo8qTWykSruRzHwwQe0SUio
3AajK5JCrtUcsb8yaYZkwnt3rj3cLfvErpSHIQ05HWWOn73UN+4fxPK+oyCqV+SX
TEsM75+H/QNEbyVnffDVCZJmLsfh41zgsEx0LeN0CqJ1hfd3/PjF/FRuz1VrMDFU
1B6dZ+S9uNYwLVZ4CkZ2Gt6Zjdq4Avq95wP+a8stBrPIukPqj3iPcjp3axoC1kbr
jot77UyuFKh97agRL/G9UYdkISOVCmKaaMmw7E2imkE0hqzw2aI+XODIyvElzl6w
dxMYUuKsChsB9DtriVI/0Gf+zYC+w5bokGAb0yf+tpB87gBsm6N4JthVn/gcsj1B
cTZYjKDmTMoLc7WWSVosjzdtpG+RQap53RWgaQpLeg5q6zlbexXDA4xdWLiyq/tx
kmFLGqalEz6p6mKVX99TFYVjPMd3cLcgKcuyphasGAFrKuelalwzrfAuOuPJ8fNO
DE+6I2V/wpDkDFfXJaanpoeTVhL3jQs9s9uI5jdKIc7e+sKkYALWnfKR+6QHtmT2
hNH/39pAoKCVG7jR5Qkt3OpMgc85B0WpfkhQhBb1mWUtDR/sDCQRIiF+vG8fkbtm
gIyFkBKZ9kwku0ZxfRT+Mo6hKRlKn/3ZMURxM+V88zTR3f7HGvsKxW1tZPfredST
EDSTXIuXvaNivtz2Rpw/7hlGzrMDmDYGa3u5M1WmI+hPZWkbfTiPR5/F+cFcyF7I
ndiCsU8XTZQd9fmeyndqiJIVinf7B6FNqp2eE4+KdNWIIjuFV9TmMy6Pjk5qdB0A
TvnEuldQlGi81xJP6cnEIypwuxs5rsbasn1SiJa6lRhvGbnisfjaX00ijBYFUc23
MNU9v7Peoh/B+tlSoPInPrdwbG0vyEyoByg333TTM0H2zZ2EySmdz421pNwQV2Jh
VQ9/PmnQRLgirriqlnRrhxSGG+vWFxsCMXDpl9WRtJbdr93p/IP8gftvyoD4dRJa
uBUdKvIijQp/VkCr+8kFqkXRNju77KdAfmjaU/Kw8Lbrr9d2sFM7UL0wKXnqcuWR
/UKoG2ZMduQNzt+cRcn6Ca3fOBfn6KPpgzwK3VRySyqHauoYt6SxBUUOeImRa+H1
I/q6VS6/yHvsAQMPOWPkoozYZF2Raghl47ugcP0u3JTYDMfoMrX2btSrQaYGZjlH
ypAU+R7kzbuTCSSzdIBG7pY43S8mlACEdB3KDY2pFQ+smGNkrCgxtLUPwfT2N/GH
weI5fPP2MJOBmalQY1LcfoH6+1gOGedgzAvO2lWgujTchw4WoY6xo/Gcquvil/e7
ovBR598jDaVoK3gCsiqKHGAlG+dyy25gocpcqxXpiCbzB/qAjEWMJN9IQqldwtHT
VaSY7GCXFEFdF2kKEhWkDERwb5GWeqFz37pLCg+q+QT7TvowDw1ZDo3dQlfWovOj
27Qwi9o6kRg+xprxABHqyvfYQOY4mQXyQbU/RheKg6XhjV1YAGYbGdlj8h9SJ9/Y
H5sNgzJeFJhiR4B+VBerS5trjS2/7w/tIRoCuDLLHFiy94poA86rJvMSflt1T1el
xEF5i635Iu81wp7OGx6wic0WkxTVX75Wk+RE8vVgzUIX0YTgzI/5lnHlxpXrrjPQ
ugHDk5mKK2duS9dWOt8b/k5kf9K/JjGGdz3ocJmcpI8fS6JZ9tZLE4kxfPbNchu7
41LtBptP85ixeN3DLihIjafCo3pERUgEu7VDU/LgIQI/V3TWdiZInMP43G9rSJyc
zNtCEKGr+O1g5CP+rsMLzwysayf+BXvQQnIV2ZpNx3+eC5LQPFp8aHCicnqIQ8nG
y19N2LmrXvSq4HAjppvzb/A5k+UufY2gdqT3s4sQsROrKyhcg5s8TcsJ3aZO0JM2
B2ZTo7nnTjsjx8zbqMb8BkwZbLiZyHEPfItNLLGVkFIrUyaNjQCey7VBtADUrPZB
L8vPsmr7WX/6/mHg+D3Tg/jGJsoHNJuJxMQsCQh7JnQPsnn92XZkaIwzwH1XuAod
gyp6O0nG5Bmi04FltOewMsJb9n96KsXBmXl7yFzlM+BUvqoHcQ3x0PY3DaZgNYz2
m+e4ABsVyx/AL/Tj5BbsfD1TsexaMhL5nCW5qFzIlPhLMSfXIBjJBh0wnwSxjlDs
ls8ogEtFnXLtnXkWAkj9ATzadVxqKeGp/HGq9Yb/U3c39P4QXQxBF2nlKncmBrZN
+B8Svtwnz6hAD3Dt2yN1i8XJ/pKSlhPcOlGoUbHB5djjgD4zrX73dUxosCcxhhMR
xmNrKq1DtvUv8sbGiQySGON54l/sxO1QFni5L6W2I/w6CtK0NkFtsfki7n7xLBmQ
2x5Zk9jrpZpUuf7d4FwupkT17YSbAL7Sx9+oxCgeV9i2JFxkZPb5eW8SCT5Ag91j
e3K609XsTEbiTFc4Z4nxEtqJWMImDJ3xC53mLA8I08+Oecob7N5B+Oj3HaJ4NUGU
TUI14R0TZnu1ZLeokZBjmO9xBtpJ9yjiwkZ28jAfUBd5OjcBlW717q0pxo46N9y1
ZIHwFPMRFP4AfgMGBCBE9a5qxj4Kf+ZuzZa4AFiJKM0x/SaesP3HK2v/OoY0H7Nd
mWYGfGqxjnnkLoQpKHp9iyKMaOh6O604ZcjPWPPugMtV/KwcJGkPfmAAW+vDH1Z7
99+Kcq7KExSU96+xIZb+Tdfmt0I1qtr5WK06Kyvo5baMJEBZgjWjxUWnYJIdgN4B
L2n7KYPO6ejlcuyF2IYZ9gWY5Mnu+Ix7p3pxBCIxDohEPZimJczZzkmPMR9vwn5m
7iM3wjkHUzsb4xyVaVCEncItl/d6ZKw6AMFsclCLx2qYYguVymiIQKBmTuc5BJVs
ylA58mCajQ9YWglOfxFgz6gwN+Q/QFBY11GcMqKqi708EpylsPYWWUIH1lnKDtbK
w6Vq6ILKDhfOTrCH9duw3qWhniX904+32Bj1u64k3Fdm5u2h2SNbNrInkYMhLoHf
TQU3b5XTZHQM+XqCbhycMwiIIhIAHDSspAV3oIc8CcwT62j8sdEXosev7z2+OAsh
sdTjMqSrnIr/ii9IMSSPq279JEpQCsHLPJ5xGfXWT9VjGxEi7MkvFbss7LLHcHJp
fPLPYLg+N8hOB2e0GEBAoy1xWu7CxhJNlJompwGmPt8XPl8xwuTu1QhUhBHBRwur
AUltTnjNDv1JCSrYtBBp0IIupFNuHbMbRBWGIq3QCvzWaspEr0jBVGpbkrS9OCKl
W/p/LE0KcupXBVPzWq6FAxO1sKkUv+nXPSRLLQ4njI8c4QIxpNsMh9+7iomOqTP7
Oi/bjRmMmVhJmUtrqC4SU4S+eglvcoX9ARZ/YOVBNp8lqtjkwj3TgQvPA534OXfR
EB2CvPSCBLlQ/SXS7BQ7EBVxxPD9y/wBhZBqEQiut2g0vvzHKPkQndtHBEYYmLT1
Rss4f9ivd0x0R3oMaVBNy+mMeOtUpvJdpsY1TWOdeSDikYJSq5YUkqdd5j0VSpfp
uLj+SV3U7nwGDWS01pz3p2m87xOeq+eGNuxOGlaQTalFjy6aEmMV40e26iU2IMKJ
FMrk+e61+vXJFrs/sx64VqpIIg98Nkf/SiAtEhx+7zXruOtENWfXUJZtsO83eIw4
Vw2b8Q/4XwUu7GGT4itI948DPYDGovqbifZs4pSuT33NfTd5AmkZCDdbLGF0TaK3
6OpnxuohGZCVYlUWIpuCTvQwXTwbsD25afPifLmLIriO37tYrC+X2k7EQY4n9suJ
Vkdr23ZxgjJ5Zw7L+d7sYj0NRMYdCMU15U9t+zkCbtUVlAtbqs4FyYvYqLivhpHR
YnzwnlHfGhdlmK+MIAnIy4FlC225LsdIbNG81H6eRqU2HM76qJjOCrXZloCxuTWK
fVviicB2RMkOZes/0AercEBbSmOz5JEMw8I4g1l10zKQtAjFMMw2hhhEndm01Bci
9BX6Xh7bJmGFD/LTfKbGuwBop1hPn5FX/ZMbut9yOuW2N3V5yCD/UERVuxlW3SQM
rikYa258HTmp2OjPDPMsJqs3wdmnicAhxZB3/GGqaW7jT7AQAK1LY8iz2kYSsJyk
MtbIjaeEsUXdrEyOCdxWVAUSb6qRX987lhFLogDtuq0oh8emyMxRnSitWIrrkcZG
LuyiY3ihCq6rkIQJEYIE5tObgWwU0ESFBGQqLX3nrL99AibCvBrgYzokZbuuA9xM
1s+Vg64Hjp8PRmQceKud/Ub6WCMaOqTAUP8ILx5sqVQHnNBQUoRHpoX7fkV6A3Lo
mRttG6qv00cj5bDHSaWwQouhDMFOWRu/Rws1ZMBgGvUbEoF0ziqUWfy+ea5rLPHZ
OFgOEVm/tN5MaTCc+PfW3dQtM1laevCPE0Z4KZ2gQ17YfnR45lGBy0WoihuzuRMM
BNtBk4WkWLrPScP7r32gJkwYjGmgMTK7jL1d1HXouIlcpyulW1rocvkm+YAOAE6T
oF/aYEv6dM+RiWQ33jEhGqzxKSTf4V+mS4phnmhfwAU/yiYl1rPrRia18fIWX6Vm
alIGOaQhnfNslINmhFLnNeRbyANnhoSt5CHhf3TzNDIWUmWdSoS0YqnnAKaCKjfa
`pragma protect end_protected
