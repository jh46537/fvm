// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aR/5yBaEZRvNgekQkjiudC3HJEoUDOfzinEhbzK/QoGBfpiZlcic0OAP7bSv6S7Z
K903Fb7wd1fD8eErF4eXWPkSkcyq7MBFI7BzFZZVeGkiXaqXlq4/MKIQKpgbMxTi
lnc7EbHv42CPrqQSwWdBGGojReT+VvSPJ4KH3XVyupI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2704)
wuOA60ShmjIQdXZ/i+BLEMPoWog/uO8wtUhCd9CmXP8Yhg8HcgDg0GjYASwBwrIq
DXtqWGIbNQk/C48t6axOVUZABjyjWkFgz1gixYAKzRpSyuaygpbHbjU2GfRbEjAU
c77oPub318qBefrRlT15LTr75+oKxjXZ9SzmAozv/CIPqmqnZqEAAe7E5Ek+NS64
UKQzYeYFOYgrhGrOyZYpp6XUC13sO91VyAgKOYSdSg+KbSd5ITwEWo1fc0H3ju3j
I3ZMPHz7kW1eAQPdj25R/B5CRcUeCkbfKJd7S5YYEmylRkNAu9qGVUakaxvaXPIt
SefiL9pK881h8I/3vrf6r3AEH5bhOE2aMWQ4K7B4AD3NJOdDu1bVtGQcbvsSVAlY
PS2jAuqJiRTsmJgMe6Uh/iGtsEcINvz4rph+KZKSMAmy6mFGf6/ofhnuCDkmeAWr
ieZex5KwRELA7mrgBhFiwIFjr6MZY+CUdZs2MJ5ZWtnxOzpg5/ZV8rQgTWZb9nVN
2/KHUDW+ScJsDYsYyKOUYl9RGTS8nLLhenjfjgwlB8/C8clr58yxX9LhBX0cFIWF
TV8gSwAazLZhX5NK4b6+msJ/OQhx4bXFNja/dRUE0/T8b4reeFB9E9DEC1UYseAt
D0XLHlxFmzmWXQ+cFW0hzIP9OoW9OSvMU2dn3nPbqE9euGsSwM6UCAhkTATuSNfZ
yvgKYkulCSykKtyO8kSjOgKHIoOcAxCGSUeZ1YSG6yt0ANUW6u/f9ETf7aYXTj4G
AyUCwzElHIf24qdfXkF3yO1Os9FOpaV1SXYieU7BroHC9Nc7erCUSgTdpZ/v/jhx
lgu7+CnyUaTZPEhMeVFWu2GyqSgsC9J0QxP3tRNa3GeznQ+6HjfuiMq0uqC1Ds4K
HiKNtDtVBtr25LeUSD5UAcy2rqxYK03sTom8ifVR13V6M1ycqXdFE7fe0/0m/7xO
hvgYogkYKvXcwZAhSc7kmJQwg3hfqDYvpEpGysA7RylIqb2YEwT6dJWN9YIR0cxw
SpsJZTLgJQH5MmvVomrSnJOEnDEemI9xDnVGj9A0l5jkxTzkrBersIRBXX9HT57r
tATr7jBvBaV7sorIsdn7Z1x/JUgv2kAmbNQ89Su9KM78OVA+0wnwNIT1CY/7PjaN
Qf+KpqML/QEjX7/Qe0DMkRW9862HaUvnbyv96aHPN6fw9kgGfHeIhTMmOz1ahRm/
mEWRoZiwmuOymJTJm/EGTpzxuozT4p71we2fKNwQVTKNy0kH7WbBET4pOIdbQT96
KyHOWEthYa5EbtoCBG8EVc+fEWBkcPu22PVCn9EcCU7oNQ6w5XR2cuuNWxb4tIuY
wCN74ws8MXIZSfT2HHUo9ygvpOmtjKw4MOpcESQkDkOwaQU9S13RSIwWEAVfyUgr
94pDlyu4pBZigiwErBUvIhEDAmEMcVhzfdIH40WV7E930eQPrla9kwKGC9gES4EI
yMrr14Jx3h+FoSMc6IfC6abPXbmh+1gNWTc9oUFkz6wFf33WKqiA1GrbKLfcK+Mo
DOniXppdcBQuTr6TCFJtDOSMOcScoQhZ+PSd4JX5KFZpoioXlwf20WupVkKJDVEO
eyoqPwy3g4xtpjPOz8OQA+frNjuwL6v++2Jwie882dwkbpNivVOFsQLWzH8hTjmV
6lySjyHfU1K8nMIXBnBRHdYm8CrcC5RaAz9Tq1cZ/7fW2EfTK+qPWmM1nGy6W6KF
GCQPWlWjjW9Wzlhax6rsko8W6lxOyjsMsEgStAA8hpm7kvOxZq1Fm9BkjZ98xTk7
0wClrZHGUFc26PGlqiKcI8U6W5Kgk85ioYzmAJ4NLv/a1Qw+tYM7FYXQihKVeraj
fwmS4PRiZL4yD4sAr6Pge6/lmJ4fSs4GSkNj9wEtR9KGWoIr4AVrIFNToMWnQ6mu
3OSoM7tOqkiXHmcbkqhfAT2kwbeWgOhYu7mLRBpHp+dUxF2ImeB0RLSvNdTFac4u
NYmx7cdJCQmvf2luFaqg6lRfP10DD61p9Bdir1Ecp78x87sWuMGEDncjSD9nSLV7
nTL6Oj515kldxtfwZ+2M1p95pW0aAm8ndMRHAIiFJzJmiI5Av/ihAbb0Qju9nSwo
G6O/05EFxRQloj7ObtE9Z+P3Z24/z5vzhXy8ke+YLybcEG27uc3Th8wPT/VNVinG
pYyiKDS6UwaHK0Oi+libHL2Aeuk/5qwOXAx/S8Q/V7aS8DpcFGvtoB99CD77cp9u
4FcURfHl5/Ss9j6N+oZVm1mrtpF8eFbIg7O9JrsLpQiG2KYt+gM90CCzOhK4uZUh
SjfXf2GeSjxUhTSxxM+34UD5MVx1pr3Zff+u/WyfoyK0Io5E4dgwS7fkAlzDW87u
daRoVG9LQydzzjH6sHl/v3w9IJOdoQbe0P2mZl+ogF6nbaGzRYyq8ins/nm+ABWw
2wAIpZ6K4G/WC+xHrr+RQxatpZEPsDhsJ6YWA50VtxJeUgtCTyfNun3HBq7bVVKc
y0Wa0+P08suhKhNwQhqkpG99Hw6ng0fqUUnLV5fl5/lx9Yr16BKtjUGT4gyYSMxw
xeIuP17H6R1ZwOhu27ST2miraG4BcDY+kP+hLi9J9zwW1/ia/RVMidk6V3wtPOWz
eNBH2REhqNno5gKk9YhLXHP0dJkItkeRQJYz0ZHokMPpXw4CcnPvK3sfyzXNDxmc
xUgb6e2JTslveh4pV0laZH2JrU7WUGNZUdkz1BjXnuAR0L2PhPA+3U3jH1eekzh7
4EYfgxyMXFqvxLcgOaTLWzxInw7ENBi7EfjdaSqU4F4HNElsXHgKlzRsIz19Kc3a
bLBRPmlG/4d99HODE8Nt36MIH0IxY/sioal1/u63Zvn67TH9FeqbEse8MRxygst4
HjlbLCOyHJjZ4wr6Mj/gECH10U6MK8ieSQdXTjESS1jgoSrX4DW2eADCuNy+ZFYU
BKCsQjd0aVEAxim+V86nrpmcnczWU99oTR/mexVvx8U4/LXX3L1aH5QYX5lJGOfK
4XatPu2lUVW58e49x3FOaxnEO1PrsqCWvmD/iD7pY2ngCpy2zUbaTfAlR63p5zJ0
x8yy+ktpVaKNdYYU0DCrYaYkBp302RYh9bjvWaaQmWmRf7/7D9rJS7ETjxzHdZd9
Nt0GNzve3DgMyywDTJYLsPhtb2tZ/3geiuq5j0vBC3rqYstLDjSujYrM9CZyFzJ9
19aYuZYnUCKvqQMEWdGRxWjWCSUpxyDQ9X3NbAKc4aFvxBnsbaDG9f1o0CRgr1lD
tVZuhojtCptdoJLp/OVX2duvs/RnHPHw24STP/CS5cKf/n2Y+zJ1Rw6pTjNO5lYU
VqewnINYaaFUa4izs7yJwUra9ZTXKnzDjNlfoX26679x6dikdXR/qnHf10EX/Kqa
oGW3Kk4/tcXeG+XpxgRhZ7fZxyNNWgrBDhg9A94Hs3WKqcH9W3ch3ykS28cHQI4t
OovK04V92pFhAE5qifRhnhldTsiNoz5Az5CFCUSNzgGvJ51JuKR3mjuUq9S4BIOn
27EyOe8eLzI7MARlYMaZVmgCHxRx2L4vt/EIEyaw2Jxp+mChBAvMGvDNvIaXCFo4
bgl2mbbutU8vGGif7C+e2w==
`pragma protect end_protected
