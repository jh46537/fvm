��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħP	�(<�%5,i v1`��Z��7#��kϟ�,�����:���mΎ�n���T�-d2J���C��^��3שl7�7JX�'����z�Fg০GA�"O���}u����P��	��!O
��u�Es�#��`Ն��l�,�w�6A��M�k6Վ�dl&*lw81f8R���T���'������
��u����=�i�ާ�������G�w�Z�������=��j��h���4M��_�8��y�fn��t�(`��ǣ���p*����OK��v{j���a�j^�U�$�*���J���d�� TM����IW0+ �����%F�0���P�uE�����B/������8�^������^!�B��Zb�9��p?z'���-�2nHv�6����A�R��_��'>s�p������8t�c��SpG�iB��<��6���Q�X1��P��8 �7f�e��ˇ��@Z�~XD�ecNw+"��4�3��3�O=�j�e�9�>��1�-�[�7�R�f�짾�ELӞ�z�Aa����}�gJ�F"����{#F��#���r�X���͍�E��}�~+u~#+<�nPN�� 7���_@������!�pa��Q�H0�1�	�o����K�!D#���d��*6Qu*ZQ�f:�����n~��3�Z���4WA��\ϯ�0��� \�jPf��֘l�l�4SW| x��H�����s;�
\v���7N�Y��)g{g�gL#�&0̱&���q�!�)�"W����6�h$��E�r��X�N�(+-�8�ϲ���1�@�7��*����ۘ>"O9NϠ^XP�z��/峣�[h�� T�ꕵ�O_�=�?*u�Rvs�3C�l�V}BY]�-�Z`�v;�
���~��_����R�ъ��p-;$��>���"�'�[-��!�R���:��*}#fR�} sw��}}�q�3��W��q�m�[G�N����ߚ��p&������N�j�u�����J�K1���G"z��Ѭ$�W����N���7Y���FR��2�8_<�:��� ������f�L��q<�P �>�w��*eZS&���me+��F�^��Z5�qI0��N�T��;�p]䫭��h���;�W2���N6�`�bg���y��ʒ���֖�4��!!���,u<�V�L#]�w��-k�$��<>�y ��zv h���!YN%���0�!�{������Z�{ƪ�kGU]L�A��+��ݰ"
�~�ʳ�)h~��Ͱ�y=�OS\�b���(M|��)�*��3��S�ߌ]��;F� �B?Ek��Er0do�Gb��)�,�eK�h�cE�A��c�ۖS��G���9	+n�jFwăF��N\l9�)�R��{16џ#�p�oC��H�/Q��f���?��ļ�KӸ<gd�4�l(M������
P���������N�n��8�s}w3�6CAw�l�>^B5?�Ƨ����`CG�U_
�&��RQ���ϛ��0@��pV�#�]Ԧ�v۲�JiaÖb+
l�Cݎ��I3n(��ES+L�^�צ�mN^<���)���N�"ױ�2�Wy�2��ֽ~mQ9|Rؗ�%����B8�9nD�i�~	k���}Y�z�J�bq]m���\˻7�­