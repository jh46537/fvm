��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{T#�5~O%�0���tko�^P�R��h�8���ƕ�� �� �T�a\�,���E��3r��=;s�;63hzQs�͋�u_�6�5���k���͉�sl�n:���c ?L�F�fR����/�H�C��LgY�Yq��y��2��9��O�鿕���@9�t���= ";�ϼ$������h�/A���j����Gp��� ;�@˘2Qĉ���I�X�$
1����|��1+\�]��q�J�ZbWM������/�ܲ������\@%A������U��5�KE��1=�*��~I{� �t{"��.�M��U%Lf���D%>��9�t�%j���#�{l�%�`'��䖝�`<�;ja�k�6?����:~�q�媧(�	�6b���{B�m�y�$@|�W9um�즏0�@Gn�r�y�W	C;���
�nD�Ar�}�
���kpl3����Sa߱,�"�������5�d��Y���U n^�si�U����pt��	�_��6l��ɤ�u������ã ���w�Mݠ�c��/ſ�2�v[���S���8���off��-�ǵXH4���C(����A��)g��A�,���x������R��Q�+�}Ѡ�D�le�ɖj��R#��H�ޞ>A<��W��t��G��ȳNS���I���
ؼ���4}�/�LX�	�7���^`8������+�p�/,/3K��'T��g�����|i	�qAq���s&�XO:�[�+�q�?�NI?��
]��@��~7b>�%ٕr+(h�7�b����HF�XQ����^g�ϣqeJ�?�/���w�˘S�pE";�<��\rN�l�����<Vm�̺�,gĬ\��@o
��~�pg�b+�
�״V�L� ����c+�O�#�g��F��]��*E�OZ��C�u�쉏���e7�k���d;�
��S%gd���,��D��Ku�2��NeJ���xs����WT�Hr���~:�2��aZ��oVC��ɏ8�/jl�ۤJ��7;GG�ܥ�Vo�M����<�Z�r�>x�<Nn$��lv��NDG0�����z�R��� "��Y�J��� :�ro�,��`��"�Zr����
���J_�N���k%��Q��1GϝA�`��I��2��%`�Q<:�����-�[��E�ۣ-�b��'���'�FYAӸȾ����JN�����\ඁ]�kׇ�ϋg���8m�ǒ��O����`�x`���Bk���P�1A�����X��@+�W�E�
͍��VN��3b�_�t���)�9!D�Ki���t��RlM��R�*��7rZa0!=WT-m2H���<��[]$��2%��x��^�}��XY�_?O&�
��G�ϣ-b��j������z8Y�"SpE`�V2$��A�|��e�8�SY�ގ���d7sqj��?�Xb�E���po����Vb>p��� Rb�#�y�7�� ���� �X\Bu��э��.�cLnjn`G�� a�9���{�d2�oRT�\��J��R�!�T�ʠ���~xH�-Y'�8��;ޏWQ<����f��EvtCHQuї8���u�s�\M�����Ɇ6��'����|MT�X[lT�C�X�"�=Cmz�y?0>�@��4n��{=��K�s���)��*o-���� P���6��	&�pzYᮥ*ԍM��G�R��SA����AK*_Y-�>/~�G�d�藺{�_�[&[*�A��='\�W���87B+K
���~n��ے�VN�h"�I��|ڎ� �U�؋`������`�LI����m�W���)'����&�q����� �)^*f�`w���ks�GFHO�X�S/]���X�2
�E�ԮD��4�
�Z̉�X�M{g���]E��������tQؕ�q����ŋ"��w�L�RK�e�ou�L~���Uj�8�%��}��p���U?x)bʠ�KpΨ�GwA��j�	���A�(+��ka�U_��ޟ��^ۚ�2]��/��w4^*Y���F.xo\U�b�A��d�k��c~��a�ol.K�;�9���ιd�5E��WW*�z�+�����mQ[���R�,���b��hS��i?F���a�`��J�!Bv$���n��g�e�b�����s�vj��� É�0�Eѩ��^�2���A�V�A�v���l~$��ɋ�74��a�U._�}�x�yۉ5Y��B�J��n�<J�=��k������xg]A�w0t����9���MŦo�!bT/��9R<����,�dM�V8���VL���:zB�=�E���^qoú盠��t@A�A�|�8���n�o�٬*���+����Ö]0����d?┪��2�j0HxVgf"��e��?��G�sG�+Bu�4�<��؛��H�%�~`��q-M_�ӷ��-	��x�ٓ��[|^�Ƭ�2��ݷQn�b�	}���+`��F`Ϝ�~8�j�w�u�<́Z!�Ewy��؋4~��%,���40��}*c��v)��©o������SʖD�]Ug`ڧm5���\%�j��qQ��o��ְ��5��FKW���9V����eL>�6�,N��U0'FJD�����繃�Ʃؖ��@4[������\��(�ҳ��D)�`��������A�`�(�MP��?i9��]zDcIf3��:��a��u�$}�#4+�"E%�y�;ݥ�p!b��O	���`n&FW�/��},��f������%�"��.u�=cs懻o{��96�{�wD5�>A���.3"��g�Vs�)hU�#�A�9P�H2D�#��ܬTO���S�j{�Y����>���8v��_cd�q��D����ړ-�*\�Ǟ;h�� d���+�ڪ�W�B8JZ����u@����4��n9��c�h1��3J����H���ίG�~(�
b�o]9I�m�`:F�]�8R��^_��8���P�C)g�Ɯ�N�ӿn��/��e`=l	�� ߑE���8V�d�Jp��!�w��U�8��і"�����&�Z i$���b?��h���L���������~G���z��^>C���'���(e�(k��P�b~|Ge~��Z��ɜ�'M�Z��/W�^�w�DG+�[_=�NES���+p�e���;P����7f
ҭ�jC�����c:U=�/�~�2&^I�?6�u��eb!94W���I��=� K��: �~�]� �Ƥ�/�qH��\�Kܸ����2��B0��)հ&h|Kł��<ټu��h�� v������]ʸ�J,1 L���$�x�^�sИYWM�^
��l��h>���7/��m�:��@Z�Y�)�G�GF<����@f�0o[�