// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:33 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hkRgPbn3Hovh4KdOhKChSB6gZI4VD2/sQzaHwuwrYo4HwQXlKIT+zDsGJZaTt7CM
uy9uLceH5DVRLXuwThnsrazQbQYxNwr3XphKEgi/D9RUlzXeDFyNccOqPZ12fBHC
OdfOQDrSB2lOUHjQyK+tSwe/j6fveobutDr3R843AZs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20304)
OsJUfraBmQK+M9Bd8vsmam5G5v+opgEYrQYV4g0hCxGtaSall4feczApQifhKcNa
pngok0joyVdvBDWgdljQ46ASzSKZa32uPJGadtDx+FPFRNVD2LNsEcNT8FaecJiX
sDANjtyh+SH08EpO+imtHUnjWiAExW42QezzWWOehGlqS3W6gtrcFW6+ovfxPrG9
swvgqo/f6AqIud8Bt6VhqyG6NPs4MoyxEd67K6TxSX1xcIewtE1DweOV+y0KbWtr
Oy12z5ZqsLYBAlnoM4Sg867caaI5GNV6vk5G1P1HXNIfmd9yHGncGQrB7IBI7ZJQ
KaoihM6NABSvUdOiWT018dcCHlK7lHyaXSjBTrpZItSObTNPZUYAfqFBmAirhyzg
IhU2bJY7ow+L1OVcFcQl+Fp1O/eX9bOJt6KRhGOvjbGEDglwdi0864Y95abemcSL
9Uru5cweyrkKIeymrIrFF0yiEYaQqEmn+SNvE4zT3Qiu/Q/yJW+isdzHlNpFTR35
t3S6RVAy7FcRqs5MC6ohzEN8d42IfNNe/T9wgziRlH0y01+KdXV0zy/DVXRxi+m+
s0UETT5RP4uARHzdL8K8IoDcDEnflE3TmsJEFbO3vwqK7Ys5rSX3690I2iE/cIL6
PULKIri3B+q+y/42g7Qe9QDb/f67ecsTXQQEHdYWFYrfRMXY5NJNjHrCu2F7Sx0F
aBXgexxDhJY6KSfqha1OAHVXPOmIS70U/HXMO4Kk1mhf5D4tFtq5UQlkGCKpHbFL
jS/JbAreUvh7REKDO5eKWxHQX+BJPbsROIfrZEc3ZrvA8zpQpeeX710N/gkEMZHE
XUN2fnpO7Vc5ZOH4gfFILj6CztUdxo7XnDC/1njbXeX5wVSQJhttvoiBtGi1qK4b
G0F+NPRhlzCDhISskDPA1EmP8GUwX5H/I+bAc3HbQtlpYWsLhIYKn6dmFRpV0IgM
vfhcfTxHehYikiUU9XT7fJuVkbQwgQ5dAau3Rezie/oLk2Tt2Gt0b2csxZ+tacOV
U84DeeBtqyByA19nZ2v7uy1VNfg3UNTlV6IL8Zd93Lbqzj2KbJK1MbxEhWsh9uI6
Y6tYja9ZWmScsNNq4pPDPumuGAZljgV92rraQQxMB73crysLoHxTvzEdePFEbS/1
kRmHmdfR1PqmRYT7gyuU9YnenymEUSKGqXm4dWBfmpjn2Eoi+0VZ3rmHF9k/oVZj
Pdplx17sclY9edW7udD7vwTkK7FS/I8m75fiqa1P41RA7LQa7O4XX0qSZS/acw1p
Yd6e+qiOVaLLQ5Syo7+DQqjHCzA/Haxb50H61LsJozro21l6borLe97C5WVUw5qc
Eibo90HpcDbSNnjQc1NR84ISTCs000R7sreazhgtvLQaCr12MtG48ZGjGcsJo3NY
pv9IR9z0is4OE581lI6Cq2QVOeV3M6vADSLX1tpU10cjClbWMKRomqX+cQ0JT2PJ
OXP+LaZzJX7b9NWBFNMdeIp22vjB/vkZDdSyEOVC3nqFBis09cKCztvbT01k1AEM
1ajMTukH+0Wv4XonpTF0jKiqKZwXHTO+g2ntahG4XxEMSFZW9cUNwfarH+7S21L0
xXDze0U7c1fdqQsQp1VdBm/FDJ99fpNfI7oy5/ipytSJv0YwQxv6ZV5uLnEI0iRH
z0dMlKCo6eqX/k6ldMjIfDmxFIpAwjXLp0xNBMr5Hvlpe9GqAQ2WbF4yhO0rFuHU
IPJksbuGEcFg5lCzh6N6vu4u2u33zmSYsLevZGqK61hcYzanQKZg9Ompbw2AI3UG
D43/EItwJotP0kVk4AU0cb1WTdMFhBLHPGGeEhbyb9/ytqO+C/Kj2Dd/TY+2iCAX
ZdjeigujTJEPq55GKmUvY+TAW7Dy54cUt/4aruTN6RBdSF9Ki0k/81b9Nd1IerJx
r2WP9548xb+aFkI9g8UnJpsWlq3XJL87xcE5axIFwfdQn1HUIkAqfGQXB11vrdIO
OnPIAPdkt/k8gKFQ/JDonalllYHKtVzXKH9H1pq6hOtNnhOG8BS3kmgqHRozFfDJ
EpLLaHJ7eAALgMQrMF00IsQ9elJLQsTun+gPIQ1GiGNvMWNJxNogscqImDAj26Oc
O/SEKEUbvs4Vbkz+sGZ1sfgfrtIy1OG7qgzhRsB3hAsX50CQl6wQJq35n9JQLXkL
b+o6lJn2h3H6tCpg+a7ImxTQX3z2fFztgTKjQccc8ZbBdBwM+KhQm/wvEFIsJmjG
b1QP5npyL9DH1etepPFCaXCDSh7syynuD0wm5sRgzJNkdBU7+B1Fs2CxFIG5hO88
RAbJrKJsdm3rf1TBiljsYrkGnN+qRS/7BBUyZcw/+Udl7FmyPc/RjIO+09qkVmKb
NCK8eROReUsKliaTaWcE+SNZB/dI+bX3ADZEftuAzPuA3vscJ48APDHVd/Hirf2V
AbHzXd/ofbR7X1Prt1gw9iUPbENWyjtU2zz234CeL6PrrTvfLYx2NsMI3LwGmeI7
3uApkWj7t3o1z73CkF119Hf0u0Zl2cQesmeGXDnxNAvXH4gT12keca5XnC7jr5Dz
9Mdw0bnrI7nuuJ/JlNaKBgN7ELSAiEMA2GmFhRZGyj0WDwukllmN3MMIDiEQT1GX
S0ak4Y+UM+TKXrAW8v0gS8Q/YRAmnLlQqPPxiUZ0ieFl5djlixoQMQeaQdtQbc6P
OIhecy7ZHZH7T4KIMs9Yi+7T3gMopcjW3rvrH29J1IW15Rf0bmEHhP+GAyw7734e
wdF7zZ4AjeXZFJnM9VP45dGoL2z1GTU5rz+l74vw6VVHuunnqIimRfbCChPfOrbf
gd/h3N0lwpXpEJq5hdvC8Wg/Oc4cZyVDJvaBdfYYXXqT7ARGsG4DiWDDJ/hwkfDP
h0Iz6OeJF31wY0+7+tnfFV033i4f6OAXdjlhaaikUeBWlLZLequW+5T11IL6h+W9
rzzjQCO5YKGRp6V9ZbtKlmUCBfZcDMpYuXOBH1bDyt2rZ0DAkvJPNBK6PjhgFLb2
oha2DGWHYmwQYLiaIMLnYrbvRZ1hXHs4k/nQMUS6zDllL3+6vklT/Zw1+CZQg5Mo
KgHKf0oWLTd0yQTwsgTqLALhPSDkYrVtHxTxOrQ1mG0UOSZPwak8rc+mIdkqPZx8
wYlu4+ie5yTnTlkTuuPoRmE5mSsmUHxKa6jJv73ptYX30jUz3/tpDOOySfTHV8CO
OQtAaN2S+TTHSdcIMbV6pyNhbIxLBtx0inU5SEnaL3gBjpx04sk4CW76E2fUKXfp
wTtIEIUizidcUO81WEXbqiKSkhN7jSXKmaMkvY914Or2buTL5xyo9rvGzwDKUqBt
oFkSTfp0hLhNWGaOPsNciQaU8g+ZKHhqLbpKO3d6SXZUJmkbAsCZd/ru8eFhTFj9
QYVOMo8H1kooiIXMwwmSt6dIRcITHK8unGfGdZG9i/LRA5zNGRp49on78OYi9C79
GqkUdPloIY7BicxjlkEJaP6kQhWoJUMNiLjKi1WtSA95d4vE87XxsBuTm10ZTdDS
Um5MXLmPtuCb4bUmF8oW8enKZLiw4Zi4kPww73wMEAyYzLVsWis1inWlpm5eE8LE
UyW3jGvdKcb5KIBztGlnXu5gZwXq7DcH5v9YnOmmVy7CgR9cJUwj5Q9rj/08bffb
hOVmKtX71rFR/ce/mYhIcx6HxjSeHC/Lgnq5EkYTtLgzI0f/cJ1OHqEqWZPLlKoJ
nbzwMapvDKbSjydpLuvPBqCa4xkFO8l3M+OAqpQbo0n79DCY62H3ZryIsez/RJj5
leJ7FoAG2br33oWFhudiHYinZFLcuFX95OC1BG+wkdejmVTMga+0cjL7JGqwAP+r
c9dPcVzRJrJI5vq1H8DV1aDl2jwDTFVjQ5Op/6WslmQuC5R3doJ91qUGtl+aonGl
IuC8mEOnxv2aBXOCZIlrLj0k7G5M2P7aRvjsc+dRXalkgv7LMJp9heX71EbsBCYy
mbL4JRV+sn8MZHopG8TGCxRPtDNEyjLHzVH6qwfP5cH2OiqEp9iF4knAZaic/1eF
uyFPbrLwJK0ad9fLcFq1Sa3kJprIulCYT4Xu1EeEgCWAEgBQqH9/uVG780Y0DHIS
FPLTjZXXkuqBleClhJSePIZu6cFm5xSkEDE3mtjtCotNsr5Z/s8xiVQIcCaVSPAp
ySQEOQuCJTeitRocQLljYQT9t/o9a1e7k/1HYVyQ6wxpWJ3tYrrByTQ5b8Q3bh8e
RMVLun/fvYf5d4dDMsv2Ihm+FZHWrG3SI2zNvzhmK6Q4UVl+82PvCKKLmhKX8MVT
WQKfx4XRSFnrVD1BO/F9JiQm74RKwdDTuil5p25lxKsPb46/6O6TbTKaAW5Wh/B2
3kjSL41C7aIRTBTX38jm3i+f59ku0oN4YQy/f/bHiIcfKQhNGGaPmgjOJ1MtbxbB
bMHpopiaE3Y53gCogTbxP0gzSFWtFWGBR6OIB/FL6BmsrL7iiN3XWNRgVtNax2qg
NSWzRwbPyaPuuGG7pn2l+T/AaeuRZXaEZP6wqsmFdAC3dTnFWLhja5v0RLLMvXf4
Hh8QVx2D63m80xV7N5BWdcI4x6qr+Mb29IWuJTyGxZFEmHn8wuB+eopViQ3T8wCr
HqFzAirWDHbV1N+sNvlSeYybFuDHbVclarQUGVPQaSPPHqPUGDrS1kBNJEiRUPrO
HssIATZSsI5869y25IYv9Rz4H6rxcmdAByFQdG2M95Q8nlBniDKxGDaeupD8NbMQ
r0DG+yop5mNFfpUpiiupHe8OS3kXBKKlfF8/xlm0lxcQbnjNdgTQSlDsckHBh2X6
CDiCLva5fZrIuuC0rCHEYQn+pXKV2/KG+fYUe4zlf6tdgziuUgVy4P5ZUbLbgAV5
7/3h3Vo0v0/GqPI3qp4XQxdkVyGoZEujsS1ZjTDLCm/InOwvPtSPI2AMerUYGX8s
CeOmLMRx/PC/7BjQ3yYNgMZKVTPGRFQA7IS2JqZj05FpeU1s6b1Z4HNdg4U5OY48
/5qPNcqa6SeX5X7yVyR6IrEAnT9qNdxrgT8gcEbLddAOWwvKcP85GqCCUhIiJNp3
lVWfODglxYNhOso7EMJu6Px6ICrLqN/laB/sWLpj6+7eXIPuNO731CuQaVnPi6RC
FDbK2F+BnZ2fMrRr3fvW/6txkwDduznVOpZUAFlDoJ4rsViQsO9dNL/hXdUEYHzX
F5+8P5nSKufnG5HZKDxIhe+2Y1oy6gEqGP/q7kMO9tmC4hFi4Ld5byHA6wUUGRyA
WRcXLo7jubhFJJpiHQjf3XguDRbcuyEkYmadfUcen9EXaeXyYJMDhBI641ZFIX76
Yv7h8e82Q9X5chzI16Sbpp3Q/cnpgvoc29RqI1WBY3L6ig4ckwPEoLGy86B/fdaB
j6yxBt9vPVmu2nM3Cp0JUu8oS70aVrcWhqdgqdTyJAoO8VOfeTwGDFr+Qe4zCCLU
7cGVpK8pKzXIEXbvN1dX1UIL5koNFfPqleR4GFK/XJnOTeIaSgQpqvjUpGC4SHuz
WVEKJ1eFKmLmAVfqLzfyJC4JSw7z69KsHwFAzlJCBTYHyz3kqV6XNJvvujo8U7pG
QnLfmv0kTai4WkwZTChHQr2nTo0FEBIHMrx0KORlSP1iIM3m0c0h47iz4dZUKvu1
G37XDuaoKsM7AU6CbOAevNS+FcS2zDf/grlGInqaEy2ahcZhIGTBiB0k+qPFFtgY
3u7ORmzurdkJwKKt2kurdXmFolp/7YZVegNhMQoLSJ8997K8vM9F1h2bf4QhobrH
AZ6dodREi1hXjglgtSDfJkcNhiMbN5VfiTX7Qwo+FkGdOKyeKgb7Qns4k9VdsOAo
cwLqYKNa2IEfeaT/FELe1fMIEasE3ZzlkOveR3YsRORZ5vV6kvafBeHtbQ6e8hpW
Ct408ecOXpbw93u162z0j3ruTBEZvJ/fjd8QdFhpdUlnMQ236/Sea6MZAH50a2UR
aii4K8lFLUi28ApJWkcDOnmfD12kWenHmEw0vsoJOOvFxVw9G/Unzsx2uip+2E2p
d3aAo0jg/OWZIC50kHra1yaqqGO9I0ghH04fnZynW1xTboIZ/gIM1lqCzDhFhBV+
Anma9BX1/s+cLiT3Y9Y6UrnuGMrCHNXzIwxItkAqsM7oZ/tKc/UnwuIlCaEJL97v
44mex3i6mGEP6mr1ZxUO0/Rmk+FLksyYh201RJdsqRPYiJs/fLDhmkWLDuE7FtbE
suNXFhSlGQdhtU2ITPNNqatxj3la6AKA6zIAX2mYpPVBoOatxkDitlNejb1pnllV
fTgp8aGewfdTOey9RMZUg6WAZdyZNk1QU+x8nqkRo7koSHc6kTVbpe5WshZC6tph
Q9Q4Oh83tcjOPIBITnXX9MADT8Dyi+D5XlP6jB/U8WxrsPiTjfhmWxjSlYPUSd2n
R+CPgUM/3STHvMpdwHb/DCG547p5/1TSmEpu4C9mb4+sdN14+fTTcb7vzc2HQDfy
ZCO90Sidxb5SN2fwWZwRxAdKKku+Gps38H+bBSpDIND2PMBH5sQdAROs2WFsvvCM
EsAOns93LWtc17l97ppXYWt8JiAGLynTs/cNFctayKn6QpePB8vkjDJLS1SPIKIS
CNNSVocyOv4vcPKK0kw7cAMgUCfrwYje2G/Q1moZ7nUaQ8XvzEnVdGDtyTyjbuuT
BdmjpYOEJi9twXEWTxTRVhA0cL/MhEnQdhekDH/dV0qsOiHRavAHQNqd3qxUXEk+
TNeS1tUIHNBQiMhqlFERYco6p+uEhHxkOEo6270y1wy2rLtb4GfmxvzZLKaaZ2SC
8QWFmjzNeQxf+S68Y/gprmO7rSzu+yrO9Nkz1FTOE/GYSd6yUThH0xalJSwwqdbq
jg5xk65YVTHTS566dJx2yoRSU2eeEVT/PTWo25ewQyO0OJzVUY56TyErkjte+aNf
B1fVGkOzLldfnvelxnY6cbFwAwyVDG3ANOJ0ujcFcYzCstKEHUee6AtHb/R05VbG
JpjkuMM6EPyrpKHPs52QbzKz2wuB5DJM2YgZfBVZt88lHMWyMoqD7Mhq5AOcQj4+
RFkazYUTVdDHJO5fD+uUIhrYPAPiQmLDHIMVOP+GYMWUiHPHdXeMswjjoKpIQ9Ex
5Jbl3PBs1t/mksDsjUrmDn1ZbtGJM3XxiukiQo3cQY2c8uIaCfekshQ2o5jGA1zx
miTUueSTMuOfqFyXUELlwPy8yHeS7xL5iv/QPb4wVFyx52eY4dBDAz4Y8FsF6cBh
WcWc3lyGKhqH0Afxh2NOORO5pDSzWaVXnXZbmQ6ei29zTwqd/vL4xuzo7HzpAQL4
asFeEEmHQJvLK8OEGWHWcJoQXE7FT7zCznkzW26VpbxDWMerzwbEHl5nqlOxMGGX
1jXZUNTXUryhcU8/plC2j4vhs8XcziipeYy19oajcpIB6YVTaPPd4rbSmKhVsFCT
z5sHHOn9BqF7YksQMLOZH5vMsv0i/bBTGQe2mQvztYBk/F4Zb7CPiBPGrqDtFHWQ
L/fqq/nk24qi3zKMBG1gaECdQnSmnJS+o18M9TJM5PAOY2P5ZwwEbXy9GIDjf+O4
ORiSrmeIh1m7nYaYy3aweY/Pbe1jIYZCtY+PSy267MiQiAU3/nYVouTTmA7WumfM
bknaiqk27Y8D+oKeU1MgnAkrW6YPd9iyPO6s8WDOFmqugLhMZcd3gQtaeL0Jrooh
0EUHCwoSOyxVZnKujUFJ49uaLFQ+ivQL6ykcO4w65fGnUyJITzZFdgJ9FJPB8RTp
frOv2tKlVCdKk1U0NsbaJiPDKKZfwbMf7bFjZ1J38pteR6f7WIKODUV0MlzImhwr
7iDO8AVVk9cQGZCUiYTCm/EbIsFmNYAH4e/lusIIeM54VrYiuUlAZ4joOERnYRog
K4J3xvQpMX5hPenRQu8blM9fVg321AJrswMPDc3TXi13TGpvAXvHeMQ+25Tsz97k
Fch8jSKXVvEo5pTubo/lNJHmvPG3NsniznUrYeJDshxRpRbdFBKceXD+FVVOUUj0
1P4f5/7dDfBnhP+aPPxQ+N3gBaWAOB85/52GHEKNQjlQEYWJ9Qze1PkRZ2ryb9I8
m2aVLnL94naWrRGttyT5Jo7SaGmJh861+guN0v5rkUCKi2ub2ztUr6o71N7yVp12
6+008LLSv2FjhZ7e27oVeglCATySbTN2fmc7TbGB8myCKuMEaTghXoYRRba2FRPj
G0t75h9ka8gYo4F9WTabqacu7sXiJzmZucRNZEZgKgEi8iO4eoPh2GhyGnRazRv5
9ltjynnp2SMHYOTZiBslol3UXTogriumf01TXFlPlJfo3fZwXMNBrFE+ygxstHcS
Yfgrmh0LP5dtiR0QcoXkmVFQkwCJ93rPehUs3n+ORLwS6h16NHssTlwrKUMzd0Wu
nH2d8gs0V8x3SzKl/pf7l5SZBUMVJxtA3I9zoZqkz0qqZtntq68jMPfeOqhIUSid
olNUOBIeXwtsMoMja+vlSTCyEyyfNKEQsKSWqKrVhN9Q43/qZpYXujXVDWKlcDIn
Pl/JMCQlICW/lnkOLkUZp7EDdIDzakmZnfITpx8iwRDDlpoC4C7rKh6Ck5jxQTXQ
UZJ9gH3RZyocF9cAsQ+litRp564uz02mSHztAKau2vrz4dKpaDzChRHzZQtYaYyd
fA6JU4dR0gNSySlQFgq1NPUcqYRWuRtpoK0poF32krFsZi/lhTuqWOvpjRGA5n7e
nTgexLM1UuqQX9mpA7V+n8xSqMngCYD+YjMngZfphm7nwPUPY2JRedwOT4T6OGw0
hFyZjYONinkCAAfuQ4u3tMluuIrYXixk4773vlzOjOqzTiFNi9KBp6UTIqba37Sb
nO7ygwcgzUApkziCQXdYpb86vFyJYucl2fTh8UelVtvkweB8ByaJb4WN8mFfpvne
BoZdDGS/0pefq7iO8s8AOawogQA6SkhCFTfHqXekd5whQ8yFH2q6kGCWP9d69qL0
qr7vGvCKkO8VVsgGqrC0w9K/owJudLvWHaNnKPr5JxV1LcErpYeFE0oYoh3fUVoy
rS+m4TehkojmE+mJeChgR1NUb3QAHGHrXgPFUSv3CNQivehdxsFHCHOqAR1rrXNJ
pXLiyPjSPeUD847q/bC3AZfPnxmUszrUMdPPBnnK6bfjk4td8E78sneW/iX3vQXa
5TeTNtrENrwI7wH5/yZYxklfeidZaFx6LESMd3gmHts8fVt0eFwRgmawrd6VRsKG
ui4UBITkVspymDSJhJ9YOpD0OgqAqDA5xYY+XwSKGPgyQ0gV58XpBXirgt0tP4BJ
asWmHPg4jzLqAXtXO7G+I9V3mF+7UO+8QKSzU9y2A71amSDc8yInLPRuZnIwDD6H
Lme31CZwL3Rdfxg12murUEwHiuZmvPS0owKRt9sf0xaQaUGknQFPqXBYXO3qxAgI
nr+liMUUOKOkzmUIPbYhYzUplOclx05HNxQQEGKKJlz5wnArgD77E+CPrOkOG51y
/xEg5TMyTPugVW6dQpZRrEcUhTLE5+q4bkOTRHwr8zO7nhlRsjgz4Row+Enak6vQ
jhn3dHAadG8Iz66Jf4cYVwUxYqZHAZTOvKAQbymnHyu1h0s3I7iJqgg7Ij3Jt+CA
8Hg8KQuZ6wd+iaVsWkBlsp2f0DB6qCjtWGpecgrV8vNyNdoh+NtQB6kMqFgIGOII
k6LwD3G/+ofphlzED3yljawOSgVNr8KB455PesO/lWuEijt3lOugNt6y2M0XPjoy
hzI7UwyD5wx4O6jH5eG2gjvB/YTXwIHk6MuYDlA/PLEIJ0c5TaaU0/IDOFUJ3NpJ
Cv4dEk+iH9tLll4DBDUzIz7h7uRZvcRHJh/X6voZRGCUUHXAKHMe6HI+ReM4sDZD
nLO7mpgAXLIRafZ+f/rne+UN0awp3t8Yhg0wTwV4iW2O083yWiDxIQxBvSTpvoPD
1C59Z9ZGhZMDZSXEGkBNA8NgrwBOTxZp5icHDd+22dwN+DPR9Vxnc5UpxtV+FA1J
sp9vPkO7j92rWSeI5r9wgrRRi5VZJdBNSOfsZ1zuhHeAwAg5GUVRhNPTLQlFyJBd
hu6EUYCX6aaIqUxKyrJDV8XWqNZU1No4IY7curBFpuq7Qv/FOQDkXtScBo/CtF24
uI+de1/UJM0vr9YQoPkXdxrKuQ3zkPo9lhSZFnvhfQfXKfKdXOIZPQQLUnV/tBEV
DTZWfLBbKlTPzJeDIo6i4u8MAYhROZ6krHsaKiyjT3hPcLK3rL5JSXRxeTcIgC80
F1hUTXT8+xmZiiPPYNhfA93a44NZOk4teAnJz55DX4Z+ljZkQtUU0HSn3Gat1dIa
8te2nBSszYCrbrR+8RhPKXrxeAttbPTW/fZUbhqdOiZs3VhCcHY6Kj1ideQJhfdY
d+UjRITVqsVVnSgfU4d0pBAJUsoocem5op+qTO7DL4XXv/eyzFJ4nDolNiVKxX73
UbSszk3vpdqy835nR0+iUXv6mK8nmJeU4+E8wmLAZo/J7RrH0oVozdh684F5hBmr
n+4bbsxX+18tSwpAoAbKahmW3jasCMafEAXGrHtJAGY2eFfNrwr8zpdH/x1FXYJP
+lTh7Wn9gmnstfx8k+iabnAun+TCg5dyTAazLawebW6mU/XHpNY27ySI+y/f/StP
FtFYu8aNuxE9amKy+uet6SmdJ/zjd6EKEZb3LkHvIJuFfjlPpeUvI8ZQkmj3gIv1
GZDh/r9MR/qc0UmCkRRjdRF3LyVQXwBYkDzhUvjUGTToDYOWGrcnVUWeOGaq1KCK
gNNIbpgLvJhsiDPj2cnWP8OHDP5VJV30qjELXntiTOabuJ1x6SWiYEtyaLJw5Nut
hGYvs47DdOslLVkrcL9G4Bj1h3HhkscAJKIf5YJLWQv9hwylDTblSdzXg6r7KS9x
dxaHb/hwxnjiF9kR8M/PeN2foEH73G/mnhMw0kz1gqxizrj56qcGoS7P2G/M147J
lHJ71Umjwq+nczmfGcDptGc6uoqzv1bkpE7xAkU7n16ZPBMmiKk+ZZkh1bHbmuzP
hbScwCpBTeODx/3m4LRmzf7jhKyorG4/Fc0p6XFYyAiNU3s3NlhAFzRokzMOLcRI
kxbYZvCyp88hPmSppZChjDHL08Gr8Q/mjvZU6w60VyjOEoLymOEtvCunnqfcCjYs
Y4eRgxAh2tMDPvNc8IgXer9h3KgW/x1jzwF2upOlziRqbXMqQ3OE6P3xTQ5NBtnH
RuVPhwfj2ocb2bHp4f7f9Sdpo0JppHjrx1+0Kgu/vNahnDvp2nFocpAy2ZiREZfs
KWoFzEjHtaxq1ZvpViCIpIy2lPOjkYVsNsnengWd3MoppuxufK+zTBEMy6N3gjiI
adNg469E0DOH4foWcHIro3yVbMH5Qnb5ZoS8ImPds7oT8ItVaPVXNW5x5DpGo4Nf
VNqGtD596syeh2nY+oSFf+CAhJgmxEl8ekPCC+VzEsd07m9XI4RgJ3jAs6ZxyaCi
1Yt3bZFY36ancanznlmngrHNKnoFV4HHY6B93g6A9z+Yw9WW0ZXHD714k+RfNGtz
MLrDchcI+J112LyitmElTlkmWFe3bmxev8GMAeXDwO6eImLULf/4AIq9ndv9tCI9
HeuMiPoLMphvn7NplrLfxSFifxphITRJM/Goo602vcPBU4DXmUe8cOLOUbBkmi+G
CYsD1qhzYM3lPot3fP7aeQxiH8N2ZgATMLrZoEe7E7yBMbYM+/SWySM3wFyFpzVy
HUzVlPDGehtIN2t/pp45gmO9ZsDy+dr+wilKNAILqXu4lqq9p0XxHUqKBZ9nwGf4
2bW5CmNaSPD6A1F41EUxrVVN7hZwjACuvwFYb7bDGd8i6KfXgP3nxURZ18DOMoUR
1AkElKlOf/4zcz1nYAKNn9cpDB1PHDGq5AoGdrRL6RFBHBTtzX8vqY7VSTu7oevR
RvxrCaL2uWIbt86+eazHisiD7l1KSNiY/xjff55kWhSiSCgHoQ+PfMcJGN78PQXa
l6Yjt7JZPsVwv91CgzzrhnbrX9vX0bco05gsiW9HjbFP8udILQ5DLlF2VD8vnVjD
qjA1bQRFvNSN9bFt9dZeo8LqIx85Gk4w+roAiq7CsUu7hBMDPWnLSt7tcWRWkPEc
fNEJ1Iflre2EMYUZ+dy0gVvDerZxoYdGFrJaIaVtVaVDFqSrIoB0NEU2P2qqEWYz
YDadCZQfBCt0l0u1Iie6kC8oQ4G0whpf1SNix2fVn+D223IJij7vHloKTu74aCa/
IYlcYvwNboC99Sy9vaGH8jE4XR3BFVKD+RXK1qL5Q/sqeMpUahk4W+oEkLT9UFmv
EC6+ewGIiCkWcn+OS9GgTawxKYeDvAhb9wQON+2/KddcRvhSMprJ4so14H8IgDLm
6Np+UOda9N0dLJvwHzJjIqLgys+y73bZhsF7/Eby2I3qhs8YUny9rmuWLEyaHyvO
ZjmiKHk9fDBYiwfEyLD3p79tsIpAHzwwXAGg2DJsgytcAnGG6H/ZfSU3G62BkdmR
9vBpzdPEMj2afV7MN1f0wB2e2MmzqO6/sR1lSmVJdIEF16GB2LWquY+VlWmmzNUU
ND+/Xj0ABlKArteW0yvxTNnGKqDSFHPxAiETLvWU4WhdZiws3q5KVoO39X2SpO9+
tYQUeDh3LEHVFPn5DhVhBxE+2AheDqhYQyhcgusKcexAGNgj4JcXnGWfM7L996fl
qs7LvLTPKYG/feUrDhcZmaeVcJLDlt3Km7OwhJ8csI8TN3v/V0fg/5Yeo9U/ebXP
2qcZA3A1xRkLFli5+Di2FJPtTGOX62hRpR5xVIdajV9DdCe1E1vrdK6rbMlf3es2
dRaSklIrOPBbKhcff+ic9HIUCe8Xt7rCyI8+FoY0QG4cUM1g1h1IJcIsN6NnnB0U
NM9yYFO0LHi7q4g1D0VZDF7SyDUrT4RcMZ2szZEItHroUTQR3h043simznR8apZl
tuQWM1DJ2vRHiJUBssqtKeKlUX8JhU/bOlkok29wDp5Ec/Rrbh8CfNPFaFTFQik3
JxzG02u3EvyMzGitRW4qPVjgm0pGktaFyJe1xFMdwl1exn/whb4M/HGiITbdoll2
WtIKmyE+cD/vC9GyIRwkNiQ0pSQGZ1boQnMvyWZS0+bohgxKnD/oaGmEv99dmxRc
7ILwuAnRNLkmAWPSE2VbFh8H1p1YLa7YSKaG36SX8eknuY5LNDhORoQtH6h2vNIl
TphO3IfUMyOPAxEZlC0Ip0I6zylnFwJtEG/wx4u9iUqhCU29fx4xKI0+cve21h69
WgLaACZE1v+H5NI+BqTQeAkrsd2rwZcT4qc1ZktAXK2ic2jZ1GwIa7vb2vksXG3u
MHa2U7fhmixzZ5AWKXodesO/9aziARVqsBak2j6/6xattn9qKtcJj5uDIJ6OYl9E
PXibtF825wORcui4/iCK/dnFHgfIhpCSV1/RI96lL6eAn+kArnr4CI6QAmK9zHCW
yKN6YN4+IC6TND1TeNASTHHNT0peXLv0R3e3j2XycKPh+IYgPfhtbe0pafbIpy4f
/y+FY4NTkptcUgT3AhK7yobchrfydf1Es93Eeaafja1DbpJkFrPEWsMMv+owCDQR
PovdZhPk903oQeTKEOq+gqndaPZRDmuipgCJVT32f0kLqfNfD4PmSS6enw7hhTDo
vhYWTUp9XKnJkbvuBWT2T8ty/Su2gnaPKqzybr8BiI67lNLFyiidxuRlDjzgEn0O
dBeVP6pFJDvw3eEajmsTzq3M3OkhMdUyUa9bjVSh+xdhR0oUhQZDjBm4UBOQhFaK
07+BLnS8mamfYYX60Hu8GBhwg2tr7wnCqOU7DPBUnX+K8qNU6XRSMiLZlHwojm4j
zBXMSuontaeGjj/mF4ul+LxGJ8QnJHOEqSQm+7s40nG6jDjVzMkgfQ5diZ5Da0yW
9msv1pgJdnEIVBhOrCKhX2T+33y52NfkvosuUPsL1sJEmFLpj6JTUZFtALQmA1T/
NoqRRJZbjtWpsHhkbkorMVkU0Ghca7TEdCDQHuRPKqB08XidmNtu1zZbbQJan2U+
G1FpPBeB6Ln2lotGBy7SoO3JtG52CNjy0JQKFaouBSGX6y9lx/Tvt4sbLhwQlJjs
IHTUhT7wxfXndTVj2PwUscEBMk464cfPg1169FKHpj8Hbm9knUhfFZHpBvjmW5LD
YgJWXeDDWJYA+ozOs71m4mTgy0Ig+f1Uzdb0AUWlOIOxyB24ssZEyt5uO5473UUS
i7qSHOjLsBO+hBLf90O2lRO6Dq3ajqFd+MfBaBxT+HCXyQgtezRJtFZ44Mt72JC2
w7vHXTaNt8ws/45WGJEIPeLcynvqpd0On8UWQ4i7Ql033gtCgswkcAV+dwbFBr0s
QRl3T4LYYouX1s6bN7mxMOOhfOo+wVvDuky/obdKdEyo7qwoXCG3NRbFdmywJCAB
gGhm3urkR7aOZEIO3OxszqjYe511BUorSSKSQgwOsRZNomQn71ZNDGR4b29eOe9v
cMG3NzltPGPse9BsW36mQP4RYxHoykHHUz6klrIk27Tp/VqdZymvNQ6kcHB2jy7J
P0edY3S67Ycw5djKMcaiggVMgmUpmlWMlynVTVRQc3pbA1cPlVIwzE9YF4d59Jpt
h1hzJhcZMvOClSG6x8j4nN0wUCRmiAGBruz29NMfkTnt5WxAvUyLcYEXRwVhcRDH
OiowwbZuPVUd8UflPJrrIfAz9YS7TaR0c13IeJ3d2uQvmB1ERuXHShbu3lqktDxC
Z2ljJWWdAsOEhujET95c5FXHOklU1tmJgSaNXdWm2taj4+r2A1nZqIoAIHNldVv4
vOCLduU5cpGDR1DpRY1PmXQDYvFDDt9DIMqGHXqI4akcaKP9lzqkjyzZiW5VuaUR
+wMYdZnUkHew4Iw0IRa9Dxtwjmb4QYOvhL3AvHCXyw410i3uf4spqUwoQ70sQZSL
/cwkvY0BfqTbn4BRL5B5DWYtyHWgmSya1nTjsk0BGWgRptjO00w7qy47XOISc/74
L6kiCBkVY9NkDTiEXCmeH49+Ldi5Xad4sQMQhp2VTDgf4Myku54zKOZt5aXynjPF
Gq3MkeMnPUuddox0vgMqXooDdpanuy6tokcthsnlMG4qMRUExeafAj6WBtekwa9C
Cks6WROQamceQsGo7nEbqTwunC54bzLgHYAs8PEH4k+AlLQwSvKnpavgAIOxRpWo
0QLG0yNBwlWTJz++u0gd1qWcyANu/7GiZSi6/tKoRSh6o+kiJBCYEY1ahhgqWOu1
VEakxIbx/HGguoCsXpD0NPLBiv++ujdbyUhLL6sIffujUA5PXZd/pA4zF+HVFKMu
szmqplzDH13zjYcVTwlC+E4qnfp0rmAGIsyBVJAiKWvJhF+LqTzC+d3QrP8iRM2h
rxhF5Vco+gXBbCOFpbLFLvabfFsSSxbE11LK4rnOXOytzEuHpsToqGXKrK5RMg9b
0qgvmXoHOMXCxNzrCtAJYmSZqk4Dwn7XU+pdTfmjDCOKSxgSLQPbU2bf/kXHEa7n
MJ3e5tV4VKAp0U3Gz3BY+NhCDsIVPBicqMB5I9RnpGxsnn/JXTP/lEQ41N59FM5z
GsqFXQ7Ky0x7XeV2YVtUUASzgpBsq013kPW0LnlYEjdyWMp77ksemW/fFDNIox+o
MdPYvq7yDtwyhOi2TgOhkVoVW2YrH0zeOXaCmDy9RC53tjy2Bimm9G3yfROEQf4Y
DiqS5DONUwqf9nnOcbuKkbyEywSuz2sPqLIGnFcGBJZEpAjlnPXIIAfTr4H/JVuf
LLa/CCgGgfVnIPoqsGLHvwsXWttOTCXFpZwlQnEUndcZ8uu66jR+TD8jIWcbKsjQ
vqHHBs11Y+Z/MnF6T5/TyINvjMrq8FXwDlQAW545QGS/nohRXNhfeeMvzV40fKWM
kPa5e/7eHAJhoNOnl1LfXZFamYLgyYffwx4ek/Efp6eLOG26cgcSsYOuCGp8DW0J
8Iu574EcyeS3XKEEcfWM2W5zWiDPfitj1p1xzOiY+rE7fhNHqPu2eqVn+F9xvazV
eKzyS7jpn1diSgk/34XRCne4CspMsOxoY6Ygd2j4/dNVvJAwlm4VNeJzFfbPw9xj
XQd10Qs80V34jNLQZNycGYoBA9ng7pBhRi1nzNz76QS+/tPl7+yNYh/ZtpVRWRu8
KgOCgrH5g6M8bkKI3boEDnIwwmYnTP1uZi5KrUKOlzAYTHatynZB7lMLfJf1cU0a
uKRZ9YTXYxXrRAb74A7575sm+VB9b+p2JIXKZpJfONLNVvme8AyrebRWqHv3JgFE
iTaYy2fkvOOXXn/+mFDSSSjn64m9JDwyEWriNR8EXCHXGhnu2L/U93p67KPqLMi3
a8xaMRerudjRDcAzOWox0aWrP3FHry4D2ImT2SDR7i3nEc7163n0UTr5vthS9emu
+Z9pOS185EmfQ7Sj6Lgt2ZnehqrRQU1pRbhRWPMVSQ3MoPAdZzJpINLl4VBD6wg2
z7FgIld7vyxrXlDURyVg3Dko38aAyV8wP2axRdsiu6H2fINitb8rbSrliB283b1P
/zTlKeSgCI7nDtXTh8vT7D4ISpKzMgzjXpUpR+w4ny3btHdVVV8pwhTZHgaraD34
stfNT74+hkRFtFO2s9JXHHmUyHQIB+jkWUWv5GoxIPcy1R2fIAfH+eRvTxfq7GFS
gu2TZD97xFSTPNVQXJwkSJhrdDuOhFe0P36wDY2DH8JWDdZDrwDsI+yn2247XbvI
VHeVuXLM3xvqtOXHW33ei0gI/8mkuzHnbx6E1+KIaxt1udhTS/QkHRO62ntNyYeU
gHNgmFXFPbxyJObQFCGym24Pb3ImnZRpJMYCJWbHXHVFVAw6ayZSjWWtCII0Kyue
Zra6Vfmd7yZK/5L9CKjT+hAm0tOBSAm1vkQlm2YmZdFHX5HyL8qsPriapu8KlVwU
xPWLJ+TqaasSk38jGk3xUxx8cBl5Uk4CXf8Y6AHpL9QfHl40ixbZ5xWXj3XOVupf
mnHEZo9LVIpP0H3p7dFcYFVrXUMlJqvaGE46C2ebjOhIcHO/S6n4me+l1DdWO7LV
Yth3X7oFR1zQTG+orzvJXV1bJnN8MFI+cv/w83PQGJLFF2HCKXHFT2HS5+K3y9kq
NtkvzX03Y7F+PEH7JOgWvrcW2j3HgHyLSSqdsNcBVhrOrcwiU64Z8ccCICM7oQ48
DCqNet2+FHCT2SLsnpTwhZnM9Zg3bVmbKhnNaCsxI7B1Utk87K3PkSkIEMVkFt/F
GYyqG2LlFsIiJhtNxAWAoWnRtCplw3IGnKONblOwBqPLKJH7Sel+MfkqLQsL6j3U
+KfbbNaCDh6Lu3ZTjF78o6P/q0BGd6QlhVi1jfYJuW+yAmprvSumcA7qV+BO7dRy
b31wuk6A+QjLYe7ur31lQm3NRyfIGwsZuhtK+eOqMjiAfVtFY+TVz1uWSLvBBQjj
bJ2nVhpOKHSQ3uTGr14gWDIdlohi4sycbDHEzRr/t7v4+w7JwRMvEchBWItKhYjW
Rj8aYW/p7Dm80qo+NdNhMekkQ7ZVbcehfKBE49vUqEyKh4TZ5G/VZdhPUViWy9li
juqSYFftJ/PGcklbcPFwLMRHABbrLewPHhrjDQtz22fi9wTBBDDJZ/kj2uPW1Gwo
VDHEn3tpZ52CqdPnEj7d1UlNtxuOjNcyhW3Dt9jYQo2KtgMayGYhFUsmnDDnw9ai
l5hZYWh8TlvZRkbVtEdPxLqw7zr5D6nKo5ANqjMfF/be94XlMuozb2efB0qQeRx6
5DjNxclpLctTdw3ojE85jBDNk6T2Cdsbjh/XpsGxcKRY3umRqoP7xyIqVvsiPnD4
IzZkyBJ8s3ss92zyi+iRaEb9NvtDwJGKPKGoRvxozx2wxiSbbHMBlXtCPQN/OV+1
LXWJcs771B9nKI7SSnzjzmdVq9zOrkN1VLwhTLwmFLTTUIjsia/DMKCaIgGhfGut
4OY8HYUmCDyUS/focYNi9RLZCgQhqbeXEANpzyftcGjZDgFte0vgqdh16nbCdpRi
tDJLNCaExoPteMAD0M5pAsasfftlFae1/yGngKJ2zMLPyR7+OnXL/TZdNtFKl5ur
aV1s/v6c/ug/uJZwRHkkgdkmfao012JCpV77fg5YBp5ejnhO8iZFc3so3DUze935
iPrMwCU/TTs+WBFrZV8L5Q7/t1dqlWCJMUALmtBJiBtvGH7xs9dZ3BHq2/k3xjih
7Vc+4GHQCPZnsQ+Kte+IVtxU/srtfWvTT4mHAIlmngB2vEFrUGqtQWDYkaAFuEah
sPLHU4V/9+mgmlc257VkCWz90mmGJ7RWdBw4abbKYkjvcEfAXcS8rOLnZYZ0G9Kn
JpMaaffuTlLnM25hyWe/zkO9pgSvaRODBsz6+jS+nGaAbhgZGrSxRZRPbJdQ5nT7
ycoqJdjj2cigaMvQz5vgpoRbfAISx29wPy7n4dCPW4uuOhm3bIY5AxzxbhFlSxg9
W+8qnvSBE01jZZjCWGbBD3NS33pxIC6FB5SEsTi+6NcRHxCTPVfl12y4MDGGzy7J
JPZLQIIzv/ZpkFs2J0231bfYFJfPjYs9aAyycA4qcc+53zYub08sdlv2f+KLwC/N
OFh1ouqcqWPMkHb+Y6YbJsksjJBwjhmLkwPchc/G724Zq/KhxISoNE6KAAol7qdJ
BJv0oVvFki4Zr/CQOYt9O/sJ7PuVpWMsqu5zTvDVkzDhONlAIbtH3OFnWOulmkZy
XVo94K1VH8dphkh5/zUkJS6Bke4Q7v3ZeV4nNGC2yo6IhaKfZ3QKm2nytcjwgZ28
sDXNpmDsunt5brPT74wmriv1pxEQlM0wIDkh5KoYzpvkY+zQKzLjWAndtjrfhClc
ufLNZTycs3ElTt99iyM+Rg8GS3Scpds/pK1B/7vNqRYT/hIMgeXiCw/dlHJia/+N
K1yvDiwU+hBBJVqOutuFF1KtuM/E09vWjGbOMELFG41fslIcczo5ug6wptDKQ1II
U+qamPNgJHoqV/hz8asXpDtdNpYnHH07bqvaXY/I0Ih4lLcoDsuO4mTrypFjwjvZ
ffr2uLJfrDBrQwjteifjnP5+OTZygru8n1KykbMbj+12JBQ3iLv2jIUhyOyrP+sR
v2/u63/A1qNh1ybZ/BxhgOswfQlyey6+JtsGyvRTPtGZl3nUU3D55wc3gF5PjRM2
1JWokc6qpp+qIb+RR8JKTjvyqVYyjhv/hwQ8WMKFFgBAd7ZIlTKfy3tuQ96s6cQp
C8RpSelm0GysgqeeK2xQsWau4CCnqYw5BAFpUk2+Mr2Ay9p+BaDqlb1GHNoT3x5I
bcrWzjhXkwGTbocIB5xA8JypXYZFX3Es04ZXy7rz0x7tWYyRRQ2B13/3c1FHOvKW
ukVLH8xg1xu6K7rN7SMEFTGj6aR/gkoTKbBguHhVdJAkuEUa9M7Yc+mH6dejPijE
TnmvV2CMDLC82ccYJnb1XXwRpTnInpwDVcZdl4ULT/VH5WqQOqJ66+2RgDALCgg7
20xDOHGy7fzQcey0AJZiMrf6aHNGGVSZw950eF+HW5+knE79iTHYlE2UYq2eCy5N
z/1BoSEhsA5OPaE1995uM9T3jDKYVOAqeDEMnZ1lzQSUwjf4DEVIakQFCk63Idf+
tihJjg1/SQg3/daL2CxOFvaQUmzeju7rod5eXlOnNIfGW6TXaxON8R0gFy2MccLN
0GoUn4zZyJs2oN02YhX6byyJIvwrJKtY7xujUbfIyp7LGK5xRfLSmobHrcNttNWP
e6TZ8Ax5p428iJh9iZHYaTGTa6JrVUc3ppC4cM77HnKop+pUwxLikG1tK7UqZ2yj
JUv3xc+dPrDUjlCz0oK1GtnBAsYQuZrY8FYQAxBu8snzt7HiSf00khSHxRmrQoDt
ZYHPNP6/Woglrgw6sG1I817RS417kmYMn1yal3fSTH3ttGrK/HsCqDIeaKW4Wxxv
ecNeJZ/EEO+5NaCEH9Jl7YcB9Hj7xkT7oLv6W4qeOEBZui9+agRiIFa/N7j0YQDp
TjIuz+PpQ0YSa0OkdHJpfyovDSb8E97nBMkJO3VDHtfGr3GOuOuF+RBHwai0w4b2
HGbshlz40Ny+O3hGWdrPhJ2bNs63z9ot51ZqzCHc4mF6FnT2OsWoFwVGMF7I4qnW
1PricumBgweGaiFpQf2m98N8NCx9F7ZgJhf6nFrUnM+aGxFlNWY3icq44Jroh4ls
lu+kTvF6u4HoiGdJ2vkUrkf961NAIPaj5QUSjJjiNyADi1FBFL0qJPxxQs5ns3TF
K3yu8UxdVeP9OemjEVq8ab96OFXczf/yKIzIiO/XNCv0FIStqLkW7SMUoQCNrwQu
DVQt30XD97d2ObnAKb6XJbhbpQbStiqOe98B5nN0cS8kwkAaD7ZhLd1QCoq+Z88g
tjTDa+scM68MtjilCV7xUoZAylmjt9T0HJwBhCaXpTe2MpXAsy+Du+UU6aDDchrr
HXvHg4GOwj0xvl2gXwEOtdBDpm/Pumzb8upxTvcoMccgqnJKvqLGVRbFA/BlZm2P
TdxZxa/lz1Etd9DI8kYGmCkBkdP908Fcxg9f6O1U0c9/wfU1ns1jYxtMyHPYcTXs
ygdS16nZ0A6zYMLyEcSxGHxGDDSV+a7VpdBIy3iwXWa8ymk9DKgpnsxlqCzM+7fw
ssc//s50u7JUYW9N4nZY4NytkUj2+WoU1BwORX56YaVksSZXog5CLOcPbIsp+/Xs
9To7OHWDj6wjyhJziVaB7RRI61zVpLmb2qnmbeYbrugM8ChWWtrTEAm7uq2YKOVQ
I5xd0MOLW9zyXwLl//o8z592IL9gYV0Mya/0dQoH+elqGUg+9ww6jbYqOXgejoi8
eUz/6rl3UwurqaNwZM4Oh7LEqh76XFliUVRvMG013TRMAohchpArvtCY77pO6D2C
Cp22U4nd8SY11O7JcATDu91/EV9Ojey0fts11Z7xbj6BQTKIahec3xuxE5tB5VOc
L4UQrdeN6hrSZx4BHFMztxcIatpuPeULwNPhfj/rnpw1ZwfdHoT4LGBW8zDN35AD
VEoBoCzI/MzFEtsWxZPz9BSt32cwsltOrmwYLJd+G8Jf0D+I268ctPCeaskTREfz
ljmrtfn7FB6jTUUkV8RDc2zQSQXZNmyOscZBvV/bGikwcBdZ9rzL0W3HwggMusOZ
sONklDSb+Slgyw5dp4cvNHpS4aAlsHzw53qRpsFIAf0PIrJfnl+ybKfAO0o5Qq8y
swycowS7CKCHLru9R6U/cvT8O/tSSQMHZF/dT5T+RjsZTc879EELPn54PSwaalPm
imZkBav60sqxMIBprsoHv64XiL+MQi4m17Y4mlKGuwXM5sG7vzC294fHd4b43I5D
QsNTF+CazTj82i8g6rv1q751DxVlg9NNLDQZBF5k2qKUZ1q78lYgECjXXlYR4gk1
owA2gGfRejEzYxlp8VRp4OGnDHWfMdsqdVcuuM5H9GgIOE9bC54uAUPdAUHfZn7/
vXCpQ3untVH2vIXNG6DVSB6vtyhq6VFlU24JNV95a3sjFV6YmiZ6BK6H/PIU88qE
s1/SGugC33CcfErApXLakGvTeNLaPebQHTxVo2V9hnhCM+uK08rtcgCqmTk64qtZ
9Zs1xUh4219ag1GPycreRv3LjD3OolBiQDfVikqyWb8yVwISDrZ74ADDlKJmXvV2
hzsVchqzP54jVCbHIioR/JjkFOV/s0uNoJF459pM1XWckaiUkhnIMAViAuQipiQr
jI2UjjUGacFXtT/cNkdHD/yyI5MVylbyMzOyK3vJvgZOJkgS70rQzKrBAEy7AYxU
wIE8aa9FEs/r9PATWzIu2ERUKKUfJ50LfUUtS5/t14Sl5MhnNS2LoVoKZLhqMH16
ICdIqEiZE1Kei9UOhKfLISRe9vbIpAgU5yMTcxjpeqrU+4p6uOwl43HE8Im7dLAT
QPMWBV4kKOAPa04bNQbbW9eERo6s9Wd63rWVyUofKjXbTuL1eLhLQxmhkVLptz8t
LorBuKQOB4LVvnGnbPtxAD8qVzy1quc7qa1QnAEZVxjmHIbqOBVSfxG8BUHppZde
eq/ZRBXL5HBh3EuDP/HNEOsxT4IP37Xt8Ehsk9mMqe2+b/9jgeFUJnWNgMimhXq5
19KqtMnICQbdJEb3YNMAopEXzNJ7dcPrN3hJZg2Hk7/4Ne6k6wu9xPr9J2sZhD/8
VAI/5++30CiiJNCHzbA/rSnsrs59Xsm9OXH5dDDs0LqjO3JSLHlpP4kC8Ykg0FDo
uw0rLucTStI1mt3aHKahe7CeHKIJI3IKX/CzXCjOJxqr/r+z38jfITXaM5ri+Ot+
xRqi4ZFOc9wyEBzdYYkft78/AL+ss/0ozVx8GB8sd54WJLkmCXr5/B991A+8FZ2m
R5yv2rsaVuVFPTBGeV5daL/Tuq58YTAed4HTRerBjiwTmc1ECA73/Frv8IkFMQ4P
uml+5okounZNpNET9Ctt/DOw6U5dBagL21MLhvKbEUxrXCGvGY3lUCff9DRtw4A6
oHC9ot9B5GGdKKEAscMf1vR2Bxv9djkn6D/0P7tff2KBpAUqyVtsXc5GYUARoqoy
Bi0TlsaSeFvoE233X5YqmLQwJIfFtLFcI9qDCMJuhUgE8q9Jrce2G5MSTyfWtwla
nrEWjfxxjL0PndaUuP0bql6qurb9VTxl6ThhrjRJnL55gPAeyt9BDjSOwbRF7ed4
YW2Uw4hTRwzq8wj+WSZYmjDvQJm+o0PEFtHcNuChWRUWz6ZM1kCsDCfNIUu7EmMG
Hi41woqdMv0haOzCFiCh+ZItiKDYq3HHa0gcof4Oo9HkJ0PKaO0Tr6zBTbb7mzLT
IWOhugb9QRZMogsmbeoAh5eNig2P4RwpDNsO45LhJhI1ZFU5BJ0U4lFXL4JXI7xS
zDy/wX6UyA7yyZmcAth/+KmujcTHtmxYLL9VBMoo1RiL4Agq0Sx0BbSAjZGV0tDN
lPRhcRWaS/1iAf5IGAU6ELPtm1tnXRhZemYk34eT+6OAWddHlq5WWHqg/9+TB0hl
tlhneTM3Ahw1oQYjfVCuyx8tbAB2Gl0GWReuy+KyXaVuxlevis5DA4PfgwKMj/+c
eL0AifVx55TXYd+Kwq1nZZShQ/K3uMhRYa2N/KGWbjeoLZqD76AsVKz1GXz2EcdH
bAUHvRvHZ6CKNLotmUwS0riHwHq0rTu4yVf9GWDN7DZahDhPXziq8zFr9LizAa8z
3FE+mmtpktAE5ckbrU8n7K1MrLINAUI4v/uHJbOMQ5XU6acH08kRCvIuDVFx9VxV
BNi8xmyR1cp7+ucEgl8M7RWRPI4cqKssQbXTp+jXFlOBaKm+yIrEL9gqpQFwyEvS
9sAxm2A0gBJtUF0YAmYzRwegtWd4Za6kx0OFo5Wr0MJ2ws/+R5MRihpC9bQb7CYk
BkkwXuNVyB1/aCYimBrECAmrfyeo3T6Ieb8szZ/JHQRTnEvWtwdC872Mqgp0Kr5H
Y6fscqsvyVp3JkBhVGOdjnWGXGux8+f/0n3hqO/8u2ZQyFPdT1oJRNrqXhaUgk+T
hZ9r9rNQ6nMgx8sNnNyUmln2CK3Pf+vHdc5tuTcJnhToW0K74Mn9GJ62gC/l8tSu
C0BTT2tBvuC/JSebZ7f5rH9WaboAF/R6/fnvu6hA/f5DKiste3zReaslvCYRU8po
v7sVoySYDM/dBUHJyMiNn/O6Uzui9c6q5ZpoVhQjFzCjaKFt+esyjTRxlQYFq0BX
6NqsJs/9WS2sLxFkkyZRJHvp7HshUjdiNFgWUbHjRbq8qiZP7GbX6TG+a9Ng0Nd8
9wTaYT2AZbzjuSJzBSgq0+QbrE2HJW0dtwzWt1CjYuOZpwarr8JXvlyuZk/BoyIC
mKDgSSpoKQT6oLYUae+pkR++aBoQJIhi411CfUxjctHIBKQq9kLk2drOJPzQb34J
d7sRV/9HlaHlaHXUHuQ0ZY+CphWIuoyz8FMKfljm5FKZariiw4FmhuttD9KNeusK
72qkuE+aWRzhOMUXAwWaxLzb0qYaJI9IFmu+W17dKVonQyqErMpXk+xOeitr8b6y
7gDDIlODFDPdjKKGFCTpvI0Agr2ypNKH+a49DPuG8Iwm+MoVgDESjt62M+GfOiiD
BLNbcvBbVZxS+trNhv46FhBe1/EOOn/ak1OoUgVKfQDio9LdhZ38Em1C2+0SuqTA
5C61xfclRJjXPm3697Ndc1veMSv6B52CY+udmBHKSzHJB/4gwf8s4J2AkSTiXbKG
f6uvHolSZoPMlzS432OIMNVoI++PoyjVQPYoQ3Sm9Nj4X5BWdMS5qbbXy2eLZYBo
jgEoV6kKlqboL7cOSCspqk5Hi0R/sh68mkqAqzzE3HOopUI1Zz5W5p/NGS0Tcsxu
IUX1t1F9MEgANd2PIh1vCAWYWMgjuSHZSnWpE6N2zL5QowEsaO40kzw/HRMDRMZL
KyDxldcgsaeTtsidLsBhYfCuOQVM/6ZHODqqInu9/hjZkCP5Iy8mHkCxWRqZgXMr
Mj5JTDiIj55vYiAyS1m7kOW8KZXYBgNBK4uedhdfMBrL3U1v/Tyv+uLciLUl1ILe
VH6A9vJT8bx5v154uVTZUG+APYsdTFWEXgviMyHofB7v+27/PG62bLnnyXJO7SJS
LnpUM+fv+/Y646RkqmRsNjBC3lK288BRe++s5S83M446PEWvU/ZZSatGnhXaRP06
oXLS56DW6BUtRRIDGDxuyaY8L5baOVEfB2jC2xGGep2rMT6Xp0FWzpmU+I4uDgKx
fuAS2AGaB+a0zxzg75u+IpvOh+qbNQ/2xcV0TcLehMh/WVZ/4rgmhyU+VZ8MKfUl
c0Q8dgqL3fLnHEj8e2oheyQ59wtE73wLkunOWSngEMB6YCJ+KtIHSVoroHvUd5w4
64/8Wl7t1fiDqXbq9XWl+JfNn698zsBNRHLvT+AuN08x6kRXDuTxqzjiE+4wRaFa
2HJ+ZqQIVQVrQK/mSdt2696Ua85AqQIX9fxV4L2wRvI/XB4krtoVVjxT6w61EyYb
08SqayhZhgxIzFS/XsngQv83hDPX6ocWO9VbUKJfHUmPsaCHffE6aYiIPZuGMZfL
UqjyO9QOwVvorlkMiile3BHEsgMuKD/2ijrUPO0br8r6WrGMYzDz+Gpp66t0TbDd
fFJKSZ/nkiE/C17nHTMYov5wPQ2bJAdXQAXk6EgurskNdAGSEZgdoCAMKyg7oVcE
MDe4U6uxEc3Wqzi7UoZlEOWiMdQf/rbcn10vyf2G6BM2yuHa/vk+fOM+lmelJOtX
b4A1iwtn/C0zXdbnzAsk3+ddZSXEboTc1+lbBfPlYa0NLz+ub98eY4rZmXKj2yUM
ySJeSsrn1xix+sbYfyL7g22QlU7y4LXqu+nOM0yInfFKaXbejoEKQLVdqX8JM77Y
xGOa6OHOS8rrDhON2yjz+8A09Kw6FGmapBpO0h8EUqyEFN68ubhaiyZ1dvlHjemi
F/k85ITUHyz5q88vKXdmfIyVBIgnuKSuk6vyGH1Yvpk/MuQe7VgDDiaZ2RdkIRVY
c29fzSq8JMNg9jrU4lz+9GlBK7TxG9lgoZAVTfkqGJDfNixvnonLROxr2le05vSf
ZQ2oIPwusPUIcJwoJqfEvuhPitEog3nbvSyNy8TRpJtuvKhPhfBpttZUDxDonz16
26TtoPZr/K4dopqctMsi1UgvsoAXL4tESlUYMcr02t+SEDxgwor6K9QpIAEJApkE
iTXiSdJXYArHasbURKILNd+qKJYMQvmibaBzJrGBDuVP3j55s8VcjutphQJYQi33
O44uva7elSI9esxEj2Vz0YsgSTHfrCfMEGcUcj7yhJGSmJEgPZJQJdbnrj3/WH/6
CzhqIscvU/nSl5Sa9TzrxZliBg+uQ6lQr+zUeFdGFEDJ54pk8IY+eOQCVirKo1rz
BGaMiFzPgDOW4Ux/uHqHLR7GHT3koHi/PN+vMuvynrjxsJ4tcklNty9d9LkuILiz
bYLlHLIfcSTtywGwHUQXly0oXjTKzGHkF8wgCyyrSwr/dyA+I8+ckljRMJwe+2La
Ocr7T1Rs4Siq8Ub7hrssPSMhdkGva26CivyDnPJJOJcKl7oW0YotEtGXchgLNBMw
/5nY8ZW4evumTmE3hQFuDkk3NuoXbgKTWv7QDaC8amu75YzNhABt3S4eUq1hsveK
NR0ilpENcUlT3dWHzHp4hBkcyIG1BB3sh0+a7wVJE5KB23YgM0Ktj4+27m3R6CuE
ETGmOag7tTcx1Devl/kmOwDn8HWPkMwi5uef1KT05v/KFoFg+4J+FlIuUIHlRS2S
TJEiEPrKqQPqgE3by4Mu+9tjnqWCEpM5P5/DJgWzt/idBsDk4LeE2aM+9A5UxpKh
ztxP0xwnDvyvBH7E4FXKUQFOTdXecmzRXybPf53XdiwtvHtSzh1DxUn3+Cyqjr+G
+SoZMa6OigBdnzfjEjfkaE+T/wS5mBWHhE/Onh9DKtyrzaBfdROhGC/bNDRQ8sAe
R+0rEV8UllCENz/sI69C7v8cMkknVt2OIDA710JO1xBjQZH4J6GRJx6ZZ6SXvDjc
PWIp7O2Ia7oG8FRKWgDPYMDMdX054x7PRf2VkqF1wOZk/Khm8/+FZR4fJ/0988Tb
56cKMowEqzxoH0Gc5pG6G49QexXJgZLKM+Xjb0OOyy70i/zvO9HjCn520B3wIPcW
xUyWtsCBJ/pzwyetHAfEKlUnv2hx/NyHSEQVcpu05w+2UULv20kR5c38qjcwheLL
9A2Kgkf8l+eUKVzBpZMmNdb8JTZZ0XczfQnDwLjQPMQSYfZZ/1dka8ll/YC9Z2/X
IUn7axQSB8ee+thdNgr46UfJn5HFTXEt5BpS0ObHlPn0hrOdTCPNkKAWNtBuwWZB
KmOGizsHP6Gz8WoqAAfhFjIM9nQhB7upfpwXIiAgqtc0RPTX1ybGzK8/fRftEL80
OlOs9E4sO9Lxw2t+8YxlBP2MJy5KrDbG1DJL/PzPgV50omi7aOaRuyrF/gLW+IoS
YIfhQXKSMS4GCbgx2KD74OXZmy3pSN9Zo4s0wlEoKiljFSv/vXIa99tGJ5tHnp8v
MIS78I3I+L2sXX0o8HvNlV6e0Dsfpxp2YT9lj7eXaN5KulxSwvMLj7oBOiM8Qxp7
`pragma protect end_protected
