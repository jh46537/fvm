// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: Status_Mux.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.0 Build 162 10/23/2013 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module Status_Mux (
	clock,
	data0x,
	data100x,
	data101x,
	data102x,
	data103x,
	data104x,
	data105x,
	data106x,
	data107x,
	data108x,
	data109x,
	data10x,
	data110x,
	data111x,
	data112x,
	data113x,
	data114x,
	data115x,
	data116x,
	data117x,
	data118x,
	data119x,
	data11x,
	data120x,
	data121x,
	data122x,
	data123x,
	data124x,
	data125x,
	data126x,
	data127x,
	data12x,
	data13x,
	data14x,
	data15x,
	data16x,
	data17x,
	data18x,
	data19x,
	data1x,
	data20x,
	data21x,
	data22x,
	data23x,
	data24x,
	data25x,
	data26x,
	data27x,
	data28x,
	data29x,
	data2x,
	data30x,
	data31x,
	data32x,
	data33x,
	data34x,
	data35x,
	data36x,
	data37x,
	data38x,
	data39x,
	data3x,
	data40x,
	data41x,
	data42x,
	data43x,
	data44x,
	data45x,
	data46x,
	data47x,
	data48x,
	data49x,
	data4x,
	data50x,
	data51x,
	data52x,
	data53x,
	data54x,
	data55x,
	data56x,
	data57x,
	data58x,
	data59x,
	data5x,
	data60x,
	data61x,
	data62x,
	data63x,
	data64x,
	data65x,
	data66x,
	data67x,
	data68x,
	data69x,
	data6x,
	data70x,
	data71x,
	data72x,
	data73x,
	data74x,
	data75x,
	data76x,
	data77x,
	data78x,
	data79x,
	data7x,
	data80x,
	data81x,
	data82x,
	data83x,
	data84x,
	data85x,
	data86x,
	data87x,
	data88x,
	data89x,
	data8x,
	data90x,
	data91x,
	data92x,
	data93x,
	data94x,
	data95x,
	data96x,
	data97x,
	data98x,
	data99x,
	data9x,
	sel,
	result);

	input	  clock;
	input	[31:0]  data0x;
	input	[31:0]  data100x;
	input	[31:0]  data101x;
	input	[31:0]  data102x;
	input	[31:0]  data103x;
	input	[31:0]  data104x;
	input	[31:0]  data105x;
	input	[31:0]  data106x;
	input	[31:0]  data107x;
	input	[31:0]  data108x;
	input	[31:0]  data109x;
	input	[31:0]  data10x;
	input	[31:0]  data110x;
	input	[31:0]  data111x;
	input	[31:0]  data112x;
	input	[31:0]  data113x;
	input	[31:0]  data114x;
	input	[31:0]  data115x;
	input	[31:0]  data116x;
	input	[31:0]  data117x;
	input	[31:0]  data118x;
	input	[31:0]  data119x;
	input	[31:0]  data11x;
	input	[31:0]  data120x;
	input	[31:0]  data121x;
	input	[31:0]  data122x;
	input	[31:0]  data123x;
	input	[31:0]  data124x;
	input	[31:0]  data125x;
	input	[31:0]  data126x;
	input	[31:0]  data127x;
	input	[31:0]  data12x;
	input	[31:0]  data13x;
	input	[31:0]  data14x;
	input	[31:0]  data15x;
	input	[31:0]  data16x;
	input	[31:0]  data17x;
	input	[31:0]  data18x;
	input	[31:0]  data19x;
	input	[31:0]  data1x;
	input	[31:0]  data20x;
	input	[31:0]  data21x;
	input	[31:0]  data22x;
	input	[31:0]  data23x;
	input	[31:0]  data24x;
	input	[31:0]  data25x;
	input	[31:0]  data26x;
	input	[31:0]  data27x;
	input	[31:0]  data28x;
	input	[31:0]  data29x;
	input	[31:0]  data2x;
	input	[31:0]  data30x;
	input	[31:0]  data31x;
	input	[31:0]  data32x;
	input	[31:0]  data33x;
	input	[31:0]  data34x;
	input	[31:0]  data35x;
	input	[31:0]  data36x;
	input	[31:0]  data37x;
	input	[31:0]  data38x;
	input	[31:0]  data39x;
	input	[31:0]  data3x;
	input	[31:0]  data40x;
	input	[31:0]  data41x;
	input	[31:0]  data42x;
	input	[31:0]  data43x;
	input	[31:0]  data44x;
	input	[31:0]  data45x;
	input	[31:0]  data46x;
	input	[31:0]  data47x;
	input	[31:0]  data48x;
	input	[31:0]  data49x;
	input	[31:0]  data4x;
	input	[31:0]  data50x;
	input	[31:0]  data51x;
	input	[31:0]  data52x;
	input	[31:0]  data53x;
	input	[31:0]  data54x;
	input	[31:0]  data55x;
	input	[31:0]  data56x;
	input	[31:0]  data57x;
	input	[31:0]  data58x;
	input	[31:0]  data59x;
	input	[31:0]  data5x;
	input	[31:0]  data60x;
	input	[31:0]  data61x;
	input	[31:0]  data62x;
	input	[31:0]  data63x;
	input	[31:0]  data64x;
	input	[31:0]  data65x;
	input	[31:0]  data66x;
	input	[31:0]  data67x;
	input	[31:0]  data68x;
	input	[31:0]  data69x;
	input	[31:0]  data6x;
	input	[31:0]  data70x;
	input	[31:0]  data71x;
	input	[31:0]  data72x;
	input	[31:0]  data73x;
	input	[31:0]  data74x;
	input	[31:0]  data75x;
	input	[31:0]  data76x;
	input	[31:0]  data77x;
	input	[31:0]  data78x;
	input	[31:0]  data79x;
	input	[31:0]  data7x;
	input	[31:0]  data80x;
	input	[31:0]  data81x;
	input	[31:0]  data82x;
	input	[31:0]  data83x;
	input	[31:0]  data84x;
	input	[31:0]  data85x;
	input	[31:0]  data86x;
	input	[31:0]  data87x;
	input	[31:0]  data88x;
	input	[31:0]  data89x;
	input	[31:0]  data8x;
	input	[31:0]  data90x;
	input	[31:0]  data91x;
	input	[31:0]  data92x;
	input	[31:0]  data93x;
	input	[31:0]  data94x;
	input	[31:0]  data95x;
	input	[31:0]  data96x;
	input	[31:0]  data97x;
	input	[31:0]  data98x;
	input	[31:0]  data99x;
	input	[31:0]  data9x;
	input	[6:0]  sel;
	output	[31:0]  result;

	wire [31:0] sub_wire0;
	wire [31:0] sub_wire129 = data127x[31:0];
	wire [31:0] sub_wire128 = data126x[31:0];
	wire [31:0] sub_wire127 = data125x[31:0];
	wire [31:0] sub_wire126 = data124x[31:0];
	wire [31:0] sub_wire125 = data123x[31:0];
	wire [31:0] sub_wire124 = data122x[31:0];
	wire [31:0] sub_wire123 = data121x[31:0];
	wire [31:0] sub_wire122 = data120x[31:0];
	wire [31:0] sub_wire121 = data119x[31:0];
	wire [31:0] sub_wire120 = data118x[31:0];
	wire [31:0] sub_wire119 = data117x[31:0];
	wire [31:0] sub_wire118 = data116x[31:0];
	wire [31:0] sub_wire117 = data115x[31:0];
	wire [31:0] sub_wire116 = data114x[31:0];
	wire [31:0] sub_wire115 = data113x[31:0];
	wire [31:0] sub_wire114 = data112x[31:0];
	wire [31:0] sub_wire113 = data111x[31:0];
	wire [31:0] sub_wire112 = data110x[31:0];
	wire [31:0] sub_wire111 = data109x[31:0];
	wire [31:0] sub_wire110 = data108x[31:0];
	wire [31:0] sub_wire109 = data107x[31:0];
	wire [31:0] sub_wire108 = data106x[31:0];
	wire [31:0] sub_wire107 = data105x[31:0];
	wire [31:0] sub_wire106 = data104x[31:0];
	wire [31:0] sub_wire105 = data103x[31:0];
	wire [31:0] sub_wire104 = data102x[31:0];
	wire [31:0] sub_wire103 = data101x[31:0];
	wire [31:0] sub_wire102 = data100x[31:0];
	wire [31:0] sub_wire101 = data99x[31:0];
	wire [31:0] sub_wire100 = data98x[31:0];
	wire [31:0] sub_wire99 = data97x[31:0];
	wire [31:0] sub_wire98 = data96x[31:0];
	wire [31:0] sub_wire97 = data95x[31:0];
	wire [31:0] sub_wire96 = data94x[31:0];
	wire [31:0] sub_wire95 = data93x[31:0];
	wire [31:0] sub_wire94 = data92x[31:0];
	wire [31:0] sub_wire93 = data91x[31:0];
	wire [31:0] sub_wire92 = data90x[31:0];
	wire [31:0] sub_wire91 = data89x[31:0];
	wire [31:0] sub_wire90 = data88x[31:0];
	wire [31:0] sub_wire89 = data87x[31:0];
	wire [31:0] sub_wire88 = data86x[31:0];
	wire [31:0] sub_wire87 = data85x[31:0];
	wire [31:0] sub_wire86 = data84x[31:0];
	wire [31:0] sub_wire85 = data83x[31:0];
	wire [31:0] sub_wire84 = data82x[31:0];
	wire [31:0] sub_wire83 = data81x[31:0];
	wire [31:0] sub_wire82 = data80x[31:0];
	wire [31:0] sub_wire81 = data79x[31:0];
	wire [31:0] sub_wire80 = data78x[31:0];
	wire [31:0] sub_wire79 = data77x[31:0];
	wire [31:0] sub_wire78 = data76x[31:0];
	wire [31:0] sub_wire77 = data75x[31:0];
	wire [31:0] sub_wire76 = data74x[31:0];
	wire [31:0] sub_wire75 = data73x[31:0];
	wire [31:0] sub_wire74 = data72x[31:0];
	wire [31:0] sub_wire73 = data71x[31:0];
	wire [31:0] sub_wire72 = data70x[31:0];
	wire [31:0] sub_wire71 = data69x[31:0];
	wire [31:0] sub_wire70 = data68x[31:0];
	wire [31:0] sub_wire69 = data67x[31:0];
	wire [31:0] sub_wire68 = data66x[31:0];
	wire [31:0] sub_wire67 = data65x[31:0];
	wire [31:0] sub_wire66 = data64x[31:0];
	wire [31:0] sub_wire65 = data63x[31:0];
	wire [31:0] sub_wire64 = data62x[31:0];
	wire [31:0] sub_wire63 = data61x[31:0];
	wire [31:0] sub_wire62 = data60x[31:0];
	wire [31:0] sub_wire61 = data59x[31:0];
	wire [31:0] sub_wire60 = data58x[31:0];
	wire [31:0] sub_wire59 = data57x[31:0];
	wire [31:0] sub_wire58 = data56x[31:0];
	wire [31:0] sub_wire57 = data55x[31:0];
	wire [31:0] sub_wire56 = data54x[31:0];
	wire [31:0] sub_wire55 = data53x[31:0];
	wire [31:0] sub_wire54 = data52x[31:0];
	wire [31:0] sub_wire53 = data51x[31:0];
	wire [31:0] sub_wire52 = data50x[31:0];
	wire [31:0] sub_wire51 = data49x[31:0];
	wire [31:0] sub_wire50 = data48x[31:0];
	wire [31:0] sub_wire49 = data47x[31:0];
	wire [31:0] sub_wire48 = data46x[31:0];
	wire [31:0] sub_wire47 = data45x[31:0];
	wire [31:0] sub_wire46 = data44x[31:0];
	wire [31:0] sub_wire45 = data43x[31:0];
	wire [31:0] sub_wire44 = data42x[31:0];
	wire [31:0] sub_wire43 = data41x[31:0];
	wire [31:0] sub_wire42 = data40x[31:0];
	wire [31:0] sub_wire41 = data39x[31:0];
	wire [31:0] sub_wire40 = data38x[31:0];
	wire [31:0] sub_wire39 = data37x[31:0];
	wire [31:0] sub_wire38 = data36x[31:0];
	wire [31:0] sub_wire37 = data35x[31:0];
	wire [31:0] sub_wire36 = data34x[31:0];
	wire [31:0] sub_wire35 = data33x[31:0];
	wire [31:0] sub_wire34 = data32x[31:0];
	wire [31:0] sub_wire33 = data31x[31:0];
	wire [31:0] sub_wire32 = data30x[31:0];
	wire [31:0] sub_wire31 = data29x[31:0];
	wire [31:0] sub_wire30 = data28x[31:0];
	wire [31:0] sub_wire29 = data27x[31:0];
	wire [31:0] sub_wire28 = data26x[31:0];
	wire [31:0] sub_wire27 = data25x[31:0];
	wire [31:0] sub_wire26 = data24x[31:0];
	wire [31:0] sub_wire25 = data23x[31:0];
	wire [31:0] sub_wire24 = data22x[31:0];
	wire [31:0] sub_wire23 = data21x[31:0];
	wire [31:0] sub_wire22 = data20x[31:0];
	wire [31:0] sub_wire21 = data19x[31:0];
	wire [31:0] sub_wire20 = data18x[31:0];
	wire [31:0] sub_wire19 = data17x[31:0];
	wire [31:0] sub_wire18 = data16x[31:0];
	wire [31:0] sub_wire17 = data15x[31:0];
	wire [31:0] sub_wire16 = data14x[31:0];
	wire [31:0] sub_wire15 = data13x[31:0];
	wire [31:0] sub_wire14 = data12x[31:0];
	wire [31:0] sub_wire13 = data11x[31:0];
	wire [31:0] sub_wire12 = data10x[31:0];
	wire [31:0] sub_wire11 = data9x[31:0];
	wire [31:0] sub_wire10 = data8x[31:0];
	wire [31:0] sub_wire9 = data7x[31:0];
	wire [31:0] sub_wire8 = data6x[31:0];
	wire [31:0] sub_wire7 = data5x[31:0];
	wire [31:0] sub_wire6 = data4x[31:0];
	wire [31:0] sub_wire5 = data3x[31:0];
	wire [31:0] sub_wire4 = data2x[31:0];
	wire [31:0] sub_wire3 = data1x[31:0];
	wire [31:0] result = sub_wire0[31:0];
	wire [31:0] sub_wire1 = data0x[31:0];
	wire [4095:0] sub_wire2 = {sub_wire129, sub_wire128, sub_wire127, sub_wire126, sub_wire125, sub_wire124, sub_wire123, sub_wire122, sub_wire121, sub_wire120, sub_wire119, sub_wire118, sub_wire117, sub_wire116, sub_wire115, sub_wire114, sub_wire113, sub_wire112, sub_wire111, sub_wire110, sub_wire109, sub_wire108, sub_wire107, sub_wire106, sub_wire105, sub_wire104, sub_wire103, sub_wire102, sub_wire101, sub_wire100, sub_wire99, sub_wire98, sub_wire97, sub_wire96, sub_wire95, sub_wire94, sub_wire93, sub_wire92, sub_wire91, sub_wire90, sub_wire89, sub_wire88, sub_wire87, sub_wire86, sub_wire85, sub_wire84, sub_wire83, sub_wire82, sub_wire81, sub_wire80, sub_wire79, sub_wire78, sub_wire77, sub_wire76, sub_wire75, sub_wire74, sub_wire73, sub_wire72, sub_wire71, sub_wire70, sub_wire69, sub_wire68, sub_wire67, sub_wire66, sub_wire65, sub_wire64, sub_wire63, sub_wire62, sub_wire61, sub_wire60, sub_wire59, sub_wire58, sub_wire57, sub_wire56, sub_wire55, sub_wire54, sub_wire53, sub_wire52, sub_wire51, sub_wire50, sub_wire49, sub_wire48, sub_wire47, sub_wire46, sub_wire45, sub_wire44, sub_wire43, sub_wire42, sub_wire41, sub_wire40, sub_wire39, sub_wire38, sub_wire37, sub_wire36, sub_wire35, sub_wire34, sub_wire33, sub_wire32, sub_wire31, sub_wire30, sub_wire29, sub_wire28, sub_wire27, sub_wire26, sub_wire25, sub_wire24, sub_wire23, sub_wire22, sub_wire21, sub_wire20, sub_wire19, sub_wire18, sub_wire17, sub_wire16, sub_wire15, sub_wire14, sub_wire13, sub_wire12, sub_wire11, sub_wire10, sub_wire9, sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4, sub_wire3, sub_wire1};

	lpm_mux	LPM_MUX_component (
				.clock (clock),
				.data (sub_wire2),
				.sel (sel),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken ()
				// synopsys translate_on
				);
	defparam
		LPM_MUX_component.lpm_pipeline = 4,
		LPM_MUX_component.lpm_size = 128,
		LPM_MUX_component.lpm_type = "LPM_MUX",
		LPM_MUX_component.lpm_width = 32,
		LPM_MUX_component.lpm_widths = 7;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "4"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "128"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "32"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "7"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: data0x 0 0 32 0 INPUT NODEFVAL "data0x[31..0]"
// Retrieval info: USED_PORT: data100x 0 0 32 0 INPUT NODEFVAL "data100x[31..0]"
// Retrieval info: USED_PORT: data101x 0 0 32 0 INPUT NODEFVAL "data101x[31..0]"
// Retrieval info: USED_PORT: data102x 0 0 32 0 INPUT NODEFVAL "data102x[31..0]"
// Retrieval info: USED_PORT: data103x 0 0 32 0 INPUT NODEFVAL "data103x[31..0]"
// Retrieval info: USED_PORT: data104x 0 0 32 0 INPUT NODEFVAL "data104x[31..0]"
// Retrieval info: USED_PORT: data105x 0 0 32 0 INPUT NODEFVAL "data105x[31..0]"
// Retrieval info: USED_PORT: data106x 0 0 32 0 INPUT NODEFVAL "data106x[31..0]"
// Retrieval info: USED_PORT: data107x 0 0 32 0 INPUT NODEFVAL "data107x[31..0]"
// Retrieval info: USED_PORT: data108x 0 0 32 0 INPUT NODEFVAL "data108x[31..0]"
// Retrieval info: USED_PORT: data109x 0 0 32 0 INPUT NODEFVAL "data109x[31..0]"
// Retrieval info: USED_PORT: data10x 0 0 32 0 INPUT NODEFVAL "data10x[31..0]"
// Retrieval info: USED_PORT: data110x 0 0 32 0 INPUT NODEFVAL "data110x[31..0]"
// Retrieval info: USED_PORT: data111x 0 0 32 0 INPUT NODEFVAL "data111x[31..0]"
// Retrieval info: USED_PORT: data112x 0 0 32 0 INPUT NODEFVAL "data112x[31..0]"
// Retrieval info: USED_PORT: data113x 0 0 32 0 INPUT NODEFVAL "data113x[31..0]"
// Retrieval info: USED_PORT: data114x 0 0 32 0 INPUT NODEFVAL "data114x[31..0]"
// Retrieval info: USED_PORT: data115x 0 0 32 0 INPUT NODEFVAL "data115x[31..0]"
// Retrieval info: USED_PORT: data116x 0 0 32 0 INPUT NODEFVAL "data116x[31..0]"
// Retrieval info: USED_PORT: data117x 0 0 32 0 INPUT NODEFVAL "data117x[31..0]"
// Retrieval info: USED_PORT: data118x 0 0 32 0 INPUT NODEFVAL "data118x[31..0]"
// Retrieval info: USED_PORT: data119x 0 0 32 0 INPUT NODEFVAL "data119x[31..0]"
// Retrieval info: USED_PORT: data11x 0 0 32 0 INPUT NODEFVAL "data11x[31..0]"
// Retrieval info: USED_PORT: data120x 0 0 32 0 INPUT NODEFVAL "data120x[31..0]"
// Retrieval info: USED_PORT: data121x 0 0 32 0 INPUT NODEFVAL "data121x[31..0]"
// Retrieval info: USED_PORT: data122x 0 0 32 0 INPUT NODEFVAL "data122x[31..0]"
// Retrieval info: USED_PORT: data123x 0 0 32 0 INPUT NODEFVAL "data123x[31..0]"
// Retrieval info: USED_PORT: data124x 0 0 32 0 INPUT NODEFVAL "data124x[31..0]"
// Retrieval info: USED_PORT: data125x 0 0 32 0 INPUT NODEFVAL "data125x[31..0]"
// Retrieval info: USED_PORT: data126x 0 0 32 0 INPUT NODEFVAL "data126x[31..0]"
// Retrieval info: USED_PORT: data127x 0 0 32 0 INPUT NODEFVAL "data127x[31..0]"
// Retrieval info: USED_PORT: data12x 0 0 32 0 INPUT NODEFVAL "data12x[31..0]"
// Retrieval info: USED_PORT: data13x 0 0 32 0 INPUT NODEFVAL "data13x[31..0]"
// Retrieval info: USED_PORT: data14x 0 0 32 0 INPUT NODEFVAL "data14x[31..0]"
// Retrieval info: USED_PORT: data15x 0 0 32 0 INPUT NODEFVAL "data15x[31..0]"
// Retrieval info: USED_PORT: data16x 0 0 32 0 INPUT NODEFVAL "data16x[31..0]"
// Retrieval info: USED_PORT: data17x 0 0 32 0 INPUT NODEFVAL "data17x[31..0]"
// Retrieval info: USED_PORT: data18x 0 0 32 0 INPUT NODEFVAL "data18x[31..0]"
// Retrieval info: USED_PORT: data19x 0 0 32 0 INPUT NODEFVAL "data19x[31..0]"
// Retrieval info: USED_PORT: data1x 0 0 32 0 INPUT NODEFVAL "data1x[31..0]"
// Retrieval info: USED_PORT: data20x 0 0 32 0 INPUT NODEFVAL "data20x[31..0]"
// Retrieval info: USED_PORT: data21x 0 0 32 0 INPUT NODEFVAL "data21x[31..0]"
// Retrieval info: USED_PORT: data22x 0 0 32 0 INPUT NODEFVAL "data22x[31..0]"
// Retrieval info: USED_PORT: data23x 0 0 32 0 INPUT NODEFVAL "data23x[31..0]"
// Retrieval info: USED_PORT: data24x 0 0 32 0 INPUT NODEFVAL "data24x[31..0]"
// Retrieval info: USED_PORT: data25x 0 0 32 0 INPUT NODEFVAL "data25x[31..0]"
// Retrieval info: USED_PORT: data26x 0 0 32 0 INPUT NODEFVAL "data26x[31..0]"
// Retrieval info: USED_PORT: data27x 0 0 32 0 INPUT NODEFVAL "data27x[31..0]"
// Retrieval info: USED_PORT: data28x 0 0 32 0 INPUT NODEFVAL "data28x[31..0]"
// Retrieval info: USED_PORT: data29x 0 0 32 0 INPUT NODEFVAL "data29x[31..0]"
// Retrieval info: USED_PORT: data2x 0 0 32 0 INPUT NODEFVAL "data2x[31..0]"
// Retrieval info: USED_PORT: data30x 0 0 32 0 INPUT NODEFVAL "data30x[31..0]"
// Retrieval info: USED_PORT: data31x 0 0 32 0 INPUT NODEFVAL "data31x[31..0]"
// Retrieval info: USED_PORT: data32x 0 0 32 0 INPUT NODEFVAL "data32x[31..0]"
// Retrieval info: USED_PORT: data33x 0 0 32 0 INPUT NODEFVAL "data33x[31..0]"
// Retrieval info: USED_PORT: data34x 0 0 32 0 INPUT NODEFVAL "data34x[31..0]"
// Retrieval info: USED_PORT: data35x 0 0 32 0 INPUT NODEFVAL "data35x[31..0]"
// Retrieval info: USED_PORT: data36x 0 0 32 0 INPUT NODEFVAL "data36x[31..0]"
// Retrieval info: USED_PORT: data37x 0 0 32 0 INPUT NODEFVAL "data37x[31..0]"
// Retrieval info: USED_PORT: data38x 0 0 32 0 INPUT NODEFVAL "data38x[31..0]"
// Retrieval info: USED_PORT: data39x 0 0 32 0 INPUT NODEFVAL "data39x[31..0]"
// Retrieval info: USED_PORT: data3x 0 0 32 0 INPUT NODEFVAL "data3x[31..0]"
// Retrieval info: USED_PORT: data40x 0 0 32 0 INPUT NODEFVAL "data40x[31..0]"
// Retrieval info: USED_PORT: data41x 0 0 32 0 INPUT NODEFVAL "data41x[31..0]"
// Retrieval info: USED_PORT: data42x 0 0 32 0 INPUT NODEFVAL "data42x[31..0]"
// Retrieval info: USED_PORT: data43x 0 0 32 0 INPUT NODEFVAL "data43x[31..0]"
// Retrieval info: USED_PORT: data44x 0 0 32 0 INPUT NODEFVAL "data44x[31..0]"
// Retrieval info: USED_PORT: data45x 0 0 32 0 INPUT NODEFVAL "data45x[31..0]"
// Retrieval info: USED_PORT: data46x 0 0 32 0 INPUT NODEFVAL "data46x[31..0]"
// Retrieval info: USED_PORT: data47x 0 0 32 0 INPUT NODEFVAL "data47x[31..0]"
// Retrieval info: USED_PORT: data48x 0 0 32 0 INPUT NODEFVAL "data48x[31..0]"
// Retrieval info: USED_PORT: data49x 0 0 32 0 INPUT NODEFVAL "data49x[31..0]"
// Retrieval info: USED_PORT: data4x 0 0 32 0 INPUT NODEFVAL "data4x[31..0]"
// Retrieval info: USED_PORT: data50x 0 0 32 0 INPUT NODEFVAL "data50x[31..0]"
// Retrieval info: USED_PORT: data51x 0 0 32 0 INPUT NODEFVAL "data51x[31..0]"
// Retrieval info: USED_PORT: data52x 0 0 32 0 INPUT NODEFVAL "data52x[31..0]"
// Retrieval info: USED_PORT: data53x 0 0 32 0 INPUT NODEFVAL "data53x[31..0]"
// Retrieval info: USED_PORT: data54x 0 0 32 0 INPUT NODEFVAL "data54x[31..0]"
// Retrieval info: USED_PORT: data55x 0 0 32 0 INPUT NODEFVAL "data55x[31..0]"
// Retrieval info: USED_PORT: data56x 0 0 32 0 INPUT NODEFVAL "data56x[31..0]"
// Retrieval info: USED_PORT: data57x 0 0 32 0 INPUT NODEFVAL "data57x[31..0]"
// Retrieval info: USED_PORT: data58x 0 0 32 0 INPUT NODEFVAL "data58x[31..0]"
// Retrieval info: USED_PORT: data59x 0 0 32 0 INPUT NODEFVAL "data59x[31..0]"
// Retrieval info: USED_PORT: data5x 0 0 32 0 INPUT NODEFVAL "data5x[31..0]"
// Retrieval info: USED_PORT: data60x 0 0 32 0 INPUT NODEFVAL "data60x[31..0]"
// Retrieval info: USED_PORT: data61x 0 0 32 0 INPUT NODEFVAL "data61x[31..0]"
// Retrieval info: USED_PORT: data62x 0 0 32 0 INPUT NODEFVAL "data62x[31..0]"
// Retrieval info: USED_PORT: data63x 0 0 32 0 INPUT NODEFVAL "data63x[31..0]"
// Retrieval info: USED_PORT: data64x 0 0 32 0 INPUT NODEFVAL "data64x[31..0]"
// Retrieval info: USED_PORT: data65x 0 0 32 0 INPUT NODEFVAL "data65x[31..0]"
// Retrieval info: USED_PORT: data66x 0 0 32 0 INPUT NODEFVAL "data66x[31..0]"
// Retrieval info: USED_PORT: data67x 0 0 32 0 INPUT NODEFVAL "data67x[31..0]"
// Retrieval info: USED_PORT: data68x 0 0 32 0 INPUT NODEFVAL "data68x[31..0]"
// Retrieval info: USED_PORT: data69x 0 0 32 0 INPUT NODEFVAL "data69x[31..0]"
// Retrieval info: USED_PORT: data6x 0 0 32 0 INPUT NODEFVAL "data6x[31..0]"
// Retrieval info: USED_PORT: data70x 0 0 32 0 INPUT NODEFVAL "data70x[31..0]"
// Retrieval info: USED_PORT: data71x 0 0 32 0 INPUT NODEFVAL "data71x[31..0]"
// Retrieval info: USED_PORT: data72x 0 0 32 0 INPUT NODEFVAL "data72x[31..0]"
// Retrieval info: USED_PORT: data73x 0 0 32 0 INPUT NODEFVAL "data73x[31..0]"
// Retrieval info: USED_PORT: data74x 0 0 32 0 INPUT NODEFVAL "data74x[31..0]"
// Retrieval info: USED_PORT: data75x 0 0 32 0 INPUT NODEFVAL "data75x[31..0]"
// Retrieval info: USED_PORT: data76x 0 0 32 0 INPUT NODEFVAL "data76x[31..0]"
// Retrieval info: USED_PORT: data77x 0 0 32 0 INPUT NODEFVAL "data77x[31..0]"
// Retrieval info: USED_PORT: data78x 0 0 32 0 INPUT NODEFVAL "data78x[31..0]"
// Retrieval info: USED_PORT: data79x 0 0 32 0 INPUT NODEFVAL "data79x[31..0]"
// Retrieval info: USED_PORT: data7x 0 0 32 0 INPUT NODEFVAL "data7x[31..0]"
// Retrieval info: USED_PORT: data80x 0 0 32 0 INPUT NODEFVAL "data80x[31..0]"
// Retrieval info: USED_PORT: data81x 0 0 32 0 INPUT NODEFVAL "data81x[31..0]"
// Retrieval info: USED_PORT: data82x 0 0 32 0 INPUT NODEFVAL "data82x[31..0]"
// Retrieval info: USED_PORT: data83x 0 0 32 0 INPUT NODEFVAL "data83x[31..0]"
// Retrieval info: USED_PORT: data84x 0 0 32 0 INPUT NODEFVAL "data84x[31..0]"
// Retrieval info: USED_PORT: data85x 0 0 32 0 INPUT NODEFVAL "data85x[31..0]"
// Retrieval info: USED_PORT: data86x 0 0 32 0 INPUT NODEFVAL "data86x[31..0]"
// Retrieval info: USED_PORT: data87x 0 0 32 0 INPUT NODEFVAL "data87x[31..0]"
// Retrieval info: USED_PORT: data88x 0 0 32 0 INPUT NODEFVAL "data88x[31..0]"
// Retrieval info: USED_PORT: data89x 0 0 32 0 INPUT NODEFVAL "data89x[31..0]"
// Retrieval info: USED_PORT: data8x 0 0 32 0 INPUT NODEFVAL "data8x[31..0]"
// Retrieval info: USED_PORT: data90x 0 0 32 0 INPUT NODEFVAL "data90x[31..0]"
// Retrieval info: USED_PORT: data91x 0 0 32 0 INPUT NODEFVAL "data91x[31..0]"
// Retrieval info: USED_PORT: data92x 0 0 32 0 INPUT NODEFVAL "data92x[31..0]"
// Retrieval info: USED_PORT: data93x 0 0 32 0 INPUT NODEFVAL "data93x[31..0]"
// Retrieval info: USED_PORT: data94x 0 0 32 0 INPUT NODEFVAL "data94x[31..0]"
// Retrieval info: USED_PORT: data95x 0 0 32 0 INPUT NODEFVAL "data95x[31..0]"
// Retrieval info: USED_PORT: data96x 0 0 32 0 INPUT NODEFVAL "data96x[31..0]"
// Retrieval info: USED_PORT: data97x 0 0 32 0 INPUT NODEFVAL "data97x[31..0]"
// Retrieval info: USED_PORT: data98x 0 0 32 0 INPUT NODEFVAL "data98x[31..0]"
// Retrieval info: USED_PORT: data99x 0 0 32 0 INPUT NODEFVAL "data99x[31..0]"
// Retrieval info: USED_PORT: data9x 0 0 32 0 INPUT NODEFVAL "data9x[31..0]"
// Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
// Retrieval info: USED_PORT: sel 0 0 7 0 INPUT NODEFVAL "sel[6..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 32 0 data0x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3200 data100x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3232 data101x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3264 data102x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3296 data103x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3328 data104x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3360 data105x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3392 data106x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3424 data107x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3456 data108x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3488 data109x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 320 data10x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3520 data110x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3552 data111x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3584 data112x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3616 data113x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3648 data114x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3680 data115x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3712 data116x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3744 data117x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3776 data118x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3808 data119x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 352 data11x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3840 data120x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3872 data121x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3904 data122x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3936 data123x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3968 data124x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 4000 data125x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 4032 data126x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 4064 data127x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 384 data12x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 416 data13x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 448 data14x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 480 data15x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 512 data16x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 544 data17x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 576 data18x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 608 data19x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 32 data1x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 640 data20x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 672 data21x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 704 data22x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 736 data23x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 768 data24x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 800 data25x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 832 data26x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 864 data27x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 896 data28x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 928 data29x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 64 data2x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 960 data30x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 992 data31x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1024 data32x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1056 data33x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1088 data34x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1120 data35x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1152 data36x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1184 data37x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1216 data38x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1248 data39x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 96 data3x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1280 data40x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1312 data41x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1344 data42x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1376 data43x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1408 data44x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1440 data45x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1472 data46x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1504 data47x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1536 data48x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1568 data49x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 128 data4x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1600 data50x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1632 data51x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1664 data52x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1696 data53x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1728 data54x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1760 data55x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1792 data56x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1824 data57x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1856 data58x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1888 data59x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 160 data5x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1920 data60x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1952 data61x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 1984 data62x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2016 data63x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2048 data64x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2080 data65x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2112 data66x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2144 data67x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2176 data68x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2208 data69x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 192 data6x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2240 data70x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2272 data71x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2304 data72x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2336 data73x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2368 data74x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2400 data75x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2432 data76x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2464 data77x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2496 data78x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2528 data79x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 224 data7x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2560 data80x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2592 data81x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2624 data82x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2656 data83x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2688 data84x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2720 data85x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2752 data86x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2784 data87x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2816 data88x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2848 data89x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 256 data8x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2880 data90x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2912 data91x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2944 data92x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 2976 data93x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3008 data94x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3040 data95x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3072 data96x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3104 data97x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3136 data98x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 3168 data99x 0 0 32 0
// Retrieval info: CONNECT: @data 0 0 32 288 data9x 0 0 32 0
// Retrieval info: CONNECT: @sel 0 0 7 0 sel 0 0 7 0
// Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
// Retrieval info: GEN_FILE: TYPE_NORMAL Status_Mux.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Status_Mux.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Status_Mux.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Status_Mux.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Status_Mux_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Status_Mux_bb.v FALSE
// Retrieval info: LIB_FILE: lpm
