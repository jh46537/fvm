��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���� 6�:$���mQ�$��z��˙Y���A�.�.xn]H���H�2��* ������<�7=}�ȥ������O��l��ni��1�F8^]���c�"'�$�ԝu;B���L�t�y�G�J-�B��\�ȶ�y)�aL�3�T�f��"n��?W�\nzL3o�Y��f�9[�WWE)�S�c���ە�gQ�>��'�cu�Ā	�}4C�Kj�kk�
��b��s�>A4�M_���>�4*�e+��.�~
=�~w'E�y��a�}�5�b����"��"�m47�+�x.��8� �˜\l�	���tB��c�Z&�`]IS��p}hC���/**���Lg�.�0g��/���k�H�Đ�(�2�/��x G7��軬B��SZeL=��4kDq.�$N�*�(X��cv�X`��UhR���tg�Wx��3|��}�3�v����R�JLh��7��h@_����o����C��Ȳ�8��KĖ��o\>(��6����P�)�Os�`�і+[���<�6���UW@̍,��tU ��> u�KP-�:Э8���m:����/y�|����H3Gs�y40�8�t�����0��Gi�dAH���Z�ө#�&,q�F�v��<���J+�Z�Lƅ�jk����#����N
˃�5
D
̦Ƥ�B�%0�,����ݮ� # u��Pk���#
"y�js��;6$�Q��h���
#ڕg^�UJ���_-���AC����)"�H�EtN�q0��Ζ��ւȐp1��F1S�@��u�a��h��8G�BKYK�Bۮ+97	U���ᡉ�x���ˎq*(����ny�=��>�^Vb}����G����
vT1h:u�H]h��E��.�_ӴU@�nf��2 [��=.��.��^��?T��g�?��j��� 7����y�A@A/y9qJ�⺤�́a�mc��I���q��s(���w}��w;��*}�L3R��d_���Pi��)F�/�)c�d"~<]N֫�*�ꐦ��?� ��P��Y�N�Қ =^�1o�{l<��>�σʲ0��ho����QF1���b $H�9h���~Z`\���j�]�Fm>Y�0f-y��5���^z�Ym��=iu���FU�L��Q�v� V�6�O����v)�|K1o�P��b#�$�U�i$��� �jX�O���Ui3Ā�Y�EL�%7�WG��A�D鼔�O��l\LB�Y�O�?�D�ۭ�A�|����wǮ���>��M�ܗnƔˏ3O_vMMȿJȿ��>J ��x���
��6�F�;�-P.��,��V�ע�t�u�8��I>�"��͖>Ms���j��}�6��&����/>5�ĩ61B/���m��J3�R�k`g�+�o	4���A��\��%��&���aط���ʼ�HM������b�h^���Su��t��B.��[9�Ӣ�:Jzk�����]]a֫��/chIm�|n���v����b���"�qx&�8Fv��#��l��1�jp�3��|�:/-#'|��ɀ�P�P���X�"U�
��;s c"�J��t�({�|j����ܥ�`��U9;?|E0LF+_�� |��w�&U=L�G�__kb�:2^��>W�ǞK���]l�/(k��r��fs�<�,�᪕A�����OS�+"QTosU�k-���I�o��?Z�BU��yl��a�S8��15�A��6�b�.<N�dK�o����KK�������)$�ES6��W���X7Y��7j ݪх+�C��yF��TP����"ݘ��`����]�{��g-Z��Int4���7����
Y{�R�$<	��v�!ϜcY�#X-�n�:�.0�#��0Jے�,���`g�E�"X� ���~$�9z"�{���<��'�HΑ\_E?�Œ�[���#�|i�(?�=~ʕ
6�ZP~bv- ��Do��t$vI��J�k�.��zS��Pl��U����;��l ҧ�|xP����.9�Ck//��=r�p���~]<���B�}�7a-9��ʸ>Ӡ�J���@��u!H���jp��-�I���ǚV�Pa�;Y+�D�;�(�/��Ϩeo����٢�h��E�v������-�m{o$��L���?^E���m�N"]�X����\�9��be{�h�ʹ]��}��UhF�9�����c��RN�'�v����������eg��Gٜ5�O#�M��V5c`i+6-q?�@t�~ �����a-���'*��6�P��e�Ҙ&(*�v+� �q�8���
��>fiux���8;�&@�͏6��)��\�y��� 2�}�b3	?�&L��H὆q���SM�!3���3I↔�p���fM`�	�6��;)���\qO�W:ePKk���3I`mS1Ȟr
@�N��%��yf��^�y�l(�bՒͮYJ�*'�r������Rc�!9��68\���;3" Ɲj�qf1Uz+)�,�����`�-���n� Ѥ��]8w��l��g�l���Q��r�i,D�0[�Q�� j�lݘ��M%�v:��w�iA�%M}�ߤ�o�����q)���
�ݶ�S�����21���@��y�����<΍�?=#=��dA�B�n�����C���9I�ɯG�s�j��v�R�l�&x$��k�S��9*�~R���=�-���e�!�-h~����X�L�(��/O&,~�]vZP� \T2��\��#U�������s�t�QD�s����!�<W�Ҧ��¶�|����1\��/��y�z}.R�Rˣ���f0D�:U���m���>L�{�r:ĭx�r*�~`-?|��V~���ٟ3��N�9�1�)��w�I�"H�>��:���έ��:m�>�PS��^vX�����r��x��5��p`����C
�wo�dě�ta���X�\W�A�QT�w,�rR�"������8�P�d�6xDm��h'I1ho�ꐣ��L��B�E�M�c�89�C����Ԟ�#X��EK~-��V�H�M�����mV����q&�W��v��;6��a4��W���E}w�<\!��"��_�Y��"���?�Lͳ8�R:��B�Z����d�E	��O�����1��4��%����TۖM(�0���UI{��P-�|+^�����7(sbcdMI��-9��F�4=��(㦀RW�����cgF0Nh���ߍ���x����ᚵg��\����Qg���A�j����q|h���DY���ڍ�Qaa&CJc5?�'I��r2���%ۃ��U���8G;B������E�4E�߽�]���
�ɶ�1��
��.�%���YlNr���$�D^/��rG `��#�U�gӫU#��cut	x�5