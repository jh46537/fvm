��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	�����'Ri�g��
�&v�/�'&r�j�U��
?��A�?��G0"L|��Q�I��X���iTsɶ� �
�.�u/�p�	b�(�N��Z���἖�td0d
$�Ç��X�FN��@��ش�F���7 %�_�犅� zzK�af��n�פ]î��D�]ʳ�n��S�".�A�	�u�!718��m	qJ���N����צuTő�Q�lV�Ï{W��/ܩ�uM���φʨ����,b%(��_ţ�~��v�{�ZǾvg��X�f�Dm����k�����qB�5��-3�P�hK��ɸ��eT�{��͟���@D������ڝ�3���PjQAM��JW��O�F���mY���-)�ݶ�)�^�L��X�7y>�D��p��c�;�3:��1���
�kK��'.W�h���.��tTܤ:ddC�?扑�SZ31?t�4�醀W"ȱ�%V#�b��$�|�ްAF�qg7je�ߎ��Ƭ�7?{����9h����'A��8a���4���y�$����pZ�z��*�]�k���U�!���C�0�?8%���E>uӨ&��3"럼��t���í�MPw����7�vo��Wtt%H봫�9%�~�����2x�-�� )�)ae�y��uT/tI�Sd%>U�#�;o2����I8%iR��*����@��E�n�ZU�f�/Lˇ��z?6ӯ%aY%���ً̧�+(s�<}Z��4	l�����Ìٝ$��xin��gL����Z,��� �J��\>�@YQO�����;��@�>���q��/�����<��^e��wy�.i/�A��_�9����S4���
�s�n��-fp�L��S=�*Cd�A�@�~ˉ���tՠ��\���>���`���a���a������ʄ��֊�6T<�*P��ڬ^P��Q�b=��<���*����:�Z}�u]�˺��!���@��bS,?_����)v۔ni⍓������^f@_�[J�I0s��`���v��0��׺��?^����6�n�#׶�K|*�X��k-�rw�<Ϗ��Ǟ�w��`0��r9����R�"���L�����w�h'���)��͍��@#��jW�"�n���>�n8�zua�Uq�j���O>t�����uo����1	���1�͒�D�7�,Ճ�D,6=���)��H5�2Z�K�Ef܏?��f
1���#߆*jⓧOy���Tӛ5��z�WC��:.ac�B��Z`�A�3%^�!w��':,���J\�W�@_�4��3���Q�������� @��N����NAw1'�^.ƛЈ{�&�2��qL�$��/O�+��|  ��`���d�Іp�)&���G��B|B�G���6?�F��!��3k���XD��~v����+`@�4���S���rrªh����+��,k���i9
��)�V�a����Vo�#�r�h����/�[��/�:����4����t�A��S1 ��tiے��cG�k�b�>�a����v��D�$�)7��y�!� ;pZ� E�8	M�eË5��f�l��p�2d^D(�ډ����|��t!�����/V����k(z�������|l{�6�|��t�q���%%B#3=��I)f��O���ǋƺ� ֓�eD4X~��< dQ���+nI �/	9�z�¨y����2�2���%yOU4T��ua��7>|Pϖ@��ȐɮX/N�%>��{�3��pв��;6�'�q&��+�2ƒ!E���@~Zc{(�	9��[2�����(��d�
F8V�綰��U�J��Ln�n�u&!d�k��[�izc
!�,����qO��]�f�积c;����_���Ř��7 t�a.�v�]�v0L�-���Ϝ������l�9���g�C7��{.�-��oDA��U��5�j>���=s����f��-o��:%�l��� ���5E5g�LA�>�����_�C���&j���Uca1�}�+�К��hL�� ��7g����V�?i�ś��<�|h���G7tF�d�f�
#��Om�A��ĥ�~J���T���ٙE`�X޸n �%�u_Y��"��^�[�V0s#g^�I3v@(�r�BB�����z�Qe���)x%����1���;��o�����+d�j��,|��� K�D|�<#�v���S:��R�-o#k�[�MAq����C�s��^�ڌ�U��a�i�M&�z�4rJ��S��*��%��Ul���3��&,#^�hU�=�O�F�Ϥ{�+=z�dG���y8G��(���cķW�<���o�U��-Ԁ�[�����dDL��n+@��5�ih�'�3�	.k<?����q��!EDh��j5�bş���rWL���l�H����Q%rW�Foyy� ?-_T4���Z�p�����r�]@���"J��qoL���T�|����[��W�UJHH��i|Ⱦ�}x���JE6��z.�?�ynm�����嵩�ca�� ��Z��z͗ٳ6��q�8f4p���~_����O��{��&G�8-<_c��Ng�n��b��M=���u}n.����ߢg*�R��G<_��^x��D���)�|Я�P�A�H�,��^�!�� ��L�X�=P�`
^�֪�1ɴ�h3�l��!��!轞`V�]��z}�T�쪂"�_�0X���eB���;��p�7�s�ι���&z�9|�"ts���3w9Fj	a�rU�P|^4�	��[�ow���Ն���*�~���*��e%x���ԙ��1k5�� �Z�J�J�۽����Ȧ ,$���,�D���%�|����'�>�+���t
��׆��M��7����~D=�Ӣk�G�7b+i;�Gd�"]-����bg�Fzua�grJ}��a�����[��x��cǚ�aPЖ�u����+��,V$�{J���!
��GWB8�q� 6c9�j�tډ)��S�M.{���9�g^,׵o�~��4�?Z����y80�v=L����@����Gs�#�o���v�(ɩbA���$��t����Jz�p������W�TH��f��S+����D@��-Ҧ3�6M�}a���7��U����,��V�JY�z_m�}]d4��V�M�����"d_�W��5�8�}���[����<ŢY�D?��ތ)�e����r�É7�~��Ql�t��Ԕ��	�(ğ�2�՟).`l�	��V�G��e%��y�q��
����8`\M����=�>4��{tLz���V�l��<�I�����������Zj����Yf��f9�7�M�M�&a��+���u4��/]"���<�؏)·�`^�,�(́Yc���~e���X3ow�4���{����*:�8�h�MF�S-���~ڹN���8�ą��Đ`�F>�(X+e	��zNb��F����˳o�	P�J��
$Wt.м�f�ȨbK�H8��7YoM5~7i�/��ˤSV�"���gc�L�r?�?pL�gϲ�*�5����Jge6RY��j��!Z��/�S��qR�ғ�AE��u[p�Ȑ��fd]��6����~�R��`�)�^�YH�S#g�bx*����R
���r�,��>ǻ�J��k��v�S�eTmI3���8^�c�s"�x�mx8=��	b�I=^<�dx�c�h�n��Q`�C���Jm�n�\%���n��n�s�j�cg)��ܬL�4��S���c�%����!xH�V�)dQ{|�q����C;�	-� W�	҃�J�J`�s�G��6�LT������������4YR�,��r�i�?>������ӎ4~@.p��>v����<t���єQB+�8$���p��[��j�й�������"x|����n�V�e:�+!K��=6(�ß2�l��,3�RO*�ȿ�{!�v����*�HҚ�mA�+�4v�&3i�f}'��>�T-���H_��FP��>���~l��D�W�:�m�H��w�.>Y0�.W��,���^�yP*ʡ�¥#���+���6��Ū�PmW_|$v�,cf?ؓ(�^kng������g[�IOήK�cN�-��X�^`�B��l;�=�ԯ�	u��餽��