��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~���y�,����p�r��i�u�&�[���W\Q��0�����	���#.��b�F��%vr�3~��M��`e\Fd�=?vb����4'�$k��&/����ġ�ǸS��f��m�ū������4[~?ᓘɚj�}���5ԗ4
�Q�-����Bqf�\ݟa=�����T:K)kq���%�����֠��9��8�Z�_.l��ͺU�W�孅s��ʠ��#eS�����ѻ�zܩ�$��{���!�65�O@�Ң���f��XAp�}�O���1�Q�n3���箲�=A��)�hΙ_	?�E�c����}t���Au�.4ů=���O�E�^.��5|���d:��3���Ánp)���OF~���o�c8������4~c�a,�n8'M�*����mju���)�x�yci�Qŷ�-d���|�Ө&}ۑ���$9�ג��_I�F;q_I�%ۼ�N�-P���8!䳒��|�� �}ߢ ������	�)��gm�))��R����FV>�{��tM$�ћ��b��ٝ����u>��C�����p��_+$�f ��hd,-J�FG�M2�_yD�|F�5��(���ۯ�������LZ��o�>��3_�d@n�7��� l��cq:*B�7�fӜؗp�6MB��ee�=O�d�hhl��b����#KE\��/8d�N�*n�SZ�&���t���m���n�@~�X��(��� I�,�+�S��QU%��+"pmU�ȗ��������C�:߷�=��@D�B_?*���ڬqг3j#��}�h�A�8
h� �d�8�F����ji��w���8���mV�X?,�3�H�����r���n���b�]dC�!q����C����B�|«T���R+�ل �����FЖ�\��ȁQ��ҿ>�z��o���6bڢ8f��/2ə�Cxh��orO���?I��o'�o٪P*GQP����*�4�ϕ֊e�t�h�>�~3Gt�?-7���v�!�D<��w��Հ����/�4(��t}����ހF��u�����`�[�%�A�����LAd==b��W)q�5v��H |�|ģD�Kz}���6�y��ܤ`w)[|V{�ѧE����T�8�V[C�P�(�Q����zeKuǇy9�+�Ͷ�04����'j��DGN���P�����z)g��ɅR75_�-�d�ƽ���UE�V�U}�I��黴~2l���H�	B횫Y�
�B�6g,ѲJ}l��*h�(<�S`��:�����j��Y�΂�� o8:�)D�MU�7�Fk�Sx����������D�*�����|��$㩕���,�?�!�����_}>�n�_�I���F1 W�6{B�Q�7�k7u�XXGQ��o�2��f_�J���G��A�3<Y�N��;8��ٸK��\0��r�ঃ� -޷��٧�Ѽ���p �lX<���n�p]3JjlS�PN!Yi����Ų|E�xw�#N�rw�G
)B�!@�Y"����}��`��_��}IK�hj|�{�������=37�ۉ�	�Dݿ�Ѻ]Ga,bæ3l4�r�u�idG�½�+���1
�|[�˥�>����8£���v9�lP���������Pw
S`������2c�Z�����p\:P���t=�Fx�4����y�*?�E5��Cq��]�sm�B��' �
�>&g��#Z��� �'���>)X��D_�l�R��n�-�ox�k1rt�!v �j� z���i��E����*��u��?9��"r���J:rΉ���G�V=v��r������
�����+%
+^LU��Poq��fKY��	��)XS�4���>b���љ���df��s.���*��9��"�=�J� ���	���>���i"Ȧ����:�.�y�w���ቪ�E[Zyd;��Yd���]eLv2�#8a�̞oc�E,����[���T`*�.r�a����uj���	���'� a���Y��&� }��Z�4����z�w/�g�F�� �$A1���^��>c2eڠ�}�a��2Y��р�Ҫ�c��T�H�#ʮs��x�����S��j{yș�R����6�t��k�B�R�"�u��	���%�M�`�t������@��i^&��<��O��RB+��J�Q��{����]2���ܿ���8��'՚j=�c{et�Zr~)��9�T����_�F�M�¨��=_�����I����b�گ�yOg�ۆ���h�����>H���¿B^� Q�ZW�.����5@�U�Ȇ�s�L���2��\4Mc���0	����܃�<��j"x	ےѧ��՟�]gg;�`�Y繻ơ�Ϣ���r?H[�-���c^c8�Gm��R��jD��RпYYe�H7g97��hN�_W��f�J7��<Ձ&��7�ʴ	o���|��3'Y�A��D8��"t�����V�j��9f���f�����o9��5�-'�Da��u�����a�`���z�>�������۫Wk�Ә��_��m0G��Lu��q�ijp�6v�����>O��D,"�$y�]&��Tӧ4��ԞA=з�� ב?[p°�!�����x,\X��JK_ �W�`��]Hf�GQ%d5�l���?��qpE����I q�Y����li9�hƆZ�8po��l<��	r�S\�"G}7�!&Ҥ�Ll�j�"���\o[����	�o�֯%q�b� I-~+K�.����	؟�c�(�gxq�kP�ȡj�+r-��:HǦ��ca����UV�:�5�k��i8�+����K��4���R�%��SP���N�����{����Il���
�yQ@�S^J���ˈ�zS�1���Y��-CX�0���S,	-Ұk�f�'2@q�'D�H��3Շ?�2d�����)���4��`v�Kӂb��3�~ծ<���f��깴�\zr8OO����Q7�]� Ҍ�<!j��75ǟ���djz�O|�GAm�7z6x����B��k"�)x�,1��[[F��+���Li�RT������3�<m��'uY�gK��\䷀�5&�TT�f����x�v{;�ʰ�8��{�f�e��i�ų����Q��)�p<�S����_�Μ���k�|a2l��5�'�}�)T]2h�&�R��[�E��� �`G�Uv���^l1|����c~���Ɍ�S��@]���N�њx/�\�O:��_��N�o3��Z�H�.�4��ŗJ�@ �7�]*�)��V��0���%�x�;x�B�W��j�f������qfX�o�����8����@ u)�jH���X\��FSjưˋ,d�|:���; #�����O$Ӎi�E/"u$ԘX�N�g܌X�/��C�#\E�F�L�U7�`���ϕ�˫6�T��{4��^!���ZH��2T�t��mx�Eq��~���f�"L'�*n�����T>H}v��Qke@�S,$����L	�G�$%�*�z��iEW؆��'>C�]!�h5\�<潂���칧��)gcD/z ���2x@J	U��F&�E?A7!� Gi�C�����"�g�����>�cJܗ���UNg�X��kɮ��'�-:�$WXP��Jr5AV���/�������::Y��Q������Hf�g�/v��=�jGҗ��G/�u��{e���K;ǭv��d_��/��À�V��p�b^��&��Gg���|A~�`�k3��g$���#���:1v٠H;��WN�r���Y����B��S��J���똄�(���8�2FGj�?���<�"�6�	c6T��uv�l�,�2&�z	[�1v����s�T�h����jC�cc�����gf�^F6��_;k����|!��TjQIS��T%�Q���oa1�Q6H~�(l�>�����ڻ����T����,&�*Iwt��˪�;�&8��O���]vê�:�#_c�����h��U���X���,������v�o>A���sN��$E*ɣ	0�1��=��[�_.��+< ޯc!�Ɗ��/B 5�y��6���H'���� ��1�v6s�I߻'�����4�B�d��쩵��>7�nO��A'����V4��2����2i��oƘ�=&�գ0��$�o�1#���TA��C�q(���W��J'�=�/QJ
�v���gׇgvv]��o�mL����|ԴN�����eX��(�2WXA�,�*f�8L,��؍��޲Y�~E�t�h��z�m+�]y(�_΄4l�7���$�7t��_ͷ(}�n-��LI�iW�v��Vh�a��5S�J�}�����*%�|��ge9��m���3_�q���&�9�gZ�1/��ȡ�K�X\T�wb�4���ﯤ�>d�6��C�L�3:����_�'PȤ�!�7��v�[v��k]��\v�ބ��{�륹si�Wq���� ����YD��[�f[��!��pr�tͽ2 ��5�9��b ;�Qz�?5x�+��q���|�pE�/��}u��w��{wK�4'�ܦ4��Szl{�;��U1�4�$SM�ې_8u�+�\Z��Ǩ�E`\IF�_M��v�+R�r�x��_u�J��{D��\9���0��dt \�'QĚ�N�!�у��ˀ}�v�����5^!8Eڲ��˙eĬPtXr�w:��[������fEo���B��g
�xƖW���隤
�M��x6�ם���l:R嵼��D�S!���ӚU2��JH%��L���h�8z��j�f\���Wv.K볟_�I���gl5r|,k7�����-ÄLV���Dv��ތ�tcS�u�<%���=NP��`{�I-�k�����9x�2|���u-Ƴ�����7��A��э�MQ�&	=cu ��H)����1%o�cʟ=I��1�G����	�ǔ�Ƈ>'���3����J�~��.����y�B����<���ۚwʫ�����^i����y��E�C����sx4�F(�wq��mO�O���"�V�QN��Hy7�h��T�qi>gW:�
�d��{l��(U�;Zo��)ݽ�����!@��Oo��#~^WPA9�	�>�����cF�è`�w@xPO�h��,s���zNH�Y�)n.UB5���|ּ�rEq7���2B>�Y��9{ӗ�J��s#�O�D56��رw��� c�5�	ą����\�b�����l���]5���#SrZ37&E�]�v�SiPU&-���0H��d�"�3��M�2n��R��rK��(��@����҃��;���� �4���'ҏ�+b�G��f��>�_H���%���|�I�2�h�(*[+�U!))��A	�><E���_v]��;7����Ϩ���4;�� b���I��IU����F�=������2��oRT��Z��S�o��+}��x̙)�