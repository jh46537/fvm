��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}�����)�p����o��FI{�����i7bvx��~�s��y\��y��3L�FF���ePQ���W���n�����Y#Dx}�����05*�鴭n[�R�.�N]WD9���[���c#�����p"�u�]	��U�h�U�H漚~Y�!�[�:l��M`S9Z�EŚnə�i����0$�:��1,MG!�-�Hv��ּ�m=����K��/7����},B�}0"%+P.�W«�Gat�U���bZ�u�B�t�k����*����Ns�)���@������Z��PC����})=����+n�`;�oZ�MqJS�,�X/�B�ɎϕΤ*�Ժ�$�m��ʐ�-	ҧ���$0�A7G�[���rE��fע��;����ԝ�]<�#�͋�VL[U�Y�Q�~��=�����i�0)���ǈ�4G��Y+֬��2`��.IC���3�u��x�ki�z��_�5:8w �}�x���A+ҎYv)��k+���ϝ)V�*o#( e���+��J�>��0�$'>=d��4�p��4����<�,� 9�r� �<_��3]�V�]���S3L�AOAaG �a�s�a4�^�'�̨�h�w�.�ֆ\������apD�Fq�Pr��E6��h,s)�����]��X�U�/�������o:�����F�DE���/ ����YQ��:D0��k���[�����:�_�:#�qZ��jU�iSL�?QgTS�����V�f�hT�W`0����^�������vm�j�Yh�8}�̦�L�;!��^8ݼ-ͭ��yp��2�~�Y����T��L1�}��OFo�g�P-ݠ�dC���A�S>A�v�DD(�(l���/��H.�aòX��jAծ~�<h6%rcxm�h��qMZ����20T���~�Bi�=0ȣQ������ơ�Ur��po��5O�5��|���iߵ���Zw�(,�_��Z�loOQ��p��M�1��k���ee	��E������ч��4,���åD�pt3p�V*,y��N8?���~�� pi*�[�r��� :Ǎ��1Цh����B����Z���h�x�"1]��K�A��*�U��я3�ڲ��A��0��װAp%��6�5̶��Ӛ��M[<O�v0L|9<}hՀB.�5=���X/U��9�	��:����3҄Mp�8�U1x������^ǌ2�7�	0�$��o}����u�/켴h���T��I[8s�+R��q���3{œ��l��ջ������^ߦ�I*[q�U�s�z�څ̅���DP�.�7��yJ�S� tu�o'4G#�mE���K* y$O�臭;U��}��Ku�Jm�˯Yu���խ�����B��c�.&�[�c#<���(G k��K2��m���Y0�Ɯ'�T��@��V��()1���6��6��b���mR��j�ǘu�!��_S1�G�cn|�b�3�
�C�n@?�IM"U��k�^`�K1�I�]>�R]�xΝFy�|��(�"�߉˔�h�j�hf��g�X𾆙=.{�A�R��P�����J)R�#2�ˀ�!��P�v�\20�	�>��$�����_�hIp�M�Pu��_��%��<�"�����=wNU�����ɞ��+��ځ�w>1zڎ	@�r\� -�r4�.�Z��A�+�0��y@?]EQP�AB#�~�h
�Q|{�5�,��N�Pv���]�a��T��4��k�%�:����{�!3X��O+D,1Ț��j�C���Y);
���>X_��EW�T�gJ�_�ct�"��1����\G�M�2�o
�N��d��a��W�����;U��]�r�]���XF��\d4�+R��m�*��/��`������02T���\5�����W�7�*R�E�vК֍���ܞ]��"�S�+�%�۷�AZ�[�!8tf�p�#K8 N��s�
W����
�S_q��5���U���e�ɑ�T��sZ�JCC-_�0�S'n����m�?Ja<�����z~���1������"�}�~l�G>as��j�ٮ�Yn��7o�~�C4A��I_�� ���ԁK�e�e��2��'oVV9�b��fLd�K0Wh�йg=M÷���I�Gخ������b����	��\lhcg8�&����+�6���-��=o/Wܢ��d[跥� �����4c�Į�p1�4�A6��`� F_���JE=ʼ�s���j��j+�,m(��4� P�Υ�1��@2�cA��H
'�Kّ�0��V�\����8@ �|j<�nH��a�D$oM�HE#�T{GL=��{�"9��1�D�埶�/��L�6�g �'
�.��I�WGt�r�~�Qn����b�B)K|���CT���Wꈪ��:�<l��K�lmH�:v�I��UB�9ץ�?��į:#�H.�;�/�k�6D�݀���ڝ4��gݻ?�҄ͨ(�r�t�kZ�_K��֩k�~��/Ӵ�x���h���
��)��b�mF�1�<�X���ʊ�9T�"d��1ZSa���\�~	�{��~����̕?��ۣ�J����K�8|��P�|���2�����P��7����9Hx��S��<�T��j�µ��>�;;G@=e?���^�=��ǲ����l�x��j�����|Yw妰"�zd�����l���������Yk�}��٫U��%�K
�M뒤̨��5KYA���=��_�ěb�����e��fi>T�ИzS����?����!�JM�	����l��"#�I�k*�7]7��p��ڛ%��ʾ�ٲp��xI�	��Bt7u����l)����o�f�@�^ԅ�+ܑ�>K��u�|>8<NzF�6+L�/a�ViN��q g:ܥ;�r�2�w��Z{�U�� �;��À�m,����H�S�o��+x�h]�/�5��\Q�^���	���my����t�ц8���!�fB@n�� Q`6��>��@�@ۧP���Ier�'�(��W\V��m?92��������Q�䄗�{O�>p���T�kvʵZm�s����hhnR�� ����� sE|0a/�?1����D[��V[�1�:>OK��F/�#���n]nA��K���o�Ҽ��'\-�jw��>��3��!Y5�,m��`�6��I�g}~��uz�bx�]���H�k��pF#���l�#��8���~�E�b�Ϗ�&�iEM�,�$��M$��u�ˮsor�1 �#�[N�,&�cY7V�\�� :t��[T�d���hR�:�9+*���5}2�=yQu9Q�Y�5�<��qnL/�g���Lqk�� �$�b�a0DL���U�Rh�kqԉ���t*7�<�o�R~�p��H��z�X183����z�Do��CN����!M:�b�>y�Lx3����� |�=����z�^ҫ�h�%��ǐJ� BF	SO;�u�!TN�j���?����$FI��m�I�ґf�x�s�[��*;�&�F�IS��	�����!�i&��n(<�S<��ޕ֔88:��;�F%�=�A���$�V�'�������am�s"�-��c��m�=��%G�X�ڦ��<*�+�k��;W�gVLOh���`�)p����\6ʉxsιK��;�h�4.��o	�>	����|t�h�9��Dh��lYs�pFƆ���}G�#KW�u0k�/&�[��5h��jH4&v�deu�dK�@���iGd�v|O\I5�,>��
U`W�j��U8�"L�P�y�>*�(]>	m/�|6	U_�߶Ծ� j�~H�;-bP�՝ C�|�כjN1�!�|��Lv��qV���x�m��E��ݷW���V|]��Ůhj�h�O0�{��%�9�l�c�	<��3b�|�~4��6SY�p��s����~��zt@A�K]�|� ��X�]Am3,��J?�DnƤ����R��+!� 펖d�J�x  �{ �D��7�[���a�҆e$���;�ɼA\�ُH��b��!'@��|�/��z��(���fm&�U��{27(��9�/9s��TQ\��|F�q�E�c�c���t�`V��i�o�&C��d2�t�Y����\�[-F;�[�̕�4}䶑{��uN{6�{	�G�r�%n�\�ܳ�q� �;�b�'��l��U���8�ŜٻB��n��"B�
����֯o�M�����;�qJ��[P��Ɓ�k��҃�z�-]3���[�<f~���:��U��]�I==(�)	 @�N���]�[@ ˭iT��_����0�1����I
���)� q�t������5ڥ��{���h�[���4���T�sk&�H؝�#��:8�:��I�Pp�~��*�pǌ"`ļ֠�u\U��<rƌ��Pmxg_�l��c�(a�Q��� ��I��w���M�u�s/z�}�Vhk�/4+S�k�jY�������k��¼;��٩�2��DS�^=�N��*�#CqJ<�x��_���O�"�[z�ObQ#L=�1IG�Κ|7���P)�+�^;L(��J�L�OEw�,'�����*ߓI�P�� s/����?�P�j�8r��b���_��pz,�94]�7����]a�LBF]S��f� B�I��ç���Z]��j���V������PtՃ�Y�d��a���zȻ�� ߍ�*��Z�U+M���w��^��Y>31�(��w����U:ԑNq�N�ffcL6��z��!�zrv&�ݝ���7,n�+���:��〔��X��;��3�eY2�~� &�����r�p�C=����x1�^v�d?7�� ֩
~�����s���m�l2��*&l��m|2{�Aş5���\o��C�;�O�d�2�ۅD�u��]�����Pt6���7��W�-�%����o�d��@��-� �f闇����Ic����#����'���v&	-B��Z�� �;��G��Kj���'Ͻ�ߺ+��6����Pt=Ƶ6��`yȉ��I�Q��@�	ݨ%j�F�oh�q ���GT�U�w<�[��,�������v�,>`=�9f|u�������~le�咢�����rꗆ�l*P���Buh�L�����#��fZX,�u��b�igO��xK��\�G�\ ���,���H�:����;]FR�vK��B�'{aM4�P����0����M\o����M�v]:M�O䆞��,�9�hWb�L�[�Uw��&�fH~:�H𨬕4��=%�1�Ba�r����w�=$ Ӓ\̿��W(���y�Q��6�4���0#3-!���$���t��k0�kL�ٛ\����[)P`P���חH��-��}��#Ǆ�`�n[�(k:���5�i�����K����9i�����q 뇑�2�<6*8u�!XF"����uo����6	+�u�i�J-^�y�_�p6�l�r2���S� c�l�3�>]OR�aε���`E<@�jEp��Xޏլ�!�y�JEk���m����f}�!~��U�I!@5n���k�y��h��
|n�ZP�ق��w�b����8�* ��$�_N��&C[�d{�2�5u���g��MT��ĐNm"3
dX2Ȇ�y�?�R�C��`m��N��<�_�S�S�n�0QL7smi>��Lɜ�S=lA��oT��.&�����JBC�7����m�}&�K�e[�MMakW�'X`]ٚ4�f2���:,����L�w[TJ�(ߡ� �.;Y�ط�|�h���>�
t7e]o&+��bw2�#q��J�c<�O�z�j���N�.
���B��W[^�Ea��U��J�2!#~�4�`.�y���|�ӥ�v[��M���	�RL�>�~�=�(Iw�Έ��({t�T`��q�Mm
2��8��:�����>֟��2'K�%���6ܷJ�lt�_@� ÖO�{����c+�iB��=��}�'�_�����N>]���Kn�|	`�7�`t����	t�߱&��rq\9g�ND.���m"+����F���bb%2�`wiCM��Cr$kz_��0qS����~jn���BRTV4%�^uA�DY���&�c�D&y=`f����	j��4������>�NTݵ���+���6;�N�ZU�@��r@����U��)�|�G5%��������4�i)H_����3�!�Ml=	�.�ܻ��5\ll�b��s_��Z72�j�`�=�l���/,eo)�P�wђ�͊�{����b��}������s���;\�O��M6������A���l���������,���rB���)w�����E6�@jARB�N�ȉ��}�Bv�ڢ9`��`.g��e`��dFVM���}�[�A-�g1�MA�~�%�N�PV�����,47�a�p�}a� `*�4�
�!�Nd�Go�ah�O��2��#�hWa#t��(��.��b;�W�-^Y#h��1̺�;�="\wJ��8d5�S�x��
�w��*���Z�����`Z��ݥ�t�F��22�D85"]nʮV��o�,K����C���~���/�ĉ=]7�^(A,���ܴV��V�ϙ�S�����XTu�ra�yk���4xwQ)b7���8Ǳ���#,���i��P�L4����3��9���0)tML�옅%q�a�3��+�K����@�.�P�-.�r�x,D��;�K�Z�{A�w�Yvچ&A��\��H�A�v0o��"��Q��a��#z7ġXtۥϕ~���{ս\�����E�2͏PGj�
N�J���Թn�!qKI�=����t;9��T� L.��S�Q˔][�|-s;O����5�&���G2;Yg��)����]��yOz|M^�y�d~�=�#>� ��.�ɑ	�0o8+j-|lX��b~_��7�cʻ:��V\&��9����	~�nQ#w�NDe!��V?|1���o���A?�
�@c�m�:B@�G?���^Þ�s~^��A�<@�I-� �*�1UQt���9D�}N�j+�U�!�͇�H��`k耣��iv��|�PlO�!
%��>ږh(�h��s����x��ʫ�dY5D�e�X�^�"���;���<u�2��
��(�E��o�9ߛ�U�v��.�^�j���{9��9�9�S�x�.�nT����S� C�?~_u��	b-�B�#_f0yy(Q�h9v�ڊ����zg��y�嚂?�L�F8F�^m��/�(���v cP��8
��n������D��u���4>"�m��N7����$����
�h(i쉉)f\�$e{�er%Q��<.��$�/[ȿ���sDK�t%
Jq_�<�}H,0�_��Ǿ���g��i*?�z6 ���o�P~AOu?-IHlZԑ{�)'�IxD���k��M.KL(��P�4ɯ�2�F�S�cCM�-�SE�_���-�-Z?J|�����qF7�o͉P.x�G��
����٥8z�Ϩ����$"�_��G�K#$;�{�n:�l��L�]ƂY<md�.�@iIUs�����C̙�WARq�Qn���jP�R����:J��o�@��Q.� 2D�Z�P�5�����E/�	�6ºc��$k%,���0�ߥT.�rREA���+�@oGP����%$?�d�+�999�<t���!��'_���={O���s��4!�ݢ��T�d�ʆOꕥ>��S�$��@����m�����^�͑�O/�Y>���Mۢ�[X���X�M�KS�rp�l�'Qf*ƒ2��nl�׶p"w�?���re�WL����`�.1��{�P���E�A,|=�W�P���Xd�h/���"/[z�ΐ8�m{�Ҳf�%g��1/tnE���T��36!�a�Y1���2'n��] W��;��B"o|�U����9L�x ��A )��Q��:C�q�FX8F#� $�Z�X��^!��m���nxp�Ej��e��F���."��V���{ w�"�"n���P�$U�*����V�	2(�r�5,1Y��q��±#a�~�3��rg�)%����3�>�x9���Dn� \�$⌽��[��l�Hr�?E�P��R�ߚ{y��C�h�L�~��e��Bog����I��/ܮ`0^	��ɸ���G�D �E����h�O5����|���F��V#G~�z9G�f4.3�a�_N���yO	Z�1�w�q`�JuH示�|�#��j��ڼ�(T�]����~X�S
�Kj+�� ������⼾hJi%(c[T��2�nr]a�=���mO1�x[���>�"D]Zۈy����)��O9ۃ:�# ư��+��G%�T=��@�-S�����JzH�����7)�¦9v���JMm�ě(t�ʤI�EDZ��g��7�..��&������T��`�H����E%šM�ǰ�A�tf���fs��	��Cu�3�~֠{3���b����Ű&J�x�T(
�Ιۆ�}ЋNZ�s���X{G�}��Nǣ6@&�)B+�"��Q��r>-�D�#�Fk��5��.�2 �-�B��:C#�\�yȏE�8��5�g�E�d���to���J�a%���X�� F^�%/�����@������K%_Q����$,$*E� �����J�`�@���Ģ�}j�<�:�>�j>۰���%� �]�K4�s3��s�9�Q�BzJ2���Ś����s�a1�ғg��=����vJ�;����M0,,=�5]����&�]WV��2y��ɼ,d	���|*������*m/���`˟��g� B��F 3<��)*v/ԲX����-����k7.<c`r�#'���8�e�l<���M"#���HO�xT9���+fӮ
8�[.%y29�g�QV�?(�y+����n[H��w��T��A�|f�y`��PC��.V�S�F���_�2�p�[, ��1T���>yeCm42uc��w���,=sM��|E���̭[�&�Ei0,ۣ�kS�ĔVJ���}���Kz������Y�S��3gK`��\Jq�K��X˘r��d�Xq����>QV�u:�*��3W�'@�\�N�!k�I��X�>���@oN'H��/��9�"�bڔ��9~�Z�
��S�"��A��Ilg�#c�
��x�������N�j�8������5���xr��"|65�l��(�ɵ<�uu��v�&��
MN��	~p�uN�lzȐ�K #�Q����a$�=��e\&���G�`aS�-��=9O暧��d��Q `	�p�cNU�R�\ �O�^���U'}I<�7�"�"�,?��!��;&����Q�Y����#X�+£���W��T�N�tz�]���/�ɞ{(���o������Xa-����c�`���&[���vVS��?�ӗZѣB�2�fz�P�P�~�T�O
�HE<U?3|��T��k��"�W�!%��iJ�@�zx��pݟ����V���W��x������a�)ɂ��Lځ��H.,K���nz�%2���xHh���G�!m�<�\	�_#�Khm�� �����F%Ƥ��5�<<W#��7l�n���%��-�wf��C�����y��_�W*_�PXq���{�{A�J#s���S����{�w%�����F@-K��=���yFN{�=�[��F�n�r�v�	wjǉ�%�ؽt>ZԓH*�2tG�UPS��Y�@F*(�E�H`�C����/��7k���HN`�h��$F��oAz[��]g6�&V��x�Უ��8oQm�޸t��Ѫ���oEoI|��z���ٴ�VPX���PM�[��>�*���d�LBٞ�?R�˂���	�N�Y�bL��1Ni��)z��?,��*;�ꔛ�$ �ĉ�	�4����	К��r��Ր��iꦏ���[�9�f3�L�\r��n܋c�)�IPJ'L��"���:�, ̱Zf@���߿��C�k]����HsL}��M�1V�#�04y��6��[3�W�Y�5V�]���<�!0�2��Z���R���g��������Yc�I�2�3h�(�g���"EƧTa���-���9vp�F>�9�ߍЧ�,8FL���h)��<��SM��Fl��|�QMw#ddR1�|���#C���}f�[/{�?��W�b˰���v8�A��RQ����i�-Z�8%Քt䦢�$p��o+�z��y��� 6��(9�Em�:r�X�Jd�����:$OsB<�3�x��̜�nD3H��b��Yd�l����&^J|4��|�M�?amZKsƱq�9����ѽe�Np�6���F���޺�s��$������
,����b�G|�Rj�wM� }���T8�=jhz��j�� �bVP�H8�$=�4��Ê<̹c�@ߜN(��p�0r���y�7-<��c��/\�`Q��Ή�ZF�y������븽���=���N�?{e_�̰�\G���zP��}ܦC����(T�S�P��?g���v;,9ÆBӡ��2h�l�Vi��,�FqԿ���xr��y�ZY/��+��h�5~�iY0趽�9�羖O�j+8��!u_���s�sFc{��5q�H�8L�P�J�N��qW|��^�]k0�ȵg��{�eQ N<�@�����҇�Mn?��	��4�����~|��PZK`V5�f�Lꟹ��ݍ 9U�~S%��+fj]N��,���<����a��z�[��<��L�ߊvb� ��y�OZ�u���?Ҫ�ȲE,!�)٪;�N��\�f@�j`��A-O6f��H#�����I����s���(tOD������C
/8*��2%�����&I­���e<S�Qv�E4�c�P=<tgR��������^�	]�G�(*hӻ&�
M�'�������Z�GV�*pfzi��^k��$P�e��s8Q��Z:�sO�3�⸩ev��n)B%������jh�؏��(ep����j�h�m&0�z� �����̒,%���Bo���?Fڕؓ)f�j�~~�����3�&�}�~�}-L?������5���C�����%���H�����FA_�����^o����}�;�G���&�Ǽv~V�����>�B��=P����¿�$7���4��[���{2��f��}��lzG�~8���9�{Q�@�_Y���/����r�F���Ğ��*n]��SM��E�%?:5�t�;��'�Ϸ���Cd�@k
���L�@�?�&�&̅0ũ88�a\U�D=7,�(�,������\9�
U��&V�{\�l�;����}�@�ECD��)�0p��}����q)�Ż/�+@�M	��]1J��bK�ڷ�I�	���O�`�y��9
�?=�z5����謨��j~��L�Yy׎��>I���<N�+2�	8N��D��oyJڔ�>ßs�*��<p�
�Sj>�^�ާ'W�����|h���{DD"`�w�i�<PCD[��ku?��t��8����:���c3I�N���ϳR�#�*ʱ�~3!2y�Pĕ��D
�(!���^�ʊD}�n| ��ѳ��"�j�Bt�6.��xn�o�1��bӖ]7Y�0}Ņ�4V-��lE�"(����4&N�|2����>p.�y�p9�8�+I�4��l{��4"�eJ��:6��)J�ܼ9�|�'$U�?ؽ������b��zɾi0Z$e�,;Z��*kI�WO0]�N%\{m����e�F�'�6V��`;������cs�T�=��D��I�/^g�w'���٥��ӳ͉����'J/(V��h�Xa	���e���NcA���;��щ8=}���V��kF�2V)~0ML �'Q㾢EJ|��}��d���BU����v�bh�4c]����������}� o���L߿=	��R�<5��ț]�86H�-��¿��i��8{�r� -l�S��+�`���f��O��-^;U�@C��P|�*Pkq �LFW����U���ԄdX�P�g;����9u��'�5u�+�6>$�EJ�ċ|9Wݾ��_���ݓFv�k�Հj0um�����d��|���,�J�m�Ei�Q6O�f�]qV�dP�t���5g�?fJ<d�-�],'R��8�i���MqeS}��5���
�_�3�Tܔ�����f�� �\Rm(�Ez�w-����Ѱ����dZƨ%�G������ޯ�+�#��mx{�
vQ˭�����Uv��,f������ˤ[(�!)v�rkAI r�48;�	��敠�A�p��$�J�+�Y ��+m|{D��P�!8����;z&�����atԫa�ۂx�M�¸e���Pbd����ݓfJ�	n	��B��nB��M�&d*[65j(��8xTV�'|�Y9B[9y
��t��D"�]Z��s��z�a(r=5iH����#�aC͇�:��C&�~���EG���eg��rc#��i��P�]yk#<XE�҈C��@�����H����ޛ�Ww�:4�{���s۾=qI�f_e>h*B��I�i����� �ǯ,Y˩�O�(��uy_������"���EW�@m5��q�Cd	���1V��w�'��s�[w�C�S������C����QL����hF�I/D����\xF���H��]=M�;���Br�<�DJ��^�Ͱ�]��^/Y����B��"�κ^|k\�\�ژ�p<����DC�����P��V�ETJW�^���2��
e�F�� �?�N<�����m��g�6=���*���0d����wqK�I�)1Y��Z�G��f�s/�H�bivX�W����i"�|t/�P3��xI�7���Z�އ��Hs���I�ueJT�����Z0qA��1���t�.�i��&�*Y_�Q,��w��y3�i�9ɾȪkZZ�p���J��%_����)Mo���^{ ��7L��Oq~�!ee��4�;T� �����o$��Ɯ*Dm�e�K��ٍ1�Z+�C�\�^����C��9�/խX'�fx��]�0uZ�qe��cHIT�������{U��є:p���M�'2�@�w<���v��S%��Q���X�����r�&auk����@ΚRf�9�ٺ�9�N�t�?+ys)Ec��l����r�=U��g�*�0�������{���D�~�g�lR�`�t��`����ݤ*���أ@�gj�I|�w��:8����� �ڬ���(;}UE����-�A�֫̓Q'����Ѱ~��  ��k�m�y�a�.,��gc6�
��<�L?�j>Y�5Yp�#O$�/D�.LE���}PN)P�[� D���Y�ۼ���y�iQ�o���p���G�uk�KJM��h��T�����T�3��D����iR�^ �#�h���&�YW7t�Q 	T9��F��_A��;"++ܚ۱��Wu#K�{!I\`T��|'�W��d�7���UCm�Ms]�|;��t'X:��(���"F[���f�>���
��Ġ�NJ��
G:�0vNUs�JhZ>1�k������#.疹�W���i)yjW�4�8g��NCe]g-�S1*�I�*�Ps�8Qʚn���h?��v�D"̒��:Zi5(=��
�	��b��U]��s��:��i�qJ\h�&�Ҍ��K�Z�l���?�#�ޑ,V��@N�
c��]�o+�1�;�;Xqh��>����Z�\9�ӱ6��	v�}�A"U4�XϚ���e������.s�kqv���ub�ī+�.GN)m�`���dŵ�	��i�t�Su����E�۾� :���3sA�ac� NX�8�b^K���rU1I�Dt��B%�7]"P�gő>�
��0�`�
3,��GxŹ]  j�7խ9��0B�-�&z�ǋ���xͷ��,;���t#7��W��IK�y�证�5E�����O�`�$ w,!��rcv���Wz���#D$�pcp�iu�#����Hz�V<OD��(�'��ʳ��q�u�y<���\x[��9�Ӷ�q΅��2��37���X���0-Dco�X�RVu�C�k+�d�?�7Ç��,��lڰ��nE��k.{�י�����'.�%�+�zO~�*��M盨oMC���Y�(x�l�\�"�`( ���ә��I��hg�.�?zg�~��;��v��,-��ӳ�Gy���5|�$l�u�6}�f!�a�|2O4��z��@�})��߮��v�:g �rۨ�1M��JqQ����~�:�\��j��;_�c���܍bJ�E��Ԗi�{����7گY����Z��!���S��m����09�8���B��N<N���me�s~d����}/C�aN������%��O��N��*��z�?%s4���.�Ѷ�;�����RWδ�z۟�0$<>�N껅� �<і��,·*�Z�x]����5Cʶ{|%��cW5��`P�-��D&=$�<�:��4�3�)��<�5#.�Bi8)a�E\��U4�B�]/����u�A��/�����2�5CI8�O��6}�?ηϚ"��pC��Z7K�U�D4�����0^3�K�����).8�:��h�=s}���#n�,pcmu�-��E	Ĥ� �(�8�Nk�%$N�~���4�_�r�c� dEz�U�N�r����P��kӃ����qH��/CW�����J��S�r����*�>޺��QB^Dk�[���j��|N����Q�TϚ?i'���7���^�do<��杛4�@%A[M#��O"�A�?
��/_�s���5L c�7Î	�-�^ݦ��IV�c;�`��֗I�ݨ�I\^�z6���cX�\��ӡ��r��{�RyEB��J�i�n]�o�Y	R�|ޭ��A�PT�*W��M�c��[>N�x���/1����u�j�T�����_�hN��Qf8��G�����|�;���� #�G��2A�8��Q����D)�0��Rɦ�S�bhyl���i�Bje���+�	ܼ��N�9���n���y��)�s�m�ِu��Ǳ��D�o�5�<BV����%w\�?r�Gi��R�9>�4�v֥G�x�<!F߱�o(�g���ʮ�<箟6����׌6
? ��|�I\��P&�k�6��1��N��>��������� :(�]r�M|�^�ܥ�7��!�$/R9��R00.o41��@\V� Pb/J�M`wN��6�D�<QWn�b���W���9�Í��[�Yd�J�Vn4���|J�itĿ�K���#�;$�[
wK,KN��q�H)6�+?��V�3h,��&�?ؚ���_�Ov�L�3�Ɉ��a&R@]�]���=Hh�<'���Ǚ?������ry��J�E*!���f1�&S6��6�q>�D8(�i�W��Q���$W�`�x%6n�7�����Aƛ�]Hܩ�����ސ�$�J�dNw���)2�G��FmF#�Z�ci��;L�b�|�;����R�lS)���J(��7�{՗�'��T_��u�.��������b�ZN��?� ܮ.D��ެ�v �����C�Q�E�l�He`�Y�4����V�ܛjp?K�Ot&�Gs D"u�Z����\tw����JՁ^�-���[�
�O-D^m(61E,�t�=�T3P���0:m�l��i�� }fz�јQ3ڃj(p���X����1i" ۣ"F�����8�l�U�Dffl��$���@E�$�ʂ����oH����[�����l�`�!����e� ����l��Kq��%	�Ac�;�:8��E��׶q菻ֽv�7�w+UZI�gѱ�޽�eu�p-%��r�m!`���RLЌ��E-y7��v�-Q_X�%C{$_@�8ԑif97*�9,�iZ��Op]j1��.�:�Ae�"q�u�Ͷo�������[]�(�����p�o��ze���s��4L�E$z��-G��A���S��<|r���usP�W���Zi� �CX|�m�Od^�@���>�9���(@>�&�s�TM�s Ƭ3�"=D�����V�cF�mߎ�E��A�0�G�#:��Q�WPz�˻ 8st�E�.�XN!�"WX 
����͔	���n=��Z䱝�����^q4]��q�?�W�(�E޸���{/w��|�G?�;�iԘi@�z���������E���V:(-Y�},K�O1�n� X��zQ1b(��GO���{�*Y:(�V�F����0�] �wď�x��5ZQK�;)�q?�m&���0e��]4��Z��g�g�8Hc���$x[/����qC�Ԫ��Ms��:Nmß�g���[�X��K\�B��g��E�-M!j)���hA�n���աz�2�ż��6}��-n��,�H��姻hp$]��n����"��,�G?D-�`D�uOV������FE��&/r���pT����t�n�6+�?�p%�©�9�YWK~�<&P)���"n[�c[BhD���	C\��t���H��f����� SB�G2�f�i!Ř Nj�F�)�>�ݎ�,��O/'MN��2'�ª�*b���R����������d^^��y�:m��AD0���H�0c�Q���C=`���-.hq�q_�1��k����J"A8��꽨������*�Ψ����C�y�-�I���W�r�}h9@,U�"�C�/:�	�"�\^?ĺ�{���I��E���z��ɿ���tlh�*د�{�s����uHӕu���(E����G: �%#C2���<��1�֣A���s�H�F,��ILi��6�
�jFm������̀��	WE�����V%�����{P�x@1A�\Fч��,A@l(�B��iR����66@ֵ�>�D�AD��aP�l�P�Qr��g���/f�C�魍WST�k"\�w6��<j���n���7yl4�C�VH}�C��K��4��e���r6�M�^M|/w�������h��	�����AdJ�� [-8��NR(HᰦR[�&
���{��m�QB )�&�d�ɗpHd�|,�}����]�(��}~�\r�
�L���[�{���7䴰�o�_op"�eAsE|x)O��{���f��]�f�e �L$�Z�Ty�JD��ު��F�����9�g��\`�ȵE}M���˿ݑΨy�z��T�2"�QA����·Db�% �B}:X�0Ϟ�./*�~��U�A�)qS
���*n.i6����j�$�o�d��<��KZ�1V����B�vƢD�3�L3K��?'Z-�N�-�������LQ�9���A�����?u<]���2p���5�}[�l^)#�n��7Q�t�gAVS�ُ�2Sn��;�(�*�2���׉�Y�y�-H׏�M�Fg9�4��Kh��p����X�r��@2	<iÕ���@$���1���?&D�,C�݄��(��*@>�ct�Z�h�[q]<�D{�d{����Ԉ`�ִ"0�MŁ�>V�k;A���Y��i|�.e�2��NAU�J�&;a�&I)��)��!���S��
i.�њ�x8x��ŧB(�/��{󇢿��e�޴̒xu���[.P�����c �Sġ�4%`oX{�١R5T)H��5��Jc:@�{}-�\c�믄��
��o��ko�cѬ|���t����w�Iv=5�
��e���&��zIN>��xP���#.8nGz���l��g�-��Y��Մߡ�P��-���yҸwS�9bZ�T��5��~l�	���_#�p���ʌ��{hV1����|�e������y(߼� و {�мkꅎ�y5��8"7d��T�i>c�� b{�xn��ΒD��� ��)`QF�`]_c�����,Ҟ}��zI�>����x�$��q*~:�� \�kRQ�Դ���l-��y>��&o� �q�4��\b�w��k������k@���~�`��_p���B�+�N�ҫ�"�8k�������w"�3\M�x�>�?����}���[Zg��"o�xK��1ESl�ʃ����� pW|��b���/�;*�ڈ[�z/����l��ʿq�xbr@+-�q9/�T�0������B�;�F*�6 M���js�����������Թ�Φi{� �-R���dA׃�(6`' �� �irT7�.�m�j����E�x�qy��
�
����#���Wb� R��vU{q��#�ad�靪�?����<���*/[.���҅�|��Y{&��Z���}g����3�9���A��&Ԙ)����,���Y��e� ��L��?���X�[���'^d��#�gT���{�G��+x�
��(۸�;h]DpU���6��S�7��z�j�p;r�Na4���skGo�a�ï�tx�ڪ�?�C��!�F֡�x�e��c���@kOLB����R�+�z�Y�YM��˭|�ӟ�kz"�n���1D�vk�Oɂ�]d���T��%���i���� �Ge�J=�p4,���5J����;R���J�"��צ+";IW.q�0����d����<UOjSdpRd3N��]䂄g?N���Bqv��x`l]�i�_^�"�p,J��%��ԗb ��B^߰����ң�,7��$]o�l�d�?��zܫ��W[�$�4�ڨ�9��i�� SZ�����w��/%�7��9�P��1u�
"4�e����M���8�� *��&��}�
m�k�-���nsF\2��a��=.s�z6����g��%2g@k�[�h8tk�� ��G���+�VQk>��"��6d�-�>z��X�q-a8����?�z@�9�lv������M�h�X<����Z>oW����g��	JO�:����G��%������	@�.*�o��3ѷs�z��Gz�[�\|�uv^H=������p�Qe��ï���t��ƪ�& At4M�/>WL�:����-�i��k�g��g�6H�*�����@9���g�~��-7��GR\L��L��eM�9/֘�^E�M���s��z*��3^�v�I�KףH5�<)��>�/#�s���@����1�ۢ���)š�$�za��8�Y[H�I���ż)j.$(�a��p!�p��zbl��aC�:���G����}�@�H%��c&<�������v������\欌��
�:""�7�%(p�&��?�JW+Zh��K�Bʊ�1?��n�C��F'fA���ҥ�%ۉӛi�����հl�Vl �G:b<�`Ř������RI���P� �vS�������ҕA��>�>�ᶓx�@'3�Nb|ޅ:	�nN���������9UFA���:y��#Ѯ����y�� ����?lO��zHtҭ7(�s��
�P)��m���B��1�������"<��"K>�37�m#��b��A���oyN��ʽn�z�=��i+63})�R�;!����[���!*�R��GA��T����/L���iV"E+��.���o���,7t��i:7�-�܋���N��u��6ˡ�5�$z0���7���"�^�W(���3i�R�Yӎ2��7���r�<|x����7�%��1˧X4�t��k������W��zN�P�H�	�y"����7���m�Ɏ�i[{�0x`�ur@�K4�\hR_�~񐣵����
BHݰ$/�#���cI����ܗ�*dXj��<�)�=[d�g0���+
����1���z�T���6� z{���%b譍�����F�8	���m�� ϡm�c�n�ɍT�ߧ#�)���Mkǳ��*a��_�%���2K\S� �4K�5���$%Q��h{���vk!&v�汤J`�Co����I�'�b��yלچ�r�$�ڋ�+����Ŭj��ʢ_����AٍD�=���&�s��G�GJ��.��k��o���	m�j�)��Nx�J�d�!�r>��1��� 蔩��.���B�xG��}�O�ƭ�@{ ���YǉnݰS���xxB��.�r /�pA�C��K�#Y	O�k�\�{p���nط�d>�x�ű/�
a:l
Y?����ɘz�IFۈcD�'�v:y��6�)h����Mj5�s0�ú �ЈF��P����^���������9�-C;�2�7	9��OV�9%`N�������?�{�>��U[T��݄_��_�J�A��GDBh�����O���g7u�"�(=܍Ta�Qe����̡�c�&=�j�O��߽[v���4�����%�]X��� �ť�@�DI�~>m�W��h®E�2���B��>���G�'<��3��9H#��6�ˣ	��=�!�O�8%�M��-#��>`�xZ�D�����a(V��>�����yr&���4�j�@���H0�e�a�7�p�c"��xQ㡚��z�V�*{|��J2�S��Ѡz��M�!��%�xEU¤�Z��b�3�%�2^�F�Q�u���J/9b�*@����0o+�_�a�e[���J>����w�T ���dI�0�� <�kZ8�E�x��}�|��Yt�N��.>>���rd|�gY��V��7ii&��������Q��n�Q^�O��T}�'W	4ٕ���Ti���,�'�FdF݄��U�D!bZ4�_fR)/E���@5��ϳ�%�ǚ�af�N�\�@�K׌8 ��j��m��}_b�Am���[��]�cK�t�7�����u�L����]���o��)��l7����s�@��0"�v���y�,@1����\��Gy�-4�A��	��w�=E'�'J�q�ֳ�,�	7�������Hy�|Q�Mͧ�oK)����d��Qo*�g���s�jZ�f���=) :CNj8^���܄H���� �J�Mґ�s:�`����(�ݓ2�L���ް�]��N�3���Ij�U�l�ó=8��2~�	���{��VY	��G���f�7�������9����"���0�DM-歔��
���",A'6V���U��J|_!��ҏo�=�4�B�,�N�1��$��_��b_�S�I�-?�w�FC�����I�C���l�6�fGD����EA`�
�@m�:��-i�w�mj�>9��9+��{���sI:�~y.��	2�;��;@q�*�[�4p��9u�c��*�?�|9�tȞ/�^��i�i�b���v�1�q�(i)���Qt��GȬF�x�M9r����Z��zʹp����j1l�����.��Ó���,)���_��$�D�l�GOo�p�
�"~�;������<��?����&�ۗ�4����B� � Q?��6��ܬ���2���a�=����Ι�}'���n!���,{֭� ����z �:�v(�=�%��{������\樕
���hwFA�蚜*y!��=ӳ
�°�/A�F��H;�P�T���c�!Or����'��x�`��C鿪��ƀ��n�.9*
Ҝ4g��Ꮾ|/k^I�7�И����@��v c���`W�BW�&Hd0����	�&\:}_o�Z�S�c_���Q��Ή]/]N{�~r>9ꦎ�2�^4����&	����z_��C�q҂�Ki�(��zT����~2�!+�	Xഠ�+�cP�+���|�㭞��a�z�>j�#��(�80?�	�3yt������'���d�	�l5lT�Y%�A�{��_�@&�,�X�r����mg�{<qN�;p���}:���� 3U���&�'�>;)g�1�F�+|i�\�
;�q�kn�_vIf+F�D��e]�K ���[��%�gp�B�&z{U(4�oByF���r�j�,��sm��>ŕ%�z�B�yf�۴;p:ݚ���U�g�'ڦ��X4	%�5I��E�aXVc�2y�� ���\�(�;����x�m�(ץ(����t�)�n���O�. ��E�G}J�Np�l)�9�~3S�\���|c�1�a�y���my(����(K9{-=sr�}8����Vu�N��!���\X�/�R�����4���˜]`\�=+K��tC��u����K��ҢVq�?��X<HS��Q�Q��DTT��<p��k� �FH��hY���=�b�Xk��,m-_���R�y�=���%TR3JIN���}�~g���,E���ȶ�%+������mp�{�Dp}ޤ���;R��&��}��߮7`W�_ur�!�+�R��s�`>1"��o8J��CA�F�Zs��  6��j�j�n�oZBi�1����"��@����·Y��րP&�Ld3"�5�U�51"m��6��n��X��F�	�C�56�����A�W���0�M(������A/Yx�a$��v?_2H�T���՝�>^A=F�;��H� ����w.��8؆l��B�����]�N�����y�'�W�G"���H��_Ŋ���R�2ꖯ��K+C�=H7�� �9֑�JfQ���b�IU��Pڄק�Wd��@}
�^�-��3���>eW;﹪v�̸�!Y���/齓�\���S��1i^�������]���4_��zv]E)���7NՇ���gm��W��]�%��p�j��o`V{Ӻp|�Zh�����V��/���� �h&�0i��8�7��^��ٯ�sԉ�LJF���"2\A(�y��� ��k��$��m2�V��ˈ�X���.W�eђ�3��&��]-q:��&8�����A����A�y;2Qz�#�hleq�V�~�=̶�}hS7��'� �T�<�p�[D��(fQq�'����-c:�w��'�X��`� �h� @*�$#/3Ꟑ�B�Pf������ ��\9;1!םԋS��&U]�Y��d0�<�'�^�}Kص��I����L�I�DlU8�m�����S�s=緸��$�p��̓�Eb�x�e��Y�H��Alh6"mA�:o�8��+��X��a5�0�
��b�Q֑'���#�����~��O�׍�]��m+����2F��t$�X�_�*���\�K����?�wC�8�N�e�]�@*���5b�1L�P��e�U���x��g��������'�H�꜂ḑf�tD�ى���������˷Q(�@����.�:U4��j��v�����e���6�	��W�����cD�H���k�
D<�7��[����N�l�O@�5"���� �닄��.W_�Ia��<����i���-�f.�Z�(Y�dK�9�%��\��X"�c������?P�r�DC�~�Ef��P��?G��u��߹����N���ȱg��!��@#�����!�u�0O��br�ɕ(���^tp�-�s��P%��Ǭ@ǃ�2�����A^�hsbs0.�>��R���z���~��Zf�A"Ndcs�ݖ�~��D�1���3��Sv�����ո��l�v�>���I�` ��q�~֭�;Q��V�$;���
D<��UهC.he�/h��l\�W.&s�t6�u��ā�W����+A�*�/&�E�4�I�[0�`����{�W��n��3���1y@��Qh|
@���r�5B��H�aW>:�<���pm
�pN�T������l� k�=���#Pj��م�>�L4{[�e�����1$=��tٍF�Rٞ�⃓�0ݾ:gJv�C3{"0pP��v�2��`���`�Н0�C̴��g�waw�߮f�ɿ|#'K�����-_� U��J==�=ЛA
e!gp6>͂-�=���C6�DI1��Ȣ�F�׫b�a9Y��H^Ô�aJ�X>3%�8<��6q�	�iDѓW4!:�쓈)��X\��ܺ�k
i��>�W���&h}�#�@��V8�6�I��"��nݼ���53gVi'�x�3�a�5����?�R��{K��ב��r&MiY�4�W��IWu�_���Ǫ<w,/$d�YD<�N��>��I���"^{.)~�W����l��;~�l;��������'��Y���<�E)�F=�4���(�F9r�Czb;k��'��e��ȱ
��Fv�t����\��&��9.�� 0��ES�}��d0�y�qV�Ǟ��[4[��x���TNDK�u��yu�t��L7��l1	0�^%�͍OhI5Ǿ���7��ޅ����gg7��!o�߸�K�i��"�ü�Ae�;�� 5��ƚ������u����ް�6���9;��	�BT�@�d�B�u+�3e��]V���P��ӆ�E>ٞ#�A�42��wm{UL̞�^�k3e]��I�$��)�_�����Ft�!u�@��(tW�סbb[��	���Nv�aj�O �4�z���7�;��7�@��R*X�]�9�,T�Π,$
�A�Z�s�zX�^U�ؖ�z�f
����9ԔGN����ЕIC�A$�:��s��0�T���
�J���W�.���k���WEPȬ��������b�����V����TB��I��ra��T�y6��[?��\�	3��v�����@Q;��ݰ�d��f�/�B�48�I�)$M�F|)��H���Q9Ln�/���YϨ�@�7%Q+y-�4��Ƙb�fL�)a1��%<*zh�7��Ζ�U�ksRz��*�q��ۅ۟ML�lҟ&T>��t�`�/�m��Il��ŗG��$]�>�[�6<�cf����C���&�h#�g��1ٶGPq�^!��9�o�dS畡;�#����N�z�G=C3Gys�]�]�����#�³��k
̔*1�<s��t }H ��'��\,�l]� Q� ��5z�ߡDm�7ΛkJ��9T�tR�؉Y���ɱ`eΥ��M��&������t}����+�	p�������a�q�M���$餘��OYc6�>������	�"#�1C���+��d.�UYZo���&�K0��-����E�3��:�,<V`W�;Y|3j�����A�T��֎�G�!(.f�����4�j�n�����n�q������Et%�}K�#�����h��
$,��Q���̓�����A<��!Z
z������߬��~f�w $v�.�J�	�*z���{w�(&���;���N��1@�ٟ�i�:�'�p���.˾~�]�W`��t:�J����)��7I�#�-{{*���Fi��-k`�4�r���D3m��ž�BPYx����WJY��N�%��k�BX^~��c�QY���5��hYsݚ�Ã�I���aQXX�:r�����=�Z�A�Nؔ�܈_�J�xtJ���Uy":����&)��[0�̜���y2�t]��5;��	 ��ܠ'�� U�m�A���\�|�[eB{;��!�Lo��z�����,]�!�\�U8L�Rؠ^î�7�aҘ~��*Vo ��&6��m�����ڟ�0��R7ܢ���>��%� �*����ٌ�a��p>��xb���,���W拓ьR�m �b��; D@�vV��=j���Ј:#����'�Þujoa}�+���dzC0$𓐇����,\��H�l����"��C����x���-��gdC��8��"�YE���R]=Ѕ���-����
vlEt���F�9s�J���"���8.�d`7�Bױ�u1s4�����.�������k1i���ࢴ���!��T_<���|O�:�RuGx�%j���J�
��_p��: EP��\}��;�����C�9�#�i
ɘ�5�(lHJU�-�~��9�DR��H�&R����xH�8�t�J4|f����K�8�(�v$9*�]fv�xS�B���=-1|{��ڰ�g�m_. �d�S�S�j�Kd�Pe\�Y� 6���_�@�$p;�ҽ�P�+{�;�qR��T�P]˾䮏�#�9C��̶��;����`��Np&���!N�{�\�2�C4��"�l��q较~p�՘:Վ_�9XB���V���fr�0(��l��g�3;G6�G��e���,��1bx"HG着�2����)�"W���?R���6H�rD�3/sd9��Xh/'z�<��C�4�v�Pq; HPQ�2$o��'�Q{;�3H�wg��]b%����N�� ����r����ڴ�wS�T$�!��jʌ,f$dcIls�[��ǆ�[��9��
�Eb�����հ�馚N)�j�gJ�wBzOZrT+#�T�cxEpr,X{8���Y�G�H�Ly�p��x�����Z���D�\����m��ZK��$��[�9Y.�;]~@Ή��&�Yo�;��[R�/q���:� Y0xV���쓥r�
�ܸ�I�{���Sh�]��c��!%5���|� �~~��.ޑ��+ShB��?=�`R!m[��'�N�=[�М��b��2F�~�z7��8m��H��$�`}�3�Z��&Ǳ�|E�e8�b7v*_��.�H�����L��TyVN C��[>.�~��`��������^��n��!����׆����7��������/� vn����a����v�8���I����Cq��I����|�����l0a�}Jy*��%���µ��S���3̔�0�?�J܏	t�� ���l�Y���������!�` 5��"*fK�/^걣LwA��v��D��?Ra��7��/FF�
��qi����t��/n�Oyk�٩��|x0������^h���+��c��p��R�#�������@�%p6r�uB�i5<�j?�@��w�~��-����������^[��C=��o�y �8<0q���P��iu/%Y�r�PGPh���	��o�J�+�����t�#=�F��t�!؎�o��(���_\����A���]�����@:��o�N@��k|y��.l�#cP�,&$&SM ���y���iܹ�����Q�9�u���x����Ői�$�[LI
IB�¸‽Y�����!�p����]��
n�0�e�)T�Ã��^ ���!}r��u�r3�0�y�����L�w�.�1���yγ,�Zmu cW��sI�UE���MYσ��.9c��> �k��]`�N+Xg���J�c��$X6V����ĩ�K�Ԥ�<��ǭ��gk�c���?�.��~@+�_'�;���6R��ʤQ�nb��ҨrՂd�7��&E�p��u1��L7p1�jquFW;�yT���VW�
"��X�@KtqyT�$\��]O�v��-�d�zsqѶX	�݀��.������8[fM�hA����p���i�������f5첊;��XQ�^l,9�[Q���*�{v�<?X���w8ɛ�7��4�m۸s:����?�4�Ig &崞e(��\r��ƴ_Ep��e [-W��Ib�ף<>�s�{�z'ĵS<��!	�y!QD6���N���̓"����fI��{�ɟ��t�	S݅bN�4�tqƹ(F���KD�px�x�<�^�B�R�c�K�q{�~�5��vu�|.���PV�&��o���a��dS��_fx91�����G�T	H]�Kqof� +o�&�IH���&��C,_�s��׿ɰ���h ���Eꙋ�N2:�[�������6�M
�2>��Q�w���+��حb?4���(ʢ@�@�D�tG����}��A����Xة^�x��ۀ���Ɲ�+^���>�V���@�[�!Gg��vpq�׮R��K��}uz
��
~y`}� ��/��x�0>yؽ�V���׀���h��$���2�n
=�E�8+���o7���d�ꋍ�e��o���
��9.v1N�H�,�`T��Vj?���^qb�L���_81�9d���x��#pweKd	R�k��D�2��B�6�s���L�s+�`���~ \o)��ڬ��BtЗc�B㵯��W�1P6�Cb83��h����N���	��ֿ�ꇡ�V�����n�/#ǿ����<�r��"2K[W|
0�5�OH{']X+�����je��5�8:��}��sY7
�(��������h��T��}�J@�!g>�����?��: �0M�xsF��Gv+�+]+�B"�*��o����!?,R ���($#������}�=F���0�z=?=��Q���@�VU�d}t��z���~���)>�w֍C���?�#�R9�z����ܝ�YϱRU�|;qBro|��`�^�V�´yy}X�~:O���lo��C�'��� ���?��e!J�Lc�!�io'�L���~r��U!�i�Z�p<p�a%�xt5A�(c�i����7cY}���g��?����э�ƿ���1x�B7 xn3���;Y��ߙ�5G ��eѣ�blͱ�5�w�Z.3�F{��LL���eA���]2 �&Ӡ
������)��9���+{�*�H#e7ք)��g��c��"���v��������]l6X?ƺ]�Nj-#���sD�ū>�=��K$X���� ������y���Z-ǾV��@9Iu8Q��a�X�t���D�����Vb�����b���*�h?�+����S\8���M&�]�*H, =t9��_]�K�!��� ПzN�S�����Bڏ�μ�����KSP�!;��>>��MO��mf�8��QL�~��G�$X	�X�{Xz8�=�װFJ+uv��
]?j԰�(���|�,؅�GS�~�������n���:����A��\dF���bo�k�ژ�_l]�r������7�K��wߕK�,$-�;Yo���y�XY��g3׆�\���l�y��*׀i�9�s8k���tG+Qۿ����ħ���>qQP�Fg���f���7U�%x�}�a=��1����*�!�o��l�b̘�����&��<@W|d.v��kyӲj	qT�5�*�_�H�k�a�"�t�y��b��G�oVS.�=�/CZ�K^5��;���$��|�)ٳ6�k�M�>��8	�킁m�!��?�~��� �-���4�u��R��؅ۘ Y��	��r�D٥��T �̞<��om��"�������%}LE��URp�'?�yU��+t����IW�o�:�h�A���qN�i��{�~z���a�h*�� R�$�U(%<�wY�_(D���ټ�.�W���=wƞ�׽�����d�&H�=$����iˇ%�����\��9��)��Πe����$��	�m&����ƥk�Հy2=L��,;b�����:j4�M�J��o��ă�(i���?ײ`.QC��ڝ��KJ��[��U�P��v�g��e�$ �j�7�U�ts�c�p�KOs\�XH�\ʚ=�"��)�n=�
0�����^ܩbi��pY��]����������k��\�j"婈�Q�*�=[�|%9.��Yt2:"�B��Qn�\������;�e��(�8}�T��yzK!�֒��fw�E T�q�ۋ=��	=����?+��
�Y�W�z$���鞮�`�Ib.x�:�I6���?�S�:�%.I�:w'��q��a�q�,�0�(����\2/�a�:s.d�?W���p�I�����!�=|�w2��%=,K�M�%�ܳ$#�g=��M��1����*1�Q�-����S;Û�q)�K�^��@�V��*O���)��:&�<���������E�lV;'_9j�ɉ/t&c��ǫ��gt�7~��/�^Uڥ���yȿiJA
����<e$���asİ��[�h}c�ʿ�&�� z������n���ZQ��*�a?_mK�����h�7��T�;�
�9��Ls<�IO�5Z�i�4��G{rJϵx�__��Ӯ��C�k�
r������f33煗��Ƴ+o� �x �����Q�w�6�m$�c����d���DKuw�gX*�5�QiE|����1AعZ�(ە.��X�-��`��u�ܖo����U�O,6tM7��CZ��!�?ra����P����uV�߱���/QV��t��̀Ӂ�h�-{����N.J�ڳ3�0�aǧ�̍��ë��.���Wy��e��GC�\K��sу��dl�X�r怢'���$�V�8(�:���?�O�Ya����b� �X裠[qnC��L�'~�x��/�o��z������=��a�5�%�I69���q&���о��"���H�����F��T��,-b���cԞ��(#��~"g�c=��è1U��k���R$��N5윶���E�\pd�0�=�r�oD�
��ɰK��w�f�ʹ�%+`BRs#Y��fP1U-�M���n�h�9xKi`t������� �ȘŢ�Ȅ'`,yZ,�;�"'%�l�Ƅ'��^h@�6h$!;S�rDt���1�;oKb��
�:����[YR�0��w�,v����A)��t5D��o�+D7F��O�p{�2��6�!�7�����^'3��S9�i"�~�vwGK�l��b`��8N���Ҋb'cx�~��_|�T����W�<ᑐn3�Vd�'cO��*�j)�����^��'�)�?�#��rb_�ѳ���;���f�"��@����Y8�v�mh6�z%�I�R+��MXp�gR�i;�$+���?�b�k{~BF���8��m�����B�8��N��zr0G�ʭ�ݨ����0�S!KN�>����. M�*I���772��	15��#E��>-�f ����M*�����ӹc�P��F8n���y��"���e��nƄ��	mgvx�	�h�jks��V$��Ӑg|TH��3y�8����e�G*E�cͼD��sWb�tG�T��>WP,�"*��J/���Ď�0�}���s~������޺�M���0��p8U�Ɣ��T "%�F?J
A1 �����d��V��:D�X�5'fC�0��ߎؒ��+�PM�:��2��/	�oސ�f�#��?��Ϊ؞��O�@�nޓ��{5U��Ҟq��5��1�>R��DE�!OI9j��	O�f=Y%�ٻ\���ؕ�p���`�0\�H�䘵H�e��A����X�DA�$�k�.ay��պe��._IInvî	y�l��G����v[Wø\�5�!5>z��mI�b�g�j��f�M�zex��e�UR,j쟮B����v�/s1bV��=&�YgⰃ7~\�[�6�H��������]b�?^����r..���bZ r9}N��I�\@�i��������w���G;bFν��+��L�����{l��P,s�UJ<��ɝG ;��9�R�@%��q�4O�>�޴��VK��{ɑ�㞥�OU[�(�<gQ3)s̒�{@M��� ��W�m����G�ZU��mh�޻��8������cAH�{�cR4�Ά�'kqy>'-|o�.Ft�)����kmcR驙�X���O]�s���aZtoD��_[�c����p��6�K��;�%�$�	Ͷ���hJ?��������U
�k�^����qZ�����JoإQ���3��6|U)q�՗p�ڣ�b�2��{�Lt�:�Z��c�E����݉��[-R��׌������Q)҇��Z�Ѻ���!)����p��e�DI��Bi��M��p{����X�g�'�q�S��*��|�n0���Ɵ��9"%�ЀLM� ]�"�h��A�wr~9꿘�@���T!Y�����M�e���`M:��������������.-c}�0*YvIۊkJ���!V�R��e ��6$_�[�;r��{DP�E���$Bk
��%w7b1�D���\���d^UX�0ȧ�y����}��忀X|L��;B�:�E��'VW:�ĳ�o"���%d�d�������_��蟙�EoFRX��/B��1k/N���}�v��_�9��J�d$�^QO�v�Sj�W�
A@ъ� HԖک��L>� +�g'�]��Jgf���E7�|�Lw���-�"~�Xz�ĝ�b����wETXY�*����XV��wΊ{突��� Y�fRY,Φ�-����$�7��t|}�/��Rղ��J�'aP���`9Q]7\��F%���fMk[L����
�O?a���ɮ���$#e(�$&� &Rs�m�\<TS21����|���/��z"B��t1:�R�����hhEx�- z!�;O��Ӈ]�������]�I�7�^�I�I?eQ�c����?�q�����	G��`����_��$�� ���P#_��^n����?��wǺ�uQB6{��HEj[N�A��IV�sx9T�� ���\�5X���e��$�L\W�f+�qʚaS9ጺ��ƶҒ��x�ˍV�r9��[�@^8��4��{߰��S�R��5G^���朾{��i9���Ӷ[��2�$/��6��;I���'M,p!��,kxd#��lh�9��C/^�#���L��xt�8^�U�9�C�s��o�ER�S{v��"1G��Qל��,�� ���^U(�R�A���i�Lqnב	 L:`�秚o'�+Z<�L����2�v{k��6�g_5��[KV����Q��-G�����6���b�Wg��P�k]�!�P���O'!A١越Ɩ�C���]?f2v4�8��A��Bh4˱�5�� V/���MF�g��E友X������;��^W������+{g�- {�dq�L"�]�Z� �t���w��I߂.gZ�n��j:a�6���H!]��q7QR�׮D2IS�2��|0�u9�{�)�o��@�$��mM���Z ���H�KDnm$�g�X{"qZ��n `��*҇vI+6k���n��~�*���y�4[�r/Q��H�d񻅻����Zw���ǰn��E���D?��zNtAd*S�߸jQ6N���]Ī?��gN�״�tr�u�����y���u�h߳Xe�+��-5�<I"��`����W1�&yɆ�S�
ֺ��"���J<��~N3n+�}z�s�'HN~'5*��<�׊2�	!N<W8d�\��^���<�[�ǖR��)�axu�W{z#��O��UF��"��K�+B�׵7���?��@;����>l�
t�o�W������3�.�7Z�Y!?��� ��������s��WAژ�3e�4A�\�ћ���*3�$(葧��L��{�9�
��AK?��*�C�7�r<%���@���G�[]$`u�RHn)州�-u�d\2Cϝl��ԡ=��UŦ��%50����i��rz��8���+�Y�l�{�q��+�&�e��-���9h�o7�G-_\ߴ��A�7uz�*����&V�I��GE�������ݚ���)6�{=��U2�,�� �����W�����;�Xs��OGu�J����5�!i�����l�˥gn�^�˶¢P 9��&!��6b܀�[���lXy��,%-WB)͓X�j��HȯݲS���U2�sI��l���w����F�fy&��e$���{�ԝ���ڪ�"����S2�F�H��z�zɽ�Z��t&u5�,J��u�<�I�`^C:(�g���c���1R�AFϬX�<���w}�4J�_��cmS%Z��|��s� ����U��������|��݄v�������.�?*/�C�u5�?^�{��Q1�Dt]��"T��y�n'w� ���Z1臼؍�����h1�Gh�"�������uZ��ۡ8�!�v���(�����g��ڃ�$p�^�z{h4P#�o޿`�y T+�FԔq �;E��Y�S� �4!����Xe(LDQ�+n���OR7ݬ<�x��7��rd�檮����P���n����]+��~@�h ���ጯ@�!T����Mo_~;�	7�k�4f�4�`��,�T��d2eދ����U{0= �ډ���fM�*��$*C�C���G$�R��.� ޝk>���F��U�)���`��&�H�`|��ha]��X �eW�4�x�� �ú��v�:`��CzI����;����-M��@�bW/��/�����*���r�����F�ⷫ8����B�>�	�Q�㎔YmE7���s���8CO��3~�9lB"��奱z�ǯ�L��|}B8�D7௢�3r��4/��W^& �2�2'�hy|��.���gX��m��H�UE���Gmڙ��N�������\�GЍ���!��5�!��3�w�0���m��艆��טR����.�IEb�0�����!�J��\ޏ"�
|��N��eR�²ޜ�ea�s9��kH^+�N�'o�U���ۦ��eM/�����sm�b�73���Bs �}���_P:�&>^_�_�d�
�-���4R�$K���b��|�B2�"�F�w&��i<�Z�����e�+ð�)!��IDN^���<a71ؐG�	|�W1�Q����y?i����03D~]˻�Re��za�EA��]��te64�4 ��O�8�<kA2lO�"�s������$w4Ӵ���0�XD�U�H/�[���y��ꭝ�'cc��D�ϖ���[��q�[�\W<�7C���`�m�5�iN?�X��M�i���n�y֜�f����u�$�I��>�i����>��|��rLF�9�1��~�#�J���gJ֊?r���a�#�{�+����\|Z��Z�33��/�bm�jvi��]�?d	��и����'U�w��y%3p��6�ܤ�`IG��2�K�X&UP�y�4=�ʱ����E�P���Ҵ]���|3_����t�ry���6Һ����4�u�\=�
3��^6H:������S�#��lc�f��D�k~(e6�A^�Z�"8�/9f}1�lz�$z��Z]�Κ���%=��HBn^W<Z�k��a/�_J2K�	�@;x���%>4��ڙ��?�Y4*�fC��=�gFqH� Y���˺��-`�/x�����N����z��*T�B��^��C�"5O!��/LU�h���CͲ���V��������8^�SǻL��J�P�',6���&'����Z�X��\3+BB��&2&�T�
o�C���˒�v���j��e�v�V��A��M�''��{򝋇�z�Cwcq�Uo�L�)�i�dI�nMT� 5J�z�$]�]���X��<���A=ΝJ/��՚l�_�r�.i���DSNg2���/0�����g�e1�� ���V;5p�<��ؗ�:�7�w�Z�ԦŠ�[�f��|�t@�Z���RH�b��{\����������bߥM�� ����˟�@��$� X��4�bSUfv�g߱ ���������F�2�]�T4���;Dɞ�Y^r[+�
OU�Љ�BKR�;�cT�S�����g�T{E:�������KXߌ3���� �$Ȭd�S������w�e���R2�_|��	ŒO��uB)��ٓ��}�[��$�LM�ԊB���C9��3BSI�ep���K.^y鰠E-O�2�AU����&]��X!�>O6O�aHקP��z��*�T�>m(+�d�j�$�G����zW�,��s��K�:#��o	�s������f%e;���Z�O���$�,,TD��u.�Q'4�w[����h��%9S�&��L�tڅ��2WQ���;Qz���_k���!�{��������߃/��R��*� e��3�Yo��k~�OO�X�����5u����dÝ������2p� �
�#���y��y�^�ӑ��2l��D�!e�75�-�\y��`s�R��|��uM�#2�4�R8�)�UJP�5��aܽF�ԭy�*^\n
_���� V@H鯝��}B���n��?ױr��ct����48 ̼����RDY�P��#2��U�.P��qZ������� ��mK)��v�jB;[���+L�b�}��~��@��e���%O���o�?�2ڿ0=.y�%�]��^��j���'����R��}%0{�Y� T���ָ��]���t'�����{h������޹7��]Ю-�<7��a����9�g5�v�(7?L��?]�5.���B��)����v�d@'�Sb-��?E�̣��ÝA	R�:`�R�=p�D[�`�</��fvM�:��V���@�$e ��@o�������V�T�სU�ͯ1!��cx� �"s�Y��g\ef�5��n �2�&7��srȃٶFE-F*c�c���8X����i�k��α�&�Q���h�eN�MR�b��t/�j�`�R�E�P���jޛ�+�������ے*x��:7l����?m-��<C�\U����9�,�=��ʡҘǮUK�Fv���Հz�̮p�A��5Q2�>p@�`A�K
0� 2͐�5�-f
�a�#S\�����9��eN���`ʧ����������7l՛��/��V�����m�*4鄂9_�M�$�0��|�1�'Gl���,-������5�ْ�k,���+h�(b{9�f��z��ٝ�'H՛=5�g��`�@�0}���&���K�C{��O�/������I��(t`���;y� ����6�������� ���텭\��.s���O#Bg�]K�&�?k�o�m������S2�`�xwz��mm-�|�e���O�5��vވ���=�4�K�=L��O�%)��%�J�~���T��3t��Yc�|mr<)��m�����D��AV��R�>�����Rq;�� ���B��

���c�x��<4���ݚ(���X����M�Uu+Gsp��]N�!wA�?O��?HT��&<N1�Z�>��85�
Y�0�?C���7�sSkm��u���Զ�����j{ˎ�8:�0+ˊp=��X�w�9J��Vk�ҵzc$����Z���̳k�A��=~���"Ϣ
 p ���L�ͣ��9�����2�z��  �i�m8k��J�V��v�*N�\�E1��l���Ru�B��Rl��~�T|#/��\	�����ru4$)���wé����ZU�)�<w�Z�9kx�&�^LDr$�xw[��+�E̕�n�|�������8x|���tǟw�O��`��<����U&�(�gIcl��T��*�$��$�*Wp�]o0��[����((=Y)\���L����S�pJ�T� x�I����\�,iU�<X��|RB;��m6v��3�[XA����PtD��]i�(l����Q�m܏o���=*���Q�Ǵ���Q,C"g�z��qr�r,Uy�hE&Q�M�L���u��g�8l���<����N��3����Ι�Ө��d��@��WP�$���t9�q��3OBp'v�+ܚ�H��W���oy"C��.ם1t=�b{D�֒/S0���^�q���1����p���}��<��XOhP:�Q�(�3��-N݉��J�R�]�lF��ړ�(.y^��[�'�+�pE�v��|�t������(��lHr��s��#.+of���զ��������So�xv�F@ �g�3�c��W"  �+{h�n�Vǻ��9��.�$��� ��hf@vƟR@���G����'��ˑ𬂆��^R�l��4t�D�.��wG{���f۞�̰�>Z�y�0�6���x̃Sĝ0��PM؜�b��=+h�U!�:?�b�g'4i���0�oޥ =��	���p�&�p���������o�Ön�|�z/��������@H�O0^+�����Ա��Vj�ة�-����,!�ł���T��Y_/`����.8+�E�5�!�Pݟo�^�m�a�o��y���:F�ȲLG�-���u��tX��x�F�I��VV��� b`��z��Ҩ�%ռՏ������$}��J�¹��
U�����=o���u��i xU�K��r�۱ ���Ő ,a�7�5���yJ�V3aǚ�"6�Lo�׶;����K8��ED�6A�J�B���a�#fGu�TX��	G��׷ �hճ�Z���:��8�9�&i�����5�vg�,ؗ�=����&޿��\�\��=�0X{,X��Al;�
bJ@��7�D�W����:�&����������H���:���O�B���Go_.��|�m�Eն�縁G��l��[�j��� ��C6T� I�	'h4�n.�\�����u x��C�}���3�ü6�����r*I��^��\pݧ⩱�3�j�4<�'���o��i����yQi!��@���#�MUebܑ�	��Wc�d�Ki�"�*�7?��?X����_���T3�FM���8�"w�c\=���t��Wh0��K�G�M��'�2�m%�O���O��H�x"��-�d�uX�4�q*��H�R� �6"`ejdj�q�ʹtAmҀ,�������� p�*��}߽C�%N�C�SX���07�잦K�Yi,���+!�,~ޠ,���� p&��F��\;��&�P�E;@�$���
)��Пq�s�F6�L��];�!����}n ���ĘL��<�Y�,�5��%���/p�S���KS���NVy7�Z��lzK�\�0���P��g�)6�q`8�8�*�-��grDzT�[^�ߪ�����A�n���e0;v+�ċdUW���ݠ$^�>X�O)��{�ۿ��!�И���\�M+�/�E��W�~Ы���m���J�l.��;���	���8@PO����Wl�/xQ)����f�p�g��=I��9����3�����5g��2�p��1~O��J��KƮ��*_oY��AIN������kўڕ��T��_2'��P	�6��o�T�ӻl��]TD`�J�eIxU_@�*޼]K�fE��J�^�Z�8,|�����qq���{"�ˏfޜ���y��aÓP��uA�r]@�bo 37��k���ÇN���C��G��	%WL�W�Cey�l_��Y x���H�'�s�t�
����&���y{�yP�5Ԗ�N�p2t>�2P�!"�Dќ$l6�Wyz�
d�9/_�(:h��2�kw���U���y��3j�{��#L��xJ���7�y<�1��@��ٷ	μ���1�A °�
�#&cm��>?�����e��	:^9�~F�N>2sԣ����j�`�գ1f���W-EV}:��a�O�̌9d2OЯ��؟�~FM��o�Ʒ!�%'֖\[��f[+���:���8%���01ĆILw��Iݏt�����U ����{�?]�N�I4�Z���|�3r͝�����ܱ"л���B�X�'���V\cz�9*�?��p��q<[��ȍ���PB��*�8��*�����B����9�O��]5�?�e9���3��㛥 K��in#�{6r(�o?J U�҂�ns���M��Գ~(����ƶj��� b<���NGewagI&V+E^!,���߼+��s}��e'H�w�F:A4���N��Q~/�y׺V���hK#lJ�b�l���%;�L�h5C�xYժ���x��>�MB�f��QO���4M��Vh�A�7����:6����=��챰o75�F.�e@�i�k��eD���t�1������XC�s�'��7��!��귵��8s>lf��Rlngu%K�1=f�әס�d>ZE��ɫ��ww�k����;��v�И��2�&�$��!s����^ٿ��LxkZ%��SQͨ��K�
��9�����uQ��0V�.�� Cj��>t#��[;���w<Z�5)�/g �װG�$�!i;]Yˇ�"]ؿ����GÀ|�UQ�r�n��VV��$��f_��eqB��L�����E*������s-�-�fL{���y��}����3μ��`�j��Q�����C�g9I)�T�lN�%ங4'��V�������	��
y>(���<ڲ�UX�h���VL�7�6�~������N��/l����Y�Q�=!%|Ԏ}��\TkA�����S9�$�U�@���s�մw͗��?ݾ��lPY��K���I�)F��>D_��|������,��:���2!�)�L���^.l��4^��!��{��g7�+���6�j���>�^��E ��X��<��A �����H�&���]�C5`����%�D1���ƾ�!<�oM8��O�\��$NX{y�YTT�PTZ���Q�`�.䩠�U�;HVK)�����18OH.|F��CJ1>!1T܊p�	�@W��D��|\b�/�ߚ�7��oWs��a���@�[��(�lSNp�]1$�eZ�
\��,�o�*��w���䲳��sB�m�6��y~��E և����Z��%�N��G֪�3�H�C�Y�Gf��#�_���3!\#�ʉ�'g%q�x����ϓ��6����0OW�]���m��&;��eq�����r��I9��G	�xЖLx��� ȶ�Y�0]סּ��6:��@�����ߑ�O��g�����ǮMS-AK��E��7�K���"�&��\aZ}�$¡����
�K�2�0ʼ7���,ǀ&��F�s�?�f8r{�UP(���j�t�w|y@������C��/��5��C�����vtKϚ�����%#c��� C#����3��7��m-0e�f%,4���_n�*o����?ř344���Xw�湫��D�u�t�H u��+��E�")���
k�V���\O٦�|(��.��^i"kצ�DJ)���Wۂkf����7&���"N �(���:��pvo��P".!`\��v��.�Y�]�e��g�^��a�u奅A?gr|J˓�[<2�<�r~���~GC#i,���n,�J�v�2�7B��'a�1@s��ٻ�ᩜwZ+�l��$��(l�D�qAY�P�F;Y������_��;^+C���&˙�7���Uй��}�S��h�tw�� H';���#��j�O9z����*���=�����P	���d����Y���X���P������RP y�
���>������r%��j؜�Ox'`'SOkh�O颛`��|Q�e-1�Tj� v�,$�8 5]��͗�Z.�EGQ�e�S��0�E��4��������B7�M#f!'ze�of�3ad��#�'̚���@��gw��z�t�ѓ�4C�Hz���ׄ���K{&i�p�Pt8U��
A�]�����Ġ�jL��0{5�'�P>�0_���%`o�~9F���N����I�8��d��B_M�B��6ש����T����QG�3&n9V�gl�-��M�q��Pi�^�O�y���]�� ؙ�?��  ����~�	�k�Y|^Ey=I��M�����(���-���u�����:�}A�$	Q���L#R��ݟ>�k���c@d��.)j3ZC��l['
'k��ܛ��t��}!�ʼ98:�s3e�&��pA�o�Q[� ��J�'�/�@�)k���&��2r�x�����:R���c]�@"���r�R0G{�4
�ki��a�:4�x,��Zʍq��0��Ջ���.�N���>}�0z8�<լ��B�&S��2��`��W8�^�Я׫7���s�!�&~RG\Q�p��>���jNlm־<1O��a��x��GT��C����&S�X��_��G/ ��R�su2���p�IĬJ�ED�M߂;Uq!NU��<�bE"��;��q}v��qB�6`��T,�
|=	ё�f�������y��g˙�AN��7��V{�;��Y��fq>��u��߱p��T�6���1�\�O��ӌ�n�C]��_�Θ���M�[n	m*��r�f��Zx��n�_\��W�$e��/����ޢ9r��N������6�0�zH$1�\J)'�TN�tn	DoI�c��3��ţ ��ȎC�b�28�m�Y9�Z'�=kR�fHbFvơ%�{��B.Oj�*���Q��D��2eF�r ��L�|�Ȉ��*,?Ɋip%�ڔ]�Ab6�2��>�%�o���R��7�	�K��`,2ʡ��4��)�=X����Pӣ�#+��~�r�*P�LT�:3ԃgpi;�69kyߺ�?p�&T]uo�oD^.$�v�H��:��(U�G�i?0U�?�+Jh����0�m��R.�ݨ�,�ٷ�0�fM� �f�yr:I�N�'����K��r4�S���Z����H��BP�ؽ=�w+�m'��L���{%��]t��w��z�̻3=�~���F	�VC7w{������Dv�H��9���Y��$Y
��J!�rY�෍-y�� ���(��j��U�"%Ĺ"h�1ۋ��,?38��%�[C�W� ߸�e_�24R���LM�.@V�����'#��Fo�s�!�U�����@�v��Mvba��WGQ:�ĜI�/�q��A6���FNYx���`��.\����I�����C�$h5E?ժ�s����:�i��7�p*"�R�F@���<5� b�&4��UЏˉЍí� 4Kn2����	N'7�]V3ݶ�[>x;��9B,$RU[��Dw�4�������Ez8�J�oC��?�� ϋV�rr���@�RM��%�p=�骨���L�ɯ�$��ӂ7{۩��s�,�v�q(�E7EJF�[?�1IU�*hLd��[�D]j�Nԙ�;���s���ϖE�y��R��t?�NLA�Z��R8���V���C��3�h(xϡqɻ�%?��c�"�<���u�Y�>v@�n�J!���&}�0��ч��}����l�g)&n���~�7��	`;� g�|L��p�뎗=U�g��P&x�����0���%:�k��� h��,�[Gku:��~��,$+;��%|�������r�~
� Si�mO�Z#^����@.�` !GE}Xh![`���7W����Jl�z�%��{��� �,5��?o���b��Ľ�תj�^U�� ������Y���E{v�%�"�>K3q�<+%Hv�D�����M��S^��km��� Ff��_M{t��{�����s@)L�t1'���ud��e��
�=���Ɠ�4eX9�Ν{ц�,^�J��r��*��e�H�b��°e��s�f��m_��P��P�B��~C�����GO���6�MV���Sw~�N��{�4�@wK��z�ָ.�򚻑��#����i+^�;�26�f`j�j��&�����乿��Gn�"���AC�����ɻmq�蔡iI7���k�W-zj��_�*�y��
�_�QBG��m�ut��t�^+W@�s������i>�tm��\��:�[U�a��\��'h��H
�[ P�7�r�ɓ<��8�9J���PP�2���v���G�=	��&�Z؀Uk1�\�w���f)�a�k�x�(Gb4(�0;��K辿=ؼ�{��.Ո��R�fE��zQ��<ߍ�Q�� �i���CE��m��z��/�S9-�w��U�[:���j�m*��{��ǐ(1.!��rx�W�N��3��ڵ<{��ٮ��ܖ���jk^���ŕV^ �v���Y��໽��Y��@E%!�8}�)�͹�J�Wx@ˡ����g\��z�O�>��*��˵�p��.��ēaF\�@T�ϟ�F����>�ujh&����Ʃ������B�����h��n3��seٕ0���������i�E�Ixzq�W�_�!`�;C?0I���Je��>3��cw#�\e̒@�S�j��ԃ�����oz�ԒΡѳ�kr�w��'r��IӲh��>h��G�
o���́�=��"�� �f�|�R�����ܞ�����C�|Ә���j�)?����4��B�?��K)W�V�[���dJ͚r�������>>yk0�V��fU����L�Qt�SkX��������s���X�n
���
�g�2���!3=0���^	c��Y�ߒ	hP�����]�y��Ӂ4Z2���*�⏴8)���:Q�-�+E��^�}����/�l~��$����vzw4� ,�)t��?z�L>�66�����Td{;��#>N4�k���	���$%����C�q_����y��/�*OeR���S�[�&{S�.��Q
��sډ#P�v��|ѻ5�ZzXt/轧�.�2\�* m ���ğB�S�4쯁(��\�n��m�1���`j��mys?]������_��QTm��:������S�~�J�wQ�����ss���&�g�G��Sc�:k
��V �X�ٵ��&��G&�]���K��^Q��t5�ɑE?�v�坱��=���]��z�%�L7�1�aY��h��#0[O =����BJ�y�m+!�)��T�Z���'mކ:�)d��5껹3s[�x]:n��@�=��s�+J}� Mh�����:.���8eƀ!�@�n�=ˣ���dk�e��H- �(m ��vcTl@"�J75�<�ko���N3Q*yJ�$F�J^� �KM��r�<Q�t��x��kHx�3�E�K�qC���7�Έ�Й��[#dg�x�hUM:t��h�����N����K�2(���S�@���i#&1,�}�=4���1�"���"�-"� ���k5�8#�LW}ҿ�����H�GJ>�A���P8&L1�pi���Hd��`�)������bs盚V�����p��L!����h؊d05>���OM�+t*!?�6�X�>x�JA�,��쫮�R���3�{0�R���/�gA�j��ouF�cK2O=R�;~3����:ܹǏ?�HQ0}Su�(7�ٍZ��qM:�R�o_�L��~�JF�N��{z�����iU��^��L�����t�݄�YMd~cvj���B&���|�>1�z@$&���V�~ݝ#��SJ��!����.R7Z�����me�5�c��[փ�ޘs�He
/J?S��/��:�&^���Ή?�E�Q��L��I��'@#iz�����wWװ23z�����9�`Ҭu<��ǁ���{4Gz��m�۸W<��,q�/���͎�G��$٫��/������}��(���������~O����&۱p�e&���p�C�̊[�����Z-��ָY2� cS���.OU��b��>������_�Tr����`l�@_O���+pw4�_ �ƣ�S�g�,A�-���biF�>�'��(�	��p���O��'�E;N���O�]U���C����7s��&��M7T4�=��>a��51�� ���?����YF��M������N�P���±{zX	:�r0�F���1/l������jso�{@��R��aۑ���6�����d*�ܓ�	ujU�V�1����]�M�vҋ�G��b���R�yл@cK�����l6����̎�s*�g}�v���*�ܟ�z�տ*��܁���0*Sx�ѐ$�`����|	�~i��������w�=�]�{��{�v��@���-
�{L�7�x�~H�j!]1�j�1�Ã��)Nx�~Q5c�7S�D%?$G��"c��s���݈z�B�5�ц�-�V;�٢d��jaC	�x�m ���Xw;d璊��8( �t�g��(%��=x�=g#��[���:�[�|n�/�T��린;��]Ke;T�x��2��ޒ�:B�Hq� ��"��V�~�s->����r��!�T* �ӧ��� �!����ؐb�<��sz�Pg7��,�4���ׄ+����B:�z�,��E'��]�^�#�*�;)��N��m�ˤ�F�v����ng4e6�i�tɳ?��np*W1u��ǜ�#�ԫ
��D
���f��5oEUa��q�a�����2��H�y��Lg������p¼��u���*B�"K���O�Ɦ�&�G�tbA���^6�ZLuڢ[n0Z-biI����^V�Hm�r�P�;�N�d�ict6�����|l=�WX�8�+��r����D۱�k��s~	S��k�����F&��r�r�~��/{ٝ(���z���)DU���]#�I}T��n:Z�1[���S�Ҍ-jW=�v��oD�w.U�@��[%���X
� ��$���t+�2�Z��n�^���J[��i瘛�U� 1���\68.PC콳u:�3>�{Sia�� ��$�ޝ�C>#j��z8�i�S
�J"�cƣ>><Q��J�f�4�eb��\%\�
�r�� 4�ma�F�D���ڠL�3mKz�v$�8���Y���QJ�g8����Sc�n��Z���nEUKܥ,�+�'���Vs&怨~�%.Yě9���I���J�et7�-���J!~���5��Vr�g`��#g���ɑ��t8�Q�H^����A�;(���;G���C2�J�1{�H�R�t*�}�Q��"�屺n�ʸ\
�U�+�j�	��6q:�#��bFZ�p~Q@9�t�<���6�ew0���E�&�"�����7���`����a��M%D*Q6�q㾜��gb5���>Ov����e�e����!�[��X�_٨cԓ�pZj�4�[F� uIq?�=��\8��i3	`�V;C̆'o�{_��j!�^7HT����/�Ə�6�v�9&u&�f�'?&�8�i�{��I�JQC^��+)��S���Or����b�\�4R�q~4n~Hg(�
ms8�k��q}3��"�1܂~��ڸ�ÿd�]�˩��N��@ͭqm�u��E�d0�E�@�|fq��w��	�O�@{3o��;�;��n��.7}O�L�&')��az��D���9��u��4��43���>s��P���=�7h����}_Z�O���*�}k�x�������4��<������c kQHK>g:	u�,v�3��$�4���8�����(j%:C���?�JfI��to<;���O��.�c�@��扔ց..e��~0ux�	<�k���� o1�S$��{���i��%Ѹ�l����tz���$�� X�Wg�e���Y�.�Xd�=p��!��!DH����҂> m���e���ި$�T�����6���<	�}�]��L�P��V��UH�B���r���p��������.�l�Ͳ�&�QgDk��l�$�F��qG���r�`�>��'�t�1��_�lgL�ۉ>h>���e�_;�Hg0�����x1i')�����b��"f�������ֆ,�!*=�y�v�l3Ur�$�'1�D��uo`��EiC��U�l�U}B�Â����q�ʐ'_���Wi5�r�[��C��p=�Ӽ��ZGw���ä�V9j9�A�Q����l�V�w���X9�/n"<�'�e�|$��񫮒Bt�X�r���Q�8�7�Vh\Oomc�
�WWI��_G���=���7�]`��>ymԺnp=9}�
S2��w�@�n1�U+���6��bY����j��z�N�XA�	 Դ	�9��h�h-�ܶS��%�UK�(s���
���`ݷȺĊ�ř��X�^�K ��/~E���d����a�����gМ箯�5�e'�F�R
D�Ol��S>#m�F��9����w̽�$JҀ71��9��t�����O���dd��|8?8��t���y�{F����YV�F�_�����s*�u��X�)���nL�6X���O��>�弐��$���Q�b��.�v�����6p���N(֩���#�i`|8����įW�]�0�q_8�2��q�"�����4p
VRZ�q����&\٦���
�Q��H_��a%�W�l�"Z�\A�B��5�G_�PT9C�{e}�xw��o�ʹ���� ��
����;�wNUZ�I���󑝠�X�-���4�����R��Y Y��*ݎhEˑ'8wU�y ��z2ۅ�`%L���kV8� ��㑩��m�ഏW8��_{�`b���V�?�!���t�/�D�8��Y�a��S5����t|D�n��B��H�����L�~���g,例Т6W��{W�G�k�cF�K�y-�v��tC���xjf��*`��W������6�7y�wZ�䤝�Q��݆~�cD���}��[S���n��	��c��͉g�!�>0��k�*��o�f0����[K�=��Z�iN#��9��c��SV��]�(�Q�2��	Hh�_�Б�Y�28������ GF�w��G�Z9�|u��i��F��[��r:.e�Ř���;��/�7�~lJ-��?��!k;T@��
(��,���S�R���c≌��&�'�������R4���H �@�M2��I����sjS�B���<�X�/s84?Ke���y�m��������*3"1���B�F�:�^�/�v�~|8}�!Q<�/��ԅ ۶80/]�&�
S�}���J��$�(�,Q�r�6H.�HD��IL�8k�.崃�:�2Fl?!^�n[wi�d��jZ?�-w�'<�V�7R���W�F��i!1��i�E\�w\�|�`�^���w�N0�2?�g-;y������b��ˏ�p�V�O-��Jt|�Y��یη'�>?�h�8�~
`~J�u�91��A�h�����oNɷ]	�~(�c�y͓���9�/pߋ3L�ŖB�X`.Z�d�wcQʖ	���ؕ ||�CZ�;��WC�»�V�i�=�T��9tol~u{�)����N�/w�X8^��[���ᵇi����w�ܠ�,��v���eM��� �f�G�c%�c�ۂߙ��u��$�V��'K�Hl���ޒB#��1�@	�/;�O�u���u��g�;��Y���-r&juU2zIf���y*E�>F"�(���N���;�ny���A8�Rr��g�
\[ ��qì1�E��efOr5[�[6E:�<߼s�Z�o�B�����$�u'I��^�r����`x]zd�4+�ce1�=}yI�L������@�jڛ%��e�g��ʷ�<��_�c�gkS�C��ⴁ$|��rI�8��0�Z5��2]>��6/�Z�\ZQ��:�4�0r|Z��x&� eW,�q��oL�˥$��O��g�8+N��y��j�u6�H����P]�"Y�O�{��^ 
�&L��P���'g�rg%��9�@��^d�Wxj�̨EAG�#�9�[IUx?\d�݊�����CO<
m0I��:R ]����ig�B�G��tf��T�b��
,(aH@�D�	L<�Q�rw����ȑ����4��aY[:�wv�pZ�ۡ3Z,K�DK��-��ΪgA�.t���z�sQ����Xٓ|,7�0��;B\�BZ�5�e?��}�1�c؅:W#>d,�"P\DGc@xW)l���͋Z�����LT`�K2����͔���x��'h��?�[�&{�,��$P\l3��kSy����Q����Y���T��Ϧ$�r8���E�Qm<7�������9�5lM�i	E�%��h�8��S��Υ�v_����1s�=6�m�)_Ʀp���u6�Ty���q!�ُ~e�O�����׀���lG��ױ��=���`�($9��AqipQ�#ׁ�,q�p�)�Ip�mf3�x�������R���i�=*m$�����B b���!�"�ۡ۠+H��˯��ܾ8@"b�����&�i�a;"�S��;���y
H`���Dc}?��C+l.n���}�^����;O@���:���s�~�F��˳F���Wf�&��5$Pk�����F��R���~�uܑGr��'י���=�W���_&Y���LE��_;V�?�B�K��_4�i�w-�7�L)��Vc�6a�:�nU�j^&h��ڽ�x;׆Iu���x^��=��4m�sB�ֲ�Zq�.�^�M��R�J�����H��ưk>a�H�!�[Ȋ\)u������p���*Q>X�z4�1������e��;J6&Z͹�( ���Ƅ��K�
#� ��b�	{�� ����c��`r�1<<����3,�K���-�H�c%'���V"�X��I����n��I.7"sS�'&�%�[(��Yߌ�����G=,��×�ց�L��8��f��i韭>�ԮF�x7q�Q�0���6��,�"cb~\�OLEX ����S9PM�0�#���{�����_yUH
>�'�QH��'r%u����r#-  yiV�N���k��5�kr.ȱ��J�� �6]������+1L��'��E������eJg�D��,(��,v��,��vN`B��I��B=��e��n�n T��a3�0đ�;K{R�z�{�uTo��:[㄁���2`9��a�ܸ 
k�T'yU޶�����̒��)�mw=i�md�ȏ!	B�̛�7L�**�����7yMaw�X}��u�vf'zh��^�+I#�K�ɬ۫0��&dƧ�x����[kB�``����+J�OO�rf�=%�4���RLI{#�(l�u3�����j�����2����o��5�Vg�=����PT���>Ur7%I<8?1�h��
Y}}�K��X ���F&���9�����R��ꦏ`<pW	T�<��z��a")��Dt�s��z�����d��m��$�;�6�1�-���a [QPL���U�2(9���5���̎���v�G˦�G� F��'��΢5V��jbr�|	�3��e�E�M6�o���J�FDQH�ۣ���Ʌ	�����]?"������>G=Ң[I~�(������%��g���U������.��!����NrU8E>�53�U��.�]c��4� �s��KZC��m�a�����GdCU�b��_���7��l�j�C4܆�+8�
��@����r�6�	����w��d%ÆDD��u�n��Ofl���������Z�wink?Ѩ"����<�X"ց��w�x����dnW�k"u	�^s@#�����j�>�5F`:�rz���n[`f9 ]��I�$q�'yQ�L}a�;�Ƀ|���aR�9��И�#Z?%ʊ�S��"�c�M
mzP�m,��cW�����O�7���	*�5;X�[��9[Tnz8�kN���˵101�j�N�m"�>�E�$7A�U�b��ɟ��Ɛ+��Pg��_���a�,W
�X�B�U��*�?�Xl�7��S׿$�����PѨ_ص���QH��d�<�
qPQ�e[]��@� Oj=LIiL�VD�R�h:e��]f�(	V-qж���+��3ےV�oz����úʟF�6DDh$�p��oU���!�D�o<�N=��'�k�PZ�u��q�#5���`�í]�$��M���r�Tl{��~'�A��!���㍑�����)��~�a��ö��X|V4�1�¸]Pu+Yz�\w�M?��
���.��oT�je��A��q�5-�u9��3��p��k`�N�ʘz�&Y�Ӡ���%�b�5��7�b��6)�����yscLH�����S+t�lH��Q�-踲ڨ#�̣-����y^��¬�ސPդ+bJ�b��#L��#ٸ㙱��̶����q�GX���41�s�u@'���)@���ᰵ�B�9u���1颶�/�F�G���[6ϥm��_X�"��6R�xP���ǁHtc�\�;�^��gS���CJ�srct�G�R�F'�����j�;?��\�Y�F�,#����TB�S�Y��r�9D���&ȟf����/�#���=��=]��,`�A!P�t���i��E���]��X k��={Sep�h<قhЉ�I]��A�B�i�@���0
M��l��i9���Pb����,�	�;X��Jv��{"�O��U����d��z��7%�ǧL���*c���ĥ��Υ���OC�OAk���)�G����%�9M^n����PuG��,<l��l4��� �O��"n��>������ \Կt�1�;�ݴ	�
������d33waw�{���,wƨZe{��3^�MZ�{�C�W�[.�E�K���>'=*fHw���B۝�-{=U�;n�}a\��swx��24T����	���BHdL*Ü9Ww�Ha_} ��2>���y�t�ORF:�z�<���N�~�6~�n�-����Ns ,�WW���j��{�!ɴ��L�<.;	v�yl�\����`��=���*��[�ko.?�e	cD 穠>�%kY��ʸN�X����ͮx0���O��.�y���v��A���2��*5.�r5��WK'�Gmd��R��`q����*9�!d��[�:�Nt��CX�$���Z+��y}�W���S˪��/���5驭h�ɨ�X��bps�:bD�$�|��	�o�����]��w�O!gD8��܎&�ק)���_<�u
���]
,ضvY(R�]�G
��Q�[E�8^Զ7߸K�s7$T��&B���	Ly��T'kN�e���E<�hʤ������0�f�l o��sf$�[�e�ɣ��=�*	�Q��ߪ���f�~�J��+��0���ht���]�j����� �K����]�d��Qk���[��J9��hc��ז��/�n�2>)eh������.+����i�F�g����9a����1�����R^�D�:�_�8n"�T�X�/_%�YP5,(�\r���~,�RC���)�;L3�PY�F�^�j\G3-��ZR��h��F�t= _��"�0�]J���ǼqOEv8�Jtx��ꎐ4��X�q�Ò6'�gr��GgH1;����)L�K@��ZX�C�%H�sV�WeAbg��٧@�|?�ҶC\��xq��#O7D;����o:��v\Uȯ���7�]�É�9�O�+���'IA���hI|�9�@�J�B-�Hh���2��
~��QHvV�{(\p.�}�T������p�!�0[������M�Zi�c=��[� �{���hXv��е;�*��>��Ħ�cU�h`C��ϣ>D��)
�Ɉ ��������4��>����:�
wϚ��%�2h�ʳ���B�5�[���0����=�up�|�Aґ���H�xȣ�fWB�SE��Zw���IR�j�-zd�^�L�!���8�}�f=�*6�jo���b�²�)z�6TCn���N��]�'�N�!^�1�=p���F�A��{�T�rODY��9L1H<��I ��w$اUw�Α��n���q�y�D/�%�Q�y�0�i�N�,��S��5eO�Yi��BZ��Fk ,�u��mW&��|@���
f�j`���������_�����j(.�d�x$�81���-<�G���+H��r�P��aы\��LX'O	�	�̊���`k�
�p��*YL�l��`����?����	���0[B��ʃ�7wX�ޕ��*�!e�KG��4VS�m�[8wÐۂs��:V��:�}[�;މL-%�v��o�p�ͽ,�9��R���xjl�F)K�4��[�B����]n�B9d�ltlL���(@�}���*��>������b6|y�1/�5�F�16�x��aF�ѰZX[��d�ހ=�aM��m4���?�{�+�Y���_����A���@�,/+u]	At��˻ �آ�D���b���@�;b��2���4-�W:���(�f�r�
�!����N$����2ma ҶW������9�}��wԵ�c�Ѭi��	]~o��7g�Y7ݫ���ؠ[�
�7�k�����XY������z���-��_���v9P�5��r��]�2h�xF�DY�M,���!/��p g�^b���D�*�����vW�"x���^R���^���C���ܤ�݈*/��LN3�+�X)$h�{g̖�|]m�7��X;�2���`�u�9�Ϙ�|W���ۗ.�t��`5(k8k%*�új�ϬDO�c���O��3i�e*�P�ڕ8�C�89��۩�q~�⓷��SI�̒d��&���"�Ӛ�j�yǣ��8"�s�3��(��;n2���ks&�f\q�)\�&YC�_��0�e��k(p/M������d�9��Ԍ`�@{L�!��z��hYi{��ƙ�)G�L�iIW%ѥ���m�;�N��	��Y�W�;W�"O���.�Kw��q��{r邸,Y�//&�"Yx$��'��mk�l�B��g>�Ѿ�˚��݅����o��R��GN�ލX�z���%f$22h�,��>㢺�WgIE
���d[��$���vS]mx��j���Щv�[�*@�<�l��ز^���s��nb���n*�P5]z�]�մ�-��`	�����=^��&HkB�ώ�Jw�IY�ǰu4�dp��L��]�/�.�s���8��h��b}�ii+�]��2e���<}6���n �ζ�Z�.�VT��y��X1{f�~k���S�%ʵ%WF�x{��ҽ ��3����Vd��]q�|�_O�ˁ��<\��4�.����	���o�1V6Ǥ��]l�f%oZ�2��ȯ�ͨj�r�GM����c-=�|��Y�/�9�k'�D$�����ڈ�K������6��*&[�K���qz�6�&��$z��Ikȏ���5ʏ$�ߗ;�ச�V�8���B��0�|�<����*�ΉQ�~�� �K犎z�^�;!x���j�VC�2��~%��)�f*�7,צ#2@O3a���Gu�� �9������Zal�s�kA����Xc��ʑKIg������1J�?�Z�����1P�i@4����b@�'����*�@C�N�0��� �.v=P���v�'1%��������˽]/���`�¤`�AY���1K��F�{#���V�$.�43�PxǕ�_�KIh�3��F�����a��դ��"�i����2mp�7C�j�`���uL��J-&�N��r�-���/nMο�~�V,Ǌ֙A,5��`ov�y���Q���,�P�§b�iuG<��t-�ӿܺ�π�0L ��%F�\;q���K��*_-_DXeМ���Q���a�,�WKG���Y�<o�r}33��U�MpH����=�ݡ�?K#k<�Q�x�B���Q��>��LոfG�z�%��x!&�2d��0TE0c�]'�$S��)-��q��	Y���,e���/Dlc��$g?e�@�/�E�1�1Hr�&�ߧ$�*�T�1��s��G�h�t�n�۫z�Xr);��C	Ȭ'���sڶ��l.�Pv��rH��`��=O����N+�aB�%�f�v�ų��nT��Y�Z���Q巊WqDƓiӭTf��Y�D�KF����/��nм&v��l@��O�y'z�=fT`1�3���<8oh[v-�N��έ��ZN}��ݸ��0fV�Oק���;fB<2GV�'���Kv��W�D���(��V�K��̿Ԇ�Z�4��|���7�S�g�K��\d䘶g��8�I&]�ڴR��事��ݟ��^�4#���G���v�ez8?��
� ����Û�c�A����*�s�hT�]�Q�C2DnE�A���C���R�t�@�x�5Tt��.CٞG��1�Nt�]i7yI�������Ѵ���a-
����ǅ���gNe������
�����EW�ћu��P�)��53X�]N�!z��V@xz%����J��h��=Ea�c1)z{co�6�5�9C��=b@�8����?���z�@��(����Q��*���X]��-�[|��q�(��B('���yR֍5�ލ� ����P�*F����k�ǳ�6�z��b���w��.�Z�h����򆜖����/��ޯ+ �=����(���K�S"�'FJ�V$���C@}��'�8f��!,7b��C�3���8jDa6��ne��)����)-�rENiV���"���B���7�~^�Օq���,C��8�y?�SC�i�45!g�M�b����T���ǡ��C�?H����骹�(S�S�����(v
����~���!Z�a���~�x�BJdļ$s=Ն�I�у(v��΀H���MPO�@��)�"�'�S��!�*�������w0\�{oUDI9��ʆ{�Tf�H��S�9���͔��e#.nˋ����w;�u5m�������3<��� �`S�L+���o����h�]hՂ���:���� ���Q�9Mg0
���= ������7G��sۂyȉ�A^�p��Y���T2`0�b�}�f}a �f�ba�n��x�TR�&E8=٬ﭕ�L�oI��w=	1��lIB�.�4�9� �갸���4��1�릯��y���9k⚱��������C��lzg�8������2)F�FM0�8�O��NJ�Po^}󉸞S�"fH���}~��7��pn^�4WXY�+;�����y.utߒ�F��H�rd�X��R7�z���q�7���YWxt%Q��a���:~���}��Ϣ��AC�q9-\d�������"�<�#E���[ `� ��:\��loh͡���I&7�����Q�)��j�:k��zKF�`!ϕ��w�4��<�Ƌ���`���2���a_ӽ^:���3e"|z	�5����z����BP��xp!+}jK��㓮Au�w�du=��h���]ia���rM����s���U�����{��vq���7���j�/�{��]3�~�=�?ן�c�A_Eb�q�&"���fԐ�X��Bva�}�
!z$��3��$�����m|��"�xgMſ�ԕh)�b��|@Pf:\K�����4��dC���c��ZU�"�}b�1�#��l{�/�h��"�#����F��I����/�!9����L�G���������6�
ǜ�@�w�է�&Q� �:�m�P�3�fV ��F�~����d��t+}OUkf�H1�b����Ք��S\�
�w��U��td̙�9�m��o^��$��0?qH��+�����T���"xe�:�(f�n߾i�͡=�Fq8�ܣ4d{�%x1V�3�8t���d����ٝ�7Ȣ�
���\�����$���aj�.�D��(�9�T���@t���fum� ܫ���}�,0ڳc�8���{�J�s��S��۞���qCM�5r��������X�Y.�d�3 '_�0�HU�m����ߺ��vg1��mo� >mr�'���(ϭ��G��<��CP��%��b��2�f����X� [I�E�Ok	:�
n��*�R{�щԣd�������	��B�ľ�dP�2Պ�����	{�i&��c�և�׌�u�P�(�)橽1X����Fv�?�DmZ\��:�k �g6p0E����R�D��<�gs+9�`��D�ô�f�0X���N������no�e�-�ێ;uM�����j$��i�h�X$��^�_��[g����M�����bn6)���3w��Ǽ�'����\,	Қ6��ܛ�`��/�xjk��z0�7�|����2���V�O�CP ��#�{T�Nۆ=�*Er���j��[�(�-�/	ρ�ܷ�U��sn�����w@�|�@?�P�R���/g>���1�qk����i�s¢�B���ؓ���Ҙi�fR7�ON�V+#��ǃc��#ߋrB���v���ʨ��џR	f�����,nN�I��Q�I6�%b6�WC�螘�2{�i��%�O���s����oX�������|�	�r��)�������^�H��5N>���WԴ�n�>�Z���x\��i�}�)sp) �.V�*�	N�
K����B7����m_a�}^Mn#�F��yWn����:����*��v��NT[ޚb����kʻH
�ǀ}D/�B�����:(���k�%�ƒ�
��0�t/>�݁�΀^D�wE}��xF_��M�e<X;������˻/���q���[����l�\�XG�W����1���3
T�N,z���`��I� ���b@��A��髪��A��LaD�a�f�T��%�'���ܳkb�p$�F&-V���]C�u�>]�*�O������RP�I�,�M��X��h�XHk-����n�>Qn�m0� ��z��ΘP�m�U:"I}'�Ƃ�>j�N�
���e`I�yl�\�I��Hn����%���4w�*�a�۸�&�����UW��5��r����x.}1��.Id1���tH-ףW�������!��fr�~5��.^w�Y�N��8C����F�	S"����N-ي�b�W�U�e����n ��ژ�f��"(�e��z����c�i�㽀��8=l�)�A\r�~��˕����z�MƠ;��d���)c����HA��ow�mъ�/�vIy*�N� 80�ٿ��������#x"����wѐ"�T������� \J���M�5`?��zc'o�� ��V��c�-b��2"�FMᑍ>K�W�u�j��t^�0������^���"���^_m+�E֭�s���'PS�,�F\`�Cғ�\D�,q�8����X���`�>Pf���6y*�4 n�c��X����H��^9�e��~U��,��y*�-���o�����t��W1¾�yۮ��`�8�FE���E�x�9���5���_�h*��(��Cw�x�؜
 vӷ���\�qm��0)*��*��7�]QX�~2�	cU��C�tu�޽/��i�!�gs�_t��\rȬ@fV��Ʋ�w��;�0�"᪦�4��m�<p��9��@Ma�rlg�v��g/"��l�����]|M%p�E�w�w���xyq��WG�e�؈�j�o�����H�L�%$���C�-V���f���7�n�5�?�#��K���7^�W�ub�]Dm�0������8��� �#�'�b�iYt�����;P~�$�d�ɱm	�jo3�:��>�;[�4U��W�=�ߒI����P�c�#�kp#�DM5f\L�5�G{=̪�k�CW4K��{:j>Ȅ戈��=�JqA#~˗k��p�&�T�.t�\>a�!܄����n^xg��֚8c�k���(iJ��y���j=���wZ��8�=��D�n�g3��#u�G*L������D����*�������f�}�B.���s�n�<���]v�P���<H�epp!�uox�GdOT� ��l�dFt n<q�T��  .�q)W�?��f96VDD1��w���m��U�Q{mdD�h*��N(�W�M���Ԭ����P�{CS��T�폕|�	p�j��U�\d�:%�V��ur��L�(;�����]��%�O����G+�7�!P��J�(t��[Q
ؘ6��(2@���)��p���g��"�!Sø���K�Q+�ق0����� ��^]�?�-����T+O���;��R�{"d!3�f;�A�:���)=y�-k| �3�5����x��N��I�EB>��F1t����R|I���	2���/H��ٯ�*��2�"8I��(�wz�:��Lnj,7^���ܣ������j�k|��_�R>��wV���`�}�k5�\�Kf�>֝�/�j)&�+�Ke���F<�z�v��ʂGX��ξ��O�_2S�^5S�1��伽���FVD	ң��i�(��J,#_�[#�ׂUҰ��l�,0<t�T�6i\Y�R���)P�e8�)����/
>,��ѭV�1B�/g�l����p�54�,��5��P�Zj`Z/���|L���,0���*�X�x �+�����%�	>�� |��S(�j�J��r+�e��xeޯW�����z���ጁ������Q4<��Q�z
�z�V�����_��R��O���G�	�r���p*�ٓ�F�oiՂ'�X�F�cTa(s��kB����y���R�Pq���
K 9+�$���|�F�Q�n{�i(Xu��=/ }��_]�I��/�j61R�PO�lĚ���ϘD�1Ձ��_�;���-P7�H���S)���A�77JM�b�E��Af�J���(s93�e(�����T��M*����J���v�����q[��������Ƈ�c�Q�4�',�Ć|w�oIc��sI�	�o��j-�e�smMP@	��+n���*���ۗ�9�*!�և�ӸFp��w�~�ƛX{��r())1�wPh>ݑY�&�'X0A����-e�8ZrQ�ߗխؤct��QL��qu���� f�c��k���-D`R�㽲ٳ�Mg�JS��n��dN�*k��& ��uv�+���c�c�E�û��ڞ���r�����/]�T�D�����1�D����%޵H��b9�H�>}>��`�XXZ=��45��Y�FN�r��	[��	2�'�`��;�uͥ�A,��3Y�j ���T2�����E�� �T�H�3���w�^�q��@�(eƀ��� :H D�{��Y	��望�XMƔ_Ԯf�� ��CX{��#�hS8tԿ
K��t�`K8F��azw�&c�sm�S�%f�_dfz�
13����*���%��f�������tI�i�������J��+/r��A��V5Bg��
�� ���e��nF���y�n��>^�x���a��fI�L<���S�I�P|*`H��ɩ���@�E���B__�XƦ{LU��Zz\� ���-�{� h#@�G>Iѣ߸�\�$<�k�u̵��PXvedRPR��c��r�5bDj�9`��C�@�1��IK�֦���oMM�% i����]���h���:���zFb��.4sy5�i���9�������Oi��\�s��H���L&��+.��=��eΨ�k1UL����(�#��TTHNϰ�B9����\����� �g��T��@�vF���p�%&���-���`���穽M@��p�*9[6AE6�u��=#�\g`�n�d�V���ߐG����ɣ�� }s����1�������l�"�߈x#בå�5���z!�[���g+�Y����;�!��ls�Ps�X�(%����ø�R��)xX"=:�Z� $0S2��tA)��49/<u�6�E$dX42��~![�gv��ȑ>`��6Z�~دk�ꚭ��WLq?YN���?o ���"�R��7�u��Χ��vy��~w����H����tf��O�	]-���y��|��DyH����-J�l7���ѭ���\�ds���<����Y����j:�]��fY����1g3�ڏ7kÉz�-�.����5���P�oB_N{U��r6��[�����X�3���Z���k�8k\3�����1�X�c��;s#��ŝ���<�k9�H�|�q���䔇9�x����'o��2��N�%��\_L �x��}1z6�� _Ƕ��`����I:V�x�h���'�k�И���VQT�D&��FO 8��VD���/�A
�I�H�m�%5�����<�7rz�'!&P��!��P0��5I���,��G��;�U�^&q#u���5�J[͓����%Q ;��u���PUf��Гa� \�� k�G�w,�H��z�E��k`�W]=�������ܨh�|�р�x�n���M��7�5SM="���x��~#2�O�g�Z�MmM`��P�o:"���EgsM�s袡��r�Q=e쀷OCp���7@�4���3z�W��ر�Ө9o��D�6J(�	i�v��(�z�`r�����m�8Qt�-y�Ί��Q�:!#H`c:pN)���E��+0���A�`f�����F���	�Ă	�o�f������U��KҺ��<;1�����0b����'��;*��D��abA�����5�.�b�+������'�����l�hw��R������R8Τ��IZs�)[S��V�����j�1�$��ν���U�}�7���E�[S���:�a( ��������
�,!��
�K�fe>����T�6����h*ÝT�LG �?KqRt��������D"UlC�K�ֿ& W�i��\��J��xd6%�wM�
0�gS�"��H�Yɀ�p=��Ώ�N�<!Х�T1Z+��l�u��z)@���)��d�r�޷��~eht?�@�5zJgd�*�Qs�Ahk>pD�7�s8�;��!�t��#��=�ًK��P�V����nюM����!�ꑩ���0��>���M!�@x��8����_�=��7::r�X/��pX�[����6��y�@`:����m'0.�;�+o�fxD�>���%X�V
����5�ծ}�� ;�q,�,5��9�K>���NH�Q_h��+�"`	��-VS���p��*TDw�ؒ� ��c�2f�b�������\���$ξɩ�IO��Mx�L5$&�f�=J�NU���S�|5���g��.	I2�6=�����֊k)@ZQ
g���L��7.�h�a��'�;���/��.;w$�k�ŷ��W�D�v�\L�r��XJb(.6YЖ�S#��%:d�w#�+�iv|d �Ɣ�/ ��)zx=�%�:��=��<1R6���6u�|�p�2u�Y@I�zC��$�!}�r��X1������$�$�>)�iQ�¶���?GXD2As�sJ�QɂѺ���S�DB�y��O�Y����B۸��f��:�5l���H2=s=�:,��������ͷ/?71L�m�;�xmiù�"��sK�T���F�.T
�Ud+W�7�p�xЦE:
��S�$�nطӝ�>#w�O�=�J�M1ܾ�f"l)�n�]��_+��Zjn��p�R&��=�O�g�� ��7�4���u���T��܉Y�H�r��}�=�袢�.Jr[U�>U���X��$(J��g:a�=� �:\`�0��9*���Mzi������*����+�z=Zn4.��UI���!�U��9H�|�Z|r\%�&�����ǝO^ң����%��!��L^� ��M7����?yMnF��F;�TgLa>�?v*�u�*V3���݀�e����7Bo�*X@�����z�3�����}�U�wQ5`.�X/��]� }̳t�®�^\��j�K�)R��n�')����m���P|���iڑ��1Gl���Ga�I�R�~�1�֑��_!(�����L�#����C��R��;	��I��K�ߏr����l�F�wCQ�7�E�M1!]�іj>�^2��\c���{��7�I�,��`���8M"��҇a@��Y�u�kp,��� `	��7�^Jm�pT�%�%��)��5�*ކ�7�<tŽ:%TY��$J��4,��5��"�窽��a�wUs׋�@ѝ%�̹=�rL�$�S�5IV��嘇��.�]4��f}�-����kE`�B9����_/,r�=RZ_��V:ԏ�i$m��z��Pf��.�{ 6���[�zh�1�LV)�ܨtU�l��L��<C�BM�V{�hS-�q�*�1�\|���E�G}ߥOH`�2f�QJ���`cEL?�l gs7z'�>ϊ�6]ν�c]��[,��W*M��4%����xj�M��H ���3�D$#]}�|�E� N#�����E`��'�h�O�3@�]Y������֨����(Q�dvSe�P|X@�i]�b1�����H6�2$��E�~�u�`��U��W������,��ԫ��oiJ���2$eJ�FY ���G���O��&��Q 5�=Q����M��0�3w�ip�zƆ�R���������u	�+��!fM��=��7�
�%�R��7A�x�}���"c�}�,��39�O��~�! dB�W��"��B����T���8m��e1��)b�8�I۔h�J:��g��4�o�1Z-�����X8���*���+��O��¢
�7:�j���h�c׸��'r�z���?�ض�3cyB���%����7��cU��!�8��{���o�L/6�}��{O��f��Y�o�ʠ3���@�������Μ��ӗ�!=�b�ѳK��T2�6$!�[0�ה'���ʸlV�H~���k��2N��o������	qi����	3�������{��%�ˎ#a�}����*
�
�4	8�������oZ�L���`��R��>ň��Gq8�Mɛ�ְ>�Ns�lS��qG����J��ǈO�<_�����#�O��;z&�)���6`�+�c���7�K��;���]�zF'�DcmS��&�pM�j�����@�F�}(����u���j]���c��]ʚ&i�֒��UM����y*D�Q�W"�����c6�d"%�\h�ȝ��w.�J����W�����g�����,�g���%��nK:e�z�]	>��2%�gH��jꣽ,	���u4�C�Y�V�.��|P8.�{
i�ǭm���Df���V�J�V����hG�j ��̿i4��1-�D���d�?������N�SZY�;��6)��( ��mdyR���]�����<}�*�-����k�/�v�:Jg��*���0j���e	16����t���H+wtp�8�-�?���H-��\���)�rT��t��������.�����9����]@~�I�t�^�+
X<��ǿ�ǌX��Ə���Zq� ��|��F�=�I�0A����֥a�*<�1�z{��3�����5�E�K�4�)�V�Hձ�0�cV��Y_��bw;�u[R#�����@���Ӗ���ȷ�K�bQ/p�0^?�r�c��6��k"��V����ߟ`���TVd����E��k�������Y}Ɠ�ߖI�gT���#T���4^�L��)��ƭ!����SϦ�R|z���Y��>��.�)�����頹�`��'�[�F�-��Y1+��hz�6�N�F���b�8�F�D�A��@���AT���v�xV��d/L>�`��K��s��w3�ߍ/�����b��{z*����y[M��^�b	�k��vI�j]^ ��G�Q�z�d)��ԧAȣj�E�Bs��4{�����u'` ���3�5������s�L,�����V��HD��b��MhWsyhW`�"��96�4I@����n��i��/�#C��7�fETO�{G\t?�D>��7���ÃF��v�;�&�{E��P���*f���ߥ�(A`ɹ| ��A=Q]�2
������pK${ �ח|���o65KK�W�yJ�n1Ӌ�?j�����ਫF�����_��X�9����0��o
�t3B�Z/��8���,Ck���$&��|1^��'k��y����Hä2@�9����˔;[�$���̏) ��27�Q���M+t�Y!��-&R��@- �l܉f5��R��߲m����Z�D��o�H��-)�@�r�5��E�,�w�Jx�P��q��dm~�Nj9d���1����j��)�ȿ{�������V�!�Y�	�YISD-_ �P~����>�8����ITu��-Qɺ�zT).�Ђ��@��xc�ڕ4�b3 ��Y���m��!�~�O���R��SEe�CV��D=gvuA�] ��U��Tjw4f�lhY0̙wm��I��\M���¯��f���t�Pp���t��f��u���]��.�y,�76P�4G�lp�j���Y`�9�5q9k$ԏ�{{�H��W����۫�\ʖL�u�p��<�f=.B��"��
���
^-sf"v���1F��N���"��m��fE�၆Mگ�*�F�#Ӽx���������z��0��?{[����e�څ���$�\�yϛ:�/s��j����y}���d?��Q� ٶq(	G�`K�C��h{	����n��9X=�x,˞d+�9��&E�S5W�[��Rcd�1�H&Kxg ���ޢ�s�x�=�A�����/]Pm�9���Z}�	F�g}�%�r��<{�ʞRZ��}��`;%x�-$���Qޑ_ع�sD=�fc�
]�����n��vZ(��	/��L=���1�YCF�6�+����5��2y��P��N��|��聶��Ў�r��^���ө�zR�� ~@�����9=8���Un�����/��j���*�B�t��'g�l��� ܑ��C���؅+���A�N��m�[����o�Ǝ��+�J}5�a䂀�9�T��*�~�&!T�/Ҏ`E��$�����@j4P��Xȅ7ۻo$a%Z�.i���T��aX���hj�(��m[BQ9�۬E�[~����Vo�)����t9ۓ.ߴDS�����s�GHtXK���*�%H	R���9Q�9,8e�`�+1a=�>@{QO�Ĝ�Q5��.QB�BU?I�"�aE\���, )�i)»��Cټ�
z���oq�B������� �k�������>.3,x `�yJ��v7F��X`��n������V;
9� M�w�{ZmM��z����3��_��:`Z�vE6�L���YbTOz�S W�dm�kMzP��5<}!���Փ�;��`%~!S�Ԓ��u�#�ґ������G�ŗb85�
�ĉ3���!`��7��L-�o��k��^S����3�32�F(�87½�焓�R�o��85q	1����z��%������n���*1g�3J��n(���H������et6������Xq����o�<j�b1xn	�,�@��_��/Ik)����묙Q���u_�u�ʡNFi��E�]섭���r�,Y���1�Glu|J`�~���},I�A��l�X����A �%���|�tdR�����{�h��5�Q��'��z[PRE�M: �����u6���*���6�J���\�f����K�}�{�c��#�=�^D�_�uUgs8��F6�h��r��������6E`��1�z��M�Ы�yOIҩ$YEsy@�lt��e�}��ʥz&c��OY|0O��`�g�]LZ`�1��ԥ�B�slR��y�<[*P�K\��n���.�5\�?V�Q���h{3s�h�?��Ң�(�EAې:[k��lj���ҙ�aQ��Cޅ1�C����3vH�$����S�����=P!!o��~I�X
L�p�/ҿe*H�GC��P5j��C
Nb����Q+���ZO������0K�i�i3s��"CtZ/��*�����_�Vȴ����} �I�U��Q>�[-	�$q'��S� �y�Ðd���~�m�f�s��@U��-6�q&�	��e��VC�q{rO�f����"�sz��4'Z�\h$fy1a"��dx�ո:E�������YU���(�S��}hK)��;�%�0�X5�XئZ�h�0]�h�^.��-7���L�����\MqMst�I�Q�09} �l�=8T��)�Նm����F/)0�Jl4
�D,߶�y�"��YfRs��z#=��Y��DZ��
,N��ĕ2]Y	2(�i��������f
�qU8��)��4�"�?g�x
�\�>�5�� W���Lа����5��9	@�\I�;Ԃ�er�����X�r�PL�&w��4e��m��[;l�q5k�(xl����i�8��L_j<Kv�t� ��0�[H&���\&��Э��S��Fګ�����jk���|�'���� ���0V0-�Ts|�����:�����Jtg ��x8䀆���s��� h�q�l�aXM�]jl\
|�˼Yƫ�c��jT�f�����*���08=� N�1�7�r��+}�L}�~҇~x5��⢵��zL����~�v|\�����Ȳ4U�б�eK5��W0X��b�lN�9���54�u����plcU�Qb��;�!�ʡr���0M�N�1dڧKd{�:�3z��]BM�oĳ���]�
�����Ln )N��Ԛ�&:�g�V�Q���m �1�ְ�`��t	����hK�2'��8#�Z�Ց,o����\���Q�M��@�\j��q�Х��\>�j��ڎ��v)t����oB�q�m��|���e�HҀ�y�@�`���}�R�5�5�8q<3��l!fek�'"�(����\3���Aj^��D+��p5c�� ;Neߥ�vaĨ%�������8�-�����qűS]~!�(�����J�I���]H��m^cg"`���*[�a�J�KO=��uu�uL.&ݻ�o�� XRR�:"j�m�������@�$͓@�o�࿑�.�/zO61�O����ƕ	��9.kO� ��j������%)���t}���n�T��G���#ϫƮ�.��|qcG������H�R����K�/���JqRJgf��P��"�=�[���}�?�.BzP?Vϑg>�u!TݻoM�U ��᭠^�F�"Ctt␽'��+R`��yj��iv�X�����ڮ��&�Z�O��8�hD=NX��w�7�(�!Q�_��2���'\��ƀ�"U)��J�3l�/�4G���^I��[Y���~��Ƿ��W+�l�_(�~H_�y)x�zm�^�F��Еi��N#"�o��)%Ϗʄ�ܷ�Ɩp��9�@�T���t��F#��jx��sa�����85Q���ї{�qth���r7s�gI%��C`���g�u(KJ���i��&i��|ųj��5���iy���L�
q�B�&5�G�I�N9����s�gwOw�.���u4�Ԑ�*�8��I|˜j�zj�)��,骳�~�J����1�����l��̛����)|Dq�>-�S�B2�-��<(�շv�9D�u�%�ux���@���8Е�� ͆2Y������0���x�p��(9ұ�(�]r�Y��od�fˆ���!�����L��~�8�K;�#���,�������=8���,�t�8�d��+f.�ni�������~|Ѭ�_P=*5�(>�g��&~t��>� Yn��WJti�"٦Q}��&׊5��i=�����M����ַ��ۿ��H�O��\�۟��n�Ï�N�I��qTj�9��P$���զǗ�R���vd�����)�'�WT�ڛ��>	�O},4S����_2��)+��S�,:�N�U~�5�I�������3��,�U��aLH�L�wZ���τ��ɠw��O퀖�fJ+yյq��:��0�<�c�W��y{�X��)�Cw�����^6�������#+�"D<ٲvNgwc���4���O��E`���&cч�	0M��k*(��ڵn�˨��e���D5�.��H̒�ߔu���D�ّ7s?���yB	hyM�<�&���^WChp-0`�N�}S5S2�Կ{s��SgH�)%No�N��8Q@�Y�7��.��.�aMx*�=���4�#-���cc=�a��\37x4�w
���uoE�SV��d�Q&͈Ȟ��5��k=������2���5��kAUE_��P��`|����Vř�m&O�ZB
X�	~��<A��=ӛ�2��[C�kB��B��U�ڀV�_Ux�=��E�!��,�����|m%�溨�=V
��ߣz��9�G{gY�c���ş��d��r�i�$r.�ʒ�+륅
yu����sG-!#���k�~�JzO�|^�0e����"�B��*�]�$��w0��;A,�R�*��#+��wo\�8�6�)��N��S%�	�Wch��I.8^��;���+>���^��(7�̴�ZMy$�ƨyM(���8���_K鯠Ot0�}�,]h��z2��*�3�}�Q�@�'�QJ�?�I�#f�g�������\Ȩ�ء�Շ�l�pN��V�@����>��~=�� �?�s�
�N����&9�������4tc���2_CI=��]FC�//E�S=E���1l!��
��O�� ��;_!�yYs)''�x0C��2�u\����3l䁅,�v�+�	��2��Pqc��]�9k���]C΂�QF�:���pU�����cQB��Sh���4��#�[i��n����sTJrf��mc_�Da����#�׿�"Lk1�?�w���~<�pQ8Kۅ윟�<nn,��*iƾ��39��zc�lŷ������K���y^:�I�k�3��w�B�VG��UܙU�M=B8������oxgΉu!0�ea"��6\�����l/!�k�b�f��/\�5�|��4��/aa�K�:G��՛?ϣ�H�YE�I�I�4,�A��]����f��H�s�z��<��5G��\�,'�྿�F/�,{+.c�Q�lB�`�K���b(��(뱄��/b�j#�P�/Y�r5�Q�<s�j`t�B�_L�/�;���c��,�*�"����1�&�{Э~��[C��-K~❰$���z���9ٺ������`f��7!+&�u��,�m�s�$>� ����[�2[��vl��=���ý;�)��X�n5r��y(�����g�	Ǧ��I~���T�)SJ V	B�
C������K4k��[��g����B�$��Z�L\"]�О����u��2�,:N��^X2|�[ �j�T���Pa:
t����2�_2��4O�����:S�Z�"as��Q��F����x1nq���-�=,��)�~rq����G� �x���B��8�W/�Z��1,�L������8�,�W�Gc.�7�(�
�-h�X�ӫ��D�Nm�␜��/y;a��i	L���-s\���,ˤ�?�'R󘘍�A�w�*o=l��df�1r2<������:b{S�n���Q��LI���-���9��z��\4	��q͙)�J���j�@���*[�[m�iNQy	(�d�:x6�x)a�|�P������<�a�-���<�MT�E��p�7��	���4"ɚ��Ϳ��'��#
�ŊۦD@�'��r��^~k�;��$QH��N�=8`B�TOuQ�4a��3?�U����bI5w��G��1���w^$D�.���9^��h$��]*�$�%�=��ʹ#鬂���O�{���O���y��V��q_�0�X�R#ju~zi�G}�?\�~��5T��sS~�|g�!���ޕ+w�k�&��s���X�f(r����m|%)F���Aۮ���f��oF�Tm˄C�Rb°.�ցV#���6� ��g!��E��Ƚ��/�Q���X��	�^Y -�e����εDd�(�M{���~wF��¯6��ѥi�=sn��IO؈X�!'�ԧ+I���ݡ5Z�>�b����L�&�w�O�7
��{>%AzR!R ^��������z[�J��v<n���8���t�Jxh��/��<�oU]$���.<�����W���4@N7v�` �����1y��Do��L�K���k�*ҋ�p�N�
nW�-N;�����Z^?��u��j	�`�KHwB�I�	l�����P��x)���3��.�6A�]$eY������c�@�DNa���?��B��_M ������UL��z�7�²� e��B��}s2懗s�$��+wzp�we����]�;����W�ϟhu&�A�T�E"�"np7��z*�i���.�_�iIϏL����&E�5M��P�P1�����b�8�8L�w��9q�´&�s	Rn�a�Y@9�Q�ݓa���Ԝ��9��A�ȁ��VfSR�B�(�qP���:�������'4��k���`�G�U�Q�J�� PΔt�aP���Y1���K8�6dIQw��@܅T}L(�T���
/H���G'��J)�A���?D`�5]i�U�;�3�Z{W��.�"j�I�E�eZ�>Kq���mn�Z��{����ƾF1�0֮����u���]��	��Dw�5[��@9���zD�y|e�K�O�n�0�}�E�$������%
6n��匟�~�Sn)c���N*=f��z�(��p<�'N/�]��H�-��w�rk�Aj��@�^�3�B︟���g/�roy���a�̙$��}#�d�٧��.�S2�i����y+p{��j)�-O�u����-f��e*��ڬ�oT��נ�P���������5�=+��(��� �f�R�xd(M�>�Ch$���O�(���']��7�F�zj���E�͓�%�]A�P��;Ě�+��P��.⩘Ӈ(�po�Ō�M�'i�a���	��uC$jb܆E��~[J,��Y=z���AY�`����*h�\PK�Atځ	�C�.��M*�JX�?�C� ?>C3����Ϋ:���F�.mV�b@J��������� .�L��M9�l�<yI$aR����%������WY`�[2K�-��������KT-A[?���|l�]���E��y�}$~����R9܎��xJr�];P��'.л/n�w1{G�O�j�F%�{��;Q���'�ȀF(f��6�Cκu���N�4�<�`������+[��l�#o�yp���J��Xz{����5՗p�Y�H�d���W�?�]���5B�)؏ɖ8�F���V9�3�㟸�z.5���%��,8s=H��EХ9�1�׽F�<x�z����y=l���_�f2�e)��O�kJ���At]��)K^}r����l�5���1�8d�1'xM,���|0��Y���d�`��. �i���~\�x�1��NT���q�̭E�~�Ć(� r�x ���N�̆��~�Ιϻņ	���H�_O���!U�B����l���D�ml7����A`�>bt*�$�{�"śҔ_��ZVz@A��S�J34Wx�*���S�G��t6������/�nv�f3��I�3w5Ǒ̠�.~���b�t-n�6Z`jr��:��3>?F��%�~�w{��{2v!��^�iIӄ8��aUe�3���l���O�p���mD���0p+�k#�&�4�zOK�8����1I�_~W�LNf��Q��B��_刱Vi����ԭ�hU
-��p��ݰ�GLCk��.�~!�b?��)
��n\-����)-
X�@�o�u�������k�/:{�rΨ��.����X5-�r�n���t�3�H� Wp�6��1�&�M��6�x���K^�0�L���T?[M��1VXkֹ@��g6��@�A�?#������8�'v�4)��sBS9n'{��zV�t��%#�����=�qڄ&�3�Z��M�!�g����a%nM7P��#��zM$l;dA�p �P1B_d�ʨ�~Jy��Cv���G�M���~э��0��6����b�尰$о�N������Letĉ�5Y-܌��O��=lv��m�aށCMQD��z������xD�H}�Jm-�MS��橃?f)uV (�A�9#1F�hX��
q����S�~�s�>��T�W��rH�yٮ�� �=�sU�8��w$��i$�H� �(E�w@����G�Y��*/���zy#�o��F~>�]F.�Bm��%�]|u�J��J��{~Q~ȶ��q�g\�~o"��vT+7�Ю�r+1;E^�/�e)��eؽ�`�c&`��~z��(�!�pw�m�ޯ�����2��䤑�uFEWH4���5�,�� ��_B�Eb8f�yu��	_4	-�q્���mM�.�? ��Z��Js�Y�$���J3&&=��C��Y�Uu�V��-�8H6y:=�FY c�=����ˢU{���PB5�C�&JkҰ��.E&I����X�Q�p��a��j`�h�M�śo�o�\DҸ�j�C���a�rg�[�YN�u�����6�<�7a�갬�ǟ,Z�5]i��q(-����7J����O�'���O�m�@VA��T0$��y��ܒ���Ƀ�%��ݩ��4Ʉ����b�.r��o�E��.���@u�Ak��'S�>E��������"�ޝ�,��ہ͝9�C���f��2�!�Ѻk�U��'��-8��?r��0� �t�eկ'�CV�F�&GB�v5��;b�[~�	���c��e��Mxfn�c#EK��m#C�*���R�����Up�?do��������_�T�Z>�fZ�b�D�`$���ϽCތ��t��PԪY��~9^��)�O	B���)�v;�Z���˖���]&�\gl��_Wv�#>�h�Uk��0<��(�-�ʙ��ޖ"8�H�E�j ,b> ;�
NX��{����4�=�7Rю��T��� �24rԸTKPJ7���|l8^E�#��$��8���y�) �s/Z�=e����f�W��e�bPN���oW� ;�����'����Y����#=\�S��3�����Z �ti��WJ�^Z`��������@���嫌Ը���"�@hp~�/:P�N�:aF�N�(1�Ȋ8���w��KU�U�mK�Ո��t_s�,�r�7R��A�D�hz��Q���%������,��U�Y�4ϱ9Y2�dJ0<�?�3@�@>�(P��d%v�M�#2#���� qO�E*@��ç�p5�i�9"�~�T������9��J:H���On����L�̡��r����Z��?.pA����$ϵj/.�s�1��	��!6i_]�@��776��\�e�6x�ep��y�O��h7�@Qd�O\��@)s��C��ɏL�d�C�XiR�1������c�;���*��x&}��}o��qmw�o�	���B�kK�K�J�H�@`���5���o���ZYmv����=�m%��"I����3��J5���0��C�O OGgۜ����OH�a���ՐX���@��h �#�O�+^{%��O�ˍ��C!�8��L3 ��?g�5��Բ�<K���7\�o�<��5?�����~]CHW̯�͈>��֚��}�s�';&�7�3^�L�&:�������������Z��=��x7��y��a�N{��0�Ռ��>磿J>9!W���~�.�5 ����N9_�
�Dt�mw"�Ji���*�D��"f!�+L&�\��}ǲh�`��/���� �~��qٙ&�|�u=�����+�����)���<�(��q�0@ã�ϲ8lt�c��t'���R:u-itf�o,�6���̡]�ŝ�e�L���i�(�| ������~�İ��oh���1jOS�����kyZn�w���w
��}~��Ů�6�?δ?i�����\x>ma#�^�˟��h�RP|9,��:���Y�'�(�_K�Qr�{>J)�,��w���3;O���Ĉ��hU{���R���{h����7�WPxm'H4�3���� #���T�v-��f�0p���$��1{ϸt�W�DB��Tf�9��"L�=�rh����`o�Y)�t�?�+�w�/��I#̛B,�V�~TU�|�I���:��C��t�I\g+)����W��C#��,�j�v��G:� OPp3Z-h@��H�삊V�N̃W���м��q�нwMξ�S��x����cg=	�1D��sԿ,���;]G�ڋc�����ё�@�b5�H]9~�U#�l�R�G���n �"5ܑ��t:�*.>Cfe���i��Ƭ8kߏ�;PR�sh��P`��(bIe�H�:5�S<��x��)M�C/�<�룺(0{;o��Ǟ�"�ˁ�t��KV�I"��K�W�"� :?�4B�ۚr�(��P��ϕ���)u(#�ݻڿv�}l�7ָ�w,3z�t� ]~'���e�k�u��'�Sr��n
��_8�%�l��
p��G�M~^h�*R6�?����Nhl�h�"{ð��7��SNVĺ^Z"�!N䧴�l�y4#�Sǰ���/D�..��^I��v�{o�s1���`�uS2_C�gw�U��M�"��.��d��X_����N���V��S��#���x����9�vU咰�kcy�\jI�}�پi���(E�� ?�>}>f�FR��ō$��k���,~�k`Doo��+T��bKɐ�]�c]��Xy�C"�:V	�)[v��A����@&����W=l]+ha��Z0���+�05Փ$���A)J�$[��
�8bdD���7 �q��7A�ԗ���*X�������������SG�E��,P��v�Áϧ��4E�ò�M�]�)_N+� I���&��f�)w&��B���G9���~w����ǞW����T���J�8��YI;�$$L6���>�AL�~�)���^���5V�������)���sL��jW��B &�;�$V��@�~�/'7�Ɲ(��	���d6i �F�u�淘��o@�:��[6��
�J���;�+u��k�򇠚�W&���xkS�Z�	}~�Tע�Y�ۢL���⯡Ҷ�gi�b�-��=�:��9�2�	��X�pU��J�8n�1�I@�p���O��3R�Ȥ�a2ww��S��Z����y���L��<��L�r��o�!Gk쓁���a��dF�~��S9=��g�������l��0c���:�h�@��AL�I�
j�@�_5����Q���l��5�w�[�.Ɏ��O�;.tU(��w+=E']�h����W-�M�_��S�Jʔ��I#�tm��o�����O7��1J���vm!��p�IA}��;��������8�j��eK/X8L��&EY
�7��]Y5����X{n~�ኹ�����*��)���30C�Ňi`zUަ�C��}������i)��h��\N0i�����j�0��`u�7:9W�?Sfk'��!�J�*ہ�,��������4ф��RL���Ay𯱍���4k�M�w�7mv��Q�v@�VZ���&q|�'r�R�  �X�e�p������G�{����81��G�Оg�H�w�Ǝ����'��l\3Y�[3`�/ܴt��)�Fŵ���5���x���3�km+`�N e�p�9�U�Y\ ���x��}d���Wm7Ń���W��m��A�?��@�!b���ע*�\^h7�Qy���%Z��u�x]���(��a���j'�xM�N�B�1��'�I� �ؿ(��;��i�	�$��;{a��oɊ�4�6,������B��t�o� <�l��0 e���Iߩ�X|2�q���]��#�d4�TR���H�K)ȼL��1j'9ݖ��۶L޸E���b��RF~泗uw/D�L��Em�J���m� ɇ�T�8��^��9/�&A����~��CP��l����Ѽ4yC*�&�@�(��F`-���	�� �Sq��e?�i�Q�j@����9cD�t�~��Ε?���;��Mg�/�pvr��8�1�]�p���h�̷��W؉ʒ�T�J��<R�M<߾5Í�q��/�Nب�VU�P�s��fWG�,A��tx�X"%�k��� a�dϒi!��4���G�f�7��`w_=چ2���b��;�B_���b�jB��iV�A�"᯲��)��˹�|9�)X/fB<"�_��I3l�q�k������oC�r��(^�[�S�>��㮘���\1{���;������ŭ��R-�FVibi�W"��z���3��A��]�i?����7���(�=��Nnp����O!1�9ޅ�K;4'pbe����rr�\�U�ZyI�"��:�<��"����Tй�%�����.j�@�w����hc�s�h<�|�D
�1 `��|�r�G*gx�L����$�3�����oK��igW�n�!"	=9�}���۲>���9�Z�H�:����V޳؞�+h�B����Z|��Z|��AxT��X���p�}�0K��Ny���ӈe5��' l�W($�f��ݠ�PAVR�pzq�����ܠ8�b-S�ޟ�VYc�].�A�Di�Ii�;ާ]z�[m���0L�"h住Ȭ���9Q�7N@�����r�TQ�.�!Y���d0l�]ՄPU�3�
e���%y��{��)����`��"nV!��_��cd������~Z��!�>x5x����q��at�^L,���D��m�g^`�$N��b�n �ŵ�5uO�vz���Ϩ>!V,�G�}��x�i�2�Y��2�j�ϓ e%b7*��){������ ���M(�-��E���_""#p���G��sS�Y�{�I!j8�ˍ�aI*3�&S�B��"�'�P��]z��+Cl2܅��=m���%����ɇ ���Pq�Ri����X$>�?�����~C �)؈������[�^���gSI�2���$[�8:�ű�5��w��Ed��Kʵ�	�x�9���rm�xX�#�:5:��i��^�A�_������n�l#�H����f~93� \y�e��u��V*�b�]����>�bJ�<Fb����B�E���Gycb7���ܨ�����Z���6���_���c��Q��v�_�NI6(�5������~&�th#o��~��_��:�K�k.�W�ԗ�����x�N$h��fD�����!ތ
���}6�P/���_i�M�M����s>����B�.�U��s�� ���pZ^o�G�^;F݁$�g��#�@j皺B[3��T_Ë/'2',"HP�-�+bv����a'��Rs�p4�������_!i�,[��`k��|& 5ʄ�����H�ǭpg�uH�8Z����l%��FW�8CC�����
WY]i*�� 5��ʶ��j��e��ݏ;&�/�;��xD����C�5�>��Ԯ��4&��X�����4�6���w/Y�G��П���	E���jKE��6�8\2�$)M�Pgڲo�rc�;��a!ԙh�9Ba�??��&��_����Ҙf���p7�n55�9K
�O(N,�*�Z&�;�n �ʿǈ$�ے�\�K�&��� ڊtt���e��i���`�lUɄ�U��|�k�^��Q�Y�֬,�)�2��PZ�e4A�������1\�.
(�s)D�u<�N��aqOp�!�9��k|N{�TEx�M��U���N=�ϋ�{�i����z�Mp�����ӆ,��S��NХ�ZD�YM���gm��Agڀ��ꁨ=@�C�2s��T]� ��nS����ౙ�h��+���z]D�j�.͍݇	wO2
/��jH]�O0�\����k�W ���Qa�Ƶ���f'/���;ϛk ���V�]観F�ln�v~�E�k�_����C����v	=Tk)�ցai��z/�Y�8��k?�HQ��F��h��z4i-m�8�/O-Fӝ.6%�vd�M�t��(ɪe�< $P�V�[~���k�fM�Z����2��D�)tݳ���?[�d5gܶӆ�O�+�*�T������2E�5)�Wb]����	�D�5���ֳ�����ꐓ��R�ՀB�)`PqWr^D֙	^آ������Fdt�(
�I1�7FB�F�ӟ�,@j��1@�4���Ŋ":s�N�g��I�S�(01EhX�����تc%7�{�?4�}5(�����_�(��=N:�r��Vؚꗭ� �����s��?���F(��H��������{��]��P�.M���x�Vai��?|�Ħ?��r����fa�bFHzh���E�"R�̓@������|Ʊ��)H��� ���M;��~dQ���<K�&���(T��q������.��r̓|�|�u7��)�w}(Ӿ��U�[> 8��ԈX?����Q�`HǿwO�?^���=�Ց(ġ2#�J4��r�3�S�?����M���عv��V�nUxg��)�s݀1"I+��?��1���GH�Z�k.�8�ճ-WY��CxE/E؊�~�C���V�G�>��*'Zl<5��`U/��|>�Nn���P�\��kK#�i�D����&�p��
����W��G{���R��jڱ�J�Vrqr�I��;��k�坟�hqϴEI���^� ;";�J�A�*kv��p|^nۆ�]�}7�7Ɩq@.Ӏ��fK� #��n�:�q��d����/� Rm���W�p6<D���uɸN>�Q�0t�+�8���l~]\�/~ǻvY� 8KZr��Q������Pvg&���F<d 6MEx�"�\��?2:�]�K]H����J7/i%H��J��D���qk�"x��`�z.sh�\��HQc���&�_fKwČb9p�MD��w���4��,�GײO:�����J�HZ��;��d���ް�`�	����n"RIp6��1.\6bh%�)��/��}R�ِyI��[�}np�c7�gKm�����R9�>;E?������0���k�2>�z���.�0E	L��屢Sg��|���xHfRW_��R�����ؖ5;���y�P��,[�7�A�!�"LYdb/���籄qmsZ4nX@ �Uf��W��
�L�(L��@���V�(�¬�mh�'x-jD��~ד<<&�B����	O����F�#Kk��  �ev��s�ݖr�%א>Ӹ�����_�Xp�	�#�!���py�	�m��QD�\��^[�C?�����G�e�)��tO���ܸ�QD(�>�������.됅+���ɵ�6�Ǝ����կ�:�MS�K�p��>�g�=�02t�t�r`/��0�7��FG���ײI��4q��x� �g��,Ŀ@����&�<�F����'���������
X��%�/blt#��L\���lN��%���J�(��:�Zq^"��P$��͈�B���?=_ @�r4����d�/.�ߍ@l�q�u�1��/��x9W�TW�<�3!ꕊFa7�D�~�r!k�H�������c'o�ih�l��_�Zfы>`���M�@"J�+���)��K@����x��m
��5�}��>G����.�%����/ɝ���xs
��֨t?#�Y�U�$}A��o��
�%�Ȁfwm��m���|c��0 -��ꋢ�@<� m��O��e`D����G���MC�zH���k�R�j3�����%m���`�ʖ4Zwk.�6��"<�:R; %�Eg$_]��S�|�n�1	^dq~@�T���u�$&<��~�_f&��_�l�uR`B��I&�<�l�N��E�_D���q�����8IC��	�y��%*��G>+e�a�2<t�`�O�(Q�Ē�x98���$É�7��K���9���?^n.xm/����̩�H�䃐�Y^���q@�Le�\�%�*U獫8,�b�����V�@��þ/Ɵ��ɭT����˝��b8~�a>`�)�?��6&챡{��L֏ 8d��}-'���$d��\�ov^�h���K��0�>9���H�/`OZ}����J��3�Pڐ����"eQ)�V[E:�5Q�dM�_�����K��U3;�銂f�I���7��P�:2&�Ni�W�Z�Zr`�3�;r���C�gU�@+{P��uE{����Z�ֈj9��-�g�~���JW>(#�]"��n����g�e�:�h�q�殾���5����z%\�(�x�Ց�z���vy5�T��98�+"��&���e$���ʖ�cMoC�1��液?��0�������!F��]��F��˘aDY+�k��r�i�>�C=�Fo��t��tpxv���N��UM>�@�GEa����>P*���1\������cB=eB��=�t���q-ǥ
�S�h�l) R��1ޕ�U��`��07⠀�du��	�q�$�t�L�"�D�� ���~6��d����V��PZ�o�h 6u5뷒]�&�Y0���I��*�vAOՑ�E�=����iw�С�l7'����"�~�	'dG��1��p�T�B�̅��:���,<���֖ڤ*�+�>ؽ8��!���6�^
	��#�)yY�G;'�W�n�K�s�B �2���K�+��1$���&\>	6��XY2��2k�Ev9�k�:i�����ƴO����dP���U��Ce�w�v��*=�)j���}���u�ႬJi+�{�L�� ��?|	�e��c�!�5�\?>F��;Q��,�j7�D;��|��i���*H����$��AL�-|_��O�Zf$��F�����J���FXP%nA�.�)#
�擪`4㙸c3����ť�W��}�35l#>gK~ͯ���M�$����꿝:��;ayb{�fL͖��;��c�{�7�||��o1-�D��E�h�٭�����d*8Rm���M0���r��KV`N�:N(�Q�����$(f;��@	����C�{(޷o�w�0��aA-Ϯ�C�oʴ�eFQɀ~��������6�b����6E�ް�y:�#$aH����O$Q�&��Ȩ=.�s��vPX	��#'�[t/��붰���j�Q꽳�ڠx�tX���Ĳg'.��*=H�{�XMQ8Q���<d��|��Z٩ߘh4��V���r�B6b	,���I���H�u�J���Ӭ����ǻom`��]�.ݞ����Q�G"8�\�H(m<z.�{E�_��NZ�� �=�I
@�~jUA�c�0
�"�KG��mԩ�3�~�;�)�sI�˱�B�S�m"*��k�z�q�BG���m����o�N� �4Ƀ��-sg��e�@�jY)����PL$e����(Ii*��1��;5�ah�4e�zU],����9�)�,U��-�s�x�B���_L�J��́��i2h��8�HGY"�U�:��g���2hhyԘ��S�njb\}���2���.n��J���$���Pcν��@s�.6^�I�x)�R��4�Le�$	j����M�Yy���qͰ����
(��K�����/F)�3;e��\������TRY@�߻�g�|�jxkd��;S:t��Q�v�͏�pk�#�%�}�LɅK�`#,O��E��<��5b��p��jb�|��)���_Fŀn�	�`������{7��N��ʗq`hw@=;w�m�K�@���z�ب��^����lH��~�L�����X%[�$��*��7��>�xHFS�_���7w��<�
j�,ך�����Z�\Bip��3/��?��`�R�O�I��=KΊ��c��K�s]��kW��I��; ����Ϻ��e1��
��I�ᕶ�w���]����us;_��sU���7��w3�`��߶��rlaX�f��U?u���a�����TҊY� b^����h<����{k�Z����������	U|�
`�+� 8ś���܋��GW�݄fV�˪^X����~ts,D��kQ�� ����@[�H��;�b�GE���]�g�3�� E��,nN֯o����@6>ςS��	�/�� ��|�Lg��7�g3\)��H��)�O��$��7��xv	��#��7ۡ0*�Q�s��*UW���?�R�Ǫb�� >Ř7�3V�]��fE�G��.�{�7�ſ����N����$��E�h���#Q��:���������������U�o�%9S����ٿ�>�[c$�R�?嗢��/+�:T��Zx�������|.C�z��S��0��r��{�}8#���~��⩸Ek���HR�n�Q-�\��CY���6�.g6��
*J��~�~�$/�d��������E.D�!i�Q����FL��>y����"���)�_�rL;������r������4���}�'���T�0��E���-�S�鐔�G�5��nH.vf�����ۦH(O�
�<��ޮ&��A~��t����D��˫g��ԕD������<^[���n%��"㍾���_�Q�^�pK*u-�P�]Ɓ�Ş�D� �|�Gqy^C�?_��H#�1g��ꜚ���f���ž��D'�Ǟ)╊ ������+L�]N���h�Ɩ�x��{	,}��uGx䴇���sJ���ڌMd�͏4���Y�����ˮI��S��.������* k���:T��#���2�٦�]Y.��$a�4�ΰ�.��9L�N�Js��rp*���z���/����&o���eN�L����F�Zj��w�6���|��.�����"�?�V��HƉ��(`.�9��D^A�ԯ��I�� H��,�z� ���H`}DiI:@ؠq�n�*"2f"�˓{{֐�D���Ւ����T��iVPe��j��b(�m�����MZ�2�/`G��^���*��ټ��+��<u
��Y�>�V=eϚ��K)�R�E���e� �v|��M���9��h�3���y���k�J���^Ƭ�Y��v�e�X��H���쮫�I��a��S<+U�x��h>�F`�T!��rJkP��l�OB��+�./֚�4���8RrtW���$C�S�ް8*�G�Gz�D���œ��>{L��>/��'a|�oY��}]ow�e�$�e�M&Ȳ��1'�5ַ���S 9�[a��'���woIm�Sc��JA	+n�~����?0��he�]U}��|��C`��u����R]��4M�dO�پp�	b}���t�[��9��
j�r��0�~R"�mXi�\=�CP�<���ͅ�0���Y��p0���$�'!Z2!#s?G$�=����#p�sd�?=�R|@N�+�i��̡�u�̵CTn	zQ�U���r�~��I�s�?+LR9��k�?��RGk
�	CN!��	��u+K�15��;;���9�G�UN�[;�\�*�9{��U�/�F�{�~�σ|�թn����n�;.1Jf�P�8�ª��[|�)��{xZ������25;�	׍��m�tMBf��K�lioF[��T7l`���?|Ӂ�~���r�J�=Y��#9����*�7�/,�+���ٱyϟ����8��p��*׍B�n=��9��8aIr�%�Z� 9	v���,o�q�R�gT"&���+����T�C�O�)�Pu`��O�(��z�l,�U|��h�0ޚ�W���=��n����yg����Z��Ԁml[���>�ku���B[��S��%q��NSL^ض��\��Hg�G��������P�X	���S���L��s�A�^a��R2KBP���d,`0y��I�A�u��VG�I����y�\���ܝ����������j�FQI����9���ﰡ2��e�|�ǥ�_�<WC�(!�O�2_M�]��f'�֝�?! �`F�cN�z�f!2�6>�-��V�2N���=`���pp����F0��-��k���HC�טzy�v(�GCF�7@+b��_E٫#vN�	p�q���9��9�N����ƾ�� ��+^���@� �2n�#~���ǅ�٦;az
��C���xQ�� ��-DWc���M����¦�'��A"�����.~=G�h`����6�K�a�g���k�?]O-"U0��,.��F� ��&��r0B�k�V�N�Re�_XVX��]!��zc�Z��H�%ug��q��g7��e���V/o�z��L$���.;��06v�JBX�0aC�{3�++;Qb��Y5߭�r�0�V`��^�}V��,���n�	ZX����R�3�ORU�Z��S,P��"��`��Iv���{7�^��?�K��%uv+	�E���Ȇ5g-֮P���"�;gͻ�sl�w����k����P �[�����ݰ�J-h���$6�����l�yL{��Ɏ� D�=�ꔩϭ�) +v_#�� �+��5�?���dY�k��&�7�2��L�y���7����k�����5{u���8.8���F��y��9[`�Z՟$����D��ݧ5cp&�F�~���l}��m��|*.���d��$#ݫ��Z2��������M��m�r7�)|�<�H��;xL��|��5U0A��S���J�5���o�c��F0�"  �\Q�^81�����'��~��谟#�qi��f����u����4~�h9B�-w�G�����m�_t9,"5끩R��P��$BAh�u#O��PLc!���xY�����8�)x�0Mq}Yө��]�2��[�r���sɒ��5J��������pp����#]O9�K-1}Tq�-&N����(���3[iW%��bV��71±*W
��"��	����jL�B�@x�L���{+���&ܰ*Di�������?K.�Z�?�h��.6��b�	�--�_�W������C�����6�dw�R��m/]�Џa��P��X�QI�ci.���Z�E�Ɍq/OQ�+�*+\azڡ�3�k��#B'�ݹ�Fg:���;���K�"�5�p��4'�?VO��EN��`Z�����q�U�q�c�Bp�����E��=�=���LN3��'��N(�5��q�Hq���u4�c:Y�p0oʽH7��x���C���R6$��`_�,��J*=���[���s�L"G�	 ~�D���%a'p)��"�r�����7 s	�[����L�j�;$�\+� s	��� z ��S�w+W�G�&=���f�˻*%���p���}*u�pUA�j�<��A���5�m/���҈),9�Am��&�I;8揕�h/T"0s��~�����7fR5I��[3
wT�9w�C<�ݕ�Wk&a�b�Eb���w��X̪ǰ�5sJ��s�D���Tc�g���~9?\B�Sm>�������
ҿ����c��-�o�r��̖����C6H<��ź�iGdw~����!;s�Ƿ���e�wOV�&Ӭk��~.�%7��R����VY�� #���7=\(��%�>N"İ0�;5y�b���[s�w�
�����:(�s���$��x#c����Q6k���D���AH�b,�B%�i���WU$!礸\{� ��ʴ75�tkM2{�h�At� �c��MaMwW��.6�a$T2h�r�D��?��G�� lD@U.��h�`k1_ݭ��ka}��ǝ�0�(�4�]7�h�k�W�G�n�;��֡Z#ʐ��81��}#�P�$�5j���"�ӽ��*�Hd;���x&�|*>�e������uG�+��u���_�H��Ց/=��ISY��^H_昖LM|Ux@Ā0N�u���A�յ v�d6������<��ly���س��e+�� ��(x��FKH�0�j�tm�Y��X�^�Ǩ(��;z/�2ؑ7�HF����C%n+rx&�=���s�u-����3�R՞��i��ƃ1|Rv<�/,��3��sU�}PS)/�ؐo@ �A�ZW�Ԏa�d�%#a�LD~�J��[w�����;f����̹�.�yu�r�s�]
^�/3ri�\!��m��@:�PE���	��5W��;U=�"�OL�Gt}�]�Q�	M-���޵���8�^��[����ʆ�A�:� ��:1�3�$'�)BXDzYT��b^67E��K�
���E�{��㟍����e�n|_F���"Ʃ<i���7aBs��49e����2��
UD�|#�殮&Fr!��ArY7�H8�%-˧���[���Ig�j��3��z����0�:��,�ݬ�8F�������U�Ӵ��.�S�WZHF
[������^99��?�xmbK�F���Sa�Rt��qS�pb��q�M�a�ڻ9��JS� ���l���Q?��,P#ր�Qv�
N��wG Kd햢�V�����gf�Wl��~��ݷ{C���8� ��v�Np�|ЬR��S�"L�~7�f����uKF�2��2\ЙW����FB��u?w؄Prm�	�ɘ�>�ts�F�ٸ�A�m�%\�.:p��#ٖz]���ΌXPR˪�?��*��XX�AAk9�����aSe��`���

��#���g���km����5\-2,́��1�X���sxT��U��4��N��f��K*�ݶZ�5��W�ƛ̇/�y�ԖY�Wz���j>���t��(�?����7�O��"�3�#
�f���]"AI�}���tp�p�}Y��;�����J3gyB��>�Є���@4���̐�5����GmO ��)	�%c-���c!2ϲY�|��Y�H~�mQ��q�]v%�a/޸ ]rdC���E��!.!_<\ߙ�#)��DX(�S��:g�Hg|[�7�+9�0܋I����|�א���z�g�Ɂ�g�����?�D+�j5�@�?N2	H���Ň�l4�O�E�6=��#G�g�zf�ފ��}G<!���zͽ�2��^�9��������-��|�I�F�9E��n���O�*&��Zr5�'�8�3B�j�Jz�#���������g����qk�Sd�-r���h����؎��{�<���$<����B_��,
��O�9�hx=��f���r;�.�i?D�YJ��~_dAs/j�G�x������O�=V=�7��`R�u">6v�o�ĕSi3肐�jQIH�b^�^��Ú�Re�~��͐t:�� 5l��Ѷ���r+�>��.�O�����Ьd�_Qy�-�bu����e�k�xq��)��x���H0��q���s_�E�#�_l�˹�o�Œ�,q�����V�F�C47.��'���o�����6;M'c�/A�g k�daJ1q�ڕ
���0S��*� �mx?]WՓ�|&���A]��s�CV����TLC �L�i�)V���0l���Ƶ�0�@8��Լ@�.�9
ъiˬt��q���I�\5�1���c�B�8�"�n�e�Ч�ќ�H�8���ЧbG�&I�s�J���Sne؆5c�lB�T��Y"+}��%q�Q�f\��E�NY�.V�H~npxVYw[�c	`�i����)
+�CgU~io[�$3nWSU��_�2��^T� ��uw!^Ai!T��*h��N6CAӤ�Y��h��S7$��i��Ǽ�[2�&��'[w�^�IlJ�yߝ�tKn����j�lkх�ҫH'�*�d YrЖ�^/�׎^e9�6��P@�U�S\ב���Ԡޞ�%�)N��*(`�O�s��!v5`u}!�U5���QW?�[��܁��c��U�{�:�?�����C+x��}e��vx�V,99@u \f��>� �~2)���=_�^����͖[G��4Ҋ�;��=��Y�&�ũ���J�=e�p�tUsW�o�/�?l�u^o�3�&�έ�I:��8tN3�`�eT�Cg�xl��v�O��JP/�c6g�s�nXv��LONԉ�g����$�+��X�EC�gӇ����Ȑ��-T�i��!���Q*�l��o�8.�*')�v��Eh�� m]�:� �Ùv��![\e�c�hq�:%*r���|�X���.B�������e������^�l���p�el�g�Z�T�ƓV����)�_} �Ҫ@�7ՄZ;=�ȍVgŝ3 ����C�"�?�*^�/j�h�T�h\��EՓ�R����ܬ����Q�Q�wfT���R��8�@��g��L6#�/�e��1w��ή��Hf�a1��w���l	�����\; U_:���T%�٣L8V;C��>�cJ��/��Rs��f\�X�u�����y9��&����I�,� Χ�NDYX�m!%��o�Č���[��^!��st1,�C��E�8�o�n0�1Wߣ�g3M�@ѐ��!,���u���b��
�V�O�qp���u-b؉�Ҳ�k���a6SK�ʺ�|���]���=i<��������
��mh�x���J�e�dY�DMH��xȎ��3�	�%(��@�,�-�KK������p��\���|R0�i��
��߼��	#�\���+����������6VM�t��9�Y���iV$F=ޑD��(9ЍYx������)4#L�@���Y
�6�탃���X-dr����˙�q�9k�7�qf���u1*�޽�]��o?�vy\���:����#8gȿ(� o:���U�$S"��%����Bŗ��\5��~):57�3�ظ渪����cNxxE�Z�0/$��V��ݹ�h9�a�-/�miI��E�ŧ�G����ڏy�ƿ�;�nkp�����F�?�OdV�n�D���g�#Q[�E�k��X��Y	?�;��������+ C���ihhP��@�(�m:ܔ<�/��|��/����3���4��!�����<��&L�j��]���3�n��oP
�#�u�i~��V�%��]���2��|�&�ܸ�B��>�q,�|��0IE
�\��69�v
��Z��6;��_������P��$���9�J�H]��|����F���T�
E`�Ph�@�*��;*89��cn�Lc���ʣ^Ax�~�8���"�m4����#/��'s�\R��;<���^&�xW��Q�Ƴ��&[�I"�Wl@���9e0-Qq'������x! c�`�?�=�O�~=e���u_. ��0��,ٙ$���{_�;_ţ�qn����a�å������O�5��nU�hD^��n��y�fV'Šh�AO+}�ox	�O�{�ְY9�)96 V��?={b]f��>w��g�Qﺈ���;5/t��e�+&�G��3~�2�ߊ�a�^��;�%"�X]�����7��r��{�	�ɿ+�>7�� (�j��[�ڱ�>�����o?��O=��N5u�,	ZݏN֫V�$w�.vd�� <�Z
�Qۢ!ݡy�I,�}R���&"��M�<̳U�ET�}��ָ���kO�/gDPw�;�tfe~��!�e�"&L��{Zav��#��yY�{+8kn�X�i��Iޭ�
���[��M(Dt~����ᎰY�D��둣�1�JSvv������o���Z&ӏXր)�!�}_l�<?t�f�Ӌ��u4���W�)���%��Y_�錪�~��l�n�׬��%b$����c��;��mxn�1N�������aM
��c�\&!&��2����k��>�!p��Bk��
26�p��&U?�Ue��`H�KMs����8������hn,�$-��c�2��J�e(�:��&FUZ̿��gBK(���Uȼ�X�i�]&�g$⒰Ey��;$��g��#H����7o���:2#���Z3'O1���WW֥��t�CJ���m�,,����XOݸ�i��ۜY!k�`�i�E��k���#����[��Q��c�<9��$��b���P{��ݵH�{z����=���(�H��YȰ7V��H��U'�%9Y��!�FA��K�&1�r^2�2.�qf�� m���x�DFi\�iX3�gt#�3�ˌD&��#4�<�{��N�
'���b����]_� �P�!J��g�Lce�����'��5Ο�������{���
}��Kcc�;9IIΜ�����K̅n�`���	�I�g �>�l,G�W�6�;�0Ƌ�>j"�^+4� �
�����Ϯ�5��1]���9�bF�)T��琰�_pB�V�i/�![�;f[����P֟���q��t��I�:esc��(p�7o�	��=^/���Y?�:���
�8>����-x����S{���O���?���W���%�nnoւ�)�c<c5����`�O�jC�l��ɛ]92)u�+m'3C���<r���I��R���ꁳ87�"�f�F�ĲsrØ�!�&Q��-�;���S��y���u�1T�d"ei��BC��&h�o�b��+�_���~l��w(LQ<��U֎�;"�}�!�����{q��%��
�Mq55L��ۥ�o�MQ��'��6k��!�Y�۪`�P���+�	�a$�u���˸RO͂F���5�h&6�,�w��j��
܆g *�g�I�,l����j�?�~[�q��6�sN��=�]P��M�\��d��'%�ғ�<(��=7�qZNa�7d@���]q'w� o=����pؿ`��^�,m��g��~mх14�q#ig`��:߄aOg���n����?��7�颸�Xɹn]$~�f<�S/�=y+�͞�gp����OKE� Ӻ�>�Hk8�M�)�|�2�U�)��_��Hb���*~҃�}������^��v٢?e���AZf�Y��D7���ulG�p5��K�½��F ��Lڽ�b�r��z�=ѽ� R�]Id�hS�;�J��H�AȷzU`c���}+��y�HQCܳ�T�Ƅ��ɢ$���t��O�8�R�V>�<�S5�ͨ�jk�i{��M����*�a
��y�������~O��I�`��d}�y�.�:���/�@�yvd&L������&���zE��S.�����&�m�E���FSc�dp1��7l���ވ�#71'S����Fo� �@�h�Ơ]��l0֚-x�W��������6��p�:�l��Ș3>�31���\�>ܾ�QK���иhF�瓐��1���id����f�w@��D��������+Q���@�@S\��~��R a=C���P������Ȣ�`�R���9�}��m��s
{v���ݸ�P�U�JΝz�N���>s�/>�f Xǒي� ����&m�P��BcT̿�� ;�\�*h,��2l1�Ba2E��s����<GtJ��oto\�b��`��CS)��g�Ϧ�/ґ|&�����a�/=��I?j�©��m��Ѽ8�y?�@�T���L��AМ��f���6�m��H�5���s�Gk��f��<��u'@􁕢=B���a���ԁ΅�ͻD��[��@���(�/VI����T5ڄ�l(s�)
΂̂	���h+�{��:��"�s}ƾ�a�OG��N՜#O{��\]���hE�3��S�	M޵�F4C �; ���+ϳĩ�!T*��r�����+e�� ��dk+��3�]��٫WZ����)j'W�Cʭ�t���P}�EX���z�a��e�l<����/1��N�*X: �5��
�NW�i��]p����d� �3l>J;���L�u㬖!�-߰��%K��U�!Gv���#�QB����6
���Rd�-,W^>�p����$�]��f2��>;d߃A͛�~�M��e8�}��(i�]����ᬃmZ�
��z���E 5��#&h���Ҵȗ�~��3�T�����~Ugh�4S�R0�N��Zƀ��
j�典�]!p�5���ju���a,:�����K� ��I�a�wa��]+�?��PAd�{��	F�'X� �x��_,E���4	3���"�s��W�٥�sJ�\ ���`��H��VQ'0_^)���ʆ�9E#Q�?�?ٌ����z5��(D=|��Ѻ�R\a��q�9^��;�!���΂7H���C�Z�s�k�!���	~8��VH�Ό�E1���؈\�Eh ��dI�'� �Ę�6,B������f� W ���.��\��~�RjD��jB�r��"�2���0l�ҁh]��S��5>9�3�͆�=;���q� E߾���!��y;�KG�eYk���������:�.�.�݁�̵�2q�ױ.;]ߘ��c�nd���f��*6���7!�?$(VZ�Ċ�.����� u�A$�j���	C�˚�c�O�r/A�Yݛ����E^��#�<��[|�RB�)��g��a�\��8!#�>�e�<+�z_T���$K�³��e�Ŝ�����j]� F��8³�T�Fx|!;�GZ� �cv/�}��ڌ� #�L�5\xT`�5����(@���ٴ^��M���@��`f��g�= �v��?�搔_���O��4���&f'���*��-um}��+�ך�X�`�+\���BzbY�� [�g$[/&�a�|���n���QW] ���I��� -��n�{��z���<����7�
_x�!g����)�"��]}J-��$1��Y&��/F�� ��E�#Żݾ���dH�	i)��(X!h�ct�6��3���CAg����̤��f�`'
s=r"��&J�8�ռ�&a�MZIK�bU~*I�H#�ƪ��a�O3o�P}k�����U>i����>mŌfq�.���P��� �����%3�I���@u�q����&��`���Tcåi�}/�k��Ub;�ߨ�!�߄]��Z<td�b}@�k��r��Rݢ�L�yDA��
a����a���[{�e��5��3�QK������d	.�X��@{����ǘ��
�ny�ҡ��
�HBN�Xɬ���C�������A��(͍r��zaҪK5Vŗ�]�9�|��g5���Q�T�i������YJ݆�Ĕ�Y�8�x<�=W���[� VlTlkVN7�谗ގw�cfq���Z�W��T}�ArY��W��gHG{6';�^�������pe������@�@f�г�!�����c�<m��\�=�y�Dˣ;���;�5�>lD|�8<�t�+�X���+��M��h:7M��f-�l`+�(�Tm︦N�� ��{��8���\�<�f5�9����Ƚ �F�i�T�{'��L�vT��;��_�`,;���y�d������4�[�8۹RP0W[6Q;l�#F36�x��3z.$k���HSH_�����(���įe�gk�B#��fH&-~>�@!���7�[}]�E.aH���Jϔ��#����D)H����)ꌌ%dջ[���r�fK��P h}瀴sѹ5/�*���<���%�\4מ���	0w-��;eT�D^d�.��C>̆�5f�v-�9mq�>���ca�!!��g���͈�p +SM�<p�1�
P��¢�Q���Ǉ����7�:�b@w����O$��p��`��8��1��V���;�}�X��p�θ2ƈ���X�yϣhK��XK��]�fݓ���*�9�B�ïS��|`.���!6y�BV��v�}W�}'%�6?F$��1@���>i�+��F�m�9С�x�{?�'�����[*$���Q�O���eL�sU���^]L[,���p�u�P���II�����97�o��{[�vV��@F$���	}f��ݡ:w�J�N�Y;r�f�@1����䫵�(q��ӣ*�e`U�q�sd�8�����*�QB����͂:��7T�;6ͪ�p]���K�q2t=�YD��28�K��z!�0dz�!.�q� �Wj��Qۭft�N��:�c����V|���R��������iX�6� �{l{>qO�3 W���N��k���)<p���]Ibvb �xk������ c��K^�$�wbt�}�R�����g��<-�[���Ѣyjo4bd*��n8C�Z���A��2Q^�ր�TR�����F�H���%ŭ��	���*��ޔ��[�m����F\���ɷ	���ѯ�GH\t��^�gt��?���3!2���}�@���>f
��]qdQ�V�sVG.ǵ*�h�[d�8���ql�k��	���Й�<�"�W�h���;�j�
�G�[Iq�1�|�7��ԙ-�����LΓ�z�Y�/���?|�!E�c�t�W��Ȧ��4/�Gze����|�H8ݯgWwx� '�J+;�e����/aNO����/�n%�}��#�����u�!~�|��|K�|��ợp������a��b��C��y�DQ�c>��Nc��3����ƈF�-��	� �R�ξ����1����ϑ~S��e3�3S��(,mKИ�����A*���'LzU�T�>eWҖ3i���dN=a\�$���0�+���A�-�_s�܆�ٴN�_���2;��������;�I�.��9Ә�d��G�k�2W�D_��p ij�)�A��C�: uf�G�(⦣�W�T��پlNJ�R��qU��썾#��3(ϋ&���M=T����x��L�^�f�2���E2�z_���\�δ�r�#_&Y=�H����� �}�h��ZG�����}��Ϟ,�$%ۉ֑���wϊ37�aC��]�>�5�,�J�S�������lI}:R}�e��rF�(��a�eĂ�/7�܍�
�C; N�Z�ş~�{�4��7�{��xə�j��D�ą�"\�@��I]9�&Vr�V�)ke�� Q4k,��v=fxZz[��cs�"�%�YdoC����3f��E��:)�(_{�v9�� 8D�Q�t��pߵoh�9��?n���Zn�+�BQ��cH��Ӝs\�r[�����n*?;��$��K�/bS�����C����W�9D��>_��6��渱_����9�:�q9�[dk��9a?�lH�S�gfTj�͞�8h�~�~B�d-�s����.�\��ө],���Z�t+c���g�A�=��>Sv9���n��0���4���]��}���{�:vl/�h��3ɜ��-�H5�N�A�9�;U��0�_d�`�;\��S�bW�7��&�'9w<���BI�M\8S�N�gQ����Ȭ�,�
�� ���j(�aܱ�R��y^{��NW��wdD�,�#��X>��w�5	=�H���,�I��7���k���Y=3w�c��-�7�sIB@�c��:��B�!O�2'[�W��k��NJT���5�����/Vߴ|mU��8�.��0]�)���6��n�7������k�.wW�����{���y�3�.� �C��n��
�d�O.����p�f۱g��7���;�ޏ���#^�q�ԥ��x ਠ�tn¸Z�U�i��×���˔5R�= ��X�T���;�ux���-r���h'y�����R'�?%:E�`S��K������O�\���Sv���7bR�+.6fv�sc�mgvtlg��^Y����4[ׂ9�Nw�.M�����p���; ��;d���f�%&~��#��0 �<�D~H�`ї�b��y�;�ř��u�U��i��p}(5�������Pa;w	~��:�ܥyJ�l^2ibD�w��
{��FMK����h��R���E��_�Ol�Lc��FE
�L�P��wUp X��%������J��ɾ(姒�,�5�L��V�f!E����%�����Du8[���<��
�~�0q�Ή�����S6be����P����Jv��b�'�\5wlٻ"(�-h��Q j9�
*��1Nʨ�[�e������%k��EX��~ ��c�:�!��#��R�]��ħ���]��A��7UǓ���98��Q�#��eo,���)�7. I �z'.A��]��7Sn���J:BդV-#�|���.���n�T��>�H0�.O6���S�wxB������c.�t$!��]��s[�����U��Km�=U�΅�
T��/��.������P�i�˹$שג�������BǼ�\���u�8����Fb5���UEof��z>'��o�y��ܝ��t
1� �r�+�r��[n&���͐�}Z��My�K�0	�Р�3e�!�9���;�� F��Z(�U����l8��hN��VL�}���;�t	U�I��R�3�<(��c�,�N�p���_#��Q��&Z
��K��Y�����3�-��
��}<�Cǧ� �۩�I+
�/�{���U�ֺ������&�b�S[є֑�/_�_˛�����؅�U�n�dD����4� ����@��؏4���M��L�1���"v�VLOP#|���kԵm�����4����b7�A���k��0�?�Ũr�1��	|`��e����O���v]����s���P�g��'l�>!jG�@	$àҠ��ĚDO����M�n�#:�ξE��Pl�D6�4��Ut�@qbE�]��sE�)s|2f����ɒ�`N��a�I_p�l�^�����YU`��`a�(��LX�^������������"���9�>��<��QOoV��(P�'�of� Ce�c��|���=7O2�3|�S�R��>.��,�G
sQ^���'��m��c�Q�T���N�LL��黍_*��"n��Fz���:zB%[��Ö�H"����8d��:#b�çgJ�f�<����V���f�Il��40.�(Y������ٱ�d����z����3�Ӭ-��E0���f��0�2������Sǳ����;��L{C�M����I�J�`k���{�w���("��P1���3O#5�R�
���m���ֻOsͦO�op�Fܐ���5�V#b=��a ���a�U����>����	���='�J�@�I�O\^��Z �R9���rL�[H��.�����官)�̾��8saG����Y�h��(�pn:��_o ^��F��,�c=�:4�;#W-�ذ�	�W�(��=T�-l$t(��
��buSd��(�7[��)i��h=^$���(n2?6�q=\ଥB�b�$�n%xq����D>��Ȑ�� ���ܢ����h� �G(��T+:-�ɋ�ˊk�|plb|T���R8v��{���gp���^8�����+�[E�8�Кb9)�[�- �ʅ�$U�ۛϘ��3�*9* �y���2Y�T��]wE��ӈp�qabf�tcj�EվE���_��_&����=�/Zq%=��0��_��*H�(�y�lį]ۼ)z���;kX�?���!I�Wޞ���y��E4���E�GZsʕY���S$��@V ���d�&�DC�3:������G폾��t!���-{�R�}���̫�}�Ys�w�r�7갰�Y�s�*C�G�|�<RYU�����~e�V>�40p)<���ͺ�aQ�jw|vmK�ⅱnr��d�rV�ԇd����j�e8�&F6�ǣ�i��Hk����ӮЩm�u��^��h�:g�*�����L6޽龿iZ�h��U�Nɀ�r��Y� Z���7�T/�kn$i룂�Q�#i�z��
�8z��6��]�HJ��Bxԕ=h����s��F���������C|?��R�e��a3m�x�WUL֥_�	�Xh��9L�Jd��<Ғ��'=\R\���)� Ⱥg�+��6;rRtH�xX���W�EE����[$}Q3����Ѿ�:�S���/��Z�*h�>M^W��4ɵnH��U�9�t_M�e-�� �*����^c
�P,/at܃�O��R}�E�@���,+]G�Y���K��>�G$
R����@%��v�s���`vF�ͼ��\�QHv��z��Q��3�������@@��p��@���'���b��
Ӑ���f&���Ɋmg�LR3x��J?�Ɗ����߸����!D;�Vs~�J�/i5Pɺ���X�Ts����2&� ߬NB~�g����n`L�5I&�t�b�)R<I2����7�!v���d���s��NiQ,��@Y�肊/;�it=q��Ŷ����%�o1xj|���E�H�~�ߑ��jI1F��9?�Ds~Z[�����X�Nd+o�2�cP�8ێ̿�C�\a5m����&�Cd�k߯�T�V�;�^ҏuo����-?#=7oD<�Li��@�I%Q�����g��*�ԟ�l+Oޙ�IvMC�C41
*�.���#i�ꛨS��e{/��DQ��[���ƎhK>�jR�x�t+S�X��']'́���°�)���ߴ���{*C�sЗ!Ы~s2<_�!?v�v�7�d+��D�п�)]TfV���!�5�����"uB��a�~�,�*8��<M�Y�&�G�Vһ���޹�m�/ �
���"��-�c��6�m(m����Rq��p�@	Y�L��E�������+��!x+��|8��m���$��ܹs[���� xn��!{���h\9��_��Ӈ'RŦ]2 FA;DNE�5H{+,�C}�'q:�ir$Lj�Q$Jr�D�Z�DA��bË�+����y$���֏[��_NW��y�}}��;Os�"�����92q2'��j����dd�}}��D�Wֻ��u��� l'ii��&*�~�ը�z, �,i��4:�+)�w��VYpr,� ���"m�B)E��w�5����ms�X3��x��I��Exx�:Aec�*/���ò���A=�[�Ti���Y^xK��N�W�v[������XXT�y�5� ��zӆ_BkIީ��ȑODw�C�,G�I^��ɱ.~�T�z!�n1%�������y/��X�ћ���؄Y�KT6�T�l�J�}�?A�g8O��C�N�6��Ƃ������:j@O��e�K-A��É�)��Ȧ!��[�U+]�LZ!��m'2 ������yB��������d,Ǿ�'�����y�blQ<�ʔ������(C����wtg�B�l%���&��<D�H��[�Ȣ���b�5�@�D�$2�j�r�f���j�K"�P�uN�>��()8H�i0"�t���>�3�/ )��8�?�6�
�8�|�M�.1HG#{7�a�^�:'7,���S���yU3�%�y�_��Ѭ�[e����}�d?s���'9�2'3}yIo���G4��5Ō����N�Sm��nF;�/��9�>���X��Bܷ5�8��㓻��.�3�ߘ��ӏ��x�z+����>a�y7��� \:Wu{1�N�@���$�'����[ܽI�|���r��{�(�ՐQ��Δ�r��n?t|)F�E #Ty�T$F�.�D���Bbђ�fǺ�#��݂Q���H���v*�L#����w��0��jP����p2�q�w��vt{��}ֽ��6[(A���$�euh�G|�x*��I鸱R/h�Od��
�F�����@��L��
9V�y���r�Z��p�Ѓ�,�b�W?� |�Ee�U�e���=�����ų�j^���ӛ�~�����@&�_�%A��-�қ�'��p#MrV4���<;j<��-3z�K�N]���ͻ���*q-nj|0U���Mr �k-n썐=�oq��O�!d�d^h��Ch;|��|�u��q�Fc�/���n���ܬ�NyP ���7�*�]�ݟ#yienNG�f�їp���ڎ\�!VOØ��WaԄ+V��W�T0�����B�:�A~����JC1��T�2o�4�܁�����`�QkDTD5|9�d��������h��D�$��1�6O?��v5�g���(j6l2�<����:7��6���r�J��kQ΅l�p!Aɋ�9�"HC�F$;P���B��|���Օ��YO��UgK�P�lB_N��C#��%�v�ݪӉc�����r	�'3py���iJJ�J�ae-�u�����;���9Ʈ2���N:T%��y�G���x�J*���}4#�z��BE��pԤ:F">��^{U
�����ĝ��>#0E�^)�4s.��q��
�ڊ����豣IG\����.�7�.��ީ���<h���ϒq�U�]�����mF@�y�4��t�G7{q�wS�J�TV��Ʊ�g�9,���zs�T�/d�l!�X�`�,���̊x���a�{�IE#�8F���
&�r�ફ���i��$;"\�=�睿�ЕB�������7��p�XgM�q����uWRu[j��QuZ�:��r��P6P�T�re`˸�\F^P\����O��. � u���<���^��ȝ�.Ѷ����I+0��).��Ѱ2n>т,����z��k��#$3��29:`iWx-�ǘ?<9L�,�# �UE���>�1\� rQ�3~?e�?b���c���@a�^�۬���#�z�t|����g���É%�yٱ΃4V�d..D�^�����a�h��fͨ:�.M��v�@��{6� Q����S��E���k��u��n���y��jZ�9T��dT��F�TN�Ʒ�x���mA��C������c�7)}�)�z��/o\yYZ�I��� Y�.��������%��K�6-R�9�v������q)b���H��U��=����Y��u�������[�L�Z֭�,�r�ݥse� �u8|�8�]��w��f��Vu,u��32��|�W0:���u��+�uI%��=�Qa�PMKlL��6��j1k<�Q���;>�eT[�`2�ͽ3��E7�-G@ʆ��m[��?�-�*�eKC9t_E�~.(դ��b�����%�\^��5��#��T�+@�Z֮|��i�p}�\��83;v��>��_����Z��3��lt�z�,����s�qB�r`O(ꚕ��/T�R�0�Ȑ��X�ն�Ua;P/AO�}�����Q�Tc|g� �
."����`7Zo{Lj��]i`,\��&>�>C3�&�b�HyiF�r{�-H���g���2�h%��r�����u)���P���;E����[�:�ts2��\_��	:��P�K��B/x�4�4+
n���@�ؿɭ�:�HA��7���8X���aͽS�X.�
7�ڼ��y*.��JEd�cF(����s	(K�����QkmI�Q-�������X�sV�6+�;\�w+i�w��}v�T���G4:ǟ��U��y���0bH7Q0O����u���1�/_�E�z��\I!��.Y4�I�į�b�o���|T/��8Bڛf. g�^�R���8OG����J|��܁'�R9��Ht�%�m�D����x}�ZM���
f��� ��>�۠_���p�~7k�Y��:�]���������]QNr})X7+{�V��e�/A�y�J������o�]�F��$�v�s_��<����_��;�%�F��;�Q�l�(�2��h���0�#���w!�&�p�^�j"�+��h.S���T�WX0�M��>���~6:�[��ZXv�������=�ড়3��p�C0�	M���8�V�`CGY/d�<LZ���=���3i��5��7�,jo	4V��Ǝv{E|E�f��Y�ZO�@�]8����e����V�^|���F�@
ƻs��� X���b[��������a�T��r�o�s�-]�&��R���$U,�e��^/��}9���� o��5��A����K��P
Qut�S�D���uhI��w����8Csc����g������� Y��Љq/���o�uK�B����y�t�^��2�`����.���[����.�2$���3���/2�K�vO�f�9o&2�O.k{M
ц���XЭ�K
~���BVv>�Gn'L���/;��s�`]��?΍O�	1Ӏ"��B�A7��HV/LwX��Q!\	¥��'Y�V��J����j�t�b���C��H�#��#T�������1�7܎8N�b�9AN����O�*�M���x���b��AS_�#稏��>�׾_B���=�W�"�����7K}e�P��{�s��z-/��7����QJ�L��a}���Yb��(���h���m�4̯�I��{$d��y4i�V��K[�a魶��1.�,���xD��D�w��fJ���~�GdB�'ūw��� M}x��pYݑ7zԫ�P��.i��o�B�C����x��#ܹ���G��xai��3%�n$Ho�r�<\��KZ
b���{e~�- ��@�f�ؒ�N�C+\*�M��+��"Y4vNX��2{���V(K��8<^����9�86 �Ƈ>Ô�}0�2�H~��E8E��z��	ݡ�۷�=��&(B�|��)��76eŮ߉���z�;�������=������{{c��ٿ6<������nHp��C�z��N~u��э�]vq6##Iv������ډ9!��m��h�ά2��9#�]�5������P�i�e��N���ߑ�8Ud�C��.�_�U�_1��=�}�s���Bp��:ݫz`�~@��Vξ���QQ
ad�^���J�]��WmD��Ae��z�oZ<����?�'���}�כ�મ�=�mBc�G�ϲ���4�ă8���h��a�'��4JV0�i"M�w-��+f��������N�Qރ}FE��Q�q=���2��/=����������p��]��R����,�7���:P%�����6����? s�V�$w#�k; ǣ�噷��G7����BH�f�$sjK��K�Ё��;bR	�3�9<�x�Ug�M}n\;e�&�hi��%48�t�ȶ��i��V�p�<��t���qn.n�˲�7�w���اLO�X��QO!�E�ʻ�*P�b$	�n���|2���;Ƨ�C߸8wȇ�m�	9K'W-Ӗ�n?�T�w����6v�c�V���x+��y�A��w�q��C1w��-������%�	������O����v�-�]����6@�rқ8�ڳ벸l���Q|/��>��ݦ��ٯ^'�:�Wgbђ)��P"��r#PWe̻�����_a����Q'+}=.N1�U���{�daU��f�>q�%����E�.�)�>X�>2��DE'm�O�_66�B%u�{Td@�Mk���Y���ҩ��O������,
�LK
a�:i2��{��Pt(8������	��6�'���,��'�8OВfM>Fj���b8)0ȓO��,dCNI��խ�]�xHj�O.�=گE�C�|�c�@���[;�:����E�)�f,�g 2���w,�+�<]�xcŬe�#��{2��1
n����63~"��x8�֚9��Zn三(��!���{�������D6�۽Ie���qԙ�?t��{�xd��]�A��KU�Ca��I��P�e?�U����5���l.ߜ��f(x�P��E���є�o��<1�sG�e?B��l"犾�먳3"�r��U��ȕ���j�]�Y���A�j�l��5�4X�H�!��lg�ϐ)�{�������U��x����q)'bq���l.�<�R2���tvS��iOɱlx3�VJ(X���Un�ɸM�?�D��Q���G�|�Ӂl��$�~�����ǰ��rJ"�פM*��߅!���ɸY��c�:���$�V���m��{g2�7����e��j��A�$�"<̧��8�/��Uƶ:��� ZI�jw�f�VV7��^�=|��j�ߦ�L�$�t1VrHҊ��G�Bi8'|<�Ӹ�f+�PZ"Z�z'v�ў��T��֣�!l��&��"����v�_�H����i�R�/ڬQ2�$[.~Տ^�8�����ז���"N�+���c`3�ƹ�@��hԹȰ���2�s���+�(KO�UV=���O�R߁a���v�X���t4ę�K�z ������ǝ�����_z2_~�����.��}�Y�s��e�7�D�܍���=����y	�8�w�ޔnö�tNAZg��)������]�`��%��αT�'�Le�݄Ե�8�Υ��[�%0�Y�\��2"�>��B582d�m�����-��t���_ͦg������3oq-�`��Ա�lE�t�o�����ح=���T�3���j��L�l~ePR2�n��hJ1��-�5Z�U����@�;�q:d���S햺���U���S��C��p��1Y�&{=�n4�	�4�_���Z��O�0恧���e���f�o�#1���
�+��=��8uI���u4Ȑ�����+]^�i�i��Mm%G ܐ�'\E���^�j�)+@�n���|�Qy���yyV�sYP�@���Ū��Vp��Kt�\�>��1,D�d�ґ�I3C�}#y%�����+�G��-��z��	oW�ۖ"��@�4��	K��t�¤�C�s�v���C�0sCra��8�"�A��c�kP2O�cu}me*����T}W�����Ӧ��r���71��A�u�H&����Y��h���8^��)���y �}&��-;�,'gKpm��;G�MDM�m��=+ħW+��v�qh߸��I�O4�n[�'�.d�D*�����ƴ͎.����P;�H[�j&�
���Z�s��{��߷�2Z?˹{
�
�o�ņ�3�ҽq}�Z�,Ѽgbwu�#���5�Be�e���	�M 2\T��ݣ͙n}�B����crй�/���o��^�R�,B����Dn7�#l�~��Kf߂Q	Q�$��1:� ��
{��BҶO�pdzz	���.��,�Z�Y��!�3���&�Q�Z���H�OSJ'"���`��ٺ��ް�P]V����W�bnNn`�p��-��@&&��0��r&�k��V[����#�>�M�u�+�vfͬ��̈́�t�L,}�����m��֒(�*C�����g�[�&�F�8A���K�ppK�a�s�C��S�#���R�KsJ������/�ͽ��k���;;�f��:X
���d1��-�4�I���b0%�0��B2�O�\��G��<�>��:S��#�؟!�1�]�zc�o�D8��(@��s�B�ZK�Xd�N�+�@Q4��b3 �oi캕�#V�EO��+�L
ަ	�f|�J�qzq�������ض�"I�9����A�澹ȱ���CƼ'��w������X�7 �3��n�0?��5nȫ��&�����A�+.�<txD���b�Ѫ��s�T˺r.��b/C~�� �؈���O)�d9&�ړ\Z�}��[�3QZ^�GBjI�e���V�ﻆa�bE������o��6���s����X>�cp1��bѧ��c���g�����)IP���|�N���)O�
��Ю.9Ų��S��ʹ̺�U��dU0����w6?Kf��6��uO��$��_��m��>t�A�W��J/����A�q��vIo��@(i��Pi��b�jД���'U�Szf���@%z\sz~����Vp�_k���	���9v�����EE��P-ϵ��a��y�� 0G��0�`9
�Y��z�
l��b��jõ}6<��&�?8to�H-�x�dK����7��{W�ܨu7��/7܋� k��v�_��"����YWHc��ʹ���Eo�p�	<��Q!���Cå����>��J�5���"g�������zLc���j,��x�ZW/4��YEK����'{��S���[j��oW?u�)y +���wl��t�'����x��P5$�iڗÊp�6��f�!����#�]� .ē�[ ~j3�˱�eb�!�8�	q�i��T����-P����@�3^��Tf�1J��ި�j�5�#Sk:�i����n�F�M4�&5��vw����n>O�K,�*�����<3V������Cރ��o7e0���~�7�J ��u�^_+'`��B�e���'(�\ژN���D� �zB�?H:��T��ܯB�eEA�YZ�x�jo���Sg�f|:��IU���a�-�[]Co�-�E���Z ,�h�R���~�)C����;��θɘ��f�P1�SX;�6CF�;�\� )���DsE2Ιy�5E��Ɂ�k?��`%�y�I3hS�p�E8r/Qܝ�l4FW�P���X��ß�:N0��/�%�&��/�ރ�����$�J/Ե����U,W�3�*����+أ��=�~�[��F�d���r�~��u؍9t��,���NL��c�~�L���n��]1*�5���*�z	��w�RK>�������Bz�q䅬3�]�����=���AmAm���r�E�4�gk\r����%�9R��n^��C-V;]z{0�����~��\�e�v<�#Z�E��% ��t"�I^�R;Y?�_��Y�֭EQD���uT�)�����_���J����3:�~��~��7�w����EK��!?Ne%/��#��ͳ�_���ge�^Q���#��Wm�{FD���3%�;NO����2sMRP�����i��S�w�G-Fw.��lzקmƖ��g���-v�+<�o�R�
T^���m飹�"�LG���{zBm|O��3y�HF��@�\(;,�,|�P�����bL0h�`�[9�m.���	���dE-���Yj���7�u���WN��d��9.����HK���]9פ(��_r�%Z��~�[����
�o�]$�)ʽ^-�ZΌ4�n/�m�&/�k�4|ߨ��K�д�1��Iu8c\�*�z��5�sq��4f�4�x�+�U�g*�hy8��@J�~����S*VH /���W�2Vf����,ζ�yj��� 4��I֦�V��|dg�RyK��m`�B2��5�9�^���ު\\�Ȼ��lG���(�g�ݧ`xЈBQ���&����ړ���~կ��k`���C�9<�3��U�d�%&�/L� ���@�JB@l�<����<6�pn펙i��rB҈�w�a���P��*�����Et��4�]g�֜��r�a�v������A�GC��Mx�G+D�$�y,�i��a�^ۗ�����qN�O����i�"��&,���E�N����89>��MJ�7�b���O��,|Rr�\��Z�*UP�<	��Ÿ i�[�n:��U����̾Er�dZN ����d*j����ͮH��]�jn9�g�0�.+X\�Q���^5,�#��h!�o��wހ�Ml������U�"��)�����|$��	�T9�6���G����q��_R�I+�E��3�O�0�>���[�o_��Zd=_b'l19bn!킢�Y+���w5���:K��ON�8�D���"���n�sP�h�L����׍����n�è9����`g�炱R? ���b�Ю��G59Ny4!�D�A��)w�Q�y�H��tɞ�>�t�Y	���qN�6<��0�n�)Y�vʥ���#���t�+���d��j���@;�ݯ�1���Y`��|��À �].�ujhr��>j���q+����h},��^=v�M�,z� ;�,'�F�U�5���ozO������2���n)[=�P&v�;�z���_/`X�� w�L�����p�"�!��HG�~��S����gȰd���q�0F��Dy�D#�7�����ܮ~e���%k�@�7^9g�7�!�J�oGz�0U�p���3�K�37� :4��9�!�Gs��.`���bB��1�qG ԇ�1�\���[�<��ʦNΎ�r=����D�4_N~�@!������<�ڎ�'��$OM��>�W��~J=
@�8�'i���27L` YB��U����}�,(�>��֜C�b�.�,ݗ�����p���q���1�)]�N�Cn����BLΎ5#$t8Zzx���4�;�-�uқ)�1s�G.I1���l%Z��������h�膎Dy��LI�v��׵��+�12V�:�s��*���
�LB��ۺ��3�-9.H�_t��b���]b�֙��و]^�L!��n`F�y}��^���?%�O�v��B�S��rD^�d�����u�QX�� �����E��<����^��KV*��� ��I�p$)h�P�$cƻ���~�q����:����~=Jz��uon�6��~y�o��pBO@�_�&8���飧5)�r��W)��}�z��������'Ww*���2����_�cP��\��b��<������}J᧋�F�-��RY�q�L�J�&y^_����A�v-�+��
�Ry^�X�ld���p��{�oQ�'�a��
�w�������RL�&�xE�X;��8��%�߱��黏E(X^n�:�����R.�c�����n�$PDEgS�QS�v�����2�������`��S�y�Θ��ĶΏl�I*�峓^?���[,��{�#�����R�q���q:GN0K�,e��XJ���k��Xd�_\��	�vK���~����Xy�����3nD��;W�>��`ϭ��,Q^Oi-a/dG����#�aJ�VyK�Mb�l��������Vc�=��
��eB"��L�_�4�K�7
U#�a���SNJ��S:W�J���9��e����������f �h��M..?���Ҷ��eyf�(u�Ɛ�6���U$����{Xs���mWJ	G�xx����(��&2Q�����$���'��-�Y��Gͬ�R�!lQ$��ؔ���L��lAO�Z�瓫�EVD�#Թ��BgsL�!����F�Y���#kr1��ɓ��1����z�!�լfh�e�*�T?*���fcC*z߮h�=��"jk�`=���*U]�~��L
��n.��0�ɼ8U�}7Th/�h���B�_���b�e�յ���l���]`p(��CġM~@ V���o^XC8@��kQ�f.�^����ܐ]Q-���>�t�*l�����UɃJ�wd��1���̏���GTl��O���Ů!���,�ڟs�ԿXT=�&�{!��4��L-)��Q�k�\U(X���g;*G���1����*���PB�`;��A_���"SZ�^v�x�*�������7�T�^�$��Z��-2q��ß�ٝ)���"�	�����7�x%�� �W9��B�P�T�z�D䳇�U��XQ�M���;��.�6�n�d7�=�(�v:0;��]?��07O_��YcWK���D�}\x�1](Ȉ\�uɸ�Q���%]{g��ku�i��gO�LJ.��j�F�56��,2��x��B=;��c�ݟ3��O�fP�	Ȭ�����S�7|�0������|�b|���m�s�պ)����O�[Ox��c�Y�6�Ө�{L�n>�H�h�'�H��P�-˂��
j>$������]�8+�����n̿;0��������9"�ث!a�����X��4%u� ��X	L��3��Ð��?Ca#��BM�@�G����L2��L��Ce��r�"{���4F�X��3��zj�t���c��\/M�C�i�i��͂+ �&R:r�Z��/!ߠ岂�3V�Y1�^���-�<��M����J��׉|�,0�+g�ڝ�Φ(LF/��{���؄ZI9��HI-�V��v���r�����S�hQO��E�<�v���m�։��<���-�����s�PQ��7�)���ŉ��U��Cl�BH�#7��P�B&M��9=4���[;�����E�WÛ�'�F��3�Тr,eV�֪O��x�"���T(sdۧ�;=��F=Ll�F��Sr��\6���ֵ$*�g��W���f3�}�׵�D�[@����Qκ�7�ޱn9��j��L7L�{Dr�����O���?����	K�MwȥP	z���#�;�'���M4F[���;��膬_T�L$��%�|F�>�e�����Y0>B��ި��=��%�/C;�o����z�x�C�,�ߣ�6BK�?*��P�q�!!� L��؍ 	u��|���� %T�6x�k|������W.�9��u���d`;���*�#��C�l���ԃ ��Բ��6��V�ſ�a�w3�m_�Z����ԡ�>2���:��&���hnXK���Zv�D�k�W`���2ɜ;�?R�_o*2BC��(ݕ8	�^f|m�&C"`p�6�;Ut6J[w�K�H�WE· q�q�N��D�#ب�W��f�W�o���ѐ��|�F�s��i���$�>�%I��-|̳�7�q��Q �USض+����A�v�㵳��y9�t노 $��ד&B+�$�6X0�͝Ry[��5m��\M�@[И��[��m.�k�k���UP��g��=�v�\�5�x�߅�c;߂�2�@�Z>�uA!^��:������9(�
Vx����B$���~�,�ރhK�fݛ}ա�l��H�>��d��Kݾ�kS�ӯ�^�Ke4��(�c�?�#a7�Au��a���lG��Sy��(��4��$V�Q͕O��z"���S:G|��є�������,�B6a;�re�
��H\��qϚrM��c�2q�E�j�l �j%0֞)�yp(�ػ2 T��Fc#�O0���%��]3h������Q1��vm)i���D9~�������A�&j��\	�$N*!)6ӆ�	�/�~%O>����5ԟ�_�Z}7�{���bl=�7�L����*�����Q[��ޥzܱ�H5<����f�4j�L�A��ŹB��tѰYiF� �(oU�-�ᛈeK�'[)��l�š��J�s�P�EjV�����Ԟ�(f����d~�+;�i-�&-[�y(���U_O���+�e҆̂VL!�9U�e���7,�~z��Su�y�o>�&�ڣe]ÈB#(.�}uy@y��vI�{��9��[�Յ�M�y2C���)5R�h`)�Q�/lKHYDv�-3���
V����!����P�l�ݾnl����&d����O��)���P8
�����8XC�ԅe+6����a*)"<����X�m�R)\	F�"��!}��g�lkTH���Fx����8qj���JH/^�v"o�~�%�!��+]�.ŉD�����P�h2�0�o�,��3v�	m�qV�E�!<�+6�Lm��Z�ۂ^����K�׮����q�ʞ ;��.hVލ��?	��n�������d��kN��9�	���>Ah-�Ǎ��q{����V�:J�"�2�P�P����d�6�a����8s7�k���7%��UJ�bT���W�	�r/��rD�/�X��p�g<�T8��y-��"K+څl�7��$�}! �3B�R�T�
�`�H�:R�U�+������E3\n���h���rHEp������,)`�,�
�a�����)��oN��V���{�0��sJ1��n�d0DT5)]�lX'�
�Sz�_�8�P�r͹TUB�����ڴ2QYG�s+����j��m�S�)D@x�mQ9bSBO��8�0�a����]��g$�b����֤��&����6>,(��AB�� o��i=������d5�>�>��7������ؖn7yՎ�Y`��b��� �py�(�?���w����i��� Y)QGzY���a��2:SRP��;��q6��E�g|#3މ�';^}���ꖝ��ךK̤$B
ktFX�P�τ�6��@W�C�U(G��O=J���G���==^�pu7ӂ{UL��-��h�ٰC�g����;�B3_	tI>�DRRG���I&��㡢�aN&����~ħ�a4PE� ߵ���ꎷvm�v��+�d�f`"o���Udl���N�h�v���7�y��R�=Zӟ�X)�˚�>Eb$E�His�Da��{�)��G���]u#�A�P!!�2s"$�sq��^��w�qTK���U2��i�ep����o�`ɮ��r��J�Ju�T{s����~E���Zm�v���F�yx��Z�1g���/Q�h��W�8D�3���ȼ?���X,�>q8X9��Fz�|`��A�Ċt�g�gΫM`<��oȩP!�"�,N@�����FHF���鿏;�k�~���j���_l���R�]��q\=¤ P��|Q��0�Aߌ�-�	�i���e������]���2��eէk ~u�*�ĥ�\r�ɜ�^�w�s�j�(����P�/�:}`2��|}��pʘ��v����YegКr�sV�Z��zMj5�]�sv�D̓Ũb��x�!���,re"�������x�@^3]�n���� ��|(�i�+m�B3`VH�:n�3�����-�FS�]v}�J�1���kCDb,%����>|��kmxG1G��1�W4�1���o�pL7��$�Y!�n���(��hi�f��e��A������+�-ti9��}��j����Kt�	�ǬJ����/�	��N
0�Ңb8�����Yڑ�s�Ԫ$F4t�Hd��tpn��6���؁h���v3���̙�K]HA�_.-���Ŝϩ"1ˢ���+-���Ё��	��-F�$��	y��݌C�DgN��I�/��9f���00�v�d͟���������!���q��t�q��x���'�K9RLM-����a���v�Tdz�r��ƴU�z� ��}�بse��rTS�3�P��=�t0!T�zW��:b�Ӭ����a��F	�Ѱ�9N�����k`����<� ��"5�
��~�h����IK,��m��5!/�S�L�a���}��Mq+���%x���e��;��>���� ftٗ75b"�9V��5$�Zq�iY ��kwK̔��#HY��|[�7|&� \��+�i$~b�bXy�����mҌ8�<�3����'���Z���аi�Kժ ���_>A��(a�YB:b�H`_��3�
���Vɨ\��yp�=��
�F�@������_��cd�c-BҚ��ih�@�x͡�+\9t�[���Oɷ�2;5Y@�\ν���F#�%�U�`P�.>�W��P�����c�����\���y���Av�=J�r�J�"^��T�i��(�V��ו��?��z��I"e!�s�7	��Kj�^Ђ���ukd�v���={z�*��:����7�C�}/3�r/�s����"�LE
!E�Av���A?U�|E�lP"��vY�^�Spx�v���)0$.V���oK~�6x�'�l�k~�&��l�f
Io���P������ı��T]4�e�z�ө�ڷ�3���Z����xv��Iz�,�, �:8YE���������5<��7{��O�����q�{!F>�(�D8������vt�%ʘ�?g�l���Va���Z�wlr�� "��C��$�f�e+v��P�dMU-�����,��^�3��@0>��^�J�`V���E��l�>�Z�ԙ�xMB�'�|ހ�V�K�&������(����N��N:��J�%wJ�h�wPO*��lτ�aq+���	��m*Q��l��T�r7ۦ����y��.�\�3jn�ǍO[���4	�3ˬf�4~������ �.8s��1Q�4�z�o�GS�D�RE� й�Fh��MU{�\�~;#�,��0�"^�_�A�\�eD�J������q$q�u�fM)Z�O���^��P������SGI�엢���DA�6�bg�0��:��c1	�G�v8M�pX�#1�8���mc�X�_�hչ�Om'�P��L뎾uu���ax6)�����}�����| ;������](wi���#�W���&$ibAQog�R�:e���zU������cAx���O�b�ʣ;"�l�N@0s"<������$�ᴯT6.6ZO ��8=^@�_I���ޒ-�|�D������ "�~�,%�j��3���^KI�N;[�_;�xX���[�I�(����"j];m�g�ӯ��gz»�F/��^�1�̢����O�KSi��uKR���]���M|��G���Wx�@2^p��c�'l���'-��:K2+�=���H��o{�~�=TN|CT�˫@Ob�1ë�$�/'�ڎ�7F�����j��W��P�������O���Hƪ>ʾ"~@~��k�Ұh� ��0r�f�Zk�Aj���/�����l2}:|��B= ��6LX�G=�V.g?�&Uu�OH���M�C�򨙰(3zb{Џ�X~���α�\[6���Ҝ�]����f��gdB�E�i��+&'(L29�Z̆����ӥqנ~���P¿UM�|��C:��*4�Yk.�1���k$��Y��}7i�_��*��zD���q��͉?-�К��~���hU��qFo4��E!S�
.R�j<���B���@eV����Z��{�Xg�S����J)�'�V$�w(��*�?_C5���]�k���sy׸�<��#Գ�*���^����o�Q���i����:��%h�_�d�q�(+a5�=�/�$�W��gU�\B� s��Q���5�o��*���w�E�t��rd�#_�äkXE��*
{���(�&��Mc@��g�����n@�K�⤐���/ǡ���r�,�*ق9�=���>�z	u��%w��"I%>WE��b���:��1$�3��0��KQ��c���e�S�UE���8���	[�5����#�ZPie�5���E�N���p��JD���t�7��_�f\S/8Pj��c�0��_t��Hǿ�����~$L��ʍ7��2o$�0[���T⋼�M6w}��W����V�{#	����4�<�V�/ț���nI�c�B�t�~v!T�|GN��+���J��ך���t_g�i�ٛi>�b9%�D��%߻9�n���"�ɥ�]�����H����Kg�L�H�X��͖R����{�&�,���"ѡf2^��.ί���Y6��P�&Z���V��7�?�t���u���F�\�/�P'q��R�RQ�k_��nY���w~v�t�1��qrev�k���nx���|�Z&D�`w���Bp!�8-ʔ�ң��z�[�ֲó�RA&�߈�b���t�,Bf�p���
��jWcP�N�ȅ�O��Si�x�חl�XaQ��[����u�i^�����e��鱊_�k~�V�g�S�xƼb������u�6׎,�zX2�S�g����S�h�b���W��X��{^D��M�
*gDC�yHP�	q�|��P{ʑ�E���S�C�i��Kb�^9�TB��8�W(��v�_.���]{��b�PN�q ���z�2�3U&=V��Q�gV�I<}�2�fQj9��̷se��?6%�����=7�7���[���jx?_]5[��`Fa$��	����Z�3�=�\8�z��]�i�1�#B���
<�����݈=^�D��6hS$�R�İ"���bj0P�XP�W���H?f��
=DA���+LӬ�l��6����T�jKWI[`���徨d��z3�FlW1�q�`�f�ME�WhJ�!�UXqG~d[�  ɑuBq�7�Mf�� ����xҼI�uAe�]LYQ��!h?�㶪O��z���MbnZ��9*h�rA���L=$�����.��ǌ&B��fu2��ӎ���3�0B{c���B��C�#i��D3:h��D��r�e�?i-'�Z�34�"^�،8�\6;ժ�1T�kބ�j��PmC*�1]�ִ�BHi��y��5��|����dA`M(=wTA����N�1��|tv��H�d���u���#�/��TD��u�����+(��*�a���/Ӭb�'��/�k��G3.��q�5�A�xlI��D�.dE��b���`Ć_qc��U��[Zc u�/�T
 �����1���$���a{�)Lr'5*��,<��2¸3ط�C��V��-j�x�\��e�����*'�%�$�V���*(���qiմؼ?4:Vn�͟n�����Y6z���s�u�vJ�M�S���	��Fk��SH��t���U�(t�(L^t�����N���w(n^����U0d9(�F�����ut}�X�i�~��"A��Z����b�V�n��q0�>�7:�H�0��D�#���������?�ߥx�+��m[�0�����	4�G)��'4��8�#�}�����Gg�#��vz7O�Ң����^h{�;�i�(v��lU<�6B���j��n�?ĭ�ͤ����n;U���ݼh�z%B��L�|��s����4���ρ0VKAʌ`!܌�F?����y���8fr�
�A�(�s��|��3���c����jH�9����&$�0�S|V�@f�x������@PIA�y��C���[��=$�*S|	��`R��=E�w=��~�y+?:�����.�dw���l}��)Kr��sIt��J�}�Yg�.�W#s+��Zj�w�B�����.d?�e���y-?k;�R�N�Q�J���j�^��p�W���VN�/�@X�����jM>��t����d�a�e��h���x���� �rf�6�����#+ž��B��-h9�Kw8y�s"^�Up�Et������0�5-E���`�8���qb���o�E���ؙ��&h[OFD�9J�x�O�x�lh��~�f_��{h��s����^<�>�v[?\*	�G�q��	�v` �P�v��7.�����{���ՙ���'5˪��(�c��'aʃe!"�E��xU��D+�	�B��l�����6	l~G�qtd=��#��Q��*f�s�z�O�z���	b�&�&�[�|��������zct�`u�jb͈�zdv91��<�?#ϻ��Bl$�Ά�)y,�cWÑp�F���+�ܦ�U�)Խ���KF�-��R�Y�%/?P���P5��x8˛�ê����5�,���k7�E�c0��2�����>��po�Љ�w��� ���"��}��lҺ�+��4x�W��'�2C��b?��v�,6%r҉�����V�ڜ�r�~&/v�O[�s�hؒ�y�Ay>%��}.�ˍ�����e�R42�̽�X��;���7��%Y˫WG���K��jAN�[�N��'��,h�9u�ڙn(;��������\=��H���N43~��ڱĩ
't�(]���б����@���BE޿���-�����I8�;	���O��.�B<�ȹ������ա����X����k�E��0柏����)VA�y#�$��"8�J��Zu&���(��	�P�	�[A�-�������b��K�-9��
zvCF
ҷ��v`t�U����Mc=���z �6�kz"4��d��B]�Hc�&�˰��w�i;G�P���^%���C���/ΉK:|�'�I���Q`%�� �t�����&�z�j7d1��o�����mT0�}�-Z�R?��q���=��`�sg8�s��QtnH����򱏋�� �;�Z<U��W~�8Gz�S�c�޴h�Q�����)�5B
�������2 ��B�_�$QH�_d����Of��Q4c*��5�Fse��&�̃-@�,�(���W���,|j=��Vm5�����+����,�)�������i�#R�[W����pa�㥟v⮙&|����Kl)F��яV"�ZMΤs����'8�H� ���a�h�8F�(B��p���,%Ly�2���F��RD1f�O����>�8<�H��GV�
J��:6���F���]5qIN!!YW����c�&DT�(�@$4�م������F�s�J1�ǜC$p�b܊B*�"2�����ڹ�g:	�d �)��k�9����#�����AP��R
�i��6�I��響���"gA�ץAR��A.��L<"ڠ���OJc���g�@�p1��>n�Q�4`��9�K������iB�n��y@H<I6��/�@��S�&=�~���ᯔ���[E���� !���O�!��&��H9�YosE^� �{�a�e��f���o>�=0�T#�1oc�d;�|���r�O-6I�����f%׀�S����1���.����lH�	�6���2vi��f�yh��V��ԯ
���i��
F8���>/X�:Bz��P�CI�R�b�pR4��
��X�gL,���xu�6�� �$w��~�`[h��H_Gn�;�	��8���!��W��˻r�3�r�ⱻ,`���Hy�����AYG�x�{N�It�������⮄X�n�:�0Et�Oٕ"�,X�WC��H���&/V���ɟk�*���;;���:��^LJ���~XԊ�\8)3Ǥ�D�J9�G��q�kF��̽>- *u�	h
,ڋg��z'�@�������ᎆ��|�P�H��=Ag3�\QE���M��4�ֻn#��%t-Q���U�B� Z�= .N(��1�H�[�ֹ��E�N����Y4�Y$��-�or,$J�Zi�GY�5xd��1Y��'jGK-mlŦ�/38r�3)n��`�~���t����Zo1�։�e>��~����5�l��\�R�Dx�w�����r���#e�'����5����ѡ� ���R�ͣ����]��w)��Wa���N=�G$�A)�	#��O����B�Y5�1

B.�2�;�n(�(�$V�6"�-N�:/��"�m��#��-��F�ˌ ל9�N�}�K&��X��p�>�dh���3R�P�{��'o{O����6��3��r�,;���)H3=��ȥ����G�9O�S�'�,e��L�>�Y���u����Q�d���q4�]�<vm�l{��H/��G3�@��%�(�e�X<�L�C��\�f��yus���z.�h��7�r������ >�.+o��|2��dF�.A���?�{CY���!j(���%��5tr䎠����sCn�s�����9�:��9��@�㏩ĺ<&^؅��\�b���py�\�]���р����
�Sn��r��_��g�/���*��:̻�X kT��-�]�[K���v�BX$=xZV?�eȴ��`�4J��@c��p�i��]��&d��hj��Ef��a�v�dR���s̃w&L����_���5�V�ї��Ԧ�S��%���vI6;����P��{��_
,3{�[�s<�;qɆ�7��O
��%�Ӻ���G"�4��p.�*�:3�ǾL��3���	 d�!�P�<�
%�84�q���͔Q�n�`p�J�K���;H�Z_�nf��a�
Nջ�����8� H�l�����fÐ��U�ۛZe,/q�j]�v`i�~�`�����*`�C��-����C|9C'�I8ݹr$L���5�D�u}~��myܞ4ym�-{^�$���Ǟ<�R��U�Aʝ�1���8��i���gm���r<�lZQ�
ި@&~١4��#7ća$�3]��ߖ �c�/���*XT�y�:M��Ě�V���Fn���I�O)J�����y�k��W��+N�*���o	�
9k��P;��P�b��3�m��2e �$|��L��њc�;���D�pf$`ء��#���m��R�>%J�n��|��px�89���6v|DKtA�?���S��Т�~��Z����
���iW�H��Z���&.7�I3�m}�|	{�	_\IQt�WN5���]��zZ���Ǐ#�*���I�SJ,��?�{�RNY"�ս����Ⱥ�0�5�Z/�輘�г7}Lͪ��q<e���hTv$zM��f��[Ψs���u��O ��T~�E�U�}���M��l�j��!q׈Q�6nN�eǢ�$Z�-~�ex�*��b�Q�K�,��^h`�=�#[�8��y~�P,a!�~75�b�J�,FNNӤC�Z_�E�b�Psy����r���Q	 �߀�*9�m�����N�p���]եb��۪���ŀ�g���P�;���Ae�iu@pV_�9�4�Fi�*	���:�/����s|��گ�t͚��.�&�g0��a�Y[�9[������P�2JI1���
=O�]�� ܣ��N'���4S֌�D4m�A�׏�0 ����|�V,4|�Q`�1&�%u�$���f5�a2�bF�-.���%�O ~<z�V-�'/,;-N'�eQ"%5d��7�HV�.�A9mdv�HV�����p\)�A�nN�}r���=�|�a�aa�)Rv�0Y�VF`hO������N"flV΅85t�	�I�bT�*�;�9��u���65o�|��B�WP6��h��a5��P�8�.�{��[L��l�����3�$u�ST�������~�:t�T�6��P���ź�Bo��H�v3��H�ZE�H.'O�,d��L�Ot�v�b�H��}���:������|�=�P��մ�kA,Fj �;<�ݓw¨.ہ�I�05xCWy{��I�A� 7оl�m.�`w�j��C�i��7Ȟ��Sl�ݹr�V��ȏ&Tۜ��Ř%�/�$i0)MR����%� ���K�� ��D R�NDB�hʒ6�"�����KO>�4���)8�5ϓ׾?�l��̒�~Y�?��vf�Y<����������̀K��:�jە��A���_�؜�>%Y�TlQ&���G_�77�/�ֆ_;_�����w��',��e��	�f4��w�����,��&�_�f.#H��ɘu/��%BARq��e�$uZ,�k]h	��߉j/z�$�JҪ9$n� �y���������F����WK�����	�dd���d�m0�t���G�/ޣ�*��L�-�q�U/8��-�iR�Mr�*�1�Jlb�ߙ�4)c�>k��}��;G���d�OV�F�Eqs�(��3�I�!+y�͏%��Z�)|	��򚳪�		`��$�zg	��*)�f�R&@I� �g�a��I]줹ŭN!���) Ɗ��`Y���[HD��e��2��HN�b���}�AF�ƕ�#&e�I]���)��3��6�M9���)�wq���ԙ����#�{�'�?�4A���WFJY hm��S�6p�-i����DA�m�o�_�0+�]�2��Y兂+���(�},it��
��Y=���s�s=�sp��J#�F����BW��3�jԕ��7�T��o�-���=Soƨ���ז�V���3]<�KaBo@C��t㱔�r��	��۸a���٢�k��_ �e)R;��	�塊�	JP3���у�&�Ɓ��'�O��(���6
|�T�(f1��en"6O�J����+
���:�2�d�:!�
�� kT&k��DЦJu&��A��|C�T�Mf����ڕ^,�d��`��tg��T-�zmn?�e9 �Pe F��(!M�w��`���o����J9?��SI�31T\R�(T�\�9;�ܿ��W�4A)�9t���SZd�uT~�m���Tb����v̈́�KP��x����P����� ��=Jcp�;;q�k #\&l7Ѻ�K��~��U'[�a�G��`�������>�B-�����#e����fH�yb�Ni1�蚃�`��'{��b�P�@ {Q���aaA��������ZC���;�;h�QP�:@�E����z[�1�ZO����Bn]���(�������n��(�[=��G�C?wǎ�P(�{y����:<��4�"����o �l�p>�/-3��;0I��� h0qj���ZFM�Zw�%*�D{�A;H��޿�)�X͔��2@z�␲���NSyv���)t���r��aBZ��S`�ƀ��\�ϊ�ɇkF���͵�w��Կ�[6ZB*56M�=�	B[bd>je��
��d�e�#V+�8�Fx���$nR�������^�!�+Y�:Z��i���H�?��2�'t��ɅC�����:<��_҃�Ѹ���-8�L�zf��}�Y #$��1k��N��٠P��Jͫfڣ��J@J��<t˜ԝ�&�`F�n�`�<L塌�8M�!\M�����	����&�f_�?��*�Ĭx�u�ֹ�JZ�Vҏ�i/��� >�9��j�����
��
G8���,��W�Ɋ���X������T��f��(!U���Z��Y�S�*|�;��`@=�mX�rr+���%W��B^������i՗��b��Ǌ�_5��ǥ'&�fưI�����3��<ٳI(^Uk0O�Ԉ���vv�x��C>5
7�>��%߀=mG36w�(cl謨�B0��٫VJ^��"������a�,t��������%�[��MU����L�c���؞T�Txޤ]ؽ�[�c�A��IS�7
웝4�0�Ŋ����x0E�?���1��ZFS�a��N�~�D���VՊI/��P��j`�t�#���4��Y�3�iN�4���� 3��{�}�GNԕI7����
��B�a��.������Nӆ����L���,E䵙6ܼ܈Q�|�6�(��Ek����`$�|��/�Q���JЩ�V�t�(����$S۠^��!*��_/F�����z��F8۳�ʼ�������BAd��^;��Q
�`9�H��4τ��v\�xy�9�hC��~���A��`F�����A����z��)i��<�^gp�]���p�� J;����x�l=��m@����0�lo�Ź Ϙ�v�PTd��qUW�(/'���"kzk�;��N�
]��h�N��N*�>�o�'O��r )��ru�I�,
sF}%F�f�!]�<&!�t���SY��N;M��p�J�����)RJ �b���7���^���=�(����������^��|��v�%������x��������t�Qk�J�>7}��x��X<
�N�=�Rg����ï�z�L�|2�u�m��ωe.��f�K{��y��c�Μ۠���V7h�ǡ�{A�	�P}���`��1�#NCH+�����M���% ��7�r�Mj�t�~�l6����2#��^Η�ۊ'�7��ZL����{���'�B���QTz|����1GѠ��~�Q"�G�+(���~<�����Ĺp��3?���wZIx��}�)���?�,�7�c*�j �e$�r�xd��%y]V�t�����QG��Z�l�00�"�K��Ē�s��5_hǻgO/K+v�0隞���m�`�bJ�ěǻ�=>O��.���=d��j|	��~���/W�����5�GA!�$�T��w���#�b�P{���f�u�m�l��g.�kS����t=ְ��ʰ8� (0џ��xNws���r���YZgѮ#�aƟ��d�]A�f.�=_LU��BF�5����=�}N�k�"ʓ���"[�w�O�~�6dv��8��R�}Y��|%iL�v*�d�1�u9�@c�d�~)d��|	����+�q��(�FXa�o!��0����YL�G��S��L70�]Z��L,��'�R?a����x��~͞+���6�T� t��7��>����A9�JG"8 v|S�%�h�Wٔf)?�����dY0r��5����m?CNz��0�1p�U/ב�ư�'�����I$��G4��j�v��l�G�nݰ<f���S��{��©&|�â?��>�v�"�_<��~"��#PA�[��@�[�)��k\��:�
�n�]`���H�P!Gq9���u� ��W��߈ (�3�b���hx:�?�����0?�[��ˏ��xZ:$|=�n�Y���("��
g������r�31��G�(��a�������]�B}M�w��0�_���m8�	�����*��3EC��@r���Vu3o�'Ͷ_�/ˠ�`?77���:�H�/�oK��E뤏�^�
����������M��M-���[��:��mg<�1������}���Ɲ����v-[0�nɯDd@���0��_Pu���i���C�&|6\�׭~i*�Z�P۳6�n8u}M��
DOo�㑘�}Uf/$}��W��)���ni �S ME���i����Է���y�=��d*���cbV��M���S!p�������X��4�8i~'�57b����^ĝ���r�Cɱ7�X4�.ߥp�(l�&�ޛW<���Vr�Mہ�F�.��&p'�z,�LH��CR!>Z�ą�3W�%��Q�b��ذ���yz�deW'VxSY@�(���zK�$!�/A\ s��:?9-d��ϴ�n��#n���^�&3����4����iΚ5�I-�.�'d�67��.�Z1[��B�,K볃��*�Q�2�q��P�< CMmn�}VÁ�=�7����^N�QTM���N�YL]
2a��ѕ/iKOq��A�ckv2��;�=�k�եI��,a�`����k�g�F�Q@(���:�R����������:|~�����e�eUZ��}B�S��	{��DwtZ���yun���M� �߯�ߝ9��VTw�2���'(JDq$�(�!4�d��������Fܸ��%�,G?g^)Yl"%J��d�KQ�J��Q��E�`nީ�!��O&d2�=`�)a�"��Pt�V�:�0�
��h�x5��Fa&>VR.���z�:�
��񠎥�9���=��=���;ξ"-Uh�ʰH�ѭ�f���PB��0:,�ޔ�-�u愥T�@�V�4�&.j� a_+[���uP��;0��l������}91�S��Yrn4�;�)�,��WWn�d�?�ϣ��U�M��SHߕOAtcɂ�{�S�{J�a��/Z;�!밟��Vo�q!HF�����g8��?�G�`����.n%���M����ɏ�zU,;��`�GU�R�������k0b7�?w=���u��4�I�����.	�����	�u����o*�E�'��8�U�#}�T�pͱP8	G���̊$��5��n�����/��p�vӊ(���u��Rʱ$S��^̱��@(	�x�R"�"��Ž�M�/Y$v7٧��|�%o6[®�gE��A�*Z2��+�����ud����H�W�(�@N�}�|�}��7�h��s�����Co�(�����*ʁ�G6/�.x��&��g���
�������*$���>=_O�*<4����|3���7�	6�w ۝��~�gp�7'G&^A6<��a<TKvDx�Œ��=s8�����9�B�ƅ� C
u���g�xփ��bc¢}�5`�~��n�_5O�E;�����8L:����' ��?f��r�w���R<2�jEc ��L�j`����*
6��f���9��$��|�v�w��ԍ쫑W�E���`8���{s�J�/�ma��27ӫƌY�Z�xk�s�
Uvq�.�	�Ļh)�o2θ ���ܟ��C=��F���8�猦�?�4�π���Y�=&���(��f�-$�%A�x=�(Κƍ�$�lf�볃Ni"���+�
��c`}Ч5�]+$0I2��I5?x�שE�9�R���(��QP��!�{ -�r�VA@�;�C�RdN�����.Q����!�@�U�O������Zeln�;�����7��d8^��ɣ����ķ��eO���L���6�A��WE�?��Y��+�ٙg;�}{��}�[�I��	�Rj�q�'����7�6$Δ��yL�cƲB��#!umB�J�1�g%i�&�xsĄb��J�C��V�C�b��}�v�J�G�	�R\���2���T�_zN�����`,�3*���kuJ����O�
���L�a��tL�v�[�ܫ��A)��)MlA� ����n��1�a�`�ihp�$����n����[l�0l�|�|�!]�����v�@�/ͼ`��8�	�����?0w��V��qo��Be��|�읶w��$���������N�)��٦?Ӳ�R����1P�wB%���f�*� �y�p�/a���^d�B�InNh@%�fmb��
	�#"3�	� �}�{�vA>-]�n*-��uK�L����Nʆ�8C�V�T�?s���|��q�C�+g��绀�X���نjQBu75,6�M���S�*0TK����Y'q�r�7o��~��^��e-��ѩ���sV:�^�4�7�18��m�j9��ҋ���.�$��#�y���Lq�f-�3���<li!����uBm=����P��y�Fgk[Z���w�u16��ۻ@D�t�t���l|*��BU�N'�c=�R�v�B�v�em��]�z�Ptl"n��]k��e���}b�f�C��)�ܟ �[��&@��C0��XAV�ȹ���"p4�����
�m;�>��"1.�0��?�� Ic����	#Ǧ�[2�����c]���k*O� M�TB����s Tğ;��Ocp1�0��#���E����+��(��y�$�(���NIEq�*���~/\���[�`��h��"X~z�ߓ���k
��˃�����l����&�F�'2E��~�-��
fZ-$�8��d���Q}}x��M��8R$�Dԫ�yI��*�d���ly����r��Y�7+'��qqG���ӟ䲪iZs��ۊ�O�:��A��n�ŗƪǝ���8����0Kw��C)����:8.��q̥��s�Lg�!S�?i��)���.���%2��>�yq��[<jv|�'�_�Wk�y�}�n��f�%��b�`+��x�X�/����>F��T-��ߗ�QE��QT���yX���s2`��;�Љ��}����bI��$�%yvۋ���m4`���S��;�-9 �8
U�G�VYy%������/��7� ���$^~�������f.Tq���*���Z�ǊL�����͐���)A��\y�/"�����F�����y��x��4	��'��ҿ5�Xޭ)T�W�����t*6ˠ^cv��0�Ǝ�����q���oJ�/M����\>A!I�_޹��8�D�-�Ѻ[��y�vȄ@���wB���2h��[(���>��|BT7���*s�Ɂ0��4�b��&J��q'JA�).�5�%�tXb8�(�& ���+�?G�!�x>K��e&nʹ�{ۛ0+�7�n�M�_�l�إ�ĕr�����s'����&éS����������4�h���j�87����Û��K�XK5�nf�9n?"go�b������^�b ��]�,Y�O�S���e��,���,�,	�%�%c�$t�O�H���H�$:�Xp|�}[vSK��Mf��Tg[
�B
���ӊĉC_t(�A�k!c<�d$t�M�u&�1��g,��2�p�AI�zt��kT��ocK�',��L#��ѕ)�k������1q.A! �6�P��&��˄Rͽ�SH?O��-��B����a���&ߘB�he�Q��4G��ƩL��ؾ����=B|9�V�3�Tϔ���rR�c���7Ǻ,����y8�*mI����2���|�:e/7�yQpBW�$�v ��g6Ux
c�CA�m�	�=?��y\`�1M����s1H�ߜ���F���"NVڳ�d�r��q�Ƴ�����.��[�"��[*�b�X�%}�1�����t�ٴ�v#�I��<��8 �؇� џ����,��
��b�[~a�fh��j�YRL��u�[CT�����w�֪] C��'C���5��i�zE�G�g4��z�sM��P�u������Okm�(g�"���;ݏ�P�Y��"��xLrY	>�xVD�$�f��^�"'1�l9���bʪs��7
��c+wl�;-�����Y���?B��'��D���|�^���K;9$��n1<Y�>q	ʖz�cU�X���+l��������٫�n`3�׼��v�(�b���>�28?j�;��������A�;�Q�6���9@��]�R���;Z�7��I6_0��]�)U���2����Ϝ��8m��s <+t��Q;�r���3�P���[��57_i�r�<,�B�(��y򀿬�E{S���,���u����7�k�"]�ÝF顂�	VN�����|!WGug@m�gqN�����62�g6Ţ7�� Xq3eFT��B�����fB��黀s��������r��S�r&�p��G��*�: �e�����[�2&��r|9�5p�^�H�l_����^��]H{��mt�ER*T�(["�X�@���H+�܄���	2 ��$�b�J^نn� �qP�(����M�|�l�a�x��@��,*y�r�<!F��t�|;��U@���Q�����9TP�`�vv``��}	�h�_��Gj,��.eJ�+Up���z��6����|h���'��}Cg��o�.�N��~�ܱ�N��\{�Qc�h�YFְ3�cGY5�p�a<L{,dv�`�8��G�n*�-W�֯����=�ƜRy8g��D��QۺN�@�m�!2��Kz_%i(�Dd��;����Ǵ�V:�C��O�ݟ}Z�S%�ouCC���W��bRk�#٣`%��D�T��wӻɮ�v�Ц&n�%O�}���X����V1��� H�����e�U$�}@(�/q�8�]e�:�s��������g������y 0=��:aV<�k���8MX"��
��	8ߖ菶����+��m&'�Z��h�ܨ��ܼҽ�_�Όro��{�O� �@�(����ABiA��^-�3ղrJn�-Hפ��ר0]G`=d9AVf�0N ��0di�nە�<�ǔO��Q�r&'�|����օ��,z���#9���=��"yLތ�$@_�E��,��)/g���7u�����~� �D���4�u�J���`�4�ۚh4<�pTc�9��A��
�o�^8�=�Iч�0B�[𘲢�7fcQ-�b;�`|��ljD�Z-ɖ�d��")%f�[' .���2pu��U�i蔆r0a���Nu!�eI�V������#t���2�+�B��U%��/��u-�k���,q�m('�/�hyU��������H�{�매Qo&9��ŕV�����K���[_@��^���jʽ�:�g�:�s��i쵩���S��m]����@�|9K�6,ׯX@븺h=���HM���uړ�I�RM%-p��<�����'@��;t�I�4Z�?>���[H͉a�h\�a���ou�^�N]MW~�
,/A���&�`̚>��/�;f��5�$�w�ϩ�{�b� ��F��J������1V���khQQ�?|����Hc�~]v���I��h@D"7*�FRgJm.���NV�S���H|��a��Q;�gQ�\nȔ��T�ʻ�<���=��q�!��_�"u��+�ˠ��f�6�r"�+��nܖ��( �M.R{a{��܎ܣ�Y@7���h{��)R�)�_'T�գIEoluZ䊂�R���:5]�:�2�bRM�R���Ȋ���3I��~�8x	G|��ֳN��k����.l�����1�z��3�H�ZӃbwB��"-�;�h�>�3��o�QY���Ѻ'q��u������lcA���\����a���d߽G���?FqjSv1�2}��:ٽ�Ίf:M�|��,�˶I��u�PȌݾ��o>��U� ���%A�$�'��Y��~䥑���w��UVf�2�=v]-J�Ό�Q��X�����S���r��sj\�zC��4G��7*���x�{��ʡg��图ө1�:b%�*֬��M���{���q�`�9���%���tE͗O쩋�~a ����SA�:�V��lB���O�j�]E
&�S4��w|���DU��o(����N���HK�,M��t���uܥ�#�L�B2�~��FQjpD���eE
[&�F�x�".:;�m<�fØ�����t|��n����ݠ��#��K���%��P�=mD~k����,l}���?pBJ���0�i`BD�d@7�(�H>3Q�pЉ3%y05�l)f���G������97.$6|�)�͍�yգ�Ձ6}�ּ�����3oGP���
�"m>^ex�%��[)�����ي�4�p����4I�N̐��K�tb��G*�O(jGT'�����X,8Ubt7hmZ�R��@>B��ܶ?��1�U�Y?H�dI1�����g�ö	Ȫ�Nh��`]�������s�c�Xn��]���@o��tym�؄��\QbU>���z�ȼ5}��y��HhX��׌<�CSF�t�:H��c���l��w)��"���l} b�5h�����g a���Λ�v/fm-��(��7��b����H_�o����,� 3���[ò�Y��f�ʙ��0��]�7�l���#���[]H��d��K/+�	�&G�B\g��{�߲!�w��v�e��IZb.�R�sk�C&D-�,��:��]���ަ=��TAB�r��������:XyF�̸l1ebi����^�{]:�`A���l���G�"��Йmp��T(N[,k�)�֩/��FC��"ka�22��gsJ����������S��@%��!�5ɥ 88<��э�>��5�^��Y����6�Ek(J���=���yX�f��|ۚ��+����<�W�G?�
�é�*���Ƚ��UC��sTa/�ͯ�ƔD��c�-$?��4�_��n02k��Z�S����i��� �¶�Σ��9`��iN{��.[&b���[`x�� ?ol1�b�����u	��--m�!J*�5#â�9�J��{!��w 뚂�;���}^䇖��Bmޒ(�<~�0c��
#�s��>-B���d?�9��սa�x�.&F��	$�5���Vfjy�G���n��흙��9W���GQ#���B��Թ�� g�j :N�s�(2 �䀺7�꠩~�v����"7��`s���ﵟp���^����*f��֌�F+�)�J�gz�sӭ}���w��1��m��GR�iY7H��=�!dA0j�Qӫ/ )P	�����yLCjʌQ�R�=����,swt�L~$(�𜨝��9�9ո��	M����G�����k��tJ?��ݎ�i�<!"p��z�`6�����h��Rai�1����ڀV�2л_���\�	x�I��d�����fup:p(����������@���Z�_�OO������:�R�O�1�wVa/�<S)�@(b9���8d��;�d2?�EN�Q����h���W�+H��zj_�����. 5�K�̊��s�A-g|y;n�		�vj��ӵp�f0���]Md
�oF�f�˲zYe��o$ �blB�k����v������DX�I�����#�ᄿ�	��`�nz�gB�)�m�-6��ϱ|x����b(���q��YL5�� �o�z�	�O�������*6�R��pܠe�x��դD�\��Y���J���\�߲1{ �h"Ål����Ԕ�@��**�� ���\�ag�J���>q���HP6�,q~����XL��C�Mf+D@�`Hrw�����ق�R�X �EҘ���O�}$�K�M<gwܚ|`1���L��M5;��5�/�S�:q��󸌰I�_S����-AM�$�?he׻+���۰i��6bC��U~�0�+D�����6��:hxY�=�)���C��c���ޅ�d��%~E.����:gp.��V`�78᳧��m���D~� ��IJ�ԅ��2eH��!7�GS�I�*�m���V
����l��ND���b���ޡA��[�U��lP�Og���5
��U*�#_vQ�Y$"ei��v7/�;Ea�V8���%2�d\��������G���3�@���+��(z�j�i��̻=����r]Fmh���V��:gRU�f,o�ޱ��� U�u1�;E����*����qM���z�P�i.,�I)�REwc�|��W�~SL~qn���nW��FPR���f��D0���A�_p���4��4�)th���b���/-�5d����U���+�������m���e���tnN˘�ͬ�Ljp���;�~��6���m0���7�a>�q��xV��^�0��d! /��9�

��INP�p�AzH�ڠ?��e�[B:VT0��4�GD��X4-p�]+��[�ՏJ��Z�����!:k��Ѯֵ���^���+�ڸ��_uQ�\���WY)���Z�{{� y|�ר!���c�G� d*�9w���H���B�����^���+�zO�������v<̯�k� sKL�ol�T���y?�6f����=��/?�����W.M�aG����TmE�F+�mzyW�o/T6&���;W��h�p����8��G�D ��?>Eb�tH�����h[֯��G��T_�HH?U������'�)S�㒉/.̈́�����l�_K
��e�Mz����x�>���^��?���Y_Hhy��e�.\r�+jg2wщ�S�7\�����[�_L�F����̤��Z�?���?�3��S�FW531�y|(C�,������e�n�z�nA1ԍ�M�K���Ks[�3�
𔾥�rwU�v�R�/ȯ4lsK6!d4����?#+;�Tq�����tVO\� r=	j&�H����F	(�H�N�7;"
i�!(�(��0]x3�č��(�K��Q5Ϛ��b&U��9&L-���8'��;3����"Q���BD����Jdv���EoB�y�K:��6X[f�:e/B�vqƢ�MP~�i��_M���\�0����SKi�ԅ�W�1�4������Y��	�m��_%�9�c?=��c�B��3;LA
�y����'�r�5N�m�� ���7�o���p�;/���:����:��m���z�����i��Z�Β!e��b�\�����Wj�����x��ʥ���;�1pf����хc�\��O	>���Vl��l�t��T�Y5�������\1�'�c�h�ߚ��\X�PI9�6����p�P:$)pLʺ`���ש�O��XT'�e��r�A�
��Ұ�!��Ṽ�^ٖD���7q��P�R�ܦs�Ip�St�x t=�0Oe�	�Ơ�g��y��.��?Q�w�E���'Hj���9��2�s��&e~�W=��GCn��V�!�rC�M�`I�:�Q���Fƞ�W��e'���[�a�S�p����!��2�1]���);`�g��8[8�3�'�,�EI4�T�yFh0n%�H�6!t�M�Sо��w�;���z�T ��
I����bQ���A�?��ˡ6�<?yz�����nMj��x�W&�k����l���Ng�m�yj�4��o#��Y�c�Wv����D��Q�l�}�ųi�gF�(2�U�o�����)!2wII�i�NU]'��5Ƨ�REk*�$��,8�`ƈs�󻥦`�ǜ�o�z�o7�zw++A�'�Z�zN�o������'�a}�KY���0��#��p�:�2�(#'�KGS����+6�P/�9��[ҋ㳗�Y�F/���e/���2��XM���&��]��ҝ�$E\�*��MR�Q�KH¥9�O�}��`�v� �*+���G��*u4t�hH��L�k>p���K����эL��z��u��T����!���-�$ɬ׍�۳���QS�p{U&�K4DKB�8H�r�2II�HE�r����{��@����K�͛�6�����˘i�c�%'+Wp|=wpY3�QX(��ϴ�ZӢ�a�(�ݫ]prA<�Yo�jP��f0B,t|0�����;�=�I�X���9���6e޵:��!���W=��:�\`��'/k6������VLn�Kdp���Co#0�g��թ�$d��L!�;4
� ل4��󾥭5�B~e��G0D�)wp��X�qjJ�����;��ɃҞ̭�K�6w&5����3��iQ��^�&��]�ѽg��.�
LkMgl�ޙZ@G�þ}����½��x�]�V~�NA�9 J��j]"���h��,���*�Q�]�m����:ޭA�G�Z|�����^��v���V̕�2$��P��FB��&埧py9C>���
���k��S.��l����\�~#�KL��"�5
Cs4��hq��~��Q~���%�.�G������F����I��l(�}�S7�b�sgS��ٕ��Ġ����7R	�Ǝ>З�¨'NtC(���"���9u_	d-yM�"��B�x�[s��*�8z�Lv<�L�y�M@D���Q�50�e�;�_��[NNU&�B�����P[��@�i��E��Lo�{A�j���og��.@�
�K�B�o`G�G`���2��e,M�1:���9.�p�ҷ/�����>�1�N�Aq�؈m�\p'y��(me��u�]����Y�lrr��h���	��B�"L��QdgO���7��.qMI@v��a��f�f������m�n6Z�4U}����\��?�U6���g+�{��Q�S���PӨ�!]W�Oϲ[MO�3\^"�I's��[�%��i��ںD��i�R��q�3)운ڨ^��6)͝��N�g:�t<}(7�`6C�聰��E6Sd��!2,Lc_xY�_Nwn3�^E��7�X��sZ&�\|D���cw�O�B)��r��R����DƐ��44i;�$�����8��vϠOņ��c.qWDL2J9�s�Ϊ�锄$��}t���;@��08-쪜�Ԟ �<e6aEZ�g�m�&G��SV��/{����K�oe�:`Пf���XV`R|��j0]�R!;�05��;�1���(��5��1�R��A3N%�$�H�.:��F�a�§ ��K��I���
�|�n2�Lȓ@A�ǣ�օ�N&71���>���i�G|�}�3�*)�{Y����z�A�y O��І�qx��<�¦�?����>6q�[�18~4����� �����y�t��nϨ�D���A��J�:�>�Q�|�r�\賗�,��B�}*7c���9���f��2ђ0͈<�P<)Q�kbe����%�:a���e��'�Dm�|�.4���Y����{����\�g�
K��poN�u��h�A��U����vĕѥL\��)���/A�6 ;@�Hj��F����c)4't��w��|Pō7�Ƃ/� �T5��k6�kŃ�ȸ[�FU'LrK��l˄w�d<������@���z�}(�a�1��O|����M�|��̸n� �g���ޟ�1='ܫ�%�b0"Rh�������Y|���� P��/z�\�@��UtuҔz����xb�I��ۋ��~�]a��3q#���?��ZH��;����P;����ez�X�Y5Axr�` ��!�'97������0���i�����.3V��K�j>!�0C����D����ѻ�W�P0�A˵��+�v�:�����2���^~w��.�����ӗ���k%2oj$M:ϊtt�^G3��8|~���=���C�q��r6�RjSoz�����1��6s�C��?3����e{9��~�i���=˖��ٶs%����DCaX�GVlۼ�;s�+=��bDk��0���[����|����W3\�-�Rs�gnIY� ����O�~��-����N�}y�6��d�Sֶe�
�p��o�{�E��f8���M蘒�K3ʊv��I�|-u��X�|d�J�O�sXfYu0��C'i��cb�O޸L�'@0x�yn�Ȝ��-]�8J�7��;4���9�����r���@�������"�Gіs�)��E�%���ጾ$��{�r��j��4�`]`��D3T�H����+���v�
��*��'&��M�Ǟ�J����!����'E�-c��Jws�0�p�֬�j$W[���>-�{1���ж�s�Sl/ə���N�\�}���d��K�@ྲྀ���A�^���]IQ2�Tm��Ł
d��
*me�곙�p�`D#
��N���	�	�6@��� e���BJ+����� P�]T�2���b�f��"q��@�B��nĈp;�fEL�F�=t�O��.Σ�<��<��Q��2 �H S��Ҷ����_o��ӣ�q|��J�8�~f[����V��3�g%��YL�r�x<)�"�Ǐ�}����P����45�NP�i�k����Sׁ��6	Ew�=ܳ����г2�b+��y�W��:zopU�Q���+(��=Đ4�j>J��&�ܐn����A.�u.�<��=qÚ��$w��`�l�{�w��7���2�Y��:�ে�k���K�&~�M*"���Y���Z�� �䚸�NІU4�E��颫�UB/~��F��l�!:��(Y�@���k=���������r��wV�sc��X}�/K�W�7y��?��EoC���H�Ӝ~B�^�����ykl6P�h9��%"n�պ3L��T�6����.^x}��
�1p�6��n
�I>�3���D�"�d��q�N��ұҡp�Q@��m�3.b5��cO�G�-��3��ҭ]��;��jk��n��կ�OG;N(\�=u�����$�I&����K������s0k���H��#��I&.ٳ�k�l�ZT.�E���HK)��$�P�咟5����z����-u��_��6ۻ��0�WUo���dhw��Ö��ȭ�4�н�h^N���&�%���SFJ���P�g�);� w#�_� �޵���k���Rh*�y2�hn�@��+���}�)[_2S@�H�]��A<�.+��ɤy��@kw�Y�zA�f��ͱiwv\����,�6E�:�OI��m�{]��4���\Z�kR>,�c�Yg�N���cP8z����ы�|�X����>�����u����;<rv13���jg�[����lQ*D5�83Y��qdv�̆�����dI�"Er~��p��=^��h��0_��E��n���O��z4����?��p=���|����K�;^��(��"SYwB��eܟ��u_�1�����������<��b�8�P%��valW��xk:���V�
g����;�%��,����4�K�ݱ��~�����`�����;��e��h¸Y����תJ��/�#���O���!ރ���r���<��~~i˰&Rp$3�����������W��Y��m=b1p����O�4��NI�pR�Ϯ��L=Fg��l�ǝ��| vs�?<�V6�D�Ċ�λZ����^�ޛ�
�+���hMZ�L���g�M�N�����U/T�|!�+"�uк��K��Q(�$�r0�-����A��p��F�"���Lp���_J6��Ԕ��|b"=���裩C�	器�fV���V��y��䂾�)��#����s�[t��(zI�ua�i�+1��|ݙLq���T��^�*�=/yF������v+uX�̍�!]�?F��s>n@L<�8�d�ۿ+�y_!���~aq
oڃ�BA7/�Y��HX"��8��.z'�d�q����g�շ��H�K�M���t�(�ε-I��	���uq��1u$��n=Bg�d�^/�L�@�8�l�����K��|�%�h4����B'�.�|�ה��M���A=w��.����~�:�A�Gj԰�*���w<�i3�l.�S\���=�#�-U���=a�j�o����H� ��# 	_�/��Ĵ�H����b��v�YONC��5 ��,�ji�����e0Cys��*y�(`f[e�ȩIK:��~��҂�b�t��=rԢ�9�{S}�
D�/CӒ'��]�sq.��*���pF��1>L��Vk�x���'�8謄ۄ��R�[�B6ţu�㒔3hC��M���$|g�P�4/b�q_����}�=a.�}��d$v��7NA�r(�������71Uգ�q��:��e#�X�snXl��gɳG[bsnM�#mt�^a�An���|�.Hs�Q��*�d�C΋�/L��<W���3���Ǯ���S��>0>��[9��'M�G��9C���M�z`����9� ���c�l������I+���q�� ��*��g�4�N��Ik/V��5�e�r������i:��3e��{�Ԡ�03)V@�Tw��"�듋8�Y�נw�NA@x�D�a��g9�CzjNQ���ܜ�,aL�"Ĺ58�[�W1�c����^~���#AJ�C������.���E��7���.�k{�����-��>��{�(�Y�m\\l ]$m��^��F��nk{��S2��~ww;�.��ph����;�:U��]���枚IT��ϵ��,;n`]@�=P�5��?uR�����#�]�u����Og>�Du��������7E��v}��MwO�'�`����+˲fˋ3��u�z���F����Zᮔbj7��#��D�����r�3oYn��Xu-m\E>�(4u�,6m?FK%�}������O��:��{8c��5PWH誝p�OثTV�v� �V��U�i�.����7����d$��D]�1�g՚�Nw�Mz��4������&��g�
�ި�8������m�� w�I�'��ZZ	�F6������ȒEϚ��OH��5�RJ����s;��7�!n��ImD����&��{&��i�����t���7_�,��Э�?���ǋ�?u���F�=.����1m��d\���ֻEy#�ϻ�f�ŋ���K{�����`'���
E)�|�W@��_���tu
}�8�c�1��y4D�p�vc=��J�IY�eg��/��cY�����"*��K��R�9�WMG�����X�ZtNN��p����
ygaw7*<W���Ș���Yϵw��K�3D3�IQ�W�o���?��3|c���֮X��^���Ӟ�̇f���������V!�tIėd��uu������S\�W�妮4��B%���Q>g��F�i�*��Z#D������o@P�7�
��	|oF��,U9��ۃ����e��;��<ao���85������fM�ʬ;��R�x�͙o�S�F�����1�_��2�י]�Xh_���e�`��c/+G�h�
���Q��ƃ�@xH��e�����~���T|�v /�ŗ;v�J��|qHè@�KF2�Sg�i�P��K܍ɋ����g0�an	T�w1�ԩ�(�mP(ͣ�����*���(f.��&�c�y���q	���E�8�b%������ 0�V���-��ƚh���>�["l�QNBt���>"����� S�d������R<�y�un�Z����	P�NMيف�f�G9��&|7�\�(W��<�ш����E*)�jҀ[ʓ�A簉7�`Q�$��C!PE����T�sq�ǐ� G�IנT��ґ����H��S�_��ב�1<8jz��)-�fIƜ�.�����a�\m���/�����J��F�AKFD�SP\ȷ��UrZl�Ⱥ������8�iNf&���op��c	a1L���3`�G_s��Pd�姚�tӚͭ���T6����{����S�,��<cxW
xc�5�u�cS0Ii�K$3�4.+u
{9�q�[4vX=mpc#�7� �2B!
�N�(}�E���F( g�Pw�+M�h�HG�G��� ���P:���SU���~�1#�W��>�p�ph%}��Z�Y�*�f�\�p>J���c.k���F�
�����z�Nu��w[�0��/S�g���ǛW\�X��.����g1F��<U/U3yǳ�7c�Z�\�V)�"�8�e͈�iؗUo�<�\�]X��PcCJ��U�S!CAZ-�\EQ��V���o��u�m:�>�\9�@�C��
K��t�hSqA��a�A�{������MSu�M@!v�<W[L�SSQ�82��+{ĳ렀�0;)d�;����_1�w.�F�ZvS��iE��M0�K*yZg���'�-�
�+R��.8�a�=d���8E�c�U���'��\K��b겪���Pp�4f&�M���7�Pپn�V���pK��&�x��}��_���Mp?q�N�8/�m<I�i���Z�^gr3���E�A��dp�ˀ��⬆'�=�s�~c3<�@$�%� ����ayO�Г{�9(��S0A��k���rJK2C�PE�3����yh���0���Y�#jl�b�	L��pz{=i�����@P�ǥ` ���Dx=�k��� �4D=�}�䚏Xo���ߎ0��E�@�p����TIHY��.�.�k
$ N&p�;��y�a����)���c7��HB�� ��9QfM���s��!
w#�h{���V͆�1RD��/"�Y�Gl�XǻZ���W�\	���|��ZUH�����������Y(��~�_ w+���*\�w����[[�}������!�:md��z+T4~���Z@��m�W�9�zaR���V�L���<p!��SB�`nla4	h�q!�Ġ(�Kt=��kѽc�L�9}c*��k>@�QE�٪1��y��ǆ%�����˚�dN�d��o��t�/�����ٲ�H��е��z��Oʦ�r*�-��(�|�}%Z��H���ߡ_1r�]#�.Nwxz�V:L�q�����t���	1�*0�3X,^��F�=P����:sJ0�c6�k�G"�B��" c�5"]<����0v������Q���u�#C��1���ۇ�h��Q:�Y���Ob��\-���I1�i9���yS�qwlK��]���A��#�	cG':3���~P7��x�J�6�EV�M"^o����Rm
f�Ђ�JFC��e�J�h��A$�)YM/f�����{U�HvJ��-X6!�y�Xz=�ig)E6>�l�����#��e��@�	�����4�vSVT'��/|�hgjG��ԏ���`ؗ�8�W>b6�#�[u�a���V$'�u`m��I��.��lә��bB��}b�&�F�;;8�KA�E�4��6�r;X砋���W)#�Z hm�p<�A��T�qb��a��d|G�k#����i7�0�E���=��5������t��K����� v[;pۼcn����Q�Y��G�R#�!V־P�}!ʙ�E���=�\t��jY��+��LI�x7�i�{�\Y����eo���w{��iI{�~ꔩߖ�zXv4ZZ��b����)cƸ��(mvX_��7��M������������
�y߹`��g;<O"�1�G�/0*������K`T�jP����M�Dh��^�:�I�&�>~+05�!�P�f�&��7�-L�K1�4�*5�a���h �D�+�gn���Ӯ��8f�y�_�9N�M�m���p��x��q�G�@�G�Đ�/I��
9�Rڒ@~������jN�������K![�.qLb�Q!j��CjNE��AS �k�
�]��i~�^������=1�B{�bl�X���vt/�¨\�1 F���wn�Ǫb�%1��ڿ5P��
J�4��L�!� l !��o��7���B*$�ރ(�	��"���rnY���$	@�ב�CQ��c��U���(�����ӆ׋�X��_���VQ��K�`�y� �GC$�l^��]Y�U,d�{KE�bi.�E�Z�㑟��҃-4�	h��ڙ6S;F�N����g��Dz �;N�� u4�u�������*�(m��;��Do�s��>D�}�5o�/�,R�ʱ�)
�HH�%"�Ҙ��y4�Tv�p�QudII��*I�`i#��_���Z"۔���K��b�\�c8�*�����=�E?�l�Y��#�>@kMڈ���˅{?�6�?_�����Qe(%{a��M�?o4B
���}�Z�U��oܪd�UZ�w���t���]��θֻK�J�c4z���gZL�@Ť��j������׼<?S͆�l��ç�H}�l��!iX�q+�<��A�0�$
w>�~]��(
�^u4�N�_�^A��,��	^���0x�<�GZ���'�H��5�se'hk��ɯv֋��R����J{���n��8|�ʧ�y��?��*BU�<��so
i�!Ϙ��v,X��q�ڄ�5M�]������䴎�xOTN���5�H�f�]����,�	�?|�b3"yՉB	���-�s.ز[������~���ߖA�T�w���n���s/hn����C?�H�a��r:;T6�mr��8"�hA��7�	7��Jן4�!��3?��1��3�K�C��챌.�q��~=�<���疷[8�^��^u�W���P��&:�%G��$ir�Uf�ѥ�s�ܞ����Z��a;Ȁ�"�r��b@@��R�:�m�[w��v��z�X���bhT߼:�BK�VO�Ę/ki,����F��4�Q#�j����NKf���Q�����cArG>�蜪����]M��m�n�����{+w��v��9��x`�0l��7�|St��tM�ӫt��#�݋���0��%z6�M;i�������R#� n�"�w�q���՜��ܽ�@����H��qds��m���v��;��=��v�`��y6E8p�\��բ`�d}+���ϑI6G�=u6 8���:m^F�@}[]����N&N�e�F���@�R�F�f�2�[�Rrn�6/��J�	G�s��TC�x�^�Y#�=��b鷠w����&y�}#�zpb$#]~��J^(��@Ѣm�/%]����?�K�x���4E�S�O�����>�93j��|!,6���E �c�pg�^�s�_|�I�-RV#>���*�j������̳�Fn� J�v,nl�x|G���/0G�-6ȭ��%ٓ〡��w��*�����4��� i5���qz�
Q�g�l��Z�W0�G�H�ξ6��uP)�C:��M�P�'���C��׼�h��(Sj�G��C��쫠?�A���E��Nk#�b[��O�ONX�Elx��]nkQ�*0�E�n���̸�`)���_=���l�$�shb��v3X�ZcnUj6�ce>��4��h$�\� �(K[�����Z$ɱI?�*F�;=��S�w�XT���p�1��	X��O�U�����QLmi��;(�?A2��&p4yOz��Z�抎�t�G�a��� (i���Ť��*���߻�x~M��~�^�~�"a�!lJ���W�	�9L�0x.<���g�S� �Qt��W�-e�%��[hF9r|�W�o]�y�{a��	��OF�#1���f3�o�"�_z��?tJ/[vk]9�έ-�����.� -�����y>aFY��;9�:���:��y�cO�^B�W�a�&���nX�i{ �N����	��C�5�R�� "SR�Ʌq��G�K#���#>����O�
��1�aom�,E�%F"P�b���-��{�D��4R���U��W��O8�� )�� �Q�@D�6����'��ok��{�֎[=��,Dӵ�����z4��fH;p�|ɜc ��:gQ�C��պzn�-ei]�t��:�}�d07��SX������*B���E�����,�u�C�3.8�����������=@Y�f����h�`ε�4U�O�[ ��������@uᏨ��(�����Di�I�+!l��L�'��h?��%6C��g:SFN�p[�[�鮞�R3�0
���(?/ߕv=�����#��$]n��i��lG��o*ʹ�/�n:�nA�"m�!����>�s
��h����%�2��VO\��2�G�W4o�Cpjs&S�@���}�/��=�N��?�ʟ�����^����e9����I�� ��2���p��h>ʡ	�8hM��go� L�ێ��如fF�ʄ�2���-ip�����Ǜh���ysD8�d���b#�ĵ^�����;r��@#yw���>���?N�@-e3%p*�U�������Q���
c��`g�x��f;�@��֏S��M�
M�����gE:v������8�rRv� q��g�4��x|J�	i�Y�ݟC����`M�l�_�y�Ϯ��:��P�Y���S�����x���4[�
��9CǣCA���U��#��'+P/���"#�B?��>h�I<�ɩ�Ob��s���މ�����2#q�@b�͗q�Ur@O�:lc#���F�W�I���;����|��B�ij�����>�����Ph���O4W<P��~�IÑ�H���a�i�:�*���yl��6,���.�i$�4�~3<�xu�!���%(�sJU����R��3i�[Ȉ%!��0qq�aj�9���A��,�I�ͩb�	��E��:j����s��煅.!λ��K�2��pa���f]A�d���{��t��`��࿈�ߣP�M�~�r��{	[�	��4{�I�������<|c���'�wF�X���%#��9���M�6S�	,"l;C�2, =%+��&d��m`����I�b�P��{�?��ӡ]�$��ѢMW��˾�&?��(_FǶ�Ln��D,�O_XG�nC�ۮOIQz�ƚ�+79[�;�nÍk(��$)m��Q
5�.��h���f��X�a� ���/���#�{�3y~��R�E�Y�L)�k}�,�.�3w�>��d�R��юl�8�=��_֦��}B���R��^�7�M�\�N���<x���ɟJ�A.�V����Fq�N@g���]\W���˕���ڵL�6�O�.�ff�,������)+2�q+��i-Z9��^�Z�θ�UZ �(�0�߁[y�����7+,h�}�z��Q�iNRc�`�:���@<�PM8*yձK5\:a��VO�Y�����O%��
�:Y����ヘ_z�)��)@�BL+�fa��̩#1^Л%�1'��CZ�zw�o'����֏�b���R�j��{�Kwt�FNF��2���p"j�t�E��%�t���-?.�BL]�?^�t�4�kV�N���i��"�)�Q>��dWAI-ט4�爉;�w���9��p��{BLRF�o���b�TGl�`XD��	�pU���6��"���C�p��T�矊k�on�����4����M+�T�)��i8)l�t.�1���ͮ4�5��T�����&'_���Mq�k����M?�\c���L��!#�Wm���i�8�T	�`����-K�˨i��聳�tb{��4����aFN�8m9"���^�Q9V��M���K�$�.����b7Տ U��3iMk���fǖ@g~I��uF�$:��+d���V1�-.��z̞�+��B�j���GzQ���{; ��l���FY�Y�f>*�_���E�vy��.:�v��I�Ǉ�a��m(�ge��Y��9�k�c���1��8)���G��������CG��ص��U��>__h"�@�E*�b�����
�1Gt�	�����ـ��W���L8��4�W�5��-1�1L�`�D�x���9�D�MIu!yeM���Ag����Z�Hy��-NJ�Ȃ�Z�W{�/| ��L�u�9N�!��4������Yf��ÑL��yaC{LH�B�;�6��'X��o�0� (��UHzS.�v��aw�,�(�|㨁�I��C7�Yt�()c�Y[��m�@����w-�1S��jzR����0kx$]<k��HpVW���j��P�7�c��Hn,�q���r��á�C.��z�T�VSz�3kr���:�Z���@��O�l��c�mPA	�k�ح�o2�t@�$��T��Ԓ�i"3Z���p��|u�*g&����\{��)�)��Ā�;�[�w�"�~+hnC����ST��o�5+l1D'�-�1#Qbzu��$�.%>��첷ʐzp�]���ˆ�����	8����Lm�5��|GX�._W�oŖ.���#�"g#|9�Ŏ.����H��+0}$�|X��U�V��p}��S�	�D(�Tg��X�_ѵ SL�ܕ�(�K�0#nP�rdr-�W�����XL\�L��v>���rps2�?5�3�0�1��+J���?�K�����P�
�qZy,3�{  &��;g
 Y����k�CqOI�����q�����SϾ���YLskKE�b��U, ��:�x��~*߯�Ga�ˮ�+
�]��E@�~al5k��b|U�W��̵�1�ug�Dn;H��:fj��#rh�y�7�	���b��ߗ��"여��B^�*�_�>6�\M�&���:~��D�r\hí]�4x�����O�G��z{n?͝�T�>�?��L�˕�ǂܲ��5�y����7�p�����$Z�,�Vy#�B��w�e.�����?���>��Q|$�o9�؊�2#���5���=�B�AC��(�uH����C���ge�c"Th	Āz7�.�2>rE��{�j ���y��'`b�=Gힱ��V��!r���nki��)k��?�y(�lI؅������#B������XP:�9K���\])���Lt'���~��w���'2٣b�/���PD�"^Y�x��X(:�4DiD��hh�K���{׎��ID��'Չ�%��T�L��h]�><5A)x	U"�;�5��C :���MC���f��� �;�"�N�=-(Τ��Z#�s~W��:f��C=�U�o������� _q�o�,��V�>/�9E�
"�L�_}��U�DHz=���0��vS/�=��<N9��rV�~u��tI���)đL@��k3Z8	y���&�0�zN�]17Z�,M�{"=>T�r����H.��FtLM�z�r9�{Һn}�k��c#��6F���IC3}x�5��;&��v�(û�:�BL�j���P��Zq��)q�oB����F�X�(D�!4�Υٻϋw&w|�!=� ڽ��rz��JMܛ"�SX���*M->� }�p m��
"IP�>(S8� 
]��3Lw'����XDWV	�d5��A��_���$/�ۍ^([�J�Q}B$��*6PBMw$�c�Vc���[�_9���.����~�;2`F�Y8x�
F���zb�)�8PBd�_����!�uH�{t뽝�t��I�X9o&wHm]cbs�1≈$\�&�	��0��7!qM�h��1�Q�+8H��D�q͢�;l�; U�kS�ϐ�]�@}(�6ж�O��
�Mb��ExS�d|�4��3nb�y�Ófy�|�rd]�P�S�������eD��p�^�l���fpp�ǭ�k� DG���Yt\2��`�d1y4acV�|�?�&�Vm4�)���Ӳ �7����b�Lo�����
'Y_g�a("�l��H�m��O�ˠ��cfk��tw�4,�;^.D�� @���Y�Ԓ: z�������|���S�K{�.�LO����1�O��6��_�_D�R��d�F����؄�k�lEа��ڞ���\R�QdR,�xY�����僫n�����=��"�Ib<>��Q��-�Br����y� /�G��`ݝb�]��G)ߚ��L��Z�?X���1�6����u�o;a )�lo�?�ޓ���S�E�<�h�G�QyV�?�2��\u��H��
�:w�_��$%�d���n{�1�0���p����j��d����Q�;�)j������X����GS�~�߸����y8�ƛ���
ٸ[��׍q�Ja0��3&)��	U���s��u��^��(J'�v�wdi��t)&����ȇ�y��qCG���e�CD�|���i�����4���Z����S���YOkg(�@P��d���Z=�`�Iq煲n�Q����n}}MJ��А�@nx��zY��s�L�V�N8���U��b`C��܌�0�d5�=3;�����=&�A셲Or�Xg�Jw����6���u�����{��V7�@���K�{��[ O�X��C������a���"�]%,׸�r�L�iA��=g���4B�,AW4��Y�44���δ��(s��
�˧�٬){p$��O� ����u�$������
Wо��S�� ��9L#-�`��d�1�
��}I��M��Xo��ț�0�5SAg8-����Qx�	k1�?����F[����C�Y�'ۺ��g�8W���1��6NF�~J}��@�C�K�A����e
�ףA�`Œ��ѝ�)f�)o�Ee�X3����m�%ף!oa#�XYz���|�\b�#����}A�s���KH�/o�鰪�k,�#ӫRL����}õ�d�b����D�!Ek��{�Mٳ��6��|��������9SUGr��<�1�6[Lz�%��2״8�@/��ԅ׭�~3XDYvY�ұ���o���o�;h��HӇ�S��
�[��/��aZ){Gj����髺�\�Sd=K��;y�f�c��959	#_O~��N��}��aB!?N��*v6iݫ����l�hb�1~�N�S�kGn;w�	#���K���^j��r'�"�3��K=�#C4�L��*�m{��4��0l��� ��o/q_��Rިn:	]��e��ޱ5'� �?e֪�:ʗ��j��C�tU%�ql������i�/8�|�[F�H.D��ӵ��kގ���Z�K6RL�|ԺbںP����\�:��<z0��0��g! �R��������h����
�}]�[Y��4��i<�5�H4��A4��O�q��,b�N�@��(!pQ^�>��߻%!;�h��B{%>e�~{Y��X��E�*G}:IP�쯠�8L���5��)��>�)�4|aޮGu�Ks��`���+��m��0+?��#י$�o��p�>�V�r ؟R}�4�� )	-ß�!�-���'6 ��p�pA�1\�bDIDX�|��dJ�2��&����^�^������m�%��:U�\�7��bWre�w?jW�l7,s��Vdd�3,'�C�~/�W��v@��L�:���'�=�+��4U��_#7�W��]4.:��S��%6��'�[����F�Q Gy����l^UL�5[DJI����H+Z��e�
� �Z�}�#d��u���L2����=5#���©w�r�[��|-l}ũ�A��/,~{3���#*A��+Lظ�G1�X�J��iy�)��ŉPz��;M�՛��;��$������j�P��U	"�	���-h ��z3=�W��D:���F���4F�i��ӞD��91�O�
�	�7�������J���*��t�>��Zf��1�i�uAh���w�֦)_�aᘩ��$���i�7U&���l��p:��Ư�J���GDak������L=��_y����⸋5����-���V�x3��7�}�$z�����U��˅�%�9!���S�m�a��˘�[R������B��ˈGW���Fd�<@�)*U}���hʑ�D���g]���y,����8 ��;]�Ы�s���0����{]W����i�4�w�g�N
�܉�+D�&�h)pB�<�)݁*]�2&B���[��������z�;�X�ys��ή���	�����x$�\�^�?d���=#X	���6�����]T���(��������\�1;8�di,r�"��YD+�q�sVJS�!N�ϴ�EA���M���gG� jT˥�(������b�>@"0Ci�:)�u�����F���u�Ōc��vx�$𧂝N��"�!q��r�[%\�ɔ[�t|v�S����·2-&+���oiQZ�3Z�䢄�Ҳ��i0�����t��#����N��p �- Z�\n[ �{�Yu�_����MWduFK�a�-�իI}��4P���^0�?D�I�M)u(��@�"�5�W|B#����)�t*'��>SN�P�C�F ]xǜG��A��1����rDwk�Nkb��iB <��ϫ$!>��9dr0񌔉Di�4���O�wBV%<Q�G(�>⑳/\�I��z��&s\]1��6探/�} ��0\������E��2��w �[8�w����c˩�(������k�f�����}z����(T�ܵN����%�r�����:����
y�\Y昢:˖JY�ʦ	��'Xw�p2�������C�RQ��s��@��S 0�l#���x�q�������?"�J�Ov��Ho����A��-q�3�L1`��~0Q++����G�]6��:f67\�s�P-℃�;����V�	�	��a|x�D] |_�Om��>甾����Z�k?e�"�0vU�����(�RS��Wk�����bu��~�t� z!��u��SX��)�<ǒ�:�֑��8�>4|V!���A�_��1ӟ�j/ O\�Fͬ=եH����!|�$;��33�cp �?U_GDo�m<	n�mA���؂GB�(���س8U���ro�J�]��]�R9�i��# C�素E���ir������睱�:���R]p���q"�m��{�.Ұ#�\�[��t�=[aB�IO8_H༫]7�p5�I/0)�I���.���ξK �Z^�hxL`�v��t��+�Te��[ipb�=��x��T(mq؏aŚ�bm�����2f>�wԵ�[$&�G��AǬXJ9D=q�4����Y�Ѯ�e1�;C�~Z En��=��v{K�M�>v���"�����WBJ�V:�m}� �����$ͧ}H7�#k-���?gY�Me\�q�4�k:��r�+�Me��DH\{��'CL�q�d����r��a��Y��H&���{��Y�h��]�$�ջ{�=�փ������?'|!e9r;`<��y���~�����7��K_fn}�#���dZ�)nAde/a����JA.3�Z����"сOUs_o&���E����<�/��i+��o�0k���Q4��i�&~�����H�_[ �!/j&Yr!3]���.WK�T�dɯ��h�OC8A�$��y�g��^_��`�t�B"T��z��f����r݂���^��ZZ o��H�鮲�:;����^�ޮMu�>��w��w�䌺��)E���Q��N�X�f j��K �&K#-߾�T:i8N�>kZ3������h�գ���A[rZ�����Qn+�ִ�!���%��BZ��@:^�oo�=�{���� l����#����E����isJs�@�2
�0���x���<G#�1�&��zm���b��&�!�D>�|%}]�k��4��b�U+}��$ /RE����E^���J�<Zd��i@�2]a*�M�����RS�s���(���l�Y���4n F�gC5�t���Mo�{mIQ��7hWAWmIqL[GOh0�WNGI4 ��6*6���ÓĬi \������*틣Y�:�eM/(�N`bak��G^{N@T7.�.��dm�H����R��י���"�ȀkJ!d��Y�ҳ�r���r�Ҕ�O��6(���%�@�{@��=�v(�(���t$����� d��d�w����?��zB1j
E`a�Yz;R���E�da�ɡ`�@���[��EL�Z�JY!���\�߄�,[�=�,��t���;�����ѿ����Ԉ���*��U�x�A:|GC���R�����Xa�T^`�Ia����i::�PXd��OF��)���=�/����b^(�Ć��}��
�JK�iD
���lAQP���[�\����^z�J҂�����AN�/�$���ɢ������tϘں��]�H{�*����\��fvڔXT����?x��p�����d+�f�udq0-�(A�r�p����h�����*������'5�>��_=��2�ن�1$s~����{�Ve�&��p{q%��E���LW�_�.]I˰��P>)��S^{S'|�w�+�� m۵��(dAW��.L��D�38:z��VNhml����t�NϽQT�hM�v�b��X&p�E���d^io+�γ3I�a��U��01:r�XIܼ�|�!�/�A�2���	�]���?����
�<��a���J#߸\��Ы*A+�h���kj�X(�����G��N�8�P�ڰ��+�����e���x7���g��n���,�ՠ?��C��Goch����+���מ�hа�^�z�
��qy�yx�'��dq2�lN�E�y�k�>�[�����qb����5����wDZ�XN�>�r�{��.!��fxn�g4���o��ѢS,��O�}+\��b�4��L2��T[�8�@�Ϡm��W]6=l�I��e�b��V�rU�N2E7�
-����9������_=����ʖ�B�T����3�sr� ]';�.Z8���=��0D����
߇E��(Oc�,��]����ժ�	�����4c�8��.��h/�E��D������sFٕp�,��:ݓP��"�uQ>��܉�8�HҴ�'�=1�8)ن��H�K��"�����_�sD|U�	Ld\}?���7�1���Qa�N������f$�*@����3�}M����a�xb��!����s�v����E���0�[ⵖ��~�n�����P�K1��$��,s�6�=P�I�N}�H84d�ʰ�V�f��8l,&�d �_\�k��7�J\4�,u����j�d�y����Q��8$N��T�H >Q�\QՐ0�-N�wvd����t���>�"�l==�M���{���8ٺ�?,jW����qI��?@/�lN�^�^��m��YK�"�2�'}u�d�Y�;c�a^|�8@���kߢ�(g{(�d*
�t���ɌY6�t���W��P�
��YCZٸ�7!��2�v<�9ν���c�D�E��P���C���]7���G��=!��:�P�6����f�+�C�;"�?���~�kV�&��7$m����g��ٽ�M�U'�ei���?2���ٻW!� ��T
����&������˴%7)����ɗ6��Eo�p���-S>���p�~�s���¤\!���-�[ϐ��0��T\�dx~���hr6�k$�ل�r�v��쟿Y>8��g�w���_�r�"=:A(n}]�`؆���Fl�o�fM���	2u����]���b΄���2}�����c�$���M�i�r5��X�2�w�#Q�&��YĢƗmtp�'02�l������m7Γ{3���;I̟>�ץ�~��S�Q��v�����Y�ܽ8�l�x8	Y&5�8� z�ޣ{x�����~��A��/�#@�e�q�,��xJ4~<�O7^AU�@ 4yA�u�/ƍ��ښ:N�4d>�-�ܖ�$o8x�1�K�J�"\6��=Z���T�j�<V�fӰ6���C��1�E���4������g����R�Ĕ��Kh�Jn�w�?B��/�?�0c�JE�L.�cR�\�<w��.��s8����bT��vQ3\{����&���ǌa��m�7�����C�H(i���g3��O�����,j1C�!3�$f��1!nq�T�����k_���
P��.r��L�@�5k���U5�WJ4p���$�}��Oo�Lna��9 ާ:�B���=��-��Qf�)��m�3қd�-Y:��� �D�G�k26����l& _��x��Q�3���8ly4d��������Umg4���C��6���~r������A��2�8�����_�M�z�\���B�����i�L(+���T���!-��?Z�b%�F527%_�)ܽ&j��#Sz�
�Q��$aj�&�34��1;�	��*R�L-�m�ī4���^��v,˥�]��*9�L?�d�C�[���]�`^~(��V;`G[��0�8"跂��w��$C��5��.�S�M�����J��w�e��Y���-~�F E�mq��n�\G�V���Tl7���Vg�0�Ơ�,�_���#n�F�c��+��dz,Ү��:����������v,ʴ������ǯw�w����^tt����)�ק�'kIj$���U�I�s��5��{�6	���^O�	��N���#�v~��d��z+d��b{OC���{����+�Z�`0��p�\W��pd�r[I�54N���֜� �\��zmH	ۑ;��w�J�L�ýu��٢�t[��� n�z��k�L�$9�Av���^�>dOu�5p� Q��B-�0��B�ay]�(�v��"����Sf����6��!����J��%��x�c�d	��Z�|g�3Z�A�݂k�;�A��o�£D9�X<2<A��uber4�eyg���3�$ �"�إd�r�eD�_�Z�FC�~J-��ܿ�����k���պ��k�A�6^�"?����g�I�ĉH�n��[[o�,�=��L�q����c����q^��"���W8ֽ�o�$:a��}��Bu���%e�Dr/����'5ȉy.hM���k>W�s��e����z1�����Mɍo�z(����E�Z�xT
�<�o�M�HC�=fqТ(��xڤA�5Ŝ~�O�"0y�9��5�n�ܭ��4�-�+�%b��� "�.~��� r?��"7]z��4�L�pw��������aÜ�7�	��Ι8�]����r����ꐊ�vh5"I�ѼC0Ty)&Pt��t��S���3���gZ�A�1�ޢ���J��P�@�u��	ϥ�[ȃ�s_��D���0Jd��c����rB��94T�P^�q`3��D�hK7W����_��f�+!g�À����M��y�8D��'g~q^r<�kS��J�4)��
���P�q�Ctl��Rp���|#������I��Āy�\]��]�4�Y'?x���AW��l�Q�5�{�mU+Ǽ������U͙�B��į���KVw
�Yj�����P��ІWv5����0��t�iZ����^D�s]���u��B�+�Z�ݳښ׵��3����;�l$W~�6j���F�o'Mʃ�%Qb��'EFM�9��v8�;�y�h#⡜�%eT�uu�z��'}t򎳕nJ���gMa`��ܯlY��k�'�N\(�M���6%r�����q�XG�������Jg5.iGd��p>f$a����H`�Q�q�]%h��^�`Sޥw�)Ҷ� ]�dk��Y�����μc0S����I�����)%m�!Р���~��U�*��W�U�^KK�k�f�6N�� "g3f�/��H����z�H�%��q䡫Շ���2�g�^̍��bTe���Z��YNޛDkY��� ��]Ö6? ���o*	�����,�M\.9)M�E
C2����*'������0E���?s;Z��,פ�y� dcN.����zg��Ȳ�fX{�E�}����o~���Bg�3B.�G-g'mk�Jo��J~���P��b�@/	G��������v6r�zq�a�f��5>�>E��Lh�(k�A�5�E�z���i��K���/@��� ���"�5�(�.O/��MU�LP4�P��5ǒb2]X���58�-�(�����XKcO��F�0�3�b1��,^��N��=���˦��N��"=�>��,aàT���9D�8�'������HǊ�C%�4]l!��g��t��.�4�5�b�W^j?P\D�����!���F�L ��C�>;K���2�qk$\���`m�u
�4��8Ed&����K6JM�}�ߩ����@@�`o�������s~=�v@'�h׶,�6��Q�O�`�i{�-��'Rvi��w �����u�-�D�����rIdK�_�=��d�yW���Y!����=d火�� &�p��UW"�D���z��_��Q�F��
k��?�C�zw�]���"vH����|(j����u��e�����~)�����%���[�>��#q�_xC�q<�[̳	�� U��_"9P|�N��X�i���/�%�W�\mC,g��M�`p
����n��Y�,\� ���貦�4�]�����jn��X�U�$(	2Rǂ�/p8����Y���l�VsJުJ��I��:��v�����^3�nژ���tA�I9��\���e�����,8�pG�oI��Z#�ݒ���3ms}�N׸s=��퐥�� �c/���P$�ѧ<��C���*̝���ߌ+x�N�Jg
�Tl������Gꂟ�=���k��0��<���wCG��-��Ǡԙu���:QN��cլ��D{�Y�����Ĩ�f���CM�"A�0t'F�(}�2� ڕ���o�+�t�_���k^���zR����î�0�Z�ɪ���V�  e���HV�I`ބ9��ɮ�ZJ�@���so�$�ޗ쪍M/;���Y�F��^҃<���S�9;9ѽI-������t���g��c	T(�e���JO�xFF���m��JK��K>�!����v� c��
�Ѧ6�9K�$c�}�(�5��Y�P���O�],j���H+�Z�GK����b� �^��{-T.��Jvn���Q���=?��^���b!$�Kg^�qy��M��4��{�$Ǡ�Rl���=s��3�{��@����Ex�8E*g��n���u�bS��9X�wW�+ ���@�2+b��������v��"�Z������CLw�O�e���BV�����������l�9���s/n��/���]b%$A_X"��qH�4�2�����,>���ad(}c��Ɲ�� |[ܙMSz�`�}�%p�r?N��@.����#�CyPV�!����.�D@��oq@d��#�a,:K�ޗk[�OLD�uuN���D0�S��`�(l���Y0"�b���9�������M��쏆��=�t��"�p����#,�j��I��j�a/&��)���g��*]� 4������j
�@s[�����Ep;��B3Ëւ� �ٰ�eɣ��mI���R�F"w(�6n���lCݶ׵ߣ�=f��C�0{%_�i�&�wA�2��`�_su���R�[���A$����	�gy��8�,��'��[M����RW�cR1�HYnk*�J�}�a��]�b�1�gI��e��}�[������}Jѹ���!Cp��$=�_@����
�Xn�*D"+��IF���٠��Q�h�&T�L֜[X��b�~:��bOrÔ=���Y��dn����N<׏�M��`*�^���J"!��GW��Q 1���~΅�=���������o�3�kE�˺>�R.��b��� U&fST�x|��ȟ6{�J��ܛ[S���uP�4��g�os����Wi`h�p	�s ���Ae)�k���}Fe��%@5��Z�ί���h�5վ`����f���W��'2��W�fpȣ2�C�T^���\�Į��.�Ȑ�~S��C��O���]��k+<~����(� �4cy-7+��M�P׹a���F���	��eɸ�ݗ��A�D���� �3l:)r�7�lb\&7抐��r�ʼ>A���R���i��F%.y+ ���T�idX�!���=e�1G˾�tY#���4#q�/��3!�8�Mժ�e���fUɧ�B��{Ҵ����^�����[�m�U�`��Ml/�}�w�g@.5���#,�
�?��kF��u���x�Y�=jN�*��%�����;�M���s���S�
»������d2��L����LP��鶟�$�~����$ٷ�0�Ћ��e�sU�`�<��q�,��2�3K��/s"@��SΟh{����ed���2| �'�fи��>����I��)�ۜ��>�`|��P5�ej~O�r�8J�b��m�l$?��8���}��ֿ%hDƪ����h>a��;������2j�!����si��-�6� k>�U�Y�?���"T�{K�?��t
�=��e�*��
�;��M|D��� ����'��Cޢҍ8�E�}(cq`@ό���B0b���O�	��7�wѵ�m��(z	]t�Z���~��[G�e6�Q��#��[���^�D(�~�͖�/`H]�]�[A|�c�0"+&�UԄ�^�bG-F���7����1�e����2�;c�z<���틍cT��W��x�V&8�"�.���.�#6#��2�4<�C���O��xڌ���]�$E'Ϊ9��S�q��M��k��xeʜ�'~�#��?�Sg��	�n7�K�dFR�3�́?O�cAvmI���W���ZI�l�?㴚3�hcCF�1�R���_y>赎X���A�hv�6+�_�Q���:O�1��_�_�x  ��6��}^����@�-�r���4ɰ�[���/���Ra��T��<�9HM ��z�"0 �+�_m�>VPB���@iK�%�����f��X�Ϸ�b+�G�U���%�֞�O͑QL�"$X�Wm��f,U���o�AD<mJ��Q�k�F!b��B�!��hg	�i��L���U�5{.�	K���e�{6�$	>�mH,ľ	��/�>�"J����K'�|wN��,P�:�g���wC%H~�0����˂��dl̘�*i�9���4ϴ��F���W�X]gb�ز��L��W�G��X���$%6����c�4�ݥ7�2�F5t�=W���ζ����k	fL �&V�ԥLgl��kU[�yyW����*���G��?�C��h�+y"ltd���o�@](��4����[R�����F�Btd/#���"g%����-�Z���@��hm���0����Tݺ�h�㬦v2��!B�S������hY�t[?yNyؗ��M��EJt�D�������M���%Z��a L\n�F���\Xݬ���@��9����Z�gc��|�Ŵ�����]J���Kp�3`pX��];��`7]��-�]���?���Y!�~��W�.1͵���5���U@�L2��3�-h-p�2�^J�R R����3n'���iD�_7�`Td=�mL�p��\���"��������e�O���)ܡJ5H.?t�(y]o��Jp�z��]���`8�աP;A���vd{�gLM����@|@Y�>��4S��ځ�V����{+��?��6��T�j��@>�w�;A��
�g����
����?�0��.Ke?#�VM3�����,�W�eV�u��6�B���Ս����}�l�}��X��x���>���05J<.�nm��<Ӭ`�R�9��U��("q{��{��%e���Jp�Ƕ�I"���갹s��
�!ꔊ��0�FEz�^q�����a|�z�D@G�C8FQ�=5tkti�h�e�/O��ZAH�Z	ƀ!*!H����({��.[���!�h E"��Uε��¯�U�G;�����5��$����+k�9K�����;� |raG�?uf�c"K�X����y�,W���� ��'�E g�M��:��3��k�B��%����:��
|���DbDa��&+]�O,!w���1���FZ�"9�z�^�)��(b�����X�흼=��x՜��1U�>�Js���������D���u�냌����V�`�I���=h�O^�&I��W�����	�朕)|r�;9�l�c�� iސ��w�td�:���<��P�%�yE����"����������29�Z���հ,[�i� QD��kgg����2E�3�gI0��r�9{�k�M�.�:Gc`��s�I��-}�A� ��Qe�������]�יk���(�E�l7��Pw�V�q��/V�F��1��VB�	�f8nQiE�>�O1,��.�˒��<$\c�O���v���N�ǌ�ۊ��_�<F���N�+j�Pa���y��l�Ģ�J��r��������=x ��������%�م��ʓ�KP@{7j(�j�ht�K��$��B
�s���~wcVx:c��2~�<'����:P���9I�����F%,d&De����~(��w���c=�E/brs�5�y.A�]p�N10�&.�̄V��Г�K�\&��K�'�)��X-�&욕�p)22ָ����oR�����?jȾ����Wp��x-a�*]������L�p����މ����f�	���)^������{���V���s�;D�PEv�)����O?Y�u ��yA�m:��{��k��^�|+��-T%2r�j�ѯ����M��ωxsgş}�l��RV��w����"�e�a���_��^4��OJ�h	zl�cK9��*ނ��׏����#��4"A�s��Ǉ>�����Ռ�w�����ǘ RoQ�D{�L��Gs�����S����Q�G&�v��ꇲ�%".��a�1��0_@��)�l�ʋ�cq��fC'@����p>����+l)@f����t&�*dU'������z�M8���Z�yC;u9��j,��T��Q?x3�v�'�� "`>�v2Xi�>968{HR���7�.\����*J5���LF3���0���X�SZ�MD	槿�w�J�2B� 1�{�p5:K烹O�wZ&�'�N&}V�rۡ ��E2��rJ&���n�0Js�b�T+ӄ���6��[��z�SNg5O�ޭm�Ϥ_6Z���k3	'9�:�U ���|R����m�n(2ڌ�!j�`3a]Ptn��lV����"�8I�ƫ�1h�
�i?���2hm�A��А�Ƭ;�K�u�=L��L�Jq�t��g@W:�>����_��!ig܄Y�c=,:������R�e�ǫg�J;���[E�At�˃P�����O ���?�=��G�D����aB�-�Y*xԷ��꩎�+�AW�+-�� >c�#;f���M���p�+ja�>��<));Y�&@v�A�sa�O�O̞Ի ��0<F��4/�= 8%��s�t�!��z��z	Ժ��Y�8y����E����~(��F�,F���L,�[�q�v^U��]7$^����'��5H8���$|`$�][�zaD�'����c�Mz�N����d�'7)��[���6B��>�D��\vrh�v�;�Q�������u0Ǡj���9$��#��$�8Y�I�x�=��&��Q �?���)����	�GοW�ɔW��*X�F��G����dC�u�*S��>�r8���/�J��'i��<�/ij���t����V���9����3�W��8��w��۾�њ@���TI��++�ȟ]q��������<�Q�����2��<X02�!��TO9�1����V� ʻ [5��zq yn��KgO��K3��8��o���o�¸�~Bey�2�kRg��?۲
�9ߞ�+�uz ����7U��D�,�+��jv��Ɏ_7SM�c�u���k?Q0FQ�������8�)�m�q�h��,s��l���k�%횉'�ejS1�ų]�/�_���u�m�h8uX<*��i���"h�v�� eEgUh�zVN�=7�C�]FU� ^��ct�>Rn�Dd(7
�.�O�{Q����ȘW�&�� ~n��ϸdJʃ*��&�O�h�����Q2���l��L�;����5�=�nD����s��y
��;�OZd&7�$���m�I����P��K�zT�5a3�.���_�W<���<����4���egR�	�|Ͷ����̕LIV�IB{K�F�x��s����ФeBAH �&�΁ҩo@���6�e�H���B����F}��^�ݘ��t�~5ȯ��-�����z��ͨ|^�2����6c�m���ݕ��e�k�
Y$��]�u����Ok����[/E�avS�o���qm���\Cǉ6h�������Hӫ��枖/`�>�OB�O%�v�M�������������8m��������MY�ɔ������H���"��0S��x������a�����W`����/U�~l2�����_�RDGZ��7��N_��\cz:\�4��b����r;��Kz ��L1�Lm���?Xf��H������]�X:5�5� ��i��O��b����:��i'���3t$�6�����|�L�`�	�Ta�Vx*�;��6q\-n�m���y,��$`��<zE4���m)�s��Dkf�mqt.�5)*��A<;�	����!G���	����cʱ
CG+��EMj��RHortYC�R�i�76��K��<�wN��B�1��Ɖ@a9r��V/���6�	co!�@w��b��{�%������$�H���:���>�w�*��39�M�8M
�䡂�樀	��M1!`���씒8�ny���-?�G�*W�`�������aqܽ�kÉ�0��!|�#V<ݙ:�YH$I\�q�X�kpM��b~�·TLD�o�"��	��$y��U�U�%ᢗ����BJ��\���q�L�د(�~��-nk�8���Ur>�!��YX7	˩+�X`
�K�΋Hwd��i��o��Ѽ�:���)�AI��uN�D������2�g�šbЌRq��P�/���Z[Z�G��66߬�}Ƽ���Ѯ�K�8Y������^Վ!�A!����(�~�84�X�.c;�j�s�=6~Sޠ9���ES��ش��V{�����I��!�L�|�<Z�]�n���CL�]�$Q��z(JnW��P�!G�9Ek�\L��E\d����9�.%�Z��l�He�q�8���@C5����Y>���,t#�V���E(��Y{l��ú#0`�?��A���z3���ߊ�o�����vFe�6?�Iz�"��Nv���U �.;����'�Q�'��0���lLz�,ϔT�'?�'������
����3�8i��?5���V�}��}Vd�z'��w]7�:v��]�za�q]��r����eB�I	�G״�����0���j+�5��m�xDT�f@oƙ�rsdl�m��w\0[�M1����ME�6Ln0S�Cz�3ip~%Sh�^����Q�ja�<��{��HF=e���4Bw\��h�.3 g��=�-�7��G�Σ	�t��}J�g������P���A�u�����#	y�s�%��=�.��衏�Ժ�a�W�6���>n*k����
4���u�|����H�����o�mL�w��F*�|�Q�<�-�[ ��+��%��u�K�M˕��`Z����,���zS*⛮������T	}-�0Z�x3l����7��fϓ�?2��X�o,Tp]�Z`Wdփ��ӹ�b@-��J^��Ku��~~�)�/�t 9+�gǆ["j����@~.�p�~���I�D����G��bJ����P0v�w����:e�t�e򣺵USO��8o��5:�T���4�3��dNl��U�Go��TV��H�ӊ"��*�����}Ѡo��_53,�X߄BH� t���l�Zǰl�]!�Q���y�b:�>2�#�t�3��g76�P���4�QĠ"G��( ����ٚ-A�`6e%C#7O�������O�+f��S���*&���L~r��m>��R3��� -��;�Y�pb��O>bU!� n�CS�B���n9GNw�4�x���ݧ�ɏw�<�qu�e������w�/l����8���!2�zq��h��g�L�Kd=j�[��4�H�=�8Ƚ�tIz��"�T�xmE������.g)O�^�U��I1A����������q6 ��	YXƜ�����&	���׶d\wlź.iB>vœ��o~j��8�3�&�K~Ưı�vGZy?�Q��Z��a��a���Ke
�F���T��̻u�5(�}47tn�u�D�Bk��;��ҥ�����B(����9����%�E��e�^=4��+ � Np��ŀ��&��n{?ȀJ�)�X��ċ�BJ�S�\q�¯�.m���������_c��ÿ�.�6M V#g)͕�ȳaO��}[I��Af��Hҫ��Z?�����ڎ[�Y��fi^Y��:*�{C�����Y���#觿��Qє�3�ͤ���-P �ОLн� @�ج0P����(�����i2�3S��7��(�'�U�a2�r!{u��h�%s��R��1)�6=���})#�E
�I)��&0��a�8�}����Ja�CP8���Hڰ����k�}[<�= �þ6��T2R���>���&d�ƨ�crDo:���SL6'evl�]�ʗqpq��*�gj��@~Z"oD����^�J-Q�y����q��W9e;19i�gF[0r.G��ؽf?�n���#�g��_��"k�l%���L|ЀA�8�<��I�q��b�-1)�.����|���`H�4��,�b��˿[�4���UW�tnւzC��Əe�oz�1���Φ5n����ps�@�7,��:�+7����m>�q���MҞQ"s�@e6�]H�Ẩ���������']2 $���ȵc�����N$�H�췯��}n��@��0�S���8��B�@��V&Zѵ���қj�
�J���[�I�nK�el���HЃΊ�V��[+�TS]G���F�9���h����)09�NN 
s/Ng�!&�`��X�!���]�j�FJ|13��S��3t�������ߣ�'��������x�%
���/��k0�3��`ȝȨ��.M�r5���3lu�5(�?\�ݒ�!yw�K?t�'��)2�jPym�rِ0���cg�>r��h=��kDf^�BBW4%(�O��h7]D���a���Y�U%�ʃ��P�P��)G;VAi��	�~�"ixL�qѽEQ`<��p��3��^~d��z�U�TJ�7�4��C�C�a����C�,+�^:����ol{x'c���#�V�5��������C�%����_9����\Ⱥ�x�>PL�����^E��W�m/w���zK]p�*א��it�ȲNb�-O��v�Q�!�WX�P�o� c��u}���'N������>�r�}�n�@�a���W�r5�u�o��S��O9�p�\���U�]X�M!F�%X�"����nm
|��jw_���?qeP�����|;��O<��a�lױ�(����z�<8�`s����`�>Lf#���F�$��^蟮�>����X�l�+`�a(&H�ڦ3#��Fa�4Ϧ�l������������T��+�j���)k���@9�{j��?�h�����n`�tp�2IQ*M�Q����`�������X��`�0 �ؓ�N��leh0���JvG`�T�����!`�f��)���^��o@�N��"䔿�EG����k���xT ����]b����p7�`b{��� �:�"���p*l���*�tS½�k%p�Г���d.�,���;n/����Q�O�_�o8ac�哝z�1�2���=�}zz�|,TŃ*�Y�l��P���Jl��<�D�9Jq�B%0���r�G	���3�S�#��KDn9�>R�.G�u��rqV�po��-� WB���X��^V�h����y����q#��!���ɲOUWZoE��JOi�j�5��#��Y27ϰ|r���\"�N�&��L�z�	��H
	��S~-K	��2=Fh,�u@�`K�~jH�K�\M6K��_�C���#��tDd0��q�q�g�^�2-50^U�`uZy]+��𳢨:��Ku�usPo�2��)����*�ɿ���lR���)��j�{'�5�ǌ��k�;�x�ai�Fi�`�1:�q?'Än'�����hS�X~�C��c�|^Y0��}+�a�A6����,�D3{�B��"�6���ؖE��hr6y��"K���m+���(���k0Hu5���6�M�O9��ޥ�=ǂ� gGt��趈�`��J�Z��bE����`������'�x��E�!�倇���䑀K�J�y��������O���:�����������̿��3��l�Wk!u��G&�8��|���)�^������Q �
8:��QA��!�~_��`
��!���5�X-{!2gW0b�w�Ff�������C�gQ�C�6���,��Ʀ�֡��%q�rꄠ�$�A��^�B�Q�Yc�����ԓ�4K�8��?���Y?��0e��R��'��s�Am�L쵗>޻=��O�.l�Һ��~��D�)�5\&���18��3w#�[hi�/T�,~�D���C�ʵ\�2�XQDx�V�S|u�Ts�|�n�9n�԰���E<�<�$�����)G%�B>�]�QҊ�G��� �N��oG2x��/刎ǫ�(����1;(H�z�����|�� HN�
����`z���eG�/�aL��u�|=1�jS��ǋ�)�v�f8I�$��	����)�9��\���Mg����NK��a3��� �Z�Y!hk�pAy%ު�7���[�y	]a�6z�&�LLV	�9���S_��f���>�.�r�O�~`�]
�%zr(��X:[�$M��w$�� M��x"�KR�D5�.����ɞi ;t^*� o[f�� ����t�c�粏� �%us�|(R�S�x� ���-��k�����Ѷ�&<:�� *�A��7��Nl���G�Z��'�o���>c�_�v�R$���}�t?S6!mg��DQ���϶<��ۈ�kǮ�1[�����E��}�_?�B-��$�{�4�-�c���,�s�
�$�=�W���}�M�B����"*�e/լw�]�de�iuE�_gAU����#l�>n�6��kp�0��&��U	��U��&�7O�_��{���g���&U2����Ӭ��Iz�b7q^k>�g���t����0�G������2����h<�+��/�%&�a�0z����8tVt)�?�0U����~��<���Y�P�%~�B���N��a�D��7֢��#���e�D���y�����K�@e�ʄٷ�����������џ�:�~�Ҿƹ�gZ�	a/������4�o���_��ǵ#�זm��O�[�S�g����3i]�ɇ��5�Zj�{�vZ\P> �j�u�˦�|�1�>��+a!�Nղ�9j�@���cz��~��H7�.�(�1�/���N��*�p���ѩѕ�yD�?F'��`�ț2�w)n��ʿt�=���-��i3�Pn��^�ߘWJ	��8��:�|�t��V���_־~O5��&�u�|��v{���z���	`�7�s��H ����%u,\?A�z����Ή��J:?�Χ�~����Z���U��
9|�v�v�gA�`n��޸'
�'4:��Bx��U@���h�������2���b3E�%OFBS��;pu��\� 7n�P�J�����%~�7��+�t��<��9�튊E�����/rH�����k�?�|O���JS֐�D&�Blni3�i�c�M������3>\�m�K�)�n߬M�ǈ�(11��D  �FA��
�Q����'�d�����05v�}���m�Li�1R�i��dyt�c�T�䄳6t��ɼJ�'@ �Ш�Q%������>�g���4,��1�o(ii^(����u(�bq˖��Bh��TysB氦ZF�݁`9��7��M�i:s|�u7����,~�P!��1�w
��PȦ��R��& N�T
y��׌�GW>�
o�^U�k8�l��+X�;!+�h�'�r;3�X��뽫�q��v>KFc[:�OJ�?WG8ɗ��芣�2�*��VK�?�Ue�3޹�:��v|Khp��O�*�7���jReV-���MF���-�s�N�)v;�*Ն�e���P��t� h�^)�d��������^o5r�j@4�͛NS��J�u�/��-U|"�H�|�2��C#s��x��%C/�����U�T@p8�%�j}h�0G����|��q;���#"@�L. ���!�	
8�U*���uL~�-5�~�GH`���R·�����/C�ց�������ը�������Q�F$6��_���ڍ�ԛ7n�Q��@�8�X��+�c�U�Q��'���3�/f�;;�+{j�а�r/7xP�Q�A�c�Ab!��IN5����&Rb�8q�E5�� b���^au�LY�'����tl���|T��%���6�����we�@z���T���FȀ��^o���<Bs�'�C�,�DU��U�|�S�����
\B���;��+B���L(i�c����un �&���^�s����
�kLn��4ەM�Mi	���$�����4�$?�Ge�DXC��W	Xx�7�cȲ�q�N�k�56mII�����8l��7\����{�v�T$�P}��b+��d�l֋c�E��[h��~X���r0QqXB/��婷ol�ǲ1�ee;�v��3N��:2�0�M}T����<k4�˥�&����胪��0��C'�RSD��>J݌S�6�l��G	}���;�I�iW�a[���^�@ݿ09z�� 4Y���j��A�ǟA|F�a2��i}�Pw��%j����_�Z�����hn�E�y�8�2o�޿�I37���	�%�V,�)�l��pc��ނMh�-^<�TJ/�b��\ Xnb�ѯd��)c�&M�Ʒ�3��g�
�at6�&��<ٸ��ޤ;1�&(�%�����uEd�d���z�U���<�F���.5Ƙ���bjFl��X���@\���]�*T9@������&�S��i�c�	Bf�lHq���o�c��zѿqb��3X��	�J"7�[=�����יけ��!��C�6#���M>�
�0er���� �.�H�3���ir���o�S�a(�?�k���,�AE�
d��|ɛ���\'��@��1�Là�7�L�96�þMsВ7p9X	!���?߲�ui�����v�(o��8JW�j+��b���^���:0!/��W��}ɔ3���+s&����F�I
R�����6�'�-�M���:����0�.1���Ҕ�O�{P���L�e��T�Sk\�@�7 ��É� d�(e�v��0�z@��`L]ȄK[�>��{kn�N���=��(���>B �Y�߽��#ɎK�A�bqu�Wga��8F
�^*�5�n##5Z8�?4��wyh6=�᱉�Tq�,I2�Syi�L AH~f�ߌ[AQD��E�/;8� �H��6\�^",u��LW1O��T��V��I����C�
J���-*.�*J/Z �`;���6��NK�����ޔ0o�D@5Z���X��+��E��;f�O���S�˿���#xD�tsd�r�R��U;:3D"�̟�|4E�-����Vz�&Ͻ>�ˋ�xB��.��1*��߲G�T�WH��A�}ޙ�5�?-�μ�Q�ݬ#��z=��<d`Ƕŝ������i�����pO��t����i:Ҭd��&П��#�{��Y״�5�Nϋ����^��'�ʙ��n�9�2����oL��_�8����M�D�v%���_`P�f�`��ǳ�4b��Kr�n~$��:Q���{�*{O��.#,ګ�-�7_P{�JޮNu��@iƠ�rC�˞Z���ȇ�{�ߋw!Z��S�r��Ս�9�{�2*799Y�x�g�_.%��;p``�RB�p�(ɾ�:-'��}�Ms$���YmaH<˕�z�L��Y�/��-I�ࢀ�#g��_j2��ti��X����&���a	��W�MR�k�J�|$��+�U�.�Ki�� (-(/��մCC�����K�Z
���t�=�;2[��x�l4�.�O�_eQ��M��g]��WX���Z<.G��B%�rTI��n�J^<�zd��q�{�<�I���[!c�QHGn���[6��Cı}#uwO$Q3.{�#�L�a��A�F�z�������ٸ���F3/*�=������1?�-�-���rN�%��<����s%C�n��T�j͚m�%��8}4:�����Y��`h��urB���Q��`���#�O�{Q�kDY��F�:����-���u�����m�+��{��p��,�MݷG.� �QA�}�2��`ySC�7FĮ�8��Κ^W6�H���d��x{k��P��p«N,�kU�?�7T6G5��S{P�'�� �]�r�a���??�d*1�2xl��I����#�4�X��qYsIA��{-o_=��b���!*a��W�O}.�8 ��a�.$t��c��
[s+��/J�����̮ߵ��z�!c`4�C�S|
�����m�B�!͈Ɵ;����
[#m�&r�܀i�x��K���@Ϭ�� �%����Z��aSЙ�]�_�|f	����N��k,0#�b���N5CP�)"C�ߊ�")�71�:2@�J��U�_p`��	�����#\=��:��>�L5���g�t��2y��1^�MJ��>�:.X:%�_���*qy6��q�b��(��j\�}{�*��`���Dm�3�v��?�p��$���\Dɱ�K3�J�G�o�C��� W28���Dc�+�u�DS{{QV��rXf2�಑��ϥ��tw�ϋ��`8't�C���4x����t�H��_��݅�?~_}�7_�����E���e��W��y�i�2���sL0������\�T0]��G���3�U�А�9'�?��h���K����0�p(����$8��!Hd�����+�- cc�3>���7���	Z'WȐ�p��ֽtm���p�J���A)�p͟w)�Q4��W
~���,T[����OW�|�=�p:��]��4UFS���s�!`{��n%�_`��\��������OPY/L�mMx��G�/�q��Z���&>:��>A�Θ`��qje���y`��o�n��6TC�t����R����W�[k ��#&V��o���� l�8=��a�����
�.׼x�8a�M5J��VBM�C�WT�[;̠�I�/$@���K$x��"��c�|8��[��Bt��0]U+�f-J��+aE�`�H�H �?�p�����mI40V%��
��c�Ϩgx
������\�!�ϰ����4�m�5N=�7�y��	��I)U��$�1�,��R�=��_A�>�����xS���x^�8�Y�q'��^o�w�A&����x�t�.z����+s����23��9F��,Oj[�׼e��O�t$Y�3��Pa��#�/Gl�u2�H7V'] ���#�w6�"|�P�i�EӋP�؝����1��*wNx:�)��ɱ���@�I�k��d����3V=:{���O`����Im�Q��©��Y��D�� �6�D�����G�J׸B��=;~��r	?� �6U8��o$E��(ڱv�#�i}�425��#��T.�������M͵F�����8q��Z�u�V�W�i|�,���`�(T�COҪW{�g�Ss_b�b���P�J,�Mr��%8m���z���X��ٵ���լ0��v0mץvo}&�ǜw����|D�k�h���`�y���n�{^�:��}�R˺���&e�ɍj|��#�Iح�Drxd)�RO6���q�����xԻ�Q~X��-C�xwqP����^z�#q�e	�5��u���{R�&�%_���h�����*`�է^yn�@�>Su)X���y�u	�I��_BLC.��	�П�Ӭ��fp�%�|���C�kb%�e�区�K�\��6[�B�N���w�����"���uZ�9��L��o��X� =������pkJ�9�ӕ���U�#�'�� ����k�!/N/CI��Ҍ��L�F�2��z�ḶO���d����i��Lz��sS�}'��^�s�h�Ֆ��v,N�G1�����1���R�*(9�9 �̖���%�_`(����$���х�(l�5K���I������|��(=#niv�@D���8<��azb� >�h�0�w��5J��)�:��n1����u�V6�����˭q��qΩ�#5�"�\p�
:y�������/v���E������-�ԋ�7�+��,رՑ�
�?�96jeJ�_4��fke�6pV��^�9Ͽ���O/�
�C���퟇�L�W=�3MFX����q!�2�'�m�ᛶ{;ip͙X�B'u�Nt9s��@z�CO�d'��j/���h{��ׂyf����٬���*� ���bE[�h=��U�d�>���� ��2і�19:R��w����д�)���v�N�X�Qd�.�sI0-i·�D\&�?�.���C���x�����?�*+�nae�3ȁA��W!|�H{;�*��� �ɚ��w�ͅޢ��w��<�>������8VNX�Xލ��Zpّ��p}g�s%��2����y&�yG���T��Е�<Jb-Y�b�/CF���m��v3cJ��D*;��	��t=&�K��k�X�Z���L;b(���Q`�c�X<��p!-`���숉ϻˡ��sp���(�^�5lS��ϖ[|˦�,HH`��Pe�n80�����l�����ǷS�.�(d�b?�u%o�kJ'�)a���{vax��OK��(77ɡ0��k�"�<�)iK~��U�oO�s����\��L���@U�dTz�VK�6����3��2�?8�-s��MpM�R޿��Y�&��>T�Z�T��e��~w�����7zƃj6�7W|�m���P+/����Y��R��0���8e#?C�[����u��= :�p!��dm�!���rP{���Ln�6L�����[�Bp�AB��tL뉗�c6)��*~�2.�7%Jǔ�C����wlH��ՠ�GB�	7���b	d앦pQ�s�=�O h�)2ݽ��i�5ώ�q��>�܀�LvRM���#�
xI)���I��a�[hGN�cͬ���/�M}��r%��������˫�Q���O�Ls"�q�6�,(re�Y� �x�(�&+3��=y��7v�����op��&��g�g��4���U��D�߷�h~D׍o���9�=�����ԛ��e��2�Xs�5��V��h���
0]���'vxV���p&C	�\�qS�g���og�����WAϣ�����J���� �B��w������^iꛔm���7��=����YHM��1gъ׶k`�@m7f�ou�������������Ƌv��X�v�.	�2�y��9�0ƹJ�$�7xrq���/e�w�#�vm��1���"���I�:����&�a���|u;L\٬T �uG3��9�jzp��:�*���/�0��F�k��r�A{{�a�Aj�φ�H�a�#�>bi�赀%1�jw�3�j����<����\�	�ۼ�yC��u��2�`	ꏗ��ch۽wÍe���P��k��	�v�+��	cы�NT���;�,�3E��T�R�Ǒ�2���V�6Y��47�(�j=��_��/��"a���+��U��F�Z�Q�%��J��"�ܡ0��� >:"Ű��Fߐ�q���.o&���O��H�)��\;���0ʡu��-��D��?�Y����@
m�:�NԐ$
���o�ڷ(��"�	��e#�	��7m��N������p傛�Y����gV�0Ss�L�{�}O�.�'�Kk�$���ئ�@�;���I��*`vS���ۼ}��z%��(��ǣ��uS�ej�d\.���h�0I�E��
��,��g�G� �v�|��Re�:����s���@\\N�������m ��X��ɹ��N���T�V�:x��9R�nX�m�����@|��	(y��C�&��Go���SMW�����r�~��gm��#A�`���Jb��g����W�cO_׊��|�L�{��C�!��G�U0� �:�E�d
<Cc>��<s�s4���9��pXq��Dn�8~W�HB�о���y�L.�TH���L5��S=�1j��g��ֺ��s�������b����]!A�f۵�]7�:I�i���?�v���Xq����7Gk4�"�{���Yk�P�0͋6�>+����}�k="��3�vo�7�6���	"��C1�:�i]x���?���5�)RG�	Ô;�M�ɻQ�Y�D�)�W�A{0��)c7zc0馮����#��s���=�%���|h����|j�:�5͚ײJˤ�d�b�c�*�a�;�N����O��s�1�qrc��P�S;$�h,��x�iːU�k@�'CG98�?�̵>Ç�asS8�~�{����!