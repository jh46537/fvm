��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*�ũR��KE��1Г��,���'ˏN�q,�9��V�D��˙��{���!��Y���I�9=������N��U�GuW��p<�����"/���#���1��d��m��isp�uU#`T�ȗ\�q$Z��وڬ�R���і����A���j`ҙ��X��@@��0�ļ�5u��~�W0������tx���_���&�ѰZv4wE���?ѩ�;L���$	0���~���U�b����@��R�ʵklha�c&���f��<j����!��<&�FQ� :/���F<�O�M�C]�e.��s�pÕ*6��ɾ+�6O�J�\�E��L�,���$~�I�D��Ƶ v,@�5/�`,c���LSE���3� n��"T������U�H���t`�����C���woo�x��� /�W�Z��݇B�`$R]Ȟ�I�ctsns|�<�-ej/ԔN&"�QM%m�du��4��<iB����4��Q����q�plar_'��桲��\Jw-�>v1`Wĸ���� :ꝺKOy5����iFR��3�Xag��I>�Uxf���'*�*�-����v�(���E������D�Lj����b�+�|Q�͵uY�r���f�߫�Ɗ�}���(??A��}��曗��2�:��W���F�u��0&�U���`)�}4��gr���F������J�O<��L"R5�hŉ��V�p༦��OHQ����
[��'櫁���G&uw/DKM��5�P�ѢX��ާ��0-���Q�b��ݳ$�F��D��^G�޹d6�ז�ᒕ=��n�e�Yj���)��#���++�]' Ԅi��bo���*�xuO���m�S X�<�%�Ln�������y>�!y
V��7gz�y�u����� j�m@T3�������c]"KؘXo��2�~�˽�,CB~��F�N/�Jm)b-~=����A�U)�75�A���t�{�Jd�R��] ��
WȀ8�����G}����_"�\D����B|dyt����l��S?fM`uWt6J�XC��~�bM��JR+D���ջm/�IY����0�o� ��v)4��vNe�;����z����,9�*$"k�/?����҈zNqp��9'ݣ<����a��rPVZ�8�qy��MZV����m�@�		>����kk5	�Ϛ�X87<�fg�R�Ə��,�a�n�֭tIw����c:v[�<�l��d54f��۴O�T�8���p��j�n���I�@���"�ɂ��H�3]�s�v�Q�븨�[�i��͇.,>��3���� �������:R��Ơݓ��w���l���#tE[��r�X25$�Ta)U!�ႬVǬ�=�.&ꮱ���{������-�%��z�� ���?`ew�*�H�F��i�
���u#��a�� �CYͩO�w��#�)�;��Y��V(���Zm�짋�ӻ3�[�:��Ȫ�{�c=�_��47�{����?@Cn?�Ñi� Ћ�A��v��F�0��h�9���ٷٚv@�,^�0
jb�Dej{�J�}̯���F[p���d߆\��|�ՌI"]��i�ډ.h�n�����0����X��+a|(VU��C;����<�B[�o���(�$[y6R|��e9���x઼����vy����Ļ�H��`�S�������Wg������M���X�\x�R�}%�<���~�u��;�h��$t,)�>W�$�,{Ö7i�h�yLGؕ�<�o+jL�˃�+���.mXU�r�P5�7�,���J*���'�C�}`ץ<�o21�Z�H#:��j$�)��6��*Tc7��a��E'W�A5�uV���w/���I<�İ!����y_D�y]��s~>���Aw�ds{Pg��$@�LB�@Gwl�.�a��p�,A8�Q��Q��ɖ��$	��(�;��Wo�J���֙A�1A:c�N�vg��6��)C6gQ��j�}\�Qh��7?�5�c�YQ��W��@��⋱���R����g)ν@�3]����V	Y.[%2]b׬��i��
j
#H4��9θ_J�¬��4�	f+�z;������0��0P�I1�m[sL�2�I��jnL�Q/:6ZϪ.�_��4k�$5���Qr�䅋��r�!jh����
Fd�p���*��1#K��O�r\[\���e�iG|/iE�EH�J�	Uh�� }��Z�>	���
�+�H�-�?��M�wL�_��a�t/������j�qR�O1��p�|I'�K��TM2-��p�0�5���>Bu����!E�
>I���I ]��;l�-4gM\?�̀��ٍV��A�XR� �t
�Y.Z�����v�-M^;�o�`�5bB�L1�3V��	g�)�޺0�Fz"o~�Ŗ,�0�=�V'�n�`ժ���F�WV���F��d���u)'����Au0���� f���L\ө��{� �=���8NL �M^n>Mo�=<_����!�*�d��l��������c�<���|_s�*�4ѭ��'��l���9j�
��2�.��e�|�̻S���a63#����d�� �-��)��ƕ$d�ןF����(�q<��a�e��Pp����(���?�p��R�<�7��b��.8������ ��瘕�u	����T�&\_JY��c�9fґ�]�苸�˸ �V>reg^:R�s��4�9�9��C��A焆@��+�D��I�&�n7����_��3� �"��Szs��)M�_L��+
uɶ�m�c��	O���4�>��q����K3���N&0�鯆�|��o
)�X�=�ɯ������T�K7s�?YD���]R��i��Mǵ�,��<ļ��ˇ^R����"��;�r���w;�~+������i�ܚf�b	���m��ОO����	әHx����T�5j�`Ғ(a`
c{�b���rM��#��|:�Z�2q��� # [f����nz�h#7_z+��8F�E��I*����pD��pدp��-~=�s=ֻ�>����WQ7��,D��A})@T���U�׶��pb�m{����X����RK��vsI�v�X�ϛ�
��" ���2s�t���m��]�BV��"W���I
cm^�\�o�ސ�Y�R�ih<���%M�#z� n?^T�ާ��Pd���&\zI_C��k�j4�<p*-C<]G�G�ً�k!��E�!'ԏ��a�Pa��Ƌ�o�LZ�Ikd��	}��ac�I��U�V6����l�����wu��)C��I�H�q�j�n��w
6Æ#॰��d��)f)��$X*zy�_���l��������29_������Jl��F�P�,���v�\\r9nf���������;d/�3�*,i���݌�h8��G�y])չC��	�f���W`�?��NՐ��`�d�Jz�6Y�4bs1	���w�i6 ��g���^@Ѩ@�|d�V��%Y��N	=�����Z�ꎾ��u�h
�	Q,�^ն�ў����3G�K����b��l�D�9��sC�y(�ҋz�N\x���5a:�^#sT2��:Ď�Uj������
l�P�6�y�#���V��[���wr4��8� ��-f��i��
} 5/3O&������f)���M[R�����{��a��nA�{�t�B6?�5��;�1��r�7uݹ��!�Ǫھ�Pj�!��06ebMn� �l3�)�lJ�t����q�^���9�O���}�B��㙤����u���ĴP�~���U�rw�Y/�N���R��N�2�7-;���o�� A
����3��fD�8T������ܬ��e���1�x�_�����g3��V&��f�R�j���G��Vjs�Q�"n�{��B5)#�*��}�]���}l��������.Z��Ɋ��<8ࢸϩ��X�S�r�	�`��Fb�պ*�+�Ff��$bB0�h z������Ҵ�(��A�P��`Q�\��+E�IIt�ہ��O��lJ2�`�]8^�߄��gz<�UT�{�)[������я��S����7 ���5��Tdl��ջf��{w���s��:Bww.�&�͚0���`m��T��J(�exx͇Y$T��)6�߬Yߨ�Ζ���C:��׵p����p��F^��탪�>�u����劒fá�#$t��[UVT���\�����A}��% �@���E>l���Ѽ򴨞�dʎ*�
��l�E�l�����5���}� &i	�6+h�29Doݲ
�a ����mԝ�S�Uմ�]�v=-�,;�.]�AR@�VT��xvDR�4_��s�������{�D{�
�?l�]9�1�����(\F�c��sȷ<3�1~�iW�N��ɘ9ڤ��G%�A����!&#�&F.���pDj�T�"�z�|�*�����? ���E8}?)��š�/�û&dV�W�D�*����D�PB,=kV��=A*
����%�;`��A-�շou?�0L�r��,��ƠJ&�O����Q`S�`�蕢ip�&h�ARq�ߑ9E�O4[�i�a�<� 2JI��,�*8��N2�z�(>��$����+֓�������4v	��<]�-V{��^�c���9�e����Z��������6-��oڿ����9޵���X�#�Ua7<Z�mYޯ���B<��&�<��="r��q���¦F���=��yɷ�<���'x�0gm��u��F�{=ǹ����?�cg{���k��"�%V�Ӌ��gK���m��h*`�:�e�e@Q��K���.C�x>��J���K�o�5��l>�főO�\�	��n�s\3P����!�kY�uSl��	ْ���d�ph}�B�J��RvB��.��}��C~�b�X._$6o�e�|�������ވ¯0��豴��\co��e@Q�R��GM`=O|�]7�Q�S��4��8���lG{?���!�Ue# ~��8t7l����6�:����g5~��`2xY�:��Zn��% ���*�g)Ca�����D$�4�p�@@�!���G�:Sv��t�9�����(�V�����l�	z0&�r�����#i����/FM*W��n�i��7KK2�ٯ؋b���
Vv1�f�"7C�1
