// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YSrGusU9cE2n72SX5zJ4GRB5UnfxriwkzryLi684g9JTcv5TayHKL/fRnyksN/rV
WV4dQIhFhYie0b4PZ4VaaasOlWChO6jqG1wBju5a0QIB+VkAwVT1ILYeWVWzjWB5
WlUcLZse3owfTrSb+Zt3HVzQwCR3X+jHwNbhd3R5JkE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7232)
Ajz9vvvuLX1Wg6vXOsbHueJOU4ENFyEJjJ4xa2eT4uGrqu6t+JTifQ3/aakJnvYk
u7hU0tot1F/XSCeR8rx9CtOyKQ+90/2h167osizpHsuIoNqnTozG2qJvUBPbgkJK
Mla4f5ABxsZI7EXypY07JA7tH190j8TEzZff25hUy5BBaNnj8Edqx6V1+NkZCsAM
0ikw186j/R6UGZLKqexDBlVjXX+qXu09cg8F2oE3AMEZA4hNd+GDahM0SVRePe+T
nuFgbGzfKW86jczoH2CY6blZ0Vu2oyAN3HLnIxMY+Fe+7P4Kyc8XY2KtA0mMCpKd
VdU7gtIjzUnh/JSgiWXw8gCsYW0IlWGUydRn4FqhQGt4eqRVSuL/YVmBc6OqNQCI
cvamWvWPwgdZcPLaWsv5H9rarYS0aiAKY5D/lEOYShg+yN8YCsfCrTnFNMRvJfi5
/n+fVxf4AnLs2/3wWX7z2rs31dyJ5m34dkjGKNoqIHl2bQ+0uNac2GPQlh3WpdZP
K/y9E4RiESpWUyQemD3UWH+w50yPO5V1jEBObr8d8D7jDKETApIPS7BnGjbmk6Q5
lyZg+Xk0zoVYmBdl8lsWUhqbaOBcNF8H/d2806EOglvnYC2uyJ/8Aeb6WF9ihMxf
ElNIE0AdHmRD+TJMSn54uoACC+ahu6/YlJnVU3e7f9F4VO+KGsRbfEW/8tSd01I6
iucMlFMT00XpNy+1beALnw0BDpHATCEHHBARNGkooctdi/DUkYl18fCzUXEe+k1T
aMQiRpco3K8ipTqYjZhrR7L8HVwxUTsVpSC9ocLuEkcxAoanSqr/qIfsOUt/u8gL
WkkNXZd2K/sbu1kGtGb+lwl9fVOsgisJ+wbQ0QB+HnTBS5boWqkxqPH0Bib6qBaj
JlFoH4N5ZgHddOc8zFEHi0izdu8IXOGnW/7K3c/+C9kXp5jrArUJXZrdEs6U0i5a
OXTkUkTXy+TeoQAL0DJvTF+HRAfp0KuFG487lP+Ft4JNwyidJt37Id547v6qjOdF
av7z4dIMOi77AEfo99+/f4y20lLVUgI5WF8MEZ50WE0NXWSnYrtD6tLz57eTdUps
gnEb0JXleL1vqAnt5mB38C2DkdYEDjAQiAIg2wgBB4gdqMVMS8FY9jKptHnvGaY6
KWE4dEnSXVhNQCS5cSVYn3nERsuB07+4dbFCQD88tXviqqsLou0hLmvGq8hPMz5n
TCoXP6vIejZ+7wPQeqPwhbc17ea8m3caG/9NM6alddaVf3c75GG3duBpFdSk04p/
auAvNMSsQx53QX1IAEcEn+t/V9iCcm66m41rydxhhPxbAJVH1pCwvWZUGNk9PFpD
fJphyh1x0X38j/nai5iolCrnPSUE0htg1fzVWWbWT76MvVer1dwXGyQlVPQnWuhe
z/AwSAKS/PMw0ECKrwAdlSYup5yDTszO7sSiMesm/1Nr7WidprMRPgbsxR2TQhBQ
DkEifJUqUlcZ2Rw8xCd9hw8M2utdbXK4Vae3TLQ6LVQlLLrqHmVMRgpZa+tUbz1j
OCAF70Xho6RgtjttWwMnR9foJMRPhBznaroow0HM5Zlwvm+pN46FLVCyIr+19oQ/
ET/XKaDJ5t6DQEv0WksvjPYUuLtYD7QMD0P+PATkgczVTadDEXygwSn4SduS98ZB
vSVd50Lz4f6tTVjZ/UKoo87/50g845DtDNeSyEhuyZvm5YK9RJVtEGI13LkdLkfZ
F0G2Eg10SpWZNq8g8vu9a9yuzZQabTK9OZEhldgeo3YIz0JxFtohJxld0/3BYA07
oOb/oFhrdKQOBG0Vtn9EexeEYbnoamL5UPIAEE1hunKlyKm1eDub0S1boPylLhQf
P8H4F0F4397tWnX9bLoqsGLInS0T2tfIBqX9cGdtw8uB9KJyKwMw6nGSUkFGnS3k
h2Qk0pCw/vjlz8XujU4VCQNHR2hH8A0BF+QPQvOhOtAFLEOJkKk9OLvr6zBn9cY2
Xnd8+2L8U7Z252lHa6jQGa6X1+BkUvKlN1v+hgrBKVXyqDrn1wbM4zrfSd/0uG6r
o+eAs9xowfBhRAuXnldqqrr3mjPO5ovjfuZRpJKnk7qd8tTiuPBDhAg1YgMj9JTR
uRM1GbR2jelOEkPI7aMrUL/ClPUx3Unqk45BtE7ub6sVpkHOt70S1WDPTgJh9LuH
gDyyAP6NZaNJj8XiZf/s1uniLh8+K/pgBreFbs9xQYXOCVtMM7p9fH+QxRo0LaWW
h9f3g3PcyJAuMB7VZz1MnsJ1r8V3auMC3x/sKfgNslo9jwqXIG7jo7OcSuv8DYcb
NtXUoT2bnH1OBfJc98GUQNi1YFNYMCSgU0GDsRKVZTF4X/aGRtmTQiETpKIskrkK
OekLAqqvJ7QYxEocdZ2wGMZRc/09NJrRCOemGbw+ROCi3OLiYlHrsB9NH8IRTSGF
4LJ3K9+EydC9C7/Pf5BnCGnjV419CRcqb/Qs6ysCLbQi1qzQFrBeNxs0ZpZgqNNA
FHKacilZ6UWTPtzMhQOwL8c+rAJU9VrBgLgDULLcvazaeQcc4cRd7BG7TQ6oU9JW
ERpFaktxS/kEIXziYD8wQe+u2+v8NaXp7/KAeGh/3kd67h5lCDbfBiT+2kuJKoc+
e2Fw2M+3x+qWQpwHYuUBTPX81TrMau2XYRfPMmZ7aGQL48vouf0RZEqVyze/bCqL
MvnZtNiIbbAawru+6aYuEg9mufcBRheKHql9jm/zkEIlInrtOF9nFgQZkCPwQhXp
1Dot8cjldrhPyXgfqCo4//b4/0jpylcFpCqqETqi2uJf5MoDU+8rgzz4R+gg1zUg
jajQtIWi2I+bn2PiH4Q3XYL/ODGYlUwNWnpWAhsdq2Zksbqv6lX8+j6Pe2icEFj1
vRhPOo0hNi/Z2viq8Qg0eX0ta2xOKlwlqOihZupZxH2nHSgkaaysZJ12Xr+uhfc3
Xx97pspZOi6iQqSqMivdINmlS/EFLrNAOBVUP4/P+JF8l2twQj4Q9DryGW/utImz
dHJZMbwkXQ4gPjn2bGgXMXp+apF3PXGtoP1QJEJ6l34BmNzIntBb3Gri3zO6QcNx
t4+/hmV7K2491RofOmVdM5NaosO+mFqULQKYuciLbiGhzIIfgWBG58qzPy7GFacf
z9wb0bO8sv5O6W5s2CpqQQXvzN8gj0S21fEtpUl8MqTiE8K0s6sABU3nUCBz8Km5
lcibOCBAgyQhELg1l2xssEyiUVlPSB1nAA+UfAwAVu+1NGnnbSMCxIKjCXg/Pgll
pzkfTLoAFnYRFaJZKNT81LL1UTFq+IgUA/3kRTpztXbLCH018ZpWtpbk802dHkKy
CTvTLnVcz7eTOtx7qMuv2DoSm51K/l3BpOy/TMBJJWFtIqcZ4jQVgqydU9GD7od+
rtC59WeTU7dlnvP9TbyNbyQHAFTPtl8pRO2dBbSu0i0JRtYGQgezvW6MQGrfZlDE
+YX8y1yvfgtAWA/n4yYq74mXZDds2ezi1fHAR/qkyUU0ANmILgvd5tnjT0G6H9dK
YEWVT7pzaRNilRJUifF9EAt4pq0WG/syuUbIoJDTEC9mmPwaI+b1x5bYMsmnpAcH
r9vhTQ/Fketv8yQQZ0VtvW5Y49qygBARpLgxnKwgdmHIVvmjcCQ0QQfCAzg6nOzR
Vyb9rtZCJ90BTZGK+sd9HU8uoMHip9Vvriepbv+GDNvG6NJTmEfL1F4JdY5MOMvW
42kZlUSgLe989yHqtcgfjwQHMDLKVwS41w7OyEO7hArNp7N76O2BtQxV+7aKgxUt
v3gZXH9j9hk3GmQEPSwMmUuyQBRLh9hluqaCey78AfO23WLEO9cFp7kbVTuoH/7O
ycKcsbSoIfCpslPya/KYjNpdYS6IHCXmjTJ7TWXyFnbVLBFlVfM4eX1C/C4P+43t
UNoiU8/HHMdgT/imf/Qzb4YF9qVayTfCUYbU5//u5htZtoFM+xPFRtxvCAwmUEUh
OxizxvMOU+GrFYHYc1LY454CqZ0KzqPczPPGZspK9en3QWq8vGj+jc/GFUDV7NKd
Ttm1UKDTmj8olUrWr6sf4r1N41JG+cIagbsgl7oFSxuWbIasgJyt29bA6F2obemM
/b+7TipTvIaeZuqXcvm1ouRoTzg78iWFISIR/zFoifVYcdXbUqF7qoNrA5wuCrVe
Asf3Px5G4ZqtIHvleqCr9E7Mf81d7/7qmsPUDON581PNhW5W8mYqRE2qtIzU1YuB
z+HJnVNrU4ceaaShMcy5gYhYJFi0n6VJ+7Pq/mCDvkYgngaMTbJ1dxDC/IH7SOeB
fRLxqHUPlLiRRu8fFu1P4GOvyW03dg8JN52bnUWmnogVbnHdgFcHjQVZkONi8Yr4
RtbNYVd655s4I/br6ZoOfS8dAHT0BTK5Y1g9MuFr6Kzc+DYFyqqFlT/tbZpeEqMm
1tkMujWrbXzwEIXKT9I34yWD/SqcRrcfDVvn5xhtlqKTlzVBsGdodf07PYL+i+e6
ZNx/PlPYvFDqiUn3qNtx9eAcXIgVgfEcYHhA2h2eZwSrNuUL8WhNkKDMnfrUq/tq
mL306yjZUx8Oqase4pJ7iYihgacWljhWWOQHPZD5XJm4LNUQZbIphhOYWVmAyQj0
LiqyIS5fOEqJExcMejcamo2x40OfRtIMF6UhLMKhRAAjwJfqnOk9Us5ybf0uWWLl
79GX0JqQVH0etbG7c/gYLp/C7Al3wvoFf3yZjauMoa0gzyvG0QQsgK88H1yRC/Rp
ozxsQlszemaHJeWK4mP8QE5gmmsGVFpLqqyeo7aGV/Cp+Q7pvKRISyFHollgQlgB
0FnSIPzmWycHhux8j1tw5RdH0s7C71lHIQugWXAxGgmVEAsAVPE2ZvKDrrygCDvt
OMvBSbWETGvEMLYA3UmiI/zDYwMU9NeBv+Yo+wdApraZEYsF3s8s6hIqVBqM5Ry2
o++3YWmD5VpUYmLlaKzhJKwk/x5FmoxkGbb0YViKXmf5XpX7k2Q2OEHSYYDCkARH
hzj9SVusQpx1pchEFnfxbRkAy50BDLE3b6z18qi9NqNtagnpH3UsCQaMNFyxSCJY
hs+ji4oJZzLdvLiIyXZYn6m/kIJM5/ulaM46W1f+QTPJCkeIo3veMz4OhOXGhZ7R
s7R5hzJN0OEjU3PiCBIDC724RYT24SVlgs1ZijVVU8YHHLt+FS+YPww3U6hj+SAI
v/2Q/BgRNFrHUmt8JbQjKij/ZKTnKkCsFMMAOyp5/OV29Al/XMgDn0ITuMCvbxSt
MM1S6vs7C/Ytxa17S8sLApVuKSesKkP9I3LxKf8hdKYtSpYYa4ckCZ8uRO2WBaNa
LAISEuOqViLe9ezGG9RwygjraDuFxE+cq2nD6ljVPLGPJBa9E/fEAGvN2xkLxiQB
HUQret2flKipqgBYsPy125shdYMsWuYI6Qa3ZjHoBAZ2EDQGjmkyLIZDW/ufcj/u
WdO0sCECAaMDb1lsyMmEK1SFxhMVPQaqms7qYRbnqNbjDkl0/niw89r56GOZDkIn
z51uPDKrGYqsezWVg1C13gUrCP4ZpSir3KbLf7SciHbYEd6lEUdNBBOI1L7TSTZr
V2R5MqAYiDi+PM3btMkHN76xu+TWlRISI8ALqa36MVyLHCCwxhNgN9C+RmjLR4rV
vYlZ44DBkDdI5Yyxrc+Y/WKaPEnSXh9YGgbFuPZG81lxTC5kl5GrkZ7nKu8rHOEh
9+bY1DFXGDNSv5vZVWHsc3LneTl6SbgHvu9qQCYKWvUlWglqUnzMXWZz4kdCZncM
mUtiz1By7ysY09ojnSpjMX6XJ8E1blg9R7gWZrKDSCYB6qGyK2uPUPbJ90Rmbqf5
l/Uu/nfnHVRlbtbZOWq1qe9S/e9pD0Uymisy39H3tlCi33p5UIp4iqJI0ygbC3FS
Zm5NXFo4wMl6rI1eVrbORloAJBAPIXWKEca0VKXY3lTDuImfXDTy1nCcSMz2YsPQ
Kho+Egh7iRGmbSUa8+behOUwaZ99H694SY6zRKDg3P5JSxvlCdhlMHgWICm4XFjl
rrdlpXrluM/D268DgWVv6siZR+DMiZ1ojtAlxWJsc1OClKBi/g/OmlIV3F/C643K
TRF/guYWgJ7co6AaCzk49wA4eW/iPmj0ir9VXwZg3Hn5XfGyq5EdSdLZNHZK1gNh
dHNBks+G/RR1hr7LtVzSCTa4sX38sBguUOupXLtJEQueqDjjhBudRkEdkeXunOn8
dFN/mz3XFkg+AGe7w9pPFOGt6QxE7uPFDNVIqj4FxGo2cTJiZ4p7wkQUO5HEAGGL
6QtOcsYpugsQhDTrh7aabMKxsTO3baFww0RWEZKI75VEsIafQtv0t+eB1nwxXgTe
mE6I9UAHVrA7ESH9k7c+qJVhU8BRnNkunOH0u5Ij0GEraJiqDCwU+fAoR3q3Xl1c
KzAPIGJcxYLHGMKZ7NZkTku69jJdeAoZgh5HmgED189GBf86cQLttOU2ArDwm2SP
Db73APrXl6UrrKSoNcN/wv9bEcdnXmOCqJwCtEMlIJPeH6Lfg7JB+5W8/hc1eTlt
5rBC1YYtmhqmgYx4JVzLy3yZcRXo9EzSxO4UNVR3wza/4Bp8nqQl06Jf8i90b+y3
k1ia6J2GsoB80ekpFv5f4GC4axX6j3+ZhOlvoGzL01hnEmS3qnqGIX2OBxtjNLJx
N1ZduKEbBSDIE7Lpwz3UyezT80xuLTUcN423spQ3ZfpiGSpTi8iHhFzESXTFRx6n
dTJP7JysWI98oadPi9QEAj7Kl7AKFT6kXrRf9I3Cep3/IVMl47m60Zm6F3gBH5HG
qprwrCRXgUbtWY/oxkWDQERGwaOZnJQzAVYgvhyoJ9VAmlT8mUWD8rgow9A3sZ6T
7HEL5fso7gO1tJusTBTuCDljQvtrnbNpWRAX2xjD2AbZDwz/XMLa70wOXWzyX0Wf
wUaox9MOwHS0oZlwCNNjqcF8o9NVhrL1RRsslHq1w/g0zYnOjyfr3he3xS53KTxo
1ph3iPROd/y16AIiwuvA2EQtRPd5EFAIYjzjiNy7cu8Xm5R75vTdYcYm1MsvUPDQ
5IbbK2yID9k794YNejqqg5UcmHzcrNQXvRiiIg6CKtkjpMzpkpDrU4aniLiGy3He
3diVe6EuvVW1VErfcl7atG+xlKXsWFQLRXERQm0AHLZoz0EdLB5En86IbSJ9CktU
k+p5IWSwyDbP5OFSD6TohYtuqexwfAkyzddVg41Oc4+5Idp+4BbydjGhv03IJ8jH
A/6pNOVL1mUTMfB/F2aqvyxp00lS7URa4NNPIcAxNQyanx40KLrVd273C1Ojv7ht
lJlLRtoqA46C/LqIeoSiV5VLWzKy6MJJ6akrm2fMI+5FNeQPwAfTb+7CjtfHo6/q
3s9uTfVgTJpQ/h/hQ+loIKPuUFepZ4WH4czl9KJxPieZFLDqhn4G5sutMfWNZgC8
9qaFl0WQKAbkoOMuG1CaXz+f8sGWMUjNXk4l1qyPZ/UA4MYZKxbH3UUSiIaQD/eq
wNZq79At81usG8a78GZtVLIrzweU8xMzU0OPNA5ikSEgSj9K+tX3EmM/a0TqIVOS
16ocO+R0T29ZHHPEQNIbRwXgQbcmuPKKchtOKhv3DkgLZ4kBdIwHhERVPN/+i4zO
syhy4CMThJtKhH8R723xjn7y3/cz0be4BDAGVs30UZ4Gl8rPD3P4BXgOOEqQjiM0
fFrI4PM7ZMuZLQjVPQjxPfRXMlAlvmnqGQjHEIgFi/io1/RkZLPdF7b61G6Rzo0k
brHuN2G/GMakFy3lVgy+YvOTuMsenUNSYpvU8fC5kG7XtQPmpWmqk9v7IqKNtbFO
+bfEEcNFeWcsUgYj1+wzFJN9dIcRT5Ki4wTHDQhN0ukFLlga4NZUWlAVTrYMLg/L
oVYJUx/oFeJpbzkkEmu2lWcpx4BIATrje1MV4UzC4BpBv5o4HoLzgdNZwn2J5x8G
MRgdfuDXEIEewCMSTP55MKH2CCnAX0FuJW1QufWntDNDsMWEigoelUr0CH9p25nA
92AbRGukIYIopSy5n4yOFTRmhKSnvW2BkZQEUjcJ0BNReuOoyBNVDbHIgC0/gy2m
im0j/ZwjjTR61LkuQTdQX6R0O3yNAXats3Y9iN83ipnFDZDw3Y0sFdp1O8H+MpBo
eLrSqz/ohCerN6OBnWJ1Az4uWYhqyBG1mxJgqm+NYDqF4IkD5/62NCIAUmrpRdNn
o9oIpHTGKGslWhpUgM+iFlgZL07+bTJnsuocHHmqQTVoLzD+RGRt9tKyI4Ubczxx
iKE40dfkmlJCbWWQMZHsNxGGq7JJjuPDqPuGgRqbVb4VvfdLdbLUzSXmYtbeR0Rd
cMIK/paZWfMN/znM6UrYmvR5Obm117OFKj4UOOGz7PdCHQK5ShgZTfnuo9qJSP9k
4qYV8nQiIPf9TVZDfVWtAtiIGIiLf10ArXyqOsAs/c1swU1z3yOFueQwXa/GOY/n
J6zg6UVrqfF/1gL1AB9FyjX9wZpS/n2FWavCSzC28pIKdHE93eUcCaU2fFJiHbr8
OnAlGBu+NBch3WtH8FUJsjS0AKE4xRv2hAZOf7MOhypLaJ0HDAnwNPRic2+epjng
XGGbZVtV5ZfNmtTHibRPbhkez8Oeeb8cH3BKvgTPP06xMlt+Yw6F9ay9bNACWJ7z
xfm7PDC2tb9oLaDRK1XRknv25NfoiKKHaKUWvTd5DGoc8Qhnx9qOAmCxXwKen/Ih
twh2Rh+F0PsiNS+CV/JCSDyaLC0TTIGWnuh8Kp2thpRsEdJyB/ORjT+xzmlh57Vg
7lIvu/yWwVfwycnKRc12fNLFig/AOAT1ryZklsMVPNV6SVAoxzaWcbucIEwB9nkV
Wvza5mMvcagz8PDrAvf/P/scFZGk1kPolvWQmPvSudbBeH158KceSj4GWJQI/IWi
rF2+MobqwgDoheYnpLPwat1xPXi7ILFIGKq4JQhrcwLs/U72adXNKEAabhzoEx2I
7cbe8YNi0i2pdF6yhTSqFoGc59II3rJmvphf2NvN8zkAXBg/jjizcuydXYvi/lIo
9v5vjlnoAoaYZQs1Zm7HsCZvodEZDRu/DSnqIo3PxCJjbWSStoWTJOSpGZGilvy2
N/KdqQv/+RBI+w4+0nKFfvuTFYfwdv/V8hrP1JeccRsj5Ccg/r25FgvzsDjb1hpk
rrs8GhpDdaSPZIJPl6tn3q1rojcFjrYTazrClPwHu+NbGBxDFQVfrokz6+41q0hL
0w9eil8ZtcIGE4tOtsiRTV5Qi+9ZBjxk9QOczKr5XffIkjoJUrk7cGv3uvKUmdgI
z8+Ms6Ifa5NpSwCZqxWLZs3C6o+NzjcSUETiRSUCKKgKSTwlAX5dshc63koDQcoZ
gm1MPEyKX3UAjUcWxzarcru2sExAqFZ8TMM0wzvRuHC4YOhxeihYossAqGdQqyzx
ma/XR2AzAjOM45HtiYO0qP3fxxLNsEd4XuF/PGESDxYf7ByjEbvl70xuCN/3tDxD
4nc5+wby8A0ePV2zIJMY72iIG76AbU3Xor9/ryAkGqSYNtiE2STXUZ8e6tZfbJcP
s6ltCc7cgjLzJY9oRrt+vpNUiCigHvjf2i+paEDiOo5LNBsFzXDuhxBChWn9lXgm
45YgzoAmTmVSAzrn9LShcx/+IgtV0hVk7eYpGSOFqcc=
`pragma protect end_protected
