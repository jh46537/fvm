��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O!) ���Y�Q΄�O��*Ȣy�dsuQ���`�Q}SA[�.���(��<
vɼ��;4���͋s1D[
�f�T�[��h�K�"HO�¤�TwƜ|�J�tR:����p�#��;������A&�K��HȮ�!!@<Ȍ��VV ��k��ko窿ae����ZS(�F�FO��2�;Z=��t�)W�{yo��r��(�K�StcN.�����s{P�8��AN�C�/��~Y����[#�z�bEB97�'���?�$'�����ِ��ǰ[�'�d�X�������%��`r��`���8D�]�At���w	V�򴴌���R����F8[4Nj7�-���ιFUEp�]c��$W��9P�|�Ԝ��L�?�9�8	^rA�Ƿ���.�He���n0�u�+}@I�2��P%p���-���6��f�8Џb̝h����喥e n/&ρ�1��ue��Fw�����s���Sܿq󀷀�	�~��ݒ�-i�Ȳ�G���S1	�g��<�ד��f�t0-I���:oۼQ gD1M隬it�;y����4_���TB�چ���thh�bL0���]q~�����4�Pw��Du,��8n�,�045��u�3`G��볮��"�W����`�hR�u��yI&n��xc���&����7���W>=���Ű��T��+�ς7
�73�ȥP#�lm��"8:�K4�j��c��<��d�eA����
���&c.�nP�	�hy�Q� ��l54ꓭ��ٶ���j'bz~�������,��������&l$� �+��D}�4j̢�0��)z���#ef �2)AuO�3�ۉ��p���s�l,��p�J\W?��sk\���k��}�a�.�.i]�q��W���o��9�����^+@���T�ӷ1m�$�X��<�j更�UGk�y��b��}���8uw�h�R�b"㕑I`}�0B���B��v��u0ۇ���A@��D����N�Zۊ5&] ����I��-�K���_å��HҚlL#��^�p�wo�O!�`'����^6y1^��m��7���s�5���"����BM�&+��#��_����'k.�A�$ʎ����ąI�4Nj�^��Ⱦ��4�e�zg�J �Ty�hL�%� 桐e�L��ɏ3�jyBh��ߕtͼA+�)Y-��Ż��/<� �q�:�gF��Z�>�I����O��s:7 `P���-��H_uuN�~>�k*�(Z3�Kx
�r��_:ߺ���
\	��L&������h]G?S�3q%�D�5����Y�3�V�½ˎ��X �t�g�l���ȯ�����y) �'��(m.�<����|���y:�;�Mj�,�;�m+ �{g��T�c_�T{b�2�'A�o�V��[����١�2s��8
���j���e+R�<�_Y�lQ%�t7J���F5��{��hj�dR�0z��n�VVWH<=a����]C�3l��6T�g�+����!2Ρ��V/���������x6���(4:)�h��Q��S,��p�v�D�5���0�k�������x�/��{?�]M��bDtbg��w��ڻh; g���v1�r+��'�:bv��O�0,�a�-5UbZ�%1�6��vQ��>�6�r�,d��T0�6%Nz�����uGGf-> ��f����W�̣�=�ʑ�]�̈́��&�|�1o�ПWZwvei0�t1�ڗEg�$���N���/��y;y��A9�.G�a������'N�0��\������X�)�UA�?�O��*�d�ֻ+vkM�~%O��5�Z�vOwam�T���%A���1�$���9�O�������1�fuF��)Fp�t����_	����x�)La���꧍��#
-�3�v�"2��
/JiS�#��1�iA��W���<z���y��6�hޘOø9�d��T�G�����Td?z,�dJ�JpVZKM��Qs����9�V�����k�PJ>#�#����E�E�qw�d��v^u��ˊ�@��t�ȫZ����4�^��-��R��DH�@�Ȗ7W�s����d�-o�j�d���D�j�V�3��7U�2e�]9 0���5bo��=Y��T^λ@UFŮ���c����=�;.#�J�����(@,&�(�v۞��bs���8�a�=��ݙ�a?��c�7�R+�K����*�8{jT��(m#��u�^���7�Cx�$��׍ݛO����{���o�n�� ���5����
� �� _�
���,��{��in
�)��j|�7R��F
�x�D�IiH�g�t��&��K���\00�$_���@�S�fH��(�O[�l�W��wd���B��t����G͆��O�At>O��3Z�5���c.��мnT��_t��
��,��C{f[!'X<4VN�gܱ�5,^�I,�8��c��Q����O�GR���z�ڇ�#w8i����d��!
�>�zQ)��Bɘ����:�����cÄ�/K"5���o��8k��Y�Eqss�r)�65����4i�l
T�*��U�J�"l�B�Kx�H9���C�]�p�q� �2����0��F��t��ݍnǧZ�j?����DC�&�!,�4cij�*ZeE��8��/�� �[I��S�i5��65�z�d?%Om07a#�����hWM����ZH�hF�B�=�r\#��b
���|{�-�A$(�W[-3�g5]�D+�8$,��gh鷬U/_��']�	�l4�=�J ��_���R��|B[L;�^�����} ��q�������7/�U�d���?���@���sQ8��WOY���f�(ң�G=��iP7�73y�R��	@�0�����~	�I&b�:ڔ&�Ռ��HT�:Fa:���=��ka�-��"N�q�5�V8��骨��7s;;�|/�܆��i�[�0Ii��[���� z�
H5��9��ߓ�k+Q�/��������΍!��Zmѫ���0��G��M�6"=�����*�Sg�n��h uv>��J�4 H]�6��6�ou���{��ς����G��G�,�j�?r���L��H�`F��l�bX��L	�:c���c�������n#�@~�W�ΑGE��#�ۚ5f(�f�祋�fU*KIMM��%��M�W&|x����[�|����Q\:f@m%�DaPU���җ�/m1�9��>9W�~��0��Q�H"��d�C��R^%ږ���h����]�|��V�aă覐�29Z�x�EY��-D�&o��x ������-�|�(p���(
Mu�p�-2@6a������"Pulȗ$[�<�EeĔ~Õ��`�� �1�yʙqu�"]a5�Λ�3u�/G���d��G�Q�'RX��8ר�A��a��|�������i�^�ۗ	��B�F�
F7hF#�w���u��T�F1X;��Y�͙�d�� ɦgJ� �(���LZ�دG��&�=E����Os9�A`�yHm:ڕ
�I��x��OFpj��t��a�\Bʱ!�rJ��`IУ3���<T��Ģ�Ϣg©�@#5,(��٣��ۜ��_}�Y^ј��[4�[^a��|ܷF�Do,������B�v�~$Q�ļȣӒ���@��n�$(v�Yf;D�gJ�(���^�ꙛ.TA3xfjj�ﻝ�I}2��\�\QQ�Z/�k����a��+1���N�,�v{>�lB��k�|\�b������f�҉��q���~�^Bҡ�3�O��%��굁"�&�����k��E7.��<	q��%�Ѩ:[*�L�C�6ȰNg��ѥ��Q����W}y��6+�*"`�/o��C����b�(�.��7�v[5��B*���?�[(V` .; f"�� Ϸ��*��ǣ>�)�U�Ŕ	�n p�RN��`kH������ J�~*!�K�Đ���9�J��ظ�M�l�СF!D>,o����(Pq�u�TX#�&�j�{؏���娖&�G��᳜4Aؔ���C����
�U��1�y��$�B�0�o-B��R}w�2@�� wj���tT�&>��pI	
� {�P���;U챎�V�w�P��1�����qg�/3+@�7������Be�s�9_�Mq����wx���=���ܻG�@���b�ɺ��3W���'�&d��d��m7��Jϛ�c���ΰ����NY��������m_�&��҂����JB15���z1�D?��X_�Z,�(�tJ���%����,2m�7���o�z<�r�����B[����]:���
��FC��dT{�WQ�Y�U�Q�
%�ko��\��-"�R�ƥ.S!�GL���Gj�pS�`=�L�[�����=��AL�hnۂ]8\o4����mhwB��b�ZwJ!<������e"j-��`���)�Y@�ڝ#�!�6jU
&OE �C`���2��U,�����@5!�l~F������*G��i!���Ј4��P���Њ`�f���7��<F�.qWX�aq������gy9�u�?�#3����7^�~�d��_?�h�W�#	W��I}D�.U��m�?���?E�莜�V�shc�P��;Hm�uF
Q������[Ƀ�Rt�BWޤ&�t<�.�Y��Fץ��k����d�I�e��^6��ɇl�B��k�˔������םǖѣ8ڡ��X���h^M�SC�,eC��Dt�-3L-/��{������s�d���e�ʽ�A!�%�lG�:od*Y��-�
�o��x�Zt��@ʟ%@���t���X��ˑ�rh���xeQ@ېņܯ��/�:�mt��'���ӳ���k$6��=�)'��m_�X�� �c,�:�2��/m�R}<�>�K1�Y�����TK��ckE�e�3�]��":tq��,#�&
��T���ʩj�A	 Fצ�;�,�jhR]u�B<���#C�.5$]���f�ݡ꟦F���b<�)�]}d��\ԩ�������E���9W+i�g�LU���;��m�
g��1h�1d-���P �UxD��f�-��rC㍙;�$OC�h/@�~|�D*�c����C>"������liI�dw�g���j�>�/���k@��O��O�?���Եy�&��6�O�oÔ��)5O�fT������3%l���d �jGP���׃bB5�-7Շ4�;�|k���E�k����_�s$�e��!Śq�+��	9�GX�����j:�5�s�v���JZ���է��[�p�c�! ��>�����Z>[�w\��x�d�7�I�Fb��o��hl-^^	>zB��\^:�i��{����r��)ʥKOXE����ct��љ��w��c��Rn���ߎ��OX�f{�)�w������ղI̟'8�߳�*�বP_4n�F�w^�<�Aa[)�:�i���_��*�d`��`��^����#Bd0dB����� ��Nh�M�����'�hb�V	����dK��E����(Ⱥmg����)7N��dΈc�wx=�Р�:坷sz�G��|>��<��um�wNḧ́�=?Z�Ý���$̓#�Ӛ��*�xil`����J�g�f�NxQ��S�|�UTV�o#��B� ���|[��K�$�PB�1�il�P�M��Ԧ݋��h�C8����	%2~�s,'���fxR��U�:���؜8�1E���r�6T\׾�+�c�,��� 
����1���M"���y3r~g.�b��ЇOԊ�I�F/�g�U���̘��Y�.�*��+vH��ڰDP�����;�.yV1u?p"����V�$.���g�#�5k�h�yV��2{�Bb�f�)/��y�z�2�K���U�qm㯯��bs��,�^�i2u�.z�ݦ�{��Ri��jEc�����Ү���Uxߍm��
F���mR�=�6�5,b�O�])�Na��6�@���p<(��ٵ��;R�B\8<�����q��{��\�� /��o7l��a�
o���5��������-;q����@�(j]9 &��,�L\�
�Ժ|��W_m��$#-��q@�ӆK��x�#������s����N�Ty�7������#���B��֜�R0�R�|���܃����<�b��iD�Bq��_:���8�9�E��d�`(��װQG�f�k{�jC�;������ˋ׆�SYIz�]�@�ƵJ�34�Љ����m�����g�+�6k0E 	�9%g�f��iI)��q�����>R`�3(m�34�]d�G�G��Fэc<99�.vOʹNy�\��R#�?�HPw�Ie�� �yF��S
&���=���8���{�=�4�.��*��V?@����[��<�ZB����<�Gf��v�m�@�i�+[W1&z=I������f������-5G�ã]��J���/�m$�)s����t��W��9�r����yIE�E���b�s��
I�,��(�~� Lߠ�5����Bh��@p쁨f�?;b4�on��~�N ��0�%�9NN�´�j��i @�զ;�����P���7f�u����N�W|�P�Ԍ����Hԥ��$�5/��<ֿ(�?QU�Uҧ��M��Ld�ʷ��
}v�.j������
�I6��u8j�m��zj|e���d��ԙ��I?hs�ɷu^P
gFfF3����q�u���c��Ќ�7��Ir�2߾l���Y|���_�&c��M��O�z��h�+U�-�ڴ�$��@YPb^����$R�b8=�?J6�G���䑼ܲ-ra�G�Q0OoK����d}_n��n>��U��#2�_G��`�-x�����cP��d��
�NxLh�],��u�_%J�o�� .wٺ�.c�(�g�o�o�b*��,���=qT�
L�k߂�H% ݳU�i�l�WPR0xA�(|;]����&�C�pL�H0���$h�W�FV'q^K���A��Gm*�P�7��쉤4�ӕ�eۖ���nÌ��T"�<��_U�����x����@���\j$?�O���m�>g���%�?��m�1���2!�2Y��H"3W�5ɂ�.��.�R��Ji]!8�(4o�um�/z���8��-:J8[��	��/d�>IE˂p|�s�d�g���0AP�װ�k�c�Nދa��
���
� �D���S��K�����XNz�?ښEhO|�u�{[!�/n�UB�~�n��,i��/����FW��#[̓����eS�G�d�">�#k ,�����(�ZZ&���<��n�@h�vJl�0H鿿E�-Vb�֐��������L�vh? �g8(����s
�ӄr�q�{��F�Ѷ�U��p������k7�d�����<V����kLVO�A��*�9V��i��B&��ņ�¿�/[����(�A�B�r�T�/ʛ��Y.?"Y��6r�����`ijWy.�1�Ǳ�S�â��	�
���?r�Lup�EO/��97�Kj�~�Y��9/���J�����mI�Q�N����K�ab$�J���9+a�_g@0�Rk�!�w%��S7&��B�?`��
���sS�kZƐ!�i���-4OB6�o�/-�P��Wc��"��>���jC��ت<���%18�dݒ��Y�51���4�k�P���=�*�=�.�qu��0��[��¤��sj|QŻ޶�]����J�o��s�.�� ��yu)��E�6�?�}O�O�	h������'ߵ�Mr���iR(�c����h�:V) o��q���k�$��9�i��s]d�..b&��
��L:�,�q�q��r�0��5���˚ 7i׿�n�L�&��"������}����dgO���!5��#�&��N��N�W,��j8�6��B$�l�Ш˼�ǕΉQi+xv0�-��
�.�����a��ư��U/,�r���
EU��1(���\&EH=�+;f�N�EV�]���ͮ��P��`tW�5	lO��w[��ÜVea��i�Q/~�.�Y� x�2��ٌ�~p�E�-Ǭ�z��~�YV�Ml��}U�9�q
�
%�*��l����iS��w���e�ثQ�x�?�̿�HM �$B�d�R��P�\�&b��UR8��K��冭<�F�[�ȥ'ſ��:@,�O_�~��Oh#�Gh4FU}��ʹ��������8�,���/Ϡ̄ �����.�m8������;~��i @�0��Nlzc�9�	nr���2�� ���<T��$` �'��W�0^�����%�������5�zU�ا��nc5?&�Ѥ,�&�+޶�b���Ʃw�QK�/"��>���ׅq(E�ޚ?�-�lu3*����[p.�5Eh~�E�nk4;s'j�~t�Oc��)m=���e<�T��
Ny�8���g$'�me����6K*ؚ��H�	*d�l�n��g6� _�V�:7�{g"O��Q"Cl,��h,�Q�6�5���Dp�~2�~�)z��e�%�k��0�f@���<I �K=��@Q������_T�%���nv�5̭��'�E�@��J��WQ��35�ۖ?�g3�<mU�r�ח/J=����Ѕ��E�:�}� p>�+
�N�iĺ"	��l'���kW}W 2L��W�o���:QҘn?g<����R��Jm�Z ��g�9;n3��7�4̘�qc��ߜ9�0����v����(�Gzq�,��.Q�5�U�R���/��6�o���͆[q�#�f���|t�n,)"	�@��ݰ��`P'�)y����7d��!A�y�8�8	�e�?��	��t�����2�@�mP�]�o�&��m�Si��HZ��_��"N6����,(�%��]zh��I�u���c�m��؂�.�Ө�%����t:��d�'ކ���q:AT��x�s���F>����ldf�,�F&�����8I�ܮ�q��@ �eDR��X�#�%:@BDǑ�?E�=��\���KTcE�&��l4^���F �q}��+ۨv���a����h|�i�^����C��r9d�М$#�d����A�H9p��ilA� ��ʔ�������CnB|j�KƇ�`-2,_VS���F�Hj��E5��bC�K��sl�DA%��Rm׺灹��qp1�3F��dO܇D�kAOP�2����Ƌ�nHB#ִ��Nۙ
5%��'.Ng鐩+���$��Y��f��H�،o��p�ڢ��{�&���;���O&1��LQkH��Z0��v��P�I���]4�U�Hg�M>������o4���:����+os(�3�!���t�7�ѻЌ�
F�������}5iES�C `���R����~
oYK�ɾ�WW�G��s�q����?QCI���%���:)�q(�WO8���m.����ꮆ
[U�1]����,�$,*@�%��R�~Д.���-��P��'ڑ�u|]��O�B� *W�\p�i��زa���Z��IUT@.f�p-�uG�*�xY�x p���֦�"���^8���\�I-����ކգR���Oe�+���Uk���+i4��d.�݌�G+?�E=�,���3��LQ��x:V�߃bXI���5��4�Rl��
�p�J��w�g>I@�)Â�X)WГK��eON�����������Wwgx
������,R.��Y�(c�����ZleE3��2��o�0��b'��l��zw�.��'�O����0 r��@��z�����g���?���37Ѵ�8ư�=�cߢ+R�
ld^��z���0�M���k?x�K�A�� �+,��D葊�J��:�,�=K���[B� ��0A�0$o#{d'�܉� �7�7�p�c4���͞�H�'ÍP�S�����G{��yE��l Y�<lNh��������$���ɐ�N��}1M��2TAGE���^�p\�ʺ������o��}�t���%r�>�\X�L�cOɪ[!��h����059� ��5_������_W�%}�� ��5���JS����e&��T�z���E���]o�Y$���ѿ��e�������O&�î�j��W�աiU��ט�_R�v�