��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]fӗ|��"<+��s-�󤱋�#��,�$)��Wʛ���,��,�g\X!4B|	�9B��:O���)oT��9JeJۡ�X�m��1���c����Zn��_n���;@��e��Qy8�����x�G�W@;t���� �$��ݤo�����h��08A\�L��1��լ�&Q��k2�}G&�^!���-��l���tvU0VA֝�y��y�H����F�:5:R������ƹJlZr&�`ғuT�!@W���Foh��\.��1l{�����r��_Z��3OZ���P�~�ji+$�Yf���d���.\��S�sF�:2��(3R�L;b�����3?;	"g:'/��ͯ�O�N�c	���NF��9C�:���N�p��(i�N�-��z������ Ų�v��|e�3��pW�k�5,�����p<��z*��hr$;U��7�\Մ��;�@�.������ ������ ��si]{�9g�(�Kqԃ��1�%s+[![����VN��L䜗U�[��!EDgoǔCKR���q��u�����:O�KP|K�	��7��]��ܨ�[�I"9�����Na;nѷ:ȵȊq�Y�F��5�N�(����g5�Bfs�n���Y`G��k�oU�1������\Uu��}�;~ 8~����J� o��C}f���w/ќ�\�r=sW�죒)t���� ,���#�����#��N4[͒��)���s:鵏�f/G�����o5��-&0��uh�(��E�^^�0��N̓�:%3�|9VN�d.��\�4��il&�P����nڧG��mr�u7�u�3��lć��� ��G3oD��Z��/6�rNu0����fݯ0^2�����?6�@'�l�oX��B���[ְ�R{,��G2����7{��W�YB>Zg➥��K?���߄��K�/��<�h�&^&$�_��n%�K��C<�WN�x�a����-�U���/�r��ٱ/�r��gua���J�M�M��\����,:�i�%�w�j0$L��fkw����X�Ep��J�S&�=ГZY�C1o�h�5�^H�4de6sJ*�u�>֣ܴ�����8�]8]�G,㟝�����I3���)D=W�܆%A��XE���s�@�f�`� �"<�
�������n�pg��MIRvD��j�r��\gU