��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħa�gU�]@)},����ע�����0v��D��CI���O?\�ܜ�0��cc�y9�į.E�'��}� 	���iG��	�c�7�]��^��V�@w^��R��7Lх�a,��=�Q"�̴Y�%c�����7j*u���L
�
�G�����g4.�6��5BYSd�1�#Ɏ�\�ֳ��8�gl&�;֡��=A�4�I���?���K��:��,rM���Җ�Կc������{��۹�{�17��~�ɫ#w�O�}�&���_��u����P����Еk�1�,&�]�j�P'�{�%� ��V��5G?����Bb���l|`L�A���;��1R�jTl��S
w=����fA�dj���ȃc���"7)oW�& fs6�MR3͖�U��<ͧ7��w ��"��E�
�S0�4O��ь�'f�����׭g�~��{�+Y�5�-.�)������{:'o�`,Y��<��l�AB��t\�<oQE���0ɤu�䧁Z�_��_�L`��b�O!���ڌ��
�ڍE�;��I��u����*�CJF��*q�9��~*PF�5{�&�\HT���#�d��z�9s�8`WU	�7?�q�,VC>�������).c�=�����J��Xn�TOɄ��L���7�C��%b�RF];T|j������c���F0�1�حR@K�&cvKɠ2R��n;V���3�G�$\��.Q�˰�[>nBX㡸P����kYR#�E1;F��S�x��!%����?�\������)C
2c�2˯����o�0�&�q�bz��ؼ}wi�7����rԑ�%P�uA���p�Ɯ����@�)L]I'�i����?����`c��8;��,�p�.WJ��jo�� ��Db\>M� �����{¯��9�<,ӻ��G�����.��$�T��W5
��
acCٙ]*�1��W�44�.g0�X+s���"I���5en> sS���վ��)�\�.�t�-ׂP�s�)]́^g��R]`�w5O �k+��e,M�eEj���P]ǲz�2zw�mv������j
�O)Ov����.�TFk��	Z3�
y҆�H���	��c`h欺vо��C�M!Ք�֒�l���#A~nߝ�E�`�?�w���}#�����Re6�����y����P��^H0�SB�<��1��L�� ��j�9%�/+ǚ��R�I����FF]J��.����ԾO�Q8d�_�,��=l/�S"�aEH��QWE����	}��r�=��d�8��PBqJ�h���<Us����I��ׁP�!�hŁ3Fc3�hb�)��>T�_�vH1���qbĪ9� ��V�xL�=�}`�j˗-�t�j.��	�{sh*����3�`����ݶ_^5jA$���.[v���?#.�l�pER�� R��D��A���x�)����������edY��>!�w���x��a.�@�8��e�뇇�*H��9�slPt����o��/M�yҐN����.b-��7�kH�^q�K����W$էf�A�� a	�ᄈnd+2[M��b�?hC���{�d��Yw$g���� tԑ�C'M�|ƝuEm0��qE���"���5�oü�h*:y����`�:���,|�iP\N� TO�m�h��V<E��?�W�}z-eT]\�{����4l���$����h`s���d��>4�e���F����w_�-�$6��i�ZP�q0m[���k.�?c����������@o�]r���.Q���!�6u�����i{kw�.����6�<y���'h0[�w�ybI�I�7�˝��|�H�;���>%nʧ��O�2ۉ \vqq⡅mϟ���y51��3�3���`J ���
&Y��K���e���4�7�|�O�}���>m�����R�'���F���A>[s�Uƀ�3�����Qk����˝ ��$/�RT��I.>����* �uC̔��_
X^x$��Ec�@]Q�ԓ��{� ������'��	��'���M)��1�<���e�|� ��W�T'�������<H����7�-�	�<�����t����"�?[�=��,�Ĭ�D�5��.�O+��2�Ӹ|c�c��U'��Bc4�n}�]�&�:|`I2NSg�c?[X�) �W� Z�٦ߎ�|����A��o��A��Y���
��~}JV��m|Ɍr��4�J7�:�L�F�9Q�bfA�[}�\S(Fj�j�^�64��V
�Gk$�4��DӾ�(��ޛG�҈�V��W\I��d9��a^?��Ĵ� `B��㶼� ��T�Ys}(V6�����{C�ɨK��rⲐmő��.dcҒ��r�&���.H�j����x�Β��9j��A3��/��p���=�	@8\w�KD�[���OP����һ��%%�!���x�������-|���?�h�Q�
��,�"�fm��5��5&b�o��r.�O���p����f��P��R����"�1�3��#���Fi20��)����H�Ad�J�7�F�%�$v`,9���ngk�e���+�[3EV;륩����	��v|Db!��FIa��4f ���sD�������j`��zݎ�/x�Ȧ���͖���fD�X3�ZB#��y%���r$o����I��P����a�ߘ-5�B}o�B���	����f1�o^-[�c�6q�a7�Xgn�+D!�& �R[��r��&ѻ�A�wR 1�wY�6�3-�P2��	��~|c4[m3����c�~'�����o�XB5��&�ߢSA���a^$5ڬ�ltf���{�$�����2'W��H��++�.)�D57%��bH1\���['p6�o1�4ŝo ����i�N�'�� ^��w�,eq���x+�QM7���<?���뤖J.\.�=��;���q�y�~��v����am�t~�<��D�)b0M�$$b/l�A��qċ�D�lm"t�{�T�	�M/���>�K��.�Fh+����5i��pƗX��Ty���E� ހ:�;�>f��v�#�8.ߋEd`�*,x�V#�g0��2bO�1��EB\�
�MF�ؔ�rکN�M�p&��GV�8+E�=�b��>��=W�kN#Lb�lf-�"�geK��ͻKe�$\"w+u���E�m1{�r���I�2��' ��<�?j1b����h
W?@���&��;c��14���iz0��^�e��!Cu�S�ۨB��W:��Yq�Ȏ�O:Dv��CD�#�|����
��^�EO 	�͏q� 
Z�|�wMV>���-�Τh�Yo(���Ai�&���N�)���v��9G]��!P���C���\�M#җ��+��M?�8s�I2;��b;i��'��n_K�^N\��Y�ta�l���B�Ÿ=�$��Icdm������B·&H�Ow��Q�Д�=��|�#0�_��$����r���d[�3UD�����GT7_Q�M�ˌ��BJ#�>D�WG��%�T	���Қ��̽@�ۣ;���>t[�ù�鬒��;��!�:ӿ&[�����YN"�l�#+��[��s���s�y\�37xFy�6��4^n����58Ѱ[�^�|z}�L��7:Z��ʖ�oX>�Ʀ���п��I�xVz��ڰ�����CT5������2]�1���"�o�k��\sL"�XvA���9�]�<Q�W��� ���qgO��+k�ep�Tʀɥ}e ����?��F��^6��X��%y |�22k5�\������H*:"�����ˣzf�D`6�1X��_�������C�&�౭Xm{�d:J�cuڡ�/��CN���/b{�	�����_SX��b����Ȅ���Z.�\r^���ĖxE� d�L��>1;���0h��5-ew�����IP���z�۴d�����EJ�̙��"S3R�	oD��t-Zo�آx�\Mݿ+?5>���4�u���-b�M��7'Y2S�{��\Aژ� M�B0��G�L�(E�1O͘�	�D$��.����A`J���T���� �}�Q|dl�'��d�).�.:t�'��3M���`�@؁�m>�הw)۝XS�	(�S�e��3lz�^[:Gb�Y���7���v7��Ň9�xr	����\�`%#���B~_|>����N��@�Ǿ@,��e�-'.wH�Ċ7D�YI#�˦���|�kAZ��Gvf�R����|#�pj�����j���V����z�I��,�4����f�­S�S鄜#JDC� �rYIV��8�'��l����O[}b)&��`��L�~@���YR�U!yP�/�sK6Iq��C�>ă�̿��wYbB>�G>�}��)�߲XM�u��?)��p�=�Z$y[��XM�f
'�������e����A�_Â"�LA��(�k�8�H^wA�VR�{���Ԕ�����P��8���k3�V	��N��:��o��1�S0R�>��U'0��E{�q�Dف�mb�їGH�n�a(]�rf�ğ�ʽC��vj��1�I�LDR`�p۱��y� �z5�@Lߍ"e��
�ۯ�+3`R��R� �7�	�]���p�w�$=���i�(�e�fR(�c�JY��+,>�: �JO�,����J�h@G/� �v<�HV[���b�
�����_q�p@�9�����kbGN[�Ջ�DM@���>���5\�RG6E�[���t�m*�Qs-��$��d.n��}����Wz/��&&r>����
��������A�t)�c�^X@�\���~���{mb�c�{����/��p��H��3MmK5V+�Ǣ5����s������]+��C�q�����^�*�#jf��]j�I��g�!t�)9:�78k��$f!Խֈ�L'� G�7�5vA�¦�
-�]_&�p����u�;1>�о&�����<6~��N���󥀦R>�/�o������l���~^����V�NO�����d.b����u*j��û��a��XҞ��o��w�O��g�NM��f����o�����P)�#!n!����C�k�23f*>�~7^�\{$cW�Q�J�� � �>�G����g|�����c��/�i�z�m��纍�v�=KA��4���b(p�<�l����$ЇZ�kdK��Ea��(Y���佊fSj"d�֞��i�22�������!hw#j�v;O[��C��W.57�CN�+��R��ԯ8�E�D ��4�O�k����cd-4�1++���>K�K��6��`�x��UȬ!�{	��e�s�	��I��|IpmI%�)KīRg�~�R7n+O�nAӣuN�� �K����=Fu��S-I^'�7��c�F�mK*�U�M�_4�Џ�1��wW*��
�y���H�,� wuN%V�&|�(�6�]��wIo�i�L��?wc�/��c���+p�����7o��\Qy�}B �alU�����Kꉦ���� q{C4�G�\��~�� :�ݛ;�b�G�A��y�瓆��o����u����F�<�%�'D��a V
�sX�d�МЭ���\���C��I'Qs<��5+��(�>}F�vk��ʁՊ3�qg�v�^���Z�16��eG��&������켌͂����p�)��6Sl�ilt�f��A}���r *���<{��pgJ�#���&��l���	Č����e
�]?,�[�1��T�3�c��mRԁ���p|�|kC�OĎ��������MN��w�E+��@�&dŠ�@'I-��ȗvl�~#V�J�v�N�{�r!>�t�F�>Y�ʊ0��=�C������^�X@i����"��*r ��!�JTgcJ�ğ���g/���{ ��/�1 ��&w"Hm����}7��`�6d[Yӆ���?H�@��X�/�2oz0ca��og!����Ý�(#��%����N�h��B"�,}�*�۞D7ڹ[� ��%d�ZY��|h3q�}-�O��i��UIMh��`���R2�wUPZ��?��_l28�p�b@x}�tnI�	�ZY���Mn�$�5*pAdU}%�:±O=�(��hR/XQ����Y�9ǚ{~)�U�	�Î�كi����CYsa�<���@���db%�
s����]!i�������QI/1�5i>����rU�=�M�ZvJ͕4��bdZ�sog������y�<������1$��Nl��ȅ�9� yD����W]ҍz��F��WT�����'�I�!����6h�ė&���<Jo���(S����� 6Yz\e�H��A����v�Я���M�@���]E1�L� �@��o>�31��t	����s,�0�����Q�*#��5��v���OJD��"�mD���k�{=C���̻;�x����TJW��W��^����"���|7�������@]%c���
��>?e���S
��D���5Ҝu�[Wy�50�Z|(oW�9��C=7�V#��	�$5pIJ���e鶉��6�B�yT�ul��!���T0��2�_�,j��|cӯf5��8���xr:�u�$���v��?v.o'`�%#x����D�`��3G��Ӓ��:���M��30 W翏�z���Lo ��/����r�C��ؽP%7��T�5 {<< ���.��[i#�+>4��W�H_������B�wa�SR��yC=C�pnAmf{v��%���6x�w��b}�!��i�Mm�B�0�{��ԅ��業S87q����t,²*�Ze�;˨p��O��Ӄ�_��!���;�����h�h�t��tŢ���zu�>D��x=��h�0�Aw��f��w�Ib���(a)��O��Ǳ��y�k�BK��Qk�Z�c�SI��7���?=�a+\�`g*�}����cLϏ-�GI���E��cZ��6F�c�����B[�}�/�����F����5��Ω2�M)w �`�@������h�i
��Ջ1�� 
��^��<�c'�e������!�m��<�CJR5Y���i�EQ��0�t��zƭV��eů->�sAxo2�n?�Jo���{���*�`f��І���b��N]J��)��7ԣ��p�3�x�U��;�Z����ہ$���%#�,z��$�O/@�K���\+���"�;�$
�$��2��T����	�{
�L�5�ë�w｀� �N�o���#h���4��]�]��g�}������d�9���4W@��l���=hs����tb�eB�w,�X��:w+��}J�i�=�Oֶٮ��o6mp9��� V�>�Dm2���-������MeO�\l?�����a��?�W���8t�iz�?+L)�k��4��W��uF'�e���R�vUǠ�b�x�S��+�ڨ��<
�D�L��C5~��un�M_Q$ju�3^���[�8���Z���^�'�p�<���Dۆ{P��$����X;��Ȱ�.%�u��T�s�]�6ȪD�s`�gM��ĳ#�/����{�(ѻ��X��+�-ٯ�&��u�<ը�ȋ��`������^�qm��v����~��\���P��Ipȡ�	(���M>���I��5�h�+s'�Q<���>�۝%���N�$hԿ�cO�? A@�L��Ԙ}��INߙh��g?T�g��b�����)��l��V�oY�_������ 9�A>�qd��u;��Ȋ�'35[r�~��FF/�&��z�#��BNF��/{G��������=���(��1�kX�D;v?%�|�T���r��S4��k�R��u��'׵�HOp���Ǥkw��V�M�{�y~�b �%>d��m�"]���%Z�l-}�q��<������-Q���8�,�a)��U�q�R�dn���[��o{�H�Q�Ykc��Ƅ������]��/�Q�8[��,��D�8
Z�I��z��IRu���x�������%����D,[af�&�3����"�)>��f(�n�NJ~Y�g��p��O���'#�~n˙?f�
\��������{�ꐚ;�ï\
�O���w�&y.h�?�j��ȑ$ϡ�U�iq�E"	`k�����Wz	�A'�{��!>��h�3&��Γr�s�B�W�g���8�������*̕\�hTt)Tta�
]��dψ �[���>!2$r��ĉ��O�14�u�Ax����G��IA�S|��#nuh���ds*�K��m!�$W���a:#��/�ݔ\{-FJE��������:u̸���|3�3�?v�%�����v���7�*Z�����إ�˳�{���S����-~��+U���>�ן�-��o�q��� �s�Є�&o�F#��x��и��-���Ժ�t��/�I���b��J� �A/���^ 2�N�z�[E���/�(RM\w/>�pH���cҪ8U.bIH	��K�bLy(.U�ˆ֪��� �Pb�%[��|��&;���1ka�4.u^3��3���n�w�8�JB,��	��l]^�3�~���q������kTa{��V����|!f���j����C��4T���u`��}��&�|��Y��ec���ej�a�q�5�ס��r���{�b����G��~60kq�D��U��'���wW��^����<#����zY�)F����A d�Fr�3I܀n��2�R6��<(��Ig���*(��`��|�<�U�t��CW;�T�bNĂF�ΰp1[	ؔ�I�8�RB�q��̈%+o8fk#�/�iV��o�3���l}T��`�l�Dhj�'�Qd�yn����h�W@(�� 1k�r���R]�R�}�g�y�u	BE<����@zz7���Mu2��o^�dj�T�޸��۷�x�a6��^V��hp
1%cPy�{���q��
�}�����6��P�$s�[�`�ٍW
pv��6�b=o���0)�AES���$�����B��l���<]u� ��w��i|�-bN:�20��mJ99|+l�o�=�"�9�L� �`n8d w�[���BB�\
�ȍ?ELH,2ܡ:�#
�u��J����h�܃i���?�~�tJ6�Oo0��-~���$&"�_BC�q�ޛ��H�&Oib-O�́�^��{���.��Ʊݴ3��8+�u�ؙ̢�"o�ϝI3�[֞YC���;�H���5u�p������j}�wݚ�H�  �~�/}́p�\���ݼ�m�6K� ξ�ڎG�8�H�a�Q�����J�۾*< �	w��^��ⓉiE�ALrJ2)������Ϣ�IG�ϫy"�Mڣ�4bU���J,e&����S{��e����F�c�v����94�7���m�v�+�Ӟ?��G
��'a�H�E�_���+�Q�v
_�+r�]�"^y�����B�(��斠���w��q<�G\�H1�Q�+7��'�>^�� ���$JD׈r�����Ȣ��nv�O��'*�\2�l�bH,�Vϗt3��عu���@܌6�3pz���i9���!>`����=ʺ�^c|���Q��-�ä;�r��%E���@\���Z��NpS����#�����Mȵ����<e����*����w�n><A
�A��#�ș*=�	�mG����+�9�CK�*zʀ�O�Yl:�]�?�1�}]��;ٛ.�I�����2�\�^-��l�*�~������`��t�t>Ȉ�M�f�twx�/[p��&�����I��S�#֑u�;9S�F�m�T,q��_�|��ߦ� �\�E�ns.ax(D�