��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7Ɋx�!�g���I'k�c�Jӳ�xz�:�-94Q�߼<p�bj��vC7$=��ȭ�B�z��'4��PNG���Z�*k}�&����G��.�}Nw\�{l<����fd�qf�u ]�[,�/�>Fm�EUx��`�
n�
\��WFO��KwL�9�P�.�- ց���u���$ |�ɏ��$B��W���aZf���b/�@k]T�H%��?���l��O��G�5R��L�]r?.�<��~b@����*R�vp�͉�d���rj�E���A:��P~9u�N�}���6Z�p��%��d�v7r_'^�]u�f�e�dδj�/����o�>di ��N=��l�P�r0���^Y w��EZ�(��'�l�#�F4;����	�I�৷
[o{�}U� �K$1��{o30.u'J��Y�<MX��!����L�?�
'���U��j��t���qO�dNT��l�~(zi�^��~�"rq�r�����w�Ζbr'����$#%DS85l�X{\�5�l%��Bn�+��yt���ɒk�2=��V��
�:�H�fp�!25��������ϧ'wh�b��(K�Ja�=Ӷ�#)=N�bg��~D:o�����.�3S����B1�����O����!e��L�J��[(��P�5�h/���p�.�L��{|�ٚ�w�x�o�$�0qnZAO�st�8�éF��!i��{!igq�����ed��c��Ϧ�\V����;��N����9�OgE�Q�Q&F�vE�`��>���2���-��G��Lf��M��w!*?J?u��,�QW�U�����-O�v����^Q�!�����ƹ5�� �s4W��Qyr!$�cH�����HS�)%bH*�S��֡9Y���������X��³�!y���ˈ�_&^�	,S� T�To:25xǄ�,�U�7�<B �};�K%�5�����O�e��џ��0��g�C~y��m����1��]�ڛ�&�fl��|�I��ãz*L����Ol6�㱁�.�[�/�_�� �@��XHPt����֧��D�l9�9z[�4x�i��sf�.��{���u���\^T�·��W��:XI�a�˫�	Rwì��P�����j�,�^TSE���f�h�y�oufxn�8��:g�t�,9�(�^bK�#
���DІ
�b+�Fкb��5b�%l��,a�
 �|]��C+]�h�� v���aI�y���&6���H6�X���D��u�ǎ9��|�@�ME�g��A5h-^��}�<be�
1t�Eѥ�����g����i�d��*�1N�e��NɅ�U_���%��/s�� �77����Ţ_��)l?j����Έ�0�6l�>���,���	�?�a<��wN�	�ʢ�h�-Ȁ�+�Ƣ�eJ�d4P�H�d�OTܮ��$��_�~�Rc�ꬦhS�*QYe�_t���A<ޘn��]G�
R��*^$ǃ
�ȅ���-S��
,-��N�^oU+Y��GL��!)�=:j;RHy�IgԪ����5}��H|r����J#��������cdiCt(��r1�	�S�)l�@���2���d�<�Q�@M����%��Ƥ�{�W�ϳ5�r!t�/���E¿��*���p50qɇEL+�ɫ6<���a:��֐�����&yB���v%����Қ�_���BL}���1�9}�CԳS^x{���L{+��k`p�Ih��:)�0/xp��|�3�]!h��%�����,�;H��Ž;.�=��ʃ�;*puy<���Z:�q2������&��z��h9:�-��?㖠���qd*X+�$ǁ��z�>�|'f��҃lv��&��'���{�H�D��"[�EB�"���zg4���SY�X�^�'��%e�Y����'A�:�@�{�()�y����CX�� . �l���ܩ� �����f�'�U��qY��P�7��xB�Uex�ڨOw;]�gF�ΰ���+]?"�+r����<�� Z�0P�E��&j��zΤ�����@z��֨8\2�3��0��v}�]�[մ��_:M�'�Wa��pS��0l'5�W�7�Z�d�`�[���Rp_�j������9	�ʈ\3�ܡ��DSᔷX��5|s~ �g�Vf+�c�� ��=�:ld�lk���G��û�=�}��Q��qN����a^�PS���(�#A�4�� L�D.�,;U��g�_�.m�Np�x��7]����|�M�Y�/�s*�oDb�wb}(��fS�d�Dt�ޒ���&<:�>�粩m��?S����ˈ?�hpD�H��{��	Xo�B� �����&U�����F�Y� �{o�ʽ�?�K��́������"a+,<�������ҷ�|��B���8��=�)�Α�t�}�.���� 2|��O�	ќ|�ZƤ}�	��gjA2�����椅R��/,��C�*J�mwĹ���[�c�D����K�.����g�	#�%�!�\<�_qd�!s��M�*57�ܸ�8�u~��\���^�ŝ���vzM�M�&�n%~�B��r5?y�0��7<0�:�H_c�j���d����W��DA@��kk%�~/	�aT�i�U�I��(3^o�z��#`��ZSg��>�'@�ť���Ё�X��R��ƚp`/��X	���p���, fgrA6Fk��ӛ��s+��Ɂ���Qj�u*}v�A:Ck\���w�����mDP�A� Édt��t�ê�����}z��2�>�������Zj�a�;�D+�4�?	%���f�4Xfko��w�l߲���$����9<�#j� ���.�G�S���H��9c�E���؋Z� �6Gf��j��A��Qx�Q$��:�ld]q-N"��"�ft�N�`#�����m���6�?yL����j�lr�����a�ݚ��%�zŧ�������А��=�.����g�g�=K��:Y�Q���p*���P���l��=`04D2�w]�Cx�����b�����ކ_U[���T�q䀣O[AW��CSmOj;�������T����T�.�I���$Y"٬�� ���
�bk� �˕++֐�L�N��xž�J���!735�4�M[�d�j\��{o��V7 P�},��PRI�:<DP��Q����3��5���Rl� \�w4>�=�����_�˝{W"��AGHhtg�f�{G�'�d7C: �
�̍Al��h	����˃����I΍5�������B��@����
"8�#˗͢5%a�C,_���y8��~�q4�9ܓ�$�Ჺ���@A 0��ߪFA @�k8�r<��𸪶�$��{�J8��-*:��O �"�}\�I0�B�J~,3!gJۨ��(��>Pނ_:�m�hW��$�����r�Z��d�6v�	�p������-E�ׯ�oϱg������ۤ@�v�B�T[���\�ѥ6F�芲?Z��,ڟ�/��;w����n�E��g��ٲ�#�\8��q�v=26kP��}R)�_y�p0��R�2G����/},&C�s�����}�#��O7݄�Ք/��X.2�(���+���6��K�Y��2�o�2�j���Q;`H(���K7i�h�9ϔ��4�ty�]���-{��2��5�f��c�@��-�Q!�Ǡ�I�Q��6(�:Z���Ä*	[�@F��\������"N��zۅ�q���`�e���x����� ���ґ$�F��E���@q��\�6y�$+C��9�:�2�a�A"9���/φ�aoӮyt#���)Wl��ը��'�ɜ��疇��i��#�?�J4I��Fm,
8
��a'}�h��G���1^���įv��z�Aw�[���ƀ��h%}���P�7�b�hD���H�B;6��I{��;��x�3[�H�%D�������f��S��G���&�7��BẄZ@�U#+yhЩ����Tu����g��}��A3����?"Dv�þ�4�3Sc;�����k�s��Ćg)z� E>�Ě��hE]��Uǩ��,/���Nf82�2x�&At�Vc���/��:)��D�1/X_&<7�q��Y��w�)���THI!V�|F��s�*@��R�	�.w"��4̋���V��x�x1�\_\��<��K�Ma+|�7MuA��Es����,|?�m|���- �9�K���zp�+IޞU�M`^�i��<���T;��@O�
\�:�x���x�[���5����J����>�q�cbp�T�xgZp)��6����q�`c�5U�"@@�rP�kw������%�,�8��e��۝�<&�<��5�)��)-BuH�z��_f�����oq#��N�	�I�5hI{fV���	�d	h���n<��3d^��S�R1�V���rx�9�_8�U�͜Yf�L���O���oM��D�y�o��碛:z(�MCHV�2��M�.����r|� 2�P�K�[��X;�28d����I4(�����oG3YQaOϸ�M�9�o���K����	�>�4u;�	�j�	$��z�0I,��`��qH�}�����K��r�zN�KI�Y?	ל@�o��Yl}"c8T��5��'�����
T��Y4s}g-z�Hi]�e���0�j%ƬHms> �;
&�����Q?i��G���@�1�U3iv�2	kWj2�F��cvI�s�d��Fb���~ݐ��_��u�Z0�����U`Z.��JY���j���<1۪MW���?����^`������0ө�,�!/^���$���-|��z�Mp;1����v�Pg��"��dz=<���|쏽�f�n�@|tf�:$-9Z��Q�Y�kf�.Cۺ�![�լ�X��in<���챃�����~.�!-%�E�7�1 �����sUp���
zt�)����!i�+9��F���=~�wVJ�TN�Z�.��S澐�kw�A��q��`���Y)�I�An\COg�ˌr),x��,[�8����`<a@i��%��9XW3�֦bE.C�}s�|�a̦o3M��e�>�-�pOt���絈xh��(�N2�ܼ~�/�Ι�V9�˱�Q�@�I@��CXI�Il��6?i�;_�b=�5�S�U&��G|���Gy�fΒ5�B�0y,�º�Y�wx�}A���s&*����1�v�&Mkߧ��AQ��/���W�o��zG╂|t%��h!~���Qd��F*�Y���P��2���h=-x�Qq�$��cZ>`��5�w��������!4���j�q�Bٸ�;��_  �.H�.HJ��~o�<$c��^�)�"�@q9���O`���5�j�mƃG�sQ�>G	r��Yj�YK4�P^?�+,��j� &0�r�4,����B�w����0j4`�琩7��S��y�se^C���t���~j�,#b��O|�р��^�n]O��a@-��a����OiJaO��QU#������z]���5���xGe�$���WOlY�|�iM ���i=yq"s�*���7�(�K����;z�E_�;{�uH�T�5��
��FY���Qzo�»!j����w��25���u�]���" ��s�8+~G�����N�h�����cGK@�2��:|�]T���+�iI(<��a�|!f�s-Q�)q�r�������P���ڬ9�����ji��s��,���7f �����3OʽM��a�\�˥��D�E(�4P=���U�a�PiA�<|R���;�5���yځ�u�\6xY�̎����F��͡o�HF�WVezG�Wkr夋��[��>m��ƹ�v+�9��a�#��ѓ����a�	��JUm��L���Fb]�ā8�ت_���7������I�r6s�j���-���Ȓ�5�T?���B��"��&�*�蹨Eࣗ�v��.AG�2�a�qi\N?�J�+�P9M��å_�y��9ӿ���P���t�x	�IX� 0hoͩ���p���{a��՜W�*�F� {I�A'8��n}���Qc�J��]�J"�4��GT����&��}��FN��^�*<ù(�)���2K�XW��~��Jᐓ����p9CH�ΣY�C�W���As,�v����˯���z=��Ǔ������CW�(�m����0�?h
��	��da��B�qs���V�2AP�f� t�#I�C��Ԉ� �#ƃ�E\�/0�_g��H��6���<B}��@C�f�%@�<c�(ɫ^Y ����Ia4�s�B��&�ab�	��Y�j�L�l`O�ݛɴ��{��^3�r� 9�a�Y��X��)\W�Q��e�dt�6���ȇ[�-�7Ӫ)/M�MbDR=_�_�5a�>9��e�ٮ$]��}�>���((�����{UH�ʯ��̒���U/f�6�"
����>>���Ԅ�K���.�����򦯚m�j4�y���ڥb۲$\~kGr��7S��=0Y\�1-��	���8�ֻE]�E]K瞭c��%Z?
�a����{<�N�x�x�g>bUcl3�v��{�h��[�^-O+�����d�W|T4i^�MP��)�5��5*�`�f	��-���a)����\�A���
���:�X�e�K�c3F�KJ�ǌ�o�G�yI�̏�n *�2��z�d�r�aQ4��%��*���CmU����z��>vذL���T�[H�;KS����0���6pn��W�Ŕ�!P�p3���=�����aN\�\�Ӭ��_
�ȎP��(&ĶI�jgM$�j��>�}V�c�^W����L:p�J��V.��r�w��*7!`u����x�i 0Q?�e��u�S"l]��R�З�_+�b��8ɓ�>_#q��+���� �`&z�e�y>
Θ*gf'S����.���H��[]��1����}�5�	�2(�!
X@�7��En � K������5��cwZ����O#�Y�"��c�K&`~�*��<������Ōе�]k޲^[Y��߹�'-�=��Ǒ�z�_�ݫ$2��3۟MG%�;u��hǸVK��,�L	k�ay�}��J�t4 x�L1?�v~�F�	�������.m"���ƶes�~��]�	lI.2S��$V>�66�V+�J�B���ϣ�RK�<���ҋ�>?�e�i�!u�B��-�d��Z,բ�G�S�b=��v��������`�,ό�S��)�f�f'�� �TzP���SF�n�����n��ٍ�a���y?��\��U6i���q̛�V��q�r|<b�#�����M`�|���fK}oDd������#QU�\x���%EE�3�?:�r����}���h�h������l�Qƭ�LvP�]���Wy��(M�ґ���X�6D�bz��k3<�y���1�Ʒ3@���PB7�u4$v�m�B��#�Jr��1�=���j�G�ŕ�B� l�ښ<�q�;��&rh�+$^�A݈�{b�'Ӫ((E��ПmMp��%���p�/P�j<���7�*1��l�S��O�J���ӧ(9~?�Rh�l�MQ-8ݬ�Q�:�2ou��7y�U��m�9�$!A_���6�A7#� !�''��\�u%�k��5 �djKҁ�o9�2�C+�YVƑ��x��ߓk_DYL̯!Y'y�?��k��Z	���!��\�DT���J,CT��ʟ$F�eI��D��:�a|�ݽ#0�u۴ ��;����O6Y���ٓ�j�|��y�K@�����:���	�����tЛ��D�F�+�dG��m{������Z�B���㛰�P�m5m&��'-��W�)��Sh�9+^�ѧ�@|��*6��w����\j�yZ{�biCj��Nǐc�%���c��ǉ�E��w��!�hO��ƙ&��X��)2�I1��u����+Ɏn���j���|¿Noe�;�Ν�V��oZ;�����������&�-�_�`��_Z(*�),د,��!�q*Xw�e�3�,�=�����c��%=#�?�I5��7�F�����'-v�R�ۉ,tF�>|�z��jb&h���$`�^���Ω��tzTS�կ��XrŰ�<�7I /�Ƶ�ԁC~ -�~�^LFL��]��q�8��Z	�^ɕ$�ymO�1�K����5�� %c��^�,�z1~&�� ��C�MMr�4�ُ��j�z��S��(C��:���`�Q�3�'J�����X�f�n��_�����s�؝$.�����N
T��W`'9"����+���rO+Yq΅��@L���M�n#��W�<(X[:Zסb-\9�h��7`b�崩2r�I5���y��L����}�7.j�#��^�a��*���~�^�z���'{��Qتv��c*�C+��X�G3$ �$�fJU��su���*S;�������+�W}�w��ν���>uo�Dd��b�JԦ
��#��OQ��L�wsi�}�O��Q��Ѭ�ߔ:��<i�A]N�D����j�rx�����k��&S;��DI��� ���`�����B9;-D������8X<V�MUy֊^�[d�`J�M�ɕ�(���ًR�M�,�%%��\����*TXpy��.��K	��hF:�G"(�a��ӸUq������v�zg/�}�D$.�)̇�������f:M��`�-%*x��7��hr<7�M,�b:�h/t�ZҚ-��ڥ;���o�7+ԅ��d�=D���� ��ĚEn!��@���^�O�v(�e9E-��W�ʚ�<��1��[�(��j�+���˙Q��Q�� FP�u<���D�� ��K���@v�d(1�"!.~�����
�}0�;�{x|��[y>�r.�+k�~���H��|H��H�1��9���S�&�O��Ca�^��=��	���Fu+)��Y��]��y$+� ���xP?�-ƭ���.��:4��;��J"���
 ��:E���b̯�a�T��?�D�8�ʘ�llL��f��ϵAb�roQ͚�"@9򮒡�i=��aG�#<8����^��.�K�֑6��PԆ�m�c���Z�7R��9�M�09c�_��A�G��z�hrߝ�|lz�<7������C*��xhz����dV�a\T�U4�7��Mlv��28k�K4��޳\�qZ,jx}��#��.,RK-H'�cK<@�]}qQ��x�z4�?������Ғ]g}IW�7j���?�Sњk�5����<�՜>��WC����Ǔ���aI� BOT�-�7+i��)��I��fcQ���͸[��n�}��'����Jt���ba���R9_0�1�E�>��$�Ժ,OwpQ���$��_��ee�q����īOܼخ�W�Aa:���m���9E��Y/��:�#��9�я%�Q+6r�GR���By8d�S�_k�C%
ѽp
Nb�L��t�f��ʄ�6��&�Br ��!~�E5%NW����,[HN�5h;�F��d����QKں��G�A'X͔���(�4�s�o�{��?����ҬqiQ�\���oP�H4��b)���"��X��2�pr����O:Z-�6VR�rT.��v},�<V�������u38���Ғ�*E�/#�@�(A��w㨗F�I��-<�8f��9ե`XoV�i�n��%;��rc8�c?��6��� %q�7~�S�
�,�b�'��k�k�*�d 3���D��	�p>��y���m
t�J�'�`@�cy��� j!]e�R](���|)�54CSN[9G�bw`�vO�]3�:%�4�+Y���,
�;4�r��	��b���!{.2yd�H"θ� j4����C�U*K�6u�:qDS7~��u}Cca�qvu��6�6t�J���=�>�>wY� o6_v{�u}�@���X�fz����=G��P��s�Ko�z�4��h�IL��3\�3XyH@�c�r�G�K���K�j���g3�,"a���,���2��������8�!�҉n`\_�Y	�~"���Jg`%��R�$���O�qU%�yXN*��٭�/��[�#C��_��o�ӓu?&PPd�p�R��!K�NX��׽[�R�G��N�ϢD�97����P�~��G>�*r����85�r-�j4֎B�:>����B�2��9��e�c����2K�kV^U$Q>� ��X��@:������_�Stv�����p���-d��#��)W��:{{B*�[m�[YTc������B�q�較 ����r��M�c�+)_��S�,��4w�v�mې��$d0w�����fx�3��؁T��U0؊�>�P��β��&�n��j��)��Qd�⸛xw��گ�Ay'�R�oR�k4��cTO�*���ư�V�����s'_׎��!��iµ��x�c��^Ɏ�1yv��"��3.1X-Yˣ]p�b�r>�Ș`�E�H��Zӷ|A�!Zӳi.	��{��-a�����C����GP���f]���~�Ɔu%�dE�	r7�F*��:$7l
�$�Ch���L&j*G>[#ܬh�	����}c<�k�R�@zފ�r�N|pN���nd��ò�d�6Q���M��}�v��v�	�g�7��K\�܃{h7�d��ȁ_ g;���\��z�M�tZ�-1� �A�C�Gh�3}��7$��v(�ˁ�c���uo��6f���Ûo����K����8�"T��ҡ����BH���V�?�����n�`=l��Zy4�g�26i�&����<�y��'^���9��y�j��`%���7 �z�]]��3�Oz��	�M`4K��;#����I5_�W��4�`��f@�۠�k�B¦�ff�.N;%���Wۣ0��tMe�8���\���U<�L�Dm1u���mK�u��u�L4G�q�該S�(c�U/DmD�4h��� ��(Geۣ�V36e������sw����)ԢG ���锷�Ƒ��VuЇb�p��K���7`�L�A2�>��:H~����SW	�T�6/��՚f��
��%��L����=Ck(_�1`����O:Ƌ��	�Ͻ���=��0��4�_�dO���l0�a�^�����m��wgCP�^Do_�u�$���,|��/�2���(����Lm�|Z�ț�&J�[V׫tì�j��E����ȯ f ,Tj����T����g�a�,�M9S}�jMrq�}�,!��² ��Ţ
G�R�mFB�%.�rtӰS}�B -�A�6'3�[=cf��N��T���;�Q� ����j�
8GA��bQw���Q8Fs���h��g��@)o�����e����w��V=VA��1�"�;m�
)͠���Z�1��pnc�����B�Ѣ��o���q0��U�p�/��CyIQ[�6vV�ܗ�4v�!�W/�/<�g�0�3d�`Q0�)��fpq�STF��h��1��xR���$�o����4㣪��$x��T��;+ߏw� Ҡ7�bt�z�D�/A/���1xس���IahZKt��9X'm`ifkօ��vkfs��PID�$���FzZ�ږq�����A�@n��2���ܟ�Ć�qN�t���'x�z�Ũ쿛o�[��Ğ�,�.��=i�0Vj=��ڄI�����������7�p��U���s0*��h}�ˉ2�J��:�P����J�Z�2o#�d���S���
d,�!�����*ۻ�S6�U7�e�A�CJ�f%����F������V�	������K< s�'k-�ÿ�d6�`��+�X�J߸g��-��m�I"l7l����m�>��;�ơ�2�s��'L�k�$ �u6+$�L�vZ���=#4�Xq!%��>��zQ�Έb��<>��6@܎�S�J���
����^��E|������k,�m�U�\��_�L�C�h�y[�۽YE�^~�'{�5#^p�9�����]�k�F��y�;㥟 ��j�-�G��[((��j��<Ӭ�����GS���B�
���`L�]�����zܞ���RgQ����9�t�{�4v���&#����q����,n�J�p��*��V�)��M"&U���L������U�:��-Zu
��9��Ù9��ȫ3A�v돮=��m�|F��"9�����=M���Q�?@���F��E4+{a�SN����Q��������k&ٳt��C�T�f/�yz�]��P��$5{Hb.KO�mE�5xv�'�d�Y������e-�(��<��t���lY�!b�q�U��nЏ��eɢAOڅ|�e�M3�c��!w���V:�}+MG�>���Z��^H[|�����?�.�6_Z�����Q��8)�T��98a�P'�v�s��*w��lg��k'�ܲ	��x�&\O��e�������]{���K�f��c�+�"�P-aU��زm~]'*ca��g��H�!7���jA�fXPR���/2TϿ0�u�жjQ��-��@(jj,��~M�HR>���^U5�ܱJB���ۂ�u��3~�11��D)�Zv��m1jA*uY�3��������3��p|"�<N����	�7,�a=�����h;p4`M��R���i���x>Fՠ FQ �C�S��{r������it��0�-�X"d9��i_}Q-V8P��@�d���S0��(���Wu�~�k�V�q}
Ff;� #̍?r^8�������h���佣���16z�K��d�
;�2�eM5le�u�"�kp2�x�-zѹ��cG~>e�zg.ߠ�,^����ʀ�N�����k�E����b��F�0�WU���!�'T�V]�aj;8�OPQ{�{��(�}�T�T��Q��Q�=��&z4�l�ڬ�(�j�|qL��I����,��Y�w��$6!?��ݼ��M�J^q�w�*�KC�����m9n�_���E���<s����L7��A�b:���3m����U�UF��Ps��4O���2��#Ze8TPExA ��]�m�?��f���nM�䂡?p�����~�
ٷ�^R���/�� ��zQ6!m��	�
tF2����`����$���Y}*�4=?O�<��ʧq(���U|�-��	XTN���թdz4�C*[���_�$�ϩ�`��g(�A��|���̅ïܱ�y*5�%���E,y�� ���b����P�#�+3ee��O�L8�]�,m�5��0��H��6�l�������wd���Ӊ@� ,�E����ktl(}�3)��1IfA�\�#`��S|hq���(��d�JQ�/��1��hJ��Z�dv�K<��5ڡ|�c����d���vtNl-�:����Jw�m�هm����CUj�gy1H$�WX��Z=�;og	.2��^5�W��'�^�����&xӤ�;�.^��U�Ҏ`��T�����,.oA�,ۓ��P����}��>W�u� P�0	�a���}��]?�b���
�G��'��'�,q�9���O�G��'�����읽\xY^���n�>a���r[y8�"��	���k=&�� ����;̬��.�ha�-]���o�`��Δy�Ʒ��t/Q�کQk^�f~���a��66���B�H�r�n�j�� ��R�ܸ�Vw,����*R ~�:(�hK�zΨ�Z
Ť�4L�\hy@"����և��F��%��l�uA
�瀯�;1�"[E7�e�?3��u�xG��@�?���1����9��xi��}�mz����`nE+8P< ՞�*'�N��[] �T��d�l�z�\�N�A��֬�D)��"E�� ���)&��N%�c�3K��+)����SeZ��	�|4�2�B�yg�7��|dm1@���.e���ҽk�JvJ�m�7����Q{�ʼF7�W�"��8:�[�d��y�4��6d����<��܁ߛ��t P\okE�(۽�'��4���#gY%y�+��
���݂7��\����5/;ۄՖ�2:��a�)�!�SN�A��� o��1���v/�)�ػ�ƖP`$A����.m7���AÃ���p�