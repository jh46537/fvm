// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:51 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ciZCNbipAdqgaIf0iPHLTJNeIPt/3gcW9NKDDdHQpCQyoCwSP6GZAvdTnJ4EH7e4
V0Rc5gyLrsLqZZW8je5p4k5H1j7UxUDdpKHLBanyF7eJ513QzmmRxMYqAKJCDs2r
IkLrulA4EwNhXw2bEJYuhGWzHPBIZUp12uWVzwKlgMo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3072)
Nwy6pYK0m2GSOWYt1C9qMNUome210xutTWlODGM10sUchDFC0MIsXRM9c1lehjp4
y31zm10sk0hMn4mU/StD8KDcQ0HbInPs+iogjyZMN0GWrMst3UQplTKnRVvoL97m
TR4ji2XsWcOzB2PKarJehj7sbgfAz99QTuJDPKSR1n+sxRpAzTLZpcOsj388zkqB
dJo4nmSlLFP4j34CIfZ+0jagUN33HC2gW81FmVVU/yhmLxJ87jvvOuAzk46ngJzh
xWCNMMpGCCw+PQFmFLUoWYi+pbEJ6g1kZzO30zXhp6v5upRtyxz93BhC23jiUhAi
hEyB6kutdpkiG2as1/y6z6sdE5IR00fKpM5eIgnXQkeaCsYjwVaFW61YBaEzVLTM
rEiqgNx4453RzjSM1pJuPebXhOuKGVvulsRTRMQuQYzGsCb/SjDMtEgkQQXtX1lP
VMHDywGJSkZqroYqkbDO6zwAH7v4QOpBoKago+J+tK8RcLfOBk4ltH7ynilfZJA9
caXL2nx+2DeQn0zgNQahQP+g3Xv8lOAibqywiPgEGAO1AkDpw9nOOjnXjGSOXekl
iGiqC69jZh3gsWl3voDrXprqXnjm9TRK5q+kL+hE2TT63wREEeyZqXPnN5ixizbv
zJbzEBC/9lH4fhGY0mj8WDUMMUZhU7eW3gfUontldFkrF8jxZCgTQctoabjsgg1f
d063a3Xsuo1x6O72SFu3cpalbKg6HW27JU7kBW1NzNvSB6HJyUwKXSnVbQh8jcIg
NvxpiddD4kw3uohG/nJFtWb4BbHSyaKl9ljao6YwGEUI81igo1j1xrxeoyUzVir9
zT7DbBky8SZCAMIkYxZjeUJdeNPceF7d/nNLXnE7zB1VkW2Te3GXzx7GgwbO/Qlf
vxKiqtOY2ch3mP06KiY9HurGuSfYl2oJpd3u7F+AZPXMzewusG93gHB00sX3WdGx
N3wROe2ZBSSrn+sQ+X1lK42wfIiQkZ0MjHtfPNPZJSCZK8pn7DUnTsVFtV2+845R
YoEuTgKRB4htPirXINDYIMfKLdUjVezSTa+dfveTbahp4MdYtZLZxhs4OK/2//PY
t/liddebTK/9zS0t6fq1ZhXfd6RGyN8ypRp/02E1i+D8IDqY/Nln39tVeluDifRF
2rMIcM+f0L8rvNy1c30qWABVfTDjGord3lKDZ24fKwowmJa3OlCImPbbIoqSkMpW
p5Z+owmsvyEuXv+0mhwFAm7n2T2v73Ai7lzAa8o5q5Oe5oK97JEj2xmUBQc0Hyat
LVno6bPVx+XoSn3Y+eKuIcDe1WdjxbgtbRblfJDnqLoMH/9ygtGNy4blsrOaesqO
zEYkc3EQW5qkp60twY6luMHuz1kVL5J+AKfALSk1GSiwExvqaUnQpc8ZpYGs4dE1
f/5PK3cTlLZtgH7Tfu9ZMt6lMEUWAkuSh3nPugg1UQBVuAZmwBP9HDQv6j6htb3y
udhA2hlov1iEd2+44h+sUHffQk9Ui0Vlzc2k6i2pBHrBeI6tXLCri0Fw84Mz6emS
QeGmAO1YPcDCqgfyVrwkpAw6G1i5lXVOI1sVxJWBt/WRDYD3ZHI0vObDQDu+ON+e
NwYKLtvYLp7fdcfVQctUq4d3TIgDjbetf0U6D5NiWhRbi240sMXM6OIC1QmeCyS/
9f/wF2xLtNWckGsmEOKasOrUd3HDPBssvS/TpvWZdwIddvC+iD7W+IK87L0yU6nI
dnfBfPAJO1mMbXgFJtPY8ajPCUOLUxzEU/Wt842oLaKb5YvJ7RJ+/0hYD3Vc5TX/
YlbeQdTJ9zREiYyCkoUWGik+4UTSBBifQ6vJW8asua0ArZ6umBXG2xtlvZ7LN+Sb
mj7bjioKhwgUPphl+aNk/8plmj8d0PgZC8enfsCz/VnV9xrD0LoLEO2Opqm3nGhH
T1ZjYcxWtj6qVbojek/W0fTPzQpf6FiBudEFVnF29SeDkfKDdDxaiiBwyfrtULY7
fWskrMsFqDGNZkhq1aPy5oXU6VkODf4vvx+2vYCGwU0Mwt4XiBtYnWnljAbIqf36
BPXSFjc+Vw2UqYBQYaFcKOea11p3WrW1MPSL7qOEDVU5oQTmkObQXu18C2qoWSSE
pgKLHl2f46y0ODi2l26BXvfD46LQ+9qks28JH+cqNX3/h89FzdOOLG/uYdh3bl6K
EhwLrxxfGWfkcIA06SiYeobMigNNGbtwgKDlqyRp8FeGmomJLEtjZ6tAYb+AKm+1
oPDdwdCOSc4kaCsEeMGEI/2jWYrmB1suQHFWqoqQGQzIRV02RLuM/1lXuyjjhXj3
W/8W4QqqDVJWNpn5Ee257hqzqBZDFG0s7jdBP+QUWo6r0oCbWlnN43xeXDQVvFZi
BEPvpVxTrK4w7UkgcC90WSzjubRdOuXhYljCFPVowuIVdcZguRGZ32Y6eMw1XlsU
mJ3Fb/drvblvAxXwgFphIuni9b+VqZJQVVMdY+UlOP6V/speHHseCjR2BgcklqM0
6lcTg82UwYqr+kELhGfSlI3kr4QMtMdbRZoB09umFRm/wmH9nXVUdg5pznhF/wD/
y7PeRcIw0SmcJJg9WhAKwKqoB9ut4T0qdT4SJhi66/dSYT4fnoctmKFm6Jzfttkz
QI0Vx1V202YwNQ48RkFAN5X5SBP/wPGlY+avxVG7K8gTWW5zZbs9vPx9ZjSVE7i1
cSWvXscTBWUBhID3Ddixy9zXPjok7ZEPc+43qmVvt6wvIqoppl9FvaGauWji7rBm
dH1BuwjcYPwI8UGKnhRPTgayETkvaWWIPrXkGWVaE4d0mwty0tccwSOtDPcjz4+a
4+Hfj+2N52xqyITMRct/iDnTkpAAjxqrxTST5qRO2ri+v5+vBbTam5W4LO4vSkMn
LdEPpjEosTv0NIaSQE7CNuYM8U4a2cGZ0TuJ0SnW+FDoJ3a54p4v4VWXjvvi9Kbj
BgeM375l/gGc+hIwwrbVWBYxQA/DsE2B36ATHXqT4jlNOfQeNKvSZC8j79bOyHWS
meYkEqvu7mI7z0c1Fx3cq+3S6o3a268U8FuiGrwBLYfqtXjDegP+co/EaHWIdUkk
7EyagODYYo4ot6hLi53OlD57+nDQb5+xErWylResePpRAFvhH9uGkRr4F4LKB5x1
81eOEklv9WWJCS/RAY71P5j2IAkv9UoCMV3vItaj6Q7CkCz7lNCpRXu1HYHv1Owd
pVOO76nTJuDNUXL8urvoSIv3uLI6sup+va3QCvfPsME42C4d9TwsHmhPcSNszCD1
9uSQwnQyoKCqa3MfizDx1sQGQHQjbH1scYVshdJv+1G2gZw91VdJUFD/xtps9kpM
ISRXKwT1KkvtWlSDMRPjPWWyOeQin+ezuwDf4i+ZT5jgyE1yKaleSHANW+BaKklG
x+qLxZl2MRz21hSPh8QOxadUU7pcZRmtm+AmZMguCGJYdwVtomNbAlIQmIddV/Xz
2a1ug79JkGUsB4aN0ZX3hb3WCsRlZVd7DgdMXNGG3FGas/OUPVhjsqZIQfI1nII9
WQiWFKdDFXrgLU3raL9jyBergMZu+WWPM0/h5TRfh37l4je0kUV+80ERkwG4joeR
HnwT+AFKa98KcVfXK8zuxRI7AR6MKwdEwQjTy05eKJbY3ujBS4YFFbPQ/vtqwTmp
h59CnKUFaVbPnCtvEw/dJOEZF07Tf5DFW7wHMMm37ATT3/iFubSyOjALc8FluTd4
8dsTaBe5cjo8kJ4Pn48QXIhgKaIhTtro2IIld4PDnwGDFiII2y6ZkBI6F0QHYQtN
N4eSni6PQYsbUEa8ZGZIGk4Kad1O/m6AgKZSpcrDJsqnUdjgbrdeGmmC4BD/30nu
2QkF5Hq8pIMCcMdkVG5u5kp0jpSczoVVYhpBJwc/OjOQoWdT0U+1TuYLiiZk/PvW
gJLFuqyTd2iLboYaKOuXT+GHk1FcxkY0DiyQyepjr+LFJd+zluitYZ53zoxPUwfO
RP2o8vBAhhTsSqRw4s4H/8tMgDxUkZGdfoyFa8XisyA6CD3LaRtjvMyZ1Cw+QhxI
hAuGSC3HQQ/00Dd3xn92NKGUINCS8LQM1J0VkZhiw2Mi/ccuubtDo+Y3pZi3GsVr
`pragma protect end_protected
