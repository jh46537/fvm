��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E��`!��O���i�*wX��&��m2�)j>��X$�Fv�Mfca�e��q��1���:�vσ{��e�b�Μ��f(g^�}���S��x0l��wp��s4���圱�I�����@(rS�wm/�.
R�Q:2�3��>��7.�[e����r5�-�I��N��L!�V*�\�P/�t&���<�d]�:�pC�9������M��
4|�8%4�ҳ+;+q��v���[��pr�����dd��+m���	����A�Q������	ȭ%��.Gr�����|a�-�ąX+	W���5�[��oAX?�G�^�L_�_�q }�B�*�-�sJ����0׬Y���l��E��)��! &���>'�F��4�rO'��F�~���dy������K����rmW� ��N�%=oP�5J��~|{��F˘�>����2kRS�sZɋ��uʴ�S?�S��j���0$π��,͋ ����b�hB��!��������흡Ub�y�觋�9�K������g�c���u���i(�lƩC�t��Gg�|�����dk����,2���^�^O�𚙍��^��-�N��K@��D��|V�8�Jf�B��1�l��2����	BN�	�3�w� �?)��+<\)�X8���'��d78��[W�"E
ov���c����F�����K_��C7��ڙ��BN�!���<3o�ǉ���	uR�������Y�LN��m�� tY�*e�Z.4r4)�覡Gӑ��V��sAteV����#�����Q��WsN��=) ���C	��D,3iy�6�a̧9<�y�1�"��m��CG�a�ċ��UH <n;�K�3�.�׌��0�r0m���r-��~��9��Ui�ñ�p5P*d/�s"PT��;<WBFBs�8f)lЮ����NVS�� E$ڡ_y0��'3�aE�6J�J%�&� ������Qf۱��c�Ӭ��L5��B�Jv�����fL89���sz�n����&u�Ǘ���B��9����K�cY�|�{���O"���mcl���S�#@�<NK��a[���w[Q�\��Gȵ�#�
GB.���O9���i����P�Jr�M/�6asx"D�~x����a�u�V$?��=;#��;�!�-5�\- Qy�"-#�m��R�<� Æ�Ԙ�Lmn�y~:�=��P7�� O�u^I*�l��3�t��R	&�y�C�1���-�|ϗ)k�&UD����/R��<��K���AWpA������,W7�9����	��𤎔��}Ɠ��[���Ԛ���!+�׶�;;�[�a��Y�{�
!
�#nb��%A,���nU��;�$v p��.~�֊e58��i1h)ל�S��:oPG�^���֠?�5����G5�/�ċp<�gx�tr�&�`IP*?w�(���_JH�?��ٮ1��Z`���P�/�-%��#�)@e�r�|��#j,����J�U>��/��K:Q{9�p�����A��.y���t&?y�dyX ���^�2�z+(u�;҅:J���y�%��4t����j�5�<�����!,�ǉK�߾�&i�Z-)@�X.O0{��Tz)wI���(���kRj�FfIL����S��F��X��*=U������1�[%�L�B���k���MB����ew~�m�褠A���Xp
����L46�"J[Ik�TP�"x�B��/
!����TC��X�:@�������mcl�S�i|gB���PY��O?���q�6�Q�R益^��/�*�y�E�H��[���f�#G�]�B!+��5rW{u��7�_�[���#�d�z;�`����[�j��ew� �����~eC���� n'[�G�����L[��M�����oԶa��d�@�6��$�~�d��	�_ې����_Q����뤙1)+�sR��'�:!%�Z@z���o�t Oϸ�ˏF�@��6&�`@fB�&�鍺�� ��\��|��o�נ3n����h��X��h��L�bs�e�=;�4X�1���eV�i"h�b'�HMή���Z��� 98�v����K'G�s�r[H���i��/fR7E��d���������4Oe�R�k�Cx���<;�n6|�G�A&�����[Py�kqf}�����Id���ÐLL��S@����Z�w��������R}	*GӭH'�;���z���Vl(Z�B4E1;�ա��wd{�Q^-�g�nW�d��:�7�o\�%V;C�E�������g  3�C�E�{�٧�(չRs�J�v�-q����R���������G�#��4Y f���bDe���e)��4p�b�6�����g(�X�t���v���ZRH5��<���d�]+�����϶��m찖�*''/�Y!N6&Q�%Nr2b��@R���I��Ҷ��Q��؇Q�|ʯJv�*��K���nFIJ�<Ԩ��@����%����F;�k��4"�&��Iئ�iƢ�GÆhhg��pțd�/����*bT;�[y³�i��d�9�c�I��ߊL>�N6�(�9F^��[���`ELmMʞ���^�4hqXq��w�_�w旇.'^�y����x��ha�~���!8�g8Ȼv�@��tn��}7���wv�?���2�9���b��Z�!	�oϐj �i��OBE���S��!�np,�J�F�`��A,K�^�3��}�M�/������-8봁���n(J��w3�ֈ1����*�g��Ɍ����)λ*> K�O�$�Ư�O�Dq�K�ï[�^6�nX}T#�?�gpW�b*.\ǚ\
���$�:�]z���*�	���##�#�n"o���L��!Sn�##��=T�0���YOl���/]�,/uX�r��%�kj�U򳊥�������'�˖��F�n�<�v��F�;���}�;V���8���C�w)�	��;�M"�?��+Q����Q0������ �����b�����4������4�T�9ȧ�"�f�f��]�x@l��ިxU\�-\�7��H~t�Xw�6���Q\�3����'�Q��з�XG�����9ޒA�Qʩ��t�׉�9b4T�RW�=��\�ܖʝd�8f�	�zqi�"���5R�;/kQQe	��bg�i�����v(�؈�ŏ^��3�k:�%um(��r��-���<�ØāO��Å��#��J�4�����7�l�@1)N�"z�(7�YC^ò�Yr4w�6�|&|9���l��q�4���`zμ�U�����E5��9+-;��Q5�3+��7�+vI��#�/_1b9���b~⌒W��U��k�5K�b���S�8��}�dN,T�l��o@Q!�7�o�l���6�exy9��)�)L�FRxD%�jj�k�׫�4�s(��ټ�%���jO�A�?�=�<0E};��X�m�G������|Vw�l�*"O�bL��=%�֢A���W`K��&|$��S�-��1���ì�5�܋��V����u۹�j����&F��� ����H�����>>V�_'h��N���"��}�siU��Qz����C	D㨘a��m����E�*<��¶r�<�j�"��y�,y�E���9b��iҍ���)J`�*$Hbb��0y����FX��!�"�Ͻ��z��g4p1��9��ܶ�0������o�_O}�`lS1����<Pa���A�D���`�<�<����3����8S�1��W��^:+P"�P_3q�5���.�?Q�	B�?2�
�P���h�2L��Oː5H`'�@@Ԯ�~'��f#�ޝ8�*Pġ�s9%A&"�}���L٧{�Ǜ��b���s3<c�w�f�c��$�ן�*~ة}�h!���X��6��3��E�럤N�I�na��'��� �芥|lĨK���A��G��*�d�����N���-�tz�2y
��<�f�>�9߾�4'��_�[d΀�vst#rNpE|��_����U*,�!�d����R�Q>(#g䗸S�X\��:	���7��l3Ma���;�� ,�	p����|����� ��s�8e�����c��YԻt��� ��7|����;��E�b|�L���*ڙj@���PXOᙝ\U3E��G��x��<���A�RC�S���Z�K�3q��B;=�2� �����)��^|��e%����q�2<�$�gO�k:�
���1�7�[4 ݇�Eڣ�� @�v����:jQZ�ލ9���gi����GQ�c���1x��Sa�.;��7[!zOhG����o�ƔS�p\S'1�b���8��+qt���!^@6	�r���E��R�3����V@A�ي4gd���/)�l?� u��HQ\[YI�y 옥~ yZ���TD5���rڋ�x|�g�=�����w�e�[֯��k��;����o�(��^2�
�C��,���%\�qw��7�g`q90;�u���}ʠ����{�k�,Nl�׃�����nG��䀥겘T���R|�z�J�,�
�F�Mw�+h�Vt�q�r���3��|�޴W#�i�8n5o�"�5��b�[�8�, �\+�3�IG69}d��	�a���1Z�]��56<
���]V�㣦�ť�y_��72�HS|����`�^�p�߿ug�Ӥ��;tVs��<K<H݂�7����GHk�2��Pʰ�lq�\�dNP��h�r�'�Gߣ�	����6�%��O'�	X��V}/Q���/�kX��W�Ң8�w&�����ʡ[�s�#?�[a���h]g�>������B���h
h��;0Ӌ�8�5�Qx�F���f���l��Z�� ��v��1+c�s���,}==[��qT�kI6r�mhm�e�\-����[Pd�ה�n;�n�im����[y?mS��
��v�v]"$��=~uZ?F@%����\E~�P�?	f6��cB��{&���1xA�t��}�8Z���A	���Vt��I?0��?���y%̈`�ƙ��q�6�\�"�ɣ������Ha1`u{���}����݋��	簫+�I���4� و���Y��`Cv�M�����=�?q��S�Ř�_�lx]`����?k�U[;�J��ޞ8��f^��="X����ă���.)] n�z�
"ph�rو�F�2V�k�zS�<v^�� �%�5mZ�Xo�0J+��8���B��qi��a�F�J�.{CA�%UZ /��9S����SEZ֐��j�a��s�v��Oh{�$����➓�׽=�&���C_����
�g��ϛ|�XXݖ�91����d�~�?���@+�زn��+�E�j.a����Va����ҁ�`�Y���F���,&��Y/���R�CW4�Ri#�(��Rf�NL;�΄A	��#{�O�_��ޟE��WsC�C�
?�ty�k2���_c��3ٯ��[<��i/�0�7��fbK��"� ���
	mJ�sL�hVV���v�������7�:��Ȗ�?�z�&�u���oR�!n�	=0�ĭQ-F����]9�N��ˠ4��s����B��<Y� ���2�05A�;��FmT���	����/mŜ�/@�Hz�����A�u��b�Y5��
>!S��u�����J)��⼐B�A�@��u���`}��N)?G�u���{0�~�rc?�n4�y� ��8�20��7�� ���əձ�:ʹ�l'��r1(R>3��J�~]"�����<�����C|��bބ;~�_�i c�2 Ԇ��Ӆ+23-�N��B����'