��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�0�w׍��SΪ]�����E��>���r�0�n �7<=N^[���|k0x���J�"Jm�%�O{u����+���m̥�D��B8m�P�W�u#�B��������|���}Ɨ��Jt�����ڻל�]���F��c�0�-*�&��J��?~:e@�Uo�P�\^?YB�F��O.�3�펛��J?��I�G# ����>��+��PW�}�֡V6cn*���y��WBv��E���U���ƫ�-�
�������������tp�D��.T��e|����W$��	y�۰�
!��P�!f\	p�4���!^�׍}�9$�muk梧D�7��s_�N��H���}���F{�=ۭ��㩰9�ed2/��bX�\d�%�O�б�I��@dm���}[����pV�E̦�%_T��J�??�V2n��G�˪�*n���u*;��{�P�$��7�x�%n���>�'8H�v�����T� 
K��J�6��
�7)�FSհ��j�,{��@p�~(����\/���h�m�)m�OL�w�RX-��]*��.�,K:�!|$QPX�=5�&�r�@t�E�X��t"�*��s[��|q�C��%xj
h#`�`�P��y)`�j����k<�p�������"����ӥ�v�G5E��d[�m��S�)W{�`� �꬞$��w�u���L@��ԍ���s�h�]�}|�,�:f:N&Y!�?�mf8e�Fz���^+�Tib���"ŰvШ�������+�O �iÅ���Ì'yp^�~�nCߖ�cW�.YV�[��T7�8���iHt7/����y
qz C��~�DNC�T�����M����m%�vpJg�j0\^*L^������VOj�XJ*�׶�\w�D�����w������1��S�+>=�;NP����n �i����pb���:ǈ��t�;��ѫ����Z��ox���1|NA!�g߻��oɻRp����:���X�%�8��۸����6*:�!���r����Uc��X�&�<�2(�=�P`91*����tu�,���tN`�r�ӽ�6��R�u�4�w�Y�����e�Yǣ"�E[u����u�,�a��'�G("�!���v�W�\B3��-�(u<\��ܖk)d��}��Q~��,+
I�J���O�6u]�@�y�t���u�͘�o��
M�	�LFIϒ�Y\EG��g̅3��S8G�61��=Tl�D8�%�2�.��ka6��	Ѯ�/�W)}�ha*����K����C2����ڧ?]:�u�&!}�<��](�����R�/X/Ӟ�b���Мah��7�a@�r�SQdĖ��y����`?쨌{�w:O��3$H=&��_��J�m���GN蛕�� ;��򙰖o��&b�_�f������H��6�z��3��71��Vs�"*U���{Q���Lg���.��-d]R�D�O�߇j2����_S�W�'>c�y8 �s��h��_i�*��f��"�4c*��`��� b�z��(�l1a��r���eB?�>���-�U�o:���'t�����+�B>�WBL�����6�5x�{��>���|HtP�Dc����%��W���l�t(��&j)T�Tu�������H]�^�����ܬg�=����LI)#�Z��Sl���z�^lro:G9��B�SS��H��̣5���?��R0�����Sq����A�؁����tM�m@jj�$ك����j��:Z��ϲG+N�����	��	�x�p���\G��9����e�b.Qb��
�e�mxk ��I�'� �&}@1�B0�c׬��zMi���Ptkh\�,l��f�MʡOM�(Ȱ��,�ci���qл��ae��Z)�����k9G�ެL�&¹BH'��4U�"m��X�/�"��>�h�+š� L�3wp��_V$ V�Y%�ѣ���U5i�����fM��A��O4�kGڰv~��\��r�2xsa�kذ?e��;��$eցMFe��t鎗C-}nvYGÝu���0&�)���A^ҏ��g� Q���ЁŮV�d�y�IE�e�����Gg#0���H`��P[����4�8���ո��qB�]c�
I����H�-yڞH��Z���J��x^���|����B{�g�W��겉)�I01&����JM�+����z�dwWh����^9�$*�� �:��2���E�pN��4������)���1���c[��[$���#��Ç�<؅
�����;>0�Ϙ���8��4�ٶ�d	v%�H�g�q��K2�d��d�J'sQ��Dt�Yx!���E���$�/Ic����b�`�w��N��l�<��;���T��Jr�^�Ң�,d�8!�͇�0j��\c��E�9'��󅇸�O0��\gZT&Y0��f�zR1�h�:>J	.fcI��R�S�8��
�zb���>�J��5�>�;����G2��Ȫ÷)��6r����Xi�_��c<�t�3�x U?�SP���SJ���d��_��Ki�I�I_aP
���! x�x��N�Bcӳ���]�e�/�i���
�c7VO=���x:��4Þ�`'���˴��Q��jS�����VG����tH]�<�u��z���>0h �nl:>�r(R�����-����ZY}S,��~�/o�G^_!G���0 [,�6B�)A��j�0�nbyd7�WW�����4ĤN!�~�O�Ͽ���I���	�l�(n�_h#	
�c�c���m��"-�A8�tq��RuR���� 8�.:�>"�<��@�ި���hBt��Ϊ�B�����w?�7urW�M�|���G�Rڞ�@BQ�F�ދ�y���v���
�#yU��'��dmT��lϘf�^
<�$�/����&לJX��W�#�N�Yw?WS�m̗��j g�,@H�+�ۊ�D�<2���و�
j��t��G�/�q�d���>�$j�Ʈ�f�A>�*�J�o�����nA� !��H�{����8;R��JO(�R�bKjb���*4�Æ�Q�M"�1-aK&|y]�sa���zvҺ ��E���2�-(+�����E�P�c����.���lFNA-��6߱,�O�鷉b�vp�򐸆.(��m�6�~��CLW�w꠼�V��I�`�u�o��8�5w�>���|�^n9ݳō��Q��o[�����$h��}f-d�4+��լ�k%���LGj�������g~8^�)<vd�x��X
IFh�C��Зg%9q?wt�Ng/#`�7��$�*�U{a�ԗ���ơx
T�T�+�6Q���B�ܣ}{������yp;�c������F���F҇@3�q�A+5
n��5S�B�A?;@����� ^�EfQU�&D���/$��\Q���'��2E�!�fs0sB�Da
}%}E;~��r�1!���(���|������Rڼ-������$//�{LY[���rP� 0��p�ʬ���ڍ���X[�P(A�#/�pp�ŕd�����_�t�1dE2��8� ��a���
,glx����ͯ�@��Lo�	9k��K��+?��ƎZ�2c�t�ڏ;�x�c�����MV�������;=��8TO`���	#�"� �p�J���mH���� A0��os�J.+�wEY��"�s�ߤ�],�L�>���/Ja�{o����'���Af���z��d���[�����s�eRM~��X]�Βt�=��zWؿ!`�e6Y�L0�tP�&O?�ż�R�2
��z	���`g�f�<�X+��[������#��#@� F���ȥ�{Q	�ā�7L2�ɁZ鋨U�f�v>HM�:�$���K�����q��H~�zs��U�C�_��L5l#��}�T�L�;釀���X�u@K7��h��0���X��cv=,�J���Ws�~������y��G���g�m�Z^�����	��o} ��e_3܃z�!�4ib-��)�:�jF�s���$�J�  6�%�W��[b�dcj�ʭu���(A|S��a �(Et���� ��_D�|�p����C���W]�p����<�J�@�H�*�������%��I/�/t�kݪ���� ��싊���ք��� ������[vnmg����2�ϭ1Q$z���>Z���XƦS�|���PL�n�M��EQm�����K�K��A�	S�iN?�QƳ`_K� �+'���tЪ2��f+r�x��̧ͺ�	¢�;O���l�OVO�6��:Q�����T2 ������G�m�.Y��:�?'/������[��@K�����&`�pK(#N�Ez8�3%ِ!G�l<��4�ң�֏-s�u���uh|	[��3���cO7���