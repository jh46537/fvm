��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� ��
�˿F!����i�xL���G)35�У0�Y6ɓL7ɶ�4[�Z��K!�Rʶ�������*�r��ug��51��ڬ�v@H�f����yp�1r��^#�����6euo���\��AMR(��=�"�Ms��HY#镐�r�)o1iQ|��]�L��|X�@T`���W!����As�MŊ[�6���%�|Df��2�v=�4����i�9K��Y@�Ի��25}�)vWv���{���"C~[Qt6'�Ftf�h}yҫ��/�c�ʍ����~^5�5���L\1) ��f���S�d�J�W]*B���L����F%���{�`y�UfS7�ms=���&f�sB��Cp]c��G�k6o����ƒ�=>�gI@�g �gWg��-�o�W�5h�ڣ��Σ,B����U�����3!�a��#t<< �
��o��iE�#lPZ���q�A?�]��z;����Pe��P�o��3O��	Dƃ/9v|����$��N�Q�1�ap��MQ��k>��R7����L�{?���%����E�q���+[@��	4Ɯ���^Ԣ��'+Go�ZQ�T�����۬joR�h]6�1X�	�5�'~�C�P?�_~���C{3F?XZ_��fB�4�;
;M9�+�O�[>_�fS����qc�^�$A�GG�굮��5�T//_P���O,�v�Zb�!���j�r�\�� �gH��?��ㆣH��Z&
%���K���?���?+?�cd�d�/�٭F�IJ�:3ne�,�!��ϸ���{j����
��%zܞ`M[��E6zt ��F1|xc_�0��t��C6�#׮dȌn
�Nç�B���Ɨ{��ԣ�8c���q��X���{=�j9� �mKw�~5�+�x&�ˌ��ʹvn%%�j�����lgYr�&C[ܱՉ�fucg�f����V���p>l�W�0�=��bڜ�LFk�eAs���9�}#������J�Ѕ�0�Z�����=�kr2����<������C�k�����Wnf�$���^��٭Q��ލ^�SW�+�����dq�L�&�l`I���T˒�2�M����DQe���n]���g�7�m�pe~՘��W?�0�>�A�sx��#L�/ɦf�X�=N�[�S)�u^%��$�{��COE,���*�_Q�2�%�y��@���L�V�Iؚr~�*�SZ��:��\������WLG�P�i�"�N�,��~$�μ�-�;�f3�6d/�Rf1��!��ۡ`c=/^�0ւ�K�61�aR
��j�#���-bL�l����<�z��u3���\�����:֛r9�9�hD]\��:���> ����Ԁ?�_?�a�1�� e�}4�E�YYL�Ȉ�u&��D�n�(�dw��q�峳0�r���@�؋��->S��6����J���mN��yޜ�)�����.���s	��n�{}t����],�3�����a��p&�|���=�o�U�lS���e�MbU�2k)ζ.�&1�E�W[�b���_����oi�u:�jd<Lb��	��7{w�t�M����3\�)ep�ϻ*��`��T]�[�U��� X�T^��_�Q���ʠ�i>�o"��
�|�3��&V>�t�_ ��4˫ߌa����n��'繙�'�&��%=T��E=�̞)mjLI0���4����:�s�ѓ}4Hr`>�~��˹}�j�J M/�1�%�0���i�<�.�Uh�H��V���VT�����T�<;d �3ԅɫ+�O��1פ��Ա���v.��3g.��7x�����&V"v��x���}��91��w�K%��nV0Y� ���z��큞hV�,�i;�&�"%o��2��Ox/����t�V��x�V/V�D?�]iN���nТ
�6o�4�'D�Ykz��d��0u��~�&-�
�l�%�ePgf}B��AA�;v�9�1�_��E,-�ё��o2'�6zr��Ţ�L�S�����C�������$�qLK3Ic�-�I����h�T���	|����ʏ�w0���#�/��/����y�X�x�m��*ZFu+o4�>����n��(����#��	�D�7�R�WvS��$T6W��%݆��C9�q$��T��xwNP~4�'��m�Ρ��0!q�����,ЧE�s�.��o}����_����"�r�Q]�C�hzsM�wx���`��i3���-��{ 6��3#�s�3��O4	����>���G�k�2KO�2'�C�$�� ���D}y��������B#&�b`~#����I����+kY_�l�%��,��s�2P�q��_�D0FjY���L{��x-UJbÚ�j� 7&v��a��4�h�����Y�|䟏�M���lA2��]���oYM.�i��S�]�m���BV�ķJ)��q�z�v�0u%5������x49o�G��S��{�����8R\�;�Y-3�G<Z���c� �̿rM�����a=ݑ@7v➐��OVYW�T�E�B9;�!HE.�1S ���l�ݔ�M�?��mdgM�:�!�l�w!
��^;5��)2{��.^�� ���彥޻�|BG��i�
G�i#���� pRƶ�����d��JC�x��Uk�Bm(W�o0��Ց^�趟��*���ڱj�,>�iX�d=:��'y� {��^���@�{h�V�=�@l��)[�Ͳ�.��54�X�4K�;P��h,�v�ƺˉ��9UVVXV�����������֬����&���,��Τ���A��h�)TV3��?I�x�+5:���k�+x�^�e��$䎅H�|"x�_M�jI��y�l�I���'�Oh��6)����T���&�r��>�*F�?�G�;�������y*u\���]�	kὖ��D�F.{|l���>��X,�������?IHU�-�gb˶d�ζ_�|(�kр�dV����A���9,w���o�Q�%5�i]Zď�4C*����!b��݄���gnj>�Zo7gRR�)���·��b7�(J������Û�;��]U
7@wVq�kjE'BWt1�˟"��W�?�W%�u�䖴�;�1f��.�5m�3�l��p��*Gx��R��v��(թ���ƣ'I�����t����L+�� ��I��)X^T��I��:6u'�����,)�M�"� , g*�z,���R�>���%,a<�"��_F�dxY��.�5�D_KeI������m��U<�/��Sۜ��DZr��d5���Az\$i���f�?�����M�}�T$�w+i^J}Ÿ)���/27)�zn� �<�|�K�>������b>�|]֦o�r�Ħu�y�S�QD�p�K5-��ݜ����d�3������~��Ƭ����[�W�sqO�m��1�)��F���AdD���B�	�:=�ʔ� �2��������j��S�O삷5s�l�ێ��ﷃ�b�%nP�V��2���ƍ��ʼk���	MT]�ϭ��^[����b����/s �i"���Γ��!�|HH����Vۦ\O��t�o7؟�D��
f��I͒�ɟT�|��ll�L��q+�^��0�)<ݖ���+SOqƒ]��}���d[�A�BG�>̗��FE���s5|լ$�eV��F@D�f������u�JZ�Fv�p�6��iQA_�4�o����]o���i��H�����>��g�����<�3O��e ~��&��M������"�������L���|�kN;N�
Y���X�I4,\�y"�]���޲��p!�N��ە�e�ψ��ɭ�0������#y��'�H"R����WjNVY}�T�c����x���z���
H��n<v��P��SHj�BLւ�I���mR��t����b�2<ї�Uc��8��J��gG�}���@�o