��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�@V����B?:S���/��݀:6{�#���cH�z@pk�����+� ��N��c�|�v��i��oZ���i%�����b���O�eQ��[��5������#6��&�E���'�2;k1ř�1��2��!����23/��N�D�����c���.P��`'Q����q��pzjсH���
�٩�"f`B�~���U��9�I�ɨӷ[�=y�q"�k�2�R9�k�7�ûj�tf̄IZ�8,��Ff��P&0?W�Y봐�N����.�ئ3�vi�c�[��ڛBE#<6\�W7B�������)}�#l��*-�i/v��b�aS��sP��1���Ǡ#Y���cu����U �1ѩp��W�󶙬�%V�����\��TY���������5��O�2����� �W�K�j��|����}j�$�i�����QE܃3����s�"{��'�4z�/��sC7(�6��q̾;�Q�>���O�?ےG���|�v�\%}�cpo�2v���a�Ј:U;BAJ��k��[����V:8��˫	�2�}�ԍ�_u%E�h��<X-E*w�-m�u~X�����֔YB������p|ܴ~�Oe}�7��LI~{���OM>�n�ϟT���
�5r/�c}��� �����K!����\󵽭��mO=�f,	9�-G��k󀄬�G��>���E�����UA��t��tH�G�F���֟7��_�Ĕ�o�NQ-jLU8���K�"�OH�����rQ�}�A}	���� �V���F3�J��<c����}����l�8�w]����f���c��}�p��T%=N���=I�m ��"+A6	�N��׎s�z�=�
X ����}iH��$������V�>���[6a��[�[a��o5���M���_�jj+���9$����� '���~d���랸�Э�H�
��:�H���0ر�-��� e|���m�@��W8̄ś<Vۼ.V��-�S@���J�6s���+2�8��8�  `d�>��̞h�TA����H��#&[p�x�lq2Mv���춨�:a�SMҝ�B�Mܩ� ?�T����"5h�_S���1�-�(�*�jX^��CO��b�ҁ�!ʆ�lyM��+O*��V�t��H+�nȍ�C$t��!}Lz�ZzZ�Ӯ4������M/����F2g�N����%�Q�?��7���b�E�7@i�w���=�`���,��E��N�=P+�7�c�%��X��/�uH�@h��{������[� Z3�ǝB	�]$��~2x��Q��y�!�y��s����ף���K����>1�4h�@I8oǣ����/�!d�[�Ouu�u�9J��d����x���Ѱ��-!�ʫ���E,'��[���	t!p�R�M����7J��S�{��,��C�d�l8�'��</��V-�.�0T$� ��z���t��S�-���e���a
l4�(�٣(�5d�Y�7�8K�{qL���7˚��}/[I��m$�38�����������
�����s���� �V.�7^�xB�!�-f_���f�V�$@�Ƒ� 1�x�&�eq���w�uj��-&�\vv�B�b����3���w�g?Š��.]�E�>�N6��
�'�g�� b��<h����e�;Y�9���N}���`��k�o^!�U�Rs��!��"L����O���:�1����d�J��'��\ӏ$w���`!�.q�>�b|��X�7�+�=$�]�����y�j�(�~���� (n�f�7���cH���)�<5T�_+�A����	B��E���4��JI�(8���~�&:W���(Q��Z���dvF�&���y�j�X�n�?O��ab��%P����UW/�ǜB���'�Oe�46�(6<C�N�eq��	+��I*Z���up*�@��_g�yL6#�K5�oT\���DZ��
e����R�7�w��pS:ph�#�xT.{��#N���L�@��?����+Y}��[��+��ο���2af+0rGg�"IqG\�DT��[���{�w�eo(g{�KV�6�J���A�|����_�x����0kC��
�񯄹1H{�,^sM>���J�	�ЅZ�9����D�P�3b޺H�KT��FAv��[���E_���Qtc�Ȯ�Àgq=]~*��7���k��[�	pi2�&��Y�h��s�v�.bc�r�5�M�v��"�W��� q0Rbiƭ=�b��K�J���	��O��쬰��\�����h�[=��^P�����?��:�H'�\#{�B�5�+�-����l������PS+�h
R�W<��1{%��+�3��fvdTv�c��B�����F����U3�?|^hg
������_�T<׽\N�	"��b(�~n��[j��Pr1��4;���P6��٫��$��N(,�d��.j�]6��Dk�s��Q��݉	⏾e�|�@w?��)�A�7����!Po��,n�1�����M��0�٩���b��O-��|�!�~�?nf�)6F�AN��2�o%�Lx *���2$HdBI!٭oh½�,&C�xƶႏ��E���z����3_E�)5�3c��^��
�vݕ��--�z"�I W���k��`�����&	��dW�y��>JJ��I��W&�(��q��d]A�����bGm�����%��ٙ�C��詡���������B�)��L�X֠v�G)��U¹��R��B��Z���[����)��5JxwdQ|̓���ȸ���#;	�g��iF����X���� ��厱���-"���!`��ѩ�����7b�<��sS^�h�8�?e�a�n]�_���A^x�P����ŬY����@��Ȼ�0.�!�Z���H�m�q��I�[�K:���0��Ht��D�����/�o��&/vg��t��~h}V��1W�P���BUđ���0\1�����LT�D���=/��y}��5��z]�mH��q}nh3���|Ϭ����z]/Mqp��p�)�����5�D.s#2O�CK��/=��殸�/0��k16��Z���69(�W�
�����5�1l@{2IW8��+^?VJ�)��e��K�]ffUo�� j>HLm��@�}gv�j�?Xd�(k(q�/�uo�'A����1ؽ
�z�[H�eX?)��C��E0�eI8����I��>EL&/�>�+\����XS�T�7X#kA��4��aa�~�{}�n�lH1�X��������\�c�gx�U��6\��Xf�;K O����*[|�44��g�4��v�n�S����%��hK&�Gm<�����yi��*ʴyB`�`�(�Ek{�'e[���j���M�bg�O܋��K�.]j���	���[#����UW��_�Js��7nt��%GT�wW�����na��'�q^\�HQ�$o] �`�f�8˅
����H̍5�R����D���o�;�-���	��c=&I`��ʠD�]�:�]�a����k;�:�Tf��U#� �h�*(u�n��3�ɋ2[�=�׺�w����h��:��x<��g��J�׬s#��e'c!��+�v�T}C����7Dc7�3�9�#�A�f�i�:�C�� �ܑ	�%��1۝�9LNpD��m�n�,�Lѥ\TĎ�ͨ�2����p6ف�����wG��Av>p����xh�����u&Nc�]�栟���q���D��a�J �X���֑�p��97K�YO,�6f:g�$\�j�&�,�� {���1`;�ͺIZ��W������_�o��'1M�4�}��O�m�Խ�=�N��\i%�)�w(*���b���&���ӡ���h��;�����ӶH�8�4p|���Ztd:��X�:nh�4TE�	�i7)�L����3�2�����/c�(��d�ϲ<^�R����ӽ`a� Y�w8�q�H5�N�,�'��4-�m�́�R��^m�Tb^�{S�����}�l���!�T�?��ʇ��i]8���l�Cx�c�8���҇2;z�����CB��,Lɧ���P6:'�g�H*�zwɳ��ү�@'�s'-�Y�|���7�eK<�+ݹ�w�����}ݜ]@X�4 rd��,�
nL�g��m����,J���^45]�]��7�*�6Q�/�3�ӝ�@:T����!�s7�6$n̶q$�^�.:B��W���&��̮�a�W ~��3A�뼧�llQ	��u�Z�~ҍD=z�|IAZ����1�O�5�oe�𬨇����OA�"�Ȑ'�o�G�	0��Dt,% 2���2�����oE���ϏC��R��h�%uߘ���(G����r��jp%��1�Tg��5jϕ :)�=b�!0�Uo�����a�k�4عy�Ȝ����ɿC�����X��jX�(Ӡ��N7ukv��V�P��"k�Y�5kk
˪��@^U��6�n^[�|	�SnJwQl�NlU��1{��Äޖ�p�ӵ�L�����!��O����5G�o5?Y+�eE�_��[��a~y��=�B3C[�R@*�O�i� _��P��ş��Rֽο�^�W$opg�d�;Y�B�0�X�=���Ta@�?�"��͓f<C[��Ĭ����?������q#]]
N�����v��;�V�GD*�L�nR�P~����a9�J�YK��P=>��n5�٢>��Ł7}���� �A�I���f�DE/�2�H�>��*����7T���m�u<��x�[:ts�9����Q$I(�G�[j����,��~S�&�����R�p����G�<�oQ�^�/`��{Z�����1Z5�v���Z@���6�^���23T�Y;h� ₃�%�-+vvĚ	B&9��#������j&$����RqT/?ޙ�=��F��{k(�o���Bf�u�Er�Q;��$ʝ.j�QnLU�Q4���G2'�;��:��ʚ̔6�U8��꺒�H���p������H��9&:���t�JɆ�^3���a,?m/k����)����d�%����Kl,s�5lK���IÚ�q���Ÿ�N�̒P{p�Q�c[ ���V�>�]}{�����T����u�X��Zc�O#��^�$�N��w���S��a�F4��/�yɭ�=\7�돴0mة/N_RH���GUZv���h򗬫��մz�\�