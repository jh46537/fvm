��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]7�2���cDP�y�2A1y�n��#�e�qI�/��u�e��|��;��|�2q�"��F�c玗�{�)�x!���9��g�tT/m�*a#�	�^����	���c�Qwa)�Í�����Uޱ���U�m��V#���o�O.�m��L��R�g�������6և/0I�C���t0�������à=��BJW6�&u?��j�_3���O5�
��X��.����X���^�|���8Lb|��˫��\��w��Mh�o���iU�$?�a��u��{��n�D�es���pS]
�.*�F�z~|��<h��)���S�A4��enKMm}ͣ-�)~��ğ�I����	���Ks�C����q���(�T��W:��e��gi��<R�Y ��U��@�7��LQ"k�̀���NW�q�6��kpV�$U�n���x�r�.�t�0�m�c���� �����)�y�&Pժ�i��T�A٥y�C�;Gg�p|{Nc�b��@1����v��.D��S�%��'�������Õ��4$<'�X�V�����i\mMf3r`�#������+�`(M���oY�aw�n�J4	2�;���"R�->t"��t������(̍$zJ_<�ZZ[��&0�u����-�0�G6]��u���k�"a�0�W��r�!���ݗ�Wo��xw�I<#���YE1�r�Hb����@��W�;�T�2n�ɿg��R����P�=�R���kH��RP�߀'��Q�ҁ�C�'?l	���Q6ϟ.M��u{�U�X,8�_�eCg%� B�v�6�?B�P����Z����Z��oV�(Qpc�\����H$,�	�)M7�U��;(bũ�
�D��g:0�8k_Ojڵ/A�8A��پ�����`&� h����Q��!kF�k���(C?~3<�L��G�%�4��1�(���Uk�*eS1����*�J�Y����� �7
g�0������R��Hf<DF�v��m�x��&P���ˎ:=:�%������0TZ)���'��'J�B��ev��D�3On��M�t��ux�D	|��9Ѩ�F��x����P��m��a�쬒�kb!��p1�Y��FR��l&1�hGo�����+���~~��U�܇�y�C�%�aBL�@S�2��׿T�����V7weN�p���$+��i���5��hK�h	z�m���`�}_��1�I$(*�{!vڏ�����f5�Iˮ��u.2S��CA�v�wP�	��-ٮ��_Z=�M��]��e��PR�,��X��,a��
{��#�돰b��/�Xퟥ�k�JN	��C˔��(��P���c|��0�Nv��1�a�&�	� �>���B�˹d@��9'l&��R �5�48e��G4l��O�o�7W���A+�k����0�:�,��蕫�̈́��^�6��0�l(*s~��B�_Kު�/�*�ަ����!�?���&VX�4����z��C
WC�(F8P��[��o#�3�f_|Y��>���ADP�`':��l��\��co���������Fό�]���B��3a`.�8�u�U�g��e�,s.ƻ�, j@:t@߂�r\�e�[�:&��V`:�\a��l0Á�������r����gGs��ü��W���<�H�-Ҝ�$a�'?�H�"�ʄ�ZUS(s��j,�z+M�,+~�O��:�[U� �Q����J����ȝRQt�@�:�y��fȨ�[رeF��}9�i�:�b��[�*��ؘo
p��+7��=���il�;�1��iTa��o'�¤���4�X��h<��D�hģ�NSWx������RV�qt��4v�*b܂%;�N0	b������[�2��s�1��7��/�:3ɋ�#N,7vc>z�����7B��	��5 Sa"̜��' |M����y��ჰ��j��lf�{�(�b���=߳C����'�Y����90�Bͮ���<���JEb?��G@�!O�~�7������;Ժ����~@�v�;ͭ�������c$�^�׳H,��Ҏ�gz��=좣yuͽ��Ʈ��P���a]S��9����?m.�Zp��R��ǬX�T3΅�.7�e@�6S��\�zW�}��g �T [����
Ѐr��}�w�UT�W<�y���G�)�o��P���r�in[z��R�%�o�J�8���SE����4��h>oJ���v�#gQ�J��w�#����F.#Vu-��/t���žR�w,}M�m�܁���o�P���9�h�mH���;����s0"�X= !
.
�C8()��M���Ӓ�<12�l��D�m���M�=z�\()s�W)�b@#>ݩ����O���r�!�}�D�n��u��C���KM����>�/�#'d�Ỉ?SLȻ:��Rbj�_�O�Xu^����:�hދP�����7F�tMI�?o�HfF7���F�&�*4$��By�J�H���d�%?�����U��y��U����\Fɴ���Ѥ)�q-�o��)��#9V��$�г�3v����x��<����h��Wg�Y�Ak�P����L5��_�V��n�rv�K#'��;����z��	N5<����e��p7�G��DVݔ[�)?_9z]�)Am^b��|�g ����;C�Ō[R��qmH� R>1Z/ܗF�$�4��+�b�MfUa �t���r7�����s�kq��p���� ed�+���-�Me	KL��F��ԕ}&ϭW���4?;~h
�����n�+w�����2���s#���&\/�C��b�[��ol=?��=v�=Ý\1��S�Sy#¼\�{ۥrI����C���(��ڡcؿ�5Qܤ�
N���(/�U)nEM"�.1N��~���
��\�㲐����k�+!8~-�B1����((��V8"Z!0@A��������{����xp0�"yȝ��� W{�Sy�����>�<���s-\}��G��ڊ;6QPv�]���l�;Mq/b�{(�p]�@^�#���t��?U-�[����8�?���g0��)Jgf����KJ���J��3L��DLD���y	��g5�=�
�v��V>���fnn��Ӏ��ͧ�e�5����+��~rv����j5�D$ڎ���s���DH|T,)�����˟+��6	��-��9�Z�U�zuay� �!2{��{Y�ps���_Y\�,�B�YM^wN԰�8�4����N�ީ��r��F�:�[��
+k!��s���
v�4M�Qp:��"���۷�V뒁=���X!���@�ڋ�DM�\Ȓ^$����#�N�TYoO�M.'D[��A��U_��c���~�f���y�8�^��@�4�/�L-�tϒ��k��5����A�Ti�:�HYa���@�>U�ж�ue���C	�m�F���&ws����.X<Q���$�Ap��ov��WbԚ�䉧����4"����l*ڣC ������5��b2J��M-#:���\�$w�tMCԧ0�Q����������L��8�'�*�����>� Tp��x�����ԙ�BY�z0Z!�I?���z�(f# @[M������;��03�'�g� T�%μ��@�Z`�#�)P:�����^��)�c�m�����t��ŊM���Z��Fn���L�g���׶(�YOr�ʨ��~�ӕx��N����,x�������H�V�Аm�����!����S�k�}{όv�o�]k�dr]���*�fX'�;��n+r�;��1�Z�#Hp�<�:������V���i��~D�/$K�����+�y2�B�|���_Jb�h�j�[���1��G����z[�n����4��-��7 ��kMlh��.{x+#���g<�$�Կ�ZLx��*�A��ܡ-Pc��a�����&��L�ۂ �m���1[Ϲr.(Rp���n��X��e|���炡����HA�K �Gx���ߖ���a�F�[�`|˫q*�jP�T3 ^�	+�57����I�3��s( �ө�9�
���TdX�0OfHN �,�$�����r8�F&�s�6��9fz�ԌozS�������ۇQv���Z����E�{�d��)���t&ν��(��9�'� vǙ 6�j�������4䦗�o��0	
�ҋ��Ѥ�g9��v��?#��ϑ�
>b1�d�����kQ�	NqI�+c�)�_tbq�տU>sb'�B��ª@������>Z0�E�k�^��N���3m.��W�
��b+b5���Z��T�I=��$g�$�a���^:���̭��rZ��+`�ر��YF����Ti9�U_Ee�g�s�l�Iϡ�B��l�Z+���ߙi3o2]��:���(�q�]q�h[�4R����Q���/z@XB������!#���e;H�8�V�e�r;8|"���3d��`EVcq�dX�ٝ���ԍt��:�##ZQ�/��M�)���/'�xY��Tb-�C�,m�ޥo�����W�n�P�^��� �Z�����}n�m��7��wq�WWBlu9@Ģ� f"���m�6WD�m��B��zQ�G�z���m�m�X�����XF��?)\2��[:�{��l�Aw�ۊ/��`�A�k$��'%D6�ˊ��jAz��	Y��m��c֪C�5y�ǻ͊�1
���\=�"�B�`'Q$B���@mF�ۜ��"�)eL���j
������P�P�^�ݙ{��Ӆ+�+|x�#`> ߺ�\O�S���4�'O1���
�x��V��:���\�KKV���6^���x�"3���V��()��vI��EKr�Z�F#c8��	���[�W�9~�U06ǆ�7�o�h`p�!O��SQ�����;�QE"Q��E��y�ݐ�^�?����g��4�Z�����J	1�}ջ�G�5���JT�v �{(x����޽�C=����nI�3:eJ��t��-}?�:~�\���Nc3n2y|I2�\���F
�~�X�m�aؿm�{\�W�3〧<[����:o�(f3j��Il��l�*����H�ݻ{� B�>"f7�[�[)������Xy��{,P�Ǒ�Q-O>����)�ma�9���JL��
��@
�d�X*�s�+[�cS#�0�����H��ٛ�:D~�%v���KN�J�����{���"�|d��֞&Vq�o�#Ϋ�y�)����?=F,\���n��������%��s�F��C��ư�I�|���5�4���5j_��)��x���k�匆Ώ�.�٫/���n���Y�RF֊;�C�����ݫcĨ���85붇��gE�ذ��~ܑo�ϒ3��O|�V��4��6|���E2��,���|yc���|W���'�e�dGp{��5Ѐ�6��0���/{����ݍi�/��]O|������<����ﾜ��W�L�a��
<��э�	���ܒ��&�:��r�S�?i�����l��b(���%���ɓ���V�r�@�9/�"7�y0���(�h����7�h�q�g�"�G��4l\b,,-dTWg~��yQ�29H����yӏ^�4?SV��5��!4D�1��Z�-jz��]��>9%���������z����EY$7lڇb�c�q��\�>�Bmz���KYq�me\��h��� ��H
)z�O`���gyFA����0��1R��s�bʜ��uT�ڧ>Z���sH��G�cG��U�;�����*���K#�� 	8�i�mv�C�p�":=K �9 t��>>�F�@��V�{���=�ѥ�aN�q�a�/�բЋ}Cؚ-��K��-ib[��[��2�V��9Ğ[B�S�q��>XF� |��A��N���P
4��Knӡ�����8���� OPp	�&09�ontY�6��Í�����:o��<߳��.E�C� }Z~Es*i�V�@��
�U�%DT�q� ��*G�1yJ�����C�6d��[�r��2�:	��5�z��;�0�$��B�l������PՂpZS��1���W�������4�+y�{'U�&�} r`��sb�}Zz��3T�I>��T�ۓ=�s�f��)[��)/^�eT��"�e��ԕ�賅����!����ؽ��	�o�
B��&��2]���C)}��i�z
�]�o ��ݣ^��Sa��]�c��4&�'���Q�sQ1(6��v[�����#uݙMɶ�/M�>�2��Zϣ<�8�%.�W��bxN��݅_�Y?&ւ.�����H�7c���2(�&��
�q�CC�F4|:<חx�i����%t�?�Y���f@>��!7(2Q�]�w��5�K�_�t��k��\�����lq�A�`3��hȇ�F�/�R�I��ԖH��ה-����c#���[|���7��0w�DK�#�����w]�l���ASd��uW�-n��.��u�㽸�嫞
܄.��Kq����K�#�X�Lv�V���щ�(����<���}�~8T�����/)���wH&�G�� �����|��~��kv0�p��1k��\����� ��z+��Ò�_�YGG�!�ĺ֢pB��������8Յ.~��{�R);��T )���n�a��(w����7^�+(p"�߫�*wE����eY]��i!�K�	��x�>mQ����Vu�����?Ů8���tK+z�Q4��P���|x��=6������o9/f�����-~�d�L�7�"���/]>�<?ȍ8�/�1��@��`>�c�#�2a���	����вv����ҭ���Y[����O�%cJ�L�X<C���5�����c��������-}o��d�4M_����.��)�,��k�������=V9��$"�	ͭ��L~��R3���H5rL�v�y�A`FE�G���k�S�/��s^˵e]z|3�Fq_��w�K�m@�b�[g��Z�+;�9-�N�����>@"�&@�!�;�z�>A��3��Uh���=�o�fIF�� W�*e�N:4�BX,{jo�{���8�!�b*~X8�P%���/�������4�a��L��5�_6]0QOd�:n�WD��������H��!Bj�=i=�N;�'�9Mi����P�y�D媽��d�`�n"�
�>*����ڍf)���e%`;W��.y�]+�����Br��5�+e����İ����ǿ;��t�Ȼt�,�'e�I�>��X^xg3*�(m���
���s��I;����J�%�P�I�OEȰ�@���.=?jb%��5���Hx�����MK-(�"Y8��3cж�j�A-��:"����!��W��py�	�S[R�DB��D�lVw�\m�{��JL��&�V+�-f���a�	>eb������"$�=:�kDJǗ3%*���� sۿZ牔7��Z���,�`1x���N:�GR/��
| ;sv�,�>Go�L�o@���:�>��#�����]@>��FO6	:�$�k֗��%x���D!`�K���tv�k5±2�m<�����]8	�5K�E�y�V�FG�g��qA�B�4�vP���;J��Y;$��;����J���bv��'���X]Z��^/@^�F�W���1���~�[��C�=uĺ�=n*�������`'嚸���"����.�V�#�IMV�+!7��T��s��N���ؗ��[��n�A�f�ë2��T�灉_wi�0�7l�Ui}vw=�7]�y8PV��q���j�6!�hj-N�;���:!w*9T_��˧�u"J���3�R��� �Q�KR�|\v ��ְ� �w�:хx���F�eZ��ŏ�L5@��n�����f��IɌ�����Cvv�X̣�6d���m��F�*L���B��Z�Zd_�C��n#01��>S6�)W	gp��J�!�ŗ��*�=L$�p�\��T�;%I�W�S�&&�Mf����V06ߓ� �6�tϊn�v��$ja��&M�J˴�_�(����5��W*.?|��=plq��ꎻ������J�a W�6���
&���`c������C�@�cpnF�@�l1mQ��(�;#�r W��7X�]�d�Z���s����`���#���.������ێf�T�g/�W�9	ܵ����f'���ET��z�7V"z��AiQGչb� �j;I�m�.	_ކ��ЪY�mg�����Ѳ�N�ڿ&����>��!�ϗ z	�My#��Ϙ��j�J#sa���.l0��._aÐ/{����ee-�Bx��~(�/����n��+�r?�l���4����]�k���Hݏ���ΰ�qI/6�pX|DgSH&(�9�y}�[��a�'FD����cp�`HIn���� �]th�H�n�e�8^�7�"�.Q�wb*�j�+
��f��.��x!&�x~�����#����A�*���b���N��g,Gf�zWT���lQ��"���كA�[��H��md"��ŝ��Rq���) �[H}�;4p�T���p�V��Y��ћ���?m�7?�j��=!3��5U˕�t6K�K2΅��qNt/h����H��̝:��v�g]�J�peM*��Z��*AY.s��e�>�|-��`;�˱깛�Ip��9V�e��p,�~���n���͚bg:-u~�"���S� jp�NW^�WF�cʛ�b� �|�}�ؿS&E��S��:He���#��{�X"���ݸo�9N��2�β��΅�򡝑� �W��*m�cS I�Y��e����2ל�؉t���tZ]K̳Gj��Ղ
�t(�?,��!� tuXF)vq��(�~�XH9����?ez�U.$tB�+��u#>[�����Z����k���;m��J]i86�'����lz���-���r�N�6^�
�r�����~w�:����c=8����U,��T�~����D?Ǆz�ӏFR��ފOqY"��$���Ck7`����*ll"Q�`=�]voG�mWa�����K�::�1E�a�\�|�4�gc���PY`�n��?���rB�n��{}$�Q���vہ�g6��	�s����Wj�"�Q5����-��ėLV�t��Y,ޓ��}"�>_�~%�����3s����R��N������N�k�!���N5�	�ձS����.���'6���u�5WZ��BB��J�I|;�\��T��(���Lu��~^[W�g �~�.��7���<�b�P��oir�#1�@̝�!茡qݖ�Ks]�:���+�]�E@�g�{���z��H��Ⱦ|�4k����6�8�i���H؄����ԆY:s��~{'À���E"vȾ��2T	� z|�~�F��чi?'���px:N����َ+��f� �[�Ȏ���ج����Y�� K(JedƂ�[��������8��:=�A��?b�O#��‷�����/~�g\�nIm_�r�\���j������$A
�Ⱥ�������A��wgq)�g�} 4�I���~t�Ĺ�d�>'�]bs�Jj����Ɨ�},"���
e>�>���f��tR��,��j�RW��=�g�2G�c�w1�X�X',�q�&9���ku8�!L���~�(wor�� X{#6�L�j�b��p��-6�2o/��^�'��]��pQi��� ��G�ٍ�+���*�K�D�����Ϲ��N�x���_�/�)�2��~X\��Sǋ�fb ��4���نR��R���Ѽ�#��)��^�<~_mug}��(��-�f�+�V�$�V{]�=��Sf�D��Ix�O%0D�uW�HF������q��Cϒ�1E�DC�%_օR�Efs�%Y%�s�kqch̨a�DƘ�C��nQl��u�-@-%������:�^WNt$A�~��&ސS5�r�'ٮ����!�=7�����g�WJf�����{s)r�XH��}Dj�\ef�jǘ~�35�Zur���m�(ܙ��k���<��<$<w�%�Ԝ��L
)�H�=��������نn�Z�&�N�}O�'lBJ0}\r�֮|����E�"&�����ڢ&���v45�s0�g�e��_�r��<W	�L
��0a4���(R��r�'c