��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM�
Ɨ�j1�]�*7󨎯c<侤�ǩ�] �I\���2��i���8j�N��8�������]���`��)VM�����8AD'�R?�_s�ǉ���t9;M8"�-JƩ괟���ChZ)���G�:K��]R@E�q�K�~��C*{�y)#��n��5������G[r�y�� �Q���%16�wL��V�R�a2y�����9s�c�)����mu��V��m\�3��$�H�?��@��W�� �uJ�"wϾB���N���H\4<r <I��:`1���NdFÌ��\@w�ҽ�a侗i����@��G[�'^��J�*�3$nW�E�̆CZKÜ����x�(k�R��
:`b����e����C#Sq��e�\ZaM�w�2� �˯_C:�7m#4�0d��[��ю����0��=v+~����2q{s��u� ��p��!.ѓ����Qc�A�!o��m��ma�8$A���t���x.đ��#�]#�7lq�2N�;֔�J9�Wh'.���x~�ġQ�:w�>3cVNr��9�cH�"����F���2�[�ྺ���;��g{c�dl��e���Ղ5<����8`i����g��_���-_'��\�kπ��#g�+8H�/ר��H�ee|`�{+�69_+�& s]��]b�<��H `��(��%��au�g1뵒�+�?�6���4�B��s�dH��7ؑ��.�����=C�tی2ᢦ�8�s
Nf[)ъp��_�Y�>��� �4�>!,ɓ*��Y~�,dN�d}�5G *)햛�)9��X�7�ˋ乶j��KB  �?P^{�n"�Ҥ��No���f��x�!L$�~����(zܖD�ۧ?0im�v�,G}��է�|7���p�-~��!eŔ���0���m֑e�R���Ĉ�JA����{V�]�<Fl�z�4�$J�]�II�b��2�q�[H���?�sVI��{�=2RjR�7'�f�*c�R��W05.fpOZ1��:��y�����m�)<���h�=V�U�[�ӏ��@��j�A�S�O*o�����E��H�Hu�v��gw߻:׹��}kz�q��*	��v�&M0u��OVbu���٬���lN<j�і/t��𚋋A�|���Y.<�ĿmI��@��:�m̊�mb�p��A�f*?�ȵ+�w����A�+~6_����#����P��|���� ;_�j�ȘqN�r�5D�lɆ9r�[�1~ɘ[>#f8���8�4!��K+x�m�����&�B�����z#�l�u~��B<��{U8���wk���f����M`'�[\1C�#q'�e/�r(B�EQ̃�T�2��z�U&�Ỏ���?m��:��~BO VU���	xj����G�p���੪\J�܈�t�p��3ko)�^�-I]s����L�_
V��L��a��ހ�m�O������.S�J�X�pá���f������E� B�$M�Z�֭�v<��T�S�?n�W��Z�]�ν3��,��S>��z,̔$�E����l�oZ�d,�c �7�E������P4J{��d֑��X��u���nI��a�bI�G?�<�Lpb��h�[wc�J#� D�h;
)w7�_ `�0�`k�����_����qh^W~�}lޫ��-�ƴ��o3��?V :�
���6���g7)�U�:v}���`�6������_������d;U��d#�Mg:�I�V��5�� $_Pe�K��ܵ���fߒ�D}f�� ؛"�x����:�P��(H�
�-���L��G�5:���_�B�.b��
M�����.�QR����	ʏ��h��G�A� ߣ;��!W��+�����M̯��/yH�4����k�uc��:�(-���um+"6��cJ�j�s����*��mA�����V���ۧr-0�����e�B{�
���1_E��H�d�D��6�h	{
��#��&&�W���-�|��1�P�V���e^����W�a�-`���Ea��t�H������XYL%�og��8����l� �����`yx�ˣ�%��?5�}�/��`��j����3���uCo�?�n����s��r��J����]�k���l��Cdz������aH#oc���9��X����D��H��'8�����k����K�!�~�Ssy��i�G$�0���n4� c!�)�SD�(�`��a;�wz�s��^��կ�VGo�o�q�
>�¥��ţ�^�{	��T���1��q�tM7���A�U)� @��(�:�� ݪR�g#_��r����9+%��j��������]��������#1E�JӀ�7�n򤨱a���Q�)OAwNl�H�AEg�(I�D�<9���|q����=Ə�yە�ll'r�(*6Ҽ:���bז*&ޱ���ד)�T���s���e��m�Lߚ ��j+�+��Ų�~�!X���#�rf���}��,�@�hA�����y�`2�)XP�T�4���(,���>�O������ <;�?R���Y���l�l��\I��ꆳ-7�Z8󹸿��Ut�!������?�# ��&n�:/�Α�:��uŗ��>?�\��$Z��c�����m{����[��8�[�OمCG���!�^J5�tW�STyJw�֭��s:R/�`�� �v�ii�����)6��٤К�(h*q�L��}*Un�\t�V��o���� �D�h�z���T#�1����+�p��M�]nv4Ɯ��J�T�g�qP�3)� .�S3-��#����ݿ=1eOv4��r#�MF����Y�Q'��|����ٍߦ]M�L�)8���� m���Z�<���Qq�#���W���v+�J,,l"�N-��ؑSfʱ��0	�.�Oc��BWl{/>�wx�!ZX0��A��~��̂�椂V�R��6�s'��
��(� 
�RU:�x��=GQ�����O��Z��f{������8��I;� <�s��z?�+���wQ���f���q���V1h0Y��"2���U�J9z�êr�_$}���a��Q�ȿ�Ome0֎)���cv��\9��$��0������嫗h�V�Sc_�9/�5�p����>W�BSB��W��N��7�Ԓ
�jd
�|f8��&��{�$[s������!2U9q�h [�qܡ�}=�]�m��=����þ�;�����<04��b��`�Z�L�5�^S���
�7u������пG�+|�w;�럛�e�Y0.�0��b�.�\G�o�=���Q��?���	�+�
ʉ���t,<d���C��'�p��  f���U:�S '�[)��b�����.d��	��eiM��\ͩ&�_���x*�������+�����`\��#���������o���H.�u��ؾ4���a��Q�4\ns�s���v����g�3��-�y���X���/�x�#.�p\=�ϧ�����s��Sx�zM#�f�f6��bP�`���cO�� ��S��i�a�}!<�P�ZD�i윘훴

F'�j�E�GLLi����7>����%����0��ߌ`���)��(�B�:�V�/g�A��eYay�"���Gi�B�GK�-�1cn�K��\�S�r�\����bF���� ��;	=����v���P�zL��eq�B3�i��C�@����@��q+m#�:��
������rd�if!��BI*ȷ~V�&�F���飀���R��ܟ�{�HT��<X�2.������>��zp�?����@:�	Y�w�ұ]���:������Lx�(I�5�l����J?��.Q���:ol5N�.��h���(��$���ft�\�摥��:��e���0�(��\�&��L��t�}I��G�P�_��ٍR�[�'�~���:����4&M{27�2�}]j*���[t��v�_�&qGg�� �VM��V���-g���V�;����ѺMhr�^38���	zA��m��&7B>���C����9��+(���|q�v�Y�:yi�*�2��ǁ85o���A�ݤ{o[���.}]a�g�Uk6������/a}((��)E�� ��P-eOXTo�����	�,<Y������S��[-jd,�"����hb���/+ ��G��#|.�\?;�4��3k$)B��[��6V��u�梅8��-k�Zp̚�8�?��Ԛ���$;	$<�Y$i�4�0IM}D�jP{�X�"�y��ه�̓��'�B��cڅ���/�5i��E�_[�Br-%��C��T�wb�s�u��Gɤu��
�d!X^�������z~��x-Jz���H-�n�쟦j��Ů�`	�N/Q4w��u�\/������d�/��8�\`�����Y��0�<��yL��wy��]�-����D��ob,������(��m��.X��WRM�#%%h;��;����<Bkp����T��)�>U��{�Q1��{$�fSԄe����F���x��]v�����zf�]��JE�#I���`c����z���h�����F�9��b��p�T���>$EaR���=N�TW�ߞ!@kJ�T�죵���'0�]>�T���۫v�� !�|�V�n��G|��DR���Uy��j�f��a����-�T��
�tT�đ$���&t`��a�.4"��W~��E���e��� O��|�N���1/+��zV�?(2�����y��VTO�L����nD��;�h]Dⷴ3o��/�2� &IF{s��"Q�� ~�9 �_SA�$B���lD���"��Ε�W��X�Lx�a>�x+��#e�3�S��_9`f܊X��[�����dܼ��4?$�)z���1�"�].�Vs�0̔��4X:S�.�@�,�mwQkX��4�U=Aw g�.F�6��U8&�Q(�8�@\��Zk1��GLg���F��n���*�k���(2�	'�y�1�Ψ�m~�U��G,(�|78E��B�=6��k�g�uf=l��D(�&/"v��h�#�$��I�a(��Ţ�*=�o�'~�������3�K+!�1���G��������~���8��F�TJ�ŤU�I�k�[E��F?}@=����
�� �uөZ��WE�[�dQ)��XC�O{�����w$t}��_�̅��Q�
�>��BrӞ}�@�A�г��jN��,2ie���k+��S�N���}�>�5�)�~�g�h
����>��s+��g�N�2�`BAN���LG�>v�p���(Y��oJ�^L�$�Z�K"�;����$���5�z��Ö�v,� _a�L6�3B����E[ۡ;27�$ڥԀH�{��ubG���&�����Ŋ�.vZ�T����������@#�>x3�T�sc,��..:��}�l����E%�{�Ƚ�"���ʚ?:=u�=��,۔�|�md�dU;�	��c����Θ3�	�[I��8HU����bN��GZ�%�Q��>4_Z�y��n��6 �J��C���d}�
+C�*��L~	]�Ȁp<����9�6=7�"��,���'+*s�N6��x�؛ד��e۫M���Dt\D�^ob���W�����Y�ȹx����k�Ά��e��)WA/e_��w�n#��$����8ѹ�v}�?��K��<}#��Ɵ	����#�	�<d6̆.�;R�xYXt�п��ɞ^�����	���@��zt�+6/6������:�M"��y*���2[d�ƫ�������j n��tTY��tN�2�c����^S�R��Ydj�yF�4�����B6���WK������oT���"M�����*��=�H�Y|�Hب�����h�_���v�{4��d%Aؕ��H���C�|�����ٳI�8{����a�*�Qe�s�R�	Őq��J�7>i�>ߡ�F�䫛�S]��	����Z�Ĵ&<�TJ��z �R��e(tz�
4������B�":w�rS�m�2B�&��Y���n4:I+5�r��0Q��5�,�0\o��٤�wh�c�1�Hm�$wjB�����1H� X���������xɊ�	X���lkm�ɻ����������p����g� �`�n*����vS�Fu�՟{��cn��%���ڑ��>/�kf�w���C�� ��mǽ�x"�Lo&�$RG�PXe���lt�U���<���C`9j�]���^oY�$��U� ��R�2���	���dI��AMT���^Рפ�r?	��zOu�����~���� -IN����"�*��]�v����U�n�[Y��C��|�s�v� =9� ��L���}ޅ�'c�tS�rZtgi��XPN��?�*P(_b� ��ƞ>(�wBt�N�W��d&W�q�`(�hef$-)��	Z�g�~AF��yR{]2���J7�>�g/J�W�%"ĘA�%��4M�)��h%KT���om�.���^�\�z�OW#�����4e���v����<��z4y�QI��A�~rv*����Vf7�w��ݨ,M"
�/�I��n��DV�Y��(	�c'���"�� W3Q�ֈ�wR��?�xD��'��� %�K�9�6���2�r1IP���c2�� �ޣ�7�E@B�h(�W�$J���F{�8�%E@��R���[���L�{fƨ�8aE6Y�=,������� �[_��Tڦ�~����p�g��}�mi֍vK0�Zg�@����P���'���cPaV_�K=���x��{r�pm� r�bi�z}����I���Ë�p*�~Ny7>$��JĎ���4	�?��o,�C�� ��<��23�#ν��2v�$���*�t�;�	d�d����Wu���x/hD�߅�2��vZHF.v`����W pKn���Sݚ��s;��Gה�E8U���NAWPhR8�a�o��0m}p��)x��hϬA�w$����AS4�H^f}���Ǫ���4�~X�����"�J�����B�p#J��*���<)\zq�(���-������g#�˥��
f�mr���3�2˘��O�h��%�R2d�S࿛7�O��;������=��0�
+�}�I7�N_P�x�ŪK����Nn�|��
�}G_��z��CaRS^z��,�v�M찌7�hf3j�6�ƠJ��`'!,s��"�@�>�u���3�D�	xmi�r�`��,TĜ�K�����n�"��MA �Gw�^{���
Q����n�S�!_\�w�͸��/�	�V٣CgP��B�q+�__o���bZ��;�Q���l2��+tQ�����v^�nk��I�\ڿ8�ĩ�q��bސZyR}i�I�>�5��Fm�D8�vLoY�L��\Y��s�f�����7�������1������ b����mh��}�!��8�I��ؐcρfC��6)຅�w�W�A��:�
 �����
p����4�,�T��Љ��J����%uVgusnU�t*�w�;d�Sq��� �
�����Z�:���z=WgG�؉QX��YSTt͈N�5��3�Ե��T�)�E�i�I��rO'}C��)���Fֱ�6�J���(�T��jx��'��*�t��.�2��P���n��1��=dD��	�m7uRa�%<�[ׄ��t����V8�wL��ک<6��H�g��`�M��/�����IIP=��o���o'U"X$���`|͇P�����Ľ���V9�ۇf�ua��!*ޘ9pasF@��5�e5���t����,�X[<�
���� :�l%�3���ǆ�^'uo"t ��2��2v;yִ'$���a"��[X�B$�Ɯ�(��J�'��b��P�`4�5��Lr���3�W_��������n�R�*ZY܅�?ԌQ�I��o��
�Z�0�j�ng޽��� ��o��m+��S�����S�������8�=�=G�o�Ѷ� ��RIށzKD0���X,H�:H��*C�mc� F�����m�r��cIE��s(- 3���e\��b��8���5�KZ�0��5]QG�a�����M�#](�b�x��;m��>R̋�'�r�	��`u &�t
�Y���Rw�3W:��;��J�p�,� ��8T6�
�Rg��W�6m����	��Z>�@� .��Ք�ґ��V!P�4��G(H� "Ŝ�D>��V��!J"�>|�����+�3�Q�*�������6\�e��B}$�����˝��K�8�+�����6S?�%��k��z�"g���ȓ;,��]��쬚dm�+�=��8Ѽ�es���:i;�Pg�mL�5����.8���k		1a�R�,H6����H��硯A�<�4���}������8y�6H3S�ށ�.S���5��}Ž+�=`���3Z*q��X=�@�Ro�_��-��4"�[�_�`�a��A� ³�Ft��>'l� 5���~M����U�8 &�B�bQN�E�s�g����bK>ä��Epת���S�hRrVrH$Dqw�8d}������rC*o=�r9�gn�{��R���rr{�'t�m�n�b�C|��F�*�:���g�uV���e�i�~ls4��,�&���K����5�z�	h���R=�Tɉ/p�ӡ��V�&��Z_�<Q�B�a�����'~)�sv�1CŘؠЋ�k.f/;�.�*�T��-�F �U�c�y<�s~� � ���� �*_�"����z����J�������w>s�3'j�����wז._y�(	��H��RJ�1`�O� Թ���]D����)QNQ�y5'�8�x3v��:��&Lg����\�r�Oe�U=W<��GS=��l�r7&�E��IV����b'��;���y���T˴��p�Tn��fm7lW�K�a��Z�M1�ӵ񥻿X���@��P��
~F�6�pp#z���:�@%:J���V�E�H�i�J���7f�`�q1���+V��(�}�'_Y�K���xgSv�lH�e�����e�pA�D�z�,�m���%N�P�ݘ�/�Ň���� '��1��G�֤�<2
�?���`<�泙��s��V�S	ucY��*��#GD���J�?�$sK�A�	���-�=��S�#xm�K��|O�lԒ_����:���=[�f�� ���`u�Y�ҁ��S5b�>��D��?sc����n�uf��}}�Ҍ!\<�A��:w�gT��i�eUźmP�����]OŻ($���.� ��5v�hB�wE���7��M�3���2��}n�_��v�R��⥰�s�~$2�㚚�˳��݅������}���l�����,�
�p��(`����x�ᩣ :8J�8�G�9�Gn���Jv�!�9���
H����mE���Ş����K�ݴ����\3K~�F�%z)\��ȿ�����[g����%
A[���14�i�wx�� tu�v�%�V@�6�[�?�e�^8�CU"\���G
���d���!+�`^�pvt��f�J�^���bg������/Y1f��Ĳ�P�Ē��l�q�6�'�_%�P��L�b�8�BF��2P��'j��wj^q���-r��X V�cM��l���v�n6!��w�G�7>�)�m�8� ��g�n�_�[���a�YX*G���~�aW,�n��k�y��*��j]�u�\j�U{G�_Q����Ce�[��EJQd�*=;2���ν�1gc/��2@��HX�pڡ��e�)�S��`cc��:�BƑ�2���h�(ύ�v��P���G@2Y*v��7���E����$Qy�2#��'>�Н�2 53L�9��������&ʁc��*J���Gz��ѮN��ߜ�(����oS����L'����W��WiAJ���lU�n�צ�&���L1B�[@�\�&�X�>?o0���jhx��yOը��-��-X�*�둸e��kiG�:wK~�2-P�������@�XlT#Į~��E�� ���j_�ZK�y�t�����K<&�#���"L��+���p(��i���/"P�����}c�8��꘾��2��;̛���Ct�����PCҨ:'է�2�-^���R���G�0��#CQ�P��q�6I�����Ih��E�@�� �t5�� }���3�2$��&=�.�<<!.0�+��5������U���.���A@X�k=��m�D0�kUY�� qGθ��f"��𾕻R���A����-��U�����#�sv�`.(Sv��ް�f�s�@�q�I��S�p �r� �ų�8#�䎓D�e����d�+}e��W�/����ԕ�"��-���p���DSC�3��(U|��