��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�ֶ�3�4q����}��{x~�� s{��TFҫ��J�^���n�AH��k���s��#_�;�b�O�u�|�������֨��#�:�b�\77���}T�I���kX�ի@�6���12()�|{J�4�&"�}M3���_���mD�ی�`[�K1=%"�T�3����j�;&���%l�`��:��zAjG�����.{��X%Q�Ͳ|)�K=N|�lw���XP�4�@]��D�����2b��"u��eg���J�u�%�4�^��2V|�]j^���
,�9�O�1�`.�2B��9��5?r��7����։rmf��퍱��CP�m]��}���&Cw9Z]����u0J UO��t�i����i�O۱/g��@iJ���2[�LC�(�$sZƌ i�jw�ҡ���[�c�"�Qjw�cK�َ.�$�]ɒ�\N{?��/|��� �C��X�?8c>B1����QO�K�6��u��������ur��}.�O
�������آQ��~�	�@nFJw<{F
�dU�|���(����l	�
H�0�utQ!CuR
���]�d����䣙z���?�š����*��Z�J��ISjK'��'�eӞ㴪������ʎ�3�>� �v�}�W��j��[>��peu��^�l���3�iIT�,�U�>�#�n(){Cǚ/3������ط�	�
׈��BSK�$�F�_&� ڷ��nX�1�0(RA�@]�R�[�l{O��� _�����~G��bx_t���H�@�,N8�@W��O@$שU�O6���Xࢠ��9��?��{i}/-ҍe��dΔ��9^��k<�Q�HZ�v��e�!ը�˘_<��?a��9�|�1��|&{'=j8��\�,��0U��jP��q��@�Cߊ�|i��ِn*�I( IK���3U[H�KO��c B҆���}z �Q7��
$-g���3��N<v�]b����{�l�JgJ���j� 꼎��-g
�����9��Ey~�$(H�����zl��$�Ԁ�0�Č�#t�vH�7���[@c-L2Q��N��UIx�u�S�χM�>ޅ�{�yDn@]�dX�8M\s##t�t)P_;.�/A.X<w{+#!����v�)Sr02 �~\��vz"�thD�Fj�v2%>.��#�O��E��/?�����?K�=J3�����L`8]�n��r���Ѻ��wh���r!�-�~�ث�1��6|�U��s��lAGz��5�P�٢g���)1ͺ����2���(���]v��������͓°	<�(�����c���@G��uhS��\���0R�h����ܲ�B�a��؏���i3��0b!���nH�7�Bd{H��j�%y�Wi*��s'h��6a0�V��,ϐ�aZ�@Y�.\�'�F�[�x��˺��K\��l�f&\�6��������E=,��H���R"�Y�lby��U�KD�0a����N�l���r�NN��a��8Kv���dl�E��_3�$As�?��+!yI���RvLs!ϑs�B�� Aj�k&X��e��Q�� �9f�EH@���[���1
 �ݔQ�A�� �0_���<�ئy��m��VVy�Ly^��!�F��F������7 ��G^	��&�W��+�܉A�	�%Cm�Šea�ﴥU�=���(O�M%^����UL}�V/"ޥ�R��[ߝ�~Z<LF�F "}��Ⅷ��y'9C�`Of_[�Q�Ux{e��[��I08e����+�M����9P*^�,T�>�\v�j[d@8)�Rݩ-2��z�%3��w�Ѐ�0	�U�]{�n��g$.���Q����^�?��ܚ5O������$V��\���cGڃAv�j(��CS��+v��%��f$���J�J����{�����7�	0����i��WИ?�.]yE���X��#~��X�&V"��x�א
�l��^,}���^��;ޯK�.E��B���d1��q1e5�l�	��䝹�1dRÝ�3�0@��~6�n�j���=��-��Jj��RO��
SR@�'�6�c�J�\>�LD�% }�����p����]R^�t�N���P�<0����;mc��w��1���/2̅��^_ �#g�}������z����a%������c�`>�?�5H�	��-�*������?@�(k;�k�yx'Ãp�M�1\�]�	�hK��o�Bq|��\
d���N���p��0��?�9h�;����9F�ڶ:$�;!���$���n꾢2�]��\�P���ɛ�(%���l+H��k$t�L��qc�����#�b�`&�pA�~{~��=��_=m���5ׂt�?o��h�IΈ�׉�sd�H{&ZyUr�����,�����&����-(��A�3nd���7�.�����F)�B�=�܊IZ���ĺ��<n0Aޅ�5����j"��\�_���!)tW�#+��N\����ҡ���W�=p�;��ru�w���o��<����g� ����B-�h#�BM��ŴY>K Wiz�j>��o5�:���sf�nM� _]F�
�����d��U�;?�(�����ntΎ�[�+rܙ5�EǕҥ�V��N&y��ݏ��/��hz��4���O\V�0H(���8�"\���D7(u�����c��q
����i��0w��fG�8=m�b�����ŽDs�7�����3$�u���o������U_��H�l�q hu�Xش5��π�HcPa�eÇ��e-�>�R�sЊ�k��*�.��w��Bm�K��B���t�?_L�&��N�#�7�Z�縪{8��$z�Wʏ9��!o�c�3��� �ֹ��qs��D��b�g�!�`��Q ��C��(<C�B�e����]#]�*�l7}��@:(Q��X��A���<�^��G2��6��ݏ��4i�G�l��+���c��7�
��`v�)��ۓ�f=�te���Ez��K n��9����}�y��.���m��PY��l��R��])���!	[�_嶋1E!��%N_�~���n�T�Ck�}21ۢ��26�$�5���)�-!�oǩƞH��A�ڕ��eT���ů_&o��'ڐ0AH����o�I����,��H�V�%)���t�q~���
��Y��eM���>w�f��5=eG�r���:S�<�RKc8�_%���A:S��^�"�Z<��t;Xx�rs_]"a��ћr�=���j�[a�bcO���$���Z�H���[2>�f�<��j1߱b��"9^�A$�By��)G��zp��Ttͱzf�4�U��W��n��2�sb�Vn��Xu���4��9�<����g_׹�\M�yH>��v)�k�1��6n�'�jK5��u��y#[kK ~��Hޟ�.�uV�x�|��t��ϼ�����(8�?ϼuY�
)ԣ�ޟ�H��%Q{Z��q�w�,`�2ݰ�8μ���JQ�-=�l�o:�d1f���Es�VO�Js�E��OS�2C�KWӔ�nSqQ�ˋOW	"��m����vu�q<�� Tܒ� [I!��3)9#���!��t���	�~Q?B���í��D�͈?*Mx����k��5e�p�.�H���2��_|����.ș�vI:�KO��w��Op�b��T��j��D9+h��[/��J'^F��c�5�.6�O0�9�81�i�Y
���\�2Owӿ��z�Y�c���(^5������u�\�f
���z|���ܕ�lye�/+,��k��*ê���1�{�!(h� ��(����Ffo�Y�a#rz�Ƽ=�����K�}8�Np�)u���]�sC�~~x��b�Ж�
��]}�͌n^mN?����^0J�v�]�-��Q�f	��RO@�ͫ����;��ZW���Ri�Q��-:��/�wqA��gx,%I��]U�*�޷���"�t�:M����3x��|�h��BE�J,BP~�}�v_��>2`��jG+]""k6�Ҩ���dO�a)�>��Jp�	}��~����_!~�1ki~�|{����˛圈	%xR:m-�F?��]`,.� ��%�6sdm�Z�1�Q���)�مI{.��LM{��`p���׷�����Y����O�D<���@�?�E]N���*�����[wX���L�w��ЖNN����CQz2X���J�0m٤�Ŀ "�[�����j���)ӂ�����a/H�&$�߈�
Tl�?د2VؿC������/BlU"X��`ԝ7���>�3��l�ye�$'��<* Z����&��� ���{�C[n�<Zc�0+A��a�a��J�|����u��o<a�H$����B���d��kYB�{()3��*꘥w�}�&\�}L|1(mTe�+ +�5y�'ш���
GSk(�j���9zQ~069j|(n�����Z&K|(�ߙp��9nʜn?ɠʄ��uJ���=ϒ����'��>������b8��C�c¹����I ��Ԣ�H�	|Ay���-�M��U���!?V �]�O/�;�3 ��>�Cz%4Ax���q��l&�ڙ&��1�(�N&��7Sv�m�� ����~c
�|�`��^�\���2�\t�BB���j�����7^�6�6_:PZ��I�F�X����L�����f��'T���Y��})1�a��bn��PS��{*N�8X�h"���Ĵ�/@X��*�n�7�]x�}X�	���o��D�p�n�գl���!5O��{����{d�	��ͱ�ᠳ.O��,:��t`���= �>E���{�G�uP�6��h�5xY\a��R���5��/5�p���De8��9��{��!K��;oٝ�+�sE�,�z,b��j�X* �Ny�\+�ܧ4�(
�����1��6������5�S�gt}j@X/����i�:\�C~�
�3��͎ȯ!�/<��#��B���c�u�Lb#Œ�K�<QKA���� A�)���0q���=��W6�ZI�$~`�2@y,���ɮ�,dXT�Q�ܑ`x�6ȱ�	Qx����3�c4h���-�l�)hIM �пUX�>�Ձ�Ѥ��p�K�i^3U���f�|�o��|�7Z��bs��ߡ�~c1߫�C=>d���W�vE�%Y��~�!b�%7Ӣ ��a;F�������)Bj���x+�:��7cR^�*��U�������(I��4����w�{�,z�
�F0���	�kX��O���BD!�!;�ف*����EDIm0~�x]�k�D�l�2���=��5����K�^�5�9��q�[�8��C��l��!��'S��j�#Q�޷T˝ZQ��4�"��I�dg��"߸L��+!��p��H}�w6N���h�:c���*�W�H�^��{�Ĉ+����d�V���랧˃2��@�8���b7�'��$���6����5��7iQ��T��*���fw����ȵB�JxQv���<S��y&$sJZ�p6�%�[��uྲO����؇�T��i�VWN�sƓ�:b�Gۈ�%jSd�1g��dD�mI��vnR���$��#M�d���t��Ɂ8�S�`��z�9�ܾ��L��A��I��ڏ����1tY� D����߃�ƽ��Hz���<b���vo�b��ڌ�$�#J_H��-�~�Dl*.r=S����Ca�]F?M?�|JIx��\@?D��p�g�$��d�i:�ks ������1�[Sɼ"�x�yv�JZ�s`�q���c�P����YZ[׆��	�7�(*)��h�a��hۧ���zLo9����}	m�-�0L����2���c9�=j�"qh�ڊ(�]��-?F�i�ED���>�']� �*�trhF,�g��$$2.ʧ��ac,��� y3��C��y)vp �a�m���|P�̦�f�R�05���GM^@�C���6k7��B$�� ��� �Ny���jG�����=S��J�P�e��:�\�(�c��M����2��/F�c,_r�0���8:t�W���D�g�U����}�.�0��.�P��Kg�M"�����k���lLC�PN'�{<P�ǁO�1Ï��#�8��G�^W��KLb�Afy���mCc�[������R@W4�dI���|5������f�����L:��q罙[!�<3�#�jgk1�3Hp9iq[���7ݽ��.�3�0�qX��1h�i����r>�0�D��)�BO��E�V�P�Wam��eB%��xK4F��S����
��+���#q���d�P����'K<wDs<沦��&CN�ڠbX��.1�90E
��]#W�ɩ�-��9�7JT�T�]�xd%"Bh�olcB�^�ߦƉ�~�?]��Q�s�#�wq�=��p7dyٝ����Y�Y�Y@���1'/�+^R��U�ٌ�����It@<���;t�|���F7�2��yۀbL�\�"�E�֭���S��O�7��b�Y��ǁP�Պ@@�P^ޏV�����B<چ����Y�J<�I��6���(7�P���U|�S\�+�U��^�=U��ی�L�"�^�S�n5�(��k.q�M�o�8A�֤2�W%(ˢ�Z�P���.�^{f"0e�X\ջ��,�񯘰��r��9��_���!�3��~VY�U�
핆�ץ������bŒhWV��q��1c��8�2l�F�R[���BKm�-=g�2Q�$�&�g�jW'c4WmR��Y1�`*��썮O~��fO5/���^F��_���T܌V�W;�t׋�V���~+#fN�hv8 b��'8&����?� �%�*6D�>nc2�^�B�彭T���${���Ք �N�e3|��1{�:����hr�+��zB�|4֬&�/�r�/�@	��z˓Uls��D����P0��KU�>6\jY�͔��W�X2��W�Q��ґL���
Z0_��.GE$�a"d�QѠc���i����\�+V�8Q荜�vP!$����Mu"y���?�ưt�`S��Fi����;�J�%1��Ό��H%	��_�%���ꓫ�	����U��:�����Ln����K�k���Y���[�=�	e--��+��ldv�o(�8J�9J�H1f��`Zq,��VuɎ����ݶ�Dm��م� ��6U��=��^o�ep��4���l��NƹV��I0}�$]�;�P�LE%L�@�֛����A�X%'�ԪU�)/�L��9��Vd�މֆ��'Ղ����Fba\�j�9��5V�Lև�ĕ��r��[%3�zBK�.���yM��*�W:T;���Y�b���?��8qdFq@Y5�����5��[�X=<�Y�4{�$�0�,XM�2qC��k�g*�2�m��5)G��Q
�AH�j�&PP��C��#3�]��b@��d���^�x���e��&�b��*�-g�a�R_IVN}�Q����qӏK"��MY=�G����ဵ�v��@W��P/�s��|�(���D��50>ǲ���<�|���Dmo��I|t,hE�Q�f� qk;��Ϭ�ɲYk9M��m��a�����,��q
�RZ�«C�l��y��� �e�i�3�;�<G�S���Qd �N\g։ʢ��l�X��
��=o%`��P��w��^퉄<��_�LR�,1�W?�yY����
����2?�p�2��u��Q��//��|�	��Y�a���[J	�G�Gw�߬�ܐ�ӄ7�!�&9_��7"��^���n
�]|�,8��q#����I��d�sWiLMMF[���y5�:�|��;E��u���(�@_~M|VQ�9��qz&���P\>o��詖��ϫ��Ao��d��^hMwGV��E�ڝ2�����.�;����X/�9��0M���S��� H��d=w�*Ua��:F�~D}#�C��S=_���{'Ot�b��ˇ�8��H
����(Ν��H:�<(���& ��\Qw�)�T���.�����(�BL�� n|=���No��z�YA��E�g��g�*���Ɯd������&u�u�r�6k#wn|�wn'�;�����3��%�P�>eI�4'^���c��DgUo����x���[	皷�3���8IAL#�9���c��C�������a��'-; @>vٛ�C鏐�`C8��H�1c!���:�3���|}�H�f˧�"SJrg�
M�o�w^�E��I�9�g)�.=&���IQƓ��&k}[�s�0��(9�§wVsb��-!W�x��`�-��?7��1ȪQ�9Cd�}A?�� )g5svO�1��$D��\52Ɍa�pr��ԍif�o������ԛK�f���X�u8���Gֶ�e�I���*�M/Z}�e�a��x�E���!վÿ�H�/ �ٯ@���dA㐆��n̏�k�z�#����O)��g�V���!yz�R�f�N6�N`�����y�� &y���M~]�p8P���Kw�����X��Q�F'
D�9U�;�z���5�HZP�@SE�%U'���h�X�z�R�V�.����2��|<��4ˊ>^������l�b�x�s�̡�g�#9� �=�����������%N��p���0Z���������vdff�G����B������~�C��Z��;&l���p�L�v�kҚlš8�0O\7z�.[^e�枴k�J����-�D�8�ф��N��<�N}A�N5��!�L �-WɎ�$ܩUğ��+���m7�I�Ħ�)�hF��E���pGDe�%���݄4EQ:��>�_N)���h_/L�wEv|T
���ט/��s�mc ���#�8;x(#��Sӫ�{�V��l\*�N�da���ġ��#�,P"a�~!��l΍SA������WW*Yh�2�Xr��40�D�P�� b72�A����SE]�^5�S��4Q��WQÔ|^��#���/�O7W�j{eٟv�u���C����>��'��?{����q��4����� ��6�I��s���fH��T�k����\��p�F�T8�ĮtN	�8��4��ף��>�hs�+�s��)��\���p��t<X!�r�$��
�[Տ4����
����g�R��s�O�ʩQ�}6Aؐ_�q�h����ˏ�������:N��"��|�c"�P�|gl]��O.�7����4�3��# 0���U)^'Y��<�U5bi��^�D�uyz�Q~r�����CG�%KB~kN/ �kMz��G2s�/_p�&����J (Y�W>�`AA��G[.��ʅ��EO���H����.	*$��?�����ρ_2��k�eF�*�W��@×����7k{��� �\C�	��a�� �P�6/1�N��·�����.�����&�z>'�6�υK��)`��3�Z|�t�zg�2j�ۇ���k�S��nT�(t�? ������^�[���B�!�du���')�ZOo������n}/|co�ρhm"��� �v�&�R~#���r��:�`�E;p���-�I�3�`]�C���5�,�Ԝ���X4��'�����?4l��oA��3�ɩ6����`~��K��zQ2����Ԗ����́�,��aK�'����0&Jt�[�R�KZ[�p���l�o�2��d�i��"��IY,�<���,Z�KvW����>Ȇ{��XM�YD��P����+�����la
Q*�L��ȿ�(�|k-k�.~���k>|�������2���J�(x#}(o�i`���R�?����bC�j��#L�$7Ga�O1���0�x�"&�O�gt>nз�96��O�[�U��vP��E ��<6�)�YY\�S��"W4���|x�	�Y�!;O���QE%�c2��L�)��%�S8�׭�gS��=8H��4Qg׾Z2���3���� e���P�@^��g��7�N�D�x4NY�����OS����	�e�M��xo�*2�d*��Bf"��Q����O�_8����نdy�p.sU~!���ё1��$�,��������ۧ:�d��^��iѡ�VK��g�i�JzO�D!$el0�.�|<��k���9��-З�	zX���㫻�!��W�$�1)��CԳ�3b��$#��X�I��6)|6�k�Dy��o{�A��O	�~��F�ϓ
���u��aET��dn�9,�C	X�Y�me�i��qϏ�Q��Kb�*~��T啠�Uh���5��9*�({r�Of�m�>ٞ����>� f0�/��]_q�%��mwFs "\K k^�7/
V�����d�)c#� ��5�9�TV�S������0O�v<��Lt�Ce,�4�iȘf�-a%�*kj�}_[̚���p���Lc�[�:���g��7S@���mY�x��M0緊ZU,O��"d�&�\';O�ڳG��d�wׇ�T�BpG48BJ6w,x��@~N�3Й��c��p�p5��5�Fl_٨�]D�4$���-�lqg�k�#�����9�t5[�W̢��紅���L���F���0rn�.�!�/R �<���Z
sǦ�b<�i����ݎ8���ՀE�WE�#�o�̏҇W� ��o�}'P�)��O_b����')�MoV���7����![x���n;�a�z���2��#>_%���c����RY�|��R�a�鎄$*4�N#{ 56̪�P��ֶ���!	W%I����q�/@L>�i�	.L�#)�6D�9��@⇙��D2?���$���䋦�Z�9݁����@�h�<E�0]�1.�etpnϯlv�0%% ��;�h!#J�Y.�R��\TcF������,��.�'��g(䤽�m�5�����M�/)yd[ }���	�U�y��m�`���̌�6Q&��1��Gesg!����$ڐ��K-�=͛�vg�'��}EhL��"�X�W-qU.C[\�u��'v���W2�e�F��F9@�5񺬗�Ġz�VD�k����*u^K���d6�^И������,��i8��� q���tI\��)1G�0k��w������4���! Ъ���ޏ������"��x�%o-?�]�"j3A�����y���o���R%����bD�~�#�_Žx���
�ߒ��� ��`�73R��&#q�@�nKL��ê��2u�ʖX	Jbq3��0�m��%��?���c�:����r��U�ߩ��ƗREO�p�qPv#�Nӵ�Y��[����7���t�ҋ*�l	���xl�2� �x�'A.�1��@*��i�[�	�Q��P��+-�$�B�6q^Y�漇�G���]�y�ʧ��HJĹ�+v����n�?-��m��ۂ��%�b=c��Vp�n�|co��7o��.d���F�ӭ{zƇe�=�����G�ŵ~�'�2����%r��^�� H���������o����B�)]��%E�nϟ���4�^��*G�=�|�jn|�Ars+Qh��d(v�[V��p�r�]�k���-��	�8���SML=��jTr��%QD�1�ҭ�����n�Q����ݛ?#�'�Mh���=�:l�^�8?�*���i���/ÅϠ������\�ة�3 �{�_Έ��ù�� M��z�$
��t3Ð�4�|Gƅ$fɿ���as�UӺ|j,�6�UU�>�)���<��(i�3��*JG���#�̖A��g_ZR�㧅jm`Zzǒ�t2zO<�^d|�rIR�p�	0a2�&�W;������(
��ݧ����e������n^U���"�^�&W��+�`/p�� �k9ug��f��r�_�&��Fl	�A �����E�������;��	�б��+`�:���f�w��sИ!~���Gw��L�o��n{�� ED��~��!L�I���轄���5k=Z�>G/�+��GFܼ�<�Y�`F�t���nH#�a�-cJ|��C
8ܢ9�H͆�z*���[W�ȥ�z�%~UiZpQ%��QG��X�7���g��;:�)�Z�O�-\~�9��[̮i�e\լ�+jq���O�{���,%�?>�M�^���7��0���p�;b3 �.E&�0�Y�4�M�M����Iҳ��~�8%�=�v�����@2/�*��c��x��+ѧ\S!(�Y��Ϫ����LU�U���9bD[�ǵH{��m��I��-���*UH�Q�d'/�͟����.%aЩ�m�ޱ6��@{���P<��Q��Xh��WP��x�S���Mj)D�O��z��,p7�hg���:�V��B�qPr�T�druIb�~B):�v�j�p���Q�d�M�x��|F���~�<�>&�OT��*��Q�b�T�(����<=[o8���B+{� ������L��~����w�*��ԭ��Z❖=�R�O�ys�*�nX�@��GNJݼٔ�. �	�Ϣ./�-���m��S�F6�� ��}�iA$$Z��d�T�o�3�U�r�#���BbcA6�_�X0ب���I-DO�j]�>Q�`9ЌU5�H;ݗ.o�'`ö��,�8���*�=[�h��b+:�zrLo���݂�w]����=���Wg�6 �ib�mV���I�h�wb�d��C�'����?x �?��d�>wCg��Z�^�
��+	�����
�a� ���(�߉fLX�x�C�2R��Ԍ�m�T��0g�v�W�~��ws����Ù���ne�7�Br{�aH��&t����TKpS�߱��-�� ���S,¿Q�
�ʗ�M�"�@w:���-����A���1(�C��nS F�\S|	W��.RR�L�
~�5~�Xt!3�g"9�b�.��'���$F��@��Vb��ZJq	�O��3�p!}c�6��h�W}qS��Gз�*𡮼�-����cP�q<#l}CqM����mQ�N�׫��#�-�1ጪ�?�����u8�w�Lܼz:	Xu,���fE��>��JVѼ.z�e.?�(w~�4�5�5X���C���<���n�!��g�y�7��~��n��Sp
�4��t�i7z'r�M�Ϣ�)W��b?�R+�_���h��x��!<�!��ð�S�ڎc�^�	�aP[�
]]�i1�x�>��6QE�K+X��������e��P�!�$n3���`7W�#
��'��� ��:�zv��3��[̣��,sR��ۢo�A�����~��uA�+ 6�fE�~ۗ�)�Y��c��y���y9� �e}�����y}�l�� W_).}���ꌁ]GR'}�,3eǼT& uw�e@eR���8ݫ��p�Jr�C+i�k�7R�S��>,bࠩ�m������7�B���~���H��οR��no$)��)�,$��A}Ѷ����Y�ST/C�k=y�զ.�@�.�TX���ˈt��<�Pˇ�1�A
c#�i�����?x4�Lc��Z��������õ���1��R*���Ø�i�B���3��%���܉6��#O���޻C�Gr	{QA�R�S�D�N8��ٝ�Ey�.{�0`�7�P��F�m9mpl6IM��DݍY�f����:�����8�.�p@��B!?b\,���&ua1ֺaW�N�"����lk33�9D�%��hVZ,b�ѵS��g��q����0����Z���՛sC�_{}�5�n�1̀���ֆ�����4�K@�x�0��::ℱѸ#���*��
�þ8���I����ʀ����N��Ob<��	�'�8��I%������q,�DP�I0P�DIR���c�� ��i�	�m���%�Je5[�z���.B���|�����T�[��f 45 �=K;�`.E|�/�6��+�jv�K�GI��F͐�T<�Lr������w|�a�U�&��ǧ�5����z_zn��P��w���+�L!*)҄��U�l����
;�5���b?����kW���o��3$3Z��e`�	���H!;V$�vY0�:qd>ɩvJ�A�C�됤�
e��20��� n��.�.���8j�)��;��N�P��`nB����.����H#�p_$?�i�qk�j"��
|�jVI6����7���!��P\)hy�+����s��bS�́+��]�����E,�ڛ��RA��U�^��턽��Da�R�Y��d%_?(bHun���������$��rJe���
1�I�,���+P2�3��N�d�s�T���#P�)jZ��^M�=�\�M$��)�D>�o��,�����Y�!M�����Z4�F��z
[���1�R�-�%vB��0��r����|�X����'�V�p�j׭��c�%
��9�J���Ґ�����(�s�T���TH"	dV���⥉�0���H�sٱY ����p"�:A����ݫ�&�V|d������c�p޷x
;1s=͟s�rL�k?�e��0�I���*WF����Θ����k<4�������A��r߫��3��{)�x�:�����e�%�:�������8N��m��"�8�!L4$�"�Ψ=�{���=�M��ƶ��C@��ן���C_�ǿ�0�k��s.N����;���;�Nn��q4��ʲ";@t|�}9���z+ڼ����^�2�w����G��==�f�>�/�P�����s��i��)�d�z%`_���xh��9��xI�y��L�=�>p�Siq1�+�Z��1������t-�`5�%^���W��-�iǟV� ���t�ܣo��n�c{�S�ў��6�WzeB%�U~�*4�T�T�`�o��:�lh�"YԞ�ʋ�P����6����A8����t�a���H7L�=\�_ �ʭ��x��ˮ��gg�<���r0>ea���ߗz�<�Xc���*z�_��tV���+�9%�r�G��&�O��6��cP@{ p�d�"0�;>�����|2{�_ٜ��0���/����gy�7�W�#j��)��Tn��{�OȒȐujҜ�ť���`����<�"В��Z��(�"�#\�1���dɏ�^M��8����8�:������Q  �݀�i=�OO6��:�����o��,D�CV&k�x���ohJ�|
������
�|(;@@륬�B�/-�XDJ2ob����G���h�\�����f�K�nv�7jbp�#�ǩ��!�Q4L�98.�>N�&��O@Ï���a�9%g? �U�����[I�ѧW���Sg��F�^%�6��>�*��,�EX�&���t�����ơ��*���|�>JJ4 �栉�G�W~BC����p��"�q��������4�.2	9f���`'�1f&c�<޻�gm�N����/@���p����1����8�5��N%Mn5isC�2��:�Ŷ��mj�<�o��ٙO�>9G$ϛ�)�bi3��R��[��Psy>��o<��i��$���:|��Ef�7ypW�RX��ז�{\g]��9����og�N_[��ţ0!��f{��@oa��#��%����7L�R��mtPछ�3r���E�')E��R?-h��7�8�.��f�]mČӌxa�  �G�L4�<�Wy�@�dP����S
��\6��RCңc�>٠�� �Tv���1��#�T
��U�k��ɝ�ŗ�I)UE�D�^@"����7��-1��D6���m�ߟh҆��}�LnW1z������i)�5uz��yf\c� 㵲ec Z&�����"Ns�Za���Ĉ�dAU�$����pzۋ���}�-_ux�	��6PF�_Y�{�mg]R���6	$N򠗾M&����Tɓ�5���ڛz�I�;Z=P��T��۩�g)	�b�T\%-�k;���e�W��欦5Ll�ݡ�.�����6���hq�=���;`�a˲��kn$�x�f��w~v7NL��r�#D����Y�}@�oK�*�Q��_���ғ�'#���zpYtzku�	����S����U�B��ȉ5񶒴�w��:.^8d^+V"ː�΂��|���y�ϳZ��bE$Vɜ�%ќk���\TƐ��ͬ�L��w���~��܇�J)�HJ�E7�V�*6�&���ҳ�Ma%}�{d�jy�"����S�Nn� K}�_���iJy�2P��^��)��th�΄�<岤-._�+�\������Z�����/V�{T��E�yɑ�����Lb�L���l����c�'\������i�UA�*���8gw�:Sm�):��k�QYQ�y׭\I��j*_��iL]���F"Z����=~Vu�"�6���S����G��U��075G�f�9<��ԭD*�~�宍�<T��E�a�F�����2�sы��2Φ0@