��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK��N��.�) �A	Z�y�9�Z&����X���ד�/�0 P�u�����?,�;�b)ޤ9{�ӆ��;J_�x�Q�u`�,Ȃ�- ����ڵ>,>V��s���ʢ�3���"�&��wH�
x�6zzd ��N��J��k>��q�H��&�'܍��q�	N����(~ b��p��̕�[�	�o��_3f�X�{�x.}�ap,���-7�&�'I)��5Do^s͑5#wIou���)������94��(uy�0�q��W���>&>�4 �t���9ݩ�����{ٚ��5�/5-86'O�13B#�o�C�#�	u��t������@���	�ӗ�$�t<Ox��2�����a��W>��z����xDQ�"���(��$5I��*z��P���ť$�he�Q�(�Y��s �yۆ�o��c�5	�� �s���$�:�<�VA��d���ǠJ"��{$P��D�r����g�����3z]ذ��G��2ۉ3	Tt��8��y*a���U:<�f�������9�Z�o|d#�^^���<#��@���,G.��vQ��%^4��Н��uG�a��f����,:GUz�Z�"��}�죚- ���/���䛁
r��똾�Q|��W�fLlقbA����wg�.��飘���.�)J�/��PQ�-�!��/�4��?�
��|�k�kW��_Yd{B����.�Q�"z �����Q|�����hPdU��d��c�q{F�w��گj�w�>J�%�yT�jK��f����nf�����U)���ĸ�8�����Kj�/PUp� ���~3�w�	!���@+�K3��Gy����rq �D�pO�IYA��������T��$�����J��z�x����t9;~�:��2��S�d�9�(��^�h��_�n.�"��ՙp
QLf�6�<:�L�T��/��}��q��nѰ$�e�h�j�z�#(u�⤶E֚�3ݸ��J�����x]�Q[�>��Y�!��s@lg~�3�"|KЩ+ _WR-���l ���q����|��Q3s_d�T6�gʩS�����B�z:P��"���-M)L�m��h8�4��'m��#bǀz�:�|�4T����^:c0�7H;� sG��ʄ��;��z���F���m�JZeU�|�\1Vh��|q/���X�C��Pw`VO���ͥ�����-����v ���r_p��;൓����<��l&\�J�P.�)3X���"5���k[9�ҧ0�	��ӏW_��H�����O�I^A���˛m�EFH��6e�+j�d����@t诈��f�q�֓�����m��|�i�.8I�-�8�tk��A���e&��xk#�}m��^j�qQ��J�x�lF��Dޞ<�>�P�@D~D�Ň�e�tE6
�7p�͊���r`�(i�4#z�3�y&բ��ـ�׀\��w`8��虻�D߮�㔩����&\4���3�$w`�I�UcPW��Vf��d������nW�%J+�("Y�D�:�oVl�4ʲ��%�`�ܪp�k�S��Q�HLl��6�BK�����*���Ħz��)��M'p�,�3`�yڬe�r��#��#Y6Q;��حMݧ��q��_���0PB8�1���U��������ݪ�)pշ�Z͇WS�E�����a�&�� j��l��K=̿�v�ѣ�3�0�pc��*��k,MG"Hi�z������E�KS�r���eHʸ�'K�-�5��"��Dd�&n����R��8�L�;3 ��X�/�^Y�Ч{�k�#�[�-$U�o޽	��B��ou��vq)i��@��t����u��F�Z8 WY�qLF�P�U�w�J|g�٧�2`݋B&F����f��#�	)�V�@hvyջ�O��c(��!�\jP�fʷ`sd*M�x���v�׶UâE�H_,�j��_�P��R�O&��B�@f+$����V�z"�EB?@9$m�i�p��A耩�~����he�B��]:7��c=�ω\����_�g�$$$@����G:<���"W�m��@�Tq����	E�0�g`z!��WT�R�~+F���D���|�?Eqӏ�Dj1�vH	�t�"KT�Ut��\�âI�k��*薨�u-|iZ1؟?& �w3�;��D��G]�VU��H��>��q���}f�U�Fw��B�X�<ͣ�a:]��5`DCR�&{�١jwU��9R�d��V�ll�q�ŵrV��s\� 3ـF��Aq=7;�h�0�UYh��5�a �o�9��:�nA�!�4��^�k8��)���H��7�#�z��34=�J*���jS�M��6Vݶ�q���d�K��tv�l4y�(��;�Gxe�`��F~���g�rk�	VErc�7$J/J����:����B`ຍ��������-����=܀El ��B���'	8Eb����Y=C��~DxV|JB@ȼ��F=.�a�b�,x���~��\=pM�1-`V��|�0�UN���!�L-���k���r�����@TL�0V~I�~ qu�:�a0ߡ\�#P$U�0R�1�3e�JG���G���j� ?G�� :��k�r ��eQ��6������NO�}�Q?���,��4@��c�|�>��B6H��c�[��҇�(�Q�>��a�SEU\�J�\=?t4b"ڻ��,g��:��G�sǬ��gUrun�)��ih�8��k4K� !�	�� ����tޑ�81�RiVʯ�>�vs����2���I�B���+F�9<	��M1��Y��wr&A)��\�J���k��#P�����.�|�s�9�S��6 O xr���
Җ�O��%)}T]/�m|�#eШsH���[�8+}�9G�"��R���A�*m��P�<ej�N	ct o%�a��x ��cf���/ѝ瞇,�9U뮷?�`�
熖9�C�C�'X�M�#��1B�gk�$����0���I�f||�4�(�x�,7Ob�aw6�%*��q5�P�����5�B��"=�)����BXӺ]1�+�*�OO�i�֤�<����q�mV�2,�所ȝN�!��5��?駜�n��YJU����
�hݢ�%��L���VK��St�:��v��8�T���c��k��܉�6��z)F��Y��͎�����X{�A�nZ�2�&�t<1��w@L?�5�ձE"Xb���j��_� ��E�mF谈�1����ǲ�f�VV`H����a�D�P���U
����j.s�؅�W��# �����FR@Q�/���L
���WYtͮU����˹�>fgp�kӓ��~M��0�:+���8�M�  l������>n⨼Eo��y],���ġ�`�3��KG�ag�K�������s]��_�sxD/���.1|�pd�H�w�_xQw��������jE��>�H}�\"�U���9���g�Q@sO�Q_s���E�-O@e�K5�zia�Iu
I����>�w���zITUh�Wn�m���!��
P�I׆N�&��G��F>ܓ�ڱs��=m��+�@�S�}�jqs�Vjp7|r�aQ�����Q��]�k
_��!ͼMu˵�F�l��x	ؿ�X��+�ˮ]>	���&����M�U3T��[����[�;m��20$�fF��!P�j�y|넸�Xm>�G���D%b�M�U 9�ē���D�}Ԉ���X>[����?��)/^���������ZiЬ�'������MV��뷡"�yގ�G��h�p�i�ٮ�n΋Z`��� F�,,9׊�$���N����w�����61��[�8S0�d{�b���
 h���y��QHy�Y�̮�.�'�kxPt-���<�F�ή�W-_ɆXI�Y���TN��o�c@�%�<r�eҨ;�9�e*��F�v�%�Bv�W꧜��G\-��bС�Ε�J+�T�g+4�Ͱ�������)&r*�<�F>�������i��p�ķ"?evl�p3Ԉ߷�`e�9��BH�f�AΘ���� Ͷ����y�
�;� �c�SE��*9<����_~ �_f!�2�jͲ��Hl�SRX@;9a�Ԏ\��PdH��X&&�l;R��l,�!Â�A4 ���Gb#䳌p��iol���/7�;L�q=�c��@g��������8k�.̥����l9�)��d�i�'+�	�;�4���]����.�����y�눝ëըxx��*H���\,i�r�fD�RX��桺�H�L�xw�C܆k^��t���=cá�M�l��M
��DZ�y���2�M�H���3��W�t���g�h�DVmSDΒ:�M2��Em�<�J�|�N�[�Z�]�`�#�-���^��(���p���7���/��ݠ=/�|ЯU`l�d�; x�6}�j���,�g�a��Ή�m	��@���;Y��.mp[���,�j�M�	N��8�Xq�؄]	;���p������{y���aKP1�=(S�bS�!�0Bo8��S:�+!}>R8�@
7��s�r�C�C����B�k�ix��P�lM
�ֹuI��|��?��.218��tk����\�Y}�I➵��y��HW�` /NM��Js�5�R���(i`	uX��2�>�=��7���6I�W�kَ-c�&"����G�5;.�D^7V=:��+�~������Pg��l�w���yT��H�K��I��N�rvO�e���+���Qb������L �v}�2�"{5�y�T�J_�u�C3!���5� �]�����@ͯA�/y��wT��%��R#�I�K��I�H����_��L�B���Up���3)�;f���	h�?K^��c+���cu�_3�ྏ,\�]�B���Cv�����0bvN�'	'�7���yB�(,�%�����,3H���6Ȱ3�G������v�x*2�]�j���?V�&�&	k�"]̝�|�WFA�����C�|'�8�+]����}��=��f5'�o����9�G ��>e�Է$'u�;�q�q����t%9� *-׀�!�0�K8a���?�J��˒Spx� ���:�i�r;�.��K���~���.���[��\N��E&\+�3R��,L��$��ݠV��u�Ղ�fA>��z.�����eYּ~^���e'=�ǥ�e�ҏ�i,ꉜ�qǔ�����>�T^���).��I�9����!�WÚ�Z��!��zi��ТoB������;���7]�Lρ���
��S��fAE-��w�Y��ײh�S�\#<�7V��$( �`�d ��v���Lx�/�_^�u_�&&�U�E?A$��[]���$���O4��q��+Qͦ/��B�$���(��>��sn	����t�W���w�I�\�K�J�c��'�q.v��x�)>� a��}H���À�uZ���g�XJ����"��GzG)g|�?'��N�98���Ό�mB ]��2ٵ��*����֌�	�����=�Q}V	$R�����p�Tg �T��]�B	o�d�nȦI}����_4�����?�����t��3�i�a�0�W��q#��ȸ2�l�l=ÿ	�O	�뭮�a|eJB׮2�����%��O[�8��ff95tM�#bm]3#5��=%z�7����_j�y�~)�P�kt�E���-t�j�m����!���ϒ��\�>�]���Y.�,�	�p���G'��| Z#�UT;2�RɩH�Z�y>��E�����<;�ٞ�Ir�`������'|�T	��wv���"����z#K�\���%k'N���b�
p�������Cpyh��X���x:�n�m�{���{� }����a2�Ɨ���Y�F�r�R� Tڃ��)�gRE,���t�����̸5�AY߱GV�%V�aG��q��[�2g?���\�.��FL%q��l{a
���g��p1�` �+f�D�]�`)�{�mu�3�h��S�3� w��N�+�Ћw�$q,Q��R�NI�EBiEm��6C&��t�E���Q���S����$2&IU����ߎ�Ҁ�m�����
3�f�8����r8}E͊�/����iv�!./�vb�����ѥm;��7�LV�\��xs�1&H���&#��Vܦ��\�;qh�W	�Û֏�����U~�d�Jz�o�p�d�$�1�mc����+x;(���(I������'�C�m��x�	�ǻ���I�f�R�X��E���X�����ɊlfM_?-i��!cԧ}�����kBx�!��Io-|��42�q<f*Ov%/� ���vsAxL�$<��0j�0��
�i��e ��n#�;Ԇ���m�={�h��R�l�8J\yތXݭ����f�i�Sh��:Q��������t{e��k�#�l�� H{8�Egt�m@9��[C��>-3~U�N2{`�0i��%������	�}T�]��1�l�(1�L=�!�p5Y ���U�j��[P�9�pѦ�7�B���jz��}$�.y'`�{��qju07�Ǖnv��Apx�U	N�dn�/,����iM���i��?����;8�� �
�mWW�G����
��m(�@Um�mr��A���	`�ۀӤXI�+�"Y|J�����,�r�j`�!�=(���MX�	t����ӥ�7���ѻ�+�����Z�d��#�%R�S)��ɣ dU];4K7��ȆJ�.����K�H�?}�	�D!�V�xcw0%�����
 ����������}^#�G�d�A/�` ;�zg2c�8�`<*8��_#$/t>�mfo*J��>��L�	�O���3���6aԔ�����{���(Z���y��hK|�/��lY�Vj/e�$�ʚ��
$2���\8Q;����~��1�����^mj�UB�*Q?��č��#�g��!� y�W��d3봱��Ȃ��)E����p��I����P�t��^lpVDw��`�hf����ki�y���Xk��؉wq��Ž������a)�-� -��Qo��_��-8R�c����!�T��N��5�,{���9��Ju���@0Ҿ8_C?D!u����4�9v�˦�M�NƣwG=*/׀�[�����A�)����orbY�6W�NU!/<�
��ߍ�����P��b���	�=��$O�"�|%R�����dmWX�.��bh{H'z�*%뙸mU�L�4�H�݁�KzB>���W[�*#�cY4�h��ș�"�/ Qd.��q ��5�Q���);?��溾+9�:PsP;̩?��t�7��~t)��0\FrN�H]ƪ�F�^�Ω�9#�a�0HM���.2����Y�N41 N��|��/ڞ9��W|f�|���|��c���G��'�E0��u���M.���@�!�U�i�����*�r��C���4e��c�&]��נ�n�F����F�x	"��<�Cu�T1c��.8����Z�k��ώ��?���?���^����w�ǈ(�z�0j(M��ר�_���z�كG�E��uN��&�̀M\c�}C0` aI���O����|�R���t�L.�����Ўǵ�]� �vc{�Ţ���o�(��o���� a�PT!�����~|nU���B�j4�8ڜ󋁯�ǟ���M�K�P�7���ɨ�cfeG������L�DIRe���(�X�e�EcJ ���~�1c�W�HP�C�.8���/i����k�U����oǾޚ�Qޤ`��w9]��$����/Ϻv]��(��{��?�Nz|BУ������t7R��"�K��%���p��nzMc�m�>&���8�薗��;�/�Ì����KmQ���<2���� �(q��C,��@#D5�Ԁ��W&v�U��H�z�c������L��]YM�hxG�:#@;�S�y�*�"�(9��{�N-���c�`�~}כP�od8{��a?�v��-�3*�k���[4�,�mJ�~�c<�v���9�U���Cu8p`g�(�aI�v�h�Lk*37U�"�t&&�-8U��6�r���"�k����La�T��F߈�*YfUG.���b�B���fg�����u���um���BqB�FU2R��1.��zQ�8�v���2j�E��Gl�E����p�h�v�����c}E\%�xU��`��E~z�����8�'�6}Q.+i�x��)��'�%O�t�]�؝�ލ{��� �B ��7���q{�����-���O]������ݢ���ER7���~���]��j�B�b���!8Xʯ@y!m&�Z�!�����kp�x�0b1I�?G63(���s.��(��E��������*��<�
�����},tSG9��,"�aZ�,!�U9��S��@�2erIj��3��e��|����3�|��gtʐ�-�d�/#��#�T���BLQ�0��-�:ǟ�K-��+;z��j���`��G;JD��n`y0�B���5
=��^�K�� |�I�\X��r�b�Ɏ�.&[�����9SV��`?7���`
n�0�=)�)��ٙO���Z%��ɷy/�.Q����>-+�ސ|����e�V��/��o�0��U���뻅�::�>��o!2�IF�l���PC=�y�I����8�yyK9����x�i�l�j��P� ����+�8��Q��J=��(U�㛚��r��xџ���C�w�,7jq;��5`��J������s�}ׇN8�W�O��h��,�˭E��}T�A��L9?��~$���rW�w���=��ZR�Y�o�dl`�z�7�M'�� �8x�k�D�=EA�$2�w)g�g�J8(��'l챲\���7�wR��Z��Xz�� E�۽�hk_E$i���U4�7�f��#����AT����b�oڜ���3���#2:�Ĭs��7+�����¢uB�
!���q�]*Yxы��f�7TL0	��D	������ќ%����y��q��Ē�].�^�A��XA�����<���D 	Zs�+��f�_������AS�$��>!�7iq����H��J�Z�`�˧�F�ô�SO�R��'$��k����Sa�H��>ʝ>I�?��
;���#���.��b'�PiZ��A}������*���9�R��uK8�'w�9A(�$�9mm̧����8
�C]眅^������Fۯ��+KJ��\�_��l��ǔM��P����?��������'�B���{�hT�h�uO����7`Nlk�(�R^�{�v���tU�]�Z׻���Ï�sĭ��a��1��|S� n�Ð��/����IǨ�\��i�-La�˩�i��PYHz!=�2&n26�W�F�)�fؿ�B(q�fh�� V�5I/; ��(J�'��Ո�ͨ�a��V�gW�����_�$��>L}��"Y���6���t���F���4LA����W��p8"�����Ъ���z��~Ǭ!Q|#Y�b���s���eo_�0>�#@��ަR���Wje����hש��u��)�-�����⳰5��"kɦC��&�T+^�s W4�0�?d�~�ݑSb��
7
���N�!�UtMW�m�W����O~��C�VMnԘ g�"5��Q��eCW��f*4sk��ʄ^naF`�y��ߑPR㵫���#�L6s���ɚ!3|�k]g��Er�����m+�0Ahq.ks��}${ݥ�V~u�g��6��&����3�W���y�^�.���[ �V�[�b�@��LB2����u�Eyp!��-�؆�¬���:���O�X����+�6Sk!�����[��w���hPD��bMll=�mv��������H�	@Ћ�b�T����Z�y�$�< �^�V��k�f�ٺ�-J��MP��7���4i`%��5��V=N����@VؤR�{�-��Q��=6�P�bV4w��Zތ��F�7׫:�P����!}�.��C
O���eN�+��K���gH�,ڽp�[Q⺚J������tm�U�=<�U�&@LRFv�!�do?k��=��ט��tE�1�vd-���yz�w9�(BG&�n���*]8�Nմ_+�p�Ǡj���`�~���Syo��Z��dE�A�dP(�brk1�Ǌ/(c��[a����I܈�+�uf�Is��D/�3�C�"h���P�(�y���r��31�{�f`ރ���8vX��1UGJ����T���#�q��{䉡��u�M�������������ߏ�;toU��� 탡ɇ�v��Ñu.��os$цߝ�����f[;h\�g+>���>��]����K�e��A�\�d�<����%�)�z�r���I�8�μ�a��"���C��_�۰�0\c�
דl��W�2!]m�K��د�'_����\��x �懄���5�rx�h_��bT�\��U5*տ�1�q-�-dê+��Ϛ���6��ڣ�]K�P�>�A�ǐ�4�[��T���o�����v���7b`�i��`R�Z�[�`~�6Z�������/���F��u��@C��G��t�Q��z�Kj�Б��Z�}6Y���C�'e�_㟿���V�(RR"K茹��������4UW��ȿ�h3?��c�F=�ʟ	�:��ƽ�(D� ��?��r%�bul()3W$k(v�TS�s�.�F.j��gУ	����j	v�{s}J���j�����/��r���� g���׭P��
����P��^i��m�ˈ!2b�7xQȌ얭�U�t��/�����B��qV7 �vG� ���v��|[<���{�~7Q�U��=���nXq���1?��β���t�T\��7.ײ��e�o�m���D���9mo�<13s��vZH��c+�x���I��e���U��SAI1�����֧ae�SZ�Y4�G��?��on�A�N��=�y '�I��|p{d�֓!����晧��^
�,`��a�V�
�ax�RKh.]G���O1��?��R�M �'j��Ͻ��F�!��,�(��l���>if��C�Lf�5���i�baqC��r�6P�%ɗBu�!�韤����A����N˒���od�A;M�fԳTC{DSn"����U�+���y�״�c��~�w���gT���;
q���o:}�i��yK��Ⱥ��+]G�ޕi�&L�\��[���Sv'�����g��,�����*�EZ�GM;P>l�ᡉ�1�c��ؗ�������7b��G�<5]q���&���;1.q��)z��v-w�w�lR�/�ر�����Rhѡ�5~K�#o��Sٳ(��fԷ��34;���ٲ� :�}o�AtB�R�<���#����2�3t��}�P���_����Q�$����Y#��Z#(R�����w��M�n�����˩ٜZ��4��R9���dI��ɺ���:__tA�4D������$�E�3���+n�9��O5�q|�8��O�ʨb�C�E8��&��\�	�Տ� cJ;����îO�9�tQ����Q;.���C=3LW��L(v�eAfJ/�����Td�:��bO˳o��l�fw�޴_,�S���rJg�A��_sV�|�%�Oh
��a�)Ժ.joƔIAԨ��$}�*��8���*�������iU��K$j��n!��C�5��ق�E�X°6�����#�Bfn�SoC	���dq�:Z'A��0��h:+V[?&���ܦ�|Vt�17�`�_����3Ƃ"��4���+���¬��Օ��s�ʦSgZ�[KH�+8^����