��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��!N;�?'ǝ�{9�1�\��,�L�B�8��V�R?��[6F+�+�4"p���n�d�#�$؍p�����.�{¯q��ěW�F^��A�S*��|��Ea)��sz�$��O�+�d(�W�n{�|��C�:� O��U荈PjZ�h�'#��}�Z7��-?D����͈#�26���1�o%3}V�9M5@�����s���F��	+�5�������S�/	��;;�~��g��JRyyҩ�M�'������Q����4�1_A�<�����E�s������?�I8��6U�3[����[we'C	�De��m�!L�����;ܜ0��V�~Ջ�r|��˛a�1X�=��
�M<3��(&�<�<���U�p�b��)��+1��+�����=�	�"Eβ�,�������pR�Ry�+f߮2j�۞o

�,>��������wX��2�:D�J ��� ��<���h�S[��h��-(��(�s0�9��5�[t��s�Lm�����S����f�fQ
���3��?�$7I��Vٚq*�T���8�!yxɕ"��f���&���4Y�v����^�re��F��������]���g��D���?��EH���2SM�>ZT�Ӷ����k��ֻ,��9p��3��XoS���,������vtD�S�Z0#���:0��8��Bk��{����7��e�ecQ�6~�|��/��8������y�dgO��4Y���S�`�_�� �8|C����6 �N�.���]�S=W�h��5_ @�WC8��#����d���.'4����'5���@FjL�D6)$2Ctc�,?������	5��f �))�\<~	�*o���>_v�N���ZU��9�`�ly��.l(]2ȴG�
vꑩ�/���E}n����'�ZG��b�U� ���-fɦH����eÁ����&�"w
0R<�{����-.H�b���r��.�6=�{���5�3�?,ۇ��;ր������$�6%j�r�D���|�ֿ�w�3蔀�b�pM�-1�3�vȨ~/��X=�H̹j��.�V��������}_�����4���ѿY6�_0
H����Q�9�֯uFE6>���P��9Ԭo�zD+���s��1��E50=�+�����sG�(��SB���?�a�o�C���q��W��
8.����G���͆lb�٩��2������'/~���~E_�I���p�'k:�M�������ƃ�S�z�S
��ƺ#v��k��؀t�N/?\|�qe�nuT�l�m��B%��.��F���S(8F_����W��m,����&��sW|,fT�1�Ig��m!������~qb�"�|��G�l	��R�6B:�� ��g�r�λ�0���,�����0��/4Y�.��_�WM0���\��mo�\��K�葚l�k8V�u ƛ�i<���v^ӏ����߶��ҥ���s�K��W2^=�T9�]�|�z�����S��U�=��:�5ߴ�8�R�b�a��Y�ܦ�]�]'�sL��-�S<s��}��a41���L��fvWVڝ�8+�;����f����WW�B���>@�^f�O���%'��թe�^c{�tҁ��@n�[�.}�3��%�4.e���@���	Pg	�q�l-�'s�m�J��2���/V�$�u%ђ}�J���ܬ���� 8B5)���B�v7b�`_y�T���=�,�i�РA�=� ��é����'e�{j�B]2�w�D�F�H�Zj��;��W9D�Pm��*�᠗ٵKH��G�O����4*)�7��ڄ=�r��=:=�_^����G�ц�	 �W��Y>g���x�t��h���h�Z�����a�)�ƴ�����96�h��56�(��
�[���Sк�e�}�b�yo]"|ՒG�ͤ��Py|Q�������+	�F����PU���������1p��A�F����]x��gaA5EO�F:�.ꛂ�:I�%�/LU聁g ����t\J����X0;U/���dУ���w��]m�bH|0M�K���RQVL.��_%��W����� �5u����	�%�xlH�5��ĭ�,[�}I���%pK���l�m�֫	���e��x��H^>�������fz����%�� U%N%�
Mͱ�2�������x��k�:�ź������_��ՍpM�M/�m�4U������rlu�Ld[�9�Tx���7��%�9ķ�<P�"�C���ݪ����H�Qz�K�㠀�x�9R5�D��4<FN�ܝ�r0���u�H+`4iSRyyVsVR�%ׁ�ۏ�$�Cša�V	t��=�!8��6r��[�� �Y^ƺs^�'���ŖֲP�2�H��4���-7�u��ṆC�!�� JWϳ!��=�������`|��r���ɜ��Q�Z5l�bN����\S���r0�;�c������/��%�s!�Gۙ�CC�t�S � �[Q�>���BL�A�w�4�&�!���rî����ߑ�)��ZB}m�� V�"/# ��3���T��L�)r`�0d �?.��ƌ⫭�4F�N������FO�0���3g��هd���ȱby�C��=r�/f� Z>����0���7��Ѭ;�0g�/&U�E5�����&��v9�Ʃ�(��~����O��I-^	�8��>�����g�����d&F&HC��D��*^mr� ΐ��21�f��K��c0�r�d$�v}iV��$��έp���{�/���C��)��N��JAvͤ�P�(����n'7�
������!J��e����*סl�#@�XZ���۾�#H���C&c~�9*#����P>G����
?��&��nC�CѢ����Z�䂔7�@����P:�f٣g�i�Y��L�����