��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�"]P����'�*����,*k{�D4Y�JW��<Tdi+N14+}���:�_w"�΅SO8+|j� �"��\�od�x}�k@CX`������;��T��d�ȥ	�8�) �ǵ#W���gㅪ+Z�T�/q��C�,ȷ�h?���5�8��濤�iD�޶}��9iX���A�^�^I'���7[=����.ץdM+�o@�.Vq�CPX�6���m�ʩ�I+[�Io�0_nCoe>�L�z݂���'xy�R.F�}�|�҉$~��]�6��%�.@�ɋ�����������gq�YiO7Ʈ&����lM���C#;˔z��!��?N�n}G�wlД�D,E)qT� YJXD٫/�V���/�b�{Du�k|�0$�L�Oq��F�I%��q��?шg����1��JԾC�7��Xr<D\�o㙥�x^i�Y"��<pF?��c��$�80��p9_XU$ݰ�,�j�	.��s!$B�N��{�m�n�g�2q�5��,W��gLO�����t�)���t��%�\��ݢ��D��� r{2��f���Y�ֻ�x8�'�{g誛�&yQ��|���'����8F�ݜ�
E��J����B��<G��O%48��|����k�)�F�T���Tl2D��;6a��tP���zï�9�Z��N};Dx�8�v"R�"��N힙�K����B�$L���z�@��1[R9�@�#gȡ��Y=�i*I�ȉ�I���Ď�ϫ��h���֌�=���Dn(v�&��PTt����X�����Q4���fɲ�4^n�'�©m3VI��6h��:>�+֢����W(!��� ��U�%�{[j��Fv���K��F�_�1%��;;������W��<b,���.s.Z�86�-�~�b�>�f�lGx�>���� P���&��6�X3UF����X��̑�{���"G��#��t=��;o8R�*���Ԁe3��s)k�Qk�5M�0��
�C�Q�b`�p�V<`���X�P��sC�#��_�w�.���s��
�N��(��О��BN�]U������Y�-F_,�y��H]��ݞ&3d��f�ID`<�eS��_W�,�i�Fv���L=��2��u�k���0�Ͼ�`�}M�Ѵ��J�d�o��d����X����!6�"d��_'̩R���t#F���NXd\�V�#\1��&��D(pzɮ�����(S�J�h$��uvY&�O�0�1�d֏��$�>�8!����z��,��vƺA3�t1<���K��M�������I���J��n��XoӞ�6�X^�:��\;%g�p��1������6�������+:�y�J�A?B�r;�%��|��Χe�k�>�H@3���M݁e׾wT�g�/!�7����A��1���Z�N!$$s
N�c	�F'�� T��޿�dX~��}$�z)W͌��am?�L��� #Lm9�ǻ����<6��ك_�m�d����t+:r�DM��9s<��r�ʜ)��x��(Xh}��r�+E�"Hp����X u�e���:th��}w�|��"Íb$i��}CE>#+0��,�Yc��a����pa��=�\UH���b;9i�J���mrM��t�E��W�O�Q��Rw�Y�jμ�B�R�)f�j��W>hɻ�`��_7g8_l� ɍ�� ��rт����p��@/7?�3'YҬ�ȹ�;�O�?�RZmC�Tv~d��BSkئ]�:�8��cg�	 ��=�ϝS�q�dV���ٽ�i�{�bX+�js�^	)�#���QI��(�t2� �mk;�<�at�.�,�-�"c��QW������ߡ����D,e��\�}�n�BD��.� t��K�t�=ll������
�4����Ξ�H0$ʳ�T.�O$�g%F�������R��'s"o'���[b�&��O��)��%k���,>�8	�Éz�d���n�B��%̲���r��(�M���^���ÀP��Ƭ�:�f��*we����r�����X˧��j���<TA��T�P@��,Ԉ'qR��]�Q�ye�r�_��5mur��.L�p�H`B4�lݣ)X���u.���<�"���&"����렰�m��m?˥�AoK�*\��cR��}�^iː3+}�������<h�zb��@8��n�q�?!#B��0hGl�dR�Q,m�Uz��Rq�E~��f,��턷vd�!Z77(�$�)b�پ�ůU�H����o����˘T��BG?^��`���glE��(k�hޓ����M ���)�V���j��J��h6%#�]�@Ю�Q����Ɏh	3w��nw�a�`2&��)���f*��[����V
�H�	�"Rڟ�&�FL����N>x�eM�r'��g3�QR�eN���=7�;I)`z������4ܷ�o����<h�ʥ���LY}��W(p1|�����Т��I'1�$N��`�"�q$�������İI�.�1�����>�s	��p�7��ܨ��J*����S�Ʌ�Y�4'��w;]�&�翲��s2\-�+LP&�D~s߲��4h�
�V�����e�*"Ud~#�A�A�y*�V*���s7s�z�P�Uk����Z��� ��v�\��ekK_�U�I,��_��Cj�TV���5�UC�Ȧ|�y7!���ֳ��ߧ�7���
�m�!�-
B�w Qv#��N"j{���J����*$�����͆��HO�)��R(#�P����V8�Us��al�=ѳ�am�Ӣ�I_.4HL�v�d���z�u1$���������E���n�@y���+�^�0뤵�l�X�֐�B�L�!�r���ωð���5��q��������FYO��5J�3�A�6�kJt�X����$�K�� �Hɏ��8JT�z��kq�瞿����~C��z��A��Y��-��j@�8�2��>�Tt?j�B�Kȕ2j����j��&�.�X������"e�^�����l^䩎=�c�4���"�k*�|�'DΜ�ҧ\�>+���4�|�Ƒ����9���n��	n��#�)���vD�A�{�i��S;�B$�`2��z�NǏu��>�cu�D�n�&f\���E�r Έ��䁨������΄���se���	� ��У��t_�6Ӓ����lϜcA�7&iܰ>����(�R���Wð��.��n���c��ߌ�?A������3���
9S��N0�&����\M��5��B��B����mF-���\�����/�D0%�ֲ�q�>���S$+pP�	���u�a��L��2"eA+