��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9h��=�4��QDG��D���������6���Zʣ�餵���j^<�y�F���	B��k�@r��Ah�B���y����SZ_|s�du���@�g��9>0V��L�
��o(J(V�r كk���\�K/�J^��^g�5G��U��qO�~�h���M�h%8��r�.%J%��q��x��_�:�8������8J��=��������M0	�����D��H��[Di{�Y��	9,�C�|J�T9�Vb��e�r�3�&s�S*`s�(~` ���z�7T��t�R4����n�#��J}UR�Lj���f��H��J>��q�C(�D��2פgi���@8'e��a��<��*��Db_~.�������^ô*!:�OGd�;��sۯ�ݯ�ޣi�؃	[�'�Q ��/q��]4$��-V��z%ax����[[vJ���s��N�3렸<h��K�L���7�@G�Ǯ�i�B"bn
�Ʈ4q�0$hb�+��Z��	-��l�����!��!��%øI�2���Ι^���P �fO����!��_� $���Xs� "U�4/8�DMǬ%nQ�S![��R�����{LT"�қy�x*Z���r*Ғ�j$gi:L��	��G/[��l"l5[5��� ��ĆJ�k�9�����^Wt4|��~�o�hz�bH�W�H�R<��S,�SW�UĬC��lH8qϥ],�[h���f)�Ðw�Z4���U;����]��ڷ�S0��u���NF��:s�doC�Xͮ�^`�upW�'k��ޙ'#C�Y�)M�|�9Ix�,��6�NN+F+do�����
�����vڽ,?����`�H�c,\��t	����}�n�A�5Y��z�Z��\��R�{��e�iC��7���ɐB�GE�:q?���{t������3��xi*?�al�	�{$74�Vh�労�@?����q��%��tj��d�L��DK��p����j��7�+�a�aG�����9�%��Ƿ�ǋ6S�t:�K� ��߳��d�6R`+B���+R*�����?�����(p�k���,��l�Tl۠�C�nOB1����J,��VoK�!�����Ci�: �j8T���_&֓�~a i���)e���
���2��.����RQ��t��zT�Z1.d%0��r���4�!�^�bt���?��D��ҋ6A��T!��y���T��T��#E;��XKۓ"S|:jvb��g�$�}((��96���^ʁ�~��l��2"�b}`�#�}��V�GμH6	x��^�D»�*j$��G�:�2���<Z���9��ָ+/;g�-R�,�����@<�
P�cg��(yu����L���_�n T�����?
�,���1��$�s$��Y	�����P��l���\��R�-3�Ѽ���M�6�6y��-�����xͲ��������������Q)XR7��D�ўzS�K-��E���C�T�����ҏ���;)� ���I����C���L�_�~�\{&��-ߡ��s-t'��ǈ�cVIE�A�|�[�tv�GBhΌzǧq�KYq:��)����9T�_=�2�.7p��J����&�?H�t>������79�˧��LG��XyP;�	��D+��㛓��i��	
�N8/��u5;/�?�����L�
�p�5�#q^p"BO|;�;����Ĳ4|�4ɒ���f}��@)\��=A�F+,_mǏ-��N��;�4�V|j�h\/�T���������������{�J�HGG�il!�̪�ל�I��m�C����6[��^Yd�y��G��Չ�L�������[�"B�4	�O��[,�m2�j$�;�H��������������Y㵮V���l�yD�S@mM �l?�_��z���s��ɳ�C#�)�=��Eȥ��,��u"�y?\���u��q�Ǎoe[��s���W����"��:}�;/��5�i���2����(��Ө�nj �V����l-��]���Ű��!�D���4��B=�"���{�t<�U{�ۙ��I�7uGs��.X�}�CWD3�v��u��pu����z�T?iO��4Ն�ne~�O�?�[B��1���&`�a��N#�D=�S�RQh����j�?
�7�w֘���x�2�V�:�Ϻ��������E%b���
a�9�C�v��В1t��"���4�1��H%·��(=Q�w^�p�H��*�:s�&�4�|�*F�0/N��~��~,���s�!�3�G��fgΈ����
�k��(ڿ0
���k�} �����ܝM��I,��9V��k�-%�a��s��*�"�1��΋��N��pC��T �jأJ�b��^uh������I�@{���`��"��k��F�� ;1��=C˗��3U��?6�T���4%-,���ɯ:�^��(�Q�����⠚�:b���qxS.Q�����邭)��X���˨�=�|��:�V�9��A��2�d���T<����+���Ɋz��l��L9^��Ԟ7��i%?6,�#B�9��%]�������	��bPХc�e&�g/0�s��d���襓
I��4C�|+Sv�KD�N�E�[����e�(~�W�Lds�0���a�SC�K$1��4��减�7s\�������1\!���#��U��@�� yq�X,���6��"�%��}���*�xM<u6e��'V[��"��l,��m����8���$g_��ֲ�y�	�b��O'N��:�5�ϰEN�;}���z�g��C���X~2q!F��)V�}l��q��GA`wؽ�J��`֔H�m���:h�+��0ep:ɓU��Zl�AI^�:\�w�}�̯����{vk*z�aA�%@&�c_�ySO�M���fN�`Xd�Z���:�v��}E�X�Rd��q�"O���,kH/�:B�gE��B�K��D����#���;��Z��+N�m��U��Si��	B�o�ǅ�.H/SC��͒��G����2@��)����/�F�?�O�❻��&�L!�>*�Qi����l#R��0��A�6�a�-W�Y)ܐ�k�=�d?��o��U���lԒķ�I�77��mɲ�������*s�)��t�?��ip���,��I��*�v�|^����:F��,H���;�w]0
�1��W���B���l&����!b�wo��b��_\�-�C.o���K����a5Z�7�ک��ډWt�b�e0K��3��%2gA#��]$�f�(�` t����e*���6��Ou��#��O�����qW�ݏ�8E�uٱx@�}R4�{��(B*��o�j�Td��ߔ����1$����<����}��5�&���u 
�7������{�C��
�n����}��[H4Ef1^$���aTM��9l��;�>'�o�#��)KJ�_R����i��|v)7� �p��[��|进��� ��&�����N=�����z&֪KS�rއؖ\3�`�"���a6�Wy�vͩo�E4R�JL���Lҷ��)�_̟��4�`5��[��4�	��1]��<������:�����&WN�<���(�N�:t�ZH�������Ƚ�+P�������N�4���\Q���o�ʔf�h�V&=3���Z!l��xU_�P�`'�;X�7�[�
�?��i���3Z��mpDR+#�e�(���0rh���	���/+�8")W�":6���3`���X��	�����eE�g�Ҫw"64:���{�1j�0���qk�.@��( ��b�=�W{m�f���펭1"�~� ���,�V��]c9����(�|{Ǽ��v���cc�_�L��4�i�ě	��H�ֹih�-���[�F��؛/��.̒���玤� �V��;A�Z��=x�=;��%��M����J�P��.��bZI�#8NQ�� e!�5�U݊^*t�M3�uKkc���w,C�bv�n��X��r-ҳ����G�g�;�h����i$��&It�`����)DI]5�fy:U��A�E�K���_+qp���,g'v�=��#KV��r�UK�+��S�-�LF:��mk� G8s�^we"���L�4Oڇ�U���7�~���S���T|�Q �9��bi���<YILeO�	���63A��|��fL�;r�K�fI?��׏7��Fˆ-��Κ|��[��8	�qZ=yf�e��:EuR���m^N�N�!��,�I��6X|	q����Q�࠮ܶ�D"��p|���%T��Y�&�0�g!����<+�z;p��ܩl�(�K"$��W�P��x��I���0u�dbb��l�s>i�no�z�)!�hC�:�E���9��a��y�������x�������sJx�ΐxr+a7~��!k=��\H�)��T43ø�{��C�%��y��,N���u���
�_��*���a�Qҁ%����E�U]],���w	��#��B�d��o�Tg�O��m>���+��)ɱȗ����j�*Y�����_j�Gc��z�	�uÒ��$�#OJ�N�Û\��6�v��C1�U��,��
��VB�yk�AðH/��؂p,Y�=�a��ȓG��E��CV9m�]�D7��WA%�� ��Sa��r�f�-�Z<���ĂWK{�wE�a)�����1�^5�����x�%�ka^�OP.
so7e�j !�[wi�᳽c��\�[+��yd�`�㷂�������|(K�+��e���,C �6�Y�Y\�y1XJU7Wp�כ�舞Kڈ�/�x��=e?�SP�7���x�2�Ζ�y����4!V�)'��q_@T�^x����`{<����&z�fw���4&A)��dF������G��6��v�W�F2�U���/�~�p4����Yu��`o1�qF]���z���m]P��[f|