��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&6��i��N�� ���r��
~G�+	�&?��D��� �Cb�v�	mh�b�D+�o����S���^� ��O\a�V���� 7F�3�Ћ`�Ρ -&Ϗ�M�\_���`�H��y(9��Q~��M��g��$��~��`�p`Rm���&�[d��&���m
Y��7BvT�M7���!�l�!�����d�s[5z��
��?{��]T��j�i'lE�4�u2�4�q�|�\��S#�C5��!3{	h�c��U>1�Җ)5G(��a��6;%
Q7�-7����ͩ՛���zA��˧�� 8�ӿ�pJ�JJ�A!�F�F�Co�x8���f��y��W��*��3��#f�l�͑���P�#/v���[��~ׂh�S,���u�O�Al[���O3��7p�FAݍI��C��7ґ+���q�[Z�b��"G����@��P9����Z���֜�}0�d\5�pN���h��{k�W���j�}`:���B¬�)�U�״#��*O0y���y<3��Xџ�л5�G���j��F�it$�:��u��I,�� _H7�d1��@2��=�C����Wʄ�=�T�+��U
��ħ\��о.u��I���nI����������Mw��lS�֩B^ g����&��Oy+̷)B�[اaΔgť����e7f���zN[���g�hD�&�7�ٹ�>c6�+���_A�sO�R>�z3��e�H���A$j�����ORIA,C�SטJ�U����Gݸ~�3;9�Ԁ`���J�aec�L���g�O�8�����a(K �z�H̱��^������[����#T!���Dr�y�D�����<ZZo�eV��J�a�>�f�4T�TcJ^ �ٕ=w��*�Ñ{x�Z�����F�^�oV+�9j���u���π�h]` 0��"/|瓆D� ��s	������Nhp�3&{�k�O�$D(b�Nʓ�6�����C>����kN�T��EZ�N8>b*�~��;�����x�$�}&==%̾7��j����1����~�]�*��[lرu���!<���C�AJ�"_2���O7}���V*,=(��k�]��[y�J������c��4Pr�X-m��Q$��"��~tf�l�� �Ľ�3`�;\���.��c,�Y��ajW�������p�/���K��2=r��ã}�@9��W��&#qO����Y���F���
D�?�eM��a�r��':��N�XǑ��3\pVm.
�������g_�^D�fT�"y�Zml~���K�������ʭӔ���=�`&���$6��&����e0X��\�W��������ɁR2Q�Y�=�M�Y������8�`XK�M�bhxͮ�}1�UoC�e�Rp�
�I~��yYۦ!SX��/lT˨z��dX��wbB�=��]M����oA��z���t�_���}�Q���ރK@��iX����[�XW�sQ�J�o���Q��(^�3�����mI?[B���عo�R-CZl׏��m�C+�x2l\���dpj��`3���*��r�2	L����J��j&�����I������^W%��@�=̀�y��r�%q�񣅆~e���c�d� �p�U��*���dq�[,s���Goͱʃ�a:������վ < �i>DJ����\}��"Qj��*5�iz���I���a��.YF��NZ�xN[{�z+?wz(P�4ѫo�Q�(a���ءm�rq�R����[^�05t�/�
I��'�+������זL_y�o�nYq�����Q���+}�2������'�3�D�����ii�-s�¨,��L�
w]���TW�_���X�#Ƃ�Pm˽��9gvȺ60x2�Yj�^~w%��)�po��π�RYw��P�Hѐ�I��'4�h���;:[-��$���3N%�bQ����(�N7�Yj�X^hIB�yW�Z-�3Z�WV�yD�v�.3C'-;�h�a[��;�)�ʛW]��"S%�@w	H|r�8wM��gC�h&.�h+�g�Ҹ�P�U�(JY?�c�e��Xd�da1��]q彀�I[f���Қ+`���?1�~�hv��wγ�]W��?8��w�Z���4g������ [�(\���XH��(�r"W� b��5��f����5u�5&;��:Ѳ�5�܉��ar�&�,��_�$�E��e����<WH e��k@-b��
���H��|I����VF�_%+�|��ҹ��035��ħ0|w�g}&�*J`�VlÌ��0��$�oo%�V��qxɣ IWX9�̗;�W�z>�q��3먐�O��V�r��MXH7Qz4GN��Bw)���� e4����z�e(O&��m�K�9��9M��|5�e�O[w�	�Tt�3�7�[��1��b��ϟu4���Hyq�~��rPⴀ�����8��.Z��mp�ZT�_��y�M�H��;\�|���CK��DPE�K�l��I��#�Ċ��qJY�VMG~�3���eLK���foω�����} ��C'����h�
�YP ��a������LdPT�"K���{�g������p��d��.�p%�;��!sI������o�t�|�Tbi��/����j��>gn���j�w���P7�ZH&h��9�1��Т�dm�6�������F���#���LzU�����h� ��5Z<~|QP�(F	"{֊��rG����O���Y*�"P�Rl��W:������v�+|�R�s�;���D�iЇ�FO�!�a.�'�������ᐒt��8r$�:2�14��jP'4Lc������
�&<P���:hC��d����A\�w;�a.�ڼ��1
,��������2���R��w`��6�k �-�`4�o��uKC:�9���>b,����
�f����k��Isշ���WP >�����|3r�1b	DL�<�F5���2���[f$���Y�$s��I��\)��bI�#5��k��6��x)�������v{Z��N	9ݜ;x�4,y�6o�+��� ��B�G�ҴS��Lj����=��<ޒ��"v;Y6ܻ�֕��.)�>���yJp��-~	ߥӾ���[v�1�Tq��d�2=ۋ��>����;��q����0mh��8�0/��2�.r��nk%J��V¥�?��2C�D=�#y���	,��5���LU���S-="*l8�Vt��TؤJ܈/���)���'*�F��-D7��uC-t2�~�8� �*#Lp��M:������K[k�3��O�M�j�Z�x���W�(�����h�O��P$?����h~ե˯�:��Sz���+��5O?�' 3)�܍���zb�$;>�U�|��4,�{4�#��2��Rg1��]�j���޷��D��Rt�m��@�=O[�}��)�-e�O^�5��+\�OqT6�:�<�Rm�1(8����d����g�>H�#o��~�F����?�7�ֹ�A���̙;��YƮ��o�f?�˪Įڐ�%�Z%3e��5��9���y|}"���;��"Ba���?����3f�o'��e�ñ�\ݠܐ�(�����q��b���
è�6�̄a�������3��������V��=�OVk��ߠmj	�6B�Ū�/�DOqrmo_���H�`�z��n����	ɳ�-Bn�� ��X���ދ�l���	��(o����a �\ 2���x���=k�b�!E��/�/����ϻZ�I!�z:<��(~���
���)*��g�Kq���">��EJ��n@�j
�����#���?�+���%�d��l�τ�	>��z��D�-_0����Py���8:�N�Q�ZnE"�����.HL���׾z��RG�JNI�X9�E tC-�cg����0ߗ����jJ�YYP�pP*k�To?��;����� E˼���z7ϟ
������vQ)��]��6c��,�-^S��w�!?0�A�ގ����B]�,�1zg$�`88j-B����<�ћ]U�
�"ڷK:��Az��xXWb�+�[���&��J��jP�!ރ(�ߠ��<`����������8���VK1l�:Ӕ����JJ��Ҁ2�s/Hj9�{�>C�X�d�� X�i��L'���*k��4�AaV>���Pye�{?(D�ƅ,��8�z��9Xª�|��gǜ�\���2ȃw4Z���B�f�E��q�,PمԺ=���'�²�$��Π�1uk\Ve!Gi��>����I-k˿b�e��BY/0K�7��ۏ���S����J��z��
�m���� ػӿ�J�^��[]�ktM�h{�kA'����8*-Y.��f*��%����T���ƋA�Dw�r�w����+h~-�����ܽ�*��@\#�?��Y������[�5��
�h1A�<#��-�`�1i���O�b�ur��_� G���������α
|�~R$�S1�����z5����QdR�::�W[�[�:5۟gB?o������C���lx��*9�ߜRx�@W"t��*�̷�od��N^�z�0 ��<���?Dz'�A���8�S1�l��]i��7�XsR�Aa�g