��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7Ɋx�!�g���I'k�c�J�]x��|7M����Lb3q��������sq���>B=O[���c�Y�a"s[T��8�B��s��7�?y]q.[�s���ޯ��	�ooe�bx����%�&�u��lM�����������;L9��o6�.�gb폔�'�Պ���L���}�@�v�y���:�Pbׁ+P#	u��kʯ�g�o%أZ���ߢ5��x���{�\=�_r�²*�Y�1�.?�)kF����P�.�2R.yX�s<J���Ƈ�9BIU9QT5^��j4ě'�S�)^�8X��8���AD�s?�!��S܆��O�6
/癧
g�T��Ƶa�q�����/1n$�l��v��.�G����	s$���^4�
&fW(��9���FSĻek�+�)�7�C�)ꩅ-�6��o�1�6�F�^��{u�T�1����0��y@���ۣ0�IՒ����+�8�¼�r��n��ڹ����_Rܢ�=I����(k����n)��H]6A+Έ����*<իA�iq��#�����I��5���OjyL :�Q���'�F��3Ѭ�������Bݩ��Axz���
������V9a21H�[v��>�Dy�x��$d�����`�&ǐ�'�@���mDw����G���I!>KcO!&C�D� ����{�z���Zͺ���GG
����$"��dGm��V��x�S0��n�!%Aժ���4?4n����|2.JIWl���Q�؃mZ����T>�������A�Ϋ)ë�e�ӕ��)���U��<�OԞE���ߒVͮ(�&�b%�X��D|Ǆ��6jb��yh�_q�SԆ��ˆ�uX઎�Ǽ������k*pA���iߺ�ma��0�};op��|��{#M�!l�`��� �����_2q���%Efࣴ�N�Lq3[3w~�HR�ꒌ���M�?�D.����D���2:�$,�;����h�a�k���sP<o�*9'��M5����#���x۬���DW^�n��
pW"�#[���Ω]��߲4$6�t �
aj���(����14�k`zH�k�G����F3���7p��.W>N�*4�YyQ��Q�� �Mc��A*�\n���z���}8j@����������E�4"��T�*�x�9P�,0��M`���?4ě'�U�6l�yo�/���u��5�Af.)	wW'E7�}��P�3/�0��7/nTDq�*M�~��G��jxT|�^TZX�~�ί#�-~�0�����WjX[
��vK�kL&zfj��3L��� e�Ё�|�r���&⮑_*�$s&�Ml�f�C�����]�7x�xa���{�	'��l�+d臻�W
Hi���3�1���d��Hu���iL�&S6M0`���_*@��s�;�p��5��LkR棫�`i�����2���P��;
�,�qĦ.�I�O耇�i�uP_��?^S����5cZ�1Jt	�ªz��7����+�0=�"��������u��G9�
6�&�u����B�{˵yy�=:6N��EZ�^�b!E1��i�s������Z�'���씥��e���eLMD��g�CN@;�4`7e�/�����C�8�G 6~$�M�PF��(���R8�f�i(B�� ��_��x�(0��0~�)v�K(���r��k���ї�7aɤW_Wq�ŀ}�(�ȋ�TS���<��5��Uq�&���#u�9,���@\�aBu%�Z�{oŭ��X�f|��,J���ht���I��q��b��̀�^AN�X��Xo�\�J_X�a�<û:��s���嫿Jܔ8Rf�V��\h�.�ș=P����9j�V��WQ+��mƆ0��S���:������ _�� A���� M��
,�#�3W=B�4���|M�1���f,:h(R��KʑPєY��d��P:���~��Y(�b����Yj�̬V*�<j�fH|{�La6_nࠩ��� �\Dtl\�j1�gԢ�^KF�ے��z
&*���C�F�5���`���
�!�iM�I<��Y;��P���}��Yh���4�Y5�u�
� 7��Y'ڛ�t)h3*C�������@Tۤ7!&���������p���j^��P��+D�~�B�ɇ�K�����΀p�9����a�A��Oq56�^�m�>�	Ks�5@G��3��~�6�;l�zѴ�����^q���{*:`a8F��?� ��8�1���)�j��l�vZ{��8�`=��/�)�h��������u�Y��IE�',pW:����3���ӧG�M�t��N N��}aW�`J�U���j���4�Lu\��8���?���"�~������CE�qgzo<5��xNA���p�U�JF�m�YB����%#�mw<�dE�9���D��v4��8U,MN<م���徿� ���B��-��?QE����uC<D�O��W��p��4�G��GL�ro�*�k�|4"�1]݂��D����E�`aѳdZ9��4���c�F�a��Tn<�fPj?����U������Npc�¤.�]�}d�"�c
X�$�� :��,v�>�IYLZ�Nl���]����`��i49����W(ǚ��BE�* ������y�@�A�Oa<���V��U���8��?x��@�e�$u���5Q��o�sT�Ш�W/w��Y���n���+�>�Hi��8��Y��!����YKW�Z^}1�A��&^�`snw�~5@��E��m��>��c����Z�h��9$��W��6i	eZ��,/�Sby/f��ݬتj�Y�蠣�_�3�.��O��Ũ��e丛�Im�{$´�y��o�F C�7��E��}��)������4X��^<(���,V��G��<'���'5&N�j�}P����ݑ_a��-m͵�Z���k��:���y�(г4H��[춝:i2.y�wc�H�� �z -���pj�us��\_O�~�/� �F古�>\�uy�m��X���x������1l9R���z�W�l��	Sߠ8&K0%�w��]��z? �_�"�R���\���;���L%�����Y��D�o�0+�כl�`�De�s�����:?��iԭ&bs�<v�E����tW`�`��٣���F�v?�iBo~lt�(�1��,$�
8�-����At[�ϖ�>���@N�7�"���c�/6��t9��C��@�5�W�Ǉ�me�m��h�x�z��r�h����Z*�d�(��6;�9p8B�5��_���<ݝ�B��9�Q�����K��3�>Ҡ��i� E�+�����Ms��@�%<���l��o���Q�^��lb�^߼����ɼ�=��.hdY�T�G�Zf�P1ܔ0�����P�OO��
�}����YW�.peN�N�y$xV���kC(	g���?`cr�c��N5�naR�l�a�É%H¦���:��WZ�	nV~�)�ӣ��e&����C~Xn�tU��|��/=�=�s	vw�
�H���8�3^�y���.[�I�	��� �B������X}��1����Y����m�T>prG[�i�?d�̴�k����	���ˊk��z��_U�S�7��h��"�ҧZnR�|,{E�uW�V|�96Z��i�E>׃�Qu+�2\�]���H��_Uj��2H�}��`�,sI��C{�����gO}Rob�_S�<s\s#�mE�$S	k$M"����8Via�wѓKJ(m#���W!�xNm߆��6�U�l�3Tdۤxk0�;|Ыp�������M̰YG|I�Q���_�k�<>�j�H��b����\����kkD<^���x�l��0�C�P�a&�K�&��s���1�:R�_)]xyw$Q��Ջ2�
�b�$I��vQ6����Ƅ4�� }(��Z�N�Ilm^���5W5�2ܴ�	n�O�m;q���m--/?N��5��1#_�|�:��ZY��"�`ʖL�?�	����(�+=�dy���S�L���
���/�My@k��'��D��o���'��+�ll�@���D�Ilul(����{SZ�=�dA�?t�K�^m��RŢ��e���$��F�^��b}�3��aH��%���U�~��,�3���kzyz� ���]��������<#���!�Scȋݿz�ZM��9�E-�V�L-�+"�Řn��'�Vlv�@�oB�$(A''	P��A@�קv���jo�}ۘA2�w,�R� � �n��־(�F��Z0'�bQ$~�~��6�6Wy�P,�����J9��O�	;��B1j�)��u�p��&���EPЀ8���E������qmh�t��k�c��?��S��ߑړ����{��ca ���raO�b>���l��Xa���$p��AD�����2���:U}oKj�}���n�sǶt�3p[9�h5{Q���6oC �C<�!��S����P�O��rH^��G����G��4Y.��ܷ8y��+��0�z�E3F�[��"۳Y�D���j)2��(FlƉ=9�̓��Am�=d��	���ڄ���<1�$�;^�ݖ|�m�6[y��b~Q�]�ۛzg�o�a ,���nS4��f�%��\St� �������C��1��^}K�=��g�~���O|s.#e��yG��j��V1�X�B���TM�Xf����H�`�~�z]5�j��m�}H�@'����%�iNX� ���'6HbR	��]9>��q���j$<��d0����b0y�����.����1��x�-O�W�I�5XF�(�<H�]+��в�?z��r����=6��P�YgW(s�°�mǁ�50��wwC1Wy����oM����qo�w�2�:��) �VMՃ�/)K���T�1PAz��7o�^���P[f�r��҇���٪D�}C3[���N��Uʎ+b'"�ߎuӾJ��D%]�*$���\��mc��p��T���a����i�ֺ�A;�Hơ��`Uk/��TD���է�����K3����x>fj���	��$Ϝ�E ͼ���S�C�4"2�<ȍ���d
����*OP$���n�>��tw~I�G�r�y�J��q�'cŮ v�r��ԻΒ��i�eO�tГ��,���8.����S1�����{��VZ��M\JN��q`!ýQHX���AG��?��[M\���1�T{�}y�ƭ᜼@�j�%�o� �����}c����:8V���$hxI��\����W��2xX�1�ߟ1=O�Jϵ�l,�0v�������!*n�7C�����y�]�4a��#,���`f[X�:dc���S�����ya �:�̈D�,s�Fv����uDi����s�S9W�9&R�{��:��{��g�+PZ��*������Zf{�E�m�L�9�@�6��%�[B�=z�?0���.B���~7���L�[�).�_ݪvP��м��T"�0��V�B@�ˌ�&Yq�"c˃[�R����Wy�f�H7���]�\� �j�M#cz|{wv򎆘�>�J<����Mj��5�߄̭r����� 6��R�ɵ��e�3���0�#��%"��ST(��F�fW�`���?`~�`^���C���]�p锂�3�az��o�O$l�r��,pw�go��G��4CԿ	]��}�({�5��)�h�P�[r�	�Z2�![��|�~[B�%�sE<:]R^*����A�!�+{v��J���]!˒���Vc�58�&�.�	�#�����7=w)�Y��G�L�q�=�(el�|�ͺ�MHcϥ��<��o��dP)���'=/ZhN�mq��(��a�|0\�Ը��j�1�4��҈VJɃ3��A� �V����L3�T=������60Ur��#4���hU�Q	���3��� `��
l��c�p��� ہ	�p4_�RT���+`�_N��|bQC�1t������+&s&��@	�=,�L*�t^%�4TṄc�.Ud5��K�⩔|��TPS*2O�#X�_�N��m�e�Bϱ1�n7�G�/L·�4|��r��C3�J�zӰ{��U����]V�e��Of�T�u��n;kmV�k�x�&����Ŵj��B��U�hD�Z
�� k�*����������������@�RJV�t�=�XUv��������v����ͳ��5���y��~^�"�`~��ƗO�%K��t��I8�Ἁ���~T�s�kT�2�3'�$��\M���n\Tf�O��ᙒx����Wo�{u���h,��a*�}��w��L�=:mZ|�ȵ�¨��E����2��T�Ր��3ɇ�lh˕%�.��؟�A��F���@
X���h�zsV.R��|šF�"6�Ԫh=u]�q�������?C�|���v��~�M�yصRT
��):ΑO�Հ�.�
�;1N?9���L������x�Se��ϻ۾�	^�|K�%�nt>9V�ۛ�-�!������Н4����Z�$z��g�k6N�����~x�oJ��n�\^��Aj�O�,�����Jp	�o�'�X�'��*��U��f��y|�?��C��l���qa���]S�J9� �|�m������F�d.WA7z:���Oی���T.8���]���G��~����n����v�RV�p�k��g����9��Cm l���3HG��e2��ծX�ʜ짙��&��0MM�����ɠ�������m�ӣ�,��,�"1/n^41�Ys�����9�h��aD���P}�z6ڏ[wO�-�����2�_+P�F����ϋ?]J�-í��>( �����4L�8z��̵H�)����{{�o�ڀ�����Mz�`o�j��p7=��7\� ���x���^6�;�*����	�AR?�f��㧆�3\��K��B���߳S_�LQ^���������L��?��c�J��3����(�c��B�-t�*л���M�(׻+':�Ɛ�0DYѹ�?��r������^���/�d�Y�#�X{r��	`���`�q�i��μ� r��uz{Ү����u���b�[���	P2��6�*����~��c.��J�����[꾾�By܇�OчI�L6��J�rT~����x��#�n0�C��v�6|D(T�|��j|���
l��}h%Q;�'p�"B�"O�:���4t7��H��C�i6f�_|Ջ�noЍ��_2�n�!�,_!mXD��*B�?������wk�P����n��Kq�ܦ8�f��rH:{���^cd�u�A,���J�%|D�+"�>)M�dڇ2Po�	�ŉԅu4��)*�[�)r@*����m�q^�W8$��94�A�.@v�c�1ŵ	�c�݉��Z���͕��񯽨3;���h?�@��T�ܶ�0���>��v��Q$����	ɦj;��0�*��Kzր�9#ݴ�*+f��|����OM�#��3�}#����C3=��HS(m��a�ys�������SL-�ؘ9��-t�h�}\ڄ�^o£z�?�U
"޽4�5"S�-H�i�f���'s��������
u��QA/�++�Wj|��
��|)`�~��K�`N2��3?^�d�z�a{�&R�O�mN3��T��uEcIF��)>����c��u��-��.�S���W�RB����c�&�aO�$��:��l�i__��Kd0��y�M5R�?�F��p)z�u��Ԅ�e.?�z�,�\d��<��ύ �;���U�f��l�x��XE�:e�'��S���.���f����*�l���zR�{i��f�;�_Yd|�~�Q��QlV�ט����m���~
�x�=�쮯�ZIT��q�ZW&�Ze͡�p[���}�����{[�Jm)�2����]>6�I��p�� ]_[~q�/8���`�X'kH����''Y)��|�ܘ�a(��d.��~N^�S7BGTO1��o�%��A����2�q�>���W�f�?�i`|RW@"��H�<�U���ѮΗ&�aW<���k0>2���k�$��z��H=���(�� � 
<n��*r�d3��y{�#�A�Q�C�����Ro��k���N��G�U/R-�J>ʙFSgv��.jVq`k������<գ��X��ß�u�\k��FD��3_gu���5�������d�)<���5x��R$u��*�^���e�tB��	�����n&���Yۥ���@œ�(n4m�am�Y��v��y#��1B��f��Y��^{���3�� ��=�= ��1�Ѝ�߃)���$Pp����
��?8�$�pI��?�Pl�9ȑl*���"
��5��ݭK��ˠ�]$�"���z�����&qB�S��O �q�0
�
��Bj�H�m��+��ו&iN'yY�-#���� f�<In�C ��BO'��3���'��������0L:����q����VDfv��TX祾��L225��ami�Ou�R�p��)w޿�R��'���
2���h�CӞN��X��iZ�2�	�d����� ���3�O-�
g�+X��'� �\����$%\��(!��U.|GU����S��5
��h�F�D�����3�lب`&>����j6�츭cl�%�����[�˩;/��7�Q��I�wnJa�č|��;��h�D�!|���R��͍�}{5}�'@��m�D �&	m�zN
'�}����6,[�[<�y��ba���[�
$=;�iA �P�!��a�?r��e�T�ɚĄ\,�C�̜Y>m@��S���XsGߛ��f���׫���O��#�$���Ӆ琴sT��oK��W6���YIFW�me?��\z��D�~��R~9�r�G[1z�o�NcOv�Y|M�;����f��W���Ns|{�q�#C��F�xx��J�RC}��%�,(Y�x	CC����S^�`�/�ɚFG�0��U����9Aضvƍ:�,2���M�����
¡�����Y����uC�U��;����Ѐ*�SY��[�4���Eyu���L�a�X��O}S4���V�w��"��q�V��OR��w7��'=�G&d�xX)f@�Y��}���p6��E$��QEL�� ��>�3��7��C����m<����>Y��Q˯�v��R��H�PŤ����)�l�:s4m�>DB��w������P��R�;��N8�#pM��`f��zQ���o��t	����S��"i��{:�
]I?{�q��g�� S1�|%�q��9+���~�q��������D�;� � �~�]�p����$��-�lI��1��	0+�c��_p�����\�<�X�"��|��(X����ѤS�En)Cť�XH��
-u��	��SX�Z��MN�@�+N����$&3F`���rh���Z��RSQ�.�j�	�Ş��`/�+hc 5�s@m�+I���>"�}Y���Eo2�}J,�����	����Ml�����X �Ʀ��L>U{���u�*y��Ze��m��%�ڈ�W[:�V(y�wf.��.��,�ί��f�� �wwӅ/��v����)�?麺N�Ia����RB�s��k�'�~�9���S$�y�� Z�I�s>�5��<R��J֝��嗑��iN���he%J��º>~z�����������%AHv{<|7���
�]��DLK*�^j�_D3tmχ�SV�Mj�Җ�\:�Ě���[�4���obX�p]X���MB0�ȍ\�y�� z�WB�
��j���I1��j�R�����V�5蜴�������cO��޺�f12eS'��c��Kd\O�x��_�|���joK��^��?l��|JR�)��#�3��;�ȏ���; �Nz!�x?oB����w�R�;�1���P׶�U�X9F9FƁ��y0%����1g����X4�ܡ4;�ń$@Z���@�3�L����!)��E�"�>ar�ށ>e�X矇�5-��T��V�E�άB>:�&؋͸�V�[�y�I��pdHqTK�P�,�`9(��8�ކ�K�#">1��-��oK'!e�,����wx��v���[h�����{��W�����N��xA�(�A\�z}��� �8��	�o'{�-	|��ݢ�%�IT��&�<v��w4�%�hz�I��K�Xf�;,��,�+� }v
���䎰��9�9�S�Ȱ�+nǭ�(l�-׮��Z?
v�D�+n��Ԓ��n��Z��M�>��tz��p秺LRw�M�8ae@P~y�f�+�A7�^�u?�},�� �՛xB��?80Bt�-�	p��4�43�b�!B�_xa͔T$8ͼ�DF�7J\����6� G<�q�+�S�tV��_�L�_{;�U��<i�ez(�0���1�Qc���_�=���BCd#A� ��"8x��{�֎�d�Y����p2o��KC�.'�Bh�>�����`J~�C�In�1�T>oр0�5|�-��<H�Ʃ��қ��s�
�A7�
zFz�~J��b���t��.0M�>�\�;���������{"�Z��d���҂�Ao��Y�O��ƚ��F���co�)�_�b��6��{�>��z�R���k�?�9]�*�#"�G&�-��8�y��JטT �t_r#l�Hc���c�:�f�Yi�pP�\���ەp���)eck���|�� %��� ����5�V����Z=�G�^h�)֒n�אi��rp���9����A]�~�MT��,�	+=��>�ʁj`h�ө�r��ZlԶ[&=��~v������L"�J5�@(�r��ݷ�QR�h�?��X��\D�|��%�8E��V�(���:͌�D�x��ޖ���:�νԓ
R1�- ߔ�I��ܬ�yDS?8�H�B��]r%��I�*�>\��L϶P��ն�����0�����*�>6�k$�K���#Њ�pÎZcJ�c��gSw���͐��G��&���q��{9$xKަ�V.�?�7)��;�o+�{�E�/F�%�%���;���ъ�����yF�+�zߎ?���� �;�F��2դ.N+;瞍)��}P�v:���Ҷ���� ������䣠���V�&ivB�?��c k�O�Q7�Ö�,�enbF{��bMY�F��� Ģ�c/�P:i�A���ĒuoHF�n��+@�j��7�˝PGc��=/��:�p�a��c��%� Zwf<�ACF^,����*O����ګ>}x�0e��
!�Tֳ�G\ �m��c!] ��?�g˒M`[�4(w�)lB����5��ˣ!Bc`�j��P�����V
~�-e5���0�����	���Z���-WW�am����/�����@4kĒ��X���N`k�b�D�?S$WĆ�,���\*�8�ӌ(��*�AluJ/�x�wf����'� �ѧB�`|���$�`@ٵ�Q� �l>\��AG�]E�jy^0�*7��@��aM&w��1�cqI��DT��d�+�8�M��"8ߗ�Z�%�9(++:�
�E���'@[
o�fG���Ȭ��Q��m��.y����!�>�XA Re\��Y#T��	e�},h,�#D���ޓV f��*����_��|!�W��.�s��<�+`ꍌ�5��+��y��V,,_FĠ^hᛗ���ڭ�6h���c�Y�����w ht�J�w�%�����|�KבC��|�>�Y%���`���}V�%�ъ!��v��_�2��i�Q��
)�R��@��$)��U��Ϲ�<��1j�v���z^�?�hQ�֊g�(#����d$��]p���p���>��A��g�|"(��T��"Ց�� ��4�
]C��#.x[��4z�ޝ�k�	��(/�}Қ:=w��Ç����))�v;�7zB�m9|�M�a�������F�'������+�-8p.uN�k��.���<�-~��`�0�)	�&вN�ES,�`�����`MY�i2�I:\9x74�T����wFd��;�e��K��B�*q74Q}�����Ƴ�a��i�8�6f�m����O޲��������C��s�dEu��ul���n_�|`�g��ڜիqG�(�^�B��t��h�Ȕ�F�B�/v��ĭDB���E�&?�6��`ʙL��7'��0�	�P⎗����j�w�O�*B���?�����=��0���c~e�h�=�8�19�nU2�ꍎKFF�@�yL�l�Z+x��aCMC˪9��,/z��8�*}3�o�硸!S#T ���WZe���%Ӆ	Jb�Kgi�}�m��>*s��b�F�q;3�*�_��q�۷��]���Z��%H�Zc�椾�M *�uo�f;�cle��K���tA���)�[��w����m�Y��@&d��k��f��H~p7q��e���ó�z��r�Q�'�E�c���u�g�5v^�m�2�B��y��^\�(�A3��Mrn�q/�V�(�G�x�7
|@��dz�>�U��Y��+� 6����������a��n߭����J�
[��Ә��%��ܭ�L���v۾��K�?s�D��%���A�9y�j䁲�|��O�6�N���� 2ͧ6��d��J��N$����Q��f-���#��T&����MJ��G�d'+p7Q�,gp�[ɓp�-Ѷ����uxO���u�ĺPՍ�Jk@���jvH{�%dGS��c��:����0g�+�M7_�;���g��.�(��mfrb�E�Ǭ��?��b���f�@
�(q,�Rf��kD�ąن�4`\kKm�V��c��T�����/�MZGm;|[񳕂���$��l	�Xo]4�ؓ�C�=(#�b����Ġ� ��2�^MLה�P��Ν+����m�Tm�ďnLD��@�/.�~�-��󣎁-�[h�f��+U��91��ˍ��S��k����i�����b3��c�W�@w�t��%��I���q�̩���k�������Q�ǾT/Y|(���&S;���f⿶kd\�S�^Vq^�zG&-�It�G��>`.F�!+6\2I���G��g��9����|��A�H��P�8V�ț�>~�yY�x�t�ٴf�ׯaZ(��Yہ�S��>9�e�N�}�U.}$#�B�?���]�NW�2Tq�Ρqz��� ���v0�����6|�:8�� cs����k9�7$�"%7����İ<;�����3�0��6ؒ��΁�>���^��f���dK�)�U~`���Kq2o��'1$��`^7��^D��y )d*�}Af���b�M�B�#�����A�6p��p :��a�\B���[$�WJ�)�w�%A'.
���[m\zvi�1#y\��P�Ⱥ��;�G��;�e��d�0�g�J?cKUCf]8��\�di�\I����X#YS��}�Ƿ]�5ȍ��J��� �2-�8ɭ&�>d�����;z�AZ���b�盩��+Us�dsD~�m�:���c��:`Y�Σ�W�قuyP����n�=j��8�jV�4y��|��ͯ@|��謅�O����V�N�jg�F�5t6�V��隟��.��B����!���9����NV��T�V�
ax�qܽ�m(�m-o��|��D+ ��� ��,DT��8-��X@ ���v!�߻v��G3��P��₿�n�_�`M��(��}�9o�FAi�Z����e�T�TBӊp��A��L|d�|�pMN����si��IB�����@)�O�vd'i?'�1��,�`2B��w���u9����Uڌtľ��-��p�T%F�u*|����?�Nm�
����`��%�����B�9�y0��5�#{\�"B�%�|�����W$�-��;�25"�>�(�.��}�a,��~u 7���
���d�s���y�d����)ׂH���}A��"Q�#��]��1��������G���,�7.��W)ꄼ؋�T����vVT"��T���]��Kmx��W�U�t�9e>�K�;���w݃,��H�i���-=����t𙆀�Ɵ�ud�� ���� U2"�i`y!1Alr�Y��X
��M���@&z]1~��#L����ۏ':�"#z�-�:Ӳ0j���,�g������x֊ɯ��H^��΀��Oi����G,ol����^��z&�+<A\��Ͻ=:yl$��J�bo��R�<�p�y5?�1�0���4
�,ö�5~'L�ء�J�p�9O�"7� ��K�/�B]FX�0}9#�G��}ŧ�,����Y&��Ԡ�u���Z��$f99wס�i���f�z,�N�?�V�f�����+g,��:%����>�x�K�7�l�t�Či3�]e�.���3�J=@i�&n��;�P�+����0D���b?�qa��c�C�*׀�h-���_.�$Q'}�m�;�lZ��[c!'�/�K��N���t,LX��C�khm�`k�ꈗ����3�&{0��,���V
{�Y��{}'�
�Ѥs'zKϡ��:����-*��/�¼×���j�S�qnx��؜a���y.��c�,Ix�ǂ�CmQ��)*;��5��p�z%���vazxY.Ӫ�2��)>F%�&0�@��KP���7�����N��ά�|�t�/���v�؄N��!z\���`�����4�2�Õ `�O�!%5�ݥS�:i՚45��/�̟ 2
�F��I�n�7@HZ|�.�5��ۼ�Kا� �̏�L�3@�)Ȋ���9q��w?��N4�[��+3�y7��h��J��Xf�6��@�݂/�w�F�GA�AH�yt_��wf#�@�4m՟wn ���E�lnA(0�������g ��m��j�T�[�E��	Qe\Q����� ��#0��-�=�u����ع =f^�~���>�1K��6�3��vH�U��4!������Vo���uǬ;=�n8�˿	��I�ՙ�{Q��d�}U���T�]���X�&>m2����w�^�gS%�@{�i�ی�q$��j%�%�ш{��G�A��d4�pJ�X,<�ǣ�ɰ)��u
�pT�I]F~����=	3�t�_�$8-Qr��
�`4L7��d�ܱO��������*��-x���3��lP�!Z9h���?$���_m�;��yĂ"k���L��(A�H�'Y�V{�v��.�4+1|�$��T��$�9��gsU-�U�#8\����+5~f��x�T��JoY���k@�d��t4�J�5����_(<�&�� o�23`��Oh�εѐ�[�?�����^��hI��/��e���e�s����m��U?h;�h��0��%=��`0��ػЅ�V�\.!� ��X�Rj �M'�!��E�B���
�y�ꇉ��A8	Q�ū^��e�����_A�|�Q������meL�IEknp<x��\�j/�J���|�8N�D�4��=Zl�A�:SӜ3����6ļ]&��D�z$>Z���50���VS�ڪE2|ܮ��ILJ�;�l�E�����L�~�P!�1�_��Z}��	�uUt��`r��f���N��Q �IЮau��
I[+ Қ0�0�K�ma�0W��$<��rG���tW)rV��2��<��e4O�K�D[PJft��GCM���+���Ğ_��$�������@���ؽ��ﾱ�]���6D-�A�v��px����K;��1�m��?��Gv�//�s�ƔYK�x��k��[��܆5:@d@-;�@㠛��+�!�ڟơ`������z�����ց��"�(hjs^�b�fs��:�#��릸:���w���4D22e�!�c���ww�_U�̯b����O/0��|��W=���ـԡkY�O�^����5b�tɌ�B���!T�{��`Xkq�7[�y�^0�l�'��d�PN�F�lh��0��-$��iad��c�
�_���R�-[0W���#OY�V�}�wn�� �=���g���gAC��X'�h�F���z2n�B�����Xc�4Q����7�%�)�?OlZ�*����E(P��P����R\YȽ�&������?��6%�p�d�g��7�7���T��l`��ioU��絸 �2m߆������'@��QX0q�Ai01iSǼ�Q��Ƃ&��_��W����@FL�T�(R��Ψ���4Z����PCL&pr�ž6+��~d�~����4�sl<T��N`ɜ MɜW[ϩZ�d�$w�I�8�,�4��@і,�P7c�C�w~�<u��^E�[��)����� r�������U�}�|�M���h�����"�9b�0�9D�s����q]�t�����=1%GI�� ��l��sn�����~@Zp�������K���������rg����\��HO�ǯ���R�m"��8��q́�c�]�H�p�8�����J�ؘ�3��Ҥ��V��4ͣ�3_�3��dYF~��z[�⨷�I'��v��:he�}K�$(�r��Q���klka�(�/W6��fA/Fݣ��z��a��T�%b�Ǫ1h�PSr�T<��ub��U��������w�|_�/�W���j��7�A�?�Ƿ'��D�HgE�a~&������AKY&�Mf\�R�E�z'���r"�(G�|*-:���E S5�-.�x�c�&4N+L-j�f��m�|o���-9P!��Z�'(2^G{̿�����~�Z���{����?0}���u�mK�\Y<�;�[���u2��BL�"��C釜ɠ$Va�^�m`�NK2�_�:��k�"�5�;��GtȽ96B�Z�y��>�������CX�?b�K��>c#4U����zxEKM�?��J��џ,(}|f�n�)�[�z�Au.��n*�7�u����&���%�pZC��v��F�����!��r��G�o w�Z�ڵ�{5*5B�K9�|h��Ӷ�"�"`��Z��o��G��¯p	����B��@��%�V/��{Ej��]%T�
�@f�nPh�-�s'yN��o�m���.�m`n�";᧬PB�>�*�0����c�z����	�\3K�"cՍ���5a�~�`#�S����b<�βkp��r{��?����1Y.`�<c�$����[�KD�n��x���y�5�Kj���W�fLc §%^�.�I�tU-D�gǿ��$'�|���=��pWE�qD��3��20(5�3��
���lW�Oߞ�.C9Qa���*^�b�Fٴ�<AKz?�j��\�(�����G  �ZM�͒��M
X�vM�o0�:�@Vx��;#t�ɟ��>7�� �qn�wE.��V�D4�I�@�h!`��^Fqh{�	r��Wa�7�-ӉEm��3#���Od���i�!}!�&6&3&�����"�0� <��sΤeo�f }ގ����ҵ��ir��!CE�d��FF�q_b��d�L�cs$�cDO�/����'�m��$f_4>�\�@��-��l���+]���Q�>0g�pd�����s��w��k#�2F�6�a#�c{n#&���໰����%t�k,�2|�aeDC����|�Q���k$�%2��\��Ӎ[�n\>m�V��w0�b�����gB�Иd��4�w�s��|j��/��i���+u �j1Լ:X�,��,A���H�sP�n��r�'ZGҸ��Fp��ֲ`3é~�P� d��#���>��)X 'C� l��C���s���$�?̮�b�W#��D�me�CM����4f�uJ�R�[O�-�6�E`�N����}E���|H����1��zgjđ���`�F�tׅ6 P���HǼ4��Зy_�>a�f+v���X��B�qP0�uY垒��.G�ڀ������+L#*K�as�v;���e�J����:�n��@[�с�C$(��D�����Ye�^ 9�� 4�x�V(�[�r1)I��f��l<x��wid�v��O��T@��BA>�?ʔ�/��Չ'��-��i�+?<S5gl�v��z6O嬨��\C�K�Xڶ��o�I�H��6�����Τ����ˋ?�^�^�.ϱ@�#�'"����N^b��F
q$�!��a��3��yJr�{B�/q��5�Y�Z���.�(7� ��_>�Q$e�y/�cV���֥��S�=����"�7Z���>Z���s%c̀!����oD� ��,�Taw#��!qA�3&�c/lj ms<���1ˑF�oad)�r��@��y���88.6�)���U٨��_����Ä��~r��2_��
��h��K�w�����Y�W��b�{�^Jy5�X5hu��lh��~�ƚ��ftV��2���$w���C#�zҞ�U9جr��PD��nZ4�g�/������p�-�s/��-^HO��3����M�����{�?���+F޳��FF��f39��H�N�yGo��+����[�'l���Q����� ��<D`�ܿ��S,�>0���v��֮m�zU������mM���@cŻ����L���B$�㤩s<��)f���SV����d}�u����6�� �<�m�kq��>���t+!��?���n��3����`*�x
���k�=�e��C�a�r�pV:��ݷ��<A�I3���dR ��1��3��
!�s������s~H��Y"9��~[.�BXJ��^~L����Z����sW�J�B�X]�In�����B�;�T̗�Y,�c�ugc��xwб\���S�%����U-�w�P�>I��uj�J��:��偉�1��O���F_�I�nr4�T���ޱ{���Z�0|��>��lvXQ�C��1���kՅ �W�Do�OΝ^d����Tw���S���U���^YR��tC��`���ʠ[�K���͐dd�Jqd���<��~-�30��dڒ�د�Y�	��nJ�źƟaM<O����2��G��uI���#�����O��j��HV6���o]�D�p�[�/x��"m�f7+��,�!����A6_k���l���5A\�[�����h�"��'E��)V*���M��R�r�#�Gy�O�� ~�V�O��璍wr���B�,M_�3�ju�5B���]��l�������)w���*-�QQ�&����9�!>����il��>c��ﻭY�{���K!�ѡʡר�	V�B��;^����Ϳᘲ�2&1�2���:*�ʅ!~��s�'9a�'�.k�(����*V�H2��٬��ˈd���Y�$�0���=��8�*/YޚD���a����G��/�L~���'�o4�!c������N�U���s�쭺�T�wC��|�!<���dw�$���W04�6��`_��\�� k���ya�|��B�B�H�'6d/���ʈ@7~b�f@��gz�V`����X�-����F����-��u��hm �hd�F�{̏���y��a1l��ـѴ}��O�|���O�c���5��bc�}G��Ӽ��ph��0}�D{�Ȅ��燾�{�j3a֟�����ϱ��R+���������	���6A<�l
��b�e��@��q�9j�շiy?�ϕ���[��bl  �2�U��7�7v2��$r���~��dŧ��K`ʐ�pz)b��R�)֐@������Ӧ0]�D�ba���1좚���$�5E�pH&(��@�s����=+��C�[�_�d�|X�a�{�����dR䳺�W���HyB��Wh��?*��������[D&@�,��+=� `W���s9�.��׿m���Ewlc9h)�_�d[x ����M~����P�����J�xZTՅ�:&X�������9-� >g��$��+�+J�P�U�2>B��ͭth}�A�b=@�Cֿ�����H������D�vip9u�	�6T�{3w��xyB�����\�������)� ��ą�)lt�$�A@[%�5~�J��Q��'ы�' �� �Ȇ;��h�4��/�{U�r�����z6w�΂�+�4���L�Y{���9/�H#��X�{|��S�mH*���">�-ؗ8�E�yBr���Ɍ�L�g�>4�q��XBcB9���4�!�x��I�3/��7���	p�&�z6�^��Q[c�{�pepD��(qj��RO-���km�zK��ޛ�.���}qwFk}�q�ƨ7��K��@E�5-�� �M=��v��A�g�=B��X��D �]��YPS�����vף$P�D��<��έ���	�7v���H�)�{�#]<2�2�H�R"AC
(���Ϝ;�v��l�B�Y�)D��y� V�����N��d��ja�<��衈�SD��r.�g�^��[ W��GC���aP�F?��3o���L��iQ`�W|I�W&Y�/x���lם�i�d5+�e��F��{,�ӳ�*��B���25$}��/J���Y_ώؐM�H�ϊ�ˠ��$6
����^,*R>�i�=����?������T��?�d���+��߶I|_~���r�%�r������˫��X\"mT���$���;؊��e�_b����oH�c�tƝXN@ոۼ��~.q	�V	�pG�ѣ�`��m��������%�����;�Q��l�M�ޠ�A���(8
X�^ٹK׌�����%�R�DG���섡�A;9�ó��d�X4ϵ�N�*��' N8�o�#��B&�Tq��p۷��/X�ôB�Gɶ�l��&��ԉd�`�nm{���,�<v$N�;e-;4כ$���$��d��^yo�n� .������*#u�?�-�FS�%3�yV�ξ>���犞�㹀��S�i�}�
|>q�'�ͮ�Q�^\<�і������������>o[/O%�����)͞�d�w���R(6!��Z6{,(��"#��["p�V\ ��d�i+Cm�hqNxO9y����z�D�ގ��Y'��Y��z-+x\"���
�]-�E��6���l�$2�KǏ]��s�1�sWz��u)E@��p�2r�ET�	�q|$'ΰ���o$#�+��~�|��[�tB�Bj�(oS��$���q�c��V�n7������?�k���g�R�Cx�'�>�����C��q��1ʴ�'�yE�ކ
����E�o%jR$�l�W�d�s9m�۩����#6�ɖq'�@��<dosn����ͭ��t1�㋐����m�R��}5I ���P���9��g�[4tްU�I�r ��e��	'���j��aś,�G�`�6�T�7�FXH�Zԙ�ƸC�i���Ϫ�(�ŀ����o0�l��	��8�>p��U)�l�$ �B��:!���B�ooZ���� ����b�鈻��v� +�g�|��$8h������ ��y���c91�� E+�,?)z�y�_V�f��]�[b��0F�T� (AF�m�%�^@�0���JW�bvj8>ϸ;+�|�����N�	�z�^���_Y��}W�D�j$�X3�d줊[��^(��R���iYC��=fz�pݜP8Vr;�8�u?�i�$����b �r�X���H��y��Dq�OߓUl6p������=?�̛��o�kY����k�� �?��K㞷�ǹ��+��]�X/�0Q\cR}��'s�϶2� =Np��fF�ڢ]{�� J�d��j��
�O��?9uk�a�F"�]LSx����Sǌ�s�y���=3���),�H>�͡-�6����H2MA�3�s�F�ʉ\�y�"kH��1�z��?�[]	�r�����>��]L����-��izJY����G.�W��ܩ�������ݣ��䅢��m����/5P-�w�*��F�z.�[�m�s�f�R��+��:]�x�{H6�d}�]�:�����N��¢����1<�CFS�g@��	I��C��S�>���ݮІ��0v���"֗PCb�k` -�����̜{)�X�p苻N���Z�BdO�c3x��D������ּ�=�}[��,CgK�;[�w>eK�N��u'��s�R��'U�]`�����I�漪��,4�I%Ï�N���C���1�6ƦN;���^)G��\؂6Eu�j��Z �I0C������I�w�>�ŘV�U/�4�G/��3U�UsX�W@a�lN�]��j�@y.����|�&���9���U��|�)n#��(1����e�4�$��4�E�t0���{�����VLl������
%�p\1!<�DB������BG�����噰K!�1�f{U��u!^V��CH�	�~���k�����C����2+���^[Jj�Cm�k ���d�u��q+:��m�\��_�\�W��0�y�i�
I�ԉK���C���������\dP�K22������׻�u�_�\R�gӫ^>&�T|yǫ�7�-"\Ĺ���0�6Z�Z)�E����᥄K	�Ao�N���wߍ|%��Os���t����Y�1G�Dv�@�I�G�!���iC�!�x0פ_��#��o+���gy������*U�P!<�C6���C��|�x>��Ng��A�j�W��
r}�������G=5���39'�*	i<�J��]!c�8�Š�t�	3��9Nj�(o ~�u��Lq���7� ����aۂ�,R����\��x�R>�[��.���*�t�Ǒ�S�8�=�\KGhԱ��'u�:�c)�`C�8G&�z��,��Vg�N��f��t0M�Ha%c(��'5�ַ��c�N=��/&2���x.L��U+xXU�Xb�W dFtL�*�q����47��ý%�e%�^R�0���x�5�ô*4	����$�3�����Ct@y� �o(��bƘ�I���,e��-�����l�!{��
�"�7��|5󢲢SjG���ɝNS�h��D�X_�Ձ�V䱩u	�<���v)�L��s2�b��QdM����B`�W�_ ?U�U���9=u�.	�AބIė�+�(tzB!&k��6���`)��!Fl�t�|$9��{a�a���E�Z��Z"��ql�u�bBKt�A��Gÿ���Єӡz����<a�`����p�ڔ��B���;q����w�>i�:��m�=�,ոq磵Lp�@���/�Y�qE�H0���|;���%1���B�kg�x��~p	��~�h��{YW����/�O�Mh�bn����]�3�R�]��9������<:�ږS�-p@�d��i_�1Ji�x]&Y+�Y�n���U8���pr�u�F�&���<�_��Ur
�'�o��]*��:�������6?MR�~<���ZA�8��G"?�׺����n#�ͻK:�0�N�%-�`9�a�@Wʫ�/�E�.�j7�y�L�m-!�����-?)kL/�����2���y�ͪRd��ו��E�\��GO�>xa3l�t��4wXy��������Bhm���-�i��hT�pg�"�G�����AO��Z����N����s,���k��"�5
I�	d���x/Jv|B\��"#VE�C��l�R����
�\t�������7�ϣ↧Z�Rň��Xa�F�nPw�剦�5���}��۾���r�#��%j��ՖpU��sue�/ `�����@�y���4ǈuլ��7�O�?����:"���;n�"�Jޮ��$�~�@�&r^ �nb��h&dT�f~C���YnC�N����ݮ��&"+��2[Yĉ��V�sbڌ���fW�������{���AR���]UNK�x�%@x�a��ę�q$	�z�������;��i���,�lˡ�8.�n.�B��/�!�"n ����T�vG-1��m���"y�|L/2Њ���f�yc�m�7#K���hi���Â��wo�ƞ#�ڸ��3����Hz4��}��F��m�:tK�qԤ�L���f�݃�t���F��:ga��*�j~R�4>�*��D®�[#s���u�!�����w�~<F p��4 1�y���:N:��q�����o���mF�i�hti��a��(w�>�ʉ�����T�q���o�W�b����~hy�԰�O�J͘d�Ԕ��j�{���|��1��g^�{�^	����)|AȔ�ń���¿�@�씽���z9�D��C$Y���.ݭ7ʍ�_�1�`��GM&�2���K�E��%�e��u��KRn7�c��~�f?o'B�q����kƷ�Ѕ玀&�2��13�tY;�kղ3��,�;�ǹDx74�~�u��v���,Z�ů���`{NY�Ӎ���&�Ɖ]�5�~�o��ۢ��
��59�3�g٫1�\�lC��C��f��X.�����DIK̯�~�b|�7R��N+����@8C�%y��%4U�$�'��2>��1_��[��D��ǃJe�H��]�p%բ��6*�guO][��﵄ ��*\��PtU!޴������_���_7�M}�����9�G�<˻[6�����P���"�D5�z=F���^Y!8�����Pq�(v������a����v������¼`��X�I��Fj��d}힩O�(Z7��t�3P���W�r�X0
���[O4y�����%�_��/%�C�+)� V�E����f�ǋV��Τ����3�Q������@��A��2MF|?�\�n�Y ��pǊ}��¯�>�o&x��#�d�d��Z�[�!!��_=�ԓ��	R�|���D0���ɰ�k��|ߦ�FV�������r�I?�u�U���F()��*úq:�ģǷ�.rB��DoC���Oֳ�s�I�'c2��*�tsOaS0^��/�6t�C�m��6�q�h8u�3��iX0y��&�0p��L�4���W�*.���/Q���}�d��$��	p��ZU��NB�o�n���5��/�o�zE�a(�VP�,nh�nY��^ b��n�%���8����[e���o�7������
=�¶v$��rn�-�):��uH����vz�7�G���P UP�R�E�wa�طc:
_�<�TX�!}���BK8������M���;�	G�A������_������)^��7o����bB-p�a��Hd�"9�{W0J�igB�O�l��KdF,{
l@�s@�8S-e.��z��)�=�p����<%i�"ǅR���`�&�;����X�0M�#���V��m�m�.P��x�����<�O��P�EZ���W��d�-wץ�]om����߽-���|��<]�\��6�{�8����B�L�����{.�O�g�KN^i,�i�Nd
�<c�E^c��"CuNRڃg1ᵑ��w�*NOc���I؎'%�]vM_I[C��ؙ<! L��������ǩe5{FB=b�i��#�h�Š+���F��v4Z�~p�B�P~[��b�B�i�2�(L��R^!!�9������!�_|��V2:��9����HΙ�`�?���-�}�H"<#h��t�9��
[y�o����U'	7�j�d��_"�\��9�+���6��~M,+,�)n5*��e�]������pQ�Y�K��������Yj�A٨P���/�����B�[�'�v�	��*���/;���R���N�Mȍ^�[GRYt<]���z�Y�-�e�p���=xT�����ڈ�V.�G��bO1Э���wh��4O��Mw�|qv*����j	?#�n���o�{bb�˱0�b��	�J�&�I��I�^GM��<��WfN�W�?��/��?�}b�х0k�0�/W��b�d�.��*I;X���)gyJ���a�3)��V�`]�ɆFv!yG�b�)�g�x��C8_��Yߢ��� ��U(g�R�u��L��~|c�@�#�3N��t��� MQZ�^Z��vm��s�
� 0���7����u���!h�. kZ��\Q���]��� �q#���9�N�)]��Ku_������3�^��X���e�g%\���}9D~.�?MQ��P�	V��4? At8f&/m����-�GD���l�m1p� �H� ��oٺ�*1Y���E�2@E�j:��E�"MIC΃�|`>k�Hq"JD6��Û/����e�!2D21S���{0R��P�L'�؅%iN����QE��U�O䂑P�U:��t��Ob~��'��ᒝ��[���L�!�f!���PE�a{z��'�]��W���'�\��>ݵ��@7��7�PSY�|��>�M�QX'?Ъ
�H������)s��-S�j��6�#�6�qJ����_3��=���˙ޘ%�sf@[����V��i��4&}R�X�(��hXx�5jzN�0(�)�dm�_��z���1���0>����D�g��>We��m�x�n���[��H�˟���ļ��N�b��:'YNŊ�@�3�``l����:��x���oM�������lO����p_�!Ubo��
�D�V�h��*�������OI<����ZϬo0�	�1k���+֤����ŧ���T���(!~w>�±�W�i� ߌ��{����:a$��7�<�����������0�v����a�?>��P;�Ĭp�r$3%e���L_h�μ��EA��|j�L����h.Budja�!���֔'f瀤
?:��W�xb��Z��3���ٟ���9$�^�!�b����!tVց�ŏ� �"g�Up^�˝��5��#���RL���h�����7Ԭ�c���j��b.��}���0�CM�q��6��5��d�&'攬���Z*=KܔK�S-@,H�-���e,��*˯2�&��o̪d����=_]eJ�M���h�!اͅ��⁨��"�Qh��zmf�ӻO�%�[�E5��MM���g!����M�`ZS{��K�uh��	��?�7��t��ᑿ>4�b��ӟ�7d�PHݲ�RnB��VB�۳������7��q&��v�^���寄- �&���>|��H�܇[����cIk �hذ�~��AyN���ݴ�x�1=�7	c��փ�N��d��δ��m�����i%�9�22�m.�`QI����I�AP!Y
0p�&T�r�8[�ڬ?s���[@�	� �l�f@���a�]�,�m��
WJ�2�$��ЩY=[�Ƥ5�� M<����%���*g�W����5&����ݶzނ2� d�`Ӽ�D��˔�2J�z@���t���1'��a�u�%��h��B1�h��3���N�Ӄ2�:�\"�d̠L�}*8��I��Ч=>�c+���-�g���$�*:��p�ͫ��'�Qg�>^z����5C�V��>{�ؖ��Z��!��w��K����x�% k4ӅPE9���r��Y����,�M����?��s�c��rc����%��lR7l�54N�{Z��_��{�f��B
�!�"� p#����L)_b�Gi@�o%O��q�B1jފ�X��.9ᮘ��s��6�R^T���KBV�����s�}ͦ��^^oޣu��jƢ��c[L���Z5LE�"U�l�{��Ro�ѷ#}�������Ws; i=��	H�N�'`��5�ּiFH΀��������6h7��çYp����4�XGJXd~V�(9�7 �:���>k�2)�r���Z~OP�:��VYd��H��9���QKI��HR�GٲY䣴����<�eNz�N���]�ޖ>�R���� Z	mv���h�r*�Pg�L�\�y9i�MG��S�U�T�8Sr�KP؝@�"(>3�q���P���2�:�y��
	�bOᥚ��4�XE�>�M6�+�cB������2!9{#�b�di���9X<f`�Cu�DNثj]z�h�[�H��x�
R&_��G%�"Ƥ��~}HA!;��&�S^�<�k��eɂ�l[��?�@�=�"���vEETGe��I�-�v��0,a�";]b'��Y��m�=��`��u����)\�f���
��h�OF	k�}9h�0by�)��r9 � WԷ�EW�+�B��^Ɲ�P���u��ps�P(�\��@چ��s��V��M�8=X�oo��Z��%K����\�Z5]�3�m�Vle������ڳ�"�L#.Ƭ{_�!%���?�P��g��\'-p�Z��>�߳�����A�K��yIXs�k���sr�=���]"�G��	�q9L,�{��V����
S��e�� r�t.���+Ogۀo���#�u�U��@Ͼx��TW�W�z�d^��0�� �{	���Xb��U
�I��f���@�O��g�L�>L��}P�}�
��}��w	2Q/����K"i4%޶?�Ii���Ci����hw�����������?�K����ГIC��]�.t{��߳vm�� �&|��%01�S�K�W��rH�T ���I�ұ���3���!�8�"��*�0��q�+�{G~tΗ�L՟�`^��R7|T��k�����&��V�#�77��g�����Y~�<���Qà��QԳwޫ<ħ�yN�f�cz���%�ǟ�Z��a�c���yO�6�o��Bl�d��ny��[�_��K�!�����g"�eR&�#��Y2t�ʔ��ol��k�*j-�k�`����kx�&|B"t1����w]���S��b�n~`��f�$��W��-�(��q�w���>~"��-�yI�{��	�?郢M] �I��#.��qT�*�m���|e�]���g�n#���}C���j��8�&ϗ����4��B�_�t�
c��z�25^��5�1���WC�v2�
f����K5�_Xtm X��k��ݥ�� �*r0Uk!��±��V�ڝ�ãyd��!�p������<�Ŭ�U��i;	�?jU|hYa���ᣒ�����f�.��-����Ѿ��kl>���x�����~
� ���,U��J�^�4�-���6Oc������X)���s���?�j�az<�6��4<��!//$�O�9؛/���7�N�/j�{88�������%�fhA���%	l<��̗)���7��������SxSŘ�ʅ�h�qX���:-i��,��M��_�4~������zn�d�9m�΁ц�*�S����Fa��7V�ye�J��d���@�?r��lNX��ݼ�X��B񆢺�2}L/l^�*�tgb�d]6���� ���M�����~�	��|a!5�|� ���3LT��
q��	¡�x0�7w~칯�tma�K��2mlB��_d[F�J�]��wTî�ZVhΪѩ�%���|&@S��fy8	�F�[O$)G�����H�)1��qb��ގz�q��_�m��w��T�X*����Z�~�cDI�z2�AQ@�����{�E�bk,�DX��ے64�:[���3TM��(����WZ�T�;�l+�nQ)�6��O�� �0WE~�U�l����]��l)p!��Z�E���G�ǥ-�kw0 �o�%؉�-��;��z�N�T2�x��L7_h$�NL��*Xԧ���ݘ�q�TK�^w4t��>�]�=\��#cd��k���`>-�<�t��h�h�*�Y�WQ�kV)�#bg=��T.0q!�rb(~Y?"���syӇ��מG�dw�za~nMtY�B�/!��������I��Ǖ;��`���HD-��HZ]e�qa@*�y��T�XkӢ���vm�m^s4멢�=c�z<X�8�@r�rA�@����$v�?�P&�ݖ��������GY�l��6��|{b�?f뇝�0�U�{|~���Ki2�Ё�$Ǆ�p\s��������`܍�p".���������s����J�� P0��cR� ��mlڬ��������P��P`��Cgr�/�����v����X�8ͣ�+&�R%.휘�*ނ��B|St�^N{<�v�x� �򩇰�����w���K���(`����{�-bRyCX�qc��
T��I�ք1s�l��k� �U�9\� �q�R�� ;*c>G`6@�?��1#ܳ��䌧�VS�/��t5�"���c˿+����$S�a���?b�etf��_�i�]ióE{������	p�k�
*������(�>B,yn�q��?��e�V?�I+��h_��Tb������Wx��$���I�-�X)'8�@qΥt#�%xщ-�O�b,��>_�b3�rpxZ��VKx�B�_}p��U�3��&���|���C��o_�*�v�6�ւ�V�����檓ا�[��݈�ݾ���ٵ��B�_-ZU�׺Jh�:��? ���ǖQNz�?5��=>#�Kp")z']�F>A��cC�G��0#N6�/�P�����ji!�f�petq��� Jˤ��j ��+A%.�Jy��J�%�ֲ�O��%�7���,-#ɏ5�o�s��#�u=yz)۽Z��-i��w1���eP��<�C}�6��I:�`F��X�x�Mt�r�����m?35$q8o��&�����=������`��ź�"A۰,P\�Rn��"�\��7�\I�Ҭ�����꫈�M�5 �{(���e�{�}��&W�Z2���α|��
�GG"5�����-�!E'k>%�>$����Ϫ�rM��ߐ=S �:��3$2�H���L��^���
^T~Z���� ��-���Ǵ�ϓa��-5R��`ѭ��pw�z��M�K����ۤ�[���帋���{����A����Ig��n��cn��j��响8����r!��Ɔ�A�c>E���>86|<Pv񎍮|�
�����=ҁe�s��v5������"m0�b��2�u���9�q���5/T�a���h��,#D��伱7(����>H��q(\�x.5�d�����+f4(UT*^��`�9�4*iT� PM~�;�bb+���#���4���_��0��,�f/P��Dty�}&�_��%?B���̚�k���UU9�MR�-߬�zV%hz��j�`���Jg �a�F���t��o��n����}��Z�T�
�
�X��J�39}���F*J[�����ig�����<��5�����вaΌU��E���+����
�Z��ڽ>�U�������S��lR_���[���L߀��Fs��[��T ��eb�
���^\����m���KF�$c�����W�����d��Ί� K�S��������&Nr��3�rٲ���8Y�5�i(x���H5���`���65H"l�d�<½�
%��K�Ӊ���dc���c7���$ˆ��<��dC~ڥd4�ǓP��m~y�2�89���9^{�k�z���Q(�/d�*���Qk��E�}՛ָ��j�5�O�ۏ�0v���F]�w>|LG�R������aUQz�CAШ7O5>>,��`{�'�
Z��?�c5��ֶm8'�q�1-�˼>�JA�4Sd��Z��_F'���!� ���Z���������@��LȺ|�����yA��Ҽ��鶉�k6�K�m�S�h�ُ̲��\�&���pa�J�2��Ǌ ��U�:��!ɘI������3��LƷS4�^��0g&K|�*Rv��x2ZGW���,`�B�b��;�*��M�q>9|D�D��@T��R�$q��E�i�s*��~px�@�L�%1�Z�a9������	��2�<��kܯ9�m��<VF�u'N�-�$�n����(7������}t��?�+���vK�?�$�v-T�-^�, ��os�@Z*�&�T|�wt�[�_��cq��|���
d��]r=�������ڜ�x#o�6A��!	��Xm�N.qI��ȏr���O��a����BT����*r<�:d����,z��!�WY�B�Ɓ���)�� �3�c���Nƨ�m�
t��w��K
� To���>��;�k	�M��U|�Į�]�ׯ�[�6e|���!��7 ;̜"A�/�������ﲞ��O�OE����޶^b�Nܡ�6; 2����86����{�0hHf�z�Z;xg��7�]���~L�,W�� c(�b^�,�(�&`��B�
���X�h�k̀*0�|�W���G������U���`��գ��DZ3q�<���6�q0�r$��Q>u���5W�4�3Dz����w���!����݂dP3p�GGa&o�����ES��D���.T������$*��n4./etP�ha�N���u����c�C^��*ɫ!i�]�'�}�^�ͧ֕ %�W����~�)۲I	����Ȧ����4poh�Z���4R����E@�/��#����<6�|��3��#���G\�+A�:�5��|b�ii
�L��쨍!'#�X��r�������GLr�� cͪʼ>�c����՝����Z���'� N����sra*�V�cA����]VmZ�|XZVf��(r�(��2��"�`�Ӻ��U�	���(�y��V�RA�l[=�J������� 
TFĎVK�~?6��ʨ���I5L��v&o�Zf��0n	�a͊vO՘��mA�����N�m���s�ٛ]-Ԗxi�s��L��E'�!
��>�z �*OI$��s���VtZ$oG�9wK� l���&�ʡ�1Št�ϔ�'�ůjC��AF�%��9����b]ށC�Q����4@M���C�f�ؑr����g8�Ĩ�]H��ɆQ������(қ�L����Zɛ�1K"!L����|�J��I�誨�z���ѣ�м��me��XcE}���~��l=�#�<�k