��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����}����ٛ�!"!�:zxs��2@��=@Їe4�e>�B�����NM���!�զ���ӊ����{!??1%�yO��q��������<��H��,��fC�38�KWN��vM	���٫O���ܼ4���2­���W�0 �yr�*n�rz������̌�,�:��Uf+6�1��*b���[O�o	
N��̴� M\1-�"���{�V^w�����X|T0�q���*\C{��;�%[�jRR"ax`(����&�o�oUSϴ�r���)��1ȘXGi�~'N�R��rSRѲJ� �X³
�<L
c��O% ֮�Zs�f
�O�@
^*��� �	��DyE�	��ME@� �>��җ�wQT��dI�P�Aq�Z�Q�֫/��_'}���B�4B~�z�'����	r���� PE�d�vM߫��WN3T��]LNЅKQ��ێ[����0Qs~�K4�͎�A��E+�o<`�_��o齜��F; UQ�$�6Y��$w��v�Ԁ
���dӗ�>J������������g�Z���AƟ�β�ܵ��7�|Ʒ��:r�����Բ�B�'��w�y��q_0
�4���g����0|���銝ݺ�d��-�sS"e@@�a�Qdç}�!���@� �?)�z�+��D�)׆`�0EWH!L=���q7�)���܊p!��U_�`�]�̭�"u���'��L^��' D�tTC���R��#lx��EC2r�\����.�"$ ��ᱍ�!�����x�;\D���$L%���ڝM�ϝ��S�N��41�&cLE#�[�矚����u
/ߘ
�)�F���ν=���;����a�,�<�R~V�n�ey�Y%����T����(�s�g�T�&��c7����	�-�;<������8J�\4����?� ���ԟp!�����]�5�ۈ��+K���U9��A�����t!�\����\�Vz�V��\�k9�Qc.yk,�y�[���V,��>R�x��v�RK�D4H
���A]ht��,e�Sr��+�]���'���`L�(�jZ4S\�*�c�rJ�С�z�64�-m��K&��%+� �H_OhU����"���~1O5��j"6��؂�(��į�?Qo�C��� #\��c��_$@�]�[d�P��Y04���Z�L�Wh�;����h������H� ���E�I�'tLpv��.��%@�{��T&lqo�8��W��`3!f�Yn��V��o���p-,˭^w#J���D�3-֥L�t��O�UL�Bm0���>�?���/�z�s�lT1D��#�b�^�V��lW��@ε[�_8��FT�vd]xb�_�"4mB��`���b`f�d�l8�d0�RVG�9I�qx�r���S�`4*Y�3V?�L�׾�3h=����0���̪���?�������ޕX%�oŬ�h�_�UqG-E�������h��%,q��vz�Lr1\Ʃ��GECL��c�O��E�j]��8Ӛ��(Ʈq
1vi0�fn��l�݅��D`+9RNTR��W���'�s �����-C'U]�BF�v��v����S��j�5�n8����1@�U���l�^a\��� ��0��S\ԝ��;,�l�9�^�Q�\v6ь�p��_���j�]M��K$|9��M]�/ªT�D�%���;�� G9�����n.�����+�^�ܐ�"8��!�yܦ�[>�h��C�rR^�^$vo��_��Q��D��ǈ�g�k�z�]%�Gɧ0��y��/p?*����>�A��]�=Ʈ_�d��g����[�Q���
Z0��ʳ}����E�7��h+Ǘ��1j>��@w��Գ_ݢ���;�����u�z���1���7��Sۢw�Gf�6�W�J�̩&�4)a%��:�>�(}�0��mk�ή�aӫBՉ�ńXm{:�FZъ�Pp�TPS��pTm|mz��Oi���.󙽵F�iN�_���H���a��0b�ލ#�J��ͲJ�	rI��%ۅlrI4�y�C����C /�N��.p�$]I�Ƹ$/�ibA�"�%T���B�i��ݮɜ)���ZH�m` ��D,�Ra��b#$��8,j��]�/{V:]���!����7t�̒r����`���zmI�:-�FH�jh����9:�0���7��>1�2 �<�	k�R*U\4M��YF�����K������5���ms�jԴ�>����5aޘ��C[)��N�]M�}В���(�(��{&�i���j����@��E�p�SeLp���8S�]�s�Cف35�`?]�_ؘ�! �EUf�F�7>�^f�Gย������� ����%���������'@������Pj ��ڿf������z{\h5�����@�ƭ�瘻ˉ8�$w���FAn 0vd!Y�=3��O��^�{���J:���T�f��t�GN獏�p"�r�毺(�t� g�HЏ�;��o��L>�M�S3���T�n7s��Ʀߏ�ңajm��������$֯��s�٦� ��@��'����Ӧ/��F�õ��g�?�y���h�����_X�}.�WȂ#y����)��xs]����:OQ4�!=���$����V���/�ꎰ�Y	�ɻ��#X#Yk�{'�@���=b�NUC��q�Թ�>)�󏃈IJPi�� #1�����N�%�F�K�����m=�w�>e�iH�/���"T���RR󤧥�[5���e��e��.1��A��؄���n�Cq�Z��q�X{M#�
^	n)P���Ɨ�3w�95<��L�r���d�?�]H�Zo�+�b���q�#Ƿ�8��B/k2%#�'�`��Ϊ6{[��)�|��Gq_���P��{��J�����Q��ޮ������ )�<�V�р!T-�0�8�p��V:y���gykƶ-@���oV?��Jb��*�"F�]s �3*ۮ�Zd#)�> g�������lYJ�~������Z�6&Ú�ԼSy���A(P�XЈ��6���ɜ�G9&.1�����kq�I�6��F��k��6v#��Gpq9�✳Ҵ^���\�//�r�6F��fHU��e<�f�v6}��� 5'h����:a�ε���%�=w������}��<����t�Og�X�z�6���F~櫕0z('��C D���(�
�]R�h{<�t�&�(ͮ:��u���� )swPu4��0�庍#��Y5�P+��F1ss��E@xi�D�z�)�w�C@�.����=`�bX�ǥ?'#Ѵ������'�Wn�f�no8��xS£w��x�+��W{Z���5��u�����:ߖV.�$���$)Qƚ���e��'X�s�{ǅ�]:���|F,��rKQ�;�� Y ��J����wDdCb��6�g,��K�l��=�ro�h�_��<8n��G�7�Y���X:�۷��xY����pui��3��ߓ4�W�
�""H�L{X�/P'�+.��@p��ghY��[�	��^
7/��$Ӝ�51`��l�j�+H��u�C�5�"�]^�45[_���r��67R��(C���q>fE ���MDMe�`�����f���ϝ��Y�������k��@Q��)�U$��p3ح��_�r7�[����s]	��SYԢ�������n8b�v�ՙԺ ��$:0\b���:8�F�tD�M�8��[M 6 �z%|�X��dlOvA������̎�ib(sJ��LLw�(�Π�o 'Ȥ���%[20��E$ ;t�T�\Q��A����kv�?��VM�ax�SU�ۤ��ͨ��]5�:�m6ӭ�_�֖.����C{�L����#MᎭ�"��/`��L�l�8y&���{iUS~hX������g��3M�p�Ȁ�����@z9��ڂ�.<ջN���-,H��܃��F��Bq&fS}R���^;[~��%�)lW5����5
=��3u�ż}��$k��S8q�Oϸ�@T�k�:�K�a�Y`+H<R�{���`���N�3����V޽qg a{�<���^�)�q��	�@y�ҁ*�!Ѝ��EM=�Z�osD��Qv��vZ
b3q8�S�� �CO5�z�߇���t�ǳ�>3U��;�l=sVx
-z����˰���hɧ��6���{I��Q��g��b�$w+�jø%�6��EW�(��#;*��Xu�!V��xI�G�죩-_O&�>���3�B�[,w�?�G�ͅ��v��>|�pp(��̆�S��T<�N/�]�����H%�k�1kj64����g�~x�,�f�@����b-����\~?���d�Y4��m�������@H� �}l���ű�i���9a/�B�]-��݁-��H��\V˼Fϊ�af�y@�oD�� �F�[,�#�R�2Bz+W�zb��8�'h�-� �e���8�k]&�Փz�j�2u�����DI0����6�;�咀��jj~��ɽ2J���v�w�n�Gǜ�JZ�t�B��)�{�Y%���aYI�O�y�yi�IZ�2uM�,��8���;7F�~U�7�$�$�ű�S�Nڕ��%j����ܝt-2�+��!0Ԝ�W7�t��t�2��ved���(sl)�T��+�t��Q$mb��H�\�V�㵥 �2��=Y���wO�`�%��&(�z�v�s�|��k���F�P����Ǻ�:�T8%@�v48����Q4�{1P�0���4j���6�>`1�V�dbꪢ��DL⇗�Es�W&Z��_�HZp��N%�����\�j�cZ�(�V����Ox\�"u��$0�.�*����
�9)��u�b��.�hj��P��AKC2��9����-B�Q��]	���ធ�(�QtMV2��*F��5�N�An�2xL(��t���=q���Qk��Ş<�1t����;��.��C�"�85�}��;���"�+�J��@��	�����#����������b]ߙ}FwM~�"�ď<$\3����	.d�#&�.(����t�0�sk-Y6W���þNt�d���/=�+���ESt���F�����+_0����D��MwC@k`#Aqi���cڰ6V