��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm����질�95J{۠�0&LnS�3�s�ǖ)�*�X6F_kS��J�O�[�˥�Xt����mS��pO�{��J aI̸l=T�E�����J��DW�Y�ǻs�g=�9��tAk&`�4�3E0""2b�M��y��eò7K�&����G4��8n
3�ɕ���Z�J�"�ǹ ��;3?�Y�b��I
ZJz�i�,��`�1���(��� J��U�Λ�(�7"���饞��PӞQ�ah4�ܼp��hPf<���v�����������:[����h�4��:y��UZV1p��*�1��^p����
a�y�uz� �l�n�R������9S��|��i�(.�vx?<1*)�(�_��7��ض�NN����iuV˖*�[��H��Y-׸�{ؙ��ej��[�_����]V:��d��!��(��7K����f�1����;�ن�n䯦��y�7����f_�yO�=k o�1_�_l�^�Ι�WW�<9���Q���Z�c�Ʋ�>�t:Ã�8�Gو9�W��
���J �jJN��}Sk���d��|ǁ� ��Pΐ��FU�3P�h�򆤒�����S�%0���c�O����n� B�1�|�@��;T�7�P��������;�_j�m�&\B�ꪰK��ql��RKѯ�j܆����xv�B�7��6�Z�F���`Q������@[��q��A�����Ak���=&���!	C�Jщ��O߇���]�p����x9)�|�Կ�z���%bD�\4t|�j$lƾ�+�;'+fs�d���P��M;���A�%l{�?	lDB�����В�mC�܊>�$)����
�sjM�1r��$#��z�Z����B�l�|q����k�Q-�_Q��w:��n� ������zB��������fo�z�W�QҞ�.�¬H��R���Lِ�_�47��{�֩��=�ʔ�
�#5�N%��Y;�a���5z[+�Hy��Ѡ�z�S�N��C��h��κ�|2�g����K���-����
ie�~	4��1&��P��X|1��(J���U���f��P���g�I��2Ѣ,�"W��G'�9���ٴ���c������5�	�`l�l���%jn\ؼj���0���Iu�Y��a�qW��o����:E{��.;�ɮ�]��ݬ�F��9���ؙ��O�=��?��-�̃���'�Â�S3���7N���M.�!���#�����V�zfR�D+e�GN{f�f�
�}�l7'��v��|I.��oI����,�>Y���,���aX��B�/�T+)*h�)P��Zƌ�p\;uܜ�ը�X]�}i�W���|kēu�r���nD��\-�(m��, �%�a���W{��+�Ew�ry���siZ2h�|�k%J���9Ѫ��Fܗ�įgZ�*Q��.��Dv��  ��/Y��L+�Q�$1�Z�T��Ⰼ��@�$��"���x[t��yJ�dՆ�Y��Cy�����d:6ae��ĭg/@_'	���n�-����}U,`<�z�u������M�_�=ʐ���+f��5��n��i�Nr��~M�erbgΛ�e����
�|˯	�8J�9��(`L���ʕ��;�Χ<H��Uc��ٿ��Oh�-�2�لFXY'��&��1�^�^:��żBC�Fm	Rw:�����ݚ������N2�6Qo���!3p����� �X#{ڠ�.P��Qx2�.���������%Ϟ���u盒]����|�[�ɨMT���<>���t��-)�;�%����S�T��"������DZ�zF�!��5�o�x[�NK��1�����{�F�uT2��Ψ-���fF�>l��x���z�Nٰ!�?�b*���, !�mA-�3F[�Z�c�\y(˧�,��]��,�jN�����]�a�)��+h�O	�9���{F
�'w�~��1�i� |�����bW����[�]BE���D9�"��j���+ژ߅[��$��W��~��Î����-��Bi8�0�!��(p�2�a�bpk����-UE.�P��� �b8'X��$��Q<a����Ӳj:�d
�����#�x�g��'t��0��P��b�����9;�hr�b��B�u���ʶ Ii��7����!em�;:�:*:AuD��;/����}��e�ٽ᾽����T!'$�}��^��a�|3�;�P"�ru�WV��!��� x5d��*�񂇧�p�m�Y���*nhTA�]�����Jc@��.�>8	���Qc���dB.����2)���x�>Qꔯ%FHh���ԅO��\Y��]~������{l�]�y�vis_��2��M*�xc�z�l�~7���Yldg ��m�a?[T�� ��aߏ�yə�-6
Ұ��(1Į�U�u7(x���5xr;�#�I���PɃ˼��_�UE��4ǔm��{(0S�_<8�?���iq!D�:��eaaT��2���j̚�]j/K���Z���xC_�&(��x��Q���@[̃��>x��yb	n5LY�- #@Xʒ.Ѱ<o�G�_J�?�X˨��$3���R��rVt��73|��(`D~�m�BI&��n^ �����W�3x��I��x�f�iA
�5�({y}�--�.U����F�]_u��^=b�U�J6s2��WH� x�����ѱ��Sh����.JMl�����s!�KM�?�o�毡�	p#�.�]b�C+�;�>A^T��j� ��1 H�֩��[�X����JP�]Kjc�Й���v،w�卤m��� ���μ:�R �� ��qS�~!���E�-�"^g��I]�F�a�y�3�/ ���"�k�|�`�<</+U��j�W�I�b�8�,ϣ00b<����"��U������KW�c�)��B�Iu�JH�fS^�b{!6�W�jGx�5S���n!DɫE��ӎ&mU��&��(��qV����\M�뾈���c^�e�o�!��O��7�Ca(gn�����
�Yw��m��w��݂}C�_��ϱ�|V�t\6��)��@�;�J�P��	dH�3���.�L����tIE��5��"�[A����G�J�U�!&>���u�R�6�E,' ����W��#T���qBi{%������j3��?Q&U�"�!�g.�ck-�A���l�ʿ�����6?֟ma5c��������_�A�k?Q�㇠c���7�E�u�f4�B!(��Up	?����ŇGh�ԊL?Ɵ���o����)n�ZUw�6����x��4��Ҏ�v]s�Uu�XU���E�J]{�mˠ*<���0�Zk�d]A��m��M|�*$�y6Xg�x����̊�G��3�A
��P�Ңi�هt�y��$)�BN}[���H�\���8n7��`s�kiVI�֧C�#�'k�K���r)}KqAe�9�Q��҅L��/K���'���%`w�s�N�BL%����n��/��̋s�M?a�5p~��I��d�������?X�G ݰ��E��%�(��M]S�a��ze�H$z�
�	<�n�V�Ko�r':�`�ѳZ"zz$�*tJ6Fpf�y�]�з�%�0@����W HVY,�+�l���2Qvr���?Y�bYm�q��쐖�C��t�Â��빞����47������C_��J�y�5�jޅ��C�\��4���a�TC̸���$��e��qW���!�[n�̋1��U4�)o���
1�Fx���q�-F
��e��
ݜ94��mj[�����F��W��O(�k�f��&�_\T��\�\��R>�������u%�Y%��ؚ��ҘT`5Y$��W,�Jjm�fh�'�$�	t{�}�;f������;���*˚��죌J��rh(�A�*W3����^�ttK��+A+���`�[$�S��	��o�U�L#�Wn�h��S��k	Ag�d��J�"���vl}��ІJ�����biB�=��E��^�~� ��}�ymœ�)�ik'�̮%�O�(%� �@�2�̀�p78F&ݥ�{ �HE��Y�ݢʹ�h�i����#��^1�	��!����h���f:*y���Z�S2��p�F'O���R8����u��
��Y%2�j�\�uhӯ�&٨�D�P��5�[��1��x���֒H��K�I�]	���U�d�;��y*5F�7��CT�H)S혝y�]�ES[��f�(�}O	�G����C���+�NF.H�)�~W�Ղ͢0�RMT��:�H�r�p�@�kɻ��Z%tQ'���D��l	mx��3�}�^�X�kM�v��W~\P���7�1*.�df�!b��*�y!�@"��������"�$�_���静g|��/fـ5�׆�;�b��
|+R���\0�\4 4m�0��vr�x�*@���_�J��v�*&�)Ă��._��j���T2Z��A�R*���O�������v��wՙ�7.q�m�dc���t��
sӘ�1���c�8[����}[/�Q��(WITH�Oр*�i�f�yi�"�H{�o�O"B���Uki^�^HC}����_<%�_�@�"̆&�B��SkFD�Z5X��)pvF$��jB�����wS�	1�*I�>T2�[�l���{�	:f��-5f��*�$͠!֋X��k>0znJ��J�F��.��V������ل�B���3��ArTj��������Y{y�ǫ��A��B;�[(�.�T:FӻZ\4�������AT��W�燏;��s�
��5�?�)�!�}Ig,��y�