��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{�I1�+��:�M�cg�D�
o�2�/)O�3�UP��q��9�
�8:�Q��s�Aϓ�
����>�֎Ҙa�h�F�[Ѽ�b��{�IL�M���BL�h"�z3;�ȅčuJ �H�Gu<�5阃G��7�r�Hal��ݥ��)����I����°-�8_����Ֆ�`j�x�׶��q8f��W�L�A,ۣ��_p�&E��m�]l����5�o
.����n�'�Ȓ[�	�SB�q�rk�7e���5���R��pA�|��D?;T#�!�Z�r��)�[n�*�P�O�� "��M�Vam@��G��.Cn��pW��&B�n���Y\���)$�Z#}����NU6�MC��;t�t���J��Ln��l�Ž�4QSt>`"-���﹚+�L�[.3e��I�e�f�����p���]�����D<�"���A��NZR�wԙ�O�R6�=�����n���B	�����H��h�1�oJYr�˪�A���߾� �X�cL��j:����V�[�2��X���>(���:D��模'Asl����Q���#��u�e9�4pZ'�������K��m����b~��R��'���E�)�G�c�+��-��E�s���,Q��Q
V<��<ه���!����lY�$�	�@nu��$�	��7�g�g}!̷W�F��
(��y8`����o�}��'�Fv���b�7Y(����N0
+)h.x�/f����w&\�)�+����3�`X�bJ'X^2���\�`R����\Gw�
��<���5���0�����6�ɀ�r2{@�SNUƇ���w����w̺�SG�Y=y���]�� ʼǏ�����ZlyK�:w���@���pI�������$�
���_������,��.2��rrTHz^Z�f,��,�ӡ�w��懋�4�������us��T�'�YFF
t-d���I���+[/w���-�����r_z(*H��b#`��-����'�J�t�����(��i �֖SYڮ�"���`b�6`^C$i濃�
I߶�v���	�M� ��IQ�o2:�W���x?�9�F�'�����@����[ӡ��3��nh��*/��w�n!>�X�B�*����p�L����Dx:k�?6$���߷ 7���jF~�갫��h���إ�^�սRֱhy�^9�Z �/� o/��0����^FC.,��
nR�S�an�)O�Z�p��q(N��̓B�c!�B�ثFG����&3 L�P����v��m��@��_9Ub{�FԠ�&�Q�%�nhs����rn�&����b.�+O&{t�h�&��
�"@G�>�g�i��wĸ��݆���T�����ԭM�)Ί ��՟VF�o6�-R؟�Ϙx#�X�>~�<��u-^��'U�x��r[�4�K�k�7��`�WQ�3�l,E�����,����^�X[;.N����3������4��G��q�ю������;��6������E�XT��uN�����0�̹@X��ƾ����BB�Ss��|�!��ƨ�!�ЊX>����!�Z���-:��z';��`s�n�tX�,����4�T��(�#�l;̶��3,Ȍ�j�˥A77�$E�Q�<�}l8��ws��>���ٸ�b�5?�n���"^o��<��/�q^�k��Zd��3�eo{��|R�Զ���j-�'��k��Z��!R'�Fz��y1h��r��5tD�'y����9%񌗁\�A���i�_�LD� Â���J
��\�k���-���9���%(6�j�rO�Y8�+�[��W�s��h�?�I��R��#�:ӟ[��Hnnh'(�g�Ѷc N�~�|����r��<��7����%S�F<����.�w��RߏR_M�oCW�������u�X�f��3<3��=��F��]~M�9�Bi����zJ���IC��K54��wJ���ѩs�`r=�+���A��X����&�H;CY��ZCS�3�2s�B}jP��[D�P���oُ,�d֭|��R�u>n�=��1�f9/�b��僰jH�R������f%ͭ�m;�
�v�)���2=Dv�??ҷ
J��M#4
9�l$&����@H���Si���v޲��}�*N@�:�#[���ƌ"M�vsF�t�	�Rz%�ϵ��L�\�Ⱥ#\a����!���:Y���7�S�mȕN�GlzP���w_��i�9�q־a2�$k�DC�\��$���Z�J�~�!�.����zB�t�SI9��q2�F8�4;/p����K��#n�ȩP�o�Jx��W�&���)����Y�`X��&��~=}]�}$����`̨yد�X0��+�YQ~,n�K�5�+m!�\�5�|��)`�>����v}�?Et���˽�w�W�^^�w��} ~��n���E��5<z��)��Zt���ͩ+��o��� ���:���R���*��{�� ���uD�O�
�.�g��'��=�F�I�$���Q���3W���A4�$���.>����e�x~'P"p�>-�"�u]r��n�xn�5���eYҕH�R\3�蠾VDþt���ɣư��9fa�ǈe���>���w����0���$�0<6Ɛ`�e@9tA�K#�{�ڧ,�$�Q�V�,���67xݐqn�7�{�ʚ]���j���V��W�I$��ݤI(P<���y��f���]G���m3�0��NO��[M��9�����#����Z����?��W� ��C�]/�/0L���<[�����	:�S��j���ePGYC��F�7��tG\kS�z�����>���3�N�0�'�?���gՊP�TaS��M���(�4p������@J^Tx��иV��Nm�xC,�v�ܶGA�b�)Q�j���T
���(CK��O�wOY<0��dHB��M`��Zdm��Rl�Ŗ�mf��ay����Xij��|�L}!*�,�e�'B��pAt� �8��q}}8�W�V7���̆�e[�#d�bJ��U�D��XD�l�U��zLžu�7	\i�Y���~�&�ƍ�:����gm�/��_��Y��Z4E/��Fz�X��Y�OaL4�[$1��E9�86����A�d8�� lY��������6�ٗ�����,Y`%f�2���h���y
a���S:p�Ld[@[#rL2 ���K�<�Y�Cw�]���_��rv���k`?*4�k#�u�8M��)�b�dt^� bTp��g=��;�0͍x�}���:��e�k�g�ǋ������2��6q"�3�e�lX"�3C�*�,q��?��_2����i(�������I���	�뻗�P���af	. lX��HݍF��1
}Y�7ag�G���b���C���2^{���������3�W�l��ߥ?k�����R�9P^��1&-��B���.3����o��u�?�����a��u���K�a�]��(���T�]��<�Ւ�?���l( �(���1J7�|bx8�2qoسRV~/�0��FN���(6H��(|@���7�:ƅaiX�3py'��B���&�3��CX��B�WjT̓Dr��ani@hT�.6�!�}���i�L��١QF���ޑw<��!���$��$��l\�Ƿ*�*1*��*|&�k�o4�Tup�n���C���o4���ǝ�$J�4���גX[V�T>�9�{ѳg� �l���f8��+���zY���CA�޶�y�NLqab��7/dў`O��N��7��D}��A<��1N��K�d��|��Mg�&�.��a?*�^�������8������c����o��'��������1z���)pa��7�,
�ٷM
! ��������USP����#�R-���&�k���Vs%k���[2^L��䍈۵�[ce��R�`\J���=}`��/4��Z�!�T@�!8�%���w׳�^�;��Er	�{ě#"?���Mau�%�A�����T��.� �̅@{?GP>���}5
Oӆ�F�;v8 4��E�!x�E��@���q�Q �iG�r�T��ڗ�`�	�5ex&�a����,�koS<|Zf�!F�/��A�R �վX)s H�������9=����Hy����^���bA�0��D�\/�����7�H,.iG�H����>-j �)�/�+����y5n]L���#lW�T��akֈB9��vt����B="����~h�uF�=3�ܐ�LZ+|{���Q��]Y�� n	��1�����z���D�r9�Ǒ~
�p��3�����z!���;	)����,��J��T�8i�٦֤���b�����)%ֲ��;���~(=���,��j��Zr����B�]_zF_܄SN���'<�X	� m�I��a.	� �sE�7j��A,���	ߐ�1ٺ���.���"��e���q��/}�v8׀�Fq�%�_W�@*�ak�}u��7�(V��|�NX��Y��W,�p�¿Z��ʵ�Ŀ�T'l�-@�m��9�2ZKke��4c,a�̧���L��~ف>��|��J5�#�1�o���6H-w������]�Ǡ3W�ϼ���8�UԔtO�"�'{G�-���3i��/?|:�WsOR�
&�@�t%,;��y�x	�3K�A}��a,E����}��:�q���vϹk�R��Ͷ�팻��XI�5ca�r<_���q��ғ�}�B�I@���:$�ݨ�]���r���`�OQ6Pj��H�\�&�yx6�}����)� o>�"�Y��q�Xs6�1�L�=����t�S�[�
Z�H*P����y�WV� *�?E�=jNm��(�O% c��T%�up��^Pc5�����S}2Ca���&��b~��ۃ��}Ku*�,̈́h8�����|��t���������Lv�EM.�70�x�q1=!ɍss��gt͟������^}�U�j��;��+ ��JÂ
�)K�Q��Z���R���C�Q�S��8�&1LW�땰9��R9�X�V:�ir=�T�)������z�vm�)>�;��9�'����TP�M�lGOū�f���c�ʧ�(�\�o�"����ɔCI�R���c�+>�� ������t�aQs��"�rtV%M��>Vc5"v|ǜ�D�x;�v��ׇ���ϖ8�n�N��j����[6��Z��M����㦃Cis,�>�'��{���:y ��m����������u�9r%���Q�p�1HW��Ai@uK�#�S)�,_dh��I�iH��U��:�Z����Z}���<�1�)�É��I
�1�|"�^u�I����hc��d���[���5[)Qaf�-���x��_Vx�겣lR�SVt0&�e�"x��H7�xq�Y�\m�iԗm��W��D��fC	Gw����:���^���qK����`���W
�o\�H��[6�<7�-���ܜ�O�}�r%4!��?UT;���ҢU�_*�r7@0���&��G�k�܊	�[&�T6�r�2�t1}��P�^?B�Fy��")es�q��Jk�MDy�qQ)����!-�M�AJ�=F9.g�d-��L�:1�RS�՛[ۢ�Ұ�e<�fe��W^@N�r�����a+��m���c!{)�g���|�����)�a(�8.�5��
vr04����T��n���`�����O�Ew�E��WiӞ��b:4���,陮-o��1D�k~*��,<zvP(��VXj'M ��Wa�
hh�B����;���C��a)�{�B��Ā�=�T�SU,��?�1���.T����̬�=Q�ś}�_;�ݙ�T[��gً5ڪ�	7�N�;	�T�ו�8���NI�P�(2�d�6c���,�qpO�ρ����R�j�����,5���e�W��5d�_�rz��ml��`z�H�ɍ��yL�S�)Q�yNM��UX�2r�]T��锱�����"�P3
.���P��!+M��kG��D�d�r�%�t�v�T����m��[�vI&�K��F7
wyƆ�wcb���Q��́�Ϛ���Դ1+^��/iL�d�YiġZ%��[^�ے1�͋�^�u�aBݒ�zb'�>/��-w�S�E0�dPc�	���b��֑� ���b,Ki���o�*<��D��{��>���^�������]p��N�̋&�� ^#����~�Ao�Z����WH-���&O�4^��o=�yM8@�3!z<Lh">���� �xF���&�"���2��V	�r��9nG��ϕ� ʕ��:�E���>Fi���$�������6V�c|�(�r���xY�U��47�������0��|��3j�g7o]��%�n� �3��m�cH
q�1��w�t��I�y��Md���9M��ޚ-C%�UM5%�� ���g��)��[�_:��kq�
�������Ǧ�|05���-d���K�Aɤ���e�s��e��' n��s�����CE��l+����fIǽ���)"	6��2�~`�/��W�~
s-��͕lv�F�>�Qy�ZeK���k������M}9Y���TvB;Z_3�v�2�ϯl�I����s�V�}~0�,ς��Z�Ǵ�ہ����K���E��?��m<c$��c�
�Qc�T�pĊ�8�:����R3=�M������ ]%i�����7����嵬�=�݇T�0N�=?�]Ss�K*Cm	���b��+�JPғn��3#���T�=s�T%��az;n��͏��S��jiBtfT����b� �����3��<��-l28$�>#�ՍR$q���Θר�t �&>C�[��v�H���vs5iRW��vU��9H���!�8�S�~��3�v��B��'�m�n��]b:�L�9&Vaʦ�� D����R�����T�o���8��&��JG�vaJA&6�����6�>�n.|�H�Љ�KYQ�X��P�Ji5^2K�ɺ���\;ym�"o�4h��Hc�����\�lKC|�R�O���5�[Q���c�D�Ӈt��ԚD�(�Z�р��q���/67�@9��H�aݫ�E&�O��h�ji&Eb{F?a?�������<�ɹ����#U�f=�9P��g��˚���s�=[�B�)����[���yxW���Mv��.\\���A*�iq�W�SQF@^��cG^���:$�δ/��a!!�K\�"v��%�L�B+)(����#�m<�����a����&9��n�cC�T����峘��a_J�4�y���� ;�<�8�b��ZB�`c1t&M����`Ue�_�
∕��\�قc�X�.snZ\����5Cz���;�����cƗ�\z���K(�X�Ŋ��!����<���+�X����pQ��,�X�E�\ݖ�%6W�$��T�d6Mg|�^J.=Di��������w�<���g|�a؉O���/�ʫ��c�ބ���B\��xx��}�����7ǕYF���C�
���fRW�����$1t�=�h��矸xÇ9�u�ߏ�*���~R��y�2q�S?�x|�J�r~�k����"�jW���%��[���W]�oעO�����TU���H�%�=��FG�'�F��B�`����g
A��N������u{����@�F�؈��G���T����tZh������1���	I�L&S9�E�sM��i�PZ�!�X,�Ks�NO�j�?/nB!�W(n��l�Y0	y���-��M��hM���;���`��BI1MD�	����C�A�ι�D]�E
(���b޴��*�H�j�����v���XZQ�"�k��[�ZTQF���	��L<E�p�i5$M;=�����n����"cI$%��,"��~V���^�B)ᣌh�����z"5[��R�ȅ��-J�oP�����Oh�	�AuG>raC�Ȇb^����d
�H��	���h����<SP�=d����"56E�"<���lë��e�ս�}o�4y1�.��
���t��G���n&�G�.�R�*��%8����P˧�߹�7]�ِ]#��q^���ɨq�\.�j&x���ghr`��P;�����ng�uy�~߳)��y�)�e�0��4|g���f�j�CW�?T�fc�GD�&0��ѧ���UzY/�+�6!�1��'a\��>R��%tdJ�Q>K�f9Mf���is8�K1>���.�E>v�hA\�ټ�fx�=&|��/wQX�o�e<X���ݚͲ¹�p���(��d�Q�@zg�
�p��L�-T��=�9��ݶ�q�o"����z���?�
�?�d��x�=!'j����9��e���Y&�S�Yx}������o(8@��H�/Xn�[,�u�+�i�Wr&v���MM���M�%��u�a!��?'�/��������Е%��(H�����I{3Q�k't"�5z��,�m��s����	��bt�H&V���?,5��d�8E�V�쳐��¶=1���!c���%k����i'Y
u� 9.�'2	h-V�}��a��7`��j�EX,BB�2t[�����y�����6Ԙ?��e:p�R�	��+,_����ꉻ�5���)�C��.����8���\Q�<'�[$�B��~�t#fp��O�������q8����!l���Qf�A��m?+T��R����h�pCx��$��wjf=��cZ�c|�+����h���(�i������LD1Mԭ{ dp�X�l�����oj�� a_~�O�172�(y�6���4�Z�� ^e{M
Eee⇑��ɵۼ��ӫ=�G���N����!M+P�ŕg]
�N-�{����He�o���ο��a���:j1K���7R-��jޖx�n��4�)�er�=��~|�<�mN��Ν�g^�K��~���q2�y�/&|��{c�~�a�!o)��Ґom�f�CS���oBıt���s�\����p����ի2m���v���}�􁳉.`�c��*s��T����*!�b�����(!�v�T�Bz��~��5��Ҭ7~���ײ�
8;��~�0��C������-;?�7I��T��}���3$��MS��� y�cc(��|�eA٬-0o�T�������i��� \��9��j �G�n�ʶgq̏����TH��]�Mz���i]��RmM(��Ӛ�Ii�o'�����5����4������C$O+��
w��>�����'��5�m�U9���Y(��ob��Y/!=D��b�[�̳!B��9�C�~ڇmw���>��5�����1�
�[;9��o�Cb�e�c��A��e(�X��VVuJ�2Rֳ���`��j�M�Ț���_�	vxQz+����y
0�gW�k�f$b
�[��+��h٠k�����t����z;�fkl�~d�m%����<nڢ���?���]��^R��/�:��p|67Y\�;�;ٔ!�M¡�D��ǫ�<#e��y�&�@���]=cb���|��T[&t��;�FgY7!����s0����1�=SĂ,Ay����G���O��_P���JTv���]���[��y�K����S Ut駟�l�s>G�e5�0�e��2Փ�9e�»E�_:��M���
�l֍��n�X�[�v��P�jqx!M�]�z�8�k��*�E���1:nPV� ��c"j=I��O��c=yЦ�^|��W����^a�����},뾟D�O�_^�dh"V/N�E�w,�|i���X}2��4�����F����Tw7�W��w�:E�ǓPXd�����ҞKF�)!,e>5ٙ��8�4�2�f��Ka0�hh�I@��D�y�f��UO�u2�j����ò��Vj:4�����-4|��d����	A�>:���U�'No����2� y����-R�}����/����L��^p5�t�~�]�֌�BE���Oٔ�Q�^�`S�����	>���VB@s�,�L�.������N����]f`.|���� �霐�l,�={��ͼs\l?�_���f{#|�HZ>�N��m-���
l�?]p>p�Fe�Iɼ�e�5�1�ulVb�ұ����Ob�*N�p��l�ʜ4�^U��E}!��S��с��jՕd���\�a��WzR��T~g�t���LJ�ųMѥ���t�韈=�������u�����e��(�����=H>����o�x��Wx~������2}��4�?�T�����wiV�V~@(�$q�C������fn��>W�^�Ɯ vW%�w��ĝ˩���|�Z�<����9���z�/���z5�������I����>�����'���^�WGW�jSm^TE*|����H%C��91�=^U/���5/���[�W��{ۉ�52>�%ݐ����*e�%���@�����
�E'/��Ͱ�Ǌ^0�#g��P���nBh<tHe>x����&��X�����Ҭkܶ^�xk��d��J6�ez�t���^�怩�ҳ���S�_�z�b�_z�	��3���+��^({�گ&)d��`�)�r���m]U,�w+$�W,|�H@VW�&Z�����ȋ ��r�l�<���6T�C��4�����T��-v�EӸ��O��.ø�H���ѐ����jɅ����c� 7F;���td�(@�(�>&ȶo�#�����6`]���^�/ @񺫍eǆ*aYЀ���}�L��7hc
�"3�����4��m���
3a|qtiF�e!�)�����[꬛�ęv%.�7X�ҙ�b�S��_2�{qM��(�
�2�㕩�E��=]荺'�#�]\H_ԫ-'7�C>X������崞dfSH�<i����vE�.���Z�Ճ�ۛ4�e��ጒع���!m��ޅWqO��?��5�jAo<�ʻ �&��+�%���:C;}ږ\�q������D".@��o&��ц�ڠ��� �6��řܥt��S�c74I��o�ґZ˦U�&���i�z�O��;�T�L�l1�9����Z�;�R�zs�B�!��[I"�(v�	ҹ��j��z�Z��B�ߏ�R� �B2��)K���3���r����_�
�N�r �Gq��x/y�?z�C��0��gp��pos�o��'"L�|AS�k��������?e�Ā[�о�FЪ�q>=G�5��K�gg1�