��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&���V�Ρr�fm�?�`>O'� ����=	珛V����M�����s�h,H�ک�M+U���h�:�-��,���NP��0ҿ��oZQ��z��[��n���L� <����9߰�n��Q�%��O��� Y���K��c�rxl;hJ5F�m���J�2�W����T9�o������u��:��Bԕ����0��������CpM�ˁH���Μ0��[
�l�9��Y^^��,A���A\�Ȋ4��|�uƹ�������" �r?*Ͽ��|k�a3�;�3gj�
�Z�q���gS ��f\$��yB�o�Ә�E_�� ڏѠ���7�M��3���c���R'[w����f�X�C�x]�e/�Lºc��Yo��L��{�㑟��	i� m��4d�X�-���� ���Q�{��Œe�ϡ��U�� �i��^���HDn�8�;�9�y�%r��'��Z��Ѱ�ڻO��>�<�k�02ӟ�е��dX�i��v��r��Tq�~��O����rew��kx����S_�L^���9�n��p-���~H��'0��C,�����x��O��ƹi�V�_Gj�����8�p�I��i+ta4�]<���*Kc3L|,p�:�8t�EI��ɖ
]����Z�W�*|��๸<��K6�U=��A���:���
�xQȃ���ߢ�m?b
�J�G�J����M	�f2up�*�K���/���j?_�1:$X�7js�Y�l��Y�;��aٝ/�
��\m{�a���ff<6��O8�w@j/I�L��������I�\(a��]�.ƾ�E竾#�ʧ��/v��$m��
�_0:� b�������G{�`.�sz o���?���QLУ�&� >��^l%]]KI�4@;�rܽ�*�dk٫����sZ@�nfEM�S��(��Z�gp��G��H8�m��h�2��mQ�n�~���Q���|��ɻ��_]P	�Œ�6�]>���!��M6ʏj�D3���4�T�3��;�Ͼ��Ҡ�ĩyU�:�;�[����)$��2R�R`���OH�����ݏ8yl��b����}�L�v�NCIk�Ų<����h@4�e<5�a�ʬ>�&�"Γ<
�3���p�Ĉ�.%N�}^�==3;n��!a�����	�=�Jg�%�jyr���$!<?>���*d�&���b���U����5{���"�S�P��2+�L���R��Vx/m����tJ�	�Ba�5��_F���~��g�J��fvXK D-M ��ݓav�4��UO�ew'h%=�ޔ��\�x�#�xԃ[؂�gr���Ϥ���×n��E+��1-�~�������08������i��pt��'m�D����o���n�R������·ą����SC�a����A�$��-2[�^����P0ڲ�r��ǭ0��ڷ$XIgL�̌� �ܻ��y�B|�b�|}뾨y�FPe���w�!^!�I�GHJYI� ��q$V��*g��>��w���"O5���٥�E^`&�K�{'�����[>���!�1�������5Fdt[�B~>la3m�0�wI�:�wNz�P`�)�}^3�D�jo�A�j;���K_�,�RV)�~5�]�z�힂��,��]���G��7f�>�Z4QF?^{y3�J��fL�է�ab���"~E�i
�~��~j�|'��/�S�}�%��X�C���TF���	�Y@�}�"��k2*�G�y�<mFs\��c�T�,�O��ӏ��d2S�ُI��f�4�����t�_��,ġ7V1�~��Ճo�fD��������M��[2��P#�a�k���<���L�a��쏍u|�+��l�/ʮB�����м�����4@�S��Z��+*�d�`�j��l�C�q¼H7���K;�&xcL>�Q{lK/ЛV�������An��2Gܞ�er��S�\����jҽ⬼���|mT��U>�)�S�N^y�I������nq����Q��Ό}V?���p�ɵ)��U��E-Ti�|hr���A�I����Vz���$�o�,�c*�g��yV'+����.z�t�¿�����OT��A����Xo��������M�CMl�3�_tz�b8sR��Zx�c\@ ��J�&�ߍ��t%�]�G�sN�u �9�7@s��A���QlxNv�!�ɉ��8�P2~��3jN%5i5d~��>��Y�OȶB�QU;Y�4�FJ�_��|b�@w��FCz3 l��m(�IJ��@�Ӥ��@ ���n�������BYވ�A��.8h�\{s(_�Č��P#E�Q��O/����e��FBM����7�PK-5���im�As<��8�4��E�k��.�]hMp���2�[{����TM��%J�J����X(=�C|�E�:8��r��;��ٛ_v���eJ�� ��㤓�ʲZMY����(�<�-o�m�1i%�1��O=����c�
���Q�aX"eO�W�̽�X�%���(����`C��@ݦu�pw�8�*��Bc���;��)���x۩�O�2㟶s�3`ie�m`��?��&vȍ�	·��&*/��g�C
;�*��q���gX���5	7)���vRݧ�J��1���f�ǖ��Y��~p����J����V��9��<,�=����3������=Α1�7�'"�u�	���?�W�A��gL��?O(�~����]Meq F��3����8��sM���UT���c�Vp�o�hu²�+�^�%/�t}�r�g2s�6خZK8&s��z��|�H�A���T+��l�R8�9>�㹔O���ח��,v �dc����ڵ&��s֮~dR|��X��XF����6���h5܊���Wέk�7�������B�k��)�@ݠQ��Х�m2SmG���kg�վ���q �	�S�5~vڦ���#̺V��<�Eq
N2��$�ĉ��U�L9��͔ikD�:0M����`A��ȍɦua�e�˳���'�I��l��E�&ZPR����'5�N����u�a%1G�s�Ɋ�]�q�H�-@�fK3i�q7��K�4��+>8�:��l�Ʊȭ�j�R��MRu�M��$�ƶ��@�ܞ�.����\򝣍�R�Z���{c�L��(�릫�����Q�͔z���H���^���}�E��X��]!ۥ6�`��Me�ÊA���U$q�����07o+�J���s����@)iLP��z���Ć��%����RQ�K�Z ��<=.v��0T�t
�;H{9,oڱ;�[�ȃ[d�-�)ҍ)n��}�0�g�g~�#��i0��	{[�PƝ0f
�̭����+��@]��o�÷����ꔾ�#]ߕ]�J�𵯼�W���d���i۩�Ճ�ޗa!v���h��6'�I����O>b%�&O͐���s���|�fd10k����3��(t�b �8��^��K���u�n�ő"=q~=8��/T���2.�6y�WT�@۪/�~����k��d��i�۠I�mk+Cm���qZ��=��-�W�ȳ*������`��`7�����e����r���G���7�g���f�m$�?���_�a�+O���L�'���m�y��!��������]������ڍ�k�D��h%�W�H���Ș�!����Dы��+��Ȕ[�$v;���[I�fE4�J���W�ѵ���G������oW������м <t��Ie������θ�@Ot9���9=D�5Wm*Hp�S���qͣ��A�)Jp�j��	������](F��U��݅޵�0©*|�1��  �m��������C�t�| }b[���W���T7�B%�`�K.���M���|���	ۗE��5G�����fχȜfUN�^Ԗ��a����|~��V4]���>0U���O�������j�~��պ*��Gu��(�]TW�����IX.��M��p��5R�A�󻀤I��}��3��(�=��w��\Q�
='m�k?���.����&�׵���x�$'5L�EnL5oZ6�f���pA徬�9ᆻ7H��XȪI�}�W?Z����P�� ��w��2���)���	,��� Q��M�(���؇TG�8����5�G��LTL�"f�]ϫ!s֖Y|Lʃ��q�L�-6�@��\J�h����ct9��[�k	��h�����ߨ�O	�2I+��qU���5Wt�8 Hs�:쀘���0���dV�e}�T
3�2�{�v�!|�ۗqg��S��K��3O������'+IB>]9hkq`W��URT��8�!������P��?(�D�RU��������u ���
{\o>5(� 
o_v)�R�;�k� �m�O�Y���A7���@�}��z���'�^Fj[�4��o(���I�U�-r2��� �
�g�(�}��"��<�	`��f��Bt��_����K�?�D�ġ�ݜ�gwP\�@YR��׭9�o�*��/pK�0��0[ɑ��:�ʜ�/�`�.����g��F>W^R�5q�ct��~-��@ۆ�r���6'eb�uG�U���Rc|hm�bƩ��\����ejvr|���W���Ly#z�g�	��Ot8��d��.�J�lb@*��KJ�Z☱�yy �O���ugW��|9��V��@�=�G��g�G�2*M�C,Xþ/��U5�e������V��&5b5}�/�!1�y(�BƯaj�?eOMn��1�,Z�>y�(�j`o���+�1~�^I��3������2f��&=ͪ�w���T�A�_�bTOp�Va/��s����˫Ƣ\i���`�j��r��& ��Jr���f�w�Ց��O�%����+���,KK� :���v6H�ۅ���!�3��v]��S����bx��j-�}�X�3�ĨC=�A|!��tS3�4��m3��X�oi03`��a�^�z�R�o�|�|���g�KI�s�R�;҉�my�l*����1��D�(�D!؎�����蓂y� HR%?�+����v?N��Ǒ?B*�d�;ۑ�(C��G �>I�G��n�`���m"m�z
��ru���
�k��i�U�J�_ b�W&6�[v�AtU{�)4uϞ�0 u�E��u��4�kKS	�)&܄����oc��6(�Zl�:���ɮcb�D�_ս˖���7��ӨI�W�W�KG�8�Z#_
E�2k�o4�O	�'@4wmp���[��b�g�����!r�����up+ :�n���#�C�֮$��Z����~{�셟���	��uYyy�U�w��OR�AJt�.H���_}x'�h�F�X�ȅ�e�Ӥ�9� ��w؞jm��I�J���K^L�v�����!�^�S�(wҷ�"��T� �T��h��A���: ����5�o~P�7��Ҹ�0�d����l��<����F��a���]�O��R��Y��t���/����u�w�|� |�i[c��\�K�ɓ�C�@�R,�^]8* P�=���i�Z$��m,����.�o"�����ɖﾞ�ɑ�GEF�� Ak�{�/�CY,4����3�K�|פ�ZfJN�o�^6=�d[�߬�GBJ���έ���#eY���Jӱ�&l�D]��+�����^�]�_�Y9
��iU,�PZ�'d� "����z�f���6���(gr*3>BXB��<�m�PzD�f�$^�k�nZc��b����D8Bf�H�����ـ�Zo,�94�ks�S��-��TtJ����+�5�:�{pR;S�\�^�۟�� t|Yu0��1B�����b�QOM2xu1�vB`�-�
�Ưx�'q_)����,�o=�iG2��[��f��0Ä��@����°�n^���x�a���x�+R-�\v9]?:���,`�V��G�;+��RJ�.Q&�,aXdOS���e�º�2�r�.��9����P���F�s��P��-@dn����6��)g�z٤�Ӭ���y'�͓q�h��1x�O&D�ŉe`�A_��l�����"̠1y�WWP��ܒ�TE�s��Q,I��-t��]��O������$��}��?�d�i�<gs���?1*�z��������W�n�H��iŸFȯL9