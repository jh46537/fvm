��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{Ns�ȭ��+{do�;��F�0�S'X=�2�gП�5~��P�~ǜ�U�\xW�D?�r�wF�@,�_����4%@P�Y�Eg�ع<�Dz�h�]�J���{�I�����:�_1�s)e��<��ԥ����@F�\j��V��w4q�t!�Nr���0������C���),E!�]h���9.7AE��t_W!8���I|����e~q��z�h;�7�й��G���3ɭub���n��dw)�a�dOo�y��̑�wn�/����$��h׺B�)�S��V�����44�/���k�'h���˙��PriF���5�t������Fj$	�sFX�6�y[�H�r��FY)\(e�x��`-X*&�&��H�\�
G�a��}U�	����xS���|�y���d砿��u���N3�W������+����,�������/�,;e�� �A5S�E��Np�����	+��Je��L����Y�<��D��I��IF��z�S4L���rN.��=��v��\�����R"�j�s� 7�L�.���K�8O��Y6o���m�Z�xtn�콟�Ͷ�M�n�./ϓ-�7,=���x5:���J q�n��_	���Fp�[-��ބ���C�jv�����zgh�z|!�: d�8�1}�
�7�uퟁ\�%G4���~�b� �o�c��sbޯ�U����>.r���:�Bz�	R�BĤ�%ŉ��T��1��^[?|{D~gk�����m�����.Ͽ=���M"f�)��'pt2@��"8$K�jFw\���&F�Ѥ����L:�۲�)���E�N �S�U ��g��,z￭�n?^��V����8���W��\d���k����{�2�ؙ����~�Hu4M���D��4�!�i�f�找�F�6�Uv�%s��1g�Љ���R�Q)����$	]9�er8c��VӚ�W@`o! ?	:Tܸ�v���?��U�+[��p����$���.{��(��Hܣ�_��U��a``�u�/BȜ��ؒ�p���3a�"aꞑ���ڀ@�}���fmp�����7��HT2��%68 $S�?:���b�e�|U�^R���w�a�4q�*� �E0���B v�%&�xc��E�z "�e}��� 4Vn�p�	��@!�ԊW�Ǵ؝�!_���!	z�!�m� �.a�#l�
��'����E�#�
���O��w�!!�����LJ���ۅ�A�:{��սE7;!��1H:��E2Pz�g`�M6[ʬ����:��L斗��8��X��=_$�S�w�C����	�b���$Y@�R�jOu�hD���}4&3�Ȥ<�3�Q�;@��Óq��%���q�����D�t=�)���Q�s�tK�*��ma�:�b�6%8!�(�3��Q�ʏ�p��G��3�Gi�<L��;�� }r�1���֜">�U9�w3�f��L
|����I'� ��/�^��(����h0tl�Qo���$
/��"���3n�'�k��
��U1Z����l^��4y�T)8EK��+�i2��ں ��o�0�৩���v�/��tX��{y�^��B}̝�y�����D�0s����@�Be����V�|��B�f��/޺�Ml�`���Ts*}�в2O�/ėK�A�XN$e���9��XMN]���c5{l��nT��E/.�ˢ͈�l^8��ˑsʾ	$o�q_9���V����\�]ջ�OJ(�2�X��!t#D(`�t��G:2x���8�j��)��he�>;�F�m}��B�Qc0<CK���ʎi0�Z/ h�\�KXcq~��������&�6��е=�x�k?�^���NY�r�b)l��\��\�ƣA4@����B��"C�^ns|\���F��l]r��^~Q�C�K^(���^øh��G�{��.A1�[��nB���4::�������N�&1E�g�<k� �ƛ�K$��@����|�(���]鹮-HH�È����3O��{+|��}�Eq�����=��h�������$�X/$-���/���r�QE�t����X�=i=Z*3v�+$������CL��m*�O:#'E9��F8a
H��Y,"�p��N�.X��U��/�Ve�_���K�P�����\��q� To�[�/�&��kڛ����=n9ſ����������eHz_�fFw��{E�L����϶u/�#/��-��Lc.ɾ�BS	?� t���W�i�~L!FF�o3�n����z��O_J��,���AW�)	4��.�N.k#.���z���3=��|�����!�dQ�or�>�������h�8k$��O�����Y;y3���}X	�M���oNX����MG���Î��n��}Z��h菌�xw�2Y&0��įz�覊J#����&���H:��g ����8ݺ
y�/��v����������QI�(��N���_������O��?%��{�e&{YԿ-�B��7��o	%;�W�ǧ� ��[�/�e�D�~�j���/UǪk�M�N1�'ڔ��W1\a��Zb�L[E����.�F+x�	-������L��j�S�2�yYR�E�/,�p�%u{�<On|Ӵ�g&DC\ff�J����n�1�S1���:�H��SaLR�a��ݙ����v?��ñG<֒�4�[��(�T[)<�����(��Mevo ��8�{�y$#e#��{+	����,4��^��̏HL���Jn}���p��XХ&������51;�޽M��K�S�cS�dhzC�5�6��]�(�}�/����[K�L�zi^�_f�EBK�\S���Q���I�c�8roJ��t�ۙ��AG����eS��@��*ٿ�T���@��"�Y�(��C�:l�!��rA��U;p1x�V�>:�m��<ISMƠ��XLb����QW(� �l�T�H|\���&��k����`� &����F��������x^�h	��+���Wn-,�d�g��I�K�}����(G���n��p�( �4��5C �������#�Qp��4i �g���"d������]��3K���?�Ӓ�ފ[�W�w�^�%�w3&LJ7=q1XB�����S�hk~��c�o����B(�h7��a�m��L�j�P��r(�5=��v��ݩ�'6�c�n�{=��}�%��˩�O�ep��0��plz%Mq7��}ߩqQ2))oT)��*V'ګb�T��v�&��f�⸿cdZu%�E�pt%��$�ms��"=��FS��վiA4�f2���ɯ m�C(�}�+���f�IU�6V�w��1�ڜ��/�:�u�審X@s;�+z�U�=��4Q@dG��U������/�?G�V _][�z��