��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-��A<�b�3gF']߯i���q�ʖu�Q�91]�p�>�	���_˲
�'�5g��Ə՝���v`�ݨ�����¯�ml��	���d��bi��nnwq�%��7��#Kޯ��ҹ{��͐3Z��~���
��:0�1�ǵ`'Z�r��v'��ՄC"$<	y�|�?�����{��h~k2��4\�����<��J��%�Y%��g�6CЧ����\�:�o���}��)hR�ïSoW+�x*�����*��-��6��	"���ڿ�l�{ f�𒻂Y�T� �W��JЀB�"X��&,���}>�.q�`���}#
b��p���t���g� �{e�����.���$Ƿ>��z�I5�:��>�V�h�j�(�-�VJ`G�-���)�jE�[�ז�R�4tM��TZA�D�)S�oX"Jk�kL`����|f�A�R��	�Y�v���z0�~�������0�,Crxn��\�ꕀ�V4z��� O�]V� mu�m��z鹀@�e7(�)���]����g4��B���G�ՌZn�(��0>Ŋ�$��������`o��J����88���q-'քK������1ZK�nq5Ψ��.�?���b�-�m�l��#�5��'������#Sfn�u�3B>pş���v�K0|RL7�w�j��͘������k��g�N5�:��kM�u`�_���!ܯ�%|&8���	�sQ�=ej�賽�v��hm�{n�Y{��l��N�>Iu5ԣ�."tT��d4#�g��0�$��˴��ʁT�4jd�z��vS
 w(UhFB[k��3�ֽ��8�s����Q�ѓ 0,ĸKuŗ��l�Ͳl���!���;Á��U`��l�Y$�%U��N8�
�r��(3`�Y��#��a�i�.��~���p��"ݎ\�����;C��>H���(2�w4����yrzWr����d@1$���C����?OV?�Ig}1"�њL&�>&������ڱ��U���r��/{����}%�|Ҷ���L3J��uA���G�7u��^��Ö&�:�8�7Z`V���m�0\�g�SV��qEss#�K�A�Qh%�fle�7��?�I��gT�9�����UG*j�������8��e�v�,���H���d4�2`�	��_<��(Lb=��d�8�4���L�����c$�UR��N��?�Hm�����n���Xo�`��6ﰷ{��N7�o����<�D4|ŧ,�8��ݿ��PU=��B�['��d��<9��ȅ�:�ʝ[��%�K�B����5i�!�4��m25��Q��������Q��@pĘ����/y�;g�����xhE����6\����0�V�3�<�.cJ�X�lf߅ϳ�mBC|�+��=:&����m ���91q�'n-��S��׈|��y=5UCuM�t�����6�0T:e�����I�Yz�ra˲�+�\��)�1o �.es(9�m��e��8�Dɿ�azˁ�/�'�_WR��Nd2%�o�Bt�ɹ��v�U����wCc��7/V��kN�=A���|tF�'�%��V_<ŏHa����h�I�Eh3�Э�ҿ��U���O��f���*��f0�s�֋���BD��:����9(�%o̴��0����a�w\�N@�̓�������f�JM�U��(ݕ�9l��V+�.rL�d �-X����s�1��ĜλV˹;p���Y_N*�q
\-\&5��O;&��a��S�܄'�U8a}��b}+�V茬R
���$�QWv����1Y'U��(��z�@�`��?<go�8C��$�e������wIN���.�{Ǜn�d���΋7v�3zz� �v���F��I����l�g�����
H���¢+�Efy�]��^`eJ�ۋ�����axp�Ey���)�r�.}���í��O�='��(A�)=��gn�k�G�Y᧣@䘩xcxy/�3m�-J���f��+ث�L%�1?�+�R?�w�nI׍ *)�VQN2��{���$�YDm�X��B��8�@��ؕ�Шvs�����-0�a"��x�C�ؕ�$����B�+�>�ō_c����}g�O�2s#�$��U�%/K�o!%�I&("/���(<@.�ɆÖ�,S@t������TY��{aq9J��q����׃0M���ۈ�ռC�	�	���Jr������I���@��`�M�]�vjzX�N����"]ٻ��S҂����E)4��fe�� ��H2�L���$�d�<I�!f5}�"b���}7�a�.VQr	$�t|m�]�I�~	6�3�>�������Q�ʃ�WHfǠ��Q��8������r��2��H������D�n��N�k���ͭa2%ɓ>OyH�����?�4�ѣh� 7F"�P:���"1�4>ޯV���~ͤ��]~;��n�8��Sы���D���e^�桑xy}�<$~ 0