// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:18 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Hf2/LgsWldK2WUmI5jcCgrgCC+ewYeCQXg8aDTP7LT/UYjGeBEIeWGUl0CUAl/5Q
sCG1fOwr3MwJdtmAvrkEte2biHT2gUflmfcvPyw9TEgwHEzsnNJTBusbh2M2rPyp
zyHJr4HzgCXhw7IaCXQenvm+cgytqL7U1QSdELHvJk4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 26160)
O/tcQj4ipmfNVWJyHkLJ4zjI7bQ5w+ZbgyyzHsCaVlgy3zlR5uBJHun56X0/KtwS
TOY6mrR0JwvkQQDKQY9REEsW3c69DkNhREAe/MO1tFe+iox3DAxYik3mNwTDP7CX
TrDEpxllXipH7ALm36RPCuY3Vbq/Dp8DT05yfeVjITWHmVJ6jyP10O7ORC6/38nV
a8tTek963R5i03ctzOI+177BSxUA3TQn+ha5YGg3XbkmHjJ/EugVZBUeYUW1gxdC
hDyQtQmhY0BLcnS0Q2Sv11uxudwZ0Gv/9bLfXFQO+EIfk4n8MH/SeY4cyBiHcvr9
y24MBarGhq9tOBVuYdLkiD2nNEhUOZpwftr04gFtlKin2sKJW24k0D0SK1RQ0qbv
UTzOJ8wTkhDjqnFTzR1jQRN0x6d1mOMuA5LORbORP2liJagBqYiYr13i4FlQHoSR
wMcs7isPFhM0MNNMUIl0PzA4C4zTVyeR7Xo7Qbj3Z0fEZbtbpjc9l/m/gi7XZgVo
SOfRQvvCX1DMB/lE2pm236I/ao6FNGOpd+fvgIQmnb4Axa+tN+mtv88HyQmzNBH4
RLkZ5YWnxdEZSlwwD9yIDTvm1UADTzDtRuhlOPq4p051mywJ770ZuKs1PIDezvq9
A1uixV17iJ3xSUoR2fS1h8JCrbnmbPtj67VWepyzewU/7++ST81u/tAY5SkNMlkj
C9d/OMum4TqTF6YJ5s8dQyed+7/TL1OLDokkSp42RBQ5GOjGWXYTL4t1sVx/jAhs
P9eQ/7YLYwsIYXnrs0q/I3Y1El5+PUxUJVRr5WqyaiuMcueX91fF2xFZRFSsfL4W
cYnyT7kFLI2mM4nvKSSZXAAsefbfNc4ZWaE4Tg1PJahaTesNqN5/y4jm4xDcnhdj
JNTNQInX1r/jLKipiwbKdztYLYQc9rqFq9fjSDrM6e562HVcs8950h32yUQwd/M/
1mQv6aEwfYDX0+6D0CE9J0wsJYJqq+qStmetxs0xqtbKwzAXH05cABVxIV7CaJcy
999FPy2WNDkLiQ8BnUxu8zPMs99zVxDf3nYxHXOMMbVX9OZRKuZ2LTG0YEIAQ2lM
yLw6Qp0bB7X7lm5B1hlDOmUm9oQSyP/m5AZnuVeiBN9RYtwjZ710fVgpipjEhWvb
iFda507Df90dAO9fQyPuj1K4EgUzGOITWJ5sY9nSpVP8r5mATduoegdxLK/DCkEH
KAvW8wvqnkCdlZUT6WyaYwagUlK8Hc0U0DzaBzrPXfo7Hsw2dxkJ9tGe7t8XolqQ
YZViMWDbP7h34NjSahadsfkZLq1uUDYb/YwIpnBbaNLCIWIXoqshtZSMRySrucpz
nQIgXsqZHQdZE++LdyL6gkQVXJz1B0DvE18VyPOtg8CtjqRlAXK5d99X1RGrH/eX
V/pU5Taj1UGddRsKXYWXV2lNtzoQR9b4QriIfDu+DnUSpsAHgwn7U0W2qkmNPm+5
idqnGjN+iRyboVx67uhgmUxM6xAiRIOHCE6rLUDixjXY8quUAz5133KfSyF2ayW2
eAFU8dD/zjBVH0vDkb9ELmzvEo4ZnDkJR1O6NI0+csCT3sXQdgfNsEzVWjj0d24c
FIAK2M5G1ohtPlRMcpm7BrAlpRVtqhLdtZwTPUC82rmBKxZKU/thagHxbmsFsCbF
OY3JtdTTOQqsyzrWctqet/pQKlCXU4GDeKnZYXA+SryhHgjM3jmVwLJQCumMyKFh
AP849loEpRj5MlgKnj61E68fyemmRYmC5qqX4bYvwWMeTmNa9vPfsWsT3KGTUgdF
eeI02iuokCpkQRv8IzN1JszHQnTiErmASiudiKLvbNlK+ziOYpOjYR6F8P+rYvtp
sjYUeL2Ve6AWg+nmleT7LhJIAH5Gi/ImYjf7on3qmJYqckqTsFdxiXDYyPNU84eD
D85FvyFw6s5qRKhwyc0YWL0H3E7FvSpMF/t2VU41L2wYxRGl+oqEOujaSoFhugt3
EDsZOc5IenU8wICyDlDngYmTcMsjxKeOIINAoZ2SGJfSj+EBQD5wKmczxkH3m8gZ
fNV6C3UMJ1SJJ4EBNOauULb+8fzoxy9UV3WySb1uZ7wZgNIUKJ8a2YsHHfVRcyqw
H40LD18fu9ib1OOB5X4o3tqvOaGT8KrWgOuyu/E4BrzaiAPDM5OowVkV4h0MT5tJ
9RUPcxE+rfuuARkn03EJ4MMtWWzR3X1KThncmVVSIF+UqDGIC8fOupMUq2qCi62F
c2NMC61ejF7R9VXB9zsJmx1Lik01q/rkyM57y1XDZI88M8SReDLns47LaS6NTRyP
Za+vD4lTIgLOgrQUGOw35yHVcicYnqirqdTX2taY8Q41QI3O04Dpg+A6Wqx1y/xN
0DRy0C8Xf5dkJaw8JvvrgOXSLYCWQkXaB7e1y9DUwKgrOohp/AjRAhmGLGpgQ6NB
hNuTGmaBW88WlSUcAxKIdiwjE01EMmNcYbOzVMh6T0viM/++/6F+UqtzlmuwZf/F
d+qLCEdrAD7ugLN6l1M9K2aaz7QP2D5GCo7zaoTgC95/6a8jCktwcLpt4VsPrswc
/IcFI3vvCaD/nGspCc8RvG+PEp+QvWgAQQUXFlPXStFhILesqHzcdlpMLMLMnAvz
GpJib2lPm6j//cEyVLHeIHIXdXsN1tsiOzF3xl7lGaMA54YnW+JNalFtF+YdOkj2
GcdJ5oJKiVe5fGPMWnE+O6PBjZ9PAzxl/gsylNVn7R+RX6+bi1JAQJkuT6bdt8e6
kLKhjzaVzNHCB2UOYKLO5zg0uPnunz0rDSmMFjjJga2M5FpKoJIQx79fb6lFDOwm
LoEGqN2zYgbL44N/xQwjToMo2YgnoY4DVJf2UiuWSIl1fpvO9Ou4OGICZUY/cwZD
E6FNNOb259eOij9R7UKCFTV9amxwB+xlmeSJVZMnzdVS7/em+yJOXrGDCQ/7sJtt
PXfKcVYuLm0yoeA0d65K+6Da9VY35D5RLtvXwxV568YN7d9d9ui9s2nPEU3hSHo+
1XMOAAwTW9QpOFF1+ALuEcDS2ZFHxDDfsAXIvp/ytHy5Kc/YMRCumBF3O/hSvFPd
0L+/ftxO/OzAqBkcny5fKSztZi412E06XuMX2JB+yYhyEvOvqgQNCDto30PMYXOB
08iekfn2ZOqp7foaMVVQni4h8xXYmwnujTJ4kJhkRXHIZbCs5Y74/gt+DjEP8/rF
pmxqQnjXn18NTG92E6WajP4x9tMPpGYGVSsexKoJFMlwFVfHVPUYXZRfftrjn+kq
usSQkCHaze97H1SNL9g1Ok9obl3oFDZXIlN4zUrRtgSFq4674RO9GK5JRky73xQa
8z7xF1k7QsFwWORzRVa06++0B7y4tc5wYzHiM6A5IoYsE0+lzb6zPhIv7aD465E2
lRwb24Rq4UDIjfpJWAseY5g1geYCJSmIEU3wXcf3QtT3FdLdiltVPouB75rI/Pnm
cXqoJj60VaCtyceeqHUenTNBpYfKbRnomnyJ8HmU4JB8Evn3gOFfuBlgg0MIudBm
aCq5T42V15SBu23GQsTTpN2Dubw0k9u8w+SlkR64fxXj8YI/3A0Wfn8Pg7hMYhT8
OVGP+/w/eJGkWTEU32kZWS4Ck37XO/xP4vycnrTebI2rzDEu+xhGQjHhruik78cX
6Lgg6d0EGIwDUVaRDm+hnDXzQL6rpekn+TgLdsJ038rJBrjSm19qG1qJgdY/pk5c
ZD3i9pqTi3NveHKyyMcGd1xXQuWVFCQi9Rtpgtz31H1NBviswIWmP+TJHvmUPvso
VuVnZ9ODmtU6oC/bt0/3NGBBWi8/AUcGX6xRC+C1ubJhL5+JMIbeXBvxS0/qh66J
bC60c2HENQF8y4tcgC9wVT1o7QP9L2tAxp47hh4d1ReTc45kU7p7S1VrOP6BrmEf
mA0BzfDa06Wwq5ku9Jb6GJdYA9bdu3/7a735i267hwwyscB5aKaYX56JT3eb+i5y
0QqE9VaK+EKOiomNTFVK0Nm+RitFHbWO1UQprvn6qxyyVs+EsCCw4n6V5ez35S2i
EEmEcB/fiCWLtvoFT5uqeWgRXkBweeVJz57BeOC78K1+3qi47dpY4gxT/GuXkUuk
runUfWXfn74324lY7hJ/26675CWyd8PYTGTTbf7OXa6thN9H89K/gecLYTw9qrtG
o7UvKIxTPVsb/P/3WVxEIodsnzT0S750So1t0lGh23sKJYdg/yfI2vG5a2aTQKtW
qi7EU4qjWZIZQml5CxXVm33W2iv3hm8Prz72VM6AkEwuJC5hwjy5Z5cgT4Uff4GX
5/nV6PRxEDcIeNnqFTFm0U5L+TRXoQ5Pu5uetFWpQmxJ2X+8eBHllidJcn6G2kay
YgXoQXZ/obVzufR5x4RgWKKL8jfahdlbLUA7UceCOO6OfYL4L0bMlInJpUWXYhVu
wWS8xdJ4rCD/+rkNVJruFTsYnPBaDrohTxuJm3S/lRlAlg61BNQu1LKKRrK+NQQj
3WbYwmmd/syuETL3BE27y8QkszyQvh4N2ebT3+ROXgL4Q385t04ay6zJ4W1n/dj+
6t5uDk0HqS8JnIeyn0UCbQ6all14ay6WzNDzf8VH4yU5qEBWSyTExVw4aMGqiSUH
4/Hftbe06EJUUJQ39O79o09vgDKf+XYXbyJbtn9cQo7iioVl9Il05F9U5q7Xm93d
rs6o87N2a9WmNR4/wHxeYJXi2DeH2unkkXSABBodgAAkKEGoeOfSaEzC67cvNdfD
a1cpSAfgT10K0wvzGnSJ0UUvq4Bs8LzBpUQdrBhyBBuy4aZOXS9pYpvXsELGj1wG
edtCZKTK98K3c7pOYJwAZOCn7QiZBWLf46pKuqyJdX81PJ0AJZ03wv2l1Q2u3R/5
yigJvsucLLkgbforBCTmZo85GwhXZhOBvqXYo2gSgzxP9xq/+WawJx/TZQ66ZSr6
yQ3mblhVkGVS67AAeKsKDDAg2E3OKLh/B9Pd7lWfdzLsds8TOkHVAwZFM8scP41G
LJT3FSYLj6lT34CAiBN9jiQRSaEzpGPrIScQ+lqTCDFtyZDdHeT8qjhz6rC34a21
QhfTTS9SiPP9NatnU+Y163lqrKb6MTQ+j+4GgzinObuN4+CrYzrPXj+8LwUOD9VW
jaQEkupmo9maA+Lo1imtkEEqtejfRdSEGmw+0wgYZ+WBwP6YQkI9iZYu766C3uXN
Ft6mgEmFyVWNr+ZhNpOlhm/YiCrVeo57H3IfVx4tLcCwBNy3he43Kfien7vkmCE4
ORrcIDwvTI5NspEjuGcL8ul/j5PkOAxj7kW48CD3JZrGm2bvqVcNO2Pq24MbzYrk
msIveUuvnUgF8Qh3jLlnK5rL3v0cfin9/Djaig8B7Wx2AV0Q0NbidiC0aTPrMOsr
l2U4vvVN+ZJ4D/68IwzxlrW2cefSPKvDZyUauhaEz0d5EplEKVoTe5r2y0E72bVU
I8YQWhyk8LaZqAXmmLJbrLWF8ylSmtoebRWCHhUua2lRy/QaG0nj6Jj+OP27oLZs
/2kwAnlobT1C1IFfi+Eu7ZXg/8OtI35m/d1Ee7X3HrcBOoa6TPYVxzOTalKb7XFn
iofnj0MhIWprFSsJgN0XDtrc9r8l1etxALyx2TuuwpBvV2ozBYxxeR2xv26nhioq
W5FiLFuc1jpH1SVx5H7MTh8D0s5xWFmhsfLmcxquCK/UKly8Iuyc4eOM1NjtPQWU
76YlpiYZtjJ2mmcyWt42F3aWtb/I1eZgJvaq5Gu57q1WvPd7mk5rIro1wAAc3Jjc
YiGXbeYGpxzqAyPZMskR3+iyv7b3MYUBNtApiSBqag6Ii4CKbSeouBbdNLRO/0iH
YKFZR6kNQUstX9mllX23eR+lp4YePQkMECaxFy56xJ5y3rX1eApDeD0nzM3yPsTM
2ropkJ5iruPOVwts8KeASlwBy8lAGHM0AD7zuqhah2Wk1liviy4GLXGwnbw/HBQb
GEU5xGuJbCgTHXZL5OThtREVeA6IGvdTCEVyBRvgXGhtaLpbFPSE2IPJZGTlfkCs
AL+aiwKN0ExRqF5tS2uPtgbQ/4GhfVVQAKZ9jyXnbgKbqlg4isqXI9UTtZt1jzKR
ovTrqmYowic18SeD4kcJhpRk1bmkCc1246/+eIyDoxo/3OOrhBVe4i1qT9qWbcaH
ojCQN1pVo5OQ2z9gZSmluQXGCD6X1qpM+9U/85dLQoMZVY8zzAtkpk00a8/zD2NM
jKXmXK5DbAAQI0pZpLOebm3bChqldOG2SHwLzwrll+SgXkrWX71D/XxVZoupeQ8t
FCbUGzqMU7M/Lx3MlHdCxdW1Hu4tUZXCqVN2N43Ft0SBq4iQvU0JrfR2/2EI54mc
TFoHk3c+hV3hH/Q2B0NoAQQjlLwU0x/EF2Xms1bjNLLosXNQvMejc1TR6IMrchKt
y68UxISqFRu7Pc+jwLJaso1dczjRH0VwmPEgluC5bdnoM73qfgCL5Ec55wTI0BXh
HV81xiUqCRwrlgx2keV7T4e0U1D/CHFyzR+choY6nFuqgWxZytIDTzXnkMmd9ZBK
zvByj6hpC3zjS1Xve1pJJZc6BXeRc3P/TDgP3uAfjJRdpcCZBL9f0NQUbBvjhqOA
s8ZUEYbMAyGTjvld5jeLtgwvVa34abGQnQxaMDsDcltSAz8Ri2TCKsKtZ3heUZYj
C+Kmla2Znct3/jMc88Cz8W+8Xju3WJ9j6p6SkVWHFfJjOCrR7W3yBQxB3cTPl7C6
hZsSMkrMRow8g6NYZyknB78ckZGZExm2MjAJn1S+2j5R0UMMkkKkiKd6mXXnYPpl
3Ey6Tywuq16pHBiO2XTDlhEHEKIRxhxNUX0OUDzNDbtnZ3GEs5XEKCeQZn1mtSn8
fQC9AzOW2rjCcwv1z/YnLIbBiCvh49sx6Rx9BHiWuLwuIZl/gIysMGjBYnS390K+
Q1cU7tEeGRM7KlVyByA+Hk2GTqfqYIlySGwlpRSMMHhF9+LBiwsLJuskp120ZooV
rWh4fv8hB5nXz8dFytagYlGZ8OQow3v0AYqzrnVZZlV1nRl2bEdSoweh/P19mazy
NuK4wFM346Bo0Qks3j3KVjghW9Y5bI38BXCRYDjfZBJTzRSXo5Bf0fY07yIv+mB+
JYPJFCNXrBJLWO5jkr3If2zWtjLOiK5w2V/YHqfVaC84FnqljIw5WyAhJTFkRGVr
6ktktbiogqQ6caJ8qd6yPU9WYrbnMiYmQhHaPKaQTeJZ6G6DqIAH8M3cgK+dUHMz
+pvOhnye3x8RBkYBeDYxVFkBOvmWt0eLTTaWUhWTjgj0L+NJGgq5nPpwbWh7I1lG
ZYu+gmLUjg1eqQxpBK7NKz3X9Y9IUGym/FSlm7/89YJVitQiLyly3YEr344NCSYQ
fdizK3b35N9JUEVCLefwmOngIkse5aGqU0ODK07aWtbTHYu0B68Feuv/p8TGSSUC
kkYb/qNUY8p4J9Wg1rYSbPg/a7tjkw1oltq0Juxy0wPcPQnS4QxD+3do3K9Apzqa
KmoVNG4KZZTRSb5puJB6BY3fcOSZhCeJcPVR8tsPdwEq0U1T/YmUveIROOyViWxT
iNX3HoJHjN4LwiCwpt91axRGuKj6PgD0DWlrlhr6RV7GC95ChASQOr7a33vQL0Dc
266r3dzYzQOlwLTaGPD/CX2sWsmQX1cFsKAyxvsYpRN9CzFLGpV2r3OOziZzIgdV
lB08Ab06IaUv1MbUVhiKa+mw6DMXKJSCZraRcu5UF4espUZ5DqOMER5hHNj0Wb6P
EPtNhRnWHa3xlAysoMY8MregMHFBvo38Om8ZYFade407zCLV3F0/INNNciOYaUIl
3R6V/Z+7W+Cbnfve79RxZn9Pq+asBD09MPGvZ7C3FVkhiYRXCHE84KFCLBuwGMOi
F55lB1vDt8GWZ6bYdB/tGmvFJJ9QPWAPxsHom6UgvhRmsj6Z94MIddeEMklFkGnu
NOglWuL/pLd5BoYrEVcLhDfM5B4liAq3LTliTeSCzjCKwYyS7EU2kuVhKP+8ohvZ
K2zLHnCfOef8HursmuPVZIT9YOxz+krBaQHBW3kGy6/fVgf1acWoYoMqGQmRFTk3
emN+WDdUX2WHPTKiHL9EmkUQGUYD3qcYxF+UAppJYeGJ5ZwSxqQRrgKcTUZ7plAx
PI+RFOj30Wba/ppX4ujOX5qsHwRaMCv1Z/zMcSy/5twlKnrMGTrv1ye100/nGgrX
oLyQXC0oZBZKQhr++qVBI8V63aqeQ3D6J4a17iWfYToFujaQ2Y1GmlukmByQ8JSd
rUu5U6SjOwK/eNU1DwYlhqtH17fWw+kCOEpaeRMnZXVV4YAMYZ0adzTD1MvhE2ot
NZC2tZS3ckREI+IID0s4tdnl6HaHV78BoZeTCXjmpxkSgEBTwGqLwSpBqQG7Ztus
MsaiKLy5APLeQZFnTK66cBVhmV3aN+Q9ek5DdOyNU2G+yPT6HJYCTtL5e9/WsNpI
dGGz+mOOR51vj6f3tVM0D7JYLuh8ICo6UpmIAjRe8jENfxPFKLCFa0xKp4/BV4AS
Kudt543BIh4f2D8RWhzICJ0jhgKzg77w9zoxBTStDLZaSr0nKzqS1f74XpK8lUs4
M27qehg/lq6opk2g2APlfhLI9DrXCvFh+gF1kqgpXMwzlcXodCwtaI6waaKL2DcI
S7ZvpU7g95O7YAXd+Av6oEvlRh6VhmgfOUZ1FvNkp8kWtiknzd79BY7fX2ogaDFb
S++WdxqZSKpEoIocNkyDTFbJtTwFpfttRWXsjBtfTrcTt2JXuj9Gpca6DM6MycJv
72fACLXmzIGa+x5VEs6lh7Jr8hahNZy2yiwBFcuP0tRLoCb0ehF6IcGL+Tx5/CTE
2GvfQyCRqZxLV48dJ3ksCATvTqP5MdkR91rtf2LCq7TxzmBUndVkd4mLp1S9Svdu
SmhasnFSDwEg72il3z3KwLyLN9+B98DypWjwisRngcEIrjGepu6fWDVhPxkjtidv
y4OJCvMCNxiA14lHkk8vycarX1aSKPgegdzcJQJOX/dTVi4LYfvyt+2sD1LvOoGe
b8KdWSPXAjRms5PlK0YKszJqNKgDRx5RiU7Ip8srNJYFgYj2PASZBl1OvTnvLkoH
fgo/tEyXACgQXkBi4dSpXbdDkxdtoCfnaDVorFLj1Ho4WBhfiXYVlXAF8+2SevUA
vdkkf188FYtCbxSTSA/lTdhL0sWNLKh4ZOIYWQQ+GXmsuMgCJQqO0TjXVyoYEfA4
p34MS8CB/Q+948/xAVkzN2sJIQpKw+NJ4vKw06ok5G4nULLD3GTWfvRj6DjfgD2V
XRqQbLsH4QRN/CkOnjVNVWoBQyWIvdizSUkAggFD5bjM/oH8i8LpIf5AuQbFYrVG
4PU9ySBj7Ys9GzGwUpq0B05MoiU5Og6fQipYrdDD42nzzsPxKc/ggP297TnxAnlG
RlPJIB+FxXtFUBdrmcq77/iOL4k2w7RDZ24Dwjt5miA+qnbCC3W091OOZtfeL0L8
R0FMo5+7XXKMtcz/SnwG0QtqEUoKIpflTgR38TMY+e2oGgxlbz1jA5vVHz77zm+8
/viKB4ZHBFc2My2dkEx3087iCwDwu0MOSpNOE+I2ojzmuOMwmLXVru7DfKyisB7t
khzmQN74nrZObLXVr3Cv0lsAtO2sA1MJeVypZkSsuH8pKjrINreCFfGaAH0Yr98h
X3AuvPDVNFljbovluMfFAqoaNrrahNjPFjlIYCRTZFzhwigEebgoqyPtVRPPF9up
EXhJlVt1Aw5qb1+6ORxwqjHyeD3AsMOsCXnKU3ZAr+ciaDBjmc0CdxRmIoKVinwG
G7lRDCYgkmATZ9FpBLGiFRs2HsY0aR6nM1ISBEXvi6ptnsXQW2V0zDd+ZPllvFTO
ve1cgPSxoVnvwYQjJ1fAz7B/y9muBieMzNibg8+Pqf3SDqQMC0UrAndVh4C4tYZl
UWNyFVxpKZgwTBFmbHV1LmyP2t0XqKvxEQGe5ZBtFm0yAshqHt4M01SuwwTE1W3t
cXqZ3ZDRC6fcNOZpqcqASldTwcNyW0JjjLd3v8WNqvZO5gaCnXQ2eR7NGdt8ELbL
ukHUfvAmndByyt2u81EglbVvdPXsD0LS0OMlgMhC6JmKEclHc4WM1a2/TR+A8WD9
e6Yk7NDuHIW/bbErzfa1EChJpBlEYAW8g8DmICkdrL/ksrT6X/QDhpqNdx8wRnck
74/3aiT7A33w9dEnMA9miHArp5ujCrXcWy536UjSPUIRKE4+ZGS6I4ImUfXe0NkL
ASIaHT7scwPFCXpanpT7pd8X+hH0TGozDNWDRGwtmVLu9zx0pYWiwpHVd92HA8C2
28rlEO2M3QQYX96t4kA2O70wZyPMu0VMaA41cYXALRzdryk9q3Xfx9Bdwad4RVsu
eJfyLaLnwQgbDtKyJ+9qbmIGfHjK1wpryRt5Mp6S92cgutMpnJK0ABh7Be2RhB0R
BmnHQMbzT9OE5i7DwUESbLvyfwkDuCtDndJ5Pe9O6OawGFfaT0Tub2MwJp+sUZNs
Vako+nleVqJA8CK5pM8RAr76mdrNR/yrhI9lm/LKlv7w3ECwGmkT66XJK6PlkqB0
oVrq4RJ3HQ+stWSqi0aBN23AmExU6ZAIOAChXxezXmXAQ4HDZnV4yyV11/GrTIhw
nigPOy+/ctx8F0+hsUR2Crtfse5EvQTuzb2q3ApuLmz6uywmoicZWudo5IFx79sb
qurGV+30Wg3cLUHfMGj1N0Li8lifEAEbYmmCVxk02ZRac0UBt4w2XuqzbtMAJCZU
E4Htj0BM2EAs6ObX/K/3EMdQeX517aDu4/LD0WD5zYWuPNFkTF9h50xWLCLebpXF
6TBl/fCF9VmL4hcYDwfM3cCakT10iGHp5oGp0JDPoFYWRw5DwaiCKd0YU8YcjZ+7
Pz/tVovYH3M/wZIahkaHMStHc8p69Jvc/tjlmGZsDpt/LVrycRdrSMXqR4voqJcB
5xDwfdMb+ykHEcOxwq43hrP4mGXN5V1feFchDni5JbBt0CFQN6hXZyc3v5hWLUv8
avdJw3ebFDynx7KjTlUQHQG0Hjdxx5FZBdJTApyo07sf5vz3abxprUfsrBYjxhyQ
M1ziz9NrXTVS5NRw1RTKkRIb5ZSm3EC/0trS9u00sD20ZPDLIUKR66zksb6ENifa
NQSsT/Eh5FICx2nUErwcQ/pE2Qz3me7CBEwMwuq6/X/dlL1MIWKFCpAPLFwJqV2J
2p6t9hxFZyppibjdITHdTb+UpjaCWZpaSIedd+DdJRGlb4Isn7h+2gvFBm+7MHW7
AfJqLuNzJJTU8pOjWx4Sqtq7KhIEYCo7L64hDtaD1LIAHSTmzWRbB5UBWJ0HTv1P
2FfBn7mrHHDDAxrLYWPblHH1w9C/GVT7XLihV6ZkX34yS6B36MLm3rp8E/uslC12
kg15mItdErU3jZMrtxkv6J+osySHgxfJq3wmuaqUG4DiCo5t01Gk8bSkxj/ZTu9z
waDQY7Rq7KIX7XNVf0XyluZ3gat6OIzs1HyyC0t/1oczo7s+AbeiVexOr0sz3Rp5
JVhf57J3dcJs4mPr5QoEP2WTLzCa6hxjw4DnM9XwahJdOJGYLUuMkSftjpM1nklq
eAaZANsDHp/8EM7muOmPtHCxEZ4VchBUKN1qX/thsv6uu9GOdEC7W6RQB+EoSqkB
IFAb2pOIV9aBJunCECS7BkOY2Znl1Un4vHBvRIK/CB9wF8paxxcod8WLTe3uXfzq
kEmsV1v4BKta2S/Yt/V8Ghjja4obhwoCpIFNlaZG/vpo+1n+saA+AT5Khq6KWvZH
Qbosa8xI3U695FE34KDCsVUrTiEBnR+akEEWPrK7P5NaH2RceTyc3/lhaVPENmgF
k6ThzntKcAQ0p5nx7mbI1IDIt9pze4R7B4siN9bCl+VHUG3PfpJs8PHgkCC15m1t
3Tlg9sECCX++E8d4EwSDJ9067QM/dvwRYFwc2nqmMZcPlJDBdbrfpjX/BeMxjctA
w6EyiB07O5dcSgqGo/ORQUdhMK5uC3RjE/ovzsI07qfk6fMYuAe8FfG8/swV5to4
i2wfEiy7QseSEqcCpLkWjLz1HzxhqW0lsHRD1UDtBtD0+X8ZZ4TTqMesxus5BFcx
7xlmc/kyWTChJJAN2+rZk2HEqknSEURRnQ1m83emh+Zy2uOVNiT1OBB5Yytw5lcb
5U2uMLMmB6ZVB57xszoUtG2Lrf9A9D5gHy/Oj7mfJ3H+XlziKvDy4dwoIH8dJVdL
O+fgCpggXy+BV51IgFNZXRvVCVdpIQm6MHP1pcVG8uLu6ZiRG7P1XSiZdpttFLGv
9uiFX9aV9KIMdsWEYy8kcwGuKiU8mSDDNDVQiawipw74hwQFNK0KjQ56AITT7WyR
fTR+G50L6nVaR/ph6De2gDoHgTn/ps/9fwLfEAKo3zUr+I3oVfyKWgAaErkywvg8
QoIPlpvLuv3RBaEMPaqzGAzqdsJdUynuXc5MCt7kVeCCYXp7c+1NaQNyKiRuQuN5
FM0jG8ubb1xmZvaSnbkix+k9xQL8yVpgj5CZUt5T2T9IJMBs4KA0COXVInp+fw88
QY9ld7WpyA30Ou4NRWcg5e4TgnbBNMhgomUrGhC0epWY9SJsO2QYnT8DWEZvPdfn
p1KfujgTVQMbk4u5I/W1F5TyqCxc4o/fY875YCuZBqiHG72J6/ZNm8vGcXEywMkp
He4tjmaGSNvuR0yljHFYRAyI9ieDtwtvVlREFHPEmHLQJ+xwIBwQsr5rtFvdYqYE
4thUJCqlztB3Bi/u+GSc8CfzPpADk+Viy3+NKm5K1pHe2u7eTMJ9ieFma5HBX4cj
Po6WiYdKWAGXUVvw0jJf7epjGI1cUEC7Ldei4LrxmSHTYT3cvKCwQLHzzj3MTZxq
RMa1EtarEauXqJfW8T1iZ4DU+RwSxpLoVWLKIf8zuY8kg2z+yvJ3guterVsKho59
/Iwleg9TwxwpLWOyUWH6uy6BsDMj1DzjkCYdWjKa35/aZonbS9hvRpJs0pBgj3pZ
EhWjVBE7S2Sc2JQS/NCnha4e+9Y/XFZppzR4q5wSCJD1NFFhlQPwNjzZ1CwbokKk
dMSjrFalktUmD5nUK2peOw7JJJiQ17DnlB7S3lw9pkuWkGamq7ku/mpzl2vFpnkT
YU6DSkQG8+oRVwnEk3ViLWSYu+Sb2bHb+TqoqBIFP2kMz75dcJDgEmPer5QgIHXD
PBvE7jaV1n1JF6HNcNuAMUSLb96tQ9hNLRLfc2xGzzLs5yMOfUFMh76xVTT3BbQs
mZJe8GgICNQ+vvKTwvWAsxc211U/HbRW1CY3l/m9XsxP7h/js5IvDDls/rLIc4My
yjD6EO2FosjgDlc+LDvpvFpTDgDr5B7uC0KJAFxvFqUeqwQuFJM9r9uoYODgID2d
mcACA+afBNY0+YVt9n9QIxRgfQaTTmMcE2Og6LLr7EmoKY+Np74CMUvzOX5LrrKZ
Y7TOrle9LKRB3nk7HUxNTIAgosjZoK5362zPqBmFjN+mxUZBQHpkRZwkvbmR3eAC
TW+fkwl3YdgozLYuei98z2gSCkI1eAyLGvHbScyFS1y9TC476VnAb7jsodTqjeKe
7UTphvTYtcKjQfYa08wZqGiEnNnJ/CqJ3PRfLNrKDWD59Y/+28E/EX2oWsqUCZZ0
Obkfg/2Mec+3ojDQ2JuNmxCrwBpyaXLVtvZSRzsGBEu7f3NdXVxRqXs5sEcwqrFX
aXl1+E+vXE5FldwDoR5uybGbd4Vtv5gS58HgX+DXBDOE431c2DdYwZ0rD0DKeJEi
o2GxU5Q8GfABg5f1wga7ycFMtmJ78CybsTohgaxCe0ROnRcXwkVu223AFdoeLM9o
FCP0MKZ4IqaZYAIPU/i3g79OJyKDdFsZLHTqPa2Ejk8GUH0sr4sagmGqv0SBXd9y
JYlcY2vbNIuP3j1ko7xXdTR1MFo9T7Q23Usn9cgVeQoRX+D//at1lQVM0CjgcD0W
MiQBAyy9DRi6tFBPAXeULPlHo8h7ddo2ur0xYToiBKo8o/xvp+LqN9QJKvpS/yyw
FwfJrsS6N7yVqHy64NI4Q9hdIlL1MFeAmVEwHCW48D1w/6B3AbHwPVwUNqvMMab/
rjs0TtgPoxi0gCyWAZFuq6NciL791NFMIdmlsjZ14uIsrpysfcMT1rDmPd3KkdHw
XMsXXpy5iEqbr25+aCzbwTM/O6MVwKTzg45An3jJOIZ3AYitqgSKZxhLVrHV8YV6
CyVhUzmpCReCGf3RzPftP89FVnXQs4+RctAZpgd4x1dvEAVarfHimvmvcJEDq58l
edNeLpF4cRUHgqPMrRm8uOzXnKEiUIGQTRiDGdN1XMOsiWl5mS6wXWjf+VlVJ9Tz
hQwf6GpJ24G9RIjZG96RtCPABbHDuHaNcZmHrz4RGp7mo9Vbbs9YEqw5Lw+H9tNA
T+5zwLZUA9I99EIhR/Ndn2MOPg/+CJJBjOTbZmYXMLnU1VpeqHZWPU8cDXQ//H2t
EWktzMhJqEqcShN4JMrulV4L3ScTJGWdKGFBJPc3Tjyjbf/zXUacTRxkdBgPtXGB
aGcrq6YEqLzO+QeuehoTy+DRWp3aw3moHX/qU+s74+yl5wv3lTS+IuzLKI/V5JEs
YrY7trgGqWuN1+I+HX6zU85iVU6f3ISlWjU8UEtj10Nz+ZDmJiEKGI1ifBBbezRV
xTep36HJrDwGbWrMV6ChRKm5z4OQAmc/jZh/JSWJy8NiQwhd+ceQRkULvFTxcQnw
ifEF4loNusVJ4SFB1P//bjn3Gv5GVbZIQAt2HJRpO4A7ockxKJip9JNgEsnP/tBB
b3E3E6wEtpToAJWSjz7YeVHoQj86aFNzRwNIDxRkdeH2TzaDV6H1OULrOXTAf+Ie
oo/wsw+VHr9/0m9aTvchKdJlEVey5uA2BJCHO4wG8aviYvieFMcFdEvoX8VVA/F/
PHHYDbwyF0RB0L6hHn6z3n4j2cWl+8A2VfqEtd+tYnBHUlBLCrau12SUAndfsQb7
P1FJuxvF0MwfTGSx4gqber6BbkWvefoGADvghV4gGif9WbxtViH6zrHcjIiYaKA6
ylJSmHXNqDGuXAN7qM2mMr3haVSqPmsylcJkI8IygNpBzDqs2/NIVbnIKs+WPZ+T
UO+kxX1iQUdNQhUHRQKIj50zlIJ+rq3k1xOjGnwZsa/ftLg0wrLXN7CAva9LlojQ
a4XeBzPaFyxQNNeviPVpqakdNkl1K2+WBC7DOd36eLO3BigOTkruRewDxnMMdlQ8
aHrKQetZkNGjzDizcHEcGYa9765u6hyCl1+9AXKIvpNL+1JZboeiiXKmrL1/kl0s
WZdm9h2FIjpax1/jBn7CcJTFHapiaNy8DrJArIE7kG+nIDJu/xWFiEfdVkPnpuW6
I1aoKtyjS4x/RwkD7FTkEYiCPl0z7wRt+lbqS+VSiqtdt0whxS5I0ppL4z37qRW5
LU6b6nG3MNCsTxGa21Z4RP3zSLMd70XBsWkWFoPnUz71asacaD8B2JuV59PTGjEw
jpoBUbGq1/IAk6iVh69LASMOe5q7paAfeVe1A9N/iKiCAvCTkZgpgxW+d5lmyhCg
CJ/XTL/+QL48I1raTl5sDhWI0+llWOLKrhdKXvjTmT0JfEoFdGa4c50robRNnS4D
hvX4ICqmv8P9jCOJnvlOCAx/s/zWqowYCBNIFKbgnvgi3xSWvxwY46k4jyFKWqs6
l4cZRiQ56xAbS07l20l5YWoWCMH7gSEXT6qx2Oihyrhf+O87Y1PhN0Yp9yasja5/
WNbeCbFXLJRZhY1QE7PAfgR7mhPQBrL8ifs74sspbOzzrf27dFl8tJGKPV2z5Erx
8Wjyu76NKIwfaoXLOZ5/mOeYF9JoU4ZXl2g4jR6ughiB42Hq4N4MPB1wUpolHt5G
3UJbEPr1LtOAifJcQKe0yUDQr1sxZTVI68AMn13Ru76Ol+p1waYx3fF5S8p3OsbN
T3CwHfzaZqLnmCijL6aIn/0XY0ovevdE8xv75egaJvGTaNa7WMbEXnPXtn21wS51
yTWj/ioxDI6Byeikn12m2J02+mg7cFR9yoKB59z0EtRYPpnbpbRwphdtmG8VTjjM
+anccmh7RO2X6q9WclWAT1uoMv4wGOmCDeSrBzf7zyxtgTtau4oz3/1itP1MQrTA
51lhpMi0Lm4Ng+eZHNGR9s+zFlZvB0dp1wIHLMMHMMT1Lb2ACvcY4u97xkWD8/G2
DyZ3UP9fNgLpVdRbtmPZ+URYR7VoUQLd33cGBsadD/EARYqg7NucfY4zmZjXCI+5
EPbRLw5TXV7YBK+RWGhk07hGTla86ohoX54jY4W0LyHv1fL/1y0lpeeb5tcZ9aZk
qBLnNjK5hYa1H9B6k3AxewrwKbGIexfwiyWOQiPF+AvGAl02PvBCfs4CnIhE6cDI
xbx6ec1O3lucYJZfolrYb/Rn750GEE98FnkVXgVnkUqEfNh9fxP9cZ5bwvNTkmUL
c3swwHgz2eKFYpipbHtP1qNymnGW3Tb08DeOsPmuFaXjje7p6DT06rILdUeDEtur
7jl/OtZmRFu0JmuKdL2lwOXZrWwjrXIuYDMYSsZxRkNv7XDGd0T2NcR35jVn0ys8
g8bcikS4vhg/Gn2H3G/1Xf74jELsvLyuIY/2Z0aY9qSb/GUPhEdXk44780N6y9Hx
hUwY+r560kr0JtR65ngsYGfAVJCLb9ETdF/2SbqGgMjRtRXCCnuir7Lp7X+CbkgO
s0xlHBoUsYhmVIF8d+PfjloHEj7hRW2nElqwAuE1GX4voDoBhITShQgKdN12HAaO
k0XH4hhj4cwaeakmakN3HJ8BlXPcPT4ZFwUU+6ab0o72XKCaVmm7QVf0L3YMcIzo
Xxi0XYXTHdMf+53bfqt/OItAiFb+8pIZF7bO5337RrX+oPjoRvZatuaMV7wfXAQJ
ae248R8RoNIflPxDFUrplAA0Lp39jPBw5bXv5m67KA8AOFNppT2gZoq7bEQB27He
VUlPlha25uXPr2/uudzNHx+xJKyRrwqPT29AeNnGyeSuk1Ee9NcfOH/bVy5RTqSC
ChFbZTbZ0LTmc2IZaEwCbRU/mJczoTwfNeT2STs1sSyr+LcfBiMtHCBeuick2fAp
fg+aHNAkeYqDT3HsJBH6UmYgJj6cAHKGtAlfgkVjpI87DWx91cHhmTSlJ21j2RQk
P/RkHV4fKS15ASsv0nCE0fXDixRAeeP3ddUu4taAWRyDHjHD/hzXXc9XkwitRIY7
fM0s5kaTbH35ILAQptmWzHVDSdcEWj4HaM3G8LQp6Wb5xsksYy0JzUy15plRNs8n
IR4mtDg0CO+j9EGFB9kTRu5/WiDGFRHsY6Jh4AA+ju/v3bEqSExf5F2dUeIPPrHM
q/BTV9uv6q9epMZDxLPW+oIZYj+lRuxnrQQX/F7fNC2kYaB3bGP81fc3U+Xf1Ymr
zSw+JMcRu0ws027rZk2ZHpqG1Ux9s+8eLEYYpia3CMZPuZUuFY1JAVQ9fP6VDLvz
29dS8C+Yt5ze6uGuTnXjgOEyXtDmvt2bbZ7MWbJko8NB/3PLKqNy0dnAMN8PsClY
bBoTzMJUeXr8iWE7K0IZ4XRn4sBIdNZYFeVBL7yHd0QhU3Bic3XdO2fiTPxltm0y
7fun0cT7eZvHqU7m7ZRoCK65g9ZDl/ADBALTNAGSeHd6MLw5pXNwTWlutmX06kbW
sFmbAqdPpgGcje430nqvzMUBfPyQikurmBtnWqNUDtXbv7fLDRm0pWkPo3+JNxio
3C+iLYWeRH07baeansgsLpUUNW5h4TKW4Z45c5v5TcFc/VPFgM2f0JEq9vaiF/4b
ErBB02eVoo2K8kfXOr7J8D4+ffZAIVI7wBR6OpFC+UmT0COOfD/zHBlTKnQTV5FP
8QTLGdoIlc4wjKNStDv/1L/94mi0rXruz4+6KKiPbnaSvlR1EafO7KET6YnPJH0V
tf7H3gv954RtX7tr+oLJqVOIUgEc3NTlrl9P2eNQKKzcJcpqJu3iWs1d7Wzo+GSn
dk0+/YoynG84wVIjfTvgqGUcbS2/jPDhDzCBgugFH6jITSkX0xNeHJmujoQXv4Wr
uE3xT07PORq82NEX8K3jjD4AShAJ1aI566I2Lfbf2o2+lNPNdfcVZ+M9esQMAVzh
LB/3YGA9+mpDIc6tIIS4sEzsOFzNHbt6BqR15JUe61ZluRaAgHD3lBo5PrRxxNXQ
rHw0vbOYYZzyohW3eqeIf9s7OpekpI9r6cdOTyHTGBATZO9kmmALKBvF1TtxXw7+
25LzSNui4eqe24m9IvE8dniwyM++xluWOUS6tTwctX/mCQIwkOBjmQJ3xKwqdhZn
3i6MjjPoX43eGynajEs2Pl36c8uOkNUlWPX+eA1y5afNpfpDM4gnDW/aeXCop+dF
YVz3s8ezI+zXl9F9v3RwpPuDISB2mlsSWjzR4xW2GIzHZGUARYsb/94hFRso2RPN
09Akwx4S4KZSsnSR76Y1ZIY1GMsqKsvrKGYs1DP48HNKZKoND1ngMf8ZXU2S0hHi
Bmk1zEr4BobSK1MoPDdi+SB5m1uix9xsJQTV6Kj8GbxpFQDUY7gVMnKnxIiJ/npr
CZxvtVDod5GKKK717XyTMThcuHZYrQN1DForSl7DNQwEqisCTim6+5viuRnSVBNL
4gu9jtbXNGJiXPnZs/z+5PeMDaOJeAVJiStSAPz5fRzBHhZgrM7/Vu+Ai717em79
SBGqXdcHfZRLXcpuYtmvTORetU63ClsAfn4aOWbnCR2ZdOIhmb82Z978gFSOXEmD
FXmTLndiiJuiOR8ZJys7wnUtevAh2xpWvseILu/8Pn+3271b0AaohO/jSDY9IByc
S6OQUfneLhwrkqrnxjoeb7Rt74d37nOsHGh+2WJ2Jd04TdHjxNhKu9qB2nK/ihVk
jzKPqH3AaYysXbT9fiaQiGwhCljcbEfC14kOof9Zyh8g4sOx3RNSlQwnRCVk5jvg
DIIxs85xVqSQPH57dS2NSY8v5Kzwe+nKNIKSVgrKHEIwQfK47mpfOdWeZoZ6+Qqo
+r5Xk7+lebfAtFMcRr6p/qBmArSEzwd5Dv/ckUI56+siQcSvF9U6cUgZdcNb5Nuw
BpnqJfbgy1AWJYuXWQVa9H729NBG1D2kKTAcwQjSq6h8xIIutroBHkjuvbmIZ/hI
Lk1DxG/zKaVJC2BHjvVHaO2oawfySopGeDAXz8dKORH147yzOgbTgTHGDDmoxSiY
Oz2vbt6j7xHz2QQL8CNTojBPcmZdBbdfqk9VHsFAAu0udd5fYdF/G0c4U36coX/P
jnh9DK2kPs0c6z4m/WJuSchpFlx2A1EFhSXfPr7tQqIiXO2ELD3et20l2y7qYphH
MP/nlJKsZYJXFnHjmJ78T6B/Rree1ESzFON0Lt7Zxhd6DxLS8HBC3oqLOyXNWx2m
FYNQDKfn21I5W808uTVhEqZ6Gqj17J5kqhCWL+yyOoHzuzxxbgCYoTDHpabnlW1p
6qYwCh121Qak4bRJGCfuaBM+QTLaawGjTbEtyh9TEvNlixSKWxlXlMeuMaIiovbv
0Th5cqOQ6liY8btSqTddp59/zDfhdlekZw1v65hZygaMcRKUsyP42eaWXEaoQgzV
OJFSR5M0sg3wmbfY8U9gLL3k2XWAmcKww0il2f7SOyZoGlCAZ/KghNtrYOyn1C3O
OWHfnEheAmZYKV9JYVJBKjAQYshAggeDzyJiWMPf5r5y8gnZEcAeRd+b1X+JM9aC
C/UZcAklwTMRp6Yt1cFysntYNZOs325CrRvTm/HeE0a3usR1zxcnV+E6QAA/3LWD
5CtJbUdXQIqa1KF11bj9czwiZCHNMO6ool3e6qkQhjQJiK7E9eBQOaUhHKqwcLj2
gIRMdA6VEabiHgzMABDfG2zCyuAVUIWN3N2rs9DkezU6he4XK0+d5UGLPyOvnjY+
L0ieB96cvn932Nnc/LbIhEJVlce75WZ+KzXS1lU0/C8YPm2os8QvfmDqaw4dVwU+
oyRQzIF8Qeknx+g0NSX3rHG2D9gOOStW/NElmQL8AsVhjJga2lizdiFGYR6hjY7E
5tu61bMbg2vGnZQlT/67N6cExRuuNefe5aOwF2CtJxAH0pZxMlKkFj3L1CuWjGsD
kT/1/XI4zbbRk+eAJkWAoZfjNU5OPLV9vpX0KLELiDnkrb/gHcOaTnwIKZVM3b8A
0X7tnVf0eGf6977svPHxlwml5Ry3zrLNHGLCgCZ+Fcvw4TOilvRdqrx7if3XDKY3
L0pT1haXs3HnHjccZmLWszvmYt3UjHgeAO0M2rrybp9+x7jyca2UMx0RiDHRQ/0Z
aU2hxN6zph2Yl1ZsL38Lut2vJMi4r+/CsYYP824uloKpReYYlEzh1fm/Zj4U9DJb
enSWB0gyRou6o9XKtn9fO4p/LWyf2tHKnhJEMWEdyr/CQB2B1nZovr1PQuF8LYgM
Zobb6ri2VcJjYp15kbsp0IY70hmxiBIMq6/i2M92YS+GVPFbsNrYoYCmmzpCrYBA
HbGzJwESGuJLBx2j7OomHBJoIgROFQSzqsrL+hIYWetPRnVadeQ38V7voq5YZTvR
S+htmH7gMyb70Bz9MCG1GAOxzmuL8o/+rFiqApNHsvpcW4xE/XJpI8Ywxw5V/BBU
CzVclxSMGLCNpcjf5tRTo+3Pq0YKUVcyOA5Kt2ZEAz+TYOTH69F7P9n+IFLToJfB
Eb02zElgm4AyPmggUNSJna15GzpGI2MfDP+6HNcCRKzAmfPvn0KQ6oVxYAyRfLT5
Yj6AutEBOqVXOMVZHCHoASeNjvDEYEngIyzMj58inaWXiCjLkXHuGFYIcaviYbtC
MemI6s+1q5dvMwKrt50EV8q1soqmCH7uqeOkymv0SSbN7ULe05f/nzcDfR9h4iVT
IXxmMVMuj6iYWcRmr1YChMtdlcu7b8geoPtT1N1gnfVLtwN0V4sL5lB8Jqmh2G0U
anzr3Y29cqVQJ4i/kKOLOwZLje7fqa4Z97gwoMeIWygKUlb8tDIs4cLMKTwHj/e1
uityIC+qTf+h1MuGwrgqPQfKhYbccUKDkvXjZ6NMGLNaNDshDnpw881ur1dpgXEi
eSpA1dJ27tZtFVLQrnnCz1dxxi8Dyl1pCBFkpl/N0e3rIOw23VLoEKVQrlqpHfJV
qcYuJ9iPkgneLs7HAXuVwCvL0Joree2z3p+rhmVVY45O0C/DVOPfhtOYxYeIf5Ek
4YWWZ20+Rrlh96hG5AG6mlFgErQWp+oRWRz1JcK39uojAd002Z2WcGaYIUf/+dx6
PXlyUkD9Hj0x2FV6sleFKy6DbPAqnrRxoEW1N4tAp1g+EOTiHq/YVHrGqtu9+kis
ESXZeCTYBOnMC/hZRDRBChZ+jythZo8wuusrpF1NBV46Fr023NRickNbxSYE+Q24
kJ802Cd4J04yLhuVGnTjYHuA+OzPoHrO28XwjcqStTGCpzRGg22Xz4YbSHIHIqQF
S805Bb1vx6QaPf7E6exhLDYjtyEuAbKM38Ngg+BQPgtbMzP0JaQaKVKcGtdO7R5/
VpIl//xGoN7+VsGbl0IaTcGSexNB+Qdm8Hy3NnNo6onxWPUEkG9tnuineGsgcCUQ
+M0Nuql04GFlRL4bsGnWTDQA0sT6bAiR1OIUdXWL3denuYzN/gRjiozSmSP7sZkw
KKqN3MD3U5XgbmXBeQXVjm9tZ+RQ6ODcqIgvJq1prqzenEQBAz14jfxLTNwgliLm
txX999TILDMHWQVIuaNVCGDwQdN0l0GBws45kXz0tLl35fSdqXy1+C4L3Cs0H0rC
9lCYQ7/HoqhT6ub/ZZU3Rp3Mvpeo76tTyxU81zeVBde5DLAY+pZJdatp0KjL0fx+
oXj89AllMtPB1omu3qvLHc/GpzW53D4N46UqiYNt5GAQWWWbsVNLHFId5IRrdKpg
Wv8l2hvjOzwmw/46rbMwlmVStY/LnNlr0hBbqwcVI3PhOE3jHFKOeFwQz0Pyvn78
Ci0BhqLB9YNN1nekn0QrLRTN/RoEaDLBNoOTi0X1vSaBFdF1zZPwcmL3luMG4HOi
e66LAqopIE5gwxRqPaLHud/phGo1GsEhiS49lQYvXpbppJQzDLK4kleFtWUhc2Cp
6AgkPnxokbF6TAsL9muCI93+7eYVQQ1SzBJFk15Cf7BOFKGNSNF5Igzmf4B0tana
clumaAIg8xfuRihsBAp3NJlMgiVmVmB5Rh7dalhETNjYSER8BvrOf8YRzLgwyzPy
/cxIvu+FsEz2bW79l5A1pY2pX4V9XqhUZxaL2yjCEIVEdySrUPnyc81rch0oFxpg
mUsvioNtqi6WOUpUKzQauzNtcsr2AeiBHI6HhiycF7cq1KMCYeMfGGP0TV939ilr
enPqJ/K9E8IhzGm16TjL0fRvdCe5BFNAtKV/Rl+Wko4xS79acu73EPROOZv8Ro/m
5faiVsgHjLWEpYNkzPcG1CtarbgOWs3Fo3vB8VbVLmDoMflKZBL+9e6aPJZWhfwp
tWJgT5dk4MdXqLXOlTjGlkGu56GImymVKzdM/0ZPPjHg9qPeK7Sez56fPm3sgHn1
5fUIuzzertzq9GSWz/YQ2dK11uie8MV+rZ3+ecwsNANNy/RC7olg7BUVXOPPkcsi
1mVBqascKU7938ip1pp9Xqei510EqeYz7qEw9T/D1qRScfFEcA+oMjvK/gEqrYzn
1p2CvVUv3aUM1hLCWMiJUzhhBzzME57D2NdVJdAxPcSFCzMbce6rMrCkpeweqi/I
o/T0cXChmeA+eaUvxuM41R55gQ7jBNJIt1SqBCl+U3LPXl5CbFsj+6OPfLpFj5GA
3bFalkE3NzFuNOMkcNpAzjgMqMN1zRjEaixxM5aj3jI4jpZMbY6+ljiuXtoEp74P
YwL+3ES/1zbiRv1Kkwc8Zf20R5+KWOI/Pl3+uxF4uPkC9aUuqP8HQnvpFqU6Ox/z
CQIUVDdEVw27CV8TzsJpvNPUnFeyf5Kk5wYzWbuJqyY+hza8F/9cb0gs6WM/u4i1
XeWQdkXagAaHOgK2mwYClrvXLm6ArWp5IN2UqscSFERuNz25xmoP2OUnTzAhiJbC
Dlht4f1mfmOBySnbaUQPXD5X2omKT7x0GipCXHY/tUuO+jMAbPCfj2VaZR18mdTv
JXhClcHxWXR6Qk4Dg0GwgP1zcCDsTzRp5MET78IxSmJQ8ZducAIGVg2EOT4D+DWO
LGYlKcyhFiTII0UmSK5zLUh57Pv3jTmmMEdLvggpviG2KhVG9Hnr3lX6+Rb1or5D
nFjFCg1WTSUyr2lt+yHsYa/2TejS/iyOsjnBGBZUmHtRGDgoH5Iis0zNqFByZAIY
RQAE+j5aZGlNP68xA29IYoMJqV7PB7K9i2UduB4KgRS+4gnBzt2tw9SvajZuQYdN
GlicsiprBbjB5f77sNc8b8HSso4xRmk6/WL7owl+L6ml3FoyonrI/a1neTsdOD7e
plu0Y6drXoBjK9t5bYOfJMIyJZLir/8l51tc52GGMXytk9mG6uwpO0na0Xt88dyH
YpsJIEDNsw6UEPOzH7Wncme6zRMGTqSsGE6PoehR8Zphl3Nf+RFxriC2taQqKMCy
fdFRbO9vi1RHZCExXjuhwpQKihT8CfCW9B4zfJwYeOhrqZtKiKpXXsIWGG8UHkSM
ZQ8XODOh3lbuFdEWapLMDMKyDKy8vM+e/WjouwPk9KtW3V2034RhbKZ18V33c7l+
ciSwnKMRwFShM2Ectz2mbBi0UwymPUmVAWOsWseaGrixey3iNtcqbg+TIfKMFIVS
46mVP6wcBOck7+UmwBpxajEmxUO0vsUoAF65xPgofHQz5DHn4anQ5DOCWSEFqqGp
qPbjSTW2jafnN60nTaEsXgPvMtU0JekwgvLH6UY+rbJ/xr8O2zmiSQDKJxY+e5ot
eN/alihUQk/lIfUi1odkkTearurMWOXKIbN0KH8d8Ld/79YLeq0jHu+U2H6n4jhk
iZX+QbpUiJ2Y0+l5jGIxRrDL92lWFwZLIUMhJ0YmybdBi57XEzl5XjbXvXL8YLld
fSkAyVC9IBK2PQqcgC2MM/YMT06Rf+FIeDdc4Fma7QGSMcrDRwWPC7CfbCwPVR0q
46Ptu9tKbtadfYozcNUqJA+avjWazlIG55kAJc0aYmSpydgXPRAhJPSO8/H7uGkd
bL+rVNqlZxU3qFWn3lhA3Kijz+bcfiaUs4oZoZhkDRVKNPLO+2VLtz6TUqLeTFqp
KpSwPhyQt6TnoW0Uj6DhWKLZH0l14zX8gkeYM5ozeD5jOvdSDkfTD5nhtopT4Lgu
Lrocl2vsy0d8GRxC1GIsmUofc9CgxlodLmNGeKNUrAZK0o6JG9Nf8uaj/lm/7xzz
hh3y+cWlz/ImlQzsoxxAxosHFBUbY+Y1Pt31peFvV2y8XYx9+KHDGpqoX3J6dp49
PeqcN6mnNlfcMAMFhle/Q274QcGpdzJW40DKmmRYf9odknGU1pzyj6VhBPrCa3iB
cU85vvMjmiS1xQSzwIdCBUkBs5i830YSdltJRhnQrHZIE+NIVa+J5O6XASO6VgA6
2UH4EK+0AXCynRnHeqQECRFZ7slYUYki/v0n3Fhr9PfbwCqn4rZJ21AmpFQpnucu
YmPTt7R9pA9UzdCeZzjUBVqsAmvKhLgjqKi6EB8yhgPc3Kc2YSE9LsNe8wmtN+X9
yK9zLvJfWqJ2JdWrapw1vxzCSZQ7eBwa8rAFkx2lv0ab5W2+B+cd8SJ38ecYEc8R
9I/NjOvhC1gGxhtJqfdKr98+3QPYW5o3ucJgIgzH8jry01YRbB5TvjQ0kG/lAKxd
MMXxTqdvXig/IrX267wFn8e2WVChIly+19wHTxY3UbZztVkUBvqGi2H4Ie4dA584
TfDQlzLJ8YgAYhXnhk0pVNlO0nPzDpGWIJ7sOANKPIIGmGHCPSFps0GypzRExezM
iDFvTewXZZv+NAt5Ob8UN3OfY+m17GmvxA3xcPv5TSlg6nDSGowOf62ksPQMLn/9
B4grzcVd+lCbrlISQt826elEdV9H8JxENJqHL02d+goyzODpUUB5WorvexrCKDWq
/SzUuctqNyjORCnd/XgQsPxnqQ6sqLaXmBnwTBXOvNn9+IltrwyGKcgjzB/1gyJ5
v6bYY6ZlmS46GqKvopaO/rMy+5nhPKauOspBWYUExYR+k4ZmMli2kQsJCUiBsu0K
BwdsSNF4A6BK+dZxTsehBeB4nHU8U1SOPTvATJe+shwIASskqT8ww/kkG85XMQvS
lvOjrqUiiOOPFkMgwjDkQ34CLdlbOVJsypiTPIeJoz2LK5EbXnlOIGsCSyjmXeFj
JMEDt9PzVaAtByZ8dc4BHTUETY0MJK8cOiuiqaPf683PB7tYgrZde+DQFm6bB6ED
11eqQHcqTeMLYToU5uU52YdZWa0pzaqNOMKi9zpgXUQsWAFnBuk4AvH5dZARAFs0
CF9nHOM2FpG30cbEDxu7awDz/4RiCg2gdVx771akHU8WqAhXcyMLKzUdphNHPa44
/1HSsMMAYSgN6lw02PKa5oIgc7ApYNR8vrE2uHaTb90Sq/+XDmieHJDOKm23u84P
RKU04ww1v9hGS4p0+LIomk9kROKHn2zO/13JtHNT/6ZvFIAE/MgqlEUGeUA/qZkD
EZSYh+T3TF1wJwhJy0fGdi1tdeF4ZE/tnHdt+QE771Q0XzbYR6wFYLh2YfWJr/ba
tOhkUEd28gV6hBW+qCeFE4dyvIju4XmChvfakyyYSnR0Hw2qklRRb1jR/LlNo7jP
q7bQ/L56/9MCfP5/2Cj6okzTJQ/KRMh9hMLSfPb7VSGrXHm3JqPCWvQJyPyE/X48
cZDkKLvYSrybpvqF30bVEWCFQhe60tK7/sm39ki1GBASyQyEuQewlk3am43g9tbM
0OnFoMxAdWReOd0UALrT+Ih32xA1G+Q9tQtey9Z9FaibRfTtJaHouzODfg8WD8uN
qW8jIru+XDuoNLuj9CQRNz8ctIT8otu0KQDJd5v4RB7b2HVSDNdRHpjrwybgQxDO
M5zfdsXq2FU3jR2zprZyR8fTzRU5933ZtfgtyKZ10TKKxM6MheKMM3+PL1opkEkU
x4VgYswpghv82q7X5d0cj4hW+S8yH3gDkZxmHXVV2dyRRPqL5pV8YjMdaOAYvTCl
0iQ3zdEvkAUdwVrdFmhnQUi1M7KBHbIaJtoz61Y6JGj/ecC+o6Rk/Xbz+vbzZHkj
/bPRLaiNawvDqYlMNBrxsjYQreni46Ye+RXtf3oYasf4CdtPDK3AXSexvRBZZ1ZL
CQR7OVkdSE3j/mcAA80TutNY6HD7V2Lku4xKOarHZ+ZTrypY190b0zIwEx1t3jEs
UdxujJPgbPt6gV/uO/eBMvGVhASRCAr3uhdpFmXM1Pf14/5AZqsl4WpDSatw/3tr
ZFRAFWJME/jhgcDUYwRQNmV96Sj4pRDs8Fy3HRHBLASti/hYM4oNTyPh/N3lnByK
oJygIEvTFW2b90Y5AAqJds2a7gW/T7f5oZMiGqs4qbQZkXwA/4oRkA23FsRr3+Ah
LBotTzBp+mtWm08vYn5eDxvJXJNJ8zqExsVdwUBOP5I3GflukEyGMtDSH86+50Zy
CP8cbigPWgEbMTSEPv52MrBZ2OFceTNdorJ6oQ1sUypgBsTPdAWYjYWvuM2MtRUw
jTUHiJJFTPvHmRJjvcP1RKMenelaV2gLGbDgwWQ44UyiiJ3IsoK1i/Ok0Q0/x5ya
ywMwWJ4TK5oD1noE67I7XDM6reoFLCvnQouIBMpg7taK4wsvL7dkqsoKXRDjaE3i
IqHLit8RrBSxIVcfq3rjSfB+AmYLXmPpYeh3NhxlMzoFjY0e4fsAVE9O08fgnjih
SoEiEInkFf0hEs5HY1qZFMMCtJMwlDYyJUWiJpZo6OQ7dTWSOjafaUQFu4GCAIif
9WqfU3qVnOeyV4tXIJ3PK4Vtk7gE/Z1WoSHrdt8qaIiyrbC0MqC0T8KiYraJeLYL
+/3XLy5XJw0Z0DvhkOUp0zYWSpqOPLLLRhuobjlGgY9pr2846s9DOxGhRV32vyyQ
FLLfpwviBS7SkPoyHNI2FAJoN9LX+HSjqXuMGgiHr4B6g0zDiFeRXkPXdwPsRyLc
9m3DbTlyF1RDS5wmQypA4u6ZAZ04xg1dDvMOMbb2jzidtRVoS4mHrvFPcMqdxf4t
4o26WlCrG7PEwI771KipYibk5y3uQbWv0KVI69Hn4hcY4o9Un192cPrQBHbYB3yL
czRlcGXUoQbImJr8dpZD0p5w0Ucg4gWC8C6cTPI3zag1Jyl5lJF1A5Q/Q41NWRuY
x8AwK3s7/8DZTy5fnloz5Ik/6V+UzKH2FAyEgEeXH13DrX2T7Fi96vi0OZNHQJLC
knXrWOLk64o7GacLmQ0heWSf52yP65LcnICmeQRPvpWoV1rUfSzxzLzDfb0g6yb+
bELyOvKK/FvgdBvV3FWq3QnJu4b4tg6Zlaq3wppSaUpe/bg3CTJ3meZBogbNt7R/
bbVJwIokmCEdNbQ/W7IJkGKfKGZPQntyj8F6UbDaQoD5MttgiBUUjT/XbzxhPLLJ
eTdHHlIztySZLhRnCChFj1l3nx0VimXx/SyiosjN81Hg5A9jETncOsJS8dzvs0DE
NzUaU52eFhcF1FNAqDTlVNinjIhXvRxw6mQhABlGf3s+fJkFCZmX8LxeftCzWUHZ
d1YEScyrP7ycaLYDlbbLIvXC0xbcv1GuV3qZRbP36DlLlLKcSIiZOAOume4j1R30
j6jGKm/BNr3bulsbZaGdAfZEgInQ+EfnQQsCsPggor82vc0/u1eCBMLs6pQg1F0L
jf5dsToKBeGCrbCL5lE5qlqDboqUn8JmbgyU/JCA1vjePctfHj5hyXX5OQOpD+zX
gyJR7tHpqfMJguY35eMbfDblv/gWEydX8nDDonCXo+7zzFSU8tgKrAVVKfxnw/dd
9KO3YYjBGbzHR9YacQttaU96S+qoGgIzQjWYl0lSGZWLcfo/tn4iY2d8z7YOw8Ed
P2zca5oe/QRXq+gWl9rzcWWzNmzwFFWtZMJV91Lp0ngyAfdLeHe1n7Ks+1mfdEC5
aSvSqztTHX7mTOQ+W8eJUN7OMxkzFG5W/udXEndV8YjdDnhBbuiAl2T45cUgiETA
SkQa746WzAyn42aRDrCcI1kFgHvA2N/CzujTDOu47D5lLzQgeOX3gxX7Iqtkoq2x
OnXVLp1Nu8neJi8SZFnGngpzQTBkGWHCekCpeRMJM6hrDUtJZ7wis3PLMM+tzWPb
JgVziuMgjdNY/xMqmKajUjH5Vyp74xF9yGDfaB4Ai8WOrqzKA0dIS+BauvAub7y7
4f+2pBnN3TqelNq8iIc9rswMxhvu4RcRRoTca6Xw7GlSDXQdQQe72BJT2BFjECFQ
hIEAToKYMEZGJw6wu9bgNrQEVgcH08dO7wBEqwYj6UczyZwb7ay6S9V143Sbxuc1
M9oW/VulOUJESQ6hPKWZwTVN+ca3cHEcyuevcIvziej+2CSBeiyJKB35MjVdO19o
AfvlIuzCXZy9YD9csv30ojM+u3SJ6VwsmMkMw8Cdl2TH9JICchhY7hOWOQnV4UWh
imaDM92HuvYpXFEtbPi+J0dkwbdVffUYmpuJ8Mbs7x/70AFmEjSuzqwOg1OzjZ8Z
YosWWb8Vpgs4HGTGGeIbuimJe7ZyKjFxn0MeLASNhoH7ygY5wxstTdwaFbUACEjC
uCUKf0HGXiayyrpGlmdCj42U3gR3ELsWI+uKxh/3YnMyOoJQMp8ev+bB2bd2WDJ6
ZvbBfJ6Y88IOhWmMNG2bmaEBKGfrYzdjfUNTSXlHM8wdlZamaXSXfa+57aXBsMfK
YeRkyfXZ4DwKTyL0+cW+jlZ77z6daOHFJUKyFJRkq3YlRFWfMIyKLoMndHqcoJ/H
j+Aa03fd/zDJezk+YT8mPmJQYryICbWycFv/0ivdphNvmzKYXPf1lDRrFLBUrZwS
07n0XooPOEroOI5nuufCur9BZHjQkYyJAZT+j4236xUzx9nXsoGWni6A/ds3oIGO
6/0qpv6uteLPgoENyw2cTYBIAcKyA+qucyuu8PfW2cqtzkLYoK2g/sRBNGTF812t
PHygUnCIdTG1ilCXU4iQHVAgojwk3F4qXxVdMXc9xHdHR+EM7MhizCVypSBB+lZM
m4gLIKGQtz3YI2ALnSBdVV4U8hDfSlE2q5w6KPX1dFvg4Vfx4YQjMZcCSB0RJhCz
pwDYG0t4chSjp8hZ/lFRq2vQkchUi5iNvwEkdH/kuJZaWWKGuwvhA3Ttz0eaB3LD
OI5iQNNCoLGmXTdFMhRRiP1EPoP+Mmh6R/k9WkZp7QBtOUbEXDOo4+s3NcEZ0E+r
aNfIyoFydkzUh9ejPhVNseQoHf9l/0GtIhWcWheCTIiTmL4ML41t95bF8q/qd7ow
4G8bXxBFbuUGEDkbR1iOEnu29ITFajU4BUTLijGpKHrXbNtTf0Rq7b5vyQHA89/a
QNVSZvOkIUgxhboZfQ28UMQk7p9mhizuvwQaHXFqU83oJ6m9j43T3gNt7QsLOpXD
Aa9uEdEhkjC22LzleZBxETQyBpA4DRW4O1duaYbamPvPQIHmvlLM8qaedhk0DNaf
ikIged3z7r3cwRKWyzQjeJ6/gh+mCduehPCq5LqopUDfz/1zrmVGZpZ0XD0OlKZ6
1gjammA6xltBcCbm/lkgNvO1rMmHcKZpo+OnhYWKBP1fzzMHvn95RJlwA6buZk/E
VbWvGd+k6Gn2Rr414x21u544LXINjeHkl+9Ek/ypvyZLzE50kUmjdDjxO4PmpcNf
MbCjSZGhX//5BMR2XjL6YSiRG8sPnN+CaFFfvsN66oRvSrBred8xTEnLXsfpAGA1
WK+BpPc4pEMcTQDCFlhIwczSVyqFswWF4a/UYzPwvhO/sxrgXc3fzsAsXUHXZ60H
faAq5iO91kOx6OeE5IqhBCKiK1b0b0ZDLCqEBReT8x+1fZ0Z025zUFti0cszycV1
5ZaTtfMTvibaEzp1hi+MBtoks7VRYntjH5TY/V41UlHzYr2AY3f5AaVuKpS+yQxj
XBRUkfDhStin/ExItpoO1UVjTvu75D5Q648NsW64VWLi49IhD0hNFQQfdbOFI6c5
SqXRg5pKxSK33FxlpPElJCeE5bp1v3f4IFjaTRzjglb4/oFlZEzU4E6sqg2BymJM
EVoXEdAkkiJCc3nuGBUDX2kT6+UFY7zxdRnpHbmDXreTZLp6rrr8coHXBp8p3BIL
bBFZQr9IpVhJD+B7zLLylqFVe0B48Y6QQkFVNRZdScJiyFB3gX3MjqXeCpJV5Q+c
Js/fYOxGf2hFuMn9Kd1rC7eiWUNtwiG7QQ7N4aEUyy9MnMOSg0sF1kdyN+8oslDi
UJBLjPcZo3asMDbt+asE95hWi6S1w+bBWzIcUfaUz7vBIv9dFB5tTDjV8Qh8E5HL
vi7gXM9Y4OTY7jRldwm8N3peA0tp0SiHFn17LuosmBON6uHLHGwECyT8CrZ1B3XK
dEd7tImVaQ4opdlzeHwpb7huex1IDnuLI7l8TdTgfszD+dHGDejlrUQR+nZbWayY
c4aHrIgS8slbJ8o7K7UQMVPglgQw4MqFz7007U+iBwAJ1xcehOX5BGirWU1XihOr
N0g2v3976xmf9qGkuGD3/ZA9O+KTFv6iVZ6Czk08NTvdXBRp0VCcz+YSGTgn4rS9
lMBkuJLHETVvM+ooHH/L3T5W3IeDi9UM/nVv9uMidhUpHAJzbDYkDtP90eEMhO3T
79dFwmLPGlu7VdQ+0bpHWJLkUFG5gfsbjtCdhozb2GGSmSYgxCj4cfGTR3qXdPUw
xqmghwvoleXLWcSnmfCcKk2N2bibSNHoNlgz3kcaDmnlh0tx/NupqozWTjZW1W5v
rJsc/kIbtjNhC5vmkFYHiA2s0jY/+s7B3xwLqBuvVKbBYPbyGl/hxsUdWQcjt01r
tLn0v1399PTGDa1chEKjzLSUj3+WBbPp57UV44e3YOXm0lyRkOmfqzc5t2+yTueV
+rnsOyOTSxvtd9oo4fHTuyroDl2o+tszeijcfPSLHvJ6MQZehKitrlqiaj48hbXm
6QLRCU33VMFilUxxx5BneNal7M6bBRen0UUnUPyr5N0GuVlg2PWag1eHlcx5cGz0
XJ3sxj/nJrFLqSbna0gK0TU+7PpVE1sUXv71SSYFXusPEXueCrmxMZUu+2HF+3ag
cIjIVasWTcWY/UaWCJerSmcT+LCVhZz/hsRnfeKbKldTOtLhOq9+omNRwgeXIrJP
5NpJ6kBmJRu7MNdIBTnB79Dl3ZH2aTfICKdHw3p23HbvZjJdAFA3P9ivpf+IAGal
V1fX6m3EJ3sRj+3a58Z3Tu94gBzcuRDo7LRZG60lj6p+DS6Zofpf5geEINRAO/io
etike/Iv1pvx/UEnlaxZi7ol5+wc5+MsQrOV9klwISPkUeMx616zMqI9EmmAvYd3
Da/QDkcJpQD0lGmMc3Qf1tLzRyPQumOTyOhk9cCLoVt728ew4yhlP/ufO37KZikP
zXNOBbuhKe8OQe6ctoOuDDoIR3t0PGNF62XY9r5QMgJF5eactecHYBQEDjvNY6BB
xopLiB6dAGIdYgH1DEzyR91KDH+tKH9cSE/dg3uc7dVn9iZP++pP+kwoEnHxST0s
GDd10VNbCq2Jln/SFlKilIKYCLHHg1Y8PygUi+uCXQPVjfQyY+xhQ4jUmzfTcTeE
f8CT8fV/NH3k8BZnRLdT6jOsXdTbtzoLyLxDFVx0LCm0nkZ146fB/csHGeJ+bXX8
tQC1aGaUmI1NhIJ6Nvx9CTfEZOoj3ZOWHXaOr0CUQxrOGx8SvTOhonf+cSX4cGh3
meONAysYHGu+4bkr0OhIhv4HEUwz9Lnd+IXBc1IMXoCS7r4OuirVUPQ+5/82+oGv
vTW8u5GtDHS92/i14JxMBugLXcGIplyxKg+fdrQv0nnlf82uZJuHC5N1jHLvXnKB
pkwt4YywVn+qMVgm4KpW69WQBOONTqvXYyYYxjYwJ0fqEOqYUQnOFIBMrY41YBc3
LHOxQQdGdOiEr7elzM9FkG1Bfftv7HNwWJ18eJoEAkrxfP6lE5Y+a/6rla0pOZCX
QHdx96Oypib5iKdMxn/LrtJD6w9KNhVRwTX7P6hRscrIIVgfa+ERY2B5RrRZHwLS
1wJrCMuK05YsjdNRBJor7zri6bwN1k3Im501yfHdy9dpNHyFK0cDlDhx0RkwwsZk
OzJg+CDNyMWi8zDd44cZQzqGNd4/VkLIevS2rExtHL/A0s5x3QyAKDqWkFUXUGfY
rM+xAl0Od4cmD5hlMEhQDrRP2jPPBHQAnOBUFQtR+gMvCPWBP0FfumKBPC0fJS4l
7JcLzkTOdsMiBXN+Wc4XvDVFATBBAF/ABLJls4S52W4+T7vqGPkRJ+9KoO3nqNcu
19VxUjqZgoJqPt+R+UZEaOWkoNsLvaFF3HkxHlaJ26Dg7C7Eumhb4C50Iw9IYcwS
3w3BiyAUYCulszcwoBaRDaImjUCf+SpHZilQMJ+CsV5C5hrokx0Z3EawvKhun5FI
i6yyEO3SrYRxBm1woA+sSN1GKx09MUFhJdhb2Kdpbtzbn70ooJDqEquKfDklxNQG
4G9tHTuGjWg0+ScMwbXf/lH8TV2PNYz5uXnaCmo2Q03YKLQa3UidgpE9NbtSkUbA
vUJWm8cyvtTHqimV4NiKbkrqWw5koKWF3zxlx1kZF2GzEuV/LrbOXPeOvEMbkwKw
ZoLR9pxKOiVec7fenwIgxWdfA3FrkIoDXYFrRAdFtyOL8cLVSVAIBBHEiJ73yDSe
SjuwEwyiu/Q2x6LehPoM7Bz2gDjTrQ2biSQ9Yw4rSsPpwj10JayqWn5E1ybaWrTi
0WOMa8/Jn853pvYGww6blRr+MAHEeDTcgMgzSvtqG61rPu78wWpu1mYQofMifyYB
vnHH/EIZGUhXJZamJACUgFmXEmTtZNh4LeK93VUGtaQbJZWu5bkB6G07uUqT4dKH
5o+psF+kCroJQbHiN8NFi7a00XjuirM8TEQxyYsghFCupjYYmIa2IroA+xm85I1r
qSRODfDznEToNfMWu+xShYyXPWchmmCG6MDvcBJ5DxsyPsJ0xieqJj5su0vLIMeT
WLtO6T6AChgiU82M7ixDGRL5dWLHLrL1FCO/nppNeccAwfXI2CNv5eedegQsHjV0
m7RbZhJd1InGpgmtUIf+K3FXhC9GwbaEQtkiVCz8u9XvFL9UW9fMnzExsAWnYnWm
4TvV4RPx4NP77U18ph8UmNBjIWQY/dWluL082VdJzRTNJQWVWOJZviJQp0ShGS/B
eyilmknGtGPqP0AEAkRZMBqQg7ENmJze420Ol2IgF7i3WtCZSkoXD9Rc7kL8L5kt
xhxy+8vgPEF93yH/PDp1vmOCb2ETGhnfjy+PROB4SlA/f3aUrLFvuBe2f5IOhjWp
boLlmvf1ig53rd0oQgvnZk5wmzpjqIwb54rlmKKAB4rehaz+jsA2+XAcCPFsFh6N
F0msw0dc8NyI7j7J8Y7Jzd5G9WkgoUo4sDgLheBUEFh4fQpPJ2hSACQjRu8sEfeJ
gJtKfVQgYnksbUE9TeLKkGM2EzsdBv6Z7Cn11TK6EIziJz+KCejbU6S8w2YfKdEe
x1OxyclWox/4oschBEu1iyDCLoCGLKOjApGO0U//UK1ymO/lC3WEHoL7RgYg0J2v
bM9apMjyhjrutyYxS9kfh0bIZhQD5WTl/RQS+lb/4PsfTfI4D0vsLvaKNpCqCPNZ
inP7IF43jKi3pKgh7PzmqOLvyyyjB9H8W2CQxC4vzfI8zxiJjH/4CEd/EE6ammfC
kxU1uEcDWaXghaLOovrDwKVdOIUe0TWnwigwfWPhbwTOHCcgPvzGKwLRWwvkod9S
PXNC/tXtfU0VXHBsOBp2104mPVJP+hqPOjFw5L+JS8NjlAE8y+FqqQelgFzeuELi
LsdGu1VQrwlVCTcDdkrNQvD3KRvYe+VWO0rPr5gbUzs1mtoGTCxpX34tQ3nRKvat
LQrmAGXParIcCls/Zy5gdFcvk1wsa+oXcpGRJbfjYfHEgX0HaEEjmwEhz77Y50KW
VhBopcJbh/YY1/2K4hL+m+EWxWSMzmBKuiZUTi9Djm1JqsWhDotrybq3zI5k1NkT
w25OYzNx+bL3cJGLfhMqnVLyX6sPVw+Ery2Houzv9e5Ir+HkNsDGr4oO8qL57Zlf
WEZmNbmsaSmIAqdGfp0V81v8ow5OIp+gUXKXBbpNeejMEqHgwI43Pqu8yNfJDdZm
aDUqsur9XuwTvjmeASNgVx4alEyNxmkPMdtzyg/yhGBvHGe7tsfhaRRhyDuWd/6R
tuDW0NQMGmYzr80cUk9Y+/46533dJpKyJ2UKfvfNN7jASPuWnKOnOrcBU5OL1lJt
oSFYOp0IwriKwLf/tGKer9+m7kx1PPaUmjgb47L8FzQWmb9Jqi7OeivIzNr5uSPk
YZ335AwMFQhBFib9dhi/ZoX+GRjdHASn8QanAm2rP7XqP56/G0bP2+ByHEznBzNZ
HpXUV5+ZIuGtbtmjU+fVaqLU85ryDrcWXVFiJHeO+g+VCNFcrpfRYwJqch2w7VOS
ap1oCZLvM1ZdkChZ4k/ozG2GfP9TPw1cb3Stq9OMycI4tUeQ3nTmFbHsb6v5hu9V
zasNeBTgzgQOozYTz6wBqxKwzTcGY79kJmEUEw/SPycaSxddNfhrjRkEVCkHk1uG
qGdC/X/lM6vfjaWT83vbbF04YbUoBVIl2Svo3Rw1OoyWsJx1Ju1HxCZsBQKoo3k5
9aD7lb9xA9O99mrSdpzkENYzRQgqd3655WQ/b+3fPIscHHikJeuy5VQQOzszaDVx
Z7q0H1CZUIwdSohcfRVOluWScmANNabQ0kPNub/yZeCqL3H6MuCXhqeOzDvGmiNf
`pragma protect end_protected
