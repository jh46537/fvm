��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"�.0�у��u���D��@�� ��1���į�n� �n}�f�%�;>y�p�si(1���h��-�풀L�7�~������J���㭿Z��Y��\T�cj�Y,>�U�t��>~���$i*M�y�6q}�w�<t�]GZ{�%��e*n��T��T6ʂq�mo��(ްc���6��{Yv�5:�>�w]��_w�\å��+�9�R���%�L�2f&H὎��r ><C��=��d�H�$�m)X�~y���4�C�7T����QX�~�[RN[�Cա�q�(qļ,�n.�k��iQ���*�,�GEa�ʧ��,������3�(;�HH^��^嫖ٺ�\�=E� f-Os󮶊�{Τ>zt�Ը-���Tp�S�3�O����`�7J6�1N��]��̼�
̥8����Nu2̈�+�M�>( 3������t'�t����\���q?���a���<��������5��fc�wԆq�ua�Ҫ�r�eW[=��qy{����_�'��ڙ���^V$��^s��:d��mՄ6̨�͡F�`'wU1N|SdJ�Hܘl��h��ص�ާO8a����wI�Tn=S
a)6�0 W{��5�m�~��.��aͻ7�-MV� ����kR��%�:�Z��)?���c�I{��+�'�U�&�=sا��;Ato%GQ�5t��i~)���'����J���UՊ5S�h?<:ױ�"<r%��-�wl�dI��H��ӑ��Z�͉
���:��@��~�m���p/�I<���u��Q)��|�$�Oi�]Zn�A�u�x] 6�p�b6��y���)�BGG�eѩ�@3���z�e�M�Ln��R��2���-�D����(���߈a8�n�b󯝿�U0�b"�{�*Q��q���xPdӋp�����K#qqN�v�;��������V�$������|ßU�$�*���ZFV�#VQ�9$��0��kC~\t墸�9N_��`��V��'h+��7��	�^�/t�n��P�+\'�CF}��Ok4��������s~��PsȮ�:��
g�r7�1���5n�)�n��%ߒ��1�@��@���c]��R�ß1d����C3��G�q�[zF�`��N�<�/}5��K��O�3V��]����U�EF9G�ҍ�45�f�	c~�7[\|���p��Y"��^;G���C*��y�o���p�
��=�}QQU�@��~�<a����I��uD�x��S[�� Dt�lS�w#�*����k�4�W�������F�I$%�u�(���髛߮�a�l��R��J���Sr���#�O%���nS����
�-^�190������
�$�C>�*)s���&���P��T<xJF���J齺y�F��/7�%k��e�cO��MJ��d�qb�=��!�:���"΃�@�۞�Cc����KYo�r:�&�j���|�jMa�!��A�kU||������:�o�t$�Q������~�0�8���^
����)-,b��1. ?k�-h("ā���5�l��'|��Js��߂Z�7D	���!���X�}�b�7J�3%Bxu=����3���^@_bU��.��V!�]�f��V&�.Kq�zݖ�9D'�*
�Lܪ�@�osŇ�X��M��b���o�u�b�V�ƟB���QņƏ�
��I�Z���uS]J�d׎�?��A�M��0]K)X�����!`����:�[��p�qd�����XWt���M�@�:�����m�! ��]^M1���������'��H���o!�fe��ѡ�$}7�討�p��9�qBT w	:�,Ip�R���)����)����g���4�6���n'�=�`�g�h#��Zn��o:LÈ�-"w��H��c�_�=@�JR*G�:>&o�=���g��n"�N�7'lj��"_�,�*���?��@�~�J���oE�v�aӌ�d����`��PE��\�#9
�Q`���j�f�c����a7��Ì;�!�c��0]ٕ�e�X�'��Ѩ�:#CQƹSs{�Xl�s�Q�B\���g�U�R���j7�#�1�B�b�A��@/t�;*K�4K;�N���P���[����,6�$�&��f��%+�*F�����^f�U5Z3gƱ�����m�{��������<ȥ�uB]���"�� �e��aT��P3~SA�M�V>��*cU�F�T.��	'�����F<J��������p`
��"��c���wj^b��i���sǖ^X�h'	�Y*�n�Z�� �<n��wj�5n��˖��O�c^��TX1�6�q��p�F�r&�!�'�n�B���J��U9TD8��qz\�~�{k-�����O�$��Wx��c�����nr
S�Ex�h�s��5�0ɶv����#	��79��=yߐIf�4�����Zh}�0Kٶ|^����R'�n��z$�o�����Z��D��ۙ��������*XvϹ̳X�U�A\�����]�Ȑ���~�E��eP_�d."�R@puyN$����Q�eq���6��hx��R��Gd�U�T��l�d���=獈���|˳�R#>�n��q�rѦ]G���A��ןq�S !	.���/l�3�TT* ��~�]:[���*�*�,r�+-� :�����w�	N�ؑ���	�[P:MA�A�gr]�.6��%��0y�5�u�ܢ�9��B+r�C$��a�T�8��|o�$��"J1*l@8����2�	�c�M=�'�S;��r(��^6����';�0�d�S�Kv/N��N3Ar��K�l�W����"����b�{yV�F�kQ�%^j7�z���As�Ӳ��)R�W��^,�_�v�/3z�$�3a��L-eCS�;�����rP���"�xc�/o�\#L��S$�vP_�Y�P�o1(�G��C%�_h�@�T����g ^w��H���c�gʣ�i\pݥe��6��al`�|�4Z�v�D��+D=S	9<�m��ˮ�ep�i����W�8�����=��0*���������bE8^!^:�z��l�h��1uS�a���z�S��_PeGI�&\��}����䣅�N�T��M�8�|-��@Ihc�i��3^3M�gǱ�)���2�iA��"��`���
O�Z�<�����<2e>�B�|N���!;6�s+AY��t(��uUZJړ�m8n��2K�ka"KN�,��
�I�)���?+`�'w�o9�L�/�%ԁ��"����B�|]Ry��hs��J�>Z-�R�'FJt��Ӌ��N.ƅכa�$FO��M����/��zW�fW�I)�6
�X���*����y�m�U��<���@�W
�$K��ߨ��Y&	�H\3#cgLy�& ���>T>�4B}M���(�p�ic�;=Ŗ�5��T�n�wTD�R>i�����*����x���S Hӵ�v��=w���a�XY_��~u�)��@5��}����r <1����T���E���m����ծ!����Ɗ�]�f�����f�Rܙ+ӵ�Q���J�'@F��l�v���*]����	�$�a�'B&�]9��S
���X4�P��`�o�2-DKT)�1�����?E��YH�y��p�\�О��L7#	{�mh��N2~��m��o8�����" �O��8�<�K[p��=ۨ���o$��@Z	D���A�L<�2(���݁�����g�G�� ���L�����!v�����,�`�[u�y�\媯O����y�BW1b��q�~�S6W>A��C�z�vu���+C�Twe�ޭ5Bw���7�6C+�?46��=%NvO�#�&$dݟ����;6~��R��I�տ#������W[�S�䧥�Y�7��zBA�n*3(�f#a��{<�O0��qw}"q�$Qֶ�c�H��H�m�c����9qB�3������j��h�w��Xh!Ķ��ηu�˺�
4cZt1Ey���T/��LÞm��D2J�ߢ�j����
v/�F�������3Ԓ=B�(�(s�7ʈ��#�e�L��LV���m(�
��,H�S.ϥ��wA��4!�Q�k!�ﮨ^�N�N�k�s���e-�-;�y�ӯa�L@�?�EF%��I�5&ЁΧ�� Ϡh���;O�Po��V�kqV:h�m8��P�)�0��L�d�
�
�t����
�.�l�J�X�ޤ'P
љ��(��-���#2�V<Lq�*cP
�3\nlMί���'@��{ą��+��/z-{5~������/���r��$α�t�j�*�~��� �>
а��o�D�>���8�[i�	7���|%+M~*�f�x��2U�a4��I��HrTFU�*"m��:��uH������.U91Ņ4:S���?`��q��2]؆lͧPm�(�9�`�8ʿ�}�hC�k��x,�����<�W,����襷՘0���O-�R*w#��W�j'F��)��u�Xy���\��+L��&�}�b- F�YߢA�\� J��_ecƩ���q������669���H��9���m���d)�%gee*��5#�84�2�~w��=Q}��|��N���(�l��}�� y�(�B-8tO �z��؎^�@!�QDx��R�u֩!|�����H452�"�N!��;�z��
��Wф\[o?"�x���k��[DP�P�SF�0Y]>_t���e��!B3L�܆��u?�#W�J=L񈝾\��Rv
kf���\������32��O.譈��rجiX�p�~�/hV3;7����H�=S�i�)l���C�nxf�u��g�X�8u����R��=+=Qw|q��<5��J���*���;��38����:��|a��9דŖ���*���O�B&1ͳ.5&]')=�˚P&m%��c�t1R�@(�u�������P��sXk�<�ė���Y^f�:h�8爓y��$
D7�l��7���rT^Pxc�靸c\��`ҽ{���-��`�v+!
�	|eSש2[��ҫ��\y��~�'o<�
,7�b�xy.;���s��'Z��	^��<�k��ֿ��+Ht�I<�ӓ��i��8��=D�#w_��rT��A}�W��F�
����!_! (�'�ö7F���" �e���nӫ��c)vv�X�L��Z0r�ȄJ#���磪�Wr+�}c�
?�_��oŞIN<2�AR���mn��m���8#��w�����l����ϱ,�{)���M�Q�\�P�Q����7M�ٍvY�����ʉT�t���l�):�w��i1�doiϲ�B�����Td#y_#�&&�N\;ߌy}%��)���F��?¢k���x�J �ah�P�����T#�HX�f��b)ޅ~���5\G2�(��ޢ��|c�������TTt�7y��/�u�e���_�������>""cv�Ji�д���=U�fL�j[�R$����Z�$tGH0^:@iA�c�y�y����7�s�3^����f1*��#}р`\'+�#�ԥY6�$z�>G��?@�����:.Y�*yE[�s1"������ZZVu��ǃ�Rn	��Nh 9��&&��]@�97NL,����o��.��}�O"H<�LK�r�jr����.��(�z::�cb��g�Ϥ���}P����E�@��.�*d����pmw��_��7��8�4�&WX���f��ۨe��i��|��Z8W0Z]M8�h�Vx�HD;?I�x��߽WړOO��"X��V�<
�]�IJopr3d�Gj��*��R.܅��2��v-wo���y���סs��0��f��ǰ�r����t��������["p83U-n�x}�P!U���i_���c��oG��?��W٩JMח��W�"��,!�v�R9[Jh��s���n#h�	"=�[����N�bh�E���^	���|��c��?%��ƍJ�$vq�`4�IڳL���|��ś���.]v���$@��>�WƄ�bd��уa'�s��a�UJ�e'��T������5�N���}GͺW;ٗf�f$�-���!G��-vM3<w������_D���g�FA-J��X9��$ԗL�I�6|��zwE{���,)q��B�g�bΙ���R����M~F4HA� t:=�c�;�?)�[�DҒHj����|�������so�Tϟ�)���g�r{J��C��s�ׂ�g�N�2[ir�8VIO�.�&���|�즜��BޗiM�������þ�)�jL��[l_
!%�0�sxԀ!�C;�':����$#�7�a���8Zi�8�G.�d�Aao#��ohX��&�;�YC<��읧�{�4�YNhD�Zfؒ&BZd�=;��j�`4�M�`������5Q�Q�|cb"y�����M�n�G��b��	�u�-}��1��8Y�Iʝ���]����#o>��ٗ�HV���_�݂�Fm�פ��oT���
��2���O=R�A�
:�m��C$)�c~IF�$[fFV�����$,��u����GTہ߷��uT�_�8�\�
����$�`����*�����e�ԭ`�1<4�V��'��A���
ms���Q�B�3i���q��|��Q���	��� ��ph�EF>�G�3X� ƿ�����E�{p�8#���?!Q�7����p���]�� �gKzԺ�].��9�_O���itwJ�V��a��(86�K��M4�i|�Z���ۗN�_zq.��i�dR[�Ȧxr-D����VZ.�	3���Wnb$��/?����;���!k�k�~��ή����O�OG��w��s
W��/�P\�l�_�mu��>�T7�z�G�\�u��Y�rE�
l+1F���.��8:"Tٗ�Yvqo�bz�ۣ���t0̀�g�])�J�r����b�R�%���{�K@�v�v� �m�S� �xH���n�ǐ\.-��##� ��A���>^�֙��%6DE�T�bb�1K^ד���w=ؓI