��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{Ns�ȭ��+{do�;��F�0�Sa�K!�f� b�|oݓ�_��\:�7�'&�6V��mU+��S!ڱ@F��40�ї&�`]/"�c�'��&�e�Q&��b袔��@#Uׄ��Qui���O�?�����S~��~����������_$"L_]b��¯����{�j��`t�ez���h�z-
��>�u~N�~�,�uR	x�
*I��ӠHQ(��\d�#^�*dw�*��(��B;!cBh.ei�"p^��؇6</��Q��r1LQ0�
�kl��������� ��Ip`k���L(�QJ�؞��Um�%.z���z6 ���⏲Xǂ�^˿�qB5/�Q�]�J�4�[=��,ZU�^�u~����qņ��Ѫ��,%{oJ���fcg������>��TK�ʌ��Qf2���J�$��$����Z���Q�����9~�I?������oF=C+�(�(���t�9�D+��#����O�҇p�;�eqȅ�.�'�O��p_���,����m��H
P���Wd��;��[g����*n/������BT��ֱ��.�Z����;^���")��c����n�1�RӁ2k�fץ�,�%��3�'�M�P�Z�pe�'C�9E��o6;�-	�.�~�̀�~�R\�5�5�����`�I��x����d4�\���1�P�c��V0~�B�uN�7q���_N�F��zj��tP�f�� ר/0�����z��O��	?%��>��(���؄Wv0�~�/�h.MWT�D-j\Zp��>@��w�7����ʐC:�v�!���!V��]�%2_�@�*�S�Ud�sKV9&����Ř��#�n�1|��zU�3�!Y�*wW����	5�~P7�Uspi�w�y`�9"W����kپ��ɐ����蘎D���K�>�MZ�X^��!ӟA�n�4��ˉ,�+�9���"4���,~+�m�+Y!<T��]螕��ǘ�U�خz ?�m�����s���ʙE.;��\��mnTl�6��ꋋ��䃫�NA�����v{Q0d�HX���������r��>��M[O���N9a0P	d�Ȉ���.��4X�$�H� �R}͓^���|�t�*@���'��g�M��͢+��(n ��G�r�eBB2��2%���ݿ����XkJ��B>��"�ES9u�U�:����C��:߽s�r��42��]T�9��].m<7������-��	�K���^ ���Q=�2Ӓ�祿$5ޯ�U�効��?Ǡ��C�.|�8��l��(`�v�6����N_-)�y8��h
�T!A�*��Y�v}����i��(fo WBo�/��P�H�=�C�R
�����.��.�i��M�]�|��9�v�_�p��g} H����o[��^ )�z
I�9d������	Dݾy���K�:��ǟ-hzA괾}L�tX��#�u}��e5���7����="P;���E.��(�rZg���p>�'�?:R*�� �S�||�,�q���e�c]"'�09����s7V*!b�A|��;T,��Gi�=4���W X� �x�ۺ��VR}T��8��[o���)蟉��egM���f���ߗ~]��Q~�=珶��*&K,(� Q���T�9t�)J���4y�� ��vPҙ��ݜ�	�q�B[�H��s?7L�yOb���{�֔f��"�R��{L<�v2���A�5Ç������V?u�=C�D"��T�dݺ?�| �ݗ�"�D:,�e�+]�
�sGo"�Jz����f�>�E�������.�2k%&;G���'���6h	��1�%ʴ�O�{��D��qW.R�i���9�v�Y~4�F���J_2 ���+�L�}��P�F��@v	v"Yc��� ��qr�\�3x�@�;ww_��8p�.Z��VY�^Ru�7t��/x����$pe9)���iv�,�n�����vi���ޘ�-����~�n!�+]����U3e1��<t)T&|�c���VCY��MN�����]5���5S���tP'-R�_���AU/�o��g��I�y(h#�pl
o���A@��� X���x�#0�j`�zz�=���k�s��l~�Jlk	Pe���A����1�*<�'41��wGs�>�k/��K��t�iS܍��R�lw������h�")O�:�Y��{�9�4��5�z�.ces�i:�dş.��IJ�|VIflp9��g A������\�$3	M�d���P}$�I�\��C�w4��<�����J�r
�z�Y�s7�:bu�Z�qn���y��Y���r���4�>n��X����I�f�D��;ֈ������R�~^kފ�4[=h������g���9�U��X�;�g��1{�G��t�Q���ʲ��-W7�7��'���[����F������?�џ$O�R �s<�h�8��4��O��$�K~����:��3����l�<ǡraA>}�IوVf�,��߅
�n�N��֙���ig�`='%�T��`��P<��ٓ�k���S!/�?-iA�R�3v��4�1��Kx�)Ip�ь2�P��I���+=����*�Uq�S}�Ď׶�'4�a�n�g�ti�d낇wT�WB��&>K�v���#��QB	�?���aƷ@%'�A`�~XS}��t\�>�R	�	��U�G����T��"�S7'�S|攬�'4���uƤS8ysn3���(�\�Q�Xh�r�p}T-n��