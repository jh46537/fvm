// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:19 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kg85J9hN5p0GDTp7Zg0UYPJfFkeE3eeSjU4AgmVkMwqpI3YafxC1mt/x5M+cP2tH
7xQB0OP0ClSCFCZIMzG0hE9JrA5x3T0pCn0VoIZErkWwG82+bGf3LXP0PBi0hFiC
OJ5HdtFeb3rbxrVC9KZsG9efGK2ZAvQxWoDalsehKyU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
h12lCf3Qsd08pnXkP68szAkTf2CJCo4OdR7jDiLo8i3GszaHx9HfdfdGJLiTg3YP
eZDG+JmFx50/LL3Bv7n3xDBuSIcRuP5b+XdCODUmvLARMHzpReIlGS6++fYWTX5D
eayGeqqkYrFjXYfxYeabZ9Ld3GskeXFPsQ0GI9iIlZP6gME+IpcyEKQgIMzcVhTG
0N2fZSRsJoZJgApImC9mxVpyn0mpOLRvxkqd4WyXS/uPEp2yu5oAbTapF9vkghHi
nK/kR8g/eHC63bE0IgmkHdjCAQpOY6p38bqMd3JMQCtX/cUruTkfG6K2NUrS3w1b
/uy18s7fGhtFtBUPJtbtN199jVYaC931NMQdFU9DO7R2Gdlv5H0tJBYFvwEKnl4w
mmorKIDpfmSitIjG2QZVqeQXEkwraZkhi6fVrGxZRorOS82SuHhwlWOZ1ZL26aJY
ZLiqBiJMLO26XXZXsr6YREcjEZiqaKbtbzmMdN3rfxxZ67CNepz696ZwZbRRAZsx
QuFAFH3eacC3SILGwdbhz97cwpivJFYlJA9rds043b25Kr02Y0pNdxI7zgUshgBY
rDGPTN1qrDT6qWNwf9c0bGL0em0pdWSSYYwTmQFTqKuW8YMEb8cCKZYmvOk6og4A
/AyybEtjP/4WM77Wc2SdEnjI5N+Ad5jaraS3C/DcLMpvzvPB9htLAYQMlychsJ24
SCjUNWkL15CET1PMbvSpR8OXlSpOewk2bo5WpPYtwxuz4cTPre1g6UZTzYTk4QlQ
qiA/PcvrRbcHnMrPH3lwpdDYuTlswOriFUhDcvyEkjEzDQ3MbLlGbtRnQgoTyces
Dzz2v1hkGAFkALImSetKbPGAh/oarry90wHwItkmDEMw+EhI3LoMuRPdgzcLKbhp
SMpAuHxRQQ7qdD113JGFi0+V64l91RuZPvXPtkZ1+w1Uyqna1NzTh+GGA9ctt000
MxD1peyU8ICndtNv7efRjTS3HBUcGUZLaRi6Nszc8rA+wtOWJsryiMjD9qy7noue
hVLc3y1FItAx8I/BVuwg8oz5uJ4Pcii9nXicNREQSmVkdICvo5IK2DHDk4WKGshr
W+GBoalz7mrkyib7FhdTHOgscYlT3+C/TuQSOSVHZXGBxtioLfXfEi0mqNP2PBli
/VBBMdxCZR79y5XP4ULeTnm3YhISnZtqkuIrx8YvR8X31GOxm/zxzg3kObVPs06I
DwbhiE17cj0CAIQU27goBAANN6Yxdi/c+GgaTzlQYnkY6azKPsPHUbp8LGU0EsTv
l+o58qmHokKEbQPc4kZEy9JI5ZkH60bd0WJ/YIoF9T3iOiYNLhBceb/Im3As9U8D
KMw8NC8rmgyJNpJn4K0eQDeRtSbwGGOXugxlkcD4LHEFq30Y8J+yi29E8FVOM6hu
xwUTQTGIMZSM7++wEKPqDUxKQL7Sy5k6giVBv314aXwhXoE40fjWp+49od/mBgHE
1wXd88RHM/HmXrE+tKkGb5FjpiGjm2LKScR06mA2i3VMaI6GIjifXZ9CWxQSREVD
cVitwdC94rnfS5l9IpCFRIFszK+WI7JY2X1hENAX2P1W0B1Yye9HzGE6laRV5yRw
Xa42rS6TSlsgDVxklZMbOHrobdndbDLfdfIuAWIfDYo2D8ETr1rFh431Tf+H5btb
Poo120LcD5ZR5n9fUzbcrp7DgzwEgcThMWDbnjyYpXEUoQRLEkrAdTcd+dBRcPMd
NbIJoBuLfibAz+hBXL6c6SjXWKfaj1GfdK/vpa35n5MvtwAoSyx/x2eaQiTJT48Q
sdtnuEY7Q7EDtl//T6kHMcub2DrM+hyb1kC907c0E3fMDoUTtULZJdfErObSzJ2S
Bwva3kxG07vSpkk1giWrr5WlTkTC1njKBMs8Yb/2cVDCCchlddY3E8CyatTOKxIX
k4Yp0a9v+B9c1raxohW/jGu7QMXLths5BWoOZyZha8pwljYsg93h8QqyFOlj8VQ0
P8nttK551kt8uBzMuIgowg6bFkthwm8ANvtrYqYfkVUyaQaMEi+W494Kgnsuuj7b
HpLjLK8Lcmq0k250RyFtD232i7ZT/sIuzulKKa38yX8TWqbAZxQ791aUN4Dz4qYH
TPSxIKJwI/NmMKwgTe2ib+pU8Bq1r6/AUqlWLI04kpDhyJQIyp47vIdTqbf4Ma+r
WeMvetA1xCv3BvtcDIScV6TZgGk0A/638B9JgeJe6sbvcoG1CHnr8mDo+cVsCJ7l
V1qaICS7KvpAGJ4PkrjD0jPKlv5sJGmI9MU9Psgg9718aUh0uey0MR+OpM4yX4Ky
lOfBWLGmHDVbmhNp6AjLYnNVl30+Fh1uy9yWTHHNSnjgQDXR7KXTMROcOSyIDTT9
uez0e/VbfIQoMfm1HnaVnMiV07Qa0ytQlcY8vA6puDEIekpaBPQLJi4k53LcNow7
npu/ZubbY16Q6nuXNBssA07vYRd6OyEgutj4SUNJq1SOXMEFGXRLfw+SrwjVZBh+
luvSWF23+NFPbcHD9c3tSya3xqRtV4IcgT0R53+sJtWQOAnYbtvdQNMvIzJ7mO1O
0e258esXKbEgP/C1+CBjSSpHqwTkF9+AH5l6+9oQDwZJqndIxVWTtWzzUKB8s+Tb
DUKTSpG27eP2Eo9zvrNNZmhywIOyUiEaC8s+exIv9mGIfqqfRsYYY0An9UKGzaVQ
IdOSnUy0yYHZ/qqeInllTksKN00PDpNHA+W4zGmRna3M+Sq9oKG66FbfAoGsHbGp
stciWbok4bIqCQQt3qSrUJPota/ynwgKGCEvKJPvHUCcUGArhtUVPYLKxhkF3I0r
wXtuqDe8uWm2+Jp7KINbEaJmBmtLi8nlluBqmYkv+zQ1krlAsugYJmEfHwZtlT7X
84KnfU6e7f7NqKpHllgBni5GQSkO5fqVlTAXUiN7af9c3GRypZxmkMRbYPsaUIOF
QMwZEB4dxlIRTocd+cXL6lezbd8hc4qS8vZRarpD1N+FrLJp2r0xtx6iZLUCfPva
AeG6m74QflcTPU6Turtt7rA3cu9pOIjIztie5rz6cUJPHSW6PWSa3+ubIUiAVMv/
x9gEAaCRfyj+mIQ+rSxNdJiGccZ+o2Ogw64Cfz5KOBpU/tduuipDRFYb4gd5cUos
cxYeTER0+snbovPMKXS9/JLl4ZniUgNmPUOxcmcUinbDtBegrD0kuUv45dK48XQe
PTbRIlfk9go1aYZil58t9x+cIIU6SgY76B9o9zuj/cMKxCvk0VqnWBCxn6qD9xo7
j05MKQOXY/OQ/JC12Ercmt3Wj+q7mtzLfLmDUZVPmNXTNIu8wgDJzFOC4kz0lRVN
lwBzFn/aVG+wUyKSy8U3EOX0Cexcg8cYjxsY94pPLVR3WsQYr+k7ta2VH+ap0JcF
gnY1UI/ZndZ3jtnBP5Yk4qZareFz40n5Iu9Nfx4GXLLgyu50gvoY4h/Ro1l2rcNu
yt7MAD3TU7t9UtMRFfEguayagMNYBEqJIKoxqiAUoMPmrNVaoHa5fR1/YJmvXAgV
cj7ZmZniDmUzC7EgePtMX5XLDu3cTA42fpqNQT/q6TlB/and3uFllceh7jc8UBch
+utujD3kgK0qaLMwOrzlr7ctPAA14NzVOw2+Y8qay9xDV5noty26vTzGzxiPXQ8T
J4ApnZQukzZtqNhTMkR9kWLfTvInFa2d8wq160Gs9xtz2gcCgO+tZxLJVAHlhDb9
I02C7aSslI7FNNBxsz/oWb6iRyAJPcDJME7+Toomk6HNT+Mm2nnxMfjoImGA+CSj
rkLl7+0bfQi0rMQOvwIo/WPY7ZixzyduPXV++1IZEuZtr5SCIQNo03jEURv8tWtS
imfPTMkyU2MEdu4x/pNs3GY84BkNvQviVYNH5vxJfJTmsKHrmuoC64vnthUYtqXW
KXWIJh4U6dV8XF2uNYhViPr5YX8ujNDdpbOldGE5y44d5G7K9H6uAY7VwrTQ4Y7r
uMRfzvGyACBGIFDIsJM+E2bL5UgE7/JFeqHx1u6jDoK+bmOjxUZFifalxC0Za3Ko
sA5BrAh5cDvBTtwA2nAyGvPHNstm41QiEZD/IhW+uYH/FXsgWu6sjXOdDS8WxDgb
1ooyNSXfuVauHnB3TAeFIgquzf0Xtt811rxFVPcWehmwULwmK6PZnGPo5l7mNvF7
wyfgjfq84bqdpZRApmd9zRikv9pdxSBL8h0fPVOeG5i2mn27fJepruyDlOJ4OzIJ
wHtQ+ONtBHZK9G+RaG3sCpbq6M8LCAjlWl1VDBfQ45O53L9Xs8gn5R+KL4qKj3f5
2fl6P+tRd7ICeIMbXx1VZrHvXheV6pkcL0GZs62Hb6r5knLcf+UT9irXLVhXpsff
r+WEL2Qm32UChzskqxWwq/QFu2oGx5IPfjeU9tFe9/PvU3k7yjQmdcMM+B7cMPKJ
8SwtdZwexSUJy0JvPP3dPDc4wlyUSGzXnqWNrTIDbg+0dAWiqG78yJ1tYdXlR4C+
4XjSiVbXYxeZmJNDElr6/ix8ziRx4sT+Er3HiNbNWQqXhd27o3Dzc8sOluT0NwzR
c0+gdu5KwgkseHdLr/CDUq9JGd8WqcTaA0eEVL2k1Zq0F6QPab6rwEe2RcrxLktp
+/HwuK9EN20Siuqb7NtfxuHovlO/rFfiEd4Cgt7TYCUKYNg8p7pgAjHG31sAEYmH
x2y70aYKlMLUFHRletKb+sRi0oBjRnMOi+GGGGagTA3VrdpUORkmKwD8Trvp5pNX
0kapk+mRj54fxfStaQktPgA0ICptwPoLp/K/qZcxVI5Y8e0wJ691CDMl84avWgmz
8pKHEfoZROFeDBTKaTX4fzBi5ezPLDi0SQ+M6N+1JS6487MEw+DeXZVwBsQtEr7R
5Fb+KKjjIrVlU59H2cygeOApH+6U/X9oYtZeH885AFVbeYv0pnof9/ZBMRtmoioU
41CGU5W8AKJ6BckBs/akKk5v9dQxqbQtzWZOKCqzXbSQIEOmJCNsqldK7wF0LOEB
12a8N1z6V4ZKbdbqAELl/DS6jnWh0klwm1IYTwA8/FjK5vYNsndItUcyWrHbYBGD
61TkSV2B/0mjlznmKcM01Cw8npP0B1T5tyqUWDHu5voAkdUreSO+pi2jg8q2QAdN
sD0wV4cnAfFfWyWkfPA6rZGJ4k6HSgEmIL5b/ZV29vQTQgPAOGt4emKgJNe2mizg
rF03w+zwV/eBZNiMlBEmNYxMZ7OnE0Hpge6OxKFqFPRMLl4klzrieEVTU+UjZJbd
xa+y2T+xoz9MjGXrvgr5rkcaceFs0wPT00h8v5oFXiJ2CH5eZjHBiA2wslMemGBR
D2er0jnbTr/hbJTovzkEAiVGZ2btLZvEXzHGIIRgfZuWE3jtnUoQlPqc5OBRX2VY
z6E+lK5RIVm2WWKjCcdlf0WP8v+XgTd2/bHveL5oC+Je+tfCJAGhYgvDM6zXftvJ
GRgbSuk5KH+OwcWxogk7rB0pLWslEB2ZvrtGrQsID0zJXc6haUfTDM/XX2kwAbun
SvIqe/AJoqLVCLlP+0cE9LLlYp/GeM7O8JLLALj8uE515RPXlQrI55/mBwL+KQ7U
c7fPm0InzW2VUEFVn9R+wh5dtXMj4HQwL9C59VXfEAlU3QMlNIcpQ2LFXh+PQwNQ
xX9hi+ESA0TH8S8io+7C8rzUpA0ZKlkhEivNilVVcXYN6XXM5aMExF/eOl7OeS4F
qbuJ6Y7vbVc0NLu5JvX7oChj2GbnNRtAdzEGCoZRgo1K38CRZLkkjjPsepW8RW15
PjV2FIq45ke7sB/9smtul498D60184361HvFZ5Kj1JF1AqeIJIESMNsESma5at1H
NMh4LgU2xp09H4SK7ZhYz2TxL23LiBCKZ9E2VA2rLsN97y2vyCh91Sm9Z4zicrsY
kzkeSD67Ys+QA9i4pROsO+xSZGTnmHg5xnDhuNEUJGsTV9YB5MI8RTL2grAXRRVv
eV8HvpFdnb/G38H2KaJxaee/n3qdqPrD+z45xuSS5XC3R2iFeBlRfJmEWmWMDwwi
9sf78Vv0Ez99QvKrgvlrwpkB77RRCzeDF/FXjGPmK9jQ7BZZeKgqBv6KhrGRdHYD
ziulfzgBn81qN805keEr2np0bOf40K939RKSmPPtyl12FBkO3Lrn827PqJRhX6jW
zaaBAXRuFdGNBTkguNV+t1pBpqiMqSeV8gY0Y0XeLExCA38E+t7t2tsq85FhKwLI
3BYgbdr0vG6utgukPfYcmaqBDCPNJy20jufureeuvTi8SlE4L1dmz3VVo0xuPhgG
mp/+buNYmIYvGQPsZqOW5R7wJ1ETelTC95JeYoh7wF2deibgS9XO4Sce7a3htwAr
Z/KWTcDGmUoyU77ePXfs3u7GwwPYJkJsJxA3fTytn2jRD2rRPqD5JlQ9IXyJjzF7
T4qPnISQ8c5BZGbCu5XpoaQ2KoR0OPqwPRm/EU0SljRN2wo7lB+mgESVl8BYO0ho
1qevsE4+tXxzDuppKqqW/Gnx48SGWWfBA4W2tFWKLMLvGOPwuAWV5AzERWcEc0zF
u/4YjNH1FDB0isA+hBzADXWuacKQyywSSZKKrL32OPHwjchgujU8OvwCYA4B0iTk
sKttvwzYsYbR/ghHL3lL9xKlAq/GRFmW1qsxMkiR3Tqh+A8931IjvaCFbwjkGRku
Cq3BV9V2SYaLvkYAEGeceRrILMSCMfoUK5AZsSKQ7eDr8AKCDS0aOXcdLyA0SO5a
XW4QqEwnaIAIqbhoRxZfZdBvdwCI8/btVrtQHyNh4VpMzvBcFKFPoXoKgNhj61gk
XjN6kYF2Y/RZpbABiih7OEc7qaGQlfH9aKBrWy+3UEphZrVPbTPf7idiKkQvhuBr
THgVXxdVRdylibAyaYmQ5HEcxjnK0x1MTa0akTqshZTLZ0++k7skQ5+pOvJKw/z2
Qgh4IJr5rKamj6en/ptOXNri50IOzDyXKvJyZg+7gkuvBsfQRLVhBwKJvdlLhCKD
XMRlDNNCPGZxvlG6lqYZvnA2rh83chTFT6vYTrmYwyDmq8oRqlXxXT36N/3sPJeP
9uS4XkHxLyQq1KGG14Mkf6RJc8QIHSdMhMO8p7TxykYfPyX75iGJ4QyloOw3rJAX
BFBNt1WRVc162pLbj9Gx33wFxXqjQZWX8521BAeRe6+vrpU644lIcvFCvAYeaMJq
1WIQWkiCfPLmrfcZ5UkUwM2HGIiMM1qy4LlPObcY2ZeSdj+oLXVW7IV+GbzlEXRi
Zg6qRpQSHKsPuMpr0iCiddA4/EQNNRbUPkkLmXS0fU0Bxh1QtQJJgs2/Yi6/b/NH
nIvXGSWpifCqvkKO+rvuocSD+0fYE/7JNMFk2JAn3P266ImbcyjeUu43GNiRfnUj
syHxbtgCRjNhRAhTnSJ7Xzr2CRNsS4Gxjng2X/nec158H1LmyXsDmdNQL0eWLq1t
qnmQGoIKDQAcM0DJQJuTI+0mtOFY3KZaOctrxyak4R5DrqiCwt9T/BepHB5eHE5Q
qjxrd8XpbOaMfMDNBPCjSgtBQjFTaefCwg2DDbj+4CDWc+1/szIBrNkoNvbVF/Yi
QMkLYASN8mq+72Oqg2DY013paQR8ADJ/fp6+RpTl6PI=
`pragma protect end_protected
