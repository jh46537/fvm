��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�{8q�]�{T#�5~e ���J�	)��2Z��q�����������y�����M0஘vi_|�}�؜��3��Z6.l$c��-/j#(�\����v��C-�~��OKl�F�Y��z��	��# �E���YU���j֥��?�U��ɲ����v~h�,Fr���_�HX-0�HE��`�n��r����y9�jA0� �E')�Ҫgv['��'�A*��ے3�0�R>��\�u^ZD�
�١#FA(�k�q�'���S�8KVm%j���R|� ��SM�^�ȶ]zu�>��Cq�����w���ʨ����sy;]��5J:.���/B��N���.��y9Rִr`�[�〦��ZJ���gI��R	��{�[����(�q��몣{=��a�G�`����U`��V8�)��̗fC�L
�VF�G�[�D�o�+D��G!р�"o�q!cW�4�$��Z�	�^�~ۉ�39�B<G�*�n����ZZ��_�0=�D0�΁�yB��a��������g�מ�	��3�9a�![�,ʐ���=��7�@��20����S��;ҷmHRU�Ska~|(	��(8�AѼFn;0A�A�g	l��j�G�ys�=J�~F�P�
ҥ
h�=�'�B�z$�6y\Rg������%�8,�,,���D~�dz��[�#\��q4�2��Z<`�!����&y�w�.B��w=��op)��"��S���(���1��k�HcV�#��a!�HR�;�J��T]��&�c���A��_9��;2���/�H�/���|�%���w|a��.S�ݡ��nM����I��;��(���ۯ���m��7��2��aܨKr�P.��c^v�lB~/�7�Vh[�k�-�Xa441��D���i�TT+�}>v~`����Q���~� +��;���$'E6�i�r^��)P 2�N��q��p����7�6ily���_�Y�*�$�T,����k��_9���:��C�4��{wO�9��qeaz�b?9bXqr��a�3"���)o�*r&8�Bsc���[S�yۥ	601^c*N����K@J~"�a�}S���B_M(��8%��A"�����3O�l���B?���^(�k�FLU%��K	�t��>N��'��୯�V^��7��YlkH�\�-*?������Jٳn�A^�e\�s��������B��g�8�]�Bę���e5IF����� ���=.UB��K����0@�t�?e`�G呕/0�5�Y����;�|��z?�3������5th���T�A�8ݟ�lk���3y�CBZ���1BW�qppU����r��š�"]3N��Zio�l�R�N;}�6��pEV�n#PW�U(�÷�:!����]caͥ(Ӡ��?Z�p]�����\/Y�Ct��s%�dۦ���*� :�u$�&g�O�GLZ��f����`�p��5T� ����Qh־PG��F
�E�z�[R�)����?�P� ��N�(G[�
�r
�$��{�|
�D�)fR�L��joǿW�_��<�K�+���^��|�����T%F�x��yM�8=�Or�PY:�~�a��y�S��xF���͕܆����� -V�mZ���ټi3	��b@YZ�'���)��]+�wV
�^`��(�3yʄ�0x��#&R;� M�	�m m�٘�,}T�l>I��ی�3V(�w&o�=b�)�:UAUbȞ�n0�C���S��GT�?��<u{8�5���X>�.�*b�[w�fŐ�g^-R��n�[����Dt;y���< S�mQ�X���~~�/�ͼ�lA��3w�4�f�(Ȉ[�
K�!C/�ڥ�, An�Z��\F1[v��tU�o�����֬s��I8	=No_l��V��������w��ˎ��`�r<6[%I�� &�ރu�>�	qS�?ᶲEFs����D0�I0���aD��+~�,���(��5J�P��=���8�=ڍ.jO�IC��"e���
�2��|��qz|LJ���`�ԜuEȏ�?�7@���AIa�S���d�����6���F�2Bv�w->���o)� ����H���&�t
��nx�'+J�����WO�5C�ϸ���u��D�;�:����+�%��'2��aܪ�|��5ß��2��ئ�+�2e����K���,�C���%�oZ�T��X�ԣ9�a��q�u�~f#E �R?F�7	Q�8I}Wnm�N�k���7��ޠg��)��`��v�c�k�`�$6|��l��I��`D�78�/~p�u���+4��a���˛�Vy�(§����v��!����f�C<-:�ˊ��u��F�mF���/o��fu�0�ES��F##�Vnb̎@��b�A��e�.4B��),9����)G'�����6��u�'Z�4����Z5��.�Fۙ�
�e��-�:�fI���5�]�2Phw�&�М�Q!RWG��J�CX��R��2~l��a��������^U���i����!�ICIҲ)b\��<e��O��j��1?*�i :��'��/W������	`#q��8�C��F��I�a�G�����i:�Ī�������/��i��-�M:�ZyDZ���L~u"c|�4q`�0>a�Ϲ�@�M鉶*���G��"�����Ÿ�x%q�Kx�0OX�H~b\�RN�FM���&}�U�[�/�!����v�
�)R�Z��E�ҤM�0H��[�$l���5�k�h$��%D�Ey2b���R�İ�g�~�em���ES'S�r)��F��R��Ȟ"D�;1� ���4�X��H��T́0!C�J�]M���}��pS�5%�M�(�'5�y� �!lO�5�:h���t�ݽ뜳]�l�g7R�>�����}3�%��ݮn��i�} c�K5&��$����/խ����r-�ae!ƾr��Ka;S���EК�ӽ9�MaL�E�.��]wC�
Sm�w��1���#~���}.�Y���z�g���%N�DID���vz2�ɎKp�đ���HD�9���8�5D��2r ��K���N�iV��ޚ5�#�g��ȮZ����H�>��zw�C��v�U�>�t�-���� �$Ʌ$��˛�T���KBkK��)]��n��g��S��݇�L:�������ĶdOS��b���e)/ژ$69��q�����fc{;0���b3�d��7]zs��u��٭#���/ɷ[��J
* |J�i@~Z�_~A�F3Rn*��;�\���-O݈��b� Y@:Ҷԁs�܎�[;-��_`%����Dy/gu�T;*�8���x�o0�QT�f��>9X�ݜ"�Y֜f�ŉ���Z�b�5�J!7g��bw�Pp�V�Rat $*�rb?ܲ�Q9�.!Mb7}�O�	��N��Z�id�M��4$�/����gMg�qB�eW"'yg8�L�A[�#ƛK熃_
X��o�[�F��歺30��,��4�X4���lO{�(f��4���,��l��;B��ٔ��,xY;ʻ�T�v&�u�e5���=m��	"���	V���oZ�EKck���ub{�pu;6b
�-e�һo��*��\�s�;ax9���H�˜d��L�y4:����u��隷���n\�����\H83�����h[ .Xw�g!�&l����|4E�H�A-P�1�wr8֍阀k?>��X��yX.��Z��`=�e��ʚ%�M�RY\�ǼI(HT�ǅ���vY��s'MJ��@\9D�ЉZTK��Ď�v�*D���M�7N,�d�Ģ:��	�|�H�B[}����w�~QCPC�h�{�*Q�{�����J�<l�e��~�W��S�6��Z:&�҅noEa�< 4��s��:�nV�q�����^YO�Pִ��SSS�C��疺��O|10���h�-0�pl��C� �x��97B�v7]�Y ������ʇ)@���Q�R�����_�Do�f�2�>�� �� V��AMEe�q.��90n֑^f�G�g3�q�6�1��6ː�Q�F�r{u�G�'`�D5�J\k�\��3�X�L�}����s��?��[�ebt�р�4�/G��Pނ-t,#|:A��n�p�iƨWq�7��L�ӡ� �f>��&uB3)WC�5�-�w�	���N�DufOta��m�(��ڼV��e=��0OO@,�D�H��>T�e#�Ȯ6��&UffG���C6
�f�G��`e6=�K���f�I�wC	'�ֻWa���@l����CP�.4�c�{�`4{�;�f �rz���֢ΰ���_P��^��Ȃ�ꁵy������i6�9I^k�|�_��m���N�zfv4W-�'�J��"�U�D2��,�ܚ��9c'�W	�!^�'�,�H�)&#�j���9,:��pF\��)�o�a9D텀>u��*1�xⱄ����2VjA��!�Ofz|�+hL��:������8�;d�S'�7�K�{�up��{& "8�7�[R��t8�^K��]�KJ�X�S!#�[����{.�����D�_�m
z���q�a����H:�� *\�����i��{ �9"���X���H=rO��pG�#��\C�,��О���L#�U���Y����5`��q�:�=�� �1����|0�>3���p��"��g�,:������zΕ��z�������j<l���# ��Y�ۥ�WP�G�Dډ���o��Kf�ި�����\���['�Z@8O����G�
��sH�E�";M�a~���ʕ�G@��e����N���&(����@u�&˷簿�Ha��f��ٵk.� ���F�)�Q���
���|������͝#�)��@r��9PG(B�i�C�y�wpHK2x<��w�4�b|U���i^ZGb�V�������|�p��х�Й�$>�O\��m<�x�[v��o�ߕ�����'cI&)K��/��ִ��u�!4�: �X����5s�-J�G�b9����5�zy�J��}��2Jţ��������JAr�UJ�2�OlO?WY��T"Ws�v{]�n��� *X��� �ƽ3B��lj�7!p