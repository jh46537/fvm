��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�ds���=�FO�|uܬv^8�T�:�_F�ğ>b2˕@J��+���Qp}�ń�9�����k�ۖ&֬�%P��[-?�c�$qqc������2�'g2��Pέ�Ü� ��������S��=���>?2,ÝҁC:v�GQ4�b���{��U�8z�F�t���g$�C�ȶʇV�p��^�Q�=�ԡ�]�>z��*̿��j�@<����1Q8�2%M͓Ә/�윎�t4=�+�x����v��2�Z�k��`x%��Ϭ���ٚy3��>�B�d�C��-�3��]n|�d�;���O�ؒ�͍�x�sI��+��ռ�W��Lʉ㧅3z��	�O�}iNH�i�����=�"o���̠��yz'�u,� ����"��a��3Qμ��ʯ;c����^W�f�W��L�iAɵN0ŒB§~L� �������J�����*�ԬZd�,���P1�����5�4x�=�}�{���,kH��{�Q9�aDT+����`�%�Lin�P70U�v�@W�(��kC�<�.���F`����Sk�59s�����:��azB���Q�dK�����Y�E�JؾȎ�e]x�1�H}%;�I�"�Y�{[�u}r�W{*�Z�BQ�t0
&+��A`��Je���~������q���s����fZ���t�6�>�X[eK�Զ�Z�B���Ӽ��Y�칢��	��̭�m=xz��0H�ݢ[���2"t�S����t~�?�d�-���B,�� �l�r��tϿ�T�n��XP(����m��������m�o/b�Kۊ^|����!�}@���ZP���A���}�S��ЧA�49���-���,ʭ��P�-2�n�(~zF���]$;Jp���b�¥��5G(�F�Ѻ�BĘ�U���}(��`-W�����+W����rb�4��er����Y�����f�pg����S�{��ɨ�*{��JlK.���6_e��T[-��0�:g�٣m>r��W8�;���������6k/wNǭ�&E<�}^��+�7XK�ߩ��sqcb�IjSB)���3��)�����h xXYgR���
s�6���	�G�uq��/���"��}dv�\K�y"!C�}߸G�.�g�y�Q����댄�����}Qt`��6Rۭ������Q/�,H�N7��@�e\�
Y��u�<�����$�G������⛯
�5��v�?ee�~%�8bh���ؘ�a;&*^���9v�f�㼽<���7K�۫ag�Q�Y̬�紝!����"X=��8��J���J�Ra~�1Wmi�h���Ŝ�u�/�18~�2�G��z�-�j`KЩХ�3,Z=�����wf*�����z��S��<B+���o��20�j����t	�aگ�!"�%�R�is��%'GB�^�`�4�wO)�V(���P��E.�עT���r��\���rSWr��tj�-fz�v>��˸��#Oͻ�.W���������No��9�T��!��Y�\ ��m�a�~��b��u���Nӫ�̌o��R�pY*ps�~���]G��&g��L�ҁ�b��v��޳����Xn�\D��B�j?�e�7v���ns���*t	}���T%� �˹���ͩF""_�8���Xy"WK��Z����6��&M�fK�1T)�Bf�.t]���O܋�\J�� D�m�"���;V��?��w�xd(�Z@^<�!F ��{�� ԧ����f���(?��[}ъ"�`�k��1�QB���t����5؎�WKld'�5��p���}ͯ����ы&��^��H�9@����V�̪+���I�:�|�:���n��f�%N�,�r �*��g��b@��������ۯ�����fa�G]ÉQ���Y�诅�i��[<��w0������F�3z����?�뷴�ܝ��KP}c�;�Oo�t@�����#c_�/�|@�0/�e�:
Q^ 8��Bx�x�+܄T�9
8$��]�푴}`���&A�C�׶mV֒z̠�V�.{�DWW���A�ϭw�k��UV�|8�e�}��#�W��Q�p��f-hY	ʁ���5Κ=s���p���.^Zk�4n��4]��W$8'���;��|����u�f��߻�%�q��<��"�*zf*$yГU�"hA
���\������:,���Cp�>S�Cl��ِ7)cq|��,n����ʗ�?Z"��Q�1V��0?��J3��sS��)�S�%4Pg�z�l�(�û�ӿ{��<v��Ι���|��$��Q(��KDPC~&m������p��M#�G�����=�/�&e`�:ɮ�]�_��u���,�qa���L@��\թ�0�&�6�7[��������7w+���� N�X���if�]�r��xu���#��5�=��8M�W���QN����:s�tr0F��h�Q��%9��L�j�3����X�0��sO9s+ɰ�Z|�'�*�r�f��R���iEˑ��=�l����N��怾-W�őe�U��\N9R"]���@���1g+^**;/s��;u��?	�s���!�&��Y'�?C}m�s)�GR0 *�H6V�i'ɛc��b�9��Y)�yC^��#��yp����4��}�y���?@S~��$;D�2��Lw7�Zwx��9SѲ�r�S�bk��� ���!k�����'ҵ�J*+|!�Z�<.Y6�5p2||z��P��T2��H�Ӳ/�`������ކ�eȥs�O���嚐Bm�R>C���T�������d��l��5K68�cA/.S �}䦵��;��}(��ؔ{h�Xd>���93a��:���3�*n���m��0�^5
9���7��8�9Y&D��K{E�3�͝�J�FV �e-/�d���rT}��S�3�(��_j�����t��I&�#����&M�����2��`��h{����Lf���"����zH�^��i�x`��҇#܍�{¢/~��L`�ýI�j�݌Y��)�b|3P�(��`�}�/��r�p=���kd����@̒a���6�~�I�'l-$|�dq�Y�kZfS�E����V��i%��*�&;�G(�����x���l6�9Ձ����P�oD4W�\GAcv�KJbh.0~w�X]GA�κ�&����0M2m���Ț�Ƅ���ߪ�����rN0��]v�F�P�3�XI27$y6�������VO4�ĳ�fL
������Z1s�������[��Ӗ��L��]$/�D+����B�fF֡�9����9Q�1����,��PC�㏯]�tJ�bu�0�)?q�S�;���W��^OR�ݘ_�ӆ�Zظ2��D@=ҿ�d�^ʯ����g��y���V�uo]��^��p�p��@/-d���r_;�z|1�4�bPf�wU�K�۔�?�YLP�wε{�ڙ4%�C�9���Ƕ3�v
�ލ�Ȅ��"5u}�}��u!G6�O�g֟�������%��	����gK�������`h�҉��oZ�?ۗ#��r�a�p��4I�	����)�t�'�����m�D�#-8��¥71�M,���1_��`!&
]��2&حe6m1~zj=)�ܧ�2���B�O�j5�n����)�}"��sY�������Ka?��6�+��+SO6V��*���R��tF���ʚ¼��ȭ���}5��m�U��Y(��2�f��'��T��������}��L�}�Y�|�k��}6)����s@�z�Gd�ieBNVa_b/>(��: 4�+�g%Y���.�H�2�-o����z�u4p��U��	9l�)�*� ���Ly�N��}Ӈ��(���vv"bȬ2|�m5h�}�g���/�u[�#JՉH�E�.�
>�����U�S���Tޙ�Ъ��E�tw�0߀��=� ��$��
���lLE��e>��6�^Hj���d�����j�����dO�����I瓛2�/,L<�3�d&ܛQ�d�z>`[�@V�t�?Ɋ5�Cҳ����,�l'@���T�I��}��� Y����Q<-e`�gIp��&���W)����_�7�RJ�@��G����;�>2|@e�Iך���N���M\�z��*d�4����S�.�%�����s��c��g�ڱ���asYk/�v �`��p�D�Z��3��F��gǖ���ԚtS�5J(��� _2�U�s���a^�U�=����?��a_�!�=�nd2a�j����X���I:���W�����?k��k��u{5�ƛ���e�~�~���[�2<������:;���95����̬�Rx��<���}D$��8�u�銒[���
�b؅�C�Bڽ����y�Yޯ��1����G/�++�Zp�Jo�&�y�v�د��7��46���p��o�朽/{s�BOj)8�ls�Ӫx��~�L�m(����Yō�|�zt����0E�R�1ےlp��H���NB��]����ՠ���8�Oj���U8ގ3�Q1�y��ѧ=�朿A�P�i��PҠ ���ݶ-�i<	�q�����]S��9�
̭O�d/�I���7��-&��Cx%����)��ӟ�EphT[��m���"��fҸdik�爵ū���8���u���R-��x;�>;T�)�n�v�|�Ɔ3�K�W?0�J�:\�Z�cC5�<�M(��<L�8����*�l�nv'Xt��7�1_�w)��ϛq�0�H�t���~��j"/Ǚ����o�H�ۨLb�+"<�Z�sZ���-K�<{O��G�wdή���!{��\Y��G߇��խ�׼t�sb�%P�U���l��BB�c
i�h�u�N�1�s�O"���>�vi)H�x�ﬖ>��!���-� �Tb>�Z����?)T"�"�@�WD^8���=
@��EU��lN-��4K�����1mN�� I.��a;Se�pq	|�3��|"UG�l 2��>L|_�f�Tn]o#�i���@H��$�7�0?�6ͣƽ�"8D�	>{��IN6)���^D����$�T���(�~���`+������3�w�Lp�@H�W"~�M)��e�c��Z[M�������Q����3�����Z�/��=��H�j4�u�*y��lF-:��-k�LC
�t����{#�]�o�D`HQ�nA��	E�]�n��������T2�K����1�59��T�����������{�A���-��:���q$��s�R��5��~$����@��_��%Muv��?K����lҦ�����~�l�i�>�y��&-�%P�#��\z��V}E-yg���U�̘OO�l�fhY'���1zDuR)a���tl�6���T>Q�o*ߩq�����ٓg^b��f�B�mp�^:+��6@���p�G�uy��*0	Ӱ+����/���қ�d3��?�B����$߄��ɏ�M_�R`lS�B����5	ŮaA�[�8ϕm�wqp��!���IpS\�b��kmy���Y*�u]���<��]��3�(d����]�p*8� �O��#���b�s���c�0K��P%�|��%+�K%���|�R��ڧ9����e9|����:��rܸY�'7��"�4�y�h�#����GW�D�>���xx�:��a�_��#�i�8�����K ���}U�%��G�~�q�$�[��=!j�P��"}Ւ�Ĩ>k��O;>���p��WQb'�4`{�>�ӎ�������=�X�~�Q�>=�X�DDƕm� �F�8�)����K��A�0c��68$���5e�*����K�"�"��ko�{{
[���aJ�Rt�*x�q��I� KU�-���~�׍^���ì��w��Q�ZW)ܲzsp��Q��}�BoB�N���д�l����Y�I�E|y�9�
y��rΠ��|��	��g�n�WB}P�b�
��	?�=J#��V~�r,�$O0�n��/[_u�����>;�-9Ẅ��G��:�%�Gb[x7� 4/=�Մ> G8+��)�7�����Vv�6�`B�����?F�P��#�o�����B_(�~�t��>���9�J��x`��M���M��0^�b��	IvvlPIM>�g��+V�쯃9(���{(Tek��?|�����֢��ӊQ
{�S�� H>�C�Ǒ*6��΀!1p��^� �Q:�]���@-t'��\���e��6�qɂ��2�K�~B��[K����QԾ*e���(s��G̍<+Zq.>���ޛ�e���'�����z�.=qi��PF�iȰe��ÁR]`������T_&�g��p��D΍���K�E����v0Db�Vd^��?P�g&@>`��^<%��@��&8�>�{8��iRAczh���u�������\�>��R�d����#5����"ZlZ���g��C������=�_�
D{[E֯3kE�K�S	��*,�A,���NZ�R|Iϥ��C��]����
�\��	6���<�/T��#($M���{@��o0e8�$��(T��hd`�J����NA}�Ua员w�v.�`�}�K��?*C��NV{��