// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:28 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
js7ymKnO+KXMCHMtbP8bM7uSwXpn++z7OwZyXPEBjBH+CZF5s64iv19cDQ8tg9Ik
2B40XP6O9Y1MYkWtXSg8XbxxWpeEkuyXOxpvHijYVaw6acEy9tDSdk6A7BlOhBrS
uBAlYuFm5KT+AhT+3HZ4njA7I10AQiX+AKRmgHz49qQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5856)
1xa8j+WaTzz5suyrerX7PubzMzrKcVlOtlk8e9gd54J81rf/BgMBt4FoF3DCxIko
XleLHTH9vCtEWCMNhY+t9XCKrgKCiB5AmF2iRVAyYh45CiMY2yQVt2/5hev0jGrU
iD3KRZ1fp6mopGZIxESoiXommSuYMkk7yktg8+25m+iuP+TKlu73fwdwfEPGaYq/
z2J1HMl444VbQNn083SwgrDvRdVjGJrBkn/lMN9aYxLzK+fzTQtv0P+mojgxH8vq
ZNq7KjhA2gA+i8CJDl3oNImCtbX42PXU15YxMxgWjuM0Lqp5P5sQgIlqy515SYBZ
iwpWOPjneE/EGSDrfxP7yxoy0cez9i1jZazaMekeZe5f8zJtwHpcHQQ7k616eBeT
m963Z9ijPGCt9kkY4NzZTNNzxEraf0UCb7VlsP0I0NfE7FSnEPSq6+v9MeNyVc2f
jf1MKYMZ+gumhYzgFlf1nk+r54AqIQ4hTUqMlw9SQ57Di7eCrQDqhxoVe7m6Vu98
RRLWj9ylATuVJyCrzQoF4EP6QJ6zlWPD1LgOWOhERXj6z4AV7cDt0WzAx2iy6lb6
whhgUnkqBlRwb+s/aLZ2u58K+b1fI8nWXH6M6rCLiUkXIfiURl3jn9MET6xrdOaJ
d96acYmWYZcjoma8mkZ1hRf82yugL2wrGUGsjwsPJaEE6u8h9hM/gQ1oya60wnyX
F/lSi043aaXDuIA17fggCU4WrNmI1ua6CKeRKY8U+q3Iehyb20bjuW8Q6Uheb9Xm
SmOevbJ/T2n0S5PLS+4Qy84v660nmRU32U6BqprOVwl64bBB1CYStLeGzw5ClWK/
8y+KTBB5MyvBjG8Yn1x2WF7BpcbZJtIIpVb8vLxjaO6SI5DRj5z43/crv3noB3Rg
Ew1luxruZ231Pv3JRDaWE2f2RBw2BxNPoauGg2ww4jmK22K9P7VP3DItXyetacMn
0znK8e03qpA7mE846EM0rZ/J4Xp64FMllNwsQw7VKYMMyCHAD1jJy0PFPwkXQv3B
dMOTCiPw4BexSJPxeV7mpJCyplPMfsfN9VUOkWmUgY+CIrQF/R2fWDXj8vWDaaUy
Ch7qbFeKgaHxB5zpLg8ZMIatVR9UNQ6/YuG2gRsG5r2eIXUIxei1JK95YBxCw4sv
KmOqUFk/iZTo27DPr7mJgj10Up6zfkTv1qqHXRjUMS/oUmkKnPgOuiwO/3zs1NYz
N9kQk/vdu2fe8uYevp/KoBG6Z38WuT99LZ3zkWHYiTSScFQ9IRPpyO88MscPrzKV
kG07ZXI+gJfMdqCR/RPmsNlNOrVrw0pTnIJZr+8YlaTofdGQFDhI0DuJzomVpbWs
sqqXPac10BugqukemcjWaLYpFwQUJCVk3SLIcrthR4Hd97f3jCSw9oC9sc4pIaA4
GK6pIkqz1qtMGCO41U7u2hkvZLlT/si80MECFRTnsGig5FNMtluwmZSZZrjyWNz2
u7natHeMnXYQlHwqAeyujBXq4fjWKzZXkLnGxLK9NcSm/lLLWa3G7UUnVIMd7mSo
jpaterTX1r+xxL8CSZn5Zdy3ZA0Yidt2rQLWHa29Goy9XdaXJTTc5abHW+flu1Pr
wmT7gqFqAzJ7kAO9JOE41zfJe2FMUtb+HozCvDyDnuoQpN4fEz6Usx1mTQ3uIKQn
nDEGMfFITJnFhv6TicYc0mLYT90ilYi0X69ZzzvNEISMEB/1+V39wxgp7rqrwHxL
Dv92pw8xvWV35bwq4m9MYsB8BJFxsxB3Y5kuapcskZcBMe1JHzCRWV+90aoQbJFg
ZQ9aV5QPyZJ9k3sHM8tGUAmrXmX0/rckSzAHFLf3GKf3Kx6ZUf5+SRnbJkPQQfUS
9sZDSq34gM/T5ohvNCl8B7XEPfdv25OHyHRYuwYbRBoi8jM136vltRh6m61jShYu
ng37icE9+/25KQYOdQB88ddub1QL/j0EvOvaFVl6L0L3l2IQA82RQD0+tcHvC/TC
AGgmL1VRzXTlGb7y0pd7EkewMy/yo/iVJupwphaQ0D3zlnl0Dk5KL05AcUltjQH7
VPluXytgP7P+HQ6btAJaf8NVIumLPzPejwDz3vXouVB0BiQlE4878KyCv560dhG8
vx3choVUeImkwRZg9blNOcAEWlHADq89KNG++Q6GrmTf9rPaysfC1UvuCcZdEFJU
fGt1uMC26eQuoImI+lKMqzSVDKNo3U2EqmiSL2En+4qu5rU9xRbI9AHe95I/3utU
aRerVVC4yLlTEh6xiqKAg8Zp1NOwo152ltPSjwHhocpjcyj66zk3j9No8QgvqT/1
MyCVgz4HeJyP5ZH4n+7huIH4zJGSOlsBEAnGFbZUpx4oqkkqs5yeKPik41X/aITi
NwoocidgQR83dboU2rovz7ay33QCKoU+E9fGbz+jzczM4D4jSA5Gx+mlzn4rH/C4
9cP86GBNzRRBLSsS5ngYpFKHtISSNvIMTz7xd+W99Hhf8VQHxUTItpbuFB+YN1Q3
1B2GesG7aF13CtnKi+B9j36LMiW0nBpYUSo1hIQ1hbU/TwGCbLH65loL/Xp6yb98
IA1OcLKd4knf/F9Qf0ujqVPhHwgIoI1OCPKKaV61idHTqBeajjuk/w1h+mqtCebC
u8NJyWWA64qJV86xAf07Ss1Cbz5naJkms3sskp29obvbMsHQ8NpU80kXWPR9xboe
hbyKY7lUObyvND/CZpy9+uJGNQf6rEZTnoE3yN/AiCp4A0fpT3AbFn4TqA+5Vqbl
9W3AO/6X2a++ALLuZXDxDJSzq9dXEnMp0UtPjHah+e6mqs9+UcIj/y5d9Q8ub+ku
Z7gK8EH+eNFwvtnMMHXKvR2mW2viPHiKa+EP+ZyamrDms58gOIjdJUEpG3Q2jA2o
AIuIE5DQQ4Y2orBu7ezlficuQ69ZeWXs8m2zQ4TqdI+JlBMII8WKiwf4/w9YqekX
DY10rdC7U8g9nT10FmnA+wpc94RwYw0H+pYWexmJQyAxBEwhjyr4GKF9qZZY2Hy2
d84QlRLUIpQfAShmhdGXpO9QwNENJZghg2C44hKLHwbYBMr1/0YSG6NCYx2EBrIQ
lR+7C0U0Wfc7fCSyDQgjGtxBjgvar+Y5I2Rnekd1slN1rv/8747MUfs+D9M71u/H
Ti/hjWUWu7ndck87k+pn69GouOBvDDOoy5wn4RMT2f6oa9DcOByIq7f4SkcQZRUL
hhiu/innu6qLeSNEL4s6q6YEm1+TJofGXAYqjicDHv40yMaLxG2xgNfCEXDPSz4k
+TBZilSNnn1msZWBx9iZlYDSJA1d8I2LL/3ukS13cg4NXpu3SaC+y47wkIF+sGpi
XEuDgoM6k1ILUN7Q57t/aB5G+9z6N5Te/iP8hpAKVqUfW4g2jxX0vVwhxRLKUxWK
F8eDlpv4xRH2IGe6ibrxxqaHul25d9PHQ/264BC6CgyU+xBYft8MZ8a/zKhmBgKi
A2LFPteP27kgw/yR33crGcyldjP0lSABsp7SDqgsuxWCfKawJlApQQFhpocQyM4j
5xkLwEcgAXnyJjYv+flMQ9SGTwowcTeUo095cPVQIfqu2A1FirElU18iDKINN69y
1mxRuVRoFoRaCPTHPiCcst6kshsez0Euf/FK+oWTbLX2l5TnffHP3X1psSuGO9ei
odk0xxNckftVO8RX4UvQltan2LnO3cWIX75/cLGzX+D5fkcEgMvJCrxoQ25ZX9nW
oOmfCe1dfpLI6mIDT/5crUAFV0oJ6zM1hslje6k4x0O9urc1QTkUpRVaSGKonTLb
BD+PecjzTMA3yoRvXUbrR6DHG1U0EyJiCDhvXJu1oEW6X/ntQb733sEgPwnIz4AI
/c0nNtN+43fUlNYJsZiwLCBOL4qPvk2aQ21kZtQ0bj0aL/EQbxxWamcwnCZPwAP5
3Xaky4pA6V0IdnS8hl97U6zFQoXJSYE0do8G2rXIjEOKnu1/52uiv3Ywyaz+4fYb
MTJSINWZmgSToLkhk9mW4BVJ+GG6+WeVa9tXGbvRH8QT1CrCfKCBgroyyr5MW09t
anSvPuFboMxAlEUw2WPHRDrGZY5mLKYkwuKbl06CWq6LtLGgS2Qowb0gZ7yVulE7
0Xx9sX1UNdF444fqxzVyGijOcN15BIGrd0/v35p1MiTEFMSNONVjSWE3DEPU7UDV
yGCLZwTgKvKKw/VTKkB01xQKJM8Br/dbVhXjuX0VdqX6G/cG8TP5ZNdAGnZZr8he
VGkdKMyNSBUyNGYVJA00OuvFG9wkLPgMUDlQ4xBmZtp+rRRdxV8AWxNHBchfLj/1
hwYK07RLsGM0exsBC/dgcKUn6keIKmNyzCvG30qui3UbTmBnQhc72T4JBUuqJqKP
06EgSE+1VlpAwKMU+AhjkGgG0mousQ0FemhpUXZnXMA4S5C+eu5pYg7vQ4hpj1Ne
mNXASI98yQY3n7WAXcP52N4Hp27tIkpwJcOfVsc8fx90e12RwIIVriD6kSHDUi0O
oqBl00VxSjg8yMf/SLjUnF65EQ1itKxEvFTCUBaHdv2D0OZaDGUBDk3fEpHc0Wx/
3QCTAvhvOal2nUx9wFtKWjXjlB47+1qZplkQIJtFRKkdh1BOSdh4II38iZrADwcf
2JZuKIilG/EhTUt5maBI65ePt/JLPK3oAW6BKkBwGh/WthtfTozOsXcZwk4hgws2
Bv/4KqxFO5rVQ7UQCiqyfwJjytj8Zv0d6HYp6SKepx+IxmVdhBOcAm5ZSw3ByUF3
63czstd7DEWmJCN/rAtEmZpG7KsPg4yglhJ4pmGd4sYj3/2KIiTDoZWO9X9dciN7
QNJTqj2HoLvKFq3TcH4g30C9JOAP+S0piN0+xJH5yS8DtSSOwCjtgEtz4YmGfjY6
J3lX1O/1/zK9jQah1kEftu8Sm+4yzCswVpkde/dF9eIqIsyQUXyiyfGoAHC5u1i6
UprTzAoSNzSEYksvP7jb3tLJnSk+abtja5XtIUSs/KOif11buduDjcNcS9AY/Qmt
k7++ss3pXkb40EGwy70Yees6vlaI9uimR96UDPHwMvo4sUGyB6KxtKfeVjphowPl
bj9rGQypmLhf1p4+dVFITZXp+R4Qw/2vMhv5QmLygrqaCXg9PtLamys9W4+BomP5
SZHwajESyGTsY8cYu0Cz67Mp92NRuNXb7R4bDpy7x7kba6n25BOuwd+FgFGiXjga
mABcY9I8JdFHmgVM0cojSsmJIu4RhseX2rRKG0ntlLQpme/sMpTi+ACGDtri7D9J
DrorqDch708eQq6nZuy8fNNCHg8c5GYLS3I/wKsmtrSjx3afv+4RKg86v3RQib/e
iL66C/YmNxbxu8Az/pE/EH3kYdNVGAErB5tqFDKEDVytVGJN58LrljOxcKptufYs
iRzDSiIIC8Jbc/dbrqP98LtYgmkL5M5aujjiU5LsjISPmXQitOUx3yo0DWf/KsoW
YFbiETdwV4f4QGZzajlxtfJPd57SPhYrKqMKHTQnlINC7RDAChVJGBWQlYRj87hI
W1uquLqnVDPVIH3EAI6inU4Y3QwAsnD/WkXgEVN8PXpxoDkq5QndO2yjCefNAtKQ
mPQrWVek/d8rxJL5c9dvIu+7VLPU9jViQ05EdRen24DEu+7Ac+g5LPaxQQxu7ukw
XJKxxM6hYbMSVCipEVuudWy2TtuxY5i3qaxCupvtRVGKA8Uf9hg9wWFZi4srnuK2
sKF419Or9bJUDYYiZ4P8I+hCU9jP/eiTHCQeeUsss4blb6+xm3XfBBtkhYVUhAd6
zgifouxp+CMqx2sD6UtyribrEMwoXkpnfilBW/wQPyyKd0N5PjSRunSYEW2BS6T/
SknjntigxsUbnvvtESOizhbQnuhQ3lfr58plOakIwmhWjTE9MreeF91aTLoFg5r3
IaH6VfDneXt8HCVCFXT22VrGINzQM9GZH7z0J+xVfSrmeffHj6DNUj3nJU0l/H2i
B/krrrpTaPkcf3HLGAXyKTG6ZvtF77Ly7yMzA9WOrxj7G7FqxvxB0S2XYn0dC7Qh
RSGkdPHSjA9khB08xWnUI3vdKT+iSyw6/nmtbQUPOoemWcymGq5I9pHupfjxcMhG
DKLLN+207bU8PliH2V80CIIf7/mR9mLSOxF/KkibAAwY9j+bN/onGg0dbm6Dxd80
uME38mWINrxZwbpXDQFBpmiTWMv9F3BlJfVjejETKQLpnDjAxLs4nJ5nb2BYx3md
rcPiyfg+5Pqi7zX78XB0P5Wh5+ShvFLxjgX+Y6hIGXpI9ZaXZzAcbg29FcLBlHcQ
p+Txv0TftnndZV6vXTOl/MV9Y5Ox2ZBr7PuwWSetp0NR6zXXbZPdjsXfGSD4kxoE
8xRh1xYVuyrBSXAXniQkGoGY/EJhXcpe+84Fps2WeKqbTg7ZlvmrVdet8QX1WSEd
SgqM9gNegWxXOUMFVm1dht0eu7/+10evImAMmetJSg/x0nj0n7GrM2mOflARRJvq
fePeiRpiPW7H5Fucj7JeXNMBt9qWmNykPw0goxsTh9FIWmVFdd0ObsFbNWLw8eX0
Grrbe5nSKg32It68fWGiFj6708cvrB+4ow/6N/7lNC8klsmG1sb7IXUenY84NVMl
sUHHDGzCT+Gs9leLZZMxz2XhLKkiLzBJCrXhsbyLDG/bwkzz9j+FsPFLLradu8XB
0t8sn0lBq2JUa6+hiYGUjRIXAyresYxiC5qX9tzKOzelB9kvoTayGddaMIHo/s92
lscIsZR7P9bBtIyGyG3s4WXfcciW8yt79bQa19yx4WuZWuoCjt5GFVgNqmCtgdvg
HkrJxZxk2yyhh+U5562UA+CF4hLfj/NTItZxjCvRb9dvrnxX6i49EdxuO0mbAUqY
nIRxk/4P6Wy6MJKRP/92e/8omDqHtU38bP4AIkZJow+ApubirdxmZX4zTLCMXJ+b
YKJLINDI/xUkcl++BmDCxancLTaVjHhOrkJsHwTjP+ij50p+MQK8PVPi5oGHhpUH
6kk/mK8i77EpOD9JyjfT/RP0739BfewoDnlGi659GN42K8Q3kgowcV9f7wR7j4jj
jmb00sj8+QOJZyv77UYib1fe/tGisk2g4zKCp2YDeH4z9ww3gWB9LU6NeL6uPVKi
gnZzcQU/zxY903AHAosuiOHsMCfLLAHdRwcPWaY8LrxqrCr9vCYeeHOtDO2EZmmR
87rR6aVPmij6WbydMZ7nYGuwvNPvvi5q0bKYQHxVauyBfdRVWdHs7qY/cBC7hEd5
R6Z4FquG0rhNFP+PjZ69PSl2l1ufyC09Sn+XexMWtBCml7rfsYrjkCfFyzPi8rkf
uT+6/bT1mqEdz5OWmjmKRTQ8g65LO7v3qeQjZxO6zqI204b0Dk4FuT1y92xxTeRr
g0r+9yPzsbyV/hZxJ0Hi6BfKktAfNdjs8WPf0B2OOW8MAEj6kHQKzGxK0/uIMICJ
Rxp3jihzb+xsLRWuVPzRN7KVggyUzbktiETBg9NA5tqEeHgIQX+2DTuUND+2ZEkS
ciqvMv+MT4dYOkUtIvvfyjwyJyvdv6gG13tmOK7OIMTuqdsbNbjK8N9bsPJwdSBv
eeU7XvyXRUpdc4++4q6P7dqFrpspWddlVVlLG5kYGr2R0Mbe2nFjqxBaqmIfNZPa
HTzQkzcFWowxmZbKoOQlhncKYX1xHZZU/sI+s4iKUuTVYMabTjqA1L1T7y2pUoVx
WWV69CxDTQ5L/VS0xokJq8WY4wtMyDjwWPaz4nNisn/I9mN7N3OTd89naQxU+BtE
/B+6t+cUTrU0GLptGIDsMfAPEFI1obIAXDRQdzwjsqzWjjKKTbcYu7cjd7KD8Pqj
`pragma protect end_protected
