��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħa�gU�]@)},����ע�>S�H�������P���2��=���@Ŧ����3>�7��$��f�\�Z�p�(Ű� >� ��)y����\����`��N5�?A��(Lރ�*�'�-'Syn�xVё~����caK#dz��#�"9�HuJ<�FP����W��<)��K�UD&�|7̐ڐ"ݜhbgxM3zPG��Ľs�|��p-.5
UF�	V��;����8��kh�"�u���-�j�҃�������>��K�h����4���B��̪ah��Fӷk{s�_[TxS��{<m6Y~NҡA�f�0aO ����ֵ�����b ���l@��K�4��n�5�uL��N���5\c(�(�БxS��K�^�ƧN��F_*�הm�j���Ƒ��0��&,I-{�#4��c����
.M0�Й(�iK<Bm;�9`� S�g��y��D\���nLP�����"�.��9Q�s�SӋ9�q�8���ӹ?�H��8}I>"����#��C#J��%m3:��ɧ�mb��#�.�J���E#쀻�@w@���Yt�����Q�N6؃5Z��)/��)!������K�W;* N��p۶	���C��I>�~$m�9����J�:A��>:�=�L���������� �f9R��a�#��s5Gŵ->�Els�r�,rX�a�1�X$� �������� �k�Vt���1-��=R��y|~[�����@|�_I��v�jl��?p9�o�S�Rg�
��::�b(~lZ�VX�7hTm���śx��\�m��g|�� �7Z��S�H��`~�{)yA^��R��N���ݿH+�������܏��GM�`U�U�wx��y�̢|�'uN������Nc�QF%k���u���.���r�L��)�zj��)p
f�Q_�1�#��x�Q���gx[M�����Ew\@����_�O�M��X�H�5XӺV��ڞ�=�߳���F�6��NV���Q�"!���|���U5���&$Zwwr�?�%|~_}>"v�ʍ�%�rV�Ĭ�[�ڮ](�,-+��;��R�e3��n��ZT�~j6���{~�#�?��a$�u�"�'�t^��Sz����,�����i��{Op����<)Wx765_g�k���u�M���<j2�<:�~tqC�����4�i���2w�J��/^���){��Lc�,�����������a�x��%��@T� ~��h�ܭ�yB���K	�/ W^t�">G�i�^Mܑ�͌3���0��1�e��rx��H��	d��	%�P�=���£q~�"p	*�nW���#�YJ�{짜c����;b3��9�(����-lQhs�Q�ݝ]'y@t͂�c��&x�ԓ�x[�M�t�K���2��q�[�Q��/9�s���+�GTA���+�&g��V�l��+���.�KV�ct��p#�lC�R�֥��k/�A�g�L/�q�mND�c��n�Gc��r���o9Ui���;r0HJ��k�a�fߌ����?���k�sX���!�@'>F��Ϯ�=ǸU�#Am٥�z-v�:�0K��oEk�����(t�U�$W`��c��-I.��6m�"0P� ]ˁp?�-���稀>`E%�,���D^&�І�