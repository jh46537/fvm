// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:32:15 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
d7zZ1Ce/KfFa8AAytZ1C2KTujzMaF1vqdZUuRqyke6lZSMQxtZjoM4WseIBiGsVY
dZVRSyZ0Q/1rCvR7rk9Q4yx+F5xWtOY8PnS9vRFGJ7sFAqfMQl3VWDhq0Gg+dJmb
gvfHsu3UDP+xrne92uq585zI0C6RuccxFHtGrbORH8w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 74896)
aYNQ5wwrhXKzo9FI2fXp+/aLrVyUbIVbreqvYDxTxC2cg1ck9muBQRLOD3qNeSuy
dnFey2+H3oDM5AErVRhi6nxg7aSfzK17VxJtrtayxn8M+Vhn46KkUJ8PSVPBcokb
99+GGcxvgK6PDKTgurlEZfm4uMINQGnRJIhpshjTg0VNQL/T9hTzJsEyd8KNhKZ9
K1yeL2R1CZaWh6bQwtf+ydoNGjYMoKOVo63xfgTZwgv0xf6Jvzm8BjfOLBqT7ykg
aA3+rB6oWuMLm8S6zA5DGHkZNm9d60GDvo3Yfcv+Izunm20L5CSB00GBglx/9iUp
AUgFQovO3Zx2OB2mvM6lMr0o4p+F1YxzD2k1WqnkbUkMc6UBInLjScjky9vket86
h/Aog5/QhwOoJjtnDZ5sfrF5sAEkAzBPrGK00tMLfuhQaEhIj4w2XqUCU1P0nuHX
DiKchiPoFTo1EHFQ66vu5cYAQBMzTCvjDumJ8fpiAELfDf2ZScy9xyCq9EL8ujQ/
Rv3+xGAsoY35WSO4iTELtYft8AES3S1AC5ZKmWBv243txs13xFPcUgCXHDO0DEKk
wfy9bkCnvldRnrzmbcYO4yJSxTL7ADRsuqokvmz3OaXpwZpzcM4h16I9enjYr4Ay
EIzYDIaDqJ0s7CTlKXsE/TSGgq5p70+DE4hum7/dt4d3y/7cxMCG8CBigGGwut8+
qS6fBGw9z3jis5/jbxD2yT9SO05FeGlKrF4FEcButY5emcl43+cnJuI/HsU2Gr45
W+4NlOE4q6OBY1YJvA/TMlYt18SOPh5QCYMi3iGwfxPJvfl0J+WG3+GBRiCMbfHa
4KlhZ7I/abx5vlZlvRUaVJLgzOOo1Cxut/x34qaTPtI48eCDrWeHY2ZlD0d9a4rA
VJEv92V3wvfhS5GtvG8va6OCyu6fCkV1yZTvECzLqz/9oc4RZ6TLTj+baP94Xdiv
yMwYIq6iYIkZ+ganDZflSeXlpxoEymORhMIVv/j9BvCudk/8TcSFz/vXlwHSM1y3
ry6eHHKxOIa8VDk1CcVv4kg8Lih9FosJcuMa5O3J/rbnydI3FaNB0mt3BE7yIalf
snNkMWi/mEMniBnGO7PdJVYsFLUNGv1zJ5o7B8REqtAUTQptTeavgANHFOnYzU4+
f3TO8/0S5z5SbBXSGf72csJo7kCEsXXKsteeuh9ZDoMl8haDZYu9SPbdhQMEpRs5
opnVTWix479ctnZlnwQiQ52dDYqeJvhfUTEBbW3ebv2pCpoVStquUckkTG2hLPpQ
370xHK+VwJZg02C71TyiSyPYR2Y3mZblYA6CWU1xdRs50VqyE0Rdobg4cmsTGoKL
9yxAnviIR4pg585Z+RR2Wu3zgIgklpA0u6o2hk5mS2sMik3+6v6aIoafstfCpySy
Rd7DtVNtJrcxqJinJboIkSUlsMrijGrQ7g4cBInT+dzkUBLTy6LOZ+DcZLPxJ53w
NPn3H57nE3t1NHv8AG/hJB4oyRtyBeDoDO8dvLQJqxuS3v/M107UPXakX4ecScJ5
CzkI8b/rpO3oFoUChbefYd79OJZqRZ8ppoDQe++bsecojP7/GYCznzF5pGQyDjo7
2tzNJasSiA4iaCY4JnC/t04U/Dx/VBtDKdbWIiEMLNMf5xXdeukwevRbWRHR9hsq
X9Oj5JURoueiOzIKBPEa6+0Jd8AqA73aTGcYOLdhG7vO+gdZi4LUimzwS5NieT3h
PJOBj2qAhCYnt5JatseaJP+0YZEKZRdn5U3pkFOf1h1MVmrLdfzOmbiA3UugePdO
26Xdgc4MTyhx6ZmmYb8j8cNcmm6STJqf1eu8pASGd2Z/E4QU3t1YEy/OwJpuIcJm
6JRELXc+jiuGqEkjc4C1dHg9GXs4mSUDIwMGpqqvF9/YcOHtcTVYgPKQU8oci56c
UIcA1+sYqwSE/zQZwwujwoS0BCwgpox0l5vNAP5dpTuJQCDuyDHj+FclVOwi85t0
7k8Z4YnoqUEa/l3VTXB1iE56UalUjyd7dax3aFJ6vKTr7vsXNzkLmvAf2uBgVoXt
m/VQfJiKnHJxQtBN2pLnV5fx8bJjvvtVcEPfEwxvICzIRJxl5eXT065Kw+fnhro3
dFUipFBsoHQlYd1/xaQh/8A/EwhpxQc+4xrl0+PxeIfmbU4e3jdmtVyAkGjSH8fA
lE2nbhYM3Rk2GP22lzsnt+g210Tjg9AjKaoBDVL3tm8FqulY9YClk37tgysitQ+Z
uLjCPStmxL3JrwfygwXrFbvwwQD429x6iqAangHtW3Q9dEToF/SSdVxyePLWOUWQ
vzSp7RBuiT4hqeMZXZANBFmMN3pamTmxHDUhqMH9XaENyiVg7CA+JN7Wxlec4LwP
yyEkLyRv1BeTMk022UXelYUJKQS7rDee2XF20RwbL3zVi8GaIFJHu0irXoEsFwph
4hjlMCgQZufyrFCU6nmyMM/2pq//kotxtgDjydwxAo7Skk0yffk1ODs0da83uMG7
1R5hEVhCmWx+NPko7bZpclrCF+Ly38aNhIxg7XErtPr8bjoRoFNJPTg0IzTCWlQD
hvZDB7BSeWDEvgIW7paKNak9Ol1Du26Lefxykl+AEkV5agBzrBlElmnbrNYeseJ9
TbN7cIAw22SI+m4COB/L4ZZlWBtvP0AkiF88ems24bdrpfd0Fh+KWBlwpFbWYt4f
zZkghItICffQdFddvyebedWAwZMA/FUNY7wLK4pnySOpQnazq3LELaHhjDfxsfPI
xlf6Rr4ZHLm49Oz/Ytj2Bym9oXWTrOsMF1zbPtdTI/GJuBpsLgmWhpfLK3TtygKn
/mBSMDXv247+dWmUUDujPWOskXnaam0GmI0mmHmzvJcVIECk5ac95OlQ4tsFljPH
SyxJyU7XHatyb2vN3akh8oYNDueu1klmVTtwoZVD9bc/onX/BvvHWE7vPTtMyrd+
l3jIan50iQX7Eyf1dam3wwkxmei77L6k29cqwI9AOPK9mXIWAUMgRT0F9iChHZbu
rt1El/56YO2xZjtpoSPlyg1i6zFbA0VrJuGXjRDy9VnnI+MqGMsvZ1IjusKZPyvU
CfTI0gP+423cSguFDo0mn8avQb3GeJI3JmCf1h39VMts9Yskj/zYnpAzYH01FbLT
7TBBjZLl7NsqDmK8/3Uz/dmVmKaPcsoz6memEvuGMLWnNexQB5osHH9Ff04bR7QU
fwjcaIdyOUGgke1eFxgjvx1wueSWnJlVIPUDSTRqszLbmmUwPXgq8e29gfhjry1K
crV0yWOycsHLqYhDvo+gPgMh7r0BpTpX/9PN6cx5CYZPtN3tbLu9yoDwJzPlV53v
sKjFqrY5GFC+yQ/o1Qhpm6/tiFX89CKal8kBi8THdvtUX1f4ntd21bu1xkwmydPG
X54s71muSIMi4fFoU0qRpOC08LOQRiyY1+ciZSrAAD/IJKE5invuXac6oPC1hkaY
Dfr0Xv+fS+bgr5NZ16ek8PTaHi0VHsUq7WfSv8Rmh9/NKMaIgjnfRqLESxCEDdFB
BOqn85LwsFCyUvMj+M1G5tK3B8YTqzFYhLX/VirpMfjqolGJfNnqNtDx+NaCil4h
NXvkusSUN2DWcq+xQsX6mIeGL7yXs/m0+T4HSDuKriQ4gzb4KOeC0xbW76ehtOlH
uD63hV1HK2RGqePb0nNniByZtJNXsZSEtoZdbzkkNXrwOK6oW0JtzOz23gx8ZcHe
8ivhQZ0O7P0Dro130KhBB88iM/ZW1mZJW/YsNlAUe+zbvlLOdM9Rf0wHDqQbCO7n
hFFYgXPNW3u0RVm7NzkVekZZhZHc0DSlOve6m5sIA+NxBl3gKqE87jgF3b24WlgJ
25YEqAq46RIB3p2TSyJzTwxia2P+nQApm0YGbdb4Tfunhm8NxpFRU6O83kSLgUjt
Y6gSCGa2j7zhS8aUuMIYlLGGkBO8mixg3AXKBJuYD2gaWnpA9o0RJA/6Ub5hGZ1P
PlM3szgby6W1q13QYczYGyNiHdywYCJ0VJ5KxScNybpougqjuklGtwF5sJtHZTSw
DY6AeJZAi+oeiucjnrp+9/56QLeVV/IX42J+u24ERqwiSFhP2OWeMzvNUQSmkOba
3vPFmx1/TszDQc36FppKuNyZFpQ+1Pxf3dAqKC3y5+sITC94BsVjAMZNknPfifXb
Y3qt+hgwdEeHzkH7WYUNgfOY0rYWq+oH9sH4AlHtzUAG4xkuJxEAhI707D1qmfgY
L61oAiWVsamCJxBUUPYHffrkAIUUOd5hTE51RzCulLJgPoE4/KsveqlwE7uV6uSs
NWvf0PdFF44KzcK2F5RGVH2QVRiXEm2iKsuZuPw0MxASSCfOiNvnbZahKIzKwiBE
MxrWUyZeqTBUwlPo8JuXYh/eS30E/BrV0bloXZ4Zj51e4mrC+o8xsl2L5sQhtxUv
QTsw2/pwYprakA2D/IuWiaVSXOanSeLRfDwnaDCOPgVR5bbiCde2lpIyyQzQ2qsc
wBUcrY83Xq+3Dxkq72jlWId1xj5aVk78jZyIV1iiKqkjPaaGk9DGxhyOGYCAtQhP
cGbVCk66jX+biWAi+iKnxFFeX58qfrXhG/7zwlNzcRnpHswJ7J3By/M/evw+447e
ZStDnLc23X0cZFBvXR2o4KcGZuJwtq6vUXX9QP8Qi5nBTSgqI2TM+8S6VvOAAnwK
1E1g5opfHs+NPHaMP3EqQh2ZIUka6b1jzilBvCilyTbACOt6twyOEvjELO1gzCrV
jSfZ0+u5dceTfoi3so4xEr8DxNWWnPiawQgY1GqueyLMi3zR/c7MAUZ70SYJAy0H
IHKriT8t+puvijXa64jO5QGRKsHCEw9PD2uat3MB72yQZx/DXJgibMD8qqV2+gjo
ySg42QHxUNz4H1FBkzoJuxLUvu1Sxz+PBY/r/h8wwsH17JjgIFDv7QxAI9Vjg/6p
peqekB8ihnudpgaMkcriIKo0C/KNXAol4xWdzrE8fX8yzgtAHo+52uPQmWJRh2D7
JgHNy8VVuJvyikLk+k1qdlm/hZeNGbHLY650fMcLk1L098YD8Ao9C4ThUfTMUFZL
jhWuO6l3GJeqdDvqROGenoi1OdCmYOuRetDRQV92hd3rRziU4S6anmj47ox/MyzU
UcKNNwQ3P4gimVXxyvRMVCVHJywK1EHvzVE71O9SQyZz2K32aDahFJt/glJb0g+w
qqf3/ftUbi1LxZTG9N/zGWCNMbAsqxmVBvJ6uEJ0n2K1kPL5PPHH+/vowaOwdEbU
19P821Ali7ZG00SDSlvJj1ildYWlicLUo+a5+KbSAx99a48+pWdMiLrQEBLtRHko
9RCE3uFTnqd84eRAwM3nrMXGIHag3XwNVmgasoI8gufi69ojRgCyegEsNmsBmqle
1Pu0d3S1AQETmQLqAVtOUslymK2759sdSXvP30ZEsKeK/vP3M7j1FdmRlDbW8ht8
q0+k6+gFP2bWQC9340tf3W1alfVLaZi52EtT69MPs3Q5+b32vaII5+yukC4J0J7c
SHv+gDxsF6GBrEQUXSnSNfQGM2ycL7RDX4LElEuDAqF+4oAOS7S1PxRwE1gkXBvo
IFausKUQ6FkQ/IDoVnkmKjqHxB/0/hxl7qER/15Dovvc5UtefeIGv2t6sRlFUAoD
E0YHchnVDmK0mkjbnho96lJs6vSE0fF9VR5FAaOpsAJciI8z7I/hGxPOjW2rhKPA
AqpRM/XaawAf/uKxo82CRpjtAH2qg1svNpVbQeD0qPBxXKqVtROtLPruIKWLZBuc
JaO+resMba69s7qRht1BTd5gTVTmQlrzdN+wVQvFdzGhEXKLyeUaPsDNbLViv4oZ
xBplLW5WpQC8rg4ijZlbCDXC+ljKlMld9ifpTwU/yHmy3hR5riIYUHUSUNAful1V
fBQvlOJSbTcUdOy4OAG5PFNmA64t+LhfesklCoauABghkeH+uAuVw7KWJ3WNvcPw
4IIrYouDZ7ofVvzR7PPNQJ8ePBlx9RFigccQSJhmCIevmHznXVXQhCaAh4kBT5Tr
QCkyv5Obco5DWSx65/IPqVEcL1E1M3XAwOgY3pEr2h3uwzQtNttzGeoahfzuBkZo
wnIkBOwsqCPuNwHCy40kdRpAGihNkTxpZJF7yVUNHut1yaIb/UWBMCHzOJ12fawZ
llWAez8UIjfSJxzQd9nlX7pnH1YDun3ylPeYjGGLasujCyuGk+F12aFCP6y5PCt8
IZ3nGFz7mDDd202Jvh43BRM8OHpXpNzKBObvbdaGjzKt5CTv4Y67dG5qVivZJ9xP
/3yttyrUODLbl0C1sgb5ml0SnqAU1vFhxQNafwtS9+2lEOj4M7ZEiDU/4BFOPKyv
vcrFxIAvGZUg2GnwqI9GPwD/GheGkTp2ew3M/uuffs/a4jkBylQLo7ocpXwh6Fyi
pP1eLRLXvTl2p7q8ou6amdmGJhG46qtBDEFi+HOzohrdpF22iYsefns2L5/6Iua4
UMGIv4ciVEunebgXKxcb6d5GZdTHkyowvhOYZeVH1T4X3pcuprmgXmzDtFdjSD4y
I1HiDZDJHoFNoKVyKxzHIQJdsPQ1DPCE2ZXAEIzykD6j8QPFxusqYu+whN16nbi3
Xg0RSSW2qg3oQAJ003V8jWy2lxKPk9C6qEnuDIiK3gPOaexO7GlBjemLzem4/cUK
q/Xe5eDh/nSSnjZhxzwhdrSsc3A0U+fXOklXfBtbz/4UaAJpy9XJAQRsNJaCwXtP
fDuGG0+4oCloxnEIpzYpN/CFVhdsgUCou6FJqPjNfe/oKOfkpvOYjVaF/fFD2KeV
v4TnM0uPN7+MTTmQm0mbOdzBslehwEpihmAo/Dpe3g4CpruqetC1nJllza7BLq5D
OsYqb7gafZCwX/beEvNUgim+wlLeqyE/2ULNvQ+pY1FIfm8xEOId6qHGD4dEZmIJ
Q8PPEJ+glM6HIKoMePdBAUrHpy1Lmo9FIM5E0ftbMvg2nk/hCrhbWtI0/LkdqRS1
8of9HRBiv1J9eVN2NLcjRdtg7mD/VnxGXFP1OUEdo264JYtdI0T1iyr4J2rVN+sg
ExwZZgI5fLvmnc74O/xZi3l4dsVJgVxmXQTU2SIxd3VHnPPpgwqu6GkFL0q5hTLG
c5BohuM3F7ijxd+40qVvKzvNwrFMBanKsINZ4JRRkoJxjaXpMunU1EMWZaN4/OOz
mxgFVirQ/POMKD5dKarfuqv83UbficCoG7GhM1IFUGg4I9nMr8e1gfodwJf1aQLA
M7tGYSXWGefqa6zSwbxTqI/oKQV2+dXT4uAmNNwLnNO8ksFT4Ai1Prsc5s8JQf/X
aRv5IrHnv+3VWG0Vw4QytG+EKsWAMEh71E6s2w9ckkOwPN60c48+BQL1Vz6U7Ph6
Lm1NM3XKrssOEvgLzjGv0lI+h5f3K9F6BsIrIuXpcK3zSsefcRuQXkm0WpJx1fF5
Wo9IzyB34t1mAlvKaCgLtSkwLrVIf13LG+TinB+ifsVUuTDHhM5SHeW9t5LPVoJC
q5qcxHBe/8e0F5CyDcs5XBvVX8Eh/hdwW9Jr7tglEcCelXjWTueRoP7259pCBqZ6
T4GrC8Yz15zPg4VQsuahxEPq/MiAd+xokG81yM/z+xYpUORC4psxiMauI7xV/Vqi
2yotYD8nHn2T4cbgDp9wnFVg7yLBoS0C4BC3H6yCBM2HqUSsEigYaphJxzLAxAPK
rzKP46ppOH/rDbTgI/oajy403Q2xsBbLqRMX7CTVH1e+V2V6OME9relvzpfx2urf
x8ikwnid7Nb9gLNR6o3SccDZbbB30eFc7AwR71hoSF0odHDHMAVBIsiNjdOl7OAy
G3cnRtYV12W2lOowTDT05KWY4pwaQYrVMjsWUaAS9Cs+9QB1mXuYHfgT4uy04Vjc
OlDg+/5G1MhTcX+GVwoAyzKwclm2TVLU3ZUdjaq1MMK4JxZn72gvAgoNL4oqrmcH
3mD7SWBBrr4FCgGHQNvrtw2quCRffRtPmQn2/C2TQVFKeChXHtIxlN5/v3N5JBie
/191cLQn4szMKYQRV4bbMJuBT3qis7c4O3QTJ2MNr7mWuZLjrFqiSKOrt2dnYGw9
AN7agvGpips5/M5ASO0ZGqCtXndw+U6R8J7OJL21GKi7a8YIB5PsYHQZYM2mLin9
w/TW7ikVvAuYTcaDUiauirhY2TIkz5ReNjCern4gA5TSSdFnA5WGWBD03/xRn5Ps
BozEk4ukjMVYjkjo3ZcLbN6PrHJmrwkIuzBE61x9NmbR+kgbx/h57KPJP70fDJe6
1sqCF/KMb2yyKmPd6LtOidUXyzuJd4DUREGVPr6yDopRDYg1gS/ro8U+kcbQ/uA4
lgx3atZDURFeMsIC2CQDV+9JT1Ymyd8q4MWaMryYkelJ6fsvZCJvi3yNUHqrpYZe
4ObddwDK9pSqYKBAi5yJVnXKfjb70MiaOA6b2g3l/X+BpQgTZDlmue7X8IpRNgJS
jy34aJsaB04goxP5+FiFb9QqiD5yaG4GU9i9xBXMRRLJiC3UXnbjYxhsWcCng2vy
8kFh7lkqwbY4NFQf0yBvN7RtzV4sDoOmdNbSpsgcgRD7S+Amfknuho0GT/NxEYdF
LF5qbYNorL3xsHcIjIADLB8z6f9PAUwixvGRdU0nNU+ABT5UWsF6SP8FAVUsABIE
dED4e1hQCXBMOY6/vdoY5y53UjjzZsKGMznJ9oErds3t+p3GvOpoOFR9NLl7nBmX
UQHzX96RH7KlWM/s53hdKz12mJisE7fPVWH+tPT/J1Dp3J8dNqrRPbbWdWdZ+U4o
FFCtoVuIJ+oasb+1516QdHlgPqLNpWp5UlvrBbOzWrwBaBRQm5e1shRr2mUmKwwR
PSxcksfeBwal3+8AE7PKQFkFj05YE718sDahwG7UGntHe6yV1jV5c2SvkGwTO8Wk
vNl0QnDEnbVJxky701uMIWqtipPS9IE2fKZz6Aahr/5t6uIyHq0Bq8YkLE9sGdvM
6X+3EKc55SO+xa/Mvn/PCfvLrGsKHbtYFUxFaOyo7ba8fMKkv61RruQ6TbJwEZTv
da/pjBnREZRcGvUY5T6qWUVpHvWcCQWTQx9U/zaJbZeHwXD563mbBMzFezZZ8Ggq
BFm+1M2paxyxWvI+nBToOC7abWp3D8yaRl04kgVQE0bEgM79Wkue0lgwHn/wCkfJ
NE8qLAsMBqwEUvJQHxv0KjuE9YuHerg/zSNnslKdqIpwp2XEiuYdTWPfCcc8t1km
t8rfGKO4T+4yKqEMFo4IiCUgXLZhvnG5J5FMQNLG5YqxXdE7WGLs8iJBgkqUfKge
l7vJd0DesJ1KgGy1LtRzEP4Od6eYMG50bz+c7E2wWIZTwEk3eqg6h2YgaUNK47g/
uh32jMEJUsgF0yRDKckQBZmTvvosraeW9DL6dBZ9YaPK1t8hcDkbluNtKVainTCx
xT/2iuaQvMu49jXzKRwpJax13Co1Kmss1edNNeOvDJILyjT8l8cDwDiuodbFJrEk
NbfQiseJk0Mqars/3WvczSlBv3SM0+LidloS8davRDw17RW6nrFD+0MhSPXLBeM4
+Do2jl0jRL/pEmfZsgco7qBwUlkK3WnEr0CyrcvC0FB93HZmaizGGhwL6AwZAd7m
TJAa9vAWhZJt839+4DTDZwGDJkqkwCanwA9elILKdw/c+PD4Rh3dhaow628xNun+
ffyYxdrKhplIeVZpDDPdBcXx6FwQXPG8RwKCorjE5D9QayaM0Vrh/89xFf5TtuhR
mV/6A7t+ilVG54IqjJ5alUj84ZP9FsKBwaCVMAar5mSACg7+Cmdsezx4zb6KAA7Q
GV/TTrlKdWDSukagy6W9R9A/SQY+u7PQGAlj1D7y97jlLLourULVzqbKygjnTAuV
NVDojMnamDW8VEBZfCcEGTvMqBj4sUGqXLRsidFh75eeMQOe+HiqpN0Of2IDmwOr
1+seoajIZ5zZLEJ8bq221eQreC95L83hd1L9+2DBUVSycI6gDIFLb414ZONK1vqA
ZLlDnLSnbJ1KFaD2JxExN8WJOMfPC7dvzNgRpGQ2GSRjcUSQ68+sw7o5DAkkVWFP
NNKNI3cQyPZaayYgnMggOyN5b47vh+0zDOr773Njasg+dUAnve/BPK6VjLkFlWUb
jQX/8RwgdRRn94lqrDH+0B+DVK3R38WNCnZtOW5Dtit5vo3jKgWrGKs9lAr6W40s
mKU+bxwmfxq5E59PqZj372hp48HWpmevLsUxqMa4KMPU370kyeNtA0hvLJYmL1Mk
2hmNIgQfcd0i1V8msoPgixDmSjSirm1xW5Yw8FuSTKJL0shjJ8v9XUO2kyNvIo80
BoLSWKc58dp58vPuhp5/yF4kJKuhf6FLJdzQun5vPP2J8PmCsAz9w64YLOzmCLTo
2oFKAcnfxAi6w3mwIGp4UNHMBvk7zSnKo8Rdk3NADXr8rpLsLZixnqkQnhFGvqV5
BjmPwKG8E+mtQscwYHHtypfc4sobu5fsUkwiM6xZkY18Bz0HoqhTj3T+mJ4M0fnJ
HuyItVntw24yYld7q8uwCV/9ufqbN+Mh/ytUOPoZ/xSCLcppmPIMErAkNsH665Og
WI9a6e8UVO0r9enFoYGNvVO9mpPw0ttVjPXlVqQgZkKcefHYjSUOmLcFRz2ShV/H
r+mjMl+l/I3jUn/l9sGzHvE3VRlZpDdbcGpBuF/v3KlYKpLhqaxU+hV/cKEKHMld
finpSqKUvqtpuwQ9DMUn0MBj8RLR4v03ZKB9gFlxWkToyp3I2/WIwS7wBJn2/gZc
kqI8xDDhQs9KaPs6JjJSabviijFP8erFHu3vkaUcuFNCiTWD87jA0yJMNduD6hHX
SOOA95natX1JwLZe3VFspBvLbJGW5rKi+P3QsTiqacHhIGBpURq09tcUUoEBJUTu
hy/OlUvpYV9xL/n1AAOZ29E1SW5hHmUFywmbjUXPG3bqXeIkhWys0Qgl5BnY8mpE
2tl0zh/dcJFpxA0845Hr7hx9enhEydHMlz9pb3cwj/tTYxIv704TVbLnB+jgSvsu
hxnyZfO6rlynJRCFchBtD7ZYdN3FNqHl3ijDoftj6LxOrBPB/9FOVXdtVWdGyf21
965AJwHnYRqqUWPGD4lGW80mkyQfJLXx8GnaBEF7rZNH/QpU0ekGb8oO0ew0OZrW
AGLyXYR0YoSdnCADnvzB/xNAl3JtusxOqLXruVv571Fg1WxiCV0EJOvVcubU4zcA
TUnHLvTMRLq6olvyI9/3KDDB8XZ8bwlpBui7zzqJqXAVEqggnWyWCTmi1QIWAS8x
zc3uCR54KpkbMVfZlRAYHOlr7Pri+5xWzVgzJM9zyv1pJQM2sn7soyQMqn4tb+BQ
B4RhOAUS4+kfh+3P+tmVN6yorR2HlJobk9l/T9PK6VFiJD3KtL6gdD8YlBtAp/vB
/ID4gMpVnWsuXyeARpIskaWDGFBh5rmT3nsWfLVlwPODoLzIKA8rVyp39gNKfcNZ
eOqlJueQy+BLfn/g81iXynKVDTbU9Z+cUkP8gDY01uz2rMrP2ovbZZ0x4i1Xy/AL
QvnQhSiJfkp4t8/l811YAIbkp9RHNR73Hqdk1DWpkc+YyR80Uw0Qrf0zT1LDUzDm
6naJafbrXwXXVAhGH36j1J9TwkwuAAqB9iaAm6RJes4k6LtI0yc3Zp3gOf2j6sOe
Q7AKfcjErxRcKy9bZu4U+StdbIcQ3xnpXC9FTFJA5ySCUilyqtwKIpPKA3N/XuKa
hAEESXzi5UKd9+uFpOVsCHuOSWVwlD3CFAPgLOE+qPL1P+L2p+6a77UxKc72UrDN
Xy5qBOwoV8x95DoALWEh9rLXillpJuMrRjvRuPpyBbXOECF6viQd0z75pZl/PvAK
T5AQbeYXSWs0jLMmS2Y4itA/K03Vd9RpM2RWNJ6A4gc45TUDU/lQLsOEz2YZruNF
GX0XHVUZ5UTkN8fAJY5tgMSrl2gPaoiIJyqQM1zLcATRcDRoCBIw+RJNYxN6Rmgy
GsHhzo6qBOkRFieQZOsquhRxkO0e7JXtLI2PgH60t9mfpiBh4QKJ+PGmLAGYkoA2
Xd5C7SFWmIcZZ0tPoVh0LzlpDP4NPZuLVqMBnRVxkvNvEYfQjZOv8UsiLpe1WV+8
Ck93ZGfRBmdaw/xbGCSAJc7Fco1Mto0eY93ydC50Gh9OFmYjVVVMES5gh4nh5bpZ
io6JaOGxNGat8XYboaZrsUrySESLMUblueIzjD0t2PlUP1kJdbXLjPUOBOTvL4sq
rjKLfGK9j8xpTpstTEoQ1ciRdnoqmmCezLRhObD4kc+obcCm9zE5cE7zfxygoP2t
Df1XPmFsr8GdQSIKJSAtnLGclv1+MZ7m1oVxXNskPaUeA6+mG89Z7iA/gW0rJI3p
3GX6bTqBTwQbtRBQD1vNaeMiMwle4/h3AwbhmfSMQSaDhQ5VIaFwsZ8ahb0v3uww
zetSN+2AzAGzg3VuNorZkrZFoa3j5whgMcAfJ8sxsVT00vUZN2vVO6ObFj9C3+h1
BedRp/eT2La4Ap/5pKdXE38dtig8NlrKAyZ6tNXj1HjHYiFEw7P//KUX3KaTNa1E
mHnjFwjUcbSjcfWa4deIcM8WFydQcgvQTIvb+P63t/Arw2eme0ShxwagUfC3AQtF
y3i8Y5U83TAiUP2uoQ8EMwXNTdYYl1tWWtO5YSN078sXcm7Rvvoc9LfPYpTJ3yGF
v3KB5p9qTTGS/Pz9YVTcWeaelU/dM+W1RkXFETi/A9ob6aNgo/OW6Xhr+QHXWhRV
L/GZX7+yMVSPLF36ZjOzPIF+3osDuAV+4pcnJa3BKatHNIV17WbRFN/45uPMA2eu
Wb6xOpDUmU3ivdbD7fg1J79RgSIt5MCamcnY4vuC8JWQuuOIlWt1qQzGGaOGCH/Q
Y1ImQnVb+WiIWVwxhSiTCNT+R+7WAVYD6YUx+g2f4B0aWRP4Ngq3PBEki+BlJm6I
SkqV5ibabYEScXEz6GP9eT7xZafdTAZUSecgpecCIbo+ZBnHSOh9Q+L1gmiBZSjv
IlduJ/GONDgksgUgyQtk2HY3FIfFvauxM68AF1LHuiJYJ+NHERQWNUpdpFeNbLp7
Qb8jL9y/2EgVYP7Fy3s9OHkal/KI1wEIAx5iJk7ONNrt5bdnHYKhKoGU4HIgijDI
KqJ/d5rOhhV3+zLZtCE8NI4JNyJYgy5vRkyGQu4CmDATrmAziB/lNo9bPLd/ndys
AnZzL0n6xLgX7sFgUYe/B/3ZCHh+qxXp7uCsxvLMNNSlfgsTTmTbF0iR5lAzY3Xq
k9Nz4/ykvSQBlT6bGCiS6omIdqRT6OfhqkDQaouZjXVsHQBAIdt/ZInpCWmQUNzM
dJaK87PfABMG9Q50VJ+jWj0wsspYbhd/valavgynQfMz4TeVWKyLmCzlJPkkOLu6
yPdAqHkvhGcugXqN5WgGlIJv0I8e3BhND73hDCrW6mvfZLZm5xzW2QBh596qJUuM
sGSmJgw0pu0AWjNo+3w3gF59Y5etRFEgcXDLY1oQepUFlzqLJKcOZZ4zzBlo+3OV
+uJqe6MshN5CZYroiWRcZFN2jyxX8VIomwfCkJwVDnwyqR90i//8cbLKDpMMHcBk
tKYBTKTKTNz9ex5s+tSDSRvR8d9BJyiSgcp/BX8y7XBvXT88BzPxLxs2oW1DIrT7
Sh5xNHAognRIP1QAq9XYftr/Sndmw6OGgRP2jeZbDKNeiMwl9sNdrlFz4ENBtMMm
LBxNR4JJPpTfkl1Fg+IGdWrnYflb3LuILpWs4PwWm8/V3b8Rnej9scGrPGGPCDSH
EgzdIn2X52E9kgVJhBF4Vh3YRjofcvl4EHd0z5Q6mr4gDuzqj/ZU7b1GzwfeNLn3
USGH8hVhyPZidni//+mK4g3nF9A8LYAT8Vl/BEZn6Zt3j3ve1sSohST3qIBvo+KY
dRLyCHDfqKruLaZ4bXiyuQYEKNgQk8w9DX1raK6ElxnkZgX2TPqWAt6clZiABa3q
gcG+4s472uY+CebGAo6iRBNr31w1GrW0xFXJH23V8vHDqQEK4NcRfX8kA6QPzySr
DXXeIgGq8KMKj2MtOnz/xF3bL/Gi6qCNjZbGyVYrjsaIZzErsqBzZAjv6sFYMNOt
Ze450replufqFkvHldu8WZ4ELhC3AwgpzuqnWi2bcPscE/ptLx2dHRD7nYMmFfxy
EEFzTrMn1GwQxyfHiQEUYL0CV/iwSjloArMVZTYxpgpBputXJhzyF3upjDAl49VY
MSIiBnyXKmp/2VxBTt+3dpaNA3zzNdTd1QBtyfMSkoBStdFARWdndQXNI0CUn33/
ljLQ++pi82AWyAqpK7nUrd8D7/BZNiMyMNa6ZoUR1h8n8Ri99AwRfWbOaY68b3fb
wGfQQeS8dt6ot2N0UcDLj6UgPmcKmz9CtJx2NMCGH0ve4KlIGdCj4ZaMTnxV6Ro5
BlMfX63Qtf7viaf5efuCBLajjO7HOb4NRWZqEJgtag2N3ZDnVrvlAnVvJbONyLP3
QbxxZk7g0OwFIVPBa941p0wJJuB5+8as0C3CXrWb8vfcOzBsjJDFk5l0ohBCs0JI
2GVFR9R5g7phCQQ/WTI8yaqZUBcczQFlY3cXAoQSL+mGFb+HiYii6DPU0gUuikKv
lSeOlNUjOZV4LpGIcyIMKaaL9ee8npa29ML/2fVZX0CBXIUZVRWu9SvqCVMZg+Fq
MI9gZbuYiu08yFHKPa/6QnWGmAJ9zOmzCM0vs5vW2p6dRBs048i1SWKVQbIXoHSH
oy5AoQR/ArARyRvkxG6Z9wEG/v65N+UdBMVYVwJviLUVqcta+NmafmEd+f9CHoaq
gn+uiXmowptv1eKaDcgcikAUnT2pKc0fQY1OgLHFeKdCPdU1Pj2PE/upnhFW+Azx
awt9gzbw9MDbCoGkpYCus2bb9pJGUSDFFyr9QE84cH0rfDtKSUhOEZuwCJUlffEt
DQ0zvVjsLxv8kipNy3F/fpNWZqdXaZHlSFQU7aTxkd+AC+D9vlGBXRjpkMt7ndHU
8jRCyG5VuV3biM+lrzDFilZ6W4Wpp+Kg+xaDod4/QmC75pAnTu5vc3saraG5gVrC
woo+WkfGLPqoAd/Fwtp7VQADAmvztnQBup4GtbYZVuLno77sjzzmtWylSV4VELdZ
bYEXeb40Xh0lBej37kQJoRjnYn6VyyyKc7fLPnXnhCWskBOsoLnDZ0xbwDOEulY9
WBaaqwQcWl4I6r78SZrFd5mKA4C4ywEFn0isJx/k+05+WPV9vw9giL1l5i/QPjZ0
gYiNRN/59WGtEHGRLtg/pA31m0aosOSbSzCRTU/2XlJwoqtQFYlaz3vOoeXgXiSu
4Q+ALL3E5jsbkRs+ZmGEAxSElEkgI0lWA7/SCodZIE5NiffKjSSCgA3kZxF2OK8S
5sxILj2MHUys5jpCXOuaVBfU4Y8ve4T5mW17LBXwEyGmkYFIaSoq82adHzIZj2UJ
eriQ9ZJ2Y3xTZZD/1cxvuF9cgx7NeiCTpc+AtlH45GJWV+vbV+8xoD9gx/mlmY/O
zeHi36zKKjpIzQqFmBa5btRDFMQatc8jCkGJb7EwZ7SQMvvbhQZu8Y639FFNh8eP
vN8D8/jKvMY4kX4XEs3pDT0hssJGNCPEuT6ZHT8rsDhZx9cjGY/vRTqG/Kzd09da
3RNSALJwwgunLbl41qc0sImoF29XSG52MOilu0EDoA4b60LdGVCmyovCvbktLxfw
6YS9xdtm3W8e0owNyJeMUDLbguaQkrHjCAlmjoX0MhkmAzLjWAnGywz0ZB+I4TxR
HgZXgV+7SoHJ17SyT7pGZHGelshYHBwkDNnWf5Rki1piKMV/bbNKYQLmYFYRVjPH
FywQyPWX8octeFLM5pwiN3gQ3/vQhkSCvSY5uCXYlAlXY1MCwZMDGdutbIVvmcT+
8LXt/byZ7Ot8RMjYMSYFHtGNvnnxJYTxM1X8IU7Sa4ho6TG/FrWiN0gBNY1dEy+g
r1OXMZQt9+pAmmaI4V+6CcF3a3SsZ2312y7o+hBMmQEQTrrhimZSr17W6WShaJx7
RZ7vE5q2jRqOs8295JsXwAJZZKzVbJoB46EeMo+eUxoBEpZ0WseMU3kED5yPSLoC
v56uhMeDoaKJC4bRgiaCoDCOAOklrtuhrOY0s/qqeDlstUA8lS90B/5a5pWjpcj3
JWnZibMUHCen4zBnPeKBgu0WisaRs8wG0KWYp/RGEZREz4tYCZL0CJVQSqAjoGvB
H30sdsiCn+gTsc+mQuYXCPEWGlk6hcWYeq4jgRhBw/AuO94TOMEjEBcfw+uwve34
vLwPJHU/4a6VtJKcMKb5eF8EJ5OjVLfg4r0r/CRfCkg+0DAv7DrqpL6TsQNDuJH+
BWnMhJRcMDv3bWMRdQBVvzea+tmE1zV50Sa+ZLRDDi6dyQpiN1sE6dVJJmEE3aNK
VgSACTX9Bv3MJndKlE/AgAV8zjHmZ4LCbRzlBqlN4yOuJbMwSv8tyaJhkp2cRKDF
RmWhOQvcORX2fwwoR2CaZCOQvQPy1c1nuE8uemBvbLXa4UIo7dFVBgXLNaQGpeRP
J43ugsbFs8VpIzS/ZzB0FwLaMjcNH7BoaUvvSpIbtqCtE70CerLO5d/NJtz5LScR
pVkQnEnLTbONuE172AP0Ra3baAb6i/BSuHmvZ8u4fXgJ1sEte0em1Jav9no0txqC
zkOJ7oNNvRvBUvZuikukgwElf8lj7pFsoz8q3uvuBb158gwc6abW/FohCrDTIdO8
6CoURTCO5hFZ7z+7mGLb4ysZaZW7VrlOLpOlOqkiSgtjDunc6z8oBQ14uqH9phz5
fUWPVSjM6uM8cuDkPu37hSxHQcux/ejHqxtws7b4DQilbWSewei3IGN4OowyKWXI
tD8kwwyFlh6L65WngRxSRemfchtxm0E+hFuXE38CetCo+bKPXHsbJQwPkfVhb3KW
WZJLuPTIXPAPhlEE5kA5ZeeEWUYQ2TGn47ns/RWYdulX0dzhVrGs/lkq27+hir9V
4lFWRYwUgfM7WV3VuKoT3aHPD/nI1d9s3x/G4BTfJEVOaA2SxStRoiMlD7sk+9L/
LnV8FTvR5wJbpO1zYEUi7TeLvHFPHJ7bxJTpioJrYERfHB/8eWo9y9dQFSR1I5TB
/YHQZEeAbr8noeeoljdnJEMJ2S8a9p3ZjZjt1WcxmTYRwm98V1PpKt3kbJX7bFBC
TATkYPP3VudZx2WFTRsF6acEspR+vjXVlX1YqUJ7VyJFmrbPdRPPUU4lDo+WBs3i
c/qMtPBu7io09knS0rH7UO71SII/S0akzQz0wtLZEI5dN+kYamOGa845EjFTTPKR
0HrBGRN5Mv7+gK6DFLsWjJ711lfoN/WLgDBSPjg7sTfTGslKgiFkPzdlMILQyQwf
JbjqXoFwA3CconILnQA1r1vn4OGD62J5lhb+w+qtCpN093Gqze4No3YEIfouhadW
PHN9iZhtVNSVLVtKmYwTQ6guhjX2l4uAOZnaEK1yq4hEwBCAlTvHp0PCCnuQAjT5
Ul2CQQyCaAPY4UfL4BU/VKIZZQNCSoujAlVaOps/wfPfsak1Yf0H0JFKGwlJLfRb
5cbvIO7EJnO2virXuJ8kCfJJbVQEy7oya/0IxhM042j86TkXF4cBAejwf8zlGOpq
67vWQ0ldJCBfESsF8AOP04pZ5WdRTr7Ep3g4egJOMbDTkDbxa3vOcYHcFpWeeuNX
boswrM4Cn/reJHkEpFPwuY3CPOf/5hKTgAxw8ThCLpG7PoZBTK1oT1Z/uMbdgh9l
fxNzGlUKn0S7CR6yebPI2nhOkTAPkBXVzrgc+vlEzbCOJ6ykJ1pjrqRze7Hb8p9c
1K+j7ht/ZRL0MYXYXEk4tXk+1NcT0UpAalUs5WKqPL7UYuu1wCRSBUAQSLiLU6a3
JsQZAI2zBbVgrB2wQTHcdUz+nZEwS1oFqv+t8TFYl4OkS+6coZRKC3PFjUBIrvEI
Yvwn7txtlQXoznh5i8OPLjs16LYekd15RGse9FAbv61rwyayIStlTRqhT9d657IL
W410B8gTTF0dovYcRFwxUmXcLOAjFZRD3diZ61xangpIFcw1XhlzPMNaIDk+IcpE
JBO/yMkY733E1+AAyoqyTWElRD+jTJuPmsmHu404QQMnP54k0gbhCoJGvSIKotgG
cLALkKLIl99wujv3f7cqNeezf9JVQfrQjzEUi4ugsicPNmyyxSJrAiaFl/oK2b5h
eBWwThlobGRSNdEkbw50+F4e2y1KfES1y2PoPVldSSmJyxhMHomWna/adF1DahXi
bv00J4OuMYyGwtsPA2TrYlS1W6NtrExy9fNh2Vg6sdOB6hpkEMOKxiVa31ZqJIlW
tDejKzguu6YkKdOHnS2swGoFdfGnFE6l7K4d06zeuXtuuf/DmdIDq4YPLKZQcXsM
eQBUKTXiIeoY2Q8AS6z7VSFLi/v2Lg5zmf52ePwut4dp+O9oye4JYDutkxFpTrHq
8lvqGoRZWGo5baDs7R5xy6gOX5rQRiAHUJhilNvUTSG6gAworpH99oy7wxHMW0Oc
dj/3JpjhHhDmYiyuxY3gBSJgn7FNRp4JjJe3j0LmPaHJFm38h72zgV4479lpANSc
ClZ8sq41sPAa7/PrR4z2hN0mtLE0vy4NqFgPMd3ig/92Sn9aqAtIdYASGMPJMdKF
o8o6C+KnCvUPtmQ+f2IpeBDL07B63uiMq7sSgz1u85vwsWjOCJfF5b8qxIXwyf/Z
HcttWMIKkWSSJuZd42Fh28hogbImANPdB2HrIiX6q0pa1KOgge7Qs7lQcfSYXHmo
JWv4Msm4Yg6Thv6FzV6MLNZXbs3JYniwKn6H1htYxB446zXPeKG37INw/V7cey6n
TiafBglv0bDVchVqldGi8MAw4KI12ekhKnVMW+7Pgn3Vf+WsLanUogXfZ7ub2fcP
k9sczDi6x8ngZMY/v91WP6PdIGnZqj/gBHdgSDcWOcLtzc4T99eNIeuxOx3Kpp2F
ULrnersgUEBbUnYZLXx4+5jhWyLnHhBKJzPxDTKekPyidMSjyoWYluo2YxABheCD
gCHCikpQ30r8Rcm0T9eqQvP99qIScZ4R5zECHYRh9ku/FP7N+FlGqzG+M4UuZmyY
X9pu4NSxPgmMTav3zmKj+CshbEp2In2C0h97otRp47Perxz+JSn4xDnx+NeEBZla
ARtzThSGGFCLH06GZNoGai5HtqNzVxSx/4Xgk8my8gCqyJsz3PXlwLIE9vKVs42Q
sUCMS/RRxqNUJWXwKU+EBLn284XarXkfetdVebzRe8O+b8rBFGNI4f0e8klTgxDW
mIwezZr6RXsFHiGeHLNReZm/pFotoZJT3ftRIFkL3cwxHn7JP6g5M9gV0pUNaUSk
hmb2fwyAzI7QQ1pMWfw8F81ViLUXFYQ9L3W7sEHeDw39Nyxu4i6cotu+zgmqUEjg
U6Sunf18FKCn+Vm5d+F9E0EQcsEgJvKMP68Mi98w0maARB0gBRelspWBDnNZAsqi
g9DhsTRb+4CH+yxex7TWpe18Sx3LBy6Z3sVlUPXvMiM4pgmgY75TI9bCwnCPeMMw
xm1Me1LTSVQu4p6dcnMir5wQpKWC60fYWLDaHYRIqit7FSbyYhZzQj4xYpgiOuSU
USO9lwHyplYGRS8ZVRFFsinaRZ0QbFVKvwlr9IhLKBFDh6t9dVdUeWpru5t7bwjo
5yUZqqsGe/2rndze81CGN2M+GGfsaGOBbOvXXPkMMXjPw+YmEffV7Y95QWb7JQ6Z
f7k5LRFHdQowBSm1feAt4V0IEp3o3E7VxfVupMh1ehV00LAWQJhlpdMoSrSKJG+/
pIT3jxb0Tp+GFk1r4Vh09EmuYofTF1AFmdxAh8xnr0gqzEvnxi+47O/GxE63G/P5
5/Cg8EvXIVPctKc8u2ZpXKChvPlGMnnjxwPQbxTeY3SyGJuHKZxezdWSZ+T7LZg1
tMSBjwY/bhEX4ozhq5IfzYqYdkNbxMnxk9V+9HmrnT2u7jYbpLpZBe/ZRh9hpiSv
KDcaTcnAJBo/UF3PPgKW47Tmu5+Y4I+ldPTDSvYn0d98D2LpWc3/D2Xt6dZ7I274
9Cdjf2ehj2WkJ4vO4ezBN+/Ie4sstTaRqJHkQemM7Aqv5jsTAQLwUZlL5q6Y8loq
O9/9V4muX3TZTe5bjdRRUrb1RPBlYAJ/1grwvJQG2MlBQLyqA0yNuz0hBD2o9lhn
Oo/v2KsePWD9Zlo9kZZR1+k1hzqflMcREqdnUrsJWUNmdaEvoIi4C/cIFXhXGgG1
qWomBCpGa6MuL0qwh69Zc2D4D+NkohYwK907IUyuw3lotOj5Hn2GIU1y0jxX6oTv
Kn/BPxImwhNQu9Z2d8hH09xJlJwjzvsvaSo5f9GkpFSerWibhGtLiOVePTVhpILP
j1jKK2/3e/aSZ8eZvIQrAZVpZ060lM7ZPWwTTiHtLaTmX7JUslbX8TJzAdcM+LsY
eI8/QlcsjKMxFUih8mkvbjuqDkV+eDdJ1F6w+yI0RHRJoaJo19PzxyFy7KqxOnb3
aWlWnZEdMQKWoYOVMsbhy/N87hXbZnMUJznylIf8ZBDp0vXz5QeZ3BlBb6MkBZhb
N+7AmcEtraA6RTUbXMY9yb0LPiDpUZ5iFOTYRcKRhnYSMbrm+CSdR0FPQ4BV/pQ8
UWEWoURY4Kx4z4i0EJ5Zn/3VG9hqo8GdBMqZ+Hs9LuT1vm3WwaSKsRRt5/yvDBr+
q8xmSmhi7B4vxfP/TlSX59cPhIV3cOgqiZg0+oKzg8/nZnZoDV8kLPAbkgA+M09Q
QMoHWzeuMuX7k6OpqDR/dR91sO+jEJXGnZ5eg4cFEIqbxswqOFC6R4mOOV8iDF7c
fj3Ka5ij3rcstfSlNDdBrivIytwAoMgGAS5zEWkcDiDV1W2D6PxZnFcrIZ0ET3lb
FCLC1CP6FAsJT3BdFdjHQD2sj+7q91bjvQCi1HPBB1SJhmf2AAbFQLSZcZw2B8Sw
bDWbZ8rYBN3JgENwCBSaMHtl+T6Xm9Wfd5JgVXN0P5IMHrFEqAnCT3DN8CQNCS+3
NAwSFIgWwkJwY2shGr5a5z53uTRkUKIkV+o0MnR3cEDNMnX8Lii6c/3XgiytGx3m
PcNhp1iAeY6wJQgiz/40Ww21Q1sWdRC1MxJe9a3vBZQLiePBArEGlLTrNrMZ7a93
3i95I2AmlnPe35GNxrdnaz+1/GV2dTxbeXXlKPiooNAXwGIrhfyXafhENXeNWbFN
jl4A++1UaIeM/VL5LPuWDxPsIbRl/6tAPADp/WvCl4tP/seDbIlHL6wUxB+uPUCW
HUur6QSXtMiOAuWC65COmwSfm1UgfiJ40BpJs0H6N+6s8AobylDR60CgZcr9Zb7R
4lBrMdj7Mdmzl+/jX2AwLY0kodj9w3W4eQ6v12DbK4zTM22MzAK/x2seOm4OwRFB
PEsp7T5UXIpzNgl6Ql6iWeB+namwrJB8WtZodEZaBwOqLhDvajnGAP2946utPMwl
nc+Atz3szyoLQlzebVAeaTwr3Wkf3Lt4gUyo6D7AkUrjVExRWKtTSoMaeT5pT5+y
hl9TFnEgw6JjkxPwVL2DCrfirIEL2us4cweZntFXg8H9cFlq7geRzewm+w7ux87H
qJZ0fCr6/t4EthJsztiZFM2BcOKVw/+sNLaV7PLRS/pmhTec541NX0OicA7lwOBq
lEA3fdha6Z9wi0GdjnmJ8OE9j/b74HmVHsWpo+K1sYHLRteMj6bsyGGT4L08gV71
FNchgAcFKNa0HAEmjz2+EZIF9JjNP99Gd8OVyd7tX/Whpuvj7HpCssWD3owv5XSj
TLb4grbajjSXtQGP8Xc7JpbNw6wsu74BuuQZAzks24BBrYt6TrsRynG+rwbCMP4C
+lsbf1KBnOgUCDnKwgoYYaMRkzGlN794jyNO+4+E4U+io2rvpStDxkrv4AHlInZZ
vTE9EsunmfkpqX/Ot/e19cQw9R3G2z+LDhVRU2onjG+ortxz9OVW870rcTPmHJXZ
9YBmbn2tSh4IWZP2vDE1JD/S/7N9Xh1PtPaLnOsbd91ouyD8NKvblIieLZfuMYX/
1xkcwWzqVjUnF5Kx82WwmZ+lZYkcWyLfYvzWVixwr5NqrmoJXUGfeoZyJMLKTC7G
Oeu8dsGDeNI1a0E/1ZNSQfKFlh9NGp5SPUBsekfJmFcjrKdiC5ZK4Cbi08PBEaxP
2CZcRnoUR01nlHi3xIKU8k/EsvJVJbrgU2E2lfZ11e2la+TkWiJ2n/LRFhEflY3g
Fi6fEzpQ4tLhNoghGbkPsAVcZ4ZTzLdJ+4Ftgppw9aVTokwTI+ctPmz31Eu8mzDh
Y4vvmqrSK35zO9LltYusgcX3L3Z6RGsKAbL5D9dcWzu28xcW8j1bp3z03Vd/LhcT
3FbEZmoJn1xp8B1uNAHTu0OiPfEWT6T/bx90NalY4jHatGZipTTuRZaQPytSnutm
DBOWb0kxlOq1E0PlNSkmXLIrx2eZUO+Dod/0+kleK+xJZX9iXctcpSWrhZe0aMph
QBZDjYlPKtdU+uoFgQrx0jDigOtkdrP7JcQiApoUkqisaDeLjfBfSvyeUdOIEqSO
w8Q8MTKxYmUUdLXdRnAeuNJuys/PozOhQSVEp08x996gdcQdvjv5GLQBTLwa1WVd
8Ysl94cBZBlBvRE2JHtZ5ZdHRDBwGs7sxGGAQuCuJE7+xBSZzj4br7jdTBzvKHYv
6OHVhvAMz+H6Fc7JpUGw5mBq6Yzr/AqPEc9GQCgxV26mrgQxR8npjA/8suMO3H2p
gHonSczDLo8TVoKKybz7bp6R7d1Wv8ldIrScKPBkwZOkww2KyNWXSAq02M0mgeiv
+cKPzK+6wp32sbdrIg5I1TRa4MNgy0ZARWpDTMnx9SmhoPpE3m0IEvZvgEXDFrWP
4dYV7IOAA5kShh8MwhldqkBzQ5Wbya5Urqg2VNF5TiNcZ2qbdU0MbGT5IIFSQEnK
W5U1eR069hUgkH17YZa5piCvjai1ZdZbWQ9+/wCrG4ww3s3cKGZ2HfLM68RWMsp/
agiRQ8fOch9Jt/le0JvdewVq/fIyQ6cGq+6LIfxbuHFlnF7cBV1ki9pc0KVoAEU/
s2JvZQffOPSKUq42pZFZvzVTFEyQCHxOXHDHGrLIU0YyeER6rID4RHbbofhOiU3p
UkZ2qM9fFD460NPE+CCxdSyiq/SfqKw0HZuZxGT2DbevdxM2sTRLapNdP8Ye7jkz
cuIr/MDW58Hv6TYxvmeBat9sDlC0RFcky/gN7E4VKiIisTqyW6oKbhGFzvyZW2g0
0BVSqO1kNaBI9e/itJxLlrOa7iapuQvoitRjwkxTNA3mbSBj2jyHZ804aNH5nAbW
RoPo07rdTIYS3lLszRDhRHcXlHaiw1eugUMCntbEY5mrlq0J14wpV/zjSI8T3o1W
DofPAlByTGMh1bCCYJfvUMOqnk7SQZkwxQqbay823gWc4PzpOr/8OiDZVmruzP7w
36UUEp62f5T837WOa51zQfCfKKHQruphMO3k6Vd5TY9TIpxBzDYQxeROn5OhchCR
xkz3jmz/eR93oXHicQV7lquUAUvGPHLZj8JzW6v3JuJk6/7vK6QW/MjFJlxE265I
ys3vqO+j/etvIUgoDBq1RWpFXfFxjdm4bAHseDd83uJi+24OoywC3c2xG0hJA2C7
6ZvKNvv5U0nB9zls/VaBaHid1rlRe2jj4AE4HkRnkYgN9fpo3ccn+cfKchawWzk6
mR2jZ9r0HD0trpXwGyc2raDmf0V2mQJ3xqw1GSKrty+W+xd5/guBIZwi1nzHpP7b
VlGggG7yMdTS2L1Wy7fihuuVBjs3s3nGu/D/xhpndG4Lqn+mV3jNCpQ6R2SFV74k
TflzN2UUkOwZcY84quZNgw/12oRmEuNNN5VU1dXupKgx6eY6b1QDQCDMX9VpKC8U
pSxAus8M8wd7k3/yjhonhr/zfYwL+LdTRaTAB9eaoTp3Vq+a21Lue8q/hgotNVZ/
I7GaO+bHj21BXLElhLwN2WSfUzkQshIQqtjdQTZ0A7qbxarK6dGLmWhiul3sReiI
Bzz5vnL/6sqhaqJiTgX8XJETrhji8sx9x9PdXXeP3BD/Y3dQRt5eZpe+K5ljII07
IpS3s1/mHKXqmHnrhEWSqgSmjxmryyLLcffkK3ywxXqsJVgnu/n3W9IkIjZZnZTN
kSdhq7VEfTssG9nyFDWz1Ff2BNezoVI6eb3TsaonXQwaGfH4q44FZKzKLaWK7Xji
soMxNUJz1l7DTx9O4saiFoDDoKoq2gk55TduczPCw1GvcjCBUvVsw3ii8Rtd8DJ5
Qtvwe96JpCDoTOeSsPBDkQ4fLv7prcF3BrV27KlMGxaeYfMwanc2IhbLf1x1SR2p
T5p5+29ACwcUamLHuen/K0p6zJYD5VUZ5HVMvfBMb867Z8DETpLiWqRZtL0CGtKa
7sqg8aZ5Gyp3+WhFC+ARrbDQTTybdPUU49L+HlbjdwiMHVx3+wL/lwCvVjlGv3rE
dWpR6cy2wiRDIYnIS/tVjzH1um5jtxdnlZyL9EvfUJsYzDhw6aeoDoENRxZQX5A6
FegxDWel5rBDSIidhSKvg25hz10FPjWqpEuOYlCN4Yqm/kEjp1Rmw1KJI9Ro6xJu
SMFHuS9QZ3zKrRIzhb03ezpNeIvIpTz/3ceheI7Ed831m1abjWf7unmZpAZ/xOEi
vb+CJKtEnB8mdKdHDPzIkjWD8YMZ446r5FfKDJ9PF+ZBTLcDBX0DVT4+tu6KehgK
bRxVbRXoxFHabXLBJYFldXkeSedEWpPosIcv9ZHSQLnIc6zQsHJkPRpCuQ6458NA
ya3T0bVaQfpIO1ow1qcbRaTJOvXd3t5Ke8FQfU98es1x32U70xaV1t4FRA03O/6r
hSKVW8CamT1oyOxY4uWpKtMA5MDz4x/6GWJ7xlOPFBKEKBj9+lDtlzVk6FDCbjvz
aaAs9/6hziBe0H5eLTbKtAH2fbbFhuW5oX3IgIXyiK0vtlP+ZCEDXfzO1CEp7bMV
Bj+Xti4dQI+VP0axM2cEtalUD8EuwYbcbXNvJlYyxiSZcdSrO8eWlFe866YcnOVf
QL8jGFx5K5nVPu8tTWtCgvUF20F3cE3vUCc/wXuvdwlPt5fa3/FSJ/U4yFIQYfgv
zzH+5VeXuEOYtBoz+8z02WBY2Px9fEsE8MWYE+baOm/kDa7Pb8l/ys/NVtOqD6iX
Qk3JkmuqZrwEivpCa7yW5sPQ8wLLFKzjWYRnHDKq8+Qz1qrBObqcfSV+bJi9QxiA
51Ax96XCNnjn6f33FxFcnGQdkITmhFyBYJfCRfCGW3nLlNzgqeN+6ExqRJ6l7vve
Mjzwcgee788FoKcvO9yFpqY9gMJ1aDNZiBqnZ1xdhXsSb2ytu/fAmhilfij7domZ
SP4n9PKmSksESD8wBSsAFA4WnLxkZ+IwD5kqc7k7451CMVdnUzIfk3DsyNCzJz47
dIz4PnFPhxqEVLvuIKKhxzlnZS70JNYGc5zPAWGwrdruM/fBO+cpKABsixc7MLye
NUyByY4X76rkFXUWk31+z6h8eeWVVwHR2QG6h8i9VDxqH0FMYEPs2fWyIm0j8iWP
MYLbTcwcKHWT4a6Xsc+VnEweSYCOClZQbwkvReAmP1Telkea1I8cFqOnol3BOP1F
/7OQaukyNKhPbhJsm97/sN2smuowhlu0+IkkrrEMKHq+omBoNGMSbvBUUM7PmBzN
+a8yA5v//dcNncG5THzrjAGz3j265OSavNnOzDCgjAj5MRiE5mlc0/0nD84cB9pp
kmNcx4EsmdBdMGhpmTP3MNwAlwXr63yvfZd/LJitcq0uyvGAl0Kd83deYin9OpgI
0hwkYxtlmuGCZmPiorB5CPkT70+QB5syarEvNyLHBa2aW0kmeQUC6Bo6bw2urWrT
DWZU2g+S3zZTMFiHS/uoaqbkruqpmT3ptiWVm0oQBlOw2FONh4HBqfwRkqaQAcFK
mni/G49KVDYPqw55cYuY6EnVNsm9rOcatIQOyjBeQPqfZIm1NSVGa1/LOruKoN3a
R36N2+dQ6ZaFryCjlLW4pvFKt6CadaqZll7bYDVC3Z/+cK3YP87k/3bS1v9z2iLS
/D542GHigpC8hcWxGhkkGJDFoZIAf3pIUEo+EY5G2/sEUyeZUoTPZKrYPa4R9nhz
8pE0rY7V6ojA54ST58WUAgNRNtkYeLaMC+v6XEyIj6G285ROicCf06I1o9ozXD6i
kW2LQ+mm1lEL5S44A0fsAQvZ8M4i0orI7qaRF3o3mS36cXQzjJ2Y6sx3ljPE3uJ5
EiVY6UedrJ+6LJ0mhO8A8mcjN/kJseYoh7RC3QliOlpG/A+OAS/IRINwKY6SZcMV
53XnlFn+yp6T6U5xSUr90mhRJ3MKQncswT7YDLFWxqvjysQTK3uFGq3tPXeGdjOW
GyDA2SIFv4fB4OW2DLMG+WTu7hhTDX1JjdL9M6cBFPJzV7cZQe+uQnBpEZgnvad/
z3vsOVhE/kU9Ixdl9OG4qjWjKnZkNIjfdED7/wO2tGYKUDb5UFZ9gazUQufDifdq
atUy6LMzwHNWCqlz4pZkuKuzbCoeAbMMokeaKDcssf6XF2Onb38PHO1+uy/DKs5t
5IIheY1RsAurq6blJDgiddQELO126JOgebquWy/LmgBeOzCM5fUVlblEJcFfSK1s
DbziCh0beqJiM0txZI4QEuAf1x8l2zV5a6cp2g30jZgJA7TCB3RLknZmMQfVTCWp
skNYy/onqbIxkeTo6MNKsKa4/Ew9mUOlUi5qZ1xoHEy8PPR9lLCZtbbmoyNi/GcR
+XPAxKT105D8wTYMZ5X9M0KQZQw8/iZX7w6KNrjMTIm2OcZ3IogWkfiMtDCRDXtG
5L5hOas+fYtzIw38DY8zV7xMjH8jABNqFUC/5oExhHMC7q+72h0ugUj5VeWrJqD0
2x8Lxc0LobfyERv5GBFebypZPIqM+iIF2WWSEgkAG2/RgGzZigW0MRnPlLlnoQ01
Ib+m+dVDyDanx1YQgvBO4IAi07c1d8uGhJh7U7oPesU5iR/6Dsl0JXNU1ppsR6yi
7oExtXsAUBnLaqZBbr6UHkNDftp14dC4/xvW6mLxarQHyZBW6bOD+Nj7YhYaoZpQ
2NCYPv0eCcDHG6kzFvauVBcTplPjjjg+8KFeFpU9BTUXPOUCztZomseXBGXTFesl
yxqfV1ttWttFEpiN8734pwcxXFy2UQ+8fgmWXKlk9OKA2fatXJwCm/H22tFnE+5R
BPR7eDMNQE9jADdo349KYB22WCiBxIwgNL8bl75NZES/Oc4C6zaVbCGaHbsV1wq8
I4YQS/pDuNN6JjpnrGcOw/+lFAYbwA6fJuwTSibTkhdYzOCKseK3EoJbrqAiivGY
DsJfcojI3D1DswNzWrczntG7KWrDroIh6xARC/9V6QQ3aeSzAHBcFkQVhVsGYiBx
CAD/0bzIxZSHoGiQ/+tugXKmwJpJKr5yoGIcbp8JsYF4f/F3xeneSFSkGK9Mg9pP
ci3Y2odUWq6nykGEvzo/eRO44IZgUGkCbX3+BWXqfmjdr4422yaTok1xaFyP+NZ9
8Xwt1WJZ2RoEW9RJU99K6NeZUzAQqiWU5Z74AWecbrUvDUianUKTi9XJaA3A+m7m
OO16m2JHJguhB07x0eyvsWK3idNDxL6p7/Oa0AD4p5KdSkSQIaQjMQjMPi++91oa
3wWK9OXmEinbQvkg/EMknRsWGDfdYKHWhKOHY8YmTc/BoWWdvu+lENmUR6fKMpsB
Ccwcfevk0qjZ8HBdPwAuzLgKsxr2RI48WYROgLiJhBtHvjoYY0uXh5P3yqWFqNEK
kD0fxUDXPKO48CB69vrEVzU7xNsGQAiwZXh/uuR4VGWXAsNE4mIGfKaPZUPfnBMY
TKi+k3ykj46flDxbzjImSrdgCJBNjGhFMut06nJ3jRhcRIdNyIhglLST2yqFU7zr
oDm0L+WEYGtFilPRFVk164q7jzVJn7jMeDBljDMM2M9+gia8/IHDxUMbpN0iDp8E
ESeWhfrm6sDba9YtffoLA1HwoSLpuloIDAiIsCHU1L1fnUN0beNYy0Bh1a+EA0/A
4yHL+WY4LXJNoOMYPEJwI1fQHx+2TBbtN0hT/+Np8v6rap3HAdx0MRdDNI+SQI11
OxpWBVSz9KjeL50WP35peCnSxcqoplmPS8OUbH9v6SCg3D2OFc+AI3WqVR7GZ9YQ
kDymXrasz3vvp/mrrH9JD/rqliiuIyNaTtqY+O7RvMJoHiO7lWW/uQBRVlA21EDx
LbwNBJHPRnuUmuBCA6gFjqFUFY/o7ARH5i4jfPQdWpnhOQ7Lxw4NezZMbd9i12+Q
Ua9kX3iVpsxoffKADL4BlTK8eiZfETolktfR8VrMwTDslPGrkhRGHABbl5X00/AX
+Fy5vX6aIAxi2wSCRvHS28R3EuNxpiHVm01tTB2Yu63Km1XOPb8u2JTqXhg85r6x
xS+XunIDjLZyUc41rI3reSSjQ3PRO0VpLE2a2144ssDg38TBiG17ocMsgl9zrVe5
BmiLHYkQUSD4jnKd2Kp9LttzIwCsJIrZtUAGjErSXD3JrEdOoh0IMh6hh89O4Yxe
VE5NKUResI2WBDOksX1jfFOHgZi/c72FqYnzqZ0Xl88LVXKpwpsAKAnmfc71DN92
/4r0h2AWqyZrTCt7nnWYz6PbWHGRDtkxT5+YYbSCqRIvTC4sWum5SxprekNvDpvo
VrBXnOEGQ0q01x3ZHgSXwIuwFoE38szrof6912P9cqgJUoZjlxxKtrDllpkCeIh/
Uf2OIgHXY+fHOzCuVYF2fD5iZYwcrkQrf79oq6kWWcx0gxw+f8nNnpoUC8X/5xkO
/516QO+UUm18JBEoIr2ve6QsYwxLsp8wm8cC/0ICLge79fD/eHNA/Yf8kcDiiHiP
/By1TdiB2T3uX8kM/2Bvt6+wwsCfxPWkvbdSWu+RTnEY+jemTvLzJI1NNf7esbth
q0A7f3LOpmuSjExA05oOdQSvNfMkHYYXrEeYkTIl+qHm8u8YV8S/H8pimjyUlfCT
803/k9/fegeDI23lWaNgeXhjMFnC88zjfYNgPRKTA7IqbqnN/3sFGHve7s4SFqcV
B2s1TW3QVQDcaRgKZjWesWK9d3d5q8NiKouq799v7GnEJczD3Ltvirc/B3jLaVPo
4ZTsq8tZ27h1VVBI77TleG7L1VcqF0pFqekUk+r2T9MnP6ViYAUGN6Ekr1qwlaIj
EjXUH1lSOXCaffxdPhbI4ZpOagXRf22RWGnaSGXShxsvPwU9z1AkQwgxmxHWZV7B
3c7f8zEE9dewrE5IYe2XKyMLxUY70xvzdykVe/1QGJqZFvol1e8QYAKRzk1FoXvu
XAoOAdMz815ndLrZMFZ28Q7rUD6mmxytIQm6J0oZ6bKCP4ws1BGkebv2eW5QWHLF
kJSPxFx6ilnzOsDflZ/OxbzLP35bwd6Xx23Jr0xD9lk9oEzO0ZkZJk5Lic8OVVuu
y28NZ4T3n2n8QdwlXITjpjhV+6j1GNzeDEHlhIFhqdlexdnXBeZMJjWGon5D+8xP
HYU0Q8B2uRgn7fIzQyTHogSPvm7VoYNnEBLVoXkuO+LThk6RsL168CXpEdw6CXcy
QJqmO1yr8KemNKP4KzFx95YmgJuByNwkOO1SVWI2A/Be7iK8g0HV7ZyfYFCHheTs
Z8BiG3AjAB2/r0l/5EyQ9oJZzWr7fc7XPoYS9HO0NSEheT/jI8ofX/mSxvcq7Qnq
fv+rlyRBl/27SSQmDmUf2JaS4B7rpL6LjONLetxQhJBWdABm/yCP8sE6Bm+Nyqdj
zw0tvbgEmOCa9yplQS79WtBCHyQoXaeh10g6fUB5sS/c8lojzRpVAd8mca/BKHRg
aJGLN/NXE+eprERa4CQTmJG9NM4YcDH606zROs64/qZY3SbOw7FYWHAi8wMcqQn6
ZSXoE0e7kwqtI71SiNQ5ZCQVZ7gvQ7kSbsv3favER8xoDcaP9ACgHjX1vLxbieqE
qvvKsjhD6Rj6p9E8Of7aK1JwhaXvvOxs5+9q4FjB8nXN4E14ySWq5AIrbCPfC7NY
zMzwqavRwHE8y7GKH9ZaXFsXA1M6pKlhufNxZVjxKW4fmqz7tEl6arlP9cPeAFYv
9s3ms7jAA/9ggMVp4xCE/WBe3DzbMUcq3YcCPxBc6oeQnySGTtRa57YGlFVKC2ta
rd8Q09KwLyVle8bFG/Xs1Wc1X8NLop4hBj25c48lIZ2kba55r/Cjho5CW1BSsxEf
XetB6zR+RTFIMF6jcbPcGlqOd/8A3Yjfxxh4AknQvaF+vShibOfU6aBcYPeNZ8Zq
5ue5aMuD6LGxkXZW3SfoGcjhpkMWqt+PmciN7A1vwn8zpAKJOrzt2KjmA+HHtiiZ
L+i6HKvnsMQda9tBpQ9jpXQY+oKA58tlccXgTyErtaY4WKJildumqmRtIdAR8CFR
58m0v9Ood3VimFt5oqh8VwpOqAuq/437zBGxros/370Z9tyL/D9cYurBJvs5hq9I
e5ef4g7Vcn8TKr1rgLmn7XjNWsPKHgInfjZE8aSX98zQnorTQnspaVJfqcL4JVJF
L7e9MU/F7XYA3e4w8nQirlSPvgLLZcCPkv50XVKTlP4AlmUzI54Uh7l+KFFTyFaW
H/ekrEoW1dBnl1Rr8d8XrUnjd0ONsp1CA0TXxQ9KUvLKMWmUDURzyf8JX1udC0Ds
2H9K81lTQgtJLB7TNJwenTIW36p0Bkg8iWrDzpNsbgZvISNeAan43sXTFjvd++QN
djLsQPXhX4rF8mqDTpOkWuNVYH7r7CThgzSPdBd1n+jh1JcmF1MWaG2r8vYGMJtN
uCSHiRQmaSWGYXvbk4gxIX5whEf56QWLWjgqII9yv0GaEX1B0zTORw+RjdYXXz69
+e4CPQnV8itbe9G53hwsyNjDZOa2tW4xwkuf8u6uaz7v+mEc6QfctPbFVv+YSV06
O2ZmFXJd2EBk1jEESdK+GxZzEzY3u6m0Zm3heMi6h1ix65ylgfCpVmTqWwkM9ySB
06QXCWP/SmFHGFt0VvwQCFeGD4KzKKZt1Ie9aq7Emx3MKJ8Hp4VQHbwiZM2Bynza
O5XINApRk4Jl9xWLn81rK3wVKoEprjjj5ddQYsjQy+YdsSQ7LgWeueEEe4pY159E
Wuy4OcssHf/pjaR+j/m6IEFAc55CnNvJe3n3RWhX5fRRnNy27t6dgR3AGfi1zkaG
CWqR+YYOaD52Ign/wFkdf+W0ibuT3y3Vp5oWcgRuHJCnKkJdzRLNgrGNKTgB9Sxd
vRvShfKbQpbolijbPeKrKwL1AZpU5fpcHoCPDvTN08IGeGtk8wX1oy3SW2oZUxbT
6I+hNTs0WlAutx+wTGjM5BP959XLROwJjMujgV8Yk9zx4UiaZrNrvaFM+GXrFLNN
HgavFfwjb9YzJvLbIfd8Ibqq5I8Jy18MqubChN8K0QC3waoX5JTAcvmlRUVX+XQp
rhxquMj7wY70fCyCJdhszywgXfuFMTpJ8yyv9VHTyNRf18WygwqMw4ObMg+S/fA1
SeqAnF9RiDvbnoxkTdaHVMOeLl0Bav7pgVRBagMVrCPX+N5BOLGNz5J9caARVYUb
gdG+ZeMizXNujD8Rh0A/94EoGLeWI1DuXK4tWxF61HMZWhBFj4hw3UvbiWvmEt/N
ItiDCC9kyXwpPID6ATERaJhypXIREAaZXzHY2fht5H4hWR+rQ+QlD/2kxbcramkK
Oy3OFJifOh+RLZSPcS3D79kGd50YUuPweW9srmSm3l0UvKjvSELMwwNZ3DNg9rqe
RDXBv6qad/d/u/fEkRVgojjLuzrEMwkyIRaWzTODyKM5l36o6KuDvYeugrcePmed
NaeSSuhFUx5vR83xcyglmlMMm1VTRILiPisOqQeqnUo4w3r5CruI/otRaIkTBi0n
O0aygLMhemtKsccODzshIBWlVFUWLmZJAEapP7tYEnnS0UcasqVWWA4bgCV0mJIr
pv2IlaqKyOqydW/y8dZrzoUjvAIISvFkDVadhniN0ikyJnmhY/OVBTimZaeVgbqx
3BDcRslIicliQTvqKTDPa0xTAOKq0E/XxWdVXAc13TFPh0+4/kHUYfNs6PYkhrqz
WUpoiT6QlXoXxjW7T+btyDsHQoWTvL6jUIJu43g/oo4StIVeoNxtAA1/B/cj96v1
QiKYbla7pw8AE6c8KaBkfe0YkyZje9XKM8T3VpIc32W+Vvflv4ZjreFW+CBMd6U6
r4jtWtz+A7jnRWaBEuV90p66liAG/QXgyZ3p8LIgm0z5YXH0HkPraMTzR22G+C8L
IhLLia6KoxmwxKGSSSQevQwr8lXQBaeA8CR11AeJdb4eCcZLQnGvkn0Fsbj6R9y7
RveY45djSoktO3qoaBmfbeXyxBMkDnHk0ymRFeK1ylWm9CJzMi8A7GrN4IsHxgx9
3XKHomJilPffia9XqOVLBHVjCpoEQWFjE4Ze0MJXxPxFIknerORK2hAc30stLmLH
pCd+Yefi0p/6HIsRnFOlJHZVvNZC8Q+7SYaDw7ixLeUXOxB/SAJiUPw3aGvZNWvI
eUy1XudrF4Yky6zc/4FgHt5YYB90Ts6aVr2vq/29gF5xeumHQLBo5hZe5/C4/39O
M7dV6KEopJwDlZSo0iWhkusJr+sEzzmR6j9Hcc4H0YvjoffWyurncHmk364vlQjI
Bfo4JRv32E81IeKmIdO9c76giDa3fABqIWx5bQVL6TEi1e6Wk0iNvgO8Xv5xaEYC
7Y65/JrfenpwLsKj8ILtas/+wXW4SCPrg62r2+3PWWGZYBJHIWVU0iSg1v5Ij8JJ
xGRHPr4cHAil+xG3ufFfpEpl2IfWh46rOTpUAkJz26ic7gJSMt+0IqnT3+oGWNkh
g0VC3m8TGgcLaPNFB+a54Tyn4aa5s+2sv83e+PtoZibYRnrxK1pjtpUCfhBOAvY9
T9mT6+/lQwopyiXcNn6qygJwux3YRjm8oZfu3u7CoocW6AWIi2/EOV9oZN3cZtNB
oPT+dmcVZsyTAPXG3En+jp7BjPuPrcOHQa+3lChzxKjAdXU4XVhhWlWMt4//0mpA
JzxJ3+L3f7LL6aeZz5RN7uoJsvbVlxU0mstGoJgvqduX2CoyjmuWOvA+XmzzAt4H
OZwp+kZmj024Z3UZQV2H7UgSZ7296KBAYK+nCyusPtj60dQJafEgR7mH9v7Mz31r
91WpiRrvT1s0iGSJ8HjqJTYI1YYDij7VSetfi8Kpq0UBi3qCpevIH5kSWLONy0Ku
T3sTOUBGber/5dhBm67AX8mBuSzSW7g/owblPX8Mjk5EGNIkFKqZRutMHWdV1rli
KHwdnQXr+VHDd2RVuymwURC5YTGyWmcVNPdczlnPlarZIQwXtkqsUHlw1vfeIlLm
61SgBPAXAHFmElLEJ/UA5g8YylR8TF2zN2D+MuC6Bla799mUTHN6ixbeZkpXdcgo
A+v/AQcSvFaOxGMe2DOHQZqgJB0NCioBREDPj72BhBCD9nS5AkYMF92AYBIsOZaE
H0MGr3OUooUzKsPZfu/7Bca+QOV57MbpFXqizJ26lkaqljj1GlZ3RzS5msaAA3zs
lIejilA+iaHp7yObHOf2mTIpqyffT1HJ3otXoxoKQsIJWhVuXCenizmnmpEHc1pT
SihiROiGDEsJMi3qSRFKKt5GUEkXO042BtYslAuQpc0XjPK2JasWlxREJ6AJ36SE
F74zhidUPuSujn6KWwwEB0ylJ3x0a/F+fim3t2cNc8yQcMSdJyUig2lemOia0Awd
SiaRTxMix5i4LXbDB0l1BKIPAckmwM3sDX9asRxYHSscLARRH1UGYd5xoOt+HFos
0CDveftyE7Oezffuarrt22qhTo2XcRib97JMt6UoJvaR6ShrOsIJOixXGFyC/NEV
Li6ukY/RZjNNCH9eciTGes3YNdgju5LmgCdg89Tfr1aok/yNPj8jgw7Y1xwCnjLm
ln5kOjuAF+sFD79ZFYm9JLweEK+suiLlOQvCx/NBCrNCzIQKPyy+ooIwaXtrF+Mw
ZtDU5cUIixnLd+nqw9Ym16bA3QaMsjAnshZ0/mmumip98nnNC2i86Z5JCzQX4YVc
sphV5uRY9WrSXVfgVjtUl/I2ZOoFM8Z1soNuB0g8T2wDAc9zoDxTEgmEfqmVC8Vt
ySjczcp/xB9IIq2EzlAoQYQB1Ic7Twv4yFTZcv5PZ5bCOOkPecwwwfXnSJDtiFZT
XgkKQuEDn36E7QaNCs9OVbJ1cuHSs788NGg5mnpyBNzlklXlMNCtlP/jJOENoTZ2
W/tPFLogyrViyXLHGFAFCyDBg7Y/5lhApkbcBdkEpZtvxUESY+jkMEdFFMfXFdfN
2IV7olu8fX30Tm/HK/mvoV+WxPzI/UnEATg31JNtKvaMe9Wfnnk/s1Vo7vMXuYmR
0EJXsxM8EJb1Itp1DtDK9ax2ftvvAaEO6GhaUBisSIdf7ninUGk1AEGzS1Ji/MJ5
5ZeOahekYx1HgZM00aeazUZ0Bh0PIwwwiSbXMu4v8opqhQdYV66aFWZtBU377yTe
PaAvQLD79bMQM4jaIOk+gled3moxXUkiEtCsfi9jdZMjPNNQwmFAkjU4v6do8xAg
XDQb5JjChYI6SpcWVpx1h+oTqp0CgyD9pouu2ena8eF2BLZHNFLf6pFQBAZmJuBo
Fw8F8aVwfNro1+i5AiqW+BUkdMCQR0m404DY8lC5DQdkIxuBm36YajdAHaqhi+Gi
/FJpxB4GixoL3Y/u16/1yGe6TMHSfAczMJrFSFzpOAe8ml+ridCo1gdGTcrk3brG
A869KWBP3r4aM0pidE9XzcEoWxYwQWcQDcQTWykPMZWgBPhFtSU+q7hfVCnbWMy4
CxZHO7P+qRylluLsyB1809ievmtf4vJffepLYYki5aEWAh9iAMmc9ORS+AfAcF6e
LxAXzBmQLz/fsAMVkjaBiNy0mSzaGPLjuVSSyZJNPZ6/fiBrHVvu0hAZuxcJ+y2Z
X/2dOU1F90jVPyXx3SdYemvtQdb9o8241j8rzGMajFPLKHfi7EB+kzlX0zigyDoP
uSVXwlj1Wjlxg2OXns5fEv/gKQQnlTHrNoqK0QcmD4aEuEI4qXCnKn1HHHOB5Yc5
iLDaHfYawN1x8/Rtby04sEWC+qW8oTIUkSpDzLn+tmteCT2EMDOkcj9vaaeRTuih
Ci3utWlMzpXrXba8JNWhv2LP4+ORuQBrQdW8d0deLjbncMEeEQNSWQbJ7kncUTM5
Sym6ZuwYenUfE/UnMu7RyCEkqh37ymHXCjzUfj7XofAdF3fAyY8qu/clCIHR8jU2
NA5GrDK1/e6VYyrwq/izdNRvmQR9eCl9ETha6DJsBHs0EBllNSyXdeI6RCxxUh07
e+Uz2SorCrPnFNPrLdouyL8XrSwyWILMqj7lRAJTeuzbVxaaEkQ89MLGdir65bV4
jUBW6Ql0HYVMWZVuwLZ8/4boqY2pNrOZq8kjNUF5m6m6qh8wqCldEeIza2IOibng
ebePFGINVi6PcQyWoHNmY3XhlqUsHkFO3OGVqySarCHR2QEJGfDB3109tg5XJTZY
JHRJ0a+SSIv5zF4OFcvCkKeg+q9gW3FByx8+Kuynyc/ad7lR60uVdnaZVCTuKZ55
CMX2QrOefVqqt/r0OmOKrpXcmSgQ3gET3hXKl/0PuSG7h9bDg9z0koaU2msWKjcW
VV75e7GZfv2mp//65udD6B5ub58edTLIAOMQUW4MTb3DXRdZ/dQIhOE2f8w51ceA
tjQfNeO233QOOIu2fJzLqkLroJ3SE6o4euR8UpCUUGMdPUxZfrJCdlHqoSbWNxt9
faqIoH/6EJNGPkxtF6l+fMllOv7IqhMypd/t2zt16DQeq8KzCKGqr/4g3JXUhZOG
DFj507nVo7iaF0WPgTrNlVKxVaDdD5nmyfnF0x4dGnAX6HOCiSEPt9Dc4IhTTRB9
tgRt59Vu7v96D+XQUxxj109TC+kWOdQwM6LdfBn0IzXqerR7a3HDyUuZJqN2ungp
ZARxORtkilQ+71PMeSXR4aNMudW6WWL3f+bGqEyoUG40ldO+iS4TZGuvAUme5lA7
NahE4x+nZ2SaYLVKkNRTLw9CLIudYHmbub1ZBnBKafrmqIeRz5vtKT3aTP+geUw4
SeGvTCN8nAhrvJj1GL2KqIyMLj+LcgTcsLNl5+o0shwQv67ErfMUzOOWsMGbvEXL
u+fnOhhuJPo8zLeWi4Urp4pfAqD5mPLs9m9imrDYT9FIXUGWg0UAg5TjQhayw4BJ
d0aYE0zHY7/l2Vg6XUl4Ma4ZQ5ObbJGWMYmmSi1uQ7JSAo8helH+HI6/SRZDq/MT
7svJEpmL45Gl10DqCyORjvSnGFTXAArTzb476isrhuRT4MFX9D7SCe0YruF6HGzs
Hdj3XUXfmIwV64aDVtHQ8S9XBz20Gw/ir58uCrKKzZAbRxvJZbSsZx6WbuR4952V
bXTqAYlH6ew/nsWec7ilhstQP6Vl+bOEMu7ZcjFaTfDReaoutA1+qk49uWVB9c2u
eNNEaJqp/CryNMhknaANkh3mvUTylY3nXL5vRNXzXQSecD6N02dhcFWLIeNnYS8I
DRCDXTl0Y5mCyAWAgC+6m/tANfcpMxY+JTvMSrs88OpTcsIUPxqKLIKFb3RSe/k+
MCoHvkVXYt3wTOcvSJjsD4+Cmu820ysRrbJUd1TffiGKGyEhjiwKNpKzJ4ZkqEXR
NILdRI2hZoL1xLQkwR6DB61bpkAFHMc0ymC+1sMPHgCclP1gF2P3Olvpj0DBNvI7
wbgf5eP4trJwuo+vSz+pC3N3l1LPuD9F73ZNw8BXumKQBWsO8/02xkTLFXVZMskK
zygqswjuri+1dn8Tvplx0bJaJ6LUEZnOtTxShptq2/optW5XgKj7co1olMmhBNcm
RKZ89ZMPwHpxB78mgPQayWmMnZAaQyQ+O0g0aK/x2HKPa1ZN+SObYCk9YzGkb8Pu
uSKvwymvoCizeZDdpvV58wuc+1bL3ssHr6Un92yj0RFIN1jg9m0ZcYDUYnHmHhOW
cvwT8IfpfE2pFKt4gX/ns+OCflsm8CBNCcrM6eSv/WDcREJkLItbIdqlxgnK2yqw
Z0lLlzFosUJk+knyOA4mTTr6nXNHS5ALBMKdRPNLqqPwVwjlEdQuxkxCOlX6yfVh
uYa5Trho9o/hiMRpCgKkrvyIR65dwJyfybDvS8Rn9JWpOD6pVpbsujjPwisZNJgA
TilrW77vCvhzv1/9aunBHkmTPot3w0Gz3h9KyfASpCGiqxmTt7/zvF0uoyjMGRrf
mXYGnUNiTeUx756AQKbkK1VD+nKxYjri9B28+WIx5imUwmchBaMs/24Wx69b3S4n
YhEesCky7oIP4bsYUomRW63azUVk0zE9XuWiabB7NM1ZuDcEluWloonWc0Vmh4Ei
iGKwgxnXS7Yu3PYeit59kunwSFDAg0BlCb21ub6vir0o7htDAlBAof/Sg2V6gCIV
7v5qUg+U0T/9jTDuSLqB1pqNQnQk48gU/JB0rD4Fy09vzGdRlSzGiYg+2Yaro9k3
1mh7vTpdT1TTuNJFr9ylMKl7YeQsnOhQsQGBuBQhXdzfMEKw+Wwr4VjeSt95WT1X
nHpVjXHaQmw4MNkqFxxMh1IehaIPU7u5ZaTazBRRAaZ/wckazUen0zVLfRhz0LKa
r+NOYEb+DVIUfIoLKoPPpfg2IWS2IgXqIgKitP8Jy+3ASRHuWHZitmZA73K9bE90
CgyDX2wQEItWD5aN+AVv3SaChOAWAHnCp0/7SzUZQZPqsi5UN2NhX03d9wc07WSz
e6WfKH8jBp32WLB8JO0bDbVQRIVwS0/AdzAAJllJGuopqoTCjb+8O7WjcuPWFQfw
l//y1DS8NdjkxzAK6GY3t7VQ37sqDAqjlVEh1tVx/b6nR/6OdmfLcQCQN+qs3U5m
YEkefDz+RZhZvj5QpPnmT6Vm0et0t93A9COPDwF/EgIciBncApj6sUbgjRaNnpuz
0fCcwFePl/C1ycPGbMkGReJuWqGZ8MUhSBSXvFMzqesHbNQpjKrTbfvA3ZqDBKJB
DAj9NyM16jq4Hp7rXMLL7qhN03s8bdUrFlMR6ClrMBUatCuifpzx90r7CbLn7ozi
BbPeAFBt3Bm/jAt5rgtVggAgkdU9TXY9BoFRCd/49vAQtDyGFKqiEG9R1CXK1YPA
AzeTy7i0nJYSMzd22+1bxcckC/4Jc7dq16KRoUVAObs9Iz+WI38fjLl04B8jc5Z6
J9FroBkD6jNElZMn3Q5PrN2kqbnRu/Klgt9lIkd5pRybi+uYJ32QVlEK3plPcoRH
RsXqueDl19sNlHIBB0wUi/W5bHmXQCuiGl5tPTYX/FifUTubMyhescZtzhKNJQ0X
/sI61MbFhxWpdI70xM7zbyagRGieZUods99x/3w0OXDoqH7RjyARQC5u1A1DmZ3A
PfZn8UsFkDaMhaqNaOAxnGd+NTsN3iveI57ROVI4b/8rlQD8soQh6B6BhKnpC7JD
4JIUZ380ID3afTxZJRRMNTMpkZq+qIr+uK3h8XTKWtCArTGBhzpGsL9FafhxMWx6
t4zScxbwNzbPStIZlQAsT0NWiN22xpQ6TMSoaztpbcuec5cXMiPAABq/oCquGY9N
bozm5C9EJHULOOIrxecMYNGPYK0A8ZNKZHN0iFzAGwMtnIqwtkbwaXw+ppJqDWtg
FRFLPX3+l1mSQbWshamX+2paIwouAuXUByh8fRHoVrRswxZQL5QMpVndNDLoA1Vj
d+BHrQAmUQkwlOSDxP61qlrUQJttEEFMD0xBpZD+SJGixaO0/1HLqPINTSM/zh8l
Hoh9ZINF0mKo9+tnlDsHLmPw3ou5f5cy+/UGV94w//kTNa2ubcWmUEQyddyz0baR
ihVAXiFthxDz0Z6uEb7FTvPs4oxpQ3FueW0iWknp05Ob1GwA+O5WPGHx2qbzvoZ5
CbP8722vzRbIIDp2An15KEqQ6gVJ/bde/VZ5gGmc0+wF43JrC5fSrqEwWBfYPiX+
cG9sl26aREq8ePUVIb4AbQAUFa7QGioCT9GPDFgx+ercMMTIdayfn1xMMCVuz7jV
goL37VCRGNpDhYMYO80zMDs8IkXYScUVHxg4uXTTZYDGofsCNrcy4g2ya1kQMIwY
MDqAitDkAOP5hNmVFCuKvdIEkRbgOVhyzk+mkmrWqKjndNuR31vBTKROe8liPvdX
oQePy62MUA0fjt5YarIA3I7HZodHlUbIKTvIMF6RTJRqtgyHx9o/YxCq8FUb3JTf
2odcTgXD0h6LbXlvQmA54D1eOeu69ieY4+bhpByqg4E1DAGPsdI8KY79OAms2wmq
uEt0R1/Vs3fVd2XUVRL9ldxupzVGI2f8uzf1i4v0nt5bhVd7eci8k+bsxYnbbmxo
1svMXl3lcY1Uj7LSW8sjXBiZy3n+i8naMm6ahX4ca1H0yNfVTb2y79HyMEoriWGR
nTs9ADfZWe7DHXdY80gCQrNiwu+cWSLnZ5HbecLJ09mmdJTyrQYVrdPQKEgAsHDw
QNKl68sZhOzaBQkgLE23bbQGZIRoY2E/IdRG9e/ZvhcWzmPyNVtOvxJ7//GK2itJ
jLYzqAzAVjijqOTENQsNwj+9UtmftSFuqz4GvGaJQ1Uo0Hb9JUAPcVWgVcRi+HeG
SwouLGZN3grVFDCzzM8vWJrhTq2pJuIwGOms8peuPLlYmqvYc5iCUYd9HL3sdIXI
hOM/G1ACdx5IDYoySfmsF3a+JPBvVwfL/4bvb/oR/RTPn/gSy+NG8CwBkRwz1PkA
Nmhdxbd2hM0vWpDMwLSt9DkinEtoD0GQzEpEvGnhZiuFqppKMDs/XrA9HsalfKY/
5Od4AnB09Tr8Uxne8mmR0gSVFRBVHtec9O1sh1pfw0LkQhfEa+n7B3atnZ832e4V
4f6QkRbImGR8439bq8z54cmQ1+4zKZpTizhQKXZLViQt6aJpwBPqUu9m2EweU/ze
1Sx4HSz1p6uVpnU9IrnQtQPpX3VBzFYQToBwSVkx/E+al59BXTxglvyS3k2FQU3m
HHjC3Btlv8YU7uSppzWhtkpKGpT6UHxYSS4o+JC0FAR+dhj8glXpWUUdOhVB9LWZ
DDzb4n+1MiyX3Am0NaGDOKI28LpbgSwcVRH7HDIYbaLmidHE2gnwFPKpaDVQbEWq
YF+UULjliTJl+/YupBxUSLJUYELduX+E3W+0c0QN6+wKx9YODNOKtJwRtQyC9SvF
JszLelehiFpNk0NfP6q9ANOz8oPUkFo5iJX68N0Dw5DmDgp/mK6DmSZ8Zx/lAclJ
u/Li2mKCXwz4gWKFdxk+wFlBbBBUgMlK8EG8NP4t+io103tzuRmhBdhPMVvr/ppM
ID1qDhrmDvuKpYnp8edpSjrv435KXiiE2zH+5eys3ZEJ2cnrqKCoXTEhDhwts7dN
omPAspOYiTLCe+jhwpavCSYSM3NxMtHILCuR1GnBzZM4Yh+6nGXKHTVKSL+Cj1Fp
BFFiq2gN/jcZJmJHET/+jMNvj76nvASyeLZRO/1M/7WzoI+iO8jIVesgCjoUyLxj
0jPym2c4jknlHwV7pj6+7jPmFIMT/q6i38zlWoHCm4A2ryQRtiS3PlGeRed+WSht
i+x96JS5TaqM24+XsO68dQub++wkxx+qPAM70wbUQcl+uoGCs25AJQ0cB7upZvIL
vGnmfsbF9yCsT6i7hTzk+Vgeb1UV5nHPYGHHoLS6EQcIdj8mEHZ74JKwNkPEdJth
WQCIaVGyqHm20xKeIoHOAZgb3RXOQR7y3273Ga56NIZ+vNEeUzJbWh5K1bP2IuRT
UpZkNhuXZgGMqxZulLRcAFbgURbQEOIql23+nAk+9sF7vtT+kYNpa+Iq12lEErxt
3D97gCYYyEHeR6/3cOqywc83wOpzUuadZCY5ioQghn/jEO1dL3F1laz1V+Yd3aaw
Pu5orkRx95Bx7sZVmOMYX2BNiM2j2cRZjvcEThIaEEpoaF1Tq5wubgaL3k/kGpvd
tGNIRClyV5kOeo6M3EiIoGvbP0V56qlqHu4vHdnti0tTeQMFV3wJ6XxE/M+KM+HB
XKv57wNSVrMuLmIkfCWa5el+BdIBrz3nvQ3R78gxPwZNhDaA0f+jENosYC8+JP5v
cQ1jVac+LtXwe3hBUvblplBirpaW5j5e/2fQYDESdLFsda29zoBmZoXrVgNRtOjM
pkzYNY1oT8YvqK6Sl3TjyLu9LcZpoKXmThWjNgKOo9LOUtHp1ZbeUui4n/v5/bHR
8gizxqYwuL6JhBFzzuhs0NE49aNl6o0+DOBqA28NlA3hcjgAma/Ik/+fvevvsMl/
B6aGjEt+Hqw5WZWPgXImx/Le8lcgmaOn9Fdu4s+qMP6UrDOrxSLzpOfFoxdddidX
4afnGSiBUcZTWY+X0ap5zRXA8w+Q/df8x58vCO+b8gOnHASyt3VDpoBLQdueNDZ4
1J3d7j5INc478pHZUZ1ep+Xunu6Jh7qVuIHaG/7LVw2P2ie2Dcu1pqgjp3AjIVad
w2Uy4avHvz/Wo5BuWRZuWnKXQbJ6V/ipJ69mWnfi+iv0HLnw26Q0bB9RmqdQz+xk
gEWJPW4HtBNb7hUpFlTsGkmTKWaW4sEnAw4MPb4WEWjqFrZC6AQJktLVv8qHX23Q
ZkEHcMD4TfbqwARwxYRhfpWLOliXWjbnZKq2sSxpwNhJpQm16RhRjZ5OSrG45EzW
SqaWLWN1oWfPDXbNVSAexNMVrLJb9VJJ5/GhRczN6ldPTD3FUyQHb93Zml1k6yZ9
gl8SsVJy+X6VA+VArpltFw6LcHixx5DCEITmTxl3VnLdykW7CE/y7hUi7kkoGn05
oU67tIPKYF4LbWgAkGIqdqjmai8K7Nd9Zak/tBQK8il6SjiPkzLkEneX4SmWjYP7
h5sdlalufp6ZU2FeV/hSqmMFeiAncqHRzbaX3gABiwb87/dWk4u0aSJcq0rtV4Mr
p/+72s/52jtzyytcCEZmiJ77AikjWaXp8SqFAiGmYvjfSIECpz2Zwbo5ffeHPdd3
nXYqmFjtpUfzU/qjO8UXu+PMEIdojifzl5Y5FSt+2qiuAtLqIQpUGqhI0gKwSTQv
oW6z/PiiTA6bJAs1vrud2kw4vvDgPPsq9ilpAnLRmio/jqQWawwSH0THk5YAll7+
EjjPkc8orrCTXsxoFj3l1KpID5yU3LTnU1r5uJ4O04mCHChwe7kzQbz4HEFldrOC
M552LyRA0l8Sk+N6ed4UcYqCSwiKULgGRw7b8/dK4gydn3YOq5K88qatWmQwVs15
AT8smiZqhQ4epjVlLO2ZFuuKBUiCL3dzON+KqExGTFK2DIWZhCO3Y0j+dOnpnjf2
xXCMMmrlN1kp6EnXvNipbCZBkQITohoBkQEVPDCr8ZKCc3Ki3BkyWc0L3f9tx8sH
pmO0q1BPgYPzd4R+A5H7SBKA6XFgSxCrayxXt7gYpFkrnUuWaSElBZJb2eJKHg4c
QOz65jayVX4AxkSDgoe9gK7YdX7E0M66yWliIlgbNUFFPsVYw6aanueeD4Xyh8EJ
eoGgtOt60aPKTm6Efjjj4o+JV5Ber+uOJPFFB8b3ca4aBUcBtiG8GVgKe6ld6dhP
GeFCFZv+bMrZGDGNj0WV7x6a7FK2t/iLKuOb1vnkqmZgOihLpPPzR/2zaTZt2H7O
pDo+j3tdcUAPLg94iMFb9wMzc0V6CtzfJ8+B0JJO2p5I2uD6nAPXpyBn8QZEdBxB
YMhtAQq5wFpbLHBfKdzfHKRRRiuKNAiGGjAU1qvKEYAgCeY9rx2htiHnNyzJmBYu
4YPAalV27H12OHL8y5o33D21CjsqLeoEG4dybBShXQI3FaSRxvpz1Uu3PACz17qp
pmgQQ+u3tZxilMbPe7c68fVZ54tSfszL7NB3U2WPmZn/60arB28f00bEdf4tSefo
Tmh6BUwEiZ/xUDCVuqQQLx6WcGAJ0kMmdkJ4q3Dtjv8ka3O6Ti2lmS4B2/BDiLE5
6HI4ZvOJwa833t9GrJnea4BrWb3DXuhrPOD1MU4hf0zG1QgLcBhtq4SZyuN0ifT4
Nj4lo4OlRAdSKs32zw78Ly+RzBF+fxAH8dTOUcpoStuJ+AMx3cU9LT2aF20tbTRI
D2no0W7rvIGFl3C7HVy7Wp9xT19KF4Y3vDoAkOELZJOuen1PiY/+beUMoReGggpN
4R2VvYJmg75t/kKw63VeOEgqK+vnyIEDAlJu0FKrq4ZLAMFlJKRIjxAghIVL4xuG
+24h5NQhSdwC2jyONjFfmd7kyKt5xNzpa2kJbICMDKs06L41GLqcF8yIcoxByXV8
GJDjVsvBp8RQSjNV1zNrPnWCvifh2YkQGng5DQPYFHA0LKedG5yTyo7xmUKxpNUs
skOnPS4DVD0lyGdTWMBudX+qkwXeO8rs4sbrk8Y3dgBxp1jYp0y8cAJ7FmCbxojg
O7fCzby3bJZd2DUQOykhBxRcXiwe1mzbhN6LOm8DYlFZAJKfo3Q583WsA3CaJve4
lCFEyYYGz7m9aZkbPwC8O6sa1z4iThFuwlsL5AMKsmj5BAhI2HlbeuHKK86IRmrL
fuUS1imQunvKKYeZL8Y0HzZLo4xLvXTScIYPbcX+sr1y/JKHg1ZQ+jd7wHnjal8Z
a4BlEFcZDeiB3s5vLhwxdpTXuiPHZWqEvFcJUxgcMHCedshvGgoyLq5+7CsUSn0S
TlBpbwoJRnx26ZEt9FWTcrpJqbXp7dTDZMzpSknw5XC25SLqYfZdwvAWfYw8izk+
CCGLqni1c4n0YPdqeK/Ue3oWNmQkGOLiOur3MZl+pJ/3zeR8o36kv9jvIoDkVOB+
0OSygojYggJJ9xjZjUbd3LhFi/uDNtlv4/cZpdKkztqpW5FxJ9HqNd7262pXj91O
/Adl3y1X1mMEyjfDS7YoTAXiyfEnGGzNS9ZW9dMUbznxRgwhZHAFqg07LoHlI7Ub
jT9kGoVnYs3SlKU8aHDUzJqgyHVvB77l3rhT344QPVx+HqNFQpVrAZM43ZYKqJSV
AfrfFAhLCsa/cFXLxDjQfATUhPCFvteK2HB72qGLkgV25qgP/S6V4/VdlDbdb2s2
lfq4ZOXnSf7X3bOxtk+VL7ehcuZZVe29hhsRgD6XA7M/BuVGpInn9dx3CV3UXH/J
rA0RaqbPKC78sJJXYxqzqpRvuXEFrGDTWDNVPj8u1WNjBigs5UO8zU72noa/1IKU
vZrv7N659YxuZRUWzWrYl8GViLc6HDEKEq4TXw/+OGahl+MH/kQVWC5Y6RfJeIon
SWSL8JwJLMH4quODbz3UfkW+LS49rMBNhCBP4w8deIic8pEqz6zRAfqIb+J3xeIn
MQEdnSgz3d+XrfGXsjwlsy6v1SQfVf/0ASrPZBQiScr/Rbvguo5L7IyDLl7U1Mil
OhwbWKULN304dey18OuKNpLnpwtw0GfRA1qYdLZDAs+rbBcFEQ6a2ALLJ4sJ1Mn/
KlEE23EIqJDs0t7rTphMXfEkrCajx6xP1jwgr7CCWGBx5Ox4t/nTlDpQoBK0rtDQ
YLL9z8g9DdRZJcdib0B24O82e0UfauMwpIwU4oZ26V2qA+HP0JPP+LUmBfrC7DTa
jO/mZxdpYQdWwiw4CXw2xe4vhceDiAqAN/EuE5zXfcTuoDiSWct2sPUl051pWqm0
TR0yNoIFg1PwEVBDDxHGSsLnRqPlhHjQ7HbYXzqqEBq7avvIWjp3xK2qMmk6dhCE
bITlt5FTikgtHmoYsYfYec3UbQqgjGhO0sirMWC1mVSjHtljBLVeFpZozl2InMf+
fJDhO/GxGihD16OsVI51ZqHKFsJk4Kvpi64TqC8CAZyNotUiWt1TcnHP+Cynzmc4
qvQa6LC10g0mDu/iae9FbrmWI3RBM6IUnmH0FMMxtJ6BYWZSZ8C7NqPGrJhZVXBX
O79Gple/oxdGpHhGM5nYaloooloaNAauk/5vX57G9XZuaYWvoi+O8UZesXl+YwRO
ySV0190CC4ciWMx544qa+6ZigSb9U7k4+jeeDfJFzpSbfwQH9TAtWBt7TAJG1abe
/4LM5o/GGOg3KMYPXmf+/WPITr29gnxv6CLo8AVam4FyylIKTrN7G2Ev422wUxmr
pwvdJhoPBrfy81V3h/GSnvLndfiNZ3wbrl0URQrCYFA9NTmtrndAkq9bLgO1+cld
ucFvlRCA1DROFoOson6R74wv96NoK/DSnBzw7e8DzWDy99fcgAzCzBPWfkpjwn0D
gT9nSI8NuhCxHQk1GPsr+LLPl+nn1hLomNZTYBHRgXKsuL10kzWWH+P1HHXKg/OA
djX2Wy+g6G4SvX0Sndpe9KzS9cLGjJ5Xdjht4v2NP1GO5ExOwzRAmnzkLOsS0qQQ
W4d0GoisxNe/btyC39lPmTKhVfWaMn54kXT61zI4jUjKcAHS//5hEIW3HJE11pYB
jwpa7GOcW6GFKgtrHtaHuZAaZnWV5LhrnJMuDLV5HzCQIMKBexD1jOKu0ThjqL3f
JvsSTOPYflpBSKKTk1/dQ/1JnpZC4c6tGDI3WsPs4v9V1AZjb6UBBkeM3vcJcHoe
qJsQCWdP3KZFV2rkkchxFFPTugIZ1zKKCYoARx83Buk+wtfYuKjEqvfTYkHFk7hz
VCWNv7Yngeyfhxm54BuL/eRQS6H3NYipVctolpMo3ZWaNQTQ5Po2kx/KA/UkDYZY
sFkpXhbxRiGKVtbQ5BNGjVPItwVpCnUfuSM1GXByt1IdMG+zLAbXo4pG3rmq+X+F
sEle++aNgtzwvBn7Ls7ppfZak5+vipSCdERiOtArCTkDXbZhCOksfjPOmmS1grMY
d+CjakIS7wak5qf2bXVTNOwdK5WSoJbr6DEhnrELcp+++iPum7D2vlR6jHgssAIB
4rx8dpz01kapZCy+CjgJaoLNVIl/JmGfIVfVGW1XUSjQLA57a1tCBRf1RrPK0Y6v
G2MBz/rwr0xtG5kvger8s7OuHz0XRK122AQG7zWSiJIynPIGQuYoutXc8mZsP5uM
DKscayXqNXfkuizvN1HiFsyBm52puT2XQqpeYkrr20CQShLfQbLpv1rnNAU8FUga
xhicNLE4lZfjFgenRhR1RLpmegVgJq2SH7Qf0u1MbqhF/PxDbp8O7xVhQMjSxbix
7y1GyU1InX6QhjvxHmtPxHzjfaTkskPaV6daMkC4j0bosPpWyeGsESIgApHMsHTP
HrGluCWNgeopJn+xaxwSUExxYQlqF6DSeWEGCqaBcjKvxoGqQ9ebjj75lQ/O8CBL
EqGoKoHJR8q+6lSFQe9wO7qB4XC4pIIqwo7ebf1uhEK5owEG+QHpt0X0pDpg2aI3
rmDZeLz613a+mkb1TDQmKbEdfWY2lL0uqK3DGcCaSb6doiFWwLVoRmJCL/naTacn
FGuPEDxqGTrrQqlSDPFSl9vI73sLJaJF/sNnZxb9ecG5em1hglraWRkD3l4MVTyV
6IXpnD20zlKQn5kx35hLt+VcVMYpLQCxt/kMPTmQbD6vaSHt0Vd5QJ4K2ybQkYl2
Xu3XO5l+8s1elNIqFilUynQ6D+CixVBmz2YD9Jd8/cKLyG1sAH6Aa8hX+D0E2m9N
XMsxwlHszu9/VBAz6S5wAyMb0nWSP6bS58mcDHLt0QMrLe3Q9TxDtDGaQtX831X+
7kKkacH95Xf8PDXgAoJZomDAwM+QUYDuv/AATLuRqHAe4r1/FqPlmPbhOG6Xlb1k
BLC8ImODCV3PahO2xLSBINwYVE8YOxUfdqo/bOql5qIVI8Tj0T9hG++yHbRmjh73
YRrQQAEn49LLjlcimI1j0ryxiYWy8Tm3nyiJUrLDFYbvmlv34pz3eJwkH+98yi+x
+SaSsRUbsD350ExnUJfLTalOCXXarQYFZFf8Wp7/oMQsW5oMmblOhq1nNLrBEx8N
AqaOn87euDy9C6ReBp8WQ4wAma4Dzb/zdWtmAjZPVC00yKfeNCse+bTACV6PMacX
gqJAanQvANlydPBWTdskDuL6XLacdZyWArokVcrk+U1g2x4FsUstUyxFEmzAVUkM
mVqoV5bCSfTUNraC8/OAUOUGFkNBUaxWFc7n7Ua1kMWjBkMQGu2Yn5XG6eT6gDYq
dD8tePyfuZlRjVIYrxM02VYoF4zcfmiyREkuZYqdoTMK/OwZ3YKeHm1D7qBAzoND
2o2i7OecHWFTaknAS6e7CmJtNnJq6bcbAbz7ds3wIB0BInysJuQ73u8Z20COrf0E
43z2cz8wtCe1wOytagUG0bGHeBh0PAvn318FG0VQTA9asIm+ZC3u8MWn2QuNf7jR
4t8x36epL9md9VqSz7DDUX6W3oOK9aIJzUAe3rO66PsZuSazgJyOCbivuJ/P+cc3
Pd9OQQM5hQEuhVAQXlLIgLspJYpKLXGLd/CBQD0cCzhY5x9iqZbyMrpQ3W3beLAx
0o7wumX1RmiRCqYzrhzd1vKAs4BsPCpZqj8A34O3HcNpnQact6oMPEbzPbddCW3W
F8WqYlmTDMm7/GM5ZUevyPNE0AVkmrtNP5/dG+7QO4uZbtEV5f1BNs4K4P3XV1X+
qQKzvEhAhN5ZNqWY/2hdzff/wVKXgmneoQmD/eTgMMtxrz6f2KIRx0fCCMpN7Nnx
2LusIl9l1aTMc8c7xgbLxJMnhDcLWweTNrTKjiAMs+XRo4CgtR26CLuqV+TWSbIh
7QC2pb6mTXBdS4T12y7hP1mxUnh16SofBa/eWjj+R3KOQCq2j2Oh7f+Lpd7e50JH
roQVh92MUBvIX34VTmRQTwpqTs6BVJIpoNfg5q7mfSeLjQYyvr5fj+xDU1H395Zb
Ql1ub50FfS1DQL+u+PgacfSqQamjRd8cnj1IeZ5i5ec98eY8AyJuq29key4AWvxn
w32guYWGT1C44zQ4V6G+HsCxA1a+YhAqkoGj6FqVsSqH4Wzr7Iz2aNNNjzq8vFNx
7HceUgqszHUA6z6epkoeb7wlv/wqBJk+DWggKBHLAt/nOpYEp8FXpyDzbmvGDsOF
PnwIyyt6Fm6mzd9nPUtmKr2KgHvzl4bQH8itYxNpOTWRWPDP+IJEYcEeLb5CwJbZ
5U759RGIFIZDdRNCkGMMZpf4zpNbOVovgzF+3rWOvpZwXVReW6Yghz8BSE96j/Y8
pMuCxUlYeUJKtUjA7/fq47HdJ2vQi8fodh1ppArLoWQgDFlE7WMruAYqGH/4Ewcj
PDJp+pi/6fnh7xABOipHdjE2zrT8WLH4gipRE/fUVUhmsDR3ZduTcIB7vDd6043g
OCqiizC20UzGAKdyGlrtED0oOoU84zfsPk/YeTotBeec99GZia7/6Qi0N3S19Fi9
y7s4Zywm+Z5hu7jOEglFzqmzmmJmf6lez6FnYGhEx1ztFx2S8VapYtvDAVAy3rsh
PXYnU2GDkCzd7SpJx6Ay7WTiuxQjxQYkoY6O2K6rVBx+ZFbEETng1V9RuXFp+z+7
FiZWQEzdfL87cpCCYlrFC9YSscCCAFrylp3e+sos/JSdBt6IsbzBASKfIQ32yfsJ
6il+eOrGGuoMmX/arjrImlBC+oEvnmH5MIYJ+qp0Cqj5FCK3dx/+oMUIH0muViGV
U2ZhAsc6sxiolUzckep3Pjh9BCys3pIZDh1vI1TSh71xj7UZJAo8J3viBUxp0UKS
1jMsNFSXsKlzTLtw9pA/MF+a2NGl/jqcNMiF93efme72sIOaSlk+I3OBy5Avi2WB
a3m+KqVLyYBljGWo2Z8y1Rf3IDHPiYsB0h6LdeKiApUrnfWGFtxLrlZZU2j1lH/9
eVfSfvTFsrVqYWzfvsQn3yPJiMwL1bqyzgdF3F7rX8sL83hgGahpwLuPlm0LzAjH
0L23ISqfyBRamcgDvHHLO6hUQGoz6xcEXBgKUXfQtp4+KucyzS9/MPaHoswmNh+h
78ab+79oN7Czzr0A7G9CS+Fg8c064GbXWcVP2QC2VArmnO4fLbVdohhHDB0fWNZG
lTALIMpltRq51CpfsAOzxQW5yyvcg/La8JocyHEs0HdcmzAlfjTpjTo2y+UdVR6d
ZP1rrbqucmwIz3P7/nn4dOCpzLiXKOmjwkfV3dE8jPH8gCRYGIrCFFa8bPzOd60J
qlJb/1sOZQUB/yT9ltEYcaoAlFiudIuzWqVXxxN7LIqh+f4cfJutoHrwHL/iymOS
fpv2PkVOtHuUPWAFC+nf4fuh5inMuGHsjkxxnIN7W8PU18zqVZNks6OGJaLN23KY
RgDD0j2fvD6NmR4C2NIlM4LVz6W2pFkgSCzXEfBBJDoxNY02QeRwMsIZCRnaqBc0
EY+28aJiKe87eq4jXGKeyPA8DNXn1MSsfhLZzLKTVIKDyAfd38wiITIY6BF5qQS/
6ITYXhLEGnXPs8feIeYg3TvU0SmwkhHkHB+IkvKtv5fCPLjQ+wwdKkPGcIu80KPm
MCbuzkNfJEE4jIFnF7zay1A79pvm/pOjEQxOAD3ibT6QLtj/Ay+VCxP/mJqxCk0N
UXhy4ssiX2cAxjyODINWPUSpyMoaft+BUTNhqDyAllh/57kMiqrv1B1p6chIFBef
flaGyBEJiLKuSdElyhTs1aKInlA8uZ+/TV8+igbmonAWsSgN9fTFzy4ZeY3LRsS+
dmLFj96L9i9h39pDIMelIuVBlLD+FKfL7IPeiWA3ZSMYDl3bJLHkd/MyByVZMbY3
QQsva7GBHWmkr/04/DcuCyON0EUjrQbadB3P8qsyS+O1jU7fmaV7Z5jyhEUXGBqF
bmlBj09U3HBwW2A13RBSOvfv87w8rFYcMgzekV2dE343iiRmHaggfwPxsXxbP2gj
PGfyiu3oCOvbfPqkUQgbsMhSkoGUDsG5Y7TTUnZo3mUntTUrzOhl0uKfwx6xUu+G
E0MkM/Tdq9ttkYojuRavSpwT7G9YbiNDC+M7BQcPZeva5d96G4G7VcMabaD4BKkA
tWkiRGMfvD8p51CGVXncInosn3J/zgl0Q4x9LiDikVPDK5/culxjBPFlEvg+DnjZ
bDY1A8bFRkEiz0vGkUQKEdaKixG3agelxq84TQ3hEpEPVTqXprLyDeHt6Y+9bJbb
Q4BaTkPOzOJ1zu3f25xFoc0rt5piCHaXgN/L8aKJZCw2xj9+AORPfsqTBKM1rSkK
epNrF/QnqxHOI5WzIgdf9sL8FTZ/uItw0nQhwm2zsvYlrR4HfP4rnGQL2tMxNBf6
HBpJb9GTZg/B2d7JDFZfdQ+wD09hsdYFNc2Fh2WW08yF+6XcAFMETQd46fQ8yLlE
Om+j8OmFXTkC5//GqGjDTZFZHUgRlGO7oCAjlXpzhaq9sIzl3B2ZM40iYioi78KV
KyLv2HwAXxX9gomJuUoHKL0q7UdNAMULjOVuTY1Q8xpbXYjK59U6KfJukGwHiARp
WEfSysJWJ5ex5ukz9Aa/r38i/XhjT2Uf4AECc5KBh/ZuJ5SW/VN4cBo3vM8vtB2M
rVAB7XklKjQXSohjkcQ3kAMs48Nb/whCQtBeKDE5b58wLvoR7M1qg20U+fNprpQk
2rtzflgQ2maRVGfoT9tHSPCSjMCqmtlDZHAq9t/aAZX8H9mz0KclW4Tz+7NhfW9D
LFPFLwa/tMYA0f5SLnt90XqFTOqThwNwWsXs2Qsx4hOP+SFQO2jwJfmoosXBFoVT
v3OZRYa/lPLima1DE96PXQw0EjzKlHsz09ftKdcVV5UQ9cqWxY7PIUbv0oWzSyKe
rYwZ57DeFx+BnSNIAsKZAeLTZCiK2h4YaQ64F7x3DztIVxT7LXseZo0ftlXGSZ9Z
K9XU22lIoKFgDuV7mW17m0ZAk6bHDJNPwoqTCE/KqgAk8czEl7CollZScOgAJSRX
iVDAmLnYFjHvUqZTrmfShBpk6FGI3+pyYowwZnju13Ws/YcH1QDlLMg1sxBchKEY
eKaLo09xEgvpe1I0psE3b4jc+ZupYbRtILGrcXayZtDyhzvr+pnuqLkWhyhYWls7
3HYC6KbabFdHsbZrouZ3OiSPhfFarRypvzwqZHLY2rgeaxNN9kZv9YUG1bwpwK8O
r5m5BKcd7A7O9YEeD/X8qBbOUWllL24b7RImbmpS1QTFW8ipEdN/GaQK/Jnuq0Oc
u3pacFfSePDtEK7zNox20k3smJpB0CbiG8xdiTn6mcLUIZXYrR/v+wwXqzFsie6S
t3MrHxp6V/oU+9rzTQY/x04/S9hQgVTupK/LZeBTsU5ZbOYYMfMcof+j7FYnyDID
TCmUmfVG2AEG6/hhPQ6i5KiJZhv3CFumuC6boogGzAh1FaHwqdZqFmM4pppK8e3M
v76VQ6uCiIqOz9C86f64T0LByBr0IOUkGWfy0fE14PrEyJKlIGJa5TLnpC71NJyI
Esb8FXDeu4ZXoeXikgi+DUdU4BjZxX/HjcoyqTgN7nxakvfc04+qbexWB38rx3f2
k7pu/ys4rVa9WLoq5/A/1e/PkgmIgwiT4BFOBcmeaftDdJ5Zwt4gu/y1kxMiLdgI
yZYVNPBhZBtL3Y9pfmS2FeT9+Hq1EkEilXf7l4BoZi5DbmszJI/uwwaQRDlEClCS
WSnKrjYPoEnqUe4JOQczaOy54rXyHQDcSbFL/YlQYFaTwDY/7/Go1M81fXeuQiRg
IJBqe+VyA8bxTNj24bYzy20tMpmYo9OO3ZQsa1f0cLVWjaGGBIaefGqvHFU+qsJT
WCzegX/hNI/pyKv/+wh4AugEWrWDbXQlzrhFIrLUIpkNjAaAzfp8v+MH5kCtb1ZR
4vhr+2YVL9w0Yyl5AVDUF/S3aGmSQISOnXj/EZGTTVZbkn+1NFAZ2vynOjAWn8yL
WIPf+j1VbYF3T7SziWVFtR8VxAuZur2KD7hw7o8KtQ3WqLRWPc921fMpn0RHvYxV
DtN3TpQS8MFziDAcnW1xrTPUOzkkK1W4WXhwvEtkexkRwRa6Csyi7WaxS+bBhv9W
lxGsbGI63qiWQ7UdXBuBPSM48zKe22lBLKCoK1xrNoIowiRozmGDCgxilyP5Ej+5
UIiWsJXwb52M5aBe+87Pt4thH4bvl6NN7tyxFoJYl1+hZ3VSQpcpDwwAJtS9Hg1p
ONx2smH+Qkh11V7dsZZdE7fu1IGOzEztC+HmOWAej29TdhrM6CTmu6GLSuw3bcCV
Vpx1mtc5/easO4CSpUFFj2n98kFrcDooWIik94AI/brtyYU6YemYpH16KpsLKejH
+i/90GD2t1L8pZZKJeIWXlUYh2dkCCy39zsU8SGZY17HmwiwGKYX12nPbQPVwZYE
Dvz6mviXvezn0PNTreviNcsCzPKgqJqYm8F7O4AMyAcIiHNguNXyYvLn6OJnZlnW
2KqtlsZ8szgCw/Exc+ms9CyB7bRjqwBrnBLTySGShZWz7p9qYGtblpiroCvmhZF4
Qej5xTHa0+Nb81aG0buWAYFeFsc0NoYvC3OdBr4Rvdc4/AS7od59v8cPf+5pwBnK
Wj8rIOhUw5rxm0oYVa6cpa1fXjFtc268WgO4GP4ZsNo60IXUXcQDRukavaRnpv2G
DS0sY9kfr2vARf+Z/7SQliHs+37gBWFWptYv6zUru8DoM+Jy6XWPL89TwAfqPG/J
92p/GMCdnBHHiGHa2CKFidTNlYgYNPAJb6zs65tVCOhiUdoK95dXuA3QDMi4KGC9
FIBGHMAufNT71XvUbS5EbFeMSUdFiGNYylPpPeCSXPlBOOwBDUMXZ4R35h8fcKU9
MYApzItHu804pTCC4gMWlkISUW5Qt24n9J5V4GoxE7SfV9LiL0LrRIYni5sys7hf
p8i9JOdlqoDh86iemk6vZ2O7fAaWcyT8bEfdERAcpw4JYupssX02GLfLyFd7Wvr1
dxkmY5IvMdhH0uWzBGvejnj5VXGwG8TVDwf7Rjpmdc/5ub6PawMBZK2quZLUQ/CA
saiMb+xdnpvnestpki1672YN+yJgmjL62ncvPAFoaRelv1qQHQqt4pB3ugDrDuEd
uZJ/V31CxgQTcFPIr5IeFj7Seui3VlUmwzBiCv+r2omuNgQVr2/yA5vyYwE9eaWh
a6L1s6qP4C7PpK46ax3LEu7Nv33jJd7cWM9XHTcvePnm1mq2EV3o1dl/LUqj7Ujs
4Clab2wCrKVTHVqhpLC7ToOqjJTBbkVEMYC3SpLYZl1cd2VH4/KWTkZdfFpshOO7
sAzsnJLIaWpjooQKGM6vzWor7KhIBW/smdw5GkCHOABLgqs4+pjCvGMUMugw2fqk
KM+wPCRg9pDRF67e1ifZRJ2PFKRRsTaYxwDNPustP7dYp6YBpRYJ4I2gcOtC5F9I
eKpbhqCV0TR+CPfP/5f0NAEL0UAnx8lI/8boXvDKofx4b1QVz+OAYKeYbPgSPz6s
4bBum0riMfSBHuFyBrv56+B2gQkxR1NnqYsV1loWZAHfsAwxCnze/gZUpnKl8zQE
xI4XfpCLXQT2VxFlzF3LWSQU1EHh+9j8O4M1/jGcxazm505xp6U02uemWChfZ/Ng
V0lXMg1ZzfVV6lwPw4sNz/s5x5+kqfecgkbAZjVMgjkt0EthTd0pHyI1gg3HRg1/
hcpFK3BOdCFJwhaDW0O+2qgIGASPzqOId/SQxiNdG6yFyekBt8qQHQriEpOW84Iu
rhlwqpwfvtQEkOkN6CCgvL48P44JXtOomq1fXhr3AO+m+zJ5oobkzyhm440I6q93
PwpXBADEKv7UMdkQgYkvnwRpFV2gqmn2+NYR3iRGDXQ8wyA+A6LAanxWWHeRkShp
q280W1D4LGtbNdKSi6JSUktj28+MozaU1DLXg9a7qY5dCGmwKJATA6jcPFeNCy6t
gYaPp2k3UwC1B+iBJ8gBGYpwuJ8Y8aJuaZ6zOsTCk1x8VqJ96WwIn/Sx+XbodqFo
K7eUkISFi0I9eVJkpkYBR4ndZuBS+sCqDGkp2JqIrj3uAWYUrAFxPW9GJlOaEIQs
yWwIRRNGiSWtbJyPU0VcrLVac6MEh7hRcK5afd84KtWtJBkDSfmnWcRAJoHqwIHE
Tp6WexZFklztI93PfF7IUg1OzVm6PxsY1bX2tC1C1yN4EgtZWSAZ3tFzrQdZiX5e
7HflyLQunSSn+yGOGhfzLfwm1FR2W+N4K5iY/otZF545xQI/CFgFrWa5zMuOh4hU
1nJAlWM6pb/5mCWBwhkzqeM99f4146ePzBV4+E/D7u03mtuLxxWt3lA5zH8Klo1H
0EOa6FT6fv3I69nBsyYr0O+YsPc1WQVIe8XK2MeqHZ8psRYbDG9f+LDLf5hPGHmk
Q8desPASQHezggWxI5pibuTKeCWAhb2KRMO4EgOWaxskOBcIhp7fC6jjOg9oY9AK
pw9sTix/sXqr6uDxMPs7u5/4yGQpSz3h8CxHEFAU5XF0pKxtqQOQSwlPkWTHSIst
3Zicg+WpGITZ8A8l9os7FmhmBsLy/F4539pqpkprFbyEDaFL42dGOncCJoVShxml
57Wtu3lcMxLpEh79gCZCsx/WjnnuSRaMO7or1vjbq45tJegMan5bzhr6S07KMpgr
x4+7yloc/77b5uDGDopiDmfeU7S4slUsC/iT7GY62rTW3Spqh7Jtq96J3D0aQs3J
X4ZX047PqCtywpXqck/FPbQ/JVcy+o0CPnKbQBhOmOdprt4mi1bUj0oyyK0eIyF4
rLADfi/IsSM3hu6aP/Ymy9BXPNqEgmGsJvnt5CeW6WKKXTdDZ1oNblzt2OoW1AkY
iJ3rC6EmTPkuq3U45+R3wRuoQKJGwNqPwtvePWeCAMRqaMbzr7S94KjCVZuwAXQU
zSlKl94iGoMX2vHAZqlt657r9XPjKvcsemC9RO40vM1aqvSpG40LJmdQmOKxSVry
5Fs+zhBMzDiXVRg3Qe094qZmkZuP9g7I1GGEtEM1Y9pyk9AABmJ5as30GYqFfwtC
Lz2C3Mk9UlRLRlYsViHkjXolBzWKS827f1Rd36BspRB/iyTNFCPKZNhg4D2ydUW0
R62avlxTUGaAX4uFMV1aFhIvJSJbTgpcXO5mFgexLwkqNoGsysfErLuiMnsWTK4H
Cl+HUDD97FCHAZeAJMmkArzMNT7MKUEMwTLMaO67jxYOid85R+3ulOgRh0WU9WZ+
0scDDlAw0teOzux36swPySbyO1GaaUbV8P5yiah73hSOMVug3oUirqUyenXcD1Fl
+B+YKnDNmRO2lFSKBbc5gspEd08c5wLNcnOi2x05n8BUnJWHyBrO1kEgdzKaENCV
mS8EVadwKg4z7tWpm813+2yb+vThjfc8pM2c2o6Auusanqej3oLuWtF2TSR3Z4LW
Y/bb2dZWDU8qWF0XrypgLTa63pFWDwk4QgbHUsJOVVfmk+oVGQwFlxoKzDSFYiCu
onCYzGLxezVXmFsMAAtO3C4hX8hAM+h8MSxbqwc2B9pgFw99c62FcPbD8Z4QHYkA
gUTVmh7vjT9RDG1TI8nFcPjVXOCtBRyb1pNnzk7BgeBG1KgxfUzHqXN9rtW2AmlM
JjOgTGBGiBbIy2HxWMPpn6/hcUg4Y7IyzFhup834mYEzY3lZ35V0ZuLUnD5dmNYZ
SgZZYvYOEwAMegWy3SO9rc6hn5RutRW5EEZQk91qTgYLjSbnnb65g3+iOfipvZGo
MZrn30iqavo0yrvvpB+p/pwzRQM8qr+gtqER6LN/mYrhcOsA8wfsRzAjrEx2RrE8
+rXx7G2vPPj70K7u5MqU7+EyB8GCMx6l9qz1lHymKZ7ZCMg9maRfOtdLkGVnXkUO
XBRWiKlY2LoPzoovglm8Fr2ICjCmYLw8geoiwZQbs6Wy4oMGu1IcN1KLefN46Pxq
HdGGqCBMKrSov1RECIlipsgrLH8zrNLxNvZZEIH2RPiUcgeAXRaAtwR/cC+MAALT
8VRq31m4atIg4MDf8PdDbW2l+lLooEwpWoWmzg0dErUk3IaHoWhUnqEc57dBUUf8
8YJKVmBlJtHn3FrJz8Xs8nI0ncYDhpolK5sDcQ2YySUaqxSL2evFlxmi8HRHNJIC
/JilNA0KKRrM3OckVif9mqL9jkTnql/TeykV7TNZlxUlLzoyStSPwonZ1iaIJvcE
g7jmJQuvxiYZuOuAlce20zEWLADRC2X3CcIPaOP0ryvRYewk+H4VRosJi1lGwbMd
5eAKS+G9ZZ0YJwKFdbFlE7UmRymHdJ7bOLorsYz5QO1w9NAhVCYjxhtkxXDbHbXN
6afEvmLwqstDbWcTfJDP1PqlicW9dnrIjnUp1hVl06SNO+EV21kAJxp2mh5XfAyL
8vHm3mNijuuWVld1Qr31DJJSIWqSdFuW0HoYSWeXqqRkexx50G4IcuSC2ta1AyM9
UidRekbxmUNreTUZCPCU5hJbYrpmrZfnY4SJ3bZeSQoIXlClV1tI8V2sfqQ59Ih7
oTEElNCzgHcDdRCnmsltesBGwxrXbytJu+/wOzeJr8ksTCK5ow8d5n96hUynKuFJ
j3oZvkvk7mHLkvhp/NoYvCKRobZDDUc3rFbdcTcF9AFJp9RcFaVacdMVXWhef2fZ
R5BmbGTUu7Vd5qmZEqOBFjI0DdcPz2hYZQCUH2O//kob04IRLJMlXT93Wixrqe0e
sREJdCNL63b5IWBH1Po6pjEB+5z7T+aot1HaOAzs5tvu5ZtLwh3QGFN2vm0dGorQ
qPsEkCkS9NOuJ686+/yIV8qrmDwgEZ/Dz+qrq0TAqQdQYiWcFSiark9PwUOfPOdY
MzvOvVpMlVMPoYonyejJY4ckwEET4twwUW152nE9mFydf58ZBJv0CqT3Jm35KobX
L768WyjL7E4qKyyl4iJomNuB3z4ebzBw1KZi6duVYkFgUh0WoKeJMzK0Ij7FuEe8
d2XSGyX7I3T0yP7I+pdTsb4OJvksfWIZK8goJ2+bzV1PlUEyAhk+EnZPFjqJ45Rg
8lN7tNJ3Tztp/X3JsYzx8fBTfREpzyD802jiHuHIq/o9r6zMk59P4zXTqz2HjWc6
d/+NG4ppO9GODXPbBS2GXflM1ERCvFmaRsoFzWvsGoP45UM+y7Rj4ZiIBPvctJpP
mYpgnYbx2NT3+8WbNhQ5jrw784USLMT930rc3/bKTf5dLFEe3OMwZ0XfDI0T7Zbk
Uk5d2tqhIr4S4bMKH4hupvjuWg2O7IkHbXLnpxPSY/4KQUDfenB7gEh3j/Ib4TGM
FoUzCUSb94s6gEz8V1maDrBF/+0pixTvJ6UCAQcEe3OksvfcTd//X0p38M8flyix
OWPNrexW5WmZIemBsl4vV7X7aisU3WIEZF4h/G6q9eusd5nHtmV+7egqM6+6ZjL5
CELkpZIkH5zVz2in6f9gmMtC/gOmzv/p6KtFc7sfceZMlk/YLjjcZVHE2HX2U/x7
VL5e5VRw4esL5NdR4/7ad4L5f3FOIdsRW3zF0MLXiUruaeZ48oHI0rJLAACEYCEQ
gdFM/WXWbmcfyvxeimV949xuEWqHuECW83vYqa7aTBUtnoOgUlT4/u2DFS83JRa5
1AlBQds6JK9fwJ70Txovs4z5rRkHUmilD3HB0SHXXsYw9xBpa2pdgYTxIl3m2UvN
No09TxQf7qXmql5poyDgOsj81Yp1a6wB6+10JelyLjL68+ZgLMOpbHoCAm4TrlC/
dzAXXg5/y7cyeChKkBa4c7Lx6ycA/ePongBi+S+cF37TfsD89Q904op8soA8K+5a
vee5qwK7tYG59Cb4HcoMRDd7cg5IHv5acptM1X73yv1+wDYoQv3C6pT5JI77mlRF
iQPN3Z7HGcnHNyz8B+qAe85VrFnj2vadVDGsB/w1+StZe0RMgQ8G0XxC+RGA0cGu
QxLckHlHriOxc3mUSG5+e2/JOrT+/Jqiox9PpvRxeu4+plEMhW3bswJAYzEZLbSE
98MFoGGTXQFTbu4iODiTcF4IWOMH3kf91GELbqpA0Nl90ei/gdcMAjmc1Fth488x
3nJ9t4IQvRVpcIFF+1wCtP4ZA9KVoyoqwMaf/s0xjEF+jbEAZFuCXhUpVFnXgoTI
n9LThMzpV15X6yC2SpcMhHWgRAh51pTHEfJOaN+Y4RTYq6Z9Pae3fDXVY++LtP3J
1coq97u9BQMWgU+Zbx2LNeyttLbuO59nHXPYaLQ02xpIQ5mgj8+X89vDWdVoLfP1
AMFOFqqehuj8ugRztt9dw8nID9+myQbV3F2TlxezzEpYDKC3BbyaJ5PQvzXOiacp
77wuk10rvzz0x3RifCP94MpRERqp41XJCI46Yr9eDkWbSQKCnT7SfGGkpJAc80Q5
vJFHeip+xPChhTE51mwWD0BjRV3p5D/sE1DZZB817oReCJdfKRdolhOrkSbtvaTB
figXPG3HfeMLTcKxp5WzlkIyhClBxqnwaB6Ws45Uc3FXmF206uMvLnoFVePzK/T4
tJh6fuE7jxeYnru4j9YLsUW8lW29Ep8agbqYEBuGM44Y3leRkXOTS6c2ZaqP5YQ3
M5v9HVxJCcfy/AaTc9ZWZ+Skytk0lZ+tCzEyC70oTzE5HOZS6GMUUBLj1TG8cUpt
xzEvPdKAGLfOpDUSY16hlQLGYC5CbV/e/xJewiFhO7snBluaWKl73sIV+8pDtr0E
cHroqmPbp2k/6vaqHCzJuAyDy35Pe8wHFqKnZ4zlLQxAlCSJrVy7QxD5+Xqcbu5q
cv8DZO7Iot+mTHvb23YWeXlt5cohH7xwEwk3+GZVRUbygumGY6d1JrR3U+mrYXxk
cvVjFcMuVQN2tYHeAqY+TuGlHzwhsWWZ8ZZSpZ893uosNzp/u0SGA03kKOdQ8IIQ
KFNbIEyeNxZmxSY7pjOZ76qWTdUhd+SLRQMjQR8L3LwQYvPpbyHa/YOubJFXFTPl
cw+/ux3V7Qa1eKxB+IJLOD+cI0JirZUPAXfBC7y3v2DxyPerJjxCbsVs3z4w4Fm/
RdTqWw4b3weJ2/btc8NacMk46s+ev1rry6uEQSw1B2k4SaOr39Hij7U/APfn6Lic
wI9wmzHH7vFS9HwKyfdtm3ZRHHE/i8+8LEyV8i67FGnTCZX8tVLAiX3jSkK4iN6s
CUPh5lVTFu6r39SG+sy64qYbOrpnp1SJgQBDNIFjidusQX+OJyURSQA2jn0ti2+B
mtha1EFd9Z5yjBWUeKBW727fg/all2Xto1BVzNUDIGasGieWAhyQd7oL4LFH8zB1
i9InmdZkzYaBGEYgMMFdkdcyNEcaBvQVC0qoSbByyXBmPBW+e4IDwStKktj3wobX
aONwBiYIxKQz3XYQCAkM29uz8sYtMvg2AD7Q3MHNTAyil/VJuKXV68KSg+XkvG3n
WWOOT/sNM7HskQnUaE4XBZR2bOhKZgl5KTvd/0Kwg1EI1kCRd1pp5tWLpvHgOZGc
mc+rOpD+gIIucx3HFbeAxlJdLwCYVibkkHjGhKG9/D8usRiGu9GHrGZxFa+T6rMs
O2o0U+rhdpguefWJluGu22FGyL1vRl3efUCpY/y13MI/xmt1LUlCvRcdphYvlw7f
6u/JUexpTUoqvR1oUprAAgLiZ9s1Lq1qJcwayHvyHSto/6vCF+v1T9yBerFPa1tx
S/+OyilmpW+I5rkWgQe5bBUEp7ZgIdIy6u7R9Jsnrdl7mqKdao5mttNmWcwyidZb
gvMB+MBCQAHhZj0ab+iK1a5Ug/jaBJlAovgNQJWotlF4fmSr6mDA8cqhpR/CK59j
wvMUXuEvUbttuh412f6E83NwDgGn/S6/fVyIWHThwCntHHNG8aYJaSh2xf8KCmgn
o9Kp7rf41Hho9dLXnHw6IHGNVl8OseJZ4toSqkEziM3Yfd+o5nONFAtENnFWff9u
dgurTRFXm5rxv/17dcqDTi0R912CqQwYGHSaInplBodG3BaiW38jaHBVRbOPeffj
Vd+2a1mBcn9TikEEan2lHLal8QyMKsQIqnsyYjbJyJLezmy+Kpvo7M2J5WKX5+Lz
fOVA96adjez6gAj70ycbffrS2wkCeLF4ugeFjtNGTyv03bbPP4vCDGoSUaYJe6sE
7RnU+WOF6Wl9B/QJd4sl/2LeIAgdRwfvpX/3UOtlLCH8dhUAmiQafZQtXP6vT0Ha
jF3nYHggz5qDg0LAkkuaTZFrPe4nEPaN1gVankXAbkLzMUaYFWEhudWSv+hRB574
RVZidSGNWNGT44qmQ/11XPkV6hte+JknTRUNgp+AD7lhtPuVXmK59f1INLZWMDG8
djyXQR7PRWLB8ysqiIg8W2I9z0igtiKclBEG6iVT7SbF0Y2+qlFVRSTWBG1rxy9/
5A8nt+TBW+VSex0ugZtgrmgKUD1ZX1h/S9Hp4YOlDQbJ5C+YL8j7vHJxXhjqnLwk
HnaNo3ntO/hk/M5tl4D/3kZPoQx9EplIA9H/4hUiOJpX8VFpohy/RFVK9u+AIPEk
QfjApDdutgpRxMuMeBy5XfaiDTFh1yoejxOwiHFVciBw+bm5Sa5V5uDXKKMhhISn
VAQijTB8+QWCuGFt7KhIl+ToFa/SbQ0BUDzCPg4LTHUxL9ijncUv5M+JPfzHvfw0
2FAVBgLKol46yvbr9mvPWi8qCcdfx0jRcnxqHm3bFe5rP/wPnKfVSh1w38cHH4PF
u37EeqWm9sPgPrBpb5jt5yWKmq9UHxUCXCHgdYPU1HIkvQLl9hlhig08Fu5ynC34
udZWd/i3gQ3Vlz9WP+FMMMC/v12oqcD+VX7H82Xi07gOnwY5m9geBLmTXPXUUNBf
H8Pmii+688gACyYhLbeVu7/OrC/s6lZc8H/fVeTOzzaMtwnJ/piVMfi2snsQl/Sp
3IgJBBz6U5f6tQoZ7VKy83m35lhstud0iWFUVzTmqEHy8r5hws4iEAYfR7e1K1wU
J3v9px3gGmjSh2PEKN2Jt6up6qcybbwfj5EKKoa5n9tKs82W4m+uRQnOAhHAvKT2
xFUnK7D/rnLrz4/bGpoz7EYPHoIqwM1GXzc5taWpMz4kH56MlNsVeR8hh8TCZAv3
80+EPrv0zMp+naoPQ2xyYlI/Cmz8ChIG0jx6DKecxod3QMJmcOl8XTZtaxj8KU85
5w7+pdmSWHmwW7jS7eIqEfQ+4fHkza/GRFqUh+NebEv7hlzUzwBbC0od9SJLrFD1
xbl7Jthq0WqbJaghmZPg/wjGM31vccvCtareuah5sIwlvl8Q29N2dpVxy0Ss3GR6
FwU5X8g+tk0Nf5n95duLjqV1SIHgns1eVc2dvPoTrJV/l28Br/okWXo2yVqMpmvI
KmNolAuWXnW3Kih8p6O2ym7gPat9vBewC+ghMJvVTqVFupULoEhAubLHedxRTxHR
ligIMWA9hgy94RSwWEhHzUrHxK2QFLCYtgXH2dXuDEkXAdMIe5H5xiYG+6u4tnZ4
iJzHRJVodRcCrAX+Gkp8Qhn/7IEeJzYCdEMoGSndYathm/qIORsimJ+mKtaMxEA+
z6rFjeAFzwATKSCyg/Af+bhSY0pAYAg/uW/SMvy93zaFE7gRMJd+rdGOIXtE9JU7
/QvufOoS7t4a9AbiUJQ4gTyDqMFtsZbZL7/+VuCMp3lJ+T42hvXxKBGL5xpTpvb3
uzfHRIdXaY6M5u1SkCYYdQ0/A1fQIzilG4nCt5Z0V4kAfjvTvsTIciZzHgPafM4C
k28uldvwWiMLVaJIPpNpvWkDKyAzJLCgMg9+4p3EiOtWW8dOKBv7BqfFqANLvz5x
+kARdVM+ce7So9XwdZQ0AmekFWfi32IFktSgeq+gTHg6xwL/TWumnGqAHm0C+fzl
BkQXWfleffy6IKAwciBHViIIU2cWkCP8HHSeNbIHDr/YPzsXNPk190guJha7c18R
KqntSk0zgs2Co80ynusXxsrgERfC1Jdhc9h9f6WSqKGM+ZsbBicMo6gNN/Yexb/d
6ciZljVfJrbvtN4b95y+8REpX2kyCGv3jfGIw+NGWam6VMScBPnB+XSUUDPrX5Ge
K5KWDG70/xyt8Zavxa88uP9JB7Db1RL9+u2r10aZc6MjsjXxLQsMljXcUHsTWp5K
Uyi2Xr4+H25PYheHwqK1jxUgJ8TSncZ4EKb3L0SNfFkoMabSJwpskRubxotW2mSQ
5xdt3gIRCM1cI3EcjWs4CHHc4ky3oaN2e7QVJh5e6DF4vMvwyof/Lb0LEc2w4wwB
bpQLQTc36xWocaRaQqIIMAB1hgvKwPXOlcuj+kT+BRZiJL/uxfZVozGiwHjcDQYA
SzdMnGbvJDjXkJW+zbrjYtqqzOCQhAXPoiskpQBGI/5pWhk09A9VNKYjpaLirgMX
tSP/UcuGeNXoFxocY70h/xh9xTl5caqVT0G+G5xlj1j2/5ltmAya8fRJEOOoUnBw
U0DdwlSAVzHrg4qZLx3lxZVZJFhVwh0iZLzCV4BrJ4vLTZmaVW2yyIQqxeFS7uxC
hvJdwhz76HPOUp8Qmchi1VQa+g1RSxAeRoRpcXMypAZE6lQBs1lrgjOKIu+EtHfa
Yoqo8D0RN2J/VIVHGVjY19HkmU+DKkOfcCQPuN4L3hiq/ASnrK3ifSH5AJQeYK5e
2iAG+w95842wz/2mSvVo1prHGQTuKBSG/VuCc/a88M631Qr7gCQdvSUun1z1XggR
kbKipWGKV7HUvIKBuz2I9riOmjqlLQc+oGK5tEa4UGeui+si00p1iLWWfIlSc7uq
CvULEpsI5DZ3qjUN6nKXKJOx6GyiVzOXUcjTihdVLgn+K2mG4Wq8TxWs3vp2Fd5u
aag2FMIO2IgLJaCoh4addYmgKER04PuS0HOYPQUvSYbEuBbShqbSr2VlMYmH4ysA
NoqMm3fJhDMbfAIl15k5i55uXkCa30UthJLsiRU5DHlUADz5OE/oxQA4ZvEMawn/
rQ3i+MmiAbnGwyGQr4fexmp95PhEh9PAvRNaqc5oPEeDE6PgfwGF0TrLOCLvpKop
u9cEQ+vDeW1PhMu7xtgWUJ+ol7MeDm1y7+LEWhgWJn/WfPYZu7o2959Rpa31ZVjL
5ySpXsIC1jfZcdmosGe1bCKoDoP6oaI6l3TGWXPZ6AbmQd6LsQYj9iCt/3gXemhB
sw+H4k32UJIKfUgL/AtedCHzdXWO+8cLSXHghAv8Ww+7L5mzLggg+LmRa8Q2RnQe
1LYl1yAP3NNsnOltP1ztFL1DOUfbsCsrXztRaApZ21ewt+rO79Mnb2bcM8vpURWR
ah27Iy0Yog6XRia4JXH4QnLWN9jndLsh823fZN4riMX7yIp0O7Rkh4xN7DXoD42u
fX43ONAW9OKxxsb+EHaPSCPGD/4iESRKGFk6iM48EwV6QAay160g538mVUzm027m
YjX5d4z57KozZB9lCo1CG3tqmlxLJbAE0NNncLjrwDAXmUFb+gi5VTEHP9VTwjnp
LG2BgCunMUDj8EEzZjwSRj8dtjo/9phWq6HWdjp9kSkA4bEB6pg27cJT0Mm10Z5h
yqobgHoeGZdh0Cinr+eZk8GAGmo123g7l9na51mA+O2XRjsFzfHO+fFvbuNfFREW
mCM4axjEFkK+5PB9irrfgfnz4Snge5T0uzetF57gjT+kAhW48NKonSDFEgAinD4h
pKAtrlYGrf5KE3KFVa9RzND0a9puigyrL+h3LbfZYCePcx6WhzB34B4DT2bXsUxy
/LCXLTvM+0yUFkP2apNOMfe/UusAdUSRnb8QL1Fx4nEedWCBs8oCRoplp/cYOn/3
czJLNVweTHHU7QEn3aK6MjmVr0+JnCpPTnQ0+Pg2X/s+IsCCOnPUm8iBeZTeeTgN
AbYw3pm5wIy3OMAK07yFhD5yrUbJZ1a5CcNUFE86eWTdSmrrcroRBf8MTXakeB1e
rlyt1AN1Ra2w/LgMMrLdDW5Kk8+kSAnF1QtHl02WQwiFYhIprqhjYrgf5hFJwqUW
2Q4Vco7LViOy/lz01ckpLpVevgK+0VU4/GSedEGA0A565kxGnPOij8DMpuFYJJSe
VNBgz3G/bEHqClk3I2NPAxZZmrZfkz0O6cjTIBd11dbj/RIHVaSF/iQKkxGyptRf
TZfb296gf9sooOiIfpPke9klyAidRvkSqttAc6gdb8FCPaXH7M+2coKW+EvfxPj6
i197R2j4la4pZynSxgv1caPlIFaBCTUNR/j2rXIFPBPOASNjIDmKLWIpD9OSykxU
qiLimncHCig6G+U3CLP1DWeah/rcUNyW3VLF2Gom29x2v7u9XqtWa1GWzfjNFLfe
4BxZFDtWg19c2AngTeMD7w7ZPhbTqiSdfM3HtAM2T3Vv5bO+Ea5UlAW+xl26NyHr
objlhF6GEs3D6wQ+hklpLkzWRxLIwYCWpdhlYzQ/O4Yuj+U8twm7XSiFJoQGdyVl
vB5UpkEBpcCghd+E27RAIeBfIc8HOxEwfA0ok02uxAs4iRVnw4slX8nw6hUkvr2D
vwTvk1PZWXFTdSm/mnN6r4ZpXReHhPcV0x9Kh9WotSfRvVZGZk95IwjWTQ4qkQtS
vpwIkXMNPbuW04HCJTg46vsHOSMSDGIVkLUZZ+1ydONPiqoixv/CQ/wo+HpNhUz0
sP4ULkI6KaXHUujP0vEIr0WZmBjvoiSwJbkgx7kSCPbgGbkcrTtaGsE9KG2DKri4
P63YIxJezColW44XYc9ge0Jv4Lv9spJWkwIb6vzSBNqIMjFBh6ZFy3h/pNSJSLT7
oi/TzkHKATzhMOPWAaukQhSZK6sdS/8oJ0dd9dm0XzzwEw8toqphkgZi1tYpNDkL
3iwjZ0aXyFrt4ptxjHC/FWWB8H9MfChhMU1DS7g7ZqIdzeDjn12qa0U0ULIXInJr
t9hyCKNzeS/0BDQUAppWDTsFdkc2c5mMtCgOJk0egoDdvlJF4x75EqLJXCRLLtbo
vkZUJm2dRS3CthZySEOSE2Ye4/XbGZPiDrBWNfPdJrw17pw015CY3nCqw7EtHenC
+/q5eT7Fzqm5yXL9hEtMP9UB/i3wXKdkbiTSkhXvGi6FRydx5RJYWkEWThOqxm1T
cEsYtx+/WfYIrZ4i0UmwKyGfWzEkj/VpXm6f75hb2F3fr+Qy+DwNXCJEkelx9MH5
kRKIehRA4rfE0d2aZs5vSWjZL+tb2WZPgGWBhhL+GQpg03p6pP3iVBfbCEHn8TTc
iKP8jw0mgLHQXrug6wQHlbH14vhdmebjAE5QLOWp++m1SAXcC9OF3Ltp6gmR2GG7
89Dk3zo5SZL7U25jnmaC0L2rqhaCWHVqOj2QFIG26ahcXcTEVuovM6KepilNuHY0
eODUS9RhwvahvEuKTgC/IksnNWa6zX3HXJR1SVaWUkta2KwUZhmlEekmDBWhD87T
7/rQbPvDvA/b7hkD4eChukiHV/ADfv+5MS1YcpCeuMIbfasqe1Ut/bofU12WE/uh
wA+2dlvi/7qxv9ng7NgNH9x+HL9xb7CQrLJSk6GLwkKrFqX++eLOC+KSlzqkRusz
Z6rDsUYyjpLdT9LxbsKQIxjIPXUoBi16Etz1zcqKQrflbwbhq+mleNv3v6LcvdaN
b5HxLiLuFl7tEzCwPpifI6ECwLd2bRaDWQ7rNyZVjgUZ4R/vTQDU/nEIJDoO7Ym0
Iw4WINcvQNRVFaaoAE9tIwabuOudI+iQog5YieNPlVA/7Mhbm30Q2cIMrdAS7Y0Z
y67NSmeYM6d6SpG7hVSEFMIeCMancidZWTfk1PGV8nqisBTreOVVhJ1hPAtvvmhV
FyEzXFm0RbVfVJ3LcTYkqv6LB5MHJa7jirH82Qj/CuCbDIhAgt8L4fnpNXWAhOXw
fBoKLVzshXLNLZ3pbVP47V9dHhlsMCIDKilcSDTN23uoqUr+zOkxsoKW3A/g1kSq
pNZpQ2vjyGFrSDRMTKobtmH+Q4VmvjQk8GSs6qL2qh2h9MBnOdGOPbOBPs+RZedG
f5wvkvPWQQUL5eZyJ7MEY0T+hrRObIkDnIaTIf+QtY4Jox0aZlDx+chX8MEv6TMR
VFb3cRgcnMLDaZGDYz0lSO1tM+vu5wMeIGp7ry+M+wgqBiTkvc55frVV6dKzuJKG
9q1zeDhWHHj33dZF06jIRMa45tc89u1GeO11M6TkP/NIo4hxOUaSTjsVwzDVd5qc
Wb+ysfNJhBPxm9q08Gf5h70t4i+V5rQgbNdRaWbpMNrFy1c+yEj1fPUFyXYwN+FM
KznKi67dRfeCvh7s6JOlcdHL2oJdLcsOeLJGkTMakei6zM/06rvqfMwk6FNUEexB
e45zcKPfHAD2CMVZxPQSDi36f/u3Ao1UmnpwNObSgAP++pP8ByMdXkgzSlHbT+E4
o2PEm+mi90RYx3JLcHkqZhC/KcHDndEc6yn7eBqaKAz8NoGyIq/nDAm4UGDzWPnA
iiTNJoCgcyUquH4h+j3SJs9XQZIh59b36/1woyzI7X0L8NprJE6l7fCVKPnlm4II
gO3QWj52VIf2elREgUw0KoK7T+nN27zBo53AgYe3jAdmL+CW/PdB+FFfpcTpm3pf
yL3x2ODlbqpFVzqCYam0cRE3BcQBNr1i6ACz4MA055VPlj6hCrhPqw1u5QX2gjH/
mUTF/okukAl/ulpAQ2vMMiHu1cSc2kGjyQhAT1cKyiBJN87ISgo5ceZY3AqV6Kv+
T2lob8H0kBjMwnxs+yuINk/PNHQBrvpPsUIOQcwRfSWbcyrEiA2f4O7tatSzguh4
bh0Omw+ETBMotqVeVtPgoWCJ/BnLj+471v0xxfsjSb0ulLWgsxdu/Lgb63q8pid8
e8xtmWoldy5lQjY8FfTtcstbPmiL10fPibvad9PnDNnWqUoY5W+qbD8bjgNVcCKb
G9vqT7eEZV3zxUGeZAdktKiaQJbFz4XC5bnYCL4ilbFDinfhN5KcCAV7sgWxhSfr
VvmqCu9KZ38Ib2EKTgLsJp8vFtTwRz6n9BmkeNwZvrAvOoxxAs0IUT/LH6e9LD7e
OPmM4uH96AUTUyvkHQoio2cVjODBY1i3VxPcmA/9tw3zDZxVBYKM1wbBJ+zoHkyF
AAqujCFS0/Hs5OG9zttq8z4RBZjoyaEBxHmCwg2Pdz4K+YNcnF0QB/NhS4gFCkuX
xgjgCaMng0c672koTau4RVqvib0MGk/EqOa//uny3iMGdSG3C8T4tzpacgvXfhe6
3wUhcv5rKLcaUTe+Al95Yn6UK2npyBnbMOd0hhQ7pszLd8FU6r8sf4ET8oM33GT0
qxWh9kGOT1oqDqlVvN4vGXQItg39Uie6rNsy9jiF0sz+6WPuHFKuikoe1OyW/EeL
ew6LbaO+mRugOD7b/Ug+7/jPxpQdbTrnhCyy6QAzc1IVOUrt2u9I43XvC+S0bdvP
YZ86li+Xe2LrqCebgXifi38MlTtE6mdf1C6akr6fUwlMgvmWGi8yAToWKAnEhAVZ
+AvnePZL/rg8nmB4lF+rYHhUgGy9AQYFpkpDpwJ+WtoMRNgP/DuzsQwwSM3AGkoV
U/rnY9TEz49obr8CmbN58hSfoYrRFUAolCJNdgMrOFYADuCqy3rHicMQqAWaqq1z
MXt4Ao3ZY/1OG+G1JwvD7xOCq+ddqm9ardEihrKYk05d0H8p1S4eIfwX/fVNuNm9
mB9e/9z4Gc1mOT32OcTeFgt2GmMO+leZ7CGCMSDHF50Hy19EI8SFbs7HOQPiiV7Q
AUspHGHFf6FQQ6EL+SenEKgVTSebH78nZ1h/KNuYv8IIHZFoqGmXIgTTf2K2r3vw
UZA4mtL8wnOUYF38KyHEnrgVC+J2B3iT6PK0Nn9XQpZxcNJr7GINwNApEQ4CGnSa
KVw08MVHUTqvZMYGf/C1pUg8HJAbqkKFp6RnYFxlLhL9Il/m5a/WpuhIr7//HV7T
PXjD4WBDGDijk0rjsHTMLodeacOLR5QLEwy+oobfaQDFxqKbjHWj/9yapObJFjZn
6OCWFNdZtePMjTqXiNdzjy2psQcRQtUxmtixiTaH+k6nULRAcFCIdXGBagC/TiLk
XpF+Uv9XKFxEBkChH0SsGZD9GLq63x/9Kup7mPQlKipU5Oae47ZBPcGRWRn+hFCQ
1ZhGuqKMQ2xoy4ACq4dne5GFBiy+sfXiCsa15gg2jImlqEQSnV/8hD59jENDI1pK
XsnRZH0nyEirZxyNZ0OI7fFamzrEXBWCLh/k5XNFfYcLPYXhGAUbp7i/tAXX2Dky
ixsa3ue3RaOw8+jQi3mwtBQMGdrcezHEqZdLysx9/nLCPfXCDfKnY0p5yUCdCHnx
s0fr6UR3dpKSCFXzvGIVJPam3e1UDemjJjI5Vvp5zyN6CjYIyl9haIeSFCpstBNu
25O9mfKVykeb/+lHmMz4P8Al9K1/U2Pwpox8YoeqLyoTWRb0N63+QtGRV3m4yukv
GzywNwcS+Bk+rBi2jeU+cTvnowvCr6lciFEx0evT5Gt+q5NPKw5+wTtIdrA9xTET
xmDJ7N7t8SQAvx0Or84e6ABu23MVg0Cn0zT+fpiyEkt77GMKoSZEZhYmaCLr8F7h
2OJn1lhbHjsrGXAhlbe/zdt2GpPxp6yQDFKAt66T34KeX8rT1CAQ6AXK87rbAiL3
ZDk+MFRVl0L7RfH83quu6/CVZhWHc1kDgUvVhLEFgFCBFhjhkm5YUb4fEWWOCeS/
pv8dEswYUJYRedO8vlW40tGJE7t7IXFrTaE8ZohZyI7xJlz3c1NI2G37dqQgnKUT
OaoZ/vH81yvoxxP5y1fzuo+WDHlEnhM8/yte3HB62B5qK+t29ZPTS53pvGUC//eB
VTkZKmAPhDszXZu09yFm4tXZwZZf2GPUqOItTnzuHRqwGAgAFqWjcZywM2v7EgZL
EHla8jgJrGgZyP//4qKqijm8vTBuHb7VVbmWV7LljZ5fCy8HYWoZndzFhhqC1+cf
/9FzMcT1KfMro3G0mqZPhHiHemERLNzKndxKUGF5iwUFt0j1qAsi71wg95LZQjaK
VpFg5GOuWYsc3deDXy1CXAxkEXGWuAJiYKDFv0WMax4Ts3qrF8C/QdGpSEpb8XoB
AbLgYbEMXaRdfDAVHrW+dV8jAmPcxen5tZWASsLMjZQtQQJOsxd8oicAPswTVe0H
qmsbLuoVmV2US33XHoEDft0uCBhLMRY8jekaaFl5+5NdT4+MeHBwQPuHZsyYk1w5
u+DtQrNZzo3D6wyPeOiyXRCo1qFchGsbodZZDAit6mPR/cta5yijtsinShVY7ZSr
9uSxIDp/C6xLAOJQhHP9gPjYWatPDfo9R7Whsqf18gy8fzDfi7eOgdN6oDwgcHav
mvnUmg/EU6I2M0qGBDLfFUvI3NrjHeEFdcfTaLj4z5297gdWdNGMqNHWWIVD2Oft
lb+YPY0nNTQ/1843S2lgphjACZHLMy/dLRkbpGwTYZ+AfmWEk+vKa6ciqFvh/F+o
TcOfnxfELTykG5LYgwaTwAay4uw5js0KRgDmg7KBizRdL+V2ZlqEA8eKifkP42TR
L0p8kSnlFM9qYv99dg1mTMBn53lt5o1WtT/t5qotVUB4hAoiyieYdZW8ymuSW3hb
/PEtfoxSKesij4neRQ+GrAF6Ct6gvyqWnhS68sLzrRJoh+8o9IEaA+cJCVSjTO3B
q8IK58MnBY3i07VW0a98V1FZ4KmbgIZlwO3uySPlSraYiM1ihPBojlk5fVKuI4Zs
l8rF6LhGb2/z40kLBz75DH81yyTP9ZltwXkKG/Tnn2Ahn0ilQNys/61PTzedS3Cm
wGNtZ1JZeUC1B3/3xUkuaRZBvXs2jnxQ7WD8bMQO+TUHMDqaQw8+sSXG1cL2FYLs
J+2zUpVLK0xPQkTuSibixv8AG26523kTKgpfuu/gcAjS5W/5gljXmsPm+Yp0mKTT
bIRMHDYo0BMTdFobu5V100KRx9gmoYUUu2fBjnmc4Gx6Uzb8511zRL1xYUM6cmhW
JRf0Mssz23U5gvU/RcPtEl+t2nYX+PtCX3vO49AwORMWhtsqlkhdM1qIZKPyH+CZ
EczAc0FSyNLj3svYNR3pS9LYtyDcwdQfutsKIQ9M2ZEXq5PcSPrv+ggSXNhuTlOP
lfanphxT/oCXTzwMErKkVvQOxaEzFe6MbHGrEyH9h4Wq7xxnTecDoSB2wr5MGFga
s2w8EVumNVs7P4hXZRUKI41n5PykZhqItrjjtrk/6QAYGSVFqAiCDq5AnxC+lpwq
t7eFhw3WcW4AJD8SH7PBuHAK5kVYYqmcRd+Yg9NSdLF5p36zGj4Li0K7flr+s0ca
IQDriQxgNJR++lf/xIfoAFyRG8mBDZl2TI7zXfx6sU1pF5yJXnTz4JFONMRV6EXH
w6d5jIkPAykc8SMRyiiTW0wOGPiyMBK2j0mC6281y2306xhJ4IflqPv0UEBHeMVd
CzChioCUdGYgkw+OPEEFNgRxJJZC3q0kGb3qpSp0gkRivupACxDeIono6KWWxCJw
mZsnLCuiyQDNgY8boFidrvsYme2aLWpfEDOvkid3esfjOxyJoe9n3MB6RTIUqloV
b20SP+aV4mj2CxuOfCyG7/JuXtFNpI+O1Oz9CL3FNaXSjgACs2icR8BSf+I7u51d
ZHfR24Qk5hnceVD/k7MfDMabtay7F82TunbYqz/ATzT+qIWqiDbW0loexAsEEj2A
OBJBr7DZ9ClnXF2c3mjBaVejT506Ux7ey3I5Ay5uG9sKJv9KNxmGqFXr6AEu987r
hrqZXLC+/8Iaaj0nFMhztJh2i1CMfNbTY6deUJFvv/vnd1TNiwWTzJGNw/TNeyPB
hX4rA45Tayly/8dqUKI/mPujf93tyN0iOhqcDzmpXE41FEN3efSTV26t2i02v60D
zpGXor0mz5XHjkGc0Sl8j87xnmMFg9/61D5gRqyJv/KInMuEIAoLrYxY7Ab4xIAk
eN6SEQoPIzg0MnHCnoMwvPTujanq4vAiRlieo7LDNU8QibOQI+6Jfs3k/nO0PhZ7
owJvWQJV2vziKUGxpmkaw2G/CrBE7GZGWXpTv27OEtQJClGUthGC6S3trt6D67XJ
8RRCvmcQGhNLq1rC0c8McCQJS6Dfa2Bdw3fmumvYxoKB7GDT1h3qbK1Y0flzAg3a
D0jGpHWwjegpFtoGLNg382nNkhR2pZWhRjaD/Y9f6IXY+gjmHC8rl83p/xmTr+yg
m2KB/wxoUTgeemjhu67YoYXsvkxo+F81Wf41cfBV9yP5rFW6Mzwn1CVyAhznorKJ
jTsBH4vu4uytypIbzDanQfyMgle4efNfHw4TCrkyHrjqfqq97+Kwg59e5bYBJgtW
Kh7p4KQrS5ru6VNzdZVftHx5nTEMRCa3Ub4OVuoPdbcCMwOapSSUQbvqPMMPxXTN
S9FdQLEfUYE2D5K7i1CLGChcRxY7IGymcZdvTRwe0g/GnUv8vGKcc1EVbpB+oAm6
AzuaxVuAJ0ggu/MicjO0aoIkNoOXFOzboH6k0c95gfozAjhEZ6419vZ2+zr+QaxF
iAFyM44sL3NQmUWGrWMp69wN6ZAPa8R+70UHYXwoZUzS/pHF/qn/LXQi7ElvRl5P
092K/8PLiGIEn90oszsLnDfcVmYpq6UI8aAEKmlkXb6tinDqkwOrvpfSezhgdwOt
OgaMNPraNqqbF5hIwnC9sQTw8fLSqUBFOn1vB+EQBvh0z8rdy1DUhv9/ULa+v6ay
X/fwo0pizkBh+MNk7VynWwdD4Gsc52Gc0Ii+04rEG7qFiDai5LohYop+le8IG466
5ffcTdyC/+JYT/d4qU7dmLbyJ2dJJ2LI6bc+obD191WWiKYp2HvXcQGUMuW6eE9a
/D3VchMwjOWrUYOvDB3n5adljdLXKAxHB/xKga3zVf7X2I2wMzlJKF9sPigV03B1
lmHgy40wMOWLRPAlwrDaGSj91YDJWL9MxDqfqDSY1KQfEm4htJwR0FyKJdlE7O8T
pitz21+Mx9Mk4In58GkLibmE/QUTPvIEOIJjJ6IAkdUqNUf4PGvvn233SKJLaI/z
Knfrx4CS0G/2MF1RLBAhjUPMcyEkkEUygixN2S3WcbQSMZ0bIkkAp0ZlYR4vpUsS
u4EedQI1SGtB/xLHywHHi937NodpSWMKxv6BOtBywuAM18RJh+a6Mx6iLlD8llsD
TioubamrH5on3GjiJ8lce4/NQYbkSwY1LkQgAxtj5/RqWJ0NIRXA1JqSXTHxpd35
hXjwreKTH5nbddzj9TJYeYXPMqmMMeSRxcODORqfMsJO7D9JX9OvebB+PQcOajK2
9D1wHM/xB68YuVWrrkO7mn/v9wTc6ELattdVgBKJfIpaHvldcOsdmltBneN8Yhsx
t13xn4qU8D9P7fYHwNwz6mwKP+Fl72muUH2AOQXRv10ZubRp6MX50rWZyryY46Pw
fFVwpzxdYVIGz7WyAE75yly3YxN5eY8FHmWqX34V7Ou+3Lx1/dffoW3nfxVaXASS
mpoaq0GJJPtSAgPes1QJoDqC/XUYnvR/1dHeSkcwLZnqoSUprja81M0oq0ZnYZA5
d2LGJUOlzqPEIcLd8O8W3Ln8DDIHQW2ao8DSvRE2M51PCU82BbZXjDOo/lZfkagG
I1DRNpBRMInDGM2iqFHXKRfNnAuXoxwFA3lB4qLRRsS7VdGoLz791IGudG4Zq9KI
hT9CNp6KQOUUsFfGwbcDyVtCrFaADMxa95hnx8KAjd5fR+jl+XVh0tKXU8MB+dh2
hd3A3wM+NYkVAdc4GMEHpvYliCEepueGgiOm63us8ZRZeC9Gup/9Es9ou7535jeS
8tMyuZnXPXl9krLbTmfmgQrXGgZOYqN+L5VsexT1iEacJRpgp4IXtx1ZmLCde8yJ
FfVgORClGUDbD3Wuj/xaysNttGMYDoL84Cwu4V+YOMyHprfwqSX888PAjDJ5m6WQ
6e1XYRrvrDD1zpXl4KOjFAWdSVm/WTG82X9S7fInBJXQFr0877ksG8b1JQlEKyii
b/mZudkXyV3lheL/PFvv2x7BYN7rCm7VBKUSOCSOYPT1tp5b7fbRMRcDyQuYkkB+
qm3LLElKQ/dW9Q28A01GuAwS3lpOrqUDypyroY7F/4RkkzS0t+AcznDmxDOy8h7i
TH0tqYBHpyYw0EWU0qNNM4rS9JsVBbzxNvya6F5VbXr9Ed79Jk6B8bV2XsXi8cJE
lVuY0qE6ru2tbcV93q4wQIsDs3nTm02jFLo8aJspmzjArwdGoN3ZVMMb59sKynP5
3v1y8yNf9phGtnVVYo/987myK+Wb+rhPGpJKYnB9QojeNdDK4mVdY2WTggKhYKFV
dTOhL3O1GHR6NxetOahMrQmNDa1opGMK2vb3LRLtB6j3YuBE0yCSiPlt3qi36A0h
3qMDNKndBk/uaDwv1gl7QZfX6LnVEPN/lUHVeuHup/Tvnt0uD4FDE519dRlnUy3Y
y/h2xSidyTzjVZJFssplvEc9tljvdvCF9ew+BgoGXlhaOCrEPr+/RTrxG3E1nEdS
hxvK0KhvOhWDx5CyBesYsn5cCrVPrw5Ou2dNp5sqBbOskkzK11NX88jiUN6yEaKQ
nF4Qw/BFSdjZSCkXx/yGC9/O88I3VzU7Vk41/TQpaz28x6rMADyVOcInLMCdqCzX
Z7nPESXT64T9cvhRCZbZuHdfMnshK9cyyoByviXRz1lUI/23uCb9PnTH0DMGPwc0
iZoMPP0+TNrRenV7zR8j8oBRI9rE1LfJpzt2Az+Mvo4hhJMmk1q/yeezqhtfIPS3
+30klBw5nUchAbwR+Awks5uxN1ndc5NiJRBVkjZTs5SKe3bG6b+B1ZfHxYR1i1Bq
xygqKO+r62+Qnk1BIyNKaxxXhs1MFKMi3Yjqj3nIS6wqPamlQGbMHlE7UfsrWeF2
CM9+f17ly2KFr72+VAgd6O7M11fgbVf5HFucxxI+fRZCNay655og5YUGzATeF+iB
JgafhXjZONCXSxQKltWJkKmq5AJdiDWPmrKIXKIXIHQpcP4f0cpGdYafUu0r13lY
/5gdChc6C/JBR9syamGqb8iuGWmg6Ynjztu4edP24fpkbBhI8QpZSpXnkF03Y6r3
9fIcYzIIJN9BdHhV+/ElJljjhZsHnksuHLe1HMQItnLroQGBkrK4IOxxRgYcgGGx
TwV+phXyeQ9p3zoDEXarmDlHfOsMX4hBcDT/WPIbX4RgYlNcwfYEPoYe7S3HpvPx
Nw/5wWcwIgF/n4z36t9UmOg7/8wxsdGziaCjmp7++x7qPgs7RqgNWJDXc7olmh6/
5X+HsbX29rOaRpr6551dnNsQPNqqJd1QCP40pGhjD/oKwAOyESRQObnBVMM6Uv7j
fSzeBRpzY2Z4NFPwnospoDJ40VqG6nPJO6O5ezSjI/W0jN8dmYuzAPH2ckXo1X4I
SyYmMTxbJkMxzAsL2aL5Y7CgjH9txsHYWo/0UdFPIWlgoaFAA9Hw2C6BLfMvE5c7
3/4jaEvsAUN1zbeDDuPcyCiKFCSTdvi7kMvEMkzCk69mB9bL7b19RujgtoCv1GYJ
4WqGO4fue/iIJbbQRoyrjzBkfOyolEVXuyLY0Vpz5OskfmukWif9bq7I2arpudNi
Dh3zGoh5yvNoP9Z8xDsueRhhDO9q/TN7kPFSKMMCMa/sW62/D/kbfS9nHj1T5L0M
Exp+WTtKR4Ko/EPcraEWlmsC9KzrNu150lhxN2jWT840mrnk5iLfnAJ1+5GMkQYI
LtLfwk0qcr9k1Ff5WE6bQZMhPB8jmx2oZDR2ZncNGfqvZm0ogS/gyN0edGR3p/3m
JbG/ZwQejGizqBgCsk7KLb1gastScjKuj2lB2lLuEKBCEHg4mXgC8wCh1M8FjgP1
4r6X3l4TEeOdAMffMfAMw51I373S6xVp00LlCx3eJCm/MGUkXz6N+W8yq/dSoUW6
YZocQsV++WFUuxS2OcsnCaugZ85JwkNqdzpoo7RIhhPwRFti/Up+rq1AEqOfEB8w
7WulH3HcBi/lMwotZv0alBh79vOpdhoBLI7P5PmPTDiQjkSp1bK48aE/1V5E3Nzk
FdKtzK39aignCgrklpXWybT6o537mBGD7+21WljxGL3BVvr+TfGEZTrTkE2AHGly
JHiNlgYGm+cMd8e1u84likKs9IclatwAS+3g2pI91wNqbWdPAuFjxieB1yg282MK
n4EEPMj59yRDy4tul3F7LKVrI+F45FKwk+xOCX5tUvYt5t/EzdNIaUbgQUAlMsKz
/vc833KRjnPNo8gfqB8O1ZS4Aactb4tt4YbDevKfhx6rFWTukOEjHl+E1dvhHTUl
3wwEWlk9Biz6qMv1AXdX01MYPKTJ5jar4Wtm70qWLGcr7+h7mOzUubU2LgKq52mX
GhBN7OZ+p3QVJJEF+br9pqmFLPFGu2b+DgUeuLag8XX4JPWRMFTI+vJNunOx8wTz
ywWZglfdMxNe74LaKJRL/VLw3Kc7QoV1M6i3Mb5TbX5Er4cYlQHw35FuPE6Nme9k
MoyiaKN+rsL5Z0ToWgQqTp9AgRSBKoPK6fNpvoXhssjwW4WQPk4iejNqgyySucm/
nKCwIFR0ry7k/XOG9NW6v2OzJwoKeebwUpf7yQH1MrXvbFohyvYMctVkfUnbMByU
GiF3IeLnFZHTd12GbDb4LSCUGT50FuZO5M8ija9a8HjonZlmLqbEP9fMOoSmyeEJ
+Mvd3MWsQdzC3GDjEQ1IKMrkIJx082+yzIyJsihOFfKBc7TQNlakKe/XhRfs9NmX
fd9Z39l9I0da9F1qw/hn6DOhRe6CToSS9ebhujr3UHA0i4yifeA1LOlHOaTMB+fq
C/PLd5T6bGjXcVFa//Btrt2pVQgBEYeclqdfsTS3FRV7+U10p33cs1tVMXg4RU+i
jigBzX9Vmu6KsbIlYV2UI51CrNWGpB9rcmNtcQQW1m+NUE+B7homh+Oa6JoP8yz5
wzdbZsz3anK1YJFI9hrFexsRjZFsS1QYR0j/RX6qEz0c47DLi9QFr+9WKuuwdeu+
0ReHqtBboc7BJASCtigR9TL8ocN3Z32iIABS0tGEVQiux04G1rt0qMKrIBMVG5ii
oFKKAg/S57UTi71mEHroc/EC+xigHCUczLOTsataEPqsijhRQ9t2TFWWOfHGn39m
2gOn4ixQEAfDE5wU8/ppCln9qYTorRHVojQSVdntAT3p3QtIyNlyquZ/YApvnths
xlT3wO6OmdTgAqy/7pGIN9oseaQK7/BPJXGa27qxqbC8cEBN7RdJ9LXMEVTU+5Pz
JRF+1EBWykxd4Q/LszaRTDdKGWPw2zsaztzSVQ/bsFSyncD7POGmSSLSLKNuJUag
IKN3EoqsRffgeLOw/2gGPV15L9dnfkY9aTkXCPvXW7jsdDxgxPYruIvUN/tHCIrJ
ZUN20mMM119ELoegZ/oW9qaQJ+GW6w9CwPQiKCMeZsdFGq1C0N8VXpLzPmM0Qq4t
LdgcRdi3hhnP4oF9sfqIqVOdqQIuT+WiAFM3x1kDaXlU6q/yDFy4VlTu85sfttGs
8vMZvIcTVj6FxkYXGKhX9QVqxafnZSCAeNlMZKcMNajTyH/7YccWrJuFiPTMjV0Y
kndhMKVc9Yedq3v46Lv6+/FK05x9uDxuCEpx3/TXTFORzAhT6GuasujBm+6/ddBz
lRKFtASFXyZybtO/z5usdFnywVvg1aw47vPdsflnGImCJ8VmCULcswckA58iQcPV
gn7aQ/k/4TDcBQiaR3ebnmT+5wbKPtkbQByGqdeDMwLmnnpiWdCAW37YEfeddyJ2
3BIqYzVIb85icNu9CGqc3IlLP+XLMr5moBIZ35vZ3v9sQWNaPghww76s+sNzfgSN
a8HJYvs39JfrzwY9Gw11kRWsQXyyLvaV6v6PkmM0ncsAhbMtA7rADkF+cMBfxNmn
lkqN6HvRat21OG7W5RYVhZz3xay4W+sQ8VbLdSFDmom6sj3DBDydSpQXgQLG4E1N
WjkFUl53psZOQrd5amgP5ToiMSF8wcNspV8Fe+u2MW4e006pY8v031ZZcpdMCyWw
qZKCT/MoUaIBYHXqYx4V2Acyyn/r7p+vtUjRB6NcT641IoYysnuf/tmhOh375oFL
lhUjPex7kj+yN6uqbiyRtanHZyaceoDsZvBxYQCw3ibSlaIwu8srIH6HdFjnpj/d
J2/Q6NwJhaowj+3D5IS297n1pUCxlV0txU6ZJAxsKIx7PVADJu7+Q1pnpEfP6TFp
FFGCkmWDnsx370ovq2P6T0S+WC5sQOZsIIOaiaP/E+pdbQC1C5kh3y5onxsHwELZ
3RQiezFT6PKv13EsSpIa/iVa4xPBEnOcNjYNeFR49SueyRrCWmDpEhCwOzpKiMRX
RC26JcSuLY+pcF7KzNwutfRo98qMvropWsLLnAm89YkW0JlJ1a4j0oHd1rkl1fxK
cm6MvqigNaYcAjccoE2T2TlzEj1NF5uYQGRN6/zqE0w5ikTEKl/RmH20abr56MQj
6WtrmTP53UaMC7o601wpASFJGg0ZI1j4gVqt0vp+K47Z1IoOfnI88uwK+nHjBiMr
Oqe+1Y5/DHloLXkvKXySuTFjLHFISzATkCSB2E1lv4mnPqURLWUc4Wc57JCGP0td
0yeJKGikaKct88tJjmzUujZrPwAVUZVWQwXWaxnyNDXKg9ICCyBtgnx1YRDWGWYW
x4g5iQiqXrN8AbnD+uMHCfwOUmUhzzBm73XZeOAJvO2juLR/PdMnoA01jj/IVQEM
oYb+MntAR4oK3cl7UdU9zHlKgM5lcb5BzBnbJafWNYAkNtkuJDektW+5Y4QVLd4r
XN0dUQOcLZ1g4lT8Yb/mbs0pRrQeSGZtARM6wTD3srS3nzyyTQav+VACwVlRgR/y
oO7L2DUn2ReaK1HY8cdsV+DEmLTOicZRYDpWkW07nzw2a6rIMIsgrX9DxnKVeIlG
IN1sKt5YxjV/kRBIUFWmfoBvAkeKEHeff4Db1PSN/SJbajcGNPZKINN7m+56BXce
dn1xJWIff9dZqCDLuKKcMNqIF5sUgTfWU1trIMnbJ5f1aKDoDsNjqr1Z6AiIsREm
OEX7apVA3Sx4Im/Datn7wCGAMqdiP/rvPGYt70gxlW7BxjYMD563Z3J7bMxU+B4C
aDfFrwCXEYjhojl1P+7qEin7tDeWx5zzPzNGTjDB3Vmp7ml9aOPFKnrEQLHiLo6z
g0mCHTThLw96NmJAcCOpjC3QynndJVIctQqTKd9hDl5nq6nsVI4wZlddp2Vr5vKQ
4Lb421TLFj4cEcrBy6+1XCQuzWJteYmfc0mOr27e9CVRSBdZFpqB9A4GXju4TE9D
d0KwXB/j0arrVG5e4COvppAUmVc3lTrnVEvO1DjeVwL9QqQ/kF7/vvhG5LhMbx7m
fNnNfd9EM7VrrqWaFAXUwx9rxCAqU4wJ5E8CTvUa/T5ZVJgFTjEnJ/vUdozqjaa5
VQKkuCeETlrVoeU7maKmjSizZZ2BfNwyBqYIUqgMOaRmNd3VyOLQqrXYQIxuoEYV
rH802XxorS35BdO6IrePvEqbdZXGemgLqcCH5HBgMzYEX5OyhKT3WKJk+JWbUdqy
Wbv15kT5nXcXWCzJ+tNd63ViSLtTcNRwk9tj2EnXe/wSA6ucW6PR4+ujr4+sz4hF
6QXcrpXKRICEMnkjq263aHDQ4c6Fi9bzMPoTbAPt6xaCZI5/dFMchVMo7ADoDU+e
i+k6QITkyxFrTfBhDK1ZgYpzooQFIMO6EGitrgpBZPNtl1E/rhYv+mZ6tb8V6ALy
J0pKCJwezrL+HQy9WRnCDGiszd9oZV/6zUansKgLiUfXgYh3QSf+g949cKr+KMJe
8KAVS6EkLcSALOLhtoeN4QpwG7119zOfPDFEP5WL6FZRJmNws0deaQf0tS+UhiJL
7di0OafneYy5PiVJC2Y0eECJ/hIFFw5aJNzPvnsKKuykD0cWb5LbdvrmV09QOdqk
xDP7mkvIAfS264fHG8uhR+L3HbSWAZ8UEptRRlpw+h3VVKlhZ6yVqNZAlU79mWQQ
ClvhNMu0GyRCqNTuJM0Eq4z1jmjVTmKJ262t7o3mqzPEVr7snpPRfxRR34IFVJjl
Gn5srW7gXZ9sWes2hm0TLtH0w9E7WwKb/aSjpVN5U1g2DovI7ajL8EHwM9X194fQ
9yFD+MehaZZJfe35XmWbrv9BThYjMJOyRMlm6zeKzNzB5xiHWrmhv/RKCo7kC/dF
HP2QPnPdkcnEbjAl1V1fV6gMK3vUOB2YicSW3quh0caBO2keZu/LE2fXB5yTRU3w
r53FAl6WHAYP10YtZmyUHpDi372mDA6X+CdBgsZ63mdfM8S04xAaIJj8hircDRTU
wx+gC4I1cB1vmndVBdTdssXa4GdZ42A3MnC01SO28/mPzht+9CWW/R19keA0WKRj
UPD1avtTVm29Q+EwV9jUy+sfeKw9M3ZSpv/yhs4+JBs6ecCNlhSq/u/ImVfj/M0A
V1Z8xRSJqSJh1IG3vt77ZdZBsbrDkAedQroliddQTd+zj6mg9hITsI40ZW3BN0Rx
n+SpmZtCYrZZ+6sIo2s+H0Dpxo7NcJ+Rt20yZsAIMmiTLqldb9ryled+gre6uxFt
HiGDId3WOQVCEW+d7/mAuTwF3cbP79ErWXwx/Ftb9FPZL9AqrTWqvOc9CBwqa00x
OsrAIW/G0qcGWAcmMfRHyaFaWaPsy4lscdPLQtXrW+zzfgu6ek1OuVa07clbXkws
PbtJ+aPbUgDsBwcOR1E7NgS4CnDZntNDRW55+07FomrDoEC0C/RJ8v1LCEs64Auw
7RV5blAGouMVgAUhPasZArJfug09xyzNeUXnYmStM/Dm0fzv7TijzrAgNuUS3XoJ
tkzaYtZRRlWqAVn8P+sqI8Q+efbtqThum4aojXmpwPyuGL5QEKxeb56HMwRMPbcs
R0asfkBOkNCdV+WIur/WjbmBcdw/Au+YST9WKxlclvBnmesIwSG+gZddMOKCsgIt
gEIRsgBv+n+xdSY8WWj3sMGxw20UVk3JXuqy8CpIetjydbAh/eHpGHmc4M+t/gNr
xiwPqU6n478lp8d/sLVbcLkSOupSZLNjkNJJWS7nwcgKxQR6+jdqjZFk60xQULWA
GyOD0kh0rZhPzl0Z4zNDel3LXcLXeVCU+O8dLZMLzRuZLQFz+sqZEwHYg2iGgXHG
OpmrLbUbm78uTx8VBK6JxlbhGmrYrOoYcaNo81PCLFp+i/96D0lQHXlty8UOCwdT
htoZm5caDZ6XVQfJRt0mONQpRytBSts1jyBhUxuey27KuWRCYLmJ1TLtz3vDWEaP
rpSdYpqWIpxYJ5QXoKHy04l4tZvWGZXN3qjC1g2IVXLonmpZQgdVh4m3CwTDgUdS
yNLKJmhY5+XMuotoDiR6sKyf17K6/YIebhUUpIUU2XdmB/0SlMG1FzBtxXQvVCYE
6myAoeYdJ3BI6MyxL+S4H2e7VTrhLzAHsySbmCsJ08Enjf1IbSUWh69EVC6BsHMi
oKQWVISOG1wL6FZEVBNoe5PAD2XQgKuSGQVzQ9TyUxGVlBWl2GHeT9PMg+qa2uV6
bOCyqRpSuvE45caCeXCD5OxbVaSIWkGZfLeBYwUH23G5p+9F0TC/TuO3yMUzcqoE
qT9gvWAjd3GwXmPuuxbt51/RPS2TopmtMqcHDhK1sCJbg3NmVT6D6397LgcbNU1Q
+32XbHNioCXCTVNA36z6cSyyi/AH6q0p2s0TuJEnDKsaKfwCXK/kkQdqA4J9ehYd
mDpEGLIKCTdnbceVrGpjqO7xlX2w+LzCFprr74OsKrWl/+lor3ym+TRWeg5OFBri
jzYKGWX9rXJ9amVmRJ67z4+Bw8sJxKRUIq2XxEH1eXJ9E9Upq+ZuVxvRnsgBIfJ0
Jm8hNtziJBWwd8gtqI1a48r21fmtKAir+XtZpIzU7y3+EfrV4jOtAEgv4THQPfER
OG1jpFrKqdZ6yFs3nRXGCCD+94v/gg28aGH0m4m5CpN+el6QkotvUiNcfYsQatrE
HVl+taqNzx2t5a1FrYE05sLmPfQbOvMMNtuWNp2pDd5L0OzdpMNYByDqp9xPpf4X
sC2+mK434Z8mL0RtJnpgTr2a62V6rw7eu5iRlofEuPsIyA8XsWmESEXVvlljgxGI
YjZaKqDDANCi2zKFjhq9VCBBpoxUzypSvI1X+W0Yzxww350JeCJEMf4sCm+QIY4a
iK3M2tiTksZrzzxkyojW15rnDaum1RjTn6cVOkf9tkzs7fvL5dWBe3QzeWGlnR/Q
xwSC5SqaaNTnhLudRva5vPl9GSC6dZVpMEcVdPk3GlHwcURgVVpIzqfIEUuY/kMQ
ZYseBBRo15B/T+Mxka/yyS+6fd6Quuga3+DBPdWgzpVhuvyzZRqShA1SjTUaDRQq
W5semuUY3Iq6q40tKq78Qj9LHTMo4WYGeYMswDho6yswHlbI92AwxCrQmS7Qhq2t
cEQYo/+UHF3zviSyQIuCbV3kovwGWRyt32kK3BT8HG/bHkkHvxuMRxjRPGPAyB/S
LfL8Zd0CVkv885afMzIVGavId4mCghr6op8vh17Bt1XTEmHQt1DrnPuyYCCPtyxT
A8gaXvGeIuuyMAUJAvvhlIHdniBgv4/jOwABJbV6s0EkCC9w2LQ/tq7t0+yssHmb
T65C1pa7rVdZD/f1quqstR6nuw5/FJWEunZE7MQgvwsRTYleJ+p15K2IQMiVGRaR
bX+nIgsSAG79i5kAc/G2jv14XEdh4nITdRKiTB9JbJQUvrO+MiYM4+cRUEBnimaP
bXH8aL+SRw0sCARgw3QJtLH8H8zXzXAd2AIcgMh7XvZCczFXVM8jCAvs8B1UcDRL
TKceNCvvujhvKPLXE//suFhkA6bJLpLb8VPPxO5BB9QG/8TBSCV9F9+pEMB07RGt
1xjkcFeHIjL2t1Yot1AkGMiTh2MreMvGMaplLpBRxhwoTUuoo0K9SFqWsz3s36oa
Nw76kIQrmXGN7dh7HuZ95gTHUuJmXPxZOuTQ+0Hmyz3ZDz0XaSZ4NeWbrvPPw1Qe
J4NlYULp7nuHiQ+R8ND/5QG755s12tX7IaeT/y5JjttRPa2s58qCokyPiM19WXUS
CdPw1V+ODNGXMMxjlUKYI9svVbhhvq18b0ceeJ5HyCTsWyUazVl92piiWdx5tk0b
Iv7alBQ5olUc+LmCYZGcOzegCsdIa1wcxvxeDZ6YJYRnV+3NF9Ydr5tMKov5LPEF
2bPLczo0GZG3HAec0SorOzhAjvpnsKPk0KLUTAECSz2OXDPcHSNtixuKSTGWnT5L
ruZGQqTE1C7nwIvnpOwkrfv9fSbqPPOpSIyCOt1eaQ9SVFakw60v+cbyh7v9G8in
YueJCloj451H6EiYLgFFSrdhy5Pv76Qw2QaelRFnmNhxrOlVgrvNwLc9dePsSu86
8ry3aR7LebkxVHdf8lP37DRYy6ZjTH3tsbwaLTYyb3uKpJp26rqi8mnqU+Pb5lTs
rIGCqRtJWUWKyLivNv1oYwnGGncI4S589R2Xf2Tz8WzXVpCOY0PnSgLoJ6XjfZy4
Fduk2SqJMgjLlmaGS8FDjoFw809qzvZmbYt5g18oUVHTNXcfNRRhnvtkBrqbTf7g
juUax3HBKrs6GmyehcJdqAL0MgAzJsk7oCpTZt9Z/wPoAo2EvQEP+/Q3Ant4OYqN
RGEH+PROZH3OmJ/HO2DxElH1v59/enq1O+oDW6Szle60VrLywYCoq+N7B6ulg5Va
No6dBEkMiVnsO7BfhE7skSdjCrVZjYWTSe+W0XhG6gA3aACVaq+8W0AI60h1jRP8
sg+PBc3o9CfjQG8RGoT/5EfglicxxHq1BH4RSL9GDdkHIU9vNFUfYlUl977bWBMV
Z7f34nTiv+4APNm2zh8fXhk0dS+Z4kM5mHNr/NAs+diutuGdi0pVtEj1BA9vW9mb
JeiQnoVk7x2oOTiM2eLQRK7CBT2vgqRbFX7/mrDeFhb0f0aeF2WRuUXlfLMxt0rG
kImgQCCXR6/VzjofPmhrrlRgspEAPgWnKtBFe4Ji03z6Ed7J5tuMgj+o0zBAEsZh
VjH+pWInuUwDUd24HCGx0UPvYG7hZycOk5CC5v57vUNVLw//SbPJ494ABopoQD3h
RRgflrrBboSZWC4yBgQkUrD17JQAjHrWv/wRtO/of+SEIBAo4Vbgogw/gh5Ujk6C
goW6Kzq7VUNE9S00UnMsqiQAC7CmgDH6sC5rwjQipWbAP7iL4iNZAeiIeVmlxFc3
DMcG1Lgugck4PrfLImchoIU8HPKC602wi1c0RicFVuUehEwS8ciaCbqFcYcBD8vm
CV+y4ySaa8vHm4+bB3hkY9cYxIG8oEq5Ly8QjAz88tCbbi8lWqS9dP2eSrvJSthS
VeoC3GBu2qIZ9YYH7MN7BH6kDHOlLhQFIayOo5E8aGHOtob1z3sqb5pMcT5VC83u
jrcDkzo9NkIIbvy0uERHkPGsZINcMYKcq0GH0l0H9jB2dp6uid1Fh6bNvoHTcq7B
lVFCO/kdYllUm2RjW29nv5XoIdDAIPfnf3eE0NrikzpC6RZXjaBf++HJoL067+vx
noLO60BwK9ysTXSPWLMU06oUvRiID6Y9LVy8wss66vjy4j2DZP1Ro/qK0CJdfqG4
E8DUPjmEDv6VrHTv4qAKegD2zSdpJs+xZk/Ryv90KfJ1qK1NDwrB2jrjY9bcOY57
bSletdA0jKsufUC9DEuBItbS94zqwISnd5+T67oyV+j0JZykmAvDaO39qUcSVCpZ
WaJLkce/GHe61wtIhftDfwmBGS6N2G1nCLISxmvVtTFZgBwa+edOmX9olfexlm0d
R9G/Ri1Z9lBxkCUaAbsktiQe9rW0K+52L80Wj8rAwtc3vUv5fpWcJtjb9udPvC0p
HadoLOxcSBhG43ETzg20tNphD8U8qL/ZQTTCspeZDwg+EjRpj0TLg7C/xjZe7Gy/
iyxAuLq36p2Os9mefmwYKT/d6Vr1mzlcu3nc2kw8pFcjcNCQI2fK6ASJ7OIKwpOM
AdUa6Cr5shvb4q69B8caANnIonbRoWlqGWT6+7hMqVVWOx/EOwhU42KpkKgVy1Z6
Q3VjdKMsgD+Hn9oswNT3WmYxdGYf1dWZeH+2xP0JsHlImD9BGvJWOBg6HqOkv/0P
1KZ8DJewTr6exDVscTdSJjVcu9QUAjT7QavQQsNAwZDlxbk94u2wL0UdO9PeaD9/
Z0I8IdAkYBLKp3r22Tlvx7rUTNYZWEEsM5XQGL5R8cm6CrQeI51YOHn/oYkCIgRk
PSnnhGHIh5bPygqsffp0BnbI1x094OJp68SX5HIMPGLfyt4A1WrmrlGtkOH761rn
b3y2ggRseInZJsn+8/L0eNRn03LKV+c/XauozjJjfcwc0+qmbIXN1+c6B88Tli5U
Rbk8J5CbO4lj0ZfsTTWWjd0X2j8w/5lc9e7wOUOmr2T4Rz+X5wCPQEQ53wDQpI+j
0r4mOoqZdBKn9svbP2Z2S5Iv8L2xX5QOudmaxQtK2o+MFX+63qYEHfuNCgm90Y+a
tBofBKxu44recKdOtX5IXaPjZDcRugLPog1orEZhdudol2yWJ9y2BRK3VSjJ/zdj
PQ+ePR/TicgRHH8P2ND22kDhZmEZbZzIXRCRmr0zfjNUNSe0/bgiEDQ/6IQonVdJ
kjJ33JS0osYtBQdwQOVb2A9VxjcV3+15LMXC3H9kqAMmq060TCJcRVrts/OO5ifu
GNjC2dDGOIygp8pJ17z1CWl7LghB/lt0sHBAlnImRZEexaOpphDH1fUJ3itiEHyQ
pR9ExeKmB4eSCSpbl6H5W0xmxxHZSxS+hyTI/Al0uXidmDqobS5HoI6L3ch+qESx
b9owvQ5Lja6zrPACsJ20vipIpwgYuIFBvB2xofq1UzKerte50MicfRAQXFCh+/B4
M6kUDWWCI7lz8P2B5FGNbv4gE2IjDHurnlkEMDhfxGs/TWcCWqac0iV5x2h6w0uT
Re8rrJTaBeeDpDPEvrQcjVv/IlctSX15u4Cboc3GNVnAQseJcqPZ4chbcJlH2Fm7
VCOSfChvItvxI4ZDs/a/b3Km34/YRpmgCURonrD6kGwMriEHqeYely28qHKMCgHR
IKmxQyxoWnL1iisuOyaqLO5+TsNbYJx8weaHixdvYERV+4iSs26u6RMnU3wxNwcb
q6fa4NzgX+/oGcncxp0scGA6JGWA2PDY5Ve4f/Ae78ubbC9l6A41yZmuG9fWJqdX
8JBvfGrz2ZxRUyxIN7xsuz9X4JgtA4GdjXP6KAhqt0Fi7NYRozWiMlEceKcDrSEC
wTnIqVGDlNvOy6ysnS0r2G3w5N9ZXIxnsKM0cP7ghdsDV1Xqc1tnMFHgQEN3Rq5W
XyFC1y74q7dnRvDqU/glfh8kqDKBtX2yMQERtLNx6CyedXzhpW8QZlM8tYDwHmU8
av+LftE6P/FpKjXN3w7bpnl4ZsDY4px/ke0cnnyD1gaZCaXBpUV47odIaAjWjE9/
PJggNdQcArE3qW4BhLL+2co35wIUISOLg6iCLO5hK3ab7o46XQvU+LkO/FKFye14
Mz3W5kmO+XhT0hiSiASAdilQkG8WyHQRWKCk8pjSnRYEMuysZPVzA6/oj5zg+Zjt
2vLKDMmbuRIrcjtF8317+wOp/sfP2COEoC4pJRHOsMAQnbJUjkE6oZyPsosQRTFv
G3/apZKYES6Xu23MhbNBMugBOBujSokQDN8KFT4A7dZi2XhHNwoxtYYLK23DO6Vb
l4XByu36JIDZVp2QdeScTazdRKX2RI/YzYZzVCvxK54kfKP2AC+J9D6apnmHYCXu
kZGHWg3n2ERIMBpBTDP0dZYXh9425YiG9NBfBfa9kNifDqQKixGzxu2uqkaXfknd
QY3mbEV5OMD3YNm6DyL/0hwhUwiTx5MB8pNsPnxUmzZPKx07cyeZF/K/K1B1203m
Yw76VKitFlErIXl6nq+0r4S8RQx630zuabN1ho36gAuIaEy1pEsm1ajnll0ajgnO
lwgyPwPggIj8A0r1QuTCI0tJu8NVqB5R8iYaSr2jzheR20aQ5NnPYNdltnW4rH0g
95UvYdt2w93wwE6gd0YzwGYprGCiDSLMFeMrnpqFTRPFliBcWLTCNvHZP3Ornq+d
mNzhrrzkl/BAUmtYQtYiEXkSRG6z+qRBpYh+kwoVAJIoEcp6NDpswr8uk4Y7KFsd
jjxE3yHiygwTcA2KJmhsI3jJbJhsYhGvyiwTPrBEXC7Zc0KvL6m/Sd8Qj/WZFrf1
NSiVv1NdB2eS281PgOtYA3/IQi48tXLx886Qfun79Y5QPFlbv+tNSCEAStVN5g+r
rVXJDu58ifqsSl4kOA5cQ0qaf+WLw2GWx+Jk83q7hH2x73BdyvBiuF98EkiP4zcO
EpRh2qXDZgrQVOpYs/CPGM314N2pmdyNXLaAio4Ne87qR7bn7pas65Uj2bH+LKYc
555N5IPtIQXTKIWl1Qu0IAq5UOGhPSGCoeCG9r54qg6D+4L8BLIS6I9KmGCt6OUT
twDZrENdxVX5FKoct1poR5OMDZPmBbovvli/EFULA41YXisDcojLe2uCRHwFY7bH
T0+d702NLLhKaDMFvzTEtWseh6lz5MVehJxI9F+GFG7fFtQ9KTsZ0a5eufzPHmDQ
84KTJ5Ce1BZ4qY8HbLgbV7ny08DMTuwUHOYee5EaEaCJlzhVsKpo+ybWaX5opvHM
FX2rz6cbLW7cX7T80a4K9ZyEDfllNKsx3DhpzTdswJJlBkqPxknhyxKYkF8T0AF6
7CYIULSSgnJtq0bRXFXxKWYPzo4LXsRVOIcsUPHrx09xm0l6GX1aVPsJw339o2l8
ZsYZaKRym7BgjRDwqGvepVMXsUnPshH7bZRurbOtsPd87Jv57JWshH3z2yoRZG6B
inv3+xDefeTvgYFjsZ1mpIYUItUuc5NNV1Ie9xsqM9XdRurc2YZ+u2tszCLPgh+O
dDgZWJnBFaD54D9B1vKQSwfR73s6oVIt3Ggf+LQej7xuJJGsW5ZCq6UIdAhIH4CP
MtNSSgZVxhtAQ/WbNiHLOb5kzP8otrh5RDL7WDJHyze7RPF8fDuQsEsz+fekPE2k
h0ZPYuB9Vu8bM/+vp18OYKh5rQ0jK/NrK/roycnOZQzrcXzBDPUA86QmZg17WH58
dHgAMJftnTXLGVCwX0fOywy8IrR5G7SjBMFNCD1bWyO6xfTdGR+fG6AjJG4TgwhV
JWAI8tU6r8pPpOS22dKe0i4PJOLPA0EREebDb5WisFgivxdfvPbsiFZwcJkaYmJy
IhxfYpNWhrExHxTTViGFKe96XknkeDvSZDGeHPTRRe+gg7Vxpbdg9rwd3v1JRxos
8f/yHJpqsZmYwvov2qrk3qVSv+7E021m7dlr2lRugM1PY9j1VF2WZsn5aGSk7jY5
sr/IHjoqMBlm/77016in0q/BGgFhbvBh2+kGEw8JFVc78O8f3YCobH5NWe4w+ZLl
yztef6AeuY8B6rYVYZfCNRY6qKcEz3d+TDmxRnFXwKtiChRAIQhZlrFyw6ZNF7Sz
0xsSRRwCb/OybZPmQ+/MJ5U/s/+pxsGtQK+9RjmicG0CRTt2L8QWYHxhJYJdBl19
vezCGmaEdPmSb5sR2/xYp5f9sjF5Pb55rcdJ67fYBdgcoNJsiUmaQ8TFQYABhGFn
UIQ9VwvPQgiwz/MqDpFo9Rr2VP/NAMfqhQgY/rDV+MKGrd1HVEbZOHDFa6Mym7+X
1bVunsl0YtZC2UGgnoHrJf+CPsNbjXEYxyRmXc1j0L9DD36GfMJKJnvztK0MqHXi
ZYDl7fhSqxTs4CfC4kmPHCDv8F1cJnmRuBSkvKFcdquJBHmI1RQfqOs5JTkjpL2b
fHWWe5Sqo4uqRuwsEedvcmFeQs5g0Kof4KPTqQHHLEeDWnDVE/0WbN1qd7oMgA2Y
Yd1MhmSx8TE1DFxHit69zImNpOYkhT9ONNJH/Kfg8N2KY3OvcwAo7MwIEu/1DhXI
QAWlv+O1+zFHCDyZ3sXO3WOEO0Qs/xrkI41RaCEXpijzVNrX7V/It6p+I+WeFIVS
IQ+z/KxIZtRXkXdx467pZdx5oO93t8/areIBxzDQEtZlC2txzPMb7y+wlMLFpg0W
pSbnrpWldA/ovvyeeuRZ+cYVxmdntwhuwy8wC1CdO3aBzM82+UQwNR9V5cFicLu+
h47nV0iPm7Wrs8PTef8jZOi5+1MmjVc1oGNCtLSQ1GMYjUbeo4K3Jx2K8UFQcyoj
05wDu1CPVpQCT9VRqM5dGgZl4ijHIOewIib8mUxduunmVy0WSslvLXxRHXb49dco
el9l2E45RHDQYP0nT4rRNFLtourFgz/OLiuJeRV7dDpjRj1va1jUMjJVbYMqVVji
NI8f0j7Wz44pIUzDP2yU9LJOR+ecC+wXrrmhxoJ+YM5pzYU/EfC4M8j77DtYkGsM
tqtetef0hcDIGXVwUoPiprS7hPG12o52pHV+jhBRnHlI9weDoyjys7drB+I4DvOP
Q8c7XRFQ5/YmioMRh8rrRw9qPasAG0N9DRFgk0DQVW6Aa4qcrhdOH3FwhIE0ARpM
GS+NNjK2WJEHXJZU7pUjkVWduIOU7WV3hpLcywSyPCqr2ONG9YIxtjWGWEyaiidP
z3cM41Oke95mxLCKD2zOvwMR4WxgVcALGI+7xOFJD/NCZJpUJu7jRXiLyaBQflJr
TaP6WqXJwHcIjs2O6CHEcjFFa3m4n4hVfThrTybWplLtk0qm2fpB5gaH3ffKOByD
rnC8EuIUzJfdPWJF7zNdrkv6UcVXIg+XFMF3ApIh+ZNfSNS6T20RfQtjQvkc5ll2
DQ+zN3epf5Y8yp2exO1K/XD8hHE9nalk7a8pbz4BSmDj3oWxWpKK/1BWJelynfrl
Dmkj6duy9nd3pk341GCuZ2cyUBpWy2KtELOe2DNbZKYBAZBoxtmo9WF7CxCR9bOH
371nTB3/renD8pt8NsfUtnDY1o9BwvCxTFYAMH3P9pPwn+k4ash02OcgirRrQv4h
217DCX9mGgan9wfupH+nPjHKgknp3yX5gmJG7/NUhVsR0GSAgnRh8PUWTb9cS7Vo
F2OBR45/M/bdiW2Kyw8q/2PYvkmWLpRkcNDZGs0cAhjUCRCI06FuNXnyU5a7kFYo
JXv3aVmZivqbwE+XcA7V1giLGrDHJyLL4wCL8FOZCtWLnR6O8DjUZWxuxJ8dHeQF
Vo3rD5cx/AuRJJmPHlWo2LhSHXNoBY1TbLCvngzIozSibfg2UWXX37JYHEGLTftd
Ez/7BFE42rtaNtFmFfSvm9YeuMI7u3keuLkGa7NwGB0RMZCqmg0AGp7LdWSQ3Kqy
blDFrAv/YAwDFuX4sHHj8/SecekIe9t88lVZjG54YyIrCBirY5pwmEQqEGWR6DGH
12s+GxehY/fYfN7cwyzeD89wy+jal2cwWHdwS0aVNeCeq4aUIwUf/r/1UQt9vAK4
D9xw5lS+K4oRDkVv5QqMvaStM04Z4pKiRRITDw/XhHYjJDwlvL6eqoagDYkXCRh7
3qg+PDAViB/guIApydYBm+wVJ6sZ7jE4HumY0HrrZlO36OP76xVDTi5296PYHmpB
iZ2GAZpZrLRRVRLMrW2QNCFi65vwIHQs+Xhj4aSs6n8MiuY4xog5nYpWJBkeUMwb
oaJ00X8Gc7iHKAKuiPjV49C/GRPNrH5qrREanTvjRQLY1NjZY7xNLN9Vama+WKmt
cX+UOLSZQp+n8wcSuZl25w3mvB7Xq8Gyqs4CTwD5ysj51BzeubihZdtsLqR38nrI
xyF3v8GNmu+ZKgsrVq1C7iXefiW/LhTuvGujLLF7Q01bVBZwTAuxJAK8liIUc+Zz
wYSdnZK/8ZjhkSgRDPxdXlniqzg/5zxDQ5zgKLn6ohW8SldmbdoPA+Bu6Tr5n66b
u4GSfl33iKdgPjZ/98Zpr9WGzv0w+WYkIwkSv1FHSMsp/y7/v6r+7HcjdsPuVwSu
DLo7Yy1iQWdi0ul0s2M9RZ5/zDV9FjF8tUdPAX9wDMXvirHmwI/Opa2MXoayubee
hgdb7/0DhwVo0xOJvZwbHs4oiwYNCwIk/l7D+4mozWEhlhhAoIFe5nPtO2a9vVGW
q3TgFecyp0Jh6rpCFDlesMoRLubFjo0ZrIJW5jRZpg8OAb1p60FLKdCVArLsQFWT
FniwCcgJO2v+5pj7n4EEjI/8JTHiqYgDyHJzhZ3ytUzHxbVxe/XA7gpBHsaPXql2
94HiAehVzLLXkHA/0iKjwyKkQasH6rjHVZOxSdzN9XmcIAh5Wxdz+x2Jd+PELase
VWW09ILHV2SVspbu3kntL+ltByMwkl/byqXpPEN1yOODLyHAMuzBsNaysvuuSpz/
84LrPcF6PmP1Wzus3Gj0inqE44fFWNofC50VJxHFyu/jiW+eZ/HHsE+prFSFmWZv
4WHGg8dG5Z6meHNlQzLxLLLY8SgiuLzWkwOpCE88+8NnV23ICA/SPxi+5rrMQ1OC
dr0Nc32lzVFoNZR1hz1WwoY2wHzvF8byNghy/+3IOZHzC3y7yDvSPXcbar0z5HSw
UNc/DixH55LTkUvIUpheMM2+qY+OqqKngL4L0BHOiFrRiQm75v0UkjLq+8104Ugy
imWMkJ9ohs5nDU341cKjDFW8xIpBLW5yA7hmfKCz92hz8CD6xxTduu9fzmvMMM/W
5H/iOFoDq6wNuAzDZ6J4g3vcTO+tlB/SZAAKHP5L+32YtgsNPEo+bH6yPjly8Rc6
nxvZn1N/NMcuIGd4oGMwv6qgk5F34E8VJ4dh97TFKXIJt46WznOJH3a7n9qt/sQ/
0zY7UjQrvsbXl85QR2bAbVZGtwVmSFdJysZluR0YmgYzz2DcRd7AodjLfuhTpcoE
gMLDoSricRW0qFkcq0q81zp/EajZL/Fj6QLWh3g0sXv11LBhc5cM/nyWi9StTj5h
1NcM6uT0Rr1rzMYfoOjF5CnRhq6iBSVPB9bnAseeVUd/e7jg391+bKxCCO2mbv1F
b+/d1RMcGKAQMpvQWWAdsB7e8bfYTazcceYUDPK+W2LfOtbo7t5KHRFfiDyzfLU3
PfBjaX2G+D4AAErj5OirnUVh79DejyutCYvS6/KafgtWinx3jnnJu8gssvpnLlcM
kSE/3pjjOoSfVKhTyXL6co6bvE/KmYRRDn4Mzg3z9xgJVbx8WJsYF+/stpRdGbvR
OKNZF8R/uLn5ujFgoKRFI0vv6c5rCgM0dQXetYOoWo00DwW/ux7kpbArfRVHPbzf
7Mm9ngxwX9Bhi1X8m98SvHLuMjs8YljVO942ICCRlwIPSRUCStz92uDWqo2WevyU
y2OEeCUG/4WaEL8/adukdm6SfCSVDb0Ogw14FqtMeq3aX0WGxBIqYw+H/IGrFbXL
CVhjB/87DtgV7XyVZ57mBb9f6034pje5CfZwRah/LQEEvOoXQvwdMgs+4V7FqcxO
lQNKaHwXnoAOvMjBrTmEVqWYVHjtwX7s2C/TV5CHnyw2NYbiWkyurNi/wiRiVfOR
e5DO4rBY1RxgP9vg2C4tHF8KcMJJPzOBFbf4Wq1fdETFdycd/jD4dhsTcYcDRfwh
bgC69FN8WOi3Z+Y+yQQfUdg6+/9DiR1Vo53xJ2rEtfn6xHNkxfQSZNA2aSIqya5B
Gz6U+nXJ/Z1JC5cxxMqvCTo5PR4stzZD1OhAhJrhCEG1/UV6WF+zcDTobi/04KUc
FwnwzrUl8JC4u8MucEBeJXRvh9A8mFCzNxr3aQ+8TFb6uGVqHLvBFun5H/Y+JDSm
5GNuyNfHuB7a9OsSsar7zIWGOncn8hBSHEQFNBBIvxpaArcL8mpHVapvUQJaWm6b
MqfXSwkJxwQSn+P67NAqAgiPJUCnxmz5LX1p0NfwxDfSxp+Qf+n0ZAO9xZ/SuBkV
35LXRfRLBQHKqxOWeLeaiZvjCFR6xN8I0yxIfoBowGWOjseNHcS/8WphSk75mI5j
uKnUL9z15VEgaUkcJ8Wr9Bh7Y9cRR8fqET2mwpFUN/MpNn0MVUCsYTNmKvig859i
CJtEe+Vk80R1J5lB1ayQFalBnx4dvNY1bXYouCi5AKiDWGCTQyj2EJzcnUvTqQcq
xKwud7Y0o1yh8diu841zy1DYtmjgel499PKgKRcPbiAG6HwYh6cJn1dRRQYbK0XE
Bse1DPAhyX2mcbPIvq0hN9NUzglL43s3FYUd55nmrKQAak4RXMnsKqYBDmbez3qP
CZDA68isGNFbq/yuM5U8uHpMYwmdiHmwO4bQ2a0u4imRnTQYpflusqAro4OmGLd5
0sijrwq2yHs7zxDvH2/oYUeGoBcJ91HtxuWPrfD9yDKVJVgjlGSt/iH2+nEZpmh5
IL70NrTWO9NeUj1xf5jjE/N/Bdy0fdtoXTfRFSHrwFQMwm/A+SPRj/vGlmaKfKnu
PMRBlctDBfX/iKHxW0wIHXB8WxcEXxEZNAzqK/78/La99Hgg6XuVSfLh/fJYNsTj
vSF1ht1NpN+oLQSLTpzrcrWULY5SsDNoQ13UYoo96jisNtcINtYZ480M/cRnghxr
LFNbzYKduQLhIOAzt0ZmFSUuVFJnJuz1BN8aO5ASc22KvmdoYeYnEcz7mxGgRTQD
E4MBL9hS8PX0xuDG/IbmhT2FRHdqbt2RyDJ2d+jHZofps2ev6teLTlNaq8XGDnoC
eawtcyOamAK+XJDYd1OPMeXsj2uV7dDNPArj+Nb1Vc8zUGJG6biBqRGxS+KNvd1g
l46lEnJOAJOY0OUUX8A1p/BME8sv3lBMnSITU1Bm48FBJ0Y7qNX+FslJJE/aBmJM
P2NFpJQGwy5NWTXaCcls5KDi7EEHR5Io1yakY7gReYNzdZR7kavAmT0HxkMGE72W
v9C5/XROFV3opCcZ9jD8+/YwOOGNzYqya4iSUk31SKFUeCcLkNzJUvgW/DAIQqLq
8fPjsYYtgybQELakjmJr8EoOs3gNCRdTJJxyjhioP6YH/GpcdyKsX0UMcjVVw5cD
4mcvplP/fWhla9p7ckFteWM41tbzg2UfiC1oRXL5hOF5Hg6fOoG/6V0B/d1EQYJd
MYii+NE0eW5v2VDTG3YRLABQ/Il4aOi/SKKIf0wPMQ+AQ5LR10KvgeA8dNMgU1+6
kPQ0nB8sqXn1csoG3qxqGgCr9UZmi2+/Gxav1U2IdmQ/oQ/whZ5zoHZuFsuHKsay
p8Geh/2+XgjWathq/x+xxu3l6qHl8E5uuXf8eEqAjY5/hE2gSESr6eeo1NAuUicR
lul32u/GcTf1MUsxKsRAFnVSHhYC0xb0k/w0721U03NFeNYdJXOk2FENsNY8jhz6
J6ZnUSW2J3wsQ2XkpX6SGJenGH7E+2hX+K+8pILUMq64FUX+r7/GNJSzvCrFECkK
5SSoBizkRxrQ34SK2DZ/YfWfL5/JsbLid5PNcwk8puDbb6ZFs5F5+/OWzah0LKUI
bqwHd05eeG3R3U+nO/wPCmH6b3QJ92MvwI32KBERWIjORd/puPIts6/fdvCv7Hj1
LyKTrXzqSQ6BlwQSBRyIimGj66jonynllwRU4NXdowHksPS1mRc5e2QB+3QjxkxO
S84rOkDg3Irbbfz8GV8z6Qu3J6ASGPT1iqJ4BkzQGpQM+fy3gItjYJkC6Z5GZ7TO
UxAgKtGHfAX2/vH2K0nsXV+RlOz+tylc1ZgAf4Q0Qy+gXS2JIEViMxeHupCLB3oW
4j5XZe/kO/Gbmh5qhnhloBL3goAp+fR5/MAkzyGvnN2Tw188Rm7bjCVzKhTEnUW5
CcC7z278H5AyG4j/td6wGptbOC0b85tL72goBjPm5ttUvjUCw+pfpF/+BxvKPvWH
TEAkPShF5UVhyKSgUleL7gYNNlI8Cu4jqiWTW7WiZLefO9+U8dzgwYgyv+gwF8XG
ewXniKx+u9cy2DLWetEXRHeFWykigvScWL/sMvLNz2GFkC1JvyOdiWudieaoQJqe
lzKg5VYZWRwd/B3yaBwY1KCGEeOGpkmP0JjKf2KzJJMBWPwR5Ro+ydCSIaht1+gq
Fv7/eiSmh4shefK4u9p01psBZp7bdcXhrEaKjx5kfLv6GvLy+jY0EKugk9LQQ3/7
uybRH4Msms96RmnNFI3Bpj/b8+AEDtQ11yUx2uIBOps+mZPzHktkUQzDdNGPFc4J
qEuuH0C/+Ww+CxGQpiy9GsA5hocO2EiajL/9jVO6HN6FB2siPcqVERv5H6/Z4qle
0TC4KyYGeUSlWQc9bC0jUH/IUQH3PGPc/fUmB7/McBZvIfMnqDFbRrbt3Brdz6zo
UDxkW2ueWPbqF2aDisXM/Ec8NP3DY06z53t96eyFp3H4yjpgTtaeGMfJVcLMxVcN
elstTRLzHIItYqmV6suwBLs5Axf04Gp/SvjcNMghdSZiGq7JUEAVB9xOej4cbBf+
Yq9IWdSQKy1j80QYRK6hwUDk9cMds3lem33c7969XBj53/QvQOjzLcsnTCJKhMgH
2sxIS8ue0h2jzhdCCyjl3v9dDyhfMSgan0nDirV/TRbhaGO5nGSb5mZlQmZVEYGE
DdiViSon4YZU4PbVcehJR/IUKEQru9JzxbPm9JSInUJIjWrxpkRIlBBKlSxx5L7/
qrszvqEwd2T5ZHSwQIh5ZNx1CanLD1fHkkLd2DmvTaopfg3zV4/Ci3vIRR/noUbd
ijlkC7GUPH791vhkcfUcvcjtDsjV7tHUuYhoh5T2BMhwNvcqCWssu6gC3r33nXbj
IGfHnGu3i6DTdNEulW9b5FuwQH+MG3TRqOj0Uiq/kJzKNWPSjSl1xmJ5tAELtvcX
mVn1xvckDe/wd6oV+oPSOpvqBVKpBXKAKeQeRomwkq/7oZbBsyTYSvv7Ineaywd3
CW/PB2joRgsu0Vm6trs6QOAx6Nv22L58HP3J/032cuQQyDqktadj1GugoMZOW8kt
WLSPzXSX/ogZ+vmzXSm+Uo2tetzVDi82K+VDLuHEAFXTnrcDzeTc7xeN6uAVwz0A
PDZ/RNm2uZs6Lg5S/QXjKjYAeIS6bLGYX59SPNynEUux1LmXg+xo941Ov9a3go3G
2HzK6j4EecFxNmv8Pw+HBy/TtX9MLfJEeNiYzog5fS1bTEtrMGFh8RwvGvrYjtC1
Ep4BMqyyoUWHglE9+5xTo1bvTXC8RttvZn1JA0HtHi+157Gzw5wTa4NNHqCmaiX2
dyM7OgBj/Zwh1OyJxaNKxMBn4EyQNpxsu30Gjgd2//64YY4GhZ9CIPYg17HfU3G6
gA+qf0SZLShYDlBZvnmhzmkAyTKw8Pf+QMvKbrRhOui32Xz7v070+WmChaPaLftj
A/KSvpBuEDcRUcUyMdMDc/kXAx1WmR6ntXNZfMpCifZ0KrP3qtoNR3vCGi1FTmKo
P7IvZnG0dobbArnfbxgvW7meyzg4+qzDAZ8cF9EDCUNSk5Brj9cIrqbLRlq7vUQ7
phQsjBaxuLF3uj9WiID1Qrl5yn02Rhw0h4+jZsiDZnzsLobQqwTu2r8L1+3W1mCE
eLJRmR7/Vj++dheJHnsQuAC1Pn87Szwu6UXC/9A0OgCNlu7qJtM6O5JufjXQFb2s
b6bt4kSE7FO7hTw5FagFuHBj/21RmMaArtOI20Jw+00QB0IxRPln/SpcgNnnrC+2
eDy35+17RuJSdxrzP9FW/txrVJjzKfWsWpyCCCLIlzza/iqoADxC8fJdau7TARpV
9qV/wBQUefDSqD6kDjSun40xSR5Z6N5FMskNs7VgXmBVi7ioADU3VUquHEO9hm7c
ObnNb1hYT6S4jaOPO1Jpfz2MP5V878Xg58Uj11OmiCJsHCdC3MQqonRs5p3ZCpWG
u9uM9ZWolj/FyIHX1Uzsy+1BF8U2m/5lrZdlk26BiPGrm6GfD+W9D6eGQidZkg/3
eZ9v/fG4ujD4mfqYVGS+6rF7fQAdVbHaiiHazXtBaCDjjBES8ET5zNRpoeALMw7e
8eKvJI1+7YQoA+S9orJuUguLaI2BPQiyeSYXx1h5k+G3yx5AjnZ21rpb+5JuDDUi
GuwiZqgqj1Y9tt0Zba+p/ybKtm8mB7P1w/k7/pxInwFTy7R3PWb53fzK1ZJuaeSA
0itA0C4SEn5/KYU3EsOocTJjcgqZpXLlc9WCSyAOP8LgE3B81GVaTq1vMOKvsg7h
SIgO5HFNCq2tlmMuL/5DLT7AzCbWpZ8gP2X0XtcJ8jDi01qWCPBajxgoAz71O1Wk
wPN2YzsMU6OcQoDsk9wAMf2i29KOFoRUzrLDbDWbi00X1/BjIstRawh5JYvIBbt5
gPUzKytJMDHaBpSq3eCc/r+BVVN0BGs0dNZV3/e8Kz4pB6nBuRLew7O20SlLCeXu
lr4xhhInmWp8wZO5ykDVwAsUtbHAj5Ryl0Moe5+DR74qJ68xbsuEv6wd9inIiXAK
qz1BFWWLYcgZRxBjkdACAxkb+ZjHzogRDYV+1QbKlWzeeKRhaV5JzT3LnDl7MgUg
A9F3L4PzGWWvs3RHxAtkX+G39yR5rspzpVgxMgJjBj0/d8OxsI0vZHjUk7AZs9Lw
OF2zPjH2udQDiiCyPXgTOBbPkyLfhUMKDqcTBbePZXafQ/s6wO7y6PiHDKkHt8l9
7pN1XzjxalfYwzEFf69HMcwxdV6ElBQktkuxu6QT07kfMwnLVfb2ZGOTQS1wwjU+
4pXktDSUy8gTbh0yO8+XXLxmy9yCqzikFMMf1Dk0LGH1cyf5k+L1BeMbaTLezbWb
sNEVhW3d0enmqY5gBE/GnAXqrDpS150eUDJnxibvCoUzOim4jw7ICr6bhvOYdPuT
SS0HeU1RIOOdS0jX7KoRH/TxkWMbU6yucPGXWjHlpaE9WgwexbfUj88DN+c7mrcV
LcKmnVaK0Y7xh0UVWuMYJdnYwQf9+pinXzFP60xe5xIwtoNbVAW4Uhe1BRdhl0hY
l2NZaByndozOclUC9ZaJE76AUmYs2wCAn45VGqPjTpzC+AsjlSdxHDbCRb6DD+PB
vfUKG8miIHditU8rRIntcQXH0fiLr8cg//RnwZCfNK4UD2YZopA8MWD7v0P5FSJ+
RBT5HHQaqP8u9/faKOZk07GQ62DvY4PcYnX6HjJpH/35N7wsJ+9W9t6HhZOqaTKr
3vEaL7V/t1ybPyuIPC9/9jdxQFHhydiP6lFDT5k9tDhB4CzOP1iRRyn9uER34svg
zvQyIVprkUlvWhMyAS9TdKl4agHmVh0a0RZXNOepAWubPfV5Y4qeT+8szzmN1tAK
hHuMPNoCsEgOn+FfRGeoHMQtFkBjYzf+bUdqb+uJMP8JkziWf0wnRXr1g/Ovy3J+
Ty4pcVBSvzRYItLC7GSSssZygqEr1JdwJvkeMASw8WH7s3R6tZCIHwvsLXQEjDvI
sPJxKdHnFCnoNn/afsZnb9KCW9spiOQxdc19i0qW6R8LWTYTC0KwvzQV9oWq7kwq
3iemusFYPw240xOCWQgmkeVPGVL1L6iC+J5urTyQ1X8tXca3/KABKfShKpxIyvWE
oMlredn9n6uBWnWBcMRtg/nmhEeN4Mq2GoNDfcjM2lzJpQZLKaIIMS+5VC2IzSl0
SFyHh97qoiOm2TFJXLRBhvKtYozOKhOmPATwCtkAIgS5i9aNiGQ366k7pMBECwCE
PGD0pMixjS9u5r+NeSdfJNhiBXiKuIIs2vheO4v0heTX5Za/NrYjmGOP/u+LSHbc
0Sb5opPnfPDNjdE/SbOyPG1Iqqq2eDgzwbVEzha4bZw2HggsIZrrxuYyb/DvROLU
qkCPNVGPfeU2k2RmVGew0RyQRstRyBVi4BmQHkENn0OA4E8J9ZCKPodGWXTFYqd0
pcqCB2WPGOCkpepoPgtd0l++HUnko5fbEuxMGVKEU8BN9N3kkKYKrNfznzgc72Xs
A+GXrNgy3u2ZBifYjS7SfDTxxKa0JwESOFjS4pirQp0c1OOrQfJL7347fQFr01T9
wmqegXF0vZSR8gY6BCc3lJI6JuF3vwpAfJeEexH5EmXITBK6Y/9w8JS61g+5Hn40
uOg2toV3xhyz/0I6FQCGJYgG4Qfxc0Vgcy69BsuFjqryyGlD743xfg1+4unUNlKo
nldppsmFAoHR2rTMh8jQYBdRDKUKjfvl4Vieo2HM4Ymv2KulJOv6hV+CHe1ZfIuU
vG9WAO7cBaUz9vpLPgbjVwIj2AkNzg/vaHqpbWzLY68Wzd+L8cQat0cs6NvgFhRu
KM6I/nT0rcLeQ0m1OpyKR0qWdONccQLq/PHboSQJyC8qeplg715vFY+Gfp9tcAyY
ebEJl58pySxTQk3SznOIyU14uGRkc4Orrf7XOpNpJQpMtgD3zCRMIabwpCRQV882
9xb7eZPlxXdinJNeZbn9RcSlqXdpXd+6NjMlJ3sFr87q+tjGX7G+t9Gn8yxZZ6nf
J8y/VPhH5j58kiZbLBQjC5MxnBo/lo97+K3NRrbhzLlzkE60S7q+6fXgra6WKUhm
x8bDEqZJK3cC5m541B+xZJc2S+Sh1foEBlAmyGt5hZxnbOxHNlVSwOGS4a6F2ffo
ffFcvJnRUxaO5yIE3s2lNhH6+vQK1H/CsD30CknHRW7Mz5RUk3D+NnurYSzr/SsL
mSJezEJpFfo5jOlOF7FPRk6A+jYPjb83/JnwTjqVZEueJGDRNC28YjXhkiQ8h9l4
wcGOPokNH6zvo75amvkd6HQothX26C1AA4bJIOGFcO120e0FY1kAAD+G44INq3Av
Gwle5ejwRq7/3fcG0HDnT30qSmuZpdxGYhK/hXIpDp8ivQ89wV77opm7cNc+sk99
1aWReYB89Xy+Q3c0NfqgN+JnOBKVvu2dW4EIJdmAfOz+sDn3CFL8uon91YdWS07S
0PM+4/MqcHQ3zFC0xpS9u+gC+2/z40X/pwWmsWG6YWS97foXbHbvIbTQfe5KoEKH
A/i9S89WDvJMWFkjAZfrswdW3uj0R2ntDv1jraPxcPkcpdLdBTx7yzsOWWYXcaKm
wZMsJ+1hbYk77VnwukybTeVafkPIfhNifSQ3Emtw94qTgywGpQCXpDDwCnVuly1s
PDTkIjwhmVu7mhmfw3pSwIylPPP74QNuodQlCrr2i7B4HJ6MPdq4lngbC6hOwP3s
uk0odiDL2rM2rUk6qhMN2zTeYte/XzjLGCNAwzJnNuZMhEtBM5R35YZW7vdjD32H
wHNFRAVivlNJUj2B8SqSLyyamzb1vs0yVIH4f9RZrM0jEhAD5d9WciqQZEK6ZliU
Yzq2h5uX5McswSYx0OOv/mpPblQI6SuSSzR0p6LqrE33pd0aodSlMi/OHJJ4EZff
YXmAVGrHEpHmAG22KmAIcGRiCaelYIyOVJoPT0DlaBbS8Y/oSp6me6akqNwrzaoq
rvAd6ouILWg1vjf1ChS04XL6JXbjXtV65DAHQ/IgHbbDTqs2ARNwXg5z6yfovlZ+
zcHBUMmKrQcg9N/HImj03KRxWA4wxdEtB2HsxW9AQvt0xeBvz6ImXRFjbGslr8/Y
7tRKx6nSn/blRXzsKgNpocUrSwCqGeHHZK8tpSrZYVX6Gec/dor4ghDtibuyMwqR
Pg1jxdFIHZh6/WPbWVjWPEr04KwMs1H7020GheiSYoMnpDyWIYpJ0OtncDjDzyNP
oD/kYJM8Cmp9tbFRErLOJ9V0h2jUi4vqnXQ/zyG7Y1YLJDzsRJ1kDQmbBJukVSXt
b7i7v6dbM4CRxfqz1j2N9mvs+HoSd8/UDSmPmimgw4mrgBiIIwqXkT1An0HOLUjh
7CMeBzti/bLJU6nZV5zHdSIh+8pnkGteescK7mT6+1RhbG57RnhZwAOkdwVQh+8x
8wC7/k/3kT+xIx+Z1b6EPMgaBWGKt6cY/yR/qSb/54xD/SB88gFbtuPJZFZRWp2w
NSju8IHGW615jubHzF0yG9TSbPnJlBpCamGWXWAfr0c4ZzCDfTKe3VwQDx4UGY9e
qxnXC1dncZO8v0AziYGDKr7BI4p9nvIXM3oBm2x6oUu/xDUoM0CpvX3m5jqJoUNH
jlHzjPwlRmA3ltXbOFsMTwAZ2k8SLX1VRscKnLaw48FAqtbM2c45aQs/hJ1rW87S
fdgipDjff89JcoTK0SzCBENEkmb13jo+y6T2qbEHdtlPgwtVskbkgzEhkH8k3ygH
KA4K4l5fJ2KRjGxl1Kw2YVx6LgvbLSdVWrKLJW67ymQZOPnxYjZ7/GCzpVo1nYG2
z1PMlrbO98AnNTbslrxqHS1CtbtFZPQvbOTL6KE+a5vJZx0VZt1JUqL7DZXun0gF
Jom1zrHyNWP0QF615gFflA==
`pragma protect end_protected
