��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���9�{RԱ[ж�8�����������/a��:��#Շrb�,��Y�)n��M��Ӡ�5H�������w�� �Gx� �Vg~�r�5�t���5�Ш>@�t���57�s�f}U�������2'�k�l�E�g�ܒL�������(B`#�%��ǩ��b�y�ّ��o�ka�0��4�~u���͸c"�x���3_�XlB���J\f��E�W����	�]��8� HI{�s�zq ���s,=�G�:F�V����Y�e>�V4e�i��_�F`�mg�_}j��&���\���B�꼗5�%_����^��Q��q�o
|�zyFB	�9{i������ag�rʲ5Fe��Eó?T6��}��K����JN>Cgc��Ӛ�cH�`��(B�� �l��j�*���gjdų���\fٙG�%���$�����tXS)�N�����f�td���kt��*ؽ3��t�����-w��^XY���L��K@�Y<&��F���F7=��g���=�p41�z�Y~��%dh~��5���$/_,���\d���b�J�Jc�i)vs�L��]�U�Z4~,��7E,�~�<�bЄ��
c�B�(/��kЇ�6+���?'��X-%��,*Cd\�H�QJw��Y��)�>d*5Jy/�����֌��%�G(�^`��R0hL�U����v�A�k�3uNh��V�3SIK9�X2D+�����ٟ�`3ѝ�6&�
*��G�ӗBLc ��0n���m�:Ҵ|�Srv��?�Ь��P�[-�?��MW>!Oq�#���gXݤ���LL*�mZ����"�5��y�}Q:���� Xb/Y ��!e�ӻ�����ư���l.oLb���"8�22�U`7����L�[�����,d݋�0��ċfjXb�C���
I�9�70���Ivr�+�Sx�����N�k �h��fZ�Cd�t��ӁuϮj*{�Y���!�V�铴J��z�5=�f �� ��|�}����g�l��X���oxӸ5-w���]�m� It2��F�
�z�@����ݲ���/1c���I ݢ�/��+�p���rk�I�>�[��˃�:�2��ߚ�vԔB;�w�t�PTUo����@q���
�~������1�KRj9�E#^���MZ��z=�Ϙ�j���wQ��K��oNm��ǿ]&m�:,�+6�ͮ�:7�#���=��P��>��ܲz���v�^ ���U����z�rq-�>�������k�ߎ��R�
��%��V�9�y�:���\�=�yPR�ץ���v^[[+�zL�ite����͊P��;㏅k"����Z�j8>\J`��|��g�˜x$II���S�)![�َJ!s9GF�9��+��<9��\Y/�@3V�\˻H�Cn[g����ks�����CylB����7&Zؕ���0���sDq
2��~�R��uĊ)��$����e�@�r�vVK��]��2j�Y3��L���Mk�������Z*̛ۖ�1b
�+q����DE��\ȼO���`�λMN#�E��z@�z�f��0���얫fD?��g&��������]�)�,�ˈ�\c;��J���0S�ڮ�,*�
<I��P�O�,�7s���las�;{�Xƈ9�H�i(������������Hp�6����coV#�G���6�p�)��
N�'fQ��.���&$)V���bgV%^����lhWLƹ�碞D��öWS�w=Bn���k���#�T=r<��=��������>�@��g�̴0f��!mS�����ń��C��=�oi깚���xA�ZL8���&*�*��R�c_,�=M�/Z�k��V,��:�,K� ?HY�͹��w����I���2�cQ�ia�@+�B�,��|ȑ��ЌL�J�M�?�^Y{�� >⏒ڨ-,�YJ�N�a���݈8+�	��F~�T}�Ѳ�H-t�&��]y�k����*�)��(o�
�9��|ʑ-W�L<}�
��$ps�t�ګ
����0�5Orү4�0o_L�քg�^�N�=�W����4�J>;`(�|r�0K@I�qg�7gc��{]��t3�9RD���M���|Q��5(z0eq"��%kf��<��h����H5�H����
��Q���,��~O�%(�\?�� �*7��z��,�%�Y��蜉`��k��=Ėh��i�J�!���t�9U�4_����WW��c�%z�H�a�ѝ�(����`�u�`o9@�2Ia`W��䈬r:&+������+��e�8��Im�Be��^�ߕpx�g����<�!'� r JC�j�֌֤B1� �kb��_U�Y��n"I�g��e2}{�#u*�$>SA��זV'�bBG+-�y� ��;�S���d�{�VVʳ|v4��La4�D}~*�*��ĭ��H�wr�;����q�{n�!k�+1������ `�� �s��k�>�"y�-���p�!�;��,�V���?�,ο�2#S>��G�4�[��i�js(�eQM���5�~��&����J帆�{o�c��9�xqQ��M��g�X(,j��7K��;�L�~���N�d���`�J�%���CI֓L?x�S�*&kF��U[B#'q��1�u�������df %��T�.�����`�ZnT�~\�Y�=��ä����b�	��l%5qvy�A��>!+��hul���{!���K->�g�ʷ�e����Q��f��~�M$e�P�h��f�
��&眤ӏ*�*[������mZȩ#��s�+��[g8>�������e�I�On��f~ �V@�i-��> ~�'A��'|����R'L׊b�aH*,�eל�F�6��V� �uuX�n/�pl�߫b�BC��Yb o8��k�fF7§۱�*l�_~���`z�m�+�����ݶ#g3CI�<q��[�*u�U},���Nl�b���,֬��&"��(�f�. j���ZY.H���CB�;�?��[���za7��1 ݆��6���
� �*���%�Rh�t�Y�|��!��6�̚V"*�P*��Ò�3�f1(�<�u���f�mIY\s,�x��O+�U	���=�����-S��+�~�ơ��!��}��H�r�H)���4��<���Ѣ���_��7����,���1AQ�*�[ڳ��a\,��	��"�3��*{�,ap�t2��Gp�#q�)L?�Q�R�����Q�\��2	3�`C&
�A���.x׋'��Vo�CR��}��}!>�e/K#���b���!�z�b���u��{=�BA<��F���({;q�\8=���+W����ή7(`��|@n�h�ǠRf�dMn�����
$[��!����}�f�&�1=�y�l.f���Y���\Yϗ�U�� �q�^iՕ<^��h�e�0�������ɶ�k�z1��t�_�%-�?UK��ˏ�Jfݭˉ:z���(d��O|�f�T���������Y�!3����ǅ/%����,(&� XJ��3PH[sĜhD2r�F��!�^a�����l>HwQ���ґN��d�%^h,�ϡx�?"�
m5u,�!wʏ!��,��i�c��\?�� +fI���!�!Sy����y��l>��x�.�I8.YXs��w
�������
�!d]*��X<�]����4�|���6E�]kYI��@V�r��+�d�k:� 6��Ka��sd>�*w[�K����'��ַob���&;,��H�z�U�g4!�B^sb��ݘ����.����L����ᤤ��*1����|���r º;��H!�6I,���=��cy�p�pb^j;����lmz��;�E!�.��>�-�>��T?� TE Bխ̎����&�<U��������&c��W��B�Z�.�!e��Am�wyY. F�t��B�S��Glh�i�dg.�Gӫ�m��$"�tq0�Nk0ф�'��NR��w�&��<P�QEr�D�%��1�v�cV���C{h�%, ?/6�9�J;%��J�~
�
,#Z�:ކN��N]�E����cW�|��W��`��="r!anE|-p�n�NC�)z�Ֆa����o��.< ��4�TdD�XZ�o��,Ј���!�%�9����ݎ������Q��6��6�������½�����K٬�F���k� s��\�v3Y�9v�&ʆۧ�[�i�\����,�AZ��13��~w�����	-�J��_J5�2H���E�N���P�39N�<�gus��#H�7�ɌvY>J�Ea��$	0;,CRN�40��ݓ��$e���4�ye����~F���LH�d�Ke��f����a���n���e.��<&��T	�g�R
�#�=���6�0i��}ڌ�04��_�D�� Ld
�3�P���{0��v��a0Hʒ	�
3W��>2�����o:����A��g>��K�w7c4nP����mB�sR��{�v���o��a0�׳���J�o��="��7�S]�8�������aU�~�������L�����.
�頣� �p'��S��ApS������_�?~��$-�"�o06{�ތ=:���^��o"u����o�� �ZnEQ'z�\p��^X�cU�;�?scwT7U�Q�[E\�B���Z���{)�\3xX����I>'�LL�{�F����e:��f"�j�ZNW$B��{S,���I��xl�vt��B1Sa;An�aȐ&�&/�Et����Hw\u�k�%��v `W�~`+]B��¸�M�Ab(��Ev�U�hE`��H{C/twpSɃ�fL�rʥ�������Y�?��s?f�b��X��!�=��9f˦���b8�.[q���c���_�V��2ެP9o;C����EPڤ��.�78���X�{gx�P ���b�^�z9x鞮<��b�L��^0�6�Xl�!w~!,;�*x#�B$xӽ}D�x��g�qz�F_��.ϑ��yIt?K�9�=R�K���/�1���؎f"� ȵ�A>{�v�2�@���&����O ,cjI"�x�/�]U<Ԋd���9�S�_��J�z[M )A���0NOb7�s� ]����j2���k�k�Gr�,�ڬt�`	X��]���4yC���ڧ� [��׳�7�G�
41�j����Q�������o;��'��QJ�SH��W��^��R,@?��0<�]����tS��"%��WB�LC�<�V�\:��*x񋩫�0�UE'?��?X����M,MO�5yg��
n��"�0T^b�.5(�[�b���
�;,=쒩��;c2N>4���,���L�x�B��8��� n�rhT�� ��Bg��t?�'�!p���JM��I����8?������ ^h �A*���A`A�K�����|�Hw�4i �	��>$�Bg�+M�-��?=*�+K_��!��J�g��^p�x�8����r��2���W�}0�u��h�:]YE�3�6�M���
 EZ��8Ҵ����yI�t6[wu�&���j;��t$-�Z���ȰK�O!b�FDs��{���p?'����H2��`Sy��X�q���|CX��v����
��љᶟh�ܽ�b�FS����w��|�&	M�2��p���u���I�i�V�t��p ��4�nkn6Ҽ%EJ�ĳ�Zg��?�V{7�eS�iJ�s�l��r�������4d8��4����v��V���Eo�t�م�&Qc�F�E�9Z�u���W��YJ*�����'�}9c�Y��G�6��Т<�x��aX���ү���e�B~��fV�?�J�>��o�v���j~p�q(�Mk�u�ip{��T�/�
ЀK��4I<�νo��P�t<,S " �S<�k��?&y���COΚ�Q��\ˁ�Y���!R�g�I7�UR�=��Z-9{ءb?o�.�Ib,��_i��u���	��y|i�C�����%�b��=�gufK��fM��Nӯ_���G�N��y��Nb�SW~�d1e�6q����T��_/�2oZy;�����[��E�k��k_á����np`1�~�iO��0�,���0�@�-��������r�Țu骜QYxQ�{t-�3Q4b�׭m��k�IL���3k�R��sm��U�Rc�70c��o���?���u�����Ĕ9���ك\C�o��R28-�"ac�!<�gq��$��Ϧ�il�)~S��S��M�Y�X<�j�d��BC�F\��(�k��=�%;��{7�������'�D���+�ZP�_��3�"��]i��_k8�<NP��S���g�����AH��_�L�W��ԅ%�S���`7z�m�qf
8�O��o�V�K�.����^�V՟F1�sp9g�_[��ܱ����)�VUE��Y*�z��=�=z�?HH쮈��P]�����HN�z�����*�͐�"%@=O�r�z�L��7����V�e��4E���_j��D|+`x���1�	����9K�W|��4��f��'����j0��M�*�o�HS1�/��
�I��'�����m6F��^�r1,IR��>�Y��&�q�@3uS���P�3I��uC ��)v��}�>�.<zfi�7�6
��S/ch[��߰U<?�Vk�<�z�0v�(�G�to�|c��� O��e�y�ZW`ԤS�C��=rܤ�L�Ir!Jqx%"�;K~���U���aQ��A�LO.��8�(!�(�����dtW�!��Br�x+��P�a�`���a0���?�A��m$�f�>����3���UΓ�UO�ׅ`��fůö�v��K�ŎM�Wa�T���зQ7錜�1f_�������S���e:�mȍ��,�n�)əoT�s�9��My�b�yJJ���E����|%%^7�8fPZŠ/k����7I\H��R��o��h=[��n�G�$Z`q�45��3�w�ڣ,�b�Uv�1���0�h�ȋ��cS���gx���v\�.(SS�C�Ny�Y�'ЄJ�,Bt{�X=�`y>�m����c2�&�6}_�؇.�M���C�	�>B�9�w�|�d�ͶԼ�9 l;,toh���Hc�_��Q�����7��G$q1�"�7���DU%�%aU��f�W5X7��_yo�A�:��c���0�Ό�(R��}]�
{�Y^k���yQ$���.BÖ]���+��l��Y�A�Ѩh�����.�~*oP��É��q�"�4��
G	� YrDS�㧷�`�:)��>9Z�R�-KRD��!�_ؽ���������$^�t���ppM��ߔ�}��At4ǘ�%F�l���>��r�~�T=�S�� #ѿL�::$J���E��o��f��;W�4���������Ѵ�%:1R_�l��K8�r����jWM"[-��M"롋�"M	��@u��ʌH{~�����m���P��ݣ\����gԥ�؃tu�a�UE>|P]U�jP 6�|�*�h~��8��P���+��hg�p�4i$���9Ia�������;dBC��T_Ȭ�xĘ+��z��-��,S�NISW��J�U-ns���@D+���>���0��No-.�{xgI=G7�����4��H��-�s�~�;}	Y��掝�3 R^CP$�Ξ�uF<.��GOv��쬂�"�{ E��ޤ[���H��坟��U�*Z�{��P�1���7���|�n;�r����B�dE%~S��a�LΞ�A���u��W�Wֵj+��px���0��LQ?ݖ0��T�n�_Q����l��w}]^�X���3��� .�Ԥ���y%NH]p9�ް���!ۂ�%;��ЁU�3���4��ptW��0B`��w�;*Z��W������h�Y{�A!ߟ9ΝC���W1z���yL�>��)���ȝ,'�a, >�T���9���p�M7����jG�2c���<�EM�g}����:|A)\�p��,
���MU��,1J���*hk���+���-��%��n�t��R�ᗖ~EG�D�wk��g�'�4w��i���(�]p>�'ȐE��,��+��7T(r��}�1�;��Y������:�=.W��� ENnd����Ʊ�޵{�=N&�>����Xhm`?����x�).��V7�S�G� ��m@Gx�<��R�৐���ܩ��7�Ѷ�m
}��zq�n�t��H&ˡjd�Ug�K�|��� �!�(Ȯ�me���_�@�g%�g������V�pb6�{������?�p�"��>�fL��"^Ɣ9I.T�FS4���Q���#SZHf����L�+���3!��y��|�!#���¬�^��҄�����dVO|l�C-��7#8!��m���'���>󖸅@3�R�o�hY�6��P�ʸ�l����t6���+= �7 zB�W�+/mH��nBFb�n�5!�|9-�<}뮭��~G�.`ʆv$�h�R;�p[�=��@o��)��\��S�w�:�=��S�* U�dH~�qw�a����]X+`�ǶN����6m`o~o�E�ʆP9���q�J��d`mR>���S�H'�А/��ݚ�>$�lmm=�{��0'ɰ�������:�?�f�rA�1q؛ĉ��(l_�}���tWŁ�vD�/���(�`-���F���ɷ�>\�	�$�?#�̸�JXo����U����@�=!��)�'<��6������7i<A�����)���m�Ok,��{�JR��>4UI0��G*��̥�K�{J�;�%WoH�L�1���v^[Gwg���.w�g���?��Q1��+H�yT��{�()�7��Dz"���8���2<'�����/��z��Z�v���0i��[�S�s�L�烹L����Y9	&A`C�삯���:�W�c��6�u� �VH����6��=XqG�W����Ř5�M>88������E��\���*� �X�1b���4윂����U�����e���[��b��JUE��o�~g��rc���i�a�]��Fy��^����«����X:�lX'��@FS�u<�n�y�Aj��X`VL�d��Q0�`G��^4�]Ҷbvh;����w�wlC�o��3���I�Ո�z-�/Fg�X��(6C��@Gm�JO�e� x=V��Z%E"[�)Ib����o�,�"��"�+��.<ȩ�e6%j�<?$Y�%���v;k���D�Y�>����=@�nS��I�Y��>XV.O����,�n��
��O�
��yN����)�y�G��$
;�J߿/��(I�2o�L���as^L�pI���c�=�.)� `Y��/�a��:~��6∲E����ҿt�K��q !�}�T�q�+�3�ҡ��;�ɼ׼��� ��Չt���{���s��b@�H2�f�l��Fbξ�FIz�CU0ь��41XS���2(�,̋\��0�GOn�#uN�B���u,!��\/����Ң�;߀ft��Srԑf�eB�~�����0{ȁ*T� �;�2Ee��n�>?M�.����"��)���Z3Ǐ�(���ad�u�I���x��|��cO8U�	�,�L���c
T>|a���E2�G[V� �/����_�vy��y���p�^��O���*c��Ϛ)�+�x�v�����;{���!:J�N�'����k�W��My[�pt;}������F+�" E����j�����Pf�
Bb������Q�R}��4��<���5���7x��MZ�+:na,��+� �GBU򲾼�ҵ�>��3L�G�tbe������6Τ���g�o@�S$V��u��!��צ:�<�e!iט΀öL�3�~a�YθkH��u�-���I�4XW�nM�B9SB�ዌA��l�+ذ��$��G�-��'z���1�Yֹq�8X�ӄ�O��:�	�����H`v��l~~�L^B����_�iʗO�7)���G4��GQ=�ѡ��������5��ڗ%���e�:�=�Vf���B��\��F�$���#){e�;>-/��V�;����;X�4z�