��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]ǂ��O��˰�	JL��	���m�T]Ïx�R���L(t�����~�x���Z����Z`FٙuM�.�-BOS`�I��|+�=j�f�̏�4�>ANd��� GF�73r[�
z��l)��V�Ʒ.IH�F5P����@M�JM�c�	lt�Ӆg�/�+�h��U���ݮJ��o�n0��R	�Zv��cTYaQ�vaT��L'�E��LD��c�K����A�g]��� �SI�f��_4��Y �=V�[�ũ�#杘C���6i�|ı��T���g%�t������J�����t�ii��&P�9�J�j<�4��5�ї����͌���Ҩ�A���-�{��'�1}+1���'}������mEp��~6#�Iyכ}=
c�@��迮��ў�kn�
P�X<X��ɨ�dc@Ps�UI���j\�SW0B�����+�����{؞4�I��j?