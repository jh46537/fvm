��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���_���W=1����o �6!�z�O�]E����6Scu�Zz���6�T7\˧��5ųkzO�-�b"��7��f�pC���i�N�ϐ���G��ܥoh���<gԎ��o��}zuM�M��ק�!M�ِ��;�U�dg漍��n���|~Ad�!�ġ��&��q9
�o�)���#���f;k^�l�2�@��z��æyv	�`̶���NH*��A&e�dS�S�gE^��R�e�L|m1>������)�L��<�y%j kZ��5�N�|ZJ�����+J4Ї�&ĸE��Ӭ�⤧"�%�����t��B��v4�Lp��>����<��.�F��K�M�����K��؏i �~<"��z��d9c���*��L�s�7��P���o7Da�R�O�-d�I3)r,:���%��GO�2�üC�F3�{\N�^;���y����RE�z`w��<��[��A��B���w���w<t���Kjw��+��@����% R���J��X�T8 �I�R��%|ń��7Ӿ�� $H\�M�40�"��r��|\%����2��h� ~�";����*��>��!�F��dǀ�r����3^�J�S�-+�]�-< Hm}$+��D0�S�Y�d�,�m��yOq�3�����,���	� ��|Ψ���[�Q<�J��,��(���~��#��e�i�;7�p.@�z����Ҝ>�,u�o�ۯ���P�����K��Ł�g����z+5�^�M����ە��n�G�I����,GBo��c�F�6*x��浿@�E���M�,b !���8q����ߧ�����8��J�w��v��\	�F���4��.���󑞸u�S��M���r}�I.�(��T�ӈQ��������K�.��A=�آ�xŚa��>6|ik�,�Q�J�5e
�����=Jƪ^s���>�K�s��0yS��\��FBb�Ef���K�]Үc}�=�� 5�_��y}�L������e^w��c:R�t˸�X��/��j�d�A�d��F�(���s殣�N��:�H���8��hy )^�Zޏ��hں�������)ً����� ��R`��u]������Yf�c�&v N��4�:}�;�jڔ5X��vXG����=�p�NQ�Ar_9b��j��|�����	"N��� xSFȆ\��6��A��x�m�����J���qbȞ����ݤ�a�60�;��ȀZh�@��]�� ��;g����Bo�"F�&�9���g��|[2T0^�%�Ds��'�D'F��gm
���9Ls�,L]�����D����Tn1?�.��<�*#UN�7�n��J֎��F���Eˊ�."3
�2��Tw+���P���0Y'S=c���WUV��5��ƻ:�V�������~h��*�a�����S�*��Y����C��S�m����R�H��Q}ŭ,I�D
[�ۈ���V gܸ��ڇp�ˡff�,y����/@���_i���^+SMJ)�60c�\? Z%��G��+�.E|���Q9�Ly.�x� ������c��b^�h܌`�ފw"���9Auoɉ���7�S�$<����������d� C:��2�}`�ߦY�f��9��-ʓ�-�e���4Z"�;�Vr��8�:������X�R�