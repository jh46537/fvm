��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)��k:�ث�����$,�:YƚN�bK9�p�IV�UC��$�Gǣ8�yF��D^��a5�{S�&�`l��ve������ӄ�d�=lے��+��j�Y^z�]w�#�k����u��0�]v���ޓ��#N�ݔv�"�GZ��>�:��I��
>�c��6|�OI�����Y-d�S�={&k򶾌��禩�}c낪��3�Y+��k	e�����תа��d�K�%�0t�X`)ϕ�H�k�c�f�������bN�H;L�ɻc�DЍ�ª= 5^�	��f3:8Qq�Gړ��^ߧ�U��@cFj�ط�	�C�?R����5�`\�1Ǵ0Ie�X� ��[t������X`�.�[�]�fTۦ�B��C�W'߭)���⚚�YȰ�ǁA:��њ6����R��;���p�;#5��|���"�x�(	��p�ֿ���d����@����Z�8(ם�ي�5�12QHKi����I𕷎��	����&#�b9 ��ܬV,�P�"[6��[��tU4��:�{i��8w56��b��_׆�L�0zXܬ�1@M���mB[�ɘ&��:,~vK���߰�&�������X���b�c�<a��y���7$��U��b"�В���z��Ȧ�^��'�۹&o�L�'fz]'�,,)��h0�K����Ϋj�5(rC��9��9T����;��ƌUtg�ԥ9<�f��v��\�ե{3q�0��s��¾�"N����QI�,v�2���Y����G���jL�p�"���/Vm�1��w��Q���3�24a�����# l%U����JY^.2����ǉR`��)|��\y3|��m"@z8*E����5��#J�^�D~T���b��R%c����oL���9��g�����M �ae	�_��h �����p�]4���-���z��I�S���q�b`ei��
��a�JV��Y~��=\ȼPQ�Ϳ�c�J�� �����F�:����:h���f�M���	�����//6i���Üﻬ�[=��㉈t<��4�p�OOΖ��G�)�u`g˩�I�E�V��w��	3|��H�ҍ�����KiBEO"�|k\5�*[s8qPC���:������O�|���W�r\~�Y���i�?+���p��0N��׾o�Ci>�rj�;��/Ҥh��������܅�{�J�4褎N��ܩ��-s��xH�_1A��rӵ}0W!Y��%<y�%a[�|WsC�����X,y��\�b��_��R���oaf��a��:5`Q�����灝+4�TDD��9+]?C�����gwXt��v���BU9{O����+����z᜔�ҋ��o�Ƣ0���pJ����W��z���	ha4\Ym)N�d�˩b+9mW:����%�� ��M���	-�6ily��O9� ��F-��H�+��}'�%�C��G�Ö�S��`�b��Zh�r��%%����X����\���6���sÚ�>V������z���`j��h~��
N�N��7�Tza�&uYW:��+��I�͐x�(kH�>�L���wG_,��EXD�T��;ܻޗ�nj]8��_,�$6���&�������^�8 ,~��5+"�h�`�^���X�z��YAL���w}�Wě�2~�t�����C>S�=<LC�o@�R�		��[n���x��n/��%{�}V��ՠ�p�lZ�E��{&Ϸ�np*tf����H�4{��G�72��H\��T���Eu�X��-M�V#G�4����C�;�&%���-M�H�B}^� Y�ۥ��E���[Ͷc�Ş�� ����z_3y���0��y9"�H��Cfޫ�!��zz5u�i�W4�w���%[	�xwHA����D��Cq��ڣ��N|.ڏVU����uY��Ȑ鸍F���Ġ|�[=kpP�mrب�%t���&ڙ���1�3��jq���~�4��~�\�jݒow9di �C�i����ۢ���9˚����EA��yg�[�i��!$������5���J����P��(������USd�OI@�:�_��+����������֠��(Ag#��8�-�y:���۟�h�=q�u��l�N��`--��Z�$E��k�i���e��%,�I���@&@�a��f��L8A����� M��_VW΅���|�&k5a�؂&S��vƢ��3\>�D��ۓ ^=;{���`�kd�b�4�w�d�k%y%�(�(����U't�b>�����?��̎���|�r(r6eT���2�U�L_&���@R��<@*�ԥ(��;Kxi8�외�����5o�rNF?^l�E��`7i�ф�w����v)Rx�D��s�Α�����g1
+g!O�4��E�RtX�gҪ~�h���5�fv _�1�T��
[omOj�����nP�o�%��ѐ]ł�1B�����NX�@e�ጿ��0����r�H�xx>�}0��I��Z�b�H����#$�'�m���`��[���cQ�#��j��_]��`h�d�P�v�����Hק؛�� T�	�b�����C����=�d t��E�^��.7��
ܨ2V��Hn���^ X��۞G,8W���l�7���j�z����Ƞ�XU��P���rǿbc�n�<�g+m�l�L+cTģ{�-[��f�ue����#��%l�_~��C�]��`PB��`�O�?��Fz���*�"�E5����[� Ӄ�4{V�O�j�8Aͩp��^Y���V�}w�sP��-������e��o����St��sDؼCVֶQ��S����D�N���E%����z�).f�dXk�E<vy ��C��%5���䞟|�`���Q��ChY�y��b�� =��L�mS;j�[�S��ik̢��J\����b�������뎨Rw{Ot�{�:>�4	
i���!����Ҽ�n!)
���*I	��tӄ�f�?4�ն��eϢKھǐ��K$��|{�TU���V�~�-Q��?�n*6k��ؤ����9ܔ�ۉ��6�}�m<�j��:�������^Ѽ�)"��t ��J]�wd����>��_��}�J
'��b,�:F�f��[0~�A���C�������{yw�HUw�����:��n�a�V�k���˨�$��1����j�d�@*�<cn�����y�_L���Z^�y��s�a��3ÜO�z��@t�˄��et��5�]P-(&O����~�y~Yk�  �v��� ��9��lv@�"��Iq�s���]+!<Њy�?/�V ���/)K���9:@�u�xL��5TqT���m�3WK�/������"a��[}�����K�;�yc��mQ4.��`ݺ]��~��(o}��3>�֑��f��07���G�lp�*+�\����4��nQM��I.1L�Y �T�+t�S\�u�H���1ru�e)q�����N�����T����i�ᘈ2N��aZ�H�Ơ��Ņ�f�{T��O�׍3""�����W�P9��@�{�kF���E#C�y�:�!�2��te�M��MƤc��@�(v�>���Lz*¦�+F�k�q�Z�Hۂ�V�������"f.�����<k;B\Q�}��w�Lb���0����Ϛ�4�t������Jڂ�ӣ���m�M��F���C ��z�6Ҷ/OZ�}~�8h`LCٜ5�9$�łQ˓����Ū
���NVbByo�b;A�MrN���S��
1���`Ho�)w�O����
rT�V��Z$��=��y�J��Dg##��UG��h6)��	�^>�]0:6�l�+2(��^m���Z������8��1\�<L\T�,Z��/����4��.<)���A��:�t�ߞ��U��{�χu�A�?�NT�c7{P�#���N�X��Y���"��[��D�V8�7� ���r\�#/�_%��Е5X�z�9�cU�fA��uӗ'�qRoc���zgBC�i������yTm�N.�8M��H��1T��I���at��`�N��괺%讖
���G�q�����$���͠�!�o��]ſ
0!Mtxe�Wf�۸�We�+�S�McП2籙�°�������Q>����:lDgh���:�Hq�=����<��Zc� �8�Q���:5��i�\�׵�¸�{6�#��c�b�:��Ѣ¼is�{M�F�C�N%o�߿0�ȷ/�Q���,O�G��R��M�Y�+�8d� FY�1�d����&��vI'�/o%���pL�-���B�<��<��Ҋ���xmU�(�B	7�Y_[57
lW�bE\nٞ�|�]�n>�)�Z�6��j��9��$9�������*TY�Y�4�H�J5"�j�@����G�O4MLE��m�a�O�"��97���{���0�)ڤ�����
�n��?ؒ�Z�x��JYaP�C���e��A���a�AAgK���|�����a�d��4��
+����*M�b򈐱�;d4q��!7���)3|�]H-
[�s�*�a�`�#4!��MY]��y���8ش���=���7^���Ϯ����+z��mt�|nA�`(����"<L�c�d6�;�M��_�3M���$�hfw��X�ڣ�{HQ��8���h엨��=y�Y�tG�2I�Ш���)-�}�,C��3��+,S'��16[�D��d��W�3sc?
T�Iy_�l�0���xg�űe �p��-9��K�
<o� �����`*�?{?�������7�o�;^�6!���	H�K��Q�),���Q;�T]�0���X.IW��c7E�Fq��n��~5��)c��>e�E��<���o>��ԵB�}PD��BY����Z�k��B[�A��{�Hӂ�j�vf0Q���XVc-�<�
-7��{(&)܀�q�@d,8�Qꮣ]� �+��`C�����9A,<��Ӏ�<��%O�bp��sX�A|	�o�Jͅ�EǶ�>6�u�N�֔٨c��^4?���6�����'�yq�79/E�O��1(�+�	[N��V�J�@�9U������m�����n�6f�+(X�HH�;CA��/>%$v�>�^�|,�{�_K��/��-�IHRǅΥ0��ZI���Rb<)�lvݲ�L	�16�/j� t�,F��v!1م�\F▝�T�׵�)��-/���<�������{��b���ia$�<���%��mEޞ�%�I�	S������C�����
Ǽ��ќ��Z-]R�zh0��2 ��v[���/)�˳��x�N?/_������i�q�3^�e.;tH?��}���C�YHI_<^J�)�Iӭ��r\3�3� jA���R~1j����{Xq�������:��*DK�fk]ș%g~��8�p%`�
l/�3���6�����3����p� ���1���zO!C1��n�Ͻz<m��#4��l1=�qk��*V��L�|F��3���<�˖ ��^�C�~�����C���/$��-�r�̫P�r�ʛ1��qK(��R2�h��"��(=���o<��D������c�u+�+���à�U�:�Ë�\P�pt0�`�*�;�_�=T�y�3������0����`���l�s��>��C�yj���$#G	�HH��²)��h�+�
|}4��p�[�*�T��ڏ�4�����>n;�^T��0�<b����AjH�oܼ`��+��:�Gq�F!�� _�:|9��� ��ے�L�)D��??H���h&Ν�3���u]"d��LKA��
��/�d�����>�
��:�l.ʰ��yO1���nH��^F?F<��X��	����k8wy��6,;���-Y5eD<��螦U�4���:�v0���������À�4����E�l��"=�A�=���	�C��&��%��]�|m[�`���-��t64�섾�Y��*lK�AuQ�,c���3��C�EM�L/O��t�p|V�#��H[�Gg�7��r�3�b�R��C�������߰�d�������ҿ����³z���h��0$����Tl�����Aˊ���W�/3�*
���(ڋG��T�(z�g�!�h�FQ�_�����7l�{?Q`IXd(ܦ��m2\M������75g�k��jFfKi�Vm{�m�E0G@�u�*0H
/�x��`�ϻ�!��$Τ`+Ѽ贗T
��e�X7TeB�L��h옙����U�	j�R����X{l�,}�I	�����DE�<�J^"� �#g�3���N�G��K�d&1�_&	���,}�B	-K��U��'E�$^�>J�)�\�ޤ�︣�����F������'���n�st����S%���E� 6�I�$\\�7����K���!��c���:�