��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8��A��t��
�]W˱�ӆo �I{�C3槏��ff7 8��6���7�Y)`6�-�7,!�=�f�&Q��"�qiK���ﳑ�ɃnT:��J����""ӜJT��Ʌj����uo��]B1��IJ�P+p���Ү�r���~$̬�͇��!��||�XG�@,U���56=�t�we[�Ax��mԧ3C�d�u!�R�9У�X�c�m<>$y��l]�
�tf�?�� ^��fdT<�n���r��s�?��Z*�����)��Y����:�v���c��0�`X���}m�z0\)	�/O��Q�J�rV�SK���&�v�!n!	�!��z|�M�%.�.�\��R���Y�q��CN�`"$�T���9�w{��˙�������m�![�Xxug�i/�~����ʠ���t�s<<��3�54s<���\0ΗT����a��	�ֿp'���B��l}�H8x�99Y*)�ڔ3Z�S�q����1=UY�.WQT�ڭ��r��m))�	h�Yte{M4�=�#7�|�M)�Ӷ���A{�Hx��� ��r�P��믚;�-�#嚄��0)��+x��	��D�ʨ|ԳP��
_29����-�$�`gS�Ӆ ��9��VA|�7^�F!<&��G߂K"2S��l+r{��X�|`P��ޚ:	�y�U61��{���c��'�:zpFC~��Q�A��ڧ��^�=~������`�1+ҹ4��TbN:��0O�c:(����g�8���y��}��
�3�Aa50�>���q#o����k�@�+gt��,c$�Y�����m����ǃ:f��Z�&�[J������O��t]�;ǘ����vk��A�������h��'xҠ�(�]�������þ���>�a����~kx�ј..E�<w&���3����Z��������x���
��ʨ���P���c.���֡[��%��^��\5Beke;_^2����k���AX���`�&���oA@�M�!�8��dDB�QT���c�߬���To(�e���'��#�*-Bb����<=`r�p��&��7��د��M?�=YM��qU�Ԭ��y�z �]Y��O���� b���/B]%W�嶥���2�Y1	�}5Z�����7^.x����d~��=H�|�K@�COx%ap|W�Y!�Ӵ�Pq�z�!�z�=�B��|s+�ry��'�ߪV�v��*�y�#p�����Ql�\���m�%�c�Vژև��edn&�7b�^'z�\F$ߍ�*��D�<�4�4m:Ӓ��>.�Qr=�B4�V�.�v�"
f�8P����������umNI�{Ӂ���[G#�R���0�jo�t{�
��3��ݍ����-����O�`-GO?C�&z#J����d{$� �lb�F�s�rdA�̠AK��)A�uω�&Ձ�-�1��HcH:h:���=ad�퓇�|�_���니g�k����B6́Vi�%�M�"�����3�k��a�M��d�Ij�w+V��0�W$r���>���l���"�>��꯰��Y��tJ/�WaZU������VhQ�i�7`q��[���׬�B;������x"^�E� �0�?�n-6�I�Z��1cr�7U������LԒ��E�����|��x
Ef��녕�9�ۙH.=�Ĺ�\Kv�q�ܢ��ۤ�i��Ά���L�;�:������1�/+�:��ŧ��R�/޿� |=;���GS�M�!4d�E[F���͍}�˰���G�g`
hH731�m������6�F�QIk(*4C:]�'DH�7]�=E9Th����Ƕ�(��0�s�2�TO&���C�ѝ���G$Z6���y���5�����F�b��������a�Eh���������z����ߙ�7��m������U�ծƸ|٠�y<�A��א���:݉a����%ye���ܫC��:+�P���<>q����p(���{?){���pA�ݝ��W��~��#�`�{1S�H�՛E3�����9��AL�W��{O��WO���'/ɡX�E�A
'�����	Ll�e웭�2C�_�8���������7��I�i�1܎�}�����
�5a"�5E}*�ּ���g��^���_9���|N�MB�c��P���m����ژ��^�>�h�g����L����c��X���g���S�)	�Çn�����M�D�^UR~���)�R�Ȓa�.6�1�5N��{Q �I�x� �o��+�$`(|;Y�\�Z$�+q��� L\hD�n z,�������n|�����K+�-q�����������1�V��w��� -'�J��AhCD'�^�l ��x�d�����:����^� �>=��0��Ň+M� E�X]c�)4jӱ�1V�!
$gvh��*9d�{
�1�LR��AUP��晧�����<j�
�)���T��ۏ/iA����]�jZ:�ȩ�Ǣ�ae����T��mhK���h�j=[ .nx�E<*�b����o�f�������Q������J�:��{9�/~������˵G7 �iS&�@�ha)^�Ŗ4��:U���r<�wK��V����ي)��WF>�e�HC�\v����A6R�Q7�\i��G1�U�zt�I��0q��a0���ޢɨ��G�RWK0U�%C�o�~=��\a�t#�4{��%w��R�Z�wuH\�#U�7�;�x>����+9�O��k��r�-�#D`K� �C�a��:����d��lƗ��q����l2���S�VG����cS�fx�HL9�D�VO�\��b^� ��L�gs,��aW&����WT`�M�D�gP�D����m�nV��h�dY�e�I2_'������$�a`%"m����h$��m#���ҴK�E|eW9�e^�O70����0��n����g��?�$B*��N�K��(� �uaz��N���h�j��i�ع�E_`3V��Փè��\0�����t���*~*e�e���  ��@V��4&�y���ϭL�:���L���_�s����
'�����5��A�'Vv�0 �s\�0�����K<"�B�ٓ�S�[�7]�t��6T�R�Um�r�~O���{�.Z�Sq���,�ͼq1�$��l�J�GBF�D�w�����v�NG R�b	 ���a�*��;���T�,�3���=��(T�逄K`�9q�ؖ���k��xS�M�-[jnz�W����D��;�H �wsŚ,'��I��l�X��X��)n�u�g~ n�t�GJ��]O���Q���vb�k)�Ro�>�;����Ʉ��[�	z��J�.���t�N�2�&̫�ڽ�$+<#s;|�#� aVZ+Q4���N뵵�A����E.�e��POo0�$�m��e���ſ�:�ZrC;=e�f0�Б�i<1@=ãN�?���-B�3�2A5b�YE@!`�mK��%�	?f��%Knn,z���7.9:%�hSR���v!Ɖ,�(�%o'P��zx�� ��[_�����ȑ��m�1G�p?�'{!��>c
t���������nH���L���)�s�fJ,����*z+s���6H]�d�Ps߽�b	YN(�]o�Wc��G�~����T	��MZ%jQv�d+D6�~�)>#���`:�����	�/#��zVKE���e)��:��6���v��y���q9v��X6AB��⚳��DX�[�x��C�#||�̢=Y����%/����o�r��J#1פV5D�E>�o쀣�����ǉ|-�Y��8��+���=�S�<=�#<S���=�����?/0\��I�m��\OC���O� ����A�5%�Rڨ[��E_�8*_~ĔTC�D�!���s�)�0��\����{r�	;��n�l�}�܋f
&!�0��Br$����B<.��I9zܚ��	���6��x�O��@�B�?M��yZ��}�� 3d�گ�i%���:�� ��+f?���DP.��y���lqf)��n5�>�=$��������:>�y�8��n6��e%�T���H����O6@a��U����F���S��8^�Phx��I)�,�$>*<�\�u��ˤ��{��ȅ�q�[S�̭�*��C��U ��o����$HH���p��A��d�v��Ww;�O�dٙ\=u�W��C ��<�\�}� [t0��ZР5��e�����ӊ;U-$�{�7�0�Z���H����%B�Hn�6��|�Y/���ޑ�ǅI*��䴝�9�f"��W�"ٮ�9 ���֙��zm��^�&�{o��D[�C�,�,���f����iF�*1Y?��-1�0�OF�9�G�vg%�w��_-�=Z�H�\y���.5x��`L�L6���A�?� mN���c'�Bf�w0hj������T��TΉ"y�:���lu��o$M˖\Qx�a0aU���)$)���(i��9�O����$RM�zŰv�W�{�ȝ�H��Rkt�6�V ��n��9���A�w_�lŃ"}���[Ѩ����VDF���=���Uꢺb�:
'�ꡭq���i=�ϙ	콌�/N��o�Q�^q��O��l�V�mEB^wk��6AUپ�i�@Ȧ�A��ة8�X�����Rg�����S��v;�G��������W�������o��W��E���?�+����4f`�O�d�L�>��r�Ok���_�mfE�G���M1��p��"�ڮ��V�����5�x�<an�����*��"R `�]tZD2��W{(�M:[k~�Qh#�������:&��y���l8���*�ޥ�@$,��������!nc7�l�H]��_t����Qq+�R6�눩! Q�3/]��bIvq�>�ٲq���
��9{�����SWQ\�{�'��iv���X���]�\�趖D�{�
��#,�).��ʾ
Y�A,д��L㥔E��	�g%�0����u�<�N�8��7��	�M�sed��06�5��=��&%C�0�G����so��ji ��brg��1�@|7]ym���C�/#BLY�
+K*8#�;$(ؚ���Dpb�'��%{?�`���?�ߦ�d�_!0cM*�FV^�!�}���)�p��޾3p���(=H��>d��a�A%���Ԯ�Ӆ'�[Ρ1=n�~+r����:��g��+�9$7�7n����&�/l��e���Up�ې��b��&'�� {��K��*t6��PK�I�Z&�U9MT���i��<w��K|�(%�O��ch伄����,�VKO���=p���]�T{4P`��{�'o�)�`'-*0�$��5����:m�Ofq6�ږ%; I<7JH=�j7.�&n��������)��P���}rk�§��nTQ��#�u&^󬎡����</=uG��Vv$��	x����Bt09�٧NAل�zMjy�/�އ�Q��T�id}�GxF�_���!��!�z���%k[Z�E7m!��kVv�c16��VjY��?�tVɝ��	�;�i�G��y����HF���>���[��,���X��fd�1t�~s�kd�P���f)�_1���ZJ5�}�a�����!𥌩��=��<�'#�v��d�T4@�����Y�|��l^��g�\�<�ß Ep�˹�͙Q�D��f�^8uq�ۧ��� 	�
I-��/��w heA�U�`�����R��I�(Ik�D�D�kVƶX�#zbN��XW+�X%)苄'�άUi�.Fk6l�c���4Ih�4���U��cxYփ�7���� �݉�������)���<�O	����0AϚ��� M�ќ�'��a�����'��<Hkg��$-���]ʠ���h���"CS�)�C��i��R��d�"n%|oL�����
j���Bo���At�7�#	�Z�ON'�Y#����O0�,K���0�o8�T�¿"��2��ǽEK��'���l�"�K@v���@F�Զ���O�`+2���"�a,^�C���a�_�w��;V)�k)�I��m$�{�'��\l���979���Y�!#����7�-��Fq��?���L�b�4f��:�Ω0��R�V<������Kn'; ���������lH��B��MҘ>����|�&������x��Y��7K����\�AҦ�>F��Jt��Է+�Sp֭�$�Q�:�x���Ϡn��B��nQ6F�J`���lǲ��4����s/�CBF0�qdb븻��`����k���:�F�l}��������[D-y�R%��k�G����&�7�eNLu-t�I��\���w�x�-j� �yL@��S+e�w>��_#@�jꐗ~sq=N٫��Q�����hh;P�m�I]�*B܉���)�QF6�!�Z07�rc,j�9�1�r�J�8׾:tn�-�v
j�B�dA3&�]!L��ѵIlL��У��eK�ߨps��'#ô��)�
����Tc�lN%u=.�U�"-�"����EU)I�F�@���c�{�?t�%X�3����� ��q	�ͻ�t<���~^��B:L
I�Ԓ5�(N[��t��f:.eNd�w�c7�O�rv�X��ʮQ���e��bt�TBEH|fu;�E�N�'VYpC���M܀B-���I�^ؗr��&�t]v�<��,����Q*c�������
�����*S�ʬ[hް4\���>�u���{�K�Rc*k���N�$�@��Q�q�  ����SO�����s��6��
�5z���T���^����(_���݄�?��h�ikԇt�u�t��G�K'L�v��NRf�*��|u)-��;��-����Ȣ��Z�EFAn4%���&^B�r�D�����9�A$`i�C.EO��i���c�>g$@��nZ�ju�e	��m.[�D�C��(c�:���'ݜ&4a���P�������'泇��� L���%�p�&f�?</ݨt\�Q�G�������Ĩǀ��L2Eg��-ۃ8�������������s��(�K��#�'^�5������@��f*y��(E�D�5��!έG�P��g��)�T�u�; �\�Bu��)�����h���i����X��>��4��R�CA/,�e栬����F��B��m`6�oKܭ{Ƙ0EGg®p`���l��yK��c��=e�~�&����O��B�ی�J|��Ǆ]؈����3�FT�,�{��縥�#����(s;� �l��Y�G���_V='���;K֋؃OA��99�>Tj�K���	q8?�ޗi��j���'m�{]��uQ{t���8���>0��<&��S���C0E	���q���%$ Y�5^�m.,������T�>�'�|%]�ȭV]��aX�B��^�7��ī~V1�g7�o¤Kg,�|.l5m�3u%�|bp��=�	M�{(`�ږ���\�7�R�BŪ��,4u��aY�~{�����6�}�y'T�q��B���C,�d�9���h�k��#��_�N[)(��,��"M���W��a�j
S�������&W��N:�:i(W9��l�N��=/r,9�?�CTN��sT�_�`f�r�%�{�hc�+)^���*�H�V�q\�OӨ���I��>����t R����* ��s����w<��� 5�ɸP�����~�vaO��C�\?'.(�Q���b��Rx�T��N6��X|t��a��h;*��V�9m6B4c4����v�ۙ׍�V�9�����̠��a.f>�hB�CN�uĢ��^s��9*i��1�(�%<�N�f�4Xp��b�ˇ����eD
06<�_�{�(2��S���&h��'� yf��a��Q���)��� �]��=����A��h7?kRw�)hX&�.2*��o(A,1+�v��]��24xr�~�s��j(���PP+LB�Z�h'���9����Ujv5�אC)�����WXG�bP��ى[Z2䩣pi�ڈõ�0]u4�h�,/`to, x���n8�62�t�]5&>���Vc��n��Ҭ��k{n��g���u�L�v��T�Eߢ�\ ;�S��!�ἷ�����v[?	���V�͆��^�-rF�m찈c���,U�g��FC��;�L���z���Bl�E9��/�F�� P�/;�I<T�rCJ�3r�f������C��I8�f��T�A�%��
�>����;�|���(e��=�x�q쭛Ϡ���gw���<:^�؟j��eޯ�Ptu�`]O��[y8�]�n��N��{ �Ņ��ܨ�e%5Twܫ�;�
�7j���8���,���;6J8�S
�2��t3�P��`�����Q|��qC|M#�¿��vth�YW����s�GG7�����|�T6��_�?��9Con�፨\_���?9!̣4���x��$���<�E��)���e�k��>B�V5$T��\P�Ph�%Qv��{�'�`[�R!_��1��+���F0i{�oU'�6?����>�Fs�t�E�1ZVk����(E�o�p�Ϣ$)Bm��!���7�U0�u10a�-�&���h�%a�wj���Y�z���8S���1�b*)�C�7�I�oǠf8�u�e��Mq�0o,�J����oqpz+����p�P�w,�M��\%�;F��I�����Wii;�dkW� �����癝s����Ժ<評L����&�il��C��w�N=��`�����'���E���|�Z��_7�5�*F
YD��t:��zp���;�7�P���ۺ$G ��VM7�(ZaHO�X��۸;p��#�͎Z�^ڝ��WP<L�Ȑ6��i��zj����(�7�u�kv�;y�ݑ���t
�XO�F>�����~�N���,R�5?�]������D�3ʖì<x�R�Li+��wM*ㄗ�Q�t#�I�!� ��\��,�q.�哓��$�̖���gmo��E?�}��ӈd��e��xږ
�[�@U�D�r�l�-#������9c�����4^�65C�c(���4��P*������/+b���s���c�gD��n1�@LE�X�MP�0.�]�k�yt
��x�=.�1�O��U�_˷9���Ww;���ŗ�3v��*�݇+L��>y����qC�m����7��i�����f&�'§'	?@ӛ�w/��}���� ⮬�p��Vm:�%��_�{޻��vP�Y���qe�-/*�B�?*5��]j��K	�0�=�E�E���ND{��/H���X��8��f>p�s����,x5
�{���h��*� ��"7�=22�.	�*#���N/��N��Z݅�^t�vZl��z���U7_�u'���~���l�C���$Pq ��kөt�h�Bww����N�^�a�ݟ�����)5�4殓4���4tok�Q��b0ql�C��*�~���骧�j~Pc!/@�J�<�T�#J.�uX ��k��i����r��z!�Ww}
��s�<.fS�U}1��/����m��"IDs�99���%q��u��Np_INa7j�J ��O#T,H��f�:e�ȟ�?��i�+Y$���Pʸt�\89���_8���'���WrZ(;�<fU���W������D��c1hH<�-��/_���:,��4(	љG�A��n#D.�r��C�������'M��o�Zm2�Pz4�������m���ʸ�mS�[�.��
�C�5X_��#����UX���`S�3��I\�V;@5� V|�F�X�(�7����8|o�fI;@k��&L�I����+��;��k��ğ��rW��N1�$/>��^,��,n����2{�c7��M�U�aQ"m�:�$��b���he���,���� �v��Cр���擺�O�52���ͫ��x��@ޥmsdE~�;=HL�׾7g�d�ۂ��ޗO�ʔ'���c46NԮEj�����*SfC:-+F�|�		D� 2�v�i�Q��!ɮ�iJ4�W>������ɼ�^��:�/"�I��"�H�|ځ{��S��}ӄj��$��ȥ1�Y�L�ō�{:
�E�2�"%М2p�L^��8	������	�!����H�:[e _q��F�	���lw�!f��mQ.�w0���
��ޝ��F�{����x�R)&	c�
<�F,{{fۣ�橚+�z�@����N�&���
���
f�
.f�S ��2�-�s*��M�a���S�<��P��}M�z ��KS��E��QS�;��ċs�2���[������;oD��c�:tǥ}���v<�(y榋�e�2Ȓi��v���l1'�=/?Q7j��P��?�����LJǋǁ��v9�SCŏ�WE҆O\/da"G%)\���E�t����Ý3< �,>:��lnJ�Iv��Rkm�7.�˜�H��E��Y��ko,OZ��eܱ'�[�$��<��Ed�c�;��#��~WL���i��#�[¶k<̰(�� !c���i��>+�A1X<�#�Г�VS��z��{��9��N�Dt���%Z9Z���m�C�r9s�;C�#[Mt試TuE�B�&�t2�'C�u�H�S����"Y�:ӂ���8~ݴ'��,��XD���pnI�ϭES+r3��Ś���f�Au�Gu��/tL���&�!Ǭ�*#�,?�q��Ҋ�ý��w6@{ ,|���"�p��p���ӏ�&��ŕ�����7�G�R��Xh�4��Ό�+��߇-���2�m���u�j�r04�(�wj�,��w�Sօ���ذ�*-�}u�w�Q0�6~�����n�x?�B��?3����9c�ǨPI+�?�����1�f��aH�����NyF4������5ڜȮ:��g��R�U$;F���d�nG!	��e��?4��=�k��;�l :5�&�����	����'vH{ME"� \ \� xR4��y�DX��튷���xm�ډ�k�F ��z5!}1�"�ח�Â� ��ڳ2�%�Tf��^����{�#!3�dq�W��mv��������?,���"�9��]�����*�c�2��+� C�1A
��Y������.[�F��c_/�ވ�������_�|�ȉ*���A�(�´M��C=��d	��i�V%xM\+Qu,���d�.�s�+ͳ[�Hs�"�Sv�lg�q,/!��r����=B꺀E�XG�m�2`5w�Ugju�B�=��.�F��vI`s�y�nd��d���IǓ�dm��=[�,7�����X��.
�-�J->ݤ/�hkO��p����$��m�g�v���Ģ��jMgќ,�'S�A���N��C�?HMr�G������?�j����ǲ�Kr����2�ގ�m��u�5/k��7`?aפ�	�	�����E�.e�pÊ�a\��)u�������(�Y�s%�B��X����`���l�e�=Ʊ��mi�;qD1��{��EcZ���&ِ4��C-�����G)�f.��R=�Ҟ��n�r��}�J!�cY��3D|�������F��Aj�)�f�	���1���ī�tO�}E����.�F�����3��o�)(!:�֬U+"7J0߅M<e�@X����(���W�i���]��J��!�iBNϘ����C$���f��S�϶@��f�rr�'�:�9'\�	�����3�ƕ�1��L�KW�ƚہ,_���ꔧmzD|P՟$�������6�ɼ��.�PZ~�G��8�;�,\�(V�c�̄�)Z.G� M��6����{�`���PB?!��1����{,i8d���j���C� ��۵�;�d*��UQ��:�	hZw�	cOt:���H�<Ȉ���I=|��Z\�n��ZU=�N�tcŵ/�H\�&%�� �����R1����>��[�h�ls�S2�k����L��ۯ�cN���G��J�?\&/�m�X�ܤ�uݩH�P&��p~���V��Ad[�	�ͧ��
7�����2�wF��w�fk��H��[c��G�R�7`݁ �]a��p�����Ts��_/;	f_���j��2�y�� \�_C�Xd5�����Lc `�  O��=�U���83�g���j��R[����t]���t��&GU���;��U�C~��u����b�&RC��!�%�b������D	��S�����$V>�UvU;zi`�Cn;�"7ʃ>�����
�/��(b���#���X����[��x�ࣻ��8zN�}�n6(��%����P���_�k�Â���DM���kvn9�eF=�}�K#���BWݜ�����-�K J�0%(�v>Y?�7�hz=]}sm��4L���7nʬV��T�����h��h���e~�&���Z�D�����1)������n96�������na!;\����s�,��eRAP �(x&����RVo�P`֧Z�%ޛ�:�\���K�ע�&��m�Щ�P�:-��G遠@SN�u�9xe���@�o|�~\����!���7<x���z�O�;���ң�&Xqg�g��e��J��7�w�j7KU-���2$w5}"�!�e�����x�
Xq��)�|�M7��;�=/��R��#s/�������B�o5��ϧA��~�5��/��'�设qZ#֫�6_�7k0(�*fѸJ/���kDKd�}�t�3�(D�ʆq���7Wب��}�-P�Ġ(����߳W��z &�t��D}��	����X�A;H�M�6-�X]lf8��>6�!�
\��D̠��׷�1M+j�zF
�5=E`�����ښɿ�~wq�K[U���vw����utg��H��C���i<����0E��X�a�Ӎ�';�h���M��B����/N?��~4��`@P�	������q�3Q�?���&�_��y��(	��<+��f���Q������$�t�O��}���,��d5��-����Lp����8jk�{�FL���k�RJ�N�Ƒqʸ	��ۅ�������A���i �#�i<�(dY�wg���/�ͳ�ya���J��K������X�*�Z�%%_1P}�>�z[���P�Λ�Qd�I>�.��ـ:K��@�,#Ǡ����o�5���v�]���K$��.�X :��8@G���h��8���_�G��X��+��]F�*�=03�-��5U�CQ�ǔ���
G�G%�*杙��/�yS�e�^�{(�p����(���m�d��U��χ6�bl|�cɲn��)%�y���U�aF0P���;��;ѴIz�,(P_�0�<~ܟ���v�M�i.`I5AӫB�3��{�z��ˣ��9;Y~#U�!�w��΋Dq�h\��85ic�n��t��b�RQ���S�v9xIמ��NZ�5pJ$��!/#��-y鞧C�P.�"�L���h�.�����g��*�,�$��n���fz)����ޭGU�~���#�1���XeC�����^�$�u#5#�/�TE�yK�5@:�<.V?G�����-��g��:���V�9l�g�^rZH���=E\����H����\y%�	t����j�ᴟ�䗣�1ǫgN�e���w!�{��w��ป�|�����~9�g����啣�KN����!�ގ�~��ʴS��֍��F����M�ϼj�
G&>!G��Q�2l~)�������W��g�ఎ�����e=w�����{�8D"��AMJ�� �sx���eǂ�ص��Wv�䭤���j��S�=S��/A�����z�\�g�-�����g4g��C��+Lg4a� �A��#F���Gj�Q��1�$������){c���]U2>8��:����kh[��	/y�
��B�)�F.�ȴ��1	��)�7^w�*9I
�S<�F+�C�0e�|#H��B:����,�|��`����֌�XX4����r���wI#;�Խ)�Q�<u�3�6��[[Kn�'���ѱ��#�xG�nԢ�[֢/3\9*�Nf^*�؅���șo����(v��'�M���7���o���߬%��Ug޹B֬758��r|_})�R�p�벻�������@�᫦c�qF��9���F���<�?T���x������X�\�������H�.4��R��w ���[��c��=?vI��|�Ο��4B-s��-��#�	�d:w����|;���U�,6	_����E~��hi��E>0b�̝�תg�@9�f����싄���"��x�\Ω	d���{�LQ� u