��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�X)�='�L�.|�w1h����ȆwE4��f�����(�p��4\ ���1�Mmm�Nu�=���s��)�ڢϼ��xJG;i)�	X0\� �}�KY�����?5=]���9��|h�Ӫp�b�/8�I��&$[�n�R����_ F;���5N�����&�
��B��ۜ� S�������w����M{П�I@h�0���E0uW*�~"��\���h���:a���c%->w�C[����_J�Yі�j���)T�;���p��A����SJ�CЪ�Ģ4Y�f4���8L��esY��[I.��v��Y	´��(��]�Pcۿ���$E�y�,7���o$7���3�	B	׾V�k�����3�eU��$u��Q�ǒ���̢�:�IH�>���S�E�����BiT��>l���>R�Q�s^��N������[F����$�l�?��[����[|Y���o/�">�\�^� KVslq�~3�O���(�����\�A�4�{�(\I��qc�7��K+*~`M���b���f�#,jS`?Bԟ��q�h����PǊ9��L+�]Q�G�D�^p�6��KI�>��%!�1�"��J�R2��7���Z6���ɓ�Hi�g�cL�ꌘ�+��?�K�� $�%���L\�k+՟��Z����e���O2M�a:e:�'/)»��˳���M ��}�?I~��BWoI�R��$ǲ��z��4�����Ɋ���t�Ń:�3�� �h]�H��"�7��3�\�}5��@���3��W9��oPR�o�$��m<��+N���|
�jߒ�CM���p�3N��D��ˈaK����iЯ�f7��<�u���D=���?�B. 'DU�����o��C9�UF�%�w�4s$�B:��0��$hՇ�FZ�!��1�g,�@�B�?p��JW��sQ��y6d��BU��ȁM@־4�x�6 R6�A��#.V0�+�����-�P�8����c�:��"���e��������,b��X#l��Vt��4��*Yl�k����
� �d��miD]L��\�D0+��3�Z���f�Gj,��[h�:�^4�����pt�ԫz녺�w�h��@��{$)V=��J��ߕ//�3��,(�R�,��Ut�J��+U��A!����hH���dI�H��F	�KPD�����;�BW��4_S���0$����z��j��`�fl�� u�(X�s�V�uTn�C�Q�1��X���_��d�_Ie��98�q�c;y�s�e��7�5�'4�A�7�%�1��❣H+�j@�ET�T�Ô��(�u�ǈ��K<�U�MKv���aD�f�WH���br��b���o�7׌P�~*�9��4ϻ�H�f�&xg?�)U�C$്���%���(��h#�� {�M�h��y�#
�����?#P3�󴽇q����<t���-�N4�-3,vM�t�(��Il���6׼?�(�{�r�	;]`�<
�_CQh t�/�IQ/|j��lZVc���'�w�T��h���dLQ������a�����O�����UU�7*��ę��kZ���ۙk)ٰvx-���Cjl�ݡ~�.3���;��wB� ���ҥ���F��u1�T`��1�O�w��'��p�"����#�9�@P�w2~]���U1�F^y����P23��J�{���?���C��(x.
rx���T�՞����TU�`���Z�9�ʵ;���-�I�V���U�jJ-j�b����7D�R�®^�W��[�`s�q��3��zg��	�_���S���#���n��՝���Y��,2a���1kN��\ay=���n�=�5&����D�ĎB���X�����D�G���2����6� �"�v`4͹�ݾ�^m[��y���	�����![�i_�'#��4���+O�e�3+7�,|{��ҙ��G���6�b�x�'�ې�������_85U�dl���*u��A��>��hi��ٓB���y�ޛM�[8;���t�	E����A����LO����`0����$�G]o����H�َ�VM�z�)�0�e�T��;��J#��^f��ܛϧ�m]�L��SW���k�'Pt�+�z��k�m���\Bd��_V"L8�kʦ~.:��1bJ�b!�t Jc��u��k��&m�@���Kʨ��)_Ᵹ��K�{~*;�$L?����ظw�Ac���yൈ�DT��s[��Vn�S�*K�^sJ�h����oz&���h�4y,�|��H�e�
An?�lN�_,��]
�k<�Ӻ����Oz�y�|�x��HC���7W�0�{Y�O��Z��Z_=���G�?�Ϋ�p��__���Q�,��ry��PKd
V9���G���5?"�1���PX�?��>��"	쾙v����y�''����6.���uk:
;.�6K_����s��+��B���H����Y:.t����V���h����x�K/�K���.0ƃC6��ΐh�Gþt�2�Lz^��+�!'��4#�]y޼ݖ��+#;{��2���[�\�!��v����u�`3�n0���*h;��z��wX�¡��)������#x�Y�&�F;�i�~�!ϦS���NY6�Z��>��-�c�Ү���%�K�rl�������`�}T���/1���00�Pq�����K'�Д���G�t�{��~��ؗ3r�X��:���'�c��� �ޖ3��ϑ3�ob�T�mNi��5G�M����\��q��^:m���.��44b��G�	���&pKL��m�^�s�������{r��TR�l|T�h�ۣ�iD�!���KK�#�D߸�����Ů�t�Ol�G
����BSeN���JgW%xvl���f���%'Ra[t�iW��3����T�տ�<,������\�G��+>-�iF�W��n�=�#��q��E�Ͱ�XM��q�e����c�Rz���c&u�5	��Е"r�z��ʦ.s�Iu�a�w�b�|��C�N�X�t��/����h���`�h9C�A�lʅ��JRYy@X\�՗S<�b̒�H�G�T�ҋ��bT�WZ��x�3T�8�Q��n��Ն�s(�h��8=}�&7c�@�4�״_RQ��I��'��~�l���͢����^�yJ�  ��9����o�hx�|,��҈]?�I|�x�Nw�_��ԉ<ݗ�=viTF�bh�-�ez� �LL��|��ɝ�����ݍÜ����`�����B�59�I����G[A����סØ�{n(�W���S����$�P�t�2��A��G�`���@d�S�v5��