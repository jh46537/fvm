��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�H|��6	x��:Rg�J`>�gPnLG��Y4d��R?�¾
�p��8ϺX���a��D����*��C�*�x������N�OF3RY����q~>s�-wjj��x�LıۨN;�_OV�3'8/�O���"W�ЙU5&H7iRN|ߪ��ϑ\ ϯ3'�� Q�9��o��� @H�jHa�)[h�W%3��4ީ��ī���&`Wʧ36N�/�����2-�$�X�_m����O�yV�ܙ�̋���/"�Hzxd���ɳ9%�}>�� �E�RM�@1��f��.r!�awPp������$� u��3��v���r�!����s�P��N_w�^�+��Ӏ�pQ����8��]�g�qӢ���	<%0��;��v|�6���a���-��l����ÿ�Y�;�0݇qEح��q��bҁLQc�f�YҾ��T!��Sf���Y���<�eI��:{��-ދG���Jȼ��2=��:Rh���z���o`�FN΋2p[���OH�����2����א�>K�vu�b�9"��K��^Cb�@	��F�/�� �t����\��}���duk��(�}��Ȫ����q��_\E^��@�Q��C�xt/��l��6�1}ª�e��[�Ì+��E&���<�����Jqrz�f�@�(�e����"<��:����A켩��1+�50�7�/��F��@��o�[ih�E_�g����t��}�OL�;�"��W}5��"���<��.٢D�Ւ�Rn_J=b�SER$��ErN&a!ݧ��z��v�QGC�W�۱L@ |�ȅu\��
��ݜ�J��P_R��l����'�gpW8���Z��)US��<We�1Q�9jJ!y^��:�����֩[���O�4��2,���'�Re�N�;+�[j#ÖS櫣[�6���9N$�#�]S�ڸ���\���M"��e:�[^�|�'bt��	�P��	��XW2�g��+���bX���1���z�4t�\u�o&d�ʼPj(�a	ln�?��*�k໸M���Ы������G���L���i���^����\��a�Z�}S0�����wQ�T�Emq�K`�+s��&�9B�fo%��FQV�U�`0*�{|� @���hA_��)��[��{G���!i���ߨ�m�ڰ{י'#���r4 ʿ ��W�孊�ɣ�/q9Ћ�U�i�٬R+��R�~�a�v�uRW
O?}����A-���=0��	gJN�M>U�4^������h�UX�U�݁SQ)�s�/GG�cj@�����$hlA��
�^oj�#��~�E�)�Pf	�ED����`�{���-k-`��C]��O�����|���K�Zs�� �����_c/�&Ki��Y4"�x�\K�M�i�K�m��h� T��o��NJ�)t�~�z#�o`�E�q[1�n5��D�����(R��E���U+=rN�l1l�P%f34�镑�1"1_�j�r�����c�iG�m��{��ȥL�s$�ց�7�n��)���/��)�X�'���5��W���;����t��W�ƀ¯�#�\�G+�=��"":p�w#��IF!Ӵ�#��Ӻ�����~E�� u-�3#�_���>ś��x�]���O�L�V�dG�=ZQ����:��X���:y/Î��~?��q�@�ƛp�Kfx�-��ZV�F�T?y�R����$o���(N��
�V�Ѽ�/���@�|��	4gWĳ��?��%�kV����ǜ/>�"B�Z y�ցy�;�)�\��Tk����Ρ��!Q��������%�:�F�ZҦ��v�����4#si���s�	��8J/����6MђVS�i���z�㎎rK��R����\f)���~ ����dT|l5I��O��w������r�K>?����2��WӦp�� ��2O�a�f� ��;>1�/�d$	0f�h���0��i�Ѥ^�����w���w���=Dͭ�!~+S���i@S�,�y4�a�����o������@�>>�w�ӊ�at|���~�K��fw�Ka��H�h�	8i�EX��������������^e	��`R}Z�*�O��.g����,7�mW� ?�?иt�� ��b�P$N��
7�c~Ԇ�})�v�܁Z��t<v?�