��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""���᤬����[���%r���dY;�uU^	/���D�B/9����t�.0��	�#���ѭ��aj���0��<Cݤ�2t�Q#)�%�^\�<�?\�l�j�� u�c�"��>�G����7i���z=�s����̏���VK5(?��؋�Z˨��<)�~��Ϻ�"�y
�º�/�%>iI��vj��?��9t��7l�����A�sG@ϐ��i0�AR�C�N2񢄋$���~��g6��K���7AÒ!��Z���r)�˨�E��DK�G	��MԺk�V�2ֈ���x�2��=M�]:{�޵�s
��"�|x�8�;����d�|�6��{�범iw��
�a�9�	�0m?v���L9O��>���h�)A���TJ �w�}������oƽ���3��A �uϕ�ɻa;~�_T#kRׁ�&��M����}���vuS���x�8[*+�9t��(H՗���.�����L~*����>籦e#�|�Nߖv��-@X��o�����	;��v`8�	��PKTu�Ms�l�p}�Z�VIh�c�k3��A�~�z>"�^FT��ӹ�� �����妅����{VGa��z�xDB��)/��������[�8��՞\M�`d��4�}Dd�z�|� O�ƀ��״g3j��8�~�yF��׶��0Uݱ�1c�[�u/��; �<�%�&jft��?7��p��bQ�T�ts0�I&5k�zޝ���A�q�H�����]u
U�[�Ո��w������K��Ǖ.��f����G5 z��S�^�j�/Z�r��b�ѓi�if��+��XӐJ8�aU+U���,YaՅ����Ɂ���aP���G�"8���jU�j7�#�v�)��m���Y���@�y�s�Wr�ĸ�B���X�]v@gs���| �
'V�O�	&چ��>���Z\5h_���q��0T����Z���]��x ���T�q�6���DWYȕ�&4��d�e�K��s}��Aj�',��:2x�m)�+�����@�z2�+I���2%s��M�z2�@�\`�3�S�$6+%�>�{�H/iN߻�E�Xl3�Ae|�(׊���P7qm=%�_w��β��zd��3��;�WՈ)�7�/�l{o� n"$ ���=�9�U��F��+�FF��G߮};%��*�0Զ�:@�5���d����g��z(ft���	Bw���71iTei�>����,��4��e����:��0S#4!H���X�"T�_�X���Q�
�)|�p�+�¶qXN����Ԙ3 fH����,�H�\���^D������ˡ�r�M`�1Cg
�*�L�Q��ڣ��Rj��)js��"D�<�f~<qzJP.g����5K��Ru��qu�QjbF� ���s�t&��ǔ�=έ�b�"�C���V"0qǷ�؂$B&VZ+�U�6D�����!WeA2MC�,>^�����gcu��h?e{�Do6'�9γE��t�x���~�����ȧ"������kP���Z��CA[oQ,G���
᫵yn�����L�ц�zGm�T7+��~qH׷��]Y�G�5�u�>�Q��nJo�n?�Y$O���qT0�,2�ZMW<����p����%v��­�$:�6���k�;�K��±�m\�]�<�!�熠r��l]�?�Ypޜ�v!�2؂��:+�y���r�� 6����慖���CI%v�"��Ȩ��'o�9�K�����7�@���o�.��2�{�������q���>��'Y��8b�?#IjB����G��up�	�y�^N�`�����'�r�N�����=��tm%��2?��vP�b��4/��$T�	j���+~�ڎ�	K�������&Ri7��L�n�n\J\܏���r-Y�B�-� �kn����y'�W��4J{���5�)C:�苅���SA����Jx���4��a8�i�VRT�k�	4�;�97�c�bؾ��ƑG&�;7R�ߨtbU��G
$�����h�Ay)�l���#m�s5�p�����O��:�zi�W��g�
d��	~r�6�V����;��T0��ZM8M�;Ӫ���/!�ǁ�xm��k�q���__`]C��x~���z�/_MQu끤R���J���lS�0�Wh�o�\�]�>�=MP4�5�����(Z��f���P�[=��P��G.�36ʰL�)�sg�q*v}J��oƣ5lwVt�	ju8�4��Tm�%h�L-�puxᤆ��"�X$є���� ʟ��̵I��T�̵��*`Q�]��*s�|�L���}�
�1�>ךf�}�1g�J��10~(!��l��g�:�*�ˣJb��J���߰{1@k�������žX��5��	�mDIY�̵�gG�m�&9��Y&ۀ�e���U1H�����>���aD�DA�+��{���w����j4͂���p�uE�w��S��^=8�T�+Cb@�z�t�_=��<���KK���~q1��z���;�"2���|�FqW����/umi=���=zg�3�kcD��� �������@�n�ֳ@"�=C�� k�*+�υ:`�&�%ٸ
T6*,��
H��"o����?��G�^�Ā�D���{ɨ�6�Zg�@�9��Bi*3H³�`���u��
ՕA�6���89�ܯ���:�g!�'�m��hi�Z�'�k���+�J�y��@������_���Tp�#Ң6$��R��O�-�!B����E��Nd�r�/	?_�P�]3<�F.�ӵ�/P	&�MǇ� �9���I/z�Wyk~�d{�9SJg�f�M�>GhAju��s\w�+�{U%������LT��1j����m�u�[I��s�O�*�\��ɕ�|U��0_)ʝg4�i�t](���Y����0���0HNH��m��L)[�3h��NL���U�{R� ��Ћ+m�X�[;��q�ڇ�{_a��b��o�5��RT�9Ueq�/$�:%d�	� a�o!�4��K��
�%b�y�����7h3��I�C�噄M��'+�z�q���+�]2�tx|xl,�#½�~�����ZWP�s�:?��ԙ��ʛ%���-\�C:\��w�[,��n�"���꿒lJب�S-t���K��!ȶk*t��X��s���?Ǎ��ͻsH,�'s?M�6��5ꦿL���})9Q��1K!E|���������"�Y����(m�����:�T(J�0ղ���wVY���L�����	ʹ�*s1��N�%!���w����M���?�'���L�K�q�u&�Cä�=XҨ�h���yd;5p�硩����2Gb��8���lk+/1�"�܉d<X~e�&�6��*7
߈E.ծ��~M'8�n��y�:�.��A��G�GS?��`����	�p�s����,���fZRIןO�`���N�&��H�`}'ot��mv2&�M"����ً��<�GȀ;�HHWPT}����Q6�!�h˶�]��n����������<��O4|{^�����ϴ�>Jw��)�Jy�� W(Z������0�y)�sn�I[��=�M���n���"¤\,��fh����Y�<J,T4wr���W�~L�lHn�w�"�gD6�X�Xe����v@��𳣷�R1j��u9ش�ǉ	�'Z�[������%���ݵ�A�E%�T%)ƴ��s�Y�׮U��}���:[����G >�@���a�x#f��A���9q�Ռ�X����:����}��ԲO�~��MM�؜���M��(���f�Î�04)]�D����>������8��!���w)���3]�g3RJ8H_y��{���`���PY�F�A�_�3WЄS��2v|� ���'WL�A�n�k�ԏAL��[>�3�W���d�*���L�l�_�Oؾ���@Y Wd0�咘�,ƛ�+9a�O�Ow�@�u���D�	-N��?6�c�z�V�fw�'=�x�J���[�)�/qa~5 t� ��!|+��/�>jB��j2��g1E�r�� O��g,��f�c���L�P E�Vbm:��Azh���1f�,e���\j-��R�N,ҧ�Dk����:�r�������VcE�I}(]�J��*J��U��������cs�D-��&�+�Bt���L~f-k��������2I��<L���у�ؼ�s���K:��v�E��?� +��>҇��nnPg}�p��� ��!�C�:�Vlq�hI	6n��#�����٪p򂇸	٩�uo��.@D�;�2��ּ��h(�LMvO�$t�5�}�<Tԭ�iKh^X"c��\n��\���F �ˌ����3U��s=F�P����Rca��n���^���σ>�v��:)R��4��*����{��)3e�=EDG����Ӵ�F����m�#^�|�9k�$s�����:.�?�*��ܷ�70!��0ʲ�2S�B�熁�6��!��	���Wz\fv�F��dz��VPm
�XYN���Y��"�K��̮��~_�fy3u�?5Bֱ:�<#����a2������s����b7�:i>���9�M��tw����F��p [y��k�=�і9xnRֱz�E��Q�;��=&��w�ݢ������@��zM���0ѰD��r�aR�4�gc�C���x�7�õ�Z�3~'�&����V�����P"ٓZ�0C?��4jf�&�.j~\�K.�Co���ES�����Έ��E����sH��h����@(O7��/���T�=���OW�A� g�_�b�Ӿ� �Ŷ�)�)��8�ls��>��D���<o����ѫ8�u���O/�T�3�c�So�y��\�������QϖF�Ǳ��)��(o<����`�(�噩E�s���q��iR�������y��Ū�}ݍU%t�S�^ؑ����o��$L��7���F��<�h�iz��Fgz�-W�o����@�p��a��E�� @��0w�~���	IP������d�o�iJٶz��|�5�֣��k!��8K��̔$	�-�IWw����<_U�B��؛K����I��V9DAk�@ n��E���kA¡b�%�K7 ��5J���WbOd�oD��M���B�30;��=�㱗�8h�h9dr�)1i?���Q~ޥ�G���������M	���A����\�5�wbpiH$�ɜ�0��1����,��<^@ލ��4l���s���W/Z�	���C~�&̠��!�
�A��J1M�Qm2y�7�#>�\�P����<�v7,�0oK�?q=�q{Ԏ��|2��Ԓ�'����x>|S�6Q�T���p�} ·Yl����?���E������h}�u�@��g��g�쿏[�4�t�K\�Λ��3V O��m��K��*���F9�zW��0�]ܗڨ}MS�ċ��O%�B'wx��l� ��o��٢8ЕI��>11b�-w6G��>�=n�
�����E�t}s�S�J6�_&��H����I�}��+�򱻛+�(�zh%v���ZѸ�7|C�D#�:��|!�!� W_�?��}l��6����Y�}��sӭ�Yj���g�E[����A�d���̰�! ��b�M����&�HV���$�>)�:�@j��/�����ez�8⥷j�k
\ٔ�B��+�W��']��NO�&Q�VÉJ6��TXGdz-9�UBN�q"�o��Pd�	W��$��T �L��+x��/� >�Ϙaݺ��Nn�h����Tn��@���X���kி����r�zU3���i�mUK���,�bY�x~�M �f�C��d����c`u�l�8_�.�dr�zx$�A�5H�`�����]�_@���!�@ή6��	�n�=�����(:^����4�6>���m���]���|0����e��*ȍx�Eq����C�����<w�n�
����W�Hm��ƇYPM��(��#�71I@�q����k�G�7{P2z�E�,hz39̑4�		�q�<���^%��ô�]I<%z�;3������E�9}$��S<�q�8�&m��"�{MkJ��Z�i����f(y�����Z��F"�-�q��c"�h�Zi
,3�e����%O��Hǒ�溋�-yO��7&=�v���O�(K��ښ-gd�^�:�ު}Z��Tz.����W�Ԯ��e={�n�o��+�l2��"��K,������Ը�ЅF��d�Ӈu��.YI���=/!�Gj��(h���M��āQ�<(Q4X��+���d��s�m�G5&�O3�-z�?@�Y��,>��I8�P�pi�g�x쏬���Q�͌F�Q��=�d�1˽��譯X�����#����m@A�wd:)J��՝.�
~�A��CHY)�ﮩj����ş�j��AZ��f��@�
��:��f�{��>Gjh�u����8*���G�N�F׎j)Q�h#�&/(J/f���XCl�f�|a%�	��㽣����7��~Vz�8+Y�}�\!}����w�S��8G��z@8:;�(�㈁_�Y��D.���Jp�����L�s���B=���LP��<|ͤ~�ȸƇ<�j
�Ո+T���#~`��Vj3^,�X��Ԙ$]Orّ�Ԁ���I��Jڛ%����d�2�E�8�CoA�*~4d��7��/JgW��(RA����E�=��N�>\R��$�W^eК��5є$Fe�����P�$�ɹ���Kaa�K��eb^�ĺd����H>��j׃��/(���A+�T`��{;B���Vm�	UU�IY���x��~�H�R�T[���(�$���p���[*�Ǿ%(FZF�~oR%���Z](;^�w�Ꭽ����,d8q�k���=�`70������D��J��XՁ.��B��&�0�}�@@Եgŉ����AV3��@z�g�%���yV݈��G�?��}��jx��Q�9�l������l�ހ�g��}m��3
3s���Eػ�����v^C��F�/	+Y�޴Rf�"sBfCų�:��� ��'���N��%S>�0�,Y��#�H��'5���H����E�j�T�eUa��"��`�AG�6�R�֡4,j��Z��Kq D��^p_`MwT���x�`��E��&Lܟ�tYM��}��9���T��J����%1��`"���K��R5�J|<�Gtn���ܧ�^�&m�:�fLUܱYhb'>?���+�{a{��0>�,���3����F�"|�'*�O�J��#�jN�?�u�S∫צ�Œ�����Q��Ԫ�)���#�lb�T�5!�w�tl0�#�ſD2�3�FJ��Y���c}eݢ8� ;@��6_?M���O�HcH�"��P�+��Gh#'�ܡB?����ERE6d�:��1M'G�>@#����
i�3]�ei�.�1������/o�D-��&/D�jf� �K=�v^L����l��-�1홈�^+�>�����w:���-j!zb���kN4o�2�B�I�l1-8�Y&Y��Z���=���.��M�>6R�Z���{τ��4-�s��� �>�f�J���q�q����X^ݩz��8����f���j��%��L�y=�Zf�H����[ ~��1iv��I:��wS�B�nk;�Y�-fѝ�6��#D47uKɫiS�$�6Ѱ�blTY��nD��/��Bl3x�ˆ�>$=��qk|փN����Eϗ��V��<�f�/�ڼ���w@�fcvɖZ�8G�Iu�1���~Ș��F�4!)�������I�K�}q�6���NlL����O������g���U?����h6��/x��'�������*�e�7T:�$��j7z�2�g������}�w�VxnoM`|��R�.���֘��o�)��X���$d�d���%=���6�w����19���t�G-��9����Y��e�����;|�țG������MNѬ�������|�1n���FP�Xh�VYĬ���M��,��X���J�={J�-@{�,�１�.m~���Z_w1�KC�.÷�[`�D�-]˕����.�F��I(%�'�_�i⊰����\
��Pս
�r�	��i$f���R���d��D,� �n�Qt�C�:��Ap�]W����;jT��j��	���Sy���T�����H"��u��]|��_�&D�i�a>�T�=XV⤫�\���M�{�3���*1� �asl��r<v�f]�'�[@
�ݿ�F�G?4����x�G8=�tk=�7�z�V���g�ӱYn�ġֹ�t�E��N��m>�-�	�������/G+�/�3��Bb����*�d��A<�C~'�����[و��.�PJ�4�Iǝo�r���Ң]G[$U�����z{J�і�=���&��VQ"n��k����x�ډ<�Ǵډ����hn���t|�����������$��1ez-0�C�*k�T���(���b'��l�,����r��gTg��z�Ib�8���'�0��f=�H��n���Y�������C����1u�,�y6�3S���O�g ���T�_��.�~�qdK�R��rq�x��3l��+��9�� m�>��X��3ć|Hu�;��{��[�y$nV�/&������)����ك������}xy5SW`�|�SMA��}�[h��д�-1Pї[�]t/Ӷ�*�s�o������*.o�Y�?���GK�nR�}��[d��M�JU�RE�w1��!"�;��Q��V3��+�9;����P�:�e�k�����*hV<�;^��b���j^ ���\nՔg�յ�5���׳0�̵��p>F��:��J��!|m�U�:'��cܑF5���=kl�'��q۷�MGHActr]��S��Ui��������
������6X���|ݛ�9X����>���/:R�u�j7}�BQ2��'gc@4w�b<�TC��2��z�ꍤјD��Ҋ_I�8�"G��͈�?�U�;�U]X��3��!/Z�U\9ї��Yb�V���k?��G�ab��Z�AL��*�W�I$0�JfJ��ٍh��WM,��P�۱��do!*6d��+�O5�=���P~H�ᠦk��_��]�8�W*���6�s��)q���7U	����P�]!��G7<���p�ƿ�r�p6p����^{��5���~����?#��Ov�򳽲,q׳�g�����iU�h�?y��H��Vs\���q�4F�uk�B�R�+�|<����0���)�C!� ���G�9��t~k5οF�<"����]��No�cVd����ȸ����<ѧ��&��,�,C��@z9��
7���~�͈��λ>��|��Yz�2p��1��b0�8\�R�UVvpXᛠo�D��#����>����%WMvmYR�vo��Bbd��wہlӏ3�v�4�ܛWy䩭h�iRJm�@��|�mi�[��oB6':4�
χ��齪A�1"n[���{��C��3�'�H�VXu�u�����i��;a����==��;�25��K�~��J���q8�*���r؃��	�m�[����tb�X�+Ч�B럻qA9��R�l��Y%P�x9�r���n���mv��?O����p�V����LyKk�P�RmE��l����c�2=k�0��~g�~:b�����{a�Σkk3�6�$�Ry�ْ�Ƿ��bJ�DMR������|<`���#-�?��b��*3�)E��hH��Ț@/�٭�?�>�1������0��IBb]
��t���Jg�ܗ��Z�Vs�/�/}e���I��ᶸQ@��TCC�ƥ�"c�X�+�f&6��ZM��kw�-9�Q�c�H�O*h�	��)m#��A�5����5V�jӍ����)�Vt�Ѯ��5,�-����Uh���%}Qnv��^��i^���m�h�l�?��j�*u�MY���8��NXF%��P,�pZȱ��eע�vu�6�}�*�#}W��E3V�l'V�ԅ��<� K稊'n��*��(zWxM>0�I��PpB9�@�Rua��8��[��y+Lz�YW�;4��=Te�&����>��(
�D鄈�q�����^�����}�O��2���o��ٸ�' ���� y��5�w�jS����W����������1|>�J����-k\E����~K �7�}C��o�˂J�z���C� KU��s����i����=��#(}D��e��N�5��|$�,�߬�jL�&�R�j���� ���T�7��0�]"ͱG�ͤ�F���mŖ?�x�����J�O�gjya���*�C��pX0���Wz[���*W��@���9*V�9�v��
�Q��֊�)��U�\L�b� �`���	�>3c��������~��