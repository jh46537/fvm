��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k{de���ӱ���!B�C��S�
b���p�V�13ρ�)�L1����,dLv�Ļ��c-d��t*�+"�����/0��7����"����Y �k��e�)�<��M&+��()KM�?�ٿ5/�90���.5۔d,�]���#�^�uT�!�]�Zӎ@D�񲺯��א]�B �PgG���;��Д6�PL[X1i���2�Hb�C���T:
wt3���Cbװ?��c�;��:e3�Ŗ������#]K�5����F�bdK�z��[��D=WIg��s�p��,
��0���/R��`(�,�2C�U]�¢�F���l��Ԋ#�w��*1�
�ԓ�"M^�K�b�d.A�����F�ڰ1h�Ԡt7�������!c��1KVI399����!����I�F�G,!�o/���H�k��!�P:���[9r(�!�Ȯ��
�C;G�o�Wzك��3Js�.ǁɺoQ�n�['�#�d$}������n�OF�K�~�+?K���AV�bM,`�!�f�U�,��� Ԯ>���.1�	*�Aݡi~y�8eݞ��s�N���K}�P��8E��ԧQ/��{��<��5&ܨ|h�Q#�LD����.�7:�+���:2|����gQ�u�N~����I�- {T�,�� �k�������_�}4H�7>�
��QiuSR���E�����Ɑ�T%�Q��϶ץ#-�~�/��1KR ���;>���PfC�J�4�5%aZ�!� W1����	a��T;D�ӱ)!3;�N￷ Df��p�I�]�W�=�������ԕ���CE ��$�^������<̄�Ne03s��UY�%y�0n⬾����;(w'�?h��������g����C�	�/,g����M͒�c��8j�ӊ���LfP�3GH��a��D%v����>�)j��&q7�4��wB��L�H�uO%����K�Z�2�E��;��6/��Va����:�+��#�=��_��}����#�A�ӱ����eI�d��ՉW��%hK$�,;��魺����7Bm�nv��޺L��+l����M�?X�a k� {����i8e{�eE��i�?�-����}`��\��C�{�<��W@Uhf�b+���gX�mԖw��#qh]W[N�ʼN�U8�� _sd*Pda� 83�A�7��WaP��[�Qtl����a,�v'�}��4]I�$ ":=�-�jq�p��}�ќ���h�������諑+�o��bR.� `��1d��"3�qJ4C�PxA:�����	U�sSK�ܴ�����>X�A�U�
����#!~��d�1�[i�wUy�.��P�<4�Qj�7�>,�fo?�ǎ3�$�o�@�R4,���(F4�