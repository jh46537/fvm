��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)����0a)|_�O'e��,i
2�l�:Sq���-�8�\��Zz22/E2���zZ^a�l�n���$`�����/j)��23�|�����̑Ƀ���R���p���Q�^��'�0�[e���r�_掹j��0`�q������Ċ(��R��hsMȼ�!��JR�4���:5\?�;�ͪ��1�V��ȗ2)�<���0אl��RX��w+R��F��,����Xn.W���م�D5��I*>�e�����5�7Y�ԅ{�E�U(%�j<0���7%�#�}�-�O4���&�Ǣ�}�v�ә�jEV�U?ꐙ,��<!jl��֣O�t�1:l�ə8 q���m��l�6�<ӼO E��&pTh�(�w翍�j�ſ[#c�;�qm'C��A_հٝ�������!KP�=T��-%�gw���n)Z]V���8a�F���K�J���R���U4/�@�_�wV�}���a8���P�L3�qh���h4�uy���ߵ�	7�z�wo�v�3ſk�2`�ǫ��V3y/�j�ګ�$�Aj7ѹ�S!7�cpe����ݭx�*��Z����������/���k>�f��_�|{ts��)�FW2�u�N�����hH����y������X���,�����,2�`0��۷������$'�Y�$�k� x��p����������u�=�*�f�c�4̘�V���<�M�ju_|���V�=}[����i�&lf
�o�r3��3f
��;�&�J��<t�q���`����qH�,��Uo}p=��Ϫ��E�(o�0~�D ��<�]W��2� _TP���z
�s5��g�k
��}���;�E�>�\��i��gG���/h�������ě�BDQ�(�s])����a�;#O�U�����H��k��.�2���4�z���_/� H�I� �����4見\��#wMg�����8FS�Hh��c��S*��VF u������S�"Yj�������� �p��^XΦu5\��>^�K��0�ƈa����.�4�Z*��o���t�p�;C扌dc�3���X���x��%�\.�Sri�p��;1m��lN0~ue�6$�>�zlW��xY�؊�Y��؏��V \�7C�/�f?�5?���Բ��rډ�9�kt���Y�����7�t��)b�v��������)'�n&EH������t���KۡMح��,�rr�7��A&b��Os�G%�e\+�X���2��R�;	M�XP|7�#�|N�]�h<Q�_-����;��#(��Y
�,��l�q1d�<34��KK:������Y�5��Q�7k0��� _���6`�9��
�C9���фPTW[˿�7�;C�2�<Bm�;82M�W��z�Ox���*C@%���<�${�L���� �8�UG��L�> �m���Pɾ�S��ơ���[�# �wJlbfJ_���0 d��nam�U�3Dc�\F�c3�e�	���"�Z)��o��p#O5�dnSS�w�H�ҹ�(�/�t���ݻ���UTo���35W^y1l"��}��-��+9�1p _pX��:sz J�U^��[�Ѯ�B�  ���}R�XJ��U�����\&�IEO�R�o���.��,TQդIK�:nR%0��$C`�Z�&��C9q�.iˏ�:�ӂ�St���n�M�!B0�M�ٍL_�Σ8L��6
�Tq��J�"�+�I���݁N�IP�mIP���h >d��?hrA'٢����Ƭ$p=cơ�[
�z�QC�F���y��k��\Y�B!��Nx������5�N_�ãX�VD�9�s��s�G����v}��������rF���4�(�-*����C���b�0�e+J}�f�[jKjag��$�X-g������y����g
���|��Ot�/�{l��ghT:0A�,�KdNۓ-�I�5��y���o	ՙ�\��ix�u@<�r�Ql*W)���.ήPO����x�A�f0+����[�Ut�w6��x�WK�ˁ�C�3VS��2���/b���C�2��s�T�2`�]���s����H�*��O�	��@�����!�S�h��͎jG�y��Q�O�1~�(��'[y�*9�*�w�!傂���5B�C����B��o�$���5q�,i�o۸�(z���n��1m:�C@1ya�X%&�������ά�%����}�k���e6�xi��Wt߮����F�{�w��J��K�ZIc�?����d0qTn�C�L�J~���8��3�� �8��o<�����O�Ikg�4�7�T!�P1gG+x|E�sJ}G�m|+?$|؋pT���br|?Q%��н�>��O�8��+����G���o�8v������A��RSaW$�ܧ���	Z%���-�^���wa��=����JU��k��[�v��0�A�:�5�c�����6����(��T@�rYI�2�+��;�!&�=U���`~����:����1P�����m��rQ1��M]��~I_�[,�Ǝ��C� ��Ds�"�+J�u�+=%ܪ�<�8�c �����8�Y�@���3�Kw�&(��s�?+ɚ�E!S������A�{��T�#��z�|�����CK]O!H�Nk!̌�-�|<͢� &���'�,Sy����'����z�������e%_,#'G�P	LA;xM�;\��	Ī@#��Kc�qI�gb�0$���n`������:��>���}��M�$F:JzR��h�KW;tIw|1`��d#�����Eݿ�ei��-��*���(H2�o]	Rg�0�����}˔,'�=n�~WвP4ջl~Y�{����,b��ƿ�83�#Pu�)�~j�F���F���NQ8g����jk:!����SD
�CKt{�S�ԃ�k^C���D�Z����o��-����د���7N�4�'��CJ���N�Рa`ژ����/VyB�p��2��Rd�/GM�a��i��VI�ǥj����ƷF��(	?�1	�)$}���0��W����n�7�@ٵw*��D�@q9y4�d��w<����Yw��D.�(h`>S��U��o)"��n��:��}��v�]tO��d���6gYS�<�l��e��"���Z�n���ܒ�z9ܸ@�j�ڈ��ᤚr���O;�ϰ���vspǥƨ����p�|Ac+o��|�r|�ν��{!^�]L��W]F�����,ɨ@ړ�^���G�k�k�a��uap�4��5L�)�d��~���/Z�ͷ$�5�ͼ:-�4[�a^S:ӌs��1fH5����{���:Fk�W�bM��X���}6�m�2�_ǳ=���4��T��y�D,Uu�lujC���LsR<5C�������5�4��OM�;ZVӈk?)�>f��Rm�r�䤎�M�	���X��z���+��tE�����U_��@�9z�1J����=���=3��9�O��5�/�_�`.p��F�>R��$�Iw^����G$����UQ��l����3Rz�*Ǘ*���OV�,"C7�e��H�[�@XV#!)������=���>�$M�h�X�����CV_ù����R�?E�n틞p�W��!�Ǉ q�i�h1T�a�`�{h�WjZ[Ȩ��v���}�o޵V�U�t�la�e���	A���h>�otGŝ5UK�	���n�AJз�A��&�9��$���,64��\)8=�,���<S!�1�g)�f�@ڱ��AB�o�p����&���I3�|��["9(g5��V�|r��
�y��j	Ů���dwj����GY�t>�e�s`����~��5�i5�W�}�& �؅j�n|TH�7_ԅ�%�@Xʦ����Ã�M�t6J���Q%C��T��qE[>c�-�lO&E��c���!��K_n\F�����MNv��Is�M
����܆�%W�}y�x<�yov�ܠ�}B�<��^��AC�^ڃ����p�G�l�@����+���@�D�O-�>�B���C-l�;+�B��u� G4��h{|ID*$�2O�%�]����`���b,�Em�Ht�/h������e�7�ُ�l�����e��i[,b�,� Ѡ���7@&���� 2w���0�2�Yj�ͥW���{v�����܄�А�w�n�(�����B��:����:��)uq�u%]U��+h��1�G`�g��=����.��?.�cz��e��sQ�y�uF�D3[���m2Y,���۾�ie���s�-����}\�v�����XB}�Y�Ũ4�����YB��]���{\X��w�A�Oy�ו��[��v���X������sY����De: p�M)F!�_%�
"B�~Ne��۸���5Yd1���		�{�eY}]�0�_��A��Mk�`��ꅑ���<e���R;�c��׃5�'�h�H��}
~��e�k��ԸHj��0z�f�@�¹N�T�f��-Ob�
D���f�r��ʂ�
�(8����_�`�9z��?�aM�uK�-.`/W� Z"����>o�"ƭh~�=xPT�^9/c?Z���ogر��K�i�'�'���O�PH&�u�ú��G�sZ];���"�'W��7����Wf��z��ν�n ��|��?����2!?(���G��_F��&-��;b��1.��%i�_ ��O��x�0��(�Q�K1�E��]a�*|ʢ�z��}a�����f⩓����Z;p$�_��M�?J}Au�C�x�~���|Y���)xI"~˯VZ&�ۈ�Ё�zi��筽�����iF �Ҏ�a���>2�4�M��S��'�\:}g�h�ht�UIx�HO~=��� �1�˗#Bʿ� ϩ��f�OaqC2r��}^;@'Ջ-�͌�j�����"�����,zș�����0-��w�K�)(��L��)�'�2@��CV���9C��_6��0�(95*��uz6��x�(�����QB�\m!���xO�ňl����m�<���k�I��0���j��CmƘx����ʝ���C$9Ze����N���W��D/�B�'��,�N�N2�ނ��#L+1V�x�����8M��t(�C�h���ʅ!��aD�ͤH􂔚����c�%�����io�0��?|�X$^VI)��,��D([R�V����g����hNAިݽ�ϚM#�G�]�`��dWŀ=�	�Y�lS�&�@�����`�Л�eON���*���`�j�Q�M��Ey炾��z�*����;�p���$�I����!D��pLʪ�l�j�TA���_�x^��	�p��`�Z�7Gc~�xڰ$X�ҡ���P�W� �7�Bzj���1�L�#�6���;l������e!�����jY^wdI$B�a'x�����"C�0��Y�ɕq6��B�05���H���}�i��d1Oc��4�>�q-?���w�)�a� �{f�st;#�\q��I-P��
J>��n�k���|M��ܘ�_�^�%��;��8FJ���|5��C��R�)h�CP�f���oG�bc��50���x�1Ի��h qK�'K͛w�Ӳ�}M�>����V�&#���+�������/,jK�J��(]���_�b|Ř!�j�A2o%�'0�B��m�}r�rɾ� p��w@o}��ܙl+b<���\!��
J�f�ߙ��̡۩"���N+�����$KH�4�$��h�Հ��3v~Vf�XGZ�������]��(*~�<�F��	͕���懞+��efZP>�P{�eZ���WH:?wBv�銣v�>:l�/��D"WM.���1��l>L��:�?���ia��;[P/�f��ڨ6��Q�wc��������}���p���nI�r�	�va��t��[Ua[_3�5�^�ԭ?<��t-3ɂbp4��Z�<B��~F�}���+	�%b�nR_�}�	�\���:�����o!r���p �N�)��RT�e���!�7J 9�U��d
���Y�^_Bw���������4����=v<��E�*T������ު�vቢK�Vx���ēn��˝��T�p"�Am$wba�R{V���fS��c#ag�Śp��lu��2���\�r-mD~�^LwK&�|#1�}�{$���*�2l�c�OW��A4��æ�X���Ly���J=�����b�go�����l5[��Awf�dI�ˠ�V�w�m���/p��M�g��:9p(I:O�̝�y�"K��'X��zS�����c�Ck�'�Wq��������!�~%sYr{I|q�/�lX����YP�~MձIH��4�v���ש�l*�\S�`;��v�lCﰬ�s�Ӭ�A���`.pZ��? /@~��M6��	 �U�c��J�S�y�S��ލDNI49��|m��P�=��E.��]Z�O]���[vc�=r� ��Yr��5��k͍����jJj"}c�eFh�T�'�� :\�^�E&iH�j=1�NLDG�M���v�fÒ���3�t��^�;�-�|��@�=��vK��!�"�S��i�p�Q{���ұm��0f�L*L֨�N(�!�M9m�}�y��n������0�r��T�}�cH֕�M�E�&��56R�:k�W������(�_��7�>%7N���Rk���-V�����[uN�cB�ۏ�S�ض�#�I�n.`h!M��-�Y
����%�ZD"|y]ps;E�)B� a0a�)���6K�唒����C	�x�D�X�Y�N�d=�#���J����Md����!8yU�6<X�3�S���*]d�4jSJ��j�	�$��gR�HL '��X����)hb���.��s?Kvf�V�?�R@����L�I=�6�l�^�ߙ��>���}�����+7���6�}�W*�H���3�űL)�;���N=�d/��WJr��g����vYФ�2�eQ�ٶ�<K(N'ĚE�&��?��`r%��(A��e
}�	M6 �+�6��BOW&`����okc�"k�sw< D��à"^T&ks�[B�ٗ#v܋��X�8,h�gEJ�jb�uk��8I8��!��ݝ�W����l�s�q���8�u�>�_�_��30Z%���1e��� ��K�+�����d0H�>V���w�����BMS��[߀jCO�����#���^Y� �=�����B��'�9\V��'����ʧ���?�Ɍ���ܱ�g �#0�|��m�����"u�׶\I�&F?��ŵ.���2 ��p�����ƥ��] ���mz,�Jd9�4���4��e�<�+��N����G6�k�]2��Y�,�>���S�x3��;��:��
fV�տDw�3!��6��I��Fy��|���;��Sx&���(pO7UpA_�|7¨ubɘf�?�X��=l��탴a. ���-�Z:M�.�l%��GGN;�r�?��BJ+9��:!�_��]���li�X��k���@tF1d���e$C���?��ӎ�e^�B{=[�?wV� �t�X�@�3L�	�J��e�v��rW2�M��t�.x�E�U:j�K�\FUP��>�4��Y]�R�r�8ʚ3n��u#1�%|b��܍��Z�@f��wq��t�Ω��e6�.�1S�bM�
�Pz���}ڍ���g��N���^Դ���|`S~�hg:ꊄ0~�(m_�e�%�
�3l�,d�A��*!t�,��JnƤ�;��"�<�_�u�l:����e����k�e|NĄ���m]�H9 �)ECߌ�k\Ä�;��G�T͗2��S�K	&��vǪ��i��=����w6���;LI�Aн��iZ�����_*u�q�6�(үn&e����9t�]\B�\���X��i���L�W�әΏ��h���,�?�Z|K�@�8��?��k���|P������6tN�ǃ�{=��p"a�Mt̴n����oY�YU�~�_���w�o��"k��(����*�K�81�Q��Yv����R�d�5k�w��/Pa�Y���X����O������L�{U=g|љ�n��a�����M ��zق�+O6�@��+E��D
��
�T S��lm38�B����w��uˈ�29�m�m�\���5x�g����}�|(,�F
�X����&s<uU���U����m�%S��w��:�(>��<�n�ls�9�s�.�9ו�T���6�N��l&��y�mL�*�T�D2��FW[��9-� 5����{C�\�/���k�a��e�q˯Y;��%��@	�3�fV��5�@`�b̂	�\��W���Y<������G�E��]�럆�o���\�*����	s_=������ b����И�����Z��*��@;�Tb�'��Z��b�� 7���Z����9Lv�몼s��1�2a��"`��&z�w��ilf4j�Yqky�UĽ�E4��k��u��������1�Z���ٵ
��(��m�QMIЛZ�.�ԢT�L�;\�M+��� ةej2���_P�5��[�W$ܵ�i"isX�*F(
`1�y�9���=H�|��>d��(݈�>s'���	z?EVtC��K%���[�p)_$Ԍ��n9��T�yK#-:�޸��P�K1��-�a\�A$��f������|�cAiR��/D�_sg��͛�Ku�4�G��40����Y��oNQ�L��|���$>�r�)V�����i&���CNgS7��yD�lM]-����ԯ`8QĴ����ڳ� ���N&=��������`*����q��9��I�&�|��>��QcPv��·�.���C�g5�B����uk�^�CKq����GG)�4,��rP�4�i��(�A�J��Ň?L���B-�Ņ�ŋ�4�j$���̽�������S����sp� �'䷥M�����G/.�������̦��fbwt�j�:K*�v�m)�hU���D׫B�^���֦��K:dU��Q�!������.H���J����˘M+�s��=��w\�f$����A��0�&��{F$LB�d�n;��(\e�����4'	�:���P��Dt���j��}j�d1��"'('����Yqp��p��X�6!'o~ѱ���g�U6�r+H��(G�آ����-���,����_G�Iý��
��q�#Y9v�d4���q�����<�ߚ����T�f�.m�,�%d*�1�6�ϴ:�L�>*��y�l���ԢdH��Su�{}x�Z�o�P�d��:M!��u>����;����s׷V�2��rK ��hYHD���Xk�{RMn���kM�8��5���H|��Q�b�a�a���r�b5��Xg�s5���K����Ƹ�9	BxYZo�{�3�°���x>-_<�h4���=Q�jЗ��=vlt�K�f�xf�R�u1U	�	��ԑEz�$��۪�M	����Ǖߊl���5b�׬�?I��7X���ؼ!�qU���+[�kc�*�Q�A�mE�wJЯv�_�T 9��)�͓
���jx��kz��w7}�3��P���A�fF0K�5Ɨ>ǲ�Wh� �|�"�����N�O�rlqm�f�=����Ӑ�C��-��=�S���P�r�%�'��b�|�F^6\��_���&�M�A����Ho�_��Gc#�h�c��k�a���\��=iL�\�]s��x�J�uˢb��DX*&7��XF��.�qf�NQ�t�� >����xk����*��Ch��>��ï2-��T�Ádt��[�������.68ͥ����00t������mڡ�C@��w�_�''ց8���۰��0d�6]�,ubr�m��Trl�=Ip��##�=�j�T'��{��-�)��)�U����
��.:�'���~/|~6����&rH���i�[��n;�e�'r�M��,�� ����+�=��̣$�~�2$%wT��k�O�����+���=FxRQ��[��/�l6�	�����W�4����n�d�y�_�\��4�f�fh~�,��|t���?I�+ț'2_2��?އ�������3�w?��2���0�$�L?���*���u��$7/3��r%���7 8{��%f�c�+k�i�a��ڍ�vc��d0=�����b2+6;O�U?E���Y�{#�|��)K��A��x�L��D~yDvNH�
����J>�7��$e��@�
�kc��gB�R�R���(�^d&1-G�.�ș"�dB1�A�`�eF�Ymԯ��e�VJ��v>.	X�kc�bZq��Hl�LȺ/���U0m���T��͙}��E6`ʤ�Όu��UW�:��&��E���1��|q� ���C�P�!�Rg[�}�)��=����2�Q��c�XBR�6��@�cXL�wG�Gc`�~7~8d��b��kF�D��~�UR���#�k����'g7�����2���v�f|O�Cv�-�	W ����o��@TN�Ȧ0ky7"��cyI���;6[I���?��KA۴�\��?�(��h�d�w97n�^&�-������!`R.�:�v�́�5��ӌ��	kJ(F�pmpTxS>#���F����g����U�ER�"k��1�ؐ��o���{L�_�� %�{�S䫑@q����
Y�9R>k���r��@���e]�2���xB��[�˙�Wv�g���V�D�
�TT����	-�B�X*��d�wpe�:7��.���U�w[��ĺ�{�[�6*U5$�3�QG��
,h����Q�yxX��P�^_�Bޫ�O��>��������B�m��Ӑr�b�]`��I�4]��S�I�n5��t�i����z�4�N���<�)�B��')ѕ�IX�0��	e�=�7!R�6�����µQP��t��f�s�ms�s��!��ar!~}�dDt~O�i8�=.j}���!�uU�����I�ޒM;b�K��9i��W ٚ��9������(�[P6+\s����92�����q��h�f٨C?��PXdДxC0�S�������fS/����[�ʒ����~�9�3h0l���,�J}�=���Z�on�nS���ƒ�z^�\�/#I�ZV��0��З�D�t)R�yH��Kf�f:J�A�;*��"9��T�����3�.�=��G��s����[v(��6~tE뫈�ԟ�I{Ϊ�&U���⌽���:��=^�ڬ�W5nԇ�v@���a���ޞ,0g2"���+��8r�>Q� WT��TX�!�Lky]��fߧ��U#g7��z���pC�Uv".�8�r�}�\'/��U$�T@����������2��p���5��+��!�>52�>��UK$���k
��!QE�R����I׾���/�)�C��C)�!�@����� -{P��C���,0��Ƒ��mm�:����Ն|�NT���<�=Z�,��Q4	6�u8P�O3�¿n	ߙ��ay��ȗcI ǹ4�5�߰���n�z3�*�sUF�"���F���^"�ݡL�,Ü0�X�#6�rB�ЧȰ���op���U���8$o�Z�+�{���6ω���&Ǌu��%��pC|΢��s���'.��;j�,@ ���76�b���5�����M�����ѤM����ǦK�
סּS�����w���_����h��n��� ����0�����r�߿����+5gH ���M�cj���6�j�q�T�������_�Ԓ�eџ�Rvc��⥝s�P����y�O�`�Ws�~�H�T��+��2���@A*� ܛ?A�5��b
�����%�6���٦��rG�H��&�j g��|m�&)�GIӷvG�L��rM�6��h֓d'��qIՔ#��"\Q�9��{�lt=��t갡�gc"Ӱ枱�e(��k�A��S��q�E�(��O�`ǆ���;#�8R*͒և��w��&KUݥ����BַV�G��*C�j�W <�lO|9B���L/A�n���Tz�M_�:j�i�8��9STO��T6�	zѷå���4�l����ν�R��Qv�Ʈ���� �X�����^�=8���s�cqNT30�+��h�X��]���A9Pc
@���ڪ�RPy�?Po� u CI�
+�p�z�i��`�s����	C]���iy�#�G�
V��vQ��Z����L/�f��K��Q��QZ
���N�:�4Rh��(��7�<&Ը�f��W�.�����N��nN8G��J��( by=I��[���z��K?��" ����Эl)R�ob(�!�i��S�$��3t�4�2��Ծ��b���{	��<Ie���B �O��;6����'�D��f��c�%�]3o�}�����fUӿ�r� m��N��KpF�A��a�m�c��j������46](Eku�Wg�e���|����A��k:(J������=@ش���c�^
�3#�8�N��o�wD��&BqF�Wog�cA�R��gbiJ�Ҵ.B5�g��y�f��=���J��uװ44N����!�B�\`"�t,;9f�ळ�� �J����l��/_����eU�f�P�25fNbz�=�WXۙ{��zb������[{l��l�M�Aq�sob`���Ӎ�9^����m��h&S��|2���P���Y/��+3;��t-vL��Lu�&b���l�l�V���j�Jݹy {��j�3%�v���F�ƌ
n��_	M7���(�v9�΄���3�z�L��a�_��{J@�q+\�Y^�V�~�Kw&��&��\�8�j��y� ����i��N����r�3��_o�f�;wV����x�OH�.m�k�k��A��P$]b��7�4�-}����G}�5uXe��bqJ��F��nz�L����y
I����5bů$�����%�D�*�++Evt`3ekbE�@����������� �솑xc�*	[!.�a��(֚\������^���W�d��=qd��Y����^��bp��o�g�N�;6-�EGZ�;�}���yz�=h�CC���;y�Fg�~a���\����w_�!'��u�Ύ��&8����l�������!���<�`]��eo7�
>���-�(��1��t�P�t]<O�#�2�m�$|�Zu���ol��t�dQ*�J\���sD��bI���O\F���}(a���k�\
tVuKp�٣��kh�D��k��$��%���Ho�AJ�d����܊@zT�4��q�2N�u��:���F��<͘D�ga�%�0{��3����K:ƛ}�����_l�z��jG2���"�²��et#���a	�����^�Bc����S�`7;�X؋f)`*�5�C�r�Q��v�`��sj)㱰�q��MKŦ���F�B�C��v��1O�'�'�N���\M�Q ��(�僒��FE4e��D�����>�j�xM�E>Q �^�<����Z	OZ�!������O v�����5#P��%~���n�M^�)�UT%}\�hd�8.��ұ��A��f� � ��alF��^dR���zRO6����i�?�j�c߲.���Cx�Z�\Ba�����zP8I��HM�>u)tB�ɿ=������%6����c��P��l��>��>�+��r.^f�jR�F�"�6䨰�O��y��]-9�f!���g���ɥy3�b+39F��y+�.+g/�;%�/�9C7��P��\v��Y� ����_Vԏx�|0��\+�3|Ť���4w&y$T:p~J/O@�͋8��LĦLG�����R<���M��@7b�y��` |�*6	�Ѫ�:�<��tg�<R\(���g�Y��j��q���9�#��|ٴe9_���mYS�,b����i'x�����B�qLW��PR�m��m�h�0��㨻9���j�^JP�ȓBO�x�_-����xQ�-PΫ����̒��#'��;A�_�v�&۱QxP9�0���~�9̳OG	�:	5�_��k����[�WJW?��W��˭Ɨ��/S�����IR��չT=]?H\w��G��o�ea����7}JF��Ѭ[h).0�E����s��Ǚ3�����$4T��٫��zF,��>Rq�aCk�YX�(��#J��׶�n-BY��᠑��$5h�|�N`<�(;�Q>�J���=�e�C"X�ť<�6�M��qN� P��3L�� �ɠVw�����9�+��PO��@����A���u�(0WrMA㩠.��6�yRa-�A�PJ$JuZ���8alTM]o��z�M�~fm��D�t� e�g0bn��J��]�8��~�Ƿ�Zjv�h=��� )���yd:�L���+X�u��@w����8Y?�ה�� N����� 3��a�h��Dr�9� =9��Yη�\�����gmfk!��44����l��nc���-i�j��J�{���N�ܭ0�+P��4�A[EJ��;ɱ�K����!O*s8��x-�cw�!Dl�VC��ȉqG������7q����3�y=�;UN�Qٮ�u���fR�����a�6�W4	=�k�W�`clF�vDT��a��e?��%B�9Љ-���a�:�����$�(��klL��}u��wR���RA�Hy햡cW��Ta�U$����9(����f����iWw]��P��K;�8݊�e�P �6�N�f����;�(\��<	I�(
�˪���;�T}��-�Wl�n'�/5����H��!ے����%P��=�xc^��]>(qN�RQ^�_ e�>w��8Y`����2W�=�+�ď��K�*��мw�7����N|8<0;��濚�E!4����q��-�~��qZ��D/�P�/�\S�|n*�M ��)�S���z#|"�J�^8s�o+����jŲ"W��t��ӋN�.��x� ��L����v�6��#�~�\�x��rO��> |�(�4p6jB�8WhW}#��d�J�Z�(Q�t��'��gE�)=opN�U��Cx�N�c��S}�@*�H��w�rYq�)����H�}�0�B�'aS�����%!�{0}����(׬���5jM�mF�PQ�{�r����
�>S��3w:Cx�爛��E�~�M�!+t�N�p�/Ћ6:�u��#�֌�Ώ�d,��ܟ�Of�����|Od�]ϗ:(�_:N�!���ʳ����� R����XÈ�Z�:�WY3O���Bc�Vӵ�v��EC�0s�M2�o��HZ�vQ=ː��w��E�Xbӱ���d��|G�_H�2��k(��30Ch�w�=.�˔����Xp��]�C���M�����,F�Eū,��B Q��@�b2)��0�r���t�� I��Ll舎Ï��* {y��X](PF{[�OЂ��$	G'��{��*�;���%�yD�]�(�I��T�=to������\ʃ����]��L'����'����}��=�p#�su1p|;T���O��-�/!5�śM��E���bB8 $�5<�\�������PGс�i�C�����F��Vl�\��z�A��cs
%�L���Q¿�������ł��wA?pn}�pZXZ7{%]�7��ǮD�#�QX�ɆN�?�k}�	��^���}vY�5�t��~=r6��|R=����X�#�{�9x�*�'}�њe�6�7��j,����JM���i�T0���,�@-����U�ߘ�AF.KlA�5�(O����E�[Vk��d�@��(E8`ʪ�s�I�zYo"@��q~R���9�ux��d���zj�{�f��2d�hB�o¡�G������n�}߬�%���o璔Z��j��P��D! ~�#'�dH>k~=���G�.�� �?�&�$�-ςF��+�����AE��|��!b��?��|/mj*����>����Xe���^��x���r��a����XwƓ�2h��מ�`��4�b�ȫk��l�>�����M���V���Mmg��@s[B�/�� z��_dOB4[�Ef �fC-��ec]tyb�pۊw�X^�P���Ԕ�<�3���λ8"B&/��A�M�+m�H�ߟ3E���y1���ܨ��#gV�O���*����wT�X����YM��Q��LyAQ��@2'�̴v�A��7�.pL��.�uW�զ�[q��D���.X�I{\�[qa��cF��vZ�9�\Ps6f��n̒����$�O�g�m�21Dݡ�j���j�X"y�`�^����v�ī4ŕ��]p0�^� ��;��.Ws%����K���Ԙ�uQ��S�6��m����-숱<:M:��[Za�G�}�����.U8�;�g@��̓���u�a��3��w���1����W�殁m���T�~�aX��Eo����c��2���h|\;AK��)T�^H��F�J�#>X!wSp��rt]�͢�偌�E�������:��B�� A:�r�H	I�����������:�l���(�2��8��:T�*�a� ��Yx?;�]YL��D�����72}�g��͖�i\������ˍ ��G(Z�D�3Ƞ�o,o��-���Viu���%d�&�xi�߄Dj1��0����`݃G��X3A�j~�t�����f:�۬�.�
�/�7�[�.�r�b���2p"�QD^��L)�Q�l_�s�W���!�G*�'�r0�/�y��p#ۦġ\�/K0�M�<7 �o�f�S˫>�hM��� �VN¤�k,���S�+[��q��";VDlP�\��fʘ"g�
�BLkx�_.@��V�{�hތ�I~EaƋ�:�6���xn]"`Ƶٹ��޴?��;���m��7@���Mq�Jh�Դ�)��>
����e�`6�gzrm��A���_k{��B=�Gv����	�\"�r=� �6�9�#���9{rO�e��R�P���[iB�\ ﷣�w�_�q�ݵ�>c,e��%��k"^�}�o�5�NfR-��
�}ۓs�'.ұ�*����yO�2Ѿ�s�M|�`���O�@d����ê�-�a��g����X ��l*�3/DlC{V=��y�(L�M�P��YC�ݩ�Ͷ;aF������N.l�PƊ�k�k{u����;���ܶ+F�$8zj-���ޡ��,) 1|�Zi�JB$55#���W��z�����ߦ�ɱ\���m�ރs��=���;��=iq��1�5�S�I�M	��!��9���8�R���ys�_����R�a^��a?�
��Y��<����6z�/ա "�7��N_��C�9h$��K�_$�Aډ��W���d����̍Z���ܣ��zءc�S73��7���D�W�|xC��0�27��e�;t;	}f��n�tu��1q�P m�&���Hm6qG6Ք?$a{e�4����pl5�W��r ��?O˯�a8�K��s���+��И���,|��,Rt
@���m�aD�6���1�Z��E�tlX�����C��V�wnu�s[�}����w4�g�,E�@$k��_���4���I�$���1XF���%�y�j�.E-/�7ޘ1VT;a��A��_Z�ː2�dQP����'4ɦ_ �ЭI��@�J׃u{((\�:^�B��~�_�v��=����#Y���V2�����Xc��">�O΀��V�I=�';��!�A��3���T�ϳ`�@�r^sP�~���}8��+�]��lJ�]� �����D��0}�?@�uT�~��C���d/��
5���<w,J���K�Z�7Vr�(��A�.�/V�涅$Nq�|�)�]1�g"�T�S�XlO~�@C����U�l8����ݡʶLțhVJ{�{ ��Lo?��7@7ޮ�Y�oS�j��s!���Z�|8�Д�jN�v�#�V�Pl���`~�o�g��Zb�q�COR��AJ[��>����ڜA���vo���t)5.d��,
Qo�<M������zT�S0�MbM��L����&F[
1Ϡ���ѭ{ �;�J�R>K�AK m�9J���[i4��N�c08�*� �����l7�u �����#*���Z�W4ݮp��yr�j:-�dPL	bA61	���pT���No�B���P'n��?6�V园��T�>U1��YD��(/�C�<��S9��5JJ���r{�	X<Y4�@�K�`D\T������\ԋZ9�jԒ���*�ů�9�"�'wNå8-���rR����.�������_�.�YʀJ	�S�dYC����p�N+��Z�O��ث��.4q����>�-N����<�Hn�%��r�C�a�fE�qݏ����~k�U��x�$L���,���Y��C�˱�aI�e�(�A�Es;<�~$��Y\����k����d�m&�%���E�q���@!���c��u���6�y�2'��j�%|�]����C���_.v��k�V
��X�f?��PJD�4F�T(ZMl�y�m�G���R�ܹk쁒����$M�Ŏ�dܗ����c[;������wd`�/hk�eUFP�K�P$M���������Z��s������lp�� �����DՎ��*Sw���ۂl'�yb�3�%-&	$�\�̳>�ʉ�j�Y&����#���������I���p����6Ր+e��Uf�T���c_��0:���X-�kq!lǟ�>	fgo���2y������3LR��Z����m_ӎa#w*:�C��X���|oG�3}s=�����0��������Z���*��p%)�I�܉�̝2����
���1]S���F�a��6��"�7#]�'-K���i,����+	bCnd��6�$�|�@%��щ��Ԁ��B�S����7�Pw�׫GF�.Sr��U=� �W)��m�O����5���Տ�UG�	y(����$���A���yq��Lֈ������ֿ+��@@_<����Y�ٴ_G��Z+t���]r���dn���e[.\�5]W� 6�V�(�5�?���/�o6�RyD����Y#�3�BCa��$��>�c�B�h��#�}����?ao���Qs�1� b��޺�A_\1_���濠Nk�w7z q�����h�B:=�����{�ȿX�M���n)6Gy`��Zo�����*�8�aO��
����5��ZH�[��w�M��a^��{,�89���t�+�	�#-N����I\i(h��:s�/6bIM�f��Ow X4�4�!�D�˰a!���F��*�?���ה�I`X2�OB#�5w��G.�%_٥I��qm�o��ؑ*ڍ�+��������n*�2|�D�gJ������P��m<�N��w���jY�fO�\�J��DI��47B1�ȱ6 p���cS�d�%�K�1T��` �D2n ?��d��ş�g������2�ң���.��)X��Zܔ�]��P��x�mDj����Gu��}����A�9�?��L�G���ӱ�����O�[�g0�J�#��>���I�zf��Mi����� �ef���p����\+�W� ��dR�3�{�ϖ�����*���#a@���r�d@W#G!z��rЮ�%�3o˔b�߻�u^9��L����w��^���#x��+Z�> ��y�ૐ���>%�n�ZS%X{$��k�ifۆ���?��>�Y,����	��h)�Ţsu5mK�����đ�y��B��"��o9[�/�-`���Ip��#P��{3ܺ34�k��jƟ���'Y����3�ڱ�r���M#��*Y�ʵ�2U`���+�ϗ;2ZW<5�n�ס��i!ӗ�*����E��k=�!�u���B�R�h5�Z�]�@��nP���B�|�v 5@��3�������q�����~�?&�hC�ʬg肧im?3޾H��U���1��F`=�wp�����5�;�m��]���GMP+��pPI�Ȗ �Q�c�g��C>�9��v�8���ѭ�l��Ϳ�q](<4�3�s4k+�¶{f?�ÈD���g��qw����,la��q���fL�C$�YX�>�Rܙ�vp�Ų��Y�>D(��S�}4�=���*sߢ�������t��!E�H�c�D���s�mE�)�?���=<��.��~h�Ŝ��#O?+���{pĜ[�hz,�IC��v�ͣ�K�zy��©��"����(g�Y���!��O�{��+Q�Բ��bJ��d�I�ɑ'�����f?��v����>�|4�p-�(:�鸰���!�<[��[�B�_Hw��#���1X��]���,$�^���8 ��0 }͖�2f�q�a�|j�\����N�4u#��tT�SL�q�\�<�@��T�#�c/=������O/�AX�*����g�D�HA �(�rozO��1wc	#��*<�uc4jbp2#bf!�]_�R#I��ej�m��)z�zB{���U)Q�����%P-��h�B�j�G�ʧ4�f<z�Ğ����?�@��t
���E�ߜ��v�K#;n=;�@�[@�U^+��*��Y�����W�7=�SW�-ΉE�F���5�N	\|�G"p<e_��sS��Ѹk���j�vMO�	yST[�,<7���`��/v.,���!4����8Ͷ#(B�<�V#��g�n�3�ՈΝ��$���w>�#z��qp�&�m֡�|4�����v�zm��4