��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb&t���3Ii>л����;�n��ѵ1��BM	�{ v����<n3v6�Ѕ�dcH
 ��6�_��%�l�ˣ�IWۂ���f�O*q�,֖����6	���i��͝�p9So�����,���9-8����Q�8:.7
��O�3�S����	/��,I��j����s�����s�������	�]K���WT%!Ϯ��s��3K�q�����9�����g��P��4�(}��+lV^�?�*O?E�@��ɢZDF��I�Mɀh��x7��B�E(
S`5 _�{�Q)d/4n������w�~kM;c�t�|�lʏ����pm"�����^�(��Qh��e�����r�C��)�~��Y�.O$i�NU}�֤�]�=-�����'-�N������f�i�r�N�\[H3��W�	@�q2�#~���:��u��'[�^gv_��H飣����4�.��u3#oէf�'���p�> ���.Ӹ��K��}J%C���ĕ�� ����o��9E3NҴׇeJlY��5�h,e�u���o�2��&�� �6��{g��߁8�"�(`�䈨����?Ԇ�8 YB�?����َ,�ٲ��,LȤo�����Xe�(��=�Jū��Fj���:�W_���)MEpd%Mԗa@���#d>���Vث�|`���q�}��%��*B�,yhȁ���(��:�����߃�Y���s<���/���s�K���1�(�4qJL7!�)�
V.�Oo�KY�D�@�M����p;�RV��k����?i���s�J���@�~II���Y�3T?���yT�q���b&��ad�?�^ �-cu����z��!׊�3�U�a����eg�������eeT���u�� Ӯ\���łYKir3m��hd"\�d{�@��0T}S@�2=���ߒ2R���ˬ$������1s���PO{M8���.��͍�"`U��8� �}�wxt3u�8(���dm<i��؋�t��e4&rO��$S�-�-�t�#�#Z�M0G7�H�� L9i��Y5�Ѝ����{
)��Ue�򪓢1x�=i=�uf�҃�'^��Z������S$���`O�0QX����$6']g�\"I+�nW3m�C���k3�X�	�vi?��X���������5�d'���4T�X���M]�y�(�Q��_R�i:42S�BDl���ȍw��&�Ō�<�����G�_��%�ZؾQ�u������� ��O�8�Uj�d+���Vt�K)�Y2Z)���eN&P��he��@ۜ�#�g��a��Y�A6t!���E�#tѥ<�c�#$$��E�x����гA;���f�|nƝ����50:qo̭���w����[�7ْ}��D�2&2~��ub�g;{ 㘄[���s�&���+�����z_����W}B���a��u_��B��24;ܩGF��Qu�}�����	N���8���'�[K+�	 e��M�r }�Li޴�3�U�����k��`]F�s�杞@��|�Q&����	�=�������j�M�'>_r�G��y^��5�0V�o �v�:��٢��M�E��L;nkq9��x�F��&��\ɡ�	�I���Q���.�~I8�+0B���)|L���OP�F#�X]�,�sj�,ز��ڙ_�,�,H�������FLa�o�j¥,�ڿ����r1:,˦']c֥��ܠ�q�i;9 �:p$5� ��h#��H�ĝ�HS]����h��tV���I-�IU3��Ņ�3c@��K�u�WC)H�N��[�6VA!���T ��S	���j�IX���#ɂ���f��� $z,=&,��=�Xm�C}� ��s�if�<R[k�Q��,���؇��FwBIW�B��V!����k����(��0
��l�:�+PX�*c�ߩ��վ)ݏ�XS�#��p�C��HQ�d�S�Vm�C���q�4�1���;����/���G���oH�BZ�ٝ��{]�D���?ʏ�3���BU���j��V���:Ǽ���d�o�5�����1/H��nCϲ��i8U��boL#$V��8��aP'����>�M�/`����z������FX��N
Fƿ�񈻟X�U2���^c�qPavu��~�����Xej^_�5S�� }���r@�~�)-c U�"6	��+�+�R����;헉Z�S#N|����dmh= ��uc^���x�A�K�j��� �N �=�n�Q�^e���u�'7�o�="�%���ð�Ćp�`���ǐ�(�x}.��{3޸WM��2Xp�A��t�w�U��(n7+�U���6���v��o&f Ҍ��8P#�%�,5N�bZ�/jM�ѓ�m�6:9�\6T"T�*�
��u1�IN$�k?���;6���0�ɓ@�X)���?��V� �BP]V^+(jp!��/��w�ij�6ID3r�E�1ガ
hmXL��6)�P7�]~ϛ�䧧�+	Ro�~�h���]���}�Ko� ��;��{%�H�s?��0qʪ�.�+��<�����CzW����2�6�ǖ���)������|�d��iA��^���:u�;�/����z$��#-�񸚴���_�b���jW�4�[�r�x$c�^��\?�/������0Ӝ�L����&���w]l��g� �-�7|Ұq�TE�m��p�M��_���"O���������˲�D�I��5,��D:�#`�&o�Ds�\��5����W;�/)���O��Y�	���I��R���V�a��ą��K1�NR��3]��ct1z��@�Vֽ0r_�c��N�ϗ7�M�I�L��Z���F
��n8d�*>���������Yd�|��J��s�:�M|�x��hhiT�.�'�.�Yrh�VB���j�S37�f�R��c�dAL4�4��$�yV�Tmy� ��F��آ���:����5	F�/�����?S�`Z&NXp$�jOJ��A� 3��7��S��6P9���N߸��`�@쩱;�њ|�3?u�ԍ�\��1���,/�4J���')�ᑮ��-{�s��W������X��t8���w��}�}!���Fi@xE��Z�Q	�=�"ծ+\d\3�l]Ȋ����E$2�}���װR�I�f2�B��2Q�v���sQ%����abn�1T��,x:+�������R�&3��� K�*��wK>�NOc�ak�ט?csGW;�;W��4�
�s-k�A�b�J8�)�Yd��F^W��Vr¬R�,��ۡ;���2���R�5S�;�W��+��)˄7� ���5�}��u�$�Uմg	d�IH�����
9�T�|�w7��r�^���/8	1�/\���9Ip�J%8���
�K���O��JV�x�X\�R'�f<�Ƃ�0��qn[��wy0D��G��W�bK �ҍq�\�J�������T��l�%�8�H��ȊN�WaU�
*��┅:��h= �:띫t0��RN�Qg����> ĞQ(R]`��VsN��v����'i��uNL���25�X�YV�o@�{֙�^��Yo"��;������(r�"?^��Q�a#���p �����򐛟��v�[p--�
�|#��\
�΀���o~�_	�����LA�S�.-��)R6�a�x��ȳ����9%��ד�Z�x;=VB�ʣ�����C�4�����;�����r�1U�p�̼�X�R����#񰀅~��$ekj��h��ofm�u�GT��x�\��$���c�� 9��O�H�qb��1ٔ��E�=�lt�dw�G�̴��dQ/ߚ'��go�q���TS}{%���/&��_i�KX#.�1�����W�~� ���8մ�9�cCR��������;ӭ]��#���nR��1�K.N�!��� �oq�mx&�^G����
�+d��J��Ԋy�EJ	���8k��V҉ɇO�q�0g`�}G��P�&���qń!Ã�6�U��rH�i:�p�رp�k�"pdl��t��;�z�:��M�ߛ�
|��!��b�3��@�y*�:���ս�0r�pځ���*�"R��8r&�)�8�����Z
5�H�I��f��|cW������=NY��)'�,��U���I��R��`��6�.��y��{���F�G�����}6�(��fN`��EM�.�q���)�M�P|{#��ۧ��_9��iך������:#��59m�_�oN� �|o�3S'.�<�oms��������#6�p��ⵝA/�ߴ��3p��#���Ы^�W[�t��n���K�.o3Կ]���)�^��zP���K�xR'�N���H�zZ�T�q�i4�J�B"�G{���g��u���<�%���Q�����kF���%�╺M�ǡ�`�f��CaG��<�[�$w���jE��Wt�O�]�iqL�(���󌞢���z������#
�)�"�R�ш}ce�F����Ϝ�ru?���չ�K��<��tRvi��d\�3�WЇDr^�b�U9,����-�M�5��{�av[[�D] =!7Cp2,9j�'����}�Y�hS�V	�˰��B�4����E��g>(�,P�B%?�AvI�dF3a�I��k� `B��;o�E��s�5�ES��TE�w�q|ʬ�ϋ���f�nt!�Ǣ��J5���St��1{4��-�-�yX�Fj1'oR@��a�Y����3���]�=7�]��ƻ*�� ,L춘o��B/g�턑o˵��\��i�i�,=S�*�K���y14�f���)0���[W���!���۟�b���6��|��-0�����Yr��=�ɲ��
�hhG)Ti�"����XA/���Az�>��_^�l&�f�W� ��r-f��E�u��k���0�_�!u�?��yVx�K>�ι���t���zI�9.���
N���R�d �v[2ľ���#>�Cye4���*nn�<�l�%�M� Kr���{��2�����l�v���'�ZCk�FS�����:�GB��!��w9W�ψ��v�YPBd;I3HJ"e�0A��=������R8)G�x�Ѳ7�ѝCFx��P�DF�}ƕsa5��R�N��[����wN��f����8�b[�yOgȖ����M�8�Vu5�Ǯ:��K�C)�hnX��Ir�R<rYQ�g�:��ʨܽIط2{�u�9���h<�������U����5���r�i�l,_���) $Y�
xW8T���v(��o��S�ٽ7֋�Mbh��hOȚ3� ����SQ��_5�s EK��#hx/ȴ��)f��R4 �$�Ӧ� �-�(k�c��A���/�(:_�\#4Y+?e���c�D!U�P{���9g�s�yI|S�γ���`����/�(�p�����nh���V"�=����ϪLC�g�{���un��1�8�Tԛ.H�ex��P���^�M�����0�"��u��̛$���j	��1ğ&8#Nf2��hE ���S���E?��e�2�}[Z����QgT���`��VNE	�&��Qɨ��k&m��zl���3l{�=JY�����2�ȃ�ziS�7x��XF��cȇ��L'����1��<�-�eAr=�z�v�/��⯶��]��(�\�ql�-�Rzl�)�b��Ӷ^�o�$�lEiǵ��aMe�w�rF��~�u](���u�^�9җm��NxdV����P��h�|�t��=[���U��&�gGQ��W�х ��x���Q�2=�s$-�%�=f.z��P5^\H�O9(#�{H�>�|]A3*��ak� 0z�`^j�WW�r�=u��bL�� �9w���j@� ً� "�(�|U�2��O��	=!�C'S����I����� ��Y��+$K#��5�g4V�z��VC��  7�����q?0t5z�/']�qe�pDû����W$�
�s\�b�˘1SQ���5�p��|�`� �3���cwF��ZI�"���M���j���e�N��ܾLGb��T��(����&l�Ժ�����LfL�s�W�t���p�\����`G�|��Ï� ��X�/��$�����'G�/��$��� �?�|���ȋ���VB�N�3��[G�E��F����8�����G��j��͞��Q��F�HI�B�v&��p7�R�vcT^�k�Z�W��m�8t�v&���s0�=��}�� =��Ic��XE���^R�v��"����G���M���
W�Hp���bma����S��L�����]��u�=�u��k��i ��c����f����=$���%�"3؊�a���^���ѨXg�޿ŀ�z�������~%���t����n�l��(��Z,�%L԰���]� 	��l�X���z�A$�!�q��S�Qf��>5"6��u�Gw���/t��L�:g���^�� [�m����,�6Qw���n6}��F��E6'�ˑd�� ��Ho��[�H��8�|����k�L�X���MӐ�D����ę�%���4�Ƭyu�r��E컳;���� (�4/�4>�J	�����������#�U��)H��5+����M�� 5i� "���,������B��g%s����R��e��³Fx���`�"(#�� �V��P� �MÛ~�+���h;AYDؐݚh���w�I�/�5�)�󉪣f��Iρ�*���t��?��VWE��33�r��:I�Ñ����3�Kc����C���B�/�l�"Up�Α��P��3K%����D�W��-C�ௐ���E�5]�SW�/�.z��q@r�0�E��.���
�W��� r������郃��_�U��JS�u��-|`�� �XR���2C�����+9e�t�-L�6�eE���qG2˨�S��� ����q����m�\R�������O�Z_�Ly�*����hAv��q��:��|K�*��8��=*��z�I�-1�5��Щ.�����K;�hȼW5u�L��:M�x;j�~���?�8j��Z֕ޠP@�Ȏ�͢��wފ�"T�W�+����]�X�i*~"�rQ��#������BF0\=3:� ~�R��:�ir+�?Q6�9��EB�<P{}�
O��lmi�ӸN�u�������W��N_�L�R=ua�*vsL:m��f��*��S}�G�l��Ԅ�T:�?R�����ӟ{L#?�E�
��O4%�Ȇ3&% �a���^��%GwH"�N
=u_G��)mw{���3Qt{����\ "�,�ޚ�ek��C��E�	�pc�6r�*���>����X���|Ϧ�|������ �Y�`�Ln�	����<�㯶�V_z1�8􇏣/�I�|���"?n�n�e���(ZiR��Հ{���J�$�ت�����š��@��gK4�[��ZUo0{�$�17�������ȡ}�g��S
�A�G�Z@�ւ"ݴ�ʥes��y��~w$�[�B`��U`OOJj�PEI������,iȒ!F�i[MC�_O3����i\�C��O�t�l!�Do�$��p���jx6�f����k����@v��T�L�Wi?x���c{Zq<�J���vq!n�s�^9?r���Z�:P@�@�r���&��Q>��	A��"��~^d�P������R�Cqz����3�p&Ё�S�6{ږ� 3u�1	�n�i��,s��o&H!��,ZqDҌ�+��0>��S�fh����t���@H۝DIy��>��y�����$�e�u�N��
�|��Px�ɼn*�����>�3��������h�����\&�%�f!�ZZ|�p}�z���E���S�?��&�4���@g��:ӽ����w�E��H�����LS�~Yx�m������%�#�ib�ɆU��Ys��E��Z7�8o*B�ݮZj'EHnί������uɠ�+�YJ�dd�з)'���m�����K{��t��=D��tٹ�u�{�?<O�x3U��扌�%�j�� ��Y*��k�Z3�To(tYP�KД]QSg���tdL@=iFn�e���Kڃ�a�h����!�Q�}�JӬ���@��H�f�E^�=���AH۟�[����"�q�]!c��E��U�+�^��H|�‾���`L+�ݚ���bO�_��I���H�m���y�e������!�v��|:�����Oiآ6ZX�ܥ���@���w5��2�m��}�py�-=k��]�~C��YT0#"FT��>x�>��ڧ0M�@�g� �2+�PV|���n#�{�_�|��|)3��udYЍ�{���q+r�릃N������>/k��+f��&j ���O�^�D���BUh���c&���vc�X���C�D�j���^x��W�pH��_2��l8&gR�7P�&ʧ�Î����K�Y8�q��ֹ��uR�//�2	tr��4n�q�����,~T�D�D�1}(<�O'�A ��!W[Gh�葭{��m{����Q2s�(��l�Y
=n�+V�c��GB����Q��/.`XŖ9��mܓss�NA�ǬF��:�����s���<���h8�3�.� ��Q<����]Dz�T�p�|�7��:��jW��dp�Y�/��ʿ�f4� ,Pc���'C�{�817�+��87� [����#�q-����\�8��4r�
*�~�ǻ�4��q:��
	l�	�ӬbWmlJ�Y��5�ܳn�l��B�~)�:Gj^�������J���W����x��Mf�T�}ʬw�ظ��,"r�8c�z��u���e���:������X�f�eb��׭�k2C	и� �_��>`�t}�o1H�ܾD����e2��ӳ�����Cn+p�}��p��٬�I�j'��
pb1�h�AW tqKp~b�0C �������f�,R������1WP|f�.<S�U8\.��+I�L3ۓ��1##&[�����d/�7E�K�T�r1�s��^GBYG):��ԗ�
Ӗ�`�IU����[���B��b���%�J.�� ���4�4K��BT�~Qqe;��?�y�Ծ�/9/:����׏3��.	��E^�'UXs��9��v`�qZ�%�J�L�-ʧ_�M]�X�0�G��� pc����Ԫ�D�C��	�����U���l��@
r�^!��:� \"�늌Ɉ��ڙ�N��إ�"�~E_D��~��ne���"-H�#֍���+\�T#ܛ^B.�#��d�������=�M s��͢d�灔�%�g܉�gO7�� �se��_w��%�0}M~��q�vn5�0u����^v�eWp;0�|0���|dAm����ps�ʖ���}���x�x;Ow��1U�Z��5�c��B�7bJ��O�[�"j+t�ϓ��n�>c={|��+x�8��s��-��L��֛��Tb(3�����R7�jn_���\�|-��jE��ǻ$���xe͇���
םg�+B�9M�K�S_n���N,4������ ny �<�LB}�����u��1Y�7(��0��%�Gw�m��;���B��n��<Ihqm6aT�L
|~F�����+J"�Uej63e`���._}���9Pw���A5���@6&S(���շ^� �2��C��u/0�Upx������D��z�ʶ�9�8��N���ʥ-�q� y�������1��O_P3ᾀ`�4����4g�m�����G���C·[�{16@F�_]:�dkE��]/���A�h�}ќpʇ�����j����%?@q�&�>���q7`4��qZ�)N�ц8�ƣy�e�	�j�n�]�G�''ܐUd��t ����Te`{S�ԏ�߈� {K���	��HLF�r��u/�CB��|x(��E����d�/O*�`����^v��h�A�%��m�,���>b�
��o�N/��d�1�� �#�\�d��4`�����J��e/q���c�W�V/�I솆ʓ|O(��UL효Z��+Sn,�F�L�Ĉ����ȇ�;��ζ���Q>D����~'����%4Ywa�� �m�IYW)�1�7J�����2vے#b�=��L�������"�<r�dB��J��	lbE8���=\_�ߥ�P��Qī��o9���$P�Գ�^湎'��ʬA���$S���C�1��#h|��)�����3C�ϫ�=(�|E���f� ���nxs�R%�z�ͳ5p����3nP��픐BG4�bY�>����������������¤��]#��f��T�t�d�6nW9�j�1@c8 ,�]��fT�lB�	�R��F�5Ќ`��T����)߈��S��}��zAD�c��v�]���~s�B�@C��bO5�=�?�/�e�����.�IU���jV�jbp'E�wC��/�%X��n8���D�LװK9:y3)��<\��]h��~a��`���	���^F��Ck1����7o��m�ԋ3*}X�Fq���\+vRχ��^��'l�f�,�=��r�E*:��)8�"����0�}M��������L�XN7Ղ+Dس�Iy|��,�M�J�)ؽ�g��,s�2,Etȕu��J��v4kK��°�x��� ��3�I�X�m��Vs\�Gu7��a}��<�,�R�!�+vb�af�Ow���� ]g�C'�:�$��I��ʁ���O��L�h��y+���sd!3�0O(�֍s�O2\O�a�c&J����2~�%Ɋ9�{� �[�D��gv��e�|��0��&&6���꒰��������Zs���e���K��Ţ�]��hl�NP?�!^`b��^�M�yizH{e-4�e��|�4Q�+X���1�TßYu��:A��hQ��&�х��&��� �X��_�;#�A[V&�'�t�'��1�Q �1	����@Hy��P��c�r'.�����
�>��o��W�o�C��0�r��b����B�g#��6�´���0���l ��m� ��X�/c��8�:'ڷy�Wr�'���JK�FͶV}qs`�Z�(A��z#��E�U�ț)����^��Ĕ]Tt�7��6�Wdp09�rl�N�'��u�?�i��G����B+�ʢGgG�#���Ӱ5u\�I�&n���@�f3���ʶ��:��eΕ��"��e�]�%r��e��~W����r�j�\z}��=&M.=.�1wе �vS6���_G�����̛t�;��YD6�@��7���Xdq�h��z�y�~��f璨w��kN0&�й���D�xT}�X~tDX�n|���6��2v�-TO��&y�C��1C<��x��C=4�T�2�o�+W�٪����k�S躝�SL�#Z[8��Ց������#ӳ����6�wѬ�d��3�َ�r,tN�'���l����j���Gb�S��K?|EO�N���8n(wo����-�LT6�ȣ��/�p"�o���r�*6/�/ G��GoG@B��1�ͭJ�IU	��h笰��;�h��޳�0ӥK1 Έ��b��0�KH:ϸ�c��E��/�1��j�q��+��mm�%+B���^���:�Je�-񬠀\��+�n}��c�cf�ZU"RX2�y�Iz��+���ta9� w�6����e����s�뙏�
�� �̠�9�]LNh�������%W,���lwO���n�І�!K�K��V��;=�r�@e�(w�T�`#�fWUZ�됹6Y��Ym�CJZ���f��ɥ }O�{U��dc��K2�w�z���rد���}%
d`�-��^����z�v^^q����A��� ��	�
���@���7��đ�%��UA��G���L%��/#lN�_�{私���n�=ao�E*��#m�;�;m��*��T��6L�qM�����鱗޶��s��9�=(�`�/zul�\/I��TB�����ǡ\~l��E�Q{i�솾�'�kr���VH,� ��rl��4�n���+_z��j��T'�`p���J���zdؔ�O!��p"��o�o��dn��姷�����]�e��g${�w�S�G@���h���� �nV +Ͳ�*�9�,���%�[1��^v8�[�����g���y�V���
T@�T��`��pp�|rD~��TS��!�5���P�̽Ԍ��QUoq5�/oA=�vC�?wǭDm_$~�*dJ��G8#x�zߤ��m^Jmzz�R_�4���ju�jR���$�{�	  ��")rW����!�����7ó���n���4O�����_-\��]x��,��W��b��GK�.� H��(��l�Y��	n��,P|�=?�g��I�;�˼i�%}S�إ��Tt��l�^��?{��Z��c]V����V�'���iA洽�R)C��;¨�f��n��E([��"��EV0�0���V��lf����`��*�� zg7���g����r���eq�z��6�H�����z�x��b�#�M��i��:k��t�v�7�u�0��d�s5��-��|��z`�z倁��G�0ɜ�W�{`����.��I7�}�ٖC���W����6��UD�y����6 �ryh�����@D��L^�憦 no��$�+�;�BI~�/�HXw�"dG�~�ˮ�8SX��DB}�y��P8wcW���.<i���L���,���a�oOR�]��%�Ųͨ#�ωXM2�sC�pp�KQ�K�
}D�9f�E� ��`�=��XЀ���GӁ�⥒�(2�4��̫��)��]��i ��)������;mA$nI`�
]���:��Q��/F�~6P��Qe��D�Sѧ�;+���k)+��� ��"0�O�\�4������43+�>�_�M�5[��	q[ �(R�O���[x�D��ﻉ�{Fv�����5w8m��$tv,7���N�p����.�ȿ`���E]ENטÁ0�e�)���h��C��8D]�\:�&�|�*�P��|̮v�|���2�_�;�yS��M�%�i7�2�y�� �A*�4�!��I-�ƻ���g5d�_�ƾ��r$C�A�d�?-z�k<s�y�d~)N�쩦���Rl��#�̐DQ�?]�o�g52��M��!�}�Bٓ0@ak�ʬ��rVS��l�cP�&efs�����ݸ��}�
ҿ�I���֞8k��*{�a��^�&e�x�D��6� e`�p�3�eMyA��a���tV��"T�!���0;��/8"@����b?�7V��RX�D��ư�G�oՂ��>Ů ���S���AJS����Tկ�����ª�'�TA���Ы�T�.r�y+���]9z�j��iShjzP�U2+4�4"�k�=����d�� �
����ce0����7�z4���g�gЉ$�H�I�!��0�X(����[�G��ҶƙhnrBY4���[	>������૔a7Ƒ�alR����0[�0�ݴ�v��Y�ڃ'c7G�KU��,���6[��o�HdV�������(�G6bee��8��Ƣ;��#���=ߌ�����¯�.lOyH��Y��ިÜ��Y-9��μp�37�'������ХaXtH�mD�� ��"[p�n����,(���/X%���E�����_��Γ�5Ù>�)��0��y���ת�����i_��G���t�9q�jrs�	J!Q�r��!P�2V�DN�̶@�M��N]f����^��a�;��_(���8h��//��R85@�F���7�6V���v�.��S-�0]���
zV�����L����-��P�K�oQ��k�L���FȃC��!\���y�p��`[(���J��H�Ã�γ�cV���s�Z��!/mUN}=����OZ���5�듭�ߣ2i_���U`M�~�:�xc���XA��Ub�V&��wߧp�X�M��2�8�d<8_����k��������I�X ��j�M�=�IZ,*�������w����:�"�AtN��:��4��u�p���L�b�a�K���sѤ.N���AF����F�!������`yI���~����I~�T']a��
.�����!YT�������QOs&x�/g��^���/N����7���0�>��E�ɠ�<{ȷ-3Q��q@2j�J�d|@�1sUE��N۬�͸���`��/�7|J��E�Z���g�	�L��n!����1��*�<�&`��~:~/l|U�ʹo��H����W�81�`%	�bT+���!�J|L���> .�q"\h�m���7?+G�^�L����e/ ��`t�c�k���#[
����hf#'γ�֑�<z��\U�S��"�93�\ ����5�G�����k�fy�7�˿`صv/�ڷ.]����+`�D�Y�<	��X����P^�������ڦw���y��R��`��w)����V�c��M4��5�E��C�K�>�φ$�f�Y�N#Q��GK�����c�6t�`��tZ�D/�v�{� 36=�b�ݰ(��}j��:��Mv��<%�kœ��W���n:N�Y΋Ԭ��)��F�����۶��z�Eͤ�O,����a�7rw�v����
�?]Hqb�����M±ܭ),�3�e�#��t�b�6s=a�(�H���q���#s}e	3L}W��F����~�h��)Ft'QҌr+8%��q�<�W#�Y��J�O�?���Y�Gu��i*��!�V��ួ��v�[�*۪����Z��<P��8�����8��QӸ�NĠ���@��bk��a��vTXP��8[�w}�)��Cٝ�mH��P��-Z���%�)��6m�	Uu�%pyc��aa�Rn�\�DBsWAtb�Eq�':��?H�A�;l���ݦ7��B.6��/`I����5�b;�M��W��r�M.i��=�K�����].u`=����Y&�Օ}�I�A�-̊�"n����Ai�E�J��v�.
��^�:f��KGֶ�Ԕ��֨1��\��|g��ը�(WN���vv@��;kA��/�v1_[l�(�>GT��Q�����<+<��&/59����pj�J���0H����HO�/��>�[@��nfu����C�ǘt�j��m��̽��u<�Ө����R����(�U�n�.�<1�W�V/iD����^Dx��\�^�^�;��8��24黖���� @����nxo���ɶDYV�1�_,ޤ�wV�����^&�C�)��:@�m]e$�`2���u�M(�~O.Ǥ�˖o[�����<����Ԃ�4+F� ����bc��yk-�Yt$Br���/�g�y����<e��+1��۱�����9�1Ĺ�TV�v�ꈾ���e8�!��(����Pz��_�W8���^'�z#��ԫ�!���e�nbC�{R�(^O��u�>��w½X�[`�pU�L��i&A	H�	W�|��X^S��2��`T�3J�"����\�%��fPx^@�)8T�1-��2?cm��G?�.�le�_�݆0�p��n�\�]d ���F��v6�B���-���	���Y婭��-��)���#<���;k�M���
�m0�B+��&/-��}a��ĵ��������ky�Q�-ƨ/�)ݏ�ۍN�b�MsF�1!r�+�uA/"�@|�q��m��}z�9�<e]�
]o@�?s�|��H��ѝ�.D5�y�͎�LZL�,�����q�a{�DM�͔3�z��b�e��;tv��c?�o�����{��d�9Ι�헑�)n3��ך���'�W��
L�g�`49d�^��� �o@�����E��p�$+��s���\�*���d�eUw��H�aU[�s�Hv�L���Dq>��g����[����M��A,�z�5�*�x��jo�EPk�ǡ��%�����>�s�'Oհ1�$�i�9^����)�����^^"��/���O��������TG��Ich�_��"�}d��2F��W6���'��ДV�}$���a'~�J~�i%5��{�J��~ ��[eߔī)d˓U�����	�_�4�JF,��9��U�p���q�tlxF$�9BN�]�k��Wm"�&&A����W۪����4��T���Ƒ4˟�}A�%R��(ү~���g�Vgw���$���x�(�/�����od���Y*gA�b�i��(`����g/A�74���id9nsSN���`�G7�����j2�wUJ��/i�	x��7����9�`M�P��r����1��68�'����Qߏ��o�=!&��� ^�k�n�����)�l�����P[�[o�y�`}Mi�����]To�=^7���з��w^�� �� :,7����*�u�J����R^e�Vvs�EMd0�oے�l� �-��qh��@���vE]�Q�����1#�r����d�r���6�Iuү1�v�("���w8��v�!Җ7�s�
8w�c�x/��f/�@��O������j��3�B>ۮ�����˻J��3� Sm`�Ʈ:(��*2We�ñ[�	@�Կ	a>�*"f2�J�՟��b�&�����hW�WU.��)�~��Cf�
���1vA��Kw��G�W�=��H┎s�`73�q�Ε���YU}��1�7�L��)���Fʤ��說��u�E�ho��5���� �[�&������ڶ�lg��Q�b�2D���(O_"����X���pV��Z�"[��`=����'��wG��GT��/ �|�����c��l���� |� <<*����<Y�f���m����3ӷ��J}�:Pj�`F5x� W�~�Z�eH�Z�c�|ۤ�-���I1R6*Й�е�v"� ���J/�����a�~��P2-�����o���}A����e����}R֠ʽ�(��)��0�ʻq�q� ��\o����#�~��cT�ę��-�5�!�����S�ԇ��������[<����n\H��X�㽍�w�

����l8�_�'9I��h�@�ȱ9�� � ��^���'�-�Ŵ_y�s��U��5^Y��Yo����$��8�*#3�= 9�vYb�eX�"�:�(xt|�'d_M�����瀆���������'+�E�5�ձ>=*9އ,xX����񀷖�<���v=�^��� Q�����յ���%�j��vY�{�@Ls��v��|�C���P��s�i�7�w!ǧJ��{���M��Q�|&�qwAH���)��B��J'h�wp��B���;�T����V�x��Ygn2p��ipl<Gf,]��zEA������ �"�+n���?��y!��<�\�C��y�y���c$+�n�ve�G���s�&�`"h=�w*G�Y��������~���d�m�NB�'S��0tY�����J��"��/��:��	Vr��(�\��?��%�0:��h�@�K��7ބ��a�i��2�]FMb+P�6����sv��q�w!M��>���_>�Q��f����~�âs��
�?$S'��?;7�BH���b���un81�L�	���}sE�91���H�)%�u�ҏ�.�J�AK�e5mA4�a�j�1���Ї��7�8J�yG�99���Y[q)n͋�**-i���Q���_��bN{��	[Ȫ�b�)��x��A�3&<�ց<[�|�]�g��¶3���1P��U�ꬒ�v���&��0:U0�v(JT�V�,%�M�����{3 �a��DVp��Ͳ}����H3D���+<��Ҽ@��4�ދ��!��&(s��(�ʁ�l�䰪c;��(�6q��RԨU��V��k��/�{i�&*�DǠa��Ԣ��H؟�5/WR+�����'PD��6vǸ\rI/N��ݰ,�tp�I�CGO`��� �����oΒP������e��ӒxM,����{}䡊���)��Œ��WQ�f\�aIa}�9�=���j ��2�DB}|��Ki�,FMVa��䢱ET��$ļ}
�$\����"��$�P�M!�Б��f�U��8����ط�H��4�|.�6t��I�B�R%k����RH� u��֊�,���#�rxz�<����|'�U:�ĕz9�**�"p_Q�h�ᅽOI3y5�|��ua7����,�~����dY0ֈ��b�.�B4^�`I�'V��}�JY���F뿺���w�g'�5/N�z�Ⱥ�g��h�-�m�'������D���Y'ި�z��?����4���ل��6�����S�y�a#�we9�|��΁��`��xcF�� %��Y{����S�c�����\u R���C�o�ȩ=Ab������%^�٘����h���;��G�����S���a��csFC�fTk��4��=,����oM��/1���2�[a�)L@������I�SpH�9=�� mq��
sk�]/XL�*¢]�´�<[Ũ>�b�D���B+��&j:A*R�����2�9I�)LI\�5I��������O�D��]uyeTX��R��6��)����
��

�<8�|�`81��4LT|c䐸(���RhTed�N�����ԁ��{������[�����XS��3�r��g�J����$dKS����n���'`���8?�|���8	ul�?�ؑ�W��1@��p�fu����e ���O����-_[k�����ٰ�Y�A��,3�j?�7�Oh����	���347�I��̣��pR�[�Mb�_�<�-�@*]F��P�le3p�<BV����>��~�C�����c���h.��/va�M�en��e	�s.z^e�T�̂��&���O��I!殳������a����?�	[O�C�xP(Z�~m��n���^;������-3�IbB����L3M�������FB�y�S�A�-'FX�r>-�W��i%������RW���J�^��4�����^��Gk��E�ű��YΕ`��4J��J=� �W�}Bf���Q�����&8�,�>�Xk8�v�Pc�z�{�L��Y��ې.o ���)&n�k�iv�(\��=�˻-c(��W9Cg�v^p�77�.��R>l&�? �'H��[eal��]���2�J��̙%�-�ܗH�7e�n$I�R��쐤cZ�e�B���o۔F�SWL1��u7"��WG���[�C���]��УA�Uo��W��3عQb����|�K�v��?bK���\�����������8�d���<�/�e�قRዬ�fU��h.aLd��TٜD��/���D��G�+2�Iak���J|���V
��������v\����
�M�D8Y$��˲��#�_����i�9%ؠ6�����h�Ү��E���x�Q{ӂ���)�2�w��W�#<�:����Z�X�*�zU�ɪ�D�S�E�mJ���q��$��.GNr"+y�e�Q�`bV� ��EnAͺm��$�?(�!^Dq9��Û��]?2�~W��1����OI-�vI(��Z���8��hk�f������Ђ5�����g]:`B�S�H�U���w)9�}3԰,n6Tx����sz7�~j���+�Z�!L��܅e�ʃ�jp���h�n��0��m˘xk�y5	�cuS�<��&8���y|Ո�����,�e��8*��xn��)���IR��7 7E+�a)))H�[ڍ��JgJ��-r|���qGA4�A�{Ӯb��F�̲�;t!��饺�T�L]��T��Ru���3�k~?���bf<�K�X�E!�zP<��o����z^ �uÙ�|MM��s�^��>�7��*���CmA��U�G�ލ�=�A��:��ɾ:,`��(�u(bf�orפ�a'�.�zVU��������o��t�k��`"=[$���[uz�*���� 'l�^%���MP�/�'�?Dנk�1�q�'��'ed����>�[��j�{�S7�m� ��_�+�����	�,�ߑ��l[��BF�!
�H�
��p(��Y� ��"��]Ip���,|���:�~qs�x-�V�j!�[Mj��0ƶ�݋�����r��.�G>�����*���Qx��{��_�;O�|�q�)�]�t�)��W2wY�	�!5����U �H��Ìk�8�芞��w�������_RT	H�)��3��V�zm�
b�`�l�E3*����䇪��t��8(��ۦd�}�s���� 1J�:T|2�-�l�	fL%P�ʀ��`�������'��8�c���gmйbx�O�)�����á��^!cr>5�-�(�4@(buGJ|�{��P)�����B�*���c��[?��'[�d�LG���BI����9�
�P3��B"C �4�BnV��e���6����rw� � �� P3�>~���x6vx�盝{��$�1�{Qÿ��/�*פ�6u�i��˳��� V�3G�� �$���V��M�<08��'����S�5�]��$�Xt�{�1���|�mA�	dU��DOn�7{tM�½�+����w#�ERh�3�ff��uQ�_#��@t��j�?��<���XEI��W�âCؾJ�Fz!��a�0I��k�[�+Ԉ�)�
:���	U�1ݛ�G�<痠��X�:\JX�A;��ve[�n�$�/n�C�W��f>��wzD�ٶG��>�=g�ޛ�PW�z�P{$h{��G��cJ�S���C��hu�bR l�f�����,@����+�����1kM�٨Nl�<ۖ�����O���!E��?P��c� ���T�F���D��_D�]�<�k-��� ��Z��u�Ąɗ<�b�8`шa�l��2#?e�V�����N�o����}_fR��6��l���|���=�)��ה��h���!�=�0l �řBe\k �P�5E�j`��p�W����4�����@Aq�lڪq�6C9�Wtt��䝪����;Eo:�][l����}�S��yGw�K�7@̏7ބ��>=XK��i��;	�g�G�������Ic��v�R�����)�λ����ubo��L�d�lX������A�1}ZxO^Z7h��'�r�6�ה�.��Ƽ2[�X�\'�S�R�8��EXP����5}`t��ԏ��|�oĜ+���aIgJ�H�ؔs��Bd��4A�#���!2tc�0+��'l��B=��Z��T�\uo�i�Z:V�
IG2�
b�����O_%$7 R�zG*~�����|5#�S��F��t�_0+�=��AsN���TI ���â�^-�̑������2�	֏�`���=�4 <���w&�Xr���SWG�饾�U�������MR�/��B+��k��.})8r��9�,�k^�쥥�ji��"���뺝������%���d��X��!?6�"	�����D{�q�zCʕ��#5b��������6L~K�}�U1��:��j�K[<��0�������`4тu	}�z�!7Za�H�#�z����R�� U��c���E�+x�����ZS�L�4Y$O�՜���uf��J���r�^MS�
�Q<�s~3��~K�	�����O�� $����wç����q�;����1��\��x���D�(jV2u�{$Ȳ�rEt�k����AwP��R�Jm_�L󽼧��(l9�^��U�1�پw�/�H㟇�� c/�$GK�nm��{�����<-��͜W0BAP�p�.o���g���~9�Uƨf�K�m�-��Uz0@�*��������l�1FEJ	�2�}W�7
Oo�غ�"N���"���k�h�l%���� *�e��<d��㈋��>J�ķv �^�������'�����;`G����h��v�݃�Jf'�h1y׬1�v�F�S�S�QZ��~j{b �6�=�@x#���a�y���YQL��{�_35�}N;��a��Cו�:"6գ���珤��j�2���>x����8��>�0��vRa.f8�(����5�vL��"���R!���E�!��%�(ظ�^	���ijJ��������?�\�A[�x�_���
eE�|^���m���@\*m�R�K��M�^i��ڵ��_כ;N`p\���������uUT��|��B�D��%4&q��8�[:!��F:y��3,��G����#DBr��!Ȏ���Q_!3�������Db�.�~U�a��cB��0Ȓ�����j�0wɋ�$��3~/%��E���m
�����y�jT"�X������ka�%��S���`iՏp��ݿ���.�n��c�t\�Jܢ@��2�܈ �Y��L ?��w���>|��	'�/�j��Z���B.��W����p�;:��gp�Xt`�v{0R.3��N��xA��5��%�4���A�|]�Z>@w�������t{$8}c�~����1��iJ�"%y���c�mj�*߄G7+��rS@���2���n�<x1����{��r�I#����>����:0�y�x��r�a�dj<�5l+[�k���d��%���$qߤվ�9��Z����7V"1��2�Ϫ���1ˢK�Չ]h5�A�X���Z0]�jz�ŧy԰+sR�?MO^|�۬H�������82�;K���*Y-�{��q:��X:$Z�sG����h �XBPɁ#)F-���K�����{����O;!������ ��D�,���>A��(�/[�K��V��g8�ƫl��A���	���	�����X��ۘ��������3���Z@��c��\�EQ�0¨���r��q���5Q�M�����e�z��Z�h�Q��V��X��Ŭ���0L<)�m��0�u��Q
?<2`z=6�(Ӌ���	��a4jVz���2�	l�>c�Ng�X�fW��^e" �pI�wGc���9giY�]����9R;�u#&�[�A}ϒ��P�#�����嗋ڟ��Ès�iQ��݋����2��<���v+=M�)F��y��=� �b��G�Ѵ�������9��u0k�w�n2���p �L�*&�i�P���(OH�܊�)�+��u���X<'rvyw�e���׫.b���,���;P�ۿ�!�S-�?s�I~e�=��3��4��n@��4������y���*�(�Vj�:�\�C�+T�_���\��@f�-�M��������~C�=�w�<ԏ �A{�d�Z����h��ɜ^<j���+V��<���A�D�����Y/Z�Jg=��QL�i��Z=����Z��c�ꔶ�l�-��)�ȶr�K�{��lg��cGɭT=���@�l�8�Ԑ���q�9��*EqU��%�G�����o!�l6t�Rl���f���Y�<n�� �1ᝰP�Ǭ��ik�b�c�q��f�~b��8=m+�E˃���[�!��6����P���j�^��d���>�m���N0�ٯ(]� ��Uva���}�}�����Ӿ\:|�	�r��Z�����Ax�Ù���0�c��9�%qbҠ�S;d�ܟ7]��v��|�ћ�@���;�@MS���Wa���c��-�ۘr�}��p�7�"DB���3�:��D_`�c-�� � \�X�ea���O�^6ޏ򚍃�ݴrԌ�@D~��H������.��Cq��\�nu{��(y���r��J��c�l�����8�B��;�`��ړEgm�P`�z���K�i8W^�u)x��bҡ�
O�0H�P����L�?ph�}�oX�D���|
��i�+�7�FI��#UOuX�K�u�J�� h{�J�/�m� ��x"���C��M�7���¹�?R]p)�J0Vw ��}�n���'�)�3%��������0v�_Fb^F��i�2\&��-`��!��{Hu�L*<���lI�-5EX��<�
�:60SSo�������v\)Gg}�}�jX{�>����[I��e9�>vܦJ�4���W�e��@cF(	󙅽�s���xD3U5#aE�kw��0*��NϦ8Eu0&��9� iϰ����������U0���b�ʦb�	�zO|Ws�6E78[='PM���1�c]�,Z�Ή�=�9�R�:�?�D�Z�����]�x)�8���	u�����{�{��p�G̟uéd~!�Ra'�!�	�	p�劀�h*1ze�>���V�n�Վ3[�<�ֹK�Q�]u��)�|.�=6���;ֱ��I�XI�B	D�vn��l4g�0��{*�>�C�����'�	0q����S&�y�!*��C�NL�u��| b�o}}cs3B�k�#�-�a�ݢ����aW�9V;c�/�4o}n�@78g�����
�.�*��_����m�̘s�èw�6���Qÿ"�ί�Lm��1��O�Qs'��Q}i};�9�!�2�t_��&�֜y{!���A#^� tXf?�^ �=H�j�-��xN��ƼV�r��o�^C �o�[@k�����d0XqK����l����7�JK'��_5Z��I��?�N;���&�/�U�\�[~"��&xcÑ�~ðfǜGF��H�'��ok����6v�j(۴Z��rh����b7�<|s���#��mn ����p��҇��\Bނ"@���A�3�� ��@�Z�׶&�Tx}�̒�E_z⃨����I�}Q6p����H��F�����VM�ͺ�f���eS�hz�'��m��sRqT�c���Kڝ{�3�p�tR��Yi G~�!�A$������7 ��B1�~��~./�H�;k���-s<�$Z���kDnHo��H�'�H�-���k���

�x@
�<�苯��Q����	v����;��:Y�������'��U���n(��~��]3�!tv(�L��괓���������	�΄İ�!G�;�G�)WP�R��.�K2�Ͽ_GW�lD���B妮�2f��	I}
���`F�=���r:��x��w=������u����l���!�K������	P[U��J,<�r���Q�=5}n�L�u
h��|�;��=t���i���z�z�n�TG����x��a���^��ce(��{�iN��ʌڪQ_�G�uƱ4qIqy�i�8)����&�9��
xx�IC�`ό���`��ڏL�}Uݒ�Q�}Ƶ�4�������xK�͋[ ^h��
��D�ޥW�;����8�O���G�uLV:UB�'��4��c4�G\B(��q� Us���
�����o�� <�`�	:�$zb�H�76x�f�g��v����&�]��w�m=��騾��ӈ�_�é�(����[�|Of��A���]��\oR.�S6-�7%Y�õ[�[������C��4DS����^	qXDcՖ>��-��x�(�-������x�扢Gf�
FN�`�`�����ہ*ǵw��Z��|C�2ˊ��$�e��Ҙ�I���.L�����?_/s��8�D��}{�D��E�b�������.<|/F]_�D]Z,�H!���+4�A�/�h�x��g�^G|�|�P�g�D#������D �C��9��y��7F�u�iJT� k����4a`x�i@͖D;o�]�g��1)֞�S�\��u,U̧�i��k���AZ�Qy]rT�?�.R�,��M] c�J4�I^6�Y_��U��z9��w������D���1�l�٨F�0����WԒ���?	7	�ȫUЦ�V�t��Uj�	�Y����B$ĸӭ%�	V�[���L��,|�5z2�=?��;�$�ܗ�\�6��kݘN0�5-ڧ=:ߗa�Cۓ�f{m��A�	��o�oO��k�~�t���!��:-���v3�������~���M+���:~����	'r�0\��y�5 R��o0��zҋ|�� ��7mcAw\g�[���=�8v_(�b\K<o6�>��e`X'�Z�M�,j�1�4��_^�� ��H��d����TcW�,VIn���o#�}�������E�!)F���5��E�%R;��}�HW��:��Pyg�������5�!�`�R2	2��Xe�Ŭ7>9�-�mMA�GG�T�Ufa����������CM��=�z'��� g�'�T,�2jWt2h-.Ї߱U
�2~�w*m7�*GPq�� 	��(�d�Ë'�Ou�jt6c:� ��b��A4BZ\a܀���!�1��p[�E��	�	�iF�;�n˞�~ԑU����h&�1�F1<FICoTH�+�ː읣Q?ċ����꩙����v🹇�j����&�;�ǅ�����̀�����8����m.�&��L�-�o�.�}�-�+#Z��� �|��
Q���ۍ��<[v��#�Y���05ב�״�`.�%�?8��Y����Z����lU8@�"O�vH�є�qO��s�z,=>KO�uP�L��E�Ŀ�K�,E���#	=��H�.$rB��Q��BW���Y9���d�����cG�+4˭�@��v3��<�ý��D@��p��d��aP&��Sd�=��ya:�o4�A*����a�%E�%Gb�Q|>FVµ�4�އ:����L@�� S���a#$�:y�oX��/�����v}�?R��(K9���E�g{��$M��!�������ν�N�h�X���b�V[��=� �ݍ.�Ԛ��'�0��	Z/@�N)��s��!�ds��k`hD�b01<��1Vj;�����Iҽ7PM׎ʃ�b������C�6
���ɦ#���~�"1�/��&Ԝ��ŗ�g�����|?W�������}���Dg��V�) 3,�L�m/���,��D�j���Nq]^��z0_���unXbs>�S7�ɓ@�Q�:[)��l9^�	!��S�k�{�*������ �EU	��lh�V(�]��w�ɐ�e���i}<Q3#3�bI�����ץ��������192�
��Da��·k����!�d�� �>&��^�v���J�fo�� �4��#F����Λq"c�~n��`Z��u�3����=�+���攼����L��9?J>qAܤ��ll��Gh�yY3�����5s+������*��RAda���Mg01�E`
�cߌbv�]@]�i�_�2��@u��-D��a�U_r!���
��Й�����VLO���y�Q�[-7=R�18i]�MH �}��a�Ą��4�q�K���$mCc�9��.�Ӟ������d�<���\��K��G��[A�y��w�˞`�qxP�$e��N����fx|�E�!nij(��tz�Y��
��ކ�U�F �+��MP��'B��C!��6������fI�����0��@~���n2Ǔt�JSO���%^?����?4O΍:�;����/�"8��}Aȥ3�d�QL�舖�X�e���������ן��6�����sd8p�7��S�Y�nϨ�D&J��+�;�ʏ� {���%��B�5"a�/��i!����Yf	�E������h%�v��Z����n�����Xd����&�C �q��Ҫ�"g�R���t/����F�,;m�M���I�B��>L���ٰ�ƻ�����e4忩^5������oa���#��Y����O�5)f.�����`̅��G�w��Q��uW�g�Ҙ�P�/�޹8��=B��>G�kc 餪��}I����w��W�k�����ؗ�8�uRO T>oNs��t���j9媏󣂩�w�]���_C����nIHR�&�h^_��H	}̬�4�0�����.�N�U��"V��$���_��x�6݇��{����ܾ<X_�)E�S��脨v��:�F9��s�֛x�o��ƻ�|�$w$צ^'�!�&^\^���G�/��;@h��`FI�2)(��7�Wj��\� =�LL��E�_�e��5���D�t���$����,?�Π7����PϤ�����OkO�Y��Xy��S*U+0�&����_Mj	0�{!<��78�^aĮ:k"��*���\{	O�3�������d9w�\ٌb�����	S���@�4n��C-��*сCZK֦�&7h�-���E<Rօ�m;�S�� �f�I�v�X-:Y�N��A�H�(��b]͏�����~K�K+�}#��
�����o{�ne�n�80�㼕�E��_�y�R�\��-o����K�ɜIs�N��yb�R1(�L�3��4�Bﾬ��;��u#Q�ĪIE�����f�r����ҮK�p4u`U{�	�K>x]��_.�u93��B6����+�n�&��(3�G����["�ї���6��r�j�&��C*4Q���)�X	u�+Fy_2�N�R��r �A5���1D��E���+���D�,���k�:"N�����4)��� �������6Vƅ����.SwB������`d`m�\ą�}�T?����*8��-线�l+�;�u�����Ky�/�[}�
�'�IG@UоAh2���u	���r�'�0A-�ؐ[�t��°B��,R���UN<��cje࡫d�?
`*o���o���ܚj1"-�i�~�#��rg��S�x�D�++������,q�n���Z��3�w�ė�W
)~�	2
ZYQ9u/'I�T���]r�[4�k�9��|�okI�PacM��=jX����ZȊ��6sxk����:�l8�M�AB�2�Q�#(�p��RL��F��t����;�%	�C�D�蘳�ls�r�qcj lD�6� ���dB6M�B��;��Hi�B�qqϛw�gg��A�PT��`7����^^;ؽ	�}Bm�7�����3k��yj�n����e#��hQ��/J|��n-?�NP�h�p+r��8c���ĕ7k�?J愂׊
�����~WjX�.��`��ʦ6J���e�-ЊU�"$&]w������|�RP���r�b�DΠLS�d]��-���lS
��Lb���J��iN����[hP��P����	��쥄�fV�U� J�Γ�4K�ۜk$ĝ�ց�����v:�:�cw�����@6W���N���e�`�KǈƜ<C�ς�Q����!����sGD���)y� ؒ�YKa�d�X�N$	x��?�1��������&�z��Y{/Wb�
&ue6����߼�Ъc�O�����F@#{��apC�~*���V�]�}R1�����F�hNV�JL�w<�����w�(	�H7j7%�չ���bJ���s$u[���*q+k�;_���Z��s>���TK�2�������|��/����_���Sv���p�2�a$ًr�#�ju1-��c�CL�!S�bHr�_��
�y��	�v�W��u��Bɷ��+��U@v(5�S�޹�T|ݠ�X-�4�
�R��V�Ϭ�����OeLUI�I�,��]{��]�Q	��4Ђ�����0�h��!���{��ܴλ�C��.���y�9���c3CD�z��W��R�b���8�7�"��B�L�/Ox�&��5/@�rłw�ف\�ȓ��A�G�LD��$��5��v׍���]DH&�M�)��rq9�lĄ�ib��tୖf��/h���gs8B�'�俲��bϢ�h	��{t�#㖛�ԂL�Ps�!�(0TZ��)e�%3�J��Z��q�G�<��f7��X{����m&]O�%�)�5� ��]qD���ecF��>փ�(a?�=��	mq��>-�V����%خ~ ���_{1�f��ڐ������%B4o�L���a'�Ҍ{���.F�̿�ɿ~�����m�(պ��4��و�#��V�@���>i����Ą)�b��������Qv%��Z=�Sn˩Pӱ���yx��	��cծOo�3���%c)v�Dǟ����Q�=eIѥ��g�B�ۧV'�-)g���!�&�,v��ax��xp�<Nı�?�	DԃP���F�a���.?��Wk��z�2:�|B�r�⅐~��n���7�}��Jϭ\����-
g��6��@�*깊-��A6X�U�?$ nת�)�V�Z�iB�I��Ot�v��f�|8�q�+/.�[���+5�
����0T�l�l��*��N7~�?*ʬ�u���;��0-?��|�qP����杊��ji!o����a��_׏U��p���d�o6�� �*�E�{�e��gRȂ�Ǜ�����W�wڹ�JE��U�X�j��k��L�QY��iqq��/�x�m�H�d%%�Tv�a<T���M�?�`Ǜ��ck�:���8P	��8�$=���h�a�u���<ڣ0�z����t�*7J�������=��S��jw��X���T�>�O��Om$$y$�\~J�j��Cip��ea�.$ݘ8��BӪ��h=���3�L{ˆ��B*)���J�.�2�=�}���R��)�>�����]�fC�c4�'�hy���߇�o1u(O�)�1�J���{��ʮ��R�G�U,�Fz�l6Q��5	b���YY�*���_������)gM_h|%�̌�'I*U}G�<��;�4^j��+�F\�6&�����jj)_&mۂ�;���"q#�=@Q�6�{	E��jZ�4ol�l�2g'	�d�����ă]l�Ø�e�|��������(�+�w�c��t|��4	��]�b�+]��|��p�^�3K@��ܸ�B�HB���	+n1�����°9f�K���M2h�f�<h/�a��TO��&���n�I�d8��=�|��>�m�ixm���ѓ�?V���5b����sB����VF��7�����:�0�\5,;l���M�Ǎ�0�e�G�G �U]EV�5�Q^��T毚�Ѥ�i#|ѡLZ�u�Pʊ��e�כ�d&�H}�|wJ����̳u B�Nl�B�|;UN	������kÙ�g���d�S͔Y�v��a5L��G�����Ro�x\��/��G/g�wM-[�8��M��53�Ԥ �	��/�ڎ�Rb���<��M�%��}m�k^�n����Mv�������g���<8v�	�N �wĎ���՘�[���&t�
�xE1p��UyP2���"ɪR����O��BM|�~�z״��G�����|T�P<�-k��WA����'NҢ�!~"�^U�ی�f(Ε2���ۖ�������h����P7����9-ښ*>��@���a���[<O�%�e�]����O,���A����0=�9��,�%|����O�׬���fM��D�5�����1,Λ&K��a���B&�w�F���"��`oq�P���:�o͞z�Hc����ś9���K�?3��=���KoN4���'�fi�ʀ����r�@�v����5aKP�Y�>���m_|���U+��.֌�m�������|�-��
ٺ6�J�Cf"�NQK�!�*�\3��o�ìn�=�����q�Ю��z����vqHIs)�����[b��q���"��d���2Q#�����(>�ؑ�L�^�"�U8�+�M�i��P[�%6�}ƫ3�u۲�H�]��8�ʘ��� ���Ѕ>��ܶ��$��qS��x��6��	���ϐ�`����|%̶b%���z��W�L�'�]y�����!K_9�,��f�3�QU Ifq�*&o�#�q�4��Qg�'�,]<	��2FۣI��y�����p�kLz��C����.C4�o�b�d+
*jvCo�l�q(�/�S;�bN��Ő�_�~����7�1f��@��\��f���)S ������ѼҤ�nlV�"3��pp���0�Ru����z&��e����}�H��Ջ(J�о�=� ���AQ�,,���ySUXѣ����[ �����4����Ą6�E��D�P8k�޶pW-��K����� �OL���N��u}�2�ʭ �u�֌|�qO�w:S�n?z.JVg{H���s�IN��)�"O�#�0��i���;1&��9f����u���w?8�߁)2�TfT�%}��?fz#�3�s��k%�� I߰���� ad	y�[�K�
�9��5��t�@��8��oէ,]�n��;2�c����+w��2�
1�Be�Ki> �~z������AAU�z)򨅻59�_�� ����\�ݞ�ӂ�,����fۄ��.U�2����Y���]&�`hJ�q~3gc#o��a7�-/�ݼPh����Fh��%d�^���f5��®��5�e�Nq�Q��_8��Bs�Q��y$i	�S�p��kj�lj�'�oa}|�����$���L<�	�|B�<�������S}ت'ǉ\�u�~�&��H��a"�"�p�>�ӞT�7q����u0O [�����Z3z��`UyPvja<�t�?�-p����f��j&��*!E.,�",�H��������p���y}������9^=�l�e�;s!�Z������F�w�<��c�Ր�;����O�v�K�F4�*	��0R�������l�@-�W�J�ut��ts�vq��۝�|��T�L]EY��O^��aDܮ�e�
Ʋ����ˡy,.ȼ�4F5rޝM�}ê��ĵaBGd��1ՠ��"̅`,m��|`�6b�m:Nk!��<y��H��Q>�H���5������|�-,�M�"$����)?R��y��g�s�����қd�[����;��M�%աEM�vQV �Td��Pg�嶋h�5����&Q��N|S)��U�ƫb5�%��Pq�-,���M��'n�Ƴ��SNY�8/��	4�/�ƅ���M#��s�ǀNsH~���,�鶦n�d��3��w��q��~)|A�"r�y�������e2g^֚�wݭa ��Z��ޝ6�Ǣ�RN>,t. bD� (���#�RES׉B������$�cE�T��u��� 'U�����͞�
w��eB�*k1`�c�}�P^��9f=�t�.���fy]*_35(���Y#���N[�-5�^�?�����-Y78|N�w�`���Y��䡘0z`�� ���4ʋ�x	��h�.Q�6�6qp:����U�E�&>��n�ɞ����,���%U��e��yj M<���о�];H���{��ͧ4o�f�@C�L�4fN8��@�#��7(=e?���QJ�
2`���4�o�I�ϩ��rVuCw)�؇��U������y憑�N%�jӲ���6&G�;M�����b-8v"��=���� ix�
lL� g�%�^���|VŔ�=��Q��j.��Fj>茤�� ��>�͘���&�k%~EZ�j��c�u����ы�K�v o:�7�"j)���ղ[i�K)�,"������|�J���H�_�l���o������(~����d`�a�d��.�lK�k���X*\i�� uy���l#.%�h�\�L��l��1����Έ)DZ�A�r��{�l*��[uDRmCTX�t9ͩ��e�ٻ@p�>�������찕�c�21���^_[
Ê����d{���m�j����sv�$Q��魅�'F>(�ΒD����9ৠ�!��{]�JlC&�uj<�����Q�dF��/��v ���f��%L�J3�GTu����7Uo�v$���[�Y��\�5��d+U�ˣ�KR��օU�%���H�����#`]b�����H(�'��?����_nm�3���#���\3p�E� �/�3ԩ�|k�R����P�s_^�BZ�� ����t�aC�30܉��h85r�,v���9��3�'��f6J��~��(��18�r�#�����|�`��̄��q���e����2���UQڙ��Sm�KNUXh,���ݚ���^��ƪ"aZŻ���dxU���V�MK-E�ۦ���D�,��vYH���P4ݻ�F�x�>�g�aD��#n(	�I��#� �Ylì��A�����y��qd��O�*�K5�A{�Gj�aШ��}��c��z����ij�{��(:�қ�ǣY��kj6+\�j��m0�������� ��8V�Ąɤ����z?��e`�K�~BK��	�B��#��M�X ����'0ߡ!�Ą_S�}������]�h˯*[�q�~#<�k^�n�i�]�x���\8ԭ�9�@������\���g��mIAArm�4yO��D+�h����ng�o��PVK����%X�͇�A��@�p�0��*v�h@׈����D<f2;W6��^K�!�b�i�E��)#���ؐ^���F<9��r��=��5YU?P�uhg^��� ����nnM(����Ia��_��T�t��P-�v���G��!���b2ⶑ���QbZ%�������9�5x/��U�i,}�v㿫�s;�� �rI��,1l���҄eW����Y��5�*}Tmz��uMH�<��(�xfP��v�H��|:��n2��눙I+jF|?��#k���{�į4���.���m�T\B��Q����s�B������d��
�!7�������[������I�A�灵5�7>K-2��p�J�2$�����Cߞ�-g�=`�#bx+��ߏ���f��h������cPC>�n+�E�m�פm���O5A��{�tҖ��uXm1m0�}?-��-��v��L�`晴��O_-]�����O��샅��_:�����z+R�Q|�$#,o_B���[�$�|��u�9�.357�͇7��.1c/��ac���E�x�b�ݑ����Kѡ�PbB����/�$�v���#��E�C�Jy���5H�c<�Aݴ~׮��wN�y�vM�ⅾN9d#�^U�6$m�����6sVQ���q����x�����W�Zn�N�4�KXcw�2U^(��u�mU�=^A�]�-��ʊ�~�d$2�� ��
#��Q�l�����de_�H���$ ݥu~�+��P�:|�����p@�(K�2|̣VF�}�t��R&x�D�13���:��M֔9]	�JʖZ�$_J�AY���9J=��e�6	E� ���Dڈ�AMAr�*�r�3�{65/�Z;7��HT���)�{W���\�ƻ�1�=���wE�ɭ�HٟU�H�Y�.z��>�����$h����G��5>��Ti߀��i5#���t���7m�=s/dc:�x�GwF��jj��Q,�@Io:���f��� >'!��~����\�����1W�@Ȇ�~dGl����C2�>�r��A����`k�;��������Z3{`���x���5h���:�M� �\r�9�$9�V����umװ����vX@�I��7#P�g9��#/�b��9�2ూ:Cw�(x��Cb=}<\��
Ӈ�Rێ�j'��0!(��C<��m�`�+��nv[4g�![�}�©��}d��%I�A@���,�wSJ��9�5:c&�>˺�8���G����_����_�o���Ⱦf{;��e�>P�uJ����'�k&�8���3��Ph�/��F����	���w��qՀ�͝�A�
P��{�h���C��	�XR�E�6\�*�]� ���cBNB)�Q^�6]F7�Ƒ+R�2�D��<f��������0�bִ��u��_l�!����*z��b.b�K|�Ү��n�>�;�~�-1H>N.:q>����<�P���8?T�޸��S˜����r	L�u��OC]�":�s@@S��Y�(¶�d�W,��~�D�̭��!B��vv�Qߓzx3�G�jBq0Fv�c2�3'2%߯=M��Y|~ ���Q�D�k��16|�M��
!2n��^�?C�~����7�������L.�	���b�'q�W6��P�	�g��~�dѹ#�-��ֺG D�5.R���Ab�V�M���%W	���W-�܋��+�Kye:q5f�|�Xsp���-l��ԎS��O�[V6��nS8�w�HE�77��q�_G[º��0#$��@O��.P3�ƚ�(�>�vژy�=�w-➹h��p��g������݆�KRƟQF0�uhD��3��a˽�Ȯ���~��(���j�v��N��7�l�uZ|4,4�$fP^C
V�~������K�%L}�**�Az�&�ȇ��<G&觞�Ch�?����^b--�U<�8*��t���]���]��`N��;�ߋ�&Cl���F��B,M.P�#?d�z5
�'G&*b��͛S�v``��s`r����g.w�s�k�^M],����(� J��Tk���B:܇c���`�C%�����3@?��*�O�����/w+�����k[�#T�'�#����������v��1�>ѝ��c�u�}�f���=���3���)	`����F�޵���f�MZ�����N���/�^����?�;1n?���^^���>ě���]o;i)8'��N�E+���ޕo��x|�r�$�#|~���nh�?�$;����ߌ��M��9�S�=lm�n�=��ү�Dげ�~|_{e̦�Ew�7)��# �b�%a�|�~R-�v�_|��`-��s���
�D���<��Q�����3�H�o��X�=}���'��xF��+�v8)���j]�����9����|���7�]�O��FK�B����f�~u�_��%�����0�%���e�p���r�;k��hk�.!��guʎ�恗���!����$z�Ax醸ۀ�Nڊ���5>�qs�[�ʲ�.��H�_I�n9��)��7o��Ƽ�zoJ�g�A��ѫ,����;��p�غSKq!��5�t���E�-�������[�w�'�X�)���x;̉�t��Կ���\!ye���,������C=���nZ�M�"|�7��N(L�@��+�J�5��"��g:Z���ĭ����G��ܛ���>f��U�X)��py��j�j�M�(l�����+*FU�]�?��@��ǉPK�O��/���E�S����V�J�:�w2OS�k����3(�sx�<�eqѧ/C��ׁ�q��d
"���r�^�5,�9e�B��/|G��ֆ�\�c�CZD�+��03+<,���V7�fAʕa���E���p%��meW�d��ڇ��헅�'�X5n�|t"�R� �u��x���?�=Y(�[X,�.��H��5����K��L%�e��w��wA���	LD���[�������[a���H�pPQ�v�,,"�ZZG,!f�[�mPa�\��ࣁՇЧ>: \d��>L�����7��VH��P@��i��B�)��o��;�	e���<���p,ܣ,B>��P��ɓ 	����W^��[t/�2�n�T������(BҢ�Cy�K<>.��0멯K餡��96/�g��<#+��(j����r�&3���/�"��v�s��ΥOdٖbrqH�KjNp���Dأ<���O=�ᢤS�%6��Drm)T'x��c�Y�>+A`j5鐨�r'��	 �����Z���]��H5V]E��x��'+��U��G��M���) ��bH�cx�a2��U%@]�g����C�%��9�e�+�Gx ��42O��߼�8�_�{��C��[��g�G0<9 �|��Q��d�fkؿ �"��i��E��G��$�l[���A#�#��U}?�{���N���3�����`I��;��~My��Vx�Vk�tx�D��tdlK�@��r	�?�3-��R#�Ov��_5]#�Cݛ˴���JDb���Ͳ]V�K߆�Q!M9����)akX��`��&�_�ʥj�q�X`M���d�@����@�?^���5�#�oR�[AMQZƽ��4�ie��_ΰ�����ˇ�8+N��CYj�}��Eؿ���l�����>ƾ��Ŏ��rۂz�Zo'��I��>B�F�م�����9��%HP�el��}>u��u��Kz�a��9^�Ƅ����Ѿ��Υ�k���+��E�]
釔7��n���RD�_�4��Ց'��&z�6^���d1��Q�3��J��KS�w�+�H9C��Z??�	O%�j��Oۄ+>�U%�G%(�o2��(<���s���+�J�W�zx�-o�tV'��ׯ�
��l�׏g��+��1��ff��y�i���C�U2N 4�����X؍G����M�3Z,w �=0A�|;���
蛀�غJ�ϕТZS�CW���^ɲ�$˃p���1j�z<tV�8�h#�t�����Bѯ��߽�y��f�y\�x�ҏ��]H��>�@r
�28y�j⧉L/'�M��f�t����˪��gF��Ǯ����P��?n���}��� �<��ٚ"<�'��oCT����G$�
��$^��M���f�ĹU��&��Ŀ8�4-h�.R���JR�>���suc���o�[�:m�W.#}Z�����׆�z<qz�M
�~�y��)���q�d�In{��o3$�Ph�=R�f�sAF>���p����|��"�kZ����V����K_�%���� �>T��AB`d�ZD�J���pS��+�p9�2��X�� ms�1��D%����c�|?�V����MP���pZw��=i�_	�K,�J9�;����i��!g-d<q���nu�&�se�̈o��L�B�8�y+���9���-z��|όS�?�fM��,�`Y�|�X����v����G�Lu**=^�ᨭtN�֫�<J�Ҟ!��L�B!�OtJ`a���z�'ˉ������ߙ?�Z�э�W7n�v���KP��b�/|ִ �7��(=[H�U�{ ��B"�؝�:F�3nF��-��<���y�x�c6`஍�渖�b0�H���к��+IHmΕ��C�':�%N��u��X��*\�oN����dr�a�L�U��tg��|�����I�x%�4�B�\�x��%N��MkH{籧����~�����Q�F_���:�rz�rqLG���'� iY���&D��㌾Yw��Xn�,�-C�U1���A�O}c$rr��b}�@V-�M~���"H?�ܸ�r�.irD�aF{��Ű�?���>t��u��v�MA���J��J%��	�?�Cd�%�[��<(�$+�����"L��,q��iY�I}=�I�=s66�3����_���K��R��W3ii?o �'����`'/�^�a�I�]�RB����Fo5��5c�����_��\�&�}O�m�������F�m~(D6�T��������ϬHz�e/j�Ʈk���!HZ齮�z���De�kqA�X%��DZ/�u��Y��e�l
ծ��F�*����=���9[7�� z5��H�焫з�������k��j�� OyK��*��H*�e���r]�Dg1�p3>��K+�z������,Y��'�$�ؒFɰ�R�_����'���L.]�Ί/S�m�j���"��ac?!�1?[�J����T)/J�ʁ8B�$64�j��ud�k�Mߥ�*���~-��v���Xa��ޣ�y��H4��������{��b�i��Z7z/t\��N�M���n�	�!���<��D�Q\�u���/~�Q�Tgz�	4k~U~��/k�uQ�R��A�,�?O���N�ENQ���s�x�A��( j��1��4�F�$�q&��n'M2�*K]#*��_m@���!�~�o��biw�0��F�svI�cYD..�9:�nR�ou�[�c6�����6���*8�3�EsT�sEV���ƖRK�8�,���5���9l}��|Zw���$U�R�b���T1��G㑬�}$&X������tI�&�'��4ͤ�*2a�]��!� ��b`( �=JY s#�T�NN˶d�T�����,����5��H!��mw�ݺ:�Ӕ��9��6��>�lv˻�J�o�Btl��oJK�l��׸��a����oNw�H�^��G�u��2%�$@�Q�/~�o������,rs�/������kJǰe�a�j95�$��]!���-�K�������u�HJ�+'�<���ȼ~ދ�>v
Ԏ闔���ӄ���a?B�����B  ٔ��s��HV�?�t��BҴ�@]:���>!#�)��1Y�\�b����c�!��lM�֚�=�mQ�"�O�}�>�[=*cޞ	�_Q��?�"�F��e�ɀoϼ<���������Fn�m����<�<��f�Ή�r�G������3�}�7!�m+'�u��ͪp��
��=�>��v�]��<�'���x��>�;�m�� �6���=\�Y.h �%¼�o�'�����>#G�uJ�̙�&�'cCD�R��O�ͯ)����Ѫ���0޼�H�sDs՟k���m���Do��^� cL���(�r��>�~�����}w(��>R�_=��'�-��f�B�R�Q�Y�lqY<\r��I,��[�9�}��b�H�7w
����f���:>�*��\HtBh�f�%S�e��&��̕�~n7Ra�	�X�N��64���bW�����*?=T]���#�舀zn�?>��.�-�d9�Q���� �;sf�~h*��ƕ�9��K����;�
��*�z#&n|j���ծ<�.d�s6[m�f�j���f����E4%����H^?���	��L����"���G����J��NZN�Kxw��_	��;n�Ƞ%mfW��;��>�J����-����dhf�[@q1oǹq�辁��H�i@�A��0mJz��A�P�'�*O��������Р��ەMg?��W�@l0e\IH��Wwp��/���:Ah��$F��lv�:q7��i�D �,�v'��q�%Ѐ�3�ͅ\�]쵿"sr*���/5�3
#H�8���b��/Y#�/�Ҩ��͜����[~����/d���q #R I��ټV*G�$v�V�.�C�3���Ur_�2� \Լ��rCd1�J�lz.��d�<_Ը(��A�)��1go��vD\��;|�K,g�N�La�!�'��*J�R���bI�z�V7��prF4�9T��ҭ�a�����Y�6��wT�C�ו^����M�V�
��v~�^��� �ؤjR1����5����	��q�J��G)z���!CT`�fs���줹�UԀ;5��cZ�P���,~H\3� [��'葳4�Y�y�>��wL2��J�[u��PE{`��8���,;��w�ԥ��d�lB#2��R�'0�X�2@\��D�v΍b�  ���Vq���U@��T`�C�J�����g��qa��zK{~���G��D���Qq�+U�ɎM�Y$^M�S&c'���6 ��"k-�I����Z�ض?9�J׹��}�ܾ?�Y"w�b�-k,#� �I�����XgL��Q���K��"��!ia��jM1�?�n���V�� �1Ko�|$|�0`L��̤��O��K��t�߸)q���S'����G���Ǫ���5,sz� @\�&z�Ŧ�J�[���8���Gd�t��#�hY\�Zq��A>���C(��hq��E�w��:���T0�q9��z� ��:�彪u�&���qM�G���$�˲@ɵ�g��~��b�ީ�=
��o��;������9�2�q��m�2ε#�E���5���h`����c��Y]��2Af���!
���V�Q�T����S�z�<���<-`��ͧd4�K.���4���.\h�S8W,��W,�d�Hk����e���ushj��}�Z�+��G0�)���s�_��|k3���'��(7S#Hu� �+�^S��w��;0� ��2l�� �Y#l2��n�̖���S��Fq�q��t.���Z�p�������O�R��zV�P�flٵ������=�7UO~I82_Lvㆯ�Y$�D�{k�H���U�b�H�ً��p^n]1+�g��6�>7��1J$]J��̢� ���v�\�ۛ���]��co:�h��\U�rE����%�Ѿ�֝���m%�V�t��wj�,�K���s�'Gw:��y���=_���-\��Pb�p"7�V@K��cD�WO��o�c��v����:Z�^�B��0b�����+.��P���W���'-�Lv��� �8�CE���Wn�/��_�߽H;���5��7���6����Y���,���M&�7�p�'GU��q��6�H��R�$����M�M�Lg��x�ơ<��s(Uw�v#�)��9�F�負wSҁ8�����'�ՆXU9�h?iY]p�n�����(�'���`(�g�BC��� �sd��,�@V��i@����5�i���<���Ug�҈� kت�T���]�Ee@" �z�N��4GjB��_�4�l�I������h:����jB"|�"�tt��L�8tt��κX��%7���F�_y�X9en�1Hu	����|re��/x3є'�~���1��c�R�9�Mq�^���a�����1"�g���P$I���):_���7Έ̈Ft��pk��w9@���E�62�����1���L�jLշ��{a�L��X����"�$���c� T��+�c�Gx�� qE�K�;�i�G�s[���`ڼ��i�<D{+���i��{Xg��Q��1��8�;����{���_{�h7���t���I/�Be8��s����[�wߎ�Ug "g;�m�ԸnRJc�U�&V��l�B+�NW�� bVw\���.+�q�b�8�&�����n�j��~��{:1/��V6�J'��9#��ב�"��&�!�W�\�S+qP|��a�s1ְ�(Fq��R
k;����͠��[�-��U�-J\BN-�~�2�i�A�e<�F7�i�H��8(:xs����}E���Tot|,��/q5�WF�E�w��z�L��l���=�\�������+�0"�)�yK��-�������&��=�QZ��2�Gm��_46m����zr���a���!�J���Ny�7�oyӘAV�w�^�����ި��M��ײ�i?v��Ӕ��m)ʫ�y��N���z�<���w���Pk����D�ĭ�X�!S�f}����w�1�>ɪjb��՘-8��m�j�Q`����������Ã��t��M���B���b�*�l����c�E8D-ǫ�Nw&*"0�u�O��S	���k�-]��\�9�G�e�0π�2D|���	c!�|Y#�³�����R���ݜCT��P���][���*�Y�x�N(.�Jo3V�1��H�a��395���Cd��s��gݬl�����q���6��B#C]5;.�64��]�r��R�ɹ�=�ikfR��pxL��⯼g@���TV�Ҧi�÷&v��yd�}�,�bx�D=f�g�l��2� ��1kϫ�`�Y��V��H�zD_R�?	e:~�A��,A�4��_:!� �����N{�`���[Ev:�^ܾ�:)�N���C�y�DF�Q-��{8��6�E�楔"]s���iq���#ڄ�X�M�A���έ�ҍB�!�dW~����4 �����vɒ[Y�]�j!���o���ڈ�ϭ>/HBl�5ܱ���OI�A'l�O_��y
<k�p.1�hv�$K��i��o`��6���=\�z@�e��]�����k���&����	G��Vٖf��W`⛺���x�O�m-:'��$����<H��t�m �E�L�^nt9��5����O<��J&�I-}Lt8��铱,1$ W�.�MN��m���5"���J<�lR}#9=^��c�Z]}���,��k��&�p�Yb"*�����>*H��t�'�ì�LmwC���u��KP��0Qs�e?�ϳ Q�G��5�b��?��§^�yA��I�s<c���.�"��v�(��T^ɤ�(/���"R��S:�֢!~�S��p����9U0Yc��Gw�:����&X O����$����w������?�t������T�����8�]b6��SH�����A�K	����F���q��%׮��\�\�u!�/�X<��,��z��ao���eܾ���p�@�]88��8�q9��#�h#@�Q<����^`Q��{�}Jc2��nn�;�+�_A���[�r}#;@.X�:S��M VW��-p�\q�M����q� �
�n��n��{X�U��`�� �5"�:m鿼Fc��q:��Ħ��]�z�����̨��6��������8�&�v&�#/�U!UO�����?-��Ql�>O�1�r�$9�w;&�9g�/M�yo�!.B=.t|���S5���}rM����,�yy@w�D}���J�ѯU��s2��K�x���X���\6����e��:f�?���@�#K�� {�WL��4i�Ҭ���G���0޻ ��8����m����J/���|�V���_���њ��V\���#� �PAw6T�ﱤQ��y2�כ�zX�H��?�|Y~::0��JF���9��������?����/M۾t�j��Z��t/b���keױ�p�������䡿�����ϐf���գ�b�u�J~�g7B����5�5ִ!�q`�3��m7�'�M��(E����f�`l������ B�])&vT��
���:H�E�Ov=�wQMb�S�� j�0��U�g���f6TH�¼��+,x���;�(a)>6Aܠר_Q9Yठ�~�*��YBG�.��zRb����7�4�jL�fWU�d#r~�ފ�����w�MW��&0�:����Z�PT V�G��:9��w��u����b��l���������ڏ�%H�)��d��Y���NFRMg�(C�8�|�{�i����� ?&/��`��A����{��:�\����u���ⴋ�b=���TX�ϙg�-j[�qlHȯy2�j�<XSO�e�W�T����8�	�����D�<�T�:/��+�I��7.��QN6<�4��G��)'���7����ћ�p�BQi�[+pJ.�a:Z@gqdb{��{���"vjo�\�h��F��=W[�����:�L��mEe��2SZ�����lC����4AD���#g��/��"^��涧oJ�p@:l�cm�D����Pb�/�a�+�Jp���l1ET�1�߱2�^��Ѧ��K���Ұ�N�Ryo�����o�N�n��d��1�>�����fV0V��DBn�z��b��XE�B�H�fu]~��K�V
�1/@-1���G��e�	���wPL`vB�U�YJ��*1r��~w�Pb逥�T�nk�͍�_e��j��(fJc�bV#Y�J�~�TH�Y��&���o�p��z����u�c�Z��
�f�T�e�2�]��#��l���ԥP���{m���e'm~H����{�y~@Y,�?柠��R�þ�I����W�ʴ�WC4Te���Ȳ���w2�>�Ö+9�ȵ[!o�5�י��x�M#�Ir=A��xY��\�*ۯ)|t��p�*�V3���`�
w��Gxp!�Z!�_a�,����''57L���~g�`U��d�U	k	h���.��z0fp�W�I���r�pj�y�����50���Oͥ�r�o
�"����w�?pz����WŌ������|'��#������������t�F���:�Y�[���X�k�甥�Z�K�]� ��N�IO���"م�)�I���8�5��4E��Ɵ�d!w�n�d�Q６:#�9�H|�6Ba,��N��|���V�xQ&Bo0��r̔o�;fWg�:G�9�$���D����+ Z�28~y�Lv��k��|L~R���	P���"?�t1EY���ké�`�a���(A�u:$ԭUAA:��õ��^ΆY���
�gPD��]��M�����o�x����1��W<� �Q��(�r����qY����sY%�p�z��a&�������zPWq;g���o��t3b5�\t��/��$���O��`�6,�4S�ڳ�l5yO:q�)��\��ϖC�Phʁ-E�~1ɂ����<6�oW�^�����EJ��λ� &>J�x�6�]l4Q�.������p��i�<�P�MO�ZM*x���������ZR��&�C1�	6�)^<�LC��w�&l�/��C����Ж��3H����ga��{!�`��П��{#�W���r��w��X���C�!'v*wę�����-�7	^�X��þR�ߔ���$����"�ޡCc��/!<-��u����X�L��Q����)����P��!���$�B�5{(5��^�&U��Q���ĸ���̼�[�9,��5�\(�&�|eu����(�W���Kr;�R:Vhz�|�c}v����z��U������ݛE�F�%�Y�,+S�p�ѧ�o��\J	��W�@Lg��*�K"�5B�-�>��5i=P�khb�84s�;�bFV����(���t������#�Ɲߪ%	%� Y�D����@�M�C^<X{!v�\?����+)r�Z5m�Cn�p"��H�x�=ΘB�k���w��E�x�+0����Z���uK��4Sv.���Aq�CI��K�"ϩ)<���'���`�/B)�FS8�/��]�
�ړ���=��p�Ys�v�����?H~��N�&k��ObY�k�Ͼ0����?���ήa(�HY��494�O^�wa���h]��[	��"�23WJ������	ؕ��s�p���B���Vm�@ҢVȈŨ�)О�}���9���՝E-3�H��]A��ҋ����Q�Mw}ѧ��g�/<�2���3�kFY��3u������B��0��R?�J|3�R�˙x��J�A�d��ܤ��Q������I/�j��a.[o�u�0���=���y����/W ]t��X�Z�o��T����[��Ǐ7_L��O�c8S"i�x�Db�/-`�{�h����߼=|h�$�3dV�\����X���U�%;q� lRk2�����A�";��&Jql�K����kf�Y�����G;:sm������+?��ˌʍ�V5���^m��"��������S�uGY��ե�V/m�Y��󼤭��H��ⅅ�6�P�S��E��BV/�4�|�z�F�!�+� =����^h:I\Ք��	YV䄭�ۨ�_6	o_k��2ԹN�� �<z '��Cu!_b	M?D]̚����A��[ ˛�����^_x�N5��zA������TU��H);4���|����Uu4���H���Y%��Aq��S>¸�<.�J��ϓ��	6HN�y�֮�ui�l��55
\��Q���ŗ�wf��<ZbK��*!��j���+��{�D}����N����zC���'\ b����|��JE�W�T�����f���N�M��:9���SPl.D��Th\T�ޠ��P�j��d�\g�خ��'A,W$�ƐD��c�0����_��	=��,]M���W-A�����i�
��� e�g6�<'������G��`�FV�qBc῿�1�Z����ʊӉ�ǼNͩ��y����B�q�V�}:�4y�J�%0'Q��vT���>��0��K�YqKF9������wYFƴ�{��
�#��8g�!�R�����)}y��s6�C��X����ۏ�P{[���`h��N>�+��Vu�m���M��r�� ��JJ>�|��!~�)D����K��#�	�-^�����YK g����!Ye1�}X��-g�7_�����	�X�Lо�������@Qcߺ�D?J2���8�[1�3�s�m#���56����]��EA}��/@�����!���:e�4��q����N��D�:�d�����f.d�i����wi�3}����S��	�W�,��:2�LB�r_������e���؎�`��N<�u��^::��Xe��cb-��`�;h�$-b_2߀�˰��@#�Dh]o��*n��3�=g�M��8�@�����	\�+�NYD��yk���
'x��7�nS*|�}S�t;�����(:��5D��$��%G�Q�T��H���}k�F��B�����`n�`�J%�F��S����~ 8)��x�1+��c�������Ξr���J��S�I4�$Ǟ/l�8��C�T^�}6Ѩ]&�D���	rN1Ƿ�v'�HT�y� ���a:0��40�g�N�?K�x@�&��oz?�_�k�6^�r��C�]l8$]���E}�����:H;�+���w��s7ɟ���{�Nfr?_���.$q���CJ�{�#uEs�F.��9mI����+Sj��vP�X��;��`E�w'�\w���䔐�=ɹ�y�q��+`���UYx�WV5ʡ�oV�!�<����s10�2���k�?���]�l ���q��Z{��\֏e���@��:�3�)�=3�mH=4�S^���V�X�A,�q%B�9�Ŵ����?�[�څ�φ.��Ҝ�v�y�%�6��A��<G�eI�/j��J�u�4��&���7�o'�x)�,�c��:�Ԣg)�~����a8��U3�&�����M-z��~,��E˲$}��;p#�֕�'|�{�}��){��M퉔MSf~���D|W��ޓ�4��m =��<\��h��B5fj�_7( ���0ZA��զB �7�o�`ؚO�s<Sy��a�3�9�@��VU��Mm��tO�,]dr�\�gq��w�-���
�zlk@��;B�Z�
��P1�IC�38���:\�WUQ�E�?@\��cZG��Ǎ����6�����q�	��6�>�� �r��ي:��c��ßʍA�	��Y/�٭in	����(�&t�Pd�#�@(�2�0XWO��(��UЭ�l�3�qY<f��!�����6Ѩ�]3[��G>ıG���Q�i�o������R˩�=g������ 2�k�^���(m��F%A[Xs�8��߻�k��<��,n`L����vU� �k���pWY�wbẩ�P�0��f//�%r=&�4�o1�plA�(PYu"�]wz�<��G���[�LtV���=�5��@��]�&�$��8F��`K�C���������Vh��y�VW�����5o��h�	��>��4�t�'������&A�H��h��Ϳ�ՠLު���������m Ý"�Hk��s;�$Mf$l#`�Hϧ�m�.��h���	�2��i�5�7�X�y��0L�t28iT�\h�����aP�m"���V�@��/����L�b��kB;'���xh���"7`�[6�n��ѽ%�}ޝ��
u�Q=l��)��D����NaT�4�պ�P��-h^n�+j�il���L�x��CA���,G|iiP��Aj/5�����ߏ~94;*�}
�'/��}c��U�F��O���&�f���3Vօ��<'x��{\<���T4a������t*q\9�.�8u[���3�s����O�U���x��KP| ���xs�ʕ ��E:�X�WP">��N���x����L���p44�� � -�1 f�E,kX��ye��3k���ʇU��K3���]d �ۛ-��"�T,�L�WA(Xe��[�����ꦮ6(�+0�K�"
DJ�o w#1Ut4���50kū�s_b��y8G&�(������٭���9�Eq��Ӕ�	-=�7�?�!�&���u�Ѯ~��BuP�i��%�B�
X^��ſ��WO�%4��D���W�'N��z�E�c�z�]K�����u��,NȎ�V�t�K7���<:�i����*��K�gc�[;�h���`�㞱.hm��[���5�R�菾~����?ee�	/�ݬ��@��H�̲�<��U}U��*�b���«%���3`�����ur��j��>*쭯��`�FF��B�Ɉ9�+n.t�<پ'BAt��	��������  �m�f���o ����r⮣��]K�1���A��q#�#~(��*�G��a�k�đ;WC��.���te�d$��.O!���t�7`�}�2v�}�k��j��?���B����S+*�d'�_Bu(���ȅ�Ԕ�[�Y�O_%�
�Q�e{D;��c����c���n�yَP�Gg�#��ŉl�Ӿm%4��?��7&~𾹴iP���Ϫ�p�Ю�����4��~��ľ�-9Cg_X�5��O�J:qҼ�}�j��6�D)\;~��56�ș��X3��3�H o3G\�ť\!�ԤgHs��m̩�t.����/3t��5���7g���q�I���y�N^'��v���~=�C��+����ű{F�"� �����������Op�P�Zp��L��k��~=�:Hv�0���rzk�ֱSZyMnKdG2;���(�U�pձ�c�[_l�|��dZ���Ln��t0i�P��h[��3��r�OS�B$�5�}�����ȓ�ֽDY$^��m+���]i*v�&�pkPh��g�)�)���<�Rd�'�Q�wD�T�2�^-0]Eu�ǋ�ߝ��eÁ'�7�|�5���˒���$8�S�a������7�G�H���pB���tJ���=���_�6��#<�0�Duo!��6�eUb����>:��$H!	5�����+c��s	��rvd���+H��==۠�xK�o��T~��p],}(,lS{B��?_�ۜ�;���K̒{+�L��wnӼ�^~��](�L����l\u^Frͭ���K7@��D �~8��M��\� _����qa��ǴZ�A�iY�OHT�F���ެ˞��|^���rM��
TY�D�=r�]EX���*'�UZ7��!��$�x�y�q�.�?_"�xug�|��{��_5!�A���?��gX�@U���+�XoN`���_8�H�V	����W��� �E(w"=�����A�W��D]G�k0�$:�}��)��M7� K�O��?M�v���C�M�
��E��Uu��̰��OE7j�qot=�ʍ��Gn#�m��X��'������G*�{�t�� #MeJ�<_+IQ?r^��0��U����g�-��8�E0ҥ������d�U�J�B�咤N�L��uاЋi�b��7��wȜ����Z߸�!��4:�N�%y4	�����5I����W���[F�yʽ����:��������{@�����Nn���V5�^=�{V�Q�W�jF�U���^p�F��9,��Y1�f�����G������ �����$[˺�Ǫ�fj�H�c�Ǳ>1s�	`�R1X1L\��%Sd'�N��0�|]���νXZ�[Wx�\ �%�A��I�X?7(ɇ_ķr(/E!�!�V�r�$�q��1]��<|��$� �!�:ϕ�9G[��`��{M;	 ��e �Ϻy��.Є�#��4=����K����/�S��r��Y_FW��ui��/��`�T�Y^��%s�p$fط;bCm���L���p�i~t�,L�5�����$!p5��I�F�}D�#�����U�N.WK8�Գ��ʌ�l���#�*���4�_9�6�m��vW��b� `H�+x�=�P���?	��' �ʇQR@�;T!���T$��;-�@ܟ��Uo?��s�t5b^����M���T��1u�W7\B�OЁ�*m����j6	@�1Y�����l���(�:�1�i������ǋwcq���dE�C�X	LQ8XB> �9:�:�ȬV��oL�A��nٗ��?�II�0%�o\$�p�;@�xeR�)��#6���J�n���\�z���X��r�/�l����Ӛ����I���������`��*ȯ6����f�f#�:w����:;��:���L�o+3�U��_X�qÎ	k����J~�1�dm������-,�-I�	o]�tg�>�a�
y(�(<��v�M��A �0���͓72�Z���YOǔ��*�L�7��w��$[RM�칖xn�!��%��{��/�o��U8Pgjs�%�`�j�N>�(���F�{3v�b��-��֬ �i(-��,�����<b�1?����R~9vن@�u@����y��^��AݲIS3����{�J;bGLދ� �Z��߮�V*}��a���� �A"�Q��jJ]�䏺�5;+ep�Q�8����
+>x�O'U�4������ǭ��q��.��49c;侴"����3ͅ!�����d7�I�����C�՞<ٳ'~0�"�K���d�mAcή{����Έ�~�y��������.��P@(c�<j{D���~BV@���NW_LpU���D)��K�ͅx�%Ŋ_@�sD�DG-Q��v!Qs��b(c���1�\ *����d(6&3�q�H��}��ȟ*H��a4+~��i�������#�^����|^OS���ŝ.c��Gg���#E�m ��r@��Mu�3�>�b{;��,���T�D�*V��raK�����\��)_���k�#=(N'o�ӓ�0t�coOQ��E"�l1b7�~&���bJ<�[��G�
"iY��j�}=5��|��c�����m�f7�g����ݩ�=[�:θ#���`*b�?Jp)�eO��v��ܗj�@qA����@�lR�4����a:����K�o��*%w3����ќEX��r��LX���z7 L"{xf@j�i�K��~�xُ�������Ȏn�����,̰l�l"u��rR�Gm�&5��d��0	����Ra�`/�_���e�As�Y�w�0��H����S�`��LP�ƽ��Ħvh>D����|��7!6!�,H? ��?�>+�v�-7|1H ��i	{���5�;�
�w���K�y�j���)��X�öћ�Ju�h*J:R�U�Ʌ� �����ڔ]�B^��!m�O]V���V�aXΖvʴ� U$����$G�G.�n3{[]N�b�Ƈ�\w�%Q��.����]�f{�h�:��MUܧ��|0m.@�����nΫ��8��=�.��Ԋ��,5C�*'؃l|�AR�1?8 (�\XR���M�(��������0�8P��\��
9�������q�1)z-zD��lK�d x��+3���Z�|2n%@Q�@�ƫ��].IF����M�^xknQ�aw��I�v N
�\�����wW��B�+_f���h�� Х)�&�K�@�Ҁ`'C �T�"�r�=����g8�U�I�5|}*�MM_�Z�kuO>Le�Pk[���P��Ojg&�fE)��<>G��(�T'~������9���\�ZU���6��IP��oHM�v�@�̍)q&9Fu�CMO�O�ȝ���2�:t�r�ʏ�8r�Ę�������f��!L�r��!�a�٪�W����������H��@�C� "Z15�Wq������~X�Z�-��®F^�ۛ������^c��fBS��D�v��/��̫�~�8A�E�ѧp��Cv�@3�H8B:_
�\^?�-b���T<����� y�z޷-��e���$���W���tr�\m}<�\@\��Χu>��K���oR�s\��El�|�I��͈� !9���S�O��
$�j���'��낻��fO����?@M����F�xJj���i����#�+�]�������.��廈*W8��f�g��7'�A�ιi.}���_��y�2�OE��x�Ij�aI��c"'(�G��Pv�����E��{��7kV"<�l�2y;ҘX�B��H�^�LC.����u�����a!�߃N]n[ 1G��V��ԸȌ �����`&� �x��+ҙ)of7y��;$�<f���r���Z��}�FK{ON$8����)c���o.�4
5�d�[S)��~,0�	�ƥ'ԩ/�ǉLy��������ޯY	���_�]�Qٚ ��C���P�������ꇭJyp�R��۔�񛽒��s�,���Ɉ,�-�ȦYqKK�`Y��\��ϡǕ�YS���ѓn��\0���W[n�v8ĐS���3&c'�n)1�ͦU؟� 4m�4 ����s��k�;ǭǏ�N��yq2�,PH���>�Pڑ¼��yr.����1ޅA�Ʊ�A�j  	�L��Ф*%�V�ۭ�\H�;���w?�L6b���#�VN����VۿY[�e����Y7��IZ��z�@&�&�N�
�������$�.��*,\��Z�q>l��2�h9p�w_���پ-���B_����(��o��sC�Xw���U*��B��%��ɜo�Si�����,>#����;aX]� -[y�� �����a��և0��a6�͐����r�Id+I��>6��Y�q�CJ��n�(���pʀ�3!r��!��d����"(u7u�̉Y���wZ��0��"�V��|�F��(�q�x��v7=��r<���gzd$1@�����Q�*�M�n[���@�/�{qh���֖�2FoR~���#��t�Vx�\��xtv���' ���'@�I|��4���Ka�^Bl�w�v����υ�~�5H&�rz��e����ZF�t�_je1��5�Y2�Ԟ䉲;�>,�Z�h(�e Q�i��xE�����xo���j�D��`Ɉ�-c�qy�)�@��{��R�3.:�'|BI�V��(o�n�,&�P�:�z[�A���m�\�/�%Ġ��٘�~̥h1�����m�_7���dy-C-$���N��#ᰵ+���7	�����Cbp�%��z����L�{����$�:�!m�]v���FH')yG�L�hB��O��ɷ�|��D�[ż1���i�<�;�~|�'M��߳�����X����D���
f~��p�g�t�3�U��l�Н$E8q- �LJŽ����e��*P�7I¹iBd����_+�D�ǵ� "J��N�.��t��~ɣ��|i?Z���ο�R�	��2�9LN�� ���o)/h��z��[(�^Yn�\��������mh��o��#C�6��n:�Y����f�!��r���#?�1-�}�-�Ґ��7�xvvR��y��>�yՄ���P{��L:[o�G���*�b�U��eY�~�&/�i6��+���ح4��a8��V�llwKz�h6��8�#��P$f�·B��C��ԙ�'���ɀ0�%���E[ ��.Nc�lw^Jf�Yx ⡈K�'}��|y*�.�<;���,�N��%���CLA�n ���zL<g���		*8��~#ť5D�P�s�����
n��9�"t��w�[_��l��O�w�7�A��`�t�	��ޏ3�R�hĻ:Od0'٘j;�r�[h�2qYތ�,q�nR\ݛ��k��<>�����(5J��f:��zbI�-ll�P���{���P_���n������s�ƪW���0�X*�ɼ�A4<7ބ�Zq�1���_��V,P��&�t�Y�u� �}�x�u'f�8�
W��*qgS�Pk���d=���?���2�$�F�<Ad���2���ô|�0��o�W�����
=�Ӯ1�Ҫ.O���r�����i���]Y��L߯
��uZ�R�Oݼ����^Գ9�&�2N��� I�|��M�U����Di8�;	j���oxgy5aO��o%b�ӂ}FS�p���F��d�jZ��G���L������L�	���r}�F���[Q�I��`h!�w|���R�<5z,�m||sp�{>	n_Pȗ��1�D�#���ۖ;'wZ����\��B|��E�9��"��q�`���M��5rP҆7���1��ooC,7��؈G\��"Pi��"s��C���T����e�5@#�����~���hP�d[i7�\3˦"\�����T��tԬ�`I��
]K��|=��v0��Eo�����W �)�]�S���!s�yi+ܭԵ5v���T��o�����k�A=^^7BOXV87M��!j_ˍ�R�,#�dc�*j.����.p��t9���Nm��E��H��<V�������4�=�����|�X�۱�}��ə��m�����I�kv�D��e���;W��2�����]��
�u3}5���{�t۱c_p��h�/fYjʆ��y����y���rb��8�7�	$��FtZ����;�ԥɕͧXiut��ԇ�C��o�|���Rn�mxo9�q ��I ?��*�v���
��q ���+qi��d��ɾVM,b�G
�y�l��з>=J�Q}�;�"M[s`5\�Z#��M��y���;$+L+Z�Ǿ���7�㔬�.Շ�w�-W<�f�{�tN&�ˑ_5֥m-/���[2f�q��K�G�q�R�Nӵ�?��xȑ%��1��҄��{������Z/jYH�&�T�p ����+d�K軾{� �-��\{�����"lo�R��"^��!�F�����)�p���\8i��O %HXcx��R�����76�FNs��X��e`>Cr��쿃�m��{�@�c�1my�����}����@ޏ���	��|>#�`�_%k���lg�v@�ǜ���7��èM�!]���#���8~R��'{��}i.��Ѿ�uS_�q�Ƴ�k[	/C��P<��v����"i�|�
�X�sl}N������˾��|��˷�8q�]ƺb�6�;x�"��4�oE+�����ϞֻF�Z��rr�+�3P�U�b��<��
�Ƣ�~FҌ����[;^E?:�����C7p�!ӱA9�6}C��q͵�ud�M'S�o����gXY���s��Y�;b�|�,�ĵ��B�\���^��
;��Y4������1��:%J�� Kb�q�F���/W���'=~����;X�H-/�q�穪	�ؑ�0far��O?��������~���t�\�Y9�xu"s�V�Ѣ���x��0�5VG@y����
�@�п>̳9������RH�_���w�'���#�V��iC_�c7Ր�]��x崗�SF�=��kz�^Ţld��g��A��%(a��rkeNW�YY����8:菏��Y�!rg���(��^T�X-,��?��}U�8��YY��v����lј��$�<�=:�d�hߕ�v���_��TT�#�4H�o�P�&���Ӻ���s������AI���=+	3dIU�����&�Q�BO#�u0@�0����9��U+��m�⯹�+���
�W�^����|�M�2��/���5�C���^�Jd��>��yˏ�h�߷CL�M�a�~�R���$ZH���K��x��ׅXNR�'^�qc��������쓷�Fnlޤ@g����E��s��`�S�Ũ�������&إi���L��]}�T����j� (I""�~��o���ׯ�:��Ѡ}6���Yb;o�Y�X��TO��������g#���:��鎥T��$�5�m��H�
��=6s|�#ӚPb�h�X�_w6>���{�˷���Q-�f�ր�� lo��ܙ)�`<+D[�nϸý�F k��D�b�(q�����Ґ���MB!k���eA�`�yH �0i��8�A#�8;�����xe|����eK�%DbdP� �Q�xV��@~u�qr��J�p�lb��V1�;o ⟀�C��bE=�l�A��:M����D�I�f�9�����<?��+^9��,�A	���,��kC�.|��n�?�ǣ���e�@&�d�pˠN�5 wp1��B}��<8�?�\h�p�~�� ��v��� h��6��ﱌ��Ĩ0�+�����
F·��U�,gR����$���Ž�$^o��ه�!rvAa��`2��I��Z<C��7�j�p+�����'�2��yJ�I=�˷>��g�� ڟ��{�������}�`$)H���#$�Js�[�c��;vTm3���NϜ����<��Ptz|tjV٥bRcͅ���L?8�Xnjԟ5�o��Q[�)�ʟs@kF�"䍑�5x�u��&�� �wT�z<�E�3�O�8Ƙ�Ġ��e�gK[�&���"��������i�GFg-3Ւ�'�6VM��l_]e�j��m������"���=epR�)�N�S�4� J?��YUt r�|���V�J�9�0-�9��E��{C`�Bfk P���3(�3��3&ʚe,�%Q�!o��D�A7�x��k��g-�8���g�	��X�O�zq�v�F���(�sݑ����ɤ��}��C�k�M��u�d�J�)q��sݶ~[H�-O<.K)c++"{�j�Q�(_	�FŬM\0��zad���Mz	<`�YANbD�jֳ��P�I��S�*+4���t��*�E��|���z��ա¥mgq�?�S���%6xQ���YK��K��6T)�BL7����gB=�Z���%�	CY6�KO"ze�����K�)�aK���ǎ9�z�gށ��ޗ�sU�Q��KPp���)�� P(lM�]j�T�?��=+$>8|���(�6�^* �s�jGo��"�� ��ԉ|��e��6��3���f��Y�Lt�!Z�N��Le��o���$\��Z�����z�fW4s9�"!�m��|����&�(^|���<�Ok"%�V��ܲ���+�����`R��'ΆqR�o��P\��'�0�7j�#�N1�Y�,SW+��UE�U��as/���A�^WwC�mg�O�����5AB����J'q�����<dZ�m!G�^v���}���<�-
�W� �0���d�K4/M"�3��@R�F#����{*i���*��Ĉ)�j���.�T�	�r���SyQȥ� ����̀��d���6[1Nv�k�R�YBo{Y�]���y~EF��x|t<^�<����[с���νw�^ij��O%�!��	 �$ �U���0�*�Er}\A�A%�t��S���T���ec��Y�����&�΋��KBÃH��-E��0�i]���~��d'{�h�j>Ķ`"�����p�JT��vc��t��:?�(V�}j̱��\y�ʹ�u��N�������9�N,b����V��3���tG���j-'O\���/�`�<�}=u��8��!A�c���C�]��B��6<Ё��o�6g�Bʟ� �� 7�o��?+�1'p�1]l��l��_[xp�cf�R�x]t��iFJ�O<z&��%�I`��}�(U�	��V��Y%���+�M��έ�Kh�83��&��xT�������l�;�u�P�;�?���s���5=�t��U�>���y���O߀N���L�������T������A2������;�rс+˷�O�W�k�1����Hv}|q;#�B�����\]�J햻�Ҹ�f��@���@�`��^S�`Mv�䡨l�����hcC�#q���#��������l�Gm!Eq/p��������nȲ����-��i�,�f��?��O�ɢ�K�X�Cг����Me��:���Z^�3�Y��A����YF!?a�WZ�%mpP I���;.��g>y��[tke�?�>�Mm���c��F\i�e��Q�#��:|�g�8�*gSZLw��D{��<1����2e���,j���D����1K�|��I����@�{�~��K��?�b����,8[vA ��f������������d:|�f����)Foi����B�7���_-x�MN�^�_y�vk���Te��i�f��. �Y����W�9�����^���a;8�
H��/���2���7�veؔ�y��΂� �&9��iGM�_v��FJ�&�$>of�GP	� �� �^��[q,�m������@֏?����ˠD~�Y�U/�l0Щ��S���7���=�M!�I�i����/�g�&�7�;2^���.�#�r6�����n����L������]�D�����iO�/�6��rPz4�>����yQ(}[�9���l�~��������ʆ`';�׏J�$���z�ƞ"u)a��sԯEL,7m!IX��<Z�%	�fMl�3�z���s�SK�ѹ�F�X���~��ׄˈ=GN�1P��z@�]p������j�?{k2MG���[��S=��N���	JWe�C��~I4���BA6sA�P��G�To<���|s��b���<hF*�Y)�K���%�ĘJ4��������G*d��:p�rB?�e��v���}����:��3�lͪ�Qs��L�<b����:�A�3�Di3E�Z�����˹�����0`�|cN_�kB�pjA0�H�K��L�]6�z-���d��0�沓���scp�֯�;������O������+֦���u�I�/�/�O��F�Fm�J��E-��`��w�C�;֨2��1���M�}_��@���O����]á���fɯ%u���xi�/bB��.�������Nq�j6e���8|����<r]��$��%K�g����,��W�W��t^�d�����J�'��6���xp;1��s�&����x
1x'�K^����6��b��hO+E����,F?(m�#qk�L�1�;��'�䖕�%G�:�^��۳W��Ȃ��u��u�e����-`�W9jD�|��{% ��U+�OfU�6)��U%h 0��L��D�ʜ�)DJ�T��q�s0Rֳ?]���NߧT(e�`�sWi��4�[[�ͩ�>znM��Y�:TPɦy#��5��u�aY������:8���T�Μ�ocH�^uS�X�O��,��b�Λw�5���()p˱f��ʜl�c~+4}�(S�t.�y<�
�rv�)f��Qi��v���fU��.���)w�����u�Y���ttA�)�"��[H�7]�Q���	����Jk����|L��;����;sVd�`תZτP[W��F8�o�DŦZ���h�W9]8Qx2�V5�݂d���LU%���Y��l��V����An���L�Z�o���5 X?�SV4`vhaO��{)h�6X��8#��h۔��-�'�L���{D�rT3zW7c�a\K�)2�m`� �|�6���G�h�e�!)D������c9�t `V#��k��ƒn8��8������
@S�q��8�� J���%�ihα�>]-K�̅I�ֆ�(��$�.t?��j16V�&�_��џ��p�A�β`S�o�l֘����v���q�2��j��r*�<[#\����C��99�����գ�o\5?]���0��2,h�k��My�:�bU��-����-/�P1*z����RΕ�<�+M���Fri̋r\�=ҜT�,iT(����c־jGz=h81I���Eh$jc��m�۲�fb1f9;�G�����rY�Z4R;7"��ѱ�M��Jbr��7?�9Ӕs��mƄU�W��	t����	�־�F�`�:5�*�[�ȼ������K	�_�u��D ��:�]����������e�C�z��x�7�'dA�����
����]�0-��׮�T�*���&wn��.@OY����:׸~���:�q	\�Z����W��xQ�l��=�n%y�࿶g���WH%��]�&Hp�-%��t��`�0Ӛ�S�и����c��2nأo�1�_�F���=�*ۼ�w�S�4�m>��dz1$ь	\h���?#�����O:$\y:�N�����ǎr��S��i���#����QrB�Bef�Q	�4N�o��"�:��H[Z���k<��^���bw�����8��Pqz���p&5P�B�����Z6������k1<ځ�/m��:7��b����k��cQ1�f�CY��	��'z��Q��0�p�6@U��r"$� �\	b�E���u�.���Uv2oDآ���F�@�?���żUhq����ѐ|%��}���g$��:�BQk5c�Z�?BV������O��e�?Sӈ�"��l~�Uj	t�����>��7���-�H�Vgh6��]�N��דM��ۈ7lG�l�q:^6�vp��F9��O<�N���8��8ga��K�wb�T�>u$��3W���[�<�w�'�FR�wv�(���\�X|B����>�9afI��11��M�'�^q�	��w�,��T�����.^��rg�V����������v�؃Q�#<K:70Zn��U4�9j/���ʵ6h��~��H��2�&���b�&bR�a�x�
�(����=�5�'���H1�B`�L����dvM}��tb@^�3yA�?&�P�>�VZ����u��(�9�a5�0:�&��5=qZ����u�T�hr�NĽu]�I����WnA���iP��x�g����ڽwΤeƦm>�ބ��eD�g߁�`nR���s��ĉ�K��aNJ��ܪH�/[}�U���إ9q�U�
)�f�&�&��4Cڦ��|!�e�V���$������)��0p�&U����5)9�Ȃ���B�GaX9M�ɱҿ�)�ߕR�$����R���/�W���;Q�Yyw\��[�T���(eo�Q�PG��8)�̌%�6�*��h*�l�v�n��u��]|Mw�oë���$��*��TB��`������#�I/2'���6�R�MK��T�Hq�Q�O�����8`�9Șw�嵹wt7o!5�9�*��u���6�n�'�p/of�#�i$!軞3�kGq�C����[]�EA
�m�R�Sm�UA�BBu�@�oexwO�J�.e��$UL%V�'/t���<����^-N����b�H�&/�Z߮=q紤�&�i7ٱ�p�Yt}�����d1���q3��1q?�ö�)[��g�P��|�[�6k���q��1\A؎{|y�&��IC��8�"�y�&c���Ga�X8���U��Qo���A�Q�K�̜RC�PS�i/��^0��&O��?߈�h����PY �-�X����b��|Ǎ�(F�{f����M��q7��s1�RU�'������3+�Q������H��܈z��0o�@k�/ϚH��3�`��E��N��O���%=�^�-SO�`�
C�F*7��z��P�������?m�<_��� �|9r�S����w�$nV��$�������pxV�%�Fb.�H�n�L��*Ç�&H4�8��)[���*�զ���)��m"��e�0��,L^[����tk�{[r��q�P�-躴n߫a ����͢M�Q���ʝ*��)t��+u��At�6D w�ح�߄q��FpWI�c�2Z����F_	FTǣ��`A���\�_*�ܯ���t�~
�����b�M9T�g�р/V� ^�������V�/5?`t4�I��X�n�pp.Ez�Րd�\aBv%���x�:�a���y�!����ea\�P?:�+%6#�7!V[fJjl�{ú���9C�UL�M�.��&�ow�A���dY�~�k-����O�6ˋ�~:�3�L�I>����?s�}�!�k\0_�����|���z�!G6�ۃ�χ��.a�t�����`%�A���.��r�|N���k��C�  ��hI�h�b3� ����̔^?0a��q+�������,<�0���4�3�� ��!���~�_�����Rm��MY2ι]	z��9�:�w�h�����k࿧�T������"$�@h���l�}��B�>��	�f��lI�����o����ٕ�l�>E���q4BP(�PH�/��K�wξ´QX��5y
ݧ.2|:��7Q����0քG+��z��v5�'Ϣ�, vѴ�!R���7�3�0{֪�L�/lɉ���{0����]�t��t�8�,s�rA?��$ȩ�_��Ypg<�>����oF�џ�W�A}�!�i(]YѴ>�jE�Z��"��D�}W���|Qе�1���W�;�j蜝�=��Q�S�;P]��t���|�yR%�6�O�./5��K���cy�T�ߑq��O��k�� {JP����2*q�W�`�G?�$m+Y�.�{q�ޱx��s��\�|��g�V^}�����&�.��c��f��9����+������+��
\!ԕ[:j�#�Zd)��>��(�g�F�����8���6۝@�Fd �͐�
��BI C"-�(>��Y��y�	�| �>àD9�0�����P�(�	���ªϖ�Ų���:_˃2�|���/�-)�	��+�ڤ.~����$��j��M�Nx����T�\�S�h_0��Z
�ǥH@UK� �9d_�b����&����X-0$��./`:#E���Q�BE�iE�^�%����h����5��ڊ
/g���'���� �)��04�|#'
 C�9�[��O�"�`��:��s�JH���TT��f��r��!��´�^�㛳t���u�"��}�.T��!����;wu��D ����2V"m�!M���
W�E%P7פ��i��
O��.���9���3��a�� �Ԋ�ɏZ*DI,��b�/��
���#�����Mf��Q� ���Ջ��d#G"q+M ��쁤�Q����b��ʺ�P�=��޹�͢�{�;w#���uN�����b�c���q�ŢѪ��z���7��!28��@Z�����}���r���{ȩ���5��?��L��3�*�4����������� J�w������X6>W��U�bD��*��-���dpyS9qS����f"�rZ~S�0ӡ��Cm��ZG�&eS����v������$���3��HѰ��>�����S���]M�A�Sާ�Е8,��Ę��ѾB/T�+&���[�Zù�N��-z��D�$3�EiÎ�NfO]�/@�I��pXp���X�=h�),V��O��mJa8ۖE�HV��I��t�"���b��
^ ̃���[�~���Z�c��el�J;��M�&!���E�@���gbIڐB���Ւ�b��R�fg�2>�y��"z�5j�(-V󓎹�.�w7�b� J
�*a{�d!�$.�=lnG % p�N�D��"����=� ���N��z��lA��ʎ���{��1z�=�$�oW�}c˲4Ⱦ�� �{h��R2�����**l��m4R�g2|y����2���2���ޒa�� �?�)'�J�L����������\�ث P�����w���\���9L�Q5W��b�j�G\7��e�#q�P�����4($��D��:3hi�/9q�b[�!�e����qH~g�u4a�4]�Q*q� �y�L�Ͷ�	�+�a���H�U `]i�H�'�1-](�a`8��H��������~��]'�6�c��>Gˠ�y4$ |�a/jz|�[��n���	åI�̮�|J ���_��(n�n��xወn��t�z��DG����U�4��C��F���~�	�4�~0�]g1���  b�)ǀ�&/:��=�]�� MR[Jb���݉=�c��2�����~q�W
?�
&Њ�$�)	�I�s>v���c��Z^F�8\8��^��>VA��
���e��}�����S�qi�`�k�� �Y}`F��V�yDH1=��X���(̗ �Qoc�͚��S|�Q�[Y4r�C>x����'��T?-�!'��5^�a�
�P&��% �����3�|�g�B-2z��4��
��k���d,T��Ln�ԭ�q،R1\�2���۵&{����d���V�/t�.�%W��"#"�1b�U���4;k��&nd�����X�r0V��H�n����Og
B��C�f[{�/�3��Ԗ��
_q}
 ���t���܈Uջ��N����dӹ����*.�
QW<o	 TN	�Sԭ���1�2�pH�t�ײj�p�� X֔�f���=rhi=�gS%y��8���v>�h�ǯY��(�!m��C���k�H�R�la�����w����|�F[x������D���O����3�z��aמÁ~�q	��ãǘ��c�4�����#���/��"X�~��
ҞW�d!L��v�ػ�Z�~��M����k���<l�ͺ%�O���9�aHC�g�|?+1D��E�v�4ή�c�о�?��2�U��Ef;ԣp����� ,N�5ϊ���<�B
��k��zj�X�����B�z5�g�
_�����f\'���ت��my����6$�A�5Ǉ�-��7V�k_��ShͿ0���_���D�G�Y�`�����l���J"��ߧp��U��l�]�78�^��,�(�4�����*)�c����;*�#̾K�w�XB���QF�)�}�_\,�G7YY��n�n����lg����{D!�rY�\8�>�a��r�k|D���+��
v�<3�W��'Q4�eP
ok����PI��㘏$E���쫤��*�F3Լ��KؓpX�}`�_#(
�<:����T����,$3�}�
>)5?�O�xs�`PrLD��C(�3WS6��0���R�i%[u_��m�Q*�Z��i�+���fJB�9ܳE�p��?.��p�Qw��X	�ӻ�j���k��W�52JYC���`?�[�\2f*6�0�4S=:.fs$='�-%Ӻ�@aR�W�M˕��@��w:&�0��ǐ�j�`̖n9��^��dJ;��IxH����Mě��[Nɖ��/` �M-7��bfy��+z���L�GN����f���]O�\���ݭ�, 9�O��`��\48.E�d8�:MP���v�=�����=i�_��C;.T�X�Ԡ����ZB ��UV���)o)[��k��� ����+���@������)�#\�j��2tN_��TO�zLٶ$ՙ���J:u�&@c���d?#�=
I�7>���03�����d����ډV=Z'@KDp���)2��7�gxKu��j�UB/�2��O��d�I����~�f����nm�ÆI�␢�<ɻ܁d_]�����^W��u}��h��KJ{��ypE4$;3Fd;e���vR!�L@a�c��}	�
!��Յb��n}��q�fz)9d�����P���"��nX�ՔQۛ�~UՄ٘цq� Ǒ($3�)�����%�����ۙ���Y�X�{�Q��݋�Ǿ�o��!�c%�Y��5�Ss����ո��t�Ɂ�_�-�v�3� F��V?p)�n"�)>�}�|�L�����L�3k��(Ͷ�E eb�M�_Du��u�c�"�7̇ll���EJ|�n�L�r��郵3�O��5vs7��s0�v�ҡK���`��`F؉��d�f�MC�LFKڻ���j/�X�bs
��,J�j2i%�^�גoG���6��_�Bїe��l֡��U��`�tU<��똦�DjR��{�H%^f5r����v� �Bx�EY�/x�G��c,�r��&dȞ*HE���U�)#hHpy�Pc:x�x��9���6�T9*cH�e��8u�-@����D�*)Ѧǂ,�Y\��xy���	�_����lSPn*��C�Y�;>p0� h���7��)��`�����Iۜ�O��Gܙ�/�H�;l�pW���k�Bv'����?JFNo�k��\�|c6�E'��R]�K#&�6j�QC6O��_���-��u���;�A���D�2�!�5���x[��s:�N��~lI3If�GL�g��-Hr��ik��xr@l���o��������Z>˞�/��v��ϔC��4��ײz��Z��!�>(糶<��d�d��VǷI[�2�W�!�X���6���;�R@@�����BfZ�����j�65�M����-n*8ĵ���Yy�$;JR�Q��k> ��A�{�����aMfǎ�#lT��Pk_�{��uxN�h��&�@��_U�m�u���z�|�C?*��a٫Ux��&k�a��B-�cz�zq�>��S�!7���G������2�Y��|0����e'(�����}࿤K�o�*����|��ǈ[�בV��v�zJVS*$w+�c
C��~��%�^"�	j8Y���V�xuG��-��8aO���$kk>��Q��x��6��8���v��ܿ ��g��n� Q��5�me�$DNK�X��@������[�A�-��t��he��^��R�Zj�K������
�bv\�&�W��]\J'�<A)���-~I{�e�k�o�����|���n"�=��ͧ�_\/GRDu�n�Ȯ=gtR�Bg�&�<x���c��N�|$
l�zO�~9��N��8~����ӴR�(�H���E��ZhC��g�����5�A�}T�Hh�����}�~��k��H�����*��,�;����\��=�sC���j�d�o\�����w`�9��݇Zs�Y=�Ȋ�\!�`�,��t����%���]�L!!�~4~�44��W�J.ZO�}�����Sse ��a�ӥb ��{MI�A<TMG�t�×>�`�}��
� �AV�	�!�������λ���v����y#1O��r�q��������H��:C+P��M�6�v�r*B��*av��,�c_�.��v�i�<g��*�@,��-��#T.y?iqTP�v7���E��*�\�(�Z�
��,�>�)�� �|.�%ּ~�S�I�td�o��5%I��J�$~��"�8%���c���Q��rU�<n��.+N��W�*����/���`?���*b��%�F�Ӯ���m
�ҊV��,�?�U�b�,��h�;��LI*G�;	^a�H��N.�&�?����Yk������.?V�wM�?xK��\���{o1|��ȵ��{қ޻�g��C���y�b[���K�Z8'IT,7�6g��� �Z z�M���f� �+QᚘB A�7@Ԣ'�X[7L!�V&�c*��j9�U�#ϋ�#:��+v���S�?�a������/��m:�7���)	r��Cj��C*���R@����;\v�.i4~�1��4��6H��`�#����Jr�j%���$��$�_�Qsg��d�[As��n�#�̿����&¢t�{mԱ�[zTW��}�����<ڪ�B�� [倳��Q{I�W�[���BuE}�	ta��eE���p�+�:?@Tu���ŷ�S�����Kޭ5QV�x�Zz��BmIQǭ��h�@)&�&�o̕�+����I�d�vX�	�17���Q�;�5�K�P4��5E�����dB��xU_4A������B���C�ޤ\��lV�Ryeл\�-���SP��k�;�YIw,4��؏�o=^�'��]�����łwJrn�[��SuS���II(��.�S|�+͘��W���]i�xϤH^d��y����\�@sc��oaaLh�v�o�]H�Z3v�������x�4[M�3տ��f0�`�(�6nt�>P������SO�UY��ψQ�]��(��[[�ӓlzq�JE���7/ҢE�u������~;;#~+�^oW��DA��̩�PC�Ȓ�S�t�!���˝�z��]���Lgl~)1�Y�7Խ#�Xk�\oH�4�����__9���i���C��v�v�#m:qH�7�s*��(�$�	�Da��O�_���� >��X�j䘋!�����b�=�G�?�g끧��Z2|�+D�*�J�>�*g�Z��1Jv-ՙ�'�D��%��%/�f�a/IeG���y�:"�Ã�Gr��c�A4���qGu��G���柧���"�^�2iл�M���V�R�fW؞6ҩR���rm�vTPTq�b\Q��T�����q�mtT��?��\�X��#��@*�L�["G��3�o�p�y�!_�������"�/�s]��t}��N�Ŧؗϕ���p����C�[P���z���S��7��? yq����fBz"Z�>���+&`����&I��Р�������kK��4z��N�vy��P��?����Ogi�I�R��T�<��%@�9����6`���������^Ֆ�a^�G��L��"}d���߭��=���WO�������QӼ��̈́���p��m�`��OW��#tS䢙'��k�Xd�͏)dجP_\*��ĺ#s�ট��ݑC����76j!�i4q�lN�Nٙ�/��R��F����7r ���B*��j^G!�9�ݼ��8��<���+ӏ͸�h_*�}�"�>t���ھ==��n�_�\U�v`����2Ϧ,����e_��h,���}X<��7�QSm�:����i-���U�
��*R�������̘���,?+�~�L+WЊ��J���s0��s��x&^-Fk:~��ʞq�8
d�
��o��7�6J��I�Q}���(r��0���Q::t��R��צ ��<٨�����T�+$~��@����~|���U9�0�ė�D/-)� aS�M��0A�L��c ����R�}؅!@���R�R8Y�]H��L���h�P.�.�Efڦ��Lԧ��F��������QvF�G�7$л��dd����y���\�@��t
��Y��/*��S��i�O�cHF]�&qza�m���$v�颪YS_8H��q<m�li�u6��sc�$��<�O����X#p*w�����m�H=R��@x�����u(���T�P�>������ŭ��X��+GK�xeۜ'W!����)�/.�#�O\Bv}/�t4�)�:���$o���X�ݰ���OG	���@�Pe��5�[��[��%޼Ȯ�$�>��dw=�Uo�ѕ-F��o~D4mx��T�o�3��1��aL�T׵� �EN����B�`5�'`M{�E`^���UP�fNMl����{;V����E����� ���nW�q�5��뷷�W^�fq?�>��a�i����@ܵ'�]Y�k�3ކ�<�*���*�����Es�����p�ao�M�R,N~f��Yrwe���i��r��ھ�U��>��2�'�D-Ն�?r^����pUX۟���CR)��|G9��z��zLjĕ�vV��UES3����K��桄���AduT��P�$
�R2��=b,ŮU
рXč�ФH�� Q90`�Bg�6�*�^��>��2)
��|8'�)�i���B8{�q���bS[gA�兡k5����:Ko�7��B�'��	��]�v�8�݇��h�\4j��#�h�>B�����{,�YQ��Xx�6�m<�X����j��5����9\x�vn��`�]<@���$."I���7��}	KđI}S��u���e�!�H�]�P�ZJȃw.ـ�uZ�"I�����˰�!�(�_>�#���6;��V�d�!�b�H��D-5X����D.7��$��X�Q�
im
���D�W���scv�KL��4%��U[�J�ꥊΘ��g��jߛ+�n�̰��ؒ;���c�8�1B�ڷi�M��W�
��d
ɶϠyu�O���'u��}���M�ް�c��xB��u�l3A�"���)o	y$����dEޔ3���r�̔�G�""���I50B���m��{>俑�[���	��=�}Q��Eδx���a5VtEQ��!v�dہ[j��谊q#y�QK���]��YG��d��z�˃����Dw����T;^>}V�E*P��[W�P��^�͎̥�B�U��;�ò������Q�E>�����a���;�-�
����t���f����>�����!4Z��ߏP�Ƴ9������J����fKf���t�gD���3�c�����n><k-l]5�8ޭ��'D��[�]���u��e���/��oc~�S�ac�C�8j�O����cpjVK��{�r�x�"��n;t.zS� *yݽTwA �Ф���,��w(���E4��Q-������=�u�3��4(9h�������ʑif-W�Y6��|8�?B|���ua�u��UZNI����+k��5/C׹h^n�kFa��M$��c-�Z���(�p�n�~Z�29g�O����k�f; �#e�Αb�S4�SV��[Q��÷�
-�}9X�F��l����4S�X;���oj���ƬLv�fnrD���3 ����A����E��:���a�Ef�QI���k1��%#���p6�F:^x`Z���̓����bW��s(fa�|i���LH��+p�IP6�#��w>dL����8���^���Ș��<c�z��˨.��
~������{ZUX�3:�CQ�oy��A�r�Wy�}ƅ�n�P�I�*(�:L�Ѯ�Z��%�����W�9��oYW�)��F��L�>;\�Kg�1T굵�����L�'Eݑ+��^iQ}����sL���X�n��`lp�T06B��ن'�}M�s/���I�ְG��n��=�|�חm��d����h0�lҪ����4HB�s��<���?0мd+�����6�ۑ��g.=�s�P ���qw2�Q�I
gu�<B ���_�$|�"=��9!��.>!V�����A�Z���RLJ-��y������M��?qAj,��$�� m��}���7F:��O��Dݑ^��4d��F�;�}�y�(�+2���Jr���9�iPD#�-> !EH�,-������cc�
��T����Џ���@�Hr-���ȳm/�%�|l���P�hǔǼ�̪Nc6���
f1��;��UI?��2�B�!�N`ޣ�NV��U	lË��w�ډ�R2�I<��m���; `HٹW��$6U\�;���o�P���+�A`8�\P�@��%FC�Ps-�����=(��s*��:�
�M���A�j�d�����i̝���6�b
��� /�O������ީ��f�"W]���ċk�����ϗ��lp�*���E$���6�a�"��/VF�k�糝�<(0m3�2zuY���Ca\�w�:x|����|��ݒp���4GH�U���l�a:�US^�2�j��B����<�A:�K�z���	۪�lMJSY�Nɶ_X�^L-����H�f R@5ɍ�~���t�=�%H�F(K�Е�xpz���+�:9���b�S@��)
���4�{��P3�U=8�������B�˺��é&�M��J!�˫yjz�>��kEl_���'����-�X�-!nO>���N��W���i���7ՃW䦼�9C�N��,�#�Q� Oi	�?�y��^�z����A:�#@ys� ��]D�A�
�Z�-�U���tׅ����^����G����!��_�V��G��H�I���3��	��������(�,��X�#�">����/������J�i���
X%�����SZ���C���[^P��Eۥ�B� >�w_tQ�^�o/����-��8S^[`b`�M�e1�E�!��i!5������CէNrC��:�H�04�R@��Z$�J��!�m<�Ĩ��`*�f�`e�;*��4�v���v#���=��}]_9C���p��hT����#�����y(KO�G��OY�r쬄���߅q �6�]�����e����H�M������x�e������&Ӷ{�};]@Am/���������
�U�g9�v��&j��C{O��+EA�VHq !@5 �	�� ��Do���-tB��L⥤	����@�]��Q�:8N�a�t��,�[�яy���1˞���;_;���a�O�>G ��r�4���W���MX�B;r�U�����ɕRE!�ڥ^�[��cH�dľŒj߮}����E��
�����:P����!S�s�M|Z�͹�#8��f���h50n)�Kid�L��4�����L؉�i��ڭC����
ƷUH��y��KxkӅ?���"껊�js���w���������A�ݟ(��Ły���p���ߩ�]���O-�W�颒<�X�)�S7�{��y!~9%����x�`�7ST[���(L}��!^7\��Yd����+���?h��I�:F�jP|��@Nh������o&iz1b\m����]�,0I����"�~�91J��m��
!�<�֫��ӎ�����
{C��}����g���h��B��L�Z�~�ܥ
��^*�b�i9nIί4j�U�@T���GE�����x���'�:IB�� �@����O� Z�j��d�ܟ�s_���X�3=�(lsk����7K�Doq��x^���G������hɼJ;�KS����̯L���g6��4�jO�).�&Zk-4��:�K%��^�3�l}�����r���]�  �7k�@8�5՗��}/JU��P'U��ݍR i�v���iG3w�|_��H�^�Dg�~�Zg�/[�+�7o�[v]���3�/�Qtwϭ��	τċ�O�|Lω���T�`��w�S�kcn��Z��E��w#��x��@��&� ��Xj@�q3�H/ ��+�Gz���7B�X|OGL
�0`��p9nê�k� �j��ǭ�M����!�k�k�Ê�*s//�р泀6��|I.�R��-cPؓ�V�l���ӑT�?5�H���=|��|˼LWQ��w�PZ�j�do;h��=����%0U�Ȼ�Qfc�#u��T�l����KY5 ��>t[�@'���c(���>p�5��^�S_�i=��O�����3Ԩ���]���` lhժ���]Ef5�q�nW�º����M�c3%r�P���F��CP��X���;�$������?3���{�eԎ���dK}bR�,�S �fr�C8�@�)@%�,^L�QNl� �z���J��{�6�C�9��v�-�v�������m������g���b��R�R��(�-��������Cz����ص�toK8{�#�,|N���#W��pJ�v�U챕M���ft=+�#!���m�Ͼ����-7�E�bԀU����$�U0��YXL��$���y�^-Wǔ�eTɩ�����,(��%G������WS�r�?�������d�%1cϩOh�T5��8sW��+���@�S�u��$7�(����U��q���.[����S/A*K��RAz�� o4��	��4�55-g+���=�%��*�J\�MZf��_�q���W�a(ԫ"�W�!vg'V��cU��P���V�N$���u�֞�x5m��ro��Z��7t���]-8
QV�Dr��θh���V��#=�e�V����
ƞk�][On-���@G�n��;�#�d�׋�&��zNNC�%�l?����<bP����࿬Ӝm]�m�^[;Qºy����mS����;~oc�U6���#�X�G�b��\��I�h;|l��k1G���3�K���?�	�L��z�����Pr/hVe���Ř֔��E]��k�ெ.���i6�~��^S����N`���@`j��&	%��#�f�i��Xf'�c����Ș+�x?..X����X�DK��W�AH��E��E6���:�Y�$d�+�R�8F/�¦c!����I��d����RL���s��ܷRot>�n#P��!&]�2 ��X]�T�����5xC��H��a$��@���WQ�]�pҜ�0+�bT�y�!ˠ��%ç7���Ľ6��>���BCZYl����?�,�:Bq�Kۘ�����\f�O�݌��kV\���р���y�4B����.&��n�
G@D�%�t��%�t�w>q���+'Xb2���F���XErP?��z�~�V������sJ��z�0HTZ��`��y��g��;�LG��Σ]ϊ��'@�ix�5�3Z��L�4�2$�I�eotS��ej�6��kW����Z\���V��[�iJ�����,?��i�B@����S0 �J���Bÿ�H�[�ڗ52��}X��oC�#�Y2̛���@;Ő?�L\5~
�s~s���Q��Jt�����3�~�xZ�X���u�\O)ٺMg�+�g�"�Z�W(�k��y���-4#!v��z�[w[�i�^���iG�,KFk����e[�����>���e�|t@�}i�q$#�~h�#?�V�j�
���w�K����=�nAg$Zi\�	�wZdTTSo(�PZ:}���-���Ґ�?����C�8�A��X���;�k��ka���c���XNL���g����m'�������#����f�;���v�/LX�_�ݎ�#t�K�K�{mr~���j����?rA�}��^�Er�3>���TFK�T�e�9Y\��9����?}�&�
��ѻ�I�NP��-��5�"W�փ�@h�����1Q���:}0�M��KR[z!�k�y�VG_��MFwv�LԎ!����h2ݯ���=Lk��D�$�Ww�="�<�!��/ 2��)z�Ae?za����k�l� �4�351t�Ed��_���#bXz�������	g�R��Gl=��u����H'}���ѵ���e*����G.M�����v?Ym�6�����]qRεI�B�*� �ꩣ���R4�T�&8���E��;�=R
3���������Bu��̤���6�"]&�Ȏ�n���t>�p�^]u��g�r�y������@��M�ȉ��"<�\�%���?�*m�oW��(��|BD��̗Ul��)7m�������`��;q8��i�B5�q\+c�D2��r&lP�+��>3�A��vCD�%�[�@?�m??��)�GZ����V�ul_-��v�bU���⡛�+-8��F�o����c�˔����,64�HZq���EV��xI���;_�ۄ��H��Bv`�%*�mS����JG�:;0ٜ���A���R;���T�[cbi�U�dh�Y���C6�D'��[�02��6?��Q���B,_��W�B/7ڦ���R��4.�oE�oH�����q���"����C໋�Kحڐ����y8�p�M��~�L��]��x�0wd�BX`	j�A�j�=�0�>���?_+����B���v
Y�A@��Fĳ<�m�mo~3�A��u�N��lE�:[��{��'ΐy�_j$���{}��Ɍ-E���$ꟼ�ъ%�]�@ښIXȥ�L�
/��M^�'�F���W~�Ox�vՄ�N��#�fDA�	��,���l���(X��t�h|�9���N7ī�,rM���hFSp��w�O��Hd��/�<�v)�+��B;��P��<m��B�Mv�Q3u�ݬ|�(����t�ٯH�n��s�iכ.V�1Zk���v[T'wu��s*D��[����D{��L�����t�a#�F�c�DT�P&�@�gԩ.d�3:��I^۵��V�ҁoG����8y�k�����9�q�q>T�׳�"�?�P�c(8��d˟ ��k	>�i~��erg��3��D��f~ۃѼF���!�q��4c�y�B'���J��Q*�}�Y?,4Z)�R}tN{j4r�[�,�g@��ې��e�<��\�-4������\�U���쫁����v]}	6�h%�z_ob�� �d�{M��A�]pXJ�p��	Z�W$-����tA��BS��!��l�;[�h���U�\_��&ߪ��~Oڸ�ph���Nα�t��)<A����=���o��Ꮘ3m��>��5m�r*�>&�t�/����!�(�7����X�� �(��,���߇�VK�j�Z��Լ%t_[��E�-K�:��4������0� ��.�y��RW�8�K�9~�6�;`̕l��ʥ7mnG��n�^�HIuFL�k��q�$�,�ֶM�Ȝ����`���o���c͆�S ��ƸnI�)��Ux�t���S�b�IR �?B�=tU�1��.�2W�%�4?m���u�2u���~ُ��j;`R.J�xruu�~?��Q��HS���@G�`���".j ��V;�S�ۚ������$�� @hЭ���`����\^�g��z�Y���ۊ����aD*�QB����@d���o�g�3��)���K��M��1����\b+Vˎ��h��h5�dI���2_>�i��w�&@x��2�SH�M���sL��1�|�g�ΊH��nʒDa>J��dG����k�N��Wh�s.B�0|���y��S!�E��!���i�u�N�`U�t8������C�h��<mwJ��3��("Y�s%Wo��+�ƶ��A_�a&^ ����%�	f4�*��=�2g�/E���u)e��%+���� g��D�<�6��B�x&���C�+t��Ⱥ�]JB9-�[��"A"H�1��#�w,��!��@����Sr<\O�6�)�
�ׄˑ���S'��aiy%��8�w\T)�Sy=ȼ���������]& XBי��+d���խB���w��GY�:WDc�=H�TS]�A�N����if�E�+�j��7.�����L�ΑM���X����$.�>�;dA9FN=���z-�/�V��Bxv�����\hX�Q�\��9�pK�&���,6�K��J)��#E�dW��Kyo}�9��0������t(��J�3���6�*`���l��ac'-���"���i%�����z�-��<��#�bns}Z���tsP�ϴ��5<dh�g��c?�`��Vvs�n2ˍ��9��
8���8~��Qq�;���3	$oY4,�G���5:zP���7��(~Nl2ݕ"���r�[WD�?V�`��H%q�<������Ș?�*�5Ċ%r�f�sF�(i��v����:�ؓ�KA�Ef�1?��4��46���t���M��J�P�cYb��'�G��hS��`4�z��
�-$��+L��#x��F���y�5�� ���uhȑ�ϸ�P��Mv8y�f����h�_~a^&'�'�X	�`¢�>0z��y�Zj�F���o� ���_�7�4�N���/Ȓ����VPh���I��q�S*5�1K%/u�}�՗Z���凸��n}����^��}�C��2P�۬c��3%i�C��9w`���O:V�Ðꚃ��.jg��/ǒ���LG�����#�b�������k�}wˆ��6�biܥ��f�1���(���R�Zo��\̑�aˈ�7Nld]���Z��T���Q�N��v�_��9ؘ1��渖;>!�]+��be�ɸNu��K���>n��t�6;�m�V�s>�1�I/k����?�1�c�����Hh�n@e�����] 'Ѭ�52�Y��G�g�^Gtu��\peؼ��Q��&D�(�5�Ń�h�nQ��{@f��RӍL$�CEwk��3����z6�{���=O0�>��������v����?A��ښ��0�g�n��s�Gq�u ��B���"+?��C�Zw�#f)�.�i�w�7¾޵�\�h+U�ڽG�]g�����lu�ҕ�«��{��7�<fizƇ5����MH���g��9�t~Y6�$�I��n#��Q���dl��{�ue������x7��ḫa��S��	Q�iN�ۍ�|�t(�M$ K>m~� "�#/�y"��3�y��N��}�!,�ʉ��<"ʙmh�2���G'�0�d>�G��z�rN�{�n�d��<<�Ml5;���^]����|��L4���f��ŀ���:�:R�>���N��4ݔu����Y�R^��>噸З���0jl_k)x  �K�>v��,iD����eB��~��P�H��%c��nJ�2�����啡&��GUj�������]�K�P�K��:KMt�[�!�\���1�sMp o�u��Pb)F�*�Y3��봫è!���\��5�%0���lA�T>ĝ��&�{��!���J6OIj������/��n;�p7p5��U��O�P�C��f;��]J�m�ڹ r"j�n漏D��t�i���h�/��֏�K�w��`�s�6r���`��m�a�P���¦��
��쪠0.�uo�]԰c�O���$��_;p�Xs�<��5�2BG���w�����u���)�>��m��$5�o��JT�p���pqM�B"�<Kmt�鋶�Gp��O�-�/gu�����s!p<�L��r��ي��W*!���m]�q�E�/63^ޗ(����a��i�8��)C�i�@�����TkK���|ZOR���X����>X��ǣ������������x�A���*����;���m�>�U�͗�ވ����@��ݳ�mOUC�:�&�W�[�� f M��k1?x�]�?/"Y#Е�P�6�98i��Gj�>L�����
�% ��F�z����U�ݪ3��ǆ�PD�������Q
�J��$��LЉ���`b�����}���W��O%"�{W^�4p�y�l���7�U-��M��!����������=(15��Z��������,�F;5��ޯ�!'��Z[mAi��Ϛî(2NK�'���n�ޢ	�I2�	�E��!�;�>n1ƬxP\���o�DT�'Y��# rr1����M/�3̨d �B�c+��a���,����("2�H��@ܒQV���I�-�#X�<�W�ZY����򟚹�>�2x"Ā�dԺ|��i�1+�tD6u:�2��;��Px��nE\�m�*#$����h��ȓ<b�)���lw�8��w�����������ӃU��q��Ѫ �V�P 	ٛr&�V}�k��:�N��k�aJb��<��M\6�a�iI����ε.��?��<.P*dz��y�U�R3��dx��x����.�{���9��m恼`|�y^�M[x3���-q�C�|�r�W�P�ŽV�>�M5�\�V�?��'�C+�v&b�ڔĨ�zV��"�l��ơ/2'�wh44л3�y�ν�O˰L76��TT���S��j,r���Z��=�h�7��8�}`q�!
���k���枎��Y����	dפx�BhCXK�J=f�6�`{JJr�Ib
7�vE�os�z��v�G�M��xh^��v����S�Bsʫ�8���	ӯ�%�F5�;�o�
�!|�1�m�S�6�xbv�Gٟ�}��7[�8�%�.�	��w�e�}�i�$k���}O��0Ʊ,o����ac�4��ת�r��P�b�u4��s�w	{���9��H?�(V��l#�3�[eZa�q0j������9�.m���<R;{�pe񇔩T4�_�ܦ.�XO�H���/���&Y �A��f`98�L--����*�`��ꂲ"�@���a�b�o�nq�Z-ǝ=.`�u'���.6�qnΝ�\î�)ɮ��m���Q�- �T=��q>LQ�3�!����p���KrV�$�����3�@����6��)W�/�+��H�^�;䂀�H�;>�BJ�1н$�hq��ݞ�[����nNǴ1N[շ%o�N�{�du(�~�	�5�f��T�#��^cB��md[�4�Ea$*��?��e������d��cSM�,�b�KN���!���?l��?"����#��"�nE��T�c�S$�XkV����G�x!�ۙx��Uz�ǲ�J��ӌB����������ޞ:@VȭE}���/V�:�����D��Կ��d�^dC�� h{Z� �2u�)k��D��	A*����Ý�G�c`�c��.Bݓ'b�*�)/�1P'J��7�4����e�1NOw���	���MI>k��]�/S�[[!�y��Eʪ/Ĭ���H۠�I�3��̏S���G���y���{��g��v+��X@;����g4p�Nl� ��5�x�9�Le;�8`�I� T�#!H8�`�֝�JXeִ�!Π~37�Y?�NV��Qo��_>OEF�{C/ňj�����>^���n�pE������>ɋ0K��u������z)uEf�0�U q	�
nC�1h<��Q��Bφ�q���� �H���	�(���ҕG��L]7@��J�ȶA\�[�m��V������g�	į�T<R;TZ�u��ڵ���^�Ni0�ߨQ�~K�����ԇq�M��Rf���A
�x[�z��ܖ��v��]��Y>��SEJ�<^�ЉU��Iy �Nj���O���x�=��.�����U�r�:������?fĆ
9��E���?l�ܣ�fu2�u��v���׹v�P�r����,�z�
�J	�y�M?�qV��1�C�|t�Xa�d��O��`�re7�,�ܑ��yw�4W�V�]^��ڠ�矺�#ݸ��$�e��T=y�<ڶ�Y��*��*��Q�e�r�=��؍v�ƣ覕^���$Wz���cJ-P<���\�!��<�H8	�*'���<��U��E���}��~e
W4`�$}�j��Wd˪��x/Fε������A5N���cLS���/.�b~XwB�Մ�!ƒϗ�W.��%��3S{|Z�4ZU̺E3/�$h,�)4�8��w��dV�,�Za|���汝�`��LW���j�&-�bq������_��q�U�a���ԃU��<,�U�׎��]�?�jt��P����y�z�gv�(Xu�|����bvS�YW>\�s�7p���k�{�$�.�On�����YT���zՏ-�L�La�pE��vF7C��61l��@�0�1X����+WT�1CP��B��UD�]��^�[�yR���c������d_6`O�1ґ�m�B�	�����l�w����*�DN��!��y�ٮ4��L�EA�yF���VL�xZ����C�q"���3SN���@��"�"���
��~���kl�D�C@Po ��9�.x��jЫܺ*���>S�"KX5Zc���o�)��Dx�C�ӎ �F�Z����Ȓ���J$���Fqiy��)���!Vq�n�/4�T���uote`��:�K�0%�肽��,/����s6�����P�vЩ��v�����d�u1��M�֒�� y���i%�I��rE� �&�:�׺���c(x^m+1�]s�q��@(9P�x�g/p�tW�F;��)��$�hD��y���'�/��ja^'��m�-Ak��q1��n �v�{-�6zxU���`�����3���6!��ٕ�D��mnCb��0V�
���-��-����=���K(�w�-*I������a���3��ͣ�h�ai� ���n��ei�D��#�� �V�$��#o�ζ��n�'�<ce���T�X��.>��~��t��J�0��F@�����i�p1_�^<�A��K�e!��ɠҎH����X$3�lx,g�U~�`����$Ip�kҩ{�oޝ��V����P3r��9��,G��!��!��6�߽)X��q�,��S6�g�dچ�0��\D��F`�m+�W �&�,�y�� ��/�Y`���*"��P��m�_�X����	!��#�+w��WF��r<�V��%+B}%��a�vS���#��1C���|L�yo��ٹ��nʙ���mU��Ua]6L�l�����o��	ғ��BПeC�(�{��S���4鄨�5�y�
�
�k4��9�0$؞	��<���LI�`�(�+��zi2�e��kI��P�P���FoR��(u��^��>5��R<�ݰ(ḻ�(t���}�O�����ɏ�lv8M�Q�}a���b�S�![y��p�Q,�`��Cu����z2�P۔%����&��g�H��f�XG�gEZ�Ͽ��-:�
D�Mb������Ff8j�>�y�W��cg�_cت�#�܃��Ee��%pEn:�Lt#�,'P7x��Fj0a�:��9��WQ�e�
��ͬ�Bπ��co\����o�?�8aōt왡����O��Zo��^2�ovrX�^(�����
��2�5���������sF��(P����`��W����aw9G�����h�C��|!���~�/(,q����<�9H��.���L��$)]�~����8�{+A��]���ЧY��Y�w'�sa�� ��$�Dw��\b:����{�����sw��hf/i�q��g8�Qh�����ČE�C�aӮ�R)󒼍�O�\�ƽj�|�K��J�@�$wZ�V�8��l5�;���#:����C�w�3�0���:��y��׃Qj�;���� i'�ssfc̰��j�R���:�D�x������*�
!��T쩑�])�QtY�g�M^v�"�T2���Q�a3�L�BDywx��v�<����p��m�(���|�����G�J�G1�N�[�(W;����\4c,��o�I�2���QB��Wf���p�,���%������RUs뵿;rV��W���=���O�|A%��`�~^�!�Kq��w���5�VT�&���^c_�p��",c����[�t��Y���?>>�OB �Z=�����鯂q�&�����1zm�?
:M�	��<�C��}�5��A.���B���b=�s2�� �"�8 [DM<�\.�W���ǛCMr~a�+�@!5Y�����/�k;N� 4��⺒�� �<ԇ��+?P�.�� M��]*ŗ,�M�G��*�@/&��Ev@��h"H��ὓY>���i����?� b��<�ܢi;ۄ�K�R�����#R;���H��罎�"nD�&P�$�y�+rE$��w$�*��b�n:���f�@�kAY�.k�hJ�ED�FQ�y@��I�I(�jW����Q�
��o�4���`� 32�u�B���-��\B32A��ĢH'�H�D4y���f�mY�/2�4Yo�E�`�[��=����b]��M��U��pZנl�	�_:���!@n��U�Og?N��=��)|X�::�X�CO�:.53D�g��7.�5E���0�	��n�]P��YU~�pQ��X�{�k֦[���X5�N_��Q󰯢��	��6�Xi�jx���)��F}62~�q��TjL,`#��nhɊ�!>2�4gm0:��@U�&�L#��>΁b��M�s�+�PJ?�uX����?r�I�R����S��&�'�8ώF�G�ۘ�����I,c*-5;���P������ <|uEBn� G�����a�1�-Z�2 ��N�K`��D��AY��9d[��o���<Q��-�q.`(=-v�`��#r���	�47Sσ6	r�Q��i�.�-�d��sW��}'���N�~S6�%`D���E��]����b$�}{�,��O���Dm�m���F)5O��x��NyIDAʒ�M6�!L��eK�F��oWo �,&����s���y]Pf}ܵ�.p-�E���ݐ9m�9r�|!����w��`���j��,���j��/Y�g�J��3e"%�ӽ�ˏ�dR��V��5��ӧ�	�@�/ϭ-(�E:�u�7eH�݄ؖ�si�4q��K�X�O�����y���, kT@W���Xc"���س��J��>8��綷�TN.c����҂�9Y���v�A��{����F��[�@�0޻*�7>�"?bUB&��b��M�����{���p#�E�i$.�H�/0�MySR�q��� 2�aѢ?B"bb��>/����s�6%�FJ�P���I\l���E�[m��Gkh:I �����K�:�d	^��O\QΖ�:�1�-K(%�X�	��bv�X&�Md C<hK�<����MZ�:��X��f+��,�c�3f��]g?�vNN_��}5�6��VA�*�4��!�Y�A[naj���nu@��q��|�G�@�^c�ڃ����p;�Ҿ�P
�^!�\?����Z�Fݰ2�Ep-�>$,�g�`��%���~@ /dڵgd.֫��	o�Ģ�����[����S�n����!�A0}����4_�0�9�Zp�TKM�O�x���� Bwii�*ԝЩ�+z�W���!NJ��Ų���0�xh`� ��b�e���Y�>C�OnM�|\�$�_R�"&70��6�{p�+�Vt��"�z�����:<'���)�"^�g�	֡��O"�z�v8�ë�&��!��&�2��:��E�O֢�ƣL�u���8�m�<�%��5��?oh_�ikE=u
U��3���-���)LrA����~����q퀅2`�	�2�d�F� sh�H�r��nf�&@+�T���dh�KUeK{����=:\��ɗ���Ǻ�e�&�ī��ߐ��V��P,Kp�s�I"�-�|�h]�4����A-I[�x�u�.c(�{Lċ�d��L����A�O2�� �̰7��ߕ�$�*��1�����4���Bz��
�N_�B�*O����-i��
j��J��jI���5��Cbr�����%����g���­��X"֖+\9vVԾvk��g��RO�=����%���\�䀪f-x� Q� d�W��6ƻ��F�D�vb�b����'����%��5�q�������j�	/*�p`o��iw�����S�x;Ejd,Z"��7�f�jhPX&"������ƞ���C�|�<7q?�q�ē�@���S}�%LB��w���(}%֙�DG��{��d�f�
�8�tt�w�4�:�Ɋ�=e���b��1�Y���z�c�\�)L����F]�D�����q�x���Gau�Di���ߍFw�Wn����x`�t��R]�#zw����;n$ص�D&�כ��m��&Mf7U�b�`��C¦���"RԵ�H���w�Z�a�K�4P�P/k	Q,� ܆T���sQ��Ɖ�7Q��:x�"E՘�M��Q��;!fX��䪮K0f)�K�s�*��!ߔUA����O�h�D��4U�^�nz�i#~p>C��oI���6Fm$���,7/fF���n{e��NY�"���߀����gXg�v��4p��S ��i�}�>`�Z�4Zu��Y��U��ւs�[���2U���e�sq��e����)5�i�����f�5��N2Kz�Oq�Ao��-�ؙ�2�
i>��� *Y`x��'h�
�eN��n��}�2����wb��"���gK���R��ѿ9�R�q�����ͯ1.����傥�SHh��Bt�ܼ\����De����&�h(�Jn��!�e���p�b������,��6�����s���X;z��& ��ue`0/V3i-���$Z�[w��|L��]��!�K,a��f��na�y�������d>�i����4�|X3������+��%l�(x��G�I�ݷ<jd{��l�:�]J��]\ˀV�S�oUiV$	OŴ�M�D�%]ǧ�/H��v�4	+����*�`���8Y�|ot��y�=z{�����hb۫������T�X�����އ���֘O��X�%�8 ݷQ$m�Пh��-��u9i�B����X�#&6��PFw�F$���޽�>�$-r� {d{On��&ū�OA�> �a-�)@u$�����|���I/�16֔�����W����:�!����V�m�f�X������g�p��Cd�0rث���F�Γ���΋�6�S���g�h1�g�I��7�G����l��$��[��Zw)ž+�����.�c8N �=���Ֆ�M��}k*>�J��;��` �1i̷�W�J3�	�3��:�}�I�ֆ��������4f!�R�=1*(T��k�L)��&^N�q�HmRa����i��yI�ݭom20�16,�4�1^�f0����*��d\e���5��ǎ B},�>\m��8E���[b'T���nлoȘ6��ȉ�CݳEq��~H�+\���1]�I �J�@sP8%$[L?;�[zP�h;݌2(�|��O��Z:bbH_?{3"�Vj��N��2MEy�(�d��|h >h2y@輄�PBl��l(�Kr�rЌO���ޤ��+#}��DQ��<�9��"��eR
j����i��N������I�5f��V������ބ@�.�
d���l��D/Lļ�#�>��-�{4�`�4ȋH�|8^9���_ʥ���,M1��*k��?�(l��,kiz2-[5�IZT�A�&ON#{O�F����ǣ�/}�2J0������n9NG_#<�S�un�#��PV:���_�k�2kbRA�����q}4�5�H�a+a�k-a�~��~�͉j�l53j�#K���@�bNM��}�W\�mH���_Z��yb\JT1{߮m���*�z�9��nsC��Y��:����rg��7���(��B}!��[A�lKh>�����ş�z�%*!�7���#aК�t�� >6n3�c�́˓���,�&�P���7�hv*�j������k��.C����
����4~�0]�� )d錾e7�,0[]���n�%���&�tMiͳM�~�'���IV���d���7��O=W[
�tjBa���l\�Ohf�t2�W�u��TcO��BT�f������6�kWĝk���~�R,��ng*��V�-}�Lݖ_xUu��$�f���$g�8Sjk_4��|�����b3�-��QfǉB�'^N�ܹ0,���>	2(,���G��Sc8�g$�b�쎜��J��Y�.䷚E.(�����v�<k0?�������[���h��{��M­cH��JX?\lNI��BV�/��ŭ���7��ۤ��3��3Rk�v���f������x�#�Z��Ώ1�ȑ���2ӛJ��	02]#��Y �ݳ�*��
$�|9�����A����G���3��].ڻ�t����P����E�WZs���dzbܚ����)�y@~ �F�Lm�&���j�l"Yq�e���8��qޮ#]���_�џ���郡ٿ���O��/P�_�Q.ѩ��k�҉v����>y�F�ϴo��Zi�����b]g�BFA��jL=��%E�Z���V�����
D`3����Ֆ����3_�k�H���@=�p̭�����Էt� �mHc�S�)�|4�9���{M�3��,:޹��k-��ˉ�3��9���YkK���%�'���%�Ţ�Ie���{�bQy���3�}ԇmg�p(K�1��4��x P��Y�9���!����Q�o���H�`�r�X�m�m2,�DN�Ґ�4 w�e'^