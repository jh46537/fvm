��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0�����
����'a���en�,�=y��~{��i�#�sS�Z�àx�WW�Bg������𓇴r�b�ex�Wv�c���V[�4+9o]��\�S�������_���]U��J��]2c���L��<e�@�&���jX�3r|~�SrOa�{NR^����y�R�ΏD�|����m�'�m@�q��S��Ƣ,(�jݎ�4��>X���w�j2�)M��&�wU�=�a�;�k����K���b���ʎ�\������E�\��,D�`�������A\]��J�o�A�����^�.�c�mC5�h�9����N�
�.�C�!�V ˘�٬.#�]�	ޔ.�⏩� j4pTMt��U�uW#�����3��ɐAw����/5���C�اDt�����e���#�h�e�W��QyG	��,ct��{6k-���w�Y&=pK]kS�g7�̝WJ� �
�Y�X�K���L �n��ӡoQU�Iy���r���o2k�aYDx���v~WX������+��xe|F\u�R��0?ked�1G���U��'i��Q8{���=X��c�H����Մ�t>�����T(�!��ݔ�K̨��c��p��U�HF+σ�����u��֫������k�r)���{�J[���.�y?Z����톗���Va�e12M��M�f�� ��^��,�OCU7��P��z��˾'��0X�V��G��A����Ϡ������;HD�}<TY��HU
=�g�#�IF���*2}w�£m/Y��<5aKdATK.(�)�lԞJ��o�?"��{���nd�͐@��$��ltn��۲u����hK�ut��i�q�k���ꫳ��ɷ�Q��$�(�۽7b��	����fZ�������+��,|�$���j��ߐ�x9�����^��^�h!QkNR&�:�?�IVG�L0+`4�p\�F�?R���������e!��LV�~a�Ӑ��ߧ��|<¹P����i��d�L K�-{�	yM��j���#�r��͛_�s�0[ȧ
���B�\��9�.+��Ҡt"l08.���:8Gy���܅�(�%������Hs�1u��0UF��(1�rɁʞ�a�p�u����s�����}+RX(g}9,"�����LU5e��+���~'|%��T�>L����2��j�wRi�ί��x��uͦO���u��_i���W�T5��!��5@�&��`;�k�Px��?p]C=Ul
S��n	]<JÛ�^��=C�ş��j&~�]�ܼ�s�Տ.�ph�;vG���?���I.�y,�T�î�����m)�4�y�S��{+�H�U=I2䢶�ׅVc��\��[��X*fz�"�B�#_�毄��~��%Tc��b��,`��4�U��ܷ�����Bz��2W�&�������\1#���G����)�bh"R�-�B���T?�ɏz's�V`@/���b"��U������&��>1��L�Z<8C�d:�Ĉ���E�<����qmB���~t56Qy!Dm)��ݢ��\���$�$�����6Z�p�4$J�4\�/T��xUlPd����zIq <k�o�O¤"��2�;荘�<~��$X�o�Iw� U�6꧸.;{�{Xb_:l`s+�ek77K�uȌa��."��{U5�R�2�
<B�Vh�o��Ы;�PHh!1L�jQ@P���A��M%��H*l�V�֎zy�i� ���!,���/�x!����d�~�J"J��7�f!
E�)O��ľaw�Jk.�e%�ډ������^����bcY/$-s��Z��[J����0:mg.R�#�:���=�	��}hF�y��$���#E e��(�
����k���%�ł�4� c�*O���aދ>f�:V;��k�Ɔ���������c�-x0�l�	?ܑ�
�	_��!��6�>B>�3�{��Y'K�>��Z1�P����W���>��o�U��l���{*md�J�ɹJ��??�<ckW�IN*�x��u=������U`�t��ިJ���������V������u1_��}d'��a���,�@�c���f&��J1�PC�c$��L��ƖĴ%��8��&�5`@�������䫋��Nව�:���/t�=�[F����Z�q��o�A]�q��[v�B�=[gFn��Єm��������f�$6�Q7!�n�n����>����ތޚ�ݹb�&9J9Ϸ|��ރ� F6m���}����q@0űOZr"��ڥҡ �=I_�;�N�%��b�����f�j�����S��=O�4��I���7c̙&!�����|�OYʀq>^��Y��V����Wm)2��'�]}rln���~Z��ggI�,C�p/^�����L��`K����	�����ҭ��#�r5���	c�(���lux-y�%I�m�e�v��\������@�s0��{�u���i���>���W^���K:-�J<���T�J�4Qf��)>�u7�=�d���J��l����������N@I�����j�l
L����M�� K�hy��R��e�ų�DHC�4B�g�?�<�QM�x����G�u#�=O߬כ�ty�@������nz���H9C$	�oEulзΘ=$C5t-���-�*J�V�G��5��#�q��/�dٛ���?�$2	�Rr�n�o*l)�
�Xx�rj���
@ĵ>�\�&�P�F��j]%<�0�ȿ�_�>#���Q��c�6x�]�N�rt����I@8��77i��b��ߕY�!�j���	���0J��N��w;N�\`�G2=C����}Q��ba�[���<�� ��Qyyg���y�I���xŢ������v�G��|���Y!�9�6�����a�<K_��m��S�}����1�m&:��P���?X��g���Ϙ79�z����Ћ}>+f@T�6BǷ��Z�Z#�q�f�H�R�Ф����l8�hH�m�����K$i��^�@܂>������@�Znܝd>�q�;��M?�V��RuSA���5	��J�Of�.XP��iz֮�)ƞ	�GAis�������Q��ʠQ^ל(��F=��@�[M(�;C�1���>;�� ��S��:!aM|��a�@|4����ժ06�LO}}�d}?#� ���X+Ģ{�V6�͜O���un���R�,<\��	�K���1�ew��$���� ��$ʍM�H��*x��ܲ 3�K8
)A1�6MgW��)����i�{�okV��1f��b��0�鰖�!���Qwi�Df�5��u ꍰ8ݛ���p����M/k�r!��Ȝ1�N��O��̎b��.�杷9}�D�8���Iq�-��׻���!/-�]3]
X�9	>vm�>kKk��������Y�K<�z �g�=r�ڈ�A�5�}`%A�c�`}�?���-���˕��������X�-�)��љhKЭ`u��Z�Ѳu�/�Q"�9�W�%������KZԚ�"�=����cΩ5���L3 GT�M�~m�ER��.�)p���c�]��F�����T~e�#4 =c=��z�$�q�C�"*oi��k�$��B�C�ՁM��+7F뱴�F�=���e������SR�ia��c�5�Nc�X1iEYn���傀Wn��?M�X�!2	�U�z��˜�W٦?�0,�g�5������wVK]��~�od"O7t�#�6�i}��#�_�����T^#�ڌ�N1�id�鐪SY��m0��V�Ъ7>�]qEE9d~{�itg�)�{H�2��P �Ǆ��>܄϶6ě�kP�v�we��	�?�&��|�d�x����� �n�]g^�@��?NpH�d���{�؆�hU�~�4R�Qj��>IY�=Oω�?증#w4�Hx#��JZZ������������J�$ǌ�▓}N�T�U˿4��A@3	��D��N^~��'f~���>g�s.%�Qt\��G�ys�;p2-�ר���P�҅v,F�]����S���¿��=b��1	(�n(��!~����5���c!��L̦����7��)��U-*�l�ᕋ�x_��#��O�o^�j�X5x�syܷ�+�yB;6�5N�\����H���lW����5�)6����.����e��l릦5�;_�1W	;���?S����=<���]�m�vQ�L��j/�Y3�v�A8�h�v���w�:�����?�ֹ�5�8������7�]&l�!~���ƛ�]�)����0��A<s&���M@�%:6��_��O? {���Oj�*��DFtD���;���,�4ʾ��&lU�_�*�_'�b�-5�S�;ê!���2ۍ�ў�z��2��	��U�: %�_�;��?�R��n%