// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:43:38 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mMDc2TfpK0fXv2MmNBapi0RLZl3rwpRdibLSCSs7DEigF8H/ucxdo5JBLL0auCxS
yuC0DSv6pndp5TmmPdqYIWloxRorsVMsw4FL1o5SvF9itOEJADtwOX527Pnmth2C
xHH5nHOUUzW24NixvS2HoQHT/UQK2ohgyjsZhS6dQMY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5424)
DiQLXAIZdeKqcec4YlFLzoAHrZIfWFxsyHbwY+k1WZZBHJZnHWQ2OVxd+MP4P2Lg
SMG5lRK0p2F4dxr6r3v6QoUboin+gjQG6ZWA6sCICFY/IrhXBR64cho0aYkYSMwJ
VPHZJscVd2UdGOhX1zdAF+mvPNGDEAalC/uiIDeGLpYXs3t8Xd92IzpPcFiOXKbS
XaLzHgUjQQlVLzloJg73JTNO4JJ3Fh3o5Tq4ce8vZQF1BITdeuEG849+r/6RuAU2
oxb5hBWlCkLP8a5KHsSGTQF9y+vhQlvxvCoCXg6ORoqcQJuXuyVfvMi1OAn9zEJ/
v6Fi2Qk+/DE0SW+jmWiKJIjk2Hyo/QU3Lt/XWTdgqMbKlUR2+y4Axn/HSLK9Zi0u
RKXyjJ50WM+ANI0G1igF8kdPFYALx1S0BuJMYbM1l4f4o3M/lTcqwnTmuFsxDYgQ
c83za5J9yeH7fXVI5c8cgL8uRcGrOmfbAptn/+fZySsS/W2zDYqm82QIKkIf5oyn
b0Svn7JA3KCoMaD3Qn58srdJZN9C8+4lwgVEvtYUXUUxTTTbUU8Q8lUUgPh3J5Ll
PGjgsy05S8mWHxAZ10PLOSZuMzLUQCfUfu6VXJ9iNARM/4H/1YxnQ3OzBG6gsKVn
ywZlf4mx9S4T8jkbpy0GIqM8zZ+YTjneitn354zz6SeJ2U5Vw3qrzyTZBW2fvhft
wqK7TLe92q0UNELS7JGZRARwyl6SMhjCADUZhipF7tZcmtZcrNpbJgItLEzHtwx+
wXFuGAXbxbJsnV3n+93CY/CB6ATNIs5NUMDCrrxEonz+FVvvSGi0puHnWroOtJHB
Lq8EADMdPFZgAKGMJISWl+B9DqSs0qezhhz8SSQsTij4SqauPOYgx4kfFwoybLSn
1W//zb7BPRvFjBAr26w8IIxvEQQRKkg9p/0dS5zMhFRo8zPxjTuoKoKq5rrEAZX4
AMgMaqs6Jv1QkpwJS9mxH/Z4AU1WU+dSucTs5mmbN5mNCQX9q+uW6KWngKPnckOJ
0YuP9+iWGjQLqWl9EyIUKJ3GsXnHZ0b29xXojZiSmHh233TvcHI/y69YoLQC2dsF
n1egy2rEgmyTssEz8TylpDZOTV7YYM/PaeEMJ09bA/o0FNJacPIoY53hNp1sAVX7
vdcF/X98R/f9a2d1AIZGuyKjrs53k4BN0zXk1h8Rq96+FNKbEU6yAY/l+PoMTEhA
z+4li3Z0fBGNd4FOGIznyGhMEE7l04/JxDsv6gSI5muUvEVrkwKcfZP1+nE/VmFj
sT3u9xynWHZvJjtEYLeKNOWj0Hcr1HKv8eQVcqY/13EBQXgGAuzbZ+q8ikUnUJfI
5oE7ZgiBglaxf6x1HLq8tXbGjjvD1BNh5bKdgMwJliObEZdAhb10piAvhG4FPAfU
RkilP+LYt2PcDGsLtOnbtYu2+/TO45Wu3SvtW5Ff7TO3e078pf1VNIuzpxhU3J0N
TtGOKWz5sDInM/Ippv2cyFXc2yuSJoL+xIF1Fv0X6IQDF+kFgw6FVoyKPt+RQJpF
DXhwqAA+ZM+YUjnFwtS6gCW7jUlkzuqSdej4Z5XCHVP43N7OS9EoPbmLqa2pDRlv
v2c7dMwKVRwyz4Fpja9q5rIvNqkncrM1icb8P0NEtR5vCdCu9qETzX+wklXu3Xo9
6JRQZS1+5D/wY3ojiGMdztlUZxhmar+rnJVv3+4q1anKPlPeR1AykEug/XPj2a/Y
DQEsIpOGzyLrGLyXCFe914GyZGdHD5pt/5VkVj4qpctbiAu1PGkn/ER1GMVuUcNY
BHkfrsOZOoH91CZhxH6OdbhlmiIRPEHw8Z6AWbA1yE4y29kMbrzNXz1YcS2FMram
2upEwYrI7Nm1ovWJNCWrfj/w+VaK7o3JdYEqR9qkMguxT037Pj7DSzR9VsO/7uhk
j7jRppK3W0iI1y5TxZ646L1ZYaaL6qxrsg6usvtC9usibunbz2u49mGaRuwfiyAK
/PaSXPqKrOYrPwl/sZq9I349LFCMv6+NRGZCfsIzGOUvAWkDQjivpxotd6QxuxL+
SAMJ9ab6rYEE7KSTMynpihDxs9N2xk9xjuVoHePtU6neSx9KBy5YzFafWIEAta+G
9UppBkz+IXtVaXFRAVizdDjS+emx/I9ZhmjiM/ttS8Wb0Jf67ADyDKfzNFyLfajl
ls/i3En/oaXt8uKwQJ38o9/kwGMYNRg3glSyS4cmrdFJXDltzG5T+FNsNEFt152n
YCYwFwjsBHKbasQIOg5FH4inuO24pHCIjdu4rX+R29ZpoGSZDDMXOUlAZYsrEC6H
QRQiRDmUodM4lWyl5tB7/c2Lf0Eh4s+ocCrAtiFRcKWd0UJ/Mqd9y3acrWivqZNE
VXF5PbRnK0td/O9qRl9yLMgqqze/tHqHjeOfsGlylnL974ikLrBjdarSEa6k9JhK
Z0yzcI6AOjFKNA1esA4WNvB8Nkxm3UaW+Dkn4VZPaq4b+keM7dKzIX7jPOQo0AUE
dN2WSHnXlukE0oMNZK/H9DhhlntlhboZzZyqjNfG1WtGoweTaf4Q5oT2mIq1ibmW
VC11MQonMa5mWIoZjEsaMli7M7Ou6sxP5VZVwoCC1/Sl9/kq6HAPfZCHSEKbbmcp
hPzV94JWDLjSorWpF0d1hM7pUsEslS2Wlf7yATbsHXt17VLpz7uD1avotCd7B1zn
BWdAyqgbytfxYfPocbjnlBWJFQM4gk5+mS4PxX1R8ZMAvt14/Vz70S6OmwTevsMV
T7fznhkRroALZFJ0uTCHSkaf8i6GhehsPaoAHuv04FQ09kuP3elNJj7mjKa6vsos
OwU0YjtaL13VWTSaK87IXvpoYuyMKb0w0i3wCnnltXxb71/0sixN0FHAIhoxoj0u
D1salZ5jKAiBclC3jj0Tmzb86e4+7oDFhI1VF810MTN+Ljf29IruFkQsPkD7lKCC
lT+JqzsYUT+FyfbTIn/LGB4GatoGj3I+prXTvHRbAOf87J90QhCsNoHJYQSdkjp0
4Lqy+uUPyt/1uUx9ZRriwLCQeWMPR8HgE8w7gbu1nV4+CUchko2KhKg7y0dErb9t
UKyD9qawc75XNWnnihSmbSIqF+my1u/kZz2gDdnraW4HdfQNqwGFL6NUCc1bIV51
WLzojELv1kDqQrjUWgIgZR8Om75e5cFFiPoGkiPXIk63YFJ72BJ/9h8w4uhDwEEF
TaTZJHSYo7ASjxAA4bviy0SGSdejv5AuirFxzbd0hG0wj7p8RYn+N8dDabwB+4+5
el1NN7zT6UmU4dpGOscvUhL7xrPHzeFCD9yRJ9rlytrXil1ZeDbYW10m1TfS9Eo/
b03Cmeq6D5EV2dAxcde4QI+i2QVh8m1tojwt5mGld5LSWWpmeYafXvmUJXn2mzAq
lDkqWhLNg8aHCROo8i57+DmJAXFN8D7SjH9Bw2t7ACy5MVSncZY8N6BwvCZQtOMK
RGZwaiYEmUrknyzX1R7EmTSdn1GX4wkkkx9OzLeh49J56oNrOw5d/p2P+5eIXmfz
D2x5SB0U/DXNC4w4JQ4Exjv7KmkSkob+Kaz5EBc1DB7ru14H/L1Gj00Oqomf3VrM
WvikDP7aNHvObtswBjTocBmPEPwjaIs6tlb40QikR8W7SkzSKzyYs9WEpnV4xtaW
uIcSgUnyeDaCkxW603/2XuKs90IVl1AZjhKCNwmnxq7DVnu44PJYjpZEOrzXg46e
ncVuiEI6G+gHf62fp5+//rMBJrETr+wUuOUpjj2uFAYC6/pbI1FO54bh2L0JnpsW
mgjQZ8yd/1aL/oB2GUNIiugS4g2D/193E9lDFR8e7Y53D8VcJmpHpTaosbFe/Zq1
0uHzdnYuCEucSe7ArJP8plp47Wnws2RFX1j2sf/sn0dCz0ImlGhE+tutHmiOYCu5
N4I5AuERTzXKc/cJTBs5Q1Q2WICcZDJ7UfS+LJ9cmTQGKXPZ5iErODRiDuqbmWUF
5Nr1VEfgbsXPUOoYbul3xFBM9d97o+/Hl8wUf/wPLpRr2HxhWMMH8losG6+XHPTZ
w0VNqPKSr5RDpjikKXn2jmjMV6MSQE1QpFvogg/sSWo5yosuFEA9tj9S5Bt3xcov
s9iCWWAyYwjWOIiqoNfDrb6fdi4vfCAYIPz3atjjlhKTHhXAfSYZHup7SqhRWRxX
mZq8tr5haPsQHZOyBR2vyfLnTmBLhXNdQqD14d9FSuMqy6MDYbnbqVsTsP/YJNLE
kg7t2299KLuYQi7zq9FUb5lgTco9WVehr4CyH9o6dXZ6N8aWzD8zUGkY9Aotb/AZ
bDBmVyLtSZPY4e6Kx+T97kYpwc3E3PlJZ3tbyDYW53ud1hRPdI2jxd8kSV5ZI4dH
zOsLzrDm1o80lUUgc92vN10wyvrkuFpaXHptvAC+gHwxzqUeRM/G+k9DgqkGekGy
lpc9WPSl/Hf2yNlqk2tPnmoBNF/kYiEL/Nq0jiVw99fI+BVyrsRheh9yltFKA2Zu
yAjNuCipuy7Ba/NjDkxtQwHIPavTAJxsAmnEGrHmrVZ6nJgFn58cmJA9IGPZ23VT
ul4uQaDTtlTM3ZnGtCiwBtyT+ZYhzMCZW2ewZgk2IJ/CO4Fkj0A5zwX3fHJHSHJS
4trSA0OVXMvnLd9wjX1pF+gHVy7XF0HhX8nh4YjWBvoyTD8zfzEdrdzpo9zOXwI/
jTdZTFUTUA8yTjRoh0d85Xlz/qZJX5EYS6vo+6bvOb7VqmHXdvOBFzfELMmKmAMp
HKOQMZuASxgD8x9Z/bhxe6h+FXbBZxbfddggxzVYIVDkFp29fa/10DDLG91Wy8DP
34t7dl63FMgwsQxCf/P1gSBbWDbdo/eQ2gTAqMHtE/wjprlb1YvKukVQckI6pmzo
M0wwlQSsDK7mKxiX2ofj0S3K1GEfVBUiNg6/Pf/geSP6hnWrYvnDL3zHqzt+jCnd
jGPPSnOpCJp6x+EGR5i0UZYCp+W3KCYnMswVE6ijF0HKvCb/HDCthyGio0IEJlBA
v1hfLjv3TLPcmwRz9H5G5qhit/oauCtR8HpCjnn4JyuUr1FZQK7bGwTZmFnmBRvs
kzbrWt6L/uVSUfMZOLMctZMma1RBs68vzib4JOy7AAoqPS38O7GiGjOC4uBXE6uB
DQBpKW+q9lcK52HD3USOHrm91CNpt32f2agMpWblucB85m9uUH3Z9BFOPHFcwHd7
Cfwxy62I3h++SL9eRLt3KI57nGp3cjVgBPT8CsZfN8GmxnGBqDpUpl4p79CwWDOI
5YSH2eNZe7KWX0RIF0BrMA8XBN92wf8my4KlPMnHjSsh0j3br8yeP7ozT4PVTjkP
8ALxzdj2r1tzStzJhWLBfG2FKN+LbYIdLo6Wm8MxS/H7Qw3UHwfBNNTvLDIMgNIo
WDtv7O29QdOwOGOHh97LKJl2yA6+vHmmgm3WxLfUS5TJXOYoDs1Oc/ErFejA8UR8
ZoJKHECdZjdcZ2mB7x2ZL2oKhQOLM2IJcORA6Njpx8tOWJeTj9b//z4oIW4B90W1
NmBjnzF47rRZb7C6PXwg8SE5AhqTaI+8RRY44/Z7AJtZBuLZlZZyuP1qOqCS4c92
KufeCXxMq5Fa+9kYopoo3cECgFcQHNWiZg8I5viIO5Srx662L5jHNeAdMd6jhiq9
AxswBdprINdy1H82cB96anAyungsr4fFG/flaYzjfbImleM1VVRsYkgfZbUPryuC
81lH2TprkVKvBH1ClpSz7kFvDjdU3oiZHVgv0DvsrGt+yX9bEuvQ+l/SYAUUa59u
6AvQCmvpMjkrN28MLPxMlGZAW4OL7uNn3k5i46WJ2l5WHCnKvWamsrUOqCnWVhqn
Irzv/y9WSo/vBJPYQKPFto19v6kxtg3KCY4onTDfoJ4H12jE76LAHG/OGD7w85BM
wP8pkmNx8xqTWYsw591lgXXT1u22xMYJnY1km1rNLqvgvaRCWeDeHhdMhzCgODRH
/22rA2wAiaiOyjlO4gW+/KjXj9LtyVxCks4+dGrw36N+9T2e83EOaDBWr771+lvb
msuUd9AzMwseaQPTyF/ZPQwQd5BalnRQpb7tRPBgIkgGUHKwnjipO6PKtOs0kK/p
iP/l0Fqcj5NH1GSm5WlkuYwR3loS3kuX59L0QD0Na114lbXRcPLSKQws3eCAVHJm
G33SDiab41qlzEnbij3SWAEY8xtnLX9KjhZPpiL+s6albgasU+5zYLggD2mD/S2C
RABuH5xxIbNqSGWde8B1rX5nV3FqLEIcWk9wKi9honQFG9KobIhxhFjYrn/fJsuE
dy2yet5GRR9XXovJCgPvMNVoMn/7FBQUYqx8uNN/m5syuFaNSxMIu7hXIlrfxpYJ
l7lYCX3xJMz4TPz2P3ZZ08BTQZOnYKIBrLbPpSktsdK2WYxr/Ox1zrsJdf6yiXZE
2Y37YXM1rhA1RUByLhZzbCLQ0HRUbIKNWKPRhOJmruaawizAYdt64PSjfFR3TBIb
lgxKPJa0l8YB+W3nwW2sDpad/FoeiwqRBZ15oyuIHoAawihogKpdgI4ZJLFgsdTN
1PpgObQzs5/ZNR6M8/EULuvBP8vCGArd7wup7c0kgB2und9c/7WQF9PWQWt4tPYk
xnrhzkEDU9x7uhZl5jcoo/CzqAmG0JVcor1ngRZWOhBqcWVQedv0BUVpJyz5N8Cu
viUgGZ+6I4QUV5TLAY0VXlZWQfVX3FI9hybmlYEWO1MA9bNtOS3TMsoc+PVyp+Nx
4htJ5TuKCYufTgAAq/w/yTHDNNRwUloS+V1YacWCE8FxIA+7jpOhAMnXQFQRbjUl
Dbaidt6JPn+qjN1Y709c3nDV3r66U5d0gC0jfW3I4wWw+vD02W8xm4Ql9Y4KSMvb
XTxl1bp8qIH43W6ecQOARtD7gCevzes3g8353uN0g23LAHA+IZyCPSX4/eY3ly+t
Fcg0v4G2Wj62VH6ZF/KI43oQlXgZ248MLEer3T7Ueih/8jx8VJeL/qpNiQTNWN3K
4GtONMW7l/uZGos5LrJN4macrgi/yO8w/GSgWx62Jdtm4UU4vnPKPGsNc3P+FYwU
AnqC4KYAf3eJ/oMoHsCvhBK6Y0NvgSz1+vOV/uHz2Y9/NsNVm76qsKPqUQtA/Sfm
tq5PQWTWJww0aDQ1dFfui7caPo17TM16fo5QPA7cDscmnuPbuxKsCU6mZkJqLMGw
YerPYxSUvyUcUaMNPOUAfqF061oUIWlVG6IltJZETSdVTvMjk4iyP1rsN6YEFcuB
`pragma protect end_protected
