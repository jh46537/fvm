��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,�������_^�6�3�@�RU:(�3�у���aL��`3��0�B�u�9O���Ě��~�W~�\{=�ӏ�Վ�o�G.͘�O�daX��?gJ�����0�rl��P�P�s���.Bd'�e�_�<��r'?{Aj3_�N@xi�н�� ~z���!(aX݁)��o�B���#K�"Hx�_�g؊o�@�j�aL�%^��&�e�x�i��CeF8�t�f�DO����>�OR��颏�)N�l;���@�2M�[��l.xh�,{���6��9oOϦLNkdQ�m��Y��*#�t4�}�P�;��#�~��F\��QL���-{D�`�R]�?�gu������~h��B|�g���_��Ft�%�J^OF�KM|7�%┮����%<b��J�J�&KG�l%ɹ^�_�+�(���jz���$��	(��+���C�;�А�4Ş�[�	���.qn7�r�2���L:��Z���;��-|�։ǇDJ*ku��N����Vv���@!j��y�24��#v�����:��z��%�m��[�m%u���Ծ��\%P�T��[��c���71�b��b���ca���I/,?������#�#��������'Ge	4㚍|y���ӓ�u@��`R�o
�|�-�Gj���W�� ��u�G,�B(�h��/<�c$�O�ۗA*�C��2�$p���44D`�<QU(p^鞍䗣���?Ě��H��<��E��{�� 9����U]�4<=�|p��Jq.4wX��zK͇���2��"��4���	�i}�����S 7꿨N�����;�wC@Q�����M5x��k�9R%��2O��n�)����:�M$܊(�Q�/�g��j��o�6j�S�b|%+�Z�#�<�:�{�v��$��R0�1AEJ}�
_���V�|mOy�ǭk�0�dr��.r���r���ewl!�#1t+C̺YkzS]�#���l\�6����	ڔrJ7�Ҭ�6d���S^�) A��혫�Dx�Ek 2�iSH��O�kE�]c#�ݣ�wb�}�b��*�d���n��̉��^I�7�����A�'C���("vi�9�t�Fʵr`vh� �ƍ�%GͦǛ=�6e��t��$�5H5>z� �A�K�q �FII"�tƶKGV، �\4���ԭ���f��u,�L��M�K��W�v��Q�h�eZp��?��9r��\A95�����e8o/����_�	���0@��ԁ�&<ne'`��ʚ�X/����j(.#�\�d>缺�j�A�'ZN�TA{ 
�7U�j�-m��E>Rq?��G�A�r\,9B֝6"������Hl��Mj�-�u��h\(���2�Ь�<���򁩠��I���v�"A;��C��Ff�~��tfa_�7xx��9\�c������k-&� )�6V1��z^���/��w�-8��q�!4��3"���6^�j��d�(д�=�;��=緅��:Ss58I�k5�%��訮�V�J��(��e	ji��ԭH~��f"U|�b"«���Ao�Zh��9c}����2Lxꟺ�˻��^��&$�o���G����m��֤Q`��LX�f���o�H?S�~���7\�])8��a�� �-q���������iH"d��'���|�P��ȇe�V}@_���fP�������ۈ:�[w�%%���u,���:���K�xmU�c:�N� 0(���?	���J�|>���J`�����i�a��GU,��w���ʷJEZ<�%.m��Ʒ�x��@ z�]9�$�T�6��Oj�u�<t�
˷)�������8���K.��!���V�&y�@�~J8w�M��wΓ�Co:���I�1Q0i�"{������X��O4�
�u�nc���ǲ��8���;9��ҝ�q�'q��B��I���%�M�Eu$P�䩭/B�)D4k�mL�a�D�s-�E��m�K���n��fz�>m��W㴕6kB������XӇ��ӀЇ(�����N���GΚ�?P��@�P�)7�ϩ�1�� �ʪ��U%s���Э��7ō����9�lT?:�<q�������ɠ��3Zzs�9�r������ên
.8�4�OBZM]#f���W�Pp}��U���z�QJݤ�&�U����
��k/��ܖ2�-���H�b-F�&	�m�D>���l><�& �Jq��&K�	��vAR�c~�d�CF��k�`h��Γ|��>�l��[3	��+_�ŉLњ̥��>�*��dA�(ξ.ZY�L�Er?�g||��~���J��)�A���)c��Cזh܏"@���s��9w��:���$$%���;ac�2�W��CA���u��'�f�P�c���g�!�j��6��8�78����(h/v���yJ\�V��ѩZ� �^+\�,��
U�?V4��	Lڣ��U�"�R
���
�3�������&��?J���0Ԃ��O��S���~���!��I�˵����͞�%WG����r`/ǁ�$�[o�`�?���G����6阹��y>��@d��pe�E�$&T�'0�� w(?D��I].QT2�SoU0=�@q�X�6�`?�Uu�
�0�o	��Y�{ys�JD&���Za?��3*��V�O��c
��X�2�5ZQlD80CE?���5��2�R�w�	�8��5=bj��W9������sݾyǆ �G���U(Q/�Qa
Zl;Ħ��h��3�1�1fo��^Ϗ�S*�-�DMͪ;p9``ĦE�qð �pU��d����}����:�ac�_li>*��f�&@�#�ZƂ�x�ñ�[�.��Y��7坹�XG��[��HE[Q��=}�����W�g8�E�Y_���V��>�E�UKU(�����J�_k�:g�{��i'��Rx���44CmxKRد�ys��[�U�o�ׂ�PlM`d�b��nAFk���љ�Ĉ�H'��S��wa��K��^U��cj�������C���`b6d(��Q���އ�Weri6�$���*�%m���{�V��nw��wW~��h�.��װ�+ �6� g�MK����UR�(%�ٞt���S],���U��P�N�����P���ŏ��"cT�\�j �6 ��h�Rxw��L����`f:���	0+
���g�R3��H ��Gw�s��/������,����n�B�S�oL�M������t�ec���J���j�]�� �s[�UC�����-dԽ#���`0��Z7]��vb�h�6:=��!Ө�'��!cf�(Ӣ�c��SB�� N���D7K�\�fu�폱g�B���<o���YCE��q��MX�Hzc�>G�¨s�6I�㑂��C��Z�`����؟����k�C8��^	������E�\r-�������(�#�GGS� k,��齽=Ħ��x��S���@�4l�>�릮V1�G���ֹ�;F�0���Yn�Me ���w�����@��v�l�G��>[�'*5� g��)�n��i6�:�M��s���г�Y�x���<sn%A���7���c��
����ņ�@4�6�Kv(�~D��Q��p�:�6��0����G�-<ަ��;�ߕ��c+�q$����R	B��̼t�d"}�%L�b�e/Ȧ'�C�L�����\d�5�ɂ��7�?i�E���r8fe �p����d5�9�"�).)ĩ�gN�A�wEti�"�ϴ�
�|'��I:�{��D�8[�O
l��2�4�b]t��s������V{���	�Ś��$[��qP N�F���"�-�Θ˅�.�'�hy�?�X�9<Pb�V��5��j�bC�jd��Ix:�g�b��T��JI�DG0�L/X$qr�vk�x��e:��ȱ/��[ＤP@��*�Ҙ �����`ħJ�i#Q�އz���	?��stm�(4a�i���#�]{��yo�+kF����Ĉh����P0��q��)����+Z�YbF��>�1�1t��r�;�fn���y��������t[dX�;}�&�5܊��~ .�R	,�C�o��W&��T#̙ج>�G�����-�u�BN�<��1��s&�2�늓ǳ�q:'3��^6Y�4�P%�3�g���2�-)jӂ�P:�=���a��S̾@��V�E;��%{Rax�!+��<�' \��a�CJd��6[xp��ҜaI�K+��w���tр*��ӌ�,V�8��b2oQ,�@As��&�*C��(`�4���o�0_�4��� X#�np��*��j�� �}4���toTD�3��7�f[��M����n�e���&yb�)��ov��S�T�e��<� �1��
m����>���Z���Y����f=�gp�^1K��3>b}˗Y��8���=g@����ۭ<LX��V|9�7��=bՇ�ӄ����0@�d���a�]"��'�
[�qQ#4��~���ʃ!(jn��[��hFqc䔵+[�%[����p&�xKK�Os���a�JW�Sg�O&�˥����>��B�]��U]Ƣ^� �;bw]���by�fC0�V*.
Jw���	Fr V�xy��?��{���F��8��P��5T����?�,d��]�]�
4D�r_���Ũ,�|���z���dVØ��N4�6�u^p<*%��%�ɸ�꧲�j��N�v�\U�C�4
�ݭ`�7vH��T�<�_7ƱO&U_z\���{a������
�Pq>�0uŔypW�bg�N	׻���'j0��ռ57Q��[�M��O	�pV=��u�!�=���5�IU�Z��Ba�Ʀp�bz�[O�`.�3���w׻�	�oJ&h�8c�A_�H%4>�e���z����'>/�ɮq�����k1�,z�O Dڗ�z׼���=�[~��hl�p���.��Ǡ���*�50����G}�@�N�Z�9CĽ#��;{����=[8�c�T�l��T�#�G�T,�ЉlO,&�z�y��J�S�mbb~��fx*��V�ňx��34@��֏Pb�U{��ԹO��
>��AGݪ}wK���z�9����e�6:9�4zm%Q���(���-�@ļ�<,~;�����x�>tqW��[h9�Ӗ�A����>����}�j�;8n>�b���� r���_�[Ny�He ��Ĭ�ڳdc�04~\�С����m��'o��롛�� �%�����h�K���6���#���,+w�w9�)������������,A�u���^��W:�ja	�:����^	c�4X-J���A�Fo��/D���G�l9I+��ɖt��T����0@�O�ּ&Ni�2�ba�����3A����L��$���'�qdpԾ��)L��u��ܿ���&�lx�48~�۝M�����x́"���e�`$�ǀ	Z;C	�Xt�b���(�W��xX\�x3�J���z,5��+ܸ�U<Q��ګ�N����?-����j�h���٫���Yj���{p%���XL��b�Q'���ެ���B��։DR= {F���+�5 �6� ��V��o�K��vۺ`�¼O��Ki�FpT���@��ߙ��P�-�x�aPC3�ر���oD���	��w�揟�����f��W:o�`{haA���"�^I$��\�rz���K�j���\j����Q�n��g�&�}A;���G1bw@��5mc�{����/Ð�=���u~$<^�>E���� /x�Cr(�Lv��ߞ��z{QkG�'���:�*�dl� ��b�3?Gq��@{�w3�0p4Q�Z��Ѱ��S'�y9:x?)��0T��ڭ����4,��� ~S���8����=���d_ִL,?H�%�'^�"J��e��gr�B� ��s�W���2Dղ-�8q2����8m%+2�PMfA��j�R����(��B�S6�T�,���m�}�o.,�!(�;[�&�mM<�G���~K���9����'r: ���E�{��i@[_o�b����{k�~��Uy� M��`��[΃:���ٮ���t�A;`H3l��v(�(�K	���� �GI�'Q
ckM�`Ѱ?���X^נ�p�4ʹ��iK������o�ZP��0h��v$��	^���c���&�W�{�G����T9a@��M�R�x�R\i�3V�4��V�V��<:H���p�`=aw��a�?���7Z���w$1Eqd%1bkQ���뤡a�nF�S���`z�`o�A;p��!� ��;4t�P�E�$�7�B��u]ɡ�J[���x�O��d-ݗ�y��&sq�UKz�L.x��[e����}���u(�#R�B&�sg�ːX���l��"��ܣ�S�o��ҩ��*T+S���C���A/[]19:�&��5?�|�1�9��N��#��@x���b� ;�<gքqWf��Ȑw"�X^�0l'v���ы�F��lڗ�	�,fș"���/G�Wn*ݔ�u�h*]����O����?u���u�.��pc"Y$�O{s��;{�!����T-�INZ��:�\0�+�A!�,������P�1�<�eF���Ў�!Ѫ�b�~u�z�Vp�Q��_�K*�*�si����y-ۛZ����C�{�$���MV��º��[x�!X̻�jbٗ^H0�W�n���Sgw�;{"C[&�v���dM[�*�m�i�����j����Šg���,�Y��n�M��ET�اK�ˊ�Ə�&�t��c��x�Ȕ��A�|�}v��k ��P1n�@���Ӵ$!�f��(��b�+����鏾�F�ΤH��4�Q4�Bho�mZ&�B�8x��L��D�Od����:rW��Ԯ�P2]�������!�q8dԻ���|���CT3@�7��`�1@%���U���齈]�6�Db������"�ȻC�/i���Ƒ��X	jӝ#<C���6�����O���R�3���p �"�KI��e++��RO��}���L(:����ބ�j�R�=�i�_Q�m �"��
�O�p�C�d('Ob�Al�- ��"�Ĺt���ի֦�^U\Ē�<}W?�ͧ�1"�܅y�MLo3Jo�j��y�T�F!gq���m6�eJ���vA͇ ��@�lA
�������[�u�w[����zD�3�3U�V�b�W�0��|�4��&����z3TY IJd�B_���[�Z{�B�3pA�3�lc�<�M�swoA�tg�01��7ɿt��n<�kM�!����W/��ќ1�����Ւ�1�g�煮�:��m���J��b�MP��(�EoY������MW�=vp�^r)�ŔE�W�7.[�{������9��u�F��>!�&�8�2}vC�⽤S�ى�8�|��|7sׅ7{�2pL;5�:<�V��j	D8�Ϧ�L){G������
�'y�!����V�����F{���٭�ͮN;���̧%߮�>�]" �+���\�.��ă�-��K69t��kw��+�zdV2�|�5`�[:���\�b3i?����i=r�Ba
��m�z�o]H+ ���p����n��6���|�z\vx�m�G�x�����������4���϶/�N�����Wr���aCz��i�A�u�+�_x{CƼo�%N.��Y���U�/9�B(݉]s��n��U���y����[�ѣ�D���N�����!@��ӌ�r�6�x��G
��6�ay?Umi��"�g@�l���Bk�r{�� ,h��#�����;Ͳ��E��S`Z]S��c%�>�L}\:�߂lqֹ�C��9L��<{����:~��XM��/p�ȧ�5��x�I�� 8�W1��Xi'��>�@۵�(�Fbkn?�4Oy�8��=���Es%��DO�t������ﻐ��"4J���:�U�j�|�������t�Kv�� �X�7$S�Ba�������hp��/�Z2�~+�Ψ@݋�-����4��-+�9���s�c�Y��Y��Od3�<k,�V���.�F��~�)X��Ί_�? y��ܖ����H���"z�����m�t�?�j��]B���[�<�B�7 ��]E���S�F��~�:�"��֢��j���4��.yc�=�ߎ6b�l;�x�-��9�#sN��7R�T(��ʠ�q. ��>ʁH'�f�2���0589��a�S巂%E{��UZK5�/׮�������-@�m�DRX�x��"/�j�H�*(ｴ~���}��W�b��,�r�tAɃ)�XE��;@iȏ��ٛ�D��I;�$�O*�0����Rs���MQ�F��0��Wš����Ǟ�#z[�G�����a���D�����b2�Ѥa�߯D�I��o�Yš7�sc�Z��d&��KW��n�S�қB$�P��3h���Ƌ��#Hb�T1�\�pd(R�^2n��)�ЀV��[L^�n�'�+��q�����v4E��E��:�'�̷���`�f�Y{��O����js�)�y���!�T�5�6*�-֣�]�r��J���l�F�Ǣ������刽��@V���̣�����Ka1rJ�&I�oB�ǣ=W׎��&<���������R	�>:�u�l���l���|��|�N5}�������Q4�o��Uv�8��{`�����L\Q�Ϝr�,x�G�jv�Ilo�h���ފ@`�s+:��O�:�8�)�:<�`�9��+�l\�AJ�"Q�kl��2�.ۑ1{����߶�/���eD��$:�u�]V`�CJ��t�C(d���r��Q� "�E%��֌��M�Y��^�����FCqܽ^Ǳ�^�����Z�!�J'S:c$讖|��aY�A�r�Y~a��<	�1t���ߌb��6Q�2�nՏfXƘ�ƶw�P��	ic��K1� ��[�,�(��W�m�.�m+]�����>���xDڈ%¡��|����>�#V������8������|�=@�oZ3L��8�@֚�륦�%�%�n���W�T.[T��
9��;Е�����3�wo������r����9��)��\g�s-�a���w��^Pd]=�H@sԒ�����">�������kH͈�>�/��.���`���3r8v���P�3^KxB��l`��D&�X��u L��8S�5D�@��ך�?/�*\ �,����ܦϻ�=�F#6�����&ӊUR	J)�F��~�oІ?D᡼���l�>0�|�����l@_�_iR�	[;G����F6��aq�����΋��*d}��a��._sFu�h��V+z�1�/�&hq��m�d'�YDYU����,3���=q���?��AۛBă�"p�s�B�qUm�GOu�;��8fG��X�.��J�� ��.l�X�|̻�T&w�NB68��5�Gd@���Y�³�m}%������a<���c#>j��!_*��
��!�T;�P,Y
�Jlgق@��z�q�� C��d~_����A9��s;�O
�0�bF����x����f��=",D�q�Bi��a@���z��p�2m��=�rk�L��Q��+ꮲ��S�*X�|_
I#�x�P�f��QHςfaow�f�'�F���6�[H� 3U�w��gL`����*�l~+s��?�_�d%��=͘�TkJ(Y��Mt�d/�A� ��Aɶ���<���|/�D�~��n,�G�$47�G?Un�����d�����7�IU�9wq��X����=�v�3�_B��g�nV���#{hE6