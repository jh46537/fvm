��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��xzJ; !p�-�ߵt�Q�וi��L��:�� �k�=�!Rտ�ↈ������'IZ�m�#p��OW�@�^�f~&ߦ��|�@���	��Q�)O��0���<�;=߅�튃�O"I�t>>`�I����_�Y@0^Ğ6��U�*eE�I/� D~�|���+��0]2�yO]-'?~pg��f^l��J��=hD"��P��P,zjz���*3�h��WQm���I��[�rq�pV��<�%ƾz�u1��j��7!�k��)�a�+�hGe{�4a$z�&�O�J/`��o2D�=,���n�9��]t'����ӸF��mo�X�DE(�^�/1�W@�O�����<Tˈ	��A,ˍ�[]�T�N+�b8۸�	b�����9���ѓ~��r�
>y�7����U�T�}8��w2�:���y���==sX�y��?�g0.݀[8��K\���>��dD��s1)�c=�,Zw���ӆ���Ê^��%��^�,�n��I�2׼!/����}�C�gQ�;�D�_��
�̻�PӋ����>�bI�X�#cCX���!�
����w�:�
P�*��k�3�1���S��6Ҿ�j��Y$.u�*]�?=k�!,K�db3���p#X;�4��Ǟq!���l�{�7��#"���$��B^~�'��p�mp����ejI~��K;�kY���MI��=����i���֜�Oh���q>3��5����P�����jP��P]��#�qU_�	l�$d�Q6�	d���u���WO�7Q2�	�Կ�+���E��K����F.Q ����m��4Z:���⥽�D�Y73@�U3���՜m��e�2#�
�LҷO�&�:��0�SY�95O��4�`��$T��F��a�_���U���g�\�Wk�{
�H���C?���t�	n�r�� �d汕2��� �|n^�"J�uo������-�{���V;�d�����Q R���Ձ���n�S5�ȁ\�э;�����zڶ�;w�/��c���ҹe�9{�y��28B�Н�sR2"��tλ��Q�e�|I�Q��M���[��3�����"�q��9��3d
;{?��+�+�۔��)�E�#}�l��ow6ξ@�21����o�Yk��x�5���Y��pAS�0��٩�+���e��d��ZZ���opEY���LA2.YV�[G<�A����/c[ ?�
�N�F��s���+��ﹳL;80H����KSf/s�2\ 8�̑���H�?��o�O������?�>+[�ܗ��R�����K�	AH5'5sl0� ��ɝD�Zo�j�d�{A\�CL�ᱬ]��K����IN�d?"\��y�k��7����<'|�+��j�C���D��u	���F7�k p�ޭ7z_y*`�#K�[-��������D7$}�$�)'�]�A�	;s��3Lkݕ~���7����8�!��I���l��I��`-"��u63E�o�  ��㪽ʟv�р>|w�y�~F�(�����$�'"i��U}_:OU�����>�ڍ2�� ݹ*���pX�q�}q��<����0�����
�sfn��~�)��^�
m�-��%~ͫ��3ʳ����AM���4VL�^�R�C�]E
n*���܅�%
�*�Od�v�[c8f����0��9���_s��`s�����$�\����.=M��Rj/����ȵj�/�{�x�"��Υ�_��B0qI�$
��sofq�������`L��X�Xgz�,����h�o&����w3؟=8����i#N��C�r,���X�l� �l�>��<��������6U��k��[x�朏��l���r�h�+��u��bpx}V?��S��*����d�C����� �@�	n�c��K;\	]�6*�4J>/*(�m�iSl��w�1xQ�����&���5����:�1�k���ݭU���'�V�ԕxR�as� ��&dX���w@
\��џ��L+�n��	��ZIǞ�y���b����S�������݄��o��YBS@��
��p�Zi�2L�7kD���z���������«U�l��J�}t���K*�>Ț�����@��w��g�K,�-E�T	��#!g�=�n��=M��r�s}#�-���D�H1	Y�`b�Fď����zѓ�f�����ם&x5�j�����s	�}������S��0d{�p��I�Z�j�o,ρ�U�E���u�:���/�)�\͉����>\IF��2�>�)�R�#3X#����J��BχC�2�dJٳo���ͬ�2������iqg%낈�KN��)7��e�a�W�04H�>37r�D޶	b�,h�"jS�ª�:�=�n2���\&ep�'�?2醎���֔�MMZ<�E?J���`��0�:�Z=��)�80�@�o���{~=�����:��}��
�'�W:³�/>b�8��Ok��a��8�3�L�x�cX\���m���#[\��t`�.la>d�-2&�f����@wwɢbnw���0�a�jdY� ���T��zLY�L�Vn��\�g�/W�*0QM����� �ǽ�:����yS}�]\vOV��6��B�0SP��3k�W��!���rl�囉�]���^�!=��r�^���2.�Eۏ�v̰A 1t��W������c��h��W�[�Pa`%�w���=ӹ�ji�ⱽ�u�"�vq�R�"�i	p��'����v����e������$[(�W��z�{���=�+��T���CG��E�f$�]���R�g{ ��4y0�g���,~L�$��ӽ��,��(@m!���5#5��ZYӑ�5T�<L�!e�������qq&�i�1�bf��)��ݴ�Q��ts��$�<��G,D}����{t�Tg���U�
���L�΁h�m��=U�y�cӑ�p��	H�6	j�����QS�Ѽl.�� a7;��J��0�à!��.�� c1+*�.~�"Y?.��w;r��8׵o	�,�2P5U�9=/RЇ����Ib{���l!o0���@)8��;/����}���j̏���S�-��olT0���0eq!�Vѷ�/Sy�P������=Q�5�ɵ �Y�΂j[�Z
'�
OqlR��C��/Vk\��
S�q�u!�{Ǹ̲ɝ�JbZ��Y4.�%���C/x��A���v2���$%��_�ݾ����[��	,�.�C���G���آ�ֺZ���Q"���@��&�`����+]|�y��i���E8��`^��^B�k�b���3p�]$�/�v�Ҕy���`b�6�sG����t��q�\Z�����t���u�6����+"''K�������Lm"�Z;���&
��T[�eZ�ʻ_��%H�j�޳r|`�8Ls^��,��84 W�@z�z�h�ZK��C�/H�e�]
�b
ޔ�=���CbZv�ˁ���򥞓�B�)+E
o�9�i1����i���S&�dG�`k'a�Ư�
�g|CpXuP+)���gH��|>�I`.Wry������yRl�	��o��~��V�a�v�%d�H-�_t���@	jw1����s�ԟ(��W�o��J�e��|�:�<,�wc	EN�PA�u�����|�qR�����RxU��?(�{6���*����_⻁�ٻ6J��L���df�V�B<:Oܫ5�]8�ʿ0������n�m6�Pޠ����7H�l,�t��:���3��I��,���S��-mRm��������9���_Ez� ��r���B�<��s�/�Al�8d����y�jt~�jA#�e���U�5���{fS4.�_gdK;koC�a�g��ǲ�dOX@A :T�
-6�eM�,b�Y���_��`����H��.��9?J����zؤ}>RsT�=m7�z�Rߏh�� ;z���A���ݫɗ��`��٧�߾\��2��:��m��b�C��c>
<��FT�Im�դY�wN�
��YϮ.���I	Y�[:�R�(H�b�
|�$�CO�ƾ�1��i� ���Ln�P�[��g�	^+Ō�[``J�6�ǫ�G F.g9�y�cU� ���Ms�w�������2(�2�E���>�d��u҃��
L��
�Q�B4�WT�<���%�8���E;:��8=��1ң�
L�@�cf@K3 ��bBiE5B���6%�m�e�z۷%��]~�5nf�ĕ�-�' ����yt��l�H��� �~:�#�I���RQ��]8d��-�]�X���_�*��}�v9#��<ٕ~G�y-RL剆�5�+oW[�mp�+O�m���TH;�>v\�Ƅc����I�p�`�:�W�1Wc�L2�1��.�0��qp�
0�K�ִ�RbBəc��Ĩ�f?T	��q�O��Q��*!��C��!�UCBgD��tg�
��M�I�H����A�UŌ[ ���e��F�"4�$5�W�Fm�H^���B:`��B\e�L%[���J`<//��r���O�h��\7� ��,6��j�n��ǆ��6���;�Bl��D�_j�Y �y�L�A�YnnM�	�,TH1��@V�q�������P�"��Q'|E~(�@�����G�^����j�h�zE.�](��_����ɑ���N�pMj3��B��5�k"ů��=�e4�15�q��iAp{�-J(^H�H!������FqS�����j��~���~�9�Z1��q&RQ�����_�D'��&�>��8���;�QGJ$�2۹�����&��~�u�n��?]�n��Tq�/�Tf�I$w]Yե�b2�ŃX���)���;^J('I�^zP��F�-n�W@�$���e5��*a�#��ћV�`wVP<��BX"��Hu+��u��*8���g?��G�
)��q�04�� ���r�,�b��
2�0�����j��d
3���!'��!���u�[�Y�T,d�5��NJ�l���k�4-��>���[�76}��b;X�;Sn�/?��<�-o�Ti��@6�kj��e!7�H�%������2�=�=��.t0e>Cu��\��ڠM%���Ѭ�r�z�M��#̷c6�'t��{�P�A2r$��Z��6q?�z]��1�~��Bn������*�w��=z�;�u�S���b7��������SS�ͱ���DT���(^�_^��u�w*��^]�U��É}27�)Z�����$�N-5���O��!o��j
�ٟ��2�\��.���$�Yt]0��İ��uF���ɇ���9|�54�;Ց^|�)��O�a~�H_J��m��;��G�Ĕ��\��Hb���[V��8)�$0�c���}�N��q@�t�0xY�a����SB/�^YB3	����T����-��y�,5�ɇ��� 
߆#���]�,�PO�yQA�f���(�٘;��W�B�#8y���4��,���'��R �B@�����CC��%��Aw��$���%M_dR��Fk,cd�۶�Fo
��9�aA�Y��yX�_��%[^��w�%�<��kuԦ�	On�n)Lфw͎.(�Nk�.��V�(�6���#j$C�?	�+д%n+�X<n�BB��/X��glo-��]U�~յ��tϠl�G��r<乽�������a,��8ЖvKW���`�M�:Ϫ�+���U���"���f�Db��%OӦ�>PTݜѭy!� "��f?��|��H�H�hZ,���o�_2I\�c�^�����4B����f gSE0W��(é�������Ċ��^��9�И�n!�*�p��3�4��V6B!}����W'h�_Eo9o:��V�v����W^]
���
 �{0�E���/�kY��q���t����j�>��1#z�N�X��Bu�ų���5�;x�F����k1�ը�H�YƳ������R��WX��e�ڧCq8A�%�Q8���7�t�e�ϧ��:?����LH�f�t����S��2����S����q�f|_�C���l�:mԘ[>|����X����C���n�k2���41�e��|Yz
/ʅ����XETf�T��j'P`LFhvf���Z���t) ��glm΃h"vp-A��E��"wJ?/�魅□�����`(��/�|������$a%Y�8�ǒ�x�
T�Sa��2~(}?� A*��r��n��)�ȯ%�ޘ�����;��i�y�ծ7c��j�+�_���O˱�b�S
�J�]Y�H�!�v�(��G�9� P^x��Ɏ��ث"��P�&0^ �{��d;ë8��6�A�'��"YiH����q=r�۴��2�.n�x0#g�bo$^c��}�I����)}<�	i�B����BR�&x�dAk��ȷ�f�P#љZ�gd�p�	�%f2�S�05s��4�ZuPaJ���������q��>�X���b�����P��0�/5Lj=�^�)#�vd�T���:��"��|r����9,�������k��-w�@%��R�X\���\9�KxsU��_;��(����=0��@l�\RDm ъ]K#z�6XB�,���"�@���K*�ߖ5:�c�������	�[�æ�/B�g�D�:T)cO�e�;�ݏUd�S�;�XKM��7�[(3Ne���kf����2�v��O��Mv��TP��C*ѹ�ˁ�-�g�+�v-9�;�pơ���W�t} �"t���*B:<-�nc g�Y�=h{g��)�Z�7M9����
,a���O�T�%��_\�C�QT!��im�WR���P�wR�l�Q4Q�k��m�Dg����~���c"��T�c��CTǩ�p4�Nedq2!5���I��`��T�����Z�e���r���t�K��5���~����j�~4���H�ꁱM��mdgd6S��f�-�CV�vG9 y4�2�;C%�/���ޥv47m�ؠb�r�l�m"�,ߘ���om�ufy�"����1,�ͿޤZ62���>[؇0��i|O�ߪ���G.r�+A�z��������,J�����sH>\���m�H��� g�.��C�[������Gjɕ��K�|�|~I<bo$:�^�x�\~T9���6��<�Ï��w�*�di�n)YI��<e�Vм�D��e:9j"���P��Bi�5,��C��vw���.�S�r�j�.GR�Ľ����/ċUi��󛻽�����NS6�Zƾ�p�0������=�ʦ�P1
�P�F?o�e���l�y��Sx��NHk��Q'�\���T�'v��>*�n���  S9T����N=c�� �;R��5*���
�݁����X�\����'����M��]X0?/����,��EN��H�x �����п�2�@�� ��ѐ��0��<G�&7�bvF=`���\-|��,j��(����'�������"�2i�rD�".(I�Y�,ٕLJ�	��'{W ήZ�ϚռO��*�:���vBO#��O��1?�G�<.?�ؽ)�CT z���V�����( ��x�������a ��{G��iL�J�#��h�X���Eٺ|��w��H�6 S��^Ep���Y���G$%��gZ�Ќq�B��]4����6[?���9�4�$�C��"�K��~8�N�7h:A�h�A^��tY��X�Q+��
U9c�j���E�����X�$  Α��/cb�5�r&���%R�=l�o �x� "�Q�nQ0@�Y�^�? Sl�iY\���;�?��9(���w/K��_�D�xY��~E���%g}x�'���Bk,0��;i!Y�>̛	�D���D1>�9g�f�TD��R?�l]jpL� ���C~Є�hVn�-�V� @yZ@'�b��]�oeZJ����Kq�z����MN�U��^�j�I�E'��Fu_���n����@�6� w@��RjS�k�9�٤*�:��#I��8����+�i�_�dXO}����-C@�S�5�pk�5�Щ?�����v��=�xV� [�1G������N$�Lþe��
b� � ���f��W��a��I��f>���@_<ךp�"��4~Ր_� �\��p ࣝڄ�ʼ%�<E�L%�;p��L�LYɜC�e��Y7�������E�jW~��C�ˬ��"�=U�Q^{M}��,o���p���?A���@�Q����7�.J��s��8	6�[�<�]�oӟ�`N���y��	��Ĝdoe��1w{�8|�.�~~1���䬐����׶M�N�j�(����]r{�]*h��Var``
�^W͉Lf��pļ�/�}�̌�%.r�!s�8�_|�~�&X,cM)�e�����t�����KKz�Z�b�l<E��t� tۇ����$�cD5e1��'.#g#W#s����y��e@����%��`".3%�u�u3���s�������to��>?;α����1�d�żM>nW?�S4p�W���K=ۥ��j~@e�f���,ȸ7�[�v���-�h,c�8�I>����pL� �%�j���a��p����W�]����i��9WQH .��	�k%�E#yy��u�n [G�4s�X�����o�D��Uô.4T�`6�-� ��B}�T2�-G������^Y�������arB�)�0(&���z�
�;@}�,�\9���j��|%�SJT���\d
�Mv�v�A�AybE#f�YO%�k����LF���z��p�?6���?���/�a.1P����~�F��o%(�ЊQ��8ߟa�����kV�\tjw\P�Ҫ%g����v]3�xQ�1T�u�K������«���'c��������g@h�	,��/�8��F1�3�u�
}�ӻ w'`�j\lGo���w����5�pZT�b!v����E���몪ׄ8!$��ƨRJLr>�y[3�QQ�EC����f�
;�r�9m���@�#��o-�9���4_���֓�XO̔��gc�}֗��Ƒ)U��Q\ZFE��KטFs�/�C��ϐ�u����1+�	�6��F�Ň{�����9�k�������/�4�������:��4Y1_0�Q�[���!J�
���*��W�`�&p���8�zw�������~��H͑�j�bT?��%驼BxFL�h�?�T�P�B���?H��s�h:�0�Igګ��\v�.��dr�Q�L��~�J�!����F�&Ol�B*˨�ZƏ�{� J��}oni'��߱��[A �[Iz�%j��^	�#��s�_ӊ�K*���ռ��ݏhx/<h
HK����~o����V�L/���v���X5SBu��*�����Y�˦,Uy=���Y�ЄKEBQC(�AZP����ڝ��p��i������ʊ�tQ���Ճ��&��-/�d7���nw�N��]�<�{Lp�vl��L�8hd~�H��������fƩ�[�KA������˅(�B����`-��PÔ�#�~?	uI�(CG�?fƂ6\}���v�P����S7wh�'��Y��_�=:�,�w"�.�y�-9��p�~���´�S�O]�$z�Rԉ�m��a�������Nhs�l��/z+P.V�w B�]A>J*��X?ؑ�;O����X��{`�l[���2�8�i�wn�����nD�Vc@��Jz��%���݀�^�4����DY��KX�CqQ�T[J'����Z�����[�r��;��ũ�X;#�_���T�D)=��Ċ���g��pyCm�3�a�a ���3�����ܙ|��$U/�-<mҫ�7/���bP�ng�6�l8���a�FS��H}�u�y��<I;�l ��/=�������i5A����m&�A[m�w�<�}������H�W��6A�4)�0C���*�X�_����L.���]I�"@r���Y	��mA?����*�-�EG]M<Q^AR����	�[�ό61W&�r�#�`�5�âK3&�K����D���Bx����@[��t^,��k�qH�>-\~h"��]>}@u�br_����Z9���Z�� �mɿ��W��E��Z�?o�Oo��]��e�@w/�G���&�/��ֹ�2��^!1.Y6������t��>�PeR���I�T�8q�j��>Ou[��h�YQ9��֥���pܲ�	Uv���t�ڔY����(I��ʵQi$@e#��Ӧ@!�:��s.vI%�!��(0&)��DS���?Q.�5��W�F|Z��`��L�+�P�[^�נ����}�s�d�V�Bv��U`��<ƴ��`��^���m�6�H�L����O�V��$K�N�������(,��&b�K��#X#��58x<����j�ǘ����!�1��ȥ���ۧ�L����0iK��c=���|б��-V�U�
è��T�f��.	�^�`�I�j��-ƌ�y�BC�\|	� �=����u(�&$�C�f;�m��Ɏw���M~�P�<[�
XYC�U��R�_2b m�D;4�!&Ӽ��_>�6��M���f����V��p��_L��}��;m�:�<�c�Q_�C�>DФ�
<YF,�qA��\�[�\��`Ԃ��zJ��k���=[�tg��3����2�mk�:�ח�-�v�9�PP����b㎥���&H�?[seՙn��ÿ�P��[�to
jˍаl�'����k��.����z�堙�1��Z~��Զ���T,��(�RSX����.�lc�tC|��5�q�x����7{q��,���<ͮF��=I�ܳ�����/
2��t�v_�ꭴ4%�"W ���dz8�tW����q���D���̈́/�\n�>�JP��H#�>�?��]����+��4 �C�q攴7�	i��ii�eX.S�r%��%�^�xU�_7ʯ'Z�yV�X�IN���6�~� ����7����R��0U�0|
�����UX�ߏ�x�V�{wqp�k5�L��82J�'הt�# �ZF3��%��`�k�FCG���b ��5���F����+:�_q�I�����$���J��W�^Du}�����ȣ}��9�~��c߱}���))�xk�/<����8)��F`Ί��S�wx��!�o\�՜��;���(�p~$&�;�#�}�͒5օխc��Q�Ʃ���(��j$屙"����(�Pb�b%߹G�ȍ=�S�$p�S�͌�d���w�|��F\�
Yσ���f�Z��Z��#bb<�Ǝ��Vױ:+��6�/荸t��JL��>c/�>v���9�^����Q�^*ƪ�d-��j�91�� j6M��o�I���9"�$P&���{��W�i (Rϑ����&f":/��Y�{�XB�:p6C�3tf���Z��'!@���*(5��&|Q���ڲ�r�k˄��ɡ/~��<(�_��8`S�<��Fm����F'�֒*Gk?�Xij�Y��n�XM�UD�9
� ��a�R˕mfa�hf�(jR]�+"�:GQ�R�&N�F�Y�"}��tH,��TG���M���8��B4m���R5��ԇf��
إZO��c]� H��d�"�O9�^�P�������,�j���s$6��T-<�+3������RYW�͍�b��Ft���܃�
�4"v���Y��Y9kQ��#�0pZ)|V1Na�����!�U�������ȳ2[C�����Ȏ>���@�2m�Jeǯ���fd����U��G���D�f�z?ńVX;�A�TV�d�0:���h��-ڃ�}.���P�V�^7jx��9|��7-N6���P#�Dl!^�V� Yy�&o��Z�vj$lhb�|��SU���|g��sZP�~������_��9�!��R���F��	,�.��2�a�e������glkgM�`�������X�B0��������� ��B�Jk��c��>}�"uݴ�����+��y��4���Ǖ5�<�
��O��0c� �Mg�`�_E��ٵ^�MP?zݭ��t	k��_07��o]�������V�� .���3p�-�D��x[�^���$K]S���,�O��S�#����`+���	�c��rK�H݂0�4i�Ͽ� M5��)�$�Hz�v"[��.6fū������{ ��,�f��4PJ�~�M�͍畴&�lt5���K���N2+��ɯ�MFk�&E������
�%B��4Oba��2��v���4v����
R( �����%���*��NbT�Y���[�h^���9T�;�p��ڎ�kk���@�1�r}Z�;m�&���\ʧ ��4`�K���Qg���V�⅗^����E�{�����>����va}�p��<X���`c|6D�K�v�xEC�P�q�������z��x�i�훣��B�OM�C0�o�c��w��1��nF+��<�c�XKJF�K�Fy��e��?S<o9ܰ]�%�#s�뫋�cb�� ��;1��7�JJ/ix�0	��V����ofGZc���߄\��U���0; �훑C��RT�,�>��\�K�?��� 7}V�]��:v��oKMj����-@qi���e%aZDZs�׎��h��7��;GH�
q[����+���� S�'a��^�8�+o�jG개���4�E�\z�x� ����?� 1F���j���%�h#���es��>��Y,hҊ�U,���,8^���	PJ���T7�����w���,*ye���z0F,��G3�����
*�?������F7����{#���(����y�²o]Ɔ7��(��|��:�t��ϝD�).=�x���@�r��ZuC֢ab�޵_R9[QX�Yhq34��(W8ʾ)x�,$���Х��RV�N��+�d��`C���*�vn��9\���t�����$�k-q�P�����+`�G�b6籌$�*U��$��bV�r�f�E�z[m2�)����>e��נ���)n ?_Ɓ�=	�y��6ZJqibb�~a�`Y*���YIh��;Sm�I��kr) EW�F"y�'K�X?§�d� �_x�%5�2�C��0�k��+a�B���z1�OCU�P�YE8n�6����9@�Xl��{�l[�.%WP���DyJB���gY�VRS$��0��!�R�E��
G"V{��Դ&�?�������!G`�0p�KC����m�?��R�]�`�Ch�9��@X�'/�I�� ��u4nҕ�??�����:�:K�A��m��ʿ��kE�,�,*�n��5K�q�d8�!Ջ���q�O.\2"~dcG�}΄|��x�Ԓ	I�n�֢��8[��b����M��D��K�&�V@�y��F�I�ތX���g��;5��Q��U��&}d�z���yq�L�[wJe����loJ��A)'�]z����R�P�R��N�n7��G�}�����v���g6ߛ� �K�tZ �j���Ld������V~O�&���'J�H�1�vtTҳ�	�OX�L=dC++Lk�+R��1�l9C2aLW���"�J�e�R����?j'e�푓>fk��X6nL�U���(���λP�]�w�c}S*��N��^�Wl�J�VC�'����#�
Q�aпш|�Ȁv���<�<ST3�G�xx����{���0�BQ�v�ۋS��>�LT�522� �1�v�Զ����I���l2���U)�����B�G�Cĸ�
���[C�35Ŧ���3g����bvZ�!;b�?���)u̞����sS���X�+�>`�����L>~Ç�*l��x)�]��v3~�Y&�uȯ�.	��"z�}���'�
`��3��ld��<!��{�إ�z8�i|�c���B����ˑ`j���I� ݥ���Z&OX�)tt��L$P�g�Ac����2�Lw��nxk�m2�Vu�B�H��9�|��y�m漜���]f�9�?����#�ۘ�h�%A��UN���O=E �ĩ�,�����O#})\+H�)������r�	��H}�p�����]�?|q�|��ɒ���6��hŁ�\�Y�;�jz�Ax�~Ȕw0�R������O��X%QW� hx�����˵��X�������1 B�;2��u��}�"4����.����*���U���pV_)�ˬ����&��h�.��!IЮx����r/L,l8*�1�:��䫎�~�C�bf��U�H
K3,�2�t-c�?�)�V7Ii��Ơg�Z�1�hJb������h�'>�����֠jU���wɇ���ry����Y�u�=v㖈K�D
�CFbz��؟�fYj�N`��dw�d?��]WnS�Az!�U|�R*�c%���GSȴY�h8MC����<L����?�����EG��d�󗭵C�:Pd_!���
�0��2�=ti=�����F��F?����R��*��������ڨ�f��� ��g���8'�u�06��N٥BY��N
�5�a NS��EOM�VFU1ikU�o��e�5
#��QGd߶O���|�S��ƾ�:0�R�6LM���o����@}�ݶ_(榉� [�1[�rW�
ƈ?}ZC��CK���j�������+y�=�6�.���9�O�����^Ձ��m�pb���؃�|@�d"|4�:��G��p�h��O����0eϱ�H��ݶ"%� �1kOy����lt�<a�����d $et�TF-��9���s�?r&3=���Di~3�{�XGb	�A���@LXDq�
��͕�۷���0�i�#�.�PSU��==k���hqLQ�R�d���2݈��d�[A��~|�2�
��W�(�|�&>���W��(⧼w��Y	��C�l���`���E+��������&���~G�)������d�u��D�b6̺�Fu�T�L��ld%���������qze�7!����7�n������ \�˩4S�)���ނ�_�Y��)_Du"#�@V��5⬺�@����vD#z^�w0S}�q.rf�_�F>�ji_�o��v����o,1���t?^}&�?z�g�HQ$=�����,__'��K�P	>�����(��L�l7#~�����Ɲ�d�z��vId��o;Ldw���;X�pEk+�bR��`Gض��2�Oh��P���:�p,�^L�����$L&>���/GY�y�uH}��L��-�x�'k�t@�6�%�����G�t�#�9=�M��O6�{�n��H[��6F_Ɩ�W��"��r��RZ�	������9e�`��m2���{e�2���R��@�
Gi� ̹�=�o�C/i�y���}>��m�����IJ}���tFq�ݍ��8x�柔����̪G�D���uz��� (lf��zGF74���MsS=f��3�kt�.-j���S�������j�[��M��$�!��+�H�Z��@�S�u	poy@{���K+��o-����/�O�9:ѩ�0h6�,S%q��0���k�6,"6'����Y�Z��&������3
.��S�i���s>�ej���/4�FH���J����,���}��盼�뫩 ����?�X-۲�˗��L@��1dA>����rV{J�cEZ�&
F�j� V��CG��s��٨ڊEi�d�#v�@H���pqyЌ ��rᔮ��
XK82�	�Y9�l�
�q><xA����������K�:��i��BO�T����ڏ��0�Ҍtג���6 �#/u��Y�ڡ(iG�\W�Gp)޸ۄ��c���l�r��a����ߓ�eW���ەw�`Q ���u��en��������Q5�8��v�Jk�;��e���R,����=T\I;+�%��>'�]��NKg/����xy4�j�=��<��rT�vZ/�|օ���̰��"녱mT򏛊SM6o�H=��Ꝯ���A�!H�t�Q�OZ������>SX�l���{>�4�vW�:��.� W-���;�\�����=�-)��n��	4��X���Q-565ވz�@����?�~��M��f\xX`�"W<S��i:�K����|�b�	,I(��C=<��:dg�g$�F>����P�Y*�)�⓿C%�Ld_N�aK��<n���I�=(+)��hΊT�gj�Vv#�+�5*��Ʀ�`*)i��a��i�NK A�=�W��ۊż��_8�H��k9J-��3|�ycY�}TSb덝"�.a�z-#z�?,m�1��u����C��S�R�ű��-�_��	��S��e�(�p�ʥ��������~ČRQ<�@�(�Ò��� 	���X%��o�s~T�N����L0=np[�]zN���y���y�bm�K5����?�W!��5���]B:��=8V����ē�!L��{���;���x9������6c���	c0� 2�g��<_�oS���L��R(̈<b\Q�VukSp���o(��R���h*,��A�r2g�� ˓�tD�_�>�=;�Vk�l�Eo�cE�۟���!
�����g^>�MF6��y�-+|�L䡥o�x���P�+��T��.Z�&��ߢ9�T�q��}�� ����	4����M�@�tǽ�ڢ5�rㆦ?��gI��uN���=ݠH��3��B9�����lNSѵ<���Z�b�=�)���e&�`�9j"�y��~'�PR�c\�=+����A	2`��bƇ��8�fx���ms�ױ_�B(v�w��7M}�� �hV�"MEF��q��:����KG8`q�~|Iz Ow���J0yѵ P���?9�����w@p����U�ϞD��QQ-�Ϩ=��au�$�������9Z-=�$%T
��ErU�J8�J�{X�i診#[-1���85��2���(9ܯ�{����(��\�˗��iQP����;&�^5�j_��֌�ًk��.�A����5�9L�&4���J��ɤaP=
��8�~f��FE�^-SHU� t�-�����|n���c���\eڼs����v>���Ȼ{��٪)��+D]JM#=,���w�Z��u�8͇V�_fë�~HfJk'������6q��DNBI0Uv����p�N5���/P"��T"�@����4�G)	�)(�"Xj���<NN�K���=�iF�����-��4~�wY.Ĺ��E����6�c/p�u9�?�9�ȇ�A~�މ
�>���1�"�@��RLOwThܼ��{�>z_ƭF>OX�b(9A���k`�>�>�-�EH�]V�6��1s��@���M6��9ި(oA	��!�������.6�E�\��ߨ�݉C���/&5�%�����֬��Nw�9ͳ�&P��p����xݦe��I�����G������1��5�̐,�ٹuT�?��'А� �M������x �(�I*j��f�Fڟc>H,�OPty_@�[R%"5�8^�o4��I������3��61B�����,+�hy��2�3��a4������(����;Q��J~NF4���㾒#]�� ��J@��e%ɶф[�R �~ge���y2�Ơ���
�	@}��/��AeD4u��ptL_�B��`�.�"������?�m~Hg��r0�B��?e;X�!2�OM
���d���X�,Ȥ������^��D���x��3������ Vu�A�MG~��0U�ed�YĔ�e��@������`���i(����4�"ݰ� ¹�����6�'�� ��Q�����-�6��(>�nFQׂ(������mNى��yCUDQ�1'6��#��X�=�S7��}�D8Y�@(:�:#�Xhڽ|b��
�4|�򍅦Z�C.�����9"�4��?lY�f��I�w�y���岃v�[!E�YKS��c��/��j��߽��J=��r컍*���etm<�D,ck��KON9i)u8GR��0�g���Z{���̱^���ȥ�mr-��*�㮱
q{���x>!<4��>wQ�p�3�2s�"��{��24�9��h@����(���j�n�T=�E_ݝ�� �e��N_jc���VN0�G��O����"�M~��f�O��:,�?e�� �Kt�Y����a�>��!#fWڪ�l p(���#hv	�`%�9�ɷj�"���l���u��h�栄-mGV�e��@�����Y��\ؖ��n>�~��ͧ�H�D)��⣩�����Rc�f	�`���s:���X�Yg�ӑcT�{��G���8��	�5��/zi���cB
!Ul��Q�w�:@��d�~E��?h��j<�8�F�T�q�3�;[�	�'3����������8i�>�N�7���%@�k1z�1R92��2�"�)�u�{���Qc�����0�)�X����9�]�ݜ��k��f�j��9m�)�����#궥6����D3+ݶj�S�ɐ�|�׎����Ҧw�@��
�&�bP��|�y��,����'�n��IET�����n�ΎU|����'�Q�4#�g
/�Y^���Z��7_�Y��E�5J5�5��3�Y���3�L�n�L��wG��'��R\^�.@@DA�.	��)5Ӹ���#���hs.��.���u���w��}�Q��`��5 �x:����mj��\A�K|9�ŉ�P����Dє�t�'���8#3�2��\���������,��Gd�`z�0c�^?VK�y8.Z�'�7�Ǽ���n�f�v���s�[Ϟ�]�B�.�³�Y��4xN��#d�ČN�>#Q�	�,���Tf��Coǌ�o������[��ѥ�]��Bl�+�
<Q�NQ�χ������9�V�@0ɬ	�� G B�Q��"�zG�!��\!��^y@�r��!�<��gl@�f��Ye�t�v�67��r�bw�Q����j,X-y�#U�Ϳ�ƙ��N�v�)+#���o-В�F�/TL�\X�~	�,�y�W������ϬKx2'%�s��D#�ӑ�*}�������~�,v:\PbWkp�n.:E�I����0#��ya&�4]�zȔp����"[�wT�s9,��W�u۳�d
�h�(2�ܐ�T5z�;/\y:�5���V���N��d	x�U()��+�n�*�V����/��<T�8�6����F�kp�F�$L?�%�cd����.����߻�=��@(����~
�eSGn��5��֥�d1*� _�_#�I|���F)>C4v��Ko��!�M
�:XF��w[V�^ת�_^q5�c�y���B@��`w��Wõ����o�:�qy"�*s�3Rg;hB���;ss��ď��2���0�����$B�g~�e&����;��[Xj�6�G���_���y簼����>��z�BA+����[��l]�Ges����zG�'�����r�nJ؇��`�XѼ���z�Z5�,>�O�T��Y� �<�|�J���c�R% �Ω϶�얖�V�XE6�@2V��\#�q4>���Nqb�} �7�+� ��Yq�|�v��7���V�Μ���>ٴ;��ܪ�:�=�:ʵ�pK������ o\e����&�oZ�Np����u�R��F�n�Z�[#�2O����P�S����MO�x��f,ϔ�C&W��{�-[�̽�H����T���I>3��C���@2$I��~��y$\��-F�#�������?��,�Yw���~���̰�NQ���+W�(��Fq^��q8.� ��n��'�ֺ����P?��S�ܵ'�b��@��3��ű��d*�_��/I���b���$nC���R��mCHl,ř�����΃�ǩNb�.�� ѓ���b~�'���"�{�4�LM_2�㸿�g�R����=2���
��(�b?Hũ��J�r}IAN�ľ���_w8���Y���%uZ72���R���V��`�^Km�)1�՘����T�
+�#i�dB��� ��K��*`޻��o����_�gF,�*���!�O�p�ԑO��'�c&F �!���V�=�)H��n
���0��2P�	�����pi|�y�0������`SR�I�v7��<L`�f��#UĳD�����l2�E5*���:�ۖ)���%��_��N�J�#��n�� �)�h��.�<{l�,vQy(1P���U�.�Cl�S���� �:�Ǚ������>���y"�d����fա�ck|�!B�	������P-��E;D5\@��K��}���*,ȶ���ƻ�b����1��c�Nb�J������Ar0q��q�`���J�`��b�x�3P���Ά�[<�dm#�|��6 9P��Q��ʨ�^q�qlx��L���GX0j���]���D+޴>�ī��*�h�;+��d�#L�N��ϴ`+���,��֓s�{���'���Cz���y�����;j)V�8�e���V�TP.?�k�I�V
tH�-��i�1����E����!��v��!wθV�7���f�(A��5Ѭ��A���"0�z��؈�q܉��r2F��蘥-��d�������zޚ�|Ej�?a3�@�ŗF��R��i� ��7�[?]������ 5��hhF���	����kJ:2�=����޼��A�:������%*�Y�^J`�����0c���z<]�+�t:��ɂ6�A��� &��_B̗�7�W�s9�G��u Q���8<ź��#6\B�ل��B����=���[5Y͕����L2����wb�y��f��"��'>1 �P"3�J���%�u<��R�L ��s��2]B�]�����E�O��Mb�s��uz$G��R�5ٰ��:Q:�[3�LuE�K��.�	�w�M�Z|�l�{�%��D_E�x�:�5Wuu�8��r7HU0Ʌ�4�͝wˇ�zk�:�9������XÉ��#��N	�����9x1iyƂ����tBEp6I۹�z|b@6�t��:_�9�������������"��0���߫�o̪��e5������(����������Ϟ���0@۳�dw�=X� ���'�w�آ>�6n��0�I_����y׫C 6O#������j�~kOs��$�bQ
&�HՈ����_X�RX�� ����H)�\��G�����
)�"���m'��Q�ou���F���g�{,���J��qn)\Aܲe�6#N%@��i9	^a��29Yͱ�1Z'��ʩ�l`�c�壏��OG�s�$D��#��ps�_�����z�R��1 �o{��T�Ɩ�[�ϯH��۴��|z����d`�$�������o�ţ<@�7Tv~lœ� ���_��}�����7��?�[t�W&j��.W���)neT�~4�G�����Z��\�W��/a�Jp�,�� u	�㤣�q�n�0�pv�k�(�C��K�N����
LK�B�1!�l%,�_+N}�F7���Q|�WS�f��څe���%�7�	��T0�� ,���ͱ��ߗXƇ�#�AP�.ܬ^�7�Y��SZ�� �3�`�.sKGX���L<7��w��y�j��n�e�6"�e��ٽ}����`-�'+�?�R���N)�.b�o���A�9R���9� ����4�#���EF�Y�l{�73v%���S(/�����l��ދ��K�O;hL�=��X��5��ӽ�9X�7��cj�<�Xʅ����z�.���������]=�A���pT)���9�q0��u|#p�rX�L��>K����k�`���}1�*���q ��sC�2|��A:?���I3����ق^�p�ac�]%��\v����ob4��-&�]���ą�97�����>��D�d�
U���L�k:H�K�<���M�=��U���M����:��j0a��9�Tx�W��bR#ؚ��i�Q/r�-�ߡ�C�l�s�HH�l��k�`�]�ί� �]bT�M�V���͜���쒡ςqE߲��y�+��sj���_[�{(���H ����^�pE9��@Ͱ�j��L�uO�_�p�,h�2�x]
yW�/� ��~��JХи�k�,XCD]�:�Q�*�Bz�DzÖ�i�9Vߕ)*�����%��ׄa�}��@ؖ�whvP�"�\ZW��愪v��q�*��'m���j
a�����?c
e���{���!��]���,� ڒ l��J	�.%E~�p��1Z�!�2���R�|t\���r�a����A��g8U*V�?�@�;#
R~v�K�V+,���$�������n�do��2}��q�.=��U�YBT�H���BO���ľop)��Gޮ����za�t�����H�S���(����J�[ǅ[�e�3O&��@���Z���
��	��{W9ǅ�t���t�
�ʝ'K;��_~G��u[�
�j
E���xk�9�![���U�|�9	\_$%j'�������@E�ߓ�L�3%�+��[װ���^|����)�g��T+�*G6o���O��v�~�ÿ�^�;1�BM�Z��*z���.�`��jd�N�Ȱ��y@Z��^iN�n�L���^w�����x��]�����t[51a�6w���;v�D�W-z�`:u��~��H�[��M⎉*q��W4�{C7�������� *��K\1Iq�<�	�7���[���BeF���ǵ����2��J����'!%�{��a���5�tH�z�Ik�}��`�D ��`�p~���"L�����f ?��D�Gf]��[l��O��� *���~��b)J�M<\Ǧ�����Ԣ�z�Q�+�"fV��.��@��A~E���'E���w��Q:���o5'k��u��-o$a���6�_o3�L`X��ɢC~>	{
��: 4v$���V��R�՟p~ų���8���ua��G4���:X&��R��p~yLR;�R�b�����©���tx�?�*��
� $D�E�K�p�vO�������~@�Z�K+����}>�s�A��
�+�j@�5�gH�5�ey�8[�_�Wi��2�^�����X��|�a�y??IX�i#��}���/�q�gXL�]��g�H*q��pF�<�����q���D1�A�Y	�����`zF�����M��AC�_��i0�d��"Y���S��U�;4�q��Vt�$>�S�.�D�1U�*
iV�'��L�=E(��NcPYO�V7�<�0� 5Ma4*�N�u� ����Q����Ζj��,�`9�3"��^SZ1�-LB�hk� p��]���Hؚ*�n#%��~0^�_�I��Ċ�ͥ�ԫ�>��:�@sv��2��;Y��#�4i�EL��#���.2K66��<ή��)�m�
J:��Mn����|n�=�G�dj1�J�f���6���D�͹�,��{��A�%n�a�:��d�����17� !Uf4������cY�'e$ �&K�W�FW�cY�w��zX1XK�#�/N���$`���wc<�� l�8��<�2=~��!��񓠱Q4'����U��a�_@�Y�;3�x5$Z?2�;}��!��+R����\��P�^i��=�>�mJ`�h�H)D��$�]F�L�u�����1z����8Ӗ�K<���q+l	n��@8Ν"�w��w����s�r���<�$��X}��샂=˪�cx����{0�־�f�Nk�����q���é�Y��v��n�UjW(���W0`U����X��Lr,�H�M��;EQ�RT��W���J�	Ke$5-*ǸI''�$͂�S=0q���粬�ѭ¶���v��F6^ꬽ��~@1���U����zK�{`���T(�H����6BÇ�s$^���ڧRc�I­YXk����x�X�c�D:�\��������0�S ɡ�|�����٪0zu�n*��0��U'�����[�h�d���X��:#vA���P���suc�	�AC��g1uVI��Q�F�����'�@ �lq��GZM�����k(�M��Y���\|���ʑh�ȯ"�:,�kY��?�f̙��.���w�߅��]6�wڪ�+ˡ0-��-��,g+�]bg���EJCSn8c���7&bMI� �UB�������I�xA�a��˳z������-jW,�cÓ�D�I��`{�J���j�Y���eUC�߱�����v�c*�q�DH�q�5��5�Ӎ��_W�?��8?�h���< ƆuX�+ce^m�-���yc0� z��y8��f=+E3������ º�D�Q�G�� �#+�)��E�ր!W�a�H���"�J�q(�W�� '�cِ��әD��帣g�w�!ui����o?��L���Z���ђQ �<a�Q���i�qG)��)���j��lF�	0���hY%_���CO�����1y2�׊=l[���i���9T)M�BMX��xb�������@������۴<G|��fô����:oE��<(�S\��93rl��	��̇��S��3�'bI���כ��ߟ-���&c��P�SX7����E����9k�7�����t�B!�
���f=��4W�Y��(����4�M��?�>�"�7=���	i�,@�Rp�eiRu�V)MQ��hX��:����3���	�@JC�(��q�J�<a�]t�<�^��D��%P�g��9,1��]���)��úN.��?����4�ko�ѭJ,""q"`2�n�X�C/���d�$�*����a�}U��̸�ѫYM���m�$h�F:d##6`;���%ejuf� _��������^�\!y�����l���Y���\|�$�N��bM���#���B�����;�AV�6`p�:j�Ǹ���1+v����^��m˨;��>m!7fg2J����}�t�i��{��@�3E��\Es��O���f�oɝ�yH{�+��z�hEb�0��M2I�pc[)�K��D�v�İ0x���d�����+��u����1�t<ڟ������A�0�Kq����	5_����,-�H�֕��yA�c%_8*.+�Z�0��|=c�Xx��\�nV)�n-kZ�b�d4�+���\�{�DWaݦL��7�B�宠m����{�����(X��ה6�k6;w�~���ϳ���ͧ����~OB��@�C�����|� M�!��)�50 '��/����F\�0ju����P��c�O���~���_�cB�sRC��?��5:��z3S-?�C���D*ԟ4�e���~=�ݞ���� >YH��|�@~}�~�z��a0c(.M"U� �lT�/���?$��z��@bȭ1"5��h��,E��t"u%�(ɶMb��j�
`e�V���;�����U�E����ՂY�G$��#p�Mz1��_o��KB5���+��^&��^x���7L��$p@��aٙG윀|{���f
�q��X�z��>�t�D�t��؈b�=��Z��m�bF��WJ߁WY^u�+���΄7dZ�1��؏���A��1��P`�$�W�0t,(��6�t_�VK��Rx�#�L����&CBvv�b�qB�d��˒EfA���n��r�S��M��ٶE#4�E]yUW�:�T(%<���L1*j���h�����F$s�m���������7�L�1��Gy������y�4�a�X�[�&���
���`l�Uɨ=�\K�	��ua�9��qĘ��"��Oճލ�+dMq*Y�Ό�0�d�ϖ������>�g�U�w:ڻ���1�L�j���[V�M�蓵��pTǳͶ��`��r�m��j-ƛЌ˳��G3kb���Ӆ�u�S�D�"���%�!��ۜ�qR�b�uxȕ���L����]A�+:�� O����v�
�(Gm	%4,��2�UVPX�˷rS�W̒Ԓ\F��w���� ��]�{�l�10	Q�� �K�}?��[�95�꫾����B����͕������r��	LNU��!��\���\��D��`C}�h����3�de�����ۘ�:�}Q�7}�\]$MxO~��I7išB�r���3n�h�M�y�"��zq�:KL��uz�[�Ƨv�;�iY�����12ѣ�ls���Ԏ����ݚ�0�	!�,r�vQ��[�e,#j��OL��l�S�x�T���Tt&�+2��~"����@^T�Yݴ[�pkB���Ҝ�"�ʾ19/j`2������Bz��
Q =�SP]��k��'ׯR蠹�\�X�A2ϴ���8��`�͙�8[ؓ���.�?�Wo~�"^_`<H׽5���R9���jN$���/�X�')��VN�њ
�r����ŉ2����&��n�K�Ю�~g�DP-&%S��9����EJ\�]#BPz5VC�m����^�X��5Oڴ�݈��虎;d����j4��|l��"��u�������j�P����P*��� z�_���M�h��ǋ�����	c۟囹W*��fZR~\��(�9�Z<�*g23�s�DiF�[n�Zv��������˿�)�V��@1P�Ī?A&�lYY�^pf�9ی��rb�AI^���&~"^jV��h*Z��8�t�*�7'��2�e�m�J�T!��n��U�g
���-{압�Y�lF�~4����X7�H<n�'0�Wp����O�	��=��̳*	M��9�y���U����V��S����|�))ե�iKDˣKk�4�0��3_�(�i�0�_v��i�@�4���
��81�ha[J�� ����M�Ǽϐ�L�]�{���n�fW���g9�g_H�*�D�<b�En0��	�Т���c��:?���cØΘ���9̀M�ީ�Uv�t	�w���3�>�|�Tb\�-�5 {��q�bIeWcV �zq�n�$A���5p�NG��=�Z�1a������o�P_���J �����1���'xxB3���,*�ˑt|xo����~�Y}VrA�Nu�j/���+BۡR���z@T�QM�eKX_W�w@��&�w�b�*%]�E�g���	��YվѹefQ�q�g
�BD�������\u�1�[e&uA�Z.��!�1��B\��[�ׁ2+[���B�ÁH9��w���`���m��~
!��PG�� J����lGN;� �T�`7[���2�p.��"f�2j�[�L��!$��](�9w�!�a�e��ic�ש���F�����B�?��7�Ix�N��+�4L�3���!�S?��s��������9��&��`�0�����EA#�XUs�&�Gx�+=�[Ӝ�A�g�wT�[GO8�Vz��m۴o|�B͹VH��f2(�������G�Y�tG%�r��=2_�g�O^�-ݟ�\ҭB� ���q7�.�T3�Է�8��mV�2#,Bhj�k;k�� �T$ o��h��#���6QZ`<��])�k����SO�oł�~�����_��:zǜR�.���ֵ��D��d��%ǾZ�<~�܈�$j��'q�yl�U�Y�g��\��zi�����	�~�oa�SY�p���dq�]�N���\Kt�m�
b��s�{�ʀ�z�ÃU]=��l�w��<������_d2rt���U�lڙ��g�(��a�5k��٪4�(�l'C��Qe����l�Q�>�\��߈w��#�y�-"�\��s)�ල�WB��SY�����[%�
:��l���R+�(��AriRdKeO] ����"�A��@���ńN`0gIhG�1�|�k��[�2�\G���{�.�~8nnrJE\Qe��1o	[Ai{�{ʠhQc���NJ�v臼�����5��X������\;�����zߎ�K�n=l*�.�F�J�����X-���c=A�Έ>�������Й%.���a����"����Ck*�4�qP%��wX�n���c0t{�w�Ȱ���*�����o�b#s����P�^�v������;�'^O.�,eF���r