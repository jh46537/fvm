// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:30 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dJFT6MIA815wQXU+iopM/GUsNfuTYqIFSO7FjpSgICxQafuFZavEKB/FcVhCfxi9
Db6aaa+rAF63zBshRt/l6/FqJl77EGYYSHRAlJrZJnEx1w0BYJKZLvYRQQ+l1NPs
OzxU9Kdqsg2Ft8nkEAUYyXdyYw80rxc1AwZBqYOTpYA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2896)
pEEM7Oig8+w1Gb25EkMHYVMBya9yfpJhL8uIXN/vTUIDfF5zjElZA3WoXpr5JDIa
AjyLvM4YH/rXfM7EIvDQMXUAB8XXWiaAkIpNLheY1FbcyzcgBQ9eX1/cj4CECCNm
Bo/oJoOqi0WdLbzXR8amJf1S2keFcWAY9yEUIMbcVptANfPTPSA0766HvAFZ+6SD
7WDn89r6tB1f6AJOis1yT8OIIJWgUTMhips1UJ7ijhlZy2D++D/XbQUnqg3lV8+g
AtyIFnqHBsBMFeAznw6tD8FH+So6Y3mNX5GLLyc306lz6pCGUJO9om1vzwZarSVZ
aOPaLNZR7RoQW9ioZqR0mtLt+O12F12aKPSNoZ3U/w+0/fGsYA1RTF76lMYODs8w
ozoFnDRyyPMCqgAtlkg3iRY1cSKOfeSx++0Le3UeMZEOUu+EO8fxcssGwPq1sQ5/
Uwrb9e8HXJGg3oLRjzC6w4j6xq1vPnCWTAjZrc8xjP2wcHXjKNSo49j8XoJoozXs
0mNPumgD+anKUD6qbc9PjOi+KCku6OJm97NqdDJs8tp5tqhfshURGEpC56KvqG5S
5maE7Cnkzv/m8sBOs0K4BYZwGneq7VsjyZAi7jw5bUWVPn0+msSdG5S1vJzKccms
V9lpkO+nKAdej7tzKKqqLZarSp6jTZfelKZUAgCFthbCRkWGmJD7C+hZvT5d7lJV
Gp09Xe1+lEd/70g59MQ2V/vjj3IQJG1qk04R5xdqUMugAnspZhsyleJerIRy2vGo
I/VNRbcpF4Kw2eO2+Wjx8g2+g3DJ4jTTF/kw7ycL/0blJGf1/Bn7M1+whdBSNjio
MfFxE0p76fcVKVMJsMYbk0pmH/X4uRbR3x+ly1enGYPZ0C+ZRuf3re+hZotyeNUH
9HWIKQfVpS7IFSnv09E7krp0d83Ep1lcQxC5TpjENbQgtDcTaQ0Ra/wFkITPLt/8
GdNrrnOl8OKJwDyJUnVVdVq6Mg0eY5GPb1bWubOeEeqtb501jjeVa/hJV3F+RaFU
Itmh2xes8GNaQbzrWCSRKtrvNqF0ruaHmko01Clyu5dpLcQtBKcFotVjqD/Xz85i
jCKaes3uiDHgFwturhuDgQJ9XyIBa7zoAVTrxIaUv8GuIu+XM3FrINyt8GDfU0y2
N9UvusGpzahcq6oJZo3WBtbW69c8wyVDX5Jvo/p0nGmNhrT5M3F98eEmX3YEIlPu
aCUh8NDkPbC+tvyGLkpaLLZiHAaYQ9lz5W2ryVzvRVoOZxqa/oKyUpQeFUpLJsQv
oicU1MmeTTwLaU2nVS7aUfh6X9edgLZ2G01C+BfemmcTJ71zPudbQRtapsQGMQcX
LL6/bvHI8FlLwPIj07EWiYsrNz1GHpck8SMPvmywSaWOm2LxH8kOMeN+zWzphnkK
mgQVTWUfC8FHKCaKJnGjsP5sFudbLIkhgTM4GtaZfcBbgZzGztbHApXVPjGgMC4S
usOBlfg8CilAAxTuVR/OEKlAphwNu9tXOlCpptzUN5h50D5+LqwqJN91FkntT5m0
FofGiZMSpCCvy8jv4uBKaek1GxG6s6oiAZfKrqPUNWRHlQ/KZ3FqrcsrFFeP3UOo
jOq/qVuXAGvrNHgpMOkE+pSJi3BUNBamkgQcIjyZ5ijk0FZWbRvKhpsE+/Eehxf5
J+6qFnnry+Q3+ydkRcDcT0EyPlzdDqDFgvw45wiJFaWhhfS+weCJqtc+AE/bgYAi
MpoSd2mEHB5EjR1H7uq014rwo0XhtSdz4+53Hbih4v7zT+Na7j+60Su2dP5sUwBh
d2CSRM1By6qZO/+/rYU4FXzXeA/NbwHTMjkh+b3m6vnYoC3eCJKd5VqsPZ/EDfrt
chpj1uayla6xKZ/iB+dXKq4fWoFlRSaij4/UO/mn6mlJA8+ISXdfn4Qo85PZZurW
DDfCEBN9hNzrcZNnR+KZcmtNhi/j/EtDGb6r0CzZxIU76jmvBwUB5KZhe1Zwsy1F
WkVaUatIA9+2TmnCxuTEPTFio6/0cVg1GeiCneAVIQDdO2Wt4m+Av4jV1IgLpoEN
JHu738ePVmqAfohISC20qUwNcYFvGzzyyDqzP/MeRtt8wK56FWTr6yAWF+CXdWAS
7C+Z6KMVGa5TnXURF1T7YGTr3hCMAXrysG5whNGII1ELl70fUcsfBaN/iE014Cw/
7aWFhd4oYoPULepQlDcxcad2Xi8SysGSWWfS1pICj6yD7YAkc5e3B6ltM716Rcw6
JK6P71ktkFqQnYuyq5Y1cgs0dfAGSGl+cJDzBlL8fSP7L8VneG0T09CWfRrMnU5x
hjlls0d2e4xgaO2vpV+sTdSFZXrAFgXTnv1Ja21xlDxLJ1Za9w1oJiQSIGRKDsT8
SD8I/ya++iL2xxYhRS8lsCOb1qsG/SNopO5vc+r2WykyuKDTExakWxquJP6amsEC
J9vkZTFleQNgloGC3qofmSkkHS8KPCVZWFr2LicIcDPVHwks335o8AkXDd5bMvX2
prbUTbjuyQoK+f8kBG/ehncJ6tndo/PooTxI7V8P3qmGvPhvJ4uAhz91X5i3LITx
j+ppPRQ4RpoZrqUzCnRMbgrRRY9xcAQFwcrESuvZDjmxAdx+7k+Ztw21jVzns9wu
d5FRgoMqfn1a5uEgNi3iNgVyBk93HJ6z5yxZW3I3hZ74yPbD/SSR3RFKHH2WpxZw
NSNXh0Cv5UJkxk+hMzAz8Lmc8xD7NhAqW2HE9YIe/VyZBE1F1BQjJQJIPBEszENd
GTRhizzqXmh6o1RCcqpr9/m4Da8ZbfkCIcbtcNIO7nnJQNKUSGRZM8e4qOXd595t
JhY8HrzgguOtU6i1/k1Y+wNG3Tg10KBoN0KmxW3lrSy097M38Du8yWYnZVBNYexg
Hf/ABzgCE9O6/jzVhE0x/4I8LtJf+d/xz9iSSOrDds6JzNklGdW+RinMY+uVOeSS
2/0yWYz+DmgHQsROYQKfCdig5kIBgypquzUMld1XOkIvouvhtkPjA5b32YqlDyfC
NVNvKWDgv+OSbkUQ+U50IRdJGyxec69rZh/nyG6+e96rI+335tJ0y12Os8iD9lNy
SgrjmSLNjI4WEBYmNlTNEnDe43LlzVFLeFLFLhAJYiN+rmYeCvWtAQBoaoluArZV
ea3jaicbCL/Hc6OKNDW5ZtuTSEHkMJg6bghi8uUAimYeY40RRkD9x+RTjsYxKmJh
j6lFmHFZKdgy354DqAeb1EO+5I8AtHJBodO3lmwIv4gWGS/MEnYo4h6nZHvyjFUX
2IsGAfBA9MQSxBUjZzqBvvxKYXIPo+Bj1PrtN4TnTkSCZ2AbPn84vpuUSnjueQ2p
YXZZim7vq1E2njy86G/ATU8eK8rAngsqCZ01miF5cLXLhHeCC3M4rbrNDTmgW5J0
He30fji0c1ax7Y6ZIZMl/OvvMOHKuI27nTumnhfmM0bPInBXFbO6tCUNE2rHsiAx
QPRt/QOQO61KP74GgMMiwSArkMfGnDTGeFv5OXZG03kjfM/ku5/OaEUfD9+1GDGI
q5gNgL7Qz5DtcF9eJpuXncbkNSBBaSRjMnGDatOrz19vL4zEtgXM7+a3pFOlzBTj
nGzu5K5rkl/FxYV4IbYmZJjfDFJLjjbc4YEA4JEnKwm/Mp3zWlCAUYf0fKmjrtcL
rqS4rSXrnAGUgkxIcFx/XOtxCBLmo+WSVmVF1nU30NtVN/MuTzQD4M7Ypp63faPd
tFVpYdsQif5pYEB99RinCEwi1Rj3MnE2ElJpEx07uJE0zkY4auLvACbk9Ddp8KBe
8FaznlLvYZ7xJvoeYdOPxIPEGaqNFWNNfHOdOdxIrfSnjrNbxdvb26ksV1UP4/tF
1iONCzHXQmSik+67aWgiQA==
`pragma protect end_protected
