��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{�ףe��	�A`������I���6��K?Nl4	�#EBQ9bq҉:���~R�\y�o��=@O/,73���`�f|�F$��wu	C�`�03�5���ʇ�R�C=H駊#�j������!Λ�F���� ��6�#�'|b8N�)\ܒ#Q����4o3F���m)1���Z���_� R)B˕�ʵUa�3�Ek���:�V⺩�Yߨf�85�R�1B���F��ߠ	�=��!{�~
��<�ͪ]sR�A�u��[�/*hU���c:��@��<����Ĝ���A)�ւ��cG��ĜQ��2t ��
gÝ��	G<'_t6�	d�!Mk�7Tb�W�d��d+�BL~����̹����=d��,Ik�m���ߑ��rO�2���~��;�WC��/QDEZ-xt�u@��~�L���:�3,E�t���'����3��.�X|����ΰ�j�,[�~������|Oɿ�z�.9#\�s�K�l�i����o�����b�?o91CF���Lǟ�z�.�i1�I����ǐ�.u��[
iOA�x�,4���1o{���y�Nu�/?lF������9�f�j�?��	���H	�C���!�ځA�Bb}�a�UL��Jb����R��������Y���\��rt��IJV8�0g����A!沇��=� Z	x�S&-Ѭ��/�*�c�+|�2�dNX�T����k�mAl�s��M�$i6����\5�}���F�6dI8^d�Z��Z3	����嬅P�vmz�M�����"g�`s<�6d
V=-K$�_)�#ʾ°N����V��MKoD�;}E���3�A���'��?zLz�E\{<���u�����rn����u��NH�9nFԌ�˷�sɴ��8�s�T��"ؽ_}��m�S9;.������,U��UjKP=�]��T��SU�ݮG:��7Ϯ~	��I�I��"�P��S���Ҩ8\�9������4c���h��l*�R[C�7��DB>dT6�ƕ����$4D_�/y*T�Q�˘��#mF��V1֋)d�ȥ~'�**�D�.	�z�͆~
	x�즒�g{��E)3()�А5C�aM��ÚoW�D��WG�0�8M����"�,ţ,��=k���ÎWD�ﲳv�5��hE������й���3û�	yP�[X���bkοg�ƛof��o�C�I�y�;e�iA��'���ŵ�(��H2^����-;�Bj�B����ʟ��-�-q��� ��M�Y7Q��|Dҗ��6y�D��ww�����u�� ���P�B�-g�r
E�lH��=� 	���g�� �_�Ceq�a��"�[�P�,��
�Ặ�4м�:�W�HH�D��u�Y�M�N�U���2�p ��l��L��N̅(��Ӷ=��v�!��V�`���pz�q\-���V�ðJ��ޤ~7]F(}{dE��0��m�r���Ҍ� �.��eG�`��(kf�SE�l�Iǃ�k�ϥn�t��8E�k4-G{�X����[���3"ѐj�`���*d+�l.��I��M���76�/�BxBc@�D�K�l��������eT����{�����	Z�sڷ����&��[�p�@Rk�p����UJ��&�-�JXj�Am��`�{WN�N�2�Bة���|�{��?;�U*��]ɞ
K��v���V'z	'U��>bw;5.�(�����YzEH	X�-\F��rD�A)�L'ؚ�
�?�&g�2����KL�HL� �j�g�$E����;�i���N��
��63~�Qō��<�L8;��ϫNSA���'"TC��+����K?��L�ـW	Q�{	�v���U�O���߆�#�:x2X���h�����4�~�HN)����U�$>��q+�񅨚��&}λѐ�M�ϗV%��ɽ�N�=�e��
�<��iǃ� ^X�Aۨ~4N�܆Ao�r��两|�L���d�����Cɵ%6�K�٧d�����1�B� ���D�.�!��N�l$���,�^�E�(Mm�J�	��'-��X���9��a�+�|�i���>H�{�"����wC)��ߚS�h��)�Ɲo�zY�o��d�v��[�:��	e�K
4LGi9F�rs�A�3�<c�qxA�sZ[D��	_�: -%n&z}��ՠ{�4�l1�=$�Md�e�PP����v@������b�PH1�a��uߓ�{-t���?�U^`:��y�� �����;���z�)��&���^������sw�-t�3�m0��<�GsV��E���0}��)���	�eU(�7�ހ�#�]��i/���X�G�֕�;1�Uls�'L=I��7�ӛ���c��Fd3���&�It0��5�/�ϒz��F%�a2�yZ����A�PL��Z�K<������e�ʼ�e���WuO���	�ީ)��*.��̵TÉ\4��r޺�E�?�ɄWT�����k��+:r�C�� _��z��M�ݱ���r��'a%3�OA�'�"+y?�ÉZ*6�+��:��mp'uGtK�*�9��\��2E�sR�ORz݇,S����p����;�-��:��s��_`���S�>{i4mq#�n/_��*���`�d������qy.���M�D��$�f_�d<��<�k����C���x��jqI�C�N�\A��_�s���fC�����Qv3೛�W2��94}��l�i�U�8sg��y��ew�6L��s��G�߇5��+��������T���̙��f��)*�B ���	zm�S+`]�["[	2m���I>6�G��3ʼ�-��`��8%����k��ÓwT�	k�پ�79���U���o̴N��%�j��H�"	JR۽�|d�{T;^�`U�Z0Rg���x`�l����߉S�$+K��=g7*�J�[�Nn�$^E��y�\��U�ч�����,*߳[�g �?O�s��_����up�?�� k�٘�����P[ե�V���j�-��o��#��B�(f$x���GiE2aS�(M�� �n �R�@��?@7[�uۼȆ��5�q��ob���������l��2�<��el��v��`�_�N�wb�eD̲�X=�ސ4\O���x4�h� ���;��W���ϛ�p�A `Q~+>�1{ϕ�s`#	���=��he}'�$��f���~���C�nK|#�Z� {^�~��}�~��F{H��>��UP����lq�}��6�<�0L�N��=J������9V�Jl�m26B���C$�0S��c� ���Ǔ�ƁI���E`�	�:>��umǶ�@D*�u&����R�&%�k<�����zH����[m����M,����&B�r