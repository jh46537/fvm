��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>��������ّ$�*X`F~�������><06�L���\�D>�WҎ�����r�.~O�I�V�X;w�G��ts��K�5���t�7��R��пr�.r���x{��}sbeq�XG|7 ��$�ڳ&�e
�=r�$��!錋"���ۆ[�8����lr���8Yi��9���eIE�(Z�)��VJ�j��?~�	��c��R�6���/�WC*��B�����-~��R���$=��&����O6�F�~gh��\P:�w�o"Z��{��ܪ-|$�EA���ٔ:�_JFJJ��S�B	*.�a�ꇔ�@�/~�WC(���&q����?��V~��A������(}�b	ѝu�%k!gŝ>�I8�s)�u{��>kp�Syʰ+�� 2����=��D~0.i4��SJ~��U�h��ERc;��@�p&)Aǳ)��� hU�`��ߨ��a�u~�\��@��	�L�L��*3?��l�'�&��rgRUu��������'��E��	�o� �í�<�t�����"	��bnz�nS��H�v#\��f.6��y��/6�ٍ��]��0���I�`�>�7��X,Tq����{"}��W�`Sۛ&����8������Vѐ��CO��T�-`����~òn�����s��	[eO�`�2�����ۧZ����wD��_��kY5��?���qZÚ�k6�B>�����U�Qg-#�0J`jxx�:���oj�y�����3�8[K�![��7'�^��fMm���	ac���
�wES�q���� ��$�;�
Dk���y��;�ת�l�>c顫GR3�J6^�.U�����.�&���g�~,{,����@�n8d�f���55@Z��%� ��4/D�w{���@-ľF�0p0"���Q|�=�F�"Ɖ ��U
�~~�[�0&�8��1]�p8�2��t�Y�
�3t�D+[�/����VT@�����g!*ue�t���ۛ�B�pƊ�7�J�7�E�.\��7��%Ft�]Fu��gt�	�����7t���ՠ�V.nM���H� � �3m:Ey˲w@��Ƅ}L\��}]bo�~����e��,[=��B�F4x9P 9!G{�:5�쬚ӊ3 2��pC ��I�t@_(H@��ǈ#2j�L��F��v������$����G�,]'η���)����;�X/5����+��>c������`��2����3=Ql�5����8..34�q���U:���YWčK�uPP���2�x%�����Y$8�?Βyi{�&� :D?f�Z]g#F��#X�s�I��m�cm[g�M�����W|�����հ���6�ۘ��Tw8�Zh��1J%xf'�}��a�U���Jrl�F_~^�,��̜�MZ�ʍ*�� H�~�~
���lgc�_y�m�K@����n�$�839��*�>�i�~i�		��Q���� Fs��`�6��J*�`���Ɋ��l��Q��U�þFj�{_5
������u ��p~�M��s��Jm��e�?�e%6�4#v�1?�{g}૭ڙ_*��j/eL�>��%L|�ιF�J��[Q_��#��[��έ�`\�^�@�w���?�"�D�@К�m^�(u��o��
��y�.��x�Uuw1v�U��>|HM�>*d���ڽ/P��ls�q��?^mR�SX�!~���
'?����K��(�o�M�M|�M���KQ�h�~9,/-�̔J(E�jM��u�[��r#�(��b��׫V2w���Ukc��Y���.�>ql$4W�m尪gl+��h:�N^).c�}k����o����=����5"$է��Aȅ�� ;doZ��+�/4	�i,�:/C �\x��f�u���)@.�cL-��Lu41�1_�j�z�h��+�\^^��~/��c�a�tP��?ʝ���D��A�w
SQU"�U[(���Ҵ&	^e(��@@O���_k�g�"g��K-?s<@"D�7����s��p��P�]�{�W��z��K?M��g�c���;_����Hc4�׼���&ܞ~�J'aM|NW. �q1޹��S���ꒈ�]��w�l�5��.8;H6#�N�P��d3`�ήY�D����0��w6|����{*�����&��F^ZF�����Ҿ׬]B|�TNa���iv��RuP�l{嘒-��0�sB�s���h����&a������&����Rm���aEZKݒ0@m��th���3�#l�Ţg�p�˖��;��l�<j	��Ti4y�zwĆD@k�c���!�ԓߢ�)�����aT�|�����ʬ��Y�T�?�^h��h
��dCO��I�+$
�٢�5�N����g���qhq"�f������{��o�0�ʦ��P�p�����Z�2K��;�����K���&���Uh���hn`/+�2d�P!�}=��Y��6j\�932��YI�F� �8�D���i�ʦ8V���.
?o�J�t;�ʷ��!}���1���3rN��T�ER��������wsq�ud�;x������H�cz��*M��/ӥX�YX�k'��1�k;�^h[H����@��U���ԛ�+���_�4���2v �m�i�j@� c\���ki���QS���Y�i��h4-Ѹ��90�|�
��TC�ij��Rf�;�h}8%'��z��|���OL�}d�v+� -\��d��~S�ɏs�k�yw�x��f n�R{��PP�)@�[<�a(q�llw[g�#��~��E"5C�ըO< �S�f�HЬj���R�@�@OE���=F��x Q�0]
�`��-�Mh<�Kf���B�۩���݁�*�}�r�D7���v��"8[1��a��"%dh]�cP�>[�{e���xf/��������^1A�H�[�k���Lx����G��l��;85�ǈb�EZ�.����|mvL��Pp؎�����k=��_�nA��Wla�h��L�Gn��qc�/���`����n]�Caq�%����<7�"�~|%t6�o�i��j�i�V�Ӑ��N:7�.N 'P�8�Ws�dҠ����R J�+��k�,�Ue�F����9����	)�H��$�/�-�w����PmI�<���ԟ���?�5��f)GL��دk� �#�ob3]���I�yxL���e�5��.�28��~�ԍ�rS��EU�tG���O��Vœ��g�� �j���-=��|&����Vm�-L,!@z�4���JѼe�b/Q<�vF���g���ݢ�"��' �^��C�WY�^g�\�eT��勣7��b��1`-&y�!��z`��/�a������
����j�A[GG���Ѽ7�3?�cm��y6���b�@}�^b��f!*o�z9�M^�k�(t��f��&�\_�;
�Lө�q���t<�F�Y�2��й,���Ϣ��[��������%M~����D�O��JM��h�L�y���ϢJ����"�"��^�E�K�lꖇQQ�$�@�=k&�(��4�	�Ent��(�D��_|���(b�+¾+}�O-��D~��iN��d��V�/Ɗ�Abw���ʉF�H�%c���F8s;���Gs{�`=��3�]��ZU% d�E�U�~��Vpܓ���
����[�IO��,�.i�I�&r$�S�H�~F��Uhe�!�@r����6IZ�ʌ����A�����v~���ҿ�����u��vDy���&�t܄�ĩ$z{k��e��%V\���3�M�|�1������6;ɿ�I	���˹��;��5>��,�PdFE����Y]�l�R�|��	 S��G>�e�����h��n
�3�.��[1?q+4����N{�� L.m�@�9�Q]!t�k"0a�:���w�]XǄ�~qm��D�̪6�E�B]V�wI���ړ.��>�(�@+᥂D>�b�����#�70Z.	&1� �����Gy�n�Y��c�A�E��]E⸫X�ƽ�ْ� �Ķ'd���=^I�(���9��	�_z;\_M�ں���a-����U�nl6X҃�Q)jU�0tcd�\������j�T��˭����k� �z��s�WЏ�b�	�>��������Ֆ���Ѧ�߶��!%�y��M�t�'7~��kW����s�"�Xd5#�*Cgg�M�@#u�}�9@$���$�G��;�?e�K�K(��S��o��m��8_���]�A��=��	:�JY����o��z���wZ�d4zٵ57���:��3<Vej����Ʌ���X��S�����+��ZL8;Տ�"���%����J
S��,_U�K&���@S.����w@3F>�̚���a2�-�����Ϳ��P<�޺�el����<����!Z9��<�/~�`~<���w���RJ*]�~2�nc)�o^����t*l�H8��u���� �Js0���#Ѿ�cǪ�Z�1�Qכ��q�(L��E�e�׷���fT��m��Xm+�xW�qy���� s�^<�6ҁ��l�ː�]�1&��$e�KeGƻ&�U_��.M�Ta�0D�8�& M��_�3��M1�y7��;���W_�A�ے�R���,���nn�	S(�'�=#bh"p�q�L����l`�����l{U��^�nIhTWǡ[�\�Mo��<�V�yϏ�>{���P�������	�"���s�L�b�@h�!}�SŐ[K����
Ow_"z�)�[Tg�<GKW�U�q��U(�0��״������~��&�Mᜣp�2��*w'^�K��rK��킛0�7\V����d	��Թ�P� �q��<��%��DB�)�L����
�p��k{C'�c�)d��w&$p����e&$�Suf���8�[l%��/M�Xkw'"�'e�H�%Fa�O�_�91S�qd���P�A��1����ya��^��b��G�p:ʦ�a$ ���_��>m�����b�[2���ߧ@��F���Δ�1�g��Iq�����*���5>@1I�R-7?���"E�Kk��o4C�B��.���A������mG�n=!�"H��;���ޮ�,l�z�.3s�"�+ˎ�nJ~X�X���'��sٿ����b�n�ԋ���[�l��g���F��T)4�3�%t��� P�"��