��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"��m�?l�3����9L��z�#q��
&Q�����c_�����.���@��贂`�P����-q}���z�{�����q&� ���|�!'f�<��h��$X�U�U���a�AI�h!w#�FÎw���D˅OIIT����Q`'�}��;����(A˒?I"r|j$��f����#��~�FX��%��7|�w��r�!s��	2����Xm������u����^�	��+:ab���Tjn���eu����, ��������z����gn�j/�%Ge���m�h ��JV��W�	E���ր��덒'��(�O�C֝�-����K_�8�8*`�!��=F��A�i`;{{�ᛅ�j:E/L^���x����̇���(�њ���,�����evf�:��̥&q�Oc�G*{tV� ͍W���W��Ҳ�fX�%�ex�$���˅|J�¶��*�1��9��\ɍ'웏�q{ēؾ7���q����� U��g��@�fX�q��Z3���0z��zQ��O�VLP��i�C�Psd���Ou��Q������~����`�$&��i���F)�6+I�H6�:��u�r����E��/�C�Y��L��kT�΄_����h�z��_��+!�6
����k�ڠķt��/�s ���t���������M/�$b�;�#��!�7 m�hPH˘=���:Wi�w�$�Ro-Uа�׾ߔ�e�T*?`p�c-��r�{���ǜR�	�I�!�ܧ6 	V���6r�4�K��AF��2r����-%�<�ݴ�М��kW���3�a�W\�C\Iŝ��S{ۻ�؋�6�%n؟�����\F�z��Z�gD#!���}�ǉ��-���t�ܧ�=04��&�������mLc<i�i6OK(�Y�,�$�2��fD�����8�#Xs��m�\�AЩn��>�U�}CY�,��1S�#e.A�=x���-���^�����sb._�"��4g����JG�u/�OWJ���X1hCn�O5�\c�(j�|����[�WIo��[��T��j���q�������͹:�f��L��#�+}�L��k����>�R4�pM�!?d䌎?WG�HO�J����T��'�(tX�&Ӥ��:��/���_���:��A��/�j�!ðA4$j7�j�����CAR�:0�,��q�����)��o�q?4'6��'T �R�C��T��J����4�w�rD��
�Q���{dSj��|�W��s�ȹs����Y�.�'���05�� _�ub	�f<��*Wjӿ�vݭdg4�g���d��	V���ŝ2�b{$c<��w��X\�Kا�=�����M�`7��{RAQ�38��c�,�Q%A�J�����W����H�nc��0:��� {7�ܪ2��Т8����wVA������K9h���41z�X2��f ŧ	П0��_T&�����؏��GcLG�]�p���)V���O���#�d%$�if���ކ�Z*F�W���6j��8K0�N��`L��2�b�3O�}����ŭ�=��y[���o�b�%��*�Ek
e���<V�).��b5@w/<ᴭ�[��FF�f$M8R|�s�.G��ࢄb-ej&�k8�V��U�@���T��D�ý-��ܔ��6��!s�_.���z���:9n�s��:�e%Z��`�����C;�� zj-B�	~��Q��C��_�ƪ�|���P�(���[qX|2�?����)�>x������ϰR���~?�Gr	��`3D(��P�(��V���uc\3ϝ���8�bXu��љe�@��nym�F}�B,w�E��;Js���`�Y	�j�D)��٠Or�3]�DL8ٟ�1��`�	^o�C����/�U`��3!�UQ5L��19gsm=&r��d�2t�ŞB��H�.��Z�g!�Q����� O���<�7���
�04�1�+�\�Ajg� ���Ĵ-��g1�o��2�7��8��ev����/�ub�����ka.�՞�B�����]Q �4>��	R���ԊV��6䐌��*��	e��g���Z-�d� ����D�_`� c��g�c�)	���vF��~���!8U�4[�R����I����4!i+c��`�`sa��V���d������x�����*r��9�4R��at��hH��y=���1e]�C�/bfg�ys'�'p�e2 C���<�I��}���*�>Vם�o����ч	]L'"P�z��p��$����f�7�yϫG4"J\�a�'J� ZN7SK����6qo\?��(�3�ɵ��8&I�m��~4�"�	��Z᪢�b��8�E�9�J��n8�Kȷ�}Q�a@]�<�X�{Z����+�8��+�#R�#��m)�
ɱ}���ǰs���a��������k�wG�2�`��bT��Y�Q��0M.f	�EW���n����*hU�,m\��$�+&�b����x�9�7E��T���ƥ���#Ȏ���A[�B+�ya\u��	�P�N��C�V�$(ڄ(B������c1����OO�gF O7�,ق��x���,�}k.r���ڃ��Q�D���2D�Kp=e�9ҖD�X���"思�7�H�(�2�n�Db�Bl�[������6蝼T*B�)u[���� �m�P��6�ښCͶ<P�@h?'�)Gt��dc?y3*v���=b�� -|m�~8�8�^V���Q���[�fYb����E��x(�]���zs�2����:Kd��צ	|ī��"�-�4��p���}���揭�ʻ�����S�(��L����)]Cp�W�lK+����%(��f[r�~�Ч(�ش�wᮥ�?q��~�|��������"@�C������Ύ`�#9���CG�U���oD������%�w�8<4ĿH޶U�=�$лz�)�ŭ�6dh�Glg��K�uD�҇��t��p��F*Ȍ��S�(
ǆ��7y>��%���1KSL\P�_����a�!�w���$�%�k�>�?�[;4�@�X��m=,�n$��G2jU	�Tҹ]qM����O����ov�K�Bcif'�PL���W�Δ��$���ؽ�^���f��랫8��+�붰���G�&hȥ�%�AFOE�v٬��u��'����0N'.�¢���4�;�%TDEG�'��Q!�X������º�����<�N���.�Y��K��ũy�|mQ�$$V��Մ4A5����tK�����Ԕ2�T����I<J��G��<Ǥ�!P�?֍C�
r�Hx:^��Tk4�7�_j����W��,o�ؾ�Y~��r�O�������$;�S��F�[q)o�)�S��)�NW���)?:�r�f�)��������
fU�L
�u�KK\7�(�
����_x@9�B���A��8�ckqk��v�ƽ���}�M���<������R�OB=u�p�G�Ǵ~"���DNO.=������m8�BY��tօ;�Uc`edj�/�-��U�g���]��V�zBiy8-Ő$��u̲�Ac��i�û��p��W�'���q�� *�,U3�S��H�ya|��Z�#&F�S�a�Z���UC���9� ��b�"�����.Y�~�`d����aJ&;���K�9�1`(am��a���d��.��˱���3'2����)*P��_L<�˳�$���;����Ҋ�IÅ��#L�����=2t�feTO8Q��H��d���������_���?����!^��S�Zvs���0l��?Z��uG�-)ji���K��,�ݐ�RU�/I��F�|��J�3�jK�2�&%S��8��r��J����o�ᖰN��pE�"�6�69����Ϲ��ݰ�/�)09�=��hMk�RZ�<8���:�W�L��C+:Sօ��(�Jt{̥L�d��8:/�}�4���3)C��B&8g���l���\|�����;�_�5֋G,�����[�jXA�۸�5�c�ڳ����Q9�}��ւJu>����H�]F���C�(QY$�u����Q�e8��y����f|��v���1B��d���}���c�#3��@�}r�P,��D�k:s����_\q��)��0��ʛd�ҫ�&iPYn��k۴����Q�d�R�ñ#%s�K�8ɮ�V�">�b��+y����=���s#ԏie��hZ�6L�L&
�+�w��M�y#i/�:ߝ㗅S�e�V������m����F@ T��@�=�S��g�ͪy�>��U����Wr��b�� ��u*����`U��w9@RY��0Kf�vԫSN���U��X���v�4
%�(�W�n����)���c�D�{3����^He�ÉF	,wL ��t���M�!N��,^�v0\��M�X�(���&�݌[�OH�n�	�.Ul���=���h�Pӭ��ǗH��x٢`����|؉�Y�&,�c�ڿh����&N�ؠ�N�Rl��%���Pb��0����������D/�&(�&���L�;�IEL��1̎�Ӿ�s>������S_10�2�?X��v7��`�ҝP�Ԋ
���Zl�Q���O_sg+B("�������g��V�{�6"`�����$)D%�*g«�^O6
�K��C�[�*�B��:"z�v,96"��,/�q^�my:К�[:�(�F=_Sg�6�ݥ�s]L�%���yЂ߿��O��7�7�f�ȁ�Sr�l���W�ޢ���G<�{����X`��'~v�{�zO�i6�զ8rRgg����3Em��������C2�K��2u�
(I��T�h����3� �n�X>E�< ���zc�&�hK(*G�T	Nn`ɪ38XD����Kg: ����`Eq��,�%�]�*t	8<�SA�lk>jg����e�Q����P~�\]�<�o�aF��D���q/�@���ۤ�͒m�F����b�Y.��Ԏ��e]7�f5��F
����A���1K���ۿ��z��~A��N��#����K��`~2Ϧ�ż�]���ͳP�������yU�<�L�����́������s@&|�Wh��o_@��W�%}b�g�ʻ�1X�+x�2�c�U�ě����@v�7�B�B�3φ|���������:�� ��4�3sP���;�S�榯uՈL+�,��h����Cs��M5��*0ĉ�4�e�A&(����s �����U�H4�WP�zk<���2:��H�0ۂ��~��c���s��*�G�nЯ�hƽRȭ��F�ߵ�9o�yj�)E���o�z��t�謃��{B�͖5�[OE��|8���E���&��\^$�aqz<��U�x?�%yp2@�4�����{#�+Rո��w>&?)�3�1�KA���c�܀�� ��%F �w�`X}�3���fE���8L�U�^��z���|U�1�y���`��2:2˺��3ُC+N�\ۃ�-�P�k��;"�~�ߩ$��y>E�i�"{3���N��{!#nxl4s�@�L`:p��E�ˍ�4=6)��3��C�T���'�7�l�Ժa{�#�=����'��RU�<�v�71��~#@ի��ܛ��Oj1w�{î��T��e�{$����,�/��p˄�� (eIi���/�}��)
ճ�PKl;n&�w��Le�5"�����ϭ��UE�M*���F�����{@`��h���@�G8&��g"E�g��S��^���%��<��1��2��E��&�n��	A
��D�IP3zh��v|�떏�r;����k����*AML���a�{��}c̉i�I����Vn�oڬ�ݾ�`>�YQ5���Д�l�b\�[�1sEBw)'��{�_��fv�������cEk-�����l#B5O+���_���-н���匯�ïƐ�����T^��\���Ӥ��g�O?	�l6UR��+����qգ�Q>�;�l�T��+����Xm��x�
:�3�$Z��D�TqPL����%���]�>tȳ �r��ʦNG��!�~�J�:���������L.��s��i�
����xo����	��e$<�b��.����EI=/�Û�N��?.��$W 9�P!����?����_����1��ÍW��>��^�&��xV#�g)�}B6��,Y��ٲH5�H�-�u����:GMJf�C�Ǯx���H?Hl��%��3dv,%��p9-<nAr���_�!Z|�3�Ni����cLެ	����� ���8l$O��T1��Y�lE:X��Eܡ��\W�����t�E�ӄX5�`,�H�ѷ�xs�
��֜�#�7��yk��e�|*�p���
}C���F��T�kiכ��8��RK�q*�&ژ���C�}��Hci�3�\oi���&-�0��S�	�t�+��!�B�A�ӂφqc��_*�\M�ѥ@���\�j'Nܮ�"��=����l�^�ڑ �
�3�)����z����m�C�%��b�K������v7Z�<Q>(�I��hm�N��������0�aI=5�Y�{D�;�uA�MT���m���Eh��y���KXx��	p@�[��T�R [O��XZ*K�wH�J����E��
d�x��!!�|���~���Ӄ������e�<���9�2���m�L랧]�2�-�@���Jc���A���{-̳)�Z�̗D[-%��D���m9쿭�<���#Q4�3�#���|+���$p�Ŗ�<�<�HvL��j�5O�*;Im�{��KZ������&ǃG߶��p�ό�0Qt���Z�1��T��q
�cK��V;5YD�x����tE4�H����r@�"u����С��0��Bs/5a����HOk�K�W=��<��`�T��yxC����b7Euٱ�I��*�1ĉ�������x�����nV�C'TQF9К��V�'�� DS��4�ǵ�d�������As���c|`�Ϭ�n-�����S����F�PWW�`��*�?��#�7�Ӱ�T�*��a�~���"��W��`hP;����ˊ���,�	(�{�yjmW_�q����V�*�3L�B�%�m�%N]խ�)�&�ɰc^����ڿ-�0��3�R�|��7o���4��A��h/q}2�[}Q�83��nQ/$֝�c�"�׼ۼD���~GQ����ig��=+th�����
���6��� z���6���A�^z��5QMB"T�H�A".P*w�3�ln�L->%�M1�@��f��w¤���C��H�v�/�>q� �~���-\1ؼ��kS��N��D��:�?�e�	�(���^�uh��e�@�u9�C��k̉Z1�5�}�8�$�0���J^Z�l�u�g7ъ�W��J�N�j�&2ব&Q�z��rZ���X�	�ܮy����c��^�jM� i�Cp�SJ.C��t���
��l�G(��4O�z�5�kX{�����0�կ}�^S���Q�@�i�shZG42�?Ǧ�3�ۍ��J�P�xE(n��qKe�&4�8�yoA	�O���9��M�&�N�������Ts�|�|�q�¼�R�iOFx\�����݌��^��q���L�J�ut�KA��5�7�������χ������&��3O�͍~�7l�� @ڟ�E1Wk�_o��j
�&ru�}��t�����
�[7qtm|#6Ɍߐ�}�{�5�,�mj��� ����h^�ަK߹��BF�������$���{@��O�hQO�z�F|U�#3�ǚ�QC6�@��k����T(�%���J�C� ����i�joٷa�@͘`���u�}��'�Gy1������*�@z�f:�l����[H��r˅Z��^u@R6B
s�tӺ׈�kU	��:'��&�ߌ���43�az�H+���G��S�a ����J���Ð�W��A�$��H�dt%�*�n��,�?�^�i��Vgg~x��փW��_19g9%��%���-zN��u��C�_��@V�߳ǟ4��u���0q}R�Q,�o�f�l��]�=|�.s&zNr����RӺC����l��Uh��q�XK
�ӎ��;��"�d|��f�.�1�̫�po)q 48��U�S����h��|ϗ,|���ľ�a�D��'P����.nG�������7M.�R�s]'��F_j�B�ߥ�X�J3�d~t��� G$�p�D�N�3� g���&k�A:�w<������B~�5��i���]��1�.xT���,��n�6�d[y/��6���;+!��N�G7}+�?ȭ�g����ͦ�Ѽ�M�n��N�|�h�I6M(�{]�aE2��,�>�v�8�y�B꫌�g3�9�(9��ѾM�.X����t��m���kh��MPwM.�0E%ɕ�<\�c�6K�&�����[�Mo!�)cpK�H���Xu&�Ӣ��F�9���h�&�)	�*w��j8�1�9˓7̈`�7	w����h)Rp�<�֘>��m�H��!%͘�`�@�rO�<a�ϑ_��10�V{C�XY��hΩ{�]�9y���=�����`�
�f[BJu���&��ڭ����v�}'o�s���h�<^�g�Kf�rv��M��!)͍�����y���f���ifv�*���ؚY��hze�.Zm��Q���!�"$b8��(U�WV�Z��k�C+���tJWP裚�)���g	�t�O+o�%1�_*�c�6W�/���κ/�	fsB����+/�a<�Wa�$����6Ft���闸Ԑ��w�ڠ֎-�z-��o�3���&������FŞ<\�-�)��t���0TX��]��z����"�$��;(�'��T*�&5�3��a�q�7<ѧI�P�O�
�삞VV��-A�zD� ]�����u��g{I����lL˥��F�V��@:����s �0���������?���@��Fū~�]��Q7_�ڄ:N��f|n�|?Z�̖*<`^�@Z��؍��<d�_%�t��X�̻���ģG��8���et��i.?@���Nc�kjL�>�'�6߸%�R��-��<:���������;!���L��?�O�❫�_iy�طB=��Do��KFͅ��o)�9�O��%��Q?9@_�Y�KǼi|�n���CQ�3V����G�t��t{_+��0q!(�DGg���k+k�u�̞24?��/�Ҟ��2��k�0M��=a:~�eyeX��xL��m��1�p:��	�����DA����F�S>[���Τ���W��t���A5���R}Gwr?�֒4B4�a�r���jy�?��6�A2�5ٶ%�q��Q� ��irT�pP5�9�˱��緄�ܝ�5�Sj�S_>���xOY�UXJK���mw��fׂ���Za�m�1�/ �v���M�A��g��d�N<9�Lr3�==�S7�Y�����Ѳ���B�2j�~.����,�M���tqn������]UѢ��'��N�nF��_f������<@v��s{�+�$�ӻE��<���pH]�ݎ_؍ޯ�8q7�b�}��~�U�6�-������4[d�M�������W8*���
������Py��Ӥ����0�M���*�@�V0�d&���_Ճ��o�&�<�iƴm ����H�Ȫ/%b�l��J�+��b���o�WҔ���z��$j�6����n����ˊ�m:��AG�A���0> �_G���C
�(�U+-M�R?4|r�Z����]�4öp�6҂�;��-^�~�?�0 ��J}�Te@�������\�r�J�(K3!$�i�@|{h�F�U-[#�^�KQ�`d��;���H"V5�F=�Յ&���̦��ۚ���3��K�8/+:ک���� Dx�YQ��a����QN��w	�o�K��+�jXX��Z
�_��nF����	���; 7���A���?[+n0�*sY�u�� ���,��n�d�otY4�]d��<���2gd��S�W?X������b�j�Nq�`�}����Nٹ7��� D칛1[�A�T�t&�kOiya�@�oƩ�-��&�z�˖�@��Wˀ֪�zZA���I��/�hi��-NZlR�iB�z��J*��{ ����cxs9�[r;�z�p� �=��T��7^Z���n�����BC�Ќ�(���`��������jJ�@��8�������o)�{�ޖ��|�""�CE�4X,��M���
��Tt��I�I�:�@�,`	MҲ)s�51n���{LA��A���������8��b���{��0�#��2����<�L�2x��%��dL�3����I�!q�r9q���7r�)��Lc�� ��u��t*"�bF�����fV��<���풧%�@��6�!	��:�O�G�*j��|���0C칈���}l67�\�XR;6�¹sȫ3�/Z۲��H�ͬդ���t�f=�?�aWB)|l�%����w3������d /C�Ai�z�qл� 6���[�����/�m���w�ޫl����r����w����H⤷T��e����d]�5H�g� ��;�7	�M�k��C(2�Pic��t�`�f��[o`|ȴ��)	0��U�>����n��hy�b8+�N�nx����c�����:F�������e���o� 2��^E�8T����(3��r��*.ˤ���:�˦i��Y,�m�7�^����^oE�}v�㴌W1Fsl��gs�Z�r�⭦�PY\ S,�����xA��+�A�ێ �I4��;�)�,�R�>:_�@�Q�dK-g��܋#֡V"�w����")����1��Q�/Q4e���K~%�;X|@��*eŷF��Ŷ��R��ŬN�Q�� ;��rPO!��7�'��s���y-�J�x� �^�4��t���W�wYl�#2L�wz#�jaΗ�"�~U��^6�*q�kH���/L�\��*V-�«�»uV%U ��&ϱ��OHMӵ�^�N����>݉��b,Ǹ�۳�!S4���dʓ�������?CS.�)J����v<ǋ�ޔ°�81.>�YU?R�A3I�ӌW¿�f��^�}�y]]\J>w)�:.sx�o}����x����m.��U��߁ߴ���odpt�}�'��2Y��#�^w�A�c�Ŕ
���~:(N�(���Ɂ�W�Sռ�j6`,\oI�]T>j��7��>=^۔�,c�ȟ���OA)�S!����؃�K��h7\x������8���.i�x�c�9*��Z*�T�$
�H�#Mq:Z�%�P�?��2��*0VV.�|���r�*���\��x��-��6$�hڔ|̛?S�-��O�����:�1@�N��˝�!tہp�-ey�?���W����pD�!�v3�d�3[�]�L��	�퀼8��T����Z��j����H���J�*�྄Ҷe泑�uT>p/��UZ{�Go��=.���YqV��	w_�^>���-F����u��� �ˮ� �0�]��*<���u�"�Ù�<b�νݠ"�%;�U��o�ܼ�����$	i�ʑp��o#b(&�L�[�\����=��**�'��;#�ѧ���5�~����&�Z�(�pv�D��L��q�d�-���f7j�R�� ��OP�M|ꍒ���dt�E:�ˇ��!�֓�9�\�� �T̴��4H��x2Iӭu�������Z�R6)�Tq��D� _g��D0���h�.V��AgL�0+ x�|4�M@�};fRx����X� \`���L�h3�ٷH
�����X[�6�|$#��x��81UU�<�Z�8�dH����k[�� GK�IgYA�[4K �Cj���Vɽ�.+�%��JZ�s2'�C�F�_@�G� ����T :T_w�I����hz�Yu����j%ll�ͼ�(������L���,���_D��A��B�X��9�<��C���1�r@�Kb�{�Zf(�Fd�G���������K/9���ϣhEN;i&1�m���C'��ɧb";������l S�oW�/6q�)����g��YNi�|I��ܲW�bc��􀼃�����"-��! gA�a��%�!��>���y�r�o����3!��l�y�H�c"/E�6`ܷ�jB�p�⽎&���\�q"�oK明��t�G` � !Gb��oib��`�0��]l�h9��VQX!��͜�Ǥ���wm"�`	�}���{��}Yؐ�"�L�׿Jø�{+��6��0�6~-����%�@�R�է@yB�2�����˭�J�;��ж��5��q�0�t��F���+t�����֬��f5�����/��R�^�EG/�g������b8�shJVO9��s5��z�������-�Uj{��@p���_B����m�U:.��O����d*�O��k+<��B� ��^��|�w��Esr"��BA�4]��R�&����7����ٛ���:RA�gy2-NZOG���|�{������|���`���
��ݑ��o��^��Ş?9�6���)�ޔ:��}��A�L��E��G4�I�iT������I�n�P~�9�K#�֩M�l�:5�^I�����_sܢ�$��p4JL��w��7���>�]��2qy�2%�>�se6}(�u#�D�qcͿw�	b�O��fz�6��VT��W����U�`�T��!�[mj]��
k���5�I�N]Nar(A�� ���æMY1!m �x� �tQ�-�|��`�B�Sq��!�ݭ)��N��E�]�^���nepX3�@��m���v[��¥����e�$�[��$�}�]h��h?�~Ir���D�^O���(<�^���@�4��e@N��ޓ����v�ɪ'Aۇ�ŹvR}����5��JH[��C�d~`w������W�I�&�-�t���kI`C���_}l�Z�HD�^�g���4�8�7�_ ��=�ݢ�ށ �""�����@?^�X}z�l���泥E$�6���~2��6|�ě��X�+ɝ'*��5���riB�!Զ+�Ju��D;7mתT����}[ml��)��^tů����8�^6I�+f&�IR�J�t|~��m��a�+Qk轀��6�0��U9� �*DQV�U��nzo��i���DH�x�y��&�ٮ��ua�e�?<��G�+���B��uH�BCQ�UG�<i��[�2��g��ųSx^�F ����>�~��Y(o��A�͜ڀ��;U����>�ݍ�T{�Ej�Rђ@���]���w8�!j�j];�ͱ]��d�jD`��Cro*{	���4�ǵ��X":�М��qd9kP!LK��2� d[t[����U��ǻ�6̲x�{�P˘�0�`
C��b���J��WbX)�_hs�ǎL4Q���~ɐ�2�S����f�*l��n+��Vj�*��r<TX�eo�M�7f�v}����2�7]X2�Hf�ò
�(�hbX�fQ[�ٞ�>u��U
Cbʊ�n�4�g.q�*�]FCa��p#�;�����LORg��'���Z��q*M&qҚ/m�<��Bҧ����z5��&��ɭ o��Sb9��HhE�qsF
�ݐ U��&Mwr0PS�B��4�نyc�Y{֘�V��
����@jS�HX�.J�i�
�芲�<7�M���C&̡�)5�&�(���]M��&Y�vV��7�M~
)���y��3Y�c ix��7������yb�r�(��5�R.<a#�|��*�`��������_f9p���9"$��j�#�P�S)k��V�'�Dc�n���q�B�ڙ�3�����6a�������Æ��d��eh�K[ck����媷G$�[SV��R�ؑ���V�P������t�i%i� Tn��{�V�s,P4�W�>��W�\��J}E�tN	��� ��Suq�u��,@�J��򋝚<"�����&�RC��o�M����	�[������r�t{sn07��8��%��
M ��^�VN��)�t�ҿ�sw�cY�G��H�!�|�š��^ߚ�మ`���`Q�Y�zI�:ר�;��شΫ)�V0�����oeq{��1�k|�5��w@y�7�ݤwI���-�ȖlIm�fo�Ӝ�(G+dNb�hq�`R����u�i�b&M_�w����;H��(g�Q��xf�A潤��r.���%�U��jɛo��Z�af	���w��W�y�\/d
�z��#i���Ǎ0�!^U�>�qȷ�������E���ن6�Bcb�y����4a �G�bn�[�,ō0�U�R\n���`o�I� �w�_��!:a�s|�����:����h�$X����$�b�^�R�
:�Ⓢ�M�'E� �N��f�����yq�	j���|>	.�zQ���p�+9��}>�V��\ ��T�����+Ӽ4F��zr�G	2��|%����^��uQ"��/P��!�Gd�=X�- ��p��,��Wu���:�8`�W[+	6��w�o��h���2�m�e8��9_@es!U����k���+�9͕?̌W�(��ڒP:6����%p�Y��fB�ǃ�!�C@h,Y+�m����c��WTJ[W������,��/Y"X�I[�pe�hbp��R�\��a��_�*�D���B��P��ō�ME�)w��i��R�0UI��'�U��L������߬�iȆ�E��kFoS�$�3��������W�%y�ڴL�$k���VS�"όu���d�[�F��h$W8 ��������Ѱ?�dRj�Љ��=y��1M߿�����PJإ�r7'����3��� ��z5�_(�H"0?��~"��I���gR�C 6`v�G��@|�uvQr� �Z���M��W�J���)�����$x� h����ut�W��5� XEE�*�L����Q�b�g��4˨��r��J�b�����s�)�+B���x��PP#K��ѿ��˽?D��Ea���&'r�n��=�M=="d�#�@����M��Ojq�&H"�4L���H�ID�u%�ă�v�<�W�>r?�NK'�8�K[ކ�pU�M�)�a}�����q�r�U)��?�6����J�5���+�O1gw���=�B��O�e��dL�90� ��ݹ,���l;�cQ��E����E�S}X3���^"���hؽm�ՐmȪ?
m)_�5���"�	��$ڕQXg��8<��ٮw��Td��I�w����c����x~vv�!�ՎaejȪ�WꖮbTV$��U
��l��"�s�W��1��@��(��/NY���]|̶�%x�<�x��j�����۞����M�n��F�������Z�ͦ�|�6�(kSX�ʓ0V��f������_�L�d�=���#�TqI���� �OmD��d���=���_�e�	j��7�<k	s���T��2{Fr�@0�n��� ��+�\(�A�b;Ӝw�*8.�I�*�^*Bq�HS����02�n�?aC�����R0O�by'�<�bD��A���"�%�ޡm��ow��]6	Nҙ��۷�?SRou���:�๸.���q\�X%�������E�aѺ�c�r��)Sb�Z�g�ED/�"�&�K�⒠���J�=��� ��n#��(c�$�.���Ir+�ߞ0Lr���Kz�^�3��	��/�h,*}�j���^�Ӵ
�`|c%��/���p���t�A�A�dV�9��1�
s�>`7Wd��Aq"����.� *��ゴd��9��ع[O_��S�'����m4�`',���A�Յ`���o�3:�]r$��"���Ou:\^&;9����b V�����^�ۘ-xx�@|�{F� ��J��arrjd/�3�GC�Hta��~3�����6V�ml6Bx �9��~Eq�@�?A��k�t�zdLf�:�$�����I��qv	Rn ��ʩ<�%��6G�>�	47|C!/��ZR�/������	"p�fpQ�d�0�R��8ȣ�>��t�(Νspey�ȵ���&?'M��+�4�͉��n������q�iYGj�����-KEU��wW�ѭ�A&��N�1�!�z�B��x*������FZ���>>�l����MF�s��U5�h���WMq�R�;�
`��&EY��e�,��O�V;4-�KIx�*&���l���GȬܰ��+!�N�K��<E6J���q.����z���}�-;��1b6��Ȓ�-��H�G�$�8L��R���2��q�	SB���%>�)�	��3�S��N�D��I��
��%�M4�����o��aE�>����7�
[��0���(�/Xgm���#뗌�f��z:�����_A%M��:!;8�z�u���BA�[�V�tla�J�J|��X�5�@���f��y4��R)I����N����O����{�4w�.B��1��%d#�V��f��a(��A�a[��RrUIy[��[X�,eȧp>l7wy�P�Uؠ���q<����C�*��>Z�Mb�����26v�D�:�kv����<A`��Ӄ��r�n��I/-t�����#A�_m��첻|T�Tdde�^k	_�f�=Db�����9v��g��O�����0l������\.����ڐ�78I���?�=i{َ�3>���豧�) $�kep�����dؽ����a��t�ڧ2�~�Ȍ��c6γ�/ult�_�Y���ӻ��nbZ_���0 z��	�}�"�Y�� �0�Y{�����x7+Z���|�ěa�qNx��UI615����a��c��3-d�2�����AJ7.|�/X���������>��LZ�;��BNF�H-�iV�۶c�;�8�(3�м��8��.���lGR
����J���c�14�ۗ���Æ��UiEA�r��-D��%`{G,���ӝB3 �͎%g�Mv�TiيwQ�W���xƱ[��V�{M���,��mQ��*C�;��*���~�� ��%)եO7h���%���ֽ��c�B���е�tՕ���3I����	���?�U/�3/�[^w�)	i2�>r�&Xw9�J�,�u[��+��s@o��Z�C>�m�D�ݗ���*:���k#��ܠ�4��4��k�[�ک�pP�J"Ñ���Wc�b��|�d�=�kV5�Ԋ�B��.	)w�΃�<�
R"&��S�˱8��S�6~�3� ���~9֕ ����jqj`D'��:?|+�i(;��uї��+4p�au�P����n�}�����Y�}$�dU�lh~��z�O�C�=Cm=8�)����)ggy���J<��}}X�yB�=���S�����I�JW�`�fႋ���W�&Qꓡ�	b�	N��aao��dY\"�E�˕��SǑ��?M�E��f�ɘ��ȃ���-�Ư\����o��^-���1c�T�m��v�s�#$������rT2��|-�<����ŎvF})�DA[����P`����@q��\Bo��!�����ش[��+?����W�aڣ����������*�?��XK �	:�,a�1�1�lO���a����pc1@�tEF�D~�u#��������oeZ\>.�t�8��9��,@�_@��p*u������[v �'[>L%0�d' ?���б�┳D6u�\�_�SPA~|�Tn���{3����C�ŧ��J���f&CY#�����,��=Ej���y�[)�^��9�|'?�]���q��Y����e�rfZ��F�n�F0����Z�p���(RDj�ⷚ�q"��g���Ax0��l4�=l�"��� ��o1s�mc��:�IT-� �l@��Ѫ;8,c���|b���T(h4���=�t���
��>5Ӫg��o�e��L�;[J*?�B��$��v�n�glFb�9���e���(�~�17���P��*�b��O�K�n���m�+<:(��5o0 � �W���Jx�!�E[�;�n#n���`�e�N%���O;����S�d�ꧏ�wm�|Է!&j:�Fd�3NN�qƸ-���=�e���ꡣ��
Ȥ8%+�漜)��+#(1������Z%7U�� G�������P�W����@zcr{\�X������`��l��4�h��F��м��d�Ɋ_�Ps��_��_Z�_N�+ �N��0 �����j�4��8��P����i;[�A�W��~�mԐ+Ž������!9���.��"�3[���5������D`vW_0 
�7�z�%�D�$r-��,��\h�q�e�`E�P�6oK�<G�y��6��0Ħ�,�r1���z��z��ǂ=����TG�ԥ�a�O��n�#������XÓ�U�����3��Q��KkX�0�?��րG}%��#"7\������ݠ��J���Ҩ>(�E��BsBٙ��=�ҖH#P�}'J�K�]ٿ�k)�;��l���lp����,f�{y7�yu��<}~[���;)�������M����t�ԔX��ۯ��Mݹ�PS�K��k޶N��ݪ�c�)���#P���i[ڔ)��!��V����X���L,��H�:�J�.7��L�_q=��äT�?s
e_WtF&��:��Hf��>���}.E�L��H��tToR2&�_p᷾��}��	4UL�}�p�d�������Q	'}J��uV�)_�s1�BX��,�˦d��T��<�_�m̔������M��"�f�G�����`/�����I6�7=�_����Eue���E޵�KFາ�]��~m@&����"ҡ~���p~�q�#gv��J�U�	�i�`�9W�:uwA��֏,Qm$�T�;�?���v�y嚉�y��<n�D�de�"ft��UXY��k�Ή̄Y�Ϫ�!ek�GL.̴z��V�:s�h&"��wq܀��R�0V,�<�4&���%������S�0��h��P�nn����l, �k�0E�E�����h��hQ�s��[V�#����DH��/�$�:�F��i�>Y6�j"��CaY�R@�M��s����p�S��˝(R����`4��B����O�����U��-c�J�2�����݂�O�}�F�s�~u7�K7q.�:.�n����y���d&��8�WuZℌ0:񘻻
��G����r|E%^��ؐy\[�>:�2x��0>���|�.$��.}��4Jڸ�����u%�:����K�ҟ@�R������c��F���/3t�;��)���O2�YM�ۅ�{��'h�0��z
i������}���c0 {��K����n�C(�?�������V�R� '���Nr��	7<���:E}�_����ܩ�l�K(iǓ;rB��񃦋�LC��-g��)�k$�׾|�Ɂ4`d7��I�����h���v={,�֓-�&������T<�U����	=|�f6�0� �������*�|�o0�_�hu��Q����+��~�?.�"r��� h��E���Ɣ��+���M���G�r�ۖT��I-����Of���!;a$��m�.ji$��\!��-�Ƌ��ZQ�O���(�I�m�܁�Z?y�?3D �J��8j*+N<�3���㘟�F�QLy�DIŽ)��AdPvb7��Č�izr���L��;A�O�(�k'��̘��
��*�;��٫* �6�1*q��^�����N��h^����YI��eS]�|r��&R�/��H���M��|�7��xa���n�=��F���]�����i�����4Qg�+���A��8&��a:��ǳ�O�wя��e�ϝ����_x�����eu1IE�E�?�E�\zHR�cu؞N�2��͢C(��7�Ҏ*��=�ò��44�gL�{�aN�{���MB�����LK�͋��fVsW�[��[���,N^�ާ�@$ڭ�	�r�b7��<�4� ��!qH��D6��������ƥnHo.V�=:M֟�B ��n@��O��ڍT��5�{�fAN`qI4Z�0�8��0c{�~���p�{t��݈��{�k��>��u7K/Z��(�0�W��I��;C�=�,�]/���b蹈{�|җ�J�3�m$�s��ES"w���u����
7���D��[��T������G�!HT�f��u�z��bUW(rH��QZƔ*D�����O�ۃj���x��V/,��E6�~�z�g���P���.	=�X2^.�}�r+��yz��I�P6[ Q:�Q_��_%�O�юX��#�Zz3��c;��H�d%��w�#�Z�lI&�7�vi�Ѣ�4BW�Y6�^	�0Ej8�G[�Û<��5���~����q��s llz"�?l��7�$�j�GҊ_�	o���s�yx��{K��P�%��q�Vi�B����L+0�a@�D=��K
�{�lq�C�E�N���Z��ǧ�1q�OV-�-�fZ�QQ[ߡ���n�?�nd)���}������d�L�ڕ�
��
���;3|ҝ��1��,v�����ɕ9�A�������~/Q�[j�C(�5&
���[+�A~b��9�(��Hz������؆c����+3�����d�;h!A�����6��u��U�@�o]�T���ZQ���l#�խn���b���2�6����v��}���ޢE��أ�}�*n(��\t�"���V���)���������UP�g�a/��6��@M��V9ZC�OnO�8�x~�fn�)-�yo�h\Z^�b��}�TPĺ�պ�pv�c��W����P�n�\���XXD7��ƅ�-�9�*��o3/P�����ܺ�B���r�kA�1�S�/���iĻ�t���wR�g�YW�2�d�6�*�6�.$� ����_M�H���˩0.|������s�Q6��z�`��l��-߬��5�i�DT���3�&�����h�3�jZu��������3��g�Q,[�̥x;���߬�ʷ��,(���Ĝ4E����z��Mұi�E�Kp�����2�*���"`%��Θ��h����.��zc�O�������&����tAP�b�ց��
��/����d��������Tk�+C�1���5
�	���sg�	v�v �)M
�V�0o�*
�06洀���J����Uw�&�;�"�Y0ن��l7E���f_r�f؞�+�+�Q��^l3eӝ��I��@�3��<Y3V���Ը�g�k�(�YS�e���4��l�f���R�e-�������Eo%��T�@w8�	��y	��,�����1�\~m�L�I�����K r>�W�:.��е��Y=v�x�|�\����m������a���Mqo���&VʍG�� �ȼ������+�[@\d���%)�pP�+nq�QO��`\���XBѭ�z�h������>:�KK/��rwjޜ<�Y ^B7�
:�����+��zv%��b���[�����(��
�G���%��!�7��Y���1��B^�(<F��OJ�2@�g�n5���AAa��jmR��,�F<oS���܇����@O�nD�n�#��V��Ǎ皒G����p��y?���|ީi|�A:J9EsX��B(����7�-��۲"v�Ą؃buR=P2 .ϯ)�����l���.x�E�ᶖ{��(�m6d-�f��[o?L==���M���.���y��w]����_i�ü��(xh'�WXl' !�� l�a���l�� ��8)i�a9����m��s�!�h�ȌՕp�q�n��I�U����+�B�`d�Qڕùl\�s�\��8��~��^�zC���W �5��