��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�z吴�)b���ΡrϷ���	�J�*��hm�E{�Ի?1��A@9VRt���0\A"�6�o����g��L�Q'!���y	�y�n{��"��shJk�%����Sx[��w���v]�@�:��r��J'5�S�_l-��h1%w������*Jm��'�se�<�Cg�x\�I��j��
��K����	���LB{����B+�m�3�W_��7��Ҕ�hnoF���;�V����aoa�������]�;�p^VKC�A�=Վ�!�Y��|!Q�t.�7��$�JC�*�S�̹�XA.wA Q� �:���1��lA�P�cgAf��S����11�����4�Ep���F�J�+T�>���$xgQ�&�+x�F&JJs���Qk������If�}í9�Bl�cR�K�o��&�,gn��)A
��v��=�I�OC��X��k!R��B�̺���Z���^I4���̂���	�
��o0�m�V|�AB�S\����۬b��i���8iOk����B��p�1�5�r�t�*:d[dT�߄��_d��o�ehfDȲ������r�*xD�_�G+�k��[mr���d�,�+�S��dZ������Ѡ>�ݮ�^
+����ɑ!ɸ�����+��{��t�` }Rx��U���A��Mɏo��0��6R>�G�4SX���ޓ$�y Į�')��P�pۼ�v�jL}P��~��r:�C�J9�35�"���\T�v�J�.2���с��BR�h��23է�5��?�&�J`R`��fY��i�/���DF������%x��٪L�OR���х�H���r\��.�W���{@sv(.<V�t"l$�����+��E��pŏ  rr��r��@Hw�hfFn����3m��y����M}�����0Y���7p�& ��|�B.ƴ"^W����+��xgҘ _\�	p�[8��I���������F�Y�N����D!t�7$�vA.�,����00�B���Ns��z�M��8��1�v�=�aXP�U�l+ =)��m�X�����ʆ5�.Y"���{җ#��0ޫ/���|���q�z��L~u��x� }�0m�6��]�TP��^�רb���Д�B&��(S�C���r� y��>���)8�+���$�%�>c��qh3 \�����ሲ��sl����B#L2v���Fb�� $*vpGے7�
LC�+�Yb�
i�]tP�ʒg6�=��T�&m�k>U��PIZ��Y��s���d7�B�Բi/䥣ф(��=9���\q0j|����˦�E�&�?h�|��$�M[�M�.��Ԃu��ޙ�v�q�<�?֨�\���FvG�c��^�c댍Ng,x�!u��V!X�+�M=�=� �x ��]�m��:��'k긦q�ȷz~d�.�<"5vK��
��c��@گ��+GZ��P�͓�!E�9�������Sd������K
S6HqF����v�?e�0l�T,CN�?xt�6<U��M�^ޙ�~³��:?/���xK�'�ѢK�Y��҉�Tr��`G�����5�z H����D��p�Do��E���q!܈�l�D*[C\�Ӏ��Fx�Z�w��u�b$݈�	H
(!Rp9���4��Q׆���4%"���I38��M�W��@V�5�Lج��z����lt���8O�����EO���4!K�9Hc�%�@8鬂��J�v}�����4���.�&l��~��a�zϏ���;%��@Co��,�5��U�r�t���TU��{��Z��OO� ����]{F
&�`�+!��kE6��-���:����ωT��Q&���Ke�i,�EU��u:O���� ��O��u�}�LOg���.@�EKP����!�J��Q��}�یD����^>@��Q��9�jP��H?�f�`>�*G��Һ,l���~��c�-��~�|�vڛ߶,9~�_ �q�)k��(�$C�X�gl�"U�mSS��s	��������i�{�tTQSje�ګ�u������c��ݘ}y�N.��u°����;N�j&�F�l���l���xy�,���T��d���ڨ�#�+�n�ꨵ�]���]����6�jU�mTA�\��%P���{?������5]��)]���盷7����:���)DM�'�&�ω�0T ��xx�n��X�2�qtxA���TNF��!��y��U���n��O�В�s����OHKS)���o��q]�����#���J���<���������S�������ٷ
�P�2�st7L�o�RI�����gBeG]����K�ܛ�IQ�Q�+�L������-W���3������N0G$�n�_%J+:c���ЎA���]a,���m*$
A@n����Io�;��о�~���K�ɋ�	/Il!e��Alw�	�q|.ٞ�b�\�ՏDX��h�Z�0��N��(	Dܸ?�Rx�q���Ǣɥ!4(#Ë$�C�DD���lX{h@�ϵ��Q /ۤ_���Yu��$�RJU�&9���%��O]֩��ki�מ��ഉ4Q�)�M.	Q}�>{۶��E�����D���0\��նt�{�%)9�a��u��Z{4#+�+��[Ff%�b��g�R��|��$~]h����e�}�ަ�W�ċ�dT�B `��?���������͞3q�x=r��V��M��$��-�>���X{\��$����~�T!������.�%���j���2\/�w��م�e��?�r+*H��OېL�oK��~��#e��a�YG��n��,|�;u9��K��� ��gfI�u_�{`v-���08HPݝ�.>�ͯ�w؝�6ɭ"EF�s7=��~xTX�lR�`���&J�}{%�o��@����ї�Ǝ���S�����É��n��;yq�wa���^S�Ƞ^��@S��k�Κ��Jw�o������ֳ�1Y
<m �0)^1��c��H���F�����PC^إ۽t6a���E�\���:���Se]�!ҹ��$��p�m:�g�B{Y{hM���ҋb�X�yr��+��m����nLY��[[$2��$8��P�D���s��̴��8]eP��*ؕr�s,d�W�� �~�/��Ȭ[]Sz���t�❇"l�C��3��0�T�~�)��|� b4A Nٽˮ!��[&>E2�1��)��%�*�hu��Rm�d�//����+"{?��1b��W����6�������l/�k8�O*���M�WD.�6a�J��l�f�ߜǩ���A��R%�n�������O|�ߨ�L�_xת1�H��fX��5�j:(��d�5��$� ����r2x�0'���~��G�"�k!�r �;i����{����&��2���3�� �'+�	��Ħ�:��+BDMbOpL�|]�"��AW���W����XJ��n�P��5]d���(��b��5�M7=W�/�f�#��R)���T5_���|z��}A`��$*��S|�C�h�E�
�����T�+pP�R!�*P����@"��.�9gaO@c�ѓ��'�3��Db/�Aa�#�CM��H�.	����g���qʄ�N���1��:wgf�\+~E06E,�5(��/+%m���!�O��-���jd}��sn9Xdt7w�?{�[F��'7���!�V�	�nl�8w}@d%�Y � h�]����1`s�����[�I�b.��9�;ެ�(�kri^�b�'z��vܮeN�x����gL����=�)t�fRZh	B�����U<Vm�����R%c�O�V��ܚW^Ci̺�+��{�m�l%�"/:��V.ת3G)5�,R�<�@X,�N�������x�gN�V'D�)��Z� ��_e���@5�^���\����_6����|��ߣBA�|���=�[ZHi���Ix��I1׋��9����c�����u�E�qH���_�tY-b'�ᣒ�2ޤ���Gu���@�:w�ڇ�S��1��ˡ�����^R�If�����Xޯ�V�g��D��=��V�xn0`��D���]ˈ�쏱�2P��%a6�4������E�	��Yde�|?�fGv��B�so�i�Y��>�B�ZE���H����Z�vt�peHֲ1�?�v�K����c���K�����JR���z�?���n��T���e�睃�����P5V��;����y���n1�J��rڍ��n2�P�1�#F*CI7a(����2e8ł`�<�椁���$�J�h�k�K� �EYa� ��o�w�(И���J����"��}TWp�/�oˮ�$����{�C�c�Ձ����=����q&������ZA6L�X��V�6��I- �%<��6�؃"��U���+��1��	�z
SҭL��M�z�Ѷ�S��YEiDK����AR^S��ɝ�]���1ѭ�jX��D�@�c���R���b���&������t�he��{,��E�
1���� j{IȜF�cM`��Ҽ�@E'�2އ�\�~E��j�'�x�T�P]+ᒙ�0�`�։��
$��׺��!��$��Fv+[M��8r|0�Iz)V2=܏��]�߷I�tZ�GߡЊ���dYu��;ʧYE���@�bE��~K �˧.���Lͫ�7�˒�5@�@�6�<�إ�#V�!�_b���������k����l�����ߑxC�hP��N�s����ep���:�͌k͍�R88IXP����t����������IðL�$�;���w��t�Q'u���6�U�Ĳڻ �\���ĉ-p�)rz&Ϲ��Â���ʈ`�қ�M���ᚓ��J�yV�*G|Ň��E>� ���/�w���%���g.0-��e\+Ķ�Q3:gIg]@@����\o���<�Ɛ�Z�B�u���fO?cH��M���|Kz*�Ë�+
�-ji�.�� ��FPG��f�1D���P�#F2��a=���ZeX܇�70ن���H��n�`!�#�f�F)��f����������*~<Dڰa��z�����ƞ $]j ���˭�1)d�
X��W�ϼ�Ҍ7g�<X�=��W�P�E�Y�$Ta�)�|Gq�ሷ1\I���-7�қ`X�'��|,�$&�u����n�x�C_=Bﵨ����nWZ�i�W�
�Ҍ���g����Z,������L�m���B=�LA��؞*IP'�P��$MPe\|��4"Ly1�Ec2��X��)R���p���{�UX]��~���3��ѣ�C�+��*I�<���Ͽj�щx�Λ�lO��_�	�g�@��(��s����R׍"L��*n�|}ǐs�X��ME�쾟�]t~U{�d�,>���'l�r�,�*3�vn�[i��f��ɻֲ���YGe�pp	N��n7%+������y�p��G�b@t��{�ay}}�j~�l�eso�k-� .ek�Ƶ~۸��M��ݺ�-L��'d�f�l�/�3E��6k^�Ϸ�����\����|qtv��z|��'�u�T��⋍�E[{�p&w|�bD�f��x�s�d�;�������������erR0y͍�EvY���2ힺ%C�����h ""Z�z��9�e$|����/��ܣ��l�3%#���(�� �abS����K����o�*�`���4c�����Ki�`$珦�>p����X���[��Pg�ѺP�ft�{���8s����y��Q��W��/+[s1��$f(p��G����M<�/�q1]0\|mQ��޺(�M�E��!o0��+�+��D���#��*��0F%Ip)��b�Go����	]��[�����ϓ������:�-c�8�a)V�,y�ޜ#�>%��M����xu	�&a����z�E��΄9e�"kӞ��MKE�s(�}t��}�;aT:�,��E��3���c'��`,^u�Ub�HExWdh���Q$�gXnux,,b�,@!�u4������F� D�zF�s��C�#? *�׶2�4�8в<�"�j�.8�-��T���=�� ��/#��*C[N��Ho�j:T����҂�:�j�GJ�u��'��z2v�g����miE����D�T�\�$�$�*e�3�E}χ���(]0�nf됻ZfL{�ܥ���v�*����}%mv��7��t�J5�φ�j1(j<>(��*	T)W��	��8����-ڎՈME� Έ�Wg�A>am��/�Z�?U�]�f�
r~$Y�ća��.��t���F<���s�ȢoY>�������e9	�1����=Œ��|���U}�fi�~IT"�K��(�u�"f����mÿdXx�2ͧ~��A�u�W��)��{�^�cg�� ��x�)H�@�T:�엉H�_a��4f�A�\��xϦ<��0�
��%������*'�_bg���/_��M��*���'?���?5O#���ښ���U��"�n!���I;|U�8�y��y�ծ�I�UDD�5K��o�4a	�n��'�S�Vv6���/<.�<�t7觖.��7(������~���s�t ��,>�D�dO!��^�>1�|A��k^�ǎ��0����4�\K4���L�.�{�F�|ߞ괊�m��*/�Q�@d��Ϧ��Ls	N��槍�c��zA��Eoگ�O�?��"�H7����D�W�\{�<xcV��"�mٜl���Н�/�z(��r��zRg�g�;4|^���gű|������l���2�1J�C7Yhl`��v�\��"�٤6�a�
�l�!Z�b}"	��*�O$�&~ɹ^�3N��ok��I�	���W&`u�������)�2�|��*!FG�3ܩ���F]Buk�RnI��_��~�(��s<�-��=�f�ri�����7����!����A{'�w$�CU��D��<^�����Z�c�.v�.�q����Ѱ3kxG	q,�í0D�"H�ފ��#��S�_6i����'Ka�2�x�	˫Qz�n�5`�Y5�-R��Ć.���IOdzE���E�$�_1(�]i$�c��ue�!�T����A��~9�s+���$p���)2̟L�Й�� ��~��
��S�?�Gxek�Ɏ�(����������\ǹ�;��$�P֙>��܈8��;}{�_4}'����[5lL��'7X�=��a2P���O����/=�]�
.]�n���(y�R|�,�>��Qev�#V� 2�5)���ν��`ޘ���V4�	���N��<E���bf�0м+x,�)�Y�e�����&^��7�q�A��űn�bK�/��3�I嶙gɸ�>F��T����_�p|+���/��8�q�������~�(^�:�xgZ,=��t��IU�0s�������d��L�p�2�^�t*�� ��#�B�_���"��C?i`�o*�4�%{����z���D՝��4�23�3�uLIg��rЗ/ ĮEʈ��d	���2k�_J�恹?^p$W��[�P.{?ҷb7�R
�^3=�oa�
O�2�ح�f�8���)
�O��j�3�s��|�h=�I_"�A���aك�_F����0���#���WJ&�#i6��E �C�&
e��=��y;?�E�-T]�""zIо|�Ү�6�`oֻ��7����]�+�Y,�^j&��[��jxD�Э�?Yt؅s#.3�
���$-���rX/\̾�k���r�F���P��&@1"�~>�J�ۯ�_�;��lm�$���n�f �@����2���\1�X�bޝ#�n�]���Y���(9���U�rG��oxVfX�y�x,c���5���T?�*��H�=/��ʉ�>K�>{,ϸ�%?�L��*�:�ꥉ�3��`��~�5J�}�^|[��V��P�7��ȐҢ��-K�<\(�r�P	{76V�+�X��$�v��U�4�a�̰<�����O,�]x��B�8C��$U�����6D����f��y�~��"��J��p5��z����{Q�G������@�{��)#�a"Ƌ�
�E=�Y����O��ݘqL% ��.�5���9Ǹx3J=X�t������Kl���,cw�i��éצ��PڇBK����Ry�ђ%XI�`И�p2#C~�3ƈE�7���S��Aa����5]߼O3&h���I�DE+�`�)9�pq9��8.3�	GrM��y:5b�n4qLc�(����U��oT�լ<5�F�;����� ��zlK2�3�h8��Q�p�:����娤 m��}�n=�Dn�qNxp�?�X�F�=�g�!:�A50�;�e8m7J�V�o�R����BE%P��8��/����F����>��(���:�����.O۷�tJ:ٛ+q;O>ӝ���[H��m�����������%�#��)�E���_�>��}9����-Pǵ���/`��D~62I|���CjA�,��N~��?�������w��23\AmC�f�w(;���Du��0��H�[��T
�I.��D"��|�0�z���s�o(=�A�Hv�|/�k�X�9��6eؖXR0m<�%9������c������DnտLŸ��ihys����Z��-���>���X�Ra�R ��Τ0;L���O�ηf^��R������נ�u	/��S*Ç��sq"��zl� 1V'i�H��S\�&M/�A�ƕ*��\����A��ـ��7퇿��E�~ț:O����x�_�m� 
r?�|��_Ă[��I��mY(�6{������@������
P�#����
�y���s�t��Pu���� *�SP�h\�ᗿ}�T��x�#)��<����؁��Cg�Y���ŸOęT���W6�1ʨPS���ymF���	DH�Y���C]��6,!�贺�6������ν�hi@�"5N�;���M�Ա���O� ��ܚn+e��{�x���Zw)\N�F1�]k�*�`��GQ�L��ZM:kQ$��~�rA,�I᷾�P�?r���L'���t�dśe�~�-[�f��zGb����mķz"�+)T��:�t%�~g:��1ICl
z�Y!�=ܘ��c<!��JI�R�I�ϥ�"����^�w,��b"�͐D�~A��
���%�����<�Ϻ|����o�ɥ��j����㎧ ��"��ZF�Y͎1���;9�����@p~� �^��@j�F�Vd�-�ϗ��^# /k�F��񊟑�>�Rud$\�+\�
�c��SM_��B'�b�-~b��o���OwX�$ �Ka��f�n>��t��pCGI��o]a���+�����Tb�q&�͢��݉DC/��p���z�c�a���aȭ���RS��.��P>�;wr���������#�� U�C�+�(���d��1y�	����{TE��@R9.H�EF/i/3��u��qP�Fr��C;(/i�R�E��B��2��f
3�:�5����C�S�<*>G�^��_$�D�C<�(����Y��51��as�Dq>��\>���íz~�iB��`�?�ACu�<�n�w�F�9�~��*}P�3t���7I�T�@mךQ;j�E� t6�%d]�zra"��6���1Chwg���hd�wlg8
	d���t�ߣ�GyCK6Aw�=���;/��/�+m�V�]��~�I	�遚�����sVs������/�51+}-8$E%�l%c�vwul�Yi]-ٮ�e̳��_x���g�׫"��HB|��3~v�j�V�����Bͯ��*���)����+ː�u�1��Q��?��ϸ03y��f�6�I�н#�]K)}}��):�����X��������b�����R�70#����D��W�u�,��Q9L�����y�$@��
��,&����?�2q���o~���R���-�j��ʩ�")�@�Gf+P�׾�����w��e��ƕI�JX*@�#3�$ڊ���ϼO\��s�Tc�sr"�ǜ��Ru�
��[��峳�O�/Q�p�䎶R�INl!�K�|�Ұf_��o{�R���������7q�O���W�٠S������-bY����4%k��bgx>�=��P@���(<;���D�ʃ�=q7�GV�t����i�Gsx�k�p�,2��8��/��_��,��r{�woj\��OQ�`��0ZH0y]�톀q�_�B�e�{Y*+5*���/bP	�����������;h�+J���XO=xi�!H�⺺n/�(��b�6o��b�� ���ebK�o�S�\6���Kq���㔆V���ȗؿ|�H߇��^�0s:��Kr�Aߢ0AӘ�j�V1�/ռ��)�5� �D�����]HL�f����%{��<L?�*r|i@��5�ـ��&-&���	��hꐳ���`.�Q
��o���3�q�/�|�֎�h�́Zl�3!Ȃ��_��t#]���j%�+0�3��~S�iXjՅ-Jl$��ҹR��Fj�18�(�dq?/?6�hٞ��r��\NDv_^R�C���C�ppDE0��'���b����p0J��w�π�{`8{9��ˍKDw��-�u|0F����=9pqh�Xr���PsL�?*?���{|��Y��k��-!�Z��s	�k�H'�1�$��
�V�w�f��
!Ь�Y�'�aV3�D�N�L��ٱߐI��"�k^�2�p�uX{#�=/���fC*�	� <k�V����co�M��5F����~t�r��z�R�Č�<�O��CbD�����nV�ρ9v��h��Wj��s�t��N0*x���>��zД1c�kI-��B�����gҟ*Q����^���s�����Sˇ�:0i�.8UP��W-L�JЦ����5�!��5�r����Z��T�N�V��Ij��Mу���&Ҵ&�S}�<�WF�˙�ĥ���i�_�S���P�ú�'��욛����Tz7|b��5��p�%6l�]��8�Y�п>�g�XR.B>+֤;8=�����)��}����\�%vo����q���y�Ӝ� �
��8f)�{���"��NC�{���Br��J�ˣ>���|�n��g�y#�g��YtR�Bu;/��.V]�f�����I���<0(�)��|֐�^���t q���E�|1����-6��Ə�� z:�SF��<�7�<�!��hi�uZ��ی�P�/��_8�R�'�t��FZ]s��NO�V�v9��P� O(v�*cy%P��M>�9έ7�R�(Z6�%�ۡ�n�d�}�á�/+��X��NM�1Af;���c���
�YT���!G�T�r�c���oY��̂�{�/��%�թ�U��-�s�?�M���+ɀ�iX6V�3%3=���J��b,e�_�䢰�Jژ.Zw`�;��;!1?,G�U�µ;>d�&i��ظO��~R%�~'�G0�긣oLv�M�s�)98�F$}I-����#���=h�LI$A	K�!��YԺ��M!�Kk���ɟ<��4"|�.Kp�=�]��U��Ҙ��y8��C���z�(95�z��ضX�1�f�Y�Ǩt��Nơ�b��*N�7���Z��fw�8���X����8��7HF��O��>�ߨdK�|Z�E� 7(�go�Ȼ����`4¬��H�Ҽu��nR�'��<�W���mu����ɮ��p�I*��t?���օޚa�1��N7�!>F�Ұ��s���_vq����3�����$�t����μ�--�]ۀ�Q�F�	�_k���]I��sT�(shӖ�2G�+R��v�]�)i����:�z��+$�6C�v)�E�$�WM�[@���a{�i$���|?̧0�0?����+��l�y�G# #��r����(4����40���6�V0禹NI9A�N����5�+n=`�!�8��*��K�p��-$�����w��ć��V�MZr� �^�y5d��3Ǩ����v#��lp�Ge�MV0ə)�`{�~Z�=cm7�+)�VQ�4�Q w��~s�o5�Jݒ�л�lUT��%'�bz[�L�B6ϭ������^I�����՚��Du�6A�ǌ_��iG܎Ycgѓ�,����ky��wm���������O���a5C���:/�~���K�D$?��6
4��B2Ղ��d�$��q��6���~��~�,�iCp��N�Ŷ�,E˅�;�AL~��?xn��Ko�C<������A����z�gjn��gI஄����6Y9ҺR�d�`�u�(���u��^%�V��LN����%J��,ƹ��Ĝ���1�ƚ`!Wk�X�'Gk�q�	$"J���� ܪSC��m	��(����%�E�g��R�~˴���_�-���M����Q�LB&z�{B��s�d�Z������*s��I͏ �U�Bġ�A�#c?z ͍g���ɒv���)��f��oqjǙ�J�+�J���5�9Mvyz�VWO.�pծ�Eal�D?����}����(p��I�1���	�|͑�v�\�H)S���ڂ�hU� دcVH��.���s��6��8/"���;$��ϙ��)]�~�JĐ �HN<�t��%�z���k�&��n�Ԩw��R?)��<��J��%���G!q��D�N�O�T�M7�r��3Irʠ�ȳ��Q吅5��S���X��v�e+�N���Bvq���Q�=���o_<i�]ߟ����I'Eb0���������'1�@�T74�8�kFN����#��w`6t�}�MU�a!oJ-�d���8.�:v$�f��W��G�b��s�^3�B�&H�BAt�cѶ��k�τs�]1�^}�{!z�"�@jb)�