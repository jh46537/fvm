��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-��j[w�_��}��͠Y��{�7?-�"xd4|���j���oIImuz�(P&ԘE�#MIB��4�[�"2?�ߘ��b��
�	o�ID ����P/����*��[�I��e���Q'�i��H����a��Χ�F2�Չ� -kI����D��ԷK��Lhñ�������p��k�f˩9��޶�G7jk9۫��E����7�	���<��byq
J{�4��"�0U��;f�Iw�P�/�pK0�B�|6p8��/�1R( կO=jH%ך*�ƣ���f�a�����T�ހ_6]d�#�4��xXa�E�ƣDR
��	O1�\�FȊ�(���*�c���r�"5[�\��y�7�v.�u�"WlOH7�QQ���i�qX���"��᫜uP)U�8=º�^�u(�k#;�@�,��ڵl��c�&���t��<��Y���hW�r��[&M'��V�hNz��,ˏz�`���d�!�ad�P�o�t����$��rLmp��.������z�';�����i
��o��}]$�FX��t���w��S��?m=�v�);�Z�+�:���eƵ�@�X�S��1d6���2�e��I���9�9�i�7��S��=���Ɨ�&�Ǣ�L��,̪�'L���)�6ǫ�W�r\�_�7"�$p�--�����V�e�vйԖW��� 7�.O���ێL�Ǹ��1!�oPT�����
��Л�*�Am��4��>0�K�5r2N���z�L���Ҥ"-"X�B�%-��Fg�H���P��Jv6mz��y��/�.ZE�^V2`}��O��Z���DB���v ��|�נ�h>��;}ڠ�8xTrM��h���ɂS��q��g�Z��UH�q��Uw�r;@�m'��N�(����p�F$	K���u����&�A��"?��Z�av%��b����
��L2����jY��9�O Gc=�{R��Z��(�r�Ȣi��&���\�d�V��oLx�����x�;���oA��\�J��9?(��.-C�w���H�V�](���~���~��s��Q�J/��o�&^���.�W�3j�p�N�	-����6�AI�v߫]�CLT�O+`)��aí�(��>��<���q��2�w�p��4on���F ��|i��6����8\�EP��L`J��}��7M��C�"; ��<~��e����<\�������Ԝ�"��,�V�I)�֫��\�M�&	���"���i拀@f�r�_ŵ� KF���V�^������<�>{����#�b�4����g�/μO���Ԉ��#��*�^a.5a�ѝ,B�I-��{Pe���?	B�8)�LfA��x-8�Ul}�W��  Cb+�?��e��G��裑Qc�TG�@�{�qrSCe[F�.yz.�iaC���m�8� ̃M5Ȼ�7��N;�����h�p8$+���ќ`�7f
��Z	hȨG�Ro��18m��ʔZ�/��ϒ��­�����Z�,u%*���
�Q^dd��~4ه�8ޙ���gUX�Gt�l~�bo�'y����Ke��o�S���S
X/����\;^kd}p��h�������FV�b�2D�]CL�8���WF��7�2`�Fsb�T�g�w:��EYqt6+��F�W&����O�/��&�2S,�+{B�e�2.~ё��z�Z�lqcp�S)��K���/Jα��ɝ�9�H���30"�b�b�O�s>vA���j�7W����)��k�]�4O{]���^Me뽟c�>�S���Ӄv�q�>�8Y����4i����$��tМ�-b���qpr�oZ���Gp�[����ܰ`>�T	X�2��P���YGe��e@��^�W�S6����|wh��D�1U@��Z;��`]��ʩ���
�QC�:0X��Z� `�OF��iǁ������Q�-)��j�f3�vƒP�Zٱѽ�ѝ����u6�n�L%�1�[�A���g�"t��I�'����g���R֩���`��w�s��]e%D��I� 7�������`��D�1E�Lz+�{?6ƣ+I�I����	X�О�`?ݼE)R��7�jt��Ï���o��wX�axV��Gm�r�2N�%�S͋'�	oﭪ�먹������UKs/~���X���f�J�xL�E�.i�
�{�o(""n� |����F�&9+�o*g 8���L��w]�]. >E��[�MΣ��֩4�hxO
�.jrS�>��_��;.>�u�Eq��WI2}��mt�uk�/�JW���Jr"�+�GX�~ʂy�W͘c��=c�̬R�iT�"�g������2����O��-Є�q���\��Rc�؜�[{��z��?�K��䠄.0�t���W$T�>�}��t~���x�����C%, )���2����ʥ�R;��/͟��%��)����dT�qhK]c�1�D�� Lи�ՠ�WN�í`*�����]�>h���; Tq��Т�Ζ��t�9�#Z�jl�@�=z���H�H5ܬ�cp/!4���<��I�X��pJ� �LJsdٲkJ3�LEV+(���xa,$i�s:K����FV��e��4NԬ-��Pc�\[�d
J@�F��G<����������˸�u��F��^ra)