��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,VI�0=�E��Ӫ�-N���=��_�@Q�:�7�����n�KyJPq��QIVC|w#�18������c
�X�e�n��8��Vgdz`*}��LW���$�s6�j�E�r�bǙ�����.A:�U<����Y���:�*��^#t�2�U��0��d�	�Y���W`�A�<���������(>s\�#W��Z���XgG�����p?[5H#PuD��SW��������C�|��:<Y�L Q�wp����f)�:��� �.+E(��[��ӛ��=�=*�<��}{/����-E�3t�d��?N|x�ڭ� 8th?�m#��5`�*%v��7�G�U���PJ��=���D��qPS�d����/��Z�W䛊�D�6hfe���r�M�=�H���)�C֞�(�q��IJ�b�U�8^?a���k3L���˖;ya�{�1졨����M��<95�IsE���j~M��
��6�0��,�u��_�l'7Cv*����]�[��}Q�8�Fۮ������|SP���=F=���x��{k ye�m�u�@�܇1��Tlmi��zN��q���pXɳr{$���Z�׍֋�V�?r��H��ӡ��ڨ���h�B��/u9��fwJ��n����M�E}�ա:s���ep���G���p?���~�C:��b8C����>��������%�-����_	�Σn�_y��
X'���}�I3� ��y:f�>��!��<]JLFf�i��I�0C>�=�ah �O�g�^~�-��+qE~�W�
Ke�TƎoˍv����L��j�ekؿ�|8�GLDy��[��.*"p�(^'��a��2��z,�H ����V9�߿�����:t-�Kp�08�]8��[6W�U�)EUשil/,\����qCm��QN�BfM�L�+���:��/ 6B4y��J�����F�
�(գ[u�6��w�&�tÄ�Y�LW������41ىk���C�P��;^N��j$���oڶ����?V�Y� �d�����'���/�t.=û4�$U��"=�0�*�yT�'0HM]c(�������6(H$[߷�%B���x���%�'��w��]|���bT_�o]PGf�1�������6�0�!YMB�����z�I��(�R��<�D��gډ�S�Jii��[/D�o�I_��;�[h#�E��#ё��|)(���%7D_6a gNi�u>�8�9�i�r1�Z�1��*~^�b~��2�+%�٘�\�@V�)�",����d�
�y�#>���󊳷��� �*̞��ك�����7LUM��d0����Y��n�
��;�!��yU�u'��ؤɺV���̅�v�̞F��M���Ͳ����3\�q`�M�<�c������`Q���G��}cƴ㉕7Fb;gj�
8N�����<D�oa!��BkO��_]��B���QƇ����I2hDwl:��ieb�=�O�n�U�!{K[��)���W�҆l~�A��i4)�P�m��R�^*fbƄ5��`*�K���ǭ;aN�Y�-�b�bd��6��$}�Ը�4g �Js�$U��'l��_a%:v{�~"�������q�N<�@�i���Re�FɆ��Wg�'��D�4�
�����бG�#&`X�o�f�����{H�KO�`��eK�0m���&�7o{��3�qGȦB�E��?;�h�G�G"���&&p�bXA�ףL�G�BS�E$e��� 1�0�I���+H�e}�T0��U���N�.���J5�O|agJ�V�9�g��s�"�<��{:(l+� �76s���_�|޿s��/���{����\j�v
�%9V��P1�m�ڑ�Ɏ�q�IoK�\ѝ^g�@V0=k�!MN��s0u]�b�Q�	&��`lL&��W䴄چ0c?���b�ܣ������5���"\x-�Og��b�z���4�1VQh�xQXC�i��Z�T`�y���n�p�~��E�U�� ;�RR� :�̮�,���UJ,��܋8z�>m~P.��IV��Բ�
��xt�����;0�%�6OK����b�';�Rw��(S�`�C��H=ꂵ�q�d�:":��
���M"��<4��se�de�Ʃ�6�3xe}]�@��rv�Z{���aD��(��Ɏ̡��L��.}/�Ō�ރ>�����+Tx����N�ʆ �X��G�zf؟w쇛�7�yGA�<c>�G.����媖��!KNR���6����Nܓ�5֏A��^�,�/�
?��]R�2K��c��.	\�JFn���Np�f��3Q������v��%���8O}+	�#���\�Q�e|V!n���'ƻ�:(V��T���G�i��s�n��i��!C~��1�b�1Q����2�+C�m���U�굹o�wAD&?P1��w2��%�b5~���C�&@=�S��5���ų�/.ЮAt��q��Kڲd���K��	8�`;ˬ�o���-���X��ɬp��ᭁ]W�k��1p#�..���YMg��a�jwx#��)[������ĬZ�h�"����1����|�Qq�L�J5U',B���Z�:�(��%�4͂;��ka#�T)Y
�+12g�Q�C��w�+�<Je7��N�%y�~�V�g�q?\;F�p󨮷T� ә3�'�ώ�έ��l�wä؋�v f3����Ф�G�ΨH`�A���*w���IO�m�[�D��ܑ~���m����f�u��+� ��9j�`�+6݂(�+���+�j���#��2���o��^�r1T���[Ar���Ɵ�o�Nz��Pǚiaf���]�����N������,�kA���S����H��������gO��	�vO�AL�K��I�"�I��MHJT��3U|3��"n� ��w�;˨���I����Q�p�q�_�'��G8�Vy��r0N���&;�3��/L�@���\
A�ǼLS��8���d��Sj��;�
��w��	ܺW����f�@{)f]�A~!��&��FDb��(=���Y��d��ţ!"�w���a
��;w֩�-��Ŧ9q��74�G�����2�頮R�=q��v3���6�8���멎j�Ysʝ>��6���}	2�y�޵I?�$M�$ԫl�y$\��JP�:������~��V:�KI>0�>�\AUL�Lj2��y�C��Iw5�L�������0̾~��i���,/>Vԇ1�-Sй������Z%(�|(��b|G��T�Z��Ű|ko�
~��
u�������7+&���N*+q��*�$mC�AX��Ii9�`Ci��
���ݸ$-_°{"���C�f␈�Mټ�py�L/�D&����3%�6��e�hO��׍K�	�`M���'8*n|��F���w� �`P�j���hU�|�8�?��u���̑�л�F�v�8�+Pؾh�ܙ��sb�"Ke�	繅���<����gvI���f^�l����wX�iZ�m���
�N�;լ �ð �ʑ�X��e ��w�B�$C%ԕQ�i���%���*�`&*��.�&�sc�4��tC�"u���jL�y