��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�\W� u(�=@=ͺ��*"%S<E�E��r�YY�HPb
�^����S��E�P������ᓶ������W�d��%L��E]���g��'=�}ޢgP���x�w\n
�9IR��z�o�O*��V�V����'[�+�}�=j߮�01l�(��
�#��Ī�˺f���H]���;ۿ_�,	�	���N���Ӏ1����$7D��;�~F0��n�AH��  [�⦇��
;g��F�Z���Xs��K�yٞ���P�� ;`� �3z��8y�[������/s���#V_��~��1֩��1���FD�8.B�I���sH3��X���j�a�ߓ�+$<Ug�r��I M�xS�����!C�yr�B^���v/��#����'w��H^#�.%�i���Yi@y�|t�����{�� ^٪��R���a��2�O
,���۱�G���z����]L��M:��s��2���NT��t�h\�F�!����%T�_�C�k>@m�Ԩ(�5d�{2Q���̃]ꟻ�D��h{4B�P�U�%bߝ������
��Hќ�<�}�հ�mq��fᗲ2K�\f�s�bO�cl$����p�GO���:KV�S�3��)�hp�����ɒ�4�f��U�פ0��C�P\����4���B�p<�L��� �I+W���ydm��w����U�$s�>���쬨w�d�����ܞ�B��?�$���ʝ���f���������<5K����d��\�&]:�t���K����f˅i�zƐ��޽�N�+9�+r�?s�מ����o/��dpgԀi�C�`';|@��C)�d��6�ޞ�E��}��߸{I-E����7ۙ�L��ၼat2�;��jj�j�7�k�R�N=j�'��pn�dY�A�c�-���I��i��T	~��-�s[/^Z5�=��A�o�Sٺ�h�C�~�aP��KD�y5ܼ�޺2Se��9L����+8��4�+'����n9�{~9B���y,����c1�ֆ�C�t����]Z����j*������(H��S�M6ժDH�}��na]$d4�\���`S��s�8��c%<������������몞|���9�#�k$(�؞�i���]�$%b7l�c3ѫ�И����c���d耕V�6�/���V��Bm�?kѡ%&�;�s,����;沩��/�9�$R}޻#�3��q^7�;�+�UA�Jq�Z]::p#�����N��BB��HA0��AGm�,��1�f_"�����;���`��D͈m�gY ;Hڞ�	qm�r������J��$�*�})�ɣ���uF��|�qJ�6�#�w�I�=��:jd1��e 2����}�ƝS��3*ҎQ�g��}C��L|ٺQ,�o�Sr(��F��t�M�6�¶Qӯ���my�ʤV��;������B������fQ@���
���{:K4�q�{����4W���n��d������R{���66���7�%Z5���������6�3�������o���n]�ft�j�8�e�������&�cd��Q�t�ѷ�Y���x�h� WX��X�r��?��xG�ܢJG�/�s窱ww@�G%�� D3ŢB:h��I����N����q� #9�,���H(p���W^f��*ShC���	���@�)���	f�8!��	�4��Z��5���������(1�=ӟ|����;��d�x�����k�0Ϝ;��3���]U*7iK+r��Y5i���T��X#����B�/$)'��DɁ�;���U{��N	��T�}a-�����o��b�X����Ǿ��5�C��zf���'������]Ԭrz^��������ݖ5���A�g��	-�3%�hm�2���G�{s� ��83U\�i��O�n�΄��9d����J� � :cE�����5��_.��y��j=����f�A��
j>O���/��$�������tiEa�[�H�-2A��ĵ\aEb���0Sz��TTQ��%O%���*b�^<)풍��ŦwA�J'3�@���B35�A	�IVѩ6_������p�f�Ry�yם8�fD�L���W�;UM�(��b�~�l�g���>�6}�r�Z��W�Z�:$���=|~lMY���L�k=>V�n�����V����I��v�6#K��[ϭa�~����>��� X\�N~���?���`w;=W�.o./hi�(Nm`%��]u2ᅪVĪ{K�k�s���w�"R�!�?�@�п���;0��A���25�R��N��H17��;�;�R���~�W�:�3�V6�M"l������"��m	wwV�ϛ*B��@]�zh�zμ�6����[�3K����dw؄���K�׼Is|���?�%ޖ�ζ��/�����W��O8�d[����4�X9�)�0�H�y�M�V�[�Z�`�$d a����r�o�<�����zy�0 �b���T&6��ҽ��� ��w`q,E�&O��w��@���o�ҘN;�U/�(S�U�{B|4s�@��L�/�����M�O8�;��F��_��Y%�	(����S8��s&�}��2|8�8u~4����X����2;q:�ڂL
���>;o�)N���!��:��^��n}0��tjn}��O_�a��1�o�T��>�"N� t�y�t@�H(���A��&y��:���߇����E�����9g2TJmf�71�$���X��=�NL����&8 '��x9Uy��h 3�ͣp����u �g�x�D�W�UR�Y~�7 ~F0��Rc��J�^�?��q?����:��4�'����qm���K�BK(�N�fA�(*�&d+E�r�n8�^ElSC^$�J�q�V��?����Z�s�CѺZ7��_B�3{��ч��;dz��A�`���!�d�V�Y�4��@Q;(���^��h��!�i#ϪB�S� �Y�D�Ů��-���T���j�K��U(�,m_�8V�{_�����u�8n�3��4�+�[�9Ȃ �.�*.~�z�6����5� O5�]oͤv��H:@$1����Gh���N��8����W�r�9Щ����8�F�k�U�����~S3g4�ˆʮ�k�^�fDҺ� g�||u�I��A�HEz����%*mV��I�'�oTQ�Ӑv��$�]���Լ��;qᆁf6��'����t߳DS�U�	������0 �0��ü�T�����DG_9�I^L������̯��hP��Td�j��
]�V߅���¼�\��Q56T�QN⒭�Hi���_�|�A�����!�Α�4C�]���)�*��X����(\Yzz�a�'.��wA��hwAH�W9So�@��4�UqLnd9���{ŨB ��j��kbU�I�%ޙF �O�_��%BD~��C{,z��[d�2z?=�3|�f�K:�%���Zz7�h�`-�\�3�o=cT�����X��u�8l8e���N3T !���Gc�0��u�0
����X�&������Ecb'Z]�����f����(=�����C���Ec��xE{w@l����N#ȧ�7<�M�`�}�u�ǝdl�H���䣺=�kȑ��ۓ�ҫ�g)`�eH��O���)�6��n :d�ě��^����Q�Mr�W8~�X+���˲���|$�5%����z���A�m�]ң��V���L��<�g�����]_Fbusm���\Л���a
O�����iǾ�k:�0���8��w���k���K�a2Z����02�C
}tN�5��H_N�!	�C0k)9�Ԧ��SJ:���ܯ=�^d"�BG�V	��^ʘ��J�t�'* �3fDw��N��L%�F}��Ӷ��&�j�T (QR��UF�0&�m�k-�t�"!�����)"�<��I��~|�`
��:zk�iKzA����h $N�0 ��,\
�^�4����Y���x|��ގ&��|Y���ȁ�WN7�{�
�#t՜/���[�VY�i�*$=�}ka�!
�,	����O������Etqd�jՂ�;J��.w������R=���Gu�#g���x�{+�Q*���>��EwGJA4a3_1~wȠc����&vM���#�<H�f�Khƀ
e4=J�X�Y�|��Ӟ��Ϥ����P"B�0-D��Ȳ�/7f�7�}'FxRO���� ���nW�P�Q�yΪLA���I���=���ۊ��oֵ�Ah2�hP�._��&@��We?,0���d9�zpK�C6�hߛN6j�uzTQ!��J������������G���bn��n~��F� \ �ɫܸIi�����k�����{�S�	���~f��B��g�8v��;a=�@�|��Ac��������7=���M0��zBoR{����"��A��kr����=Z(���j��>����!%�I���h5Y��}��b�6,��|?�&�j�/%�Ca�3,�t��rМcv�4����� y|�8%��^C�f��?�Ik�t���@�G:4I����"�j���p���;a�j����.�Z�H;}6�f��9ra'^�I
��[��m�npB���#�b��Qr�($��
�@:�pdq����p��[�J�Nf����(ݮ���
�	��C�5�}ꋲKɷɉ�������Ј�~����u����|K�aPX�`�놨�U%�?�O�׾�y��ב�Nu�\�+�V�9��*ڽ꡶�]����Jڦ��\�0���F�K���,��{@Qj� �K4�J��(��"_*!)(��7<j]�o��`bB���"�r?L�D�Y�,��D�}Ψ��:����y(�P��$�<�pm9XH�I���ƻE�6�2���ץ}�4�I߯��J��%���t�?�л<K����S��R����#F��� �S7�������'�f�������I6?S�;�a{ջgJ:���뷕�"b�]q�G�]����!���T�,����[�Ii���]�W�l�����ӗL(��l�A��G>�ʔ�>���!g���I�SckT1�?�s�����v(���Qq�M͹d%��[�[*�ľ��"�'��z�n'�%����%��`�=í�=�OWz2����` ��[r�?�[<+�4u
N�Yy���3��d�B�>�-��=��h�6\o��
�k����Uw��
Xz�?�ÙBW��1�}��E�9�i�<��=���9~�Ky�`A��p�z��,��m������2�i����6�1����������"ֻ���n)���*�1�d^�8d�]������{�%����btչ�@�	OF����V�q��ۍ�dW�����@p�֣����<��1 �����aZ6�G�������	Ǫ�_���Țw �E+f�����Y�0�$^�}�h��Mp�6��XQne-tF*����P����է;);�俩|t�����:���VACE���M�1U���w*�X��Kc+r28n$��1+��"$۬gu�חs�~������d��g%c�1�{�"p��ç���׾�E~��lN�2[/�^Y�B[":h�?�k��6!�!�P�T��f!"��$���ap"���~k�d8j��LW���L �>�?7��@*3W��O�xj`\�ac!m��E(�R#Ƿ����H�|:ru��������~ GC/3��V�u�P���x��CL�7��E%��r� 0�X�vi���MĴ�L�/��ޙvd���X��zD0b�ɑ���π���ex�Q��!��`j��e��S:|F>�>�ߚzaSބtIԵR�n�ye��_|y�.���:zn�
�+�#��fP�eD�u����-����ph*]���~��oo��0N�F�a!��#}~2@�� �v6ܦ0@��бJ�L5�k�
H�H��y�n�c#�B�P٥��rVY�t�'�O�ٮ%�����>���L��L�4�`# �}X�x�'�&/�-��kۭ���DMo1�����p!�అ����̯4.N��(r1(N� Fl����8Y�<:��wXs#O1o����<�!!s9����M�,���x�%���M�x�⹝݆��]���>s8���Ě��>�tDQ�/X0�HdU%$��.DH!�r:0�U�Qw��Ff�Qf���|�x|b�M�ߓP��sr�a�S�M�"B��{�cX;�p��{�a�w��MlŢ���oC�ך�<���BdU.E�$�E:��"1���\$˶���+T�)	,L-�K�+�+2��ùO<犬�����|]{�\x��O�;�/�7^gLz��lJ=�?�vx�e򘺋L����G�m�T�>D�-�$r�T�3�t��Ь�#������TS�z�d��!S���j�ҳx����R�}2�ޛ�m�:Ñδ���ݑ�I�����P�5�#��P�0 W��We��LZ3�Z4E��Gy]�bƾt#��:�-�P��]ܰ��VKԪ���k%�}�e����n@r6@6cn�?h{�۴��v2u~���	oas����G@���-%%ˬ��~[9�,Ve�o}��c��d�o������"���P��%0��I����[�Z��F= W��io��ȃEYr������JuH��[)���>U't�%����67�X؏��5��"�ly2�{���;g��)���&����A�-�@���a�&~�a�S�.У�r���&�bx���9g�ɨ�(�r���ʅ�h�n��IUe�Ϟ�c��9�c�����.?D2V
h6����'�fz3�y����-�X�*
�#iU���~�lZ�~|f�+�(�M�(�@���p��9��-�(Q�
���h���W���1%/_PIY)�N����@ ��ap�ĝ��FÑh2�1ІӤZdz������6��{�4��H���|5����X��uƝ��U�����.XO�����Ň_����ռ��q.D쓰��Hہc�I�P$��n	c�{"�Q��4���������A�U�?���q-re	�K��޸�����Ss1^�b�V�j�����\��ڠbB��B���l�*:N��o����WX>��ß	���qC��d$=�p��6)��H9!i�����Ҧ�m;7��7����͛ˣؠ}�B��`��QK{.X�J�Qc�$k��Z����@}c$�b�F�v�>숤��Nk�n80�Te+�b|����E��$@��h��˔���e��<��Q����a	��@����F��p����^I������["}�����d��~�,�=4<�F�F�ҥ;wav�%�|K5O۲�Eݒ��N+���I�Q�ajo��Bz���r@�W�����7�������	�o�)�p�h�u��	�����O���t3P^�[?�0!$�� r�{&�_�W�?�SP/��g���nŇ�Xx-�d�+�;27b�$>��e{|Ҥ�rMC]�q��  <���	��#h�%���z��IA�� ����2���#���b+!����M���d�
�%�Z������Y�v�N���ڸ Ё���B��:�v���\��\�e��IתH�]��>6)�߱q�"W�`�	^��{V����[��`��Ȫ�1���0NM�V�r�눊��e�a'	��FfɎ���������SQ[Ou"��ܒ���K�4|nY��I�1L�E�W/���Y�z�&���}���)H�M�!���������/Z����C`�آu�����h5�mzzlf~�p�+BifO4�n?��>����s(Jh��Ɓ"�E��?f9Si�['@�ub%��G�Obf�����&؛'�J���p�<��k=���ܸ���_�<�)
��I5�K� �X�n'����oV�P[��A��)~#�p!"E�Лm��w�n�B�6 "���J��#C��V8����v0$=].�/�5ۯ�??!����
`�?�B^���XYe�P�!�J�̢\h��ʬm;�InA�+ɛ�}D���g�S���q^Sۥ��]J��f�gu����2�@:c��s�Un���-��q�+�~��o�M	�ƠVe�٤}���R�	���Y����{i&mP��b`-���hתe=��H�^�^�J�v<	�$~:t�=���8�5� �F&��V�_^FK�ּ�D���=TPx�ԕ�=�%�gY�9c�A=cH��S��ଳ6��x,o/�ō"���ˢ�j�M���d:Jؼ���=B�ه�-�Crj�(��|��m����Q�l�j\N,���;5���'��HC �-+v���T8�G�#���Ǵ|���Sa�x�t�ͬNm���p]���a��dB�9]�;4����$cQ}�L���$�d��p냁W�K��������$r�A��V&9���U��z�ϧ?@td�ĥ�zE��t\w��Y��m4^i�hɄf(	i{ݖ�5l\�m�fʭ�{�h �F� xD�)�B�͟d�	��A���nӣ8���ma�(���⪏���X��C���N�*<V/�����+[��̘��n���\�+Yhv�3z[��i �`�Ã2��'��/t�U+���:�V�&�r(�WZ,�" �+5X��P���z�>H"<�sң�V�"�
��+ԩ��~��c�M�B�Da�p62tE"�x���NhtOU+d9R�!U�0��*f��9A ������t��%V9�W�0k"fS�%R�f��ǣ _��I���A�v�=�*�l���֩e&F��@�wɈM���M�����v��]zQ���F�����V�vzSS�}���"���A�U=v���&\�2��}�L]U8���k��ȟr�]� A���*#�h.�#�D�e��?������w+O��U��$k�C�褈�d�>�ŷV��qz�@�O�/����T�@#�Z���=���"����A�B�C�E2D��5���tj�����9�����u^�!$Z�x��[���}L@�OFw#�'��S��z�����
����d6�}�a]�eLi�a)5d^ů
��$� 0��Ra�AKv%�Rn�;`�wb�+�ku��X2�>K3v��|?�f>x���;��4�Ĝ��{ѭ�6��i���d�~�tK��|��;�
v�Zp@h�'�����p��	ȚcZ\�����m��(�[���.���͆��媔i��`��%�0��t�(|:]��lSj�TЮ�5��26]��\˕����!�@_�r�榭e%��I.��,JS���������Qc������}�V.�-�) ��d$R�u��s+;�����r0�{�Q�J�y���x�|dW��y�~Plp	�r�nUa3��x�x�y�|�n��W�4( +���-��6�(#�-�܌��=|5�6������!h[�;;����
���0�CM�Y�����5_�����C�I�0�)��Iּt3�Ӑ�\���F Y��8U�\�Zf ��g&m*3ȕ��t�ftC�~�/���`\��ml�R�w@m2�SV3.��倧�J�{���<$�EIF1�ٱ�;���]�
Q��ő,Z+������xK����ʈ�~.[dT,
����A�(�'B�W�t
��g��wo��/��'��^0|���QO�zq�R� ��X"��\U�<� oת�\�IҮO($��u��X�I�_��q:�H�$dC�Ї"R�#4��(�Bؠ�*o��8lW��q�,��+�X���4Nq�I�B�ՏPÅ�����Ӆ:�wt��&]�B�j���R)˫S]0/�b�EC�9�M+jp
�K=�9�W.X!��ذ�����V9�?3r��u 4,����#Ʌk�ߥ+�u@l�:�]VU����׷��ܫ��_K�[��v7���P}]���}�!���*d^�39����-1�V��.�\���]p�O_�9��@�T��+vƖ/g�L�"�L�Rc�0Е�͘�P���%󼯽G�U�Es�'�@kCa;��`hH���ɦ�
���sV�r1>�����b/g�Ἲ�;M�3=Z����Yg�m�L�ۻlo�7���7y�F�$��z�����5���\��v2�I�I7���槇0��>�����W@�]*�Jڭ�6�uv��E*�`�I̙^����z��j�8H������G�L�ٜ��ct��b��߶������z6<H18��ż��#�u�4�s�[Z�,	�1l�n<>N�}�P���C���ؤ��.|�`�۸<ן{�"A:K�Z�E30T���.9�(�5�5�[ ^�{��^���b��������	O�)�{��~+�#%��MF��k#�� 1��0D��h�j,i��qm��e]q��v�����1����hR�!$�~�G{{AG��<���F�b���>#��\��0�c�̍5��o����{���ƻ��
�Y�>5��iˎ�����V]~O� �oo�l�4IT>Q�7e�u���o�v-_D5t�)t�����#���vQ������� �Ll��,����q$�K6/!���TΦ-�KW0���[���K���|kLS8���Cd��Y�[`�w/+pu����`���p��jϷ����l؀����R�jB��ݰ?S�=R�4GE�T���*��;FT�@���y���w�detM*E��V�L�|�W���#���$�����,Q+�/�S3u���k��x`E�k>2Rp�8o�������}� �7����+o�0�)��?�9L�BWTB>?��:黆	�zmɛh�/�a���iۃ�^D�|�Td�I��*�P��k�L.9�qϴAI�F����蘵\�O�����e�c��U,^�fv�gb�k�~�[$���M&�?3U��ш��&���z�u�y���2��I�^�����&��D���qƆ�
=��%D���$Vf\9-�Q��t?/\M}_=�km�ג���%��9�HEm^D-W�%�
.w䞀Na�������:FH��
�B���O�~���u��#����x�(��\�����+�,~8�3�jˣ��~������$i��ײw��H����ϵ�h@�=zl�Y�[-�Mj����2z7��4d�W�Ғ���̪�� ���L�jaW��`7�7��!��EwV�p���!!���}6k+0��XK����&K·9\��X��Hi�.�J�_�ƒN(�"�!�]�����V�̆�A `�y��I�pn'�A�Wa6��������L=�8�ȹ��8��\:�
 a_���D���eKT]�)kwo
|�������Y�F��L@mA�F��Rی�5�=�I�v,{��cM��q��"K��#���:�>bA���lX�8���ً��e������D��&j�@��2B����i����E��+���P��<\Q��h7�%,C������;ҝ�э����a��Y�5�jia�G���l)
�������(pH�+W"�~�V*1�?�	����6f5D+Y>�3��zsI���s��;k�`�����Z�@����j���}U�~i<�����]�;��2 ��1���( �qJ2Q*F�a�U���\g�P7�}����bT ַ��=������k�]Kz:�]{��,�A��h�Z��Ѷ{Em];�n;��C�YDQ��6�lh�@��딺A�%���\�B)7����g?�2���y���N�ޒʠ�G�r2n���s�k5��zּ�ٙ&��2�&"I�L����J��؁�/>�b�Јk��l�5��m����ޖIY|b����7��[��:�T#��e�*$\�e�j)��O���"ĳMb�]���x���/����U����I�=�#^v���!�E{5-g4�鹲�KR�F���Kb�.Kٲr�R9��h�'ޙf(��Y�H�e�����W�Օ�ud:R�zl�3��P� {|�>G�4x�<4��b.���Ar��#�����+Xt��!�3�^@�L�;�oU�\ ��JK�$��͇�G٣n �%-��O׳����{K��x�o�xl���+7�� �X�t6�}��X�H{�	����-��н7��q���2�"�=��՗�V¯�X���NP�ybe���􈛱�9l�}]��c�@uLi�p�B�v�9��`x�ƛP���"�c�)�a(�Oۻ�=������H.u�y5}9��>�ZJ]�C:��æ�aE�H����aq�НOQ�7������"D(#X�^ږ�X���A?B�#�̢u���`����r��U��B(��i�c�yꥰY�P��G'��4\�(J?>�X���wI���J�#$p�vi����O1k���N���hC�rh	����TNHY�α:;]v�nJ3��G���ȫ���0�S D��!�)�o5�^d1�X�Gt[tD~�"��换������L�*�L��|���|�,X%|BѧK1|���'r��d^\Rs�0�ٚ-6�b.��x���
YY���T�:�s�������k�0
�́��;�N����������be�����	'XJ���=��!�{NZ&���UMSY
�j��~f>��7�����J|Z9���h��.�=�V=�֘_A���jbp�g�� �j���aL��Y��1���8+͘��U̴�9���3ɐT�u�z�u֒���1�����+ui��ZZqZ��b]:V	���n�Y��,���8�?��za�v ����8g��xYm�Ą�rB�;���A��B��D�Z�p�&����cV�l?�t�Wpꡛ�%n@Cm�v�j�����y��*|#���P�����	5�0�[v�nl0�����AMdG�7��� ܞ�\5˅A#�Ԁ�ʐ�W��e@��-:E�"D�DT�!<C��둋�d�=�-)~��sQL�K�+l�`��뛪gѯ�D�(?�K�1:�h �5a��}'t�`�w
5�Lh-%|wwF��(q�I���Z �Wa�p�(P�84`�L�h<�R	o����Z��j`)y3�M�5>|��l���� Q�xM�xw��s�<)����q���q)��cϽF�E�?�]�@1��5��Wڀ-9O[F]�PӞ�;��}�;�YI_��+ZX��QŠ�+�u��=v
�Kz[�S���w�@<�Io)���6p��}|� �j~6��U��\*��	�5t����Rw[0x���B"I& ,3��{C�$��H�Ɂ$�,I�fa��ˎHk�#�>�=��կ���<�qg�qG ッ�H��e�ـ��w���d��0ԸB�e�B�>q�� �,sf���d�)z<��I��a�W�$z̋��
������#�0$�_�z��/i�A��|]L�{�����Q�N�b�"��ӱ&*>K���!g���
3̔U�?Nu-4 l�u��V��:�C�E�2i@C^����שћ����0�� '�ڲfw��~�����/L�7xA�����*�� P C�>�_�m&j"�T_t�՛�y��L�S�)C��<�?�j�Gp�zj�,O^��`be���y!��-X��yf[��F��c����c���۾�J�=������㕏�8J��i3R�_e�]e��E*n����.��/������ۃ������#�ZYU/>^YC	���{��e��ݝn�w�c�w�������ʽ�/a[�����?4�����7�4�C���c�1�P�/�X�����`��
�)p�=b0�2č�f�g��z�}�S�Wy�*8��%�NS����I�T�t��p�pf�FU5���{��Dܪ:rJ'�M?��KC���@e�f����w����N#"�5P��5u�/�to06p	������k�:��z��*��V��=�GMA$kZ)M~M�8U+x�ǰR�����y�N���*䴚$k�C��0�VN
2.2����gt���wS~y���ŨO��pt/�K�Ne@y�������!R�I/��*�Z<�[wH0'�K��M>�]-�cʙ|�:5��L��(�,<�����=,���G��/*�������?	ʜ}S���Ş��|���+�3z~��>��~@�HD�j��4#��IfT�V.5�����%�*3eJ���Z��I�wg� 
K@!t��<�������u�+��a�SD�ǐ9��;@�9}g8Jͺ"��xWJ?.A�eK��1��J%�3�tT����Z���v,��>�1C�Uv�t2iMUL����7
� 9�E*Ñ�����l��@�?��Aw@)�=�R¥0�����B��]r(Au7��#��,\5�5�[m���(�PȾW�x�	Q+Ň ���&��D^�Q#�V�%ql�/]:b��9O1��Ύ�jY5o7�~�&��� ��t�T��l���h��ݒ�|��G�g�"�����c�24�c��R�3�w��U��du���<��W�D��N�n�c�-l��|�5�����=	�b�2��M�� k@���4��g����[�p"bT������XX�ؐ�� �WN��U��@_iq�n���§�����v���1z?�b��q#�%G�������-�Y�D��'�r���@��x]�q=���1����>=��
Q��O�G�����d��E����]��F�l���N3m�T��U�Bc���R�4W�X��\�ԫT>��Ď���x@*��E�Nذ(����8���sĳ�U0>lUZ��$�%,�:�&)R�>O�*�@���?ev� ��!E��Yt_8����Ҟ8�#Jn[Bj�K�����w��M3�BCzAվo��jGy(�k%W��E���T�YE<ɻ��,s���O�)����͐P�+	[-���ğ�'��P謦��� �R罰�dr(]� �#��>SI����5`ZCr��D�}v��p�5��s�	�|�>�H���~�uQk��e(o+ϴ:������+�*��߸}L�)f�8%�9��a�1l���R���i_�����z;'4M�ש�יG4��6ƛL'�����1Q�73"��k���%ٮ��y�gA�����0�>2�r5[��,��0���O���BꙜ�E�T\#_7+h^���7���F*�,z|�t�[;u��
f�l,^�`5ϩB����]��_�x���c10T�jQ��k�c��׏����I-��l�9M��Њ�.�k��fv�"����+7-�fz���vS*���v�����M�-?��8�0���V������֝\�~J��9?�DicT]��`VԌޟS"�����X7��)�L�>n>E8��s^�}A��܌�ʶ8�`;�.eu,2�����]p%�U��Dz#ɠjmPF�?��E�XZJL;ˮo�zGL�$���-�?<(|�T�%L����6D��A�v�"-�����E�l�I `x���e�dK@��`�?a��t�&�ŞF��ݞ��{���y����D�2^u���q������ПŬE�^{�