��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)���-5��T)�uYl���hP�LZOn�n�H��l%��/N�*'��@��t�<����'�B��L^�U�:�,�%��&xc�'�}�xk�s.?P�|�JG����b "g�e��-�I�3B!="��,]33ZM̽i����.|+��cêJ��d��B��|�-G�����y�>?����0�2ܕ�mm�O7�l���V&����s8��z[P%j��99wg���mV��)����z���8��~|�3�K��\�z, J��o��[�$m(U��%���S/	�^9���Q��G���X��Vk8��	c`ς�Ņ�p�-)Y��a�[�^�Ӎ���Ƴ|�"e�,�d@.�VD]�a��u��~X�ǥf%�)V�Ƅm��	�wU��P��PZ��a'�4������ ��c
��n�|X��ɢ�$&�x5�raP D�rn���G�qPz\i�VLXw�Q�}�(�}7	
���f���g`l2�����d�� Bw�4bܶ����Έ�/��QۗR�(h�X�Op�Ѧjɂ�_*�ݭ�D��~5<��&km�����{ 勂A`�O����/pB�	{�J�۵-�kt��K��b��u�F.b�.�����Ys�Y+��1�H��9@3뤫��g��C?��/���H*���w�����*��Ġ��bw�Eͬ{N
I%�w{r�����x����Jd{�CJ����Y(�L9_�6:Ϭ'�AؽĬ� MRU��zm�E#!�Hk{ڮ�Vl:<���ń�z�Co���J�S�
=l�K�G���y�kߧ��s�L_5rQ��Τ=��<U{�T����PT�-�6�L�3�a�|�s�Fy�>�kU+O����,���s�6/��R�!�Y�p{��� .A� � i
"v�Ŕ�� �T�vNIQ��հ��s�Ɂ�LyW���ky�U��ˣb�'`�h36IU�~"�_J"$���Ӆ���ݹ3�t�%�,�AN�<�`Zؤx�C���z��㞕��
@��4�2��՗��x8�%��?�t�[$�ly>H�Pҷ�qf�R�̝�8�E1�i�ו'����Jw=9IZ_vb:ja��x�㆟��="�"����Z�9�T�{���Rw�K䲮j���(l�xY��F�ݧ|�Y�2������"�r�fSd���M�7��U�����|_�u��'�Gu�p8�~oRX�����o��Ȅ>s�%�B�1ܥk=��΋#�Oō3J����^d{��Z�Va�۠�׻��S*�y�!�p��HW]4��o�Q��
�B�J���Y�ch,#��vS��ޙ�I}{�Ht���#&���|�
皢T�Br�d/��"e�v.��6GM/�);���~��$��p�{�\'KQ�:�dgD�����/q�ߔNm��������j�<%Hs�U� ��G�r�#|�c&7s�qz���6�X�1�V:<�g����JOp}{�0[WJ��'E��2��� E۹������(��h�D�b�،�d�81:WpO`����Q���^�s8���
�SK���d���B��������gt`nG���sI��3�2r��]�a{���'��-{zg���.*Yml�FW��sr�v�Lf.M��^&/`V�H��1��"q�qe#Z�u�K����Z];���+�wėz��8f�'�JC!6p��Ԙ�,�H�s'�"DIv�2�b1���3�x�,��ZP��ީ�H�!S��`�F�ټ=��{�a�c$�}�6AS�R1m `H�'� z��M��0����ۼ��=H�C�LH�@φ�����a״_�_��LWkJpܣA��[/Yt�_��2�BJ��TW/�`~�g��p1YBHõ����rGq��T�!�^�Xk��%"�w�	��
�_pG.F��x9�!A��V4}@ٱ�G�F�E��<ϼή�6��7�T���R��x<E�mc��4��e��U:{��r������6��>$���,Ƴls���ʻ��⠬�Ғ�6t�5]����?�%�n�X-m."$��C���}`��(V˃�h�,S���OW�C��HQ��%٤�D}?	���_.P=�G*�(���bUE.����
�٭`�"����ĵ_l�J�G�(`ilby�!/yQLq&���X��}�� 	��r�x�	�D���X�`��.o&�D�Po"��#��=N^y)���}�������r���:_1(V�lK�w�դ�5���=�Q+:���� �'"_��MH��3^+I���LsY���)V�;��R�U�AU�" �5,37�M�R,T.,���1�R�7������d'�B�I�3�r�@����FUQ�A�w;�s��G�Wq�����T��ЏL�tP�2N�����[9	/_��vT~˚�l�����l�5�O�dBd�oo��d�'z6�q|��L�����	(J&Fݵ_��vrY��Oͫ���ڄ:~rL�g�8��Z��ǡ[�C�[À����ll3]/"��s%3�}����4��qW�욻���,7=c�1Yr��gօQ.�rU#�5)p:jD��%�f�e�&&���&�`��`�� �3[ t^�ɡBKի�MX".H�Hyi[_ni�����#����)�jݽ��r� �Mug}ONl�9"y�ίU��r����u�]t[����F���khӇ�(Bʋu�(�W*;�����A��JM{�p�{DL��1eŹ3��cǢs�ԩ�����O~�^�҈s{���[,�f�W���G���M���������(������~��.��W���7S?϶���]��o�������z�:�m��+d���7�+��-p���{T`�� ^#b�^;�S��O�Z-M�����J��/ )��u�[��+�s��\d	����"�܃���Հ�������h^�[4^n7�K�v7��+9�ߩ��'l"�x�k�Z1_X;�8=�.pm=^ ـ��!�抁6\YHn�>!-m��#�x�a����u���EE���,�r
u�F;N�lH��"c����{Z�uk��d��K��GK�:���e?:C�� �����^y2�(�����J?aH��K����+�֥͂�r���T_k�S���7��%g�^7Jv�Z��b��x� em��ƃ{�b��v���5�'.j��7�����?4$�|HkD:�ʐ�;�l!6�J��-�-�DKnVZ}��HP�Q�B{2�-���-4��>����N�/{��=��?��8�+I*˻B��lG�o]�ugֿ��Ƽ��]f��k�r������C������;�H�0Q��/��`��@��WF�~�4���V_u�JCԯ:�������g۳udͷL&'c��u7t�0��F�Z4��Xw���H�C&9SV`�>]K�ٌa��U�|l���e����*�gv͆c�;{���0n-w��D�o4C�to6)Ŏ�Qq[	Zq�cF�J�B�Z����d���F�M��Ώj�R�w�%Ct�2�l�Q1�2x��o���f�B\c���t�8�xE�����[��k��V&I����q�;
�����[|*&V��  J��9C�|$��[��~�r��^�ME/>��2����}
C�(U9S���uKI˭2o��ѬY��<l��G�b4;������c�0�Q>�Pe~��6��(G�;��#n���	 ������΁�:VY�u�&y�tҰ��]���l��a��A�Kp�e)� �4{�����$c�/�vT��7ƿ�i+��G��p�b���
�6�������N 2��DC�!���OFG�-����o,'	vGz6��*q�ߐə�Hӭ�vnIoCO7�"4�r�q�����i�Hٴ��P3�'v���D�8�������nNdy�I��O��3��՛$1�m쫪uʼO�eM��Y�2piHp`]D�����@g/-�"��-���r�Y_G_�S��nmZ�j��rX�9�[��"�q��'/�$���3�F�����/k�Km�&���k�VW�1ZV/y�T�1��j�-Ԁg��ۻIx�O ��Cd���Q43R�RN4y��2��ic�.� �4!�5,`,5��S��qd��ހ��V0��x�!�K}�nHʮ~�7h�SL�KW����I�<���s>]~�O�`�5IB�,�<��?��o�#]s�#��N����-Cx���;C���[ﯳ�l-F(�\����C��"o��^�t(��Ĕb\#���Xl ���Q���d}1$(<3����UoOa�f�����P	�v�wߢ%Y��9K�O������2�D
+����H�=�j�P��w���Ө~Z
����u�q*2���>�}�r7�����>�.If_�M����Ѯ��5	Z7�R)~/r�Ӟ��^f��J�>����韲*|�۟bi�LU^�J׮����ץӗ��A����ȥ� z��Dj��m2rXc)��p��=�zmi��}��Ե�gx�@?�WN%p�����t�h��l�ɷ�fNڃ2����ͭ���5�2v~����D�`�Sc��0�&�������\4���c3~_
�BZd���f}.0�k�o��	voc��mV����N�Q�<����#}�A܌|���e�k
L7k�{��Ȟ�Iϸ�g�5�D��]�4�Z�$l��Tk/��[��#�~{@qU �-���-��ocJ4S��U��R�Ɯ��BsQo*jO�.6�=�e8$>3�z�dR�Ҥ'�3*��R��1�zL��[�x�,�o�_�.�s&���%8��f)7��5��|�s�5�g��bA]0yAJ�*ۯ����eO���\�4�^G@C��u�;�o�m᥹E.�ttY��$���O�e0§A���b�$M�s�'�g"�n��K�GvҞ'���6��s��Wl1�,�8�S0����v��@�<��������Z�~���
Tj�}k�z��:�*k\F0�1�@�)�S��+�[CD<C|9�ԩ�ð��E�dж,�F���.O�N�G���\Q��f�{���1.F����d�h��8>�l�i6�x���8�c�|_�o������qo�U� oȮ�5����A��0J�ΐ���((�'��zi��t�ul�E�WV�����@}�����[�7or���ۘk����fK�א��D�B�{����H�x*�˫�:�f]%K$�͇�;�H���1#�u�w��2)���y�TQ�w�:�xٳȟ�2:Fw�ֹ$!��xϩ���y��$}T��[���������XX� G�#v�_B�w�g����e�$ �����o?i��=N�'�Uk;H��Yx�fC3������W�����3���s�!�=؁G@L�� �!T@�1��Z	��gx'�X �H:����0��g�&�/~�s������2��)���f9�M�қ�Eqw1��' 8��aen��/C\,
������hb_�f���O��d*��
Ä �����8�̎�7կk���-%��)�{��CCcba@���uf�Zr�GH���ks��o9A�/��(�*.�p/0�U��b��O׮�P��7"K�&�V�/_�W#J�G�j����7����ˡ��ʔ�ҥO����{�)��\�v���_��nLl=;_5�Y;�������ӑ�1^r/���D t���<�B��s�{y��kQ��Jpȵ"��&}��9H�*(T����Q�S�lrʈs����<��U:�ڵ��F��߲��̞�.e�1��&�P���L�� ��-��0��ÿ�%�ۜ�Q>!�(���S��R|?��1��hamYl0�O�C�+�k�m�ڃ�l%%��\4�V;�ٱ=�X�(���
5#�?^��LkRߏ�$�9=u����.��L�2�|m��t"�f/\��nY�ǻ�D�&�a�{@5��n�p�x������V�?�^tg~�x��M]a[;&�p�3e%��脚S,�$��r��
@�<R�}��ýB�G�QV'x�/g� �ᕎ�<�?z,�)�;l`�w^Û��jED%�5�t��
<u��_)<4���.�PB3\�e�K<&ݥM 3 ���Re`�"Q����: i!V�>p�\$�;�����F�FiP'� Q���Ԥ���n�C�K2)�[����5�c����f���~������7��h���Ѽ0��x����ɮ�[^,�ݢڮ�P��IF3�!�+����.������V��B� w<��h�N
/nm=���n��p;dZ�O_"�Ӻ|Zy���>!$���A�|QS]���}�aoi�����X�D�D\��z(2���/ q�����%�:�٢�"����Yy�`����l��^��2�\{:BD)-ٍe��\�����b��l�$��Ks�[�A���3(E����ٹ�{�Z���k��e��e�K��<� |� �e�l�lʌ���z�b��n�Q���r�����]���m�!doI�.[�f�˾����Ď�����MR��e�W��L~����V ��1�+g��x���(d����\!��4K�/�����7��/��m*���<���������@Ǆcj� f�̂%v���T�,y�!{FѲ<���2L���H��öGƣ�U�g���t!?ݵo����#O.V���E9sW�m ,WGum�gk!��}1�c���'�G�4���OΪɢ��̏�f������Qf�ৣ)�h}n�XD��>��6�K3+�x�)&��hk?Z��_���i�ŲdaF�pH��FNZ�5ym��q��]N3jE=��>ݑ;��آ4��{���@,~~�S�h���kf�:S�D�PP�6��O�S�Ċ9y�+�M؀���*;���#m�������s�9���P?j�������U��Ƭ�Vi}N�%^�bO���v,�}Ol�����mI��7���� �%V�_�`���T[:����c���7��u8���+Q�eg�@F�)�X�Ҝ�f�n��Z�5� ��
�|-��В��Qx���QR�1�;���G�+T@ҝ�`#=0�[��*$�6��(��ŭ��I��0^�wH�_�E��V�t�7���q�o�fh��G�L]\��b�T����.�
[�z��]^���UCȹ��E�� f
��D(�Mº�ӧ u��H�[S�q*�((K�_��u�W�1��."�¹��!���[f%�]!��ֶYK��.�@ܕ��"x�Ŝ��
۽����kG�1��=U�� ��^���)Ls�
T_��u�fqV$+D� �Bs ��H�@]U�YO�Gw�*t�3�㰖�~Џ�O>�_�r�������W�9>��So'Z�v�? 9�M�����K��A������[2c->_�
̞��	�ܱ�M�$��:��ݲs�;���63��z���q����0��nz]X��I��$+�=-Bl����qo`��[�$xd�B��-<�>�mƩ p�C���z�\E󪁤�F�S���7(�M�+l���+wJ�sYb��zĥ䱁"#1%6#u$��R,�9�!9H`+���%������86�k��o�7's=�ȋl�F�3 �$(?�%,n����	���2��H~�.�
�
���eA�i���JC�BMWw��fF�d�B��݄%�V�yJ���̨M�
�{�c�rq}2V�!b��$ƈ1ַU��?s�����i�5^�/���X���bX�N���mR�3���S�
Yc>L��WJ�~	c���F��\i
�6�R�İ�:�
�.��u�8���1^^������~����*��9ڄm��!���~�I
�p��%��K_���)�IO�{����BwA����U���?~��x��e^�@���6��c���NC��&�y��B��Q=T�)�+DJ^0�|SEE��\ueJ�@��0��ݏ]��TZ�w�H�)ZS����[��9��%%�,�!p!�td����:�QFnM�!�}�g\�a���ȎV�5��OjqZa�u�k;!px<�Z񈸬�D�������&�sOⶐ]�/���B?$�D��2����E���O�vOP���#�����q��{�pB�s����}��B��ڦv������4"��lTh���B�#������{G��9_��*��y��O��Ɂ
�Ց�0��KB���Ӛ��X����II9,���-���&�ǮmA�`.�胂�+A��s��Q|��
���L~��C�@bO�Y���,���Ȣ@�BV����Ex[��{z/ �=�H��!+���-�ǁ�u��ٟ�����e�C0�}�I�֌dVX.�ɗ�g�r�a��eZ3��f��Bb(�C��<R���U!��w�j�Blj�����N�� 01Q�}ؚ�����vN��q�*���tt���qw#j&THD5W:y�!qÒs�Љ�~����Ma�cP�d|`?���0ݻ�ΰ���oU��(Ԝw�d�B����r���?sp�͍D���;(՝z5j�5�@��b/��j�J��Y��V�a%KB���w�������z�=��ŗ.�ߣ���ڶ@;�5l��eo?͠��wG*P\�f+��<�iԓ�w�m�-ְ�G�)m�qc�ui�69��j[������n+�4[;��@`�K�g����!��H�5W�x�E����?�15�V/�S�O�_Κ@��Eri S������yf�ۣ)�ԅ��' ]�i������ٲR��ӂ�v�����Dx��vњ�j9:�l�_��{�~T�?R�����C�k�l�!EE��Y��`��B�z�ԗ#S������[Y*:8>Y��N�z�Y�v�,:��N��{��dca9$cx�,, 1G+5/���J�����}X�y�%?[� Ð`��(�0S�뛹�#:���8��c����*�&���9�R�4��{X�ӌ~���"�GT���M8�{�u��YL��;3�S9ʵ���w]o��'�m�t6�D�2�R/� ���� �2ԁ�㙵rW��~$���.Cm��Pu�+�C����d�oU~6�f�b���ё�ʑ24Q=�uV���o3�ki��I����2��� 7tt"�h�ӫi�:�N�Q�@��r$3����t^�������(�j�2�	�$!]b�$�?2#�u_:�ྔk��<  -�+�z~*��}J���d��Z���i����L
=Jh��z���[ũ����ǜ�Ȯ�U�Ny��0M���q�f$4��Hd$Y�(����*��G��`����߁r�zRA₵{�<�/!}�6Pvg�,A~�i����u�%.������oĸ���S-<���|���������b���xHyIѭ+x��N���Z.d}CB랤ףHAI��>i�����c
j�_�����B٥�~�ܵ=d]�HE&�!���P,�Љ��ĭ�`I��4̌�L��gz����w�S�D�{��L�G���de��"��`��{u',�-��Z笢��}@dC�Eh�s��'s�du��C�X㔱b��/3�aL��of�����=�zu�|�@u�A*����M����(ڏ��e�0
��O��l�U���\��"�k3��r��Ђ��e�����M��u��>�D�a?�6(��R˿]��R�N���(\@Z��N��hLM0�����1�43��k%8����*Rn�vx����|�c���)�9N����V����I���AQo~�G�	�s�� y�����΢�~�j�K&%����: �A��ע��D+|��������Ě3�>Rz��_E�vp���
�`��=���Ak/�ӽL��:@�˝�~��p��ww�VH���>�ns=����0�b�ܬ�R[9����QA;,j�\�N\E�f�z����v������r��ۻ
J��e�D5FןĦ}��]��忝`��E������Pi᜖�ZG���N��	�ˤ ���%x ��A�`<&fr��.�G�����'S�'�9K��Z�\�V�"�XԷ��^��"���I�g�͸�G�ć��3� ��.���zk���/7]�)��������y����ٕe�t�Ճ�W����d'�	�^i�`�W��q�\�w�d�������	�f*r5^P�L�I�dSH�w�g��[ݚ��64.��Zb�V�˿���}���{�M��w�%���A�-�<o]�_�Xž=W��6���5�պ�r��M����v1�#Uj�PY��$z8t@�ZMԸkPN.���c�rZ�1K�Ξ�O��U!�ߪPw��_���Gv{���n�bDD�\���q�%6+�<��� \�I�y�0���p�� ��[}V�@�.}*{G��#�GT5u��T�"Ӕ�s%-�BxSV�w��:�A�qe��$I����`�{��ͽ��Vam)���7DШ{��f|&	R��|� v��iK��vT�m(��ag���A?�N�iR��^�1;?")�i�'cĦ)��\��_���QKB���7_��D�ҸH n�&s�����QCa� ��kvp�A�%	�W�u{���gƊC[���d�Gs�� іީ7PDb�"��8��Ú?�pZ�Sfs�r0~8~DL����ʍoqᨻ8R%�r�O;�jΐ��J���(,���^U�`�T�t�p5F/֕�n�M���@��@uʑ���*�>݇���H�?0:��Γw&�.l�0��	9gz�5su�x��\$���b^��.�ފ�D��(,D�4��K��1$2��e��S�.񒏮���A��� ��;�O���M�ޤ�׫�i�y}�`g��:.��zB ���=��Wga��[��'���u�X,�I����u�T������v	�hw�r<e� op�Qt#&�ʭ��2�}&]��E~@q���� �|���[�7�����#�$B��6+m8O#NE�	˄�p�v��"š�����/��8j��ZGqt��T�gH��0|�U>Ёz��༻p��m�a�kA�E�C1ةg?����<�N&�����'�O�A.+Ĩ����G�s!�y�ő$I9(���RW��DH���o�mX�w�K?L_�d�ꝞI?]���B�~)�Jys��Es ����OxQZ�\�0�n�*�nK����c�4׍�`>˄<!��hT̹ٚ�d_kS�����9����.V���;�Zۨ�_k���s%��f���� �ME�C��x���\|{�1�o_HV���Q�PO�a�ZXZ��i���׃[��j�:�����Q>�}�6�PO5i+�����vϱȥha�aՙ���ʏ�e��CW<���.#Mr�=��Y��KP�ġ��e��U��B�m�փ��ˏ�YK��A�T�QKD��V ��P�w#`�+Y6�-D����f�H�%����A�Ѥ/1��g��SzQ�]�3:��nd3�ѸaR�h�Ȃ�������S��,E�˒/`�]��\t�v����������v�S>�����}�R��p�l�3��󜊄w�؃l���f�N�����4�|9���׃�˃0h[c�KOț���ޜឡ��rG�[���&7�2�w{y� �椒�
Z�{*^/��Tb���˻\=R���������{�o����L��74
�g�^��Pg�±|dj�|�9��>�ͧ=aхI�����>�����W=¦������?wZ��]�� �v�A�k��m����~,hg�����U��Ar�3���{djE�F�r���d�k
��t�x�w�!q�VnVqPf 4=��0IJ�M²�`4X/y|z���-�ݍ�d����`f�ﮮkϐ�(9n��t4P�>`��Q�i��A��
R�Jܣi��:qZ�<�pO��Y[5弒��kI�n|� ���Q�����,��6�\. ake8����'1x$���O��2��K��I���>���!����㪧�t�hdy�=�N��3/�OP���6xTz��Q��R�=�i ���Qh�K�;��`?~�i��؈D �	#���/E����f5�"�x���e�e���/��"J�[f�4�^�
�o�qK��
NF��I�A�9�$���ITX�Wׄ�J��R�y�o�F#M[��">jUtV�-J����bk+'�>S,?{����&P���2;�7�����@ZR5vqaڏ��z:h9����o��~��6�c�P�ۘT�P����7G�>��c��rdPTODT��� Ҵu�˨XY�<��s|�@��k��zN{|�)S��g������}@v,ֆ!���I�6as�f�l����>��݌L1@PP`�3y2����[L.Y�s���8s���C�	������ޯM������Ħ�:p8�
�ևc���<���eNdzI:q���ͮm�/A2���CB�P�"اU�i���O���喝H=P0ʫ63"z|Hʑ�5J()�!~Pg]7�"�$�n2J-7d�-l?�n��?,�,�TJU��C���s�-�ͬ)�ݹ��b�+><�A)�=*���i���#���>#����t7�vA������a�\*�F��6�	����uʻ�Hh@�o�����&�Z��L�� d��J��<��_Q��e�K�w1�[<Ḉ��7Ė��Έ�J �=�Xq%Si]��ٴ��e".8�E̱H�n�7�(�<q�����c}�k3#~F�Hc�)(<�k����b�dP�t����d��r��E[	�r���_�^��\�a��2��~�k���J���:Ћ3yfȪˆT.6�����@�Έ���Ni�P1jԎ�`�2|Gx���<�8�2B�|���`� ܩ�2��XX�:DR{���ܰf�����V3AeV=�\'�<���k��#
�Uv�ٶ�sNT,�Z-�����}��{`Dֆ�"=�?/�eM��l}#�"~�Iךm�Us�Z�;����=��in��Q*�z���>�~0�T��=s��ǳ�h4 ��� ��]a��b��Ec�����D�:.�����1��_��ϯ��T���-KZ���KB� �:`�0}�ki�&�n�8��|��{h��w^?3OD���8�{��5%5�
�>��o����2ٗ�GT$h���uȟ���љ��2i����Or��H�����G�4=�a���f��s�ӥ��4�����D�#^�Ynim���k���6�V)s.O��M$W�+�U�͗]�@�C�W��>J�}yZ�V7�Hu�ͪ�O�D*c��`WgDh~̴�s��p��tJ���3Zzv�"������O#�YB�
�!�-,�R	�~�i�`2�-2��cT��������^�F���G�J�ʊIU!��4ST�D��Av�����1�b�yT{meu����V�Q�A�'��ܼ���S��^��EEW��VG7Pᐃ=�W�Ui	Ŋ5��ϛ���,/5��ݳ<�k��|HMB�d�^�#�E��:��O�<1�@�D�s[�B�s��n�7ۅX ��NXh��¼LA��s��w@�o��٠�=�=̧+Q��az��YW������-�,9�E�;�ژ�Y�}�:���3�޼mx0��¿�3���e�\tz���<����s�+�NaIƅ�t`7WXCsMd� ���I�UlxK�	�3�;��J�F@zg�a�.�6��������ћ~p�;h��lE�5�K��W�"k_��h�\ǵ}�2�Լ+���O�gӀFk��O�6�"C����
��du��t�A��7�-��K��٢*���sO�m��Z#�mN�qW6Ӫ�ɔ�X�,�}ȏ6�Db�x�M`�ެ����]8��rJ�^��X|=U���Cakg�X_1����)H�e5)��i�0���$��DI�?�e��l���l�{��a��~�Քҡ���<�5�1Q���f���,m�VL�ƹ]��P���e}�����CC;�nTeaM_�@������_�J��~
�8�����f��<r�C#�L{g.�έl���t�쿛q����]�m��{���"����d
�<�әGm��ՙ`gVߢ�0c?���ć�/	�V�s��ed#PkbP��&����ﻔ���ˆ����\J�4x}���D�	��AQ��h����+�*�u�ժ[��}K�d��B�X�O
	H�_�n��>��P��x����uLVA��V��}U���Y5�r2y��v͊h�[�R��y��ny��TK?��-���o�E^#������,�jM@�і�l`�YѪ�AY֚n |X���4	���I���%�o^nHv�L϶x<&	,""Zh�*�&F���h�tQ#w�G:��!ވM�~]�	��	b����ɏ�-�K�4�ڤ�O�ѐ�A�/��W�����Ĵ�ٓ5�r�m�$۶L�����#?R]c=�3}%l+�n���+Շ-��h��6��4+����e����꽊:�;��/e蛍��[��(��K�5��{��P�, H�[)`	�*u!@E]OLY9�͖&_�����%��2#"c��k�ŕ� �>���S�x���F�1��=-w�*{���(x�z�'���3�Q¼SH���K�mfy���&��50�S-ĂEb$�0�1KhO�k#ĵ��ͦX#e���P��VHg��0�m��;O�:��Ap����䂉��J��hh9�&��Y��7�{��O���5���(:�IP�A{.d��x��8ޱ�w�s��g�gIy��k��*5Js/�l�
ڼ6^��cnщ;;$�s�i�5|_����J5du�ͷ�5�~@�o�x�ӡ��gH����H��@j��9����,��R���C<Ľ��Z�*�XpL�j�St�eU�K����ӏ�]M=q�m���ތ�!df���V��/�%J�D�=�dy��a��4��xͯ���Aq����G��8��Ŕwh�;�p��)s},���v��G�j���3���ѭ�;?�ľ��Nl `�%u��@u�����af�r�0H�zgȗ�	� qm�b7��(l����cN�e�q�]���|'~(�3��o�z��jG�t�t������D|[�֟��W� �;�?G�n���sٖ�5Zz;����rٛp�'��5o򣿯�G���C��$��L�L�����K%{n�� [m��x�6j�oi��%Ʌ�|n��Y���g�)�S����6A�B��u�0_�=H�<��rʦ����!J�����ٰ�ۼ�y�����;����0M�T���8X��ܰuj� A�`���`
Y.�qٻ����4t���d}� ���|==������Q(���ҭ� �gG�ߕ�W����R����2�ק=���4��x���¥�|ĺ��}O@txdJ����%J�>�GR���ӵ](d]���`�E��"�=-� I�T����j.�E�V��'w�����%���R���.�� %���'�ve��x5�;��*�ӗ����G�E�����#�WLiˡ"�����ه��E�8��. @�l��boZ������oy �� �HV��R��Q�'�p�������í(!/�!_�9�&���b6h)lt?�/�_�	��A���v�\�Eۆ�	�8.鲤M[�]a�b)�>i ���<=jO	!��␤;/De�S4|^��bV�����K���,�E ��8��0��eb�E5�a�,ZXV�%(,��\^�;�K9�Y�}+,L׮L��'0������9$�(���"��ό�uV��M{�c����UR�S�����]IkL�����Ir���}B��V}����������`�(��R ���"@����L]`��&t8�z�0C��F��_���j������^2h��י���!�*��U�n��'�E"��������yX}�swWB�Ǵ�h����ʑd�������2-�R�k8���~I����Q����7��W4m8�ip��Ս��B��jzn�`�D
��Vp v�����
�nq]��X��G������s��aڧA��ǘp��do��2b�5R�),:|3�܏aRAPy�:LI�!�QO^㈥f5;7��'�|�Q�J^� ��@0D?��z�)8�*1:�C�#�dvT&�L���E`O��"H������8c.�5���h[�м+�W�;P��Uۭg�r�?1$F�{���[����wq��u}g)98̖Jx>+��b$ nȟZ���\��G��B�	1Ǩ9�_��k��&����i{܌�U�;N�ϲ~��\��.S���y����=GM��y�	5��}l���=�����_������n"�p�"���o��)XQ��R�zA�B�nqC#����q0��[��,!���������X�.��սN !t���kK2��I��.���R%WQܗt�����+,�y�0����S���&�b�C2�)u�e����Q2+g��Z@����u%Vv�����z���yBV	'6HC?1 Zn#���9�G�q6!хRj�-�Z�pV�[+�ܸ�A���3�^�o��(��h�s��܋,�r�U�͈�Rр]���*�N�z�L�$}���g��Y]{�Y�ŭm�[�r�H�Jَ��$��7A���0��Ep�ڃ�^Y��:��ns�\(����@r�-���uE���Ugs�Wúf��䮥lҎRs�G3�&�&j�ק��;$��J ��x�"�_$RҐZ)�	�e���a� ��v����w����n��6����D%�8t�55�ׄf�������^yj������B�c�rE�^eXg]`�Nԯ=���J�z�N��W�%�!Oe�g0H�9f:�T�21�c��_�|�B*�T������2��_?�y%�B�A��oB"���,�`�	:Z��Q2�3�����ͣ�#���/���_������u1����1��B�ô��5e��t�d=��?P�\!�I�����l[�#�զ�=X�(�k��d��z��(�W�lF�cP7P�j�]���Y���ZB�D��V0���V9�<t%U,	���:	���ڑ�a����{����́���іU��k$�/��ԑ�A�q+ �%�'@��1��e�;v�� ��l����F�)Cv��,��4�F�\Z�ڒ=�ɢ�2g$�r��{^���Ocv(7g{^o�E��ޜgl3�i~Rq��e�\��n�o�s�!5]�7kU������+�����e#�w�*��=[�|�"�1�~ނw���<��c�f�#�p��i䪤#́@�}�������勘�c� ����������yH`C�|�^r��ł�����6��^������:.�ܳ������Z���d�}��]�7���o�;�@}��������]-�� ���p�H�:�F2Yr�
3���C�C�� bs�*-u���%��=�ܵ�^���hO�?�r����|�����@aO�~3��V�$I-q&<(�U������ȼ�;LN�C�|�×yWo���*X�~�0�[2A,㒝E��s}��y�=��^�Ꮶ�Jq hP��>��)��9|�c�h;&�:T�`B$�V�y-�K܎�f��@m�uqUS�#�Y"����ccI�TLyxםml6?��R#ãYMU�j�_��ZT���f�#�lG$8�����h��!���0K�	�8+^+*�R���C���w�>�<������*Tc�����ׇt�k�U�|���5�v����#.�p���"��߸��댒Y1�#ΚF�	����$H�)%�w�#MT�[,3&�&��i�����Y�Ň�mCY��H)��!3���x�����< �fK������Ci2�k�S���p�HR%ΎP���<�v�a_ͥ5Y3T}�7:��Qg��b�;��.�n�RBF��̨����sz��gy�Ν4�3��w��cۡD�K�H��y��T�j��5.8�L8D&�����l��iN6�H�?�ᅲ�b������ٲlz��,��)5�Ĝ*.k��H��ٍR�)�$h	��(��]�q�}�"���d�*���N^���Cb����f}�7e@ʎ�-����b��]�āuCY��HVA�8�5D��Y����.K���
C�A��6G^��1Ojr5������r	����fh	Q������]�D�m� 'O��)�[�M+}_�?!�ߔ����N���SJ��2p�w�]�؅��A;Z:;@�-mD�'F�;J6G��%}��_9'�X�RĔ�Lz�uk��,o#c�P.�Mu��v�Pa ����f��C�%���̶�9��o���;��kK
Ǔ�*?9�#�P��'*_�����~й�e&0�Y�<�C��:�;Eb8��NF�"B��г�2%ΐ�	�<�5�h��}�#d�f���\�'��6���t���#D�s*r�Zm��(ˡ�JA��l�㭞�&��4�|wL�Vu�P:l���:3�Y�TFƼ	�Z�����1�xg��Ĩ&%6S����Ӏ	�-3A��A��)��f�X+]��v��(�����8N�L���u2�릑#��S�`u޾�A��.`4>�PR���["ms!���5��/��c�wjj��W�mE���상�)��,��C�?j\��-=���7����H�=E %I��^NJ��@�	�͕��	^X���	w
��(�5"H#NuM�tH��k`�n1�0�J���5���#�҂�L^a�hTF5�{���I�_���� ԟ�H�!\P��'�C~�6�]#Az��a\)���/7��짖TӘ�?������_YE�~3@�p�]/5Q�� /����ME��%����w�6�=}�iA�Z��d>#	/j����ʩG4��>e�Ӻ�����˚:�K�w+e��Jߺ�銪/&�_q.�ڗ�D�0����ǢBb��ȸ�O�p5]�fu��S������v�u����O�XtT�3��Ʋ	��/K�H�/�+�b
9f樯�Z����k��u�\>dz�>����d�sUW/V�òN7�h�N%m�R�3�O4�)�;슉I�ᯩ��T6OD�h��3�FA��ϩUc�X=k�GZ�u� �P��1��!��Bׇ`(��i��4���X�W��J��t�W��6�}��]��C�U�83�ڿ�-�'z�>��|��:aX����16K�C�����1�|�1�up�\��F~O�%�|Qn��:Q���m�W.��R�}¿�����tnj�#U.�h�6^u�$(|x[�R"0F#�͠H ��D^o�tI����Z������ڻ�V�CW��>d���%�2�4ٟ��dJ�}�虎��~Y.���O������S����ӗ�v�7U	:��o��=�n��K;��d���hl���f���<��v����� r�;���9|u���䇃����H��H��������-2Z}�|�ڰ �����/f7[|o]�G4��5��Hp��O���	��q�����ԫ��F�yX��@��<����nv���N�x���ů�c�$�HHy�E�����5_CR�\\��_����
��k��tQζ�`�A��w$�A�7�;����>֠��ݣCĨ)�����x��?W�����b�Ar����"��(`q����V��fqa�Q�!�;���\��u�̶��)�B;*{KT��R�ۤZ��L�8�����jOj$ǒ^AS	���K����ce�~Q�Q��Ɗ��!rR	C���`A�C)�i��W��Y[x*�A��(1/��i"�}|�Lm����n:�*��Y�$FH��fl�R(���\���DQ�=0�|�r�^�)z�@Gu��}7����6�y����� +8�z�#O���6��������v_d��Q�iڱ���zh�����/��Z1kam���1��U����9���6�í(n�7���)�֚+�i8�/YZ���J-^��ϒ�U�}@�ܲ�jl9q���{��o$����TT�e��������آ'X̴����.U�m��1T�����'0�[�=6i�6W�����հ�Q���1�:�#ت��Yw�m*~0��(����6#��T���������~	u���x_�?��
�h� �Lt٠��r��;��ǆq%\��<v��IHe�����Π��v�Aj��v'�Q�,/�`�#��mh���䈥w��{��:x�Ǔl����5:�S1��gr�>"��K,s2�П�4���]K-�y�s5T�{^���!Lb���
	�
��O�qe�/A�C`�c@$%�ל���Iby�H��Fp����G�C��Q�/�N�T�a�L����DT݅(���Y�Rjg�G�/��md8�����y��O����,�Q#p~
Rڿ��e�EvT�r���F�cg��p���s5�en����ؼ�*��%( �%"�\\�U�]�Z��	����#���p�d����^7WqT%�[~�f�jw�/-��8"�-Q	c��ɍ�.�,�Gn���Z�� O�}+�Q�-���V����gV�%Nfھ��K
����P�磛s�<��U/]���2��g��W����0�*�B�ͅ����g�ˊ�3_����]������Ni������?�]=�N
iߌ�w�7�mU�ǋ�M@�V�����+�s�B���A�?t�_Z4	�ZJP�DJи�o�pj�5$^�}@ے���zwK���naw&=E�������d��&�CG�s������WT:Z�gW\�Y W�d��
�^���QP"�����U/H��!AWiO67Ug�1�-'���D�@����������fE|����H�b���|��CSSl;�&����� ��n���y�㜸��T`�5Cw��Р  זB�9$7
t}�˛Et���<��B���'�]4X�����P�W/ѐ�b  X�r�ZJ��@ΐ�n����Y'7;�~5Ԯ�P(H����@�;�*0�BLV7��2@��>-����04O������!jKU &N0g���Ӛ�*`nݐ�&��	���n���a��=��UU�++F@��J��p?���mW&�R굠�.������񔖚����Z�*-��'-�E�s�7�g��Q/F�$�����f~5�v7$]~T���58�+�]:	�&��h�#CМ��"ѿ	1
��on�J��(�,O�(���?�<	�P��z�.r����/|)�O��KQX��g
b�Ċ�Bd���T��P2�y�t١���g<���n���J��\�0�<+�C�$�qܔ�ˀ���$��m���̾��9�焚]62��Ǫz�k�����G�ZlRj�����7��ᖺc,�'<͏7o!�x��_Tuw�%l�䷯�}�mq�$z�&bɯE����)�K2��� ���)��J�7ZC�0E��ym��<��ȞE6l��z���w>���f}����k���@�[�5_�� }�6H�Z@=�o�H.��!-/�a>§�m���m�����1�)�}�<��F�c�qc�
�~;P۔[aucD�[ѯs���%Or�� p1^�[|�[,,��s�]�N�(7E��{���	d��t*h#,"v\oF� =/��G%l�R������Y����$�s���ˎ���}(l�]���a<�V{��f:�g{��GC�Z��r���}F�QDp"���N ��1�T�"IQ�6o�d�J��t���-�3�bLLI��aB$o7�T��0��K��p��fT�а���.����G��i�����i�WP:��*�4٭� �(�%�Z闺a��<�j@�q����+��l�u�S�4 2ynR�r��ꙶp
�`�����{w�a�����-�O�4�a���!hp��_���?�H��Q0-��M�E��̷Y<�Vb�I�5�,ϧ����K�H�H���@mi�U2$$�G��gh��1��W@*����u1���)]���7QG�
��'�PK�тE(N��M��#_~H`�T�͸n�[��E���|vV#�ֱ��0�0���*���#/�ն�d�EF�ݚձ�O�,�@�B�*����	d|�[��3�a��[3ؙ����pٌN]u��`��\
�m�t�x���n��IA�^��3:�]E�����fz��\����B�DQ��㏼0�[}��[y��#�l�K��I�,��Ͼ���։��y"��b+e�mB��h�e��k4�ڭ��"U��fu���R�
�v�R��J�8�.���4,G "c��| ���E�A�\���#i��{$!������2����݄�k��迕FO�I�i �l�
e���L��0p�&Иݕ�Yy���Y�D�P)���?&�9�h���b��q���m�7�������bF�1�~Ț�┟�ѕ�D�H��%�Ѭ�C�=+w�g>D�k��$ҤA������/Cո.ظ�1,2��&'z肦c� ��7S$�?/3�n�!Z v��r�0�^�U��^f?v�B�F�)")�O&�ш��&9R�rnRq����;���_�OA�|F ��{�E/]́���8����8 D;?��-����A��lhkt��"ؘ��s��_�iN�Ⴭ�D��ǵw�G@��$"âB=���!�}����j
b����t�W�V[����Q��L��=9������B�K\ϟ8�X&��P7�ਇ�z�k��+�V�1�>Bu�fsz��]uF�:�O���W�vo�Zq+���*�:�x���g$���S�:'O��'ǽ�6(�z�9���O��5p��lN�?.8U��C�#%T��j�.<�Ζ�@��6|��(V��%�f!�͹&�B�fi���6�_]�֧��F ��܆�X�5%�?;`t�ۓ�b!;��5�}-��j�)X�w0�p��dN�Y��Q)H>��U-�����[��uSN�A2���	yی���M>�J�D��_v�C,MY�˪��ح`���EQ�UU�ݩX?���U�;vO���>�r�������G��w����B�q"��K�Ц����:��h������qq7@��e$�M�$�QDx�d0���ጧ>_|�Bդ[_ߔ(��m�T�c�%������q����>q��R��A�k�,뛢p��|�x�hQ(ʤ^��g���u�H[k��=��4b�5�]��Kd� -z(&�3CA�v�u` t����A��^w��D��n�r�p�||�ӗ�������Ii������Y�	Տ��*>���>���S+^�m����,Iz5�W��^W��\]Cx�uJ��q�}�M�h1��7�#�L�S�d�c۶�e Rɨ,��96/��N��>O�C��n���&Xq`�s��Ҫt�e>���-/�Wzh���`�ʗ��W�P����A�r������ޑl���o�i��lK�f�C��dM��*�O�gf�p��-�j2��M���{���B:_�ª��&�x�6Ϗ�fJ�{��1�{�69����Ue�;�s^��2�y�8DI����i'=�s��t��s�y���V���9-s��r�'�2���h�{�y�y���l6j}"�_�I��M��0�����?M5�"���O�X�)̉r߇���c���� ����r��t��9�=�.��k�]���8/��{�ݸ��>��2��蟩ؒSR��t��0�'A���Z�8�qN��7U �bf��!H��?��4��6��X�`U�+O�B!�~"J�b�?~*k;ݡ��7�/(�;���1��b.�g�egCy�&�R6�9��M����1�1#�!�{"Kl|E�p���^��}�U��^#h��yh[��;��3A��X�-�����0��#0���/m\yl{�3��IB�g={`�0Tlh�Ҵ|I��C���΁�'ֳ��<�_�N�9!x��LP0(F�3lӮ�l�0�I�O�=�t���[2�O�x�Ǌ ��[�t$h�9x,˴��#�����٪�^/~�`E#�?�'P��J4�F�=[�=IWc�s�jT��Va�Ѱל�y߾0���;�����g�� ��M����o���T��	.���jR�&$�ZH�^�D-H�`�IU�F�a
S��&�q���i��>��;M�P;�q�ᄾ^<b�k*%�k�����+4��09�X�gȸ(��.3 *�����Q|������i��J�pk� ��ƕ��dvL]�Ë�On/z�ȟO�l)n8T�U�m!�V�������c�&���qK�M�x,S�MP�T�Z����G�d�~���>�2:��|���N$�p�ƻ��T���������I���NC�^A*�6� ?��p>Ǡb�n*}�Sk7��K{�	�I�}WL�� �Xug�p���ʳq昉��D� ��S�y�lӰ��A��)��M�<۾�7��Q��9x�Ze���}"�_%�J�y�ex2u4wH�ï��9h�3xNsp���V����a�kK)�<�ܫ�B�Uι���*K�=S�s"�Pp.(�Z�n���<]�2{Wˢ���v�ɛ%��_l���S�w�.H<�ޕ_�bOpz�Bz�!���HaU��5:��%]B �ar
^�
��� ��)�ZE@�^p��y���ȧ��'�/�B�q����]���u��Z��!/����k��:���M?�5vFǜ/�,����2&��p�1&���x�����k��Y��"rxl�KEg1�:%>_5B���T*����kc)�A�/��yH$Ш���^�E�&_�4�>���ace�� ���Z�wD�8EK�j��BL��>k�5�J-�6|�t<WA�äw�۸,���Ƹ(���J�c��q�v+]	��p���D�#B�N-�V��a�5&���l��,UmB�f�b�Hܴ?{�x�[X ��Q>p��4M�%�������h�q��$%A�ϩ�"�?���0�IŽ�D�<Q�������$�aQ�H^�y�+��������Og���_�dT��^�����&�*��@u��gx�jk�eb�Sj��:�)J$�aQU��:�8K7G�6lZ�?��U�tV����Ъ�TQ���:��f���T���@�\�@3U�û���fm\[&��lۋ�\���3���Y�G�*���B�,΋�.��Vj����F5��O@�}S�d��&�ՒQ?�C��K�m�& �,���x�B�YA2%��F�o�"�sV��a�F��{j�vH\a��Z�v3�� ��
�8 ��Qt-ɂ�KMߝ\O�߯s-6sL��첖=�21��S#$�",�ȁ�I��T�l5��0���\E%Ȍ�Irb;)r�����N|�P"�0�}����������îFu��\Wfq&��M�����\Xk��juC)(+
��-�71���Y�PR��%Ĵ|j�@9�D�~�Wڎ��t�_
A�
���2�s������}�
��r(�X����Q�<Z�]����$�"�ø��V}��b!| ��H���S2H����MC|!�
��t�@CΖS	So~�6��y�&̊c$4� �(�`���� g��٘|]L�l!�8r��7�M���
���<ɞ?�V��q'Ř�֡�_H��ܹ�U�ɛ͈��Q��A~'�|
�:q<�O�|W��0�	��̞EnG���fS5��%�Ia�6M]֛�L�.F5�a.����r=sc��_�I^V���'x����6��#�7�F	l0�&��O$+�F	�������p�D�ޘ`��h��q'�sh��m�F���Dߝ�gD��U�J�M��[���$�}Z�.\�?(��ɩ�Tќ������nz>z��d¹j�UY������f���ʑߡjD�9�#4D��m,tS{�6�e4p���D9`I�+EAi��B!��6�N�����
N����(�x4�jy���T��%`��������2-����[�i�Bk��&zQ{� ڠw7Bȝ��e�&y��O�颱VwHY�Rt� ˆim�[����k�Q�O�Zj��"1cͭ���KFtw!��f�]V\B�&�>���b<Y-�j�M���f~X)zq9֗|s�Y�b�a�L<A"c�`bn�����q�a�V^��[�S̙�8����XF��0��,�a�����E8q�#?�SI)�XMi��!��;�ǄY<� ��{��>Q�5 II���U��' �u��s�%p-,��y���,�Q�֒�������7���k�,�#�c�X,��������N�#0^���ˋqJy�nYov��Y�0v�nG M������xg@�<��  ZMƺrX�*B� ��klm	������VZ�
G����4*�=3����Fh_6y$:�5k-��Y��J���v�À*��xLAM@�IS�
X���[���ޡ��D�%� ��q0�)#pgH~�4���Ű �IKo�N��
�eJ�����@���'����	�Dz����8���Ҝ�@�4��eա�����#�)Q�^���~�\���}�4c�{
�NDF��h�~���D�,����d�����B�r��'�Csa<j6���s�a�ಽ� 6����W�=t��s}1�.i`�o˰ڠ���Y'�i@��_I���T�8Kn�'��r���
~B��i�L
,����leXusPʉ�1p���FA�[8��f��/��Ka�Sl䲋��[�� y����M�ݏ�ϖOM�RgS_�8�[���1�oϕR�Hݖ_]�
��XMK@��-8�*�v�iP�ֵ+u�����\A��+���r��B�$�*q�:��RWҟ�����w��%ï���K�n��<4��1���X�X[i/��ո��w�Z ��;A�0����ok��WPe G�Iֺ�ih�!������c��X�	י���9���y��3��gco��T�G�~�T�D	M$���>y�+`�&���*�'���w��MH[�f৙�?^Xs703eэ���\�ja��US��'��S��.�Pa\�5�R�*C��/�'�Ncv1����^���7�"����Zٴ"�Z.O�xDUj9�v��)� z#'�� �0�&�:��>�'ӿ	��F?�'0X�3�B�j ��p�[XH'Dpٽ�x}zA���Ӥ��m�΍�prpfզ��?N��Kq��[7
��Mj��y��QL�w:���~6-x�g=�P)����O��|�tN�NOwk6�:�l�����ر�ıy����BF\��xyv���X�!/��OB��F/B���|��Cp��Fw�"�W�<�O�W����MGHgi�������:b��D([�֥��˵��u^h6j%9�rt��G�� �Ѽ���Uk�#�W��+�D_��閟k��A�Y7���~��y������g�N�4��L
�TƲ�,�f����*>���Vl��2z�y֥��@� ��t��Jh�����DsK�m���}˞=�C력JT���O .�=���L�a����Y�X7\��`�Cj9� @�1KOz�[*3ÇP�<�mJ�*��T��8L$��6R��Q| � }Ut��F�)�ǋP�v�[�g���Q"���K�P�N�x&ǭ���{H�>5#OdFܢň�;�#U��}r���de]Q�����*�V�#��c"?��Cu��ڂ��H��,TU�A�N�!ڢI�����6	���̐A#K����P#(�k6��/0��D`6y�a�B;0�Q��]+����'��4�n}ՑSj�GYA?�Q�&���'���*�9��B-���q+QU�nt��Z�����ށE/Q��dU\����������wyp�]/lWR�L�I1��«W1��xF���R/2������P�����)���`��c�,с�=���F<ς�:�9��1�^?�V�v�,�;������M�&(�i��%/V�5�4�|xq�L,��]'K�*�M>���!�؍vJ�r��`˺&�}��T�r��h T���p��'�*����2Q�h�;w��e��گ'��/ժK�2&ܪ�&����i�i����-��{����5�]���n/��dw�rqv ��G���b���>G-���8p���- 0KW���d���O�Q�k�ol��v��"��\^m��$�;���"��` n�ԝn��.b����t�G���U��.nA���)����(z��a�5hҊ�z;��/+9�2^�bS�d���a��]��ƀ�S���.�L�@�^�@�v��BD?�w)�[}�����@V9ᾀ��&˶�n����Q߅�27I�1���E�m���� e�:>W������ .�6�e�;�s�<KC�.�|��g�>q����z��ѕh��h�+�z����$�����5�bd���O2�I�D?c�C�.@��c�u�T��0�9����˂岞ȇIZH�5l(b[�Z[d���4����عX^~�I˯/��bz���pe*o5��PG;�n��^�A��v�k�@,������]��D�o��������~����J��9iXS�h��Z���N-bp�&E!w���>��buڐ����6Q�4���[��VnV)��p�w���`�'���#I ���k�U�?6�%Q�u��/	/ﰖXЂ�2��泬q�Cff�jf��;�1LC�e��h��������U(�p5��Ӟ!���7���G?_�k����6s�7p���o��$m�ȌZ��1kBZ����5c�ȅ@�j	�����Np�l��j����Vr�oޭ'A���s���&�">Y��������X�u��wGo�A'��Mg�}�Rh����N��E����)wx]EY�0�U	Ms^�
�MI�g8?��b���8�L���d���g]�����>|��P˩��$xsx$h�]�1质֌{9Pl��u /�*v�1ߩhrD����ui�A���;^��9�%���X��3��1&!]���x ������T�����KPg{ƻ���]~)Lh�@[E�睌� ��<��ⵤ-i7�1��H�u����mER���&o:�e�E�z�G��8����}M�+�u?sn���"��������9�]��h�y@	��2�x1��z�֫$<.,Ƽ�x� 3�ʉ�D<]�'C�(z�ğD�v-/,���Z&~��\C�!�&1����B�D������A��a�Ϩ�C��*��G�p���B9�N��O��8PB���h���\w�B�/*�,h�'=yd�ޣ�@��>�1���`v&��""�����G���Ig&b ��Jx�_�N���>���B���ܤ��I���j�I�t���V��)	9���l��wm���TsAIk=#N#�jCx��)�|N�D�����)��#1N!d��e����S@rD�V��=D�x�'l.�m�B������w�Ų��u[� ?�̓+S��S2$�-g�zn��C�����m�en!]�փ���jӲ���{�l�~|��w��a	+� M0�46}��a��=l��e�����C/�ΆQ�<rX�5h�t��Xu����2����E��.𰫳�%����ձ�/�'&O_ُb9�З�8j"w�~��e*)�����~t�>]x���otF.و�bAѡ$�Opw���<��(̛�ֵ����1م8��c�0:�|�΍��m�_��Y����q�8b1�'�O��t��t����{�`���}�
���R�
��?T��?6�o`��,:����Ҥ�,c��,��H0���貮�7��'���jAAZ�2)�g2��X��m�������0d�㟱J�pcB�%������8��� X�҉i�TF!J�%,��t��_��y��:�`ZJ�B�n]��u��5,���S8�t5'�C47�s)�T19���<r��q��JN�ǎ���д�敃�N�i�r�����Э���0�ě\~�����f��0A��R]GV�w�)��#�+�U�c�+�F�����7��n!Ǝ�|�H{*�t'��U�i?�|H�q�V�(���r��H"��d$��(��S��z��zaI.����hbp>�z�QV8�Ĵ�R�OXH�͈��iN��N@xj�ݤ�(Z;~�Z���[
ۢ�% ��|����,�T���Ѥ�h���n�4��nV�%o�`��,���6�#�?��\��$]=�Jm���5���N�xNw/�~x�ㅶ������u*#��[��a�ĳ��d���j;Y/���1��v�j�@�9��x�u�`��042~&5S��x��U��t��э��׀h���uC.=�Q~�����6��\��Օ5��GȘ	+2f��un�����CN3��ɝ�>�6�$|���y�$���+c\�g3zZi�,���y�m��1��1}�����^�u��e�w��Y�r�&�4dG�����<�	���CA`�H����Ќ:��6$"���:��Z�S0릺�H�<�+eI��']��� O�\���g�R'�W�Q�bL#�d�R���^�ٯ�`�*cxM8���\� �m˖�Y[L���J�{H���L(V���� ���X�>`�#�]�vO�s��B�;�ow���Rp�% �EQɵ5	�ɩ�}C�@�>�Qq'��	�O�G�W��F��?�r)!�u�)hSI_F#�G��(���R �-*
K�e�A�֍p��G%�z���H���L<��뉼���c`ɤY�~�Ŭ�d�'��gZ����Y��J/���5л�>2�O.�4��و���e�1�qjq�d�;�6���{Хk	9q�Z?� ՈK ���
�T�5�.���f�7O�jQ5ǋ~��fEı2t`���=����T���d�FT�|�����删 g����O�\a�*��T���p"�,꽔��Ǩ(���H_|�( ��h2�����Jw��;th
Ȇ�E�@p���{Ɉ)0Y�r�U��>ˤ6���*��!�3
�5�*�ћ!,j��K���3~U�d�ά�9%W�#�\�@���l^���^e�q�'$1v�M���V�Ol�m^ifzj��H�c��8��B&Ґɷ�*���"/�*H��l�͕˛���交*Y�J�ťXf�W�� 뎠�Q���-��|�o��jt,hE�Ãö��9��JaYJ��^nd�/xb�U��H�l��Fb��}�W�>l��{�~�h�	r�6�|�5}"�nr�O4�d�F�$��W�R�. k���0�
K��]�6̌ĕ���.7t����)�J0�mΦ����@�9|O��9��qWВ
�~�}��љ��t����Va^ɴR�ȼ��Í5��3FCK�"r�h���p�/J���k�  ��A�a�TN��n+���B`�*Kqd�+ ��]���@�� 0@���D�;��zp�X9}�a��@pIW4�{�=��M�����I0���Z�Ce��E���ۈE���aQ��P�屑4����I4������t#}ew�8T竎M������	�] @���%�/ƞ-��\��]��� �]������[&<��?�3�?�%Z�O{v����$��e���;N�ϊp�
hOa��'��W�١��6���	�K������$(!�z�.f��D�S�`�ZPZ!2�e[����w�"T��~�|��c0����D\Շ�"{�"S"���,�#�V���1�S���"�6q�'���c*���C�9%'��Y/Q��f�7�$�E:�tV/�ɤ,C������oD�T�$�' �$r�~��5~d��Bvv��S��v��h3����i���5� Y�"y���E��|�,Q������T��O7ZM�	_��=5݊Q� /~rn7��7����2dک.ygAz��u���'Ok�Z��`�`�P�9�ֽ*�~a�Fj��UY=�G�1�WV�o(��ڍ���V��y�����B�U�W*�o��T����" ���~e#�c����|���?�aa�̑�x���֒��H����H���@��\��n+�ʙ<��4Di`�b����n�qi�d'�]��u9G��"��r���H(��\D�7 Ĳ;��H8���{��5-\i������kN�&:T��Kn��O7�������N� G�$���s�Z39U��$�D�T�\�����C�?�,$��f�蝁�]���"���!�.��m5���bq�F���C�t�t�L��Qr��5g�Ѯ�X6��%-���6ݎ���\~� H���ʔCʋH�Q"�;��E#���tMA�/c<�B^�4zh�*��IͪڄA���o�>}������F��Ns�E��fO���9���T�`iޥon-���4�k��P�ˆ#_�G�,�n[Qq�Zkԭ��B�SX�$�H����W\�_j����SN�$������H �"�A9a���@\񊄎�i��q�m�+��#a���N}iuϜ))����v�eY��r���B|�z���r �_!�#��9�a#H��H��ĽmC�!�^��D?��6咽`���RU���&�wY��wC������	��MT����ަ& ��d���9�~
n���ޞ�
;(�H�zv��-~�̈z�'0<\��i�^�ܸ-��[�<|i�u�C� ���/ŗiY��)d�df �t��(�:=g�$������R^�7{�~�����D�;��H&��N��A��g����dX�V+����Kڅ�'r@�X�a� �������귘�t��zȮ�2�҉N��j$��A�=G���O�@��$��2"y� ���Rc�*��%c���k�>� 9a�jQ]3�0��+e'<R����f�}��S�rv؉�>���M���P����1����+ ��>&�L��f0���c���8=�H�/�}�)�&�I[�������e�ۯ^�Rd����ұ�s�z�p�Nt�|q�)}�$;'I�U=W �rǌ�{��l����^1ͬ=�"!l��<Y}�*��bY����&_�#^��Y���W��M[��]�~�rYov���2���Q��<4�zv
�{��A���-+o��
:D�6p!�@��x���F_���1�Ulb��'�Hy�l����4Y��Vh����$�f0�r�@}�o��Q~�j=e-ɫ��;��-L��l@>lJ�0?/u�1X�8w�Fu�V�����f��	���c2�Ȫ�����b?۟iDh���٠T��;ɫq�p"Ų�5g�I�-�}sNj�#��m��ZT -�{�I�u��{1?�r����2�C��|	���X��׫1  �m�%r��;ns 1�ɮ_���8�����@�\���-�|o�-u��M�ߡ��g��-��挼ȕ T?�+�rz��C�C�g��
���X�.G6�,��&�B|�\�����!Ԇ�ZϿX4���"l3�� ̄��$�18=d�$�@�V��㛢|�c���J��Ao��2|���Ȳ�X�އODժ�`����͏I]�r��)��N�g���koj�,��҃�4�%��&�.Z��rm��!>��f�N��N�I���-��R SJ�=8y�}�!�l�3y�3���7;�X�?��<x�-�/�vO��z�rrL=��")
��D�i�<(:9�A3WTp�� �P�9`#��m��{P)��@��k���zh���j�ɠ�ЏT��7��l��N\T�dqa8�/��]����~8j�{�
̸@{o�h�-��0B2� .PRb̍`��D,� R'��r/&�]�/ilut7⯻$+��Sܮ�a+R6�lfA��v�������2���T�9��@��t��m�x�{"�q7��4��+���AzwR5��?8ǚ4ś~s4�㢩#��^�n�?F%M������t��̚0�Ya�2�<\$�����4'9<Ӡ�3��X�N��ͪ?]����v^�ێ8�/rq�GU2��	�.1��4��pB���D9ŋ⼉��d�Q����7��:���jfSiFL��{���3 &Hr���F�}��I?�Ä�4u���r�ف��m��aI=��ۮ]����TQH�Q4!�T�*׼��[�V�eCl��R�C㔋�G��y ,�S[`U�Ĝ��ʰ:e����.V�b!��!�/��p�:q.;ʄn!�+O�P�c��ŋ'd�Wz�*��A�RΆBx�����Q��a`$��#�-�%\�=#䧃��T�a,Q�B�gRD�0�BF����ߩ�
3�{)OV���j]P��y�׈�~h�f��,���$��{�V���+��/ ��ؙW�ԇl���v�VW�c�h|RG gy��-���Z7�O�Y����|��ݖL-��e$�ve��W��pa4Z5����&�)5)����h�&��\3;�#��i�c������IG����)�|G@�+|j\�y�	۱%I�;ӭ�{<3��\����p�6a@�։��"�5?k�Ơ�!C���X��B��}	T}�'�{UP	�a?C�7LB���,6��H�V�)����b!���[X'�#w�o�Nۦ�Eҧ�C�5�/�-�y�A�DX���_2�QˊژQ�i^B��3植�x���"р��K�J���?N�l�Ȩ�h>1�-_�j���n��r
'`HN�<y��`�J���3�g�%yY��N�)|`�`�B��z�˜z��|�`��R� ^'ċ��L󻰼�x�?�H�- ��l����-�|W�
�^ ������x�Q��3�����=�p�*<;�ʠ�!�\[�1�갅hB�Ng�3�GhY�E���>�f�vXd��H��������&���%g\X�#ѐ���	����=���t�_��#�U�HB-G�I�,WW��Hg�{��q��u����{�Z4�UNhQ�W�uX�e���|x�sΝ|Ȟ����[(?�����`K��H�����o�hބ�
z"u�v��.���g��^m\4��)�Y:L]�	�wx����V�0�B�# �Y}]t.��h�B�8�|%��pm�>���(R}����ɥuoE6e�!W9��У4Vb#�H��y٩BS���
�>��[{�B=S��+������3��*���z�vc![���ţV
B?ϋ�P�����b��d�?��\yN:��ivh5�fW����d@�Xm�D����D�LVF�=��<�Ag���D^�H�V@��nx�&$v��'Ni���!t	jN��]���e���X��(vVa��&�!�CQr�ƭ�L��?o�9	�9S�ئ����`0��,����e������y͡b�r�;��~ڶ�H7_�L���z�s�W�$ϣ�VI��Y9������:��D��TS��Z�4~�RӌdA>+��ߴ�-��^�W�<��	���V�Q�����t�~���8�����p�4�¥����E3D�άKQZx;����;I˽����L��8���
�ʮ��R+\?Z�����?�ֶ�M�m��hA�����Ij��d�SVBE����U�+\c"�*�(�h�B��p
�hH��Ǟ�g�	��LhZ�rj3��j8�Q�'��jܿF)�m�O��'$�f��u�޶3�ƹ��N��8&�L�[�L���ױ	j@qg��p�_=�4�� +Π�ٞ:]3��'@#6 ���8;�QS���WM�j7-����-R� �w�e�~�)��p�̼�
L�����21޵㴿p\98(�z�G�� ْ.��K���F���w�O���Q���3+6G���p�}��#�����/�N�ȏ���%���,}W���I�6�?yh�1��N����gU�L�N��'�Ġ��m�-�6�X��iTνK�<B��EM�p"��Rw��y9t��$�����v�>���]�L�9IoQ��E��w�]��,$�s�GVL8�S����;�?(��a�r�V*���)��� U54�9^�P(�_z�A>���>�ʮgrwo�&a:ʩ�/^�.��sO�c���!Hv	:��OL��3 !�`�Gw�u��EJξ�K���9(�ʠEo/)R��h���ϳE$h!���SQ�_�k�O�೦���6�-��;����I���uL�c�߬�>��w-��b�iϏ�v�)����Ai(�$�hp{.tp��1����c�i��#����j3݌'���̘r-��pv,��yQ?eG��ψ���}z�t/=��v=�+n&�B:�5���(��]��饆&�� �ڝ`8��O�਎'K*��TіN������Y�ivAwoi�� ���,��J����Uat_�c1Ί[����7���]C���5�!�bUz��+�j=g�>� �H��)�5��}w+"��T�9k�Oo8%3;���0G�D����P�{�a���HC���+]0<V>%6��~���]�̯�^a���,�3��t�v�?J����B鍘�������L���ۑ���E���(\����Җ���1�>�NZF��y%�_^N(p[��A��U+W�OokSRգ�j��F>��՘iPm�ks@MX��Z7�2|�_q�a�^�煍ak;����@>uaN�,AE�k��uhn�,5�0�y�n�x:Nq�{�l�ؙ���8��xT_�R������HyH��-!�����x˕󎎘Pi��3�`/>C��s�Hp,�|�?��(��D��*�W����<�.�T��z����%D_����
��Et�[q���+y�����#j�jw[�k�r��c4��q�r��w�](��jW�m'�y��=�H�lڌ;g7h�7�O^+ѳw����q �zc�H5��5`��M8Q6�F���e�F�ч��P�]]�&7o��F@e���4l
_- �d�F��t6j��kt�O�0��K�0y��h_2i&r�Qy���qS��N{��-P�Vx3a4hvsZt�K�$�c?��!��eNg|��D�8~�˖���	k�V�XqW
d�-����G���P���<?��;�� y<^���R�@���2�~N�+�"����)i�`fl�kn<����E�n�H�$-%���Wģlw�6x�Ҋ�)�Zn������)'��82��P�ˉ�W����Mp�=O��`�^�%�c�H<cd��T��MS��~:��@���wf���4��SS�̞f��n`�-3�H�p��y߼�W��i�&NcP�1�u���|����0COʩ�ի�K��aSܴ�>5���tG*�~�v�/q���I �uK�9��@<L[3����P"��x��7�
{x+�K��]��1 �W'F%��S�.5"vbΚ3��4�a򋶹�9e&��o��/����r��o�S��ߟ4v�MS�;/��̀H��E̚[n�A�4
{u�pc��Ka#!f�wb��ww����$��O�+�dR̛��C:�5	A�|�t�yB��/�^�O� Ħ���z�lR3���+��,k)�x&o^9��"G�|�)n���b)�V�~l�m�����+��F�g��o�v���?�:�|�p0s���W@Ê�+9Iö�j�ᔿ��!
�h�ƣ���\������W�y�q���mH�϶�m9W�~Kz�~^O*��)�!��� e%^?��h�����D~�iQm,��Y��w�S�i���+�`�0qu_���DlD�Ϥ_�-Z�{�su���왣o�])���A�G�K�i�\��L�J�����#�x��(
��>�R�\��Y��[��~��~�ܴX�$~/Y+��d��xծHqm7N[]�&hIv���W*[�;j�#�P��iu��F��=�GG��f�<���~�f�Y�7�ʁ8�#=�����+��[v���uޭX�=疉�����p��
_19�]��dA}�����	��6f��F�~��7#�V�Y.�r��!>���A�����9;4~�8�.�/M���G��
�+�ò6����aC��Y�C@;���^�2�/pq�b���9��`�&KD��$��
˛��^	ɴC
����$[�xωG ���Y٩��?�Lt ?�AD�¬s�I�dt't���b��=Mc��1�{|�BM��4��c�7K�*�$�i����&�6(���3%j��aSz2$�8�q�L�0�FAzrܐ�{b��+ܨͰ�J_	ֹ��E}��3�A�i]�4��w�W`�r<�
��tT!��� ���5�Q"Ӌ��DX�^<�c���p���4b�,��0@hͩ�ϵD����o��8��c,cj�#�u�b�$�Jl���s3!v���-��0`���h�Br��i�5A_�p�;�G�R0���Sk��E�����N�h�H�B1�*Q��5�U$��yU����S}�.��a��J��=���\�ÔS��n���x1��t���%.����ܹ��>��
�(?f�W�w�������<g�K��Y�����  8�6�����8�܀kqx�.�Cǒ����o0XN�+������ϔ��i���w߿���8v��ǚ[�l������c���c�>̭+��̢��x�ϸ1q��\��hSr�{s�C̚��%�P+���!�'vc�	�.���[�`�:���w�0��EUÝ�J5��:�m+
r���f����GȔ����p�,,���7KFť@�����'�w��I轐X�| ��:*��P ���sB� �X1�/�"��� �u-�R'Ƶ"����F�Xf`�0p\X.]Z6Fږ���]�pQ�%�0�aY���iMn��~rh��<R��֦�U3���h���m����j�<��'��V1s�kU�?�v���)sc@ ����7~��m�m! '���R�V�e�,���N%#�� �g�Y<8�[Ѡ����!d���Bw�w��d�Jo���c�b�i�lM�e�}.f�;8G��I���p�Sܼ<H��~�E��[C���T9cew��ƴ������r���ψ΃"�9��0&ԡjn���O��b���� �L�&y?}���X��(� ����y!rY�E�����வ,7S��p�̆^��B6ƕe{�d��@P[!ǖ�Mp��H��EC��A�+ޕ���d�]y��V'�?�����r-)�|�d<)[��>��-wK5��uC�m�5��k�C(;lX���ƥ0�Fd�49�]L>�5U����YG��?x�2��H�$�ؘ��TX�Ճ�$�K�l��*{�.��ױ��G񛼊��ϯ���
�7�mj�״l��s�*��NBF�5w_����0�e�G�߀U�G{�	�T8ZS��6��x旝�����v�$�W21�ɿSРnH��@�Su=R�.�������(�(gϏ����_��K��=I��[���A���a�>˖� I�I�G�ΆZ,gNhP���c�	���B���,"�=��ŭ�?)kԣ��>�}R�d���Uj� �'���=�,d���T�'���R�썝?�l�zܲ��8�`}o����<����W�
i��u�7/'��^L�f�N4���7���V��e�s"6q��+x��=f�{�s�`��33�?ig����s�����J��t"�<p����u�ln�n���LO��������?�3�W,��L�ߣ/B�Q�5����������"R��8c�x�{�Br*�N��!y����cj�Bo�2�[���'�F��t�k�WpCpYؽ����%�1�p̀��`+�2P����Hq�i���V��S׈��ܯ$D��[Sdc�n���k/��*�O��5�0���6H�9���&������m疞�X��4��>F�6d�u<����c՟�gf	p!}U�V���鸓�p�T���*F-G�{5�J���̈m!0�>��p����|�p5i�:i���A��^'���;WW~��8:��Z�XI��}�U4n����F�s$�s&���PP_�ǎjS��y���NP#��)����f!��t�uO��ΏFUgGTsJe�v�9�q_8�݆8`!IrR�e��g2o� %����^"��Ē����]�/�	H���<��F\< q댠����J�F���H�VQ�a��ͽSs~�Ej�H-P�]uT��b�6
�bzG5�a������>�n��?l��i�]SI)�0��d%&M�~_���5�kn�|B ��=�k��}AErӥ�~�*�:�r.JVT�3#!Z����C�(g��Ơ�W(������A�>}��{�{򑢘vB�/Ң:V������'���_��h{I�3&���~ ����վ���N�w~�'2�P�f	���;�U)=?�čI���-��4y:��5&�_�B�K��AYdה޽���`ba��V�� �#�8/�v=jn�h�<���k` +k���(�ƴ��yb�_�Zn{�SX}�m�	cbe�������B5]Xg��öw��hr/^���-���Ww��4��@8�V���p���S��f}$��u4��Ƹ���p���.�i�� h,��IN�O��m	F2R��F��d���ķ�C �����On,�'�U�U|h!E��
�������M����H���3�����P5�ڡ����{BTjb6,R�;R�tx��9�LY�A�g��)�݉Ǘ�Z��1�D�d�_�;=-��!J��[�H����Oo)b�+li�>^s�<��۱u�l�W�P���k���|�J���i�tPl���K���S�_r�|�⽓0�\Zk&��S�w��}p���imy�
�2����8�^F�>�f�wt�� z!��g���kJ*7���AW�UNKGT�����DM�}���6�A��乑������2�g�X�s��uMz��B�ɍ��E�K�Aޯ\.!n
� jElH��s�k�L��O��f�4���p�0c#zGR��Fu��������y+����:�O��h�"h H�j�܍�OZ<��y�/�t�>1�¢q2�h���1���H�v�AY\cW��z��|?�J��u�M qyg&䜀�<Ȃ'w,�޴�5����$��)�|^~������r$f����&z�nl'�^�H���H��u#f��T2YK�_�o3��갑�膚��}[y7EsU�o1�@���Ǐbs`?੎K�������4�6���Kj�NF��F�7�!��܁�w����+�^ˡ,#�C��ý���G��-��(�V\�Ml����i�"jj$���fD]����= ���^9��J�woR���y�G�a�7|Y� ��!��~y���[��9�XEJaSN�����~Z=c�.K�8�u�q��(����z3e����|�.|�:U�P�ͼi�&F;��֓�u?3�_+��i�jj׃hB(<}�`��t�R��<�����r����pW�-�̜��-��6�,�_hٔMy��;`x���3B�A\�uO�x���RA��Y/r�L/�����!�d��	�,w#.�ӌ(iCp�j����FC(��%�RԜ��Ĳq�ǎLT������X:�0�4%�H�ɺ�H��E���a��5��+�i�.���Y�՘�B|�FHuZ60�JY�Ѱz���{��%("���_2�K4]`Kycx��y�z�ɴ'���k��8e5�=7�G�w��J	9�a�`��%���&��p

_8bzy��l&,�ٯ�,��r5I��*��V�rj	/���kg��ٺ���$�C�2�[+C����E.G2�'9^�����
=CrbZx�q547T��:����t��甘%��LR+�бqݬ��FlѬ��lZ���L�mȬO�!3��fI7g���#���R��������+���l�[�K��Ns�� �t��w����#�$����\oL�0���^.�+��n�?��&��%~��X�e�)�N������ޞ�"�^�����_�T�K���z�P/�G���$�-'C�2����'�W{���X�tH��V����;VvwU�B��:2o����,a�ob���b�nǘgG{ߑ����>إW����a�	@���Z���|�.&9ڼb�����N�`�ɂ�#�8�/7��y{_w%0���Rf4C���Uy+i���Hrj��  ?S�O�C�% �1N=�5����|����cકf����9���L3���X�2J ��Ln�u�F���Ks�.ԡ-E>��S�T�L�q�ݯ�Z
��A3J
ڏ�7�E�d	��5�h �2�1�t|!W9/���
�څ���eV�D0�� Y_I��˗���[E���n��!�4_�
�vZ�cĺ�l❑��(Lz��,� �o�m�4��;�6�{Yi��8+h���<Eu�U���~��ܝ� 7��S������r/��\)Ƕ�G쭰�=�������I�ZuH�H7/*�{mN��Q��O4�,|y�����G�h4L ����y�D�W�a��ݍî���\�*|Xs��£-���E�F�az�n������b�F`.|)[5����`L)*+���rʋ�և���W�ۧ��&Pz9Z����٭�!�^�:m���*7��e��&m����N���$����T�1��(7��{Øӿ�Z	۩o�$��vi^wx���Oc�Y�N��dTp��t�|��@=<�fw��ʣ�.�Ww;�u��7|�L�ZA�0�f��&&d�;��Q���=^�9�(=���C�H�n����Bu��x�]]mO?Rk��t"\�>K�)xa�;xL'��m���d��½K��NRW@:��e��##Rx�7_�4[׹O��2:4�L�=�eWI]~�%@�S}dIs�������?���N�<Rwd��dM�6b�ѮȦ[��I�k�&����4��A6�ɻ ;V�n|[x�6Ѥ�[�;lsS����aF��0� xG������$z�j��ĩT[V�"g�^���6EV^��x���H�8�?t��X�@��^�2���M������e ��Tς����]�� �ȑ���+SՕPd��[-���E�i��o��Eǅ��
x�%�ip�J��*�_���}�� �n\�s��m��u����<V�����7#���χ&�p���،o��H��B������ި��D�ˋ���1�Ƨ�T��}��逈�5�5�G!r�O 1�N�t�(AW_O��7
U˗�rj��(J�*J�*:x$�{̆?�?�c�!�Y��_̣V���^�JX$��]�c��D�k�j����u�����Jw��ȍ9��&��/�r.�k���Ű��4TO��b�^��[�+��d���x�1>
 =����+}�LJ��$��w�����X$�1\�[
xO�^��7��S� 0��耥r(U��Kإ'~6"��#a{��q�Tk��ߦX�R�?Q:Kw�%԰���<5T;YC����p�&�Q�b�d^I�Vx��8���B��X��;Tg�fY��K�w�۪r�a���W�H���r���9�qQw�ur�b;���s��?jM+gX,�Y�x��4��!e�X3N�hE<BD��K.*K��q͸�x �$Jw�f��Gd�_�Z
���7 ������M����Z~˯� ����;���hP}����z� ��~C��=�Q�o�0��Omo���C>�q�z1yD��㽾q3�%H9 vj���iB�C��Q��<e��U3j3[�[��i�d���*ݕ�n�G����L��n@TE�7֏��'��3�ݕ�tE�۽�8.rZD7un����P�]g�<��W�TP�OV�f
�9X:��m��;�5[-
ɞ R�`t�4�Ou�Q븆q>64���y�mY}�����d����9�U.�l5��T���Zq���t���q�=���kN�wN���pV��0֩�Ēʾ��n�����5Ph�	��kdP'3n�!,�$+/<�/ñ��W�@|d7�Y���=Z�����6
+P�M/�cj�܀iQ�O�I�&ϗ�)��F���fC��	vz�4E��(�K�����"p�/@�I��p�\U,�
��A|nW�Q�K�lڭ#�� �LFSp�14
2�=���������i+:�Swg�w����-�w4�r�:�A��$<���fs(��,%Ӭ/�\��5 F���%���x��% �Lֺ~�	��K�a�>C�OS��[�, <��"��������͆I@Vm;l2Dĉy����W3�O�$���]�����d1L�w���PgRl��uP�W�[hp�JIli�1ҥ)�+�����^0$��*!���kLٺ�ľ��˿����%�|*Z��C^�