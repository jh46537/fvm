��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k{de���ӱ��.�|�2n���Hx���]|��36rJ}�}��dE�F�Ԗ�W���h�p{�{�v��?/B���75J�l���{�)EƊ<Po���������U&��&��)����w"��<�;l߮��k��D�yH���D�j'8��\��f�-�m����j}�8�vU2j�$�i=�~ج���a�1+�\�&k��ͷ�#����Ƒ'T��z��l$O�9�J��é(�7������X=XͰL�vW*Ĥ�{g��m|����U�%���8����Pמa#���B�8pH*��1I��n�w8�}��w(�zl��fb�uE�SM A�h ��"���S�Sm�-r���XR\��!��u�KOM����p�Q����Iw��Pn�%QƮ�hr��}�e�^��"��}�,��҆׳�yfK^����Cu�8�\t���i�|}���]�x2�&>$-[S#�Yk#�I7�񓛤'�F�K�b��Z;6���YA�,��c�O�����*���G��;�p?����U�5PG�"�h��=ϿL\���� n  %cO'2� �^7_����ٚ����X�׷�'�S1�џ���;�$�;pOk��6u��D`�;RhGi��p�DcG�rޢK�'B�ɂ�&*���FL׳�V��Sb�$4n��#���*u>�O��9� 8�c��I�2C�0�&�����l:�����@bg��g����D��n [�������F���O	�)���Y�^��L��{^D<��b&y3��Q3=��c(K��ė�����ϊ�@CWP����Ϲ׫� Y5�W�}5�c!dmle�<�:Sϐ0G�l�)�VG�_��1�A���* �4S�e{E�W�Oᢅ�>pѯU5ёU�FK�o�`�kWU �W��f�(�H9��6�z��w���K��ޤu�7>%5E��~�`�H[M�c�#^XE:LUD��ȴ�F�,�*�O��`'�`>|g	�DMT���ͧ�m$�;�f��kW��A���#�y�I���a�|@d�oE\Ǵ#1�!!�����'�I)D�H��Nɧ��[ ���L���82@�K����o�["��zh��"��]�ͅA�l�����x�!��҈��b��x���������.B�-��R��)�Y�W^�z����4(�{��6�ެRvR�s-���%��zK1�d'�y�ѶY�Ke��T��1�����z�㞾�z;	�%��+V��s�Ɵ�SJ��5a�Db<D�Ƅ���gU���ۦ�TOv�j�Z�nÂU��iI�p��R��g���;�a!^�yjg�L���崼2��}��>�pqj��yթ��'�l)�:@����Pb��~)غXG�Ѹ܉�!S[�ϩ�S��
�<Й��e�u�OD-K{l�&�S0؆���8ӟ�2��C��p8�	���Cw1�*No��;h�J袼��$��W��s���5�&P>I�a��T_ź$K����璌���\�۾=�Kۋ|�dq�#U������*��mB+N_U��2�q!��0� ����0�š�_MS�yw��|�BեΙ���i�Y�K��;O8�:�6��ѿUo�'���`��nq���=9|����%)7����#IQc7�̈́�o[Ks�ۡ�B�.. x�lM��^�F8ᅾ�)�M�����n�M�����2����A�
�7��w��镵��}�Mq��^t�s�= �+C�4������bmPm�М_~bC��"OgB��?�&��t�<}��!ɇ�v�!�ɝ�*6��s�]./]f�u����k��C��e>�c����%�N�:�%��c��ޙuN���R�~pR�O���֢�/�43Z�L��v�u�R^&�ܞV66�A�t�e"l<H�R��9�7��$��v�a��k���Ȗ��roɒ��^>�1�%�4��?$|��I2�)��tj��sQ)8 F��?�}z;;x���l8!3w�YI�g��+���P���y��n��y�"�3�:V��}kC ���ЖB9v�����\��s�rau����Q�˱A�ô�P�|/��C�(r�2{A"�FĔ�T��u�s/�i��җ�<K�)�J��=UW8��a9���Z��3h��+9܄w�	C��6�fk&NW�*xa%�X���Ŷ��c7hV�E�	C˽�&hSt�[�5�,8��t4�7�C����C���A���:��4���]>���Nݯ�	CKV&�]��]e�����}=������b�L�檩�o E�V��%В��k���`�L�qa��댗�/�|��Z�k8S�e*��K8<B����4�zJ��w��6>
٨*#�U��C�vjL���u�Z� c�W}��R7Q=���sڃL<����Y�v�+"qo"�G�