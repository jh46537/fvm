��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"��Ia�W�� 2Ch���E��ʡ0
<���촚n�/qo�����>��i��3�ց�'�Q����%@C��ɥ�X��ݐ�K��/>�[��3��7v��i�|�\�S�qGq�~@@8&���T(Z� �8��.G�	��$�KBzdX�M#��7hU���*ǰa���'�^�u����I����= )�8.����f�q����|$f!�ky�ȼ�_fz��}���L�fH��B�Q�=`5�y�[ �D��w��#�G�|Ŝ���V����E�y��/����fx��i�`�:�^z]J��"���Ns$C�0�W�g�k�2l�ꩬ�L�� �y<X��=���A	5�QukJ#���^�Yj�T;�(|�I��9�{*��%M�4�m�$�=���h���͗������_�*�7��w������-xu3�z�#:��e�+%��ݾ�๳0
 OR*�����CKoQ!{E��#g��P;7f�@�c�=FK��2hg�%��bji��3-�Ī͕��=�I�m�䁄'���E���C����f-N���Z�eԈ���-��}f|󼾝^t�4ū�N���NZ1[���Ńp�E�m�#��ϕԟ0&u���w���~�PyP(���2� �	=�0�]uS%�=a���س��<����i�	��S=����Xd�׺r�u��_t�-24\��H��u��f���^�"Xc�uP������C���Hu�V��L.���T[t��8�d���=Q�`�J�T�:�J��I���< �7Vh���"��h���w� EWc�x�_���
e�W��P�K������YI�߾����@d��8��,��FF��#�
/�\�(���g"�vx��ym�j�n��Md�H��P��Ug���Ә��ީ���:�<sͳ���):������ ��d�d���,@���mx�U�6�M{�_�.���!�֜��8�(�#w���̖[��0�7�L&Զ����D�D�:�d���Ӓk�킙!�7ЛbQY��[�t�v��G��v���SD�ƫ*L�Ҿ�6��l�?�9ܻ����i$7��7��A!���r����q\_y�������C���*��Uf]Z!f
1J�n;Jd�Ү�H:Q��}d}�;�aoǊ![d�k�Rł鷚��b��������4��M0�S���}�@�8f/V ��Ck��  ���CC? ��!-�������"�� @&�\6?E�Y0	�ֻo���X��Q�<7���9cW"S��R1J�/獴��
˲�%�^ԙ�3����������H+�`����V��r�>�8��'�/���M�`��b�%h�S��Ws@��雔x�Ũ��C��u�C�t+=�&է���;�Jjf�����(���;�i�<NQ�W���S	������$� X����n~��'*�>� ��f �^�̅�U����.��^Y��%�o!��;��JĢ\-�=��N�:˳�'6��K���0�>~����5�Q%�9q- �{�{���t��R���[^<��"��{w�1k��z