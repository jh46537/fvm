��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����,��f9t���3>��Ձ�A�7M ��uj��M�0��{�ơ�Wa=Kg��!洭D�2�&�6����2�����X܋��x� ����G1���w�S��3�C�1�9��1+CH�<3�vwN��F�T�\#[�'I���ҒO*K��V�6�k%���D��Sn�&$Y�au��Q�/���OO .�XS}���9��k,[=0�hj��V���w��:g�!,;�(���1��+�\�dn�-�],L+߿+����.Y��67I�OK�^��^^u"�g������X⛚���ݱ,��t?;�\�����ϟq�0<j������n���r�^}�3���B;���75�po	��l���a�#Q�8,�;J}�[��M�ob�^r�:i�O�P�n�ߠ���%�;��%z��P�b\���?�;n��V������Y+X�t{�,�ȼY�����
���K�����y�,�]E�e���DӸ��ם���+�G_��р؉:��	�v��꼴�d}o&%��!�Y�³YUb��I�;��҃l�(̝�����|�6��^d+! 7��+9\Ǹi��g�M�N.��g����ɓ�������nC	ЩMB�:v�sb�9��X�[
�������+@��٤)�>_L՚`u�| �F
�mj�Ͼ��Υ��F/N\^Aa��D���6њ} "�]jG" DǓp�7�J��6���ll�#İO��'O���T�F�ۆ�nP%�98��= g��X4ǳX�`4ʿ���/#��/��n��ޯ�a�LF�ku<��S����abm6�o�ȫ>�w�N�P���}�u�O,2�k���d�⯈�H�����P�+����$��Ⳙ8�& :%ԋ�5��PģkI���uH$6�/R����S��T�x֠�p�3r�\uG��������$��s˫�.��^��Ԝ�b

:�@�vU�1C���a�젘_Xn���n%2/��M�~G���S][�����O��e.��f�Y�م�<{�#+�:�����T��J�����_��!{�j�5��Z���a��c����B�4�=��sk����W,��P�Ž��`�&���R� �d��@��\�d���ң(Q�s9�O�g޳�UƱ�2n[d@�!�NT�k ���
��v�����uW�5�{�ގK⁉���(�gl6�{��vM�������������T��c{be?�ds����s[J����i���а&�|k
I������X�]�Dκ���D]��:�.	� 
+�W�E�?�����/AO���V�z�9���j��tf�u�}T�|�*�H�L�T�5Z�`���S��&����V'�54h??:�V�˨�%7���]P�����3�*����d�>Q
C>�e�f�]����k2#.X&I��Z�Y�=&G�P$�z�n�m�V�]�B{L��+GB꫏�$�O���,����,������e���}N7��N��u�$-&���8�B�V4�e��y<}��y�Z�?b�P�?�,�?����Qq���=m�9h��f�6���e0'�%����[��tjvO8�;|�5��\$w��+G5�H�<�ޥ�Wp�9�»�t�b�Ts�h��R���j��UW�T�E���LA���W!k5��C���jp#�[\�3]��.^テ2b2wS$�ԝ�S�}Zz'2UMwƻ�_4��?��)���1�3�*��*@Dh��� �vt��O&v�ک٣�T��l���"��K����\�)<#*��H�������֮`N�%���^�x��?oM)�]�!Lh�U5��W7���0n��Rm��>nc�-[ S�p]�͊��r�E��b�4gB� ����� (����x�g`���9/W���U`�0?I��D�ɘ�(����!T�S/���PVo���J ������\�x:��])�F��ChZ�,�HC�X��{Ȉ<�,3'-_�[�a�n;�"�E,�d9b�؋&���
n�]���y}�P�x�+�|�B%���m|w]&цx(
ab:t)WS�9��˯-�������J��2�G�ϜN��R�ܦׅ���_O����S���X�0 �Z�������Я���,5>	���g8�\ctm��Bki24wµ�Z�7�"�+?I)�j��{1�#(�sV�%����|h��y����Ў{b�=v�w�h���˯H� �Ծ&d�1W����B��[�X5�7�@ʡ���`+���z�
-��C��(Cp��hQ��w*�D6D* ���tæ�nB2@אN�F�b�b��%�Nƺ�]�����$���ؗ� ΂�x��\\��ҝ��+N�Šj��*=�lj�Ed��r������;:O���^��:�����������1��hI�_�T�\L� 
,_�(���s��7R2�ϲ-����:�^楈����	�/�װ��徎�z��{T=�C���fP�Ka� �h�eY�ޡ�"�E�󻢠#��zaX�|���������	�g�d���¹N#�S�Y�8�U���#*$�&o�W��_s�&��_�5N\S�:��\�C�e��:OSۗ�+����Uܔ�B� �z�}&���G�So	iw��+F$����x�痖)��)�
���c�i=W��H΂�N6H�C"��R����oWK�I�_��������d�ՐK{C����=�հ�G�����f����o�J�!M�a����t�P+ūXgL�(Q�Z�0���������	��ν�Si��Q>�.��d2M��O|��p�`NAY���0��B�{���9��t�+�� ��'x��2���!;�[�e�Hⴻ�J
�bNCH��LP0e2�i�	%��tw��Z��Yt�.v�yT�q2#��(�u^��|0�r%^컱��zq��mN�B��gƗ�-���s��F?�B����J���+Qc&��\��:�Sf �q+6�?:S�@�r���
+p��3xW���S0��EM�!�O��wư�f�˨��$�u�����5��U*{���Z�zg��e�QW���+�l�{�к�S_ej�txʕ,�����j�~mq�(Zˏ6Y��m���f���� ����p�9�/PK�C�}����ZILK~�4�� fmf��e���@��;e!H�B������&�����x�0��`�!�{��E(MǬT�Xv)�5�Qu/�P�}���W���1�l7*=Z��#YN��vh
9v�0�����~�RwNT�GA��Z��V��֝�#�i���=gfے�a��2�I\�I���Jo�W���5-���P��^��Z$�9����7��0�,55����q nL��18�OƐ�d:4n�e{���w���حr��ºǕ�r)�F��dQCL}�<�Ժ�: +�e�<��FK��c�A���ð{�_u��S1�L�ă�+J6"�x����D����-ڠwA~�����	dr#�THŻ� 7���1�±��f<�.͒�}��ʜ�h9����SgJ
&��m4ĸ�u�}���� Ov�p�b��!��
u���a{6�+�&�l����t�N�u�@��l7L���M�@�MW�*.Y����됿1Kd�SHg� ���z{m�K>�#=�������l����t��v�����_ZX�Mlde΋�c�Ո�9ʺe=��z>ʭC�S�pU�����7���[U��~��.	�8T��kK���h��&Zvl��|x<�c|��D��R�jG������_yIod%�bjCh�Y`�/z�>��r�{љ����Z�
ݣ	\�ޤ�`�v�X�]
��a\��2���W�T���YV#,������\m"Q`�F�l�ƶtyi�M���,*��� �]M��rD2�@-�a��)�(ƱA�d�-s'��d$��>��j8���'<�JxoHp1�w�h6�1�ט��c�R�E9�À�-T����#2G�b��G"��1�uŶ �/�IGv�-�2k8I<�P�T�6�'��6��,j^�Q&�:�cݘ�Y�dY�p��|̅��]���~5�͗A�j�:���1m���2�-�%}\��gg����z�<��������dˁ�S`�T_5|��njV�����N�/�'�Ȩ1`��N�a�p��Nf����W
�pS�f�TX���,z:P��K*[��y7�"�;��Z<W&>�A4�~�J_Fbu��U���&#e��}�滰�_��kMS��ɿ�$!�7�}��q�q~���~�᩵�:�_�*� u�␠��WS�&̢I؀-��u�iG�1 ���Et� ��8!FxZ�u�)i��e����xq����a�NT?C3�L����/�bZ��
��ݰ�m�p�����*5�Kn�9�<|�%�j��t�܋��U��,J�=$5B��<A�uj0>"Ss��Wg�غ�pi����5I��s��!D[��M��>�bNm~�q?�3�U,U�$��-Qe#�5�t�.g,�N")H��7E����Px������H�(��ם��#7�<�j��s��c��<�'d~�F��1��x����@���"��~�?�X���n�0 f�����A�	7�e���� �Ѧ`.���:|��������Y����A���һ?�+gj� +
7Dd�2�#��U0b�G6��!	7bd���aڥfc51��L�W����6��r��L`�@���/��F�e�[R���$�t�]R$��6+�t������s�3���t
���W@K�m�Y���XG�`V�?#�1D
�B�'(ց�p7p�b�3+�F�4}���p�e�J�imU��]	��� .
#~W���|�-h
ӂ�5��o��^ߴHg�uf9��.�7��&:O��!�I�f:��o@�܊q2��<V�B���2�uQ�G�@��5|�o��q0�<iJn#?�B �����<v�;�Bs��Ԁ����d��&�7	���ae���i�<�u˃��� {��J0.�����ے��e���}*�G[��ю�٣֛�G���"��xA�G:d�|�O��������.���8��VJN@P�OP˩LU͔v��K�U�;|*=H�n�}����J�t~�.�����h���L/�༖�RzQ��VEj
7P��6�4RH.r���җ�E��d���am4R�6d�=+y��c�[Nu��t���OJsKڔ��߬e#	Y�r��̑����(�bg�:l��|V�}'���������'�bhTA�^�Ĩ�b�pZ���v�=r��qʺ4�J8��Ia;4O̶��R'��%�� �_X�B��Η��9���Xɲ����h2�p!H��H���~��o�	��T�Lk����̉:�m�{w��R�N��c���^8 ���y��ٮKpn([:a���������5���3��S�c<E���[�]4�a;g����Aɧd��%*��K@��O�T��s�Ջ�;���l��� ř ��p��$ �DT����r�����E��ɕ4��l̶6}W-M�{W{�۹�����r���ӥ�z#qä�)ۗ#H�D�v�����'�}rv�p�*�����'�Z?@�^�w��5�^��Pw$ū�I������g��n��0�������$a9b�t�+_�?���P����;������s�q�*�*����)걫���X�`�[(���n�$��c�B� w��|��u�?���n.�z���*����PC;��+yϱ�E����uW=dJ>�v�Us��s�eP�`�.�	� Uk���ㄹm�Oڐ���ai@z��"H&�AnKa.�1����Z��Q6�D��O�QJ�9{s�����������)��'6��}���V
\�w� |^f0詷����ϔ)'U��Td�Rc6ϐ�/0&�9_S��Ȥ��>S[�� ���q.8�.��L�+�T<L�ÞϫI�nc����^mق|0�T�sذ������ʜ��	n|f�	�wK��w����&ú��\�����*�o��T/,Џ]��}���g�1��c���[\�5+�<I�p2�=L�6�^�0���E�a��a^�-�E��"�($�`n��I��@,G^�J�?'m�4K��3��Z:IK��;�.�JD-�>g���7���H���Np��2v����������lg%����z�dzF�U��"�ؕ�M��q�]����R��B�c;�Ɔk�c�Ҭ���Jo������<ׅC����j l��qF/���
?C@$�y�<���^�F�ꍄu��/L�T��Ρ[g�?���ė;>�W�|$z�ݲ�a�ޔӪk���NHo�����{C:�/[�����z�6Lb"�tN�\�����}�i���|#�ܤ�Mf�=N����qo��7=|��`��}�wnc��R�2��6Qq}�I-l��m{V�-�G����@��"E�s����1 T�"��ե��-w��6 $�R�2n:%��k?�#rE�Ӄ��q��4�����p���Hf�?��
�X�P\,����e����	K����Ýn��Ǝ�0�̐p����4��!x�&��QBC��!A���L�|���Q���	|�i"�i�%#t4L�8�!mі�\����;��WB���g��1��v`��)�����v���!YK�H�O�n�b�ʇ���#"@|����kن���Kc�����h��*�/(q抔+�z��Eu����%fB;�R���BR�ޛ����M��B��
f�`q��vN�iA!s��K�D�Br-]T�gj����8ǞL�)�:�)Fe��D~~��������S�'`.�W7���`żuF�V8�>踋�įy�G@<����T�ܶ�td�>@J��m��%2	���<����S=�s��H�n��ہ���"��sX����O�6���dئ���e^�l �ʿ���:�-a�I1ܤ��%���W,�h�D����L2��ұ8��>�K��ݍ�U("D���9��XI��C�O��(Mu�92��[�I�>�9���wY}�d�ƆG0�u-��)�ǛsT ���(�.�sJ|!����ȫ�,q��(/�O%�~%?Z�},�����Y�NS�Ҭрж���������̸�j��AC��R�5&�.����������7��r���*���C���r��ĺ	�i����ڵ63-B�
=OU���v��=�A�%:�so_�F���#��ˣ�; ͒�����~a����2���ꩤ0X���}�Y6�Gj.<	T:c��FY.d!9N�q��9uK":w�dn\�i_�@c�O��X~�jO[�"�>*�β�虯g�A���Ɛf>(�}��2|�7ٸ�LE�B�SC�7�Cj����	�����u�$6K�;@��Pp�.Z:��D���Xd
B��!��&��aaL���mg���d�~k4�����"D�=ܺ��v��ܨ켓7�|n��������C�(z��S&s�
>�Z3���`��V{f%���k��x���$��G�
��r���ƹ�I$[�31�W7n�!	���-�ܾ҈v�k��#�˃2:�Q�鲒�?w��!�n^����/<Su���d��o:)M&čeZ�eP�Y�Un`ʧ<"nD��&��F�>�AG��9�TUb@dLh$��ř�^��%��l�	b���U��Y��S��G5�zY��\V��Ԫj�\ّW#�kx���XF;v�V\�oہ�j#�.��Z@O������ܡ_�������������l�Kְp08�[�=f4��z��0GX�w8-U�̝. ��=���A�5��T���D�g��#�u�@�!:�#��zi����U/��I.��� �����h?�C�����P|�#V޳f6Z�-A���Ѭ�*dT��� G��Us�9�PZ�Z�XN��꾕c�|(Rj���= �"���ڦ���DlZ�������mqڠ`�	��P�%�B_��X��{%���x�.�R��*��owZ���{�A�Dg��K1!;��F��X�N��?�J=C�R����d��=�4��p�0�{��*��i��ǼՀ�N�٪���&'�wcg.ȠIt����*9���V�e��\8�Q~�C���z�Jtb�'�TI6�t��=s�Y�@��S}�7p�߃���:�޻�#���SI�1;d��@h*�;�~Bu�S�qU�>.8za}Jɧ����~c�Q��aЮىk���+���Y!����:��dVh`��y�F�>��Z=&�/��.��L��o��'��D`D���=:��;��F:�(Yܺg@��$A_�8��	6<�{����F�&ڥ�n�+���rpy�B�7>��b��+���䭹m�gpK��"�o${���\��.�T6&d]`�*���|G�
�,�cfs�>{&��K��.��|웵p�c`�f��.��P��BP�/=����qQ�w��T�$%]�gi:���J��?в�1	15!E�*ǌ]f�y���-AV��h�ؼʣ+l3����q��}ØzR-Z-��vfP� !C���&�2���`9%+�$ ^[:����i,�k1 f� ɤ˿���� ��` ��nZ����P�d��訛���T9.g9C���e�z��㺐&AՌ�ُ����n�����7}��Q�j���ׅx!?�gaʝ�UA£+���W &��E߬���T�$(g��%�����o�OZ����־n��s>���4���ܠ~ O#�Ѥ5&��JtD��}H?���O�#)�<~*x�3�SuE��	0L=΅?tỏnB��!(�O=���37
6u�*�M��v˅:�z%�Ng��A��/����!�@o0�tu�I-�io?SIW,��P�rw�p-F����x:�?H:�&1�R(�H����A�
��.���=о�:���W8��jW�o�T���a����ϡ�-`��h�8�c��#�F:Y�CO��nV�h���MV-�"�Jk3�m��b  ��Jig���Ӄ���ڦ�]�&�s�,��Y�h��K.�\��a���������zzj�'踊ʵ�@��_ք2�y�p5w��T޿l��^qMLj�*�-�Ev2���g�O�, M:��]�(#[���,?����M����TpPiu{~��30N/޳�����~���n�7�q5f�׈䈢�4m�}T�"����wk�(�������p�<��X!��|-'zA�m/-�^�����t�~������G��`���lq�,�dP�-�)�P�v�+�� �����2��D��W����β�I_|�E�}c2���t+�4s���,��W>�p^_ȕV��{�h���1��7�8�; �(�O>��y'�ƻ�;�+K������7s�UPj�K��9 \J{���d�T�x��т~���T��p��>���D	�لh.�\�\.�v����@��N�}�M������$}�����z��OQ����<�K���2AqQ�舒���1��d�hO�<��{�/!cF����Б�\�V_�
SsG�.8P^/���k�al�/����w���C2>��cX�p����w��1	�g�:=U;�@�9�-S��H��]�H�wH��*����Y�\3�w�1���d��$�"5�4U�v{�iæ?L�ľ��'�'(�lU��jjR��Ne�(=�8�d��ɚG���:Y���T��}}~3��B�XJCB�����96{�J�z\ �F��T�6����Uy��3�_��PE3@��s}�1��`���4�ױ�2�?����7	b&5�cz�= p 1�*�
l�o��J�
�8'�?KE#6�X��ɣ=M���$t��m,Ώ�2Uˌ��E�����R�M]k�$vp-��Q�N+�)M���b^S@3��y��2I���w߿��K�DL��"��O��7g;v1��2gK�L�E6'ϡ�m���c�T֌�R�!`7��ۗ4�_�"iȷ��h�1Q���EpԽt�^�A�;r+Gf��ם��诮�f�����c�+�iE��� �|i�O>bt=7]��<��������\�x�5��2#��֊�ʩ儿B�B"���é�C^W @��K��]���+hRN�T_�i�3u�Ф3��B��GA%踭ai<�ޜ�b$r��*��'��A�����tgJ�F%�nV�iQ��P����t�����I.i�cٰ�d���L1�L��ؙ$�Խ�[E�� ն�; �m	��b��Y8�*I2_����P��T��U�_hm�>A�"��m������G�𔆿�q����&�j?�V���t\!?�����JÉK1�������;_-C�1�WhT����XN6R���A�X8�f�A��T�T�aw_#
�0o���r*�D�K�
�h	:��J{ܘ�C�^�KnB�&����6�z�O�f�/�|E},����=�����h���K��,�+n��\���mU/�:�bX�"�O���.	�c��]��:���u�U8o����}���$D�f�[�]v�3+=��D-� %�F�+=C�JQ��\�P��*�O8� ���?J!�c1%Y��ֺg~��sd���'5�-�;�V�^R3� `�l	�ܨ�_���=��ÿ0�9ϭ�:���@���u�h��/KW
9�����(�6[C���b�p�����+�W��܍�������K&�dk��(�F���) moM�*_5�d���~F���u��4�@��ǃ�.;����[�J_�ُ�ez����t��U��އ�$XiЅ��kG@ ��|Q����Ƌq��Tk�w�T��Ðk9'e5~ZO�6�����&��n�賥%$�}
̹M2h�[zw�dC���.�<�Vq�*�ۇ��;�Q��]ykF-�ʫ��$�$��1U �0�J�sJ���^!Z�����lL��Q/%�}��������J:�шjA�	���[����c�R��0j�G���4.�i�S��L�{�J������>��K��ώ��#fq��m�f�#B!�VVձ�+��]�Y��L��Fu�!����{�t?1��}���w@�T�v'�@��Q���G8t�rX+ˢn��k<W����v�"p7��
Y��M5�G�_s}� st+8o���H�g:����	�!e��݉i�R�����ڱy�M���o�K�fM��bI����朏�yP�#v*k1��~v�&�/g�q�F�;��_�����
�bPb������A�����,�Ä.�t!@��h�Ģ�on<'N�����c	VM/Yޘ�1dÕ ���>��'�a7�
��1펆v	��|q�:�9��~�\���S���*�E8vٰ�%��F�U���!C�P��ަ+���%3�D�y
��,T�OS��E��5�ZFJ��_��E�T�3aUi���0��c���=U�̖^��������J~-a:[O�]&�{N�)MQ�aN�����c~ ������G3f�P�Y"�`S�в�	K�b|Ǹ�Ճ5��y}�E��1��u�t���&�D��k��isG6͎k$\�m[��)�x�]�`�C͘*/ ��4
�w�PH=�!��h:���1��X��+0K��ߚ9}b�=��\�ޟ��5Dߵf NI����1�|�1��D`� X��At&�W�$&�ߗ�'[ښ��=�&��e�T�E���� �M�44K����Ӻ@�]kZ��@=�S����˪y�lr�����x�1|Vm��<9�c9�`�k���Rv,$3�},�����,�!"L�u�tط�92a�A�x:г�^��J3sy���Y��j��F�*w��A�ۂ;+���Q=�+MQ�c���a���I*�Bx���0��
�pc����Ǝ�v�"�����DK�4\�c&v{OSs�e�W^�!��Pj�Id����_��/\u9����$R��������ɰ��)�
q�3�謓5���<g�yc]��a/5���Z�~�ҽ���XO���hZ��,8��)� �	�%��>S�j�,��*,�� .ܫ��� 7P�zH��(.mr&7�˻�7,����.cί_�ҽ�G��\U�T�t�RHe�H�U��1z,k�������A�4��@�X�(�ް*W�És6�� ���B�rʌ5��sE�<�T"C��@rg�6�N4�Ⱦ�|�]E(�\i���U�ak��|s0��-�(�:&d^�F<��9Qli7���-#~aE���ܱb�2'�H'O�k}4���Ԝ����/V7�� �����"h�Y9�t��w֗m���s	���x3\�C
2��2���^�h�$��4@���τ�BmuO�� g�>����t�2���ӎ�
>�GI�L��{��H�϶9��sT'�Dy�vCt����blgH����k�Ʋo���V�zJ�k2��<Y-���N�a����;H>^�/E(�v��Ԥ���k)�Ǌ"2W�-VL$��ד�D�C�Lf�}��>@�t��RH�-�?j�7m1m��wI�A�ti��$H9B5B�ُ�Ȝ�Jbw"[���I�02Z�j��p�p��)*��iDr���7��㮤�V)-[�e���Kp1��0�0�p :.�Z��z���"]�ٸ��F��yw��g��e���p�|��z�*��&�i�c��8�7h-�"�`�MW�Ƭ%/���Jde�LG^S �u���Rx������i1����K-��"e㜶K��;�~i��H��+/v���Di_@Rs	a��%���?g�/%nh־�#��l]��T�C��kP9o���o��l��vAV�}��[ɫ$�����8�XokR������Cd�ĝp����fH����*�Ó�ʛ(��%���eN���bh���MV��l��;�������88���F@��O��8X���m�K�3`-�PGōg_9N;�\�m�N��q+�Z�U��	[%R����_j(�85����.X�.���
d�֗����>/Y��J��.�^ �3��ظO��� l��A_e'$�̘W�MZ�@�:3���n-���.�!G����h�Lg����/��[�?|
�e���U�>_VW>$�t{o:�� �"x[�O��36���w?m���m������ڍF��wI�o��D��/�E�+;�Q�������4O�O_��y����V�T�	�g��tg)���![�~��Ly���i�Xk�	���V/ԧsn.��e��K�����էpv�A�}d@K=�_�,u2�^B�S�������𧱌����i��P��&���X?��f"9��|犚�V#x(2{/ǗᣍH�$Y�ޏ�\x�����} �����ѿ��\~8�E��+�y �����2*��l�FP:3����}g�o�^v� Iz�YA�`����tQ�&(NZ`F_Y�k�@��� �<-�x����/�/��f3�J*�x&�N��N�!t�O6{RDҐ|�9�QTR�]���N�"m�����5�]��j�]����d���$m[�X�/����>G��',y� ]���9�0;�p��$�3`)lƎ����b���;� �G�X%���ܠu�3�LW����r�;�<w����s�h�9�Y�A���7bQ�[~ų%�`T�V+�k�!�9�O3Hr�ޅ�7gM��)��#��u���'��a�˲Si��p ���Z�aꊾ��6%h(c�Eqm��3��p��]��#��ˬ���Pˇpx�\�x�M���~N	Z���"��{$�2�?r�
����`�� ��V�j]E0q=|�ёI��޽٧�6&nC��� ���C��ۺ��=%yTuo/���&�L��{�+A�jR>`Un�v�9U��k��3,�h>$`by��z��P�ӛ�j�Ĕ)�%�f���M���������� ~9w�Xˤ�����
cv:�!T�y�SF4Eϥl xHhNT�|�-��e��/����Ɖ��������H�ox�0A���P+-�@MX	@�.|�B �G�ai!��#A���r�{a��L=QR*X�E�؞��1{����^+tW��e�M}�KeƐb�6�eq^���9M�Z� ��Ĝ�c�즡��}��s�+����w���w#���t\��7�@�lXRmt���m�IQ��)3��W�T4�pϻE�l���d�YO��Oa�usޟ��rF̖$�,��_��m�y����D&F�A! ��Ǌ�
��Ŀ��]W��_�)M��lh:7R�n����n(	F�0�`�����`E ��XN�~\�G<U`9�H�$��ΆTD���7J��z��	�ɽ��2^t��P��+��R��":�ŧh�)p
w����~��vg�&	��&�Rm]�$���;��c��Sq���k����v�������yY<S��~��<]������3u�۶7§4����:�+�|�B��Zh� 9��yG�2���/|�V�7xT��-:CyK]�\�Kp�q]�T��6|n_��%���6���z�?Z����|�h4��*��(�����D-�J팼�8��u��p�w�fU���f�9`v�no�:�a#���
GM�oZ)�\�z*��!��ک��!i���l$�1m&�>~��1��憔lC�4�g	�7#����$��A�Z	�IB<��+�-l"8�Uj·���Jئ`۽���9���ۻT#,;p+��6V��Qg�2�/�u��2YV�wDO��+�.!�h�;}��~� n4.`�"�]��F��-%��dB���������R�;)��2�����NqX4d�����+~]�|�n`�>hC|�����#�r�X�O�.)$@6M��p�EJ������M�)~��gʄ�Tō���}������9���ғ}��{������:�!��g*�����4��<����>�,���ƦHP�b��G��(I?����7�5�ִ;	$�}�b!���g�^���I�`�[�i�7i�8v��_�t��t)8�����nN��xQ��������&�R}D�n��ل��P�{���8�ϝמiNq|��Ҧ�|Ӂ�+�cz'a*��,Ęp�\g�~�`u[GCd;��,wj7�{Z����Hņ%�Ӊ�үx�U��U �`�_G��ߕyH�ʝ�1'S��H�_��'6�0���g�B�]�Ο˗k"�S&~lR6l����o/p�E�œN�S�Y'yi��B����}y�cɍ���	���fEK��!c	���,m*�E�I������P��L��c0��M|y/p��k��~�.�X�7��c��	���2o����uݜs�,l}U�u��t �)l��kD��Rl�\}�l�zG��oI�+5W�\�5d���p��O�n��gّDS[]{�h[5ț�� t���T����2��:Z}T=i���yf�]��'8�XlW�`�{���͢���#My�?W�>�͢DW����nY�.�'�����%�K�KGLOt�KҢ,W4{���L{�T �Z��k=+T��0g̺깄T
��Ոb���B�:�9�(m����4�dqapc+����0@w7u�� ^33��Y��*�=��r"'���	c��NDF�z��.Zv���w���pŤϔѯ�{�mۨZj��UmG�Q}*4��_����G.�.́!O�s������V�wq 2y�
Mwz�����"x�[��k
�$�sJN�cz˫,�FQ���2w�I��T��J}������IW3����� ��ЅH>�Q����3�#�z�㡄V�Q�kP6������rAaߊk|�Yq���]#��P�KȨ��qC���8��΄iT�I'�ȟ�~�m�8�qm�*#�G���,^�C��w4�|�$�3�f���]�h �����œv�}sq��7�8ng�i���K"_.�!����v��M��1�sj���(y�i�n	�0&��,:��+�U����IqU`��M�d�����ŏ[s�><"�v�	�Id#��(�9Q#tS��3��tDn���s�E�b�ۻ�]�Z3$7ϱ��>%d!LrW��TX�R��"�`P�N��=.�e�U�;�_��)XJ��!6B����� dL�g��t�I�k^n�.6��o�g��%���4T�x���*dr���k�-(�)���$��^T�XZg�m�s.G�Ў�'hoBi�Xm��0�I�t�M�w��.�^&��q��7)G���P~��" .�s�U�"����Vw����c�;��Nv�_�Q���1�f.�Z����e8�HӶz���y�2��[H��T�kRֶ�\�r������"hG��7�x�9�h��K���W�@�~Y�3������JY�3#�bom�n�K�dy�k�*3�=�� �.�S{�'o��T�4/oa}�(�s���1�F������F�1����G�(?��+�&e����ˏ��@�)�Ż� Y�χ�����D���(%'���ZO����(*Ma�(|��@�Y�1ᚌ�Pd:���P��ּ6 M[V��H�q�����|�9�������w�M��; �	�Df3�S)�8�(���</j���Zo�,.�VW�?�_���p5���6A����~:�FW���%�cf�'�,&ޡ�+K͇��4KpD�q?�#�,a��'m��f?o�tV�����%���&���K�L[F-TSO�֞ҿ,!�ӊ'U:A����d�+ݶ�-�������'(���Q����������4���4�	�������N�&ɍ�MU�[(�D����Ôm��A�2	�h{~H��Տ��^�$"�9�!���)��!(�"�>]����~����f�(I�����y��b�+c�S��n+@��%�3�o����	�d�_�Ħ������X����!1"�:�F���<ޒ�q<�*j�8 #
V\nrW��P۱O9�r���qЏ�>�@Z̡���t��މ��H�f���>e���]N���~u��BT��*td�0�9.��z��;#���ӥk�]��ya�F��	�ur��fW��|�,F3͈+CP�f.[��jdg����ɛ�b�I���j�K��c�-�P-Ee��W�|L_e^���M���ij�`�~�+nm������5�ח���.oI��YE�H����i�V�s�rt��N�w�r���?�!��ۍw�MR����LKs���F��4QS��U_U��"d��,��c�fhb����k�)�yL�,���B$ˀ�@"o�Nh�Y�|&N��RӶ��٭�!�*���/���EF�/�mH�K-"1M�:�� uj�V�o�^��(�IIBr��]��%-Z1�Q�]��B�b&S���uc�2l���u��n�0К(bʉKR#p �T�	1Ě������f�h�	^����)��am#J/�_��[�S9��t
fWi�Б'�0`���I�<��^�<��m�0zrl��*���=+4�r�����.%S��P)Gx�
�4��|,)K�᧠\<�u��m�3ڟ)�Q��jڕ��& ����R�;��.� �6���qGRcc�8�G�W/� #���QbD1]�7�}�n�!�ԅ7�����"�fi�_����rQ4!0��^�N�2��K��������񌾦����i��&N�p2Rr��R�#�V� �#4�R�� �O˷k���`��>{!?i={>���:Psun���g	T���%��{�Y�}�ܙ�m
'q��'����,"�]ݿ�"�^Zt�1�3��V��Y3�FrC7!UhBaFn��?�"��������1����'�X�dj��k��N�);�1w6J��"�)Ƕ}�K�_�A���F����R�m�X;�O�;�t�®H}&�Z��-v_����=���g�V\ܱ�'��_�׮F�	���e:�dr4�I���=��]�i��
��F����?O�+��3�=L7�Uylbi�>Wbi<������aP�P5�Ы��[�o�]&ͣ�3nƺ%��s�H�#Wm�_��v;�߃�Q���vn�T�o=�*��ȍq�L��kf��@HoF�@��_s���XI"Z!$��s�����<�P��a�K{s_s�u�'m�ooTTWC	�~�n��P�#�M�j�v<�Iq�'l����$�Qɓ`t�����(�-���R���Ta����!/.��\�2.��~0��q�a�yj@)w�Rk^���Y'X��W}�ۮA3�9t���7<y`�ZL4J�e����#��/B,��ZW���{Xx�,&c1����;cS� t������A	7	��u�Q��&M�!�����ή���a�#�l���[��cKW�Ss.���;A���0��{U��������͉������!�Z##B�h�y�G��R��۹~�l����Im��9��$,�i{62T��[������X�������DP���RV }��R�&�)��	�x��=@O�u��
b�f��u�Eo �[��,�K�ܽ�4N���p'�|�s��&�G�K7L]Q��¤��yxӋ�ӟQcX<��d�7e�"��S������/4'��_x="���\8d�'��N:P�\ۮU~���
;�@bE��H-��}4�x�8������=ao�l6Ƽ�p)�G��
�/Ͳ�pk�^$�f��7��Dq��>A��"}a9FA�/qjT��9��-:�����8��xGc<0�&�X�2lU�0� �������x��ɣ�y��	�閁�\C���Ǫo︧cd�z(���Hv���r�c�
�R�T,`?���B6L�w3��L;b���ir�|�ۧ�hp�B�Ԅ���G�?��2��т:v�WQ�T���QX� ��`8D�pD*p�����O�m*�}�lu�O�D^��)>��#��;��������a��݆�D��`.�`��/����eD�ѭF9ĕ��J�-���a�{rW�X����+�$�:f��j ��k&�=�#cx�s־<��B�^O��E��R-�u押�<�PZߋOTqy
X���`���-�s]��=�_�;�M�����;F�B�Q�W�h�V8D�ʂG����?��7#v�<��d@�y��Y-J�OTu����:��*y�ʜr���R���hQ��Z:c��Wx�|�^�����XmaaO*V{��^\�H��ʵ�2>�/��;Wy6"�..m[El��Ui��W#RF��.�=<XP�/*��- LI�kV7���Z�MCJ�� ��I=���"Պ!��_&���IwA�wGI�#8.�=��h�F���wqX&�їQ�Ya�g�@%��k39E�cn;%x��]p��5��&�$R���ǇO�����Հn�����[�Tj���v�UER�W�M�O�>��9-/p��"L��W�y�[K��{E�:���Y��_"w�7.?_�m �XJ�Ŋ��uY-�ƒ4sn��ց��F���Qp/���
�ʇ��2*�`z�������Ҷ�]t��S��ց]fO�DL�����{��J1�3?��]{��d�V N�N�3��])�t$��dF��.���܋�d�=d]�Tq��]��:�%!�}�]�'DX8��f�m��p^Y*�yq�#��mҪB+�n��-�Np�RV�J��-e�ye�������nm�5|u?1�f�S�t��4x>>o�{j�����{�|�M�qꉖ���Mr��>3��n��t��F��N�FIYF�����V>PL��3����O%�GӅ�Z�T�o��>/W"+�KK��z���]xqr��KiO8�C	�Br�V�Jynfͣ/<�Ow0�������g��8�	�
ɜݸl����m�S�"E�t�(:(5y5 ��;8����)�rl�4V,�1Z_�	V�� ėfs����k�����O@g+<�b �w��0/����6���d�Z3���.�qM���F0�6�{a���$Ե�M֠�v�u�4������BM!��0AtM�B���#וu܃"�\�)��q7_���	?�s�W7ac�r���2h�/�RT���s!���| :��!0.�eį��O?���?ЋB�����6�q��\�F�3@p�p��dU�C�Ā�-�sOomp����daE�5�d �5�����[�,R��7lC?�+��Inʬ�w��{��0�ZW�������0)�6���cx����x������i��j�@����M�����@i��n_0�2��-�w����1�e
�s,�=�G�jȋ��Ҍ�FuA���B��G~�ͮ��Mz�ɫ��M=��TA'�g����F��c�r��IB-jҦ$K��]5�
$�@z�%�UO��6(���_�qmv�{� 5�^J�#����~'�4|�jV"�ٯS5�W��:��H{ð:I@V�B���LlN�#�e{Qc�����گ{J��O�h��=@LuN@ۇ�m�Z��=��8���������|����E����Pl��$���3���bGiñxS�q��+bM����h����I��G��C�w��b���@v}@Y�x��4V|�:2�G�ex�Y�/�L���Q����]lH�ྍ���8�e�2!C��O��e����W����)1��R�HUq��D���2�O�ar_�N�,��o�}�+m*i��\TH���qs����S[����J�de�iUZ7���5̛�g?#K�����T�y+:��%S���]�[�/*��	 *�!vy�٣�Q�JV+^�i�N��b�w��D�-t1�-&t1g]G�P�-v=�th8!T&�䙫�)��
�W�yD2)^�:�$���b���Ԥ3مg�gΆD��^I�(�Xkzy�2]�+�f;��O��O>`l��(�Š у���^�䡵��G"!3��R�J���P��4T�8�l}v���tlD�hD�ޖ�re}�4�NQ�j٣:�!���۹\J���C�4���M����qx�Ķ>I����2}�?�`��P�t�-�(+b�dYO�y�!�j̇����Bs�:ѧ��o	a�$�	h��r�RX�������*h�m�����_Y���L���y}�a����Q��c��{9��i��]�H8Kz�ۇ�ۭji�7T
t��oU��BӦ?�Wǋ�4�C�8'B�5Zj�H���4�����;�&�} ���Z�\��m����ܯ�U�t�%	�k#Q��u��G-D(\��v,�/�a�W���_��2�%�4������=ʰZ;�J{�����}�n����E�Dy.�4K�r�p���Rz�_�}� �x��M:?|��¢� fKMAԙ>��+����E9'���7�>�#|
, �6�[� ��Cc����9���-�1�Y��V>��&�D��D����$!�I^@���D�g�r�D:^S�f�\5�GG�e>~�����T1j]S�(ho��E�a��!�)-�J��Y��E�z���\�6&*k	��'�}}������e<������&t��rp��J���U@aGݾ�n]�]X(�L�J�8�+-�z"���N��)_�ĬO�2�F��R#HC�9�/�ׯ�u����^g��H
���s9n�;�o{�yD���Eq�k�";������Z��ai��מ]��&�t	�u��[o@���鄊hMG����$fޑd�f��/��j����d!�U�L97�㙪f�7������<,���\����?�3�;������H9�b+�}A3iM�U]�Ԕ����L����O�,��2a�0�CH[G���_�D�"x1�R��m���4U�X�}F?�B����2@T	�o�A�� X�7��/y�tU��a�+ı��L-BK���<���g������t�/^�?�3��� �TQ�"�.8��:Ƽ��%�i�]O|ү�*��@����(N�%�q/�s���#[��ڞ�V]b�iUߔ�!�I1O�mh�ŕw�1Ej��Ӧ3Ƚllk�3%&#URh�;�ɝޅ8�w{�.i�<C�p��S^�NDa��o}-���~!�X��`�q�T�ت���hy�C��;������T�� PS���%�G�o[Q%��]�^��Hڳ�� ��F_���q2����۬�"Q�3톸��5����Z�Ia���Dx��?�m.iM+�z������ɔ
���իd?������).Q 
�*�����ۍ(�����]|T?�Sw�ǹ��$�8��Ϩ���Y���~�ߏi8���F������iP�U�-��*K�qw�懔ڠ��f8�7��{���@	�a\����9Y���������Z!� ���ڝ9ŀY���<�\ǿ�ĵ��9~hnI�<� ����-�0���A�hh/�ſM�;�Sc;�V36-Kpu)���gtf}B�#YJ�y�=��5�z�/����{o��9h	e�R�����-f�Xo�(�E�������8���s�J6�)~[^�@{��L�k�b��_ͪ8�ŋگ][�D~��4��� �fT�����o��U@��-?AW7{�da��!������N~l^�N��u��f޵�H�4+p:�镣$�!Cer��D�&���F�E�H� �8���M�8�5�cH\���{؂�bFǵǳ"7��#7�������k*�s�x� }:�E�H�2H�/�F�^������,GWU���؎�E�\��r��|o�Zg��k�A�ĚJ�
�Z���쌝ZCH�Q�� ml7SnP:��«尓3��5:(��n1�&�T�qg�n�������*���?�0�[�����T�3����G�2ըĝ��W���9�]��F��pam�^�$5�9�԰6�r
�������ˤ/z����C���3�Y
��m"���<���̙���'�����D-�|���k�
mXվ��cF�ڳ6\)j��A|�	WaU"I���IvZ,��$���XV�+5�B��<R_B�U4�t��&�zP�GȾwP�\�q����$4��Y��3�6v~!�BC�כ�ݺ_TF��[�ƾj�٬��Y��v �,;�s/g��ߖ��c�9]�%L��y^�XO�9�,�MNRw!��C�A+Q�T~}���X�|�d	�Z��<�˦x ����u�jrŏ��`�HOx%����ZU��:�����(*Dh��v]v,�I��;FF�=|>�W�[L(܀��(Y�ʎ�I�~��/<���� �G��B-S�: sg���z7A�^���s����r]`���qKFb�#���� �*�hY�+�U�\P�5��;el��Ci�2��&���m���G֕;ly�Fj��.aj����6p�At/��MҘ��>�%�zWv�qC��q�b�wsiJ��,�Φ��Hf�"�\r:ҥ��:RN�g�K@�p�e�M���W5"��4D�`8A�;b�SB?��ws�CWi|uU�O�C���ך�ù��H�N�����.���=����  ��J��|���̜a�n�}�|:�0�����K\x��.��($
l:*��^�j��w��A��K��C���?,P-:���Nbr�^O�i��u�$y���TWk$  �������z#��Oh��Q��; ݅��	z�#Ƨ
���b�Ϗ��$�g��殝�L���$��H�Y��Crb���Pv19���- X={�d80xv�[�~jӄ��T�0r�|��F/&���E�AƉ!A#U/���Q�E�I��� z`q��yY�E�\ҋ+U���i�lNH�<60	._øs���Cl���|5�Y\���Mld�Mf�`\D��- ���]߈�`�ɦ����W�ķ�N�O�k���LY�|m�Jl� �#��N4�,����v~�n��e?�=�4����r�������%��M�.������7���m݁���WT�_��c���lUz�4m#ⴺ�v����4���^�'�{�/��$��TBN�
p�5��}96�4G��럓�V���\��D�}t�W�G
f��WYF�~�23�G�	�	5�����>ES�����@Ki-us�-f�X��[�:n��� nYV��%��j��o7�l 4����V	��6v��8 .��$����Gmq�lzަ�!\N�`Fͻ������Q�6����s�J�Kl���J��iA��z!LzC����1�] �̚�Q_]KL`:2"��Kcm?���jF����s�M���f��)����^7e�T���1����#K�[�	�#�žs7~Eɉ���|��R�^���$�FF��c�+�1R^hn��?�z��e0P�1;�{��]t7�Kq3����u9�}���(�\��������Ё:}v�/m�ڡ��bl?	�n�xe�J@��*��ȟ��=@w`d�[���Ǯ�X;��23��;L����(�&!]���1Vh�:�ɰ�{�	a�o*�Q�!��D�T�3@�D�T����t;L2!0�:H/s.	�d���j�dZ��������<mٰ��Z	st�#�.UaJ>d0��m�"s�v���8n�M��M��ڪ������1�׭/;��r���s�?XP{]��j�>����e�
�5��_��.;�B~�����mf��1岰yL�������~b,�\���&�<�#h���C�'N3+��X&�˪�ɐ�ލ�\;e�kF��p�I�l;jF<�����#��G}�Kz����'��;��C\/=�O��h���Ğ,����g�N�b_jO9ΔB!j�g+3X d��P����D���C������ǜ�����q���a�	��Z���c�^�X���EE�'���ӢWG��tD�o�~�Í`)9ww�cէz#���v����Wo��B�A5������tE�f��s�Y���4H��>R��8@�)��k ��EIgA�5^s��k
H7�܎�@��Ϧ�P�5�rKbp: tݘ�ӑb�Ե�k	A`��N��(Ŋ�����$�Q3�hȰ#��.بTF�7�^x)~�j�BZ��r��oKu <���� *(B %�*����@��(�o�+I��"�>4&�>��%M��( ,��v�����_��|g��)��q+���3��ڒ�����(~����Զ�Nrn���˖�W��؛w_����lv��rj��J�{�D<�z\�#x�UjL2��M��My�v#J0}M"8�2B��q�4s\�*/���Q	�ԑr�� �0�ؐ������X��V&tBс�Wck�!����0���ע��C��\�Q4h���@"��=��������IQ;�PIZ� �٤W�3̷��!p�|?��(�-(�$.����7���,l_�I�N��.4��=.�L2�]/�����v[Jc�3�=SO)t�e�0s�AhWq��]r���:�N�w��9��ʂ�:ӻn+�<[��#xB��{���y���z���m{���������ؓ��	�.;�O��ʥ�Z očAi���֢(��|�ʡ U"��fiH�#�C˕���MlA�f(�w�R1�y��=E
~�sBf�"�;�4Q��� �(�ʚ7�fz�J��;
1t��\B{��lx������Fp ��ߔ�6�m_�?�?�%�qo�?�̇�9;�Ɍ8oZ;h�(e����c�U������*lx� �^Q��O~C&'׳���p�L)�n#e'M��E0�K�h1~.�ƛ"��:Y�K0@�p��{��B?)�Ε�8�z�)e�ˇ�pg1��\ҧ�,0q5�a�$��f�(�@���x��4��,|R�V35ߦ����;	"23��8��s�M2�wϚ����=&x�I2�2+e[kdMN�S�'b���(�V���3&�,a�x��z�ɣ��[\�Rh�M3��f�^S#���]RZ��S����3dWeR��N�k!(

Ƙe��R���(cy���LMn��فp9�^���ῴ�����V�[!�~E��V��4.��C�<��S9��B ?a��G@幢�w�J��|���f�?�_wnJ�5���+�nU��z��Pׂ��#���1���=�QS\�X�m�������΀������p{��(��TȻq;B��l����r����&�D��0"�� ���ׅ����g�obu�t� UX�qh'pkx&R�J�dGȥ�w��m�����Au�54܁aa�2�U-� +�����}���u=�Q���֡���Ӄ�v�S;��)�����D*-9��f�E?����_#3�'���V�QUĝ,����i��:�E^f��Kۮ��! ,�ɉ�Q�M���O�h�Cc��q �d���f� [�N[t�����g6�Yq��m38i>��d	�Ƨq���`�t. ���<�^� xvk���۹���հ�8놹��4���/���v�R˻D�T���q���W���D*�u��Ye�&��&��PQmK'G�4�?c�6���\ ;��̟�\dڊ�9��)�Ԁ�p��z���e�P��1H6!����v��O���QJ��S�p��"�(���������-��)܂������iYE�/���̕`��J;�"��x�ey�{�*e��{�g�gy�	s�}����61��~�Œ�\�w����
2H$v%�XeIN�pw�o��
�d�%�omr Mt0u)�������e�
�]�i���6��[������uH�n�ek��ܐ�"��Ix���~��}�^#%{���]5J|Y(.�eL�*uaR'�E�f)�@%!�`2�@e5�~�cba���OLyC?���e}}�{�Hԋ�6-�G��?s�;�Ai���,������1���T��-�SU���e�*Bx1���~�����rg|v�O�%�zFݰ?��^4��������ٷ��[vϱ{���d-����N�?����xL��p�f{�9S�]sY^���<�������	,kg�^�Y����:h8B �f�� �秎6���ȹ&,հ���0����F��j���+d�I|��Z�ה��l�VdtY��.�2��]�����~�`��7u��~:�S||d�S�h�"���Q|j�Ys��;�D�ޛk���8%\A�l=9�w��'Ώ)Mi�X]�c�n(?�o�U��&
���&�0�q-�-:�R�S�7P-`�WZ��"�����^���}��>P�N"���РJ�Z0��;���厫�j� ��
R�aI��|%D�ˠ[z�ߎcc�KR�Gx{�&�n}�K�A&�H
�&G���m$ˏ�F�ӟ]��iO����ߡ�E=G¦��n��P���vhJN�^���|%�cnMW�iK/�i4�d��
�22�6P~0����Xh�5�s��F�L��H�0e9��<PLR*o�k��R�@��c�I�
��	�������ܶE���/�:B�>IYm%
�������e<�Kv�b���J��f�4gN�Y���f�H�+�ˈ��B�����Ru�0?��F���ol(O�_�@�u���� ڝ䌆�fa~���O�"�Jo>����7l�K�ߊҳo�Ȏ+�,�
��_�_w�q;T4o��-Uv#�iÄ��'�x3H`g&E���`��ڏ���M�;���n�v �R'�X���:E.n���w�̑ﳘB���.���m��í��b������o[Pvm<?־�$3�ԅD�����l�uv�r$��`��\U� v��3Z�����"�/,��}�z�Z?�Xۉ��q������/���;��w�N��tҳz-�"��
�2.^��t���{�!G)�JB��7��b��7��h�skMz��t��S#���݋��D!&�>.�b�{�
��Z㑮�k#�d��}�� [�eWW���~�x�tWԂ��>X��-�?Fs���p��n�h�ÄqO���$o�J k%��`���?��+����APmp'|<��#{�+2u���ւ_E��/+@}p�E3'y�$V"����L�	}����=X���5&��	�@U�B�N�_�~�6�ln��^v>� ���$D�6% !O�@Ԩ�������>�C��2��z�T%�����s��9�5%�P�?�'}���*�R~�d���Q��%���o&�6z�%�K�䨬�6����Q�#Ɓ�<�^�q���~�����r����7_w;�Ř�#�f���)p�����̐/A-	���Ǿ*�w�}���Z�e���6�|l�[�W"����[^cr`�*�k�x3��)a�ē�f��uZ
Y�W���ϐ�*l����m�����}(%�d��&ʟfx0�jӧ2R���C�-=Sz1�3�K�`l��+�{�Z6�pt��M:�j��QF�d�~R۳�ş `�vå��-Q���}���a�d�q�%35L��cJ+-v��C��!�g+ߪB|{e�T�!��wՃu�y���o�dzA�G���LL��CC�
��ySk���r4Q}�"��a��]�����"��S�{rW�;<i�};|[XZ\�ۊ�pϳ �QGg�4��.=2M��I荒�
,7:mb૎|�[/.�2ގ9��c<�7ţ�� F���Է�R_Y���-q�[���� ѫ��qr��[#����]ZzbaP�����2�VcZ�e�pF�;��]a�5vm�R�S�D��˲D,�>M\�����$%�9�컍r���]��k�h����֠�\d锼O�(ŏ�:�Ǖ�_KV�(�/�TY!����yL�D<o�}�:E����T��|Y?���@���	Z��kC���͍�m��G�,f�"����
)3	�A�N��.jyo���ńˑ'M�X���3��~�Z�R�ڔut�P�q��>�0�l�k3�R��"��C��&b��k�%�ɵ:�S�Y�΅�ߘ��
��<j0tM�����+�ު���A�3��b��6ѹH��(�3��S�yԒ3G�����ɼF�Xh�lO˶�T'5��:X̯��@�l*C����h
Qu���L�'e]X]a֚誊�Dz3)����"���^ɪ ]ǣ�޶>L�����o��v��h��h�����3Yr���u��2���6����W�����R�An@0�%�f�>�X�fɡU+��5	��t����I�<�ά4��OBy�B=��(~FkռB�{U�L3n9&���(w�$�	�w��a��}��4�r��~�Z�0'ш�����y_GM����'�P4`��O`��b��� 2��+v���{xT�;W�Q�g�>��)�Tn��� �y�v4����~�����MfvA_���I��ւZj�mȬ�f�2����pK��^�S�w���ݽ���R%		�ӕ�UkT�o�׿mZZ]k_4o�1���m������p�9mm$/�N��cI�}���8�[�p�#�5T��jm���[LV��	�BM�����b*��c �D�G��Z,[���A�٥DJ��٣M��-'@������q�-�܉P|i�������6b�n{����ni!�\��<4'\Q'-�I�-CCP�/�%�7��,v�(���J.�h$K[�t.րXNWA!�K���Ug��`��̹x�m��W�AX��w��Q���;�WD�f�#���9�Ωx̌��M�ŀ��4g�*��)�{Z���K�����R$D�F"��R�K$1�jK��N�e����I���h���4��A�\��Cꦼ!�e���ha&cS���&r�N��|Sr�k�VQ���������vc���j��ȏ����1Dά2p&8�??�]��>GI�_%�"����c�G�w}��Fs��W��h���@<�gb7�λ�DB�Sx�>*��!����P���
�!7wdN[_ULYȰ��nc�kc[���E�(�JGK��y�����[�.�N��^9�p��T�t����Z����^��a&<��iz�cU�V��9�)�z[e�.�=�+���dNq3U(�J��]{?�����( A��i$�^d�bjujB�?C>�����:�� 8w�Y�M�<d�d2�A�����;�%OՔ��7��q���<,;f�Y6�țv�px������ė8#��+�Է׮���d�*�s��߇�QY��@2X���p�?)�"5Sϖ%9�z]������`�r��%k�|zL;��rX��S�^ܚ�Ju�a(x&�o�(�Tɚ�O|(#<�m{G
�[�|�:�o.�^;�4AFM�-�⟃É�u�&��1��y� ��H<o�r����_	����k�7�뮷�!���\��Y =Q��G������x�ߘӮ��3l�u��ҹ���?J��;e��V����D|:��Dņu|��y��r���t<+�{���d�T�U����!�kQ&��ЊB9�n�	�v�LF��rs�b��*��%O[�vuK�鬗믯H���>.5�����Y鉶�����eU*��qv�!�FB�A���0E����(י_�E�� ��ε&qe��L�1�SL�F2���h �Y�zVZZ'�K-r�pUgVQ���R�\�*�c��xQL������-S���P�9�׷K���d6��Ji DmsG��2�B�5�h� :��[q#�W̩�x^(J�c����)&�2�KS>��X�+�N�*o^ǻ�,p��&�x��ؚ=��셂u�0������a����+��K�?�L�?���a�퉗x�Kh^[���`�g?�H���?�̴?`�)P����͐�\�uSUs'�k�_f�'�ƺ�ܬZn�Xz����8@�:䬌� ו�(�8�Gj�W�\�7�[��3fР{͔IN��Ӑ��U��r�HCP3�p��5�z>r�U8]�3)c�^�ߨ�r5�: .�����k�F�YX7����Ą���YLSbv�_��<��QT��M}��2����Wӗ<R�l/�|G�jMc�D�9�/^ <�A�֢�>�^.���ԝ��2�T���-�ڲ�ۻ�U�ъ� F�^��2�Z J��8 >T@(���jWdMg�H%�����G#l���u��.�(p|���~l�D��h נ@��7�)�51�`"i���˗oű�oz�W	�!-�:'�zB$�X�O�X`�^?�!-��O1�#a�L���i�Z�G�A��d�{��P���:	-ʇ��?,a@�����W���&Q_�l[A+,��q:)%�!���B!��"�1�E��Q��
�VLp��5h2�;q"�o�/s/*�(W#J���*Z<�����:1�8�2��)puLz����9�j&ת���㧄�s�$�`�HB�3����͌f��[k=,����-d����K��
Y�;���\����Gq�t�ڱ���_�G&F/5���z6)�Fy2	�^/S�Gv��ѣ���)R���F/�J=��I�s �m=v�!(A>$�om��8���`�]�q�jA�7������R��4MP���T���[>��D��B������k�>��a�0�r!��_��@��ڦ�>�QC��k������^O�.���<Tk�D.(�X(>wĹ�d�$�#�ҝH/�lVI��]nN�y����S�X�Y ϫq�5�D�JC��^S[��u&�ț�3y�5φ�(�u�#��bW|i���.���*����&��桶��C��0�J�K�J.�#�|-mK^-���lu���GCo�'�0�@��F2�@�֋k���A��s��FRO}xV�;��}�ҩ;�S�r���v{n�IY��h�F�~�Ӡ�X
�d��V��SP��Nd[�lP���F�����fM[�wv�����$R�R��a�)��i�e�T1/� }"]�6!�2�X3=�B��
�)�,�����\-�uՑE�^�`V!��ٍ$��K�%�v��Z�J�����LU[;��I��|����yQ�1�B���e@����1�~�.Le���ݷ���畀KjI�Hj��-�E�<>ƴ�M��?@�<f*@�wL��k��a��y��_��PH����%� �Ҩ�͑ ��^LS4��/(���g�-�Ѭ(��<%���t�>�	�"'�ZɄ�c@��"�D2�͛�aug��VTB�̫ h��/
{�Y�S��I~o� ��Q(dAj��6��u2��Wlێu�)��~�9����z�:�s����xZ/c�ɧ
�l.{|�B	�/�.`��J6�f�~����;9k��i�_B����n�ڊ{$�	DEK�dF�DU5k�)��#��M"~���e�����F��|��l��P�jPSݭA���m��C=�/>,٦4�F�9����:(R�}+	$&�W!�t��ǫǢj_��m��4�5 C�B�����E��
�)^rì�mr"lz�N��c*n��F�1��9�}�r^�8��ddeUy���PP<���33�%{�LP��=mNhH��U[�k~�(�Y����n�S�3ꥦ��j�K[Z��я�/�����𕴟{��uS����E&-�i:
���=4iT޸[a<H��w]�q�Jec�2f�n)���6��J�	�L��V.� �/�^��6�����݈G�D���BP�8Q���h��*=-G4vB}-:��N߶�~G��=Ǆ�o���{���@RUtWe9�ݹ���M�DD�w�j�����>�l��#b�O
o���i@�'�S+Y��_�c�3?�
�|0��9���hCc��_��G��$N�,�З���J��Z��V/,�Uk�=U��J�{��8T�� �����F|�>���VK���;5��[�{V*��1�Ư�I�U �XE��+0ߛ@�t7�3� ��t����KJN�POn�ШaF`�*P�8����<R,c[�Q:WF��B��zt�O�T[A�N�DS
e�x����#�ߢ�W�1DJ�ˁ��L� ��lC����4qV�z�{:���C���_7p�3���y@�OY�/����%d����BY�7��-�y���$�$��!�sx�H=��
�p������pڽV���l<�Z,�#L}ҍ�?t�vRC|}9ir#�F���o��s�@��FtOcF�����e>�fk��=�?���xw0�6���]�9�k��	lC�sK"<���ՇT����3�vH���F��B�W��w��b7�b��.6O�	u�}���#9�ݩ�$u���Zu3퐄OVc���l:�g�(�~�Rz��c�]n�W�=f�U߹�ƶќ�� O}����XZG��þ
x�)��n{!U����� ��6{\�������o�ܓV+$	+���H�u�IA�5�lԁq�:��q��(��L���Q{���}�� b�=��#D�<�ewhN�'L4Z�J�t�)�� 
������"����dꁚ��V��L�)Ȅ��s���k��&�M�e5�r�Qɤa[g��,��S�WQ�D������G4�ˢO�;I�Ig�F�e�,��:팦�k���(��d��h�����gx�3��Eu����������§��"wU�I����R���%S�Y��fbO�QbBY��'^��YF_Z;@8��������\�5�1���8xb��h�n�������q��-E1 4�W��d�[eA�Z&�j�,D����ZN�>"�k~�k���[g�Ɲ�n��Ĕc�w���L�=�6m���F��M�O�>��R�� �+u	<��6wְ,����DO��(l�חZ�zS�̲�~X�Z�$�"D�]��߀��ֹk=�i.�͔&��W�C���?��RvMK�'>{��'�GE�������%\��p3���ы��	�8!�(�w����p��O���ƒy��ŻF�S�~���ǚ�45���o\4�Q����%LO��i:��]�b.�I�]Hj�/����OW@h����;�yx- z�*�	/'��:԰�ے ���8�u��*�#H���c��n���6�O&�3����	����F����w4��:��D����z�.�Q��gDNS����q/�Tչi7�69���up�6����8���j["���!������*�\�*IlT�0e�y�cy�R�M0	��P�m�gT^� ˻�~
�b!�ɮ=���k�
��zy�Xͷ�Lh��G�g���c����n��rg��[�`&��@M]�-��c�U���$Uǂ�d�_IEh�=_cjU^PV�-��ѡ�LTE�e������hvl�¾�XσCK5V��w��ZׂٳA��ݘW�ӄ���w#��.�WWr�ߧu����45�n)6�>�9��$�gL�A�A����C��"r��ms �����F�|����M6����y�Z�ب�n�\J��{\'=��mI�k�"� x�V�G����dֻ<h�J��©�$��(�L�:ֆ��\����RK+������З~"�����$�ن��+�^��4K�i�JH��@g/��R;��u�p���E[+�ꩧ�u���gU%��ԍ�4�~�l��EMi��kz�
�-R1>í�{�I��01|25��%{ȫ$!Y+E��������T��U�7"�J�aS����H�dV���3����
�Է��'�q���J'�!�J9
|z�:L�Àk`�� ���ٚZ��0���"�����и��y��~1��(�OS�����rE;l�z��{��BWi��Z�va�"�moެ���/B�ꪽP䝚h]��R(��(�wp����0ꇆ�
n+����1���V߲q}΁�G9��_Z�r�ۧ��{����*ǃ�40;�g%&0��!
T����v�S�������VC�U�&F�ɗ��'��gPd�1�l��o��N��7���b��:�~�WIf�S��~߼�y�=��x��Αw����฾����pZ�.M��5�X�[R��b��:��2nJ�c{f%fMK�,B�ޅh�P6�%"l���MWD�Y����2P�S2�am���^�g�4����B8R���ǆ�I@��_��_N���~k��tMJN����!��!��$w&d��J�6�v���֢�q�����hh�� ө��0o���z�q�і~��j�t�8�M[3�.�O�TS�\B)��K�)�Yi��@w�,j������5���# S�R�ݝh����۬M�ֻ�o� ,���3��<8|bQ��X'�g��F�����g���[�	5
o�K������IU{�*��x0.��|U��
� ׏���o����[�Չ?S�y\��\[и[�
Ю�6r�B@���z���J���A�#�r���y�f���o�iots��"r.�`F������D���#�=� �z9��(�H8G9�v�[�kSo��?(W�����1���(��#�'ԡMc�q�$�FSx�G���3���rP��^\M��Xr���.	���GXA ��#GQ)A��:of�Rliv#��9�{��V�gb�T������-���7" �q0Ew�+��5�v�ҹ��]�gJ��&�X�6U���G�j=/����&$�]a��O��������풳oS����Lz���ݚ�1�oyu��`UX� "V�/�v��
$M�L��Xihs��i�5�Y��y��葞�,CI_XԾ��[pT�3��/`0�Ф0mD?Z�C�hLr��K�UJi*U翢��*����*ţ�F;v�Wi�!Z`��m%+�� y��l3�B8g�O����|�-)����HH�SV��5��"��;��.I��{�G�I~��z�f��8&nx�W�T��U(V�NBMn��b�x�ަ������͇8L5r5;jO޿�<�ZΖ��<�#��ل��_L��A�����ҁ ,E�qڶ�4̓�%��ܜ^>��v7}�di`#b�֐E���e`���6�����P�t�l��f�|���=�F@����l��k{�;��>"�e��>[F��l�����2�A1��V������Ͱ~�=�9ZH���{.���35JK >/S�� N���k��:�tܬ�Lid�1��	��� *��DM"���YE؄�z��3�#���z?��%�>ˣ)v���[��
b�?9>Q>��}Y�����&���ґC���hj�������ɬG��x��*,\-���β��h�C~p��R6�<���
r
˨\]Vᑺ?\�c�|�O��?<��E���h�a�a̢n%��K�,=z�S�a;;=Iƪ����6r��o-�8-�f�U�7��d���_�YTH�;��FNI���ҁ!qeh����_m��X��� ����۔�K�s+Njd�Uʑ���
��Mi�� T��J�?�Mw&�S�:M_Wǃ14���|��=�CO�fY`LUŀZma��=�W;�l?nT��PJB�0���|�@��</ì��>i)2S�"�Ŧ"�!=<��^ID3ya��~s@P?]��u���JŦ*��_*�T�D*����T��o�K�N�$�8�=�h�?����`tn?����/��b��ZuYhctM�7[�"uO��׏������պ(jG�-�΂�=��e��~�C�k�?�h��a&�|��ˀ�2���m2��;
_���(�z+�U��w����g� -l����G�Q�5��0� ���W��ْ.ʜ��5\���2;�&�Z������/3�t؞9���c��Q�&����LX��p��!�ZN��۴wױ�/I܈�������Ra,��hca��A�X��$�c��Cٲ^�KR���f��׏"��z��=�,;<:�����