��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{Ns�ȭ��+{do�;��F�0�Sa�K!�f� b�|o�Qy��\��ºQ20�[ '�����u���y�K��<r&x���\�X�{?�X-u�~2���J�:	>@Z��A7$���d���Q��+��?�+�yJ����~S�����l�"��е���}�-v�F�G*������{|�ʒ}���Ӷ�c�1e���<*��pA�I�o��B:2>�v[�F挸F��-�T��a/�.�7'%^�um=�n�\��i�fx���!�_j�[�fbb��Jң3������/hm�
��u�/>}7n�W�Nd�%DCCm~���lh��?Q��ԬC�
�BX� �c{w;GʹBi��|��P@/,n^�b��}��F@Fw��4���UIK]`�vp+��n����(���6���sݵ�@7{>�nQ&��/�0+�n���)��eW�<)
��2V��:��c%��i#6����<�yo��4�����;߅�ve�;BzurloWTL;���/����Uv��Y�L�q��zԬ��Vϣ��4t��º���
�GV�`����R	�8����p.�H�"3Fm��ꐢ�kwj�@���b'��~���,�hH��E�ǉ�d��}0�T���00#�cA� Ϧ�&t_�3d������|>s�?��`C���gH}'�o/���6������hq�^�d/����-ÎR��T�õ8��3�,����`��shX�����y3�	�&L�m�ͤ;�h��dǛSm`o�.�ƌK���u�{�؃URj'���toQW�Du���.��Ix �����Gn���rb-���i�I��4�<q�je.�dv���UR%�����P�QRY8����oǙ�)f\����̣��#�R��@o[`'���s?<��~� k5Ȇ�g���%�'���Z߰Cb��{����8�|�s7�������8бisxt�$!#���=��OT�B�~�\����Q�PI���͞J_���
$,n��0N�+�JA,Ȇ�d'�%�
���ӵK��8�*Kzn)n��pƓS�����  NZ�/� ���E߯��!���(���۱"#�qgF����j�����ټ��,�{��}十�4�@��_o�G��̆�A�C��n���V޷�6��.�IY�;�^��3���=����B4���s�YUA�@!
!�=��Ol	�<$P��ɤ����x<���=DXԯ$!��O!�0�����8z[�A�5 ���n� �HE���b�������|F$����6>�8�r\����~�5�}u~k4=� ���Ob�J��]y���!8JX����r���;A�����WЌ�?��z+'-���s쇌m�X�Q��H�ɐe�����n�u���m���a�=�{�k�26)� ��2>A��AΘ�)V؞Ű�'z�,>{�5A��(\Z��[4����1�[i 0zA��1P���P�%��!�2Z~���D����l
�g-p^����?���]���#?�,K"~�"KݩG+A��^p��`�r��!��=n����Mo���lz�4q<n�>':e�3ѝJ�I	��F�z{;o���)&�h��<���I� ��L`�/Gp��P���U��� ���b8�Y�lPy�.���q(�� ����-A���L;&	��6�G�C�6�_Gb�e�g³G����f����u����4�/�-�|O�udʆ�'RS*O�������D�1�*a"��h�9�L����P��pX�Y2���NU����i��	�w��6�`��m�m:	����U��*�I��j3ύƎA͂<&�B³�<�H%)~g�%�ՂӈA*�ZȺۈ��^�	�����}��R����<��m��a�#���PMy;y�Po�F���*�DTC���8�!����8Ŀ�(ل�
�X=�,(��ڤ%ܼ]����r�c։�v����j�~�g�gTO�ʠn���u�u�q�Fsc�0Ф0�)��|bj���k.���
��pl#��GW��2��R������R;(c�m�r��	�a�]U0�lLF�.2��|>e��^U���П܃���\�&�^�X�h�,R����vظ��q��5˰��e�����7*̵9 ���Z���kz� ����cYl�H�]�����T