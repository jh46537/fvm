��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���tǐ-a�Z��e�l+�H�uW�Љ��Lk�p�@}5�[o�Hݤ|����j�{38��/qlW04\h"��=7P��2.��[��,~�����d���4�o��3%��!�:���&��G�Q5FJ���H�(�m���G	.��I�I�_���]�r(1��k��0��h�&��b��j�����Ǘ�g6Ԥ�f��*��9dS�>}᝟�i�C�C�����Ó�����RǬ�]�BU�����po7(gP�ݴrsе�7�V���~'�u�=��Y��<�(�;?}��Q2_�����-N6�R;SK8�n#1�d��0R*h%]6@�Kp� #�|�S�nj�C���� ,`�T��m7��O볻�ʗ���lUw�{�\�����pL����@��pEkR։��h�����,�Bf}'}'zM�����b"y}i�1ʤ}|#~
dSK���l �ԡə�����-~�+�*
.�;�����",J���g���|���P�����G�:*�:_��fNah��%�߂v��9X��Ϙ��� 6���gx��o��
f�x��^&N~Z� ��4�Yw���~����O>�y��C�ۭ1/�H0b��U��xM�C���.�AD[�ď~�Y>

����4H��zfq�o���as.)PD�3�Z!�fr~�� .	b��J��{
�b����.���	
�:/�t#G�F����S��G�z�@��rQ���g�D�ɓh�q�j�&)[	Ҵ7;"?��	kX2�!<�e�O�-HR���f�S�,��П�g�2qҼZn�s��w�]���#�-x8º��yc��R(��E��-!�U�%M�lO���~�Xr/3y��glK*�gW���9��|}��c���(JPkG��Sώ���q����@�:��"�T���G�"��7�dk���ǎ���=�n��-`����<�)��W`X�#�%��(�:1IU�Ř�V�4'�B:�5�n�vJ�G�Ӿ��Mb(��&`����Zx�]b���"WJ�v�l�:Cl�"��udN?�	����S���Z���)�3�O�<�S3 ?&�r����@qu���nS�P~�+��u\���Pݕ���3b0�%�2� ��q�kƕx�6�{xQ�D����ʄ[E��b��i��|Ι	;��>�4Ds s>H���mQ���B�D��jמ+~�/;Pj�>G�,�H��P��ӄ�����D�!F��H��jCB��DxWs��P�Mͥ4���iZFŸY�|���ׄ�qvG�4��Es(=ő��6������SC;�i��$GE��Q�A�Y��c�h�u���5Q�䂹%�4C���FgϘ�V���s��2�>�+a��؛����S�V�:�ܶ�z2�x�N:��k�Yd]�`e���6t���7�9=���>�}r��:7��'�H��Ms��w����־��d�븥����ŭ�j��C?�u(��D���� �>΀Ad܊5H��B�1O{iH.�H�&�&����>MFo��9%���K��gr���W6��&>
�X�/Q=R���D�����I��������&��D�]��5^덫SL{�_�ۓ&�_����F0 ����.K(����ݶ���������K�-��`��'��n�`fΤ���$���a�7|�;I2q|��N�~ٹ�����%$rr��6>����nt����ܾQ������]>�h��"���?_V�.>��X��X2\:f���E�>���촒!a��Q5�� ṘK��^l�R`B��}ѯp{��fS���ђ��УL���mn���6��<��zW(��}UHx>UO;���~�A���5ubl|׊�U��*�P����
��a`�;o-Ec�W%>���K��q�����D7o��N&�>��c<�*�$I�`�l�-�@1���>���/D#�����S�._rF�h"�����w_���|���C*�~����JXir�f%�n2��$@��zv]��d����=v@&��%��WX�s��b�p3�k�`|���j�).f��;��RC׆K�	��N1��������>�uyZ>�{�4���c3N�{h�g"01�:ﭮ�k�-@�?�Ƈ��1C�������-�,��:�Yu���"C$0��%�W���.(�l�>��a+K�|�ﮘouK���A�owd!ݝ���g*����jD�=�i���O���=EHf�oYh)�dH���G��� =�x�0=GR�$��'x�w���_�n��f%yl鳃���)�b9������ wy7�0n˜"<�jQ��� >�;Uy��|��9���'�gIF�㭂,�#֘�����2�=q߯ŕY�@�i���0?E.é�r�%C�x�'аw��5X�#��L�����8S�z@>�טf�"ީ�U_��H
���iY9��ج���\p����~��p�:^���Nu����!7R��n�'h3CI�LQ�L��m�*�(t{Msi���=${Ub��)�����-y'��m�+�l��{~^��V������O/S[���o#Ρ/F�u�9�H&����i�V�#(DS�~˃�-`����c�Qʫf���_�,F��	��}L��R�q#�!;@�_^��%�Ү}Wo�d��"M r6�l�"�q���j��ղDF�3�Hҏ��(�\y���~�ű��E�ʸ˞@�%%�A��J҆�U#h���e�iZ���<�p�P�����z��㍩V~��l�yx�H��^��+�)6uo�r!�/��*G��{��h�O���'��WHX$3�<qQ��	`��e _�2���L�8)@�� �Q��1�)H;^�w%
Vf�ؕ�Dh_��p��֚ H�50C�x���)�bgĎ
�s(�.�N���i�����舼)�����4�"�|_�[��k\���"��0�a��m�91x�C�c�T�Wx�G��Su=��&�r�h�w��ÇZsW�1Ϩ�0	mJ���o������o�������K�6�6�]��S:��*���X�Z��8�~�B�#���m�&�@�8�ԒZ�������Lg%>B�&�վ�����Q�-M�t$��AЉe�zq,W%��g��ӨvH﷒�Z�9�O�)�� �;(���ݍ��"s=���h�����J=F��;/�[�#�@��P�)���v0D���D�U/�틌�I
2$s0j[&>�&��=���!x��N�b�{p#��@����?�QL{�������f��;@����WOG�V������);�ƆW��A9����S����Z���!zQ�ȥ�O,�kd��J��3d�d���$�y[�K�<�1.㩷��Ê�TH�S�h����5��;��~$I�nO�.��k4rL������ܚ`F3e$@�F��k�tŮ�.���qY�l�P�3�h؃f:~�e{��\��g9dByf���)��W��<����N�g�9o���8A�FY�ߴ�t!�Ujj,1ӝ��(��(6Jv�y�:2���Q���C�7]���ǯ}�\�m����'���e����m�ŧ�G��kX|!��nt�����I��0*@��(���ݮ9Ԩ�H)L�k��˪�^Y/�������S�Fh~��:TK��J��΢UӸr�f�h�-���8�*���6ݷR�K��oc|!�[��x�{�����\m#G:'L�<T��<�`mM��O��~�p�s"3���Q����/orZ��݄���7����|/�P�/�f�+E��L�P:�dK���S���/M^�[Y���$����WaJR���U8;%S(�T�^��ǜ�#�����l.�
"\*�I�Z���?�oP�E�EW���jX^u�֏s��pg�y?o�ߜ���z���R�g����9]��bdK�6A�|�*�7��1~@��3�������i�
�0�+I���c)3ã�dZr<kT�����4�|�2��NQ����Oikv���?ᰴ3z�Pa�R�U�L�;���e��{�#oS-�4����b"+�V�d�+������qd��C�<�����Q^���:+�P(�,��&����1E�J����t�TvU�����ώ�|zL��awr�AN���I:n��U�����b�2��LS+g� 7��t�q���:}ܿ��`�γΡO���5�9�&��k�m;>�EY֥��+@	��]�A2s��&�\�4�U`p1ը��>��O�p$G���U~������^��+��i��&W,z�jl�e7�q
 5��<ސ�rE�-�8,5�����~�IIX�[TNV�M��_�u�2��H���ùg�,�->��B�ͮ���#��6�`,a���j��;����v!�9K����Yl���P@+��Y�AH��7s6�X�X��t�4@��+;�yժ�FzW��{��p/��L�h�0z^ڴZ�K��sQ��xs�& >N����!�U�O�}��2^9ơY�#��`�5�S*oD6Á"�r<�'fָ�O?���)�mzq2�T=��{S�ecᱟ�!� 
�`9��l�ͬYk�!��dE�aWP�g����]�[f�LȻ��l�Z\{ڜ�1���� ��� ]�!ol�!gӜ��S�|���׫b��3�<���&����}z�`+n���2����`�P(M��Ĭ�v�lR$�`q�˕�`�.�ɐ�[,�yJ�_Ö:�.��d����5��#@+C����U��V� ����q�;��T�d������Ѧ�+�_!�Ac-�4:m���aQ��@��E��x��Y�M�l�q�`�ڝ_�F�a��:k�g�.G�_�Vǀ�B���� a�>5�/�_�R��aC��
SA�g�!�A�F�\+&��a��W��ێ�?��k���;;��n<�[H��:��+rcV8��.6I7�����E��ڻ�+��9��vv�5�w%�����?K,���e��9��ք>��˰�'���"56��|�
	]@v-1`���,N�_��d�vĒ����~3�� '�d^*͹,w`�*��Z��杓|D4�����(*>8��(s*֤e&<Lr�V����[���/���'��@duV=�i0 M� f��4���C���}��#E1��߇Y+�0�{��ۛ{����lW�gE��_7~i�L��������eЀ.�� �M�O(�{"9Ώ��Rؽ��H���E���H�E��s��YA-n���賬bƛ�ML�G�o�.�Q>q��2N=�\�rv��*��@�:��3.�]ux0E�gq|&q�ʋ2-�s�Dm��s V�������|.7���Mc���/]?�EZ��0�=�`������(�L]l!c 	>f����A��+ԫ���rv?��J������R�gѦKd�P�����x������=����-_U˄e���ı4ۜ7j��'>���5T�jG6)�&�6�>��="�Nus���खC�?�[�lT��I`AY��H�� �V���Y��l9��-��1�/���$.�i�^���_(���ﶣ�5TYMQ�>�I� 
U���ĠL�6��Z��J��q���a��Z-����d48C���p0�|����8�n��
2<1#a&���C�Ҹ/dI�4��]F���ذ�KiH `j�p3h�z�T�Y��/��.�2
Fh?w~��&������a���ă�ZL�YP��-3yCgVg�67�|"W�j�3������,�[-�2�5Pv��R��v���_��Er�Qu��_1�:�g�Z��nD��u߂r�����h�t�ɠ"t6���?0���24�����ߢ�e���Cb<߈E����2A����NF�F�_I���lAĀ�ʿDd'b�1�MZ�BF߹_�����I	bᷫ�֒�e�C&J�=�xTJk�� ��p [Q\Cv,	�g qB�(p��m*c����"��'CC�}@73xO��~Q��#���4�z����U��
W����6Mb�(a���%uXd�Y�%Iw�G/���i3�����v���x<��]L̊Ǫ���7t슫�D3&�	��گ<7�;�t��Ng�(� o�Q�d�Fߜ�T�m)�4�����s������H'� E):k�|�<��׹~���hv��eYd�5�f���R��׮W��&��\u։�D�mh��?;D��>�X'�*���o}��u�`�(��o�奆���ؔ��t�@��@0$m"'���E��� �]��,[.�?��"x�Jk5���vN���Yǁ���#ǥ���؀B�^N�r�ǝ�m@å1ȢW"$e������H�\��ĥ?P�y���fɄ�<y�;��]��DԎO����;��](Ԉ�}�A�Yaͬ&��L!��F7gc��8�৉�g�Ʌ��mWH�N�W�հ[۶cCsB?�J��R��p��%P$~�r�������Z�VT�z۝]%�P�s��@��+�Δ�V�R���+��<�*�r�r�o��v��oHu��+�騀�F�O�ͻX����^z�4�7f���jr�\D�����d_rfP,�=����_ݲZ(�*)7�=�Ur���Df-�֮�L
������Fy-�W�[�Ԝ}�v2�T!�cI3uM?ܝ�N{�	�V'�|�5J�qIޣ���"�M���[�[��d�'y��6��[+bZ�EY �K	c�q�օ��?�K�sQ3�~���{�q&A�d�0}E�h%���J䴱�-�>��-���F$���հ��a}�.��&�{*��V�AkXe�U�'�V�!<�ZDR���v#7[�d2�3ӟ�+�.�X�k�%Sc�^<�fqf o,J{�YS�i}z���(�9o�&7��/�	s�7�%�:f����p��/6��o���i�u˄"�!Xl�nr�Y��脪�^�~��=��N
�<�F���T�L��L��-D(>O:������R���,�0�<�iVD{�z�1��J�sF��������9�����!X�ǅV���);8����BT�>S1"�[=����pA��N(玻���x�.�g��O�>xA�+��H�9����%(w�Oe�qho�m\�Ha����P,R�_X�z���r�KVx+\ht�g|{%+i��0�a�����6Ҏ�Z�DP�ʽ�<����)��&�Y��=�ǃ��=�dԃR�5��"�z�Ӿ`+�2�>Q4�/��p�b�M��]�vR-���g���`�Z��E��'�g��Q� �c��p�H�x�
/��*6*+�H��/CZJ��_���2w�����sW���2�y�o��:� �8O-B�~Ow��x$�����GZr�m褘Y��ط���g���nb]�^��:H���Ԩ,*%;(�N&�sm݄�Q�z�/�+����XY
}�6-�[�d�
	�g �|N��>>�ճ
�t�{�Wȸ"Sǡf�bW�s�Dt}A�ܡ�)�}����EHBԑ�7.�� �5���s����?/U�=�)��8��Mztŝ6;R�	0#͇`+�����Cxȫ���� �+��ݴZ#�u
6q��m�w]��IEg|.��	�i��U��Ǵ�Bg����I�l2�c�,����.X4��B�=Wa��d���l��Ѻ2$����՗zo��+�[2�ͽl��qlK[��(ͩ� z&V���rrۮ�-bɐȷ���K����V��p�fRɌ�/��dz��b�(� �z4�<�:,_Uj��t���DV��X�&C�/��a�n��-��A1�t�A�/�t��JǶ}\�����\�e�('_(�
T�{�Q�("r�O�,��7�7U�N�$�C<#�R���pҢ!R7T�����=��3wp�k���Et~r�LJ(�NvF���+�q���}�;l�+�
�$��eA��UIh�J�[�D%ھK���֞��B���� �����P�1�=*=ǥ��@���y �z�_ՈKt�C�_�)G	��Cz�@?���tiH
���z�+�����VbV�M�6��	==��zl�����x��?����v�;�|X���1�����6�LX��Tx��i��::{r	i��8���(pl:�.�Ї��E�髳Sʠw����k`�_��^��?v =��⫗+3���#�ߪ��p��c°���	/�:q��>�d=��Y5�*�����k"0��ο�~���-��50�o�	ݞH���s[9��g���[�h�TB��0&T���Ҿh�@JA���}��tmeD[��J��1J��塝nd Y���1��f��o���Ɓ]�]b����6�KIS�5/�Ϛ�sF	Ŏ�����5Ǔ���b=��=���]0��7@�͖?�&Rڊ�����uŏ�\�˭����<�5�E���2Y٬���.�p�S�
J[XeZ�Kɸ�hН!"�?�Y7%�P�t������@2�����]<�v�8s>p��<x9��e�G0S�^[����%��lN�[{�(�=�x;�1�+#�=/�g|�����pͤ��'H�t�p��/�yX�\��/���]T��=Tk�Qa\����`��?���/r�0s�~�a��L�G��Z!���G�Wԩ4l�RJ�YF�� X�Ո�����̜Tmd2�砫�$��Tq�)�%	��Sk`��?w��矶�5su{���eI��A�3�h�5q=�ilo�2Ӑ.6k��8��Y<���M��	� ��cx�&�WB(��2��:7��;$8Gڅ؛F�ƈ��U7Pw��ŷ�!aq=�u�G���}�S/�H�*;zד3߰�*��H�h>��؞����½��Yc�A��+�c�U�@E�؍*��ޛ=����˚�+�Щ�ӂ.(C�e�e)l�&��@�E�B�[�b�4 ��Qu�w�S��r�����Ҵ�5��o>����û!�TG=��¸%|3���"cZR?�<�"��T�ʙ	�`q�#>��ո2�uȐ�6�(�7#�Q�_Iޒ���������.<;����ʋ��K�F�f�}ʨgJ>
�1`�GQ����ܧ���8�v2��hY�˰+�1��b�:�d2���� K�*:"���#1�����X��zRKm���@#��<��З1��Ü0zBZ��jyb,H2��j6�ޔ���Xw��ĩn�5�I�1#�I�Fzv��¸y��TYG��ۑ�<+]����nD�� J#�����t��S�O�X�@�}@^t�	��Qki��h�kz�^������Y%6|3Q�ZHO��� �3�_4�����0�f�B�ٸ�"]5����я�� ��;���L��Y������H@/x�9�D����gvTd~%cmp�~G�?²2rFGv�T3����&R���iyƤ0 d�b�żp��ے�+�����xP7RD4����vf��epTIx���l�诸s��=P���@���q.�����% *	C��u����,������>.�=t�h�.���&��.��x[;Ɉ��}`��&�Fn�I��O�4�����P�<f��v�R�t�p�\ba2(`#�[x(�8��@$|>����em�C��� ��-�GO5���o�x3H��V9>��*�I���dp��2TǕ�
�}�M~���.���؎k�ꖴn��s���S��X!_ˈ�4��$B8gF�8� �RB�Lל��c�d�7	!5��i��rE];� �t�!�g�� �Q�d �֨%�А��j��oV0��\y����	�M�����8�D:���4����ʣ�Lb��ٌ\.���Iu�d��B�T�8�C�D���7܁����y'���~�U���xf�;iؽ�"�x��n��� �\��z.�e�
���%�d$�:G�����9��s4q-��y�	����{�9�y]]>�9ʥ�w<@��Z uR���fpH�W�m*Ϭ�	cK��@9�~�Mv���m$�E� �&۵}��� �����`�ɢ�O"�d<��PV�MN�2��h�!kbL������u�ΜH�����2�FK�u�o�W�lX�>$z{�^�,��IH	�y1���$/>ч.��2����*rw^��W�>ԗ/��=�Y>�9.a���%o�����3v��G���v;�=%keȅ��i<�\�����˿Z��3����ʜ�d\�J�v}�Qr3��I��mN	��d�o��Ӱ0�f�1-����R�7�;����Q�+���5�����/���-�RDH�mZ�cuJ\ݓ��f�l��ifgiǁ�C�<%�O�l.���x:7�v:I@���"�j\T�0���WY�J��d�"����\���X�$i�xQ��(�S�7{�Hk�/� ����6,�Ԓ\$�� ό�U�RFj��i���|��%[�"��5�G*:��2Vᨳ9gN~���;b��)�s,@�9٧��D0d���M$�"B9��"H:OS�9�d����{҅�T8�T`(~PO[�!Rlڿ7�w�a�C%m%���H�v#m��x�F`�r��d��Bxj?i1lb�U��P�.�+�?~tzN�B�M�$�Ǩ��W}@�ק��ו ���n˛O���#�v�э.��ѡ8��0��V��Wx��	LyX���1��Q�q�X�lu,>�a9mϚ���X*���ÏX,Aa�O�Գ&E�qY�oX�!���!�,i�w�'fw��<�Q�����O5�����D��R��QM��!c_"���f!g ��y�O	M�צ�n�xz���� �7���0\�gjؙ�Eˠ������V#��M����A$�dI�$�w�H~)�,~qP7�I��ҕ}���$���Ѯ��E���θ\����t3����d��nGP*f+�E%�c3|������e����b74ڷ}�D/�tqT1��*������&V��;�u��N$�D���Ќ�|p��Ƣm��Bn�CvS�c7T@����H8��7X^��$>��L�UK�+��a��=��OA֡k�_�JUYk�v�V�z�U�W+?1@Θ����`�r�iCgv���_����vI�h��3WZ�����o�"G|QI�	LӘ|�:����hj,�Z�u�Aҹdc��A�)���^d�!~|B)e��7U��������2R��0f+H��H0e%���I�|F�2E�{��ױ�=��z$F�,j�>�8u��7�8�Dc}F��9���P����,��'���T3�$[m�JT��u$!�,(4z|�E��FN�^s�-��+RKʟ�t�a�$B�>��].L�����ʚ�Kb�g!��˗����`� ���bխ�����!���/�?ok|"� ���a��QU2',v���L��Sđ�.��;����8��M��]!z*z�F��Q#SIX���S��Ĳ�_FW��7�,=���/_�G՝&�m^���MAw���qZY�$:�N��	8�I4�^�j����TM"
�W?�5Q����MQnm ۷��D��ҫ`�P[Na�S6�*l�r7��id�Q�67���g��xҒ����e���lͱ��"�oǋ��}�|�p�v��]��"$���ǯ��I����XQ)����Ǚ����J.z�=ˁ�Ya��p�F8���yPY�1�a�Y�,QA���uY����
�E(��0kaO�X_
U��) ����I�0g���~�c�L��I�c�(��8�ᅡ��/��w՞u���3V+Y ���Us��Q���a�I����������˚�-mMj������c4�;M�l�xXp�2��+ͦ�C%/��],�WO70�7sm
j�S�����ZZcڕdG��'Q�N̔S��c�Ʉ�9�"b~)�n_����@��ܱ��9���F���U�`�_2 a��M/����P�f�)�0�	�K����GI� �0���$,݁�;�jzg�=��Y�q]k�Gy״�����=������d�$��G�o�(A1h��(������6/,�$j�*{wA�����K/�Å�4�0�<�rq���}e;��aX� #�J{_�D��\j4\L�E��>jσ�h�uWn�D#�>&�_�	���b����m�^����m��Q*� w��wb�:Ch��Yr���r0��ͺ���H5<pGV�]����gj`d
�R� W)��&�8�.߯�`���q|�W�ß�r>�|uM�Io~�{?٫��,�36�5XB���	�T���~y�#r��)SH/9=} �sy��Һ�O�����D{O	u��g	�B:b���}'&��c�.c�p�ہ�)�m�9&���	�GN��W�10h[;S�S~�W�d�q�6����`h
]�5��Q[�� VQ:^�b���S�;i�U�Q�#���-f���[��Q�l\}�u�ib7k��p�����1��i$��S�O��A`G�[RSH���M2{��yeSgv�����on#�,�� *w����q7	��l`E�_�;����X΍���cd`�T[��fX��DgH�9">w׿�[XNH��$�z���E��ZV�N�2p5E�G����:�P�d��FK�\4Ġ^�]?��R��ކ��f��#X��4�K�H�U5�xJK��!^�����[�� B���쬹�Е�]���IG��牌 �7[dT���9�d���Oa)�չ6��X1��_�7�կ��&2�����nDę���-s/�\�iء��P�;Y�ml��ѫ:�) ��r��Q�n"˔����*�T,ս�~��O��u)�ڏ������<b�=���UD��aG8��g3�ߛ��S��Q܌��}�g�4��]���\��@N��0V1��8`$MM_�w�¬;�Ȯ�<���| ����
δȹC�~1��;�9���rl��@o(Ww�E�=��t�1��ڡ���e�@H��IX���!a�tbĔ�����gX[B���r�tKQcuxd�])����gR�$4�/�g���0����f�$8���d�:�� �ڠ�B����ț�C��h%��mj�]������"�K����nr%�S�J����4��p�ᖁ�Z�����ۣ�֮�t���\�|���I���jq���꥟�sW�T����
�чS��y���rׯlq�r�-�*笍Η�R[Ԉ1��y��&�h2�ί���y�yH?3ۿ��v�剤�Z��������_@Ig�F��_���h�x�m�������l�R����+�0�=`se�`j2�;	���dQ2�]�/ �r�ɏF.A2l�k�-�z����Iǋ�0˧��Sѕ��=R��[]���B�vJ�\��?��N_m��RĈ��F����" -�&��Wz�6"fG}ߎZ(p���^IL�J2Ԕ�� ��'I�^zW��{���fbI_/R�ݧcKҾ�B����V^J��-�,H8]����Henw�2�� �gnyB}]N6ی��	�4?�y�*��
Ug���d����L��ӶG���ˢ�B��<�C�pp�c��x��[�g��L�Xh�;��o^��8��ÞgF��9@��(]Ds�N�Rٝ�N��['(������b����<�U^x	br<_y�[��㱴��WW��#x�N��]EA0u�_�nMK�
ZH �x�C�Tŀ�+�9�	/�\�Z��͵$���xA���F	�N?���3KHD�U�yS�C_%m�J&l�[�F���6ꥌ��Q�i���K/�Xr�`���������z,X�[Eb���&�,�tS� nD�+�5�{GŌ��uӕ�qr_��d(��=���iפ�G�5���#�;>�m�M�u�g���g���i�	�.�μk[(/&�t^��,�y�Y+�A=R�/3�A��t]Ó��U/��|�K�]�V��?�bH_�S`�LM��H T�ex��%Ի��B*�d�&�s��;V�Pd�á���N�G���~�a6�`}F0���v�:��"��IG���%{�H��"���眖�D�P���a������I����D�IU��o��`�V#nC8�C�7�Ԙ��|�Z�1q��W
c�pI����R)�ވG�1
č����y����e�98�rOa�Iy&�1�y[m�ps޶_��	��:�d>�_ȋ�Z���BM(U� ��wj-*��N���v���`Y�HZѨ�\`_�Qf��W�4Ԍq�c{��%I6��[&�t��ܼh��Y�B�#��FN�s�.s���f��j]�L���K^M8�K ��Є��A��mX��0��|i��f��M��'�@S�7u�c	A\{�	T�e'6�S������w��q��g׀ ��ǝѧ$A"r�����L�����/O��y�능8�����`�>�.u��P��w�|[�ݫB��{�E�6R�6�Cr?Ur���|�R��S�Խ�s��0\Y(�"-�&�U��u�aH,mw���m�f'e�����xB0���'��\.S�s�W�L�&}�f�.
�:
�B���V
�I�����i���.󠐏�8B'�9I�c�]�$v�Q2 ����E�l�bz��܏�</��x�)�����r,_F$
V�S��k����ç�.���T���u�� ��6�/�U��w
�7ㆫ��GY�6Q��6,+^ӊ��	h:��^�{ {ז���&�	�@�}
� V�>׳�/��F�`w������+�|��LS֖������.F��@�D�j.&It�e�=u24�nK��a'�����:�z��U�\�i���x�׬�T�'�qN2�۝nZj�D��0�[r��b�"F��r�/f��4m����gJ�콽Y趱Gd5�� ��+ ��G:1���UN�`J���]r��R/��Ԩ`�� ��;�]PT��|t'T*�O'袥��	�ʹ�|\q[�§v��PײԅTj3��HƲEs7\͇�tћ��6*֬���v���
�޴L)Lώ�4kR�c�X-0���-NQ�r�oe�Vk:��Vз}|-֛����>�ZV5䌢9b�8�^��O�.�$]dcC����?)� !٫?.���k�h�ެC��TH�|I0Z}�,e6�+vv��3���^��8�v�?��Z�U��kFt�$e� �C�R�Swj�׿C�we0x�o���ȱ��-Ggö�!�~�(��t�`�������|�c�K�\�c��"�-W4��$C��� �~*.��w���udJ�ˍ�L�`u��@�K�O�QK@�7��[�Ϛ<�Ku�k��~� �g�,�ԍL�R�a���֠<M���n�\�d��s�L��P��8s,�Ε��Y%��'|dS�,�H0<\n����d�ZBW��1��[�J�`��z�Ґ����g>FV��qtp��W��n�l���:u;�Ri���N�Z<�UT��Z"�H�TTn}��qHlf(���n����?��IW_��#>�M2��3�5��A�jI+v����@e��<�_4�E������+�`m<��r�ܞ�j�7L�9Y�!�J�9GY���۶�%�ǹ-!��hE��F�ٌ�@�9�ш ��ѩ�"���]$�;4������&?���՟"ڵd��~�(q���ʡ}�A%�%�E-�X�e�w$0nV	�=�$x6ئ����,$z�}Lv�T%��M�|��[}�e_[��Wt C�)2�N3�.�Г�8X��� \�J�|A܀a���O]��+���/2U+�x�!�~N$g��Mr������H��t��BMD���׈=Δ�ʽ'���W�\��	�� PG�
a���-� ~M�@���=�����L�V�����Ul����� Y��q��ٵm��f���~�r8J��ӥ�vh��S��Ӭ!��|(��/J�W�jBr"��T�=H_ێ3�|
�k�S�W��`�`������O�R#��X�&��� �6����􏔄�	�J,ړq�!�ϓ�)��[�i�H q�M	�p[KVg�m���5]�k��9u��c�5�>�:�V����a���}GVs_ձ�ԫ�x�������MN����;�,~�U ���/b��i8�/u��C���u֬V�o�1��WӅ}/����T��y0;t,�E��:�s3tl���F�K`�Q3��V��7��c�ȝ�"���OZ����%֩���4F��S9�߈�9��|�geQw�������! 7�M�?��y��Z��f�]ș$���2�Lŧ�(���pt��s���	'�3�(�ƽ�'�y�+����$��Zz2jT���J����t�Nl�4�!��V�].�w���	��b�Z�S}������� F,6�掟r�?u��l�Z��V��#T����I��*T��w�B��EuVxd��l�՞(˞�s��&(�=��Ǵ
����5�_.R�϶F	H�>"�@�������N�7��3��p�]�&�²>w �ޕ���v������R�w�	�6��MY8W��WfC��55H�#r&�B=2���H���^�DH�K�������!t��B���lh�\� t�"lEWt7i$�%�����a�o�R������ljS5y��y���6ȣ9U?�0_w`r�i��սPQ��~�,�����JC��A�#�'{c(�1AΓG���iZ��A�BE4&!��+���SfC�ߗ1�#�j�]y �@:��)+�3`T����f�Ҹ��1��]ZR�)��b{�>;�&��d�!%����6%ߘ&qJ=��n"芗�ڌW�Q�=����LȒЛ����I�/��v�N����3"�/�
�t�Bg���t%�m:�+T�y�w�y�זq�鋋���-�����K�HRL�R���A+eه�%���6W�P,AB��%6��E�1��|C�Ԁ�?�*�U֞����6��Y��/ȏg"_Em;Ǉh���ljH�L�\�f�_�}�%l�ZN��I�t'��,��T�!�PF�i_�������D�]�}=riR.�Xك#��I^?<�p���&�=���j+��o�V9騿��C���̔S���Ӯ.�䚩n�+.��+�~yNM(@IU1�������@�T�H�`y�kW�䪨�{I�M2�A^�����z��f�\ n���)�En�4�1�Ka$��0��֤�y|�8x��1T�4�L_�?���VAm�Ҹ@q�z���{Q�P���~$/�-U���3��ջ��G�O�F7��r�V�	a9ߙW�2g�[����a	'���b�砨|��!AhR$T4-m�|���jй!R��ra-���rwn�j��p�R��7��,� �����g �H�ᷛ�/��׆���\��V��2%���gf~�j�Z��:1�'�2����-)%c���bMd��ʣ��:i����uK�.+�ІԤX><T;�(�E�Ρ�������'[��Z�dw��yՎs�T�d"��_���44�2YB3a�w����l�l�`� �}��|n};P-���\���h���-l��+ݰ.���������,lNgG���XSͯ�-���Ї�|�� ����?�z�2+� �� ��ѧ�/B͞��pV�x�2_*�>0��s#e��t̩��IL�6���*w[Ϸ�YK����
A���N� �"��-\fIO�
?\������hڝ����,*Ʌ�Յ�Z�ɿN]:#�W����M��q�̗��3��8�� k�]�l#�o?'���hTH����t��H��661�Hcj?�k�ZFT�����'�"P}�H�2v��wkE����;X�����]�Y7u�S�ۿJȱj�7��y��5��.�?[��ϭ�,/'����ȽD���ӟ4b���[�
�Q�lzW��x�٫����,ȣc3�nA���#��L�)�q|e�lmL�Q�-"0�<�.�h���"�_���WTy,�{A��O��uI�߬�ici�,?�����x%M&�q�lYu�6ģ;�~}b��_T�	���{���Y]�>t�-��U�M4�s~7f��(�ˬ��������{g͸��s������J����{���[3� ��u��*9�`P�����!�g��dl�,��Y��^BU�\/�9I�:���r\Q�!�۪�	ø�5%��C2$u�И��kN�� 3�N
��� ����F��A�\M���m�lKu�@ĸtHhJe���!��ƿ�4��������7���:i�wΔ���D��E�7��c<���awqr���#<�KV�y��}f��UqOUf�����?YS�u�����Cxޱ9Nҵ��V��f��{;/�ƒ���o��xta�H��4'G����}�����B'� �8[��t���
�A��*A�nBP��c���/�ӊ^פ��؀�0N�� )-�;:i��{YQס��1���<���QkҞ@M���whW�'A|��,��be��>��Y��l�
������%�b�����:@"lj���������f�JYi,3���d�����=�+���l^,��4:LH��F#��TU�^R�RR_u��H/=��`�^���5UY�,M�~��;�)�1���5��.`��5XU�Jh����G���g
��ЕYF�}�D��x���	8a"�;��z\���S�����Vk���I0j#��?����9qZ�)����>��~�⨤�J�X�Ǒ�A0�=�M!�S"xp���b�E����Ĩ���r�R�̥�!�z�E��D���a���-��}�V��/!r�X��z��!�ud Ҋ�4��n�'q�O���4�M/\��!C�����, �dj4��^pA&����U��2_De"��q�tǔ��a���P���>J��F
�����?�N���L ��l/��l�[Gj��������&A�h�(|�����ѯ���A�^�6��C�;-�ֺ	o���Hmvas��:
�CfQV�Rtŋ#Ъ��^�/%��v�H"����8����841	U�K�Nb	��/�9D���s��O��r�V �`�O�.̹���F!�B	k�#��� ��G��00�ׯ�9ߜQE�=,R&�w���4�T_!�t[7�Ȧ�{P�0X#v��"P(o��o���UWY��@<Kt`�1d��%�-����4���ih2x=Ėr&�xQ���r�g	1�G�@#ǋZ�>��^ig�eA��Oq�����`裮ٔ��QT:5���%�a��!Uۏ+~ƥҘ�?��T�{��"LIX�y���d�m���� ʲ�oɇ�9�8�S�k�<�ѐu�W�K	����	QV��&��O�P��?�P3��cf	!�k�ǵ����'�FJ �9$����bCi2R�ڷ�=[�B�؊K8��}x���;���(����si���hniz�{��s�5X��D;�P]p�f��@�i�U�&#�Uf18!>(�^�0N��Q��ʳ�D���x��� �8�r�4%��@�T��ҳd��X����Y�3m ����6F.X�d:wsLMO����M�:�-5�����C��"U<��X`�T�l
�g�P����g���d�˽�`�g�a�2� 
�"|R���ׁ��Ѓ��6N��_������A�fmi���h�7�D�i��J#F!�~�0y8\�C���ނ�TtV'�(�&e����D�g	���X��H9������ȕ,���WF�t�J�.���K���+=(.�𓯆+;���
q��{VA�S(�Ƞ��h��I�i��@T�;��DJDT?J��Mt)�M�/�f��'�c(��X��Ji8�F�?���P�r|0�9�hS�ݎ܎��qtD�L�oKM���վ��A~�ݻuW���B��{��&8R�%�����I_K�L���ұ
��Ɵ�-�`E!oi�r+I�*D�b�k}�8�u_���n=A��&�mqq����m����U�l��<S�p���54j�F��m];�niCfe�w�t��8���Gҹ�s���<bpĀ{�ޘ2��I��D���r Q�Q-4��s#�Һ��v���A�yY��7
�*&怽a_=j{�zP�"���r���C�<8�����d\�c#�s���K{�%�z߁`N,*����LZ��|�`�ϖ�Ԝ�'�a�A�6�����F3���Z��������+��B�C����}f2�
bͨ��:��PY[=�	��S�?� T<�'�*���䆰��#�1q{��K~+��p�v��/�"�W+� ���`g������N�f������W�v�K9Z�n_�˔7IA�w*E�����IÚ�C׬Ta��<�*�{A�;�n�gV��lEZ
�{�=��Di:g�׭ �9����ͳ�Z� �|��&���%���W�<#.¼+ V
̳m�7�w�I6K�:%S�r[�9Z}�ع�rW�tXíD�I�t���%�fM{���,����+���I��u_&U���n����4���=�@�5���0�]�y���G�3-����5�
����Lf\s9���Z�1r�g���x���u]�m�Zˉ:sUi@
@���B��O��s	�[]E^�!^�\5ޚ�ѓX֮{�8�G�#����?qb.l�uE�s:/yd<����"ZkQч�$$��������q�W��"�hZLg��敁�1s!
y�|d���y3ųCL��K23�R�^n�+^'옹�%	�Z\�/cg��Xhf��b���,'l�e��$�R�����sv��a;�p�=��8���9=�Y��#�p��y���o��4?xcs.�WGf��_8 �r�D��{Jt��$WCo~@�B��Ğ�m5�
�/k*�㍭v��6 ���u�9}J5yR=��F;�wm�e���Bq6��#���}�"�h�Gʚ�D��[ć�����I���1�&�}&bS�%j*��]PE�E;��9`\	!�9�5�n�
���d��\����O�^V1�MA;�Z�I�Wߓ�Y�R�sA2�
唎���!cId��0'g�1�|Ͻ�5�m�b�þw'�he��X
iif�!DL��c;�>�ۣ�+�(MHy��׶�1�a��_�����`6:k*�/���E���4�.ˑ��D޷��{����w
������jD8F�6J֣k3�TH��#�uW�:M�޽���5�2��4��8Ȃ��ܦNAD�%�5���$H[����е�g{���J��,7\��8i�"]����H�'qۇdf�G

�5�J��y3������wZ����ٛ�g�3�b��%}Ո�:Ԙy�"�+��H"�v��DBw���z�К�{��X��P����Q/���ag�5D,bb�zj5�~�����M�n!��pX�ء��'Yɳ�j�D��
����Nh
6�}'f'�����j�)�N�e�y-;ӕvֿ�����p��[�,q�bA��$����
"P����ȣ�������TpA��c�<J�ʹJ-%��f���%-7,�l|�+9��
�}� xwV8c.Ѩ~%(OU?b�TvLr�M׸C� mt�W1[�7*�� �s��A:��i�"�M+���Pe~�-<��
��C�9a�,����ӕ1k�Mg�j���PDm$���pR��,I�Z����ך�;l�.u\���z� ز���X�th-Ӊq�&j_��+�8,�ۙ��3s�%�}4�2}F5�tH,��Fo09��A:����U3�9&�"Ru_���1S�5Z����1�JJ\��[���DǕ���I"s��z�=V�+z�	)���hݢ�~A�kG��ćݏY�W/D��D'J����y���~&���j2�ސ�`���*�5��T�<U�y�5�� �\��q�.�t?�q�5"k|?Z\�/ٺ�$*}��!T0��ݍV���C�M�c�!�*�Z]���sH���%v�>.����X&w�\�η4�.&�U7B�j������-C�s�'��$�nf�1)?�xx�\�-�ޓ"��h6񫈲'����������S8'b	�P�0W�T#%����p�1�g�h
�3��>nO:���1���@֐CR�Ud���-�|��4aa��>a3N
��3�4�6aJ��y ����P����x��׃&��{��*੤=8n���/󁄁o�7���� �SmP������i;�( H��R���67�Ng^-�臸�V[ ��W�QU�*�ݲ��e��O"�3��R�2�ȷ^����5Ԡ�j�̗�e�&�Jit��2]?z�3ѿR:0���(���*�����W믭��caѲJm&�.��������h0�X�����c@t:��=QV���E�o�)�kQL�1p ��£����֦4��X�E� ���l�q�8x���˪��{�E��-�@	�r�2VM֍ⳮ_�1�o�[�O�rv05�륽�u�v�X2Vb�PqP{@n'�L�~FI�s�Â_�u�E�y
����Qb�T��R�F����U��[W	
"-��˅� ��%�
bs��S$Xb4�h `s|y�1��b�!UJx�Z����N%]ZJ�����I�s�QiY���K��<j�e��}�ۣ��*N	M��<������+����:�ܻ���&�)�=G#�_�IL:'~?f����;@�6=̈[U�eL
������HЙ脨cn��X�Ñ�"��l�E�ј%�t����M<�:U
�X�W֥�Ci�#�ʹ�ЎH���[�^Z�0y~*u���ߨ��(����y1�jP�<7��X�L4��'N3��hӓ�2Ջ"8�vv�p7e��	�n���0s�S�ǨN��ʙV�ӽ�|���җ�/���`$�8��|O�p,T�t
�=�%փ�ߟH��(Um��m� T6I�Z��(�1�ƖW����9];l%�t#�`-�v�3���l�M�J�Rp�9��nh��c�A��!�סWXd�W�s��=�-Q0ė�*1o� ���؆�T8^[%�����`���o�M�U��BL�cE��������U�&p���@�9o1����k�{ ���ҝLB�#ً-́��OY�}֡�����0U��?9H��,@/�%�$S�eD�#�d�&H��%ˣ�"��
Z��7��T�rL�B�?B��,^�F�|��䲱C�+!��]x_�%i�Z*�������_�f�L�W4'6)���B��ȼ���L��s���EIĚ}I�P)�>#j���@UVo;����5`�@�®V��mJ�`]���1�aC~3�8���;���WS��̋ګ�E,��ͮ�ѐ�f�u�9��d�Q�����ݮ�w�0�J�K����0}���H`��^���FѦ��t7��wA���!��1~��ۼ�����Ҙ��s����JN�Af�{��WbO�Y�nA`tհ9ow��_�y^8������ps�8���W�a8�B��^��z#$��IbMKo��(�S~�:�2lfg���|����@�V�y6k��z���2�9������}��Pw@�O6 }���92A�������J6��?�5�������}��Ad����2t��Y�����P�*=��dm����ZL��{�n���[�t�w�^s��U�3���� y�H�;M� �Ac�^gȯ(e������@M���Ub�V�땓C��P�5۰W��PcZ�o*}~v�m�k2�@o�-��;�7]�1��ً�b/�i�"�Z�W+��N��e�����hƕRV����hp���|
'�&
��t�Z�+���Fkun���N7�A�έiCm�S0�7���y9�3d2��R~�N�C�|+���(Ą�۾�0I*)a��ѫ���z_���=O��,"�����S� �4-m�C�/������)���gq$�:�5��T��K3#[�/����m!���r�s���砚];nݽ����N_����L�C���mM�B�:�"TCL��/*2�N�@rgF�+,~�2s)s���8�����j~�|i��K��f9�k��p�L�K��Ja_��Y�tU���������;�'�W��@ؐ@�;qGr���3�P�gl�R|C9���Gǥ��Ks��BN5���^��%r��6+����s.LG4�xG�m�B�����(.l��R椪P�\��,>0&�f>ԃ����Vߌ[!L#J�/��w3�k���z���(s�P[��~����]�S���tʂ�F��u��R����kgޜ�8F�Qc��`���=�H��Q�c��GX(Ӌ�_�+l$��	���˫�|X���.o٥.����Y^�lO�
R���m�؉Do�4Ѻ������
��v�)��=�qo_��W�]9��؃��ʬ��^.oP1���0�G�Ʀ��;��xf^;��/���^�Ǯ���S�7��>���.W����C@�3����g�:�a4�X�s�8�*zE@�\sd�b#���r���Z�?T���ɯv�u������bUN[�E�]���b���i��ߝ������y��u�H6˰J�@9���2Q��1W��L�RH�fj�|'4*.C��$܏6��e;-C��A',�8�p���ex�F�m�ЬUDX�W�C\Z�z�˺�r�x��XI�zr���m#=u�"k���TL�'�'SHLN��)��d{I�]_i2!Lr�̰K����pk9�]ğSĨ�����u������a����Fh�=�Tv��M�ً���$9gf!����� $!�.,�7�(W���fC�zZ4��}.�M�'I��ۖ/�����n�U�uq�֛F ՠ�]�W 7q���+z۱JGe-�b�دdӎ�1�l���C������O�1Ge���]yY��ؼ�{�HQ��t�1T'WLa����o��a?1���k������I&Ȇ��9��I�m��rr��� ځ���/5���>������1�˷X�ވ�_�=J<����xJ�B VQp!�v���Q�[.5�9��������)4[t0�Q`�(L�Rz�����d��,M^���>c�˫q�))L��3X�gQ�]oіYV¥�E��4+���><*�!Y{�݇��.�:��R�#T>_l�G\0(n���-j�~��T�(��]_J��p�+ֺ�*bvΨ�_���>�ȐX sױ��ۊk5�9��!m�qC����
���)v�a��v�~����xX
�1$�h�-H�)I�7��2�&��!�S��]u����	4�IQd]��r����-���.����ׇ,c�Kω�c� �.�6��%���m��'M[L�%6����Ņ� �a�"�<�}�R���f�������U�{��+�ۗ!E�����6���JU����8QՊ��Xo�T������0o��XA��*>�⬢��\�'�35;D�o:���-M_ ?É�i݆󤨫'`� �贯 �`1�Zly�����R(�i \<��}��L{���|^�>��f�ʹ�~Fr������Nb\�7k^/0m�Xa��G��[K�|�1|D�b��-��9��p�]ZG���&->�k�p�ݠD���(�OْE'��dk';�]����Q�!rVv/N^��y�᲋�q���b�md�����D�g�~�4O�o��Sf��$�]O���e��V�䒲�����D��T����*�2l���#��|�&�'�FG�{����X�/Uω���Dʶ-fttF��
�<���_����J`:C�	�����ɒ�b�Q`=u���7���c�8�r�_���qFG3���c}���hb"��YM�:7C0+L�3�w*���zj�hZ������ g�&x�/F�U�Ph�4�D�	D5�A9�]�1���v/m��9�ig���]�ZX��Jvfj�?�S�}���[�\ 0
��"`��fHk'��ŷQ��u~������\��P�>3v~D���0�������H����H�8`�ρ-����e}��z�C֨3�T�_��M6��(��{d̘
�{T��BՓ��=l�<}�<��Z<E5#蒘	����lX��5�,���2��i�G��hei����c�dt�騞�J��e�V��	N�{x�$x�{5KX�*��B��z"Go�.}��E-4���S[�Ѡq��[)�����L�";�UA��F��᫔8�`�T�xH���u�Rn�?~���~`g�͕����#���	�tA���XY�HY�Y�X�[MAn9�>�� �N����Wb��]t�?؞>��r��{���J�J��.ya7Y�g�R���m�V�/E���N�|ww�K����J+d�mpm�$"V���F�~qk�ʧKY�ɩ��y�~�du��p��W�7�KbNG"v��0��M|3�]�C��he��Q�x����FZ-��:@�Bt�&	��l*�ҧ_��2.oc�9~+��}s�;�2&��Q��\)~~^�����C!%�3�t�@��ܹJ���aE��
����b~��5�}]����<�?�+��0�Ķ 1RY���z�=i��r���	ߨ�Ӑ��a\��@��-�H����Ehg� 텸b�Ɗ��Ҏŭ�܈���F�)âڪg��Ô�͔���r9H��D:B2�E��$���6�<������]%�p�+��MF~j4ءNWp���&y�����٠���#�G�u99���w-!I{F:+�O�űޱ��I�}/�e�!Z�z�0�r�aŹ����A?ªf[�9��o2a΃{�[��(�v�WՒ�y���yS�Ln�M�Cn\��Y�c�H}�<������DH=�a����>�C�����ˍ�$�� n|�%�}_�0�����S�L� ���M�7�me�����Y\-e���jz�*;h��a�����1x�l�)ү��8�����[�'~}l|q��z����G/+i��C���H%�����eB�j��u��GN�}*�'m~��·������9�?8޸L��A�Σ���%�>'�*΃��jg�
]���v��Ti���]!���hb�+���ǶS�5*$�'�Þ������q��"O��AW�>�\�u��b�K���ܭ�y89�"�@�(���/e:ݎQK@g Òp�1H���D�ǳ��\E �7��Y�������.�ӑ�9H��G��f���|m~]��N�icJ�:��]6nB����#[�M��}K�
|O�g���%66��6�H)��qZ��O�"��d=�� d�ȟY�'��CS�f~���X\Ԅ��V��[��Y�����K�0ȸ���TG�䩫�G`R�)@��u�(N�(��O�+2��	v�w�b2A��6�F��m�Aݲ���w�Rр��5��5��ۇx�>�����78��m�'ʻ�)���T�0 J���� ��~�3��	�����OI���A�OUN!q?{<��z��o{J��v��̡�9�3Fv���]�ҕ
��/[�B��\ �����S$
ι�
��,5���cI�`N�fz��ɿL\Xk�R��:�>��WPP���_��.Y�'�6ČT���e��̆���> �_�ͤ�e�\N4x�b��_�2���"̈�6(�#�����8٠+��H(Bd\�����P�W�5	�*zj���ʓ������ߒmx4�7�9.��<�c�������L�����QgVL����RY@�Z��4!�497�D��㕺�������p*{l� !�@�TO��l�ƫW����Kש]$��掚��MRjOo�fV�	P�9�r������� �sQo�(���5��le�0nTc*a�E�g�J�qE�0���W�Qf��wn�&��ma��މ�x6��.��\�\��kj���콞t.��6�7�z�L�bK�`��a���t�l�>�C�X�c�΋I��e�	�W�3	��o�G��D�	��3jH�5K����}�&�ߔ��_�tp8���{���9�i��׽.�U�ҥn���F�����{���'�o{����&�������_0�<�쮝 ��ty�ZL�t�D*ħ�s�}�����Lx�dJt�I�~(�Pva_��*f�) ��J�V�r@5���
��\խs�ю$EY�����XL��8��	wxT_Cx%*���;ߋD���5)�j9��@��aJ&�H�b]�"�'���d�\����
��G���%C�bi&�e�߭�i3*,��D��%��u�"��|T��[����W���?�<1٬�v�r����������>8���0CDx�0��_�y���{:����-i\��:��I'ɇ��Y��%��Y4)��ʉ�J�K+)�V����ޫ ���ڲ�`67A�NsF�\8��]�8W^*���L+�Hnu�Sg��/Pe9�4��(N'��'�Yݬ���z���n�/�M�W��\m��<���%��!�̒�m�rm���I�ͼ���b�8��uT����|9Ƿ3z}�K�f�q�8�����x$E����e)�4����Ss���`��J4Y��xܛ��S�A�F&؝Q+&C�]~بR�t���Oq'\�՘���?iځ�se�IǛ�������&�&�MSTv�I�44�F�k���~�w�h2ܼ�S�*��n�6��[�f�^'ѣD�#��\�!��O�X}%\:�[��q�� W7t��
��d��a�%Ε���؝=�F�ݓ����:2a�P;�9ԤvW�
�q(�Euz�{n�d���oOe�ϛ��-P���_���}!緶H^�bqӓ�X�1�F4qcT���H=�)�;x"+H"#�瀏������;��r�H�!��d�%v���z�u�s�wxLwC��3��F[��@���8-�r�G�h#3IY�q��Y�F����<]�H8k�ϟіXX^,��3��D̓Ls�2޿{I��Q�/��>�k�ҟ��� ��	����DW�
�y�q��x3��eW,����/H23���+�r/�`Ϗ�aXү��'����t��S?y��&@���ŧd�P�n ��}�h{W�h��ЮG��>}�q|���{2�s�x�JրR��^��Bn�ԋ������Ѓ.�Ê�ND�A&љhT|p jgu�Kg�m����5�h�ĸ�H��J���5HsPc�"Ii�$�V���T6�8��R�����L�98�∁�TW
:��vGGf<r�[3os��Rx�Dw]�0���m�w�u��������C&2�������1�������9�'����Kre�Tg�2X�V'V��o 3�+����<zzuH�~�?X0���&����C� ':�zx�wgX�B��S{��M��KЌ�E�Wq~o��$v.[����XI��}��
�g�Z����Ok?���Z�Cf9:y��O��)�p��� [��ҧ���<!K.=uM&�~�-�_��������6g�h�綳�YP�����=���u����6���ń��Q�5D$���zY�w�����f�d�Bj@�Թ��.:��[J�2�|��=u��]�L���վI�lؐ��.�tZ[�;��[z��m ���ˠ5N�7��������F�D�F�5\��	yo��7��AwGXf�ฎ�S��]��$2u�!��:F4:�c�$��$��	�YtMO�Ù�=_��g̺���v���+l�e��6��@	Hb���[�;�φ��q��ҏ�$*d�g��k��_[��AvG��L'��$���z�rI�l���3�� �]��$Bh���D�O"�g�
ܙR��i�-�"�܍�NGasE*�����ʄ/5�����
�0��B�5� �)�K�����`C���9U�*�pmʛ����8�}�2J�V�c
��Н.��������b��冩z��ŃEJdfZ��1b���N$��Z������E��hW��F6<|��A�5xy��C*���S�%����F��m����kܘö���xjr���=��	��)b�E�-WAa3y�-;kd����%�'?��vuo�׼M��ٌ��[��,&�Z0U���}���)f�H,W��s�'��f+�Qi
t+������L;�B�C���ȯ���	RE�&�ywZ^g���˄a;�|��F�!\ ;������X���A��C�ҀD\�;摣���1� _ �P>���܄͹ sCI֊� ���X�Ӗ%�4��Oq�SC�љ�gd}���Ź[�-�����):��H��*9�v��!�B�gT����O��㟏���^����2�y���n��КLsf�rJ�m	<{�V���'8�a�Ylmx�c�`��(����x�u��4�p��+5��!�I��-����������sY�/�Wv9���rCK��X���������O'�\E�]W�����>
3�b����Rt���x�:	_.�{cw k	Y?�\�ބ���G�k�q_rP��}�G���WM�\93��40�����K&t6��P���(����q�1���$�z���8$R�4��H��I�eo
4(�F�����#Í�����Uh~��|�T@~�2�i|?�c@=���d�C���+��~��q�()��B$�w���'��c0�v��U�Y:�ʲMG�
U�_�C�L��nQ���w\�֗i�[ ��"L�~�Bs�EFy�J�g �-�$�����>��t��/i��VK��}���t�x,�����<��a�d	������E���_꘸%*3��C�Q�^�L�ܼ��8�S����-.�O������}h{��6}�;^�s [$)W.ƪ�,�S6�nP���Nkk�Y_U����B�vQ��-��/�|l��Nd�dU�=Re��Q��b�#M��cP�]�k�+۵��?���+�Uw�g�S!����,�	��t/�yw��[=(�ͷ�E���Jx�%��Ud%�7Kjrpո�»F���j�i*��e�Y��B�<rD�(�D5:�:�Q�6�}ml,�_"�d]W�U��QL� Gv����"M�Sx\��6��l|�B�*��:���Tn]9q�R*U�YW����	��7"B3�02 }uL�l�!�'ܢ�s��[���{W̊�m� �A�Z���Av'j'Y���+5�hø��T�}�[F^NY��z"�� 4�C��t�bn��c6}�a&̽~��q?
�gߢ�2��k����{B٦���T�;�p��^�����"�R&�¸���	X�.T��`&��
]�l���Fs�rn�#��&�e��=������Ba�،��0�y ��G��_�)������DPq$��+{��pv�j�钪	H;k��h��B��mT�y-��A�,�!���+�sSN��$-Q_]z_]����ք�<��f��F��l�7wg��@G��<%�W!tʆ/K��3���Y^��jUn%��#F� 賚f�6���=ֱ����xES���\vJBϑ'��uƍ�b���')U2%Fx���X�^��N���W�9���E?�v�kA�`p��j��s0����SR��Z�
�NvR���D�z�XcZ�r���;���4�[�[�8!׵����:��a3�QH��K��y�������8�d����L�u��u7l�$k��-�����*6��t��no��z�`�0���clA�??)#�?��>nl�>�\D.��[P>%d���̋����*�&����<;��&/��F�����ɚ�3k�6{�2\+uX��r�#%=�~b�O�4@S�mx�GŅ�`V��:�Ku]�:����ϭ��%�mO+;��-�B2V���+>��� �$�����Q��$����i�b�^^�\v-gGp*��:!�����:�p1
�JNw)����b��v��ߕ�18�[XȫG�
�Xd,ʣ.:QxW�KNIz�0�*�!H����6ZVȯ߹�����Ϡ0��LA}�������-Ҡn�H�qǶu��}�R�,�g�m�C!S�vG6n=�r����G{�=����+�Z�J��0{���W�]0ؚ7P���'���J�ነW�L ������y�sGϐ`x�s��2f��`c�L�CF��7`�	���X�\�toh�%t1��C�/�*�w���ʡ,U���Jj�B�Y&�J2t0�獛&��З<�P�F>)!�d��W�Z�ރ��+R����bK3�r�`
s��HL1�2?�e#�hwK�ꎤS�Ad�M���fu���𪯜���tiO2?P2
�1��xU�A�f��֠��B+��Y���.����w�z�[��\qR��>])���]@X	�e��Caa^�J���bcʘ
��5�Id\��	�6{BE����0��e��H{���� ��&Z�_)~XK8��,ǟ���m�]��]�]^8���c���A��j6r��)R{ \��E���:k��1�����e��:��L��!*뻪�oH
M��B�R��;�u�O=VDK{���Z�������\g?|j!�Wvp��cv]L�&G�=�JR���E��#? �8+,`�5f v��\�gfg"��IA������UCL���z�}`Ʉc�@�2M��	�p�9T3�C:P�RGnX�������ɷT`����pd(�#���
���]?Ϯ������cWw�'�k7U�V���Q@O�z���.g��>jǡ�3�����L{ (�K��}xȝ�oO�J
B�����81��˷x��(���S�)�7�������)���6F�٘F	񜚜�>���:'ˑ2hE�vKMlڽsiָd��`��鿍^���|1��X�5I�ʮ1[�(dC��m=v�*���7ע}8���W)������<��W]Z/,��5U��k{ڀ�d@Q�{z`{Fy͗P���!(�`7�bЌ���"o�ź�X��BgmGb��jݿ�S�$M&�*�yK��s%�n� $	A�X/,���Xp�S%&�%�LiOF�sumr-u*�Zm���M��xz�y�2�NA���q+Ta'�U�Z~��ͬ��<�;Ȍ�87�6Ϣ��o��Jm��ӭ�"����_]^e���S�F�a{���+_kA�DE�u��,,�:"R�S�K�Ǖ"�r;�}U٪;�Q)�@��/cOy]6#�K��Ż)����ם���jquCa��H���ǧ$d�}w�z�R��^2���t<V6�����wz	�����m�i���a����7�2x0%�Y�`�K��v� �ď�HWXL�ۓ�z�O�}�w �F��LW��Ui�+S��餉��ƶ�����e~V2��)�G$���m�i�VKH|��p�OF��`��`�3�r�##�N��X��y�'1n�N��S��9��
/��$�:���""q������P-d����8ת�|�-t2=����mb��)'����S���Z�ɗZ�����0ؐ�OP��w9�4a=�r�s�B�ӝy)n�.�b�r>%70��(���ʄà�z�(�v&H�Ma!Cj�:�NS&5C53˛"�6$���������U�Rդ��7���&��!G�;b�3�)T�������od	�c����N���-�f^��4�1�c�$��H���>��XHHl՗2�Ş�ws:o!?�i���i���q*�niJ;�n	��gZc���֙߆N`����@�A8u�P�Mmf$�g�q����5�˅�'b����J��b|F�}�R&_iҏH���-�����ិ>�O��%b��w��4�׺���P;<<�|�U���
���.H9`�x~�e0Fx�h%�`D����9�IC>{�q���;��I>*�g�����S�F>cG�.\�Z�j����&��t5�2�XEX�y,���"A�Z`����:CFI�6�Y�Mn`��R���G[�`)��m���Vw�8�5A��6�؁k�7��^ل&��OՍ��Hz�P��l�q��ָ�~5��F�h.�xz�*�0�2?5m ���o�o�Y��E�hq@"�ۛ�;t';z��K��P�ȷ{��<Vؖ�,���`��� ��S���)I�2?�t�M���9���Z����k��|�9�ԤU�
�r�JT��N��mA��!�CP9~Fz�x��.���)} �F�	2&��'�X�,��!�	`�bB0p`q����H=4�F�	~�.H��C�΋o���r�J�?@�L��e�dĹv^_V��q��\{���?H�Xp`eFdq�ʇ��,ُ�5��K�ң���h�#���q�N(�l$�j<{�����P�g�m�c�x{z�{����/* �\L3��җ��:�ꮺ�: 6�H$�-!
���2Q��%���py�N;�t*�d��2_���/��C�rrxMR�4��A��V-��%�&�My�w;�~R��N�� ��\�R�6�poJ�h�9glߠ��H��Y?����~px�&����PC�$Gߡ7BR*�_���g��k�%�v�����G2��~}G��Ó]��>#&���@��U��?,,����ę���|�"��9K�<�9;#<+�^�)ʖ:�����ّ<�|.X�����~��t2�r�y��
�M�0�s�ݿ�R��uQ����lڃD�.}T��~��'j�PZ�4b����>��5R�M6���k.&�wyHYm^(@I�J��V�o�;��ѳ�sP���6W��5ml�d�# ȱ�\��#b&d��F�N*s�-�EU�n�����R�� ��?۫�Y�R��2�p����\�c���:���NP��7"s��4c!�e�BD�����Մ���uhg�_����3.����C��z��sv�$�}�l�Mi:iV*��FM���ݢ	6�p}O<����Z�ֺ�f\Dq��T����ZX�Ք�v���7��JuK��?XPg���`�r!�m�+�
I;�Ge��"`�K܈�
�*�WJ�a{����꙼�KEF RP��Hc�mT��¼������)���Ic����AȺ��߅4%���Sb����\KA}�Oy������yw�<�i<ͱc�����w���}>஘����kk7�i&�C�AW�m��E+�ȥ�?Gڬ���X옥.�x�5,h����a�ߎ���ݧ��l��B-W	��a�Ǚ�΄b	�<�{��4�v���2�j�p���֍6�>�
U:� ��;�<K8���t�����>�/�������7I���KsP0'�д��?��T�{?�~�m�2����^J�z��H�!��vvo�5vǠW5�tH�dk����7:q}���A,�,�~#�-�� ���ߜ�-=��bj����}�ȺNe�*N@݃���ҡF���Ş8�p��C6�nٗ� [T�I;d����*W,�X�{:�I����Mx2?@wQ�Z�7�B�04�H��Ftuᢌ��&��΀R��l���n��Zs޽Z�n��F�	3aކH��s�oI���Y�[er�B����c�~����D@���^�4AЃ��?��`���u��D4;f�>��?�}�����گ��zQ�W��O��:�ߜ��Z�~s����@�%�^T�sF{�[����h���0x:b6Ldp�+��7TYV7�ޏw.ԗ��B��N�:E��İ��wab}�VTN����@���Qy
�)��+�6Iy����~x\��e;�k����nU�8� q2�E򫁯��1�+b�d"ϙ�U@OD�a��;�	C�?����PYK��}r��u.Ul�����KA��/R�ow�=�*���|�1�M��Y&q7)(!���<x9�at����2�� Iq�_�7� 
��7�u"��km)V�C��
��^eQY{���f;�)=p��3)��敺};hj!mV�ϩS	����v^iu����4��T�ִ��Σ��l2���W�y�NnV~cBy���T5[Z3<E��'}U���NҀ�z8���#�v��tJ�õB*������-I���{t�x�vF#o���5w[�5��HU!L�Vz��w"C��`��C�p��o���-j�����:����/6AS�+�₾}�H�'-!�B�\��L(H2�(�a��&��T_���r����d�/�3�>!~s,��.8��d���oz�f]����f4� �����$0�]w���4����� Wy�=����V%��$JG�2kv����&�E�C��F��=�&�T�U"m��y+�K�D�f;CK��MY7l/a�UU�-}�
�/�	q�Zڔ��Ku�hB�Qc-�W�*�\��iB�伉�5sl������j�SɧRvF
(��VMbW��y�mM!�+�	Р���'��,�|�_�͓�u3⊡2��yJ�?zpDH�0'_TY �#��m,�|h���ҁ���b�k�I���Ǧzw�p�y�=�Fh�����*Fq�S�V!d���OÏ1'f؃���aw���3��JN�սҋP���!�O{d8H�))�}�yl�Ɍ�jD��]&/t����U/���-4x�z'�Oy`���m��a�׃�԰�yy-�a;�S"~���S�AM�[�/��Ɨ)����n��y�����񺷾*�Qv�6�H�\l���L�w��oD�U�����pPm�BJ0^�q~�戁o�o�7�ГoM����k�κ��LF�� m�˰d@*|�[)�B򼈻[�)�����7����BY������K�4���3R���7��먙!�)$�iU������Ǭ虘��'C�Ǚ{�����q�`|ƅ��B.�!��z�����1�2���5��ޗ�mY�x��S��āR%���uсCAJ=��~��CeSoCL$N�yD�z/d�ћNɜ���)�3ɕ*,f��j���Lys�ոd���Pc[? ��i�){���3�Pϝ��t\-j�r��<��5ȕn�p7��b�L��U�����bJ�~%�G����d�oǚ�{]��{t.RS���=��a��H��q�x�6��[@�p�_5���5gN~Vs1��)bV~P;�6��I"a?I�C� 8r�\�6ǸI�M��H��')q8�(�U��L�$���7�/ڃj�*l1��������ǳ��5 �J#�&��߷Z��U�}��V^��x��A`'���Ǻ���җ��(�g���;K��NO<�?<�j�1)&��_,PA��^��+u��'6�g�r��{�iͅ�+ȒA��F땗�z�a��9;wz�B�g�wF��F�	�(t�N��>��`j�Y%��I�G�G�Yq;�>���~��)��N�!��Sң�|A�]�|-
g��l8�4�� N�fǀ2�4�,��uJ���ջI+ �%����p�������Ľ�xN�(�X.JV�YV��:c�Dz}�frE%ĕ��g��ڷ�0 t��;w���.;����9�|��`��s�x��=�ד�A���n��
B��G��b����g�O*n���\I ���ZN�CA�WL��R���e�fm�+����n|4�Z�^��E����D>�ѡP��]d�$�f�^^�>qf����b)n�<τ��$s��"�r��]��w�(H+ �G� r�-��6z�t��Dq�cRt��G����%AUǞ�px�?��l�m�%��ߦ��Ӄ��g�L�ZC˾��>xT�\1
��&����*��\�S��hK��]C���ir���*	/�1τ���Fn)��ԩW`�hP�=����{���c�hD��ٛ �҄�U�Ġ*��/e��SV[�/6O�h�+�� ���l�bՕ)��)"��-��0���p��K�:�>�q��/p�(-��/�=�02pB��I��-lgWLh6��X��S��%.��6w��5{�[Q���yP'�^`�&���M�y�u�k*�q���u�g'z�h&����5�Nb��x\����*�jA!3a{po�F�6%L��2�2�B.��-�n�8���[}�(%z>����ֲ���[l��8z�a���&`{o��jq�=��
A���G9PȎy0����T"+�����&?���FP.,��Ο���}k`Y�| !K�A3�a����Z���z�~���P���.���e��_\̖��'������E�Ƽ%㼪A�Z����~�-�����SV�|������۴��1td�ۘ��0�5 �+�uc^���p�gk�s.<��3_�E�{ T|�u��,0&o^�mX���@���a���8x���"�Utx�c�n�=hy�����P�5X�$�l�XtL$�F��ޒ��_ghA�sB0���&J�`��7��ZC[e	���Q����}d��^ `���H�)Lm�	������[:��"O�1���p�/���#(¨�f�pر��?������{�x9Hъ�Ṇxū1w��L���u����G�1�X��+����>�bB4��+r�&0�r5�U�[Z/���5'�+�����U�K�(v�<�H�=���1ŏ<�+8#�0�r�X7�(M�>�B��݁��B��G;H�e*ܻO��������7�`{���!戋�e��0�غ�q��0]�) �Q��G��F�.�9�*�X��0 g�/
O������k�.4sCA�QȟE$Ť�HĿM��O�V�\$�������=���B���Suh�0�U�4C�1TA �ss[U�m�h:f	�A��ـ|݅LX�,��9���[@P�Yt�,�٥)��+Y��?�����?�w�z������XT�Bmh ���z|A[7.:�|T{l/��8��QJU��ZAD�����wA�%@��tL}O�������k?�2�4A��S:j7�b���(��>&�&�݁DA�px�J�t:�~Ƚ�07\*|8�HW� `l5��V����0�%�E- ��(-���8A�~�P C�ː�o����k�5�>J���n���.ύG��\�	8ZC�����]#Jɵ�JU'z
KJE��W5ח���HKfX{�ܢ~��.�`��8a���u�)�K��|� ��2����_����3��aſF�پ8������<ˆR�5���q-N�5�u�MB��vr�p�u��2B"����Q�p�����o�)�e��)9�����M$�)�|����JK!��>����;Q�e�y,���@��ʲ�HOs�x��s�u�p�S�F�vt��)Q8W�}���x�z͞q��P�<���'�:�
[N��2����Q���Ef�>{��n�=�H�!�t0j��j^�����9�52W��ٛ���'��4�_UT#�{�&,J���of�brф�4@0�����H��"�nr�&���L㾭�PN�!F�Gۂ����;�p��Q�����)�<�[� #�E�l�$y��������qG?��cP D>!y��ZR �2y���yv��
��>Q�q�?�E�.�]��6GF��Kً(D�[Ves	�N�����-ת��"�����j����y�X������W�����Lowl}=+QH\�3E���AXM�� ��{�ˌQ5Z@����p��I�W��&�')ᛲ,{�]����f���[��U���9�䉷�rܜ=Za����[���]>a<���s'�@��'��K�ݠ���1�L��������;���\{0���0C��]b�W$��g�boq:�/���ݖ6TLd)�)�	c�L�ũ����\}ѻ����<P��z���Ш2�, ���-d3�K̾��&�3�4���o �7����V�7J�է��s���F��%�.�0�$�zɳ���R��_i���ݸ?�%f��8~�4l����?
^���4EnD�Ζ��gZ&�)oEnD�osg���/�b�'�i$���cIdc5r�զ}�h�;a<�g���ie�����E���w��N��d���!��@F�Bs�-�?l�iH�hst��Qh�#?p��Q ?��d�ZSx� �nv�r �r���d�$���s�}N��
.�W��Fl�YI<�w`RTi�Zq�єN.$O77|�P��i!���u ;�,_�X
�����Ǜ���"�=��i�.ZU}Oɴ5���  v�F����!$����>������_";'�P6A�*�eg�h��NW"C�<e�n��ct�V�.\57�����(\�ӣ�XVqv�!in���U�ʎw����K���20��rV����#�Y��Â~�Q;�{�?��S���`�j����|�]��K0i������ǃ~�K���=ç'�r8�:��\�O@��) �>��T�L�{s��_ϲJW���'��.wa���|��ċ���LTɗ�"��Ĕ�E�?�M-�V������hơ��|�*�o/k9D0_c�>!��)�Sv�C���4{b��Ckd"��7�V���(˧���	1�a�Қ�L����u�Y.Z	����r�b�$8���A�{A5�HLȂ��8�r�b��HO��L���zN�*N�]��{�,W���r�4�̶������S�^���!�e܀UZ�Т�S���n�:���"\�0в�J�X�#�LG�^4����Rã�vd��0��n���
<",��H	8&����u�q���;@SGnu�_$S�։�����J�$��^���rʠ��C4�׼X�yn�SJ�'bw���nW�}�R�s��}Uu[`�-��@���&�PЇ�/>䍍%AN�~�*N�����,�x����r�T�&4�/U�ً؊1�c��Q��.���U�h;��1Z�bK�υ�1�l>��%�
7Q/�ƺ���#��m��:�Puhk3����ყ+ͮa;�(I�kJ/u�3(�4�;��F#��re���܅�,���+o�2;l��?Aj����ΣՊ��<�-�-Q���xT?P3������Ǔ� ��2a):����m�-���m�t��q�$�h�$	GF]s�b�,�\n�kBs��\��~TI��ȓ/:	4����j�P��ƪ�z�$%An�`-�qW�h��j���N�KFY��M �˭qA!�tދD�BŮ��"�h�ٹO����[��@�e�3YѨ�y&m�x�MG�&;*��;��b!���>,�'C%��1w��U��Ջ�v�3�(�5(�x{h�ì��5QWm�(X���8ߩ�+���kn᤯�Y�k,����L�;��֥jn�� ��j���i��)r[g���5��q���$�G&_�V��^��o+S�B�M�,�X�GZ�P�+����vO��d����K߹_^=
��s=��i���H��&9�D�܌��*���<^�g�Я�.n�DMzU��x��KbG�}�\9�ξ�> �'Cj��C�|���:�st��"N�m	�H9ꕭ�[�m�����Mm��*��Q��#�@��Z6q�Z�`�G��}�!z���N�v�N ���tF��x(u0gv����S�:�و�$?��+߰�2'+�no��(�D�s?��۫���J:X�?�L��j�sP��"���B��ZA�59V.��X��J��&��ۦE4{�7R��	TtaN�Ԃ��Og����;�##�������	��n�3�C�x���UY�u�?֢������Q/A�Lv��C�Vyݫo|V�hW� ���)�|ք���cڗ���-N�6�Z�Yfc�ΰ$����MƮ��t@#ѭ���~��&)�5�[�l��3_i�q���[��a����� u�Yo0�_4�0�fN��e�q�l�~�[0�[�Ї$��l�[�qH҉&� σ���������3G+'d��=k�s!E��,Mu��Ǐ5��|��P�����6 �[5�i�d3��May�_��2����`]���L~����l���ָ�e��C{������ڗ��?*���yP[�L���b�r�%bU~�>4i�ؒ�0�����YA��x-�<�Sr�;��u�;�=��;� �2;����,���虚�W�W;��9�,�\4Ƭ����u�BC�	E�'(b��L.6s�	J} ���w�ZBB��Lm�����J(�G�Zn�	����־��p�j%�@jh�U�e�z=�x����K+[e@�b���byN!��ǲ���C���͔�
pÜ i;P�K�ܱ1� ���9��I��O��=�G
�\��*w<37����x%�	��e�e�py*�T��;���O���J�p�����u���G��|�~�z�,c���
�ڵ��ٔ�������Y�����8C��Ԑ�����OGГ��9����9�}�:���0��c#���w�ѝ������;�U���;��"Y�e.��2I�ITi"�R���|�`}�4��k?��o[�N�4��4?m�NPظn�wt9�F�n�N�z�����|�'�bo/S\�E�]k�T��QL�XW�q)��<��D��P���%zJ6���۝s'%T�	Vlmt�5φ;=h�ur�����e���t��:�.t�`*�ߩ�*x�Ҽ�GMl��B͑8���b�C�5g�����_���6��
I~0���!�?�����՚�C��y8os�Љ��O��M�����c��A�l�յ����?���tֳΆ����pi@g�[{�d�� �B�{�%Ώ)��6�݊~K���`;��ڜX@�%*���@nrطmҫ����e�!���s]��}�QT�M_�h{źn�=*��ra�r�Mɵ5:�tt4g�-�5�u����eN��S=����.!��SbkM�*^�1=z�q�Z@l��JV5{�@6��أ�a�s��P���9k�P�f��F	���I3�'��A�0�t�~CM6����EL�P)���@�\�F����ҭmyV����i��oԛ�a��ނ���ϖ"c'����4���]���T ��&�+�-@]��:�DQ��y�	�y �R8���%BU�vk�����,��=��E:>�QO����Kq��I:��=r>�niR�Q�����Z8\���q���4�c+��T}i�PNa���B5��d��oti�d'���(���1����{��/�c�!)6�O�*$Nō�A�,+��ݵ;/w�y"��U�Ȣ�Dk���'�l�ֵ����Jƾ�<k�D�.�$�+U��J�}'l���y�a���3���!8�G�!�0]tO�ȴ4�������l�$�
��kcq��w�W)e	6; ���u�N�s�p�"���4W�R�5���u�`NQ ��
��<�ϯQ(���!f�'�T ��H@1>?�$ma�J�&b��"�$�Q���^ja�'rRW&2����m>c|M%tN�E�������|���Ӣ䛦�-�ӧ�8������čQ��dm����W�L�=�z�������B�C �}�M#������r@����E��z�F�N���"w�+ُ[#i�]�cq��f}�]jՓ��#��~=ˮ�e���2'���to�ka��������;�Gg`R=s�%�v�Nk��2�a/��X%�5��6��c�ؗ?W�Jz4���t�\bߒ!��%�G�=E��
�Hy�G��`��/���6,������ùx�23g����1u�t��b<���b'�6��0;ٚ^��*J����8���m�c��])�b�H>�'}
0�ћ�X�mh������mF��W���V�e'�^R��ż���@���I[y ���KS\z'.dN���@��J����i�t�럋h�ÿ9�N;�?���f�����]��������e:Y��4.#����R�e`�\h����x�㬊�ґ�3fR@�d�`��	�ř,(/�{:��{ʠz���\B��9���\���姼