��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
�u�,k���L��z.vJ~ 5&�a�+�%�����n��=c�DS��D�K�;��.��]�W)5��4jQ�l��u���ݕ)$���r<��p��f�0���G[�
�!������2�n�c��Bl#�L���(��T��
��$�˳2�������O�Q���$�j���5���4�\l`<$S%as��^��n��=�;4��M�w��	ٝ��İ��T8��y���,��k�ne}�)s4=��x4ő�t,�?�~51c5��`�2��hG���ߏ���0SVo��@�+Ht���g��xV�/�f�51��6��fk
������d͉7�q1&�|y��p�Kʟw]J���{��u�ȓ]O�=���\��!���;L�po5�G�4f(�|�	y
;�lQ�kU��3�3FmTo�pܪ6n��<݅��L���h�滊�3�F �?{��o���7��9�A��fr�_�h(�-h�إ�}Fj��K�)��P#@*LM�:�L'�u@4i�':�I�7,�{3�����\�JkX�5��#p�nvEz5�TD�
[~q�qZ/0	�b)�3��vV�s�`eȢ)��-A6EN���c�; ����/'d˳6��mŦ�K�A��Eʔ�=@�������G'�O��7�\����F\�V�Į��vX��3��[%����j�����x������{�y����P�F������`}�ݗeC����2��s�%b x��^��͔�2?5�C��I���dRtg�+`�?��,_�\6g�]SH�2�׭µ�����ߦ�ǵ�P��u��m�\�n��	�Ũ��}�1�ȗ��B���	GT������x=��
�̃e��N��;�G'�N66��<�&��z
�r�h0�}����_�<�t�}y�ƚ$ڸ�1�L����7W�Wg	���]�ȟ���p�ѽ����:XS-���e"tG�`�~��J��ł�e5Ձ	Z��e�l��@7ӏ9�wQ�� ������õC��A�4�_���U�%�I@/0�恢2#aS�+�[)��|���~$S���uJ_K|I3� ���x���]$���iO�y�9 u>K����]��U��9�p�qȌh]��<So^�Fe�?��`��SOHӲEK�t�6a��ƲJUj!�}MO�ۅ����n8{�{�����Ɯol�8"ټ8���h6�R�ظ�W�v>�vV5�!y��$�|ψ=͡���G�TL\�9�2:
;{eh�³�o��4����|��9#��/�cO������*y�H�@�!�It��ܘh[0�X}�x��k1�֘5��$}�F���嚲�E�3�u^_�
�[,���r ���z�|�J��j)�!X �Kfs�ފ��m=�����$�~G3}R�r�1ۆ�����V�FG��4/?L�y��K�b���F"7���V&�1�M�a�A��q��ÎO��U��ぽlt�$2OӉ����è���3L�y��No.R�p"�Ф�J���X��J��V�.��J��%�Sţ;S`�<9�{�!Bp|���1��XjN$_6�S�R�BN�O3�
X-�T�C4L�n����5�C���^����'b^�la[4��xUayx�_����0t�� g�tax�4�q�lg"�#H���2�dْ�Np(��O�aj�����݈���=�):��r�Vդ�b5�ce�D9�>�*��'�['c��#d�PgF��Xb8N;:t�?S���tg���k�F�T�j6�,���hT6ƫ�b&np|�-$���:)��xD�l6Bo ~�a�"��ݍ����vD��P�z�v�i���nY`(ot�W���-��z0�i3��I]��6YBJ���C��/�J���y�g����w{��ur�z, rE���T]� =�ڳ�&��u`M��L���َ��0>�/x��3t}���Ǌ:5�&Ҁ������%T.�練�5�Ҭ�;u0Np�E�+v�g���|u�]���Qm�����Ă�����PT	��յ8+`a5�c�\7���"�J�*��ց;�S؀����1	u�;�B=a�ܓ�9�I�Iq�ZW#3@dD�S��
�HR��ZI7�5xa��B­� ��h�g�����'4\��	��F?R��xcf�Z����n'a���Iq	LN���c×�t�kbE2 o^ٕ�dU�âUH��0f,c=>�$���~ܲ�x4�(��1���Ttm���pGhbs�����X8�e���Zn$��*d1˪�qY{�%Q�:F���C�1��U��Rc��9y�^'n|:�.�
�&�ca�`9���B�>(g��m���`6�Zn��^��<`1�#7b�d%|�����(_��C����3�6��w{�9��h8ɮH�ܣǮ�~�����-��@�w��Ew��5�w4446��3�����U/@Q��\lq񧸴VͣD�����[C]C���1%�Oǫ��Z�o�e����7}t�����SЯH#�Y��� �K��r�ۤ�j"��E���gj"�� ֕��<�����S/_KqU�<��p�3��?�p�\Hz�m�ܟR�Bn���9�r�s��m��x�2\��Wr��*�N}Z�T�f���&,�r!��A
�k�A�u��EW�k�I�������Κj�G��Er����}���/��g�p�����	�C�"U�5eç+��P'�<�����UAlE2����Do=MU����j���Z&���W��?�C�.��EB��k,R�
��� ���#;��{�g��8���T�a.��j�y%ͤOGMT+v�zp`�@��ˍ?�s9�$CE��P<ɸdvZ��0�R���E�P%L�i]�*�t��G��͓�1UH	�V=)���W�$��6.�H�G�-�k&�/?;����/�t�O"�!XHp̊C���sQ����6q�|�[O~m��|����o�˧\��L��� H4��{8�n'�+� l�
)[�=�������^2E�iz��h�c�U���?Σ b"�A��9X�WٓU���#`tK��N��������F�w��W�)4���0_�$��Ҩ�����'��ϖ	 p�6"���C¶���Y�� _d�mĲ���ڶ��0�k_D%8�1��%X�良��C� ��d�ev\cx�y�͖G�w��΢*~Qp�a'��s;�q�C�����%�����w�,��A@6��1��RG�������ǥ���dgex�l� F秙����-�7䡐�Y2��!�Z�P�UU|���M2��,Q��H���S���>}��6�}��T��6���r�u�s�4��LYg�	����g+k��-�ۢ
��GB��fԱ@�M�%�/�̀�׎V�<{۫k����Wx�1X' ���*\b��7���q)�$=�Vf�n�s�)MIyF:�TWd��.�j�=z�)���~�0�L<�r�e� ��Y���&�ur����+�y6y�H	�bTq#��"6pt�-��T���i��چd����r@�
��-��]F�I@�6,��l�0*���-��������Y�G�B���V��?��=�a�����k2���� ��tW� c�ZSan֑�ǅ��u�!���;\	%�7��!����԰�\l{E�d��
�\ı>�R�oEx�T�3�����A�m�fč60�����R�l����R�H���c����@W�V�5"�ms�x�kΆ�x��!��*\Һ���*~�c��p��w�0�u�E�]���K1Y	�pC�-1RO��W+Ā~�6^�U��m���L��Ԧq�$�!��-.ge�0
x�s]L{4�ztag�)�x/e8G�U{��h�p�\[<�1n�:=@b,*���j����J�U�og��_X|�J��ͣ[�O�,�m׏���N�ѕ�#��k�a��գ{��(���b~R�.��H�맄��.>TIc
��@L�!����eS���b�bzd�X��e/ո6�d��`��@DΤ���!	sGH�N���h
� �P�k��/�%��<�9A^*02<5h28��~�nԩR�C���0t��w�&A��g�Lf����� ��]�N�I�J�VP*I^�)�lp
֠q���&�O]��E.��9q��>������ b_���c]Ҍ[{�q�|8Y�"�w*G�7zj9�h��/�)����1��v�ix4�6 �]TV�����t�qT�!))ڔ{��*u�"��b�WCJ&)��	��u=tl[�ZJX�X�ml�O�l�d[e)��#��������J(� ��H ��R����&�hzu!�I���Ә�f˨�yY�0ڠ� .���옛0d���K��cN��:�����d+��(ir���B35V��G��j�o���-�tl��o�mqf�
u\�ð��N��,�$c�g�:Tj�-D���A��nF5	��R2k����jitǠ�F �i���qS�r� �w	<_c
�_�!���$�ݷAMZx�-�_~D�r���>�x*E�#a+���1����	BM���d�%�;�j<kX���*kP�oѩ�B���dC�õo ���?N`�]�.�I��3`�r2L2�j�bf�:��bQu/�G��c�\��̜�����kw����c�iE������Jp8;�
j4m�4x7�:�J�#��:�{�yR��3C!�\s�Ʒf���ZT��`)&��M�9/JD��kŜ�W�e��3�4_��vg���R��� ʷ;cs�iO�ul�f*V�tt�̣�Ud�6uRw�Zں����lϻ��
�6Yg/��t(��o����Y���9+A�VW����_�<�&�:�������(�w �Sg��8�x�ӹ-1^d?�~
 �za>�VJ歅�Ay�-��*ŌI�,���ꉠa�Rʔk?q*�9�nv���*��?��̕z{��Q��H���}��DI��6�oɱ�u���:�e$>���S]�q�p���k-U�-���bQo��;2!�v�^��g�E'ĦCLғ��y������#�l��EW���o��E6�'���#ۨ�IJ:�-BhS|q�"�0ɞ1!����S1}�k�Q��u>�h��Ԅ/鉲��/a�\��V\q7h��&�M��J�iW�fP�_$�X���\�N��u�	 �%4��
����ژW
�vy�� e5�`���q���M���6��1���)yˢY�53�"�B�UQ�$|tV�_)]}�tA)C�%
*��w^qVсP�n|���g�:)�v:���3/�޴�z߆͸����2gbN�j�>l	���a��.��%�`�g��j0��q#�V�G��f	r���p~������%��=>�˽�6��ץY�|a=hx�7I�ȊD!���ő�>���.^����u���p.ޣRj��z�`Y�C1ja�𑒃iY�hI)-��]��2R�Y����Z��D]dDWr���'��_+s�b��������;�f����0�6<�(¯Y5�+��%��0�B�N�n��!i��/TC�5�z��Hk����|,M?l}V����F������d2�]�E�q|q݂a�?z]�A�,��Jw�BP+XF�ke������1��U�����]���U����xm��=|r
c��M���͟���6o�\��F߲��Tl���g�T�qFםD��n�D���}qQ�ɸ��$o�i��twTZ��*_��u��MF�+�3�����x�����)��h$����������?�x�9uv8|�N;j~�N@w�#i �p����խh�r��H"J�9���k�I�Wk�K� j�Z4"�WTyCS�OqL��2^Z[\�-�0�@��'��!̳�W�:��g��;`�C�|�91g�m�v��N�[FpJ:�ѨR��RPF��(���� �����C�
�u��I�TN\E;�R (c�
��x�N�|,A�a

W��쀞ەj��Ѭ=Wj\ ��{.㙖�mۼ����[V}�/E�zwA7E��&��_�8n��U&�X�̳b���ܓ��6>G�U��{��}#�XGx�5���H;O�E+���)"�i4�O.��opc���?m������V�5����_pJB������C�h���L��o����{�S�O�l�գ���S}��H�@\��[�e/"�~�r�o�P����aI���6Wi�tjZ?���_l?+��$bW)��=�2֟����JD�P-�P+� �\bPn�	�&�nc%'b>A�Mze�#�?e��u���49%�+���8�=�*�}̕�~�n��ȓ�!6���m�FO�I����;��Ȕߤ�#o�������qt��ˬ�>x���3�l�#��Xbg˷��.�+��9�Ѯ���(2.���xDѿ�/K���?���Oh��9$���X������(Ťx>`_Wn`�@G>��8�~o	�ꀥ��{��G�C���u(������C�Cwl�<��W8��e18��'�b�<.��W8Ѩ�A��/���EG�#
�j0\.�{I�*��ӳ��d�V
^������蔴��D�is��~{]�����K�'ÏM���o��-L?d>`4T�eq�A�:
0A"���ő:}8�-�C*=o�iUIR�Š�=l����.[ ��y��>L��^��k����J�� �m����Fċ�j{�M�,0��S��ϰ[�����L_81�H2F!�V�uv��L�:���m�I{�d���W���-���Ə.�a�w�De�J�4�\�������PH#��O4��D��}u�=���<R^�k��bo��TuK��r1��y���>��qb���͢A��:�בyzo�D2e���`����H�KZmu,��K�l�H0�t޼\, N���9�J\���;�ڈ�'�y��^2�<����>6�57#89��MF�t��^H�Q9Lf.34�1bjm)�_�Q�X6�Ǩ[��D`DV�2����~��`0)�M<h���P�"$�#^�Ya�	��b�����f_'�<o�n�NN�G�G�<"�tZ�؊����Aj�]��'kc%��C���'�Iʇ��
��n����5u��D�L��L��{���1����*��$,�CK�Q&k;T�q6�KOz����0s��$�[T �]�=��D�HΘK-�t�{���m�^��k��u٥���n���ȧGL�U�\�1�����~��"��ѐ���A��%��ox�*v����0�[�,��Fg�{�ӧJ��d�f�@R^�5{Y����a<�ō��0V���"�YTo��������ȑ0 Ey�n^�e�o��l|pɅ*I�3�pŕ�j@j�Ƽ����>������Oߦ5�Pbҍ�ޫ�M����`J��^}�r�D(�(2���x��]&����{�*��*|�c&���/�E�Y�~k��
�nΦ_ �� -tI���|(;6+�z2�s��u��x9���vf� ��t�X�>������D��:\�F`F�^�8��h�`�a}�p��a��AK�Xx�s7
X��Bs"J�C߻�x��l�Zf<MM<������Xx�KT���>_�mL��~��-��Sk����oCz��+��qy��6q��)CLa�_��X�8���+�O���4�e�-�W�x�Z+}U>�~S�HD�[��)�5e���D�� x��[��Q��b���e���%R�7).�GD��<�:�9hȻJN�#���V4��yM:?�(x#�o��13��6�0�Kw%�1�N0�jӗ��ޛ��$tl�� ���\�lwf�C�wDV�[$�pE>%�k(.IodD�>͓���\�`�9��e4��Y?�ñ���~/O�Wf[��
�=%"�#|=�{��vE#A�����5u�Q׶hF�_�R2c+�ؤZ�)����s���`t6��K�nn헪XE�D�V�I�no�H~x����H���V��-�k�t����,AuL��ϙ�:J%�M	������c�8U�,L��c�^�`|���Cm�0<o,����<�vn�������CCZȉ��שMQ?A���t|�8�R=P �&�~֧��ՠ�쯥[��l݁�]&t��)6KC
ܔ14�bP�����ͳ��C�&�퀪���uz�j���$�ѝ5���߯7�4�#�TL��Wj�
�Y�A�z���0FaVy���������0��~|{$�1:\�6<��i�^���4�q�-;�q�B-���zl../���m�ꐯ�}���p�I$4�8q�����,>�g�3�N6��q�ɤ���3�fba���D.qv���x��CE"��nǋz[(D� c⌺t�0��j%��z����k`e���f�X��~�E�c��]@�Cd���m��.���;r�؏z��
��88#�h,f�;��V6!��Ϙl�q��t0$C^��& Y�$[��Gk�+ԉJ�W?w\5R����^��jq���c����>2H/j���/u� �-���}�c���6<~��fu��K�jP-��	ª�KT(w��et郭�Q�$�9ؕ�FB�2��6Ń�#j��k�H6'�\M�7�´E�5<ч&��a��e\܋����}�6�/�1��u5�sڗ��[#��-BIKAS�����hA�H�ٺ�����b����*ܰ�as�&�(,r��F�P<�)�&'%�O�h�K��\}:�vv�d����8�gWF6�D���B2�j�׈�?c�W@�5�.� �w�@��a�8G7���v�����ŷ�KF��B-r�R%)>�1r�0����1�l�ʛľ� '|x<�@�3с���l��|2G[�"\,}E%�w�軇Gb	b����*<�ʽ�[Cc���sP_��c|�ś�L���(ۓ��
�t�@�ώt���!QwJ��J�Hv�9K�k���.��Q�[���{<�c�Oj<����m�ș��B��Y؆bB��s|��ȾC���w��]z��})Ssj����M򵞶;
ܝ�nu��¡l���;��(q��p�m=cf)��-�\UiE嬄Jh�Z!䌲��Z�+������+i�6b[+��� i���;S��c�8�O�I���\�K�̟��h��1����.|kno_d���4;G/�0?�xy+"���r����!��M_4;�����8�Q�LS �k�*�����dMA8�z;����B��O�s�tuh�����s�����C�o��!òY&�«�t$�ݤX|����&~؋ʆq���q0�s�,^����#����ySW�ļ ������U�v.c��y8���փ-�j8�d�?�S�O�4�t��K�y�}�m�kv� ��������p"�Z�(gr��?�(7Ƥg,.�L}�`igTPV�n���Sen\B�������`V���a�Ⱥ��tfl�r^��Ѧ@)�`��Y9;4����E��,26UĄ��۾�Sbo�|�(;�=9s��ˈ�Kb��2�"��j��F6ʹ�m��L�������$癏���lH�#>UL�Vj��q�C�ic���~M����{9?��/��ـ�73y��q�,��M]��+��J6d]�S2�'��S���#y�}�T��$;��)Gd��/���$(ݑA��*q���<�[��~I��	�oglL�!�����_��|I�?�!3	h�N�L�6�PlZ?8�j<��,F�ނM5�Ti��8���aʞ��$��ԑ���s�`��{!�A�6�Q�ȇ��� `��d;�oFJ>�����㚯�3wzk�͏8gp�q�Q��R�7ԣ��]� 4$55�^'Y��C�����E�l:Y�ۈ��\T��6 �y]�ʒ��~()�d�?�����bt�?G�8�w��<Nb2[O�=-WX��@��?|/&����Q����`��QA"�(]��S�����i�M
�}˱+����Yd���:y�UF8�)\�G�ޔU�w �p�E(�T$7�]V:䛛k�X�����N���B����;fӬHp	Y�;;�t��~^�A<t�h��¨���U�����oQ{
]�
�xȺT�i7~��rj��Rг֠BW�`�ׇ����{>t���@=ZQ1��c3ޤyAš*�z�`�~���_�. �c�8�oh�N',�+��X��2��ٟ���b�Q��
-��֬��8���6�)LC~p�K�����t��j䀫��U@V%F��YK_~7� ��=}B��
��eq.&Ƀ�6���YC`A�V�g���k�m��ܹ~(�O.�VZ���5<�(*�3	->t�4�1g�Ju��w���^��S��fzfA�&B9�#,S`�ywc�'=�D�M�9M���=!���C8E�(�� h�g�=`���*��oY�����	<�S�ڱ5�X�K.��NOOdB%�&tv�'
�U�>�P����e�P����,:���2�$� ��t�N����"���~��"��i�\�Q�D�q�NVy�P�+ܳ����������Pd6�Sn@�Uo�aG�+ �Õ����>n�3��,��L|���	���~n�?ь("��ܲ�M��ēbX�|��<��i��mO/D�e��
�I�)�{����4�N���`�l���EJ輒� �M1'��A����72AA3�*P��Gs�ۂi]����;U����� :���GJA��$)�SE�eYғ|�u��{��d17�Gz�g����C�@�8��G�N���8y�Q��}�G刊	)Z������4��E{�C���q������
����_;�o����G�׍��"d��>��w!�x�T�L��m�s>n���w'rB��_s��)��[D�Խb3�eI:G6-��>m#�RJ�ȍo�U�}Bp�K+m� K��U���/$�����}�^(ǭޗڱ�"��ݦ����5��g�6��BN�* V0�Q���9��<�C�`������xH!:�לN)�hO���^Ds$�K0\��y`�-q��9���q�<g��H��Oa�?���PN|����`c�����_��[-��6��HYz�u�϶���(��Z��/G�����Ofo]�{�Ԃ��T�j�e���wT���X��;�&�J���qAǺ��`1��O�u�vj}�{*�7�ͧ�s�l��>�u_K���*�	����bV�M1M����㸘N��a
�?Zf,�/�Z;�?*��]�Ɠ��9��������j!���E����2%�;D~�J��y�82���9u�&g�ԋ@
)��'*^��������`_tD�h��Ʈ��a���9L��kSL�`���"��n���_������Hlp��eHOB����@��4G'-�'`0mP�]���(@��S���|�\��ͦ�$@+�k�g| �˹Vy�^WsS�I��!՗�$q=]��f�!�4(���oX�'���f�o2�W��x���႗��N�tD���۝�,�P����!Pe4����>�ܼ�^P���A0fY0\$�.2��9�>q.Ш��f"��sh������ @S耮c2U�RP��$�5��&�x+9���ϓ-�2#`ޥJ�q��爨ha�*�%��YS���j����I�Z- f�gJw�3X�~�b�^-Y�H�kJ��N���[��2w�D;��4;`���ϗ�O>�y��S<Oe���P�jջ�Ew����ut���+澈)�H�)E�Qk������JQ�r�< FA�c��~���X��P)&�>��J�=e?�uX���z /�i�u0-����n~���Ɏ����~N��k;��Ө�,�e�H�2;O\���ʍ027>����]��q���`lE���[mm D�~!�&Ǿ�8�^�\/�V��G��>cX�Fg�Lʨ�����k�ڷ�����z�h�K. I�dm��(̫p��<,t��J�2aD�8��>wS��z �|��X�xl<=�~�_2x��eZQ�d�T�c�?1��D�{Cd���>d�u��~���Cb
�2�%��v�
3M�0�h|�� ���[����s�?��?��:_�V�ɵ��̓&4���;|����Q�>��)�Co��_Z�'-�>�:����}>Y�>[	����^�e6�gm�2++y��;�� D�/�����_=�Kt�šPl`�4g X��y����6�-�U�s+ԉ�=�
�=lU(��Y��mK�
?	�����y��鄈��|�gto���C��z5��x��d�)�SGt�j�"XEXk�w�3rʚ��M�{ٶ�a�����H��YW$ Wz/�Q�U�&V+)��0��e_�ϜA�c�?�x����U�GZF|�	5�_~��m��AĶ�T��y$73�!0jM�1̘D&�s;��
I2i�܀ԁ5ܶB�uxϞ/`��X`_#���s���R�t�w�~!L{|e�zE5 ^�D]0!]|7>麅q�GK��y��6��P��y�oD�D͘i=����FW��n\�]*�3[��h�$[!�������/��w/���sbO�Q���O��#�ՍO�4K9V����єw43M���OpY���$��,�Zӣ~�y
�R>j�+��"��-b�4�����4t+�w~���a���9(��X e�?$9��Ӿ�ڃe���Ƶ9('��C������>J�N��_��T�vnW�		�:�z�uM8�Y^��D�>%(pɗ����r� 2q���=*��{���¤���Z�AÇ��+����t��j�yf��F���{���:�i����z��$��8Q3�g�ZQ#�7�@��??y��A�L����4�K\*7��賊!�
d��0���}FԄ hЄ�y�IU��%~�>M����X�*�@�R6?jz�7���I�(�	����c1��B��mF�آ�8�y��I6�i"(�W"�؄ٯ�)8.��a	80���$���H�i=�$D/�[+���qd�5����˯˖L;�r����]d�aj���#jHh���<�@���4G\9զm�����&��S��\��!�s>�G����	_ٶ����n���#F�$�#L~Vh�u�'����>_J�00��� ����G�_�ͬ�&Z���;�F^L��$N�?}�+�0���Am8	�S�/;���X̡��N;<�v8�*�RN�0@ꒂ����冀<^S5gk�����mS��|��Ucw��=L�����@�ݯ��L,�^_@1�lZ��5#�����\���z�b{�:��P|�S<Z�OY�u�e�őS��&�*�XS�"Np5�뱜��.��XF	u�ȅP�{��{0�If� t��g�\![��h�t�^g\gh:�*J���i03aD�T�ʩW�6&[Y�Sԋ���D1\m3g����VN�=��铐������]��;�j�0���d$e\�T_a鷮�g��B��׍J�O7!{�QyWܽ��6�m&GTa�4/�@P�c�/j4Q*�����՚�b3ƻWr�^�0��VǮB�h}Y�A�=1ΐk�����|
���OG�m
F�� �&b��9��
�k�e�Cy����d��%��ۑ(ے�@a�tx���_ӓ���TU����H��z���U�4k6��3���*����&B�O�*�R�K�Yn�w�zx��u��~�>�n]{��m�k�t�_�ɚ��P��s�S�Nx�I'���)'��?ٮ��z��$a+�?����V��Ǵ(�F���*S����aʄ��V\GE�"��7A��J�P'�k�	��j����;�z�[.O�`�΁{Io��"��*�fT>+���Qkg�a�6I>Т%X�t��܌��w��pM��dv!L'3yA�v�6�ǂ-�7�,�?檬�헐���|ƅ��8��R����o�P�2e�K�u�戋Ґo�pS���@ 1��i��`����/��7.��V^���^-nRmW�Gm��R�<�y]X{V�K��q)��
�h1�N�N��b�6�ft؅ԭ5���0�����%=)6z��z����u٣�r)G��#ɔ�H��␆��z�������+����d\�Q%M=e;KB���V�!�^DO�Z�e��jZ#|�%�������ʘ�ӓe@V��� s��="{l�M��Y��S�J�X���%�\����$x 2�m�$��=m?��dҨ�m��i�Ic��4�\xEk�<C3΂�����Z�t۾x���`����tѵʹyusנ(:�?�3���v4Us+�_:K��K'+(�㙞�&�d@�<��|���]h��󩘴�{�~3N�'��o"��36�|�ѐ���H-S�4f��V�l�7��(�>����e�4����|�ߦ`�#"wRr��<����q(�U���c�XH�pe�gy�Q�˨q?���o��7���]�d'PYD�D
��B_)Ŕ��Z��6�3dv��l�ߐ�G+WFV�JQf�p�cZ=Z-ڙm㗿�������0�8~�#eRY�,ME��r;v�s��v��E��W�mg�a1���v��e.X|*:�ʯ+�V���|_��0��E��`>g{®��W�1;��rJI/$Jh�
 �����]������֬�/�U��Ɏ×�a��WA(�^'�4�Y�����Kd��:���
����Z�
�"�ǡK	ܨX�`�"t��Cx ^���Q�
��!����׎��wX�/v�Ƌ �'�Q��@5�
�^k�*�j{�儕r��+��CjV�6��T�J�:z[zH�B��˅D+�/�l����]f��g:��F�+�B_/�'����bO��-�p�Q�:�S[1�	D�'��ф��<�ᩙ��B0��H߹�X(ED��ɟi|Ʊ6���;l2Uz�m��F>Rn�h�t�n�ɼ��o?��Gp��c��x��h�ǡ#\
��O��h��l�x���Y�6�����g�FsL�c�����_NP�f?�2/����O^3�K�BGT�~-��=��r�6?��u�S�v��O�ˀc�x���Z� �ʔ´�Y
�ꊅ�$��H�qC:D��d�R���	� ��m0�hO�d@��ZГ~i�Ƙ�J��$�>�e����H���Z%��A�/4�Ի�Rd��nնD�Q������?��w,��f.e/¶vQx�~�⮈��
W���G��(�Mi~���d錓��׈����ZU~`�����eEHG �A����[!������@�j���e��j^=�Ι��V��oB��BW f����N��u�w�z�@ �b�"*N����2\Spӯ��#ʝ�r�f2`_�g�	Sv����)��;��Gs;�����A
t䞣��PB�Gg�M�]�����Җ�Q�P8L���2&�Rq>��$D\��� G$y�nv�2��Bj���?��*X��op�4-�?x�@��_��@�f+�h#�
����cV#�'m��L|���UG-**�	/砠_�k��9(��U�Qo�D��jK�̎�[)�����*���'=�fY��uK�I7�r�^_#���eK7 ڝ��UDZV����8���RpV	������H�ml��P*�����ui��*%6���Z+�*4A�d�4w��&���.�'���Êu����<��4Ƿm5|�<������m�93��T+24��E`'>RSZ�Ef'����^�`���6�| i9�{g���sK���/2+��[�{اo*��=bi<�RN�"���؊��f2�Sݽ؜��&x����o��zh�^��%�W}�E���,B|��
,��Oxs5?E��;>U:�軸 ���*""7	ģop57�Wd#���$�/F�Vȓ��-����L:���A}���rg�G�>5emu܃C�P"���/�T����Jͺ8J�C�1U�|�JY�%,~��۰f�����-��3ԏt7��ot�>�[���)^<Gn�Pd?��g#�Ij��cx�h`�k*�V�Vlֱ���Tiͷfeė�qIP��A_`���1��u�i���� �����x��A]��+���u���8*��P�k��G�r~꫈u��Ĺj,R��ɖ�'6��>�F��8u�|����,��P��=����u�Y�����u�wK��vyyl�|��`o;ӻ�ŋ�y	S4�b 3 ��q�S���߷���K�� �WX �[���e���4 W�1X�7�H��#���&����{��Y\>@z�GV9���Ղ)�S�s� b5�8
=���4�2>�:��i��a��Y�N�f��	O[�h+C���$CX8�K�B� !��| }f������C�Ϙ!?-J��a~�3��]��,Y�ʃ*��9=, ���;=�����a?Y��=9ѣ&�i-��ƚ�D�gY��˦u�i�����u"��S�Fy]���r�_,��a+�Š�3�2+m��|��E,::hJj�TX`������VW��n=8���ȥC}��pDI��+L��p�ʒ9&��� ��.N`�#\��!�3��n�~��G��Y��+�sԹK�*E~A\�Y���v�:s��ht�!�z�� Y㇘{��'���2�6l%FYkE-M?/�;�籘��GL'R8\�z�rq�>hI��֒�N���>r�~�4�D�_9���H��+�$���k�}�l�0*'=�6*W�&Z�-�dߖɃh�Y�� ��&�H<�s}�h�ǔ}w ֑ 
ݖ������+>�DZ���Mª01�I}�&8B@77	�"����o��-*����)I��S*)��5���H86�J��S�� �As����V��?�	8Kzu�J���t�"���7���8U�B����S��K��Q�t��á�|̭֨�޿t���S�V��J�~���Ĩ��  �8~O�P�/5>��7�#�^��f�@@8��h@F����<70��0�HL����՜��o�y�I������ 2�QEy�mC�0�V�~_	4B��q�ѿ��X���\��K]�&_��?�I��M����ӎg��[���7���G�x6�.t?����GɟCm2�9Ws-��i�NȜ�c�ĄO� ��~ _Cb�'/E�����3뙇��c�e~QJԀ;c:Z	M�="E���=�y�:��ެѳ��P7���m��4�4ܾ���b5[�lw&�5h2���Y8��6��N��ac����Ȣg���oiH.ڡb<�϶C�8�kޘ��3�\�
J�ܗ2[M9�Ո���������������A���^d Үu��'@�*!�z��}�AM�X�h�Gv�*j�n&Q��γ�a�������_H)"�wG'�l y�/K}[ۇ�g����$
����Nit��{ͰWoH�����~�|���m�s��
�W�xT+^�G����9r�鲑D�����}��~�^��.��Dy����ߑчO�ٹ�
M�#�-�4��k��Be��l//mu�3z��4eN��'ɭ�$��>81h�v��~�{�6���E��ͽ�	(��s��,�^� � �A�Q0|i~��ӓg����k!����[Vo4��ţ���&���7gڅ�F18t�,����l�P��vK�<�)?厯���A�� ��u[<���K6�����ߒ�
h�ۘ����t5n�L�QN{��̌�����@���+A�W:Y#}��i#�2�C�����"��ۥ�+(Dʺ%D���'PN�u�A��,�����o'�VUu
�����s�"Y�����g�}�6��^��P��Y�����R�%�e�������;�w���iVu[R�Z������p�+�FD��8�����2��`�LD.�,�,�YI��Rz9d�j	�z�r�S����sH��+=�Lu��q�x��G(h�n�BO����F��l�����l0S�6�]���0V�%q��@���O�
�I�=�W&�Vΐ,��c$rx��2[�;�}�jH9��?,�h6�s��.���=�Ypa��$���~O8�_QN\��l��p=�0�i@���73���L�)�����u�!��Ʌ��S�k�S�j�����2����ɿq2�1a�fS��->�M6����\n��o�aE5��L�8��`W���o���vA���ˢ�����O�3{46и䶟�$_qE�,������ߡt#Z��8�n��%I��^9����V&)�I����Ì��A��G�lp���A�/q�'j��%��@Mi^3�~M�Hc��W����Uoj�W�r�r���/�7� �$.fk8g �@:��ëa��w�=0�Lj�����
e�2=KP#�/���8�7�R�F{���?F��2��畧�}o6����m:"F� c�t�;��Ur?��"��=�u�c1J���v�==�8q�W��0P�}0���S?�c4�_^�N�7k���3�"z�	��I��LH��_�Q��GLjo̠��m���:Y���=Reʢ��K�[&���Y��nQEy�	����H��_��'��^�R�f�7x;�����g�F]��4^���Bt��<��.R���|ZČ������