��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{�?�!4�.o}��0�m��"��w�#��c�>��3�����U�6�1��_�`i%��u
A���;� ����������.Ȇ*-oh������+��gj&х�	���e���қ:�y�H��K&���o�e��������C1��+�Dnm�+%��Z��N?'�Q�:�%�V�������8]WX<��3.����B'r��G�����a�ٚ5��C).���{=����^�!F���e��SL�~pPmg�\��c��Guخ��O�u�|��٠�ӭ��9�=�&٨�c2X]�颠��"��#�z5���@��Cm�J���,��:�7�{T�h�H��ב�/K���bȿN�j,)��к��q���5zz�;���_�.�a������?�&�uo[�%��SsRwsBOQV�"��4���7~ �)�����	�E���tȲ� �gg<_&"%Z�>C@'���v.r>����/��RQ��K&v���.n��  ���u�+\�81b�I�i' R!o0��ƭ�@����W�r�"^F`�]��a+�*����P5���K�������z��%k)��Hg��_�
.ѹ�����B��}?H�l�By����ǿL�ۍ����E�ȭ�g;3o�~�րa&�R����Ћ{NO�ou9^^/�] ��~a��=�96�zUWd�\	u�o�a���h�~�A��@���mU��L�wpMN��@�b+�8l�S��7͈`l��r\���օр�X�2a������L�89�ް��h]����¤��x�[~�X|y���%*�$����l%� ���X�߆�`3?�ڸٟW��JT~z*�0�O����,����Օ�w���5����a��������HN7���_�d�H4�u�M��{,b|+��nfP�ѴW;pb6� DP{����KZ�(d	�^��N;oJ�;}˻�%�U�Q껔�0��y��1�)W��	��v[ac�k�&Z[��	�}s`���:�?\�[q7�ޅ���|�C�.2̉"�A@���&?��7n�LT!���:���5���lb7��i��j�8F
ýy)\����	���6��p4)&)��~*')؎~�F4Քe�0a��8��1���y1�]2��5�����׳k`hO�A�Tp4L�y�[�itr��R�5'ý��p�3RO�Xs<�����BZo�3ʎ<S�����/1~�Lu`Pyux�+(a@�����y6��搊�denՄw#U�.���w !��G�>c���8��<�Fi=CA00`U�Xуa���}1��s�����b���ω��߱/d-<��G�ܗNB%�9�L�0�r�����<��y�� �N��N/�3�L���
[�B��= ��o$��$�j�\.���.�^CK���{��<�W�3��Fw�(�k�O�dQ9�J��/��O�ֽi�ȼ���U�}Q����Y�l��mbӘ@�f���
���k��H��l[��YM�v%����fU"lo��'�}�y�P��*�h��?�`�
��#���I1�H�@?Mq; �\9�}Pf{�f���N�IŁ�V� 
�V�4֘Ϗ�CY����`���)���b���W���F�}r�:�}|^������CO�+�qe!����$�W��Xz�U�V�^7;%1;�B^m�n���:�G/F� ��'Tse�WZ6��Y�!�·Y�Sx��*U�uR�&w�1��X�]�w�.o�@�g	j_� v)t��oG*y���JF��GP�[��y���qx��	����><./+�mRI�~LL��!�Ы��찃������r�,�;�;�a�@T�������<�{��l�Ǻ�2%����'�g3�
��+��.|(����7|����z�Ȅ��g�m�2�\�-�������D>P"~v[�7A��;d �{���u��ZW%�:k���5�mڝ#v����g���$���pN��7,Z���ͳ�V��;�n��F<z��<�^���mY�WYrs�X~ik
	��e�;�𵦐O�O��d&qns��A���ټX�A����s񑱈�"��{_1��7P%�#�۽Hb{W�Q����OtE�;�pb����c��o�8�oL*�	�����%�w�|����5��)����ݮ�\���<B�§�u�U�� ɖ	�S:�:����,��2������-�>gJ�/�R�Ǻ"Xx�:�'#���: E2 ���d����w�ĉ_�˃���k�@fp���r]^sH��7f�t?j��_�H�k�C�G'1�7�}*@��0�G]F��Tj�
ƾ��Y�X�4
����}wpu��sɟ-��5���vqq?A��0�
�ҷ�W�@>�/?1�B�쬬$�lQ���e�!��LQ�Ry��E.����XQ$]�:����l��l�W*�'���դg�5'f9��"����v6ؓ�#Y毴��G���x7JM�
��3�k#8I�3�o��%{a�� �BӐ��|�A$gIr�)v�� �*�5pW?�����ut>73c��N��)�L�R �f�0��Y,{��I��\�x�#Jʽ��3@<�(⑚I�&�ˈ��K���̟���C	IܙaMФrO�H%�7��[c$���|�E��wɃܔ�]�����(�ʁ�5� 0��)!��_�e@FQ���3D3�W��fqGrMx��7dDU��6��\����S
�f�Y*'BHu�8E[Y������u���o#��HtQ����X�xb�{$
G���]�6$<�>���G�(�.K��ZE���zY��b'��-� ?o/U[T����R��m`w��8��vƩ��3��_�$QX8�م�9 &=�cQ	��~��e�:z��)������ScѡĹ-u�7��B�M̬�o�,U�
��݋jE]�0���I~"W]x�F|���ԫdR���n��L�JH�<I�J	���M�3��;����t}�%'���[�z�Dh�R�h4	��Z�ڏ�����#_�=-X�!~(�Zi��G�αfˬ� ����&�ўX=�*;?��a������z���E�������U�! ��~�abe�/��& &�L\�~`g�+$�9�Cz��*��#ն%-�X�ް��A?c�֒��C�mv��{�L\��MD,/��ך���T�5G�/`"�iL�V^��l�������('r�^�д+�Qֈ���<�_o��,��C��$��l�����}����S���f��L�v�l��9��,X�5V^e*������	��HQIjT#� Zo��d\�|�TW��4�r%�?����ēq�+��P�6 !���̡��Ty�l����"֏���S�[�
��'��6#2L���D�T:/hF5�)��K3�ç᪝�p�&��TN����9h�T�@�v���b�?�4�j/�\��B���sZ܄��=�M�H�<���ۥ|8
��Lb5+Um����A!�~�\2����Y깫������A���s$,���Pb���H���(��d��9��Ӫ���AFސ����Ӱ\�\(7�*^/S�, A���/޴��W����J��$D�.�u�� ��O���k+c}Ji�ޤ����Cނ�
h=\�X��D=�6�s�,ؤ�:��zWo�/7���i1O_ E���V$ɾ��sj�y�Uf3�Q%#��/Y�?�P��+x���9;@K�H���
���UWe3J�̀�D��LF75Uؐ�l���ֲ�:�_ꎊ߁wE^x�>B�3�3Z>�|�c&]�4MA
I-�N�[���ʺ/�2>^}$bZ��OS��xu�I��K�`�z����Z7�P)����n;�ue�/����������U����ٲp�|E�h�)s�R�u��4eb:�mɹ��Y���(�������"��6Q&q���)��Kv�<\��钞{bu��B���͸���`����M���*Q�?e�'��}%�:|�v�����T�kJ��S� �"��G*G"�T�7�e��.��P�G��r���+���^��gd�����|�ow���S!���Q�� �	+�ٖOc���u�C3(�+ӂ���J�C��ģO힥��I�P��f��/�X�n�1�CL����kzZ��c K#�~`�\A~|#yO���.N����_�D�Ӓ"�#"ހ�c1���a'S�Fm.]�ˋ��������f������Z���)�-}@�*���
��[b�6��A�v����`�o�&G��6��.dP�j�+f��	ژPyZ"��-���.�h�~�k���p/_���҉�ꬡf� ��0e#0;(LO��PH:��쉪:|�� ��tM$�V��0�vt��̪l�¦�ՙ���r���8y7)����)0Ъ�2b�d'�UƸ8��,�q��V;5^�s�$4
��mA�: ��uL�X�����GW��::}w�$1�[�vq�>T"��X�Z����Ɩ[��P��������
�̟�=�1.$9A5�� �ĸ���ˉ�<�w�A$3���W�t����
���>�uA"���?VV�S�Z�ߚ���޿U{c�߻*;��C�������������N���C[Y��8^�+�����N4f���Ua�N\�U�U��7R�_���x�r�p?aq*�x/�!?��17�(��uG��B�]�lL���c�GOB7��B�!��P�g��9�"�5"� �C�1�U�'E�%V���;�VZ6p�,j�}؎�B�rX#Zג}�O��*�3�6/zD)c:������{4�[l�s����I���/(�#�D�Ȫ�9��wR�u;��.v(=��Y��
|t��Nn����Q�=R�gDi�D���d�D�`?�;�@�&�m�:�n��I:���R��c��)W�K�T�����Rmݡ����TA���������g=����;PW��NW�}�]�������8�?Hi��h�Jn�*چ/��@�48���2��-�T+X���(���X ������f�u���� �S�G�d.w�(K���!�{Ih&�q��Oc�/!0V3�`c=kK������5�5{R�]e�P����MP�Xm4�~-nS�C9�� F}_\U��%�V|��D��hl� ��QXY���%�W� hn�Yd`��da��q;���q׵�p��Q�����"	a�i9�����?�Q�+�$:@a����v�0���yV���6&��HX���&ΌAsSI{�@���%��;
 �*��˩{�
�����k�~`�%/۪�J�N
�~�J�N�f���4Lo���]��3���`*Y��2=t�����
¡ԃ@��4!v��Б��dkD�-bs�o)9��v�R�5Z�,��?�aQy�Z�tP�����~:��n���-�ض38D�|N�v�f�H�eM��R��+Ô\�b�{��<�� �[ڞ=�N�/�J=�P<)J���_��UO��� �3������]�� �798�Fɱ�f��ݗ�3BqS�\q3G8�XӄlZ=;�!�c�xӋ�xS��@9raCb*\ ���~��=�hTi5c�A/�ҶH�Xx���Ѡr4�rZ$=������b�������-O�ZT�4���8�����g�����N�*��q'�ZH,⥀�VJ�.���cv{�P�z�U�jӵ�v��{P

MR5lX���q��kq�_a.�0�+�K@-�098^8�@�cb�d�p��ԬN�_�ԋ�k�� l�}��!X�m�+�6o�oX�:0�[7m)Xh|GD�O�����9F��Q�ٟ����\D��s&|�]q13ED�}�Z�_����HXz���U�<N1���!�9d2h�ˎ
�G��
|hI���X��:!��戂�O�O6��������u����e�+��c��YhF�b��%�N;Y�On�r�lN1�9�N��w��=�X�F<f���8*�� �s�n�vX�QH92�^Z~���\^����$�g��7�����1dv�!�V����J__������J@�*��z����2ລ5�	�8�]Uk�|�A~��taL�5q��eB)ץi���#�.�J2l��鬌p�G�+�]'��+7���<W]�P�C.�xԡ��0^VG��Kin\�b�FH�A�q蔄�k��.�1� (�G�sN�A�o�yTioq�F�8�t��l(����\��X� �<ߠ4��E�
"�8Z�pg?��{��?&�Ì��$��o��}�ʰ��߇I�pM��^��J-�g�?j.s��*|�E�kY'�q�K��'�-f"��w�\Lu>#,��l����J�A�&�j�{`��>��C����"w�������!y�w��؞��U�]���P�'��A�Y8D*��z�<��sR�]F9�Z��Y�A��څ�̓�Q��r�l���L����0�1�5R�K��Ɵ1���	�������P�u���T4��i�!��e2�Z�'��T.��82�����t��`aFY3^�I��nh��fan�nx�u���þ�<ON-n���<�R_��8���g���y�`�ҭt�/��bO�x^�����0��þ�2�=��z7!�����Q
e�J~�Q�<e� �c��P�ޓ]v����[�`~��%�}��
�]|2��H7^T�v�l�ٞ��t<����I����Moޗ�4�y�3.�Ws)v�8�]����FyS��ǡ/� �E��6���T	���/��a	���{u��]���i�Jw�}���8PC�'9^�8��e}�;-(��b��B+7�f���A� j��;2́+/�C�OF�^fG���/: ���(�&��ѯ�:�y��&?�d9��:��}��X�l�9�>�U�۵��m~���M����l�&H ���d�R����^-�Z�/#S�_s�`N�T��KD{�U㊙�7��x��Eh8I�?mh�!r:�����y�.�86L(�A�&���%iD���t��h�)�}S���ߓp���-������1u�Z���5\d���x�����b��@����p���f7�~��\�o��	۲�9s]���e�C��X��[�
�(m��oꌔ+y��V�V��Ќ|�s�@��>^�_��c_����Y&�$���:;h���;��]���׊�B�O���wp�#R9�p~#D�
	M������v�0�M�4d���,����9#@��,}C7�IZ��ӏ\�	�q�$�۪h�,��JDy���q�7���u]��b��s[1��q�p�L�Vv�㍟�`�y�-
ݮ*a8?Ṱ�ko`/�����t�!"#(�-�u��>1�9Vlkz�02ȶ�7d�aFLEّ�o�%�P���ɉ�ǩw���'���+���[+B����G��_���c�o�HoT���+�P�%T�'�p���
��n�q*yPV�I��Tp�g	@�v�a,~Ck�p'�m�����V~�n�8;x�|>@�o�[��Ҍ�s>r:
D2����VojuB��W�6b1~�?蓤��}�o�}��2�p3&dNM�?��o�����۳U2J���7r�H����3�QM�уZ+w#��<�D�R�%���X>8����PXw㜸^��`�)�����	�J�:��I��	�ޕrY�w��z�;���[��h��+foFI��d6̪�|~%��A�s7�ed�'y���v���"^YV��Y��YIjJ��Ȟ�H�l�)�	����� i!�	 7C����7/Zot)�SVH��E����Y+�@g]gJ��L\�=���j�T�Ti�ձ׀!6:^���VoXƠ7�J����ѣ��F��Ԁ�qAD�e��n�ŏ]���㏓Y� �(�Pf �6�c×!0�Z�&��䁶��py���ˁ��i���ι���Ib����l���ğyg�������A�M"��d�A�E��"�V8X�c��F;(��C��yi�M	�����i3����\�� @&%��A�<5@�'�*m����.o��3�_i��qp�
u!���;�����2~5���t�I.r tP,旡��H�'� R!l^��
��.��dx��~N���d��aO�F(�Y!��6ߖ�-��p\'��PL���f�6h�2�@FŌ{s��8ՄQP��_�����,V!�Q8J��{�]�yBoyfM~��jX�蜛E��V���F�O[���i1l�`��_u~� ҄�'�5����V�ޟ<�@R��eޯ�h��a��N��[l�����uqg��F�`#�vG@R5.3�e��%6���	�|�ױ�k{�l ���H O˜Ŭ�b�ļ�x��{<�,��Q];gq�8!��;��TqN񼂇��Q
�;$�T�6�2�XnH��A�j���.X�|�r+	�ʓz���|4T��O:wq��3HhjCoG��n5I����+�e���kKG�3*�c�3�?
�
�e'FF�3�Ր�f�(TE�Bq&]�F��p׸D�W�R� �.�Òk�wp�G������\7�t�J�xR�B&ncv�NXn1%�b�����h�?�U4�?� i6 �� iiV��vmp������3��d���EY ��R��T͜���w#-���j<Q��f�ϚG=鷨w���Ԓ��e��v�wZ�T�︺��hq�V����L��lQ����/¦Hm�$]��S�������(�.��g��@�o^��2 ��lL�ӆĄ��B�v<	�t���|��Y}.v���D�]���f:5?eT,�$I�@;U�.C`+�X���2��Oe�t�z��g�����_ɍ���L����_��əY,4�4�f'Y�8q��ٔk q7,���颗�*��#�%��'��9��u�VQ�۷;A�z�x�U�%���j�u�8��gTWN���HB���(��'�F]*[3�ȼ���H�v��;k��פ_][+qTWc_���m��se�����k����v��v�v�,R��o�����08k��0��N�9�U��:IY7=%�e�����#�q�H��)YLκ���Z��ڏ��ݦr�mS�z���G<(P�j�B)�j8���_��=�g"��;�	�V��mp4A�_�^0��rā
#����F �;+֌hN_?5�?��:�ߩ�n *.:)Gv������OK��tT����� J1�W�G�[��HD�?��������<�>��0�����a��_g���v��=|dC��JU#�r�d��������BN]��n�U�u	ԏa9�$�78n�.�f�<�?I`sl3hM")�����Z�S��hx�u�]�W�P��8�l�-~�h����^'���O; X�JbCD�񠫤�K�"����8ْ�������]�� :o�&'�q$e��L��6<���
����X����,o�4�?&��]WN���w�s�Ν� ��[`��5��Rw_�'�U���[pߓn2��y��J��c�Z�^]\�6���`/K�z��y/k���������EW�^����G�ŀh�i��p��tz�_C�ؾ4��w[��_�hsr�Eͦ����f�<{���� �A(���o=��+gPӣ<��e��������p���5Kw˳������_���d|�����uefo G�B�*Þ3<���%�2��\PJ�|b@H��16ˡ�Xsίm��L��v���������o�*4鸍
�<~_[l��I7$:��f�+�@�i��y�GA-�^�C