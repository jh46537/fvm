��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_y�Cz3U��� X�D^{�lW%�:�j
&�tN�4O��a�]�;;����L�S~��%y�A�tw��d���2/xT�e?&�
�W�@���.��+�l^[vhw)Z����-���=�(ݍ\���Ֆ�(�H��Un�����PT�Ϊ�f�aE\��@�ߋ�D���`�w�8�
#��0�A
�~�������ۘp�u�
u�Ծ�~�U72��v��AQ)B@�~Da��U����ٹ�w�$�_�K�	��*��;d�w�p%F����_�Gw-��6CR�dk(���j�1>-����L=�b�2���E�8D�)�:
{��`ƞ<���dѭ�*�/m[ ?��}�=�vA[6�H
�gޥ��t�Iew�O�)�1�.���iu�Oqt1�X_4]~O�d�e��DOf�?�AW�ˣ�8�5��{��פ����s�T�>C#�[�=D�o�/��!%y�zׇ�������d��u14�{�	���?6���V���YYw��~��a��Ӫ���l2o3�Ÿ	\�����H�#V����$���N>}⺴�rD�l^��zr��K���M�~9�
�yJ��NEN�j��oō��"���Vt�fU�9�2����h������u�O��	�YD��#�ˣ剧���Q����-�u���F���c�(�c��Gr�aֈ��mia�Kj^J�m���#)y�7�"a�*��^���]_g�� �K7F���y4I��H�3��TB�.��!f����k�)ɺU?����'��n��%�u���v�*��)���(��j՝����J�4��7�J/�؄��3;��q{�iJ"�35Ԟ ;�t<F���w{�/T���ً&W���J~�M]���U�	�tJ�G���L;�hArI[�v�*���j}��N&
�z��J6��v��/���>�'����4\�5�H��Cn0��yz�z��v�r���v�8I?��e�	��rzp�ݬ1��Ac{w�]
P�=��}-��s�Ze�fk<���e��[�px:/}LwQ�iɤx%�GҸAg~�6������݈z��|]�9��D$6�Q��vQr:���k4�B�|��<Z`I:��$p�����ψ�R+��Y~�O����C|���4�q߇�~ ��9�ݭ�}�iUu�0�2	�m��|
�=�j~����ݬ��������a�3�-�>Pӭ��������?���2Gٲ�U]�j��D�ꐌ`i��a��Tq�kw�bV����ݑ�`;�*�7u�
�*hV�����mטQ��H���:��w�A�8;��M���}�*���[�ۍ�5����"�
L�Ղ��O��:�7
�|�!m7����=��[����5+�`�זƅ҂�"����볫q���LoI�߯nP.qɃU��ݍ�t����,\EG��B�9`�F���)�l��k ���N�kB��Pw:d�]2Η�{ʖ�l�~d�"dYd��\��}e W<=.s#/6����yV,y
�+f�������(@j&��u��T2?ă���02�K�~�TrDL�~|ΫA{4�hyY�����&�8�	8��S��fOO
;�wD�.��c���9�����.�n�����}O�z`M�K���+%!�����Yת�/f/�$���ǹ����(ar�m ���Mp��حY�r<J����$j�kx�z^�ulW9ˀ�U��s+�Ѹw(Q��)�p��%���!Si��ܣ���O�%��3BzQd�v�%ky�"	Z&����"19�ػM�o9�����P<��򳰊q��Ҹ�)o��CaDcς�E��}㌉�ى���ݽ�}��C��L�J\��bA�0c�AM������+���V�,R��@0x�P��*���WѪ=`��9�(4+�����n�0�N�Z+sG��;1���E����Ȇ���8�k�Qd�tK,ĺ�u�H���30_C$��FdDN����C�%�؁g/��Dr�����<�>D^���j����KG]��D���#���4������x+~�4~���VX��	��X�5//$pe�WX�S��]�,i���9_�O�H%���{:���P /|v���~E.fe�6�q% V���1�L�~�bB�u�:��	�?�$"^�A��j��Aw���Yѱ�=<��l���7L^y�(���S̴HF/=���.���|�J˧rt��b����ٖ�tF?p����Svx<7����>���M��ʙ!�[ƀ w,BcZǆƿ�˦�J��ơ_wb��;�y4�q��R��:�M�T���a�5�M)�Ɓx`��N��֝ɯ��4쇂�[�C���^?���%�o?gei��[�.����-�4�|j�j�x��#���1�3أ"dǕ=v��zĀ^q;�1��!,.��&�-��� ������K��{�PP&