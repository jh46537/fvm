// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J3V7eKyEK3AbjKD3mpSQ1JDqLJOHPVLZBWUuq8GiiI9k6kCAdXHmPqR9qfeXfAKl
Pwk6zdy2ctWPC0f7m4Xzv+HEXBxOaQclMAOhnlPGjcROtd1w6KHJKR3+r+XRaTWo
wAVfoy3urn7lSPyU8dhqgewoDD6M2+k9Ytt8MBjKCd4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5840)
shRIBl+7abtiz9cUrIhy/LnRZ8AAtuwz1ZbdH5RVDldOPN6FwyIT9fIS6j5yQodQ
lWXmZxyey05Gfnr/TgDLBzMbGV0psqSRJ5ZMPaQX+d6mKZFOeW3eSZe7/rW3pwM2
Kaya7B5NEJAMdgK3W4KMILH4KeATLHYHwd2frr9nGMiea311GsBBuI/zb/KbK/eV
No/KqeRbAH7d2r4vAJ/OidkqMnxkfx8TZ65EpMh7t9C7uLQ6cmefZQKsIO//KasT
UoMbNc80tXU+b03Fn/kKM4x+EIgWgBV71aN8cXDe4jGNsHvH4DgPEw0oPLq1GH6i
wp4No20Tr4qMeFrqzS8wPvNnRJwaTg/Yat8JTlsMcdg3WjomlfGfNCxZwXtwagd4
uPQBPkNel4IoUE6nt7jjbuKZjPlwJiszhT+DZpT7/AOatBP781G7Gk2bdjmHei9C
EEWqwv98ycQO8xrkHMaYQa5Qrt50OPq/Ju8jAEOzTknf04sPKmMNPBdeW8DDBw3C
NwWy8iwOAGQzS4MLpKyRgfwErZaJoGlkADqKw/TECzaVt+qYNEyJ/DijKHp6Ln5u
uYK24I9Z05lQqvSNgslWTo1JHXsT+VpKIPqds4Hpr6YKo21pXEA+iahMbmpcvUow
4tjL/1OVGWrQi+LafOD3i5UOSKF9mlfx7pgjUF4xZ6XNE3/Fw9O/5VkWfMr8xa1N
wWeTu6Mt6VfBwjqYNqem8jl7Z0dRHtWYHrPMik/SGt2LOqxoJ6SDHVLw0B4QrK/2
PtOtIY2mAn2e6/6wnTNYjHRrP6hXPiZmyPQUqlkKIAy67JGcOMLyDeFbeLCHYWAv
0psWsB/LXPKNfs7tcruFtEVzgXuxoZOiTUdDdJlRHAN+yz/oXtrZVePv3rOUgh/G
jWMWnS6ivBecfH0V4Bds8bQprake8xhfMrg99P1PgQU1J2tGOlpK3mV//MdFxMZU
VRTP5omf6+9YAubBEokJ+botCGO5h/lTBS3NoC8RifPurMLlkMzKs4LJlFjJ8NS9
tVxBJ+Pq/FDeH9+FHH2mxbscxWLegF/LWPI0e+Z8jXPicUMh1usIjMTv31PGZ6Dz
tAS7X0NhyxGwbDa4a5Xl3L8iNi5AAZ3x5mIqGzh5sHGrz8ZwNF4d1yxzVVdfl1xu
gSq5NrI3S3p9pnjCp1Gx6aIbz2uXHUcAuGzOH8JCHgn/QdluwlHf41iiiV8VTuJI
Iai2SEcUfZ0vWKR2DLCxVxouZL4qfOokDTMQ+PfsYzc3POEDnY7m/mTP2qOLZLqC
ODkZQMy7RFmMikxfl4rAk7KMSBzo9/0wGW1H+bvcvIrwTqSh79O4zbIGICaku26W
GdbEFT7M95eKgtmA2ufMoAu1pEGuCxBvumTHhRaxWYGhuE8ATkomutKztj51thvy
BWC1dLy/Mf4FpPl85IjuqE3gUeWgbz46TGxIaA3pgigjYE+pXIC3ADL84wmHADjY
GCi5A0xV5xbDsS5KAjq6/+clrp5v1SrEq2ZQ8IqaVWvhle/izOmbnGGkvcU/TAY3
tJmEi69yQ9xoBVqXBmO05aP6xiTYRnQm57H55P7+Ar+EIgMeIZRmrfrTqmkVwLx0
rcK5tg/gG0W2Qqaq3fMraI4kSjvuTF7JeI2mLuPwntVXvc7bY43HHyJizQKN+Pfu
am0PAGf9XIHHW54aZyIAQpe31ZhsOBPUNkqEm9qf3ZN/fYLbGmnSySlEy0rMxYtc
knORWOsEaDDUnTf6IGGSGj9jRvTscyFsQ7VwMEDU3qPTt0zuYl3dK5CZXzZ6Q9qd
1+BYTQpdWKFqrPMl4HHQJF771/B7sEHgRPCw5QpozH0dw6ZGJJVtp4GyQvvH8nl5
hPveqGztsOamM3k5MfSl/r5MZJalIynQW9GET68DA8M7YYxApOXceqt+yGJliwCO
ZZNkSxBL8wYv+mcIgigpbY2Wo+XyosL5a+6vSyc68aBhpcgpiiCH1VA8ObftYpfF
Prpe8ZikrtoehIt3HKp9raa7ztN+CPNQKsTv7XWXJcm296FlPHlMhbuHMvmGtjZY
Rkfu6YDDR/Enn3trMgTA8G/7+VxPR8JayEYz9aweNoK8La1iJko666O9w6F6gpz7
H1whYsHfmaa99WXid/YK7fHnHgmF8Nj/vMmDe+YPedtZtlgIxGB5I9ceG8WuHvfl
Ms6keZn5qBJyLs/vF47QSQnWRv0t67POXolMYymWsjlx5+1uwq/ADRnIXSJHwV37
DYvUMucz3uN1/G3WHm6AUEC+J44dLPrvNRieRkFQuNifpAmISh5+SAmYOF1dDIYa
x2bCxIyd00qRrmTvmTd2WpGke3DSXPXvL/hmsahpquayMHQS6pVmNB+EkI2L9vhs
4OhfPAAR8mTrK2GpFf4/NdRac8R8KgklHWNeDVB8jAPwoaUtIL27izW9Nim6OINW
M+22OmSrFr/Y5Di0OUOE3qhh+IQ0roleuaSVGWJpDtyNdhPYf33FQxWX4ed86JMR
nQMRcHUwxb0telrMCfnIskeoYg5Qz9DiVIiKZ/eISInj9mQ2/7ulB872LyVKA8/y
78OdgRqXiiqa4nu6dPRbjqRy6meSv4g+0yrfQaZm+JjdDKuu4TyVBrhV6RIobgt8
MGKsZpAajqhgvHfeumV5Dvu7wD3OEstCiVZqKxVLSfa/pTraiGH4B+b+xqEsJsZt
nstUSKM2yTlQRYbsGO5/t/lfissEvbayC2pLBcQHEUVrROp9W5wRUz3reF40yPfP
WzQ3Km3meeNvd2yX4E4kytR+xhkJKbXQtp+D/2lsmr+nCDb6t9mxUKAdA+bJOvbL
JIH3Tx/sKwXhMlj305XvJhPUPtuPLJknatXE97Nze889TyxwNiJfef2GIItAmXD0
LyJzXxIFf12rZ/gx1wYCNn4xD9ZLyeYtcbXaonRvpZVxp7+pdfSYN1xBA460zLsZ
SqoYz2KacFSGsmJGA7S7qkDNGXDFDw5ZNzqENBByeXr/+QhZ1X6eFZq0MNg3p9gm
NVAAB/Ovz/QGkplgVgmMAZBYs7w+Ca/4o+q7nQ9PMvqwL1tj3TKjOCKP099rumOy
3SAmx3y6br7sM7pFmFbunHtULis/jmjLJ2RQzhVRj+qZca6VIz1vr6FI0ynupdqB
A6qaw5YcYNwwis68w0Sv0ntE+mBJX4ZlDHyayRfZNZNFQ7MJ/QUR3zWq5IjRw95T
5BGydS5zCIcumx+1zu3EtO/Rf4wMxxlCuuMyItX331msOB+aMO4rgTdhwcJcipJM
VUWKKcBTtDR4UZZUaTIZP1FshGbuBTuW9azCQ4vdCC26M26hlQRPNY6P+5z1Q3wM
CXT1WRiZ1oS8WJW3MDhZRm1G7RsNRV27bI+X9/laXKtNykHhmF1l4xce/DEaCm9g
wmnNFAkgXlolhQXciMmZojztcz3tP7IyswulzPsuF6fm0Wdim5PlnBo7ro5TwVCi
n18dSYJqlb318bEHtj/6qYRqj0wwwf/LiUQlWfn2QONLuairFCHxpRvO17Ip3PH5
hT9/nOxR1MlChujRBLSXsipJuJHaNoarTWJQ6i3T3Pv4uUybpKsP5KT+WnKxMR3D
bmQC+WEcqetQTEzl5zP5UfSwJC188uaYNFubSMengmO4Z2WurHPuEaPmW4p5+CN9
1Rw2L4f7BM2wDJi14nDU/sZZtspvTykEeiZSVUMPG/smaWcN/H98peisZuBALR/D
/2dTgoPJmFKpMckFo6hafmqXhWk5Wtak+Z9UrCFr7tkCQpHJ5wn9JptbGXpv17hT
ijqxfLmmbnfcwm1BkSXvMIV7TUfFDEPCbCxQQm4aoN4U3Y8sOq7x71c35NWJ3YhU
1osDioPoxwcqixbk4qvw7iEukbPImv9Up+YDIp4XNK1iq41LM4ECePJhl/WHPJXx
WXEoyB1SwMS31okOAmJ0xHkZkAj9ZybJC1bWuYNkspWOHFwgTghRHiUPOY1vdtre
FQ8fITqcOkwPFISRgU1uki/ufius9yY0fR/qtg410I7VgGUDveqA9eTcV36xrLpG
zMHo9uCKdSxlrJ6POzffKVMHyOOqUTpDUns0fzEolif880+eolpbdRBp2dNxgP9O
87f0bnK0SavyXpvO9n0LVgqRNGwaQcKmgDcJ74DhpkOmMO5yoaQhHT5cREccgmU/
wcJEnicPb9YL0qKh38lc8EY9Flo33IOkGLIr+W3dhfk+4NrZCbu4NWb0ES3a8eXY
DReq5ibNqvK/A+EeHlfDR8RrX/JlqxLfv4GEvaPlAcR24i8zWfiSUzDadS0pFCq2
mcR3bOrOeqF0BIH6An9KXNE32/9L6b12l0kTUL2z2j+c0tmLUA3qzScFM3dWjGxv
qVkTNcRXlrOCR6CETBlwdh1kPwOE+AAIQRWMrohIHxMO2Ixv9LxGPznWSG8iS+iY
ppZdN+hbP91zmxO5XKInCglgGf09q6RI9/yJByeKxiViO9M1xf3JFzfksL4bPgSN
ZLaRBit237j0x4Wa3LUh3GF+dVy+R/fmyar4Dyhg3NDg81VfFfrqiNqPDgA+RmJR
/seOx1h3z9J9AZqhNuNLP96MpW2bFs1PQmCmF+RheeHORz+M1TpjJbkWDrXJVrpS
EzV9UgJqCnbVk3H0PGaIL4mNYU6xMgLZmbwtdlFzNGSbgjcwNaVBOvqtWSy+O39m
WAZB/WzzSYSmJDetJPwKX7nnzqGhAOvyz9OYg+TRA/eZWVFHtxu14J3SDShjiSkD
kdUoYZI2GeWo8GwwTyOnSmr14PojxER60tX7rZVMpRmhxh6VuiEgwldQ2Ps19qVu
3e6LcsX49DBu6t+XcJOdwNqnS2q0MzOHV5CZail17QRp+uSouRfr4X3h8c187onE
wP1R9XVZ0v8eRfEBzFkiU5uzvX7HntbScebzDuHNJMlvyE1JBPq9r63lsygCdfXG
RyYWkCLkCKwQPs+ZdqwbxVc+Q6PfsdDzInmyTQXQ2nqzz0FB/0DFwiztIl2k4Spz
m4hMDvAHuzhfCK+fKQaDn+2n/Ak4sZaMZMyYZdGAPeDJu0FAU7JYQRUDa9yvQC34
sox9qbeYoPnGK6oUy+gBBgLScRtqp58HmhIV6xgbuYwYjXRJJHF+H2UwQReYTyi0
zNVs4sKE0LPRlRN2eIxR7c4k9qwzPZgPIA58LOrN+qGCKMgEQkaW5+soZS/EL4vG
qLup9WRugh2xvNINvj1ZqLW35wENV6jCl4uzScxOm0uNvNvaHEIJyZlHPftLQK8v
9ajg476RZI/we3UoRkEDPiqKGaMj1KpxOGvFHomt5Hf7se7J7Hh60jFTBqTEEp2t
hcPSNSGA3UtqhlYoaDAtUkzdFG148qgos2OLRdFuyxbW+g2HqXq9/TtudVUzovSo
rTCNjSkbIN4sxvVOFCRExbWut2HAule762YD6aodA2EHvaHKbKnZ9UodvddGqLJu
3XVU8XV+0nD1hJHDan3gnZIM5QA0Nb+2F/QYuRUc3Sf/X37+m/FWSAegtGLz40ON
ui52tVpnbJ2M6n212SxDmwHN79Ylr094xQ2vjbT3Fs3S7vFn2tt3ASA1RrKVkZCo
6hfbtetL2RMG2uswkwkb6KVCu0ag2aZnwGSGf/Sg69POJssaEpu5VNuEllZiHAeB
LUcfQcshQ61ef4XqAdwSdFNDgUMXP2PlKsNsGTbYj7ZthPWK66MOJJa/ggSgOPnD
yaxtA2p4Svqbxbj9Uc9AdbXXXKL3af5Xm6acDamjFCvGOs+jMmsPfBc8DfqcoYpL
jqPhWed898DCsRScoCJ4LIH+SCeKJ/u1picWGRpnzaxsywyHmTGCK4f/gR2fHrdv
bxv4NF28XAq6uir5SyyQB5R1rzQTjkHYLIBkNgDNuXyNkIGrYhT0y/QBMez7fZIl
cytpXvFTuqMy92YmrHjDsAtzi+Vd8HZqqqE6QzPqigIPg2QtV1Vl8GMaPCy0b23Y
jLuTm6CfNICKvNkpVHEuBoeSW3fIuVsM+GuMsGgdX9SVTyIwD13mdA3vK86B4nc8
e+SlajqKJI02VXhENY2etNveSmPIxca3joeh4K3X7dQb8gXSdAtve2SaYHMJ8bgQ
QF4t+b00L24K1gGL8T/rlez2KyPOOayuCp0w9d4eng0/g4Id0UKmR0Ntykqo/cYJ
fZRQmcb2n1AU4pg05S9Br8txlsFqzaq75/Csg64lPcwK/TBK1ESCJqsDEx8k0MRp
F2DmIWwLezLrprtKUtx6wem4705/GQ6jAUcFM4lZg7+95ljbczj6HZYScEVFuZ/1
taXMX2ul+NlnR4+366wSLuwjI3zG6tkp9vE+mFgGUfyRgX2eDedX8F9r5GWdOrT3
JJGZeKZe4xkTMzctTL5UxIhtsy+7PNc8omynX25Lzfl+CMHNT1jspP5Pi63tbghs
9SKUJmKIK7KCGhHBz6zLNAdLDN0v9tUqn/RHRnXNxabHJVqLyqF3CBS8skQondgJ
2s3oIHd2vpiXGD6iRSeFltAyQUooCbxrdj9Gif1iZKGguFdNVe0WOh9+BE0iXuhu
BaalqVYUOXX1zOEEGUS4AEItv7J4K/Wap4ZqErsU1a3L5cro8yON1DJ5tq8lRas2
Xr7FQgIRKOWTNGGPPWBSvH1N6d0ee6+7toufd0kAkvSC023r4KS5ppGbPbsUnk/E
ThRcvRoWuFchieKjlknIJrMrBoV7w2qSGrrUcso/JgZJPD7oUmE2WSpQz4afMOZU
Ue1Lo/bxoQy8KyqltXwrgmdt7WZI0O4i2MFIYz0Yb7uXKYd0VhHVg2ffFyFNiTtx
p7WcecaoLIDhoRRuf60LpRjjUE9BC/qXchtGMJoVLLx9l9DmI6CC61nPBgKYmACW
mVenE1JHaSIpNaxEB1NcvQvTEjVvTT1N+K6uuZi/LIfFrlZjkesP9YgLjwabliN7
0KJCYLOmCaP0AZcNZ8jb1YU+QZsjKnGjtxXjYUVfH0Z1rdUBKrAxb2DjMH+RAya1
e4gIdAFX4yepwKRj24UM6n6lt6tgBpPX94f6KSG6cI7Z27LKy1bkvfqg6izoBbLU
0lRrUtyu9VgNsfT+Tic76D/gBvv/tOVtT3XtQWOx5s5RPYziAJY7htlufPzLJskC
RZBh2FPQG9yL3NJXM9Knj3fubrwL+3j0p9TTQWOW4f5engRR9PYpzPkqyTnfxRLj
3cMNaf5tFMNVPF5M/Anv6SCJwvMIBvvXprYIiK7NfcKWUCV/v2UNjyW4b3YfHEjL
+oYz+F1grCL3b2H3Z7qoL+Shz54Tyb0wbU65Jyrka602I53hGYxCWs6SRY71JVjW
f+B7B32tkYGuiQZggSZd3pd/pFw/5VsXhDehLFhmGjj2yrXa0fh7/U3NvxuULiIP
FGSZgJ49Weg/FB/lPchoIU53NWnmXAWqs1rd5umUdBoaMsA1YZ8zlbhoZ7V/6/Hb
ZUDb7j6OweRnQZMXZQ7/wt3Mny0GmMrjpwAOcArVs4fEEPgasWy64uMZ8kne+b9E
MAHXuq9bMVvAeu0OmD9ZqEJmyByua+E5unwe0JIk5XdrhDZVy1MboLRCK/LjYUO6
uVTV6giMwrOPFI91HM9j7KyO6fVViGKVFDBP8lYwWVVEUVbCH9Ly5BtFZxibVd/A
UDUjMJE16Gua8imQrIK2CQf83WUTmYh9kbSqhzQD3FpRUS/05KRAOA5Pzy4d1swS
ad4AJPByPr6k9ZtBwKKGH0qLP3pFeM7RM2/i0t4kJT/E1gaXTf6dKtxycRijgE8e
ADeI2ra8cUFhbr4JkQckMw8s+8WilevyWyv9S43mxV8=
`pragma protect end_protected
