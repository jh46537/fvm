��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{���b�e��_�@�*��Ht�'�>��j��vK0�N�z��D5|_�-�ڐۖ��0$5��=[��ЊE��6s��k��Ƕ_�V���gxy�=і!=I��bvZb7�������qw�^ͣ!��H����֬�T���Ƒt�MrW�殺!>C��� ����ߖ�܄\������Ȩ�/���4>�R�g���� 1۰����2RKLE���FdH����4g�Kw��T�����$�Do�3ᴞ�?�$M��cba���DU`k�&�V\��An��G植'�i����ź~@i}.K�4%H��?D��)_^J@���u����Oby���4��v��;1��q���"����d�g�u����1�2�,���d ���ޜv^�j(�7�JR)fhg����ycpAF�e8*������6ST$rLP�d�r���4Q���ۡK�x��E��n�ſ2���A��O���h�}�^�,���h��
��٨Z�Z�a�G3��81=1�ލ�OH�d��7�"��W�
���O�A�fv'�ae��49ȉ���D}1���f{�l(2�d��_�����I޶BĤƙ��hHC � .��i��\��Dx@�f��a�ڐ_6>G�N���y��ߚ=�%ճ�O�4��&�$JY?�6x��YcB��t���_����y!�q&SY�^l�O*F�� ǽ��������H�T�"��=8��_�����JwD�P6�_�{U�	X�n&����y����9��l���Œu��*B�b<��RD�}�20{UlMR��P�v��T�m�n�A��d �KoI+��6�wGOŃY�
7G�.���~BS
.a|�tJ�|����od9�+9�G�"�L��ucU���Z>�VۿNF8�t�o�6Qz��, >?%�L��1�r�޳>�A}Q����������u��&�����A���' w�\�f��P����&!Īb���	I��ju�#Kb���3qnI��^3�t�Ꙇ\n[ˬʄ��!"��-Ŭ�m'.V̝Z���OKv Q�/��1���Q+̐��JU�a�νEZ-d@W6��	^:��A�� �&Q� j���F+�=�L}X�8�A)l52Qa��7?CP�N�E6�" ��\�I|)j��hg�S&7�D��V@?(v@E��sk���!]#��;{���&(/�`8)}A�Jd��I��vR7P�������f�����#�>o~I�gι��t|۶�B�Z�j��}h�-�6�p��(�t�2O~r�KiMA�8w�x����k>k�t�����پ����N���*�k�9��5d���= siDs;�����M�y�[W[��]�<	?K��1|S�v�Rr�<LohO��@W;�2����uo��<�� �4\4*������$�h1N��0���V+c(T46���6��3�bV�;�2���SӴ���	T��x�+)	���M$���r��=�I�j�����k6�1��z3j�Vj�*�!ַ-{�|�㚯�!�<�%�\CJ9������0�v^CAn蝱����)���k�7�������'"J��&�Gk n�������1��>�q���=&tlUn ��*�{����5r[<)�%�S���(��4ע�۾o<��)X�Q�(C���"�QB�,�z��R�^Z���i.������,��u"���gPV�+��ߢ*��NK!mkX�#q���9���ʘ��J>o�I:S앮�0����)�6G���-������l�"��1��Rl&�`g��f_����j���y ��N��ۓ$�����12�z�\3�$�
̧�|�s����"����5=h <%����HG�X��|���!L��<��5�}�Qd��Vچ_���O'�����^(^��}����Zz u};<���	{h����Wp�Tdb�4���ˍԛ=]�����&#�++l��la�D���d�����/����h�����lzP��' �h3&�j��}�x�c��Gk���s`;�MIp'�G�Z��}Kp#?�1^
p�1���\]��ѳ? D��ȧM�S��g����8�A7}�����nr 9�cB_�����v(���e��36ωg��j ;��e]��C�e��4�y��H�$�8��⦾�|����Ԫ�|�NЯ[,m��>��Ia���+ /I���X��Zf������]!&�}3P���b�Ag�M\}�0�*<���f��$0F>�H�Y�
t"�Or�r[�,���%/BUv�|q6@��gM�~F�Z�c� 2>��y�Nɚۦ���a�4����-�hb�%���u�����~���tދ�W$�>��h �������a{��-�����{��̻�&>\y�?�i�$U����մ�_K�_��Ҥ<ɷ�\k� �@N}�	��w���� I`ⵑ�uk1-���������8�)u+��)�\�+������­��|q�#2�S��@GW�����%<�f��a�#r|h:�Eb��K�h�x������&I��e?�ޖ�,%�?T'�~��p}[}��Q���8�'��*yKo-��E}j��'u�ћ���u k��|0�˗�O���#��C�
Yk�phGJ�®��)���/s�]�ǉ�;�ӢVw���-q�v4���!��Ԉƶ&>&�@4���ȉE�zR���r P�-�����F'4lyW��+�
S��/����҅?�_�<}oR�:6S)r�#V�)��?�0�d���%f�J��|�ʊ^�	!ou�W��@�Z�[R�ũ�j$~�\vPZ���>��s@j?��(u���46��Ӫ��HU���i@ ��hk�1_Z0F1��/�8���H`#�N�?��6?���\QӍ�����贋��E�C��~̋à��x"I���놵Z��7y��]\��}�g8(��?�e�]�un�Qi���/�u(�})S���}����s���Ϥ��"c����G�j'��G��Zk�PR������W��ؤ�(��󧇿L���H���a��_+������Z-s��>K	�,�`|�/$4ͰI�G$�|?� iq��T�-է� �\�5	U	S<���܃��h=����Ne��nK1�o^���+zK�l��9ϳ! ���nT�j,����BM�7݃��p�3�h����D�b��?"���
7��b�\"gy�o������ߎ�4�3c��C�(�	�X)���x@��譡��(�Ƴ �%.��?GxȤ���6�T[q�e�	ku�J�O���!���LuV��6�2�4�������ԵT(�W����O,z�6�+7"W���kLxh[�q��)�~r%i��A�p�4����`ZM�q=�c&9�-�A��fJ��Z\ܲ�Kv�՘���F6�D#�6�QJ���@�8��#�ms��W��ٙ�e���~|.�10J�H�U? ��슎���+������J3{zh\���3:��6w�Q��#T�>L/�N�e�Χ�u%�kV�$��Ṣ����l�3=!'VӬ$��Z0P������V@��=�ʇ"�x��+ �K��2o��*��i.��=��+h�dj�£Ykq�.�=�z���<C��K�}f_��A���% U^v�0�L����ض)�~�93�voF�cD#t�}Ӻh�_|/*�����q����H�Ea��4N{�w7,��?%���7�O�h0���t�c֗عF� ����;�@~Q�xfm瑾W=�zHg���?�{M�Ma�1g�m<�{X��|�����3+ȃ2T`r�{(�J���%�,���2��>Ͷ�*e�.�q�j��T��"�
��������MQ��C*^�f1�U@�W6�*���h����*���� ke)!�����BViA���2w��e�(�+tS����9�Gl����'����B竗�-�z.�h4>��`�&x7�'�<]��#5��q���
�ڇx%Ħ&�*��O�-�)Rh7 �c0^�[?F����3vz>} ��,[U3��.��`�P��䄊���E3�6��籪ګw�Zm��#���[�����3[�p^xӒ�D����h�ޗK��
NBdN��G>-���tE���#���E-��VbX�mշ8X��&���l�v
�ݚ�qJWQ��0���^�f*�P����GYdH�O���K����66���^>�=¢zt�ˌ9���Gg%�>�P��(��ER�u��s&;'�1�������ēD}F�\��]��t�(��R����I
6�+����A�FS��_m;Q�7R��K�����V�S�o�Qe�}��pR='O�e�xoX��U.��'�gh.�~��z>[���_�C�8��W/Dqk �e|�����#�~��� �����g���k��r�5�.b�c���u�*=���yh���tm6s��o��:剼i��Q(ԍ�+��!ga�$�������7sF�d�g����Ȩ�O�[�m�<����Q��G-�\�"�o:..@���6�������l�
ǽ�c�#6�G7�!4�Y(Uy��K�֪�+����O���v\i6�&p�/�_Wp��a���������\��*u5�!��U~y[<k\D4�	��g�J�~X裞�w��O���W��.��N�?�]I̼���@�2���6�l��G��U��Ś�(`O��u���hj��b�B0rU��8�~BK�,����B�B����[m�~6WX�v7��W���	M���;���z(����lؠ��}AW���Y���գ�,)�( ']�ޑC����2���p%�t��Sw�Kr~x2)u��
��z�<���Y��r�ӑ_a��H�5�7Z��r�;�q���y��4�Zn�/�ާ��\"EigϢ_�C�6��U����E�u��W�4�e�	���B��z=D�#���o�sW���Nx��)�����h�o0�e):�{�(���G�T��q����=�����'x��T�%t�~Jcv!;8[c��	= _�����n;͑k��]�
��=Y1��MEM�J�6����vBl��7D�Y�[w�WKZ�0�Uy7,&�g�>����(����An�;�I�+��#��;�8�U�ߑR�V��y��jĦT��'�7�`���O�� ���@�\P���s�H��/����8