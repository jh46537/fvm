��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�~�������8U�� ��Lll,�3?�c����~#Rl���ю��Ba�ĥ�>Ҽ	��a��v����'��p��`9�?4`��6�&��Y�B�z%�,7��/�J/4�ǑCZ�-�5���z�y���Ɣ�k|Yџ��L��V�C��ґ������H���ϲځ���U�s�����g$��-Y����9Xr����`��+L����a��(�:Q�c�&��,�e'�B'���T�RAu�O��'���<t�7�T�L"�6����0P.V�5F�I�N�i�.��x�c�ًӌ��ߌ�˯��tbW b�
>�i����0�Rk�8v��b"��e�F{��$�qk,�%����'�)�'��Sԑ��u�˕���dV�ǍCa>3���6��C�J�����7 ��3����K\�� �܇AJ�	z��|,ŰS�a�'�C3�ǩ�ŭSuyC�}8��!5�x�3��#�޿�� �،�h�<�*�e����o�"�I��"^Q`���^�m�J��D��BA�0����|���w����~�n9p�V�f%�A6��*�x�i�H����A|�Wuj� ����9ģ���L7S��P���\�E�]��^�s��0�xC`>�����6HƃoO���&U;/8߲�$�b�g�Tr�M&y���a��@�h�ރ��������� f�K8�R� �i��1��������2���	��� ��p�Qt�?�"�Ć�~�����9ޔ�f�/���5��?*��8��T .�B 6Қ$�q�Jm�qd.��5z�|���kIݜ���oFX�7���p���Ϊ����X��ɔ�����WD2L�������'(k{�%�> Ī�z�{o���zI�m�<rQ#0���v25�@�������H�5YW#Xa���4�h�6\��i�־�3ü��~{j��g*��rVM�UrT3F�hςL�eX�jH"o��>>m��dd=��K��|��ע�G�S��8�X��v�>������H.IzUȆ6X��H��TG�d����`Ka���S�N��N�X�p7۽9j���c4SD���Y'mn���/Ɩ�ކ�8`�{��&��\���g0W��P�̤u �q��@�RbF�ym&�|yL���w���+�g.QT:���uoz��y
\��$�?� ��g��~J�i�#ɇF�f`���F�w�b�|��рA�=�t�m��2��"{kA�	Xʹl�k2����d��L�3|��bY�5z2r%�Ɩ�F���q�#�-��u�3,���4��b--z�SO%ĩ����^a8V�TM")+y599�
i��IiK)�̸$����6YFo�%�Zd�*�F�z��TϔL��S],z����S�[�mM�ۤ(םx��j��.dtTbg&�-�0Î�#b�����Za��y���C�QfK;�i�3����z����;��>�u��4�������˦���[Lt� �,�4�2F:�!��k�<�/R<��%�cX�B����is4NЬ]�+����;X
V�sB?���g�ʋm��A�J��/�!�Q��3�0C�ӽ�'��v�	���^c��.u�R/������b6+��Dޅ���N��0ao?Sx��H��v5mJɈ�w��-͒sES�ym/vj���&�Ϝb�n�=}�ʻ�F�-¬MTg����@�W~VW�u��Y����}'�3�]P�I,�qI�iߡ�BY������!�=��1�>��ȣa9�sˆ}z�/�_&���H���@]6$���J�Y.R���ѷm�d~��S�^F1bF��:����MV��1��ɳ'�� +���>�����>������Y_��V��о��z��p�g��3% �F?u��JS�畨��ŭڛ
{�fr%Zb�i��o-��9��j�#s$Ds��~61�Gk!(�Q�e���8��������+��M���k%E���B'�t;�2C(�i*Qfc�Jb��?���ǿ(�5�ψ7W�O��5��(b�R�cJ���D���9��=��bX�����aDN�q��f��U[Հ���w�FJ����#,P0\q0"�aߴ⪡�E9�gΕ}ƵP)B3.�(�1� N�siNd�	5�� �~|���	>��b#I�z��9�����ND�_6?����@������!������Y�RK��ѝ���n%2���7O;���:���z
��R��r=]#�ۂ��c�_�J�����D�h�ݦ��t#T�N�3H3^��RJ�mĊj`�#J�\����	�M�K_v�)���h3����G�K�`+�wy��<������{�*�k	��;,��<�瞲4|J�@&�3�i�"B��X��s��	ǎ�R�\�vi76Q���֔xu��o�l�`����OF
-@��T#�ҤZ'-	"������������WW�(���E����Ь�I,��?���}�y(���'t��"��R�/m9EBW�$�&խ�	�~V�LE���R�J©�Y_pT��E aB�k9�p���tEF��A�(/0��L��ii���K*��ߑ�HA��V�.a��d�/�a�(K�ǳNԲ��Ֆj*kJ!�dI���Ň��Qk:�{����3�t��v}��ny��c&�h�#������_��n���g������Di�ڻ�^�e6A������HD�2�_^��bvI%�r�I�'���H{���&��8�_<�n��FIr���;�⑅h�����j��g��Ŀ�;@�����]�A�����]��~:P���Ш)��P������H�>�KB+�~��
��с!!��L��=�� 9휽�ֻ�40KF��F=�>Q�tv����E_]	޹� �:8���˓��
Ӏc^1��a���E����~V�sv�>Z�_��o�����O��/;�e��	{�L�x�h�s��xE�����nS��$6������6Ր�v��@��Rbu� PP ��bc/k�Q/��u��)�C2������h���,�CC�Zo|4CY�X���P��2`|��T6�y����hֲb�-��D} ë��D�͌n�� h��w�@6�<���o�m���W=R;:���c����ʷ'�z�Ӈ��7��M����Թשw��(_����G9X+\���l�~4����~��c�oW%H�=�/�p�lN�Kw���ڈ���{��D~s9W����x>�\�����+ða29�z;ng�I<�$ޱms���0��F�g�N��1`�����)��t��/ '��ϗ�}�'�/�x������ �(x$����\�
�U`�c�Ӷ�a9��� *��/���p /�g^���}D�]����XB5u��7U�a���JF�9t�KMK�TJ��js������E��.*��!�]�^l��sjs"���:���?cӽ��Y��r��Zʪȃ8Vy@�~�q\!�f�L��ҿ㞑 Uf�f��=�	���
���j%�J����F�}�"�5�8���q��'��\�)Ѫ%m�3�B�=@���u�_�7+Aی������y�O8F5rR�v�����}���D�;m�!�+���?<�'�l%��:��˜�e��()�&�����-�9�s[}R�_��>9�f�E��æ�W������5\�<��@�Ѣ�`��U�P�r��#��$������6��,5������<�u�1��!f_��En�/��9�/ �3iu�u�^W#����;�������u7�o�|�%7��Z2L!�/t��4��cYL�&�y��{AOW���9'H���l�yV�7�e�қ�Y ���t�@����f׸���`@ q�m��)Κ30��X8[�3�<U�һ)��[K�h�OZ:����F'�I@����.&n�N��%얉��*�J�|�\/ V�U�A<�͠�e`������BB�*��N���|䔌�L����f��TK{�RwT�t?����j�0�	�Ϧ��ծ�L�,�$푞Dc_�LO��*�<rx�����e<%�K�����q�f���G(5>h�r�~ MC�&J�C��q��K6H��U�����*��Ȕ���� a,�hw��<µ�m?f���`K�{����rI,����M�}DF��VՁj��˽����b���(H�6���+��:
�Y�����enz�_�Lذ։9Q�����_d��cS�딲JX>d�����ZP�{�0CcŞ/<�����w/���z���Cj�B}��_�%� ϨeWň�YY�T|?%�a�(6Ëln���r�xslu2��K�oV*���^��a�1��G$�B�Sk�<������:/� �5'�?<��@��/{�ߪ��F��6��8k��B��IZ)�LC3]/7�B�p$�C&�H����Y-��?6q\b
��H�F���g�!�ʟ�,j+�nFo���7�E������ˀ�V�~�"w��(e����7�o. �
�`K[7�v/Jd�!e�76F�Sen���$eͷq.K� C�e\�7�e������W��I�u�;�X׀�-Ob�.�%�z���n�T}!/�:��mHo�����G9]8� ���/fP҆�-^,P*�ԭz���3G�����a�,��� =.��?�ž���"S�ZxX�W�4�=9!(���w��yAP�W�nс��e������鱟�v�U�h�}C��H�q�rmr"�_����9�i�-h�ԁ#����bM�9pO4E�������0�Ḏd�&��2F���R��i&5��E;~��$|��TIqP�S�M���"��R�Oӷ�W7�F�/}?����S�I���fO����<H�|�j�R��#�ИؠC3������UNP�B��
F��{��	}x�Ŧ"� yK�W�0ԵՆ��V��=/���0������x��=,������7�شȕ��,�� u�mZ]ƫp�1XΦ�K2>Q2��^�@VR��ӂR���5��.����ޏ	�⮪S�aN��F�B,�J[e�X�rd˰0�w����}n���pfqK�vq�z��)4�'0,��0��(�ޅ���!�k,X^BaX��u�@ha���tZS�2�� ��1�4�����D�V��>�g�fQ3�ޏ��b\�<�*�7�a �`+?#��&�l�&d��*j�˄�.dx��I�I�4 �*��ͽ��ǁ�)�Q�Y�qek������q���SZ,A�C	IrÀos������Om�I�hfĄ�ێ����"��׈��W�h�^Hu>�S]h��n����3i{�vYsۑ&xLѐ�qu]��h���y�$���8l��F�2�Jd�]]"��?E�$5m<�߄
̩�]|���CU��߷�6w�iԗ�|�ܾU]aX�"���6z�*�U74�ta&�]m85���;���k�LR+��?�rr�8F��@�G�9�b�]��$�i� �P�������%��t�n�0Z�7������
�̭1>��R��z�g.0�\����q/|��	�c���M§N���g���������򡽂g���~E;[2%��KQ&C��J)��'�P�r4"�,�/����)!�K�ܧ�pE�c�e���t$-\�-Ml2��l��S#�Q���ȲjidY䖌���'������
���[[P��Q���iĺ����}!��m!�>�C��)<�3��옘��V����Po��NS`s�Ǡ*�Aࡾ��0�Lf�΅�v�����Ci��9|`旂!������FK�����;ܓ��I���N��6��ֿE� gLI�n��;[�ݡsÍ�dRr;��.�5Q�jt�ZŸ�UA�!�3F��Ƥ���aIbC�o����q�$����𜇣D�^�=�a�����^�#��7e��_���Z&^��uSq6�n��(�&ag���Yh42f�T �a�~�Ƀ��3�8�sl�Ĳ: 4O�ί�tI�֠�����V�0�������LN^���ׁ�<A��/�s��G���l�8Aاʣ�+3��Rm�\R�'W��&d��k��ʾ�z�ANQ|�֦�@r�k#��g�o�m72Jn�B��^�z�a/����S�����Ot� �C�Gߙi����}�A��mG��ֿ�RMήEӂ)�:C�Vg��5��r��p0ԧ3�
�
}�R�>�.�4h��	B-v�u��!":�bZ�`��t��� �=n��l�Qə���JXC��A�5l﫫 ��\��	$'i45xRġʻ�U���v�9�,�G�13�@@�o����W�Oф����X��T��4B�;<�]sn�+ɑ��ˤha��G	N�v0Rt+_�C�<����4�M<�s�),�/F�qX����_ɝ(0����1������F�!Nf��U����icAc� :��,.D�"�����ߠї���/\����U �\�d�H����Dx�Q��?U�w8�K_�?H�r2/�y��.�w�?��bd��X��;�t�Cx���vj����Ê�Z�%��������o�ɇ*�3f�C	P&?�a�@E�	~��t-U�� 﩯�؀����A��=I`�p�Ɉ�L��ڲ�[8��bF�A �eJN7�͞W3����Y�tb�>���/�&".�ɟlaW@���L���]0إ�.�ã�����\��Ƒ%FL�C�~�A@x6��CǏh����$�ţjI?28�"�K�	ef9��>��3`�j��(���ӭ&���=���m�)��?�0��jr:���n�0q:7ÛGn�L-h����JtE/��E5�`z+u�/:i]�"�"��zreL?w��Fwe�XN���!墡����n���U�<�h<n;R�^R�
�����[
�	��ڊ7������_8B��-��+~{��(Ji�t�Q�{��?��'v�k��Ŧ���z#�I�>'R{^�N]Y{mE6�w~��6	��2��!N��5�T���p�w5��4����ZS�`��L�aZH��a��]�^��5���mU��v扈�G�\I�:3�
�T�B�U�:����z,D4�d�d��1������A��t��HH|��u���?�<a� VZ5�	:4*�\-��:�#�[.�e�9�$9�c�6�=��.��SX�t�ϸ$���2�Do>�@�[���Icn��SXe����|�t[��6��� �{��/�%�r:�O�_��q�4���\�"�Q)����f|��'}㥠��W@d�e�g/v���CI�!�L&�ʠ�ʨ؝҆�䌋����~KfB��ۊ-��2�����US2/.�'������R�df%S9X"~r��S��g��C�ĭ�-��J��~�RC�ؒ�?�d)xo�	ŀ-1^V�e�Hʧ����Y6�3�p��]J�ڽS(r�	y����ۇAr�<=L�	�d�`j��QQ9���?k=l/ù��i}A�m^�iZ�QTW/6�mBV.௯�(��-vy���Fy�z��W�1|+^k�q˽j/�i�b?�`Q��'���d�%�L�_ 6�TJ���O��kc)���a���(���?L]E�"NW�ށ�����/��Q�7�̪OZ3Zv$Ot�B �����)}��?熭O�C�١:T������5�'�q�ȟ�X��}�\�)����|��l����bG*Bb�͎�r�+���9�� ��6�"��f[|��zKz=�(N6;Q3��������Q��RڎE>m��`c�~u�/����g$Aa��b�B�e��Kq�R4{ �)g��Y��
��-Eg�x�E���3l>ޥ��(~8=�덚x��'�*�Bw�,M��O�tS�h(4dײ ��Z��S}��N}���87�`@�hjA������H���-E�݀#����ت{إ����8� ���+nЭ�[��H�V{'��'�Y�w�Fk �Z_mϦ,�x��������v�D@6�16�������O�3]u��Br��D��
@�|��#��,�_��<�w������\jgAY�$�߹f=ZZ�N�������7�u����n�)b$��$�q�~�G�>�.�ˋ3��c�{ǳ�m��3�L�A-�N�֕+��:�Hf3˩�y�7�-F�L?��	�L�2wi[��5��?��� ��W��u�E�r|��i͂؋��
kR,��$fV�AdZW-��^PiS�8N�F��l~7�����M�j(�K�m@Ŀ̯����d,LW�~���=M��D�	H�q	}�4g݊��e��']�x�Ldלd-u!\xƳR�fi�D�RS��땿3='����a.��|He�2��VO=�k����Vrn�)��l��jӃX����ھB�a�V��y������6�V�����H�[���H=�����)���ϓ��,HT�sC2b?����<��A�"���o�{L.1��7�w�vZ+k����Ë,��$�bX7zY�Q�{�e�V�Y�M�I���H	g�`ؘ��K�$���;�8ZYR�r���Jf촴7�nk/9g�F[b�1��Wv��%p{A�Q���(b�� ��q�Ɏ�Y�A4��@�u��
㸪F�L�s1)MGzf�X���C�u�.[)m(�j�Y(�G�\��Ϣ+� c#!�WU,ݐ,�1n��UT�`"����=����}��2���1�0�G�1��(��Q������D=�I'��eQVZLFY���&fb�[܄"5}���� .�%�,�f�U��rEI�8kW���,�!�Dk
K%|
Kj@��!����WY+Z��e��i����&���P���;�J*�G;��\�/g �c�1��� �̬�[�N$��������Y�K�J��\ǀ�� ��)�\Hg��\Ȟf��i0�����׵�b�E�ێ-JaI|S�N��� ��n�Qv�ە�Z�N�V= �ꀖ�,��5m����y�f��q��@`U���z.��f��[E_%�����Fr��(�]0H�u�1l��f�����@nO����#��%��H�������Ev C��8�0��12����;P��l��Z{�f��Θ\=��FV�������y�6{!���f�@"
1��).����;;2�7��H.Y\b`Z�c��L��Pn�l���X��B�k[�i�,�ڋ�<��α�a�ݙ��F��$暪@f�]Kn-��i���kb��<�ϋ��������X�:%pg}!�='�tD���H/�;2�� ��z�Y��G��ݐw��A����m<���e�8Z�}C�?�ieӎR��ZL�d ��u��Z���.=%�D��	�4��x`&��*��+�*�tG�_�;��I[��됩 UP�Z_�f�	�t:*�P���-�0�2�pR�,s��E��i���p�V� ?�be�F˸
fdI�1��w���i�u:i�����
�0���\�F�-�K!_"PZ����C����v#�̨�[����T���m&<.���jco�s��vk�x�������t=�~H�wZvy�Η���bvc�TA�o�ZV�$u��<ZQov�ha�g�2������dd�w9~��d��J�\�ҡ�X�����(����������z�fx�a�����w=S�q�Ч��� �'�vМѦtVn��s)���8t������`���5�����@��B̒9goO��%2��t
z�-8>}�Ƶ�.��(��I��R�O1��'�bsIm ��ʛ��z���l�53�~�i��T�At�-i��̩L��1�mу�����lcx�+�4 ^mC���HO�#8��dY >Rb�Ў��WY h��d j����l�C�8���0�����LV�[�1�!�e�5�R� �~Fœ�5��dDg�l��_+i���k���}���g���l+/�,-j��[�X���Jc˧����L�&�4������`�̋�U)���d���������Z���ަ "-̖��y|Uv�x4�N���P6��I�=�Yl�Zt�T-�-���&��y�Ӑc�����^�B�B� ������,��o���G�0��PZ�p")�.ib��"9��N��D҅�V�e�2���C��K$���M2~�e!p���F����)�����д6�|Ȼc��
c>��s�$H@�?��5�&^v%*1�J�kSgErA�������5PL��yL���3�zl��+��$�w!qō��hB��1��+��,�3)��Cҡ��� 	vf���f�T}��>���i�7����A��6���2H2�Rv�v�Ʋ�??p�~��t��4���}���ӆ�@�d�cY�.�{��!H܍Rvp���w��l��
�≾�O�&�ծ	�]���=�]�Q��b���T��B^�:ĝ ��
��}��hfC>Hʮ��2\��<I�ڐ�f/�-)1D(8F#B�Q昡;�p	YGF}+@�9��'<�e�:(&�� ��?R�O�}q��2m��Bh&6yp��u/U>��42��23�����+�sE�,f��_���#X<�ыΠ�n}Q`
b# ���@O,�S�1�8��n�N�G�x1Zn�K�3����M8����G��>Q>&{v�y��������[��#���+�;�����jiZ���B�O�� Fè�#;G�aŏ�׳v���x�����{U���隨L�s����G���H:f�v�A�6<q0�g�3���4kJE�u(����DJ׻��Nh^<@��N�*" ������ӳ�1�[� ��#&��|�	����s6���?Z�Ϋ��+ �^(>(xCՀ���� ��a��W$��a��:G�(.��L:H��V�X�������'㜗$@�'��;s���f�`c�.e"�����c��`��G������m�ϛ�g�v-�^�到�-��|I�u($.���L֧ZǨ���EfYGVX_�⤉�J�?�M�‧?����z��o�
K���vu:�ͮ^�u������wK��gCR��R�ȕ�M��Dڔ��.�D����UF�c�S�۬���m��!�s�u7�٠Տg�/���7�H����yn��X�n�O��K�D�7.,|��˜��fJ�)/J��=:���,��"@Us����5ؾ��Gc=���R��}�uHvy�yWPIS�g<��W|)�F�H ���#?m���2���*%uh01�M�ۉ�Hwi��j�L��DW�\{9�{ep[�ύ5���ؘ^�'I����J%-`Lz1俩ۣ�ѫ?/���u�s�Ӑl2	�R��e��c���{�T
�?0i�>��5	������ �߼pCC�̦t����i'q ����Uڇ�5�>��SOpk+G��\���6<���|�2{3�Qͪ-�!�lMß��^������P%)UP ���dT.��C�aQ������Y��`S&/�e��+��������(�=�h}��At>�f��-���a�lM�����NI�ڜ8�=�^�W�?g�n�U��l��=)9<4
A�[��*�sI��ј����d�Wڻ_Y?��#���Q���{2���\�L�эz�����`���*���ų�����\�	?&����jˈ�G�m]��	O�M�3�X�M5B؛��i�
H�k��_�x�/��=���Y�&��ػ����l]�z�2U�H��y�ڐ9�v�q���n�q�T�����K���Q��"���DD: d����)�-�>��'{�h"]#t,�h�#�mR�.l��3�ŵ��$#�>O����e���2E�8������q&"G�?�{������e�k�i	$ՕQ#«�7��g<����r����WԂl