��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5���r��"tz�a�N?�@�8��^�j+C�ԃ��9/w�B<������H~�O�>��	� �nb('^lDp�f�Tuɀ`f�u�	�TO��b�
-�o���ˡP�k��C�� �B���۫��V㻐ME�� �����N�JTW������a
��F�c��^�J��ܐb{�?� �tf�!�/KYc��FIWuq^���m�����O�T�1eH��<3s�7g9Ӎ
<���ݠ�u@Ab�YHe;"p������։ES���^l����(N���D��R����W���xW�#�1���q�eX��o��q��w�#�
���q��Y �:b�2Xc0�)R���ɂ�D*189V�W\b4���u|Cp��|;4�����%ՒeOg
�#�JȬW�5�~��W�k��)��-(�~���/V�'�_��W�
<����ۃT|�՜�mmC�	��^�����7�2�йN��sj�5rlml`�=��}V����)�ƌ�� ��Z,±F�TK� y^+��v])�S�H�=+�@�5:��w�tC*/aSk���4�4:��ͩG@�ĵ1'r�#P�Q�YĨ��AViE�?�0i_����D�~�8�,��4�Ό�`<N���0nEkC�O�w1�8��l�6�s�c4`�A�{��Y�QX��"���N/!�����B����1'&`���b�>���1V��9-H.a���H:�*+����k��$��`�_N�$4��j.��@��*;�Ѩ���n:�{��]�\�N4e|p�v{j�{N��nPf��1;
��w�U��쪁��*����3�bf���a���u&|/H�11��&��lBeV0������圜IM�s��Y�q��BǙ�&軰a�̲$�!�5%������EFn�!jttI��Z��y�o?*�Ӓ���
܎�á�rQ��d�]��O�;�����1���y��Խ��0{��_R�=l�Qݲ� LAP��'�G^$o(B���4�S���K��r�7ӎ���-�Υϐr�'����W�k��I0w'��R�Fx�D���|�����*Z�%%͋/σb����cw���^��@��{�uL)�,<7kR#+LKj}�J�B,�J]���fwb�S��~$*_�NE�A�,���;�n��1� œ Xj�X,�gd����{N&i�4��l���"�����ٞ������i#m���+�y�_,��j7���} �)䏌�r�4h)qGx4,�6bG0��y&:ZJ."p$_4��-������ ��A����y�]+X� ����eP�=����?��#�3�es�9�T �r���̇�w^%\��#������J׼�.3c߾�b���b�o��M��zd�a��f>�&�t�[p^���ĕ�3Pc�h�;�ʺ ���L�A)=��V��H��, ��ND|o�i�B���A
@�ՎX�tg����0�_X@�}c�`���1�|��pJא���>V�yS+Q���H�1o)��)O�l��g
�;�;�tp�,�f@�Fh��G���]o�znE�!��KX��n���x}RN0A��b�3���[��n/������M~$2�*B~��]з�j�1^���E�a��9��?��GVb�|��RP�'���܌%���&Y����g�!��zg^?�)Z ;���<��D��Z��lI�'i�R�&�	3���~��=
t!a�ӄ-k�g�O�����&'(�fd�](��)�,����\�8=u�
���"�zu�U�߽��U�&�������ƿ@c]��l��7�o��Z[��A�����;gf���m�9�s,3RN(h��K�? ��2�OH��
d�":�y2 ɐ�!{��-p����pZ�:e"�
�!&��tJt�R��i�a2sV��3�
�A�t9!�!�&ϢT2�Yye�;J���b���n-g4�7���:����s<tl@sM�
Rm����V�0D�|��r��+=Ww�k����%"����*o2 �C/�c�6�e���~�:ȅ�#���Y����UI��k�6����