��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�D�AF�t�/Iq=���z���'5rÃ֤��8��e�I>1�V���*����ۅ!G�a�M�"̐���K��[��Eۢ�TaYI�U���h�@߮/E��r{wu�����+�)u�J,\��d��Q���x��y\%����I�q���5F�mƣ���n��\�e�[��0��A���P)�[���T�8/)�M���W��{�J]\���x����r�|�(H�;��`���~v�f	��?�����n�R���Y$v]Vq��;԰��3��쿒�[�f���� ��tt��M�#"-�k|� >���s"�!�FOQ����~���X���Q��-Op.��w�h-B� �C���S�(�e�?���ku­�Yu��jc��ͺ>���?�({~�2F8���#�H�\J������QR����}����㿡�F0E��еpu�7��ӹa����V�-č��v4�G;~oBmS��Vvc���)TI���_����=���S��8uł[��\�EȢ�s-�4ȟL�o��t��?X�.)�Dd�� �4�Φi~\���3@/�S���^�V2�j#��p7���V��Lzr�����E4�&aU\�n�����&{祃�}6\��3ڰ��H��e�=~4x�e"S�i�Y�b[���ɠ�a���C}��9��fߍ�#	�U!�l�B����$F��y�Lt`G��e�b�2运E�00�B_Xt�D(1�Y��C��]t��ɼ%?5��}�=����J1OU�Å$��2�oN9�(6;6�H���o����4��"NH;N%G���߁ zZ�9o�9+�v�W�:'��N��Hv��_ʪ����S��	��656��ޓ�LB>�ˢ�B@\j�ߏ/�LO�m����W-U2��td�'E��j:���!��2<.��"z7A縖a���叿=�Z��Y�|������Ǹhe�� s��2�;w�?9��q���q6����&}�r�������[#�~����^"��=w�s<�q@�R��S�}���+�p�;���bȓAZ����y	_Aa&�v50s��8Aݩ�7�	�n�
�s�?�9��n�6ꝶ�WV���h���<z��`o�.�i�2ї��U�׫˘1{���?��H�����S�������٤��M�{�]>+�5�Q��{i��M-������d&M�(�MX�����X
��R����#_B�z@7O��06�]|}Љ>��W����3<�U�K���l���ǫ�4��"���2(�g��*gB.v�V�� �L:����!��uWg�-{��`O_�&�fӵV��a����dPK�/a| ���]R*���T�r�?�Ou��w;��q;��!N�l�q�h��t,�LȱK��:��K8���v)�6"V���͜ۼ�xlB�QUn��d~
�l����9k�I�ѽ;��q��`�Pya\Zc���V�c�@�xl�� -�m�Ҡ52�R�fg����o;�/�b.�-S��X����)HK�!=����au
�v���0�8�9/�p�`�&�_q�됂�2�+a�x �Ӣ8��ʹ�n��37D������_	��W�#��j�T�6��9 ���C�F���Q��\�jmt���k3�P/�%�Gf˧��^M��C:��̧���7�9�`%�X�8q|��(/vݤ�Rp�$+Vd�X�4n�����$��w
�FK��Vl+�q ��| �29���#�,��h���<����`1|��S�V $~����쩩:��k��Q G�p
�:br����P��8��9�V���4�����쪐��T�G��i����	�P�qA���Ɣ{�or���s_ˆRXr"�QXe��{�$��PV��M*�d92�����ɷ���
�s�̀��]x�l�ȴ�oM�j�j޽��9���X���r��T��4�.S󐢎Y���n�zs�D{Y>T��ϝ�xq��R!�@!���o#	���ۻ���kJPz�Z }C)���8.���~��fu�ς��A��M1V�	�Ǐ�7R�T���CAN�_QQp�}���a��J�A,~a��YVN��� ����  �(�2��F��:Ɵ]-ǽ�����0�Ñ�iQ�T�_/t�_6: ^�͠X�zZ� �����0����w�K�����}�2�DH�D����Q�I��9����'�`�R�e�s����1�Z���W�w8,-�|.&�Z���+?m��P.ڢ��I��r����D!9~��ݚ�a�t�)��eu�kXp����s�B�'M��ߨ�==� �o��"N�;6s���6T=�U#`�����*�u���Y�t��ε��[�	�0��i	f����b��5��_]�*�ן�F����Q��LpM'�)����-^3?���x	$��۝��"g�hϏJ��	�9�I�%�ґž�,a�I�y7�2� ��P�x�
0��p�4!�����z<";Ev�^�� '?� e?u|���ֲ�Ύ���_"  O�
pU��e@�s7�����~*5�R�
F72*d�O
bП�\KX1��w)�iø'zo��I�������V$c�ٳ΃�P�Y��y�C�&�epzߑ�>��X*�N`�h	s��L�l��!F[��N�;����h\2m�#� ��d��5R�JM�Q�z�ǭa���]3�YJ��+P�ߍ�H��6��|��&���uR Wh����bb��_9��c���y����a�8�����'�T��6lbV�g��x���-��$[���$Q�`])�\��Z�ݕR�^Tb�WP��*0w@!3*����Z�a�5f|�8��i+�6�mW%�F~?��@w_q�Yf���j��D����b���OϾ	��"�H>Fܣ�:¸8�g��i�suJo�(.#)Ƹ���ƩF�O=�-�C��Җ9B_i,fFD?�[n���F��17���R�L�Q5���h��j�t+�?ν��~��R��Q�-݅D<�d�`�9���Hֶ�]X��t�`F#Ee�(�`��9^���c�Frd"(8�����?��r����B���[T:����(��	C���)��Q<� 7�����o{���}��O
�T����MY �|cL�Q􃙛�Ƨ�𠯀��;�����5>��~��������+�o�|��T�����HC6���� ���Z�pL��K�[��B�v�'y?w87f/*�GB���(�,&���&@d*�T�f�-�����Z���6xv���`4���B1�mV�l*�,q�oq �G�}���0������R,�I�w8�ԦD���.He�[G� ƌ�e�MNƳI��X��$B����8q+@`f���;M�g|�d�#ꒌ�f�QR&|	^����MΈ�T�50�.8��h:��e���[~f��y:|̖ԽDJeG�J	�	c��t�48�=�$� �ҦT!� ���(�6	��ܼ����P)�wߟ+�`ch�nN��bTt��a%�6��x�-=IJ<�_��19�8�Q�솕���E�l~ǁ�)zT�����x4f�|��dD�!�N���]��/�i���Y<��GKǔx�7,^(��EH�!�ٽ_�O�X �M�`,S}#��7�b�7�a�[�+�Ӱ9y�5���P:D�d��YG��Kk��)w�.RY�����=ԃ[+���E����N�[�춅�NҠ��e%��{O��l&�~�/-�8Wv�e���)��.�?���1���	5��N󫝬s9�dKiN�s���s�b �+�A�d��]=��y���/]�i�;��DJ�N/�hB4u�mT���P��b�3��c��Y���>�D��9�����_k�����-�i!����$��אvC���5/.TrT�<V�Bi94M`�=��{���E x�MA[.1F��!��64������to��Xd��2��z�,�T��0~��a�k4�1�G�Or������i��G}Qّʖ��qm�h���"�t`�i��ng绰x����<�J���0�<?8��޷U��/�aC �q|��������Ɲ��޸���S*>1���ܺ�h��J���AV��T<s��R@#��ٵ�4�:��$]n&���Mߢ�~��:\��G��i��F�4�r�O4S�� �}��è���N������ڎ�5�u4h�-��J�p96?�!?=@�7J�&W�j�NN��G͓i��g5@W�H)�3�1��0 6�}(V�A��aT�gMU�	C� K���x?�@�0IdJ�i��i(�?���,���D�(�Ay���Ǟ���u��8n/g���>��Q�`ȩi�\�1��sv�ұ�Z���c�6R�L���D��W➋�T�zF���(,n��x��1^���	�db����SS8�'��}��*�7�v셺@a{��!]玩C���A�E=(ky�$��-��L�g��CHw
��g�gq��8�)n��m^�T���B��r �Tbsԝ��|t����� �b�a�=9����4�c5����8���;��xg�ɮ$��LI��NC��AW%�A�4�<TO�H�xZ��4vn}����n��P܎	���Q�H����_M��EGjcBv�d�-d��N����maX�c*�2�/����I)��jE��w�kߡd^�7v��n���F%?i���R����*���Hx�\�7ig�$��*�����*����q)t��iu��*��k*�W���hmo�#�<������V��^
�U�o��@Πk3�ת�k_�l[8
~�؋@��$}E���S	�&�H���a4!�h\4���Q��E�M��pģ0 :����z�#Uu}�ʗ���M�@�
�5���JVگ�=�ď�S���1��F�_��Q'NGQ��$���%��rw�|��$R����M���HC�ޏV�������D���P���3h�3�_�Q��-?��#�{;��lr�����Ts����d�I �/�E��Wt��(�)�-����ϐ�����7Ґ�7������.��l����@p�lӖah<K�Y����R�����>^�������oV���>�f�Q�?�tw�W#=K�`�U�,(�hlRB����/���l���x����N�I��� �����{�eI.Үy%�-���Vh��~@1,�ǋ�,�Wж�"��c���t��"���{w�*�˰
&Ux-��[��Mp�m%���[�
S�lJ,k8)F/�]��$�g�3E�S��j��E ������G*��I�=tuL��Naܢ.6�)b@;&Q��
�yT�L�^���o_}��V��(k~X#'�B��C��d22�����G��(�J0ݷ?�S�9k�P#w
�݊�6�#���C�v7O��ra����wۺ�Cr��:;���O[Hb�YCgh&qK��5� ���E5�0�	p{]#R��\X�#�e9�hJ��)��ş��Jc�-�"�򇤳?�H��F]oh�k��^���-�㵏���C��;�h��D�����=/��B���@�Ɵ�U\s�ǯj���\|q��g���o�{��gGAڎ���?dpz�>�aJ�:�85|7�.�bm}61����&x,�!EY��A�2�g�g��	-��M�`X6��������t�#w�dw,�_0���௎�q~u0���C����ʌ��W�~���C�fi�}��h�Cԥ|?'ۺi]Wj_��zeo��ؤ�%iZ;K�"��\����A��o�%��ï7tpۿ�RM4b�u��ș2����_���J��ǲ�ب��6�e���Yrx�(�RNpmʅ��-H�k�N���>7�(��@�Kz6@��K
t���;f�\���cN�*z�\y5
DRy�K��*�0՝��r?����Ľц�����QZ�e@./lAޕ|�흖�Ge��֙k��8d������Mϋ�F)Ik���������`��X�n����:u�*�N��e�s�g�WP/��x�,Hj���d���
D;}�`fAL)#8:�
s奮��|:���zC��+�f�U	\~���aC�����P�X��h܄
�&A��?U@X�$����WZ�2�=H�M��F�N���D	��^��gc~�+	$�:f��k�y�/��6�Y�Y��nc����j�*F"��6%��P\��k�9�Z��ӵ�S\i�-�����iM���!��?��E���ד�xP�(�`΍�kԔ�X����ʙM���; �!P���8�3���ݰ���"<�i�
��b?�H���_1L,S�+�⥘���\�'������R�]d�r$U�j���w�6�ӫ+o�呹���U����������3�8X��䧐�MT���S'!�F��iEg0�c�|����E0�Yӫ�
��2����+�Y)���NX5l���*���c7��o(���JW[����
��>�, ;q��ª�ni�&^q�4�xE���@�U񚦾)��MR[i�j漢��6)@)���8��=��|W��?�#�4t�A>�w���J�\�J���c021=R�A�e�ɔɧ�\h` ;0�;��e=��o�Wέ%�]ݥC7�������� �e�	���hC6�6_�&�>�#�݆ �-�(?�B(�4,Y�����b2�T�ڌL-f�D8��#��h����y3�Ŭ�ߨ�QV�|S�������T�C�i�M+�ƾ�^�Hf��`��ꭽnk���o5;�ف�;�9�%u�P�.o:�Y��-<��u#<�|��J�0xv�!̲!4��]Zm�Oq?~w���&�ǡx�!2�fH�:Bgv���?�
h^����0��{r�ņU���iܐ�y��@����1�ƭ�5��F/&�K����_W�N:�+JP�z�'�F1O�$�D��}ZN�9�j��{1�}��k)Ϯi �f�λq' �����o�+s!x�H�`!=B3�=;�z�s�o1�Cj|Ov��_u��k�\Hxoe�~8Wh�c\oA�I�����͆��×�\O���cZ�)2�G�[��W5[
��r%g�q����B,3,�B��*�<6�_�/�p�gL��/$vGO��?JB�uy�~;��R�+�d��`0���-�� /�0���	K�z���J���*7�)EP�,�������/Q�?�Y���%I,ה�В�je�..�&���g�����*�St�Χ����ra��wW}���]��x�D8s44b�}���d���U�+5@���v���A�mr��%���6S�S_Ȑk:.��q'JG��c�w擁z@v�$�D� ۖ���:n� �����u<�L�n�`��ŋ����b�iYȽX.�+�cE�q�2�q��f�ؗ&�t1�%��H��rK�(��s��	@1ya�����]ߨ�}wl���!Jn�?z��BIl�p�d�˕_����Xovx(���#�xFn�DI��Y>,:��D�L�.�/@����:C[������H�ש=��/2$5�-h/`Ɲ�%�!iq������Vsۦ2��_[)\H9#y�ٍ[Jd�� H�9gU'8z5����(b(� �ӭ�@�c�0a��Q+K= ���nU�
�|H��S��݂�8�a�n�s���zR�
���1�� ��@��G����᠌MH��Y��,�3l��M�ՙ���=v]�c��"�b{��L̅�SUn�}�7���k$ӼNo��1X�<&G����3]��ժí8 �FW�k�݈e>��B���KI�;h(T\���p���*����+�kg6<6:��g��.T�M&�0�c��r�8vaY�;!�iډ�rhw�֕��|��`<ݲ�$��K�e;8�%^k��D�O���B��UFP�<(��@�>�>�7�U(�x���9/*�D����JcG|fX=�ƃ"����躔��5�Y���C�en�q����̓5�K�����x5��C8��*-�8�g(W��(�Y-:�щY}KTw:�.YŔ
�>~��/��*���4���Q�s\1�+]��>K�&���>�y�0O�8�kG x�	�Q��O*�J��v#H��-�}�QQ�\��T��ܳ��#�!�Ș�щ�)����PZ=jT�I�8��7;��OG���KL��pb4���)'O'�D��D��֫�����83�Q��H�1-�p�1K��ܬ��U|=��5��i/V=|+c�흊���PN�y�S���i7�>�T\�ʎ��W��Qc�6�5�QAN8:M4+q�ݍ�������P���$i�e���i�ʭ-��-E&&�U�-�_��h܄�y�8ϖ}�Rcp�q���zt-�H��6�r�0)�6��5Ι�[}S͢ؿ<T������o��n�A6[��-���[�>��@!���O~��"w�����4�
�,~Q6#>w�Lc�>���J�3:!�ɢ`A&��)��,[���	��d����@��|����'�$l�t�F�:@'Y����ͺ6��fMW�������ٞ��i�js��:BXk<�}�����ZH(\
�=�_/Gv��
�b�/����a|~&�4g�fi�B�i�&*d- ��寏%�H������8�sӊ�E.��R2�ؒ��7�r��h]_Ye!m2�.�~_���Vq1nDV%v̍�;�m���N�h{�[܅p[�hk��J&RC^�ϳ��L:�C�o�����O�4�5r< K���_����6�97�6��L�ջG�|���A�c(%�$n�S���؏ư��= %�"h����8{"��qj�DZEg^}��ŬW���C���(�nb�[>����h*;�{�Z�a�V/�k�S�b�����T�q� �>��I�
��_4���{�g�����ܵ���N	��� <�ݯ�']��.�D��e�rmVP��,�Aʡ;����Aጇ:�)?g�&c8�I�t��G`Q�7�ne�1��ׅ�Z� �7[��m ��d�r��A���5�T��)5^��nW���G7c����?.2�gn[�>�C4ȱ�q
����.t�-|��iҁ���+�M�[�;F�7Xr6��
��Y=�gzIFM[���^����f&�������")���Mw��m	���z���h95�.���Q��-ñʤ8�DZ�5�%G�,�7����R�V?�߽��z�Q�M4^���I����O�J���B�>����AR��l������f�P�O�Jxa�x�����}h�S��6�j�}����b` �g�����OI�k�<7����;�_�:�n�w��f�7��
�%�dGC.}���k����m�c�]�T��g�6=� ~)<�o���OX�A�F�m5&B)����X�\�-���\����"KޚhHRv�8���]{������O9 	�8A���ٶ�����Z����`
�H7���2���%ˁŽ���
<&�!?ff_.�Fh����d�Ǹ�y��"P��Czy	�(���o��O��y�cV�$S�4Q����$��(ENu���6b9�	�ᮈC�s��L�@O!���Gr��wr�@�
��*��h�����U�Ax�#g�y�~���`�縧2�9\���A�Ay.\N�>?*�$߼[
(+*�>ͳ�yyɘ��]Y�;��(ih�r�k��ޖ���_�gA�A����N~X��曆o��sf�8N�:o�*�K��\�_My	K[�P�dQq�C��Z���Ld9���磬�U���wgWF�C��_���Ē�e�.B�7�`�q%ʇ窨�3��,˗l��K/��lR�ђ��|K�R��g�ZH����WE�	٭���6�c4�?����))E�J��#�+E$I��N�>8KsiO�z{ث�(y���b��qT�����-���n��
��p��Leu��*���n'~j�Z� ��}�*���)�"o�����r͛i�+6�����4�GZ�mQH���0�N5v!�E����j���a��Tʐ�d��E��S�S!B���mx	WI���w���P���k0|����J��r��3�M	-�k"^I�498�2*R�ȝrp��c�$�aRx��6v��R�� ���P*���QKH=���8k=9�=ͷ3�f�tT԰��\W&�mc)9_��zi�V���h�Q�jX8�E����MH����D��ݾ^= �i�#�A�f�AҢ�C��p�ȚF���_v���&��+�z�@\2˦ۇ�GD	�i@W�ʘE/#��'�E1%�ծR��V�M�r5;���⵱��v�$h�C�X^vg(�o�x���b���L������R0{��d���"�0�Oݸ��ꈆ0
�
�uv�+>�~W��,�� ��A*�1�C7��1����@b�
3��~�r��~{���xk�c@&���B>�:�	�.��J�캛L/t�jv	�d_�%p�[� /4üsM��`T���s4�>�#��)Z,պ�5�!�ad�FC�H�� K�Q�U��8tV�2׶�5��+�p�gƊ�X��,�GJ�Ճ��y����K [X�]8[p�� O�_�E�QG�M�PJ��;���7HX����T^��D�+�hp�g ޻=;%��#�D�l�_�#/*�0�{�ίƁ�=p�.��y7*9���ї��=I~B+�ƙ�C���Z���h~
�hi��ҍR�<�#��+�-$yM6���A�CL�쳁F8�/	
�S?Kr����@�ơ���Ij:��*��qש�B2J�$Bxe�- ��YW��@�T�5��?Zt�I�i���j��I�l^֔ĕ����(����s.��V��sֿc�\6{X��<��i����: �t�lӵ'x|)4$x\l`Q�F	V|���`H�LRP\���������J}a���b��1����L�e}G�0Dj�E���w^S8���i��!���T�\OORw�e�
^u׬Zg�RrsL6Wc�<���ۓ	�����4�̝��V����zpq^d���(�����(����C�����-��Z�� �����|�zF,w��0�	i(O�����27|�!�,P�ү=�f�5܀�w�D�D���Y��[������Z&�h����Ǆ�Ђ6���a�̆=�*��=ZU�Zr9��;y{�|{Z�c?��ڗ-�e���߽����gt