��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��e��8_����+K>�e�&WD�v�����d2��~;Е��}d��S��:��|�����x�O�Zʎ�:�u�%$�UKn?��H
�~��qxy+�(G�c�}�8B�!�>�s����1� Pđ%�B�r*�/�g�2��� ��Q���|����h���p� /jO��1Q/�eQQx"�m�7mhѬwu��Y�0ѓ�I��U{m�OѺ`�����|l<^iu(#�z�_�Zl"R5jw�B���/p�؀�h�T6l�.����L���s��[����;&#~etEA�ES�US�^���;X�g�`c�/�������i���j ���I��5�<���z8;��ĺ'�/_Z�D�,�)��J��#� {�rP7@���ZxѤ�L^�Φ������� :�+�WS�ut(-�>2r~�`W��[$�%�غ������4Nq���F�x���Ox�
Mo�%3�΅&)Cx[n#SZ����!�C�p%�<Cp�o>���(��j��j��io8�~g�$�����I�F�N*�VF0�=��C���#�{k��IP߰�#	���<;����� z��~�J��Zf�_t^Fޤ`�`�q@bOsiH��V��?��xE�Dg3��O��f�e�4�!��L���2��G�6��h�P"�Q�Y�ԑ[� �f�QԺ3�[B�q5ݡ��Ǣ��ݜ�G~�#�Jo&x��
nP��� ,aIO���ڨ �\���M�S��i�T�C�?��P���)D�&[�]|�/��Nlz��}���f?@ax����ʈvX���P�^�#j�JsMPyv^�v��r�˓=��3�^>�ئ�*4mq?�>��V�2Ge�m�f�=~��R0Ke�XHp�zb9���3-M�&äG��1���/� �n&�,��������$FD����x��μvk�pq�Ժ��4{SB��8������
k���L�Pi0zm����l�g+�v�Ǉ��w�;�ƺUc�U"E%	�@�v@<5�)���`ES��8j�ƅc2!*�Ű�&B]��'�d�7a.t�Fn�ɭ<�5y��'n,�`������)1���u�ůt��F�1\�+G��{ُ�CKW�ه�a�jɇ�����
Cc>�D�>�8�O�U�BN�����q�[����*=���׭.3�1�W�w>u�;4�M����]7R^D��q<`����4n՚���^#5v�	M���fW��p`b��8.عE'��e��U��
������۸���Z|�R�Q��вK�.D#����)�/��bw�7�c��O.O���� \���bѼA��X�~�������;�j$U�4?�6r��Կf�-��t�:bw���SV�X,��k}�o1oA8%i�f���Y�k�T��LU+yEӡ&���*xC5��U�T9�LpH]��=m�|����߳��]i��ݱ������EyO�V���n�%��y�r����f���0k�ŭ����G�����}���x���Q���2҈R�Z���Kԭ0�ԞZ�9l�8���x#�����2F#��b�#}�SkI��þ����d�,"F�=��*,�:2�?�I�-�{ɢj�uo*%�����kf��6X��!
?C�� ب9�5&?%f1��1���VĮ^?/���V�ك������-�7d���:Jj�G��|���0Y�Y���a��J�@�g��J�\!O:�C7�ѱE�����[Z�=<O0�ZY̈́u��)⚎(4����6ϭN��~��mqw����q]]�$��c����mb4o�_7�fiyi�ͺmG�Y�-�l^1}��i��D]�������N��̞K;�תTvIw�Y�#=t<�ʈ�	,h�lTסAv� ��w���hz��m��G���RxQ��H��,N�5Ҽ�Yap�������f�X�Kl�W�=.�zqubF�l$�ʣ��8Qg��Y���a�Cʶ���m�෮a�3�#~��BRJ�4�
��Ȫ�vQn��C��>�/���\^�Zn�����C׺��T���4~��8�l3�_����5�():�;�E�0k���-�oA~������Dɚ���	����A��ԭF�^��{��c�9[/,}~@m�^�_�߁�e���y*�`?G��5�s=��9n	�i��`��5S�+�G{���@��5���l�K�}<�H���#:e?\ߖTMմ�.��"3C�]o�(���f�׶�0ݘ��O,��Q�	�)Юa!8�a���sLW���8e�ȭ�R7��g���V<m��E���s��q�y����j ��4�f�[�9}y~��ش���=�`�~����1_�|Zf��v ���v?���A�� �V����vyp#�*����'=pN�l��3J��(�wN��-���mc�!�Y� R_�U�P��?f[ku��FT&ݶ��4*\ܭ��+���Tݴ�W�g���v:�}`کԴ�8 ~�QƅЫ~ h�f��~?[�,�s�,�6���d^ k�;d����{TP�����ғ`��x�A�C�8��7��f�vzU��Mƌm1%8f��Yks�&yZp�<b��X�F�D'�9{L��Ĭ/�FI����\�N!�~��O �S������r��ݘ���dɽ��i�꜓YM|�^�ە�x�q��.���0�ǡ}Q����D�щ9�@K�s��<��3(����cĩGQ�#b�>�:4�i�j>ʏ'���Ezʦ�_�(��)��S�e��Vz�y2>n�zĉ���B��� �a8�g�Aj�*���@���U#���h�?]�)�5(:������a㭦-�5�$��w��I��+��K���:���?aU{J�����N������yX��n�Kz�MX}#'�]!e�{��3*���#�������"'dV�&k�@�4@7މ_�z�����j�o�]GQ_7�ސ��%��Z�c�l5�`ҭ��ǓOL�� [+��l����z'��<��P1&�~	��V�V$�����U@��h; ������ϙA)�M��;���G���f��f%��[�F_~�7�;a�)�+8[Z�X~�|B�3��$�Z;��^!�摥*�N�.�;��iħ�JߢB�Z�6۾`N�K�����m��Qwk�CŹA��E�"~c�
�EDV�g9���t��ZJ%���'�'w~�&��l�����k�����n1TTQn�}��m���4!b���DMhW⺄f�}�YA�*0�҆�(�eٚʩ���E�ct���}���\��_�E�� �!�&����D׫C'"�L�2)����~����z7?l��K�q5/��?�o|�l�y��J�t@$o3�^5�&J����SNZ��=�v]":s��£��^z�xؠ�9J�̸vJC�r�w�g��Wӑv��6fob.����qq������x��՘��Κ�P#]H���wza�(��H�k�b�lR�rq�^w�Q5e�ڽ]_<���=e�¿)�~���ui ��O��#,P�������w$��3�1V�%w�Ŭ�]�������]���s�͍^�^�Qm,�UsDCv�s[�
��}�G�