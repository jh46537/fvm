��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�^��h�����mb��feE���0�8GI\�VE�|E�T	dݹ._lR<���<ߵ]�uj�x i�%��K_nl����Qo��
�ٍB	&��jƫe����j/A���� ����J�7�K��j�X�D�
��N_�Ū��`�@��=<(dM'<)+���\d��+,��_x��l{���#д���5�p�-�~��N���(1o/��ctj���}�y_�d @?�Dt�PZ:Պ�N%
Y�~�)[�~�&wt%獵�9)�w\S��6��Y��yfӸ�7plj,�}����MM�C/�(�CA���o��7U�]n�l�N�l�P̥�e�枥�&5K"��TR�J��Al��:�8;;tX�q�$��d�EG���b�'�k�ǳx�P�Pf��`L&������0 1����6'��?�}�7/��$� ���0�s�;�:����oK�1f����I~t4ߝ�7���uw��xC�(R+9�r�,圈K�W���������!������ܕ�q�*�{�H�:�"�kj��0��	�D&'�5ˈA�D�T����><�I��~�JP�$��;P����aAH���tS*7T�Q�B����<Y(�vufN�������`�thM�f�� �5X��b��jm�pq�Фⷯ�wA$��o� )��l$H�V2���}F���1�˗�u����q ��BU�2��V.<�k�֟�w��7Kߊ��ؒ�[��b�Z���Z��dTe�[;m��*%j�~��v��(mm�{�3� "4�=dc1Ķ7DZ�`,*Z�Y/c��� T��
�������鄆d=�2x@o�"|�b���Y>nVGOU����0�����g ���_�E�n���W����J[=ŷ8Q�b�qY��X ���S|�bW��-�S�(�ղ�')Zֿ�Z�4Ys(��Q���߷�a�W��RQ���+��D����{	�y�ldR�s�g� 2:<}��Đ B��+��zob�!$�7��<��(y�s�f)�ԁR�Lgw��iSu�w�O���9nh�>�4�#D^�3]��jLߔV��7�m�����15�xh�V��i7Q��������e�GG�G+����7fs���]�hV��@2���8�|T�wu�\�P��_�!�E���8i��_�mV(����O��ۇzYI�������'���t��8�?�"u��+d0��(�*RrعM�a:9H��	�K�5��!����v�tù�f��g17eP���!Wƭ�����	s�E�e�)���z����ֵT�s0���Ĩ�`8�����V�S�@��t:v���l�o=��.�ô�܃���(Y�l�fG�9����U�n8T�����^�,[�.j�p8R���Y�~m7�����b`yj=9��[oY��*�����$��:�K|xM�Y���D`i�Mѭ�#�`�"��@}9|0��ͅ��W��Z���w0�nƚ7��~.�>��yp��j���Q���9hr0�Z�H��Ua����`��6���x���kS]S����a]P����n�fE�����tρ���eo�l�|8t�q`�?��Yt��x��/^�$:��9�m����|�8��+�x��`�����-��,�Ak����Y�(�����{`'�9��p3�M!y�{ZI�K�l����Z�HH�{��.�/�L�Y�V�(���g�[���Y^��HI_�+�h��p�F�m��!V4+��c_u�����u8��Cx�Ju��K*�l�;1��X��C��$�4��-1�y�`Ò�_�Ňv�:	>����k��O�S�|��<�Q*8zs�w} m���3��c����ॎE���]�қ�RW���� 3�=*9�_^a��Б���c�Z-�?5��X�� Z"����FJ�?�P��EA��
D�#kD�r��3�"���Z�\v��#����<�X��,�MP<��h���� 	�0�;�)�_�d��̫�F%���4��-?r>�!���\y�Ž:�P�TK���q��K �\Ph�jX�D� �u�~�ua>Ћ.�R��\2�R�4P�����"��U���	�b�9�O��&�V:G����ic( �R'+����oE�?�	+Z%Ϩ]���dc��ڥ��Z�1�۔�~�
��'��@e�|��[u���ա(�!�9���w�l=�]zTg�7�U'i�.�;Qv4�ΰ'쀃������R(�Q���Ӈ�Ʊ�k`��.���o����K�2s?��f乳���^�|q>ږ���i��¦���mW��z�ˑN`kf`jKwxK�����v4>:s��̞Cɺ�Y���6���r��7�3\�x��-���.Y�T���Y������ �*̤4�]ݲ+�E�,a��]e$.��#?�F������ǋ$A
&�t��1��T<l<�i�//�L4MM���ɇ��y,�<D�़ �B'�s`�s[_�э肻�]����&Cr;K͹�Ċ(�n��@�X��܄�] ��"?�϶خ.�6�z�/4