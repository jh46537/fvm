��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ� g�I��Jw=���c#hN�j(r�y��l��λ8����^�[� .:{��?�'�iVj���+R�pM�sU����*5���A��v�T�V[y�,+FP.p/.�^�R���ƯH{�2R������//̨�DR�����56#��$��3��N�Ԝu�c�FSGd&̤� ӫ2�����ۋ�"sv+;i�p��۳�X�ʀP�$��Q��,�Ր�y|ZPԊ�ʫ��&�FjDQ� ����{4]�
�����f9��w�p��kն���q��wT0�	�[R�ٺO�>rP��gol��h��I�-T�=���3���ɦGZW�4P�p|ө��X������o��:˩ZrA\��
�͑"��0�8��MY�A1�����t.�w��ꃆ�������s���;Ȏ]k�c�AqG��� �}����O8��^ r�͚�cY�S!wa�ָ�ATY����{?-��� �}A)����+����}��:�Gó�#J<a3S�a�y:����AoK�G2�l�IV�|��.=�ڛ�848v>еP�m�E��M��cy��[6��U��C�n�/�$ߖl������1O�H_�����~i��k���NN'X�Y��vٲ��?a��/���)#�G���L���a����"P��g�lU4������ �M����������lu0�WwZ��S��X� =��;�H.��K3�w�#�J���@��H��V`�(6��޵Vy��N[Gq�RY�z�1!3�i�����o���
�T��4�����<0N����^s�}��9 ���i� >�A�}ѳo���rt5j�$��6U3@O��5���S���T��T}�
��	�U����R��n��@�m�Z�ݯ	�?i�h��^�����`/'�fp��V��T���j��d�}��ͯ��I�������|p�S�4�2�ʱLW!�c 2�/wBJ�OA�]g�x�ħ�|�Q�M��iˮm��C����Z��fđ����ݤ�/��q�*;z!rtj}����xp���γ5c�;����yз�&�wpA��m�aj6����G����=�H6[QJNRUii��!N�SO6�2Ŋ���?��m�h1�e(f���^�$!�Lt�M�NW�?�1F6*?)�d�VG-�������.�5��n3�r��OqHc.ec-_�]����()�rkʚ�IV$h���؁D}L+�����S�oܔ��Ź�Xjb�e�w= '���J|��iw
� 0ŔJ��n5B��ik�/���@Hr�ܓSϼ�6J|��~8 ���h�M�H�k�(�`��N�*G
�&�MV��2zR�W�"}�˔����,\1m!��o3
���_rp�š<�|���^���~K�}?	����Nl8����Pn�L�D�|���'��>��^�Uqj��"���5��sd�m���qz�X�{�[l^�6#-��/iŶ���0q�M�rK����5f�|q��y^�$��b{�SzXxF�m�r�#�Us���*�z3Hf"��c�o�]��YcS���$��l���'~��{��1���%�E�'�2����c*)����]RA�,M��3�x��8�OU�g[_�vN04YF����1�u��c	n���߾�C� @�罜�)@r���H �K0���QEc�]���f[���0r?b�mԖ��3ӻ�R�I�_P��cx|����k�h,���ժ��i�����l�V�&����f9[>��圛z.�ߍ��͇[��|͊3|e��<Qh",��yg��ak���@D�̢��X	/�o�G6Y�Ǟ�~��0��$�_�=/�F]� �/R�w��-!��¿��\���ī(�'�A���Z��k;y�сew�ّ��u�W���39eqOB*4�,!H?&1�B��%��0K�=
j��c��/�L�c��᭞}ӻ��X}�U���f0t�I��/����/�"�X=Z��G���Ƕ�[?$*��,_1�	���|�6����(�eV?	���`�[����䓲�'k��{�&�[�)���)1�!Zt`����n��{�1�j��$�珊�VH�Z�tc5�H��"��X���(󳱦�3t�$)G�V��&u�l�z���\�L��b�G��۾�yq�H�[һ�zHN�����ۈ�S$�J4�F�ak��U9lO�H�:� �_�3hx%I/��5���p�q��|UY9~z6�t�M�@�ē�Y�@�AZę�ek{0�Y����dM�ٔ��g<OA���Èp{#����KO_k�&X�pv�RQ�K+�%���˭��R�>Fc|�T�3Sdܛ������{U�`Q�P%{8X-o��$�^j����[9�Z��'�N�GxK;Q�pH$N{�:AK�z�ҋ�#i�����a��
�����{�����Y嘝E�l��i�p��W�0h��obSW!Q���5f��4x/��o�n�Y�����h��`�Qn8��|�ێ?�-D�F���?4S`�u�yz	���vي��$,������P��F�����'���K8�4�����*i[���)�1F��ѓo�Ln#���4n�\óf}*s�jK65r�'֦M���¯oY j��G_ͬ�n�\ؿy2�f����e�E�n���B�S4B��Q.�M�θ8�5/�!�E���Er]D��ֈdOI�8�Q��1�<�M%��un�X
 ��%�I����K��=��
��n��u���q�&����$T�e�2t��쑰�evH�3*�_S$���`Q��;?T����%�'�c�*�a�K�	m��ъ�=��*��G'2�a����N|���b.C��zx��:F����qM>�	
EM���^vTI?z������a���������EN^t���D��J,��Kb4��7�*�
�]�V����L�?K�x�����#��ꪨ`�mK�~w?q\���q����:�؞�X~����!Ol��1�/�:16%S�m+�)��1�Ƙ"_c;!h�fշ�� �s�����Q�,�Z�V�����;Е-���ut��&);@38�/�;�
�C}9>�R���oI����+�[5cD�9�{�N�g����Y��H桤M@�X�K2z����)��BȮ��������Kt|����M8F���h���~�<js�ߌk#m%�n
G��P�#��df�!����=f������;{�r��a4sWpD$�~GR��1��~VH�!�C�tI(y+>��א\�	��Jc�ɢ�8���Z�aG�[�?���W�sᲱ�0���W�V��
����Ni�Y|14i���o����%���.G�H�^�#��������6���m5̒�Aj�/X��Ta=�t���:ZW� �_��SV=w[��������Z~���ֱ������T���i��G0�K,Y>�j�+�!V��[���$�Sr���icR��\? ���� 'q��(������%����j/5�ۑ���$����k�`[l$�&��I��!�I�H��Z����;���5�AG�'�֪��\8��'{�_��lN�7���וl�6�B:����gF-r�vU��h� �R330�]��ֱd���M!g��:a��f��܎��_����rs�D�=�y,~5+#&ȑ� '���<e�w]j�,��E����E��0��d����w���٩��|��U�;s	�ө��f�i+���}�Ԟ�
��`SwX���>5嶄��Va��p����ۼ�Fsd���
��镺�߫[�w�U�3�䪦����>���M�Ex@�*��}��v&�N��c�{.a��VH9��F�>����q!�⭙���T|�0o?�R�sxt�P8��N�h'~9���۸m9�����!"@�$Kl�9�lW��8>j������bZRR���z!K�D]�oz5�-�\�������i����`T �-�5[tFJx�t�S?�]���M71�:��<�nq!�^�z���%HFr�X�-1Vꛭ��d��`8�'bHs����&S ��� <(�V�R�i�4�_r�d{��~��{�pEc~��\rh�ʊ��?1��Ck�z��bR����-����s�cT����z�ݐOISw�p���U'��*E^s
�� �H.�X��.��ۨ�u8�n�{��*�%��H�2.&'P=�kr,�E���c�^�Wc��^���U=2�ٝ��s�B_�t����1���3%�u' /�t���վO�g����@��<6����4|����Sd A=���Nf�NWOB�M�j�=�ط6^��rMD�ʳ#\t����������j�Ox�O�)�y�f&��4�?$���\4'��/�p�\�Nc������W��<�Fa�M�>]�`z��e$�1/U6R���{ ��@sz{�Ү>_�G`�Mj%���խn,� \����w�P\�&���ݑp+N%����Wo8X��ϣ��\Y��)��z��w�옟��la�y�ۉ=r��^oA�1:yM�z�T��Ƽ� �2�n��\�.����?>�
��Pm��~��Q��K<Ku����iВ���h7 m�?U9n4�vO<����^��>v�����ō:��.�(�����r�<�`$Rs	�+;Zz鶑�7�A���ێ)m�z�d��3�x�2�$�Req)�Tg6�c��RQ?�p��)�E����1Ĳ�����L�^��F��I�޻R����N�E��.�w�Iвq�6T��Ǟ����fM�eY5��h����a�Ӡf�@�\�t�<#}w|;C^Z���R�ޗ����7Y���r��\lp��_ր��<�5v@+=v\3�4M�x&���Z��1S]T�@O��ȕI(��=ǂ��:=��0G��^��]���P��Cw�g�-&Cӫh�FU-g�vr�����o���7U݆����a�ɿK)���׈,ВM�Q���A���Q2�+؄�%O}8�=��X��@j?�ﻹ��\Ar�k���锎�*d ԏ��4)����kGs��Rx.�P��J/�3ϲ����ؠ��g>ia�%�މ"H(�T���&Fd����A �r�{�?8�*&��O���A��T�4{m�M�(��n	��o�|ϟ:�g�"��烅 ���j�jG��:]Fl�-9$L��~�DY܎;S�[���l���1��+^(ND�����-�/,gBG�������ZLP�u�ܡ��=��x����Ne��ph��5���+���䪫iJQ�c���ⰵY���;��쨟�-J������ûo���N�� �?���|�.:ē��gj����TB	�NΒ�Էo�{"���qN�+E��۶�f�G�Q����hl'��J�Af��\������g:�_Ry�"�&PɎ0B�<@;��
P�s������X�m���5j����Ì=�
3��U��C�a9>�n�ѫ�լ÷ُ�N�:mP7!n��U����C�3 ƨ�s��x�&�C��'�H��y��^��	�����e�?�s���O�J�O�7f�����l5��R�#��Lރv�yFz�x��N������d�,z��"����/7��L�J�n[�)��n	�����M8�<�`��g��Z��Z������0DK���T��dR'F�F�]9�;<�؝Ar�� �9'�fL]1��2��F�y��N��Ф��,�#Ksj�n�g��ڴ�B����୤�&�7�2��1�q��$�kS����P5d>^�l�G"����Fx�]*xcg*�t�Օ��ǅ������0J�K(G��:/)��#=/5����9��[,b�������u�X��3 c.�sp	�k��}���'2�K43�������C��mC�}.i�S-�nҨXy%,bIOހ����lC��E�_��E������!����I�>�|����/gp͑Sm��"�O-�}H�x^ćn��$�&)w�|_���yl� [e�����rk�ky����,����'�5�}t �m1,�qNm_�WR�;ג:v�v�"L�_9��aSnõ2v�w��T���Y�C�e�&2&�!Z�۽�k_M��D�C�f|����I�\R�@�VӘQ����H�;��T������V��v��S��q���d_�e�6ftiP�*�×��7�n�H���c��	°NY�(��sUZ����d����͓�%2�L�]�7:,Wd=�z��� �<'�Ԗ���W� 7��4�?��E���}@`�~ ���Ū
Qu����o	�mB�e�v��e�u�H5o�Y1���{����p��������1~6����`�'yx��Ԃ��N#�74�p���9�7�B`�L�"�:�@*Μ����B
Ӷ;[�j�|��/�,DS�BW�>����LY<�3�./"�aQ�Tdmo��A+���� F�%�`G����D7����������H�2���{�o�[�a�GG
Shd	�Q�����"���yi�7C� ��J�Ou}���~�������Z����៿�!�%��oDg��,�Ӵp��E�����e�ό���V"�3i�����I@�iе{�gܕ7�}v9ҒhI}n���,$�n4�HV4���#���ۅ��c����Ң�e��9b&�;@�0��.7�?"hI�u�{4�ꪣ��4Lي�z�G�/�DO�_C!�U��{��-������'�Ru?�9m���4�4=iz� ���;���(�i��/{��ye�P�Y̥	Եh'A�<^i�e�2t%�����W Q!����/��>�ޥ�S���|>�D��bҸ��zܠ�R�&��|3��煥�3Ʊ�`"nW�A�O�{�,<C�W2��﹅��+�-�xy�>�hJLﱙ4EC�iy�;�P\L��*���Z�(���B=>%iT~����@��^�W`y�螦����*�8W�pru�}�0�������A��Ԭ�����Q-�ϝl.U5FfU�*u��PRK8V �]�:��dN_�'�ҧtV�S�3��_��FX6�#V����t�d�RI9/���VY)�����z�8�^���l�ׅ���6Rag�E�twA�L�Q���40�}��*��dK�����N�T�RfqR�.�?���<���a�H�>��J�+� ?�3G���Q��b��W���K��>@#D���v��Esب+I���~j�գ���?ӆ�Z�\��i���л�(K�A4�]c����g���hy�"cO[&ˎ�]���o�P��`��*�'�g% ���_�
�`$8G�
�T��V%�<DW8��&�[1��.�ҙ�{��ٹ����T�k���U�X�BF[�m0�����b���YCO�L�I�І���pݗ���m�S���p$?S��y�/�3�L,?m��>hԂrU����P`�����l��RF���T���QM������R��6`M���'������ ���P��a�D��(�\��:j<�j�c��ｰ��Y�^�R!q6c O�i���`ǃ:�_9B	*���	nP��Z�����VQydaۑ_w���=���ȡ�0���~h�ٽ�)�ͫL؂��-�1���c묃��c۰�)�v�1{�*n��+w����w���7�k�Q���F�GRe�?#�$gܵ��mB��cp;ղ�|�y5��M p�U��t��-B��Л�e�f�����I!���УI�s:t�xRh/���/ʣ��1&�s���La�����گ�:���J� �Չ� 'r�>����Z�%���	1�:A��9#֐T��'F�P�����߂���E���6�͋�m��E�COZZUY�g �K.zs����>��k��$�ZU����}����v:�e����Mw�,����Uౚ��e��
~�y�2��κ�߇ЈT�𔗱C$�
��G�o�r�YE��1��މP���xX<�C��=��,ה�&+�V�<�j�����Pfx��l�^1~���9I�]8���F!�K|�3_��]�T�#d�Yi��0�����$�B�[ 8~u"�w0C�v��z{E��Y۠��R����Ä�)�ߡ��C�6Y̯����T���z�*1qWw;�,��U�+,'�kJ7�ӳen�|߾�9l��o��l%�:,+�HjY�>_oA���L������6���_Q�(���T�K����Y�4�#����5��ܧ+;@H�s�bpk��������-�%-�^ 5X�䡊�ܿ�$PxG�y��ra��`�ᢋh���t*B_�����!�cN����Q
�sm�)P<�\�o'��9�Zȿ���g�>��Nr���1*���ԓ>ɿ��,��R�蹄�m���������d���"O�k�ԇ�A�hS�W^6��O�Ɖ�h&̦������A�>)���f@@,�YҒ�c�:�X$����(B¿8�#�K��8K�}6իơWԉ�8ň���Aw]>�A{0r7���3��RF]�h'�N1�֚F������^ <LL���P�E4@�ܘ��%�jx��NQ�,��ܷV�W n:l�Q��:A�_6�<H����r+z�V���~����!`0��tn��f�"��k�[\��z��R���c�����<g��mR�~��3�Y���*um~���OWV�@NN�גJ�'��K�^��j���c �m��%�O�Ƙ�C�`-&,e��qȇ=bًM���u�&q���]��c�m�0q]�\�j]���z�O|��,���U.w�
ԕ_��"�'�u?�L2y�����|ʵ5���0i�<5��u,5�_�β�X��y���x��Y�qN��+��L׷=?�p}�b���8j���\��q(�e�x���p��Y^�L�S�):Ts  NwhI��(��A;f��=--k�d�j��ͪv!*z������{�HzB��zu�mϛ����o���s�,��]Bikw�����iKn���)��D<(λ'�I#��N��+�B��0m�u'l��e�_��M�m7�F��F���:�Wy0:V|='Sp���^��l��1�_�dj�C�h���q46n��D:�Me�kdI/t�2�~�|]xݻ��P�'P2X�r���ړVsQ��/���=X\b�T�<.z�߲'[�U�I_�����<�e�"���G8�nn$9�Ǵ�Ϳ:G�*P�o���0�ԅ���zҴC1&��[E8l�Qڛ��q�	��������]�y�6���@Z���2�V��7y⹧wLU{�k�2b�7��#L�*�+��9�ˎ���oC��Oc�����[�;�u�~{��P�Y���,b��ӥ������8��:8�>��Z�B�f�����c���yA�9;ُ㙋�>8j*����@����0�ֱ��NN�]�/�L<�1wǡ�s��0JO�'��w����֒��������R��QD���ZSc$I�k�TJ�v�]���[<@�_͔,ݫ ^�Ͷqr��!���%�O�[t2!s�S��R�_��pD�Fk����Zj��}�A(s��ox��L��k�U��;w�i�F���6�6Q��h��$��R�.� F��;+]��/����t��S��Fa�VȘ�\����`�u6:��$���s�k�̥��Ej��]��s��00����0���//p��YGѪ�o�$��^&9��#�i��Z� ��q�Z�\*p~�c�X��<�\�C�1e$z��f_���\��D́�4�_�X�x��