��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���_���W=1����o �6!�z�O�]E�ŕf+��З�\�����`9�1�h^��Ј�J�/����kٽ ��h���Z�|烛�?3Ԡ��n��,g�Y?�K\'�Vً��7� �8��>��������vHJQ�= �1"m��4Qe�����>�O���{:JJ���d�y���5Ap�3�,��|2�"�Ed����<��_���2ݸ5h�J9HwY�`V7�"9����"{?�C�g=j���S���2�|2�r�4��Tby(��79{Ψ��j	�6(ea�u$T?��Z���"�9�\hķo7V"�w���(�큦(W���6Ly�<��u1���]��k~�M�~F��0��Fu�+�����%^$Ua���{��l�|GVH~x����o� ���и���C�l��/h6�W"�{����ؓ$��B�K���90�!9�s�׹������z�� 1��O����`�O����{����0{� ��c������*ɼѱU_d�Uppk��hh<쀁�jÈ2��!SA���N\J29=�SU9����+`�����ο��y��w��<}�p�ʨa@�%;z�vߔ�1��Cj�Ŷ\*�=f��R:$�����Ur!��a(���lB�O��oM�'��i��Gs����X����O~�m&|XH��G�q�3�W�(N����@��FPźKb�B���w��Uq`�R�;�\/�Jzo�Z��5Q�u����5�8Q�§ v��v�ݴ'���)Pn���T]G���P�}y�d��lζ&F}���u��ܤ�[*�)�VdCgf�0��yZ���߁���M���0{���C4b�p��0,?/���V�{䣚��T�%�Rw���4��h$BJq���4�-<�s�G�fo���Dd�YM��A="�L.����G
|�x���i�G_c��;�
:&����$J�-|�ѫ;(U�g�X��c3��2�ٞ<HQs÷���@����M���P�+�E"g�9ћ ��ƙ��_���l�QR~[5��W<���x�Z�ҼZ���_�;%Ȩ�j�3"{�n�U�-��� ��P0D�6��/�Iz��r|$�����Y�Q@��z��Y�B�nZm^w����tsE{�W��$�����斥E	���4�z��嵉�&9T�6�ːy�_�q�4�/.�2m,�H�:��N#ӹ�v<���n���'趠�;ZI=Cv�I�F Zd�-�Q�P��~��Fn:u�z-����OG.}�M�-~I�D�?�;ؕ��1���:Z�H�r�MN3a+i�+�8�]��b��0�TW>�f��ł���" �7�^�(nFD��&��]��*�R�Z��#����NRGw�'eh�{e���6�K]P��|e�	{��J�(�����d�^�� {Q�J��ML�&	�����#9* ��>�$�){���2��)J��Ю������b_W_MZ5��H+���·��3U�Ժ7��^k\���0�m��d���9��C�;E=%�mG���U�
�6����~$ٷ�,G�k�{����Cs�GP[Ѓ����$���m����h=�GI�W��j�\b�7��C�?��a��2����|���`���m�*���d�SE:w�w�D��>��wB����9��
Om� UյSA&GN�"*ef�ʳ���/�I��n�A:�q��8��KRb�pU�����T2��(�bѥ���_��O=.���R�	�WD�,
� kF
t�u��6�L��5k1��ݏ�PMR(� �r���+%�Rh��D�th�N�Pd�&'-����ۚw�-����tp���ƨ|�2u��>�8��KBd�i�?$'DD�� wCm]�v	�t��S��9�3Y*s�@̃A)!Mq}��!_gƫ�z ]F:�?�l�H�7�7��뭥�s�^(J�[GA��Hi�?��D��`�o�T���	B19�?�'�q�Oah��������|w��@��K�&��ݲKt�=N��G}��_���pŗ4�H}L���R�WN��<���� ��Fݔ�ʇP�ٽ8[
d-y;2�^�T'l�4�������� �Ř25�����mY���-�ǭ:�j�"��0]�`�z�Xq��;H�����\��,O��V-���S����}I�İ/�&�����M6�A� H�Y�0����5��ՒfcW�H��6�֯�H�#��T��-�mtUe�,�!��"ѹ^��r�W0fv4ݿ~�ٴw��0>[�
`�\�0��ש��d��je�Y>�ӝ�ޒ���Q\e����s��d�L�8�}�}�W|����p���vOG�ݧ�vh�`=�WPvHu0_o`P0oķ�s�Aӗ,0�N�aW_U�Y��D�C��Һp[�S�p��>���ˈ"��(q�m�>�n���M;��ì�.�שU뼛H'\l�B�3.S+��h�|�Cx#��0Rlqb�&�4z򐌒Y��]nP���?�� ����O�M�- $q�Clw�S��0�Å|���x�-,�Z�������3Ǳ�}>љ�"�s�����*Oa�<�Ʀ����Ue�����Q�������H���	�m��qM��X��O��l]#�.t�M͈l���b8���e%���	�jz�xs�7p��B���Rߟ�W�Z�:�+���ygn��28r�.*�d0�M���=���/��oڬ�MW��a4��5��v�C}�l4e��6�6K9풵9b��J��~"(Ԧv��~I�~������)�(���4�+����M{�V� 11�P�g|92���0<�|kh����&d�C���S����9��k8�����K��x����a.�/nq�VʁX��	
W�,:s�4�YZb��vK�Ĩ���2!n[={q2ݟw�X+�\��.�-"���?�>�m�M��@jz�0�p��Vi�_�=FR|;S�[��w�'8amm�D��mmQ8���U�Wsĥ�H$Vl�J�6|�V�[ťz�H��ʋ�A7����d��p��	����]���Ժ-�a�d�ǜ���ƔP:�a��i>�&j,���nZ�RX/��'�s��ȟ	Z�j"3���'�5)��;��,��xl�/�ß
6���"r��p�#6� �(��˃�Ey� �~����UvT�=]`+�W;�~Y>���Ć���~���-��G��E�AI{�G�B� ��@]�^�X
��v�� ����R�f$�Q	�.�% Ynn�wF��b�_��)Y�/�p�A���������3]�7Z,D��y���/[V�,t�g�_���!���������̙D�e��DKݧL�UF���O��]p�(�t�~����[Ϥ�K����)v�X�X��V�S<4&�−}�`����}��'.쾌��k3R���(��|���o�A$���� -w�=��$�� �ɳJ:�8�rȟ�<�I��)}]�2O0�¥�a&@}@i��Cb�j�����^�p7�0Y%^)�91�į���
ss��r�3F�g���ڒ��0]��þ*��N-�� ��+�:��q�#�P���r�e�NB⌳M��V��<W����qe��.�匼��L���}�a٧������������x��[���	���r���
70j���g3���U� XN�R;���RTd�K�x��z�B��/jC��H`)ߑ�n���x�(7<���T�+��T������*2��������GLC�+�T�Ծ���I-�G���e��EUP�����&9(_)�!m�J�vͬ���JA�-��L���xP��k���9�ʹN%=>�--����u14���ФA	t#�I�G�]#�T��j�.33��������xbO@م��b��+R��vX�[�j]������Z����t ,Q˞Ѐ7���T�$S��?����{��[of�C���t)�������������v��#X�`{Ҁ8����g��[|�ū�]x8uHr�)#%�E�L�Y��ѳ�����1�s1X�mf�%bѩ�;�Z�u���Y:��M׻�������5�Y������D����+6뷠�Jo�	c� e
��Kě��AW�Ac{�>����*!�Gt&]l��G�B�������Y�QH?�XW��e�o�Z~�@�[�'�;��r˝9��fH�I�_T����	�@Ӹ򜕗��ɗMoOV��DCnL��S��?�"����cO7��˽�ϱŧ�f����=��Ps|�#�C��U�[I�o�jY��
*�ۘ����?���Eyź�F}�9�j^d�IO�3��Nd�l�`0L����6���1xIq�,�/�^�\��g���rV� ����fT����V���$[��\�/��������N�gǃ#S����8���%���$u�6Xl�\�f�v�6߯b(��9i�ō�r�6���!ԴD�7:Y����%V���+JXGH��ď	��,�,�S�U�M]��P��� �P����ss*�$��;4��ܫ5�x�*s��D���Hj�/��ac�F�Ү)�(q'��?i�m*�F@���XX
�����U(I��L\�r���G��f��^�8Kw�~�s��������K�?��B�����L?�m����.�ev$ƛ��qI,Z�!&~B3QP7?<��s'T�٤�5P�øü'+��ٕh{Ĩ��%z$ML �����H�7��$^��g���3G���� g�4��`݁����k(�~5|�{�N>�z�p6�2���-�ˠg<����g^�K�c}��6���>�G�[�L���LG�Z:�NO�M�ޕ}ngZ��A�xDyC"��ZK+-��^��2�ϾxYF��*�+�O���CI��=���B n-2M��Ē$*ɷ_���]h!a�N�'�\�"��v�2[��x[�C����O�`�/ut�E���F';Z�za�!ӎm�<mS$���;\�4�+��ˀj�[�Y�M����c�#ב��^:��	��'����ΐ�M���R�x����A��QK��c�Hf�&�p�Kr��tPCY���'z��	�o\�;}8n���h��>z`By��4����?5Za�����t�t�/��w#���S
��I��U�"�\]�tKh�*I;]w�I�m�]��r����>$o�����S�K v�jF��:��棬�����yx�����d��ݧb_�8�O�A/�y6 �kSBV�S�a���������.v�T������4�-��
��VUx|k:��U-f�c�]86g(�:�7�>R0u�[?��K��8�x���������R�+�F�m��WA���:x�Zj�b��1O��Z�G��BG�f�"I��"�49%��.�U��J{�T!}��2b��QA����T§�o�&���88҅pkbt�NXw��d���ч%;�� 
M\ݚ�1�
�6jkL2��n�G7^f���y�h�
Y$����Q�s!ewKGn:�=-�%��t̄]��6�&����y�\ �T$)i��q��s2���gh,�Ǽ��-Gjx�}����/�6��r�A��1J���'�v���l �A�HWf!��$����c�V��ж�ԟ���%8�.����۱��@U��Z.��:I;��}��İ�Z��]:a9(������Q�zr���cz���=i=�nXL��,�|k3_������t�I{N�n)���R���$����O��.���&���#��7�=��կ��S�cL3�œ�Ru���^"�ע	�m�U����W�^�f��G���1����e�`-ւR�+�A��Ee1�0�r��6��B�{�K��/�[�ï\��/���?��0�o��$�O�o3�XXa��u�fd��Ez��E5+��-�._��y�q��O��)c��$@���Ȅ%�J����b��V��+�}xMxJ���& $=�_t9M#���R�'@�G|l��2�-���ac*��=��ayX�_��	��vPX{��u��eg�n���v
�O�9����9V��A1U�D�1A={g�I�t�"�=/��UJV�0�e!���Q��+,Z��B��b�>��=W8�8-5���4|����a�.�)1�t{�B�?�=m�L�%˒H�!�fvZ� .����xn?����J�I��B��d���s􉇴�G !��O�Y�ICj��k��(1!r��7�6x�m�@���Sw����v���
ԣ�ӗK�~���F�MfN��6������
�Y.{��S��Fr�=_��2O�>� ��P�z���{�3Dc(-P/kh�c�G����Q��fFka`q���4 7E�2����!(]x����P1�i�i�Ӂ�?f@p�
�/�-
�]3� j~��RP(2%��	&�} &x����wE�!��	�3�S74��B=y�ծf�L�>-�\����u�8t�^���MAm�HIS��᭄C�p�K܍x��Z�����g��QaB��D�f�FX���j�V�=�d:���?r^��iӏ�F9�
wA�22�ߺ��?���|�0irJf�F�<��㺧��X%�h�3Q�0�I"�x�Ǳ]�j�Kr�̙bKW�6�%y���*K�M�`O:O���m�P�do�٠�^;c�~�la���%���,�ap����;�2rL���M�ye(��h��<����ר�E�TޤzKN�x3/o8�m����MQ꛳�K<\vl�i�(=X�k�G���.��C�(}�HK?���)�������.�;J��f4�R�PeV|�6�/�4!�����[-��Ma��b��d�߳=���j>�����Pf��ve_�{���x����+���y1��R���}Mj97�̐n��I�2�{��H��ent`Yǐ���تa��[f8�g�н��="/	pwv����L���U�z�}r���$�ue�rI�q�̓��:$:�M2�nw9���4�^��v9[�UzK���/޽�o'ރ��I�~C��5�=��n���l�@1����G������{�;�{�s,��	H0����+fR�f}"�d7�"��ti2�h��@���VĈ���{���e�Є#�"6��0��7�u*��Y�����p��V�N��׿;h�@��g��~�̎����C�@��ɲ ϲu`�)��PT���n���I��Ȅc�N�o�Ty���+���Cq�lc�[�V7d[Ou>R��/~�UGgV�<�ĥq�X<�bK�ӽ��j2(�F`���2�?�,�L��vm�H�'��ʯ�ًxj���'xrn�������`���i�� �>��H�V�$G�}$>{�N����<��0]��1��H�D��p.�x�^�1�<d�f��Q(A7���O�q)n�D.Ags[��92
k�4N��57��#�k�����y����2�P�6)&ڌ�<�B��r3���`;-^v/����w��@
���h�ѓt� �B���1}D9/2$�w3�vIU8mYW�F�8�F��ʗZ7��n�M1�d1�r���h��ke���O�D }�[	���;<[ӛS �[��$�Xa�]��H��/�T�p"��� ّ/-�^s"9������|�Ā�X�S�K;��KA���n��D��A����f3%ll�Q�G���2.�G-�)q�BY7s0�f}����7B6笏J��s)��cI����߯�хsc��rv��݌7l��(���	^nc���QW��nU��	��'�}�;�a���͈PɵW��TC��|zb��I��<b!��j�l������4D��d��0�J���ֹRZN�'��!�vM?�0ʸ���o���8�8����ނ{��jt	��2����~b�����O�� ڟ}[�<I�������A,y ����uƽ�(I���j�j����b��܁���έIo���9��H�sŇmT]م2�2��ZF�}l�1�ڕ����������f�|-�K��֞������N{A�
�[�M��>g�`p8�]`<�B�N)��=��Fl�jZ;�לR���ƈE�D�%�� ��:a�^�0���oxI�*�,��.Sl���E�+>|������A9o���&]������q�M��K�����,���`2^�uXo��\�t�oM^CmMj=<�x|�.���%��7U��;U�@U�%^e?}�iŘx���D����Dg�d�SPsw`��&�pа�5[�\8�}���̵��O�:�F�}k��4��Ӈ6cT�C�9�v̂��v,i-�;�K���q�(���H��h��G�f��e������R*X5O	�c��tP$|)��\w��dc
o.�c*���R���x[����Ͻ���j_�.�,?;#��Df#�_�*�, c���`�Q��T�yI���n鍓9��6��G/�к^t̽��-��)'�cd'��ǰ����"=�a�dz�%M;�},�4r�\;m~���ٛox}���|"��*��ԧ��k��]�<��?�5dȒN᤾EJ�2�B`m�+j�^�ŵ
��ʻ�1���$��j�y"��xY3�ҝi/?(
��F�Y8�@�#KL�[�.������ӧA���#j�8�tׂ�&��6}V�!�'_��N�'ܙG�|^���������t�h"�=�׿٩Bi ���3U_?߲���Sɉ��������'���M���ߣAǪ7��ו�.A���l6�{]�'\����Ib&�Eৼ)���ZOv��"ُ޲p����+��d&K�x5Ԁ)dr
����?���T]+��\�F"�㏨t�B�V-ys��dLp"]O�P����L��}V�cd�=_u9Sn*�x9��Gx�X�c�,14�=A(��-�� /{\5�]UЀ�~�m����\�n�p�c����'�O�4���B��@�:��{A�Ū	�o]1��p�P9��]E�?����̩m�����3��:6DT����qs�g�ır�]##լ��duVP��jlSԥA��z�sKM0&!UnBz�B�ek�F	��	�d�9WT�;,���*�g�o��
RA�Q�ydx���ܶ8,�N**Ū�4�*��MyT<TN7��l���VFs�Ŋ��b�Py�q�9Y���`�Z���܇X�t���\�j��FA�ԏQ��qbs��kO�#�N4�V1Ĩ����5�n�8�
f��}�p*�;�t[�C�! ����B=�%*�F�����LX�4�hY���6ӎ�)�ftt##K;��y�f�PcDא�_���Xg5nte}8:b���gB��N_CDm��p��nd�X=5~,��[KJd�)�	��E��ۇD� ��i��2΢�`M���8�m����w�s~�]�s`"P
� ��a��n�c��D-�5Αu,���l-��諃����Ii��J8Q��5�q��5a��%�u⹫��
e*��`|�c��kR���jS��t��5k���2��������X��(re��G�j�A�*�~��$	����H��\��\f�6Y7�@�fo��9�̪UR�M�B��)Ca��t��=���$��k�Ȣ���r���dE��(��yx��%wq슈�g	�o�;F}�t�C�"J痓�ѕKpeT��a"�Jb�MN#�i��L�)��[�Nb����A�Qu%)}a[rrnx\����}L����Ph�cМqO��.ʄ3��Zh�;�r�0oa`]�Ҡ�V͌��
��L'��18NRZ(��� _/��S*���t"�q��~"!���E��Tg��ҷ�M���}䓋1�;|z���@������۳��-�����/�-���Lm~`�h7���	��^��?4�M��ЛN]m�Z=�<�R�_ٚL��UO��E/�����G�7�o���x;�4�fTT�'w�P�X���sZ6^%������J�:Pr�� /	z���x\�c�
ֳq�%���[�6��\2(�-��H_�"N�:����ޔM"T��'��g�Cb>
�Rd�/�7��`ו	��Q�����H�5D5ρ`=���Õ+ijQ}��U���[RB�kf���C�gL���@��og2�mb��F6e"�e�y4�UYi�_���񱁹�'5~إ�C����'O�=���J�[�u����<�zb���R2��w������	T�<�	��~*���e@�G��{;	>7��]В�����~ʞ��1p���mx~�`�K�Q�kG?tv�CZ|1���R�δ�d����P�E4H:)��aK��M1�H��m,��(:���1��CrU��&�u��Wp.�!�j%evb+�%̓X�I��-D8�����c%����9�*f7vՕ(g�3����b���2�hi5IUxǸ��>Pq매����'oߧ2F���T��/�ml�	��3�C��N��#9���c>��J�Ф*�������B���D��l�<c_0����؊��{^��$���q��ެ�Q'�0C��|~w`��X���9:fլ~e-]*�΃:�k�M�}��Q\h���8���E�j�	�7�7�aE�hteೂs���yk�D�@��#.��}Y?);���^�B{�A�����`�Zι�ު<�ٲBz޻!μ���"|�k!�e�Ѫ��&��d��PMӊ
��ع�%Q����缵rl��rdi�$8�B�[��T�!։��v�D��`��Q�v��34^4kJ��}��)@��]NaÆJa�!J�JN{,�v��:��}i�M��A�Q�~`�e rD����$����N��A�4�9;��^LbV�,� �����(ѕ�+���z)�!�뇍If��9�C5�JX;��KJy�ɘL��A��ˮ8x{����3�i�޴$AS���9�:�ټ��f$�gZ��]�J�����in�f�ѫW�u�l1u��E)Cc{)�7w��B5�Q�6�Q��r��Kӧ;�p�ğ/QI2�%���8���Pa�{��.ܲҡS*�|z�Ƃ�� �o�JT����B��`}@[āùv�3�DyJ�����{�O^�HPdP��$;��s��>����Ej����u�>�#z������%�ItB-zz����3u����U�Z �
�isM�܀�p)��<֦
�Qڢ]�=VGa�'F�E%p���:�Q���K�z`%;,Ly�/^�.���I��1��D#�8��E@Q���*��(+tc�ޏ�+x?6�_\ON�t�qf���x�~yj�Y#w��3�6~�g�i�L?��;!|���y�A�s�