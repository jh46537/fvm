��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�Y�э+�`��"g�ȓ��{^�*���;{yf3����t	�q�̕�v�(6��h���"n	�>==Ɉ�E�P����J�-">�\T<�\���H�\�*H��4����7�K:3{���C<H���,�6IÜT \섍����ˢ�pH�I+���\f9����F	5v����֡������(Z� OP�\�؊9����|�>@����������k�є��.kl"���Z��S��[<� ���U��cy���8nVD�0Γ��PEf9=2��PCV���?\� ���Y7.��n9��j�@]�#C�y��N�V��w���wX��vj՞�'!߈=�L5���fɻ�x�Үߋ�8�W�D$��0�����dɘ�s�ߣ>�-:,+"��$�q�	8\ٓ|4��|c���`���PjS��w�&�s�4�7��1�a�B/��� ���ox�h"��k��.q�"�D�b`��!�{Q��mݜ�:��<V����� �D::��٭�f���fJ9~7��)�ٱyS���Y:�%��0���o��oޟ��N;�v��������Ē1\	���g� ��{�2��.T��[^�I��,^�PpE��+~Ő{g�I��\v��̰�$ϲU�:M�I}���j��T��0�0��Ty�"��^��ɤaq���Mv��@S/T	o�Xd��� ��_�h7��7Rz�r;�4���O�A�71�Vh���yT�_tx_m��f�w����,m}.Mc1蓲�A
g�:�]�҃�g7�i�`��	څ��[P����?� �i�.7I�U��z�?j
���%�N��R�i�6�LX�kn$��,E�����?_�H���=~<�3	�hy�:U`?�A�5���ߑ7�	�����1� �����>�����P�nN@��q�co��L�j��^ۛ��(\�쀜�D+�FA��C�%�pE߽��@��U�J��'sh�E���/rfr�t�z�� 0z��h����ᷗ��X��nÎJ	���8�H]\��H0��,�D,��SE�f�Ѡ�1f�9,�t��p	o�8�Jc/�UŌ��K�]��8ƒ;B
`���T�6~a!���v��`7g�?T`W���V �;r�k�i["@�q�w�כ����w��iE�!*�1�p���W�/���}a�窶�hʃ�t-h`:xy��WW'?���?��tbGp8-	s!"�8�*�:�x����1@^3�?u .W��'孽�� -����ώ#�˲N��o��3�4�[@'i����aqB}�@,�X魯t���U�0[��9����=2��Fh�{�7x.O������W}Zuc�e1u0޵��@�᧾�!���F]�Ƀ���_����IH��0��,�kd��S'E�on�
�� ��Ji2�5tB���>���f�����n?�������f��,��xK���rqӳ6uE���*��?���e����㩳=v��N
�hj�P��CA]深R�B�*&ǝ�������}~O�!�]�p��-Z1�]Z鳥	�O�u�5>!g\D�);�.�[���o�8��DY�bc�ڱ�����Q�M�Rj$.������$������Tz<�f^��K�@�(0q�ϥL���R������������ܮ�5��}�Pkwu�4��<��ݢ&?�^3��H ���h:���_.69�91L���b�hz�	^�
���@�`\�XM���2 ��dȫ�s�nP�����pO���6~�U�؟��}�'�K��U���͵>"�Gu��p]Ƶ*Y���F����3��(�{u븒2}��N�mfP� �(c�`;	f=H=R�45�e����O��؉<�D��7QmX�Y=a�'��-z��d�3�9t�+�%e���ڽ;{Hy�2��8�2.�&��&]��z_��HN{��:V�Y��Bb��c�h���՘�upBh����ȴڌ���`=5�8J0)�	�MXQ�Ë��_�����!!&�>�\����B�ș���d�uQ�N,t\ ��H����ܟ6 %h���)b�G���S���b�t�?�Vw�ΏI�Q�0�<'��9U��[gv�
�B�ӱ��;����ȅ���h� u�i�J|��QҒ�|��Y����V#Q���@�vC;��M籠��6O!֋�"��K���5��_	a+���B�,эo f���'2���k`�D�f����
}���w���_	�=����!_QVA��C�����&@uX������x-�cA��I,1�����/�E�,Y���g�����wE��]�����קi�i�>�O,���x/��3��D���q�d-ѫAp�:Mo�.��`��?!�`�Vu��2�{���K
����Hvb�9����Đ����~9(�9�X�KMV}H�vxj��h����J܁���O�	t<���>��98X����o��촧տ�e6t�(uI!���Ǯ�$���w���0�Ș�2�u���f�7'�j�Ueĭ�r�c�Ч�T��Ǥ�{~�`��?�$#?]��lm-I����7�7E9�/�n���0�O_�C
���'�z�c=��/Q�e�,�t�LR�C�5]��Ԅ�V��d���o�//&���'_'و ޕ��9�~?��o#����3D��b�����Z���w���d�`�I:�n6o�Q�597o����%m٬�#�!�[p�h���
_EA�j@4
��0M��HX0�/$�������~�_����5e !��unW�����"h[I�'����K�� ��H�����yZV� +X�_PTa�5AH�-2 Q&����bp��5�c���1��+��(�Z2�Ѩ ����]�O�3Td3l/��(\�=����e��AL���#���E�ǜ������(�6Tz�e�����n1&R�
v�m�ʚQ]�o�ނL�aK�"=)��u~���+�.��I�j� ��h���aC՝B�7]��_��'��<o��6�h:I��u�T�CF�:�;�R�E���F���A"�%2p�?��6��=5�+����y�$N �{��יo4[QL�08�Ɗ	s�	G\Z�m��o��qf�NX�������9��j�9����	Z~
�JS�Z��eJ-�%~�b�������7���n�ZC� >��ǟ=A*ϨC��M��$͓���-)a�cn�!�!�O�QI�$����>jר��Q	F�7g	�b�K�I��yx��y[f�!�E���V3Qj3�%�G�QE�5��R��=U ���Y���[�H����SC}�S�J*Z3Ds]��uPPj�����S5oL�_�� H[ I�JnrR�E%�k\;5i�V���Ǩ�;Q{!70N�Х'�v��_	#^�j�?�z��G���ech'����Gl0�T�u7�t�҉p3^��r5�.��Y��=�+��WbF���4�tc~d&��5PT�7�<IB�g=6=�٦aq������2��{3��~��s��J����j<����$
�u\9%�[ �]�g��D|C9i�Wl�s�fQ��R��k�C��R?�rI{��z�t��[��O�M<�����.�74�R&Jd�l} ���F�6:�������v_ݩ��56w%M��CB��r �u,h���}�Uv�"@�P�~N�����d��f�i3���=U1�d:�OJ�������T�Μ��LgR.b�>M]Ž/̛��.��Gnqs��Bxx������뜐�Т���#<�����>?��;�FpeN�y�Zv!��!�O��/ ���ep��,m�\�Ԃ��2(���Zx`*���z��ࣹ^���k�&�,��f���?�p�#��@f$�
�#NψV�Tm��8~�f㤔����nn�Ӹ!FL�Ϣ�o�����I�P���5��u�dFU�f����6ȓ:��K�Y�f�-Q��9�(jpGJ,&j�`��~��@�AFe�	7�r�{� �R��8h����6u�j�Dqw��g�O�G�aqE��;��Cʒ�؁5v�ˎ\��79c7��$�`�X
%"�W�u�"o��X����+��1�k��4��N~�  *;�i�H*e��tg��pa)B��s7�쟒h�{�"2m�+ë��
��n{x@a<m����E�[s�������[D�Y_��Tz֞د}6c�^��Ut��4�k3��?�~���?����\է�
����136�Cq��f�q��2p�7|�������o} ����g�Eb�����m�������C^	��տ��\��T,���gx�`n$��3�4Boɍ��H|V�1���b	�+�k$�kN������t�ѹf\��>1�����I¨��~�4��$�	��~�^OQ}����e�s��"j����6r�"м�6��A�|)�RM�-�Xz;P�e5��