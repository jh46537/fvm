��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B����R����l�JxM%�$$���E`�����o)lh
6[#V&L�.2�%���1��(|6����"o���F�Q�,���-eQZ��m4�`�b(�I���w2�Λn�J�~������%@��~��� `aG<l~�tG&9��!���Щ� �;գc]���6`�AO鞱����r���D_?���0�����a/��3oE�p�:>�]������+��M�Q�'̌�����{	%�92�L�,ԋvm]�"3�F��Lr򱗼ݣ�65�R�?�}5Jj�%0Š������'�P$f~Ad
ң<Be�7Z��4U`oHj��3���܅K@��6��	����u��//���Z��ŉY�3�[37jV葝��;�[�˟h�ą�x-5��aDX�:�/�)���@F��+W�Z42a����G�>�mr��ʢ	k�`�;�p	t֣�>��s޳醐����Br�#n���Á�h�F�##�����޶� ���eʢ@Jn�v���o=�cY�ӿ����i�R
_�۞�u�مT�f�:��7���Ss��V�o��1@�"�@��[UV^8��V(A���Q��ʾ��D��LBZ��g-�i˞�|U���d*������As�Edn�>������@�A��o��2@'��P�V��b�"�~R��	���s-��3N�)�Ζ�P�X.�1��i�{ɹ������3���~1U}��S��J�@����VV�OX���"�.�!�z;D�J �8�C�u�D,�ɟ͵q��rpCJ���,)�>aǗz����	l��A	�����[�7�b���Y#��v�	A|�2M:6aJĿ�u�Gۖ:���|�4p�F�h� Z�� �l;�q9l�t��$g]�
�4��X���'Id-(uLhD�(� #ҋ.L��� ���t5-�f+�շ���IP��l��
{Gx�ϫ\մCU\�n}���@l�����U�QI�a���#Ybܖ��`���1&��)
�]���(4�?1�� rpq ��h,vu��Z���^����L�:"-kY�Pqf��r6�i+n�`�.n�)w<�wi7٢
�e�p��d$~U3;i��HQG:5��G5���}�7n,H���j���8��1d+ws� ��YE�+zA꘣�-Wך34��v�Pe�j��A{�Sj�����(a�4S���/��|���@<~.�i�oE%�2v�ioK����&����r㠾�Ŵp_7�W,��',��[��^�q�����/V�PU�.	Aj��{�95�EVP���y����K�,���\��
`[���r�u�{C6�B�,���6�f�k�~{f�U�;e:�����D�&M���WnP�
(� �6��o�V{��1p}��|Th�g��Yly(���ȵv0["�%ŕt���
O������n�vx��ɉ���f�!|�tn��Fza�)7c5�����g��GD�؟	,CKt�S��������)^[jm�cGx�s&pi��v��M�9��W�tLSN���rj���������hV{C�p4��`��>��&_]��c�:I/�6�v���?d��|�����Hb?�f��hϩ���	R1Kז�q&����jf��)b�t��v�'^��Y;9݉�������;iy����(|6��_tc*�șl����iWކ2����NE�?އ�(~0�!v~�퀩c.f]k�78�o������=���H���~x�֫=|$�>�7�m���L��z/��GO�h�	<*D�|���3uy��ٺ�g�ս��f���q�lu�M���<I�d��#�Wk�~~DHHv��YhK�,�͝}2�ݩ�Q&rB;�kd����~^��J���no�},-s�W�zU�:R�Ps�%��C���L��
k+��[9e�d������E랲#����^&�J�9��ж-]��y6���LJ���!����GPG��|�� w�a����
�Y�$ՊBW���B]�G�뀓��~X�:�ͫJ��5(�������n# ���cG�4?*���H�?����$�_ڄ,�%�ɯ�Hz�Õ�$�ބ�+m����j\-�����k>4n���h:	�O���sE��Q'a���5Y�1T�#�.F��h�'Jm��[TC��-X#M.{���!٠Mp��$곣�a�O�#�G�NX�B,��㕤�0�A�* [oJ*L<���
���j:@��F����&��p�u|	`���wEf��Q��̛-���]�=!�� �/���L����U�y�n[�f8�oS�	�H"+��ĉo�|
�9�u��M�Ͱ6P�����k~P��e�7�}��8�aZ�~ė}��i�^���b�8������H��|p/�;ƷB-w�V�]W�	�i#�p��eau�2؉�����"��1� _W�_B�A	���$MA���	��x�&#��P�ҫ�_���� ��H�Ի��ԣYP�[p�$���
�{�ă���Q���<�2�H,�T��mL�i�`؝D={^�Sq^ఙ�q�Z�#�h%{[�����eU)��S���5I3��l�i��A���Z����w �R��]u�G ]���1Sb����z�����:�6�8��@⹄nV� ^��G�&�������.|}�3hN�\�P,/Ohlt�qL��C,\T�B�c�|`h����^Ԫ�ghO�0����G^ʵ),�$��vw� ����3tS6`	>8X�.!�Q�J���i�N��e�y8P0��k�e�J)q���a��O��5��.y��x�G��*�5$榪6/2�a�}�|-��,9T�?��{�� #�$-�7�M��ˆV�[9�ߟ]���������\��̗%�V6&�=�/�W�J�3c���4�(}<��Y�����	#��b��:x��&��U�8� �:��cQ���*�b�I�U�u����W��u`�k�8'�%��fl���k c*�j�mذ�pfw��!�q�@պղU>����y&?�u�g�I��K��KY�>pp�xv��pS=�����X�'|�A��F���ʱ���˔�P�@qB������]��-��E��=�Ę16	 ����*�O�~�  �?�A��2�/��&� z[�� �V�*-����!���X�9�זT>Ey�&Y8)8��D{�5P��2/�����".E귨�&��Ĉ�P���!A4e ���U9]򧦊v��4��9
c5%�9�hgI��v�I�Iam`��B��X��"Nzg1�|Kw������W�mP���8�Q]�m��j�ɾac��|����[[٩�/�u�-�D*��;����<�ČS�VS��@j=����Eet���>��#�B�����u�ߝ�qʝ�����y $��r��a�`+@�uKs���d�w��
?�"�W�R���U����R0�F>�([�J�}�:�R��2۰��b	r9wW:Y����%_K1��)�: �P؊�b_J����rΆ����㉒��C�>�c�V���ԟ�Nm.���p���g�������Q�U}ؤ��/�ҙ�C��XO���۫���V��H�`���24)1�ضw�U�Á�զP5ym�}�v�l��|go�L�$���(�D-�R ��BϛN�%��g��R�M\*�������I�#���"'����`z���`�����i�����C[���OYRz�j6�-�$�:���q��n��B����ڌT,�t����yC��}�$c�X\�K�=���כ��
�h)�gs8��~�&$��J���E&5��N����]��K��*���ม�Bin�<H�Ǯ��h֧˴|L;��	����~�i�h��n�թj8��h��Xx�1@[��V�'��)��m~�&DA�d��}�����p�
0WC����D�1B1���	��T��P��66��*=e(~@�bP�<�
�t����-��#��J�Է��?��J����N�0��rxl�~���;jVt�k�c��Ro<P��GG݌�D���B��35�!7�昈iN|`��������\���aJ�L%s�{������K�����P+)#��&.l�b���a�z`L�RM�O畡]�x��o�֏(	�m�k(龪�5Y���v���,�?̍�*�~���sYu"<>�Tf�@�@���T�0��h�����#�9�=f��V�����s����t�mSh�Ү�:c/��=��TfVK�mx����W('�WZ�e����
ƺ����O���Zg�R�+0��  ��+;9�Y�q���z%A��7X	�a���&)�j&�l��55������t�����U�s�[��!��� Y|8ѳ���]A�