��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK��N��.��q�tS�LfN��7��y�����U��lz��5�G�Tȅ��&�=���a��W���9n�l29@�Ǯ��|Ŀ�t��4�`�j�MSJ ���`�->FۻƜ���T�	lU���ςrXE�H�tp7���̚����v&l��<3�~��D�6�/��crb��^�^�9DX��.-�\K�b̷?��I���Y�֗��TH]2�{�Ӟ.�ž�ZM1n}�	Q��Ey�����7��T��.�345K����?*)5�+%���jE�(�T��Ū��#��[��V��%\�PZn����b:���$L�<�n��V��P�bQN�AL�I��?(�h�>FH��r�y��oY� �����w�qH�8�Doi}�S?�؎2��X�-�W(�#�Ňk�\?�WL�>9al��� y�D�/����Rԉ�q���G7!2�$���h�,@��k�X����>7,���`S�6�a��\���t[� `\G���
��h���^~JoN�VK��^qw��[�O��;��A�W9��֘�: �,f����2q�5,��<����c-���N�G�(�����&Q7Vseo�����ump).ۦsTI%ك����߶bʰ҂����i�TC�2)!%�Z\]Kԝ���lz�fHƒ�XyØ�u���/ZѴd,�-�����7��Ln`�$*���K�F�v7 /'�`wJ�����<C��Y��I�I�+0@���p��D�V`�� �����K�U6g���`�
�J�2��v��D��ɏ����M3�0�P��[FU?�����%@3E>I@�`��F~�tT�c�w�}��D �%�w�Ӌ=��߉�%X��s�V�K]r;R�~���v}l�r0���!�� 쌎��[�2N�X�|*�D"u'�io��(7{c�\��3�k�_QT���c� Eb��y�����W@�%�:�m��tS��p��n���KH�:�7�>��"� ����{���!ƈJ�T(�uA���s�ި����ޕn��3h����N�9?Xl�2����~�זF�9QOd�"s�J(J\��0opi��Ȭp2M����� ���&̪<+J�+��a]���]�Ғ0��_e��s6iL�%��%rm��+�������*�q�+y\4EN3|[��>�c'N��Mf(?�N�H�~k�&�O:X��5���ъZ��ɣI&v"Yq�i�o��+]&sb /x��i�� �7"��iÜSR��J��p���X��5�;f�??�J;�+��Zv�p][��s�A���j��L��a!�HH������LU��D�D�������*��,>C�6�N&d�{�Jɺx�,`]�>��(�%XCԷ[_h��o�i���ϐ��]��-1��H��Ͼ�v�a� ��:���P�-z����<I�Ug��/b��Z���}��C���^���'j����E�����W�������ս�^!W%�j��>/���X/��a�}�'÷���؆gQ)a؁�䭥���-�+]�6�)6�>ۆda���˃S��l�	���D ��6~�."�y��æض8��X��D&�l���c�n�02KR|��7�/�`�� ����>��x�7a��d<���/�8L=an�5%�;�v
���%�&6L��4<wc�0�2�kܔ����Y���Z�j*����
YP�)�*��^p~f��a��WH���լf��l�m�m̝{� �}F����M�[T[pLs�*���l���N���=�!n-��ę��� &� 1��/Y��.W���/��`2���*��oڝU�:�"R�w�V���<2)w̐V�6��{�m1ZW�^x�� SI�|�M��@�)���kP���VF�yj�  �H��8���=�5Ȯk*��â��Ϟ��f��*���r�'���Md�3�4I1�)0"r�"Mr�!��Q�ͅ&��ӿ~~��G���M�GJ��S�D�v���]Mm��	���r�x�!{	GP���)V���t6�.\���k�n���m�wkhf3v��()�X1Bݩٳ�o��W����ے��qM{�4�I�2$�-�%��I������$�Tf1�+�Q�g��a)��+��y��-a��ō���G��ɇr	խ�&��)?!Qg ZE_�H9��*V\�d�JR.LD�OO���v0)��N����ӭ�u��/,�뮫�H��Y�S!��yq��<9b��8����Nk��� J�3�o���w���:Z�#/+�+�� �HU���réC�w��5�'s��'��Rј{"\PU�S�(�7���նb!u��GM�=c��*!H�<=�ݨDw35�/T`��%m�H�k� ��o�ǫ�0s>�7_jo�pg�"s{��c���J��3_�X�S���Z�� Du����C%ӁR�����U5��X��o� |�Xf����'�#�A���g���M�f����׃�a�պ�-I�V��Əj���R1���P�͏�T��w�A?d�2��4���ʤrƴ����\�*��N�Z��~\���9��"èr2��pkI�����.��I��l���tI������*��ɫx��Z��ɩ����:�؅����0�k �O��@�"�i�"��{�� Mg7����(���@K�Is�ռX�K�:O�$�^-�#�.�,��м����n��l�'��u�y��U]���M�g-C��5W:S
SΧk[s���4}9���[A<ϛ;�RHa(#.�Y^�=Ɲ�����vm=ӣ.�s�n��_W�L$�}�^��R�V�x���[�#���R�L�g���d�)���SI�`�����ga*֌�zW�)+�1�T��9
�g����]j�YF���R��W��dn|>>�{P}�Ч��H�XX�b�[|��J��T��?�|��-|�\}A�
z��̗^�^HZ�V�����_ۋ����`?[=�m ��4l��D@�'0��N�(��Z`ν7�b�ġ!w8bk��(q-���p���^m��<��Ebl�ѹƎ��G�3@uA���(��a��s��kæ١w�D�Y���VN��Ħ&������?Z���'eǲ;�:��4�%ң�6�Ř��N�@�����=|�.~S�F�b�.��3p?�v�L)�=Ι쏔���hF�9��f��������#�x3n:���̕�:^�k�"�x�#U��1�u�+��=]� �~5,���"�S)D���T�ě�1 �z�_��Ґ�B.)K�X�n����/�Ԅv
���y�K�Ux��O��J��,�֯z����wz�D*�3�!l�E�	�A�=	2���ɖє��;h	���k	�P�@١�i��=
�C���e�R�����[��U
�!aH�{�
45ǽz�/��?֢�B@-����52����|�5�������٘'� ��vՄ$1�U�'w�'�o��6sC����f���_̆����{���ʍX$mv\��� F��W��\��6��W)ɒ�`���*����)۽�!�x�@_�/�h�U�UUjh���b���
0s���/} C�^��Z���!�ݲ�Ҥ�H�ۇȾx���q*���h���X�M,�/��V5Ì,�L�^� m[ok�FU��]k�wy��N��О�ڙ�����,E#*'%̀��Z�w&�
�g1�ʺ�����1�8��9�3sK ���q���f�g����`1�+�xm8�3>�s�B�0ѯ���y]�vUۤ�o.K�h�5*���OK�����a4�����#v��Δ�p�C7�4V�
S����w�P%�" �m[�c	oL����2��s���ǥ�F�����2�&��p�>��&ctd�EX���~HFǷ'�)��T��֥�"�� N@�%L�Q�"S��,���gX��ֹ�fB��X5FZ�.����T�L:n�v����U�ɋ��� m����-����-U��� �(ɣ��^F��6m?LTB�GG�*�Q���dcp�΂�b�?BL+̼-�����	������z�����������0��8�<�.�؞���� ����X��R�UT�W��8N�pj6��.F�z0ʨ�~H�FG��������@$�bV�q^��.^�/ܯ�!)m+?�&�8y��d����Yh(��SZ�+� r��!'sy����F�2tj�J�]�[d9���OϏR��
˼D��w��H��H��*�%�t"���uሂy�w���hK��1Wfb}03Z�eGa�
=�`�Ċ���"
}aq7*��8psM�Fn��g�x �2���EX� ����s�P䊍,�YUrl