��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�/�-bڃ0���ܛ�'֎�f�:�I�gt�銡�����hd3U�&{8\��{,�Ei����BF�����)��+�~�KP�H�MD�W;������P�B�tN�fN�ੈg�q`����)!k�1��T�䇎��w^~�.��X���ƊXFX��~nԭ��2}��=PJ� �W�r!o�u�6ۻ��Q�i&�g��BeX{���?��'Rҋ�&e��@�k`E?%��l��K<�2&H�8y�>�_c�ߝ[|k�Lw�19�����?E<��J�%�EClfx�%��ya�����'����dG�e`�����?ʌMN�ޟɤb|a��<J%l��h���c�f�0�6��b���	6n���2cAԿ�w/����f��<~����n��!�n���^���GEX����r�_�M4�=�3٠�ʜ��N���G�g�E�����p�^�lV�>w$<��9BX�y]�a��#z���T#��tN9ٗ����	rd��+�HWm��k����V��4��i6?�E�1"� ے���Kd?w������K#��>�*}�)�ƢC�#�Cn����j/D�m6��ܨ�0�D�<m��;r�C��"m0��4�<�SLB��˄FǄ�hk\�<씥7�~�t�, m����
>�,�)Y>5}qlZ�
*wؓ(�G/7�&���� _\X��_��|=v�Y��嫃 y��s&Hw��ڪ ���6˫{$�%C�Ȉ#��EV�r@��BbX�t��U���3�n��Y��ce���E���J�va�'4���ŚKt�Yp���9+���$��I�]�jCϓ�n_�LC3#�)���oĦ��܀tv�f紃��8���)ܟ����r G��=W��1�&�ٷT]2핹`q���qM\�Y�� �
�q�x`�l�-Z�Mb;Ϸ@�B��D�z�[�1�om�^nU��옚~��P�ҁ�;���=��s���~Gj�l��iz:��z�@�Bny���������|�H{� F��ٴ5Rv�g`\��R�Gq'��J��D�-�8�%*:�z���mxb
�AJ`RH-�wx.�EX��[�@>@�h��B�`�4�(���Ѝ�W�ٮ�UQ�[$9�WL��{�e�kU���D��&v+�!Kw5{�n��z�|L�[nq�DR�;�򆚆�Ł���O~��Q�w��߽��L?��V�k�m�Z�}qw$4^���@�l%�Ҕ㱻�s\6CڡHp�.�i�)��,Kuy�[] �������`�rJs��ɗ�!��?���V<k�e�ӂml�9#�7��$dZ�/�V�ʈ�ox��u�H!rՒ�s�"It��ߵ%�+G�]y����;D�h��OR�9a�e\��/U%^$�	�v��*t��
#kg9{�".��I�x(��0��ذ.B�6� ��[�\�q���N��}�u!6��d�v�]<6T�D�u��V,g9I��|6���Cc|��h�I����^�5�
��Ѩ������=U(�#�����r����F;?����#sYm��4m�%L?i��:��^�QM6y�f�j�u���E����]���^0�����j�_������B�S�[0����#b\=�4#ڂmr��V�k�*ԏ8�ڨ@F�ۚ�܃	��+�����({>h���2�+�v���3����+N�TՃS�z���� ~��s����+�V�X�~���Q�3g	W��K�������%jExU��k"��d�{`�s�OuOg�YzSY`0ɮR&$���UJ��;^9�zc�+M�a��yh�~��A�o�4J,|��T����`�^�esm?�Z����\BVy�u,��"���7'4?�5�,͏�$��<��O��SOb+_�:G-�SN��Qd.�3��5*�e�k��f�
��a)�R���2xS��p6��v��S��ii�C��iq#q�D���.�TȟH�7e-.�"�Ƹ�:��w��8��I��� ,�.�Q1˱�L����q�8]���E���j�I�O_��̙9ͼ��sRBz"Ko 7�6�D��ޡ�����TF�<�'��d�F�[�Vx��>�ψ�kQ�3���PZD��M�e0�?��%`�`~Yt�U��_�DkY�C@�V|ҁ�y���B6l��5��n���-�v�yE���ʵ��P㮂�t��U�M�X�5����J����Q�Y�+WMzߡ�J�R��-=��e7%��X�/��ú���3֢0�� �5�7ԅ�a2�~� ]�;��3Z�b�VN�X���gH$��s��#���[m��2Y:Lr~lŇ��m��q	��"�J��@O�.J��;K��$��bkY�m�9!2f�b��9޲��T>!�tA�HD��DaT�b��E����r|4��g,�%��D���D$Ax16u��n�)�{T>�ݿ?`[g�ڶ�X����eu���o��2ǳ�/����_�� ��e{>*]�'��|�����ij.�A[Q�)�MMw]:�t�q�Ц9��%J&̮�j�7vh=�08�W�^�*��m'�͓�='��j�|�� ډ��j��	��Al�4��P{�_�����^�2��H�MM<��3��`��ו���_!ڏσ�rN�>*�Ú^�Bn��Q!�9\���hoT��,�Sa��Y.�a ����ʐM�E~򦟏o
�a^mL��bGP�����/P$ˈ�ZF�h�l��]h���XO��,#F�o��ӽ�tA&?1�F��u�^�~S,ﵡE��]��Ωu������/�9��Zv�V����~��2o�7*����M}�����������6$�L �n�|��X�Y]�7$�⛰�Fꎟ�mA�?��������w[c�Y��E �*`�ц�K5��<8�-$yv�%�w���P:����$����/{��ڬ�HX��"���392Kz �-��:ww�Y�\�]������G�V�o�tz��.�f��w��|�!�=7.������\aF`&�