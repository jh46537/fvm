��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzG&jI�#�aW������r�2"ݽ'=}WῶO��nRﵓ�pZ5\��?Bkk�n���7W����@T)Ry��?R</q��Ѽ���U�Cӹ3L��K���(,M��W��:�����K��o��9:�ە�У�	�u�H#/��<K�b>�?5m�^b�%  �����};����U8YO0�E���Sl؇:.�Fp�I���a��={��AtS��´[ƨ�T�;�����r#9��Nf�ܢ?��c%c:�#���-:T[{�D�t�!5VRQ��h�]Ge���_A����4�~ߩ��H� )�8\�m�e�D��	TlZ.�D�\�H
S QN{��AL�[�pb}3���(%wT�Z.(�+�a\�x�]u|c�+��!5����*�h���C�/%�̏iZ�����J��|��㈞����NWNA/Y�~u҈צqu�_G�>�T }@Ci�kf�ws�{��T��ٻ�0f��4���y��YrYt��,��y�t&�T�N�	��������c%���X	xH�=I�;�xWX������!��fX�}|��_
ʣ��Ԃx�L�<�Z�C��	o���y�d�԰�°�k���
?��,��^Nqt���ӊ�C�[�h�q�gd;��Y�A [1�_K�+�m;��k�*��=�;E��l�(�#��uc�]2w������:�N�?h��;�=4�.�0�덾�Ƽ��l��m+Riz�by�d� #���<#�/�^���E��J�A�utz��+b
��O���~eS�u]�ŶQݵ�.�5��.�h��~t?Y�x�|=É!븃�O�b����O4��[���V��}�hݷ�F���5�<���r@�v/��2�N�շFEp�O�e�;�����Ń��:���J�Dg�D�Y���(�Ԇ�$novȾ�7Sy+�xt�F�������EVV�Sh���{�R�5/�x{��$~p+X<��v���{��XH��ev6�QB�����X�4��]�}�/x'A�Ƌ�ǻ�+K�o���v��"Ýo�r~7^��m&8t�p�%7��S��������>� _2������L�(.Tn�|X}�����W[4������@|�	���}"���7�������5׬`�TkB/'���6��PxT\�2��;�M�� Yi�(-�=7�L�������b�ѽ���a�#�`��$���J�T�L�P��2�C��0�!|�Յ���,�)m�^�}��:�� _b���W�JftFSj�!q����ґ~H!�����^,$��uH/�hd&z,Lp��� �yb�;�H���m��rX�6�V�K�9+��w	7�����j�W-�;�X��9zvS��s:0� �q����=]m�83#$ �Y����4d���.��ʸ�INŐ1������������	�u�$I
3��L(�k�+����#<z�O�(���@���w��K��ª%I:'{�~�
R�z���0M�[j�k'��,�+Sf�Y&�q�9q�r$�������秇w��+�qpW/h�����Ӛ�K�FPp��aQ�Ć��	I�Y�6d�tU��'-������&�,d��/^J�q�:Y�/����vf�����DP���g�L��J�ةkC%��k�j�kl&Ŀ��+��Xk���x
:F6	������}G�^�W�Y�s��Tmʝ�^9�a���Bv�S��o���k��I X�[������%MJ��.HXpp��YsN!LfP˥ 4c�ζ�A�e�����N 
��!R�O��)��/�����q���&64%��[tJ����+�V�a)�%~��������K|�M��r�����:n��*�4��T(]xU�c~��=9�կ�޳;,�k��Y7g_�@BR]��e��-S���Jۚ���Z������4)W�I*�,BX+�	S�+����J$�/�K�?I�(y3�/�I,&�e��=6������jP!�A��S� ����tN�-��ҁ�%��yFI��bx��|�|����AhJ���>X�	�hw6i}d��"�3&�pZ������T�^������5�d� �Ό��Mϒ���sѧr��0�����������g��Z�e�>��a�B�����E.��5���5채5Z��/Ɖ���0L��{ HS�uD �Z��L�u:�W��G��TՄ]�f�Y������Y��Z}�o���4�O�o��83�+��l�v���J������C(	�z��:�3���l���R��>yчᩎ���ĠO��x������z�{�25��B�LLl/.����R�	��/q��� >�?G�	<`K��Й;�/nUv,]̍{�#~q�/�<��b
L3 T��"	�e�Y}���794��u��1����2�K��e�(��֞/����7�4�X�Ҽ.0��9Ѫ���/�>#;g�����@���c�o��Ұ��I�rC9����� N�ٶ�E4e��qq��t��9�"a�sLd��h\K��vZ��f.:!�YH�nGU�w?f�	�]�쁀���rg,�/��K{�>�����\��t�_yDx�H���+=޲d7桍5��qg�����r'p^�xL|�w����IG��A?�L�:`ۏ�?��}�� D�3m�w��p���p�&d%l�	r����$���VE4�!^
#�:X��gAԋ�m�(����J>;1�8>��q��{ޫҔ�n��+�����J߶g������F�P��`&>Q�(��,����Xx^/o��c�������9��Z�s���>�<�$�V|����cI��p�<�մ�je��ˈ󠚱(����p�����@�v%����V"���Ю��	Wu"��
|pA�&o(ﰡK�.���Sy��&q�9*�@���T�)\��>*���Ɩ&���1��6{�J��%f��rP	�_ڊ`}���a��tv�o�|$�i��X�^�]�t?��,��e6��W!�m��@�!���壈��	� BC����;)�}�B�������2$/���a��d�ծ9ާ�6_�?24�5���<��ǡC�R����G�|_�׃L��l�#�rs��>�ѩf5��n��*���b׊S����!���S?�