��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�;<�T������8�l��s��2.�Sb���V�3*���uTx���U�Y\Hm�2���d�+�(�b�0��~8;�Tf����T�Ec!�,�{�)��%��`��T��UB|�Cyjʹ�x��{x��VӉ��ϋD2P��0�$�k��;ir]�3y�o�mL}q����t�Þ@�Z�f�ǧ����"�v�8L@���N���*@q��+�o����%|v�P�zZ!?����o�s	�����ib��23,�E�FS*2ph/�*�E��۔���iKj�J1��l�����`+A#���/5�ڎ�U��;��E�<�����}2Љ4�*�HN��nr6�?鱧��El�4_�6�WP��/�q�0zO�ꛆ�0w*5P�P3ְ$�!����{�1M���t��9$v�����t�;ם���|�)2��P�U�v��ڱ���� ΰ��"T��<;���.ꁀ�������aGć����#���E�Д^�B�O�v-I��IVq�m�?	߲,��=m���1��PO���Oư��}h�#�@�|l���R�y�yl#��L?������]���wv^��7a��=#��^a���r�����)�>��v�7�7~�W�?�n~�	�3 �S��V1�᡻�����*oC��v��>GV�q��=,,�Y2þ��a���kIe'gŜ�vy�(_�"�� 3C�'�U�.��f�+ЛN��6mL�RU��קc3Ӻy.n:ű]|~F�� �Hpa��X�{�	��5���:�lg8�ȩJ�����V���Po��%��ȗ��z���a���6�Cׂ�z`G�K2�g'/��qA2�Z���U��ܹKA�HV�&�#)�A��"[�-9�����ܤ��j�Xbȯ(��o��@��Sؕh̩�s�k��&��-�m؉i��[5��:m�=I2�tU�Y=�ͯ7���w�*<��>&��[r}Z�g0i���!�#��<T�z:���-��St���p�b���������'�� v,@"]�@~��̚t��fWs��"�7�+����l������n�T�|U�@�7]�
	���`�Pj6%��k籵�ew�ᴔ�< >��8�}�AQ��b�h|e:�`W�/��a��i��m,��uINbM�=�&��<���0rd)���=ޘ��C���
Y�Qgċnr2){��*3�m�=�{��������b��9��N[�>�ao\g�(V����>��FJ�MY���UO'���$�f,J	�L������ݗ<|5�sѓ_Y��]XHA���"i9z�X��Xy2�p���F���]R��h}C�d3x�6$��D�a���#�:��V"~�4��f ���َ��L 6'4�-�F�����
!Wd;?��ދ�Y��䰿�|�z�kj��-�"���+��Dp9[CmG����Q�(^���R�B�H�� �OH�cxab2�%I$��2P� ˜��g�� �*��E:Z�-"�< ��O��J�&�4�U�q��d`��	�B�d@����U�Si�=I�;U�s_�q�;G�����yӥ9(���E5a�[v�@<�@t��~���"��,6~�FmD[\,V�=�����?J��"�����Z}��t�8z���s���	h�@� 8o��ۆv��z��o]/|�Lٌ���d��~:`��	3‹Ξ���h�߷��2-M�Yiq+�Z`m:���?�<�����hcH0���)b9:.+��OG����s�إ�½xj(��gE��v>$dϧ_K7"��|��0�'��ªz �3�y�H��M�/UmN�e��]6/叮�	��~�у[q�B+B^�ǚ�c�(��3����OOl/�^�[(������PNP���\h�4{�l�j�de3�C��7*��χ�X2��.�R�>��E�;��Β��rլx���؞:Ŗ��� ��Is�C|D�S�t��U��}t}#�b��lA8�K��l��]�3�q��%^��3�P(S���-t��"����U� ��̟L��	�pG��6��G�r�V[�m�+��F7�榱�,�n�N�=b�M5�`QB��&������&��pq/9�Ō���6���J=q� q����)p:E;�p���C���}ݦ0��_VV�2��֘�`ۊx�O�3U?ޝ<�ނ�JH,Z�LJ=�\T��L0_Ĩup��x c4-go7��B�>2^K(��9c�3Tq7�/j{EnV��>�q� |���g ���7Kp!��j�����[��Jփ���1N$bvB{3���~E�P�S�}
Th�=��?�#�[�9�,��olO|B��g�xdH4YK��A`I�o�����G,��ى���ӧ�ȡ}�����g�f��d.r�2s�諺� ��/5
�}��Cw]<���f��,��X�%Fp���G�PUu�ᰣ��*���#��ތ�{G� >�� ��Z�n���lإ��D�Fje���:"�[X��U����0+q�>�)�f C��=l�%��m:���ď>3gg$_��8�3ڳz�]�=�R���ЈN���+ţ��e1�0Ww�G��Y9m��7��a��(��M����d��_�Rd����6b�#��d��N2Ol�c��!�ߓ��e+�vn=4�-�Z4BvT��Ӱܩ�. "/��n�J���Bv.I��|�*P��=�łz=ŏ�����=O@�K�A%z)c�c#ȕu���P+����7��6�®1M�I��hx#>X˧8�Z)O��|��Axh#T��hƄ�@|�D�6T���^E�M���>+��F��3�抯���!��f��l	���� a�Rk�Oc�y�o
��;��4X�%���۰����\�ǧ�ܥ`�mМ�V�<�LGN#!�a�l�6�$�3y�����U�N���t�c�K�f2+O��7���!Cv�My} �4I��d ʨ.���2�;U�)1�F���nn���h_ɯl�|:7��x���� �Pz�y���e�Ѕ���]�낁�9�!�~��
w�SZ�*w`�5jk�Rk��wB����U�m�\"Q�`�fad��p���7�7�;2�M�`>�Zl�4��UꚣŸǛ������e�2{����f+3��s��z�e��a��������,XTJ����ә1�D�Q��hԄ9n�������5i�ցV�"�����K2�pt9ݏ��>�/�[z��h8�-�b��g��(���4Q��:��ʚ��]��2鮯�m~�����r
�e�������}� @�Fb�;")1�	�n/*��2��f��~�������?b�r�XF	�O���.�������&Z10�W����W�	��<d���q�U1��]��H�pA�#j翍�Dk|XكN,��g�Ȍ.���~gD|��T9�L���|�Rm&.�]}���s=$�1DzX�t��$����,���E���QN��>[��ŋEЕ�س;`��q��!�����N�G��m�=ؿ\�����,\�B�3T0���1��WQ߳�Y>�A$;U @K	� ;y|jS�ж]�:�z�?<̯�@�V����4��v��gs~�&mʡ�-ߞY*G�Cg��s ������(�:W������
k���ۋ2�t|يsL���t���3����}n1E����j~���r��� ܜ�- ���m!82!)���ϧX�ȁ�2�͜Jl�;��	�%kT,��)�H��'��M�̾K�R���//�D�h=w:�
���T�ʳhpl#��bi� ~LPg�p�c�f�e��,� y�^�,�Z/�8��H�?�f.�R�pN_u��R��V����Zvv>t��.������L,���q)44<�'x���+f�ʦ62�9b!@�KZ �Ȩ���v�+�;��C��^c{'l���(g0I"tk)kդSH�u:���>uAr�W���w*p�.�����Q��h����7������d�j�o�_"g;3d�9�x��V�B���D�@㖛����4�oy��V�c��uh�)X�J�Ġ�k�kگ Xj�
��\@�Ԍd�;�ʖ�V�ڕ��cY���+ߦmI�����ډ�R�o��5�N���}�~ӧ�E/�"\���lk�v�Zl:������0�h��Hm��R|?��d�^�F��}��մ���¨X���(
<b��#��o&fr]'�>��]��G��	P�Nz��Ѓ�=(�@�d|��7\
:U�>tvA/�N��}�>5[�#��%3�H _��fx��?U졕�5UM�h�?Ęky��Bc�X��`1N]%�"K�TNH�&��ŕ�jv%��$�b����̄N
Pl��r��"�A���Y�.afNz����Hb��>:���e`���w�Ą�ϙ��H�K�����7�1<r6I̎��lO;��e��O0p*�p��$�q�H��`Ao�RW���F Ճ.�,�1�$㰽�M�|��q��т�N���8�@)Ha���k=�����G0f�9�l���}m���;�*7\U@�-��c|��&�ŵ�|P��(�\T=��
q@F���|a�b8�����j�]��";�
rqV$.]� t<��/�N�h��[�~��q�]�zQ�y�)��c_.�n�SD�{�!�8��G�D=)=��{�����q�ߢ�]y��*�=�������GV����_�J��%���FH2��-P�A?nm�p$��3��Qj��U�P��>�_��*�i?�@6�H�6	��?���۪�D���ʌ��o����<l��Ƴ��������DF�#an�u۪�_ov�;��p)��[3a�~GJ6]z�^�� d��Z�i�E9ҩ;@�HL�!�E��L1�$I.���<vsm&H%��p���K�&����`��d��QJq.Ly�cz�˰,�V	g��)�G]����KV��Knm;(K�粏��hz0ENy�l@��� ���L$![�v�8��j��E	Y�ዹ{���X8�n�=�Q0؟c�BV"s�;����nP]�6����P��!tԄ��Y���]Kׁ�	�k>v��"
n<J����81�T�dO�ٜ=�O�cEL2��_I����%���{��;e3�!����_�c�98�ϰ�y&�!�V���WHt��w|5�n��x�y����
��8�َ[4��J�����'<�>�����zU˩��<t�}M| Ab�h1q�����m�>���u�H]c�ul% �``U�����T���&`=]}��/g���ԤÍ?WXm����l�t���o��m����~.�D� ��#�0�<�=�:Yk.=j���D�-��*�j�a��A�1��~ӣ6�88�9΅�	�����R�w�{i�l#��9/�H9G�rBIdn�.Uμ�8O�q9+�VtԬ25�H����&*3�t<��k=�!��W���	e�1`��)�]Z��b˲�T��oO��[O�?���d��b'�t5�O�i���Oݓ<��]�X�E���N��y&�pR�߮?�?���-�h�x�,��.ں� �V�ݚ�ɸK���K��Y`&I���4{Uojm>�Q���o�)���ዯG�
���å��M�m�
��L7�
Yک)	�j�G݄�1p3qH��9�lj�����z'}�)���B���^d�Y