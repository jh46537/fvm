��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�ӿ�J����m�`��u&�ԅ�mU]Z�A})�v`,`&?S���.��K�@� V�sĺ��j��Z�+���8��/��X(�K��*3���F$�2��k���ՠoȏ>S(z����ڟk�.as-�jՙv��Za�Xc�<����/w��K�Ƕ=j����[�����H�l���XmՇ�BS�@8�F�3^�X�AW$RV4��x�~~�%�xB��K��k	��=˼�H��mf��.å)�'�t8#��o���(n�Q��
B�9�M���^���d����<$�s��{��S�%+>�995XP��[B�&����mJ�Z��N�� ����T�9:���f�j�u�}-4�M'0�>�۱!� NVm�]2P�r�K�Jaক��E�&��ډJ�S�ƜǑ���-d���y3��H�@�q��������E�
C����]�����ݫsp(��<R�|W����
4ٶq�.w�1 ���_���Լ���}��O N殳��F�����������;���
&	W�����c0��!D�j��dT����@Y;���V���z�a+��lZ���e؏tG9�I�-�g�����sn��d{�)��T�2����w~��b@=��"�nN�z<լ{�*����)W����9I; .(���O�e�	���\A�e�s���Ew�Ö�x��Y.�f�P= n%��5�=�����#��s��ŕ}�����{�}A,���_<�J
5/*�]V��oubfm���x�n�a����"2P[�	~.G��m8%��~�]���X�I���Y����UQL��(�)��7$�����v�R3ò�MrƏ��?$���A^N�]Z����k$̑�vy'>(
xh
�E���&���J�CM�t�>�i�
UNa)�ݥ���D�*n�&r�����T�M���)!��V��ZXH`XhK�x�o�0�ւ�	���U� >P�@��)��z�%16�u7�������=�A
,|���#����2���?g���^�ֆ��� �{�s)8/�R�����7��.���-D��v���.��������=�T�?٨߁;u6��q��s�r%<\k4P,��i��Q�PDU>Y��<�z��Tss���y�Vp�����}����Kk���W��ԏ��ì�0��i��̀ξ׊¼�H��6����?�E�(r����n3+��^P	�LU.�p�C�z��K4Y�i�>π������ڊ*�N;.쓔�z7�7U���ᆫ4��ҡ!5�@�1�9P�6vFc��mwyD"� ���?pa<��j�Q�	�_�ֆZ�P�VYdF,o;���(�[Q/y���!�^��đ�|���笟�5�P��`Zj���?T4��q��Q��u����]�>���g��1������E*�/���`$��q�5�C>?R0����艼4
���yX$�31^$�k3��~�9!Z��gXYr�<���$�,�0h�Q�6�D��l�J �C��fo�ï�f��v���Oc82h��w}S�����0Y?�ْ�"���a��J��YTޣ��z ���]'g�{+~��$��17�`���^YT��߅h��I���j��.��&�K��j%���C~bw�T�U�P#,~�9�FYbz�A�d	dA֖5xI�}F������M`�̬�/ا��ή͑x�l[�N
�7�ic��AzXa(�e@ؘ=����
�����]k4e���?~�loS�kʛW��*����5�OD�;��8`v��,�W�	N�Zț#��߀E�R��.("���u���OeU&�����q�|����0t"��C���W����`H�0U�N��B���1�W� ?=�u�C^>�)B�SP+2
n��KShQl��-���R-�c�ߩ>�=3�"*��f+m�ᤎ��k�]l9u�>�p�S,b��֜j�l9��|�h]r�#%g�Vt��Q-J�4�~B�z��m�5|��܆�4#�O���K�(S��<ǐs%X&ɉ�i5�؈���dHv��<����|�TJƆC-^Rm��z����E63����6�!y�
�K�! 7�����2j��s��0��7����ӯ-�����Y�;J};��]/R"���<�)O>�럶�t���C�2N�	�'��߾���&�<ճP{�4��\�Rm��~tw���������k�E���F���6��bPE��>E��R������L_�v���;�X�,e�����:�S�sA��j��_�z��M��=��N����^ja�l�^��MB6Y��DW��
m�K�|�K������ǦĽ��h9�-a�,>��/�;����|i71v�&!��]h�{6�z	S�5�-;4�*��Se���X�6�Xq«��+B��܄��)n&��#	�X9������b����#�/����p �{�NC��-Z���;"�\g��pd�ᯪP+m[�2d�<̆"�<I�VH�~��aKK~�L�,-��,���_���;qO��0b_����D�_�.��"&C�n���pi_+����S�B�eOKY��3R�:V"q�ؓǪ�O�_��R�Vh?�PpԿ(��"�@��Ec���Å��N}�s�d���}��US���֗!���й��X����l+:��9�쿆D��c�4i1����v�����t�DX��x#��)ln*N�Mi�{5g���V��ǖ��si�o�f��l�)(�ߋ��B�_kH`�V�����"�dbHCU��s��T���o�Z�e�_
bV���?��Yq0n��6�`=�k���OAw�yV+���%c�)^\�N�������Fd]@:ȭ�MZ�4� ��Z�ҊG��;Ӝ�l�j"V�d��� 7fD��R����n�֕��&�_i�ͬ��iD/Y��e���ȸ4x��"{V���*r�6���-�"�Q��;t(tڇ&�&5�k���16�Y6��(�7� �,� �6u��rN��|�w^�=�\�U��������n<�..��@,DAa$��J���{�2����:e3���:�^����y�ܨ�v�P�^���稨^��>���y�#����ߘ�
3��Yb�݈,f�Ε5�n��TO�GT)��w| ����Ѣ��ٟhQ�2�����0[z'}'kX�Tx�.��hc��CIj�F�bZ����|A6���u˓Xr�-��
��Rr$Z䲆'�	�ͨv0�B潇�B�K�.N����T'�;;�E�iOmV�Cܟ�U�<$'kB��˻���b��[�$otl�s�So���bzu�Òhx��{$x�S��Ă���� HA:sM���ឤ�g� ����Sb�9�oJKG&��v>F�<>��r#}T+�&����W�)�:'l�ɭA��Z�/&U��a�����ZѠ���:��ġq�5�h�]~���T�����eO)��M���K�k N,n��oouQ,:k���� �R"��ЮA_	���ٸ�w��_�iaII)K��Rۏ��i8,æy!Ʋ�)��TVo�����X5^ƺ�.~൰)��=�!����&�٤A2>C��4�}.����5�gj�����5N�Lo���@�\u��2.�o_sz�:'	��`�K��]�e�,g�T��#�D���`�쵷O�+p�]Hk�N�I�]}�Ҳ��WZ�'���Ɓ�8rЛ�B����w�+O�C[�?���*�9v��ڐh���"tVᖚ)�4{�rL��|��H� 3�`��y	��K�/���A��D/�6$�-'F�σwQf7)�"�H-�L_�_r��<���0�p������,2%'8jfi�G����\�������)рJ`7�)(���ފ�
u9d��+������.6���(�6��moĺ�{AΉ!��d,>�7^�T-���筬sS��[%�p`n���mۋWW_X�m({�3$��g��N�A1 瀲��C�]D��~MX�ܼ%�����o˼<d���@>��V����4
�Z���L��n�2�V�_^��Ή�hr��V }�:Z;C8
�� lӆ�>"�-����p�<z� ��Y��Pa�����r]"ٔ���D0��)O�%�G���*V�!���B<?J�,JލpMwtW�B���б?�w��]\��T��Lk�e�h��<������������}.�z��nj��y�Rc���c�e��*7�~����	W�~-����L,��Usvq��v7%9+9/�O�kA���� �9��(��[|��/��XJ���Sl�6�x�y��t,�6X�Y��6�+����]����@��Gȏs�T�%�u��ٛ���� J���g�{z�ɲ.TS��Qi;���|��U�-�VeG��h#��5���"��"c�3��h�@a�w�ȩ-��F҆��z���!%�3o�������al��<�ߺ	d7�>���;/z�o�����\�e�6���\�'�v���3�+�FT�/Hpe��V�\c���L=C���������4)8/��V>�$�xj]�4�kʐM�3D6�t���c����I�����h����p�0���OW!�����#������e�~J*�W��(������}+bg?E`	fMi�/[�zi䱆�xv����TA+^��IO�˳ҝ�dl��T�ɴ�����W���{�-�"��03���q!{`%�G����W�M�:��J[טk��k�i��p��8$��$o~*a�o��=���xl*"�;��XtƩ����������U���.v,��y6��jp��f@�)����x*%��x�'�6u֪��6����p"y���?a��7��
��9���ٕ)4�QTW!_��#��h0͝ow_ŊRZu~�1}o��g�*�������@J�0�/��.%���9!*�sV����^\Ű����[QU����>m��'�Ѱ�`,���>�qpقdg~s^�U����%��=�9��D������Kb��c̰F���S�q#�3�#�ȯ[ɵ�#�&�L�͒&������߀H�b#�pqOȐ`џ�{]�N.0{��CS8P�=&��q��uF@qj ��f�<T�z�_���Υ����7���0��Z�C_Ml�ڟL��w�������e���:��O��k"�[~_���%��EQ{���Ф�߻,t$DE��m�o�Z���� ��/�=q����%�ۓ���U�Yw�ߚ0��-�=����P�cv�hY�z��ܴ�L�C�a��w��%��8��7f��ħ��=A�S.`Ki-�M-q�����$�P.d�dv'�ab����Q�b��:�u��u�)��W�˺�G�V�iF����j<^�:�w�\Yb@�k1����}�nO�q�qƗ�F_�6&��#U�QW�&Oz'@V��G����~iу�J+n���8T8>y8S:��D������yt0�'q��D(�~ID���9��Uѷ�
��@Oq����nB0#��ln�3�{L릣�/=mo\)��CP��m���ާ� �D3���DmP:�����,٦�9g�����׬�����J�ol�Y�]��9�Uk{ׯN�Q����&�7YE��U�%S[�É?�wV���NFn*
�qt��}�Z�o�sa��Y��1�H�K"�.�7Z�Q��y}8}ui�$+��F"�dd�Q2��H����]ty�E�-���]��_��U�1Vl�?(4���9�$@m������b��Í�؄���#.�5����׋�
�WxrEE�F�w�٪��崌}CMn��w�ԁ�[,����}��ů\EQ���?��Ef�ð�"���qK�a����&�.�i�?���
7�sϲ"�����?7�h�>�vkk?�?w6!%�L�ԉ�D]W�u�N{���P��ǜ�чY�5k����_.Eڔ>I!ϻR����;(Xp��yy#���u,�{s'p2���)j(�	��W��j�˽�� 18l4\�R�}ƞE'8���HWJ�D4�hUNY�E��#Ś���7m�ΎX��P�o?��Rn��������p��F �\C��]K�\�z �����VL��Ha�|!� �UZ`�	'
��>�;|����Yvhv���C
㍭Z��y*���`kb�n��ʛ�OQx^��N}*X�Z����i�����{K����
�����*��P6*�Ш�Mj,.,l�+��K�}�лɃ���D�����l3F���g���a�����W_.I'XP����8���qT6��v���d`�A�pI�8kT-e�.��02���rY?e��p-�Uނ�k�
C5���Nn#�-匲#;ڂN/��.�:_����E3�08�4!��}:����()0y�������s��<w&Z�B�smn��b�{���Fͫ��%���`'��W�q�?uۇ!ǯ@H�
<B��ɷ;���]��uTj�~6V{�2_Y:�3#���Z�H�RS�� ��w��|N�-1��e��%��Fg�;��30�Z�7�>�oD����s<$8]7�8b��40�C'<�$7�"0ʎ�������X�a�N�z�������u��>���!����^�C::i��X�gi���4��8r�`��b�G�.+[�Nd�B^"�WXZ��ױ6HW�?�IcH1��\���q���,�u��̓����:s=�[��	O`����X��>�֡����� ���Rv�t��	���F��1�ζ|�w·f��6p�rDW��C8���� ��7�zz�$���갤D�_4�a�mpbD�� #`�HD ����a�6����ǻ���dm-C>� Q�[��#�������<KI��+�[�VT1閽�Ѿp�$������`�͎�S������z�����K�Ջ/��jdF�p�\� cM ��T���Q���b��״`i�C�.��K��׿)�e,ǌ�q�F\΄Ie�t@�p��,u��,�4p��cˡ�G��7S7�KK���|ۓS���B:����?�_Y\���60.)��)GւН��KC���qϮ)��2��3�`3�@�ISɗ�=-��N&9��ʊ�z����x����`�)��\4b�.�&�d17�IbI��e���tv��!`�E��9
ѣ��+����'��'*up|詷����<��FR�kfN=�
���jPs*/���T=�?�!���F����,��f\��39jw�b���2�gf%��l*� ��&*UZr14��y�S��f�\o��V��&"��X$
b-�T��\A[�K��+��Ӊ�r��e
�~ʧG���p9F��M��n�98f���ݶ��R
m����}�W+"Ռ�?��y"�v�Y��ƛ����w�{i�q�"�7V{�Trx?q;D�E��E|�!6�E��yyz�!�{��K��àD��gcӊ�|����@O��Y~i0����l�2����'غ,��={.3�Ik�)+�87(\i���2	��%GBE��Zl7M?^�Q�%�}3ٝ��OF�<}r ��Y�:��"҂�� ����W�ᩱ��g�z*�	� �@\J	�Q����n�s�"��K�v��M����}�	����,��$_��P�0�� m�$�X�B�atiO&^ϩ��-X,�sVҙ,B�� ]�"���ю(����& 7�J��ojfs�T71g�'!��!>���4e��(�v;u�7Wܲ����3H���B�ذL+sF��:ׁ�H�p��U;��#��>r�;��f)z��������eC,O�pU^)�ܜL�؆4���&�>�k�s���w�a�:�}jYnE%̫��T��M���z	�D�P`L���K��d[������!ag�M�a��{�<�R�WbXq{ ��3��^��*��φ����iL�Uc"�P��zl��M��%�:�������"��c=���	��3�eI}��p82�O*8�T��ec^��f�ỳ���Җ@�2Q�T��(F��u��GQO��W��	�s�N�^D�!>�f.�C�� �gS���C3�q�$�v�5w�"�c������3��Uي�
i�1lҿ�K4������#eƯy�$��������v�g�i�
�&�4����_�� m��)�d| h\�e����i�#���ۅV�}Լȃ���#�,���-�~	�G���6��U�YS�c���Y=��Oo�<��}4y\:e�~��0ep����b{�[d��!Չ/p��p�s�>[�qy/�lgQDikV~�J���7X�շ���~a�Ro��>�'���S����]$��_��6>�W�5e���ۆ���4�ۖ�����D�r�¼��/�Ɇ���N �O~�uZYJ+a�
e�Q��ɰj���󫤆����QOcl���J���~_p�*MaW`"(�1k����4�ЇO�U(��O�	w�	m��*A����L;*��bl�"'�5�������#��׀��:=���AU�?�̞_*�^B���sI!��ؾ��}�o}h�tm� G�	e�����_|zb�+����t8?������h>����?�O�,�j��c��Aĥ^��jþ�i�����!g�DSφ	Y=��1�-�m���g�1W�cM��-��`�����U#�)p��,�7>��N'��|��}t���f���$sd��d8��Kא�UFg��=��BWZ2��B�'"�0���՘f��DVG!>-��t�۫3�k,�E��8Џ���`��`��s��1���n�D���Ps��^m�ys�ɼYxEvoEķp����8���W�ĭGb'�&�\:m�
|Wk2�m,}8��i#�(J?�{Ÿ�yMꎸ$��KvΈL1(�j����E@�����;�������w�����Ҽj�[M���X4z=��Ò>z�`@�,0�?�wd����H�s�Z8_U~dZԅ�E�����*3���d|l��bBX���O�>xq�2�C&�f1��
�߲G���dK����1���,_� �<����4��g�`�E���*�[=s��tNY��?�2�K��_��k&W�S3�/7G���J
���h������8��1D��}u\H����%�~V�Ts��M���9�����e�'����&Z�����xh-L��� ��y<>����׌+T5�74�cGO�G����o�by"�wb��^㢎�oEWu����*QM\���Hޖ���'_��9	*;c���XM��mEu�$K��?��dGKp��Z� .�KPt��<*P��1��"�΍Z:����P���Q��͊np�� n�q����za�<إ�n����o*�R�F��g0<�sBЕ���$(d&��ѻh��}1^��X�aT����w�i�qƜ"
|��?���'Q�+�c�c2X�r?lR�Ӵ��iL<TefW�`�i��J�U�Q����I�_T�J!-¨l�*�7�I	��t�����r�bh�ۈ̎����^hQd�A7&ݘ=���Ԍ5�T�fs�+$n=��ֽt{�h�����%p\�p��c��P�7����L�5��󒧑�x�w5'�s^k����e�4-�x�>��D���s��j|m�B� 3B���!����w~I>Bb��8���4�}6W�H��8�|Z�栊�Ϧ�E�>���@f�FRr��d�C.������q�A���i2#���!8��R���3x��	(��.l�\�������5��5~���(��Nd^�g!k"����v2-��$n �1anu,�LS��F×� �8(�2N��RB�����U�S��(�Qk*���Lw��f���A#%"%��jL'��YG���������Gk�-~�� >}������ �砒9����bj�[d0$�Z���M�,=?��h���y��*,�K|��ìS�'G��Y!������?��E:q6���	.$��M�	.~)����#G��oY�(u��r�w���E�=����w��)>�wm�3���\u���{`YX+7ʽ;CY(�p9��@��muhP#����S��3��}��(lq��h6(���9��u�a�V�b���=0��;�X�������Dpt=��w�f��\9b�*Fzg���KC���Ź�HtQ��V��