��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����rhhm���%�ñ��\X}"y�GM8�,�eP��:h�Z�{|��L�~�t ,������DN�F�	�:j-��u*�zn���{�h^���C��zlC�Wg1MH����{[�rx&R�+0,@Q:/��ц�?yU��g_b��1���C��M����훅�[�>F�?X�	��ϟ�]w&A���E t��/y[�x�b���튟Y}
�]�w3cGTe�����F;;�A���|-�¤��^�{�w\e�+����"-�v�E�`iӆH��n1��Z���Z"9߸���֦�}Q^�t%��$w��=6�e�C�?'G;n�F� O�9�Y�,Q���X^��"�p�񔺖�3ЄQ���W*�'0J��kq���>|6d$j���V�+�{��Yf[�( ���_��qd�pY�o�4�8h� 
��ɴ884�|�?�ͦaJ��>�ggc˲>�����^����h(�\�<�݈�*��� ׋�H��[�<��<wݼ:�۟��k�l�a�Y(_<��"�1i����2�,6�`.�q�l�@�/yŇ��NPLn�:���U�ǡx�]�:���zuѓn||�����HG�ρ�t`���:}
�$8�rK
f�6��U���᷺{#�>U/�`�ՠC-�K>9_���k~��u>�Z�n�W�	׿a{��!��	Vn����������6]1�V��'�3���~���	�M���!�Z{����~��2p���I ��7�Sl�6T�"P�a���J��f�v��&��oy��鼢��w�gUaGpו�Z-�p=p�G�+5�/�Я&��:�ͦdz�ѿF��}^��i�n25m9��羉���kP$��'�-1��d�ۀd(k��?IK�	��_�/��Y4�2�d?;@y!��XWSÝ���ɫ�s�t�8�@����mAS��F�W}G��$@��ꐮ�y���G���d�tcϢ��Y
��4~?.�(�8)�1L�`���8��B\|Wl�̭II>�c�1�8pV㏴D��p�q~_v -Gt���">%���Tg���D�'2~�����W��u>�c�1����i�� ��6��?��� P�m�bkCGj�6�4���W���v����`?�f/&���k���a,m��t�w��������A��J:�4J[!˳ElB�繰5�dk������I.Og�u�pm^Vo!��:�<^
b�/r|���F�A���Xڗz1���'�����:0��,̷��N&u�!���Y�87o����+��&?�#D�ok�� ͺ���ۊ�}������&�:֓�T��^��6c��r?N5�?��u�{M ��\�����+5Zqkl�;5�"��!P�%�8����?��uۋdX�_�;��WK��TA������[ !S��2H�S`b�,��n����r4�/܌ɠO�Y����ɂoT7n9���S����Ty��EV�s��q��`(�[���ج�w
��6I�2K��Ŵ&��/�����nK�wWFQ��t�t�Dy��ʩ9�@	KK:Z��5Yd�@#ڒ<�2�~ާ�p��p���o]T����|Eu�Qq�R\�c����%xOx�^��a����NU��sMH�� � &Ǉ;��z�V�. ���G��p���{(E���?%u��z�QK/o�����Zx'���x���\���9�0iG)	(~���q�0��x���G�5W)�p
ES��aDǥD	EwxˀƏ�聬�~_"g����)�}ʤMb+��_K^�LrO� �3��<��YhM�ǃz�"1OϤ�'��2s�*��v���L�T�$�iKb).M2�K�0���`��qK�[�0ج�
��1��XL���q�Ũ��B��l9�|>(��B�X� i�>rԟ\��E�U_R�5O�������˼A$����D;��[� ��#�J̭�������!��ybk���A�4��^�Q9����}�4b�[�w�4��{���p�W���9$����|_���wR<F}~���	Iț?%�-%}4O@B���Sڪ^䠪���9���j�L�#�̴���3~�������U^_,�\��@��cx�Z]���<��G��Cw��JQ���6s#�?��ꍣ����̞)�,	9���&+Qߟv��.K�'�ۚ�*O����
��V<� B�4��JȾ
����9�rE]J�e^�Q�T�stO�w <�n�m�}���� �z~���df�YkK��ս+��0�V��:�=�Un2�+롬��C�0�RRy���Z�����x�T�D�+x(�AR��S�Ǚ1y�uw�9dm��^���X��c�s���L�h�u0��ݒ�qAS��py
0��V5��E~�O�X�g1l�5�����/��`��yL��%����z��:�X�ݤw�b����)0�+���1r�dbhJMG�0C��L��}kep���7�}Uv����g���EP�?7(����6�
A4���������k%�A�Tьa���m�gj�Ϡ���0l��,�H���r��ܾ�+�_�i:���x��\��4����־��q��\}/�(i��g��z�������1x ������ZI�m�K<$�棾u����vQ��:�ݤv�B���:��L�$��7����Ȍ�}?#.�~��_K�<f͈m+��\���#�g�2W�xdG˴ ��7
��jv�Z��z�f���/���e���o/��>�`v����l������&<M^yz�p'�q�S9O�U���Ps�J�d��������r���h�X�\IJ*��Hu H{�ø��4JYb2GW�Է���w�k7�7/pԙ�$�D�J�S��{F�]��Z����h�,���,��6K�2�F��@��	�fR;4�����K<�a�G�5,����4ޝ'���dyTB>�V*�O���w|<�YbL�Na�){���*�Tv�f�D��WTA ����V�DP����$��(=s�g�P�bU.H�P��n�}���'NAG���R�T���*е�l8�#!a��"ITu#�g�e3�K g�2��E��:�B�� ���s�4F�n�t_Wu�H�%ɻ�	
�!����-��/�3����o	)�h2ܗ���y=�̒�խU}Q�>VR"f�AY��X�O+1�s5T�nPfe��#e1���(�8��f�$�.�"��t����վ�Ϲ'(�Ѽ�s�9 ղV�gH[Խ�o�j%�qѠ�euI�!��X�
j�`�)ǃ�֋����H�����9֓R���P� �(������)<{ho�/�B�Zv�� e���(�� ��@~�"��!�T*�eR��\heed�!��Ū���pno�8<{'"�I����ĥμy�gJ]�'(�0m����=�����5Gڟ:�T�����Y��6=����̜-7!�E�<8�6��Q��T�|N�Н���BP)��1���q��F�@ 1=
yl�H�Hj.�-W��"l$�ĩ��kh(�H܏S�Ao�x	��21�D���?D
�(�e0��������{D���'�R"]eP\O��d&d<t��������a[��p�/G��֌�wƙ����ElM�uu{��Mj��(�4#)���[M���|�P���Y�R��s5j�>�;'{Pei��G���Y�mR�t11 8����XC�--�+����@�7Tu�r�l=a�d#;�ɰ(���� ƁW��s~+���v�;@�P�9vϛ�>�w�a�n䳹���x�l���W�V��A�Z��X�*I��E���sj��0�{Fӿ���+�a}�z��%��qL��m�7��O�Q:�g���K���$�
2'�m�x�,��T#���5@���h�垐�9S�"���X�7\�j)��<��;�iU�0�3탱S�dlS���q���Yb>#.��3�X�w��M��J�~ha�:L�sn����N63���-g��R%)�4�yz���j�9��w��O�F�r��)B|+2Kn�Z�9��bs�<��+f.�q�2s��|n(�p�<:��� ���2	�`�I��}���M��W���{��byw��+� ڕ�^��3���ZX�@L8&H3�5o �aR�0y�晫�p�))�Hp�ȕT�0��c���Q/% ���j
�e���se)u6s[�=h?��&�B���%,��M��Z.���7�3��j�C�d(����`EF5�&�I�y> �	ٟ�x5e�XA�(2M;���Y%,�g���f�fQ7�;�e�	=�
	�w_ۂ��-�ku"�s*c�Yȯo�O����6ҋ�Y�DZ	ֿ��7���7`s��df $���	��#��;JȆ"ͣ�����P�0JK!h�簦���N{ ?1��^��[)�HMt�Z6���~̊�Ζ�m�A���������4��CɸE&=h����a�g�h-!�P[���`�AݓDC��93٘�p@�%ζ��SK��������dU����U���k�@b���Y���?YH/ DS"��Z��m�;��z�B��ѧ@�&	+���M�:�Q���R{C�RG(�I(�K��2�]����ir�|�"�D��	���XH�J�2��7Z�)]�A�ͣѯI��P���h�*ڜ�e!�}H��7ޞ"��D���L��;�7��M㨂����K���+�$[Ŷ0��Qץ��9�S0 Z8���D�LF]���%�D-����"J=�#C�� N	�g<��
8�_��!�`�f�����Fxj����z#�T��lǹ�S<�`��e�Fm+w�c���蚵C�}���X=_�֯K�9����Fݹ�.e}��zvT�v��l���BAN�x�{~(��_;��3>�m�_�O��6��	faM^yF:=�����g��u���D�fm-Aa��!{2cU9,�9L�f�d��Ǆ�M���rJ|I��Wm?�X
\q�4^v�F;7G����y�ʑ3ۇ����6��y�ڿ䭝/�X�L�B�td���?@y���=���%���ck-eÁ'1N�X	����^����H��b� W��Q}M�;�@�P��k�D��u.�Bz��A,؆M]��;� )���z�{�:&��}4=%��rT�@K�YI �ք:���3C���"{�V�o��q�a�@��v�^�+��e`;�� u�m��;����������"��C�!R���U
�B���}����Wڨ�i-c�;��Y�GHl�D���)�l2y���c�o�LY8�K���W;92�̅�����S[}gD��P�f��Wow�%�Ij�u;�w�m�B��bkh��Le�UO�u��';O(�Ժ�5��Z�\�O�u`Nˊ6�R���?�o�p"e8����xi��E�j��tE��W#��ڌF�_���P�q���n����lU��v��6n�@����Պ�������Qq�E_���P����d�Ԗ?��6���G5Z	u�se\bT�i��)z&=�;V���܏T2�n�,DM����7�	YЎ�4>1��%��-ni��[�{�D�L�2z9�*q��V��g��D���UH��FoI׫u�?�����)3�
�¥UO��"�T��m�X�����]��d�*V��ʖ���R�U��c�k�>�J\Y�W��
݊sh��	���=�1��H��;��>�!��"�$L�״2�ѴR���R�o��&�A�wիGߎ��]����#���V|쯞���L���Q�$��/L��mд,wH6�ҿ��"#ǣx�z"�$ʖ�����zE�)��U�?����L����T���x�+�(E��7�?��E��K�|K��b�a�G�EP;44 EЫdߗ.�����gZS[>���Qa�.dym40�k���ȕ��R�*S	C�b>G�VE��X�;)�c0<�kcT��9R�>V��%�ax��]7�s1�U�@���A�Mh�Y˺/�����7��5�(���҃�3�t��s	Z�c!�S��?����S서�����?=�4�3=m�~Χ��Sq��<"�౛��z_�`�-<�ʱ2~(]Y�4l�go�h�?3(��M^`��Mo��-v�֊��8�`��G���%�$S��b�̈1��y��f�$\���w�׾�#�� w��/��Xד�4ak���׊[�Q��x��|��~*����*�#�����RS�4��wj4J��JO?�%��ڳ0T�*K]�6�"k,Ԓ�!���D�evz�o*X�PBe���T�%A���	���Z�zd��ը�?��W���*���i�����no���x)�V�L��k�5���7�T��
.)�ϩ4.�UPى�c���C�A^��[n���ˍ�,���;� ��,�6�KS�M���՗j��jJ�B �*A��_��='�J_P���
 P�ч��X�o6k�W
�2��\9�@�~U�(���V��9 �U[��ͭ������Ђl��v�d{���>s%F�WiDo�$@��jg�AJ�=0����)�9@�4�~��sxw�%
lUa�����}B�R! ��T�Nڮ�v8<21���?�[�Q�h����'�dT��xb	�UZ�-R
B&s�nz�W	�d�Պ!ߦ-s�r-��t���'���tan����Hd��D��RM/wo�M��/We����~W\��<��ʦ���+�(^<YE�Oo���Iw��d�bs�q��Ν_i-�X�����GʡmM-����)F</i�0j��X`>�1��.�Bjܝ���ԡ����%�Զ]�Πm)�\���B�h��zV�e�M���Ӕ�Tj�c~���瘠-ɉ���a^t�z�*yejq�<�(l����H�bD�R�/ E�5�� �)6�$LF�(�e��_�����6�~1�S�>ݱg]䨗�����-�%�N��\�rö�~3v����\e�LX�0�9��c�Rh�	���rw�E�<����5m��x{�J��Ώ��Ն�k��@���ZѶ[�{i��$qE�	�"��cK^�"���q��q��K�=��]g"7��:�G	�_�������nO��U���ٖ;.mډ씼�Ƀ��KD6.*;а����l}���[4(o�����I���`2�o�l��T�E]��	.'��Z�M��������{�)aC���o7����7awYh�V���x���f��>����y�^���c�S�f��%�#~�"�0����9�DsfF>;��Q-H�5g�z/|�wT�` 0�Mk�KUO?�ޏ?�\������4Ώ��!#D�p��Z�r=G��ʳ�X�����O_�(���w����o��zNG�!�]!��+)����a�!�ؑ������^�X�c�x41ay3�����^�� W��I-:�_�~�9���U/r���]H7�z����(�B�4�!��Yj��,�A��F+�� �5��o�ȹ�@%�x%���f+�Ou�Q\S)HK2<���M/N��B=��Q�(�����]hv\)�_�6p�2�? n�
�F�\{��f����6T!�]��{̀5��_2=����N��׋��ؓ�[��ƍ�s��dy�<�:�Uhe�����ON��.0j��A�C-��&&(PM�n�7�ŚAU�
����e�F�lX���Q,��w�ԣA���e:��tg�2����oN챸+�r����&۷>wi�����;JƌU���w%5���+=�B�M��>�qr@׃�̮����>: ��A��S�lٞ<�
�ˑ61�|�:�gpYd��G��=o�y�Ѷ�J�~ ����ݖ�6a�;�~K�.t�������+(jt��QjV9h-��3�06��ך"�fG8a↧�l���h��J�`��p]��_\�M���|�.��j��_����.dv����t�n�(*%��U)z���TlM�3t�w��v���>�sO���*tQ:|x��I�8(��f�k���I+�u~��wp���H����Z��v�j;/�W�UD ݣ���1I�8ˋ�����M���ka
ζ�r4��c��7�HRR��}��$TJ�+~/{�������Ox��7��b�w��E��~�|=j�u�R;����g��������%���+������$b�`�[�b�+�c�OѶ�~�-��_Q�����P|�9��M������wP���x�9��jc�S�W����U�4�$��{t0�btܖF�f���{�v���Q#�f����5Q�&���p�����d����������`a2D~7�U���xG���-�c��bǮ�"R;���u�D��%]���=�
�2HQ�c|8B��N&^�w<��X�#�͔1��UY��
$	��p@yꀕ��X�Azd->^ �G����Q��T]4��j��௱�Ț�3�C!�"�S��b+��[ꜵ3�ɔDN&vn��D�
�^�5��`ښ�h�콎 z�-o���W��C.��w*� b��=J
�]��#���[�A,2�w﮻㤁u�)p�YL.�-�kO��fs������5S@�Gzp����V~!� KU�b�BZ�W/�|T�S���P�a�.�K�'�Y2tX����T��7�'
(��g=�2���$���+��M@Y�%�������[
��"u�U�8��Ɵ�㜙͕�#�;A��x4������]�Y�ɟgJ���&G/8�W�	�����e�נč���gl�@�_W��e��,�њ$3;0�{/�%q���>�wC^���'8�|0@�q������N1 %_2�g�R)֎�R_qt7VN�r��y�v|�>�{M}���tx�:6oýj$�z���D��/�f�����A�I�����]a0Z��T@�y�:�DC��������3��U��	9pg��7f�)�U��/K�軡!j� RG2��Τ��uTB� �l��̬�4u���"Թ�����fI7&�N��Y�|���#cٓ��"ȡ�aٝE(U�h�s���1�=�$�(���P�!��2�ҷxVS�w����y�5,p����|*��(�Z����t�/���1�'�^>��a���|�̀�:� [��� .}=�`��`
�[�Y�V]�����ͱ�h��{�����7�W8itjl�q���Di��u?�,�~�2J���4l��nJ�H�3�_X������%��
/�K)�ǘy��F��;'�����x?��3#����S��6G*��K��"�E��Fgݮ��kB0��,���ԛ<A�M�~���3��[f�ȟ�p����H:M�2��ѻf��9%rC��Fڧ�}�����ۓ����\2M�5!ep�k�U�	OߦCڞ��QA��1J
p~�ܭ}�՜F�K跛jW����ȁL�pK>ōj����T��M`j����RO�!G���t[`�]�'�8�^���4 ~/,Н.o�0�������s�Y򓐞��q��ʾ��.��.K�`Kdt~��U	�s��:&kB>��&]�y��U����m��g�0� �Y������YL&��,{/�e���]X��>�Ȧh5��x��"����-�S�+Ƈ(L俸E+XY��^uV���l����	G͡��emt��	��F�R����UUM�$i!��룀�~���HK.�M`7��d,�L'�u�d~%�E˙�N�t9u�K�ɳ� �2KBG�5�-@���-J�Prg���]F.�����zQ��"f���.���gKκ>�g��Q��EG�z+x߮J�,7%:��T��oi�Sdf+�à;��ڴ��\�pG�˦��_b��y֔�Ef&��� {�(.�/% �s��κ���Pc���Nm����\���yd�j�Z�}9������ׅ�x��������u @�w�9.N����q�?���lq�{�FtN�<L�GGS]R�.��{.7�)���6�u�����2p���L�3Sg\�4����U>��uD�|��|�`�+I�^��O�~�$K�4�u�E��>0"��r��S�<;�t<�b����l�<�������ҋ��[��5,���I�{�ٹ���w���ף�M=ש�,��' �˶s�Y�o�G�!�6��wڃ�?=1�G5�>t�*C
ࡺ0r��-�>�E�~���'�h�\|��P7�i%5���b���F��VF^��Y�j%�dMҀ�!�cV-.0��a��+��ϯ����`����8s&�.�(��g7pZd�e=@�&�hꑐ
"�OֱC.�������}/B��B�����3��!]^X�dẅ́�m��TG�5�	�D����7wv���
��������!~~��ˤ��l{@NV5���:e^#�)r� �D$߷��y`��<:�G�/�>��V�Q<� ͬ�W9MI����R$� �
���;�b���>��������H���`M-�`�TyG�I��0�;��j!&\C+��{f̶���e�4z1"�NP���6���'t���m~�7x���Ԝ�Du��ZuF��`���J��ʍK��e~.%�������ߪk�k��>y.�F%�zKN����$N���ٻ^$�7gٻ`�>R�愤���ޅ�aA*&3�J�AekEAJ����"=3F�v.���z�96�W�JB��T`vjD�yO��E�V`�S�H_�QL��� b	��Z�0 ��'���.{����!�B:x^��%�O����J-��cq�� �E�;p�#��}�Ҝ����7l�+���H%צY��
]�K��1� ��hp�=�j�=n,
��+�qފF�����Ϣ�E��TfR��U;�w	t<�̌-=7_;���c������,/��I�/:���#t�2�>k7Y�Sf��y�i�Dp���n3�հFoM{n�s�i|s��R�"v�ׯ�u0%`�,KHBڠ�����-�o����y�V��4�N�XCM,\
ݠ�WY�U'Cv�`͏p,����'jL���-U'�K$m$7R��.�<v���<>'�&��q����6)/U�	+A�y���k�]}��Py�^���6NX9Ѐk%�F���)U��N��z�1�S���&�|*x��%�E����_��A-���謤�ۉ�E<�@.��<v�FB!�e��ؤ�Z�h+�Ǳ|�X�u���]$r��r�F:���(����s[3 M;�4;x���*�5�2W� �@ �P{Rk��? ;g�r�s�7����A�PG-I��?�C���'V���#u�2G��a��M��L�	W�Vǁ����E���#ֱ��\�#��x�d2Q2˸[��G�_UeZ�ks�_Jɉ'	<:�А��Q��qQ����������;0h��̈֞ی�������yzH�5k ����Sk�?������	8w�:��>8�-Z��+��F�*�ߠF����ꪃ6��$mrSMrןy��9���+�V;Z����uX6�iJ����D��@.4�v^L�&�J�On�R�{,P9^]�Bh&��L�Ob�Xo}E`��pw���'�=�X<Q�)�O�"�g�2�蚵2�(C 9 Ɔ����T����_a���Z���1�����tGrժ���j�-�Lc�ҷ�+�1X� M|������l,G���-к��=��OYV_Z.�{S�&�K�^I�F0ϯI��T��
h1H�L&I�zv0j�?���Џ��؁Z5��L�ݙ�*�KJ(P8��"N�q����I�������V@��'��E�R�.���^
%9d6�TR��^A�AB�栗gЋr�V)ݾF�X��_\��}!��א�T�B׫��8�><��Xv�v�*�2$PK}�J&����VQI��&��b� 	�&���z8?�8d��"9,�_�L��\�ź��Z*x����S�":$��q���	�{��'���*䡑R#,����`UE��ҿX�)��08�4�$�E�ݴ�-��G��E\H�)�!���*�|=W5�,x�<o��'X�b�zk�K�*62&���z�&J��\ϯ���b�|S!<	��xxש�Ž!OT]�$�6�	d�[�f�= CC���ſ�[�GuA�O}j�qr�ѩ� O�Q����P@ёn���1~ZU� ��5tv.��ϞF�7��C�ΐgRZ� R�U����3�.,1ć����c~ <��"h��f�&ɻ%=���p�ܿ�Za�^{�@�u(���qm��*�a���@Q�T�g�e81�
�l��&��{Xzskԃ�Wi��b���kl��q�ߊ���'5(���F�%�g����]�vd��(t�xy���I��i먕�b�MD<�3�;.��uU�B�b�I�C�>�Wy21�M�@�N\�l+3!�<�o���W��#��,���Z"Pjk2������S�CA�!��&ؙ=�*�ʀ��	ɘ`�s�'O�y[�Q�S1�}�L�Z6��6s��v����Hm�K�*�鹨i{�"]u�o��#�����)��6�L^���~�w�vId9��_'=J�t���u�o�{��T��Ǧ[���w���C��E�j`$Zj��-jjt���t �W��=��rY�2�?}������:LL��.���k��eO�PLf��&~�Y��c�e��8&W��@�d�sV�n����+.��'�����?��o��R��2��DVI��G�^�2�x�v�I'���W4O_����9g����H��Y�ލD��b$Υ����	7v�h{|.�z�6��ĝ@A{���_j	>������������]3���OA��3�lP`t�M�"���7p�!�ľQe�Ңa���� $.�%;?`���|
�
0�����Lcz�I<i�`I��~/���<�iIdx�$�Z�6.�}�߳�z�Q��3@�?����yB��+{��L��l)� T;���
:���D��j�6���azO��/�Q�y�P��3u��}|+�{`@2x@����Z�BY��&�K�Ge�(�7UYa���c�6L��E�,�E�����v�i�Y��o8��s��O�1#Èf����5�90X�&��܎nXs}����K9�����}���Fj�8՘#᷒m�鯹O�TrCFp@��^��Ci�b���ɪ���c�@Z�^����=�m�j�^�] ��DXT
9 �g��pi�ˀ�Nz�r���R�杄��x.)�<
�7ǧ1d>ks�	J���	7�0���)-\K���k��"p	�B
e˙B.�"��锻WO�E.�N5{*��RFB&�u�&j����Jx۫�i�� �w 4�zf"sIM��R9D{#���LY��=	�'j�����_0�X�ma<���5�l��	YՔdcu�4e����w\ǵ��t��a�|~�Ql�)�+En��?�4.��]_��A'�2�y�b<��)�lJ����L������hdM@zN N�q�;��2�_��i��'���7�S�����b�Qx��
��P��6�AD;N:���5�6];e\�7�3r�8��\G2�R#f��mW���_�`2B��f1K�7�*�+���Ȩ	'�)���m�|'i���*��/m7��+��B�R9K)P�s��������䮩ƀzs���ݧnȽ��!��u3�s�� ["t�r��I���A��x7 ��+ 8�t.��#Č������+���)�br�r��tὛ��9r�(`8�[[�}�$�Rd-��=���3�9M84������4W#�b�%N��ӱA<��\���)�s��*x�6�Q�`�ޝRi$l�-:�_Sm�Q��̦и�:zD�v-�=�1�U�ȉOI��;A��ȾV�ƚEQch/I-"@�N�����G����7&VaZ�]����F��f�%�������*�G��K�l_ �����J.�TA�~y6���H'{��*�`K�[n�VF��6k�D�h6!��]�k�U�?� �r�c�??��%���8GrV�}*���J�'��Lj�Qf	$$�퐓�3Q������}$j+����l���K����A��6^�Wż�U�Bi	��xkk�������7����F��@�X�Pƅviz��l-��2��֒���qڇ9�rl����1�ċ�eE����#��x�\�.����j�@n.���n�e�u��)e��Ѕ�F���}X�(���6���{A��v�[g�ȫw��͖kX�-Q��u���ڠ�F�� �p���?a�?��Z���	��k!��qf�;�:��M�K�s&m���g�A�a� V�����&{��g��m#�}#�[�,�<�b��j韺0nD��L��e��%ȖB���$+h�fY�}�C��5��k*IW�� ��.��.�y;�'�6��ݘ��]c��;�	�/Q�A>R������s2��X㎣�ڪ+�O��
`H� x� Ի�D�����hē����r笈�}��"� �ó4-Y�}AS4՘�~H�g��ܾ��qYi~��x��ï!�>^9����+�u��K�
+�OK�d�WJ�\�Y(��źP����[�Ƕ��SƢ�<�Fd<n�U����ƽ�T�/�sa��FxæL�i)X��pG˕��vN8x�9uy�}9�VM��.�Qd%�3�?@��D�Ɂ���	���(��P������:�(��C����vY
�F̷(���͝��R�A���r1�PD�)Wx3�DIЉ0%]�]2j���* �H^��#��+���?��`^�ˢ!����)oY�g��+�fm��1d�3kv�Tx�78�T�'֎�E�&�yB��]��>E�$��}4�W����6��UH���&.�#_�!����W�L�t�)f�2+�wN����ǃG��[�����n��r���-q�wYY�i��&�G�)���������GJL�2c?���%�5aU+����}�� �F�FV'D�����=�EdT7@)�mj��j)�ڑ�}��ݱ5pe�tca��{����	�W����w�g�����(�ͥ�?�l֡b����2!4�*�[2�/{i*�b��fF�i��X]�\jɎ�OrG�M	J��@�]bCQ���ѩ�X����,�m'�T���tMۥ����"5�k������bwb��	[��B����\�7��-G�S��щ:��b�5|/�s�h�l�����f$TܳJ<V��=����K׽�;�B�v��Q^��[���LwO�-Y(�����Hr1��E*c\��k����9i�&ׂQ�"�(�ң�k}�I�����`��^�J����(�?Q!�/�8�����v�Lz����f���8 ��2������nw�u��iH1��G�b�ܺ���G���Re
 9�����[�E1	Zk��H�xӏ��q�kA�:���ղ�H���c�ay`b�&~^`���vOR�H�t���L*��q��,��+dC�">�G_���:�-hlc+�4�������u�]wd}����WQ�+C�����?CVC�� \|n� ��Dt�歫l<�{u�m���˒�Qة�
�"�
�\Q��@��N��:h����hӀn$\�99 �=:,w��e��	�:<�eMb�v8ř� �8��H�m�빾��Im����/�m~,�>�bO݅� ��\���)�w�u.�ˡA�d��13CfL~�=���[o���C��I�m��x&���A�A��>ǦcQ�~��͵4v�Ve$��x3Q�ԁ����I`�-ß��XW�R��B��s��
b���]���;�Z�4�C�"����o�2����ό�=��Fm$<-�����-��ɰT�ܸ�%�*��NZ�ء�9�f�1�J� F}��o����$T�����+��;Fխ" ������P��lPL��~
Pc�XfC+��K��|n)0�Űc�"ި8�9�(䶙0�!u�o�����o`�=��	to8΍�f��ꀉ-߫��c��Hf�:W x1����LXp*Z���_�P1[ע]�煁�@&Gu��ό/��f �ľCz~��`��i+���J����0�B���9!��vR@W�+¸5lqe��!v��HҔ]�@�B���u��W���*�-JL�i' V�h�`y�Ya����o���3>]Sղa�c[���h��Q��D��d�jꃃ�[+��rQ8�$1)��%O�W0g����NQ,�Q��p��L���Y����w]R�&�g.�l�$��R��O��ny����n��L��bz�S�$�5�`�m3^� �(������d��WS���e���B�z�w�j���BN$o�$��ipp-�!z4-���lW���m�J<�L�]!2�e�@C	(J���pk�9=���X�^�����&o`>�d'.��inf���:C�.�w�.&��I1�$�+����Z[�/F��2�?Y�IԠ�F����2W���\��1h.L#31VO��a�o2>觅�l]��=/���
�$rT�@<l���I�'��EA[-I�Y㏨���e�v~L��(��u���ґ�B�/�,=[7���*�z �����yνO���;���j�.ҙ���\�Ӄ�ll��F�r.Q���e`�u]-��<��Є�0~��*jo�~�>g��y���c־ǀ����*�u��F�}����H�Y*]���Ce�óG.��d�l<leep�?@̦`Na���R�r�%��������[sb�/W}���]�jfNV'���-tq����ȸ}���%�5���ț�g�w�;}��D"0'����|M	�ѴV���<���
9�]�Ȧ�,|�)�p�cR,kk������<����e�NT�2˨�m��i�"��G��Xfxpb�K-R����Nѭ��Ҥ
Z5�fZ�a���x�.���9�v��h�;~����>��r��sj=�N����uKy<�/���/�>fOY�[)����� Qz��v�%E6�5�ܓ)��Ԋl���*�_���Zs�Q	ڳ}���VJ-Ӯ>���zh��7�Xo&�g�91K�:+,9Q��׵�Ҹ�o�#di��=�%mش��fY⨂�F�K>��wB� )�^�|�F,��ms��-`��gpi�&�qX��(#"�O�J�!���A"O2F�d���0��+��.^��!/��Y`8��K��+�w����(NB&?���u8ds����+H��lxfW�~���=�Av�>>��ok��
�&M��*�t�:ͣ�������h%�4H'�sY��ؗ��I#Ma��!3��x�Ų:��27�d{�U\����/�Y�,b�I�� $��PƸj��7�Y�0^���f>d�چBmpڤ.�qF����A�L��T�߮��KA�دMW���b��Cӡ�Ŵ$e�q}�ǳ��\��l�����L�Ze��hH5�kzC�Ne���U4���ި�s�k�^~:\�T,�͑v�l�|��\e�H���{�"��8�T�q�sCȊ��n�p�����r��N������S�Z`����-������󑋥�Y�Wq�(X��iJ8�����Ȝ��x�M��q�"�'=m� ��$�.�|��w5�Ǘ�'}�E3Y��g�P8VIh-�h�T]\���yXaX�Y�c���~-�W*,������OЭ�ĭ5�<4͙�����"���O0�B�y���C��<�w�wWud�X�'�v��{�k�vOz�|��z���j0��b�)��xa�{B{�\�~���Aw�@��J�]��b/��J)V%�0�F��>��k��Oa:�i5W��,ǲcٚ�V̹��\f�u�6�Si�3�Ry?�#�9���Ry��D2�8��>�����nٲo�I������}�r����3bN���|�_.I��C��Qh�oq�h�%#�3v�s�?�Ro�KQW2گ6������+U�1���e��h������"�#HNi�� �% d>?����ŭi�ު�* ׎�
[��e���K�<s.�'�	aص�(�QY{H��u�(������Yl�"<9/fZPA坨��)H��,d���S����|9Gi����|?9I�;=��_�5懮�����P������dȦeEU��^o>/X�b<t��Q!|s[�F�՝?Y�E�����O�n�6�	��g��-e-ɚ#M��YjNw���g��%�<,�9&�5*�O�+�=N�����f�#m`��Ը,��W��fPce�]T[�����{�%���d�Y}!=�����PR����f{�n �6�T�6��yVWnY[���f����o�G�>TST����{������♲���{�T����wK���G�HF#ܪTS1�K�@��Tj����M����O-)�n7﭂Wa=o��� u�����)B�U	�q�0�R�"s�y-]�����f#�%�����AeD�W��~�c�ͼ���cF�s���E�%tHI�ݵ�Y�/]-`{���ُ0��X��W�����D�E�Fv���5�U���5hK7�^O��"T�B�:-5	dMR�t�W_;���v�i�s]��^�6����ya�|R� XDZ#�w)a3�'��±�E�A� 	�j��/�s!��\ڕ�
�[.��z{Ff�f%�':~�E�#���ɫ�����ǦN�.ƈ���
}�}a�fγC
Ke�H���gOC��'b8Lޒ>�
}D�A(��3
T2w�	�� �����/�f�昸�� �t|	�~� �e;4���9�K����8��
��U�$��+�*�����.K��Z6�,���ZH�� ���{�΁g�NNo2��7��.�,(��u~B�,�-~���*h�ثQc�V��5��� ��(���LN�+��%�V�}�@8�$���2/I���( '��z党՟2u�㫋_���N���c�H �y�۩����������|��\��O�ߌ�p<~��B�Y3�?r "�����}�LC�hw^Wj���y�|0��ޝ���7��s�L�����Y$�8Ǯ�Y)�P2��|ű�Y�͏�TH��|n�] ZħW��tش�c=�ԌL�|ٗ
���]����ƅ)5��JX�O�pu���慷�v�+�V*wj�V��.���2|r�~�k�.����}O�`l^Z���T<������i//{]�sY��D;?���p>ۂ�=��J�B���ꀈ�-/����S
9p|(%�Xz2�m���v4M��A���\_�����dP:��,��%��%@�XMߞ�����l�%u�xb�7�a��dE�|�BC-���'�l��~;H��r��C�=ms^g���ï��<��v�Y����mR��	�RM�il��޺���c�QQ3����g���HDmOd�H1��4ix���)Z����vRtiR�{�o+�l������a�^"ۭ���3L��i�Dp�����O�ic��`k�P�yc�ߟbу�����s2�\�ޣd�K�El�ڳ����qQ�pk�w�0��?S;�XS�)�X+u�z������rF�1_��=>��B�����L� ���
?(~i4=� 2�,��C}�u���'"㫔�u�ͧI�ok��E�B�?R�hrޔy+r�⇟��vkwq�W��m;�d7q���s���:6�Le 2��A�(l�w¹�ñ�?�_�S�*˺�5:6�-v���F�KT��p���;��7�$��x'gYX>��\A-��׌)�_�@���̦������y��V��궻I@�C��g#�F��y�#���}��	]���y�bl��;M�KZ LfQgX���D\�����v9��<�P���F�"�~݂�[��x�?':^�҃�����v�����D�J�E66{	d�F���^x���y�%���ш�aa#����2�D�8g�R��M�#�쁵	�i�
ˡ� ��xAm���<��~� "R��A�N&��w��.���]�:�yH���
I��C>w���l�2���G%R�t=�ΰ�g�ꐮ+��ዻ@�ך�0J���8գI�����w�;_p�K����X}�D/�6���'��iwL�m}���,����lr��V��������-L�����{mȟ&J��3�'�����m��4����C�S��W��@
���qy���v�p�g#��W�fY־�*��]�周����.�ë�ފ��\P�'l(Z����EW��$�~cWF%�([E��L�`x�p"
ni�ʚv��G�ۏ��g_�!���Z�����d�U5�3��uɢ���Q��q�&�����A�������Es��:ڮ_pHH�A
2�D��-�)�����c󷴡Ns~ǭ/l|��K_AwT>N�����:D��%F9�]}	ҢEt����Aw�|���}m<]��5���=_v6�=)��E���`c���g�R�W5v�2�=��5F�8#�XT.��4f��yY��\�B��J�׵�/�ke�-U�З�DEE �
��|����"&;�Y?Œ�����?%��Mj?6Hi�����="b��8ן�W����%rBk�0��>K����1r�����x��Rڊ��hz�w�w9�\ST_��n����"�t=j����n�}I��8�l�ƘO
Z,9��Xa��Y�e��8��6w��~��y�D�RE��o���]��;�5�3M� �j���X�,�55>�m(&��X\�p���]��q1��٢Y{fT�2Oy�.nk��9>_:�����
��b�SfZ�CN��t̗]D�؇I�ɝB�fF4_����G�>�n�Abyч�9��1c8+̺cFh������J!}�4�"���d,/I��_/�;*d h�ӽr�U�z]��x�&L���aڊu}��ɩ�����T)OBV���Š�I�%��A݌t��`xm-���r����l�|z�����Z'}O�ϑr��1ψ��R�ƊѰ��ʸ����szU�ѭ�\>,�f���M�I��Fm'�_cao�@ ����s]�'���	Q��x1U���v}�L�����01�JY���W,�� *N��[�)�0�)�pٌ���W��0,��te�|5�ÏrF� zJ{���gk�@�*Zj F�
`�)�.�7��yt"̓�.O�c ƑXb$β���Y'��;��ʋ �;M/v/EG@HЈ��Uv]�[�a��w�iԻ!:Y���l
@���>�� e�7z���z�_rc2���x=�PQ�qN0��f8��GbG��i`6%,>6�9wƘ�=��i��Ѳ���0�eA�3Ȭ�ُ|�7f���
O�
$*1���W����T�&$K<xŪ���%�M��V8d��=s����.>�e9���I��Li&
^��>��@������q��Hc�o�Y��̍)q<1u�2�W"r�ʜ^`4{���`m��b�R-�͔ŀN�xP�d�_�=.�a�JL?��b��L'A���a�a��b��뉤�;�nr��-7;��	���v�(�;���� u�z�fb�eB��H%�z�3����E�D�¶��-I""m�g�1�9��+oN���q�HDVh�L�z���;;_��Z��)H��7�'sV��"�����)��+���� ��"���;*�!������4LN
���h�B¾'�7jBS�R��tB�H�R�mw3ltqr؄����.*"��k[.��t��6g��c����#
�w����jv�l��!D�L4_$��N~>���'���{�Yc�);�I7zg��,r<�P�@�[��p
�WL̈́W�%��k�;���[o9��\8�#jTa�ö�dŉ� 碔�So��A璪��hM@cy�b�"�s}N*DInh�&x�}�W楽q7�g��e�CF~��f�b5V׎H�
u�(�|Ua���G+�f�Y��۞��%�W�8�Q����$�g�.�~H՗/��vh>��KM�1t�E ǵw�w�������I��1�Z+Ī1F��s�42�-�l?��F���)� �@R�r�3-�5�'goܟ�L�����@=<'X��V,�M��}Dcq�M�O���$�`~�������#���[#e��N���4�����0s�{�߉������Ja�m��s�����������QM���PnL:g�ԝ"�Pgk��z=��j��'�>򾡦l[��%��N%�~DK1�?�O�Ϭ��.���_���Js��}�L`�j�(ø+��J�3�@6��.O�K�Q{�`����L=vj\�ۘƷh�!�|(v��}�9M�H��{__����fN��A���3�>A�,i�MI��څ�Y���O )ⷈۗ�Y�&ir-4�ݝ:�l�{�|��{DT�q|c5Y1�i�V�q/>�����ռ��|=u��y���9�A��"\S㙒�Ni`�k�+�fo��mα�a��ݱ��6}�Fx�T�gh2�KH}�,~ֱ��>g��<��g�c��P?Q]W�2�4pT0��f�2�� ڏ�|�	�����
-},�ӫۖӇ��_{�kz�&��j��������|��ra�R�s(�t�1�[�a����M�x>��=�H����nC�nF�������FZ�=�N���K����}tx+nѤ����Z"uS��&��$����.�]D�xft\,���`�����;��F'�k���Mm��[+�ZOnϬ��,&4d�� �����1J�@��l3�ӷ�m����&7����!c��3v�y�͊1�B��`���52��}��"��H.����y��I���oܑ{�t���E�m{=9���zI�yUw�
�ٍ�掓�%buz��8\F��d�a��#MN�u��l�чR���PQT���E��㠱���n�%�oC@2"�V�]<���H���(��^�g��������A���u�4ku�:q�Aߖ���߈YL��w�{�۠w� �ê���$�h9��mF��<3}�)�7�]�@���Z6�CMB!��v�5O��t���q
�	�;Ϳ������oݳ�?�Y��Ԛ���c����q�B�r~�mZ����bb�Z�=B��Y.j�l� /|�w��7���i��͞�h6p}�f�!
Β��E�J�2.AK^^�BQ�|$(��I���d����H;
��?
�c��̜^��2"ިR��gܣϳV����y���