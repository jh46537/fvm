��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $Wժ��Lg�7!	����I 쀸f5=���#��gF������B�Ѹ�*U�i��q�k�ʰ����+
���
W��F�y6å���x�Wv���n�h�3�x^�N���e��&�ٌ��E4�
��%�1.�����cv�J��G� =�>�l��e�	cUB���N��-���oE��W]KJ�쏸��������i�J劂�j	Kk�b�q8��Ea�����W
�4�>��˱��o�f-�0�����=�A�Dkd}G�Dp2߹؟̘�G�t�X��e����!D'F�}��ʭ�5[(�ܗ�1�˙��3~���{`���J��%s��Mx�$�x��\ <z�ٴ�f4��rLwL��q�m�'Gx@�hӸ:���SǷ�&��Rb��D�r���Ao���K�ݞ
qR�*q	�5��L���qq{�N�U7dqIq�) i��9�P�W�p$�`���Q���z�AG�?�jk�^�\�1�_�K,��%���u���C��G2���`Vep��d\�(f��7�5����$�~��_i�Q�[ E�I����D�(J�	�wg��J(%�'=I?Z�j�����gލI&���L6M}��e+�э�� �{Dg)K�_��?lXK/�@!2+�����#\�>WY��)[z������b(�]��-��r5
�p�l>L8���ﶷ�q{EN�aiuz�I1�/6o�M��[~���=�kdlp�=8�<�#��+i7lQ�Tk"�h�����@tT����Wm�FM?�HN(<��=���^ ��Wh��C�K�rj�����?��@o�`·a�Ea�1�qa�PPj��@6��@�%��S�<�w���0�p��61�oc����Xs3{��R�㴽8�,\lE�"��K���B�"��hP��g��H�gWJ�݅?2gZ��0�V�Z�M|P0�u)o��	Y���n�����{��FaW��F���I�!���OFg�e�i�k�i�1���G�_@��5��f���������K�{�����]��ҡ[�[��Q���a=Y!%ݒ��LH�lAj/6��,'���%;!�P�Ҿ:&碂P���@���FJ��.��jic�&�#o��Hwv��`�!)d�e������忸��YF�0 	^��׃NQ	�����!F	������T� ���/&&!��K�eѷ�G���AyW�X>>vU�����2f��8���d��EU����OZ�Y3��fh{j�-��9���=��j�z�ƭ;���=�ס�����ކ�zĺ�v���#�ނa��U�[��������I��l)ʌ.je[�����������㢖Zڷր�>R���\�=�he��Z��>� ��@���z��@3����[���*�k�