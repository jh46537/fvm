��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��1�z��(����Oe;����b��
Z=צ_|���e�Œ|bŋK�G�{�M��u� �o.#����ӯY�7�Y��g	��_������d'0�k���aȸo�O��} ��y�kɛ�n��|��9�{��о���>�<~`�����J5 ��C�G����Z��-Ƀ�1��'�؎R5��GDaD�6����5�uH9v,+��j�߉���dE�`T���n�\�ju׎T�c���L�q1U��G�q1^j��Ճh�o��f5r.Y�ϭ�^��܃3�R�d��b����*%���!Bktp����B
8��ÊElO@�N������'������V-w��
 5-��d41�S/�U@�7��#�l�(������8��c�yZ��n�n�R�p�x�Z���q1w}`��HʨyQL^�h	W��vh`���Z�^V!J�U�[�N�☽�փ�"	R	ٌ������!Лc���'d���R8�_�;�T�0��~c
�'1G������@]�D<��N.�Z�S,�G}��.ٙ)�M�(#�3�[�=P9#
Z7�dSþw��9�Mʖ�+4�=Q��,ƒ_�Y0.��/%�4��\M>��dz���Jr^� Լ�p!����ĎXe;�И����3����W��\޳��/���w���������4�wQT�&��Y(Z�?s���}w5K3[28���}�|H��xd)�޴��u�߰�8���;/���.p�a����kI�wLظ�n~f��X�m�z�T��@��`X�F_�A����8��	�A�e�E�	Oܷ��ۉ���XY��8Ϙ.�D���uT@��#;�	2�ŸkQ�9�9�נ���XgI7$��w�%�P�����Z{��*��E��� ]3�¿Vx�Z��8Z���OG;�!jי��(uYY���Hq�EХE4�du=Gptj�.W淋��y_����r��,L�FEޯ���h�>�frp��W�{�k��e��L��g^O4&��D�������`Bޏh��T0��S�5���6Z%[�g=�֛UH$_H�� ��҂2�CA %�}�+��P1��q'�3^�m�Xg���p�s1�^���ݟb�3��ma��%���a�s�t_.������>2�CzCW�$h��������O���9�\���ހ���G���h�!l���T8n�U����^�(�,7�%��ؖ�}����X����'�l���rN��
�H� %��+Ѝ/2k�;\���K�Jvc�zN����`�D�LJ<z�7��)#���!��ӓ�p�y"��R'�|�gn^�-��	�0�t�����:�]���r�:8�<��c$�vq�L������2''��+��+��5��ǐ�xT٤�?�m�t=�dk5e ��PF�RͿ�*���>�o���)Hmɉ�'CU�X|�Q�����G�)���s��rq.M�"��p��w��>(�����+���B��6=v&)\7���q_��ߔb�r���s���C;yY:Ƽa�3��KE(Q,J�֠�b�N�pÚ�1�l)��͔�HC�u-�bv*�����	�<hr(B0��ڒ4����Xl��J�������1X/z4vi(.���}�PK�M��������+Ԭ�Huڬ�����f�vj`����� ���ߐ�uE��Tx2�gD|�o[�ϣބ�	(�g+�7��B��M�����G0� M{���Ik�8%�=�J���Oi2�r�7���8�q��r���b�iVF/2�X��M�B�L,F��Po^xZ"���!��D�cT ��z����r�A�u�>R��_ߜ\���nB�pM���+A�Y��EJꯒ�2��7�x.�o=�vc��G�%�-LVЭ�����~�}Q��J��i�ʴ����}D0|Иg~���yYe)������t�Q�X�ڤJ�`������_!(&�HP�����.�c5��q�6$=/**[�'��{?��zxg�N�m2��*j��fSv?Gc��1u��?L����p[Y�����V�rD���ǋyzj�4f��Fn�J?0Q��i��}�Rjk�u�]T\�r*��\zL���2��o�BWm���uZo��C,��>P�*�0���F;{�يȈ\�h혽�! ���O��4�hV��C m@b&�i��A���[׹�h�J���ư���ǎJ���?�d̛/쨵b^u���O=�ǂ"|.U��w2����N���J�p����/����=$䩶қ��j�.)���f�E'�ga_ r��e��#5����pO?�tw#;sT��o�v���O�:9���՛�^�,����6b���=���@�
1d1�՛��`�} lA���%ؖb rms�5Q�s�\F%'��Z����׫b�l����.<S��
�� o�{c^���.x�/�Ž�C^� _��͔s��3�FR������ ˮu�V���'}	�[����.�LC�Ti��������"�dPcN�F�3Q��� ����w�_��S8�
�14XA/(z@v���Yë��P�H��]|�l�U,�����54�;����V����j}�`��k�~Nm��3E�[z����~z��L�P\v���ն�{l��"R,<�z�'\�+�sPA|���1�Ε����������R/pvHLn���c ��l�-Ri�7$�+���i1J��
�	-mr-@F �C� �W�����UvL΀,8E��N������ܙ��F�֫	6�fL�s�� �
���q��O?e\2��u�N��d!������O��dM,�����n9�a��;=Ww^��,�𗏕�qj,�:/M�0̷"��w�J[���Wi�sֆ�B/`gI�ؽ��+�/��7�;���R�5�^JHy}�֭9��J��*����y�r��>g� *�I,�[��9��Xkp]�{�*���^��T� N�p=]�<�̿��k����Y���ĭ��i;�h��
���D�\S�A~@ߠ:!���pЄ`K$��a�]Ui���E���/�՗-�VO�g��&�;�� ��u�SF)1�-(�O�틠&�2������+,��)s��9���x
7|K����s�bT�r����qx��)�ۻ5NOc�äU�����Q�2�&�C܉*��C�2��C�(�`kA�e}�����A��Y���Ge�}�e���t�<�5�y�3f�ɞw���Ӈ���h^���΂n�������h�Һ�j~*�$Ba�4���:����Zy�f���{}��M�