��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&*���α�&֪_�ս$��C.����������=�-W�#���^�n�$��
3���o��ͩ��N>�t[���@!��U.�f
���^�Iء���P�dʿHxK�K$�V���m/b�_�a�����f�\ħ{���U�zJ��N��v��M׷����]V(E奨�g��`���P��6��n!"5���B��$��(&t�K��8d�P4&��pRB�J;����|���<��"m��Mu���mVS��<����)�,����s��E��#{��b��~�B`/�u$�go+�3�PB�083f������z�HΪ���L��kB��A�: R��l��fA��*ZXy�o1�o#��7<˶pb�
~�*7L���
^x������I^zf�#5� E���N]��Vb2V���ӻ��v�K�Uv/^��\J�-��V|��v��ǻ<-� �#aPG�{K���3j���T{�^a2�;�C	��د��ޔ>	�7��,�]���Ϛ�N�=�RS���ʭ�.&���ST��=���k��68@qˉ"n����G.$�,٭~���2���˹ >zI�Z��_"��{x��Kף� SI3�d���u��8X�ޫ��r~F�G(�=��VۗjR9�Ӭ+c���(1b���{x��!^�a�;��7�)ZK9���|T��_��v��w��w�䬄d 1�\�,83�A��b�̜(�%9���a��&��@�䐈��4��������w������#1S�M��$�i7;m�M\v�h�#zr�Բ+>n����ƯOey����tE�$}��� �&�!h�ֵ��a��'�L�v��`��:Tb=S��B���'��ڲ���q���Y� ���^�nh��آh�E���9\�H1��s`3���yS�AI�jr>����Jg� �7�>流e$��:�Q�{��*�%��F�l��
�%�����`}�@}D�p��^�p��$�\��7m.[��k�#���iG��/%z��_~��0bʔ�lʻ'��U&�^��vN6�H�:�u\�ŸV�_�Aܟ�3,*�Z���*Cg<�wUV�z��H��v�Icz.�-$I�ojw�:ٴ3���e. w!��F<"W2�_A��)OCa�� ��B�a*[Nǚa+^U��py��0�}u�q��:bsD��ᯡ�vgdIl�
�P�GߏK�?-���U��yIe!�`j ��iشk��M�I��m������l�|z�{����f�,
�ʨ�Q���(��GOE���D����B�PÚ��z/Q`"��#l��Mi(�oA�eV�RW���~W�~Dp��t���zf�L�Z�8٫_�DzZېE�A�;����Cf�;Pχ���ԇ����44����p�&�@aK6�h9 �jo�F}�.��6����=��{Z�M ���Q�����0L�L�,3�k �\�]�ezR	ݑDJI��Rq�(v���K,|� ff�@��b� Z�{�R�t��:SU�\[W������;�?�~�ۆ�>Of��<˙<��Q��Rr1%M�y�m�M����߈��i���x)��E�W�_��@:�~��J��I��4�)Ha�@-�&����d�KYm1ؔ]�`�#�i�h���y���n��7�pփ��jZ����\O�$��Qyi�gd�r��9j�,$��ѡ���ߖqy��1_����e�R�M�W|3�0�a�f� N��NU�E)�\���,��f��]O�'}���oi`���<#QKU+�+T�d|�\{;����pu+=t':�4k�Y��т�.t8GF�9��Ӻ�d��G�e��8��F���ʶ��x�cSČ��?y���G�Dcy�r�+c/4��<$H��7���ʎ'�q8��G/��-ݍH�����d�f ��7�p]�x?l�ژ1�!أ�)ϭ��2��I���D*���J7zюmz@��F���{J����A�z�]�$�wɛ�H�����p�-��� �^��O^��3$S/�j�M5S����v��.��.5��T��2>%��[�7i4�ג���P:��!��/4kwI��f�Ku~�edDE@,�u�XwsX_c&Ak��Pm�+��,�ړ��ܵ�⇎ܢ�����la��oR���A�y�A#ʇKj�h��V��U}�V�6��'������k_V�9�����%��_�S	�/cbku�Q}hG�q�(S2ڎa�L��"޾�BX���X[�!�b=ҷ��{:����b��s�qBH���	����>�x��������/�> �$�USH(ᩄY��0��9�����@%� ��6Q�W�g�y�dD��_�����Y�&'C~~��g$�^��9�_fJl��#���w�.��5Н�F���Y�}&����qg�]E�����a��/�@��v��B�/���ܒG\�)��{�~��5�P:n���b�(����Nq���S�-u���O���4�N;K���\Q&�8o4�ǃ	�?�Tf?�++�T����G�_�T�?>c#�؜��[
At ;}��f̙�ep+��������t��Sv:���<�����>m@��:�*�:����C��B���h���Km�V��u{� Ae{G����4C�����N�P��1��Ԋ$r�QB�M���B�Mw�ʶ��=������9C��*�!�S�~"p�@�~k3�՞�j�� ���*�`�D"�T0�����ܮW�]�E�Aqhbq�>��QS�+��k����|2Y��!