��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�ֶ�3�4q����}��{x~�� s{��TFҫ��J�^���n�AH��k���s��#_�;�b�O�u�|�������֨��#�:�b�\77���}T�I���kX�ի@�6���12()�|{J�4�&"�}M3���_���mD�ی�`[�K1=%"�T�3����j�;&���%l�`��:��zAjG�����.{��X%Q�Ͳ|)�K=N|�lw���XP�4�@]��D�����2b��"u��eg���J�u�%�4�^��2V|�]j^���
,�9�O�1�`.�2B��9��5?r��7����։rmf��퍱��CP�m]��}���&Cw9Z]����u0J UO��t�i����i�O۱/g��@iJ���2[�LC�(�$sZƌ i�jw�ҡ���[�c�"�Qjw�cK�َ.�$�]ɒ�\N{?��/|����NB}o]O���G�߄PUS�L�����$Y�!�NXΙ�mA޻���'sZv.'Ɵ�#%|R��Ey'4���ꤹ�|Pr)8�3���Z�9���.��]���+�\�?�zX�P�lg��feY�^�Kb��a	D��C{�b�}���}I'�x@!����v�-�-vuL�$�\�+�?XH�M��ÆN7����:�~��l��T3�Z��S����l))�#�yT�,HsAFi7����0�F�$W����HF��͓��c�={J�ʯ�w�����w��c.x�=��#��ay����^1Q
ڳ�O��,�/uV@��&a(��a���F_���ɏ*�_�|u߃r�c*a�.�*�B�tǨ���rk5�d���(�*�G��y�@�"��zB�\>PY�A <,�`���P��^�I����I��,�b���D�	O��	�I�N�R�"F�����,�0А�������߀5v�5�\3��I�-h�͡a*`?[��dP��=
�%��S���X�����V��z-aL�r�_�g,.�&��ƨy`�u�Ld�� ����x��2nz��%�q�z�B2�����C�� T�肟����w�A	�9����<�jb��@$�N,�r��Y"`�N �&��N�XUn���l������@�aI_Ouz���<2z$֐'5�K.�I�)��nv�z������C�a��ĳ#J�'���I5�A�E��_X��?.��Ǫ���EE�X3`�]߰A҅�ǫ����}��0j���0��|;ˬ�
َa\�89jøk�����D�)1J�3��������@�}��i}jy4�j��ץb�9ā�{��W�=��M)���t/m�t=�/)>��Ƨ�;����4b3Oè�F��&�	ؚUR���mw��Q�QPd}�5%�5;]��'s�͊ ��;"����Zp��w��U�b��eH�k5�����~����"�����O-yF�4(��.~y���ҽ�ܖ�pv�@�7�i�6��n�"��pi���y|ǻ����(ߪ09��R�,��䈝n�
�k�,�$i]DVWM�ѧ��>mb�҃Ҡ̿d-E��p�!���dA�j�^iҕ��	`G1X� ���n4�/��Yv��Q�G��&e[n'%� VRvf��^���1�]Qq�;d38�+V�n+�Hp��Qg�Z���������������Xsv����*�[�-�O�����*���ؤ�Eܗ!��<Ԅ�zu�f� v��6�~g�v��|��e�R���m^��m�{15lIJ�7%��йx�;��w����B>�ِ���"�i���9[�\{ݓ�V��������>�g/�ؠ\���M؁U����w60?s[�y_4�{c��?t�@��o�	�A���Ws .���xg�D��*��t���R����o8+4�a9r�:9񮳠�N��xqzQ��Ԭ��Zf��e݅Z����pW��nD�{�I����7�D��4�n��\��Xv��W�w�.QBq���]�a`H";-��	¹�y���(T�j�����ھ`���Q�&���
��8>_���� �������,� q��I����j�> j�����v��1�i���̷������}��-�+3����x1������"�I��U<K^��v��*cQ����E�+���	�w����h��<����A��>u����I��6+��$�dA��:���o��~��B)�N�����p����&U�ϙ`�}�'�{&U�I}� ��n���{*����-�a�����/H�VQ��
�~�OQp�Ų%�z�ܲ� b�~�_��������B��x�����	�_�b��ߍƥ�w&���΄A,��_^�d������~`,�)�C͚*FN��t�^F��Ձ��Y`'��M"����a���pxK����@D�EPء��7!��&P�`:Ӎ��'�=4�/x�7��,��
/�!�bp^Q�:R<vz~�o���dr���M��v_e�SR�F�@�M7������s�#z3\�V7���^�&�[��	�$a�Ǒ�y�$�g������ ��n�2pe\��%�,7��Y����pie�2�=�1��w�i�x� yy[��=&��_L2Y�
k��	]��SA�Rp������O��p]h  H�Ԣq�φ°H_�r���� ���B��iN��w�o7�(o��w��[y^ㄷP�n����
(�_#�٣
Uc�E>-�ܲ1��r�H>@�ת�~�-:�4OA�k�u���?Z�<1jMW?��d�O�n�؇��K;��J�T9JG����	"����PZ��d�)���C[6��s�����T&3@h�Z-\�A��FLR<�0A�+/�֖��'�cWi�e3�S��S%�vo9�)���,�i#���U&9�H?�2��>�*E�F2n��mZ�����?�h��{j�6��ۻ��1�jN��[��fV�B$rl����i��5�\7�|���r��f�
��i�$�[1��,��ÿ�|�)�x){�|��_�Er�p��qj��e�QE�f �
M��$]��;U)�-�i�N̅��rcϞ�����Oy:�_���cce�kf)��ԕ�PO�/ѻ&����Ӕi:~(V�".�"o��mSD�XkD����o���)zh���0�UL��_4s�����ǔ��R
,;��4�$7���k�.�v\ȂL��bN|
亅��K�to���I�a�@�y����"E7S�7�?׆u�u�E�E(�Ji;LC�1��朮�Ϻ{\��<_�h̃W�a֭Q��,�������8��s@�_Y�p4vM�z6 ��Wܰ��������\�Ҙ܃	ɪ�#�P��y*�U�wb5Be��.:�
҅��Ia�<q�X�S��J�d;��T���S�>٥Ρ���L�(z ������ɯ���=�����}P�ym~�F�v����^lo7/	��y��.���͔Y��r����o�\|NB�VA3~�D$�p��;�<��ު׷��d��%Zr��X��++�X���4�1��a<�Y��c��Be�ǱT�ϱejws�f��S'�٩+0��&��/�"�i�Ob	�j����b�3u,��t0�=ʯrގ�2�R��(2q����uw����=yw���c#� �,a���[������w�0RC0�LA~d��?�y(S�춀��<���2- ñi���ȇ��CEw��9.*{bN_�S9�v�q}%��L��h���o%ol�$=oa�S��'�B�� ?@���qk�%t���Z���^�&&�$E/J��=��y�C
j~��TFՌ`#q�����!�*��� ��p:!�vhqxA�����w�:|��(�=q
��A�GV`iB���(��; �{�i玖̈�*�*ˈ�%S[�u���h��٭�J�7��[��e
8�b�����.�dֹ ��m2���t�A�i�L,�M9PP�*>�>�n�3M�­#�����Փ{��@�P-y�<�Fs�B��ՙၱ"��7;�-[ ��i"���k�\����Zn���@�i��iP��D )�
I{N.{��b�U�=,�!{�%n�ϷW��f��^$6�Ը;0����z�J�8���^T�9*�����t�����u������@�sB.�[�\*^2Cu!*��0�a�꤃�Ѡs��^�+0齋�R�3Gi���ռ��D����sٝa"A�:��s�;��P ﵮ�Fb ��d�{) W�Ã̛p��uU��/ņd�J������(����zzZvv܄(�wf���E��ǆ.<��<��B�7Nw��.�"ye\E���c�X(�ۍ!̖TF^�>
����F�"R����'��GG��z�7����{1 ق��^�;p�A M'W ��`k��SD]�����zC�$���[�	@cw�^��a��+a�9�C��������gP��g�};v(ͩ�R�t��3L�y)ӝ�lܓ�_�FEo�)V����0���f��ag-�s�)��llƽv�eA��ٶ�0R����ȹ��C��aM8\�1/��;7B��ٍO;Q䦷���pĢ[Fp3p����-N�+U@T��-@Hp70��a��>r��
�Rk�	� _���� y5N%\�AJ��v鹺�����D�k�!�3�-�vI�U�?��,ξ_�q�ҵ]�9��!u
:9�&'�J�S�7%mHu�P s�-��t~3D��Z/��U-�c* ����6kW��8�s�wa��á8Tx�u�	�z�qJ��j��w[�p�5|���%�-}�ܹ�ޏE�M$�89>�4�T=:��\��b���v��O��p$��l|~A�G�,�Nsi�&��q��o��1�?�Qܭ�J�B��p�*�[j09�g�6���T6+90/�G�'ft�9�]��L��w�w��'a;��T�5u�7P?8�+���+YZ�����$�>uG7'�^F�J�p�v�j�>��w���3e�d�ەeq�P9��RA:��c����e��a�9�^X[���-xA0ݹA�bW=1ڲI���2�,^�u���n�+G%_�kYb+v8{!>-j
���/O�َ*,щ�(_Щ��3D��پ"�uo�/=�\�3DW9.��AI���h|!�k���lȞ��8�b�g~��|,��3�J���tP�s6�驭�쇎C�z�dݺ[�n@\���N��}�D(<S N��*u͢���!��!�&#��/�Ѣ�Z�CF|;J,g?�,�5@���feZ�s��Er"*_��ѩJ�t1�5�SF�<����5+3)��֠u���@jDB�*�!�	M"fυ�ӕj�7��DOX"�D� }��8��c����F�����/2�P)�/�V�?-���F�:^w��ԕ���b�F�ʵ]�'c��
�;vN߁0��B��\�Ek�C衑�YG�z��-�L:�ߍu[3|3@k���8�?*���?�z~�<0��J�^B�짌��w[�1���X�j�#��V���!'��s�{V��u\�Xq��"��U�� �	�CD�k���CE���9B'dUs��9���y���~3�����o]"!4�=F`��<�I"_�&��qO![�t�z}c�?�{�4@D�	&�IvP�m��9�o�9����`�ZӋPY0"�����8���K�XAo�����S'�9DG�I��� ���"v>��#�{8?��8Ƨ��r�C���ߴ��z`�y!H�?,�F�������5`l��9�T�v�M�.�nL{m~���`��	�۪ �9l�RU�"�@�/s=����qu�{[���r�Mf�K�Tحc���2blӛ�p�ye�S^;�d���S�
�-�D�ΓhX�&�� �2�pfqJ�e������t/�]F�35�kTW4:">鿱���$�N�iP�v�aݺ^}��	��+}o�����9�YK)%�F��d�Y�5�������fx�q��vy{ǷKt��MO_�ˎWw5�%/�h�� �<�D>�2&�T>�M�B'�=@�ro?�E^1�R?Ҳ�O�B�"�)X�d���+��]�Q]�E8��{�%2"�����t}\�ד�B�!'�2+j��p���x5��#�y* .�Wf��>�6ð�o�[4έb��)�~����ͅz�AD�P��l�7G���8��������a&�n��!��M^��
�!��<I����Q����{&W-���v��"�@-bڰ�2�1;+|�>�� "�Uj>5B-� g<�O��~�M�WIS�^m��cf�'b9F/��HT��.3�+�"Zpsiy��6W�b�|��Q��ut뜼%7�l �;؏b髊�}��S@�XG:��2"�N�zn�o��Z/d��e��+ž�ǣ> NY�!�1:�$��:(��+����z<Da�\m���N!����)�[}�$䦪���1�q5+$���y6#�u�O��u�vu.�ř�.I�]#P���Hr��ϭ��lw�4Tzӱ��N�#�ܳ�1�����Dm�����Ԇ����M�zʽS�?���2c�<�����p��E?v)����>�Z��֕=���Ա (olt�w�&b�����tP�[��b��ρ�}l��a;6(n����Š�g��Z���kû`�=����p�,��&>(��$7��V%?=
�ۡ�y_�n�M����/�2�r�b$���Q���+��[�g��:?h�P@� &���ĸqJ��
����k��]�b�xe��F�zJƣ6u�uQ��KD��g�U?�f��t��+Q�!���S������Y��63 ��C��	*�pf�ZH���]�-7jS���~�5�t��n􌒇%�r��P&��6�۲���J��P8�.Lhi_��C�n|N]�jS~��D��a" ��l�#,�א��9ZCϠK��ޤ!���y��3}y���﭅�P9��W��B�̵�蕆N�l��5�kyV���uDyt!(m�ǥH4�&�2�U[^��v��r�B���^�BL�z|�	>6QDjd9�n�W<�^#P�E
0j:��~�/��?b���\����u��-��SZ#���LtyL�i��:�Q:EX�q��?=��4մS�E������ܿ�ڋs� ����H����/������4
6�Ei��w��Dٲ;{��<W�2����\�Q	��������盱��عp�0id3�̅�~ʹ#�!r*�0}EQ����kd�%���{K]#��R^�6����d�7o�����ڻbl�SF�@���ur
�����/�?;�jW���5ė$<H��.�ԾkKU�O�4��"=��JD� �С��v���Y`}-Ub)SՂ�O�[�{�~�\̢S��;@Ҫ��t���)7��h(7kp����E�EIqO$�$A�|VF�p���AD���n�II���Q^!��z��K�\C�K$���#�sD,�~�q�6H|A����L����!.YL^O�7*6gȒ��DC�b$7`�����f.Cf*�մ7v�p;i`)����Q�r��Fy��L�|)Za�UyR�l�MmGLã�6��M���vF�r[Z<�%�k�p��EP{O#U�K}.j��{ts��)m!ƅKM4�.*7U*�t%�0S�_,43�`���M�&&IE5�2�{���Ҍfp���s^��Sr)�c�k=� �m�B�߾:� �S���Ѿ&^��f�^+�.��!�OT�^��L�����:;ym�Њ�zc�(!T�x&�3RBe�Ԋ	�����b32c^��h>�jI�ˇ�I#	��)�tB�F9x���k�@���|vbE�_�$�w�#���q1�h {t|��U9�=_�S� ���S��̀��T�aR�:���Au�I��N~�`�a]�6�Q��ݞB�_���1IdX���Tet��N�YY��b�Ѓ�ssd���w����>�|v�ןv�� ��@p� �(j��@��X<�%���D��9���e�O�(�����������I���ʙQY��{��+�YT��9�]>� e�w�m~:���8입�Z��|�Y�yY.��)�>	=�=�u���Ҭ�<�Ӎ O��VO����Cu��c�C�a��4�S�[$�0��������E�O�YR���-�nONw]hAw!�Y�N_�� �6�*�<"1��d��\�2P�����;*��p5����i<wq��`�li�tT@>��do��:��q�7'�<�*�N K�d���.�E����/���-�
&���=p�)��;��
�b�(q[)a�[�wS���B��*O�G��"{�\,�*Ǧ���!٪7���Z�eؚ�:�R�֮�{&���$⥊+'�덃�Ek ��E�z����j��o�� o���B��Y���@p�f� r+�^��-��V1 mNKՃ�n�&u{���N�W(��B#��+^�-���p���6�7���O���X���0>��:�4��/Jiu}�4�q�0�������}���񸏮$Sֻ������/q�2��ฐS�-�!�5+#��vFzA#�w��H�⺣w7��tI�/�b@A]�8�-�px�_���KR�.�����2v3S|���ec���ř���CV�?bC�viY�{qQ�vf��"�|�ұ�-�����k�@��)]����D���`RԏE0m>_DF�}6$����8����1P�+ϡ*
!�]鳃�h?b��n�>t9
O#*�4���L�1~��<�53���:���ک#]���{"�LV��I!�j��22#�
2��"ǋ�(m��f��EKMx����k����I�+��2?��v�ېU�+���l�B�+�Xf})��֍�zh N�R���ㅆ��-}T.�<�4�(�#lU^�?щ5��u[���� ����y�Z�cy��T����GOua��麛l��#g3�sn#~���G��t���=˪v�̣6�JD����r���n����9uP�� ���2W��9��}���.���_
�7�@�������ʧ�o���}���_`� ]B�E4r��Օ��%3t�r�WB�kX0UN���sM�a$v=q��])�b�=O'_P�F:X�D�����i��6Z�Yk�(��LV�Y?����{O{|,fH	`qw�f$�M�>q���4�hU��/Y6�����fmЈ�����|�܌H��x<6�]�^��% �e��"?��y^J��� �ߙ�C��������C�f9ES�X�Y��6y�`<�� �[�[o���s�5\x��˳YL3�B�n@#�¶6�-���G�-9��<_sZ]	��G�n��eK2:J3��� ��n���	o\2zΏa�;���a�TE7�m�`�R�]e��c��~�l������n���K�cF�V�A?.�QR2_?�H����L����[6����T+���ؤD�Lw����U�,�P���%�%�`��&��;�kt�813 �^,����g�I��5��yE�K�HMo�t�\ޗ�H���|�q�2��[W�z�A6H�4��r�1E@@�e�;����v�$P	[%}��������f�Ϲ(!�̢,�����ʙ�r��o��ε�3s8�#c�WT�Z>a��^�hN	0����\k?�'J��^�=;*"�,�q�'�^W$f��9�=����I&A�)-��^�Q�0=�Sk!��_	�g����H1��6����;����e�� ��:��,�*-��O�a�6 mY^��"#��9�F�5A���O��x�h��)����?����G/9�9���gͳ�~K��}�noU��K���#����"���?��ˢE`�6�I���`&�o��?��"�Uf�"�KX��p�����aJ��nC<��E���"T�����&�8r?R��7�!L4#�	s� �N���Fa�%W��c�<�ie)� L��>벢D��I�w�Q��1q�RٍZ'r8a���7(���A@��qʑLc�+T:�Cߖ�g����O�r�i�D�\�C�T�hQ-���a5���D�Uc$!>̗��2�%�k ]�T�ֲ���թpY:&�g�"��z�*KHӣ̽}5UNUzW)��1�������9d�b����#`���pq�h�˾wG��=,�\I©D�-'��BmAR>*_�}ؙ���cT������eI�f�N�ܫ��w����5Rc�9�����Ɋ0���������,,��J����y:��9߲���Ci+1�߱X`Hs����z=`#�ڐ޸NH�l��M��$����5	 h�ߐ��*�gR���:�����9՞��
�2� B�FZ��=5�tI2�k�c|������ݛ�i9����l�3v�go�d�
�[���e�G�~O��^���^���J�������鿫��*M(������͟p��J�l�[�*_%˫C���)Źa�ciY.D�}K	Ga&�cz�z�1%C��*�1�G���5L
#Dp�!s��qa���ڀ����"z4ٞZ6�0���Nk�)&Ɏ94���Պ0`1������t�-�?�om�ʃ��hT�Q�'N��/B2xh�_oc�r�����u��s�90[r=ė&aSF<x*�/�Mo��?)��h�9�T/��v����8`*��р<!Î�FB:2�(����
S�w�y<�-@C�F�0:�U��z�AĂ�cf�*�:S�D�_y��Kcj�iW�B���i�ŵ�t>�m6aț�:�ϕ�af�a�%EwwM��U���rZ�P�[��̫
G��d����M��P�����D3�x�Ȕ{ؼ&�wF4�y�����ԏ�˅D�'�q"diKc�o�Cշ,�?p�"#�����eXHkcj �i��
�{H@���nG�Hl�ũ��a?�e%ԣ��Zv�Ԧ��ޙ�#��`�Vg&`�����:PA�|�D���}/���|1�jXAw� ��d�=.W5�<�ܨ�3b�W�v�,�]D��ʢ&uQ��YPB����5�W|��[�;Ӥ�H`��r�lI�L��9�G���Zs��蒡�7�p�u���ھ�W�q�G���bE������:�n��d�KӉ�}
Qaڼ�:l�yc���3,�5�8�ۼ���|�(���J`O}p+��+}줔y%�T*���	�\-j��8&��/��ʆk*	<{\��s�V��֓0MR����X�i�es�v�Þ͵0�Mhr<�D��e~!Zh�n�&�z_�S5'=��9k~�8�Evǰ���Ib��qjJ޶2��l�u��ͬ�6���'b�Rq�Ϗ�8n�яP�����l�J��>sRc���U��꘺c^�/BM�\��g'�b�u[��LD�D������k�8㢲f�>�@�A�d%�	c|�wm��m�{�<a[v#�{�4������Ȅ�m���+CR��>�W��!�|�x�t"�8D���j�4!�F����r�`N{��;�چ���M�B�f���2��^	�P�R�	��SThC�P��\0�R��C����k��X���M�^�tc|����e��S�8�_N
A��s�h�+n�An�}�?����r���3/�h�Q7�U������G�!��C�:��,a@vךg�Y�x�xRd�2�7��>c�~�$H���Z��6�1,/ګh��!׊'.�z�`�2Ր$������T,�і�9N��<2�E��x�}����/��#�(���x?R����je?vi��اGghoz��W&�U(����Ǹ�j�_f�,�*Y��R��OG��*tn�ϰ"嫾(�D�f�ų%�!���?.�7���F��&�8A�~$�A@�Z!�
h��4��,κYi,�'��^���<�g�B�����+�����}�R=7���\�g��@�#6H[8�D��z}P�l��K���n~c.�)��n睮��^�`kw��&�B�O��)�x6]�5]�K����a\4/C����۸@;��ǐ� Fs��L��|�4*qԫ/e@^:�a��j5e��VnI����;����;��Q��Ȼ*���q?zΊC�*cL$�bSWe����ʑ���MՔN�ԲkL*���U�@0�ƺ�1�U�͞D��Z�ߚY@�"7����6V�x�Z��br` �n8�!����,��8�\IF���	��+X��ߩ2;y�h(q���p��r���d�
7�/F�$�_�׼b���a���Qk',�do�	��IS"z
&����y+��npŔ���Q��D��lMwj����1�,6x�%i��zP�0wQ�s�9�S:b��t�ǐ(��Q�?(WI	��^�ef�o&��ο�=��ft��4��*O��3����Wr�Ww
G�P~��b�5�X�2"b�VR���1�6PC}/D�e��R�.�BJ:�|}c�aO��x�oZ�%w%6x��d*h���mJ������2�7VV=�$zn�)J�2�VT;��P�-�}��jAۚ)��m�_n"���R�?,	�G����3�q�4���J�܌!s�f�
|�g�ˈ�@E���m�*�R< �3�v�� ���`����5P�P j¶w}@��f���Z�r\(�_���6ݟ�G�� +$jO�rQJz�l ��+�HeBk+n���CU0���[T/j�a
ЊI�#]��G~�dܘ�XYJ>ݗ��Ξ;���a@VN��6��N�BR �ҠNZD�/V4?ڷ�2bv�ـň�p��&�
Ćѩ��A�\�7`�i�7�[�mC�ޓ��]�+��(�7��H�OFP�����&K��?`�`�UF�?9���~�S�=����3�DX��%.�c�F�e%#~	��t��F��]�_�VLvJGZ��,�U�L��TvT�#(����uV�}�Y+�9Vވ&�qzюNZ{jʌ�nq�ݲÀ�ޫ�O�bZu�����3|��<���lճ��Z`�^rU���g�I��u�kz�]zg�]��*x�L蓩#�B�2TS5�f}���U4�<�\[��ϊ<���	��xrym@
�׵`�Tb̶��K؟�O��`)Z1(}�y��ĳeU�eL���>�V:��P#5!u7�����x�B]�oa ���%2�^?`�î�@�䆾5q7����E���?*A+9`���L�d��2A'^�u�R�E���^�c�'Fט�!ʕ���Zl����/ _Ը0���_������֤m�<�V=�v�c0nԕt\�L�)�Ʊ��Ni���.��o�}�a�=rs�5Ȋ?#���A<�c� �-;.�V�Q�j-/�k���Yu�G���EI=��	��9�q�����'�����l����]��K�Ŧ�{�xdZ����?#,5�h+�(N���ӹ�Uxo�g�[<g9��f&c�ї4�Q[�`��Zb�7���>4�_ßd޾��I�׏l��S_VS5��K�^k���������9"�x3��������d����5D2���(��h����gF�J���kZ7���^X�/��������ؐ�,���0�S ��w$�*�����^k��V=ܞسt��ԅF��*��X
u���0ZM�`m_�O#x�$����멜�0�sčR1�7�`C�qH�ْ�vD�N�D��k SV>���9tMw����-���ф��D�Q�T�����#�6�����0��MQ3u{*�_D�N�:�p�.�I���`���;_�<o��y� "��<T��N3�gWO����0�IR��3�@Xdo����ҋ��vP���e�[�A���S��b"���g�i��lư=��&/�l�� �#�vΎ�f#��.5��}ȩܯ)����F���>I��\~�z�:�"�@��\����7�
hh�$t՞�6����T�%lЂ�D�K � $1��G����e+���';z��3@�M�l���G\)gAy�}��"�6���O}��{`���?�{��%K!��[Қ��?��dO�\��9AÍ�q����cy#��Φ�䐕k��?#�n_,��O��d�ɄA�U:ƻ���h �,�R�L?\�{p�,rqdB?�G.Q�t�$x�$������T'��h�����D^?��r��3��Bܹ0�[���H-��ܛ	�ۛ����j�=R��L�2��P�_���D��� ��4%�)nM�`�'�rZ������z{=Sy�b�&o��r�ˑ;	VUUM���ԑ���w(�q)�X��̬��=D�t�	�Fw��oǓ�.����q�7ݣ�%��s+��*Z�Sw�=���pXun�
��VN��d��*�ߋ��bD�{f���>��W���	�4-�4Ǟ!��.�A�Bi��=6�y���h#�<�y
j�@[��?�m��m��EEC7}�e>�n�'�@G[��%(a��_�v(�Y�E�{�)�1���ҝ��^#}[����[�7����,aa.?�/.r�����,+SĖ懤�3����#�Ӭ�a�}+�>�W[lO�;��-R�̷C�H�(��9�˯kg��Ǹ��6�3�7��-_c=�-y[��h݊��$OR�Q��ؾ��-�� EM�-�hdr�;'_ad�%^��h'�����S-�8EYʥ+�C�1\#h��3���m�Ә�wC�q�G#}����=G1!�z�2 ��,7Tx3'���\n��U��ɱ@k�%�����.�GC�rA�/�8Q胪/I���ڔ���@��1�FI�9r�%�����s�M�����1��K�pWc,�J�=��Z����@H��3
`e�m���iHW�Y��kj"���6��ߢh�M�͟O_�;�m�G��M�J�����Do�J�:!��Z�������
/�T�L}0&x�8�8r�Y(L���1�����e%�QT@٘���լ1�[�$���D�
�ވ�'H�8�,��',�
huP�5{���������Qi;ҥ)��q<��n����>��Y���9Y+K\f��Z����+�f{(�Y/�Í����Pկ���0��q�Cs"Ē�r�AmZO�X�kE[ı������s��ϼ�wJ��C�D����.h���(g�Vbi;f�@�({������Cu�`*��e��nx�W˜>���Hȏ�4�(��w��{����WS���R�P�:���I��A��/��]ݑ$DT6W�J);��vOǥd��a�]�[����~��4^n
��d�6�v2�si�q ��W)���!a�p�m�7t�3�P9Fd���!��BX�(���*#EwG��8U1�4������,�VV��x����R�ʝ��
Ϫ���1��+}G������2X�<�]�#
a�it�y�<-���e��Y~q��f��oXL�4lh��f��g���]�k��~�q7)-9��I���n���9��"�m�m$&�@QF~��x�"��z��b�&���ᴻ)s�*�;�F9
�Wp�I�IpE/���?��2k���� T�3sU����t
A�b��(�L;	T�dT�=�Ӵx�lfqs7�>����A�]5m�1�����_�̐�A֗N��;�L�Q}���|��n8&�]���k?+-�9~Vi���R��*#�Awi��'�ʐpЅ�=mGվ\����h峌�^����}��PK� )�Eo+
���j����qIH�[��8�GR{��K ���e�Q��z~�r��i�ڲ��"b�ֿ?��aU�J ����v�9��P$�ϖ�����fj�F�59,�(�s��e�X��u'�Yi�>�ׅɚ<�2o�����8��Pz�s����!���0��S/��,u��C�ʦ9�?�{����k5�Rv��[��D8���%V��y|��(��0o�{/��,�xIbv:����U�
e��3����V��ڝG��bq������)�N[�z���&O��OSz�M�+G���o��A �������AK�!
`J�F�TR��u>?��ʩ�2G	��2f�� /Ok�wiF	���Q1�û$��C��6 ��
�uب`o���KR8���R��c��v�u�gPk٤�x�MV����8��0 D3g	:�fkK��Ԕ��X<�m�c�-��b�Ö,yO�l�JqY?<���1O"����:���U��PYxk�w ��˳���m�hI����$�aϣ7hx�<]m�}�$Yk��G��s3I�J�1���� ��L��5�����S"ۃ��vU�ހ.2��qd{/ ]�06�6��Q
�%�M���[o�]��1I��'��P�m�#�,,*G�9�?��-NO�o�,%�?��|��jj��]E�J���3�)�d8xNb���:
��Y��b����\�����X~�"��E:�-��B$�?(&9�P�H���-Y�S�0羅�Kep$������O�. ���͈oP�,N/���`>������o����P��@l�G�Ҕ(����2_jqvl(�>�2p�2fe��C�ͩ��^58y�U�g�h$5��1[_n"� 
S���4����X�,�d%��L�
�����ð�/;nq���2�kl�d��|�Z?���A�����M��Np�m��d�	�T�������4�"��q\�Bӆ��]��l>&k����'P�\p5{E�6�.9��T�eW��,Y;����bvĮ��:F��Re��4�p�.�
,�7�W<ck�g����EϘ+'��ET��@�Y ��5�M�h]��^LSMZe�:)���Xw�΁�a�'ߪTU�;�}�'s�x����h�����ҿPL�^�#�i)3����R�R9�`�Ct�߷�#vL�s����*߶1�Q����(o�zՆ@,6B��BB�)�`>��0|��>�X2ý�%ajɠ�k���|e���1�m�g{�I3�!���l�<Gw`Y�`�8i���y��dϬ�E���X\~������x{u�M�� �f�8};���Y�H�����7�I�dkZ7��8z�ϕs�)C��3uo��G]�2�KC��/����<�.��_� w藻�H��ƬT�n�?�����YbC�A���d��k��T/�hxI��p%��*�m�Z���F������[f5.Y�>5���j��CR��)�� 0��rP		��K����K�jVo�����`K)uJK�^D��l��ӕK-.��j�,��&J����ས�#1X��������1z��b�����l�,�\mt����J�c��fgg�p�_�c	���)���k�ݯ_m��i���g�<�Q�kl�]�s��j~�e&I]��N�x�4�+�C|��>ˁ��V�V�p5�j`��k�HNT+]�D�f9 ���D����M�t�3�m^uZ�xN��"_���^�W��p3��,����(g�w*�)���v�K�۩8�Y^��Q�C:��Smkh�?\�/���{����T3�ܙ��`��f�|M����{8�M�[��DH-�i�&�Oߥ�rB�ɪ��m�iץ�B6Խ$)�����ds�^��~�t'Ԩ'3A���;��xCU���[�x�_��JJfW�@ �.�g,^����$�f�z��uvm��p
�v>47k+ܮ���q��m���}V�I��M�z_����U��&��a)�*л&�	�����!���H�*fe{`yu=$2�׃��"���9�z����gɵq=R�o>�I�y=l$T� a��T��n�� .̑l����`�_��a(�GEv$?U.UuA��}��*�a/_�\(�ݥ_�wK�KӨ���`̒�z�e�Q�OL���o��E����t~��S�Op)G͠���}�P�a`ڏ����.�^@��7�j4e"��`G)%6�����?@4;���/��p��zA�{K��덃�H!�0��Ρ&xP�,ÿ�?o?T��Y�D��	��w��q�Y���Z����K���h*JIIо�b8ό���05��#��[c����/��o���ڮ����px��I�������V�ir� �^�Xr�P�j����P.x}2�Tr��z�8�Gq���
�w��`�s_+ �a���tF�b���ɻ+>��ڴfy��;)U��s���Q-"C�y����L˹z�����Dv/�:�}�
�Ri*�ʘ8G�S�^����v��9z��/|�ɾ#k|PaQ��NP��g���Z~L����p���6mB�F���S\�f�6�!]VJ	U�8M��#���[��$c�;��@&F�G�1�Yk�����X��4�p�o�i��{S�T�hU����$ h��a*�պZ� 	�5'�6$�H?͙���[����|�=r�(����h�Ӵu��1Рe+ᯱ��T������8�F�ȤL��f�5�P3���<҈XT)�&G��:��Th�q�izҬf��y��Z-�=��&��?�p�fCP�d�aN�9����_369����,fW$䨇`���n_��c$P�2�P3��f��zy��Xt��߹T���H�����[�;:(�cܞN���놹=3�%<�fb�Cx�H���o�Yq���I���N�dlH�����4'�0�S�x״/�Ò�'$�����|%��C4�N���r�ů�A.��k�4�h�nYP�d%���}��e����&=�Z+��
�	c���E%=�8w�-'��,������!���N��"�*Hr2.��>�|�Ǥsr<��.�'���=Ћ
e���o�K�9��R�K���˂�I�ln{�ýL�5}�����{��E�0"�W	?�3:�c�ur&���=�L�i<����(�ٰv0^������9�0 LY_��̄	i�d�dvaa�e��EQ��JY�Ij��Q�)#�d���w6����\U'6D�C���#<գw4����!��iT�� +�\42��Vqh��)��W�T[D��C�rH���H?�%
#�F4�����"��7\Q�
�#:&��D�w8I������0Ȁas(�AX�x�p����)��6�	F����#Q�����D'`�c9P�%��w�9#ĵ�29��?�|���1��:�'j��Sd(�	'�ڳ���E]��j��|t��9�`dI~�	=�٧��`�Z�M���r�'��^93��_�Ԉ�y���fj5l���`iW&d����q��6l��m@}���K�c0�,.19���鳁7^<������0fI|)���x�@����z��F�y�Fӟ�#�t'`�6c�p+�����|b�8<Ƶ �io+�-ϊڋy�pA���oR��Os�gp7�7�bsR�2�[wB������?d��A���R�-�Ȩ�<�dj	����8����ٻ����k��o��p�"X6v*��=��cݚ?�C�@k0�" ZW^� ��,>���Z���v���A ��F��F�I�v ���g��*bC9N��C�L㰈�J�y�a,���lY���b�-(��}����2,dԤo@r��;��<��:���n>1^$v����Xd��_q�X���#���|ڝv"h�c��B�s�����Re��~g���	�`IuU�Ә�b'��Pv�����8����j������� ��AcwݡأS[�� ��%��g:9c9�����I�%r�1g]�sV�8��>c�3O��|`�~�6�*��u�n�Y !�B�+u�������I����w���is��z�<Kd����LXg�_���IE��[���
0���M��x�֡l'W����������5ɶ�&�-5w:
]�0�JD���*�qA����O�i|�Z���NX�@.x�yӮ@
6w}�^[��� +:H�|�� ��� +��'#�>Pс?�؞�O��991!�����r�m���:���+u� �ERδ<���Q&�)��91|�1�H��G��E����Ȯ��$��� 2��b8p�Z"�v��*V�'Ĺ�.��c�f/s�;��;S/l䴶�\���E������ƪ�chտ^�IX��j|T�'����'�}�R�@ ��В�t��W��+g�֢_a��e��i-iϡpJ�Eb�S�xz���D��o�ֈ�A�;�&9	��1e	@��V�\�f�����0f|ؘ}���ŋ���t������5�����3N�����2�+��M҅�C�&�Ο�e:��Ʈ����AA�I�3�uW�C,E�īl%]����
�ܵ�!�s��	��u�����7����x{'����ԞK���%J�G|)�B}k�aG���ܖ�!��B�=�i�6�P�q윾/��;�B\3����FZ{V�qa0!i=�)�b������o�^�72R�W_� ˽E� 
��Č*{���b��2��� Y>|�)pЗ"TX�O!�qcO����,'����R��t+�0?� �Z��G��OY�,:��R"�x��`LU��J�5u9�����wxϿ�>���?�+�| O������X���@�7M/����^��R���C!�}= �E�\eœ=/�H�ļB���G�,8��/�7�j&�&-I@yL��01�/~�o*͑Aǽ�f�az\%�5!-��+!����{B��!�f�Y|�^V���w�G��9㪚~�ib�u��,$B�B� {�47��v~�,�T��D�^~�a�2�+b�K������-cY�X��un<�c"���I*�~g`�D�p�c����
Q�ϼ�);�ܰ�=-�����U�l��E��o�IU���/����v��y7���:�S���즭s$����H�a��< ��}LT+b>6����z���%`hy��M���{[@Z-�C��0|'�7���輚�J�3��d޼ؒ)=cl���.�}�T6S����;�-1�P��Uڜ��w8�{�n�1rV�®U�pX�e���T*�o��D�f��9w����TO#=7��M H�`qİ��"�p�͠b8&�L�3O%�Xr����XE�r.ї����"��rj8�3�>y��%���LԂ?��Q��]�M 50�����!<1�G�[ kƷr����1$W/��Ʈ��A�ؐ �$o�  /&z~D�����D�!{g��_�`^���(�צ̡�t}�O�Y��|��˅����	�I�o��>r�#��<ed���*|Q�����ͩ� O���9C�M�#lFF�T���_g�S�O`ɉ�ez�[�?�ܦ��c���u�V� �υ�E��m�-�z�S�k`*�F��&��۾���yV*���{h�klM���&>�p z�Ry���Tߎ^�5��o��tǨ�/�]g��P��n�����c�jk�-���s�o��` aY	!�⇳���̶�L�U��*s��l��M�)��@v�T��X71�;/��|��C�ܞzQTiA��"�N�W����KZV��0ܐ�;��tK����\J�s�C����Q� �dm5'��_�A��AV��jYuV`Q�YB!��:�fm����x��>����~R����$,H�{쯸�����(e:��r,�ԇ	{0���W��/Ʋ)�aT>z������a����C�md�.����g�6`���<%�i�˧ �h7}���hw
iP(���o�p����z
���W0?>�(����m�Wu�T!=��2bA���|�05��a��^_�}�Z���u[n��-���N�v�.'����Ч�������I�T�,��"4��D��,�G�ND>�`����Д�߷?q����N	�� I\�אVd�vXQk)NZ��F`�R\�����F��rUP��'u�)/0���o`���,}�� G@�H���������J�V`4��'��������6��XI�-�<y��)��2މ���å.�X��oٓm��%��A�!��@�E�|����*���
u�}@�A���
�0���Gv�@�`����vǾ&"���墨�vH�{(�8����*.P���#'�&����Y�#` 7�-���YV��b�de��Jش(���4�5���!wF[��fh��uG�F���I�O�Ŵ�	��$ �DK_��7�~��Q�Q�|���Ly�?'�~�As�� �(̩	;�Ԫ�<ln��u���	,5Yzlaj����V�B�N
�<�x4	e�ut��/,)'7h#7[&;��4���&C%���j�s1Rl�Q�Y3�7!7�hr֞��U��>�����N,�I�ʢT�&�lbJ��d���2LΒ��%o�k�ylkj���|=V��; �%9Oa -|�zyZ���b�m�X�Bͭ۬tc��_
2��]�y폻��	�=ٽ���a��
!������X��Z������j`�0�#���uc%��sƒx��Y�.���}q��bg���	(�^!�[��lV+��qܭQ��|��|�2�3a��bh���-�o/$0 ��\3��8�	!�j����Ta%�o�Jw�Z�k�-�o�å��+T�v����Td!��`C������O��-v#�3�6gW���@�%�>��>҂��=�E-2u�`d�
jo���D��z�� ^t�NXv\������]��F�ɧ� �8;�Z�;�0�6l�(a=O��A���\ <���M�溘˰�5woʕ^�.��t�U�!���3�:�����#�+��X7 I n�s��P��=A�=����ICF�N�X�-S����)$�^�щdVΜZ� ��=3&����uxQ��) �(VN��L6��I� ���-���eQ�Y`�vIֵ�Қ�G�Qv���(8�Ձe�܆IN�o �/℘(�C?����_`Hw��N�Չ��TuT�!1�]y��h��*��$���.�@y�
���[�DE-�/�Ыt���������x�F���zJ͖�J��:����E�b..��V�?"�R��v�08x��8U�F-�S+�9�S:&r[C�`��=}��?Rb���LV���L�d���������FwZ�s�7�՚@Mt(&�b���K�J����Oa���u�}Ʋ�Sck��\b&Ӻ}�0O*rT�!��إ�5���|��
X,R-:'��u��B�>R����8Gjڝ��Ή���k�xǟ��VE��)ԍ$�K�N����%���m���| 5_zøz�|�D[���%��
��2�Ŵ��Y�ЎZ)�b:��n�x}�j.K2Yf��eG�X����d��h4��� �\/>����[��ǜ�yj�x[��[�P6��HB?I�BD	d5 �9d(
k�$�d36�{Z`���|���7G�_��,Ό&��4h�a�S���9��Yd�#�nOZ���z�e;�8T\����\Ao�kz��b��Ӛ� }�Ti���D��$X�.lKsj�㸥6X�+�~��.)�O">g&>$J(1��Gw��qO�`���@�u-�m`x�)n�:��k�	�������*��3�tK�����T�j����o3�b؊p/��7���IUe��^kU�f�l�o�H�Xuo�8��L�|�%�ݟ�)���p�x�wo-`��x��_#�y�7w�����:߼D��΀�+G@�,e��,�³&�œ z�6��yЮ����`A���0�q��ŉ^�v^��}��"�4X�����gUR�~ꆪ����6��S�M8]t��n,.�d�?S��=6��3��H�U��{��<���ڄ�\���x���x�;�S�e�Rϳ��	I�$&v
vJ��Se� N�Avͬ!����L_�<]Ǎ���=`y?�Ͻ���[k.@M�a�Y�s|'�����PX[�;������s�h���fU�,4�Ӧ��f��Y�R�%�n�Qj���Ի��uG���2���m}W@b�n�6��]ع̓X!�xj��+z��ڂ��`^����ݧ�{��̸�u$���sa�M�d M���@��P������M&@R�+30��bx
�x*�
i�򷹷/�V�<��t
&[�&�t"�����z�߈6H�����']���s�2j1:؈���!�y�h�U�n_���G;����މ^�����K���U������sE���J��)�q����Q�	?���P�.
OM��sk��W.�b�@[�A�^�bH�')�7�7�_��s�x7��?�?�.�o�ꇭP�	וS�k��Ҝ>���c�����*B�p�$u����I�b*�Ǩ�k���5uL�/�TЌW<x9�r��L�dHV�[��*Q�^�s��/{6�$Ub>M���4B6�"究�Bl�J�~tAc�<���:}��)z�c��q��+{��tu����X�:K�<�{]�Q�3�O�����T��Nl}$��Uc@�:�5	.m�1Z�Z��f�ZV!¼e��@uv���{��ϴ�����	&$-G�A_���IHТ��WM�N�a)���������q�����1 kw2���8�M�q�q�{�ټ۫����-౓2���e=+m2��^]*�2��~n"��0�;���ZL9��~G��nUB�̨�_a-�^�|����Y/S�����������ٗ�������_��u�z�fz�yu�=��3��1�	���H�*j�i^�8�ݛ���uv�"��z���9�h[کgf$SnzyQ]I�:���>Z�*I�a�"A��"Q
6JBP��[�Ln�"[���ق`1l���� ��ND��)�~�x-����$>�43K�;Y�E�F~0&{���ת����捩g�=�0H(DM_s�.z�p�vs��v��Ν\�Dg�%�T(�u#t_�5�9GI��I4�d�/��ł[��Edi��t�K������"\��s'���#�� �n"\M���yxC�ET��͗�a�0���Ĉ$&��_nbtq����%QV��w^5ͱ��l�T��Ԩ��J�u���8}�Çd�<�);���L��7����f`�b�y}�+�eĒ�#O�λ�Μ.dd��W!���~�b"�K3}w��h�QZrB����6�KV��Wނ�a~� "��ǂI����EUS�D�d�|�+����&�A�쭻<�d�t�]��
�0ـ����C�kv3����2,|)'��@�\^�G�Z!`��$�3�P�J�x35�����jS�ȋ�7��|�\��K��![�+'�!k��]:,��}��W��+Y8�f1b*]G�(�8�/%m[дSFY3)S��Dˠ�Ƙ<�����}�qo�*��1�VL�;�w��1�Β�A'��S��@/Ma g��/����
�jL�L�`�4�!P�<�X�o����Wמ�#<��� R5�܋�,o%��w��x���$��C�*�e���G�"�I�R�b�;tw�ܵk���EC}�i�o�a��rFW�Nၺ2?�	5�Jk��`��Ze��ߙ�@�f�Sj��?([y����a����1�9�#�����Z:�Y����ޱ�է�g4��E<MŶ�À�I����Y "���X��#kq#������4 C ��,7|���|	����y#�ϦQ�e���w�R\��~��x�;~n0g���i4��A�.�[Sٜ�w5�����~���M��}��]dD�Y�\T֩J�d�{y�8i��B�K���".��tk��Y[�����f��$���\v8w�#����Xq�����pn��ͅ��Ux�����І�m5.��"+�<��O��4�pč�Z�y�3�X�/z�����M�����ޚL�e#����X�aG���vy�<�l	|�ϧ��N�vA$)Jo��hҭ����ɭ9���M˰�L�	0Gw#i��V��)�S[���c�J�C#�:6�����G+�߁��
��iF��!U��	��� �11�G]o���ڕ��V���X�Q?�v���/�e���i������lK�� �fL�M�+�V,���޼V����W@�r��n�E�3Z����#�Sn��ږ���N�`�	f=��M�Uxʠ�G>z;8`������&�q��o��I'�7^=:�V$��(Ni���p���ۜI�Tܟ�}�ӝM}v_�pS&056��#Q� �c�IJc��&��\Z�,����>C�sЊ<�lC�8��v����[�J}5̻S�I}��S��Z�;2F
W��s�;�Y���Q"M)���]���v�0=�9�@Jj��g�X�B����X�Z��F��+j>IBS�E�ق�n�u��X{�V#6kx�)Aq>����L���c?E�����'X�z�Y�ya�w[�-.}7��x$���A;W	ï�%����`�����#�KZ���/g�b�`���I�f1�w��)�i�\=�}>������H�w�2d�ǃ���=Vj;%u�����n%����q�˻��I���ٴ�sZ��_ٳ�J���1�`K���!��\Tt��7o�^a@���χ7�L�r�W��ݧ[��s����M���2^��jh�&@��/�s��q����^E�����2�[�1�.�eݛ7T�u$��u!�[�$�F�U�&@�J���Fk���)W�
�?��Ũ�f����5B��,yo ɖ���2����|1a6òy�<�������-�U�/ʟ��I��,��9��t?q��Y�P���t�衿2�ͩj������]CһE�4~^v¶8��<:���*�9BOρlo�l�� ����a���&o��r �*��`o�3H�5KF."�]�ХJ�}Ɲ�������lC��(ñ���g�9S(�fT��ڥ���l���Hc��:��!�����2���t6���I��[�n�J�)�J?��	?�'
���0B�����PP�Ǫ��^�X��u�;�+1]#d�:@̻{ǂ~�Z+�%�c���YA0���j�կ�U?C�i2�� ���&��X�=b��:
���X�Ǵ&M j!�B0U�Q��rw}:��.��>�����g@�
��`��$�{���� �TD�n�dQ�p�J|9�!n�|�ʯ7�rn|����#'"����w�b?WN��b��Y�Ś�f
��ZQ��z<���H�A�R�-"K"F�@�K���Nz-3��<�}"���P/�)7��˹�5A��J��"t`�� N��|�1W�JBX��T�����[�x.��"��Th�r_x׾�͗7{h�6����J�$��F!��J������{*ߴy��!J@�����$\<��o˘b���Q��lP
8,�	�ċY��<���R	m�*��4�6=+r��'o���~�pn�]C���*�ms�uߤ}�_����^/2._׿ozǡXӣ�ʅ�P�>GS~�E�����]��>}���i�cm��-��3��3�wn,�VNmz���Jz&������aLX8J�4L�� ���p���3���o���v�K��gH����[�q����G��Jo`��� H�v��ᣦ{��K�ܵ�}ܾO[��0GY�L7y:�Z��qu/�C���)``�bC@����a�6}��P���ƚ���FG!�� KS҉����s_��L��N��y��o���݈P���_�=$N�$�(�p�a.-��Vl���M*�\���VU/��_c���?�@eI�����%�h������P8����MGǤ������Ծp�tt+nk���>}Q����,uA��apNo��x�a����m�TR\'|��69��0i�$�ԧ.�z/��R�"c������=�g��\��!&�γ��'��-�&�����Vq�x@S230>I��c���Br;��§!ێj2q�g���&���4Y#�zsd��s����-5{J�No��0�~�{o=I��������W����2Î�#C������߁�����&)�"c�p�-�J��Ыt��}��m��%�%Eo�|�䣸?P��rƌ�6?S�X��0M���R;l�=�7�(��5�\4�;^1��a���灹�	P�O��l�:�
�@��S#���"{�����M�.�O7«afJRggx�$�^^���t���&�36��ЩjyWD��l����W�~nd{!��؍x��#uI�nhNA�H�z��L�����m���OĄ%�ڟ$x1s�wy��:1,i��
&�����GĤ�
D�>�j�D���Qc�<̓�Ǿ��M��I�ݚ(Z�S�D���ЌnE%Qm4B/N���[B+��Q�m����*���a-Z�
��\�8��24�V
?�-lR�1�v>�A�已�I�WYN���Ty����̮�O����9��+	�~Cl$�����U�R{�$I��,prs]��v۞KGYy4��˖�k�k�Z+�HɈiJd�jY�SV���������r�;�<�u�p�����vk��޴��:��|\�����bP|ƿ(�9#X���?<ah�q�F5&Zk�����5����fg�:�<��>�Mf���u�qNS�#j#��En�x�Xs�{�[�W	�g'9�U���7G(e�\�`�?�3SW�KC�|ED���V�9�ڜ	?��,	Yzr�������>�
�t�R��6SAS�a��(�ǰ4��D�3��*3u:�&�O�Qls���cM�ƱEv ��<�4G��{��-����Lz�;��=O����2��7E�����sHH���
B���c'bK�m1x�r��I����n:I�}�ȖDY�%�w`�d@�ߢ��:�f��N��H��d�+�&�_��b�?�V�ת�{�(��%�5Vv����K�s�~�zAN=���S@t���I�/'��J]��41�q����wr�/4#�����(� �t?y���و��8K�i�rC��m͊#��Z�b��ࢅ_�>YEw�`�c�����öǺ�y�$���^����.P�� [wB�z�p�2裣��͉�`/���1�[�n�3��Y�i�P皠<0���<?�V��S��K�ʦyz�����*�nx�,Io�H��v,�K̾������$�WP�8�P)�XA���<L�?O �	-�F�8_���è[�s9e�t��e����\��`�ܑ�J��v��O��yzRw��{w����#M�z�ɸ{Sp��6�s���Ӊj��"�O-?���Y��r�H��G9�/�|����Ə��&�0��Tג(�-P]K�%�ڸ 3j��i����������ʳk�WS�4������¼`/=�$@�^E�uK����)Y� ,��!�t�%�-e�	>����%�� ^
>?��%	���-$[�[�� ��yg]��4��.��2�徴�����iy��"&ڂ���(F���XI(:y�:x���/R�+�A�`��$��9i�(��2ߨ2�kD�-/fk���|�Z���h��4� Wwx��"�E���Q|�^6� ����o�I_�t:�d��E�Q_�*0�	gC�n �-=k�	��4�y�ݯ�g>%5Sϟ���X?,y��5�4#���4�_�(2�P�0�C�j�G&_ͯ#��s�8�={� �	��#gD{Sh��]w�%4O�A����֩�|����d��V,����a�[}uC'EDNx��!O�)3~o�g<7
����d�K��ߛd�H1�u�ꂸ�?{��0��{_;�'��Ɛ���V(��9�1Z�M�9�>tXP��3��$4���[�Y�yq����TtD��z�K�fvc����OO@<&1+�}Ye�ik0���/��`�w�.�Ȭ�0�.��8f���A���V=K����;�����:d�ʬb u2.�2U�[KI�%O:�r�C)�t�dg7����w�"q|�ܼ���R_�Ĺk�eQK�Pee
���}[�j���?