��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� ��
�˿F!����i�xL���G)35�У0�Y6ɓL7ɶ�4[�Z��K!�Rʶ�������*�r��u��@
��x�·p�0Bz��#�;V�kg����[<$e7�#��5�!��������Fi�=��Uy}T��%�oy}e�5�H��|�ԥ9},�&�?2��Z-|����������ߝBT1Vs<��s�)lE~/Smv���(d��1��U9	�
Nn�Ҽ����Mڵ�Z��O�dmˍ{���ȍ��}vT-z��s�����m�Tp����}}xAd3PeAEh�x1T�%�H�q��P�uiX���^3��]������s��h��l�X����'��.�4�zʁ�=���ͩ�p�(`;_tO(o\���_�&M
:.�q��u��M3���Ჱ�a��~�.$3�A8�M&^��4��u�Z&���@5�'��i�|��~���u�J��(j<��C"d	����u�F�*�Jڴ�d�7%!�Lc��7�jj��p&����n3����)��ہ�V�7��p�h�S]�d~��]��X�ЁV�U�W�j�JFj,�W�l���[�1;�.?Y�$2�ҵo��v��!}܆��:��� H41h�l�j��n���1O���y�Ê 䢙����iw�P��l犴d:�2�'�ɠ������!�Y�E���,m/��r��T����|\�4��H�v�wF��;\�����H���e)0�$)�k_a�w2�:'���|�_�n��2�<��#���xu�٫jb������O�">&#����>�'�/����6���U�27׎�������C^2W�.B�"NJ�̌G��jHH���8��x�Ww(��D� �׻o�d�C�}�?O�+�Q��4�V���%<+��3������EBoIʮ�/�&C�9��O�*�OC��m��X���0����~�u��h2\��ɀ�LZ:`d$l���3z�X�Q��o�ܥ�>��
#n>bY��L@��cXA�؝�M_FP�MP_w>�O��T+��Wj���
��B8��`�S�D����?e}�k�z��M�ƅ��l��S��xˌ!Դ���2nl������1�l	r���d���׆�Q���!��#�Z�����o���F^���V�ы���?�}�w�G�.�lm�*���6j؄�2���<�)^݀�2̑�dj8R��K՜snpջam{�0�{%�O���f����Y-�P�>Q��j��[vP���}L���B��Wo��q|y�)G(@�練=7�__@��d~lT���o\@˲��aQ�ns��)4�29��?��N��4�S'N�i"�6�da�m0w�r�9�i�
t7q�mD�?�
{�A�["@��E�82XU%O�O��*��f[~%�]�>��>=N�R+��n�Q����aG_ܷ!�ls��أ��3�[���%%�B��Q����(�� Yp`��Qp��ö�ԔkJm���[dD؎=�Vbf���S�ĺk�1�����t��^��f�Ť�}��X��I���>�}eXWtraCдD�$��3[wę�
ԍX/�f���&h�'�>�(�g��TI'����H�v�Y����İ>�9��r��;�N�h+���ҟ��ں�K0���T���)Ҽ(��uv_���3��z�eY�n���i����ϰ6]�c�D(st9��$sA�n��8'&ׁ�c8δ(�_���aeZ>J̹M"�7�^�(�t��Gx���훂٧�y麺�k����ת	� �d)Y������$��y��N��I`Ҡ7�X��(\UJ���r�j�f���&ܴ�B���,��q�*��_����[���%�r�~����y��&��P�lz����4�L�K����u\$:<���m&�Mɕ�OFY8��|mԫwR���k�S
�_��O�)M�`���gm���y3&J���5W�J��ey�}���q��$�g-$���ȶmgu�a|9vU�8x2!�b6�:�������N�uZ��� /ǋh*��sx�l�����2Jʵ*�M�juS<���p�H�'�M���+�X�꛷�����`ܡ��]�{8����?���hn*<����럽�u`��4߾Uz��U�|�xd"q�U,��@r��Ty��] "��P�\p։y�~�+���8ֹ���}	�]��K9�$�.}O�-p:��:�w!��%�ѝ���?��љ/v`��Ar�^g�,�V۳���_��-r~�[�lt_��2� ��=0j����df�u�|�1��2�h
�^���4m𴳄�̈K�\����Y���R�p=y�N��9[o81 �Qk6!�'t1�wL�v^�$��a��X����Qϴ)���q���q��&ؠDkV��#���a���gg�ұ�U ����3	��-ʼ�{��jƇWo�[����ǓW�;9���ƨŝ�]�c2A���w\V�6���k!��;�Γ8�B`f��t��n�.�_���?�t��I� ��X���_p���4�Ѷj�����B~	�MX_�`6P�cU��lo[B!�D:\�;'�?0�R������:��N.K��p뀱u�1]"�;m
SHG���ŏ4�[�@V��iЈ�=\����{ �?jI*�BG3`�u���I>|��#4�i�Ɍ\h���4�Å��)!�����z��HY�v�V겿���9�M�Ϙxsҙ�K(�-�ѵ<����n���}�CQd�͗=�qr{�
�ݏn;B�ؗԡ�٣�͑Q�Z1�h�0����%��m�[�ָ�b	0��"�E��6ײ�_M/�C�	dP^{[Z�RS��*��0�N�'XX	g��f��gPA͇���#�l95���ƀ�J/���q���F��ߗ�ͷ�����ӿHbŋM�tx� �}'�I��I2v��:�֑(���-�����ԇ9R��Z��^a6�c���:�nD��'d�]G�H�@�4"Hg<�WqY�\�ms�?��5iu�M�=�dHE��O��_����J��wm9M�@�����t9?�!M���ڍ����ƃm���w>���e�B	�0�1��i�ku�k��<�ޛ��1���te!���Oܦ<�S���r:PT+��V9�p�2�&��y������p����1�:2qڜ�ڳ�ݸ��ʫ��0��#������ �j�g䦰|��gԅ����&�G~v��j�
]��j�(A,8�o��j�c�- 'P~_���	��r�5/��C�NŒ�����_�4K{I�PW/*m�Ν:^AX�Pvu�]������������M��!�E��H�w#8~:g�qnC�KY_v
AV�����܉�\��J�o�i K���.���2�$QqZf�8Vfr�y��-ω̦
ȱ�V��m���h̝ޅ�����u\�(ƾ�`�nX�����U�O>bq�+�d�^Զ�3�7���Ą�O���ǡK8Q�<�vû�&���SE�9O���R1>��S�۫������*&Ρ���m����A8�\:�MTf���E�f�Z�5�Æ��y5���L��ɒ�?C[.n���-@[ٰx>��t�y��D�/��?��ſ���Nts(}��&#�-���{�!s�|��8x �6�Q�#�\��<�+�2�`�i���z��+P)��KM������a��;�Շ�vנ��d�n��7�o�r�j�t��h�:��8��h	Z��}� �E���/p,�rj#��f �Fɜl��g�x����[��I7�LY�������L�Ė����� ��/���*$��=����gd�&o<��-���&�s�kwVrbac��"ci k[��-���3a$wF�{߫ �i<W��s�c`���T��`�_J��Z��]
{��G?�nO9L�Z2E?c�S02�m�B�b���nS����O�ʙ:�'D�A}�^?�ҟi�� ڙ��L����'�lAj O�!�I����Tx�l�0�e������<�p*K.��w�H�^�y/���\x�c���c5� k=����=�>���q�?Te�a��f���'7�Z��P5̴�ķ��_��G�,��{�����B�r����$Kg�i��x02K��<ʮ�E�ҿ�J��U�ai����&}ͳZB�Ɛ�hg ��?�%b&f�������v���+e���P�TD��ޱu� "5H���T8A�)�O�M����%�9$h��I���M��~����y= ^Go����h�nY%� ���oI�&V�s���z��k�ҍz����3}�Y�$��b���qz�a>��*d��>��@���;��9�9�\���'�����_vrV���Ң�]��b����݊����m���(��W0��h�|��ccպ�a*�D��m�>�rȪ&�Ғi���M�qղ��b�`����ٵ��.#b�Ѕ�����+ ���@6�,b��p�֞ӛ�	�:$��\"���y��if�ȎY��wo�O)��K���"��������H�� wṒ���BxP��*�0��]Z��IҀ����U8�Y�8W8�F<A�S��]6�4�0}u�쳗��wi!m�FU�2�|Uus��`���ӝU�������W��,��_-#k���+ܝ�t�Rm+���qiN� �?�'Qc}����Ҳ��9j�R�G���YƆX^�������$�q�d&�/�C%?c{�������dyF�J��{Σ�1w�����bγ�h�`Ы��	3���X�L6� �ۤ��N�ɞ���3d�\l-��̃�݃?1��&_���d�^|x���W<��l@Ph(��m"Z�a���������MgU�n��7(9�<<��?į۝��Hr�K����uM ������c�#[���}4[h�ι���w��\?."���#��1R�HP6�21{����+�����F>-���B� ���ҩ��|�<	��ybB�#|=ɡ���I4U�6ʒ����� m���\|��!�2p��O����-�r]�[���ӓoy͑}H�;c�c��	�ݦވd�08�+ĮǸ�^#\&xޝ����o	D���$DKs�)"�j&M����� %]�^X, �%�4T�M�	̂�$c
���Pfv�*IǢi��'� ���Y�(��|W�d�Z3�s�G	9����ʿng�2a��u�m�x�_����5#4�Qvi�nNG:�>�<���6W�;o�6�G����}�?��k�����Ov���8���K9�x. K���Zz�T�w�{���WO5Z&[�G�硹�ۣ������0��I
�VjĔg��nw���͌ۗ8��2c� g�N�Ì�ӭ���<ꏝr�d���C>`}|eY�
-�7�]��(������X��W�BQf������zܲ�o8�"*�b6�c�A
����4?v�����([X!� ��ZKQ�Qy�3�3D�������--�9�d 6enZ��=�wh Ö��C�
V��.�j'����	�����jY�0Řs�E��J����LH|�>
��g�pG�svi��t�'�m�^�d�n�Ƶս����\�xO���#��JчdU��p�^�l��3�a�{��������k?-�\�k�6�NO�ɝ큝��-����е�*���Y���˼n�5 ��*Àxx?���h�)�����^x�I�o���I���"�n��Cox����'�3ϔÀa�)<�Z�R���uë�ĭ�_�-��'��ϗn
LƔr��Y�/����4���o+�Ri4��4�/��u�O��;�-�R'8.��iN�a�*���'��k`aנ����'3��#".�O[��Ҽ���	ҫ�2�*�E�:S�Ů��9�k<'n܋�Q'/�J~rӛ|�<ᒢ�גdϭ�����