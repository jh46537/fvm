��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���Ox���0��?T�}�D�yBl98�锛�l	`�ġ	d}�:��PƸ����~��R��o�K�jV�,R����vy���3����O���Z�����g�̼A��v�{�7
��5�¾����B�C����������r}�:ش)qqa���·����BW�4����"V�CL�zhXo�e��6kT]xl(���%lT'�W���'�N�V#�L�`�`�Xy�6$���:��9I��ì=P��uS�I�w��������F��<��s��y�i�u�����ml�G")�O�4����}�,r��𯴢}�鑪 _@�y�Tkt}��8!�JŜ�>9��C �gl���-����{���Z�*� 9�[�B���c�M�͠�+�G�Yy"TGz_'l��2/;��	^F�/	b2�ܕ�Z���./k7iǶ�>��R nS�}O�i|�y�AP?e޽���1	D�9U����	य़��n]�n)y��u��IRe_%�I�����bmZ�IK*�~R�VmW����Y�{~�VF�K�\��O�K%�p�jاb	�.�!�-��/6u\��m���^XM�Jʃc�LK>#�*��V+QHY1�Ң�F�gϵr�BG�b�]+���A�k�`k��^�MI�j�bm4��Y��M��8\��*�mB���n��-��}�/���kh���ƽ<�����Ld�4�����h�!�Y�)���B෨�qK�s4���~d��Ӳ|
���J���Y���G�"��WçU���{���\"�]R��.�}�AH,2M��i6�N1(A��}��F���C�˽���?[S����P~g��1\D4U��}wì�גB����%_��ԣ~�,�5��<<�j'(e�G�$��~er�I N���:~x�0�(Յ�\o�s��q6L���J�υ��1A��\�n|�p��(�#���c�=�xh���� �J�[y((\��mx������8j��}�߄�ڎw:j�Z&���W�E��p��.��*�MŪ��FQ��^w�1/�sҹ\S ��y�&uAAܡU��ѽ?6Iɦ^�X8��9� (��V��G׆���t���G�Rg<���Q��и�Z��\F��y���^v��~��6�_M��Ni���EH��C�6v��Ua���UH�3O��(��
���3%+��E��,!Y:�\��#���Β�S�˜�.��.c�+�E�HD��p����a۬��aZ@��x��ԥX3摍��e:R�O�,z���4�Z
�=9Fhܭ�8ד��1{�өw��z-03��@w�	��t���1LLLD̳�r���6�-�����|���NY����e:��i���߿��2���G6�͘��7�O�ik���4ا�{1ğ�(���<��jn�f'�ŕ�d�5���x�A����#�w����i8����[���L/�|�Zz�z�k"���a'������5�I!2HN���҈���:���I;�@ �:�
�T��o�E����=ZRe��6"Z�P��\�$v+��h�Lb��j�8���|�v����~k�r�z���N�1u"��P��隸�h�~��<7�D�x`�i�ZD�I�%}�E��Py����L<"�H��]�E�vmӫϔP��kl�kǕ�V�U��heV���z;��m8��q���o��\ǋ���b�]㙬�^B�t�d����6X$,�%Q�_���������}�c�R�p?;9FCl�t��>��@��_�,���e���R��z
AZMɦ�:.j7��.�	��:��qg��m�w�;�}ɅĐKb��7�P59���Du��z�+���E�����˄1j 5	���t���ذ�kYS�C��8G{�ӷ�2�j	�Η�'��`��-K/^�r��E�L���|ކR��ZBC�AT��Uz%/��!�7�v J�-���(»�o�0�jG}��I��*�\��yI�uhfK�`��խ*F�g�ϥ��@(O�zH�)L�Ȱ��/gk��|�1hw[a�AKj^o#C��׌}T�h���(�-q��uJ8IҮw�(�g���G%:j̻��¹��/�	�V2��W�#�Le�p�@0ܸ�
r�X����X�ah"�Q��^0����`�*�x&�.#,E�i��C��J@��;˗U�憼`��UZ����kk��BRZ9��C�*����F]���Y=��ZJ�x)_m��?��T9�<{�����ڥ���ݨ7���>�7��55d�����8��aB(��%P$T�}�@�TR��x�����KKΫ�#I\�@6g�{�(�\7��eC�H#]�ԏ�q�]����)�b��$�¥C�bġ�Kz����1�ؖRaR�[�lʛ��]���O���R8��W��YW 2Zw(������aؔ�m�u<S�f}���Y��ٵ�c�!i��E]I��zO��|��]�����sMէ�.�7�gL���A�4�얙��m	�}��*��s�����A��o����7!<Ⱥ��R'�j���lb�%�%
w枚�#\����qK)7i�o�~z&�oߚPAc�=~̙B��Ԗ�F�i.c��U��"�~��؅V G��}י��9pp���
�Av���N�i��wo��|�E��@���^�q�`!�'o��`���%;s�ͱ2�e}��_d#�7;˾�H��ŋ:
�P�I���/� ���k���'e������.q�	�f_H0�ܗ8J;�B��ij��`�&0_��k>W���A�;�7�>ͨ�j�{4,�bM;k�LU���	��{�F��;�l2)�j��p.�������L�4�g4�.ޮY	K`�Δ��;�= ��i�)UO�zU+@�b,佻%F�	�/��]��4K�0|٦�I�m�À1vCm\��T^���@6����_*4ヴ1������*�������}�?Dʦ$q����� &,���'����-��rK ޚɤ��k��Z��o�j
� c��|�QSVZ�n�*X�h�f��J>nT��*T����*�Nx�{���c�	��ȉnA�]��ې���*pc'�T	�B+E��q���cq^'X�w8�� ��A�]�p#��X�1,�q��>e����q��ǌ_�#0�;pߜ�@dDBǑ~��d@�����-�b8ٝ�c�!-]Y��������c0�u�C�&G��o��6f���}������}+��	�皉%�����?��@r�,�$o�oИK��ΕJ��g�ѯ�7�u������7c�ap�Ǌ�G)$�)݇Q���ca]����rc)勭������������k��*��S$r)�C�@�H�H[��,�	a��`�V�X�P�'y��d�7�܎.��l�����T}9�|�̇��k�*�Z�VV� �X+��E�P��{��K�v��˧��E��;Y����O-�.�2@�nXQ��z�Tޞ~eﳕ��҂:��z����>���
)qr9�Ɣ����O�yWE�I�٥�o��`G��:�Wn/����y1��l�@�.��[�gr����Q�wwf�3�fM�^_"���>/hfc�Ȫ�����<�N���`��9R�kp���1�&]4v���7��%���JS�
�${��D���]���vA�Y�[��\R;[��Z�ŲA�y�zu���NP�/9��qIZ��}�j`��K�[�%�*��>M�e�_�޸z;}����$���UI*�BhF{�^�g���K��˫��D�!� �]3)�����N��s��9��yWb�&��y:AF��/��44H�X�T�O��8�Lp+ю#=e߭�{H���[�����(�f������	���#���+ut
��q��7N�w�;py��HG����e��5?.��C�:Cҙrmy��o�yiƖz�˝�p+����О�M��?�cD����C�|ȉ���6�9��?YDWFi�Ժ�4#�42��?�,��۩M��&���7��0�����˻�'��c�������yb��!9�[!��� �B�������e3� @�AF��Tn�$���E�4g�� Bx-�q"g�"������bnۓ<�3���bfzk/yt��D�
[?�h�!�ѳ��da;A&j�6-�����0�0v8�XH≥Y[o�E���I���l�YՈ��ØӼ��Z�~�+Z��0|��(=������� aiص�@\YM"ψ�� ns�=a	gT��,Ŗb���b���K���$ >�ӐWt\��M�8P�6�@��m�L�+�K�z~������R������N*�����z�=]��pQ�Ey.�{Ro��z�v����Ayz^��7�����ή�6n~��3�J2s��S/�eY�s�[�H)ڔf��A�`�e���"X���:�'\�w%e�O�����/A$�����E��%�/�x��G��S��09�$)^Xԩ��&�v,�:��OX�c/(�Զ��k�M��[� �� �M��7�����q��p�h�xZ��a��\J`q�RK��O���O���w�]���
>��O��	H�N@�0�����X��M��	�֒A��{�C����"�řG�����j�����n������iq5h�Jܘ8�[�}_��v�4ʀ�F����v�c��?]�]��}T`	�n�\ţi�cbl���}n� ⻃�i#�$*ߛ�p)A�^S��Tz}����{'Iλ�Z�t�i�Ȕ�V1�`���t,h��O=vU�����U�.u�h-�,'�2=E�~������w/�ƴ�����u�3<R|��8���k�� �ۼtTd����Y��t|�vT�d:��5$wg!�V���s�s m�?�$9�2vNr�h�Q�u�$��I;���mx`sQ��t�����o �?��P�{D%[; ��ܨỸ��<�������e\)'�-$�P�~���!L�L
J��GA�I ��ӯ"��a�u<�@��<�cK_���;�K�;5�A��b<�^>��ꦯ��"���Z�`��1�p1"UA�����a�ò����|B�.x[9B�w����f�χ��;�6�R>�r�~�[�w�Q𮉲�H|p;�H�7(��1���&�H�I��]�vh8?��g�,��cޢ/�:+��H.�ŗaA�/H��P� LUR���w��B�4H�����(�<�}/����:�tf�*��.K��-b����5�3Q���ޅR���Z>9�yt�}��z��Mx*��4��8�²�Z�Qb�8�G$��%��"�n-�J?Gؾ���sg�)}���	��Y�ɔ���nQ�(�)B��#��g��=������&�}4��0}�h��lR�6�6�X�5q��)oϨ_Ӧ�un���/g9��38����-��e�%�Yw́�i���:9\`�,���t(I�oc��Q�2s���b�<�Og���X��<B�b�I���I5}���Cc��n������p�	#Q�3�˳�AȠڶ8k���>)
bvm�h�f�aa���(1����1?A�f��YE]�\�v����߂��(����/rG�7�����.��k�kNqB[%�=�fD�ҸM���l�uz�_�����D�,ů��mw��k/U4A`��k�N��銮_���w"����0���,l��Z�����;(t�oc#-����QC*���<p4�!��u�wPe)QH�$��oi^f4���+��X��
<sgBV���� ��)\��>�����1P;1@���g�(u F�$@Ps�"}:�/&�`Q�ON�Y����uS�Y'��˄��n��줃�s��,�1��t���x;v���
�*U�7��>���\ܘ��f��l���pcV�D��`sb�'=�6n�d�5
�ғL��̃ʵ���B`�X�R��o?�D+��_�5"4[�:W���4��=��yi�0V
���I3>��F�߇�>�N��|�'O�Z���Ӭ�,�$N�W#�����I/L����ck	����[۪&���,��bx�֧�҅�B!�M'vn�̪F=���ڗ7�]�D0N�uU�g>"ځ��%������I{Ue#���.�"#ɢ���N��8��2=����.�`�� tv(6t偌��[�
��"1��X���{PI`��`U��޺e{�@X�As�[0n���>]����q*r�T�����fR����z찼�&[G�8#������voH�諄�D#��y�T���*���s-y^/����Ϝ�\�щ�_o�!��V����Qk�!��}��ͬeAh���l��V�`>p�%6���Rb�P6�Ɵ���m)�.�߰���_��,�hܢ*���9s��]C�Z:k��t5�Zo#U4�b��(���Sֽ��X�-h�S?� �eK���W��-5`ِ޶E03�����1�(}GB�������!�'��U-;~U\�m�|��˷5��6zN�C%`~�Ի4��E�AOI���mut����%7�=�}���g�Ě�r�0k�r���]+�$�}\2_��A�N���j��Ʃ�3-����J���KB.�\��fRj�D��?H��ri�j�v��:�����'Xt;���f}O4�W��c�[����a]_@�D2m��iv��6 .��ٓ8�}nn�A�ٌ����Cŝ%�_FWḫ��PĞ�פo��vHt���qC%����c<1����1L^#I:9"���ݟ�g�e�$A���2=,�"�:2�ҵ��=��S�K��`�V8ӟxW M�ꑀ$��\s�s�ver�cUX�4�*���z����UH¥�z�l�J�&8&�l��@E��-�~��J���¡�Lm��ؙ<fAB�;j��_XC�a��4��	ƂRa��Is3��=�8���4P�{�<��:����M/x��Kv%�TK�d�5�_3�C���3Z5�d3�'�p��Y��7#ܒ��萆���:Q;4۩��q�ׇ[f�;�10ϋ��� _��5��*�	c��p$+Jϓ��@�?��/���6i*f� JB���w����	� �ŀ����^F�Z�&�(a���]���|������iE������ivL
QL2�r��z9\�[/j�Cޞ�o[.�*��^<�V�t�uS}�)���C�m�?�q�{������W���|�~+����bJq/�'�0Ց�=�`��S��+m��$ln+��b���m�͏qXO�M��(ȟ�}6�a7�x�R �g���]���@#b{�6����l�W�c��黟噿�ʈ�)��4�Z��^��a%NKGXa���X5�^�5���\x���C{���Y�����܁JT��h�Z���'(��AƁ�p{C��&H�Ȝ����r�~i/f4���@	y�_a!�}\H|q���g��:���|�D�ѕ(Ptd�Mα3�|��Q�]�k�)C���i,�ja��)6.�(ei0u��P��b�L�γ�����Cp����t��w,ԍ�[�N�}`ޟ;:7�S�d�M�!I�Is>n]�l����(B�����Do�7�����{9�wE�W@!ұ+�f�}5���i�7�$P�BCw�Q+�	�A1�x�~�S-��F@�/4ef���6uo[{x�v�b-���,,F=�B�d(\��^\�4��5(�^�@,}�U�Z�����'*���`?y�@�]\��B��X���/ZoV����S1�@��6n::T��C��>v�.�8N���@mpxWH7����9�
T�sZ�� ��Fh�C�{�]r{2�-x�U��U�{]�؈̕h�'��j yq������'�'#ҩ֋�x���,����{Kw��6�cp����� /&[��E@�sn�:��"�HAT�dW\�z<)X�Oߘ6g��t&����>��(;�j@:Lasm=�� ������
u(����̚�itz ��$t$x�
��C�+�J��`9���D��^XH�t_3+����L��P�͎�:а�0��:<�'9������������5vj��hƸx7�l��G���Z�䇆CR�v1'W.���t�Z����%���e9�[�4���E��ѕ�-@ɭ
�҂�Tf�E�f�!P`@�R������ƇaAcn&�5�6֘C�S���x��f��?��Z�[������@���;c�����k��V�	�U �������8�)C�^�k� y��n3���z��b(�$L�o�/9�:�?��&���c3ly�l�0��;�uke��E��)#_V'�HQP�հ��'+d�>4W��'uEpY�:�A�Q�0xU8�5X�)�NN�Q�"�������ms4��)�H���ڶ�!N��˳��!�����.���o�-�޿�G*��G�� ���pIe�t7H�\�z��P5Pj�ݪ;���ɣ��آ'R#@M^Ul��µ�;0pW��RZ���?
�Zz��!C�)�p���#����ULko�1�����\a�;w���8&���1p��&��*�(�B1c�pkZ3����m�
TvvH�˅(��~qRr�X�6�{��Qp$��<-2�fJM��Uv%Y�SA�db~ܪ1���W�����g7Ud�s!���)a�"��M�z���j��^#���Mßo3�Q�:c�Z���Kl����=A�&J	堂�O�
��O�Bw�\��Fz����S/ԩ �VMp<�6w&��ŋE�~��:L����!��V�>0�m_�Ø�d�����@f���-.H�r!Y)�
�F\��[��1\�Ҳ���x5���K���#�C����г�4.b���f�J�b���|�+�d$�����Yi���m\�Ϟ_ky6yQ(v�mF���A�!��vo�{z�zc&��]����E/�����[���e��Mڛ�E���y�:63�C�Ŀ�8xj��@�P�Z��(�7r#��}E�#��j�MO�2�p<���}�Of�`z@� e���dņWusK��y��\6%��=�I���ǉ��!ީ�ܗfƪ��U�3���i��p��N�����]j����Ƹg��0]38�>} �����8��
����(F��[ֈ�y�/�i_%��j��#�3��0�5~Ԑ>�YB���}|��6A���`���\�.�r��BqJд�;)�n��r����@d`������̀�f�����0�x�1Ҹ8)��n���.���Riu� ��4�&@�Y�t�]k�|_�o)�?*6@��$�y��Ζ���+p7yȬM�I�S�:	:`�A\�Q�l�\��[_��?���]�Ě!���[n��L"� Ƹ�p@�
,ȉk�������[*�9v��4�D��4�ښ�H��l���t�i�m�y�0.P�,�X2'�����������qd
��R�C7e ��������.�oy��k%3!:�p��$�l�8�8��͍��cz�B�F�{���!�>�:(�
�p�;)�Q����톃�<%�:�h��iRq!l���k]��8�w��OT{1�^���K�3'5��<*J�E�w��������3��6n�%��e�!�������s���~Iwa$k�#i���t�y�`.}M�&��;t�g������y�����:�h�L�`ʦN�e,Uu',� �b��鹸����