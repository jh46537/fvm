��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��x#PcJk�� � ��Z��%q1���&�%�0k��j�9¶��>�m�{�2ڳ�6` v���n�3W���ɖ��ܣ(kl��ϴ�d����T��'�0v��1��+@lO{��L�u@�0u�h�����æqP�B<�� �-��A�zE� x6�� 3�Z���i�J5�%��JFRǨ�pL��Ga�VsA)9�X��� C.0/��cb����� �r���ݤ1�VC�M�\�� (i/)-�q;<�ƭ��4���%��u�,U�����y������|6�ȭ��Vln���8�F���2�Ff��ڻ�����=�s�zv�r�cu�01v�q�K��A�k����}��	�~
۩�����/y������q<���[�%^�]���̞T�D���9��-��4Z��?�0N{�P�Uv)y����J�B�����]aȠܽ,Xu:h�#�o�6�-�'[u ���9�

Z��3E��3�����#v��~u�Ć�+�<�	e��hRS=v�^�T��`�ۯ�jh<&2U�{{��i��y����X�q�T"$^G���r.��� �4��O���7����G�������p��NT�(:��Z�aq�
�d�G�a��lJfb�|��2�Gq���.�t�K��H�n*(1��nU)��8|U�j�'�T89�� �	��p�E�5�^t]y\8��=W|�M��?�b��f�F�_���p������G�E��3S�#_|��L��}������俴/Bן� �w(��x˷ed�dE�pM��Rϗ�uWV�@.u���"�]�!�U�LGF����fk<�vhT�g$���_>d替n�掰�5��CkL6�<Mۙ�GR�
2WV��9��5D�����r[�o�If�1 Mm����
f��t��*g�X��W�<�g/���W��&�x6�j���f��S3�=���U��)	Qt?@�d�P�[œ�Б�3����N�/k!�@ֱ���`�y���:lD��B��X3�'�[x2�G����)��om�.�[|��@s C���W���Ƽ>�.i3�"�s$숌נ��bf�0�D�f���n�1�<�	���Y;Z�� )R�$�c�D&#O������8��O��)pq:g�F�Ka�N�c��;O�`��͉���m�]\������ Q�7�����P�y��W����D"����S�;�5roy��L���?ˁ�֟V����V�=).̻���lH���FdYQ>Zſl=�d\&�X��c)x�L�cG�759K�]����y��IcW���/n￫��9��#'�=�Z����+�a�[��] �3��\ Y
���9%_�N��V+İg��O^l��OfKt�|���#k�L[3��5u�?y<ٙ���y�S%��|>Q��N���G����Y�s��,��= iդ¯�=���4Hf���,�)�V�-���ѭ �]�c��4x�Cj�!:q�Z�pLe��b��8�Z���K����u����Z�ƀ~���(�U-zk�x��No�j��3a�k�ޯ���H6\�FlT��ega����3k��:_�!�a"t�p���ά ƀ��,i���_�P<\�DdN8�YEV������ڝ"ifUM�o[R��'����'�.�������hG�h�nI^�e�ݽ�1��/<��3��j������~�!ݥ}�Im��$�Y���T'}$p�!C`]T�A�~�xs�|��Q��m���~�)���D9IƚC�����L�?� 6��L�b6�w�>��%{Ԇ��P�����w���}��ݏ�ī�?D���J�{Q��dn_}i�v)޵"�@���B3SD/�󌅡���6��&���`i
V�Ir���AsL//�3�.�&mJi��^1�K�<XHkPP!!��[�퀮�(ԓq(:���m�ܳN����.2B��|G�H�9�*G��W���
����_���#*�dŹ�K�=�_�0Ͻ]�ȯ+bA��jD;���}D�}N�_���r.����Ť��I��|Bw%�$ႈ���<i�l���'3�F��䟋Yhh��Co��R#4���6r^l��Ij́ vϬP6����P���_��{�0�������P��WL��sXҺ[��Q]f�G�%7���4��B���)cR�F�wG,�1�4�MFk+��JϏ"g�8�+���B���=N�.����y�G�O��Pڅu�+N�S���V���ɝe�Z��s�Ik�Q'/R���`nW��������¯�U�&"yE�ݮ����y%�y����ϒ>��,",��9������zBׯ�=2I͌�����a~���E�
j�p��g><\��4�x:�t��(����yf2��_3����N��[;`�CSo׋��2�Py[���qv����R�S������@�i���5j��M!�E�^��)��	i�E<,19�� T���G��ܘ
0��*?�q�����g�n�o��j�g�P���#PB}�j	G�����
���u,:�E�]!�#5�X9sY�$ܠu�mD���%G_o&���[���o>"�S�<�����rQy^ul|�V�te'���CvWTD�z~�`��~~�����	=q�7ߴ؍�[���t+���*��B��_�WY�?���<Zu��7��kvIct�٢�
�9]����0N�l�)�9�I�p!4�Z=�0^�ޔ0�vAŕ��W��⤀�s.k�ո�IIl���2WF��j�6=�LC��|$l\�D�A�����d�=�BIp��RIL����>�&��+�v[m���)7�Մ�\_�m���X�+ے��ɩ]��U��7_N�?�,p��e����otj�a����V̸��ܦ��U��N�D�m�V��2�]�_�����~o���ݥ�a.B	E6���4�'{Gi�lc�b���2)A������ ���U��2��&aG]A2,TɻAn��C�T���"����"sz�:H�Gq,����C3�͛�DbDն�.�N ���uZiw�m�o�A"D�����PV��"��f����5�������.�m�k��>lj�J8YD�����$Eۖ. h��+��t�V9��vB`='����v�9ﺃ,�t7�FA^C,����<){5��c���gDNB~�P�����C[(]�8T��bt�n��)e�Ġ��^ΤȘ�¾��R���䦍��ރ�#�6����u�8!��s�aW�U�&b�y�rA���(��K�'Ҝ�����K>�Y�;m6��x@\���D%�о>��˂r��t�@bj�+�4��ø���Z|B�/t���R��'���tpFo�6_���o@��.�����>#�V &�B��8�ڔ�@�t?��n���|-�&�#�u�
��J��j�X���
��j)a�N8���\8���etEUd]i�_Rl|uc7 7�GcC!���c��I�ŝSe �2	mBCk�\m�����b}����T�(s�^?���PD�?�Dղ�qII�V]��;��/K�7f�Mj�.��D_��}�dmIR��c�ǧ�n�R�9.�E*&�U�U�{fίd/Q�Ş�u6��� �ث�w,�LN@����@}�l���0]���ӺY�.�T�=*��O��/�0�(7y���(�T����h��g%�L]�-E��7��E���h�_fʪ�*��*���\T�ӷ��45��9rDc��
�^�&8&� ,�ޢ��_�_W�tMܘ]��zT�'y��_��Cpi^�zTBQ��{z&����B�N�'��
m/���9�k�#�Rk�[�C���Q_��|N�L����L���=4;NrW�:�[/�Ҵi<��N�lr0'Y���	����-P� �aE�M���7�/�N�'\�_x=�#�{��1�s�f�En��"��M�%q�=�v�nIbs���qɎ�E���݄�)��3-��1�:	������^��GV��Tｷ��<�poz-��S�\���<��e��p`����cԄ�<�;��J�!�n[�]�Qͫ���;�#�VbTѐ����x6��q� 
�H���e��^q N�C/t��� xl`Ujt��%.e�Lw|C�OyŨ�.v�.S���
��P+�_F��H����|AD86г�<��ɂM<����cC����~�_���ET�D)�H�a
�Y�&�)w0'g �Lh��xG���W�2��7��~�QSɁ�mEA[�m!"7�r���>��%z���0���P�5��nD�[6^Uy�Ie,�����/�8VTC��M/ҵk<�n�H�a�����j������U�Y�t��[��t��	�"�^�l�(�	�H�,Z�}8��� �lH,>�����whJ�ǚ�E���Ƿ?Tٞ��(f�d4C�E�Bl^�s�{Џ�+�搟D�2e���|�V����I|w�c�j�C�JՔ��t�fԯJ�J�NB�9��oܯ[�L��@3��è��K
���>�HT")�:I[��uD&���k]�o�ś~�-�D9/���C�Ѕ�+�;Xh���|'Z��H��}��rtl��v���}u��ۧ��Q�l��R|�=e~���n�4�୶�����gH��~Ca״,j�����{jӻBq9�V�ZVR5c.҆�_�-���f�G�8�e�e5y�S��e���s8{�eAvHS�����[X�mT�k�iT�5���(²[�]tbȌH����s��Hx��cufl������/6��y�
��*yG�&���N���l�x���ܾ>p�v=��t_$�7��f�mt]A��̂���&l�����֭R��e�5�P^��/_ ��i�
u_�`�9�11�)����QJ��$2N�j��ۑ�=�v�Q&Lm�q�5r�c��;=��Y����(k�ro*�x�=#���~��"��1�������5��TH-O�n�������j�~����L��
��Z;C5�7�
+��h䱂&�j*9�a�*p��ǟS'0���<���Q~كZ닗ȋN��v�=�DA�<�3�y�)ݴ�ŭᰛ��2��6!Ap])�'
��r-�E���0L���ܓ�)�D�e.͉"����)�r����'��o^��5$C�@��I�'�!�v����p@�������n�|ʆ��j����^
"�Av��Ԟ�����zV�KV�m��\cu��E�Mѧ���'F!A���z�L�1���4��ĭH&�:��R̌NuF�^q�ٻJ���(�_��]�����)���	AԔ�A��{�:�o�IO]�=F��FN���{��J,��Ļ���J��̰)��h]�Wi�Uu�5����t+(�|��p��Ն�=��t`�����*7�
�ύ�4G�H�4�����	K�٥�3P09ߞ�`d?����9]l����zH~� �_�׮0w��%��V���c"�X��4f�av�Ai�#�"&����كk�|]�ϲ#���o@���3(,7{{_���^�w!�5e�Q�5";�&���$F1��i����+y���wZ��7-������>`w��a�����x��lU�� �|��h���0_���:�s�V��bK�r-(m{|�x�^N(�f�}dQ�r⛤��9�>R���P��_��1�,�,Mk�������8b9o����y��}��$Z�e.IϘc�k���{r
�����8w#֪�����"	�B��l�^�,�`�Im2��T 4i��%�I��/�Q[�������x�ܙ&$��n��o���5��]�ե�W�0�uji�;��Hw�
�;�Uu�K��,���S�V���aΌZ���AT�:qY����N2��=໣:ˣ�4�{����/� WW�T�(�:�ֵ�O�t�c���v^�,����Q���SyvI�W��N�{{���K��(�EMb듊�G.��LU��f(U���̑�xF��MnQG�"v�e4j?ަ�a���Wz,k��|�Ѭ~[G��T
�)�	��cX��'�ILǦۜ��_U�Ԍ�Bs�
ckH���n
�}�6R��7����1ߺ�7Ϗ*V�_�3t���<������4��ڽ5�H=#�3�/|�>�Dh������F<� �ʮO5�c���Hb�@��Z�lƫf�>-��<���к))��ﺏ|b�Ġj�p~l%ϓBD�WzR�ڛ���l=�7���p��Z��*�¦��z���c��$�$�~2%(Yo7������ͩ^Y����>�.e�q��a7j��n���%�;`�1���Ƕ��{�wz(u��*P���^�
���N|ہ?<�W��ce1��k#��S��s�ZT��Re<�܊v\�N��n�x/�-A��9�{pF'aB�]�:���E�8��W:�-�
��q����MfWo��aؿ�Q����?�{��DY<���V�p�4RUX���,�p��������
N3R�6�xԛ]~B�R���w�i�������Hn�t�6���R�[�]ǄF�`�a�{l���i�N=$�L\��Qr�Q���$xq�]]�h��{>8]�������β��v0��#��Yn
�0��/�`sui�������!7��k��1�-��^4@+����^�Є�T�{��F(�VG�>�8%4��/me��I��]md=��B~r-8�jz	*{�kZ7┺(��:�%^���J>i���5V|�����R�fU-�Sx�7aI�W;�=������<�8�D��V2[Rz4�����b��ն�n�Ϙrނ6~F��?{��^Z��[�^�Nv5W���h�5ъ��� ��o�T�oJ !~^zs�`�e �j��ݗ��_{�\����@B���*��{��I��/I��r�;W��+�����J�4;� ߶��}y�#5 ���9v1���3G�ixڇ�:Ͷ��ڴռ�ũ�̀�y�!���o'��}%+���.�/U�}fʶՆ��C>�Jc�c��8 �t��<�Q�2���#�k#�逢�WM��k?�q��m�8oX4���V%�����Ở���hv)�Jlv��i*H�s��m�>��؉�Co��LU����.#�[�>j����^Tq
E�!v��EX~���:i�h��F�j�{*��|=ņU��U�sp`�U��n�5��m�]U�pQ���	{(ٍ�/�q�d�9�ݖguX�)Բ"l�n��BᄊT(-�W�_�xgiD�R9Ё��\�4ye�r��]�t��=Z������P\ŬW�G���o�o�fmňX]�$�?ɘ��:Z%��ja"��gU�A�Xp˭Q7q���'haJ*�E���t ި:�ZiC����=�ƿ�Y5�i0�@֧��&�Z��@:�A�������}�_Fئ<[�niò��ۗ�%"�qt��P+jp�H���Q�4��\����n���7�&_c�؀�%�+���Uhѥ��C��h4�{тĤ�~��%,H�kK�C.�H*O�mEi"dO���^�N����
�|!��'�)!p5k��glr���Ջ�	��Z(]U]�zvқ��>�^�$�m�����)�ż:>��⤁='Q��s�g+*�V���8/yaAM|��<�	���|ĘI���N���H�<y}�ߠ~L���]�(��!��=�F�^�qsg�B�:$1:�) (R�fH�c�"U}���ހ�-�*<�QV��H�H��-�uA��	�"��R5Oc���g����]y�b�7�t���������-�~ϘV�N�U^d���rNF�GWD9�mT@-e�8"XL8Զ�n�������]X4s�5��9	@��ŉmI�B���U	t��5�R�N8=�$�Џǅ�v:��Y�91��FZ��#.V7JZ��;�L��m�첑Z}
�L�]gT�������a1�>�f���x��tw=�� ��8��dX����K�P�̣S�}N;;f��E8�B7�­��_�7��l[��o�Jc�pW�Ry�a�9�4i`�l ���<ZM����k�s�8,6��u5ie�ٙe
/M^O�ŔU[硔Nj�^�����toGX�v�<�+�����mFT2���LF�t��'�m,t�����8~�.-.�)�8z�%4!�\Y��`��D��̻W�@����m_4|��	V�x�2j�M��
m�E����g�B7d�kwV|���#��:�V��R�+V�}3F�\��"��7�K�7���(/�a�q
�\<%��>vS�#K|E��H��w$���Ef��}��,� k�7ĭ��e_X4�O#�X�_=,%�Y�cA,f~�-+��U�CȑrX���>����В��#z���e}`p���}BP?���;�H�7�SR����l�9���ۭo�
���7̻����1�@]�+y������d��U�2�R#~>әI�&�ދ�;��S�	����
 Y74/�� n�8�oh�:��4�w�\��#�υ*���"v�n��.���	�M"���E�-c��4���ٵ�3C�"�IfԂ���@+n��z�=_��)w<���	V��V�WmP7����Y$!6!�:�qp�Pp��Z�D�^Y
�r�j��ƿ�A����Y�7��r2��(w���Ο���O 'x��u�+��7���sd��{��(��~%�CʑC3���l� ��D���{�!`4/P��[�qkR5x���xF83� ������䜜}���B��O�����VU�ΑO�x�NӉ�K�C2���z�'cb��uN�`�!�k�79��'�GP�e�vW��!�3=b��?Q>����c1�0�zt�BJo)R�яI�X7._LMo��ʟcl��1�t`��)����}}S8���r_\P�Sg��C6�lyߡ���,5�����4~�=سP	�e%���)�y�������J|�0�.k/��b������UX�m�m3B��"n�x�U��EG'Ns�S(��ra�kd�����Zm��Ǯ��*�]1 ���[�x�S��֕#�ǬRـy0F�_���IC{<�CuA�1>]�����E�[�4=��9���{�oh����W[j�,ޢM�;YLL�U�'�w�#�fb ��������wP���D�HA�y�Ͽ�v	��A�х���6�*������g�fH��D
�DfH���!V}�"�U.k�����OPԹ�
/:�Q�TR�)�q�a#�1/�5�w�Q����=��c�_9�>��A��c�N�����ֶ7�$��+O΂>�~�)����I~F̙��4�7��k�,�R�����6Lˀ�c�&8B�N�����`������lqC=<v�ȴ�Y�w[��b��|5<��7�N��e���e�}b�2�8�vg����u�l��`4��Gz�q�L7]�y##��o���$L��ff�W1���nF�d��G��Uw��m�`�i�^������Z�;���.�6���@�!L��Ӝ�sـr���[Zl6u4�)���k<g����UR���F�`�W7xr{�4���S�;�B+����Ô	Ӭ���p�_��,@��;n]�	+�s��t�22<��¼�#�Qh�͠$���СxKm�*��4Y�°%�X����K���eb���&N�Ҏ\T��|��X����2t�;�_ҐxA��L�XɆP.������t]��}1��$B�+<Q����s�u����q&����4�V��㑬O�0>i���/���l�ͮvN��'Z]��ng(��F��W�{_�S�s7O���\$��KЅ�9S���G�c�M,X��:��u�<3���#���;�_V�4�)΍]0$6�2���}�Qb����V�BÄ�~�=NW���|�{�a&�~B�.Kj�7�d��<<7��o[7�)ZGh������96��Eec剑ikA��lf�����R7ZD�e<�Z�*��+�?@��sf�
��G�1�e���-	���y��E�,��,E�/U�L �|����ӟ�*-ޟ���r�uK��B�Aj��W��-}�`��HP{�k�l��[��-A�����B����ǥ�/8k*���4˺_�����7�[�CΓV*�g��b9#[tL��s�Q(4ڂ��
���`e�z��D-�a�P&-�q)�J=��M�<����$lQg�49�Q4{��f6HS����"���-9�,�%	����k��~�K��m�
��W��ȓ˞B͜�E���ţ`��`Z���X/(� ���~{��΀>,	�sr6�y$'��IR�d�F��]�Q��:Gpm�2���q<�!�Jh�X=Կ��T�<���6�h���"�l���`��)��`~sG�4r��i3~�U���٘d|yq��5 Oƽ��{/����B9`$&9ǍԾu�Rmj�'].9�F#�طE�(ao''���=ܺ�7j�Э�1=���G��
P��o�i�%��ʑ�͐�����Ŏ[�"M%#�K�:�K���N�y�Q�'-Q㝕��v6����x�ˈ���b������/�ZV��o�7{^2K�
�O7��qC�M��Mh��U/ZU�ݑv.������L��4]�I4����3��e��g��F� *@ڽ��!]y��9�a���5B?l�Զ�m�ycV�/6Z1���!�"9�E[���܆����Z��0�7Y��i�<S�D-�v���WPyy픀����U*7��S����E����	����<��y6�$l�<w���)�Vzخw�0��3&
�k.oC_f�>�Pl\�qU5��6��DʯJ�*���aM􈅸��m�'���C��3&ky^���E��0xل¿�����L�6}�ވޛ��v�y�/���-��VD
�PsJ�Y@Kmn&+�� �TK?rS��G��QQB˫�z����m��+�4�?�s�SX�}Ih>I��c���A�ø1W����Fe�h�Qk��^���o�5��ܛJG����#�|�	.��_�7�f�S�"�Wz��M3�:{ݪMD�0�I<y�5K� T�#��C�&�
��UV�Rr��#\<<�˳t�y����=�S����DǗe��i"��|����e��@xMy��ٿ�͹hjbSyCf�d����ZoZ:JN]�M|���!e�8Y~��;L��xӱ�R���L����m@��^�ܤ�����i<mZ��E�m�)�]:8�c�"�&)��1����P���{��.浖ަ�L�%el���X2I�f@�5	�g��WVA�c�=�Z׍{��7�	�mZW�BK�ݨ#(��I�~b�.'��f}�9�O����j�v���(8ܾ]U��Q����2i,{":j��^�_�c�u.�k��;J��n�Y�6��{K208�����ܻBF����+;ZC�ì�RϏcZ���"
I���I��;�Yͫ�����z��f����E�Xo$�m�d�<mcyWI�Q"p�$�T��������7M��7*!s�:Ͷ�0�p�������;Db���J'���Ј�OM��u��ԛeX��7�ǎ��BC3	�ڊ5�D��%ݍ� c/&�Ǥ츦��J2>f����&i�q��!���̀��=��*���W�������*�{_by��!8�$�ޏ��U=b��2l:PHJ,�������i�]?[QdGV��Yp�`��]CN��R-os�r�����5}���bQ��-$Xћt�͕����A��/Eu��UkΘ�O����������0�H !ʍ  �h��_�̘K�oG�je����(�eJվ�DB�zK(5)�ڏ���b�%�xuv��&s<���u0Jƺ������`%�ؔ��'$��^Ƥ����g�|�G�ZzԱҔ��נ��K-��� QW=��;��h)@��A����;[�ȃ���2�qT�H<v�@Eds��L2�x��%,��T-��t��y0��<�.��.����<P�=���1O������kW� ��2y�SN8+�؛P�"y�kبh�)�SH��n�&�*��3�'B{�h^����jJG�V*@�w�@��?�wW��BM� ����q��c�!g�m����|q��&0���4�Qx2�M���bן�;��%MȲW�vQv�)�>T�h�OÄJ�~�o]O���u�MD���}�7.E�vX�@dk�r�]�\��G��v�H�c1��b�X&�<6�#/*K�$u���ʇ��3M��`��^���ϟtM�U4�x�7�zLP ��[�a s)�(����gp�tk 5U���W)�3m��nŰ�0d(8�YhB?�#�?�W�K�G�	W���G���Q��Rܶ�nm9�OiA����p�@�X���7WX+�L*r��3-B��/ױN�_�S���y<Wf��PQ��&�R�j�dz��XoLN��	�u�Og�)?Ҩ{e�!�\@�����DM��g#*(m�����y�?%��=��o�G�/w:�[�Z%amn�؃b��L��t�[:+S�ƢO^)(cкn�y+h�-3������U�B�gN��O~�!��a�b�� Q�g�q�;3x�a�ZJ��E�!V�q��"m�yɦ���Α<=Q�CE�w��'�!���4�� 0b����R%CCh��3�K��=TU��	��!a�@ԃ��)��-�u��5OB+l�+A[���T_ly�9�>��dH�'�G��ܑaxF�x�C��T��<�F��7S���w��8?�%�z�g�9���!	!U�p�7�>�w>cː	.��x���#�_�tnC{�"Ga�W&�`�n��Ź=p7ۋM���]+L=�w`�r>��>t�T�� �+g8����`�)���]@dy*�'�P���C~�?����Y�G��7}l1l��~�Z��#H��R%Di���hOw
�_�ڀ�_\�"��%웭i�y}��L�y�K�ۺo{U����/�:�Z%e�vA�;j����8�pȅ��0�K�E�2����j��C^�KS�	D5�n����o�ڸz`먘����&�0x&�cݍ�W� Ku5��ƗV0\����ESԻWU�6��6vq�FQY>�,�J��x�P�}>�n/��zO��WYʖVuܠ0q����Q2�9�Z�W�%�+���.J�ʲG+T�#� ���e����У���?T�V��x�Z�jS)܁N�,v�@<�� ��ia��j���s��19O�ﭺ�^�eI����~���5Pf�LL�7� �#N
�2�&���p�������"�V���Y��Ĵ���H���5�k�R�~H����n-<7���.N펅�c�t��3�OVkJ��I
�
נ	�j~`���M������~	KW�f:4"�al�}���j�3�����Ζ�{n�"\n�.A���G��j����j�x��u�;f���c���q��TͯK���3՚ylv�x��֐qerA���*] �|>�:F?і�����+i˒�o;��u����L$y^+d��wOP�7"
��&�sS�Vˠ$�q,͝ϗ��r~K1����lﴹ��S.ץ%����;�RN��BOɃ����(�Xi��� ha�U<�lV-+m��R ��CF�d�Gq��ղQm���!w���R�O�4=w���؋�s���{^���3��ɞ�����<N���d��N�4_�u%��j�a�p�$6��pH�0��T��U �Z���a�l�P�[R�c?_�A�~�u��#���u�Y�}9�	+�Z��8	�4s�;��g�L�
��k�_�:Fx�8I���D�k�E:�ܟ2��'V���������׎�G��4c�Y܏-ov(������j�`i>�P޴�lc�M��O�`Ҟ������c����gw��ܾv�2m�:k�2���� �|��A5����M��F$���}���_]���E���0IEu�0��j�m#� Сa�x�=i��<�F�;���A��u�ea������Y����i���6��\K���ԮC\����_{A��*�d�\&9�eK�?օ��>>���ۙ�/�$yIR����>{�� �
$��vf
�G�5�ՐIl!�<�x xR�v�ҧè�N�J����LB�y�L��{��Q��y�(�(� U�����^s�k�X���G�c���`�V���{rd�f���Z�_�&�Tw.* Z���+w~�@���g`�'{�p�#FU|L��(�L��*��T")�K5B!�L��,�:P2�d.���<k6�!@�^X�b�g/��u�|�<����VS�l�=�kG|�T�BD䏰
N�=�Z��0�7v 2��}K��_\�a��oَҎ��7��0��?554F���	S�]5k�P�w�04uJ��C�CV�w����4�$E�U����׏�e2�->8�y]#��+�-�dD���W���'o�d�N�Y��G�9g>�y�
�A��[	��$�~	S��)ĺG&%�T�x��`�^�ʪ#��Cd���Bu���)�^���W��]n���'�5�{�p�MF�d�I�g8�p5	k�W�u����t���n݉���ص̀I�ɔ�bG�P�R��/���uFA��&&Z� J��>��2�'��n��	b��z�/���C��kG�؈�7�����=dX̱%�p�k�/�ێ��	��nNå�R�N0��}����a���-�L�|><����8��p� �*ZQȡ,>u��mK�8�|R��i��<~@��&���Ӑ(��Ŕ��0~��]����?�C�v]�	�x̬�i�����\��=����ǔLH@�OV�����p�)�0�䖕�o���E��� eI[�_���pmu�6���!s���b��X���C�4���5/0Uǀ��t�?xRy� �m}޽>���?�ݙ�`���l.v�D��K�RW"i~Yn��=�ˣ#A�Yp�?�� �{1�.�}�x)��C(SG��Y^�5OBҍ��
-��i�p)N�m�5{r���� �H=���D��1,���2����W}���t����}�E��d,�L��#��2���R��J�p��X�3C���٣]��y`�7�t�ǽ~S��&���n]�v�=�C��ܠ�	=E�����D�*%/���╥�DOA��3�Ԙ│�3�h�L�h�a�6�,Ul��^���ev�nF͋�����C�?�k����$�Z�1�'x��We��w�@��MT����gz��1e��E�U�>�,���
]��s�5���2�@����R�P���<�P��Ҿ�S�3�\ֱ��l�y��g6/8T��ן%y�`���j�e) �%5N�l��6�*�UNc��"�V (�������o��ވ�pݿ��!K�����d��@��-_b9T�duHr�M�������c�� �?���_s�Xr��r'D} �l;�Y�\*��V���W��οM�,��p�u� ���~�G��(�a�V
P&Z�B���{���+:G\S�m�
8�ǋ���q�/	��N�E��5'����_w��o&|)���b���}�mN���*�P���[�=Px4���.��#Mp���V�L�N$��Zm*Y[���"�!7�tej��;��F�.��ڳ�3�CY�ݘ��t�*�x7mg5����s��?�b|R��s�.�4���2C��y��ؘiס��q�E�gu%�hX�)�ǟ�[4)��}-M���5���۳�J�����v���d��D�4Z���`�B�	7��)o�D#e�O]��Y~��+o�Gy��6���"֛@2!�I)>S�3r�r|-0yT cB��b*�涹a�_r��<h2�|)`ߧ��c�Bmqg6"Q��:N��W��n��ط�2���8�p�������BC�J� ۖᜩwuVS�)��;�(�6�r[*<_=y	��w����]��u�Ia7M�w�xBۋ�HI��<��<F>Uu�Q5٭¾����]51-75\�vj��3]�����Bۨoֈ�i���&1�9�dЋȅ�ME����WOH���>'x�t�q����D3.�6zJ���h���F�>��&���;��@��b�uzG`-^��������� �<6�4ś�����pH�������;������(2�E4%���A��6�*�$V�c1<o�={�@�$�شK ���&l�`�L�������T�9�mh2q���-s��V��n�91gK����S�<���
�[t�Ã.�~�~m��N�mh�Q��m�C�����P���V�c<��
�Ν�tTYjq���@���xEy����)���XA����z���r�z���P!�O�,��Ä�����������|)�?��r�H)��*hk�m�2�"�}ʅ��h/�}r\{\����+���"I~�V������$��J	���j�y�zNKxQ>�,�^ip�v���e���h��}�� ��~�����qe����':�d-��lM}^�q$-�{��Bo�����-�~FM��K�}�B����E����~����ަ��|nT��9�iU*cie���XH�y*�#}�#�����n���˯)c�Q�=�'6�aH����`�R�21�~=������]��6�����E�O��H!��m�ߴ���������.!�+Ny��/|㬷T��ҸB����{Z����X"��ε&<��_Ȋ�ШXc�s����dǱ�C�x�1Z�(�E����ht=g=+y�)�%�M`'�A�f�/�R���@|�`ib����?C��zw^�'Z�oW�1��R���qQv1,r����lm�5����Duw���T_��i ����
�����⋠��	��vQ�'�o��}jv�MZkh����"1֦8���td#C�@���J6L�A{u���N��)+��e�2���!FX��T������g����$�J#�۲4(�3��=G�^�nE,p9e��)ZĆԛ���Ƨ�[�+�u��p2y`�_��L�B��{U�خ��^SKz9j@��Sz����˜;ల���P�c&�@1$�CMr�W�j�^FIg�7~Gق���	5�Ʌ���>A?|4�8~V�VB;3��P�9�B�F���B���n<�@d&��'�d��1���;M��r�z��V9ǰWu�zx٫7�wM��D��z�)c�w: (���H�_CwZ�g���a�ѵJ@��zY7&J�=<gN���&�|N㐬3�����>MD���!3�}ھ��O$�,��S�p�<�����d�J��Ag�,6�eT��.���#�,^��u;��2�A��3rϩ��Z'�y�� C�Q������ȇm4]ڽ����ɲ���_�N_��GW��do�F��])WB�51�NGE�qC{�X�0���v�d�
��m�������,�ˢ�Q��?/D��8��2T�f�ҭ�#Kg<���[,�)j�Cø����-Դ�@�J�_�e���������!���ĳ"�e,�������s���P3L!�ɡ������gK�H���7��r�ʕ��S��J��d����@�Ĩf�N�R�{��ׂي����5����oԃlU����cǞ
�˭�D���� V*w�����ġ0
�ȐS�0��E�m����\����!��_��囿��y;W�b�:�I�F�+����{�X�4�!�oJ���;��z8����Q�r<��q���#a�w�װ#B��c����U��,���Mh�Ⱁf��C�P|��9�����Wt�8�!R�q��p9��g2�0k5��֝�P��~��a2�)<9�n/$�4�8aYu��~|�8���n�1�!��>���n��|S ��� ����ɀ��չ�I���@ǐ�d�2����hRD�0�te=��H05�|a
z�\.)Mm�`�����
�eն�H�z��{h/��b�F�ٝBsa@r��4�+�L�·���9�G?Y�c��wzY̛7~���3D�qϓM(�bU��~�$��J�Ҍ�Z	!����ns#��^�r���)�~ ����B���!=q�[m�UW�q�N@+�t�\ϪKO�V����Y��ܼS���ߴf�~k�S��l+SD1̟��~i;�TTؗ�a�| �0c�B��>lxјq{TJ���d)�����a_��ެ��3�Ӥ��.�X��	���р�`"d�`���}J�}唩���kaMD;D�YƓ���(`ZT��=)\},#���5�$+��h�|r�#�P�+��jmx��EH��������t�������h�Q�<�dˤe;�|W����ļ�ٔ8�9���I7�5�D��'�S�&5��}=���T�Sl�� ��W�{���Van�I3Y��%���p�U�q��l�H�3��#E�����dݟJvx��۹�n~���rU!8I�c�0�g<3��H>pC�6�ŉ���b�s�8� G�������xZ�������%]R��!�k)����N�s\��El<��rƮ�iO��wZ�d�DҶ�H(��	3�>7[��O��k��.�O�_ᗈ<f�9\�56���gV�����\	 
-��vI0�w�h%h5����g�q��W���4���qNf+R�e�߀��gD�9s�T/��P<8N���F��ItDJ#�)<�B�}�i����,�î$�,���sl�������E���zA\:&e8��I��h�߻k�;�I5�ߎ@Hбf3G�V����NN�������ޏ��NR�Z���S�m��fŎ̢�ĚL�]˼�,�M���$b�u<cUG�����{"�'� i���k�8���F�-��"Q�Ko7�|�?��S��g��}BI�%.58�'a�~���38�r�c!�_ڛS�Xq��U=/l)D�E��/�یS��L3�L{��S�ţ	�4�H��5vJ\��J��=$���H��#�b�����)|�bp+�i �2?��#o*OL3�x}�};�3lc���&��?i=8�
G�eD��*��6?�P���HcI�&۾o��h���6��iI\�P�w�nP�4&ް�9�.j�r���	�+����S%������5lF����\h��tDٶ�5�-D&ko�l�����P�9W�k.� Ṵ̊����`�mh�s��S�]��O�(k}.ސ%!�5?�d,[x�r�-�$&�����D>yQ�MNkwP�WmQ��=�BF�<��c�5��>��?^w&�+�d�h2�\L�[�r��@�"�Nw"A�vO3��t$̦�x�B2`�ZkU��$�$)�����TkmQYq����Ә���ꅞO)��7*b��@�B�KT���\�iD=�b,�&S�� 0V�܁MI��f�����iCD�*yq���a1��=���T�?��A��2��!t��_3{	ŬQ�m�����җ����e�ɒg7�a�9~������K��N�O��W���{H�v�eL��
�u��� ̃#\(���=��xgU���SC�n��~��w���ңn�j��?Zf��3�4N[׼���7�RXt�{�T`C3�zON�� �I��a^br���u���S�\�R�e�#2m���ۖ��S�i�i���,�^"���d��jvaU�E`,�Q�<��"��ba��Rٰ����3���|� �#B�I�s�����V]�X7l*`.'v�2�H���*\�k6�[�}߻і������q��=q�����B�k������j������t�zI��%]ȳ��*�pw�z^��9^
R2'���;�V�o���X<xoM���ō�.��L�78�����l�8���HpФ7���
��s�H�� H�bɈ���;��.)pEgt=RU6v:l�$� ���M*H��?t_�QO�s� ²���t$�{�����YKX�D�y?��m4��S�HJ06����欦�U~�l��*�����Buu�`�?މ������%&�����$*��c�̂pH�A��һ�񹪛j��������S��i�CA$L��pk�\jw�;���cR���M<fF���X$F�3|Ϛ�|��������o(�Q�.��Q��q{�M�dD�A/ML1�w4��Yc�U�iD��yNY0��z���#����Ʃя7��B���_���~Y�y��Z�\��Ju�OJ�<�O�Oy׉"���#�=�t�?1�V)�q�Opd������4��,���԰N��a�Sr�9��i�sGPc�{5��Hn����g&���:D�)Ј0Z�e��J�R"��I4ٕ~����$Nm|z�P�͝+�$֒�Cڔ/��ú���`�޻-�\%i��T��Q��H�Z��K'���W��H��Þ��w�¯�>]Rp�4LQy,���,�O6�.�J&ʅ�e+�=fAn����x$�8�>��*���dKo�^9��r����:ȅ�G��UƦF����Ƃ�D������5>;���K�.�ѡL��n�_􀑂)��aLyWViV>���2����p/G/�F]{63k0W
�sU�"i`����fyG4��;�x�ANA���+z���D��YEM���^S�/�Q�fV�������mX���&@-L����}乓"�&�i �l#5@8�μ!x]���D�q]�k���ъ΃&��-j6��/L����x�P��J�LBC���1�اf��?(�yy�����zS�儥�GJMIϖt�\�������b�L�+���+;8�r!L�*�5����Z��u���j�G+{,,�J+Q��ٗ�WN��^B��?���q4��V݉���p=$A$�5�4�8^�?${:�2�5�^,9�g��[*���a�g�(0f�)s��B�����H5��|�G�K��E���kش�ۢ)����I&Q���d�b�3LD>v�gY��7�=)��6A�{
$�^ڴ�cQ��gU����:������!�$�ً�J�<E	"	�z��/r~��<Y˲}�hL�K��K���MwB萦��ܦSs�B���m-�Ҕl��2Gud���Mm�-%@��e�o�m�� ���+���a�P�!���:B�k���j��	��p�̕�z�Y�@Ys�xQVt�]���ubJB��4�`2+�Ns
ak>Jx�6�1֤!q:AksF�L!���Ok�
e���V��q���Mv0�g<���@��u�,����� �Ȟ�qԘ��sD��T08�L�W,�봽�S�D�PJ{�w	p��6{�����I$����$W�aߓ���m��n�l�7��V�U�P�&Ӻ�H�R"����ق�^@�WR�K�`>�fZ�%����#�"D�>�
1q�br�>��?`��z,n��ݫ*��O�y6�ʹ%ie��2��&|��32����j0�!�����?�H�g�'�xB��\6�LQTK��`7�!��_(�0�\,u���\�B�+R=�eM9y7�ĦE���2M���;��A�O��������+��V�J��}� �����dn�-����qp���Rw�k���ƪZ�ب�fm�ϖ�x�m�A9ȋ��n�~9W4`]/��R�N_�ϓW�M�0��v@���J�L�zz�^�¾D�!	�![���z���AEɱ1�Kr���W��B��t��>;�`���gWЮ�A�
�Oɉ� +�5�`�\FR�1�
Ɨڗ �~��qi��U�'�� t}�hE�Rg���	��[��Ƿ1x��a���;��PW",��,�hz9��4p���H��26�o�	��S5xz0��P�ZW�Vo��)z����T��k�x���#�?��)Kr�5E���r�am�jRl�Z*��m�jΘ��Xd���t��\"��_#�V��S1����!�b_�o1XQ]3�k�@�-��9��a��b�/����ɹS5ь+/?$o_ӏ#;̄�_ӫ��&�����L�_0_�yz����+��� �ܗ�U��x�ǘd6������k����B�u<8ס�Ĥ�w_��NLDw`gʞ���W�I�29��?��HX}�K��-V�q�#�����M�pҁ�׉�yӅ Ar�Sq�"��]�kPjt�=�ѝ�"�Yf$E�q��} d�`T�a��U���K���A2t�����j���b܌�g��G��P�R��c	�"�\��	(��v�q0A�Lg��P۵k36
dӠvє!$j����F���G
ݭ�Zޥ"ʊ:�A��h[
1k����6f����'~�Ѭ��=�0Vp�`��n��w�FY㸾.�͟���[��H�?t��Դ=,N�ЛrJ0b�I���2���[�m��}�][����*)�Y��u���ܨ�?
�Ys������8��O�� �b	�wk��S�RnV��,�A#�Vr�{y	v�dQ\������x\��VHqj�l��o V��.�ɨ���	��� ��l��8��.�S2t
�{�����,&G���ѽP��b���[�)��NҶz`A��33u�G�?��z�vxJ�,����*ʽ�~��E�k����f 
9G*	�%� q�sA���Ч��~-�D6�\>��
;UKGv�ts������ �uw�%F�_ӛ�}K�D�@�Vw��\K���e��������Wa��=�C��������&�FZUq�6A߸��-��iQ��r|����M`��)`P"�lF��m
���J��M�T@au�"e�J���Y�f�k� �$J2��j�{Vj���������v�8��-K�rՎ�c�8!���9~1�K%COM�eq�%v��hgKɳ���q�H5����^�ˉ�A���G�_��\'��'�)=C�Q!�0M�h�CAʶ�5{oa��p��9Dbɲ���}gXΦ�)H��o�M<�\��3"�4O@�t �=�~V]6ϓ0/)�;̆Q�8j�8a��V���~ӿQ��a��5�����$�9ةRF߷mc�Na�����f�B���2��w����Xa$9@Ȗ� ��E	H�}�m�c�H'�+�gԿ?�����Z��S����4��[\>��3R�?.]����3+�?/,@����Z�U�0v�;�������H�vV�ͫ�ؘ�:����ԣJ�Y~l�|�I���Ey*g9M�)�=��������ˤ����J�7�kȝfR�싟�	�h� Y��S�H�V�ƻh�dJ���Pb��dQ1d�vc�Ԫ��*G��Ѩ���"T-��;8[�����zm�6t�O�t� j���u���M)�u{�j���*l�8ݭ�L����J�k��h��U9zPB+fR����&}�DjA���0��J��
~���R}���Ǳg�/)V{{ɋ]$|e��*zz��z��-`DG���q���UĮ��`,�.�ꕢ���nX���G	��a8����klY(Q�K}���Pc{I�5!��53�I�u���/(���.�HK9���	����Νϴ��^�ąƩ7�YF�M6x����Аc�婣�q7�M��T�Ҽ��^N3��rg��[��*�D�GIw�&.o;B�됗�p_|�`���b�U���w2��x��o�ar�-I��8�~�VL�O�ފ���|]��X����⸼s��8;�r�|;�klR��P���2�.%�dt|q�";��u�������܇.d�����0O\#u�z�ֱкW� /^�8�t�(z�gg:X?L�e���X�w��=��wF�;�����s*`�ɇ��ϖ�1=s4������	� 	���J����Ռ����UH�͜�v��+�z�����
q=�G���k,��t�P�e7��WNA ��נZ�L������.5R�
l��r�E������Q��f�uZ�z�(-����1��1$��U}AL�E�tLI*� Tv�G�⨻���0u�ҫ�s��� Ģ���X�����!���P����x�"�w{��` TO�ˏXyu�[\=��I�a5͢p�wPߕҊxy��s�m���0�1�o��1)��b���{l�j����pꅭ]�_A�O�d�Q<H	�A�1�ب��7��6J����8�M�#&���p��K��� nST�#�D�UcX�pw*���� UA����1�NN���LtJ� �:8����}��r��+6��s��(�4�ܬL��*ӨQ�^�,���( t;�=KHEd�ʱ)��f/�5��͏�$�J+9�kd߻3\?�T�*OT�!ѐ�]��z�8o\7����~dJD7�ݕ��	g�S�A��{ϴT����7a<%L�r��H�I��Z��E���e�J����JЎ��H��ZJ�e��Q}dy�L+r:�������+�]�`dN�@�C-�,)�헿.oY	ǰէ7���x�p7���^���Q�XD�#m�\��~ᗭT@�� �w.>Y,�z:FO�Z��F�wވ�%�q��ʸ�m$a��ߜ�%����3��h|�� �¥�м�K��	ʦ��Y�}_����g;����S7��}�h�D�<�d���#?[L���kٴ��j��3��^���Xm�g�E �>Eܼ�VMX�̖��,�(�n�|�5��A2���zU,=d���`i�Ix���4;��(/U�՗Zݴ��!B�$�����v��o=�VV�ƿ55U��m����Z��i_\��Bm�{Z��NT`��P 4�p�~��C@",lZ*SrM�05A=��!�;4����+��[�NFΫ�4��Q��2��_�V�U�UW+�L�}m�8o��=M73�OD�1v�3��m<l�Rd�۬�㍏����|n��<�J��*����QOD���M~Aƪ��K���0� 5��ŭJ�u�X�Tw��ēX�C������{�sD�J�9��)ш�e�!��sJisT�y�����sijD�K�J}�j�x���x]U��'Z#;#�!�dPr$�6_����L�X�]m�v�a��]'r�y�~7�;$�^t�6��7�A��֢�_!����Ya¼]�d�14���k�"8�Wx�9�\k��dHX��XU�<��T�1F�4x"
�Zy��B�B�d����cm+��|�U��2!�!�f �+�P-u1��W�r�V�`�Q23�P��Z\C����z9(��v'��:�t۟62� r������ ����6���-��H�l��Y;�>}��B�5n�g޶[�A���l��A�2������D�L6����Q���aq����O�C0U�$�8�9��
�}Ẃ	�@A�sn�°N 3��K��,N�ٜ��J�-���]����
�������C��H/sp\e��*�������.�>�ILL����	�A�n��qb'�`-����[�uYƫ������ i������x�б���)"V����ΤC���������	�:�/��{����g�\XYL;��4(UϹ�����ӂ�<Nj����RF����I����������ӳ�ِ�	�/����������z:�ʴ�Fʐ�=��9����Ok ��CΦ۴֣3V�����~۽'�+^��y�8��ۥ�|�:���aʲ�L��$@��ZK��4��*��#3Ch���v��>��<�$K�cvAǿ���'���<;��dLOF����0��,�*6�����*���wզTl�ѽH�P�&_��=f ���x�Dw�o�E�D44J�WPp����E�9`�E�2B����\ɰɖ���)?��2گ�lZ0���me)y��=��j���R��(�FN���������s�y�D�U�V{��'W⎴DrTL�A�7mG��	Cgi	暖=���G��8�.\.�P'v��$>��M�e��J�z�Ե�f�(�v"�Ic����a�L�������|��bkKϔ�����"�Oʠ۲��.�$�2ì�v� �W���(�i�7'��RG����&�������S�-��L�:VȤg�3����s��fV�$a.n۫7�S���c2�g��X����o�%��;.��Ԥ�8K�*���� )��x���Y�rl�i"�N��4~qMx����j�%o�*���E��Z�