// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:55 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
YbXkvDPHXZVlaGyEfvBNatlhJfwh28xdGqY3qtPplPoQG+BAAvSXJTh48b39heRx
3xWuzAJkRa7OgPSnIjtUqenszIWrqbbif39Zf3Wwzn4IvEpxlLUpvPubLu/wOgxo
zss1d+xyOoPfucrAtF1S+GPII6rY+/Y6mZyLM6d9uGM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4112)
jHBxm9KIyGbrzW+14wsDdIEK5krIik80TBOZ4beTK8Z6DtYIBKt7Q/laK0rEQ4dJ
KtUdYUJJwg5AHQk1cRyov5l7y4nq5fShatWWzS4rpcjASFbZWDfw3jjl49OGiknG
gYd/DBy4zx+Or32nXRtdISUttSZwufsBXvQGGwQOneE8irHfMTepyBPSlxEcq2Wa
DPl8WSP+H/E6HXxE2vYelUOFkeDx/gyCGQu2NNir88WULhyqGK6OwyqkvnDbRmyM
G1gOmcKvVoVLPS+/oeAbmlvD9rs6JI/t07KulVeDiEILwOrdrsuB4sdkEnNxmHit
VglKLfg2E5Q/ispYl0T9d55n++wQnkHnhQnljSrMhRc/U+a0NvU7JjC2SavFeqPY
riRrYQ1rcOkVekSWwUBEhf3+ixOCAbFYLjh2Txik6Nf706nGmTmv4wg/N1/SdiUO
RhkWmjLXp9I4raQ9+btLnisH63xGtobnyuz3nD53hRA1t3jEiNEhKQ9gjQK8Wk1j
eaj58WZF5T68zM0Ndb5l6lPCjLDgd/J2GZ86u6PqDwvNX0fV5YkJisVau98k9Kq6
2IDmYh6fY8g06xpHia4hy42hSdPzrESrVBQBHCADJR4JvP9DU3ZA8lwInEJHo1ng
E7P85icY1z+jqCJuXEWBNxoeUsmUQsZLUkL386BjxQObyoF9zmo8I29D4hraM3wi
ysGRs4z0ZixR+PcTPYQgWTFRVOLP35ZJ1nRiVFmYoR8lZAZKQoG/1ykQf9JX/ax5
jna5eBvggviHPAs/E6aYCJnPXsPfxM2F5NA2ql07WeXwG17cchFDSqYMWKrZ0Wtp
ilovVOKI/dHB+cf19wS2iTnJZWATnt0EbE4gT/azDP9qvp0igE3vT7rkLqvfd7/N
hF67g8kIypqdSdsFQ2zYSphjOJgBKPKhRa6KsuGnKJNIuBQbU6QEMoeo+yHsaOAJ
QuTQsrBn7CFOxMkkDqlTwFK/k4VVP9IllIeoPi+Lhdcek+ESC/+RhT6pQHGX+K68
nedSbOQhSBegFGGT+b01VnbC7N0z4jBhzg3c2pGQh970Vn2qWPumYAdPfafcOFTc
MEteql/0z+PU3AQKK4/3+aHUr8CdaH83mLkMNlOiG/Zv4Bp9pEnVhWtU4nkeY99d
FkteYd7rgQ34/CjBo8fdHUaWC+SSI82dadqLIT1BadjMuwsLRg/SiBf9tf6PMiVd
tyq2xlG2d3JX1J7mN2VCSk+Ye3h97jlnbPl2JsdzdP4mwgLkhv8YiWTQLRPDY2nf
0EsKNIfVi7SE1/wz7xVZsYTMRKbju3CZEI6F/9bQq2Ajb4m4fVuLQ1AW+wloYitJ
ZDGS2RFuxAl3OEHtJN1hIstKB3IgQp4oIRUD9AskOf2hdcBZ4zksfxqlueOE/4bg
NLBmA5Uefv/UVX8STqcIWy9nhhuLder1QRM0fIQXveWArnG9oS/wJakCcRMHuHg2
bt7gn1QzgK03MEwkvlqHAkE6EpPPkOmVn0tnk0h2WxvA97oxASm20NOkC6iVYFbx
1fYcHdf/2kBjuw5uUz+R9GdDGEIsMS3QqQ+rJmd1qSaIz8VuSksCij1T8E41kB3U
R6QvOzgEksicxir5lakOOHY8sCFDUHBfLGSF9ywF3uyD34WLLM1fsz2JENnMX6i/
WTbW5Cr+eEo6qoevc/MrrUT6Oju9/zFb0AfcsraIi+7+sHOsQOfq4eQpamxRu2KB
oSvYrrAna4Z//k7HZvzWZFinl0nuCGIZk4pnSgLblCRnubhuPABaMBMthotm3qW2
8k50KSFgNhYvTDd1hKRLItXrdO16lJtTLVmIJIZxpITc57C9Z8TjMxpV9Vq0Ziv5
BORMw3EOd/D1uKpleKPUVI3U7EJQCJOB2QxS/GW6a0MI3ERKtgtVW5Wz28gcOxgS
Q913gR3vnWgnTNO+KGRisXjyiKjS/BLSEgd7oA+JNFVQ6JEWKBksRNjZT7iKNtcQ
IDGa8JqL8K+8z1Op3n2l1j2DXDnNdrKb9ud+TRUAzySljx+PXqLA+4OVjfVOvzMv
jpFHljHjl6sRGzBylPKIKPPMXqFy+aDE8LEGJhDqJWbRuSV609e1QZLHpWs5git1
+3WBg85RI2aF8yc+Gw2dgoU53irsR1r/GGiKMNPRigWDkgGmWFcuEjH/E2wu1XFi
0i2tcysipYu8mRjBpBoV/tQQV0EKBXmkCV+9rvWhB9/uu+y9JY2PJtxg+KyT+mKH
dg/rJk7BrVJYm6p1lqdxsvK0CyxraQOCBc1MNWcJz2SeCvXj3KS5oIUHFHRWBukb
G5HQIvDloHT++6sESb4TWeeZKKM/tl4D+16qvHuKSo2HT/ONgJRcPeFLQNTjnu3S
5M4rSzJneEBf9GZfhJ2Nsego+A6PhKDg0SW0+DHExKowAVI8h8rPWXRDJj51Yejl
32OsqEVRxLd6yxCdvPOu6hMGbwGQzz9VPMDzdTFuafJ65Ay02iROFgkGnjUyMLWl
FbAFg4Nh5w5LCGM8VEgW8uVsMOxgEK1E7NxXCZINj6UwfWIVYp36Q/y/OfHoC7Ol
cbtyR5hFkW8Ufnk/7SLrGCiwPPLJd7Z5cJzaHvjU3VROm/OHmHbLPNgIr3qTH5P7
4KD+x7J90cD1sSs3WFOSTuVRsyqWyn1QEWAyIIwmJFXt5JCBuAYp4wlvo+fsAJj1
XQ09nGkX/GAEc8DwsJ/YAphjzXXVBRIOTN/97J7vu7HUsgO2wkWhXQfyvPVnHxaa
bx/XycMz3zctq0G5c/WUjZvYp9wGkPL5sE9hySnz2C6Rz58imSAD5t3dUvek+06W
gWrxzrJVIZ5yQ9RklXxTYflpPxSM6jCbhLlM3iMM0Wi7DDYhEHSDLYmGpstRAVFo
C2jWr5Bcg48vrgFrUaigB4aZmqJ8UnbDUec2cuN1ibof6hQ9OnuXRkBSJAP2eTk4
sFHOl2SxHyuJ253+vXDHxmV2xCdIOqLY9QW3mY3g+JY0NwHBJM3RunmsnKX3Ljma
fEV4X13zELF4CaXVuFoef6fRXS42dqqesLuL7nclxqB3pXw5fg9c53E6m1LnjHxn
tJw1LI0DtzsBdR39J5m8uIdEWRhEEls2r7Q5Ab8v+3uqeJGS568oVQFzSTbUFCMO
h5rIQ0uoKRWkeyY/BmdXlutT93bp7y7vbKRGywC/5Jh+6aEda3fGI0dFBqxVXrPi
Uw3Yt0KvQuKMqi23p3AB8CchdlX2fgqWiCY2Xv/EFMYN2wm/d47rrYtqJTcUPu9g
PHA4q/+5hpAO6i9fJCPNt0GxFdJP0YkPLOaTUg4RTae9oOeWoytAZLSK439X5aa9
A+MbziNi49K4t9Mg11Go+Wpm60DTKnfJSlQRCI4H9E25lQdUEnECSA/j4S+qG2dN
Nb4vx6UMGUqyuou6mXmXMYNdFpgyTuSkNmsoa0nY/Z2ba53Q1jAYorp581ynlaI9
z8frrfh8+pc4TfHOtuY9z7ZWNdSQ5kRiTzcE3zPTpLo2T45GIrz0rA8UVH6tacvL
tKa6bJwbIF4b/ALIpa2ZI10IAbAu8Fz4JzUdr+jCmHJpcq5uxWCKIXZs2W34mqVu
ID3w1FFyqmOgy+N3nmVxqFkDM8RJp6OownCC3xtifWu0OaBIUrwBi+tvi9/1HsGu
tki5rZ6nZKwL9WtFkDDBxWM7Qhi+6gdakWkh3cPbUWjtZl4+qzpgmxof6jyfuPCQ
vBrB4Nn6qOkDaWjzASFqxUBsk1Kazvvq8uYZwooYZGxSycMkLMa89RNbEmakWYzb
AiQt7+PAcQchEcByPUqbXR6L4x2xs6tIw5ROTqrWk5rOw28O3QnsZ9djcOVBEStt
PbN8o1/JL7a7iF3z3XNccKkQsKdKy3TjE98VsRgqMW3+YIqUDzZeNfIhqRoGgzig
cHMHkMlYEKMGyWKYpzfpY88gi7Cmouej7yZEwwDYkZtKZZYKm51W7+j9jJG4WNIH
8uItTRMsthBaHfwwJ92clXJiyITVv74b3aaifeRqD6SD58sksKvELRWZdca92jbv
OVmqrY/eIfcXktg+PvafqXoY7O3LjFD3xTgRNlsMjGM61VBeotg1l0TS/I249nNf
L+HhMHCEuiC01cTnqXADBDeRKyGl5UNLoJ+N8zdp6gF7OLJ6ungUMrmC9iRbqAxT
H99OO6TcT4rkdHwuMQW1Jlldb5+jWAno8+8mzfSW9V+JDiEuWwseKwlY6tNLfUXD
nqLHTk5aX1hyTDNzRVHTiEZHB6NNzqzJkhG+59ERWcSArPIZ3H1edmuvK5xFb/jR
H2rHGjIgssds2v6euRNVwutgU/23D3HMiGPOdyHaDOgis7RjmXE26bDuA1lCh4nc
HBDKNNmkejnkbFiZNH0vBotuVbbkfVRhtANU08oTUnCOBj6gKyph/rN3EyLvr/5i
OArgz5QFO2cm864d1GsMt4aKKhT+PGfk88bpWkU7Bl/KqAxIfd8F65YOpo5+C/Vd
9fQ6Dl5mlWBlhCDYpOotJSCgMBvJjvqxkPp8lkeDx88jvOYcSi9+gq46Yh8d1Ic5
BiTs5XgpkIrS2HOTVCFgJ67jG8iuYpVlZmpXuJTNw+E57wExCLelMAakgnolkKdA
3KkqP5z9loJ7XdeJNdSNdjJkhmWVbwxkTwvnNzQozaGH/ADPsZnWpelbnIvRZNXC
UnGsg8j/3Mtje3jeoCTSB3M5O0Vq2SxsInTC48E8aCAc37GhIyhzT31LzTOAvPpO
TMz1+oFpuvkSgve/CUrQOp+igc9o0uRZURjJxHIohCf/dbISmk/ie1pvZMS9xb25
djLmI2FI+7Dg1upDkmyg0SFgySeVCgWWaOBeIa4njaKeqgHw2hPUsvn88YqwtRGf
a4iYID37xfntydOHZixjDqxO7c96bHL9e5OQCjYdzj1/JYvqZqxMZkYOInhyICPk
7BUVEPam4KurPMFBBbFJlNPZvd17J4NtdURM/OLE+h0EPN2ndcVwMwBYTtzHIjFY
ngKNCDAdfVGGTWr50Y+/CSsFvy7hTQX8yQzKhmcfr4QjIrmLSLKXVueZ4aFcZ1uV
QSq6X2nGAuh3rLF1uDixfiGLPD1QI4lFUEVIGhA6m/gEC/d4e8+W7Hyzr4feHhhB
u/GM1asAwwgdVhDm2SKSHOv7jaK0fHhcm0QBAFtHUiUAJHwzby6FYVf+KWFJ06hV
1O+XtUvusrdkTR44NM+4kTyJ1iM/cCPZVErUhuxYC0DwDMdcvrXH3wEk4HOKuYoa
iFs/YZW+VBmWE0/SnAyMrG6ebzk3L8j1Fhv/8D4TWq7aFqd+uVKlqd4l60BSgOki
o3qxzrcqPM72lyQJaQGXCYdq62pmdrwq99SkxQlxJWRhJwFDLwIbHbnmMiiS+E4S
IVJS1t60yM8WHMM165/Ky0ni1pEbJYSFJiIkS+1GvYoaDOdraciMNgNmcbAFFJ1N
WzRg3s7Tv2kIn6/2K8ZcjLectO9dBU1ZjG5n8ZhIar4=
`pragma protect end_protected
