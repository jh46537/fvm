��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z�D��>ܱp�w�����|�8
���v�-�IW91�_��m@��n�P��|k�������e�9��#~28V�(�NݴYס��[�m���~yw����uU��|��4�^�I�3�(SR��2`���Y>���d ġc�-�Kx|ɉ�G6և��Ǽ��j��ȨGz��)�.�3�O^�Аk�YǺ�#:!}����v����+Y��
��]a��7��إ��9
٭g�2�ӗҰ)�}�q@�<�5��L�Km&��R�{�/�(���x�&"�� �5w���a��8Q���ݞ{���C8�8���;��8�G�RW���ݿH��D���;#;ڣ#?��>xTԽ`�(�E"Tm/I�
��A�1^�'��ӿ|����E��9�#���ƍ����a×�UN��3+,��d��q*�Kt�Xt/�H�_����u }�٣U��	],'�0�J.��۩�&b e�x 0�3yß1(0O�.��U���F4�\�^�apE4M/���6ԯ~)|��Q���i�]�I@_���8����Z�C���b�GF�iZ:ΎΉ�Љ���� ;-<��g�S�;s�"La-c����}�[N�#���;	�b;�Ͷ�(ח�����AOm�b��+0;�RPi2��[�K��a�m�zS�]�^����K����c�K�gu_�0)R"Y0C'�Y�cb��(�R^�#�ci�=��
�ml:����κ�t��H�] Q���k5ܘP�ډ��L�v�b6Gǈ��3��z�ˡ`?��(m$�p�:B	#t�������}
�R�'�b���I�p�im���F�u��\e卒����7�cv���R�4���#L���{\R���~�-T+^���s"4+��5��;� y�m8�q���	r;ۼD�5H��^X��\Cm��p>5�aq#AW�=Ur@�G�5���VH~��\��o��
�i��<�p1�B�1�;~-p���k�ۃ��ɵA���sC�W��#&;���z�As��4)�eKq��s���)ɷ�����`��N3/HEE�	ؗ��c�(ʗ�/�}�ɶ��mI�y��:�c^ε���4[����nO1jĻ U-�l�>����N�w��
��&�(��3��P�En�&���ϙ�׉�M��TwD�����`j����lUwL|	�ޢ�Qe�ÀfP��ʫ�7���߲ڪ�����d^V��ޣC�-`�2k���!^����*x�ȝ��P"8�K��qw�?�*u�'�����L���Ʌa������e�x�o��uޠ'�<�g�b�E�/�� J���TKuLn�����ѠH/���sI|C�mr�ϩ^� [�m���M<�����c>���ފ����.���\�7��]R�Qj@��>�ج��r�e5W���J�֧�/���tEO�{���"�|#���OD	dR�Ҍx]����Y|�$��I��ť�{��T\��=Klc�FAv���N�� z�^��1���Ǭh�-�̐�R��1[�����%���r>�����i?�{t�ѕ]ài*s��0� �~�?����nr�e!SsL��{z�_�8M�3���)��`̕\������D5k�q# qI��F_���ZQ� 3+�0~����u���nqF1��v������Ϻ�W��yjA�	�WK�	��L�B�c��M��O|��0�;�7���;��0#�4�|��6��at9�|���]�Vis���3���x�=P� %2���Z��y-��٧��ܖ����!�J����
�@L(�6f�noz*j1������]�ni�����,�ADG�)�Eb�|�i�h�|�Ƌ�x�'��hl)����\��-�X"�W���F�F����Ղm8u�F+6R�Β�{-�9o̫��z��x�˔����������`Τ��lJ�GH��H�l�1	$��;�+J@A������%X2��d��x�$��hsQ#���"� ��FR�R;ڽ��0�Y�5Rٞ��
�����fZ�藅�#ݫ$�滬�g,�d��r�M�H�x}�|~�`=h0�Zx�h���JF����U���bu�����EM�n�r�~���;]����v�'E��<˘>p-�@◺��J�|��V]$��d�<�UR	�=�<��:��Se�ȂW�0x�e��	� #���>n<9N��I���7�<�0GJOl#��p����8v�ܭӏɰ'��u�+���m5A�p�x�tՂ��	�ץq�AS%by<*�iz�|��1��d��t�d���7 &6R��� ��zY="n�����E�0��-��VS�u��iҠ&n>�:)
�֭����/wq��}�6���u%�K!	lXN켈�U�v���$�_A����\�ф8��]ц��9�0�%ѡ�Vѣ I��������b�BF<!:�j�dvsA��|��?�Pb��BY�E��OFO�[��&���h��{�`1&�#h����귈�Y��y�w�5a����+��o�3���*�B���
?�*|$R,�Nw�O�±1�����������E��[G�^
3�E��]`�?�)��oLEa�a�a�H+��5x�~�[�"�@�������wR�����<mm��%�EM�6mb��kc�V��������Yf���Ȥ�����ᢎr'1uX],�:Ib�7'��l4�u00�x��wʞ����]����(�kg&���L>��n�kL흓떡e(��+�.*�A@',�dA���o�xB�aƦ E�w�$W�)jR@����W�s�k�j��5�7f;�m�x�������͓4+�XGr�hd�$*z�%/�tdQ��d��G�0g�m�gD�xV�l�ޔY�0�"4L��7�>)��f�R��+E,Y�ަ�vr��X����X���zB��1{�Sd
����{�ەED2�i��[AY���J���t����M
h�\�,���ȇ=�c������*��Ȃ��������e!d��@�J���r 6�%�ڊ������~W�&�Tn�@2іV~*jF)��rϚ�M���5+U���3�(����+�FK�[�[���P�9p5e��?�V�w�g2�t�)���0Y�J@����>�&�g���}
XG��a����j�2�z�N�jl�x�㘿X爣�08˙���t�r���~�O�`(�G��\�=�A+ք�����G�?ў�d�q�'Zu �Ѵ�"�3C"F�ƷJ�c�d0t*kF7�a_=E��<i��@z&!���P�
����\hk�rz��XY�������AU�Ch>XI���zD�
o<%��֎$˶�B^n�\꼧�
'0�v��ZM�r�����I���)��_.ˋ����k\����18�8�r�귛p�����5�F5����U�E�'4�c�v���Y��G�K���>I�6� e�c����%Ĩ90�Oؤ�+v�٦Ū�e��`K�!M�����ɥ���J�B��I��Ezn8*��?6��#����opy��{Y�ڷ�	�a�V0�ü�%�Ur69�����nXo�=NjN ����hj������k����@#_��DB��HY0h��f�2����5f2��5lR�К&ߧ�a����]�������n�,;��_Q�8��ߒ#�_�r�Zo�`�b�D����*O���_��gI�K�ŀۗ�����%����a$�T� �Hx�3\��󼈀�Y}���Yf1�G����}.��6��Z��l��}y��ۙ=]���C��A�y�3��IF��>c9��\�XE!^����~�Qls)ʘo����������������ҭ
6�h&�G��N^O�����.h�t3S�fs�_�� q�%�_l�K�4f��I�{�B�>� �9`��7�(n�Dcބ�i^���	e��rh8�+�&�.��C�j��_N�jD�VK�;���GF�z��ۧ*��zK���� ��2O�K>%F�#i)�R;�RѺ��:^ Y����Z#�3�&�1��!�a�
mqxE[����=�����T1d(��l+[1�?�a��t
V����m�4�q؄�ֱG��`O�E�R�57,:��a!z�{��`N���d|��h�6{�	>F}Ց��o���t��3�Rk,�y�Qݝ1�g>�qE��� ��f����SdJF��O}���N?�K��<�fxL|���2J�ګ�q�!�~��H���ǚ}<��<� :�ͣH]�@�� �*zp�œ俼*��<��ܥ"4�f6��n�0�&�S��Kn�0�S�ŕ����D��alV��9�
_Y	���(���0�+�HR���/%*t/u�%7�� �n���I�")g��2��Y��E��R�&
ȴ�af��#Eq����}���.�͞x g{ݳ=�o� !����ݥ}���W��-3m]�L#�l��/$`�#Y�Oވ�ˡ2J�-D�M�~;}��y��jV�t+��V�:ދi��/��{H
U=i�C2w��!�'?�|?T����|���ωR�V�5��S��`���7+�^�1��xI�'Ǚ�5T�9��#|"�%�j�S����q��f#�皾�FǴ1�d8�5M����#�R��{3nƜ�vq���l�@?w�f��R�#F��|�,3U���4H��P����c��!�� �ϘS�q �qYQ�hy8U#��U��XB]�C��
7�8�����L�M�߃�S��G &^XùY�ڮ���m��'�PdU�n�.���A�;�K���+kg�B��? ������ֹ����Դ�j0���<�g��m�����xV��{%�(ۑE���I����r�bW��.�^���n��_��᧧�ʱ���_�����ɖ^�Q���Գ&Z
�R������A�V>V.�(�}��W �[�o�X���x�!I��[[-Eְ�22Ӕhi6ْY �� �Ip��1
ܴ�^���l�ǨwÏ��I�#����N���.w�1*���pN���˪�a��U��0e67�bI��k~�*���M�}v��y���ۚT�4�v�J/��9َ�i����<��]LTo�0Ñ��p�O����kZ5&>����p{���g����`MX�o
�^)�ȝx˝E0�0��LxM�qħ��z�!��6%��D��
F1[�*�������� �M-��KIyqGӕ�H�����<�4��=w#�����gN-D��?m�p9G�F�����Y�Iz��g��c�-��l'L8��ή���8�F̶���]�p�o����7U��i�>��6d�{6���%�g-9����x��l��y|Y���#�ю��Z�g��!6�$y��i>\�()�*UO����g���������w��f~Iќ��8֦���-ː��%��?�C��1J��ch5Ȕ�)�1yɿ5���Ǘ��rwߐ@܎��Дkt��&g�'�!�ʡX⃚�[M߮�"�vy�TжyPP〺�5�y�;�h��v쀜>H3�F�-��~��L��t�C�6�3ܱP=�:!	o�������;4B8G���A�A�t)�{Q0��2�e�P��Hw��
���c��6\�޶�ꗬgr[2��*m|$�J��i'�8Ծ5��R�&��Ԇ-����D��d�����qQGx��[(�Փ��}��2Xa�;�F�]-p��☽�
:����J����Ai�Jg��ek=���-� ݜ�����縫�K�����@P�_lV��Ku>h 9�'.������]�)e���N�1�u���+�9-�D��tF���ٖC�+WÂ���?M���
����S��#�H�s`�{��{������G%@H:��[h&7|��;4�U��>��W8����6���Pt$��$.�� ���>����b��g��0���of�7ҿ�`��9���
�`�i�q���ժ%"䶧1�--f�&X����Ǥ��˯t�`Zw�W�km1�x����
=h�9m�s����oA�s|�kO�%�w�tS�3l�ă�f�|Of�G�&g�9G�硩���j��6��icA-���ܤ�d�x�S���SrݹH�y���	yNLJܤ�k�~�Xg̝�χg��;"�pԃy /�Ԭ0FJ;��0�k�mϴ��|��w��c3������:Q���UL�Ҿ����/5�'��J���M�	��ae�"�V-���_o�TI�Snˆ������9/6��#�SK�;k	3��I~<���4$#tu����`�x�> �힄�?����T��o��y�#��/Ln,����A<���ȟ,��Oq^ҮU�a��%sx��Å#�/��U�ꋱ
{����y$MR���NN��{-�#eӆ^%
2*�K#UD8�,Ij�>�}��Ո�X�ԭ���X�����]Pq�y6$���4��jQ9�������������̵�Q�f#�/����W��Y�!�4?fw,,ςv*�
�ver�k �R�⍆O�a��2>�O�0EBεX_�����2���$�mۨSp!�
����lX3��d�+�z��~d�:�g��W�w�s���53�C��E+v��T�Q��X=
���������-��b�Y��X�|{���l&�����%�ANi�A)bv��9��(Py)����7�G����] S�*�hD^$o����A�S�{��������DubuEޯT�'���+y�k �g�r�??@�<�,]%������%1W�����,�5�u�=m��^�cWI�\��2�?��L1�S^i<&��z�U�٠<#�i��`�H�b��E*������u ���S�����Y�8���Q�U����H4	Om��-�Ŭ6��I4�c�Ӛd�7n^�r>�ʴ2�_�;h�J��9�C���}#�,��|�R3�9��c���lR��<^sc�o=#�E�	�F�Gp�6f?�qB3� a��w`:��<M2�v�8r�8�B���. +(���y�}�J���Ξ4D�F�� �{��P��0�Ht�.�u��M�N#/�2��7���8�r��Œ���>�r7�)#1ʙ���=}k\a6��[4�'���&�R,ϋ�;��z��b\�,Y�~�{TE��X�{�����9)�!��#S
�A�Pb�g�$RS)dA�Hq��em�|Rؖs�v$L�o�sh���G/�Jm5��" H���v+�/�b���(z��B�`qZ�Z	g;��()I7�������UU���M��خ
3�I��#A�^�RB�7�`������ɱ�zR����Q��w�j�����{�о~�}�;�x�����'GY�[ܦ���Lr��x6l��{,M�y��Qܱ��h/<j�����<4�A=q�m�~�O�� ���JS���̵aQe0�X�����\r�����&5�7���^"����$�����Yf��|�P�z,��� ���go<yռ�=j�5Q���17p�%M���_i+@�'-9�WHď�n�e=�W)gQU���z�����:��K���o+�c32���☜�H���.�j��X^��*,��b�K�c}(���nw�t,�n�O��b_6r�$���@�yv�m�hmWth��c�r�-um'��Y�,��T�:R�A4A}8�M���1���W�x��ŪU�{<�R ���P�����> �=f�[u>A�S��-�N2&�Ȱ�6N֑�9'�i�kCg���23u�'51�4�s ���I�m։�.��[��pX�_�4P�A��y�������1Ǥ��'���M�ݶ,J𹦙;��<��X�f�y�˳��X�ZC���<��sFa�mx[6�X����?Wu9��]�Ե^�p.<O~��G�R<��l�K ����rZ6��Ky5�`ș��9�8M�q8����~7����;�	���n7I�D�є+��P��A�"��/h�&<z��_G'nX�I�ᑻ�b�Ѱ���u��]�Xt�K��9]�F�Z���H��
VB�e�i/Lh�-���d��,�"!=�妀�)3��ਛp'"ĤA����"V P��mȢtH��Ǐ)�}`�N�$��s�0�x�I�^v�K���"���v��4|;w�C�����#�	G/(�J�st!����%wE�"�u��BS��޶��`��D��Fn�U6�+5i(��{i�{����9��G��f��AH4�xҌ�l �� ��R�w���򒙁�vj�*�-V"[�ew�� [(�F�mK����mm�f�����snH�d�P��[�+����#��	��p=�V'*�R��~و$�hmB%�#�5Wf/������^v1@��)�'��`�dԌe,��j���c�f�_�Ƹ��Y��l���(�$'�VΈ�s6��m[�Uj��2��[�3�}m<��24��=*�T���^1!l[��y�L�k3]�.o��L�K��^���ڲ�^Z��{Q������Z��eb���R!,��cPZI��q��%6�~�����HJ�i��ev�#c2UڲRS��}�Z�� �~s|U#
,t`��收[EK��͉ϒ�,���L�6d�y=���!'��ʀ)�	�?��?"�� "�V|w�
~����q7�<��>�/�Q������M��d���u�A9������=c�	�ԧ{��Zi�`r�+ 1-=���
���w��1 Ň���c�s��rڸ!��!�&�����ë�ǆ�%2oN��L���Z�'���ڼM�X�鵒a�+�X*��U�5a*��<��u(TL���j���nUߤlh&�����ls���rB�V���eGxǹ�p`'6�?ʾ��	t,k1��Z��J~��텂��c�*�yy�Y0 �������)����ګ���-�Q�B� �.��
WD"���4bR|R�a�q�$����Կ?��΋H����}�%�u���`��,NT�w�̾2�E�%��Q��z^_��w	�R�L�S4c1.����ԑ8��#iK��\�N����ܘ6�sTnlX*�8��&}7Dυ��}����UOE�ĠWι�L��ȱZ������?P�|�D{R�(���9!!C�S��)C��ˉ��AەLa��?��~j�e)��k��Ck���g '�YѨ+%����5���5���Z����O_#F����)�1�KR��\����\h�w �A��˲����R���L�:"�a�1�tU� ���k��|5��SΆa�O�a�؍��E�)��p��~�㷨�oKL�o����lQ�ae��W~��f&���]�i[H��Xq��H��L����Ǝ*��V�m,�s$��X%�d��f/މ����i�a��8Z��B��!��9��d/]���!m@+m�a��᫕���ز*������,j��^i�?�ݭ�n�����Դ^�b�1�o^��t���]��
9:�( 9>�ytD�꛺4���� ��]1EU5��闧�W�x�?����Uܩ	L�.���D3�b�CYxȌ��3��z.iMJ���a��E<(��.,���C���t���������f��mG8�;�2�C����,+�pX싍��#Z��Z�NE�>�x��_H9���uo.KA��j ��M�Z}�X����k8�˒/��p���h};M7��Y�w˙�$D�݀\#���b��2�M�ug=���U1z����[��P��3C+W�P��}c��ܶ�)c��~|!8�p�!��c�8ǲ֛'=��-���v2	@�	8���\�4lO1y0���&,���gdd,���F�#��/D�0@�#sY�!�����WH�)R�0�%!I�2l;]"��-��!�=���Yq����?!_��F\D�������u�Ӵ���@gb�-sgn!'H�p���bd�E<00� pW�k�p���tj^UuD0l�I�CVY<�c:z�Qվ�[h��ci?y���&Qf����ؠ��f^4;�K��ӵB0�4�8���X@J?�5���(�"-߷KJ[7b��$�����N+�Dܪ���$����YA�gv���{2c�׫>��%V��FN8Ll}���L���xƲ�;κ��-ס�i&���;��XLӸ�w�M��:J�	��乯P.�z�R4^H�IV�����8'���$h,�W������;T�a]ֆ��}�<ɜ��c�s+��>e�/)?!R��H��r'�q\��t\7�Ȱ���3�73�|�цh�4̳��,7�/���>[.| 7�3�tfV��p�Խ&�	b^�Q�B��%X�"k!ls�K!خ2OG�&0��#׍«��+x��zr�L$6Rݣs9�%�M���:vk���V�2Y�#qͯ�O/͋��A�y�@�`k�C����Hf��0�Q6�� Dj4x3��蟞���[�z�2E��O��(�?��D���V7��ȉh�1dEo�%Zbʿ��ݎ���Tᗂ����_;l��&"A��oFv�((��J�F���h~A5wq�y�b���c9����A��xp)��e�c��{�1�M�L;�wv��(�lE��5EX��e� L�.�ҞE������%�{"��瘻b�%~��&ޮ� ��]���+А�K��0'�V��gj�.�wI�F̀z�g�p���u19G.G��R���`�_��E\9ў$%yS��<�R:���ǂ=��PŔ�������uj�?#�c���ik���M�l����y�X�Ӈ�|�>ʥ^���E�����iD�y�J�69�HJx�>ک�S�3l�|$���.E�w4i�K��߬D�3ʋqtp��q�a�Q �5y�v*W����Z�4b-��K0�?��2(��{�&"�bg���n6X���53�HQ]��{r\"��j�!�>h�;?1<o���H��<�-�����[ �px;��P�JH��>&�i<{ڸ"$�@��mE�F�a��D�X;�l�q��� ]�~d�\^�&ٿ��9Z�x�[��w�L��\���_�v�_㭕�A��j ���H��\mvvr;�|���T�� G�
��q�	s���R������� #���$(�v�®C@����Y�� _�p��6�^� ��e��};������w����|��P`��Ҧ?S�V�&����������2)��=��(�g�Ŏ����ߙ�eiΆ��ڋƊB��D�"x�O��Њ��H��gO'Ƈ�F��Ћ�R�C��3�?у��ٽ-��/�����NM!/���L�hPyI*+��2} D\��`�)I��I���ȋ©����|���eEƋ�*�a$q�m�*1���k�Ye��P=����u�=�˷s���%!?�;8I ��	������/k3*(F�xĻ�*Er���S�A��5#gM�~wN�G���/��$�63�n�UI�u�/Ε�n��G��A�>�ێې�/�+�aW��W9$��P$H��m<���������K��o�ܦ�A��4 �[>WL���� ��Q�g�aB��%����$
6��)���&u۸����2ce���?�	�2Vٺе3!O= ݇El�nw�G��.�F�����q�&$��_�hUz ��V\z5 ��e�9�>�@�;5I7��5F|y`OJf���ڝ2���v�΃ur�8i/-��M�����{mq�'�k���h������K�� k�������T=@v x���.ƾ;�\ޑI�kl�vܵ���G<�͚��I ܩʈ�h�+�N�����Y��ٷ�.w���D�d��}M� ��ѱ����v��S̗����{�ڃUJ�?��}|�&D���4A�.��o�ƅ�%�sg8��z�-�E��ϕT,��v8�Rq-�rM���>lw�Ȥ��R�_[[r��
P1\v�����ŵ��M��hwP�ri� CeL:�@��ck�1��ft)7�
�d�Z`�s��j�c3��	��\��v&L'���,�A	��4��8�$Q^�h2��Ң�:���d��V�O�:�$�g��� �,�YS- � �Fk֢Q2��I�*_�?�&�PD��UDTo�+�8�\�=��QY��F�	\�?��z��f<�:�9����:�����w"8��o�{n3���x������Zts0�Ս|�UW�ğZ_�!%��<9y��_c\eň�Cçvl��Ȇa�" �����ݡo�&E$cX��-3�p�wRn��g�>�pdc����+L�M�D$K	.RG���w;38c&w��k"�k��-��?��夌$E��c�Z��b<ť�7"�(���a0 O0�D"�#�9#��&�#7	������??`�È���ƂF���MA��ze�Y(��f��G���/MG���+���p����!f��$��b��v���d�k��Y�2�����:.�+|�s�g�� ;ew�0�D�SR7�?N�i6KD"����9�v��"6C�ܒj�2��*��R��1��C����u�L�2(p��C~�\���ÄS�_LA�<3�KX)�vV��|[?^�n�MU���vz-�dH��>>��I.b�T��_�S�:iO�],J���a_�]+���;�q��2�����u^c���U�ZL�Шg'��Y�bt)�}$ 
�X-��Pu�5��c��+h��&����D-�]���W86����y�3?���Q�}�h��V�����[}���1ѿV���z��j 4̖�9�ƨW��Tq.Lo<łW�8%���܂���.F9N��jV�����Ze�S&"-����H����P��  ��zCg�@u�l�UZD�T�OF-�䡭VVc�$��h�&�����t,~�ᔭ�+���<�@0��y�^}��иO~SU����Zˌh&�z��,�j�ȯH Xdl5�4Z���` &���?Yt�#Gb��G%�o;"�$���}2$����@[
��(�+GĆ��2�`P�`�f*�ׅN&&�F�&y�b��%�C��ҵ%o5�|�bS����4:ޗ�lf��2��4@{s�Id
��,ڑO���ga��{��|�:��2�{���f����س3ΰAX�‟�:�}<�[tϢ��e��}�c���_��eQ:��a([yxĬ�9abW�Rm3�L��4�Q"�(�{]k�� \�-�O�;�r�Pm	gR��'7]eH�u���{��&�́d��=��*���S5WWWv����j���c]i`��F
����U�y�E�.W�ʳ�6�(��P}f=��O��')�^	��=K�f��)�&)�G8����O=�P҇���	�j�
C�g/�+���AA{���L�
�Zĝ�1t��������`V��]�C�/&�T�����m&�Jurm��mV�웩RNUD��`�.�����&${��� ���l)=��M���#�G�Uy�"�:�]t��Z�t	�:5���
u�c��g����Y����{,�Ԭ>Bi�`9d�P���z�Ŵ����2�j_pu�����P�h�tv29=�K�(^F�|�%r`�F���=�֣��GIae9÷��b��P��m�� R1��ߺ:�9�0��5��(��/����xx�6�����GQ&H�
[O;�Id 碍%�F�?|���*j!���[�2ʇ���~���u�k�1�~ٸ��V�1ׇ6��dw"�\�҇���1�чrgv�a��|̜�lz/}�������8!@� 't�e�yΆ�(���ӳUz`,$�s�~����3ׁ�^8�c6WSM���b\�� �3�}�3���޲+O�3%�]�(4��Y �u�O`�{�����ݣb ��0#��A�%�0n���Ū��q���ZYk9��.�G�P Z>ű�Ʋ����6��P\��t���O���D�x!M��o���ќ��� /!�=t���������8Ծ/y�\W���^F��rT�hX�P�j��k�j"s�&<-�ަu=�zЊK��꠫�ˑ�E)i#ifj�����!+-��4�6v�|������@@�*���[>,I�q3�]!�^���յ-�?�F&���J�(=������I�Z*�zS�zX�\��qF��,eM�9�0ʼ��n>�e�n���]ƀ7���|`�%u�T��yBm�>`O���ȹ������Ho�6ur�S��>I���\LuPx���Wi��	�4i'�l��*;�wI*�ɿn�9s��i��i5�,�{��:��p@�wio'22i{w���F;Z�I�?�����ح=�c��?�5�ŧ\��9��vNPn��<��48b��B0���e~����`�哀��p��rŸ���Y�|e۾w���:��>`�SMH,�!�4(���(�V�w�	����[L���� ������������t�i��қ*��)e*��i����w�)��{�疛�V��������S��6B��u�.N�b:Y��IB��*�I�q�,�k�#!�b��Jt�������ق�rbJ���Z�;��5����V����%�#!6Nz���|J���{�#��zZ�2
��{�D0����%��m���4m�<�~�S+��3��sV-�<~�%L��7��"���=��ſ�ai�V�ÃW+�#5��*�6���N'8|�a+GJJ����j)���1pj+4S{[�i�W*m%�\mD� u��k}�����?�{�\��W��y?��� X��8�X�����	��
�a�JF�)��m��B}J#7���s}���Pp�j��0�0tZE���(��x	PT����]�lS.�3!L�Bx����C�������Ѥ�{N�C��t)I���[<��L���+��,�R��{|f���Jx(�.��0��٦\lS�/�������Rr/�+�O�2vǈF�uF�]J����!ԑ��ѷ�;��Չ�W�����f7	)�����$Nt��=R��kt����1;����|�]����
K�QSᩈ�A�����-�4���"W\�����U���g��:_�5<�^�s��2��?�rq�|=�a��(F�E������c��6���4��C��*c$�IoD7��/�)!z<+�^J���ġ�Ak�8�!�D���[��.4�Ä�@� �
H�_�/����b����Ǆ�s�,r8ÑYJ���gس�K���w�/�2�/J/����ް�ƗGY%_GN�ҙ�_&av�UO�T%��?����u���¥��S��ڐo�"p;� �Nd�y�w�}E�D��K�R>.�F��eB ���k�j%�fY��Ѕ��F�ٚ1������\��ʤ6k�՗pj)&�d�ٜ3�~Hؙ�n��-�u��?k!:t�E��~`�� l]�׾*\ȒKy�Nw7�tsRȷ�Z6D#�7iu���t��A�Z��s�g�Ga:�h8��O�DD`���@���������TK���s	.$j�%V��K�V��RA|+&�`�,Z�;���*��]�"yC
X+�� ~#�q������%�Y��ݏ�ʸے#'W�.fh�|d���y�.wU�@��������<Oa_#nl�(�|��Z��ͩ�[��l����m�]`o�o��Ӥp�<�5ۘ�᫣q	W����Є #����x\S�8��20�ƛ�� p�v�����x�^,�s�|g�ۋ�p�c6̆�@���N�_����6�Z��J�Q����\�'�}��@;�Z�T]�񴈒�j�N6O���k�߽��,b���F�W1����[&9X#S vh誠wU��E�28L8�����
(@s��iu��
"x����Ph�=���� b�5��k��.�C7������%#�R���lt�o�s2s<?�\��Іɰt�J�D�q��65W���8�d:�
W6���4�ېѓF
�0���)�`��:	Z��B�*�����~���w��m��� y;^8��0�40�E�R�P�AVBGf˻k��\ o�8��m�i�]?��iʊ�Ths���iᗉ���O��hjP�`�������t#��D,D����_��5>Ǌqaɂ8;�ʚ~��>�f��>zv�X���Q#f�6��i�&��ב��^�=f��%����c�����Śt��$L��p�]3�Q����N�㛑��d�F����Z/wu�^Y~=6�ֱ,ѢL���+�J^y��"��d�8�D�t��c8�:&M*��O?|B�I�ʲ1oNw�Tk���B|�x�kJx���1���gg�a���'A W�� 5]�h�6�5�мJ@�h8>U5%��<��	��zpx.�?@	�]~�!*����p�w$q�BZ�:���L���l�_-���0�'�p�����������g�q���׬2%�~�Phn�/��
"�
�7qc�gF���CT���f��A���tһߩG��v�y�=���L�o ���j<��)q�"n�N��n	��q5�J��js}6v鼼;�@lRv=�(��"��`��4
퐔D�@E^jz�n⎩���ΖGش��k���:�� &����U�������Ag]��(�WC��~W���&���B陬�����V�y�tW+{��&��:��"�ή��I���p�N�6��G횲\��N�^����B4(��x�	�@.��s�ϰ�@�Ҫ�'��M�ƅ�`�v���%���l��4|��a���$$0����r|�	o�>��8#�J �~�5��A!��?��=����Y-'��5,�W�����]9��y�����)�!`��Y��z�c`<�R���;��:�� ��Ӧ���t�S��S9�[3��/��ΐ�]���	� P�;�w�.���)�b�ʏ#��jő�r��/�{<I�g@��8�C:Hӗx��\��iOkg�+��EB)�/���d��`>����4ضD�r%��5��%�8�x]�?[��P���ĕ����[yzva�5�<�j\,��)q���
 'oPdvmF����ýv�x[��cGV�I���Ӱ�)8$<��o@�T6ip}Ƃ��8���k��=� a�C�,?P�'���m��!�)�Jw����M&	t����v���
�ۍ�lb���{l��9��ҧt���B�����@�"
��d�,��(��R�
88���O�s��lP�mW}�/�f��[#�f-@g%^�f���<�R��Fv����p�\IK4� [����G6�"e�D�IHA�m���]�stOj\/��)ݩ�a�Lw�IS�/�Y��/��S����`�vy����ڥ�,K����l�������F�DG��'�YZ	r	���bi�9�I���l
������ŕ�cQ۴�[,0ZQ��jܸ��-�%�4�g��p��"_�VY��H5:�K����,����vv3�t� �>�ڣ�m拋�qӂ~��ve[ۡ�[#DI�ocl��J�z��s?v�#���
��Q�R�Ȭ2��z�R�xF��x��S�-��
��.K�h^5!�g͒K�^v��3�	Y��A[�e�!��v��mU/-$�0�q
;w�5��T�$8��r�>�S�J*�Ѧ���X����T�'�q=��&�
�^HB�-s+<݉	�#��p�=�D��[�N��c����ٿ%	Sn��ͩb�;<���n<��Q�]%�ҪH{��z��vexU�����tK�p����=wO��Zx�H�̦�d�gC���`u�u��I��72�"UW���L L�O�;���8����k멌UUS5K�Q��!��y�����	���tΤ1���i�e�8]t<w-lԣ
B�>y�on�[9�JwQ��gy�Z���,6���A�+:o�������k��1��:�
�3ְ9���#ڝr$�>_&o�^�xTm������*��R	Ww��l9�O���t�Q��L�V)�x��7u�⑱׮�s���R\�����}\��r�	�k`��.��w��Q-�ɝֳ�����/*U��).9��P����y�Vf���t&��L,�Շ��$�qx��0]Y^�H-��k
��v�k��`Ƽ�-��� ��u��M(,��N�a�_9�a� ~&W�fh<��3i9�kD`i�%4ð�4��;��;-uk�m��'��	'r�p�W�Ђ��&�q{�do8Q��e�g_��4�t�?P|����dDm!2�������ql	i��Y����S	C�@���v���2U�Rꖲx֣8`|7�%-nٗ�n9��q�T�C얢�)��b�çbQw�v8�o����rK\��HC�3i>��j�Vz��	k*������/�zv��hvˆCwf "�;۝��)1�3��Wul�S�[qI�	�l "%�X������*i� ���+�&�˩����%�4Vik��막,��\]*��6U�1��ta�t��~��4}`cӳp��k��Q��}�Ap��憦�ƥ��;O̊�Rwc �b$5�����5�i���_�=;�V��N����K���\�MƠ�m�/�KE��h"���?���7�?,����s=%%Ec	˰�Pǃw� 	�G-�����S��w6ރ��-�;Y�q�����̨z��:a��Wu7"<�Ms����� ��H�U�ν�h�U�Y1E�@�R���V�JO���lO��=�Y@��d ���J#!�xCf٪;�U�$�+�����x��c���	3�#̘�� h�5�@�a�	���3,$�M|�)���c'�N;������I7{��Q
�2'���s���q���i��6|���*@DUƐ: ����,��8o�9�f1M���x��� ��J9Bo����ИZH2���1!�AW>�n�Eu,�=Ԓ1�=�<ݖM��q��n�L��K��B�Z���Nx�V��5���b�KȞ�j-����fI��)��yl��s+��ىuedŘs{��E�H�yeU&����HN����Ĕڸ�~oj��2��AvƸ��X�a�Q�:��j����n ��*��[� oG閆W}2� lA�6n�-1���l2�ݍ�)��O���ӝ�q����o_!s�]�v��(y=�~e[�d�P�ɒ7��AfrR^���v��&���ˠ*e�yΒ�>�^�1���"��-J��k5�*?.K�Έ:��8�5�mڑ�0UjmZ;�\���<�@�����"���Fz���虤C=�7�G�CW�rZ��Tta�Ze�@���T*��|ᤦ������3�"�do��fd���X��P��$�f)="���
�B-���3�_涆���y�������=:��;�����ď��X?�6"M�|�<\i���G�(7�+%������%k��o�� <<ʖ�QNn���J*�h��x ��!	�Q����O%����z�����̏� �����{��!f�+Xp���W� �}p�Ucͳ4f�.Ft����g5���%f�O?������}�4{�휉MQ�Ɣ]-Z|D��[u��v�,�sZ8���R*�{��͊�ų�ӷ�����yaP{p�*�U*R�X�,d��SVqk�_y�5�r/`�(1=^�C�CY����'�lr�4��җ��c�!�_��b�j\s�&��v�8(��M�%�']���?����B5ò�4N[uT�����mn��>���M�;K�ke�A5�n�W�l�L�O�hW��vڕj7�VX
]P�3tj!S�X�����*j��>�D���kO��S���K��6!=� l�qU]Zn��nYYb�x���8��һ�ш:���KryMQk`P�f��u]����$;������\��K�\1B��k[��kjQ�K�,H��_�:�2\0�բ%��q��E����p�Y#�� ���٪^�kί�<����ü��V�����oN�\�\r^߬d�*<�Q���7�3Q�trD˾��:Œ.��=@i����?����1X�ϊV�̅v��8�ȡ� ���IS
���C]F��Z���r�EO�d�=�o 0i��w������2c�Y?�_��K��B��9sK���d!~��>��G�[�@�A�$E ����N.�z�>G�M]�G���+�.+��?�^���9���a��K�,j䨲y���FB$�y^C/1�XﵡZYE5�q�5@SZ�d�ݞY"��^�v��Q��3m-WXx.�F�O��0�N�IyL�o�8�cյ ٻ�V�}(W`�D4�ٹ�D`�=���Ft@U|�}v� �"e5[��U0�Z��6Yn	T&�6�2t`�ᮒm���8�٦_�wo,�����kw+[&ѯ1mIǁgs/���*�$�(�^����K��u�cu.W�i�$��O�����ىz�=�i���� u��?�2ɣk*nl<��o7tL=�X�f�KH��<�e�����V�/�ZE����T%[�8d/�B3��r�j�p���s��*��t�!Z�n���a1��A�lgac,����V����kD�P� �r?w����x�A�lu�l��?L�P>��_����R�<���o����K<S��0��֎	�Y|�{������B4����LG�|����x�jg�f�w	u���.L.�-��ۜj3}99�il`�ҘS�D1�
qԤ�����Y�����I��4җ�M��������E[1�=i�:&�;1�gж\���Zik�XN�6�kw�o��^�tX��<��!��P: P�(��o�ER_Ɵ����R����<OSI௙�vD'iA�&?���3�Zz�Z���C���{��! ���~��� 2�,WN��NA�y��2d@���8�P�ny���F'�f#�M�F�')Cإ,c;ΰ���"c?� j�k�����T8���O�����;˷ցF$Je�\̉2(�<�L��`�ٓ~�|�0vʆ�J�	��ί����S�'K *�c�	*n�p�Kk�#����"JC\zS�E���53��#�H������V	�v�в/��`�07⍮�]�ô96�9�k��Y��W��e\��v)�" ���iF�X�ޕ.#<���H˳�}�Љ���jWug���l����։D�=OH��d�����I���BcX���9 J�Ko����p���%�Q�zm#6�3Z��E��k@�!0�,DZ����&c��� G�N����ZjHnK������ DA��%�`7�Ǫ�nh@��ʳeVxW9�n(�����:�9���}5-�(��3юA8��g�Jv"�ڶ>㘋�Թ7���������hڵ}ĳ��wR�ߍ���+ҍHku��œ�ד�M!6y�P|��� �+��n�R�?9�d�\��B��e�I=���ւ%ˎ?P�䙛�s:\�����.�O3�dbe-�gE�y�+ `#��Q�@
���aG2���R��f�oS����9̾U��Y�����ޅ>��Q��	��	����}pꟕdB��R�	�#���ݪ�喈\�<���LF����wk�p�9n��]	��ĭD|�%���l�ت�q��2�/*��F����\@��&�Ss#��LJ���H1bU�켳�T�@=��w���J)@� D����{��b���_�q��(�Fx�w��sm�O^���OJN�'����2��+{�Dʁ�_p~�R�)\m��K��T�ܢ`�+-�-lM9����e6���H���Y��P���F-#��+<��^p���*�]z�Xg�d3?��~S)�A(�~Ed��pQ��(����-�T�ߴ�8Uc=����a��,��#^v�O[i�*S��۬<�q�[��@(u�M��'xp$)�&1^uX�L%��g�P!�n�;M��o����(a�,�.U�}s��r5�湟{J�WHG�V�%� f����8�gFy�)�{�Y���FU��.	<LXsb���w�
�l4�r��@�8�E���X�]-w�����6�C�D��$S����=�è���l�r\j�����A�����b��α�W>C;s>�� ��4��p�s�"{���;�"gΓWlk��������)D������u�f�����V:�T=mr%����G_MC̮ē��yH7h��[��۔H��NF/�G��T����A\�%eA1Y�vѧ�2	��C[$�B��������'r,$Ghw�3k� �QK?����jA�g�)vͱO(~��Q3�Sy�'DFޯ^)���_@\��KM��#����Fc燠σߪ�tn)Iź�����li5p�2;UI	fH���fT�p��X�+)�q��dn�8O�_�X�O���N�Y�4ʁ��g��Ր�t�(tD�m���������nD�&X*���H^�^���~��e���<×S���-VXhNuSdsY�K�80��j�"�^���?:��n���On�����Biđ�N�U�v@?o$�j�ne���iA��YRL����x��T���7g�N��c��$�c�Hx*0��;���C�N�4t��Sg)���{��I(z���ퟫ�H'����N���i�"o��/yP�:�d¢)���kP�����
$�X����-���o��|4$RǊ�����!����P�o0;�vh�I�
	�_T´\(�R�"��vg~uP����ѻ!R}Y���|;�G��-b�ѴqC�D}Ԏ$�*-�m��gT�s�{����e�
�tm��[G�'�]=	��x�t&o�Q*z����=�����t������҄��M[��=�K,���Qt#R[��gh�6S��������ٮ�} ��Fc��k&׻!������w_D�=3l��3.Whk����g���++�%�gJ��0�#��L�h%��Yw5nG�.��H<�:��8���*x��`�@�-7 �+�׋1�{��+��M0�"%hB����5F}������
5�0#9|��rOoBn�G�,���q������c?CO+4G��O#D�5���u�@ii]涭-��MA�keI�*7�yK�lЭd��(�9A�0���쉀�Tyė�D�������*��+^M"��%�j����&/��Ѻj�(�&p(w�~9k��1G`�
�+���e�$���E�;>5�ɶ�ϋ#�yS�W������e"�dڎvA*K6� ��=!�6���z
@���+R�/
���)����6��#�"��.0���_Ⱥ]�������ʯr�.Ԗ������$�bK�ɲ�?�mx��4���A�O5�v#�*�BMiٷ��`�T��궢��b��z��8�[����$.j��sH�i�r�r��8�����Y��:���GZQ�>�P��y@�l4�b���b���KW@�߂i�瓽7ib9ڡ��>���k��O����^J�kKd�$Uu�p�_f�/��)�������L�kP�ZWGwm�ۜ��_'1�q�17�	���KC�᫷
3a��ͧ�f��|9�v��`*�K��G���H �{\��gT#`Z�U��\�v���m-�u��ܠV޶���d����E2gtX����ĥ#j�~�F��y2N���ںLɩ��#��t$U�k�7\ȀgO�Q�[�1��g�5,=
@,�]�g%��Y;4��8x��b�����.!�Z�xBY埠 u¥�O8���K1�a��Y���C�tvDy{Mp������f��
�//1��@���(|\!,�jy�M�̰R"���DnpEX���A�.D�����~4;%v����F0 ƥ��652�/8Z̕�[�U��� ��1!.��N����Y�e.�fcڷc�����lQ�9ݠ c�v.�=?[�61b>�L䅷X o�l�b	�2��ix.��YCA���J;q)-��]�ADj�`?�\���_�,"�_iݼb�X����=ki&[�4��ꭌtHž����(�v��:��k	0�9�P8��1�=ࡤwǼ�d��q̃�����]O8	_���(x}���`ї^&�F6�B7߈X�]��;P=�LJ5��q'8	�9/O#��~��c���h|{ƬI��1� ���Yu�mh����@�/T�C�h8���R�2t� �6?>f���Ԗ(Q��
�itLB�|B��^uc[�I��=��G�=/M�#���πFM�u+�C���KKۛ�1�B2�O`~�I�` m��������Q� R�E=C'>]p&r(�ܨ}J���M!����P��^�#����z�+^6�U�@?@����%�K�����Ӭ�P!��7�a�n֥D���Tߡ���1��XPH5,c�갉�⠻qT�R�*��V���5$0���voM~?a�@nA�G���	Kݖ(��_��2�ml2Ĕ;y*6�S��\k����x�Y��*p���K�𛟤������f��"+$��(q9���p�/]���P
�Q���e��_q��^�ֹ��4���y�%Ɂ�t���%?����wRv~�A�Rm��KG�rYrB{�{2m�&��ll]<=�Cf��ǐ��SS"o�K���n������[z=w���Ym��;��l�K4�8/Ds���p����(��KK]�;I�����O��U��J������m��Q&+ �Vfe�}���#py,1f��N�͏I��Ͼ^�Ȍ�����W~��28x�S�.9Ci�>CG���n�|6xUqK��@>V��o�*���I�i�u�M�7��	� s�`�{K B�iA��L�G�h����Dz��$��9�ic�8�om��ȃ����ߓ��ݛ�A������lQ��j���Z�����n:T�*̾���d5�.���IV��ǷxyE�p8�A��ޞ�Ġ�� &��1R��vI5�[�.�w���8�5NG��������M+��ׂ�J^�׏ڥh���4��sE<�,�������~f��@��l��� ���ͦ�1�^����O:�j�6��J�Fn\>/�a�+0�,P�$&T���`!��U�wJ&Q@a��e��6�����ti�I�߇]7������H�f�`��u�&ow�"x�֪�p��<(�߈E�Dx�Bt=[�SV���_P�xŀ�����W�p�A�x�x؇ �|S3���x�5��o#�^��f��E\�-��V���p[J���u��1cG�9���%�F�1�!��h��ڐ���B֬LF�|��$XB���ɳN頌W�^�'HlX�m���Q��"+�ƙp��.e�����D��f�wn�#i�>��	��}�&�!u{�TV<'=���$+sw.��JGBdk��֯���te8�tJ�S�D��8L��R���#�bq��s�q�kq'���m��Y��KR��֓0�W�������_��j���Μaƥ���i�
	#q�?�r�˯4�����X�
6�nmI
�6�ǹ�{]*�	YL�=}�g_�����.f��D��$��N~If3��5g)���e؋�f&gJx;>,a�f�?OM�S�_�n��"��j]R���Έ��W>��2-9�}1 �N>�G�P�3f�0���H�.ޏ(�j�#�3��c'ȯ�t6۠���s}��]�}�q�_��*����B-��*� ]��<�<�93}h��ey)֬�
ٜu�҉�2��3;�Ԇ�|�b�B�ή�l�ճ=����Q.�e��Ų��@��;����;Kֆ��K¶v�b�LL���N����7dC�[>�LeA����U��Q�x@шm�7���"�A /�v|���������D�hܳ�Y��̋��tj]���@���e���r��+v7uuU�,�ד]q��9F��s��Υ�?#�A͚D}��έJF_��GS�|���D�;|�a���o{"y��*��� H�~��L�����g �f���ܭ�nS4vj>"B�sz��%�����g��eBߔMOu��b�A� �)F�xW�	�Rb�E�g�k�'��+�G�ѽb%�(�9����HRm���I�v���Kv�p�8��h�Ĭ�k �2�`�8ƁsO�A���(�:;+I����+�EY�mFy�pw� �N%�'|�^�쭞��S�V�,��"��Ѵg\o�X�q=$)�+(Y���A<;���mU��HU8/��|�O3��x8֑�i|OF���.g �$T��f<�*�©) ��l����H�
mi�H��	��|[7MGإ�����@�j�5-v��廏�83e�����9��'x���(��ֱ37��P�?mF$�d��
֭*[�����&�w��q(#O��?���ND�]z�D��JÓ��+��7��,�GD�
+?���k��9�eP�(5�����M}���W7�+V�?WWb�C}&��|�$ٹ����v˥G�C�'"/��%b�I�O	�sn�_���(�:��q}p��#�I��y�L���S���@݇Y$�ߝ0#E;r�b�4�#?(a��~Di��Y��
!��{��Cݛ7V�2M�I�mT���9�uІ�/�f�T�vv�&�`�I���ꘈjWƸ�\z�lp�[���!�e��^"?�@��`��Y����L[F.��f�օz���;��/4`�/���V����� ��Jϛ@��0�R�{YS�WJ�i�¡_��V3V��Z[���|����E��) �`�tELlA�9p��T�6c��o7��ԟ��q`�EY!o �y<��F|����I�&h,2���"�9����#Uy��������K0vC���j����ᕗ�S
����0��X�?�%�ħ��J>$��7��%��6b���S�.�����t���[�<}��/��W�����
��dڲs`�P\L�ey뼓�Bq��:�@ɪ�].�@�y�E�(�	��ds��*��[�ȩUҲ2�B��2x�����BT*p�T}�gU����QO���F���Zk`<�x���a����<��j(~l᱈�Õ���-�^P�f<h�H�P����{vD��{~E|�6̓}�4�t˄��
  ��L]��O����zu���s�5*��P���㼃�
7�9�'B��/0�D�@�(�b�����a�#��~v>�	�#r� �6�ha~�O�WXɴ��!�}��6: �0a�OK���TRU�;��t�د��2�^�%	�NJ�1-�×�o�� 6�y��ڱF�����I
��?�Ѹ���8�r�˺[�W>�#�K�
͎�����K����cԙ5�`���'Cp�Tϯ7.���F��NUɫ����z�5#�X��oY���� �l[1љ0?���Ñ�J��ݱd�{ȑR�R������S�.kE"&�H������ڷ�g�����*��v�k��/�"�J I[����o�ywNƊc�v&;��8� 7�� �-��)�Z�J_@^�C%]����5z8P٦�J��#������h���������J�V�V}�������fc�������� �.�ED�xދ��ڝ�^�P�{�԰+��V����� {�#�;Hu p���>��4��)�����L�|�����d��ֲp�����[��5�Pf=DC�`��b⌿!h�Z��1
�����>�qs���c@9�"2kT��v ZUL+X��o�K���;|=PY��hp��X��}��j�X�l9J;�Fḻ��)G_&+�P���<8X!ڵ���5NHDŴm���X�z���X�=�ie�ې��^��M��ρc���E�ǻ~V;dJ �)wɊ�;Ŀ�t�-Y�8P��.,|/�U9$���
w��)fǣ.;|JN��Q��4gIc���q�ڈ�,���=H�u��O`�
\7~���eX�J�ړ>	Ϩ:�4,>,��]A��옸�������ꕨ��z��Z����yin  ����'Kl(x���a�j�P�0� �7��ty�=�r�+����@��
�#K-���AGu8�m�;�V-�?ķЖ�����,�I��7Vx��R�����"���g�73MR�"�|�a�$�䰛c�|��2a�ed�d� ��r|�oj|��I�$$ \g*p�[�U ?��VG`^p�g>E�x9��f�F\[#�6ؼw��U}�&q�k�c�����E�px��6�z`�~�g+ϡk�FL��bR�k=GL��vv!2��kY���F�}V����|��n��]F�=|/�.��U,c|�6���i];���zO�Yv+z}}2LwV�.��a�e��ԫ�d�]ڽ4,��<��QCg��i�LN�3�����u�I}�3����?�IV�S���ޒ �`��S���@�X����|�)�:,B�����mK�p0�ԉ Gē�����iޱ�O+�P+�BU �9ʇ�@��	�.�F��Q�,g�Nw�t�n<F���\}��1�~hqc�T�F�g��`����J?�:�Z2۔#ꯏ���;p�`�0'�?鲢	Qj��h��'�:,oyW$�����Ƚ
��QW����E��Ge8F�3{���_�{�z��4L��V}`<Ġ��2/����ؼ�$Økт;Uӧ%~�s[{����%���t�]Af#I"��k^�x���=u}�����*��x���_q�^�-O�{.0׏A	�ű����z�*Y��$�2u��&?ԣ�@���`Y^\M��;�k�/��v��>�kxi�Wu���ڋU-)3����f�Z�s�}���8�L���iA�c1U'�%�(c������
qIJ�mJM)C
��c�`=(r����u��\v��j,�VJdBU�?�M󥣉oSX����F׆F���s}#b�/]���JkЮ��A���]yP��V�we���$)��wy�S�B*�c:r�X5�3�� _��-UK��|@r��6�2�N�V�-���_�H�P��AH��h�����צʲl��x��ζ�	0=�>��y��뤼4&�5r4����!���^G�7�%y\3�_e�R^g���3z�'d
޽�����.���	"*�vP��̢9{�Ĩ�a��*�ڹFNܸ�|}V���JmTXn���sq�Լ�b��cG�*�@[܂�Z�c�7|����Z�l��IJ��٦r#N�5)�L�ێ�+�Ag&��&�����l�� ?�aHڭ�l�s�=��h��P2�w7���������K����PǊ���x}��lYH��RAʵt:ϓ�A��S�!PuJ)���O��w8O��=N_��`FWV��O�Xɸ�{���o����&,�	�e}X>� '�ݱ,P�8����!�O{�El��%>f�L�α��\�@�q͙OX9Ի�����]�D)9O6����ޞ�>w� ��G��<;���+�����NYd����n0C1R'k�tF�˄��
u���!÷ ��ta�EC������{�I��m��[5�����K��v�^8xx����Z1�$��k������3�_�4?:�T�_�6I�j��Ag���[���(�jJ#,��}N �V�����:�ʺ<0��׼���S ͫ����	W�j�}�J�@�ާ^�}��O��2�:�6��$�v
~ �N������vg�~�	�wu��#���"�,���(�Z)/�	��̝U�K���C�)�!��L<���Ǌ��tL�Px�-;g��e��Q�V
�Dl%E���5�H&i�1haM��5�a4�����D���^'N��4�W���},G�ח��%������s=xk�g�R	�8}�zIQ��ߌ�w��*��U�ߠcC�� w�0���D��_ 1�~Q0Ւ�,H�Ћ���0��v+��H��K�Ro��[
ݟi>�4����=z�vEU�(}N�v�ЗH����9�@:8�-�9���o�nS8I��x��`F�O�Dk�S����]�}�|�6S��K O[��29��F�S�����2�|���&�U��w�*�HV�r]t�s�UX���`��_�KK^�'�q�^�g(��OЭpj*(��&d�Ϲ�W��=��Ќ�"%q ��7۾����{�ռ�0� K�QH�w��~d�+mSj�Јn����2ݕ���P�n�Zý�6R0�Nr�;+F�?=Xn�IM,�P9A��_���G}��S�Ad�}����]x1��k >�k�B^��Ȳ�����@�����>�F�ܒ��4��V�5`9�p�q䇪��֟�|��xd*�^���^W���G��nm�t%���K�<i/I��Y� ��(}o��j����ӝB���&!]_���K��S�z�9b��v�>�Hd �U��Q��Y.7s�T�����\������Iki�;e��2��a�q[Cn}��c��&#�ݖ �Q�Gu���Q3����Y��氿T3�TƓ��"a�����Ӕ�*dB=�ok}5��g���^�[Ӎ��ޢծ�5��B'�T�b����E��G4��-D��/+&�<PSH''�M���.V�S�z����(���zk^�����zw�br�H�ɰ�njϏM#�g�H8i����#~����K��3喭�Yt���	��VGuY��DF����pW��p4sq� `'G-�wy窀��i��*�H��=���z�~?I�KI:"6>�