��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�^��h�����mb��feE���0�8GI\�VE�|E�T	dݹ._lR<���<ߵ]�uj�x i��6�n�m��~�~{~�b��D�
0R6;�a�c<<��"�UV�Ĵ���!�g�m�c��_�t!��dR�CQ���?D���wk�	����h>񪐒��n�#�E�՝q��z�&{6Q6!Q/����&Z�@��L"=��TB�MpS�dXn�vC��S��L*�<�g�I���x�,�Os�O�̴ =��&��j|��6�!��u�&�����$�4 �g�2�<���[ٰ˩v����L�ae�dB�xa�6�l�(+skh�;���_�Or&���T�_�^ە��:{�u�ujhL#-	�{������Ug1m/��lk���]%�))�.ƣ駬|H�̨��Fx%���A��Y.B��).��}ޤ��ju���@}���S|�9}�6`�:6��JУ�2��5t�M�q�������u�Ô��k�@�9�����8�JSA8�Z���ߟ�%�ׄ�߂Ϫ	�%z��X��.��=V4�K,guL�uޕBK�e�;4�="ђLz1���C�p"�Rx�O(�D��?�c8�j~촗�Rvԡ�G?-�#b�]j�.�AMx`_�j$��p�G�ω�u�1/j|�T ��\���!�H��K����e[�m[V�0c:��m�#�|<�0�26Y�й%�����L,2!M�z΂��ǲ�i�rH�%�7� �BF�juv�"a��!�F���Fъጏ���A	T�_�:
�n��!\��=�[J4�W���[H���G)�}��nn��1 S�K��~Ʋ27�~��C���3D�����q�J��?���ҏ�]��*�YmA�{~H�m���o��FyS�%���� �ʕ�����=�6a�vy�=�n��3����Q�[��Yb@�hx�G����tcb��Pxpr7�/��R'���ۋ$������I�8�6(������%Ⴘ�v:S���W��R�͹(�&�P�]&�PU��sZ'b+�vg\��BL�;$�W�*?mv�Nw�i����m=Z0�Jm�Ƌ�t8�J�G�xhmQD8.�&*@�J%%f�/
O���Naf��qt&����e*��k2xN���F���s��S�]�9�$�T��^�g��#�T���P�_�0���xpp���˿���R-��KD���|[�F��FAI��V:r�5&��6&��W�5�!����8������J�>���4g��e�1?�֑/�z��&�)��r�x��0Ɍ�{����C��N=)!��w�\��?��	D�䵠�0s8�w]�;��'��4�d�G��w�D;I^�M
J{u1{b�O8���G�|E�^k��l��*��'s���me��w�15�8q�WG��GhU�]W�e���W�0�7��3Ǯ�c|sDU3F�۫6�N�G���[.αRUڡ>�jAf7�|W����o�Mi~��>��q��������z_g��S�]&�Ϧ݄: i������F�6'�v�	[��f6+���MeL���6ǅ�/�m!Q�fh@\�����#�����+��
��P��� ��:�6h�<�����E����*l�|�3c�z��')�Ю���ޭ��� N�Q�� 1�^(�g�AY��h�0*���Q|9��=�<�e��!�6d��а6Ѻ�m|�높��
�i@l9
`�k>�ɪ�1r�wC��g� )��
�.���&��IE���VW?���0�˵C�tAZ�B��@M_�|���I�A<���K���v��@o���˒<۔�����f��jǘ8rуf))��d�uB���E��K���n�}c�E��nT�+'�%.qa���o�����6�I��y6���k�����Q��b��	+4�d�K5H�\�f5@��a#�::0�m�O�;f�P��=�	�f���s�FS�CE����並�
�]ߋ/����Bo��1�$�h��^,[���Hcs7+�.�=��<�y>	`ѯ<��m�qB��#���ޟjp��'ZEiE$�K���J�8����sf"#�ZiPf1�3�AC��`=}J��2w����B�1��X8TG������E3|�&�������Fֆ���o�`����^��t��CP�H�,j�D��tVlJ��mE�r�bP~�.�)�� h�J�H����7��Ϩ�@�2�0�t�.��=d�7`
s�?���wZ��s#��>z����<����6㺖��H���a��c,�U�a��2h.�~8�U�Q���a���ɴ�Cu�	�*�3Y5�al�Ny%�4Ax�V�3�6���dK.�Pih��Y�KT��A@okr�l�7H�� �A��K
����kXA�C-�rY���}�d�~�P|��Ɂ���s��qNF:,�w��ɒ�i4�}����T�c���L:���ow����}��@O���L�;�'u����(���