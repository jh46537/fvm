��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�{���dʂ�V(��p�s�0ZI��q������N�n�v�Ѣ5���nJy�ql��l�8�6�t�Z�DLg���#;�����O�2BM���Or��m6w
���db�,�}��`����o�z�7L�#�OhT�uGl���~~��g'���|����e���W{�ݼ�}�b0�n��zgw�����0�I1*�QǦ�I��ߛ{��ܽhr> f�$'�����ٖ�����H��77�I�˦\G����y
p=����f���ڥ櫘'���X�K�TP`�$�m�n$��b�!˵44D���x���G<��q��Ɇ�:���C�ݎ��t�ӥ�:Z{s��E�ڞt��y�V��X��d����Ȏ��ۛt�v��`��;&?�˧�dSZ�D�m�x �q�}�:M�p��b0v�a�т� %s�ގU2)��ُ#�Q���5�1!K���G�;��T�"�㕒�I����!$�c�l%j� ��\�ԡ
�.�έ_�	I�ag�ŷ2(�[D]Q�c�����c�D���#P�{W��"1dm���x�S�� ��ŵ��e]6�����u�Il1��4-A%$U���z �� +գF� mH�<@��WjO43h,���l�T��ȸ�4\`��q�E���wD1�Vj�cꭎ5�[�*@P-et�r7���`o���o.h=��wU�~��O7߹�� �&�n>|˷�@%�X
%��y�F����|�s���l�����Jp�����7��G��H ��F�-Y��U�f�ӥ~��9�`�@!���(kx�Z�%��!oL�ҒlB��Z�k hu���iH+G��[�����'$�oO���1��Y�;W����I�}�k���h�X"A&��F�-�T��@���,�NJgOb*F��kb�4��o[�`�{FT�0�Ou&�yCC�.�c�ϫ�iצ�:��v�:��Y�i��t#�nG��!�#[�>�'bV7�0�a(�YL�d׉S�p������6S��;4�]��TbD�-ڑ4�}��ԁq,�s���d�7n��� ��j�. xjT�vOk<�y�H��  �r��M	�	�ݐ�[�'vö[@q�Q�E<ԝ��Af
�J'I��Z���
]������sk��&X��l��r@�I�4<zs0����N���`���Y�ԀU�����x�N0��<^d�V겢~���b���zOn3�xvC�i�X��-HFt�]��1�UN����p&u�A[��[Yf%�9���dg.�~x��u-B��\p�!�s@g�����1}G,��<1BU��58ƞpT ߙ�a~ȃ��m���:���g�E����v{ +D�q%��)����c#L^?�<@�zc��T�Q]�B�ۧZ���l���y��O��C?�)byȊ��J��׭d��#��&�XQ�$|?��j��>�%{�/��o��o��{n����کB��m9x9G�s��-�*������1��[���}��Z�DD�����Y�����TDS�j�L����n$zkBf��
��7 ��	�(R�S �?Z����/	��!i$�����bU�'ͷ��m��M�LV��MO������nRhF0$�
����$��e��s�����GK¹���i�	~u�Σ�8�nr[�Yt�ţ\��HL81r>S�F�Ϟ:%�������Lt�a�jLl��<+�6�����9��)r��5M+Kp��͗��i_��YR���`�Ir����D66�NIw$M��]�ۺ�0$ L�V��E<���s�:s fS�А=h����UJ9�W�	����^�9��g��ü�0Z�L�&�2��K���G̦���
R(_9�~�SU�0_��"�θ]S�D+{a]��`���& 軋��+&�`[��w#|G�)T��E���**�!�� ߽����z;o�C����G&�Dl�>U`�4��#��K�'jҾnV�b���\w��P��)����P�}2�Xq���qNt@h(�}���-<�U����TE���\���J�� ���B�07�v���h�V\��yqJ�j�6������A���C<l����l�Ud$�S��'+��L}Ƴљ������e?��EՉ�T�U!r��z�3@�������eߊ��?��.�3EY6�Zn�����!�^v���h��mHr��mj����.�3K2���Q��x*me���fm/��8L�؄�7ll3��_�2�6��.��g>Ԍ���s��V���{�װ�^��
�m	�{��}l��;J���[6�o��	�G�q������=�H��a�QB��B�;����9�Y-�gY��5�x�Y�n2m��A��۴��p���f9�kji�h�®��p�6Q�G�
K�1h������N����Y�7����?Jlxt�o�oH��R@O,��'4{f r��ݡ����k9���!H�`Ù��9�pU/�dƍ�|�R���$�#���T�#���)G$oƃ�@:�ȵ���+��v��pi��\�{^�{�J��@KS��o���6
C�'�I#��.g+�>I�T�2�cL��x|�?�s˦��F;n5x��_(�V[k�p�E�������{��B���55�����ݫ��e(�C�4��������1��Y�X��Gw�d򽥻����0U4��-mbǔC\Z��j�~2q�)�PO2�w��17M��)�V�,�����^�~}�Ҟ���<P������g��H���D�}��t���g_9Y���U���(��k5* ��k�j�Frsk-�_3��������2	V;j��)39b�}���d�]C�8����w�ݶh0����Q��0�.Xt�mi:ژ,`ǅ/Mz�����)�Bd"��P4�ײo��A�������������Q��l��Cz�&-��yW����Q��ݣ��;���@������w��b�$TX�@�جey��3�s"�Q)�ۏ5~�"/�_cD�7��h>�GϬZz���	�I.��{�8�E1��3�e uNY�J[>�lP�iƩ���-Q<y���$j%�޹�P��mco)B��M�|z�V��)u7z�F"��K<,Q��+<�IA]w�a|���֚������l/������c�ic��/+[��l<�Y�����$E*g �0ܣ�
6QE�H��E���Y;qV�`�Ճ]�E ��ګ�@N��7��?��P��-0=v=�
U�Qm���'a�L�|ng"�HA����m�m��_I=��4�8U��$���~N� �c��=���`��:�s�����&�|�td`S��9�f7��&�;�'�1�+�I��V)˓�i��w�ݸ��r} �� ��q���ܾؕ�q��,����Qܛ�P^��x�?K!�cЪ���{@��g	,��S�#k}2�~�Vs�a�ձ��[���F	��a��\�_~�&I>���Wa����a�5�3����'O�.�`�Y'LgD �IO�ќ$o������'�uq��8�G�w�X������.��Z�%C�=�r�¥�RʄS_���I��� ���_�EY�tNbO�Q��QE�{����S��)�������g�O�p�M�"F}-~Cgch���m�dx|:ӏ�`3��đ�*�]L��3�f��p�aDM�G߾z�s:���k&Tp0�0���7�1�e>Iu��������4SJ�/�x�].�ϿR[�Ƀq��

�����8`��J�L��fqj��Ff(��X�Υ:���B�]
u�l���I�[g6��G���9���4�Bo�j�i^デ�V3�Y��TG�*��������eի�
R=�H�2^u��'Õ��St��?0�U�5Mˏ����ǁ�X�,̳�2g�Ve���m�����$2�+�(
���J�4��TR�UG��x&٦��[���/��/Ę�����n"��`I�۵[��ڗ�CI+Ϣ�'�j��w�|�/��8=����::W�1Ī�l���w${���;w���l,pw�:<�CW�vM�i�P�َ������w����0���(����	ç�D�E+��ŐP��F�����B��.W��H�_>8w����/�U�m��)!If1�����m㤋ȓ���������<K��ݽ�uq��S��f݈�%�]���6XVV�_�� )�4��a�ь��
5����|���|8�$P���<`=��3��I��b�� �e'Rs�v�0`�?bw�L�}9O[2��*���@Zd�x�-��t�Ęt���]��pf��]A��@R"p	u�+˫����M��ّ!�)�ǘ(���� ��Τ���%��Bwm#PDw�&|��	�,��c�ns~I��YB��s�^m7��W��ؙ�M��i54�����Z�/���<�ݶ�.ř{P���=�RBi���e� ���9��ny$H(v!7,�Ic�_���D���e,6'�	��	�n1M{/ ��mޭ:ߊ�S�+,i�tCɮOq�޸䛐:׭��ד(?h|�%�*�n`ܲ�(�0cz�F�Ҩ���}r٠��E�Y�k�p�3H�7�
�-2�gE/e��K��H�sq��n�����Ş�_(J�� ~��u3��8�=��c��8��j8�gT��[i�|���_#�
_v���w�z�@��f����K����SW��U_�K��&�`�2e�k��VnYاW0���+�Ց~��؄��+ߚ��7f�aO�& 2����4eW�ea��E��"�;~*�f<3�����٣H���ʥ= p����*w�/s�&SC��]ÃX )�.�J��~<���=6cj��'�榫�>�z%*��	��-�F~���4<+юh �1�z6����Qe�i�@����''(NM�7%(�o8Y��X�E4Y[��
�&�m�S�y��5�9�^ޕ&�<��C{8�)���YZ�����y��0͋R�ޛ{��j�9�����v��ij��&�xZN�U0�ڂ9O����?A�sQ ���Gx��;��T��}9�c�� �z��ֵ',�
���]LE��O��H�UEk�q��jo��O:)��0�p���2���pJX��˄@�ygiI�;�t��֪�����i���ыu^�$�RuV����ˌ �_U�����=@<5%6�x=�a��.vĮD�nb���9��]S�7���<�~���Bx0���3��2V�մ"7���T��jn��~D���0��B��b�c���v���@�yI��>+�J����؞ķ�|�%A-V%rt�,�����EC�I�OVd[�W��yn<��ye��Ck��e��qe�t���q�Ha5M�N��1ә���^�-dL$ڜ��w2i)t��꓈�s���I�=�HW#�9�"�s((y��V�b����l���\��5Z���L��Z9"���q��~<�bxG�^ h��'Um���!��\�d�i��v�e��d�1���>��_���4�~`K�n9Q@!�6���N9iKn|<�=�x����$p��%��2Nr,�B\�s�=S�R���������B�ѥ��aEeH��)1)��Q��M�8ד��H�U~~O��������$�L��%YR�#\� �.Bm��