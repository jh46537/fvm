��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъ��Sy/�р#���}I1o���d7@�m�I}{�(�D.{x G��<
W���T��%���	w�6
�����,���n'x�ɕ�'�*wn�1�=�f�����,��/N�D�`L[k����}fQLtw&{��q^�7.�>^�1���:��-z@��A' �U�M@;���'�u?i_@lC���8c������n.?��c-��E�=��{|="v��?���ƨ�d���o��l�~�B�aB�5?B��9L�a�G܁9,�S= �������p=u�9�˭t�ˬ��s@wզ� �{�z��<!�:8�#������潥w[�M��h!�+ͦ5�d���u�X�BF^4z�����\P�S+�#}a 1e �M}�ܰ�����1q<Sb+�L�����<�.���3��ȩ��PkB1g���]!E�0�SX�417
�k��Z+!��}�b9٥*���a��dq�8���Ck�f=d��MW�Xj�,ˋ���&�8����>q�-ܳGa'z��3N�7�M/���}0��@�,ƍ�sw2[���xs��ղ��?A�J��	'."�$��x� �m��I�A�o �L����*��p��D��fY��{���w�P�z]��ͱʳ*b~d�'�@A�6�]��$W��̣�2U�D�M��c����9�ܥ4+t�s���]Ҥ�.�[�d%.bL@���ZđQ��n�"�e�W�&����o���z=?O)`$[}&>X��)w�&����Y�%F`fZ[v�9(?g��6$�=��^ �Q�		�q�4�`�����\�b��?�5cyem��i�
�����_�Gj��aii${����Û��΂��l�o��1�[b�S�ؚ�Q=VK���տ#���u�5�+�׌͹�!�n�+H�OR$]��M���T���Aj�Z���A����{h�fs���N�a$T�w7K�Vװ����z�dmjI���묨���>�}���Kִ3�z>��k�����ȿ�0RYM�$
P������p��$��<��]"m�w�8V�X����`}��l�Ц�
/���z
�b���jdBEHrh��ћ�>�����´���f�M���!l�!$�,��a$�]��G��ȿ���҆�:��Ug���o�r�I�����jQ���}R��m�* aϢEk��\��O� ��W�p�]:�?�<���n}�xŰ/����]F|i�y���:J�f��V� �uY2l����X��H2�Ϟ�	� ��Q�1Z`�����RC�,`�n�))�>*��|��E.�//���t�/�\�sП�I&1\ZҢVUS�X�$b�\�؎ :�xp�߄�&7
��:�>���	P�Q�믜{!pz�-A�SdhzD�;�zc|�����Q4aӖA����VH��zju�-@,i�u|�sR�iW����1�	s����6U*i���^��dZ?��A��;��N��D#<xfc�nC��"�ɟJi �9%p����Y�w{~{��G��j%7W��q��v�}�}������<W�5��ԃ߲<�b;�]��b�J~�ȅ3^i	�XL7k�cB���::u���o�3���E�l�44�&L�*�+��v��m�U��ߙ.ٝ�'���d���S���c�r��QQ��c�q��y�M�U��t�:��L)����I�K�w�̀?���&˜B(��Χl��Oѭ�ɒ���"	ǎ�*b��=E�c�A�=���U�>.��KlT �ᗺ��pS!�Oŧ�d*}I~���[Ar�8�0?�D��A��W�O�`��8�N��Y\�a��~!��}�Ik�N��b?�j;�ʧe��O������m Bc�\��K^7��U?���@�t�03�?,���L�CB�L ���)y�/��W�U�����_k�ɟJ�2e��υ��ۜ����6ex��C�UN#�*��0�H�I����O�]gx�L�*�8g@v�|#�F�-�h3W���?Q���"�A^X�G0Ʋ����� ��Z¥Hcy$�@I[�Ҍ�e/}(��U	<����`?R�w����?^A�&�K�MQ�77JQ_j3BQ0-�g���b}�k|�
SM�y�	�<XQ�u�{$H�6o
������9�⛾���Jd��|���H?�$��I~*����"�K���bw6!�%��'�3���k��u��sİJ�Xu�\ӡ�r�E��Ӵ,px��n9�J��e���ȋ��fn��Q ���F����rȤc�я��cS�nF� E'	���PM��O��6f�M��LR��>.�r�fY�Z�� 4�撿���w:�84�Ʀ������2�BS7��������7m!)����#dP�c8��t����hAɧX%�HX�·�䗍Ϗ��/Q�|����*���}�Uq��w]�k'���>�=�\&S(]��Ǐ+��EH!FX,5��^��<聈�	��}����a����Mpw�WD(��5�ΨO����)�5:r����t�����B#��G����* ����p����:��-ˡ��}8o±7�8��/Z�"A���Y�g0#��~^:\� L/ڑo�,� Vw�6w�`
EGX%,�3�5 !�O�rD�\�m���P�����;�t�8@A��(m��oI �+��)�f��E������'yn��@��6.��濏׳�P-C�^ݤC����#�sjU���9ȱ��`��k�SAǿxK�b�:�c�T�`E�~0@z���v��:z�\^O�z����Hhox��u��j��h-���\*(�|H�?����4�k'��(��4�_��~U|���/6�(@_W͡�z3����R�`�^��#�P&$D��)$��b��x�DNl��@���g~6��K�B��5���"֗'�)��0�=��	���%4�Zr�<O���8�-���������?�S�d֐��S-K��k��I��J���,���Sa���Y�(wr�o	�:{҅uP�|� JycK^���F1H|����!��5>H�aO�1|?I�Ç��e�>���1/-i|h�WQ'�x���~~�Ο����y��%ۮ��I5;g�c���9�eg��x��0L�F�i|D6��5�(i��5詎�����n��S%�����:h�D\w7��E!+���h����h�d	'��:z<.�gp�5���&�y�?���fF�Z4q��YM�y-�XBKB��΃��R{��S৮�f䵍c�  ! ��jv��2"�F�1���^��zd�I`VQ?��fn�J�yl$@�,A6���}�@/6�|wb���h<�R��c�U$}E�[�9�;�KK7P�4e�U��o ��q͋͘�܌:��R�6t��ٻHK6�FS�����6lf[ȽbΜ�"|�=0��V��{5<:'�g��R��N��>kK:��D��୬�.�j�" �y\~�)�
c/��f[�t���C��K���*�����rܐTayf����1�����."R��"�T �m��Y��ݏŮ�!��ܪ��o�VMN@����"Q2��}NyuX��~N ���^��x��W���A���k#�gAYa�]�B����%��(($���<��?uV�R�q�O:*�<Fr�/���$���<,c�l<\>`�38�IL�A�JgI ��46��+qw���Tz�e�P�ޤ\���߬��V�i�;�3�����Aװ��g���CmJ���i�5�:n�������YZ�� YǞ�-ǆ'��pǭ��d#GŬ���G�E��4_%�F �Q��p8��6��
;8U���>��Z�E@�h+q�:<�Ɗh��i�$���-�'����6ؚ	^v�.���m��&�r��ǳ�dJ���x�ݟC����|V?DwT�-A�ٿ��2q���@l�;�Ͱ���{y��
��[1U9ORa�2�_��
E6ZH����i�{Л��#yT1=��������=��/���	T:
e4>΃�.��$�{�W��Zuq=Up9!,��{�8�A\�E5�t��������&X����CM�� ��>Ѭ}�Xi堌Tp�AŜ�NN������r#ν�ծa���՚#kЏs���~Sd�aA,*_�B���$�-��@����(���K^���ع�_�kܸ����mN��M�����g���@�5]�������Q�P�*"�	���^[
*k"n*�I�ry?�^?�� ����n�ݘv�`|�e�}�Txdn5������K`�M�s�[���-Y����Ҁ(��T�������g>����R��~^C�%�L2l�'FB�mσ;��Xm�
u56s�>�w��%L���
P3�ʦr���S����3���̣t�EP72ڕ`�xY����~�XZ���+KN���e*��Pa�#���j���(n��Zo`j�����/Z�Ji�}�RT�c�O���ݞ̕-���:x��fx��Sԕ�#���y��u��[��KbLe��א{���	Fۃh1N�V��a,�i�X��$dw4��t���o�6�@E�;�ů?�&��������1d'ġ�ʢPvW�&���*�*��]C_���u�S󢑞�g�s��|0��i]�%�c���a�36�~Oqtq�엸.��"�Pk��j�q�M��b���1y�wķ޷w��SM�2;������FEv��E������r���O /��_�<������M-�|���@L�S��oN�a;��5�!=ʼK�iKGD9�ֹn�'E����=ib�ی� o �qa�~�'�s�[���'�ɽ���3aZ�r�����@�Df�G��]���%��ӽi묛��Q;�5���:��-���߱�����,�<�)Qmx�#���
נ@")�3b�Ƈ{v�KF�(1i��o��ϛؑu���.Lo���e��{���u
���Ӏ��8`0��G��5<�	�uV%�zʽ���4�:>����� �O��*�J��S������= ���AwFD�5���u�B;��%��ڪ`ks`�����9�$��S����¬{��J������� �$���`��3�;�5a� ����1l�I^H�&e��#�I��Dt�����yaB g�>`�L���-��b�-kMI+R�����<A%ˤ��1��B�Q�tD�V��b�%��Xi��s�,�/r�x9�i��J6����1���9�À�{���J�(���N�q��1�R|�N�F���DV�|�,.�����F���	i�Ĺ��k,���i�w���ټa�?�۸�!��/đ��W캟O����9�_���5�)� �%��ލaO��1��P�^�����G�G) ��D��MVv�HSdCaʂ�/9d��h������E�XCz�KU�)"iF-)����v4��ȥ�jGN���P�ׇ��I>�p�y~�pL��b	�����}Q��O����w���xXm�E#)�u�v���V��ڽeG������yVyl�v����KL��⑊�?f��>����zX-�Et�V�XvK�0{���G����C��&{�{7��9�|�(%�q<i��͇),X�+8Z8�z]g��Nf�6��ڂXpo�F�Ε"�#/+3_��BPU��wY�P���6�lU�Iny ��bra�I+ �n~�z7�Z�F�:�V��AՖ�M���H���Ӱ�S�f��ݍ^3��F]Z���FnL�W�^���ܨ�}j������ض�o��� <�k�_�o~�/� 	4)��REE���)͕��B9�"n.m���h�?<�?��]ͱ\�͝�ኌY٠#�-�����N��l~k�r�e�`���~�ʨ�~�xn�'W�%������ ����1�A,���N#}��V5����o�Z#m5o��#G1����l�_���A��b��2�6��w6ynMm#E�@�
-g�/��	�<�*���[�9��Ce�?���9�c=�a��&TUid�P׌P�oK�my�u��/���SlH�o���%�b_H_ЊDN/G�x��F�����j2�y</���4���A��ѕvT�;��h�{�Ki#�
�惀yƾ���C�cݖ|4��撣��ȗT����P��*q���d�(]�pS8O$Һ�uKl"�K�/RIu�s�R`?�|T}̠��nTo��}��f���ޛ ?�������"�qz2��U�P�-��:�PX�Ay�!"lcM��*����.�R-��o����Km�8?/��]���0�3�S�|;lM�K-��we�Sp?��Wލ#�z��������Ej#3�B�#g	��܃�������G��wMѻD��-�9�M�!#`��T X�i���T?
3[|�Կh�@�2rT&����Vsf>~?'��lf������"p6����ZL%F���ɍ�B����G��0���_l�v4�u���O��T���a�9@p��k����*��cu$�j2/��`�{FQ.��N��\,ŗ���T�-��j�(�nT��OmZ�{�Ʋ+K�ؤYJ�N��U��� ����Lk��%릉�zV�_dK"���7�q��F�V�F~����w��Es���)�+"^p���}� :>����Y=c�P������o��s�D8\�w�S���{�=��B *w[B�P�bj·�㡁��o\���x	[�ji�8w�ζ@0�ܲ���<_J�Um�
;V���R�(��V����ǎ`ו\ߐeQg��i���h�� ����������o�$�W�5�${3u��X]89��6?�뿴�_�7��9�$�X����'=�>�_���3Xa�5��T��	��h��ٰ�y�FȒA0�;��	$}�S��f�s�X̃z8^P�aRj!{���-+Љ�'1��mEw����"ک⺷�}��!�1�s��	X�.IF�NVո�k腮oױ�鏀��R��
�%<H@`�H��,|*�Ż�d��ùl��'����;����AO	
MBe�ؕ·��m ���8���A���{���(q"�^�0�ʩ�W�2�hr6���lW�p