��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\Z�;�j�A�D���£�d����2��<��.�d��g�a�9`E�H`��O\T��<�MuYj����/�m�@��S{��]�q�oE�@>mo�����]�w�Bn��+�ʶ@/қ�9��d
P�G7���Gu����XA�W��	���U<�^����me~��+�Ђ�U�b�G#���S�m!�vj��,��Ά�������0b�����_TJ(UwY�A 3�~��b��΃cY��7�+T��bu��oӍ��P}�Y�X3��"%��^�:$��P����W��]�&q��U��f�=����S��r�i����4n-�e�
�/`"B��s�������0��n�?�����3��?��t���?��S<(B��Fիc�eƥA����e��3左�s�^��W��.J�J���0����"�b�^G��JWP�r=fEj��{�Ѷj$�L�C���U�1�1�*wu,u��")8�d"zXY�a+�ٸy���dl�[R�"��	+4G�u�s�ωrR�MVxB�F��$�1&�(�o�K���Gp�F�74������a�S�Ϙ����P��iR�'c4<�	(��#����rK�8�\=����Dܛ�x�!���#��r�Y�'y:s�i��=]�1�+Yl�ΠY�ι��-��u��y"��I�h�wG��b3��*}�6�m�cUKS����§��4��8K1{+�y��g�د�1���;�0-6W����{U.�rU��z�<u&A#�<1��D���OH��Nr��I���-�*��;���j�Z��B���������w�+ş�S༤Z>uҐ��c���+ԅ��wL�؃U?⚓tATD�� M(@�&�/]��[�����#&e�:��vy0��p"`�Q"̵=N�22�?m{C2��8�믗���՝�!�̼���ʌ��>����l �d]?�CsL����q�D�%�K��%����T~�������@�/�D9�0wA��3��[�j����w�
v�V�>�l�y�\<�Ս�s�F�Ih��ST�}-�uȢ�yA���I9F�WGh\;v/ϸ�ꪝ�E(�MsA�����#���H��{�0�]����+B�����l��99���"����ݭ�]��V/Yb�oj_��ҋ��cDD����q63?N�6W��2w�7�`.�-��M�&aW��{#�1F���J��&���F�y����}���nk���A&<g{��Ibh��x�o·���y���fH�����e��k��"�+}���l8ʶ"7;n1�F$d�Dfq�$��<qbO��LtP�a��9V�c+H�J���e������0De'�Ȁ���r��^�v�X�Ѯƶ}�N����l' jc��F��:��4JW2���*���6��*���A��>����?��м�J��G#=�]�ơ����!��k�yi�n�=,�,yt���I�z��a�Kn{�p����9W3a����J�ғYc���J1�����&�%׳$a��B_j����M"�
���9o�������%QÄ��	�,;���&�~�.�wU�._��b��O�S1��ٲ�ּ��+�+r����
��D �DF!ra���f�׾)�.Q�T���Q�q+��L-6[��J���V�gq�?�� R4�t���)!�'�d�Z�ł3j��2o7Z��Ạ�uN���u���GhB�0]��Rp"ʄ9>VR�����@ab�!̻vt��~(�拎�����hñ���Ҍ��R��P�h,ªL�mS�E����Q�BF�n�\��RN�?!y<A���!�Ŝ�G��cRx~���2�Z�~�a+;c�gw']X@�E�<ܥ��oT:�)���Od�Nʤ<Q�`x�?������)q7���F�������!��� m�t�x��%�r����1q9��&+�3$���?�Q�Mu٠��CW���G ��K��.�,����8e����>�a���#D�3�ET.GX��Чļ�m^��f�Z]`V��S3�M1֞ќ7��?2������HMí,�.;s��z�f�v���H�Lo�aY\n�G��% p ]+���npj���g~��蒯ЦZ|��9��]����%g���R/�O`���Ea�
d�+"�����:��e_/w!��ܮr����g'�Ja>�0Qv*����C��W�E��Y�?	i&�iB�(���5~��ӎFڀh�o�6P 6��G�y����}���-h�o h���0r���t�R�333$���М�7S3�y�r�{G{	�a�QrN/ ��!�:?��J��������}-J0���)Ʊ�� '��N3�;v�9����(h	��\�R�@r��t�d��۔o�ukM��Q�0�g���l��KȻ��ԁx�����)�l��E�z8GF�wO�%fǚ��?4ax�6V���c�U[�*�pd�b�'E�dK�J������m8����u�����-"�������λS�I�f��/3<�ѯ�3xN6W��8D����BOU�;Q�9������T!!���XL�����I�!�
a�c��)z�1bz��{������<6�j�TJ��Ԑ[����HAT��X��o}�V���`�|����e	�V{���D�G�9'�W�!�����@�C���a�qU���054MwG(Z�Q�xw��ϼ����1��[f����L��Xxw�YW�5�#Z�K�"=tB�xY
�ba�Xg��k��i�Q�H�IRy*������>�Y���j�D�^�4:��5]"�>BF�s�bo	�p�vWJ_��4��2��
�Ζ&$Si� g�c.�u8���n�c���Y����y�E�#�_�����>��)���6��NZYYF8_�}P]��i��҇V�˫KB!���'��,�f?�R�8_6�_�L�3N�X�a+�
��M��ϻc�tn\�H����6�K�h�� ���+��qs	P�����3�#��˼Y֌2�t�/Ob���Ϸ�̩�Q�_a��Cf?���6�x��%\��e�^��!�_S�c�ܤ�GVl���g�&L�3�|�b���8������$�2���'��ˠr��Ͻ|�e��Zm�ٚ[��<�;Ju�*g�A����*�p����<�&`"Y�):����;��w�/tڑ�/����-��C��.EC�W�NB���@�S͘Ba0[�,Ix�8d~Cb���@k�jlg�2%�nH��U�i�ㄌ^A���	p�!3�(��׬�o�L%`�S~�u[�4c{$�ϟ�!�{S7�V�R��&��#�c*�����Yʆ{^�
�HQ�aͦ�j���80�hX�����}�6�����(MbX>A�eU_������yW���ͷ�w�:���MQT]���sp��9�����/K�H7���`J��]_����x�W�R[<x�" !�ٓ������	f���[�!��
�!6�g�8�0t��~�~�ML���l�JOV�Ț V���i⋐��h@�:�3B�i��u/u��N0��4�`���Ľ"Ain��2�T��M��~��ZԴ�i��l�L�.�.��9�Nf��O�^F����a��&��R	5��{������]m��;N�'<]��~���F{���v,�D���͑x������+�r"���W2�rԞ- X��P�����A�]�i�����>E`Z
��&	]q�s&��Gl�#/�6�#�I��Bz�y:�_��fpc:u �|m��Dig/;n{�_��|J���j�a��H�/M!=\��s�5!S���ܠ�z�����?{�6�����>}�yֽ�5���}�z�5�k���S���4�#
�Z�(�L9�L�4��~�V�p����T��\Xi�?���r�ø9v|��y��<���t]�A�A�y�x�փ<H軴(S�We|ŕC;�B��#��`y�νN�� h~(���|�A0�!�L�f���D&���������-"�¯l�0Qk�U�-]�8H�
����l��orX򉣡� ���M��"n�������4/�T_�g��`*��z"0�yן �E�F�tN�4`SU���݅Z���⯯�p���;C�&���d�-��h2O&F+똓�I�&F[�s�7TuJ���f�ح��̀�)�7��=�FT�;Λ~��R-Q����$`^"O�N�4j���r�4�Q�G㪴�mT$C~��EM���h�qw$�ty|nُ3��g���KDi��ܖ���D���V�)i`6�UR��v�
����l��#�5��*3�tc���^�(��u����v��~��p���[��ۜ�&��V� ^뚼�{�GM4�|���/�U�w:�KtsX���`�����8�Nv�����a�����45�ɝ���6�&��]/6�S
I�?���M�����.�����<'s�c/���`U�)�x���ƴ����tY �mCʼ�;XS[�ͧ�,v}�U<�{���R���TN�:��Љ�6���G�f�:خ�T�%L�VY.�ԛ�Q��}ҍo�
�:�.p+���66�B��K���ٞ�T�h	K‽=�.���rw`��oh���+Y��n	�
�E<�Ƌ Y(>4+��M\c�$���M�Zb��Ɍ���l���VM�	Ъ�`��r˰)�����#�%���U�5`�էg��`���g��9���:��?�����$"�𥗩c��j��w ������D+� DB?�͐.Aa��HX!X�E/^w�KG���YK��1�$���Є����$�#;�'`�AK�E�e��M%�m�˻�&��n��'��W�>��P;�a�,����;���pi�'��I���iW0�	�'P�G������
��QD�	0���O��-;nL|6�|8f���? ��2=i�p$�ڤ�*� ����:�*[9��z�8�z���z�s\�:Y����뀧h�u|���7�7)�F�)~�n�Z�a�p֬YS?����)��z�.��
��
���^_jYa���^k����@�3M�m�x���ڔy�I�pX�A �� yEd�ζp�{EҰ��t�H`*o'�ƌ��7��$o�|~a�x���v��	����۾]w�R�p>C��`t�lP�N@� �^Р`&@#v�Q	�Ĺ>K�H��S����