��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���H�ي�9�c���]�uJ]�u����`����#������`��`m�ň޾�-B0� ā��q3h>���gw�HQ�#�)�>�>T �P9�i���̟Ck�xem2���.	o�ע�H��-f��r';����v�
l5V�@����F�n���}F[K�t��}D��ʚ�����N$�E�K���C�0��~l�a_`����z�(��3��E0emY�c�#ZE�xv7&�uk*9t�bB�#���IC��"I����> �XD1��`?�M����$���[I+�0gS[�D_e�R�i>��j|�S&�~!�U�p?��>u^F!D�{Kx�����NyB�uѴ�Vjs$�ax@h�eف'�K��~t�����I�A��'ښ��e6�#��a�,���{B&+I	�p�S��.,8����G���0��`د[�!X�P ����h'�+���F�,X��[z�^�B<=�TH�^<-�_&�L(ǂ����v3;n����� ��
���A���:�3���\k�D\�sϩ���3 �C%�.W�Ԧ �}�{`�r��I�h�3R����������j��y�Ҫ��O�o[o+����F�
����w���P_���C/,��-G7�@��s��n�?>�ڣx�պ�������X�<��y~����|8"�qizg1���n����Pڱ�?"@�7@�L@o���6Wػx��{�UF6Q{m�����<8Ѯ^�ROQ�q��Z�@�{Z4A� ��C�U���U�����������+���KY�e���X�Q�6���yP�;(��`D*�;���)�Ѧ�h��[M!�􂅏�y���~W�nO���3b#_�������Y9�Ci���3�r!�9����1�#  ��fc)\S� fPt}Kg&��bI:ED��Ժ��
zI�o��h5޾��Λ,�R��#����%X�I�(��l<-6Z��'��K�E�������/Cda���Δ����b?$$�.��<�pl�Ե/��D���T��k;̛�����Z�� �Y��P���CSKP��A;^\b"�$R�8���ֿ0ߛ�^U��_|ꌽ#�p��5$���i^H��Z�~w5+=�Ò�_�bU-�˟:��_��f��m1��ެ!J�K��&�����U�mH((ee�k�Vn�Z�G�+��kޔy�=D͈��=Ӱ�ŧ��r_���!x��.<�G��MSĹĠ�x3�[��9�Ֆ~If3�d�������RT�����$�EJ�Iմ~�� ���Hq������w�\����*��2���rë�d�W|Qf�q[ʜ�s�=�Ҁ�H%E��׬�����&�a�z��/�g��m��F�u<�uY|�Z�Ʃ��������wRH�ϠA ���R��o�1tM��{R�q���K(�1���[�Q�vۈ��v]�&����A���{���m�Ž�@i��?=����]퍙j�����a���9[9�Ǽ�,���Ku�<w�1��b�'����᛭U���}xK��̰����t�y�j�R�!���3pj	Խ�4�H=�E��ɇ�6�_>M8��R�&��'�� ��yȮ��?܋Y��òTj�f�ws���iJ�|�8���T�:������2����'j�o����Ftj�`�׏�X+.lr�����������}�hk��}O�G� �*���'�7�S��I�ݜm4�n<�J��xH5-��� �p���3�ݪ�O��n7��,�����H���D����.��+�>��vO��Ҝ�6����eQ�^�R7�E_��c�)���׿�@��v0����	`�kj��o�L��	!��%�	��A�%��%s����@X��u��<i;4-{�ͽ�!�=J㑦
�c�
Z���~������'�5���;WtI�,����%Qt��uM�nԓC��6�>
q�5q�;���*��� 	���Ȝu�&�ɭ��T��T�Q�s�HɆ�a{Mp��$���5��LP��`}iq>F�F�l�Y.���W�l� %���>�eѠ���Жu��挿��J�ձdA�\�C7�L�?	 {L q�<�������Ou��8Qk������Eߑ�兢+��߹�p�\�K�(��
�6��]���_�X�*��T~}ٹ��
