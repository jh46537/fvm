��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q��t�Vɨ�G�b:�e,�;<�T������8�l��s���:k#��a ��G��&k2�%�I�����ނ�<��m�V�R׺��{���������_<6���>D������"A��%�E.��n����D�e��`�������v����,`�a9
����c�U�2�h��8���w��yQ/P�����>��.���������q����`�(���q���ڇCV4��ۓr���^M����-�/i��&}.�ێ�(�@�ל9��,c�0b�#Sg��E-��X�!�U�U�Ks�z�kM�¸+XNS�:����Uk��C��C���Hp��R�kE�è�%nE�-�i�\bS����]&�N��q�#�&Ӫ��&�?C��]������)� F"�����B+��U�~�� kU@�:�sU�����^ � ��;9�jz�f�;S5��vX�[X)�<o#��|��=��vى���"ľ����d\�D�8��F�HO?47���"�yZ-�I5A} �&H��\P�SCx�+�7�ݛ�HQ6�QIr�0� &�`t��3�gg�	���'���8�e}-����/	m����18z�b2+y�{ѻ�Z�M��/�bu�GGY%n9���{�R�tTs�&��)<B����h�+
��R>�t�R��U�y�����X�{��M_��yI���do���ڿ�=c�22�Y��\!�o�]v+砩&=���_��l-�v��[q�{ �����X.hC��R1Zi��{8�U��5\�/�@�[���c)*�X1�($��?���<�l�u�#��^��f3v9�S_M�����U��@ƿ�H��#ۆ(J�.hJ^��8��=��`t/�4�_9ͤ��M��*�p��M��D<�S^�n�F
M�焅�M���ܹȵc}�W8:�$H�y+״Φ��]O���۹�b{QG�;i� 0�y�p�8��~�����u�C}+��ɕ�>�Z��FVm�$�D5��%q�x GV���5_��,!O�̃�>�^��a�rb~w�[�@GK	%8<�3�z6�2[����0�P珁����*=F+�+ewBg�8C1�v|c�Dҽ�97l^���� ZVl�X=P�uexZW�Knm��OK1IN�fr]�#<]ͽI׆�.���3ʕ�IO3�dܷ>��w�ۺ����#(�W[JS�|MR��)��������~�(�� �r��4�	F����"�n���4��y��W�Lw���^�%?�0B�g���"B�1�@RZl`�`�D������O�@�ﮒ��E8�$�!��X;�/ �*�����G��3ǛNGpV��`�E��%��WAxi����.��*I�t�5�2����޴�Üs�ލZ�0��F�4����8�ou��o��d��Ԟ�K���";�(��{B}A��	�9����0����x�9nF���$
ŹMX�5�6���$��&f��67&�m.����<[�+�7�.0��\��_z-I��0���%Հi����?�(|��m�'n��U	c�Uj��$���Y��mb�
����:m��՟���^�9��Oc����ａOc��\6�ˀ���0��VA�m5���U�*�$�fa0
��R��� �� d�� �Dχ@6�`d�B�����m���ͨ*ciJ�� ����cw�<5��I6�͎����iU�U,�^r4���D�NM���i2�C�>���;Շ���F<��]?ѭ�fE�nG���m�1�����pc�*��4�o��5��b�v4t;�	_P��Yx��=�M!�.g,�SV�!�ѿr����j�o�VX]��W�b�.mkW�b�?�tA���|��]�߻���&��^��8��^>�uP�㭽�Sf0hȪ����
E^�>�
��6�3��r�Q�]�T��G A��D���hr^cKM�#�-�!���s[�\,&8��D~��Z�U��k^�w��f0v2��L�wl)�Ρ3�^]��,�z'����T����mk�aE�.t[Z��&b���,���ھfL	����_�������=�w����@¬k�5�N?J3=*��؎m��;�?cOQ��)Bǂۼ+y6<��M��j,��#��T<Y?q�z���Hi�k���6�g���ٰ��\0�H`��3΀:�p,g%|" �23��{.%z��IO�b��kR!��z[Ú:xfs���|2Fvww�F ����3g�F.x(r>HN7L�e<�
���>ڰ�#H�/tZ"�p#Q@�D�r�p�9�Fӊ�^3w<�x��.~�ԟ��_S�v*^�s�S����:�b��.�`56J`g���y5+9�OLL��X��Z��kΥ�(�8�	�mj#
|�i(*7����o[�؆�
!@̘Wg��EXi*��LO�S/K� TzU��[:�8�hS,|�f��� ��s[��.���G�SW)R���~�r䭎����k��7����׌_��j�ֈ����d�#kW�EϮ�g`Pc�q�%�k�������\�Iy��_�*��Wf��S�G�_���e;$�A6���.�Z��Ŭ��9!��ST��X��[?Xm�!;�ʡ��}غ9��N�2��cl��Fc'�(�r_��p�.�&��<ܑݜ�YB�$����q5�g�'+�+7n��$S���������B-2��)��	F3��@�ca/G���F̤a
b%?IH���l%I�6Ij�;|��Ѹ�����������s/�rUg���~�E$�(��?!���+JJ�>�@�G���{%���`���Ep��Z	����ϣ�B5�Y�d�&��EG(/�N���z_� �W��|x���ݕ�:��n�P��'��k�"r8��K�؞ک�oޑ�d�=dmFPu�`�5���e�y���as�����܀������K��HW���QQ��m���V�$�<꾝J}��lq�����lڬ�Ȍ؏Ds��+7�
�;�nd&��i8�`����it�0����U��Æ>�`cy]
�
V���[��o�K
�x���u�-�������9�Sh�����ls�'��C3�;@��"��Z�� {���������4��L��. .$�1l����s�d���ߦ���I�+�SNQC�z���`|E4ɝ�W��1��$ ����(����'�^!xx���3�FH�y����
���k��gn��8��)_
�n#|�|��5�@�>N�x'�>[�ۤ-��L��@�T��"�t��ꡣC
�g�c���k�q���*�`B�@A�3���O��T)E�>&�v�r�ߏ<7��0�"��Lo�h�99�.�4]%yRd���s�ӛ�-�];�:�yK(�?&�Gwc�Њ����D�!o��0�P!�d�gͰ�~q�Fɘ���au���7!R�q��"�^�(.���t�y@ޑ�N��x�b�hR+vc�GoO`��_���V�y�����^!��,Ɠ�f����O�&U,xs��w��2�^
#JM-T+�W��KH��;�����F���UƁ+��Z�4B����寷>���<M��Gf|۝��i�uN*������玮Q�d�V;���z�%�!��X8E.�t�u�Z�(��<���3��}�i���ퟙ�8�`fF$����	�=J�s-V�O�Y��B�|��'��q���xD����q��?��?elO8�/��������j
Z^J�8-�]�(�-<����1��
�oL`]'���j3�C)�[��n�}Sicu4Z9%]�sXn�G��G��Y��?{���&� ���Y
�
{��ܹ�������6���ִ�i��B�-ry�u5���D`�(Dpy�,��������D���n1)�B քPZU�P�e����;�b������!��@a�D
%{�ڞYE���|�B����"҄M.��>�D��������0hA�o�1����YYl�0G�X�|�O��v��Mi7w:}(AV�����|�G�������X݁b�㈭L37�zH��Kd��~���.l~���?o_(dU��}>@�dǶ��Lw!$�L1��^����UF��1��<����m�7)��s�|N�i>��^�	cW��d��z�}i����&HE������Ako�0�mD
�[6%y.�vB?�����O*�M�}rdz�n���4�=�ucFx��1%O�s�t|N����Wmk
�� 2���-�3��x=��8ȹ=Tf(�w�j]����m��h�x��v��T��H��q��i/;�wS$,���QWqtR)A�^?ۦ4L����F+��KC�f�EUy�8��]BՉ� ��|������V����؟��m���*J�-�[
(��D��,_��r��6���j�H��/��������k������hSY�U�t��
�	!��,�W���r��!���zFj"��e�pz��4�i=�i�gaϦ��IP���!�r����ҔpX��`��,uhQ*Ņi}QR��ۜ`86�W�n�[*�J��5��j�l�W]~8�85������W|Ӆf]j��z���gPy|i��#��xf&M=c��A��������!�c9�v��c�<��Ο��۳�?�M�� AD�����_>l�G<`���i�Q�&��2%�����%C<���HCt9hO��8-���4��'��,�p�z�u�ð��4�RH2}�|��H�Z���n`-;(x˺�"�,���n-K<a�(�l�,�t|r ������f�?�������K�2�!����A��;z-j�Va~l\Tt��([k�kR~m= �#�����Z�j_��\��=4�@a��]�:�F4�9�Y�j���˨T���%��ipw�+��-���?�+x+����JgG��cA�Q�8���	 |��]�7>9��4'"��)�oA��ʵ>�{�{�Ҹvs�/��� zm^	��0���]�{ӌ[:L<�e��o��f-��u1���Ԗn���Q�^QH��<���A]�C)��El_vd��i��������wL����a���ɀ�|�Z������`������ҥS��%/s�x��4�:(0W�����y�o �L(�
f�Ȭ���J�s����u}�)��v�O>�5�c/����E�{x�5�H`��>���'7�m�F�KO��@n%�����G�?B�M��ל�A��<h�f|�ud���z��U	08��"��ឩ��Nh񽕀)��w�"y��1����۰�&;�&4�Ћ�͎�Y������ҧb,$�铰��x�Q���1j�%��D�Aֳ��lO����mXU��j�l��4�)�ݚ3����r�X�&GU`>cY�ɵ�5/&�m��%�xF<w��7�-�n3�'
�(�h���X���9�|�%�۠����Vֹ��v�t��e��X�o |]4^���ls~܄*mKY ӥn�b�w:$