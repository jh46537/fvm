// (C) 2001-2012 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License Subscription 
// Agreement, Altera MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


// -----------------------------------------------
// Reset Synchronizer
// -----------------------------------------------
`timescale 1 ns / 1 ns

module reset_synchronizer
#(
    parameter ASYNC_RESET = 1,
    parameter DEPTH       = 2
)
(
    input   reset_in /* synthesis ALTERA_ATTRIBUTE = "SUPPRESS_DA_RULE_INTERNAL=R101" */,

    input   clk,
    output  reset_out
);

    // -----------------------------------------------
    // Synchronizer register chain. We cannot reuse the
    // standard synchronizer in this implementation 
    // because our timing constraints are different.
    //
    // Instead of cutting the timing path to the d-input 
    // on the first flop we need to cut the aclr input.
    // 
    // We omit the "preserve" attribute on the final
    // output register, so that the synthesis tool can
    // duplicate it where needed.
    // -----------------------------------------------
    reg [DEPTH-1:0] reset_synchronizer_int_chain/* synthesis preserve dont_replicate */
/* synthesis ALTERA_ATTRIBUTE = "-name SDC_STATEMENT \"set_false_path -to [get_pins -compatibility_mode {*reset_synchronizer:*|reset_synchronizer_int_chain*|clrn}]\" " */;

    reg reset_synchronizer_int_chain_out;

    generate if (ASYNC_RESET) begin

        // -----------------------------------------------
        // Assert asynchronously, deassert synchronously.
        // -----------------------------------------------
        always @(posedge clk or posedge reset_in) begin
            if (reset_in) begin
                reset_synchronizer_int_chain <= {DEPTH{1'b1}};
                reset_synchronizer_int_chain_out <= 1'b1;
            end
            else begin
                reset_synchronizer_int_chain[DEPTH-2:0] <= reset_synchronizer_int_chain[DEPTH-1:1];
                reset_synchronizer_int_chain[DEPTH-1] <= 0;
                reset_synchronizer_int_chain_out <= reset_synchronizer_int_chain[0];
            end
        end

        assign reset_out = reset_synchronizer_int_chain_out;
     
    end else begin

        // -----------------------------------------------
        // Assert synchronously, deassert synchronously.
        // -----------------------------------------------
        always @(posedge clk) begin
            reset_synchronizer_int_chain[DEPTH-2:0] <= reset_synchronizer_int_chain[DEPTH-1:1];
            reset_synchronizer_int_chain[DEPTH-1] <= reset_in;
            reset_synchronizer_int_chain_out <= reset_synchronizer_int_chain[0];
        end

        assign reset_out = reset_synchronizer_int_chain_out;
 
    end
    endgenerate

endmodule

