��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�ӿ�J�fVȖ�!8�a!���x�6�`�P�0�!w���K\�<"�Ԃq�AY5X1�����ו��GFᛧL��Q_�U�� ~�^�n3�����?��l|s�Ҙ�����kfXe.32z�ܲ{;r�%�GH[�%�S��!�V+�*����×Gt�L$L�f�MJ����dn���L�(T�S��e:��e�m˗�x�Y1�Ȧ��ɕ���o:��Xi��H8�M��5/������h�����_���$y����D�,��Y�{%S�ll����)��j���Kz�ÿJR�~a�N�����op����2��ߛ����a&�W�C��+C��@�AǸ�~�����Y\n.�k�P������+$l�7�}�8������k�<�,�m;��6:r�"��#2&��q@k�.@"������,H�U���HJ� w�hcq,��BJ�L(HE�3�.^`Ӊ<f�G
 �-��eʒy��b��y��;ň�z�S�Պu+p��av��� T�ˠbJ-�A�Fs������-���ڏ��o����xk3�=�\��|W��7�vQg	�S�o�ɚK5-X�G��~�Zl��d���ƠS�&�4��=>�g��b>X�����2 �����ݯS�Zk"53ن?��8���f�E_�eîou?R��5̒����03ɵ�L�|�ɀ��z���\a Տ$/S�u�r���@�@��4�֗G���(�����	��Nָ�	l�S���4v[�%͆���<f�zf�7D�X��u��jn���JFF3fN�I��J#�uN�t��B���B��~�+�	VA�I��[�ܸO�H-*�A��|CS�G_K�Mi��"��(ܪܭ�u��b6W0���G��)x����JD�éw��c2IW���xc�(F���e3���S^� 7�Ͻш��� �����m����wu	��`��E���t����v5�3�Ss*�|�꯼pb�:X@'?��P�n�O{Z�ʖy�A��0���ޏN��pM�4�o
��;+�j?��2�"�N(;�;s���ME���M�~j�\����"�w������{mnF\�34ʭ��yc��{�A'"����&���K��_ADs�=f����$�p�:W�������p����;�v��Dw�bq�̉3����j�ػ&Sc�yх☥�'	�{:i+��� sU��ОpB�d"���i����20�C"�e���7EI��˅ջV�H.
ST4?h�U&�yT+�B��ּW" �����������c�W&VS�\ԮI0D1��&�0��t-�Q����f���Y3=� �A�@ɧy������]�'Ae\������P3R�@?�X�>�a����%\��������D��q{���[p�#�UIj^��f��h3��=Ƃ?�QE�\�2�s�w�A��"���Q�D�
�o%[�P�L)@<<)4k�`83��Ƅ;�}ţm�n�T7˅�[���ڃ��]�A�VX�������4�H�8YW6;$h'hv�υ�j@.�������RQ�?�G#��z7b�!�}O*�Ԛ�-W���%-P��ƃ��/��2۳O-A��OIg�Ejrr����?��5x�� �"�[�F2��\�،l���_08��tSy��۽-G�i�wqn"�$��s��	g���W��U#w�~�cv��|r(���Rn{���'��l��$Ib�����.�;�%����8\��?��d�0�ģ