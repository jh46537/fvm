��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�����M�+��P4��p�<�� ��L�F9H3�(���>�q=fd@g��������w�u���%/y1]��-�$vC�R$�S�<n4�h�RB��!�u��l;�uXk��#\���{+ !�4��r�����Yj|]�}��qZt/�}9����6�A�5�T߮q�H�7�YK��Y$S��(aZ�O}l�8�z%�&�k��o��sǑ9n��j���=tКU��Ke��{^���>�n;��<��h���+�6)�MT�e��/@u'�������9����1�����Al�!�������<8PΖ��� �)��_['mv�B`~m���~L���""���N�%<6�M�����i�?���Wjk�l�����8O�h�\�q3��%B�	8����T�n�w�`����R�^��]݇sΤ&�*]gv�-��Ȧ̢ԱVN�J0�Wȁ.>��Q`p�#�'��mI9�Z�9_��¡j���͹�$�����2w�J���u�cz
*0�9[�cw�� �̓<\ݚ�'��2���(9����HAmp%���[^	k �ԥmJ�gQ���Z�،.�ã*����P�ڋ<�Ō��?	>���Q�w~>�{��-��n̲X���r՜Ѐ^O��,عLUغ+�+	�d=�Y �`n*b+���M�sԶ�U��t� �H�}IZ�_��x@"��ք[M3� �p�?�s�9Qf�������1	i �n���pXo�2ږ�>�<:q�4^5w�.K9�\�4���P6��TE��y���6�)���ע�z�L����VШ�"G(�C��}���@_�(��6Ҁ�w�=�Q�"4��W�򊔮� w�8���E�R
��F�8{G�P���`xF����i?���8h �R��x�m�ͷ�Î��;zf���C�#�5>`}ȍ|4�tUf��
�~A��<�dG��$x���:R�zU��)p|�2!����Iɧ���kwO:�V�+�&�R��$���2�"sYᾠK^�뇄XN�L<��Qq�yX<��q߲,�Cy�!�q�P�B5�� 6I���݁f�6w�à[&���qS,|�?X����� ��@7OR*���*��\���j��\V�J���H�u０�
�
�v"5�I�G�4����-�	C���qz�?@��"N�Il�ʑ���iH�n>�7�U��ȋh�m�n��g:����2�u�ɐY׃�R=i�Qn���N�MN_&�r|+������=
����e�̐�He���O��'�(�ɤ<���9��m^�A�-�&$4X���u2�)M�f�B�_�p���R�#�j+�=�V]�s�9��\p�Al3=���	��<I��W���e��Zd�r#:����r����9wKڀ�#�n��9�ئz,�G�ƹ��0����*(1l��.v]�#�|��ز���i�hG$�>�*�7�l�c��G#i|B��dhȸ�E���X` 	��N�-��-T�������@�iU�@�5�8~;��Nj����bxb_M�y�B�n��
���C�����.w&CWi�\�Z��{��xF�b�%�O����I��Ҽ�i�A��� ��� ��l!��W��J{	�.�G(E� ��u�#�R�ѢCY��h2�c��mxM$�4�j:���7�/�M�v�*��+�G?�*\�9��%j+1a�X<�8�g���������Pt8��!��,vͯ�C���;�/�nx��c�H��r7<I<M�v>��OE��ދ�b�u.�y�� �ٺ�N�yL��4;���|{�#s���3��^�z���ls�sF;�8~����`��1�B����d7J�[���������&�Cs�O��jw*�
����CX����~"i�dHg@�)r����^m(L��rQr�͆���@�G)��Lhb��[-x:��r��ݫC�B��XU3޹/2$�(݊�����!>��a�T.���jd�?D�#��h=�ݳ�_1�x����uW#�⦟�.C�׆�%B�&���u���3�i#���Y����'�}�y3�_^ �m��VJ���h2�ΐ��U�	��;�����E,|XC�b�Y@?Y~���l��I��=����حG��r/G-;���x���dl�1Yw�������-�oF?�԰���:a�����<��/�N�{��o�Z��4T��S�_�ۈ��jj��ɏ�7��K/�i��" ~�N�f������00f5G{�Jnps�M^�M?0�=�� ����2&,�=
���7�S]����7B��Tv��Q�&~w�.�K�]�7	6^\Q1�b�h�/B���?�i��c���=̋R7c�ں���L�«����/ ����1��e�{k�%��V:k��wۣ� C��G�d0;ͷ
t^p&����Wv�?Z<�(��p�kV��e{�� @��C��u)�3�o�#g��TD'�.J�>2?p� ���[T��+�|>,�S�};nI`�C	16yi2�^��*݅���o��<sc��~u'��G��B�҉���~��E���s����{�B]/JC�$�6�l"�tF��`��^oŜ�5RC!�8{�,,��R��9�n�%&0kN����f��j�(�c.1�+~�:���EB����g��b��s	J�{����/D=l��չ�����m~EM���*s����J��N�c��	��"E`�g�M9}I{MpW@dw��c��.��v�O[b�`
_v�>0�S�|�H���P<q12<���Kg� �q�FL�#2��K�����W�[N�6�*R�ı����<�+�sM�@x�G�C��P��U�XL�~Mޭ����*��*Q�Le;`Ӟ:�r��H{�����F��P��D�ߓ�;^^��A+S�Q�lk誶AK@�����J���,Z�.�2aY��T�ȑߙl3��tO��jɋ�yd����<���dӬ��hн�G�aNP�t��v���3��^��!��pb�	�8JW���-��ʍ/�ne��#�!¼��ecj>P0"M"�K�^�P��+�ƬQY�#
�)zϋ���I�^�:[�Ev� "���M��=E�b�h$cH��纎1�}���!5~d{��<���%jnC��1lr�૽�#�� L��>���Fe� lU���@$�
{h6j�h��uZX�8]���N~���/����V�Z��B��B�NK��rfl�w�%([x��3�?}kvwe�usc��s5�G���A{�	�����&��\C]u��ֺ+g��,���?��2�W�z�B�
`˵��R��u���1�o��wXͪ��X�X���HG����*�E��p� ���m�1C7-�%.W��EQ*j��N�fVw�Oz�I�UH0��u�N���e�C�%��W�`�mR����
�'�ǝ@�r& ����� X�5B� ��Z)�Z���2dnLO���,�,�AV�c��4�/6���?�n�PF�G�J19�r������)���kt��K�Df���*�Ԭ��WR��YJD�(.
���W�s�����\��ES���g�$E�2X�7�6O���z��$���X�M\�J�G	*Ǯ8�ד�ؗ����d���v3aU,�i˶�Z�6ؕWx�`��ԯ�?w�dۑ��)cE��9O`V�/����erR����
�6	͐�_��5�+W�L�u�).�L�S
C=ڡHOƯ*��B��	�Vf���44�(�A�_:�0�:��~]��wq��d�5b�*.�yr��T?�Uʏ�>AW��pfuSc�ㅤO���ˉ�,� �=�^����ڥ��#��V�Xe�aCE��
m=�tm���^�*a��;SD��_�0i�B�=1u�K9��'����zħ�����f���v�o�?D���\�g�*��y	� ��?\�d����*�6��]�s:��?��;���s^���Uo��D�NC�_���&�x�lVB��o��,"��~�&#����jP��ށ|�:KSo�A��ڙ���������u������5a0m� ��z؄��S�p��h����Ұ|:~��g���V=�O��Nb���/��o�\.�uzE�׾��cH[Q�q��6*�"=�q*&��8GL��Z��0!��HK)9C��h���M�=��0�)Z+����v��[\F�Lǰ���Ŋ�2�ڱ6�"L��P��e�=��8��)>��9A���~��`l�ƅ����w���$�\��	��С=&��r6�ad���kt'MYF	�Ȥ�z_�ȅ�󗀮�&�f���,��K|��G�&Ȉ�i��=�'���%0�>�!S�t�E$�,^x��j,�7RJ�7P#)IXH��Ǜ�f�S�?����,S�LG�x��NpTQ�g�|NrI���s$M��E���U�$Ūu��ڌ���5����i��]Xؤ�[|jB�2?�80�΄�$�w,������o6�3��r �Zs�Y��#���݋ʏ�$O''�߷�r��#!k3��c�
h�~��1F���'
�F@~���'�Φ!�3#"�2uE��o��/�&AJfA��m�qb9R�"�r�Z;}Xө�,%��c\�m��1D��y7H+��f;�wk��̟]G+��.�l�b�o!���IE��-���WU\ӀeG�Ӄ�4�����|%��u\���f��ڗ�L���U��g�,��R�ɴ��� ���LqQ�g-;��C���0�c���"�G1K\���V}p��$TŪ�����qr�0��m�A
,+�m25~�䋴����_���Tu�?o�ѭbE�����xU��OR�Y賿eѵf�a]��Z�
@��[��{�#�B�e��K�履��`Q�B��'i�
js�����M���%��/J�6�W@1�[.��l=lB1m��$[I��+�a�T��]�f\�6�?ه��)m_E�M�zU� ����b&4���$����~����߀�׈�Vs�C�5���*3kP�f.�^���GLj+�-�S�7���&噊4[�	!M�9F���ꃧٗ�i+c�����Z�d�[�Q�,N�̩k%'&
Yȓ!Q#f���bu���?�+�[�=�ִ�n :�6�	Ưe�\T���B}~̭ef�Ԝ�S�'��0��0:�cac�w` ���~?��]�O:4����Lf��{Q�ԟ��).Ծ;ؿ؝����c��-����,���inRc�1��#Sg�oߘ,�f�P��l�(�S{O�ܤ�Qsu���2�Mln�Bxԛ�������J��% <q,\���(�*t��DC������O�o�>�	ȔT�}�a���\ҡ�|)�D։FV�:r8U��0~���#X�B�4}�sh\ @�a�	t]Ǟ���TW�yk/ �w�ō��W,����!�̻8��|/�̐%+�)�_܎f����^��4���Xn�S�J��)���fm�Bz��v�m�������k�ܯ��^?Dú^�nz�l��BI���\O��耙������y���̺s}M�:F���� ��Y��YV�]��(���;�S������no� �M�Ҷh#L� g�����Jê��c�kV�	���W;��9G1+�������o,Y�?��`mH��D�53�Zrق1���l>���_T��5VU��w�)Oʝ����;��Jԩ-@a!���c��w<��XY�4JSioA���<���İ�kH�����*���|��?��m���E�=�&i6��������cC81�=�'��X��,)�I���;��� B�q�M���*�#Q��Vߘ�4j_Mmop��r U:�=�<ds%t��5;�����ee�����t�D��f-�㱎�a�YXF�E-č8�4fB����M������A-T�ٵ~�c��G�T
�#�^ �)|��]]�3X��_4�ș���{�����ϝr������I&�S����
�3����^Z�^��D���%��ufȘl-SV�u��=I,m$���c_ՒGXa��`ׄС��u B��z4�d��t�X������d�ý\��oK *�LϫV�˫��=�7Q*�Y IZ?����(��p��o�z��=[O���s��w�g`/�`7=8[Ů��@A��9��%��J�4�R� �\}�s�[y�R;욠oo3�k۩/�pNGM^����	��=@�Y��s��I����=n>��SM�{M�2��?�h?F��M0N�ޭ�"��Ν�7G��2�T�=���٪�1��ɕ ,�N�C!q�{�J��0��&�����cI�PQ䷋=������KX-�J�D�[emC�ձ����'x�����E�ЗGb��`�!��1:����{詁�,Q)kh
)�~��E�F�����0;z��,���4�̈������<�(I4q�����$tot�*|��o�����׫��6��"�p�>�4B���Όe���T��4�O��X4Df`;j�.� ���?K���Y_c���k����D�ލ�EVU�9��������'��]١�9'Q�1���t�c���B�,�IN[J��{T�AFJ���Tdx."K��6W���k����\�2�Yb׾[��1�FM��k��z ���Ӹ���y��IvV=��h���F ��o�i������)��!a?T�]�\!HE�X{������a>l�7��؁���I�Y�NPr �HU�����܋������Л�c��1q����Z������֠Z�������k��#s�?��^�Oba%g 5���.�*)
��ES�}/<��B�Z<����n(��P�2>�p���{n��kO^P]�9Ҏ>ԫU�+aI��!uC])�*�R��љ?3�
��ʇO~�P@O_�,"�7X�Ђ����\�ZHr�')e^�5�?Hd�gI�o��݋-*������f�9����o�Z�m�H��E���q�F�M���A��N����N9	���?4<z�G��3H�3ӛ��$-���O�S8��&Ɠ�>������f3qrI�<�0�8h�J��1d���H��P�:��u^��cW�=�C�����v@jCX\=x��l�`T��HP �T,}w %Q��s���$:*�Ϣ��3�O���*o�a��eF��j\��4�F��ͳNV�%I��Yӭ��DL/VBi�k����9@jq���? �[����s�6Jӗ[[荟�/}�Ik�y^��Ujy���e���|�fp��c1w_cne&�"SB~h
�]en`B0�{��.�󜝫�1I�y�%��~�q�.5p����\p&��7S9�kR�Ɯ�9�Fi�a���Icl�h��#(f�,�%[j��a4�U����Eb�~������ŷ��ȑ
p�& 8̅�3܊�TfE���k��A�>�vC�_Z�Uk���o`>�yô9�H@��y@;�d�*�Q,��T�����Q��5��Ͽ2��;y�/�g)��S�����{0�������ϰ�c�d�]��j���S2���F_J8cO��l �r�i>HJ�` �}�gJ����)�y��Iv�~��;��.���p3��Ʌ�����~����:|P�LJF����3��KG0��>�������=51��x	�P��7^fu��uF�_}���t��y�<_(V����3ɏ�c��06�9�:Ch&�v�r�@��i��1��<<�$�?65���p8A��60@3z�ǈ}}�m�s��_�����H�()��e@�TP�,��d�|�ky43��5�.K������ 3R���g������@���m��SM��JV��Z�y�	�vJ�p������vܐ���1�o�A�LC�W�X�s�}��P��.������+s���Q(=��I"Lj���1oY�nn`��O�m5���py�q�Q@T;����ISKi�Ȳ�Y>���.hzj���B��ǈJp���t�ኬ���$�%t�=����|�]���r'��i:�:��p%��M����~I���ԡ�4F���/��Z^��Z��f��?O%���:�^G"��t�{.3|������yI��g��<�N�nÌ��>#�8ކ]I�M�JKniޜ�-E0L	|�4�w�A;��q[]�T�	�纂����FR��I�G�_;.�j#4�y�0��"!�����W��@{ �����*���*��~ï�P�G�v#�J�ED�l={H@g�_Ւl[��@�鰵,�#�E��E�ɫ]ɔdZ�=4q�%�s�՘C)��(��0@��l��&Jx�ɧ4C�z�.��	�
KQu���/p�j�3P�X����"���М����sd�#�w�3�U����WMW��$�uA~\��������v��B��D���,N��^\Ƥ&�JxL�ﰹ��+���=�/�OX�7֩��_�8J���ln�r���V��r�Ï�fS���l�pr����K�P8���$���-���S��\��J�	k{�	|�SD[��%�A���D�q�e�&[|�A��-��y0�b��v�U��s��z�5[� �V�h��_;�G���	�������P�D�B��b����T�%��N	��J{���[������n���
�G��64����'��XH-PhP �EU�ξ�*j�!�峅�-��Y����̼�SnF�w�!���}Z��`Kf���$ZFJ�����.��N#!V�^A&b�1�N�2XD��������̙ʐ��U(j�a�F-4�!J��B<$~������b���>#>��5�;��i[��5�ۣ,Ҍ��P�S�Kp}؉8��۰�X<Da�?�!�8�ndI�����3��>�����*�Tj���U��*��g�r���rr�K��t�ѫx�0���z��5X�¹d��B���ewY����<
kQ�)�Xy�S�"�|/_K�~��6@��J��Uk��P�\n�0�5]������V�L�|�� vr�����i�Z���o�;=[^}UڗV��ʴζf��i|��)���R�6n����W��k�g�3S�W��욍x����R}87+�D�_���H�;8�����Z\|��@����o��rUxQ@z�8.��ګ�q�(���N�H�6	���ǫ1��M�2��J8h��S�룍�Y@|���PT�ˁ��7����d�@P�����
�h/�$h,"�S���JY��Z�#$�P�NL�
S��y��nB
�E8�X���2\ʈ��Mt|�]�#�f���٫T a�C�?y{�`���KM���xD����	���d�t��55� dۼ�d���f.@w�[�62�Y���'(BmnT`�B��j�(��;��xpyvm���P����y�I��L�%X�0^�������h�uw�����r�+��g)MJ��J+�@L��.���Y�H���9�t�bTIV!�\Y�	���X�_K��9a@�I�fp2mһ���-�>Uȶ��h�ӂ���I׵�K���	�Z���.)���e��#Gw̟����*z�ѡB��W��ǅ�6��8a�Ɯ��O�NRH��
�l����Yx�=k!�s7OV�a�ӯU�"��D���/M~�DȪ�1X� >{��W�K����*���M&}(A�{�
A溔�^5�)G�S�(iP�;��z�������+n�;�q�T�Әf\�FM�z�X��h���D/����@Ԡ��_�3u�������㦾�0����0j]�-U�}t*QhSWeE�Y��3�ք�u�����A)��.h8<���ˑ'ُ�d���G���E��O�=.��JQ��F�W�&�W�7�o�}Wi�N�lB��`��o�ՕD���NC�s��$�-j_���CwA涷+�
��5V�,���jÉs�#A6$>�Hd-�rb}CW\��6�i��q���	�D#^��{��2&�x/��Gv2�݌a�5�((��ի�9ح��L<��+�̬�\3!��C�0t݉o�p�{��ub�͘�y��GvQ]8�kZ몞G.O�� ��¾0հD��M�~F%�jJ�	����-Y�L!!�d�D�����
�H>�y��q
ŀ��"����*V����>1rR��g�aoS-� ��&���V�� $$���n;�Ú��iѱɄ���p7�6��ŋRp�J������Wȧ�'� 9~n1X�2�`��C�QI-�fЕ+�V���W�)s쩗�����
���O��j��:L
qgh�g6�a�iT����y�	�kdnr1���4u�h%�w�\����a�Pg�ś��%���IŔo�%I�y��]���O]��!tj�3[���n3�39�!�K����0����CG�}]P��L����/�3���WĚ���j�d�L��MM�&	��^�����G"5%��O����x��5W��;)�~�3ڪ��J7��H�B��M��?�������?y_��; �aAՅ�j�W��r"��Yx���0��_��Ѕ�� Z��O�gj�[{r�]o?j	��0#Ct�SN��`�[Iݬ����FK�	�������a�¸2�]�N�Y>Z�fa��q�r�/�4p�	�m���
s�`^"�JÍ8T�ie�=�3/=�\W8Kl����	�zρ̈�e6�Ӄ��rG����J���F0$�`29��&�آ��f|cFW�l�o��΅�͠޿b�f�dw�&:36R�#�7p"�ŧ�� ������	
�P��6:~Z���>��>&Xp�����5&qk�+]ꂗ���;9����]3��8
��?w�]�O��f���j��f�>�%�X�@��q��@����m��>�'V������iN(���q���jDeI�y�܇�(��&ڟS�I��Blgz''�܀D*���	��"����)$ȟ���e"��Xh�D�ުXoef�U��[C9���i�1Y����<�)��	ݰnsG���h?�og��+b9+4��	H˜����!��N��7-y�.��҃!=�!��X��_��%��z�@Ci�{��m�h{8�Y�#b�o��70p����{����`�	Oq�� 1Bjio�{*�~m[�p~��[��ռ�'�V8����Y ������`��N-��zK�L��7�'	G~-ȟH<�'4�� ��3�}�Ss�=|.���	���~�w
{��)�O("MTPY	�6�7��o�]�!�]*䋻��7d�����F3�a