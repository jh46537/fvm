��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&Y�%�ddؐ�ပb���p@}y�| ݀'�2��DuE����qs���E�);s2�>t�c��L�/r# �>[qM�
�V�In���$G9_��gb)O��-��1@��I�A�0r_�xCq�\����Z���m�}E[�T�d�LAA+�?����LU�S��#k���_�+����D��/x>�R8z�1���xi�G!D�f�70�|�=��2���ůf�k���on���Ӂõ�2q�d\����q'Mg����'N�ʙ>\	Oy)}��/+�wwU)��<��0Zf�^��:�����"����\�y��힏�x��ܲ�wQ��
M�|����&1�'���u�.f��a��Q�*���H첪�O�xor��ĻhO+��VܛG�:�w6�|��������|<��Lp禚�+�e\�@[������Z�v��yI�m8CР>����|T�w��}lH��!<���]Y����rF����y"n|�;	��9l0���#�t> 	�`�B'��;6�Z�a �~��]}�ȥuJ��/3$m�����sr'/��r{Ō��&,���Y��i������s�J�>����Ʋ�OY�Gó�ͷ �=�W��C/�����ԙQ�:~���:�i��㼛P���H�3�#V�%MVB����Ȝ7��с��@���/�N�9>_#6��HY�uGnE��Nt�����$���Tuh]gϏ�$�3-��,��=oNY�T��`�K@q��%��$G��f��a(M��7[��3B��Epk���R�����")s½_1z�϶��Lt%˾P���2��J�2_B�).V0	�z�:ޔ�_u�N��Ք�����{�;��ȃ�F_���(p�<1(S�S��S�������A���4�#��	�j:���q������mH<���e�bqwa)��s�x%��%w�e���5"���7��(��V>��l��讻��c�&��`7ܝ0ݢFeԱoA`� ���9�2N(��a0��r4�_G��Ѐ�5��;v!��mpS��5��������;�sV�A˗>��'� cD{<�<�4��	"ǐ_v
M�O�.C-銟�`K�����d1�����-����k�Z9��oэ�bv�!�Ս�q�9�3�te��ڿX+{A�|��פ�e��"��[�����N8��&@{S�� �� TPG�M����pR�끇Y8��\ܩ�8��9�1�@����>,�u!���6n,e�)����R�m���R[?z�m��G��%B�%h�u�K�b�ǃ������H��@�|��P�D��6�\�wXzp{gg��ja�TQ��3��L߅�%\'�����l��0�8��jz��sAQ̵��Ip��:��QizXLN�s�g�4���m���>��z�[|=�`/u	X�5�Z��]I�_vH.��F�	��o����d��ãMff�'TNu2��8Qg!B��T��+栳��tg�(����V�����E�m�Prɐ�a�佽�
���n�4n�}#rN�oYrnҢ��$H�Y���"��	���PiX�g����O �>�^ˎ�/��0�J�"�sm�&���i  mNX艙D�@aZ����Ժ�� M.��)���b�H�yOD|G���<	�Mz�0O�Xe�����Z!5�N帬>x���wg����L�L��x���v}a��IŤ֩ͫ4�f�|�r��
�g���6���FW�#߉�F��)�vs