// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:57 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rHed4aJV+n0bjSXlRUxuR4897meCkWvAEsBfHOp7lKP3hZX+GTtvXYV4w7rBhLue
6wPVRHpukVijOBdE/AYs6kg/ou5kqs+aL9YLwy+cv8Na+vA6BVyQejiXg+mFDYIl
Ga3a4SclL9yIdbU6UxCT1VPjU8jxgPj961TkAgMA0iU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7728)
b7Sg71y91pENCqINgu4/rvraCoxDnvMmeEiCDJbiPPGSFjMGW/OvmvwqxOeVxhjv
y4tMRrUlgt5KDuiwsFiluK+hopAwTXnhS7bMIBHx9grvXgqnhDZ2MV2Rse6sPY4R
MDZvEzD6Il8geAcpetwLHMqBUj1euGHzcjASx6sQ/FkCu7EdOmMehxbOqmyg+mFf
thp48/JUMT6jb9MNnhIdToBt/dbnVfYvA5RuYoyKBEMQh575XNqdYNUfwayYTVqg
N7cwwkKwJhXJyROAvuHr4gqm/XsAQno0ziQ2IUKa10AwYHttRbxsjrLb4DvWtZNu
G6tho+QOGNerWGRHW8WF5iEXuGaalZHUsG73Lanydc+6BMuIXlVWPyLjf0XYgOhd
4mc146W7q4xLR0PzD7V94vrAK5ILW/U5DwAMTvX36syzop/qZKGABfO7nwoRMssg
q5S0c7K9pH3PIvxkiQQbUNyYP+yk8lZo3nbYTeTTRHMfkoXnyh1gDTvkwenb+fDr
V/78/JrS3bk6rzj5Lr941xMvy+3GrG1tv+88Re1Rt4+OJPwpxW+iUpiViI0dDw6D
VnT1PJbcaAzD0fyCZ76yDevz6nt8tPD1OmWdrU1emzy9WWbZFBcwQT0p6/6mA2zx
/kSzSX+HIIZjWfHEEYcjfL43daAYjbszznrvhsXxfBVrmUyvP2z2VWsWdV9z7wFE
e36uuTVqNvAHc3aXi9uNvAA8GBPZvY3kYcJvKF++YoTGDnZFm9S7X3uMtdiWJT3A
6p5jIwJ/3eysMf04/MsakY1Xu21lnjM3Ncgo8trKY0vdAYT6LOi7sMkbMGDRu1zb
L9W/ne9HanpGlf4byRNNKOyJd5plZ/CcYq6MCIOOs6AFgty5/i37WaKaPwoUiqe3
uQl01oue+mxK5jhnYd0e/ws7sHHQplTT0dw0XIaU6D+u05hSbEK4XXESmfssbAEb
tWLFDbAW6qvM8/X78JV87L+aqTYi0ydLfMZXKVh9TT23BDiBI4LsCNDNquRs5YLp
GKwddXlw/pJiS6ukaCRl64W7ML1wpB78ZAu6ojixD4JqVCyZf0u6CpZlPDtitw/y
uPmpR2dSLx5cVKuBo4ihmpQJW1xvTrThkTa79xLtkoJ/nPHtj2hKx3OLnBpCLh7k
vE02N0v9FZyCL3UOu98rp5BNu9H8h0XfMJijO5TUJNfTsOd+L5aEvvLNhh+5qw1F
64bQWzIqZ4e2xzIYc0jk0/vxNTyYP51sS2kYQzzxNoCCuBqqlFbkRrA7KssvZqfS
JiiI8wUEnUes6nKwE68c12CnYS3kIWiYe6qh8uf25f2olQpuIFd3159PiRKvJf6G
Xk9HmqGKsgrqEMQqxx0898BaM60NfLSu0hB7d0lvnEIVoG6IMrTBkBhuwwzxqZa6
x43pW6Ol9c8VBW25f60mJGpdSUYtyVTT8/vBdtz1uxscnImmDyakXExqbLcGsNU5
2w321LfFIE1lE4gAoGsaXUgem3J7w8xRO3gB9olwvvfDETajomxsgn1ighzJBrQ8
KgxOrBG6aiWt8ymUtq5QA2Wq5bjuiITUKaH8ApJIxYMhPr/15JPOLPDUB6OYQe3/
2n1dJ+9QyOXhTwQCMKJJXywhUdTHVD+EimjnauWmLnadmv2mCH523xmsfdJHbSfr
BvV4vsMZY/pOFl9jpBCh8qGUuqk5w7zQ2qBTCX2JtYI9MXjw0C8rAWglU2qWxe5h
2GhGBl86DJrHtqw9gDHyXxpfvMY8j4BsDRcUuh/jc658L1MvcPqRK+9cGtfXgByY
DN0nX+Qx3Av/x3hqOhG8lJD5/ZqvaQImwPsJT84zVucLhWpah8N3azHfiY4OFVSa
t/6ln4A6qTo++wljgyrKlQ/SLCPz/R/wBHGo0r5FrfiMPS4j6/asQczXssYwtTK3
v2fRAegvj7qgGITvaneSbSkKA+I++SUzPsrPBTFYIy5OCXSotknjTxCjsg8EvcqV
ZbjfKUXwpx6o+NBkzry5PnlLicFrL50UbkNKgbUIo+zQESiZ3cD0HTco0yEV6UTM
8d1k/OkJoDv+F9uXBcBSA2wCXDkw+470JIT49+aW4NhZ3ZsX1xcDpXvYEUn58JFa
oq8d3vP2urSA2cUrOBKHnpr0LQYTJqJA+tV/K7wqWut6EpZj6iM0EtFkXQZBE49U
pIaGNpqEfu2zcQHokDemrr5L7uRBCNXaqkClnc4IYmOQ++d/CHe5DHZvD3oFfXEv
fWIUbULTq/NKNHctHdtR4XIWVxQ2Gqrkqru0/CQNswdw0pk7fktNevIGIEjSJQKm
gf87X9799Q5h6nBw5jovq/pIGW8fEC/r+PVvIUFzlzNtX31CS4Ohbt8uiYyM5cbs
4QYIPzDQ3lnmTZGrl2NrR7+6hliANqsAhgfP8ja4s39jGLAX14RGbMQqfCeSmTOQ
9vJRZBACPaguCKFVGuSBtb02JvSVQog1h2ygh9in30CplndA9gZYIZp4q/YQaXmK
UrfOR+/aZ3UD1gjGF9an2QvA9qcEp+HFegwH3ffy/DzX8OYhhL/GVhn/562BKL3V
780oWRci+MvpBDzNQ0MqVFzrVrjbsdkg06msHBQ9abMFMZ2oiHKefNguEDfY265q
+nOTPkTY5gkEdDXRHTVK+IZDINFZOopSbCc2PMVMbCBSrTOBlzflZOVOW1JCoCa+
bUOkKl7ofoiG7jSLpkkctfssasDoNd63SCRGxXkwT2IxKUc7TQg0FJId2JkMckWN
wQi/weWCgUd7KKcAwL0PJ0c4iwK2CPA+te4Dvl4zdoc394uCaHcgs9R32er+u3gs
tzbausHNp5RsRKdJpzIrJEHgGOEWekW9zj4SweF4YYL085G7G5XhZ6Ulp8eA1wNY
1nxyHUtD1FKzdlbPUzxuQNOSy5lMIERLANnZT2UwXRE+jt6OpKWVFV7OKSIO4j9b
ToeBAsTgTtx1AZ64H3rFiblf0xPwpL8/hOj2auuBXnMVA1Fp5WYaKOA8zLtz2rPm
8t+CKEvs2j2StdqQlXce+cIzEr0XxVnIgRkPEphrzmIUk+G0hSwIduBobeo/pAZj
KsBcAXVOAoGzL6z21L/kFhNA0OtIqksinApc2+HuL4xrqQjpbEOoihr2PEPaVBHD
eAc+lNaYXEtcWhGZ72vLACIUuLzo+ErazMDOMBQS0eB+FK9gKL6ylrRHx+sSlYCm
KqpEnaGtrxDcdNz8/2YU2JAlxB7hEoL45OUgCLuCN3bVWSv+RX9O/mUHhj9nCh8/
cRTJpIHbx35UmzNvu1+MGvmOownbCkxTJyUOLkQvIGFLB/SARlul3+cFzQ9Bgqm2
pflibH2jrsSlPpPB/PweSmgkg0ahFX9c3J7IDe1yNv7kSPPshmJjqLV4CNzfM240
cALF+E0vYZXT/DfZ3C6+QgwIATXd6SLpZ0QP1QXfYA2XMdy5RPbyrW+7z/G/X86A
AHiyDFuCOI/p4T+8KRndc39W8vhFjqJQINl1b5/Mvmz7NSRSEyjqU4E+/G4aJBhr
xXRNk01I9KBhxPWNglT8lm7VJs3jWKcIIE6/hpBlXzgNBnLmx3P4B2sKfhqlehRG
gQuRTK3iWegfs9NqR8HdQ3zl+MSLlEHfha9oXeMzsFpXtsDSqe/weOcgeSDqrxtB
UfUPBUsSNcQnsc5tCLIuL4f/zsx5m3GIROMG3AmZBc4m/aS+xCwC1UT/ZfRR6UsZ
QBUt794ybeBQuc8pexryryTs/1Y8K2yo1dsV0PIJK1O2XbGdhIHcTGj4mmBXlO+y
cM1+ypdGL4ULem7Z7CQgdvu2HvvAglNfk8wBW7PQ/97pYXkFen0Zzw79i8TaYH7J
eZhkxDqG0YXL72QPbVDF8qpILEXSkOhbFECv/hp7yBjtkaDv+y2LyvQ0jo/Re77e
TTltHYKRLEpXEPjoJkBMFsnnDeaF0KM86LeYbKIRv4sTl6v3DJJQI0JXL5XV5Kd+
GGqzXAJYCXT9kROtaDLIBJkypGBLHLMkbmTDJNlRMYKi+PU1YS9SiOkky86j5neV
Kyc+WY31hvTAD2YSew+CjVHjsZ/81CUMOENuwuVlMTEhcVidXgFWFYoPsIk1CjBW
qCK5HlyEOUAzqIiaOShKPKoAGxGTtvUiyCMUbqlyWXmFVN5Mr3J/rQ8sykAim0oR
B0UC7TSljkC+ao5t+3roNoZUuhyqEVH3Q5U3NjkMIAT3u+HnTFX1bZRTZcFFSn1w
9fv5J3ZNxJX/se/VRcUhcgnB+wLaVHINh+xaYrqjOxIbS1Qd8hmGjfe5tgCwlHs1
3umFwgHg45BxeY1VLFGeN5c+KFXC6nQ7hQ1x2jx16OFVMv7NZjqYKAqVNQtn+gZX
x9gHgpxX/2FpLH61iGbZyuFwhuLKApY9UIYfUYUP4OAKby2xdk7FHrRQx/DvYlYg
192hGst6cJUvt2GcmJVf4XyNPJliYb6PL+tiA/oNeaJwMTYH/q0tPmiOw+/ylBIR
egcy+LZrXbpTtkPMKr+gpbXlvYfpXjAITxUN222NwqeSp6TGdlQKj8SltAtoo2ZO
cSS28JNFAHtDwXmrilwnhF3mgnGRGojMyiYg6ifmUIR72B5+A8pOQXEoWNEowi2Z
wMqbvUAX87FLg/K+7s0DADo/RyiNULN1xVolzyBcwT1ooLKo2TcF+IuVrWxXZiwN
9SRwYfhm6JxuAYNDZM4b0ZCawLLu8f+D21l6CD37L53YpCz907ZjmCxk8iDHX4fB
sN4w+QM5gfFnkmBjkB9uuklPjknHRJSF7Zw7SQAfM4Qrwslw8PDd/nxV1Ms2BtEB
t/7UW5tmZ/jvU49QaYaD/hiE8LeuHs7rpM4hbWW1CYisaiQJRAmwcU/UZkVYpZk5
EV+Ca8s7KNmfPpEQXa81Eoh1PkX4FabV7Fn0ikNtxz5v+yfmw+DQYWLpDMsZuuKg
HfgDvpckiZAOQQObwwpdOTuFJzKFf0HtQgWqSkqhY0C6hT4xtxIViQFDjBd9XXdL
ToZMXEgXOhAVLoCkRqQVIM8RYyp53WCvHP0DLnWwspFCVOnSTM0CDiz8+lMo13ha
wtxza28489U6eBlXNzdZBaKftQlfcPVzvXb5uUjqRgeWRgsuOIXVvxXXMUj7m+ZO
HGGMeZgM8WyQcG68qozru0K8+92+TQqvC+ayp7TOmFXgYdG6hF0Tc5fODMXIglBb
7K3Nq8jJpM1P7nTrwLyNpKou0TrclnFMFHAuUU+w6XC2FD0S69UG9e1dvh9+3L2X
tJj7rEDgKGlj8XJqE6IV2oBpgiJD6oD5WIYQEpzk4ZQ1vgtdpRjnur0v19C5Sd34
s5KQ9JdptizcyQbIz0pxJ+7kMhtxY8mjfu2qUMODHX+HhXJq/sdjWOfo5vB2FKvJ
m1eluMCgZMaOpEkrv7Vbq5Ua29br6OHVUMSrGvpG61WEmqVxRRqfJzF3nR6Y5smy
DDXFdi0fSx2FKN1CER6J+BO48hAtYYrWww0o/AY4H4rgY/i0A1sqCYs/TMgY6ubi
owZXXR9o2KmxDy+3a+4DPw8g1xIF/5a0MZI1aQCLGC8/eGcJFll2JyL7WGDK4YIA
acPQMd8lJZtGw1ciTWKmeG9R7A5lfOE2G6tMpXt52VDtEXxqtfp9g7mwy+2GRfG9
gh1Qc+X1/P+veHYNYySAd3Ewa//uinYYZCRWIzGEweRV8dZxguQjW0xEz1IupkNo
DTdm/yCv/3iM/vFmNTYqCN/3IIMAjnzGKSFBYRUvlz95H+kdsXF7TaAd/izL587I
JbNpqULMXiihC2OrWjkmfLHEUgXUloX3lSjCMwlgcyrHDetEsoUC2OktkJk2f04H
zGKt2weiozBv9oNLxAjdLHo+C1RuAtHtjYNzTu2cJzCQtKOtBgSoYYPT1EHI0p81
MAzBOOUeHPHO4hdbUe7xKdXSI0JimZuAPGJQY32r5Frh+FWbJHO/D9TadyQYKFZ0
J+2e/FwtuKbXFH/vk6mNT52j3RFfvq5dhLPa74JaDE1W0lwoRAvxkN37EsUAi+m7
nCbxr6skJ7aNVK8XYa6s5TVtjmG2YAapfS8RcWwFgcOfYNAJ0UTvKxa3TwUPmkeD
eIJIfokNDC/wn7ji3ou/rzDDk0YX9yrARTMWmg5sJ3nK1I6U3OYFieS84ITSABuv
vjE8iU87j1q7ZEAXmRWvcZtFitRfW5QHi1JxQtpqmf/DvaChORbsUCZvTwfHYFNe
6I7MxjGaicMJLX+92BCHoUpshBZ3TEzWg81VF1Tq0gijn3eQ2zOwwnP1eEepQn18
kahpjBv/IQ/JfrlpFSxNYQyeliQgNym3ONUxcBy9XnjpuwxLCkHUQ+2WG2byMSiO
m/F3BQTGvkVWo0TgGRg0E9m9QSIbdFKcjrh60UUvxX+TkQf9KkPEp93MY9K8CUv4
bTewwC6KDrMvHVcX5+Vd6HCZXjjAWylLwAoNv2mtlCw5kT59MkYPJn/A20tdOivU
/reNGb9EyvuBJYGhWeIOi2o6WzpuLe5/fLlV+PCqPYvMsG3Ov7F2xU8rDjCsI31c
MomvtjykIhjpoXRYHzpW7p7zr0Hsr7/ThpUQtIFByAKOrpkXTtGNylf46kPflXTa
RB1Yyx9ZWN4NULgc/jtaAoHZ2+SbWLxvRQQwKdBRVOV3cNBtMJGnvn2kS55pxpS2
vLspKg0Ye+rROjRFA/TfteoYTQmI12dOVTk+RPYm7iyReYtvIvU7OHdRMicICB7f
KaNWDHL3qvQ8sj/MHJF02sAgBlPm2M9+hZyAH102fkXolkERfjr187g/OwXrK5Jj
x0QAzSfb5YZSUPUVb3HgrIBpZeTPaF2XmbAQQ1RRLzM8ID9EXS8yMWuGel86OcU/
81Cm6ZcpOz1qzyJtjbw3+otBdIR7MIspa5MakPD7f73sWwmHzGI/41qxSrv7r3YR
ryXJn6jE+tZjEEV807X6ng2z87LOeqJllrw4J1t5Be6BMwfHW99HOv/LOJyBu1U3
WX9Tsg3Y6s1EP6pkJjDRfNj6rAHDuvXErSOg+Agn3GmQGUTcrZbudSAcbJqKq4xG
zuZ3AOz/iuKPTx3apLWDjyBXQdwiksSFBAFMrSKn7Kc70MT502IZk7P0q8h+Sa9Z
KEQxrCoWvE2wNvf1z5zNuxbWy3vMjKl8wwPtvGLTeox8H56+N8q8mVlN8ejqrZ+W
7ty1KQB5aEXR6rERus9arMbN6am2AL7Y+bflhW7oOc2uUvNLAGUAWdVnisHlTRnR
J+LDJpdyk0nzik3evAclDy52ixPUSXT94AW5OQTH80RCtMec3N8NBOq91R8yR9qm
7m9MiNoAFXVqCLoB3GtIKmoLqgBIj8KUkGbktDFKEcJhVE7RstexBFr7g+1LukPb
VOnDtOuJH0aTZKYM6e1NzJPAWQuFSLV7k5acr/zupVtEVgB++5uO4e2D7mtu+Iiu
h0TVtTWt+l+1stNDgkkjbbmGTjNe6moPe+0WJXjmokmUwFHewAty7fMFJBDE+5Fz
hKsGA+6JQkWTKqtrJqCfbbbMZcm63cEAgzKWmZURWfaItAuUVYdOQS3sGsC5LO3n
zwJlxoS/iawdVqjokhwKWl5hygER1zkOYegcKdjGw/0shC//CUoywNI92W4dzK2B
slb1B/yYVGDa+OlIlpIgfc2BJNuT/5UW8J8IbcOA6V8tkwFIZmGSP3Ba/2i0JfcT
/58QkPLLD5BeIPlKp2G9az2hcu5WdZmpHGgQcU4R7yU4lHZFH1pFVoOrkrRcctmS
Ok+V72Qv9gAG7WW5jPWIgZuzMrvpRslOYfiX64Z1bkg0/wPNlOYAmYLv4wrJinbC
3k2gwNPVhJKrILgK0BaucuuaqBMi9emWa8ahL9Xa84T1GK11NScvfNBiqM/uqz3f
I3lmZ/cZH48OHXidpowW0pZl3EyQ236NetNIHYmjF117WJV0mLnmpY2Y5JGG+GxH
id3Irg1hlWSZ1nF3ktvliQmILSZ8iIJ9ZwYn89KdT6EBjZ/zYztQ4m60t6VA8y7X
HgBUIMmW/83iQHcrMp6Nq14HfENAncnLUHN/CPSGe+/woPO+hpD7qbQz7hml8p+8
ZXavX/IiIpFUfdjvP5eZGx5rDIhY8p9Fvn/eGPZ2TfKO4haoUcTSuz4rLDtR2AWk
fPwQyeRtMe7CT8Y4LJyTsZ3ILcjg+9IgmcMPmi/JLON1Uotzb/DP2CryG7WD2N0J
z7yKTc4VqjN4uWaZd/YS6xt32IY8qUpT7qRZpS9Ct6PjHOLPwaAATQnD/OA7UXmw
mea/h+LoV+Fhk+NKDCPMATmo/yEL1KbSxoSFZyal5tlj66EjU96AwFmHEt9o6t6t
BqMfdE38MBviOJNHB7vwTQp0a5vBXaELhsOknOvc7RZkikxicq0tZNNQtKIo5s6i
Iyfob8pNuZ/kfKk40H95ZK5ihID38h313i263TVHW/Kb2FxYuVUbUQdhVi73iR50
O9kDIjJXny3+IwE59ST/DYqr+/x9QTG6D1QM7qKGLNEtteAmuXqLcun+mfBINObt
0IDXIor5aPWJvMLdihidA75boURcIlJWnpVkWDVmcPhSc9Ej18F2P5lBkrge8Zvi
KSULPiSPU9hWg/Jjf2ec76YL/R6XyeMJTJuZ40DEPgJtxRkg9Ti2j49XXWHP+yWE
nkAUZjiuzRF1Nh5+F56ivD0XgatPiW+1XuOF0webQbnb4qkWOj5xCF/OHnQc1U6z
YSeMb88Ev7mGXqTZnaioowj0X5lL2+fKb1IOU4v6mc/eLwxWmlxqgEmNE524lxTh
CFLYKhMEHNqX840rwHb7ZkhG09IWtU2/Ddzf0mLRSBdfstV8ako1Fg33wT45+YCC
gMFC4g7sMiO6HFlNAEDRhY28x/m9Ph9OVafk06Le5LK5E6+iMLhyB4fsGsAHheYS
8s6lpPhCs3ToPu0XDaVOS0dx+zXcXhhx6SkbMjhKVhkzxy9Vmt+zgTfLm5dF1LZ1
QjoKRvYZI8OFnzzoM4ezQue6ZAA0i/OLZ3Op6Y3oXM0Z4LNoJ2SoUmNIbDkjKmMB
qWm8KVumj+CG5fbrKeVezJSxfb9Omb9f7GyGJjqq4WIjIxeakTPZXCdphWd/dhET
ZPPLh5c3wB+dYii9PtM3L6vpU1Y5Qrp35RAOhifR7sRW9hQwBQYfF7rsIXaBtIXY
UbEcQeGI2Fr8QTT5M/WmLKMcpEDSCTkjPtnvl3VuIgzPZMGzTnwmXyKsGnfGQYGJ
pmygwZDJFS7cbi2LuS4vFdrQXVgd8LZLFIsPY/3AzEWo2Jf5DuvSjSBteBE56vxh
Z0mPkrgw4CW84dCIzUihtO0vsQkyzUXMuUEoK4YNqoHhZhUHLurtHp45faCk1plI
mOULYcrDOqGHwd0OwDxcBxeAp408uU4GdqOuOg4T5BFh4JUZOjlT1jN91mfyb87v
6e58uS8rpuLQZDu9E6ZCkm8l1+oMUGID72x830SagUtevFmhfNczbghfahr78OjS
iLwx3xIgRfEez7b2PrSFwFPUSshVzrMR0EKWXQ6FsfjG+QORAHs1ODasTePdMlYy
ugGCcYWrEvYg1t41mU1olnmuwHzq7OT4E3/WKrUTjNcuuz/H0VtlmZNB/9UtYZWe
G8/U68BznXcS5IPkoNVJu8J0b68mJyVhclaIPa+h2xh9geHo/DG3RQ5Eazk8rq8J
hIChn+fLaUOvxLlddxFxNEVhRJAvmBNtH2Qrn05mZA6YYMjYwbvZq1H7Xb2hWv5z
ZmXnU7Njg+GdeuLJik/kYmwCpv4xBnXDd394LcJEEaYwc79vEkgl1VxTeHDESJ2/
7gC6ZtJ5wSaoeI5HZv10C5HZeLvsgj+q0h1WOBO8aJlhZVLH3LCB0y7XmuuNmzlf
gQPSiBRU81sh5nNWmr42tFPRMetaoSQB0NqjjvDr6N6aKhhHumRq/bboPoGeAw2R
EaLGgXcrr94dQeVhdzjnc0rO+ir7em/HMFE9xziVZUYgKeJFc19v8SXYIySN61X7
VE3XOIRyQ9Y3frkOJ25Hee1A5gUlMQKKGjhrUJRaUTUVW39yrmsoIGoc7s3i5mfO
uY7ZNtMcC40Xewcze/3qNsQctotUHKPHPckaQDhl+HDFyDooDiduvIpQJan9n6MZ
5aNDzNZRm/hQb2qLDVmNh4Z2NFYQkWuDIaZ/6LRKCaMYja89Ikr83BdHlnu9EsFl
whlXj0DyekIldNRVrbN8OtEj1LXzhpjOFhbUi2XnmUwlTSXQ00piug+f71G/VvJ4
9bJRV0k4Etgc+JWJrSgvTXatqXJgT+jadMJgYxwAPoGY/ePXgtccuhEQ0Gli+ond
`pragma protect end_protected
