��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���^�T-��!#��S��v�Y�����I��v�����l۝$���a6�J�?��+��PU�j{�k�QL�7�v��SùJd}[�B����"-�i���?�6��ڬ�4�c�R�!�_��Q�,<�H8��<����7�q�I���~y@c&�9
x�]n��8i��V�݅��E�i+�N�ˣ�,x����(��2,£��~_�lf�U	4��f��!�%��5�Z��H�����%�?�n����&D��j�ӕ�4��3a$Z���툆��~?��=�	b�6r���/Ө�=^��I6-#N�D�I���Bo-��d@� a��4W������<���e �ޙ0U�Fe���+��-)^*���.qH5�>Z��_�4'%�xM�;w��T�Z�it(�ڊվ�C\u��om?�Li�)�q�+*w\�u59�^���zrQ�����Z��rS��m�Adp�ZF�� ���ɹ_���r��Y��/�0R�&�ՉgF8�F�f���zQ���0���r!���u�-s5j�+����?ߊK�aʈ.v&ń���y�6D������}�K�޾)X)P�#�	9~�� ����j�Zw��r��K�Z�VLQ�$ɕzU�p*�">����i,��<6Q���7��.)��WNG�� �KV�5m5���@ Ѩ���"/~ȏWj�����Z�G�s�p�N���хV���`��mBz�^LDҞ�H�.|��`�g ��	Nލ�(ð)ߏ6�
h9�5B�]����c_dC����_b:��k���CB�ws�j5�&�t<��q	���Fb�7ƨ~�a˱���#<~�C���7�G<���Z/$ݽ����������n�ZX뗅�˦Ku��^_p.�D��[)�����e�N�I�α�<K�p�#{P�<�5NӚ|�i��6��(��0!hR���P6I�X�Z(u��Z�ubg�vX�<����-���
�D��]��F)ls���d �%\dB1�tv�����ݽ��Tьĥ�����\����^%&��ư���D���(�6V�h�x��>n�0����廪�$�E���>!a���R��C�yR����ܪ#Ԟ/���3߂��w��H�"x�)��xF��;�^�b��{�s��ҽE9�ew/��[��l��|^�f��cl���0QuO�\!�[�Č0ۄ����	$
8�e���u�~����?s�$�[�(,n�%:��Ut���$:;��Kҝ��?���.���i)�I�

�tx�c��M� p�o�ڒiƨ�Գ8+$�:Kt�a�<�)��8X: �wji(��[<���L��Z��f�0�5�%�'�8�CGb���qb~v�WW#Yk���=kWx�*� ���}�nr-�h���w�٩��թ�Y.���0/��h��T0���K�4h�����1
v?�o��{
s�`�{yk;}%��::��s0/�:rS�" �}�#W��G�WA��B�6,��h��F^�E-?9x :&�]�C7�i��F������cEJ�{P� ����h�Kw������������@���溭�~O_f�{�{ɰ��g*?�""v�rACk�K:q��;Ӻ���Y��C�׵Xs�Z� ���MI9�=���!9 }�M�
s�l�$���B}B�rB?*�"sK=Jl���\���,A��R"À���k��2#E�f����%��fR`�H�[��F��#��%���}�
%H�J�ñ��h�<c��2���K�[�$�`R)�l���{]��vb�n��=ښ'S��L��X�3Gc�#���m���Ş��`9�����P���"/;�<<��e�XL���M�D- m�)ոx_��Vߧc�����~O�5T�1<ݩ4fN|yWl��"��D%t�.=9/��!H�)B���FPtTW�]������O0���Eo�Jհ��,��<k^&gF�)6b�\b������������M�x�U,:>�eqmƉ���=B�e��#n�C V!P�e K���0<��?u�\;���g8l���1��ŵ����,�U�+�/_z��x���=>4������5��W$�j���Ď�AF��-��HW��"sWCQ�9��CjI�M���B9�fq�xϷ����:vj��Rh�D E���S7����U%)V����~�ی(Ca̢�ї1�"r��VB��&�F���@��u) C�x>;a��Ay�G�y����q�S��lI+5�-o��ŝC�� ��W�� %�K��Ѳ��u�l=��C����lG|�4%��ak&/FCI�6-��ʥ�M�;���{�Y �c��6��w��}w�?�� h2	�XCy�~w������>ܮ�л�l�M��3��g2;ī�6�&�<x�<� �gjע%Q:�@��@����C�V�Pl����BN��$��d�K�M�ʜC(r���h��_$���0DHpʞ �u[�	�;Y��]����[�$�y����t�:^&��j����*����.�����\����v��é_[�SE�}���/�ۅ�4�4�+�"�� ���w���~Ҭ7S�Q��I�rQk&�ʣJ�ztYTVv�Y�`A�����!�l�����%B��WɵP�$;W�.0Ƣ�aa������#��P�O��TM ���H��Z�C^@\��[�Ur/ގ��5�Bv���^|��̴6D�O~pNm����8�H��z���I�G)�~rhg���N,������A��L+9\d��ʄ ���ӌ	�p���aW��	�i�+�#ΰ��8�[���>!ۢٷmU@����q�
��B<M�l��C%���(�l2eW�||�'���v�cn�:4eLa�9]w��S�ו>��5�O�D	�<��Crk=�;��ڼ�� �¤�4��X%�$}��,%�G@��Y,�R�C���S�46nXW �X��&�F����;�j>DW92�C�~���]�r^���O�<�>"��k��9���5��Y��T�t�����P�)WX3��.	y��\@��&t��`��x ��)�G�i������1�������)���$ B-��=��㚁�oV>R`�U����-�MQ@��/80?�X�ʲܤ��[w+�in�>�^��F����3��"�N����NA�MUv����~47�=@��Hi�x�5�$�m�owo�bt���]3�$~��� ��oi���S[�]�^`�]���$��;ܝ]��-زlpJ1'>��ԟo�BH(>��`���$�v�Z8����>���&�s�F)��΅�4�H����瑉>�؝��I�0��&q�H5����"lؐ����v�GKezP��閔�ú�����Z���	�X�[�O=|�x���렗yW�Sf)��T���^d		.C�LK���2w�40���
�)��it-��ͼM�e(����
���.p�B�1���m��(�ɑ�M�c`���={N���.jӵy��vD�ec�$mu6e˫lɝ*�/+i�kZ���T`}�)��.Bz�����2r	Ϳ���F�1��L�r\Π�L!���,|����S_���d��q�a͒��Osa�W�`F�o@	i���q:��UI�c��'�a+�?T���o�z��g�@M�������6�ζ�١"q�Go�V�$�߅ytE������M���f<�?E`����S����nY��')��S!8��KhEg�f�F>)���!�m>�q��R���;��*��	/��G�2�!}o{@�@��Wn|s봶�4Mb�0"g�J�J	��������hx��{t�sk���A�=���U�F�",䤅�ʤ����X^�������~MD�b���*<����)�N��d�X��;#�֢tRpT(��P�����$MΆ�T]�_Q��r�Gv�+��^�>�����.�s{�|�B��;�|��65u$�i$�%F�w������
�[ٖ����PZGz����o�릒���KF>�〱4�j�ܼ��!�������Fb%�ӆN��3|g6�~?��#��[�����f��8�?���J�>
����:�f&�C�:(0��Bp��[�Y�'.��;КA�G���|�x��ѫ���#�t�|���xL��c���ڕ����I����a���kъ�-�&f���B�^�����#��+t@ų�*���a�i�*���TFzє�����I���zI����޸j6��u�H(�&�-H���YR&.Y�`������
h������O,�T�v�2�{Hĝx�b��R�/o`iX�4�b�j�����]�+=ڍ�ғ�������O�FŬ{&#��L��'�p �rA�S]���w����5YR��\���=M�D㮘I��(���.��.˔�H�F-d���=o݇+PAr�],R8�^Wpf7�����@��|+!i=&��$k��G�jp8����W�a�¹��w_8���FS'���RVJ�}�4����K2�e�`s�d�/�ӹ����*I>bز�}����CdUx��3U�G�^@�c��$��<�I6K��N�b���|�H~\G���g�)��ɓD5.�s��a�o��`�2��FX���SVn����i�a|~�T�#T��e���p��8�2�����Pm���҇�?���4P����nӝ����laJ�[I�n 0]J�-�����rd\���-��߽܂屏�9ꣅ�'3�j�&����mv0�*K��y���V^ ���a�\��B���+Jm�p��aI�q�)��'�|��{Lo7�*E���i�]Pca���
�g�ǝ����GP2��0��s[��%����01�Io8F�@�"44�˷9�#�,K�������ߡ3�paj`A}���{��"�9��yL6�=w��zAD>1�y�׃�ǐ�}HD}��_�����{�6U�|�H���M1�5F	}� ���K��* Ց+^��[7��9|eGl|�3�T��r�Wɉ���sE_f��A�C 쐨�#-�B���[���j�L��r��x"��jK�4�_}wqc\Ɵ�X���Wޏ-���;��:���캴�UyoˑGM�F�1���l��cL��@��o�{���ݪ�:�؈��0��(b�ũX��=8��1z(	ћ���U����\	���5��z����Ԉ��6 ��Wv�"Df���J��E%�=�6�^�`"L.�g�g�b���`L˅�޻�o���Ō�\I�5ʵ?su�
�(��t��O�A�˱����Ӹqm���j��F"��ș�kѵ�U���X,������#�YC�*_���T^kG��$ϴ�xM����E{ūV��_ܟ�FЧ�h�K5����Nl>P�@mϐ}if��:�v�X������X�wQea#����UP�_��$�@����)��c� �9S�HxX!o��lH&b���CY<Za`�=5o&����_��+F�.F��R���t�����e(�?�~Xh����
��gzHB�")�J�a��uM�0�i��f�1C�k�E
W ��57�����"?���Ou�d��ɤfR
6OVh�O��#�ɂ�M�*`��XqEr[b�Y���i�F[!RNUg��+&���0�_0E����&w�B�%���X�~��j��dw�$q��#ϊ��ʩ�s��a9Ӭ��iB��ֳ�g*a���v��_�,g;ƵV���;�ˆ�]��-�-����v�����u�p��s��!��UU�C �pv�k?�/q��ƛu���t�'���L��g]_ظ����a������|˿�a���.�Op���F#բK[��S �cC�[@�r�\�*��'�1)ga��9Ԯ��x;/�A���V%O,����.W���/b���m��M7%ǜW狞��P�3��K��O0�&x�o�������g=.ǒ��;3q.�q-�T�Q۾��P{k��}��vH�\�hO�ѥͩ�� �,��e���8g�g��%>v��S$���X�l�c�����\PӍ��㩕ۏ(��e��Z���m��R"�.��:�a���#&��%��CC�ԣ�4�#%��Xx"sO���Qk��njQsy�	!SG��{�k���Kck�h�ޱ�;Q������a7�mw_����'�t��Ƥ���
��K��"��o�B=x��M`��9�G�K4-V��a��ŏ�(��wj��Kz� �w}��`b�4(@z�Z#rr��	 ����{2�>�����U�[�)EY�_�s���>J�˧�'f������]�y��v�tځa�����Uk�C�R
za𯾟h^�n�L}`�>D�I�]5|!U�U	�}�Կ�|(��m��K�������<\�6:$�(�nSf�H&��w=�7��?��xr�~t4�y?����9<|N4E.�1ѻeN� ꟩)��0Ʊ�ӳ��Rn�ofOcJR�4M�c�"���3��s3����:���Gwr��@/-�Y�� U������[i�O�ݪ��_Y��8��|m.���e�D�Z=�P�Vk��t�k�^(ښb�r�б�U��k���I��n�eoc1)�x�]1��G��~�݉�������V�
4���
���bZ��\�_��.�t��)�우�j--�AJ���턦�i7U�&1�o�x���,�/�z��ͺ`�,��R�2/*�0�Q�u�VF቞�UG�d��LP%u���'WUY��788X6���Ԯ��r�v:?����Y���O��*b[f޻n�E cB�H��������� �;��|�
��u����i��w����kUQ��t�i�	1x� �Q�}���r����������Nٌ���9�]����U�N���̫[�'�/(�{���Zntg���_���引Q��+�d�I+�Ѓ�h�7�S�Dg�t��^'I��okZ�X�;�::-h��i�Y2J;���B��SQ���U5Q,
���u��y�p�m�$��RB��Nh<��J:�M��]�Р���_P��9(��e�= ��5��&F�'�ב��C�t�z]��4`ʈ������ٰ�4�A_�,Ux'���]�2��j6�#M�u��i���gi*��΄�O��إ��!sU��S�d�޼{6�����m��ȞwT����ڻ �R]�s�����@'����R�1�S�G��%�<��� �OgD1p�.df��	�C_-�]�i�w;��G�� ��|1�=�$�E���~���,�Lqr�D;�mV$���vC]i�2�����C�F30�Wl�=O���|���������W�����m�
�O�܇6��=n��Cdx��\� 	K��[��t:�kxu���&swd!֖.�Cyu�ju�x!���]�x��У�0-S�v&k��Y�=��!�|'�<�¢A3��	�0��H��D��n0����f���A��NL��ӕ\�����!���4��@*ߔ��W� �L�yL6~�����@k]Y3�H��$��Ԫ�!��aG{��ű��U�x�v9�'\Ǝ e�q� ��Ìn�r�q�c)�j\I�:�l#�� �]��__l�����0���7$\Gup�lC�9����S�j���r�*R�9������㊱�a�������a�V��<����$���u�˔Jg�cms�-Ϻ�K��n������};Z��3@��_s<�1ǒڪ��!��=1�A�ۀ����zWg";ͼQ��k�}w��|�k�8f����V�:vcQU�=[�������,�V*��h�#L�P���LDXQ��=*���=��5(\����`&�aD� b�Ѳ]��H�I	�������q)�`O'���D�_�t�u������PI��:�{R��]$'��H�T˗�	��v��7�p�2,~xZF�37iI�;�Q���c�}�Aװ`���{����B�g5̜�@o���f0�?
J���ɕ��N�H����H�	b���,nƶ'k��ff��[��R}����-N�B��]�X��,��5��+_U\Lf���m��;Zڴ��H���Ɔܤtw�%NW����|I�c���5��όOw�S���'�l�1���F��*,�`.X��Y�g�[����TR����(!�[�޴�plv�o����>GoDV�cVpO�'���y�\�y�J�������z�&`� ��H)�[�Cr�^����@��M�|W��sR��2]����h��@�*ABJ;��kC"����b�`�>}+z�$��	l��AU� jp�#
�o��ǥ|.��J��xs����u84�a��'ʹoàs���ױx���:D����(|����r�Fc*���mPO��no���I�W�<22���w��+�OPV[cf���-���~L���`W��p���%���rZ^�Y'e��E1�!@��?�	c�v��9|�z<ִK�;	�K�:F'�`��0�7��E8O��Q�J��ڂ~vo���b��C�+�Sp5ZoU�v�ڕ����Dh���7aY�������U9�~�@��?�R!�Uu��u��8�<��q���]�>S�1��\�;&���=�a�/��J�j
Xp�~D*�	���E}a�<3���j�R��/�p$A�?
�����3�������7gb���=Ā��SD$�bb�Ԯ=[-t+h��C��9`j��zj���S�� Q ������p��!�	�V-w&�b�e�f}��&C���*8O�;� ["x����v�Q��c�����t�JzG����v�f�����U�*!�#x�U��t�O�K�PdE΁&�������q��r�j�?=7��ﮈ`=������i%�����/�\R�c̚n��Ȉ=5���{#k��u�j,H����@[8�oY���/�{�.��B���Lc��Xq�y�G����]��+9�$Qay�\�!�$L{�@�W�=e/��B1���N*6��`�3:I�8l�e|��Ņ���Du��~x����=�Y(�u���m�tzjR�)Ŝ��H�n�ZO󰩐ȝt��H��:���b5��������L�+��qD��&��ɵ�(���I�z�ٟx);|Z&�hM�崗0���/���D���U��p�u�F�mB�*Ag���H�B�W����7�co�����#Hz�g��"�BX�9��S���ݨp�PJ���"�����ҟӒ�������9����,9ә��p��TO��*�d�H�ϱ�T<WT��C�����R�EL�u0F��9�5x��}L�VUo�y��å\kM�Q�n�[�� Ȃf�����OT����4��'��[D`*�;��TED��l{z��?�#���9�Q)MQ`Lj���\Ǔ��3���,��)��ޔ�|Mc)ڼf��^@���[⽳�64��i��i5vU@؁����D�����K�s�濕[vI��J��-/���{�� ��e'���7�]J���>���i8����3'I�k)����w4�c���t�N�
}+4�L��9W/7�j�g���L70�g��L�_�J?1�,���֊�0>I���ڰj��D�Ik����s,F�$.tw[b�p��4��6��#w}����0$�!	�K�Mq�-F�	��m��2Pj�q��c |��8Yv����w_K*�ۮ����*�D��lg��
�����D�0cT��/��������4o}/`�;�P�s��=��_q�Rc3O�2����If���]��j����� F�ڄ	tL�