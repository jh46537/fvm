��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�S����U`��P�^��k���y��0�e��ݰ=֮�h����A�x�o��,�.���h�9b�~ֲ�O£+�꼯'� i3.��lU�eg�L��<�*�QJ>���Z?7b�`��b�K�t`z䕝>έ[��XF��F�|:z����@�Z�*��ֲl�7ݱYZ����.��
�$��v�DϷ�\�G<<h�{v6j��;B��e��,D {������Z#��I~���C� *T�w�B�����0�k�Gg�Ѩ�n٩�A�ӟ*YVib�,{�m��3�v��D��pK �/e�n������#��y�A��Ӿ�`�9	~�@��A��UĤ?�9q�-h2�v�9�K�A"�����ٝ7�.���,>�b���?KǗ��W�y�t]_�9�l��\�LK���v��k2�ʀ^l�dQe`��0�`''%\�d&�E0t	R��~�_B��O�_��kDil�U���#��4J�B]D!h�B���6O0"�L�C�G�n�)����\�㘇H=M|�C��d���=�;��R�I^8�G�xe�Ev�mx��~�0�X�i��� Hi��Ê�E ��S���5ʈ���FŹ������3A�u�+��v�uEG�����a�D�]}���	��:�p �6��/�C�h�mߺP���!N��"+��N��g��%<.���z5r���.��H�|��N�#�L��9�v��e�ve�Yf�V�³��pEeQX�$@Q���RY	с��ŃL�Ɯ�y�=h��NE�o��]��B���<b0�X=g�i�sW����W���׼]aI����f�nI�K�D�G�_V?�D��� �&�Gm�����@���̙j}]��Ml5
��D].�U{���Nn�p�^yN}b��?8��mn�y#��٬C�0���%�J�{C�P���a�_=�y��#ה�DQ�ǢsJ�uX�*�%aׂ��Vx�%0���ǾٮeM�!H����B�c�;8���p���6���&Vz���zd I��ݤ��"Hvs�+ę�L�{�y�K텧�WK��T��"{�f��ii����x���I�K�����g�7����
J��`��MZ�[��l�U�P2�4:�T�u_ņX��}c�5�m.�Ta����������o�H��i����ۣ>QގJ22˾����_Q��ne{ga��$�2��QM�	c��2t,��y����O �'��(JЋ�R�k�����s�qs���4�,��Ԝ\�/G�/���}�� g��:�ȋ�aU�R��]̃���A�S,�rU��!?�[ߵ��1������E���=�g�L�_�{��s�*1= �f�=.�z������&]w4-�=R��)6gV����۾�뀔�		�|�!��Q[��eK�O��L��3����ɝ��0�#��1%��ȼ���	����	�Y>���Q�� g,����|o�n�8z"tpZr��h0|�}��UEP�Hf1ts�۸ ��S���=b����l�?Wl��9���e1p���S"�l;�������j����yV�v�-���b?(V��<i[�"�������4�-2+}5�t��t�(E�24o����ɼ�E�:ʓ�86�)#h8E {�p�^r/���u�q��Hx���v��&����N��a+X
u�u 1#ܿD�ʂh�v>Z8'�����"�L����Ύ�k�d�$��#�LXd����݄��Go�����,H�2����>�ڵN�f1��r���Έ�N[�
�qA����'�� ���1@�Q7�>`?oH#�vܜ�E�n��ڥ���"�n=�l~�3��g�Ci�����v�����}nP�PH�z��?���sA�_k����7�j��՗~�.�֙b�O.jX���� ��)Ȗ-�DT#1���6�9S��Z9	�[T�T�� ��煐:�J'�>�ؑ�:@�L�[�l����=���7���F�Q(2�p�b�trC��R:�d����.�����=���t�^��īU7�u ���+쌮�x��U��I����fQ_�[:��w�͵�
���[���T'v�w��>%���x�2HC�����<��G^����H,�+<���9�66� N�\읱j�*�^�A��0/ ��g�}�Ŏ�rO��Q�Ob�Òg����O��w�Ir���p�/��ʤ�H�t���Ύ%)���s����a��N.e�" ���M����ʨ��!�#�=i��4�!�&Bf����7����@QD�kG�}/�����H<S�Z���?�����Ȼ�*b���VN+j�O�:��uI��-��E�� �	��<�"n%���=�/�0��V�$���<����q~��Ǥ#�;
R5W,��%̈́tSb����g$��˛ݗi �s�Ǔ�*�/��`9v���s�pg)[b�D�6�Pi���5P4]S��I�xb�42!��DQ�2���`��ҳl>�X� ���Ej�k8��S�PQ����([t����]��&�<(9�N�@,G���[;O嫕��l�c6��o+�J|��f�#Ϩ�ۻQ �@tt
�n>szf)@�vO��B-��ü�8(�?G�TL+� ���� V�(IJ����P˪:i��I3�[}Tw4���E3+��Xfᄉʣ�)��]B��#*Q��*�v��I�x6���4
�f���ۿEN��=A�⡵D�{v�޼��p����a��T.�a�������߱iG�	H:�G�.[���5K�[�y�f�?@�K+��#r���x���^����tw��n:��C���Y�`�];8p[%h`���F`��n�,�*J���t��"(9���2�z�.�+:���
�3΋u��+���/�wΡ]Lt�愑f�1�1F@�t�yf�}W�\?�n4<\#�Rmliz@���>��_�P��CȦs� L�7RE��+��/	�w�a�
��c�������w$p��QgDL���Ψs�fmƬN�q��V=�,����{85�%�c�T�~"��-?-sa�L��p;����2�����_UY�[(��./�[��&b;#�D_6�2�7M	��P�?�8Vڱ/fuE��&Zrq�L'U�+��F!�%�n�c��SS��>m
h��g&:Z���v�š���Mo��ȱ74���u3�4aۘ�"�V��p���Kgd�DX�ת�P*�t]guv�����q�1��ݾ���2� ������B<���۩�1���J�ɪ-�
�ɝ+�����1���S��9!F��F�P�U<�i���@�\ɵ["s�U���y��r��r�c8ӈ��O��8�&���?_�Or��"+�k�ɉ����4�hIc� �#�����f���cݑ� �I�q0����m�}zu�R��!`�|���\\bs��=]?π�~��<���Jj�&���aa�u�Ԡ�����P3V����I���K�Q����ʠ���3�|�Bm����	��TĜDNn�<��o�R��)auE�Ǟ+a�J�/l��o��)	B7�V�X�t�?�-�i������e�zQ�����'�<�S�:��E�m+�|��zWvri�UG�}�I�QJBDfH}z�K�eh�'����͎��DT]�� j��D�e�غ�z��j&�a8�Z�M�A�+6O��!����:���%��=�l�g��]y���������ċ�����I���_D>��0b��D��9���И��w?+qdŦ"�'`F�>h��Y�W�[bM�es�9�B_��I+�}�|��`��op�KT��E�$�(t���MR����iv�gTR�=���e�8�Q�oY$���b�[$��.�[쮻
Ӧ2W�	C G6��3s�q}ɷ��������)	M��$����@���q�EV���@��������/�O�%cζ����_�fcB���x��f�R�n??Ƿ�^{R_+�OkY���r]��a:ğ�81�� m���Pu@�4��$���Q9�D�(��E_*���$)�E�=�͸�x���p���!�2L���*sE�����ŷfg�|����H-�N�=�BX��V
i~��F�gu`�ĉ������@�v��m�#�^>�y�u~1��H"������$�tU�R,�����u������÷Ԟ�-��0;��Fx��HM����7�r	n<���-���{�Y�����5�a�:ЯK��Eɐ�n%�^��x6��	�s��Wj��T�ߤ��	�m��S���Ap\${X{�c���$y�(hm�M�ɿ�;��]�P��
��lF�x��B�H���H
)��i�P;h�2�M_�ǩ��X���_�j/4�P������v�� ��U����Q��y�m<sa�k&E�Q�xg��F��1QJ���.��9�[�4N��5q&���"炰�[x�fuS|��P�C=��N�}����e8�Il}N7d��B�{m|M��k�AoC	D{�윭D^$�Zl�%&i�l�}�W�,�5��Ѳ��=�S�d���e�q�n����I��i�d~G���,�!��O�M8���{yƃ3+UvL�1^� �j-˚-l;�����bz
p�ڏ�J�>-8�s�4-�}���u���������a�%m ���1@�L
�7:rxb�MjeZ$A�hU�1�G�~NL~��8�!�!�/�ع�~��Ȑ��rG�dl�����P���|��I�S�<���z����#�F]�I&�tm�
Zw�����\/�0M�q|���E��۠5P�C�;���YlG	�Wk�[2�:	3��o�:u�ݜ��s�T�,�ݦ)@�0M�����=�_��,f'�Κe��^�B�@H��\.�� 'N!@}�E�1�O
������d4C�P��J�f��&���S�'���*��O*�X��i�c��ʇΜ�A�q�Ϙ��[��{\�|Cc�����w���|��3	�w�dR2-�<�5X^r��?��6)⃘Idp��9���5
Q���MY���szo�8:8{(�#=$�97d�FXo������Q.~H0�'ۊ8Ԗg��X`/���A�vl�{��X����p���B�����ӂ"v\�	�=J�M,c�,��(8�B��	ҩ%9�
w k�T�I����R��g�_<NjyU�l؀�hH��gzA�O�:C��i�o�@ϳG���@j�6�d;>-C�H4:��30K�o�C�1I��/��*2��(	
\�����ώU-�A�p��v�v��Z�q��o���s&�HX�:�9��1S�~5a�y��$q'�+�?$B^^A�/�س2ߦ]y���,��M��&)撡t?�B[��󘀹:������=������4���������q�̟/��/��wح��[�fCZ�8SnAH�xk���C�O�Ul�V��h�y^�.LR�TB|'�����)��f5^PN$;t�oF!'+
�~�0�Ǘc����Ԟ�O���Y�B޽�=�(���x������Z�O��u��M=Ԟ�׶�)RjԺ����`y�|�}��nx)_(
J8�}&ʎѫ�)H��:�<�b}Q���?�m�-�]�)�iY;3p�X�~�&?R��h��^"�TɂQ��4�@^X�x�����e^��W�-����[����)&ɤ�Z����`����-	�L�E����U��R)�;��[��%�t|�,��&}4�����9gݩ3���Ū�F ["�r�e�]�~x��#�MwZ�l���}�Ώ'�\xP�0����)&�Z�#ޖLP�w�Yd���9�t�� �Yz|��r}O{7��M}�cM���N��7��
�(Gۓ�������Ñw�5Fl�"G��3��A}�p^D!�nr��T\Vm�8:r�Y�7G�{#,�X�2�b3�[l�u�Tf�$���EN��$:�3Cm�KQ=����'F�uO�誄?x(s/��nf�(�C6}�T�_?Nms���',�R����	��Jq;�tذ�EE�f�)t��]7�;���
� (�N1"��Z�c����7po�����|Z1�F��֍�����*W9��=(c�0�q���O�o�3�����jF'�|
?<��б����[+#W+�	��� U�4i�uV=�³D���p,���`un_�S�����@=��n-���5��v6���~��)��$V�udN�&�����H��ޙ��T�OfG󹍫�F75-�-Q1ꎌ.��%��vw�]@�JՑ�ńK�yOz�����9L�<{���~�+6%	��,2��r��=�EX���h����F�f��������E��],�Ӂ3�ߤ���$3�|Y׸
�&��@��e9�m Y��5p;5d�l����{(U�Ot/�
�k�rJ�[#e	��{����W1��9��I<
��ٱ�}�`�M��A��7�	��0&@�܇��L�/TĖ���9σ!�>���l��p�d\�{����:EoM3��c���lڂ\��t^Z+��g����J�C� !o?w�"��	�߇B%P^�S&�������>A˃�!�1�lߋf������(��Au�J,�|���Ql�w�'��͐�0\k:�
�5��sAc���(|�KK�xT���o�O�H��ɐ�Τ���-�{�TkjN��5�{�V�ixuޯ��ޣ~��f�,u#�;�8y9��:Y�1D����=/^�xi���9E5ӔȔ�6�$��� k������ �X�vj�T�n��(�s�N���)�!%��~l����h���4���MZAMt�!�)�-��q���[\U�]�W_�oܝ�푪$���M �z[��Ț3���q��C��o�%$e�y_8՘�P[��]i�@\M�������]���;�~8�FŲ�@��s1�g����b�\���4$�ʿ���/�cKǰ����g�r_�Z��'$���@Sy�ѿ��{&a��@����E�|�(�1F3`Qt^�P�L���RJ	0	*�Z��Jf��uОw[{���n?P���dgF1��n�kϱ ���X(@�����bZ���+�ѲG�3�.Ȭš	�5]<δ�RU�?{}�s_�#9�g�L�mT���w{���;��g2wl!5�3�_^`p�#��9���ݛ2�s�r��P�fWfW�d3E�#����&`�'�s�t2XƯ���O���L�4BqMS动����۔�[��T�r��c�	�v��4�>F	0�s����S�a�2NP�茲��R;7��i
4��j�2^6}�l{�Z��=����&w���OO�O.�\@����j ��Ir3��X�o,����c�sv�FV+�����3�;^lԗ��رM�19�R���}��TA������v�|�뿖�Q@MAٓ=3I��B6Jj�C�-�K��^����L%���T0ҷ]Ruk0�Ls�,M=k��
�y�F����(_��yS�z�ni�G��b�\={6g�%��J�ܿ�,3���������ָ
�&H^�:��@�B���R��)z��.��Yb���T����{�T_��і���7tWPI�k�SSwo>IL+ Wf1Ȫ9TVn�*9G.��}�~�!��q�w��FZP6�:<]*-�C񾆦�c?�AX��- �Γ���g���������]YG�Uwzv��� ĸ�R�'Mr���A;	�x���gk�w!��C:�ÿ9�����n�0�Y۱���JIn�l�T9Y�CJ�M��_����r�T\�V��0��A/�5�H��9�����BF��3���y�8�`�WaԀ�[K��JC�z�ESb7q�P�7�i�Bl#�l-�M�������I��i�&�:��)�t�>Rw7���f�����s?%�_�����Li:���p��t	� m�,������,�"���
��؃���һ��r��n _=`��3�ٴ�~3�c��i��'�͉c��}м�V���Z'ۿ�i)�J`��������ݲyjh�  f�^[O��W1�p�;���s���D��d/��X�x^���]2jN-4��ޚG7�������&R��f�EvS��P*���n�wG$~��D�� `m( �v�k�����(���fb+k)f���e�Z}�9a���<K��g�\1��hƀS�����~{�1J�q���v����PJ<�j�a��t9�G�d1���J�b��i$��\�K�"=��}j�ŕ!\�*�1���Op�#�;*��ZOd��b�;R�9<	��o>u�X�UɆ���Yeu$~�ߜG�!�'��nl��/�l�&�5j�ƩX� �M+G�8P�Vo��L0�jU�J�[�y�
���+"����2�M1�-��_��(
�AL~'��F2�cp��˲m��94ɉ����M�`���%�)z>�P0腛�_@b�VpB��e֤�������cwf�)o�/^c��1G?��sS��U��(���)���ܙtǕw�k�K��V}�a�g����?��E���eřY�֒�o�ȿ����x�m6u��r�|��,.��/;���7��7?��}4 Y{�<K��ՃuM}�����|��v$�e�[��J0����o��(F��	ʺ�!C��\�@T?l��e�|��ޠ���VD2�p��X}�:��G`�6� �C��2�h>Yl�&����[�g�\�_�\�#Y�t����]n��P��3�,�<�Ki�wE�Ó����TJ6�}	 M�U�1z������	n���S���H�f�������(S&�ب
��0���/�X�sT�zXǘ�*���Yߖ^r�=7P0r�f��/�ן����^����� �n�Q���bHȾX�i��Vl]�|�7
��(�1+���O"R��`���H��q~^��
5���L8���zN��T{O)[�Jra�Ƨ6��O��u@L�cf^�o5ԲQ�˓s��$�4k�+@s8�Y�����/ͦu�o��p9}�*�*�W�!�ΞH���$�:T�\�,|F��e���[�2�H�
M�7���g����$G��}�Q�s��a���V��('Fv��	��3;88`�n��N�?�����A��c�vm��t�+�C�Y�H׮�~���Q�'���?Sf��G�E!�gJ�dMN����vHF�G
A�+��5�JEǊ���T�����z�6�oKHN��g�ߚ���a4��o���+����n�Ғ:=�kI����iWe����������h���a!��.�y=dE!�����`3#�M9
����3v�?�K"����M�{�|�������j��6�&3��`9�gWV���0�3�a�[�v3?�� �'F�����{zzF���=�X"dFY{�̬�j���S�稔f }
�0��B�?���S�p�D�����|�(
����������,�Y}I�5n�n�
(E�q�t@�4ۄ�l<�3�M��_T��B5��2N�O-�|��ڂ����Z��;��Ӂ�aN�����r&�T�LI�?5Eۀ��� 8~T�a�?����M��.�U
J��St]�9��
�� U�|ųK�,�W/.�������:~�؇��l"Z�Tu�k�`̫�ϔ���\A.ۑo�Zwځ�Þ��]�_!�x~���B��$�c��;cҿW:��=`���1��at���V�l�6��~�:�v;��_����aP�.��:��ʛٌ�}�����f�HH�v}��H�验">�Q[� =���bF�Oi#g�T(e&@��4��4�v.;x��l�ϣ"F-m]��d����M��tĘ_�ZTo���ڟ�ѯ�t�e�t�d_*�q�1�ORh�=�q��C���LLh���W�f�OE�t�"���/�d��[�D�G�!��
3���R�Ɨ�V*9mN�oS��vY��)�M���=b&z���8)��_��|���i���y��a�=��f@�^j�o �OѮ��j8�5��YG�X����IU��H���^��ۂ�[j�/���Mj>re�	��.SS�J2��#YE�`b�=_�li4��,��i�����F�]bM��Q�qa�<�64�R��BKzډ7f4&������޵

T�Ø��#��H=}_�a�E��m�\
5l�M��6\���(�T��K�to}��O���_�2bU(%���Ra��QW�r�p1c:,��VJd���"�/�T_ⵟM\�/[4�ȁC���a����k�%�H�`ɞ�I�4-2���+��c���>hC��ήq?jnv@�t!�}D������������ ���%���tǝ�%y��/��L�"|BV�'�N]ɷ��d�ʴ�5��i�-Z��4B�j����<�t6���Y��J�ԇ�l��6�⶝��7��K�Эc������cTY�� ��\?�z��#�>�(����uy�AΝnG�>p��o2��"��տ����ܐ��Oj�U����7W��k�\�> ��B�� (�s��r��O�r/�9GA��E�i�A\�|1��%�2'2��F�Θ���W+���C'�-jwo�V����&���2b���f��c;����&�	�f���g*˥wJ�S[����bI/��M�*AO}Ʃ�:���o��~~�$���&�j� ·����,B2�Kǁ�^�*Fa���&�/793��\��/w�vp1��UV�h��2\̼O����Ѫ�H�&������L���#�v�sP�*����ṳu��C�A��W�-l6%�T�sM����hOP_g*;��$lU��u΅�l#��)A.�Y�Y�����*�B�^�z�yֻU���%�F�C�
[�0z6��I��0�L��3뽬�um4����m?R�I�E;�T*N�{�I��M������I��Ʊ���h['�D�B�W��u`���F=s��27�9�CIa�F�:C���c0vf���?�.
J!�R]���Y�,�!1�㘕�h�9V��d�Ҋ��`Z����	�*�1}@7nƸ��2b��pH��	@�2��#2�7�gYTI���������[[�9���N/��Yt;�k�c&��:�����r�4i�w�c7�%���+;���i.�֫�ɽi��\/�� BC��AN?��y���{^Wji1C$_��0n�st�y!����+w�$L�����d1����~����2���M$�ǊG@��.��N��J&1�Ό·����L�c���<���:Zsx�~��|`W�e�_��b��EH�G�y�&��4p_U��]���Khp���X]It�ί��TH>(�N��2+v���j��q_���S�Qͥ�n�F<{(�5d�������+�?��[f�����CU����L`2�*TTԠ�#'h,�߼��j/���o��yXm�,dѠn��TI�:��Aڤ0�'_hRqj&�G	��Ƥܬ�
:����ҍ�L�e&�"	8d��L�G�V�z�1�tUwj/Z�����!.i䆺�)o�X�r?m��,�|8
��?K�	����Bښ̧�;�ӄ�P�h3���s}U��\[�w���C��*�ӱ�s�KI�b.�`�[0Ŀ��~iW�"�D	�sXۦ���g�r������F.�o�9�Gb���O&2W���ᨷ< �b.k�����R������c�)f��D�E��h� kix�|l򜆡S*[�ݙ] �%/+{��	YS�eGr#%dEhj�ap�� ����&�2�l���ϵF�������R ��ۑĶ��+����ʿ�ڂ�*i�朩���]��+�a6߽����v\��_����K�^R�rgDT��@X_R4���V�8Uʰg�UGo�g�����֫S��~���&�Oo�OZ?���S!`����P2����W��?���k|�`q�)°�ݜG�p��w%��ȠC�*��C$l���l�r���^�m� ,_��;��[-���^:�`�����me���T�g��gmb�άѷ�4L,m�����'3��Q!��6���V'�0�A��i�β'j�l|��;��X�%�3З��L_f�,S ��
�C5~eǀ���c�l��]6C��d�\����K-64f/;����a�yG9�1�w��l�+Q���> ���G�X�BV�|jN�VI�7��eY�3���ǿ�SG�5i�����]\̐��l���Cr>�i����9��&.�8h��Pב���/��@�ް�$��{$fpD̎���\�I��҉&�X�Bf&��?�{C�������d�v0�!.���0(�>�-��|F��AX~��uVb�"	��i�q�U
�}х�a0-������J���S0����w�P-���_jh�`��5�c_���!��:e?�[��ĥ�S0���3P&�
�f>�Nɛ/Ę4̲W�Щ���uP?�y��}�Z!)	r;�h�����3�!lUt!J��"�����K����o�Sw ���J�ʀ�d��JE�$�gD��e�梯Eِ�L��XU\��=b���W[C�oTyÆ�b�<F���(�C1�p� z_��#�����E��^�j�|LW�d�]�AJt��nAn-���~��V���W�RN�b7Gڰ �Z\��HY-l�s1j�ö�O�ް?�G��e�ͻ�L^g<�玵PN]1�4B��_�M���3�q��*@)��Ǯô(����ż���X�F����,kG�A:�i%�AE\��I�n��o�:�^���e�F��x4��柺Ԙ:B6l_�'J�]�eG<��fqB�U�ڕ�J�խ�*}D�*qtl{��0k�ܷ��Eβ��@4�g�����iɠ�hz>}����_+����,��1��Ł<�W4\�x��ձ�����X �ga�E:y�F��D���)㄰���ht~R<��-�:F���z�(�w�I��*�	���"�����C������ul%�xʟ-�I��� ���'~���	ų�ɲZu?B��\?��jD
R,$�'1ԕ�Wm��:�
 g��kj�q4[�h8���-��f�c�BXK^���_�)��a�~���W�6�.!՛/t��Ouz���0f�̓�������N��Sوx��P4���.ʝzL��k�l{��«����K�P�$�ېp6 禉�U;
����qw6�[�9B.��\�4\C�`<J�ìŏ�y�HOA`������K:S#a�~d_����|�"qr���! 6w}u���Y��S�K��z�Y�Ь|?J[!ƝH���\�����{[u��T��^�i�l�� ���n5FjvR�c�CT��X_��+��MEM�]�U�ǲ�H��(Hs�;�վ:�Ӧ�+	25������>n&��ZS)~�|��Q%v�"��X��vĖ�ܣ`D6���@j�mw-4��!�X�z��S���L�!p��V�^���î���.����ǈrA/���|�lP1$T��T�G$L�˵���.6��d�ڑ��A��1�b--�2��̴5=-�R��<�in��]�
�-��@��ӓna�t$ׁ1;�ʈ:&�
E}֨m8��l[/����J5��;s��V)kȅYЉ����$z��ne"�{���`$Y��Q�o���0�لՔE��-1?]NnࠎB��`}[�:��d|��Yʱ��J��­��oEi0|Ś�qF�Y��hv�>��4l�ё�?q��9���{���c��'`(V��D�UG�w����>�B�|�������Dm4��Fo���z���x�}��am�^q//�I�~�/i����]&�ԂJ�w��C�9���:�Ϛ���eJ���-�-�Yℕ�()��M\���ʡ�<��˯��#�L�♤��5��C���dZ�I�x��?d�Q��%�ߵx��:���o1ӸY���/�_�!�P���^��؍�n�[�L�j��%��D�5rN�r�hZ��KC9Y!;(]�k$Wq���3>��a�Y\�����%����U�����-7��<"`�{}��Y�
D��S��Bc�M���Ғ��1B�Bb�S˼��	,��ak����N�������u�V w�k��yM�s��|v=*1/I�&@�Hc��c �|Ā��ցq(��/���pC�;�D�9��|1��*� 6�M�;vr�U���Co]���l����oQ�qs�E���~�w+j=�iP-���V��"DV���˗�bO228ڃº��&{��� ���m%�<;�C�z?���y̿m��M8�"2���-�����v;�j��[4�Б����C �~<R��a��z�ovp6��f~�w�U� j��}Uij��n*��=?��� q� H��v�p�`N]���̧��#c!0?,�m�����c-�nf�䡎W�}�6�ÿ�D�%�#)���2��e�zy�k��rϑ�Ew|ߕV��@�M���W	t�� �`�6"#DCN��d����7[�@�ͅ��u���撧��_&�J*�Iᵓ�]����ڑ�F'��
���'�5��7�W�#LҾY3����mIX��+ �p>��ܻ0�%���}d�W��"�8M%r�Y����M�M�'���4w��y�Y#Y��˴+9ľ��N�z�ק�����h�Fk�=�d���0B�{ҍmߺ�{��ac@���)������5coa�b`����bwЯ�]��b7��r�,P��H�zw�^��d�/��9v_��������4�>����������=8BڿvG����~9y�y]��+y�Gs�� � ��Tx��!X�˿������e`J��Q�~b�ݦ�ٕX�E���Jh����y����`)�b�u��Yr����t���<|.���M��e�%�c17Y_�K�}��>���Nxǈ�u�I4R�lU~�"�5J;��=r����|�A@w���u�M������Б&X�i����g�%	J@�.$u�a���!=8_=>�v�e�U�Zu���|�-�����Ng��A ��/���ͷ�k�Ɇ�oڄ��E̊^7P�l��c��.�Cx��?�O�bJ�C/y@Q��픬ގx�o��r�g���݌�&p_{�!��qj}��Q��1�4ݓRZ�p���|�������y�'��"d&��s�y�s�I���+�A��+��9�!��8l��ڦ��o�-����ƴ|H�=�v�i4=��~v𯋥q=͙'$�*�b��Sx�*�@�ԖƆM�q|��ӂ��UKq*]Sm�9�߫+� �,&J�r@��Q�
�`�1�������'��ok�����<Z`��K*�Dխ�2�rb�M���t�1$��
P�	�$-��(�v�������\mguO�E���ش���p {����e�N����@��`�/¶�Z��[J-ᷠ���)/HBt�]��H)CgH�� ӯ�k��-�+ǻ�����2WO	�Ug_;��~ڦ�#��|
�jJ���/��+U�	9T"�, ��;�Q� ꞥO��l��Ϊec�C�ث���R`���W]UD�5��\=�	�*�S���U��R)OjfF)�s�i6HW#B��X�%У�-�E����,6�Z�]-�h�ғ���p��?�c(��,��e���Q|v���� �����7l`�2�����wB�)g���"1'�C�yw��k�)��$� {�9R����ohsT�I(���JX�iG���o1��N��՘��̫!k�a=�&���:$%�
���ޛk���.B��T?�p:JK��B9Lz������/�����E�~m��w�t*G<p]ն6N�i^*ԞEz�"�µzC��m��_��wj�	�)����~�"l�e��� +��$��W:_�3LJh��#Q�ǵ%�C�dҠ��NhOC�͙�rlbv�@�o�Me[�ݦO�h��1�ߚڍ����ܻe�3�`��a�N�BE��抑F�:����)zՕqqXFQ;���6��'�F`�T�6�2UJ���7���8���Xg
���e2_!�1�Q���k
g�pR ��q�^��:ޤQ!(��]o5�w6g��ڞ|6�%#��M1v|s#@�>z��:����R�?v�N��}�-ό54�����ǈ��w����܋474�����
^<�N��Ь��	6s�51��z�4�t�.�d%��F󮚨_#��"�LL���nZ�
����)�z�[���`	%���Zt���g�3��^r���]y��%-��í�� �� e�퇥E���i�E���3f��xHז;j���`���; �����/�j�N-gh�JU�/R.��L�Jś�{��)�xc;P��:�ЙS�8�^��ig��Q�<d1g��a���7rS�ۥZ���(�J��3�zB�ׄ���}�.�A�"�lPIb6�h�o��;x�.'D|����a�g����^�a�l6ypՉ���R����)�S�Y�w%�!C,���9�'Ό5���ce��_7 !gAI�a'���+���wH��urZ),r�
8T>��	-�DU;nB�پ"`�pU7 I�43�`A�Hp��T&5�6;I+�\�g�8��Bm���O�O��w!�ʴ`Ƞ+w��mOlY�G,G�3L�E�ڰ�}㷈`�����ŕ�����ox�%G�r������.S�v�"<��#��B����]���[@KX!o�2o�1�SU-9+�N�����u�a�'��:�{����S4���ɫ&G�O�u�}�d*Z:v�,�ѽၤ (��^�p�V׷-c�2V�86Oe�ߡ�c�b��e[q{ �z�1o�����a��O���h�R��H� 6��F����;�^9�t��:��17�E���ʳ���2�Z�ѯЅ�'N_4�_����9m˛�k羫�E�'�0n�lQ%J����&�1���\e�&}�!�o�Y��H]h���Կ�P�G�>Bk��-�V��F�,�IS��g�{ܑ�;D���]Hټ��o���P�4k�!�u�|�w1�~��������<6!��]�h�5YBs�;�f�K�:�XM��*���2R*��${z��6�#����v<����ߣP����k�]|z���wc�+�Z3n'��TA�b��#�Ws�hѧ�D��]��A��,���]��;V���	n�	&����W�A'�ʶ�ʪXA�R�t�ӝ�!t����u�گ�)�ѧ�m0V����-O���&6Y��ϛqf3�h-͸_'������?��6*���פom��tˍ�J�c�UF+"��WΠ�E� � �a�	.����	�\\"�ZiKf�[����9
�	�)�á�K\��#��E���R`c\~q2�fr I^�:�����O�mz$���c�΀��Cg_���&���/�b�M��z�
Ѹ%s��z.��N��6��xʼ} GiV7"�������#�/�:�Lk�>�@�?�ݠK��c���)��t���5�C�.�i֎���Sk&'(��7IδDT�����Q
��k)�D���aK,IJ�O�ٛ�m��Z��+�R�SY@�g����H5̹-�Ϸ]�y�t�=����췑��i����f䝒eJ>J��������z1���d*\g'��량�-�+'�rJ����a�v��/2/a���:�e	b��;[�f7t�X�Ƣ�gC��A���ɂ~��ub�>5e7y�Ѝ'�Ʒԝ�W�iV��r�t]H9���@�v�oD��1*��$�v��W�z�U2�x��Ɗ+�}��0��	�_a��Kh���
��{H^�y�j��g{�;1�a�Gn�YŃ��:�ï��+�E�=��kO�jC. �����k>���ů�>�[���KYu/�!��/"<���a�pv�tm��V y[��Ĩ݀�,V
���PK:��1�^KDb���P�֒hC�o�Xԙ$	O^����b�y=Wl�|
���v2��H�a|�~��T�hډ��C�,à��(�̓P�P��.����<��pG�V�||1�`ՋT�f���:�,����Ə���53Y����4��[�멇������r��l��SЉ��u[aGq�B�h���U��n;m��x%�sW-��8��&/f(M�0��
�{6`{e��Q�]f��0]�)e�7O��JF������*���c�k-���<��2!p;@&F\���DQ8�F��Tc��k�[2X�4�p�����:���4B盀�(��g�~���Y�})=)�����!C��T,Z=
���5�rC�kw�r�͏!a�1�	�?g����*�b��T��\�j�?R2�(��۩�k<�q6M�gN6}6�"��^9�ʢ��PL�0���J����U��`~tZ��H�haXw�:|� ��C�5�����IB��ߥnSVo+�Xb[�G[�`a�;اc{׮�@W��8�	��>��O�!16��f�+.�MV��M�䒿��9M��.���Z2��2�� C2�x��"�Z�;��n�o���r���č;���\x� uoA�KJ���Q��u�����dS�'9qC�,�w.A���d���E^EDAq=�����^a:��@,���*���E�I��1�����\6�UˮT_Ig_���GIt�#�A�&2էU��?)�F��H�	NŦ�+ht^|�Fɴ���t������a��e=��S��d��#����'���'�*�Ӊ���)�eB�M���6;9���z�5�a7qs����l�SK-�Fd�)��/��삺7�G�w:fO��7Q��J:���6�XO#�;h�ȺE�j��ΑE�>��^i󣮍EV�Ǧcx��(�]B&��5,w�ލ���Ԫ��N2���5$�X�����	�h�ު.B��5���5��m�0������άJ�
�9o"����ф��k.[̞���P��L4����ԓ�Q���j�+����L����xR |�h�:��P�X�I����O��Imk{C����M�N#��YU��*�2!�L�X�n�e��.ӟ�� 6�J��I\FS��_�+9�q"���9�q�IC?��`�0J��f�[_K���u�K����0�§���%������<�e�$��m�܎��
���}�u���ˠz;珘m�ϗ�7B��rĭ-S�D�J�5O�Xq��vld=?���;�<�����M��쳸���؟|�	n�v�k�-f������%ݦ����	ɑ]��d�~82`������8�m��ɾӧ�=��'U�<uF��U
�R�����&�n`R8����v�& ��h����8�M�a��DU�OFI��L��,'���`���,5$Bp��R;go�-��*��tM,����q*� �E�^�q�Q�2�2IkRG�����KӦ�n���䦂3iu�a�
�y�.�@;,e�u�\��{�d����j�=�w�F+>հ-{-�Ni
�r������5�(�'�P�9{�Y�q�|J	�%-�P:�
X�N~萊$���k#�>7��#٥�;�6/�<�<�4�F:�?���3V�$�V�P{WZ,��t�\��w�1IG���~9x^'�-�海:�T֑�L"Z0�p���%�յ�F������@�Pu�����zX:������J�9oy��uE�~f��j���Y�9�l_m�O��jW܁��0�Y�b��vKkG�r󗎈�,XKf��j�����9[�SD��%�8֫{�˿@B;���8!�"ԩEn;��'aە�ݸd���I�����ƅ
x�Iy � ;ӫ�\��A���$fc���2��ah: �"1DsNMP�v�Cqs[õqJ(r��N�+7"��E�
��>�zi�=��S�א����$��ʤ��A_���<���yŜ��� �����!~nf�)�W�N��ʌ�q�D!�rܞ��*A�����͔��:y���
n���c�������E;Rb�x�=�f���r��sK.�+ߧ�ZG�`33��,%`A�?��͔9n6�t�� ?]��I�A�%�k��(�{i��&<Y}��m�
U��8}=�M��x�MM���.�J��)�i|��-���F���^�u�l�����ې"�y�^���Ua6X��/�\��^��U�aIr����_R�	$�6�u�ir�Χ�j	�Q�Q��8�\��j(X�b%�D�<�B<�M�֌r�"#R���#"�qu+�\�2F��YT+q�Z7Ĉ�����.*H�W�n�B��L�h�׀��I���������~P<D?;/t��G�cI� ~����s�{Q;u]�g�^,u��/Vi����`�Ds�:̬Q��pa�)���}<(��^��S�|%������W�Z��;�2>����<��/���!H����خ�5	���%�>C\�-�/_�z\YuĽ}�'gv��K1Lp��K��-�ۊ�t��3���9.�Ե�=���a���*%@�⮐��Q�
���yP���+0jG���~ܜq��;�Q4�Ep��Y{%Av�H%ܭ�4����]�(��f�}�6V��Uu���0��ne	��U����s3�SH�e��b�a�µ��dX��ԏ�j�)-�P?DIAH���9�-�~(�bp���N�Y���Sh��S�+��R8��5'6��M�*�b:�]M~���`�&���@,?3��I���Ek�K�k���z�z��?����2	�Au��n��Ƞ�>�3Xu�Z)H�|���Z��y��ɱ���G�0�n���v�
�3�?5Č-z��r`�ۚ) ���$�;옴��-˱��E�+�������=2��DC]#V�o}�2�'L�Y����.y��ë.�la�V���-@�y�G�n*� ᗉ�_§����PN�W>;�e>'�>��e� �8��Ǌ�\���};� i������4��Z�M������- �\^ERPE��j�D�����ns���Հ���"v�����i��p_�&�oYΐ��V���K~�*��_Q��GeH�d1�
?ɺ��c�T���pb�ծ�cܬ�D.i�����Sȇ|5N��ږ�H�������p�#�.����B��gO�/7���s��fK��fy��+��K����������Lű�W�K��$Y�(�����.�;!�YW1��N��\�'�S{(ƛq9_��u�.�8�P����T�ݰ�N����UC@��F�o��eD�z��j�	��_��J�E�H�>�?�� Oco�0ls��**���z���u�
�N��uQ��K �nN�O�kc $4��dR4�u�$���
���[g�o�/=� �hh�-� ��2�����$;I��C��.ۈlO��0���h8�	�^I�1�C(1��v0fݽ�r	�\��=�f�Ԭi����E,�j��=z(C� >�[�0�����Qv�
�$�n�U!�kz�Q�l�D�\�_(M�U�M9���P�/p��s~z�i?����}�ەT¡� j�xu9�ާ[`AG�^^��oĿ��6H�E��D�=!3��n�6KA�s�Og���>���S5I�W�4T
���\\�}�8�q���
R9�d�(wE�΁
v���0`��;�|��̍*�WKN	�Kn���/�3^O��1
?�PS5�*�?�c�_�E��I%����ӹ�R� ��b��Bg$W��	.o��|_ۻ�[5����z�쟖��1��T�[�͈�
dI1#���GP�uf�O��T��?6��f��V�[�)���������#�tw��Y�:@C1��*ۏ!�?���k	��,�3�."
�h�k��PZ�Bl���2@M�\jG{�4�ҁ�I$$��&(-A�ܐ.?p��N��J�����@@����h!9mgTS��m��|���~U�tQP�⩤��N��Z0��׳_��>Hg�L1囆6ę�dP-{�B�Go^E*�l5˞�ݗ8����"� �n��y$�5���*