��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"�.0�у��u���D��@��-5�׾�l��C(�q�����6�K��j�� PkX�O��N�ctL�>��|@OT�'��"5RH���af��W��.N�&IA������Lk�_��O��T5��agfv�a{�n�d��C`IF��"-{��Sw���<=��ݺ��W�~t1�}G��"z�⃡���?�ej�iE��ʚ2���,�Z��/B�ݦ���ũ8��������`'n^B�p��KcB	:i��VS�9��G?�|�}|�N3��Q��+�rmU�ŝ�$����'P"��lG��Fy�7	�^`����J
��T�	��*�="v�ۄ���?��{��nwkS�%��.ܖ	Ws�q��D��T�"��_o}v�sG�-��5����iGff����^i(C�9uʘ��ђa����oL`�M�'VM�Q�ɩ�F�t`��~�X)���ThjU���Bb֎91&�&��J j K��!����Q��}eL���σ�gdh��}K�F���D�G��� 1J2��|a7eR2r������ o��?��>UFs�N0��OsJ�ai :1X�\�*VjDG�Hs`�:�p�S����_���ӽ͢�K']e��օ��4x{+�|`@(!Ίݹ��a
yY�ķPWn"��DQ��R@� �.^���ì�&1;c���垎,t>GϢm� �^��&������Я)wj'�g>#8Z�@���<���_פ�L4�����W

Q���+B�C'��bcA��8bm�1�Ɩ3j/@:�k�z���r��7�ΰx�N����l]���fg��Wp��[���sM�pb����=���:��x�	J2��d�3ٜ�An���Z;�X^"��MuWy1q ��ol���r�MW������>Y�c��_DBJ�A&���D���Nb៮�2=����9 �Ǉ��Q�}�ZJ���1���b*� Q歼T�[vB�qd�㓽+�.���
(	��~�BM���F�����K���l`�Ʉn<�ǈ��?|I������[�쉌ܗ�г�+��L��G�&f^C��7+���M#�!���nݿEo�s��a�%���,-����'z�<42�ʥ*Q�@M��b]EɆ	ױA�>�l�]��\�~�,}^w�T1� l��I9z� i"ӄ߆U��A8fcQ;��=��v�=?�*�~���D�
w�8�U�M�6T�%$�����53s9�%����<Y~3gvŤ�A���QPm�à��<I֥��	.�!5nG��<�Y�	6����ӭv�O0�2$�&!��5��uM&4�\����Hգ2�>	Z6���aW������OҚ� 9ʫ���buW�������8���vn� �DO�5?t)�,��9d�'WX��<�`��c��A���{@���\נ����vl�T�axV4Ni��N�I����u�I�����5(o�������Y]�CMu��(��֢d���7u%ti.���%n>����	Dfp�Ej��C��м�>��V39aHam�i�EF�P�UU)�~���(�E%���J���*T2Rf��0��9�*SCua�Ҝ��4�v�Ίp�Q�|�����Yf������4�nH�(�ؽ���kͧ����˭�;X7V�O�iĆ/f�E+��Y�Φ��j���hs�W{�`�0�L3�=�i�v�k�Kk&��o�>O�mܹ*�s���c�
��鏂�X
��T�
:�%َ�����H"��� C�+= U&����9���-A��!I4�m�6ᖗEc~�V``�Y=�~>�%V~&��k�CԸ;h�#�L&y�}�<ؗ�&d�����'�+xV���䲺�)�����	d�|�;<�U#�m�����$�L������Q��#2�#�������!��K6�3��L��P�I�4��������	M|n���Y�ή_���*��������h	�5F�����v_�\?'�c�Z�����vH!Lf��d�p ʎ���Q�XV#���Z�z���3��.rt������sҦ��/V�Os�C�.��>��;�W�QLaZƴҊ�Z$�!�����k"���팘G�jR����������0�<�J�	U������>�����^,�>�X�k�(�&X�5��	���І��Î��S�mz�9��
Nݤz�OZ��b�XL4S��$u�S=92��̸��zD�Aަ�hivJT)���~�l:���l�YU5a��� �t	�c��&F�����0�� 	Q��ƏH������ĕ:�3��o�����s%��;^b���1� 3�ݍp���	���?��8�;18�`���3#����H=���r���U
�VuNm;�}uWb�."�Z�	a@�b�L��|o�V��_�Ԩ�-*V��ӹTJU3^�h����[L-O���Z�豒�5L8��`�6�^��d$V�UR-g\�7��nW-)d�O�������6���:~�rZa�> ����Nu�U�W����$gŏX�Z����Gޠ'xM��m��-Ň⮟ӌ���Z��LU+�=�DrM}�]q������b2�H⩐����ř�����g͂!��rA�������|.@���0�����>q���>T�������
��	׿�#�z!1 �3y ~=*^�z�L�y'9���=|�՝)��֞��i(H7�������ŭ%a��ij��i��v�
Y��!��J���(��T�k�Y�VQ 0>���)%.N�w����ژMl�0M�B�:�&��8�Z��[�\�j�A�7���L?{m��
���D�Nw4K� 5#���cJ`05k]f�:̛�?��'��i��%�Tkx��M��/� ����+x*[6c9�g
N�gɤ�˱٘�m֙ὗE9��	�VdHa�����w�Ѡ�����Yts����x`ձ�g R�e7$?���x��i>;PJ�(���7�ʰυC�[7`�6��� �5�t�B]U��j9+������@�"���,����?������'�#�.k%�e5B1�ƴ��?��7 �s%d����0��@=�+��	�o/���w�c�#-�%��}1}�(���vT��qʶ[M�H~)��xY/S���D	�>��V;��ʜ[�[����G!���5�{SE��4gV�-Ԉ�0!�8u�[9K>�!�����s&�]N�o]H�rj�R�|/[��l˨p����5��q��-�čؤ��RB�t��K�j���P�o�^�-�
���]>�����Oz���d��?Y�l��H:�.I�Fϒ&�����NW/<ԫ�a��$A:��*�o�>]�&�v��� ��u�1B�,q���� �	Cf�f)��<�RX��À,7��,�'Ԝ5)�F��Q�t�y0l6�r�M ��� �Q�6;�;���L���/�?��ɶO�N��Y���"�L�'�sDi��
�v���-���K���T1��R���'���r�0��8~����%�Ў4�~��"����o �#�kz<��C�O�j�B��O�Q�߮��	U�f����VG�}%�� �G�rHۓG`����|x�}��2ҩ%S���	��<���5bv#Y�r��1c�����OQ�\�7��ASx*�>�1l���j�]���l���<g2MEQ���_EP��f	�;���Ģ;n�嵖>*sW�8b��Ç05�I���WT.��N]��
c77�Xu|�/6��вʂ�N5s�;�!I|���cZ��q���]ʂ�=�+� �J�����Pn�j�E)�E�=��y�=�M$G��0(�UٮĿ�@4<]���kSj��1a�� �?�I,~�=2!�E�9r�+������"m�ٹ@;v��<2�ݞkoJh>4�u	��ɍ\�4/�K/f�Υ�VsF����Ǻf.��Ճu�w��-�?�����c��Y��]kH�w�!��s��d�������=ĭŹ��3c��s�e��lu� ?��E��o��QL�#��9y%�^ ���)�:1�hRs��Yf�z�(�zNS2?�9���ԛ��.�O��h���Cl�I^��Q,o��|�&/��3O��nƐ��`�U.��eK�>6��D�/8߽@�'5��TJ`ݤ�����>��,�Iz�k_\|�$&�pz��%�>bwv-�ț]�v�
��7�>?s���t����#jh����������#�6Ȩ���_��9��'�������'��?�����N�������E�a�f!�W�:j�TD��ʸ�\46�4�C.� ��\��&@+��G���E��nD�oE�Ȁ�Xm��(�
ыz.��X(,$g��ccԦT���.]�:o���͚:��eL螛������7@��+�`�EE�0��7��zn8�h�]�bm�+��Wm��pF�)wJ�nȎ����6Y��}�p*g��BD����1�.�`�T�d]�^ w����ť��`W�~D���y@��[	)H-���"uar�M�h
��.M���p�����0�vb&&,��=����eI"G#N.���2�Fa`�n�n`lg�yt����$0Bi��.àϙ�An���� �����A�3����(z�F�vqy69C���?���)������V�G��{��AZ䥙m�� ����WN(��fT��$��F�D�3��p��o �U��;�J:�����!��$�+:�%\���zr��:���w����=���M��ȒV���{f���Gj��R�R4�B�m~/��G�W�PR|�����bX� <������S��{	�9r=1`�h�e(�դF��̢e*�d���Y���g�6�\'���W����+� ]��BL�N�mxHt�Qn�n�3�D@8��w��a��l���OWa��b�.ʌ����;�"}lC�b�Պ%�fҔ��t��e����;zHRs��L"� nl�k6n��������Ҩ��8p�w1�����{�?I��@�g��y��J��~v��jq(��:v��$<or*�ܮۆ`h�%��]C��y�TCfqF��1�����Ѿe0-޵�����@��Ev8}�G��&�J��(�p/�?��N�@��b�����{�����r'�i�p�,#w���j#���t��4"�7�^��d�@;���F��A�3�E�EMĦn>�,I���]4p8�->l4�,�!ڻ�
2�Y� ��!zȼG\=�d4&��2���4��"|5�k�p�]��d�7�D#&�zHR��9�S��~h��t�/�;V��{e���S�����[���r#"�=e�'�x\ޒ������V���ӫ�w⫻'k��#��� �ٰ!/O )��S� k<�P;��ԋ���B
�Fѭ����/&��\�y�<Ç��S�������+ (����3���۔��,\�Id��d�k�Wz'���L� ��q��`Ϲ�4�=W?��w�p(�Ù���ѧ���� Ѓ7�̞�+���6HSS��n�R;��ڋ�%� Me�Od�H"v�Lͩ��b�u�T�]&����T>���	d�/o-h�>ZR�W��Oo��s�'��E^uJZFڿU��Ev0�L�"�����?=�f�y�Y]�>Ǒ2;ƞvI�>�N��]�i=ځvȽ,�j�|m�i\Э�<ӫ?h4M���#�ۜU��9W����5Q�Eք��%�e�;Xs��X�2I;1h:�p���~�J��{C�)u��N��.�K����W~o��5X�L��_�\l����[>����w���-Gö��Q���`O��_� sH4���x�(9mx/�nD�����K൱=��Vx�x�$˪��1d.���/$&�vҝƷ@O|�3Y�[���n�x�?m�`π�f�k��qfl�D|�z�5�&�{n�mg-)����@'����%$3n�̰2����Հ</L8�,�w@+dd��f�̓�ʛ)���&�>���w��B�=��U
��ZB�H�ɪ=L}"�o�Jƙ `��� �덈,�hdg�
Vy���4 ��l�БR5���Y	��+��`onX�6��za���??������^9s޺X�m;����&�և b���.����5ECg�m���gnH�_�}͕��.GT�80���ޜ\�e��S3�?ٕ��H�Я@���H]XE.%���˯����sV�S�q�H�E�x������B(@%�Z���ѹ]1@:nh��Vd�9s�]kG0��6:�7�N��I�������$��K�}���=TiA�jM`XR��"[2sre^���$�FW��p6ob�٢��V8��+����
��\�B0>�nC4Q]i�|�.�_�ݾ�����Dl7e�B�C�:�Z9]�K��U�cZ$�VC)�w�UE����Ǿ2���WK	�`Oj��qG�Ј��Ro��@$<%Mp����_��NaJ;S�>�{-C<�;z�x�����Z���F��Oc��oO����O�r*Y�3�OuՓ�F��?��W��L�`\B�c�*	#x��o�_��p�R>��I{����� ����T��.4��� ����f� j���7W��qs}�ɔKN�.�^�Q~09Xw[B*zzmQ�{'���wd"�:�*�
!��R����=H��kH���a s��ǻp����Y�����C�V�7�zI��9�j
�GDsM�>f�]�+��(�8M(��1�#�?�_��M�b(zB��(�(��m�IA`���by�!��ʘ`,�s��ݙfZ�戴L<��R������}���N����[��!1H���Gy#�4�d"���	��+PH���x�������S����ˤ���b��$Y����h���0>	�����D�w�W��]̕�IQ���r�#��+� �}��W�6�m�����:A�K��<����@5����.��[>��M