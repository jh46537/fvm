��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)��4��S�C'���Az�V���g�hN�6���~�w��(�,곗�%F�Q鲀ۭ��m��7[�S��������@e������:��m���9�����e��L� 	� ��xl���Q�
��
��#G�A�A���CG���a���+X��N�b�T� �Yr�F��J3�,x�յ�5���F���\Mf����U8в$	T/��8xO��3
yo�x�����E�Ҡ]`{?�stN���4t��� ����@�70�UQ���*�=N#Wnd k���x�^��xr��?��nm[y,@1�1�NQ~�k�����J�g��~�ճ��y�b��xP?D)���|% N�AS���:AS��^?C�$i��҃�iG�[,%.�l1$1�׬��\��)Spkٛs�6ڽ7����0�
���j;�W�F�x���>J�:�F�1�C�0���H`&�}t"���0�<�+iL�)28�\$1��˖ʊ��<R
�A��/���>�d�oc�Q4B��=m�@5�X���e�m�cB=2�܋P*�g�b��=+h� 
�(-��S�}jn�[KS���=K{��|��44	y��\�������i�=�bT�<[���Y�������.?L���Q{�>_[��?���e�0�KN	�k̡��k��c��9�,S6�@�8�2�	���p�+f����wDI�7!��
����G{���sb���q;��_�a�*�q�NЮ�g~k��%r�����K���swic!+��"iQ������?�E����gJLeGE�5��Up��Ͽ��Y� ���B)8l�I�^߹>m��(~��!�}N�T�Y��w�.RT	�|#���k?�y��P��xw�ڣn��{�g�u��IY.����Z�`���}��7��'��!� ��Mf�伫�1y0[9�9�>��5�&$�$�c~5@3>��3P�A�J4ŐC��ڐ�J���A��*j�uұ�!�h�m�:}�Y'�t��}��O����)��O���Z��8��Av�x	r���� �eQ%�g�\�5�+���mS���k�m*�2�yv�38��ΤL�������6�du�-5��6>�$>��E�Ù����}4g�h�۠v$u�g��t�s ެ%\��Q�ړZ-���	�q|>�w�y��6R�r�O��f�(�S3����H�.C?|�����6�_��^�#�K?�/���9?r���ma�\�c�r�>����'
!�cC����&b��wĵ����@hA�a���ϒڍ(��_���h�f]74�u��K��-�eU2i���
H�y��:BNb�2Y=l�������5D{�@M�~f�W}�m~ط����A�u���S�n=|�d�� ��Y>BW���o�����5yUZ,�����XC�]-��K�����z�iQ�=�B} ��]���[OH�A��Ie\����(�=�3^���R#�nآe�ra�豈�GQ�@���r"��p"�yĿ�A�r�1L�R��>�C'  �j�x��j �<l
,e�>�Y�o|��uz�c�cw��(vvoA]�V?���9݄-?h}��W��2�a��V���aU�m������A��B����Qp�,͏��~v��3-�ڑ(�#7�cp]�ǆ9(��A�qѴ�|	���<q^�Q��Q���6(SN�?xM��y��v��,rSg��&A�I߬��#�i���Ŀ�n�����}�bow)�WYn=7��J��Ҙb]Tπ԰Z<`+��QT�7Y˹ڌ��G*3���H�Bd8mi��e�>GH�"bGR�������k]�J܁��ʩ��5IK����i�
�� pȱ%
^.\Ha�z@���^��)��ac&��/�!^kJ���ӳߥ;{�_�Á�{̒�>��&�[�Ǿ]���+C�}���vf���s>�ׂ��eo<	�m4֗�% nMD��k
�����\�<,ztD�)@����Hhb-¿\�~'P����@�+���|<��&�T�:9�n	�n�J�jG?u��F!ӱI�ׄ")�IV\�n<�y�)+L'��<=���'`\���v�wle�_�^bIlm١|�E���*�Hn��?TV�)�cr��Oh�Q*3�����ɫ����}B96A��?�F�/]v�U|�DB2YiPI�� ��d�h����(Zo��|Y��kB¥�2��+R�zx�.�,K��- ��{o���k�>I�����G�NQ7[��/�߳-R��I���!8"������:�z��H�}�(z��8u��̙r"�p
C!�-�B��5�vQ������d$6�3�i�������`��^�Le8��^����+O���5]���erÚ[�v�`ˎ���B"�hsUe��`�z_�����W����BN�}���^nHw̿'a~���V��R/Lă[FZ�]�bgs�}�
ԩ�,y�|A$��-��"���ź�]c��wIq� sY0��N���=4���|z���u�OQs�
�C-pC�{P?���g�G�� ���4�!b,(�o�7)W
Qn� ���d&�ŷ6���&��S���k-N���� �p���Y
��(���t�����&ݘ�:�{���yY��W�^�%����%h��P!R�8���=h8.?�=3�7��>��9���Ԗ����b�/=�����(dIi �V���p��ܧ���m�~haX��*�>�AX�F{"��կ��((�y���D��#)�r[}��BElw%�I߮�7��f�|�Z�������`��Y��G��x��ْv�aL�kÙ����yn�M��5�IQ&�)�F���TZ��wfE�;YDOB��;��F�%Z�\!���}+8�����(�y�����';����i�qlR:�*�H�󌅜�W����.�>�x"�#5 �-`mvz�?w��e��ϩq֥�q��OG�> �������n·��=M�ݨxxtD5fb�����)q��;[@�/�z�3�������2b�fR�?�0}�FRv�y���Z>�}��z��X���
�m��G���Z�k�1��DmT���货��9*�7�?w�kD%��wz+�sǡPT8g���$�6�(b���Ζi]&砄�Y>@% J/B��D�z*gH4��+�R�t��Y���=�0����Y~�s�������F|ϭ�P��dr�)�]�E=( �nJt��PY{z�k��h*l���dj���5��푗4r���OL{�F+���1�@�p#�޾x��w 䌅��J��"H�ڳ��+Ёze�K@�$�"qe=Qx
�h�2�`�:N�$<,fn;?��L}y�,��2��"�wb��/���4J�a��=�[K+��R�In��#c ů�Tx~c�;#>�Rx:~Eݺp�#�f�F�*(�t����Ϡ�݈/���##s�ED$���+h2J�����'�G�cJ�N�XZA���{�JD��I)t�t�u��V�o���'<��yׄ�S�'���r�C]�iEs*�(�]�Jb�� �b��Ao��3E�C�&��R�&}uw���;��挀U�hKYZ���R�C���ݢ�C�1u*Q��5c�эy?���ȬR��0<����$�z�#�C즴�:�m��/�\Ҵ�Z'#���/ZU�|=��M��h������\CzP�ѪB�ם]�h� �O���sy8��߯i��H�i��X�Vƙ������-F��A	��L�Q[qq6��!�&>|~�HZh/M?:� J�Y��ߴ��{�W�K��,�7�|�C滳I�T�s��t�L��as�0�������>�?뜡��Q���T��ฬ�`p�0>���/�]���t���I����~�0ˌ���tߏ�~���I��ߵ����Vg2'����� ���5���@����>����h����Ẋـ�3����u}�J[ɝ��=^�����Zx��T�9���w#�ν��uZ���_6T�Kڵ����Ϸ��O�}o߸=�r��l��8fb2G�Lz0�O�\�@���c�Z���G��M�zݸ�<,!A���1�#OC��y6��p�0�H�����	q�2��~g.@�<헻�[�mPM�w�&��0���S��T�;�'��a㛢�7:$��'�bm�&�F�[���"v�8��<�\�w_���zAM�L:guV��;x��UG*�ƣ_0��8$$TkG��}��Y�8��&�D��q�HJ�"��3�v��9�o>�R��F�Y'�t׻w��z��D��O�P:S졾���}�w�����z,k�s�GN��d;u1}�X��7��9X�hN�h0�ɶP$n4Nt�4�� P?�%G2�Vv-�q&��l\��GB�G��f�!����i��R�G,4��U�.T2s~�|@�]�p �̀�����}�K@D��O	�"%���F����O%������]-�	�c1t�CbT��G�Us?�;d��H�c�;�f�1e@u���^u"9� *Ț0�(�y/���gt=��{�C���жwl�2"���c������+��1x*x�H��<q����@~5��������f@��,�L5���u���D	�5� �}�!�!�&,qbx�������R7�qRUY�i�ߣ�	,<��x k��r]J=��N�)�$ ��ٔWZ�վ�f�j�
��;ls��Rk)_ia���.���u�V�����P��P�#H@���m=),%�D�糞�s'X��0���ɵQ�	���! ������F4����T����4�жq�A *t�=6]%߮+WZ^���X@y���q0����x�`�F�ؑ�ɁeɆ��Z	�� ��r1�&N��$���٫�w�a����^%0Ю�,�gu������;T��Ĳ��<r�|�i:�m���ߕw@�A���?�~�w>e2�'�=��.����E C|���-�z�HT��LI2�kPJ�
��η�]�hS�+^�	2t�,�E�ń��O�h  V0^� ���h7����F�p�l8�'���(��p�uQ}:�Ci�gW�_�z�ݚ������H�Ӈןh�F�'����<:{U�HC�7ɹfZ)P���۪����BQ=Ms1��<f~�}���&�(nǤ{
���Z��8�M ۄ��M[DP�0~����u)�YF���X���V�Ѿ/��-���߶CM26U_�"	������DV�hV��m��;!�0,���^r��^���x��Z��e�Se���ZX\�>��
\������r���ǀ��o^��YSMp��ڦ�DC��<���i�2<|l;�2=�W�WE��5-Z,���g�a�����_�XA�.;�$��������Y��:h�6�r�ry]Hf��A�e��:�����vJ�LJ��u�8�E���дV��Q�$�m^</�l\P/^���?��9�)>K��X�x��ٖ$���;<�wa��+ָ�T��������6��ɟI���nx&�ze�I v���ΡI�p%��! �b�x��k����t�)}tL��
�S��U�S�H<+U{����9�G�RT�j��؊�"o��l4�I��x�=ۀ��.��k��-�9�L�ѝ��M�{��1�mI���zɠ����l���#�â��O����(��AwԌr�\a)Ai��C}p���`4{��'��iu.�Y�{��"�'5��]�4���QϯB��ay��܈��l�LuT��,1(e�8�&*�l��>� �qM�Ao�8���~����?��.�`*�J91�k�=�w��bE}�wna�Z:�.PDAy绔���J�~@�����ֆ��V���+|S�a��2�W3f��ĵ|��:'��-�1�����:I�C�����ϩ�c@��c(|��Ou��cv�^�7�in��9��ڲp��r���3=
��X��;�G�Gs���=��C�O��^w�����g��u���ۻ\���:ަ�� !��É#���)�S��{�2�	�+��lDWf��Y
�Z�S�p�#"�Q7�x�q7�S��Y���U������X�A]��}?�ۤ(T���.|�\�	�D����>!r�V�e r�/�@%�0�=���4xq�n/�
	LZ�:�6g4�us!�hԹ����6nn2��Qq�'���2_N�s��¬����^Y$�e{E@g��YIji9MÔ�yr�8�t���`�����1�:��%::T�2y�`����^��ZUu���HV��J��oqF6���[�6��:��� M�-��Jr$H�/	�o>bG�*�O,�����\L�E�L1�/J�T�� �#Yzu��Vk�ѶmМ��f��D��DǙ��e �M;1/{��w��3��4��cg_�,"Gp�h�j	�EP�j0�,O������0em�sns�{��`Z�F��7C�rO�3��'lD<���Q]�mQmf~��dx>�<L�򳴺˺T�[H�N��òDlιޯN���������"�oA]�p��Y���Z��T'A��z�P
�@� .��zq�#�A�!���t�zW�*�^���kI��2^U�XN��!h�>����4�gAAD��TjO�RHA�}�0z*=
���ڦ��~$�'�{�|z��xx=.݉K���Y���������������w�[M��u��>�9?ȟ��sj�-��Q��\���})*:t{<$�*�
FYIA�k)��� t��T�<���)A�% `8���*hs0b��ċ�'1�~p�C�w-ys2��X�7M�b��O(����b6;�ߕX� �)0��lL"��$�=*�?�/�^�W矡��j�]�˵_	�]YX���Vr^M^j�D"8&[��5�@UaQb{�n���a᥵·yF�_D�h�jg�őKc���	T���$m(�(E����1S�c���Wjná��l!��e�+�HYg�v���,�ZfF�u����<�1��9��("��; '��`��N�	� �6�OOA���t3��m�=����ВA�+q�3�6�6Z		y>wVK�K��t 茱�Z�T԰o���W�G��^�,�T�2R|�8��]��d���3o����T��S�V�p�:'Us��#Z���o����1�3q y
p��_i�����鲿<
R񫄑/럦��蝂8�>5p�戏ڮd�E���H�R
'��	��$�O�TL�d�P�Km���n�E���� /����h���/8�p�6�Wpk��#kMI��΁,o.�G�J5D
�=~���_pI��,Z�$/&D��ٞ��F�����<퐬�5&L|�6� ˮw~fQ��`�v�kv[�h����+j}i��4˫%fa�������иzi�ɭ��6Ă3�Bb;et��f�.��=� ���2V+�'�|�����E�7��Ěn���LŪzN vz�$�Q��҉�`c�/܅���Dq����_a��-� ��/VBe��i���'�A�Y��������q�Ï�8����T
�L��CaA�E'јPC�f�8�*W{9�c���+i���4���\r�DOwmz���թ��9r<q��K��9���̝�� �3��k"�!����8q '!K�5W�d��Í�Z9���{x+h�bL�|����9SH���2n��3�uP��F*S�5��;\�xH������l�n�ay���=�c��s���	�m=S����q=��Ħ���/J"����qS��/@ۇз��XQ� z���b����?��'��5��}���Ã��=D�'vVVZ�#�K@Qo���k$�T��d
�\n<���z]|-[�!{]���P�g��7����ivBEԸ]�&�{��\�=���tĩ<{�v���öI��*U��~$ϓ
y*�Hhz��.��zp2_�]Hk)Sr�y�G��a���N{��F	�is 63�p[ ��_x6��;�1�$ϕcfr��g�Z����9��2�S�y�2�t�z
\�\�:`C�(�q5B�!ލ�[��ģl��71���ᅬ��ʎW[,$1Tgڙc;4�?��3����k��e��OGk1�,���;���/Lë�x��RW�D0{+��zK��e|��0�3��J�-p��P���^���`~ϏI<����-TR݀
vO�>���Z�WJ�|��T��m,[V#�ڥ��v�)"b���ޑE��ҿ��M�>?��Uh��V�9�kє8+���u;*0y ><}~*�c���� � �1zq؞o�&���(Q��qEu/ݔ?�;{�S+:��@�Cf��=@�F����e�;"��]��ou��S�LW2!����Y�"�w]��8I�=�\]I5�װ��=\���"kz�r�3�qAjQ
ajW�0!8��5V���}h�5���7X�h��*�X:�tf�i��n/v�`�|���Iѕ:x�H��;B�v���>oj�ٸ�"[qcG��ld��
�*� �&��u����#���H���{ e������^�������G{~>}p��n��kA��T�}+��bR��N7�J�,�&+�|2��(e���:�p ��(���	5e;�t�;��9&�X]�M�h}���:h��k-��tA�x���<�@mR���G��=D
��;zCO�o3)N�Z.��+<�����-�az{[b���zP�"��į���{t���v���^�Rn�ߐ%��P<C�Z�O�@ �x,#�J�܍+����X�{ӏE�9E �f��/7�L<�����w~��S$(�(���~���Iⴼ��L*/,�[37��N1�_����'��^��x�xo�0�׮�?�C_c:ct��,GWX>�@u��{$M�@��uWŤ����o��~T�'���y��G���G���)�Z�������:fzJ�u�t����W��8�ı��(�&�����M����|�n�f{������@�=Dr��1 �N��5DK>�0�?��� c���e���Ř#b����V� ��7��GE0�~|}�4�Ol�AG�1J�\-<1�x{�yG��	jCLA���Ι��E����L)3u���cKV����xo�П��<N,�^�qx���UZu��Gf�D�)*)�ăk�Ls����4����r8)1Ғ�q�)��������p4��v2h�����k!P+�][���nh��8�jY�`�G YCvL����>�\c�BMh�e(��u�~<��kʧ}E�
�2 H�vAa^%����!y��>���s�q�V���}S��X:Iܪ�*����fe�L5������wF��Y۔e���w��6��+o5k�'� fi*�N��wa��9�rAS#*hlʔ#�%�SA
�eC3r���<MG:��lw�n�νlOngu��]���� }P�5��"ݘ�87���:���$�ǘ`��z�kՓ:�V�����n7?����# h����'��Έ�m��&A��d7�2�-�3y7�?IF�Nѣ�l�T�l�j���pl�>|�6y[.�l��騢H��T����P�Ӎ .�M�2i�e�й��r�����օq�����hGd���a/{j!���=VNy���M��`��XV鍏��s��[B�����PpS�b�8��9�I,hn�f&�.����6#;��C�ۼǮ�����2��V��A�������З%I�Ƌ��_
�]��K�Vh���f(�O8˨�m�;製���vz��ċ�\9>����Gč�xAqg��lP�����^�t�"_J�<b�(x�6U0}<�����J�=m�V/+}���,.���!Z3�a��˨}��;rlJ�uJ��r�PѶ�t5�C]KE��e� �T�����K����������Hc��g� (��mty��$�Ϣ|�Y�lϳ&x��6Qx\,�rF��2a8<4���9Ui�>i%�3�#|��p|x�ͫ��;�0��ݺ���Z�kz����S����Mx��D���"���"U��U7C�����:vy�;���u|-������͖Sڢܖf8�q�K��
����f�n�G�g\=�ސ�e����q�Ivy]��s@���K��-�g�C�Xٺ7��,�J,B���I�2��V].P0`�(/{�4D1�[%,�n���R�e��+��1�����Y�.�Q�#��(}Pf9�S�����~�]�x_�`1`��B�)� ��@x1t�!��U��4'�{v����|[{����i� ����v�W��0���X�/E�HXKH����>�t���A[�hZ�
\���a�y�!�_��h�	6�;�ӎk�ˌ��iz���G��/��y�Xe[k�ҕ/Jzs���+�#��m�؝�����~c4�x�������Q���F��id[��#C0F8��+�x�H����^p�x�3:1�4\�,t���b���!|I:���wc��U�[�٬��}Ek�e�����.`�?Q�~I�J�y��=�|���r���P�_%�h+�h����;m@?��>�{���eiAJ9�r�����+)T1�"Yyr,����>�z8c�ȣ9���F_R�`G��2q^�b{�B��X|=S�_�X$,�9�e�~$IVL��:�Ԟ#D��ow�K&��/ٗb^���i#�;\,y�W�R3ltß��ű@�|m1�ƀ?Uj4���!{Z��Gf�x�aRo=����bGZ+�Fk��!���d$V����"AM>��Ev������hV�F�i`1����t���lxA�[��"�9�~��=qd��Jb���s� Cq���ѫƙ����
��w��~?-/Zi�r�����9�cPx�뛨H��iꃵ����~:���_��'��)z$�
����̄$/�U�lbx��j6$��oV�%��K�����@�^c9.!&9����Q��������4�`�$N�F(��D]�^��@��j�	ą��7F��ܜ�
�]�����#
!�`�;y�x&��C�4�?�ڌ����6�k���9}ǕNz�	xw8�(i���X� �]�ŵ���FP�ߡ+'��A����ηTV��3�4o�f��pQz�t��'�D�4�C��U��v8�$a�y91<����������lE�Rq��=��|�#�S�~�B�u����2��9ٷ�E ?P�K�<�䴸�=�/�"�:���^��9~��9C^��0�k��'�'S��ՔS����^��S�c��xQ�\�3Wq) vq{.AV(3��	��	��w�N���`bJ+f���������>�ϭĭ�Mx�C*<�U��������b�}>&��a��#��S\ܺ|�@!lųv+J+B�9�XjR��^G�y�g���ݔw�!�%����y�2؂�u�z�����#F�ﭓ�=�ce=q�]kX�Q@N��t�l�#+�b5�(�g��:{9�,�m��N:r	�la�l�^V-rku�`d��x���SG Ev�3>�`i8W�q ��W�{�u.����:a��]������Ů��Cb�P!��3	�� �R�zs�)�PMnb��w'_��!e;�վh6����EeϺ[��磢-VLꞭA�i�FT�P�W1�����C같�n>#����k�"�p��%�0n
�<3�\RXܛ��䖪>�)�?L�Ƙ��ӝ+Ћ�<��Z�a��s'�?�as,�Dz6�9����C�*������L��\Wپ䀔�	ݕZ��-{�?_I� /ۙ(�(x՝��%k��X�q0_r�lw�3�B�+�WJ���U	iֵ���G���X����*<�ev�7���m�E�5�RVWN"VZ-A6<&�+Q�����8�ӆi��u��åZ7��f�����VK�%-�O�_ء�Y������eYZx�FatΪx�J�-H�߅��Lnz/��S'R��i�A4�����!_�(ה5��MG� ������
B�HʘȄ�y�S���o��Vd��ƪ��O��4��`S��l�!fM��3��|�^����	R� Gڭ�)LӳN��/�(�ڕ��ᤸO_�4	�S��ȯm=�1��6r�� 5_��f���_�@qo]p�	d�ঽc.\������V jzLD2��*"���t[5��e���	{w" �҇`�NU+���uH��Q�2yG�?����V�r���"%J�;�lz�+�R�-�{y�갣�*|��7�h����Z�4��� ����+8ꮇ�����o�(���h��c�Kl���m]�ef�҇ �21a��S�v�+,�q�m��������Zh�9���:�}�>ῧo�ݑ�N)ls{���q�+��K����0����v����$) �IpJ�Oj~a8�]��|)��~[�]H������O��]��I���j+��]p�Sk�s^m<	pȬ �˖zx���x�Ra�[��:�l��=�˯Y�\��r��I�y�b� ����/����!�QK2|���efr��> )���GqMwx������~���?n~
7��J����=�I�FH��aGJ	��������=�>����t�MD�J��Z���K�(i�����Y�@��g�Bd�����L��Rp�x$"/�L�?X����t��Z-��*k� ړ��/>�x��QdS�N�Q� ،�O2v��EM�K�IV�Lw@b��(�)W?�/Q��R5fYGN��HW^�TC���t�/��3�څ����o���Y7�M�n�&�q�k�Q�-һ��ϱɜsHD���܁	�絝`�G��R���'c�u��!9����ڄ�/���j�K}�X��}�g9���wV�"����e�����ͻ�A�E��x$��п�0H"?Ey�S��i|z���7P8�g��;w^j�Hڒ��z��UA~��Ĳ��G�)�7����(TX��c��1�8m �:W*o�	�ݱ��lo�-�(����e+�8��\���;Ki܉�@�_D�[��(�냕(ֺ4$�C�;�`�)�L����	r��3��h,�y�2�����Q�TZFK;1��_q���*������kc�.���|뀢�l��#���H�5�*���\�Ʉ��66��d��{0�EbU����� 1�r���������n�����	=}^o���Q_a{ H;���u  6��j��g�]�hn:$����Ed��C*"Pz@�[QnoM��.]Ojq��T�&�3��.�5� iX�»�-(V�1pNB��~�L�{/��L������<0(�����d̗8��#�w�o�ˎ4'^���0,�	"9���3|���N�9X��z��ݛ�,��<[�y�,e	���F^�	hG�f�7�<�i�Ph���1��F��%:�wxe�v����$l1��H.�omF.����Twi��:0vMe�ck����S��˧�����uU)�s��wP�Î�j��ѶP�b�o9cpj�_�����ۥ�[�7���!Oޤ�r�=ȊyrnE�kC�$����q���Y8��唐 ��i��am��N�s���# Mt���9������^���qA�j5�>�[i9p_Ac�zL4��oY5���b����<����4��x����z.2xwzJe�n�zKVӥ�,���^z݇��*�\t����|'=�xڵL�sң�^�l�}Na���6��Y7�	�N�`@4Ϛ���\�R�eS�x�d.~���r��U������Q��E9��-�1�������b��~q�Y�O�۞�4Zs�z:Jz!HL:��y�0�������y�i3�!�R�^�r�T����SJ�wF(߬�o[4��]�߶zV���,o۫��������������� �{R�9|l!���0����d0��b01!:΀d��ʘj#.��[(X���>�
�*�S;0���<������0���͐ꕥ�A3��d�i�48��G����:�q�|�UUɾ��1�J1|���m�s.�w�eK���&�z`�:'ы��4R ����eƜdC�������U�}��ɹ"�lm ���ٴ5�d���-A��Z�#�K�He�id�k���.ld{S4%��	WIX7nDWq�3���o1R��A8��-Ȍ��x�||�(a�W׶�����|�j�Y@��گ���]wyy{P�f�rz��E<�C�7R�J�Y��Ė`���
9沖��8JKD����
`�?�d}H�z�.dA�7�q(dW20�D��^�>nRݡ.���#��P؛2��_�>�I��B����HO���yw�v��@y����w��� ��O!�_sbz=Ax�����,��|d���;��s���|a�C����*�	�����]�-Ա����[$��o7�6�S��2��gU��A�X�e>Y��X�"�
���Ȼ8ZbEn1�z"�-^�7���A��v\�Ģ8�[�G��O�S�/5�Uפ���f�̦�%\�D�NK3q�~��D.�i�w���;�o@<�%�!K�z�2լ!����8
���Zs��^
�؀�/������L�姻DF#-��ϼs×�}J$��+fm�+�h����v���u�RY��^3�Jd3�^B��f�5�t��҈��M]��\&=����g�krfMa*�F|D����lL�Jj��`��a�Ii��	6��E�����͆�v,�!�P�ǹbQ�׆��"�+�&���տ~_!��Z��	� �%��/��@�B�VαFp�_f}݆��;=�P��!�P�A������k6d�S�_��h�|�I'f�}�I��L#�~P���ϲӾ�S�XN�7c��$E3v��OlEg5����4���i�S�1ÌI�n�yW�n�#ʪ٥��U 	�K���Bw�sa`�����V+�&��IA� sz:ww��±�c��Y�v!z/���m����m����^��.䒰\�bXeԢ���w�8,,w����D���4��ȜWX��(cN���}��Ȏ��ҥU.m��zN�^*�d̟+z��y��ы����vx�W���ʒck��P}��{����<�����i�9_S8���%�R��fC��:��GBrEY�����^\WU�n�z��/��:g��->��'
�:F����� �F��l�u;�����&��m�*!2�Z�Y�ӼZ�vA~�ـ�8�����E�_��"D�E�$1�"�Xh۬��K��Vn|Ǣ�>#���ؾ[	���ri�����F�� F�e��,�����s�zs}b*�fIg@���.�*a��s����a���)���;t4aȀ*�>�k�h���IwЪng����H�,�?Vf�0��!Uz�
b'�������S�4d0�
�N�P (���lUIq*�ޫ2�O3e1R0A�;��;ggu�9����C�\� �.M�:B��,�y��������eR��0
�Pf�������s3�!�;t�]�o�PQ��*xd� �x��ʘ��V��[ٜ9�:�}�~��ѻ'��`q�ܫJ���F�|���y�����߿��K�3e�I,·u�D�]�,�eJ�(�a��'v�p0��qpqs:X��a2&%�x?�̖������ܺ��J�ݖ�L-.� *���E�3BѮ[��@��)�z��Z�5AO���7��d.R3��J_�X�Sc��FI?��u���n�ܔe3~�O��,{v�"��~�����\�se�\z�
��x���C�`����K��צ5G�'�k�A��w�8�|�3bg�='��bJ3���B]i�踟V8��Z�F�;�s�-03˶�����ۢ�XvB��s��$3O[K�+�^4���r�����N�/��L����X[A�_��*(��e�K>Ey��R\}6w+�9��8���Ԗ�mm�������9���I�^8�����T"�����0aB�o�Q��;�L��M�Ӛ�o�.��F���O �A;q*�Dm{]���刋��eU_��^	�R3��V�ƴ���Ft}�-��^��ɠZ�?�����&�9�ԁq�@�Yn$O��'��O�0W`�ر�h�w.�d��[�D����k��Cv��H�fз^I�/�sE���߿阽TȎ�!�2I>q�f�|wiJ �ٙ��{Q1\%�W*D�ƙ��NA��٬4nH���Z���Ol�8<k�������?9�����X��SP]��?mq������]��?a[zeA��y�*��+�E���a��؆����"�!��wWIB����Y��5�����L�d�3���!t�=�h2�	�Ϗ�9DPh���P�?���:���8�	���/��X�u�.�`�:msW�,N*LPfؼŇTp|3���х�ˏ�j+�ӳ�3���܉���)Mc$�����yԉ��x,�o��Pcp�{Tw���4�#xV��S2Wg����V�FB�[	�r_��QF^�{�S�ϧ�2:!J�W�5��{�����b[�/��m�ɱ����װ��M�L6����ȌX2��L͵_�^����3~!}+:&W<�����^��	�8�e����~1�*�( ϗ00�YB/��bC�A;�?� �V���Q<�����ս��!ObdE&�������o�eY�+���x���C=[:��W~����կ#���V,gYL�LMe����7�T$9�jA��^������.��2\��Y�Y���4�g��]��?���ԕ��7���x�sEF��+��Ҹ��*�C=G.�I\��y�����*�����K�v�$����ʼ��p1#>(x�>7�&��e�/S�v/aӹޔ<�[7�X�E���д�����Xz<����O�?4[c��w#�y�JHt%��¹�R�u�Rl}�Nl�D�RW�W����\O��g�L�C0n�K��$����23�n�R�vj��f�q�蝫�.+���W�?O4�$S?�1�)XCv�<��	v	��íc�9N��q�Ш����Q
w��jҙp�4������G�]����k4�h`��Vr�ł�bt��ѣi�(A�NvCsZ�j|6�{M���� ����#&���c����ؔv�|��:if����GY̥��ߊ/�^,0��������h�4����E��"��y���#R"g�6Cd`�����m�$ų���[Ӳ�� �	kmڍ/����5uq[��+�o#a+"(8��</�H	�ч��R1� C��dK�<�gU��w�G@_N�����?&c��L�@�b��a'u&��zΌ,[���%L#��>��3с"�0��DO��qa��)�׿����E�z�qKjf��TP��@���Zl��ZL���@��l� ���c�������J�J9=����^�P�|*�Y����q�[�b�)Y}&�WD*0yKay�Kj<��w�L���ku^���8��t5�V�r�% ��l��#Jnls��W���t�3%�Z.k�@��5���N��N
�I�W���k��$�B�8��OJ䖀yƘC��`d;��xl��(<y���'ëf�����b�4���d".x_<ͮR$��5_ei1v�Xi�%�1ѷ!Z^#l�$U�w�0�	/ ��met���¢D��$ZwLi�o	d_w�ؖ��Xҿ�㪪�=���Pv�( t�4�_t��n�$Kh��y��	����݈� (���0�PKFuT�ϯ�g�����|ț�o��r���
B�,b���g=�;�̜GUK ����
K�p��a����~	G�76��������3b���#@����C�1[չ9�gJi�Ӑ!
d��B�
_�7�kI���-�.��9V9� �̫�q�T�hH�oe�J�:�xw��l܌`�~��;�H�C���ÒB������tM_Y��Jy�=(`��u�	1�)�6S����Gi04^I��q卿͗>1;}��ȕԥ:���m�`�v��&^eSf���p���|���Ju��k% ^cY/f�c�{������^����JD��]"��o�/~�}�~�6'{=�{�8��l�F�0�
��!};�7	%�-��p���IhY������e0OXR��/C��_#��t�~�ڑ��Sf�jRFQ���tp>z�iE��=�Y3�����WK��d�čά�.uN�*����)\��ȭ��Bf�)�Ā��r[/�
�������ᷙ�n�d�0m�t��Q�9��;D��:@��Zʭ��FS�7���$ �4�eVh����/���f�EQ~�-H:�^'꒭�a���}�*Rg˷��X�xdӭ�d�C��d֌UՑh�}��Ѧyb�D񼯮��y{��_��wc�4�Z�Fl�I��_76*p�ֆ?��I���{�6i
I�,=�< �z�,c�g�(��_���P�?�#�����z�������iI%G8�o�a&ͪ����@N9�.������K�� ��\���z�q�L���Ú�r����a�"��t���I>�LS���Z-:b��/��nq�4�C�j�M�EL���X>~�:f���@ȣ)��IY�K8�(��el�{􁭷r�.�y���˳�/�Ue�ڨ����!w��Z�f��a4��t�����
������ڹI.5���[7Kr�d������L�;����?��Nv��&��p|��FC`m.��K��ʄ���:[�;v�w��TJEO%};�1ϼ�J�O��m�q}�F]��o��h�=��(��7(����{N�`��H�SҺ��('���F����y�Gɐ��]��J2� ��݄]��R�������	NF���z(?�]*�ŉ6`�{��ӁH���8>
���4vRJ�( ��_z(���n�FVу���O����Rև�0�v�4,�B����e���<�y7�I��;h
�/}"�}�����X���n��m�66�'��PG�=�#W�(gE�˼qė��Y��۱��J#�Y]H�4�	-��CUf��[O��12[夤h��~�j}+(��ʣU�Gr��r���ȗV%+��H�pR�@n�C� ��3Heh
{p�O�B��[x�NX�ڛ�������Ӊ/�S1����6d�Ӑ�ԫ�j�x�_��X�-���="��a�XEa˵Mv��'b�Q�л�ԋ�岓�2��C����[��.P>x�L:H�ċ�v�@fCO�����H��:�^㼟��|F��(~r�*��t΍��9]����qֱ��݃w�"��#��U�$4���q��'t��謠s�C��a1e4_+��b����w�a@���(5���Z� �%>�$Z�:�#iU���T����z�"����K�.e��Xgݩ�x�A��BH����d�Rǽ%�)Տ���D#Tg���q�`r(*�|&P�M^�<��S�w ��0�+��2 ũ��ਧ���> ��	�_��:�<���I��U����P��D�7� �z�������4��a0�!�~c����;�A&.�����EN�N;Ί^��6�~�|���|xP����E�C{��ǚ�������M�q~�[e|� ̮��B,�rfqF�&�5�	ޞ����M&֌���9��H8���~����`b��b�g���d8�i�>�c�$gZ��
i��|:H���G��Gw2r�N��J��2rf�4�m�������A���5E	}h�h��0�����<M]ܱnc;��[�ąxZDN��J��R�����h�ܨ�����튇Z�oG �m�,����s��0�U;�j������~�o����'���e'u�>����n�"�O2�p�kQ�����shq����s��3	<�q3����4$D�`����R�
�qO�Ͼ�'�e�t+�����o^�����-�(���[m+%���V[>�}b"#�Ć���G�d�h�nM�*SYg�"�v7ֈ)���_X����[�������8��hn%��S����AȤhY.°�P٦l�I��u�'::���J�7��r����鸔o����q����k{�g��&�!)���R������C2�X�z�mpq�b�d+�7������i�>n���aO�@�B��)Y������.�!�x���:v`�ð���S /Xx�)A�e�UXV���D�ġ0�`�IS��A����+�:���9t�2�|7����X��ڊp;�mf�t��0ۚ�?>
�-�@��zM��d{��:S1�R��ȍ	xSC����U�=�7�bC�V���P��PT�v]n�-vSe�H_ZgG(��?&�%{���7~��<M��a�E���]�g�~D�;�k����k� c��*��nU͚��EZa���ڷ���K�!��G:�B~~b�~�;1�@�q�LbF'�R��l�;��S�g��$aS�Ԑ���
A���{��<hć��Y�����=�Ǟ8g�A�,cp�/X��i��yc ﹑��Fs�AKa�x�JE{�x An#}Qƶ&ϢP�L���5��Ha@�'�z���񦷆s��k�\�[�7&��^������������t�(z'�&#�NW2s���A���	���x�oH%�˶�-S��M��RH��o�G��
K������^��~᜹N��Q��-,����AVI�+s%^��B�G�C����b�BW͑S�iCoN<d���;���Z�#��<2+Է%7o���ٍ�����*�X��Z.�3$��<�H�Zx.�hd�׫��"�\b㪘�@�#����+� \풶d���Y��sDڴ$��u+�x*�� F��;|鍙�y�em�W`�T�����F���$q9{�"�5��]�|�<�+�|����@􉉓���QtW	����|WQ�S]��:K�s�۔[�5��C�����Ɋv/f�qAaS�W�T���T$Ur�f�n�B.`�k�
�'��C��ul�_Y:�v�`P�^�X/��4�� �w]&����6�=����Tx^$�C��S[_���>f�{C��*���P ��\��d;�q�ɨu����J�
��͏g�C��B�C��g�b���4��4/�H���+R7o�Y�2"���2�q���������0��F�X�@`�-�����")uz���U@�R0
����7�I\���x9z�HLH�L��L{O1�.aʏ4 ����ۑ]�J�M��A�,0{$q7hA�����v�'*6������
�|��P�5Z�x�j�B�(�`z�c�脆o$qb��bŒE�?�L�b�d�m��J������5����]�]��1F���弖Ũ�vh^mŢ @�gxY:�g�:*�!B�w�tv4�%�a�F1��Ոt#��B;I���÷@���}9���&!��ڽcJZ�*/�R� ���5��KB4�><&�ZG��(؏����\��;�m�r'��d}�e!ia�w�&�]��D ��h�}#���:uj��X�@��>A�ַڸ�\0��N����������k��e#�Tg�B�x����0W#BI�-�ކ���2	�,o^�V�l8c�ϱ�PE4y��������v���S޼6��8�EC���f������_�]�W3��7��h�gʶ�JK2�	��M�y�J���7��h�.���n���
���a�%l�ɂ:ňX���m���x�o������2��3��R_b^6�����h{������Y?PZa8�k�	��I)�Y��wp�Z@�ټά@�B5�n���(�:6�2����<F�<��d�(kY%$��2�l��7�ՙ�İ$bҕn�Ϲ�|���!}+3���	�����z�aj��~�OK{z,��/EW
��$���?�0 ́��Fw�?3�A#��;����������.h�I������W��%�x�} j�Rd��5�
Q?V����f��V'��u~J�վw��8(�E'l��CNף�W(�&���+Z\,�Q����mr�Jq��uGV��O���K�W���'6�CH�#ɍ���#�a^cσ��=����e����|H��r�+xŚ�k;-|x�ϻC..7�1�E�j~������b�#�&"LG���M!ΰ��P86OG,��mj4_LT���V������G�{_%2�NF;��.�|�M/�8�kn.Y(��G�0��<��Ege��Ny�M��g�}¹�z��x�O�����#�f��]
�pᰚCO��K��z}tk����;�]���ƣ�/���ܡ��	�uWc�	J�#�4x����E��$]QIf�;��O�0�R_p�nk#�ԗ@5$��q�����g�>Mu��<V�+<|�\X֎�*�0?�#�͒�>��[fo�JI�`�	�=S���Ip��_����Q����%��Z�4���c[��v �N�V4�U>�׹-dY�I�����<G���rO��G�j�%���ш���tQ�m<�/��K���Xv��k���E���~�D^�b�u@���2f�������Ft��N��n�d��~��B�:�?��j��<"N.������������x�u�.��k�Ұ�k�sj���ƏQ�%QC8�i��C�R��ض3�5ݢ.Xi.=_m+�h��_��$o,:�`i�҆�^yaI{�(i��B���0%�1��t(u��)t��lN\�����D=�����1�#V�����SX[�-,7'�J��(]oa{b��3������&L���|t�oC�I�����e��Y4���cb~�jL����#�\�
��H�}*�F��p.ARK+VMbNAV(D7�<.}%=a�t�]ꈇ�H��ь==��ܰ_�.�'7Kj>��|�.9���;�^d��������� z���(��nu5jqG���B%I���hd�~���?�xk�٤<|Vh4S|� 9��ޣ����@��}�S�M��d�$X�fI{���6��.�^8,����ߢb��&J�e���q�@kx>����f�	�j�`D��}�o�+�@�<�Q�!ٱ�#�Y�Zݮ�.~#A\�bȅ��닑��w֔E��?T���&���`Kb\��g|�u��JőՒ�t=�e6�g �:�+.sU�"�_�Am��7�}M�y���㐷�����ńdL2vS�\�QK5����^k��# R�^�*���s8�TV7LC�I��D�u�)孃������:<[���2�2%`��n�����J1�O�O�,s�T"2�����v�v�LI`����Xv��I�ν�q�D݋���m����d+��!ˁ�1X�>X1��'���݀Sv`�:��Q܆BM�g�ޅ���3�_�@�;��@��Td0�������uڥ��z���N����w�3$���u̧���L��Z����(ˬ�����=[ܒ<��s��t������2*���q�������:��
���V�<��~��G���:�ڇ|�zb�x���Θ��|:��Տ�P��C��+g� :�ypX};�����͜j��o�p��X�嬾��|y��x�R�ҍOO-⸷��g��l�u
�8�������n�ڎ���c�\Dc�'ӆ��i��&�^�gq�R��*u����w'Cn�J&^.V 3�Rx��'�]��:)މ��,��K"Y������h@ҸȤ��)l��M�:W`���f�n9	�C���E�łѸkϫ%�$^��XF�^�4�ݵ�nz�����`�t1�($��[�QP+M�Ih]S��<��w�m��N��p����D"�B��N�ퟋ=4��a��f��sҰ�'W����Y#��.���t�Rؔ�z�v�{�.J�Q��U�D%I`�~f����핡���@�K�ѹa7�*���DÝ��-�r�*����Ν��`H��͌�� �s&ds��������@�,����fD�({U�:b�탙uf�;�݄�Rq>Fn�/�@�ӱ2��S2�byh����o�;�P޳(�iPl�
�����4��闬ɓE�!�I�bv]8���e�W�Q/�'E�:3҈�20�&^�,�l�_i�A	�*�?�L�6����]fI]����)R��O� U�m�0?R��y�K����g�2Aލ�)wn�,��L������1:����T@���p�#<�"��:8���A�e�<�}?��u�k�6DO0a����0�v������X���}A�E����AuS�p	���?Gy�+u��ϑ=GcF�t��%���T�}L�.�堋�6�^z#�S>���_����>k�Q"��W���p�T��"M���MֺG*��h�GJ�B@t���	�۫�Lp��Kg�j��b_���S��=��E��}M�5���I�k���|����elY���W�tQ�U�	SM"�CYP���,#��Y�fq@�V�Y1��.���:�H�V>��"4Ct�gf�����}��<�����Tt]�̇ĖSF����?9�~ӣ�Ԇ�29=��.}I����~g<����"6�'�pF��E^� ^���R��+yż�0��]�����ݬ��ز9#�#��cz������Cd�V��H%D��D-��s6i���<P�y?��:�˱���N|�����Ew��5#U�'�����7�:���`��8�������F����C8�^�`i��Ԯ������q��,$��&h�R�3�p�n`7��I��z�Ɍ���9�x�&EY��Ow�ܪ0N��gl���˸6r���bEmA���g`�̧�`]�|�U��S�4}��֓L�9<E�Vs- �;;�L;}��"ȄU/֔���wT�`�\�H�Y�m��z�ٕnV���
�Z�w�Zi|꺁� -�Ғ u,�!�N�u�
@��]���P�{��ƽmۑ�������P��0��é>���tF���bh~�k)4x��@V1Zv�Ϥ9�)�+���o���AfVs%-����+(JR^�����7��<��"\2{n z'7�$�٫�B\4�|�CV�t� Q�?� �P̓�	��7�g�B*��\����巕�'O�r�f����z�ˬ���}o�<���}8�[��9��*G���F�˟�����7 
�x>y'��	�����'\cqB� S�`����򫾟>��]�!�G4=F�J�\�IT�_�Z�&��[�ѻkwj9�}ao�����v �0���A��q����~�H��͓�����s���&�0�<�V��`�s}�������S�����B䨼���9&r�S��a����/l�On���X}��?��Jʴ$�!��c�������Z�B� �R����'����-b�\⟎���]q89	z�}ԩ_�iǚ��q?���S��R��iT�찏85b����C]���P~o�K�)B\nx�k�U1�Ʈ�[,�sL�cV~��xXJq��k=��C�$sa&\��Ft���(%+�d�{�j��ȏ+p�z+�{gP������$��wcJ�cd� ��%�Dz�{��[��I��OvH�4��w��'��׉=E�<�qH����0�h�]�g\�r��@!�lJxk$�m���7���ky�� ۵WR�t���HG��ኢ�?/�mH|�}�w�D7�z6�M�2�DE���I�^Y�سiÍQ�V��V�X(��@&6n)Ť{H�6��@z|�	��`Zf7�=rVTl�+����l�p��֮ gU)�!���w���hS�0nRC�t��Ի܎L�����:��C_��5�GQ17�<����$4��t:P����;y#�4x@��u���C��7/;Sq��Z�~|��ļ|h���r�xTI�������1�A��_��U��W�a g�vQ��2�����+���7��.4��| �w�<���:i�@e�V�)��iRN;�����_ܶ�:i.������n��M\������x�oS�h+�x��-��=h�q�c���iƽ_�cK�vUB�9���e�����_,����k��3�����#�(����O�o�l�z(T� ��Ц	�G�� 5�2]��+��F�������'@��`pc�:�9v|���Ng������'�1S�v�{B��%���ݍ�g���0�hk��I�������L��I�T*�������?2��_8i����+�����Ǘ;c��������[~*��s4NZ��sN�3h
�?�O@��縿��)b��K�j ʳz��q�#x�	��g���r�Q�$�� ��I��Ԫ�;5u���2��i���6���
��3U�D��]�N�#�
���`�c�#![����M�$��3/M�	��P��	�&~�MK��2�O�N��&������"��:Y�s2�
Z��Ʊ��D����L�������恨R:2i��7�����/$#�
�)d���A ��n�/vI���}�!�;�2�X���}��'�s��`�	���#^����Ji�Q��Ȩ��\�L��	{����~��%�����%iiǰ���NT�W�COS�Q��"1�g�쫵�����d��E����.��FGv���#L0'%��3z���Vj���fI��L���\X���:�b�.I��l�.�~�z�ݝ3�b";�kf��w'޾�}(�P��2�@�n;��G�ǿ[tF�f���0�9$��f1�r�"�a�K_TS7�6`AA*�4��T��ty>@1�3�v�8����[R���lQ��'�u�됧s�/	r`ip3�{�7c%���W�p͔���X�i�[��u�i~DV�2���|��*?�Y B��ˬ����8����K+��}����eՔ'������\�r~�^��ٯ�U�(�Tv=�����
��5n��w� J����-=���Z��Ok"��9"|1���������+2��� l����e6�=������}<:���<j:&�$��ddw�i�f�h��/�^�_�oL.=q��K��<�W���}�%#�ٲ��޻ѐ%Gk�=��)���,T�K
N�Cx��q��.��d��4$���K_����.)��H����]И�,�{���	'�=5��
QW�@�Y%�#e����pO�R���&}�g%�Z�4}C�ʊ+q{4(�t�9Ip � �k �K�!(�e�Bp��s}�g�T,�M�s��[�Kc��~�v�К5�vn�����  �+�X�S2�,*ǁ��	F?�s�XX+����rL��"SS����p�*�GT;z���9C�4FUw�#&#�<^�2|���%=�ߕ��J��(F��(����x���8��2��A�)ܟE�d�!G�4[��n�N�D�.��Xrw	��rq�8�1�G�`��������p�>Lv��B:.��8�ym;q	'������L��P��:kP�Q<`�Y�ؾ�b%����6��2�Y��F�t����P�T	~�d�.��H+�!R�	ބ�Nb\B�$�¶L��R��l������Pނ�}M�<�<�ǭ��B� �*�nۿ��14"�;'rJ���?h�^3̡�Ƒ$�16|Ж���+�2`����P!����p{c��sE�G�p�"��D�q�jqe��fW��F�g2���X���#���K)�ǋ�~����������d�0Bg���d��dݍt_#��)W�RżYT�̈��~�M�@�=I��\õrW��E��_��'���#K�im���k�hKa�IsBb��<���]_d#��R��d�׻):�q@�|�	Af=e�m-���(�:�@�����vo��D@�����3�j�Yten�4�V�2���������-<�iX���l�-��܈!W}��64s�ꖗy�D���8+�n���5��m���y�̹}���[^י��=�Ξ��� ��8@fܧ�,��C#�~N�Z�t)a}]|s�a��6:,m��T�1�C&����7]���8������P���Io@���ƿ�輰@�c�5/my�;�>�.q�i.29B�Ly׾%^��Ŵ(���7;���^J����%[��DY�C"F�F/02�E~����J�	�� �O&?�ѷ���y�C��i��yf�1��-�mb���/�3v_SZ�{[��vf��S�"�3������7C5�T�.�e��B뱙��{x��2���6�f%/]A�`-)�1��<Q�L{�����6�@�g���7��:~�Q�E����0Z��t��+�$�s���^���,�����dp}���Y��8n`�o^�Vc��I~�K�$����Ȉ%�,4��V9�s����u������t��nMH_^�Ӗ6xWIðj�v�vq÷M����������ð��X�"Q�����M��'|��yf��ZO�2��B�o�Zrvo�K'�������9�	��pP�V���5>�����6:��x�Jf�V:��D g0� �ٝ���[[�(�N�@Ի*��6i�*o�:}?�������M�w#YD� ������׳5�<�)�\�0��K��<���)�Ȉ�8�Aś6�@�B��*���/�9�W�H+�î���ކC��Iy"�e6�_��<�.�~��E-�o��;�#J�X�2Nз;�u��F�6��C,���R۴]C]�����Lu�(�s9���<�"�v�29/�'ivi��E���f���%�v%^������͍�����y;�&��uX1B�s�4V����6�6V����ĄY�H�pgH/CR�n]��JaN3�l��6�q�FJ�/��-F�"�=���26��ͺ2w5�[JW�Ӄ����	������A<PQJ���=�p�V��^_�N���S,�/�Q.�eSZ�A;_}S�+�������j��O����2�X��5`�G�bm �# �wI(߄(q�hT+$�b���.	K�*SM��g�9��]�?�;��z|��I�\yK�mPI++�՜d�X_���8ʆ�m�ΗP`.{�p�Ζͣ}��Ґ\$~�D��*ۄ�;g�}�=P[ڽ�N��/�P��ԲI���!�z��ϓ��,������U�2�~P;䬿́}U�/�cin���+ܷ���A]�%إ2vT�R�@��y�gK���@q�*��Mt�Y���&�sYO��`��{��n3���[�W���)����^=s�Շ�����3��[��ߊ�7F�!�В}$v����~���E��\$���i�&�G�ٶa�����keT�΃,�S�^^��ɠe����N�I�A�:N:L��ω̵�w�D�P)�z<���P�A����ڥ[ɚ�_�5re�n�*�";�K�re8:�̓S�A�T]���ם��}?���5���+���x�2���0�S��>����3��Eo�=p�vv��-n)���9���!7"�O�+NS���#j(w?e3�A��}~��J�f�����C��Y͍"��]��޵̔xڸ���X�AJ���S�Tyk)M�ǿ��f�)u�=.�q������lFF?P�#��7���Rx�>-�)�pN0���
�C43���gh�#o%�S��r�����I-������t��r��>�+'���_��)��\�o��0��mCE �"��(3)s�]�^�kM�{ �X����m�iY{���b"5.ڛ��E���Ѝ������Ѿ��b�D��4^��r�؅G��C����,���>�ot��[Ҫ�=��ZK.���U�~|j�_�	8��n��ۻ/B���z*="}��O8c�Ω��\���/���P�h�#�K֜@��t5��(�I+����+�r�/z�2�^�� ��#��<��7^� a���{v�{����Aגy������(�O�l�}Q�5�Ⱥ�#*e+U1��E�dW���V;��k|%�7������F+�,]�IO0U�ߖR�����{.�y��Ozb�+.�wa�wK\u�����v���nW�&�E�H�����Ok�ICe �5o*�	y5̀&`Ǡ88A��z�j���~��v7M�L���~�O��}b�������	0�¦�D=.�L�܌�l�nt��fm�ʗsY'E���ԟGA�'�)�2%3O�c��/����'0z[�6۔_���y߳���$i2w�,u�	��p�/L�Ӳ���~wOe���1���(9a3J��iAߠ�@D ��a�G҈u8r{��4��/J� %�ƥi��>`�����j:��w=V�J;t�D��ciڋ��z����C�ڬk��	���nY�#�k��U��d�%� t��wts&[Nw�t�?L����ob{�߈�E�9��t�b�+PI���\���KICkצּ-vks������@�Vש��eo%�_-O�2����x��ć����\u�M�Y�9��.��f�U`<��C�-�*�=2���6����?	���ɯ,�l��{�4�a���A�t6X
N��C�9��@�|��;.S(;�w�1�ާ�����Tr�cV���	�<3QA��L��^#�.��֧V��@#�,z��􎍞�P,]5q�g���~Y���ϼ��r�.e�rbʓa�%���0}���{q�83<4�(��sH���j����c�钽��t��b$�ʘ���i9);S*y[�N��1�m���
��K��T5wj-��S�HE��Q^a��ӟ��>������P���o��'q���Z�n�R���d4�{�R�39��ڈ�,V��,��&��AhK�`��؎!W��k�������W�I���>�_��B��3�1��)�@p�|�nQ�����!�@�cvXx�]�P8N㳠�<D��9�=�޿�K���i��d���-���lpt� �:�I�2�T7?i�^z��c��$��f��犾G�/�~�#aO��a-LB�y�4��1BRn�g�ـ"f;��������Y�ǌ�������hd���Cė�G�]_��N�&��q��M�H����~�����5.�.��`/���v�:<�r��{. ���I+�~�Q�q�W���w\wn1Dr^v$XgN<d��U��C���Tj�Rw��9	*ő������Q�7��Y2?^|��)�F������WQ�>���6��/�ElH���o��{��z �0c[^e�?qd����z�D#o�&$�G�� <�x\�a�=S40X-!�����^!K	Z~�I�Q	JƉ�U�vM38m!�Q0�@G���-0cmN�)5w�ic��O��.��K��, ��8x���l7M'�w?�2��y�r�I`ݹ�t�W)���C2��_���*�Ƙ�L��/P�FZ��@}�z~>/~�yRnO�0��$�ڲ�����x��b����@H�J�\�<�O�pȃ�y�!N�*�lqp:[�-Q`ģaS�O����4Q���7�M�l'�_H\l>�}�$�,��k�'�
��w�*[���D�_��O��4�V#9ieȒy��q��'��G�ካn��d�I�@�`?J�"�.��ԸD�eVGO�#'%�G+dH2�%��6o�I}����Йd����u�]!��I��r��Y('ɻ���I_%��Xˑ�(p_�I���yӽ��G�]]G��gԒ
�UP� r�Ԡ'on���0@@Xt�V�jtic�t_�(�!2�83T�ό��c}����el�f;e�Z�s5/�M�Oo�I'3���}���*�ʿ��H���8j�\U')���9��B,�i��PV��8���(��t}�����k��r�g�b�W���
R=Ӏ���Q����X���d���%�|!�o!+b�ȶ��.�V�6x���t�u[^2�R{kAx&��Eab�y"�@`��i]/c�mb�!��I7�yE�`�*���7��a/�1���1H��v�o=_uǓb;����c%��z��!��F.��h�:����"}\��p�C��J-�x4>�V�AtW���v�f���O���)�G���TQ��G	�F�9�6�'������ܺihu(
i4��}�[�ڬ^�Iq�^�ަ���v��g�����7�1����ė�+���-�6�p,�G�ȒJ�T�������S�A��ۆ��U���[��T� ]Z�ĕ���H�S{&�.]l�5�"E�l��
FH>B�]���������"������7�
wOSg�bE��1���w���CEFY�T�v\f���"ȧ�����UK�d���1�jC��l��7�d��з�ٞ�B��B����.�jc��R.��>�X�ˏzq��}@�!�,G��E"+�A��P��r{�Y����k�y��*ï?�	(
����3�f��$9	���f�
�p�.�~��bL�-9���*p�4N;���@]��K
��BI���}�|!��-V���J�i�!����}�t� ��,j�%��E�������:�n<��G�W���I:M�d���|�4ڰ���|�	�K�#�9��Z9���jm�xՈ�S�a\mmɅ�Pf)��4��@��:#�i8;�.ѵ'v-��-�}�?N1�:2S�I�D�#2c�Vx9?�B)W�w��4,�p�2i,g|!�����av6u`��LCV[�A
1���7e���-a�A�E~��F���Y���& >��]�1�3A�A�K��x4�S��k�FX+�}l�gE�IqTI��I�:��*�}|D�I϶k5��i �[.U���/v%m(;�M/���)=z�䄲����Np���m?�f�O��7��o�ӫ�e���n�G�})_L21�������(6������a�iI+j���<�o5ͪR=>��>�{�,�8��1��5_����ͺ^}FiY����x�7�1��U�ۋ��%*�m	��c��b=�Q=��$�W�ND����Pbw�y\���*������U>���+N�^�Q!�N�	��0��1[+�O�lB��+:Y�����,�ځ��Ne>�d���ߘ���V_7�R��&���zt��.Ҕ�Ŀ�}|�&Yl�7�NH$~���KRi18��NRuz{��4���^��g�3����KL���^"��Ds���:�&��佗9IHl��K����=�����|wKj��A*/�,�d���/	]��T������eg����5냰83ᓖE���\��H����T�Z-�`3�B*oTj͊Ty����qd��l	��f��������w�,`q�:d|򲛕��#")���)X���??��+*}�"�c!~g���<����昑%65A�CHu��ӆ �6�K��#�%;H^+m��7~��At����rf���ak�'���G[v�}B�ŗ
��ng�^�;��k����"n��{y�7��huD�����R�DR�"�!����H,/���H�B�٭Z#e��,7o�n�M|>�tNaq0� g�GVk �*��Mϖl�q�����M���.y,�R����C���%����d=Dy/��|o� ����Bw<�|���޸�4O���.��2�3����Ȅ09����q�4�H������p�w�G6��x���k��
\��M� �)-m.����5$g������QZ{�Wo�)?Q"�B��zbt�������]�jl�l�����>�	���5�p3�V��d`@�lY~&�Q "i/y3D%5����/���a"�����Lل��9�{�pAb��O\��.�Z�1��+�U�<��{����Q�rɮ>Yr�uF����Ǒ���!C2��rv�E���Uў�/s��,�
ߓ�g�wQ\IQ���v���:AVS�\&9�W��,�$ҾH�.	�Цug{I�}8��*���8Xs�0s���|���i4�G𖜶�f�C7��*�g�P5 s`k�lRJ�<�O�=4ݮ{��ܴ4�c��
��������ߕ9�j��᏷�܇ 7�)j���^�Dn��]Qbqe�@桓Isق�5���5�\��C0l�1�ѵ�����z���$��{XxjG�b�4�B����NG`��Y ,�D�M�{�0s�W��Y��'�0c�{�S�r���O��ȭ�$Ys�S���������$�M�m���O_?�x�q�����P>z�s��)t#�c�]�߯A�r��J�w�@Մ�~-��D�{�D�E���<�� Q��}߈�3!iĤ�h�*l�Y���IՁ#8�ˇ/n|��.��rz�T���6 ��^��4�^�WmU%�]����y��O�A��mP�#u�ܤ�	ð���-S^�NP� n�>��t��U����U�0^(6%2+�k&��#���~) #WM�3����e�O%�J�%����?
է���������{��ϲ�&�[mdƱ�2���(�_�dД7`&Tx���F��Yo����|�2~ֺZV��(��K����E�%D�Ҋ�?�����?��TYu����FV8.|�.ȕ~t�8-�؉oE������B���?�Y�|2��z��#J�y[�O{E�����\=��t��u�����O����(r΍D���*�����P~i��N���=i��,٪�=�:{kM1���>,W���ఋr�3����%l�����g�F#2�����sr��>�1�K3k�YR�����Ć�Uq�MV��M��>Kd�%�����"N������r�� )oX�.�4���V_�]aBJ�Ͳ_㱁��9�
H��C�������1O�n#V��)2�?_��(�,�_���l�^��7�ᛅs�O����� 0d3|���^4����b]��=�7i`�GG�3��V�u�h�������P�rm�B5��ZMM�(S�x8A���'(,s�;�A��}��KʘD8̅	���i��1Y�%��e�#+S��I�p����0�S@^�z���"���:C��^�<�*Ue��Y�G����D��߬���)�f��D�j}=���FMF�e��-��f@m�0�C�c��ط�H�Q���
���"��P����C�s��"�� F�;� 	u�S
�!��������띌�IH�h�^��@�����HREYiW�,W�˥�e[.o���:ԅ|�T�xs]�4�ٯv��m���|��v�[�D������p*��7Y�"|yB��NOs�c�nź�5�Gҿ�#h\zӷ���3�=ZRM]zmv�+W����ΥV� JC�r~�Z������kvB.㌑��CL��y�o�r�K���w:����"��)�瘎5� 3w�2k�HL5��Jz�۾��R��>u�H�斏���.O�5P���`o�v!d9��� ~��R��7[P�f�P��&r��J[���]]� �3\}:�����cQIy�;���F\#���J��V ��#�<R ���E�"��#�r�m醩\o9�T�R%,��	؂lM��'��b�������$Y��.n9{���1B�/t��Y�hV2-=���
�v����~�((�Ϩ��{�G7�mC.�$���i�om���si�P� *o3s�e/�?U�`�78���?�����ۊU)�֖�oS��z�ԁӯ7��g�	0��y�w&�zD��O�}�-&¹���K��f Xwk�1��Z�����n#��: �"#f�R�Qi#���4F���>Y0~�z�q���M;kk�r��L�G �U�o����:(�� �\׷�>���g���V* ��%,
��?���l9~�6�9*������&h]�[*h�}Y�N4�C6N-���G��qv�:���� J��y�����1�l5�+�S��e���o}zA�X��]�M�5���N� 	�H$��N����*[t��/����i Vs1�d�5�Ti�~��8]�(��v� #:e=Q��m3�x���7%DߦI��E̹�����H�;��Q���<�����.F����5�X��Qi�f4�d���|)�cp��Ť��Z��~j*��'O�;ˁN{5}�Y`\�������:R�ޮ\?������|kM4S�Xu8��Z
�`�٪��J~�=����A�A���AP4W�{�5
��+�*�:�x!��x��@﯊(���	`f@��*Wb�|�*@�}�z�]�������)��К��x�{�����~���F`�"�qa�f���e�C�uݪn��"^�����Wbw��7Ŀ)̄؎��p<F?�X�JK�98�A�э����wg�i��]�k�D|\�Ս�v��d�T�W�y����Ջ!�5�\4��X�A��E��X)EG�8��M������Y�ة��8���})=�@�\Ll��=��A����/�}�26�,�+�-,�
�h���.p��h���h��yc;��Y�my�V�|�{O�ȃ�F4�S�f���V�ax��F`sz�P^���,�[ێ�E�J�z?�����x�]r��"�#� 5��e.N��yĔ���0ǋ�O��A�K��3��"���,D�� ��[�rY�|-�ë2H�� �{=��D�j��M%Ӈ�7���K�y3@�a��ӡ���H��#.�z�r���	Â�3�G�-ƞ�t��4D�[���p��EW�=0��HMff�c�kd�Y&
�Z��ǽ���z@&����F֑Vʍ��&�EA��.߰�o����x�<Y�I��ZvJ輵t�G�Pוo^T���Y���_#� %V�z�g��O�e<�z_[J�RI��~zI36%f$����^`�Z��F2�耡c-nI!�KLN,u�;�b1(ptq�ay����V���+����������Bz�}oDv�f�5.>��rR���4���ٕ�bj���˰=Y���v�=Gp2�
�F��s�PQR���(��3��*8\2����ķ7��U`�."Z��E�n��0���X������.�3=wDƑH>�zB�[ �Mz�Ց�2��2!|z4�AP<�i�5�n�e&[P��fΐ���� Nl��#�x�:��Dg��̏�&g�DdJ=I2��4��ar:��*��p��h4h���_�X�g��*�O�<1��B���uɫO����G��Zx1�ż��V8^�%j�:�P�;e�O��jR��K.��F�KF��K����ߖ�%��H��+�Χ�`�9������>0������D@��>'���j��CcJmEgm`��b:�ў �4�[��[��ЁF�Dׁ��} ��F��ϣ�>gE�����	cC�o���	�: ����Ⱦ�[n���OY�&(KhX'���do��;"�C�Ʉ��k�H������ƨ'�F�g�}
a��l��T/kv��+F�ϖ;�Ƚk�p� ��y�q�Ş�Vt��<�IV{8�j]���z�5�,`�
���Ǡ.�9[Đf��U^)�>���B1����ȐG!���T�x�i��r|��҅��%�dc%����y?��⛝����WFD���
�������ȢyX��"�>�I���w��R(���2�B!�������S�iU�57y�{��V�_��@�5�cNl�&KM�/2tv���\���:qϏU�v��y���ƴ�DYWG6�����(�^�Ja��@�|����e�Hy�WR�P��u�hW�-���2������I��6[u�d��>�8q�y�_��#���$�57a���7�]�n4I!0�]��δ��"om��%��"�B�9vO���t`� >S���G����*�=�⿓��X.��$ː�*H��"P&�����cW���Ô�l��]焍CkkQ/�u5/� ��h�*U�}���߿�%p=����̽$��%�'�����JW�Æ�nR"~V�^�|�PPt����C�!��Q�B�|J��v���u[��v ,��� �+$2OέX�:�V���Zf����t� �{c��_>�\�Y�&ZDG�T��@���T��dg:EX'p��_D���v�2����Wc�9ʨ��x!~�0��U�+�N<S��e�`�xFa�{5y�Ib�w;��9�D_���!66\D۝>NE�J�QV�[��Mp����%����#���V9o�7��P s��T�G�&�����eɃ��J�V�4��І�qe��c�����>����}�Km��pd�s�F��d7"��(�0�����YA{U�I5���:��n��q����s��h��5�wL�6]ξmC��$`�/-�Y��P�"!Jo�*�.�!�T?�a�c���OTB�7�5��?��b�0#��) ��`���VAK�
��v��5�¼x�m�<ǆ�=�� �Ƶzˀ���er ei)^:�Ho�H���LU�\��벹֡e4<2�j/�C���"�O�~&.����Ǡvdyp��Ez�{\Y��k��4�_��+��w1��	���u��G�^�	�i��>��c��Vr���+A��iު�l���^�}�-�2�;@��W��T�JV)w,�	xzqH�Q�
u�ܢ)}��E7����`�J�hW�}1<I��u��m�o�$ۤF�|�5	g����u�nc�9�S�,����z��O��&��R[ �"��跡
v�o�|�Y��,T�:���p.�m[È>�`����DW+�0��<j�V{�F�ؠū<!~�7bԿ��$tk����JH)M�~CK6�P�`�	I��B$1�ɾ^��~8@u����\����S�y���g9�K(C�JV�>f�@-��r*��r���G*�k0Ѫ|�{ �!��O%~%��	��G-��`AP[�J�t�I�zN���D�@PЪA��V����1���4lҫ���}�s ȎF?$d��N�]�M�rW�w�+F�$#����A�F�H#p>}��"�M���&�X�I��BJa1r|��s_��ވ�;<���w7k��o�4<G	*�w��%Ⱦ$��̻2�	�#�;�Ps�dH��p{G��$�L�c��a2�ֱ�I����Y Օ� F�9��w�z��#��n >I�x�� k,�L���޸��aH�,m5�����e�$���	�����U�g���,�|�&~��k��K�ւ�')����t�/���P1]�!�]�g��oO����υ�ŭ�L�["R�\�u(�Z ؔ+��V�Fgxan�ijz(F�"a��LUs��=+3�۸n��p�=#��0�WZ[��d� !Z�٧�$��s�O����Ѝ	�[�L���z����dar���ywN2��ִ�i���,��I��N�w�E16E�t��d��$�f8��v���SH	���cv�K	��!{�� 9���{af9�?�B�U�b�++o�z�T��)�dTC]5q��u��śI�d\`<�rJ�@1��Ϲ�NC���D�9㏟XD^���>�E3���]��R,�����x��[y��'±���K>v��E��ô~>B��P�Rd���E�y����?�t��F4��3XQN3T9��GVy�]n�!w��J�'����W�>mr�)��f����T�WX�(��U�n}��L�d=�*d��xT~�����I8��3�l��O���$�tGz��U<��)�B�p}��e\�G�������?`7~�=9W�P�?�m��N�x�|*�懓s�L5!�����Lh�4,�&���k��|;= G(�%�1���p�	3���XB�%�1�v�c��<���/G6�8��s�{�n�g�K�6�i�|��l�!��Lj��x�8'#Җ��p�f&O��tu�,�W22�,� �,;��C�ufOq�F�V��B���C��w� _��,;}_R�' H�w^q�~I�5�i���#yX�6i^=�E�Y1�E�a�<w'�����#��� �ư��N�f9c���|�����'jR�4����Y�2��z~��3�H<~F�~-�xj}S�5�c�c$��!Fe���Hþ�۩Re��=�w#���R4�v`,n�0@��?߾�n����p�${�e�C���`�8������(�[a�hd� \�A���1<z��a�a�ɀ�t�A`&*@Si�$!�]6	�� ���J�tO��|)��+Yq�x}�R޶Y�DM���뿮��� �+Vl�_.�5#�qc�I��; �xR9��Ṷ`���
>�e���5�o�Uo+kt���zH�������n��xl9[Fh�ƫ՞.��;<5=X j^�~�.F��Ѱ��}��׈��7ɱ��a�O^�G�j,����e?�!`��XGߟ%B�,/:i���2%�&�6�J���9������ ��̒�pV��k��by��Ȑ������	XQ�@��������E�$Z"�ݚ%�N��p��nH%I&�������/R���,P+W��|������5�BFTn���"�)�:�Y`5{넪��|����a1[�ɍ@��ιZp�~#Ѓ}���SH)��A_I7�^�Գd�U*�z����S��"�����c��qΘ��%�t9�/P&�&�x��ys�e%d��1�'b�x�ׇ�0��t�
l����7��b�岨sv�]�����W� �}����.XG�bHC7�;Il�b�~G���p����*9̼C`6A"�M9�lZ��WSc�Z�w�vnf|����L�ĭ�N;_R.I������ojM������ ����G�ɀ���l����dUVԳF����I�,�={C���#�ª�5U��x�	�i}����*��.�L0)��7��#e�d�FU^a� �X澾���9H� ��C��֧�$����C�΄%�	-L�j����������e�h0�Z-[��Q��[�ɱYR�v��-
>7W���QZI�b�v N�E��<>URF����)<;����.��j��T�KMΘǫn���HJ���I�G!�$%��*ђ��Ɛ-��2�� � �j} `+#�:M@%�]'��p�#���x��O ���>�F���$�:��')���_A�Ӎ����<��l�e1�{�P8V{��z�|��^�BY��-�v)����}H�j���0p=�~��7�X]��@�Y�G���AAYl��Qq\5T#��i��Ϛ}S�G�(3~F��Xq���༢�`�����Z>(r�I�z�:	�I"���Z���9��/���Ki)�
 كyi�NF�VQD�]���_E�B�FY�/��a��E@��4��C�6���m�(�����-1��<��~.8)�Ji�@�UڋF筺��JF�E7�<��y�a�@)*}�F��>�����>�t���+:��G��g��TN�:��?���ĒÞ��9�s�D����;�.��@��x��(��T3��+&�%�`�Op��O
����n�"���?S�������L,31�� {�;;�}A�������O�!tEF�1��4�+!'�0r4ܤ�{�[�xjm�o�bBj$i:���#;;���[R�S�~�Fs��5dA�����3Sx�P]�����L.8 m���ނ�������R貣����2��|��2�yU�x�0R˃Ŏ/�6i�з*��l��� �d��8� џ�Ufh�[�?��,��GE��~�U�+f��>d+�%�h��b�����\<�O4�=���?F��Qq��b�︔����a�5������C��jޮ~���)����H\�9��IS=na4UA��i��}
3��ш�1�̟�,/�.q��ĲVM<݌@�%��u�K\��O|�5��?�{�z#�'����K��J��V@O��Sp�3����f��(M���{L�j��2���_Õ�)��\�z���nE΅��ٞ���K�S��̙$�;�{�!�N,B�h�7j���0z�a�+\t�͍�`j���G�ozh�|G�1<�a(�IW�\b\�	69��I��|�L3E�+o�q���4�b%�Q�����-��L�f���hh]H
�FK��m$��vyA!����O��_qW:\# c��HH���+��nY������/��r�݁�e�z��-@c��P)�����\&xk`� #�	ژ���{�@�Ы��XP�&=�^���jFv�ZeJ��E�=	2#���OX�^\�� e�-!]�����3+[� yv�7`��P �ݛ3�F��n���=~��ۯ�a����5,���OŜG�����[�����K G>�J���3�m��<�p�^�a�,l����M�Z�[��֠��1pnZ���������r��x��#t#����6nO��a#�rI��.��s�աR��"�c��p�4|�QBC>)�8­6�<� B�GB�>!����C)�Q۰�gR �_��������ʐ(���^�@�����CHe��J4�g&(�y�g%/
8��2�!9R�6�$�U��� ���q+y�8����!]�o��Js��3�Y����|�ʌ��v+��������ܪ��YK8����{�����v�Շn[=q�Bm���ZەI���t��()g�ܙC��_������ c�r��oc�_���/�]D�(M����F(>�l1T����Z��ǵ�=�U�S�sƤm6� �2�v�@����3�C��]���B�	8_�����Y�b�P��y;R���s��.aO�����e3poE�K�Āv�s�E�ٟt�A�!�@��&�۩}��Ŷߩ���@>�[��Eb.��[{�,{*�b�O�� ��lV\3��t���2��(�ϻ��-4��I���>��Nw��=��ȗ\ĹZ'?���e\�%�(3ULNս:��6BoApo���U�<]4W8 ��9k]0��cZ��+m�Ȉ��g%�.�.����/�]��ǂ$�o�/L��u�ۧ���F�f-2>F�՟��ޱ�8�>ӿ��{�'�\J���I4�$/�9If���9�, Wn?����_�x��?�;���u���c�4l�&�(�� �by�N������~X�xH�=���+X��9�x�
.�����f_�C&z�{[k�Vxz?�G7�Q!/7�e����q����y�/]���[du����Y���M�S�</�:���]
��YN:��V�~����x���+w��9�����Zv+X�e�����S��-hs�E��ܵ"�҃�mU�����e	�d�kԆ*b�g����}��u�'Iﶥo�^�����%�4�Q�hDg������>�i�-�is�FxQ��������~�W+�A*���]�9ȶr�H9Vɍ��ȮEcO*q�X���9�QH�r�g~�C�i��G�\��ĸ�8�S�������Mu�F�j�Q]�����5�Ș)�J�LX�������7�<8H�C� ���y�[/ [�
IA@�����A�h���țTXC����5�m��XJ�@��U�.WB�ϥ������G���X���bk9.p����Q$��� &�/������ѓ�wS�J���3��&���M����,DO�p���q�V_�7
��G7l��.Z9�����Y�9o_|����ٔ=�gP$%��t�TJ��H
��X�M�xd�&��jf����ʹ�.5ˋ�F�h�O1W�Ʃ�j�&<���'Ol}���@�5�����������K|��L�oT*�a�VS?�Y��N�e.��Z(A�qm��Y�C���|!�xhM����p�+��S��4��*�^$ڸ��oAonG
c�l��߬����<p��#�/:[�x������Vw�m�ڥK��Q�:Css̺�ӈ��DO������d��+���_�т��(l�P[=�K�Ɗ�h�e3�۞a�ם�]� ����^CI�fHs�B��{����'�۟q��F��Q(4�n���s��i^�}`��x��$�-x7}E�v �Eb
�gv��z[h�{Ľ^�VN�4o�}.L�0��ng���'TZ��.���ʰ�K[S�[V�u�6��K��΂݋�ᯟ\��F +0k��V�H��[���O��Hq�[�,&Q�� �<�2��G�CB[oU�Ė����iBuQXX��j���0|�PSOM��"dˡ�g�ɺ��U��N�j�@v&��xP��;��2�"���EG�s8��޲��~��~��h�iCz�4��otyc�-��%���sϬ?�* �.��\�|��9��2:7,`��,�%'1��(F&d	T+��$��������z᲍�{*���$T���>��Z6~|/^'=!z;Q�U	�Ř�99h"�k�_���5*��Puw�Ln��!��RW?=8:'Q_�߰>�\��3������m ��ܜK��T�mc�s|H�iwGI��JUmsP����1Ӈ����A�@TX�i}c��	����|7� <��x��a�}�&�\J]�~c ���t�{5��S���u�U����4��8�r0\�G)��%���| 0cR70�2��@g9o6�S�5?/Nl��i
��+�l4�Ф�Hj�����N���iŏpRN8R��<c�Yc�!�ˋ���/xl1�3��LrF�k�W�:�7��vwԠ3���.nd�+,w	7�ѓ�\cD��H�N�ĉz��,�wfP��9ڤ7 �\Εl�`P�t��Wn�N9���I���2�VKA��r�S��ij�!
�R� ˕��vl4�Zz��BuRz0e/��Ō�݁�I��;�{(lu���+Ӻ��i��Ƣ���٨��Iu�)"�um�b�$�ݫ:�'H���H��۲��T����eao|0�6l4T�θy�+\O�Y �
�Iޡg�������T��}-��I]�J������W�a����A� 
����$���<
�_s�x��sAx�v׽j)�P������^�I�^bو��G�cө��Q�鏗�$��/$;�2[R����Ʀe��k����j�	���1��/x��:��~l�>T�����D�m�l,������ ����·7�3'B�j��J>tx��#	�O�� ܺ[!�����~�(ˌ�����^�s#��(���i"Qԣ�F�@=��屏���1tI���b!��8��4{l��¨�}�Al�۝K��!�i)��A96_��:�PZɘg���� �}Afy�GZO1���<�����$�x���e�n�v� �#A�:r_���R�8�K�E/��!��yB9���d�R>��t�X}rpSF���л�A�`?��W���6I�493.&�O�@oL�.|v|%�Bw�0�H���[�{�&c�y��@����W�,rN��G0R�I|�J*��Ž�M}���;�%\��R,��"Wz�X�AƱ���+���?I�<���,FF/�kt��m(�~���	AC��+�p����6�Q��Q}P �Pn;c˟3c/XIprq�B��r?݀z�5B��Y�R6r\5	��ob<8� :���*���j뵪J+4X�n���hJ��[���y���,��m��kA�
��F%�(6U�|�5�������$�������8���2�f��P�^cC�^/�fUL�*Zю����_�Bҵ7��-ITS׆�x_���L��*2%��(�]�iɎ���)o��������4ѧ�_���f�h�H>dK��۱'���'�<�9�x �^c�/����+v ��H�T���\M)%�q���1��ͷ�EDZ*�rօf?-ڑ�=����M�+�:��6K~1�\�������H�~{a(WN��Ї�汥�U�D�%V�?�q������Uڃ�sL5#�
x`E�v����u�[V��e��S9;��1}�ZQ�Ⰱ��O��r���ct���q�
՗��u*�q���F�U�oQѱ[<�A���dA�����w��Q:}��ь�����1Ċ���$��Y���η�+D���j�ћ�j��&�^4QD�ͥ�'���S�����7���P&�)�:3�br�v]#&o^�B]�|-�1hU�f��#Z��M-V��y�Ȇ��_�]�3~�P~)�;���(O��+J�@)f� �c��E�|������]<N���l-�N	��w=�AYl��	"��"�*�,Ҭ��c���S3��;Hw`'/@��.vҰ
�9�`4��sjJ�{��g��N�4�h
Ċ���D��*��}��:�)�@���ƶ�b:M֡���3��M|����9|�ǓVT
�`�L�k͒AkϰE/�}0���G.����Pۍ>{��7�: ���. �;��0XZ.[�1�<�v�f6����j�bI������2ax�tiTvЋ�*�L���?R�L�S���!�2�z�N��F$ˎ������
?��+������8�ֹ�6�AT�Ⱦ{�Ua��{*��&yomS*�x��F�`����:%�E3��%�ߡ�S��'laA�������hvF�*aRx����`�����,��s~�Ɗ_��򀔸�Dd�F%�x��s�r�i/7^�/�z�_�wpy�Z*�@�}�6��
���8��.�1��:�[�,��%>k738T-���;�3���p��Ζ�v����J4��]< <�qtM�j�h���*.�HOV��ߦ�l%��j\�f�U.��{�G�Q%�89��6�͂~���>)4ݍU� �
��1�8�9�x�t�w�.�?}�������0)�N
�f����}�L34y��[���h
��-KL����jڀ��;;y��>�Ö�Gc������A�:�n��k]x���r@b-9:!ș�$w8~+=e;�:p#,p�,�&r���?�Q��b���r^���鬔�W��\�)'�/��6���֌�Z/��mS�2��B�1#6_54AJ�V,o�&�>Q�gvZ�\�-(b�g��q}?���cHJ�g�� FR���~-��B�J�T���@���vw���<��Yp'Bp'�"Iע��'IeJ
Q��m���t.8������Ri���t� r����t�tǧGȲ�۾�-�>�Ws�]�|p�����ь�c��o�D"�Q%�=LZd3������ԕ��X����ox4��l�uG�,�{��3�C�G��jg���*H'��+S7y� 3Q�ǲ����C�l���A�����)b�S��E��D���bW4׶\L�Dt�S}�l����a��R��Z����/C�`d�� �;���ú���H�_#!�����}��r3��;]���l,�{�0�Y;�3���l������������V@3�ҷ�	Xt����=�����I�������s�F�2e�L�*�%J��s��s���n�H7��1b�,����V��L�ˬɋa��v?+�����"�GK���{0A�ܡgC4�L ���&�Oq:0p����Ǽ>?���h\���)�V��f�zO+z᫡>\���rM��?*4i�%~"��p{��񮅓7m����M�&ً����S���"O�'�P���G��������5L'�mq	�C+���(�F*"o,d���?�_)d}-AE<�� B�rH��x�u�8v;��T�'�?�h�ʹ]n�<�7�N@����/Q��E�*�g�L_�©���\�^�M��Y$�\�cI�SmO��2�;lc�ԹY����U�h��xЦ�JG��H��]x{�?D�B�����fzDС-�U����LS����ºxԍ4��np����S���R��u'�/�"����e�l]%���M�8v���h`�q�a�y�"]��GG�i�,h��:.BW'�
�m������E��:.�w<�����f~�o:,�i�h��C:/[����_��=��"�o�=v�����]��%$.:�@��f�-�Ћ�e�8��o�p!Z�����G\�Q%�-u4x��|!U��D?��o���߭c�"���4Q�ig�h�a
,+c.Ҽ��$�$��j�=#daj7g.�����-p����l&����b[���^�|:r�w�Q��3�3�Xu�p���d��d���֡k��2.���0�����y�����ʼ¨@�t�����X��yZƚ�Ğ�8䀍*����<F��߸��V��g�\�1�w��L��X�
'QN�F[�7jܟ�o�)W�𘁉�!%�g��/k, [r�N�wJ��)%�xވV���n�/φ����U߻&�u�}�?�/����A.u�e�D���8e/�z8���~�����Vp��j��K٫qY܇P2����#�2�o��
3�	�E���ŏ+!�.��%Ƞ�E��V���d�	r�����j������k�m��~�η�8�A�tv��R�}���3N:~x�l�S%.�L���}��/�tl-B���\��m#�� 7��m@�XQ��ֽRg�U�V6=��YbG���&M �4�;=V,]q���yW�_Ov�J W��Q=�Ȇ���d�1��$����G��Y	�x���ޯomiV���@�c��M����8WtD���WIp�E{uFU1�Nj.�@��d�?@߅�T��f��+ $� ��r�2���J��9���h�ѵ��]ϐy�ė����$f�wW���2;�a�3B�H�)��e��jJ�� �ˎ��i���z4]o�}J�H�r�R�z�*�!��R7,y	I�V0�~��%�5C�S��6l!�"NG�tV��5.;�g!��m.چ���v��/6<���P�+7k"�t|���6 )ͩУ9���y���Ș����t+��x�'�ns��Ɂm�E��||۸�C�oD��0��5pw��
�}�g��قO�s)yo��jz�&[(���D��&5��T���q�
G?b���D�^QG����9���Lߘ%��D	�L���l	%Ř�a���[cdc��3/��������?9��P�X��\�����(���ٛe���`3H#y�((��~�L9#��̑2��zyNI˨(l��� ���%�l��1���J~>,�{��o���V��h��ɾLY�SΝb9��޿�z��j��Q���/|Я���w�=��
r?�R�ho1k�Q���b�~��L��@�`{1cM�� ��d��vB�z�WG
���Qe��Kg�MP�=�����D[b��Ї8F�����s�����M��!�t3���-�!R�7���P�-��N65	�7F�dC$Ƚ��k�(yc�W��^tr5�x�	�OugM�Iʊ�#,8��R<+�(Ch#عf�m��~uI����V,2�C-�j�?.%V�l�'�ڣ�IHcV;�gVnUn�
 j�V��e��y5�K ������nU�����~������� �����s7����퇋DT�">�������K����������"C&1�!�2OLV����N%瓡�D�$�qS�GI�Q(T7:�w2�٭�ح{B�@l�C�Y����i�s�CBj僼�:X�2�q���+�E55��C��gJz�S�?7�r��Y�H��4�!O�B^T2��DJ�`{{݇��F�Yn�$����~�0~UP�� � �v�l�����@P�nv�t��J� �#�%R(�~ҜS��l�#��cM>�g>w�M��m� ��yI����ވ@Z{i�k,7��hU�W��n���hg�Q(�
�j���c���q49]$Ȟ��[��m-�]Vk����m�_��dnT:��$��%kv��W�4��ޣ���{*Mq쨌<4�3�V���m����$L�㝠��!~N�[r����Ԝ�W/��n�-~��@g��c��:�f���+h�����O]�6��7�'N���\�#~Q��?�!�����D���7{2K6N����r��c�t_ܡ����pA-Wsw��Y���/�}+E����}m�rQ��RW�x�?�r�'�!�}�WIm�O��TϟkA�����'��X<-�/`��!�ɣ��0����6�s��7*����nV��s���k�wi��rI�8����<��Q"e�n4�b���]��&O�mO���
���=_._�K�
���FA�Ǯ� 
b�y�E7ފ��0�p}��֚�%����;�7���D���)sա���#�P��%������M�T,�ǖNg��	�ӄD�C���%LຍEF�L#�ⵖ5����"p�SU&�9�\�V���v1���L�$��K�KE�c�	п����l�,k��?*=�`�+M��U��2m|�ziw@�*�{:��RD�X@l���qD�8c�?����B�I�l��aXx�
"�wsa7��*��ܵ^�|�������m�X��>�@\&��f��U�7�`�^au����۸p_N�	���\�z~Y���j�<��*r���/H�/�y���yf\�<zcq������Jɱ �p�%(�r
x����VtsX3�z�@{0�|^6�ON��e�s|v,Gq���y����z�O�Ya�ڮ��e��I"�ͳ����Ղ����߱�@{�!�迳-$|,a�����mF�
J�h���e!i# !�E"�L�\�a7���P�����ӓ$��j�����������b�i�fVTj1�e�C��p�I-��&\4ń5�~����^Q;�W<1���g�zM4�����<cзPZֿ��"� �d�M����4�-m�c��"��۝�el���/i �酓b��o}��/a���|�X�nt��;w�Vš��'�M��m�hE�D���T~e��h�=��T����0νEֆ+*a'��x��Txf��:eC�a�M'^�����_g9��RT�lA�ݵxj��+^Y��W?ٛ��Td �[x�U�28��Y-x��m+q�|������(TK>n1���[q"�����c?�@96�"��r��_]�'����B��W��G=6�}���� ], =�G���Ɇ�|β��5�Y�cM:|jVd ���O�Gl��rf���_�3:�������A-��av Ul����:���:�'|�Bc�Nϡ�ɋ�^Ӛ��t�O�8,@�Gj�)냕m�
�O^��H����H¶�v{�v:�cs�>��d�7s�6D�5�50f��Nx��;�nw��gMW��5�<�L͏ik�D����,*�������D��a�\���RSO�n~q#��1R"�Z�$i�Nޗ�Z�\������6ɫ\7�Y6p��82m�~C��X�yr]���J�tTT��B�K���n:�Sg�����I}0��|�q.7���s͕Ae�a"�U���^�˗�̓ŏ@�[r@Պ�Ct__���-*Ɣ�㤓`K�]VڕUX�����=m4�?<��k��(,��36�b�-����y����	�3�k?h���Ic՞$i/M+� ��K"r3s}֓T���l $�"$�.]x��U���1bO�K�^2y�L����o��ď��s�xqS��F���I8�]����'����s2�$�����@������V�c��C��/�&���I��(��
(X�t"O7��g?ߓ���z!L��� �S�ֆ����9�i�S�w}��8��{��I��{�k$�o(�uЍ@7��͓p�;�4#�T��p�9Π�;R-�v��j��Z���=�N�ꢿ���z�@L���gO��+�bv́:���O� IZ]�j���T��D���ugX�=���+����7��^�4��e���AP2���k_t�%F�V��JV�-Y�G�,���%^��v]����/X� ����$d���E֍����}R��A��|kE�`�7���X�v�-1��ˡ�C���e.ï.�}7���2lJl�H�sm��$E�$G�;� Ýqp���f����˨\�\��a+�P�!�c+��
�Q�#��1L���r_�܍�ύ^�E\q�Zі(T����3,��r�����l�v����z$��]EC�(6!�����֧���F)����� � +�mIo�F=X�m�g���1����e����r�*�sg��������
�nMwMC'�YJB8�1r�Ӗ�"�*u@�^b����<|���ｷ>��5�E�x��d
�T�^�hP_��@����+P
�a�oK$%.��,�Il7F��A�� `���3dk��o�Sr��=�>�*���	zC܏$~��0BJ�h,�@Z������lV
���Z&��v|,�fh�o����N� ���+���b�#�p�lQˋ���V�U� hF'���n��=������ʾ��(�?���ΝW��LN�e�{q��C�ꌜ�E��U:ÿ3$-���b���e4!fM%�{K�p�.�W�GH���ܓ�V骿�=+X��:��wC�� ����!���<��bO�eZn�ت�X~V/?��w�u�
 �U�y�Z�=urlٝC�u3�4���������ō��	�����W�H�#RSl����M�@*xVPY43�xW&zL1
w���n��]��Y�3*�X�p��i�ר$[68���')Wۥj���T#������<�� mc�4�x�=������E���ϗ[����k3U���u�뒬�Cc���
�C�V% ��]�Ք��7D+|e���#�J���q~9�U��y�g�Lg-�kOgeq���>y|�6��r�J.�~~��$�1�-�P�q������e5J߳����9.��i��d=���- t�h��'!�]���@9���p��4NS��{�p�N&ܒ3 �0M��Y�5'��'lm�T:��j�-|(����b�2��:J���U�	w��u���)K���RѝZ�[�ޠ�t��we�Cv�>�I!�P2e���� 2����d�$[�;lρ
��z��m2Q"`S"j[{cҾCHb7�g�hcoJOͣ{�RH",�҆?QCs���{�n�O�y����/�QYEi�c�,Ѽ2i\���^^�I��Q�j��Ƙ�ܙ�=R��6��o���~>��F�H)«��v�a�C{6�'�.?~��!u͡��_.��"����иbsk�e�
?��*��{:�����a�{\�@+tQx���{�H����A�z l��	���RkM��M��A��~:Ʋ��yN���r�x�u�#Ő�Tդ������u`h��#Y����+��?i,B��]gƗ��Y�q��p�!aK��k*�,@�C 9�g)}�ڽ�m؊���W}�ى�7g���4��� $Pg��-�1�V��ֵP��n�9o
������A��a�_�}�AY���Q�:�p���6|g/��0q����!p�)�j�.S�6�}xE��{��A�-]T=����&O�C�^Mn�u�t���Wʕ�9��8����8_ç�z�=�����~��$��H5{	��!�8$`uwϸk�*R����:!��!ݝR�=g�W	�In�$�e�M�������e��r�6����t��>l��ŝ��C�t\��)RAr����Lpc���b���a4C�P��	���Q�&l���y�{���uĭ�30[�Zܳ]�%n�CI��e�QI�	��ۨ�m- {X���௼z�C;<Hn�C��m[A�T|�O������2�W$��i.lby��"�`�$y�|��ٽ^@�mD5t+œ�e`�.�=���a�3�㤢J�R+�� ��^��Av���	"�g�\Ge ��H3GA6����p�MȮ9�aސv �n���(���Ls��S�p"r���˼Xa�m��9fv���0�Ox$rz9��2�B��Ӗ��
��#�a��.��<!H�^����0��߽H ��8����b�0����l�~���G�v�
���S}���d��8�T�g������o��[�Ҏ3�G����ۭ���($p�F�ѝ�9��8��n��ݿ�cvfbjJ(����_ȉ��+j0ĿzT����{�Z�8(:����.����x�YƼ!H�r6�oЈ��b�ƴ}j]ǰ57��Ai,�>ӈ�Ģ�ھq��+���M�=-�U+�b�m���JĠ�sm�������j`oX}���1�ۃ��ٖ�qFY�ΫS�����R���WQM�����ՠs��}����eg�j����fb��iѶ7���BX|+��s�C;�M<���Ż��JL�����|ɀg���6f{ɏ�{�M^iB�c��܍.puv�c�yk�Uc����Ey�ȴm�ox��oQ��m*���gaopҗJ%0��rb#î�Ǹ�=s��y��R?ű����"(K�<�ѯi$[�G[�׬�0&�,�s��BZ@g��0�͜�V%����`�ԁ�'�����q����g��cTD�C|�4�1�[/DNIar/W����옃��TqB�0��%t<�����z�]�ZS���21XX�>�N�}u�som��Yu��������鈏�e_�u�`�l�Q��DҼɗS�^bg�4��s*9�VFs����#N�|B �QxSI��H�Rz#7�����li���C�H��/ӱZz%�e�Ps3��6�i6,��_0=l���~(�f�@��N�'��(>���IG׍U���Fֵ���*H��s��a��.�&o 6 k��|�ۜ�,��,:$S|�f���$r���:F�(q.@�~��z��F������L�F�jF��-s����:>�xS6����=�����gf<�F�BDZ�r���T"ڸt�z�K�5|wg�J\��S#��{����c8��s1����-��3���g�Ĭ�tJ�H�����G��+;-��7<e�'���2����|�k/�?-�B�`���m��֬�	�q����^-qSն0��XkL!g@�9�}d�G��e��.f�n/`�J=�~=�!����U���!��$P�Pq�u'*�d���`�4�0���������%$2�$Ϋ�{�|$YB
�"������z��㨸�iPblE³�&��J�5��=x�6��I:!Ai,N�!xm�O����\$͑~�?a����Nȯms=�t���¢[�W�1�Y�M��#+i��d��hw��+�}�{J(+I��p���,�з�טE�B��8뉽���B��g�Zl�Z� �o�(���e�)��j�bL����;0��4�c�q�d�<��-Q����ޔ#��u�3S	�'6:t	��&m�&�t�%��z&>��~�N|��(�o@�m�����
��{��o�.u�<����P��e��*�)ŋ|=h�;
_�p42z��/����x/�e���L�;�,��N��ES����>3�W6e�����P�d%S��"�"�ɐ�m�]�y�dg�䃋ibaV0��������/%˼|���u��R�¥u�\e���i���.\�Ce�T�����_w�Q驟��Gl1ߪ7���Hg��(��ά��H���̝��g�4:O1奸���D�T��_V��f�����8��U���`^�U-���΋,2MS�	+7�3����ә�md���4&6PKz���)�7����eg���''I�+E�ط.{kJ���V.�=���$��ax3���PS#ٓ�1Q�ryf���WK��O�'�cӐPӄf�Q�cG,���ܜP�;����s�r�d+(�Չ��G�8��o0�{�d�h��X� |_�(�e�up�F¤6����~�w�C<�LjNٕ�~B���/.��������os�E`q�aV�x�>�J�M:��%^ƻ�v������@��(ܕ�$����m�)�}ר8	�$���E�&�J�Ͽ�#Y�v��Y��d��_������̗�~H�j�ݞ�*���Ua��1y1�4l�oG)�j���G$������D���kZ߫���e8hVHH>�4�8%�����^בֿR�Y����mzL���kuZX	���e�'��y%n�b�A���+"ES/I��rD�Dr]~�k�hɪ��$���#����6M�`>�a�32}�F��޻�Jl~Dc(O���,�|Hn��s{�hvC�>��ܹ�Cz�.���_UL΁	s�Pò�-B���Gpg����u)���E�.�h(��o/%���c��PÚ�Mܭ}؅��*N�߆���>��73И��Zԣ&w���լlI�k�-�mq(.h�1��c�� �,�u܃ɜ�dFl��U�+��J*Z�M2�ìJ��=�>M�`�8�ߑ��d;┈�Uu��/:�L���p�mm��%�{�%'�t�O��BP���+R���� �˧)�t���v�uaO��i���i�Xs�v�������{VV�3�ā��� v(�_3-�BL�I���O@�����.��s$��ٝ��~l���p�}^/sԌ"��d�ռyE��{����X��q͆#F"���4�2�!��p /����PZ[ŦW�����A�jY��|$�B�R�NM���e<'�5>�V���PK5&�?V����q�+�Jx��R�r��<����l�������]��0�Jt�I�]X�]0t�u�e&���ۡ �#nF^I��T�=���g����=4-�+�\���0�Q4��u���"u� ��\r��R�R��s0��J�2����c2)ޫ���	���cH�2GE�d�DP�|O�����'�B�7I>�6��J��Z!y��	`���8K4�,�yܴ^�����(���`?p�P7nG#ه�1f>�A���m2�И��c��s�6���ܾ�����~�U"	'�jKQ���U��K%�g
��Vc'�����H�ņ���p���b����pXΛ��f9�g~6YD�9��B�smŻOR�_�g"-���;\�����7G����O\3ŕ�-�D�f-�j��}XmfX���Kbt*�����H\x���f9��ly%k�F��M�j��&l|����C˙e�c�d6��F}:X-� ��ǈ7��BM�8��?�B�D�x~^��m�C�>�ս��5Zfq����@�+�LN[|ĩyN�g�Տ�o�ڧ��xH�;Nv^�z���{9�#.�("�W,��n;����ho�w��6� Z��������r��-��`�;��e�M�ܰhm��P���h>���bx�������4���h�ڜ#�x�iI1�Z>N@9��T��?g�"t��9�whլ���mX��P��g�+C���)Ɏ�7$�h�K%c��p�4M��|R�(2&�YPO!�n����:DS�����ڦ���C����zu����G�@ _n5���<�h����ݵ�$�V(<�R�\�v�AjǍ%���$�Ş�=��S,����W��x��l��pޥQ�=�4�g�dTE1� _-#��J�f%jA%�Ǉ�F��'1�\�Ӳ�����J���v�c�`�vG��Pi�%u����H�]g"�S�@I,�0P-��w�|���n�	�Yk �Rj��t�]ц�S[���Ԋ�_�#���{J�����T1�%���2}��ʩ|7��e�4��d�&��*th�!�4���n��4�Qfx�%���z�D��F�Α,A����3,+�D� ��R)%$o��7��;�]��9�n�~�������X�6�]Kk�l�J!.)�pml�	�j��O�鯆�S�f��9�����%�5��,������^���'V�G����%T	9��dQY�YJ�*��șxc-<������$�׉�3�&�YmY��0�:n�K�X*Y�ꮏ���0J��Hj�yT���^|�4Π>�i��G��g���h|�]���ӛ<oY&�#~��pX�A�d�*�-q�옿�����~{�ֻn�:�z!Q��|Ԡ�2��<���.�_�%�1�=^aǪX��q%.c����ՁGG�[��I���7�3�F�D��]X�AE
@n�:Ǒ(׼{�G�])sU�_O|���}�쨸�����yE1�����z�"�R�X�R��E��B�f�Wey��8�� �mN���?P��2"�s�Y��ߦ�)؂ywh�P�~[ �,��u��9"EGXc`�% �!���/V��b�9Np��j�޻B�=�T[�%�A3�Py�|KD��iİ�-��^5��E�.�5�a��*��X����mK���yg^ib����w��0��H���a�^�������d8 Ř<R�*�(]��k�����o1��}M�s zj!İ罗�&~�dx�!��5Ǳ}��5,B�U�.�c�[��ٗEփ�_��,�5�+>\s�����x����mE�W�b�re��/�-ɿ�ΊG;�KO0>�X�[�C�J�B�����a��x(��1� ���1�D����ޗ�`�J���*�Mީ�#O�p.)����\�}bYH�m�Fd����?|\��1��Y��
D��5�K���`��W�:�����f^?tX�r�
J��9��[�M� ��@���'����eX�ڰw!Q"��57����a�$�2����(W��e3�7�u=�3�`IK�YB�OLh�-��6��n�����A�y�Х3��݉i��,����B���7H���"	�'`�K�W�XP:(7��k!�M,�{�[��η# �	���1}�׆ �[�G���sI���q?���T���s�Li9�"���N�n~�Xњi��������f��B}MW�x�pB`�@(��[[�׶�⥿-뜰1k5,6��i`ғ>3V?�%�3�ʷE1!�A.�Y�F�L�K�ܔ+L��H�@��);�D���o�y	���v�˴x��|�W%�>����/��ѥ՛>x�{��R8�><�Af��w�x:��[��|m*b����!�	L�%q��[�� D�.i4�ڱh8�G��TS�D�S�wN!�ƹ!渐� �pZ;�2�|��j�pU��_�D�a���aK85�8�����`F�%/S�}QVa�X���F�>�����TE�����<5�Er%dJ=���[�y�w�#��x���b�$�7�����D!�>�^5#ʭEL��l���Sб��hR��+�기ُ]+ri�M���p>�6����@,"O=�n�)(��Oԅ6vz�����U;��4��a>(T`B�!|��bͨ勶��wI��)�����J'Y}��u�*��>����~&���զ�9�V�[vS�,�h�����b���O{��C̠�s����>�M�&/r�:���H�T���,v^p����WX�j�Q6�'<�k�W�b-l�W1N�ڗ!��J�'�X�dW%��돑'�Ӑ�gq;� X���Z���fRׁm2h�.�wɗ���j>)���Y�T�JϾ�kO��d�H�#YVa�������������{jl�2Sʳ)�ߪ�ӂU��J���$�D��`hx`�TZ��qƭ����-���~d���}]�5%�f�&,��^�,E���X,��r�8�F��vG�֨i��l�"�5B�=	^z�t��P��A!KZ�{��hr������,ie�澭_!>�F��b�n�Wnvr��&U�u5�v�'�p�=���
v�z|�{˪������B�C
A�z7eC��r��q1�ہ��c�ۖ�oY�� 4y��Eڃ��
����-���J�yO���8��3�>�{���D�Zr��n$�X╰`���L���S8���TW��~Fg��\��I1yL�D�2����IqG�ޫ�Be��T��7�$9a=3|Ln�11�K,l`��&�E�<M�Nu�qh]�2/I{�9sV~�KGW@ܕ��n@���t���g�EJE�����	b�<�m��^�>odgr��1���8���buі{\�[Դưr)W���{�DWq�9�U�S�z�-KR�=�V�@����eʼL�[��Q=|������9`�3����J$��/L�V�#�0�F���z+e�<5+ �v؋���5���=�Rk'�Fe5�+^6%"���zpك֕� ��ˎ��:�wt=�t��h���#�!�D�Kɭu}փ��9Zt�@�ZJ+Bd���y�=޽ k������o� @�pm�}�gAI�����h�9ӨQ�^<Cq`o�i��ςY2��-���벓�~[�
	�q�4�R�.����?��#![�C�4�l��b�zJ�4��5�(�f�n![����Ji)!7"bN:�DB���[u��7�� .�\���7�{i�����xB��T�,����n++Lţ�;��5���2���pƥ�د�Ɇu�?�3��q���.�h�u���(\46@�8X�G�k�$�y/��a���K̊��J��r��Hz9�y�l؃�wv��e��q���ݝ�nL�m8ܘ�9Jf,\�%G�+���)��\�|[��B�qpK�1I��i�E@�3uӤ�/�Tkc�'���~Fbӏ���j���P>7՞ Z)�q������&V�GT�SfkDpkE9�	.�Og���T�p���!�1����b�b��l�moBY�1Dm[�=�	��I��өp�E�Ӛ�A��UB�k	7*d	r��$�D�Ts��QT�qRH��/�Kߦ����=N$�6�%��w�lrJ�d�}خ	�;����t-Hc�<hz8���a��0,��Q��Y�d9���	�&�ʚ!�L/���3(�d�;:Q�A��̽����,���]HsӏZ�ZS'2Q��ѽ+>!w!g�}[�5�SBWD[�*����}G����h�UhH2֘������;��4����7/�-kwx�/���N[��H)5��gj����_�5�dv8�.x��l�X��}G�~3�׿�[]i����4��xEz����S�i/}SFt�>o��:�yD^4��^!�2�H�z�|� jR��2�?���	�����Z+�3a��2f�
�׍�Cc��O��sh���AfՙHhR��?��EP��ڱP�Z�l��䏧�Gu��>/hL6X-���cjt��'}�٠U��"�s��ܸPҋ�'��o����t���t�"P��Jbi �������(:;L��';U��c�-��2��.�8~�T=Ὂ���E������;��Ѧ��b����=�����VM-��x�{[�Շ�d%+9�c�[Jۉ�_�����@�ǀ��D�����:SC��wHz�mX	k��Z����R�e�Y��G5X�I��(�D�#�Bf �!sc��d��Q��%�]�z/����,�+���Q2��B?�d=&#X�S� �Tʀ,�(9���(�[�ON��=;1{�G7��R�`5�/g�J�2�if�r����¿��.y���s���>��tǲ$1�2�=Ϙw�R��b� R�ka���\�����jϰցÊplQq�؁?��Plުx���̎i���ח�1��XŕM�淓}I�7�f�s��/���JDgC���b0b8(!��s�5Z�/@_"����Aގ��mOc��zA
=ݾ[��{qٵ,T��߰�1	o �%��|B��F���xs̋���4
����g6m%
����O������d�A�˦��4��<�H��r9	�q�D�}0�r��#��s�&���i=�%���>!/>)'�<b��QMuVQ��l����l)@�"65��:4g�Y��I�B�h�y0(Z�4tw��G��������r�b>�)*]Dै�!'�xs����Q�3-ܪ��r� �R�K��.N��o���[����){������:����m�����	s�B��0�Y�=B{��I��΂xڦ_����)�"�G�
�9��-��{^q���jD0隒�^�7&�V�\V��d�°��ar�?��̲ڍJm�g�g.o�q�yL):(I�+�s�[~�2%[<�+3��ݶi���� �����A���xc�`u���$�}1U��:rT�ߦ�
��F�l8v���Cs�b���j�ؐ�0Y G�a��]N�T��~ l��	�)!�d���M��۝{a�Ԉ]�d�V�fm��I�d/ݼ�r��6�;"�J8U���-N��[��-�����n4��#�����t�d���$Z���)3�g��C�|�[fI�bF� ���Xj07�B�θ���� �K�����"��%��hiz}���785ak!ǝ��0
m/�U��L����V���b�w6�:�voҫ!��j/ɑy�En&a\�蝘�:�'^v��b?y�RU	�Ȋ�����<֞�rѬ���(�k?�u����|�n��[�B�"�m�B��з�3p�/��2�&җL��p�O 0���[����
�I8�sT��G�������_,��b��}�[A����ŷ���3C	�����8̏�J��F���O�{n����5)��.&�x��^�����S$�v�B��W(��G��p��Xtz:�	��=��NNI�����d�k���3���Њ>�9ȓ���e��'ʢ�&S���K��A��Jޏ���x�
�{�K������.�g��4泖�0`u�d��'I0�nbő�u�9M@f�P��<��t�M���.)��Q��O׵�m5?Z��]�)}�&^�.�2�� ˝�h�̭��>�P�d��}�6��@?-�K�쟴U��IGl��+���\�<!�Һ9L��6q!� =n�B���$z�Z�k$q�V�-+�l���k�e]d�A�NAu	�i�d)CZ��"��^�tg�~�O�J8h~Ҏ����M�$�p�P��Ad}�lMNl�����ͭ��T*q���I}�T�؃k���M��]�!Ŏ]�=�������cAʷ饁���ECK�̡Ċ�ҊUsQ�UM$�abx�oG��<�t>W�I9���-�q$6ǝ��vF�"B8��@f���q{��L��)�=+F���P���p��y�����x,\��ū�[�8}���,��mE�ߑ܄t��?j��'�űSd��{��y_y��x��2|���5��}=��uxy΍�RKY���/��n1�l\ՐP���,��R�27�}w�'*.��Md:|B�	�N�H��*��<��"�i����1�$�*f`�S�Kƶ4�L׌�gp�u�2�������7t�l�v鑰�D�GM!���T^��(�:U� +-JJ�ur_?�3 ���W{��)�m� �;�@b�덮w�
­��t� ���8c6��*Լ���H�<���[�J�L���rw�1�4��c��N<{YM��ɂ�\�G�������~$d�w2��1�����.1��uK)��	m����1��3o?�Ɖ{l�1�T=_:}�w>��G?��[�'|@�O� �lU��̮��3�؜S�B�֯�X����C<�qޗj~�"�t'����\�s�r�&�%�QJJ�W�#��j���h@�]��7��&N�e��@IP�i#W��t/[��{Pi����3	MǬ�y�9j�N�=��&��G��?b��3�����|��������܁S���T�����=�b$(�c�<�k�4Z�:��`+�C�0�A֨T���@
{25��փ2q�@��U�%[�iG�P����#�X�V�Ƥ/��������ټ��,v�|R��pT� "�G����]��(�kL)��1�����E�+Yv��L�M�[�S�PXM��p(*������I�*�,�ق#u�%�#}���z5���+��R�'���Rr�W\:$ι-��[�1�F֑��%��
�$2ej�#���)^P�� �8��my	�ƿ��dN��Y��qX|��/f%�7��Y1�豼�G���W��<�j�ס���ude�
: �����%��OΆ*]�V�j:nz��?)Ɵf�B���=�[e�^�ȣ;�@c�P���?��$v�=ڼ�@s�0 ��9�9pW�e��7NM�����m��b���w����E�::�9�D5��R�m����LȄ��E�RJ����+Sq1�{�����]zg��'jq�!���գx�l�ȧϔӜr�Q��C8�!�=dU���x��c�_��t&��N��i�o�7gρbx�QS�8�����N[1T ~ʘiۅ6��Է\�s���/��4%�^���B�n���T*g�`�N`�8I�c7�( < ��Rs9�NYbb[�x��P�\R�b!����<�E���.'�JL��E�(�;=�>�\�q�/����p��Ĺ�FcDݗ��b�N2 �]� (���DZ�Of��IN#"�ڲpT��_1*le{-fU����q%N�ư7+�l�ZW�*�'l��,�4��i�7��8��i���Q`Ί���[������-5>dX�I��u��u���Un�ץ^�ʶك�/��{Q��f�b�kԣ�JX�@��;��蠶&DvW�` ӾjPu����\�L�Q��;�Ь�&��g2D�g���,2��JM�}����lI�QM����.88C�k��Q'+����}B*ӣ\^}��u�_Kc�������b�+��� �=��r�¤�Ι.�@#���Sn���?��7�A���,Vm�� ���3�zR ��B��1��L}���	|p]�{l��)h�nq�3!uً�,��i�����l��n�!�F���~������b�����@�[�=�����!qG�,9��Y�H@Ɖ�B&��ĩ��٦��\t���V�wo��2�yA	��Ԧ��w����xT=���B�L@}�:>�_Q:c�#X���+�$�;Y�N`$V*��(i/�O_���$d��¥����i|��n�_����0?�G�U�z�F��`0�y��[�`�/���|��GT/�9D�9��JJ�GY��L7�����S�n	Q@*t0���l�ӷ�Ԣ�U�� @��y�h��G��ڃ䱕̻�FlZ�h�&���Y� n�v�z�t��@3�Ŕ���9�2w��Н�L��ρ��d�+ ��x�Hv�	���K"f�2gY�*�wI�^갑 8@#0;+�j� v���r�5�r>	{���V	�L�t/w�- e�G�����ko�j�:T	}�v�Q��+vcx@�?�n#���D��BR�R�I�9rP܆f�u�Չ�o:Y���q��Be+��1X�$8������v����l�
��+ ����!�<"��:�
�G����5����Q���R���?�)-���Ȇ���(���&�����@���K!~��]Br���2K�����:�Fz��7%���כ�(�G"$�
��ߙe��v!tu!�IV�B�������z��a�0��	�@$�����U��?�E	�] �H�WE`��%G铔�f��a@yJ��䃸+`H���x�����7�7��p�t���%��3���}Ot��j�#�D�B��c�H�ni�������6��;H�m7�r6\��wOI�/�ؔ�t��ɔ2!�CΨ,�(�L\�/\�je�lu��C�U�V44�ǃY�W����ڻ<o���?=��~��Q�׾�@��k�w�O���b5��+<۳r��0��C/��$+��x�)?�#���f��%a�f7V�bI���4Q�8'�;���̋b�C��>�q>�rL�j�O������c���3���Xe,��"��&GOg*�ú-��.Z�y6N���d��h��h�+ 2h�ƍi9d����+	�Mr��gӀ�>;�����z������x��� E�?~Ἕ�cCxFҲ:��yj^����	a��_8�_�9���໼�*�q!\���5����}J$˺m	t�:�(2�1�&C1mK[�����1�T\��)��nӹ���㠝K�����yĥ���G)�w��2��$Q���{���z��Y�㊕W��P�7@*O�ݯ�8I!{�pQ<��^��N���$�B����M�`m��jy�� ��!��R�p裧�zJ���LF�][i��������lZ[��O.l�*�Ct��:�ш�`1��� Z�0�M�:���DF[�UQ�܂`!O*���Qt7W O\���C�[�4�UaR�v����a�ezN����<m��媩q�Z�A��=�P�h��`�Wܻ_��[3��^��<��KL��/���D�Ty[rE�*�������`��q�iA��1^ڋ��CB�I*�-��m�c'/�H�|e���W[%Yl�)�S��Z�@���1�U�;aɷEb}}�R�T���G�.�0I?��m���t&~�>�g��݀z�F(��Йz������Mb�I���Ps�qP�'�~m���7�����2�y���M

��Ss�q����CX	������iG)��e�1{�g@��W_�����OV�e-�ϦS.����L��9�'7��d�v%�����
ȬR�z�/�C/�}����[fw�:�R�(���p.�ˍh+�z��=�㐙�TЧ��9��@8���pg
d��?���(EꞠ�8���n�)733����!����6ߡ��J&��][������<�sp���X�0����fQ�m�1ƺ��}�6�D�qvai�����N
��?m��(B����l>A��ZJ�=��V��U�[�����
�+u��y��ސ5&���]/� ��8E#�K!P������?Wb�6�/*��5���w�d���Aa�\�Zٲ�X�.��eDF-S9.u*��cQkI�\8_���u6h�M�����>e�a�Z�~<Ii0�0߰3��z��=�KJ�Y���A��q���KaEa]d��������N�!W+i;����K=4��jG���~�S�܉V��2�x�}��K�(o���2=�������/e/8R��}MX�/�����w�j/Jd
?�Ak�ʘ�)GD��B���
�F��dB���]cӟ�ļ���x&�{}i���Q[΂�ג�� !]��M�KXV[W�E^x$J�*�*�e��@��A��ȝ�zq��V|u��D�[�!n�V��lr ��Sz.��%(`��ᨙ������2_U����o��M
�5��ڐ֦d�Q5c�|ۜpM2{x(1�B˛'�D2�*|`3����+ǾJp3"��/�u;�:Щ9^��뙔����
���=�ʈ�kU�Yeo�׿���I��&ؓ%�+Ja~�6�nD8	����N�����B(�������R�p���k/�k<̶-=��+��������Y*�k&�G��%Y��h�+������`<b��"�-7���Gr�v!M2o}u#e����<b4m�j0G�@�C�̤�G�r]��)�s�ý�����3�e�~-�x��h�z��䡌��ۊ�n���F�ـs�.T�o�����1�Ɂ�O8Ӣ6�e[����i9p?�?��1��b�o�?��o�n�u6*����D�E��3�J9��I#��jZ�ۖ�����6��q��y�,Ne�	4f[K� ���<��n�IR����@h�>���O�e�p�����VG�=���Ȥ��\|��ņJ��NXS�����G�Mӆb��$Q��~�ݶ��'������&�b&�.�������*5.�����:��z҃F�մS0�A-��yL�'+��D[�9M�ӹ��2`�r��˖
]6����0$%xz����2�j�����~f��2�-��i���|b�á�E����"���r�%٩�X��'�$�������d��S���5!�g)��8|q�Ȝ�������i��;rq��G�hL���r���I>�pŌ3̓G���`�}-+Z�?�6��"�2�0�3���.�S�L�d �[֭V�ތ4m	�b�ăF'�C�m���,���S�άo���MP��ȭ��}-�bg�E���,�&ƭ>���@S�qN���a1���ݹ;����?�����<;�xY�J��4Îx���B��Q'�31;��p�:��][�%{͂�f�L���}-И!��p��'�͟�Z��z*r����h�� ҙ`�H$�$�,ɯ��5�� ���t�:����ai�mF���-�B�Y}�ܪ�Vk�9�)�^z�����E��KkH�2+jP�4���^IR��D����~�u_����ǂٓ`xb�M
��$Ev6�����N��=�����L.>�
0₷
4n�)�@�TgTp&9���uE�T%Mk �V����d?^q�x�x�Ԛ����S�X���bYR1�eW0qH��ݠeZ��<΄�/9��i��%A����+��$k�۳C5�Y�*5���]u�����l�X�p���B?��t)v��H�'�"l�g��z�lM��w�/*��:�<��!z��{����㘅�>��&}#��v��'-����)�/�N�~j��z�3��e �4�z��K��k(�{����v�����}������R���Ҥ���K��8�oh�������e$���y�PZ�o���p�gG��xO�0OG�ĵ;�6�TL���Z���gecq?���̝�/�)d+�N$N��/�%�A�v�M4[�ڄ� �k�u�Ҥ�C"��M̗����+h|p ߒ�2���HC�1/p���-���.F��i7�s�()8�	�������A���ay�2ϋm�O���|���P@��{?�<�����#��w��].�˪���q�zC8'��.���H޳�Ҿa�$��8���u2&��i�h��LcZ���I!xZ8�ӣ�@��V�2Բ�r�=���ӵ��F��Bр�Iv& #p`�/U�L�o~�f���ω1�\ 	��7�l�M ��^��Ӳ$h
�&#i{�+2DH���Vp8!�YQx���V�W��_�o�ݶ��4�_!!i�ӪkF6������bw0]���(M��jl�1w�-�N����f Xd���(��g��C?Ԣ�=c���d�C�v����4W2ɽ~k$���g�D�Ţ�9����_�+�FfH�&�M�8�c���� }���p�"���gˡN����лw
�>����s�=�OS�Fu�bkE���fT��Qo��aX��2���8�����/��\�
]r@��"��s{Q:��P[�Y`0�1���F�����r�h��Y� ��2.|��턴4�}@i��L�;�C�R8�T"(e'��gJm%IrD�!S�v-�D�P�k�+���)0����nd��8$I�*s���m@�~��@t�QϮ���ț�-�>e$�43�.�$*��e՛�������������ϧ���x `�L&hU�9�iI+:3�z�uVQ!a��z���z�"Ya���{�R�F�6�=�.�4?���Z���Q�{�~�_�udmwkf���ϰzaɴ���g�w�L:�ǜ��v��V�+�|#�E#�p���l���Ҵ���7�����aҏ���/��� �\�kS��+�`�Cp븕emg���]�@&�=#��JR@���lg"	�|�vkz��Ւ�9�D�P�<hꎿ�� �� ˅l��Iz��	\���V�䡐$��\Ѓ�t}%v�˚/.�n'��G� }&E�w�Y�=�u�jњ��,������L�f ��s���4��t� �S����]�<�	(Xv~ƹ������
�x�
W�ʋd���mgP���:�%A���&�.�����9��S�SӶ�	�!):��vx��E[�+?�{��6A�
8����GL��~�X"P�������^	�-���@b�T����U�m%�-��'�MC��A�9h��3�n}�۶�-PA�K����2������I�n�O�_��M�M�1��,�	U�UX���w=�6�U�˾����:���<�EMU�r'Z�Eʆ���ަi܍P�M�f�cXA�}��������/v���k�?CTթ�#�3�t�׋/ֳ�"௥�AI��雱�M 麤�..rf%�쓺j5�z���e�n�
89���:9���W�i-&O��wܲ�f�$��zî4Q`~�Xo�
g���-�P�q�_��$��W�E:����#_�	绪������e��C����,���Q���}g�T����Sdí)orm���!�I�^\eۑ&*����R�%�b��S��ox�)�����L�}:��)I��!�Q��oQ��Q��C.�}�A�p���\��jS��9�da��C�/۽Ah:�%��6L/�mi�%��v�d�֙i�'�{��[����Sy�K�sd�,X��K���m�A�*Nዐ&�%n�Od�e.���Z���,�.������VH��7o�O�����[�N��e�н�,u�Ϩa�V��Dv�*�?��潭�A�;_%�O,�K����@~�."Z5��Ǭ��≠x�������c�4�Q��N�Ǥ�H��(�](�Z��}��VA9h%٬���Tb��q����œ�ɓq��:]��T��7�-��m����ăA�����4G駖V��x<�~[�(�|��1��Kl��R{��P���_R�}Yxu���me�\/�hwرW�gl/1/t-���u�'\�)�{����z �����݁�?�|;��r�7�-;Xz��a,P��M��/v=B�!�Bo���pDr�E�N�a���g���{�����U���V�*_n'�ܓ�?�@���5�h9HXa#��Ӆ�h��}o*��_�����\rM,�jG���k�Tk'��t2�ڕ�'���4]����Ő^F�Ge�������j�� N#�x"�ܜ&�e�ޙ�[z���o�Cz�&
=O�ڪ�鱊܂P�q��������T)J'���^���nQ��7|'�@��mqa�W#?C��:����&����둖����n�%.����F�Bt'X&���{*ιQ�tUӌg�>j:�o��e"{�DP�����������AɪM��b�ٴ��N���pzbJ�&R�h�Zr�#N�H�k7M�.;T��j����,=E��X��<6��Z� �S���׭܇Л�[�8�*��į���^YD����gG���;�:A*��߾�aP��vH�R��0����h�����%���Q�WUb��]��?�;���D2 ���<~5M�P�Qv���2�!J��S�.�o��"�#��q�Z8��8M�Ͼ\��wK׎<�EVJw���4Ō;l g���Úbn#�Ҡ='�[�������G �x��:������X&��_�a5���?G$άhya�hni�q3v��f���-��z~���N�=]�c�˲�e`X���̈́��BVH ����GH�w󮵟b����f��8N(���l]lft`�KNGˁ�ԎA;�
�8/*R�^"�ؑ�UoJ��QL�.�*g3d�H�!tܗ�Z�|Oj���D�>�P;��Գt{��w�ͱ,O��[`ԃL`gI4d��Ti��&���1�%��
��6��f�������L9�%�T)\3nU��-+xs�t���J�_�dY���T���pQ���F�Yt���zZ)���	�^�r�����d��h© �c�)�&5��������z���5	i���8o��1Gf]����*6��5�1��y"�&��PD�yu�3{���u�pi�8Uo=,
u���r��ٳ�����Ǻ1?X(�� �axO�)�����b��u�*Yy	j���ՈZ
�ɿ�յ����v��:K��G�4|Z�W�`�y�V�� Rc��Z���V�|?���Q�y�aA���\ha�L͹�h���?k��F�D�P�>J�����uaiД�����Z����J�"�5���z쭄�$�E��wCO�|�;��s�U�ܧ��J�^4��@Z3k�R���Vg]L�gU!��Qx�#ܨ���GN��[h:��<�e��dW)��sW!hd�����?Zz���-%�
�^�3�h���p��h�&Ă�SP}8Q��R\�w,������hunR|"�b�Y����w�W���?�hj"�;tB������y��<"�u��V"����gij��RD"�z��H�,�q΢��~ڍ�9D�9p���%��{\-5z���t}J/�4hv#,�n��uG���I&f�-��H�
�e����(>�=g|�tB1����KNCʬS?âp�p��P6<|=%際�@�~S�5��-����6��{�+���˴è�*���M��F��vSh翽��>|����~�%v�^�����_i�#[ni%�W��R��jd��p2��l۶k:?V�"���)D�w+zǅ���"gh�$Gq}�<��M�C�Q�%x��>Xk��i$.�H>��+¨��@
��u3�����q9j��
Z��	\�緖�eh���'5�L�jI<%Q����d�z	��2k�s/��8�.t��b*�]?�F���-̣ᐖ'[�{��ʖ���D�o�#$���ܠ5P��'l�C.C+��Zr���+�m�b���:C�g���)����ý&�p��Ć�Jfu58�["�:\�B�_L'���iE���� �񩷟�I�9�/�ŇOu��L�+�jf����zʁ��~�.�%tG�t��J�� OP���,������WEU{�PA����	EU�Ǣ��`e#�m�v��������1����1DhE���4-�Bjϒ��^7�$)a\��p��D<�"�R���篇�snMH;w�(���Bqk��4���x1�Կ�&��3��%�����]Y��ꪸ@�j�`ZvA{E03�d����ΝnzW�������_ V�-��R�-���u��D��E�N�O����l��X�!G� �9D�Rl�t9�$Eee"�9���v���
�#��pV�oX	������/eb�p�i���FA�ã(�:_��;����e5����ǼF̿T]o�q��ϯW��Y�o`\�W��*���qY����{s3}vQ��y�T�ɿ��^J����$��}̓�a��I�U���ʡ��6�I�(91��.[�+NOJ��@�	f.qSb�x#/>4q ����+�D�I��D���N/��	Š_Ց�b)I������d ��QV����|x1����D�;�b#p�&�a"�.h�Y�4z���l
�\<�{����3��kTgn���Fxu��Փ����5��Ȭ�\�H�Lޞ�<������Y;�!uC~¶��w��:���1&6b��,�ɡv�*9��G�v	��T����8�ێ���Z(;��p4
R�B�>ɔ��Hh�$�y$�WW��SI�S���Ps�ڠ��r�D4A�K��e/ Ll҈2�����8wi��|;���g�]r�<�MUؗpa�W��&3f�%�S��l�Od���Ƈ�D*pتj�&�"wt�K�t�mvc��8̛�4�;�[}���f�*>��e^�5�
w6�ᾆ�˼��UYv��I�������F�i~�����Y%���؇������4�������F���[^_��A pzAA��=@�=�t�Ƞ}�,�$(�}�;��X�N���m�_��!QnB�e|L��+��.�w�wY !ߞ��k�����$:>����^�R�-��h@Ɍ^^.F�@t��њU�-�t$@BYV��Ը"�I�Xsz#��k]ɉ��|�l
��ˇ�U]�{/>��:?�[�_�5�Ծf�^�8<�o8�U�A��щa	.5V���B�q��QaB�7��&�,œ׃�ǖN�\
mn:�C/�����E��B���bv5�����V�;4�mUu�
�X,$@ݢE<g#T����*q�@�Br���H	�LY�������۲�����oLm�A�*��ё7n8�</���4`�\�f�M֖~���H����@Z��w�r�4��������g(��~�<�>��;��LS7Tg�>�\mϤY�����$��7���G� gg�;��N
��k��Y���q�#��G��F��.v���ċ�0Ϳ��@2��u0�(����	�_�@�#A����@�1��- �����"��~�z|����u�*.{a=\�+��qE���������mV0����B�ɲ�iw��Ȃc+��_5�F��p����l�M�-
������� ���E��ݯ�_%�0�I�=9ѭz�@#Q��tp��l�r����Z ���0p_��wY𘓏k�%d@%��E~=�lv��)��u��=P5�Ͱ�S\�V��EY�c���w}�������p��"��|Ġ�=L���Ky�}�m�{�T�Sp�t�V�côY�
ʊ!���[��H�9��ۨaXG�|t{�Ԭ�|Tc���,%5�ДV� w�5D�gO�u�ьB�����|*�w��:�m�wX�۸\�y���F�(���%x�H|ne�&�k�����PBS�=FFC�/f�����m�_�l;�X�9խ��w����*�z�����iUf�ƙ��,U)�<��)��&ӝ�C
����Z�j��|�dU:�'c���ed�3-%mq9q<8K�x[��`���9K8�Z��q�/'�B��� ���.��:���O����%��@q[$����5���"��M��f	QY�%ǽD���O##=�qE�d�`�~���E�XVJkk�w ������%�:�ֱ���n����lg��0v�Cj%%2(���!s���?����+���0�T�W�U UC��l2N����}R���7t�� `�0`lw��i��@�#��6L�h�$�0u�A
ܹ�m��h��͐߯PiZ��˥���%�O�9dD/����_���8�)$�KO|q}Y�@�������'U+��Q��H��������}�Ұ�L��N(Sބm= ��%	M�Gņ"2���F�����zw�A]�-��ʐPGO1��z�� ��r�\\_�-z�[n��>6T�m�~H�|�1*�޸���@��i�垗8����d�7��*~|������1����L��k��3.6n�<Ze)k��c��'u&~	�ĩ�~w��O6=�&���}�-�y�-k/�0��q�����8i���iG�Q�'d��9pk���wο{4��E�<Q6�%�k�сYI�2751��v[:n��aJ/�S�k��Ƽ�oy(����Y��&�����ۺ*��kT6�-Iw������}"R�R���#�Kc���*���l��-��y9��'o��Y(;��y��`CO_w�7�D>�I�th��r��t���W��&u?u9샰�%���l!��
�x��[I��P)9D�Z���r��:��Np���3�H�q��Q+��?3���n�jrev�j -�g�I'd�t���~P|`i�r�otwTV\�c���+b�-���i'>�37F9�����T� *`�}j��g�}
O�b]��H3x�U+xR����q��'Y��L��(�XJ�6I���Fm�����"���n'�Ï&��C��ϿJ9���\栠�4Q�h�s�$��)�7pRʢ ��'��M�6���t������u�=0��7��q]~4���5IB^�^dB���nU
�1iE=�� ����
�ӆ��˯5�)6 N�U
g\��8I�����/=�Z��OQ�|N��n�?g��`p��i�y/­]���y�� v0����"�G��	�� |3w�&е�xB�2�-NĶ���$W��qt�l,s��MbRZ����
��S��kRĜ�RK�������WK�׆��)�[�|��	�Lњ֨��$@+nK��mSg��
�s�x}6�Iq˄��v�Sh���B��q������Py�ϒ7�8],r�*�>*���������C�T�3���y������8����G�&̲�-S�^����\�8��|�Y������C�	��q�k8��0'g� � K��V�z�x��r0mjS!��+��g��o���������L<{�և����L�yv�aŝf�9����������L=�.j894����ߌl܈�����S�����ـ����o��~vt�wOJ�l'CKJ�O�}����]>���$�U�*�0�B8ܬC���P*��:��5�c�T��zؠ�5������L�M-�εY����)��O�@tJ�	l�|�xr�A�7\I�Q2��;;d؋�Ӄ��~_09� �J��� 
�b�!�Ѥ-��t_��51[)K:F�t�,�8[�[C���T�q�4߽�\�ȿY����6L�q��z���,�^�����'�#l������ÇD�2K�į,�b<_��|�n�򀟾ԭO���k5�߫!x���`7� �Ӡn�����2ʪ�pȂ͉�5aOw~�-�"Ф)������=�����Ҕ㎷��7,����~^Ov}�ԥ��-å�b���#�0x�-W܎9�����f\_R��X�L���� ���B?���j�(��T�z����g�f�N]�rtj��tH�� �hb��6���q�q��}��O�?��J�e����,����R��a���J��i-� �V�>��@[E�SnY�b�g	dF튶 i�A>��einX���6vO:�pݺu5����
}�`J�.���%j���|�,Zt��W4@<�a?�8N���G����{�m�Od�=���Q4� �*4[ȔHGH�4)��zZPćwP�Q�fh
i�S�W�����H����:��fA�O��}?ؐ�lή�د���1��'�3�䋢A���#��i��<��M�8R�ٯ*J��Z)"㐵4XDbb^��"et�ஈ�9\��mb�bk�#��+޽�š9��a��-@u�(G�Ula����ܽ������<I[�%���᎕��}�@_8�O-O��s�q�2 LԆG�]��c�q��+j/O�ږ�0��l����Q+�gR�Ǳ��f4y���ք$�?�T��+�K7s���/�>��q��P��M��^�y���2]oFه��H�yR0|�j޿B��ٞ&I�Ca�m\�(�ww*�Y��B�M��z6���t�1q�Fn9����jvFO�ȒB���:< ���3<Po�ϱ!Z�A6	f�Y:1"�uP��c�����v�.�Dz��9 !£�� ����,����z���5��Y-�������{��R��5p�7���ê��O	���?�@���A�h�Ί0��(*6>��+=WNWHڏ=�L�m4,N��'
�K�ⳂE�R�L��A���z>Kk����6��}t](��i����t�� �X�8`�k��ru9zp�T/�s%q��I�~��g�q� �V��ADx����i����
�Ti��~�q�ˋ�����j�I��(8�?�m�Z'��!�k^�^a,\.y�"��xM� �y(�Of���ZDe�'Mx�0���<�z��@�]Ly�@mC�̂�o�jeHFL�X�n�S���;��i��-W�lCyQ"�b�a�p�z3��W�*��m��j&Gd0˖*��HX�Q����(ǷV5�+���-)[�#^ZRIc{@D�wbz);��6�(
�~�h��e���VW��=���n#G"��R�\J�˖�������0Y�@#����iRr����7�s#��t�2���U�m�$x�v�]�Q#�K�*��癝l����I4.�n��3��Q;D?}R^�ܟ,��<b�`�Be͑#X� ��nd��Ӄ���#��43�Y���޳U0$����+<I�?1��v��K%E���vl� u��}�����H������"2E10�.Qs5�W�:�z����X�K@q(Ĕv����ý����r�Þ�8)���s��_��g�M��=�YS=�W)ʢ�f59����#[8/h�Ƌ�ǫ~9��`P	��8���>U�l$�/7s-fTp���E������|�I-�e�`���,=3�7�M�~Cy�Բ����T��|ct?&�e̸pa���/>�x9�B5��a����h��gԷG?`��T��xX ��YuA�G�3�-u Q:�N�99��Wyi|[��fzvP�q#�T�lu�?쎕_M����:E�.I,�2F:���O��E��%�)s��A�����Q�~ ���ē�Ը�	�:��O9��%:�e�E9�O&n4�/Щz���\�F	R���<�"?�^c0X���/���O*�����ќ"�`z�<ۍElH�T;ε:⓾� ����yۗbu�>�k=	���Pe$��\ti%�'IК���GѴ';e?x��|S�r64�֪?v%�p�M���E�?�ٮ�6�b���l���^H���+YEl��n��5�d.��|0��a�U�T�V"��S�VV��F�s�5�Ӣ�c⢭�5�͘MJ���w:B��6A,�G���.$ܓ�2�v/�g�әK�,�\�;��[&� +�~���BHQ�	<C22Q����O�G��O\���&�^Gɔlmk}�LK��#�.�����������*�FG��]��`��)�M0\l��8�,I��W�6� ��^��+�S���T��YPm��M@�h·e��Pc��}��#���[틞
E1��x�/�f�r%�ۧg�l}}�?bwG�fIMm4��#U���?�/⚀�qK#��g��_'w���$��B|�|V"������.Qw�I:ڟ�%_ڠ��	��9��n����G��˲";t��t�e ���0�9��Āv��C]HNs�����[n#�M�	�9!�2Ȼ��E���M�QZ0r��]���!��6+�(�äA��X��������Z ��r7ծa����F��cRS�;l����^_�0	>�:�A8�{(>��U���M�"�(�5mB0���y�3����KX?��4@Tg�ŗ�����,�I��Q���e��7ޛ�1D�����r_�[I��@��\5l!�Q�pT�u��Ξ��3�kj��fU�2�u4[b5�����-ٳT�<�#d$qF�/Zs�V&�5���Q��?�VU��)v���.�Ƹv�XnA|<\����EY�Q&�J�]N��B��Q��7�"�T9��(9a�3.k1�����J�e�'7�qؚR(�Ar�X�H_$��*.�ɀR�fe$¡��dcIE�O+IL_߈\c���Q����	]�+��-��kW.�Ե���P�mMy	L
U	�o"<��m���������̸�o��1;�����[(�Џ�&���wDf2p��:o�4ό�(��!݅t&�kRе�*���>�}�,8�Z��q�S��<��s�B��xوК	牿j\Th�ᩓt�|�z���4����6J�%�`��A��w,�� p��!�P��T������:]Ѹ��>��\T�h����f�cI�N�ƹ��Ɉ��-hk� ��<�c�/B,d����ª�;N�Mt/_�h�nҼm���0f6����h<Π���g:V?�}�&���͞efp�7�����|�8b�,��(g���FII�i/��SVWf�,�J���6���>��c�;�N���`����x׫�n�� �yG���N�N��\�'i�d�\�C���� c���ɂ�|dy.@�h��<�c�1�ʮ������?iR�}�Q����lr?����"���p@�Ϧ:xT� Bg���2�3˞����(es���Z���A��1���J���*�L/�럏��Ȏ�b��3{�����^z���q5�T��%������ZI�^�k���X�<�$Z㆏�2�3���Me	`Ѽ��h��U'k8#����g?�=m�¹x���]�?�{6��7x���;Z�H�Ĕ`������v꭭����h���0^�1�,�\�L1��j�<�z�K].��%���\���먜���fVs�䔂�n� g�#�8�gB1ϮIW�<^���PX\�u�ڭ_�8�!A^{\�C���6����yf�X���QW�E�F��G�fܷ����xrw�u*� ~^�PgE�i���o*��;������ |gK��s�T ��74�W"���P:�h��UQ?�اҍ��������qG�>��4O�OWښJr�7�����#�0ۧ=�F�A�PE�/��NCY�����9C@���6j���.[�3�-a5��z+NO���̓4�KS������Tv:�(JF�3S#��F5�>Pb�x�dmi�T�kv|-�o���-����u�[+krE��a P��O�<0�7�׭�	��������x_��!�.5����]�S$��S^�Y���:$��vk4C
��ɺ/]Q_$;!�x�Ū�ϔTzĩ��?�0�j���1�"�Q?��Z6�(���P��g�":����r���C2���[L���=iK`,}+y�y�è�@�E)$������$0)�<5N�V����N$��M
6����x��0��a�?S����[c�g琇��ι<ة$e+ٝ��r��
�3v�(U�O�!���;����s���wM1��$^��ڮZNU�c^�`p����Yd�$�Y��7�,���|������~�@xH��*f�3�^�,��e-��{�? d�86x�.�x�f����m���Gx��S=�֨k��b�lI�
�
CG�q|��!�Ƈ�6<�?>fsm�CP�9W��g��M[����R[tD�"r"%N ���k����K�:&� �DeF*`��~����������0�4��������\�v��]�	3��R��_�&V��F�\�*�Q�s��%å��������3�'��cyJN�Ȟ�J����Ti�6)8�Z*���EBו3�E8�<���TD�K�^g��Z!�X/��zݻ�ks� �s�C#�3q�"0y"Zln��qg�[�zG?"��Z��7^�鲹���M���f����ɀ�{^Q��Ʈ�>��{�EC~F#��R�&��I��>)�Qs���K"��	&�!�1!C�`J��\?N
��k x��~��Ɍ����G�d]����-+'�@���?+|�/}v�"�4p�5���k�=徎B��)T�ܸ愸�|�*�M4����!U��)���$FX��uیŚgVt�(ʣ���)m&��9����<LY��h!b&+��A�L�$�F�9RK��g1sC�`��s�_�f`�J�:eO�H�2I+���\�Ա�~�ۄ끡0���{TVA�0���qB2�V��K�0mV�r��#в�1���%}k|�E��I��Kz�Mz4��쐖�r�c�Ps�[��5[O��e��ܨ��� !6�S��P�X����*a�̘��.�>g���m\&�I����j��[�	@jM�Q3[H��^�]��DH�j6���~�˞�OW`����.���S��9�y%��s���sĦb��Sr�xs�v��qð�	���D�B���M�D��Єm*,�n�nN� �3���N��٢����Z�t\j�X��Z���
WWw|g7B�Gg��Y]�]��ܾӸp�󼟲�_�)��a�?�5p��6Bo�&d�fgЈz�_U�Ĕ0�����]�3'/�5�V�q?d��=pV�u��x�!��kUlD��p+g����L9"-�z�{�|��6�h!jJPa��m}@@p��Po�f�/;�
��z��1�G��yϔ�d3a*���`��k�����n���0��@�n�D4`*Tn��.	a�06-c�"h�Yp���8�~�&kg��w��@��$6�1���k�Y���/0���9�j���=Z�0ڒ���6ċE��t���˱��94-PC[4�n�Bs�����D{�艃U;�����ыq2�mi�t��g�CiOdG���=��oBl,����)0z�/��<ޘ �o}�� 
^�S��n\��=t�tA��_�)��.�0kSޏ��q�� dw�I���]���I��6�x���De�&����������tq�����t#����↡����a���L�,�:���4�NT0&n��5�:�6�����f�+�~_�:+U�ިC�{K������a�!�B�s'"{��zލ�������r�A��6]p�)#H7.Y���8�Ԟ�y*/,ꌯ\ ���n����b7����P�������u�G��ڙ�[-"% ��ϫ�_���$�x:�/R��]5y���`���=m��% �b�ٰx#:F�+�n�+�	���$���D1�lׯg4-���x%7ygq��Uuu%B�P5����N��)3�h)=��6a�)�n�7%eV(���9h��G=��FT�pS�M�?�K3��fH=N�9��^�9�WǊ����:*�vc�7�*|�u zT�7����bYk�׬�4��2��1Kn�Y�Qv���
g4u7�y=ݵ%���Q���7�@��Y��e�`��u���nF&"�����fD��e��y���+m)�흿��D#2��S���(��L�w(0��ۂQ�7I���^����[��%<'�solm��؂���E�to����l$[.x����o�˳��eUE��Z�kq��{�pޞ4��7�b`h�Vk+T��׭f���A�쇰����UK���1'E�2X�g�L��1��]3O���
jO��9�/���_1��Ր�^y��j~7�܎��(|��!��V%/��>��7��ą��W���b�
ʵh�[�2��m �����t���@F��G����6���׶���m]����g��A�8�0��Q��S+�9�~֙�9����J�~��>�
|�� oVğzv�[I��"
$���f����c��ڲX�~�3}�1�ɤ�G���g<��y���z�Yɸ���=�c�����2��R�|��?�Fw�ՕX��+�d�������E�1=DR����Ѧ�j�&f��0�F��_}���{��}V<YS�_�ꤔƬ-J#P��=��eJ������l��r5+ܯ���C{��t|��5����;�Ԯ�|wĎ�jA?Z	]���!-�V5|d[}tI��)�$���h�>X����V�����l��v�%��p5�p��+(G�yoQR����{� ��T1,0�)�$L3����%f�(4rt��Vv%��GJ��Il��x��%��4�5=,�~,�գE�7�'���ʹ�$�G{jL���Jr/(��}Ҟ�rm�M����}8��Rgf���_��z$0���&&(���	���O�Rͨո7�P�'+&+�򩚘VN˴�T�L�w)j �����Z��Ӿ�:Ҵҟ�TNJuTv�M��@ڌ��R�[/���A�/��%�D�R�|�c����e��Sz�>�����|sQ����el$A���#���V;)��a��z�_o�dts�s8�S|���=d4�$�p��D H�1ROU��[��x��1�J�kq`��S&��8�������w���Þ��$��_щ9q�]����qmp�M.�𨺋�[��i�>��8Z�F+�������p?�m�X?p����rW�����@��=���C0u�0ju�pgC*�?�a��X�;������O}�	4�菁���%�ppZ�.r�Z?ZNλ>9�'���Wf�ҘS�
�z�]��^'���v�3�8f���}��<�Ľ�&�ZQT��l��C�!�Y"#��B�=s�R�2��Zc�+�������f$�>b_=4�^�*A�UG���奟�.����.��6o����va�1ױ��=B��jh�2���	J��A[��M����X�٦$���n�¤�4��s����{����u����a��]u��D�fN��q�js	���cz|^	��5�9+)�xc%x�!�Wb�ǐaS��aLRHp���>����P�2<��-��:����.�'�p�x$D�D��"�Oױ2����-q�,n���vނ`�+��sF|P�P��{4:A{PZe5�9�;q��5=R��j~��jُ��^-��v	�ŭM�VH��g���nt�zu��V*J�#p��Y�;�3�B8/�g<�o�yt���ʦ��֏��fׯ��"u�$��2I�r����N�f�MRpE�7����b�Ĳ5+*Ǯ��d� $1a2G�1x�kW�v�[^g��y;y,7����zhȯ�O�G�:~��t� 5$֓���Z�L��0�)��-2ˆ��DW����	�IGh�����M��[���0!3��픑T�x碒(�l_Ġ@#�>J��E<HM��w���Qׄ�t���b_��l�D��Dai���'W ٬�9��8�XxFËY�\4�̯��\~�	�Rd49����m�q�bhFr}�@�ڳ����T)��&vVZ�F_�;����+<��#W�J��z��G��'��w�������r�Rkh�/mrP�O�
iZ�	cOJ�S@�u�A���:"˾N��3�"�?�;$�O�Cֲ��3�����tS�~`Jr���Y+�ٕS���C3,�K"[s��X4�^/���A�2퍭�:���Wu��L�v��z�C�z>�R���o#tb���2��_咬��(*�����^�<ty��Y�o�tc����K��(#1Y^�f��m�݋[�OA��+l0�n�7&	��ۓ1aF�4��JY)5��
]ʑ�i��7��z?ц`Ys,B_��
^�( �'u�w����Y���$�|��#srL��[r�oǇ�_���K�d��Yr�?�����BT��I0n\?�E�`^�`!��q
~�pdN�g�[�F�mD��V���w�*�l�[�}�[3p�s�w9��Rt�x��o��q�u&y!�m�Ⱦ����!'�5Bo��8nG�w�,���T��4|�sH�� 8���+*��"�"�T���u�2�d�*5�T�O|��Χr�C,^�ьnb/�;�L)�O�U�V��rįqT������L��<!]�7"c:
iMe+�φ�i�14 ��')�i�\���yc��uV�����  ���� ����������h�h� ���R4Q&�y4��,�]n� �#^3����K���(�(�!�Yl��,�u���],&�)p���j��o��Z�6xt9ڠoꗥe��#�9�����7���� 1�q	����a�=�]��}�ԃ|
Kϧ�������F�l2�>G�;����y���߈f�ݩW��c���5��_oH,䳜	jLug����n0��R�8�����J�����]��.��֮��6n�����v��w(ȍ�3%1Z�*Y����c�� Ó�5o���ޡ��([�jni�0�ݒ�9�R�� "s���{>q������y��[��4�$d�����K1G�"6�Ec$�y�J�Q�Kr%Z���-s�M�yN�Z�/tM!�޳
 c)�Ua��Yc�LL�i2K�V��U���~��p]��:��>�{f������.`z#�jW�[�J�*����D�i�޿�iO��[�U�G�ө�M�v��;<Y�{(�O ]���I�7B���K"�1u��P��	�;�4� \�a���	�/-!=d8�ຟz_��o���W���z�-M�I�a�*�2���էMOS�	9��i�V��
�Bf�aZ[�l�w���s��Hŀ��^��n�X!��a�m e蛻�U4`t��]i�m&��E�9��t��!�#�҂�`�e`>�ݼz��y�" o�f��E�R�Ap���9A��?���l���i�$��U��
�>g"wz����^��j�!%�@X��G��9�Z_�.��n���J�8;&-�|	C�:(��Cz��8�йχ��Or�����0
OK�*�0��ɚZ�ipĀ,�)���+������r���x�[qK��-�W��\�W��'g���6=d&*��+aW�Ƴ���I4 ��g���VJZx`d� N�z�k�b�r��b uc/��׀oq�`N�3/��ƩX(G���w�����o�&��E����vX��r�����E�����E����S�f~�B��D���j-S��Ěa˟�ˤWz��}�3{�Ʈ�Ls/�f<\S�~< �j+�w�T��hX�!@�*�m$����v<3�?6|�=a��H�a) �<�(E�\U� =��|�
�H7�x�S)�~�ϗ���9;6�ht�5��kt܉�7f��7�k�#���gN�"��P����"���=*6�J#jyJq������~[Ӑ��]�'��'>�='Z�3���n����*l��}�x�4�HՉZMs1�y5���ۻ��p�P�{�|�ϼKt;���O��inw9�v� �k��������[ЎQN�� �UK$L�5Cώ[q�	.d���'�:�2�Ǎ�?�t��A��{�i��o��yC_ϷW}��F��W�\#�G`.�h~�Rź�L�9�0E�3��L�V$���X��0,{�c���׵�J
���H�J�X����"X�KӖU��v���7�ot���9֛�7����H<JWn�_��J���֕Ʀg���gQw�v�	'�KZ��V/D-��Ax#�����t��<ڜ�y�Riƥ���.K17�P��z��ܲF�CŒ�8��A���|��̾oM�oY\B6p��A��Qu?�kSYר�g]v���}�I��~	�9	 �I'L'�������YD�h��w�z7�S]V��Ub�)��J�뵔f������ �=T'&FL����(ɤ%(@T�۫���J�N��:�@�MI]ð_���)-�IǒE�Αu�������O�ʔ�����-����	k��\"�����˾���I}��<G}���9��-�_�����U��W����#��D��7��6��/�E|c�}��o�j��I�6FSe�xx l?�`�}���V"z�`��=�#��E��~K}�	��>P)���=����)�N
0]7������> g&�T����=��vv;�7P��{�&ն��x pB�[��<b`��M�h}�i�Ì�V=n��n��PS_�����T�ch� (�-w6"h�Oyh H>��~�k�Ny1	YCvsD��A��x=��=��$���}`�-������(n���Ѱ��w�&M���'yy��[kB�Ó:�.�_����5�S�z�9V�^~�GQ2C�'��r?G�e�,��vy���q����'����[�p����ص��m��Qg�C���{jO I81��!H?^ާ���0���N����2z�H�]��[�
+���5�/S-|EB�J�>���Q+ӯ����d3'�S|�N�e���\�Ϥ�oy��<�%8�W�7�����E[-�.�p8{8���r-���M8h;�zn�uȢb��������He����+�`�s�u�
��t�dr^B"` ���O��\�8��q�I�:om�D�!-�c,7�Ƙ��.�Å���F�A�n�D��}��<��j0"�뻸��kUh2+��P?)�(�Q��.�7�g�~�\T��*}����%�=�(�'sm�$)�O�"��qb\��'�̘��6��c��5p0u_D�`����S�<��텂��N��^_�8��?�e�Xbesen��$'�lJ؏Z�B�u_��Fd|`�!|Jj�KP׈H.�_\Ш�c� P�#�iV5���}����2p@j\���fA��h24�/T�\��,��ے�)��0�Cn'~��՝�0V�[�e���[n]a	�t�A5"eqr���/�m,�J,��5K$k��aY��dQe�B�P�
�繲�Iŀ�fg��k7��9}b�Xr��t�DA+@M"M�x��l<�b���&�<�(�:Tϑ˫8
�K���M�s�;�12hI��)��&y��Gu�H�z|zMaw[R�aq��y��JhQ�J`��~A��^�X2�h��k6y]@
x�"K�����G���=Rl��%�b�v{�p%��OL�wy���j3��ϛͷeg���pK͍H���)��@��4��-��jԫ;iKQ�rXd�t-����������a�T�q���dT{��+{f�%���W�Y�C�HL�c����hj���9��(����(���k�^y���4�Z�^(E��R�T+iYP�ΛN~ �?���ls�g2�}CfJh�~Q�\�I���L1��_Ӟ��eA��W�p׀F��W�ǅ?��ڄ��gSikC�P�!�I�w�䥊����t-`/x7h�c��t�m�������$m�n��ӂ1�ɭ��o-RwTo7��Y��>Y cJ�	�8)�#w��)��_�jg�*������> v�{����ťO��J͎�UQn
O������/c*�&���H��u�}x�����حK��du�!���x�Y���QPH�Xg}�%݀H��mٱ%�� L�����zI�LN^��uvE����<�e>�5Gy"����J��p�̍dW�Ԙv^�R ,D��P�'Z���ǡ�)���-l�.�5�2I��k?\����{P�0beR�Gmѩ	�C�]�&B�`Xh����^�b� ��U�ym{ee���L�n�6mbo#b��Pu%��9_P�G6ٻ�h�p���d�0�:�:HK������1�]�o�~:�R�A����`��/,�2 s�$ծo�	 ?��S/��ܿ1�g|W�٘g���K`u�Wa�T���u��l>�Ģ�4�/D8k� �w�R�����yY�����n�6S9B����p��^���N�Qu洄��g,���"t�s=���S;����Ͳ9�>�jY7N�-?�7U��"s���6�;���.`�K��o�E���7�7t
�<[#l��Y��$�.�|j��� fW:ڨ���!&�?���I�G4�w��{91�������Vums�'�ed�/s2�y�m��X����V��PE �^�|m��&>ױU�F{���SV,�d��k�5�k�R:�f����E옝e�e�n�8�ص|�qd�êՃ��҆�J�� m����v#l��e*���+�g�qP��
�?�`���/�n �I(�+�fa�δ�ˡH4��+]��8�>�T�����X�`��^TT@`Eo_�:�)F)���ȥ�2\�����с�-�+���H�hh�g�÷*��A�^��[qDw����#m���qBX<���a☧$x��M�M�6:f���-}���i	D&��#kԈ��Ȃ�?L8���;g�j�'h�y[�<�u�����ڂb�����H�9_}����Ɵ��P�Z�;�e��L��W��:����X��b,ߞE���c�Z�q+�g�vܱ�/.�PE��m���"49-x�Z�q$I���>� �Ql�o���j1�|*��#=�%ˬ؀�=G�J��<��i'��g��)�g�����\�M�I���4���-��� ri���V�t�E�	U�1���;�{���?+����UZS��]�ap����$2��7��DT�OՄ[���ᬉ��S��^Ht�$�^��m�vt+DaI�3dA08\��xok�ݶC[��A�a"Ҍ�:��pyN".�Hm,ë�[�K�A̱XV�j2��|T�6Z��}����:�������3OkT���7&am���y�HCo7��x��<:F[��r�t^Y�f=5��#���a�$�2F�=?8f&{��4P�?f�7��!�]e�����N�z�:�NY�.L/X�{��>��U%yY3��&Z�{ -�|n�V�m��1!�b�g�k�ɘA�%~ث�3��'�r>�z�U�߇�m ��y�G<����[U�w�2�����݋���|l��`�c����#Y7k�6�5�ʀ���������m|�R�SOcd�O���J�e��7��$�ݩ���t�(��J��4���fA�
|î����w�G�36�d�3��o׈tȞ�u�ʖK�p�[�����X�0�ܦ���^ح�%����+<[�ZR�`���lҌizY���i\��n��C:�'�7Z54A�o+�������J�tg&��vb VTF�T��-6v+J�>X<���W�����J��^
�M+�	n�'�!~br&\�N�v�5���I	�6~��*P:b(��K�&�h{�b��"҂�G�6�M��e�`�ǜ��Մ�m1e{������,�[�Q�r�]�����7�{����|��, ����j<>��p�Bvh���'�����-tl�� -��0{tN���j��@0�[�3YLٮ���Y#;��^��%��+���/����qh��N�C�2U����}�	=�m�����2}\��V����B)���zJ���S�Ÿt1<OO���j�c��(J"S�GK�;+���5$?�m% ��o��\�f�H7[!yĖ��z��'��ј{��ڂ}��9���6Ĵ��dR0���b\Ոe�5�c�P���;�����M��|+؞ {u������X�����x�;� n�*�֦J^�p��v�Q���;5���<�tұm%B��@�pV#}���'\o�;�`ǀ��M����C�t��0F~j��w�7��'q�:��>|~�r*Ő��0���j�d���i�]2?R����މ_�q"�Ŝ���pй�J��;��� �����B�Q�24J�z�Რ�6�=B�P\m���'^�۟�'J���k�dوx�Bs�m�+�[LC������Z�X�i�C����1i3'����N�pV?�G�C84�:сB�g3��>��8�ܪܣ׽�6������*�GD�-���3��z�`��M;�6��Q`��@'v�΃|M���i�Z�݌�T���`��N�[���\�BqYc?�5�U���&��IOU|�j����(��0W��1�^�#Wv %eY�bg������vR��������n���O�N�O������﷒��kN��>˛i0|�ԋ�"'W8��9�%A���%1¿~U��fb��Z�Q�"���V����&�U,�ğ�ǆ/��j�f������D����P`~,eY����X�A?�͝>�����A{��
�����F��i��a����B-XT�г�@%:*�f~P\�S��r`��:� ��"S}�n85gLzX��0�h^���WD�B��R�׋�#Gf'VCz=@��@Ja6�!r�Ak���Ck$���Q��LГ�R�H�,={�~96����^Cex��*9ޣ&~����u�"�Ĭ�I�|3b?{���_tN��xb�Ć�t�h#RRRŷS������q-@�}�׻}k�N���{�(�5+���*:����� 4\;�9��Jg���A�՟�j�!�D�"���k��H!޸v��Fq��-��p�~�ҿ���1r��^�u�����Y��0G:lA5�l��P���"cTz�{���������.�j8��	��U�`\�Y���Dޤ��ױ�Gk�"�RL�o�g����9��N@��g��|���kx���E
�q,NEl�v���X {�=�zc��p�A�ɘ*$��Tm�q:k�.2�Gl�J�x�WH�/���1��ezE�( �6�3a~!O�=$�	P����P�E�G���nu�ط�g�6m�w�?��[�)���iQ�bڻq�+�s���g����'(.�����Q��X�V�C%-|SO��'c y'~.�	1���������}�(�?��GGyb@��+12�c��hM�u��d
�ݧ���NT!q7�+i>�	_#�B5Ջ�7����7����u�'��h��lRۂ����0U�
֣�q�Ǣ�NR���B����>�Zn�{��
�P`h��9%�!�L:�4�{�&��e��m��蘅0H������k���0���\�i	���*�TF0�^�zk-r��!i�;F姕�{�$+-"�Jhz�0�,f�J4�<�KL�-�Y}������m@��7j{X�5�0�w�g��5:"���TV�E*$@O}Nٳ�Ɲ���U*�k������5�~s�O@�z|�6j���#�a�Gi{�"5��,��Z.����pg��W�\b)9�R!n&"H�ȖO]��)�ť�����v ���>�R�h!�sC�G��)�E@�ǚ����k#9����D���dX������Q�c�j�k��]�=`��b(0/-���r�C��QE!��!.�VC2|{��B�1o�lP^�9�O�����]'iu�)� �����, ��G� tJP$(��t
t��qK���8љ+�G4����8�ػ�D�(H���>�M5��t ���p6|\�2�܄R@&�r6A9�G�DIn��U#/��������;jb>6�>��o���&�����i)�3?6%3P���M**T�����u�2�Lf3^���	VlI��iT�>a��:%��ySl��]M4�bn�����=�:��	8V��1\�|1[��?�
���󺜡h�9;/������Mb�m�2O�S)���=��lV��� �+��vF�����,�+619__,x������\�i}���h9�|#��v��ep4ld�l=p�y�E��zN�ѣW-Hmu���>r�`,{u��&#�g��Mw�ڲY�d��gd��pe��{Z��)h���Y�����S6�s6XQU�^/��lp1q����/�m��T(����{p8���J1+I�H��I��OPFc���S�{܅�g~z�jGXvR�J[y����Ql��C���#^��Wy9�`<��-��A��!�Z}�o�5�}���٢�L��F�<����,���8<?�G_�@H)�R!���)6[~ށ�&�d���1��5� !.!��8�e�:2����<pC��g�(��/�(�d�������<֛�� ����q��L�L����CƻcÔm^R��mCG�^]��ڊ��q�U�[����?G����-�č�R�''T�C4j����8�4+ȝ2���H��:L:�[��%v�,� fO�HMX��)/�ژ#��6u���B*)$[7���tzI]uh��V�̓��m�p�v�;����](
����Ia)$�d�x?�5�[��!��˷U��XI�g������Z��e)����\�����D�`]�b�dCL���(�rx�(r]�C�Ԏ�w{<�62)�Қ�<|�@�0,vRw�}g�R��N}��DOx'u~GH�vk9-#�3}X[]�̲!�?��~e��������X���p�����r��1��#�[�a��@W�ITj�4R|��ˋ��V��Wyc��JJ\��qM�����c����Ok���uo�]�W��:�7]ğ�g�&Ry�d𱖦�i1�#�?�`�5/(0S�οErO�4@��`y!���(�~ßoٗ'���V9^���e��`H��t?��&����
nH�s8V^
[�0��ĳ j��"X��|�I�<8İ��l��%�����ҁF3�/���5TAO6�W�_m:*!9�I��բ\�BV!�Q�
�T��,;ˈu��jRYIg<��$��8�A�bWzSC9)2*T��1���3���!�	c���&8�X0I(�8��<}No�W�u��-֓H}/�IѲ���V,�y8��E<�W��|5�-�V`��[�yZ7w)J�=�S��`���ܡ]��i����`�K8:��\0��=Y�~��)
��^&B2�s+��H<�Lrr����<�DN��M�<pQ��������.��+�����*#I>�1v�	���L�,���e�*�&�#$��+�."���:I���B�F�y/u0���{���� ԕP��X!��[��@��X�a���.��puĝ�ߩ$6ɥ3u��Y��W������r}��p��)c3���i��g�~��r�D�B�5מq�5��Y�u'���i�$��=U�̣�"����栛�|a�HH��x5��6��1���o��,�Fle�o���{��(ƁjLqP:v�WS �(mj��`M�>�5��'�o�F�g��RO�ASs~'� ���@cg�����0�&�]۩�7�e�eĊ�0Y���P���D�q��w[&��\��m����V۱����R:�Ĩ)�9Ng��B�Ӝa�𾹵���G5f;������~�o�R#��&�2,�=Jm
�i|�I�oy���յU���VG���e����7Ib!��'2뱞��;io1c�F�2�v��h�[&DY]�OD��N�J�?R.N��N�5$��|sh}c��"�=�m�(g99�������:X�4���#/HH��Z|܃7?AI��`�a���_z�iS��+y^U@` �|��D���s�8���^Q��W���T(����^����´�+�o@gVu���EY��F��w���(Ŵ���a��͘q���S�1�	�:�W����F���t�2T���qh�����%n������Tc���Q{9�]@��m��fz�L�w��C>��ݜv���!����gcl��Y-X�'�Z�����ym�ǘo��*}�����3�%��ӗ�m��r|�2�)2�7�J����4��=+�K�^jD�v�2�?���N�A�.W��D����l%8��0%���L�!GT�"� ��E?��C�L�ߪ��&��|X��wM�w�s�ȼ��ه�)�~��x�8Լ�HH�mg:���b���
����S�U�8Ϭ7��[o�Z�I#��cd��@G٫Ӷ~���Sʈ�9���µ�L�'�����U�v,�QUݙd�fɴ�:Ё��W��]M������|͗j��,�n��������*����)%^_���qʋ�%���[�s���t�o>ڿ���QO�A<\`.�Q�H�4wd>(�!��*C��FJ�e�������V�p@�L��\��%��GӛW����g F��&f٬#.���|���vC�:�	��� �����מ��{���T� �_��A�ɪ܂HJ@[� �	&mұ���L�d�������U��t%��-䱿T��'����(Q遉�dR��Q>i(�]#	l�[��!t�pԯ����_L�@vb� ��B~>���ϩ ��9	sdt��4EP��W:
�G*
��4"��t�H� J��6����H��U|Ӎ�c��J�L����X��	R
�sx���b�{V#L[J~s&���%`B�Z%��9l��q	��̵ 3�n{��ְ����� C�ڍ=	��(k�K�ڙ�r�Z��mR@�W�~�r�w�������fp2p8������@{���'�G�Gv���� ��p�M]KQ^}�Û�;��1�̎����O�RWfx�v����ߢPA�#xGr��	��ͱ!��#�u�ם�7���j(���3ͭ��K��@�T���]*��k��ۺω�iP���G�4�\O�����s墵ǒ�3�F��@�?����UՕ�8�k�L�!�����4���g+� "m2�E��j�yp��X/[�j3Y�"D�J�(K��a��Vf�}	�#��w������l[&�DH�
�r9	��.��r�CP�x���o;e�� ���L=��CP}�&����b
E9�A����X�f��4����\}}Q+�d_��_�DI'��F�!�]�O�}��g#(��9�~�u��.j���%_T��6�嬒m��u�1�|�u�����M<�g����8���
�m;I����l~"P�f�ZM$�(M�a&.�Y��8�����ɯJ
���a��k��������ř�G�L�����4I��Y�z#+.��<�6�e�#�B�,��l[wYx���x�������X��S ��O�\J�(>)JY\��$�/���ه��������H�V~�^��,�5N?��){Ŭ���RW���P� _J�kJ��OOw��!� ��J�Q�O��X��4�?> w[��!�7�M�\�Yv��V~���_*�b4P��<�t���=4��e�f6��g�3��K��5��O"�_j���;�\Ńr���m���}a���73eN&���P@�ke�	���am�q�q޺fRN	��$P�U?L�y�Ԩ �+������=�[�S���S�}���g{cV]�1�tOGE�f����=ݩɮ�ñ!?����g]�g�A�	�7����|a���2���Ç<Φ��֫.k��!F��1���&��Bg޹��/;�٠Ě��|����
e� Y'��Z{��T���/�{{2$��X������Z5�OHZ����{���-�����'{���~��޽�?��9����!"'7޺�'�����M]�`�X滎�'��)�dsp�$��Dl)�������{�пY\q���AAg�=Ӯ��Ye8�,G�V��]�/q�����C��`,+N�AG���R����)6"~P]S����&��l�fG�Hև��[�{^3�5>�;�~�0TI���A�i�T�U;�����+�_�D�A���(�:1��j�}NoJ,x���$�;V��y�G5\������rۿ�*��ɷ*	Ä���7n̋�u�{��%D<c#�x��V�I�RيF-ps�%��xn(bV�}�П���W@gxB�@b�ü˯al��|�J�fA(1`�R���<I�@,���3N�O�ޠU^rU��,M�Nٌ'�In���W5-67*@7�����JB�����I�6���\	�9��w�$E~	B����)�3�� �ݴ��_,:�s�7��⟿ʸ'Vu�R��[8��C0`8�\B�G��~
&8��*7$EyHb�_K^�Q��Sl�>�����ڒ#+��S9rIps� 1I�s�fGŐ�M��)*�I�9�'U0�:�J�7�3�Ok�V����l��.�ҴH� A�u�Ơ�h
IV��8#�(���Ge�YKoa!7i[=�(-9�}�|7���L�JNm1"�铘�C�+wI�R�Ρ\����~��dg4��Fz�  #�>����}�&M,��)�+�	��a<��r�(����|�}��y�Y��g�[�:M�����n
��ޏ��wK��K�"�̐c0�}	:샺"N��U���8���z���\�r��\�!2��Tǀ�n���r}V��D�҉S	ύ�!%:yېW��8��ELgz�8W#��#�=r7R㺙�Qb'�r6�(5��_��D��A3}KQA�"�	<t]��H-uE�dM�:�x��ͻ�>0�����7A/�P�Ԅ�J�]^�%�:|%|uZzqu ƍ��8Ή���P	p���O�ۑ�h�A��PDF��l	3��5�R�'\�e��ceh� ��B"oF��wm����E�g��9�'�L����fg�
l�Ǡ^�t���w;*��5�w��=s�ͣ^�g�a�|-�{=���7�R�
\�{���nC���7	�@�q���$:�����]��Nh�չV����W�0���x.�q�3]�7q?=ꁧ�X�
��&^1�����5~\�>�z(�v��X��,�|"�<��Z]76�F����P��aDޠʦ#p�QC��uV0� -�����L_���v�4�4l�F��_a��`͊�Z��KcҊ3^���/��Zx��Y:�o9c�pl��G��{=$��j8���:�z�i����P�Uu��h�����B��9�6w�P����H��(@��?:uAB�����x?H��e�ι���#�#��d�J��7��1R����l&�?��q����S�V�!y��9�Jox��ɰp�	��({;�h)($Pܰ$�X����1I���&�p�6z�61	���ɟ$�<�۵B��`Ԝ�����̷��N�Y��Ռ���0	V�I��7w�Z_^��m��DM��:d� l��L���P�nMQ�Ɵ�,E�����uv�t�����d��X*$f�mұk�"����v�BI�)>�gPڊ\�Țt�4>@��t;�W�v�Kw��4��V٪�K?�55H3>��_1C�=<�����L��*�=hnH}._��B+�ntT$f��ڬ<�u�&N��?�x�2�3�2�_�	���:ys'�?t�6�2ྪH=��R*@��8r,k�I� s�9â�$����l@��7��^΋���W2�*�>�Hi�8�#+hϘ���ݰ��k��yK�����~ol��[h��� X���u������/�xc�dtGyE�蟵�9_ʹgdI�VMug���
Ǯ/�����Hw�+��o,4?ĝd{���D��n���L��] �T�eO�a��{Ӊ�1>iȈRK�=>�vv��L:�����
(��@-)��vU���+(��,9dӹ�B,����f�c��3	��ʷ�jafum.H��

�	��Jg���|��G�v��js�E3�Q����6u�������"��c�:�g[��J4�W��Й�)F����;��>5
k��xE�ܮshf߷{ц�=9~D��dZ-�Y��������'�pc߆�,���W�񬄉�կ짂_�V��IC"�7Q�A��Q� im'.,���/ 'X���X�V��l���߾1
6��%wlϤ����hb�vjt���}AQ;�d= Q���&��dU�<��e��ҞQ�~��)���t��a�*�_Ue�s*@�y�Z���?)M7���j!Hj>���j���p���j{�]D-�k�9ȉcM��X�� c&zl�4p��"��F���ŝ)���ьVH�-l����S�S���ז�Br��	4�J��K�����C	7]/5Z���=í�V?�h{�;l�kfko�0CZ:�t�B���PC	
j`1kn�s�^����	y�V!=��[��(T�e0��!m���'e`��^s�T^Zγz��oq���:D��ۍ�MB4�G%K��I�=�K��H6��*���gF�?�1��.4I��|�m�o1$D�\���h�C�l"��jɈ|���fbC��!r�a�`��@��0�߇5��(	cfv����/��=oW?[���2p��t'�wd�g��;8G���97	���QBI����\�k|����J�0/ҞI�_8�C��~�'Ԅ�4���a.����,�,P��κ���C�|�w#�r����6bmI*��G7s�aE�qD��<ꈇE�wR�Z�U�Ҡq�ܜ��ϴ%u��I�C�"ړ�k�.w��'$ᚳ1 s�� �h�ͬb�������|gː���|��m������XW��jb�|i��
��~Z��2��M��u.`Q �@c�*�M�[%�./=�\|t��z���9^��M�Z�vY�L-���������e�.ǡ9Ȓ=5W�	4m�=6���S4�ff&0���������C�f9F~�Ŧc�wj���U��`�#���p%��!�[1k?�P"R$�w"�)��jt��1�+�:㊁�³�����!$1�_]�x_�Z*M�Rm�vQ�����2�I-kT^���^������.���Ta������8�j�g��Q��&����3�e={ɴQ��o��refQ�C4�+[��'��%�Z�m��J_�hq�E���3��,fAF�4�%��;�;�g���
c��8�&�A�.����@B�F�گ�Bq�UHk���
J��w�DȵKW�qN,B�����	a� ���*�<��Z}%����?��T��ŕ�?���,h�t��\m3��RR=B\�g5Rp��ޜ�>uҡo����ey%������TJS]	����0W6S�Qϛ%���-I!u5�c�S�܆�����q�~�j�v�r�2#:��/<[�2���_�ۇ�ml-8ݣ�����.
?JX⍿����\-H��sp&8��4��
�!5�|�w�����L��L��a�1�Wԫ�rt��.� �������E���RX�m�Џᤐ����9>��\�� �:.Ԗ,"�[a����"a�P}Ȏ���������1����J�#�^T����.��\����O�@��X�9�"��6�����7!���K0h��gL�.�R	]�mo٢P�
�3�=�Ws��ɾ�+�UN]~�6�/��ģ�|���������y�U=�p��M�S]�;E_�;���
YJ��C�w~�뎧:���a!�0��"FF�;��8j�cO�T�6�Z�@�\��ҭ�4��'���0j~��l��I��4�/�A��c8%�;�b���0Lΰ�Y�mj��n��r0ׯ��x�-�wya�Zk�UG��ji.���G�ÒE� �z������Ga�<T��5�ߺ����f�D�
M,���;�@]�8�_�	Y��i\v���~r[�x�G�Uϔ��7�����_l�Z�U%^)��Q�Njx�0��������(#i�V��+1�%YX ��:���s6]� Z��T2�vJQ�N�{5E���; ������ˑb�k�:ay�!L���F��l��a�k0�_
-��73�D�$���8K��י/.S���0�/`���٣�� SMeM��e
4%gGT��@@*���P�{*��D����u/i�Iv��|��Wn�U���6�{�t�F�/�fõ�M	�`ї�W�~_�rēe>jѯ��~���A�X�����Q�ej�_L��>�Ț����]	�y4���������u�NO�ɸ��K�;��O ���2�W��Ċ_��+�-�ߏ2�bN������tfWv��D����ka�^��I���/r5�2F$oN6nˌ6�]�w��g��+�P������g�D'��͕%�D�en���_�I�nGs����	��f=�eT=��y!'��4Pbk�0g�+�2As��M>���:�hA[�S&��K=� .�f��e2X�>���vai�4���a*	ڙ3z���7��S~��F�+v�
T$!�v,�z?X�4�@�X�54:����1���#b��P1	� {�&4O�AnZj�@�_gY�:� �h1�Z���=��i���k�ni�-�O�;�z��7����ٞ�l��w�Nܢa��_ZX��+7/����4|��)^Bp @ O(�3��l��ҹ�I����a��3��镖
kF��U4 �W���f=� �о?ô,w�-Wގ��U.��Z]��7��v_E��nO��y#����UY�I!L��0���"��ǔO@D�V��S�Vti�l�wH�5��9�ր�������
�!�
�b_$��?4��o�V�͒+'S���	X�6��@8�q�0K�6�23�,��QD�Y�-sCn$B��tl��P�2ՙ���BX3�;G�̀1�7��^�W�_��N	?���'�
�x�B���,ȩ�C0������o�{y,��Տ�����dX��4cQL��K�O���c3�)��^kK���#���Ý=����ii*��3�����o������㠙�@}mPi�z�觟���JpX�����[���N]����7"���$�2ϙ�'�d멇�x"� t��i������&�mgȻ�i�P�����>W򔋾!�X������Id�M�{p�飷j_>�*��Mš�z$�-E&�^Ȧ�*JG��AE��$�g[�a�l���dA��+%���<�w8P��7�R���Px>�������X�������9��3Hw��ܦ�k1���[ه��l��1;�R1���I��v��T�_���r뻣���m���Q��V-lC��H,�z��� T��K����h�(��R�4љ�.}z�@ZZ�7@��I�_�%3��4�j~�E^�p�5����5�n�JS�I�q͢����"�|o[A�Z,��#ţ��gʄ+n	k<L�#��^2-(f�J!�ɺ v`��qn�B���dSN���Ҩ}�E#5�Q�zͻ�@�*�+3�0eΪ)��k��ag���C��1>��3�ƛ����tL_�:ݷh'mjddt&����4�$�����S�˝�K��9b�)
Ԡ�Z�z,n{S���@�Ɖ.�`�J.�H�)���yJ՗mFiFU�3EsUk��mzps��%�kO�z ۺ3�oȘ;�wV�X<w��H��p M�tNp�v�ګb�2�{�^ �xv"B
)�����n�jl��֋���HV�'#�= �8��uu�Z7)�{����(�db�(�A5q�%&��K�?9�d��OL���&�
�*]���Kd�<��b�"#d(��{G��향�ώ^�#j�M5򳩽��n7��҉�{Q�����:JS鐰�dُ��$"�׌�k�Q[����^�d�)�hv�,w��+Q!m�D�hC�(���J{���(%���N$6�S�f!�ࠒ��wX��o��j�c-1�ۣۨ4�"g-���2�m d�c%�:^�dE�X�h5>�Q��\���� ~���i."c���0�n��X)ww��i+*��h���S�v�4U��~��$���V��U(�z�!䮠yTO��g�歿��QHd� �#�-���>_�^�뇌��Rޤ/��/$D������l��9�uݸ�	4��E�}��6E�x�U.ZA"�g^!XP��6e�2���TE�	֝�����k���s��C�#{X~Ѣ?�o� �[f?�����
���=[]�uY�Y�>�#�u�ϵM2���(�Ń�8��J�B��C�Y�&��b*|l�[YS��;Өe��I���#%�̬~�VK(��8�F��!��O
�3 "����Ǒ�������!�A)�MZ�p��.���pB� J���G�{��Tr���
�������&�����+��'��c���*�����^�1�?-��C��:�tG�3�{��<�md�5k�#�+ց�O;rk�T��la�,}�}[�S�;E�ؚ�y�G��J��l�2�4Qv��!��{���{!s��Y���*��!�g�7:�Wԥ�vN�T�v����G'rP*u4�F+�n
4ߢ^+��eM��@~ҫ&�9�(�L�R꡹0����5En(R,T�����p��{q��g)aA�%-�	�BR� ��K�+�FJf�#}���NB��0h� G�%]f�ik�z�OV7:�<�r��e"j�y/�$jl�tj�06��m��ʞ18=��M�Fh	J�(b�󏌚���"/�c|��;iE�6��C*Wa���\����d�"ȚP$XO���t��f�9� �t�i揧���p�5o�\Qw�m��N�k���~͘�J���1�����vT[�H��K���x�"��'?wʧ���!x���.�������Cy�h/m��6�Qc���ܷE�`uI��A#���'h��#,�-��A��=����"B_$@»��&|^��a<H�#�y1)Zq�m��<^�#ۉ�c�?i��I��9>�]xF](Y?�ă���C���+�=5���_�r�֏�㜲�Ǟ���a�$�y�Ν'w���Ǹ=�t| �'(��+Ί��=`��#i�B��L'w���a�{����~s� �1�/ޝ�kԫn}�mS�}5X;3/;�O��.���۽h0_v�F/��ߤH�eM��l
�&���gY�7GQ1���J ��|�2G��4ޓ�&am�UV%�v��m^%�=�2<Ty���ϖf��?#X��1�X�ێ���89E���QvĖ:�a`��Vpax�=*����~���c�����fe��}"�X(��8����>���?�{,�&C�U��8��_���yA���ט5�:�)��b(c����[�4ق����G6�o�֡�}�ʟt�������:'�cX؏��I�bŅHPd�'�@�QC)S5����-�I�H�)3�!��x��(��RL| r>�?��cড���S&CP���|K	|S˒F��.4�:J,����5'��Di.����6�-�;�; ��([iUp��9uuJ��x�'�M�uu�Ao먡��	F.�B�tc�|�}_.[E�.Gw(��4gJ�6�M��J�t��I�>r�RC�!��g�d�)N��6lw{R��=���9(��R���K�Z��m�Š�?T��@s���է.�	iT7F�������h>�Ȋ�dȽ2N@�Q�aB�*I>�r������9��_Ǳ5�%8'�Ue�թ[d�3M*nX�W�����uV��� 45�Zݟ���n	���v��dM��s�f�'�x#;bcCKd �!�N/��������$|p���fa5�#c��u~�ATv���]�N�ß8}m�����Z�b�(�ͳ �Zd6Z�Ĭ���l�$M�����uS��(���mZ�����5�H�G�#A`У7"��	OeꛂϿ��A˽D߀c�$�[f���G|�!�ԧ0./�J�M��a�GO�_���˰�������QYkU3�nE���j�3��ۭ���ʋrMC�:�hp�zi�(*hk���WzYԹaSQ���yv>=t��D����(��e���;�� p=�PB7�\�Imt�B�5�<�c¡{��X�'6� Mk2z�������|�n ��&��`�<�4��s�{C�u�[b Ep���A�5^���w	L�ND��N%q��5&����'�$=�Ƅ��� ��𨒧�Xϵ9\�ez��;1���%$��2&�p��_G�P+��ߨp���%UT��/M��as�h{#�0����k�U����Dؘ�[�G�8(<n�U�uz�i�*rp����E��]c&�v�-���-l�p��ٺ�J�s��J����9IgZ��-Fz�b���@�WeS��+%�E�����I�k-U��L�����^Ґ��zbX"D-~)�!�!l�� }I5R=%�a�
�R!@W�d��d��>\=O�/s���y(eC����b׷c�E�H Mgz$d.��	K���Vb��?c�t#��;ś��#*|��)D������Ģl�-��OCF$t��2��N~Hl�w��,���O9�
�xy��4�,�ι��v��y �v�?�L�+M�@@�'T�c? ��R̭�fzD�+7ӓjq��G�r%"=�b�dU��|�R�_��%�1'L�Q�IcȘd�e�'iL�Y�u>=�=vH)�5S���������{�3�1K.ǳG꺹����%�|w��>M��h���v)�d ��<�ۯ����>F"2=�A(�L6�n^�����b�Z��U@[��Ų��:Ѿ�Z��u�u:v��&��U�5���2抢��*�/2���)��TOO`1�!�喳o�
�����tm�N�$惩2zӋR9P��~�����g��Ec]*7tv�,|��3z��m��~�6�O31{�8�mX��,?�'#&Q;�z�7`8�~!�*�/x�p|!'�@k��/�Ҋ��0�(��!܆�EB�1\V�>h5n�7��.%����t���RѾr��bʑ���8ԿQ���w�=ש�Oa��9�[��l��O.��eHߛN��GU��Zg��6Msm%x�y��gK��q
�bf��l�?���HJ�k�5��?Y�kT���F�����^8d'bt�Ql9�r(�����v	=x��+,ifC��p��>��I�`r���c��6�ZڈҠ�M�T�O�rȺPo�3z�>a���r��π��S��C܊)A�?�tk�k�v��`�<�`���JV.�xX�KҰ�7:�~�zG���%l6z`���q������L��I�07"�- �|�	���?-��#�.��I�C�ܮ����>����%}C�\�B��*9�Z�gP���@^W�.U����{[vw���X���8ͬ��<�@;<Ca������Q����z��m)�D'�A�%�4��"��;e'�)���<(�W��ˎJ��_��i�.Vm0T��}&���U��'�W�C����t�.=���O�L�$4��k?f�I\�_%��͖i�	��X@{Y?5ϪY�����m��/+B���Yp<D1w�)k~I��N�f1G���.���Y���w���${,a�&d���ᚒ�\K]�c
�R�"�����W��L���~ɷ��EpզB���E�d�#l��¨ި�'�3-�S��a'��1�1�~.�` �#l�Uf���r��Et�N�9����D�u�2$�sK)j��X�dy��1s��:-X>cg�抂1�	�|b|��f��F�{�-��	7	l#:	5���1do���JJB�L���u��'���2K�� �Kh�z�,T���uT��Tr���%� R�$�|�$Gտ>keьfL�nӍ�(PXi�^v�*�x��h�Ѐ|J]J�����`����Z+�cPAS�!�0N�,����a�Њ�D;�9����~�L)�*;z!Dٔ^͜I���}TfyF��Q�BvR_,9������w|=���d�QX`�`-N8
�)���d�U���P-Tp"�&=�&QU�-a�]�&kL ��N��`5;?0+�M���w%Ȃ��iE�Q��;���?�"�R�S��:�z^��W=!�x�����鎑u ��lB���h?�ޟ���:�2�ٳ� ?VJ����eVQ��)u �!p��]ɮ!�R�ec�J�U��J�inf�-�'����ei�&�5o��V\��'��!�w��W�Z�X��u��F�g_�bM�<�ڲ_׻c�Z
�GZ��{J�Om�sO��x���R;[�4��U.܁�Gsע�(��V�u�"���g��f�>C�Ҽ���ۍG%��D��+�/����N�]?	�����gO�o<� ��P��8�F7���N����g[�x��hP6���+�U�Dd��k�֖�^�8��`�:�cv�x���Jo��?o�5Eg��n�v�ɀW<_�n��Ϝ����S��7VJ2�Ǐ��~YF;�����QC�&Ӥgi��������Es�%ߑ{ڶ(m_��S�,�X�1��%*qE@ӎG�;Wy-#Q����׈�~��l���� !��-�3����-̰�Ѹ�bŘCO�Z�υ����T3���A�m
�ү0{s�b�r1��0S��+z�tV�e�,~c�락&�Z��^�X��HWh^U�p��_�+9'τ����+Z ͦS�	���*t��0U[)N�I��-��?.=�kb���F.��)���&u���B�^�m�����c�z��Q�1�gD�vGp͏���"�~����|��47,��v�����#Gࡇ����^|̤e�Y[]����
���eu �b-p�\ʝ��$�P:^�+g�hb�<��X�]'Rv���d�^7�����`B�(��d�:�"	S�PV�r�V�7 ���}���<E�����lW**4p�j�qj%��^��Ǭ8���w�)`�o��K{��$ŷQ!��W�x�,D��A�Ӈv
v�`�XDğmH�ٴ�����x9��o�-��saNH}G7w�k(	1���J��y�]��}|mmVA"���,�'��.k��FjW�Cw%����$���/�WCr�pH�fV�I-�D�[�kO��s��፷�T�g�P҃��Q���j4�^qn�ǅ1��&s���7ŝ�|� t0�z���NI����m�n��|���{S��i��煘#���Ǻ��bەL�օ!�gm�b̚dvnP�Vסr:��D"�����B�<� _޼�=D$��&��y�a��1���ٴ��ϓ�\����� ���0�IP{J�"jiz��N;�*�#�嫹��0���j���?�*�
��֥�%ħ�2	s��z{C��D�����S/�|�P��`%���2�u�Z��irg@b����kce��K˵�q^_�-�߱Mc�j��Qη��}˴�_�w5���/l�U`��9ş$^׸��Sޗ�"��ƵuEx���9ín����=h<��m�
�S�����Q�~�����H�\ǻ�S����T�':��/M�z��V�{W��u�q���e\ny���Wn�{��
\�d%)a��jC�NE$шB9�-J��'+��a��>�ꬾs1�N�ģ��)CHÂӳ3m�jؤ~�7e������#�О�Yc&v���T�|[�]�bs8�Y,PlhL�u��pr�g�*�S��s(<vf�]�i<�Qn
�M>z�G��R�fy��Η�_;mh'�Aз�TW7��f_�e#.fձfo}��B�2@y� �Aji	u/��o[�1�mu�R�r[���,�� #|��n,_ʹ�v�C٤tl�9{����H�K��P���h1�%��n�⛂���Ix��
���\x��_]L�n���}�;�'�м������Oq�J,]�L{4����f�ғjfxǧ�Յ.rt$^���S%,-m֗u�{5,vəD�8�&Kgp6�"�X0)sM�k�[�_J~P��)��	��
�`��q���6K�A~	�,���G��r"˜}e�kt��?��C���f:A���-�C$	�iZ���'�ˈ�	��QwLs��E���1�ܑK1���,�:g�����赨����N��Z����A�]&�Ύ���oƘ$��6�#��"h��':]�xy�/^ĵ�;���2�F�㖠�!xwTާ��8����D�Kj+����
��.Xrq�~��S�C�KH(�LT?iA|���6�Oq�B�� WE�g���)�� ��e��{kz��
KH��A[L���1��a�L��&�5!�^К�S%��i��V��Xc������|�$���l@֤T(��D?�h�M���B�h�.%-��w�G�����7�o�� V�ȁ������Rbju��Mx����w=ӥ?�
��h��3�KmX�t�d�zs�5Տ3�2�?��
����ѶƗ�G%)>�X�!�?n���5�˵���L��)��ƺ�@�}ώ��wl�u�[񼶳v�o)���s��j�9|����)/��C� �t$;i��^�X�K�����Y�8���d����V��9�|�"�y���7bT7`ڼ42�� G�R:�{�����%%4i�Q�v�;�����`m�p�Y�w[$,/�2�U�P�s j���.�+���G���_���l���E�S�Qp�=�2�dF᧮�+��G�@ؗ΢�`��ع���Tq�|
/U&*+g���N@D_'���j��� �J��{pɤ~3P���F�}��4
�O1h�`:�2"P�ϝc�/����s���5�#ۅ�Y'�*�|�	3~X�=tggQ��vl��s�%� �-� #T:UPHT9��b�%�Ur�_1HAlB��<�~RP��4�v�?�U� Q(0T%���}�2�EpgM���&,QJ��4�y1Ў��*]<���8����Jlo�6-���N�u�g+d��لzG`yK�{l#� ��=Z�j�<oc�d����͠eS �(`���&��*4|�-��Z�����L����Gl:#^���;}�\4P�ZDe�SV�/�g�:�}�Ru�mZ�YUiN�=6ǽ��}���	%�V��D.�+�&��AXL�	�\�u� 
q[�.���Q�#��q�{�/H���g�0�l�yxA�LX��h����?TI���������r��a٧�%�Y�
���i1 �ȓt6��{��0E1~�5\��j!@�h~!|�,9��p%�?��WR�3���5��]R�ԙ����hFX��	��|�g�(�3� �<��Z��%�q�e�3H֥	��o
C��k=K=����8�aU���d�!Z�wYH7ݥ��L�M5�sB��'���T��ފ}�7gԇ�> a����T�Y:�w�H9����J�"�8X_z��͐�.�U�n�p�����2B��L��_�̍Q���sDFP��]��\��>��bi���@��47�I�\3�U����5�8�/���S������)�����n׼�h�B�}e+@�����.�����P,!˕i&L��Xov�>S�2l��ԓ�}�;�{�VH���+���{$=NP�g�`J�͸7���e�I*���A��|�^��#F��d{[��\�	E#��B�Mز�;�%'n�xh� k~�E��Y<a�c������8�5���EY�*���=���R���ç�q�7��z���|�8��(<]��G۲@�M?o�+�Z��Gd�E�h�d���Y���osS���1^=�P�1���;������~�7������;�J<XLhZw��f6c�L����퇛a:tm
:<�aB�0��r:���e�5J�$����v�3�Y
�&.�Q�A���qq�$�:��W�{�r�]�"K{���~H��+7w֟a��&v��)��y��Ɉ���~�9�y+���w�������q]�����8
}|,u"8��/Z�.��这xhӿ�*�K���|��[:i�9ܞ�B@��Ch]�X�:�&b���Ӳ�����k��?��x`4Vps�y�=���֫�̪FzX0�c�2"�d�X�Ϧ)�S�.2�r�{��r�uk��*C�0��A�5��l3n����"�r�����U�"�3��ڴ��)i��1�Q\�p���@|��;yMh���~1Q����vH�?cU��ю��͓�&��⁺���$�c ")m�i=yoM���_,�b�	�Q���n�,S���S<e�����O���+ú�?W��Gg�s˦#�M%�Ql���e
��8�Uy�a���g���&���П @3X��0�L�ݓ��F�;�^X�B�'��ᓐ�����.'JoC�$5J��Z |xG�l�!�q�1��Cば0�w��>%�z3������B���{>n�0!���\�
FP(&��r���K��4�Ө��V陁�4 A��ԍ�����z�9�~n�����d��	Rl,$B�[�ebv�SS�m�� &9E�4��P�G@�IbW �o�Wd?v����\BH#�VƑ���|��:��,���đr�ZxQxX���\�`��w�|�ϻ $�gCDa<��E����ԭ�W��ڀV���6H��+����"<b���p&����e ��v�U|�p�s���مg��Oِ�Kݡ;G~`?L��G��w���BJ��<�{l��t)h�Z��bn{7W��v�k����֝O֨��Wo��{|�kd��υT@�&?vHE��H�S���2	ݬ���0�;��:�w���>�{�����c�0�<��Y�����gE:��W�M)Z�C�~�Cn�IB�8��?:�~"�6�I�yfj`�T�x
f-��7u��hC��c`|�ª=�3�ݯ��7y�s�C�$*L��J�/4ݿm���	��	���v�����2��*�/1�L:F�DS˺u���'C�x��m���L������J�)���4���C�PM'k�wڠ�>~KR����׾��l
I�I+36)+d�X$�V��̏�"̺�6}'�j�#��m�j<6/'4H���oT�C-���ɭ�$fO @��4 .*42��%鮮���,������V��B�� Zsv�D�d<�����$M��"*q�#GK.�����Qmj.�Mw9�^&�$Q-�[��sR��VS��f�_��Mc<��ѡ�V�l����9��K�.��G�T�X%"����i��q%�9�m���
�����\��B��)����t@����X��Jf�¡�1ª�ީR h[�����yS�34�.v������٪���y:e�;�z߲�uBP�mGt��}t�� �5P�:��������i1N�S�@^P!`���\"�o��̇����^h�����䰕����i���o�3�+����7��BW��te%�׀�0\����"�fSi��O1�������	�`M��<,��P	�/=p-�HR��ѩ=���'�Hn��>���fj�ũF6@ʳ��+M���'��֯7�X!�X�򮶔�P�GZ��O���jR����W�^�%gN�n� �[���(��˷H�v����t�4�CǱ��'��$!�W2�ǰ!�܌���g�ⶪ�����{T[�Crc_m i��e.OER��0�����z-@��%Y�vԓ��[ƥ�.�&^ѭR��3��û��j�Ve�;@���n@� L�W��Wپ8!A�dYv?�2�нIM��<&���c�
���Q*�� o��wn�M���G��vI�؜�d.��d��\ְ�{�H�f��L��_���FVg"L�MTi�@�b��kd^5|ps��I��{pgҭ�^ɇ)'��b�0Y�S��G��I���g�.A�D7n�c����j�3�Liu!�F'�2 �I���}o�6�L�1<
�Og��'�"�E
ō�r}k��ȊF���D Фa�IF�|�t��S�M��ݿ��6r��d0���[AԹ+��p�r��vdj��^lF���Z�47��U繕�ޱ����u0�B-#ͣ�{��;�z���=ʯj ��Q��!O���H�l��
b�9��E���=�f+n� �]������R�N?>̄x��@ݴWAAP<����Og�]�_��2.'#�l��q�d����}f���> �x�i�Q�k] tVf�j)��ЈE��ؾ���2L��ʣOI�cӿT��r|I2cKl���h�Jc<�,���s�����zG�Ƥ�(wGBB?}��?�{w7�$�q�,��FiB�T����	�
oH�9���c��
.�mL2xUC%����Fv��;go	3��_qt��q�z (lk�g�H}��<���G��
���`�� 	}҈O
	�bf{1.k��'��(�
����\����^@=}�7ؓoH5��@���s�۽�	վCDY	�,���v��f]�#���/��,5�٫ɍ���CF]/�y9@���kƉ�- ��A�*뻩~��i4iN��-�@U< 6���ȏ���|{���hêz(���)��VPMb�vcC^	p���o�X}L�j?R�H�DLL;�xf�q�x��}��x��������uّ�V�#�4B�K�UF4ڊ���G���)�I��Y�A�h���PrAr�b�� ܂B6n��������l*]!jڴ��9+�z�U��-�� R���${&� f9�	�ҶJ�	���=?�wj��y��9�B�q]	��6�	=���d��e�q%���OT�HqM��<�&Ph���z�
�����# 7En|�	�o���ə��^%�7��K�` �^��P��L�³}���<�*��\Hb����@ݣ[�O��K�=m�(֙�c�o���W�7�դxG@���|����Q+���c��w�޳^�rV��n^c����X`��<���T�KK��� �Q"QZ׃�P�f?��Hܜ��eQ�O`1���(���`4�j�N!.ԼY[�ʹ�w�Oх�4�:�dj϶��!E�@�c�:"O�����
a�fǮ*\���98��]�v���`���z��`�b���?"V�ΑH��V�'|���ҕlq *�=K��oƎ0�4��`̫}|��dG�❀��Y64#h���|���k�}��g��il<���J�����趓ׂ�&a=���`/{tB\�.�����V�D�Ĥ�>�X�JaMZ�G^��̑hx.�R��)M�ȗ�[���Y�,2��U~D���z�9&�Q�i�H70�	B�І�M�I@y?h/�m�m��������t|A���Xs��0�U[�7��&(�ϵ�T�@,�h��%�b����*I[��d0��9X#�#ϐ'�f������R6njt�H���
����fj��=�mwzm�t��"
�ӏ!��N	�f
��4e�s
�O��ƒ׈e�.��� ���0x� :��<�6�3��e�<K#ɏeֱ6��8&�_�L�C�7I��LF����$�/��V�J�A���I�ѬR���-(��n�m�yns��y��bXf�@sk��on����� ���~&�\rc�L���U2��m�v�η/c����23^P:a��ی�^]3X�M�_h��e�$�7��L	��������uf,O�*`C�4Wq9��|�_`���K۪�����7�W�H����c:�$0Zs��Q�GD��o�9�L5��p:-`_Qz���*�O�5@&����=m��rr�0��=p@n�|7��Z��I�������p�ů�t�48�I%�Mvᡸl�H�I���D�$G��-��o��'��E������1?��،���J�D"G�����хDm��5b �`�GZ+VlY�T �C%�~kdp���l�w1�7VF�=�2:�#h4ߢb*~��t(,ՠ��;���sM�1���n�7�A����R��Sy0ѝ�)���ߚ1�JH:�7�<�R�ߺB�P�-�Z�y�⍶a�r��z\T��i(�SG ~�� i��N��J�%B��Ԯ��W����8��^�@�3��=��d�>%�ou���ljy��'��xa���4�@w��2�i�Mn�t�[v7�5���	ͤ+����0ujq�i����)����g>Z�n!|�ׅw�{�j��O�t���F�O�?��.�)06x��1"Ī�X�[Bg|�0 �ؤ�ЪE�h�GNl/�~�������5ˈP�r����žg��h�U�s�Ҡ3�U]D�I|�5�I*ަm�wDvY�.�yF��n�C�.�o���`0�S�<m�
�x��):�h�8[�t�ȕ�SLAj���!w��Se!��i���쟥0��=���3�l����;Vl����J׉Z�H�:�u�^Y�N��$���Ӕ�K%-zt������S>,�.QSH8o�F��	���
N�xF猊n���ǧM���ӻ܈лn��E_��(".{c@�11�:�{�i�u
�����2tR ?������n�<�_<q�x�ГH�rXca�Ѿ=�����Է��/Ȯ��pM�^�z?��ؑ��`,�=EP��t䚼'�aCߙ�7�R��?V�m_��5����*��25�H���¢�=��f��!K�+q��ی"N��_N�o܌�4$?@���y�t́��1V���O�G5�����@�4��=2XC��81��O׼��K�oNy�-rt�3���X�����0�������b��=钽��� '�tv�m�����s�K���B�b���f���Bs"c�[K�'���q�0)��;-}�V����un���X�GaU:�[vb9����M�Lqngw��l��D�gb�u�;�����ڻ̬[�Ψ]
�h�0u-mb�g�	<��Ε�SW"�DW(��w��%GZ~�5�F��X����;ܒ����ݔ
�(C5D�k�}gIF�(�h4���O̳���4`Pd!���"�ܾ��2�0��3��� �	�e6� m�ꊖ��9��~B�8P��+�$��wa���J`=&�'��[�J3���|/
T�6u����|��}s�B�����u*	-�b ����0m1�n�B�F��� �����J�/��!����?�Q�V�뉖D)��w���Ϩko����K.�
m��}�3��u���[�l��7Gu��u��[�Z��з8�p2a�$�R�k��t��7�&���ڮ��������r�t��c���R[վ-i�����E]!���SaFsM&���Ǩ9X�h���L�����Q;C������%O�ܑ�/p'��,CKi�Tx8��ĪHv��Ff�x��(|�>ueƐb�cM�Z���8���Ǹ�;o�iFr�+N�g1|�4S2�
��}�^^������TZg�2�;`� ����9ZPL�-+m���G���ui@�Qp�0�:�@l�ת�'\ˋ��8{�3+f���̌�sO���V:� N��8���	�uQ&�wbO,�K���s.�P<�j���f�����M�S˴-L1���J����b�+�7���Y}ٹ�Q<*�/Ӑ�Q��T{<*�=��iY?��������1��6��n�3����
�%��S4W��ȼD�����+�a���o���h�Co�9a� ,���<�����l"_A^a��u�~����}nGW&��f���r��� ��u��k��ykTM��F�Ye0��M��@
��7��&:� W��\�����d>X`s�U�����'*���r1Fr�٪�# �J��������
���8,(��:٪��.h#,k�����Ko�Cq�������1�(���ƥw�p�B|�����۵˺U�����=y2�p*m�]���'O�k.ە0kb��^YY�䆭��Y4�L�;�x�:���+���l��YXr�VH�[�V��%>x{�"��A������X4�y��M�Q��|qwI`��k��ud�3��r��0dƝ�h{���P}��_��.CC��vy��R�H:+ߪ-T��}H\�Rd�4���PT@�V��P]�,�c�G`�<-��Z2v4�j0S�%�1(�4][�]))|���{Ǫ��eͺ[#蔳���+?1�O�m���C�0#l(4�7�>��N�2��J��><�% ! @",�v��������~�-����N9�[;џ�z��O��1����t4�����Sd� fh�/�r��{�l�9�iR��|����6V�x���2%�<�����W�];��TlY��fb1e��y~O��|m1��O��͍�T�������F��_��i \�*|�U܎{IS�g��ӄE`��0��� e*��ҏ#���<��*�f�Gbp���L���aS�:��;>��0H�v�pC�P@��t����w'�	2�� ���{ZM PA�$����s�-����g�S}G;t�40���f���G�:f�8w~���N+q؞}�+�J��?��a��������w@�������O9G�GJ���d�t3�u���tγ�C�n����Et)�	�/�]�� ���}(
C��
r�i���IeP�(���Y1�+1��a@:�e�c�0��~O@L_D�?}��o����`���@C:�koZb��ASC�M$�C��uھ��������
�4�yC��U3�����l���
.�"�`E��
�(��H`AR�r<��"m��}`U;Hѳ�G�gp��R�F�4WK��7�; 3d2{��}�L���غjsq����R�k���tj��0�ɼ��7���Ν#o�um�ޮ`���`F������?���x�'�mӆ�h}�F�-��~Ù��S/��m��IŘ��'��d�؞�ut����02h��f4���tGO�M�L��S�w�9TN�(��Y6#��rd�0V��x�d���E�@z1W��� rW����84�����V%�(D<̆ ]��(��aS�}Ku*˘޳�.ޒm�P�5MՒ��}s%�ߐ'���A�j�VQj?����&&���k��A;eJ�p�bWV�̓���ܰ^7�$��x&q��F�l��ߓpR������$l���Hw��<+̋4_�#���f	��4flF�8�ar_	��<�Ʈ�.�2�B���@]�6�����k����m�p�:s�{�5q�!�_�*:�=����y)m��6C�^���R���6�&��>�,�0���F�o7$�p���f+�"C�����A�-�nf$q��&��ѡ��� Ȭ�ǜ�-x��bX:�"��x�0��s�>w�R��l?�,�SC	�j�J���1��<��և��\t�t:n���m���kί���r�V����dl�M�IU#�)(��|���v���ם~	E�R�����聻MqG�����k�1����ˏ#y��B���GTm1��Z�D�鯱��ް6����hMARD}?�p�i�".8�Ȼe��WG�	��2���\�\Ups�k���l]��ddH]�^H����T�@�޲�3�8�.��1�!�_��Z�I���50U���I�rsټ���BNQ�u��(ը�S'��	����{>L��u����3�C4���A*7��p��4z�K#1��`�����Q�K�n���n�W��+���Ǘ�u�V�.�����U���`W�:��'tb&F�?&�f�L�`)�_K��,A�x���}�4��KqG+l��p�{j��c�A;�y^`�6�ˢ2�0���c��ۯ'Qr��:���.RQ!�옍X�*�)TPd�PE�H5OŔAc"��0Kj�S�����_�.H�|F߱Nok�[�z=�S5�Tg;�2�L@�'m"�t�������}��碂�� =z���C*R��¡2�:h�,j�`mr�0�߫3"�B�1��U��X�i�	H�}����!�q[f����kD����)a�Rt��+K��Ozf��i0�<�p}h�;��/�sRE���V��	�Éώ_�d���	W��7;^Wz���T�L8�!k�eI�r���%G����Ա��3���پʾ�1�W���Ǩ���w=|�#�)ˁ3�9|@x�9�_W<mySB~<������H)>���H�\�{Ph�_ٯo�C}NsA��r`̣����@ϩw���ph9�`�H�5RQ���TI�ڱ�2'�$���q}�'�4w;��f"�S_�=�*�i����^e�ߔ=lU�ߢ4Gw�b;hZp�7ì��M�:����� p �ԏ��ێg7+g�������yÈ-��ɯCYN$*1�4i!�?͍D��`C-����HO�c�G��m��F�}��2$w���c1�v�x�H�p:�M'a�H��{S��(��,r��v?a�L���T����_r�9�Ay��R�Ņ�p_!U�}��-�c��1�a~^��峲Vd�[(��i3qDa�;(���ɞ`=�D��n	��@Ne�R.�(WuTTR�.rs5	w����7�3Rm '��d�,~�Ψ�-��%�p�L��s��mk��T	���hB���f~њ,Eo��y#w�����Rߔ�3i7�z��Rm���m���Z��e��é��?������1j���� ��G�ţ�7�F����Ɉ��˞;���g.^]D�=�ƥA�X�)��߰i�%kÛ2���re�a����HcJ4��L+ⴧ���^��ްeE]*�
���o���Du��-�r�)�q�o��j�ѮW$�9�^�ZL�qA����Ri����Q�{��UW����&I��oB'�y*�/_��!��)�6��a�Z��G��8vݐE��]�ح�fI Z�Bj�gkSq��|WO���{�}��gh�)X��&{o� %3n��k6����V�v>�E��zjs����T0�k.�Q�~[r��w7�}hU/�y��sL�]`K��o҂"�;]g��C�I���J��!�k�4�^"z}KF?�O ��13�|�4�#�xOB*:W����kg�\�%������0����k�R�$J���z�ǵ]<�QD#���(��m��gU_�r��������p3ެ��o�]��T��� B�{-�"_Ԯ�=Z���֧����������%�����>������e�&�U-����_�Ɂ%ekF�W�x$����p_�F�iu��@v�а�����ĺ/H�hTI
4�$���Cp4��U���w|+3�� Q36:bv�.[ހ۸��+�ާ {@�@��+�o�/G&WQo�#��]G��y4QR��ꕔ�O�P��Q��Ь�JY
�|6R�.Ah,�q4�$��t����`�6N�qɮ8�Yo��,Ym?��	� �c3����M^�����EF{������O/iVR)ÐR�/�u2���d�[��~p�XC�&U�(�����?�Űe��%?����p��m��C�� h@�#�m���1�=�-ǫ��<�� b�mˀ�؁>��j
�G$�V<��K
��Gg��V)�.L��S���~ �U(�A�(�@�~)�+�K����_��KйFط����_mm�0�	��b���X'��6(��;Q��V�K��U=j�+�~B	W�T
�\�E/|^p��v��
���p'���s�X~hXY)�8DA8�R.�������h� �b?��FjZ�ضV�lH�Р�\���<�w��[dK�PH�����w��u�U�JQG/d^u)�:"��"����8��ʆڋd��4����$��R�7�˰��~,|��T��<(�=��2(k}>���&	�(f�WH����E=%�3P)d�[�~+J�aՆ�̉.~>̂#�~���)8:3'Ό�*�笚�Y��O7
匢O5���YaQᢓz(�Z��0	�~��b��jɩ�V��wD�n�r35�YޔVW �cJƫ���g)�xO�00����W��Y��v���^&d����uEIW�2�ڸV���GH�έ��1^���_���v�X�t\YJ��/U�ם'�,��S<!̇����S#d���b��&�)��7(��Ph���sz�����[�#�����JE���!M��/vaRp������n�a���A���@I�T[Li!��	���IT�����Q䂺�	bmG�q�?��z�v�����D��.���%�v�0��lK�z�V��{�*1�*�l���MH���+�y��8*�ȺE�8ۘ�����L���%t�L�cU-Uޥda�~!��a��!�Fk�:��H����=��ډMs��@�#-� ��!�S��Ъ��pR��Wgi���P&x�mo-\��6��ѫ߄ nAp��p�e9�xij�)��e���pe��#�����M:�������������$p�I1��&Zc<�sE�-��ݺ#���9�`��ER��f?�䊉%��p|�*��{&�M/o�]��n�y��q��������~%o�I����ɬTB���v����XF��^��M���@�z�$�U`�4|ё�B�оS?��ZyŐ{�U���9��FNI��S�^y���`c��Y��o�^O�NKL)�W�%��p������in
�Fj����~��S	�u�4�$��D��E���Ɗ�*˫ۈ����h�ۨ���F�u/�O:���ʮ����O�Pr��K_��ʭ������^Ձ���Ɵ"�\��0�g��1�r�n
�q9n2j02����-Z��t�{7I�μ����y�,*/a�E֠���1*�TN}\�*&�Qa��L!=��/O�$����9k�Q<C���X٨����R@gQS�̯��&����p�B:���J�b�R#}�%�B|�Fr�%����ù����OU�� r����w��1�J��k4�"�Nv�ѝD�����)�Z}���p�2Ȅ�u2k�v�	�z~����K��u9�l�}�j��8>� "�9�#�_'4�K��:Y[t�F�+��\\�Ck�9���i�W�|`[�R#�F��^�8��9 ����jy��Rf���z�Cf�z*�E�d��T���7 ��e�	c��Q����Rs�Ϗ��n,�5�͓ �'��Df�!R�x�\����u��-<7���Ď�{�l�Fu�N͓���|(�3��M�@��~�U��,�EbB�ʞ����{
ZS�r����u�YO�d��ħz:��M�V8=>}��������P�uU�)��\�eDd������\���;WH:�'�O���9�F��(d�{X�A,L��U�͂���1��M&�n��<�(V-�,$���hԕ^=?$��� �_^�g�Z8_]C�6�$���ޠ��̟��d7�Ή-��C�q�C,&;���`�6��މR���H�@�U�8�ؐQ�}X�բ)Fc�'~%&���Q�#E+EP5������|f�����rKk�i=	�Z3��*�ͥ��-bU�ņ��D�w������g���S�}c/��q@Ѿ<A���倫&�)�Ge��X�w>L�b[©���G�Cfa@	?�l� }����o�_p�.�5� �\�T��H�+8�'6�L��s��i6*���V�9��|�7���b*�iP�i�n�p.S]�2{'8�yu;�%��I�F) T��0h��V�&T�,�(�~I構��-�a�჈���7"5[�X�Թ��7���Tr����^N�守��Bp��6���gg�uá�����d�v{��|��.�Ml�9XR�>��i�,�;ی&grQZm4#�sDa~z�#��w�OU-/&��Gg[ˡY�U2bS/�GJy�x+<�H�d��K��&Ml�O��h ��#���B�
�E���%�6Ѭz2S�Tiٴ�z����!���A�׭!fp��5�wI����p��Խ�h3R(�A�i��38�#�.s#��6����K��D3��6�R�˩�q���nl�j������[���18}*�gQC�f�J�0�]�Ę�a"���B�l�񾕉7�����-�	��N�:ۆְ{C
�c�Ǌ����eEԍB&O$��Ć�&�7_v��YKO� Or��d)[ �Sr��KeV���H7G�%�.U����{^�M���{�����cT~>��l�ze<�ń=�*ʟRVA~A�r�V���HxFaA�N��ͺC~\��CC��]y��G�v����*�{�Wb��Ά8H�<�Ff���m�`hZj�M�EO�8�Df>c	n	��9��	+*��mG'��7�O҈���M��7�Jp�í�mu�(r����H�H�Zs�Q�[*]�.�cd;�r����*��ƙ��(|BOu����N��
T��g�
�����k�di��x��=��r���騏�%�i������K���eR�OD8�]��-�LuO���<[RqpN��#�tjl�����M"���щQ�&}z��ٞY�L��I�ɞ����=����J�5y�B�>FO���E��|B�|����9�먿�%V���VS}�.��w�����@����o�C��Eq�ς`�T�[���/5Ȃ�� �?v<i������ܚLi3�����f�ᗆ7,Й���\��������Ìw�0<H�=�
������nŵY����br�evqh+9F��5�Y3�HGWB�t�P��LB{�5���� ��0��6e��[�IE�Lo܂N���@
X%��d�:H+���p�c�4I�����`;dc������'gySlˮ�U
A�/��(��
\��j�bj���4VpNt��tX��w��;�w���G��޲����^_~��Ј)�sBV��ſ���B���2�Q��P��6�3!�G,8Ѝ���� ~���R�с�cE�����Z�AA���8�{Q�-L����N�'FA�{jm�*���W�?Lű�S���@�\:����_�����y~�#�$�����������-�.�b^�P��:gh>	ɳ��q��!qY0���� B��=�����k��y�6G��W��Ъ ��7I��1iJ?��v��X'2b����5L���衛����ܤ��	A� ��� [���z����@��A=�~P]����}�#]7J������1���*�Y�GPɧ��f:cuM��)Z�ˁ;1�&��ə�0��7�k�f#�zf�x�L $�/�]�Y��p��2�DSyS�#�g[(El*<��5�6����%� }�ئ<�3�辖gl�:'��s|�������v���~����V�A��Z��t���\	5!���^i`/0�r�2��(Wz��ƙh��82V���wh̕Fo�����by2�n��p�I^Ck��Se~(� B��T�H���l�G��	��j�qx�N�ߠ�$��j�uϠ�/À�[+눌�{r�ϯ��WI)�w5�����;e�ʯ:�հ�* 1XH
E��Yp3�v�ŷ�x
����L�{�?}��5�����޽y���V�������Q�5ۈ͋ӛӘے�>����ҫ1k���{tC\u��{�N��"8���<�%�Q�~`wU�J��edU�|���M�e�w-y�Â�%����'���M��}[b��nf2�ù�4��+��i+ 5�N+�o�Ua��q�Tp������#��g�e���f�8��H�Q뜨ԟ�.٣eŞ�"/�%����`�U�rW���*�3�+X�C��h����L�w)��7j�lv�T&R?�_*����{}��¬����Dz��:QM�k��l�e{8rdd����'j���6�tG�uO_A8ryE�.��*��}�(�� X�����ʸ�Bbt��&?OM�(����x�h7]�ǁM5���>��+��шX[��߉1)��
rƳ�&w�]#��#p�'��'贩���5	����T�IDC����B2����{M��� ���'��_�i���ԁ�,e0�BS\Je���Zg�fs�_�p!,si�O2�����R(����O��|[�J�S
�I������و*P~�>F�E-iI����b�D�������/K�Fl�fXÃ�%G�l�~�U�uaǨN� A=u�q1O*+uE��9!|�np��b�4�ͤ��=�����X |���� u	��%��eb��Нõ!^x�-e�DXZa<���q���K�����-u�V�tA��-G\�.�y6��;Y�ȕ�Nk(��q��n�L��ϗ�9 /�	��O>�gK#,��T�QF��v���w��_v�CG"�AX�B��%�녂A82LI���n��^�j�a��YT]gr�G�䲋���W�eY]!3z�OOSĭ&.h��\��$����,�W���-YY$���QG,�ǔk�Nu�i��|U�2��i���By��¾v{R��8T�R"Od��J��{�J�?����46�좃�|/Rp큨N���1R6���귟i"y�j(,��-�H�@)�^����["�ۮ������T���}"��5L��\�w{c���b����˺*�f'��Ǘ���E*�^I	������t�N��c{�䮎�b�͐�2�,���<�;�Pj�E6�{G٩r����R4W)�^�����E�o86<ft�X����慇Y���a��}!>'#�o;Z˲��ʧ^L�Ouￏ�yR#di-�7��r���#EJ��OQы�����L�
�Y�$� �c�H��`ztd(�V��v4 d"Т��9��q��� G��[w_�b�W?C^�9���X��Q�3ݰ�Usm5rK�#h��ٸG���0ḱXUP*;:B�I��;�^��Zy�1/}�5�i��\��un+�|UI�ګ)��n���3~3[M>e��{��Im^�Z��Ǻ�fL���</�b�A�9������/z6�8\�@I�9��j�wx7�*��xa���xd��"R�)<��J#]�ڜ2}�\�a �=���^�c���aE���Г��Eț�	[#��*dwP?`N�9ȧ���d�f~Q�����㉓
\6\�:�M�)+�ù��$�]Hdn��,���յǞ��i� � |_����_R{(��}%b�N�E�6���dO؋���K�Hhڰ:�	�P�R�1�%[������Y߁D�m���B�gB�έҢN]�.[IR���Tm�[J����`m��0�T�7��M�T�	�ꚪ�H3v3�eB�9�W�]Ю�t[����R����*L�@��ue�5���j�Ny��]&k����S=t��п˥��q�E�m�Ĝ�n���"
_��ԥQu��J\4��}!���0*d�y��HTj��O81�;�`�M�,A����ƫ�O�{"����r��uȯ��Y���I����Ur 6FyTgK[-پH9sR�A��R��{#�w�M�����m�;)�l?]O�_��Obg�Z`+����y�8��Y�:���h}�u��O�Nx��<*�
��{J�~1��_j��7�-��x���p1f5�VCbPA�ۗ QJ�I(��dF,��2��?����<��Ȫ�6��h@� ����ꤎ����75r:�����>@t��.v����=��vM���}��Sȍ���_6�I�q7ɸ�u>��4�L��f�J���=�\����U>��sſ[Dr��/4i8,\f*�$C���@�V�]�ܵ0i�pjU��mY+�?�'?��}��N��5d�6;�"X�<�{,�`*��c:����ٲ��1�]�ltۢD��uu�.zx��vv���������A6��É=r�
DA��R�-���,�AޫxS������ľ;�EvC���ۨEG\�Xl���uBڕ��DX����jH�9�$ӱ��y/�r�<�3�s���̡��|#oR ,�R��Ibe����[��������7܌�R�q�m�Rl+,�* ���9<촰��M�J�攍�:�k�{Y��3U� �s3���:׉�|t�ɘ5k ^��A���"���K'�N{�
)�-/q�y"N��Q��*Jm�z�g�b$��f	��_P#��c��T뀳	d�����-ᗡ��2y8���!�Yx�Rvc� «[�=��(�~�o�����\��0yN��ͣ���v��(Y����We�������π���5�HM�Pՠ���� G��j$�g�o�/];Y*�F����l�:�SR$���`i���;ѧ�P�L�B�a��K#"ƚ��A:�~j�v*G�I<|�r=��g暃�4ƔHw��gE��c�ˣp�r���k�mֈ������[�Q��5���;��[K�K�1��@ؘ,�.�}(�YIH�`H���`�j�����)�����Y��2���zq:	H���@'"�u�E�eE�me��~A��+��b��_�)��:j2�)���M�N5���Z�#�A+�@B0��4�#R�tf�"��S:�H�
Z���VQ6��6���FFW��E ׷�d-���Pׯ|Y��;rOR�W��3��9��[�n5��~�;(��f��� r�r/��G��Z3!
*�{zvx�M�e����j�TK6�G����<�ga�������S}vݭS��_uW&8���_��I@�j �����afd�Ϡ��]g�jZ��߲�;]@�4���n�ގ{���W9���- �c74ue���&_U�SPt)�3^L˕��S���h�.�}6�3��Q&hm!��O�&p��V��˸�f������nW"���(�Լ�؎!	����L���eU�C�đ5cI����)|���ʊ��ERhr9N��@�{�n�jH��<�}� �t�:��/ &I��K���/κ$Ոs-s�_����7Ѯ�~)��8[��լ�[�Ew��J?���'�r	��6�#�P6T�oGi�|+���O@���fw�z9R�D�������� �u]l@S"K{�2z>8v�zh�`��=Mscb���&��� ��v;K|kD�S@���x[P��?ܑ�2�q��4l,Cv�=��4�;ܽ��rq#�_t[�$c����R�N��[���6z%�Җ�z��&�0��:������u�t���ފ>�a# �!���^��7�mxgD�`��Q6���k�@�Жj�/������*��V'��m,Φ��_9�X�e��e P�<�R�V\K��+�^oi����x�Y,7h�y2�U������^F\>���2� �ۖ�֪�@����W��zVH3Ev�6Y�s�R#�	��6="���g���˰�G��-��d#��Wi�7�_W2P���Eo�fF�K��<��M�S�-ʍu�V�\5��&��'&�?��y���ʽ�ϡ��=2f��ڨ��C�J�f�O���C�hh�0�,����F9��w�
%-�#��7������O���Hv���Ș�c��B��}�`-["�m\��ܢ��Y�["�.��}+��g�8��N��;��(�3����"s��1S��t3��:���%{��O7��yQM`o�鶲� ��V�5���1X�s����/~!p�{�O��UA��G��WX���M8��6)F��B��T�+��])���:�+�y
'�b�|�с��ܙ�c�{��ڋ��ږA�p24g��4��>�i*��
B��j�]w����Xn�*����TK��X�)�u�L�����ӿ��%둱�!�'J�q۫&�6�%��mpӚ���۩�G��L<ݲ�R��& �fd��ѥrBf�C�h�u��(�]��6��]�s�� ���_���M���ά��U 5��xV�y_C啼A':���%�]X6"��p�ee#^x֛��A��
j��%Y�D��QJ��\�u��K�l�(}�e��q\��̡ԾyI�.����,����yK|HT�����i1��椠J���#4��Կ��z��+o);�iCB�[�Aۻ�����|�(�:�ۣ�ݻňo����B;Y�F ���)�X� ·�;��VR���~ۺ!����(���vd�1��cSB%���T�A��Lڔ?���@�zՓ�ؤɇ�.1������-_ݖ'W�o<q��@���8�he�$����Z�Pk�����መ���*�R�lA�?0G�;�i�J�	�o9�e����2�����x��ǉ{�S��+J����kr���+���7,��,6�iV��V�n ��rcɻ}Hd��	���S�c�O#�&UӰc�b~mB8��Rco�aA��r �J���TԎ��79��f���`�i�u@\��Q�>���EW��5�f҄Ii���'bp���£!���G{Mk��-/���;][e�70�x��t�O^)���Br��]��Z�5S*��^(��'�>��s`�1�5�N�"�TG���4�a�%�tAݦT����ߥz��@�z+�i��j��6�2���S:X�&�L
��ͽ�W��U�N�ӵ������`[��,1��q=�����֜�%����/u�BY~� qZ��uD��F�%���2L�QlA��������p��B�К�v��!�H����������{�&	��{�3Z�Y��m�r*�c8�I1��&��6�Ο��g{[�Ҁ��M�@󯷛��> ��	�t�H����7��M���à'�MǋK��nC?z�~4qؤ �S�E
�Dc�G��P���&��.WT��+�^MY'��^�L9:��?�D�*Ls�k���ZK������Fl�^�N����F��.����ڝ%��������+V���̀�+�F�"���HX�bn@�'�U@�J����k����M�e.����	mToWpӤ����'�-cn�spB�수�_}��
O�,��k�'��Z��<�y~w|���e�)��������ɴ�]�#\-LZ;錈������RL�%�"�������)7L�#�"��w�N<[��ɍ�}�#���͝��1l|	�Bl����|�&���@[���@�7a��ə���!l?8ɍ�4)��#72����q��:F,��4�/��� ��r'N���g�:ax����I�m*��Mw�X�Q�c�U�d-�M�8� <kyNm�KF�3N6��z6��r�P]����]����
��t�pz5hȧ�]v)b$ �R�'�M�"Q�H���/����`F�~��7��Cw������}�O�7/H,�+E���[ғ�������8�7�ңz��d#�6��z(�HG�(
������V��\�i�pd4JH��A\�ƜK�jr��>�%��{�]�_������ $XC�!�s�ha_i�\P�4��V�4����9Y���!K�d�	6�#R���Їԣ�Z3�jY+���q`����z9#�"���s*���ї�p��$g���ɰ��f��ؙ�@"�OK@���в噘e�a�,�+n�`|~��I�<�֞�N�Gn���FR��ף	�1t�����d�̮s�`G[(�Dj5�C�G�D",Z�F����zޣdCά��-��j&N�]+`�LmB^4�ϹTՉa�!,9�`ܝ����C�A���N&Uo����t�u�I�+�2�1y�f�R�8�f֋E�m4��HQ�+�(`�y���eM��S�OF�j#��-�d��-[�����la�K���2{?�{����W��o���ʨ9f�wG��@�O"ox����F���Ϭ�}�Ѓ�3B>�~ז_1&���=��2��}�����.+] %�&[���?���j�S=���;������: ��j;`rP��G��ݶ�z+�Y�[o,����t=��q��I}�3G���=���i���U��Yo�	f3��B]X%�S
D���Y��B!��ɚY���T[%׍	��m�:��2[�@��)s����
�?8׆�g. ��X��c-A��?#��߿_F4�cz�hWkjʙ,��Q'נ�[�?W/6�/�����geaY�,F�!��J���%3���^�&�U����7��F�HNp�Y'�����r�G��ǳU�4(� ٔ�M�&UU�t5@쁦���\�ٻ�yP/<��"Ɖ"_�] ���Qu�����,B�Fg"�p!C�b\߱��a-�n�߆�!� I���koL��,��
��g~�5�rh��r�v���p>N�\< w���4*U2�]�QOA��-!�^��+Z���c�Y{<_]`�˦�2!�r�5}v�M:I��̢nJQ{�Ff��h��]��2b��	gO����~)��ҟd�v�����t��^��J��G�*�Ze��Zq�y���TO]�R�_��KD��L���e�}�!�T�z��XX�z�:»�ˬ"t����m��T��z�.��Q��
T��`cJM�·��:�gWޟ�x�Og$����n��>�S�A�u�Ν�t�"OJ�%�čiC���lS=�3���5��L��_���f�ģ.p��Q(�P�*ktB@�u�����w�WU_��@B����9zSG;��\���G��3���Ω�m�3̋aQ���G�1�w��Y��|�(K�U�e��:�����O�P�e`�HD(��p��G'�m2�/�$��hn���F��LLG�/�	��U<�2������b8�����E��1\s��~W���'���i��йB������d-If$���	r������Q�H�t"����h&���+�-Tڏ0�R�ûj�AfMo��uRM��
�*mmυ�>3U1ZX�v�|�@FL+N�w���7������u�{�Wb��G��_�H9�}3�wH�ʁ��7&�p���%���v�`NEZv9�iO�B
��0n�U[���	fc�A	��[�-�Cw�GUy7���s��h�l�*��k�q�Qк5!��(��,�DI`Br(rl��d��Q���7�A�ʝ}�F�5��? P��7�2j�=ͭ
$�w֋�B�9l;����>�`6�hp�ll��ǏtT(r*��
AdPJ��������v���%6�����l����� �ɽ-(�#Ә>� ��Xv��q-x7x=	��O�w��q���ʶ�)�K�[J��4Ay�m�B��k���3�<��ր�d(�#�6v\�
�OR��*&Q��;���=�XXt��5/w��צ^k%���k�p��MW�BB��:aM;fB@���uai�,�iX
�%+��Zo`��-�ԟ��L�v[�x�p�5$d�/gX����_�᯹g�.��N�Ɨ���\�S�Y4��u[3�2{S���J:��1�K� ��-A�%B!K)K��F�����A�Ai���C%��-�=�z��2�uM]�����A1'G��@5 5d/�)�Iǣ�1I^�s�c�]�Y�<Ï���u��SP�)Q������}nb�?Hχa�'aV���Q��<
�m���q��r)���Z���DhN�f#[�?�n�s�u��8��S�z|�|?��Vd�=$�o��fM�`�!Y�s�λ,
��q 6�u�H�����!w�"D�#���j���
�'/��{�iD"��0 �&W�T��R�䔥����m��rU����jJ�r��(�����-q��C*��l�^����Ow��
�{!�{��ub�S
&�g[g�����g���+hi�/rL7*5��9�&��Fu�䡾�C���y_�'���ܵ���k'.�nɦ��e��)di��Ū���M`ZA���:O4����]� ����aO�'�B�lA�;���X�����hf�?)e�e��r�-<���M��l�����[�O�'������Q�o�Jt��n^��rM�8Typ���b9�%�(��3����`��!��N���{�!�N����2.X)4~-��Z6��a�$g|�k�(=��!�s���m�8�e��N/9Bw�Ƶ����7�[�+V$���]2�:��4%ƺ`�z\���-����YY��9�K~+8il$��-���!tUWEz$X7i���:'Qa�]��1*�졡	���;p��2E����W�g�2/�^#����ǂh�w�ʍ u�����8���!Iؚ(92��`:k�
6�rhf���t�2��ьl�������ћ[��Ii�l2�U�&F��~H�����A�w'z�O��CZ�M)�ub�G�J(�!������ľ�ĝ7��/�d}��9���v�O��y�b�Â�ط����?�SG�i�G�q���Ã(�D��f�O��2#w��y�/ �+-n7"�`)T�İ�)se�{�BV���A>?6�W��"�u*�:���'8�� *+�NӠ"�%'y�XW�	?�'�fh�<4�oW��2\�׎�g��hXz��5jw�^�p�]g��]�r.�׮�"1w/�8\x�6Kb#�G	�&x���@8�Y�I��R�(��硣�!ci�[�G��c�G�
 �����q�;T���N�K�q�	�r���dZץ���M
b�1}����o �N��O.k�4��Rh��G�}ޥ����;>�g��>�N}�����Է��t���/�\�~�P����Q:;��x���?]V2>�ļd/�+��a�ge̱.[��'ŹJh�2�cI���P����h<ƫ�q@�b��d)��'�t!���;�оQF��+��@�9Y�'��)	�,<�c6ۧ�j|[n:JJU�uN�p�@ؐ�/��!��X*'��NLt7xg>��� �����Ӌ�U��mܿǵG.���NA2����+�.ě�����z�KB�a^��ACk��gc<�G�^���W��+�CV�<��?c�9V��9ov-V�}�gy�zy?3���k�t���8�|��݅�]f�η��}&�,mvm�O�;���E3N)9~���J�Դ�8�W�D�[U���[�� ������z���f�`i���z�>"���II�*�%�7Kn,9QaQ7��.��@<gg��T�iz��kX�	)�46��)f�^����>��
��+�q�uĖk���5͎�E��Z�=$�>}z]�J,K4�pw 12��2, gVh6�:�Y6��%�ϒ��1�<\�h�%yH�:�y���k���Gw����������΂��`��M�(���=����cj��Yi+|cǘlF$�9�w��	j׌��]�9c;����]:^n��Q���ia�^�ƴR�9J	d* �r3��`�-�����]{���~h+D;Ҽ}�'K�i�,�%��V1��{��9�t}�zF��e�����/�0q��k~,:4KJ�����N{ѐ���\b�)��:��/'�:�a_m�w}t.��k���g �N��̠�Ҵ�P��!_/&g7�ZyJ��
1?<+�2�@��$MU��MI�(� �+c�C%*d���t�֯}r�S�z\�m�+���N��~�� ���CTw�_O&�ƶ�����E'5��t�J@�W�B���J Ï��V�<����:~��+
�m�_O�;��~M�B��h��u&�d�i��4�l��ns�Oh|����q���T�M@�o���x�sID´<2�=��Dn��J�iN�D��JntK������,͊W��.�y��p��n+���o�K�^���?�[o�*5Ϧ�9�������%����U�"�$et|$W>wv���Jsg�]�q�r��`-S� ����*z�z�?N�����A2W�ȢY['�p�cK"�:��(�a���>{¤�x�p=�7���À��`����B��'���p.,nc�*]��LD��j~U����"�(��=@`s&����<M�*3��j����MVH7���V;9�h�"�Ȑ ow�|I��
�V��D�T,���)p �ZB�g'V��r	�X�D}B���;#c�<��Y^��Y����.�Ss��֣�]���yڞ��@���4%%+���z��d��W�u��@��l�6���Q��8y���k�TG�Ɉp#�"e�B�������F��w�Y+�$�7s~�1C���x"�'�f��W��5�D<�Ma�	Nw�x#H�-v� �I��6�ͭv��BN齦����K`ǭ!{K<5�@r���B�1Ͷ)n��-ųN� �8���	,��b�r`6�Q�<��pWY��4b���S��Mn����(��^5j'f9�5A�?$����=j�1w�7.�Eh�Q2\I#6'��5�D�����r����6��8�*��wR�yh���Y ��R��H�����ErS��
�ᜮH^ZH���$��a��O�w���L�v�����J%<�q�FA-'�Y��\S[{ͭ���؋��a-V��a�sA���C���[�6S$4v���PJA��;���^m�s��ר��;-�fR���bv�(��C�#'��y;�u�2�E�(
zB9�<%�[��t�h�MaH�]ڣ���9��K���u�j)�s#M1e�x�/$"�|Au4I�b��<�dDf�.i��7����&ڰ{/:s�2��z�4����|Ֆ$�P��˲�jI�q�� ��,��F	I���P�ɼHk;��霊7f�5�c(�qh���9,U�=�#�����EI�X~ˤ���Ճ�=���B9����Q�����V��%�T�
�Z}���]�eY�Ų�-����H�r������J�h�i�/�W�UQ��'��`]���tn�3N��C���X�\�-J�`��K�M�F�I�!T	ӣIkp�����f���#+���_K��Ƞ�����ȍ�α�����6�M_Ƅ��Uw��6��ቔ7��L*vˆ�����F�s�Ȃ��#��{����������v�뼠eB7��kZ��_wp �!�>���:� /soXW?���b�/r�}l �ᢾ�*2��n~��d��ID�(���΅t�T'�n���"���/��[/=m��R#�[�x\6g�|<$]S��_�'�jI9�i; ?S9�_�sn��^�
H+�9�Ɓ�n��;R	/X�#Mt��.�/�Ih}�S�
�>֫'�Çv#�zb�-���8��pD�
��J
��7e#����(�}C!��L�wZu���4bu#<�d�8�Kʋ���Y�R?{����N8���g��{lR����!/���Won@W~/멉&h�O��Oޜ��
A�����K���������UK5�s�գg�	ĀԾ���͵J�BKHZZV6�E<�7q)�t7� ]gS(`��}�����"7<T�(���4�k!8��$�(q�jA���ΧD���CLzb�:���F�s������{J9RBb�Z#\^Q:Y�r�k�4�QX�����E{�A�k%�al������)���_�ڄC���S�EY��=�} S� 5(Y�
u��ѫI�|zO��~Jthm~EC��~.';�4�����s�k�fm,g}��@�%���l���ʊs�Y�t�2��tar�������z����gi]���6��5؀<�s��}G�	�L��B���t�ƪ{�¡�~6�`Ʊ��©R���@Y�#B5�ĂD�c+�!N�Dk&��v�n]0�u��68AU�`ܭ�y\�;���Z�|����l ���iњ�3�Z�����[$r����b�:��S9��)�'jU�Su�|��*	`�@Da-�q������>�[ބ��	u���aK��ʍ�$�O�����7k�I/�F��.H�Z��R�&Eߡsfl)iA�-�IRO���'�������ɿ������e>ʆoTam\!m�J����Y��e	|�!��h���nq|�ܿ?��J�?�����k���"a�Q��yL��<кg'ufg.T�\�,Ώv��i�=�%��9#�C�;�)Ž~^-��i�H�i���/#��q��b-٭荺1 {!p���8I���me��Dt���P�����=��nW��/]XØ	@����3�"iPHW���gᮽG��Uzp�|K�8�p8՟@�#urv��j�.m�A�lĔ�މ#��7�)�w�.v����u"4�?v��ȅj��}�# ��{'�`�%��
@6;0�]ͻ�4����7�y���g0��_s���.����mXdP�	P�Ȗ�nw�*-�'�^W�)�PQ����s����"��+��爵tO3�5U��#��`������7$���i�}_�>�)�ҟV;}ѥ��$��z������-�b����q��0�� �1�N��P������ہ:I�E�cN/�� xT~�ъW=6����_%��IC?��u���܇�]R��te��7�w�H�_XCnx����(K	��Pw
*P}ۈ��{�[1�*):]��`
�f������x���.PH�`�Z	iwV���s�^K�K�(��d�S%������S���T�
m@���6���<�K�vjU�l4�L��j�Zm��t!���7��k<�-#��ĕ�\�����i+�����e��pƹ��7h6�o�� 9��Q�$�5�Q����M����U�q���!�v;���������.VH�����u�f�,�3Q(R�WI�Q�Jĝ�p��e���wsϭ�Rv{���`���t���dF��g�֌�.���%ʌ�G=�Y33a��m�f��*Yo��:�)���.�uP3���f*�ϒq���/l��\�s��%������j|�E�hv��j$L�_��o.�%�>��	��4.M�=%���U,�Vm��'B�9��%՟^*LK�6�6t��$��C���X��j+%�g�!�ɝ��� ���Ԧ�Z�C!�q���Q~���l5n�9��	�n���H�U�R��\�^_�_���(U��A#�W�;j��tf�܊j�����]$�"����%�mK��4��@�$�c0G��Mm+nA~�>ݔ%v��<N�̉����ZB	�Ƨ�h)��-l�e�Ȝ��*E�f3Dv��t� ����;!�[����3R����&Ai
�AY:)�� �޿���wNx�1�|��{�-�*�7얒_���z�|���9�s-��aMƲ�Ysg����d�so5<��N �3�R��n�
k�p���\4A�E���Ն�Yg�z�[����h����є���vRx�u�۰k*�y:G��\���������+�u�'��-��+IL���p�o�ۜ4Wg�6�b��`FLJ|�ư2]P��>�:��n� ��e�� B/�׭7`�nZ�b�va?)k�7��5� ŉ��z�����
�c���xi{B!6O!�E �M~n�vx/>�CG<��Ѡ1�c�J�U���+e�A�v�W[��T�����(�o���Y6w�f��]�q>CԻ=��1?���r��9��b�[S^,N�����+�c���-2��Y4�~B����zK�!y��)kC�i�`6�+��W�mQ��R�����J�
�R�S:��z(�i�����f���i�uV�� t��	>i:���6Quu��'���crںt~��\!�c���|�]���K���.⮞[�]���~}�{~پb�A�>��jlɻ���M��{�Ċ�Z&*aI=��dh���5D����9�E�c�@.и#Ŝ7�ܢ!F�PJk���Rk����uss���RX1Ѹ
���3{��kB�N`�J�����H�<!\q�G�:J��|��wl�����'��R��\��Yi��۫_63)�û.�׋g������-8+�4w�Q�
>�]�@���J��L�r�ᬕ�c~`=�|r*,萗"�k�7��E�5�S��������B��
�1���q8x!MXO�Ư/�f��[�z�/U��Q�^޾t�ҥg����t�FR�c$c�4��+,w�?)��?�q���ٞ�ϻ&H�K�"t_�Th�X�fF:IH�.r&��ZM���}4G6
��7&�����1!��J$]�{tnw8#���\����~�6J9E���C�Pܛ��L=����o��3܋ ���t���J�O1� ީ�̓��)�c-��o�����Q[�����6�����`���Ӿ��5�.]�W4{���4����(�W�r�q��0MJ�5��X��`�ֆ��B���(]ƌ��ev�2��,C=Ð@A�Ȯz֘T�4/r�?��M(-���0~Џ�f�{ޭ
�(�l:�����gx$�9�!k#>�2y<D���Qkt���e����L.� =B���;Qu��C7���)~���w�j�Q	��G�
OmuL��,�G�x�c�����ȳUw��?Z�_���2�-0	�H�Gb��.���?�Z��U���9���u Z�l�/�_����{
Ov�R���جm_�����2ح��?�ݾ���\i&����O�~*hΠ��U�@:��D�*z�hC�NM�-���e�����T�t�Jq���/ȗ;¤egʚ��:y�p���M��|?!>(,���z��l���BYˎ���2H;���M�@XF�rr8�v�)�zj��?)$n&,�w����$1Ή��g'�I�b8�g��0�1��p�}�
`;�t*0ry"z4X�[Tn�"��Kq�U^z��>֐�ߥ��Q�G1�h����Xu9R��2*[/�ݠ4����o��>����.K�R^�fd�oq��8�4�%��y�W"�N|��=�0S���c�,�!�H�E�K�<{��\oL\�V��M���;�W�u�b�+5��~��ReWT��Ȭ&�K�h�_a�D]w|$$Wa�>����!4`��@�ȇ��)Q��J}f5U+1�!�;�d���0�Ҹ����]<���f��h�V
%� 2���4Aۼ8�DHo^��E�݇8�K8p�U�-��ݭ��e��x�Ƚ�9v/�Lߒ���SW���t������0#�Ju\��!�y���NS��a�~v�?2k��y�����̆I��$����,�s�dؿɗ���yo�e?I��	9��2�ta>���\Z��W�>{��5j�_�?j��ʴ��<f�r�!��ErѲH��(��]�p[et�I�9�/����h"�F �:������G�T��ӏBu,�u0�L4�,������
�'"zu�'������<��8{|*�|����'�%$������v�:"�}�O���皎dht�zz�A�n%���h'2��q�_7'��S�.24�C��k�6�G���DE�d�YC��x92�ف&��a}*�,��:���O�kd]�M~ɇ��W�֛����@�?�x7�B�
��!����Q�ֵ7���k��>�[O[lD}�+<6P[��`�+���;������쀬�^A(a�ir�	�.���[{/!�fB�Xn|@������$�՛8�ka��=�cr}���1+9�H�~�P�
�gR,22��M�v�[��i�@�H����v`���\Ɇ��h����]|�7� ��/5�鳇s@�Q���S����=�����8c�>Mr2��<��e������,M帋.���-�+�z>�􅩎K|NL	P���v-eh}e#DH_�K�2�h�5��a]�JТ�����]I@?��U�eb^�w��g�N'��!������	YM-�����=�Ԑ��J���Ip�N!�b�M'C��D(+����pN����]G�aǜ,3�T��3_�!d�����e}e
*����Q��ZcOҎ^p��zU��H@�R;�d���89����O����S��������ڴ-���U�㩴�����`S^����_ �א������%�d'j#��@�cKm�;��5��H>>��\�ץ�x�
�v6v�NHl���%.�%B *j�/H�����oj��V������or�l?��q���Xs{�>f��P}�wB�{_���Ȳ�ߑQ_(l=������?����qŔ"���5s��ǔ�aHX�'3Ć��u�ʰO`3�x)�!p��Q�������-� ���u��F8��*@-7lhB^�4�Q�_:'Xk}�?�Nhd����Cn��n�>j��x�O
�t������J�,fr�VO����;��lNg�-��3N�:ѹ`]�A��,J_���Q]���䪈�
�Gءm��^L�/8�&��a`~�S~#��e�%X� w��?���/�:窯��+��� _�ƻ:~ϯA������I kj\5�V�[�����u�ZG�m�1I�ż�(:������B����.	�4v{d,B|�D~�M/����팫�A�*0�j�R�I�!�0��_)���~�����]I����0 �b�df� \Id�/|]�����9���[ة�`o	"j��\<����.ȑ4���/ĲS�j��L�D�Y�n���"'t���u�W�0�YO��T	V~m�Ge���U��0I8�2]rnэ�xҧUf<�#F`з���Ƈ��TK��*��L;�REj�A_骑ӫ9�b �ps��\=3`�7��e�bӿY��ߘS�O�"��h�W�y*�i�_<*xz!����^�^ou����EP�5���XR��� �������fK�Fq�Ѷcı3L���#�����A�,`V��j��_IÊ,*��Zϧ��E�����ǍRZ����u��\]���ޥ�6���D�����eA��)�s�N��C���N�ʀ�Q�G����{�G���u ��c���um��utͰ �蝕���I%"4�k9�t���t�Gx��4���H�!���N%�fث&<�- I{���J'0��/F�����J�3�d9!�(O���Z]
�{ȃ�l�9d������R��F'�Z��WE�ټ&��v�U]��٧�	a�Ԫ{9(H~
i���u��w�mѳ�!f�>%���c/�;�"�{��m��`�xp}���m��w��y��c��/���gV֤)�^��/ͬs��T�㠔T����^vn=�}��Hϩĕ���f�o	|��rCW>K"�����-���*T��±��k�ʮ�~���@���3�P>O �v�I, =�-P��yGAM�X�+�W�ʜo��׿�|����B�=ߟ��ULw�(�n��,�Xd,��RY|��B�"U�"�D��=��D",��0S�oNX���KM��_�'^��cǋ�r��8�%Y΄� H)�䶸C���`Ow)%�r�Wѵ���A>Q��j)���?�d�&�>f,�&�M����!]��s5#�!�T�;���}3�	48w$'t4e����`Nc��^N��1*<ǚ5���`Ȣ���J�J9��I�{d�|���� ��A�����$�,�3����T=�ݢC�P��:���Ô�j/����R�27���$�{i�:����z&vr�H�.IV��,'l���,{
m{�Cp��>��"x���=50�FI�9�D锣��%Y#��:Q���ܞk�������I��/3��r
�d=b��-�!t���S�d.�V#�J� ������n�7�H;�ڸ{Ț{������)��#����r����d
P�5Xu~�\��.&sW���}�2w�˲vy�I6��Bc��M�9�1�����vB�����
NS*O������qv�νʽ�b���z�]�����wf���h07�T���#,X^���xx�7�������΃ﴮ���C��t�0�6~/gC�%�9�$)�؝+� pg���r�.�����7�A���i�Ee�����Xÿyf�.I�HQ�I�1���@ d�L7?��Ah��������.�K��yu�f���P�ݗpؖ�R��Q������ Щp*�;�ȉ�fM9�Pgl� ���c��~�h�B�ҁ����k!����	Ś�!�Qg�	i�f3 b���J�Y&�8�Tp�\�d�`�5��O�	�����M�G�_��тx�kc+�ɏ�Ip��0���;.cr5��D���Y��,N��C���grF�l:q�&�֫����	���H���x�P��H��=CX��_K2�����`y�>6�N�7�{�YL�F�s�G���T���i�$�&+�>-��Р�g�lC����{��
B��<�ʿKtQ�+�5��u�ש��������?�;�`BםO�K=�z���S���(�6��fp�.>����e^	By�8U���pm'@���o0�p�4���O�_u_H�͡�I��EB�ڣl���,�N�����8K,�m"�	��/���{�x�� x^
�O�d476�/P@�;������&}�1,l�ɜ�JB��b��U7�^.�Yy>3.�#Ɲt�t:C����Ӡ��`3`�(0������U��|	R��z� ��bf�T1I��V�s��O�Y�ݯL�÷$���)��@�~����ʾ(�:Q�B������h���M����Х�f���<��VǮ�0ӵ��"�i��>�d�r�?<Ð\���q� ���CJ�W:��	bN���{N�� i�D"���=�0tS�ի�Dn���u6�Ө�)Yr^3���*��m����D�]d��-s�� ��9n���Q��Mߣv��Ԗ:��yB WE_:<{ T'I��a"<J'������!O �[;���Z�9�TB�%FV.��S�;�����lX¯���oU�<��	o�S��C���ikn�������M�� _c6	��|�22a��mg�[Mۃ���jI�D^%B:W����.���K���r�k�(t�c�+gL��-�Vu^�/��w&0���ze0}�>��`��|؀w�1� u����{+�j ��?�9��"��{ݘ�S�
-�w���������\�Py�@�hA�?���]�>�	��^IX�_����e����H�]���Fw��͗���"�${����w�v,G��\��S&*�4�l�h?P����9� a����n�?�}r-�}��8lvwQ$�٬�Sv�h���z�2����t�A�lr`jO䫕 �_ !i1P3+�<�N�+XL<b�A�Z�ʚ���
�.����~�4iQy�	hN�*S@��L�~�c�hࢹb��6�"'A$x57_�U�#��tn��eGc*(��������jR|v�v���*I�((9Ѷ59��4H�e���eW:˵�}��l��¬�~��Z������ZV{D�f��A��N�&�n�ը2~���gӋ3 ˽HF�Љ�2C�lVo��R�ܽt��[�Z�#�,�Z�C��b`�9�θ{r] ��In�˚�F"�s��<�Ʋ��t.�A|���&�M�q��;�*CB��G���?-ې�3[C���?�(ϒ��t�i���<(��aw��Hx�V���}@�1��N�d�V/5:�|
� 55X'�/M7�k�Z8aPSR3�r�/P��m���VRMt�G�:�����}$~)g�nϫek��A`��3��H)����C�	�&��N?���8��4�}�;h�K��NIHF��~��`��~#�"n�;�4@�E|�4�A��%ѣ�X�A&�x�ޯ�!�`)l��S{{���j����d5Щ��4M��I���{
�Q�/h����i�citߚ'�+-B	�J�s��2><��0���`�f�sC(�����;��Tf�N��0� aIn"{�Ad��)S�0b��5LlGLn���L��Pb�Y$�ݻ��A�H��w����@�0k�,�p}�j<���f�y����� �������:�p#k�� N�K&��7)o��g����S�K��߁
jm<��ˑ�-��/��@~�p�2֪��:�U]{��>��_J�o�WŜ�T�F�F ʽ�WhBDb��o)���������W9�Ox;C��%4ɔ��&|\��7)h&H��)�Lۑ+���(	����X̪��l�0g솹rH��Q*�8!����M�6��LԾ(X��0T����ܒ�B6�8��$����LN%��Ŏ}p�;�^D)n���k�~������Sq
�g������C��{��N-,�d��1��=BE���	��WL���G_1#�C?)��cg(�'�36����JL
��3f姶��+ⴓi���z���
�����T9Q��W.�-d���K8��n�͖���?�杼�r�Es�)�xƙ~qX�4
��hF_gJE�v��;�pL����y]��X�c>����Y+�(�?��PD\c�?��'鸺!�'?E�ڬ�jڊ�?F�Q�}L���q�e���Ӝ9��Og�2ҍ��*P~��8���]K����/�FΧ�v�>�r��%��̣~�⟩�(�M���뤾�ଽ<�*�|�0@'R����3*�X%}��(#Z��3�Zs�����
��o��� ;c�`����Aӈ��,����/�*c�5�K!�	���yk1  ��x�\Hd:Ş큏�ƶ�͜M9�י������҄TV-Aֳ-?hA<��ljPi�2��h��Ǡ٤C�+���A�z����J��I�N����B2��W_Ds$Ѫ���~}jՁ��#󙢒¶���Xڳ��e��R�TaT.�w����Z4���@=<��R�x�b������A�\�?�Y<<c!�"����5l��P�ˋ�B�9 �����Pj�ה�U�P��6h���m�w[�����@7�dO�X�i��c�'��x����4�ݔ�Y,�����Aӳ3�2�q.h|�/9zȦ�ڊ����*<�,|�o�K�>��)9"�ui�B���S�O�ࣳD�5���Q���1��e �Z�~�O#��Hx���/A�O�B�����g�jc)�L��Nc�)�����mpk���8�_�p�F4U�:�Nb�8�7/�~��P�w˶�����yUtx̖nq�xͮ=.}bo%�X����A�r�F��O�㢻�E7�v�f��]��7�,�઴��H�#U�i7ĻGY�u��muj	������*�D6�~o�iHZ^N%�XEі�������'�0_����fX�W�
��u���,����<G�ų���47�c)�'�E	0��So���ʤ�4=���<�9�'�**C�����	+��6e���Ĕ��X!����:���B^�T�$i�`��t�ܓ	���K�wB���};i�U�0�5mn?[X�"�ӱޮF��0g�j/�|;�09m�VܽЅ��|K;mX,�����0��_�D�W�W��D�͡�����^ӎ^�`����D�}'�f�ϱ��燦�:�27!�mB0�Kx W�p��[Yrh�z�X���j&�ct�9\�!�bnr}4�|�PP�ۿ؅]C*�j/Oh�h�!���>����5�X��-����T��DT�p]��f�=i�_�H1
d:��f��s�S3��8c������ x a�Yp�3��~��0�7�ڣ�7���_�J������7,'�-ل(�,��M�S��@
��#��$����2��E�Ï����(0t�ԩM�4��9!)���?s�26ّ�  ��0~\Iх�N[�!%M�_D��_��v�{Whi���*��J�3Ŧ�f���H�e�`�8�^c�:<�L��5��������m�P����
�>�1�"�0�G��ˣ.�N�L�! W�<���$�)�
93 �)�?�����h���y�G8�\�O���|�)��Zr݂�B�4���h�oc��1�;ef� �܆d��vRh���)��|�u$Z�:
��	י�r-L�m�55؍D�9M
���'3\��r
oڗ�c�I L��C
������"
��x�q扌���Me�y?'~���G��P�m�<fOW�=�Q/m'�[?Ȅ�0}y����f�'���5���P������s�A]% K�aJ��v��O}��6��Oqjg�kmIO��E�T,�߰@=&y��O� +U�ڡ`�����џ��b���gW�ʜ���tH��h-I@�zz�ǈ�Qľk��bc���d�+�<���"�R��ȹ,_�]e�Q/���h�P}x�"�c��_5�-Zt�eF�_őK�M��}8���%П��3e����?��E�	9x�h��B=���nX_�
���4�n �FS�R�|�P�4������(Gj􄅦>B����^����ŗ�!8u�����$�:�rN+��Au�8�o}�n<Uzt�F/-���]�{$V��'1��_^���F��~G��T%s�5M*ǅ4�M5i[�ۂʰ*k��\���F�R�,��[��%���s�W"DBC����*3�8�Ro�LfD~���)�Iu-���.>6v���g�ș�I zK�a@�hЍ��=B������������a����j�tcӧ�ݰgZ$���2�z@o	g���(O+9<6������)��8f���6:+�UpCVX!�����#k-��X2 nJ��8�Fw��Z� ���i���;	%y��6J
I����җO�Fb���#�)?
 �5��o��]:�ͤV�?#;bg����F-�柑p�+�м�u�;������&�`-�8�`����W��ݍ��D�0)�K1�Ս��������3YO5�UÉ1k�1���	�@�2�����KDu1�Co�w��<O>? �)�h'���V�����PyB�7�8%��i�:�I�P���G)��Ѭ�t���z�-��Ò�D;�-�2c�R�`+�h�J �8d�����(��h���;����63"�U��ʠ�Wq�r�lq�+��(S ���a)M(�9i��a"j�1|W=z�����0,n��%h�x�0��R�������1j^\�!}�`;qr���o,ݰ�%d���7Z�83(8���
V!o%��;㰝��Z�r٢����hS}��0lt�d�\vY9m��Yg~"�?H��_��aX^�|��Y�#�J C�jr�bCl��/�m.��6~ =�*���K���|����.~���Yu��Ym,K���������[��a���5F�gʹ`�/T��~�޿X����~�=K�d�ɘe�_��DFpZ��D�A}a���9��D�u]�X1FF��i �v'�}9`}�
��d��@�����s Or|g���(�à�]>��j�Zr�j�ĿB�}�G�*rj���6$ȼy�pT��&,Sf2c� �֯�T?����KzOt�Y�AS@!.m഻��U���Z�؏`�.�R*V���*Ë@4h)>�P_Uv0�긛�no���O�C�Jl�<�jF�PZ�/ƹ.[�\c��ƻ��OlZ�Um}D+�7q���a��	6��Zrݎx�v���e�
5��QSP.�Db~�w����8��V�����|�}�e�h�Ac_)�x*Pql1/c]�W�.?���s�.��o����c6́��8��^f�&6K�?��5�i��Br�ptL�_��U�FXV�C�h
b'G1}�/��x�֓)�����e]r�9}C���)i!Q���t� ɏ��&Nk�I/�7�29m��\��_�>�?c��Ms�$�[����JE�>-�4k�1t��o�j�i���b7��6k��x�"�\F�����'z>�FCĈ�BjGЙ��OV`�t��w��~��6�ձ�ӺIck_�slY	xgN��n�N����#D��Ӑ���f�)&�:��+��#�\��j��_��fɠ4�|ayp���ld4�7��j:.gY��4�� �ǁ��"�x�^�c31�f
'�����?�g�D�h8����hgӝ����w`fu�:�w"����63O�v,�7��@<h�"F�mG"��QS-Փ��� ]X�q��ˌ�'x����<%hv�NBO�t-�I�U��$��-/�9A,�~.I{�$!@��@��$�
��y�O�{o`������ ɯ0 ��.�30�������ln�K��ԅBJW�d%|�)��f?)����A]���i'����`�5�o*���'�R����6�c��X3c�w�`m�f�-j���e-�����K�H� ��D}	��]%���յ��޵��� ��?��O�R�� �5��lp��uhY��A,+�o�E����Tl�Շ��MhO�?���/���� +y�u���ǧ���R��
����S��r$�{��:������ʟaI�H����D��k�����6���W���,�L��ۑ����mR���g;F9�,$��r�6����i��Z��k�f��ۑ�pIB�6��D+8)��-"h�F���r�~��A�@!"��s�&�(,�B/�}��f���%�����.���"e
��F`�Ά��CK�k�ߪ��/Y4�M�b�eo ��KRL�,d�����5�F%(B<.zB�Ԡ_� i�b'n:�<z���`�	�N�.-�1�]� a���v��->�zt�?U�x�,d0|9�����)�@*�=�c�&�1]13�'0L4���控I�6���<�"�מ"&N+�
�< zY��2{�mF仸�/�p���W�+����Pȳ�@F<mO���t���,����|=�cH	{T֐�S�ߓ��T>h3��:��ڍJ�JXt1~�}�*��Z1��bTxl����@_�BC���nm%k|ܤ���p6)"j��� ���_V����d�G���X*"�<W���cK�����r7j���xu�P	{'qP pk��n�x|���0s:��o^��lCe�E,(�b=ʾ7�A�65�p��8��ˆ��/Ql���[/�L R|���6Z̙��Pl�]� �*%l�� u���&#D�R}�󤎫D񯅟��q�����op�C�t	��o�U�zM�X\��O4��0�[���0����26Y�ف
Û��_����4��/G �S���e��t�j<*>a⿉�/u, �,:'�{���ԙ�-swg.�+�g��T��������2_���I�>]�:b�%C��4���!ldZ}8��Fl��fP�.{;c����N��ˣ�q4��J�,�Q,<�e	{~?����C�i�����#�PI>�_RVBL�|�(�[�wX�#F�/�,{�F��[?Ck�U�J����y�����A.�|�%@�=�,�	���k��%)�;ɕ�(|"FBC��9�����䕺G���@��WF��
����c�l��4�wU�H�`�>?��*��Tm�I�Ss�bH��"b�tѾf���Ó��?�e�zv�1Lz����Aj�5�����3%�@���*����T�<��gV S��cu����*�)��f�n;���:���Z��o	?�6(�<���X8��u35���.ȌN�E�ٞ���P�7e�ѫCVR]�4�W��=��_�H�=zaշ�Z��ˎ^Pm����?m��ۈ;�ʝT�J�a�FH=]��e��V*=ZqQz�T0�=7b��I,�s��n@GF�t�g�)�i��I��Ono}�gN�'C�~��B�[D�۽_n��h&BxX�D�È ��5�'l[
�CgY��)"�)hg
�o;{|jj�/1t�ЕdA��2&��*-k��.9�P0n+�����(|%JT��Ev+j6f�t���iP�� ��P��$���><p��S�@R�)�n锌��0��̒�`���t؈ڿɧ{F�NrE���x c�ۙ%�[����4�C*Cr���T�[���8>[@)���G�c��Ph�k7�FD� �n}�s!N���}S��1���!Df6�c��������3��Q��S��0��fB�߿�~_�)���>�'��@,�	2�U�x�SxG[�|��Ɂ4ʊ�~!��6�e��� �8�Қ5 I�3[E=�����k�@t
�}���*�c�+<6���F���h�(p����F4� �`��ڹ�R
{L@ `� ��먈{-ԃ=Sp )=��X!ՄC���c�c �v7*M��"��n����l����Ȕ;���j�*9B�Yޠ��|�]A�҅'�44ǭOѯ֢RH�+f -�8@�u�[Y��o�7�Xk����6R�n�(o�M4FZ�/�[|��0l��b�)/�������eGO�G�LX�~g�n�uc��*B�[�Ew�dw�~��'-K����J���t�$�k=�Mv�OY@C��� z�4�3� �L�H�����7Lo���D�`��0�j�o"�5K(������FN�	`s$'9jL�).HNXMˤ�/	x���E6������8Y��Rp5-��BH���G��iG�!hu.MD�jG���|y@����$d�E��܍t���Wd`xc�Om��`��O.�jaŀv���N��ԟ�!Ĥ|E`���f?(#�E�9�BV����L�m��e�[����k\\����p��_vĆ�)6����B�Xa	������*1x��f���Uzf�N��Y���#pG��h�YO������;������J��E�{#�]��_	��z^����5�L��i`Ct�#g꠲>���tYv�M�]�����}Uԥ*4ږ谁]f�'���$��$�r'�j�@I��<.���"��l
�#�2���"wʙ��+�����
�a�KA����I#��b�	��o����дʕvH(�v��d��頻8�Z�f��OU}nՒU)�;�a&�)�+ݱ%���#�v���R,gfD�04\Ǐݛ�מ�@9�XN81'4.j5>n�k���7��:}a�9	�1��&d�m8�T����x1[Q�g��yG*��5�&(a����� Ʒ�-Pa�n���$��.���-��J�G����S� ��>��s��Z��m.��`��]�j��o;e�����k���7�yV����v�p�\2EmW�]�C�$6e�Ƿ7w8���58q� ���>���x5��à*��wj�K-�Q��X߈����)X��k�ʶk���ʰ���1
�`��ȹvn.���`���5J���g̨�ň~��Ԝ%�o3`�f �֒c�t���'Ć	�A�WU�v�\/�����q�x\jܟ�!�')�L� �b�5�-Lh^ʒC�U�}�C���.�B8h$��-���[���=:~	곆-c�`zŷp������E2J�^���eέ�k��F��f3�^��0"wH�Y��ĒC��j�?eC�3rt��寂�ٝ�o�,Q����#�) ����8G8.���R�R�����*�=�߯�;��!�)��46�q�"��|jsJ6q�$��Y�ϯ�|}�L�P�:�%o���]�bMk�ӕ7�H���9wh3qE�o����Ҕ8��&�8������g�%$7x�k*i�0�pT��E�To��@�h0��#�f���3������ IZ�g�C��F�%�{��5�4z�kO�����d3��� �)	� ��G�q�V�$�)	�1$���Eږ�2MDZ� )���������>yI1c/�-�e�;Ѣ��T�}u���h<���ڝ��?K~K����b���'��g��X����A���Sw�(��zl�v8�¬s��)�H.�C�-|���$�c����c�'E�M�g�&����mĠg}m�:qAm�\�h��
-��6 B���:x����Q0���j��5	�Ü�y@�a�\�v��oƙ�H����fΥ�N�������ˢ\1�G>��9epס�gCK�o��k��:���è�X�3���	ɚ� S��P�ۇ꛽E8�(�!V�6�əw��gլ�v�I����x���G�AkI���r��,�-�lޑ������?곙���b3�a�����W1n!�=��~����̇���\�ϥa���`	�ȣc���mdH`�H+�PhU���dٝ�(��í��/�h�0��V{���:�ׂ��:����?{�^G�7R�oҫ&K�}<	'�ot���=���c������K�����S�1������Y�Ah?�&_{��8zlP��uukI��s�̶�D���h�խ>�θ�oQ��1wޔ-�ŗӷF���l��|t�]��L��d�q)��6�Ck�W�Ǝ ��"�I�w����ò$���ٻ�⇝a��" �x�'��K��+Jϟ/�ۥ���k���]:��&���}��\�ygW~T�p�LIg�̋�K~��Ք&Q�-)�G��P�îpǧoX/�����=HRϛې�I���:R�鮻�#��]�u`�^8�{�v��v��� G�z�3�����l= �R�U"��7EFѷ������Iy)ru��u��M�|!u��j��5u鏳ZȽ�Y�t�^��):I���
��濒�+v��J����q������&n5����`a��)�e������?�;^�t;B��@y��X-[�� ��D�~�mi�Hd/������{Ȑ^:b(�0$AC��!!�b���&�m���Fx4�[I��sG.Kr��.�$ �&2%��.�i�*(����ѣCa��N��b��[3��s���TpQf�֣*��z��{rz8��Vo^���]r�y~�6�8�.[l%��y������'H�=�N�H�z���r)@�)-/�uC����rO�a
 �ga�m��,h�QB��{��h��8m����Jj�ٮ�&�W͚������Jk��ȰI*�**䣵�qT�{�n�l7�qb�3������7�����lR�v�����)�t�~�E���N�,[_Ж�ف�=�_��.�0���u���#;�Z l�!�j�+>c�j���Չ�������2�F~�ԥ�@[�JS���B��r+��:�~!z�P	$Gx��NӉ�O�N{��Ȕ/-�M�J�`�b��I(���Q�����<F���a��mE�����RKw��׉J��SR�xĸ��� Wd��DI.�M�%��]*(�AY��^�T����2�,���)q����$�)�@�>�/��-�Xk/[�V��/b�6�%��hϔ{�fiH���3D��>���;zP�����3�e��S��(�x$m�Љ�|
<���\����7�8�6�"T�Ѫ��]�e�.D��W���:�b4a/Ō��rr*�Q
�e�$t���O�6`)ŷa/�ݯ��r�Or;��{3b�Uf���IQ����XU<.3X'�Є��_?i��V�ˠg.7�R�І�>+�܄���_*YȮDb���5���ưJ��u���8<�G�}�wF�h��]P�h �[�S���퇢�M+El~�#�X\�1�Wr2�x��؂�	�|H���r�C�'�:�
�j�Bh�# ͢._��vh�:�[��vH=�o+B�V�Qg}>I���=��H�ۂcCKemY��kPM��bw�K�xY�iѼ&Xk�m�Pr6L+!�,��˽I�S�������f����J�FmRx����,t�C^��]9��J 	�o��ڻ��pcԦFX�̙j����9��. �ue[_�ۄP~A�'ϧꇦ$����|�G�$[�e|�y4�>��dN/wE#��;O"-#PHǚtHq���b�4$�N�S�̜
	A�b�!��-	<��XVr��l��1�ii!߉��2���zr��������+�&���L;4����+a.�[ȵX����TU5�(���?�l8�NJ���ڙ�ùC�.Q}�8%�hL�w���p	dE4�j�����4s!ҠK�48JqK�g�}}��%�s3&�f������چ0-mZȕ� ����(+Ht���x�v�����+�`@ʡΏ�ф���;L6�Cl|\e_��_S!��Y`ț���	a��%��e_�O�['�ϓ%�d�t�=>p�:����^;����\}����M�Br)��G��i���C��|�Z��~�MĻh������a�}К@g8Fux�t�-1*��`��5*(,\�3�<D��Y��,�;7\f]Mj��)���2z����3�2s����k�Ж��A��;��lA��?�@Ԅ�,0c��`�\����8a�M��7�z�M����$��~ ��>��S�֍/�6N�:�/��3��Ö{R�}�)�@��]x��k1c�a�8���E�ǞĲu�}(�Q�ؓ�9
��'�MJ��N��+�(Y��m��̗5t��~φ#�)�WP	���
��a�@|�e�{�G��Yte_lx�S6	EPP{�H�����r�NŎ5Pl�X�2B�Q�&��>�F8���Ɍt�O�|9f&�����˞@$��	�Ohʌ�[�h�5L��ٕ�H����J�V �	O���M=�W�`bM7��H��L>�?4w}PMhj�n p~�+��t�j�w3tZi��	���JNc$9�����y;zqۢ�w��0�O�5��
|ށ�[�:�e}��]�k�����v��.�pT�U���Ŏ�jws�=>t�Lo:0����%BT�~���M®��j�FL�m�!U�-V�Ik�b�n^� 1�1��,<���O��q��e�]^F�MoME��Se�i��C`ޓb~5�u�8n`���Ѐ�q��gKz������ 2��F�����������q�fPP�0=ts!�����W����@��؄rpa�yodW����k_�!�t�����[���W[�!���p��1�/C�^�{UQ+��茴D(�z���.��f��d�Ij?�N��M~w�ѝ-��|�X֖:��jԈ}�O�A�i���B��o�l0g<�hv���f�,�fG��9��~ԫ/���wR�h5�ж�֕����B��2a�-�ո�)k�(�2�D:�Y��!I)�M~�% �F��`�C�NQ&U�M36�������^�Cn޹�9+,��Z�)��������v�Vf�ŷ����-�H�,a��P~~u����LR� �LKkˣ1���4�]���hOר���Jd�>�gX�:a;'�Ϛ]�#>x&��G������9��F��9�]\\�<ջ��Ƥ3hL�B٘�⦑B�� �茺 5{s��?���/���Zʶ����^�4�������� b�?����2��Tdo�y�������OKGF;���h_)�������,�$�(!��[{%������f��G��n�Q������� X���u�����l��b�s��8P�g~��\B	������F�\�D3�yF�-+� �`t�)�<Y��'��qs���ԓ��@M�/o�.�邷�,.�y�9�0�������l��cMf�=g��w����Y�DAN3�	�[�*:Lhq�˹�C�#!гd\��(��.�C^5p 4����%q�9}���Q�7���g�+<I9�oA�:�Q4������(���-�6���Y9q�ͭ<�1~���gx1~��bV�Ϗ O��Tj��̃��\�RP�D���@(��Q�Td�%�U��8,2z������=U��q�$̎LX�'`���3���O��\�RK�T�Q&���#�0\	C�)�[���]��{����~M��1�?5�"��iĳ�n�*�Xjs����G��#�Va�!��/V3Z�y[}4���%�Ŭ�>��W%�K����D`(TV�C�1g�RR0Z�=F/��G8:�)���c��� ��6Y,��;�����R�v�wm��MM��|ز5S�!�	�wF��.
��?��pa�KĖWm�� ͼ��Jn� ��|���șbD�%lmd�P�F��H%VZ������,ǳ˹�g�8N��
g��D`��}�d���F���3��>h��̊#����*Rn�D�z���N_����p���w)��q >���L�����������M/�*��X�C4%�.o�]ֲՋsL��^��w����_�uW���j��'��(7G�|~K�E�7�ٴ_��hGNVq���A�PɣJ�z�&K<��	���RR�ӈ�����E�$�ǼD�r�s���7y�\m��Ŕ�}��;�OVr����r95�/dY:�&M��V����)�3UDe���5!���r���\��xD3!w9��=f��>|���f�Mŕ�/b��q29E�i~= q��if[�պ�������㽫G	?��lɭB�gbvx����p�iNJ�ݰ�O"U��8��g�^4k�JP6_���hw_��t��B1P��RJ�E�:].*�Ug�8�m�Z��n�j��O��rCj�����_�*�k�L�ٷ�
� .�Fp5:_��+D?��O�[+W�����[�qo�,`R��"{��-��V"����:��.Z�,�����Y�;A�Г�G�I*`w�V��M ��t�u�s��d�m_��mL�w�N��`�����%��NP�)�QPlO��>��D�#&�rE�]��;�]�g�B��M#�Jz�;׋|�Z����n�N���0���g��[h�O�����T��=f�Um������{9#:ζ��'-Twz�=�������P��놜`���u�>�Ң�l�d,ݚ\��`�!�t9���hA�
)`�߰?�r� �B.yh�h��S�����U�4Mh0�����/ೂ�ޔ� ���+���b/�Ӿ)�K���<t��{Z�����?� ��0�����|5��vH�*��A�B���	_n�h f���C��j�y�D\V]O���fy����AY��!�>��@
����!J �:N\�H��>uZ4�k'H�+������j���xyԑ�u"�R�멆�:�&���� �[���������I���:��:�E�n�L[��^9��+2��Z*�=���r x� #�~��d�B���[�Vo
�̞{�d�0)����{��F�%�y��RT�y2�}�#&`�qU��M؅�����'Dx�O�b	؉~A:^����u=��v��SǪ[-E�B�b�!	���`�Ά׽s#���Df�.6Q"\W��H��܏U���u�Md�W����j���
�.��I���|��dG��Y����U�z##����[��s�i�pjt�0�$�NX����P}uk$;�_,l���q�G�2��گ�\=%[�͓�-��}�����C�<�����'�8��=��Wy��t`#H�ۚ<�"8�G�Ͱޑ�Gxa$�^��{|Q�P�W�~�-�d�oz��1��X˸f�[�mڥU�Xow���Y�ۛ����|5�f7T�Qݡ�6���b�b���'�V������B�N���ڋڷ�1YO"��7�k��p�h�����I�5��賟�!�|rm>��n�9@# �@����8� ��nw�c9>A�{'H�5�R�q��h
�\��;Y�% ����4z�Ĥ�IdC�L#	��=�I��q���rד���YɅ�l�iz����e�Xq��e�P]�d�E:H����ha4`8�arV�<��  �޹������#Nu�뭟GlnCp��æ3|��)��j��y�n>i=z�b��a-Ky���q�HuG���(��lZ����E�j��hW���T�Pii-X�(��w/b�MD�w��Y��d�շ'����G�ص
�zM�������g��i1���"��՛OK:O���*7��!��a~P�"C�׉�hLH���@~�wjW@f�A�f�e�"̶i �굪"p�,;y��o��}ª*м��	x���2�?SZ���W@�7�@��ͷ]������.��e��kU9�e4�9xZ8����%���p2o��;�bbt���@��O$LT�"b�iTq}Y�y&��ցR��nݝz>*�-EFG �
]8a��a�����	aQ����W�'-��N5�-xUI(:���<5�5����tj�3����IQ�E>?n�2=Kf�V��hA�������&'�D*��<��jU*<o��ƽ���B+��7\��ū*�t��~�d���ű�Bd���;�޹�n O�3���X��+I��
�wc�w��9yۈ_��@67 N�K�7Iz������T�7��fU�5GYB�2�mǔ�u�DC���W�N(��o�D�K��M��t�խ��gS�e�r��<�����w��R�PxL�]��G]�����_J���5�^l�cذ��KQg z7�ߌ��	����W�û~�K��"�c�[�:��c��Vl�n�/=�d��t.:?װ����g�g�Y�
+�.��ΐp-��RXI:g� ޳U>�h,bF�:+$��Ő<�;��ف"!)/��5k|z����h��]J�5�	O�@���u_�������3K��R:�%\�60��U��YXh��Y /d�zh��U��C���!��K����#M�/!6�e��j�9I�´V��CG���<~vz�4tҟ��~����X�3W?�ŀ�� T��-��b4+�����e�D�|�\�Ql��_����7�֡wO(RJ��`�q�A� �����֖����B�ZԾY���(Z�ifJ
�+w���\�s������A�X�I����W{���㲡���vxL�hW��V"�`q��:�4*�?�V�
ԷόQ#P7��:�#��uy� ?VN���F��~�<�س��5����
�����H���� ���D��Ǥ���_՟�;��Ǳ8�w1^]��9q}��X��`���P�f4�t� �g@d��W��n�Y�.;	x�wN��8	cY�2�!A{�A�t�)�
�������g �Q=7���z+��&��_��s �3�Fb�c���Q�]�m�#�~�F̣y7IR7�>~���� &!�#{�������ӥ�.�K�`NU��58��Hm��H}���CU�\8������3�s�g�.��D��A�]*'���m�
-�NJ�Ne�B�����8�gXjV'�>�>�����m{K\�)�?�������Ed��Ө2֗D��䡦�QRO�v$?�)3X�<��7c��^�Zt�3Ky1�
�ћ�v2���M���`o+��K>������;R�	���<�Uf��·fE��c=�3{�B�{z�OI ��>�E�*�KĲŏ	��)�H/c ��xa؁Ժ��b���ެH���N�1�sp���1f�ɾ:)�������}3�m�f�B�B�ߋH�m�������`�^�����i��#C�&��x���YAu^���;>*��c;�!I6�}Z�Np˦5AƑ�?��q�:���p4j���,g��y�RqKk�.��~l��0�wc�8��ನ�X.x����c�8Ai��cl)n��ָ݃�~�H�d� _c~���G�&a�'~7A<\�8��#��QAyo�6�n���]�:���˙���)� ��q�l�=7���M�k�-;`t�ok*Ѝ�7=����'+SN�VC��a��Ei���Ѵ�y��'ꄻ4����Q��0�B7ή�W=�2��:��ce!|hkK�YEXS^i��f���� pv[�܌�x؟]�����o���� {��������`�Ҫ)�:�S��N����n�o�wR�=iJ�@�ZnU�;W
����l�~��,�\�g$���.Xh*�qފ�E{�Chz>�𴶘�}zbW�xU/�^�c��q��6�dX�H	C���a�<��&[���ik>s��i�*;)K��I`N�3�GX�&O�0W{�m
�����Z!6�a��go8`SP���5	���06�&��k(RR���cȶ�M���D:U[�����y�SeϮ-��(�Z�!"r��>s�Vx�:�v�I$4�C�9w�6>�b�66�],���)4�e| [3
��a�q���k�G���oOI��x�re+5F��6�/}m�Sq��L�d�����d��M8(��eTo^�2A�{�m��=�QeZ,����ԩܗ�A�$�����lH��dVK�;�a����]2�0�gQ�rg~!���tKR�=m�6`��_���;�:���;����	ʥ vYj��B�����Nڬ�Y�-�3 )��,�,���C�C�d�8iz�=e�A�#��.Ƌ�O��=�Վ�ƴ�i5�ٗi�M��A2PW@9WW�a8���Q��r��B64���<��,o�~�M�?�B)�wN�3X�_����ŗ$�^��}m��¾�^����������Br��+FA�EEςl�ı��]����e�NL��\�[bܶ�0��
�����s�юN?1�~g �:4K���脋�7 eF��ip?������$�	i�� |
���צF~EN���kh���v!�W�`�N���C^�u�ٺB����8����4��� �n�?g��"łX�^��*���eK���7�wWƂ�@�N����n<�B?��n�LM%Q2�^VFI���o�R��)V��{�6�~�IHo�XW�-��"ߴ_ ���!}{Ls�q|LخG��RI�ht?�E�/z���^���QH�,���7�<����｟�־��ލ;���{�S��R�HcG�!���M!�8������m���%�6rAEA�秗N�,�R&�Q����I;Mh�g�O�Ie��&b�I��ϛᯆ'�F��N_�ʓ�a�7�%`�'7�eS��PМ䛰��m0���%P����*��l�ٳKFuf,_����	H�A"yyTG��f�ˇ�N\��#�z�1�hO_3n�-D69Q^�����{��q�k �.T�`��2:hd�;n߾y呱�ڋ�	�"�G�
�M�[� 5F}"d���(�hE�t����u��0�����[��uA�ȓ�e����s�F�u�4����֯��˙p�엣)GmD�2�'�G#�*����X�(a��t-^CM�.�l�s6��5��S|مn���G����)�Q���7 �8�ȍo6�ޛ�8al���������{�5{_,�1x��[�~A�Xx�^�Q>���l�6��[C�0`�2�H:V0�������⠄']�4�\"����r�P4��~^��4[��u�܍���?��
켬�;]U~�[*��
�8e��Z�c�_J��H,5CX�Hx(~Y���M`1�'3���f�l{:'�5C��}KTq^�$��T��at!ge�)���Z����$w(��ӷ��c����K�%��-�p��W���H:�w �J�{t	Q���lp:���xy9@��Giub���@^,�P���G{۾��ٚojt{(�a�@;mA�~��F�h���B'#&b��WD �O���>�_��"f���| ��i�:󕉜��m�\�4��4eO�Z�?�i�.E{�ɐ?�@���ʵy!Ӷ�,�IxlH�Mɨ>�\0��ٴz��BۿQ��Q{�t������G"F��2�
�z>�&�k����q}��\���~G�\�|�iF�#������(_홖U�*��-Kw�;��o�@�J��ca�λ������C��0��̶�#���$�>�u���s������?sVY~y`��P<�ު���o'�a�a�T!y�5:�P�5�ڄ볌�����įPZ�0+mK=]o,tR	T���Y�L��:^�te��1�@�*9e>�tȬ����:ڨ����'Gq�1{j��6�(f]h��_���'�t�L���(ւ�;pҠ��8���"���T�\��8(4SpVKf�X�jg�� 2)ƭ���'b��钱$��q����3��$�0� W��Nhv�\�ک���<�WT�נPnf"��PL-�X��)잷fgR�n:��ηRP9�M� �zd#;H_A#�����bs��e�9mڕ�&7���a���$�ηfD�Y��}<�_p�O�/�:U�?A�`i��u�/�q�����Y}�:T���(���Wd�@�5�Niv|����b	q{9H~���2m�!��-ND^}j}��%�[9���G�M�v�	��{z�v��(H<�N���y�(V��bҮ�^�l��M�'^�t�(وG1�.��Q�MS�n'X�쯙�����z�I	-���D;��@`���+���\S� -hE(���+�,�|�����L?�+��)�xz�U�ިMx��x��n1Y(�Gd��@����#^�����9ɝ��I�
/<� ���ٮ��Gz���k���}S����H[���_Z�d������}p��3�di� ;��ˋ(_7��Q����ow8�q�D�9��1v�_�3�k_�{�1�W�9���J2U{b�
�R0|�,>I�nQ�.ON�`3�@Ykx`�/�B^R�@x�A���e��F�8c���.8�X��]�)X8�4��U��q\�霦]r�-2n��ܔ��P�+xv1�g'����h�-Y��]�{ÒĮ�e�H|ی�gˁĚ�s�z{�8��[rwc����pO�3y�M��։&|u}R��`���M��Ur���QW��FZ�(yX�m��au��/�"a�7J������2�����F8m��m��A-)�}��Nڢ�q@�l�>�;>p=N�pUsl
G������Rorr5/���Q��n��\��������h��7{�����3*�,���"���1k/�j��&�p������g����2ˎr���Ok8A�Z��7v�hT#�gc���`����ɶ^EY�6�WCA7A��HFN�O�|�f�EhS�Z����_�柗�h�fӦ��<��/N�7���J�N*��b�ݱeodym0rf��ϐV�şh��ר,�\�{~�$:�|\���Ht���C4ﮥ�Ҥ���b壀�et��w��vcE��e}��	q7H��Y��+�d��z�8U`���OȍC���x��j|���O�):�<$zjA ��g��;EP�&
�귆#��4��|�7��;���"�s�y����2��4/!��B�@X�s��% �9b�v��d�V:7#g�Q��`���NI��	=~	V����V���4۵�F��̀�|��|�J
몀>�W~xaI܃�������WU]��8I�[���q�>,D��-��)&w��-`�r �pz��������Ody���L	Ǧ�]�폼�?�a� bI�JЯN�!#)��Ǯ�N�$ſ�1���^�dU+�T~��]�Ř�%���b`�f�82�fv�����u2TRm��j;7�g�?�݆eZ�(M�����|������`vLJe���`�� ͱ��>�%Q{廃TgkuG��Hb2긷���!>��z]�-��qNU���s�����ܵ���Gx~E��f���3�Q�vCglK>��{�#��;��-�1�Fw�:L�!=��^N�㣞xK���W ��0�l���UkJ���Q����:��1�(�C���	�&j-�<�<����x=�X�oK433I�Ư�ç���py�*��Մx���*w��
��uEڲ$q�Z	+�$��|L��޷���z�����ѻ����$������7���9�p�.P��w
�Z5��$��+f�P�oX� Յ!,�S!��c�-=��K�j�m�����`P�#W�D�EI�b�_�>w�sN-��Ŏ�A�='�K˺?�}������;���Z�r�Z� �+!���w�~!2!�c��e�lc/Eۏs#JSv|�Tr4��9+�؊��L�b��� /T*���Z%i|�Ѳ+1��,ՎN=��3�뻙 � �8�N��X�N�9y?�7�1TUW���;!E�t�>���
���O��3uXo'���b�������"JpK�<|ى�,���;eR2�����:���	��c��h�!�%�8�(>ܹ��b��٣C�?�j6	�=�N�`'��~u�����)�� �
�a�|6��+#�&�C0l��%��O��[�Q(�b�k���k�4�1áx�gy;.e�u"���>��K��Ad��D��Z���qf軙Im��A��g��qB���y87C����S"1&��ێ����Յ,Z�"�)���dawY��s�-j�ۼo0����7H���K��"S���!�fM!_���7N� ,/煆��p��H��8ҹ}Ю�,�JQp��j���?9螷(I�f'#�\
r.Ġ�������'Y����8��֪.1�g!�/���%�Z�aPz����C����#�"����
��:5�d1~��!��qլ�6��>&����q��;� �ݭ�Nx|Ɲ������m���E����ݥ-%D�{��WU�v��!&���8��Jnb׌��Ĝ
����=�H�������-D?��E�>Bh:Rѡ�C��N�D~��L=S*ݚz���t��s��s�}��ס?_.�M����.v{���A��ѱ_��'z�.��,�p��,UhD4��O�nT-�Sa�V<��}u�S����J�:��A�g��O�#>��?܀9���?�9�a��sLn������ЪQ/eb���Zc\�;�;G��6ɋ�n�_ffOd�����<GX7[��j
(Jb�rXHj����t�4�i��m ����`���VOi�n�l�|o7��f��&z�i�E*�sj1]���'cX;��I�Φe`�1���E�2��͌m�44��#3�Cs�"QQ��mn����6Ԝ��
H#V���ܐ֕�m.p��֪���[l�-C�<sV���t;G��F��/�o�����9��L������{�k���E��|_�7D�,���9�RA+��sӰlã����k�w�3�����*� {�/�>�F�6\�W�b��C&�
{G|-�BtN��f��������(� �.wA���35&�L'A�7r�)�&�����-��ȋK�&QD0�8��g��B]gl��5L���>��ٚ#J �W�{�B�I�U�rӪle�ͷ|60h)m�m9xYt��ʅ="T�fn�����	�C�*Č�¼�@T?z����v�Ɨ�5�uV�S�%%�R�J1�3�x�bw5�qx�#:x��c0
��O�Pn�­�Mp��dy�Y
e�'j��n5�YV#���C�ͺ�����Dޫ�ص�~���hN��D&���Y6��(�E�>3���FU��~�˩6@T�=�
d.��e�̍�H ;���#���}�6)wՎ�ƙ�k�I{�0��MAt��./@�MrAb)��t)�ZI�8��d�Q��6ϲ0:SF@M�/n���%Vh{�Zuʭc�v>{�dA�V����̽o%�QV$�"+�4b�4��7�/{\�3hwC;86�E���B�'�L͸���^��R�q���X�M_��8f����Z{_�Α9�Ţ�j]q��ӛ�3�����9bU=��V9�����/��Nx�'c��r�:la�>������@����l��'��C��l��4	jI��s� ��kUl�	��?S~��*B�-�U�i	>Xn%\�VL���$l��z"f <,9'�ӭ��2�4W�gZQ��� �	(j��q�1k���¡eܔ� >�1B"D��0t:����!"�=.��ܐz�񀋅Ɯ��,S`����Q�������[RD`&]5��c�b��IE!��P�D�.*�O��a<,Hf����G�yp���r9���<���ͭ�w�
�pQrYpHї� ��rP�9vL���|�@,�R*U(Z�yx��!�D�_R�F^W�NwH}�a�;%����yK�'��Opy�e-�˅+��c�I��dh<��Eg�*����F&V���(�wu�&�!/%������}0���B(�Z7�6�LS��q��v���kJ@=R�:B���z���N�'�,P�4���OD�$����TuGh�.Ȗ�
��g*m��04}�MQ'آ��	kT"jG��D�n.�M)�&V+�E�|$��㙖�Z\SM��]݊#�htil
�;]���GSS�w"���#6�B�@y�5��bv��(	�k��Q`b��+łPmqm�E���E��f�2��Yɔ���J���z⥝$b�|?m���L�'��3����'�%���j^.jDt\�fI�?�?���		����'�}no���"q�U�;e\|��K���شB��u�1����H���`��f���%0ɬ��HG�A}����`���[x�X�\`x��;��y
�L�~���Wb��m��D�/].>��=��R�d�3�R��L<��),M��� 6��ڞg�\؎O���D�A��O�"��Oʱ_KǧN����H�4r^� �:#��gѳ�441���:�T�vV�����ϠC�Q��I����v�T~���n�b!v\~���(�/�+-��H�4��F��d~�E����([pM���V�eD��q��j��-j��U؟�*5�v�����0:���+S�v��RFE���~���ϧL�}p�Nk���Ö������Ԉ�C�lb�3D�V���B�t���K{�	�9g�>d�W56����ޛ�
��,�~\��ލ~���&��bYЍRd��:��A��F��ܦY�@�ou�;h��'b7Q�v��Ce�;eB�J>��@<;���-�^���->���nʚ_���\ͮ��#�:��z���P<���m;CT�,b��)���y�i� PӬ0ĸ�9�:�=�¥o��QU�E���~����XA��>���-C3�5}�bO;�h�AAx��?U�!	����c'-�:�7U-�v�*i�P���A�j7��^�D���H̀g�p��K�G��y"���(d�"y��ي��XD�H�%�|��J�k��߽" h�T���8Z���ɀ���z@��Z[�t�u�Z��1��ZA>k�~��v3����H��1�C�BL�4,�BO��ߵR3�ݣc������r��%�Vi�*�`�؎ٮ�{,H.�dH�)��S��CJd{�F�y�L��%���;�-����{�C�zW;,��M�1�(� ��:K�g��x/��+��?����A��$�͑~h߄����Fo-�r��R����'kA��CdcK]���Pw��ҼA�I�֏�YO	����lY1h�<E��s�F����Rٴ�I����kR�Mů-k5{�0	�I�J���
�!��GR:�tbw!Т:c���ז{�i�=��@���uU�dg������ĝI9� P�v�j#�̙+&:����V�O�k��jm&i��$��F2V˧.ے_�3fD��G	p#n@T�!ǄǙ{>.�������ʕ2�M����r�ju{sF�78�w�D{#��:ΎnrWl���MS�/���	d�,��wh)��(����m�'"�m��2T�
��g�Õb�dk�������i�V
�%�x ]Q����wX��[I,��K�0�p�1��TِK�<��B��m]��Ĺ~���L���EC�S���f_���(�U��!��w�%�b��(�\ �%5�jH�)*H[�Ѐd�9Y��D�[�-�G;�b���g��5@4�]�}��m��1�ĳj�ns���:�(_Qm��#,ӿ�M*4����/�W��ޏR�UL�>�ǯEP��n2r������計vmx����[S��v�ךT}���g�ߵZ@Dըw�2=a�rSE���P=~H��%̺H�	�*���(�ʛ���ŕ*�P7�N������N4�ʠ�J{�[ᔼ���o|��W+�.�9���&�n��崷����^l����V��I��
�:޼�}t��I�L���%�B�>�1g�L,���}+�E���5��[#�rVnC��h�{K�i۾��ʑ��b����Y?�$$��N��0�������\��,�X���<��`����u��xg�-C�'l3��pK�/<��/ ���R�+���j�c�f(�'��/<~���V 9�s�i/��N����tha-�޶�� �1�_v�7�nSL!F)�D7`A��㤽!bF!�CQ������>����ѺKIш��'_;�F�@D����\��痐>[���Q*a�ޭ�L�S�a��@^r��k����	��0�� ��4hK8��Y
jf�����s����q׉��#�*	#��Q矀��f'�	��B�$�k��ā��\���U"!S�q�RRT��,Po�7�>P�)չh�s��1�T�d��;����;(�!N0�ܢ����`�6%*1p����w���f�Uv���0^uQ����d/���<�Ri����r����hv��3�k<S����#��j�������Ƅ�r��ȶ,M`�{�����>�`�ڐ���?*��p�������"+�}���pE�Hǆ;au�vl� H.�T�_�[F%~��		��q1ib}w���Ϙ�m[����&t�s�΃ ��}���R�j6�ٞq�������/�g+��L�w��0'�l#i O)��wYv[�L�iz���܇�K�y 3�Eo��*�W�)t�M"�����喤������0M�l�t�?���7�0�l���TC���͹o��^��x�z?�P�YHe�YW3~~4N�D:���<w�	�裃����A��/��'��L�@��vM�W� o�9�l2TWKR{2��c����:�}B�0�ě�a{�סŢ��3t΋�����$:�R
*-m
�����n���3W�o�E���M�g�S�b?���U��q���~�I�����\d��Ԅ�����`�(�$�S@�AIP�ˊ��tm|�d�9xBA���o����M���Ï��@,i��Q�jl����v�f-r����.��{,F퇌{�="��z�H}��y��ƺz�1���� ��c���0���{G��9�c����a���f�ۈ�b������4o��b5��-��q�m��`�!����,Se�B�l��;���[�Ĳ�5	�}�~�ɋ�^q�h:uà���#��XѠ��0�5��|7���,��m���ۙ]��n]�Z
�*Wk3�=^(�͓��0�$T[�����@�]�B9e��R���ʓx0
&D�s
=����/��a�B�l�Q�eC�̕�}����V�Q�+K������_��=c	�S>�I�ВQwQ � ��K�.aba�1����TZw� �4�֖bc`�X=9��
�ui{"�(��D�L�&&{��!j�/(nr�X隋ڗ�A��l�����j={(v3�8�2ڗ�����X�g�W��
o��˳���.*&G�~|�ڇk��7:PY�ოҍ���C-������,P�) ��ك]�0L=\�`�i֒+���`�b!��| �
��� ��O<%��x1"�Y���PB_�Me e5�}���/);>n=XP6��Z<�V_��a62{F����U�/ˇ'_�#��x��N{uّKF�n�k��mȟA�"Q��h]�v�i�U$�0���ׯy�)f�zڑ|�ߟO���^�yt��l�N5i�\�w��o���/�X��B#^�:��p�Pqː�
��}�ǋ[x{��-,�s?�_Cl��gv�A�N�4�2>�?��ҵز-��~~���|�\^�� ��,��)��o�1�v	�ԥ��w�B���	�v�^$*��XJ��O��	j�y�18����6��G��.0�P�����ę-[���k3�<I�D�<�\Zq�iRff��܂6�8����>ξ���j�g&}�i2� �������+�ԓ�����7�q�#ύ��̟��	okq�^�z,�B�-�t�?�'1�&�gȍ��}��e|��񔫙��������UvV�*�l��n>Z=.L��~�:?d�zZ�~����7Jxj��˘��Hs\B����SU=��R�������{��z�Q�J�y	脫>���gOz1Y�p0��9X�Vk�ZD�$���E;��>���)�9?Znt#V�e�>��Cg����)�� h�\y��d�/T#O>�o�D^a�!ٷc`�v|���ː[|ˎ*���W�B�賯�hW(�����(�ߦ@n�o�߱ۿ����@�M)��Z�����F����{��x�&[��%��_2�]���B�F���!���P[��
��3\��	b#`yM�:d������oz|I9g�@[�5����"��򚝷����b�O�w��C :=,P�ñ$9ni~����vƐ�-�"+��4�<<�5��D�ц��7^IzZ��9�v�gg�����G��G��k<IVQk+�$�=�3���>3C�k�%fT������朌�o�H9��;.��||�p����!�M�����a�a��R�Ӻ��[�V���p��T�	6��s�,��Y�2� r�]�}$�n�ʬ[��5���y[f���֡�\ ]A[c
<�p�2xo�ꠦ���1y���X̞��)��q��ڀDpn[�?���.����0xL�T����&~՘4kE�;�&Jc�/H !�v;=�lֆ�$����J���ұ'�;H�ؾ�`�p�И@��
~9�M
3k>3W_��y��Z�i�?3Z�C	�.,o�#�٪� �m#��κ�ъҘ����ɰ=/����F�ҕ�Ю�?|E��3w���eq��"	G%"8������<e?x��k@ѯ��U��ȇ�R ������&�k4�}���_��3����a��ԇ,uћ'W-�6��:�:�u��W�ھ��G��Ĉ'�&`��<��ÝB�?}Ԅ��z�6�g$8����O��Q8��?��8"(�m���V��tk�C�5[6[(�C2�DL�c=�q)� �J4�̅�x򬗸��=Υi��|�aź�A�'v����@ĸQFۡ�L;M�����3��X�d*�9��9X��l���\�pTH�0�#�Ϟ *5�!�0���@t�G�4S{-a�5)��
��r��Ӻ��0I̽)��k�1���$

{:`��k͖����aN��|Hȟ�a����'��t��F�����(4���+�,�R�IKڿ�J���
\���������� $-�7�֖ͣ�D��K��y��5�����:_?@��jųi�5y��ti�z���~�u�6�+��ǌ#�M!��%r��t���Wr 7a�3Z�K-��M4��_2��m2��}�T�w����n���z�M!�Y{�b�� Qi:�n���p���ͿiEf,�r#D�I�a؝�&�E`Qy� 9w}�(��A5��]���U��F��g�epV���&G�kO���j�K R)�oE�G�u�'�4޹�/e�̂� Ñ_���ˉ�%�\��4�4ƙ���m�մ`:��ⴉ�J<��`w<��o1<�x\�iJ��m�����1�N����z�?�*�Z������V�� �"O�R��S� S������EN�����6�/�u��>��s��+�� ��N]t�r�S+(n]{�L��UA��A}0�9Yz���`#��A޸_��7Z�
p\�-�� �+(Y��NeFWLA��R��c!��[h�x��~we�������7�,)���b�i��6��Ь���}f&������
���w8�=��b��w�����X5Vw�a�4�v|���	nL#�k�V2$+%�e�,aX�q�R//��w��Bgi�A�t�1@������u*}:;�{��h2I�9�����-FY	�_��"G�z:j�C���Ġ���8`P��ij��K��!m��������k���@�]6�n�0����\�Ӗ$�y`Û�5��n�m�vi&N�a�ٲ�n�5�p�7{=�l�s�����L�6��9=q�����'��p�q��j�gM����Os��ӂ�S9��^��+���9WZ�2���l$*s���6��4�� ��G ��#_�ձ��/�J�/��*�\��j���7H�s���R��UBf�S��k<��̂�L^qe�O�[-����UL3���:���u0ҒW��z�xS�ǖ�_���aaʚr�˛GQ ��J�2Bc�HD4�ۻ8����Y]h�%4o䐃�Y!�B�ja��!*�^O��_�X<�Z�C�
��NO?W�j)�R"�C>�k�"���a�Z(�O�<�˾6�+��_�D��=��;?@R�vȴ�8A��P)��S}�dܪ�K6GӤ�ÍUXI+��0?f��8�+��F���O ���1ƻ�揖��޳Wk䵤��@����4�<��Ĉd������uB��-��ș��=RC���o�_3�]�l�\�������Z2f9�ƳMDP���>#[Υ	�����;�d���{TXs̼0���-6_����W��_켝�DF�щE��_3@iF���G�6eA�^�Ŧ�G�̇�@��l�6�
���^�I��ni���a`���%CoE�.�+�Kڡ� ��a���&]J�|���U��b�*4����J'WU[PY.��~+nj��H��F�kV���������PFM[eC&pr��N�\k�7D"p���IF���!��We+P�Aq��J��<põ_��P��h�	���W���zgJ�kEʦ�����J�aH`!C�Q��	ע=u���ɞK���������Z,"�5E��o�3�96�P��L�n��'{R��s������(����P)���L���B���>���\����a��GdS;�z~���8��$���\vڳD����X�ƿdeצʹ����=U8d1m�C8J�&�Ȭa���Y��l���$���kP�����T��4���z�=���*�H}��cc�pt��Xc�xV���B�sR�G�m%���h��w7Sjr͕va�t���� ��(�F^�w)n�]�3-X��/F�6����ݷ3��/��P
N�)/sr�R���+̱'�tsc9Կښ����4�钅���VC�qi���C�9r�ʰu��
`�@�v/��j��r�\,�2���;�������H3ӵt�J?d�̲C�%/�x��+F��Қ
����;ij5V��儱j$�9c>Kq^7 ��M������t���;��j�|���Ky�K3�H����E  �W�h�n�K��Gf����FHl�dK9˙��Iv�2��^��}�6�V�!��q����\�tzp�~Ġ�e��C��»��U���c"Lw
���j���J�^��:� �+k����?X��1G�d������s��B�u�g?���k�4��=�����i��۪�d~��>[5JF<�L�M�����d��y]��r#yKH,�[*����>Oz�#�K~=����7 ����U�+�/5���ݫ�d��0X�)�w�@�ƿ��(��R%�M,`[�ء��{�44b�
c'G �)��ϊȰ���`1ɦż�%�L�c�N���#q��j���:�$Y ژ��	�Y��=��?����M4l��ˡ�+(�vS�^�y/�t�!��!��v��|�<|�,\�;8���G��c̜a�vX�F>���B����6?N�?�c
�7�5�M �0D:�r���)�6�a���q�Lj�0&g����?��(���N���0�6�����c砣���у��E��2N9I���\��R��
�x�G���6�t�5ƴ�y�S��/�w�ͩ���!s=����,��jY���\���]�O9�Wx2�_�F6[��Ƴlv�-���H+��-X�	s`z�!=�*ҍ����`haد�������뀜��-�^_�%�zd����[7��)0)��.�d�}�����>E��CY�!�R14}���r@� �%���]u/��'��ҞN������	�8]1y���u����H�u���$��R��_L��o.hz Էs����B�O��;��qgK���4�C��p��Y�=M$+��q줏�7�\b��n@T�*K4Vo���◥���̫���Xkt��H�ˡ=T��c�e��Yh���̢^�,qx�\|����1�#�-����b���aѢ�3վ��ޤx޴��RZ���6�u�YPQ=�ʝ�	�u)I�P,'H�g-:m�=�v��'�*�u�ҹ�U� ���}K���GO��6�@���y�՝m�if�6*2�Ŋ�H�G�����3�"H�r��3�e�f�ވ�5꜋���d���_6v�d��.�d�H��Lր��o��?6k�8� �Wï��  2�z���7�7>&bjc��{��s���t^��c�7�W����gʰ`)���X���r����g��?�2J��!���%3��@(�1��Q5mk�Wgs�ĉz�ͱ�M�Qa+�F�=����m�lPO�@��2��h�o܈����Z�გ�TΜ�sf_�z��6���� �փP
es�6��Ә����ӟk=o7�Pwғb/�;wR�	?�C�� Q�C�f��S�?)Ũw��=�s��x-kF�1=�i�.�*4BD�Z�ˡ[�;�+>(7�
����M'�uh���AO���� ���.,C�v�8��D��	pK�m@=<$ҺHmM��r=t�.�}v��8��ܫr*-g��A>����Dz�W����8��>p-��	oAX(|���Lygte�'e=�Zzr����VD�/6�I;�uN������h��
�	�[��Ż������ �%��!%��Oy?����o�p��n߀Ǽu��Δ������q=���xq�T�;�w�+����Yl{Y��ǟ{�����' �i^r�j�D�4��`�f�c������Ru��#��(Á^=v�m�oi��R����N����V��<Â�ca��z;�y9�vL�d���x�¨�D�ι��M�FZ5��X&���\ZA�G�;�$�!	z��[A�=�A�f�6Z:U�|Srr��������u}�+�R���}q���х�xU'.!�3r�F�c!&����Y�9��y}�ͩHsU� �փs��a���:��Dn� ?I*�K���{��O~
��)�9񑕡?�יg���)�(P�/v��3X&YfJ	L���p�"bn5��G�`[�9)7�b��a~C�S9&��@u��q'������eŎBr�]\�1(z���ARܷٓI�8a_�ck�T��b'M���6�j��纏�U�곬���P#y*����nгgn�<a�Rc�t
K�du1���P1dާ�3��Y:��-��=�[�gS_��y࿛� �k�DN�ϽW9ߋ���w�a�/�*�"��-��wBm��Z؄���� ����ə��I%s�AR��xv�=N?�i��<�t��^E��
����Y��A!�P;�OOF�'Sٔh�5�^��N�lW���Q6�w;�Jkz�'p�4��z�?`Ι\����"�Z��@#��`������`R؇.w2�H��;�u�҉����J��Jڂ��>�U���E��ߵ-�R�8� ���^���9�	��xe�\�̶��!ٓo�q�**	�؍�� �!�>Br���� Ҁ�7�������%6��6�P�l�55����q��#�v ��_<�΍de��ó�õO�Ƈ��)�/)!%�趸M�$���t��x��C�pY���oR*�@d��Mws����T	�5�\��C�� t���Ղ�	�����BKB�S�W:b��ᘙr��]7J���d�
�-� Ox�s���&L��4 �xGZFSS ��k]�a]U�4�hd.�_���n�v D��`���d��Z�B���ύR��W�q�aDk��]
�
���� \7�� �q�g:_:�e�S��D��<�`-�/Zӊ#����!�Ժ�������l���6;G���r�ʯ|;��Bޕ|Y��k`�&S�*����b���}���g�/����Bi��+�E�G�(�ѣC�wŅZ!�"�vq�X� +���	nV�����!�N�w�r�f3?����ٯ(��+��Fސ֡��T0�����6��Y q��x_�u#;�/N��_���^�\�u�[� �Ed�z��r	'��.o��0�b�e��Ў������~�=¶�`�O(���Qߎ�Ѻ��K���d$�|��`�����8H����p���Ŝ2��u���8y��V�5��qI ���J�c��:�B&l9=�3�����	�*P1�D����N{Y��l��"��k�Ĥ�4It洪��lT��2���MP�JOo�έs�<e�	G1;�6�������IG�|SQ�4J�{�/�aI�?"�Dҕ�V�8�}�;,Oܞ��Z���=�g_�H��w�/�*H��ϳP\6/ypK�N&����:F�%<�Y|%-����l�R@$�}u
-����)���8P���X���/������6}Φ�ސE3R��;�Uv��,#�@���e��;"�0Nk�HR0f{�8L�ƂwRa�(�25�R�^�O���S�v�e�-J#Q(�h�Q���9��:�ϙt#���Ҫ62icބ.t�7t�F�ZG�M�
�M�3�TQ~�C�r���m�D��̱��ir�֚�u�d��,�,���ʮ>��^+�'��·a<j��� ��%����[՚��co�vJ�OÍa2��:h&���SD9j�!��ȵ��lUe\HA�2;L>�!F���4
ҸKOaq�[\|��_΄80�'z���i9��������]��m٣?m`�u$B�{�~���6�� ��I%����6N��'m�y��Y����d�ݘ��ia��:�}ş��뽛�F~��S�E�,�a-z��O ֐����Pۊ���{;��c��^��<������Ul���vK��^:ͽpݢ}ު�?i�-��
c�>}�P蒹y��{�W�L�GӉzЁ[Bs�r�����uaDn��+���5mIrS�\�����LRw�|��s��9b�?�glRf����r�}e�@k��!י�V�`�ق�7Dd�Z�6��;�Or�,,�ٸI��^���M�2X8ϝW]�x��5g?w�v/�1�e��BCr��ݵYx������H�͏������J��O�;���A[N���4S؈#�&O�SO%�ӛ�f]�t�u����=���M�]��C�����s>�{
)��a�*'���r�\����܈[32!sg\>���yN��0ԉ��L��q�D֙���O�9��`�#�0{;�9J\[M�V�/W~�#�T��K?��6Q�T��.N!m8�T���żh�$ZqL0�g��y�1|e3A�,��ye�r��`^����m�ޡ�ӄ�#��t��%�BRN�B������9n�t�G]�n�:���}�x���$܍�{�y��S(GF�ű�� ��ر�	zU��h�R����թ�'�0Bl*��vj�����q,$ā-��6��!����y=�.�2]PJ�[׍N:%T�a�gOwk�W�jC/JGOם��{�SV�U����"����^%����?b�a� �12M�:����VC��M�`���K�a�'(�6 �Q^��~5Aș`���1�].x0�BdK5(��~�� GW��8�vR��<�'��,�~cG���'���v$���$8��AJ�Z(��Y��'�y�l��M+E��SD���l詽��`�y�o��|{�)0A���Y�M�%p��J����Vԃݙ޹z��03vK�k�nU%-<�?�q�jJR�8�Z�v��84���"7z;PX[���~�����6�U���,hN
���1;Ku�g,T���'��ũ�V$�(ңz1����B�^QY�N�g�1���ώ	}X�dO�H`�rV!����"i�3�qъ���r<�@��3bM�F0��i�ӏ6�{�,=✀�u��w�/<������Z�7�=�9���w�q>;��/�Z�"���B0-*ܖ��_�Z~� ��%Wښ�a�)����ܚ��%����F-�b�w	>����/�}�$_����sc��(bCǍ��<�+`b���$Z�3�t�É@zzeɁ ��#��VAE�E�>���|��/7>��vaX��p�[�8�w��C�H�����T��"�R���/��6�h��g� J���U�ַA��u:>
�y�>b�D���e���G.��}�!Bdh�����ʺ��s<#��F�
r=��_Bg�y+�R�w���M䯑Q���ʊ�l�r.ul�ʵ�KH�@�1>��<�� Fd,��E�������h
m
%��}��}��5 
�q��s���C�s/XI�p����b��k
��t:i�
�){-iXD��N��GI��؁�E��0�Ȳ���y��.�Q ͥ�i�ӡ`�y5';d�,ԂPKL>���65TFݶk~�wR�J�%�n�O{���[�\�O���lb���4K�u� �G-�`c��:7<<�سx��,�8�Ɔ��ɖ�$��_��O���4�&z�t,�Y��M����c��&�B�f������c��5�W���(���ݼ� ���i��_a����������"V�T����̺�6T.Z�Zy��}
 ��,;�G�Kl�^�ebQO�p� �_6J���n�˻`�"W���f�ls�����tX�}*���������I���B!&�eRB�zKe�+��!	9j���a�^���P,�u@����F��{Q�y�(:߉1��yٌ��`��LFrY�)�ոs�$�E+�c�����Y䬆H��ui%'�1�(>��o�l���)m�.x��|�X�/j�m�;��ѣ9�v#����sd��}/b?�f&��ޖ�#/ū���[=�ۆ���Y�o���=+<dt9V܎��ӧ|��0ϕ�e��&-�O�90�:�F_Sֶ������F���vġ���f.2���p@
Q����s��T��r�?��Z��}&X�x9��ϧRB?4�5��e3v1m�����u����Z�-Ԧ9j-�y�"���I[�a�ٸ����~UFJ�VDG�P+H�u�v#�^�0��߲И�����97�)�?��f�u2�4>u]�k�� yr����U���}�Əl�p���(j:�FB���~QEvs�]aMԍ�@	�\������T�ժw�I���+�+�I&팆M��9��W�;�BR�W}<� �Y�Q7}b��n�?������XZ�V Q�,He0�0Zф�R�R;𦚳�O��` i����)�<ͫN��X��yU����#���,X@�/��� ����@����ՠ�@�����)˼�m2�U���t���y����J��5K�����y�h����Xa$&eik�c4�f��f&��ɻ���L��?������Bt$���Aί���H�F�ø�*�&�O��Y��s9�J�'�p�4<�1���??6}��D�Rb��D���u[ s)�M��f�1�ր�W3���h������d�~������G�F��-�E0Q��~����h� ��Z�=��DNq'#q���K�$Pݏx�`���c��/�Ay��r��ˆ�!	n��ؠoRp
]!"�J��S��`oϕk�ą�pz(,{{3�_�y�wC����=k�g@X��f"Hi�먀<�F9�f�njO^�qŐ�"p�vy�^I^!�V]O��O�!#i�	���k��~��6��y����K�r=�'�a'�H6_�4���oxz���������r��j�� w�^5���(s�ɗ�����h�A�'t�fw�!�|�;�2���Rܗ����3�Q���F	H(�FUq�����I�
"����-�����.d�h�<�
��擜h�H�@�W�^T�8�.A�c<��llW��K5A��h�x9yȎC�9b�[/5���4�(�8	���G�S^#��#����%�T���x�yR�"�{�ۓW~Rk�w����A}؀s��,e��H�s~��;O!XN@$�%��{����QC�N��4!fe�k0&��8fq�qw�[`(I���*s���M�'�!���ONw�PZuE<[����u�h]-�xů��ݑ/�G����S�N����K����o/Ә�>
/=�[����.g���Ω��Z�{,�'��8���z�mm]�M���'�"d���s;Ei��W���2g�*N;���4(�w؄q���!W ��>AhM�Fs�� v�P��6.�n��ӬX�FFґF7�Q���k��q�n�x�3*8j�`AǰJ#�0h�]�>�Yg�2I-�In����x�]����Kҿ��9mb�Ȯ�6����U�����_4!�} �aD���D�lc=��A���*�Eڎ?��7;
��������FC�.h)N<�/��r�/P���b��1M��+����t��ɳ�j���
��Kf�#�F���2�च�������R��D�>�:C
<߁��f����P0�8A$~ ����h����"���[��o��e�k@7&] �LXW��� |��@�}잢�yGup$�cu_�)G�I�j��d-�ԃ�~�A��T��kN�Vv�r#�7���cw�Ů֦����S.Ǫ���ײ��(�a��ր�+	�D#�Nѧ�70��Ǽ�nE�On����U&1zf�U��i&�VWE����ħ^�Ca�-.��'�%%����I�RxZS�IC��6�\�ޏD`��I�6=5t?᎞�=�6�Z��kp�[{8t��VpQyH���T%�2q��i�*����y�<�h�	��ygZʟ�o���踚w�X�gZ�a? J'b�����e��x��:�4����j�#8�;�"�}�p�R��6L��oS�n:$��)}�x>���펑��Yo��y	M�}\-�AR��li7'�)�j�V$F�ǅi�J�n'g�g(c�`q��f��t@���6�Zy
��->�������
�Ű禫�Cן(��S|��./�,��G�\�X>v��c_�TP3 ��7[1��+g�̖�	����S�&U����0�x�h�E�-p �|o�R�QOr ����Q�q|ӟr����H��-(����W�'�3�=ߢV��160��. +(��D*��[���8[r�#�K�4l�J4bI��E��2���U����B�� �h�A}�{1 O����3v���]���yp~�fX²��)�P꛶)��p0�>�kE��ɐ�f�ͦ��G�_<�3��.?-h��.~��e�4w���ky*�8�F?j�*����o����y*�,�ǈ�p����%�>�"[r0Mb��Ν�g�S�?��~��oF��N���Zq���< �O��ԩ�qig��.=5(r?٦>�P��,H$\�o��߃�[�E��β]���5������D&����2�k�\*L��踧���:t�m ��X'�fL�$1�$ӊ�ղ���5@_�qe��kIX��7���pD\�6��O,>՛���W8�)k2����nXp"����U�!�M�`l�y�S�E9;:�ű�h�ů���m�m���ɍ\���3n�}ff4��u,a��ź���-bJr����Vn���(������p��rs���䒒.Կͨ�bLw��%&��b�*���x��k��8�8܊�^՟R��嬷Un��r��E���;8�2�n�Vf�݉�������8�ު��aYr:��1x��K�����=Bh���DG�Y����~Ҁ�g����qpVorKh} _�k�G��gw�ɇ7;A�4��B@�[�\S��o!��l*Ė��m[�8�=8�������lw��KZ>�4�P%�R����b���?&Ҡ�-[���`*Ͳjq��f��i�^w�_բ�0���B��ܶ��2�Z+�~E'@ ���3͐A!�J��Ȟ���ܓ�A$�GAQ��a(�����3�L�C���K�����=O=}q�QN,Q�$�s,�!^�e¼�ӿ���� A"���d�oR�#>*����e�m:~4���KЮW�Ύ�'_o�R���
h�Er�D ��-��"��:�������s:�+�8�쾮����� ���xE�C�8�������\����G�E?��,l�e�E\�	�H��$��Ep����Σ;�w/�~|�/�-p?N�u�P�jP{�o�T}��|b���^q5�G��с���9���sv�c�B�_="�6�A���O� 2V���k:��o�1��z聟�"�Os���|}b��T�4FA�1J��{uX���Ɛ��tK�H>g�V�13�T��b�_�WJ���t�;���x�}��*Tu�9����2'��#�� a/��D�8�~9]�mg	z�H��~J9B6H�'|'��xcD�?/�"/�����U����1���q�N�Icl��������,(ُ^|,���]jD�k�n���f����F<���0��V�d����4%���9�d�F}�?��wma�^Bф5[�&a{���Ť�=d\A>��_�rn�tSl:SQ�����������j
����Y����ϮJo8�{huў7"s�Bhm����R\�8}�K<TJN�_QC/<�O{Ek�a��Џ���2�i��ǵ�����K�����kܐ���g�/`��.Hi�p�	��.�^�	����<�>��jK��%^M � �X�N���@H����۝�o�RK�u���zůe/XF��-*�������\� ��MJ���I�ֽ��� ���S :Tf���R��(u��|��ʇ[�%Ž�g.�τ@9V�b2t^>&T�#���,}ּ���)-���Ҙ�F���)���bU���k8ھ��/�r��������x��^��Z<q�$O/{��G��RV�˹�[_����х�]^s�Z�6���o0�vNg�e���9���7����A�I�U��+��;�m�F����G}O�#�M@�x)�){gӶL[i;� ��*�ϲ_VL�u3��ҾR�{jRϖ]��Ð['�~Z5)T�#���~�n)��?�=r�B� 8�~	�ؙ�A��
�����Vӳs�"��C/�t����_�ՖA7�����JLM��?��^���P�?�<��zj$����'	�i����@�8����`B�W����,闋���b&o������r�F���g�V�
Y�G-LçE��3|���ٕ�_Y�E���+f�z�D�wO�A�ᜰQ������Έ��IڵYN�ҽ�YE~ gZ�1cܢB���'��<D�?Pi�Ԃ���F��NG�Ͷ,�|��!M��e��`;>��ů�K�|�3ݵ�SyC�qaOO��`{Yf�UR�~ �D�1̳U3�\�${}*�jG<�������OV����9�u��/q:�ԁa���"�5�P��T`���q�Ah��U� k��Cp�E��j�:}lI��&#!�>a $�ӥ|��!#����Vg�����	�.<p�r�hC�������P}=#LK�97���}��F�-~�l�?�~k�K��v�p��X�
 }��`�^i��3k>����U���`<��@痝zv/����[q����gT�&�R�(��v���0P�[o�5��"�U���$@lAG�:ᣳ�?}xo?+���u��y�-f�_n�5&���U� s�,v���~���y�x>�u9q��X*�V�c�֎E��p%�H�%bb���v	�8[ђu]�$ _(�Is�S��#<YSf��	���~��O?�uvW� #����3 	h_�r�V����W4����D��I��� lӴ��D�%#��>�x���a�L���>a��`u�:Z���J��V"��0x$�+C��u(��}	1�����鶦�i�� G��W��#�#!y��-����r�VD�v��Ԝ̲ q�$�����RcɬO��>���������\r�=c��$�->Ȇ�V(���]k]PS[�j��Y髃A ^��jz/�_�X`�k�0�`����c�6�w4,���J�nB�|�=b��!��!ODS��uP�1��2F���iz4Y:���"��M�Ns��q��e��VL���x[.�Æ Vǳ�`�,�Ъ���=�J��y��"C�.=�\%�X�+�7L,�e��Ļ��(b,��᥊�%�;�NUrǰ�G6�'��yu�B���?��Y:���z/u��_T�9zC`;�g \%�ɛ��s������W�4z�z>�E:��,�(��&��m��F�b��)��R���#��fr�R�`��ԧ�rBΚ)�p���8>V7�9�s0����<�k]<��ΚJ�w� ���%�<<k/�|�=������lO��n����/�l �2�k����O�49����*iv^�,�%�`�xY3�aE�.��
��y�.��_0A*z��Y*/&�MZ���_�Z{N�{n�
�TM���|B�N� V�����du�ei���G:�r��E�n�S��}��䁡o
�:wOͳ��n����е�H-!�Qp��~/����&��ad��p団�O �x�{��
�&�P���?��v��E8����߹T���>�>�b*��Fʛ?�?�|P��~��O���%�����.5tB{��?4S�&���T�����&�-[e.��#f�Ps%��RGTصA�T[[]�Aq����*~��U�x
�*�Su�頻�z&���U����z;
O�:}ѯ�h�[��p�z؂�g����ׇ&u|�ɛ%C�V��ri��g��h<O\�L�-��aH�)��'����l�ؖ�Z���-ЖJ����K��=�Ѐ2�.*�v����'�x�$Wi�'7���Yc��t��f�w=���0B@n��+�;.t�U����C�bL�.��w�b�0�x�]�I�Kǯf��D�"&��r�e�*�QEG��d�L+;,E\�D,��̶��,��� $�G٩2/��#�so�		 ̺
��Vc���������s�P�A��p���a�"?���v&�~8��\Yo��(tx$%TǜI����r�Gu
m���'�h�qmM�������15>w�ص�]Z���L���6����ʨp1���9�B{ϫ ��h��4�����y����n]N�-�K���!#�$��D�z�����E$�@��З��������;�l���,N�2'���϶�,Z���1��N�r�����ĳ֦މuW�jt�QQ[1)D�oOZ�j/�Jp鱝���G6^�����8�A�O�ks(��mt���Y���r�4��tC�XUe�R�2��M�Ёq��h�I��J=\՛�6�X��A�ؘ�o�Ȣ���(с�C5)� -M�	d��kO��b��;�;��S/��Ws�"���3C��|���:֩I3F=J�����d���RػoCn%u�#��i�য়I�-
<�?�%��+�%3���
�ю��)��~	�EL񵔑=�,�z��ea�@�0�Oƈ9Gii}�'6M�T�9���ϫ�w������ȝ�mOx�,A�ݜm3�,N�$e*<�|����E�3�(<<?�(�DC��@4Sk ��������cO/�  :y$09�\�7��߼�X���޶-M�9$��,Ls�ja;'��iR\�
�r%b#�i�� 勳xfmc{/�F���0�"��5�44U����ۂZj��tu�B}�����;�f�{}Ykr\��x �}	צ��U�{�G�r΃�J9}�������~�%$T0m����}4"�- ������ ���?��K\��N�idG�O����F��_����{�&�5���NF���h�j���L�G�ɴP��o�}u�}^0�p����op�Ֆ�^��f�\�3�S�;�0ҹ.]����z݄��9� �;��%Tp&��_h'����q
Ď�qm}��f]`H�����h�|�ܦO9�vQ���L�+�7*Y�|.=]�9y�mv����)G����w���4"O��;:���r�fgL)_�{~�+���c�c�F�U�`���L�U�0RK��7ģ���Y�oNA� �o��n�ͺ��R�8�gkJ�gq��~2���	����mL0�è���S�CT��2��	Ş�>��5�J�f+�b�t`'�x�ku�y���}�*�`"��jC��9p��kQ��mU�%*ő�x1�q��GT����y{�`�,�OZ�[���>��8��A	y�N:r�ػ@O�ԑ
��$�P^���U��'��6�N�E#]��2�$���;z�Q�D�m��3�/����_ǜ�ւP\3�ѮC��2�2�"�IU�<�ә�YQ��Xi��Aª��b~�"���� �B.��v�C�1�[zǄ�?
�7�XL�B�eaԻg<�c͗�KҎ� w cq�!\�;`���������Nfi��<R\4 	�^c�*�"��o)�K1�v��\4�T��cE�tp�"���'m/8��<�#8j.L4�y���dx��%�2�����5u�V��r��-AN��R~&��� ��	�)�d�K<�ܥ����X�߃ ;��!6��@SؖY�0�q�k��|��%S+Sܣ,z��_5d�_d襭3Λ�f���_K9�ܣ�D��g%�70T��a�Q��niq�8��TC�(��]>z�'�]��U(R7l0� �|�c<=S+��-�rӞ���V�ђ�6d�;�l�u�9����UIe��+[(��J�@`B*�ѥtB�+SS�w�`1���ɒs���k�Sux��6Q?�f�?1J�iB��8�[�F<a���7�PG瘒f�K�zw��o���)�!��� )�9%ir��a)ד�di)%2��櫢��	�sR!ʨDCg|�3¸e�v����Wt=��@��<>=�!6��{���p��{%K�=yf����y����~��>-����bHb��:.V�X�D�U�k���P�>�����LW�)�w�L?�@z.>��E},�[��R^-��.bf�%�`/���j�����O�֕�\o?������׈��^�<����uI�R`y�皥'�h��:�N�d�|E���{Yj�k��h��U���D��[Q�Շ���������ݕ�
�Y���}�M74�~&�ɻ�1u�^"^-���>���;��)
���>.�br،дOK4������5S�YTc����d{w@O6tϓ���a�_�L��{	(Q��PG0�N<�0B.o�/�뷄p��ȯ�� `M�\��u��g&?��$��XF8 8i*]��P�u�n��!Ĭ��6x���{��F�=J��CL���`|�9�x
�I�SV�n�!���$��8ӚKEM'�xt�E�Y]8���V�$��-�j�)-&�/d*S�{�7�Y����kos�0=,9��8�Z�?��ɬ 2
|u�k7[)��|�Xfu�\#�� ���> ��OF6��v:��$��َ"�|�;��%9�Tsd�N�����"i� ~q��,[9;y�j4�>����PV��T�k���s�s��.�A��z;��ښ6�dƆ]P�����P)i�X���6���$�}��\���W�C�ub6�f�����>�wٚ;��s��Wk���E	�7A�(ȁ6O��n�B�G_���B�O*����
'g9���ȹ��>ދ�s�+�@�����ӎ��/B˘�
"j��Xۧ���	p�HS3!N	kÆqɠ�M��Ӆ�L�����������^�UI5¹�S43���s�5	��GA�@0!�c�If�xW�H��ho�
Rj���Z-�����&�7뱳����,��/�zL��m�V�Qi�`U���y�/����=@[g<E�ｶ��LK0
� ���hw��g�6�vQ����U���]�g�}/��cy�?�l�ԆT4AҰu}"���ڥ!Ϯ1�Db�.�9���,��*(�D���	{�<;Q�9��TZ�Fd�hL��$�06����mkl=��^�Df��\�cen���2#{%�PH��T\�#�/�$�4وkbn��Ɨ�v��K�*gx��ۑ�fZ!��t�>�M��A\��^������'Nx�n��wY��Sq���'�Hr��_����[��<�o��0�Ʀ���G�Mƚv�<��.�����Q���
�W���߰����57Hy(y#�0��,N����B�Mj���Rv5��f��fz3B�WOT��F��O�`����+(j�:yi�?���U�8.%]�b�����C�0�?`T�{$L&ܝ�D�:��{dM�梎u������aמ���_���j���m�Ο�c���/�ڙ�*��и ۮ��ь��le �ڋ�;6%L�R!s�"�2
�"#r�׏1H5[@�
�n�ˢ0�"��oLoi�A�[ ez%��Yzek�U<b��'�
D|OL���A?���g�!0�O��>�� q�^�c�Z��Т��$��Vv�a#�����ю��P��r>@m�%F-J�hV��'���|�����w�Ebb���Hs���X��i����(>,<�B`�r��7+>�F
�{�Ď�a�:�#sT 6��&�C����wF�����H�	;�X�*��-.�z�����B^���8s,K�^0~a+ԣ����w�y��_�ك��IJ��L���05b����z[�y��o��CE�8G�6k��bǉ�j�*'._o���}�ղa4U���й���'O�a�4p�;Ǟ�h`�Tj�^��S �w�i�B��u��G*�fB�;��m���kj����$�)l�"�(��1�$d���$Ο\�tc��/�F����Oy�Y����D���?��0˵�]��צ=#Y���ny��$��R�\Y d��A�Sg!��#"}d���x��&�T&�l�7�7$!/��	k�X�~�bz�T/n�&���Z���4�p $��L�j�yʻ���YS���ݙ��_�i���T6` ��u��{����˳�]� �-��F2hӸ^H��������s�S<ވ/��V�� D��\������hI@m�)X�Q�b�~�ޥ�r�����$��wrG+�o��U �(��2������w���n_Yx����]���~~;��F4/?u�[8�Ǐr�mYj4��y�k��w����Cj���xq�b���5��|_v[��N�A�2������
V��gP�ʦE�֬�hE�) y�+����\��A�{�Xtג9kp�	�tZ4B�f���c�7E�L&�uv���4�GO����﫦�6�m
���d	 ׷i7
)�8��IH>t�=�琱��
��6ѣ�4��0�p|I�IC�ZKPH�sV_ý)u���X/6!\4�U�M���K\΃��m��y}�*O�uOE����-|t��
�z��V��t�!�,/
��d���X��=|h�Ɏܵ>�q�<B��.Z����p�������n@>��?.�O���X�ۘ�U�b��f�V�/�[����I�]w��{m!Ű4S�E�;��vt���8>��������Y��#���:�5��:z���D^��Ka�7?`O��B���F�('�GG�u8�U��ᙦKD�)�$�DQK�W��v�\��W�	�Xr�h���7d�#�e��&|ӵe S0tu"K*�Ƴ��^�Acj[H{���I�g�+*��Z[�j���H���	��p�;���DQ�%O�m]�%B���bWod��O�2 ?{�;�|��S��+����x�<'����,���l3�#�}k�� ܯ��3�?[^�7��Uh=&݇��kS|��C\(9N�\�(Qf��N�3w��{*Pw���s��YV]�s�r��ҘQ|�W���˘���>Ƕ��Q1a?HU�������y$eyuO��d���v������[|�����1/��x�hr�K��ێ��r9��Cy���0��b�떔\���7+���"�,��߹���΀U��+�%ù#�H�_����`z�F]X=H�I�³2�r��]]�@ۏ�f��٘��j��LW�,�_�v	�A1[	m ��Z�;��3u��?\���P�pK���^誹�L�tp�>��Y��A�~�-�owU��]��9j��E�cZ6_�ͧ����e:�!�����;ERKH��w�wV��qvߢ/p}���t�m�)3�w��h��p�?t�;bHMA������2�;l��|��I����EQ��u���n�#*y�Y�{����'�ij��l�����
i��4\�ԃQ|&E��!�zT2���]�Hs������\w��������ėi?�0Th��6U��w���Q�r�y❹�����`�Ċ��TZ�qyH�[�>�1�߸�����$J۟�R��B�9ٔ�.2ͯ5��z֡%�R$h�k=W�Kh�������Ț��������$�9� ���{�T�:�$�^� �������k���]��@�GUf���Er���h��g�w���;�������g�U<�wU���+ �^��6��tm0����xA��e����ny�X�g�g� ��2�ּـ�;��B'Pj)J1�6I��� 3�J4�"�8y������~E��k�5��"E�f������h60J��K��PU_��h���W�����mW2zY�������(���;��w�p���L�\�����n����x�HL���𷽾�Kj/�3�8�_���l���b�B��3U�TL�%��I!9�eX��r "��~���2�pTM�b^
�*as�t�C�G���r��94�^��������'�%د9j0ΰ��u��ɓ`d �>��N�>�H��u,��d��89Yo3{�Y)֏\����N�H�g������r(����o��N���R�t�>nn�'R0�HJ��1{��?��u�:�t�Fo�\��v�V�"��_*�snm��Y����/˃��wj�r�&���2����1�ZR\�u��fq���r�
�� c�Ӂ�Ri�o~�ūv��`Yw�1ט�޲+���B��1>V��SJ/�}
��Y�,����U+t���^�*��ݹF�����8J0�0+.x�� �s�ٿ}�e?|T�ܽ��'n6KD��9������s�?{�1��^dy�? �G
(��\��=��;n��ec2�N���Rg	���g��.8�2,~�G{���rvm�����\�X6�+�)-e~�;{�}m!-r�-d���lƭ�!�(X�a�@�&n������fv�.���Þ= 7���S����4d}-Y�ƦDlS�QTV��/W¼�b������U�jy���/�y���K�I�����_�^����k_9{ܒ�z�{�b^�K���Zԇ�u�=ڛj����𱈋��W�������E�7��|��)Z�1L���3����8`�3�*�� ��7�*y�+���پ>�?�X�&�;̼�TW��	�w���z$j��1�6��.e�jO/�t+��Q'ш$dk�z%t�?��R���x�SR��2%�:"�%Z@��!RXr#�Q+�,�ZI�)P��o� ׎L%Z�w]t�y�%D��x����-��HJ��C��m��?o_"V���>�uj7��B�^ρg,��ʌ���,j�����T.��j�O�`OX�,m. )���	t�.�l�ȡ7���NL�|�$�蛢A��o�Y�� �7��P�]�?t����(�Ac��	skЏ�[�K�*�p;2 ���:T�����߾�M�}����+DU.>��:u7�c���$�	۵��E�2�qGϱn��N����hafd�H�]��[�ch���M��{
Z�>�&Aq�1i*1����$gnm�s�-)w�x�ۮ�-7m
�4>��u-�e��'���f,�S�D��a�4���s�
 ������_�l�#dz�I�1�[�z�O�|f���e��~m�}ͯ1oK��D���1������嫻���̋uM�|�&=J���Q�&�@����N�Y��F^���-qx����q���?��4S���?1����a1>�K�u7��""N�ҽP�̍v��LȒ4���2�1	�j�?�|���L.�mh�;��+ [�U�)��%w��{?�1E����f�%�=�x� �v��ҥJT��c ��~����y%���?s���W�󽓪/��H���lӒ�g���G1��G�T���n����'�_�6���h*&�0��&	;���׫�5�؝�e��G�:t?[7P�yA���d����5�f������Y��k����QIxڴ���ahc��b�$�)�� ��/� >�`Ah��z٠�T�m{&��e�A�<W�Eї/�tr+��,j���%i4y����i�IrӰo_2᷇��P��f��=%^ꍛ(���nq�޶�:֚��z���)�`'^��-�zR�7'�(���Z�Q�)-S| �@�uT����]���no���j,�G���3]����{�0�gb�ճ,X�+�p}���O�Jf�04�pl���>���/���<�MQ㸾�tP![ZIH��.���n~Q�B(�48(�_�Yx��XB���=@�5��h���N(��G��[�
J��H#F�F~gRp�)�J�]������!�n&iU���D��
[�����]��"d�A����M}��݅���;� �k��Yhz�$���6P�0��b񫡗l�[�r��>���hu����r�����0܊%��ن���%j�QZ+���.U�^�ƾ�vƔ����3���	%�w���/ c��J�E��X⌎�&��D��X��l
 ����rMp�4�z��0uތF1"F�6�>��{y��������������t�7�+s=�>
(֚�^�v��\��(0]�f�-���tF�R�~�]z���4[���~�������*�$��$mph7u�m���U��w��-�L Q��p���P�Z�Rx!r&��J���{6��)d��M�죞V!*�"� ����T�i�=fv �¾Ȫq ���^�����T��O�x��Z��t!Im�H�����(D=C�|8�W�N��s�#Wh�Kg�������|�?�(� ��:�*]}F�+��m�O"����}$t�><mN4��~��i� /�����q
V.5:���D�Eb���Xh�7�*G` �+d.�٨E�u�T�)PcD��(�7 �Q�Ĵ����8ʦ��1Y�̙h�C�?�P�^��v%Kj��$B��bL��r�4�@�܃�d�m����튶~�W��H�^f٤銓O�A�3{��G��2�k�=m�뜕�x�L͵S���1��P@,��p������c��M��T��/���~fZ8��̊?����/BX�]�,�����3�L<�y� ��V|����^�S��Ł��@A�$�.��m��	딑���r���E�^���2؀̩:�I�Ġ�#ܴ�w>�@���mm1U�Q]�dmW�}���q����0�ud�z�]A��g'�]<F�D����ts�2O[�.�<�~����Ǯ2B�^g9Z�A�9(ŀ4��@o�W@�w��Ց�w����
FpA\e�6�L'o����u�f��R��"��]��Г/>���R�J���rX�la8�r~n��}u�Ź?HWz�txb!>Hyb���wea���*�`�.��Փ8�(�[���ŸBrɲ��^=�%�u�ٍ
�G��<�}�-�Ԧ�N��14@�@'��`s�u���
i�G#�6H�n*5W�J�EY�qk����<t�M��Q}բY5�����c�#��l
��աt ��3?"q��Ͱ����T��ǴN>�U�)�A!ط:"��*��V�LƸ';X#�Q��0�n+�Ϣs�8��H�8�
$�!�I���Ȓpo�.Qi3��Qwʸl\�W�X.>~r��*/�C����䭽Zb~I���s�nl�i�}]r����4c8�'�].���sg�)�Vl�F��3-����T�̿F��:$y���X�;��$M��gO����1u��Tv����
� �iH����S�E�v���W��AD��[�{����W�5Z6���GI�o�@R�k�R����p�W�.5̄0I[��n  `.M��d���HR��h���Te|ϻ:�:����M��qh�<���Y���ǟ�y� w:�0~��<�q��R�����v�쇯�����.�/e�5�@�Zu�D$��F��TV<9��%	q�̞�9��=`���NDv��s#B��{�Z�� J��̠M��J|��E��(��L{!��[��j�t:0���T���U��Y������eG����F5�� �2��'��vV��b���z�AJ�U���-�Z}S���Zň��x|n�$N�D
+�����ʗ�Gպ�h��09���i�?��x%��� ���ւ}-̋��,o,D
3!ߘ�TQ{���Z̿�b!~?r��-&��10�[���S�����]5�o^��6�
m��n��� #�[�!}�f�E�M��C�m��7�Tf�=(K��[�[���/�C�CDp�~n����ug;���>��B &�j���,X����D��OƈB	4Q�(���:���W��r�ڑ:�Pa�������Pa8��>H�$̄x�\��nd/-���=��꓿(΍� ���m\����q�>��������_���0�L`�hd �P6��'b�f��~[Xr���	��
�Ϋ<��g����+1�w/����%�ͻ����9CŅm�S\��v��{s*�H�)�^>��s�{W��=r79c���%����ը�͇�����#������4��C��r{/�Ѝ��E͖�*B�zԾ�⥝z�s8 �M�6�k5����B;ôtc)��̀<�nB:�7��&�>c2{���)��������٠�Θ1��P3`Fw&�,<1�3�o�A�	�(��9#.��T������?�Ј$���4���&���ɤ�� �������cO��s2N����,^�	�61j��h����4��{|���)��7F�I�'=hC�~.�{q���ԗ���=r���m�#�oՖR���}3�� �-�qW
�Vn�$!1[�N�P0�b�~���I��=�t�6Ӓc�Z�Z�c�Ҫil�tn�{�x	��6�����>U���<�P�s(oe����"M�(���_Q ��q�+$��H�7��T@�Dڲ�V��+���)*�::&+[o{���d3Z#!<�SH��Ĺ��|���p��ÏJ2����23A�k5y(Ò���<?�Ӂ5������Fc�ם����:��O:Î ӡ�L��q6���e5]����H�\����Xe=�7�h���.#��
���	yL�� ��*���k��K.LA�[��V��}8��I��j��U�&˜�2P1�2m�H8p�S6r;�C3���j��A��%�iV�����X*�G���/��,�C$q���/.]|���rp��/[�p|:g���轱�&�-g`{M3ҫ��G�C��i�_L��<���,dm��/g��2�u��N��W7`Dm�3��>҅�Ԓ����v_u["�Eг�}rUX�`�D�����!��進��8<�c��.r���O�c���9��l.��d9���H�p��SBY���Ƿj��I�����:5$��>͛��}����M�ǡ�y�L���@)�L�z��
�Y�>�EԼ%�"�YP�?�.�� F��IP����WS�;�4H�P��_��6���m��*
������&�RCF^�w�Fh9�Z�y1}���
�_�^��p�uY#�R�.��4�!��ӈ��WːXm����]6�h���7����?C�MתفԴ��-[\�R����E�3����������[U��G���ypQ�w@hg��qw�$*�JC�3!�|h��vV���v	0�D���;��Z�"-.
���Q{�Q�s���@fX	�������F֓��U����� Ϛ5�V�����A�Px[��u^��`r}?�l�֨�3�M��ݙ����]���Y���S�*-C7��ĖY
��)�
��!k!�&�>�����qI����`��v�h�����}C��$E�0q
�Qm p����������:-����z�58�$��2�ӛFD:��H�
�V�jW�7����B��0����`pd�Ίx1��	jW/��h Z��[5�� �5�^��H�{�ʄ\���-�[��f��m��h[�Hͱ�������_��0��RP\r�c���;���z�7V/�Ni��cJ^<cw}��!
�|4�~Kʆ��[����u������b�I�uz:e�Q1�~�����B��d��/�1��]������tL���\!���$Z��K��ށ��A�Gw���d�?@��.�SH���Ā�j11C��z��eEULN�K���Y�pъvu�|�V�-�e�A�.�>�|�܏k.��'_�6����mb<q�|�96�h��Ef���1�ZM�>�aĄ{+Uk���,I5�Nx�L�E�*t�B�/aCJ�ǄRMI�������_p��iCv#k�
T��������;�����c�xD�j��ـ�Վ������>���kF����a�0���-�p��'�鵬�{W̭v�+��iY��&4�;��c�'j �S}�����B���Vڸ9��H?$D$s7�,�@�x{b%�i�2����oo���n<m�p{>48g��t�L�HM���1�A�#l�N���Xa_s��\$�:�F��������B��ty��7��jo���g]��ʃ�:'�^��w,T�����PY�����2Q���2:*��3	��ܞ덚KN&$-�D���/V���*FuO�a@��E�4]���dL��� eż�<O��D����b�,?\�K��@� ���\��})C=�'*��@�?E�B�Y���m=�\����ǁU,�b�������|����r��#��-E���6�T�ղt�b���ֺV�y�,�?
����뮸��p������`�V��k���&٨�L�B%��*B/�_o�E�J�5��M��Mv�98�@W�cGv2N������9;Gx-�f-@Z�����'�]�b�����ra���m-uG`p%%�h=Ӳj@� ��*�ͻ�?�ڌ����u���ᆆ}���`<]m�ڑ��z��u�>
��_a�{dС_�[+$������#·xD�1���/͍�o�SCf	���ˤ6tl�H>U��C7C��7̍M�r�|�KBW�
ވ8�/��Lm:�T�
~�A��ҥֽ������d(Ďl�{��}��G���N�.^�I<زMV�vF��'��ZWУ,M$k�K���P�"���N�;\$G��m��6n˓�=ֶׁ�pe�GNOG��M������fdO�G'Z�}�Ǭ*]�c	��=����B.[���X��+�4eJr�_�沞%�{��*��i�j�2��"��$=e�s�F�{D*z��P�/m%���4%0B��yv��}�f�Ĵ{T���Z�7�P&�Q/O#Z<�'�<�ϸQ�4�� �p�V@24�{�Wx�⮊	�?�a�:�'�Z�p�{Ģ?{�CA޼Е��z��8
�P?��r�,�^E�׎��Yʉ�GG ���gTF��,�)��q�]b���mUs'x�K���<b]���+�5��t�?�����~�@��[1�V�;��ݤ���p��BQSL{v�{�Ĵ��7�@��K,�F5E��E+Nы�����I #D��~�o�-TS�/9蝰���|'UB�̓�c;_ƊԵ�S�I�G��8e�=:�{H��Qj|͜����k��4,ՠ����M�?vƷ~n������>����g藨^�~��㙜�'`*��]��Z��O��E��Eu�*�S̡�$a'}6���F�/�����N�MΧl�7�h�$ ^M%���+��̒cɄ�[՝h��E ��(�xx��9��I���D�͍o�	n��:�{F�&���e���O�PF"
�!�⑅ˤ�6"Ay��%�E���dE���yK�	Y���o��6��n�D�|O��Ѩi'�_aqϣ�&#.���3��<�������+�{��ri�n�L%�<�@�Hȗ��ܹfË@�66Whh1|ZLŧ���AcE8 hC&�=�w8>���wbׂ���f��S�7��s�>z��3��]lO��f��qn緁keOY�U:�F��X|S��r��
MI]P^Of��m�_�j����Ϲ0�	N���H*0x���[��M���6�*�]�5���NGY���]
ҟ&�����FM������2�	���h��Ag����c�s��8N��J��L��1�0�˂>��_�!(����jY��Qlq�dI�s{��<�^��v��W�Q1WD���w�`��/�E���l�5O/n��h��L0���x���.tg�+w]���2�?���H?�X����\��U�nѭ���/]:2W@p�OC{X���7w����;����X�N�,�a�YN�w���WlEw�/�TU�9m��^�B1Ȕ��'�p"k���b�,��ۖµ6��k�i:Hb�	�ս��)Wh/���+S�C[1�i#�o���J+�=��y�@jhl.Y�ado|+������ Smn�#��o��%�Ó����3�|Xs;]�L�$m�z�,s�h�w��c��책��[�UI1G&���Hf*�0�dI�ߑ%s�:t����� q�W���R�;!��D�n�ۿpW�E4]<�k&�I�Tu1���'x�H���jd�eH��Iv`�
+��������l=q��[w=�X�6�n=�&��F5����ܛ�6�_�����F�l�[*�3 e�C��c��2}u���N�!�_*"�V���=q�G��V���^}��I�a���Ag�Ve�ө��݊L�ͺ��PM9���XPf���X��[���~��X7�}�)�DF�� _�Ж����xsvXG�F/��q2� z �<����3%~bB{ �Y޶fű���8�7��zM�){�3fO�@���[�	��(c���?�Q��?�3c�z:�Ɇ���-f�lb�%\©�j�ޭ��ٔ6�	�?�>���\C��p���wI���]���Sg���/�@�����^s�;���$M3�Cgi�j�����A�Ƭ8�Gȋ,=�
��4Jg��R!ݞ�����2s<d�-�H��C��8��_���|Yꛄ��k�fRX���;!���R��x�����]��F�c
�^��{[�]��o;��ѹչ��`[���X�׬M��:����w����\���kN���'�m�Er�i�na��vP�7�6��Ek1҂*9�L��bG�}Q�[7њ�d�&�����!�1�m����L�����9�EK�2�����($�r�k�}%���<�?�y��e��y_����c�Yp�8��\'!Q����Y�s;��:�=�7�.���k���6�ŸIN����*���K��Pi<�X�~����Cd��:O�|u�5+�B�$���	iB	��o���6 ���c#ڵ����{��6�@�ٽ�8���E�p�G[����sV��;,�]j��rwhL��lG�Z	r<"��&^n�}7�"�&k�x���k!����{�q�Dk��G�� j$ח9��h!�~���nQt�Ҷd!o.h��XI��/�Ů�BZ�?b�,'΀� #����-�l=�n��Am1�	��9���YߴՃ_�	Q�]���\��Jf���*�D�>?�*aa+��7	�ء���Rs�5��1��{����V���C؍�y�m����Gt�X�\ �v(����B	V�0d��z��~����#��`�T�y?���:x>|iU���!��3���$��zGo��ҋĜ+'9!�>�I�a��)��r�c�����tK G&��y�uX�m#�%o��n+��@*XB�"��=��RF�Z�~�F�7�o�?��$MX_������v�@v+"�'�c0mj�Eɰ	���#!�B_(�?�=��G6�]V���Wƶ:T;:W�}\%à 7c��|c����?�	/3[�isE t�~!G�:叭\}c	���H�M�~���Y�Z�0��(RK��X�_��e('�������HY�\�.܉?�������|��F-�[BO���3@|Q�Hq�?d��!Mk��@�1��LNq�<h������%<3`�)=>4���7��	G�G�~=���T��qhLϨՒ[~:���0��
 g��v� p���Y������r�n\" ħ�2J����ho:��'�3��l�̭D��:l�.�#'�O`=M��eЩjn�� 87 !�e��C��Hr��ѳ#��~����[-a^1\=�eZ�,���j<^��YA ������x2���Y��̚�/u�+ �;�P�z��`�Ukj��2���Xّ�_�8�N4-���pk�����(gގB��{��קQM-���ѓ>~x�7W�ns}hg+ŷ�fK�^����n����	���x.K�s(7/8��s�(kW���v9��De��9Ö�ԫt��"_!�c���$镋�%@��G�����B�##`<�Hg��Ǝ�Tr�q_&�]i�r<��4 >���~#��ݭ��Ň6T4/g�0kY���ѳ
¼�?��)@J^�;dׄ����O��]Fz���q4;.#�E^�Z��l���cUs|����S8#mY��op����Ԙf��;���d�qg������ԖC�%�����=���HLV�c|67/�&�Z��ﺇ�[z%߅;��pS�\+h�������c�I�o֓<F��٠S�����B$�Eq�9w��RZi����c�����x���������&H��	̨�މw����hz��t�&�p���bQop|�& c}E��He ?d/�L����ؼSDѕ�/e��,�`�X�1��;�9�l��#ۿm�����ޱ����r#>>_)�ε&�U�'���i��c=V/5��Z����сA
�/��O.0G��"��<@���8�e��:��d�B��ZO���K#�D���i</fM	uRq�6�m���Mݷ;l�;~���M>�R-�YoAyMt�gϐ+q'���mi����M%4����:��'}�$}�A�nQ�Y+�ESw0���Fg$����M��y?��W:��g�p$���["���C�y
���ɏw���T���7ڠc��2�'�r�8u~�G��h�٭B������M^��O^Q�J�ws����P��6c�o؇�"�Y�@�@�>L��s�m��?�2��� _rZ���4U�c
�@3�
�M�'��J!��n7���@��F7q���8s��c��7�t�]��	�e��n{��?V�~
���e���ac4tw�����D�K��լ%� {��Y�H�=J;vʇ�FK��
D|@LҜ�`e�M�3�0i�3�@��A�3o����lxy�6;������i1��gd���.�^(`Inf�xp6&���|�.��h�c�ךlP�!Y��g�$�^>�|TeO��������빪��>���s?��jٙo���g�G6`qd����c�{���&<#��_���d}�����d'Ԥ����J�W�4�j��o�bd�4&}Y���&e!�P錢S�e��&�P����I�}?c�1ы����艟�����7�'���NU��z�>�� ޶CI ���`錞��u�/�`�\�uR�^�������\���cY�b1������ P����ȱ��Om,-����?�tZ�@��b�x���hw�	i�/����=�k��W���Omn�[k�j�����P��T�j4ɖ�ĵyO��C���˅8	đ��&��P.��uĝ��,���L{��O��TL>ő��:SxI�� M��UR%�V������9'p/��΅���E��J!h�����,V�ے*�>�<H	>Մ̷5K�/l&oǈ�!K�X
�q<�g�LE�_���<|F@�J�����փ�g��r�,';��5��۶����K�=M	%{�g�s��`_�P���ɕ��!�:�ꍉ�,B�hŊ�
���> �)a��B�O�.�Z��5rӴuKő"B ���}.=tqK-ir�Ԇ۽��F�l$|���^���U��]߹G�۵d���Zw>�U�!�o#��;�ڜp�q6�.�`����h�,h1�n.ri`�Ұ;15?�r������~
 �7�
�W�go��O��U��x�A�Z�0��r�a�[B��:�O8��8�=� gw��ܠdj$�W�ɳ�-����Vx���_�CT�=�	�\:YW���m+���_���bp�r����PoC�v^��L8�v�\���^�hx%�]+t�g�&�X��|/�mn�q��Dp���|�����M)�F�L,P*�x���X�o�*L�N'�}��7��0�L��࡛�:$H�k���~�j|��c9��8a0`��I8#�&z�z��N#w�I%��Wi@�@�VQ}k�J�>y1"%�P)ʽ�?�1�ȼ��Y���dm�R��e�Aj���6Ǻ��^[C�^��˲��w�.��OZ7��)������|m%ۛ���	|3��0�1��.��ܟL��8�oӃ�.����	)ܨ.���w�Wq�'�X7"g�&t��|��d��W�y�A�	�˧�꼮#h
wo,�w����E����\k ��]}�JZ��+��R�MlZ?d��aU�/�_wѷK͓w�qV ׃5���(!�Z ��0^ѲJ����]�
ǥ%E�L~x�N�GLJE���z�]�ز�  M�I=�}$�����-V�EzUU�~��#��,���`��紝u������tܝ�Z�_�?�^j6��DH��u?Ԗ��C���ydƨ�"��~柕��˖�=���2��Tê5)�����Xεǔ���t��ّ�^���f�N��B���'#�h��;꒏v�?�}�Ř���=Ko(�g��A,���i�E��L�K�����7Ft`>�?���������~����6\9�ԧk������,�Q�q����5p���u�R������]	~����L>��KoW�����&L=`��_[��+`	�A�R�ks/_X�7��O�r��q(8����v�ĩ*|\$d	S�] ������a^��ڧҋ���]���:��Q�i���4��~��5��n�32�?�k����c��Vnֱ��׳v������
��-⨊��c�!�:���o��r��o|��:U��6���uՅ�ACw�����+�l$���>�xQ�){ $�����3;�m^�����rD[�^o`t�s{��d<b��=�:�s&�1���o�L�j��*՗�V��.h�E���W`�$��G��.�I;:ާ&�r��;r�����3E5shpe/�ս�0�\,ˌ���Q�[HiN7��OZR�n��h}t����^5]��ƪ��PsQR�`�stȷk"�{R�!`�6�����]�u�������\N��7�r�ď=�����@
�v^%�d���ƪb6o+�EH߃>7q{�]�?*�L�*�BKZ��Sb���L�W������0��'=?;jR��0�7����}K������\S$ǥ}Lx��%�f�.�E���}Ѣ������X���a�So���rd�k���/I`�)�oG��L���਩�U�!N��P���G�3S�O
�ȃ=˦)�Vw2}})��U��W_�+�龤M�����+�"x�7�$]�$��C�����:e�Z�e}*Z����ӦF��c�;`U�P���cu�0;X�#�=_3_�WA��;%� ^7�˯��QR��`����nF]o�N\���'y�AL�����$�"��c���b��!��GX����*�� f9	�[�$�Z��HrO��U6qP�-N��>�eWj�a��Ez(�P�53{K�(��E�L����f�}���	����������.�qu������N��"N;*���eql  a��\/�r0ti5�f��~�+0��yv��s����B���&����Q��"2MC_#����#���N�T�p�e�C;Ƕ+�h�&�?t�a�\�����8Eݸ�7��
F��y����"9�X@�c��G7	� ��gwPЮR=�݆w+��>����0/�ǘ��<�����+�>���2!2����g����'�Z�s����/�� B]d/���k�?�s���'�4:^���ݼ�I�U6���	��R|�cdW,#/̨oTh���K�x�ud��Ջjeഒ�B�y�N	��:����s�6�`v>e�A���,���Ә]�!�7LF�Ե8s�A���0�f<BԎ��,`��MG����_���`�#H�k�1�!�zS�?'q���s�`�9�y�rIb�E-�j��{%����{��]���be��:%�>�~\ZC�3}D~6�m��ˬ #U=X�zG��=�8�J�Ty���Ň�Z]�S�B���T�$$�y� �Ñ������GN`E��3������v�CB���#���������T�0����0��"s]��� �o!p<�4�>Ou������AɿS:i:�G����*�W�V��r?�A�H~\�S���D'���x����"js+�j�'!�{1(��Q�*���ٷ�ު-�4�Ŏ�)�Z�� {�b0Mh�J̺�
��Z�]�@��Ȑ� �������G���&�4yU�H����=�8y�%�k��y*�M3C}@~��`�>������y这�`��Ϝ�d,lh�R��s��\��(��5�kE�X'�� "�fV�B~�>d��U��?f}7����}4r�y�[`�~��m�����QcIj�ۥ�:�[�M;AZ�|���l��
��Ai�����~�(�s��^δF�W�1S`r��ՂgmP���:�p�^綫����lt��\�`�e3*�</� 87��o�n�DI��N*�e�;F(ވ�%=J]U�\$�F��C���ũ���L����x�a�PC�'9�9�V���5��3�Κ�,��n�X�搒���j����]��)�,��ZL{<+��}�0I��VSn�@��~�ەL��q��;ƟH)R����5:�y�}�ʸ�.��%�۞J�v��Yz ��r�Piw��W|+j���}���	���_er�Lѐզ�f	nO��&X��a'�P�鸣����k�AR�*ϵu0ԙ����+s��	�`�pX�1s��<y���8�Ӣ�Û���P�H���6,
����?�?�����>���,<
�%���$#�g�':�H��KQL����������P�"e�}̀[��p�`�<
�%g�)ߗ6m�|ֱV9>�t^�Ʒrg��eU_[Ik��"sv�X��-�<�)�l�f�/��:a�J�{@�(����ٹS Ch9���%��r��~M�������ԙ�{��O�N�;�>�wwϱ@��# &�WQ�%�]8������9��N����u� �Bk�]Ouq��
K_�O"2=C��@��k���zA��Cx�l�{� �I?(4j�����%(a�����E���`'���az��̢���At�|��~&>�l�vǑ�
�{ �q�?�7�-7Ur�C��sASn�Sc0�K�R���Z��̒W���z��zy��7U\�6�~_�9�����XM��1_�#z�͝��q�m�@a�~H�w~�0v��t۫�=ʧb���S����O�^.�>v�O���<ѷE��#;h�t�5���!<�ۜ	"?��e�ml�͜��؜~$jQʇ4���.�8a�v帨�h=���gO/!r�IU~\r��$z�q1�E�Q���/�.K��@�[W/�H!u9AG�j^�ϟ���:\O�M�Һ� �,�dg_ZH+ƚ����P�]� ��""�nզl��!g�j���-m<
Z�y�`�-D���[�o ��aƌ��嘆↓�t� CN��+���?��*��"�5���M�:ؘ�J�EI���3�+i|
tx� G���V5�&��":��_5�y�t!�ջ/��H;ꕼ=��s&��C�V��h��{�F�Gدa�F)�X��Z�=c���v�Xe�٠��k�\a�����ū����R��Wr�����3�/�g&��Ĕ4�.��i~�E���]/��G/���6�"��P[Y�(����!�EQ�˜�$�~N
�sB���/֪#�oa����$�f8�z_Z4t��P��#H�*F���M���l�%w��.�ݐ�}��	�����Gd	��m�����q���F���� ��� ���9�Gg�jy���6�'��I��yb�"Z�z���=����om�I�$e@ܦ�Ch��˧��Fp>�s[��Fa0��ԋ8�������AQ<��"�$�Yњܸ�eVv�?ǟ��݃XV�Px)$�8D����nQ�Vߡ�@�pN�9��d��ۖ~�is�;���Q���jRr����jԒ�ךV���|*F~q�٨��s�D'1��x98Y���S1�5$�(Q_q��9M�s�l[�#}���0����TZ_6�+sH�Ă|�L�i	�k;>�3�S��p�!�s����s(��b�q��(RA��Ǎ	D�xxo20�t�����A��.��5p����K{�V6IX�����Յɋ<�[TF�q�BÅ1�h�}��u�`u<�`���3��[�V�`3�?�^R����EJ�ڠZ�"��������w{�}�%Fs��m���+^��k)$���"`4dit�c�=^���\l~[^@�-�U5�g�(b��у�YB��l����P�
�[�A>��`!7>������"'��>�"�M|A��^e��J�;�T:k]0��"�k@c�6�(���T�f�p� �qZvA��-��I���m@�;j�ol7A͖�s�z�~1�4�Q-YB�i�EK�`����+��כ�����DO���>r����Z�iFXS}�[�����]�<? N��?�+�F���.������cW9�
� cǺ(��LK�(��@G
2�F����5�����6rY�P;�̭��UW�(|����
��|-J#�U��2����Gpw��湎��tɪ��->�H��aӮxZ>�]�)�0���Ok����,E�N�C�t-�y�a��i1@۞ј���	PU3.��0���B�'�P�v� (K
�$2�6H�G�ӆ��A���wi�/��G������*� ��XlE��y_�
�D&-�&�j��2xqw�$/<4m,�2W��(���G!5�M�@��r��Z�R�b���]�5EK۬s��:q�U	G�(�o�9ϝ"^� [x9��@���So�C𦥷H�v�nT�6��Q��b���X�31�2�.�3�7�eeQ�R�呄̧��{y����Z�Ɓa�P;�E���D�q9�z<-�����WFg�v�;jѥY�[���(�kC�D��%���܎{��T��A�q��
^��q�L����:���[�B�5.z?$]a}6,�<P
�WbٍFew���_��}��U��!�#�O50��t�PS+E���3[ ��c&RR����0Wk���v@U]
����8H�(�
�4��U�5:x{�?�_��Z�X���Uz<���U���5��@r����C��㋮oK\�p�}�oD�T��z�kL#�����!�y݃����V��E��>�����F��@V(K�Ք��Q��+^��� ����ە�	������K@����;	��Ao���A\�f��>�޴�ت���C@�@��~)��;�?�QE��T� !������
�T�Vi�����Ah=��Xx����N�Sf��_
������~�n��{���v�LZ��>[���{L-me��ɞ�c?�*�,h=�)�f�.�k� ���MtaB������x���s��Q�21!�A���Xk}�rVk�y,�L)���d?7a��t��AM�&G��72���A2�
���u|���NE�����+�P�dDn����u�\J}{�����rP�g�ţ�E�6"Q���F �ʊCM��3��T���lxq3��ot�d�(�:�7��'�7)�����@u��O$)��%^����3���I�7����m�Dvm
>D�Boļ�E���S��K��nn��8����IUi4�(u��B�	�"&��)��"a6ܹ�Z����s�y�?����Ld#�U������L�HM˧1�q�°*K�on����桺@����w銊��%�3��Ć12��_7D��S�F��]*u?F�P0º&O���?+�@4U8j>�0ƽ�](�f\ԓn��"JnġP�C�Ϯ��n����`�n����l�G�y���_X^@�`�+�@���(�j�lg4x�iqď���g4k�)���6����۳��Q#�hj.lw�A�w�=9*���t����e�L}S����¶�#�%���R%�>ކ@ ���ѡ
�����'d���Pf5:��-q��l���a`G�����J��>�g�F2kIv�Ol�w�Zdˎ֣��aõ+k���o���.�լw���f�8�O50o��M�?�d�wNa�2��6���4�T_�����OUѵ��	u$��L��>�P�h�W��/#�*��텠Tf՗/q���z(7kۅ�F���]�����җCb�!�͙z[e^���%6]N:I��K�@�� D�ӵ�D^��횚�'y�,0(u��Ь(ِ	,�a��^ѓQd��d�!���Z�āͪ�E�mEɄZ�o���[�~1^F�f9��7ј���I=��ĸ������=.��c�q�9}�b7��(e�h^+ɘV-��*<ݣ��y��n��9vm@!d��x�kʟ�b�����h�-C6��8Hk/Jނ_�;h^��X�O����PNv�i���j	A?�����?�W0���T�x�\"�Yl����b�k(v�f���� m~	Jv=_�j��^[��C#��N���ɘ~�g��,���͞'��~��m���DN��AX�ks~��b 
���7�)��S���?�y��qZ��;���D}q�`K�"�/��j+�j6��΍��,������E\�_+B�7�I�#�aDb"-����oy�&Sݷ�r4
�g��}!augI��Qڟ�a����#�&Z`��k�>4��mT�p:Xǻ�&�5��x�c\u�lw:1Y��w�IDZ�-x%2W�$��\��	/Vc~�)��:�^�e5&����! v���Z�,�!�ETZ�Ll:l�H�Q�:i��i�T��!]I8`nuv}��)��q���S2KQ���i���/"��5>��s��5P�Lx 0�ԓ?u'�8\�&e��[+��H��c�>̇�=�S�@�/���"���6��ǋ��g�?����c��t��D�ύ`Y������p���w���q�x�ǵf��7K67ɧ�a��d��-��ל��8@�e����:N4�����6LlE�W�e��3�.��b�<ZHḄ��b#�EZ�c����e�����b�l��j;RBx'Nn6���¨1ҷ�ؠ��!��r��w��ږ�FI�li�-�A�FA�E�cx���|�S��|�7����z�>fd0��DO��!ңf��n�pٌ�Q�w�+��E���i፷J�UQ]�_���e�Ѐ��!?�#1�6����u�[�\�&6c��.�ҹ�W��Ԑ�?�y�?S+�WxP@�	c{6qiVTߟ6|-�K�ҡ^M@HEtHv�⤬�bG
��=v@O���G�4C׊K�	�,r�0��f�77�g���W�bF��8�����o"51K�4ku�x�Z�ظ�m�G����0ߺؾ�7UY3y2_/�V=-ES�Fq%)$]o
����0��dۢ�L{�QiJYe�"uY�S*f��׏n��KQ���H����5~�4�i�KL� l;Sq@���y�̞�R79�I�0�z�w�;퍵b4����a&�tM&1�w>T�Ն���'���Z�m�M釩Z�5S��R��ɨ����^�E�\�&e����;9��
ϊ��R/#��ֈ��$�X�I��g2I~���u_n�+���5��M��54��^�� �.��=;沼��8v��&,�y�l�"�˫"eE�;x/{�Fy�t������A ��� �q�����:��^` )�PY���6�5U��Fi�0����+������	�����O�-f��L^ً>�R�Շ�:5���-�}��j��𬙮j�<�Ri��h/2?Cd�=}RJ�[UG�5$�r�w(%)� \�]�����W ȞD�;�xք<�'��E��4x�D47g��;��Id�B�o����6�:e���jHf:�e���]��\����vi�����Amƨ�l�2F�2`-BB�����*����	�a.�$���1�F��k�2rs�4��Kv��
8�atVm��`�,3V7��h�XwK��מ���Cdw�z#�\*�(�sj�8E���#S$����3�[~Ѧ�8�;Slu�:� �z�s���Kܹ��U�� R�����I��7��U�8]4y3��{����~U%"��	ZcT��DY�R���@�ݨI�����_�V�ٞC2����p�g<0����\0�P���(����,,w��d�G�6�4�U�T�iG}7��8c�<�m:�X"	�a�WS2� \�65����Ѕ�u�!�����^��6 �ĝdhW5�������v��T�B��k�r��	U'��?3����z�A#ح����=�2l��s��	b���S��d���gR-�*v�N��/XȌ4��5�Gi%�=g�x��� 5�����LN7;}�����wKz�"���kk��C� �}�U^�Zg��f��k[㱴QX	Ƴ09o��ϝ�c9��\�'��T�mՏ`�X*n)�{6�~�g)U��h2��lm7h�u/�-��]!	c4�d�B.h�[��Գ����(/��C��h��ߤ����P�@@�.苾�^�
���/$��h���;^2��u�#p��&	'������kK�X�f�W52|{ݱ���������^�y�WZ�ɣ�����X����@@�tZλ|�m�n�E�l���E�tMDO���J1��L��O��|�� mu�'!��G�^��8��7n���[���-(k�/cD��:�/эNm�Ρ��C�|�j��Oⷠ����ˈA���E��v�{//H��b%5=����t��{�.�v�:k�7�2Py�|�`��j�l��z��C?�՛�~V��7Ă�X|<���$��"�����7�Ĭ��
4! 1�X7�b�SM��	$5�u
;�Pr3`( T3�q�b	�osD��&�@͜�P�����O�	f��QA���Z`(9/gF��f��9 .����bW�!{������|��R�L�נMB8j���2;�F��\$p���
���3���u�Rn��r�z~J�^H��)�)��犵��~+���+Aު�&l���1�@�~�'�P�|N��'�{ȫ�R�v�Vd�Pw��V���?��$�A��V��Ep��_�)d-���O�է'g��Xܣ1˾),��љ�f�k�?�y�!O3O�4H���Px��K��É>)C4X['�r{icQ�BL��` O��	�C��#\�S�s���t��Պ}~:i����M��ȩ8���I��M�](k5�9ѰTH����t��6��+|	_h��>�*�3��Ղo�p�~}�K��l6(��W�������{��@(,��� B那�A�/ ���6`����4A�^��?g��ɏ��[��A0s|�g������;!�S�B�pm�p��Lѷ\��XT��1�as
�53�����l�r7U��CVR�⥂ƕ0g�o;�Q����guf�w7��h�w% ᖸ}�ǎ�kA�z)o��R��ߣ�$��gh'��?�䠸�?p�
~�Gg���وE���,�6%Iˠ��c~[��TG�/���j�@�����UF4E�蘦G�t��1U��잣����^qؓ��cE��-A3"8�@��3����S7�o�j��v��J�� ��Lo�H�r� �W�Wt9Ɏ\��1F,���MA�v8E���
�J�%�ÐTGU��ue����d���w�Ѡ�@h����������:9#�9t���k�c��4�H�y*�C�<3%��'9�B����Yб����v�]��8�^Ni����8�ib��ܴ���������&!+|%M�t��A�V��|�.��}z�j�μq-�H��=_R�ŗ��}���,#>��d�^EG�փ�0I��Gv�t{�紴��뚴�k&k���������l�#l���9<ϱ��"2�OEe}~a��K� ��q4�	u����To��˿�?�"Jq�1bO�ܱj��ߺZ@d\!���w�,�#����@<�s �����\F��3�n���q��9�lhc՗�T�5(�u3����h�#��U������c�n$�ߊ������`�2G�We�, י�>1}9�x�O�p��);h��,|.��y��[m���$o�D�0��}&�9��yHK��IO?��ѵ�?��:�|{�#z�>���۷�:8 �z�%&�4`L�/7nr���@*'=���1(�[�.�Kl9\��4^PD��b�lx4HR<�KQ�S�X��d��]ep�D�khy��7V
Md���	T��]���z��&#y���#t7��zZ�t5���ѡl�o̭���bO}��q�O� �6"�n$p���#Vb� �,2L�����(��'�Y6� V��΋ @��Ȯ�!RrTr�Yz^�g�aZ3���K��J~�q�l�I]E�Ds��h�u���ѣ]<��v� �pP]�ٰ߲�(���;���K5�-�ׯ�L��9Q���ׅ� FC�N{pI2��<��^���t,,��,��ȹß �� ׃�⌣g� ��O�d��=�:��a�|��r�y�|�y�/%L��*�y[�!͟m׾t�0���E\$DBS_U�|�~o71�����^��H�C�����[E`P=��$ �p[Z�d�f<�p'J�1�S��5�4��\r��VV~N�a��^�s j����q�pK0�fU���GK9 T*tP�(o*�����eP��u+�y����u������q�4�\�v88♔<���C�nf[�hǕ��^{���tutM˄M7J1J��W��L:�̶S	A��l��,�a���j�B>�(��{��*'_���K�%@gg�=�t� �6� �3?�>efF,��6j�[	y8x�����it�chr<˲<>����X�[9�F��̺���[�j���Ӏ��r��A�b���ᤥ�KO�=�ՙc�|����Eԑ9(:�@�Jm��\�.PH�6�2e����e��7H��A����h�9�?�d~����w�q]�VW�fd��ng+IO�\�O�}����m���,�v?���Î*s��XSg	p�W	"󣧶E���e�K��z'��g���TR��\M"���dI��]��(�"@+�9�����tM�.Lpqb7.C�K�v��	,Bš v�ʌ`�c閕��%��3>���O������7��H4Y���K�#�[�y���'Y�ی�fj�3uw����գ�f0�i
��t��SV�Y�cD�7�,�	pfv;����Gz�>Nd^�!�R�wc�)�^�J�Y�޳�z1c���g�{r�oH��犒)���r�m�d1n䱊ݝ��ug�����=���[ڰo�.ڗt�d 0�xg���[mT�Q���F,�P��'-������ �*�A V�4)Ws���7lT8��Й���;���Z�)� 7Ԑ����?�
����C����x�\Mi�(ɞ@ћ�m$z��G/kk�hH(� �cVJGs}���n_~�z��nC]E+(V��L�
@�%`���h���_����x9��a2�9N���Q3�_����ueq�D���k�r���^V�Ǻ�Q��},=�r0�f�������8m)���!��<E<M8��*$��"�WU� <т�\�,�-ٮ�!V9�(Aq��gq|�B���0���R�l�ņ��!�3$�'� ��51رF��{��;�~c����>��tX��V�-3`SX�H��v��cF#��A%�����8�M�$��D��ON����Puܸ���z���HS�/�s��2�Dg��P���jVfc�J���_TZ�y<D��9'�0�b����LB��l���M�ᗒ��D6k�_�˷ �-�����E��C�����#�x5	Ӳ���Q���$%�z1�)-<�A9��cB�k�=��1�M/�Q���ur:k>��:���<V����:E�ڲfȾ(�N�om%�>��K�ĝ��X�)~�'� v���@Z�/g[u�$�g-iJ�3�E�2�#Vl]8����|};�Vl͝e�{T���ހ��@bKJo��͸��0p�Թ�� ��S�c�����>�ﷸ�\oj��Ѭ#�a�����l�K#R�u�c�[�:�����HC�X�׸���E}VK�l�\�B�� /f���x�i��]��N���M���H�w�*y}*�,>�Ҋ6.�Y{\Wu,�1��fD�y$��;ڐ��JH�y�:��Mr|vj"�gi���	��@�q�a�8�MX�3-�C�o�!�+?�F��J��B�jlb!���#�K;v#�{�
�Y����K/��ŏ�;#l�����c�x��,�y,��4`�5Q�Z��y�(���%fFQ?a�����!��+��a�U�k���_�B��#o=��Y7�k����kPP��r�����<ܛ��NVP].���/-ϻ?�<C=,sw�͟�v-(Mӹ�*�������H����{܈+�6�>��c����{"��Q���?I��+�7���P욞Z��y���=G��},2����Ct�|��}+f=�e�E.B�(��v�����C,T�L�SN����{Qn�����P#(  ��J�Cy�G��"n�lT?�嫓J�9���#����6$��o���雭Ē��5��2���/�K��[��i�@&0�Yܧ"�w�Z�z3���G`�fRV�Pj��AC���*Δ��X���E,;-�*�v^����T�J�3B���M����^o���Ֆ#!C�1����I�a�p��a�����1���>�3~=�xF-���O4C�w,X$3��k�*/j�n� �-)8h� ��(OD�[)q�p�R"g�������fx���g6�W���gcԯ��!˱^SA�e�Z�����`��8m��OL�"���8�U���f-��贫�18�L�B���)(��i �f�K��Bt���g�`(��˭낑겁[�_�q���?���Ud59���23����1��Et�OP����Zn+44����#Alo�@R�9LB��/��,6@\�{������%�͟�u�o���4�W�o^��-�M[�vj?)���3�ܿE��t�GƇ�F��=ƣ�.e�<S�%���a=�\)�(礁W9�qo��ܹʀU��4���r��Z�.n�'E��rJ%��[��ZdZ�+j7g9����@��( `��i�6m��Ϯl��οi}�_o�ְ�R����<��w�� ����$:P��h=Z�w�T^#V�Ow#��'W3]��� Œ<������G�D�b6��M�;|u��c��J���2EE`ye\UW��J�$OF�}��g���s\!� ��|�c�T�wT-b�S��&�wU8�X;�s�O%�74pp��m��bSܪ�1��� ��ꘇ���^�&����g����X+S� ��kt��s,W@��N��>�P	$��>f)�Է�'0�T����V�1A���Iz��I��nk�(���#�t-*C?l�g^�i�i�GC-��Z��˫>�/O��i���uT�	=�<����*�xfo��AnM�G�%#XWTی�.�\Ի�������̳;�Typ���5����-��SA��#oDF����ou�vޖ��$9�.؇�����������,��7���;{����Ӧ�0U�����樗T�c�ۣ�����Y�'�]��ٻ�]�Bm�Ne���ɟ��co�l��Jϡ�3�d���0\�GUr�.�-�8wsI��uЁ3�+��x���[�n��g资����E&��ِ�Ѻ���R?������t��[����5pԕ;�b{vY���}��ZF�X���~@]��M[��q���R�A�Li؜ćM�5w��UX8u[B,�IJ�Ã�{L̾$[q�|U	�2Q��
*&�\�n�v܁�k�E;y�r��X2�����<�A<0mW�`&��2�:Oo(q����oN���?�D\sp��4��vӁ��A������OW�ag3�e��
�m�"�pez������$��C��Ӕ^Iq�!?�q1�ʋy^���y�E.,�����`Fm�s�\�y��(�&��W�����v"�nOb��e��̍6���	�3gXm��T���|u?f6K�j�C�~B�7�d,H'o�Gӗw8q�DpH�7�:�\��V"�Đi���-D+��U�j����kQ�,���$k�(�L����|N��@��%r��؍?�O��`bVq�&&�;GH��WF�\D:^��������rS	�/o�)�A���w�#z�&���@^p�g�������>���� G�&w�=;�A*�WmhO�oU2���&�����4���}#u}31jlkp`M5X��\�p�zP�S��7�#J�m�#������uyu�N�U�1��Y)j�.qp��0aIqm��R{�F&��ꅖBt�e� ���i G�9�οq$G�ĆX�����/��4�24*l?���Gs�����qz�)���&�����h�<����K�DV����.��/�Z��t�;�f+����j���5��J 4<�b7�D�����N�XV����c�P�l9t(�E���q�<lS�g�
Pg6���AvΠ�xU0�H�~��V��}Q��j����{2����iBO̼�k(o6ܹgI���8kK��܆���u5��JIn�6��I����	�=�*�kO��!��yS�3���A<Bbiss M������e�u\��D�K�>CI�i�׹KA� �jAp"y�.g�E��E	6w��z򤮽��t�_XO�W��,��oM��H���=�tZ?������8�ǉb��(kmgfu3�/�v󋔥�������Ň��F>?{��Ur���R��ďB��]}�d�]�n��}�c\�4�@���O������P��Σ�59����*<�fUւ��=�(�.�O��ݣl�ϡ	4����0�x��/�1v,B�oAD�E�]c��Wk�yk�_��G��,��#ǹ�ߠ�%8Cz����d��?9n������E���'T��j��4��]�$O��K�藳!| /���G�S	a�tx�[Үt���k.�ɯ�X�&�5_Z�'UPi�5���`�a�d0��%��:�����0�/�h<���,�I�[�xpB:�0���;�I9�6�1J�
��bK�������@��x��+�:P@)���Џ-8����d�Oo�����b�6�&�������-�уh��6�ح�.r3���y}S�(�i���=�Z-^���A�?�'�).�?�Ƹ)-,kzT�+ZV4�aqY0�f�p�"j����"��:�[J�,�La䠕ʄ�R�tzE�Wa���X�'/�%��8�=�������Вc���_?�n-C	��t�����ҁ�=���E�C
���<����RH%�ܳ:��� C�p���޳A���,����C��ͳ��6P�':v�F�����{iٷ�6&��6���5I�6�K֢�L�-�{���QHW�����Z�t���'Y�O�2�y�J����FP@�+�oe\�]��$�iX�w���@F��,���A��3G#o�f+0c����5��h�����t#x�푁e'���<T�tV�h�Bf@
# *�ԣ��&�X+�d�"��S)b#�4���9z��cSs�l��W�M�|Z��<R��
�"r,)�~����#�I�����-�Nw�'E��yz�m�~�U��g]q@����T+�ӃZ�F��|�n�M�H á�	Gy&,�\@�V)�^�~�$G�+����@�0S��ΛPc�` ��u<�/$F��3�6�pO6��x�P�0&���{�v�G�t�����saY��y�v�9�!�~��i��S� �����;��Մ�(_�H�y�Z��v7>2��U������'��"�.�Xl�bU/.�sg�h�*�<IxM�	l(�u��M�612A��^�Y�/2A�p�ow��e��>Ԏ�����WfB��^lm҃��
�~\{����qL�8��î��� }%�!1����vn�eW�{\��Mz�9���S&�!#sP�PX�hX�>��c����L��ŏ)��}��g~+� �+B�+�6�Ō�6���o%���x)�I;�y�p�D��R4�5v��Q��A��
�ˊ�5{��$�'���5dWuo
����r���2��S��0\�!��N�ss����9�ȣ'SF/�V�	�lz�Υ��?�w�	KM��f���m��'$[D�$D)�����h$Nt�}��r��!�Q:\�3j�Π�̋F���f_��"}}�.�~����ٚ�d��E9�츌�Nn�� �)A+��쏆]�}K̥X���Ό�q�p%DF����NWP�>G�h� [��/�{���~>,��Dӏ���֚ɴQ~��>��E dc�S�{w �V��ة���������/����̗~�u=��!��: ��f�n�Aͺ�ɧ�k�\�[�F�;'{�E<��NG�08�n(��/9��r��8���y�i�77%�W�S�&�z�����ѣI����ș��g��J׃�H�i�`�]���QK�_��(���|��{�����h6KY�~In&�z�?�{�Á��:ĸ�������>�$�d� {P���7�������6��^��؀ڲP�o�W�Q�"Z��������<ewӬ�$���jWG�73p��{��L$�o`�����ѯ�y� �c�*�*���l�"��r?D֬���$K���Ѥ�[ÆA)ګžr�Չה�:=����K�n3�n��s�Z��'F��� �ˆ��eI<�ę� ˖�Hit���SM��.�Qi( �Zx�@�,��=��YMUE��=Q���3�j����O�H%΢����4�*��$�rpK��?�./pCý@9ڴ]������"�����8>D̘�;T���Qڔ+	���;
��g��o�P֎���;c��D�_�J�-@�`�/u���>��������Lճu��0`P	.}�Co���yL�"��;n:�_�,S�/�B���C���K8S� �������E��b�λ0`����b����mA8��	�`+��?�P�u\�)i?K~�;�j���!�f�V�g� ���a�gʃ�9)�����&���<�A���_�L�i�޻��e�b�d��F���Q���=��I$ц���� =P�!�be��1��G�A��y�d�jUW�]�D,�'W���RI�6	=� ٟ[
)aۋ�t#�?���(�m�,��r�cM��\�Jmv������Q����L�L��,}��������Jp-��G��j��u�jqi"Q0X:t�Rx�(X��C��N/ԑB���U�Yu��"Jݗ���6�T������7�W��\�A=&̹�޴p�W�JtE�:��Vv<4��`i9�Un��k�\q�~IG�&�\�����+M�O��G>��B5m�hH~K�(ͅ���Y��Qe����|�r��K��7����j�f��0���h�K2�j��g)r�����������u�"ds��٤/z��I�<���.�o��bH�/�|8��V�+����������Q	?\�	
y٦N�q>v39	��~>J���;ݳ�;���se}%��uL�'׉� u��;}�-rTY�y3P�H����@�}I�_H��C��\1�$�p&�\k.����j<�k+rM��̧�q��}���E��8��8��n�����K�Y���b���L�8u�7ϋ���߶����e�H��BQ���xF�Y�	�����1ߒhZ6m?RAU~���\%��?5:!h�:��0N<`P�ʏ+3u���]P������YF;��4�u�7G �CQi0����7~ǌ 4Y_ᨙOY_�Ȳ*- �e,�H(a�{;_ۋ/���Ih�J�
"G͕3ٳ`������~f�\�_���.B��7s�)<��so-)ܫ�,%X2V�
@cI�����:Ik���y�1:��nC�����i�Ek���7kY:�
6�a3�י.ugc�6i fc�W��,�+�����w'{�������LO��izZs��NakU:�>i�
�>���Ŝ��G(ᆼ�k��r�;�8�*�Ȍt)2#�>=5��5u�����g���ХV��7[MŇe���ꬺ��ۨ��J��c�3@��� L���G�������|�R��:�,aBT0�e��%B�ד�_=�T
����p�{�(2Z5n�иhG+�]e!��H�y)<����1a��E�������$�d�����4щ�5!��gb����#A%_�>k�3�X궲&�)H4���* *�u����4kΘ���hV/�({	]���yt����`��*HIJ���+w�V"|�����`.}f{.�C�"=�ѫk���:(�*e^�̌�\+�"\q�f���(X�I�A��$;\��^gßq`��09���k,6������L�c(\��C�Պ8���c._`�W#��}p�T��ӾNe�E����x��2�[�]>%B�+��F�֏*�l`��2sR��5���m�a�0���_դz�L_���!8Y�;:ni]�B��>�^������>���ӾQ �Y�6�)��S�S`)���p�-�Ȱ�,��yc.��1��-7���zhidQC��m��3���M�� I{'R �j��b ç�X�É#Do%���?)��Br� �l��7�z��npB9����]�yb䌝�q!�����$���E���	U��2�D�Ƕ,T�^T#Q���:�*�+�5�Y2ҭ�G\E/��$��G/|g��c7�v�d���l�3��`	�{�=P�E�~B63Nk�@_��̎��|���D�p`f��rށ�Ol,�h��*�/f��0�8�V��jР8*/�WˇW`�qL��/p��}��D�ݻ�%8�}��ͺ>&jݻt�&��|��R�EL�j�Qje�C2�6A���x���ń�X6a^l*P ��U��-=6�q!L�.�@�Q��@" tG�e&Mӱ�!O��&��굾v̊�a��C�U92��jJ�(9��Λ��<�	�7�����P���i�Iڢ��7ˉ��&c�K6YFT>�A��9��H�@�+*r��Ldh�3]%� -1s�N��nHC�-��D-���ĭɱz�іt�`h���_�A���t�������)�'�L^�k�ff=V��u��~-���w)�4�H���W�4����	��Tا���Y��P0썄�y�ޭw�7s����ꅷ�P�:�S�j���>N�04CE���ě�y�kr�_���ڳYWG1���
0���S����SI.�J�dV��f��6���?�(3�}��]:��A��m
U�'��o'���m��6l5~��%��B���I��<�n���q���������CA�;����s�*�͑9����#�~`II6"4�2��>�{yL��U����8h�M�D�*Dov�������j�ю�������,mgD[�m���Y�=O�)p����0�f^o��W}V�(�����!M�~��.$��G+*��'n��$}adʸ�4����d���M��eU��Y6-��{�r	}<���pkJ��r�~2���&�����h¨3V�z��b�U��%�ٵZ�4Nv�T̈́_�f&���b�i�y��x��A�ߢ��kU5)�YP@�;�Ǽ���`�Hp��e_4�+�YnJ/�}N�u�δ`LJ$JK�m���;ˤB�rZ=+,���Չ���cqe��p��G�u���������j0�ǚ��O.�`t�3n�#XmD:D�p����k�0�5� x�j{�W[��$�9�v�/�p�>�n��uñ0dtA����ps�ZK�9n�\#2�O�U�� EI��Y�`��W�j�Q̮<DCqd�	ϻ�Pn�	m�FT7(���^���?�2E�YW<ka��&�Q��Ȏ7�#7Fp�]��cΉE��7eZJ�<��r%�&�?7�j&��K���<�DչD����i�d"X�Fs��B�y��_;���48��D�đ��D�ܦ)����0��H�i>H����o���F����M	6���#�K� �a��'���܆�G��V=�[����+�E��oϮo;���ɚ�JCB�����:�5:#�oin	����y@�����u)���}���`�^�y�vl�g��L�Q�-���z�O�сnV("@a	���P�-��6�Hr@����ץ��Q���@�_cǔ���X��f�wJ�k��	ͭ ��.�K�Q\c$���E���@	Q�n�d�%�hو��-O���B���y�:��{��H�ȳ��U�Ǔ��_s�9����6�dY�9��:�D=��u����+m��������BNb���g��,�b�Ϫr��;5��+'��8�h�Z/�>S��O�[S�[[����pr�ܘ�?oi^�)����8Yןڵ�}����g����RvM)��T��������eAͶ��f^:=I�F�x͠Qr(�5ߓ��v?���͊|Z��=H��^�D(Jk2L�u����~}G������"�t�˵�KڏF�������Nr6sܢ�b��-˺�#45�5E�:RZx�*�=>�h�y��B���8�٥;tG~W��e�2�|�b�B6 |��G�9�tQ�z!�G�4���B�>Z٣����]-���%�
N/Fg ����d�k:�H��,-���R/����/FY��9��Y�����!�C�	��ԛ��i^uR/�I1�F?�p��1�h�U��m]�x��}�8 }�S������b9GB�v����b�2T��F�=�@�q�@�r�~o%Ԫ�z�UxV�y#|Կ�Vx�ᶩ�< Ĭ��e�{���x�]ޛ��3O��满�05p�#Y�-�(4?-��Q�Vb�a��GD�>�G�A��Gi��l�G`���>ުV/7O�(?�~��zn��1�J�Q��PVb�$������83��l�2Z-�Kf96dA�V2K�F������1=A�O	��'�?�)��ɤ�!�n𳸶���,�*������@Z��o�:�?�i�0�s�:��<VK�[\���&������Y����V����+�ck��#>i�,+Z�o7̎\����b�:͞�O,ߏ�痒#���&�e�t��<���+aX��w^D���o�+�.�ݸ����*��
������ɨ=$�>fX\n:�F �:�߈�U��G_/�:n�^F��+೻F@�e�=���˺)�瞰σ'��T������GU��M�ص��]�wc�^����.�"���}�e���"�u9y��_��gG�2���rhOaf��+�ﱧ�A*
��{;���(ڈ+TSaÃ4�!h{���+H��� �X����P}B�A�V�#7��Z#�0���S�ԋڅ��O����va�5y�:Da��:b7��,aR�n�(��s��4΅[��E�b�-���A.�����e�� �Cn���>�_+f�k�� �D$^���?�:W�D�I���4��4�?��}w��0������V ���0l_KJ.h�M��!fUȉ�ݣ��(��NL�7�?X�5j]g��HR�	S8������U��,ɥ?S�u҉5�4?^�t�#�����0)狧Y�i׃/��rD�fu�0Kf�7�OV�3��~?�ʪ��+uP��\[�1�h����O�8i�S�Y����nI��S$=_}Q�������|�SAG�ů��p�m�ʳ���&"zn��㴴Z��9�K7�N�"�H�ex���q�Kɇlu���/K&&W�Qu�ӫ4W-a`9��r��h��'lB>�0�GIX�;����m����_���/�@���{T|sе�&PJ�[�s)��S����r����
�4�/ȝ�u�4�[l�J�d�����fn���JX��뻅Q����+�]�B��A��*�x��.U�p�^���T��cnv�m�XL�6Ӈg6����"�{G
^���p�}ZD2�{*J����n�bVh+�3������,�ƍ5�LWҦ��/_xt��꺬����M41�&}L���g*�r�T<�9](%�:��Rt�6��nU;�e�"�Jߝ�?^q�������[]����J����Fbr#�2)�zhz}���	_�ڄ�e�]b���}ݡݙK1�Ek�L�?,���^G�Qo��8����͌��l_(pV��*֥d��	�L�"��)�8!��¯7e�p���=d�[����Wd�՗�ЌDC@pɕD��d�.�'��tˊ��jG�����eӑ�`8si*�Z����o���hʜ�B�v�972Q�g�䥉�����Ǜ�� _�Z�?�j�=�%9d��j�]���p#�B��tq�8�>p��{Q������:stb�cG`/��eZH���8��u-(�����)��3��!�~j���Q��?x���V���XY�!`�$�)�	�k�	g��l���K��5y��r[��q* N����e�����V�]�3Q�?*:"3�˒W����qk��#w0<7x�����`o�����V�e���<qY�7[��)�@Pd�ae����˸�2m������16�@S����)H�K��A~�Z�a	k�Э��p�m��%Ίb{��@3��A�Lbޫt$9����h�s�WjY� [Rg���W��H�9`.c�O�A��Ѫ�7���aC �=�c����;�	�(k��6��想�n��a�)�G���ثN=��7x��/��,��Gb���-��buG��==d�vz��޿��P�M"�Gzs�Ŷ����܅/!�Y�.�+��0yL��^R7���)����%s��j����;Æ�<��=6)ް�2]��(��#)�b��4��J�]|Q�I�[�2�\<���3�v�M��-7�����l�I>�A昱/�t��[$����= ��(O�/!��Մ� K��Cv���S���m�h�L�'�
lx��r�|�0�1��!�5��Z��Թo�~/KH��:b����"����"[����h����E��f���\<P0�kY�F(�K�#F/���)CN-{-�d�NNh~e�^9��g'�6`��<��	R��'��g�ļ?��[�����m����~���gR��z��w���*~tm��:L'���r)��a/~.��XV��<U��tc`m��i�*!PS �q=+̵Y˘�xrk"���H��_�^�Г�̕��ŝ�ʡ��ql�w�i~�W%y��ލ�%) pk鐠��a��s��A����x���L@o�q�$�po0�FhZ��y��rR�4'�4��E0��J��:c����#�+'Z�S�):E�eS�Ɓg��v��^��j_����G�f�����/��ͫT�|�	��5抷�`��f�����-��*gHq��]=�&Э�"'"�=C�!q�����B}���=��ro�T�b���Q9�z�;��m��k@����m5|�R����oU����z��Qo�M^���K������XX%]8��0�,�d��_Wo~:�u:3Q$��2�ò.�r���v�۟�:Y)C�1��O
���hXu�D�����y��E޸
T�'\��Q��}�q�߸��!{L��~�׏"�B���3{Eˠ��k��ļ���6T�$�O�b����~�`���h�k���s҃��U�S�"D�橝#Lcn�2>-	�<�ǒ~�u'3_(��K.�h� цa�d��,K��ϐ���!��� �H�h�^a���D@@`\x	���IP�]��Q�Cq,^���n^�v�f��r#��OO��G�k�j�b�薣K?um�n��-�1]���{�Ս*��4P���aZu?j���8�z��<�>�̓O��E�QW�?�ۖ�9��.�6�q944+�һ�h1��8�F�>���*R��8m�9z2�JU|�aA|��^���.��	H�nOC{��/[�<���6���ی�g:Q&]��F�Xr����u�L{��R�h��8M���6���-C"U�SY�[D�kK{�����y��oOq^\�I62�k>킕b�F�0E7չ�ğ�C���s��N����$*i��|�8�wj���Ҍ&2�媁���^��0�N�3��e�lR�)�b���d-�^�Ƅ��'��,����B�o`8�����D�=nn���?�E���z-/�HP�<,�QZR-�^�I5��>r��p���N�r=x6ƍ�9KqI@}�e���V��F�F��]���Q�]��$����%�xW�<�6?���㧎��C�~U`U��1|�g֣���|���6E��(�vZ*�U�en$^I��*ӤQ����-��@����l�I�o:�2�s`,���hkN'��iJ��^�g��#L�o�e�{������d]���[˭�\,���"�����6��.�X�i�A�[?�R���Fw���-���?j\P$�̋�uFހjm�G����jԑ!W��AU㚰DR�7HK��ј�T��fe��˓���S��pl��cИp����Ł�9naɝ�^�'	>�����Q��O��ieml�t9�s�'K�q�Y+���F�I��?+e,%FH'�j%�;1=�Ss�(���V��҃�<{e�s\m�#�@?�!%�T�u�?�]u�UұдĖaj���zD��'�h��h����&���w'�$Kt��N)ۚ'rjN�� �x�3p��2k�Ҵ��%�({ǤQ��4�]�q�@���ςЕ�.��mP�qJ��J��-<,f�@�C���\�D5�biS�����/W��s��D��������Gi�F�*xE]�v��":4[u�;����.���'�QF!#�BD��9l�È,d��r�¬��P�\Bp���>k�xtP�y�.l��OF	L������r��.ya���*�,��8T�c�ƨ���J�W�O*���Y+z����v�\a�Ix)�������T� yi��M,��A/�j�L���o����Q��VE�L���Kz+bJ?f��Liu{G_;/�K�10�j ��o�A�'W����K����B�;=/�=�|*�#��H�����^S�'�/���':�5�!��6s��[C~P���nC�Đ'�j�t�P�U��R�������3�zA�Ҡ���
V�L��e��YBԾX^~�8)���W��I;)���?F��kv��~,̇��6��f�f¦�HG���A`IOȾ��'�[ҽ%���~�+-�4���M7Q��<��Id��p���cT��:�u�XS^j�E'�0��΃s	k[i�1�e 21�x��Ţ�q��~BL8帹����!Y�"�hu���_/$��O�k��Y��?�,���q�H�8������	��=�lM��dC�+~_i�������
B�麹%��#(���-.5:\��D��F��J�\�E��؏���-�� �RN�2�.��g�8�I!�n��E�Q]&��#|^�Pq����[���t.D�f��y|�2kb1Q1'�S�4�ͨ�s�1t�����<�b\cWyc���a��ԎŦO��!���}��Sk_���9ی���k��z�����a��t�x<�
���󡓉�1�=�mS}{��T�O 2���A� ����dwkf�v{2~��_b�[���5EP�憤�����.�o酪�1MF�(���sOcc�J=�.-0؄_p�5�ٻZ��� A$[�j� ;�������c�:�P
H�y&��˻�a�dI�����J)����^{�C�"�ik����V�f���*`�0�	U��B��@�<���Y1�]:�ܽc���e|��@D�H�w��9�A��H+.n>ћ��?Z����	%�O��v2t�t��j���v�������z�g_�H��.�yAQ�>R�0ͫ ��+�)��X	J���d>"~<tm3�!5����t��C̎M���$�%���Ԃ��Eb��w���ݓ)c��B�D��0=��}dCR `�ye�� *Y!�4!��] ���(K�d��sF�2V�UP�L�u1��Xp��/�B�e�m�Ź���T/.$}��'@��qx��Mt��Q�^�DV��eW�H��uc���h�ƶ�:{�0��s��&h��e� ��(</S=p�g?>
�]��@�����**��۵Bg��gرM�Q�k�H��8�շ4�B\d�Q:o�h�9��|�<%����
����yn�+?�=�p{�-�t����6Wcxu�~�b)�uĨs�d,�-pO�C*|I�?�I��=pMƉh�z�9`��\���������e�Q��(Vu�Fp��Ć,i�˳�!�C<u�}�̨�$>ȫ.���bk~�/_\�wa�|-R��� ����}0xT��i��9��������FX?9�ca��p81�+����Ʌ2����Kٯ��7����+~�g�E 6Xԓ����6�xo���繱 '*�a�FT��y���C��F�o�ސ\�"�)ɁH�RPw5,�V���S�d=��`.
`�/���aA���+n����\����Vo�4��U�SS��p_��Cb%����c1;�R�12+^~��<����Y{��ő���М�Bp[�?��D�3�^_3)�b���KA�n���G\��A�X7P�[\H�j�m�O��4��{�fHI`�\x��Y�����\9�/�a$=cv���e�-HƖ>��f������dp��)	¯���tQ�÷|d�Y#�V
��\�'$��+2e��)�{�J��<H�7�kkZ�᦭�2^o���Y�5l�O"��z�n}81[��R��u�u1>���b�t"�`ln�d4[
�|�kW�O�2��N��j�c��h����0��»���z��}�1d�v�?PN){��rL��	���]q�,Fa7���mu��D7�?��Od�RUx.�U\}�fZ}���a�c�ˮ��W	�CtF����\�{�tp�s9Y�06������Kf�V�C�r�81q`��S|#�����|��,�Л������T�'�}�s�v~�e�������P"̹��R�+2��5(&a��[��9�ٚ�Y��%a	�}��h�X.0Y��D�ACPmn�?p�T)�CQ��e��uɫ�zp�n/��+ib��M��]��FHS�v���..�ս�IYl����ż�{����d�\b�/�c��/P�qڞ�쀦DQ"�b�����/։Ə���(\����U�H�������9�ahu��NRH�֏���g����W�>^���d�pIh����`$0�!OBDWW��0�ڨ��f+���5����o�_���%^�N����9�տuw�����}���VW��<fQ��0>����yXE��ЪC/�����"1����x�M;���C�*��϶:4c�TC��L����q�i��4F��_��ew�A�҆)���V�9o��⋏��u+����L͔*q�a٭�*i 9J��p�S�àF:o0�M[z��1���б���ӖP�9�)�� �c�=���@�-���'T�"��'��RPT�`��vV����,�������+V����l�)����"s�;Z);k�Q�o@������ݿg�)B��8��Q�w�A��nRH�nZ<X?S���z#/�o=�,�8�t��FȾ�eq"({3ٽ��8�Q�����)}F�֌ɑH����>F�wQ<�hj�P�<s�g��E���\ \��Q}#���ͺA�l�F��-�y�'E��^0I�����q�±E�ؼԐ�mH	���v�2~��:ѭT�r��h/U�dK��)��U�	�3���+��x,������@'fd���ST۩"���eW���-&�&�Fr�Mc2�3���TKrP�vf��bl*c�[G3��@�J!���n�R�j�+��&�ҝk�vAj��0�@ٮ�������D�-#�cd{G��M��G:����!5k?z�����
�O���9j,ikn�-b��*�_(/lY=+V|]����nA ?�\�h�_�È:��w-���P��c�}����Rar����.��
��>�ŎY�G��ʨB~���֕�B�gKSH������t�`���
��^�p�AA��g8�WӾу����-�)�5���ѫ�짵�1�D�k~��q�u�`E7�W�}f�~I�lK�����"�{r�_�}�kN���嶚�3��U�y�˲Kx���[�Pt���&��&,֓���lSY����]��Qyn�\���)ӷ�JP�	(}��e�>L���r�a��<6|/f���_�� �}��(��>aU�.��>���U^��9�y��d�u	���T�d�ps�d��T(X*ȣ�W�Sw=�ѓ|qp�\����<p����.�s`�[Մ�K�����N�b�fm��)f�p��c�(=�s�v#:����G6�H��v���d�:G�k�\���2͞�����7	Ŋ�#%��b)4�g_嵪��4fi��~>E�PG3�-�@-5��u��� c7d��e4�%Ч���9G��[<�0����zWg�;�]���e1S�i���\x��	��#��飪=�^s�XLc�Bߏ�N�6!�z;��L� ْ���Fm`��Wd��N��g9ِ6QvQK�%�~}+>+ü~j���$��$���h�ߢ��p3Y�Y�;@|��	|�H� �Ć�%U!�-H��d��RVk��->>v��Q"a��>����J����ǖړ����sJweʗ*	�rBk�)�K/KI��Q4�	`E�҈K%���f�KĻ]!�'�=�ΚF�$_�n%F��W���r���ꢩ]��d�C�k���D���%c�?;k+Z/^�2R��d�7��k�x<���ah�O�Ü�]M�y��	LG]��#aJ�R�!3�ޠi�4xg4��a-Aʟw��ge�Z�o�,�Y����XQ��<�����{�~�;�y��	,m'���-ʡ�.9�3�7���>|�i���N����&�bpN~���$�ǉ��pL�L+a\qg�w��T�SRtybP���ԭ��*"�8��h��̈�ߛ>�L��!�@���!JǶ�A��3L�Ha()���X�`V G޷Ҋ��q�0,�*��S/�Yvߔ�|��d#)dG|��"ѪL}���B7����(_P#�i:+��"Vʣ�MG��*����2��|��8�Z�)�)���˘<��?�U}��+�pS�y��(����7)�oCu>�.m'ɹ�_4��Ox��}|*�H������]����˼��(o'��9�^��4+��2���A����XzےCM\��o%���F@��{J�T�������䮪����p�����s˅���=p�D��6y?Ű@�P\�'ߢ{K^|$����b�K&�V�L�IDC���8��rg�ڰK=��f�B}`�������ƙ �	 �6�6���8ʿ��T�jS֠����XH�(=��?��y�G���~����N��q�2pKo��cf_۠��^��������cۓ�K�|T)7`\s��	�G5�	,�?RY��ؤS��3qD�->�G��0�Nd����Α�E�h��(WnkN߄�!�W��9��PыaLp]�`&�1������ڜ��]�SC�D,�q�~o�M�ބ�S�{w/̱��i�&�d6��m����'vXqj��![�2���?=#*5)$��{��*��&��_�\��l^T�������Lw�Vlzz���ն C��G��X���ԒM�J��ѩ�nS<�$��k�56�<c�8+��e�[�3�9�!/Lz�x�S,��ƍf���K��/r�酧 1I���B-C��	�݈��ΐ%�}*����A���5��(�r嘘>����??ﲓVQ�#�I�L��F��Jr`�2�Q� 4�SBl��_%�u� ���.��� �'�f�!�U��8P��E�4�p}���Ęe@��di_q~�̾��+!,�H�f��
���~O`�3�zd�>$���
w �y��%��P҇q�藷��Q�g��o-Zt�G0{�E*��q�0|�Ơ�O>�ˍ�۽�����t����f�gI����S��F��Ա�ќ~�.Jv��������fi��V s���b�	�*}]Qj)ժl���|Կ��W��:�dJP��|�����ך��@+��-�^�V���z��#���������f�D�\V ��HQ�@O�*&{'�;t�&�Ɉ��lޕP��9��' �O�n����kx�L6	�*t����Di#�� ��;b��yūE� ����Kw���6��`3�t�	؂K��������L?T[q�>D��� ���� F�A:�����cKo���hCZ�A&�Ҕ8Q��s}��jh����P�����؛R�4;��C0��fn�ڐ-z��w�2��\�q���Ru�vZ���J�ϗ��4\�k��+@�U���^�U�^�GX���5O�7��F=t�Z��(��3{�9I5d�$�q]J�\ޛi�l�V��~J��i��X��(u+���Ѯ�+�l n���"_O�u݋��Q`Z��UN�3�+�XЯ��Y�^�A�n�zу�f���	}��`%��z��Z�|��R%�yۑE׊�+��_8�&k�#���'�1��*�;{:F"9.�/F��	"���
7.��[W��]KN��n���#Jq�}<i�5�5@!�#�`��&-ݜ�U�8����J����Z��o�a�Y���1T�-<�%�wg�o��_ļ�t�Z{,�������)���4x��BA��Ŧ���E��,�ē]�8��UOm�<���\eD���4W��t��]��>��<5��4�.�f�/�7����.�rQѿ[T����b>�"'r�ت5�ա9v'�9}ڌ��r��p�x�)��^���$EVf
7Jz��! Bv�������<�愿Uu�V�!��!;Gyi���RI(�Z�����½f�s��&���o�`��lC3 _	a�4r�Q���S����)�p�3Ƙ��`v��/��D���T"hht���"��q���R�pSu�g��ca�h ��t-�Y�d��<`�GD��L�]C�⪳"I�>Mڛ��͉�g<
���&�x�a��	�b`M��+�������w�?p �D*�ۀrkhx�Մ�H����Ф㠘	S�?0@�L��5.�o������� �O�.ʽ���J���4C��^�lq�7��	�;�\�o��c�dKh�,s�s(�#*;�����GG���H���sqm���H/SQw5�{;M�W.�yR��3��y�����-���o��V���et��FЍCP������؏���Q�C�w�<��P�'��C�������$��%�'L�.]~`%����^A����pO@C�R=�ǥ]��i=������".�h�`U���}F{]��9�� �q��#Տ˖���p�8�8�n�ᚩi�{Ǣ���B��p>
�H��Z�h^�D�Iy*��i�M�f��Be]�F�gr]�U��aM���1�wC���8\5���ͧ�]sV�$xX!�A�O9[)��xۊ/��v�Owh,\тE(VT �d@_��	��M���~3���9C``��%� ��Z��R��2������H�{���^�f�?c�\�5�Յ�e����4�qvE�,��U~^�d���_�w6��I�C������T�Y���Gΐ�J ˿�K���X��e�`YC��P�ruM��@티{�B�VvE%�sSJ�~"5ٙ,�o��=�M��`����+�`����Ubq;�e���bK���6��g>��8��V�a�c�иCH���Q�H/��h���T���i�������d�{,c�+�b��DzZ��՞.)��Iy��a���ZNL+���T̈���[t)T*G-	��2GɌ�QC�=�8�_��:+�|M�-���Ꝡ��̇��$��'��O�<X�͉����o�lqS'�Qό���R
f���d�Ӱ�N�_[+���`s>�7Nq�],�r_l/iw%fւ9��Rk��L�s+�(�_
���"d�B�ۚV�om?t��eB�T+) �tLv�#���7�j&��LKq��ު'��H��s��d}����`P�?�l|+���6�@Kd�jX/��
��-�� ��7����p�ޤ<�㱏[�h:%- �8D7m7+s�2��Q�t��)VѼ��y�D\
?��|�g_���Ӎ�)Ha�%�"���I�.vL��S���ⴵ�f֓k��Y���p�JA0��Yu5�3`�@	��Ȩ��m�pT-cC��Td8.�}sQJ����!��}���T�kS"Ql5�a-!f���bXZTD�52BV�2�=��U�ӝ+�J�:I�=)�G7j��`%$�1���A�b����s߮�R�j���Wz3���dtG�P�*ǎ$�Q �6�V�S��ɒ���}��_�b�q9�`����`�5+Z׬^��3%ɥkD��Y/����ۇ���Q(8Z�DiD�w�24=m��8���|pc�U���V��29���	��o���C��[�|K�.�����A��,��&���D+����Vz��l��*:n��%݀�4��@a����`@�.�������hh{�0�A���l�-V
þ<��QXh_�Q !A���5~��S�D)����>�8��! T:]��sMq3#goZ��
�#��b|�j[,���K�O
����OW)��5w?���\�tN>eT�G�V��9������J��|�ě��E����/tʙ7	԰��`Z=��"��无_S���>̌F�tz�VP�a�'͗��PYk4[���H����XD��V82��p�*��XQ*'�j��A&���b�Zg��Mt��I���(.59����ƗE&�Ц�:xv���&6s+R_�ס'(|����G�����>��ȉ�~�S�%%W��/�78O�~q�gp�T�/+��nR���'Y�r^����N�����`�/���z������Sz�@u��(╕�I�Q� �'�^4'����8
T�8_�����j=.On��D#���z��aQ6������wel��Ǽ0O����Nţ�&�R��A�,9�3Õ�ڒX*�G?���0^�f�%��Y���*��}Y!�`1����D�����R>���[\��w�X�[ou��f��iA�+���2�hd	��'r�ѷ&���o㎅:�$�Ip#���	YE:��,��i#�a�#��ޥ�Q~���X����nW�I���cAyR3A��~�������oO`Դ���]����J�����v�%^K[�X�oRZ����b�.���:�f��-�3��+��
����y���E���eز��1�V�s�L"ɩ�M��Vrm�^�1�;s���9����c �8y���0{j���}��w�d@��O���I�I�� �5q�̲`6�����x��hV���Ֆ"�:���~�à���Q����7CƘXy��.@��e���t�;A2�� �I�؀����u&��y7x7G|C���/!���E:�ts^9�����&�Q� �4�}He�ͽ�%�8.�It���!�G��Y����+$�FG{�`����-�c}z}�v���sl~+7��C��E���E#��Ĝ'�p�o��Z���c��J�]�r�9h1o�h��[�j��J��᳴p�j�d���+myT �;��ˡ�Op��� ������bN���G5�&�8�.�KMu������ۂ�nW���P~��עǇ��E�f!d��,�i�r��i4tE})WK�bc�����O$I/���)|�Sw.�.���' �q
�$b��N��⡖���c�1tý�G8~���KŮ��1�m���� �,>�wdU|d�mSc�W�fx��r^/�s2��e%a.��!���Y�Il*2�Y@> �A׌��C��5Ԛ!�c�]�.Q����ߜ�̿,!�!
�)���PA��YxY��#����Q��\���I�����jz���85-�o�T/�� Ⲭ�G�۽Ftδ���]+��~J�}��iS�IDj`t�_�Њ��e"�;-������@m(���^�h��gRl��1��OX�(�|V�Ôny�����t˩�U�U��3�!j�Ӛ9��AB��m/���\��6���e�yf|�e�]�`���@'՟$`�^����*�H�0]��4|�9�{�&'
AR�Zm�Pр����bF��2�u$L����c�Y�(y��a�q4�K��DC�+����-��Me��'��cYU��
m���Ӻ�ժ'�`�Ə��QS&]@�aM�ƚ�d1F�_�{�a�\�W�c�@e5�a��n�FR��'�ѭ��L�RX~1�4��
dڟ}J�%4��'�$񌃂$���`*;-8W�&Ƶ�w��,Ba�=���q�,������v�s�sڶ�-W��ȣ�IH�F"v��+{SA��&`��hZ���M��c�+��w�=e#3��G�h��0���bD�����B��&�َid���d���t��C����Z��Y��҅�b'��_�E���튂m�n�p���P5�Y+�_���H#)��)q4>lx�"�"�rh}�z��z��v0^#�v�&���$ug������=��1���`V�ZE�*{�ԔM��u슃a�?��g8���}}Fe̃��O�IM��t-��o=�Kqt����.�[.�kt&��dǱ�A�ki��^sH��n�W2|A��q�1�k��m����E���&�A��iI���K9��!��%*.>�+;�z�����F��#���e4��*���w��Ȯ����epy�T:��Q���nT�#�ߦ�j�Ɠ}��v�܍<b�n;hϱ��m齾gdU�ɓ"��Oi�NQ,7h	���:� �y�Ca��5���%"�צnd�Gl4 [�?�B���7X� ��X"������6?T�
ڥ�72�\�����i�Đ�l��*��q@囉I�a�a�慎����Q��s1����mj/�h�6�9����:��C��P+������Ѩ��ID�~O�w�������k%C�N���=~o�f����of�ır/�@�ԫ��ZZ�!�(�[�a��4�	[��#be�u�P�Ig'�#]O1$���FL��K�#˖[�w��?��Y��=��L�w�����iL孔�2{�Ml���縙�u�*P�I���y��ބ�qs�1�5!���8�I�L�1}9�~l�w��R����c��_�6"uwj��2���m+<,g�:�F�Md~�4�wJ_�>Vϊ_��f5@�v�b���Qd]��h1��J|�Hd6�G)/3�&�or�%y�̉��%��&�"�U&� h�q���%;w-�-��P%�a^G���q3�#�@X�y�b���9��H�% ���ך��|����(d��,>�_^��ͦ��`2[/�mj�Q(t�Ϟ�f�F�l҈[!�F�ހ��Y��8J� L0��G��/T�l�k>2�t#I�l�w�
��Ց��tn��O;�@9z���D�,������#���Wn���a|���I�D�̒�Y帝���CJ��Ԁ�h��|�����Ra=���J �l��Jq#�#��1o�'ʏ����9lH�~9y���v����qM�H�4+^�_q.��>h�eT{��,�4�O0=kB�0�!��5���٦A��,��������P �f$;S�R[O��Ҵ���0B�k�vx�ܯ��뽣�ɨ9��{E�%L�Wr��C���n!/�Ԅ�:��D�@�d��H�	��T�nł9��<(��oiɮsE��d��#p���͌/t���b�v>�]�X��rY����e3�5���d��@9����T���������7@�^=�g��'\uo�Vf�i���4�G��_x�Ź�+�ZG�>%ޑ�i�(:���B�7$ߒ�Y��`���Ҡ���@���˭_�{k�0����g�9b�-��������y+�~=��.�£��7
QB��u�H��5��JAAu�<�Q@�>���j��;�^&�]$�#��q��t��t$A(�&.�p?�@����� R>a��b3ž���i^,�XB$�����&��2cU�'`�z�.p�e��$.��� s����A��>�,�9c ��咦ýo�W*��"Q�_j� �+S���d��$�2�c��&&��B�h�����.Cbi6�BSH����D�WhG5�G"�m�u�le��E���M����e9���cG�=�#A2cP��d�݄��%�>���m.���I����p"�����KJzM[���RB[�����RO{���JX^��?�e(E�M�b� :G��9�(��4�͢v��c�p+�>���t֒aT�,a#t���w~Ȱ8�@^n������l���%Z@�TW.��^����B(���/�!�m�(���Nc�b%��\e��A^��8{�e�s䄸27}|'�~��W>�	�q&7Ihx;a`}���`�������ECLc�<�X�Bय़�������$�7��01\:����^d����r[hAi��c�g.���]r�m}�_�1�H�C�����I�ң��<�����Z���� �S�~���Z���K�NN����Fq@�����m���,^I3 e���S�sG��[��[�`(��L��iE���g@�B,��k���$���O�98�@a��x�*Z4�6B�=Z\b�02�_ߎ�!BN(��۱���'�ͥ
���^+���ed<ll�2s��v|2��R��x��� �]%K}Y�d���vQ��˶�FR��,��5�/�v�o��� ������� =N�LҁE�c*>[��p��]~ˌa �Y=���Ȑ�<V�s��뢳��S�y����nb�*ߠ�Ս�0S��yPoj����Xx%��S�}-�9�u����xR[��j�bͲy ����9�L������'C������am}�Ss�
��P�O���=�мx߫.�����D��#���J��o>��� �cs^ky�4޶��|�`�Z�����&��
=��"��)�|G�� u�`H�}��(��m�:��qM����	qR�ɢ�}`2@�R̥���}+V!�w6n��4��,T;q(v�MNa�Z���E���I�
����:ULzH��b�ͻ:&BLd�Y���^�L�B��dVR�bE�_��1���X��}Ad*ۚ\k�
k�\���:�oI,���C����tF�R4��������o�}]�<��_��Tm�L���1���)��rQ��~�ݮFU��b�&�4�~N��d�����f�_����%�i;_�e��-j�B������bGT=`Ѻ�)�G;�؝��^R٩�� �dh�@k
��;�r��x�����@���ČD٨�[B���Qf��q�ȸ��>���D�G��D�)N7u��ǝ:B�\5^��~?m��6�W��%�P�ڗ��� �Gâ;��� ��oG���XM3��e5�M��0m��I�d�$ey��j��;�.��%�2��r��o��+o51�7H)"K��[")��"�H�̝̗p�&O�%EP���޲'�R�N�� };j��8��a*�g�]�CW�H�o�ݖ���o��	_�ۣ����T0�~4����ty��z����n&SJ$�5���@K��hV�*$���S����oC�e,��.)�f����Z�ѣ����Kul>���mf��<�Q��ADv�(�3��+{l�;�^���Qϐt:�ဍn�X��0��6*j( r�ȇ�H�Y��5�gz#�_�zJ�!C�x䡺~��GC劏�P_@\��ս±r2֛���b��ØN�&

�����uT��!��ұ��N?��V�p����^FDz7�ͯ���&�̤#�6�Q�m��w��rP�1��k���L5�K�=�������H8~j�I��3݁��|&OEh�V�%��|�o���Ej4d�/� ס0w�}3��j�b�4b%�x!3��IS�Ã��	�z�̋u�͠�Dj7�����<'�`�wi�?�g�jρ��ͪ�O�o�n숶��G�K�3]	8]ş��p�E����)�p�ıB��񤢨�R�Q��a���:y��S;q^�c�=�'�M�FKX�����"6����BT��'�_��~癄���m$�o�� vrE�����v���*�zϓN9�+�\�`�3��9������/�8=�>�|=�~��(Dd��e���҂��E����K��R�����;j�AgoIn�9L��4Ȳ���jS�k�]�R�Sz����T���ݝ�@2^����<�e>�N����V��!hJt��{��vs��r��$%�rUݕ��'��	 C���\���xŉX�
��Ul߻},�V�s1+�p����-����M<b1,n��q�$~�~��w�)���z��: 3���X�ߕv@Z={�F`��N��Ar����%[y�@A��{n���MBJ���au��^�L������VhOm��@����7G8�>r 
L�����8
SP��)��ː9�f7���*�R��sTvRĕv�ȕ`�St�4mƹD �r�(9��~�C\yK)w�h����1t�)���a�������!�xJ�$�c�"��4���i��&�v��]��Լ�j���2�U	� |'>��{�Ӕ��Z�ؙ�����БGY����{[�w�Crdc&b���e���E ������<v�+���h�+�5�N���d��nJ���	�)�-=����;��n��v�+�����7G��1⽈��ǋ��cF����ɝ��h�n�� G���??��c�r��?OEz�7��ǀ�R�U�o2!Z�B�Hr�_���y;	@��ʤ���M���}u���#!��{����F��^a#Su�1�G���8�$� 
'Ol��?x2T|Wk��9��:s�<ұ�m#���`f�]�Q9������т�颕pZ,E�����T]U������
x�C�w6��ցO�,��J/GC"�UR���P�Ny�bm�]_���X�������{mm���/�c�FGI���rݙnd>�m)dџE� t��EH��r!��^�o����W3'2(�lQ��%�i�~�ՓA��s9���"S�M��?#��j��Ԇ��X������.��$���Cy�K�Mj�_F����
�ϟg�xC�ەV h[L��
���f��S䙦}�E��'U-��� �C);#���$b'�n[U���e���s�퐈?2k��3�i����|�� Y��X�7�[��]�-�C;�S�#Oz0��琒�w����d�-1�?\���J};e2j/���s�["z&T�m�~&*A#<��㋠ӳz�+Ѷ'xo�K�L\�S���9j(_u�����U�Wq�-�ў�cj��X8�{��6�D����mĠ�Ni �6,I�������!���]�M-��Zx�zw�k��$j��P.1��n���2�DZ��:���|�6�l%D9g� �{����uv�pJk�0����hR;��Vd�z�Of��w����T��J>@��D}�j+��~�8��-�Ϧ_�'9v��-�_ڔ�=4��M��	N��q�8�:4�J�Ei�}^�ؙ��En"|Kմg�U�l_R K~�S!B6N��6�c##�?�Zg�M�sWd��3;�X���r����z���>N����r6�sB�ћ� �t|sL�'r�z�
U�8AQ͗}܂�z�,a��`OsGB�B�= 9�ø����7���5)0���ܮ"�0��UTwq��$ ��t�XAUL�
�;N�u/�ꕏ^3�;Isd7�^*{2�d,�KMn�#�Vݾ�����x�ߞY#x�X����$H��]�[ȋKuux�\�_���"�d��gj�v�K�I��va*��A�d^��5#hH���y|P�(w��M�[D�XI2pi�u�I1ف�b�(�����3CF�	Aj)My�@mv`x��!j��~�Oo4���7�wn��Ǭ���c3)��e?���b����������m,��i� ��H>9k'ć�E��=��C.>l"��e� �4�B**�v�Ķ6�O}����z���:�L�36��VxD��_x��!��#W�˔������M�_�Q�b9��zZ1+0O�z�T�V~�J2��R��`f:M\t��`���c� �.$�=�[6���q�n��<����6���-¢O���MD�q|�a���zE��;*7Ŝa�FQ�/�e�Zgj0��N��uc;��
�5gA�"�Nנpvv��{��̍�@ch��6�å3�f��;����"w���L*LbJY���#�P3�%E��9��)�q�k'a����!d�ݵ�{���h�[�i] Dm��W@g1�k9Ń����V�.V�l��f?|���e:�������N�)��o6��[n����ʡ�	|��?����{>�J��=b�4���n~/�bV���S��t
�t����il��p����_��n�Р�& ��Г����(hv��yC{�PϷ^L�v��y,T��^�C����h��JcKs2"gcǶC�o��^��<;��?l.������S�|��S�ݎ�����<,+�gb�{I�ytUu�xʅh7����%+�C�#>r8my�Bm��*��p�d����M�3(m�Y~-j{�L�H��t�8o���vچKPUD����(�V�����gz���������i�u�����G�D�W�`���[��a���`�}�Bo8*o��ǄY<x��f�I��c�=^���_]|%B����#����W�ȿZ[x!-�������r0VS{�s�|{%���߼��KbU���l%70���Z1�Ҙ��H�Ϋ��s������I[[������� 0����g.1��N��&A�c�Iv��]SnBh\��	G�k�1�2�f��mT�蹷Ȭk��t��E�'툢���i�^Хjؙ^�e ��C\E�q>e�YO�z@!�-�^�����^����-���Y��2t���W�ӑ�^�����6���a�������R玭jV�azk]��\� p�#�,�}��6��ߴ�m��>ѶEr�O�/q����h1��:��<��>`��,�hk\��*W�����ח�Ue�o5���OHsOq�����]����6}"̖ٜټ�6�j�S�U�$z��ď��2��s�P���j->u"L�o�3]fP�yX����������眗�i8����b�kYsPS�\t�7�o�h�&��utbC�r| �*�D�(�X��>�X7׵�g�v��q��Dk�ٗ��}���s|ZI����m�L���N�u�ݜ�z����}��t���Mf� S#�~�e��#f�g�>�`j{|=�<�u{�_��zK	]���>]M��q�[H�Y��kT��r��s�G(�_@�� H���R�W�b�u�f�k$A$حz������%�lzo����i�τ���]H}�Nd�_#(8y����q�r�A�|LG�1=a�~!��"�>�D���3�t:��d7�� S�}��f�&�& *Q�_h��@�m�yU�R���-�ǉ�=�fQ��鰠mo���K�p5Ť�E��#�X�AM����|� �@�A˕}�w�w*.wl�����I������O)���|��^�lq{�@����V=ln��s5ƒ�������}t���i�7)�?N�'b���v�Nqy����f}
��xI�Y�_JH� �S¿����Y=�|��vX��]�k��Ù2���&Wϲ��я�0h�X0������p�����R�������m�E>������(O�0ާ㌁Ǥm��)`�W�>��u��]|�r�j�x��x��le�P��_Ahb���l2�
��N��g1�<A~E˸�"���@{��o�႔Y���6�P�犧�������x%�ER�YՐx�\�n���5�R����&���=��[n�7~�ykv��!��hc��l� :ơ���)���A2��F��ܟbA�L���zm���rn�s�b��Ag +� �d�\C��u��h�/=����5l��i|��8�čO1���4xQ�S���r���e�+\��0���n�I5|��GO^��	�ޔ�g�_R���fn���X����t$}x�沟�L~����u�O�h�n���8�-�[Og*��K��㩿C6����J���|%��`|O<cܲlh�ng�1��%����օ�1kI��2�D�ml\
�9�,�����P-A�"F=K��'�m\���3�<Z�2�m�>��I�$��n�(־J)���$T�%;�@��Y�X���D�duCU�۳
�#4Í^��K!���Z�s��C ��EP|~�R���d��� �U�)�i�>N��|�!!n�&2[M�����T��3Z>�S�2Jq�ekӬ��hUE#���]���ȦoT�[a1&r�R��.}�)Hі#5mŘ�Y� ;[�#X�0�r��!�Z�eU^��+��.��}U>�ߩJ28�
4I	��h~N�]A���e�1{>�[�
k�b�d b�֦R6�[��U�U���O2��~p�-1������n~�Pf;���63`ǒ��dǗ�V-z�>��6�YSqz��0FH�:��=ų�T���GK7����Ȳ̠�$r����(����?p���}s,j�=1��ʯE��U�l��q8�T�����;��!e��ǔ�G�{�Ԑ6��m'��`׉�����Z�o	߉��q��׻C��`
���.�����^ *N��JIH���l���u]T`�����A�Vƍ��"�K��2�\�/@w[� �!�Y�%C`�����0�˜nq=DR�ד�y-�ђ���>E^�1 ���za�+K�z99W5��� �͗#+���|rF�<��C�}�ݮ��Cq�.�G���IE[�"��;�<U�'D������no�>��0���Ѱl߹}-&��F�< r�0�Ď~F�ڋS���9���ؼ={��+�~8�&�»�nַ�������q2�ԥ"��d��u��y"ވ�`��
�ێ��dq=j�a��b�S��#�4$�y"}�hGij���8�u��L���G������"hk�Ɠ�!i4T�I�Ba��/��s�.-���(J���+j[��JO��O�>����\�tL>� fzN=�`�X�K�q�t�,E��g*�?�e�B�6�+�Y����&޳*�B$;�doh��w�.lK�L>�'	6/AV���IU:��@u�U���������>�ǆn{?&hcY����_
��~��b�Q�l �)XD���G�[;�M �G�A���t9}�@�� �Ԓ���O�d�4\G��4�t�ͪB��1FQ�B�Ȱ�J]�	����w�[�͈%+��߼���yIN���գ;��gG5	D�e��c�W��5/�L�|���쟠�2���Ob)j�׉0hÂ�8N�l��zE��|2ǃߺ�H�L��8� �I$3��;d�:L��A��A.�pc�D%]���J���g�5�oJ�����6>��U�_ �`�ɭ��m/&bZ*w�c�U��������u!{����/;
&7UC\��p��f�2��XS�F���Vɠ�*ӹ�&�s6��_�w�X��lں!+L� M��tsL�r�J)͙X��Cc�Oc���j��.M���boҟ�r�'v;�S�>��0O�c�G*�QR�wţ�Ntn0SEJ�Զ*�9 ��Se1©��1�����x����tN?��m������m��K�&�'+E�wpp	�3>}�W�',�"#1�]�
��gO��%ᑛ�Q�g���WDq��zr�����YV@d,_`I����sA$����EbV搨��}�E�C�-��ŀ4�'(2<���b�h���(zX�з��^�Fب�{ �BB>�x�������b�O�4?"��-��a� _�	!0ō����#�&f�dw�U�Cv�FE.���W�d!�\P�-jLY/���Lt��v�;�C����Q������| �,��ၑ?C�NXt���֪�x�?j��M�s�Z�z��9���M=�ǯ뽳�Q��o�n�I�Xy��Eq!^��$mMp��Tʨ����Na��a+�+v�?(d*o&e��(�dx\��z�O�� ��pT�KǤ�T�'/�m?��`vY�֝K��ў�k�9����j$#�k̟~�%�K��O���q���*���t[��s��?N��<�h��Z�"ZȖD�{}�#�5V����·�w�BG���}����'<l>�4�@so"�DC�u�5��&�� �;]�OJ�_)�,���0��<7*4�p�/\/*$_��~�8bz�J�W���o�&��5��G�l0(J�#R;$�0�,�R����i:�E �z�X"kI��C5,;W�4�hj��&�[�H�9h��XwY�ї��ă���@�F���E8��'R�T���WiK��-��Й'�%�����a����q�� ǡ��v���U�ٓ5��U�oP��H�*8r�����W!��TN�t��*��$D�F�S�Q�B��L�Z	��%�EN�@:,JG�鼈��O������ٱy�ń�<��	�wwy�?������[i�!��ײ�P��ie��D�<"�h%��N�l��38ųfK6�P�;l�*6&%{Ȟ|f\Aq<3�><;!������x�ﱿ��@��g���	MM\��U�����$-�50����f��N�S��}m�<� h��T&g� ��_K��<�@�`��C�F�6{��-N������I#�D��;�y�X�!P�}�hz,�w͠��g� ����oѮ��l��w�3mc�8�U���+�x-���[2��vw&k�;�f$nu.�xZ�I��=H!`���b�H`Ў.��장'/6�*6S蜐OZ���(f��!|�.=��������#;����,�����b-x�X�vW�i��=����	x�-#����Y�}t��	�w~��C*�t�O1�[P�����x�F+}kI���������|�@܇������߿9|���O���vV�+�pV����:��^�Ċ������<�>�u5rM�, �!C�a��n�����IzK�5�FC��ٽb|�f� �xe���4h�9��ÀP�≅�)_�75�/�`��'0�ŵ��,$�̰���7Pp��g>pÐY�qeE�D9d%��m2��Mr}!�01e�{8[C+NC�=A9k��P��O1@��yؠ��Ө >6�Ct$*�$!�@
��@+0����O�R���Z�%ס�Wj��IP�uZ9;�����#�"8�{�_k�s��z&��x�b�]�ɰ���Fnt�;��e��|�� Sq��B㮜�Φ;ʬ�T�]ĩ)�V�G�E��2Ij��K���{��~��H����~G�~d�'K��/*nf��î\;�ǜ@J��y(�i��z��)�_7=��[C#?�/-@b}҃�˳�蟵K92s�`/Ks�R���C=
��mg�=e��2�c)RtR<*f3�{˟�NG�^n�`	E��'蔕��d"x�8��gɯ�u��-O�����l)��z�0����6P��'5�|�:�F�� ��x�p zx�m�Ek�d��$�K�V=��)^
�tS��ۄlM~��E�;P�DO�T����17�h��n8z��z&V0�<㠯��cfG�%���05`�_�)֌��l^x<zݻ���I��ɭ�uM�뵚�;i'�P�ӥ����d8#.u�-�Z 
�#s�	�GB��D��aD�Z�V딝mgh۩�����?�/��[�4ש�v�3�=�ԧW�������T�?��{l�M3��$��+YiJ�Qh����T�*m6�G��˙�E����U�P`��
�[4W�H��c�D��΄4�#4�f�k���"xga���]�����T�w�_��eg���ɾj˛L����<����|r�������L@6�Fe^��g�O\��/0V.���gs��P����X��B�	P��f�/�j���c��[�(�;��by�Ԥ�p�L%��"��R�8�vS!�Āc�D (us8v�m|���Hp�E�[��G"�xG�%�O0FJ�|��PZ?�x�j�obc!�5�_���d�@J�S��6��Q�pVf�c��(��_/y�C�	v�ض�d�EO:������ J&Su�,�t��vT.'�[k7��<r��ڭn蛃�!A�N�D���B �X�0�'��؀�"���GV���Ϩ0�h�uUϮ�,t��W{��;o�w��cҞ!%u ��\9ۘz��������x�]#��63>S��2G��������_�5�R}��A���)�ds�O%gR��JHJB�� ��ky��������"u���*n��5�aT��>�v �enCK!TNrcr]�$�}˵5<$��nN��H�r��I-�T��:�r�ٿ�ߪaA,����7M����>���Ϟ2�Y����c��7\���$q��a��p?���R6�Y<������7t���=��q07�t�ʖ`h�ְ���ғ�J�\ο�0fᮼv���"I�W8�m��^�DXe0���ᅣ	� W�L�`OO��j<�'�VD����������&Ū8���ࠡ��kv�9�$��~�AM���1�o�,k��%8.8��f�_� Xu�x<s�\O�"��VgP�iq�_�^�79f��y�"�~�q���{�֕%r�����=���'T��@[�e�X�zd�S�;����0@a�O�dGz5F�wd�)C*�>��^�a<��u�f�Ϻ6�㸢������7��,�c��O�*(�C��(���;��{!;������	OmuB.�=��_�Jgs�¡��?p���f)a��;��D����;���7�&W09��I���c�5p+���떰���+'�gʉ�W�z�:p�3�E��˸�S94��3���3���mW�����Z����ԕ��N/���
>R���ͽ�VP\��&nJ��>.������Tbz���������*c�ԎBf`Hzp)������,f�?H��Y`�/�	A\����$j�3#�P21�T�n�ڲ�/�?_3>g!7��`��k���/�����X�/l`�������R/��E fm��ZNi��Y\�w{��#W0���w:d��s�- �S}}��(� ���9
�aDo'�mI��3a���d�؅?��ǣH{��vD�K�v���~z�i������W��K7۠��*��)Z����(������^!���)���hS��
��'Օ= ���+��K��@;y�ԇG╢��"JWt��	�d�_���� ��ͷ�a��?r�V]{+��x���X�ZQ9��W�܆sN""��K7���{�)N���cv���)�O��3�����n����6��9�&Y�QI�26�Ƴ�0��}�*Kr	���M���3�}��z�W�7��l]+���M�"����Q�6�yP�f?��,�P�p�Uj�	?�R�3�2��tW�ސ0��)Ѳ�iJy�]�B�>�~|���S�~s��إ��7�6)J����ْ���	����g�Q�Ֆck�m�[0��d���/��i�iρ#&eT���sP⽈�z�/ O2:�^o�!��cB�5���jo/��J'֚������٬�E@�;�I���UE
�(�r>ރк��*U@ō�+74IL�\V���f�� �r��,���yFQ��{���|�B�4����"��t����dv�Jx��BL㻧�̶��[ʈ�Q��kNb.�����eP��z��oD�0�P/#!l��/��5xz~��ڗE�,-�C��h̗��f����F�N6�k��~ņ.4W�ٰnU.2�z����t55�s��5���^l��W�m���85�;K�b~t���������ۦ����J�iN�eP��,�*�EV5`,�_Y�� (�ZJ�3%MOfR	p���~�4o����M����ܗ .5�T���d��*����F�뚙Hߞ� F�Y*.5IƾTm��>
��N�(�Ma����4��ߦlh�{G��_�FL��!�٪����4E��x%�T-��-`l!\��G<UsG�����E:�g4�� ̙j�"�|���=܃X� �X�ZƸ���.bjY',YNC�t?&sK�[*y��O��Eq-��u�h9�6Β��y~��<�a��dhk>j������nixh��ejX�Bq�����w7L�s��������^>4����߾\D����an�}��R�}&��
�4��ס�e�u�-����8m)Y�6+9�/�#���!��Հ�ی�VS��H����%��e��=#��C9ؖ��gU#�nVI�~�\5p������cU,��k��!6JJ`�Mo
4�_p!��� U��-�`ѫ
�׵a�.b�e��F7`.
���9O�MN����ul��T��v�_�gْ�U'�p	�Р�u���5��)�_�}=_�¢3�V���G���CV�+���IBD���1��������?��x�ܵ�2����0S����`a�LTJ�&���[�,��ټ/,X�4'^ֻ��n;�`�6���%x��j�1<���|�Nl8"�Q!�e>x Z�-��[�zAu�
��kT�w>�b�<s2�CL� �/�i��PG������}X~,�h�M�KX���K�Ѯ�DR���ؽ�٠�m�	�瀭��D`�S�L8�Qh�[��|�G*���o	����7��������ʱ��^B⎊�/�B���t �/df�ub��8Z>�L����o�&*{h�t�(@!�`R�o��&�G���0a�k2ci#7&�5����5�F|�h��<�7���9'�Q\��{]{D�3���J5�V��i:�̷z�#Yg)&?H����Z�x+("'���g����r��0���[�A&�t]}D�	֒¾�U�c��ђ�nۻm,�H�a<�49���M�S��-�@��<9t�h!^�5�D��x��}�d�z�i�(��Ux�Cz�S��h#�-X���_#0�S��tp.,F�ɭ$)k��c� ����}D���
p/��A#�I��g�ƍ���V���8y�qޞ�v���O�~��&�o`�N�|���x��s��a�N�`ɫ���i ��J�ʒX}f�]Ϯ�ǈ_Y8�l�p<"X��UM~�+N]���%��$t_!S�%�Lf'��f�=@]q-���^�5�p_���M'=�0��9Lu��EV��hȞ���h���+��oh�S�W`������A�Od/�!�f���j8"|����<;�Ȁ>�)��D�I6@̀� �7��<�iT�ٟ4�LLo�6���P���E� �����Q�NU���G�Øw�,��!�V�_�:U�z)y����"�`��7�<���_��n��Ռ���18�c3���nw�*$��eiⓤ<Q���y��p���q+���=`�	��rx���t'y���Za�D���Hj2��E�V
���6g����~3�9����C8�!�x�Oټ��nd�-U/Ηisf���7�PY��Ϫ����C�&�P��c��:�^r�����P̦�4�k�O�mg^a�}�������a�h�q4���q���Q�	$�`Q����\H{�y��rӆ��FMJ�bc6!)s&�f&gR	�R[��B�A�������8'z��T�SG3#�L���6��w�9�2y��̮��vn�+�bu��Xa.��
7Zv%�e��!@G�"GށTӱ����R�-��$vp���GE���E�]L�Ѡm���A��j��25fX;5.��:����0t�#���� Q vEgh(�������y��׋�����u�XGͫ�4�w�}�5��n"��C�4|E�i��2/E�]�?�z��R�'�g�D�~����0r&"b��\P9�ׂi����;!"4CJ�Ԉ+���~(VZs��s�)��@���6 �L�)z�T1tz#k��J㽨�\ߧy,R�V��Tu�=�9W��ǅ_Gl��w-��Âŏd�g1_9+��i�X/�|7�d ���ȟ�g����T�m455�$�b� .�VZi��)� ,U^��`��B_|8�����{P��\�}�'��	wAl��y(��,�g1ռ������|�א�_����+0,%��`�".��{)+$��~ARprک6Md�8nJ8��Z�����_�x�G�P(�-u��b
6�O+� ��usz��Ӑ<l�b%}w���rg|NQ�K���
����fwf"灨7Uo��H�_|��G�7�����kr�"�v�Mё�3V�;�l�"��l@(����\�.Aun���-V�\�d�����qUgg�a���@�{�7�x��� *O�ػ���$V?�^��`�>/ZG���$�@5 0�&�ݷwT�߈�.J,yZ�� J 0��y� �9��\�^e��R�������+��5�Kc���bT��T�"T&F��`v���vrgM���{��,��^Ӈ×v`N���9{�D�=�R���W��-�ڗx
#��c��x)M���܅A�Jk���!�D n��]�)f>H��lE!nphR�[,!��t՗yj��s�cf�b�.�9��O48�K�[����5f^���ˎf�᪌G�L`��j�t�&���v�ũ���ہ�IA��z���W8�O�pn�"����UE��#�>D�%g��\g'�~�=5pI�"Ъ2DU�Ғ��d1q�Q�����%_������P�����\����Tf�,�F��%t2���X�\i��:0/�7�)X�I�����Z���^ˌ=�qB�o���}}0�у�+̔p��X�V^bjԃ8�tc3;�.�&�3��(i�HEV�S��]B�`��� �G����Jg�h�
��&��B�����X<�PO����Go�cOD�]��(�hF�G��--)���)�_�Y5���/�p{��~e� ��R+5�>V;_�#V�����'ƳI?�y�__�D���5g��,���<4c���Ph�K9 HI�2�@�5��� E�K��!�q���2��٠���%�J�GK��aNh�>�`%t���5lqH|�͡W3��o�7�ݡ�*��k9DG����P:��-����utH�&����P���NG���!t�5[�t�%v�&>w�J'� w�丄�	�EfӺ���F���&�:L$�bs�)����+L���v���{��+�����i�b@���\蝤Wd�X�b�yU�3�o�U�d)v庱�@��`{��7=<���x�3%|m�t`��	��ݝuM ����j�@��F�E�(4w�m�YO烗�ۀ�W݂E�Ic�%GwW�<luB�Y�d�O��/a�@����_�&\z�M5��e�U�1����{�Y L�UA�9&'���� C��Կ
<U����R�i�Х+�8~���%y����b�����\I8�JX�7L%t��P�qPh�>��Q��A+y4?���-�vY=w$�pdѽA�Lf��e��w��3�^[�8�>�����Y��N�6��0r=\��`:�O;]�^U��IO�(���������v����AQO<1��f<9��M�̌��E�Y�Ǟ\ζD:�Z�S~�0��x���cAfl6`$0��k6az��\�AO\�����E3"��U�2���[[-F��:#�C��c�pt�*�c`�±�1�dMQZ`�N�v{���Ղ�Z�������[|��չE�V	�Pʚxq�G����a�Ylp��~��r2�vdzk���Ib{�u����]D]����8fN�����U��ʒir�O��g�^�������w��u����y����� P*߸��Q��RB��y�Ⲛ��Ԗ~�r �������W �`����@)kex�b��!� ��-��FSM�QT��m�'JL����T܌�$O�u��'����)PY3z��P�Et���\C"+uʃ�vT����Oԅ�ӢO�z�r�8�<6����^�~�(!,�-o�6%�ѯ8���)�'����,`�/ET��G3����H4�$�������.�� Q��A�_ր�8'���ozcN=�H6��1�-�`a���)�*�VKz�����À/K�0�s�	�i;�>n;gj.Ro�>~"��꧓��W�Ld�|y�Ӓ���9*R��!i��C~Ku��Sz93�KZ�����x�E��w\F!%��| :�ks~띀P��u����k�Ym��tk�8�����;: �C˪m�.#��α(��η�h�X�.�!S�o�U��� 3�p�%�8��@��R���&BξV n�u����Q�V$���'@��9�j_:gi.c����N�X�NƓ���r���m`v2�� ��Y5O��x6
�ﾙ�ǃ,���eE<�����qA$�j����Q1@C[�Rv�	t P�/ l�[B	'���]��|_qa����8S�z*��������p�|�M��C_�Џ��Y97n�H<�1�K�!�1�I��w�Q���7'�����Dz��vd�RB�UsI�/9�3��;.fu���M���3T�EB�7?�/� "�Vs��Cb�	���50��1�;����k��*mt,�p��hI�������	C��7gO"�:�lQ<k<E����"�t^�+�e&�֯�M@Oe|�?=
4�@I��Ϳ�!�t$]����&��^k$RI.��'t��!!�l���
K� J�Pe1NU1�%��.�[�Ꞃ���[�ϏD?�_�� e�[*��_�#�8z�9��Z����_�|���65�%$�� T���Q�[{�IO��-���P�~I0]�Y�QT��ꆽ�hr�x�F���{)5�WY��̩p@4t������D�� >�|��[�"yЏ�
�7ؽ����+ҩX�O,����]�s���&IUDG����T'��ma���6��D�-�Gͧ21��g�Rχ�i{ej\�:��ڴV=���L*����߭g<p*9:V�~��2@|�"]s��B��9ѦςDd�ʜ�kV}z����Ҩ)��k���+�3'��=sWt��C�ƹD�E	������o���`?��oQ�[�7�Y���c�j���T\X�?�I)���R� Rl���>vMz�2J�S0R�d�,η.�mA�}�_��K.�dqhKe���3nڌ?�4m�?����Ьqެ~��I�=��M�u�Խ�����l�l��طݙ��M%��rl�����d��r�Kd�&K�bؙ���XVr���I+���-�/��D�DɚX�I~c��QڭՃ�WCuir��թ*\��&5��D�����u����|-�� vKCM{(���Z�� �*�H��f�=�=��5��K���FY��x��vFL�J$��j��~abS"x�>&��x��G���G񹨧������\�΃R+)hAJ	�&(\>�?�e)�9k�Z�
jn�/E��b�p/]�N`S6����[B�@�>����W��������!i�Gx��ƈ�$�:,ki|)ު�Ft�V�#��⛧��l ���k,�	��,a���2�;�u^/�Y�� �;,�jT�f.�:^�3���D]8�N����m�B���ڻ��>���'�x���,\��c6L����^���Hq�ٓi4���<3J
��/7�_d��o�����\�!ΏǱ��@�}Tq��ץ�s��V�v~,�K��B��5�g ��ԷTy#�����ϸ�`�W<�t��E�Sn�fqSK������˿M�-��$=e����!fB��j2��f�>�[��	���U�(;�I���pT�}��AL���r����Z�崋�#5��2��ͤ��>��H-ｚD�k���`-c�(�\�b�ћ�����i�@×��+\s����&����v�M`?��0�#(��Z�?�Gb�|�VL� jI2RzT4$҇�$EW�a���X���BnE|���ad��a��"}�n6{-;L���cC� �@�;�i�>hS�L��[�-���+�[��4��/{H����m-�e�c#���+S*��6ݪ�i�d��I���~3`���y��T�߸Ej+��_��Y[��c�����;%Y4�"KG>t1[�� �j9�Kf���P]2qv�UDRFU7�%��EA��)ŕ���A���Q�������������o�h��\rLܮ�	/�<�'Q�7���J���C}�$Y�~��-�?GUi�����܊�Y0	�s����10����e��@r�����g-�B#�� 6��6Ɗ�x�Z"/��abٰrl{^���"�`6w,F.��(4o K�UG�D��O:���Ԙ�' h�0F�� ��6c�j@gDќ�r]��S���|9�G�#�\�G�f�e����iI�^��'�� G����5���R��Y�0Ȳ]���{w'�f�?G���=_T���2�S����Ģ�e@���#��Ǔ5�u��Ϭ�c�i�zc�,��/���;px!�X�W��b��/�FR�΀!�8�AC�N2���K���~�K)�.s</�x29 �T.{p����z���# a,�@.��M�D1�0z���	�!چMV�7��ղp$���b���TE���^m�W�3ˎ����p�,0F�D�B�7
t��S�L����ߐ����0js���$V'h��Y��XC5C*��#�����pĹD�V�Or��ā��|�:M�b��0#���%zp,�<5�����t������3�+�8E�sC��rOi8��C�d�_Mͬ��B�گ@�]�������]���b �yK��:��ce��E2�ȩo�o-E)^��B��OC@�`[��t�n�_����8"�'��\��>����y��+kӠ[B	������%_9� 7�x�L�j�����WJ�!:��R�5G���*����ר��b�!�s�f�g��v�[���e�%�3������z�fs,�P�32i�7��2��{39�}��`��08t���iذ�p&����~I�����9��<�S&��㩋��"m2�����|Ey}��v+zЭ���,Ƕ�Æ��e=0���oW�/k56��?Ҏ���'o�������
#E���w|S�� �[c�põ��R��tl�2S������C���C�%Q�6��o��P��,�n:&�`\�#���h�
0f��Hy�,�oL�;���h�4W�ŝ��q��Lk�[�;�S�!�������]Sz������n�����S�v�W;ǯ�^ �6��~֏?���B�e�A"���Ei"f��)lQ
�_�N�,d��åAm@��@DK��Td֕*^��&`o/�v�n�Eq�rͭy�C��)R�Eu�ڌQ�1�,-h���n��?d_1jc�m]4.�z�~럭�'�d��X]0��]-�L5y�����Z4|�M�f����X�H������ j��A���
ۀ���Lk�K+���0}���Ɍ+g���������}���jM
��;E���-�a�w6�}a��QQn_�S����EUdН�_� �Ŷ&�.��a�L��'���������[��;�"%+Έ���V����v-9��[Э�/F5��	���А6����Q�D��w ��R��<.`:�)�tj�J�ۅ�'�(�j�Ǽ��Q��z�ް��������8�ާy�kP~�zg�A%S�r9�VX��K��JF�EZ��������D+�-"y���Eݔ���
����1v���z�m�yP��4f���	s�X���o�*z�i���aο�?�p{e�0���R�2{S'�<�c��g�v���C�؟WPX�hcv<��V$�V�!W����o��X ��Ft���'�A���!����������l�3�-��OIm���d��Ym�r�W���d��[�܇�e���)׉��_�-^�x��7Sӷ:2w����l�NfA�!{�{^l��:t�#��v=�K�{���ؼ�Ӟ	�]���ٶNb+`��/���$��Ω}@0Q8�z9������a����W�'�X��˭���,�)@��kU����k2�[�o�n��Β ���Wޱ
�ޑ� w�7s>��c�(�tI�
�Q]�քz+&w�z��O�g�-�t�=�ܴ(�Ǡ�哦��k�<�н�W���Xf#����\*˝\S$3l�N��=0��<��$*���T�g�D:Ac4%�4o
%��+Ʊ3D��1 0���K���u0Um=?�n�G�%n�}
Ry���Q��x�1�X�#wT��ӱ�k�*�(V̮�QZw[�wZ��![,z6����tʃf$ߣ�|���J��[6pôT��A���Z c�8�A�>����y�����8��k�o��יR�����?,gVM��Q-$K�-gN�H7���$�̍_��K��{O�Ҹ�U n� �m��Km7G*|i�ol+�Zwbkπ �
f`Hh�)t��'���g=yխθ��B�*�85)D�W*ah���
Dx+GU�x�_�pH�G�+��M�g�1�C��	�MR��V��?���>�P^�J3+e&̔�y.^gS���D���!�X�9N�4q�]ʹ��HI�0�'�z�����Q􍐴�$/����~Ղ��ެ���َ������<�ݶK�uPls�4P���^_���<C�4�e�gʊN4"�ro�g�6:�y��-�۪���!m/�<��S�h�\���$l���b�Q��,$����$b����|�q=�I$�\�ȷA�1�c�N��4�As�5�&
e��"�0�?G���t�U�?(e^6���SVZ<e��^�_s�ߩ��r�UNC�U������1!�*�Vg��s!�O�<ї�!���|Ĝ-�Țˮ1��55�q���7���� {�5���+�q- c�b7�Pp>cjYx�v�-�2sƳ�?@���j����H�<�cƄ��Q��NC^�����:*�����7��9�Ș�#����E(B��q��
�)n���tVV/s��y�����f]'E��޻��ڊRP�a* l�!�@n��U3.���0�x9� q�z�EC;'	��|k��1ï�>�z����v@�M�)�<�@����q��CU��m�g�{`�J&���^4z������`Mz�Z��jw,������U���R�P��e�]�F���Aϔ[b��4�"�lμ�	<+]�.�Wʉ,��4#6]�

)s��Bm'���W���;� w�H���K��|��&ne�@��
��H5���̓)���~�Xb�Ft�FFU(��������}/F�Q%���/C���<x^}��)��jW�F<C�����#���V�~�e�tn���[Y
c�0��:��W�SE֮š�P��~�ޓtN9���F9	_�}A- ��@`*<�*�` �x�[��+�GJ�\�ۆ%+Ĕ�SS��n��v�lV�r� �h��`v?|*n���ޗ+�!��raun�����V��m� ��`�:]'�>Xϼ��3�P��y��I��ezh��2H��i�"m��u��ܟjx�	����m���a���iX��텿|6�N�$��p٩
�7f|���.����L3 ��$�n'
��d�N��k���x�h�+܏�[�	��� {A10w	5�Ix!�S.f�Y)�N�R�^�D���n]x���f�������ygf�C�Y��0Y9.Qk���kq��ä9�(� �����]f�u����"5g�y�u�4P�����Q8���Tf4�3ĕj+"�[1��UY�����kC�e�sb27���p��tO2��t/�bsPK�w���2���$��\���8r��cq�M�,,��y3U�j�Q��(�(SJ�%�R�������9t�;��L�u��������c2a�-�/�~�/�}Ѷ'��� o����X�[�`ܓN�Ȟ��$yD
A���b�$��:*Y�p%+���˭�N����K]P!����5^�pD�o�p�6�-qY �;���wL=t`;�o�1I�ي T�9��ZЋ�v�z3�Ȝ h�o��ɏ������%d��HL�J�����A���ШO|�U*r)k]������߀j����0�n�ވ
��bZx�*�{zJE;�8�|��_��q�#��u`�H`b���;�7�b��!z���4��Q������rr=�Z���W�7�˒�dD������L����p���*<��#�����C��֣s�?n���S3�I��RoQCQ ��N^�]�4���b�z�ߠ��VS�m�n�j�lqI�d��4ܴT�S��ƆO�R��b����TՉ��\L�=�v���|\��q���w�����>x���Z���
�j)�Q�e���k;դZz��uu��t*��N�H�J*q��9�c(QM�>d]1w~����^x���2s���w����]� ������?Ո�P´G^b5�`Xz�fUI����k���e1�3�Y��z�)q�}V`�CHY�j\M��♄s؄\^���N|�=L��j�ög8�)�W�+O3W%wF"j�{oz3)��.���҇6����.�^��0����Y�a�{=?�3�s�*r|�!u5+�{�'�"V4��ơ�
tլ�1!�O3�y�*S/?����6�q�7l�1���\߈�F��F<g_@f�x� �&>ˣ|�c�B0ⰾW��w��yi9�r�}{���������<y1<"�*t#���;ԫl<j��Tn���_�QO����ZDċ�Ǜ$�W��lI�TW�{�/��!09[��6��Z2�������'k�y�j��-ĭG�|6#,*o�xe�@�~?�=�V���3@����ܦ����h�s(�}��	�ڼC9>�����:���:�&�h�ϖ��s�"��&�4�d��8N$� ���N͂�DܬI�a�K�A�U}#����:%,!�Sa�g���Ҩ~b�s�D�ӈ~�d�+��Y�t��Q���w��t���'�^��"�dU[9�!�ԟ�H�e��.!�#q��@l������{
p�M���x�V����H�K�> �9t��f/����S硂�V[*��ID��]R�������+�>���>�u���l~}ׅrB�˧a0���+�e�K�_�u���e\�0c��c��Ί+Ac��/�3%2@xw*m��T��U�v�]1��M[�,\�9�� Dh��I�m��P��w��G�ؒ�۟���1$�
9��J�w?��dr�`�Z��AFJD�`�m�)�/��CW%�]�;EmO�c�&zDk���i�d�Ռ�}�9=��ڨI�Q��2����@8o���Oc %>4��.F�C[r#׌0{�uT�1x�(�/oO&R�{��fL!�.�O�"�'- V��f�b��|�w���+����t �C$J/	�`�I�(�!0�۠���'H��'�rX�Mo}�՛��_�p()���_�+�Ż�i &��|�l�T����/x6�Tp��)����E��m�e���K�4���Gm?AM�2�V36e�X>n� _ua�[#�Z�5O�~:��
F���,�Ë*;L*���O��X,��F�(HF��d�# ��9r����qQW�$c��cW�2O�Э��<<%�O�ǳ4�Z��#���x��7�V��֓>�H�J>-�;�'�$�&�O�ᒑ/WS]O�9R��H���t<?E��>	�V:y�iH7$�S�6�������L�B5��f<!�}k��Z�t8y�ރ�-����Fà�r��#�Ѐ�N"��2ܟOH�i��Hf��Ⲅ����R$�h�l��%�!�b��I��E�r�=]���6�]\lJ�������P|�.Ac���EZȏ�M� ,���2A�n&�*���7��������!��F$3o-z����X:ȏ�R��%�*��]
��M:��$)�}咆"
bn�u��*��#F~�6��*jN���M�H��v���P'9'��G����0�=vx=�'D�M�\�t)�0Q�#��S!F�J,�$��ۦe#
� x�`WN\a��Vo�T�K�Q�%��5�J����N�]��8/3>�����0���̆��.�@��n��KL���L�;�-(��(*/�i�x����z��F5�n��f�X߯P�-�輨a/���Q�j����v�e�E�凨_�E��6�EI
����Jx�eE���I����I?	�G��Iܡ),a�R:�q�L{g����9�;j�8��~V,0��yn�xաf$Ke"X%�V���pҠVbj�����j-f�mk���R��׀��.�����O�zd-п�\�ٌr9�B6�c��D���6"FD�$q��CHo�%�'M�� 4��$�*���p^�!�9i�G��<��G�/2��<UI��p+Z����
��1$��U�D�7���o+
Z�1�� \���fe��?c"1GA�eK(��[P� �B�=_g�F���n@n�K�ٳuL���l���h}ߖg~,��o��x�$�%Ŵ1^̈���d[\7�i�Ƥ�4�ݏ|c�w ��?��s�Ud�EzH�t��țW?������F]���j(p~�T+�".���
�'l�@V��G:`�����2�Z�1�?Ub�O�J��m� �+�� �F�{�(��5�Bfȍ���.0h7��<-�w���%e @����{�6N�$.��w�@����|6Mp	��y�-�{�2�#�X7��f<SXR�8��<a���A��A΅#=�طgU-U�����9��7z<�R���ȹ�¸�\�TY�Β��z`|�6�@�Q@wb�&�z��0;JG�n!�Z�x�p�	�n��LG��ܯ�����U.�|�*!G���� Xbb�(<K�}I��GѠ���o��ݫq�Z���dƈ�bs��@D5�p3��'��I�o{U���ОW�@攰�S�2� S/S�Y�ی��5옛�i��b�I�Xt�,ĪVI/\ʹV9�"l]����\���\��t��㕗������|V�go{9�}a���I��w�/[����%��I�V \T�
����@��J~���X{vM������v�\���Ն�����oa�u*��'���k{Y	,SU��	E�����қr���Ӷ�]{FW���f�p�k�T˂c��L���57����!<��˘�w��`����P�=�/M?i��he5�]e�t��ov�*���@���|��g\�2���^��ă�*�Qu<�����RU��' ��@ ��Z�|P̤��C�j/�w%�/3�Dnq4���BA�T=v�ߞ��]��M��M��9=I�t��Pb%z5�7�SS���������^V�^<��6�Pp7?��k��FRď4��g�_4�ݗo<�E�Ϸ�Y�Lku:�'Lf��Z'7[�$����f���}���H�s0{9���;��lP�F6����jn�Ͱ���IK��L���~�#)��S���>��1�gY��3�eu����;������>����C3���:�r"�3��6T�#a��#c���q�g2��˫7	��ԓ�v4��U�zKO]���\,�0J/�<I�M�>X��MO]�C��|�&$�yvR�Ow2����0I�$h��.Xf���!�B �'/��2�?�"l��+E�����������^�Gm�'�'���йC��z��pj}��l�8X�.{TҪ��h��a'*�اj�K�r�`��g�؅���oQ�R:���M-���w�s���\*cU��8�� ?���v�'�,I&Z��:�)�X ~��n�CUm��� ��~;�.7��(1�z��lsף��"��n4�Kj�pa�$ u�n���,�K�3i�"�wL�a\s�pP��K��V��A��h��:��jܙNj�n ����.��]c���]po���g7����k��(2Lc�N��T��
�"d��|V,�g|�PN�B�����P��w=A��*n�Z��r��Wf���8�:ҡ��"J�8�S��ޭ�L�uЪ�T���vYGuE�}+�VBG&�<���� J����T�����0�(��B&:F��F�)E44z�	H~-��~U~'�B�CN���-��"\�Y�/��Ø��N�Q�G��	v.��0Kݕ�U�k��%�.#za#ϖc`<p�wO�����\x���~[�_ �W|�Bw �{�|�8�=TunoV�0x��7�;=���(D�GWma�'�U�qB�'�{B쀠߶^�����k������g(��3�B .8��Z0uv���tq��T����2��r.:~)ێ�"j?/���s-�~�ذ�(����_bX�1
DM���D.���	�g���B"����n��o�� v�z�>����~jpU���0������$���O��J���9ԒO��'E7�=�v��:�@'8�9r9��EЊ���_�b �]�(��-K�w��Ap�L@,�.��5
Ԇc�i����Z��K���!���"%����?O�"یsun��iA)E֥Ck����w$������l�?9��r�	2��u�gծ�罦~�V��\*��Emȸ�����R���iQn_=."����-Lr���X�ͧg�{9��:쾡��(�'�8�b0�Vэv5�i��k���p��O�Xdr��qs��v&:51���j�9�#ߟ�c@Kyf:g��p������h�8t.��뻖���P�˦ǃW�ቊ�L5�ɑW1M=jB�����ɆN�@��D�K�p;���Ue�*�]<3o`��vZ[Id-���wjf5�q��b�־%cdP.�+(�ó��<���J﷿?%����h�ő%����5X,7h���AH+Cʟ��#�]e�+t:"a~3�i��!K�f�v��v%-���I�m��x@h��I�q�U(iF���Ï�կ��^\�.�1���
I֊'�CA�G�{�
A_�5�2U˞�#l��n���M���m臾�f���'�Q�"��aٕk�oC�{��</~�R�Z� d���(X��綊8��616A�͑�Ok7a�������˺���#�[��l�'cY5J3���\�2�M���(i~��K�O�n��R��z�f�3H�/�q/]k��y��ݿ���$��O�I��ZD�Cz>�l���O�����`E��؄�X<k
 �J퐓�J��sXy/E����ߙZ�{�Ĺ?������@p�+v�#�~ބ�~�ɛ����֐�h͝!~���9r�@i��'�x��\� �bV��Ul�:r���~�>��_�8MVM۰ͬ��³���sb����J��;�~0�Ԗ�#6ˋ`�^��Y}HN�f���]+Օi�.���UڊI`p��=���PPq�e!86�e����|`=�d��㺩���y,����;6��&�l{!��QQJ��vk={۠쫃�4b��b�����J��˟��w�TRw3ܜо9{�_[ֲ�	S	��$߃���A���;�MG��0�h�˥���l�4�{�^�K�7m-��.�X��%�CҀ3t-*���ۺ�hF�x�H��B��˞2�t �k��i�x����}�sO+라��A�y���G�N�E*?�&�K4�̙|�������cJ�z<'0m�[�㫅�]��T�p�O���z븳D���4U+�A�U�J��@�)vp4K��2�fo�Ys7��v�oQ
�8��w��n�x/��N���t�a?Zzr%#Y�uؒ+�y[xn���	����D�ag(�	/v/��]z���|ɛ��Ҵv��c������e�&?.�6���cv� 0�7��ĝ_!)T��ʊ�.-��<Y���L�d2@C6��sş�и�u1�1�a�E��C
���SnHl�N��=��S
y��Jȓ�FzpH�Rz5�C?k�;G�����N�V!!�RRG]Hx��EF�B�����:��%�u��D^ [��Аwi�{Ym˙�4�V��o�Ln�l	�A�B�������T��"�-L`��5df��W��hW��1��ݭ���@�(`����mQw��`"]�q.�gGo�y�#��rc�e�M�4F_�u�[JI,�R[)��i�)C�NGyTUns��A�������%v
��]ޫ��k��5�3�v�\�=@�?��6�
�[��K|�cI���@�.�#OZ����dӟ�)g�KD���0L;ѣô�7Ъ�uQBq������@��D0I�_<��ɥ'��䍚h&�2SJ�屒�|�]��2��4�2������Xh�J��Ph�)��fyaq�d�v����2<,>�!��Su�S��o�'��V�y���q%'�ө����F�=~�)t�'�h1
5�B���U��+d�п�~�"~�M�]��O$�^��F��3�Oqҁ:u���)�xRi{>�B�IC*lhm��C��>.���-D��UB[�F6n�TXQ>��'��C�/�	��w�\y���-�l�ވw^Px�nȱ�wipWrMqh�Q���_u� ����B��{AN���)��w7�4���A�蓘�������̳G:n�6�g�hQ7Ds����T��� ��[��E���U���yj}�<��9��������+]]�e��*jD�Q��n;|�����1n=��X,��U�� ԯ�����l@~L�A /���!�v����'r��-����>�x���,�d�w�0�-)�%��o���E�(?x���[�c����[Md_n�B�S�o�a;��8p5D����Ӿn�C�ϙ���N=.~ֺ��+|� �>!!s�_&�y"xW�M��_��Ck�%�_���}_���6�J��1.��3���b$xu�a��k%<�V A�z����v�^�Y[�{��c�=����|g)�Ai�5�˛i+�)�^yH�OIc��'�ca��7�N �^�oRzLB'��b�][K8�V�ķ2a�d�*:6��Z_�UQ�����T+{6d����C��@��O�8=v ����FJ�m�r|B���� 8W_�b]��T�����g����Ԓ�Cg��@h�����f��R���y��D���3Mƾ��4�n&<�J��+IŏŹ����8��&�B�h��L���x��TM��G}�����,�)��Rz�D�(V��������:;�0�V��I �j��%�#kgQ0ޭ�(x�L����\���]쒮bu��Y��8��T����?��*1�)�� nǢ
��&�@��JbS*�9v1$MZ�l oiq<��p�V��XD`M:�R��w:t��ŏ�S��6�E��L��T������Y� �4d��c���.�Y]�MI�N���Fu-��� ��.o?�,��Tw���;������:�I��L�B����g��qG&��	r�}˯�x�1�Q�w���0�{~�ΰO�NE�aVٴ�^lWh���O|[`� ��h̝{��e	�Ѽd:J��j_PC�+<���aS�%�ܐ7��GD��;�?,0A��l��7B���A�w�u1>��;w����9Xp�+�� !.��7"��x�N�%x�E�g�����rb�knEΧI�Y��r���1��������?�v�?1Xn�y	/�g=�%�5mD���D?A�0��_��)TAZ�-�8�B�#z�6��8�(I�*��3Pr�T��T�6����
p0����e�f�*�=I�f+r�3�?�'|�!T�Ƿ���ǳ�9�=+�B�����5�6}��s�W
0("���Z.�?^�˂~V�iuU�q�r��l��X�`ZT�Ә����-����Y��F3����'3�: ��!��J	���{���(���C1�������.p�}}u?)������:�F���h�u[p�y+�6�ҧȏ������=|XcF)AU�]���{�";�Xb�xX����W��;-Y�	��/,����wI�Vbd�`l������!�ދ�u�U2�Ij�)Y���v�x&�s#��LZ��6T��?ʵX7'�M~���,������'F�� ��ʸ����Z�SJ����=�Mes�7����y-���*�h�hl[0D�1�!򮫆U�2���:�����b�$lL����ߥ��2č�d�p�m���FvR]�����.?�*���\���(",��*��%#"0���dS>Lѻ��=���e[O<�s�M���gm{ԧo/�C.� oj
�v�"�D�1��qד��;?��lߡe�"s�eyT����4y�v�0��sQ-�[���'�U2Xv�G�i��>����4�8��S���V`}����}��/%�sfH��O<�����G�N��ҳAC��`���:�,:�Q�O�t{�X5nP�5�������Qg�1Sw�v��tV�뻑h�K��0G�$DG÷��bP��Z�����˴ZP�5�NR��.m�m�"��\��1�6�Ҝ�[�M��vy>,Y85�Y��^ �-_M�m����:qe5���$i�~��\:8׾����-�MZ��P����o��Y�[����S�f)D�8��~�ql��|���)�tn<����3��4������E�Yq��hL����t�j�&J���0��_��\�R��RW,#�s��?�I���T�ξ�1p��&��?��L���^�����D	�S�����G�0á���g��y@S�JUQ�8�/������R�	pv �A<^��b��t6~,F���W�����u�Y��	X�3�/ǞJ��b��|X�*f���C�6�/�?��q�v�0�?��n��<B��W��	,�^���\�XP ��3	��S�B:Q�	|k�H���&��h/��&!;�G7uV�M�R�h��ķÝ��ŝ�qq 8��G�����]d�(�?KD���A<w��]M-�.�U"���9�smeu����>��gQ�;�M�%U�8��b�iL*ܿp��1����vU��h�6�&`<B>M���cf�`�rgsRA<%B/��)�xK$���t�wG�iV.��vA�CW�p��)D�1)&�9-��B�uUV"K�,@�#��$^�K |�W��vN��-h��|	����y�ppWy�ҕ�9-P��e���j�\�Z0ILp�3j��D���=��'_H�hÑ�᱔�rA�Q�4	h�s�L�,K�mΝQ�&�N�޷�����N-Bha�ַC�Ɩ�?��8m�- %��x�eI˽��r1w�I5��W �ECh�~p܅�dt8ᣀ��P3�,o�I�"s묶]��8�.�M�4g���}�2V�ʊlr��Kd�������P|<WB*Y:ט�٬l���a�ԫ �34��cZL��b�2�ߟ�Dؔ�]�W]����ΐ��@�\φQ]�%+Z����^V�@�81E�j�Э�J�Z%J�LE��+�!}�����ak3'{@m��������2F�*��OB��V]�Ƹ�y�
�<�\��P`3]�HUk�/��P���|x�7�B��|쭥��O��z��|���)�Bܑ�����e�pX���x|��;��o/���8��G�-���V�:𾤎�TI	f�RSy�]Qx���M��0l�wx3����ϫ�
��+�f�D�U�<������樛��5�Wo���I��a������Х�WTw��y��,s7������Y௲ơ�Z����%�Ha��d�P-�c��i���R�hke�7���� �"���o�����R�;1��Z5��kQ݀7�R7��^��:����d��x�F�{��5*�������D����(B����5�T{����ؑU�o]<��ej��w�%�rmR�����嵊:�5��[�P����������vFh�z�P�8s�Yu�nT3d����=��V�c�lLKГ�y�c�Ya��#��=#������p��,æp�P����gT�6m�4y��I?"��R�ig�yYy����Q׋c�D2�^��40�Ʌpu�HdC�Aф!5�ƆL���pW�\�YW7�o���h�EØ�u^}��>��G�����aw�p��`�Oe�B뢕���,QR�0����*��f-��Bбopj ~��I�=S�M�̄6O�lb����]8(I����vG@8y|��x�t�?�y���Meq�)�];�������^g4���:ib.���x�Y�0R�!���ǐ�불���A��H�6դ<%I��/.5�>���|]Q?���*��x��MX\4xn[�_�ig@wԂ�Z�4�	��O�G�ҩx4�gT��ȁ�e���9"�\�`%U1�z�"�fXm=O��@¢�q�VP�W�1�,S��	;4�C���e5��w*�c���g`�&:�8��Z;à�lq"k����֨ǚ�ڵ��YhxD���d��W�b�</+۾s�3K�ըZQ�鎜�����m���-��puDG�*�Ӻ�����pE�v�����&�>���p���7��Ӧ�@��M7�8 ��?K��&R�� �_�)�#`+�?�=&����Cˬ��JJ�|:�MD�\�ܒR#����V��~�Ƙ /�Y��?�ҧ1�jw��JJst��H�6�TNh����i)����d`�}s��_��ux��z����%�p�vA̦��Kl1)5�?��J΀o�fj�ZK��)�ǃʀLBy�E���c�v�//������;j��LD�S�/�����Z;8�X�T�K=���z=H�_jb�xH�]h�c����չ�(�;c�[���l,-������/{
f]�{˃�it���V�1���Ƥ7U��h�6#8D�N�l��H�~5�Iq7�ߋ���+�O��tX������S#���N��*|���B���Y�O|�'}D�,|��(\3(Hd��s�~�.�DD°g�P3ϵ!��ɲp0�Z��ŕ���z�
/\x�g�������r�^��b�塰�Uj��������φBq����v�&;����i&"�0��	9������[�s*�ϩ�7Újn�.<�/<y�_eҩ-�3b}�)��v�֌5�)�����0Pv &��X8 �rU��C��RO'�D������_o=�(�GNHmM�~x���g�`�SRfej@�1tʥ�T�)�0Ν)Pܵm�-w;!��l/Ƿ4�Uc�%�LޣK�ݧ��HU�?2�P}k��B�rA|
�uE\p��T ��G`��;���Ծ��(Y��h���1۶���+�	�ǂlny����%�	M�n�u�g˳�si�m���Qמ��B�7&��iD�o=a�2Ĳ�8�����ޝ'��5��Ǵ.Mcy%����k~_�jۜ*Aj��*�']"������*#R�P	_�s���p  %��AVv�X7J�B���0e[W�[��w�K0!7S)>!7!3OF�H��Z�4���%`���S��^�����R�8%$?X��9c+y�)�ٸ����1�h�^V�_�M�Y��#���4��7i~#2�o���aw����=Sb�D�V�5�f�H�^����s��ͅѱ퍬�*�~ji4Q_X�
a ۾���^�������`�R�(:D��>�O�PL�����p���8ǟ�eO9����jj�>� ]�@|ͩӇt-t�:1�]�㩝�#�s@����%���ʓ1 ����S�[�Ρj)�T��b���*�K��U�?��&U])t�Wa��+�W�����xΑ�íV}Y,�s{�u�Ҟ|���"ĩ*.�$,'tY<�,n�6O���!L�H�'�끔�����N-k�BD�����"	�
� �ջ[����U�<�?�)�� 8:�ؾ����3�.���d��+�j�>�S���g�B�s����8��H!%y�p��Vb('[>�Oj���]<1YS}�z��0�|i/Z�i?����q��^-hH��w�:/B����߁2�f�U.3&�4��8�]�YHŉ�hʓ�xC�\�ń��:�͇��k�D� �I��Q� �4�J"-ܫp�V3YBөG6٘@ ��?��5��B�� �	r��nք[q_{x�x�N��,���̵��'�i�`�wu>��ʥr�l'�t{�@�>'�RDd��16����I��ԝ�s�%�䘩�(L;�-Q)����i�=����eU���Ӂ�R|��<���IK�|�K�^k���\}����eY��\0i����cBh��y_D��%��J�NJq�&ɔ��l�1U��aʊ��cBѴ/+�eQ�pJ\be��=�[�ʝk9�+&<��Ɵ"0���P�9j�O���n�E?�*�Xt@����,+,����?Ï����C���X��t�R�`���fP�h]�b�F�"�!|�����j�;���x��jeR��K�Z7+�H#c',-H}Z�C����'e��@��S��f6�������B��jG�NT�+���l5�˧�t�������0��N��!s���*m��	E��2���\Mm�J��$H��L�9_yڧ�(\hB=�'�Ϩ��0��1�m��( 1Y���(�C��~�悷��3�J�J֌�D�o���k\鹓��#L����S-�Š���ؙ5jIο,�Uȍ�l��F/�nDy��a��m%"'�N����,D�dV��W���ʛ/r����?�������u���*U��	g��3�����ն}C�Ā�K@A+�,�������c	Be;ɻt���-�|o�R����~� �?fm��s}|t��G��p��iC�̥���1b�~�["r!�@f�
�O<e�8:e��Za�76����A#��u~��6��ݦi8��^X�	|٩��L`�!ǅ�sҢ���^� ���I�-���NK�I�3��Ż�s�@�S@���8��R�0RVY��n�x{Q���t}����o��-�Jz�j^0n_X�U����á{�Y;� ��MCtPn3_g}��Wpސb1z�����xs+˞���VZe�M�����f�M9@^�G$D��v`
�r��b}�� �V��ѽ��6������I��,|H��ifIߟ{6?���^A'��R�#F�5�I���� �S�iQ����8�3HU����H�&�����,,�Q�
!:A\�P	5A)ɺ8����m%�>M	�̞?l���;�+����X_�C0����?�8��jDE� �a��j�(r5��Lqk��aK��:<�_���m�JYך������9��b`"�Xk�0J)����������Ua%S�F�&�0X�;�Y����5sa�"�������xw.�u�?G�����'�R����٪]��ȁX)��V\a:�"�0[QC�|�R��*U�#��1f�-�T�R^M�90X������7[�4��f�%;t��r5�=s��:��/`�ڊ���^�x�ʶ��t��h��˘¨�@�ݢ��f3�.����O;���*e�xu�a�������+�AE���D"
F�^j�w~l�z��0�fF���L��e2��D��\:v���CEZF�O]�ӵ���]s����y�v#.��|��9�Ƹ�!�����>�t�����	�� ��uKD���Wn&êߥw��U��K����Es6l��*�[�o���7 QP�0���Z��U����pl��U5�T)@�Ϊ��I���4iϺ�I�i{�~�8���k&7���kt-�Ȉ	��?'������>cf^(�c�rD�	��3�����/+?(�ݢi���ݮ�s�Q�9h�Y�kO�=���I3�*���9.�`L����Y�@���$�r���!j���Wm�k���P��ׯ5���	;��V�b3��y�K �X�G�1(�_|�n_�w6L�f��9n��BW��4i�Ձ	�Dv�].@��=n\q��S�Q˪z_��p����ND�ʸ'�����<�"`�"
�u��u!�+3B��jA��G4�j��H�Q���?1�Ao�����	^a��V,�r��wn�@�U�e-�3&�5q{Mu��]�G~�o�����2�	ī�}��j؇{)�X��F
y�J�����pfS 
^-��k� Pt�
P9��z�[�9���YC�����li����Iv�9�����x����գ�9�i�S���Z���OA��܆��������V�l��MG�J��$:C�����>��$��	c/�+;m��h�L����q�(,;F�T3�hM,���xa8��WL�b�]]�6ͫd�v?��6q��LL?�_��c�klr+n���:������'��_�W�쏫H��E(ų�/�bm�/C�O��c	a�8�(I1���~�t��q$�TSWy;��Þf��zLS�F��R|��]d�S�F������2�,!�D�0�)(؄�\y21Mu���ae�N��HE�6���"Ղ��i�t�n� i�L����p��6�=�;Xs�d�UL�U6S=�ý:�
^�SӘ�a8]�������hG�wR+X{��|u���d�}a��X�TFj>4d��	'�K�HW&��E�G�/[/� s�I�;�_5G�^̟�����������6ڀ.����zt�:�ʬ���F��ɺ���%`;���(��&;�����T@�Q��0�b�B�(E��#n���-Ꚇ4x}���L�d��t'J�`��T��3�W�6F�J�}��vRV.=>�z��b%���� �k�'�U� 9���-8�@�(��g@`���oV�`�NM!����ip��ƶ*�|`��-���
b~���:2�7��J�u^�������M�����q+��ʿ%X�ǲ6>9u��=�����g�?�᮳{��'u�0�mOoz���/?JqC,��bZ�	?�P~fX����0�������Dr2�� �z�`
�,��(��f$�5'B�ej^�.�D½�e��M�N߁�ؽa�J ��m>�90R2������,P�`�N�{�vr�PH��[�d!��>a�������6Z�`v.�z���p+�o��b~��q@�I��IچS��'���S�R��H��R����Z�m�}T޽F"�~v����m-hwI���6�����OJ.8[���V>�<�㇟�E���伺�0t��f ������zP���y\�i�k	/�h�:y�Iz2���7ŠejȆ(��M�p��
��n$'�$N�/����o&��2(���E���������+1��-�2��T��T��P������e���<x�;���0ȋ4���|�U�B����"-�Pm$�|_�^�ҭR��o���*0 $̱���ℏ;���4,���}�_�{�vZ9kSIS?�$YKyW��^��8S{胟~L<�#[O�,���&\f{C������:�Yv���l��FC�/C�ޢ���1�A��&H*���;�S5TD#7�O}��d.L㵈�ވ�ٖ���$�C4�9��W�b�˒�;]��A�!:ޥQa*�q[/�WJ����1�Ю�4l�4����L0��}n.�(HQ�׃Ւ�̳� ,�-|q�w��LH��Wj���U�d%s�s���yz$V֍�D������==�=��_[N�Ã�7+��7O4Vk^ٵ� t�����2�c���Y�nU�����E��^o�n���l���X�������鍶�|��a��[���4XtGiZ�\ېs��6�����v\��̎x�&�X�����ư�G�aG�!0��J��0�F4�.�OЩ�h�q� KoY�o�C�K��e~ũ��AQ$1n��������jqi�z(�8��e#$�*Ϡp[�������9e`(�=�Ր������϶��<vAt��(䥕GԺg�^������u�NLBTy�
��I��sd�4Rs���aT��f�H�kv���k	����C�V��~��d�rL�r��?��4̣:�=Ya�8��`���XX m�����˩�<6Q�rpd�Z����ed�2��s��������G��ToE�� A�m|	�X��T��L�ꙶ�=}B~�C��Qk��L�e�8�>{�#�_�1e��ҭ�j���Ŭʳo���5&/�&*�H�M���n��+���5�MB_�Q;&1����m���Y���K�z=m��f��'$w�aχ{Әd��TP����tN�5��ğ�,�F���ت䚮���JA�s�H�����鎷�Շ�O��jM+�}�������_tNi��ȤÔ�'�(�%G��?i�+��0i��ZN{�����zګP�HbvqT'��:"��U!�
E/��!̌(��C��g����	3��d���>8d6^�RL�]߇�=wL��W~��>��&���g��&�|eC�1h��4����C�.L�f���"����ܩ�j���93)ǁ�Ɍ�� 9 �1�P����]O�� ��9��x)49���oK��	�+���h�zLo���W��P4�C���
R��.Qc�Ś��*��b	�ᩨ`�(xڌ����>��,��bL>�m@��&�k�����w����+�p���`s�3ꮎ�+�J����t��$aC����u��{���>Q�HZ�,ȵ���z��pE`F�E�O����M��n/øu~���׶يµ
�Z�T�� �"*�T��@x��;�1���Z����R���*�B`��Ia�N�I�����/��i�t�g�&f
��*c"���nFrN���Q����?�1i�M��[a�k�kZ$GNJ�g�Fg���t�v[/�'��h�^��[C��R�}\!g�l3$�o��}�3�����<�i���5��X����5{���KK�<I|rc���|���G��P��׎�"�U���d\c�H��=Q�i3R�䎰"�cU:b��M@2�Np��"� �5�p~�64�"�c�E� ���lM�1�`�W����\����i�{�
�ɹ�u�滜삻�nǘ���9���o�+t�*��w�����Pf>�޼�:/�n�g�� �l�<ޝ/0�p��|:���-s�Y#��Z�ߏG?��r$*�0"Pͦq9tB�"�E��t��$�l�VO�P}d&�c�oXy4�.OPg>5�"@pz
��NS��	X�U6
��w*�s�{�A��v�.7j�B�lFsOؗ�{���%�^�j^c.��/��M 7%���D��\?� ���>yB�%	��N����I#�T�k�7�����Y�XIl����A���μ�bt��oU��8�J�1��h���ZA�+/��Y�� ���?Sr�.7��@�s��[�_:3�|��x����u�B��R6d��9��R���2��O�'ˮQ`f�=e?+�wٰ�p?����̓�6���O]�����f��>O�t!�:J0�B*Q5��z�
z�����:6��1�?��wsum}��oL`��4U5�AZk\����o�9k��B�����9E~����j� �(�߾��(�xSC�7�n� ��^�L &�We'$���W�A"Uy���*wz�{��)OP0b x�5�Ar4��,a�$ϵ�:�V�#ڂ���W���i�*x�M����ŅiQR�=��!��q�BL]�$���q~�N֫�����)>w�C�ۮ�3E��8¨ɶ��&�k��@�&v��'�����B��b��ߠ�:
�vŉ4�Y��剆|���Y�"	�6-d/�jj;p����[')�⤕�67T���J�4+�>ӫ�&)���'%����vz�@.y ������	��fV��Q�����K!�ri�Rj����\�C���z�:lQ�2��ޏ1�Fx�߳����x���NN�Y{���@a�z@J�R�R�����Ȝ"�U���W��t�nkQ��`a��mY�A`��sE�C�� ��AxX� /̞c+qF�����sp��2�����7��$���Hp���s���.,q��y��ޕٰ�H�<��]��_�l����{�q ��4����C�.�[�)�9=�ɮ�䵇!��*�z�)����mj���p!9Bչ����s�BK�qPA��k.dx�%+�;�MJT�Q��pF�9�'�bv�I�}F��Y�3�a�Zt9�J��}5*ܧ<��}��eew ��<Vƙ���9�5D80k���ŵ�6|��GO�|x�&j=�=����LI��T"`��\���:{`}�bG����K)��������*B��m	P~f�&���bL<�g�����I(�`Y|�
�+�F��d�[���O�Z�6Y�kJ��fC���y���9%�<K^*�*\h�C�}�G�ε+_��=��ـ�������g/��TҸ�ra�a4/=���p������Z��k���ېQ�.:o��>;K���lњ�3�2)yh��!��J�����駵�vђH�|�|�Ҏ��Q��f�������2$�>S�r���DV��?� ����c�XJ�=Q^����%MI�iGV"W��A65��p��xk��gT��=��6i������[]�v�y`�v��܆�w�4����i��r��I-�����2ATb5�K�F�~�3Ǔ����j$�3k�%T�VPc��`�������\��=fE���IkT	�H�GdLEq�6�la��Zމ�&�����!�LXsYZC���P�Nk�#�dt�CB%����'mݷ�&�;�g	�b�$o�lE;:Ur���9�2�#B�&�� rD��3�3�Q�V���1g�/(�"�L�b?q��7���ȹ�ǆ@B����w�8L�����	�������O�h��9��'��Q{��@��>E���l{��I�OD!',p���<��xEj�'+T��.�;�ɕ��腟�X����Y̆�]9���\imf�GF �k>�h�4V���\�A-l))l�+���;x�p*;K8��r�
3�Ƈ�،t8��Y�\Ⱥ��#�:������T�='b�F��i�A9�09�c)Q�8}�O���1J���K�s\�����~ �5�IƟ�K��rUЀC��=��Z� ,,�G�ޮ��6�\;,Z��(�� ���A��?�R5�U'c@�n��1<>M�YG��uSE`��N&'���p��~#nl�E�wIn1hW���WZ?Ɉa��G0}R �^�!n��dL��KÂ�	ꇀ�L��o���r�)�#�B9�(lۻ�=�(6D��gxq��7n�Ё�[ {�Г@E����Gq�"��cc�H����rc���p~��1�;��m���O/��M�D����	�J�&�ZLl��%yRJPk�Š�
A� (I�o��]���@$�J(nV�6�y�_��Vbw�H�&����§В ����yM��m�L���X��g~ r�s��L���N
!��@}�~�i������b"�#�$����Odo�7���΋N~�n����4�x�9� p%[YA��O��JY~����/��Jha�ԏ��!ڕ�~����A�Wm��'�>�.%�Q�۰�E\�����N�)U4gѸ#�]�J���UG��Jf6�1���xf|�!dgX���ҿJ9��Zm�4O�~*���j�l�
R�:v	�4]9_<X���OI(�Ȋ�;5�q��~uw��I��S�0���;*��S*���4��5�|Y�B��pJn^(bT��)��]�â�wh�I	��՛�F��NY�L��5����V6'N�.c����V�eYe�W�w�~x�^��m��~ ������Np�F1��@h�gx����Oc�x�8��KCŴf#�7&�99��(������N�ڗJ�t�&=��0����$�ʊh��W��Dk~�wQ�T�%���H��ZS#��n��Sedu"��6OT-H�ǟr��
^x�5<�0r�j�W_f��n�2�5\x�0+;������*P8$�c]Q���zՍlN�$��O���[^�hze�Y< z)�f�B�U/%n�-NmUϪ���7.����h�J� "=j�j�{W�[���o�:3ު��銮5�l��ăT�}q�\����o<���K��:x����#���(g라�a���� �&e5�S�ףd���7����]��PHQ����LuF�T�Ptޔ�D��Sކ�l�����!�ޠ�w�̰W�`IZ]R+���;5,��o $�~�F�$�R�U"�	%��	\#�+I\/�a֪�\�<��JhŎ�0~�Ʉ]0�/��p��>"\Ɔ�������hg��(<bf�ў��;BQ���bwtS��u.i"�d\��@��f�YgC�Y��/�}��TuQC��r+n	�ɖtAs�&3������
r�����e.�)�IF�T�5'�hO����4���(u<N'g�nw�s�Y�3�/͑�⪡8�
-#}TLg�����cL@H�)�+�7�cd۫�e�n�{�SH���$2��6�¦�;�''�wmj�l��(��$�����7�����s������#�M�5g�$���h�Mü/���@m��c�0	���>�9��	�T���~$�8�������nH�JX	�;W9�&��
C��>TW>�X�CZ�q�6>���Y;#��S�!_����a�6l�7E&���k�f��|3�����2�ӌr�:k�{G��0�ٽ!hu�2|�[����Lt�!U���R[�.�X]m7��/����9d��Q�RAZn��88<���$�Z��x�T~߱�66�ߟt7гe�F����{)����f/����fQ4n1����
2�o��8���~��\VK~��CՔ���������������{��:	�	��x����.�5Mka��`Dfs�S�L.���(�2�<���d[¸�S32�t��߆u~'�=�wn���(�[c�<mn���4�3�}O0���ÚW��i�z�w��"������ʦ�Sय़!���g�~nR*���7�#<>%3�m�Q�"#�`�����&��o�K��Y���G$�DN��+���?-�js5�a� ]������)���p�EnKF�����
y_��o�]8�t������ʕ�j�����HL�M�#|��+�A����X�)���`F��t�FY�/�C��B����Y�R\����%���8��Q^0 �E�g��6ʮ�g��;6������a��6X@e?���P�yS���[������'s�/�r����׏p�<P���7��Ў�Eu������4"O��r?j%�ІN���M���k�1��Z���-���(K�Bd���Z�s�O�����l�4 �\��_E�  |�(�g�eqW��v
����R�P�P.`��v,�1B��I5H\��| �e��U�7c�սl?o���uMn����58��)�2��Y�z#�
�X4 Nt)!\��̼ή�
0=3��X�6����h�m�Ku�mA�k�d��N��։h��;I�tǡ��a0Z��J�)�bA��D4<��}wcG7��/M��Pca�¬m�E��]���h1wǕq����р=-=�wX^��e�{6"��X���h��F�|8Iܩ�ق#�l4���d��gV�2\C��gH�u8�W�	W��G;�qZ�/Gs��j�T�R�^S���@���^�ƣ���p��������4���d��b)�x��%߳n�ǲ�;�(����~Hc���:7��b��ӽ=�ծ�64A����BFs2qȍ|���7�5��nC�ؤ5��]z��a��38����ύ{S�)UP#���
 �g�"�\F�y�4k�+cr�����n��J7�^jCs�Smjo�q��&����T�_p�r1�r'�N�z�_ꀔ�6�W�SL��
߃��?kk��I)=T*�tf��aE�A>������4�^Cm�-�>�[i�˛�9A{�<X����r9�9�=�om7���Y��0��.�Hy�����*��>B9��c��ࡖ(Kтw&�0�8�Ӻ@
��Oh�FV=3�Tl����"o ���Y8~�ع�2��7N�*��������h;ס-E�}5T�Ͱ�`�Q�
����}Fã��q�y�
K�����~-<2�6��c�O�����wv�o!>�f+�搐 �:8>�x>�ă�` ]|r86 ��F��` n?V^%��]j�i�ӣ$�M&���IroʚC�׆�p9	��B��J"�e��>�e�}}���
BX��`�]_�V�D��io�~m0�Od{���f.f�6�	�<ҫVE<g�|�!D�Xm�(�&��7%I
���
� ��I7h�b�g*iV<����9نA_��Pn��L�^)0 ��zv��*�#�>�(&T��������K�J�}	A�_�;?pn��
��� �gj���V���p��%i�,=O1Gȑ��p�D��DJ��]���&ĞJD�I;�M<<R�?.l�Q�����Y�tw���Kb��a1�0������9�uD�g�>�O�cy����E�+>c5��!�5D.!�yK��ǽב���2��&�A��s�4N��Qُ���'5��s�1ok�F�1 ������8Q;�`���R�=�� �OWT�k���:K�큈`Vl=�y�E���֘*!I�ǫŉ�ȳl�����w^B�-��6r�@0�1,�lo��䭡pm� 	����ZcR�L��������֞3�G�*�U_u|��i�y���;9���^�ɥ4�+���hߍh�m-���)�n�2q����q.-�3~�m�n�8 M�U�m�Ӧ.�e�����Jм���Q�,Y��%�U�7���d�}������F�52�<U�+�.�z:�f��h˾<`ec�)����H6Y�R*#+����m\�I��Z�r�"���S�D����^Ãz���h*������Ǹ����Ci8ts�<�%�7	\H��9�?]������]�N�\��sg�[�y��D��D��Kp���θ+,A��J���R��qSV�Q��?�|��w�"���N��Y\�/)`�'��lP���e�	�ԙ;�?�Jɶ#��B:0y�Q�_%'A��Ղ�wx�v�K�Ƃ���g���ɹ��d��tگ��y-������x���
�<~����/^e�ا^>W	�)BB�%2@��8���%=]ﭦib2�Gw�#�$"��`l���Nvvx�eQ��f��/;_E�K��ɼf�qon����[l�J��bܯ�ȣjDk���[������^���C�3��d:G,�!O<
�0���H�o�3Bc^mU��愇��Z@)7h p�V��NL��Lm��
?f���k��H+��h��4\jf���{�BrGj7��b���,�ub�?���:��0"�b�t�aq�2�9>> �&m�w|�hwm��
��c���� i�%�D  >�-,S��C�B?x����� 7擀�wa��o�]��௕�[�ԧ�E�Qƚ�����h�u�����(�<ׄ�!`���6Ŀט��R�]懢��A�;�i���>,����c�X�;s������ǃ*I�5]_����T���\	�*ȡ5�YX~E�<a�UԊ���D�O5�.�Kq�8 ��)��H���"�}X��.�ћ�N��Ùim�.����lA�}��s�9�8א���@v��3�@o���h���8�b��UuoX���O�ωP)2Eڋxbz��֗J(�
|�CH
 W_��|� {�e��
�$l�^��(�8	���Bc^��,�G�����/��`zW���㭓D�}6m���Z ���(�f��;���w�%��0���?��п/v�*Ƒ@�/	�Gq�z"���`a��k���O�ԋ^�V�}֣֭�SϘ��(�sKB��96��2��h|_j� ���ے?JVQo���[Ј�tG�����ٛa���w��h�ݵ���2����V��aE�;A7vY���v��Z0Џ�º�w�A��ǘz$�~6ɔ�_�n|6�� ��+�u�m ��q6l&Ms�ؾDŉ��p�$��;�<�[=A[,�*7x�*�k>�q��DG"�z�p'�#%�	����Y<޷l�i���'|3�,a^���9b�53�͠{|������q͆[�{'@���Y;E��<5�~����[�����w��C6�GGvB��������TV0n?CWe�q~����P���Z@��/�f�9s4rP^�T6W2cp�$t�ɚ�8�Q�B����@�,��Z,]o�+t2�PXj�ek�E^�6'Mh5P�����i�����l�y��	<��q�V8S�yǈ2h�?}mN��a���Xm��m�a���\���p���<�b�-cn�"�#G�zGEj�)���G�Զ�hǮfϑ���p��H��k�v�]��� _-K�L�W�xi����`(r��n'gu	�?	�:A�ɷ�G������(�c���T1"Mg����v�?���ުN&}ݹ'��#e	�ĩ��-<����F��,Ϧ�@��9�7{��xw����Ε���B���}�W���O��a
�r�ٗ���wJ����{�#Z��A�����w�ef�d�Ra���Nj	�f�9�����-�ِ���M��;�@E��q>5z�2�!�O����W�_�s�q|Y;~���G��30�>���T��
q��fCd����6�a޽g`�3��	5�p����.��w'�b�0�2Jo�a���1|p��|,���HJ)���D��u�x�J�Z��V؁_��f �������Q�u�E�
[�]T��Om�K��J�U:ys.u��߯گdӾl{���/o��J-��ōd��>�K\af��)\��/�m�MÇcE�j�Wt~�z&�V�mX�t�5w��L���k�4�'�L�~��<���ߡ#��geͫC�?}��gjjeG x(r&��ZɌ^Ė�_�����q�������e!���8���r��ŷ���m�@�7�t�;Þ��F��] ���.?��;c��i�ol�ZT"�eD�  �W �x���3aZ�[�B�V�{�7�Y30��WX�1���];�o�i�5IT��5c�{v38�snM�$��:ԭ�-G�BP�za���S���ƎLn�5��%u�p,6\eYM�=Y`�q+��r)�j�(���|������Z2�+	A ��)�9?�	�w'�J�p�g��cr�c!��I���*ʪ��+�+�~��!���Bγ��˾=���)��A���+�!��\$u^4��<3q]p�<M���Ũ�p�p��P�v�{�M��S�.(���K��[�U�rme%��
���7��d���F���h] m\I#��W_�[�������Aʸy���̛��貀�j�V�Ƹ.p����o[�R����?o��Yy���-(����j��5�D�ۏ��3���flħ�5��ݗ�Z�t�6;t4��h�ث)�[c�[���I]q�ap��X�x���2[���,:I��VB���pM{�A�x�wR����6���6^c)�l�w�c�ɧJ�Sr<	=.��$�D ��9�F�ﮢ���N:���V���FѤ����;!�ѓ�/����&�T��_��4�+���ձM�N���r�fP���۳Nzx�d@����V��RR(�3�V���o�&��)�)��e1�Uϳ�u[��p��&%[;O�%�CR�٠զ���?���g��u�юqi������\.뼯�n<�{i��&Yp-�/�2u�I�'a^&6���*���?|�̥7��vl];�!4��g�f�P�Z��2>~��qq�l$|���=����uT��U�Y"�l�1���`���Y��Z:O�B�AQ��X�D �o���tK�%��d�]h�|j��MP8AN���;�������זSaީr���ƙJ	��Y�������\^�xF���R��~~�	(��w����"�f�K�]8�������_�m��<�p�� ���k煗k݈�di8�(�#�H���{
|n_h����b�Q�%W�v�z�]��*��x-)�ܑ�N�~�t�:�����[�(���)�L�g��0���������hJ)�j%��o��&=d2�׍v�������~Eο�b�yzV��؃�G��u�K&LF�\Yp���\mp|��d��,���h��K���k3�{��]�`W�D����1}�"AXH0/u�x��W9ج��8&��A�{��棠i@C���ftf"�B��d�ǲ��r�f����w�hPt��e^�����HnH� o�������L�JZ�rw��u��ZJ*�<p�t1L�=���F��p�3�R�I�V�䬋�����{F<[^J�_n�,k�$��Y�9��;����ȓK˾�s Gp��F�ꩨ�K����|��)��Z�P����|K�,�w�b0[5��n"����c���¾��M"[uȶO@'��_.�N���);[��ĳtUS?0&�@]x��^�w)�:�����im���j�\��w��8��0���2;s���	Q'���^�W�`}�Toi�9w��cb�k�7�r��W���n<r1�Wp�Ym�+�i�q��y;>Q��:yaS`_0}١��(,�8��*�>�Y�[*���O�W]��)rP�Ĩ��{�߄���"{J�T��y�9�3�31ցlخ�ܔ[f���Fk���J���a�9M�]Ζ���6`���rvֻ�Ȱv�2�.z�����Ϙ݀�ܰS<��+Z��rQ�t3�a��ߦ�@_|�Yt��A�G���u�<˨6Ӽ��,/�	;��4�K�@)�1 Y)��-��� 	!�����U�z�ڎ6��A�M<q
���Z ږO�?qF�ЗMI7R�]&���jT�R��%}�6�ڊK>����:�l8�m�;�>���H���7���'��?���AD�=J�*��m��eڀ] �C�il.�	o��[tTc5R�C��ԭI�aM"�2�]#RS`5�7P�H+T��4�f����"`������׸&ھ3̷M��Qu�5�{oVE��B��ĸ�#�7�Η��L����:���p�4r�:j<�m,�<O��4�|yp��uU��A`<�U)ߥ�]I���}(�I�m�M��2a�Y�jr[øS��*����ue��8w|d%دE*vP�"��va����.�Ʉ�JR�m�8"���/p3��B,y������Y�|���I�
"�j̚
6�|�"��tʆ�yow;�ݦ晲Z�b
���@���Smq���~h�r�LKB`Nq�GX�tj�F�L�.�ޛX����D�CܶW��6��@�h2\���-�0��W��>�~rQ_g�=�B���_�S=Mk>�L�v!U#���F5(�����J�������c����W�Xn�䦮Ϥe_����U��YW��ʹ;���</���kм�Ժ�����ҡ-�:�"����������1-��}υ��=2&��vz��W�V�q2���y��uPC<�5�x�ᅅn��gڛ��O�#8��#��\f
�(��� ��G�k�CO9�����w���b»��~��f:�v���D���� &�w?�d��h:K|#	�2Ӻ�aH%~�с\sG�Ĺ rD�)���:�F*��'hq�ӝ�?�a���������Iu�T���K1]�P��3`�J�j�w�a��W��:(Pk�j1ǆP}sp�)�о¶c�v��$B��`?.%��Z���#��3�ؙ��)m���|	�v� 5�Y�k1�k�>t"����U���1�(�1�;�ƛ�����J���Q�����\��4'�.�',4���#i?UKU��+K���6Z�?�Kq3>k�� Ko�F��N�{>.�_$�߆SB��2K�����^������[
H?j�Ϋ/�6���C�O7W�����<7����Y599�)��^�}�Qi�'`V~;Ҡ~[�����p\ɏ���a	B��t�w�9��A=K�C�T�Ɉڄ��

�z#��bj���Z>�-.}��fU���%���1��|$�~�Cj9��uK� ��#���aR�P#y��"SP��I�ݤ���1�0}�7%k�J�p��U���R"��#y��]h��[3c���N�l��#���jߵdl�g/<��T�2]��ۡ��^x�
���|��{��ky��������_���+��q	J�)��d���{���4i���ؔ ޷�٣Ҫ������(�-1����;�*G�;�{�Wyj���N�r�%�1��#��I�n�z�t�O�ԱE5���^)`��D���ߤ�m�+�?G��`�2�Ux�� [qL����QH�����<��X�4_U@b�#�����{�v��һ�vz�X�F�@#�|��$�2�}Di� j�?�%�>At�2��3�Q��{��#��/812��ճ֓��V����F���E �c"�Dxvs���\�8��i�u쒋xP�QS^,�a����M+��+OB�^[�e�9��c�z���Ǆ����t:`Ra ���~=��%Ⱥ�q�m	qamN4�7g��4ܾ������@¦���ه�m���� �+�V����RϢ}V�Y^u �ćG��ޅ@/\���L�x���0�J2IBW�5&&��)jI�H\0S�Ƞ.����?{�:4h�+��4FS��F櫪��miFUg
a�`ŏ���;��}J���[��0+T��mPZf�0A\6����b��5�b�\���m/qz{�T4�W�H��۲�r�祇/�1,�,�튚���d��<�Q��m�~�PV���r71����Æ�*����kZ��0Y�6_[Eݾ��˸E��>����QW9����&\���CLe�zG���|��h���d�!�s����D�$w�X�"�`\���ϥ�iq�������#����SyH����iࣻ���t�mKK\�׉�b�Ƿ��0+/B�#& &�ɖ���cz��G�H�#;�U��&���s$o"���bR�1/���z/��|R_J�v����R�`��yP�5�\b�I��|à�U�.8��)U������4a��Ɓ���6H�'�Ȟ�SO:m�3���b��bY�f��Î�U�����6�@�i��S��y�t_�X�BJ��M��=�Q�!��Xҧ\1��,�'��1��ꙣD��)���2�c��6�Z�8 -���m�X��#<�����O�/Q���Nִ ���L��8�W���UK-��	���ѩ��}��Eo���Rpye�|� ��)�'�!���Pi�D�*�6�w����.p��;��ʧ�V��Jr�Mɤư�_^R��x�4�0��1�C��3�nG�3���c�r�ߖ4�9^v�zD(�rz�ޑ�\-?nNVnGI���Ԉ#�TSD'�2C��HEջ_ud��Ho�>��9`��4�� ���?�Gn�V�>�X��H��G�aaѝ��̤^ǩ{>���K�������zDW��G=MPqJ���5�m|���5��f���!E��Na,Muf���n�g�Fџ�ߝ�p��Y}�<GF��
���F������]Dl�a��(�6�R�Tv�p+?(�
E1*"�\عU�f~ПT�=?̋'B���|X�˞��r�&�6�˩U~��:��tG���ܾ-r<�ȩj&��X�@{�=z
��xY�{Ur^��[k5�:�[�#R3Vw�=L6<�(�e �#���"���t��@��Pg]����:�����/}נ
����,O�?S�͛
�K����X0�YP�����U��m!�dʙ
��ܛ��[V����`T~�|:��XZ?�)!�y�n��:�NY鮉��u��;�e
�k�f�tcCQ)�k�ؠ�{� T�Аe��}<���w�`D�*�`�����+�N-F�c�[m*@|F��w&����㊀T�}�,�E���ٚo����j����q#���Rq�4����5�H�:��o��&7Gk<�&�6c�����IJi(�~/��e�����S�*b�ehP}%qO�&��m2����52����E�#pV��-8�	��M����u5G�=�@0*�4�@(�(2ؽR�Tȏ6Oz	����NV7��N��|��ڎ������b]3�FP�J��E���x-/:
:����p]�h��LR�]�f�3�(4�DQ��2�pu5d���z���KA���kuZ{7�w�r��WŒ#��XB���nC^�[�\7��ÎN�5�鉇vI����������|GtبGt�L[��T�Y�0`F$!�"USQ��
����E}}����y��hV|$;"x��Jg)�;+-c�����\�ܾ�����M}�qf�(����C6Y����Yo�(1J���'V­l+7W���<����� cH�C�^ل�b�n"�#������0���4ꌂ���n5�(�כ�I�7=t���
��A몾;���NXC�Bd+uv��|�"Z݋2v�搴��hFUC��ӉcK��}�u7�pΌb��S�m5�$ G����`Ǧ8y���2�/l�\nĊ���<4�&�&�M���7�ʻ�A#�}� �$V{�A��X�z��ED��B�	��_��~�O�?�{����a(5B�-f��p�����2���hH�)�b������Hv�n�SX�t*O�&�ϲ��ߞ%�����hF�ex&*)y�JI�,���o^���r�C?���l.� 5��TF�^@���P��5��̝��X��'eo�e�1���D}�t7�xߥ[��Ў��o[O��%�=)���vQ������9U޲t�  �d�ҿ���f��������P�D>�+9ڠ�j�d��%��8}M-������<�e��|zd�]�"����9%(:6��y�X�ù�vn����֋�=�?2�ucO�~_vE>�%5�Z)���������&��}��JPJ���*(�m���O�T|����:jzN����a���f�C;�jCV���%V�.�t��P��H��6�
��#�����0����+ۣ���|l�إ���5��.:�DtM;�>�|���v��0�W�z����)�D����9��F\'�0��p��+�-U��J1�H(?A�,��v@�R"�a�S@��o���B6�/"�
����-[��K�"'��Z������������4{dO���X��:}iQ�w8m�U���6_ZN��iɦ�$��U5�W%��B2b�
]��W��?�&�7~fim�^��cm��4;��ټ�ޒⲜ��{�v���y��h�5+�#����	��j���t�����G�z0	,��*U��I��un���������>��<Ҁ�\�{��I�tz%l'Lp��(����/�7���7jY��.�ί�!؅}�4���Fnxd/��8���s�f��C�������?d����^�(O*m	�Uo~�$�	��B�9����F�&k ��Z�-o���yT��K\�����Q�ܳ�j�>n���j���GO@]OE��*"V\���]��h�3qM�cu]�{���	a��(�rNM�rj2KdQ�_�_���P����(�T�g� �c�Ix��yJ3��B��EؗO��t���R�cb;�Q�u�S���T��Vm��ޙ����.�Ɉ����Mj��g���������_�M�6CP�&_���q�Y��*y~<Z�r�z�G��0jnk|uV�ޮ�|9����ڴ�Ѽ,����zYQ0��J�b�[Ӌ(�����y�c��$�I�Qs�?8b�%V�=z;�B�a��+������~��`S����k�oA�skW3Gxo��0��$�a�Ұ:�����u����d��B�|�,��`�H;hD�\����[�~���D�y%��+�����}�Q)�= ��+(�J�l�Ͷ�we��S �T��W�o1�8�"+^#p�� P����KCU��%7�?>��[���bk��@qUm�}�V�Gi`�Yf� �/�̜�I#��j��&�y�^q�M�r/����kQp*R"+$I�5P�'��}s�����Ca�wN�ED��0XrA��
��ZZ*��9ro�J��٠�v%ʟövx<÷�Gq���E��Xެ��
 �e�4���QǇ�:ד2�Y.�F���CV�S���
�H�2�*�n<q� P7M������  W��Y�Y����x��H9��3��U�S�J��Qo�\]�D{��uw
u��z����=r���S�|q��{�D�V�ED2���gS�W����5�UH^�\�����o�5�m� ����tD��rd�6�qCφhĬ��E0GI�ڱЀ�����yi���B��__��4�^���=�ns7� rAu̡((>�$���Zd��l:����S���1��-��b��?!����We�5�"g�ӕD��vF������N���2	1CP
37��'�{n�71�B��BXo:F�͌}ʒ�;��]�&����J�m|A�"o���&��Y�8�#f4E@�O|$���DM&?�;u��"/��G*���0}��yC��T��Į
��tB�c/2
>�v-P��u�[+Dg pΉ��K��B��Z���'А���V�ϟ���6xi�=L9�b��\`H�h(�m�+q�A\���2x��@�w|9W3�AX����
D����8�������q���u�����"CЎ"�j�Aj	�ia��
'7�����Z�s�\^
Q���`��4Yڎ	x���G������1���v7A���LC�͜ ��,;$�1}L�M-MH��B��͠�;���Pi���� ���]n���z0��8��Lg��T�(X-��yo3�F��:�dU�ů1�+"�Gl��I�l�����/���~Iivu��A�����ܻ�}Z;W��#�n�A��-6�&�S���`��z�ϱ�6�5�1$�{�����ڣ��B��p�ܽ� ���kQ��`+�*��n�ڕ'b)ce-��n��ſt���N��"�ล�p�={[w�i�tL8����ɠ���|�>�
^$�����Zc@�v�U���< K�~�꾘��z���lE��
m�s:_��>�-����\p&���C��ђ�
ʃŢ�~Px�H�Bε	eZ��{!&'D�6�c����=��X�"@�6���2q:�e�E3��=��]Y��]���h%�n��%�rlw��v�c��ߖO�ϐ��� ٜ$ �+���7e� =�UZ�3uАZ�/۟�씂QgAl���4g�r�2���/��3p<�P&5`��z�?=�V�1�*�Mf�$]P��Go�'��R!�s<P<5���Ʀ�#c[Z5zl�
�^w����UXq��*���͕�r;����/�Xݴ��_�'�X�)���4�\���A֢��v��
H����Tj:�W'�_�o�v�{�.07e��ְq��hx�+�������9.0�b��%\sd}X�#�$���?.Q���bT��%�,����$Bt��#IR�V�\&�.ꭌ�'�5�do�Mz��1�O��_��-��Jd%b��3���_����b,5���D�	�s�U�0�j��<E�`D�Ŕ�u���8D�Ӄ���M��g�:Yлg^'.���R�S�5��֙5��d�(�ѫ��n��/i���ηA����o�hԥv
9U��&íd��!�N0�#̨�7��5F�iS�E*߶G[��3ؠR	e�R��S$��2��?_�y%��\���ؾ�F������ث�!�ޖ#�*�b�#�z˺��T5!@�=�ʽ�q���,�]L�tV��"n�%�x�g�J��FE�a&��O�/����M60=b>2�8N�Ťe���L�I��R�F�p._�&��y�{�HSء��*5��J��I�Y���_�C�,����#�]U?`�%!��%�R/��*��v>���d>�>s�P���?JM�y<�̒"���L�gx^k ����0}R�%��a���%����9j+���s�H����N93. ]�x�P���T �{��A^Ȫc.�n^ʕz&�"	����Ђd�ˑ�OTš�����D���r�)�B+�G7�)�kmL ����T(o�<gߵ��@�ep���o�/�˝"X�D�����p���_�jU]�7$D �̞+���QOV�c�3��xr�c����E$��Br�m;�/3��+{�(o��(��
��
�ƥ%�s�4��p�Ur�J�'�J]�l��/ � �a����d����b���Oq~�Y3g�[��ҨqA��aĶޱ_�9�D[u��o���
SS1E���y�;A,��{��g�o���]�,D3�m�.�ޓ3�J���:�����us�\��Vy(�I/�D]Ruy��u1"3�#a�&�}77N@�W�P�"Y�Q����;Ol^���Q�;���"]�H�0?B��,�Y34o���;�g����&!��E�6�����x|g9җ���u(u�H��!��Hq�����N��,���S��p��?������mIM_�I�v��KMj�?Po͵� v� � g���Rx�;q��(��l���ȖM)P� �D
G������A�����PK�1zF��xN���Y��vvF�u��+�#B7e�����jh�ʛ˫�������H�M΃�����g6]����cm���&�?tś�]Ȭ
\���y���W�^B�s�t��T�h��l�ʒUP�$�D��z��$��àJQ��V%�M��r��5c�J����Y���S��C��yw�'Bl�8v��E��
�ܗ�@�
����t� ��t�š��u����;�O˨�q����^%պP'8ni�v��<�!�c}���sZ� zM�3ĭ,�i�vm𡩁ڲc�	��$��k��׺G����d��M���8�\����`��z��߭�e/T)
�B�ŋ��w�����M:�q�(ԍ^��Go��)�F+�h=�H��%'��dzH�y��L�H�/���t�'D�(��X��.~Pq\8p�/�Cɣd��!b���*n��ۑ2tm�%TU�^�hAzewx�.��!�~�����]�J���߭]�ח1�j'Tp0�r���t�^�����TM<B�48�/�X�=����:!��Ʀ����p�%������+4�Xޅ���C����CS1���2��AdK.�f#SM��,=�#,�w��{�!s(�'I�|��/�g��#�{ImP�>�^�(/B� ��w��"�4,q��=�7l�e�p�/?Hçp礜4�eT��Ӥ��`h!|�����W���it� ԃ�)׏��:2��p]W"\
\��w�ɫ��NA	��;
�c��Y�X�o�j����FnA�m�4�.�>�s(�aH���G�zF�A�gW����L��s�+`�-:��|�ɩ��fR�Δ�>-�t��IX�ϟ�E5'o�&�sl��ƾmM��q+��,�=Hw.G�l��!"ÈM�����>G�E�����67���X'԰�k	?�K�*������d���[�9�c�j�7�9�#���P�A���3|S�슢R�Y#�DP32gL�(�p��ŹԀ�i���jcO#1����UH��>����&4����qsn޶�n�mN����Б��鄑���/��(s����2n3{�[Ŋ%\��1�<�~Ńv��%t�ĳ�(㻠�w�6��������fI����������aOtX)��;{�<��F��Y�cQ]�2V��:��ͼ�f��?��"l �XK��򻅌k*�X0� kaP���4��z֙�Ep}�D)٦,�	3�M�~̭aW�vg��q��5�_��;NP��:�����"X�j[NTT0��c>N�|�}�w���t}X�|$p������9l�C]�嶁�OE��~�R=΋�w�u2	�t���<��x (�wK�=AkÌ�TH��7�o�ů9I$Y�2x����g���N����Ӎ�l|��.��ޭ��&Z��4(����4V��DU������/i5Bѻ�t�}��@O�Ǣ��La0OB٪���S�Mk@��/mA�l�؊ųTܶF�v:WMe)lM��}Uz��~��� YТrB_��Dx k�\��ɭ��V�>6�����>j�d}&'��q(֋��$v{<*��H�6m�� ^�UG����`bQ����θj͊?*�g�a��}ET�U�	%��d0{ܣ��WoA6��ut�� ��3�VZt6���%�h���8E� �lX{��7�u�T�E+k��oc���M�5C�;�s6|�I��XF��Nm��!�ɴ� #���zK��=�z�(Lg7欑x
{FN�V����0�X�O���=@3��Ep,��	�{9�S��`ZR;�
��]m ��e#}6Z� �IK𸒬��B��mN<F���nC��R�����sE�I#�/�}���i��X����S�BPZ�+�w��V̼��w�̃���n���� �*r�7��8��P��#ݷ�9\���`	�^8��m�����e	�I�ݨ湛�4ͽ��;��'�Y�K� ���̼���>}U~K��z!�7�|���r/~���֛1z��/�lA|���*�)&L(�n&8Y�d�@3xlҕ�i3'g��l��%�ݏr���CGM�^�7�b���
�$_hҙͽ����'@�+��mM;f�T(nV\c�z?fH}Q�1ר��tWV��Ao&�A�D��ߟ�/�LkN�����~l�>&�	�����J�mR�k���g�<�I+�,F�̡���w��{W�6x6��6�*�&>[�Z�	�xF$��������;z4�L��+�L�v�&{�9i��~�!�'����8�B��@` �c�0v`A�̝�Z�y�T�R��{�
\n�o�5=6��5����r�ץ+�B����!D�Ye展eJf@���
�)���*��w�V/�\�]1&Ǆ�󧶧��ئX��������7JΚ�� _�2��9�>o�PB�X�*9$�a\��ͭIҸ�T�4�Ж*^Z�ahf�G";4 W��S�Bng2�VUv��q+�Kf�@��0Od�u1g�pg���5���9٬�%�\��5GW �&j�.��Eh�O�Ĝ-�P[��d�|�c�l���Dhd�럹;<݋�"������>���̔
�/qf��NAr#�+�9ܕp�H.3���m���Th�ˬ/&����N��e�!�?u[�X�c�2x@��Hp�3�/�_���@f8���5����\�I>���RδK2g���c����IN�E��ggzeo�Y�nr׀s�]��
��S'I[C��-oaK�!q�v�Om��8�ԍ<����0	 h���5B������@K����y N�#�B�]�`�v�N��Tݴ�<[���O�&U��0�n������:9�
޸/���2�
Kƻ���(u推�b[�(Z��π`��������HŖ�i<Ǐ�k[�A�u�@bJ�@Ɛ�w��mk$CS�EU�@�%�hq6i�}��跽s��&O��Te�@�x�bq���e���E�z�7��5�'�]`}rwذ�]�h���_�5 �5�j�N�� #����Bht���d�>�`+JZ��T.K�@���;C��d>�o�ԍ�e�5l�I�N�ɺt���Q 4 �
k(}�Z���qnT5��	�g=jU�YA����pFךF �F-�&M�z6&����s!�\�#r#xA��MP��m��i�/��D�T��at�.�;)m��
���~�n���d����O�ӡ=Me���zƁ�YZv��[og�eaߜ�d���F��0�ukQ���
5t���mD��3�m�q'х:\(Ix�hŪ`�a��۟��=
lY�ԅH����U<钝����D�*�="x}�FR����sb���0��M:Bt��c�s>�e��|�7�ht� �3��|k�Cb�
e���O~y��lwa����s�g�j=�xYXW{`������+(!�ł'�}�P��X��N[�]��vr$P��#�ơx܈B��	=m�?<����I����X�� ���̃�z]�1){1g��`"4_�������K8Wv@����q�M{�kS�	Ӡ*��Y���(�%k�|�sZ
B�����x_+�A���/m�+�ϵ=��o�Y}�P������&|�eׇ��j.��\w[�+�X"�͸��,�p<s�=t���ٙ���(n ��������#�p�E��#f~�Z��
m)�U��~��O� ϩF�y�_��Z�WFP���Yp��sV<��1e3��׌���9�8h��V���2�D�\�T5��$H����R2���'�7���P�D��щz"c���]�
	њ} '�	=d֓���E88��h�Oy5ݓ������jhP���������/İ�����=�~��໫ Q��+�&[����ԃ�4Uip���If�"�f+n�a>��OR)8Ex�镪%�}�	�ij�"4[k��tź5����'q;	���!��R�*�}�#�e�ंQH���ٕ7o`>�#�
���,^�̿����w�r�М�+�:�7{Q�Jފ>�6�j�X'% k� �˰@�V-��8�����E���녓�2��5�,���Pf��m2��?�u$
o\��`C��&6�+�&�n�A�̺ j8[���i�>��_bYS��l�	�� 6jNڃ�BHP��2ܩ��0�x�=�n�0¡�1��^D�`B;dI���s�t�X\�nl�.��m��5!����¹�'נ?������VM��($�g>��M���|gS@����'씷���Jy��w���8]ڽ !�{�_��=���ÿy����Ab��E�A8��g���|���V�>�)��e{C���(OV��^f�6Xg��_��yo�)Κ�;�<d��d����'9�T�A+<����h*���z1�Spod�n����5:CD�~#��a�_)<��Ӻ+�r��6�Xz�C'�F�Qb(o���ŋ���ԬG�PX�~�>Y��bxa�=�qq�Q�/������\�r6,��ʂ$���b��G�=7�e����ܪ�L�F��׫b)E�R��ya ��_O�g<��S�~Fe�'U�J�| 1bZ���{��SC&#�E�����#��_�	Q���~{��sK$y"Т��7�BHP]Dr5`���&��QѡƼP.�P&x9��u�/p�e=��,ɨ���r/��@M�VJ�l��@�qW:C�l'�B)U7k1	\2�Mh��M�@.!�ߐ��k��� ��xza���������_z��[�����X;�#(K�h�g�W->d�<�#{�w g%�^�������w���0>B�M��͊H�ԲF�
��ܷX��m�WZ\��{�b�V�0ĺ�����5H�������޹ZNIh40��ex>M��2Nv��A@V{�9��,=�D^D0�V��e��^�-0pC	&�l��G��V!���	�P��~����ۍh�\>tt�W��4%a�&$?����'�{��Z�q2j�<C$A����*EuF�ԉ�
��ˈ���$�^*H,�_8�� Q�`}��ұI	%G�$	���¦M��.92볙H�(�<Z�/n����������0��p�M$����b3��7���~w�}�����{7�z"�o�.���Rs�k'u�����y�'۶�!�������z�+��4���A�.��sF�.بh�8����ª�R=K,})��;�����1AB�T� 2�s3�J�h��0ɂ��:_����b�Q��-V���u�O�3(S �>�~~B;�_�Q�#k��\q��.U�������i�I���C���H�y���+ȿա�;9��M�МU�J���*�9f?��#���N�?>	-@�\�1�#6��@�*�����ViI�W#�ʗ��I��>̭���S���TQ|jXb��[��J<�O�Z�!'� �lu�,b����'�!١aЊ���Z�D��ъ!+�B�V�eg��b�f9�W���zikx��AAWn0�/4hG		I V�h.���"�vC����Qݡ�s'��|��Yқ#
q�92�!������|u���їl۠w�,f�!�����ؤ���#"��E�lQ���K��U�E��O��Wc�vK.�oQKS���Ά�����tƾ}l��j��������8���X$������bx��@z�q���n�W*K9d���\�a+��_�#���f��0��@\�j���
��C�<s�6!
�3L�Z�J���Ϊ� n������ȷ��Z�>m�È{��_��(Y��̢�q/`7iM�#:�w��W��gG�Z	�$'yeb(�h1U]�j>���i��͆�|۩�Ќ����^��{�s�zq�ne����-Pc�g�!��ſ2���m���n� �'.�<N���9��%Ֆ��JF�C�����Qr �7(�9	�)�7Z�����Dgn�F�bG����H���}OY��6-/���U�/!��]Ⱥ.�%���A'�����>csdbó@�#��ےr�'���BBT]��Xmr�P�Z!g��K�?>����k<f����IB��5eTQtk8tn�(���C�e�"�۴��k��c��%]�����K��]G���j :T��g�J�����~M��3����5\�l@�K���TE�L�߬���Naq���(��s
H���F�u5{W�h���9?�sN�LL�@L~Oe<S�����lvᴮ|�z�*]�7�JI���-����θ�n�Q�.��Յe	��o���N�Gn��C6͆�ہӒ�+l�6ۀC+Ya��Bh�32�e�w��]�og����yyM�>3X��?d^��?>=�,{ �^'3ݞ�hf}݅xG�'p��0nk6��Z��s��&&q��'t�O���ߛ>�9����YId�JF�^=l�x��c0�|�"%�v����PX�d	i��<��J�'8,]=2�"=[Q����NCs�0dq�ۼ<+7g�y5̧� �bM�����m�����@���G~)��E��^��_6J)��P��]i?��'x��կ�pmmŇ�;��0֒
WM<}ڞ}u_��%;�@v(P�6E���Ԥ�A?o��JS*���f���6�˸?��#�a�]���S�}!�mf#0?Џ��\�ݛ7W�#�{'��^�S�������Z��:���U8����`��Cֺ�d�iȖ�?R��K���]��7Na����*.`�<������u�j�]=� �\l�~xB�p�]4lz�j-�u">s��Q��L�5|���J{aQ�Ou�;���|^��F��G���X��q7V�׳j��[�
��9V<�,�b�I��l[�Μ�8?|����>��%f��xr3t]{xQ!j�^��������ƨ-*gJk"(?O�J6b��F��M���1MJ��)���h �79����M�?`�l;s� t\X��>�]ɖOr:�%����7��r!}AhH���M��|�"�G�a?߶�:�e���(��mԌ6����>f
W@<��:��
j��?�\f�W[1}��6���Dr�c��ۋ��m�� �i~�f:�L1 U����>�� G�O��u�
���݊�o%�Y0�A��k�$A��⟝I���^��^�̨� A��G�:m$��}�wG�U����ԧn�����i(�^�ø�L5��\�1����T%�	���'�s?�4i�g� |�g���0��C�as���N!�L;�,!������k�y��'��̂���D̵q��H�&z�	$����}c�3�P��'r��薆�1S��}���?Ά��,g���n$�Wg���8�����~���'���3�"#��,��6��e��[�ݗL�>�L�
�r�����r�4��΋�[�s��-ܽö����I8�Z��b��ޘ�8�0�B�9t\�I�X̕�ڃ��ܚp�+�ĖHʼ��<�ѥ�3���=ۋ�sڨBI1�5�+�S��v�J�	�����1w��j���uJ��:�𙰉�{F>$*��?�RR k��&ٮ�^��N��잱�3Ŝ'���!����Q2��<�A�ĖIa��� 4�a�X����[��43��x�?���h�[39�=���DI��!�2X�MSS�3���8��CJUw���*E-�
�Jn}�)�C-ft��Z�zEp�ɺ^1�5�{�{'���龛��&�rM���Q��n�z����� ������b�A�O����}�M����=��h��*O�EVco�\�q���{bQѠRc��&��(v�j�;*��=���0!��Y!�>�wQ�k:
�:����� 9�J���-�e�xԻ���&IW-j����|Q>C�X �+�2������K��	��5hq���l�u�&�8?ْ?iPH9�@�t]�t�#��G}�Ab kA2+�L-3n�'�{���UNP�י�TN���!�Z� ��UB���g��lB
�����
{�4�{�<6�߆}6���? �+����0Txr��r�5��]�{�y46�M,�r�|h_�b�6|�/8EP͑��m^tH�A
��@Ԫ-��Q�8��n�I��n�̬ܭ&	��A;�B,O�xk�E$`�6Y�/3%�$_�vV7����.lM6���� u	�R�P��Y�`@Z)��0��y2U>s���/�����ֽ��[!�\.�=�:K��Qz���]i1�I��dJzCW.�c���o��H&R��vJY�j!Yr;h��Yn�z�����|�^W��S�z�ۗ^�/���U�d.��Ž,Cۺ|�K?��'8�U�w���Xo��xx���Y���-�LҼ�X�2]T��[�c�;f��ZH���/�ষ_}�/0��+\���'�#迵'gzt�~�J��c��(�גr�oќ�������dݱ��O�4��y���X�_z�����������x(�qL�O�P�}v�S�#�#�ʪB�ٙ�9j�7]����BEAVt b��Hw���\�*��Ni�P�c����yzT�~g�Ѽ�w���p_4H�����HS�7����9B�{���r�>� ���c��;^�͛?9�.�O�unz���q������n��.�i3B=��a�m����p^r�?V��@��������j'��ø��D�)��;p�,&��m4�G��x���_�i3K(JdBD����RǴśҍ�,n�h~@��9w�/%Ҕl�7ђC\Q ��hJ?��3������ض�vI�m�����/�_Ƀ��O�?7G`t������Ш�f��^�/�m ����;�JU^^/�砲3�~�Y�[�
B��*d�;<�N�\�y�n����Ѳ`�4�zx�A	�>���Cz�zD����$�P��7��\z?�ĒZ���
�ͩ�::�n�dvh���42<��>�(uR��qb�rc���,�U�k#���hO�������D㞚@J�	�`|��jL�b���ۚ� � �=�M̜&Gd��>iA�R v6�i�0���7W����-)�`�~5��z�y�kǑ���Hˣvf�HLf�Ȭ�>�U�Ë�
T�!�,/$��F�T�"n�m������m�����5��rhebOӋ�H�v�I'P5�������{E	�3!'d���kcX)��RE�^�VhsU�q��u\��f���9�WL#YT�~�G�m��<� 1���U�"�Y��M��|
�u�M/)��L.2a<=bpƆ�$�r��.��n��#����?�T�Κ7ĕ\o FW���]Lc��Y��{�5[����xGʮ��=��[��8.�tCdQњ�`9��|�=�����PE��"C���R�O�87/��!���r8��+�������yu����Q�czv&��v���B*Bz�>���(WY��<T�x����vuK�wИ�� uS�fK��7�.��X��m�iن�8��a�N! S��#A�z����v�{�Y�j@H�:�o"�c��^2���2�c)T#�
������M���6��=+Fj,�U|� J�^�;��I��9�E��rX4N�`�U�uq(Z9^!��kkG8
��:u�)��M�����q�ι�!�G]Z��U�w�z:��i
}�u����n,&6��;��z�5���O��	�-�̂����F��\-7��p��f�z���~!m������Z�x������n9FJ~���,��6�(OP�B�:��JG�I|C���T��]�G�׊����HJi���G��d�z���j��g�(c��y�@�+~�8	4�)jv���|P�o���סv��zh.i��Q�d��H�*%8�O�Q4&�ó{R�n���w˕.��'�X��Ư�0�1E����o��%
SjӢY+��k��"��r�Hd���fI�<Ijw%�H��Q�=x�ޓp�維����o6�B<�,GM5o�Ƙ�˹���_s�[�`Xf��e�ݘ�q`V�<�[s�4	�{��\@kƝ-b��dCG��m�δ�Q
2�M5�"��"�A��k�M���S�*]��<CP>0O�o �;�C�������^��ĉ���tK�V�k"�~�a"�bl�M�w�}8�ƒ��j0�-Q�_q�I��ӶG�W�Z&��$9��-�#���_�^�"q��Am��sz�O��aɶ�Q�鎢����7`^���^�!*���Ox�\]�π�#���̷�ј�{� ��7\��-�sb\�wa�m��yN�0���Hl�p>��� ��1
U5����T�q���tv���fv���[�$,}���dzȉn|���VȘ{��y4E�ľ�b�w��ܷm��rz�ǥ,�8܇v0���ы@?<xMO�|�W�x�{Xc�l��Eb*�����.a�� 	���cސ�gj1�"_�6�9��&�*�U&�:�R��|��26A!01tҕ$ U ��)眈�/��1�����,آG���F��J͐���P�����ܧT�>{��Xe����}}�O���| �C��,J��-#��#ׁ��Q�*�fH�R@���ӎh#$|p�MflA	_W�i���c��!`�K�����u�\�j�qJ�H�@Ԭ�y��ZF���g���$\���������m%[L�e�"Y�g�j�B��(�����RSl�H�|Bi6>�rr#�>X^�p�K8�^�D,ܛo'*����W
�����)SZ�`l��VaH�`�7�&��}&��Z�V�hM����n��+���'}\@݅j�))^��S��U����*��|��c��lrӢ����K��=��Үd
���Si��]h[,v�BI|N}C��@xB�ӋQ��ۅ^$$��'�"n�g'�k%F�f!a�;Q�w9C%巰�4�}n!���;���=�|v#����1) �жw�N�����n�`G��v�(�K�;\�IT��\��Κ��x^p�	��J�8u�����P��	#Asw0���F6��ꞔu1ɪ&�肙�x��ES�o���\w\�C�C1�X�-(�i>	${R�o������I�omT�N�l�6m�]��[����({����o�D,:�Ee��(��b��0R��|[�	�����C��18��D֜�#�vG��3>6��+w-�}�q3?�9�c�c�9��1}�E��C�z�,����\�]2	�Q����_j����_�jJk�y�\�t�#��~h��>x]���(���r5̌�����2)�{�O?zH��#n+���-�V�n�ߋ�WM2�v�<}�<�K-Y�T��n�� ��g�IT��e9����6��kXo�߿0S�Cj�!v>��y��(�4�$��T���]���Z��tV�A�Ii#���>{\O��5�؉�	��P��O��ЁYX!N��	(4�"ieٗ�n��;�V�Z��0;����amX}�La�[�߁d|gך��:��pG����U»���A�#Lru!|w�v���!9�&[�E�	R�~׉���I  0�M=������#�;�������?�$�Ļf�}�R�X�G�<уg�p�se��O�xR�!��n�<5��m=�3$��`���k�H�3y�U�p4"��C����=%g�|���2զ4s�lv;.�Q�pi�tP��0��O���T=�p���t�����mx�������|fB["5�'Ј�{���}��I��-�2vL���i�JK�3(��Oo<Ǹs3�3�)��T��@	�;U2'v�l �@���g�u�M������l�h���a���=�Z��Ճr�[�ڌ%[ﶽ�+�pi>����U��*N}m�J i����Ό��=e���) ¯�tS����7��<�^d$�{�48*��_��}(i����Ր���Qj_�v��5_�ۅEl8��PY@� ���gܼ��F+�M
�&H/"c�v8���a��׈F9^�`�*'�k,�Z��u_�波s��̇�و�51yk�P4-�(�ކ��[[��4�^9�ӅY9E؁��(�浉��pGa�Z�C���C-c�2�Z�Lc�i�k�3����
tt~V��XM/t����0�e��=��^��l5GM� ]��8�Fdp
�}�#TI�����bFgb��g�����/"4ewئ9tN1TmP�u��]ϷU��WٚȞYWe�cL��V��
��ۨ�1��������0z��la�0��(�,���k�}9�A��j���z�I]��Qw���u�Stģ5Y�d8/P}��^0D58�ʌ'���$���p�*qpG*���;B�Jxd�S���hh����DQ�`a�ë���_�moU�Tm-+>�g�QGq�w����q�5GG�|�z��⳶u�#�!���B��V��C�8�����c9���/e={P  s����Fkݼ�Y�+D7�;4ԛ�s�����P����#x�/�z������-�~!�H���Ṽ���5Ө�4�S��I����ETR�hݪ��g�j��k��UV"��C����3]��M��h�_y\�q�ʋ'wY�r>#- ����}��?i�	��{{8p�^3��I�������(4Q�(�1��ϋ��)�Y��>&��&���Ha[G3�V�@��G\�K&�D!J������	>x,��T5�*xT�L����k^6���i�3�E����Z-�u�4,Ty6\��p� 
Cr2�S��yp&��ΪPA��L����O/�L^�O>bi���o���~5Uyl7��	��*��W-Szy�=�,�1@Yr��Lm�a ێT����%�0lõ$z�%.��:�Ԇ�B�B�f������؏�Ffݣ�[�(Qе�(|��ec̚s�I�b��ɖ,+�S���Y"4W �b��T�k �9�����!sv��~;���Λ5���Q�F����a.�M�jxt��N4׊���7yz򜿵EG��|������|�
z�I�/0�MR�eu&���.UGzX�),�������)&�Z��� �F���ޢ���W�ٰ�Ь��[�a�`N���/lY��:�N���n�]5�R�Af?�3�|�������l�$�������|#ɧ�p"�b��2����YB<���K�:�i����"q~!����7�7�#�c�i@Y�ac�W�Eyؿ
d	6�6�N2,�E�C>��ܺ��|h��,���/fj���L�$��G��\Ql��2�IϏ���a�����÷�3WI�0����L��3k��$��RJ�3�aḣ�B6ڤ�ّ�/*$�V�3){��G�+xfdC��b��#�+��pdOl d7+�N�gv?c�/�א�N��ow�-���z�慰��He��w��!�ѳ�o����P1,�b<�7Yٰ>�KB���*�!m\+�Ϋ�>�?M�*��pK�Q*QSH�ݴP$���ЯkOO��?!�Ē�+�S��Y�D���~ce���]�X�${>��. n.� 
�<�?E�ȹ�-U-0��%�k��Z�	�"�� ��o�Ӳը8ѓF��3�Y���N�S(%��"g`�aI�d�x�\�����ݟ��hm�Sևe�,PW��>�B���c"��z��6�P)����(Z.��㗲��Ѧ���CI*i����z�8��!]ґs�����??;����h-����tA9F�Pn����aƉ'�ŷa�f�,5�ay&ռVe�uj�� �0�"%o�W�F+�>+*Ug����+�<��L&N���ab�Hxf�����ey�=�����loJ�H���kKD�3X�d���OqВ=���_��Q0�u���C�ì;���=b~p�FIzE�����g���v��v��7;ȶ8��H<~c	znÃ)��Z��Me$����1�R$���25�6) Н;!%����P��$40��6�~��!�����1oFo��#�]7[�LJ�)lK�|���$˸y� �N%��	�����op`�_GH�
�{T܈Oa{�cJr��i�h�� ���y�*����z�1�=/�^����GX����}��C�o�����4+E��X]���I`��Z��D�vUq/e�ڝ�ٮ/�(g5+��f��zj�6��w:�k�S��Ov�1IĘ҈�d�l��4�f���T�l�g���:���r̖�ԃkPI{4�uBb��L��c��#�?��QN�?�oa�����,d̘G�$���\�!�q �	u'�ٵ�GP�XQ��q`�[Y"���,�6mpTok$e2�U��U�ܬF9X\�4%���ɹ=}v�$A0�����\τ�{��y�>w����Ӝ)܂��X�w�z�Us]���ӕ�����7��u�/Yؙ�̙�&��)V���A~�E�uyhB�%��������q��5tvk���3B�a8qo:�����B�ISp���[r���o�'��_P�N�aNP?%Ə�xb�T#1y��8���������z��r��7.r��R�0�sc��ArPH�7y�OK.��	׀���e��؝l�,���ۻ�ҹ�G�*�w{)=2�ܘPE7�I?&��'RnYo�T�k�S
��q��m�����1��-�s�]�ZD���\��T������a�)����xn ��>*�R����G��DAw�N���[������M�����1H�cO�D�W���w?�`���|w~�0|u��q@k)*I�X�d=�p@��l�ٵ7g�''��+v%K�z�w��7{?��3����%i�b���
,���	v�6];���M;~g���МH� ���I�$Ո�t�����&��P뎌�<A[)	�[&��A犸����%�����E��HK �#�����<��A��s �(�]��X��&�����oR�Y���j�6��"�؝%�liUp�My��Aʹ�k~��3� A�{'����g'���b�N=.�k�� c�2#���}��y�7a\��s�55�J�7������:�<�}�RS������:N�3`*9������h8DXo�y��T#qV�iP��[|���˰�[�:�;j��h	�2i��g�/B�m����VNߨ�V�rX�YQY{��6I�r�e�[5��x}wסL��zi���F8�"�j��#2ݨ� �s"�U���m������̢K&`��)]��'$�$���^[{���~Y�ܮ��q�ݙz�Yp׾�K��������=B��$��p��B�B��1����7�P�_(�ƫ���^d�Oz�nݬ�,�;ܷh�:I�4�+if���y#��7��)K�z0��\���`A)�G���~O��-�>�V�8���c�3Gڳh�A ]���/�  �������������Q#�d�����nkCw �W>)|}U���J��'�8@^'_���j
�N�?�~�`8��K��+�����U9��:���G�Р����.�g�/T��P3M-�KB���ׁ)��壃�bʞ�u��Ԇrؒ��y��!jd�>_�C>���(����y��&&��Bb�p<]h"����@�\�=�Z�*���#��k�$�$�~�9bq'f��a�ɑx��?�1��V,��@Ѧb��ݔ����G1���c�r��Bޗ�@��M?l�dá��$��~�<��T��q�t��9��SJ
�刱���,��ҿ���������U������LLxI1��'q�|�h��L���GđҸ�Ӈw}��Z��r����*m�i�0���,!2���yr(Hzv0�_	1���W���m���IUs�Ok�z���5����Sk�ӈ���D��g[k��15�_�/��޶�:nP�����k����: Nn;�<k���/f,���4<��@yĒs3���e��s+��o)��~S�#��:+�Ȋ:f^5}c������شr�'{k;dXe����Tu���-xK�/�t�OG�_b���޲�Wq�����o}�VA�2�\��߶�a��S�������*K���_�$i��9_+�����'BE�[j}���fX&,�o��J)�c�nɏ#OE���#�C����k{�n=7��k|�
D6i�5y���X�q9�P��\ �uI]��{�7we���0��[��K%r`֎�e�D\��;x����5��3��ƥ�}B�7Da������n��r��j��P�$|����隵+���2>T.��/Ґϓw�"�60���D���&���B� h:�2w��*�j�9D�,�
g�R���-��3�U~\�����U���g9��	,7�;z�?��_�C�on�rͷ_�Ǭ�tٟ��>���1�	m+��-V��(`��ss'���#��������ͽ�y�}uUe'�Hܕ�@�����H�o�Hjd75Tb�� �B����^V D�Dn�$G�`mSKÅ���4s�4;8�|���+�(4]� �J*m�Bj/g`��4���\>)��VZ���ȼ�2��S�L>-(;�8��Vͺ6�9���u�u\Ş'xQIW�4-�Su�R��n�wZ|�~���v��?yQ�8����k�}�b��A/֚�<�Ff-zS�+�=,]��M3��r�àf���
�h+�D(!�M�aq���Y\5r��VT�l����I훶f�Lݫd#����>9MS����8
~��  �,���W���
�_Pb&pq"�~�v�1 ʕo��Ԙ��+_��ͱj�~��>{���@�߷X����m.�W�#�x�|���@� ��ϥ��w���^t���"HU	F�����[�� X*u�L�����Mh�W�8y>��7(��EB�e?Ƕ��]�&
 ��7b�傣�%���ˎFP�P���D�Z��J5��&6�����;�̬˓;���o=���8(��%ů�JK!�i�U5J.!�	���F~�o���i�=���1�
\�/���i��7������=�,O'�LC�k6��z��nK��sG��b����^�Ӱ\7��u�^�̑��qe|�̱%���E1���� -Xrp)=*=�u�wm�V���Dai���P�	ϒ=%Uh��]���V�)M�\�������=\��"�����{j<�?��I�q��Ya�ɾ���R�V~n"�0:!��Ҭ%�(��}�pNe���o��#%���L~ �5j��wPωKx!����S�>D
=�~�ɓZ*/�4Y�!q��h�;��]\<Z� �C,��3�=kM��;����IvX���1�Q8�.����s�l�!�R�� U��~e�}�)�=�'���n늬�U'<DH�������0 �teN��L11�yh����ٚu uƺc?(��$b4+��qj��C0&;ڋ�N�_���U�F�-�4��晽s*(qŦ��$/��J���������r��3�6���m���i�c��yk�o��3������#���x�Io�U�@�;�ʅ<B���C�;���R�!���=���-�@�9t�J�|���\��N�b�.�ϥ%�I�ŗ��!(Z������e&�Y�Ƭu���%k�"��9dr-���K��\h�a8{��+�:� �$�?�-��7S����v���=9����*)���&�!��d�1D6����VF�{�+�n
05M�Z5)�0�����&~����A�@{S����r�/�D�����_��ݥQ�R�n�G���Q@�@�m݆��6�q�̀Hhp~�w}b"��,��E�9H���m&�J��pn�Ee�ڦ!ۿ�,��D����7��?�N&KDS�b��ڊ�!D���<Sd�?O{Q,�/	�D�`U5�ݹu� &s�/i�|#d��&��,�l�:�̓<��'�������4��GbX�~z>]X��NX�ܷ���ٚ/���M��ʯ5?	����]V�=��+�������<���ѕ�H��/����<x��hc���RL$�둢�C��6���m�'ܷwM3��)+�r�ѠxkG4�{��4���anw������L�%u�¥�~��v�����c������>�^���a�R���u*ˋ_~4�X;'�]	�>���V���z֏��j��.�-���{+��q�*�{��@QH?,|N��ݛu]��Z%F��8<G��Y��,U^Yܤ�w��=�o���3+�8vFj���I�/%b[eyT���=�����'Pum*,.G{�VÓ9�}�!Z�ধ��EF�z��^���Ɋ���$�^���c����y���x�M+��pг��r�t�C6@�WvN�Bg C��7%��ƪ]ێs�2�2%�V�}�r���7:�hק1\�\�yaGJK������D?���T��9΀�k<��Vݒc%��q6ίX�X("F�3 �N~�3�Sq�p��z�	H�zv�"� I�T�Cb%��+^�N��C<(�9�K�mԺ��y�Bh|����.�PM���K�Un[.�#v��"����
)�@�X�P;!���:�A|�P!����M-���������_kiI��:=^9��?Q %��T�X� �㣖Z�W(�o;�r�u��A!�Z%��%�l����+pK�f�ݨ#�������pɓ�8�DI�!'!"x���v���gʅ���j#��I!gP%j��T���/�sS��dC�Y�J��?�~��9��o�(�j<%�+�
��:%I��벊ۇ�dH��,�����dD�=Ȗ�7���1hI�7O��]LB�Ie��|gq4�[�n�������i, �#�ު�ǒ ����9�ob�v�����P�-���9"O��R�g2�F��}e����2U���s��y���#`dۏ�`f�)���:�Zo�u��L�q��y�j5���T�!<�K\����<��%ĒBF�0	���)RU��`$�(ބĖ)�d=�y�؍�i���2����x����+� ���|R�qn�Uc\�����2~�]�h��n0�
��S��H���Җ��`�-�ׄ_��Ve^Kݦ�]��S'�3��N��Z�9��ga�{�U�P�T�A�*s>���j���&��ȼ`a��c���r��ِ��cR�z��j�Rz������ƖY�4�]��<s�����<��jJ7�9�S�b@Wj��}�4P��y�a�9��KGWV�[S��ą@L�������hlO������\<���Y䣷��؍qi:��̟����0���n��G-��M2l+@S�1hh��g���C�{�"b[��U���1W$h����;ً�1~���Y;h�m�)�LZ��,�r�m\��½r.�S���pX���z;���.x��`x���n���M�U�V	��� b���3�tzЎE������@���
��S I����H�`��b�`LϜ��t��h�h��S��|BC�.o��X�Н!�ڦ������:��xl6C��|m�J ��[������o�*�oT��^�s�b��
�oA�����.)�S㾚���{�CN�@�3�zΜ ���@# �W��)ªRlޟ8G��9��������v�%����ɎZW���J�����9%Zq�����)`F$v�ɸ���O���s�-߼��^K�~�DS�
������'�}#Ѓ��D}������'�Qa���` u�yG�V��(�v�) k�J�:`6���Ȫ����e�b������ܿ��^E�7=�f