��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�]d�L=3	w5��?�N��A-�5�P����B�[���훋�^b�sG(�dt�.KR��:z��X�X�8,E��c��DA��G���\�9��=�����*z?��'�]?�VUv�.���Ԩ0���L�sB�Ξ�U;�[�B����gM�1�·܅�̵�$����Q��^����W�M5�}�<`}�]مڦx�|KW��(`G=2[�'J��m����5�E�0�d�ܩT�I�f�[9���wt��f>�eo��k��F�����Z�jz1���(�+־876�����O��|"��Y݄v ��#�<�;�dWZ3wP��3�Λ�v����6ě�M6Ш]� �ಳ \��+��1��U������
����$8b� 0h�H%˂��>�cxf�T=qE�Dʱy�B���	��cS��4���f#�7�dd%�z׾h/�=G,�C��O�gq���}m��Z������\s�B��H)R�:�)7^>&%b�D:��\�`�6��H1�M��d�5H�[(�|�w ��m�����<g���eb��M0xc�b�:mQ���=�[�ٔ�"�� [D���9��(L[4Du�jP�b�A+��AJ��Jr����%S��:)w9p�t�U�.�6� 7��Gt�����r7&�q���8��1��:�4Z)Tj1����V�k]S��1t6r o�T��m�c�>MZ˪n���sN	D��'�It�����qp�'��#���TLQc�vм��M߂���P��<�l`碘ӯ�h�% "�z�'1�G��*��d�p֖�n`�/q=��S�b�Se�U-����v-���qG����a���oO(7��H�����y�v.P(s��i�C����<���}3M�a�FXCz���^
������U��|��
EH�h�$$	~��Xֵ���jYK��k��qͥ3��!:nS`�@�a}�H�`*�<�H�$�).$�P�Mtd�~9({ Ea��	�g�z��|E��ܶ�
"�D>�#H��N�db�:�����M֡��za��yN�)a��Tf�#���#�F]�B��ث�
p(�N.����P�+��K���{�_B�ޑ��䛹�>�=�z7�8�l�Ur.��ӭ۱�g,b_����:�G���*Ŗ
6�!�e�P8�G�����Ð�E8|
�� B��{������ !U_�5�ڜ��?_;�о9��ozIY�0bP"����\�^?"���M�������^y��G��妻pU�/Oٟ�H6�`�?�>
�c�h^%4�ｈ�kU('J�a�{�>|K����%?��g��R�k���Wt�K�A	i��Y���3��&�I�R
:���R3�����(6#��ML_�b���	xZ�|3Ǯ��9e<���Ip�,Hz, {��Y����n{|����@o����`q�Q��1
�Z�x��h��)<%{�sQA���t��B]���:�?B*%��v���e�C#r�K�|����$��B}��4J�XA<G��Raח�VAe��d��l]J����jD���|���쉭�Ϧ  ��
 2�w��<�����]��Bnc��J�9����( ����QA=it^���̽�l�%��LK'��h�lh�X��`BEe��j�� ��6!�q��b�%��L+�L�A����8��*�D���E.�%z߶�a�e�l̝�S��ҍ ���^���1�m �Z�[�S_��4��t0)㮖��3K��$(����7��T�b�����I2���A�WɲU��BMyU^9�u�/u�L.Y�F����.P��$/	�3yx8C�a :�䰦;���O�X�\҄�ae�s�a	;gQ�~/5� 4�US���p?��e�_%��st�%�p5�籄hN�EN�)_���
�3r�Й;P&F�b3tnL�-�O�_i�����5��p�E}�k� ��8�OI��I7H��(����H݃�S���;�w��"�:׵pi(������I��x]��=�}#8Ȕ���Y��ף�L٥c�3I�Ù+�/��ݫ~.x̨0#%�`��k���<����f�������hm������b��r�w�u}�W�����8�y�G�P��_u=)бV� %��I�}č;�4��l-���g�r.�Z^/݂��;ʟ�ȃ������e.��v���pz� z�7�ȪߧRt����`k��G	)�ۂ/�5��R��)8�%��Z�B�ѵYkZ.z(&������:u�@"E�
�,�)I���3���Ta);�2Ho�1��BR�I
M�[�`A��LN��Х�b���[�=��2�(�憍O�g՘q���z������ �7�NE�������Z���h���>~XO���HFG�~��Dڬ�v��m[ �A��(2��X�� ��,�J�BK���M����yi[���ηCV��.N�c�k�_��tJ!�7,Gjr��G��<�n�U��g$��̈/�m��u	@ݡ� �~v�]J��3!W���i��,߾j�U�i�P�ʪe)=�����`
8WQ�s�<��B��̜�/&�p&9�ǣ-��c,[|��'��'��1��ew���-2:ӂ�����YQ. x���O��Qù_�x����F�ۛ^߳G1��r=�q�Q�cW�X�nuP��.҄OR\8��摺g���b�u��<�p�p�h��WS��gAzN�؁�t�EH\"��4 a%�(��it��w����p{�	���j���nc�0�"= /#��|	f`���^fg�5���7D��@�bS�
D��5��݄G��5�Ȑ�{B.���G��^IQ_�P�`Sۗz�iٓ$�{*"q�ݩ_7~� �R���L
m��_+U�zu��;%vG��:���.��Mx�6�|�S_p4&f��g���`
����ǳ��r�W.�ܝxj�����o,|p�z�@���Ui��}�o�����_������	{����+@��A����p���3ǩ�҄��TOaa�#U�ڕ7��G�3�l��&���H��T���1�@yLウ^e�� T�d�	�g��n�Aj5�2W��Z_t	%�:����*���:��8���1�7�y�2?b-�"�=QCj���ZBj����}�g8xe9Y��H��\�<$79��GM��\$��%A4Pip���H�?iQ_���>{"g�	U�a7���k�p~��2ʁhɎd&�V�s��$���mg:�	p̅��d�dp]D��]�46�;x~g%���0O�[{�"�!�j8���K��BCf]�|(�ar}��lW�VrG�j�#ǉ��O�����>�2LJf��zi �n�Ы��p~;���х�y�ᵎ�	�{���\��p0�\F+�UH����x	[نMk%q|���򳛴^7T����H��yǜ�tC��%'��i�$��m �4bhzD�z�q2@=��ۊM�vA�����_IN�C(��r�8|�n�u|��J �C�%�n\��ՠ.�ԃ��	�-���@��y������A�o���S�;��Z��GF$OU��l��b���h�`��l�Τ�f4H����z\4UW�_�,�`��hB�Sg���ΆGb�s�PHr��#���mmg��˾�30~|�H��Ĺ�FN������g=˗<���J�+��n��s{L���(W�;��;��`�5����v5H%�~W�BFC�]%+b�,�]ʮ_���{X?@�zݐr�����ˇU�����Q�1�;�7X����d�J>�0$�2U�\�ٶ�Td�oU9ME�,��>Zn�޶�=ɡM`vF���W�Y?���:��+�t%2~2�s���"���a���O�5=N��;�^h�]3���-'�J�ջ��</�,���[(l<瞁Uݻc�/=�|B?�eI���\P�� ,�C-�$HAF�Uҏ��p�Y��S��PS�w����o�:q�и�?���'}��$\�g�t,������A�]@�:�Cw-�_J�	r���N�Ԍp�`I��d�$R糖]�H� ��/_0����GOv�=�R53�zb�ٞ�{�g�F$f��Å��F����wq��6̄�h@���c-��Է�Y�1��M�@0!�t'����q�̔�,����YHB*�@u��,���pu� BFt&(���#��ޑ5l�O��(f=�%�>�-��=��r�Š�}I�D`�K��\7{����Xư.��i�p�/)����dd2覐�Y�+�B8�'�Ӫfq�__����n���������,��ر2��/��\<OI��?�J�������):Py:C�n�3/8��c�zc�[Z6R��A�N��	��J�c��/�@�/ٵ�MO7F�1_Zn@�x�d;�X| !o&zĒu9��S��ʪ��6(:�Q�|�����2���T� �y�{W��G�V��l%������V��?a��Gq.à���Y���\�6�����M"��U<<�P�V
�+HLX8����5�����E���x���qRާ��0�:f�6ז�}Hy�B+�> ���d�Y;ǫ������P�E�E�m��Kq�K�\&R�Sne3{B��Bl����7K��m�;�0be6v#E;�W�7H���(BSR����~0��ɀyЃK]��z1�5���N�l-��+����fsO��o�d�(���[E���+���`"��z����[��'i�ϋ3�q��	ӎƹBrI�I:%$��2�4�x�'���JX?q9���n5r/��.�KU���Mc$Am� ;UA>���&�"�'�7;�u�$�zb8����!�u��䊰q.��1��6aM�C�T�}Uh�Z�;��|z����׀mk#�K4���CT �������񸥺�pen?����33��6[�.�f����ҁ_��z�A���6�u��*�?���8@��]̏i�,w��~�s�9%V ��;J�IW��Jbk���
�#'c�N�#<[9+��Uq��Q�M>)�a�Խp��+�����!b�2���۸�-�bZ�W����K�5ꤩ��Tk'�B��T̦r�kin���-�C�;s���� :I�l���u]�t0k$���Rj�HY�<��0����RT�VZ҃SFsu�h"qKt��t�����݆K>���d�"R |?(h�>���f.w��( a?��`u���󔼊��G���zq<�#�#�3���ps�'/�i�[eP����]�a�hK��8ckH�*�Zt�Zݏ������d��!�0����VY����bJL�I�%D%��[}7^�S�&�����1d��Ώb��d��>VP���N�E6�/҅�1��0H{B�*���m�#�ת������l��r2;�I6S���Y�0*��@Y�����]���\�mj �*b-7-��R�*U�l.LA�#k_��jpwP���')��M�ǵ��!����/p8wn]i��o����?���2�9�q8��-(��Y��M����`�����#!Ҳ�?,p����8��/����[��s�8<sĚ�Y�����8k �
D��vE��ʲ�]:�z�%��aq���@&g�Λ�)u����Ȅ��y1�%u#�RN�<n���H��$��C�����+�!*='��sm���P�}Yn��<7��쿣��.o���nq�����Z�}�-�Vt���6DAx(6�������o� �9�/NI\�|4�ȶWe^��w	���X�ψƞ�eUi331�Jeb��5�p0e�P�Ӈ[@�������"�
�	��#��8�w�?ؘ�����Y3���db�wb�d��tb�R��b���bx����y��I�H�Q"�ii�pv��v� ��6ic�Iw�1e�>��d���p����r���b�n�����#���|YI9�qԃH%ք������6z��Գ��R?샕�{�9+P"/&-M��z���.���ͫV�Ѩ G�S�K��ӑA���Q�X��Z��l�=�>x�e���G��A,^�����|
ib�qq�'�4��ރMk�:���.�kz����n�B0�X�A@��r#s퇧t��y��$N�)���T,��/_�'�G�4��v
��x&���9��G�Aؙ�/�U�_�w�͎�e;>�ȥ��8'���?��{x�UwAR��|U�l9Q�C�JgAݻ�����|!Yfk�:;����b�ヵ@Q�`Ƭ�f-o)q����{����Ž�|j'be��E�-������Y��%]��X��n�Q��o�v�?�OG�K�_ZJقA����j����p�l�PS�"2!�$���.|��x�����kЯ�����Y$4)�C���1�UxW���]]<���v��e�:ڻ2a)��1���Y�tA�X8X���ƫ��]��}�z��W���ys���R�i���Ƈ��+�:GkVfơ�If�K,&-�LU�!�M��"�����(���6���� U���F�0����ϒ3�3l���>hƁG�m���$!�!s��7��B��:��37�	Rif�z�I�ɬ���`���֡.�p4�\-�(,(pri�G�-C�%U�7GU�;q6��B|{01�`s4G�DV���a����%��m�)�ȝ�'^��������w���&��I�����ة����q�-4�HǤ2���M��f߱�ǔT��P���G�6fw_�\�HbC��`T�����3�E>�]a�Kٝ��ʛ(��aZUh�y6ᩀz;��}@ϒ���s
�����4{������Y��#C$^ۧk�|���Gd�=�%]�ה���w�(�D�G�9g{�1�2I��,k-w� Ϡa��KvͲӸ�>�),��ᩉJZ�ڴ
����c�-a`��c��0�u�L��y�1PPc��?�x<'|r>�GJ*��i�'�{~��-�~��+�<f�V��ǐzM>+ 5�`���)���h�R��; �X��Sg.��X�����]��c�&wv2�gsV:��U~�񭜪�`�I_��n�w�TA��`��v/ߟ5�u@�:н���������9�Ϝ���s[ŵR��5�����{���c� �k�����/��OӮ�yM�B�UQT4�2WK��m�
��Ѓgb>C�ob������� 8
�w���R�Z�?i��}���'�Z��>Ɓ�9�Ѐ_:0/�5�s�a(��Atg;���G�D�@7J�(�^4�^��A��s�g?Ճ�<LQ�%�^�V�a���V���m5����!�4qF�_�^ �nS-�-fiR��u.�|��נ����u��<����J�GBg-(�I�p*�{��[+?�0i-@���$�7Y�x\Ȭ�r�U���:`/�}/@���0G�lg�.�v�o���z՛CI�IaV�=�eH$�i���	�d�!$��ǜ0E,6;UIj�&��lN���x0r~�
��}���C��O�s!\p]��0�P����.a�`c�|s�1!W*�)}_��ś#d��ާ[tB�Z*���)��_7����)D�cD���G���������3��o�<�����޵6|=�e��%��θ@�D�;_T���ܐT3��ւ��5�Y�+�'�5�Y���)�������O!ۃ_��S��K@5�r���l���
f���{3�z����esP~�R�d�-�7#��$=-*.�@��[��T5#����)�Ě`�Pٹ���-�;�HV��
.Rϴ�	K���JHx{Ɗ�ꊅS��G	�h���@�6�ٯ��}�NO�un����0s��.)Ƒy���(;��h;Ѻ�`9��[a���F�J��,�cB�����UL'����;s�b�����k�|F�/�Y�N���R�̆m�e ���4M����qc�^_L��j�$K��Q��`��(^�%m�f�j�s����q�\7�U�T����!d�j��Z�������3�ҜMޫ�5l	��v:�q
q��"T�`����eq[k����b�G,�d���(�;~�k ����UL/��@��g��u��rZ�@dX[65�u@H����vܔ���^������7*��0J8���A	����V_@5�X@�/�?�UC�+�@B3<���p!�i���[Q�{5�?�)�Q4z��`)��