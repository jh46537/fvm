��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�6Jr�����/
#����������!ώie���c��S�ѩ'���ƛ�#i�
��	F�L(D�}�|	�{����j��dP��G4/��~�`�E�	k��x9j$��0��0�Ee��f�<���L����٫�����8��b%���*D���3�h�T�5�P ���P��L�� +5��~(�M@6�!ݥ*�:��|���8��Iگr�g���>�o��ga�� b�,��Z<!v��uW��!b�!��̉��	̙yQ7l�Y����Y6@s�����v��;/���v[\�NC��@K��2�ˮ�3��tc3&��{��WJ��8a��
����{n�DY0��K��sq0=v�P&9ƣ�D/� �a
e��N�Qϛ% ���@�^�+������M6�{����E��d�L���aJ�����`�|7���,a�ފ�Ps6]�*���.�`�C6�3�������	�m7�{uS�]���AW�>��&'����wP�H_��xv\�]a��=�[�}֭¬�{�H{s���nU��c������ѕ���g/�&}�(O��v'��~~�Eb�O�l���MȠr}-�
*���|ƹ����+^�n��C� /�taL��NԂ���|�|Y�ِ�8���Ɛ����y*��'Ǳ��>���s kYF����q�1�뱒���)_���S��,�I5�����{�e�x��e�����c���'�JPq���v
ͅ�+4m)�K%3�r�E�74F�H�dt�??!1���&���~a�SR���U�9[)�0�)�V�ř'��yhwg���p�C�5|'�Nj$����ZL�r�|���AqgI6��Y�,Q;U�N����_m�-y��l���ppL8م�B��L�N��������z���D2����E��G�m��¯i;���g���O��r��i��L�k:�߭޼H�nJ���IJ�v�щS���:��%"��&�<M��q�Z�*��<|L�ݟk|��Gكȹp�P�4ԓk��*�����8�Pn	��*3�ͻ��J�\���Dn��J�ս$ƚLӟe��c��Q��6�]�6H� )�'����W*�� �*+�CJ�C*�&�N �_u]���^�d�R7Tj�;!T�W�=v#1��
$��'�&Z�܀�����Y���2��Ϋ8?
��q�ډfM	sg�F�`��1w1�K��C"����
r��^��G~��ĩiO�P��ME���i�҄�e�j�����7k�)pm�o�)��SL'��딝�3#T�����}N�!�����M��{��C��-U�~�b�_DK�6������&Lɟ�R�9�y3Rl��	B�r�;1�Y� �@��Wc^mH�\n�Ò��/��5[d��N�F��
�ݵRDS�c_WaQ�r��Y͍���z��_H&����
:��F�8��j�%���n5"�XH�=i}�Z&YT'r�IV�b��AV�� ��h�����(�wZƲ��P'��@u�������x�/�����ZFtQH�қu�d�i�=����:tU���jx}Z�A]�c�[&�¾��ELL,n��:j�0�$]֪_|�vK�x�s��`P���
�Rم�M& ����7�� p��Y��%�n���Z!K@�X*Y��o��~)��8�6%��f>��^>�g���/1�*��_���aS�(@e�ŗ��ۉ퀶��rx�r��Ss]�	u�~� 9ŗ	?�.�mR��|���9ĊC�l��ȫE�N��'�7L�}����p	�����q��̇Z�� `����������jt&e6��{�mɒ'l�xR�f�#���Ť����K�ykɳ�#C�"#��M��11��j���9`��Пa+B��t6e��5���\�(5�j��𘛸!���s��F�4aS��x����)�l	���T�����`�%�S|���5>�,���Ͼ��Zw��C�^.��Q"��A1b��1��Wڿ�x���P{^OD��D��ƛ�r�n\����[���"O6� ���D>WU��4�^��IY��t�s
��Rx���8�ZF	���o^3LHT�NCl���O�V>xU��y��m�	� {ۛOJ�E[pr�U�y�0G]IopDt]%T�?d!�����'�9�8vɲ�r�7dD���N�-˺K�.Qv���=���]�]^0«h}]̅X�ˈ��17<�KE�y�w�\�w�$��0���Y2[����h�,�k=�~�-�8L�7�C�w���2����mCo�cB�����+��1t$� ���R���<���:x�`x�D/�s����^��k:w)��@���	�O�w����kنȃ�������&CC���Gy�4�j
S�c�9mKv*|TUƺ�I���U�=��z���ւ�S������gQ�}�.�y@�9h�j�0)0�UK�H���+�h��\7�'���/��_Q`Aau�p[W @����� �L��t��.�8���W/�Gq'r� ���Bg���b^i��
�����~Q=�M�� Y$�2��^ޢN�eŻ3)���#]v��GM'{��8�Y��\�����w���?���k��e �2H�X�r	�`��TUs�.G�ZuW�ȴ�fm�1����,h;/e΢8��Ē=q����TB�KP�p��(���Ee٦��L�=�S��Gi�`����JX���N߽٤���G}�bX�ZB���$Q<�vF��*3� �I�E �G=_RAҗ9Μ�3"�����5J�cd!�*x> K\��aϰ�/'�_'B�x�PIlu�C��x�g�0��l k7I��|�8_�{?Ԧ�@�R2�.v/$$��	�#�uV����EYp��a4�~'��{;k<ɹ/�����/7ߒ0�Z+�ۜ~�Q7*�����o["��/v���8��`�UE�YK���-s9��&�1+���U�=��M�)��=!U��ns�hT�\�Mʻ|s�s=��5��,�o��.c�6:v�>m-6,�$J����.y6t*�h���|��:,@h�
�C���^������xZ���H�ʙ���:�� Z�ZZ�qy�n-M"K��4- ���͆��wV��?ȱhZ�,x|����"l³|
P�<]$F�%5w���5Oc�����$	�������2sK���EN�w�.�@��Q���d�Y#�q����&��TSƘ�a��F׹Zo';��<ѣFK�,�C�w8�t� �wk�� �d�{gZ�����������}b������i\���BR݂�����(}�S�>�=A��k��Z1���:��"�+fb)&�������Q&�6ٯbh�f