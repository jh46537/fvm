��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{��*�u���8�R�� A��R�:�@�b�ˍ�#�)AӦ��OwЪ�ۘ}�6V��;ɟ�I�j�8A���WA*�/2��WC��%:/�/0'?�xg�{�E��P���<���_��)����)d��y�W��{9Y��p3�[�A�+��P�>ئ� ��>�j^	G�pԪ0��!~����Ξ�J<�Ŀ#�K�L'R�>��H�g��E��ϥ���$�	�/v,HCg(��X��8�r����Z�r�+�/����D�/�����In�a.rpȟ��v����=���W�?��y�p��׼� �/ڒ"�ܮ�rZ��Z��@�vT�ԛZ�NdL'D�:�%JEm�5r�y8��b�_��cH�#�Wr�=�YC,����RbEֶ���=���,�ZL`�.�y/��#�	��'�Q4�yo��*��_M�l�-#�!ҐDd68��f��|�ۖ����>-T�:���Y�����U�H��rA���6�0R>�é���e4����'�n�r�]�5^@�ڙ��S�ر?�;�;�ا296�;�l��
`�����F��8(�E����3���1�(���+���ݝ��i��vHb����������@��[�#2@ɔ�1������p��3򫪲ѓ�YR,7!��@�K���ndC�����T���?
�X���C[h��L�,M��D��pLÐj�u���ΜƵ3KU8n��Bo�c|N�CsS�����T��J�]�c����~��J9Z��*���=��da���XB��4=��p;�� ��B�.ф��	�ڋ;��;�%�EB���g�
�!�^�>Y�Y9��1m�{�+_С���j=���aY�T �\m�|b�?���}+*��6�]��o��ԥyIQ�!�Ga��7��%;�mӋ'!Qwl;�ᥨS�?��{u��i����w�6"T��#�X�}���VK�%b/�8��X0�tha��$y��7��M��5A��~������LZQ�6�fCH���n�BQȣU�ؗ�.i�N];F*��o��������j6X��C�� J���p� ���N��;���8�O%30�9�".iB�? <x�`I��MҊb�~��6CȈ�ae�R��N��N{��"�,�֤s�-��/��i{��#`��H��e�)wm�0r)�i�J����;h��D�X���Mo����?O����)�˳qCׇ}�9�Ro%*���c˥�~�[�C�/e�ٜ
_�����B̝������%���^�Y]���?EhfvW+ɯ�i���3���>�čϲ���'0���E:����Jj��-[]��	�Ly3�w�@�a�Y��p]b/�>�e��n����5ھ3˲�}z�h���I����ޢI��j�@;ʊ^!����2Ί �:ć���FV��׿F��n����K����-�`[!)�t���bU����`)�����iڍ�,�Z�^�V
.o� ���5��3ܦ́�t; �M'BH�7���7��!$z7�r�ȝ�uQd�z|I~q/Qf�4�z\�V>�Y�I��Q̥�a/����9��..~Y���&B:��T(�Q���ѼśQs3��[��#ޕ�Nt`W��%���y_�qv�b��+���5M.��L�A%�?p�}��3��F�F귆�d/rJ��;ょ���������<�5��2@�S�o$"p7�j Y�qx*'���;E���|�H�v��:���M��L�4�}:i˂&<��9�Ψp&�г��.}������n}�[}dz����W�A�����'�詒X��3N�>������`�b[����N�P%��-��g��i��@�0�;9Z�����*�M�p!y"v>rgj����~5�dGlN�6�	�_�`�W���G8�θ��j=�}A��U�.����%��[KfٽFeRԃ&��YŌ�����`��PwF�"X�2�Md�x��8�ȟ�S->4�,�F"�����G����e�O�J�֭U�{��p��Y}(�o��zw��}s��9�s���~�I�9�,t�� �J���UX�c &�����.G��t�� {۵|��~֐_	-�L�%]�+1�y?��5w
���hG�P�Ҧ
�4I _��0�ˊ�9�-ֻ����L]JT��G6`����vL�������b����о�6��Ku,�Ҭc�u��F�y�Rq�s@�
�4��!M��s%3�,��#e�Ah��ް�d��0S��Ƈ2�������k)V��Ұ͊w'+����♲E|ճ8:@����� /(]s�c�l��Yp��>y.ӵw ��_y�aI��k����4�ɣ��>��Ϻ�����)( æ��傂C(�dv�Ǆc��5�C�-^6��xS�?/>�k,j�ᑫn��z�y�\aj�(��7���&���_�8�n��SY0��hI��T�zۀ��P�oB<����#Y�̦�p�^;��C���;Xt�?����1NAD`��=؈����5�Y푭�8�+�uY�8=�⨣�Fֆ�j�*�d�踇�u���_&����ͽC`Q⛆���N��@>�m��u-�N�v�>(�zW�æ;v�I$����3Nh� �ol2���� ��i#v�.0d�'�<ɳ�c����p[c���C�'�ښ.}Q�\8��<c�^s"NH�۽~�r�%���q|�j�$ޣ��L�H��2�9z���½Xړ��UWt��(�M_@D��n�*���+x<�=B��e��傮3g�+9�&�� #��@|[�ƪ�g��y���d:�x�Ws��º�<1������(":׭�E�Hb���1��|N��M�y����Z���나[~�p�=���G�V�@�@���C�*Q^�&��VzK����^_1px}���=�H'�Rl�%���T��khL�2+]0�T��r�>٨�����hLw�n~n!�t�P�T��Ip�ծ�|`2��п%�4S��	eԆ<⳰����4�[��|�	.V���YU��b�@VN`�H%�xp��g��wt%N%m��J%�];Tg:������VsH9�)[SC�ȴRE�u��v�O�VpVp
�����O�Iv�(&��]�A$tew�k@3TX?4=�Y�E3�i��q�&oIB0�Kw���ΔR}��d�{�&P&��uQ�A� ��B�ᜀRHa�"-^ �Q���!���¡g[��2��X\����2�X#1�X�"9�V����*@g�s����-y��e���+���Mm��X��n\��7���ۨc6�>a&R"5��@e�*�[���
���|�^�9��
���-�s:��Qi����c�O+�th?[�-�t�}��Ň�W`�!�Jw ���L@�>ϫ��X�Y�y.����Hb�+�X��Z�W��R�JA���؇�&͛�i��	���N)�e�;$�k<������`I����J���-�y.o��n=���޼J�,E�~�ف���͹'�/K,j1��,�W�)4���Jz0�W�`b�6�p�䌢�I��֢i�>�
��w�R�q��j�Q���n����	���G�2F|c�"�s蕝�Yb|�ͱiw_��%��L����q�'��@h������`���cyCΆ2i���1��Ŗ6C�cj/GIj0�-��1�yt�a����8������<�[�،^T�xZK�:�{FĶMa�+LĨtAy$�^ցj1.7�ʥ��N���rS�f;�0�{�v`lho����][j� ����~Ia��b,Jbýb>F��_�#@NI@̾�:Id�1'�)�F?�=X>�a��`*����:S齯�3e{�͟��YڸW��v�C���t&�r���m���>�[�p��ӠB��)�Գp"�:�o�*�d�6�#`/��S����n�n\
ն�����%��N:��$�k~{���4��F=�:��p�.�L��j�������D��k��:λ��^5���c7�/̳�axڢo+�O`���`��d��������8=ѽ蚜�auRC9��y��K��"<��.2,�����37�ϥx3�m��J�m�D���v�ߺ��e��K��zL�k< �,3V��e��t�?�̄��Z�u]�D<:���2a�8�!�v9�֢�eS�N-ݲh��c�%ITK��M.�~`�#���Ag�����ˆc����������N�\�"��<����|�DW���̿�!��u_���̵�|͖��2��>rm�c�(���u�v!}��^_3Lۊ�-�i���G�h@*�ӊ^}�($���q:u�Z�A�r�:K��ټ��gͫo������k�~��(<z넿?'����m{9��I�i� �T�X:�[4��~j;
�0Ȫ#7�R���`�hqqD8~�U:т95"G�{�π~5���S�Pf�º��i6��OV���b�U�A��h�>����.ĐI�P�?�8�0�3���U(���
S_�40!����
X�N�L��&������l�@
�����f�!�Z��l(s�!=������!żZ�e�����*ebk���!�A�ӊo�j]��r/'S_[��GjYz�|K�8�+k�#΅�s;�>sߚ��;��.���}�_��ëC�C��K�[�|T�f���?���3D�$i	q���
A���x�7��qMȡvU57�:z�s2>�z�@W�&p�u��J�L82�,�--���;����o�nפ�܆��l�^^K�>���]v(Z]F���5���4��F��Ͷٰݼ��@����p��7�o[���2��7��#�L�x)G1�'��BeeaR�F���āT������ր�[���\'���K,u�Sz�̧O(s��wa8E�|�z����`.`[d�H��q��ӕwz⨝�#�_O2�c�Wig#�֟S�F:T+���05D�=��!T#T�*E`y�y�j�n��[VUr�3F�3챳&�w1EA5Ă4�*ה�v8ӡ�p�
��7er�حT�y}* 6SV2����J�tҽ����H_�<�\*o����/A�K�\���W�հ"�J>r�ի0��O��}j[�ץO� zƟ��ǂ����T�ذ�d�)A���ŅgBcc��ة�<���H��,-n��9m-~De�|�}��J��˼jO,��:��Q��Mqch��(x����.��T�MQaTI�t.s*�3p��U�m�S����mcҟ6�O�Lg���˸�y7Y	G��{���G Bں����9D_�̹mH�%q�;&m�,Mj�8%r�@;���y}arj��n��0�rB��(�8���`W�F^�K�w%c��rRlU�Ofv-�&y�N�ڒ���J�.�΍I�J�'�����T�c1>�:�=��*q���^��s��&��.r
��l�0�,`1�`G�:�n�9)�M|t*_�R�8� F0t3�ƹ��=b��8v��x�[p�X
�����^�b)w����m�a�,P<���J�(C�.��v}�JwE?eKt�֖���y+/OYt��a�OW�;���K�\q���f)�m�,ׁ���f,��!�v���5��e	�6��pqK#�&.̟����؜wq�4�O'Sʣa��$�q��k��f��DT֚ ��w�*A��@RN���NI	x�-�V/����v�6��}��k��ϰ;���u����r������|�<">J�_�;I���!&%�K��=���е��$.���!���}�O3 ��f���d�O�;5BS����BE<��%Q