��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~3��Z�������# ��d|��̪�����PAZ:�;� ��Փ�?�}�F�ԙm�-r)��]���m�V[��zA�?�p�,O�?����5���dk�������'�]��i!������&5E��PN=����x��ҤLh��c9�`���u�˄x�]�-S���)��q�(��EJV��ϲ���rb,�RsW����g�.��6+|�{@z��'�V&�.�@q���K��&���x�:ãp��h���D�$ޛP�\�ljD,�>���]z�4ׅvQK$L�<��y��%�*����E^p�ݱ4|����QB�h	ce�dL�F��I�0԰�Y �#ѱ��uK���}h��q̔kJ���̮��v���5lq����>��4�Ñ�F�	 2�� ~=-o�U�/H�g�_�;�'� ��3�&��a(`?G��w\r�BR73?���N�����輠r#�\�;"a��r����3���&�QP;���u�e����{{䩆9D���&��H�KW�Q\��d>ǥ�q�WoA�B,��
}��{�[�Y��A��k�j>��t�����N����4F��h�,̖�����ၠu��=�(b�_�)�Hí���K�Ng>Tw�iT��H��!n\��x>�OY��)LJ�!����>�p��@/O����� �M�Z��!�m������V����:-����*y�Y)�� i?ͺ�i�����$`�� �M�梨��Җ_��BQ�YlK6>��81��/�Eh�Y�T1*�{&.��	+�BO[���PNa�ȹ���C|!�ݶq~�c���4Q4b�?�j�oRT%Ӄ!���z�n�,��;iXXn��	�twx:3V7�[h�>���v3�10��+1y?�~�)���pJ������t2q���&/wN�c�0���cS>�c7��ͯ����}�L��%��Ų�V6�b4J@����n/�%�@����yh���a��l�h��Y�ڜ��ǈs�qT瞤�9�<�\f�����ɡ��\i�n�M߼�C�}��ӓPi�
���S��D��R.��f<xD��%i�7X�\%0I(+���!q��MI^?7�vmh5�*��tlZk&~u�tK�Rx��6{��~��y[�rq{I�	7ך��.bs/��ȄD��& �ʰpISb��Ԡ�~Y��cS��R�)����u����ϱ�Ն�s�8[��}T=?�&�L����9�H�to�i�j�-R�KE�ՠMFsB{O�@�`G���&�ѕ���yB�C��9�j܍���n/��z��F�DŴ�%���	#g�.�u��`��?'~TCl��~,���֏>���ȮL��=}(��\���E��K�!"�Lm��K����Bta�����X�bx䜢�i����S���m%���O�qO�J�v��`�gL-��d&rt�{[�^�Y+���34FK�i���c`>�	3��������| ��J��}[E�}<"!�L��U`͎�����<jq�b��fPj�/��ь�-�A^&�b#=�uS0+���+��aU��
����&`M,��,lsyX���ͯ*�o.���x�\Get���>�n�3�)rK�y��w��	o�Q�����7�$���m��ۚYg��(5���6j0�h���=g�/��!��g��X!i��!$d���y���B���*�%-GԼ�֬��V$�]��g{�gx� ����_����4��}�|�˼�3�P�;�zQuek����)bͥ�sP��j!����"
��o{b�G��r:�qZ<�j��(�	�� P�`�ݚ�B�I�YJ��2�����p���?1������.i�8^�}�i��
f-��ڤ;Lpӭ��u=�(p�Y�?3�XJg��n�6�1:����yL�nŰ״E�"�_��ʷtsc�f/�!��B��Wb,��,�ǒSx�D�/�K$��NOH�U���ov���ɚ�gr-�!��W65 S���ɓFt��p��!��LY� S��ի�}�~�}��@��ؠ����ٯ�0�ش���rEP��7p��܇�N��=��sk�0�.�X�h�hzI��/�T����ODPC�&d�E;�~S�y���`<���a����{��^�&�~8)T&9���O~~���Q��k>]/�m�ͨ��Wrj`P�c}j`��y!A��`��٣���Y1}�����Y�gb^�� x�+w�u��Uǭ<��.���s8����vO DT�S�RVU���!z����\�����L�㈳��/��3X���1�=�M���bذ���ћԱ��6P��;��Ӝ��~W��ͅ���	cO����z��q/]��	��ƶc�r�k���F������jD��l؊q8:�:σ5�A�W��W�@�v"vȮ�̦}E<L��"�-��i,�-Mڝ�����	W=���⩶*��~���)�`8c����G�4����=�خ��[���7Q�"S׃�~�Jq�@Po���f���~�$���ƀ�MF�V��H��/�������\�y�l)|�&T"/rr�2)�ʍsZ��Q\V�DP���Y��x���͓�YUU�������<��a��9=N(��fe�(	{��ˡg�qA��iу3o��N;�a?9C�}�]{W����b���S��c�uGn����$�W"�2��U1ģK���_Wi��'$�G���II
`�/U�������f���PI�ڨb0�#��'r )�k����Ƨ��1��>�W�&(:U�iv�qm��{�].�Ks8غ��+-�r ��I�N�ӈ�h'���"K7�$mb#*��9� x��?��O��r��h��qY���)�/�*iT�g�� V~���/ ���ܬ	՜1D1du��|��|x�3��T��Wxڡ'`�8-�lH�G�e�VR��$j
x�B��pE��t��o.S��U������,Czf�-�?5?&�I#B�)��/�4nb��
�AI���V��ti�i�W@��c,����K�	
�7���k�g���8���hI�i�Rb�M*�i^�B_X�&w�z찚	p1.H�=~����/>N�jRK$%�k�2�e����m�@)Ȕ�_q񮟸�鮆���ڱڔ[�p(�嗶G�]�Ԙ�tg�Bv��+�6`BX ��bk����ݳL�#����D� N�f�]r�հkxA����P0:�U���%Rr�R��"�m�͗������64�!�iz��U"L�!xtIQ��^̯�d��"�68�����1ad#*귁̃}tHK�ڝ<�����p]!7 �\K3�ODEU�W=g���`���ް�;:�r��K��YU�k�v�k�+G�P��BV�T�i+-�Բ�c�B�h_�ٴ���}D��][ے��L7���z��\��;�%���΍�[�T����'��d��I"��K�gZ�ѲT8�W��v.jY�ֵ`Ұ��6�E��!ʝ��z��]�<eפӊ��Z ,b즸��ơY���"�-9{�/ -�Dᡕ��z��ڰkl�9Lw/м���� R+�j{4�~���:7�f����@�Z�ޮ[�}�9�q���s����`^w��������6,�z�缛��K� �����J5#B��Q��8noL]����&������U���*ϴlGKo�M
��S4�e���\X�m��A�/q?����p�?znb��4���u�8jV).�ܟR{���=�%/ۀ4o��a�i�O��iV\�{zRtQ`����3��a�:t��W;��3��g}�Y6&�2B�m.  �o�C�������oSD��qRa
�x���N>�����s_�QC���Ör��î7GQ�v�!�Sϱ�&�\ԍA�m|��1f�I����t�D��VI�q*�=����66l��`k�P1�&4�8�`o$�_V�
|�A�g��+E��������[!����GR����	4�+W�v�}����'q����ng���1�Hߑ9�U"c0H8�M�j�27��@������L��z��4K)��d|N�H��#;��A�m`��L^ �4�M5c΍������zg��D�!n�~ݓ?UV�3
�t;'q��@��C4�
D%f���e�&���`o[�;{Sǘ�8{ь���;� �iA\}T�T#�Ŝ��;�*6L�գԴ�Ԝ�� ����eXt�I��&sA�rd%x�KM;3��z֧���ː�<5!�0��79����8���>6M~��-%����n2�/��z���kp�?�������!���x��~��VH����KSs�B�bHf�*^Io*p=2�`!�\?���,���ALm�"����Ɉ�7I�\���Z�NZ�$EC��w�� �c�85��h^m�f�9P@#��/�%밋��fu��>��������!hG��ugtƿ�
8;��31cu��}���e#��.�6�Q�p�ѧ�3yyX��<4��5i�W"Mn∷��������Q0f�\u�NZ�]^P�6�'m�}c-���%�F(S��� ��Yγ/���S��"U!�̺�L��M�u�XO7p��-�"�y>�>Mp��|�%$ta}�-�a2.��10�Q��dQV%e�a�Bı˃D���{�D��m�$�DZ!��p�򜖜e�1�z�iǒP��c��yY��*L��h!��ֵ����g$\���7.("�����!�cZ�p������*@O�32l5�2����dG��nѤ}��kxq,4�(�zmY����2���o���ӝ�bR%��5�����7���}�L�$u����c������XD5��P�䜙��?{@#����=��I��a��g�&��>�����V��3uo$���4�P���Z��i�6�Y�=g}��-\B�4}Pۚ��m�3L`~�H7���$�~|��ݝ?�7�b�By��J�l����P���4�e�NvyO7��)�kb�-�(�W׶���� �{0EW��� XJ�� �LY(3�^�_��>cc��c-�(��#��#�~�v���ڜ�I�8����I-�O��U��Qk̻j��4���9~��^~�4�@�=L��%�
��gUҘ%�E��m���1��K����s��Y5_h�	��t�yK�mm��q+�t�g��	#��>{
	�J#��:C�+�L$�XL�TJısM^C�ԓy�`|�W4\S��bi�9 ���	x� �V���!ᐛI�KT%�����-NdS���J��U�Cei7O�&�� 3�wŪ�
�)4�B��a���BPR�S��w���Fz��X���JC�)�v���M�=�#UK��<)E�G�R��:9��͍��H�`���G;���YV�9/�Ճ������z�lGmaZ�_G]�d\T����	5�*�2�õ.*�Y���ȷjd�.����R<k�l��M���f�%�dij��UJ=�c��ű�B�KBB�n
fǉcC��u/�0���'[7��2+G�����\Tr'�P&З��ˣ�U6�J��
��csn�5
����T���V�]Vx=�6��xF�r+���T��`MUI��fI�Sm��M��x��C>�.O�W�k�U�p}��F�C1�(7251)�p2�WM���43͌�ˉ5�^D\yY�v�!U@L����38��(��җ!�C��A,�#c�l��et�"iW^��H�5��G��K�����&yA�\�2K���@I����ζZ�%R��?�=v�zQh�^ E���}���3��-��ۯP"b1Y{�Fg�:�&�9��ܗ<����,(紆��1�~�L��W��n�O�{}��-��s���Ə;ʕ�;m�t���^9v?�<~�Q�S^1�pA���ø�D�o+���u�j��n�#t�)h���C����b;�r�5�u(*d�?�]K5bs�.}���e�ʿaP���dvQט�RW�'�8b�*A�_���t�RS�M�]�n,Ch�
'\�t�շ�l
�zá����i����)D��w|Q"�*�����T?��d��#輗��[:*��(}���-c�5�(-��Z�\g��c=�փ���KM��]J�NdӅ��?��n�$2������n]���t��|�IR�z����5��ݧ���آA�(<��C�u��֫���B<&��IA!�Ã�u�ٻ&��SCQ��%�Aj>�$����mP���l��xP��``7J�wTA���S�	�^b�<qE-i��k^�Z��[	�\�K������1�ݘcj�P��iNK�~*��Щ�H'n�v����}I$OG �"fw�Xti��%���"-S��9�L�DV5�t�MժG9 f�Y���8�\�� ibe�F�r�^WSsb	7���F��-g�h\ϸ����s�����b>�1�c���c^~���r>�¦S��tS���V4������Z���;�rċe6��s)A��g��|�H]�^ayj֝L˴�$��6�����T�-S�� 7M�*iw��2�)����"��#Af�D���D��(r2d�K�5����ہH��/�8��cٓ(�(��3\�X�mٍf���33���*H��06A��ډ�b5b>�s��ܸ��� ���6$�zD"}���+�]�&�AKdb��X�$�,)���Y���.<U�]�޹~����ZB�c�K��|ݏ�G�w��ܨ>��텵�#o����韂aK9�%�CP)m{�����x$� ޤ�1,�
n$/���l_9��")^��$��IK�ΚT�̉C��F�i��X�sC�R,��#9�]WJ�0��q�Na�O&�G���Md��&��7�l��M�?��}��VY��I?���r8��N{G����i��=�:H�j����꒮� �#�9G�����0H��a a	�����ƀp���rChW��״������I���A*�5J�����`��$�(���?j!�xC�7�{�p�w��u{�D��t[�n�̒V���.��'<[�҆Q�a*=
�BP��[�y^��X��{��Cc�[w������+��D�`/>Ye^S���
&��6��$�*3�@�(�V�r&mָ_�r}�(��7C#���wi��2ŀi�n%(��9�'�˩��zS}���ȭ���[l�1�龸��U�cHZ�N�=<��1Ʌ����.k(�>����P�㸈����
R%;�'���	A�VFV��뮑�x���+��_��I�"R����9�/<+8�}ws�$g�ͫG���d�W���C��o�<�����(�np��������[-g���-��{=���E_�3��!��<��Z����2Yŀ��h��G�ڲDQhO��7k�S���=<��A)���")P�M%�3��?�f�;=&5�q)X�S�c��V�ik� �O`i���n���[�4����2�<��F�)�I7�n��(�U�'�\1���?ȥ�u+.���T&gq}�9Ȕ�h*�UQG�撱��}��mbÓ���l��24e�`�x���Gs8��c��`�[��6�KC,x��7��'��C٤_(����\��NkU�2n����*;�YIl��@���a7�7���H[��3h��j~Rn���T�#4�V�ό��O������݉I��ҹ�.���d�c���f2%]6K�?m�Jl^��1�=�\�<:��c}8P�m7�Gh��TSRz���n�!��t���I�m=i�	��t5�N"��WFbjw�\�\���+�	#�LQ1/�����@���_(Yvr���P��]���I����%X=����mS� �!���bMD'mL�W���N)`�R�ʻsa��͵LW���x��H��(i1����$���$���h�.�	�Y�X�k����~�[�.�Վd.����jH83��ݔ�V}`���[���ST���s{�V�#�A�"r_��I�I�MA�p����f�d�a�9�	$>�Z����z�A�YI>v>�]x�_��肺 0��(A�s�&�ũ�꘭a��\"k�x�1@�?&
������2BCBnΏ��z�5��y^$U�*d�W���}+펈��o1��%�x�� ��v WB� \^�� �D�p��.q�6t�V��& S2���d֍{�Vnf���\���9I}I37���8�C�y�$a��Q�����滥p��|كO7��	FU"�0D���&�ӽ1!ڒo�p �*�%}�K�u-%G�'���)�����̤���2��uo�Dڀ�Ca��WX߻EEjqGf��4�tV~���,��~�eh)��vI:�7������vc���FO��p6�a�靝���a��H����
�`�C�Ѐˬ���Q�&ݡLi�]�Цe��§HWg]KVJ� ٽ0�iW���/�݋	���H���WϕK=���nw���4�jnZ߭��<�L���D����a�!Ps�zi������'Ǒg�2пF�ձq:�3�51FA����9'���R�����u�U$AVO��T�Pr������Uj⍮���D���,���3#�����y��Ȣ9i{|�9�s?z�,��w���-�74�M�^���3��Z�ن~#�E�k�N�E��#�23��\7�e�Ph�2>U$jl�7@�u��Q��k���1�w2�Y���kL�m�,2���|UՅ<���SJG����aN�zƼ;�$dOn|[7HlM��AQ0iu������/t��^�p����� ±O���#���2�]�Jh��5�q�s��*&M���VɊ�(}T���!��Ed�h�M���|ȱM-L�Ɋ4� o���"�d����L��G��+��mZ��E�19���=�O`����kA��1��?ܗ\���>#t�L��A(�-Vm�3��1}y�=~��G[n� D�k��Y��>�ӛ`^�4h_ܝfi'��ODo����Z���YVp9` ���s�T�&Lp���1ʫ�.az���B!eȷQ�R�Qգ�$	c��v��fI���<gV �y)�Z�{I}!�=/o�aJ^�D�~��]��������C��8e���*��:$(b@���^�`����x�ԬI���g����/�*�?��v6:>G�d�;��4x�N=�`C��]yh�����MY(��H�^a�P� �"��V:[��)��z�����RDNxZ9�����W�1��P��e0Qx(���[^柼���G��~4i���z�C()��E��pmM���
F���v�ñoCF��}1]��k�x�iO�