��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�>��,�t�Jq�%�qr��A���/4�HRN��Ί��w:p��'�˷34��>,'2��q�B�'�ri�v��B>�k����2(Ahb�I��Z
9�-��I|:$�a�^�^RB������������i3���k�����Ԓ��B1��X�}�%Z����'z�_�x64mhOm~(�� '��U�B3��H��.�6��K]v�(��`ჸ�<D������Ö \��j.o�ShL�v5��SԲ��z�өY߫�%��?�'�����"��@�_���B��
�k�7�S�b#5�	�9��K��b�3��j�BM0� ��@��b"u*C���o�˸�V��v�$���,ް6b�?Ph��lL��5�V��am�!7��!A{؂�ߢ3�"=4�Ct��B�b՜H�+O�X s�ڼ�R�O�Ū��������2�p��>�N$����`n��O�����*F&;�Uo���ʯ@�o8t��ͻ�Ӵ�r�÷�᰸�W�k`���wb!9i�+�J�F.�������&���1c!xCWup�\Mk�&�����"���4��^?� <�r��-�iM���a98�#��5�q�Yl�:q�������2X4�wj��7�ҥA����>:7|�^%fE�*G�WQK0���2m��{�{����z+����Y�5�~�<�d�&mXԀ[Z[%e�㍒�I�0���yXS��c���VJW<sb���Z_rw�fo�������W������cN�8v�ݍ����%�$-j�F>���� x�E�P�J�d<E��
���Nn�1��E���P�+�����=XiU�x��a5���S�;����L�Ȧ����.NH^�����d��b`�Wȥ�4��N�o00�>�(A7�!�O���|g�kb�u���=���Og�e�q��\��!�.%0�s�MըJV�{���pp����O�)��WN�QX��uL��,Jފz]A�:{I��?�
�ެ&�ϡ�/x��d>+	0�P�&��#�j�5�π"�FtF���9�o�蔥n���)O���Mq����f��J_���n�6L|!�02rF�b+��o͡~�$�'Vj�)d�r����HW�M6����;�VN]��!d�6�U�S�G�*�y���tx������V�/�#�t�";ʰ»c��/_X~5�w��M?�3wƀ��ɉقz4WH�����R�[E$򡎒)���U{2S{*�X�Ug>EIT�ь���`��Q������o���J��1c~�m��u�6]^�/+���xb��'(�_Y6���pY�ǎ�!��s��\L��֝E�+�z�D:��̜�(��ʏ�X��2jgS�(7�jD*��n�Xbe� �1�{@��&����<U*�g���'�� ����0]rf��F!%LQ�����#]_����z�D
)�ӵ�e��vF��E?q-���W�i*_���fn��ŮT�! l�u��10z;_0w����BCL�` �5ϼ�kC��!8�V�gO'2ch���V�������~�����y6��Лgq�T�G���'B���ຑL ���4�S�\���F��T]T����Om�����*6�ْ�s�����?�w�-X�k������OV<Axa�zg�I^����F���� ��R9�?��n1S��"��jx�=H�7�%B��Hܧ�e�L%u2&��Z�ʺ�n�i8�>��{���E�K�έ���"�I��v�M��5<��y�W�4���pe��k�]�YW��P�
<���V��i+�6�_E(�5{W�;�T�x	�w�m�k�[6z��G���dY��&�O��k[65�!�Ձ�M�a*ua~���wE��])�k�`�g��T�2�W�eJz��Os%�x�E$ޡ���`)��ܕR�y%�`8�,֨�����uG�C]�~qa���@E�?��R{T��'��S�7�H��������+��W�r��=�}'�qI��q���G��^-�0�o����H��B&����H�-�G9���L��Z��i����e:�+���JD��Ѵ����m���J1��(���X�$e��i�Z�?����>w�������̍c��k(D����3�j�61WJ2��š�y�~~�� do�2��N�e�]S�|�0o��bqy�T�{�K�xδE+mX
�zm1D."��z���B�g�}���@#�5� "�&l��;|��"�������8&��#�K�Lt�*/oj�H��$U�\�����K1��-t�p�����Bq�C �;�k��ځ�B݄���o�z�`�=����Ygy�Xӆ;u�K@��OO3|��O�kB�Ϯ��}����dO�5J�����N��F+�XI�ĴYj:?������25N:������P-����՟v����l�N�ǳ�+2ԃ��H�GG��<�����"��j܊�����Jh$.������YɓA9p|�=��f'x| �T��iվ�i��#o��c�G�_���{	��j`�dr���}���a@{�.a�#'��o>~q�f�C�5�V��E�!�Dx8�*�H�i�#V���k���x]J��s��m�	���,�����&;d�^�Z�T��7'��n�>Pd�:&d�/����pQd�%��^��<R�� �vS�B�ʂ��Y�L��_`���i��(�\,%�Ő˷`��������V|#�%��xv�yhp�sL�7��"à5$�0j��Ky�0�oC��pn�X2f˛�~X��]����Wbakq�Cj]e�:�+�g�f��?�-��M���i']��k��^^����}#dz�����q�,�G"���0���d�H��o��t��-���ڐ�_>�\+,��Ck�Y3�V��v�<ı���.�e���I��X�w��+�;]̐ov0i�"g&u�s��J����?g?G�\�W.��߇��_P��U]l$c�ѻX�Gp3�Q]�=���j�#�j��O&E�C�1_Ug��lS�����e�V�����b�\��1�s�1�&�F�lV�f� b�~�٤G9����8\6���ukl�����)��)4C�o�����`*q?�Ν1թ�ۖvɎK=477��ݎaE��/M(J�5e���7B���.��v�����^γ��cu�gE�ҫD�v�,�U}�v�������A;��ñ�-��&8�(�J|�@����A��0��	Q���:�Ql�p�a�F1M�YP�:?W4�ԙ٢3Ԩ��6�Z�%@,��f��q7���L婚���8�v�^��g�ϥ�y��D� �Ӣ��0�� �i�����z"&�����6,2Ƣ��lRt]�ɔM�H��H0h�C�A3�Cp�?�#���r'�Wa�[s���TP^wEC���ǉ4�f�d�	��%��� 0��_������h���/�%-�߿��^����0�_cE���?.j��0�K�V<��"�]IC� aW��
,Oe�Ѽ,D���� `�WQ���Yv�fw�0!i-��2�s3 ����t+�;� <��T��Ҹ��#�䊍்w��ST2�o�����y�ЖsT�/��D4��Mp��jE��l!J�~��h0\��!��:�ӯ��M��ߐH�������2���ADjqJJW��Iڨ�e Xs��`�����g��'��g���E˾4VuJ�?49/0��8��}�/�o<�˗9ɋ<M��t��n@�J�3C�V'}r��LgC��~If�����H���u���R�#��o�db��ޮω���p�����ne�X0;�I�D�������Ѱ0Uj���%ǥԮRS�0!�j����v��� e|��}��%;�O�w�E��7 %�硠�o�H�$�p6��Z1+�7G<2س��9߲� �d���׳,{Z]�A���=��{(YbW�n %ʟE"�*T�*:���a(Ex�"�*�������+X$�K4�x�\�o��
n���|���K�O�2C��y|!�P~���y��nr.2
�1�(W��K�o�M��mY�^�:a �'�v��߫��XP�)�"��bfS1�W��-x8��I2ʡ�V|�gkx�\*Y�,]W��?g�(�o�,�p�q	����dV�ϝ'"��n��$�1������7)�E�@�ǹn2h�	����U�{$o�,�u� =�&�<��{���YE7���(LCt����(#� �Yv/j�P����oa�A�S���l��c�����m�c{	w�A�lsP�*W�'�����Rx����^_���[�3�Ӌ���曧��)O0��.D�����$���"�� *�����du�������ǟ[>#,��ao��Y��Y���
�յ�]��ub�W��},��/x97���*5͢?�� LM	���[������m��-��~��Gh�f�˥Q�9�;�}t� yE��� ��)�ms��6A������B��W� $������/�*��|�]]�Uz�M��jGb��\|��#�gru�8��.�fxo��j�G(��S��Ci[ܾg���c�5��m߉��=�K�gK��)SHw�nӿ,"�G�S�6����e��'��֜?�V�}�����X�<�X�0%�sF-ܰ˞c��ph6y9��!x6ҥ��F�@�.��Xv\N$���H��'R�)T9P3e�,�)��Xe�i���B!�R$@>��������;���nDҽ������3K�lY+��!L@�)�����oΈ�l�#WFU�	n$lM�zg��C�*9L��[0ɩ���� o���"�����4c��	|��<L�MX�/���aTI��;�j�B��4c�T�F$H���"V��)Y݂`VC�/�_�B�A�	�������Mɋ�J�tQ`����ԁi�F������$D�ѹ�Rh�'�39����v�XwI�Y�~ xx�s��|���U �qju����$ �l��z��4Ɇփcap��*�O���Nɠ^��Z��m�N�uFx�oFT�C��-��/'׉Q���JK7flGS�,��5EN��g?*����~]Yt�ς2�ԙ�'�{��$D*)k��(F��Ҭ���f|`d����_.�xJs������m7�R:�aSξ�A�cж�T\��{;Lwى�@~���S�}�_J���Ou�KJ����(#E�W�h�w{&�K�1�U��%7]N>�XRĽ�� �2`��7%� ���_���|�T�|�a1M���v�N���Wxq�KC8��?L�]��lZ'���q7����?\K��h��O�"�ų�%��S��1��L�C�]?���H�󱈹������,&�?�{K�_Bk�q��U���趙jݳD߄�=�~`Ξ�"�ɯ�g�=�@��T�6���$��:I)�K�G���D�=b,l/Ac�T���~���`�H��9���]#Lq'	�j�QR�Vm���xs#����mE��9�\ ry�)0��.C<���&�� b��.�<�1∈��Ƙ��L�myC�i��N���$i����c7n&cJw���Y~��"� ��Sl+N	?�i�x �hSn.b�.ߡ��p�;��ʑ�}��&K�.B�'�x9��"Ӆ�
3�=�t��N@���\4����3Z�zx���j�VC���r�O���ʠ��B��(v��֢��	��h��+��s��V�F����ȡ��
�%UOh���Փb����2���Z�,9�W�{�?�_�ЀP-�4�f�dg��?p_
GB��1 ,��,8�͸�<�$�siE�|�o3��fxv�&������&�X�R.A��U|y�oǪ�s�Si�Ys����/Y4��%��B�GB}Ҷ���=�ѣGԚ�?���B�s�� ��ny�$n8�K���?��K�2vl�أ>Le� 3Q1�/� �5��6�5�:�]�^I��ͱ�X�܇<iKտ#6�E��[y��JJ��^�>��J&z7+N�{�H25w��DT墌�����w��A�ؗ�����T��t%�ĴDT�juoC���s7��+S��a�&����M�W�$J�95XTc���qK�1x�
ehq�J�O�&�HJ��u���R �x/�M@�>����j��#T�a�@�/[R�8��7��&ugKl��j+FrUnƧ�]�z���B����ʗ˳S2�������Xj�?���:�f9h��O�c�zKe?��D�;;ܽ���.˞�>��/<b�0�*	@���i�j�->1�TXG�&�k �'���M1��7�=\��H�1��V��OL�C�ͶQ����]{f��z\�e:Dw='��7|�&2��F#x�[㨢c�A�	C�����'>�[r�/��������4�lF0������\�����rݩ�B�A�
��b���֯���)U��jR��"�P`��9��\
nUK�$��ئ�&���6c�zJ�7R(L��#c�#GJ���t�z'�v�0Ei�uM��a0#�2�"-"���G�T�!Ț�K��Ѧ����5��c��/3eWɱ�\h8;�������.�p�����`�~�����V2�_L��������Ѵ|m[r_΍�^a��}B��Ѿl��̠
�H��a���@8��b��2x��S-�]��Nw0j>��U����]y���8XH�(x�Z(�F�Ÿ=���%��5��ى�S���m�7H@H���o�U�gE�J]���D��_�f��n^��_��=�Iz�y8:��K鬹M�a������A`f�g�ݛ{c��H��bL���-E�sy]|�A�г�ಕ�q�Gw�R�DRuY�'�����o�����m`�qA]}��?慵�91iT��s?O�}��%4��I�q����=���۔�6��A���};Y��0ͷ�<�����Z���T�!��/'�٤I�!� ������?���;q�t}�?���)t�f%Z�#3ǔ%�IJ>'�ǲ�t�:�YF1�<�ǋ����!G��% EH6�r��D��=|.�O;[�j${�W��s���~f7�愖����2�ʞ�k�����P�Ɵ�l?6���j�-Gq�Co�71�ɵG:��x��0UJ���6_�ٌ��(BPC�F�Z�^2=�0&�@j�O��k4�|�.�����{9����� �K~;�B���a���	�\{ˌ��L���S�� ��#\�@�"@-h�`��	�n���c�"��j�v��Aͼ^v����
*q|̃f��!(-Ya��6 �R{B�Y����0�﹮b�*h×����r��PC�= /�(ݾ}=�
�R�=��IĢ-�����y�[/\�������P>_([�����x�믆������)R��Bѕ6�Í�,��~���6h
�W�'w�S7�-2N��s�{E�����n�<Td4��,k����T�I�I�=j6�ˈ�{�Cx���g��zz��0��I�eWRR^��J�	a�}�
�a�_���� ��t	�r�K�����=�zM����ĳ�x��,ϗ����Q�"�©K���x�S?	�'�_�j�i�����.�y�d��a~UK��U����,�V�L7�4C�x��[{ϯ��+O�����9D�a�-1���\{6L������n�'���:aSy��g�����J:�j�&�]�n?'�tK���*h:�R6���+���BQ�"��S�M�ױ��8 e=-�3�DZIw�Z�&6,�=�iX��5gHN�����Q/ؘ��)f���e�jl-��c�e��u�)���v��G
,,N�R4��Po���"�8NY��2iTf�F�*�(*���zVGG�z)'�xf�ߺ�V3��-:[�x����^�\�]����nz�ܫ��K�|��0�_ RS���bE+�1���p��|��w�m��T;�d!�O ss�kmk���i�bvWQ
�����������b�3�g^J*���nya���:��y�k8���'��ty{�?���������e���"q�u��`ZN��5^`���o�=��_��&9��񄑨(�T��в�b�c5_S����$��0�@ ��l��D)�[�,A��S^�Pc$JvQ3�z��a+y�H=P�pQ�ۛ��h��W�BۥRX}���a���p��Β�Y�D��ߵ�-:����R�g�'�څũ$f��I���c8	�P�*Cݪ�o�V �{��7�@�#����)00G��ڌÝ� .�j>=ݍ��E�eդ�AN�-A����yʼ4��j�	�1e�X|��Қ�<��+K��2�.1�Q�,C���`������[x2ц0�@g�4//)!<����E��ْ�? �c��)���F.~�Ҝ���\�aDm̟�a�
ƩLr�������<�qWb�|�T'E��c�E"��|�#d|�\��������)� ?q�+B'����:n�1.�˖̺���,�u����o�y�!Be�����>��봒u��xL����Ƹ�������i�����.���Y���&`��R ۳b�j��J�.�:��,A����J,�9@x�r�=�?���I�7���ؤ���4�(�7V-hf��S�xD7cg�.Ey�xcQ��5��]+�92�^<t���']7��	6iK�F� �s�}��� V��a@,~�/�[LKX�؞��6�ZY��v��,���)�:��R膞+K���ǅ;���U���o3"5�,G6��r��B�yv4��U*\L<)�<���d9:,��d{�h4����cV�h�����?	�?c�9��ŶM�:��{��s���%�-��p����R=$��+��0O)�h��H���z�� ��5q�����*1�>L9��~F˷G���8����<��\?�P^���KnA�b�p���|~z�C/����_���l�Ơ+�l=p���\\8_���������� b���� �ci̯��WL��YrL�#_e�o:�H�l��x��j@/��ȸA<��[=�M�O�o�����{/�
��c-�\Җ�?Ӧ����Q��s�_p�W��a�$ù� ӵr�<��>}x��[
�C,����^�3�հ��صݖ�[6�ʗhG�d�L�iδ"gg0� o��xxX|�q�6�*K�q�A��%�-kJj�q:�6�=8d��zaVr&� ᆈ���P���4�X[�ۗ��ܱ��t
Y#�]�|����Ł{4��<WT=��c���I0���6������C=c/��F�i�PI�}����}�߂���U �P%�����9��d� ����U�磐��zL�c�h��W��ƥ��ܮ�S�͂꬛P��ݳΖf��o����g��!E�]==lذ*6��f.X�"��4+q�.0y���cS��BRƱ��~�����0=���YILz�:ϬB:KMg���_�e$d��􆜈��7F?��/�~���r�S �b�3�%1D�����x�.��yT�@�(7BD>
�u%�gj�h�Q Ip
-�kU��߻^4�z���@�2pټL�J�����,���DB�}�Z&؈�k����m���;<3G��&��Š�%�\&#�Q@_]�D��s���{{�<�mjw�y`���R�#��}�V*��p�Un�>T��?.>�cpx�{��TJZ������X#��"�pU_�W�%�h�`����H�lS�Rֽд������s�-%W�Y��x55Î�J�0��R<�ԃ�[d-5�{�1� UZaI\L�3���	��7Ү)��s��'$�Q����Z)&�^�e��j�ke32&�}��Q����o��Q5�@u"��&N�_)��=d��h`�;'�:��+Ie�,
L>��r����j����YB}���Nh!���[���f����|� ��0�q)����b��mb#@�����w]�^��<��s��狵�����_��o��#@�I��3p��GF*�:��KsLa!j�J����V�������;�q�Hf�h�x7\�X!u�?x<�̡���P�m�ų�ɐ�9���ED~��P�~6!���E�ʵ�gk��3u�P�B�Ƨ��47jVD�0�6b��WY�Թa<��e5����D�͈P��r3���_)Y����F��*ԩ�<��ࡘ���Ґ�O��hv�ӫ���G�A��fC�+�=>�|��o�|XܬG�C���6��V2vo�:�y$%�i�%z�~vP��6KH�(޷hѯ�\�̫�
3ެ���e�y���/"C�;8<�9@�!g�|�+�`��ݴ ��I�D�Hw��U��T����~��O�9s�Շ�'AP�h~Ɏo�!��@H��O�ڧ�s�H��(iP/0Ώ��e�bͥtaw8���r�+�]�߹
�yr�,I��E�n0�K!�՞��0/�#�ma�d-�a����Zp�k���BT�U����G�(}��n�Y,'��ll���Zտs�2�O�ƒ�wQ��d��E)�!\ĭ���]���������9���?�W6IL
u�T�d��A��������3�9Y.Z��t�_��y�U�u�ƩQ�冓7�cv�����vNmN&t� ���M�<�zk��ԡ��#�����C�3���1/�(�	6�)�/�y*�d��ߤ�K��?}ط >� _�4�i��� �J��炼�MZc�Z�z��?��l�T�w���_��&o~9���U�͐�R��@O�󿼍P��u���Ƨ�&���	�a"ڃ[�2��GS�Ȟ)�f:|%��2���5�zIO\���uW��uň����Oi�U���?�v̞&N����Rd5����S<���`66���uB9I4�:�!�73��,D��֚�����6ͩx�$�.h��ԟf ���	9�ڇ5N��G:t��O�~#A!E�����N�'���Zc�0�lܴ��*��G�����˾�w -�#�V�1�o�~^a�7+4�0Z��(F�AE���]�Wa��ƝSW�{����Ee�Pf�N
�����/�M��O9�c=����[��r�®F��<��D/S��5	S
��]�'�܋;�z�B�X,�����X�4T'N$�6|�Զp�6?<�%������r��g��)�����V>�_0 $�s!*��l�NhC�u*bc�"C�f�h�(Fo��g�T�q0_�^�ū�sL��
)�֖��x��}�b��s)j3=�w����""����=���&6����C�
hZ���N�1}�(�M`c@�=eT���idq��	�J�EaI�E��`Wq����p�p	��N�x
o�6�������`�}�/�y�f��i'VH�����>����}[i1�O�'��V5p������A�W}�ge���9=D�x����o����CP�&H�y��Mˣي��f����B����|V��F`&b�3�M{�&�^Qyd���;̀U��;�*��wYMt�>���.�RB������F�QriAS��W�{&�4f�,&�2'Mۮ�y��lY&�DӲOb�Xj���(3Þa�C�+|]��q��ޅ�����烾n-a��B��/�l-s��}��H�Dv-±����x컿��7��Q;7P�#C/�!��A"�Y�7��ZmhW�x�J�E�v}9kT����AaZM�t��!��X��9��!͵A��O�����p�F2va�e�57[Y_f*`�up�ZC��~e��2��D;���	�8�V��+*����Q���|��,�y�K�*C��o O&�c�Kf�D���꾘%h�A��ʑ�좝�Q�z|uk	V��{�����=H�SIT:GU`�m��
����~L�8X" 8�F̨>��]������C�I@�U`�H�o��>��!>������!��� ׸�"�*f��̿������d��2ˏU�4>�CHYe>Wq]Lg�*�k�D�,���T|�ԸqY���cO%g jeˑ�I�[�z�,+���gd:@[�^&h�O=��,`�꾁��V%U�6<]ns(�kݸ�����s������Fyko,{R��:#ɪ;�E�����ҹ`y�li_��$���V�I�#�Uϕ0�)�'_�?� W���/u�2LB�k�ʮ�Tŧ|rPS>q�'�Yς>���im�<胱߳�t����O6���g_@�=/���j����k��
����Y�%g.�69�����s�.���,=�n�y�n�(*EI�U�'������s�C����n��Yq��B��w4B~��w(!�az�t����%�G 7���A��t��g�<���=���6����f���NB�0+r���x3E��5��b���*�JH�*� $�s7{���'�0���f����ۊ.�ӂ��&b3��?����.O����r	:�-c���=��Бr�������0@�$�y`/f�eq�X��g��A�x8�}a�q� |5�6 ����< �%���A���8��]��� &k�qcmǜd����w"N��gQ��8�:������%+�������`��=�����t�����]L,MdGxs}� �+P��~hs��i�GҺ��;h�P??������T�4��@����۪�
_&�Q���i��b�6~��RT���'`��&���`����`�5%Iu���R�i��a�whk�>M1<q����&˒$����>Q�=0t���d?�Փ�'~U��P����4��!K��~W�oy��g��M8a�$.g����{V�>�uk�H3�=���5��xVRΕ��vx�/?<zl�� }li�BX��U(��]BZ��.���@��m����(��*��؜����-�SXދ�<$+%p��g-��
��X\UT�Ov�{�|F����!��=�:{�jEt��B)Oz�f�h��|��na��-"��P1�&?ǘ�G4B.�eCTP�Y�p�FfЛ���Tn�<v.�	ݩ̂`���n8��M���L{�%��U�r���tv��tO�C�8��K����]>Fy��\V�b�@])��)*9o�p0|�I���aRI�&�����e�&�����Qv�+E�� z�[p��f�N�*�U�J�/����x����E �+��G,��j7�F�]$��Q��4mlM������W��;�}��@"C�k�1:_�`t1��@��:�����*V��V�II	A�-��%w�>��:6�)/5K��k��K݁�
_\m��]k/�o�.�C�\�b=�[,Gќ���tS�"\�G΃�k�ؒ�;�[��5x�#�Ϸi�x�5�!$X`/0Ɔ�Ġ?�032�{�@�К^Я7.!QC/���ê��aK�������w�n=��"׶�0Á�#���~V���ӕϵ��o3����|�F�vz�+g���( ���m�+�ɏ��Q�	���-�S"�}���*��^҃�P�2I�C�
��56������%4Ȣ�!۹q,^��0�J7�W�j�G��D�0&�~�CW�)���B�haP�M����ݙ�����u���.�����hʛ�����]��	U�x�Y
��j��L�+�Mcl#iEgw�
S����A�n��|�1�T��Y�Z]oS����� �`p豍IS���JN'-c �eP�E�)�[���Hf��%�B|�Hmϒ�l��K�l/!;�vB+#�E^S��q3��?
mJ�uԋ ׃bN��  3t��<���-�p�MGL�<��Lȍ(Sz�A����ɪ�S�Б-ޫG��~wdy?T�=�����R��t��N�}Yo���<J��ˉ+��z��7�D�8}@�y1l�M0��Mm� &'������J]0<Ĥ)ׯ;�Ȓ��:�)�0#ae��F��N�l��8��	�k�$-��w��5#ۖ糏�x��W��!�l�~,���x��ä,�u��1�D�����u>���h��2�
�돀oj��HBl����O�.v�	Ƒ���i� �?/��Z�&�Q���դ�e�L��!#�����@���J*7�2��~lP	&	�Ud��5Ҩi�ݵ��||����DK�֎�R�DT�6��.b4�	���c��lOU���Z�q�_��F�E����/�4�J�NC[�d�k�3�a�/W0{�F�'��(��2^�k����7���B����9���o��5��$�b�-l��h��WQ�;�=Rs,8�LI�-
�P�?��ll��Жф�*-�-��a��.�¡�P*ҹE�j��3 7f�lȮ��tɔ������O���Ɠ�1�(-�ŧ����dLf֙�~���7C#_a��yPS��e�н�'EX�:�(�%�b: m�t�ƕ��b��,)a���2���#��W��^�,��z>R�%��-�����C*�;�ZpUl�ߪ���ؽ����ER?$7�A��(a�8J�(�0�6�\���=_�'A̱�кi���G	gp8�,9���х�Ii23��� 6ՓwWz�xac(���;����N�o1k.=X����v������ǵ��ཏ����n�ž;}��
j��q[�ђzt)q]�
1s���%B��P5
�<�T�$LO裘?� �ޱ`�}S��Ek��(��W\��i�s��>�n��K�׎�9ǑM�dX�+����K��-�N����h�{�� �D/�R�c��p(�5�}��tgd9i�dB�f2��n�/�4tZ^�-Շ���u��w�7h>�����x{�W�K^EmJ0�A�e`��]��E­��������й20��7�8�oJF9�U���1��r�G��vk� ��a"��|��ѵ�o��;�*&㳡Ny�g��3�	x�Ed_Vd0b����<d��,]@F#��hŻ�6gTh&=�:��S8q�g[8���?���Y@��m�m��s(����v{�7���1��Ō�"�y��	'���o��m����������	I�	z������T:e�ޟs�%3X����u�v��
ŗ��i��k�)^Y@��
��`��+�/x�MɣZgd�#�L����,�-M��Ee=G-�i#�C��@��u��#W��|G�V���L��5���a�	M�}�ad�8�w�a�Leǅ�[L!�8F����&��k�j����^r&�F�Y�܍�X�rf�(*;�p�79#6�[3rL���̬��"k�U�{�����F�)y#���4}W�,�ƴ9��<5n�{p����3�$.���-`����5��X���W���>-�K����\%g��uVHh.����	�k[9�0wq�b���@�'�o�.����㝤 �y�}m������s�c�/WaZ�R9�n����K�zB�2�-;}���ַŬ��b68}����Q'Ā��0�̭��L�ު����`��K)'	��z�������x3븤SY���Ԫ-;��0� �
~|Yȉ�y�9������L�u�t��v�{�߅Z�Z4��Mv6���o:m�R���C��:O�f?����0���+���ſ��1�3�����P|��6B��4H=���N-��޹��(������LZ�mI�S��m���ܒ���hL.ܕ�.k&�d�K�ͿΜU�^��_#.��A��Wt}�v�r���'��?%�o���Y�[o�m��/M��f���J�cg^�^%j,�f�R&�8�Q.o��y�q�Ѕɘ���r�HyI�Vٲ�0f���k*��x_Z<9G8�P�����GyV<(�����*�o�`Oo �'8 F���j<;���y��K|��sg�IJLԢU�D�Bf�P���D]#��X���i�x0�7i��un�i=އh�W�[�kA�:1Z���*J���+�|�E��T!�V���>n��O�	��豑6S.NG�����]�����Q7VyF�D��uC^���������2�H�h5�D,Cv��[g�/`GO���VW��\i�����(Z��?OGy�u$�W�4D��\GKl�X�'+I��T�����}i�Q8���7�<m	w��G�n��H��Ä�ǈ��H�k��x��t��囃�W9�s���Iƕ�8>k��BW���&_���Y/|x;��q�!�C8J�ؖ�e.�[f��zB��)[1Q�,K�d��9�r4r=�66`��;��;�~��eG8�F'��A�G
��Ԧ��g��ʹ����V�*�wì�`�Q�?���YDv�g0�b���v� ��2�D\�)I>�at�V΂�D�M]��7��,�Lբ������l�?{�ܼ`q%8��$�c�t��-R��Ҧs��	���f]O:���@�a���8o���D4)��\�p�>��:n���?� p�#}C�B	����7>�SA�c��Z�* R�G���7���֓� ����e�vVlw�6��oM1Yf�s�0D%$P��'.i� �b�	�mj�<��%n�߽+bֈx�+}�;�L��y�z�oG��'�(Q��	�>#0��<6�<����������i�0�3����R�k"M��KP5' csC��o`��W�FD`��oU��ߨ�>�����5ob��#+b��M&���$f�V�I��f�8z�	T̞��;Z�6�����6{��	Yc����F�a\niX��v��f|���k�KUD��R8_:���<I��c�*�C���K18Z��&�SM���%;njz;gC����O�TF'���)�� j���*�,:�c�JS�4�E���ݳаB�+l�BD�����b�>�28V�����?�K)h!�!pJ=�F����ެ�e��^X�t�D�6��p�Ҝ���bQ*Ǝ
͕(�z��j�3H�{��N�M�U ў�ܵv&k"��U�6L�r ;���S,���mc�p�2�����j��ҟ��4�"�gHcg.�\|U�;���������CLw(��þ��痦=.�@\pU��[r� �j��@�5�_��c �6B���"0@,�"�9Rǈw"�8�]��� ;�,jLƊ� �Q��l�h.;A�~�Dj��h�i|������jn��VZ	�SKJO"F�]��NH�_Z��C��(t�G#����3N	i,ٙB̼��tƋM(�W?���܁ �*�CwU6� ��`�n��t�	4�����<3y��꽡����O,ة�N��Z@�
����(ٜ
6���i;8�;.���sG�;��{�{[�X��FD�qv����g0�������\z�e���fo��+}�Dm��5X��H�^����10Ϡe��7&��a.�1.���ʉC�=:_�lH�2���؅ZQ��v'zc�G�p#��������N"�S9�I�{�>�`ؤ Գ�R�����/�`�9T���o�c��~��#?zQ�FI�#,9�W:��Y -tcBoȫ-!rm��٤ӌރ~�g$�G� Q/���Uq�7��G�D�|Dz��\��s�} �L�>o��Cb.�3עY2�amI$�>���q�Ӟ1:cy���>K�V�F�5C�M;�@	NȘ�;���|��+��\9��ꎦŏK�$�貳6�K�����(��/wr�Ϥ7����g<�������w�Jx��I�T��>���[l�L绸��-��\	٩h��vӕ���-��$���^	�F�轝[w/��o���M�lm��a���0�\$�0�d`�T��
��GX�<�>փ��v��z%]���	+����L7� KA�o�4E;j��_A��|\w;�K*����T]�ŉ9�;9��(��v�m��湏��h�4������UȼT�x6��8�1�$�|v�87�!od�$|Q"7M�WTsS���݊�QVb-�R	`����{��K�m��#�����w����T}$؄,����v�=��2L���F�|��.���쁗c�����S>_�}����;���f$�)��jt�+���=�Ó�Ύ^=e�q	�(�%�M�$Z���t'i�B `.�µ�Ez¨��ѝT#R�{�`"�� ^'���s���j���{p�����ڇi @�6��w���nf஛�T����	?mu;�A[��#F�Tj��@��I���ӝ��;d��M����:rr�o��BI��<�����B�<!��	%�ej��m����X��������
L�4��_��2s��Pެ%��1�2��B�bqE�ocfL�*��?�@�����f�kAa��d�5s�򨑍A!6w`V`aF�5�	
-I��G8_T�4�EL���D _�z�@������"�T�'��>D�E�4�n�N���+��  �����R_���ǂI{A�t�7<�R����2�3s[�ET�%+oBS=Zza4���+�<,�*1�4��|������v�%mʤqr�~"��?�˩}O����eNm��z!a�X�-��9۶P~"�ǜ�z��o	���9�1���0s����#_�<N�����n
b��T�.p`�Ih��9�!&a��U�n4�����W�p�k3j�>Gz*���� sS���ŹԴx\N!��&��`�V�On�?f�8L��f��zs9�^�|9-f�H�C͏�x��e,p�Z��}���&����S,}�e����B8@�l�.��Ѕ'|q�	T���<I F5�`�*J�a��T 1KH��%��u���I��'N��]�m��D���K�������)�)�#�š�҅�.¾G����܄}n5���? @`ł�⹩��ъ@��Cőh�;Vi/l���'>��{y����{&��(�ʣ*�ǼȋC� �&y؇n+�rG����J��i�"�,���7aTL4Y�`@��m�w����:Ѫ��5��s��K��P�߰��V�Y�
��y��!�IH,��U��)�~ �`�3 )�&��{�VvU�C��2��4�'�z��s��0��%JY�hv:z]ƚT�GN�q)��X�\[�ϻ f �	Nhh;�9r�8-��3���+��!z���@�pt�����	�g�qR���+ ��Q?�TX�*�6�P½�LM���i�'S���)=����l&� ����O���n���X|]��Av�q�����	��	*�N;�%�-nbR��G�U5|�z�1br��j���L��"
�;�N�7��	���5�*�	��*v�9�M!��z��7g���3��,k��F�\��x�#�����+������V�na䵾��ȼJn®ަ��x����d�U̞��OQ,��� ��m-�+Аda|��d�4�݀N�~!uZ�j�ű����t�4���E
��a����׾�@�O�C8룜����,|�����ʢ����d�~�'u�� ��5���$2��]�uF/&R�M�Q@`b�\�8���q:e3�����#�:M[��tޓ8�4�J�='�x���Da����B�XGH��tTF�bf|c9Q-m?�W�9o&x�������l�PW��s��_�U	��~��D����"�F874vD�L�n�}t�-��İX�b��+��}�6�Fst�������pϞ�� "�W�5oXڴd;}}�
(3�X�~��Wo��:C��Ä��|�0-�f��o�N--6 ��2B�_�5���B�+>�sQ���%\�-����y�j$�G$mf��F��[k�:�n�MB��a�kl/���I��V?��b݈��rI��`�=����k��=����7�t�߻իX$2B��!�Ӊ�c`�1�̳���6�sPB�)X&����6f�P�a<=.�B�h,�	h��3�beK�E��.�����Ѓ���b'��~B �yGc��*J� ��CPy2,rF�@0��e�5���D�܍֡s��m�;-n��!�%��L�3�,�'&���N��P��jO�D�*s^�,���;(/�iHzq5��J��"�͑v7��-U�����.��K��p��=؝�������~o�bh�I} h(��v'a��K�b��&)�ũ9]\��r��쪮��/��Խ�&Op_�5B�i2�.����Jf��'����E���1����_W{P}>�U�YY5�5`f�=��jH�d�Ŷ��r%���%���pϣ}p�]%�b1�n���Qʼ�)u��h�o�I^�]g,ɘ�^�������������̧�1wF%̗h	�A!��`�';�r��1��L��¹$(?d����[c�=լ�\�@8�텐��9�J}]��̡���71�+H�^�x����(v5�6Mô�U���ܵ��'&��(k�B�*C�ħ:{�MS�̈́��4L�%���2���L��V�h\E#�ɻ'�L�cGs΄��HV�ЕqZ�ΝBҍ�*K%�(o��&�h^di�PD��	��|�=:�լ>�J�y/����YjV�<�����qAe�Ydց��� ;8Hu��k�\;(���!V:Vv�5A��������!dh�.սP�UQ:R.�PF�
t_h��O���`I��)�?�4+���jU��J��m�N%�h^N��� ��k:|��ޭV<�ɘL҉Ar��v��!R������o~f� �?a#��m�J�셪A]I2�dEAV6�5J�{��t�ݻ�Z�Y���nX�`�`ݵ1�y/��$�V�֮V.������{�V�'i־řj�I� L�r(����B	І[�:�ԗ�<>U0�	�jZ);�ݜ�0ԌP�ʳ.��S����2t#�SI$�MG���;�/a�SE��y��҇�,�6y���[u����A=���T���vZY��a��sĠ_��K�߁��/[X?��� ue̊��ޢ@��-�6�M��km͓��.m᡽��LMۇ�8fѩ;�[}i{A�����<���"(b+#Ѕi۰�4)�҃t5���#��v?�����iGf���O ��v��c��s���B�&/5�¥�IL��)��v�#J��k��,�/�$Z=}u5f����q�`�&4+�˦���`�A�}n,�X��2F��[�Q���>]�P�=a��=��n��QA�M�c��z�̳�AU`�?Q�<#�Dv��l��V�2��L�.$���8C7��r̕�0u�p�x����x���"���+/�Ζ9��ܒ鰥�3A�%��g=�l6	�6I$/~�t��ʺH��L2�8ۮ}p��b���)���y�iRG~h�Z��$��#̩,��C��~/B��O��FIk��%rJv�.�x�n�ҥ��W��b�m�W�>��Ea�߁�!���Z�%{��� P=ڼ0�zp���U� �9̟V�&��
P��;z^�~�6Y��$���e]"\/�k���D�@|4�wa�fm㱑iϨ�	�8~ꯥ�#�B�V�l����)��D�"�=�v�#h}��S{��{��EW���k�1�7�F��a�_,�XB*@^DP�E7�q�η:yH|
�Y᠕_&��˜��?�m̝&~e�$������$���b�U�����hTy�	������H���'%쓬�(�#�h�Q\�5��Q*m%�4�G����M����8<�9�YX(M���e%�{�YGT���7|jT��B�$���p��=%�3`�bqĢ�X��9ۭ�@4qoG���ZV�ǋK$Q���Vm�Ű�τR���D����#ԫo�O����#��y6GY1sGp�y�~���Q���F���D
�W	<�����,�n�I�7Gaq8-b��M��G�&�XF	���9$�	�.Oz��6Q�1�<�b���b	$���~a���4y<�
1h�M?� ]9�]�Z<���yo+�� -�ɲL�G
6�e�y4a�jhv3M�@R��R��둅7����%��50)aؐ�'��r���U"�_��#Y��=@f�����N
�h��
��U_�+(1vm��\Q�Q�p�E8y�A>�3ضq��[��+�d�6�k��{��3p�c�����ؽk����n������4�N2SCDZӇ��~� ����]��N