��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ� g�I��Jw=���c#hN�j(r�y��l��Φ�fT�	Z1�%u�dXw(؏į�� ���q������+dF컡jea�Rw�4Mh��K<�%�]J����U�b�C����8�YB;�R�Dv��Q�0����}e��^�K���q���lyd�>�o�L�l����b�f�h+�rLV�:�:�'|�4R��J�HJ�~������]�4:�/p8{ӱ%D@<r����47ܚf���?[���P���:�&��<&j�����:�tQY�:�A�����b8T�Ԟ��n�;�~:'�H;��.J��"�j�v%�+ub���pe;1gW��V�*���l{U�`�.E��N�M�X�kd�<*ϐd�);��ϭt�h��d�Dq�ao2/{ g��n���S��Üd���Q=�5t 1~Eʓ�ÀB`)��Q���t�u�зb�chaչ����3C�~�;�-��Dn���������6��	���C,xo������B�L�y��5�<�ܸl#��OM��Ze����(m膎� �*	v)O �B�e��� 	�餞D�D�颰	�%�4+��T+Nfa��T�X(s���7��Ǽ4��� 5q��s��d���*}!l�l!�MЋ�ٸ��
GE~�p��S���Ύ�lw��QR�wTu����E�z�>B�f��f��q���]7\P���t��!���������h�p�UE�q�0�˧9o���I��>A�A��)A�Έ��Ei@�d��1�-�Mw���O�<%����$���Xc/�ww�%��f��!bt\��2���E�.�b����7��<Y =�i��~�(d{�)�����6��/�i����W$�����4��=x�ƴ��# �#ڰ�q-,�4��d_�-���;��$��?�gܫ�����!��T}y��$s����{XW����b�d8v�@�<y}d��Ftj��bN"Пc����=�2U����!k���\�߬���L�8Лx�^�x���)sW����~l�x��F�hʃ(;�1�f2Hd�F�C��/���n�����\>��W�`���u$8�e�a'/���[4J�0]�/h޻7'G_w�)Zit���4��7#?�B��#�:Q-�A+� 3qx��GZ��MP]��Iϟ-��	�-�9�T�(�E�'�{)�lQ���S��#�bPr_�=���Y�8hA��� �R���
{I�⭄��?�N
c��Z������(*�d�$��j�a��yS��e3*l%ݒ-m�:d=X�i�k��`�am���.ɒ'�t�����v�%�@�B�?�o�e�ӱ�L�Ws�}����C��}�BJgz��.!O���9�I@�ǀ04��L�>	d����(�$�'7~wb�`��u�c+^9N���������q_��&����Us����7!�0p
v9m&�3���q��pm:&��]���`��'ú[SJ���E�"��<h�ާ`�yw'��������j���CX`Jw�J�l`�<)]K���UH?%��������#�@;�jz���#��Rns�p.�k����&�)���	���7�Vi�J+q;O�^�����GJ�`Y3���͆�*�Z��t�{�l����Gk3B�`P1b��|$Qe5-Z������Ҽ�۵�g�WXH+��R`Ktj�:{�h������Y�wl�I��ŬQq�j{�Ⓟ���i�8�]�-왥���.ӌ���.�F|L '���ܚ�H
i�d�	��T`�b�F�m��[He���~�^1�8���4���~D��EȤڵ�](�Fo�Ƽ�{⌂U��9��>�q��j��8C�����%�P׼�	9��yơ��[{ Ɠ@#���0M����v�"��%��3ʅ�eu���ha�p��3͊��W��<y	>�$/fS�4HqU.�C�����@K�Ч�!��L��4<Ҫ\�w�k�]�X��FT�=�QH� �4"�����Vd�7-�؄�m@t����^������c,��h�6�*J�=c��)ﯥVb�'=��z
����p�H��J
�����q�^�i��J��1*�ۤ�p���킮_��|*��t
�β�[5��&B�$"������d5l0���fD�����yM��E�����ӻ��Z
 Sfہ��Hn���Dq�"�Loǆ�'gO˭�%�K7��kV�`�H�1�HE{pvw����5p��˱���e�k�&CpQ0s(�dPD����'��id�)���/}-^���*�1ù¢C=�J�fq��}������X�Ͷ��F�=�~E�u��e].�,!{�����a��s��+$���;�t�]71�%Ͻ�X<S�����!'v�r�a�sa���fǰ���%U��Q�հ�5�r���S���%,C����r�p/qf�D�)�����a�7�I1ٙοTn`'����s�}'5�v|l����(�,)�Ӱ�]
W_ji��%�ҟ8������z��rqh3��HL8!vm53��O�dh3;�B3�q���$�>���ChxI*�����~�2��Ț/(�z��Yd)?���.��W\bD�Taގ)Ys}��ښ�!]j�yw�ܐ�7��)��p�QOf�ڍ�S~�#亣��^�M�:h�X�A&DH{+D��*E n�-"d���BF?��}�0�e�(
��x��e}+Dsj�Jpg	.�\x=_. g6�R�I7(��ǣ��@W[^�����o
����\d��)gɦ�b`F���C�*)Q�t�	�>ò
$��ռz��y�!m��k�ă�1����l��w�lު�H��s����53�2uZ`QG��_Z��D�r�t�3��]�Y�~�*7(d�R�>+̻ά�C�8<��e������<�IU9��,2
�'1F��o9��w��a�����a�8}B����Wp�[V"5��rZoӢ�,���Q_�*����a^E.��#���ѫ�
��3���FP�z�K	q����'.f�D�����
8ʻWq_� (��4�s^�<,KqɋS2�D}�?%�cDq�XG�2s��ZM�"s�ӎzA���"a	�Dv���I�f�׾�ȀZ5N������KI{�pS��
w�K˶�v�/< lXFI����0RC�������D�1�sVb_-�Ȋ&�M^p�^�ω�
v(����<�	�U�<�4ЌeNH�p�6M��OsEЗ�nBb���{Zq�~��[�b~"�b+E?���ìNX�{� �Rx��DL���~�Z�0�������XH��T�!4���~���u/D�"�#��@�Ӗẖ�c'�N�a�ǭX�7� խ�[h������t����m��Ȅdb{=�Z^�|�*���(U�|xdU[�cR��H\q�\G2�t���h��Ǯ0q��Hc��BD=��T|X]�I���WE&k�4<�þz���j��;�e����0_,6qtO��'�܈�L��9{��7E���鏛i$ �y��\���RG\ؔ���(�.G��%�ub(�k�1p�S	� �3����[6Mi�48mH*4@�zCd�(����`!?)@���	L/����_��(h����qRpT��p1X���-6�lk�|����Ȝ/�D#')�&%h�e�j�� b3�D�'�9��&u���l�k����I,D������
4���>��Fj�ʨz�γ��y���,;�k���1��^T�)C���btЮo[���}�����(T��7?��c�R�%N*Ǔ��?t�_fxN�p_,�ϻLͿ_@���ݥph2ȧ|u�f���R�����$���x ����6�cE`O&LkzX�P ��KLi&F�<p5��n�� 8B���<���;q&��Я��8��Z!׃�j��>� ���4h!W�������al�6 �u?Ь9e���=H"�*"�sGV��d� 4W3�?�82�
�ƞ��@��GTԊ�e8�W�N���xɑ���_�<-=Л�t6���GY����O�3آ�sb"|3+(���%�sU�&��2�qr�R	��N"��Q�����B�J�n6��4�@ <�
�C,p��xi"�R(]2��.�6�ZL�)f�,.:�
U�0K����V�X�\3�t�AG�&�(>6���.�&�����!\��i�:��#D$J�~��	=R�*~�,6O3�9�a��R�
1ln���N��YY`#�HqMw���3�F�5%}A��,��)񯃤e���9 �W��W�-t�G#J�s'�6���R�C
k�0��r��$"�+X��T���Q�Ԩ�]�V֎��ӑ��]��Q�V���=�g�2�fݓ���H�9��z��w!���a`���
�"������)��po����D��.�����4n8���D9��ua��m�c�}Kf�>a*�����J���%�36kQ�|{mݳ�R`� ��G�I��y2	��ͽ^�u�
�1_�yQ!T��ҫg�n�#�%Й�AÁ=�'](k�Շ�ߪa�MBG	0;����'��i6k�m�[����f�Psf���lJ	<t�-i8�|U9.7⠝(��"A i��$�w�m�y^�C���dA��$=�h"�J<���Ve�4��Sa
D]iD����Y2���˖�'G��	p�Z��Y��4[U�a���ooF��s�Vڍ?(�A?O�8	���0�"
���cK�2e܇���5�wk�`��`�J����=W5���)԰H�ݔW�Z�[^�f��{�Ț@ݺ�������'��S�)ѫM�����i��������o�T�\&�n����O<�Dd�,�u,��&r3P��܅y,��k#!d�{��R��?��_����G&̭�S��{l�fYEh���ξ߱�����	�@B;OJ�� ��x�Y�4���c���F]y�Hb8�s��1����}`��=�4��s���2C��"���mb�y���q�me�x���@n�j��h��lZ(����*��Փ���؎�~F���8z�����
y�vP� �K��������*����ۅ%����C���~3�R�Z���sdL	��M*�J����G���;W��Ww���<-�� �א@(!�!>ʖQ�^�q1i
��I�����2T�|��U��=�L���oVK(�_��4�������K[B����P�V���4H?�s��O`@�DZE��EA�21�Ґ�-&Mz	�r���^���M����Ū?�U��"��/����������T:��j���y����徫d���:y��4n�\.�#O}�:�������q�طPH�U�3���C�5:�`����ݦ�n攊������^G���U��V|V�Nyز��SMw�71��g��J��	(�H�+,Z=]ŬSԺ����� ��y���碁� �f��"	�}�7Z(�~N�[�"��ؒ��z!2˪�>B=��t�h��N�VG��nZ�ji��(�*�0��n6�W�7���=�3 <a���L�0@yG0^���sn�E]�i�'BG��R�#T�j�*�:�u@ł�>.�D���o�Cϥ�/Va;0�|?]%�r�pZ$9*�й���h5r/��0S;�x�5RA3��z��'5�͎�� ��S��oR�^���i�x�b|N߹c�_ĺ`"bg�]�0��|��4{L�"�vDMh;�?^5��W���*�:���eQ�z��t%!s��Q��2[ѥ�G:��~%�`�F�W@P��M3*7	߱�$�	lnn��W�3�֜���4�:�y=A#<�<�:44i���~0
Þ�1�,�E�pc���f�M:�Mi�w�E�8�9��k��曖4�ʔ��L��_�lD��pLO�KA���u þd��wN�	�Y4��&��Q��F;c��m�PdJ����0q�<R� 
>yA��8�N�
ML�>Sz7%�����Щu['�e��#o7��g�FwX�Ph	�g7U?���7.���/v���g�yQQ�8���.�KߑDz���6i���<z��I"����?�8U�fNY���"k�s1m80���c)������T��,t���������RL����A���"w�
�S�
~�/	-� q,Qw9w���_�x�r���F�7ܯkǖV�g��8jK�1F"k�b7�Qw���(�@Cw����(��C�^���Q��T�7�wk�t�!����Q:�_Ow+[�L�}juw��Z��#�|lTjd�m�.z��V�����o5K2�(��I$����UQ�v��}�6����Í�4�7�6�k�P�xK�:�CY�y��\g^��x�� ֮+ �+-�9nq>��-��*Lkt�7niaMC)��t004h��0U<>�R:-�d���f։E���S���B���)�97��2�P'D9!�H�E²�h�*i��p���<���֓):JI)����6��1��]\egT���Q����tk�f�ßR���)�wb"Sp��	D�?�XU�nz�8QV3��0��B��������v�
��R$���6�嫴[h��d!���iqx� 2�/}4�TU
���ʵ�c�7�ꑆ6d�*a������DLq�g+'�9a]D&�] �,�)o����m4ޣ�gqRfȩK͊	��V:��lD��<�i��e�p��x�T��b9���Y�	q�2�fw�Z�i�/H���J
���
�\���ri��i`��IN�(��-m���4[��Y��
�bX���R��Is���?n�Ä�s
��V����M�~*CY&t@1P����‣�YȒ���6����!�2���{�[p�_<��	�_�9�����J�͢��n�4�`Ɲ������?3�$�~�����=WDbuE��;�]����������d�T;ԭa�*�uɆ9��4� ��͙-�W�0#��.�\����.�PTx׼����h�E'���U���'��e��\�P��Jϳ�����RRU��Cd�PG�C�k|�J�a;&�h$����0��R�Nُ�bS�Ü6b�]�����J���?�

�ҍ�1U���p�T$��.��I,~[鎗]1t�-޴�\�-�q�;ԉ�f͓uo����݇td�8Qה�j٦��=�h���ٕN������I�|D��zM���B<�_�� ��?F+3"�ep��ţAR;�]^��e
 ���I�,)�ͅ1F���c��'x­�B��qK���\���bB�G�/J����'Dz|��mk� �[��
s���Gv�W�r%�w��}b]����\��X�l��}S��x�X�]��x�E���<0h��W{�ȡj���(C��E��[GE�L���C`@�����t�9����`-0Ô�&X���#3��_���/F�ؐ���da! R��i��qN�P�_��E?�6���Ę��7hJ�d&�O�ʪEU�Z&,���>�#G�Đ&���; ����mu���Z���`��ļ������誝E�;?P��x	Ú��� 
�(�p`�K�g3d$�iƗ�M[�����c(@��d3B2~�972�B�̌Z�
3�w�Ptnx�2vH~t���Ζ|�E!'�a�2��
B����Z�[<
F'�N�0z�U�l�1��R���Y�'b&ugB�
���^�sM� x�HJi�%�*�2�0%0�ƈU���$��3~��l2�
e3A�X3G��9���M`�z΀H\�<��S�ND�e�����߭e�D�}󪤷�3��Fd�4$7��E5/��h��v��)��ʋ#F/w��e��C����EU�rA'�)HR�z|�<�ѩ�p�͚ .�D��M�!~|3�ST�8�"<�^��m��M�^��>,`n���Iq濩M���w}�nW:�,,��
�?o{	Uq�o�O��|�<2Ķ�f�]
�j����m�}`�x�qH��Cݎ��GM����@�ڴ~D���yS[l���-�����_;�rN�e:=uݣ��:A���&�>a���yd��р�_�o��j��Ev���=]M�F41�%5^��ZUi(=�)�u��!�]��RG��y�vlXLf��A�AR������4�0u���닗xvP�U�KF��C5.���"}̜��Q<Bp�ʖ���Y�P<��� ������,j��{s0���ƹuʝm�Ư.�$f;FǁK�64:S��QA�zt�I<x�?;�K���~�Q��2�	1������b�5�/~
��=/Ҟ����Z�nG��$�dc9�;o�wnr�t�{�;��v٪,�&��Ǒ����m]#���6q�FE����_�-�D�¶t��[�Ʃ/�����mhV�peq@��߽T���[U�������<\����}XU}�p]s�0=o;�S���E�n�W0N�.cܗ<+L{�����	���3?i
0�&�H
8aS����!��;���T���:��jrk�AU����L�Eǣ|��S�t��s힂��ĩ� ����	���?5��!�.�&�G��֤�k,�0��w����ѷ�5&�є�v�S�H�k���`�3���%��.�ch�j�[=�5����0����Wނ��H���.2W����#;�v��B]wE�����,S�i܃�ʍ��2�QE�@޹a�I�C��w��;�7�s�}��J,�����$����ZG.��TI�tݔ};s�#ګ�+��e��m�d���U�@- gJ�����:�y��O3ȫ�v�fƶ!$qvKCx���䖟=n�8�ܒR�̯gG輠���-
��H��L��D�B�.U� ݳ�ȭ�.U�W�3�Z`�m�m�*�u�zٛ�Џ$���u����� $S�8 ���&3��H�Ɇ����5��~�)���4����Pے��)�?/F|蝚/������zr��
/��	�5�Ƥ�k�ԭ���8�IY�5�r��n�PC,������g)��K�؜h��!�����wW��Z��(���ܖ�Ѫ&r#��d�ċ0e����W���˿���zsW���� W-�G�>7雥��Qܘ�=�>�h)w����<��4�tj������ܹtHW$j��Dia������:��r�p{��+�jKJ�o�n[��첳��_��
z��@��`���R�5b4�EzwFgme>˔xT���w-��d�Ӧ��3�eL�7Gt��*��k�4���i7�[�e�����oBv��h�:��n���[�TTG p�P�����+��J���_t��ZX�����ǃ^x���9�=\�����MH�C��;Q�`�JO�L������2TQ�����f�G8�����]�U�J���t��P��*5��#S���e(�]��b}�ľ�o*4�=w ��d�� �+�x��rv���5�r$�7K�o��3wj�>�d<�Т����i�#�_	���ދ"�m�
M�Ll�7�`</C�Wo�2�?�Y{��$*��{�a�?Uȧ�&�����B=�CV�
m@>�6w�g�FL~��q ���EZ^:�R����:��i�-I���<�T���	O�D�E��-~qy�p��tdmΡ;(\8eC���SU��@�� ��A*t��w��U�2ذ�bVt>!\n"9!�,Z>�E�:m+���cn�W��MW��tN�l]��(�IY#�JK�C�dK���;�������J��0�C�Ma�^�h��=�?�p�B�>o��1���D�	����U�w��(���B�P=�x�3���*ɡ|q���{#�ZF������!Js&�<j�8�1,��J���:"���&�kH0�(Ico4:,Q eA$�$p�U@LA����~���������!���X��r|�G�׆��
��Yfu-`��~?/�~8h�P� ���9� �T��9�7%B<���P�SH�}�2�z�8Wu�zn�0)!A�H�C��(!�R)�s#m�i�|{���mZs�XV9\�R����f9�(�ԩm�;��$�7[hE����'$����c��}wY�˳�{ϻwo���1%�����D���o]���?2�c�[�V��nЅ�_x�س�\9������cW����� �,���!��*47�#y�ӘӍ�x;��x��S@�<ٺE
�:�ޛ���܉e� z_���[��}�-X��)Q�0�o��S��1�@"��S�]��?e�m�#JM�>��[�9K�J���	st��k�ܥ�� ��.�#?�N�jMFϭ���8���vB��U��F�����{�����z!U���\"�6��9���D�%�؇hp.5�F�ㅄS|I��=&/�������(Be?�ŋ���~��ѲB�(k��ӵE���C��1�|$����Ij�������8�`������{v��*�+�ѬD��%09��[�3�c�38OF�NzVf;��I���	C]���I�[�B�s�ړÍ`Dt�9���`2���m�,T��z]�6~�]�� 0�� ��j_�Zk�;�vc���`<չXO-�NA@o�x.5���6M~�v!DQS�)�[A5L��	Z2:ȼ��=q8����m޼I{R�P���m�y>���`�I@S%}�?�9^��,>Ȗ+��u]��q��F�*\I#�o'9v��v�n��䭩c-*TE�-O��g���q� g[����`���\`��E��Ӊ=�v�8��,AFK��k#�r �ڭ(�4�M��EN��,A�j�^Ryip�K���eG�����?�^���M�e9��סZ1E�c+����XQ��y�����ډJԋ��Պ�� �_\��c8�[�m-<v���/2D�fh	�  |fg�)JC�X��h�m�&�_埶����m���{�i��śߦ�L.߃��M��4�ٔD6�D*�*o������e���k���Ў�QY[�g����Fl�(���%�U�Z����{�1� I��)#i��әN)P�P��c)��]e�5�O^Ȟ����!�`�����HH0��r�{�!�`G�u�s5�x�*=�͕����K���Q�d*���4�B� �ED���R|J*{�R�)���H�_Zu�uo@�t�����rϘ�ҶO'�v���[�4��˚�B��s��Զ6�tۅ��PWkL=�Ӈ>�sDbim�ڃ@��M8=��KG�zTQja���K�+�@���6dh1O�h���n�l��7�( W�]%x��۬��K}y��k��rܾ����S��U���'�_�f�V`���|H<;G�c��=&�� T���ju^�Ӗs-^��*@��P���w�9{ jĚ.+�w��6��ڤ�omns��.��|�#�e��L���H�'�q�-��*�ɶ�k"R5֋���F�&�v9%��=:��T����)P|��#Ǯ}b��۞'�rY���u�����e x
at$�i�)������I��ǋ��\��b��N�WK&7=X�^Cq�W���tr?<�Va5���7�М����\�N������c��-��-�i�X�hwէ��^ ���p���;#&�YȀI�_�D�E��n"�c�<��Ğy��);�G�#W��9$���+�`�Y}��Yq_���n�Ƥ0��{ug�6P��Ok��g&v��j�s��11��a�e��Y�����U������T�`p:�K�>ym�3��+�����x��m%,�����!z-�guW�v�9A$u&h�"dNM�����P��v����oT�K���HQl�D:�e��t�C:�7̹�7U��?�M>Rt�=nI!�2�UBQl)�����[�c-8�i'4j�6��4Ǥ�N�'B��'`�8 nq{8!�~2u��y�:<�b.���O)�j�qP�����G{��iV_��|)͏y�z$\ש=����t�Ǚc�����y��^�U�ro�5��0 z	�_-��,����u�����$�񏶜e���g"[b��e��ʆ���52�q���@�U?Հ�L�<HM7)z�^����U����1Su�b9l#l�'��8�ym�t��d���H��jשdA `�4Tr�j&��B�ƙyS7QBㄈX�e�aw(�n0o�X��}R\�O3��}_�0IC�5_^Y�0��#�'�����������Dv�Z�$��l7��z'���n�NN�a�Os3�%+շ�f�9�ΈnD�#{3�2������Q�kv�o���H��� �Z�%V�v���Pe]����;8G1~��%�"F��ֿT_�E@��˫9��K�}�K��b�L �v�]&�3+��WJ5P+2���V�:�^J�_�w(4��B�;��	T;�I�F�b����qO��_s��a��M�f�!�8eI~���.R_�B�"i��m�ͱ�����0�� �n��M� KX��UJ�9��[+b%d���1׮n7"���������̵�4��e�q[
{�i��}.'1ʹ�m�?�k0��)R�cb�U��J����������d�)�|{\��B�f"15�K[�(��q0���d�LT�����^��z���@ù���I�r1ZIn2�R��yu��/�ˊ�.Ҧ�w^��}�*�u���8�:����&~������@17�TW�j�>������Q8`Qu2]%���i���U+с�ay5�������6}���eT�`q5BG5dF�1�O�A�O�P�]�>����J�W:wB�C&�$���|~��}����~H5��H�f%�;��H�[�G����6��7��,,0
F�ˆlv��F `T���O�	�J,�