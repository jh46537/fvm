��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8��A��t��
�]W˱�ӆo �4��T=zZ�}�a-�Z��6`�Mͱ+ߐ�{��������?��LJ���ϺQ�9O�0`���J��9>�66(�P�[��?9��\rS�\D'�e0B�w����=[3�%R�ț�(����W���b�N����c���0Du�~S�v�h��{�:���[&yrYeQU:����R�Zf&�D0�@�lQ)S�F�k��8 �[�{�i�����4?0~���#^���Œ��M�Obc2�8BW�<�!�Y�^�NL�e��٩�,r� �ܙy�I��A;;&-R_�~�l�M�3ƥAUL��Ny|��8�ДaAa�;7N���������"�N���̛pe�rͤ��R�%�A,�$���:��}��*�_==�m��r����U�t�v�H�|��%��D��v�D��sY�Ui� �-�G���J4��%�u	���>0�3l��G���b�D)��A���X�5�{�´�]it�x��r�ъ0�&Ul�|�ߘ�l��t���`�75�1t��a���uj�0��`ۉ\vk���$GrTʍK�/���v������Ҋ茀�b	ri��s:[ލ�6�I��~�r�8ـ �w3/��W�ؾ�?�]�tw�/݇d�=�؋\)���{O��K�d(�H���t�.�9Rėf��H ���ڸ�x��̿͡N����������
-P��eq��'lMm��C��-~��$YH1�R�9÷�^g�b�'Bo��&�z�WE�.�Oq���" |54����bNZ�phR6�sG}I��p�(�'w%rO{�D�#Lyi����ax���OM�*�dfhK{*ʙ�+㒛��j"5Q6|�ˣ'�"X�E��ʮ��lK��x�� ���^7!�s��
��s"�dS��W���v<�Qk��+}��f,ݗcަ��3��IѧE��ʷ^�w���O�-B�I�P�09�n��{�#��2�F4���çv9��f\A!���B��lpvV4�<�:W�8���Vy�A�e��Vӏ��?��m.01�h���੼~6�Ԍ�<5/n|$����C�J���_3N���Rb��3DHH�?�[�b	����t�8�"[S�FǨ<�H����}-�}��������+O�g@�V��]�e�b�}	gľ��-��@^4ƀ7+�A6	��$sT���;�k�5�	P��Mcm���{�7��?�,!#m�e��*�y
&-M
�#�����y�/&�T���3h�,ʛ��6O�xބΒFd���[~��i�z�Gԑ��y]�%B~ލll�����/z��q�#_�gѨ\�c�C�2a���Z�`���.���[~@˃\e`�D���b�-��SQ�6�S7 �}� �%��:9�E�910��{���E{(,��y�d9B����Oxii����N$������>�&XU�}�JT��#c&yA�� ���H�ͫ�c��ޝ������P��EU��S�d����~�#۾�	��)e�WX)'k�.�s/�]�kr����ƾX������|231[�UA2����e9|�n�cy�����d�$4m���l�	%vm:�Ѳ���"��ƶ�Mkw�T�;�@�D� �3ƌ�S{�=j���m�:}�)�s�{ƾ�eV���E�ȭ��3(ơ`�!1�)')���mEe��J�d�5q*@��d�eK<{�[�:42|�R���i���h�H|u����N�
f���}uĉf1Q��~w(]UI"t��_�?�����>���}r}��R	�8�b ���-w ��i��e?0R�z�$0��j ^~B��j��d@�4�@���],�Gޖ�>7�ǘtT��F:��/�%�#"Hk�W�U���������ǃ�{�T��*smKF�����6�	�9�Y�	&a��R$vR��8]Ia��3�ڽ�#��xA���mj�=�&­"Ʋ+WF*��	��?Y]����nH�����k��*sv(�%�	H��e�3Mc'o� �ݚd#/��e���