��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ5,��kF��#��o`�Y�7W�?Z�ҋ@���JX1dS����
��57~V�q=�]�f3@��|����#�F]�$ר_�I�A� 1�'L�:��DC޺�U)3�ܟ�bnQL��Gp�g�:�4\Z���3��c�H���E������m�=��]%�H�*J���TSۛ����vy/m�JJ���\帓�È��1�r�/b���n�܈%YP�pί*�j���w��,6X�:���E�"j�&��j�6-�$���a��؆g���/��R��g�>6�:�W�@��*X
{��7Ż�u�l���T�\��7�&���a9"�1:-z-o��3]9S�,��po`���W��H�P��&��譄O��U1��@�f�"�=��B�f�&~��ZN ���^���A�`R����&Շob��:F�o��C�%v��!)6-ä�"GTz�G8��F���@u��"�����M<v�nY0���yy�d�׮r�).tA��;�f	��ܺ��4pθ U�	�S+��_�ɗx�X%�����⯇!�I���`AI��p%(�]g�Ï�2�j��+|!2PE#������o5��cu���1k�m9�gU�HgF(�q�hxꅴj)-���>�iʜ��fÔ��K%1�ԿʪJ�@��/a<<%��L\���,��C�-Ẃ�a$�
�Ƀ� q�E�H���p��Kt����{1}8�u��2����ܨ\�~b]�Q�xA���^'�<m/�_��#xs�B�&U�L�(�ء�X�Da�ab�_�U�!�B�"�_^�#i�xG�H�Η:���̰�X�ͦt}ѷ�=�U�W̬wk���+I�0��0�)���X��KH��[-�L��lѧm�;�z��_<���,w���O��߷�?�[�[�v��)��5�L�:�pJ��>
� �A��YK�[��){D�
�᳿iA�U�l�%Lp���h�j���< ���x֜���} �!?E!��]1Y{7ҋ�ng��l-gT�ޞ�>N����
Mk�k��ۛ"Yؙ�ux�(mo�f4d靟�i������rJ���uM%�?������O�=_v�����J����>�!�M���eD��>���̢[T�4�7B�sL])\ ��hGtH\?��S�]r\ ��\;��(�d#�bL��+�7P'�Z�E�i?�xF��m�.�\�*!��6-�Z�ۊ�����pE)���y|6|��:@�6ϗ����ۈϪ	�pq����;��\��N����s ��MK�~��g/_~`|E��J�{a���C�1@��SDY8�*  k��Z�7/b�4n��f<Gp�����J���dg"W`|�o�o�(���r+��!��a"�=e?)��3����f Ι�~$�x�T;��e�����)/'{�,"�#��/�]%���e�e6�#�,�~Q1;̸q�{0Q{�75���HT�X�"G�?u��#J��F������of�e� �Y�q���!2�������A�|9߅*��F�s�i<W'M��١�X랠Q�� ��)��͏�1����:\��,���g1!�������W�y�#&[I!/��؄w�<�a9����R�1�-��,i�D�t�����y��I+ng�,�����G|Y+�V҅>6��&�T�'�͸
�2�����T��_*�Ԗ��ϋm�/�g)et!ї�O�u)\B*�����M396�5k�
��d���G&ƶ�5�~� ם)!$\X�����e��h���N:�OE���,*vuUc�eV��iӏD� ±-��X
�\����$k�)�Y�%��lsoG�*�[MD��-���������)�O�ߎR��z�F=g�E��{q&vՅ+.��&���i3`V ��L�F?�ܒ|�c��)��h���B�\�*[$ �Kq�w� �GM_�z'PI��ƾ^�M�	Ew�n^���	���T,�f�XU�i������� #��#*����wFzgx�"��J�������M�n%��|��W"�bްi����gi�%6}�M�K��B�覶e5��X��R��H4�E��<3n��K�w�&Xr#sk�R]�D��e�aY��WR�S8�L�!2�v���nu�����mM�'*�j��ó���w ?Qq7����Ywz��z'�k+V��q��Vu��3�r���|�*r8�c�I�PS��5�_ѹ���(��Z!�����ͩ60�'�Gx
�i*��j��Y_D!G/�z��-�yѱ�SQp� F*���)�m���Qf���)	��(�ݙs���'��w����׽��[.w�o�|y�܊�'c����&�
O�O�h�S�A�9��-�_@���'�Ͷ��%��������_�n9Uf�3B+���X|=�5��v-*/��(?����pq������r��I�E&�F�g���m�+<e��⇪�HK.D������:0��˫F��U��ҭv�ک&ƫ�@6�2v���Y�V�*z2�:�C��A����;��vEh���u��u�S�7۸��k�	���S�P;H���zLBE��qj���pm%�]��2tu�=��G�#���.�p{��ፑ|3�6��4������d������,3U�r�QL���.bG\�37o��Ǘł�~3�e{9����>��$re_�����YkRZY�(ϰ���/틩�ίV�y�u1�ya.Ur7�R45�jˌĕGB[`An�LFOpP,�r|���Y@�$T��V�
��B+^V)4y�q�k����Aks7�e��I1�*U�h+8��$t�
)�� 4ɱ���p�]I%׍<�ݽH1a���_i�KЮw��zϖU�Y��K\X��$���a�}����*��C��&L�O�ax�!��2b�,l3���טuX!c��	x�$�$5�!��!��eg� `�R��|}�~�������*3�>��,��)$�H�L@1|Eh��2���*�~c��XW��@Yq�6�'z��u��i؇���|�}:�g�B4AV:��kx�v�G�-c/Ḟi���*]E��K��4��z�Sj���� �����@��&�� 2��x3OQ%��o@R�[C�^f*?�XB�$sY��|=7��G��;�NYQ:!���������l�m���6=��&�Q���@I�sQe���\�S�?p�@��6���[/��h��� Zd��$$W����.�E��Q:��2�@�8��c9�@�j�y+(ƍ!Ɂ���	f���X���s���M��&z�56�OO�?Hy�>�]����OUH�=wic����E��=]]� `��������H�i��A��hJ4�k4ß(�HO��B ���V�����߅K^�<��v��@S㗅x�R'7T�p7
s1��k��� >����C�<�qo��q�җLp��RHwr�^;g/���j��(������R`?�e&�[���ߐ}��H(nI�EU�'��oRJ���Hj�^�dL7�� ҆B��-�������y������B�	 &wn8]�!Ml=A�R�����*�h�2�wN�_pw
����n;+��C��F��K)Ffm��Mm�4�k����#����R���� J`�t����B��+>Ý�������h�g�ݧ����~�����U������c�I�:��U�U1��,�_���MNԫTp�M&{ix�3�I��0z���bt���Z���Q�O<���i�/? ,$I!}����/�h�G���Rm���'[̧�Y;q$Q���_a	^I"�������/x\d�b��D+�">a�y`C�bR��Juj�M(�Ȭk��J��̸.�f�7m��*�mDgAӛ߻���M���vt��td&�*�i�X�/���y�g��6�D@͵��K�x��ol@{k�6Z��:�~?�_�
FF�!�̺���-Ģ�O�ib��r�����z����⸤��u�:1a�:���D-��꓎�_��Ydd��x�G��!֖v(\�Meh��RQ��m���$�;����0���$[FHa��8�Ȫ�*5������C4�����#1� /���m�_|6���w~�{q�x�1N�1�Zsٰ���O��v�SW�|Os��a���%�?���@Y��������К˸X�A��D|�P)][�,O- �g��!��W�e�1R"�Vo������삆#k.�0����(�K��}��,��+����`����|"r�!���6C;$���W#�ε��햕ªӦGX��L��U1�8��+C>�bC:��:�<�[y���t�Im��5�z�����h�)2[c>Ę�е}���R�*��uk���9��^E�m����Pt56�����;ZىW�dO�'k�}h�f�)=�<�2ѓ����C���g��x�H�<b���R�rټKC����v�A;	�[FM�9+;H:�ާu�7bͮ��N�jeW�3G�?rQk}2�����	6�F[(�k���˒��n�.;�����'�q��)v�����v��NM�1�T�|p��bAM����ʠ��z\r@FI���Z<J� 	\W����t؂�k���:�X��e��ǙL���(�Nm�	�e5�h�XD�,���� ۳�K���N�Ih�&�"^Vd�9k�e���{�y�&�߉1���ex����4�'5����:�N�;������,=�%��Z��ƿ��ty��d��v()Sk��!Ŕ��2�9�ԯ)G;Y��G�Өg�f~��fFӞ����h���=+��z���?ln��*�'��Y�3�)�����#% |``ҙ���~Y	7)��A�&�����?^�A�n�F_j򼽃��߾�?4C0tٌ�ԫ�����1���
�	���A��=ԞG�_�n}�V|%~�-�s�`�W�E
��D�8��8Q��kO�<���3��?ΧI�C[�c�n���T�Sة���ēm�e��3
�El�����f�þ$
d/?P�yz�_��x���� ��:d��0��(�D�i�6�e��}�5m���\=�j�Ґ�[�&�,�)�Ήڿ��u��>���h$2v�J���Dh�������,b��fs�F4���N�ֻ+ER�aGϬ%��0�=	?�ZI�aA J���=��������g���3F,\^s��$XF=��n�� �9P �^�\T�������%/��x_�Q@�ɖf.a��7Gehj���G�{%���A���>���,��~ ><��I��xg��r2+���Q�e�s@�k�7Z��$&��}��7s��/�$uI��|��),���)��|�2A��� ���d�+�E�":7���?t�fc=�*n���#��o<�t%[����b?פ/�wg���ȣ��.���E��ܗ�t�&IF_[c�!�xx!�}��gI�940U�(s"��R�E���D4��7��T��9�R+�uN)|Ԗ�� �b�D��9���S�R��'�46��ͼ�'��2ZPG�vUi��OD�W�b��������+/�U��k�[)*�!�s�wbT?�1���*�=�}�(c}�e��h:��L����)H�>�:A�*����T�}���l��o����
|��Zu��}&Tr�(�ֈ.���T����Y+�s��;=���4^��"�Z��C�]M#ʼ��(A}�J��q#�R!�$��bFȆ�u�!xN��?�O,�ˇ��C>�4jM��:)�:��Gn]����HL!��iGl8��o|j9U%%�r.2b�� �4�_ykN�$����J6@I'���$�kQ/%��X!�+���a2�4 qƘM��BԨ"ع���}��u����bA��Z����n�7M���?>uzK�W�^�DF�'{+~_��	�9D�tV,��;Eu1Id�t���(�=	܉�<@��kOA�C�gWS	
���Wd�d���IK��V�:&0��~���6}�� �=���f�"����إ*�a� $?�iD��,��ib���뫋A1΃��߆dpf��wpuJ(�T+�\q�Ѯ|�M�UX��O����;�	��Z&EY*=۶�vV�S�J�%�����Η�zJ)Fo�/���<�<�`<J�z��SW
4��w_��꫏�n��UX�=�Pi�
X�G�x[Þr�tTǥ���Z�*���?��;���	�5�����V����?�,k����OA��'?kr!�d����wG�c �ɒ��
��dQrR�'s��G�5�
��ǰ� F�4�ӹ����1�+�CC�ơ�&"����^T;�����qŢjN�Ʒq����	+��}�u ݶ��m5y�U�ݧ�Am�'��,�~�p(�E��K|�#X��+/{Fq�,i�9�!��簯��+����$;:\	kLV�3+�}�l@�/I� QN�J���h�d���T9��cΝ�2n.e���?#]��pU\�h��3.���F`W�� ��t�[��j:��������=�E�6l$rd?�v)�E�۟�Mt�t�T/�S�Z�����;P;(�5�v���^�va<g��[W���R����#� u�#��+�9j�fqw�cm$��q-����*�U!L5�~��nt��IGX�-�5w~�����S�|O-��mAnޜ��*�Y��xE*i��� 8L��� ݡm]c,]4�h{6H2c1�r[*�aa
�mYU��D��ځW��t���|���n���,�b��z6�6�,i��G���b����[�De�$���������h:j=������ZM�I��M�����VSu��&�TK�z��y�!�~ݥ\�P��.MS�l/��%��EQ<�T��؎�>7������(.���$͒|�hY�!F(�rZbz� zK0��ȷ��w�	��|/����掐�i)���������E�����A�#(ox*9z n.����h���ZR�Uھ�*w�[��b-N)˰z��6�U���ss�#?��V�6r�C�(u�x�\�C�'��!T�Jn�6N��#@���^#.~�[p?�J��UR+��!���b� zzm�2<v���V�����5�w����]`�gM�nl#�k@��Vi�����<�0�NR��RUjϟ�6�[s�ƎQ�t
��"W�S���ӊ�"8���{5tP�)��奊,���Zw�)wx�8��Ze�7^�ΑzL+>@dW�+�)o��iM���IE���ni��@;[�>��b�KAHoZw:������CQ=����d8Ƌqĸ_F�j,>��)Zp)+���(=�c'C�T	��{��l�u!��H-�|��>��10�Kt�˯���R.��J\	rH�R��#M%#�MgZoh+��!�d�����������̛�*(Q�v�D��KS�������d����k;��� �)��|��0�è�I���|�;�k�\�@�Ğd�1;��b�/V��?-�2ݹ�F�D��J�m �E�dNWnW_v�oqV�QO?~�ԟ_�L}��\0{�ꯟ������\8׷~�~�~���>�SXw*��ةN�w��v��W���z&d��j�*�p
��}*+J=#B^	����}�>O��ʀ�K(�5��W�|d#	?�xR�J���t�o�O����m�]y�F��B��&�0]IJ�Wy�{��I�.l�/I�;^ls���I��P����w3��j��P����9I����Z��?}j+�1y��Ԯp�����,��}���Oeq@Q�j*!Fx��"°�עɬ����|�U�v.�= �t�L�3���~�>a�׫g��Z�T9��h_�aԦ���狽Z��H��o��R��* (G�c�U:��%;����\)�S����uoYS@���C촯��J�R��f�ٷ[_�WiC�8�//��� }�zx4�Ly��]v�����n7$����P������SA�|(B�q6r�-o�D}FQZ�Z�?��fl��˓׃��:�]0
���� B7���2�j/nlv�)E	/�QĈ}����֚������Y�s�Z�1Y���!�Y�O�b/�U.��y ,��a:�VV9���\֣�� � L�tk�u�O���n��~�gC#��ɚ�߻>��ޟ�5`���>�j���#��%X"<	*��bl�+�dgB�@^�{�6�`v���D�YZ@��J9.b�P�d�������RA�) ��:�-ݑ�|�����A@^L=l�jWh6Ô��7Gʍ&c�g퇻o=��ϕv��_R�H*�S��b��MLo�@m���Q%'�k;���j��������D����x*�t?r9;�,��%���\?�F��O�<'�@�d��[��Й��i��	ۗr<���_�	GkZ���n鞼<���mmv��0�E����O`�L�O���ߨ��n<����9'P���;88�B���O#p+�	��.���M& "������[X4f9����]�
@6k����|n�)�|����IC�' �î�qMq;��5A�MBk��o[!�b��z��#H���������8�"�J��(�Zaq��H��Xv�t$�4�Ꚃ�����l_�8FvT������.N
^����1:9C4Ǉ[�����#�� &A��r�2��T(n�u��{@�/���K7�b�7[d�A�e�b�]FV�T�Pa!���ng>X�����k�ɍD]z�(��E5���2��/0���4�5���D~%w-X��S�9��a��������p�i^(�{Dzz7�ä���]O�T1��q���� �I$s%���Sg�۶��%G���`�V.�n�ް�Y��*�k��l��O�mtM0Z�հ��IC�:Z�)Ӟa9`�{���J������l"W1�^3�
@q[�̺^�T����:�M@���Ld,����O�����j�]��y��Y�(��Pngt&��XН-k�bE�2ў����O&|�-B��O�Tڝ���&��=��"���h�2V�2aS��g˩8o����iY?�&m�Ed�7 y�<�y�bWL��&�Q����}-��.�zW#�=]-Oa�@'�X�>;�*�
�D�z�=c?��]<��za���a�b�����e�אC7�x�$9P�͂U'5�K������8=v�-n��$r �\��$�[g
�Vݦ��ڈ��K℁\̌���H2��f�
�V��	=����6��5�'�Qdg�,Q��G�&"��pa?�B�w��zGjN8��|�Ѝ��}�;���Y�œ��h���Gg(f�Bb	�B)g���"2���a�CU�V�j3��t�T�o΅\#�Q&�ǂ�����e�2˵���T�d$ӆې� g���U\�6JC@�\��Xσ*f��Y^�r�%e��E�}8���L��1$�r��߅�8c����N�v����u ��v-WrjJO��2/�۸��%"]&�E4��� <�鷼�do$'jrT Zr�T䵯df����)���[�4�j���E:�N5�8@�Y�5����2|�P�C�W��`X�:���p�(� F&Z��d��x:�I�ip5��CB���5�kA��gN9l@"���N���O��e[7�������\}N>�>&-f�'W=!4�ߙ��xN�YPCffW/"�\B����|v��wrZ�R(}�Ј���Yq˷�ȳKG����A��bׄ�wl�^�\nO�Jq�sl#Ts��ڈ�k���ya`�k�w���