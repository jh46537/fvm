��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"�.0�у��u���D��@��'���Uú����0�"�W3�!��N��4��e�����M�.G֮Z\�^����#���w Fu(#���E���j&=_�/�j�����㩋Ҽ8ܞ0��DW|����1#F������~"B���%/�#��Z+�G�!�%'�"'b���0�:']��P�G���,8J������}C�Cn ��������oSZ����>T�1u6�b�`�i*n�!	@[Ap�O���8�5��/=�!k�W�5�q�(�J� ��c:G��q��&���8�u:=��W�#�@�r!ǉ5 �b�C_�g[�I�s"rHdw�M���&��Z�!�/����dJ��y����ͽ���Q�;v����{���"VM�P�(p��,������֧7@)�
����/��	�H�T]���|�豂�i^-���6\��)���ك�zҚ�q�ٶ��Qz���0��}YNHܵ�U��t&��bp��$�5 ����O��jO�z�k\�rͲ��?����T��XS�r$ؼ���~*��jF�!�]g����v�^�/y�+ȖS���$��߉�-1�ah4�z�$}�>��Z��_�RR��»~i[�7{p�=�3F(-�2JOz�)��"�˭����[@��(m�V�"tƥjw���7RC�XՕ�4��kƎ&�z���F�6�hV.4@X1j���7� Q䙿��BIr�M�)oN ]	Nf'~���l~�h���s���}�پ��Q�k�������������fS�鴩�<LVD���o�V~`������� ��P�r������uD��ʸ��� 2X^�"��*�B"�9hjI�zud����{�ep�3�$��
�L��EýP׳��X^7_����2��}�(5��Z�����*]zG���֝s[��C#|Лe`���Z@5�#Y^<Fر���F�9��i��I�Ԗo>�M��������k���8�d��|��mȖ�v.�p4$�=O���Ouq�N�#����_��b���,�A���	��3��iQ0>�<���q��}�r�Q���g�K�S+8��)�X�K�s��@��U�ᄆ�d[�lDB[Q1�E�#H��>�UCm��r`;T�ȯ��>u� ���Ee���{� /8�S����ش �l��Q���VR���V9B((�D�Ɇ���Q�w&J�O_�d��1���&�%��'���7��,�0C����B}�_��b*f�E�E�&G�:Xj��I�[�!_��B�z?7=l����-��c���F�D��_�to1?�&ɂ>��6�������F�G��z��o��b?]�+ڊ���C��@w���NY�P�g6�ӑ	j:�M�*IA2H��w�@`��_�4�ǟ*�4���[�q�n:�<�7RɁn`��̷��g�L��"���/���+��F�_*g@eS����9ii {��I��:#�Gl�2�[�!Nɂ�����`jg�~����]*ц�'\��,����'�� �� {����~N���Q�Q�gQNlu�6��_:���·{4����yCj���8����oc{������j��`���X�M��+~�G?V��7K:��w�h�@l������ǬeZ��Bg�&�#��f���:�+�,m�y��"S:��~���v���^D�p6(F�9ឆ��W�����zQj`�L�ͼҋ}�r�B̽L����\͇�	!���:�!���}����q.Z�a��&*V��e��.���l<7����0�e����1v�C�@�Z��0:���c�%Z�3kz�����6:M���|T����� ڭ�\��#O��M7r�c0c@�ф�8*>=�[�>�2.������3�j��DHb+�
j�
_�P���5z�'�4���n>nu+�-�b�Tuk�H͎����qzK��p&�ֽp��8˲�O�rZ'W(��I��8^��Kr�HN�(7Ra��v��҅�@4®��Ĵ��LY�s[t�l󨊟+��_�R5��8���'����o�)<����r��z���+"q�M�o���O�{����������y	� xD�Hc}���#����r/Y���Ɇr>ڼ�8��e�Ȟb��+�� �L�J�}��������N*��fVuW�U�<�(ZL�>nǉꥻ/ӅjI(�<^�-v���py��$� ���)���8���GC����F�ؤ/��;\�������+ʖ��5�
��<��Ex����<+�=?E�g�7ۅ�� �VN/;��3W���c������y�(�.g���"P<����o�V(7�KGL�$�)���b�&7�
�.�t�a�����<Y�mR���`��r��h$�Z���7���;^�$�Rg���y-<��]�8Q�z��BY����&���<��Ct��`P��V�=�QǘxE<���趴��P2て����<-�.%[��g@� ]@n�N=�N�b��>�b��.��uL�ΟuB��7τ0��yz�M=��eM�~N�F�3��rƷbc��}zXL�u��j�d��Sp��F����֞m=~�p��-����q��I��l\ɷ$6!w�Ĥ�K�)�=G[.���/~?)G��@^@��?�V�1ӑCsg$hM���Fg�x=�-2�r�մT��jD�:�(UǈÚ݅�υ����d�/a�(���n�hb��3����_���P"��X�E��=qS��t��9�+��֤���7�ʙ�?gt�I@I�%g�'�ehu(#v�H��3��*C�t?M�N(�dWj���>§��l�+� jR��)�D����v�� f�Tb�m]�ѭ\Aϵ�M�wb̅'��PF�a
�AE�,�K�I¦�w������Ql�a��Z�Rq�Y��pyy*v����6f$~8P���m��ΐ{��Q����d..삀o�����6f}��%��v�)�Y<t�ȁG�
���!�T��P���K���6Y��(�X�:��۞6f�wf[a�s0R�
��F��@6l�bg9�#ܚ��]2�N/x�~��!'m��p�K�t��y��M�qP�Ak�]����������`<���ɠ�2z���������g�Ǧ�ڀ��x�El;��Y�z.1��f�RR�>����LG���u���N礆��ej��ɊT�CN�G��:U�g6�].#�܁�Ӊe�4���,�Z���6�8������d��_�6u��6����t�|����ToQ�e�s�y�Y�᫳���᱂�%!�g��R�g���<��jM���6I�^2ucf�r%���l]$��:���I��H����W�������x1���sJG"��w3�^tP}�KZ\ѲbU�8UĉjzԽ-��N��-ɞ���A���df���gl�߬���JŘ�]�\ۋ��,�Q&Y˷�|]NZ�㐛(s���;���lD.*q估�+���O���1S�@���c{�,߼��r�$�Q%-C�˥~]�^��)*�5�鲷S��"�p+S���J?͸���%4ց�������
-Ȇ��'�Dͥ�W�?#�?x�GԄk�1�,q(%F�9�����F~nʊP���k�Um���I�\���0f������,��d�D�0R��
*Pt
F�Pyg��G1�N�&J���JX��=�+��1��63�1<�x��#���骩��+�wu��@���Wϭ�"�|��xc�����_�԰�9"�,�o�����ͨA#������I\�鹄+�s�D��
kUJes���,]1��Z>�/����6�������Z*�����Ϲ�x$�]�$�<ǉ�k������#�{r�Ѭ��!�r�& uq�e���:�i7cWј�/p��\��b��,V �ШN�~�P��Z3�Lc��ۘ�ͯz+�S�N�j�~��G�����Q1�Hͨ��r���LS�1�4E����.����l+�"ly��7<��,��`��.�Иka�>���;�9��RȦ�I3K�=�V�B�WM)L�*���ąre�;o�y)T!^�A:�Э�U�RJ�T�D�i�_�YV!Iw��Fh�haT�!�����s�$W\���wt^������-�<b�?�6LP�a��W���xvn]87 �\FT	��ţ��[�dr?Rzt�nj*��\�E?rR%�^�`����kT�
Fq)lg�1�h��6L	`u�D�깬�s��q�c6Oc�V��}�ٸ��r�Z^L+J
��L��U�HW��tέ�w���]�X ��Yc���P9ӑ�z����*2�J�R�J�$�ǖa��b�Kh� ��O�f �e��<|�;�z�C��,)��^��H_�ᱟ�	�cC�#"���"SͼL����ꯢg!�
���;��ǘM���X�*璛$N]U���ը� Z^��OW��� 59n��Ӹ>�կ�s���`�'6g����Ij������j#V7>��X�����I�e�|rĪ��ػD��[�XS�%ve��[��!�1��9UnO&�Dd�R�B��Y ���˳]��4���;D��]�.[��G�O�ς�W�'[!�w��:$#��O�i�W���� �����n��al�>��6O.���If��*�}o'^Оl"
��	Չiq�V���E@>w��^q�%�N� ύ����5�j���?���V^ug#���tQ��\���Z-I���EC�c�٘�}WFh�+~���,�(D�x"lm[y���p�쀟7RDZ�qty����m��z�4�JU�����"lª��z���_Bt��e��z�c��Vy��)�ޝ��k"�v��z������f��ļ{Z��
I�=���������q�K�1�|��9?��\8�[
�g�=�.�|�ń ��LÂ�e�������8=�Z��1?�@��i,�F^����x����S�(c�N/r�N�I[A�M��N�3�9ɭ��s_�?z1�s��d��p�98�����iH[Nj�w_P=q�4`'~������GC�r�ߝ��{F�	 C*���)!���l��h� Z�!�!\��8=��� P���]�BJ�uD�Ϩ�)�n�>�z�|��3f����-N9l��gܶ�t�#L4�y<@�1���o���"�
���=Ro����6�b�!�3���ZN_�x���[FvN5���I�20�����~�