��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQG�.�����t�������Y����qj���ߟ�Fz�8��X�t��ݙp��-���ܷ��é4&�	Ř�%���%"�>�;s��Y7�Ȓ҉�e��o(`U�WA�]ܣ��K/���u��ĀZ��� E�7���$�t���A̔����K�eT����iP����⿳�K�r��n�a^�<7� ������1K:vC���6�)K/6P[	:��4�ګM����O&�;���߲1p؁W�ɰK�[X��+���%L��@b�v�&�����Ő������V�DZ�n���F�Lص4�����45��O��uQk��VƱ�wd ����1]OC��*��RY7�I����2�鵣��~�.(��x�d����2X���\u]��f�**Xw~�*�ڋ@	����t_��́�3ۺ�.�0I�w����˧N#��H����;5*#�9�i���p=2���l��ߗʇLY�J�p���[
���s��aT��DT.���-u��,��n�&/��S͹��~�!ʤC?2S�If���!A����E�z��ưގ%`��� /b�^p�wi��i,3,�7�<�S�vMT1h�z�OA���$�9�/��͢ʯ�L�&���)(�yq�^�4��J��"+7���	��&�l�(�E�٠�[t�2ݔ�8�g7�F��k�X�,Dꭥ~�]FBF@r��4)��l i�����\pwL�v{��V���8#��҉������~A�-&�+r������X����&͊���^��:nG�T^�n3��ʮǾ|߮-�x��g0����s�q��L5lr����f�C���?�Ah���G�=~d���Y��ӛ�V̀5�Ed�6F�7��]'�n2��ƈ蒿��q~�}G�� D��u����Ye�7�����.��<�<0�����J��Wd� ���{��tH�Q���2)����Չ�m�]��jş�"ƌ�RK�D\�X�B��!�Q��_���R�m���嵐8���i�v�1��p�W��0ڥfHt�VWs�}!�c�-|�/g���ܸK�8=�����6G���)Z���r�@���G5��x���@�u��B~��������LX�2 ���x����S���8a�[�����=g�0�N�߈tt�e��g�:	��^[�:Bcr�O"��ˡ�f�5�k��H���p�=r�CC���+�.��$񪲁7���7 �ȴ�x#C.Sϛ������~�f��7�r�-��=��sp�db��KC	)�'V�6��x&��Zi,7��=�����9����餌'=�����7˴VC��z~��?��մ�ZrLl1ԗ��G�Uc��/��)����BE�
g��� �<���i!.�u��jZ�`�����n*��-���N��d�\nK����Щ�l�a<�	'd"�(?�o,�)�{��Ʈ��Q��������<��"	���?} 	�J�!�,D��:*�ңc�W�<X�pJ��}����c&ȉ�i)��4��\�j�==��ب��:77���^�KTd�����W��u}�j�%ZFV�8�Ȕ]��(9*s7��S�lt d�s�diڈ+�h�����;]3��a�Q�E�j�ؠ����E,j��v&���0��1�}�v�0˵��pimQ�؉��*�T���q��:�R�����D�	_��9��'i%ճp�9$f���Me�?S�su1�	���:�"������E{�|�D��O��%��y�U������
�+�?��u��Ҽ\�+�4��>�d٨�����aH� ��3�%���!�� ēܶ��v��
����?�hW��ܙ|?�S�(����k��v*��\C_9�Ba�z�b��w��a��b��y30�nj����D� �}��;� �wey��cM���0k�u��"��d��Ubͣ��V��C+��"U���~畩�@3��)�>%��f$Tn��>�a谯p�y��=�5&����i�<��K�\��z^�����SL���_��Y.����==,�2>�gjR�f��u�5�^LM�T�&د�9|�\8�8@Fp�x<|q���)_l-"ąŮ�Y����� m �blߤ�-]��!�oT�/�N���~��&�`"��䴚����s�r��"P_i�I��k�q}���������>%}O\��+�P��<�L������]��t�����O�8a�L0��i����S�Ѡ�Ksq���WM�8�f����<�0Pʱ�uƼU��)  ��۬e�r���&v��:=W�X �]�J ;�侗����:�2�<�lJ��#5��z��*��D��a���O�|��O�
+h��ĪG��=�����.�]���A� �Pv�?^��P������n�j3��G�����F�G�$x���F��h`"=<I��v��Z�Ft�Ȫ�Ze��ܶ��)�SPtu�:3�������w��L�{����G�Y���S{��v-�+�\T.ՠbP�U����f�Z��q��a��p.N[�dOM�������%��"j�'U@�~�W�^�����P�t��".��^ěo�0��S3�z�2~�J�����R�0"�@����E׀Ę������]1?ˌ���+y�w��+���D�;ߎgE;�%�Z���CŋF�� �NhKu�2C[ �;5Y���*GT��^�zPrvǨO(ی�����cIOf��/�5�&[�a!?z�іſ���U��3�(C?�dL)�5�D�5�0ȣ?*�S���f0�RDљ����Bi`�h>�a�0��B>+�*(�3�E_rNC/=� {���g�ݕ���M��,bIi��,�`m��{І�y$�lu	=�B�-��i��2,Pw�">@�,�'�����ڲ���)G�oJ)لkt�e7GH�_�+o~�R6�m�LkK���szKkjI�a��
V���v����o_ ���uS�k�1ʗ�"L�_�c,Wn���W�ɠ�I�P�C���T:dD�C�'d@wlR��W��F����)kg��s���B��M�Dn��3�������-ź7Gރ��?<�]]rÒ��ڛ��_���VGS<����v$0Z"��M3EK�B��6!Ǖn��o��ۜ������|��%E�G,�t'p_��VP�s���/к�(�&Ζ�)pE��c�s+ZP	5Ԡ n[����r�`N�˵�5����8�腩�q�i�.P$�S�ęG���w;��S����M���c.2b�I�:��5��݄�µ�ˇ��$>ͯ#����v�츲ůt���\�@4�ڕ��r,Px2�9�tʻ�����������ޚ���d��-��@}�o�i�G%���Mj
�X����f��������sB>JUT��T��6G
ӧ��
΢�;0�?�G���G���M�G��$(�ڔ�y>MD��H�T��}�`���1��Y�M�nl�Me)��
C�)��)UlޘI+^0α�b�^=�f�d�W+[Q>�\X�H�o&7«��w�C;�
��0�J�z�Zdߣn�v����n���Xv0?�gp��-���c,��[+O%���_�6���^H	�ۃ՟�E�`��t���r���w�+r�i����_|��=AHY���������ʆy�$�Yj���f�KR���B���fKP����,�	�9bU>jYp��F��:������*w����˪��s��7(4�c�h�,����+��p Ϥק|!醙�Ƀ0���	e�p+p|X��A�jy_Q�O�f�����U4�z��g*�<��jn��?���:|����f�����E�(m�d�E��Q���cdS��F�0��[5�\C~֟��k����S����W9�~*"�9�y������~e�(��lǺ��)w9�)���V[��{W�-����.�ZO� p�5�h����vq�����T�<h7/ຼ�I�i<)7��?P��t�kar��� YW}�#������x��~�f�I�p��}�Cq�7凳M��.�K�v��U\n�@�;�3�C���8���0(���O��J�ѱ��>��FT��N��>R��=�B\
�ټ*5ax�1렢 T�#�[ ��"3O��zm��Q{�V?����ad;U�����`X�X�_�q�l�����B��'̻��̓-�g��5���UW�;\Uh7̻!9��>�A�갴�iQ������'򍟕�=b������&����鍊���{.��O�c�z�)���x��9�����X��Z�*� �Sv���;x�����X�%3˕�?e�,��1�^�Y.@�ߧ�H��%UX�Jv�2/~{ x�Ze�����YW�d)��:1���(��\>@墱�P�Ei7��}��WYB��&z��]��xL��J43/�&O�������r ��(ԺW�k�"��e��h��H�����F���f�X�]������*�_�}�Fp���P/5��jSo]	�����E�=�^��0#v�,�<�7t�K�W���""(��k1�� tu�E�(�!���j���о��b>��Y���C�B>�T�C������J��W��犄���Me�Ҳ.����D$s)�=!Tm��W ���	3֋K�$hM�e��m �=/�����Mr�ԣ�0l�O�A{=��UgJ�ȯ�3v�+[Uu3!���4�)ʅ��,��@>���1���xd���S)3�Z��jc���D$�\�;�P�hDq���D6��'�������>.��<gwo;�L�4չ�]���;{���-�{�vaGZ�Yp%G�E�T�fȐ*S������t�W6A�A3�L;޽*�ؗ��S^��w�,t�M=���)qdT���~N�Ip�.`ݞY�,k3GO(�$�ێ�s�۞�rg���hmp�l����vf��롉�J Ԅ=l����^`K�L��ziRym�,ќ�p��u;B/j��;��FѼ�@h�S{2{��B���]̐K��d�i�_�I�	�[���o��lx
30�jp�� )-���<!�"(X��f��:u�4lA$,�+5K>L�(�B�1��tIt�N� 6���^*�eWc��-~Q`t��z����