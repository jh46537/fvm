��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK�Q���L�OX-����P@� �K���(��2�#�|'	8G+ǲ�q�-?�?������/�1�gR��ϛ���v�O�ۨN��r1�W�ϒ�&��)�tS�	=���o���E�������XP� c��>���-�;�OUp@�at2y��K��DҺ �̧VSk�)���p)S��nsQ\��N� 6H�`
;��dOW�q-S(o�w��.K���f`<�=N��lh��m=�������!o	�++�>��L���h�)1��{�qo��1�a1��
F��B�Ȑ����x��:��7;�1C���c��N��}2�i�F�{4��xUW����c<Ͱ�>iI��2�= ��s�L�H4��Φp>4uR��xy��J�I�][���ʞ�k2m�$�Yc�`��յ�P_/Tw��d�9�P��bw��M���#-<�;c�"��#���ne@Q=4�q�͞S�ޖ�9BTC����<W��S'VZZ�������(t⣇Q�n6�c����>��ի� �c"�y���ïɩS������s��s�ϑ	N����1�w	���en�,�\j����뜜�).�袨���D�g?�dp� ������W��9f�:g1q��nl�m���gQ�J����? �y1�A��,y=�*��'��]�.T�;�]38��HO�q��A��!�^��L�eqަU(��LBV�T׵Adu��C~ЛF���Ntj���ܪ���*�L}�X<�'=$tX5ܽ��eh������-��'c�6����D� �s  �sst15���	`.�
!r�m�j9�G��zYM��#�!�Z���Z�+O|�(M;��x���I���9}F��~z|e�Ք�K��%�y�}�.�'�:��v�F���-`hU�>F�~>]=�'���^VuX�¸�1}i��9���@]��zk���'�x�;�U'�C�]4��5O�V����0Zt�T�<
�b�w��㩳��P��f�ݤ^%��s��n���.XDZ�f��s*��\�d9A�SQ҇��ų�a0v{#���/��aH�m�@.NE�d��$m�D:\fVZ���u`ܽf�;�$ƴhwgZ�΂��R���.��rg㸑G#�[y�cAI�2�Ӗ��pKmy��o�� �|.��
]Mz��	��l꺦ĮE���#qM4������.��R!�v<�T�OC�v� ���ey^��cIi��${ɽgq[g��Of4"jg���Y����4Z~��v�O0Lgvl��f�)T�w*>6[߱-f�]l�n�!�5�ه�_nR�J�uS����t�_�����ۅ��p�u�sb�]U>:I��4���9[̇=]��P�[�o�`. ^˵qh
��_lr5����Z��L��HlOQ�6�N�B��;m�r_]ݎ��OZk��tM[@�� ˲����1Nⴌ��p�^���U�V�aw�g���7�_�8,ўL(�"�b-�v���bэ�%�;�����/_3�i=�ԛj�]�O������v&R��4�� �/��*R��|Df��#|�Vc&1x+���o/�FG��`5*:�;��x4��x5uu����R��нo�M�8� ��U�~��J^����n�ټ̆��%�eZ�q���p�ѯd"�B��l���u���\��=Uxt�́�n�U�&nĶmPy�=P`�*gfg�*ͯZ���2��a�;x-�������Y�aPtN�]�I�L��R�����������<jLC7a>�Q�Jӎ0������ӹ��!h��1�Ç��E�+�{��G���œp�V��?TV'�aF� ��}�I���gzt���}�.Q�J]�G;��gU�V�VP�Qf;#�s3�H{����f��?	ɣ��wĂ�Gq�D�K]��z�7�ߟ�ne�%�ZF�5�y��w}��
�h����nl[�bࢻ�ҡc�]ce��,�ӝ��=�a)
clC�6"d���^y�6$v�2� _�����'Rn�hC�B�&�)���©�>�>�Sq�O}m��I��Kv�Hj�������淲 q�&�<�xۡ4g(]|pq�h�@�����{�G���=]���E��}Xf��B��h�ғ���E/�G�Y���Ҷ��&x�q'�k���畜�nm�vőd��TtwL�@.j���M�W���p_��oK�������v5K�9FS�PS	�.U�Kp%ٳ��^gԫ)�C��i�|
���V�hVP����2\�0!��S
��{Eq�#���#C[�5�:�?��H�E�Q�i_Nw�gJ"2�nkS۩0S��Ѯ;�1�9;o��~ )b��0�Ӽ6�Î�R�g��$IG�Q��eMtBg���DS[��C�UR���T��֮�Cp�N����3�Q��jSN�`˪��)���!ٙ%^N����n���v}�3�ږ�� O?$���T���C���o�ūV1�`�P��DGH	O�;+盫�N��l�B
Ҹ���x�ꉠQ�W.->�\������E�)|�_ӡ3=��;�$'�ŧ���	P[L�it��qj<��!q������ 
���p�3���K�,�=��-vK�ZR���LSig�f�
VG�n��w'�[©>��Xd~ٖYq��z�5��q��H��`hV�*Av#�,�W+��{%�?��E�NBt��.6T�ZA[�>�4!����۽^��{08��O����?XME�.F�g�'���'"�����P־�M`�P3m�0�Ez�@�^:�6mLl��5Z����@s0�H:zK-�p6��*8���gi��2PY�W���Ō��n��9q�Ƒ����c^�|�|����fJi�}��F�H�?۠��K��(��6�+�1͆>�Ӊ�OBk*��>�I����CQp��j��I�鍝R&❃cm/��H��*bA�8��r����H:�%X�3���}�n� �PLG���!�Uv�c��U�Hr��������x�4DL������-�����UI��֍mtmi��/��<?�ZeԒ�K��}�ֻq#��=B7��P��и�),)�L^vJKs*t� CFe�*Xm�s�O	��ש������)���ʭ� �^�T�	�nv[J�8�bv0��ͬ	�S4��� $��j調��kj�����p�vg���iFgt�S�0�Rr�s�e8�=?��g}�� 6zk�-e
5Hh��~G"(u�	͗�D;g����r�WǢ�T���R�ս�uz����[�Z������~�XGW}>���Y$YjZT�2u��s]���J3�c���v+��K��t�«��	���O��)�蔎QC2�' �0w��=U���a�V��<��lSBGb�Xc�Qe�����=�M�$�p�$�v�-b@(3����]�x����&��Wа�\v��,d��c�\�^#\��!�hv���C�jg��)*��)��o�+d@�/A��aD��}�#ӌ���=�BXO2�����C��L�]����S��[�K���\!� ���`)P�	H����=�毺�Ҙm\ɃZ�q-A���t�Ad\�m�n��x����K�k���bE�b���#�&�A���y��zղ���|����L69�� �/G 9g�4�ה���S
�?��֭�[��i_>ܝ3|�v�ǾW�L�o�^���I�M�Տ���V#(��B�P�oRHx�db��ʓ���y���(l��I����8�D(�>�9��dqܔ��)g����)��'�m��]5�{F�ݣ��}�R��8J�CY�6~�i�z�3���*f��o���&F�I5�z�aR��,ɞ�T�u�Z����{}���)׿H ���[p�C���������l}�'pC=q��'�)9�� �����x��z�f���̔���o��	K��/�E�mSe��#�y��7\�p$������|�Wbt�n���������ub�O<K60��Q�Ax|p��bf���쏐�����M[ŵ��Μ�w���ZW��$G�P�m�c����\��PߛJ�Z�g�&	�L�	8�q�f�`όWd��dz��S��0���x:/����M��2!�(k�*���/�B�B�Ӧt���_���0��{E�J-�-<�$`\f�i���7�cD��|�:5�½+�y�9���I�xN�~�� aV���˪�Ԃ�g[Y�&h���V���s������E���-h�_*�8�O�͐�N�����9�B�Vq%Ax������ȺA����-���G�c��^���3#�9�3�qq��M�< $�V<Y�2�}�y,�4W*��:�[�I�_����W�6�?z�8�-��+0�fGh���șAwI�jX���"Fm�S�=���d����a�CG%�@����f7[
�>�I��C��h%�����������2�l�A��锜$I^��_���6�|QP���gg@FV�fDXt���{o�~Ti�"�Ge�Z�U��([^n}�;��S�
�̨�����<�{�2��( Z�a#b��ݥ��2Bx��2+�s��>�͂2�Vk����B����`�`j�g�h�I���5�V�q�	;�i���D �G�� >F�	�X#��� �C��q���:�?�i|���?+"6R�V���/����`�×�,��}�˟�1YX����\���~|e���\ys��+fs��xWh�J3�s�
W*�^�(�ےY`�P�R:�;R�U[�8��5��b莨b��f�t�̙�ʉ>�Pğ	{d_��/{dϛ��ԫ���E#���t<�y�D�w!��٬k�;z�f�@�a�A#;GSFO�z"o�.|*&f��X���I����ߋ ��8�y�W��>�"�*�b��ZrƔ��Iԁ��Y�E�6���H׳������v�G�l���������6�g�{����Î�;����4�˔�R��I4��LV͑�����%(D��v�����K�{{&������W�W���u�Ū��5��1�8���%7���m!��
'�E�j>��٬?��С�[��cᕵE旤�X��2H+��D�k�����Ї:x:cl�(��B>%�֟�.�4ԟ���0&��*��c#2�t��,2,H*�<@��㌐h�>�ҷ?�b��J�ɇF�������Y�H���r�;D:P���n�f!b$�Xmq�k0R0�����Dtҷ�Bܪ�m/��a�/�>Q�Y�YT>KQ�R^�W��sf�c���M��_��V���i��a�I��]��"�d����uwi�����
���"W�ǝ�j����.3�^i�f��{J��y�u���2��j�&�q+���m)a�8έ�ȝ�̗�9=Uka�
H�x�њ�d���~	�\t�ї̦���`���VŊ�63���f}�z��t�!�D3�F�<�6ӿY�s��U�x	d��@l�zs���P��Uچ��LGŨ�!7^���\{/0��b���n	+%��r,Yc{^R��y���<����:�'��	��:ڑH���թ���t�en1�$�
�����V�
��-+����Vb�E����7�n�n<�p%3����'�-F��*�G�rf���[�/��������BS��1�N���Xe�iRV��	��䫬�'z��ZZ*v�!zi��W����_?�'���H���t�Jc������R±Mm�YW,�a�D���ק�ƾ��`7�h^[fu�X�4��,��cW�_[�^��Kes�����0۷k�򮚎�WܣS�L���Lγ��k������ԅ L�岠P��0�:�HC���/���ߏ��*��54��mCU1���/������QsTx����44e��UN���u�H�K��b�6���`���9���V����S������F�{	���F[FB����+aK>o�YgnP�A��D�o߸ɷ��D�]��?WM�݌Lq��3U���h`땼��o+�	DoU��KRk�.��pg/4^v�T�I�H�ص��ͤ����s�4��Ș�3r�5RT�����Rh�m9���=]�-RI���8�8�����Q�-m��En �[͛:H�kU(�+i~s�zE�XQ��Q'u9x˥C`�X�Vk�t�F7Yg~��ԁ���=]bQ�sf]���E�i��2�i�>K����������Du�}d�'C���-�K1Z�%��4�(A���A�1��kj�M��d��'�^%�����<OGTz�]�9wAoA��d�x,�j�7�����G�2FmK.���d�lRe��������ܘ���$F��{|
Aym��4�j�E��%\��F�#I��j�l;��cF�[�_)A|F�}�-�\��)HӔ�ڈ3G����kZr�F�w����;�v�("�ܛژ{�?Z&�SZo��BP���D"G�1������>����b��	}�}<"���Yo�w�E����)['�M��/�CoKZϡj؎� @�U�����ҜE�Ol��p��M��Ƒ�k\=�����Nݔ���5���S{"��|�� ����eh�CN�;�R/'��R0#Lxu�E,fq��ʲ��blٶ�p��c��P^wD�ӟ��{�E���Tx���/�2;�D.���3����s�6�{��K�����Ԝ��v!{0u�H�ܲ���Kf�:ifpP��(*IPզ�!�b��x�cfY�����ǩ����P�"�M�l�h#����\�0���S�KF�/��嶶�-���&B@W�{O�r��#�z%tu���T'����:�{�>�*��^F��WQ켚q��vn�ZD�^7����� 4n�4dH�6�������[C)��pL�}$�|����_c���xcE���B�:p�ļH�R��H�2�k}R�$����m���R|�t%(���u��|�
IǓ����X���|�M:�q�G���$���|�O�ڽ��& �(��R����i��u�F���`~#B��b�����@�jV#�Z����aq���c�L����ioq+������?3E� 1�\�䩐<��'DC��,<�'#3S�>&e�vx2 �,��s���CQ��=�%��O"�y�p�y��7d�"�:Jĝ���m3���xu�x!�Ĵ	��I���9�؄?��#k�R����ITL��|TGKB������WWj����<Oߴ�J�
��ş7���G�M��\�q?�8��l�E��u��d�i��c��CE�A�^w�i�*j���A�V�tY:{y@��ڪA���{@�䙮�p��9�K%�Dj���%�ym׋�:�x�Ԩ � DM=�iqm���i3��S��&��?�N���̾<�"��g�A�__�j2�6s���_G��Nm#�%�i�z�V�L_�E,,����+������U'PjOIk�_8��z���V���[����s%�� Hb�v��xn��7@>����s�suD� ������H������>�K��<¶*�>~]��� �� �(�Ur>�5����&�]�@�I��>�o��⅓b�ft �i��SN���sv�y�~�E�e�y�4���R{�	u�YsZ��ż�2G�,��i��Nc�Y"����2p���Ed���`-^Do�9b�@�3�����)G�%�MZaJ=�ͭ��������C�Ԉosæ8��%���)�"N��N������4�sB�Z�Y˧��J
�5[@	���߅1��a?�0�KV�]�f�=l;B	�x������E{>�Z��
k]���-0 �PO���O�Г�:L�{���@��mh��Lc���f�l{jΠS�u�(EQQW4�@����5E��|�ȳB�M�1��,�ֵ���nG��nd�~�����2�f�$?���3w�}���2���"��Cy�����8B�l� Dl��$�g�S�'��N!��*�	��*��\u?��î���Z�37�4�ru�1c���1�HY� n�4p��ᯩ��S�'���%@�x9�E�PI�l���u�儜���kp��� m����p�8e�?���T6�05��Е\s[j������%O �F�*}�{g�d���j'$������x-����}��T��X�L����5d�r#~�I1^�W�z���NR|�@����-�O�fg�`�)���W�z<����"��T5�}�u�Ĕa��wI6b��Q��k{Y�ڄ�d�&��"�tc�9��_���-5�Ρ�{(�O�ˋ&r~�W[�s�%Py��$宾MTka�B~޾��}KX�g��]�1a�9BBʈ�"X��a���{� ��j�@o���=��"�#6�{@�?�f5�YĨ���:�#W4�*S�e�G��/l�e�Sy���w�T�F�@E��M��c�E�/���))�Ha4������"Bz�Pv�e�A��2��<ҥv���yܹ�[����p�T��WEst����Vgm����{I#� �tt�Mo�����%0�8����{�}��v��чET\���c�ք���a�-d���9*d�!�Q��=�^�ݛ�4
�Z�e�4\��30�nU��iAH��h�fJ����k���j��|w {�y����Z�@��-����#�Z��X�e�\^2�6,v�J�iu����j�h���1i���²��+θ�0�.�*���:�|?eZ��߱�����B���ω�,�M��j�����|q{UaS��9~$����yk�������<S�q�h!�5�5u�UWz�F�da��MsX�|�v�^�$�m�#��R���3?Q�9���H�eF����a�<^W8����x:�lڜ��'�[�u_;�I��섯��P�X����	;]���gn�9/�8d�J�SBx�Uzl�a>h>%�l%�	H]��JM�s_S%�LY�Yy2	]�e��>����2P��¸��5�XXJ���8�?2�h�$C+خ	;V�#��>~���-mg:V?�#�!�k�{z��Ae�h=��7�ա!���[ �:����5cl�E]�����.2��s��w"x�b��z:P[H��gN��U��D�W�EF���-���D,T�5�eN�Pc��r�<<��U ���%t�������ru�
*�o58`�1��MU ��Ǎ�6_��/�L�Ê5���ĳA�ݶ�}�HW�y5���5��<���%����|� �<��&H���hz��Q��>竳VצWO��B���� Hc&~N7!i��]L�y���<�1,�xE�\eҚ��4�q�Б����5KY�|�%S<�L&1r���hӡ3�y��-��Zg]��Zφ�ĩ�K>���p���9�*^&�b�m>Df����'�c[y��ږ�� f�
�z�ܪ��9�8cT�^�5�pzr���Y�n��f�'�T�ԅ����D)n��;�`qb4@Z"V�c"���*�F����E�� Gx3Xe��I�vYX�5"d�r̧\����;�^���8@�%�����( ��dv<��_�2�\�����L����[��	貶�|w���re�W� �*-�l�iSM���!O����<�
UKbb��Q���^c P[��d��T�C��~"�K���o�$n���1s��Oy�'%_�. ��}�4���Jܺ�9(��;]o�U������=��CkԊ�"����e��U��;��h[��ː���ѭ�ו˷��;M�����T�+�%��q�5���� ��&��c������gU�����>v�F{�NJ/���tc;��|�z�Ô����3J\����E�[F����1������w�&��~���8?��@�؄븷����j]�9���%gu����6]�ejcQ�IL����nZ�v�	��\mlÂ�r�G�𒌙U�T~���vr��丂ύ$�J	�7����>u�9�=�Ŭ���Jb��,���3��W�s�h�_e'L_�1éT��2�4/�P��M���2���5�Xl桑�}z�y�w�XP�O��j����`CԌj�