// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:25 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Txa+d8jQbo7S5TavIhWzdVCtWRQEHHZzaa389GXrOjEGV9ZiVI75eSZIE4lN6MzC
4A5adAqTXkT+EnClQHpa6A+dewTbd8x90A/327fsvzYQi3adPWiOSwKkrg0fMh3C
jssj0ZHo8msdWQHsQO9mekhoN4nhBBWoOM4ikpZH410=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5920)
pENHfLvgfh7uTUaN4aMnlIDqZySWXaYKodyrwcTbZ3I4uNPkDAwkFRq+H2txSuhC
e+OOksu5YlVzdc0+T2G+bRlxVJWQAHe6Z/1iCiHEoM25tm7gM26RnrIjmscLV3p0
MiYcfSFUY6N6v56OK5HAmacScQ1NfJpcNIgvw0uBXA7rTMfL4h6Ebzc4PUJGxx8V
IfdIf7ERBhoSWq0lC/0OiDtYGRzp0IiRRz9gxBPE/fgCQt+thiKOe09n0m9A3MWS
cVlIhMR1Dhkj7HknzfWJYi8X9rNFDoGQBCUiZGh1sHIluUU/bDmTH+qG662yFHxm
d+xAJVyVkYkad8LUL7A6Qe1neVaYSXlGCEIuZ9855yfcRklEAUuqSiytPUahnsay
hLEgTxiV0yv4l6Gff9ngRC+lsKGxX7Y1XUsR1z4+uJAc+rh7IkqzOOAQ2HulDa/6
V67mdDxA9k8TT18s69w6MzOrLt3g9FjXIH6EaCwsEmWfZbMaNLafwUPhSWmiY3/T
t6wS+ESkDpe2lenof+K37vI3pOX1mJ1tH+ykMV5VcxL9zI7eEXMD94IanbD0KbWj
OuJsKg2LS1pgGzsiMESCQUVn5PvnSj1fIg1VAw3QKP3fvVTfG5lla/EJdyTR+YUf
aH2u49dX3+7CITbtkXiOnTn18YDgOW2ClyR6FxJHCrVr+bW7XCwLXKfHVcFlB699
1fSUA6aZ2zVK8tmuLgDj/EQFTb5whokruGKNzH7TfHu25//RfGK9Uqc/cIUZoAwi
Jv6ImJ8apj/4eqVdbUjebotocwX4V06rEtnE8ABlzkQ79GTVPGQkcgmlTtsgF8Lb
FK9hyfk6SswNoRmRfkxyVbP6BTrBJY04+IUaTIM60A6lJ3SaeelE3T4b9lITw+gn
xRH8dEu/ohRNJQLsmX5QfN9jILpJIxchgHuobaziteJ1nVddnkuIN/DSQ/U431EG
KwhC98YcZS0QBX+raYKeEmqMuPtNTgKto5brZE/Ghf5PYIIyAv3yRXW/epsq/XG2
FM/R9KShAgURRgdLZOl23r9i032nkrThP5dePn40FMqr31RENexAJ5kyv24e1vDq
Al/pxtqGGbP+LGQkxFCciwpmmEXZqaCWOUM5RP49BAK+YQ2eXcKw4Rrob/Pw+c6F
ZEIliJpPUBomy0X2c+WmMGAE8LsEqLdrtiXxqSx0+qVIjpELyE4ZQRTM1WYXOsWl
60sL5q6C69YPgeNhYxNDOrgUFKnkKIMMa8mLPimgX2bvq2NElQVXWVvpebHT/EWx
nC43mPwYPWy7oxSZGHvGXRbb1ND8+fdXzQWV0pwfl6va59l0gok2v+1s7mi3rmI0
RwJA7tVez89RybKl6Nw/6Fusn8UW5GYNxSmGyMLtZL9Q3dPwTlAJ6AdrNcNwZjBw
EixWHgzKuXyoNkt3QdXygDJMDvEOD3+8UAqYe/mqLraMW1YDh559cdG6+BynuZzA
fTtB3X4WI2kMTiDrjoNhoXjdr/+oOu3GMpWQOpDgA+vAeUA7Lsvojg9qn+HAsP2g
ML/FB1Q+h4U2vyMDL750oRSC93qsqACGe2iKqjWI0Ru2QtG+v62/VAuLDKsYDWSa
V3uR3mHIMGNRGD3qsXQMgb8v1Amso6SJqwdvsSzc/LIZGRrODCB/JSV2FSpIPK6t
4UABipu/qqGqk6B5zXG+u0Mq32QFH41jLZ4hc1wPsZUKPsQOJzeIbMqK1uLclaBs
TOK00B49/GUGQkZGscoaRytr9rzYR7HYGHB93NZFWd0zRLw/jiEXEgJcUF3g+Fci
SrAwlEZEsFAGk4Mk4M6m/HE2vmczWaguoSHDtycV1Wt4Rq31Rg1BRrW8aov5806n
iMzsOb6OUSi8+09kGY8aKvX4M3b3IebruINu887w/m1NYzl4I0FMVaDvokLnMA5L
EjIpOA6fHkA7N9LadMJ7daQFD4Fh68GCkqo66H46Df27P2bzQOXDjlm9/96wTq8z
ea7jxJj8scWlB4MVQyZfNVj2fk1yjUvuyblz1SvQJVfeHoiX4mJwEsnuQca7+jYZ
hTbQnFBnfCPNKoKLxd68Hzw/P7VXVvn7W+pxS+6PQqAmDf1PR8ynKj4tqkos5kUZ
fnlnmb6LoOtpxStl0Tt0Le9LJ9TnoAfU2qCSzUIwoVOJEQ1Y6r8w+x8wBHBcUosP
vCatD9C5cfjgL1adONE2hOLnuB0U2JItcKpND4q/wILn5ie/Z+Jxc0Fh1wHZgqd3
P7mVi9Xb73AT+tCAif2Xcjf9cLX22WMB/FKDqsxKT+r1VAmRua5oBX4XJyONmXLT
a83GTSUDe0oaa9R7pIoELLsva/I1YwYUXfU9mMLDZcB7dO/lTQBJXSEJOQcoD4p+
4fkOtyP7mp/NK6u9kWZlRkwa2HJy3ORjurCwquZiA86Zt7eBXVKO8w0GNQfUQAhk
tyrFnrdirKK9ZILRNZYg8oDD7VRGeR4H7ZIojfSIfc6RAUNduEmrAYw/LWW1fE1q
sG6BWUgJtElvNjpG3BkpjhyZstcbAMkvxDi8tWVLPqIwp/qFeWzIo3mIv15MQ9/w
vSUA6Qe2TPHHkr1fGTGCj2TOICZGFt7qsE9XQGw7E7NhHnjgKdOa2QYGWm8EVCUs
I7l6XKPm5MAInq8OMyvrSu60Ml7fg661fZwaB2B2Jt7VaC/+54gyu3fdgiaBqixR
NYhNupwOQbtvJ7PO2amzewOPdADHs1m9ZSOKb5rXwi4rk/IZdUGwTH7I1cFEUVbW
pV/wIWEDUDCs3F5xquB3Y0+sGM9AfjewrE7AuMsTYgPDPmLSML+DpsjBdu69vdsB
8laEvKqg78CNuEqp1h5xorOJMaXHjL11mzwrck3sU/kutK/16QEtl1OGbHfl3EqE
pNXraIQliRz7jRN814SnLq9Qqs77bDQ+QdGd9TFtimc5VzZVqULNGrFO40lhn9iE
mpbCKeliuHT/E0ROzi2xzfAlaeKmwRXxVvWKQ4+qitSDQH1WPxgdkHPyUzN1IThG
dqlgyJgHJ3us5fMQeoRjuGBtDqUJw/qmEKYbgIOtQM/uEzj7xKugPC46FHsUuaZq
iSBT2WWqYIW0qMyM9Xz67KtwCBT5iaOUMeFIqzNp+zAptpwYWxH7ZCUWzfbQPuTJ
csV4DAUe5Cq0jvtKJbVO+3YKQv6Sn0ewcdoUyM72Wfe9PRcSMJIK8YNl1enw6QEa
iuTlwuREkaOxOma0rqTniNlTE+IBBWCC9foyCNCf2CrZmITModOSEQ4ij2iCxmrx
Yonym/hxhfnAsIz7Q942zRWWm/bdrQnYHSbc6nj+Qbor9FiOHCxfvbwSUvkvzfio
iWMQgaAUBsy+tVOAoNVgIC74FH4TBc14i1bnVeB3wLeRphJW/2rraLiDwS7qStJX
pCebIM+8N0UQSKUuXD8DpOzgHDZkjO0X2ybLtwRu/IE/0DRiJvMCycfuqgvQaqNf
sA9ADrHIst2Wp66tKy+f6D5+69nDMS5tFRKupK8jmBObv+4AqFKTOMMUcK8FkQ4T
OwORyBn/KL4kziWwZ3bp3ZQPeClydFY20LVZexJbZSzLqVS4c8Y4Ojdvh7jGNfcH
4Mya5duBlNIuOOvHgveIBwbkzZx/W+QV5ndYMkN4PVAFQPNlB9v8ILEbXGuR1I/A
46jCqjtvHfnI0soyf280anQrrOG4bZ7h6Yw0A4YVA7YmvLJKjKjX0NH1xtr2U71Y
Vn6UZLqFGYHajs+eeK/7PPQRcViFwEHtRzRwnGyQpTY1uWPz8SyuwZrZuoHJfTTS
moZjMERBauEeWVXGNhzAn9udWpv1QPPvUMqihFx2vP5FaCjQObGXP8w27xDrXQgg
qhTakFSQ22jusj0O/zI2w2gUt1G1G8IgnoI7uCBdCmvFTkKG1jaOmfiC/Xo+7ibr
6ir3e0Q/DapQNL2baNEWEg99ohbw/JufDbdMm8oewhZHzxIKq+ZIioAtO/cT9//+
EwcnORBQbfVVVYaj9nPk+xSf+bfHM2/G8XhAxrWT0/2dJPjKbKPcf4PPQQya+WQm
yBFcMoYH6Mjn89G7lZitr7c3/+dJqTQqZ0m8DCBNP3KnkiTKwKplS/7cs4M4zHGQ
z0zjc/noQe9ktYYW7+swxftMrrQvPTzL5dPBvbtlcLHa9nyuoI4XmTi9Bt/Pnqav
NUZqVEn/MDA+QzdsIaox6UP4q2u88UXY86fHWAMvl78XXn04SHQP4g6nL9I8wIMs
X8Qxe4+kJi1UCblm2oegN5sEgQiJcIss2D9F2M4erTSeBKExgAMbGbsimktJmmWw
Xqb9NqJVukkbX2s9AT9CwFN2Wt4vBd2QvuH394LJrtEtgElJChsMHi/ayVHbUBw1
mQDd5kj2W/BR+X79XuFmN3OEiBNoN/22qi+8Eoi3pok6ELCsd7yH1wslm0Jk90pi
A7wO30uBndrrXMpKYtHCBBHGevgvfCdKq6r1WSJDIDEYTI3BVzavAM/neasHEtlU
nME7472xjL2rIFa6NsYlX9CW6yb3t9SbBQTQiwdDVnaj9h/duxktS2R4/lWaSO08
44LYOwxHWsq2ENcE9vF+EWU1I/nvN8IMWqg3ys7MlCTkZA/ZsYZfPrCO3CGrlIvy
WtjCautZbVxxYuFym5TTlywEIfGXQA8WuU1zXhLOqUY4BJ6A/KrApd4nC0dYyny9
zcIGLTmZgPtYkZKscosdKpd7NJU57oLpKC5jityrrcNY/FTVFCpWFNuZzvN53Epa
nv2XCaAtKx9s5f/3+8cH4HVr4iGBiqH1l7he8Md3D/W7iAw3nxz1gE2tA0p58QTi
n9faqNsduZiO3kRX/tgt29s+qX4LawfPwHySlo69RM+2IPkD6iBvelDp1qk12pBj
ppexinQNvTSMVyHdh/CChPFCG1pb4zO9VMc6nedXGJHtkDa7dOSOjThn5PKIFAxB
Z31UeTKcJk7IBuNgiD55JD6PBOyBjskZsnS/IMPtO+iMawsskbihgfO82oSd/VgR
WY76Vqoy05e63vXJoXFhHhThgKrSnxrVTcMK6qiASbBicatGloWbasnIjpG0I+4H
6CA+8AxMJgheLWvyYFiFgkq/+90pUvs+HWAmn94WYpxX2hfUbL5U7NXvVQVAA9UM
f3q6g629F6tl/jz5ihzkDToGSHwPFAm4gN1OCqYY0Uo4fJrbRUIx/V+Hfr+urvER
z3Cn9RAzj97dPNy4WS+gGKswcz+Y+CdsUm4G3BXcWxj5MEMVAzDp6ZT2j0r5Kfk+
zzctmbwQBr2WkQKJU6ydovWX40VffsVv0EY76CHMn0wMO3/cfJutN9va+w8qaF3l
K2/s2GzQB/s3WyCCgzBtt4QBTsqPI/d/jVZ3oXBRG2i4B+a6k7NqOBIiMcqH/LY1
mugRBsNA+htlOnUhv6z/2nor+TkFkE/7oFTKjM+k1IUJTgkOv9HNSyO1IyNxVZIi
74Pg92oOGnCNxOtNBtBLfWFY/xrKiS7/aW0Wo3YdmHsZRoQa9XsSqxI3MPmO2K2G
47MIq0vMyWzPVQcKzxB1myjvqwipb8WYmgnrSTRyiny+2oea3ah7f89Pd+AI2dF0
3ufOSH1+qDVQTo1ci5YK9JNdp+IPBk7BWuo/ZW/3Syf1fISIohWwrFN5pHb9FXG1
hkD1tPXfAbR5ICewaPiO3MjsdjjyvEGS3sSU3Sk+arFvSnUh0XNDFbwbMqvOCxlB
IXtynypXcg24RYOiYD40N958O9/VG2yCdjVjJnJkFzsNkaNYyYMS2ZVL8EHnL6jB
hSiMYdJwNn0WUTFsEosZjYCV/oatOwxNWXQU6BvvpnQC3BBLUo4n8vhURNjCnDXI
M7LkiIW32PotdmzMlJH3VRN13atrOMXpu+ZwpAs7MeOnwAlkov9CjG8fi8cb3x7L
/DITlS1Da9dsrtIFTn+G0SFK7X/XMKe97OjsAC8oCp9zSrQb8duElzQYqDMyPiKU
RAxMpm4t2M86sEZGbbH6ixOcNiwb6bXxT43HetGGCht01YWdjRenVh4OaJIIC+8m
o5ZnLqF3h4y65CkbIOrbDHQSGS9ZhkWeLhZGo7rruEV//u71TUbghgl4ZgA6/n5t
UtvkF6XYT0I4JB/8L8zrP4I84m3QavOf5/nC1Dii7448IHl42EjPPqjcRxpo5cG1
Ys00oIAPR1aUnsoPjsqL5+7C6jhuyGD7p1hVC5Nx3c5NghPBLbMkZjmEAX/z3cVu
6ywFrBG0IUxXPNMgJb/Q5fGOuFo3/jc/IZOun+iEWXTwYl8OwX5ET1xqY1gIusxU
G3ivwndXjFqqYnlx/DTQZ5bJ3uCQxI2B3b7ATpNizl6tNGCx9SW+1zVQOndoo9r6
IrCiO17fBQlKJIfFxvhjvbv9dm0FAPdgIXAcuVJSKjZ1AP8XfkQPJX0KKs0GwGUV
YZ5otIpsnza4pV1MwUpgT4y6N+9JGMFGytFlQs6eZaV4TE7iEaej5a18+0pdg+ht
5RKImLzRLtn7VpbBcsPOoEq7v8uGzkEOwjhz7jdy+cwzDTaT9XXpG3PHC11KVc1r
XjKc53tfSxKNC4hCupKWRTjMwot1hHVURBwPD2T3FAmRmuqIFtNNQBgZbcp7L6aC
UQbyc+NyKH4BvA+b7bGBB28d6pOXaa8ylUSD1HbGyHD+WOvAwdBMsW3Gqa3RwWLv
YBLUVtL+JUSvICByMqT/1+zbmOukl3C814jZzpQmk3C2GEs7JxuwnMPRMd63dACb
SXjgU/TL0m8//gYFwegxzedzqnWTDopY87YRVBGYaK4kKqUt/0EkQFecCxzij6Qw
HEkKhefDPmA3xsVljjBUq/sWFuXPld5mPmXiaoErh6Mtz40IPwQ4bSQzgupQIrgz
3Pk0l7qZUaADchRf5XhOqGi0wmozKHQiID+PI/nzD10OhWEntz0W47smiqUJyZsw
AjdvmQIeGmFEW2H0FYEDk5M47gWpAVYpvLKTJ5al/eftK3Jyh4S9pAyDHXszgT+X
wmGrt2+sERBPfS+uNZ6Q5bxlhVtvON9WJ+F4R/mh0R5yszR6x4PA61yWg9HdOZFT
4UZeGi+gUajoZGMgT9yFQ1+eTrGIoJhzWT6zRnfXOnOb9lO92szofRW6oWMclPKh
rxrCHuA3fRIrIuVEAYhUpDhR9z2QTkPNs6XFvn+TCgSG8f0ItheqzaD9KOWbLxpb
dkiha/n1KWdjhOgIjVi/P81hnIGBb5y8B5MmwXOvup4JywFw2XX6hRF4+Hg4JGBg
0pRyleQVrFWTMliJYUeNnYy8r2W1rRMZ6vb5puiUw0mlfYgZNQvJBglt+uf2QHFV
nkGbvcVgRQ7fw+HQsZg1+2UWUCfHwaXnZVCRjVkOYG+jHh3RdcllyrMz0pK6FfwL
+AWYUUfFBas7hNlfXFRNhTvVIAqlBawqtAYD+uoH1WMVEbN68+DcB6EPxXsdBIIq
l9aHsaTwgrtLIAU/tzHT5Yf9UobJMd3WLTYeL9/JO3nlxZ9iOoJfLUI7Egt4o9pN
wJvgnk1+Og6nAizmNSCdUKPkfakHCzmgBV57HAJdwTQ2WUkR586Lt/DJxP9PaLrM
BnvepucqATJfpgP5YgYo1UMTvFlEPm59hpCI5/yzaJFtDPsqikLCafKiDre+pd+L
SPwCmz7goFGDT6uT7h65DhCAus4cvRf34MStYB5Mf65jnlhPJZz2Bj5uDEea4EHo
wnOHm9fVss9K0a+5K2bH5PiVJP7LT+XWj4SO5LLleowGyvBQ5RKf75V5OFD8od4v
4ANBbe/JdfgtA0hQQxSUY4Y64odxiMridOzthxFaUW7DOPsiZ9QIrtnr/WiYzhhC
FyLgNCmcctrlaxmRwdHwJAsQ7QQnlXYwmZr9xh2bfSgqYbFIKfnTSM4rBNATFlaj
a000y7ZU5+dvDvHl+NJ09Q==
`pragma protect end_protected
