��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzG&jI�#�aW������r�2"ݽ'=}WῶO��n�~&^?W�U7�>ZΛ�M,Q7"���2�!b|�Αm|5�+�
\4�al�c
/<�"Ҍ9~|�w����$��j����e��������N����(���C�����˦�<Fx�,:����)݃�^�1�?˗<x��P��Ǣj�cM��e��*ffȘ�߳��� H���5�4Oo
.�Gf)s�7��&��ˬ�%Q_"^`��'dh����F��W�Pi������m9���9���{Qbxٻ�F:}8fl��G�T��þ�c�=�`]��O܋a:��!������61�z��f��o�g���K9�cI��8�ya�]_C�����q6�#K��~;�� �N5���A��4Gʀ�����rw�1Dr�.M��n�ב�W�P��'��Z�{��|82|(�Z�Ub�$�rKL1R0��W��Y��d�^.�;W���w��I�]�mUa�(T=:!�^�ӯ��e�̣$�d���S��ϛ<Q867�b��}(�g�j�[@���g�8mF��Q��!+�K7�R[��>F�؆�(����B��[F{��3�UO�Mi�ȃX�<�7a!��v����N�V
Yw%�--��Tρ�q�r�����)��E$��7�/�����=�g�m8~�bq(L0f?�hz+b� H( Q*FS�M*�ܖ_�H/��$/���/f����G�8r�VJg29I����!F���߁^"��:A�
���H���fl�1T�a
�������Js��7A�l�+�����D��ٵ�{(��xu�%ºx��]=�}بZLsM�(�3�8�.�����NZ��0+�;4d��/a�j^���9oW �j ��E�C�Csfs��v�W�P$�8���S�CB�y�����i!5�7�Q4��3ߥ$������|�w�����jy\ѥmR$�k��
|�w{M�{��|�q �'��P;j��-�W��]z襪�&{� �Q �p-jOH+ڔ���T#�X��yp�{b�����!l���A1��m��	���~�v�/�~���iˇk���>�*��ꍞ�`�d����C?��8Xt���s6bMZ43�n}bP���~.c�^��8J������0�	�3I=4@�΃Rs%��p��]j!���I���>�֠��ɾ�+���zђj,%JI�T�Ow�U(0�g �Ԙ�!�L&��1�+�eMi��$G�g\�{��k�T����̓=ˊ)z�
d��~�z�H[{�C�-�4�e'�$�D�� y����g��y��dv$��L��B�g� 8ZF��ޘ�d�z��<%}��O ��a�x��=+Pn������"�J[�.�~CF�����2H-Ԝ��Ϣ�(C�$����:M�4V^��;��5ɋI�ñ��lօ0B#8�o%�8r����/
ed�V�e�0��G���ʅz�<(GS�[}��,:�R�vF�[�K��X�"�a*}�=���]>qd��>��RKP���v\�MXq��1
{G��cV��fb�㝻m�^���fG!"��Q�?����*v2�V%��f�Uw���
~��N"0'6Yd0H1�E��Ml����g,Z��j�t��d��
���t�r�~ZU� �K�W��r��˫�s�{��I a���'RϜX�&!���a:Q�Ґ�}8�]�]����bezzk�m��)�/�X���Ïz�<��	vC����ۂ�XA�ާ�����*�
zK�eS�n�6V��c°��4d�O�B莘^Ꚑ1��:�ΠE���������*���9��X�\��&~�Y)�2D�����:�96�T��>��oJȊ�vw:}��t�5�.�� �1�mU+>��*Y��ӓ,��F�m-�ͣ؎_�����&ن<�k��{�>W�]�u�?�,va������xn����0[��&U���5:1�u��w��Yl:��Vbcj����Y�_3-`�K�#����s,}8��9R�@��o瓂'�����が������P=|21k��=*�t{	��O�d܀�������5��N��;d���u�\�
�&th��8�s�����V��0($;�'i��$��82,�������fR�	�5."r'�l���Off2q�褣����N�-����:F�mlv����CI_�DPmy�Qz`;�i@��������R*����T0�3<i4�����<pW?&~����I>��㘲	�L$�Le�ƪ�͌-�.P�]\�����؉�+Ś~V�\��M�T�������)�*�1~�D�m2n�����9:�|� z�{U�
�Ɵ>Y�S�͓��\][Aǋw ��[	=��C��*��v�k	$�3v��L�]|C�����