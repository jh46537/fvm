��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7��z�&��`�I�X��a22}L����*��S
�8��r �n>N�ip�)'���%*�} �_쳁�3�K���è��Wq���ed�j��GB���Q�2��E�EBw�jj�S������u<]ɺ<��:�m�<��U��.�-ҝ3^���bH��
�y��0f�_>����V�F$)©�3��O|3���N�iB���L19���'���Ͼ`�g�Y�o"� ���F�y����a��<�/2���A7b�&����d.��Pe)"N��C=;�,�2"�2N@�	c�˓y�n-݄��6wٍ	�-���������������q�
d%a'>&��(	D\L-��g����+&lܮ� �A����YIȎ����d�t
w�|����Z��.ɝ#����[�G��z�I<u�F;V�0����/F���&G�y�PY�#C��FSjT���H�a�����'������3D$M����34�����
j�)]tE��Z�5 �t�f���m4܈]�vX���J��%����}փ�7�~��Z��fd��[��7J<���oo�ޟG����/��`<ª^���������%3��<#�Qޜ]"` p�N�+H�!D��Ƨr�-ϭ`��c��JG/�(i'}�%��T�����+&�B?3ɛ��\���1"��2���^G�Ʒ�� ]M�H��~�
����n������p�)@e�#_���$[��Q�_@�̪.��v��)�M�oY��WB<*оs�]çO�;���֘S~x8�r/v7@�T�U��-aVJ{-���6�_z��E��֝����F?sG�7Tg2$6���M��uJNN#��T�#��r�[߇|
9�������6 �R��Jo���/0���a�^��&>MJ�,��ᬁr��z��@_U�idcf�k:�G��d�r����7B� �#���=��=W�O-l��/ɞ�?�a�l$�L.�c`�D��O�� yB���k���?���I+�0���!{)ݹ��+��@����$r[�=��V`��]uboiyR�6<���8��͵a��zU{ 㡇�����ƒ��0�C[�8�&fn{���y��ǶI~��>S��̷������)M��Z�j�◇d1-4W1��[]F!��d�ߓ�d�MX1+qK9<衠����6�7.�&U��.:���=�E����_%�F����X�g2�(7���e�k�W]�é�~IG�W����/��ȵ�Bؐ��Y+]kE�|��=�گ������w�t��I���.Պ��N8|�`��+�ѱ�\�����xg��sE��{]�:c��A�/n#|L���G���֮���V�k�y��q���J��&n[6�P+LDr��I^Q���A2>�O��x�蟶�:.�+�/�~�lEE������Ƈf���`�8���nM�Ue��;���U8��iy}�`���VT��7�7"yEd
؝�ӽ$} ������4��ݺ�`�	T�+�o�=�fv�?�&�h�&DB����߱�����g���Q��cm�|�����b�[�
W;�Pzm�Z�t�C,1�ah�"�\���1{�����d���Q}�T�^��$����4�0TB���1sY!(λ�.3���϶�e݌�0Cn���}�������^F������'b�~/��:C�z����_C0��X;��pT��r:�~�-�`- �t_���b�ݨ] �&�k�oYv�Vx,jPfwJ%{rA����J+�?�2}o��Hl���yJ7�H�趻��rc�P6��?e"�1����u��_�^��#�j]|�-G��ɑ��>_^�9�B�3<%��NKo����B'��J�� 6N`���)2nw��T�-������;b��^&;ƻM��l7fnFl���|lH���=ڄ��_Qr���if�s�Ͳ�_��&Lm*���Xi��xTտ�s7ƙ�%�+:�_0w�ue(j̐7����Й�2LF�~��l>Zt�=^���[�k�7�s���T�j0~];m�b��}�s�]���~&Pa�V֫��=���P��=�"�:ғh�V����/۰�Mjѭග��w\j��eZ8Zb�{o�-d��*�����>��^(�G�2���" ~"w��`��,�;�yd�/뤄-����$����{��C�B�<����]��AF��DTF�����	q~K�wz�I�+���X�_�xC���(�x�#�b=���cF�W�p��<D����вw�Z΀�sn��S�e��"U���y� H,$%�G�-��߸,��]�>���Heol;�4��
�b�[G�%\?v�$��%.��t%��?KYI7es�/`C�E��4��ƻ=J�͸?�ψ	f� 0�w%���P����rv�|�F��Ŋ��¡X:,>�R�˫������x[L!�E16���3HM�\���4���v~ PR{���j�#K�-�reI6C0 »�i\�W�Xͩ�c�Gevzh0�A��kҰл��6i �𚇱��e�����FP�Y稴�%�2�����%�c�A�W��+ȵ��Y�^ƪ�����*ߏ- b�Hq7:"��U`v?���u�"��1I<J�x_�%-�u����6��s�����|� ���c��oG�z������k���4��"�!d�6D�p����e�R+��I2;j��k��`�Bg�T,%�7l3ॕ�*�())��NJԭ������1��&�����ל��EWJ<��`z�U����8jnw@G�i
�9B����ጓ���߁2�6� �.��e����ې{ƕ�ڑ2���5�����l)�}m�E��pWP���|�ܡ����sR��@�7rJ��?�t���R�rހ/���=�z^ڶ�ȒY���1	�paW�9A������S����ҝ�B�,n�����S�e��M�S~��e�v,Dr#ɜ3	��F��*�B��8�EX19K�{�$�p�>X�q�.,�|�
=��2�\���Q�ՆV:\&��f�����!ODĸ����Q����;��Ԓ�j�#rO���( ���}8H��×[u��9&}/�{�H�������y���o�����X���N��Jx�%��	-�8S�k+�H]s�)�U
�
4��9e�6RlR����ar���6ܒ gښf���#
O@�����'���W������ED�q�^w]<��B��щ<�]���r��nf,�$���|�����6���T8kC���GP�����nMC�bxvJ��c�6��ll*2��=���Ç����l�8�(2���t����a�u��X�y�^̖i� �_�}�8HJn{]��'lj`>O��tmn<lvX�;���s=\��7_石]��#
'9O<�k7(�m�\`-��"%�C��,wIk��u��-8,���5��tl�ƫ�,9Ȏ�t�M�*����Gع'� �.���&��:3ɪ&ޒ�O����j'�M�Çs���t��4�R|���	����p4l��V��5S�LŅ���!�J�,}��ƺ�8��񥗁�cZ��t;�T1T�+����:��$IA|H �l 4�C~tº7z��O7~ �i�%+�0"9�;B]	è���(�*����K8��(��'�|;gzZz����Zo��������ЯQ
�¨6�^�:�t������qe��<Us��jb�w�[���n[�1e���bd.�{Y 0\	��>�'�0�
(�?�Ǹ�f�z���X��y$A;O��&�� }Ѡ4�I ��>���W��~&��/a�"HŃkLj��)�CG?���P��.�<&��o��׺�2�}��W���Q�얫��5��n��G��˱����p�T*��k��ө@��t�'�0��"�LH��ѳ���ɃE��/=il���L�)n�g���ǃ}Y�A-�x����(y �idF���g[t,G�>C��$k��9��IZ{ΒC�=��bh����w"��9��84���<*����"�e���B'ֻ ���:H��{w��;��$<�3b����Y�N�|�M-pUi�����Fe}��F}|z�U�v�����H��H��Z�O������)��)8��+ǉX��s�Ȼ4@� <���N+�57^���aJ���#!~��
mEm\�ύ�L;�(����1A0L5���Y�|�(.
|IA��������
"S.�4U�!�Q�E�x�T�0��
�r.����W,��0K[	�vL��Y�;���	�>�PK�p��Ҝ7Y��^��&_���m�$����d�̿-�<{�N��;+D������7�"l2���s����`��Ɍ�u��o̩����Ϛ��k�P��!�S��
&�D�g!�iՔ�8�b�����ޢ��������#��i�k�&�1�.�^ard�gG-����]%J-M���9�9��t�(In��+k��=�/�y^���}[��1���t/�@�X�R�u0�y��Z�*�	��68�qF�fؐ+�Y�	޺��Z��w��"R}P�?Sɦ�������H�ZE>���V�|>����(����X��p���>P$��1�\�ef�[M;nb$BO�"���:pV��>ɟ���7��\��=.>?�"t��a�h��n�h�6UP�����?aXa�Vqj���P��DtU�i������x>b�c�FS�Um���C�R��G4��R����6!n������.ԁoW�A^��� ��
iG>͑�P����l�>F�'��d�z!
4J�QHN0�5�
����<�	nT)�v��R�y!�t@�K��>� �]蟵c�����p�2\��M��o`��ގPؐ�Ѣ������B�ãB�m��������a/~]���Q��p�-���tpO꺛5+�~�8��E9jO�� �~���3@B�4�v�ҠV�#5/���1��d�$9��j��3���U��6^����,�ǏvZ_c�(��2��HY�>��,��<��a��%1�Ў�����OL�"��䩌诃�R�����7��{�D��^ G�W�>�Fw���ZKO��U�]C3�A���)] �K�ä��.���Z�85S �rr�,�4.!�+ O�cV_�̿h;~��Ve?azP 
�C	���U�4]'�'�e����P��9�4���f�Jc-���� 8�'�R#�4�#nv>'E�o���JCi��B�z;߃�E�WbΡI"��@��'��Rc0�weQ�o����I5Ƈ~� �;���H�Ԕ|��Q�]�$����@�H�@i59�k0۹>S��s	Zw��b����y��fc��<�t��.���LU|�!Z:��ŊL�z4�rq�-�����IN�h@?*W�7A�R5�z���{���#2�����JR�I
8\�eO��=�s��yw�\B��]��S�.R��5#D��	]j�Ɂ��7I�9���p9'?�'��ҙ�A5�xnDȔ����"U��ݤF�aL+�wW�l�?�՜� ꨔ#2��H7l��FFʙ�j��U��d�h�"u����z�����k���f?�[�g6a��%!�������*�����C��>TӍuК�U/uvʳUZ�JװG�� ����:�N�/��5���jlR�