��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����i��;ݏ+��ↂ0�?�ceR
k�&��;T/�h��HKIw�|��&3.��Ů��p�!Q���i(�+��gX]����\G��/"�TDV
x; ��*���1$���'�os�G́�C2�:>�r��]�#A��]F�~?:6�,Ӱ������4;Y-�����|��U]�Ԝ���6&F,O���*Tkt�Zzڠ6]�ޢ5m�IS��Z䝤����VX��@)���t�I��Ml�k�{F^��-���2#��q릍@�BF(S��:�����jm�â.]"�	�i�,��Z��GU�՗��5�P�N���Lh�����	"���>�֞=]Kd����;�'��D�Yj���I��Kv���R�]���}
�jD�Kh-��W��M�� 	����eD��p���.��8�O���lD�Wa2]8)�b�;p![��5E���I6�����>FN�,5��y��zo�����f�_p)���P�Ey������0~$��^F<)أl�Ϥ��uvLi�9���~�B�pQ!�H�)Ie=�f�F xH�ཞ��IJ�|����Fpk��Hj�s����j����t/�)<{�&��ꭕ��ٕ;�n#,�b�&����P�nK��	^d5���/ R�"�5хS��tZm�i��k����i�я� �����Sa�����
��9�b�� E3j�0��ɩ5�<��dN�e�l�|���.���\B�1}Q�8��mco�z�F$����W\xf����`���іKk;�0�����_ςzk�OfK��-�i�����1޹ zj��/��f���z[���d=<��j
�!�]y����k�r��e|~�#����<f5��X��p$\@��U
������?6����j�Y�t[җ	�ܬ����*+>��n�.�8�gC���"�Sv ����*��ʣ�0#��sYF�Ç��`�m���ֈ�=3�kpF��䫶�G�:t�ꉄ�S���s/�ڈ���z	��Q��m[�����f��Np/�� m��a�GŊ��ޮ�����k��D5��7��J���v�3���Lʔ�AF7�WK�"�A�,����j�U*P�H��l���)�f�<�,���cz[֯� 9�/K_XRQ�"���[cֺ��~N��1x�@�z'��3F�e�:bSA�u%N{�p�۞�gف�zy��>�|�\{f�Ж�8�z]��i*���У��_DVS���ⅸ�����j��"���x�6�]0*��B_et
q�z���3� ���PdB�n)/���>�)O]�}��^��P�ެ�%^B���.��-j������.1�Ð[�׳EP�<�dŉ�f���ެ�r����Z�p.�V{�ݙF�_��{u�G0B���Ҹ����
��W
 ~��%i���1��n�=u�A\}p��[ �s��U��u����l���3��2��Ŭ��uU�oY<�=P�Ʉ��Q�Jg��t�t�r&�S�4%�H��6�b��)A0_��D<\f��W���dY##[�#��<NQ�#�������zpa�&W~}���_�SW2t�?�d��dO�g{�������\�PC��b;���\٬��4ìn'�̇./��S��:t�oQ��}��;Zw��af�b����OR{h͐���l��0'X��dU��V\��2�b2�y�Z��Zn�7����6˵��J���(j���s/.��D��x:&C�0p1���p�Vg%O�Bx�k�|��ھ<P�E�_$�5E�'8^R:hnxQ�{�4Ճ��8�y��w�^hWRH6X�D�y���xMI^����m=I����,�n�a��y����G|C!�ʋZB%Y_��f=u�׍����~���#����P�}�� �� ]j���j����WA+'�g�8XӃ�"8[�����u��8Y�;���>�Fi�!+��#?���7���� 6�+���sL{P�N��ޫ��͙�W��۹�W���G�K�>��v��-Ƹe�Tu���F� �Oʞ��T�����9�i��@��>���F�a��+k����9^��Ł��z�l(�X���r�����NZs�?��;��7�bX�/#��g+8���'3�c��Y�x�+���L���w�ߣ��\"d��]bZ�Z��S��E��n� �뱖������
�>��^
��w���\��U�RK��"��x%��k���C,�u`�j��.A�`��\C�:����$g7��h@6 Վ�V���������B��B���R�����r���t\�F���R�eAʲ���dq�� ��f�f��|��]x�ɉ���� ��aB���έtN��M��C��<R�]��Yx��y�GU�yV�jN�j콩p����=��H��@��<�.����>v
Ǚ�	>��P̿ŵ[m%��n��b�F��*<&�8�>K
�O�O�2��ȓ>\u���������z�Rb�޷�������G�'�;o���lR�#�9}�����~J�NI��̥9��!
�N� ���+��g�đ�F�U���_*TA�F�������MD=��J�?�|sf�q{�k��A{2|:����Ё���ڧ,خ�=UjW�+�k���S	���\� ۦ5��n�N*b���2�e|��ݘ�ZWF���fh-�XTB�B���L����P~]�]Ĺ߶����m��>�ŀ�N���>�Z�d
��*��W��J4��sb~-<v�ʄ�#H�n2Bcu}` �_�PW	��T5|~���|p+畉j8�iA�@,u��#D<XC��1L0N_ߏ�G��KIKlϣ�D�B%���!ΨtH�v=v�C��R���	��;u��E�qkO�2;�t��\b6`��qaA�o<�0�3gP�M�h��J㰏�rGٕY��N0�n �9�P����h�.���A�ql�B��%뾗�ygM�2!z���WI�s��|��a��,�tbC�k`X�S�`ߕ��@�Ni��b�Ƣ1q�舀����1��G�q;N���9�hQ6��/pۓ�7i�{%+0����2f8�d����p���t��+,8�v�����;���a|^?���b.��.W��%9��d��[��:ɮ9C�d;�P����3B��Ru'R��%�5H�ޤM��^�ӌ�*Q	{&y��x�)��r<��D�fq�]��lk���.�ۯL���Q���u� ���G���^�]�ۅ�(I��H^�3��L�hʶx=�G\i���@�� �wͪa���/Ml;.��CA��H�J�d앻����v��w�s����`���4_ء#�J�i�:�����	vv^���+7� �e��e�dP��ߨ��%V@yZ��ѩ��l��U=Ë��C'V-C�m.�{�����ýPaZ ��ۯ��w��$�*�M��xE�M&x���@e�R�6+���	N���K����X�B���[�Ѐ-!���b\�q����f���f�hq�5�f��g��%�Q�������s�����s[,I�+g�i�1
SdO�}�à!Ue܉�U�ľ�;�� ,���9����k
"��z7Q�] ���B��6ƅ��uf_�̌�A'��8��
�fcTy��%&�K��ht�Xv�:���~����>)�8F�P�.}fl4����������V ��l��u�B{;k8��fͮ�����ѵ[�Pe�x)C^��G����8�[e�	gNC�����7��c������ >_�����Ɲx������{w<�΁t#;�~�ªu1���5&�~.md�qbX�~�N�8/�Jr���HDQ_;�5o��7H%p�a��J*<�y$+��`�x�
�Nc꺸��uC�&���D������A	�t�q�n]�x��<�#�vr��u�O�5� ���xu���)C	O;�tD���g�x�ᲥL��>�C%U�-����^cCk�<<���o�{�pƒ�:h(�;��;C���B�)�-�[F��a��
�R��#a��^���C���`��KOU�0��m=Y�C���f���h�j�ei�
ap�bs�=R� ��q%N?$LH�@k�����[C�2�MW"SiL��k<�O�.������3�߈<���_���[p�,^%�в�eb:qB��.N�8q��Wn�1ê�:I5���V����6X!�RK��baYEHH7yaTc�:I�Hr�	�{�҄ȓ��Dyw�KM	����a"K�oT���5;/Д�?�.�b�.��S�g�hd�s16�d?(N��N�B��j7[�u���V0·�Ff��r�Ŋ�a��-��5f�l�ܪi�GM�����|�;��m���	 �-��m��p���ɖ�y�>��o)xR�i��ؚ��)�Ufu�a�{Խ�l��	BL�������C�����6���R��[(��Oe*6�v&��b8��3Jɖ׵��g�� ����ϧ�*Ht�O�z=:��b�[4�f�Ƒ����z6IN;��`����̉�d��-�d���2P��~�^�QE|WȨ��X��k�#�]cT0�@�}r	H���AP���3(��"��!�GrD5��k3�*nMa����.�$�b�󨩪�]ĺ���H|kj��T��hX��d~�ϸ�{4�I��Ӣt	F_�i���7Y�����&�o�#@cM���?��,��*�l��ޱ�ư$�^\�O�M[\0{��g���>M����o��ec����TԦ	a��v�so�E��}֚�%���v"��D���1I��*$���l��_����,�'B�'�� V�'�}܇C�V1��`�>�2L�G�4����{���^M��DߧD%Q��NZU���&�n�0��{2�!l�=qN!O������OAH=碲C�uz#h��=3�M�j� Ve���*.~�Y���.e��;��c��7���ҩ��{h�{^G�I4`��.{{#^�Â��+�������C����?Y��K߾j��q%�h���u��S��7��ᦂ�I�gC��+HD>�Ph�]�K5Ix|�4��{8�L�d�`�V-\��"�.�o����ʕ������Ֆr7�C�4g��^��E������EP�p3�#��1�*Fش��3����F�᫺��FO
�� E��50�|�#���~��1 /��>��L���vʘ�����Ψ�kt^^s�6�!|��5����������c�e�C b|�a��k$�����K�%x���sV�)�� ��z=7��� Te�`n�7�gCHe'�Lx���!@'�������u�O�u>lP���l>,��=ge?��~�6���@�!�7�--֛o���~+� �o� �5�P�]�=9%�B �k'|�����J��Q�~���g�ܟ/5e֑��=��x�6��چ�@��ΣӃ�#QX�A
���,dފ�[ݿmj4����˟�zԎ�|/�B��]����n�mi[�ar�B��DH�0�����)H�2em��V�$�H��������>�T�A�N)Wl�W���,��:S�G��B>������A�M��ff �f��d�i�"�9�'8�+���J�CNۑ���Vsv�Wc ���;��{X���/9�o�QO��7K�Äju꩏1u���V��}w,�M;ɚ���]hY>Ժ��I`�M���s�[(~��c颳����~j*B���;Ӭ)�aH)�<'��?���e�
̡JiN�����`��pd�ys�&3�M�[��P�P�����4w����	����*�xk'���S�)H�+��e^+-oQW���1��>�ͽfCi�u�!� ��_$n��N6睦QS>��$�/@g��pj�X����WҖJ������X�X7ǔ��_^�"��>�0�������%{}���{��pk���W)���R�_|���^�B�]������p��?�"�N}X).8�t�."U�~qj��|*��ڰ�1 &���tW4]�cx��'^���s�U�<�a��T�]�|Z)G��T�B��rd���-�'}�EF�Sl�n-�7��B����6���_�dZ�R�q�w��U:�ĩbz�"�`�
�g����'���moe�Ԉ�8�2��݁` 
�*�5'��v<�z� �p��ղG�����9�4s���U_������x�ӱ��g��^o�V��bFvL:��a�.��2�����O�cA�wGD�����Q�VȔS_�ݡH�#6S�5��ө,xw�Ga$<+r騡O��M��jH�!��6 Q��ͅI��3�C��S�'���_쥸�[ ˥}�=�DuF�xS�nzJ:��u,�JW�Ih�A��]�PaG�ĠOb�I��P����e)�=9q��2�9�
s��z�;�!�{C���tR���7���7Pi�YK��5�G� ��[�>[��ڭ��u[���T��rõBͪ}��)舨�%��zl"Nb�����؆s6|9��'X\zlmmV�q9�S%�0���	�P6E]��D��ꮻ���u��K�ԨVmQiؚ7��/@L��� �si]܅ە�	�%��z`dW���(kd�$�w��j���m�`�}��i�Yg�Yy��n^�@�G��b�����䟺72ذ���V���~�"�c�𥵘:�8=�^��+[.Vg��*��ɪڭ��i
~��j���v)X�q�ʫZd��پ���r��w��◴ܭW
� �{�7���&0�w#���$$"�w2%0�iy�|.c^��'�e�ШY����
�:@;���1w�>���@�D�@k5���R��>ȑ���U�z�D�u���B�q3�C�*�0�c-��X���u\Ssϓf��PYٻ|�a�jL9㾂�Bnc���y3�!�
,>K�.^U�X���"7��(W�� �g��%_LK\8n���o8��C�ѩb������̴rl?� ��_���5#���g�zf�Y*�TG�����sp���G��0K��f�hg���I��*�<)�M<$�.���E�[
G �p��bP���oS�*�L��*�@�XP���3+�F�/U���:"Dcta��!�E�O\�%���&�"ᾒ��<��^��Z>�pha� fe��W�L����a��/o��D��d���,CTTnL�+����A1C��,�Y�eq�(��!��E�67���Q4|'�8h��k�ɔ����������ߢ͊��g+�nEY,IK���uj���ֶ�E�ܩ.�j�AQUz� �j� 2_���	�2s�S�1�4���;?[`���J�=UuZ9�֭[H��`u�l!݂t�+G�b$�lB@nD�Vh�M���O�4��,���v#�X�r��.������by. �lY��u(�.�XYE'n���/r�/�yX��X�+�DgO@�!o�A���D����9�>r�Y`��;��\r\A�h5���c�x�"���/�r�9�2�^f��7d���)]����� 2di�e8^�t�t�y�|*U�U�����>�*�Ϝ��;�sȑ|������p1)�l�e��=ɮk�����[���i� ��g����m�.Y��%|�[���n�!�w�A2��S�k���6����U-�P�gj`�ٓ��A��Wgr7�@�O������Ee�٣��gP��w�a�[�r!�>���o"�$a��	������iN���� W$�a��8q��WcS�U�*V��}�Nz���1��,��]d�u�P�/���;��%�5We�qi��VEυ�蕁=]����t�D�}����%�@j�Y�!&�]�ݙ&���q�[`)GpH�0[ite��d�Z�9��n2Bc�,����6g�`+�d�NV�6< �dٍ�C/0`��h�!��M��������>�b�mx�LPՎ�N�2�9��*C�XF�[��$}#�5�&�������Mc��L�M���
�WT�L�"�F���#oFȔV����ע�M+���TE-�;|��Z�l#��|��5����=B���;���ì�+� +z6 ^\-����O7���Rm �rVO��F>}�	Іv�r@���٨�c�-Kˏ[�R����''C�s���F&�s�=���;�N7-0i�"s#�7+�e�&��dk��<Q���(DP��G��T�h�	|.�V��ݛ{�ݗ�T3�W��C�W�6L�6䵲=��m�3y 3�ǲ��|˼ ��j@�h*t?=M�A���.�����
@�5I^��2<��ؔoKhؾ�_��Z*�±ƞ�#OV}=�3L��c#�
���+�"�<���8�*3}�RVkqD��Q�c���jB�c�#_D�"&�a�����5��>��#�;:nEl�e[�Y#�!Sj�u��r�0��Z2�֙���%si����ܿ��h?�!ѣd�E���T�͂f�]H%^(�Q��_BME6��df�>5xUCM3B%�2��:cF�����)zL�f�F�̹�A�n���+���������$�fs���w^��-��z�n�=�$��U&׆>�TV�9�`B�9��\���riؕ�RM����w�Z��Ϙjک]{1�s�\x�}��_vݾ�VUCRðٞw�hW�j��I�v�"�<xd��9�W�0%�:��~R�@M�9�:c�n�L�"���&�S�� %WqȂ�7���^g��0_�_���ɴ�oI�<Z��A�b˓��1($�����ŷ���0��P]���N���ͳ�	E~�9�ͻ�)Ap��:2�O��P>��a�mM��Q(^'��#r(�%���U�h-02?�c��@�QHBJ(������şd=�q�5����uH�I#K �;�3�
�}%���,���iFm&�~쪄����E�h �6���R�S-Jz���^��VTw�[4h�r�|�,K�ڄ���@m"�!��A�L����VӠ����I��\b���Ԍ�������y�F�^E��WMD?�@��	���%܏9F֮e��JM+�lE��؅�ӛ0�u%�����3ܱK���GDG33�	���UN48��ϙJ�Q1w���T.�km }_T-�����&Q��g���L�`�tG`k�0��t��M�����΃ƣ�!�#�|a�5���nݭ�(�8���MG��>�a$��~f�a�},Qc���{{�3�b�f����%amE]��x��V���}�Y؛��,���Uf���F.�����v.=��U9��M	E<�k��j	������d�|Ϗ_�d6���?�L��7���^@.>l� =f��ԏ���_	u��ܷB�����K����o3Yqbwmr�9�/1�?:�q��$Yg'���~5�[.�c˙L	�an NUЙ�z��xs�%I�C�l��6Ր�{�ڙ�͸����N�>#�mD��m�%л��q֋����h����'�n쳕��e���������	��z@h�X(������nJ��p���LO���k�L�})7���=[JM���/�L��ƃ�#��8���?^��#���0�ZC�~ljP����q3�	����<?��㓖�k2�6��Xz�'�wS>��fS����ْR���L�	a�a�V��e��ￔ<'�hhc0u8��Z�W)�Z����J��q�ѽ�h�i?m%�d��#[�(���Ɖ��16*L�F�S����"3�H��z׊Lόx!���ݴ��F�go�Ȅ�P����tALn���"�IW.j�ZެR+�������-�*�9�R
Al�/�X��w/tѮI$6t^;�u�Ց<;#��(���l��VA�44����� t�߈���f��S�%i�T(�x&����ϲ.�=�:�44pk��O?'����}{�!�*�:
���=����MU,Cu�
��9�̝It�+tQ��*�U�i�� �RBZ�(�byy��������)�4-8 �a�IN�~{���X�>W�q ҹ�`E*Q���O����G=��m�Wf�t��k�Y���g��ED�~���9�agB�M/V4�մ��6!��ᮜs��L��`�0!��"��Ցq�L����ğ(ڀO�x!=�C�L/@Y%4�nx#�}_=u �s��c;��Qw�I�$U���i���#�1�GQ`E�j��ǻ@5p�)�:L��7��[�}���q�b�����w�\���[=�*�M�Bâ��ڧ�d
α��>Ý�����%�=7�b\4�E��}N�Ž���:����HC����h
6R����*�AJ�ŏ^}R
$l9���X��c��vS���~�ƙ ���ncK{�p�߀��yb[H��zˉ�F�a<��fGAm ���v�U�[k��)y?�����mzΓ�a�<�x�f��sO�je��&�1L�f�'�.�����]�ױ&Wxi����*$f:ɐ���'FU��J�*���f�7ix��^���1��\��x)���J3���&Y��F�9{B�(o����-`��X�n���k�u�L��7a��sG�r�X�P� 6h�~Ú�lI\�2�H^��md���G��	���LLC�`�nn�%�!ը��S��,t�w�Q�q�7^*t�4+�l���M?��ڶʬ��5~Y�/����L�����������@��:���XB:�]���!:6.��|�[���(�񌒹"%!�"�Ӊw���N�'�)sbΆR���N�'�P\H�p�N|��UU]ˣ�.+ڂS�Zn���D�4�#�᭶t�'#<��b����_գy@��E5(SP&�*{�pA�s�5f� ;_���kA��D,�dߓX��B5S�*�iUv�Z;k��w,�e�'��_��>�� ɒ^j�k-�V�@$�� �����}�)Z�<Z�H�o��fSTr��ǘt��%}�۽D����g݊�t����O��Ok�pU�ԭ�c�c�^a)zʎ�F��3 � r����KW��=�Dd���W� ��S�y9�m��y��I��� ��tO�L+?��C�p"�\����xt-�%�C�=�G�*Yr�4TH2�7m���$���_D睺��&�l2]�ߝ<<6���6���X�,�r�mM��R=+�K\�PFT��\i�9�]bi��"L�����
2���X,��h~A'��8�.71��x�m���9�2��J�2b�4���޽J7>���z�y�g��jn�g+�Scw$��pUb[+]<��_�V<��1{�:�1���Yߦ�£�h��ZH$)^B�xH���[�"\� s^§y��M<��)�-��1�ڮ��L������Մ^&��to��
�XT3�=��Tm����u�y�쓝��!ش�q<�,-�+�Ψ��^T�]q3�U^�xɋ7m���jK��H�n�*�6�ʟh�"���'sb��4U�p��յ$t�Ҫ�[oP*]tn}�$W�6�.�r���\GS�������^��v�&�Y����R���lUXA��׶�$K�ģ�8mk�ո����_�u�U̹_� ɖx��#eغ^��|7f����y/��h�&S�M��?GW2�o'�h,�3%v�Õ"t|�?@<`��Jd"����,)�U2e	�|��ˎ~h���Z�B�G����
�QJ0-rn��_�?��j�=-ò��/��4�����8�;�o�Lg��ߋ����Q�*zӫ"�K�M�J[d��wf|z�W����CE�cD��|i���J\AZ�-
�qީn���E�/;�p>�CC'��/���to��>��_����h��7C���s"�)\7Oܶ"~�y(ƊŭY�2�Q��\E���Y����"x�e�9�ژ��dƏ��%���N��M^"S��U<8�}������3�3��C�W9�a��<<� ��(;e�w�"3��P~�vNz<����%�ʟ���7��F���Yz �`�|����"{x��	@��>����_ጯ!��s�DV����(��K�6
���H���mC���������S�����{�i8,�4{���IJ} �	�;;P���e�.����̓%[���(l�޼p���Rh�����ejq��h����}!��X��z���&��10�߹ :��0G����n��vd\�򺥴Ӯ��;3r��%��/
��GW�j�h;�TZ������?b���]�R&�ּ��B@�k5������U� [cJ�/��O����Py\����g�BD�������iLph��e�����s= �����^�0�<��4}���x�r�4T�b�����E���E��O�_���S4�_�_	`�Xm�F�b��?w���a�+��+��\�Xb�Rq?���'O�z�=ǂ�H2m�����2�q"�j	2�v�3_�$eq�<ָ�Y�G� ���%p�NS��sF�x�H�z\G��ω��<���#�,װ�=�vBT<�l����
��Aa��3�i�twL�-Ĭ�\����Ï}�Z����Ğ��9�p�R�����u<��6��E����2���xoP@�[�徴��U�U���/�b~�WD:�e��e�(D�s��z@\�݌���aY�v]$��B�g2 ���F2��iY�iک?,4����͐HU	6� ���Ɨ���Q���F7����18Ђ�"��E�?'�~N��rs�3*4���-���?�S +#�q�����H��A��Y	�C����$�򚟧�<��YP2%�h.�i��p��R'��䖔��t\�~�K�O'b��s��Ǟ�t����K�޵�S��@xa7ʆ@�W�U��=;Ax|�?O[�c���.-RvF��_BSV/[/%���"JyzKx���i}7�@^ǿC��-�I���lS^y�:�e��	I�9��9�Y�Ѳy�wS�7_v��r��[7���v�(�r�7L���^����7��H�f�k�	�%�!���9�
5�_�L�V"đA�J�]����g&��~?J�����AuX,����. JR-O���bi�*f[gѮ��0�y�������df�Щ��7ٖ%�^oA?�QڳՎ�F�����������emG#��%�u3"^n������ �l�'P�mLs�$EکaT�c���%�A��1�O��a��*M��h�W�B��Y��\��_���uh��\�:��YDzC��ٺP��[�▚"g������lH6�9�06aE]�+���НА��>��C'A;�U�/�p Ǚ��K�tWoN��@n<���;D������#�H�=y�%�߇Є���;7�1P��	�`�c��^s��u��w�g�o%�fn3�00���Z��O���3�<�L{�c��<��{���)�2H�}G���~1=Un���+��W��%S1&�K@��&�������7�6��hk�H��)
{V�)��1�i��Y~Ce"j�� K�SJ\+�v�G�P�2S�]�%�l�������P{�6j�h��#���A�lx�+�)i+(�
fr��Ds��=��j��,~.��$���1��� 5b��D  Ǳ�~�}{A`�-ȱ�G�#���0.ݯ�H�Pu��>�Ul��&������Ig�I�[~He�c��x�5O�6�&����Y`~�'}:�.N)�����W�Mq%��Ud��0!lJ����t�&���ӛ��n/.18�>x���ѼåCގ�̷��|�<����V��ߊF~I?�1��-k��m	�o��I�W$����f=rRyx���\k�:���D�`hPR3�Ob;ݱ����-y/�KHٗ����3
q�ǡ������A����[	X�rw�]���v���h����,�-����r)uVȶ*�B�!Z�8�XB`ܪ��$za�c	��Vf�Z��փ��[���$�����E`�T����Ed�\Ow'J&l�,Eq�=\�x�ಧ)���=k>��I_"N?cGB��	;���5�%�u�_R �a۳�6����ނv Ld��6�̔<V�4�Y^�D�6���@^^y;���nM1`:����wVui�I�#����}]�'�N��0� G��v��{1vb�8E�>֖,*lI���w�#��F�C���~�jb4�y�����*�� �j9���ٲƧ�����{�I�պ/�2��l�|������kp�Ūu@ܸI���f���k[�x���R�Nw�)|�1.�+�0.����g=h���X�+(��a�a��9k���r���Z� �Z�~H=�F�L�8%�]}�:�,n	�S�I�@�{�U����^������;5�K_,�N /��5^���\��$+;��q�G�R��*�L�uT3IR))��V.D�� ���#5�/�z�s����<2D)Na�A:�B�&m�*�]1J���&�b/�fX����-�Z����m��?��
��p*,�'�<^��,{Ȋ�5@ۍ�_�P �/�C@GW4&����~�锣�x7�5h�`�ĢDzte�?Q���A+�"�y�� 3GzO�*E�2칽��`��+�>Ҫ,MUIت^�
���\:F(.iJ}����d�U�&T��v���_x�1�e�a�4�.a�V�W�/���9ÈQ?n
w�}& �_�i/����3�����Ll�����e� ���F��
�!zf�P! �a�<�؈�=/-r�{`������@��#��Ȱ*>��Nj*�>1(��WD����	�G�K��V�xmT�D<�uC0�t���������J���EaE�'Ϩ�bX�D��<Q�ߒy���>�{���ڽY�+���;�7��u֥Mhk.�b��%=���Q5�	z�yX�������:��7T|Lz�!�3���j ���(��f�f8���T��V $9��^�F%�3usৄ���U����X�Sì�2.;�4"\���B��w�O?�G�6���)���T�?!�?Ν!r}M'6�-�+:T��C��b�|Y��%�@�l�|�qg�����Pc�(y΢�h�X=�O1t��;����6l0Gz�xm���&����k6\����A^���V��)�b&=Μ�)Iw�bu605�^ݮ��w=�V�5IO�����~�j�X<%��)�	!�.8`F�ǋ����?m6������fr�U�����wq��W�g�I�3���ҋn��4�B�,���177g�t��Q/��K�)�`�wMӅ0�\�:��G�)4�R�ߒ�|Q���u���h�)�=j�E��Ȗ�3�Խ���6&��BQ ��s`[�3�|ݳ���G���m�:M�hp���ʧMé�ՂI���������О�-�|��J�X��N#���C9U�a/\�@y�~���?kj�L��/�?��
>�v&+R�6�ߡ�q��ӕ,��9c.�|���}w@�@S��J�j��V�����$�澰N������*{�?!����k^���w�[�����w<b�m�B#8BM[�����&#Kj!Ø���:�<=.�{�`�d,���-���lxd���r�цVY�%��-;��e�����s!��uH����?��~!��[���N�v1�G�uH��l�_�,/;*Y��<zJm���i:xc�ֱ(MnkH�wJ�$UC%��]6:�ڰ��Eg�|��O��"9{�(ٽ?��]�#��H���@+O�%_Jk�<�t�i0����8U��΢���rt������Z�AH'�@�DF�5���Q���23鰶e��[���� 	쮅�m�+�&���T�~�c�jȄ�����N �e�1���Fd���[|���l��b����.m+��mr%�E<���h�[�����xp뢌�3����o��-SU����E���O=���
gzoR���,����Z)0�W�I��2��Ŧ�vh� ���U?W ��t�
6ԯC����7��_.�'�BԔ��Q�w�/NJ�d���M�i�l�# �i��F�2*n�>I\}�1}P�=�A͊Ð6�Σ}p�#޲�)�/�;�]V$H�������*�[ވ��D*U8&<9��{�Ԯ	������QT< \d}P�.�U�\g2��x �ؒ撖	��BgLO��M��U��D�I���7���
�}�d�D�-���	�S�Gavi=i���e"�O���jf�a���Z}CN�O^�U\O����+�o%���k���$-]��M���%C�,cي#�d�đ	�iH�ɒ��/%@��E���,wPB� �Y��+���y]�޹���=ەb��� ?I�8���L�������Z���H�W���Ů�jA���ƅ��C��V�$�)�l����Oe��-�>���,�Y����(����=v�Rx0G�(�ɜc��R�I�3�$���G��ͱMS/��N၅�����?A�r	���q��~����_����)�aí�k�>� �x=��q�{^��p�?Ш���1�y�\��A�Ř9
���fݚ��hX�T�66.Q����{O��y�w�RAv�!����eӕ��kC+���Z*y	��d�:�z �y츷o�#D�Zwj;���$� ua�^jn�c�n���N\x�?��hX=�%��n�ބ�K���-�-a�W�6�����'���@BӝkU��+/C���z^�$/k��;�ۂⶪC�ǆE��c�dz�&*C�-��X���rCyG�R%�~����2^��k_r�~�-�"rQ�	/%4@F�6׬�΅�|�?,�P�$���G��~�߳��_�B��7�H�Qsn$w��6�4�ꤼ�u�����H􎛧�����ߓ`���	��T`�,%O	e��\O�g��^��)Qf!A�7s@o���Y��*��]��I6�g3Gs|(����ٴ��S�$ME6�O� ���/1��fD��#)��mg¿��ޙIa��oS��i^���@d�yUF,��ެ�]�ʒɹ����b,��Hkb��˞p!\����8j�m۱D�M;d���4��͏��I��NXRrj@��x$P��5��>��y�|O�f��f��2�MZ���/��m�,l]k��.V|kz��27_���Uo:�ࡵ̳��T�&���q�f�����5A����K��a��
��V�a�O<O�)ܑ�����&�irx�����N�#���5>y ���G9d�h�I�]�g�G"B��g��i�gw�����XJԚ�,����_�%H�·2��*Ni�v�'�Q��J+���D�h;t�bU�$�ag�ў�+���E��)~L1���E��H�H�"������	3�b+��x���L�#�"�k����!x{�by������l]���G���"��r��`�?܄;m;.f^k@ȴ��ɪ}w��ʅ�Vk��ϳ��Ȧ���B7�<��Ac�F�h����RO��x���]Ց�#�p��q�H�4�5� ����S��W����ģd�se8�6�x���n.:9bb���遂�� K����<=����*�01�~ۉ�&� �V|�z��5��.:V<tG9�3��2��a6p�|Ĳ,�8(��nj�ir��Y��پ-J�$�L��yFPG��>|�A��=�N7j���oU9�n�J����,r|E�/&+��0��bG��{L<�?��fص�z�VI�蕧C�H3���<fw��Ѓ"ʔf2矝ZC�����R Q'��8֠���ў�d��=HK��������]I�.�����S^��d[8�"�6����8���8OR\HbTZ#�c��3����^b2�㊺'������wwmBf��e���hexnG��G5�@ 7��o����zZ(�P�]1`K�n"+Q�'$��a�`YMe�SY�D�n����'R�$j�rY�.�ު�JM�s�jP��	O�62�B��)�M*%)�p/L������4��$�xU��-����&{Hz�>9��C�( �+�� .��b"&-��)����ܾ6��ZM�TO���^�Z��YH�)��� ���qMh\�<��v���u
��5�����gr%��4gސ����D����i�!���I��h��NP���:Ŏ�rAxX�U�0�f�?����@�	���(�>0hVy�*�D~�"��j
ZngA~�-���7�vTLE�mL�Ѽ$G!�N�����<	�Bj$or2ذy����X��Vt�FH��'�dh�2�z����}��3���0�u
pǲFo>����_jhu(����0~�E�KQL�`7V���c��!R�( ���U��.�D��J5�'ek�yE(Vpg�m���d�	���X���Ǽ���|�`�����ʴ��D�@����
�Zz����Mt�_4����X�5*�N6�T�����T k�3�t��z��iP�2;H�N7�#���s��Uk� �[HE.8F��DV�m���J��8y7�.lF!���T7$��.�1o��A1�'J�I��8��j\ZB�ɚ��-�uGzf�B ���y�Ai�
I��1̅��~]G̊B�� o����4l�V�
�,��>�
ҒԔt�8�K�X��U�ٴ���Ȓ �'���szk�t;A�D���ӣ��Ґ����oƙu�n�� ��WC�;ΎH4��F�./�C�捡����:���zK���4Do����բBK��+ܷ��8��! �@���E��&}2E}�zP����t�gԬ��E��_�����RQ)�`��1U	�5\�H��p R�
�Y�Uh�n*�����y ��23�G�"� �-{��v1r!�J���z�4:�/CT��P����*+7���@5��aX�YV��կ2mo���2�C<�d��ls��1�
��%B��(�w��R�H�7�Z���@C���w�;S$Es��n��r\�C-$��U���eҩ~da:
-�D?u�:����.�5`�I�S�x;�v<�	��_�	W]X��mYez���
�A��/��H�N�L5a�+m���Oس�8�B�������f�ـ��T�����.����x%��|N�	#H�T��]�uB��T���)����-�Ƹ/���|/������-&�L�:p=_��%��q�_T��c ]�Ō�&p�fD���#p��ޘz���L��
��]��	��z ��E�Z�9�ޝ'�R��Q!�f����4Uv����U�8�|IUF�^��O=�GΡ�KW�
���MD��V-����k��(�
�@��+�x��T+�%����3:n�f�Ғ`樄J��ϻ�N�1M`��Y$�YTAp��7Iҥ8���5J��m'y豖��lC�e�ւ�P�r^���p�f�7����2���X0g�.];{Ҩ�8O�����/v�]��j)deP�ѓ�ٮ��90,��}��,����%��*�ƙ�!YLr�zr�����<�c���j?T{k,V�YW�����VT_5)���>�������](ڦ�}N�Pl�NTX�����A�GgT�:�V��]���U>}~�~@+B�CT��z4�ٝ���>���94~ `�����1�t��ƚ(�e����f
׿�I]����.9��_������9<��8ݰ &`��{�fy�8������7����s..��{��G�RO�#~��݇���*�y*�9D��db��6d l�p=L�&�b����H;��
W]������*򗵜�&��3��.83?iu��O��C�TF�#��7 �����ֈ@���h��a.�e!M�*ִq����/]gO�J�̫�f8��O�*�55|��	��>�rV��,7�=toEs3̮���8@+B��9!��3埽m��ÿxc��&/�^�	��j��b[��-�&�p�1�s�f��>�q�C�ݮnmc;�뭷8���8< �������Et�l���:\zS|�XdRjJ:�-�5�ٓr�i:�_�=5F��]��J����Ԟr�h��� �^6P�t�`٬�I�Bdl��(şǘ����&]�[����G��I�8�c՟�^���y]�E!��M]�z��`W�6��G1��
��؄������K��6U|��R� i�A�(�AU��l]00S��w�T��%�y�I7�=$8�:�Q#^�3_`j��_#�#�7�qثFc�vI����5��d�!������z����kk�Q\t?�R�_�$�Ǌ�kb#��c-�)�$O/^
��=ͺv��,�6�F�d�7n�R�	��b"�>8�(��&�g���\\��sKO��>��K��ƍ^@X��ɻ�8M��nV~.���п��J�צt�C+����6'o�������K8�����b�����[�}���Ffa8�r;�WTu]��F�I$ ��>�$i�;�.7���>���ߟ?�Lk���tp�tc������P���9	ˮh��u��r��N'T���������G�.#4��&tT�ڀF-{{�-tT\_4�����{=�E�����u��a^���c߯o&{)�w���Da��F)�R�*��.��?��s��tTWW5��j�ݹۛ�I�2s� ��4�?�yQ�ʾ%e�oB���
�V���w�A8�%i�L�)����[Zt������J�������Y�W���G2ݣ�я�q�ERA��,�d�7�U��.-μX%�����Sl����[_mEɩV�m]������y�	�+CCΫ�£a=K�B�Q�L�#�0��U��e��<Bw��P���6��B����q��wd@�*[1��-�J�����P-�b����� �`���e�lc�+kkY3X�0��3��c_���TQ+�
�?_���~�=}Q�jD�\3J9��c�0	���2�.��')4��>��4��c��*�O�[S]���<�T�AF�/�&�4�;�k�W�F��v�9�
݄�$xdܻ�i�]M�z�lt_b��R�aIgr��tp�N$��[2ܽ��o�6�@:��ô�[����]�q��;����%�t	���r�%���z��:��v�Pz�u&����V#�[ύ%��������õ������|8�[���ۜ12��zfX��^˲p>0f�3���XZ�J��+�^��R�O�$��7��a���h
�����wOJaCH�@�w���jR�n��k�I獗	�~���ʇ0�Uz������ �E����@՘}�Q�c(�R�m�4��K�˝I�"~�;F`��A<}.��ױ�#�kw �^���(�ԛl4��3�S_�x��1c%*A%��o�dN��R7C�<�k�N���Y������ �c���*M���glC-�N��i����c�g�[��_��;rk�!���d�?L:0~/�U&�Dl�QWt��������u<��Yl�������)��5�,{��5�Um u��E��
�Lw�TuS��B*)����ȫ��X���uϟa.2�Pzs���Ҵ���a��盚���sZ!O[���̨���^P�v+\�'X�0��w$�U�ME�҇�����o�֤Q��ڞ�Ac+�<k~����������!��bN*���̈¯#Qm��{l�$�j�GH�ʅ�2�|���tpod?���n:h���lJ���:�i�� ӵ�����)5�Zf]�:4pJ�K'OkJ\ϺD�M}�RX]�.n�Xo�������f@~��N%��2��n�������v��׫�N���S���b*Hb�Ì�|u�ѓ��P���#k,OIk��Y�~ �$�_\��(%�F[A�S�C��]�x�8����u�AQ����I�M5d�uV�9u_k�����&�ù�?[[��s�ͣ;7�U�c#
�S����<4%����x.ؔ�����W�;�Η�ڼhj��IX%k&��5~p�N�?����i�2�E���b�&*�M�ۄV}�U�����:&������7����{Ă{s��J�[Su��[?i�^>�2�}J���=d��`=�x�1��cNl@�a������މ�)�Z���H����M�o�q ݭ釖�D��u�5�a>�J:+!����ò]�H�yT�A2��XKy����d���
���8�~�	 J�7����z�N���K�����q`YF���d�t�.�v�\X��s[�A����Cm+�@�;)n��B��	� �n\�Q�T9f�H	D��ïUx��0�F���`}�Q��[����	�<�}���H���֒<sK�(���`+wu���9@��=����
�-鐿�#+�U�=j� ±���g�¢T0c��,��팿�{�
�W�j���r|H�eЈ�Q)�K/�9���1O���0� _tv�a0}A� �u@唷h��]����0e\"��A�c�Q��um1md��̆�r#Hm��a�IwI� ��N�����u8>tϹ�{��Ae��zFl��a	h�{f��1i�8����Y�M9a(�9��-�x���h/S/�<2I�2�6��<Ǯ��m�[>�Ch;,0hI|��	��x���#� a��_8���!�P��$ܺT
�������3"n1p��i)���FʋA�Fb���C�����x�=��0�'NA-w�#}�>��g!則r���?�6j˩�n)���z�0��nڐM�Bx4��(�~�xD&
b�3E �	"���5��0Mپ��(�E��؛O��* 12��*���F���IAF�a'�����00>Ù8��m�b.1G��=�So��w�k�~���jv��#�[vbŢ�x�d�˖�������aYhcƒ��o���q��6!cBf�Oa�����x�z��~���h!,���Y<U�G����훶b \�c�����.w�Zr�E�|'HBf�߻�و���������v���Kv�hDШg�����K��}0�ݧ�	6A� �3C������#pw�hS�̋��L�7�?��}3�X:�rby�wƳW0�����a�tL�?p#��4�U�������/)� ��Mr�yZv��	�8� ��������a���(�C�5ҿ�HF
[�|��22`C�����S�֛V�����-�_�O��/H+���r����,%�z�G����o1�	T]��FK�P���a�`�S�(�K����V X�a"฾uG�\ߖ�c���?MX����Ģo*!Ock���.+�-�}�~�7����2T���a������E�Wg�9�b�H~FֈP����>8MX\��P3C����k-t�{㼳�
�G��Z1� �V\nL�O�e��>��o"{�`o;Wα[��������5B3h���3:l����I-Vfv�x�2���b��4z���	ȋ��<�:8�QP��o%]Y�$䥊���3�Geo������N�i6\۶E�ҝ�4,&	��d ��t����9w���	���/�W�x	P�w̩�l��W�[�o�����
=V%��}�h&�e��3��%��f3�OȌO%�և�̞r�l�Ӕ��GԮ����6����p��%O�;�㕵�(��'�m�W����~��s��(<-W�gXb�N^/�5}�/9��oU��0w=�wI�jD�m�7y-l<����	���
��*[�Y����A�]�J:�T�a4}�y�!8M} ^��n
�N��y��L�X1�A�x��U~�y]�v��-幠w�@�CZ|?�2:�!ʬ��B����_���/Z�$����K��Zf���[�;�O`��ʹ�J��k��u-1Q��q���i�op�P���&zF�)�6G�XiA�Y�v=����Rl#ɼD��~�ш�0�L�@I�C��J�|�Ӿ@�j���k���{Gے�p��u�8����3��霛���43���*���Ҿ�%�|��K)�X��8���"��Ia�/�
�z�ʮф��n	s�6����.;PQ����<�Di�n�GԺ+�^�Y;w#ʒ��
���v�:��P���|�g��}��?	�&�3�U�S�H�#S��X����UA�e�'�O���\�0�1+f6pUylG媴Ru˽�6��1�J���6E��P�M��f7b�+���hy[��DdY�&��oz���g�oy:�!JÖ�쌠�J�]3d�u�R2��=k�J�������,�3�%i�)�we�x!��	��ov��5�R5�^^��+�q���I��}Ƞ�����ZB�7mif<7�9���P�u���/�_pP֗�H5����Q��ٙ���0���d�]��JY�Aa{��k5x8,0�پ:8�~�y3�p�8��ǲ���z��m��x��=R��,��2�5ܖt�Fº�����:U��s���L�櫯����o�'a �v��舦��#Q��+�6Ξ�re�D7����s*f���.5�f뉻c;���biIQe ��F�WZ׀EP� R_�S��������u�	0�XDr�F�a��4Ý���c5��ӓ�d�?�\�N�f�FN��$��y�d�J@OR�)�$���V�	6p����v�7�q:� k��5�r��o��U��7f��dPD��6;�T�l�)�o���E7$g=z���oz����4��D���g��[��T����y��᷄x�G�>����-K�>��]Hf����������.̷+���_h�U�l��n����oe�0
��F�},��.��z�����^�~$�^Nn,�r��b�
az'v�o���S��9���HQ�L~���P$\�T'r�J:(dU0�)}�T�/6v���B��.L�{���4�<��؁X@��?��N<��RZ9rx�ת�����V�����d3�c�#���;��e�Xx&����yyr9�=�}����t~]��>tt�d�s�w�=�� EQ��v`�j���<2*j&���I*!,����Ȝ�"Am��+� Šmϐ[�hDâ��)�~���?�O��^��l��r�n������E��=���M��olqn���0���R|�D���)/�7:�K����	}İ �.��i<����^ˣ�.h�}�(����F�}^��#�?�����M<� �y��x�*�6�W
QsC<�J H~vn�%�q���:���32�l{���<�o��=(~��:gk��UE�bE��ۀa�b�1K�!+Y�`�Z��tBs��>g����/jv�l�X�K���ul4��]�W|B����۲�P폃KOF�@N�5Q�wS�Ap���P}�z���#�O��u�JeQ�	�#�aXD��Ӑe[����Aq��9^'˞$�������.?���:��o��m��{Z\p;���	��U�k���0Q|h{w�	
C�"MU��72lRS� NM��s�%[�2|=�/
!�^�۶	G�����s�f�'���%��[#xȶm�l$}����EB����t�5�4m斝�t*Ȟ��m�_qa��K�K����U��ۅ�c����,�;�b�r��?� �|��5������*�b]C0�����||��PP��$�J�,�̗�ө$�3�%-2T�Bj�Lz����X=p���[C~�����a�4J�%�+uNE֯�XKIUd����I��)��i-/62��v̩i��bG3��h�LT���x�s@���将�R�A�t�G�$(U�g�&��NEF<�bIȃ"��%�gF~pk$�$�*�9+r��f�U��7j�{ׂ����ۂ?�Ϗ���.�*���	l|�kH��1� �R��NM1nW;"���)Jh�J�q���_��6����=!��=�N�eO�4b<�]����ѭ���*y���#��w{�������uj�����^I��� L���@���( m�J<1([�QG�ÁnQH6ZQv	5��)	��Ah�Z}X����!��~�*�>�hSG�ʷx��/1���P��6�HVi+*5���6�`@ѿ�A�����"�-�Ls\���p�!���u��GCh�O�'ŲN혹�}��X���r�- rk����:�C��ۘ�{0wy�S�J�'Oi ���ޥ�Շ6�2�l�e�7E�zі��UNx1�6R�֬,�}�Bte����ɦ��U���I�%0��:#�Zx{;'��m����]�Ӡy�ܓV.�6w��1�����h��T�SrӒ�x��B�=aOfW����Q�"a�_#������ʭ�����o,�+	�\��7��V`D��@�D��E��C�W��J{�"O�z>͓�p�&>������.���ڍrN�o������h��݇iD Vγ��v�?{�2gp�����������E1���*�r���&���%eU������y���k�vE8K��!�W���������<kD�چ`��Vk�U-�bb��f�<}�V]�I���HnW�ꋇ�tA����@п�xg+f�Y㙨��J�sf䍠�U0�>!���P�u07nA����@Hf;Q���eC�N�q���E���5����M�`l�.A�F��-r�V4��g}d�� ((��tp&V�|�KGdô��H������;"��R`9[�]�]��Z�l�7; ��K������#��0-�d�UюIoM����df$�@��R{8��˛��î���wqaw�&��Z*%�0\�ԥ?I���E ��ow;��W�KoO�D.gtS̝)���.�洑�s�4��.bK0�@3�9oJ��*�&a=qt)�#�1���^�5��� #��C��� ����J`2��Zb<JN%��$aJ�`@��̮��k�]d"M������x�&<�j�~��e�S΅�b(����\�W�0q���ȼN�9#��g�IN����h�`$(e6�{3��/�M�E�e�B\`21a2;��P��Vf�.�=1�ۂ���n.�JAaDA5,(Lň�r絙6U{��ks���}x��!Ķ��!�<���,�W�a�4X�;�T�o$قü<~�rمa���~>"�2��O��{��m���Ak7DI~`����[��0ܔ�ҭy�2)7dإ ./�B�cM��\$�8�fq|,��4����� �3!�b��L��d#e�"�C}�}굆r�Z'���p�jŲ	��ߓH���9��B}p�З&a����K�l��%�r���c���$��|���!qyK��CsvC�$�r���PQȮ]Ş�Gؼ4���3ƮS��}�wk��̷>�>�����E���~�l}A0�c�Y�� �ǭ�iwl�E�iT��H�;J;�׵h,�z���s%1�F[�������(�Poqs�'����� 9cS����KEbl���'}���[�7�T��m���(�iwpy;�0��:����O,��� V�{a�r��24܅*�J$.����7E����z��%2�;���R�_g���,v����_�[B�qr�����[v*֚7�i�(���r����tkhvv�ϫԼ	�	ZݕS�i�=�@��^Kq~�[���%d�������:���$��f��� ����p6IU��d���z����������Y��x�
Zc�D�Q�&�-@�B���N��r�v׈�7���#��BUI�o�D��e|8�)G���x�	�����忂����P4�)�\`oDܞFҩr�S/tk���4����$��|�������Rĕ��OV������m`�"7�W���A��Ψ�M~�,��0��x5�Bt��Bc�{��t8l�^�6v�2A��F�~<gv��v�����e�-Yf6�i��>sz���0Gs���G�;i�^^n�;�QY�",1��nl�֎�u�� �"��W�Ñ����/��5�<�-���t~���Cv��`�خ�x#Ô�ԱU���xꑊ}��SJ�B���J�����<дJW��Tı<#B|Ev)Bu]j��#?�0�L���G�S����o� G~L�^���V�:��S(��JU]Z��\�n�+�ݗ'i�MTwUh	�����;�2��,4��OI��#>^e�N��>Ɨ�!�����A�fo���|�6J�kB�#_�iY��XO�j\�IJH������3�^���,:u�)K��{̜.���F���P������o�*��P��ʼ��i>�@�n`E����+%�������:�ZH�ŠZ�#[q�>r�	�2{�0�L�ȫ5��W&Z����>M�-5�NCD�^O����x����:ݶ0h���i�Q�oWK�Lz��������P� <�k5f�mٙ[���n.5�Ki����Y������@	�I�%�z��/�N=Yb(�g*��q�����)���Ӽ��i&�*�ʣ݀տ�>�$��5#q�t�0�V35�>������sP�^Q���:^�����-��((�?♚�<}���q@�fL`J��!�)A��j�"#0"-�X���ֈ`waڅ,9_: |�+Z3���$�6D�f�VB��q���*.rx(#$3ϴF�C��&!jCp���M��G©97	�5<j�Mh��'�+gsA�����5�ʳۧh��?U/K�gaԋ�e�a��l�";���#��n�⬑t��&T��Bl�i�{��A��{C�=�(-=|2	Wi�[�H��K^]�b����QG�|+hkX, #�����ø`:�k#?z��t�[v�"�d��À�)���sp���ρ�I�o�E`��[�������嬤} 7r̗�-N�����?�r�����ˆ5*X��������%(=��lX��%5�8��&}��_`�N�4�FZ�l;)#8�BPd��ឈZڎ���z��I���FAek�u����+VN��GJ�G.�\mX��`}<�~��a9��ٯ��8�	'�Ju����/(�{�0,L��~�!��M+������,�mB�}÷��6/R�	H۱�Γ9\����*����*e�|� K\�V �����Ц��Cgp�W��5��FE_*W�=���E��	�m^���JN��~G��'����.���d�[�no68�;.I�4%YGsnO*�mkn��l������1�B�_�����8ȏ[6w�u\�M�M��ظ �" -�R��b�X��vH�����RȤ�����Ǫ�����~��+�ժm�s��|_|C���X����$�N����	�T��j|�.�=�����I��mb���������kl]'��.����;=ݷ���z�8�VT��
) ��6�1�1�h�]��5,��=#O���|���nt[F��~RV �0!GL[a�i0�fv�S���>�ו��NAI�ga�9@���x��I�Zp�J��OB�Gf�����	t`���]��3��)�L&�s��'x�� P�y`��t��Ԇ���e�B�ōi��s�/����91Ȼ���1��T�7+U>]ȳ�f�6���'�:��X�L'jiP�6.g��U�&���۾N�a�-C�P�KE}�l!�{8����t�B������t��*`�7�sP�A�|&�+Q�9L�}]��b��"92ݛ�9�u�Ihh�	���pN�?���1�^��"卯�8�QV��K�t�GDz��V�����ⲿҤlb�$�4@&�2���3iO�܎�y�_��`��e��,��v���B���ME�e�\��}RdC5l�;���[\�3�֪���N���?�iE��$|�����ڹR�v;l]Ҁ��oia�h���2y�ܩ��:4�kd�Վg�poh�+�͒Y*Y'�]ǣ� ��5��Dv�x�Vc"N�ڃ�Q%na�bv'Q�a2q���<��N,]6!D���;q���	R��.A�6�K�jwV�[IxT	W����$���ۿ�Ӑ��^{�^>�w��2&�.HAYj�4N6�F\�:[�'�ҙ#5���;�<d�$��9ڀ����޿�1��U�urqZ%�ꭇ���D��^�=�D�s%0D��G"�'[�F��$�3_""��;��P�,�x�Pb4+���+�Ap~m{�Ғ3O>0�ݐ+��P7Ć>��R�t#	
>���Du>u����������<��2Us�n�YÖ�Y�(9	�+G��2
&iV�O5ʀ^dR��P.u��p�Ł���nd������R?���Y��(>�j�D�׋*2�E]�t?n��j�|d��k��V��s��O㖷�;�	�o��|u=�'��=��S�8ֻ��6��hVf��T)'�O������s�K���$;媣I8�бP}s��=?�-,$3�S� %�o��J���\���}�Љ���ط,YPߑJ~u������h�9p��j�]�8��t�NQ�r��C+����5���;����Τ��|P�D����P������ڝ��0O��UȺ��c)k�e#壓9��K�?0�6}ߘ�l<NA�h>��f9��%�Bm[~<���C��>�dC���t]��=뱷����3~y;�*��K&���%���j��m ���m �=�������~��yG���(�rdr17qoe�x�	$��1p+Y����;�I�-�iA�B��<�����3:V:�㔷�M����a��r���5� �Ù`"��"�/jб�?tf�k,��-�BVV�o�K��>s"��ںԖ/�Zʧu��4�m�ѰS�l{�9�������й�|�k�� '�dhw��C(������Ε��?�����t��!1"��z�T�o�*6��y�W�3���-78�(J��ۄ[�IS���w!%�w���nC��n�G+չƾ�F�]�C>n�%����N��w��˛��z>H�^讓��AF7^��@�<w�����*+���Y�F��_e�+�A�j��~`�;��[��u�W��U��?�MZg�X�+�F^�Ɣ����-�o6�_.`��r>YM�Zo>C��9n. װ�bd?4��ͭeM���O&GBL	��<�������p���$ɳ��#j���q���W@�iA��-��V�#���Q�U���0�=���RT����-fuk�;R��*��Hd6�"�&"�X��'���ib�~��qX�/����&��fl۳J���F�O߹�-��׶���֬��!���I��B�[���~���������á�c,ѽ �������窭w��2�#Yk]�q���2Q��o�X=����;&'?�Z^�������G/A^�n�!���(;�@G�	�t�f��������gǲX88������<�Ck-^��i馂��0X����o*��-�s���?' �yB�)v=��Hr����=����3\Wp�ǩ�j���j�":�~�EMy��=s��?-^:�\���-}����V5���J�kHD���6Q�ݬ�ׇ���
_����|�Ȩ���֜0_'�*u���(ч�ݬ�G{�%���"8;jg�^:a��/�|�|et!�����Sr�J��H���y�:�
�:t�.GT3[��Q���A��"���G�؝�O#`��.$�fa-p�~�9���g���2Mt�7"夸z�W��P�s��~�75�zc�%�M�ѥz2_��W�EGKT��qj��w�?��7�*��~�.C���ƣ'��)�حX�����ࠨy<�n�:a���C&N�g3������!Bx�=|�X�k����%����Q�alx���,����j;'��en��A�S6��D����g�9���C��@��3�%�+Y�S�L}y��� k��L� N�?��f�9�ٳ�ʰ�	�$Ǩ��������@� �y�P� �;����q!�[�E�ޒ��[}90��P���Wo����+�D�6���e�_vIlx��L�M ��VE!��Y�H��C��3��A��f�tyT�L���v��E����L�8����t�f����R���2�\!vڨC&u