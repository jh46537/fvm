��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��dm��JP. S5&�Ac��<r�Դp��������#�
���<��?�8" ���sfD��m�,F����S�Vn��8]��A4F�}�֋�;�}�5q0����J)��l��=���KN���U �A[�z�� s�:F	� ��O�*������"}\���~�,bp�(�U�8��$ŉ�܎��Q5;��E�'�y�> �z)ih&P�f�N���_3�*�x�H5NJ��͗���OxL%V�>���W�)<el�Om\��D����'�Ľ0Jt��!��#fH9�@l�8�n��b������U~���Jؒf�q��D��!������;l n��%멱�f��.X%��XKL6O&.�5����|��?�~qt�����q�v�.$���$��ҳ�Tu�>�pD��R;Z�Ϡ�l�0:�����5�&�����$_��:�eL�Ja��\t�&W�mE��m�ЀTs-�~�Ɵ��{�a��2#�N^�K��%ku��rx����	��ad.j�3v����?��4="�˞*����<A
�^0��5�'Z��\%�M����g���h
$Y����K������	Fm2��j�g����h� Dj� ���7q
��]D㹌��� m�kI���hW%M�Iq��(xg��Y�Ȼhp��%�l�O�@슄�O�_mڇ�)��Z�;~�4�kA�,��~���mkQt�<ɒ�+iB�5�,e���^1�=4�U����l���~�9��5��	�5'�w����?	���J�� WמF9;%yd�����\sq�'�%� ���Y�x�����-����ה�O"Q_do������.�&�j�{�
7��Z�c��߆���M���s!�t�1���]�����]��Ѽu�U�*`"^��Vz�q`)��
��#��h���'P���|5%�Ch��vy��5*`���[T�Wa:'��2��SUU�I�)��v�ϼyZ%��ܡ�V(������j��K��� =#��=��y�o�����P�g]��z�Zα��4'<J�LP�Z	�:��G�[�� ����w��v��v3v��X���4�1ǒbe�̗�G~�_@c�Y����MtXW!�1s��� ������35��+�>b�\2�Tb*ܣ>3�wa��5H|� A�q�WR�y�+3Ô�e��*PeM�{�ӾH`98�pP�J�l30_�E�i��)Mc�_�}� �b��ɶ��iE�2	��ne�v�I�AN�C��>X�&#�a�W���u�,^Fw2*nȅ�D��G`K�������/f�f ��r�5>��ϣ�:ɆM�X�'à�%�D��KX�Z91�Bt��n�s�ù������L�E����t)؊�ݯ~��sn�]�D �����@�j��]�^���`��g��zɦ�NԨ����=�41B��ɤ���*z����'Ve>�)���lC	:E^����Rt�;Q��2����Ё�("_<�4�l�c=���W y����Z�,�uu����Ph.���Vi�s��� 5{�Q��[�<,F�)C�8���!�����e?�TdU�B2�)a�Y��L�w��[���0W�s|r5�@���q/��25��o�nA��3~���@Y�	����0Ưi����g�z<���Օ��z�㐎d���i������3�F�fHE���F;�ih��wb�x$�{����b�&޶��M�k�n\��]wӤ���g?��k'W[��t�X>5�o�`��Ӈ�j���b�B'�>M�`��v�#��J�&+Ёҟ�Hl�+Q䎈�Oj����D��mj��o�p��P�M����T'�ڙ@����ɵ)�]wN��{�s�$�7G,nM�6�оQ��ziR���FʿƦ�"Jxv����m�Y����m���.^6FN��nK�|庫���{�������p���鬈R����ZcQ����`>��2�v�"͏gz=�G�Rp��w����ͩ�(dꑢn��1�`X�L|�Wf�
%��7U�b���;��H�=�>�ko�-7���	6bt&�Ɇ���x{$��V8]J�