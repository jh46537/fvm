��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]'���,V����i�E��qd<���2���U���ǵ� ?��K��D��,����W�������:w��|�� )���%�c��L�~&k1�љ[s�o�������@�
�+�۶�����1�LR��XI�c��x�υ�$W��N��2U�����AGDc�M�x{����~ؔ %�$T�]4�
k�>�)V��,��4}зj�}~�`�|��R�s߿8���s���+����wm���w�F���`{K��̆����N)�c��0���k=~fV��k�m�#T>��Yg��	F���7���V�2	[g/�[،��@,��t�N�P1��:k�>{��.H(����=$V��	B����4�G����㬐�X-
�^�}�������?��	O}#���Z�(�hp���v)���zm��L���>
34N��1���ͅ���?��I���';�=��պ�"Wb<)�+R�m���C��'0\rF��Y���̺�ն���Gj��מs�5����k�-��J����6Z�=@�R�O���X)�����
����S��K�=�Yw�#�s{&�q
�m �Kӕ��V��p���&߮��-V0������	q��qn5`�f�Ы�(xpw}EC�V�M�G�o�p�������N�6E&ZM��gC,g����?S������<��5�?��Ë���F��l�.�I���#��LyD�ZϼW&���#ar�czf�z�KG��z�
E��練��`6$�^ΘoKk�
����Ie��@_H�4ZCgx��%�}m^������_��۬�<��
�v;��I��,CG�(�a~�=�M�k��-���� ���u7�?,�ɶ]�w1��	c�Օ?uQ2���>��O��CPĄ1"���1�9�q-j-��^�?d܄.J_KK�8�4U�i����W����ML�;$`��� E�T�Y��'��ϑ��dxb~�!��>ʜ��B}���=K����@%�|�N%bX�U�&-,P�� z�,|�(8M��*�"��1���e����EO�=y����R� ���UΥ���1��پ����6t���U�@J}g�RX���NZc����S�LG�Q�k�-p�\��)�t�%�:���I�i^r'_Lo���S�]u���&�T��Nbw�h ���
�j*xV�K��H�SՑ&�|�Z��y�+�\3E��E�xɡ4���t�d�\��I?���&ˤ�N����A�VG����BWV�h��]m��N$bm�����b�!��#*��*��C���f}�A�D0� +Ҍ~\CP��p�@#Eq\��L6�Z���	3�l��J��'��Q�F4�9<.����䕇��E|��{�5i����Xr�kՊ"��P	�a�O���c/��Hbp�6�r�j��������H�xgb��+b�Y��ګBX貏_`�UiYPz��2�pR� �Q -�e�\v��� ��Hr��@�Qs��cdp���X�Z�f뇎��7�v˝�r|OT�h�b�ñaӰmq�qJ�ҕ
�efF_l<���N{ҷ��F.���:�o]���I�K�I�9t���+������j�w@���Y�{��T��&&��l���D��fN>N��T�{dl�x��{��!Y
��L��B�{B���� ��XDeۦ�נ�D�fzd����w�
M!b)�Σf9 �" �]�s,(�^s�]��6�OK�C�C�I��ń&��&�1z���[�&�iN��86��`l'�-��o�m�����ԀuO"p��w�J�GK���3+�Ϟ���-$�ג�����a�N9a��T
�J��\U�D��V��lY�G�p�!+�I4�ܣ����E�0�'_�>MI]a��K
}��A��&�o�:~CxR�Kꃻ�#��:�P�­#OT"ZȤ�M��*\���\U�*��F�'�*�3P!�Gy�7���E�>�.�����PH�?C�'��W��J;�9>ƨ^����ŧi�O��F �i�B4��IJ�K��uЛ����r���-�I������\�3��Ǚ�^�H��t
0[ؑ�?�o�G?�m��)�ǯ�V��/�fS��e�a�g-�#��� w��@�94�-8�ϗ<y�����>�Ξ?�:u�c4tOV�mi������68]+]î��.��70|���KR�" �w����.1�Ê�vs;������2=x��Ά��Sk&�ϒF ��`i��VAU�A���2ca�_кݙp�z�XC%��!{3��Ֆ�����Y��6��DPX����i>�|���"�����������F�����d��L��B�� �|>���y����}��ޜ��{NA�9�CZ!�����C@+F^Zk����)���l��G�&!�{��,=�/���
X����\XoT�.ݒ�ʃӚ�g�6�W���:˻��)������ʻ]gҎ��0�9�
7[o�\�f2&�L[nӁ���IBk�em�����Zt�%��BDiy�~\�c5�� �e8ة�C5i6
��c>N�񥃫X����H�`�sF�5�2�H��8>J��>��X,��<���yĩJj�=ټA�MK���6.7�b���HdSUQ�J�W�$X�V'�4��c��Ǖ�,���Y��tH=�Vr��Y�fE�=�M�s
� 9����{j�%���3�S���7� ���8}9�͵�k��ϑ�A+�%K���]:m,U���<0?e��-����"!��.�V��i��QHN��|�O�>�VG�F�� ����9M�i�mOѺ!� Ub�
�:ȝi�TM�g�q\�f���D!�3���f�9,0&���0��}�(Y�Mz�RUZS�H�%by��kz�R.Qp~�����{�qp^� u�?��5:��6��O��۾^�x��C��wE?`��[H����~v02���ԟ��g��@��J�-��h��2��6'��J?:�~,8�q�:C��-&+�-��>0Y��l6��� �~d*��c%RJ���,&�di��S5)����n#�Eۖ��4܌S:�g��Q���2T���K�6FX�<q�BIK����ۏ���F�wL�)����fa*P%I��p�yl�?8H���e�i��~¤f�,��ZL�kĚeʁ{���+����W4�S�/Hnھ0�I���{k�*�Ѳ3�.Qq�y�v��π���p�U��I��2�T���l�V�L��%�EX_���`ZK�	�JP�@�["�y}����N�k<�����^����H'6��q{<�r���3��^B)��Cv����# ���=5%F8_���JQw4�����5*�/���D��5��>7�����z����p���SN>�[�bi����(���l%��mt{3|W�mg�#)�1���Z�� ��t�p�� >�IYH���TI�����|�"Fz�U���ھ���~�$�(F�N"��p/�m3��B9=+��j^�~�Y�P�y^��E��v�F�l$��S]H�M< �#�� w�{�8��qzv<� r��ж䣇����"_������XB��l�m�m���:��|���,�������Z��J���x(H�߾�Y)�q���3*),I��:}��Gq�������z�f�K��t��D�]��cKZ��*�%(3�+�#m�p)�ͭܓC�iϽ��g){[	{03s�.��'��5?�a�93�nP:��F�A�� 
�8 l~���,�}�H�/J�*V���p���"� )X*p��=�Ȣ,�F���ا���:`��z��dѻ�n+^�|A#��C#4^+�op�k�3L�6%
�7}"l}� .���Y���ӵ�!�P�m%Gi!�@�y��?Mˮ~pr��{��#�;�éV�W���S�Q�e�Qq�PcR��V�35�����K���R@ݥ��`��+�=���4A�Z� �'`�4�77���%/���X��W{�/f���H@�ڽ�>:�y��$s,���������u�M�D�x�7/X��V��Y&�Yyhm����Isx�M0��V���ە���,{%�&�b�gQ���(��Q���H�Ε�i�f�1�hG�e����$?pt�>r������1���9�?��x�4��ܘ�z�<���_֊ao����^��~���
�MƗ��8���I_�x�����#��1_D���e�Ifg(]s�67�t�nB�� O,�C��4��a�*������<WUB�=���砕x 4}�s�L�G�Yp��4
���R��e�$}�������N�	����;@�~u�-��l1Z�}���Vgn௠���u�\	��g�2�h���.�Z�V�/���<tE�φ
�G����n<'���a�أ>W���2�7 P5a�G3���Qa4]!�c
F$:�hCyj/C�&Y�5G�򼙜����z�s�f��;z�M�FM��|����[sCF�_F�+�lJĨ�-�V.#�~��AD W�0���wP�!�n��L�sB�G4��˼Ǐ�h���W�ι�N�v�y����BT��B湩$ߑnH�:�<���Z&� ��_�� �)���C� w�����mY"Һك�����/L�,�1�Ԋ��8`:����3|@����K�,?~�H4�_�8��P��{'����bFJT��i�@HF~����b?��vo�@Aȷ�P�c���i����E��O�*�I?@�M�� ��jqMs���m������E��z��`>48�C�3���Ł���H���vm�a
aǊ�!� ZW�hđt�:_0��B}����'�z$��F5b[�X�R|#�̷���8���-v���y�c�*��WՁb!6.(����E��B�\����p����I�{g�_���p�9�!f�T�, ^�*C6A���~)�!�P�v�A�.���/Վ�!6�SF⇠Z�g�*w�튝i̶0�L��A��1`�$�3���W�
������e��ٽ?X��nb�2=Ee)c���o�"E~�O��M�wyb�&�~Й�2Fx�s�Ә�O'��<�������f4�X��eF�,�+����=s��!��냇L�K�+��D�:�f��B��9_79n�~�p��j3RK�)�pxHo��?�9���������4Mfam�+ �����
�N��Z����A-S%�RcЬ1^�6�?2Zhk	�6��L#k�t����	j�X�Qv�� E��[�K^�v˓���h��0����0���Fh��L�$Η�����o�� ��2@F�Z�E��~?#���&�'R�5�*��(x���o�1B��[�F �>T�&�,bQ�� �y"N�︛���6�n�P��K4}���1�)�M=��]��d|��qX�^�f�\�|�T �ns�̓4
��vK{�/1�z�f��A�_���JUX�?��hJkS�ʋ��NG谕y��}[iT�I닇s��+>�J3+���_�M�^�q��!h��`���8:,%�=Gk����%}���g����/�L�nQ�9�A`�O	\���/~5,;��kFǤ���`>�0�d���́'u�������3�J2/�a.��`�!���������'��k7�cR��@n.N�-,p0�+�;ߵ�}�����@�ʪI�(K�"�;��X	�<��5p!&%<�)���I�>��[I[ӻ�sB��rZ˞P"%�Sn��@����3ct�fWxP3�&<l�@m�I>e<#����6�j�u#F~�ES������xf~�j�>;�d��}c���bL�G�7ݚ����ْ�PTS4�><D��]����������hT�O��)������㨗���b�Ӹs��'��k9��͘��h<&�:5�*��4�T�j��9�.�FKu���G5OdE��˧LJqs��R�%�b�@G��c��/�YE����RE⎒5�x#�H5v�߷2�P���%ʔs_!�/e�f�O��y�f`JG�������g����1��z����	5K-���\�����o~�(7p�N�xo<K����9y�Z� ��Ӫb��7ޙ$��\c,�/W�+��_��6�j5n�sj�
o�>�bN}%p��Kl��1��E�I�/D�Lz���ȡi���y��\�K���X�p�=��ѲK`%QaY�C&�w�t��?��W+�Z��j�t�Q�uh��?	��_�]����I�'�P���7c��@��Y��X�$f�����I]%5g� 4�Ub��i<��]�/���������?�S}˕H�$ i�F�R_c�j$�,;�EnS3��E�w�[-�M#5��M��/j-"�<�L�Kk�����ݻ8+�Rrd�v��kK�c�oЕT��bRM$�n�����%�>���J��^��'��z�)��dg�(|��tA�
�{����[�$V�_�����b��w�Q�9/p��85��M.^�K���W 5�!�Ν�|��H(*:��xj11�!.Q��3�/2����-��#���4U`�3m�`f��FC=�Ϸ܂�����SM%��8��~<���f|b�Ah_�8T���)������,���D��S3�hπ����/�Xq@��k7c�=P��@R��&�6a� ���NO<��bۇ���*����7`�����Z���a�
��Ծ�ׯ~1J\ud�C�%�SʊcS��*N��`G�k�
���H��l
ʾ�lC6�f�w��i��}��,/U�7�����l�wU�F1<L������`���yn�؆mپ�F��R�X�ε�.�!�<Y2� ���y�@�a,&L��sr^`�T���0iHkAw�(l��	K��c9�wၷ�w4h@�?z?� �W��e��!J��w1�˝���.��s/�i�N4�aB�1���7$���߸ 5:���P��tb�(~�(����ѝ���r����A�l���"Dꕏ�0�n��~ k_ R������B���B��n�e��"�¢R�h��������\��
�����C�dN���N���ZkW� �Ԟwy{��#��9:1&z���?��o`h�&w�X}Cr���9>A��]�#�����}t�||ʨ��Je&�}ȫW8�I/2_|��QU7�$����̞J���B���PߋJud������t@4�&L�1�p����1[xM�E�;r=S #<
�K�� �h~ų��\���׶��z(��DR�&\D�H�s,�P�����DZ�|��_|;��cw�$[���ĭ#W���a�����>s��6C�K<	,ڌ˖���Q�mWDd��������Ê�q�ż>vOJ9B�N un��2��EOߋ�j!��ĕ���G����k��������C�~?O�~�?=۴�P�~��)%Yd,��B	k'�GL]�%h���ƌ0��w�HRh�Eb��m�e@�����=ܥcD`z�Y��?�_�FmW�
��ܳ��"Ĺ��3 ig��g�]rw���*�W��C����[�)9��`���۬,�^�9z�Ǭ��=�|����w��t�7Ǥ"��1�i�Y���q �,U(�?�狖��閍 �A�M��59[��&��M�&"�-û�4�"�3�{jU>6M!�ᐳ�t��C�۵��kmK]>ȵ�i泧`�<��Th�}G�l�͘�d=.K�`r-�60$��R��K�k�H�!T�����!;y�5�U�������h�d�P���Y�)Ȋ�0�o.�1k2��h���t����>��i��ܓ����>�H��[��Y����{�c�Ԍ�K���; |��"�(3���mV�
��9sϰH������{�%J�A [r�G�	��t6�y��w�f�7E�BTa�z�nOY<.L�}�C�f�dJ������@����.�j &�Ņ(u3n֤-��C�C��{09�]�ח�u����2@П���Yi��At�Ӊ��X�9H�ph�y[��Pl��796S���h$T��g|�B8��_L%��������X:�����7�>��KD�R'��H��%�{�yp;�!��e1O�\�!�l➳%1G��R�R�}b�v�0�����U�왯����ŭ�g�ҟK����+~]��<�k���o�����(9F-����~��޹�Ֆ�@T,����ݙŦ��tuE���6"V���YA��':�D$LDC &�������xx:ÙeJ+pz��3i�7��g��D��ޜ�?�'gS��~JI���xk ��o�:u@ q�R���U�a�.���7��^J������- Α�F�o��|k	`�}(C�\�y��k�J�~�$ ����ls�:���$=���X�nH�~��ڴ����o���  A|��KPW���j7�� ��xy�$m��_h}��Cs��x��"��7;������ 0j���b���#,iS� W=�7k'��4�4U��Iu��������B%`�p�q�U�Q-�&G�O�3�$/���~_��|��a�����9dZp����7'@z&���t�ZRM{=Z�f����1;�(��0�b6�������x��Uqptl��K���]BO���㘿O�wҖ�^ϫҧU�#�P��|��֦��P�S�L��kl)�0��T)���(��ޤ��OE���,I��?@L�&O�R+)�E���`�<yi��7)��ç�#}5,����O��R?�� �v[w�&Y��e����0ɮ��i�ׁ}������K��C���2��~$��M�8��$Jx4�'�Յ'P��/4��h|'԰�u��3�����Xx�+�o�{�┖�����P\��n�`�l����Q���Qʟ��w�@�ƽ�E�a4�aK�ɂ�''�Gw��MB�8
�~Wi+T@�oӐ�:�A3�)"�K�S�|�D&�r�[�j��2jX����?�9�NE�W����W�J����.+*��C������k(
rމ��-�z00.NqxE��A��b!��eY�J��9:���Pn+�wF.hsbݐ���æ~���'.CX��Z�F$��<(�5��m>�*C��?�t~��95"���	s\̣Z){$��+�H.}t�జ򹫧�)J*ݟ��_���
$����<O�ډU�{n������[c���"9JA,���<��P�wI��u"�4�1nޗc��Q��V�c�?:�Ԫ!\]7�>g���b}F3e7��%�z��@�>�8$tls&�Ҏ�4�-�����"Öq;�1��d̡G��z�	�.��V*���lI�6��Trj��-Cw�J<��-�"̑ϋZm���3#�q
�|�p�1N�9A�-(���$���3*��6�(4\i�p��aGV���D�T��Ż@�L���<�q7(·���8�i�K��g�r�U�֘��K)���<��;�<$��^ĲU1fu֘�0��]�l��h�Ϩ|��줨_��"��N�.N���}ukeU�6h�*�bc�>��g�:jz��9WPMS�Дq,���hb@u��-�Ԡ�f��ѵj�ӞH�ר��m>��1T��4,l��髯o��(FC���?Xm��?O�8zX���=�7�ޖ�u$J�~��]+��"��<�/#��� ģ$���]�g��m� �o�߸��tD%�~�}ė�5�a��W�&V~.)�a/�'�[�R(��/�����$Z�[���$�����+g�̦g]�!�g��}�X~���ioR&�T�.�;{���{,�[�5}���������L�9��ܮ�@04�\،U��Ҭ�bݐ��!��>`�,��Cۦ�$D���򕌊���XK�z�mDK�»�G^#�N�3V�n��g�o���͖��z[#u�:ZF������������ҭ��ƥ1M�Jhh�*�k%{X���.��[��yD��p.� �����1�OuM yr�5jNM��t�!y�_,(>��i�V���]>�V����vj�;�@ +5U
䟑J<-;� H�Y�&�D� 2X'�=���_�a�}��_�wă'zJضM��1(�lL'�F&���;^���|(ѕ�}���������H���=�a�Y��ic6֨KǼ���.!��t��D��,��U]�!���WiC�sE��M@E^	�Du�F� ��<���6���J��������\�{L�@����<�+t,=��!�_-��Ɖ2�lI��7�f;L�KPW�}��xo�iT?,"���]s�o1t�&�6�m6$,/�P�*Ζ����a�Z/��֤��Nb��,��6��agx���ԍ�ی� �(m9�(7�	%�|��+�ӡ1kB�6�9#G9S�ħ���+�c����c:Gd�(0���\u��V#gݜ��n��9��9�����,gB��b�r}W+Dy=<bЦ$�	�6OBi�2�v�@n@��g�SxLˤz����ǣ�v蝣�����s?���l��X�-%X�$^[�N������B��:�>0���@����eJ�B
�����o�2���)��w��@ 4�,߈Em�l��J�%��csY�LDd��]����Z:�A)�8��Y� � �ќh�J���1|
�FGL!���Ub�i�*T�� )��U�H����:��K�J���0y�KP|1����v_��-����"�(q��m�r����lC�f�ꑋ�΄qG��$%>Ҋ$��oҕl���v�\��,����.�_�1���-Ë�l�"O��Iq2>�l���kml�~}ڈ}�z���g�L(�&��/�A�#/dH�Y��Z��4}:XK�+�w�m"`�<���Cy������^����n��!�������)b4�T�Y ��	N��$�9b�0S���+�xbTw2À*�3�8~S4��?%/n�:��h��ld��{u�
@���$���"�pf��f�i��Rs��7 P����.TQZ���^VɁ�x���*���<�K�����:
̦J��k.G\,2K�2�Z�!2z�,ɻ�F��njJ@�ǣ�)nT|����9c�L����2�V����J`� ��i^C�����t5��%�Ln秿=^�_'C�Hʞ������\�.���5TPn$���Ҥ�~�@��_�Bn��t��%��ݷR�O�`8Ds�<(q�4�	�5��6�`n�M�0�h^d[cc�y���Yb_��B��<&@�w
������mR����хh-X�U�ێA±��w�#�b�h�ծx�{�������&�ƞ���n��^�G3w=!�� ���!��DȼJ^�3��?9�����X���!%�VR��N�I��F t7ܟ3؇Q�P�o�P+��Ð+���)�%z'p],��{}!��#d��˜s���[��'"K�&E^Q:�@r�#��*h�nYt`�����_�2���)|G�1J1����m�*�K����/�T����)�	�H��b��ў����x�oU����<Å�=LT?\�6�E�]:��v������n��ݷۿ'��)R�M*��_�<��q��F����� ���|Z�b��0�k����H��w�Fq�]��R�:��f G9�l�.7�Bd���T��z����)�-��2��W��7��#�;L�U��ȰN}�l����K���+��9L�:d5��.�}�ɟ�9a$��-�F����ųr8��]���>A�@�GKys	I��z1�`�����y�t���=�3aH4�=D��E$��xf�_�/Կ����S�l�I4 ��r��I#�TL�P6��5@���E�V,s{޴�V�>��_躖�hu���ه���`Uq �Q�a�ɬ������h���#�����9�*�^zA�/�Sԯ{���z7J!urM�	��(n^����VjL��V'c��F��e"�!�1���2ͷp���>}�o?|��(V��X�;=��o0���&�{G��h4 Ńvt�P+�*Y83)��?8�ˆz�J���W�`X;�~W%�t��);	������=K�r߸�η̦����H�j�������`T����o�l���C��	����l(���aTWv�%s��\%QTs^��&�6�VTv�\)��Zhr�ZY0�t�J'�]����(�9Q��~�S���6$���uƼ�
��5m��h�̻�%�w[�c�zm���r���� T�]�	����'YzXQ�&�i�W4h|�62�w<�_4����i�2٬�R�$Dp�b���bƢc���vyIlv1��ii�.�l
FJ� �u�5Π'��P�XY��0	�����F�Bu�=;�9��M�,�9+$lА1i��40Y�8��)тM�X?��U�o�D�Τ�#*�t{ՒJ��Fm�������)�s�6���o�˦�:��Z�N���ؙN�ʑq�d���˻���U�F��X�^������r俤:�Չ7v?�ʹ�#:�A��\�ܔ[�����g�Iaٔ���u��>h�a��qqfiz7w��G� Ǒ_*(�3��&�+��I�lN/N��H�#��\r��4�[?pE��2�^