��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����i��;ݏ+��ↂ0�?�ceR
k�&��;T/�h��HKIw�|��&3.��Ů��p�!Q���i(�+��gX]����\G��/"�TDV
x; ��*���1$���'�os�G́�C2�:>�r��]�#A��]F�~?:6�,Ӱ������4;Y-�����|��U]�Ԝ���6&F,O���*Tkt�Zzڠ6]�ޢ5m�IS��Z䝤����VX��@)���t�I��Ml�k�{F^��-���2#��q릍@�BF(S��:�����jm�â.]"�	�i�,��Z��GU�՗��5�P�N���Lh�����	"���>�֞=]Kd����;�'��D�Yj���I��Kv���R�]���}
�jD�Kh-��W��M�� 	����eD��p���.��8�O���lD�Wa2]8)�b�;p![��5E���I6�����>FN�,5��y��zo�����f�_p)���P�Ey������0~$��^F<)أl�Ϥ��uvLi�9���~�Jh,|FZlٴ���XҼ"5o� ^���p:�cCUlr���AD� ��f�������N��,w��V�\x���W'}���~�ʓ`q|M#]6(tND���Y���usm}D9x�.b��'��+�_��+�T�#�D�ߐŕ�Xpo��+e�zu�W¦��'�������ڷZ�~<����G��2���:�jt�ҋ�5=��y�=�";=莆j�%�צ��Z��M���]��F;�� ?�p�N�'�����NHE�n���0�_V0i�%-��������~���&r���;��;�oe���ßu�t�AEc�r뾁��Z�۷��F}A% ����j��#�G�(\�m���GH�>�p)sJ|"�j�?#��!���o{'qF#�~�FS��E|�\���~�&��YΨ�ðZ^�,���nC@d����"�T"I7��5�O�,�Y`����Yp������	_EU"�H��O�R���ɩe��Jw�B�L���T�e�� �6�~���*B�<�9�r�a��� W��\[D� hvu�����R��{��o��k(IV���������6��o��w��Wᒶ�nͶ��$�.�3�s��ɰ�$S��\�f����_���>y���K}&?�m'��,�"��s�>+;H�r�&�e�X+�q�{!A@�b�K�(V&�^+3��s���1Ű�LX%|.iX��2��>�P����Za�tVK�	�ᙜ���A���S�c��`����z;��xCӀ�/�q,S�����ۓT8u�n�9��}'lS\v�l�T��mB��J!�ʟ=���� >�<uS���ˊ/=��	p?G��7D�*�I���IJz�@�qj`��f���R��h�e�
�M<9��Խ������o���'�Z�R����P������g 4ȱ�m�@��I��d�5X.r�a��%Q�E)]�b-���+y�gz7g6nv��|�N���x�Ja���kl6�2�����Uv��TIE��,N��n��}�4'ȵ�5�C��6�ؕ�����Ż�m���MyM|Ұqb:�1�ۻ Z��n�g���,�y�kn H������e�,���C�&E���q�w�@��8����|��r��-��y�Z�ۍ`Cڱ�}!�h5�͢f�Ȣ1���w�G^�;7'Ƃ(��DFer�c�8�2A��3{�f'��fw�<�� @t�;��y��ʆ����2f�sG���P� ���c�=���X��ؚ>����J? ����ݣ��ܮT�����7e��֭ق[rn����;���κf�B�(�2,���������E?Fjꆸ��T���>�����M�yj�޻��X�:�� �Jz��Υ�e���|�[P,��>�������T��0O�iA�ҷV���(��C��P|3�ը��L4N �d�W˫7ְ���#��d�I�:S�c�d���c��xey7�qs�g�a��l�\��װ���7���K��,lm�֥m�W3X�U���K��b��Ow+[�㷥��}�m�m�B�	��]]��8P���4o��z��/;)n��Z���#ϙ�2�y�Lݖ
3��v��[�P���md�H�F�ͪ)����Fug���^3����yDKqw0P�2i޹��baha-y	�jV���`g��8�#�g(]��G�Xܨ������{�h;�C�����"��Ls=C�2��3�iԊ��+�Pe�jv�܂�	^'aW�P������w����[���i�|�W���b��lSڃL�i�Q눬·*��F(+ۙ�ㅀi1V�G���"�x���{�6��74�����[�A�n)���c�`)(6���-[��#.�}����p���ɒM����AS������:��>zA
'Fi�/?穾|J�iYYT���	y�m]B������/Mig�7-$7�5l��$?�i��wh��C�V��JGob;��ʣ�[��ɝ��tĎ�C���ĝ�йԓ/,P9xaA�ZB�ʅ4fŠ3�01Y�5%����9�����c�������AU��y�lT�/d7�}
��ݱ!Ҷ	�jI(Z�䘎͛����kh�'$y�b��)m���B�1~C$��;ު,D�P�&���+�Au�{��m���S�
x� [t�1֨�QEFMtV�ď��| H�X�`��U�k�w���F@jĄA/A�l ��|�09�����ޯ<Cʳ�G�ڝ���M좣�Q�V�?�sg�o�Y�Xl�MA����~�]Q�#	��Ջ���Q�0N
.a#y����&˚�D�c�;e{��{-noY$3%�����X�C�%��*�v\4D�.ֻ^�c7e�6!l�>1��vMY���;9O����h����Ƒ��P	Z0��$�,�̋A>��Gr�fv��Wl��,�# ?v���l����]�y�.W<=h�.�(@O)�n���e��Gq��꺩6
�V1�c�K^�������6/V�5؋N�Sq������`�� m�D� ˜g�=������
���̓�}�1L�pS6����z����/� F#0�H��`#�7g�m9�R�#��%P��Ԑ��/_�ﺣqR�����C�A;�Ś�����4;K�y�G�]�ۭ�p�:=�qonG,Y��"06�/㵣�y�r���_�/B�//R������Qo��1%�N=}+Z�G���j�˗�Xk��y��=m}�s���ܱ��+�nH�ly9?Ԡ��p��jgkI[�,�Կ{Y-�pc^;d�(W�vF�-���e(����{��[��hm^W��9t�h"�i�q}l��'ܺ���p�l��iH���g
y�E	��s
H��.�������t�J�#�|��dίЖ2��X���	���$dMʰ~�x�%"��衝w��2ל߰�?1a���ԉ�[��;�"��f�`4r���/u���������,��$!���F��mx�i�Td����eJe�ua@%x�R��	lRu��H&|pt��ƙL�g�)��f�@\oF�aQȩRlf��c_�ڤ���`/ד�ͥ�>)����P�a�`���2i���'NV�FF��wMx�3�x<{|�����=J|��m�N����0�k��ug��f�s��sx���l-�� �(�e�#����	�)�t4�2�ȳY��K;1e)5���~��͂'3ړ���BH!�%ӯ()iʨ�b�y�'ZSO�3��{x�gNʖ�~H����T)NfJ5PGDMt�f��Ө,�L}����Qxh��h*�,�E-���A�Ǩ�P-,8F���D�~�J�����o�6[tp2V�py�tIvwh�ah�������ѡ���$X�޿���յ?�G�7.����z�@�XNc�(`��!��8Lq���.48_P",B#i�=�1�1��jz���/~��CC�y:Ff.8�|��z\���Cڢ@7����_�F*gF���|b�D��)�z'<�f�QW鉺3}[�g쯆����Ѩ���C�蒮=9����lQ�{Q�۠!�%�- �Rl/]uA��Q�ˍS\�hTh)�{��/h�p0�ApKo�T��mk�(��GSv�|�lv0�����Z�����${�h!�$s�et^f�95S��K"��ڨ�yQq�2�Jd��=v�]^�q���h�,l3�k�`.s�V�Fd�A�Kj
u?Q�U!/��;�@�ݗw����=���z�;k�1u��Q�R� �xg��cb�|�܄b7,�����bzѽ~��++�W�D�ʀ��fSw���-k�֖}�p�@ќ��3F�E���3xjq�D�%G�0����s; IA�G�*�*�ݐ0j	u����R��������Z��.fW%���g�'1u�)���7m����x��&p�8�sچQ��
y���lF�ϗ�ܘ	�-/I��>����O$�w`
�0Z,%l���}#!3Ra .��d'�Q��h�B_�`�����]�y�\ � �D9w`���^u���ɯz"��E���]�q�8�'�
}��7�2���A����OU1	f�|t������=v7�BŰD`G���V�Qq���,ְ\��L<N�2�:-u�]��`j��\�����8[F
���o�ڝт]���3u���G�@r��=ޜ��۾�4l,RSm�M�x���+�ѩ\�i�.�1��~�\��߄�_r��^PN�mă�G��E3��غ��ic#�-xd�������<[<�+й���L�u�es+����ؽ������S_2�E�/M��7N��ʏ5xd|�|��E	�ll�o��z�K
�
j#dT]����������*<mLm˹ܤ:+ǈ�1�3A�����@���bUdf��7�9��Yۘ9��$F��AEx�m$�?/TH1~Q�1&�-����r5��y��c���χSڂ�H�S��!�)�3��KV.�5��f%�]���#Fm�qMS5B��A���!Y���~���O����[��Ƃ�����  ܔ�b԰�����cd���j�]�
\Z ��Z ��l��qjvzULB���$���9_;���;�������ٚ�mi�G�vp�N�]�	p�WK�dP���iJ�>�6�u �`�V�aZԱ��;�]��j}�՜�aD,vO���1����:(��1�c\T�>���Uz�Q��따�$�:.�k�9μSE�Ӏ�i��àJ9�^FuŏŬ;Y�41���C�����!�ͶThH7����	b������)�h���1�Ep�,�*��5�ƀ�	����J��V�XE��y���|n)ų��/.qc�R�W�mH�kV3Xo�	�Y�[�A��mغ��O�{.�[�p�BO�l`~XJ��Z�u�;����-�+.� �V����M
�n"R�P�>�ذ����f̌�ذ�
���ȹ��E6y�w�i�1T����Y]���t~&���+Ŕ�)�*�-����v�H���+�||��ԏEv��y]G3y���B���� �`�{ ��  V-xJ��	�7x� ��!�Lx�q�[=��*nڳG6�'K��w��Q��7TO�
����wG��g�����?��9��f��D`SO��,�"}�O�0�괜vb�t�X^}���d��Xb�z���<�+ҋq�J;�5b9e	�d��P���J�PdD��J6���;����!��#��K�4qˤ�l!��m6��.�x�@�!���S7������t�޺&n�١��8O���Y��[�9�bM���G�[�%����@�p-��Ç�ɪ�:���c!՛$:��4���JQ� WE��^���uF7/?���w��dA_����T��t�}�㗳2 �L���@�Iݦ�34JAs)��_r`#�xxɀ�3�Iw�og$�VFq�{`���q���k&��G��萍~>���U\�%�$�攚{��w���i�DDs�]˥ݹBb�er��ݜ�<���(�$�LU�V��k�G��v�<ˬ/�S����*�7��
@�@6��|��/?kY9��2/
;��-�"xjW�v-Pѐ��Ae��Pɽ�#�x�z �}���^�c�NSU���M"�QQv@q;��ߎ���������22��n�;o��1��ô�5o��G:=��0-Y�[E��7G?�-b�d�E�����["���>��S�Nń�-E�� �j6�~�-�t+[�qM�sc(n�C����}cXӶx�h�D���Eo:F���c`���G�a�a���~FH��V������u� �t3�Dֱk������'d.pڕzF�[�	���S�{��Cr>�6hV��+Z�T(z$%<�35�����R�˽�r�S��Nɠ���n�VۗP]ږK�o�K2�'�+7 �g'0gƴ�"{�҄��1�o"�J�YF�GC>9���I�~�p���Vu��1�������~����>�tD�q��/A������bD6<Ev�ɃK�Y���MR39Js�E֭H���	��_��5 �v����k,Tc��^X��g������ş
��܀o�F�[�c����5,�W���M��H�z5�n �i��XM�^Q�x�nV�Q#�8B��E����/�a�ՐT���}���uf@?)r�7A֛�s����!�� җ�V�B��H�jB��TDX8�@��'������ͷ����I���Ej?|G�<�R��X���J�-ﱶ���I0(=�⒰�˵�4B��~)���-]��?���:����8��tp�����=���_�L�S������/�b����0U�1d5tH�5y���9��+'%W��nn^u��j��8���ιV@�[���D��p���O�q��81O���t6�͢�Eye惂����$)��=N<5y�`�!C���QI�V��J9- :7��sv��>�W�jN4�& ��i?I1����ۍ�QcM����k?6�+ǟ���(>��iQ��bK�M�e���%����UX�f_�L�s�s-�h��X�����C%�䝄�e�c��=u��H�<�IDo�͌}��U��:�7� ��%~籌�H -�}�ծi3�J�m���`l{U�#?:o��6��wn'M�`!�49B��W���C�a�ZtN��C���wB�"��?v���
�7�U��Pdk|ҍ_Q�oe@:H/���z��+�y�%��ttD����(H':Ƹx���:���� ��vu�(��'�L�E���X'�E��MOXQ+3��5�Iݨn�Y�Xj%$ډe�3�)����EO���Z;9��hJ�c��[�
�6u��P@u��_1��_����X�C�`_�Y�j������lх&5�{@�f�n�ٜ�uj��:�%﷊u8�>�R���\��Ip+HǾ���P�{g-q��磻\s�9�N��$��5�����m����'Y�kb���FIz7������H3�4�"�o�_м�{ϟ�_�jp�>/v�^͕��2�O���tϷ�jƊ*Y@����	�#*ՔP�`�¦jY
w��AtB��Pru �+���t<�� 2�RX����y�N̄�*��m�W����ʨb��5u���򹧁�q��Rk��G���VNT���/b''Ф-���ߏ0,%���6�`���c�ǃ��M�S�".@]�׊/naD��r��yvݿ��ѓ�� �Z��Y�9S5.,I�!�"�ʤ��UT��9ㅘ��>tC��a�τ#X��~U1�3ŉ���DBGP5�7�p�,�\f_BF�����g�vH�p�O��gLC�=�\�lm�$߂��jn�咶��/gi����.c�}�
�����`�Se	n<�{"���A�cC3�I��Ԑ�9Y�xSH�.�S/Q��rM���%�bB�揵&�I�<z�~ܘ�{�-!�؏Z��r�%�Æ*�{��dJ�+���U�h�,�i%!y5�	'#�߿��ξ[U?��������`�@l�E��"1��6�B/�F����-f���u�橋{2� ����F��ˬ���(j������N>||ň��;����f�C�� ��_�$&�<!��OY�Q��+]�0vO�� ��R)j�N��
�~�~�g���@ZGzq[�,�dtR�x}���%�����5t��%�J�Rz��|�5�n��� 0�E�Ğ�ç=UR�uz���#"&`���������(X�]�x����Ɇ���UI�C�h��T�ڈ�y rq��퀺��������Y��Ϻ1~�k��|.U��� K��(����x"������"9�2��G'��ۙG��n�},�|��~D��E#<HT�������P�-���H0�Z�d�f-II�Ӣ�_�g"�l��{Ӏ���䑖��еoD�+K�1�	S��Ozӫ]����+}�{=M"��ٶ��̯˩�(��7 e���։�x�Y*�q0.F�f�
%L��#�{Cb�'�������[�RM�@�.-2�q�:DQ�mxjD�q�)�.���׼��=���𑺦l��@������+{�L��î�@ހ�ⷅh3m�"��<�ٌw9���-?}����{
v�"��V^o&A��A�'�T�3sS���|T�W��rh����r.��4��|La=�o�g61�(Y���
zZ�Vw2�����W����~r5K�:g������Vyx���"�0z��iP��K���O��6�;���ө|��Ɲ�����	�]A�yl���:���� �f�PZb�K���j�rӮ�0���apz�����%�p�H�ǯP�/>��,	0�M�w&�bzU;�C�j�=eRЄ*O,JϝL3��	5���oG��0�vq�����,���̚Q�J�G�sA�r&&�}D�����w��A�l&�{������W�ӂ�(Kϼ�E���K4w^�~�_OTd��O�eR�1�l�Htq�,��p� ��fr��T�Mu2��T�ٽ_�2��i�+�8Q�"�J_�̖;�M���X�Lu+��½��='þi>�i��
���.v��]كB�h��Ik��DDs:��0��h��4���R!	�ua\~gf)>l�K����6G���p2U�k&^b�j�_�Co#�R�����Ԩ+�2�bc����@�rp���W�i*��m	�Zߖ�<m�F���=�,�* ���Ŋ��nK7�%#�Z/&q/ی-��:�
�[����÷M�N.E�sӆ���NoGj����8��n�oϟ1i��G�� |-�N��h�6�u��|	�f��1�9�����91�wV%U	�X�nhk�[ݖ2-��&.�3d�ȋ�[�#�=s���8�O��y ��:ěJm4䓘U�L}xl��#�gn����&r~N�@�S��|W�W? ��?���v�ɿiܨ��Y�u!�ʭ��
���Q��>CT���fzU��M��/��u�vT1��l$񋩒y��}���xa.�~.(�5D�"H��v�x�CuS�M�t��N���5] ���� �Zc���$��#���e�q8�9�!%|t,Jt�4��5\N�̭&�=��S�z�*��Sh���Pz~=U8�2�e}��o���(V��$�v�9R} >[����o8(�[˰��w׊��1 S6-F�� �j����k��70(�g3����r�TN�O�l5�Rl\���}L���}��+렰�W5�Ԕޡ�i ����^3��-ʢ���`��6���	���N�K�c�..����D��o����;���=��A�v��A��3��U��A#,�_p��	6^-l%�Pu�Q����L����+۬���{!U�MV��y��a�L4�������,�}eS6��Ӣ+#�?����$�����&.��_�?/����a�r��G1���N��6���Ōm'�>�a|T��}M���G���Y��T�FN�G�4��קc~�~�����y�^<v��xӻ��Kr*�ʼ��W���m��Ȟ�~e��R�iS%֮�kZ^j���v8{}�-�Aj��T�q� ��d��u�1�<	u��/�2.�ĈN7l��]��������,m�����S���E/�e'�vغ�>s��r����V�q��])�?������^��%�Q�Xj���k��;j�TT�|��^i�o��6a�38�҆?^.TPX��M�-��ùy� J@Ue�44kx��-��Dt�v��e�����f���A3g����KS������9T@�B�_�z�̈́�6�!�S,d�����3V6
˙}9V3�(Xw(�_���qh!S��`%������},`�u�X�Bi�40�:�+v8���p!�4�S��5�x@�1��2��`�o��'��/+���O��-�iH�v]�F�o5�G6�k��/ω�b�߳��Pj12NdB<I�����p+c�[�Q�}�YUh/dYM�v����k��i��cx�I"�K9��.���a҉�SA���� �;-����g����M���Һf�e�=Wt��@.�����������T�@��-��EI��c_��^��.EO��8���z@�*�#�W�6-�9��GO���ޠtD�7��KM�"O�ND��l���J�H_��s��UX�`�`�N��5S��w�R��BON4��ϝ�UJ�H��hS���S� ������npQ��j����u��Oi���O5���E�<^��'aEW�/��R�+�XI�Sh�����/����C��^�#�[H�D^�->M�D��FԅΒ|b�MU��w��$5����k���+_c�g�Ĳ��@�7t	�gG�I{*ڗ^;i��]�L(-������Tnwc��7>I���l��}�Iú��E6&+�g��C!Y�9MKw ��ݫ:�&�K�ӳ͢}S�b]�B��
�"�._\��-��E��◞7-��{����_l����� �hK�W�.����T[؟�?�~���"l�\`+����N��*���UՐ3��Q�6��bka�&mpk�%�ǁ5N�.���V�*?�Z��i����<�+���+��E!�.��M6�.<fq<�.wU�+�S�����R���椦�u�F�h�f��i���N"]S��0�4�x�^
��{�M�f�+<�z)rd��X�O0��tԅ+!l��
��<�j	�s�����-�u�w�n����K�3�{��@�o��O��U�V5����Iv��御�I��(�F[dKL��˧)�R���əTd�p
�'��	@�vP��(��[7hֽ7��~v� F�x6�����D�[�}l�挎7�I�jͺF�q����Sd6Nl���T]Y܈f�Də��u��{����[������	�b�d��25�7骖�:P)�r�%�#p�U<3�U0�W��ч-�y"���hty��;*��H�t���K��P_=!����ҝ^p�
�&�ЙF�\�l���Ӌ�_(waދ+ښG�{n�}۽�BxX�^�QqBo���@�Qs�/k�n�{�>��jc������G�m�"
E�gm�K�e����C��J��͒�~T��[���d���۵�к�j�L��o�
֓q�&�:��� a�[�`2l���X�G�@�l���c�c$���_Ħ
�%�tO�����F��%R��u`D��Yuߘ#�}�(0�lYX���J�0�#���
k'<z��c��;��3�#�\��-�	I%�ۼ'F)�yKY&ɂd^e��=�M�������,���4�.�v�Z�B	ܖ�,=v�sQ������e�2#ɣ<R�բ�Ч�E���;A>6������nxo�z0�(<i�X�C}��q
&9h��A��UKc�t��xz���U�3���G19η ��MՌB!��D���K��+ zLF��,��V$�����1��~����e���j�|�3c|�J����\��7+L��ƽ[z�9�5-�X��#��yx,b�z��^��?��߁>$m�;
��W�C�(�J�� �E>�d�~���
��l
9������>Cn�;'N�%P�g\����?�B��k��?~���[���=�H擺��Ÿ�����%h(4���TM�-���9b��-'��KƔ��-f �]�)�Zh�L}I��i\�۪�.�/��Uow\�}4���F��E���c���+9�cL�̬�������QM�K�����	��c��?{�� ř�q}���u���}H���Ass�wv/m�&
X�`4��Q����x�P�	m�i��M�R���}\f�����i/i�K���3,���83D�it��nN^���
9�����sb_Q���/��)Ё�o@����Z.d{{���#�+s��e��Х�����2�mK��7��dj�I�=,�C��3�V�l8�!�jga�Kb7��qлQ�ƏH`g=�2,�(h��0���_��I�&��.''\n�P�m�L[n�T/V�7��	�	�N������70���g��f1cû���z����۪ͭ�Z��,�����x�H�Z������/����� M�'z(UY����[0ωG���R��j���d��5'�JhD��b����i�?����S&�3m�	m�u�z�]KԿv&�/<1$�=%�����HB"���`�	�B8��:|�`����#�RV������`$�����/�:�}m���p.�' �ae�=������Æ�Ƕ3\����<�����D�]sОU7)�$��g�/}D��`��e�1o3�}o�gph[H�&��m���ß�&ϙoJ
���[+#�Y^!$K����w��� m�8
���T�r�F����Z�3�]S4HcB�F��R�"D�O@��fQr5	a��Dժ�������KU>�t��Sm�G9@�lW�wM�� ��z��	zh�F��^^�O
pak�ɻ�g��nF���ᯓږ��%�����1Q�� Z����E�Ǵْ;�by�/��&�ٴcg-+em�ޢ=�l��4�����Ӕ(����8.��L��y�� z26��l׶��<�������IA�E��I[�}�A]Q#�/�b��,��l�:�4�hkpv΍�uc�Q ye��F�Q��?�R?����a�ҝ�Gq<Y��0+�C!ܱ%�
�u�#σH��.�4��1���ƞ75�����d�I�&����Q"�1��k�Y��/�ŕ��ۚP�o��2�������E�Wo}����P˩Ȝ��ΐ{OaႾq8�%�y��l
�h
<N���{����Z�r�'�H�	w�8��(:�E��5���fb�`P�Xz��7uMF2�5wؕ��*t�N{t����sŕ>��{�
X��1���+��l�c�X`����F�l�Ͳ�r
CZPoz�YEs2Ԯ����nn/<�~���!�\���=�޶�b�Nha�S�D^����/j.:���`�����fA���I/a��J�9��Ȃ�R*�_�����e�@��n�j�,la��t���ŧ-? ��"3|w�g&K�[��,�q%�敗��{y���:�1����sss����9Ѐ�<8>Y0�\����J#_�������%ơ!fTM�G���!e�]��?@��P <2Z�p;�6��n�~-�.�Ч�GHU[8m;}�r�-R�t��)4x��*�����Y���9�� 糪��j�L�FVb@~���<Hz�;E�r�������D����������QI]J]�����l%������Wt;��3a�~IX9�R3�>�v�*�t���ӛ��̛�Ix���D���'Q�/����:��A�G�Q��=��J�36�,��fo�k�C�.D\T+�3�6��D���(���#��)W%��I`F衂1���s��I�(����Q$}#��̨�k��|��a{�D+gC���H��b�?砸�'\��-��mG�)$��&�'+P���L����qk(����!�;�r��	�=W~S�vO|������W|E�/��GKn���Gc�6�#JY��h�uM�l4��g��ṃ��]����_��ϳZp,�����yl�xӼ_�vv%Wz�����R�~x^�n�TGD���Q����2.�Ek<ԧ�Sp�E�9�1-�CB	���#y��+�g�ga�r�G��1A�K��3W�M��zo2� ����� ΋�VJ��h)�^�@JS[�m_���?͓���%Iȝ�bp�&n��L;	}6=E�z�:��0�<�ک�{ν1r8ho0�YQ�Ph"��l7�#�ǣ� �?.��f��;��L��f��f�S�EO����ɏHІ!"��m}2�2d�rY�u����ؽD�Fi[���������h��(��5�C L�������9olax��e��x��TR�[c�����.�-�Z1��R�X�"��O�\�ρ�����σ3�|v�ݬ�Ue�>}�!��G>Fwy��:�^`�˕Mٌ�M&�n����ø4"�
ˏp ��j���i�����������0޽�4�1|l�  �f���v� ����"4����w��$n�J���-��{���6b�g�Vm�D��X,uE�Q��:+����8��|���+�2Q�4 U��/�&����?6�Ƃ�y��Fv
�.����3�ě��@����~��l3T͝w7<��E�`I�⋨���p,_e�$�@�,F=��X��4j߁�U�yE�|쪸��3Aqk�+_�C��[x!рϑ`����S�P$CT3�u����{1sv�L+N�8��a�)����O]9�C�)���I_�M��r:�h���*���7�DɎ���O\	���k>�p��;�J� c��-_}�5<A�����^�q�Ǒ&�k����|r'��b���oJ�zI�X�ye���{՟J�|rBP�l��^d��u��=pƌJ .κ�ƥԤ]0�$�E�N�@5�����/p��C3&;2�fK��W���V�o�m�&�/�Q�e�.7n����^�)�M+5��~�TU��eF<��iS���o�}m���Ё�f|Wer9ˏ꾐������u��]�����0'��a2��ؔH���Ϸ�)sk�X6��("��}	�8I&�Q~^Q�:e#�9けi�9�U)�0XZ��h�ܺ���og=�)*Y5 rkw��]��|-\�*I~-3U�<�Dl�v��}�=��B~ň!�Kf�m�4�(p���~�<��>��&�=�v<@��3��se�w͠��Y�s�!��)�K3��R��n�*7ɬ�rK���|]��T��X��J0��5�h��eT�����ȝy,�x�	G��2�u��HI�G
�9�^����2��I����C�0��-kʊ:k���|*��wq;�Qąy
�+�[�Ɲ%�D��Ḵ�Ҕ����l�*��B}����Π�"���^�8��Q2���j�?�6-癿SPᅷ0�6���.r˾����9�m���`@�1ڍv���'��G�|�� ��Mm�����&��#Xց��̎�ɝ�>40Dӧ	D����sA�SM2=>��RW@<s�k.󜻹���0>H^^�'M���b]�!�QH�, z��g|��N�U,}��R�.���@��2B='r�±)�nP@���t�d7���m��Ay��"/�j�P�zڔ������=�Z%�|��%�{H7!�w��N����Lw���n��P����(�^F��]�Q2�&�Ϡl@�q_сGq���s�082�U���
	���/�O��<�4�
��Z��	{��j<�#����j�g�.��"�3��ׇ�s��x�8�@s�ʹ��҆�ZP�c.�`a_�B�B>?e25Yg*��6�%C�������j�ph����G	y>P����>VJ�3�F�[]P*ps_G�WI�5ݝ�A�!����+n�O �I0�����Z����ؑn��Q��x��Q����Ȏ�S����p�K�� ��髚��3����Y(SG�`�P�Ϫ�=RD� ��O�l �����,cm�����`�e ws%#�BO�v�[$*GBi0d݁����݃�uć^��	�����]�ѧ�?⫐�FK%%8%��Eu^+C4l�=�&nNbKlnS�Lk5���3)۱�?._ũ���*�g,�JIHa/������bM%&ˠW5;J:o僕�^�~�R�m��>�ͺ�{X�"�Z�l�����3�}��2���a��k��UW
*a��?.:,|��L�@>�q�k&B����A��f�B�I!���4����-@7r�!5�=&nf�`�(�/��݊����M����!�L���K@jCr!1�u?|<nZ�����2N�x�N������$�����;�pX� J2A��=V��QH�Ț�ᬻ���4����L|6W�hT"����.p�Il��;�n�� �Z���"����e���>�`�����qvb��;RRj-����~W�ؑ/��@���
��D\��yĔ���w��pZ@g�ܺN�gV�߈�L��>���FB�B�a�ņT�C��n��i�o�C��y�2��~���?��ͭVa% @�a�p����U0n�g5��ko?�� q�c%7zP���	:<�X?,�=f"c����Fug�8�#�Aj*�EKFW\����2���DH�*��س[�X�_褦'[C��>MpB��z�"����,53�?%i�>��: �3������Vю�ni�l�9m�c���M��.�~]d��Z_��焆����q'$�QH�����U�B�U@!��y�׈y�2B��
�A^���A���΄�,̆2�gg8�(��}��X,�ˠN�=�E.m�1�T��W��ؑ�����y�`�l�`�Jwݔ�W�
�P�'��������C��Åu�H�c}\�FLH*PdWCb��-ׅ���dM�m�/�K�	�k��L�d�e��Z�2�6�1zխ����q��l��oO��=jj�fK;�."g,8��в:������W���2�ϣ�y��T�	�����r��1�N�[R����cLe�1���B�wx�����4��j�,A�e�	�Y����ZdNE�T��c=����6��f��`���L� �(D��*4r���^�����X؛d�e����[IZ̙n4/đ�`ů1Z� `��e��a�(K�XWD�dH%A��g�S�C��5j��? �m�QI/�mv-ߙ�F�NUfD����]��M���E��b�@{�\aGj�鈽��5��8�_}'�2c�_�� �ȝ��|p=rV�Ow��eD�	R5�)3����N�!��[������CuC��O���#�ڊ��:�=u����~"�g��d�گ�onDu���=��T��E��%z�2D*��Q�ih���e��nw��z�(��P��٩��~�ߙ������=$�c4rZ�k~�@͉
3����+4�|Xp^���*9���ZI�����^��˂ ,�k�^�b�T�7Pn;k�3*J�.Wܮ��#r����m�Hj�Q�TB�����wQ�C��]C�7�~B�h&��V�y�[=Ea�R2�aՂ�7�c����4���;0��ǿm��,�SEc���5����2UQJ�A;����(�]f�K"x+�K�?>���2��,�m�Q	�!Xh/���9�Z��W?�	�v�'_�
&s����:e�uބz`�zwM���J�[��?��G�&j�X����N��A*�~M�Q����;��3/�Bf�OEO�2����r�H�y���W�Oe���6K����h2�2�F���g�7+�J{�_�:'����2eYo�m���ڮ$����=�i&B�i����4�?̀b�}�v����v�,ԵW�27�X��v��*��ţ�4W�Z��&"��Ӊ�/�B���P����_ATc��:wЙ���?���
��̐�S�*��SQ���q��=!m�?��D�����n���[�C�js���f��ǃ�/������VH~�&��O�v]��v;�n3&��pA7�AW8���W/ <�x�F����$Q��,*4h������;�^w�b��`�/�I�@~�z���Ы��ĭ�:E8�7l����3I�D|�:K�Q#��>٨��
~�V���s�S(¯p�� �+&��P�^]�GAi�� d��R��8v��鄜����Z3����=1b �A��n�WFk
�JJ.�y��J)��^�|���+B�����ɲ�bͅ4@���jU1#��Ŝ�j���n������8��eg�5�Z�&�K({���*��]L�v4W�K&Q��������`=�����υ~�ɷ�j�B�q�}����w*���f�/�N�jj���t��E��E�f��T	5ٙq�F�u:����P��,�WB.��"Q�tR��2�`�R��ӵA��dy��ڏ�ۋ��QQ �MU�i�6z��i*��=<:M�`��ǒ��ݵ�{&�6�'��z��,�����4�f�#���|�!�/sy���sGT[����Y�"�<���6쁔��ѾaK6�pddj1~�D�ن����98̡X��B�-d���3�CoAe�`7�{X���Ŀ��3�ɔ���YfZ z`#��v��.C����5`�C^�q�8�b���)}�Ȧ���䭹�F�yT���d?�GG������	".�#7ߡ��� D��40/|?��M��|E��-'�x ���H�6�&���R1�P���B���A-���V;��d�~*S�9�A3�������@С�6+9�M3��x���i��� XW*#��co�|R[;i�"�Hǀ�T;�m/�A�,$@���+�|/�˂�6j_���E�R�l�1t�e��������_�[��4�ş3K�LIo��g�%ל�ݶ���4ى�?�:+ȔӰ�f��a���X���N3�5� *��rh9��g�Aom:hǀ �"al�&�(R��J���)�
�b$.�"��(���_�/���"�3��H�^�AJ"��H�$N����j��JLf'��7��!�M�Hr)Sȫb�ˇ�T����z�,5��Ǧ����G���́��AO�h��U�"��,@�<N,��D�s�z�TdS%�ZN��fG��9�Ŗ&� c�ؖ]j�w�8�.�G�;LE����p�[WZ�3d����s����k�:c��V�cݝ�I,�O��&E�"��'̡����v7��LE}�I����k��+�=� ��>fj�]�	�Jy@	�~8H ��T��� ��x�P�u$d�&��vyX/�@��۱�C�x�I���G��"��5�\|��{��\�`�5��(��h� "�Y��?�h�R��\���V��&ձ���������X�S]�� �~^$��.��=Ё�/��^O�a	���Of)L��v��ϑ� oڀ��Wy�,�*��1�fs�H='-1���k���]��x�ֱ� �ل�f�J�j�_�N-ю��b�����/v����zN�iS-{���U�g^����Y]�פ���QY��F��ǆ��P��Z�X��F9�UB�F���Y��%���>�����P��x�����$���df5N�;{@Й9D",�/�r��z]]�����L��S`cn�B7}�O�f�(
�M�>�3�DU��<ѾE��ra����]�p���-<�$XZ�)�>���B7@��%N�-�I�)��g8�zx��KN��_6
�o��a`5�+�PX��H��ւ7���i��������83����b_�u���W#�_t�Ax���O�6{�� �8/$�j������3$,L���x�������iͤ��xEZQ������2���f�x��ZD�ڸ���7]�ս�P��7�����~�t� KEݱ��.�s;�QՀ������ߣ�
�2�te	C�W}M١�=����B���27J�rX��6����!���l��'�6j�M^TYU���5�X'E
D�t�n���q-u'V�����4{����x���L<�N���5�W?��׸��3���4Dk6�T�oy��%Y`;z��C��)\�+�su�C2��h�BI;d�*�b�� ���p�Y�Gۆ�!�����	�T�0u 
 ��nf����?�j'��Ǖϭ�OT	�#F,��KhCG���z�*I�K�ǅ�HZ>���.�����6�?�#�i�{o�1e.����Eߎxh�9��&�=RI}
:���:;�i�.+[���T%���a�&^� &*�M|��=˰*�{bp)�򢊢}����aC�Kl��c�7�NYu�u�o}yC}eW�r�q����Q��vW$<(�`ړڽ Z�ʷ���C,b�Ō�*���̶�z���D!�����5��~�K˭�9<v�Ф0ݳG��=�j�GW�"	��.�.R�H;��o�}F��XJC��~OY'��Ѧ�҂��T�2�gwC�H�B�X�s������ �L?z�K���eM�M��^��Sg.h����J��MƱ� ��ۗ>��j_�j��n�T�G��RU�1����-�u�Ǫ�,,�v�D�q�N�Xhȝ�R�=q�,:�1��b���(�������?��% $�V!�r 	�ZUa`��;�IeY�[�M��{1	~��δ ��!�cS�����D��O���m��S�o����77|pw�0wT����]L����8�G��V�rnpL'b��W	��Ȩ�d�|��S��$#L��`���z��q�#V`������ƕ �jb�U3���>;7�= ^�4�fB�sf��5e���}p�h.t9�F�A%Ǭ.C��@�7�u���O�k��DCM
d�'��+Ju�*��;�����:qr�9S%�0>G�b�"�>��֨? v����t�t�=�}�͗璪�t,�`J+�����;�BQ�:��@/�4����5\zdx��#�;ʿ5������>9�0a��-��;d�����B�`��~G	'��J�j��e�b�r�{���_����Q�h{vX�B�v̏�U]?:�*��%v�����H�|);��(ٖϤf�m��̜���ŃΨ�t~&�~?�p�V���`]�E�J�	����G�L�nD{�O��MCf�(��zR��͎>��	]��fg4g&�[#Ȋ�
��0`�n�j�Ǧ��5�|����|����(?�����{�Oh|,�ygV�1������I*�>��b�����y(��? V�D��CY[[U��`�k��R\��e��b���6(���U���J�h�'#��C4WCY�p�)N�t����k�-�Y�� �!hz��R���\iC�4�[�n��>��������YƗg�n'q��!t��[��� ��8ɃԄfJ�S��A૱�ˣ8��c�P=���� ��N��т��1a t����d�3�1���QF0�ArbM:��:�ݼ��l��t���쨝��\{��.�=�4��Xi����N�r�0��-�X��	7C��9�sD�G�b������X�:;�*GF4P��7`g�?���\���YK6����DY�'�U�צ.>�B*:������ڈ�\"ه�NVϵ?ꄦQ	�L��C��(.�t��\��#X�LDQ��P���ת<�A@.2 
��uJv�F"zc�+E��יuQ��Q��&��v�Cd��A��y�����kQd�C�@R�"�<�3��1YX%P����V#�@}��C3l��З�p~7�x� ���/_����е�Ē(�d�,�>���w�SZ=�^O��;7�4�IH�8���&9W9\e�9�Ĝ|9��a��C�F���gR�K`qV׾	:QY[���f���"y��9| �/U^-6���bxpV{Ac3&�&����H	S��no�H����̛*y�R�rE���%
�T-7H���p|�O���������z�"�%dd8f��,�z�S�9���.�ŜK��#�A���^Joj����r ��Ţǻ�d�r7��>~�g�,X�ޑ�<ܟ a���0s��ꩦ��In�$e�ݛh��d�G���c�H�/A�����׵������
�����]v�5������e�ϻ�Q�":$7���G v�,عM��-��^�6Se�d�n'I����c�(�u�"B����`��v���k�� ���Ѭ����gHs`t/�����
��%C24�����ϴڿ���́��U��#ۮ�څN\x>�8�Fė�V\���M㧌��-�t�G��t̴�И*,��\<�g4��c�U���\�wBG0���6����8�ܸ\W�e	�+����Y R�x�(q4��;���xZ�@!�(m�`4ؽ�ET��蜺��!�L���?�Ss��'7��C�*�q����V#�dRp���rsk6�g����u�"���l�SЉ]�U���]�)�<�Lv������M'�Wr�cҐ�P2������v� 8��CwK�F����W�r�q�̿{T�?����vqE{j�¸51V>�Hm��n�����&z����E�<���D��4ڝA�9�zjV�x�:j��s
nj���Ȅ�q4�z��9+�m��ۊ@���zF�T3v��Q��T�"e�&�P����{Kev�_�a�$���3@kpO����G*,� �8���[3Oq��+�M�FТtU��0q�c?��9j�ʾ(�K{��{f�,�P�댵H���oN�}���D��GOE��0m��䧧�`A��K���n��[�J�ds^��\�'`>\��$������Rx��fLo��;$�A�����,���,�ڢSR�1�H�5T��j��p��`�vaQ���<���B�buWs'�Yo�zB�? {p�k�,6�2�0����j���c�i�C.-�3=$�BڅJB�����l��r��-��� ��Q}w���E���@��6�Q?�.�%(�C�~Eb��s���w����mK��'�frԩ�u��<,̆��U�G�2�|l�p�k@K�[�)���Pk�{��#4��<ϻ�H0�j�J>a�K�W�^Q^����W������0l���Ϳ��U�B��<oZO
H��T�����	��@O���%wx��\���NQ�b�_�O1�۶.d��J��8�KM}��x����xt������]�7�]4�hli��DLF���E��_Os���^���iÅګ���q�T�Phb���<:I�w���g6�i�R!��a�~�3h�x"Iv���NY�D��v�4-�;�V<�}_t�=�������c�������ю5L;�Z�v^Z*��w���r�M��+k�KP��\�iU�:�G�}Ð�dm�̚Q:lA�����U${���-u(&w	���@�2P�<t����u�����(�(�s)����@V�b�T��!}d�}K��#W܆yz�������AD6ZUkśԋ��FdU�_�/mb��������{��P#�W��@I[oxO�)p�m��M�%����D�{eB�=Fhz&Ŝ�� էt�W���<n� ��}��U�^a��"jK���5��lQ��̑X��⎬��Ӏ,"*�9%���^�mPD�t6�u��l�c�fm.t.���ǡ܎��66����i�F85`g�����q>�/�	�9���5�n�ՌV3!Y���61f���ȓw�����fz����R�۰�^V����nS�*�ΦxxV�$<ꅇ��u\���Z*�Ɍ-�ke����	I�7�O��r�����K(�!Fd�N�K3��IUn}��d
���K�@����h9�w���O�]��|9l�ZxqMS�|���d��-$�.l�` ��ؚ^���2+�X�,NJDU���-��_�kb��! [��E�{��q��B4|o�R��,�WskW���c�Lg���a��N�/�k����\84^?�*��J+�����9��/v'�8*u�� .� {�,�汷�|%�O[��5x�K���2���iG�@�m��.��Nl�t��RM�w�a���1,���'%q��e��Ý9ة�\���L����.�Fdc�*�WU}��e"��216��Ϧ�ouW_CaV+t	�sAb=H#��=����S�JN�"�_-��	��OPI���>������^�>Y�#O��)�W&Z���EH(t��N�\%�6����<�L�6�L`ށ�$9��]'Ez~(�e�#iLi��K�s.�����/d t�����3�P<֬Ei�ߺ���m�"��<�0��k;g�G@��1nʻ�k/@O�^	�%�����W�����w�YHˁi�?p��Gv�5���V���+�YX�<-�������uob�������[�"<v�D.Xx���;�)�H���(�c(M��v�C�����	>L�=�����S*��_���w��y�
 7}+����<� ���z�lC�k��k���r�Ϲ>�=�50��B���=��r�>1r}OcDfؚ�/���+�р�b�6�tV���,���s���$��U5x>��
���iKJ$�5�.�KoXR1�w|�D=�y�T��y�����5������9j�M�x���n��y������O�t�,JӼ�e:��[�C�����q����+P��'=�b�����(3xBS�nݤ9F)7؝�FA���#,�6��8f'��T��Dð2�$���S��^;Z<>�E��av
u<}�������^�(���?lO〾���b�jډ̘Q�X�ŕi����5	�b:�L�"�n^��sX.���i.(ѳ���oo�B�k����)��J��!o�3-�$���ak��Ca�u��qP~+�~yqdC6/��������d�Bm$��U^��"�Y#���J`�F�HRМ�%!����J�ܶh�I���GrN��,`�����'�q��XpRcg�҇� 4@�~����O��T������iE�P�rڰ�r)dpv~E�5��a�'	�{;��.��K���7P�\P�4�5�������Ӓ*tL���
o�\g�N��/*�������	p�9�H\!���<��@��5�O��P��s��T�ҀN��A�*6Cme�>��Ř�EU�g1)�����*Z�wЂC:�*p�O�������\�դi !��������N9
�P]�`����� k�r��h���5��za���P��.=<�{��U��4�kHH�ý��������XJ�Ӫ%�qJ0>�V�g��oK8����fq	(X���0���0P0���tA����A|bn��u6��D�A�&7�q�7w��l	m���$�G�X�fMmܯ�R;��Y�2>r��~x2=� y�I�)�����v��Ŕ"K�F��G m)u[#�ft�L�Sg�}��.��ԗ�(�DU�ܧ`���V#� ���b����̉�z�<��0=��W��z!�@�#K�����9��XJfh�(�>c@+��hJ��'��;���\��(z����'R��0���69�=��a���XN�O�;�~��� >��|��$eHJ�hd�lY9����ڒ�GcL�a.�x�/�� ��>��-�!�������ߚ�C4X���`V�����G�ku��3��]�wI�$�.7��
-{�6"+9X#A���/���]�����,����R���/VvT.O+��]�����E��l��>���y�G�Ĥ���]�'3�J>a��]i���v9&�����Jm�)�v7�5��9r~o���������]S�\q\v$%[���S.uh:!.-���%eD ��!J8RnŅP��p$gȚ*(W�� Θk��#qI{�{Ə�O�*����n�CDr!{/%�lʀ�8���ĂC<��A��"�U�UQq�q3r�`��;�<����xC&�l}�=�8]���V��ȯ6-DVu��&1��SH��ۄt�e�;i����F�	(E�xL`��T��s]=�Ļ@���$Sj}�{W�!���nhc��пl:�5y}:�$�r�a6��BUT�Us�Θ k��.,�w,Հ�Dۇ�<am��������4������X"z��8���z��i8�!W�B��D�p�J\�X�o�h��גYpҼn$�;�:��g:�-R�=]��S(5y_�W��-.80��	2ȸ��
FКu�O��跗H\�[)�K�&"��7��s���>��a����Vu�Ky��=u��������gC���!����B�of�Yf�Ψ��3RS-���/d��C��K<���l�Wu��@���R)f�Q��i�;�h�	3��V]���_Ku�/?�>+,S+ ��~�|�4�݈������JR9��@� ��K}�9�d9t�I3��Hnm�ъ�^`�}��/Q�&��N�Zl]HO��U��W
#�������A��b�;�=���<̕e�ڏ9m.��E\�� _�d)re{���%�.�|�p"�^d.�G`����<�#��=�+0������c�W�����Pm-����n.��%y���0停�Et�%���;��i��y�����f�d5���r�^l�=��Õ(�m΋|?�͔�<��`���g-�[�9iU���?s�s��Yq��\
��Ao-�ko��LzbB:�V�MC;"v�����(ۘ���z.�%	��J������wo���Z�!1���j_����+�Ӵv2H��Tآ�T�_7P���Q�rw���i%�q�Zl�S�ǘI�d�7#�Aho[�U��:�S\���,+`��=�f����,�H(��-BbHNv/���^��RQH�D�[M�Kٗ����Ij]i���}��	��X���EAІ��?��R�|1KAwc>��Wm��r���6�*��Y�Hq��
��>�,��=�%{�y���.�$3�;<�N��?ݰ ��ba�l��V1���h�A<>�D��4��n�]X�)~��R����7]� �{������ǹb@t�[&C�Z�E��~r��
��aN0P~d��̉'U�A�x7_�x\�/eW[ʷF��و3bԘ�i~��TZ׆#u3л��R�p��7&�J�_3��UuI�u*޷����}�{�3'�VS�/�+Y�N��,W&����X�O̪V�3B�?�I٬1�S�1�Õ�����n`J�R1C-�:��=�?�h^�%W�8ƣ�.ϵ���m�y��z�kA�㸳y�������XN�=��5����~`�?��l}W������Y��C]619!ģP�b��?F�M�r[E5�����_�P�b�`�nl`c&c��v1ǆ/#����䃟�p��)%�+��i��l�6�Ƞ�Vd�ks9�
�NÕ��z8��}f�n=
��E���` k��ܷ�I�?�2X~oYhG�����b�`�_�2��B8�������`=��2�[I��Ѧ�y����,��b�I�FM�}���E���T�H݅�4d@W�\���
�ԍ)���>J��<Q&��?Q��݋�]Hp考�RޠJH��_ɏ}�,�M�wxް������:�Z|�H^H5hqq����Z��� `E
�FY�O����:��� ��xp�`$�R���6�qU�)T����M�"hF��? U�V�D�P�om	�s)z&��?�0�Ý>uQ�z�}��KB���r�"��%ܥ��e�������ie��,U*z�����}��/ߢ��b7��`�h�o��"���9	]�� ���Ӻ��/��"?�I��"
^4�Φ^�=�yr����<�g�<�����O�i6����.�z��59@�E����E��I���ŕ��)Ļ��L��Q�BjT-����V��>Z�@^\��e�#~��%",���3����/%����(���RR�:#���rD[�c-E0fnb���d'kѲ�E<rE��k�_g͠$[��[|�س0!�����m;���%��oA �t����'j�N/�%�aZy��q����я�m��cR[4������|�'y�Ub[�=G1_7H�R��ص�ͼǑ$�K14i�8�GX?djvXe�N��!�)O�X� �����71��i���l� x<�.C?�*"�p!%�a��1�a!0�Jvª3u&'Q���J�a0�0�y@��sHT��qoغ_�*ڃy�mO���<iz
�����|��Y�W��� �O��ī=��=�񬌲c��ޙ�|c��8��$v0�Q�e�/5@�hp�=����ξ�%����;���BZ Z6�z����ۄ�5!<��V���`uo����~epv\~b�Ԟ�x�}*7h���e�u� �ы ���lɟj��}�Z�X�=`C}�B��N���}����J0��]i���N�:'D�G*p�2�_N���=	L��O�L
ƴ��`���kmp�W�3\M��\f_�+̬W#ϸm���1��z�Tbc�7�B�W�E^���Q�B���.JI.��[���rbn㾱�#���7��H�����#����F��B@��,Hg�
	�Z�Ɓ�q���89(8���m�j��[[O45F�<R����B�#����8N��b�b������Q"�:��(�S���	/��*tiZ�`��p�X�ʎ��l�x����h��ARA�I	@�xӧ`�����F�:�k�T��۷p�Ta��5$�"-��dk���A�Ơ�����Tʢ�֋I!� �B�f�iw�?Q��;��]�N�M5�p�:���a���7�}��n|�7X�P}�+�E�
��:��,	���\E��w��^S*7t(lv�{k�\S	���u��[$����Ɩl˫sSSz�XX��1�����CF��i�Z[$��� Z�<47'5<�j��q��i�I3�k�y���Xd�h����6��G`����%W�K���z9A3��!��� `�9g��/Tᨛ��bHp�������U ߂����M��B,$� H����J����e-�����+os�p~�JM��:�}�gj~i��mQ��s6�q�)h����m��L1Y��p�5��d������r��B� �w�q��ˮ�Z�V��pV���.����W Ʊ���|��	�tΛ?yP;���擔�.����4�ۂ�X|ܹ��%��1g}-�`(��������������׈����� �I�����[v\
B>*�L��M'[��>��T�Q�� p�5� ���~�v�#<���uyk JN��u��,Ir��`��*������(,�F]z:ɇ�]�K��[R�,V��&�����l��@�2��,
j��n\��D��8<"*�M*�SS&�|�u0��~z���e�(�L�}�J,��P�j�LD>K��^B��gi�RcC%Z%`��֏p�>2�q��+Me�P5�ۙ#l�'4�����f�����Sc
Ă�E�Բ�w�L/Z_��+덛i����eR7c�����R�˂��y��0>��8��	Ȃ�u(2|�Kay�p�oJco���R�n�����<�j��xi�[4�e&o4�Q3D���x>a���CՂH�` ^�f���d�"裘3ʚ/��r}X���a��vRuN���:��D��.��`W}��p	�*���9Na��C�e���m>�ot!��;T2l��[&��ק.�S"��{H:֣�����!���5��y.;���Y��\F欭�WON�Y"=>z�Ik������>�:e�}�e���Ժ�6�5��McT�jOH�Q��H��f�MiI�6
4��C�M��F�^a}���c���9�Z4�̙�O��|2���7��[��ՈI?�g<>�"�B�90�N���\���͔V�5!�� ��GW���5��;0�
WS~&�v�W���T)�0�4�8բ��3ѫ��R�s�[ry׍HO`��
�K3����j�v�+�d�"<�2�#��S�W5��f֯��޺�
��w�}�� �=M3mY�,Q�g�A����1V�䍺�4� ��˕�PF���ɩ����x�qO��J�	jl
5"2���3��n}z��<���3zW� [e�ʞRA77�K�{�NU�v��ɜ�G����I�"�*�UKn�r��>�ɉk��q�pRcj�q�=��$Y{�T6B����ަ��G�5�u�	�N�(ޖ�c/�D�����D$����͈�̙��;�{h�%d��h>����+|�uG],]��.ϊHz��@l�^�Yc�_XT� ��BaPΟ��,���>�a$���;AB��b"4�v���Ta{�+��Q��g`��o,�\���I�^�x�8q3n�L����j*߯�2k�*A�R�qdA�F*�)��m��&
�1�)��U����2M���']ףCo� �����qr��q���鷘 �"����@|�v1TtK < V�"�%�NN��M������M��Tv��۠o��8h ���(��"j�]��ND�`�Az�01�Y�mvze!�|��?�#�$���>.��"rA��ty�"�n������#�>��BQ����_"����U_�	�,������Y���$�����7�F.�.!�;y��3��ѷ��z4կ�Z��	ț����d͘�	n�^�N�r����	CXِA�����`	b��9��N��Z#(�=����&���^�J�I�	��v����Nf{�:,�뭾��᠔����N�WK�۝�ߚ�2+de�a�@Fu�ry��u�<��8�����rܥ�`����։#;᪳y��gt$������/���
@��6�?y5��g��eq^u�g�÷�敿��ڵNX9�E���{&��� �@��p,P�L�Ū��zP&�5{#p���̈́BXh?�g�|E:�򖾤���w8�BpA����W�I�2��֮�nZ�W�Ч˻5��c_���vԱU&�D��d} �U��u�	�,���t����
�la�R�4j�`��94qӭu9d.���V��Q1U}�dѶ�����!�>TNg7��Huj������B�\]�b��Bp�m%���`���A��w]qr4}ꃾfQE�o7!��2����~9�:ϝ|�Q���G	� �E�p����P��4���c"M�؊E��NNc���d��ѐ�T�����'��s����vD~�^[��4?��sܢT�H��evI��%��x���$-�b�
��	������\y�Z��Y)��Oa6�Y\�f���h�^R����^�ewmFi=#�
}?�.��7�}���m�
�^�;]��6��ʍw|�o
BϨ8r����T�M��?b(��zv���UT�����[��5��[k3Be��$2���ڢwuyd�S��{��*{p~SCp�q�S��������]��|�F��t6K�5�Nm~(�M����΍g�3,u/Ԣ�((&|� ��<�g�b�&j�ݑ>د����\�*��ܑg��$	�C�v�sIB�7~�x4�f�D=,߅=�>[���ctT�M1��;��P��$ÿ��fUX��*V�V��1�ׁ��)��)�C�c��X�E��	?�; �9��gބ���M|�>�Q�p2ʨ��I��kﶢ�Q�OFXkI�D )���$����;%�A_t.�U��?�#�Sv�f��h������`�����k�4�R���Q0�t�e��}N`��%4B���[�=ߤ�