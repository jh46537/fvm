��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}���j �]�ȴSN6��@��m�)��°����$���ٵ���\��T�iK�&D��	����3_%�.����,G���=�̷�|�݋RP���)��Q�qɾ1�`&pA���R4�_jPړ��{�4��.�D�/�l8V�Fwޛ5���]�B���wh#@�X�ܵ�)~�sRi�1�\�ubx�%ѕ��B���岝�%i����t��#�����px���vҿ���)�K���p���Q+�Έ,vP�{Ӊ�����GǷ3�� y�ߢ'����E��̐��0�9=�x�\�$z=��OdG���ʢ�~�G�'[�.�}�5I��w�`��-ɻ���Ox��(����łs���0���~�N&<ܐ�1����������0֌SF��5�;aW��I��ˍm�d�00u�;!��^��>�;2I;����I�ަ0�ڟ���b6�8��	���p��4�� �ӯ���Q��G`s�5�	&E�Fh9M|F@�(	����[�=���t��n2;O$�y����y�M>�G]��k��j������T�I8�
*�C:��b��c�f�bj�+-��.�����'X	�8�t���w���,�6���b��Ke��x�em)���"unߌV1��m����8�EKJݻ&�a�o	 ���FWC��Q��I�8|�Z�|5�&&ڄa ���
����ɟ��K�˒���!+4�T�BJ/0'U�[���;(��ա.+%	�30vv�7�������%�r���8�6� �����ɟ�30Х�ˮ*�D��G���LX���jMk��QWiᇆN ���F?���Yh��Uf��x=���c۬F�4��q�U���D������F���N8�Wk���a��3A�c�Gߟ�j ��ݐ*����*���Y;���C����[�d��b@���V��)N�e'��2��)O�"`�+��={�y��������!�fKׇ����]��M}%�pPJ%����j���_���P�R�^�zV"��p���9�TT $d,�Ԟ�Q�=�+�@4⤻}��j�O��R����D�2oX��- ã��c�κ���oQ��(a�qF�e%a3/V�:	}�xi�z�sĳ��t�h����J,�j�f���+�P(��)Z�r�>k�pTyS��3޹��ʘl�׎���� mD�.��d"k�
˦�F(�5ʦ�5�1 R](c�N4��dG�{_�rV��n��o	����6ek	�n�����3oTal�6�O��.L��>���8<�-��R|����7�8�7�������#WG4�/�*���b����P�@D�����;b\��A�����
+��e�d�a`G}e6��
�Cحe�������A�=C�G�`1�J�JQ����:��/z'��O���p�!@��Ww���Å+BrT�P�ѫ_/{���])�0�P���+�4�G��𩞠_��K�sO�/�͓ޘ���[^]a!jd���ʞ�SXWk�ſ�I�W_���B@�f� 儖;��]�d.zI����4���GA�����2Z�I^�,��DC���Aw �Z�T��E�[Y�Vu[ ץ��Aj杌o�Zg[��:+�Hc+���s�u�"zm�n��T��,��<��t�r�P����-�|��0E�H��a{Qa�~'�� ��+a�A|"V�Z��7m]�GK��;J�'�R��������M��+��$�	͸Y�t1�vV�+Q�[�Z_/����<Ki�Es�02SH�k\�0RN���PB����䋝}�̞#�򱰍�0D����<�ղJ*��o$��/��R�}rm�W
�/2��.G�#;_O����p>��f����T��`�FII�
VR�J ӡ}�t�7z3S2��xBc��t"�� �Z���dÃJ�f�Kb�7�Z���3�S��r�,]��/!�K���'l���b��5Q#.ڕ��g�D����`0�S0�M�؋^�I��p�yo[<�~y��N�K��49He��B}���]-o-�Y��]n3������>������j���S�'/��xg�gu?|���V����O�Sv��,��L{6kOV�wR#�n�����Šb�{�6���}�_>���٨U`$i�6��RM6)�����1TaF�Ϥ�֯�U����2��h��˾� �TO��3\j��)yI{�{T���5�!�a�RQ��*���(��]/XQ�riF�"�f&=��
]�;nA�'5kME��ԩ|��~E�=�t�����`4u���"���&.�n��`\}�I�Y���H�\����S ���9��N����U5�[��TrDHp~��⛯^LT��E_.٠I���I�N�&�bȜ��ṩeQJJ�pH�dg�J�z>�������K��v���>���01Kx��~ǙƜ����7��.:���՝����p�ע�@�U~�ss��H7�X6�v4!�������lԟ�A�s@������)ꓣB&�����C�A�g:t�ZVG*ܛĻ��A��)�=P�{�׆��XCi����EGh���0;�� V8�%o�=aFk5�4��K F�̂��N}����!)1��#����$�"���IY��=�h�Y�o�j�T�I�x���T:i}��*ޕ< ����\'�����6ˬn�U�՗��+�^�A�B`N�8W���`��dd�|�XHΡ��G+�E}T��*�x��!hLa�ݭ�|ۓW[	� ���G�����&��X�uUS����#� �m���`a��E&�>X��r� !3�0�c����ٽS(���>c	y��Ҥt�U[��HK�<e�`,��l�.�X>��� �$	�w�&2�aB�`r�*z˷Rb�����]?�����@R�&��S�����4��� ��D
����%L���4^z��I?�"ɼ�=�|�\�G��<p��S��w���/��j���V��ݔ��xu�:UЫ�e�N�~MmI��c6^�'*�6�s ��kF��bu�c��.em8V�ƃ&�\
�{��B�r	$t���^��-���j��к?�	�X����]̷��Yn#�v�@k7�%�F�TEAKԻ���=t�$����8g� Ocш�݄�Xp�k��*�g�����l�	J>�_���N�Q�H,l��˥��1�iŴ���7#鶄N"��ݑqd�Y|#�U�Q+ s�^��N��.��O��X���\�+�8f�-(�d�`�(�x��?/$/0z�s4Ou�� �8ag��y���8#y�6R�����nr�	n&O�O�7"�q.�!��/-WH�1��պKǘ^E���?Љ���n��B�:={�N�IV)q��\�3^�d��+
�2�[�=�メ�\���*�`5�~~M���DV���%����I��E>�'s��M�{�N���QH1@wM����@O�
�n��3���٢T�B+E)fӶ`�?�د��1b�v�`�iGHg�:j�Y�m�d������i�{��1P8��bVO���lTg��Ap����g���K@�1��;�������C�mKA��e������٪Z�|''���sX��.B��5e�m;4�y]l�C_��U����h۟�+%�)b,-�����>�li7����tQ53&���M��0��'*S�aٶt,�M��p�$jϹ�b6
ߊew�����%�(�T�u99!��()iZ4q8	!����5F�cO��+00���dS�k�Z�����)�2�>���i���D9�ա�D1�v���u���NX�Nt�ք1bO�r�zy��o��u�⯁�Ӫ�@Oi`p��[%&�JV�U�
�ܑ؍�K�~��nu0��(g����TJ-��ER@�9UKB�6�F��D|#-�>�]X���?y���iM�o�ǦG�xTd{#(Et��һ�������2n��Y��
�o�JWv��d�ۈ�u��D���M�wD��l&�/�<v � ��5U���S�����V(�����8�@9�˟��	Z���S��u.�r�"϶�D�*�s�>�!Wx�`�X����n���ᬎ.��>ҵ���,żW��C�ylV�����7�C�4O�SIQЊ�l����s�6L����1�VW��K�3S�{�v{�yS.���,$���R���lHX����T�P=��j�>g,���%aK����F�b��*0,|n�!0a3R��c.�{�0�<P�?����a ��74E3%�.��k�Ǚ�-aE�#4���C�'��{���� ~��5�q��V}�t�o�U�TV1U�~�r�/:��� �Ҕ�鯴�P/~�hKŷ*K�����j�-�{y�O�o�{uz�i�m_*��*"��):\�,���4V���ѩ���j�ͤ��kD�@��r�,���.dUB�;qp���B�1�c����Xv���n;s���$QP��eF��"-|%C��[� �C�8�.� �A�f)����\A<��┺�L��!�5��:�g��nZ��S蠜+)M�ƭ[�
�.��%������p�6gcC.�o�3�q�pw;.��OȪ�~���[S��� $}A�Z��5���,䚨��g1�������g�M���5��Ýˁ/�k ��Ąu�Y��_�ȡ�D�TJ��?� Y������o�B=���.��{�ʎ�䉱�MA���sis:���{���M�[�O�x5��f�>"[u�x�ڎE�q=����&Js��^��Z�i*�I�\u����c�����dq-��n<����L�>��V?UM=ŜO��Օ����s��&4��Ȗ�g\�A>=�b��<�
�@���*͛pxn傭T�A�߁���Y�(e��}�G�˜��tp�v�9�ٝ��${5� 0N�iA����9�HL�2ʃ[v��Qљ��DV�����8�"�&��q��d���L41��=��!e"��0Ӊ&k����|@�����	̼nb��"%�b.[UCƨ3!Yр���'	�o�
�Ɋ!�c!��Z�U�-��(�]�t��Pt~z?���h��p��π���j��$�[�W���ȣ��/����82���N���D����`�8	���$)ql�$�n&8	'�[�����.�z���<C�K���K���ƱM�J�"���_�G({�[E�)I�����s���y�8Pl����:ݔ�H�!����F��k�-5G�J,U���3~��r'sy�CD��nܐ%*������UбxC���|��)��U7gUN]�^�Ι�!b��M��֡n
oA�>��7Oz9�{����@m2��?���}A̅�Lr��K0���R�p+���l���I� /���գo�\�w��!1D`�Ŧ4e|P㳞��<)]E�^K�T�h��R(�[�Z�����͏���l�q;׮U��"IE7C(�SF_�C���4��h�BB�[*䃿�"�ǻ��3l����o&&߻&m�{����Z�-g�@��O^����f�o%v�5�5�`����&j{�N��2��a��j�¦��i�W}<�B��G,�9
������ a���v�a��Z���^�yV`���z�O����s��;&����!��Oi4����gf@��#��	
ߟ��m�G��~c|W�S��5�CH�*>�*��-d63V��Ծ�8�� D��u�Lj~��I0|z�#*F��>FϠ&M�Zf#��i�+ѿYZ�>7������=eI�0�x'�ԉ��t~f��g�H����g����|K\�y��pV�6�?�KG�2��x\��lp��{�&����2�57V|*gCG�y�ěu�r��c]������v�"��b��0yB���S��tH�?����p|�T�ܮ]�=���3��n{U�)fM���$�a���:�K@h�����aTJr����mjs��۳c�����.�����@��"G͌���¦�u�zu��
h9��&��{J���}�uv�Z�I��g}�F$IH�@r֠9�}��������R��o肝�T����/�о�)��:u���W�
�'�e"sv,P���S��.��W������'��з�6p����`�$��X�+��k.c.A�[S�Vn�@����A}�n3�6�hC��u.vjk��;5���(-�>*\0���ԃ�:�{Hyk��/c����v}��)�
�����O���*�&��q�NLXNü�� "�}���]�S�w���f)�N� ��w1�U�%"�8j	���
H�)���fx��O@��=.��H!»�*ѺQdGDp6�(J|sY9��e�!<�eO�4���f�ß-^�:�{-�����?`�n&��x����Xg՚p�ew���=���U�-]p������c���#��D��<�e��������Y�BQ��}��D^tG���_ke�jjG��d���cH��=<��;Y���e��B[�7�6;)�u���2�7���k�5����������Cu�X�[���d�n	��*��p�.��eP�d�'���ԊiGE��f5i�ZJ-�}�,���["q#�j����MM$k��.H�b�Y�����I�ky��v���E=<	n]��x�K7��t#�6Ƶs�Z,�퀳��	>vi�9�v�����h�s(���Z/�vtIϭ��;;��|�	,=/46�t�U���MW@dZ^O鏔́��d����,�Ř�g���O�g|\ZG�Z�Y�	ȫ:s��	N28)�Ic�꺀�
���V���e���A�)��xՑW�Å cv\������ $��Z�[�p\����[|�+e�x�N�1�֚w�^���[��B�#Mi@g��E�'�G�E���R�-k/ڥ�i������$j�F�|�ⷡ����iK�s�Z�H�8D��e~��	1����[CwҚ�u�G��7�a#�(8�z�	G�)��<�@.K,E�?��9�x��b�4<��v��ъgZ��[3����RsMXɬA���]w	�jg]�������-�V�1}�����]�*+�c_k*��o�Kj=6�P��������L�?/6�}^H�"Ǻ&򚃿��$��m��I���V�w�M4���[�|�B�X�#�Y>�p���~��x/�|ު��*�r�*,Ft�]�=*����Ő�7e�Z��� �,�xn���a��ml��ѕ�k
��3�5Dʝ,��jTu�-�u2�~��۞Pܖ��7��H�P#��j��:��U���y6	iA����_�90����w\*'.T&Z�d�=�,�����
�Vڶ
/B��;Y���EW�<&�'E�;u:K��8O�g�O���;e����9��DI����7�d>��2p`1>p�@V������kP��u�`����=k� �;���x�<�s{3R1%%U�׉�9�/N��F?w�G����4�¾���uG��jQ��dr�k�`����b����r7��57��n��G7�C�SQF����wU�,� -���ZAa���>Z�E��5�/d&�M�Zޣ���B6��&��G�ZS��Bo|e(�|�\ܬ�$6��w*���՛�0�,H�'��N���&_9{��M��H��ߧ^�Զ����Q�]���HB4(�������62���VA�C&��ܝ�@�'�/ '�9>q����i��y��e<4��kV�`=�
����TS�p *�@}QD��G���o޼�:"tu@n�MRܤY�m��" �j�%C���ԗ�Oj��R$l`���3͈R͎qզ�z _fA�@I�YDX���G�=@���$m�	����6���5p��[*L���F\��o�<=��k�g�w�>[u����#�|B��A���V�Nf�N�P4 �!��d��u���6{w`e
�˂�)e2H% L=P�sm�`6؅��Z��T�����j�F�� ��8�������i'��CD܍�)�5*Qݪ�r��D̰�۔�]BQJ��@-E<!văB��r�V�ĉ��xq��̚z����]�j4bx�-Qhy�i�~'�3L�M��rނzח�� ���KX�э�]��~O��NR*G��z���?&��l���"�WT:�'�(z�J�90df�y�6}ǐ����@���m����㵱)�;PH	S�KW�=El�5D�����d���9/�%�S[ n��^L{����X��?3�p�����e{-���h��s��5Lr�6�U�0=r�GY�i-�7��=���� A��|��X��XχF+1��#T�� ��%V��J+o����1�lHǆ��J����/�B��&g��6o�H�_�s�*�J3�������/MoLLK�ą�T�G]���2�uv �$�������5ק�u��%R#0c�5�c�n�UGD�.1,���I׭=����T�M�����u�����2���-�7
��_�N���Q�q���:�h�R���z~�8C�3��Y�}Z͡�͞��[���#���l�T`�麨��ɩ:��\��`�+�6����"
m�� F���
���4T���yN2l�DU�a0�L���:d��k��=��xH�r띿MpS"�i�L��H��}F7�s}x4Ң�ǹ8�_N�������S�R2`<�-��A���8��:'F��J�D ��}��(̺����'ڛ��Dr���!���T.яAX���6�F+#�"_7��[�L"��|�#��qX$C������G��C��5H��m�ԹLv]���d:dV�}�aC�I�zleo�qa�6��-�ٖ�{��AJ���]]�5jZ��#h*
���}fT����#����G�ح���ōz��uE��m�[ްqAO[ĐG�r#���Hk��R1��'>��z�� j�,W~ʛ�ԭ��ս�y�kU�3tOR͕ٙ��K*X��L���`=6��o���0�&�����ĎG��N?)�����~�d��_i��!�a�=��q�����u3�)e���2�Vw�!�C�iIV����&�w��u�� ���C�f,�����K�`IR@fƨc�;�^=�Øm��#��#Q�Dk �m�_����ہRB`r�#� o�U^"Q�&-��^Թ��o�D���܍Ĳ��ވc����0�b1��N'h��`�Ϭ�NP�lBp�(g�Q�s|��F��?X�$ =
r(���
H�V�^����G,�X�TJ��*��5�Zp3����E�N��?T�K��&�덨� T�jʶ}�1���OH�@Y�޽J�b���.s�0w �N�7�	��x8����� ��1�RO�c�6CˠZ`���)�%M0v�3��A�T��ç�{H�^?�������l7w�c����dA�l`�D��fc]��輚�W[�0�,�P�5'É�~uk���ʏ'��M=$b_�@յqBD���St�&Z�V��d����?�Ȯ��[��
.��Y`J��i�}
6�)�U����9�-�ykb�����j�"3w�˥R�5���������%B��Gl5�zțLv��_���� ���,��cК"�#�&nzu��TO�K�U�����q�N�`^*\W�;���MP�ұ ���Il�gE,��$�՘	A�F���=�9���Q��t�˔�d���@.@H������gv50}/���>W��N��0͝p�����X��s��wFM;��t ,�z6���mƕ�:s#u~d��-A�W��H��h�<2��C��n������Q$�۔k'�R}~�~%�>�0���"C�i<Q9D��C��1���D�$�}�j�ZԔ|:3tiw������ȯ
��X�2��%�@NaA��avE�@m����NZ�������+�0M��MZ���<7ebk(�FcB�0�7I�X�2LD�r�:��w��b���,�95����h��Ғ\�ىvKz���
>b"\[��S/^�a*{��_��A��6K1}1�祭���Gf�M��#n������<�x-�W^�cI�^��H(,Y�'�Ӹ��g����F=#�Տ�R�$����f�6�'�/dF�%G8�J����ٌ��&m�N \�
P�Hb���b�������b�<�m~o�!�j1�	�!�!چk�bV��&S-q���m��RU�`/��#��u@����|wE?��4�B���;��Kj��E\v���?4՗��O<6�5;pn�@����M��j�Bd0���fB۫�D�5��V&���g׊�~ ׻�|�4�|�����FL~��w�2��)�J%�ݛ�VRoZ�3 
�|��<�So��dh��z����}z�2� ����Æa����ɪ�˧z�]����Bǰ���f5���;�[�6�%ʙ��"�/�����Z�y�iBCbmv8��jd�zl��G�߫u���T�o����JRo��K��q�"?���2����2���-��mz�(��6���)��C�����cs�#2�P�I�
�q�m]��J���}���F�;ax�"8='�wq/�L�8���C(��:�WS�*|C�5[�;Nh�}�kLf�I�/c�W�7��������H0�v��O���=�0Zkg�f6��y�Ƀ�N\��\2�q`���]����� �{�;�����-�r$g6�/P�v��7�;�qz���}�J�-�5���mv��yDY�ð}��t��-��tw-�l�[����1��ZD}g���y�tV.Z��Ic����8u��(��t?3��<��q[Z��-K]��PF�V^��d���J��� Dc 9�7m*��.�C9̪Y�B `��܊����6v��;��q�)���wg���Qn�KU^D�O{�j3#����?ޤzR֟;����k��m�[��e���0�zs0-=S44^��8���H���Odz��YZڱ��E;����O|�����*�D��� L�W���8y�ٌ!Nw	?$^�K>��,��6�Q���G��/\ƛHv�D�q�I|%�l9=��|��H����,lbC�N��R��d�-�̭�(ݜ��u���� 	�Q��Y�QH��Y�_a���)���� �kr����B���Bؗɭ�a~M�% ��6��|���2Vv$(p��թmr�j���.��[[;������b�A5,�pD���
��0�0o<��fE�i����@��tu��2��n��.�YM0�Wݾ	C�[	XZ�Zu]y������'������dk��!�4�K p�ȹ��N�n�"�5���������g���˽!�.B�}3_��V�ot\���s;8b�]Jy8�F�@*�!t{�A���@uK̖�6q	�4�/
YwJ{<^�����(L&�22O<���K�˽҇�"��p�e�k�C,���=W�'�C��]3�٪�h~�P~���@;�'X�zФovk滺CGçi9ʪ�ҤxT�Y�ֆ8��waP��z4`��LR��)�x,�}Ö�"�" L�z=� �i���0R����F?�[��.��s~�3>|^�W?�89��R,l�^�l%v���M������͂�K>�G
�5�����~f�l� (LP�U8]f%A��ZD�-��)�K���"�Q��HJ^��+��5�=ڑ���w�D�5�?���uIЉ�3�$3��Ʈ��*J�}���i��+�$]�O�b*,�7s�%�6311Ve0�iI4GOcEg��2�W~�o]�?�1J~�ظ�FN&�#��V�ŉl�rԞP���5������`���#��)���|'�`kᘁ�����ߡ�z��;ڸ�e{�2�cL����ؚ���*�=LҘ�K*
g�Le^@#��Β��N����a7�L�yna��5����0���͐f=�R�o�̈���:��s���{�rA�΄�?�jm̜�e����I���2��U%�&QGm	���e@ �������.L�6��}��U����ՇY��v����F����Iӈi E��f��aȺ�u�19�V�ay�m +��h��V�φ��g�*G��u�I�=j�ܒ�rqn�O���ފ�Itю?���-tb_�-�������;��hˆ���7�W��^����yڠvh��߂�1��_ #��y��E%������m��S��fb"�X޺!����+9S�z:� Z�����D|�p3��e�K��1����j�AF��F�:�B:��шRV�
��u�g1�ڷR �-{.qD�<�V�sű��![��Tx���]>�fZ.۬��_p�hl��T�gZo<rX���?o?������%��8L�y�,����x�"b�Atǹ��ҕ;A�����5�����s��Q���Kh>x��@p����	m��f�c <����>�`w�$^�N�Z!���ӳ�Ģ��r#`?BO��_���
k�N�һ⺠�ع�Ƽt���8���^��f��&�= �7�u��QTaL�{�ͽ��q=�|Ԛ�_��>Nڏ�ޮk��0���*��%�dG���+���V�����\��9�Sy��k���Gz����?���䁿e��==�0�q]vQ�)P�t�ü�?�1f����b�@��w}ŀ������-=��T�>�,)	�EΆz��E���7�R�G������E�l��Duf:d��t�e��f�N���)iD��l��oڷJ��p�\�n��qV�ȉ|-����=ć�L���E��TxJ���E��4W��t)I?+D ŖTO�\d5��pj�yb��4���s㪋j��;�Y���U_�6��k�3����W��0k3з	�O2#�e	i���R�vj�U������>@���w�݃�S�Y-C��R��}\8�%�#�W!ˉ	��J�i��H6O������
�l��v2Y����f���iDtL�Ȁ��#�x-ԫ��r%4���=� ��3cr�(&˦%ap��;����[�n� �m�h�RI�$�?|���<+H8{�K�R3{h�v��|��)D��6�����뱚-8Z�T}:+I_�J����)�O-BV�=�-&I/&Nga>bv�4��t����*�)qr�����9�����I:�+/���B�A^v!��x�ϴ�Kx��cҠ�l�P����zv�����s�bOO���-G�h�^V,5�dL������B>�s�n��LZ�ڗ"�3R�̽�OH�Y��=��|%��V&kF�t�����\8ݳ�n]��đ���]�G���-��Y��O~X�d98/m���z]�c|�a��
��
�Wt�?��[QĦ>Ւ#���Q�BR3+��P��(5V��QO7��n��:�њ�|�����)�?H ��e�?��G1����{��jv�?h6v��yN`���`�V!
�������[u�����/�h~�$�[v��h��@���c���eg=x���]���1�ӹ���H������f*�yd�ISKe��C����l�����M�Sd���!�?�CrX��ȶ$yw��t9�4;�fan����:���K�um�]��߭Lo��бR�(϶#�^��KDa�j6����|�X��ٿ�4��  �v�j	��L���-](�I�;�^���	q���FJ���'0�f�l�2��Y��ȞS���M�LP	��^hG���ʾ<�>��1�7!�_�Z�.UL��h��E��"h�X\�
<q�3���M�	i��c�T��~�Wux�e=R�&�s6�7���z
Zjjz�����Ӻ�s	�n��<��7!06�K>�����U��)�-8�lY�O)_}Z{}����	�K^�UW��X�3��p,�U�<��A(CޚVi�]�q覸#�2�|��H9w�J!�p9`^g�D��uͳ8��\�g�����7M���`|�QB����߄�r1V�E�b���v#�,:kV\)>�1[8K�Q�������7yd�Olѧ
'f�H��[�����iE��ݚ��N�.1{�R��h)n�!r%G�����sn��1W�<��F�q ��C6�`��?�5[xP������T� �O�w5�}�񮨄�(In�@9�c۵\��N켯�pS-�4�o��/g���b�zk%����[�z���F
:��ӓ,�C~]BV՝4	i����)���5>@��N��JV5�jUE��S�8�7�~jc��P'3�e�>6��U��^a��܄����=�b��~����H�D�&��ZA�K螘�{m�tS!P)��ֿKdA*��*}h�1��b�9xȤk#�uX�w���\�	H����|sD=��nr`�	�!h�����V�I�b�L=C�^�f��d��� �w�-Ë���3�Gʯ3"l�p$��x�Fs��ѬK����S(�\^��u�{߯O뙢�P���0:I��"ZN��ᨤ��"���v��z�����r6���#�U�IT���@"��9/=@{�x%�o��T���jP^�N~����c�*1��A��e�8�R`�[zWM8�r�ǝ~e�_G��.R��F����!O}�Kei����R�[{�!���aF��(���4��ښ�=�JZ�����P�� �f�w���5�?Bj����IG��� 8?
Ot|'�`�ٝ%�Y25Q�J�G8G~���p����>��
�C�*��O�^jci�_y���d�z�-��j�)!�O�pq��n�o�<��azb(���6����t^je�-�+"^�=�.RW@�
�XӤy~����R͍�>�,�g�=��L��{�^�K �a�L��3ߑ�4��hA[䀨Ą�V�R3��0���Wl�,�u<� ���#�@�r�vW[�"��D�/�O:o�#)����!ۊrG}Vy!�2��+\�;5�,����1�{�1�\�Dѵ���=���v�M�N89����1��֒��	���<GbV�O�6�!�4,��J��\3XZ�Ȋ���M0�����-�Il����1�%��͈���b�59��^��Gu@,H;��\|�x��;_@�H��d(?^N�5���m�\?*?^x]9�)M#X`��t���#,�^]�i�R�u�H�B3�:��'�L�Jq�\]��6]�sc睧�G�A<��`�##Hq�Xo�&�� QFL$|�d�;F��+t���G��t��w���p��CMi�´#MR�f� Z�v��ZQ���.����h�1CЮ�n�Y�W�Wt7N�7�w]s?�}z�ɠ������W��r�$����,��?}f�+��־ �U{����r6cZoq#�쀔���{�5>�q>�-�ߨ��y�X������V`X�,�!���'���[C|(��T� �!J�0�A��ԛ�\��0煻p����o�� ���� ���m�bu��Ŗ��չ�`߽w��0ROO),�D�w���6TQL�ɘķ�A+�ث��)��;�.9Be��Ψ4؉��<<[��f[b��S� !j'�БCW��%���BN&�ɠ�z��ߢ��Lw�A+�D�5��r��}����\���pan�~̭1��o%�~�Q6PH�����q�ϔ���vc�8�!�O�J�Y<�����g�tw�u���B�hA�,]-b>,���[���G�pE{�O�Q��XK\C���@�F)®}�σ���$�/��y�m��ɮo��y����h��=�����z�ܭ�M��T;輪䁻6ncԛ}��ʜ�V�2Җ�sF;�*�B���F@۷�K�^f�P�|�8�9)#����sJ��	�$���*����X<�5�Sj�,>�̘>1d\�x���ݖ{Z|�/�f�]c�(��Be�P�)^�@t�\�#�%��0L-���P���U�!Q1�ǁ�f��_��N�q��rw����c<�~F�'M߻=��ؑʽ�T�.�k� �vn.AZ+m���Ot��7b�7�ևڣ�l$�KajF1�7���]�X3�1R���
Z�4�-�%a?����T�A*lBz��(�!��k��a����>|S�����+�����#�?+r*`��ʴ��*�bP���;�g�{���tZ��Vh�GL�w�:����4�-��FWZ5�΄����9��z\�c݃��������l��D	ބ��9��
aPiU����t��|y-\'PXk�Lm�3�>�sI�(�=}(i�L����l2��3)\����Žs�Y���0�M�����@��PSz�DeN7{����3%���-���$h8�P'�E���LcBvg���Z�,���t���-4��F�V���_Ow%6�?yJ}#N���҂����^����x�:S&E@�J�fe�_���^�F$j���x���Ί��7Fg���'_M�T6����q�S��0
�4�΄R%��B�W2�wIJb��[��z�(�u��}���@�d�W{]Hq��&����<���_��.OC� ���)UT|s�S�.MG��A��q�qG�E9i{�	��Sw߂�ߴ�cu%̯�&�k�Z�)�����X8��JE-$0���f�y'_tʚ���V�ϗ�$t�B����q�i�V*cX�6�вx��#0�f��j��9�|4�w�@Y���7P\�T��+��:�m$5�,"�3|I�=����F	�����t%8���L�����8D�R5�o	v�Ͼ���r��\���}���Z�@��kw\��{�3+:�9_��R��K���0)����S1�p#]��xhi!n��h�n��͚�/�ͤDhuN�tQ�@d �-��7N�(��� ��+��4��[��<�P���G�Kz��"[ݹW'�?����#�~�M�YOS]Be�?:iK�V�+ �Qpq)�P���_�F �ܶ��>���'R�q�m���vn���PO��}C��"/�R�nĚҘ�� �Ó�]a�8i��%ϕ���@`�/;td���tdV�?d���������l��Q6i�K��.�0
��Ŀ	�����f����ؓ����,�Z���Q���O_�����i)�k�Lh�&U��D� #_e�(߸7#��1��ܺ�R�a�|W�Tv�T�9/`�����������|����!�e^_�f 爾�2���������ļ&����U8�>*A-�Ġ/��R۹���fg�a��4Vm�w�\��'7%9�^{?�����)a��Uā�I?	����e��C�p�����6b͸h���=چ�sY����D.����P�}}(����2a��!���s����C'/��U�S�2k�`���($^�Z#d��cV�>Fܢ���!�ŀZ��PN�����մ
%uQ9i;�A�Q��OaL��y�:G�,m�I�����i�|3����5�ɰ�l���`�=l�����]?͈֧߅2}s�}?��2#����ڍB'7���]$�q�MZ�?�z%w���+Ԯ�t#u��or��	��'���v�ȱ���ҥD�QTOst��Ij�\��W�X�G�P��e���ca��(��9K5#~jr�a`��6%�*�g��;?X�U��&���;�
N���F
��#���RYH��m�"�z�<�D�K�{�l4]?O���9B��
���`AQƀ��-F$b]���d���[as?��x/.ɐ})��tĨ�pVQ�j.�FD�&��,��]-'��q��@8��<^<:��B��%�m"n�j%��F��_&׃Ǵ�����C�G�S�G�z��=�uՆ�&2P�>�+j������t	+��iѼ�a�C�/�a[�?����>;�s�Z�;_e��fra�&�'·�ݹ���	dR��ƾ	�L�0(��!4�@:rF�j�������e9�Ŗ�9�Q�������Ҹ�/d��F�,��G��6�!͟{T��
�hڒ�y�-u@=�����;7��ơ��=���6���ؑZ�t$�n%@�����Ч�C�n�2b#��S�C����PDw� �����'�:yh����,}����(�����ϨR!G�ާ%��8ڲ�����)7����G�Bfs��w���-�~�\X���"��������i�|x�Ȓ@o�a�Ac ;a���5u��S��t����S�;�QN��+bi�6�F���I���pB��F-&���o�0�(7�F�~t��|���g�Jn�"�=�/���z�Ec[�a����d���vN�#�rz�&��F���}�B�PO/�
�ۜ[�˭�:� J���&s �_�d]�x�ߥ׼���N�^m�o>M�����H���w�$ce��4"��bK;�YHI��.&�Ȣ���y�O�Q�7���:j\z(4{q6�z�3j��r }Ż;��c6�'��`X�1���!i0��e�X�u�8������������\rW�7����(���j�V~=;�[��ӄp�9��ä�{��T��a	&�G[��4~I��?^K��p�{%�:e��5ޟ���$��N8��Ԯw���D����f� �i�+�����cׇJ3d��'���\aZ�u����'W���0��f�~],o�R�� \��M�ڶ,��Ǳ~��AT�����ZK��4[�0�B�qMn�&P������k�h;��)�����P;�6�8�<�i�'z#&Cb��L��2����6Q��G�����g�#�NT�=�6X6ؒ	�W�;�Mq���[�'� s� �<\�:��gg:zO���>WI<�@v��@X�b��N��4s_l����d�}�C�ɱ3e;���k�Q�Gs�{�N�!�gq��ذH��X�j��糓������=Q����L��jHnd���1oa��i4���7~Bh���+����UHS�L�+|������B����-�Y����T�"(iD��j�H�O�����|���h2�LwSmF������l8�V`4ɍ���Eݰ��-�$�ϐRL1���{5���gU���DL����X� ��m����Ɲ<Ec��h<�H�P��U�,�BO�:�W���ں#}x�ק���0$!�R#+�t�,T�Y��Z ��{i��(ف�NF 'w�������֐;�9��r6.A���V��҈�ڂAq������Hz�k= �6�%)N�S���F�	������Ԫ*�<�U��`���J*�}c��$0y[ �W����=MB<��7PU�\c�}^�3]H�g��q4F��k�$��q�Z��]l(������l��������������x���n�(}��h��\�c�Yw�������a�3h��mE�����uf�����Ћ�m�>()%�6��{61.��w"�P�`s5��c�!c!*�2է_�t�Z�x8#ij�N�m(h����y/c,���ZКC����K�
�<hR�;o2�ժc_��3������'��V�Q��8�d�]t��\>E�Bо�4�ݴ�`*.Ƕ}K��u�
gPQR��O9(�^=eЖi1s�I�g^�T�W@��T<�61�)�5���<����#�~�Y���)��Ae�ل�
(l}WC�^���4��u'�%�h	���G���R��͜v��m�J���p!�VyF_�����N�.���<"�oÝoc0"�z=�4���f��%:�{���렋�����A���LEvM�J����f;�`nz��������{ V���a�?��(&��E�ʔ<��F���V`l����]�Z(�x�e���x�|���oCs���+�Tx0h�j��������˅ch��#��=�����I;���K���vFK����)�{��A,POI��C���Wsm�hZ/q�·�=t�cBL��&%}i9;��=�Ҭ|�I.Hy̙P��¡� ����=�.�(M2gn��dS�yvַ�f�nga�����@{���dJD�Ea R���
k|�TL-?�/:�ՇI�"/$�&&$m���C3�T��2<QQ��i�[q${dg\���v��S?5T6G<��� [��7�@�\��ҿg���AT[j����q#'�����/!G�b������q���:+�*�a�CQ�����T���{��m���{MJ�C���}w���?��
_�\��E������� ����^ ����yicj���}������ϥ��fe�]�S�S�x��F��1���rb"����g!�.������3�d���� ��`Cٞ':wL:�۫����ͼu���bL�*|_V��Tތ�.}���l���&�N��@0�w�E�!��9����߼���Yj�X�o�Ss`�.H���X7րOmM�����!<8�xGK�*��b	}7-��/Q��С:	��*�����Q�ˡ<rQ�H�7�M���;Sx(��[$-��BJ�b�c����k S\�O.w�_�讄� 
���+oI6�c��N5yw8,U*@�a&����2O"YcQK=�X�*[Q>F �;��4�v�b�^=�>Ǔlr(Tw��hT����)���n��5;��W����e ��H�}X���>�,�c�S��M��`�5��ӍӞ�}�e+�a�h��%�)���}3�j*MU|�.�!���n�g0,j|۬^��A>���4�/%�/��h�}6+BL8�Rv��J���v mw����+DF=s�UI���
�d�v������3��H������%�,I���P��w�KSBT�fC��QуA!c�-��!II}����1˝�J�����O��;�,jM�1�ﾛ�#Cߔ�2�:��ʥK�b���(������sD������gS��`��c_w�ǥ�TFO(����.��E��,m⚃r���LJN3>5�Q�MIΟ��1�~A5��].�j*V�2�B�;U��r�P.q�q�`a���)��"&�u�/JiC.U��qZ,|T�u�<��[�S� Mnt������>{�|��c0ܣv�%��n�c���� J�_7<Gv�@�U�Yz�����7�� �6��fX�f��H�|�����i�q����.Ġ�M �c��!Q�� 
�s����n������.\�X�7A�����U��un�ڧ�(#�wðC�$q*�s�E}w�6]7 CĞ�2�������0F-�-ƕ��κ�O����_Q�e`���a�C���jd�Ag�Kӄ_B�g�!�z��u1%����:������$�\J꛳Lm���k"�Ɗ���2����|�[T�#���]�Z��¹�x�*{R��٦`��GZ�(n��E�()�3w�מ�
~g�6_ے/�4.b�������v( �Ŀ��z=�sg�(�6{��g�܉6�lk��&��y�����̏���2����z�z1#J����Nl/o���a(H�����3�T��Hj��SJ��՝���b�>��[�î�db(��������j_HR���a^/@��t����ra�)$o��PPu����I-���%�6z�qa����-��/��
��ig��wlm�C�TҘN����Bp�x0����0����U��`�����Y��t�2���[/ů�����5�p6PN�����]_@z5�n���I���>(9i~��p��g|�6����W����ţ�����`��H2M��}�0(�����CB.��� +�o����ʚQ6��rdN�C9�-�Z�>bz|[�
�V��PDu�R�������چxWA?��tg�=}L��[y�; �d� �~���Mޜ隥ݵ�
����i�vX�tej1y�������ܡ4���d'�#a�M����IQj$x �9�߬B� �/R%nf��l�]��n����n���Q	���z0�r|}���!���UW~��&��Bolr�|c.���M���H ��	~�]mt�2����/'����+ֲu,�	R��B~$�	�H��OiF �='vm�8 �-��)�)��_w�-�6���2�n��( 3C���>�$�}�����0p�sBަ���H��w��ff�z�G�c�&��?#�YEsE�*�9@,�Zo��*�Juf�����ɘɣ�7���l&5���H�ѷ�I,(�)�c&L�
��Fhb��IVr��x3���x��]��ԗ��quK������~V�F 7��4��WZ��T�8*�m��oE�]����*	t������A��'�AF����Zu����8jy+��*w�T��^���i"��Б^���2*�������L�G3������)��YQ@���}�X]?۠���L�r#M@*zޙ��$BY��K��>_��8,�r6C���L���Y{�T�>��L@�_�8|ztB@R	�/�y\�o'}q �_l�X��o{i���$�n��o��$��7ԧ�^`/���ט�d�p�<,�*|o��]3��_�C�CZ�s�����q_c����Sl�K$���l��_2��qtY��I��Н R���0华w�S9W��{�\�x�K�G��%R~��G��Ӈ�����]iA�T��s\�g�_�!D�Қv���iԟ��ME"�!(9G�D�srOg���c40<����uK� ��<3���}g�{�L�؎D?�gsJ�"I�>������&�!���^h ���ˍ�ӒDLc'� K�#�X%[�n$��(��D=)�{H�rX(�dQc!��r��"�T��sH�;mh�4K�x���O]y/�--���9�ǒ �*E���n-��^Jzl�Zp�᎓���������Q���~I%�V(���a��>��h�U���5��4�c$&�(��DB�n������	-�!�o�|�i�7!,���C�h���X���k����B�XT�9�C��ĸFz��+�ZA�iO3��Hl#2�!���hjVn���zFل���� � >d:�c�jyR������BL4Ü�,���9"Q:��
4�څ L;_�:���tQ��m��<������ +��#���;}ػ1���_����3�\�ꬠ�C��lxÒO	}�Hqj�q/T��R��:"Y�S��4��u�:�!#%�q�Az���E�(ajf���u-�r>AJ���.*�
֠�hβ�Y*�S�׋eVCV��<u1������ !eT�__��61ΡM�m���:�!��.�������7�p�<��4��N.�9+�vc3�[�+<���Y�x�0= R.ڟ'\���~��"�G��rn3��{����>j���+:t��G��=�Nr��j����nm�(����/��t�R�[(e���t��������`���q�>�o��P5=�o����+�{?+�
> #��
�n,�p��+p���;��OG�"�詐z�I��~�d7��ȼ؃Hp�XV���nu�1���j}ւ�u-)���,����D������eA /��c��Dv�]�'��J����῎�_k�Ĳ����.�-$i$s��	�{'Z�u�ћ��� M�e��s&�ZW;6��%Sݤ�{���|�g��_� ��cJW��tD輠��6��Gs]fZ�}"�i�7-o���8L�n��\͠B�c�eB�K2�AQp�i|b��:aiP�dH|6��c�R*w�Ɗ}ү1�L�76`�B�&_��y��B�>��JEV���,p`���m�Ku�i����Ģe�{%�
��w[��4��i
޷�[�+�� ��NO����3#����դ
ҍ��ب���)�u�]�&�BJ�-N�R�r��Nx��?�����g���m����_�FG{�{�5%�e�8<覬���['��*P���Еa�}Z��n�LL�@��lv�A�8��ͰO~�&�����h s��֊��In�	����c�v�A�6�j�������y��������m�6J[9S-���4���'�T(>�L�<<�(_w�lV���6хG��{�Hf�]�n�,^(�4HpA��7����^ז���dK���Fk.f[d&~d^bI�s����������u��;o�$�ż����J؊��uҬ���W�8� ��n=���ȷ��;��.t��1�����ۡ �Ǚ�f�2;������=���ƛj�9�������+jf���H���x����v�K'�J����8!`�*>!w���������LA(z�X�f�cQm?�uO�~��vf .�m�$�H���H�>��瓷�v״U�D:�`-PEʸ�!c�h2ޥٜ+Ɠ��p�w?B�k�G�9�x��wLS:Om�&��\���Q�A�%]�H9��g�������$�K�@_ʗ�e7,(4-W4��cӕ'���m��� ��ju� �V�&����Bb���>�3��@#
=@���4�䊖���4�z��t>f݂z6؁V�-�q�jӓi5^����í#Y\��Uߟ�ߚ?�|����F�K�}]��wm�J�'��t7��c���OB�}�}L	�*����hOB�$S�?Z���.٣��5�Ώ�_pd4�l�&(2�X}��[�a��X�z	�EwZ�/U�C�#<�@<�mlK*�����鏏�(��ՅEt.�ĞB�"��)��ڂ�*A�}����*��=��w3RM>r��h����s"�|�|�WD\�?v������np���b�qI��N$GK�x�"gC1��S���hF��
�o?)\���a�%�r`�~�� G�}]E��Ǉz�$zD�|"?q�J\����!�I�T^�|�t� or4u�³O��Ȉ��6ML�oct�i��=���S�q�����!�^˅gJdo���s�(
�T�
T
�IW��=wQx:�S~�b��iO�Fd6ӽ���6?�V H5$�u�5<�>o=�dg�iyQR:y �r�
���ʠ��I�=e��j�]U���l�r��G�?\x����¦�4�3d��[GXM��K�|���z�ֿ���������Q{S�b���-�lt���OxE���;fr�s���%z��/4��#�`V�yp��6"�%]'��H�`J�S'�Ȣ��}�'�$e�&@�u��F����e�{8�����������!��YŇ�I�c��r�蝣��U��ة�C��B�~?�;R�\�D'$��T�ZЀ��q��ô���b��߸��+;��65�Z4�ޤlZFW�3]o�����كJ|_,�-����W)yξ��0���d�L��aH�*V̹�ߛ/]GH��eo/<b��t	,��{��U��P�3+�dTb?�7J��Y��,+(��q������mxx��M���M`&�.a�M�Q���NX�؛��G4�ڡ����U�t���[K�<n'-F���+��y[�G3� �*~��H�4�bj��b_1�M�v'f�6�ܳ�ө�[~�A�����s�Z���-�����C��us�y$�f�3���������T�C� ���`�����d����bU��A�i�����6��*�'[P7k�OC�a2��WȥI��*�M-v_(]9������Q�{��C��-<�F0����K�2yƮJfK�=a�� �Ԑz���aj|��ŸEsk�pLJW�I�:ú��h���
Q�3��ѣ��)P��m�������B��]5�}e
��9��8�.2o���e����*���<�B�K�el��4�;,��S5xv$6�Ʋ%�r��ѫ��XqΕ�z��BW,�8������m/��^&!5�kK	y�o�f����}D}=ݡ�yz�a \q�(+��+z��B7S
�/������O�9���:%"�����wE����L����� ��m!�(h�x'��bQ߷�+�LxwY��*��q�jd�\
t]�,R^i0Kǫ��BGqV��@��_�;r�Zd�0���;�G�ٍ��&�1��Ζ��*�P�U����7�<�.ִ�\4�-��$�%�Au�,�Į�y�m�Nڼl�Sꐇ�ۿJ�P��Zh��@[f��ruZO調�u"�+d��@�2R��m|vs|OX�g�)�Ζ��_&�'�	X"�p"K�S�+��ʖ�>���&��
K���v����z{/֚��x���Vkg���e�{JX:�P���@�~�>��:�r���g�$BFz+�w]>�Tq�ę:)�cq݆r�߿vUTMRZ`�
���K��X�@=to864�q�q`�64��a��|.���gu�0���ߒ+C�;��F�������m����&�/�&�Vhj�7���)������N,����X���g!�eU�'�c����1(%�IɞA����^���8)��YX"��8h�%\��$#;ky��gr�E�f@Ў�ѡ;�N���r����`Un��1'W���~)�^�u�]#m����j����\����)?�\t�q�ʷ��q9U�"�Q���>��GƯ����6����I E*��y���1$��bŝP:}e,%��RJ?sW����e�m���`ydCN!�횸j0�g}q:F�P�2�+�ba� �ߠG��Ml�H���Oq�5�]���#�K����}o�y��k���L��ϓ���P���Yh�Ƴz�PsMД�}��}���4��X�3�x.����C�����;�8�.���3��1I��R��	AJ������/�URd6%B�R�c`U��]�݃����4bk�*[�	� �0U5}frXh#����Z��R�4}�0��^��Yfv��%l���f���L��-[�X�9���Sw�fy�$�TV8��O������MA�ΘQ[�������r��D���_t����~�_��yg)�Yrُ�S��ɹ\H�|/�g�)��%Q����;
39w!]w��ݫ�`(tlW��a}��:�K��Ֆ�,d��DR�%V^�E��G6��Ѳ]C�,���OF��C��ϓ�,U�\�ևz�tQQ�UO��J��ժ16�:cG�
�څct?<�٥;�������ܲ���'a����94�MF�y/JR��m�b���;�/i'S��>��m��H���@)�s�o��<k�lx#[ۊ�H~���9�wɌ<��R���v�6�v��`�F�t�hD`V�#ޯ��h��{��x& �K���ޠQG�o]Gs{��DVu�lX�O�c��f��j�4�+���DЋR�/��T(��n`�􌂚���1��c���7\�-8$k3`~�$x�����*����<��ǯ�������_/YϽ7;�tV,�S�,�S����7�;��DϞ��f�:���.�,�v���El�5�\�s�1���
[��2^&�GT@�H[Q
����i��~$�7��}��U�� �0���	�l���'���4�� #�3o�ٛbn
����/%6k��� ��9�R���^p(�c�.���ɽ1>�&Ahovq��?�Xl���$%��0����(�a��$��\~	3<����܂�2�9��R<(�����.դ��uݼZ��H��	�i}���ХA���g*���.�:�鰃
�3��-�E�<@D;I�8j\Ipl
ؗ �m���D]�r���I2���e	�<6�W2RI����D(�O@~���	$3�7t��լ~(`�k����H��K���$۔�jcES�ˌV�6�٢(��۾���..%����\��$���,�#;�ÿ�8�����I��d��p�]t�z8�����{����!���+����E-�ZCq)�*��NWH�խ-B��-�l�&���L�h�r���cdG��
"��m��U2uQ-FB��8>���8���@\�;�>����[�1b������>�����uĳ�q)X��Ʈ��@U� ��/��c�e�L��,e�[W-�����nw�_&Uc��v��MSD5c��uH!3{����_׵��o�f�sY2���Chg�SnȨ��� �E/e��nXy/il���|>(�Or���J����s���,O�'�o_�D8���4ƌ��Ү��9���3�#
l9'u�����$�/��P��C�*���_��m+�9�L�0��
d*����r�[������Ϙٳ܅$mGz��d��׺ߜi)�7X�n�x��.K?v�S�߳c�zH�@��6.X5��K�}(��:�D%��]4��D�v��5�i��3���I	�$��)���4�fp�h���HL#�s���_�ܬ1;���C���@�奿x��8��G�N��x�G��Y��XJ����dt��*2�[���,z���UW�����ŉ��\��R�*� U�k!~�6w2�����,����	݈�n�Q݇��!���*'�_=��i��.-࿫�r�=_
/4{ha�����u'��9��U���p�:���db�.��]�ˢ���Y��2AH;	B:I�����w,���}�������R�J:t���՞��@,�!\u*DP�0���١Cj�0i�G�i�R�Kc�pE��H��{�z�-�I���Se���F�%UA��0��=� ��\J
X۳K�:��x�:^��O��MV	�t��M����	�0qAL���[R��t|����'�I�%�!���*��S��U��^�(}��I��시��Y8�ޕ��x[u����\��-k�����7�J22+���L%��	�x��%�l�_c�Э�Y�����x��P2,Z�-���qrV�XxŽm#���(n]�@��,�����B��=�h (C�FYƿ�DO��8�Mo�6�Z�Q#���	ZL����=C�Tr�H�R'h�c��X�Lxs������Lr�6R�+��6��}84�cGD�55٤D�W�Ya�l��4<J��b^D���u/�dm�H@�Cw߻oE��P���ԃ2D��vݾ�=)e�ט�'�5O]W��^��ș�C��k�zÆĥ�I�z?pD��#'�!R����}U�����!IѠl���&�P�]iw5x�갚��A6���Cf]��(�¯����H���C\xڞAh�a�PPJˀ�w���3����[�O��>3Z��$����wN��C�,��⼈z�!��#�Щ��;��'{9B�>31�"��؅�z�oGw�.dW��ǩe`p�!�P�FTLC�p����1t�O���K���+6���F�77�u�#ϽQ.�9eM�ȘC���kD���3 DPM���q�{�Q��W!�+v '���L�L��W���:JFO�1̱�<ݫg�Z�m_��?qdb1�ʺ�;VC��X@����^I�j��S���e��;=_�W�p�ܑ��ZH�cc~_�R�W�⮫}KU�|~�G[�_.Ƚ���s����O��RK�*m����L~��;�EXP��cv>1�Zc8�_]�In�^�����R�#����̜mc�+h0���z!i��1�JF25\��,
=�c�; 4�q�O|�ri[�Z+G����>]�����m1��"!.]=�i�������)��YP�z
,��^^h0�� �'R�}�BT��;�<�t����(�k��d��~&���)*�4�B1��̉�"lH#!�n ,� 
KS_;�O6��;>�Y*IH�^t�|�Ӌ����V�+e�?���]�0�W��X�?<薙�a3�ί����|ה��c�y;��UT��\�Xe�pV�R�?�RH��х`f�^f����ꆣ���;�Ai"3���#k���^�o�Ȓ���f�ە���a�ν�K�q���Շ�r��LǙ�|<�1 �-$8J��E�\t�RI���}?�Xs���g�衛� =��%	*,�����B:�rj����DZ���1sYK��(Q$��]��� m܈o��������;x��K��֧�{�_�Ra�ŸB��ݨHD�n�U������7�%�m��܀�"����dRT�m�A�������/�T���O0��%�d��vX�C����;�ʞ�&ܢcq��Cc���յ�,�gǠ<͌�M6�lyM2�1i��?��a"m�6T$}4wgq�%\���¬��rZ��|����9��ƚ�s�4��vİ�f���o�Q����Z�ܶ]����d���jh����sѴa�*�][k1��}@�쫠(7�&k;�NK��J���U���n���j�Vz����Ǖ@����G���ݽ
����z�p���#�d��WQ���FPj�K7��X�|�����1Ч�ڪW4���A�=�"�=(u,�] ÒG�	�Fb:�F�.����=�E�NIE;w�*Aih%A�K�y�t��L�҅Y'�p����$��@�-?��Jp���o��Gѳ��@��M5�r������KBfs����{آ���@rȪ�I�t滿�8�/(W��{h�� aJ�]g��ҭ��I����6���,��qU����,�c��hZ/f��s��EE�'���B��'i�ak|�^ʻ��BڧN�A:,ͣ�/#���d�S*]���cJ��g�m_�=��3�ŋ�N�(�S��Ƚ%}hf5�8]�P�EK�C��� ��*�JDYE�S�]�l�^���Q�s�_U�^8
BX�e1��hA���u���������Z���]��Ƅ�"�w���̛J�d|��%~�GFY�҉/���]&v�p2:&=-��2���0Q�$ o�p�3��s4z7-�a{�ɼi'�+�*�L^`z~��*��!�^L��\�+bkݷL���^^�p�����K�
ZxQ��=,�p�բ��J�촧ݏ�P��D)��貝��ĩ�I���t�5�j261���J�+��QV�L����m�����.*/��ۗvOp7�F�t� ���S*s����M;��R���`�q�^X3��:����4���h�/\kr�l��DН�ʩq����i%W>�{Ri���u�v�������᠄Y�k�R��bM{�@�����\^�̬�ڰ ��yf���P�&I�c	 ���������p�fkyt�w-Q7yS����@G��EYԺ��O$�-Y��b��=�hLH��m�H�f�� �0���e��y�]j4�������f��:'gL56�q?z��>*��lY몝�����	{�3���4�&?P�3V�i�=�+z�Z�x1�5��Kz`�hC�&�JxA��Dx8p���	���{�1����V���:���)HJG�yD�k$�$�hzm�k]���8��UY�~��^
_ݏ�ԋ�H�0G�9�>����5{��	?:3�$]P�h猯bۼ"E��3`�e�Ț�ѫ�����H����p4�G��*��7)_uCO;��ɉ�py��a�����n�"�G��j�|�J|�T&G�WD���z�#<%�"�#c{�@�B��+�XbM��~p��KJh`:2���K��`��{���''I8�Q�Ê�:�o^�\:F�`���c��nUಆ4��Qv:m4� �/��U.��-p�k|T���g�ܼW�p�:L�i�l�`x8T�K`�|W�}ޗE�=���~y��Z��tu/�su8ǯPWm�Q��c�޶�漏쵍���E���R�ԧu�AH�r�����:;FϸR��$����q��n�R�5���9��ýFc*�$Ug(5�4d�M&����@H�L��1՘���1m��K���Mbi�'g�E�]�FG)�ΚW�:5�_�A%��'�E�ۡ����FBt�]��5��MO߻�(���n8-;�V��S, �6��晩�UD5���w��iW��^k�Y:u�k�
��P�,Xǐ����]������r�a��h�s��g�a9h;w�@XAE"̬�j�E���K���24|�mY���&�n�.����� �R(����9{>�L�F* R��7+|/����1�T��yr�
"��k�U�a7+�>L���<�A�cb�C��������O���?��eJ�o�2凳� ^v��CV����nLPZQ�<M9�]YI��J�\!<�aKϦ1�-uB��[�
�"���cn����>�o۟=dG�챊�v�b��Ѷ�M=��M�%�K%,�d.�w�ݎ���M��B����������}�=��� ��������/��q��<��M�k�w�Ɩ�ܮ߆�O�pP�tu�+��E.q�O$'n���v\~/ѡ�f7����^ljTp��<����e�@�իN�7�3�
���w;���f�b���j��.�-$x��]<���y��nuѥF��P��C�($�V��upj2�n'��!`i�##,��>)��/�E�ȕ�V�X�(Yt0/���> u�90Q���_� �B�|x�d�G���"~�����|狝e6d�#~S�~lZ��n��ͧ	��?D���*���IΣ�eP&o��b�<Z{pƢ��{Z�,��+)�,G9JB��L�J��3��7��dAH��`_������}D��4@�Hu \G�K(�s��, �b�����E^>�ŉ���W�����vB��`TNB�sw��8w�B�m�&B`�	������۴��7�j��8�n�$��ZY��S�C[��?��9'�����(�_%7�� ��g�T���*�%�尿�IN8�|���7R?׷s�m�)B���N�#��7�0�)�r�ǀ�B�� �k>6j�H�~��J��D�%55��:�e��=�.�mՅ6û��lC^��w]�a��g���N�B6�֚� gב�.%Fσ#��̬�u�����/{�b�	��}K��,�����OO$V����q3�yg�4�E��񡀤����+|�-�+�{7�O�\��ᶝ*���)FX��N�16��܎��4"�xP�P�>�_���s5š�����W�+.�.�n8a���J��.�*��oh�;sB%�)�U8��P�G`��Dw��܊�8 l����{�f<��s�^���3��]�c� o�0�|8��{t��p�t1��4�p[j�n\6��hveo����c�?��1�|b�|ԁu9�W��� �
!��`��Fqǟ;~��}}�1b�&uߖ��h�ٍ�"E6Y�ez��-�J�Z��[�1����hEL~f��Bf���3�v��^k]��)�;i$"��U�H���&�Ԯp��P5�VE�'���<�<Ј zBs ��ؗ�����Ͻ	��}�q��t�Ĥ�Vοz��@'�E�e,��FO{M�p�B�#2�^��9����݋���6�ձ�{��i&�vmO"�S����#�Wհ��03hw���������T� ē�?FB����O���qO��N�E4`��B�?��|.�}r��"BZ��^��zhS����=㭝��I�a,ZT�P��K�?+d���̪���[�롴����ƺ-*6��Q�E�����l�i�o���x�ji�6n��(�ty���O�D#0��x�[�H�i@��)m��G�ĺd����3�A:��ht���^�;	"U�Ֆ�i��o�3F�le�s�+�x<�+P�b��(���'RQ��Q��y�n1��. �>�j콶ay�����B;Y7l�3�H�b���˱�y��N���ys%'�g���?=C]p�GI�V-#dp�/�^Md�@B�| B���h&��C���䌟�5m��%��+���>4�ThV��n�[,��c�Q�W��,ٔ��ۜ���-�2�+��P5.O��t{	�����
A5��׏��l`x9��>q��v*���J|"��s|����{��^��D��t��+��Ǩ��@V�\ FL9m��+Qk��QČ��7.�vW�Y~R�s򲅙�^<#�y]���=S���'�!�A@� iUY�'ɥ�P�  Bv�fal}�p)�g�[��ȂIyb;�Q�yħmk���`�zd�CIB�1���K����	�����+c.&֢�./��%�$5�"�����3R�*���[1v�L�[E�3Pwd�Q�W
n�`�L�q)��J�|�+�[C=}1��	��.E�:��mOl���30����+�RRY`i�,��Y�-T&�m+����;	���9�T!~��<���Ds�p�:�F����5L=D�zE[J���-[������������:o��l�	u�"$�Ls�ұ�%S�W��W����Q����Y.���GV>���3��j�:c�%>iI~~�P�.߳Q���[�ʈU���C^�6o���[3������"��J�`�ڇ �������` �IGKG�_���R�I�c���N��j�����f�L	��y�|֪~{h����ty�K�W<
�嫵;%�>�<h��3y���zO���=x��v������{��Id�*��qE�����;�`��7cZ��-CF���2��ao�I�v�W�����!ܕ F%�S�y��x%���ǹ��py����}�~)�R0�[a�����c�ȣ^ݡր��'G�t0zȩ�4�`�y������xe�Z �)]�İe�<����DK��J#)u<����+�������W�u�����U��i��k�C�.�^$�4��.ݪA
lT˥��r���ށp!m�|�Μ6m��d����1�ެ7M��@�2{XA��8�;����v2\2����w�Л�!��n~]���TS��b�>��N�mE���;2з�rb��qSѡ�\�M�ՑU����孫×�,�e��^fK\���i�fZ\^.l:�H&V�HB�rԑ�|BѮw���kA�E�)*���4��ު�#�����Y�Gƌ����%+�vn͟�5$�1!��?XVS���֋{��J�:qJ�AYz���E*.K��Z��.)p2��P��Ҁ=�������4�-gd�	Ӛ�_�����nN�{]������+t���l��2|]��L0	VX��8. �G&�I=�JQ�g���#�KJu�E�~r36���hM����۔0\!�&^I�m+�-#��0��6me�:�i�,�s�g/I��j8ox+����$�p�͎�"�v\R�8�M'ݵ�>R0	�9s��i)D�m�S6X�K� �~{�x�li��uB5��.̳Le���d̊�l84�J�*�݊�$]�-��B��hF8&U=�+m��|�ś�UY�z{~In����R8}�sV��р4K
���W� zl�p�v�G}�lN�����[���v��H�֞�(��9����(�e�(6� @��X���
X9��.����!�ԎV�fD��P�a���h��i��#Y�H���W��$��\Q�ŏ�9%	��3�T��}12:
!i��E�a�-�����"X�e&Ӷ'���r�[tr�&`�Zx��	�E�{j�)�$+�Yu�.�9I��I�d�Z8�����烖�����.��MW��Z���۹�/�j~%�?�4ʠg�=��}��W��휉R�	<�@��u\F"3T���ϐ�͖x�zt��C���b���߁L1�o�F&9{��8�1BC���t�'.���c�]�FOt��[*)U8}C���v��E�~�?��=��h�@�e?���`��"q�0_8�~���iO@ �y�֢RPŎ�2*�����2.�^>Z.��_w���qL� �%q��XT�t�7ڛ\eў���/N�EqS(�d�U;9NJ���� �u#�k��Ν��_�&�B�� �,��>�<΢$ѹA��)X뙚ذ��4�� ��,�"sD��8ٯ�HP#ǥi	+�M*�ޅ�6����T��I��.�	��$�z1 k^�D��K'�vkOdn�ZW��(���R���6�A�AR^{	���٨caC��K�`=QD�V!���l��Ի�r@-�uQ��gJ�l��[�L+�p`�L��C���*'X� ���h���=M�54+$F�IΕ�J�Z:l�[�}��������w�ױJ:Ͽ\U\���\��*�b,�W�͕19XmI��:�(���3Fp.J���*1��/�6Dħ�
���>З�&u�Q�V}f"t�~��H+�x@�ϥ,��������O�n���-TM�}�8�V�ev���pq?+�+Bǟ�T��������\m�{N��Qa��'~��,�g|��s�*���z8����J��f�S
�>�s�~�o����t�S9����᤻dH��v��jK}\6�R��LK
�a?�m0�b�!���;��r���,����.R��:X�A���M9�Hft��Y
E�C՗�i��!g;���wTR髖+f�2�����G4�+� ����(����8���=$ګj
8����Eݹ�|?Y� <��G��:�������n��Q�S��^)��²A6�5�g1�>i���%-�o�f:�����|h#=�isr��֔�ŷ��hSc�9&�6�{�%S>K���_mAi�2%��dw�w$��ƛi�6��y,c��Ii����0@��ԀK�iNtj`��X&˨�O��#.>��UbK�>�U���u�ZU4�-ć�u{̎��ٛ��.������)-ô,?�#:	B����|�-r)+�b�e�.<G�PY6��ig������]�kH<N�#+��s��ף�@��5�?^�r���,�%j�� ���ӠI 鬐�+Q)I_�*�����D �	nNM"��n�X�N
Ćf[�{,�6WO��C2�Â��6��߮~�baݽxŴl
�03l�-
��%��s�����Aق��r}ԥ��S������:j�e�݁��6��-���
i��
W��ZR��*@�)�R�N#�$��/ł]�â� �an� ���3���HPk��~�D�\�AZ��&�^�c����NW�r��m=��7el��n@�����{7/������/}�Z�wq,\]�*�����&���wڞ}�g�%�\Ow����i��In?��޵�J~����cK|(1b[:��-��?�G���FWPc�@$�G�����������c���6�ɋ����5� .�E��A_�-���T��Z�`#{l�&�DB���BvJw{c�����U���
��p���y�|��x"3R/h���U3���S!�Ù5w�)�pt��u��0�$�3����u�P�K���eo|��{o�Τ�0���cS��Q��>�!�=642�x�*�4�޵'�s�����\� ����a�"`�yt��,q�īi) }N�~6�Z�����
{P't��ԗn�rs��O��Xm��+����1U��U���Bb3b<���'��䉃E�l�����V�b�BB�d�I���)��{�	wڽ��қS��\�墘��W�8�>��V�~�>�^���Q2���2;�	FB�'�����f)�|Ǌ�3�
/M��B`H����nZ,��=��	��u匙sM���]��7C��z���>��<@IAvY�fM��#�Kx�����v�o0��;~�]1��E�%��1_,�I5�vs��U߽��J�=�&0�s�g�V�˂��n�Fu�q�t�%	/ڄ��B�����7dBU����N?�����Vj�L�]t��(A �R�g�����-�26�.��E����]�3d��df��޴�Cɖ�X��[J:@��p�)�4/=�N��\���ȿ?!�N��Mo:��1�PH�9q� �k�ӭ�F�!��/�� *��q���Wҩ�#hpқkCD�
��$c��5'A��j�/�������Ш^�:���\��f�F,�N��k҈�q�d�(
z����K���mn-���&����עp��|A<-FxG���8��ߛ�P����R�귀
�Ǝ���?ٛ�0iccm9w7��*d����X�%��U���M��������ϦA��8@�-Lש���eݫhDEw��d�c*�d�m��a�Vy̴T�y-zk^��/i4g�>��H;��`؈�ks����������G���G!�#�+;�����Gr�~�Ϭ�㸎^�,����#��;H�ʀ\�Mr0Hjc�F�zU���[z@�h^rВ��eO��+�3�}t���HU�r��J
���I4�@��
���uѺ,a���]���;O�R/5@)�\?�����TR�:�}�)�jK���$\W܅��U4D��ӧ}7��@���t|_>%$ �ݔ�Ʈu1BV)���d}�[���@�D͹�%N���7�<.�CK��� H�P�$BNv
�ũ����g}�ڎ��8��L͚@��]�X��#W�D<\�r���n��K6t�˰$���an�o�#w�!����ߍ�EDz=
&�U�G�9��E~�ɩ��������&Ps�T���A)Tie5�:�%�U&{���^��َ����B#�+T�ܽ�/�`�9��e�L0hI��1�l0ʏ"˃��G+�O>:{�H�OQ%ΧW�ˬ��ʨ9��PH�����މa+=f����Hb|�|��
�ܐ@S/���#�u�"�e�ol%k���������,r��}�A��Ba�A��F������:�ڇ����&���zcb?ج��O0Vq�U�F�)������͵�w��*O�V��y�	�� �����m��C�@T�0�|��b�� ��T�}�&?������Ř�g�E�-�>"����e�@!`�<��h����Ke��)F�	)>Z^]\���W��)�W�K|$i-�FwJ���[����/�i��5��w@�P^����ܠ9�8��������R�ĝ6�
h�����g����au��E�⏄Eဉ�B@�(���C���'�jH����sDR_���u��m�#�N�8��Tѩ�M��Sv|�ƍ��Q�S��M#� [�T�^)��f��
��^���f/X�&��l{0j#�46oA����<g�����, 񴐶�<Y9�A}�ҧB��7���7���������^Qέǫ�PP����e4|�s:�Jӯ"8&�!��"Y��Uu�|A�	�r.�2���ƩI6$���=r��03$�r��g��z��v-w
�E��&�Bތ�ǒ�!�V��A�p�{�ӏ7��:���W���ґ�j;|�=�;a���_�g�G����,�{�c(�-��[��1�]^ݬnW8�>�iQ�&H�!�xN���팿Gu�Z�o����<.	�6ę��ߥ���ϔĔ��PZ+),@�k�=������q���\��M�H�jo��ۺr饎�{��*����|'ie�㐂���X~N�	�nWec�2�6��O �`��Cĵ�E�ج]��Q6ņu���D���7x^|����q;��T�п�I��He�(1��\X���ai-��m�-R��z��;+�s�ݼT�@����"��2�_�E!6�5��Z����$�ތW�PE�U��~�oj��jk7�������=��#�K�c�6dL�KQSÔ���}d�V���?[���G�?��=n+���]8Y��<�\�#,B����S4��t)9k��J����t橸��Ԉ��0B�b�+�x�I�6q�����)C$ �c+�EB+�j��\o>{���Ft:o��-���O��k�D#�x)X���
�z%�Lt�|������Q� ��������x����d���7�����
>��l�櫯��zn�h�}.�chW�m�4'y�!��&cTqX�p�j۱3;F��}�?���@ɾ�*�$����
Ra�M��<s�u�櫔e�g��լ����]��{> ���b�;���s�>���5(���p�:t�I5��T+�yˮ�0�S��8��4��,N��s�IM�Q�-@z��2�k����h�:e�237���{LA�ʢ� |�8�k�zq������}�ȿ ��Ea&��mn��V�c�Xڡ�kOΊ��A]_��F|���4m���~�����H!=���
�}��#䄈	�6jH<�z�|n������\	�6�m:��t�=ڐ��iCG�WE��^�u;�a�:�w�oDU��\�
�-(��'�����g� 
��-��8��rR���sހ��3�<���� �;��@��dK��14vʆ��Ճ��D��̭��E�'���F�a�5עӶ�dRI���B���*�70޾����;%ˋ&��)���g���<��LS�{���I��,���������"ƛ�4h����z���y'xj�ĭ�����S2(�M�k�dc�e�6��l]�z�����Ap����(o����1�Q�>&z��م��L&��{5g��9�=�#��:�6�m�Է�a]$a��Y���Pj���[Z���l�N���2��9q���:�{�K���Q���4;��T�^�
a6�L��n&�$�H��B��1�M�I����l���0?���CɦÍ0j5��$�Z���aʞ`��Oŕ���������S��=U�G4nWi �ۍ�-�k�$9�T*����j���Olm58�1t�;Y-�TƔ�Q��109�f�Õ~(�ي���~�ah0)���%�R��LX~C��N�M���6��@��h�k�6p]�*kc��ܣg��B7�zT�~�=��cU��� �?�o��~] ���R��Sqv:Ǚ7K����0di�b�O-xq�|i{��#$ь
妰��m��7�U�%OH��,�e(��VRZ�J��%�4�{q�+RO���b�-7��S�Nƕ��T�(�����O����L�Ӆ
D����H�G� �c��B�#mc�`��EB�0j��^?��,=A������)�	o������	���ۅ�y�*z���f���=����2Y����BY%W��[c/�j馂jN!'� K�l*���n�Q��S��*��Tޗ������eX��z��s�b��w)g�!�9r�冷�Z�M�ә��������U;"�7������ 7'�^�df�s@�4�����ί!i�V]A�Ҿ(��	��,k{UL��o/�mg��tAexX��Iӑ �*&��ղ�^Ge��r����s��Tt���O|=q˭<,�!�PL���er^ �U:ok{ �e�������@\��:4�x�Ƌ��-�uP7p���,�5��Cf=f�Υ@?��=ڷ�њ8F*p�Qz�߬�`a���	;����= f�Ń|&"��0fd�/��%w�i~XE�V����<�_׋��Q�甁JI~z]�s1$�h���EYq3d@]3��8� \/r)��}e���F�#B�� �A�Q������ !-�E<��K�u��!�'�aT=�K��e�j�j����@��7�櫓f���Ͳ2�G6&E`�V��[���PQ���U�0�n�c�+�ڢ�@�3K���.�"��D��=h1�4�>�!r+���۲(4O�!�d�<G�~yȨ�_���
��L*uҐ)��`����AN��f�5 ��.zT5���묱��cܸ���0�Q�HL%���'~��0o�C�-:�j=2L��B��(���B瑺+�:�.LYm��ЦV�q�������8^�҅���0����m���;�x3X(M�
{V�6�b�K�O�f��3d�fo�ί�Ior��%-�܅!�=&�Q�E7T�3�#8Ɋ��Rz���q��������$6���O@�V)�7��K�;q��Ͱ�
��j�UJo�����$j"�0���nR2�V�>0� �^�S[*kY�Bw�>��I�Gjп_� #��i��(�L�r���#�iw�bʭ�\����:t�W�N\dt� ��A@�P��$im����^~��ER+ɶ݇��v�)�5��DlO��+��i�Sq�F�쵆4�W��/Z{�"�B Tt�=.!���2����oK�_��Fh ���Ji�sy�&Y���y��y�ߚUJq�Y�6�.���E@���eC�n����ґ����k	'�3E��-H�,���)"ɑ�W�F�s
Ч�tO7�a��H;t���<���6-@o��_�(Q_J||N��@�=�>N~�q0�Z��Aoi��țI���M�)n�Pکv�3�����؉+�ys����G�j�L��F�u���x#�����H���r�����}�p�R1��GW�zV4��"LC�gm0����f��_�x/������t��
oTa�U�f9�&P�-�*������_�c?yK��.o�bXQ3|��T�tVMFì��Tp�pZ��&-�I����{d������yc[!�Q�����e����chu?�.����F=U	o�C#���8o�s�#J5�Uv��V��\Y�CG6�X���0�{����.�
������?-�Z�iK�〔��xebO�8R��k������,�E���i��$�����h?:S�T\���t7Rʨ^�!%Ud��=2�=�~+�45���k?vPeީ��'�RT����JrX-iئz(S������� �)�d1�
�M�/��ب��@e���]<dW(E�{�P�Kr���O�aG:/7<np�	���\\~��C�n���
9Q�"E9��I�鞨W����T
G��)ޏ�@��V}���t�z�/�c�6��S,CHh�������k�8�7�]O�wl0�_u2Ж���N���Ս�l�G-��a�������18f����ŇySG�?͹|E��a㭃Y�C�6QbJ��(�Ǵ�}ݱ�ǂNBn#�e�7wjdr��q�3�ѐ{NDm�׺Q�%O���jZ�����݅d˧����vF��h�jO�/���E�	N�Mwz��+���2A�TeiA&^0�(�"�'6txC��S 셈��F.��1G@��Zi�ϵbe���+����m&� �{�T9�Թ H�,C��C�Ƹ>*g�b��bԽ�6Io���5�qMY�Uk�˄V���!�(�DR�gc�d�OTy����]�L~ҿ!�P���%�in��g��K�|��el��G�d0����L&�J3 ɂ���!jFG\F�r-����u"��[ {fr2p��`����UA���;�i�w��~?${�Ak���!�ޫN�C�X;y�4�N^�D�9���O�]�F%#��bMw�q�}h!Չp�|֯n�\%��~Z1FKhM��8j��:�������/�����۫�~s�Y�[\��2�	9Z������(:�[s����_�4�%��y�d�a���|[*P�c���������[�ny�z���ea�ݍ~S�~�k�d�
1�ȎhK�)����Z�`I���b,��dZ1��3#�1��?]�+����Z�͍�4��,��^il����u�Ӊ�C�XsJoB�W�ei_�P^���I��	=��)"�
���n��cg�X��O+N�o�6Ԧ����y�H�meb�HC��I��T�� ��J��э��4�1����[��d@Lgl	�iȹ��)�
ᫍ�a^5��99K�ؽ��ʏ�"(o�#���[��q�\~�pY�V3�?� �#�Ӳ����3䴿\�Κ+1~��6��7���(-���`���FE�͸+C�%{��_8?�=F���W�!,>޼�#̱EL���r�|r��_�F/�G�KC\�������*3�+bЁ����5?�T��7-xȜi��N;�X�Y���
% t�N��1Ҭ�q�Vn��u���7�ߊvQ�q��O�	5�T��.۝?�`��I���yqӯg:U6����R=c2�ټ��t�YE�*%�U��i)%R���ˑW��R���[�U��E5^S���Ş�4�Ͷ�qq$4}21�?1:LTJ�B�Щ�:��J����:t6w�*}t}�P(O���P%�B��)>�+�T�'\�V	A��^�x�kD���?����|Z"�~�����ű��O�z{](W�Qs�H;I�f.�ƭ#�͑�r��.�=��X�s�~$�F�u�;�Ǘ.�:�b�E���,�t'F�~O���8ΙB6-��y\Ȗ5jr�ͳ���_����j��^@�`��e&1��,��.�\~��܈�x����yh��f�N����Y�>��e������%|�*n��Q����\�x�X\����mM)>�:JV����k�N��cӮ�!$1g4�%%S/xE�����x���Uul�741Bh	��C�R��g�g��W}����I���v:N �ٮp���v[�q4��3*�éGq��� ��Q� L����o��m�:BS{O��]��w�ϟꢕ,[ ,uf���se�^+�{)�ЧZ��7N��-�f�.���Ys�e�i���/�-IO �#��S�!���Z�����wɁ��>���h�;3���i<���T'7M)R�<I��t\wY�%��9�Y*��>�k���{XF�	�l�y�y�OV�$&$��߸�'�����V���dO/9#n󝐓0�\�}�('��fN�&��Ob۫����Qʼ�~	�pj?��Î:ô�?>c5�r#n��NT�Sv��4�u����R�Y[�ƾ�>��`%:���m84g@�x(�����Uj�;{�5��^�{p<�o�إ\I�nP\�Ʋj!���L��)����Q���q_�R&�e���Q8��hc��Lh�?q���1>�b�O<#��$���*u\���sm�-s��B�5T�[��Z12`~���*Ls�Җ���9������\\�w[�����Ξ�"��L�LJ���J����<���� M6Zy��e�����6(uQw�����18��c�.�u��ZA�c(��nӪ�Bj��)�0ˌ-?u��2W�.zC��݌�c�ٳ����i�3A;ժ�mCp��k�j�F@�s�$��Է݀��v~sQ�4jk�6��~�-FGH��\W��."Ep�9��f(��]u�rX���	�\�p ���Q=�W�s��Kw_W�7=�qn����©��u%�(1R,oKr%��^����΂ǎ���e��@u��xC�H0ƾ�A�#���X��q)g5�|��a�Q1@{e��:�jua&s�w�+��Z{��ad����V���!d��c�=!�\)_�0<��[�����FE�k�n�?�!���`�[/�牖���6�X��uV ���ji(یusO^�b��v9yW+� ˈr��<�!)�\6_��ծ�	�#�Ќݰ�tI��7�Ò-�-q6X�{gv[4�W�zs�QT�����S�W���{C_:2��Vq?�
��t���D�%�6��4��`��[
����OdW�(h-׾�J%d��ڽa����d�q/�
9��-N͉��⫢unD��o�lm@�$�~ZC�w��f]8K�i����8a��G^D��B9([�h)z�ś��Cxv�hn�M�7�ׅ�����\���v-��_��h�[���9)F����#��)���3��s���t��<_mǶ d ��[�-�za���ۡ?p �f��~ �H��6"�'�V��.��k�yJ�ԃ)c�$��"�~�������@A��x63��Ҡ\t�j�B�C`L���>��gB��yr3�aY߂��n�@٠��a� ]J�&s����e?��m��6}R{	�&ݨFݦ:��@)�g�*�r^/���+���6�lm�j���vC񘤡��֡�21.�6T�K���6�6���+�
�*�R��kmchO7��$u���Z�W��֨�2R�o�6e�z�2�*��&�-�$"��VaM��1����0F�4�!9��ِ�������|.�*��Y�=��ІX��M��6��=&�T��U ������8���
�4��o=<�G=�v���I$v1C�(�`zٜ�̚�^ >��CGk�]�.���-/�zU6�sc�Z�4F�6�zXc�D�au'!,�e�0��������C�%��h�� 7x���4�< aM�=���b���ߊ����s�4�/L�TuLer6?����״I�po^�{�QQ�9��cõQ��j�J�qD�����0�x��t�|h��	�oA̺k��itŐM:8��S�����񳾺�Q�V�H;	�S��C}4���^���*27��% �J���,q�H�;�E� ���fC~��)�ڮ��5m|p������� �{��Qrs���CZQxl(�6��M��o�O����O .������eSz$�;�fͦH��<����`lF�G��ǒ�XW����Q�瀥�Q��d->Ǯ�+��4������u�	�!I�Tf���=������n"*��^���L�4W�6O!=�5G/D�l[}���39
�3����k�����W1#��/��8Ա�� o� �������N�
�4��!�����9���)�)N�%��Ȕ6�~��#�5��_Cp����{��jb=$�2{�yo�&%�T��Λ�'aY��PF����#T���1�p��~�"5�b�r�Z��0&����}!�Y��~�P/�e;�d��P�ͻ-]����z&ۡo��&D'���YW������9q�I-�@e$��)��ӕ��߳��C�E�u3E��:`�O��@Ǡ��,�
=�ϩzN}$�9M���0�����A����`��B��'e�y�*4��e_yn�5kIAp4f;D�I��wn=���SPՑ�aR�FQJ�Z�W��/C��P�Ew�W��Aݵ+t�+�\A0*O�Dh�-���H�ޭ���c�D�ATF�����V9��W����k�0���1r�������Ơ6�W��?M$(�b�2w� T�����7O�Ʒ%{��z>,��m���%L|��,G_��t�|'t�rBܢ���`�Z�|{ �1^ܙ����EȆ���)' ���9}c�;�SO��dˡgXyk��x��,j��V~�e� ����W�>�<�7��U�f5��9/\�V{/��M]3�p�'��m�O��Uz�^�����LY=6��c[���x���2%���-�\s����+@�^x�4�,��,�����-�h�7[�DYciNQ��񰧼�®��+�_�.�o�b���{�衤,}�YZ�}���ч��P�v*O�A�V/%���r�pof[�w?"$�KQF�j�R�*���R�d�%)9@=���m���߾��U��a�FPǚ�ؑ����o����4="��
-�˫��* ,��_ǖ�C�|�,�H�� ��!:��0i��HD���?����&�^i�4��Ɲ|x��aL�Ȭ����b%��"�o�5�L =:��+B�ݭ���C((9V�]��N�W�,>
_�ݝU����B(����N��Hg螪������EC���H4i�?�@���M\c�<L�ۊj�hƓ"�56<E;�=�Y�E'��>c"���J¹e�y����ѦQ��o���km��>��(�Q��Ů��(F{0Qc������d�5�"�E�<_^���Hkc"?�|@6���PQ�)�h@Z��u�Q�x#԰��~5�j;��M�h@d&g�rp��jY����-q��<�XW$�6"h�KD��%(+"�	�] �e�s�v�&V��*L��e-�hrSQ�hnʖ���u��5�2�>�MycW���dH^�r�cށM��ر�a�Q��ŀ���LM�Ҕ>.Yz<��p��G}&̌������t��&�7 T��m�K�S80V�}=�wC��TK���;�8��ACG��8��)�*�#�ʸ;���#����B�b�T��v��$s�uZ_f������cm�L�x���gl��hA��� �>1��>����I�:�%�#V�$��:8(���}�V,��q'޵e�hvoş��U��b����>��ZX D��)�Ak��Ϋ�$��DV#F�K�#<y�����U{w9�������7ʰ��x�
�w���Y`��5�fTV��>�kln�Y{� ���3��B�������q̼2@�,��,!*uY��WR�Uɺ3jz�Fx�
- q����D�AYP�W�c��8�'�,Qt�V�8q��?���M�d���=Ĵ��ۈ[���%:�ޟc3��Uh��.*8���W6��E�z����H��-���,���K	V
ъ~�L콜�g�dWZ�F����k����&c�]���C@e&#�By���I�Y�ؽ��
ΞV#L���OT�����W\l�h�`x;=�	���e~G$���ya��R�Y�!>R���Y���n�aח.:�jr�7�P<)VP\�T��(+P����:{���7�P�9�z�_��K�4���5�Uv�A�^-�	�G������2b��F� +���$rzT��|�O�b��06.v��[�6����MvT>�'}H�ﺇ*N.?j��o;`���=-�o��b4ɮF�3HFؠ