��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]a5^x7��j�J]�4xB�"�}IS�LrL(����z�1�Z���e�/�����}'�%t����� ��@`޾V�r\�Ɛ�_<xp�%7I��/�V���%��!�@��1���R.�V4[p�o;�ื�6�a�'�ܟ��Јv��9�ם|E5����۠���V:R^175�+3u,y0�.�I�m����&bg���d����%�KPF��Z��8�.N�tDs|�W�ۦ�8a�����E��IH���cY�f�)�����P� z(ǩ�E�0��Z�BJ����t��3.4N�,�.I�A��ػ<���Jat�Gc�ݐF�ݫ)O�da��q���Bn�	E41~S��/~s����`CB@Ts۳a�*s���!��^���7;-"�q���w�@���S�t;ś���K�>6\�A �x����p�V�(�ֳ����@u	a)�(��n]�;�����ZQ9綛CuՌ `����Ԙ��´&\���u�h�Xlu	�f�[Pb�`��Ih������e����+~�����,;�'i�%%|
|�P3�&��mŨ��a )��̒�h��P��)�A,5ˡ"���fUe��d��,�� �� IÌ��9D>�D{I5���Z������C��t�+�L'�.��G���;��_Ŋs%NԾR �E^ʋ�AD�/۪��:�����t:9��O�
p�g�����S�S�6Xy4��M�&~[��K�"XPEϬM2��U5!φ��֋w�#�yE�����HA�˰{�q�'��R���gn<����%��&읒#�f�*�6���y�*>"C���Jm.x�Ï��Q��1�'et�!i�
����%��b=�3�� �-��j����Ǥ>�S�����  ���g�6���0(h"k��uN��A�n�o]�����gD�[M��im�!H��90E�Z�#5(n�g�o�zgS�J�����_̊q${@�V� �r�+���,�i2��
�Ì2�-+��?mƥ�7���gS����5Wl�۾����"z�)��{����\���*
0�ȜMx�F��m����-�лv���v�8!�F�T��z~��b�6�R[����h#1�$���1?�jN���>� �Yp_� ќ� H f3�H���!�V��a@�锷OL�h�q�s�d<�"��I���ca�¬��e��屢x5_'h���뭭>�� !�; N4��r/�g�$�1�ѝ���ň	w�3o�ucW�1�I��������1G�H3����d����W}	����D �����&Ktd�6�R�`��"�k���J�1���]�Ș�]ɮ3T6��1eQv{r�%,���1���	����� R�<~���\��[�,�|�+�E3.���x��$�nzŭ�s5U����i($���/�q��\����ԅK��gʥ�ֺ~ �v�"-�J��r��)l��S$jA�'n�+#���#���@<���0�]yv�����ɿ�3K��T����CUe���&�XPp]�-��s�̇���>�N��S���]�������ȅ!i@-��۬(���o��<���^��f�.k*������t���b��:F1���7�Bس��#b�1K����iȘ�#�S�9a�&��pW���V��`�qۛK9c��UL�������5j�5��;&����xk^�.���x�PyXj��P͆��`�uߌ��<�;���R��9���.?W��'��ʲ)=�w�7j�O<�ja��]N�P�e�5�����-t�&���q�ߵ�*8P(�}.�{b*  ��\%�����/K�$�|yPWC[ϲ�F�0Σ�v�zWoY���D�,ehvo�~��N�lvw���9�}݃ڨ��x����R��췀�n���8k�?�7�]�\�	�1�NVtC"X#�O������a���˘����z$WΆb�J�0���{Q�E�I�!j�w!TH�������9/ 2Mv�Ydg���m�3��7.��U�#��ًȴ��Dꄮ��m��il^�|]}x~Rz5*�|�'_��r`g��Flr2Ԩ]@�L���2��8��!;DQ.^�ܲ�(}��Ҳ	Hm�8O�!�$�ھB�<j1��V���g<
=o(k����}��E��q�iP*.�0C�.s�咙�ylI��I��%�H�����@�B ��8�Ő	�<��viz�G�(�I�ǆ]�������k�Sa�P�;#�'��"Y�&Bڵ
A���q�ѽ�lo���T\���H���2�Ʀ�:�����
9w�0�+����{+��A��A4s���=��I�7�"�C��_uD�ʂ�&��`5��u�^9LVζd��?�{�Rβ�UPUv;��$�3��k�y+qHz�V!�Œ4�OT/���;��9<_+�E��|�ӿ��3�sk��h��r�ls��|\>��Ȍ	�]��
��˟+��|�ף��oi�G�Œ���86�0c(�k��������@���2���0�/8`nz5�T���J	I�Q��/fK�������B]^��-��?ި�
��$E�l��Dh��L�0�_	o!,�R#,�Kg:}#A�/��ߕk�R�nk/`2ٶd;�f�?��2M_^�7�ȋa-CB��L"�)���Xk[A�X�y_��f`@�r���E�e��mT�W��r���d`��k�����I6��R�'i��5m��1xPD�[��@j�����H��(��x�7Q­�3��u7h��NY=�i҆NOB6E���>R�� N��j��¤�����N(��{��� ��|^�wU8,���	Em�j�C߂���4܎?��9�W#M6�#�t���Jא�g!\65e�U+�ћ�6��;�,76�w�@75V�7JI�	>��$�JG��_�q��������xp'$�唢:� ��y�e/ I�Jnq�!�� ��饭p36���
���٤�MH!Y/Ň�f�_z��T�#̟��]�D8-7��+e�ʩi��MJR|��y+�R U	��;r�Vi,H*�1���쁤�Xa������T�gA/�$q���?F���DU���jX>J~h-
{�ј0� � �	ǌ^
�<��ځ̔zr�<�n�����S;��#<�^G�Y7�E�	��ѰC��͸X]���d�zE���ͳ9�Ǩd���o�Wz�G���t��~	3J;���:P�w??��bK��"�H�M+��w	���G"��ʈ���y���d��nT����������-��ć/w�M���$s�M��)�j.�*�Hw},�;5�St��c�=Tҋo��ȓ�A��F��sw��˪���&�-B���@��ls�X����wO�K�����̦�ݺ\ƈ���f�,;�F�m�,��]�	kk_֙��#������w59���B�z`����G���2�|lI�(ͷT(OY(M�`�оmφez4�6��h�;��xѭo1j�m$v�ӭ�@3�����ZE%/^Ig���]K���#�[���\�f��Az�fw�LL���&�r\����O��07�K��H�勉�փ�^>Q�i� �D+2�����}7t[��ۖ� �\i��	�i�gj�R��l��ht�Imp�8[ꙥ9�
B������{�+�;�B�4�+��e�u��8�B)�*���mV%�]��"[���(H���p/�yy��h���fg���'���n�����/��*�v��+�:g��N�G��C�\o4�AYUe�s��sr�Ep�.%�+��m�*�U����`YG��&���.X�/Ƅm�{f��s��2���r�D{+sy�Qb��.YL�qVZ@S	�v��욐��o�B�H�Ȧ�jZn��ך���#�xy������jU
,��)�������;���$~:�'��,%Dܶ��h��z%X�ν��7J�"K5H�QΕ�5�u�1��<
�]Iњ��Yoe�,�1#��?e�����_��^<��)��{V�{�r%qu3K(q��W����~x�c�6������Z��BbyO�p#�:�P�W��(���]mȞ90����c�D��F;\xI7{���&?�1̿���h���J�%^��YL�	��a�fo1�,f���p���ٍ@��3{������̓���l�g�������k�w�k������������l�H� ����w�ؾ��,�JCQ�����}W��
�(YKD��ܕ[��,���Du S�o��:{+�+gڕ��D�rJ�<�rY%����"(�Z
�@	�n4�Ҳ��}㙛�	n����L��]l�d|#��F�T�(���8I�(���~�t�˷�C?����9�o��
ƫ���'8���߿�+��,O�0�� y�1�c�T`m��������:�Af>`U���g�l��и(��V��A)�e����m�@f��D���I	����U�f������ �/hA�A�`K�j���RARzT�YP�Dk�d��W���0�t)G���N��Ƞ���S\��)�\�Aq3a���\��-���ϢvF�!ʋ�=u���+q)H�v�7��+o�����d��V�K�Bzj�I���?]BN7 {��y�FU3���e4x��&����p�����9-`��d& �@oW����$�u�=�a���Xa,	�@Q<���n��_���5����pے�@�B��#��d�u?���.B\c�ڤ�hm�_�ú��AER�Z=
w�1����FW�j�rd��A��5Ǟ��4�6P���mL�or�#�_����BB��"�ui���Y�MΠ9�+��  ���2_3z�)+�.'$<w��e!Ł�ѕ�WO�|���b�awL �kx�.3gap2@G��@�!�r���f/��K/C>/��cqTE����ބ+C�9���Sڛ%��Ѡ�)������P�I?#]E���y+!`��Mŀ}���M��|�D�7�4G1���9)���	��-M�-'�,���W$�����r&a��"i�gh�;�l �Gdº�������W�w����2�>�ԇ3#��Ř��cq/ӡ�����྄mK���ںJŷNJ�nf����i�^��&��3r#,Q�ME��l}b��ǈ��j�]_���x{c��*}���R(�0u�a9v+�i�
q��\.ZF�}����+�6L�҆Z8 餯�p\�vX���ꐕ#�6�wK��ȼ�k:�Ŧ;�UJ_u�+��TƖC<�X��m��r6偀�T��g��۩Fs�)bl^��
C���z��;L�N��Vp�ա鷚r+�eu\�%&x)YV��V�r��B��u�t!ON&Y��M,q~6��?��Rv2ހ��PS�Hۨ��š��ïUF�g�����A�w���v8%��?Z�S�K��;����&�N �SQ	�2A�d,����yKh�!u���K�t���,������_�R#�x�kx�?���G���@C�-�%J����Լ	���d��^�`<�.�eH����nQm��y�P���n݈l�HCPK��(�2�QY8����G&<X��l�����P��7�N��b�)=%�^���Ļ��.�J��cF"�����s2�|�'�$9�J�t^<1��\R��Rk��BF1����/��z鑻������p�'�J��X�m$~�G�Xy�{��gLha���E��B�`f[՛DL��͓5��\VW��aІ8l&������Q2�!!m��%�m9���p���ãeֆ2�@��7����_��~���G2���J��q��Q��%�HG٦k�6�[�`8x,�K���#꧋, 땽�P��]Y5��
����gL��3�Ϊq(!S��x�kC' ��IB�L���x7�NQ�3W���d�HA^�}��j�M��2�n