��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c�Y֢�08)��k:�ث�1��=�1��cO<������9�5�^���W���.�����<��_�sP�x+v^�Y�+(���TOŐ�ܱ*R�8Fa�2*1��k+I�,��K/�$��[�h���Prg�1?S��x�7����yj���Ϊ$m">�i�1�o*L2Md~�(�)/9n�j�߹uԔ7�w�\�;����又�z���QJ�ou��p�1�rl���<�\��~u��}T�g�]m5�8JECU#�ř��B�����M���1�8�i�}U��YΔf�G��5��z_Oi�/��������G[�~�<�06�^�A�ք�U�9S.\A��-2�W��!k�ȱ��<W��JB��F(.G��օ�y���O�D�C~�W�ѥb�&uPmUt������S��9��V�C��M'���8�G���Pz�� mٹB�Q�(�';|���/'�;]�AwW�PN����%皋��a�HN�R���eFXB�x=e	�K�����~ ��o�nw+OS������l��w�}�@������rօq�(\.�v�Qbw�^�oA8yV�h?4��_st�Dq+-��?�����>S�!�$dvtu�qx��c^���;�L���y�Zf����g���Oʣn�Jm�D����ɥ^dbG����Ц��46ϵHQ���3Jmz�.�)F�&��⻫�SC�,����)��t����;��iadH�a'g�L��o��.�K_J�0���%�#�1Wr����ZGC� 3�fǇ����9I�$�&���Ub0:<H�����΃��*Y�F�tb�����۸�(<��pe�aX/�v�|4~�S}�Oo�s����6V�ʲT��2(��J`�;��,u[4��0��r)��X�Ĉp��%�B�6:y\�w�Ѥ����6>d[��" ��P�Ht�P�r����0����X��vO˗Xs���<���!��Ћ+h��6�=]~�9��7�Z0�\�@�C�oJ�x:��:8iS։ӪA����^�4�%�p��/�4��u'���3�H;&���>�Ɲ9�:=���Ϙ�����kz�����Z�b܈���� �fm��<1p�DV�_�^x��h��ڍ/���9� �1���"�}�2��q����S!�Mƾ<��f9 >��q���Ǭ�S'e�h.0Gu���֓xfr}n��L �̂�p׫R��(������)�I�*HԶ_��{}�4��n;���
�Μ�[��~�
������g�D���y�H�Q_��y��Y�O{ ��5��y����^���ZX���6�g���7�9׃ъT9`g9�xt�6 (����t����9�n��Z�n���p9M����o��'��5G���:È7ٙ�NG��*7ٴ���e ������!��"p�|;η%����}\*<����(4�y\1@�;LXQa�1����Se\�mf�֮ \���Ył]!��(0����٨s���e*�LR(l�9	Y�gm�L>h��j`E'0�W։u�%�I�gM��c10/ǫ��lN
I��7��&�l���9�ž�xᔕ��F>�Ah�hL�)�p����dJ�n���]�P�)��s߰+���g��fc��L0���B���?���/�Ga����'�S���nԸ�0�qǁ��﷐T�&�����z�t�\����,N��������x��qEK���U�8��N��b����l*;^�L�|�ZL�Ցi����-�=���W?�e�<f������Ah�4/�5��̄�4���x-��M���2�+�h�	�H`���aR�Gg�B���%�������mcI`�{7���۟�����b�d����w�0w.F�in,����h��o>�}8Z�O��y�/X� ��߆4DJ�����̝��1�5���҅�¬$o�́WL/�"�p=��9ފE٧��N�����">���C��?P*��޿/|B��o�9�z#��%�)��=����_�F@}��UA���X!��q%Ui3�;�G��fEl`r T���a5��Q
�9��c��Ru�קd �l&�'j~�@۩��a��EtC�"q9?���3�-Q82E�UI(;�q��(%q=0�Ս<�I;a�"�J������!�㉑@�d��z�{�>l��ī�0	Y�}`p�t/�^��?�O�e�6���ZQ�EB���/'h��ғB��
ۋ��n~�o��\�jq��v���@uY��X�c��V������Q7˄O�*�M���Vy�!ӹ"�C��C��bJ���%#c�e� 7͆���t5�+5��ER؃b  T"Y�d�xj~,CS���1�R��udD8k�lh�Gk�-���Vrd���z>YW g5�`��$`d���c ����᠘w�_�L0$lҠ�^W�T`�����>N��J��k�04�vQ�IJw͐���柡}�=�&=�>z��윮�� �5fP��TB���͗?�%����4���o$�x$�c��R�ɯn7�~�p��9������� �8�>Q�Օ�r�RuO�e����F3��ry��'o'���(�*)�jt��`^��}꾬�
��Z�kn���v��0���l߱�2��M�oH�0�59-<|.G<���H�8a����Rrn@���i����W��^јo��'C�t}�࠾� &���7;|�*b]��n�}��qa��̘�.k�[�-�B�R<&�A��W�O�}掻Ŭq� A�U�o�R�&ҙ�o��F�>��5��R⭘	J���/��D���A�}�ǐ�}6G@�^��J;n�8"hA;���H���i���#�Cڍ��3��nܸ�n����%@��;N7�H�k��m���j��b}��U5'�S�	$���L�2O������(T
I�䪂��s�n�a���☣�r�X,lォF�w��c��� ��= �1�+ʕt&8Q��1�w���Z�h����5F�lCE�j�ϖ��+���=�{�eܵP�*��m�,W������S@?E���2[�s���l��kNu���d�V�i}_QD��=�XC�q����q�y�J�WgD�o܉K~0�3j��oX{��
nP�)n.l9�6EVV��g�R'˨�!�{�ujp��,>��vб���4'?&\}�)����F~��-����Ga�c<B��{��+=4eh݅?"pJ�8�1�'�QS��^�z���*߽q��є�Y�Y(r��V� ��է��$JhΓ�G�?Ĳd�H`D�%��1��/��m��Š[��I�t�jʱ���w�V��Ɋ&Y�8!Ӽ�0h��Hn2)뎮0B]PF%�����рL�6�k1�� {���[v5�QG�%~���E��������2�/	��*��y�����9�?�x+�U��1�e�s�=|b%�;�i�ɣ��]��k9)�2n/-R-�k�8���{�=a��۬�c{&���a��F&��L
y_l\%"{�\n@���ͧkē�Z�.p}EE戢�+m����" f�ܒ�W����i�b)i*���ߞr��68ѓ��gf��hJ��h�Q#ƛ���{��X��hȖ��P�4m1�.�+�������;V)�L���^-oq�eg/��]/&G���Y�`��m�����ܹ�ɦ=8�S`\-��\_�q"�?��Q���ʙ1�H �����G,���S�Bc�Eֶ�I�"���hP�'CE!�t.ʴ��x�t���^� ��q�pTCp!C9����ݶ��9H������d?e�O�G�<Q��Ө)}��H��cX����������7Gce��X�:g����T���� ��/x29Q:�I$b����˥=U1����Qc��<��0IPp
͢����+���Hm���|R���F�r����5�/���o��=��%�z���X7+���N0�Y�C���3��Zv4Ǚ�Ή�!f�k��F"fo��>f(��2 c~�C���٧R�(�a�z�k��w3#����ɉ �:TI�e�Җ�n��(a=�S6����RMZw�8�e�����28%H�P���p�����si]�Z��B!vO�_�t���$�t�O�QH����3��\�`LT���p7EU��8��t ؼ����Y��пL�N�eN���}�	��?ZG2B~�e���V͚�!�[2��G�����I:�d� h�<����z"n3�ހ,���&�T(,�1R�ƅ�uV�m��?�cM�h�=\��di�%��͕�J�頼��z&�?]���_ �W��>��׃���+n����- 9)�@����L����Ҍ��u2T�#��fk�ڈƀr,J��;�po��f��F6o��=5��y���=S���vt�>������@9�C��̥�����v�H�����6C��B�ġ�n��dpU57>���T$���p�g�r���I������ej��ϸHy��JY2�(�$n8f B��i*�fځ�P t�H�UZSIsW����)4��P��Wec롕���搓u*6��O~0ć�7*�\D��J�gAy��ϊ���9I���N��Q�8]��c����I���CbO��K�a�fw&�/=�V����)Z�U-|�Bkڽ��3�偅���,�H�8O�P��8�P<���H�*�~�������^�07�$�:���j�P�v{�V(Z*H뙝[���{̰���*&M�G�Br�10V�`4�XP�[?N�my |d4ƀL��m�I�ieT��"U��$�vλ?�������g��Itj�`8�"�N��y�u��������*��`S'(aA�,��`��EW-�6Ⲕ�P�~t��ᔉ�:O�6+YH%�3�@�9
%�"��Ǵh��g��4ծ���j�-�H�ʳ)�a'xCZr�5�w����c�(Cl�09t]���qki�^��.��r)�V.P\��l?[����s�[��p�}Y���Cj�7SD��h��p龊���W��i~�����;mA�21������.� ��u\hi��i ��g���.Zi��<�)v�]O��N���?�k�}��B&�B��[��Aߪ�J
S���_�,�6"���H��^"9
B,��qA�ړ��śF�3T=e�y���1�@-	�ӂ/<=^������0��z��-%-m����ywL���w�Ґg���EA��I�S'M���.��yk��r���/ti�~����E#����!����t�����=�LJ}�n�K},�)0�����.W������k,@m�C:�mg�y�g�V��O��c�}�xR�}��2�6
'��Խ�����:I��C4��-/$*x�i^�ŗ�u&vu�)$����rZ��˧�lΛvP!k7?,&'��1@��(>8܀�7�]�8�u�*�3}|K��m��w��]b*�D�1���1�a�iL��D��� N7�������n�Fg��u�\�&
�Em�K�>��r.T���� Rв?�mXFe:P�