��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���Ox���0��?T�}�D�yBl98�锛�l	`�ġ	d}�:��PƸ����~��R��o�K�jV�,R����vy���3����O���Z�����g�̼A��v�{�7
��5�¾����B�C����������r}�:ش)qqa���·����BW�4����"V�CL�zhXo�e��6kT]xl(���%lT'�W���'�N�V#�L�`�`�Xy�6$���:��9I��ì=P��uS�I�w��������F��<��s��y�i�u�����ml�G")�O�4����}�,r��𯴢}�鑪 _@�y�Tkt}��8!�JŜ�>9��C �gl���-����{���Z�*� 9�[�B���c�M�͠�+�G�Yy"TGz_'l��2/;��	^F�/	b2�ܕ�Z���./k7iǶ�>��R nS�}O�i|�y�;�aE��J�V���>��t1S�W�����y�4sr�$�&������
y�VB�Jb�u��22��
S�:~���N3J��H��SV#6;�b�f���p��-Y��N�f�N1]��֜�cU�v��,a1��k*>?]H�ܨ�p�Xm?I�m$0# �4���݃Χ�L�F���,aAJA��((1�^��N&��֣��JL�$�vM7�����*��-޹+(�U�ilV��p/�z*�	������!.�6��M��W��Z�G[��]M�-�v�����{�:��n�rD �h�/�<�䌜����G��U����d}�D<.q_���^��ʍB��y.ޞή�����L4g��W����[��(�b�ݼ<����H������f���$~� ���9X��C������r�3sw*vN�J�Gg���R.����;��١�_�V�7\D?!�9��&$u�v����b�����.����8�Gg�3�H�1.���a�������'�0'�67�.� fn��WsǢ�n�~OJ"u� �R,Ǿ>�]��]�Y�;��L'��r�����Wp�m̐u�1S�D�+�Q�YUB���ߣN�^�8q�
�B�f�Ws��LN���"�}�hi��l�`߷�;$�8c9�!��_�IPZ��w����������_fEHY$�d���B�)�*ꐢ������l�q�kp��&���X��δ;L��.&=%��/�l]�)%�)��]P{�Q�p��WJ �B��:.T��]��̮����I��[���cE��W�1Ӝt����R&	3��O�+\�T�w�lS:�ߣ�umǪ�O)~D���&���@�z��
+Z[�a��h~�(O
V�oW���饽�. ~:DkFZ `F�M���SK�MN��yDc�c�<�J�������փ���JZ2�U�e5��8&��k���;g}�R<J��,�
N��N-(��+�U�]�E�T�_P��%�Otv)	�V�1K���ęn�e�ޜT�&߿iu���R	z\������QUt����"vaB�-�q�ꂟ��աz4bwcK�Ar������Dpk	�$��Mo�8�P")[�M3��;.��7��LN��*�_+�&��(��2�����#�"p�
JD۳:;���$��&@+��*PT}�E��e�ȩm�vz�E&x��wF��7BN��s��mY���9\�y1�W��-�M�qC�\��ND#�p� 4��;$�)�\ ��R@�2��nG��Oê�e��SwEPu(|���[No�	 �[��X-�,�*����V"f�������޿Ŀc�b��oR.�����莴�USh�Bl!��W������-�EGP����a�`�ձ���� �/ +�%���?�i��-f2�E6��W��2k��0(Im2�v�/�~��7��o�9�%t0!�<�:Q��G�a���}S��S|�1tq�ѯ�s���O��wH���k��U��%��V�TL��]��	��\���pU����t��7��ß>��XO�B�U��c���&���R5��@��y�:'�]D,\���;��� BU����$�&�O1E5���O�����p��|�;G����]��guǻ��Ө�R���}������-QLФ���� >������1@	�D�U��a��q|���Ť���L�T�M�}���\z��m�g���]�����kg���"�S[�e ���^� �e�qu֝�M�x�ؠaI�LIڝÍXCt�ߠ?"��O�SF��J�C@���Mn��#r.�l��1�"ۊ�̶����zl\��.���۳F�fB�e*зm�}L��-�EY�%7l�Q��[�����V-��L�=�=��nP���r#�ʕ�Ut�ށ�\(�>�G=�L��N���P�j�Ə��X�i��O۩6����\��;�k|!�5���e^;)6Ǩ��>&M5BD�$9�f���P��s�{�[K��g���x_��Xḥ������{���V�o�7�:��v�t6B;s��Ӕ�F�dX-���&��oa��N|G���,T����b��7�p���G�z͍cש����������T��ֲe��v��U�|��c���3?�Nz2� ���/��OJ-;����V;�M�[�!
�,�
����NT��_1�W'�m;��������Δ�� DL�ݪ�<�Y��lDP��1t�C�CQ�X����UQ�����>	q4��!�<l�w���Fa�ӕ��sbJ/|�'s�V�bD��1=�?����='���ֽ֧��~r&��9@|!h��ʨ�]0h����\�if��=*��7���׉=���ю�6�Q�_��Y��K��D��� ˔M\W����)�ߙ9�o`�<��=��>5)&��D,��X�u#�A��U�e� ���9� 5x�pa�/^t�{?2�[!��B'0ф@�����Yɏ00���!����P�I�_iEV�͜:6捄#�ɿ:�����D�A���U ����0�*�D�N��l;��ՖU��u�0��z�A��f�%}����]�tTaV�4���nw���Z��@<~I��`����*���oA3I1����(D�TL��� |X��h<���Y�<�����$#�
$@����xH!5.kKd���i";#l�@�I�i��u3�8�dME�|�X�� ��".`OЃ�H>CŢ.������a�WfЪ�hIb�A�{f�P�SkK_��|� ⥜z��?)~�
V3��WJv�ڰ�$�N��m���St?n*Ɖ<�/wær.�	Ӽiɪ�Z{��D� bRF&��V��^�sN��a�!�:�/}3	R�N��F���}w4V���v@�2n/�6:�ᔜ7I�qY�	o�6�aE���e����~-@@�+NνvvRk�m����Z�%�hE��Vʲ���J~�r5l��~\
�Ye:t�T�m�� �v8��wn^a�[����=��U��z���&��W�/�H���M{ۙX��ٷ��*�n<DLX�k=VI�YB;m������s+��8_�I+�nV�2@�@Y�dn�:�Z�F��,�5%�%�^�/0�O�B� ��Ʉ����fAt�Pv�畳
�[��H�,lO��7�o�׊g7Ep��A�mPZ��]d^�x���-4�:�
�V�5��e�[7� �')�qcopSk���Q��|�)B�n���R�m���@eW��%�dT$���`���!�:�!R�Pw\s\CN̆�ݞޣ<��b��[���j�0sħ�
&(�!�m���h��󽑞 ����V<���=��!���c|��&F<@t�ϭ=�H�z�������8����ީ��%�R��jbDy2Z9͎����`;υ���-a�q�@GTA�ִ�(î�qIe�wAQ���o�2�.'4ty#@�F�#C�����m9E?��xa-����3�'+0=�b�/.Ɩp;* ������S��\-@h�h�&Z���5��jϧzЯі23#��ܯwɊ\ʉ��������D5-� �EF��$����H�+�^��c�v>{��ɳ|�,^J,��nExc�E:��N��b��]Eb|<lZ�+Y��_���`���A_�ʛ�fs�)wC46qF�n)����υh�Ǘ�]5v���	U�xj�QF���DNw���1�����^�?����v:���P���$�iB7���k2�	`0<Ɛ©�D:l[�=IS:�bIq��v�1l��2)'�,Y�[�u`�~�.�7��6&{���C�;���"ǭ��M�Uʯ�v��Q��D�������˹R������`�/�K���?!#H� ��D6ns�Y���7Wz�Y�3Nj��TR1[XAK���K!_�F'\�ΐ��lt`�[����2\���?��wv~��?��w�@�ش���n&�� f���ڌu/�AΪߞ/U;���V�1�@r��0S�ABWU�3�7�x3�賦D���t�1��V^K��[���q��d������d	�'t~���Y	�:����ް-oXM\��3���H�^p;B�[�m��2/q25lĆ�joO�D��p#��͝Y�A9Y\1�O� b���	[�!��˻��@��*�]e������$���	&O��a��j�N�Zr֜�|�4�����1��?|�{9l��%����_y�i��D�Qј!�V ؖ\�/�Jm޹�J�|`�GneSOY��
GJOA1Pc%$!ޚS����˜4����&�g�Rc��\(��?T�=Kg�98��|e�ՙ.�ę>�0`�і[�m��}W�*5�,$�bd�����~��i�|��n`D ����r
^�y���Cx�b�P��a�20����q�/mC
ST+��2X�,��S���X����DgLa��ܯ�j}@8��ɩ��� �.���Ε��=�TG�S�M��Oi�.�hj�\D�E�墄���+[��dqV]\�4����[��;�q�<��7Y8�>�X�U��m��҉0,:n_��
=͘��\�����[k$6��q�AkX�L��4�#=ݡr��VUq��h�o}���V�-)�x!Ҝ������Ռo�:�ь��ɗ*=�\ޚ���qġ�/I>�tu����Y.���9��J����k�Y���i�ƺh~��C-�M�)�9�ӣ���.�"0�����sN��J2�DL�Rt
����6ұ���I¦������/RL�r�R�o���`AG^U���F�ys6��ɹ�͚l�׬"A&E-m�(��T��ݵQ:T$zx��r��IKɏS�w�B�;G�ks��`C�	�C8 ��M�s���♜TU�}
N\E��&k��#�wz<�Z�q!�='�w��ܬ~/�Ċ���[0���d �5��ֳ���M(���������C��S��vٝ9�e������<w�3��ڈyWK�O��=��ZM��{��S�՚ۼlԝ�?�mu���Dyte��0�t��J��÷~���u2�&��P��O��9S� Jo�J�"�4��c r��`LaS��]�Ak/�T+�Q�\��] Q���|�N�ӛ�q,`za9)���sq�k�6r��o�3ɖj�����^4!lyl��f���he~�9X��p��"Q�Ty�D's٫�a{���a�ro��� ��q��o��ġ�C�po�2B�	y���2tR�q�%����<gI�`opgZF�醝�-�4���g!��L=�~��* #�|4Y�WX/r{x�Ի*�)��������.a��Z�1����֧�m�ϩ�rFR���׉�xR�X0�0OV�J��sY����ev�����[��놐�y�5�FK�;.\B� ������k�X #
���U ����q�3�6��J٣�����rb�J =�L�S�?�,B��9l��)�]$����f������t�����,��3>�i1����;����&+�Inܿ����ͬ�˟�f�t惃�H�rg��S���-r��	�Q�� ���{X��+�i۫8��ޏ����||�۟���Krr��$R��T�P<)e��lȾ�52�lQr�*��<Wy�����Pwي�{����It$�6;DE$<�͗2-6�,�lQʅN8Y¦�;^`#�$)����s���3��I�	�O��.�h�Ҷ��/0���U\$�"h}~ 5�D�#���X_I� #�]B�{ٝq]�I�������4�aR�6Y�#\~�/�s��m�_�#(�s�CAV�iR@�\=6�=����
ߑ�?q��!8f�Ț�����%���IG��Z� �&�Y�����OZ肞I��kKS�y{�(����~!�����Wژ�/FKL0��&��^y}�+r_��ާ�Q��� '��<�����>�>�M�bat�n���r�w�n����U/��X��b�n4�(_���$Z�Qn��]%T�!��HE�-�s�2Ӛ�"D�_��i:��;�0�f ( ��M����U�p�[S�<G�Y_F�`�)��f\E1�7L[/�;�>'�H�DE�m�I"L�:%��������ԧ+}5R\�Q� tR����pN�ȓȘ����y� ������E/�h;��/�� �IKD�Ww@<S���!��F�;����ʩ�^RbXf;�
<�}��aW�*:e�h���E��w�ϛ��S���績}O9��E� ��8�d�FI6F߳���Zت�spl��Y^��/b.*���D�D:��Ĩl}�T�\-���aT|;ֽ>:*�]�eI��w6������q}�=L$L��W��%��ԛ�M+�	b!
��!��re���� |f��K�8�(ԕ�r��Dv_.N���y.$䖙���H����;��p|�|v/F�5ݫ�|���a*����a�E.��
k�]��
!�A��Mg���O	lh(Iߕ_C��o��-���WS�ɩ���)�q�]x�v�]*à"єN����Ot��|5�`��z�\��>٤]�]q�{�k.^�H44SH�Fm��4WJ4-���Tg4�f��Qj�[3�Mo�U��׷�X�a���L5�},�>�W��ţ0@�v���lSG�NcqΖn|����
�a�ɴd���s>Ϟa�*�5/��)��{|T��-J�"��.w1v�F�z}x;���$g��cE�Q��<¹;H��ɥ��a���*#�Փ�o���V��,re��G�`.�=�^�i�P]������u�d�(z���&����[��7l�1"3v$�ѕ�isΜ��8���Vp�mq��{���<L��U���R�+��ה��ɕH�/��o�D��ST�}�"3�_����[�Zi��5�^��2X�u�/�虡1#����	��"��u�n���8m��k(��|4��`���w2W�@�^^�*��f��Ù�Q�0��t�\��ao�n[�y=�ڦA!��z�˗�m�Ba����mjؼ�!��zM)�H`):ۆV�h�=+N}tJ��@��P�! �=Yj0'���#HLh��\:�_9��j���d���8nJ�%u#	\�Gq�)*GqD(�/ii�J�fb�ӭ(SH�C����8���s��Oj�t�H��V�*����z	֮��S�5����Y	�ON�'U��p�h��p�h��w�bo��ei)��E����G^�H^�� ���Q���6��@v>=M%�gA��`�!�e��O�.Q��.�Z6�ږ�\X��:,��l�4��-3.s�y�@Brw"����PG>���:n`7~>2���.ܶ,�3w�#�\��Ҽ����KIP�R��K��t�U��O��@���<kѪ��ѵ:�2=u]S���h��޽e�MECЭ���	U@ؑH۠~���m7�-�Ӊ
0�\���0��b�w�9�d�"uz�1�.&$��=f,2:�V�`�ݦBq����YwU��Sg��s��^��G��`[�8������gՐJ��2w�fb��Y#�� Q��%�Ï��fo��%��q��������G�m�~Wv��b�x�/j�a}|;y��Ԇ~YLr�v'{���	��c��xRG-���>�B���6��vB�P�%�W'.�' L������ٚ���'D�N��E.�n�O�OfU3��c����� ��E_3��&���s0m�1_����
�kK�ќ�)$쾿�e�f�ʸ��2˩#P@#�����f��39�|�ȱ\���O������G���;1��z~���~[��<	�;�L�4�$@���-��h��H������-z�Y44����p��W�(�u[�"�Zg֢�˩M}vd��%j_t��&q�?��{S�g�8~�]+�Q�i�o�Ua5�	�G(@J��8���z��M���O�k4�4O���V�j���h_�м�IɴaPIS1)ү�&��ߒ�7SL��и��<lE���Q� E�Vښ�]��3>�R<�nm��h�++�LZ+.w.k�+��>�|��t'N&ԖJ���2B�t��ry�/�&ɝck���1,Y�蟜S)��S�_�ZY{.=[� ����v�z�����&C&Snqa] /�kj���8 ��eR�f�\�
3-��q�)��MO�ek}s�9��o�
T���S�R��;�ҪQ�|xQ	���}̡�4[�;I�)0�q�ys��i���O���|EU�5;9���3]�0��W����`�?xpw微w��v�`yn�#�n�]1�I�(�.��M�~>�:'d8]m��{�ܔl�!� �F^2YuKkM�5XrL�e������e%��~�D����7��Q'��8��{�?��[�Y���2��G�.M]z�`��	V&��L7[�jK����35M�P[��$2�NU[��G	aZ5[GtP���6���c��Wi8Q߯�����Bmt�L���h��0���	34��p�l���2~J�F+��e�8��K~��q����]�r^�����a�����C��<�V���٭��*����wǱ~҅�Pc&M9��u�d�;��F8/iz��wt!�����o�2���NY*�f���Ş$s�KPGN�7��*(?)U}w�`Tt\O�b*aw�z=���T���[Ԡ˫���-���j���u��b7$�%1O6=n����_KE�s#V��J��3:ќ�^��WQ'z��~7���|��s��d�p3��
lYv�]�S.� `��z2��M�|:G|��x/n���р�BźX�_�n��|u6[ǒ1��}
�b{�Ѹ�9a�x��2��L|��1
�])�hQܹ ㎍��&G����d-V���w��:��F|��mbeV�dwӺ��a�:3�\�.L8*���·{�-{�C���[9�fOb�Y�/��Q`�GΜ�h�ܑ�P\�x���&��E!V�75-V|�>�>Ep���S�ȡF�"<EW��^���W�U,�M���(�[%:a|�O�Џf���J�p����.��X�/?�oj���@��[��,C��SF��@���(�.�pֹD�j��P�g�s[�mL��I�\Y��Ҭ
{�U�� �T���9��V�f���z��L(	�������D��E�����g+�"!���V�ύ����j������E��,F�����u�����|�φ9rд�q��F�+Y!q��N?�n�KO�t����b��j'��C�;J.	o�]
/]Ʀ&����K��U*�k�����~d%^�w�kO�K�f-��k��g�Iv�	�m��Ƙ{�x��,`����gǋ��ȕV9�u��s�i�t���X� |xW�j8x����4:�-��C�T���'�Vg��4T��#������f{�	�K	�؅¼k��{O�&.MI�
��J6��m�(i���� ��/au�r8����գ(��kE� Bߞ�2��b�qAJ����w�z7~�H'����XUS�T}�P���A�nnF��X�KG��b�Q�.��W���:o1�B;߃L�����/�"d}5��/ٮ�����x��**���0*����G�q���l�t�'D	��ox��Yw%�Ga#?�m�P���<��x��6k}��$�G��*�[�g��Nt0���^L��Vݓ�ZT^�\�x�?�ׯ�(�<�Će����&�⑲�(�9/�~]��F����s�O���%�,i�cYK�M�߁��`���0�$��	nm�h�F�+X�Cj�o;`�O����c�D��`k��./w�Ԃ/R���p���D�'��<ӿ��Ty�I�Sy{g���,3~�r�:f���ɨ�ƅ0�;@JSܦ{�mt��^4&4�J���#~�yX��m�k=���Hk��s�3o����㈑x��,{����"�ը
�<�Z�\6���Y͚�C9���l�r{>>1���|���j#vx �)�����+/}��x8�fMȋU��`K���'���z�I�۔rKv����>��s�7�W�~< �j1�4�#�����/�1�]ִe��;�q��=�h��rS�6��)�,LXS����=�x�KM�I^,I�F��� ����k�Ƈ]�����6ܥ���q���-����v��"-��}(�b���&��w\��"=lX�&��Ulכ0���9���J��<R'(��~�H48ݏI���UGp�|����{d�V���t0wO�c��f�u5���n6}᪽����=����,�D���l\����-�s
B�'9�~�Y��B:���ͼ� �)��}�b!	�����B�ܱcP���K@94���+q�~˭xٵrle�D������KDKr.{ǔ���^���r�_�m��E�}\C���i��i'��K	�׾?��8����π ��P���4����Ÿ���4!�</y�7�6	3�������k�_�ׅ�X���̠Š�QSF�y�o��J�E[=5ʆv�������X:���bծ�1R�g�5}�I��J��;����;�X���"� 1a��A�:oUX�J�؆~�7<�ppE
l� ��9���
������k���.iK�ݺy�k�raC�f*_L;�r��9���΂}�j��z���q���eF�,�o��HkN�)򵶞��n�r}����4z�"�O��+�F�nk0򵽏U��x�$���ɬ��q��̷�>�O]��*�����\ӹ@�Y�i#t��"|����Ɠ�}ʎ�\f̖3�~Rٵ�E�k��>�f/�S���]KC�er�pɚ�~����Gۦ�T��C�T���~e����a�a��e]�]���.!ӑ��u`&X��)����^�F����2�D-}w-�jP����Y�Ԫ:bo/3���?��0>��Sa���0)S'���8�ڼm���Ām_LM87�<.e�(����L#g��u�Z�1VS$�U"�c%eivsh���cm�@�f��`�
�[Йw!O"y������n�;9�aq ���Q�{�V�8I�/	���A?���#'|~+�.Z���?�(O�FB�aӬ��Ⱥ���?�����<t$�a�����e�3�ǎ������������G�`����خ@�9�i+!+��[T>���&F�f�8�g���q��԰�e�5~��B��z٠r�Aσ,����b���hW��\\��j��z�5N�؁���|A:��D�?7�����a@2��S ���&f���q�E'rv/R	O��"�R��ݔ��yi�{�^s{t�+kh�#T���/�����_,�Y�6l�D�l��o���I�(ٰg�|�ǲ^;+{P�[��3�_���R9~>���G6��x�p`�҇�o��򫞞��[7��Ղ�'�[b�����O�>*h���O�� �%�B4]� �Kqm`�G�t���{��S���U�{�)�i��E��Tp��o��wC_���M1��Cxf� �+��D��[ �eؗ����q�~������T�8�Mb��� �Nh���
�'��>�"�ۏg%����0��F���~@�WOF��s�b�B��%�L2]dRI�t����n(�����i�}Cm=Ax��G��/P_A��Gj�FCC������t�V��OX���A01��� �v�N*/�!��	L$`P�7����<�X�^a�ώqφ�ا�v��t��s��z�u�F��ʤӰܣ���ڠ5Q�������WIq �<�<L��wݎO^�[�}p]l�2J�3#P1000���3*v]D4F�,�gzBi-�|]�$��D��~�9b��w�:J�(&HY���8��(\s[!�n��z���������Ұ��G({�^k��Ht�>NO�;z���%�u���~��3�<��Y�x��M,g��|���GfӶB�;W��<�v�Z�;��D�����7h��k��ls5��8��cA�]u�;A�H�Tp��:��������Xx�Z��SסU�6j`�j�#�^A���xw����V�����3���a�-��WǟBP4m�
���+d�����b�@<���WA��h���K)���x����5��Iq_g�Y�`[(W�s?��`�u9xr�Z��8P�]����� ��l�FE�H�M��I���ې��}k*\�JĜ,�;r�Cp$k�Ȍ6/u�s�����8�F�9)�Aàb�Y6�NFV	֪$�����k��g�A>���6�nq6_(��^̦�y_ғ}��w�s���H�t�C���A����y�%�(l�=/�<�y����Fo*Q�:;����k�9-A��a��KC�&�>��hVۙ\��+D��ul,Q�͛}����aS�j?������?gJ3b:�/1c��頭��sp�&?�s�5�"�A���ak��� �i�0K�og�2�+?����	 �^�=���xz��k`��v�F^<]�?|e�ԢN`e �\���T9�R�
D);9 ��u��D�(w�?2\���--���6�2���@���c���o=�޼�cY�"es��^v�-�g��SW&����r킋�x~�N��>;��oG����%�(�1>�V3!l�)��k�s9�1X�(�R�*�AA}���h��[p�7U��d��~��Y��#���-�ʌ���{T�T3�t���.#s!�{�5N�	��gSgp�A��X�9��掌&��c!Ȝi%�"f�A�K��QVl�b7!T����͞���T�ē�/��C������4��k�O-��>0�J@x3i��wh�`���h�0�%�[��i8����\�I���9?<A5�p��n�e��dDJ���F-���B�D�'?5w�U\�40���q[�
ɜ\�:�#��#�X����m��������t��+���S�������*<��@�@X5�����s^�9�3V9�G���/2���A����zɧ@�p[�{%<37&��j��`��N|����w���&�O��i�Pv�	��q�Xr_
�m�
s2ZJ�F�J2|��@ߡ�\�|X3�߉]�Õ�$��JE�EA��SΩX�`�Y����u�k����a��b�����O;��u��ʵ�փ��v>B8� ��5b����]�Ö�����^z'���sh2-���fTID��D��Y��Yn�$�}�Y{��q��x�H���XN�ޤ8fTl�<}JCH�D�r�棛(�ȕ�$�s�O+��svfJU݆���!����~(�|"�Mh��4���[����(o�A�5걔 `7�ՎV﫹����킫�	�ZK���&�z�}<��?r惞�Ӄj+6�fՅ��'K�q��/0��o���rp���M��fF�H����� �Ɔ���U5�8䜅�@x�;a�Y�~��BJd�^�/�]g]Gѷg�9��v���}cN�����O�N"h�O��R��
S�6w� �e\,;i)��������IEy���Q��<-��p���v^t��,>�&�ٰ~�����<1��b���i�t��,P�AH�5�CI �o�ƴ�'���ӱ�EN��EL@�1q{Z��Z%��s�VM�n�^�^�CB�O�C'�2��Z]�,80"_>���GC�(ٌ�5'�� �~�J��"摡��f�������?�;��kčٵ���9YF޾�)�q�?v�uŨ�]Q܎��E����4�TW` L~��R���H�	��G�Fƞo1K�e�}���g!;�BK��-�l�� �?y�bs"�/�8�cv3�B.������5���;��>����;^�Ϗ��Y�)�;;��-�.���}��j��^�x>��FP�r\��ؤ�B��
��"�!���W��*\�t�\�Z��.����b!����L������zrs����Ŋ�%��/�8?RzZy�d{ Kc`������r������V����:�<_s:��
h`�N���!�F��>���3�FJ�r	^�[�h2W�	�t+���<,*V* *r��K-R`�Q�	M"��Ge㏔��y3�&�.0qA�Ɇ�fB΄*`�Ǡ�E�vj8옄p�Q��\B����$�j|6Vcz�ʥ�裡��9�w5~`���8��)(M��Z�?��=Z�,�q=��3�U]���5/�3�{�'��ۢ"}�+��nބ�)�|���Α�[�)�{���)�[f�������T��`hk�˪J��PO}d��a��4��\���ڔ�%��]�5\aX�E&<ƙ�q�H2k���2�3)>�-^�[��U��q45��*@��x'������k�=����@PXla��d�>��] xQ����4��͛z�9wB0;� �?���"J0UG]�n޽|�k��K���	ޭ�2�=�=a �.L����}<����J[-��J��gz}��L� �
��מ�[�����Û��f��� �q��l�-H2���"%����&��#Ѽ9_O�o�j�i��K��� u.'A�o���˩ 
JTE๏Ѹ_��B�����@��:���LJ��gCg%�
❹C��
<M> �i��+�i�@e��rW/��r�נ����	.	7���?�pR�|�-ŎKQX&�R+)��>�]�����Ȣ�\%�������r^1�o��e������X�m�r|G�5ԩ3��*�f�K���l�Dח9
j�!U���=*�d���ΚB�x)Vۘ�ʘ»�I^2�I �a�h �UMle��d��w[�n��#�?�P�`�D2������ظ����'W��a��B8_�����2�3�!�+2�z���	Wn�S��טڜS�g��^��_��hvT1�����R�U-��T�f/�jK���dty!P�P	O�,Ʒ��4�F*���}]'�k�[�X��֕�`k��2K�]�+��w��#~������MZ")���������.�rWkK�ϊ�RO�!1/�����1��2���`���"�_iT\�^9!Q�X����a�����!h�# ��d��a�{�vq6�xIm���/|�dX$�y��
����C*#+� ��R����fe�䋂�L¬��o#��4+
3%-pMï w얢��ov�Ht*�$��:$���U��
��Tu�_խ[&\���a�;���a<��=T= i���.:�R��i/�n셩�/?PxQ��P� ���j6,[v^�Ԛ]��R��Rqr�"[��Qf�'>q� >2h��p>T���,�\T�eC9��lC༠� ��T+���#��!9��� �DJ��	��/�T�>dj������쨞�ow�������8�u��a�|c�s+f�Y��{�n��A]k�i��;%@D��	e��O&��d����P�g��3�&�2<���/����"����Gݭ�?�=^��Q�9R ���9U���x!KB�_��9�z�>�R��Ɂ�`Cţ��W��4����-��L1G����>O�7�������A͍,�
���krdCΕ�U�B����?�+����У�SY�AY�r���q-�2JC�滘iu���^�o'i�?F,N�M�e�cG�tF�}��]n���^�"U�*���(��ս��MJ�i������:�^3��dW��@	���=���#�(3����9{�fhsS[��wq��#ru��7�vH������������({H�z���>#�5y<C�U�U�W�aA0��a����;IO�R\����Q)��g3,���Aw=�����#Ԫ�C�M�/����t�t��3%D�ß�'A���z{T�U��@�eҞ���W�ӰOm�G�%P=�37�hr�A=n��+!K����F�r�S,A�F�ZUn�7��Z�>�A)n��D�ĝO�zd ;#3�H2}�]���Ǭ�(O�Oo��vC��Ykʺ>��e4������6��3�7�����ӭ�kTSOk��K'��U�:��j���0�[��7�q���xtu���4��<7hd
�)�����-s�b��[2H�A��$^���Gl���z��z��y��R�b��uCZ��.����U����E(���if���ş�'e��N���^�������(���&ל��Tt�M�� }�jlBgsP��N�� jׅ])°����@��0 L���c�A��F��vz�����t�Ŏ�wQ�����L#������,��l�}��E�F����T��I���r�"�������J ?K:� 
^�$s
���[�����������LcĢ��ᄙ��u��Α�h�8�g�A�a�Bhk���1�����$�!�ب�f�	&ω\�b�Up�� Ֆh'uؐ�4�u1o�m9���~/	�(�=�h��*%�-�hr�o܈�x�.�D$�;|�&bm�)�`�	^�E�+��o	��߄�`��
5����ƶbo�y7S<�Ǥ(f{�o�߻�2N/'�i�^��>��M#��/���	2�D�_�����Sx-��f^=B��G]�]m��P��aE�
��]��׀)�"�&�*�SY�b�B��xRD��������lC��ݾq��s��(���x��t4{��WU��С��u~��N���������h}���xl�&D�x�(Ӂ�#̃l,o"t��� ��Ux��;�[V������%�.�N��x�#eŹ�䞒k!��;<�O)�@؞B໘/Oz�� �"���tz��������6�:�c1F�cV�!蝦u��]�C^cα�~*3��.����I�~ѣ�eUJe��L�븇V"��z�*��:?��&Q�����Hze�T�����I|��k� ��_� �u)u�X�1���U�`�t(�:�d[����B�>�FqL�q`���w��v�ZW6h��Zݷb:O�@Zw�^)J�±�"5N��v��b
�>AYru��Iq�ϰ7��
���ϣ��E/1����)�[{�R�rC}Om
a��m0祘R��ϻ����`�S���� �։]X�'Bd�D汙S�i���j��랕�d���y���\�b�.#KW�	 <ꣁ�ϱ�z�T(I��^{s9Ϳ5]�떝#U��&R��Z3y���s`��)#����q�cg��3� ,b�y��m�rdk,R��6:�'��拘�gE.�^q�Er���R�f�}Ҕ:�;D0�ڹ�t�yL>.Ѿ�>b4� ��"����F�U4�I#�dhjNQ~�C�j�Hc�g�n5]S��� ��ٺ����'9s�戚�XÐ�.g���� j��V;�i���ڍ�OQ�'��'�f��P��ס̞�/M�V����-n�!�CS�b��bU��㑣�m��z�F����<���꿜�?kf��h(u����#��ߎc�AJ�r�	ܥ3ڻP��dnl[�8�+0t�F�3R�qQ^dKK<m��)��"��I�X�Le,Y sy�c�BY�]�~A���uJ,�r?[3vA�z\cy=�ؓ�;��ŧ�@4p�����U����:2�dFڹ�.�1׎�4���~��ʾ��3]a!=�v��U􎈠o��
�v�b	���p�9?[�N&.ڄ����ý��d3�v�BMjBA��ɂ��.�p�4�2�O��	>n�uu��q�m�C��(|3�=)��C��4%�����J������ ����!:�&�F'�>;s���ٷ���a;
?�x�����5�d�[����ٟFo8dc�� 6�m�V��r�@	Y/�'m��d�7�^���q
�IiQ�>3��x]V&���XV�����-ͽh(`C�b�R���S�\�T�x� 9Q��d�c3*|t[CYP���)��y��u���j����D�$Di$�u��i�㏈(s䚹�ij0����{nZ�Oe쐆�磗6����{���<?2V�ALM��t��K��zK}����~�2�^K=ӵ�Q�^f��0Z�ޡ�\wc�c�_ �+_���"���Lu���`�1E�c��Kr�
�DQ"�w��政&l(�����G7Dl��(�~��^F��u�p�ɖ���T�HC/�Ilޖ��f�Ja�Ȃ����m�'ۜfQ":�`��0ޝDvr.c���HC3�(3 ��_1(�΋j����L�Ѓ�\g�O�Zt5�!c�&5��%<[������: )e���Ɍ�H�}7��@j
{&�@}q,�6%�|٫!V�Kt�m�@g�@��O�9�!F.%�@"�=�ͥb
^��'���2k� ̀4f�����cl}�ׂ[wi5����j�>��ܢv�"���?� ��G�ezE^�Ajk:Em5
>�.��3�1���Z����}��ߛK*�6�ƻ�*��
�"s�6�Bt������� a������Y%FӶ�����S�����j��0�F}��c�9g�$W����� N�ex��>X!��e����DTߌ�oR$�[��z�c.ɫAj@�dq�	C�y�N!Ȗ� ��i [�pj�,�e��_�_�Df�Bz>� g�13x�D�Y:krV#���͋ᨢ���Jd���&���\�XR�sM4+�/�b���T|��?���֛p&������3R&u�r�W~�@7� ,��U8A���Rn�)���3`�6�� HgXs+n<�T���bu�6eK�Bk,�9UC���*��q}��<���b�&��O;q�����~���׿G�c�Xm��M*p���ƙi����^��|X�܂y�ͦN9�5�rK���Ȃ�7`,��seJ��� !��'�/҉\�{�ʖ�^S/�#d��6(�|���;�"]�H�֑��0%��"S�C�8�� �Q��e�Y�&�f��>�[����2s^`W-[c�[��p���O�?̪�
Y���������j�Rc5N�7[4�y�TE�H�0j�%������_�CrQ��1�~kϞ���d<���p��ӣE���ɡ̴�(� �_�:�� ;�>�{�oDd�Q�ޢ�oI���88��#P�@�r�?�D�pοo��4ʎvޖi�M.��Nע�[g*5K�Ol��w�:u�mAR; +'��mJ���K+`N���	�(�D�D�X0i��9@�t[��i��??nz�NH��'�pA� I�X�������[���'r=ܳ��_e9�_"or&�<婁_|Km�Jw��`�V�y�3�r�-
���yG�L~�.>AӞ�%?��wS��i�8��躤���f�;��b��:GC��&�.��#�O��E bb1a>�#fD�0<���T3�~�dR+R����� ���xn�?�K�/b�j��d67��8u�������=����p�կ�Lϓ{��"ާo�8\I�������x� �d�-l#�h x6��<��:����aa�;`�
zKz@��l�<I�{�N�	�_��|�9�Z�ek��{�A�~��i=�?�͚���Կ��+��3v�\j.�c�ݹ
`�V�_P.��1�f��0��d�r��~K�p��59��w���N�	@N�{Kr�$wO�Ix]Y��>m��}3ǨU��!έ��$|�ܛ�#��]+lYc+���&k���G�<4��?�8��3�I��R$l�k��.�L�[���0��cw���e�&�{�:��R�M*���R��E��4b�mF�c����9 ��ޏ��S���EJ
���P7�_/�ޔ-:@����SđՄ��{�g!r�-aMA�a/k�.5�#�H��]Jc�������4mB�	O����,;#��)��8�鯌Me��L5�~׍ʱq��ng\�YJ8��<|��{�g�r4�F���}$IT[���p-���tE�UX�sq�Z�N�w��W'O/�m��c��L.'�5n	GnYU2��j����83��u�'�?��m�!SNfi0��f8�ro��$1���)8Wb���c����^��M�)C2���\�	j��������0�.�
0C����xDu�w�X�Q��I�T�:�w�A�^��5/NN����y�H[�Ӛ[���3�N]H����]�^�����Z��Ϣ"����m|ѝ[ܧ[��9�P�%��T���g�_�����m�6gF5������D�����	��"~��s)N`0�C9�xy�~;ツ���߉֦�$�u;
���[G�|��%�@�0?�{��zgS C�v3��x���b���[�ɴG�Dȓ�7��|�aY˸���iG.`��Û�z ��\�.|�,h�����)������^�H�&� c��i��EKһ����"����c�d,��0���':�5��2�����E��Q����vDx���' )cOX�-������MΥdA��0�+�D0����ŭ��m��i��W��?>$F�-�6�hʒC^x�!�D�m��9�
j�W�s� ��w��ۘ��^��}�U#��8;/�{��+4�B�t^�w��9��Ư�x�9�\_Q�-=��Ƴs�ǺE��1� ?�.�S����FK��o#���أh=�#�Gr�UM��/�
��:j$�
�+Ɯ}�Ni��M�JXv���s|�fY\<*{�UH���|�z����cq!38Q��3E�v����������.3?�1�/�6IR�X��m�99�BfR����d/�0�L�[x't�S��sl�o�ȫ�cO�Os�oN^�8��HL*A207��mo�ّ
����Z5h{��{0T�З��\��+���Y
��.�E�g��Y�3�e���A��K��d41/�s��"p����9��s����*�� ��"�rI�A��+���y��7
�e���!�Mnx�gf��7H!-�� �(k�@�?5߂��-�A�2�_��?�ww	;��\�G����n�U�[���A �������j���4�{�_�%y��`���e��۵��9#�N)^��fl_{B�٣M,�뫴��8)@g�7�;5���Y�>��/
�gWl>iLN),�5l�ξyB����ɟ�a�Ͱ׭��E���L�0L�q��3��YMؕ��' &T�[ݤ�nM/Ba=j�]4"C�4ƙ	�SǇ����NE\z��9�6�x�M�P;:�i�"�5�\ ���;�އ�~M��4u&�e8g�������l�A۵^���&��ݰ������WU�'��`j��Y9�'j��C#!�,��I93�mKv-�5	b��oA��t̥�.��Uf9���#bB3x/���n�H�GL�3�PKҀ��Ab��C=�A��{Y�R���c��oT*j�uq<+��<^��:��?��K]𝛨�A�C���841�K����PB�:z���?'1�h���8UA:�{�l���o��[V��t�P��H�'�a[$%���C�=�g'����B�G@1�㼗<|��lgJV��`}��,$\�^rar&��gt_"��x��ϧA�{�y�&y��b�1�~�|q�cfߟ�6���K�c�oW�m�TKg�d����r�;@[�	�w��/@��f���}c�58{w�!7?> �\)-��Ĩ(�����\^���oA�P�����8��m1�t��>u��
�L�Y�ɮW��~k"��'l^�2��'��ˣ�8��Z �Jx�RX���'n��m�zu�\@�ԛ�ǘ{a<�#���]��:��9Nf=����H����J���;'c����/�c�S{�I*p}���X/����mHG��u\�����l�K�������\�M�h�H����/vߣKX%TZ�S��>b��D�&%���Kn�C��a��i-��d
�x�"����،���{PЧ�I1#,��	�������u�- �^���@U�@��gK:��U,���r�ÂN�:�C�?�43��\R_2���ǻ��5��@C�6o��7^l/>���vu�)+.�gN
��S���wy���=f'������?�Ș�K�۩n�"�d��XT�<��gf&�3F~�TҲ}�=m�=o�oXi/qT�i)�)\hl���M��vwʸkoI��5�t�@xߺ:���>t�c�"��t��A���/m�S)�̸o^��/�5��W&��ü+�m+pG�
�`^���&�]�,�|�/)EW��@�:��ȯ���i�xV�q�/�Jp�C�*�
���n�X`���<���n�~5���:K�����4�SZCx�I�r<:��51w�.�2�8` � ����q͜{�r�d��A?t+�������Z���.w�K��9�\�V�FS�i.�pe-�9݅K��9�
�J��l��}�&N�m�{��{L@����뤗X�AL��e����HCk I�h�+0�{m�_���44�aR�6��'������������ϧP��cg�$�j��6�=�ȧS�t�>l��<�W,_,���Y	��.��dIz�^�<gχ0A��_:�"8�.�(�e����۟��<�^�]�1z̙���o�����
�1��[X���V'`�gS��u�
�H����ŋ�f8��&���⮕�+I+[�Bk *�#5X-V���j�>�	���/(O!��tp�.B�n�s������ֆ9�p����:W�9m�SL��i2U�e�5���`L��3ZRbeΑ#�,5�5����$F���3�� �PvW�b��
��'s9o�� ���k౺MA�6F�qC�\�e�5�(Z>Ұx�X�U��.㘯F�I9�ۮ�8)e6�$�/;"+G�!����c�dl��梳)�{��wT҅|X:�}.�1[O$o���/Xx�tR)yI�� ���+�^ ���/�8���c���\��K`���0D��9=)A��ݒi`V�bigu/��R:ґ�sG;5�X���GyH~���U)��2�k���W��)�$xl�� �;O��0�zqE>c:ƻO�΁�,���V�����\�1'�|�u�`�s��ͅ����ׯ�x6=$:B�f�R�9���o`�җ�@Ǻ���x��yo��Ҫ���m�^%j+�M:�5sZ|A�"Y�c�pg���HZ��u,�e�j�pFDϢ�mPx�f�H�����	�UJe�m-ڴ��Ax��FoT��ñ^�"�Tρ`臊-�XOc)�K��gz����3#�j���u�w�ո�ma�Y#�T)��ܶ������h��&�K�����SE^I�����@�O�ə��w�E�����
����rP�ÿ��<-߼��𧒯%T@]!���w�`UL��6��d�u���Uf�zM* �>3'"������OG^r'�_�bT��
:��WʡZ��i�q�O��g�N�|�؜S6]eZM�T`72{3�I�*Zu�7lzd��b��k��]�@�8�ي��'�8qѴ�V�V+p]�ZѮ#�p+����R-���zh��O�B|J���rM�3Щr=�*6椾4���ſrz�.a+���*�LG��1�ig�����o1)ˎ�9�����~�N�+' ���x*i��M=e��;� 7�*����|��g��X��}�3K�*W�얯��;�[�z%=��S�Y�/)e�8�0�`��eU��$���O�Ɓ� ����N,��-.<�{\�(-Z�(��M���:�� {_�!�7��$נ,�b��pVl!烪 l�T��%j���*s��L���C�E��*}�v�ZD0��@6�P���D��&bJ�\���K�Zz�򥴏��^��-�\�,^�!�H��/^�u?~�`L�S�.;�����m�E��'�|�#k��I�v ��M��V���)GSs��`ԃI��4 ه���0(4�i��4��Lzu�s�c�l`�2s��O|�V�g��G�F��'����z
�H���(/�s׿͓��޻V��-����Ѽ������-~(I2- �8�$5�H'We�ׇ�.��̉(�q:�Cy��j�@,�"a���T���W�w��A��m�P
��WG�FkFf�4* �A�i����T��.՘����-�E0V��T��D]IjI�{�x��r7<�M�#��i$���U�d����Tщ�$��uE{����R�/�Ǔsmk�*c�ZOω|�I5�~a�^������zZ�Y��!� T�ӝ)�TC��t9X�%���H�&a�[����:��~N|�l;)a8Ʊ��&8L���73�9�7زU�P���m)ǹu���_EU�p�ǋMNs=G�"0T�8�/�]�J� +	��Q�V�/�Z��6冟G�Y�
2}���3m����'f�n,�ߙͨ��
�h�oO�v�Óq�j�D�!w<�&�Z�c�+V��.�db������P���X[7����Efs�!�赯�ٟGX�%����f����v����\u�͓�3�(�V�J�9,z��D���#Tg�~pەO8��0�S���KhIv�<��,D7E)7�/����/S���<ӓ���mSJ�.D��o	�U����4np0�+X�M�3�
3��R�䎗_�DJ��t4�w|��6�5����Nx7G��������yw��X��H�O�5i�]�9����}n�aw�R~�~H���J�zY���G"?
KQ
�K��X��w�_[N�G�<,o�Z�l���o5D�6rC۞Y�@e�0���D�HP�)���DD�/h�����G(���\���2±�r�Z|f����Гj����J9Q�j�<+����u9��f��]`�(�z� 
���9��Ɍ���0/v��ަ(Ȍ���8F��E�9%�ӗOW^���R���_��0fdX!��������T��2�Fb�z�;*�9�X�4�\���.ÉpD�B�P{�c�W�4O��S��sV��S�����������X�p[�vK����J���Y��3^�:4�-F�!�K����ѱ㎄Vx���!D��a�������]�����ɞs�0�o�M�hc���+osG�����i��v�M���r��cu�?��Ѭv�
���W����>R]ZE|��rfNl���1��7<��Q0kn��"��^�2��q����PB��ŝց�YNm��r�v:u��٤��і���Y��\˼V�r��[����Z�yS=�R�0��/UU�?��_X�����#�r�U��)�Ztu!�z߾�XҖetd����[>�V�bR���k/���0B��A�r ��$����(fᬳ+z���l���Makm�ڼΊ�y��F�qթ՟��:��Q�?QA����(Մ�,���go*RQ����u��3)W!��Vl���i���e���3�k��ub��^��įgJ�Ϙ�J�c�
��w����z�b��o���'�Ц�j�ˌ�eĚ���MKw�|z%"]�ʉ�
.�S�����9�`���8��[�p��@���1���{g!����4t=6�.���3!��(*C�����}�k`%�b�/��P�k������A����،~�Sǽ����ߞ>����@�Q ��3&�i*U�s��/PS�E�A0��W��kiU��L+F��Ȱz���9�s��z�/�P�M�_E5���_g�U��t�5��(r��x��l�^��� m�gƾJ���+�H~�D{#�R��ѱ �ؕk�3m~P�̙q'�c\�=M~>����^�gӧ��Y��LǗ�a����fw^�vO2�P��W��;�Gދ�4�w�X	p��8���a��'%��Q�	*ݧ�R����Z�fd�X'��}9�v��3$k7J��5.�T��\���h�׿m�3[�����x]޷#��
�v�6P����@�(�C"5uX�8}��x؍��~�WO89�h��Փ�Ɠ���O`���$��)��[R�g����HD^Hd���CN�E���;��,���W�n�XV���ڃ0y�����9oN5Փh�_  U�w`n����M�1�g�M�)R�<�/�q���$���|��V	e����m�v�]`1������՜�8$����Z�:���G�|�Y:����Bct�{��4�$��0~�
:�����b�0_�<�ݘZ���`��NL@�gY��{�3���>ޑ߿�=����1�]��J��fY�h�h�t�?$�򅡘�{~Bx��A��%�)i�\��	�M)v���?]�)מ���2�v����Q#K����,���������a����k�sF�	���R&I<�#"�e]�G���xPvVE����7���c#����罴��Rx��,v�O��j0����uء��
0>�GĲ��mm�5N4o�R2{���ktl$]q^|���jz�.�L��t�
�@����;"�"}��i�F�0b�7kS�߳��E�����L�����3����P�Ũ2��!��js���8��e�<$��w�Q�oؾ��#/���.F�_�T�e����c�_�.�x9�*��������W��Y�������L#��-��G�{6�'%��bN(B�3��V�ᙧ8�gH͌$��.$:7�"J����i�	g1��!��{�/ا3��GXM�WT
V�W�#�r��"3���|7��)��Wr���Z~��7�v<�&ZOS����󢩺�ˏ���w���i��cI�v���,�1�t��=X��'��'�ɰ�1�٣U0�y����Ofk�2�`2N��},�p��E�H�Jx��Ke�D�o���@�&�cf�/hޱ݉����uϊ쥸��n��3�d�=�haT���(Z%��4���8�u$��J��J�ٜ�����U�XO�z�|��%[�&Lt�_t����� aq��Y+���栰"V�%ˋ:��+�q#�7`u�ܻ$e�<�J��v\X1	�9�	qo���.�k���N��`�U��c��M��<W�#�CZ�W��S�!ʈ7B:چt@������t�I}=���3���C�M���ɠ����g�lGH�~H'�h�%���,A_Bo���L���3d��Rþ�A"fM̲�%滫	��{^�D8VI���ɋ����B�+��(<f9i��	KK5�65Q��!�O���)YKdى �gQ��B�I�*LF�y+k����X.=/��w�}�eɜ�+������=��!��G��?�6��6���©"�Af�8�djTM�x�d_�[8���UO���YNT�Z��3F����Ȗ�@���j
�CXΖ�)��+�@�-N<ЅvڍJ:��24����I����{)�X�wna������>h�_6b��Mtot���մ�S��O�d|Et�r��qE������`�ʓz�Ǒ"]�@(��쉌ca��f��YWq{%������Q:ڑ�W�����8j!3��#�ϟ���#C��h�PN@^�`�.zu�FU�?�mR4�5[ҽf��7OS��G8r6�S7z$�({��������:�f��U���]��Qz�V���*Y��d`���TDa�
S!�}�jI�"�@���WS���1�'���!^�ˈVV��&�O�/KNV3[}ɉ�?w���x|�n��Dӯg�z<5�A���������`����h�t,�%�/�5�L9�����c�<��{�`�.�f�Yl{Q�/Q�����
��;�+c�'5��'�Ȣ����3��3����'t>����C���!��� mnC��s���"��x�X�UtRS�u夝6����mu�^��f�W��>��pfM��GHsp��g�ݨ���x��[4\+�YD��g0���f��P�E�nM��33��=r�r�{ֿ�R��l݈%�l���j�ӥu}�?��5X�I�#P�Qն�5�P@I��)�<�.Y���SZxhrR�c>+�U�$�y�B���I�����7��LR��_����]�L`�C� >]�f��Ӎ�Ԥkܰ��T��w�Um>!�N���0���^�؞n0�DWΪ���[���@��"���t0����D�6�2dId-:�=`ոc+	_y2 fyrI�E��:Jd����p-'b�v�RԜ�jTO�!Y�����Ȫ����Ն�-=�'D]-�����9gp;�dW'��_��\3>s�?Ҙ
��Qg+�J�[����E��\�c<��g�*�B��n�c�汢˸��dD4#�л {����ݰ�{�����/R��ӯ�WP���E,�tL/���u��r�3��Cq�PVWu�>y��V_򦜡����qw�1�NAO�#�I�{�i4n�>��Bf�O�׿�R6!���~Z�=��,:v��3��_�(~�A.��$�QC��k}}ӈ��ֺ�C��]�p�bq���M#jz���}��}�;mҒ���є}"1�!��r���x��޵�t�̀��v���UqjF�����?,:Н�@tH�2��� �m��`��ET37bL$�Qe`�j�^�[@����ݶ�Π�T���VFshk�dF�x�͍٥{��O��HbObB��(_���jlLq�*W��p����)K���0����=I�n�e��b�]r��f!��\^���I���p�A��nȃ���?	'}c#$\��`���j����p����o�T�[�O���*���!�`�d���	��i��{�d�6��o���	�cz�x��}�[� V�&N��QERw��*�F�_�K�m�A 83��`V�k�h⎪�v*�jLG����ۛ��b�a��ˤ���:?ϡG��#��X>���IU��"-�mTtv�?�R���ldƱ��:���ⶒ��1�?�CA�^ѽFYL�Z�ye��&���L7���)�v����</�YxMk�o��3����|dv�8�F�&�
�&��%���9���D�����@0�� ��ʅ��#c��S���J��g�u7~���a����pM����g����'���.�'�����A��H[j��G�Cbء�tխ4�Xs�-b�0� ��I3�䛢;�M稬^��K�1���|`�#I���UԠ  �B� ������k�],�vS55���ȑzQV��;�*,z���5}9G���η]�[��Ř�Lo�p�&�ō��Y���=LG@��;��+�n:R��&Q����I��I��t,�8$��}-Q �í�d���T�YWЅΉ�@E,6�f�J}d�(Rj@�����݅O�E�\y4T�KbO{;º����H�}{Tuۇ��ܾ��x��t4/�ec���Dޥp�@oz����x��$մ�3�g����%�WeVp'~E��q�"�E��\��KH˥p�L#TND6�1O�~>�0oy���ƶHni�����z����3 ��<h"�
a{	��íj��.vo����p1��䴔{��J�������M`}rǺ��_��g�� ��a&S*��d�(ĕ�Ur����-Z4q/0c4C�����X��E�tO~���lLv_ڛ�v�w�����#$�����=����i�����-K�h[� \��lkøn� �gl)i->6�TVg՜�c��T�z�ѱ���n0K5�6�1��	j#&LƇ�H�)���Op!$s�4��-�1.s����h^�8*���vm��LŃ�Ps�����:���9o��L=��"fѴ<�����
�9��V)�D�=���1rGqI-MY���;��;i҇F�-�/��xB�x�¦a��D'�l���3z@C��W���H�2�����;��Sbk2UH8r��}�Y�J�3~O�0���G�n{A�\f%��r+�_�Q�K�.��]��K�⛑g��
�u6�.���G6g@ �h4,����{���ot��"��i���1��1H���� �Br���-�y@,~7��wP��l�\�n�	�_h���hPڊ�J�����<IF�׬���D��X	_P�5�-�p�yi� �$���\�#��GtC�_�Q��Wsh읗�:	G���-��9�Kp���A\�j#�W���s+�^GS�_e[Ici�N��;���W��0i����I&�-�0�#���ڣr�lY*8H�˥��������ĉ��'��&�S��܂�\ie���!���KaDd�"�]�4���wB��!MW�\�_��1@�K"%g�%����©�/�|%Z>�=5�Z�g}�O�؇nY�LS~�8_���y�>B*qec�ح��o-{�K#\q����yWh�W#�2�ɜ���T呅߬i.����b�u�����(�P�	8��e=�5Ҽ0(�Z:)�����ft�1�t��GuJ"An�/6x	�^��jyOf���9��1 ��n�_���s��.p�]�Z������i���B��U�7!�I�}�����,�B��A���{�	�MKOi�7��L
[����0��U�S�~,����~v)�fH[Oi	�B%�8@Ǎ�Ѱ 3����f�a�E��d���`��Ln1n�M��lk�4�J���%E��j�߶(����*�cm� Z�r�o���5�œ93���#^��hD}W䀛])!���hK=�@�1JUN���0`q�T;�BG?�9����y5�;�ڝZĠ�vP��	v�&�(��^��͹�#���6�R3�a*���J�>�м�q�7�Rı�u���n5�|�r��Qz�����0�rZ1�M����*����j�MaGG�0ޓ53�}��������4���́/ ��?�ĝ;�#���T������$6�Y8	��Cri`����H�����Q�S����~�Z<��wy����BN'�1\�r���-|2 0��v��/�j� ��K�f ����Qv��B�	g �'[���ѕ���&�:��:E�DW2�T*�\
\� /�z�}\ �a\�k���>�:�d��k&��U�=���k�)J��㠉<&/�;ŀ�2'�>t�R��f �nr��:��U+��I��s�U8iH��6��2��a*q�J�~(�ٓ���KXNgx�d��d��)p;�#�)���*��իd����KQ���������5�ᵦX[�5�~!����0m��~�c��yW��Z-��� ^h㿞nݤӉ�G�C�ː�۸nXd.���2�i͇z�9�o,-͔�.(B�2�o]Y�ם&����^��ܭ���|������2�T�=_�����z'�e�+3�)^<�<y/U�l�sUv�_����u�̡�A	�{�՞�w��n�W�ZMV$������ڦ��2{�/�4�m����$�~��b_�G\��
�)�"ԑ�>Յ��ȡ��n���>倚�� ������+2�O�Χ;��|�b�ej�݂qM����=���T{�ag<݌��4�C8�*kޙy'��2r��&M9y%T��燍EX�S������)s~�y7�/_֟n�|pi�a��k�?�Om�ݔ5fy������K>P���g+��(���[�r��qx�e];S�	DK�4;+��[_&�"7��������b�Yl�4��v��;ɪ�ҁ��{pѧvK5�TI	� ��18|w����Hh�{Y��47���T�\��!E�qdl�������?/1f�	�`��	���u��ۜ��')%� E�����Zj����!���:�R�(I�Fc�g+(%����m�_�=׵;2�n"/��e"�JU<� W�|��S:�X!(�B�i�n��~%HJ���������K�ݕUۦ�����a�����QM��}滖k���%��6*���
g�ݥ�b`gq�<"[�g�W8U(q�,�̡�*�1>O[ ���-��������o�3އN�S9���N�}�����|��L�����2��/�(#����aI)��d�IT��o!r����>0�ZT-�O�H/�"6���eW���SO|�⫉)��}�b��i/�vv2�?y5*���
y���L$~r%�$�[�����:��G>̘�����K�A�<kgU9'v%
�5�l���F;�PX} ҿLag��cB��J���J��S��t���ذ��R��*��R���w�mv�w ���hl��oǤyx��H_��r�=kVG���0�����eŖ�����#W�C�Q�T��ߵ��Hg� �I��}����@ҿ�p,i�d��}��|�_e�
:<�`��>�P�(M$�n�|zOp����m��J�ME|ͩņ���G�@�O�8�d�v`EY�K<�����f�P����EN���6�o��e���c�>�W�9* �$3���]z֮+38�nsK �!���LW�l�Iځݧۛ8aK��S��i�I�����͔�V��-�W��%�0���n����ӟ�K���o1,����~���'�(����q%��������Hi��#��(�Yhj���Co�������Y��R����ַk�w��B�^_YrT>�6��2�A�F;���(�g�@��v����+R�%Bh)J)a��IƋD76N�#S��n�k�w!�W�鶳���(���$h� ~{+���]�"��$R��[&�L������'��;���g}�tiN��V#�bԎ��,�B`W��pW�O�!i�h͆�a�Dw'+\a�qJ��f�.�[�~ء
������زM�
F*?(?��'�9������ �ʴ)�=zVQ�B(|��G�?奇(�r��$12�*�'AO./�!�Z�̉_wX����[q������r^6@	�&��O:�$+��,��+O�m���}k�zp%Iґu���+�Bs���/Q��[QK��~��̀���mR����q��t�G	�/�]�7��W%���9!����1��,��ѽ������?����_" �W\�~�(��4薺���*��]D��K:w�8�u��%%)��%e����*��P��s]�4��Y���k;���AB۲� ���д吤���=Y,?��z�W�XV�h2�К\��p�dK5�tT��
�_�^�d]r	c��-3�PX�P*��f,0"�mW6rO�7�l����OP��g���?�z]�1T�k�;�ܷ���� ��eY��GƦ4/>�8|+%T�h<K�@Q`,����%�{C�}���Xz[d5�֟�	���	⎟��~Ν��.X5٧1,�Ļ�a���xGRodh����S�Q.��m�H�,�
����FNe���u�A�b{�_k�����y�}2w���{}K�b�i���=���0E���.R��]�����+qo(�ڔ�_�"�ǝތ��sS�Պ^�%�!�U�J��{�FB�@ c��M���P�T�9Ǖu.���L�J!�.l�#v+I��$�-�-��V�cWvy���o�o��CM��<�	F�7,�g颾[���i?ع�xWM�E�z�N=�vW�l��NXty���a��hr�s��鹽tZ�3w1��4g��U2��79o��t\�T@̃"���C"oB�'>ds��)���7`��UlbMX��Ne�qC2���.m�Տ�����t���
#�.?#]�-y�W
+i��i��e��io�.�]�j�V���C��d�$W�S+�j0�VE�)��@�{H��C'Zy���)$��y����s�GĖ,�X=W�*��z�	��2 ��$)�K�rʊ��7�Q�s�	��"�Q�yJo"�u[�-�hC�o��2p�՞�G��-h��T7�֡F��A�=;e�r�+���]��t5>�$�H�s�Y濂|
��ɒ�̃I��m�oD�V�/{pwT���L��������̿�5?O"�[5E:]�e�X��������F���!�&"
�66�������Ja�[[��$d�ts�0��dZ��Ո�v���exGQ }o)��Ⱕ�$�#:��7o�p|��k�E�b>�\�4�x���>�с7>��`�,��B9���0��M$�p���_����L��h~@I�a�D���}�U^����x�����G��޺�)�7%��+w��F�P	�>B�)`W�]ֽ4�V����e��Pi*Q���jb'Y.���J�RT��~^D�:S�C 2��qz(*�=!?҄�1�,u��(�W���m���T�I?[�c�߀��/�B'�>(��� v��+�7�OI����G�+��V�=�n�.z�xlQ�����]�$q�6c��:7}���)32�	�3`I�$�D��ߏE}�a�m;C���5a$��N��z��Wtst���������q�:���TH2��G"A��� � ؉��?"5���������x����8Cȓ( ]ܨ���m�gOg���a�04@���Ϙb�	�'��)�y�兣VHչ� C�5oE�a���9
�<WaD�z�-������v<���-W���I�?G�wkL!Y��p(���ꢛξD�G�����7�����5&|�����Z�36�����=���֖g~��m�S��T�$q]n�����l�:�Q
��[���.v����5��rNw��u] ;f�.����x� ��Ql�a1���g���蔉�όx�}�D˻��@A�/5���8p�Zohf�U�{��ϝH�z��gM*Y���[��OD�IIK��]����Ri�]��Q�Bu^T
��Q
gy�ᐷ������G�4�N;�M50Q�Aϣ�T(�;r,�d�^>��]��YhK�⃒o��f���枺��e�m?>�WU�9�mJԖ�4���5�V��dIB�Wu;�(?�V�
��L�X��X��@�Zϛ��*�=\��VX���ϱ�V��y��U@<^Z�"����Hk`:���E5!Ag/9�C٦*�t�x�.{�w�|��A�<��''=�(��d�"�!AC;�������C�%ݍZ!D�M��F���뒞糯Zo��n��%��
o�ׄ�� oQ&��E���Z�~h�l�Lƽ7��pϱ�����Q���G�ńǫ�ώ���7��p��])�R�̮<��7<(�X)��#ˣy������"]t��6ua�ױ����^�b+-ol>�����%(ۥ���&�#&����}�O��ċ��n��?�R��e4\��G!����6�~�ؖVx��K������	���ď���֭��+�|���	�Np4�v�3Q=��T� W�b�u��{%]���Ȓ�>O<�~L�Te�$b��@�K����O���ʣ ��o}y6�DX�!�:��6��[��ؙy����S�4�%��p45�,ٯ�C-y(Gd^�`oL��4BK�T�6�-�+�y�}�`���g=�^Ld�:�@�"��!��YsL��s�@k�/Х�� �b	�"{���*�»��ګ��ZtK�ڒ�2Ր�ƪ
''���6u��s�3��?v)�f|�� �bI�noq :���Ec����|�>C����H7[^�2'���.V�ǿ�W[s\ ��G���6�p�a*���Z/,�,��	� C�x�P2}|�?%�ڳǫu�bH<M����mq�s�J�Dx�ڂ0P���C��5��-H(�OH�@�e�����L��HA&'8=_��������pL�є�c�YLr5������y!AR�a��X#o�P9c\3���a}��*m~�/�؝�kϒ��>Hk���G�;�l$zY�$��O��L��P^�*�7�n#���_"�ޱpl3η�\-\�Yfd@��g����N�S�*/���M�]����Mn��<�t�q	�t���'��!��#*�+1�ސ>�ٺ�ϱ��zw]�a"�TQ>�p��$酟�y��E�T�/>[	�RKu]2�lxL,�'i�F�NB���c2�>�-%t����ݼ����I5�~]	?�)��4~���t�v�ްq��N@����y�M��a�/��E�e-=�ui{h��Ֆ�T������(%�� �uxH��d���m���pׅM�Q�1m��ͼNR�D�%����3!�C\hϽ3���і�j^goB\W���}��X��*)�ܗ�,�3_��3�;���5��ʙm�/f��[.�æ޴�ը3�r���SH��˃�9y�ʚp���y����[�����/7��+���erfB����^b�-%Q ����І��q(@4\:l(�Gu���Z&/�*gd	��i6**�Z��q	��E�VE!|©�G��ٵKj��/
;dV��L�51��d����p}D�*}���� o�wL���a�g@Z����a���>1���H�9lt�N� ��?P������R+���C�hg=�7�[�V��iOŃ�u"���<ۋ�����O$3���5�����ۘ�|A�"ڜ���#%t�Q�C&òuDv�X�ɸ8.|ʶW#��l��A&��j�sT��>5�a%Rw`x��3������8�.��H�Z�9�%iǁ০�ݴ>VA�t7�S���;�![pj��z�|�r��OM�v�}zB�>N� ČYM��ڵ��u���U����H�J^��-I��9�ጎ�0/���H����P
U�Z�Igt�v�5�8�n�̈t�����q��R�l�SReS��O�^�P�E��IyƀJ�bط}��+w��o�!�/n�KG~UF�b0���h7ȑ�۝s#P\�Z����MbRT>�~�*�=�j֝[�iQ}�x�B��X�ݶ��b�O��:@[��w�����:+�����y u����c���q�2�۴��>�\�W:��}4�
Zh�ICS�n���Rۡ�hl����V�A�a �2�݃K3Y�&��uﲊ�{�'2ԡ��ol��[�&�+�SN�`!Z�E�9*�� �Ӈ�}�Xޘ)�F���dl����}�>Z�`&D҅�Qa&���{��c%ʝm��*0(E���4�/2��H��mTw.�Lp�P�mR��u��)]8�I�ό�Β.��P���ǉn� ��B1�Cぜ�*1w ��5)�S1��fX)��՟wN�K�n�Y�XcL�S�+�![)ǒ|�Ѵ\�t�wO^�j�z�Bx������L�G�d�p�s�D���E�'�� �;
����hB��������z�
�.
��ւ|X&��5~��|IN����,��,R�n#�tw���=�hLy��BS�\�'�1>4���]��&1�������ly<g��J	a���b�e� ��[w	jxf��x���%�gЀ?Fy=���f��HID�`�m/8a��!�&}b����3�	>M��2��w����ꧩ��K�r ۀ��K�r�N׶Q�%b5�{O�9��dq��zCK�i�;���\<ԓY(�-���l�p�|��a����[;%������(����7�҃�4䀙�a��p�Z�
��X+iUS{zVE�+�	#�F�Q������S�,$��GY4Q�'��1y��s3tܖ���b���\)(�V��Q������iN��˩�Mm�EB�S;'8��`����G��j<���G��MޭoS`�w��$������~Λ�$pd�S�i������f0�ug�61�9Cg�Yj}{����?�~��J�{:����˕U��|Q�Ka��`E����C
 ���?,Kǘ�.�@�p���H\��y�����Λ�S��+�.�i�.��._V�_�3�|+ ,��
��H!�{0V�����r�Ŀ�pn��˓��r���ŕWh�5�a����,++�a�Ǭ�)l?��!��"(a��;��?O�#�l�˝�:TP���;H��}n.�#ko���bU/
,�,y_#~ɫ�yN+V|Lp^زD:\b^O�$Ŷgb�y,����5e*<��;Ѱ�a�� ~�U����N���O�I2�ň�߂a��F��� &��z���,w#dK�a�1����~����9R����\�^C�.�@���L���+�-8�kك"Km�Km�qG.$��0װtG�=�飗w�X|�f��êє�Bͯ�_�^��4)^x� +圥8p�
�k�,�ؚ�D�����p)���娌���-V�K�^¿{�h{^���"쫔��ԭ�e}�����#v��Y�f~d#<�+�)v>���[D��e�tb7�DQU6Ðϣ�����<�o����X>�+�ն���R�A�?�GeM;o�Ȥtl��FA_��uO���\�Y�A���T�b0�8q�����n!�c�D�1�$�3/b�~�/<ƒ8�A$)�e3��6���l����h����4sqFHo\h25ҿ��:�4����U�WD4�2����8�ĺ~H9AO��38031�%hkL��Q��ݶ)=V��O�rhY���7j�Y�Fͦd�|g�� y�ZT|eh����nJ�ջ�mƄ^�_lQ0���B�w4\���߀�	Az��4�QF؈��梽��&,>��2�ɳCj����Z���zl��njpp�7�]��цC�Щ�#��x[��98���ą%.~Y�fj��g���xt���T�\��$7��'�y�<0�YĜ��4K^C���˪�v��"���

��s��Kc7�q�-=�B?~��X�P�p�@��L�&�HKY�Ǩ�z����Ҋ�X1R�>BX�Z��W�*��"�1�;Ce�+M��$E��	�2�GC�L�;Veb<q��g��\#*��kNZ�}��Dp��x[�n�x=�g���_�)=��G��)�\:,Go�8���Xߵ�A~\	���y*�wT��`e�#��L.u��d�T �2�g�B��8�V�W�s��H/����ϑ��\!�G�1�?!�>J��Ӈ��G��b�K
�\gT+WO�3A�Zp�i8�y��E�a���Z�������?м���K�@����|�zL��/v;$�k*���T������Gl��R���;���W�׾�����S#~f�Xl�`�ܬ��%*�p�9���P<���2�U]��9>B��	�E��W?W�	�6q¯����b|�0�w/�^�� �6��,���o��Q��������<m�)v�R���J��j����`�ܹ�q��$���49:f?kn�V ���٧�����_<R�������g�Ay��WTld+��7�(M�:�ɏe?NH�g�� �Ⅼ�Ww���g�&3tn�����k�W.� �11Diaғ�ǩ2��i��ߕ6_$�_4F���u�emf���t#M^��v��X+h4�
ظ�!��a^�� Z�۲���h�+��q�+5(��Hs��1��0�O���*��+�&�V��ζ�ۭ�&'��a��{����0��}|��>�V���\}�i f�p�y���)s����,5U�ˡ��X ��3�B��L9���$���[lD��������V�C��'nw����}R�Ϙ��SW��+Rά�}Մ��=��B�yb��d�J41��3��Pҩ�=�i�Z�-��c�F��;V*�� &l��R7hiRFeP�{Ǜ�3C���>��Q	��0���|�Q���5��"q����w=�Μ����J�KA�z�
�}L����@�f�W	qB2y�qt���uh9��#�� $s�ly�^��v!����sL�0�$�F.�'=�}��kD.�����H��?�����q�L����m	P �wp|-��~R�8p5�xN���������ց�I�Qb�j-�
���rXߍ�g�x1r�mѲR!y��R��J�o�Fy`K��@b�
Rݙg<��[Lq�;����	a��R�$
�k�#-�Gx���Ժ�d��1�]��W���F�� L-Ñ�K���CG�ͥ��Q����P�R%%���4�y�h�vӞs�U=���a���bp2Q_���2�Pr�B�U.�;�o �
"����h�P(�V|�f�ﮥ�x�p�8�C=덱!��J���Y6��4�tr`"��4F���ͦQ㘩S7U�(n�\wie2�-3)~y�
��7��8 $�����ӳ�S(`�>�[�T9�c*]VQ��_{�C'�[�K�3]�3�?�L�X�-���s��U�9�,wJk�_�U'�{�y9�[K� <��[ѻ�+�x����,�)'��ԝ��h>j������b�t �}�����I�����@�e�%%�%��؈q8Ŕ[�6
���w�q�`�}t5=ք��*֝��>zF�'� ~#�n�,�����/�LC����N���%7Y��e3-����C��e��"���I�; �����z���N2#�Ș*U��؝$xS�\�;!2���Y�H��ֳNsu��25��o��1�F0�A�қ$��_�&�w�(�_�=^Lw�uX�q1wvե�^h��r��H�1�5	l�./���b�{��t�����Vֆ0�S����
���k�Ą=/��>���̓�][6���Ph�j��i��d��7Z����5��auZ�^P�?�Ay���S���.�)�?bɿ��!���34m����.iK�xꭂq�����ߣ;�)�M�ڞ��H'�K��dF,Э]���Q��R���uOP3PS�¢&B���~��p��r���լA}�&��NX������C�#9�鹞o'@�����s$N��A�[�K���b�F���C��m��w��N��S 6����\+4X���}��*��j�B��{�itl����9+@ʖ��a Vm��3��8	�준��ҧ�@*���Mc�_<��0�sݓ�O�HN�p���'���� �:�x�Ol
җ;I��"5IY�  َ�6Q�|-;�$�F��D�����1H
,Gv�{`ߩ��n.��瞄=�4��`��3 �3�͝���[�ytz8�A����o�9hT��2O�� 0��'��rZ�tP�r���~iȏ�愇 O��
Y��잁�oK�� �T9~T;����s�c��{:SSX��=�Z��"�[��c�s��,�bΚHW/`c!�*H�K����?Xk���.a�XV`ju:i{��.񍼈�X��E 3������0�'a{�'�:��(�n���nJb��6�${�"�j�Z�Ȫܬ�������~��h	<�GV�$3D9 +��*�&6.����R6���d�{��%L���!��^=ܨ����9<�w�-���{x�ذ+�4@�0����h~h�C_����%�N�rr��k���ʳ� e��1��Bx��J���+�9�O8۲�rٟ��L�}s�e`:�� �;�P2���L[C��o�_��,��g�vj�L��:��>� ���S������56��Ô��2�Qo,����v���I�wM!�q��B�b{9��A�/�w����e�D#V��UM�R��$���m�1L%I|u"b愡������S'�k��x�g[7�Z�U�y�ก'�m�w+
C)�Ͻ��E~|�V�j��%�!	�Ί�GIoYD��a��';�B�e����e��& ���8NH�����8+�ئ�e#���H��,W��D��~�nV�^��?�(� Bm���_������*nc�WF��pцx��{y�-d&y�Ⱥlp�OC�ڳ�����[��Ia�R�^폣 �r/T7���#7�J/��_r@��ȚSt�=.��m@O˲�\�^��HE��Q/��J}N�ͽ����|�R���*�^K��`��K�0'����-�!�R��O�^�Ǳ���R�]�M;�sH�Ma�vgw��;�n3�������Vh�q���_��t�Rc�<�Ӳ,qF�Ug�=�"ݮ�o��i�fb ����ͮ)�� qtњl�y�8�������
���q!���bJ7��2�B�7�����7aem#j��y�1�%=�N��G
塟Z;���� �~�K9<!`��D\���41)�֬3������b`��ۡ�GK`Pںg�����w�b�Q�t�ֻ�¯�l|��33��EF�����۟#�ޓS�N~�0U#�^��?��Ө�M��ɇM.�ǋ㖑��)<#��Y��u_z��
��89T���rf�L)+�&��o��>Ėf�o�Y��-�~�����hU���|a��s�KO0�&���%<��*;��o%��Si�À"��!p��so^�� Ӝ4��-�5��h�Cf3�$΢�k�E:�/�$�5@\�b���<�����C��6��٥g��/}�a��h�\�~^_�nX��"�*�u���{S(]�=5�Rp�/�y�����ĩ�p~�E�Գ4���z�T�?��N������� �H*�TZ)D�h���T͈�p֎���HI�I<Kk`x|v����'o��$8$��.L���Z.�:@�B���L<�n%�;�wD����+��p.��bS7��5S�q�_�c�Fl���M����筗cдa4�^`)n���j)_�DK��2)�C�Di�k:o���+3% fdC^KÁ_6�%Ff%y�K��ܕ

�ZB�������l#yŶb�71�m�?k����u�v�viE��8��qY���{��]]��#���ڑ����v#r����Ϙa*n����>[�K�zĻI�d��[�$�&��u���;ơݞ�����Ml%��~/�T�ar�:縲�|���ʣ��9�n)���ne)�BS]��=o|���,��G*��@� H�W�i��������0X&9�u�a���=O%���P��Ӊ�3L�;���~�lX�罈�����{V3��H�n}��ҏ��D\�bGo(���S.(������b����)�&*���@�Uzr�4me�� ]�¯�׿�,3���.ȉ^�H��a����Kβ��$�ٻ)���g�����	2�;�����J�;��T2����F������e�.�\Eq�b��/�^�uH�^ -�zݪ������"�pH`����\.uv�J=YI]
P��|r�{��������/�s`����(ǜ��NL����I�t{��z��Ci�����7?�����Y�}��3qq�$�؋Z.5���+S���D+�aG	���Jj��h�V O��4�������=鐄����''���0K��߹���W��˧���`
�ɾ@M[�ڢX� �u�J�������qD2�o �`P�;rV�ɃN�FU�N�b�<BM��"T�p�D+�%>ԥy󩭓����\�G%�Ξq:��6?�6M�i���LN�9�x*���v�l��)S�n�Vf}H�óH!#ff��5�IO��8C�P7Q��Bǝ�-�+��=��b��m�kn�9/��z,c�K.⦜d��(�lt���O�ĳ�v~��I�G�0�k�/���c(��<��HxB�1�(��̨��l�$S=l�[�0M+c$z��E,�������9Z��������5��q��15FSj��NN=��d�3��@$�4t0{�f]P��(c�T- �#_&��X*o�:g2��=�F��X�kI��~q+G��VC���R�?dd����>		0�*+�-R�B+���!�6=�5�]�7��&ТP�����מ��\턝DҒ?Un�������-�����`,|�ߡVl����ؽ��߮h�d����0�����=��%�,�p�G0C %4���[2�=������:M|9 3��6���g_�j�A<�TJB
�a��]N��À(��&�*o�Q�=aY���o���l-�NV�I�)�?d%�w��8�O�l�]i5R��Ԓ�~��ᚼ��J'�
X��V�*5TU5�n�3�'��#���G�.�N��3p^�A�Lj�X��v�3&����xN��R�,W������p�
��e���D4����!e��3�XF��kH�ȅ+#��{���
����� ���+�RN}L\��C՚#!�0���3��MI� ��Lc� ��a?=[�*z4� �M��Y��h�PW���?e�cZ�HCJ� �4,�hK������\�/%v'�$T������]�aG��-��Y�������#�9�8��}nQ��[&(b��<��!�O�D@mr�b�&���L���'r~�3ّ�&�T�]�v�On7���x`��7�i�)o��M�-2�a�ƴon �7��ҜwP%����?%.����B���	��Հ
�	9�7���䭐�?���%ۢ8��gQͶ�|��w��f�1����	(�VtH��������~��]5�����uH�p���ٰ�z
K��ø,�Ƅ��&������=���S܃nK.l��0A��.Ko썆t�@����J���6��Y��*��� e�1�B�`��{������# +�����*��:3���D1$�Ϳ����-=�=�^Nup����`�S��y�'&��'$�B��$aF�1���>2���u�rc���Z���V5S����
?]��:����1�J��w��~rQ�tr��s�b���mo��/d�:N�B���L���ZR�~�H��`?�j%������j`6������?�� �2#F���|��y����QaQ>9�\2f�Өڋ��� `L�Ay�1�?�S�m�Ms�l�b7?Ѯ�g�L�bA+�3�3$u�{��ۧ9,��2QW3L��$X��t'g��2��ȼ�J0�<S������q1�O	9c�-����Ѵ�:�C�S-����;��@���
�ӧG����������J����0��Ɋ��-������EX�l�����1��!��j峕��?����)U.:���c�h-ώ�
�ͤ�#!���mO�����,P���oSV~n�4�d͕Co,)�aeW��{��@A}29h`eȺd�p������{r�����n�"�����So�����/�D�Q!c��>����3	�=G�߷2(��-h�R�C߽[H�>�����k�d��H[S��ߦVr�P���b�&��$=�/�A����h:\Q�'ի��j��R��GP����~/Y
V#Vϻg�y��� Ԣx�f�����DmZq�L�c<v֯�V�N�C�B<��°�3�@m�
���	��Q�����ȥ�Z�ڸ��J&ٲoț���G��n�;��|a���ѰB�]���D>4��p�T&��g�VD�`Rtq������e`-nٛj��70S�V䂎�]�[�{<�_kM���V{"��v�UQ�������Di��t!Q�RX�Lv��V�{��z��[�YQ��'ƥ!�+��Q
�v���6s��L�Gy��)��{?K�+��DF���^�3�+��+*�!o����G�!��X�4�cq����t+�n{�8)�JΆ�`����Y�ho|fX��7|�t 
��<�x��UJ�g�vmL�~�i����͊˕B���������������4*p�'ʂt���A���>M��ʜ���T`��%+��,%�ZPF[l��"�sN�"-����4OB��&Q�E��� p?X���%�	�@(9.�p|\O3��`;�N�n"�?�B"���HrO�&=8�%��:�m��d\EJ�wtx��6����c�is��`OK;����U����_&nH(P�dI0>�3��C��E%�������ǚf	)��M�vϘ˸~F�W儁{i-�&©Pɤѝ�h����E�@H���6�ռ��^�m���d$$J���=�#Y�ps�e�kKW�T��G>�) ���m��mF����l��f�ʬ��4v@���#/A�N<z	�@�lS�Y�P3��f�M2&����hM%�4�P����R�U�9��C�R�DT^�O�\�������}���/���'��r=��BQ^*�uYw����"`L��H����q���T�����*^%*'r�Ļ�3���:����]��������~�����ʡ.��Mز���P�����s��k��*��^������j���R$vw��J�����cVn�2NQ��<GϞ�r��4�����[�D�6|��jJ�cn��X��D7-��x�_�C��=C��
�v�	�̄ɫ��~�+%�/����qP�;T�q���ZX�p&��xU��&ڊTk�~;��/Bˎ	Oxik*��m����-�&�[m˦33X�ZŌ�v�u�� �-��wQ����ȑ��	��k���ڈ��t��f�Th�4y���g�e���öN�OYF.ul��)J���m��7W�vB�Ϊ�Ӛ�"Q-�}\�G��s�h��%3c�kWW�5A6GA@�ε];�ݻ��&?���\(�!]v��@k��f�p�z�m[ �� ��,��\�[[��� mu��c�cs3C$֥�y��ht�N�!p��g�E0�x!��V��yG���2�{X�����6�L�w�Y�U�K�_��W?i��-Ղ�<����� !g�͎�;b}{�ǩ�l��g�r$�O�t�����y�Ds�ƚ�,���d�1oN� ��Qp㙈�M[�x�F���z�%2�L�h�
8���d��h��(dk��=�#��(��)��weO�"D�Fp�٥?�CW���$�\k+��!F�=`.-S8�'�ϳ-�ƞęL�����v1N������z�-��RB�'���׮�Jo&��6�bܒ��6���3�Ӿ�F
yJ��B�͒�� t�7,���lmG��ƻ�]*}������s�>�\�F�U��`7z�x.������>�`Bc
j�ɻ�z�E��{��.�d�Wk�vBwܙ�%B��±��f�_��l�ʳ`�A�{��]k[�q+����Fg�I�#�I[C��Oh1��]�%կ&.�*�6מ�~Å��f�S/*��v	�#HA�ѯ�{w�=Qe�0ZN7�ԩ�Z�H��x`߰��>��9�i�O��M[FZE��B�pT�}i��L�HW�6�=8.&��ݴ>��)2�7Z��Y�C�]-�]\��ݿ��|8��3�4����~�	��j#��Mg|�n�u�<Hzyq���Y�h�QY�,8C-ߥ�iP�;4)��q����d�J��n�^ޘ� �:�6��UcR�[X'=�%�*�K�U�Xv'j6�k�,Xv�#�<�7��6#�	����Z��x���:��m	>?�Y�b����tS�M���ÿ�i�����E�J ��<����+�5I�?[��d�S�"^�Qv�,�@�wȞ�T���[���vz>�i��ZXsd|��������޺V����9C���X+ڛ�}���O����\�6� ��,�9 RI��*[F~�aL)�T�۫<F�+���*y�/3Rط`��u57A8U9Ç����R��޷q�N��
�%�Zv[�I�NV�����I��=�1��~���v�>�PW^�p���o�{ώa�zR$��{��rQ������9A54C��/f��(��5����D+D+���1�Qy*��x۞���[��Y�{��T��K��u.6|}�D����3�����I��l�^��)��R���!&M]�������VU�P6��9U-�Δ��p��E��9�k��2��s�.�͌S������W�v��{�YV�,��YyN�2 ���a] '�������ҫ���Ylb��ȼu2�8�V�{i�k���]C�wBsZ~��Y���ݓ=�,��e�(�4��Zt���:
������5��>0x�(3	7;k#�~p�a��jV&�7F�]@� t��Z|麿��J:��6l\�H��6���:����d,��Z�����mO��Q����	9Z������Àd��\�x@%v�Sor��i��Y7VW����9�A슫~F5�`���`�X��x�������-�vط>����g�\cu>K����I�7��v��=��'��S�DA�L�����$x�v�n]��7s����������^��v[�#��/��%�%s��>�&�;f�-6<XjS��֏�7��k�Atb��M���,)�Ic �f7_Z�Å��XGXR�^�9�4���ζ��X�x�ϋ�9�fC��EV�����J��}�:�?��y�^ƴ���&��24�n|ޫ��A�X�W���HC?�r����ǣi�t���6����IV0�k�Ő��W�%�S��ron���J�d�+��)�ĥ��3"j�f�7� M��G�&���o��ֈ��..���S@ȡ�z7��2��Q��7�/�%�w�=CW���U��1�k��<�vxû뾼PP7�t������?��]f◺��BX��״D�1������iUJ5~�w಍��)̬�&��D�Nq��|�&1�{��x#Ŵ.��j�u51ר(��ǻյ���r��hû&�=�秲F;qm:�yJ�y.G���5��!.ɯ�W��g��bq)Ca>6I�#P�'�4��&#��ߐ��?��������B��ϑvoz3������W��I���s%ru��Twh���UJ�[v��Y�f�5Nls\�a W@F��k>#�wFc tJ����^UI��\�|z��j9��w�%��;&^D�(��d�6J�)y��)��1��k�0>J?[��a�SZR�\�p/��TO�(����[�*}PL��t���l��jB�Әݭ��w�scy����Z��c�3�KT�w�\v����[S�xW/7��1��K�)�j-,ŗe�JgG_�)�X!�2���s�J�T�/^H�O\�xpUn`b9\A1;�D
p�g�z~̙�+Ǎ�*��&��i*B/�� �|��B���P����X<�#a�(C1��ܩy&�_J�i�ijxs��I�V��xپ�($�L�r��I��r{x���m��B������9?�G/R��u)� �$��NM���<��M�*�/n|H�zyD� X�K`(��c5[�u&���L��-���Z��5�_�ꍡ���F5Q���Ԭ����
X�R*z��,1%�Z�����"���h���U+������u�8+N�T-ִ̝�I���:߭�@E���� �м��>AL�2�t�� ��Ġ���C0�J�l���B�����@pC������i��2���w1>��"F`:� ��y���I�f��B�!ef}"���'���FƦl0��o���?��l�x\�V���˕^=���z�5g�5�Z����]������15Jj�NU%����&n���"rymv��Gn�OJ5v">������(�i ��c��N��6g�[�8O����ˇ�/v��\���z�o�t��q�e�m�"��v=/Y����O������6��{�Ş�[ʨ�(oaK������Q�n ˻�S&D� ��j]�ۆ�$�"]����g�׏��O�O!�~ѝ��h��d�0H��Yڵ?��d*���֥x��x���cq8��|k�d������_+:G�d�YR� #��jb��a�g��Ю ��/���������6j���Ry<w53�5�X�8�b��K��ډ���$�~�K��<B�+5�׷u[k|-�,
����5"=2����];�]~*f��?PX�7G=�x�����L嵕e=��9*�����൳.Sh��3�}�F�<D���N�������Ua
1�R
rne�4�{��s��JO�޳v��z.M�yj~о!Nv�̝-�߄ƪ�F�̐�T�8��sV^6�H�Yv��c� 3�āN'���9@wF��Bj��o`9�5~k�p/.�?����[Hvf[ŀ�����ڢ�B�%!v�ibib�_F�Bf}���b%��	�r�О�}�!��ƨ���b���;�Y:<3��Z�JP�E^=%����]{�(]��m���q`�~vze��gz��)~���@��d@�J>Ӻ99������Z�� ��b&���g?7Y4�T.��$F#�����F1Q��4��m/o{������6D��U���I��'F��ߟ/^�2��X��|��]�۩���Q/I���m�Q��dH��+\j6d��DPa#�]H7�k��"Q:��*�	�'e�اN\�?S�y�x�X�x�����B���Ny2X&_�S����ߘi�������LEшIp�� z�8ļ\�~P˃����*�z�`�X.�䖋���G���S9~�n\�M�4X� W<Ʒm��;��W��x�)gW)��H��x���G@j��^ ��C�_�-���������!q韐y0�oWc5��ߜ��d=՗�O�-���f��9VLp#�H5M���T�aL�D���G
 �+v��-G�bn����C#y.�Ƨ����S�`
�43v;�2��Z�N1^ׂ��5G�wC"���u�xb��db�K�#Q��j6�Y���p�2}��R~�К�c�utbkx���P�06�]�CÌ2)�(����«?xd��Mbd#��<�mf�ixE��f�b�\m� .61�nt�Q⊝����w*��}�*p5���H�ǟa-$=B1��K����%�RL���{��w��1��,]�h-�L����U1TnJ�iѽZ�8�L4��z���<�GVi`{��S;8��*�JNlV4�;Q.y^���!	+�n�A�}v��kl0�0��x�S�1�i>.hj�d9̔Yϱml��-{T�|HF��O�23��,x�̱o	���l\JQl���z�P��,��*�c}2'�h+;�c���y����܈T`�*�?rD��/*�^Ȅ"��>S�27Y�W�}�a[쥍��e��=C
@��X�3>�p"r�r)\�<��R�j�hy_o����	�%~[��Ћ�H�"wQ�ː$6t��m	�����fY2PD���98":�P�/��=߷i҈���ۦ̧_�|w�ZRƪ�+��<�B�Z���홾�@�k�1B{ю���n�*�t0��J����WI]��h���	����5��t'l״Q��כ��p,��6Ç#�����%@ʀU��5�Sq��V7�G���xg8	�@7���m�	ۋ�Lp_z�����z|oe-��x�C��	}��'� e[���1�vC(�X�?�}�S|����	��g�����Wt'�ts����[��`)��E��1�`�C�/x�Wf�:���
m�N�>�}��BY(5W�MoP�VE��\>7	/t������H	�����"�H������wf<1#z��$��n�tL��}v������ğ��z���5�6��J�ك4�����<�O���lЂE�9�>�C�r�2T��/�@pf�Yآ�"�*m�[.�D�n+�}$�רp����:6F��+�	�М��$���+�7p7�'L��<�	�[n�y��]�U_�M��G��A?A=<`U.���:�#��qR�*��ߝw���"6�pp��s�"�Ƿ���*|��}y�U���G ��yT=�����xMF���N���ף]?�)���R��ZI*�	n��Y|MLq��8��%z�b�J^��%��i,���U����W�!���zs	�_R�ܓ��Q�{�z�>N\`���k�1�ЧDy�@� +��e4{�x��N\��)/�X`�Lh7K
g%�_ �΁�?��n��0�<��)�A����e=й��U?�>!ob�������.@��Gt�/I���1.���}0Z�Y!��<��|�9/4��b*��U8�&I�G�������[�k^�[�����ۉ���`XӔuΘ�zT��˩^�g�<�H#�r�fY 3':��5=��auR�J������AV@â�Q����d_:QG}/��wZ�����C�34HX��=
�SM���x/X��T�h\/�2/�s�<��%XD#;v:l��T;�-A|��N�ϺKU�6�wv�,���[+�NS�c�h�|�\�s�������t�hk��I��"�R�!|�F^�݋C}O�Z@4ͩ���/:��\[�n�@2K���*:�[YH���٢C��˙�	�>)��׷>�@����9�W�|y�C�@�(��=�ɸ��${���b�}����
�D�����?5z���\PfB�YU X:���K/17K�e��FIn��k�Hd�_��R=J�:Dp����7��ۀ��L@���풝j['�j)�3��fK}b$;�*ۭ6��L�����%zui�⹯gMO�r����4B�+.C��?��,�ǖ�I��Ҥk���_⃙t)P� eN،x��5Ǜe�{�K[�� ����'�٢ͩ�u���X� 黻�� ���MS��ͯ�6O��<�<�tB����p���fk~�Qp�˗�;���u� �]�=��2G��p,ߩq/Y�����|���Y�Q�2Τ��_�������ѯ������V�Y�������=���t�h+��H��*�S��/�l�����b��5������<��J�\v���Է�ށ�0U9��nr4���D$LL(�͌a#9��BD�נ=���k�s� d��4��o�P�]㨚��cf��*�a��O������i�j�?�?�2�<^�&4�S���cif,�r\å[=*�/f��u�O�`�F�"^�˦�̠�#L����<3�bn����"�5%���-�T���rI���!���\.15;����O�õM�]�}ly��;O�6�VR��?��56��9xwX$:��hd!���nԪ�����XY��*V,C_�
 �[Io�4%3bZ����_	F	�g�*�i���ϙQ���K�x�c��v�9F�-P��:�@u��$����) �+=nJ�&V��.
޳�ǡ��C�EVn!'گ���A�ngg�d�Ĥ�K��!��n�Y�X�S��B�EF���ݫ��e��&p� >�tƳ��7w�Gm]��5��Rrn=��Ʌj��'���0{�P����im������%��z�-٧y��� 8lͳO�B��̪���l��* ��]a,G���/r� �L,KY�}�T��E��}l��SoB�>����l8�������+h ���e��7S �7l�����
��muVZ,�zߥ��@ �Ks��P�`�v)��de��5*���-�j�!GN�f)X�?�+���d9�BS�r��4r�7�O)f�H��H�"V+z�xɺ|�?���9�
� #�o�'�����	N�@�X�))������or���R��}���=�]"2jCؔ{�r�aQ�����`�#>G�� O��74j���4��`�s�5����Gu^/��67Xݥ
����$%�~��=��/g�����K�(S���A��ulH����C�����־�Q��z�ua�Ʉi�i3Nr9�Q��m��i�?Zq20X[A������M�-+���n.3�|�7L�n$��$Lz��#Ǻ�i��:�
���og�Qc�F�ȋf��o�A�LV�fHb�p��d�"�xპ:,�T�`lR�`C�A6��=�;s��U���X��=��Ox8��6Lg����ތ��X;3�U���>�
�YV�_�+l�^sF5J��p�Q{�Y4W���'O짍}���'�0��n�s�U���/]�N��4��A�a#�J��;�=�
&����a
�E T2�i}6]��,k��p��ca&��Q���b�A.���C*ɀ����(���@SHa���Mr@��m���\v��12�]c	�Yj��AQ
q����7%@�6�*��>޼�:�B7/��c�dķ.�>��=�0�.3�������],�ez���E�`��v
Z����X�M�μ�)���]GAc��~�Ëuͦ�v�P�u����~	EʮA��>{�oD��S�����7BD�������6��Ѳ 6C������/�?�ce�t�H�u�)�}qN��ۼ��e�$��F�S;Z�E}C��j$L)�y��-.9�����Q#yq��l�l�W��=���׀.!�������2���b��Op����Z���I���4��
�b�	j:`����6I����ˊ
��ʿc�&z�@�,���7�l�n�/t��?'��R�j�c>-g
���`�a9�I �	�YY��x6�B`0�(r���I�@?����_�z����)�X���E[ ������K�������%�LC�b����d�X�rDB�m̘�TzÀ��Z�9���c��c�Y�!+��ׯ����xl���K�:�-�Kc��z��MD���	9��"[X<�کn�DWl�>b8h�N����N 	|;��"$� u@��5`��`]نp�slBS����1�:(mȞC�+FFD
nkI<A��ы=q�J��-I��M�I8a��D�yupN��]������M�gT��'�s_���L��T�7����E�	K�"��Y()T� ���'�}�&��1i�������Ɓ/�M��r�b�xD�L�OK��t)�d����ƒPٜ���<�v�{Fc���������:���� ��D�lS�q��\\"���J���A��=g�� �\Q���t��7������#�en,LHڇ?>	�s� ��7Pfu�	e��ں��S�x�d����G�_ެ�y�S�!����Il6�7�����6ӂ�)���8Ց��Z��z�YB=H���$ ���E&��I�����{y�����!�q���9��Y�l:I�U��^6�,��`]�)�Ү�?�'��л~�8������H���5�?z�S�R��O������z���T�������] du �ac5w�7��'��j��N�8F9���z�~6ݩ�.JӅ�LM�*g�xLoY2I��O��-���nR|2��o��~q�\�痨�5=��n�p���xR�:�S��;�L�u���&�)(ｶ���M�g  �@����%^�f(���1<��W*�l�t� &UܛH�8��XѹW7�����������t����ncC���*����x'��b��as�
�֢�t��>�Gv�Pw�K���b1�JЋe�V�m��c俠nM?5�"��A�t���v|j><�nRA�����aAC��Ba�Y����{�fYszY6� �)�[(Be"˙ݔ�t�4���N�P�����mk�D,ʋÏ|�!�c����x�%i�Zin��L}d��eo%&����kܝ:!�ع�>�8��T!.ݨx�9��^tm[��|�j=AH!�Nd�tCN���G��BM.�����U>���S�(������,ٻ8泬�����-�,I$�GMj�k��s�e��..ivz!�ֽ��	��]�\%��YS���7,��手ʦqY�)�a���w�t�1�"��+(X�4n������ق	��7$��+��n��c/x�\��������IB��V�C��vC��O���,~Ƞ�s*q�9<�!6#�vcJ���H��vc`�ؚ�U,����*�,x���Ù5W�6F��w')��q�'A`u�4�u2��i�΢łK7\��H#�a��U*���C�Y;�ҥ >3r8	���"{Q;���-��A#��.���@�~S��(Q�IxQ�����HU3�Ľ��3�z*��1�m�A�;ON\���R�T�~N٭I@M�x/Bfc�o���i�� ��F��)���G�k��G7�=֢./ç4�.���i�I�Qh��wn�$a�f��s���Ha�W�ѭ}-f3���h��ŵ��o�8�뷿L�p�s=�6���w)#v�|�bZB-Wr)
���֘��S)u3v4�H��d�$�~]r��̢���L@}]E)���[�+r�	�G�k�9�E���l��c�V���ɨ���D�T�}�����4n��������o�:��z�6/��_D��Fj'eร�c<}��D��t0�W�!�8ԩP�o�	�3^��� �|[p����n��U����R�C�V�%��߅d�o�G��](����~����$i���V'��@�،֫��D�!0+��A�68�Gm�n�+宿��{�&��	z)%�� ���[��>���������1��pɈ%�(�uxNO�ŭ�+��h�x|���a�%�Pݚ`ҁ�Ki�'r�WН-��5]da:���\zIv�6]��u�[�R���?tw�Ri%�P6��k�B��4�a.s�R�������̭J�U�=����
Qh���j����e�wt��:��il"��q��"Ua��%S�/B\�pH��^y3Gh>�m�CF��Gq �r�/5���Sw���i�ˎ!�����c��������zoa\$�y8��`�Y���J�ؤJƩu=Ը[F����`kZ�8t�V��?��4�Ò��l}A�^y�(wX�|[6k�d��*Aw�!b>�'4�B�Ѳ5 l�������4��+-�-�*�K�Y/�{t�G��t���ZD�z��A��6�ݤ]J,��4����'CS�y���g�+ƴ� ����$
�<t��{�v��S���	����d9c!Dq����e\�3ڟC!u� ��q��ߪߐ�X��X:��pgxߥ_�+���vE�b\���P�/��ʪn���h��oۯ����)@ߛ/�=˙�x���\n��DivU.�fu��̡O��`����R��N3d��x������=��J�4u��ڼ�i�s\����:��6?�
Z���4�lb�b9�k(,4|��	��:s}.�
IS�����#�p@��lI�WYu��ƶ�-E��E���A*3P/�I�Ϊ�>�w'j���)��K�x��<����@I�x�����D���]�� W�����.Q����-�x-?�\� �WN���7���OG������
��?
{f辬��ˣ��8I'黥� ����[IZ��+r�^T����knv�6�Gq2ϛF����B�z��&XZ��HV�H��?��X���&�F�����\�3�����&�8�/�8�%�~����lL�7�-��I�~/�������d���9j���2�(o��ѿJoY��������L���,.��d�����4��t�Tݦ	���&�Z�����t	:˕��6�0օ���h�ز�#���O�B���@dd 4a)q֥H��65�55W��t�����~�0�Ӑ�H�a�du4��#��� =�r�� śC)+^�C��]� ��r^�G�˺��+��F�$g?������c�,M9>cpM�+��E�C����c���B��g�����Ӽ)
��W=�B����~�4��յ.�@��nd�)����(���)�~�C% ��
°��FcL�&׮FY���F�s�K��Qݔ�ж	%\6�v�ےk ��f�|I"��7�!>
���DQӐ�袥���؅��˵U�
쭰U��Qi����4�߁�p���dC�����E�4k��2�K�tˆF -4ǔ%�Gz�L3n_�u,o��XǍ�~�W �V
F8��5�m'��Mv��Uv���u��\~�jh@��L ~9*t�'{9g ?��ws_�W��c[6�/���p��XUNh�R˕p�Qބ�yz��rv���,?N
 F�&�x<ʋ�lH���[IYc��Ʀ�$;1������Nyu��]�Ncu�<JD��O��Dv��E߼B
�y%�V��qV�跌-���i3���}|���V�>Q�I=�e?
�k��"{=��7)"�v�����  ��7�L���l���ź��ځJ��Q�~��T<��j� �n�}m<�7�I��D�H���Ί"VJ����&��0��"�q�0���]+밼�g�H����R��c�Z:N:�S��[�8��d��&(��-����5v�4"}�l$5�g��9C�Fb���=0�ϝw���~R-eV�L�YA\�.5pO����l����&9������x�U0	��yJp�,=�*<��|�n÷xdL�
/x��3U��,���]���D|�����5��8�*����ک2��N�,%iG�uP�O���}���]~-8�+��,0�s�9����>i�ڵRo�w��Tօ��?�dE \8��2�5�1�"�MO6(Rn�Vw<.���E?����6��e!I���j+0�?y���#	 ���p�s0�0�ȸ�G��a�ܘ�L�� ծ��UΌ���8ս��斶�'lxb���"fԏ����&�(C�[#R��U��#{����z��H)=0�;��V)��yCi���?��I�vyͷ�a��ש��N@/�rN��"`5OY�����%GwLR�a��7��d�Z�Qu������a�Z��B�\��Y�@����M�ٖ��{r��#������*DL2U^����%ǚ�P1�D��X'EQ,ȱi>jK���~�^DT4q��v!����[�f�1>�eN��X�+�����3|�;q�~o���^mP4��.���q���lLb 10܂�Cpj��P�ua�h�m���D�r�Ud@c&�}�/3�Y�%���,|7�N��J�g ��L�x�Ƚ�Z����QǤK�]}<��J�={�'�������2�0rݖ����-�C������S]���E����]����Rv�/�}]��W>�0"];��
�X�Ͳ��K/�g��th�z���O�|>u�](�t�,�b��9�o���g�T�j�V"(R�K)t��n�}���JX �;靖�����,At=1�L+��锜c^=]ӣ�%-K�:)n{����a��y  �<�A`�ts)#"�^�qѓ� �Z�()C���}%x� �M�{:%8 i#1y�C��"k�CR��"铄����S=SY��Z5WQ��P̞/�v�hZ#�u?�W8-�S��좴�7@LpH-P4��z�*H�?!�h�M��&��j�zpGcN���=��|:m�_][Lj��0߹�ڡ��U;���P��A=��[�o�Yf.��o Y�%��\Ql���eꉭ��(^܈H4�L���JDH���Ϊ :������rL�ˊ�Pؠ��]@'4$�n,|�muT ���~:q�����״��1�%����J9#��,�Qn��v;��j#�&x�R�����ʚ1��N�.D�rz�V�G(�+W|J{��=1�~�m$h��̗���J�Iw�ާ����睮
7�9:�;��E�������AAPݜ]��nW&�Hb��f�k�A��@.@e�` �}
S�l�L�\p����e���_����+��$��