��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����i��;ݏ+��ↂ0�?�ceR
k�&��;T/�h��HKIw�|��&3.��Ů��p�!Q���i(�+��gX]����\G��/"�TDV
x; ��*���1$���'�os�G́�C2�:>�r��]�#A��]F�~?:6�,Ӱ������4;Y-�����|��U]�Ԝ���6&F,O���*Tkt�Zzڠ6]�ޢ5m�IS��Z䝤����VX��@)���t�I��Ml�k�{F^��-���2#��q릍@�BF(S��:�����jm�â.]"�	�i�,��Z��GU�՗��5�P�N���Lh�����	"���>�֞=]Kd����;�'��D�Yj���I��Kv���R�]���}
�jD�Kh-��W��M�� 	����eD��p���.��8�O���lD�Wa2]8)�b�;p![��5E���I6�����>FN�,5��y��zo�����f�_p)���P�Ey������0~$��^F<)أl�Ϥ��uvLi�9���~�
�w�a�?>�J5f2����!ȜF���2���!�P\땺�G�*,;�J���U��#�x�jJ.X�p���7�`�̽�E�ȉ������A<:J��9�k83���v���s�0q+6r��D"C���Sr��/��Foz��r,��#�%��?嗑�8'�T�p�h9�7�d������X�)ݯ�|��!D��.BR�����%��� t��z4X����0Wj�P��Np��P`'�� S��Ym9���nO0h�4ڒ��[�� ��aq�ʋ�t�f�_��	x��z���I��t���T}�L�B�8"Bz@Q,�M�'?{+_��{5̞��QH{S�Æ��|g���JI�<��L$\�K=>�.E���V���o���f w�8�-���t��ޗ� ���@~W�B��ɋ܄x�.I��IjK���=:z-���g��� �'��z�j07!p�?�J��y�z*�� ��ʱa� klM��@�!�R#S�xSZ%<0@F��!�I+t�����kw4ї�[�٫�up^�q���72�Yk�B�M�)!M�S�P���VXN��]��C��۔t�{*T��H��vD�T�:߄W����d�S(4ج��n�q1��I�dt�#����SM����7�����&dX�2Yd�~�½�Z1��l���c�қ�Lw�!��O�_ 1�k�vvz7�=FE���`ϟx�iU�L�:q���1�u[�BrƁ+30k�ڀ��f��&G��$��wk�w�,pWY���=���H���$�M����4��N�� �^&>>{�U�f��ݠ�j�Q/�w[����B�Ѕ��Ыx����D�hPw�H��}����� !6U"�2�NT�x�JP�Dz����w�>�(�ý*���>kS%#�0�|]>�봧�31Wi]���6��Ѫ�m��f�t�m���o����3� ��ϯF�X0���p��,)���/pmX����zbGF=қ�-��.��tp�Cס`���O��]�����vG�}+Ζ�"����6�����/1,�ܥ{&�~��:���p�g�C�qj$��������Hs�e���1���ݔ�/�J{�+����T�;G�������A` ������<��3	V9G[�*P';�,�1�=d^�
��f��xl'�cɗ��y ����ٍ��4zr�KA�.7'�X��T�1����ޤT���3z�lT�T�l9�N~z.�SƬσd�M#�S��y���d0�5��ԕ#��:$�v��t�� >���!�c�ɑ� �#�'ڡ}
��#Mf�K�����$�Z��L�S2_��ᅳ�)Cy٢L�X
���_`o!��9�6��Z-�u�00W�:�3�K��a{Gt͍ p�_W`.���l����ru�ڴ6��TlD܁ݓ~�h)�RskB�5ҷW�w�#.�z��M
6-����G�Ks��'B�IX+�z*j�tߪ��`-��K_�퐄�'/�u�}�h���Y&����?��AɃ_f$�7�2�i(�T}�-����X:�)��x� ��>���m��i�����U<�ˁ���	¸N��hj7�QҲW:}���! ���U]�S���,���\GI\��^1��> �XߚCY��X���L���a/����l����j��Jgŧdەd(��O�mi½s0�k� �k/��Cc��#��7� A��l�Z���%���x\�A"�<ng�e����W�N�Ej�w�W�$��y�S�j�[�_�EY�����z&dF�y��0��H`oQ[�4��KěcYA�LĂ�S
��ο��+���m�Ev���1���ٮE��4�=,p#��x���~�p���}�)!�n��`�3�)[��:�N�����6`�B}�c��[4���"m݃��/��O�{5�Wmx]P�$���ʥ&'�X�l_�zzU������G#r�8�S�A\\�	�Ponc^�I6I*�����q~��W!��׏�Qz�x7`��-qK�*���7˱�U����l;{bh�Os�-:�ݑ�3+X_ҋ*8��h�Uvh��7�1_�}�����������N��/;P��aE�c�0D�Yc��4(�v����D�1d~ꐷ nԄ��Y�Lj� ɟ�6�_���?wM;m�;����4
`���t��w�2Pt����Yڨu�,��$'s٠�b0�9EB+�1E���O� ��t����\'��� {"�LeV9���4�ĸ��X����z�[�N�&��$V�n�F���)�GD �@	���9#��w�i=��Pl!@s�,S��{�E������R��V��ǳN$�����lY'��(c5����B5������P�4��\۔8�c�ɨ��W*@(�Q�f�6*��˝�B�	t�wt�بN!�~N߆c>� k0�\I��+��>^��ʩ����a��*�')	( WV�H����'��������7�?ulbX���[�q�~Ge���V�I5�L�j�5����Z�̽?�n�Ϯ�O��r+&�5�h?�Zn��j����]�2�8L�n% ǕC��Hs8�*��Y�p\4�����?��=���&Ď_��3_* 9x��+���1+a^�C�X�Q-2�������1z��G��]p��ʱ����UxdX���!!��r�I��#�8�v�����{�:n�!\L�%� �|���1�&�][�}���O�S>�u��>@}���d�����O��W�EpsN�y��3�Z_X���6)���9�oy<��l�UC�ףp��R8�<�J��hJN�:<�����Z�;�$=AX�k��EKLuO�U�L�\4ܟ��>y�Q���:t�A��|�b�J7�]�j�X�x���Ɣ&�#��D������?����賝���.��5f� ��
��@�*��te ��ԑ�R5�e榿����s����K���P�[%��r�.��V���&����p*�¥gH�k�ߕ�B\"�JQ��c�ȑ|�(�K��v��!gǮ�;�f������'iU�@�r<Z��Q�#���P�F���Nz��(R,�A<��7����$����N�"�r�p��Q�@b�g]�������Q����tS��C�^�#Kn���ρDU�[�gj2}�!<t�a�b�2kg�o=5�"�D�a�|9\Ў������S�#����?������p�O�*��TV�p��ӛo��>Tp���\�����־�s�S��������f�bH��t-H"�"��wuk��_��j�Շ5����Q�G&W��9P�J���RTDS�ϒ�����Z� ���`�vi��SA}��A�2R���-������t/����dz���~+�k4�P�iQ�:)��*����� GG�!��l�=�Jj�A��u�W�!ĸ��((��=���y?0ꂣ�x���j0slk��'hpt� �e�l��B��y������g�4�F�d˪71�_��n�ڍ*��M�qÒ��J��7�XU|�ֳ���"��8n;�|�������v��L8��,���[���L�����ү_p<P�zIw�,����`\��$a>����4��-��bQ��b%PmV=d�u��Nm��x���+n*�-V�,�T}�<��J�n~�������C���1�\�3��[�_�xJ#��_ޚ�_�ӽ�iţ"7j*a����: |�z�8���>���m�?�o�hH�1�=�Q���k�����G���?ɘ��Xr�<-�z/�Q@D쐖��v4��-}�SrKs�zX��k�)(�/���Om�����x�櫏�w<�,!�I��KVo�t��j�wXo1�D����.Ff���ApFd���l�5ƞ�"[,^�$�
F�e2X���ϳ���0�#�J఼�웋����p��xZ��z2�;Lv��ZGq�J�k�þ���D���j#\ߞ0"�<�QG9��5s��_.iG��w/������=��3n�!-t熃"®�oh��Ե2�Vuk�\KV���׶�b�[-������%_���d����>�4�4Y�[(���"��ˆ�q��p�H�
ovCC�KT�.AT'����q&��8�F�[|Ͱ���Y0��z;��Ǝ��*$q��I�L�2\��jY2���3Ǯ�'���+��]�oA�u2I�DGڨ}�N�C�m�� UJ�&J
O~K�n��<��S�0f?zT�66��	��\�S�oT�;%L��8�
��R\�����Ů��
��kՂC�x'�Pq��%.5>��[�jh�A���Ƒ�w�Ԭ}D��܌zZ�.O��f����c�F|�&��{�U�6�Ȗ\]t|�3�	���]�s�B��ϒ6]�X��
r�lS�L1��R�Hç�G, �HN�[�kC��QG_��**]�@ќ2��m8��8C4����Ѯ�*���`�i�p��q���uJ։���+����%D���Yv�����*E�T�r�#���ؓ��B ���U���bemί��b�ֽ�t���+.$��B�L�>����D+Hlf����4p�Ѓa��6}�Җ���تT@-^��f�NSs�;ChȜy�"N-�Xj��X�J+j�Sr$��g����(z�c���X�.sn:���":���,����Z�)��!&?�g
�P��J�a;��D�����}���P�� �b�j�����.Fm���s�D^Mk���Z��,q;ȏ?{&�?�bk?��"s:��z�s((�1����ʬvh�C��?
2���_i�Wk��d��䔑�Q��Pdֽ��O����r
�\�/�����9�e�(������
N�C:���c�V)�Ѱ!���q�F�f�g[*tT�tu��$pf�P�s��`��v;������Q���+9�V]�[1��SR�p���?�d#�%WZ�W)nT�c�1%P͌$˪��2���K��ICi��Yr����]; �����sEu��K��-��~��`��8�Ɗ=a�t��U>�8���T۳��z���qE�U�o7�����I@j��,��S���#=�Y�s-�n���f��M���d����v��� ���wZ�`Kއ��۾ۅ��]]H�����8�D# ��9?��"#)}������eA{��R���5`E8���ϩe�89��5d܉4J}fU�ba+;�P��,J��>{���e诿�l͠�#�k;�P��:��������?;�Bq� 罿�q�k�FX��"�2j�t3����2:o�
`Dd֌��y���S4�d]��u��H9?�A#ɞ��^N7(���J����6�
�C��[��e�4�H��������4hHO�Ժ�=s���B�����V� M�꤃��g-E�3�܋eϴ�q�n�	:�u5�Yb0=�5Prz���6(�o��r㝆�$��;����7ޛ��6����!}Id��'�%�q`"i>�1�Up��v
a�2Z���K�&'�O2*K=G��ٹ
=��d;!�4)+ZLmC/�*@�ۍ�U��7Uy(M��{�����}�C��K6#d�Q�3�� ����Qr91Y�$2�+D�
�cl���=`�V,ҫ1�k���.�
�k�}5�Y}9+�M��h���y�u,PK}�\��K�Aܡ-�-JgёΝ
�}��M�$-k!{ڴf�e�������n�0b���>��a:��R���M�۫/���92|����S�W�+ 4�'O�ZOc;��n&��((��3>��P���C�0��w�����-���H�����W'�z]]�NB�ah�.�r�������J,l�	U��m���t��:	�@ܰA�s��U���c�eg��4��i�@�r�Ƕ�[Y�!�˔���>CgE���b�=J�P���F�ߒ�j��f���,�b���{�f���4�E>��0M��[ML_ �`'tdr�JT�]G�:$x�]�k�X �3���<�������Ї'��Et�P�`���b����z�@����n��O�ͷ�$���RbBw�hn�'��>Հ�h� r�	A#j j�V߱�]U���|ֶZ��gﺃ�?��=f6A,��q�����Blb[��`��xu�5���#�/��p����OqЮ����v�,�_� �v�ФRW�v�cf��ʇV��u�7�����W_�	M������4)�|rP <?(���O�.�a攞J�c6��r�imp�Ŋ�ǒ�-�t��� �ovZ��C��*Y� �Mz�Ů��$ �%J��h��坷H>�{oh0��5WkY�¼�C�����Ly��}�%!���9|-���4},��u�g=����n;�x���	��|��">�Vv�I������.5�!��<Qُ��[tu��G�y��핮B+�pԙ?&�;�LtMiY2���dn̥�	��"�V`$3��>n��o��v��Ma`����%�SoX�C��i�`�9C�n�(ʔs��0��2�"�>��{���q�b�E���+�j�ou���)� 2>'�8�����t�$�|Y���v�x�0g�_����`q�5wb�D�^T�r��`f8��Ss4҇Qw�M�M��X[���F�7���s�!��왵5�#MfK_��	%�|�?����4(�����U��W(�|�1� ��+�iNb���˯s�h�5'�k��x�h�����h��䮐VAa_��42���p���E'�	�nF'MKP���	b�	�V�v�^��>�.��ؘ�^w�,L�G�%�}��ۗ�ƃ4\~�V����	b�qM�,�@~.��d)T��B&Y�p*�Qk���xݛ��{ٲI���L:��۲�D��ӱG�KS��-\�|��aL@�1d��FE�me�� �T�QM�\���SJ�9�vG�n�.@�y��p���f �
��i3�Q�R��T��Ĳ.d���V�� ���՜u�$Z���>�%���Ȟψ}�TG�Vb��F݀ ���G'4q�����yK<����^�!��WHQ]�R�_X�,���Y4}?b¢��N��ٍ
:�j֤qY��B�`	K#S�x���G�N�khvtB]�b��,���E �0����*����ى�3Z�o��8�����++7��,';%[�9C�z\�e=�/p�L��F���9�� IFƑ���&�LҜv�~�B�}��a�����eO7Q��#+?���v1������8�b��mz�V����L�Ϳ߮��b����='*��5�b'��4q�vqb����ި��1����M@�b�+?a0�}�=]�U	&Z_��5��vTt�#�$��]d"��nR��K���4>0��C6��Ou5dq�ӳ���̲��1���09�	٣���.<g���2pcj�3�8�02�?���n�Y�[�N��ƭ�[��96��Lt;O����@ͮ��v�e�[��gP�I���rs��Q?�R'�KKT�dZ�
/b�j zs�'�)J�A�ik�.�1Bq�D�+o�Nx��5���~Z��U5��B���L�0Q�tO�[�$Yssu�%)�&�m{�
����`p��ˤXT&,���ۄi.d��P1�G��1��I,��I!}{��NU�I/ꕛ�{�t���7ュ��4��P,� ��U�{���u�(���o=�r6���=�#|�B�f�?�V��N:�
6�������)�j�{G��m�v1mB ނ�r��+wo�Pm'h���Ǉg�,����Ģ�y6��,u]r&�>� ��n^����'Y�ߕ��o�G��VWNm�9���S�U:��x~����ju����N+�����e��`ZWg�t)�����
��y�Q�cL���
mP�q/-> -C���(��o��*�J��.�չ?.>/�|��3�L��R��~��I�[v��C?;����Nqkݤ¼�	9�G6�e�|W�I��
�E9��%Y~R$.�]�O�l�#2�c�D�4��4q��,Vx�%�(�z7�Y3}��]�Q�X��./Ͻ��*P��x�qLL��ZjMNen%��nkW��Q��Tr ��fGPD��D���2@�W3�}�� ylp��6��a������@�	NM}1$u�G����gEB��7��w"�Ϭ�'�F%�⃋�+��s���]I�ھL�N���~�����z�ֹ'�t�� K*�;3jf���]�U|�Ψ05�$��0b�M$(�"5��LсK�n�=i�)���#+?�J�V#�pX�!�K�Ǡe�>/� �~�,�.�/y;J��@+K����^1~���֏6+��M|�����b�*���<4��Ӽ��KgxW���������N�*7�RUrIn̊���ɉ�w����ĩ�ps��C����~S�*�G [l���2�Ԃ����d��8RKb-��]�������"���	��/$t�t9(�&���浢�4��Pq��9�?Ÿ�q^V��'Y`SS���{B =<n�Q(f��j�ٹ�-#a|p~�r���oWCT�f��4�����ߤf��p�ڀSE��e}8U̟Ybá�?R��6�d*���_���� �>T��V7X�]�g����� �־�m��ܾ�JqeL��1e�xק$p��dk,ǹ���ϟ��C�#/O��\j��Q�Czj����A�N��8�a��{q�TÐ����\m!+%�J:�H��4�.���$A����S�&O���Bl�<G-�vI���60cn��]O�m��3�tF#](1��Y߁�=*�2C����WK��i�0����]�V�Z�k��NE��LZ'�����y��d��l8Np����Q>8�E����E�Q���ԛel�쎂,3����g�3��l[ݤ�
��	���N��W����5�!��'w�S�,�[��M���a.M"����@��C�b�p#��`��R���#!� ������(�A�v�g�M��CVb��a�|E�����<ˇ� �EGS��y��4\kf�x��g#&���Q8[2���?����L,���̕�Z��~V����)#Y�b֕<ßI�RX�!�K�/0�	���K��=��ޑ$o�L�����Uyp�a�
� <G���̦9R<g�*��P��ە�@UY�|f��#a�A�ըh�&t��B9����	T�ޛW|$䅹ΕXp���ԇT]��:����$=cE����S�X� S�'?�����^�;���?!<H��V�8�'O���یF�]yѫC�n�k?�J�;¹۶PZ� kt �؍�puP�������T�.��.�5��m��M��w���M	�v�rkn�CƮ߭�;���T)f`H�6�> �l@n�*/����D��g?c/=8�֭D:uyk}�����z�|�,@S����4��;u��)bjyt��w��� �M������LC*�� �/F .���\��c�g[$����$��%T�#�4&�ݹ8�O�����������?ħ�S
�j�!@i$���1;�ֱ��CQ�H�4����/�p�W�&�{���%�a�����i?vj����x�%��my�ϐ]��}�V��a�5o�
�f��r�~�/����|d�c��(��T��L�(r�e�2��ڝk�@ �$U��'�ӃJ���`�<`�qﰔ=�.y�p�N\�?�.j�~z��-\Y�C�#���&\��[>b���^��%M����D�Җ�]�_ę�P��"	�������V�.�)|���X�z7K{��e��!��z�"���R�:m�ǡ���Ɋ.��1]0膟�Wb.����-R߀]��L�W��k�Ԭ���=F��f}Le>Pܯ�_���#�Od��#aȇORZg~�GH�&��2�U�%�O��?k��,�L�x�ϊ]�K�ߪ���F�k�C�����_��-|=i�N�|�P �Djm�3X�%�X�YE��
W~�Q��>+����T˼��ӹ������|��?@�|J��,(
8������A���nsg��gm$nr� 8�,�E�p�����s�+�1P�-s	�C+�_@
��<���`���`5Yl�#)��ü��X�q�M�SO���ox�,GZ��WD@)�K����q�Ra�n��#� �"���ɦʩU`��ѫ��G�-����*G7�W}�o�4���9��ͭ	n�����V9��	e	�_����Bs����\c�/3d���$�/�Ѡuw��:��"�ND<���1 ��H��meq�H��Ú�<	_?�2�����9��� ��㪎h�:�."��d1 6����AzL�2�7gE�
�m\)��6)S�?�i�z�ZeE;�w2��ϊiGNf�+��2��S,�/�I�b]�`\o:��p�h��Rkҿ9��T	(D䠈�)Bq��ɂ�v㮣�J��O���JӅ��s��C4I��-+��	8"(Z"pPH�����q�Z�5wHLZ'��d�~��-pZh�v������s�͙�L��3��`�#�pqb��Xy=��@V�����A�I�3R}����� �W����i뵩�C�K��C�MT�F�^Ԛr&f����r�a�x�A_XLϜ��gk��fQ"-��`�>����~��1��*�r��'�u}�$Q����i$�sOoI���
�?��5-�O���V):�}�Q,���*w��Rx���wunoǰ�bǴF�ș߸��1��䳛0��U~uu�m_K������Ј����7E�R��^9��k��Q�]^��h7�(����x
��^���U����h�&���t��s-#����Ю��L����\�
rM%u:�5�[��|�B��]m�&�˸쮴�=�N�R�/����DzIv$��`cy���+i}�=�=[�xK��c���TZ?��V<Ӻ<����i���F�9�T:f��Y8�GF}6p��fg�|����^�s��A7���Nn�K~�1�]���Hb���?J��)�)<�d���z�ܦ��^O��vQbEN��:��K�TE>�^J��E7ָ� ��H��t�O�BV%��X
VQ[��7��>�b�a�֠9�g ��v���&6þ+�t�o�A�}��I09_�������Wc=4��׾M�Yz6�DЃ0Z���Nv���S�4��/�������A>���@w�*;t�l���F�E������AvBV�������u;A�b������odk��|(�=Ң�ƼJM��ޝ7K�l�R��-��Õ�칍^\"�����s#+��Ƴi:_D�B�3Y���o:�W�x�l�)��`��~B/���85[�?1c�FN1�� 
C�����6l�!�jۼ��"��&+���'9Z<��흾�E�l^�K�RZ𶇏�V"����(�0�:��Mԣ�����B���!.t9�xU�e9*�A��hj�>�����i�D�M�l�4�G(�v:,�EՆ�Ί;��9K��)�~��Ni��漆]M�R�%U�UP��<}Cm��a(�-o_%�6��"5��I�R��k�v�A6���4?����{�;�Z��y���Nt�Y���K�Sa���g(���h&��hS����U�D�����}���Gm\�7� �={�
� _��ZSRn~ἎQc�/��)���~e�87WM����w�/�w�a��ve%k�6���0;3�
z"��5ɵt�#e.z�}Ǣ#���a�7^#�3{�_��3�8HOXW?c�q�;%�l%B=��@C$��?�S�WUu��'h+|�$ ���;�6�h8�j�����kk1����D����[_��C3��	���MUi)��j�����2�{ :yӭ����Z��%Y@�7t�b�)��}(�;��Ԝ�4#�Qu;�Aס;#aP�o;\��[��<CX��B����D.k�%���z=w2�g��0"*��R��So�i�4�n�v��j������Dǳ����_���N>⦠����)K3��<����FT9W;ZI��w�hĔ��(C�)�	ݸWp�,��̽ ���E�|�[)ᛮ�[i�~q��?��2z�e������o���'��Q��:�L��J͉W���j�N6lF&ۗϏg>u�N��f����Y�N��9uj@\ٚ�}��օn�;]=z��3����^�ț�M'��R����Z�k���/�����l��eEq��[���|3z���y%L\����ӧ)w6��{���}����('��n���,H�g1�C��Z�3��7�K�%ֈ�Ϫ�e�Ͽ?��R��&2�5̂��,~�Q�
����L"��yD4����\�M�J]$��#.����\�Qf2� 2)Ɉ_�D���G랱]�6�#�����8��n�7t���8`u�_��Ο�y���;�ح�pu'Q�z��X�{�'Y������i�!�SF�䉯�:T ���z%fR~�U��xJ��^XH'ADz�D�*�U֒��K<����U���f�j��%��S�*|�X�Pih��0��V�M\�q�;��}-�`������!7����`M�9�}MA���٣&�%Ǵ��W}.�>�Q�{l{%s '��g|�$��'�ۀ�Cq�ׅ�
��~���]'�1���mS$4ښ��]�������`�л���Q�ƍUH�@�m�Dv�ҦS.N�7Ց��p�)rd~+GJ�ܡ���ha3g�Ӯ[�k�����I(�	�q�u��r�K����J���Q2���2p�T2z1��ۛ��5�WP{�.�c��"�9���r�����r��h����>1E����Nng�w6�7�"F+]��pi7!&��d]<y���И�t�v�x��:@62T��/��;֗�*V'��\ePL�t���޻�yN�d�;�Ɖo�1������H���h��c��,��|:�=�-�}zX�Ȥq󏨿����3��o����|)*�Ԁ�R!�t��/��<N��?V�C~7ѝT�:� ��Ѯ�s�ѐ8U�U�u�#�/=���	�m�F����ĸ-Q��Lcž���Rs6��G�/�&�|��(���ۙ��2�B1�����S�����<d��i�t65��N&�ϩ�T�NV��U�Ov���{<D�r}�%�@�5�۟ 8�w��q�d1�/���(/F�+��=��Lg��0HF��<�IS&���d��T>��bj�z�N�&�?]c���܅<�Y����BWlqI���щ򞎧уӱ�D��^}�D�.t�������ֶj�i�FT�!�S��,��3|��QH0[��%�x��
�lK�m}�F%<����n�,'a��9�����C��?��d��7�6���Ÿ&�}�J�L�<^�7$��䕰����4���A����ِۗ��X`wƖ&@{nә�vn��+��0�v�K� k��7ZZ5�i�X��H�t���z�΁��9����Pps�Bc0,S	�j���V��r& 
΄FVJ�|��>�,�7+�'�w��:.짨��=~	�`x��NWe�M6��xU�7q��;ç�������k��~���2�?Z)���;�<��s%�p��w"o'�{�"]�9k���dq��Np"E)(�[3�Nſ�\��`9�(=�����_
�q�N�����ny3�m��2R�X>}5D��T���IYvN{�m���>Շ���Rz>l���;:3���UB�O���hQw8=ߏ�^�f/�K.�%D��C�K��9����+9l��r�&V�������"��%���y���m:D0�`3.��Z8T��~��ֵ���z��6\��Cjb�Q��ҡ�)��}���]B>��w�a����U�)_T�g|2����X���S�f�9:�ϸ��7n�,�"�ҩ}BU��n�`-W�t�RXs�)�R] �����8������)L�aj�:��C�Ҿ�3�VZN��}�x�KB���L��.��2�o��Q�bz2����O{���ːt�����Q��}E/�g'bYB'1�U�b��7�[��u?�$�
�V�{8���>k)s>��&߄k��յ�;9�����~�8ps�A��aaz��D��%���"�K���I*�b��ͻb'G�ww�b�1�]0�{���]&n��R�FN=I���y$Q����ȭ9�e���J�5+�	��1�6/��#7Cַ ��d��NW(��$ ;�T��zsrxI��X��~[�kSpט�W'�+Q4�-7R��M�DkN��4�:����#닓 �B���t�րܽQ"#�3Y�D��Y�%BN���vp��F��>qWO�KEfW��	���VNr�Ӣۥg�7.8c׽�8=.A	P��u�W�Θ�a>R�r`�s 9�纗�����'T����%�AZb�����De����6�:X��`:�nIN�2���{��[eJ�B�����dn�EK�$gھg������.�^�o!�+��1�\�Fz�x��FO�' ᛁ iRe����5�uZ��N��72ݠ�J�����������A�n�ƺ�[���}�s��=�?Hw�r&��d�Ps����S!��V��@��'R q�l��`��/�~�=�dʾ�}�z��P����Q-��|��A���8���z�ۃ��֊X�S����	p+B0����J,E̞Fn�B�e5�ʚ�#h�o��ak�ޖ.��8�!����~��[�A��zX����@���1�~��*\���,��u��/|)H"fG�`��as���"� ��\�-vp��qc�uZ�U��&��v�`#�2��j�-�A�fN��<�EL@�7���+�����KA�A��$g���=�/�d ���QĐ~./[%O:�"�
����m`���Sn�	lބAw�j=AX[oLY��4�n�%
c��'W��Ph2me�P�w9�>��6�${��@*H��ɂ|=�_w�՜L��U�c�:-�x�����
,f��u�N]���E,6d���/��&��z�7z���<��f��9��)�(����/��Y�'�] �qm��(�<��O��R�|��Ɗ~��V�ɱBȍ�#�j��Yx�x*MMI�;��ۛ��$_s��1Rؼ�G��`�l�=Q�]V/��i�һTG�8�h?��B��	�2�#�pIX�WC#��=׵�"��B<��&�^���msA;�,������
3-��&�>	Q��T��Ԧ<���`u�t"��r5��\[�%�`��s�D'�p�s�p�Ƴ�{>�;����'��X��� ~��F���N����E�]2��m��3)E��̸oH���'D���ʅ��<w��� ��Dc�#��U��-C�f�&����|��������� �S�F��*��%i6'��p>��;f?�a��*�k�}�7�n�VBB�ɕ���^��" ��[[>�;_\��f��-�ma;9��;��?��tE�"<ll:��9�g��L���dn�yǳ��b,l��H^C{���p������֧M.(�Ce%E��7ٍh��xĵ�:�H��ͥ�S
Ϗ,V��.�����f��4ՙ����5��fl�|י*&y��4�M&,H�ѿ�r�I.���1V�O 1H�m�#�o�����s9[/����y��	kw�h�&�&to����"�_���&]���j��@v�Df��mN���0ظ�<��l���tZ�8<ߛ�M�%�s�HM{a۟x�s��w*��(�Ya�Hq�c)�[�}����j�����h07��?�P�Q3^ig��f����Ɯ�3���힌����.�+�΂�!L�!�$�%RR���y�,O���5�,�f��D`ԃ�1��$��:��ߎ$+ku8�K�\�-��.�7�̳]�%���C˫�´�u�a����ca��meK�����H��`qԔ=:����h�Q���]���+�f�{W�M#'QD[��H�A��=��ۆ���'����0=%�!b-;���qvj2_\6a��@��������T�dE���ܒ���ۂ�*�pb���=&����S������$��'��C�0�O���� 4bZ�\a?��s��u�VZ����=���ܟcu=Ԧ۷��Y:C	bʹ�M1o�IPrO�n"��*������`�k{uGB�)�6� ����2V>U �R$av���I�<[Ut�׬�Y�q��y�p�T(-lM<?�u�1~K�ꁐU��ƞ��G�E��@@�бjB��x
��A���r�ah�5��'P����햼��sѿxh��2$�^�8:�����~L*�O��
8Դ]ƴ�]z��r!gPx���7C��7f��ءn��r��l���8����������{�,�w�]�&9=�W�$��c�a#��fH���:�h�+&X�#��]�g����C��s^�Cs�H&L-�J�49��eOUo����MV���	C�Q�`�c�t�\��DU�h�yw+Ҩ�ɢ�2%� P����W=����C#��Z+�40�K�]�v8g_D p�� ��	�%,��-��W*P�L����+��3�o���ƴs�~�Ar��L����ŋK��٘�jw���*.;E)h�z/J�fؓ��-��^�$����� �2rV�ٸ���C���L?/�$�]��[�S���������Ĕrs�q���*8�7s�U��s�y�����&�ʺ�	�=3�l�ZG�Ն���m�hɌ�9I��='���|��b����u�9��cnx)�#%�\
5j:�&��Nx�}���g��� U���e��zG�϶��	���AO�D��o2x%��PF�+l�L�N�%V,p�Q�,+��f�mʝ����
����s����ȗ���t8���O>(*������{����2vy�R1�(�9��G�j�UTf�-F��-cTg��Z���-�o�p`>��5�
ן+�!���(��T��1��´�+6��g�>���Bѓ���d��i��.{�� ���@>�:��j�X���k����ai� fP"�T}��duN���� �H��ݘ�!b��JEHs�?ʢǯ�6M��>��8���j���6��WZ?������I`Q״�F!�{7���u�[��)�y��9/m�m&�TBg)Q�y7DG�\�o(t��O���w�W!�͉|��>����=�[z��}�8Jf��1����-�r�8�pz�§�B]֦��=�攋Or�B8�F���V�O��R ��ly�d�
�ܩ�5Z`u1m�.���D�X_-��\��9���O�}A�GC�dePYO��%� ai�*�ê���_,�S� ��fӅ�mn���n�)wK����1$N�G��MQ��������z/=���� �eI�1��A�z�i8pq���t2�����3R��W|̨��FK;wp׿�|^�(�*�7�����D��o	R�c��=��7��(����ȼ:��F����Do��P���e��
y"Dx��E'`<]���	��A4�Mlҭ���E�![�X�h�c;tE�X��>�ig:d�;<��|��?2=��׼ci�2W�!ŉ�?<�ACb�p�6��E��D+XI�t�A��+5H���q78���k7[3<�b��Ge�<p^9��w���Oڰ��� �MA�T9�MWn�mK�;*����f�{cF���	<�#;t�*Ay��5}뒵PDB'm�,��N�aaV��4�x,G{]�x���!�������J�3Ҙ�C�y��ӿuE�
�:ݵK�;�=ȃ'��r�/��6��7̓���Ѭ�zuc��k��i��VWx�f���OY$�J! ��Zy����?Ʊ~4R�>Nh+���X.	�?0{P�Ǎ�G���+����t��<r�����P�䮼�'+��7oT?�JLO��� 	X`ee���O���F;�W��
��S=��&ۗWۤ9��]����!4n	����i�tu�yMv˭��H��D�7$����"�5N��>�i�A�@���怙�}�!�H}�Ji�8�<�JN�z�:����G�HL�� ��%@���4X���e����f�xd	Q�|x���µ�|�7Kᕈ�����Uh�0;����$j��a�y^���g%j�\�(��e� |
�9pg�U!�Y�l�(S���X�
û�赇�b�O��s,�9;-�z�`N՝^ł�6�!��x����;���k��v�I NɊ/�R���4��HI�f>ގ�.	̳��hXy��bc�K�Y� }5�\(Am��_��V�)�$H:.��6�b}�)8�G�z1GE�;��bl��	i��T[�|9��1�xH�gVw��fb���<�A�����(���Ee��9�������Y~sc��>�M�p��ii~�x�jx����� 	�S���	��S_�u��3�5�6��	��*K��� �+�ͻ�N�����4�����:n3{�0��+��hl͗�4�@/�4�F��k���e>�1��_Fg��kP|m�#���A"�I_$N@��#��|��u�8���M�c�OÃi�Ԫ���N��ޱ�����FݘS9,�UX:!a���:�#�^�+ Ԕ�X�$���)����}���Pi�R�VP_q˦sh�=�l��zo���m����د
R��u�>�9A�IW3���0���j&�#���27�oN{��/� �C9����].��V�P�J�_GT�v���d_H�2�e�$6v݈��p�ot���UN��᪸F"�f]چ�wT���8����l�dϧh��b��X4Itkr�]���}|�Z��Xv��V��v`�[�k}�A���r/���f��F���E����U����k�7W� G;��'����\x����g��
��81� Cj�a�]%�����"e̤$�FI�8@�I�0X��!�"���<�S��sK��i�p��)r��S��ѵci%��s��$�Mu_�FtrC?��t�tGݭ�i� 5�.�4A���Z��[!��o��W�xN��q�;f�y����ni�E�Z@���x.n��������w��J�����$��2��*�#I	ǯ����;��D ��8�b��yS�2b��ś�et<"ԓ$Ϭ�$��X�L��I�xF�{<��4�Rx�~�d1=(~�{�c���T��LK*���G����{�{� Ц!J��4�؁0W��~y��m/h���+�ᐊ�Uꬔ�>ha��P6��/�*�v�� �PFQ�V�M�)'��F��ɯ7_h-����]��d��zkA�4ȾuT�E�_5,L��$���ɹ:�*�LJ]�#� a����*�1� ח��1�M�y㢕��+g���P⼿�åbŶ]��jU�ܔ��CNY�`+�6�P_Z�1g��������.aF��J��ɚQ��Of�5,�E��	�+���~4�b�c}�<�Mkl �$�'AZ���Ei������svTH���P��X�ӊ�f�΀X�RU�F�,BY9^6-i��BN�	-]`9�F����'K7E��|�
�_�`}]ǧ�r4Wm}a��gF��g���/��t�����C�Q�i��(���V4?�����,;��Y;V����F�=���7}~�m�����L����S\�C�&��#Gs�����V���iM�%�VP�I]ȹgg�Y#�F�b�~ű/�	` !k)����0�)H8l����]Pw�]�aW"���w���F�9*ѷ3B��ײ-�N��P��/�z{^��
��R1Z�n�g< vm�:L�6�8���j������6�(w8:d�����H�}Q0o�� ;+��GXZ�a	��L�n���Ԣn�/�o�V�Jv����x�%Sp�44�r��/�d���m dI�~c0����:�?C��f�#p�i������cd�4�v����Jn�&(�L���t�
���uN��w�"��r�(��F$Aq����t7"�F�s/�,�aȬB�*����
pKO��Й�<W���u�!�8��_���Yf��T[(87,̠ᤎ�.�,mRDP�'��63��X*����7�c��)���>���;H�%�뙀
�Um��	;���'̳���u�*\��L��}�7�T��!V�s �� z90D�gq�j%�Wт��D�,~mCrRn������t}�jU�vQ(/�o�wU*$�ǹtJ4����7����Ӈ�!n%�]g��P�' uKy�0�.���	��j/��a��EC�z�w0���[ ���'\��b�ݕODY�P�5
�Z��F�g&�~Lr_�x�8`juv���X�� ��Ȋ*�z�6'Ұ>mn��� �q��|"z�	9��?X�;IuV�v03�y��E"����_1��ohx������+Z��t�Ux4_q��Y<�)�����qx`$�XЕ}����#��\=���O�.#��n� jV}�7��/��mv{���t��h*P��v��%=�O"-O�]VYv�I������9��c�I4��ퟛ�#n�!�(�D�β�^�L�������C-?|�v���\����,D��/�#N�l��%�d|E��٨�؜�ֆK�WX��I�.*�&��@rH�b�A+��< *�ڎ�fy^ٌ�R�3��6��A'#t1]��Qp���mŅ��<����3��ԍ=��}l~����nd$�C��l�т�����{�u}aof��A��;Ѫ!�o�8ݝ������K_�L��{ז?�by�Oʑ����� /�Ƿ�j����h�5i��\EҼ�Զ�	�oX�̧kY~X�g�C+F�'��uM�5/H���l����$m��������_�	���y�Jtժ({�%��A�M������f�d��&JBkz-�F��?�����^J���D%t�m<ȵc"�����R --<�jhuC�����J���K&f���[n8��G�w�m_��F�<�nm��8N�����R;��a�����U� :\3e�yM%,E�G����Z2��{\b��ī�XE�l@��p����=�qI�_��o͝A��Xc=fi��K��� 4��(��{�Uh��j�Mc��%�)�S� �{u��U~j#���b�W�ŶbWW�EkF�տ��`�)�D�$�c*j���e�Hq�Z�xH�}fOb.� ���T=1jW�f�(��o.=2���� 4�R�u�m!vw�m��G��b�Δ�PR<�e�G����i)����"{H������b��5�l�_C;�����9��!�b��<P�K���VY$ 3��@^�厑MS?$�,.w��x�e&�ԣ#�O@�k2h/����:y� �;�e9��9I�h*�V�y�<uR�	r��0�B���t~;a��5ʏc �w��!��NG�_���q`�� �,���ǔ�W����o��0.��~�A�ľ��St�Q�_&ԙ՛7�C��SX��  �P���$����)��R���ד���E��!k�<#8,t4���s7ř���H. �2����|*��$�R��w#���s}O�����j�_E�Y�˸���U��|��g��Xt�	)���PE�L4|���GY���9)�O��DUi��ʨ8�ޞ}u=�q�:K�'v?L�}�=OI��#�Z��a��#�Z��$M�B��"�H�!�-�bB8���m0yi���D���9A~�8�h6l��� �v7�,�F�(���=o�@U��h�9^;��km�6j��j������T՛P/1-c��W q�\��ܠ.�14��!�	�$W&�h�tY��w�e}�w�+|K�� ����Pu:C�n�2��)$>CF8`��V��?tzWx|@��"���J.��#�����Ǌ�T����מ�PdZ���Xԑ�C�VJS�&76o�|�i��,�����~���0:����@^\���H��J����������ȫ��� �=g@m/��?N�}�TM���_ms;
�����n�f
�ν���X�=b���R��b��wK鸖�3L������=��UW��*@�Ԥ�Cߩ�=/z���%�?P/_ 5�b�)�WU�œQ�|�-�
47(H`r�u�� ��?��C.f��(��ͱz8���B��7�L���l��a�I�[g�6S��t���7�<k8PHf�SwЇa�Ar��Va5"��%�n��0�A�k�%�!~Vb`��T��ėx�*��m�f������;I�l )��F�V���*W�ne~���'��ɺ:��ԓ����3C�1��Wj��Q�PE�sd.��&�s����+�Kè��B�3��N���Usz��W�+�qҤ>�RA��y�8�xg���:�F���E����ʷшt����*�ɵ5}�g1�U�k*���wI��ML�jc����8I�޵�[%����mG���H�QQMP��">Z؋�oJA��	���ke��6���,��J�Ѯ6W��8U���	�,YJ�������_/�{�j�E��:���Z:�0�;� �&ӥ�^�~6� +��2$�6~	���9j�}GwQ��Z4�s
4�6;�T�p^H�r�n��S���=�	��4�œѠ3��rA�?��<�d�������z�9�;�Fxr��9ʈ�ٮ���I �@�҆q[".�2Ej=�~�(��-��j�|���Ho"ǀU�y4'�Cn]� _VZ1�,��gp��eKN#�
�ahь䝊�~�{md�d�}�X���9���ì��}8y~܋�-�t���v*ph�a�� �󱤬���4�Y�h��=�}㰕4��i̐��i,�T_���{J�:�"[�vե2��+�+�����y���K��y,��#�$��_/V��$�ɡ�������M)�����('�v~7�����)b&t�(7HMD�v��V��4�BrQ��~�"s,Y>����U}��l���e�\��qf��Wg���{ߴ�c��D!f�qH2��LZ���zg{�W��6d(� y�p����v���ʵT��DǑ��Qê��D�7������>t>�p�5�1\���*(
����Q{:?e�g�����4z��x��8ߜw��.��ȌW6�m]St�L�,��w�u��P��S�PX�+1�Z��y�T���y�� �q���Ԣ£8s:[�JF�=e����h2�t.���\62���j0Mʑ��*w��Ͷ�|�~�����"� ���r�#����kw��je����yG ��`����a�2��3UI�+����Ձ;?4e�VĂŤw�@W	�����.�S�K�Mt��X��ӈM�ZKe�b&=�=���\mȚx��SiX)'�L�lJ�fY^rǃ��z�ԻT=�����ʹf�`zs��56�ːU�P����{���Q��pEN3��塟";�`��C�ޙ�4���2����#����ά���i�����2�ksz)�A�\,�<�!ģ���Ч�V�#H|�q�oM��g�>8d:�o!�|Z�����V�`����s�	L=�����R��n�DcZ��#��l,hw|*`����MG����_ˮ���n�~q�>��!�zƢbލ�5�Ӣ����4����4�ї4��JZF耪���v>?��ߟ�"�#���;HmM�hF�ZN��Z~�ಳ��Du��v5��W��޸�P���ɐ������H%l�sv���X���,,�B1�T�T�[XJȝLQn���0;�a�it牃2��-��u�P��90J�Rє90@��=��0�b���&�:?6QND*\�K��x�n��GT<��E��R����\/�H�Bռ��(����\l�=����ͼ�kH��>�jj�,Y��>��(�e��R�^��+�_z�փ����M=1��(�2ð:Q�hCEH\!�r���|F�S�βZ2L��Y<��y�#\q��#�̠ϸD���_yI�{��sl�߱n/�Ӯ��B�o�΅��t�5`꾮Y'S�ؽ�L�Q+c��������#��& {�*�J���Dl�ό�.a(�)��8���0~F�����)����GP%V"m�T$��h��7� ��*ˍo��8T%�_�b�k_����sh-N�z��.�����pۇ����p��b%�Iz3u3פcutq��:+s���T�xئL��]�1.䏨#�F�ѓ�����SH��q'��a͈�����O^��yDr��lۓ]:H&M�<��VN�C��!1)T��T[�u"�Fd�ec���<ߺ�P��_f��PV S	,��lkhj,j\��
j�&�V0TY=��o�7�C�)���y�H�q��{��6�wF�������MK�/3�;�LT<�>7��|�7�T����1�����1�&b��&�P�����{C!���09g������t[��6�ʶϹ�� ����7Do !\"�8����?n3�Q�q���х>̡P��4zC]��HF����b��p��bp�RJ"��V�d��P;LqF.U�;��X�'أΫhղY���.s��򝏐�P��\�����|F]+�R�<(3��©16r��}G���3��.��ه
rw}b�Y�H\��ȋ��}�F�D�W����? ���䀧���"��h]�eS�\�r�PV����~ִT�٨T���B�mS�f��g�KfY��?��~h^��1��n�LP,1��@��{H��^�ʱ��L�m#PL}�%�
S	�+bz�T��(p <B�}vB=�Jz��cc��aLz�Zn�i�	̡ L �јI�fd:eG�PY>�6�"��z>�S�ٕ@�<>��e*�B����g��-k]�'*"~A�w�E�MN;���e��_r;셀�p�����om��?f��f�:��$�D��hs��n �ۓ��P��i��~���=��w��}�"l���d3( �|
t�?g���hŔ�p�t^��:�]Z!{Y*a��C݌����Aw��+q�����Wt�!�D����w�]E?W���?��~�_k��)�`�wJ�x�\#qQ�&��.���n^.���}'��B�􏧑�&	��N��_�n{��\��^Č��PӍ��\�8���}�X5���\CE�s��27���<"�Wnm�Hz7 :hp>1�$�����bV��4%5S�o�2�h�`����4P�*2�1d������͌Q,�p	�5�1`�Dk�L9��m�+ .��0��E1�� �N)]ˡ��D$���gH^*�s��'���p("K�}+����tP�UL��c����q?��^��Ӭsֵ��d.��q/lj��MT�pl�!u˜�dd)5�����l喗�\�5U�"�A�ھ� )������ ;%��k�D7��ג�B�{!�N�-��o�b6�xS�$�N�\��
b]%�t�;��ӧ/��Zmd/H���gP`�%���� �5��Zʆ����-����eǁĻ��V��h����_/s$��t�U�Ї� �#t5���2��\1��E�%��UN���-8Z�Q`�ࡡ&xqQر`���b
_2���ǹԯ$[�eC�w�Yǭ!�� q�38� N��A��r��z2?�15�4=�����7���0mTZ�9^ˁ�!��L��y�3O��S�v��Wh禕���v���f����C���g=�O����UFt�_���u��\�+��֡�6�!f���Μ��N4ߋ��3��N/�#�c���ߕM�t���7P3�R��D�6��`�!9\���g��ñi�~G�R���j��\�X��u��؏A;ʓ0���tVD	*h�y"Zi����O}]޼	'Ǥ��6�Ƕ�pC�"�p���̀$%�Wt�:��R�L��|��Eά*�c�P�@�(O\-���0����Y�Vʉ������">��������K���k0A�6�` ܙ���K�r�+�1���ĥW?8:~�����4�
��r����籞 ����R�a��X���C�o��6�	�B6n�l�x���iOg���[l�&{1��	@�%�p�`�RԇN5m�)Uߒ��i݆U���m9P����S��.�њ���W���������E%t��_�Ԫ ͤ�!���&~5�zh;�u~�A�WӜ����s�NJ)IW���(�s!ny�>�N���dO˲C��o�Ȉ�GW/i�(��U ��^&J=�x���+��X�6ۧ��
�mͳ����v�	��m�������vC�����h?��ˮ09$�ꢚ�V���*�L���H��%�3�z�g��j.�����d.Wt��M. �	_�>ü�q[w����]Cr�h+OB":�M�ã�F���gl5ա�� N���nE-���Q^IĻ'�^��t��$��aآ3U�g���� ��	*Ά�g��`���|�U��C��݁�L��R��?���pO�Y}��i%�V�)�ӵ�;��ghu�&d�q��y/Ҡ�7}��`�O\k.@�+d�5l3m�וx�|
��e��9���S�Snq0�B,P<>�)ae�����f��;�Vf �ð@f�Na�%0(�ȘŚIbA��=��M����$uf+>p�Hp�6����`)�>>��URicmI�pkO�β����(~���.ؼ�����P�"y�h��b)�k��}�m��j:�KͿ.�V�|E�<f$��Q*3U]��'�x���-*r���",��bț���p΂���e���̯�Ucpzۜb�R��C)�h�w�/.��?�s!�N;����`�<5�p�b5�1�U��1������h�\h�Ag\xvz*D>'m[	<�q+�!,}3���#e��{,i���Z ��0�t�@P�����3�tW:��8�� rR[L0������|�Aä�{���&����Kj?����� �6a5v1	}v�&`�J�N�j%r�L�G�i�Fxd�JfQ���,���	8�ۦKp��fE9�0B���;���������*Ȧ UE/E,tI�gY����R�:�9D���ϡ- B1����
kc��P��N�X�P��f�)���d�1�a�e���
��>`�^R���V317B"��h=��k8cѐero��އYD��%�A��v,CD/��k�P ���-E���o���qu��C��Ʈ�����ɯ�ڐ0>�ӟ�y����,�N���ڵ��ha��7y�p��;c��56��t���r�e+��ż.�}���'b�g,��B���y��n���>�o�8k�jsA��3�\�@�:k1r���a�@
�gz����=�tH*q89S'�1�1���Yəd��OmH��-`� %{�GڤTu�v�Y�	� E��#����te�j�"c���l�H�����x�b�����e�n���c!$���D���ſ;���ߖ9P��a���V+7f)��m��a��%���q�>?53�`��}M�x��򿷣�76P�m<�x0� �;qd�0T��弸�-+FW
�*���o���]s����fB����΅n�\k0.VG��u�oy�.u��ڐpW�~�Y�����'"#���-D�r��,���铧��|4[3z���7f�$�g͜m\0o�G`ʷ\y�U�މN���u����GE�b;��OF����%!IրV	GB�J�^�%<v��9Ł�;�g)Ê�?�J!~�����˫$���?�q��u�ڨ�d����!N�aX�q"��a��ϴ�ÈD�,���Ї������;C2}_/��`c��N��/�Y�p} \7�ƾ���P:*n�:���;�@<H�)�9M���FǝR���i�\�?�IkwR��]_��xX���D뢆e4��S2��˯~�g@[T��ua�t�W���r)��}U�~�WM��c��.�����+�WL _6&���}S�ԥ�F2�ش4���{ْ���R���S@�������wd�d5d�G3��.1�g�y�z6����� vH=p��u\�8�:����1����P�1�9J%HK3���b������t��۶��(�
����W��t���>��YhY	we+��W^�i&����䆼��y�ث|���Y<�H���̟K��SA٧�n�~��k��L�ދZ�sDݥQr�v�Y���!a.��LT׉�m��=)у-|�+0^��\��x���S�G��~�vkծ�$��lpYOP"��~!t�4>��
E�`��}���՚��Q��0ѱ�s<+h%F,@�,-�
	`'��2�����Zm#F'��j����E�%���AJ�⍋D�ý�p �@o��v���_��vP���-�.����v.ͤ3|��#5�e�q�!��G$�ӂ�U}�=��,BjO���M��*o��UaA�g��'&����!y��q^U����f���c鍥C:������O�4Y�2��$80�eG[y�.�'������(��eh��L�_~&��O&6��op�Ӄ�s�d�x���X��t@�?�h q��T���5�G	����Pk�?��L~Ļ�;	�����+���<�"�y�s�Xn�����vW9ԕ�%=m n�f�c��*y�<����:�k�����A��7�RĹ$��CW���*�� �����EQH���@������.VwG��i�V��1G!��)���]F����R�5�Ƙ�bP���,#�k\XR�n�����?'q�n��l��'�F력A��!�r�aVA��'��{tRSʹ��䯁� i8��Ĭ�^\�8k��K�z�n;W�i��?xUg#�=O������	�[~+��P讃����}Gg�ƺ7=�({m�΋�����[M�B�`®�c�r6G�P������h���<7�2�j㑕/��C����:II�e����9�h�F6����5��K��.Qn�0�ૡw͕;�~6i^o�T�$O����
�S��7�y�����NPu:K&0�4��������`�9�tϫ��s��m(���Y��:���P^�U5;��5�Y��gŚ���^�i�V�i��,�0��J$_;r�c O�_��3+N-�X��*JHl�XmI����w�Tn���'](u��S&ꎟha�c_	�b@O#,R���L��FU��UA�|�AvǸ ju6bn�!S^*~�l�����O�<C6#���/�vϨ�\�m�b�P3AqsH�H�g:�Z�
�9*�-?��?��f2� 6�A�����ɢ��,�}�OH:�ˡe�\�b��	?G���H��R|Iq��9�<W�*�y�W�@�B��u�0s��
��&����e�s;��(o�L�w]��_�O���Y6W2ش��,�&|�.��܇v%�I�ӎH�H�mR܃�n̔�V^�sl��ʣ|��������L�׹����+�c�=bJwz�0 �����]σR������0���C{��mC�]�ˎg:R%z�4_��>N�Dfյ�A�ޯ�����
��n왧����?��7#��Xf����zP���(�;������v�\��1"� nJa��[$H8����Q��/�hݑ)�N��{I�&�7��������0S�%�yY<����P=#X����忂(��h"�k�zop�Ե��n\tNP3ax�X�ke�E�'C��fG��r�t�g�I]	.7�ލ��*�� ���OC,p�%ŀ�G��\��R�� w\Rt��c�]�Vq����<��9O>tu�Lɬ����_5�3�FO��0CH�xQr��w���*�b�b_�#�R��w�`��@��foSh��g@z���h�A�{��/R����'"����Q�r�g��h4��idp� �iE�*N�m�4!*͹C(��}�/��/��8��0�����p��^��o#8��7tQN��g���=9I����5nV�琼���>�J��A��j%ɡT�׷��ዌ#�g|>�,Q��0y0
Ƒ�u�r�Hg�Q)�[q^>��
���3v����'<m�h|F�]��6I�+pJA�y��Rw��n���O�f[�}C�G�0�}'�W�j#:�{=�خx��6'�:w�챟[�]�	�jP������_��N��_���xz�ʝy�Ȉϖm"rlٹ ��C%��UjF�D��>�"�����,J���[#��ͳu�m��%��?[09Y���E�Κ��GI� +e�����j�]�/Q]����n���\:�s/����Uël�k|���}��jq�6\�b̛�^����D�R�0���6��.v�0��r��bQ�@�~|a;��'A���"{G�*�h1�d�c�mP�Ic(��O��c�Z-�q��
�?U�����͑���k�Ӷyq?8J2��]U���Ka#����SJv�bZ���|%�̏1N��b7D����	9�ŶSd��A�w�j��/��
{T���ܛ�G�R+X��L6��D�qS˰B?�-�`t(�u�;���El;Oc�n�_�N�c�Oє��;o�����]�ݠ'�|�3E��+L�n|�E���;�
���[�����&�;��Nfo��Ķ�d���]�Zo7e���fX�,m5��J��D{���1�IS&�������.��N�h#�I<�؇�c~�=�
uEL���K�_ �u����l���C~�G�C��g�HL��3sZ�^]P/MlL����kuכ��S�x
sӴ�$�^����_�!���Yu 	߻���?k\����h����Ma���"���j�+M�=�u;J�aN�{�B�/��ƫ ���Ͼ�r^a�S*Y�$@�6<d-/�41�k�RY^�9b,	�,�#@;�Ι+���#���Bஜ� �H>J���v:_Ji�l!#�0h�T��gr,"�r�5PE^Id]$��g��FdB�+h�
�v���X١�����G[|M��[�\���P!�K��
"�t��{��]b�,z�tA]���@sj��ɼ��A%H֩sI���[E��1o��|72��=����ZݵhAV�''H��ic״�xԓ�2�K9�ra��&�
���N���"�w��J@VԈG	�a�Wi��ٔ��R-��2i:��h h#ï�¶�R�.V#��]�z����&���,�"�o7�\c<�2WYՓ��CVJm�a����R�5-��'"�����}��4����ȶ����6�]rprx� �q�S����F���l��
(r_ �<'ͱ"o����__��?� �3��h+bG��-I�'�`'E˰O��!���Xk�'#o+��C���5�%�?>Q�"�UK��5M3y�XiV��P:���.�_
�