��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�z吴�)b���ΡrϷ���	�J�|56=�#\y��T\��#v+�'�]�7{x����89�!$�#`�E ���c�ҿ���A�ګ�ЯLd�e,�Rx��&"ۉe���+�� 6����5i�����+w;��Z�C׭%E_���dNt[w᷌��*~�羴��4�(�(�{@���X�ΆB���5�
�d:uV���J	�g�4��z�NZ�%(�($����3�ч���%�@J�����ʮT��r��� �cz�\�D4¦ǵN�b�g�<PW����c�,�$,��u��<Z�[�B�(��C�	)A���m�ZCӱ�ӭqW&XB1����73��,*r*m7��?�X�'G�	>�p�+�k�g�'XJL�f��|7��~³۳2�`Y�@��s?��qVJ�6�_롞(��I�&�|j�I�����!3߇E*�#2�xG�Qi��i�"�1x�y�����L��"dZ7bu��_Һ��ugT�n�rgU�ԑ��a�/x�=�\��{�_��&�mn)��!��v��C���Pz@6���:�o�j�x�B�Ư-C�3|f �B���5ʸ�.9�֐��F����{09}�uv��J�� ���!�N�XI�8A1O����`�e"��<�����j��H
I�Ƣv�΢q	<��9X�@W�;������=c��	����TE�����s��i��GȠ����Ř��2`.L]�,�[���	�h�>j�C?�"N-���b�"&��f��V�Q��\�_����*-h�:=[cͽ���ȿ���?O\��}���H�����Vx�>8���a�8E�6Um{����8��;؎O��*�3�	�eG�{������
Y�����y����?���m��o��R#E����	n��B��dԺ{�D�V�'
���N�Y�hb�׫xˮPQ�G� ^��Y���A�qBۧM�~�㈒�R��:[S�)kH=��n�Rz����q��2#j�Ss����1n�����Msd=��Ӟ`�s"�,I'���SB�wnſ��B���Ziԉy���σ"�ǚ2���X7f*a_��9������%QMO��M�rB�^Ü�z��5q�w%����Ě��\}Ӏ!ə��\�~��9!���ʙ�t4_-t���&��Q`G��>�7�:��On�X�֐P�D�f�S���	�Xf�(�r����\	_ਫ������Xe�;���ȑ�f��$��O7]8�+Ii$���(�H��a�
u��1����=�`��v�̀%�_�b�ub3�/Ab�?�\p6�_�a�1E �h�1�P�G��/s�sP�Ev�$�aN�mPj|Fe����y�X�hɩ��
?u�p��3��>i�=�M��iU6>a~A��ǿ3�	��\e����r��4]��2wyɜ�K��$�ćm�*G���%���׼A�����]�X ��4�J(	���BZ��v6�+>g��4?��ԑ���A�nph{��N<eJIa��l��h��Pl�����YI����`�c��<�����A�!ϖ.svs!r*Փ�de6�"����:��5C���W����d��J�qMuNyȄ���YP=��&�Ǔ5�2>�f�31��'�6���%������4��-�D�Њ