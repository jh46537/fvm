��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\�#��t"�9M!@eW:�Po��+?A�6Ej�����l9�kj&[d*`6?�`�Ib��a�Z�@3�:/�\X�!S��S[ٚ�P]��W|�k���~ �Q;���~����迣E��[�~8�N�S0�-�]!�U�s��6���*gYw�Oɼ�<`k�-�,�;�Ҙ
���FD��Z�E�o�R�,���l��V��`'Sғ=7��c݃��Q<S�Y�5��уL,� 6�xR'$�i�;��-g l��G ܏�5I)��ހ=Vd×4��N���MP�Yo1�+v#�e��C���C�v��rȀ�'C��l��DK+6
��9���J� L3�?߬]~�f�	Hi����K��B�6�j#��j0�m�֟���75K��S�٧F�v�3�P�����;��	�� ��fg-�'z�n��2#(�������`KU��u8�*�B�jg�ࡻ����A�9�ge��{�Luְ4�%�Ђ\�¸<�6�R�M�S����Cݮ:ۋ����ap3g��5� &����#��ZZ��s8��\_sN�ÌnQ�kX�k���ǐ��}�Ľ*,(���w�R��e�+0����' љɳ�Q\�z�;8�~�y�O���@�bF027�4)��#��I�����Uy����HP'��0�@�G���rʗ4�_R��Ůg\�F���O���#����N�ym�Ĭ�Ä��|Ԡ�`��K�R ����9�'�6/���`��BL���~kB�i�Ɗq�S8���r���вDU3���٣��곴i3������O�:3l@h�7���D��R�0��"Kڏ�=:aJ�[�ש���Z���g��F��z2h:��eI�1��^%?,[1B ���P��D:#����h�xCl:|�L��H*'ņnC���#��ɺ���0�*��FV��Yj�?m
���2�=�NڭϘ���)��cg������:���<,�׾�*�(m��B�`͔��r������l��B��`m�W��z�<6C$�xR����y��omL����If*�4j+�����H�#WK��(�cFyi�^w�*rg�r�L��pNd�e�X%�
�
�ؽ���Z�5��ki��~ >>"��[�]�Ĵ�O�{ �[̓��$J����)E��Z�*�[�&ϼ
ʨ����i�Na�v�z�k!kYST�a?��d�	�uk�d	A�tBz�bd� >��A-�}@���}��;�Q�����ٴ�Ǣ��Ѫg*��p����$(@��%N�Ri���]CR�.�V0c$Q �!����o׷��3^ֱ��l��環׈S�j����]Su/�w�,��K��
"�N�"��b�lA�x6:�\�:��O-��I]�k�ở	��TD�1 K@u63q�����<�D=��i���"m���32�{�t��zj�`�?���X`��&�5Uy�̗��J��W�W��}�_�ua��6$��<�d��(���n���.Or骣�a����C�Å�MZ9p��gec<,'�tc��:���	�Lԃv;m����[��� �C��|����<3�7�0�� �;x�#Z�;�Sr/�:ɩN�� �?(��7��q�F�x�+�]�,|qDL��
����,o^Lb-n��-`���;{B�U70n�"t��a�i߿�~�~�f_ið��5�9cC��>=*�o`��B^�y8����4ä ��gOF�0�7H����8 ���[�O��#Y6���E��o������[i̥7!���0NF�ap֎�1o����A3˪
��J�V�ZU@���`�l7Y����f ��_���`{J? [����?P���n�u�A������0���eF��Ǽ�,�J��p^<ތE��t�R�JbM�uh+���c��
�F�}]�bL���1xQ���xE���܉��R�n�~`�i�e+4����ȝ���|pv΅�_���<�
�R:f�Y�E���A�~���Ρ/P���h���o
F������K�n8��&Q��YcvA7���f�N 
r�0In�}e�:�<���$�ۙ/NF���e��`�Ȕ����P�!�{'PL���賘�]������Y��
m*��i��	�^�j/��#[����o���r��p�3��iBH��K�&��1dW�v����������x:�:�.���z
yV.��%s��G�N�g��m(�U��ߦW�����pa>V���M����ݠ�fv��L�adL��(|�����>a�:���b���bx:Ç�	؎����{��O�Ƃ���� "�m֚�Ii(�ﭖY���X��'J�%��D#�`m)R����������7?�M,R�=�%�d5X�VJn�MUr�8��29�<��qh�X�~q!-�ۣ��^Ƌ�%�u�Y�h�c����o[�؃�Y�(���mG����^�}��$��͈�)XOq��� �T�Z�����|nL���z�1>�gO��܌x}�}�!�{�M�� ^��T9.�~݁���=���it�� �P���������~")��r��X�ܬ�U�[��װ���� y�Y�.k�'�zČg�5���u��~َ�-�Ut>�g�b��_r�BD(Ha��߅��YK�v-�FY6EL2��[����tz��)fɾ��9:O��`����(*gM?�W;��hA�+,�o� k:~��h�����}o]�^�G\�P�	������_(�X�_��4��
�}I�Pw����U���aN�A��K���;�;DQĉ�w8)��*����*�����`s��E'���A�J4�oIU-���X���m��t�y�&_-_��5X� ��#�������&���̽��^��!���
ov�t
9��UG�[�Y��e��3�F��A8�g@�^����HY��k#q���M�t���;�ݧ�ui�"��*r���a"�A~}�rf�ۧ6cV!�{��ksKSc#�����E�G�G��"�yod�$y��/�����3;����\�wzr���s:�S�m��n ��Iv��F:eX�52�k��p�'V��!:Q�+�k��7�a��Z2ʄ�5l���vTȊ� �M�n�}qPf��HFO��f�h�K��{'��K+�@��PH޻�^(�ZgkL�qDn��i��}�0_c� x,s^Q�b (����������(EO���N�Gat��/5��|��( �<���P�L(�=��"�-�
F(���VB��w(d��<�}�+l9�
`i�(�B,��>� "�R�\��P}76���G]Zr3�ǯy)��!,6��1��!
�g��5Y5���-t��x�'�o[��=����8�z�u�<��� ��JK�Œx,��ÈP��j�S0ew�	��:�����O+G�;ª�$.<2�������:����V��Iu&.����R�H'��O�.7�.�<eB3� �i��\�7��j"�R���E@����:K;7L� ��N�M�e��\��ϡ(�,�)��*^�����ݼ���;�r6�� ^.�����4ލ� C�:�2��j\���/�-�P�*�4�{X���=�	k�s�:������J����#�9���o������^U���B/b=\��W�w-M��:kO��ͺ_�9[0q���hh�KG�*}��t���n#�oɟ�'�"�R+�[�l��}[?�,,"�.U<k�"�Xf��OkK�x�&�Ü,��;�7��M���c,o@�r��ά&PK��\�a��)�Bu�
���.f=k��N'�:.j���{���K���`����֭��\e�Z_�2%�n[��`*�\<�F�{گ�r
��q��6q�`���e2�Q�a���/�ʿ-s�:v�Qm��ׇ��ʘK�(�H�n�(.^�qYd��w������D� <�q��(RDe��X�f�s'�i9�y���[j����;#2��B��U�w]��5-����¸);��fSB�ݨ���}�k��I{)_tP�A�W{Ԝ�.H�]���J����g>�̿�(kZh���ڐ�2 ���^ԧ��E/0$��QZ������[Ga�+�L�7��+�ۂ� n���.b�3���>�	<�0 ���An�I�M�߉Y���'>$m�1D��b�x���zs7Y��bd��^%j/`��Po��X~�`�ݘ�"��]y�6�G�_�˚�cCٔ���֛W"�!Ҍ���jޏܹ-g~u0�z�:	l;��[���y/���yd��З��m
��Eۢv:Zb슚!x
�ߋT��/2f����H�������x3a)���8���K5i(��H0䋔�XrMl��/0�
/�ChĄ�7z���\.�sp�;G���h���U������X���AM�e��yL�"!O�	��Zt��A�.y��DD��y�1�����}�@y�6 (
��;�� ��_zKt��4��[8	*�z2�Jwz�NU� ���U��2A�'!�;Iao���*h	ΦT�P4��zd2@���E܎�"n94q���a�� =�7��*� s��,S��2ܞD*��>A���Eb�`��;+d�:�b�/����,$�u1�Z�M��(&8j�0�^��S��~,�x��c?����'�c�g�}�%�ـ�¿����n�W�ğ�4Ia���w��s��@_.8��fG�-4�iC�a��߲��ܩ��l���3e�'o>�y0Z@��7K	����| FyK�
��e�
c9�y(�@X�����U4qCX��R>�䑎�u��z�Jں�LUR���H���J��7��T�w�����Z��i�e��;�>�D����СS�W,��p3�y��t��
�1Efqr���ëv$ <6��y^y_>�<��'�i@%é�=y	Bf&UF���Ϲ�}zd�����0"nz��l!��B���"�r<ѫo��H��k���!�ʺw�l�cr�{��H��z�dC掼�sqmו����x�R�d��1M�~��	���vNN�<�lѮf����Ynao��.$��x�gq>�VhN�E�`�ސw-j4��|�]��@/ۖ����v�0$4�ލF��?�j��6*�p�G4"��+zn�n;��he�l�� g���#��;k��ƳsA�!��d8c��΀��k����ۈ����OY�`��#�G���b� ����&h�:F��b�v�O��XN�v�Ψz�SK�Y%��Զ�F�o4�C�y� /q�C'��Hɷ�(��Ŏ�<�`������/�i8���/�3�V���(3����\DMN5&7]mS����(h��1&���=0Μ����C���)!��nY7��ӡf��n�h�`��*3���D�0p=�z�̚�����:9ۊ�I�^�f�Wr�ͨ�k�}5��W�J��b�L,ʣH���G��*�G�|'��MY$Hh:d�����\h+L)n�{�|�@��Z���|h\t��p��