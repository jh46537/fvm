��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[������0\8�J_R8�C�{B�z��I{iE9�Ъ�+�x	/q�{̱7\j�2�/<^�~I -t����o��1
�Y92AY���u�)H(����͠,5P^�V�Z�u��rw�`P�tR!���	?vM�i@YY�h�S�i����ȬNJ�Q;��m�ݸgF��݃Z��^oC�g��g�`;�'�gA����v`��#��^��PD�{"�pnfN	C)�=/Sd����I�V���,m��k�CCQ�q�Y�����ٰ�]-�aʿ+���rrI�Ҥ5ՔY+�(���ae2�˳x@䒺QdF�4�D��f�@��4�P8�Jm��zÏ������bUO��Y����>�CO�e���݄0�BD-��`�K�P��v}�{L8�>-�c����3������$��X�~ ��=3�y�$�
�El1P4o���W�����VSt)^��o[���SmCƝyZ:&��񅣚�GYx�K��1����ĻS��֡)�*B�wǡN�b��h@sv���\��|�fw��'-qW�Gb$Ȫ�*b$H<�t�Ӌ��?Ɠd�?��B4�}U�uѨ4R��q�I|	@��Tm	Vs�G0Ֆ�쓖V>��w��Y��s1�]��ǖH�~@ȩV]W�e���&!���۲p���!�WT�`����L�KJOW�ry,l��Is�%��SLB8Z�!x���-��p���4�!<�2�~��&��ڬc/�V�|4�[~=�Jq��/4�!q��k�ɡ�דC��7����Q�[�0��A9]��F��M�x�}�X�}��@��3�<|.|��׌�𥫙=�"�vȣB$�4@S�Ez�m���B�xNZ#O��ҥp���Kk��_�Ã~�P"=�'9_��Q.��P��� ��<o����|+TZ�{�w�}�7l@q��-¸Xف|��S4��H�C��,��q/����yCD����q�/(I;�~��.V�� :~�̖�nb�$�Ǳ����S3�dWi3󩧆����v��m+N�G�q^h�.��6�m��ي��_�<���������g�*��d���bI!���Aͤ���άB��]J�l�u���D�b��;�����Y5����z�ǳ�d�A�P+�l����ǧ��rd��e`b�p��J'�^�J����b]#��E�֞���>�:�3D+#�#�W������9����z!���!�f���r�'y�����Y���oA�T�e{�X�3�	���7!�V�����j���)�|�%wl,"/7�1t�u��|�l ����������܀$��lU� +()y���r2�p�sF�v�zX�t��"D.��2+m��7����m�i^�_���(T�?M؜�ټC�]"���d�
=z����h���l �퐗����i�m��?)L�/"ߘ��"v�L_���S��r�uu[�Q\U����.Z��j��x�@Z����O�%uz��Y����y�9N���d���y }	��b�����n�EAỌ�o	;��5	����"�����tqA�Äۓ���R$��c��0�i*[�fG�j6[B�u��>���E����V�(���z�E[�U�Y�cƈ\����q2W���YZD_3��ᮓ�ƴ���>��i�8ݏ��u���������%]ܧ���v煨��S�GiII.������G�S������,��S��l~Зg9�3���	��s?�3^�$zT��?�+�?�rw��	'�@b��ZuF_�C	�eZ�p�(m9Z�Sw~��t�S�g��E��C�q]�d��n�O�\^�x�l�WS���[�:��/�6 FǙ�kT��j��*��~"|S�N����b�
��N$o-��Ӗ |�Zh�h����^��ߊ-?��K<j�u�67>R�Z:�1qo!6ۥЋZsB������B��L��P~.G��)�"��`a����
1ĕ]�%����F{�F���h�k�}�5H��j\�|f64��-�GTw�A��npiw
	�%��}� ��v����u<���P?���ea�y��}{���33�z��e/�i�4+u�^�8|��}��J-����k0�S�����̮1�Ώ��#%��fcf+���ķ��z��]��Q�X8&�U �ȃ y:F����Ug#�c�n���]ƅˑ" �%�\�t�Z�{+���޼)BB����e�;x;~	T��V]�>�L���m���d^�+��1��@��&�r�����c�%�h��x������Љ<�U!|N/�pzM{|販߄23h�����Qԅ�� ?����p�-^���C-o��.wI+��&W������K°h �XÀ����eaSwW�����*mV��P8��.����Z M߮���2�w����󓂱���k*�Rk*s�Nwz�x��L����;|�f��d:��Ra���jh�i!�gf�S��lqM���r���o���z5�6g��݀�u{gv������Q���L��Q�)�(Wd*1�x�8%�:��j����)�ٹ@avmS�P���"(~��?�x�<Y>YԾ������+~�sp���|���&�V�`G��O�u!���fB�m�������L�mQ��_Aҳ���8�w�-�j�Dl!��!�c�ߖ��4"��l$o�>V��9G�:æ��Ɖ��鹎�M�?(nM�@�{���@�2���C,�d����nn-j��Js�WX~���C��R+bh�vw�"����[�|?	]�:S�+0��mG�
M�١��eM:$�2?	��%����	(l.y�\;�Ps��(+I�Q�{�~qo��v�Ew�rЭhN;�I��.X��6aJ��J�7ޡݤ�b���\`��W�W�[��>Z���͋W$��"�m�r���^��`B׳������n3}O�QI���`˸�����/Q޵:�kd͈g\�`YV�=�)�QBZ�q����ӫ���/�%��@��#�����"��&T�����HȨ/7��V �1��W"\mٺ�^P�9�����3s�(: ^�Gs�ߌ_�
܋�A����i�F��y��.��_�Uy�Eڻ�A%zZSq��)#��]1X|��w@��'Z���nb��8h �j�#,z��I^xx�S3�Xc�h掬�\o�����>f��h<��k{���P㛱q��q�"'��CL_��[��q�	Rp�O?�Є9-�����s.�!I��l�KUJ�3x�w�IZ�߿��G����jb�J!>�L��ss0$4~�`�nmSԚ�l��1�^���y�>x�%�p��T�ϧ(�A5{��,Oa�1?䎴��B��E��9ɧz����ާ6,:U�)3O,���vƪf�錭��l+`��y:~�0��%�8�wiL�)��E>�S>ڮ��[�V�?�ծ,�h�9=X�6����pܡ��_	��)���1S�Úd3k�Vu�(��W-�1sJ�	P]p��~�7N�����Uϱ��G�#�8 �@���Y]
p���E&7G���	%^}r=A K,RDX��ܱ�}��\���:���ʮw��g䍀 f~m7M�����4/~1�@o$z!u�|���7����c\����!ӛ�s�/�����o�?p�V�O��3&pZ�o�9��H�W4��N�,�${-��q���%�׬_�w���Fa�VV�u0&�f�G��c�J�.^�큳����?����٩��#�*���- .�Uf�ea�Jm��J����=�-Y1�I�DA��P�^Ԑ8��N�|��Ո\QC.�_��8HEL�i"��>�&�0Вr�e��NohЉ�mʾ�t�0N䮂��z����é��$,\�xtY�[�Y��N�F������(�<�5�Ѻ�_�ڑRf����6q����t�yY�r6��	�hc|�3��l�>!�~����n#�Ԭ~�d�����cmǷ��]|���8�J�.g&�J��;v�O<�O|=5� �!��*l�òL���a2C^?|�Fh����5-�9I����}�2T(��_M���Q1��!�/"������Q�YA+�����J����$��/��4(FahSAMt�b�6�"���c�	���*yG0�4�sF�u.�d���x}8؊� �;g�������a�,|�H,������rVk�6�f�:�2��)6��B���Q�B�&�3�~�O�/�\*�|��tP"I�n�b��f�o.uV	�af��=�[?���Ly1��e�T�o=���������Z�U�J��o`�&��4ߜ�;��G�G	vpqANƿm�Bs��ڪ�6�Ƞ��h�W����7�F5z��#�ť���5�~>���&W=i���3�|���S	�}X�/�r�i�����p�f�|�sH��9&���,�F��6BRt�ߛh���|�U=<j�$���@qC�Ѝ��r���3�g �.`dר�Ѵ
�W�h��G��.�z�M9��g���-r�R�h���u6�3ܣ>�}�P�v�&�0���
9�y[2��'e/޶#����]�`�!��̗jS.TlwI�L�'����
0���%��J�o`�;�p�����BB�ý}f�G������w����.�Nn���0�zy���&����֖��1�ONb6�v�]��A$&���D^���y)F�*������0��I�|�:V�|+2�Uڙ;����az��G�h���mq��z跁��K!����8��>b�biSu�~x5�۷��t��Z/Z�۾�۳K�Ho@����Q��k�S������?_�R��yϞ��tL�����M03m���OR���Y�s��9aq%P��	�^�3����ڟ�X�l�nu����뫌B�/�@p���rȟ�Q)��ϵ��V���47��W���b�쟻�+/~�8����^.��%��r�.b���ӆs?��|�7��h��&����k��� H�FRG9h����g\~�'����p!#���\*t���:�{ 1`�fA4��.fe���[�;��03rE�^�7Q
�}xh=Sg�p�5g��+,��j�2��1��3��j���h�d~����sK{ݠ�"̺�_Z;7+cҚ�`n�j&w� �ԋI�iz�"X��K��e�=��a.S������ۃ��B��+�ǫ��Wý�hl�+�ܟ�f/�N2�]^轅D8F����+h�AT�_��I�<���Q�؋�UA��cB%�F�~a���wM��3����x?�Mҗ/�57�"#A�.H^�Yǒ'<]�0-�b����l���Xƚ^�k���A���/�>r�4�Wr&�Ml����4��F��l+Y�;EO���a���H��g��8��X��{?Z�O/c^�M,��v�I�f5�]�笩L/��%=>��n؉��F�����n���H~��9��Zh��YG䳾hpP�v���9��{Su��rc�h��)wS8��/A�c��|F��~���!��S�����t�%5EUG�$Z!��0r��0gH��6�Q�~�����#?�Jܣ��W\=��u(R����K�t�<�u.ĒF�V�f�
b�B@	=܉��C�$Q��=�g:R�&(��b3����p�p+����!�2�u����7_�J2!\�i�gɪ_����m0�[גּ���hh�{�X��ĿB�?��"y��A��&������Ä
��re����`��8ZΊ"���U���C2/~�"9җ�56�$��l���x�ҳ��:d+�!��AKF����5�G#�2���n�	4��%���[fٗ��d��%ZnmC�l�Ns;�S�S��.���!�e����S{X�:J���N1'Q�'����j��p��a9E�׹;�D}ʘC�M������%N�C�_WN�q�d�5C�B�GHJ��w���;��v+,ZI���*����3��ahl��mG���|X.�k��m#]?��@R�F�٣�X%e��)��g����9�S��OqF�&�-�*� ����2T��w�e�|U!���D�\�H��,�������/�h$c���!���̓�,q%�g6���
�H�К"\�k�
���A��'�[��~�s�L[���1p��R�ʕ�-�]0~�\3�	˅<�V�2���Ca���>���^2k��!�� �]�d�N��&D.����5��(x�ԥ��Z�<쵐(rFr�H;n`���cG�q�f}���2��:i��Nݚ�s���ʣ�������g���ahJ[r�!�W�3\"�ߦ����#+�t�8n,3Vi^$EmiR|�7��a�{�d�W;��="#k�p�c(ª/o+�U�!���J����ni�)Ln�s���G�;�̏�⑿�!�c���OG#�Ƣ(�5r��~�Ф�ˎ �V���脯����ߞ����hC��a����G��vc�x#�VS��Cb�L/�6a�nB�l�֠��K	�!�i�������̞լX��~�J��US�Fhx٥���]x2�����BHy���gJ�]���4n�-������1� ����D�e��������8�Ȃ���Wyc�Y�t�q�e�G�my��t�N�MRf��
�5���؅Q�W��TaA<=n@������ҽ� ��7Ɓ�,��,FaE�
U������tۍ�zl5��a��t���,��=Ѭ ����� ��P�P���y���ICw�C�h���+��T?��.e�ԬE�M&�z����X��ɱa��(��b��S��a��u��%��X:������o��� /����+׎��M����rRh��B�:D�����Ł���O����9��d�J�nX�#�o\L�Rϝ�Uv�����wC��F�|��^s'�6�Ԁ�8�1S���D �f/�j�>�����'n�6�+�پ���0 ��)\p� ͜�W��?�/��9z�ˈ;ۚb��L��X�Q���Ų�'z��kz߮�J��"��Tl��L��j�gǚg8s~u���x�/Q�_�N��=�2�p��c�Wǂ$[R-0�BR�1�y���Պ���4w�����jP<S����t�4�}п�H/��7�}��
����n��g!5E�yz�(0�����5�u���� ӳ�'���͟�m�U|~�/��D�D4����*�*5��]��\�*�� �B��A���<j���e�0���fj������
G�!B�滾ú�\����I�O ����8����J��=�
!=1���N��Ѹ���]��✾�5���tp1��j�LR��P���ɵK��?r�'�'���-�}��wV���]i��	$\{���n�ג�Y������|=�ᴉ�k����FXڒ�c�>�����ej Ic?�7{C	�=0�q4(:�c���?��R!���e�������PC�}�(r���#��Ǟ��<�˽�bydi�WIuTIY��7�%�R����O�5��t��6�������:�b��;�;�R��ћ��ð�>��_f��[p�r|0X3������o�\~���shn��ql%���_�H?�t�SG��4�ԇ��O�Wz�^Z.:��4�m���n፴CT�К ������<��}*>P�a�Ai1�Vp�el@���}�"E�\���j#@yߝ��#P������z��璆�p�SVI�o�M9�&����S^�o��M�7�[�a<dFȶc�%�c��݇�^�D,���Uj�1�d�l�����Z��@Km�+��ᤐg:\�B���j�RVnI�����/�V�WV���`����_��s��|�!����<��-����Pu�*߿,������ tH����lm!�/�p�d�PnZջ�{ű����x٩���D/%�<z@�}6^���b���y]�w,�p�1��H��b��{i��������n���R��_<�����2)�'�i�9$w:�Q�a���%�G�c5؝ku|���w�R:}v
٘��X��M̰$r��ֱX���5n�O�a��Żt��qN��΢'��?A��ڏ�4Z�T�0X�
C����SĢAmt
ld�*���܇iȃ�py]�y��5��.`W��n1�|�ͼ�2��f��R\�
7=�!"#P����u�3��b����)�]�T��B[{���f���2,����@����/F�Y,+T#٣��A	�Z(/�W�[�Y�U _hDb$(�(#���#X��d���
��W;b�i@�13��U|z̈́��K+մ�Ӕ�o9�38������O ��Gׄ}2���3�b�H�[�b����/��U� òҪ�Gp�b���ؾ�/FgX���'�s�k"|m�v�1��]���A,�|���H��.�渷9I�2�VE��9]pe�ˤ�����-QnFA*O_����a[u%���[�u3�z/j���@��F�g�X�U��1-w�6o����5]��U���5���;k����>� �6$N|�d�V!�����q#������֊dU�\;X$�lV�"�a"�/0��l����a��ÎU �Tz��KéF�&���P�B��n4���|�%�O�C5���Sx�!��L$R(�fT��i�Z��@S\�A�����@hL�y�0����#nt�fU ��S�`�o~�E7�!J��^/�Α"�5��<eJ���2���|�E�3$J�����gg�)X�2-=�o�Q[J�^W�)�*��"H�r�dh�.�XJQG�yU:�	7���-nƱ2����O�&�D^��v �f)�'��gkS�%5�q�
�كײ��s�s���/����?D��o�!Tw��̦�F��{���߶C`6�ߧ� ^j� Q�WHF��X�1| &���`UO3KgEK���2�ݨ/c->L��Ogw�@s{��T֋#%B�(�˝��:Zk87����$�۳���%Q��N�'T�|�q��Pt�����ȿY�*��y���g�]&����~��A� �1D5GZx�|�}��]g
���;X+�M)\�pء���BE���l�#us��Ҏ\:  �?��e��1.�aVlj���:�{f.p��Z�����lZ�8�c΃�(�3o!��^b�+��Y֦�B��oiB=�#F�rcRKF�$�*p�֣���������3�jZ��K6C���,���'�Ґ��%6�q��E��po�%�ۙ��<&����G��e��sK�L�Y���*�I	�d� nH��d��O>Mr�.�B�Qen][{'��Y�*��w�7��6oO
�����0O� ��� ���(D����+/<�-h��{?5���E�������0U��5����к*вS+�����)QF�^�`U*��"�������s��<k>^����Zf!v$�r�p�)�%3�B�
3I���4��[��}�f�QS�A뾄3���+�N͌UȦM�d�*����9��t��X%>t�%�3J��c��T�aOx��̏���Sߋ1A�D���J�t}�t:�@m��MVe�c�5���03���Y����22�����$]��w�P8���S9đ�^}��t����˭��beo�btE_�	|�0_`Q~I�6����ͻ	i.������d �t.oM6�oB�uK*<	3e!z����2����U� ��u��`J���G@�G�D���E> �.�~�8�v���y��Si����e>����D�����VL�ay�,��lVd�*�'4֨UW�QTzـO�j��oԃF>�;���o$���l�m~����[k�u�\6�"�q9P�]kg:��iOC�� ���y]�m��h�=3��d���=�d|(�0	�<j~k_�P-�d���lS-�ʈf-��'u��߼`��p(��VWEjp�����[B9w�CUX�&/��i�೘��]뮦%hY����0��H-Ȗ�S�L�VĀ�NeT/�pH/\���:��7�?s>v��}l�lVIH�f�o��W�|�<K���"��iR�:�k���M�Lc��� �{tI���n�~C�]��!)�@FZp��&G��Dc��8'�xȼ�F)�iے$,���D`QY���R�J�`uY=���������UJ' �%�7��3@?���a;9�W�+.�7�EH$.��kl�Z\�����R^�7��A
���j�i\��Q�z�
����}@��S !�w/�L3@8���IyL�O=^}�e��Q����R�
�:[7�_�(�l��sơٸ_Ô禾��<�;<�y�p�󽂷�_=��.������)l�F��$��w��I>�t*ey��nc���5IR�)<�_NZ�Pt�@��hY��-��D�Ӆ�����0�	G�j�SI��yY
W���6
�H:��!��c���qЃm�s��@�\�������F�e�#�J9�ة�QH�K��W�S>�b�zhJ|��B�B�d��9%w�&����6
(�ȫ�8ap�Y�nR�/��8F�)8��JQ�
]-6�F��eA�گ���T�2�|���05�ωɋ��cg�Y9��;}9nj�����G�5�����9x��ľfA� ũ��={��/ړP)�p�W7�"6�����+R��;L�O�zٿ3���NP8'�ӥB�Tȯ�؇�ǹ!b��)�Sf�>�rh��2<��xӽ���!d��e���<��[R������D,Ai`�3���Z���9ĕ`��vbQ��=��"��8t�;��m����F��!j5�ȴPoMVS�(���/g��GR�{���~߇\Ѩ䡎?�b�+��=�X�L�YHvT���Q��̈�A�%.HW8�5 ��kR��yT<oStB�(�_���[Q�-�9�H.��[7�o�d��]���B�����g.v�I#p�I�gQ�fR[0��!\tH�O��.��F���EJ��S�Yr���4� /��R�ez�ak��Ļ,��`����ƕߘ5V��ZG����9M����M}����z��5�ڡk8��p�x�y�;-o�����Jyd���t>YD�=�f�������#b�SJ�)*3`K ���>~�<3�n�܊k_Ǥ�i���`h�M�"�XLPk�+tt�+es����}Y�!ݛ�����I>N�T\eA���
��;������V"�{�4�Eq��"�c'�+��m�)Z2=�BE�!g%�0�U��ڞ�w\S	!d+
��9qDϏ<څ��.> U./��D@0���#�-��������'�\��d��wV98%u���0xse�JN������R��=Sn���}��T����X����㻯�����&Y��'�:�R���*��9S�	9�J|�8}i�@	��eK�gJ�]�߬�B�2I=k��ᖥ�[c@H�	�5�܌�n�|�P*�~�ǽ%<�¸�l��r�7���:O��Aa�u8������_~��.������"H�!䰜���B3��ϭN,v�[��bs���M6�>뙕�5a1���v��&6x/����P���OwaJc#`2W��0�&����e��/ɤ������0:��ϱJ�R2��E83nE��y�u*u�ZH��[(}�)�5��|A�v�19?�'�.��wȕ��0�YR�܅l�Ym�(���/����v=��"�����6�p;�3����B"�W��q�rkX�A[��K�����+�-����u,v%��>��*���JV�n�Z" �I� !�s�����r�M�Bb-��������C��N����k��L�B��`&dso�+K���+~��q+��LH%���@tܺ`�[�ȳu��̗3��M��d�H���z�N>㏼&~�P�s�S�+5`iZ�f�{_χ�>KH֗֩��L�J���8�>By�D��K�"0x2�k�(���9�^ڵIF�����9P�y:�������z:�e���1��~���^ǹ�1m�i�"�x{�2���zB�iy"�$���x�E��|?�5��e���[�jQ`N���ś����H�Os"�$Vt��7?�=H�î:C�*I�kLP*��WP*N6�ԋ[�h��-_y�Q\��(��UX ��'����٩uh��_��1J3�_�M���ʿ�W8�v�O���	3�&�����M��o�!��
?�+�V�ؠ�դغ�E#G6!V1�Bfm����c4s�u�K<��b͊��9��B�S� ����Vh�7���<h�ca�`DB�����TF�KzqW�M"q�,�MJ�H+�-ǰ���E��ԫ
�"���Ȇ�{�u+ɀ�"!�q�;�6?�&�'�oe����l+�U-tL=:���}~��T/u����c��+8�ߊ C��نa�x����vJ��d�
�mH�<��/�y=�7k�]��zO�w�S�� ��c�N<]���}g��ɂ��=q#�����6�q�p���&�������:�f��ۈOD>}ۡ���1���X[уP�s�[mj�r��!i�+IZ��)0KQ��V�j���
4���-:%�fW�P8Vv��㇗��$8<+����ƥ�:"����#�:=���ng�N�П���Z�����όa����uJ���иe�x��ɷ|l��!��wy� �g�g������w���L��#�G��?�� Xb��tEPA�5
&]"Z�z�Te��~i�����1,ޣ=�9!Ľ��Č��hUn!��B��&��Lb|���<�Y<�K�sn�3�^DE�~S41HH��#H�O�p/��|:����|��Q�U�j-��pH��=G�����F�	W���
�
��������'1�o7��)�!���U�n�C�A�s�5ɿ�;6L��W�h�
�vW-�l����E�L������w��P�}x��~���ۅw����f�M�r�:��>PM����y�Y��zZ�X�u(�]yB�����K<ڶ�x�p/m�8������o�Ē�;�sҀ�bv��q��|�����f��J�φ�Z����<��$s=.��P�ݚ��%�+m��c^� M4T`$������	 ` �$��p�㬴9/��͓�5����@��u3:�L��(f����1�}�>HKb
J�"�]*��?N���)�r��ӷ]V�W�㡑�(��o#�S�.!������E�:���.����H7<At�c���^J��&�ۆ_/��e��6d��=��z�#1F-+f1�*��}?|�F6�%��r�ߝF�cp�:�:XC8#���3�@�l��|m�4����2]���^Ӊ�j�RM�S�p�^D�%�U�>%��[ۗj{�-��Cʸ��0ɰHa�B��k]W�~kYK�v�I�#���k��Ԟ��4'�x\M�ʣF=[��+��S��Z)0��y�tjI���]~PfZ���+�YOd�۬SI4�Y����
P�u��V��Y�N�ꀣyF�"��&<ofx���̙�&�婒������N!͈����f�,�y/�L�[����}�F��XU}��뽠4�F0U���	K�2�s �}����8f�t�&u]	*�T����,���WZ'WW��cӕ��q�o�)���e*����`ߊ��7F
,��������D����U��e�w��pP��]�������}���f5����Y����q��M�*�<�w	S�m�[q���~�"�f"�?}6kwqk��؀{q��=tY��	�7/�z�mޡ���'�ƨ���q��߿�����W����P�QfqN���Ԛ,��\�i��.���|E�q�q'U��OJ��	|���a[!�:d@m��<��TZ�rK9d������2�ZMU���!+����M2�۫�xlq����؞"I*PH"��e��yֺ�t�����t|Z ��+��'�(��w|1�+v(�g^"Ď�j6 �RJ�"Fܫt6}�<��WƟ�,��ۦ�C�a�Cu������D�2P0%@D��V2̱hN�uHZ4K��K�y|���#l��ϋSS{�]���O}~�O9��<��cS3<�f���K��	��Aw��Fw	��Hi�uq�=���@�2۔o�oђ�j�Id(�/(��ht�d��;���B���*�3ds�!�B���Be��a5�Ei��B�Ӷ&*g��/�Ki�����-���-6K=�=��bٌ�"��s���2��B�ش]>�#�$���ǘ�2���yB�i��v�3VK"�0�Q{�=����ށ�y5�:�������fK������q�k�B��H���1��ԭf���E�OqM�h��1�+݄�A�[V�D�� ��[t��A/{S��L#�b��J���v>�z!½[�{%H����l���t�VeC[�&Њ{Cir|	?��Բ�w�G���	�Q`��s��������㓐��z�����tK� ����|�D�_����H1	�~$�*�{V�:<��n�Լ��T�f=7�ב`Ơ��T@ʆ�	4<�k�36I�!.��d��O���˳�k��<�L�+�aw~�rC8�sr	rߙ��F�g�3�GE��e1刊��;���HV��4yÕ�×���)I���歌Cx��@
B��#k����W�,������mH��8H���"�c>�r�V��ÄZţA	�$�bδ�on|n)�J�q�m^�m�2G!0�j;ڵ���-�_���)�UҰ%Zj-t��9Vkk��[g'��Wd
߮v�v[y �T��l/�D�q\n%�Ew�V/2\5���U�hZw~^���9y�ٟ�Y��Bd$;xp��J��y���ڸ��cm<T�����p2�f���&��D�E�}���[�	Sk��,Qu���u/zH�CV��b�*F�=�M{*bcG�Y�1�70U��GbCVZ�0�t�č�elX?o�6�N�ޑ܏M�>�
�;��M6K=�F�9i�3��G���'��o��]�IE{�Ξ;9�#�R���N+�PDP�b�N�}��W:o3)eVʋg��$���p��,��HZzYHZ���jR�H��N~�m�c}�~S~(�jǿ��hJ�%@ԭ�Ti�}��ʤ 2l(�`G�}���8j��>�A�HJ�u��c�N�W�.�ִ�`���ҥTҲ��� 23��!(6-Ǵv^o0V��Tox�EZ�3B���͠"A)=מ���?%�΢��~�?��ҺM4������,ط�Ov�S�fȊK���Y��1�5*2���o��D�P�5�@�V�*��U�_ܻ�L%�s Ø�֡�Q"]qi7NJ߼��
��1=W:��z�pD���d�_�BM=n���M}�+77�x����0
Fk��5h�������:��ݢ��C>e���i	�]y����.�����+�X�_'�~��+�Ű�Tm�T*�T�?�#��yhpx�6r�nr�z������Z�z?��w+P'\0�����|��`}�t͝<}���?��̇��g�v�����DȮY��j_� 51�����Q	�.�D�Z��Hu$h�?����9����@&<Z]��J�^� Ƚ~��4:v"�f7O��ue�rqx��@z���h�8�5wLe�`�����9�ϳ�h�b-U�0jL��ޔE#��s����L7jd -�IP��7�.�@���ǉ��Ywbq)ˬ�J�H_�B�ʙD˭/n��/�u��̼�K��`L�5�v�C'�
=뮱e�$~�>�|Ə{�ۄw$p�}�FSޗ����Ǣ����~A�}i�G�?�R���òLY@��mWۛ�BMR�T��K�u/��cg!1�DG;=�7�2��崑���X�����HH��֦�M�~�'��+G��m7t��d���nS,!��z��_�c8�'�\������c�i��!����I&��ظe�������"(1��[M�N�G��V�AvhQ�Q��ӧQ�������\A*fϠ!��cw��׿u�ǀ��U75��A���i7��@;L/UNH�����L�V�I��毠M��{ ��:��)H�⡒i�8�̺4��T�?7�)n; ��"����}�
�V��F���?,P�ĳ���>��kt\��/���l�0��In�H�F@�γa������8=Y@)�u��J�5S ��
��N��,#��|.��8�Z�w������=S��O*���z��u��N�supq�;�'����#mI���W1�n|ں+���G�� v��r��s�M����[��[�u�S��%��:�uG�Utm� (��aWq
u�n�Y����Z<GS"��<��T��/��+̜	�?��0�}l�Ah}��;�����Td����P��9;Z4�Z����9�{�\������k5-��xT�l�W�ф�a���Er��<�C�Z��&Q�yR����_Wfdr�-Q�>�X�M���I�::0U��a�o2[�pl��F>?2���H9~�*6��dJ����m%GJ~����"�hp�t���"q7�?�rnd'�M��N�0���>�v���@2['�[?HP�k���K�g��b{$�8��33ҿ��e�$�f�yW��އ���I8w��ZJ3���+�}l�T�Պ����2���[�;}������ߪ%�N�OH��2���ߡ�:�Z4�F�
V�/ǚ&�}>i�I����#{��5��h�櫨\Z	�w���l�Vx0o�(�km�B[��sӛ#(7#�5�I�0[�����Z��L�,p��Z
I@#�����T�>FJ�O��hl]��M���둼��	$?nB���F$^�v6�E�{�q���B�f��6�?��>iJp�rl����/E
/�Z�_*�L�&����7���^G誷픶�Qƌ�^ p��Z����j��2 ��� ;��(���/�E�w�+=�����а���ę
j���Υ� 7��|���Vy�PJ��ѩ�|�s��>�P^;���̡�@S�1�����Y''����k�%�S���\�O�6��W����$MIy�e�ZYҡ��O\O]�xN%���v.L�±ׁ���LG0VR�<�|���-ZSJI�Ϧ��g�?��Q��xڎ�~g������4��x��tꄺ\����kc�B����z��H��[w�9e��u�BmĬ����S���dw��$5ݰ�o[��'brD���+X���̌�I߷�l���emh�D�B�����^pSpl��h
�޻�<�;��2�.�XX��\![>I���9=|n����hGKS��n��j*p��I*0:��C"q7��>��M�sS]�j0'�F�l��m�G�n�"\r�w��~WS�X-o Q��MGY��E= �aV<Q��Z��%N|��A;\	fF<��ܲ�(��{[��㩬|�r�3��dtVK�dY����B�*�e��xbaC��8\T��m����M��5�Ka)�
��C���<'²?}��-5� �r��&�ʨ��j�V�r��2�L2<���sa��_BkןJw����/J}��]����G�K�@O�-+ۤq�ڎ8ѝ51C?� c�1CKnR[G���c��ݨ���XBu6����-f�R�/9�.W!��fP�y��ch�GX�N�j�%����v��GP�֗H�j�e㥥�I=N)���j����Ad�!�_xyC��6�����!o���5��6�A�J�R{N��4^U�_���5ϔ�{��M@��ڰ%�$�}Ob*�,[q�c����zv��BFO����H R�"���8y��M,HpA��h��K,"!p�	=s�����*�Sg�
h�X����8����tk�^��+��g-o�{�_�T}$[�vBۈ����W�	����&�C��P��0�(t7k��e��]Y
�os,�S���NX�l�v)ȡS����j�Aԧ&Uo�W^�ym����D	$A�6�:,w�"w�����e<i�[�9sIJ�j^A�1�=0�t3e�y��I/��ǅ��P�Ж{e���@k�&�9���zp wF���/�����ؔ�ڠ�q��>vbwZQ�DǓ�{�s�qWSz�x�I6Jg?�!�jP���1���8���y�82��h	Z�C,$�ڱϋZ�l��{��wwd �,%XE=8��Nd��--�����k"$�/�ԁ/�x�{.��eNa���-���:�_��;������r�-�$Vz֌����I=1�E��X,�P����m�!���@®۩L��VsscD&��}�Q�0?;���<�
zap45Z����3-v_���C�S�s��se�r�(9g�Im��{�����}�h�i5��u���g����LzG���x����G
x���.��=�F���������%k-f��H�9�����w:���Ňk���o���zK���N�li�LFc�h&�4�'�K��U*|�m��>��E���F]s9*�{3���޼���Ĥ؝$p�)�|�v��t�M���r��8���R�L~.�3+l��ϖ�iH,-i�u
,c6u�[��|3�z>�j}��CЖ�\G��]�7bzS7���Wzϲ�A���n���7��;��Y������*�k���W���aE�楣ͧ��`����o��uz`�͔]��DO���8Bq������=xȈ�7��նb]��z��j����2C�]�,��i�̨�5��>���;,�>���v�ý���X��d���M;��^��'�L���=���-���ŻCO��,_�m�
��	���h��PI�o�����_;b��B�$p���K�CN��/�V$�l��I�C1:~��c��'�.
�{/e�[u&o��n�0c��0L���o~��Ao����mO��svʤ��y�fCn�l�kT��l�x�R�;���!�H��b�M���{���}��s�o{��&�V�J^P��T��x��#�;���+2�V3��n���t�o��v�5�	9��õQf�i[�[l3 �9�Mg��X�z��uR"嫶�G|�(H��v�'�|�SQ�t�f0�
w�p���@K�Ħ�G<SLq�-J-u8�\���w�^,��\���`�a�986�j�ɚ�m�=C�T�.l.���U3�)ˏ�'TG��Lǿ��<M�ԟ�{O����t�+���<4�98n��~��|_I�Pz��c%[Q�W�do�] �1��O�!�ĕ�s��ܓ���u���1�|'���w����
kFG��˟}�/�<�_&��q����圍(7i��9"�ro��q4�3�@�4�U��K��i���l�l�P�����9J�[�ZP8e�S�AM�����t�X��o���o[ِ���Z�Ŗ#
ѥt��O|�z^��xϰ�k�Hq���|��ϗ�1+���;�y��/}P�7�g7�T����싢�vn�5W�M�����ɘ�C��xB�*+����}ֿ��D���L���QqHJ�!�<{�ZcV/�I��	��cK1\��n|�r�@��Κ�мr����Ci-�ز32	�<tq�=s�E����/y;e7/kE�vؔ�(,ȌT����-����c�!
l*Eo���k�E[�H�:����EtWe�[n�$|��J� �&�L����AR�ۅa��*�f�Kӄ)F��L�r���}-)���ΰZGZa��3F4����#�4��r���;��D���Ҙ��ۮQ�w��`��Ͱ���n��-�,}�$�.9�p�e��ۮF0��@A	:��	z����2��9/�VK�(w|M����#�2|�-q=,cV�RɫX�v�G�Ê�|<��&��{��L`q��d�QE6�r&=��6�M^�AW�+�B
d���Sb�ͥ�S�'������e<0�N���GT����Ɖ��6��.���;�M&].�q��wܰӽ^J�l��W�N�x&T��/�>�����N����~�a8x+�ηЫY�G��x�v{_ioU��Ӛ� �w�a�g�yp)�ԃy�wѠ��˔"�������Oۣ��Rw��a0}_�M3~f�R�f�9B��Sê�k}��{��'�m諅f�c�x�@M����X�?��%mM�>L�����k=vak���Pȝ��_�0Ʀ�<�;����5f�� 2�	�s'�j
m�] .��c���1�ֶÒ�����Zi��hہj���7���dϱߵI:��L��h�k�_�'ޖ!8Q���q	�E��͂\��Ew^;���t�M�4H�$��􌦩�����8�=��x6�����t4�� c�tfm/�)K�E�a�b�Ϭ.l)�NήV���yu"^��>�P>bN�r:�|B'��+�Ɍ]VNY��j����A-/�y2����I�^�f�{�t�n�V쿾��
�73�V\>nGe�	�΁]�\j
Vj�*���ڇ����#f�+'36���:��vNa5���.����B!=�cH�m��z��Y��{����V�tʷ5�Rq5?��ʤ����v4r&���ً�0�w���k)&_=�e���_h�y�et	{�CZV"���#�DP�d1�X�kLl�ޮsO##a/#y{��{A|�4��
�L�L������>�S��';�7|4�v���ۂ���
w�xN�0᭲���U��$<�iO�ɥ�{u����%鏊���<=���!��l����+U
�W��
mƟ��ZH�q����Hԑ(���"���a n��8l
�hW��'Yb�<{�l�qN��K��]c�-�+��� 4N=�$ї�>p��6������E5�օ�ħ�3�Z}"Ђ�{-<��#�v������f�1��:�aо�<�s���#�Ah��Ԩ��u���|��h�1&mrB��O�����X���p;}m�ėD1nJ����tb>��?2Y��ɷн�� Bx2��֯�I_/�1H��I/L��5[[��NOl�a�$�V�x����]҅ 71l��Fǲ�=�׭�ӗ�h��������Z:+q2��������b�������V�p$8����ɧN�Y�k��ڧ���BvL\��$ި��!R`T#H�tx߶g�L�e�NCG���i{dW�=�Wt$fL;I�P�[�:�(B�����h��C�*��~���Ȑe�� ��f>E�y�-���ur��6��
��YQʧz4Q�M
g=�D��MF�vt�����q��u�� ��Wt%eY��aȷ�)�t�����G���%׺�3��mZc[�÷�o������.H���@;���d��\	.=�F���K �'��JJ*��
³�*�s>�B��(�Q�P���j�c�C�]%.�%�ӝ1���6w}us�Kʗ�_g��F�{��k��kn�J��}����(��ԍ��c�H��������T�]a������2�W�g��^h�wH"E�8�m�=�=Ԛ�M �G4��ʳL��hӆp[���W���l9"��>��Ki�(�	٣sYKz"v��'�w�%"TA�?1i\ݯ��N,��=&t���<0w�b��c����cj�J7��5�kA(P�?D6�>ru��p��F`�B��F���,1�o�Nm�⋯�S����pX;����k>��4���J�n��E�O5�]C��ZQv�7k"��m�m���H���`�[B4V����_��k
&���wy�w�Ҝ7̃d��#H�WCS�
��pt״I�{�P�\��1 G.����I5�?: ��J.,ي�4�A�FWX����7y׀v��>�x�GG=�>RZ���"�6���b	��GI���!�@��S|V�;"�X��s\�`x"e|�Ix�����@^�݈�ֲx�3��O�����!0P�.���V����^�?ݼ��G�=!Й��նh/��*
�m]�~6+�.����E$�jL؂+��6(FoV3@5�e��d-�6�iY��=�E�y�q��|��8P�H]�-q���t�	��`�]�Pp~�R%��\0-;T�ucp�Z�8 h����3O��;�j�ҿj�e�=҂�^O�Θ\�\Ä��>8��z@�2X�؆��bqF�۶�]l,�(��d5�a3��f<� "��� z*+�ن�ﮩy���%��셳I�ż�F���
!#��J��D�wV���v����ƫO�o�Ɠ���k^��4w.#�9f���p�ּ@�����d6��Q�>�
�����К��R��,���Ψ��H���+p�O�B2��	�s)��.V����=�,�0 �k3�fc/����3@�"���s/�n�y��R�[R4�m����}*��N����ZEl�Oq�(i	�拒�&T�	N���߀si٪u�����HE-3>�H�#{�4Y�$l9����>i3�ߗ�]|�{�{ڋ����/���?}��]����f%V��l�z�m7\2ge3���]k �k�`�0W � ��!d��h!�s_B��ӧo:���J雹�Xp���M �K�Fc��"� ϣ��6������O�[ߜQW��
��:��n��O�+u�*��{��SW��������&$ �Ī���7R�)��>fjG��4�<��F�f�kN_��4$s62�Ϫ�_�u9u�:dS�v��'	������|�L������MX��Ժ[ǝPcU���_y�%�Rj�@�b
�p��H�:��R�y'>��T�Wh�C��}<c�D� ۥ�^j7n��(c.��#���trn�@ �Z=;C����\+��Mȶ�ʃ�[���G�|Y�ko�E�P���k�(���)@d��^� Q�E�x�P��1B���
0�4�/�8�V9�S��5��/c��t:�n��2�|j�N�7��o��a롭,��t�x�t���R��MOa	50�5�I��;,6��U�P܋��ŶѩZf�sf��8�U� +����h7�@m��:�kf��\����o�*�Vc@W8v���
�VR0��&�ÿE�Cr;�x/Nca�I� *��h�i��l�T�u�鸟Ǎ�k�x���a����'�v���2��{�C7�.T���M�Wt�])%?�T�*G):E"��X#h&�	��v/����Pɷ�'���q��"v�a@��Ć�E��^��x,Ի\��LA�����=����[Dن���Zc�����R} }����F: *�υM�B��
���3����T�'J���"m� �%��g[׷�y�������x�#7f���,2�1�i9M3�.���l���<�����I�Vp��6�m8��[��d�*��
$'��]-�V�SӨG���"����O�0=$���ߑ��� C l���d@����b<�3e�`?W SP�:	�|Qq��p5�;W���Y�82xTo���q(J�t[�R5����Y�潩G�=�}/����6c������W��+%}��$9��$��լ1�{��oސ�����̜e�CI�4j�j��d���,U�_�61û���y���h��#u�������Ⱥ�&A����W	f`�@-8ۂ�	v"p�p`�F�y�����L^d��g3TI����������fwz��2)���
z�Ǉ�@M��_B�$F4���#�8��O[yK��2�%6^�(���꫘8�=�3=y����cie;Ck����{0�4��K�oe&&=?�
�b�Ds{H�v�$v�G��?I�Ǯu�n� Ia1(�*�ɚ�^����wx��㕛��r!��eKen��&}���4?5�p&	�i�c���pH�ShII�c@g}��ΐ��$\�j7�G��aM����!���+c�V��qc�/j�q�+�G�ѳa6&��5^��ŕ�	/��O7M��D�]�_�'C��h��Fqo�C�ϻ��YA���bL�V,�M���X�Ғս�f��F�d!5-�E�&�vk�ΰ�=CZu�er�Vc�� ���\�(��E9	�(�ѻH�5�^U�A2�w���K=�\"g���Ҋb?���p`%#�Hg����f���;����|'��2pM���_4�F���s�}u1<2��c���X(�o)����F�H���Ԩ��Ɣ��l�� ��t����#�1�ǝp��d8ڗ���X��ΤA=�X6���"[���pv+e0��a�:TBX42�z^f�~F�?���i5&u��
,���]�q�9］]"X��զ	������+3֭����T���Ni��g�=�J�)�R"Y���!~��e�D)0E
�Q��bV���j�Uò�[��X3l�Y?c� Ɋ~0V	
���s�F{Epa�6�BEO����+(����Hd��^7���:n�D����bGQ��ꐓeʗ�+�
�+�1 ^Q��I7:�_�p�D�|b��!�%ɟ)���h�줞e������1"Q�i�[g.k�f���7]���r`�G�5J���V�5�"�Y��#�h�/-�"a�򺃶���Ҩ��E�ߑ�J��A0˾�r� �������nB3�`�l�� 3+x���m�`]�v�^�Ze"_E�Ձ��~%�<����/ңK�ޤ����L�XZw8�����>�� �&%�"]�/)�����<s�\�k��#����g\t�,4`��r�������6��hG���x��Ձ�s[�B�*6��eFV�V��#g�L�F��%{���%�`U����NL=���e�VR׊��fr��_޾�r�1't.�X�Ő��P3���Z�X�z{2�<;Z�ԅ���n�L��P��uN�۹��tS�4��5�|X�b�-sL��8��#z�a�a}��ƴ�)|Fy���0ƯBU�v�#����a"�\�-'1�</��s>?o���)�
�#���<	sׯ��@�ȿ2v�^�|ތ����� I&���C�X:T+�y]���Lm��-�d���ee3%��������$�Z�D���F��m��vx΢�w�L�=�C}�5m<=��n�K�,��d��U���T�K�Sr�����ZHư��e��B[�Z"� �Vͤ�Bxs��]�D��kqQE�e}֚�G��OK'��v����Mu����=��������C�H���moG�ՏW��a�9k[��Qc����B�[pG��υګ�����=�h�&�]��0�E��\h��.˚�\Rn8=[8QѨ�Ӯ >����@�9
��4o�ڮaObP:�s�'�PL;&#����|V[g���I`�HO�]�Y� �Ǎ=���M�V?�ی�32KF�>�|�U���2
>���ΰ�+c"4מ�Q��R�[�c�U�v��%ڿ0��2�U�ܑ,M���=�L��5�'��d�!���J^�>S�1����*�е &��Ҫ�w�/t�Z9�f�V����"�?άUnH�܈�j�@6C��B�a'��֜Y�՗w��l���y�ݳ!RHq��J����'��Vze�O��~
&E��.������͂���2��dī<5:��thjR��.?�{�6l�d�\�bF)f$����ߗ�����哗&�g�:I�AOiKT�sV[)���-��F<���n�����l��n���/�@`����f�����IW��<��M��X�cBR	$��7Il�P�(���0*ko�+^z�j$���axe���4蟅��+D��S8o�W\\yN�X�Ѵ;�m[oF��q�
�x�(�h��1��Z 8�z�,1\|ؖ���4����lsMs��-p�3&[��!�}�]�����w�B�I"6q�ͅ�!��40Y��N�kQC����b;(�"�0�5FIW}��[��}S�u���[�+YU'�O�)1(��L���2���G�����e�V�� PJ�א3U�о-��4+�aCRwe�H<O%̋�g��_�ot"��r�j[��[a���k&����=��g'3��	y��F�`�Z �@�?���L�"��9�P� �[�h����N$ަȋ')U�fĥD��J�g!{wp*��Ms ����t�%Zl,6 +H�п
�\��n�{W�Y/]��J�I	n[�
D'��&r��s�s�E�B";��z&���ւb�gէ��=$"Jwm�>|R`�L�������뷠$͵(�R��1�w%6�u�&w�K����D����vrwN{�G]
J����c�x� >��`�8��p�m1�N)���H�<���a���H6�0�[sq@�0`g�\#V2��|�3��r	�=��St�uÜn����p`3 %��x��W���Iyw	�>U���""�����
e �iE������e\c�m�S��
���O�l1R�\�fF���5����C�*�L6Z�8 �C�D�ת�V�Bt�x�E^��~��9o�v�O��ٔB��o�a���m��p ����Ǻ1��=��z���u�)B
��Z+{�3R�N4�&U��,�E��WU��/=S� 2,��k��5�7YU�k���~b�7�z������	_g7:�$j�9J�mt���n��e͸��\9^���m�� �W���񖗘�+cjN�Y�.��}B�-d�7Е��}����{Ni]�VaW��(�9���ɺ�p�r�c��X��g�Y�8�/���S�*���_��L�;>�o>Q�sw]%�f9�ә����.��[��Ԫk-���FI]<{<� I���e�*AtoW�G�&��i���E�#4�i!�s)�g^�0lh�Y˾��{��?�^3�'y&)���py4IG7���k@D�J�<0��>E��/�X�v����j��!!��ϬL�E���Q0�O���!7���*����3����T���5���<��p[h�/~3�#