��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�a�[W;���(���=1�ѥ��Z'�,D��5�N���������u����-W@��sT��<���l�&h��1
!�s����R�`��ү3:z���bi��͆��zn�}�7�IPb(rh��ń��P7���}5}`f("$#n�[�1�1u��ԪH6&���]��S*��}=��y��	���4�Ma+���pt����cfMn@B�<��j����������Ot0��䳀@8u��h�Zf�	
UC뚮���}��a]�Ak��^-����2�8B��ˉF�H^$���T�2�����AU�4��)��@Y+���ڡ,�g'⫰�!x4�k�&�S���ٛ��ړ)V�լ��y�3�r�q��{�\�@\����R��rk� �@,/��cW�s�i���t?� �KI�{��9]��.B���A�؈[��5��6e۱l�pu�D�õ�ř�� WYI���i�c�PJ��y��-¢=sFV�DOr�R_��&�=�-��4ߢ-�ٺ,��������M��!{j�f
`m�|OG{5�T���ܠb��$מ8̄G��f�P�dFt�d�d`�`V3����\�_1E����/,3#���	n��KY���>��C�)�fKNu��$�#P��(D(o��>�>���t�k䣘q�}8QUu��_��T�_�9�L`��@��V� #��x�G�x�\v�|>;�bIo��,˺�o�ߡ�7���)3��vw�tl�ҖC����J�`���@)-o.���g�&�K���0KzfXp�/�ط:��bYZ��!O�()N$��e��݀"D�q�/�.��gX<�n�j��Fܦߵy��y������0;��ޅs��D66�-�:��&R�p�&cZ���ߔCƭ� ��lX�ט��nŵ�Z�Ou_Q��#8��KS�;F�xꢶͻ�V���duر>��zڨ7�^X(�{����M�!X�fI�� ��X�2e�kK��$��%����g���AR�����(N��
��da�K6�a�t�8/�J�:�]Hvv=#G�V�m$/_�M[|m�Be
����`85Վ��2��(�ɾ�@��p�a���ˇ���=?C65������8
E�+�U��M�$��7��,�0�m���&	��.	�٢�!�}m�E00�]�{���~I�D2�H�҂��jeOT�[������rh`��G8�0�ҳ�g�ز�#"q(@��	8�� �bL�dOp��xup��V77V���[�C�u�����y��S�Z�]�q���C]�?��J�9ƕ������gp%� |�li����u��s��k��')�Q��+i8����f�� �.H2L�un3�*�	o�sX����+RQH������Pp����B)?�l?3O/�iz����o�����	R�N����i��[X�߫A?�ykp閕I
���҇#vJ{�ˌ�1��/�v=�ǃ�~�������:��\�GI��K��J������@;_��L}�g�+��_�<Z OᎪ�c>.̺���ij)���.fg�5�~�%�&�J.e-&���̉��s4�*�aA�m�F��7�\��Ӕ���OK�����G��X����r��ˇE(�Ɩ�3���[����B�W���%��Z�D�,(A��kn�`�$����!V��d�G�X�Z�?;H�M������X��2�m
/c�4�;�{����z�Z��RĶXp��:m�䪌���ӽ�əx�0$M�Z���i}j}����Ȅwr��D�`���r� ��4��0ſ�79)�Y�+�Ɂ����=��}MI� d�X�D���,�1�{� GJ'��H(�u���_q-3�q�x�17V��p����g��q�d��W�U����5ýd�K��L��<a�^?eKJX�s媋ʁAcn燳�����\����2� �Xn=�ؓ$5���YI���s�y#����eG��ae�u-ԒK��ҕ�A�B�S���g���=�=:��PU{֚^�'
T�a]\
�:	?��Y�����S1��L���܀	�:�k]S��Y�f��pEVs� Ί%t3���4�R�E��x��%�~+�<Nt�o%Y@	�Y��r{A+�KK}}�U�|p���w�_2�B�+~����$������a�E����tL[�Q
$)7����� ;��I����6�Ϙ(��i	盞�iTiKQ3�N#���JMw	[����n7�Х�GP#�+���L8p|g}yl�(��)t�Uj-fwq��mo�����{o@��u��ɪ��,�W����޿ LqסXj�V^��`�ۭ�T6/�E(a�'��@!�S<�?������Ü�����Z�ς�90���#t���x�a��]gc����o`+�Յ�w����몪���� ��ᣧ��u�.����-�H}L`�WPȜ�Z��N�����z둅<� ^U�Pw��z�%M�Γ�� �,W�X�]
���WU�a�.����,x���=�����K�lyA�b��ͨx�J���@�m��q�����FI�*�����VA�5+�� 8�pBRds��i�V�Ʃ%W�2�}�'��V���x��C�<�M�b�E�A[R7)�j��7\��ꉛ�a�3�>�_S{�hr�q�����
�Ʉ�>3�'��`�=}N���n8�
�z�欖�3�yG��?������ü
ɣ��Mw�>h�n�'#��z���h���?���y2�~�Jm@H��� ����LO��4{�l��p�N�����W�N^�A�!�O�=*ˌ��j�vdD�<w_�8��7���-���4)�����{N>�X��`u]�	��K���n����
��ye�=k���_�H���{M{�d ]�!
����HT��{��!��3%װ�y�����N+�)?�穩2Nd�P�]_ W���6�*�׈��XB~��0%�\�dqds��Q68�اQ#8p1���I�`1��'��А�ػ󴛋gX�3�Z5��kz�uP?��Cz�
[�c�o������O��'������MO��ɴ�;��9�$�2�yy��@�׼���%Q
 ��3��XIB"M���-�E|�4Q�"*$Ey:�i�O�	�5Ud����K��*T�g����=a�7]��^����IP���+#�p?��;��/^��4 �X���k���C�k�#+�l �����_��xa><Yo�����MD!�Z̸Z��������K;)1&XjЯйpZ�j+�v_��1���r�2���|���c���-�Ldr"Z���.� ��漊1P:��7R7e̢�,�ʇ8��~�L)e�grЅ��I(�}H��C���{�b%5s��DN�u^�ӌ���]�9�<'���r��ǙK�c�r��wO:d�^�iz��?�hqb6��jI�ܾ�/dZ�?')��5�����)t;>�W�.s�N!}�]�s�s�l�t}F�˃]����k~�k���K7�a}��˘���t�����֤*H�Q�G����/˴�j7~Ȧ�f(b���j�s����.��B��@}�mě81p"�عKj|�VSJb�Ȋ�J��Nyq�`b����;"6�ol��8�kd���ip%ie���=j�D���*��T��4��-�؀��	1��9/	[z̫:(`�EI<"��@G�2���(�J��ٕ�/uDK9:Dc,��p&��~Պ�)8V��$)A��#��i�*����E���w�G����ގ>I]����/�w���ˑ�GeMOZjL�x���@�v�>M�iJ����G0�� �`%��;.\ XA�U��qq�B\c�/�O�_����׆XDf�^h'�����+�b 7J	��1�8������[Q�|H�@��Ռ�ǹ��f�zL�+��	!�J�[Tҽl��g�0�w&|�h��P温&|V�a��.�Ԏ@��7��:���`~^w�pb�쌘S�ɳl��$a\M����.���pm�,�!#u3�gδY�w��W�O!�`�X���,���X�7�K�T_P� � O�em>vF��7{t;����9Bw��Cך�� M�a��p�d�cq��&���M�wXSqr@]�%8~T���(l�>k��P���?�EDe�š�8U6In�K߁H��[�=�X�\�����|����UJ�r�{�,����a'k0E��vTr}��U<�Yu���.���o�0R��yގOWcu#۪�+�ulL�(����������J�K��5���;���=i���Y��E2��D42��=J��e����}	�
7^6$+�kMS����|���?�u���K'Rd�.�0���W��N���$�/^��9�<�/���.�4\���N�OU
ӡ���z]��仦�*@7,�E�,�,�L��ޫyn�x�N� : r�ۼ��A��(y��xV�j�8)z�
�z�=�PYn�J���QbV?sQ�f�@�!EKD��aw%I����A���
��ѻ��0�O�eзˤ���C֝g�p�:�R�Ȇ<'w)'�'~�ݱ�پ~\E��&�|�e��$���w��4��X�,
��<�<���q�9g�,	azu�@
)y�4�G�	�B�I�(�8���3Hj��
��s��H�n<�P�П�("+��m)x$3�����(WAN�	�5~��Z������A5<�I��?��e �_D�s��ھpa��0��y�?��>m�5�6l�;>zW�D'G����>@t}yJ���X����5F1:6�*�B�Tf=Qx���T ��$�B� �/S�*U�U���O��j'��!M�R�7�Hs�7���e�1� �-s~��B����&W3�Re��nJ�S{��$�(��Ed�mR������37ǎ�ZQհAY)�βb�)�%$�j~'�7��D�]n� _�2����"#�L[���lQ�����t�r�1�g�i(y��X�iHy���-ӌ�v�[~������>�%��GV��Aѝ�������[�tgK��`�5�q� %g�bւH=�^���Y�ϏQJu��z8Va�Z�&�J���(�{���~Z;P�~�WH����,^�����)�����������ÛW�Xޒa����'#�,])1��`������O��W4���6OMT�TW��fѷ{F�݅��� 	wO	�Ü���Q�,��A��!�2_嗼���_��Ѿ�;Yq\�򇙔���X�]���=p�����O��M�;�Cu/#|+B?)�����ж�ްB����TP�����s���-�x��i��E���B�EnX��M�7Z$E|��i9ՋLYӊ���˒ɅЬ-��"�ĝ4��c���N�X���+_/:����Cl��֙>rN1�w.���aJ ɊvF+�{�Z�eF�|t����TL�o�M�9 �@j�Z�)�YYܕ.�LʅX�����n���c��6���Rd�������}�8NT�n�z7�0���J���΅�z7,��>D��ޢ��W�#�\�� �ܜBv�Ȓ3�PN��G$���?J�F+��P^��[��<L3�8���?%�͚�Y^J���/�l��g߿j��,�V�i��?���q��� �4�!:��N�����	�lg�v�����ÿa�e��E��:P8[�T�6�?wG���!�`T����o����c��}�7��ǚ�5aԽ0
-a�ǹTLbI�3w?��\�z� ��
��P�|ʑ��E}h�#*��F��.I�*#C�Y-�~5Q0�Os�6-<�{t��O�B��ߥK����ps�r�E{v����ֿ/���{炽 ��?��U���d&�\y؋�������+&�:�@;�:���j{i�gk& ����<�(�L��2�5L�Ė{���9��ε�p���U\��w���Z0�(0��֍�~d��vH���:�֯El�l�jQ�;��'?d��0�(���F7Oɞ�U4{��e���l�W.pZ�i��@�p/�
���Gn(��P�P�ys��]�8���$���q�GI,yr�V.��d�@#�'�Kx��^\2����8�..Ѩ#'Z�^���0kr{rй�j�0�o�m���z%.�.sZ s��&�Q�oB!� "0��mY��(��G�e;Kx��\�֬��g���9��A �@[e��{i�n��1��x7�A��9�11|�c�E����3��H��o�Tr9�dr�TDd�O���5Y�:��H&޷g�~{�l7�;���	�`�J�y�+�v(��~�-�G��q��P�ʥq��r3,C/�g4h�V�7�Og0��GGt�u�h#��a-x�.�6�\o�Q)��D|���;��9d2��w��+��ȯJ��s���$�$�������Y�H����I�| �>F�^�9����<��)�ʞi��iLկ����0�����x��>��4e�ۇ_�"�D4�:{rQڱ\������f�x�B�rI�#�������:�l�2�ru�G>+k��eMQ���o~w��B���Թ�R�����[����11���������]ִ�4Oy8-nX̛�ReF�BId�2������x��g~)�`��F��8N&A�PL!h+�8�I '\��F�����|� �P� ������z!@��~d���!LFb�0a���q�� 9T O	w���9x^�n.0��.B�K�Y�E��L4_Irj��^��9�?y��+̔HlC��!U-�It@/,w+�}� �\$�B����H�9U�q�XZ��Q�p5�,A@� t�ߕ�g�F]* ��n>Q	��%Hozq������\?�����X����\e��#�v/'zI�Ti)ْ���&&�_1o,�U��gX�7淰�E1�i�d�G[P���1��p|���;#�ܢMH7W(J���%�4go��W���5����X�z6������d���J4�k�l�ٛ��bZ��:;l+$�?����dD6���q��xk�+҄�U9���G��)��#���>6_�!��퇊�|�Uj{�'��z�Z��n r�c��s��B�H[#�	
�5��#���r���)h���QMy�?�A}�&v;MF����lٍMK��X�=�+��H
�f����j~i�Vo�E������p5����k"H&ԛ���Y����d�|���z6E��R���m��vj{�bw�pOZ���H�bUqY a�[�����������q�U�2�d���W��#X���*Eݮ	m@�ڏ����i�^�+L����1Hr�BA�g<�ji�4ɐ�`Pu1��OR���6\��HFח�DѼ!h1�^��S�@D�i,�{U�)�d���&J��+YhWS���L�R�����(4s���2������-S9k_C���>|L��h�h=��E�� �YOeː̶�
M�?Hu���Ϋbm"۱Rwk�Ae�7��E��6��K���b���lJ<�VK����(�㛌�6�P����r_"��k+S�B��Ӣ�%43M �8�7f'� E�/eHz��ÞB���{x���A~�l��՛��(C��	רd� ��Zp�[����[AGa�%5�3HO�U�6p�C�6@౉^92yQ����3��tfO�y�.�w��I�& (�}�$3�&|�t�^μ���)e�d�s�2䊤�N�
-c�l���nr�L���"��d�*��ź.gv`}�&�B�p�L:?g�jP*BV���x,k���=d]�x]s�I�g��ǘ����Z	J���Я�����>����Q�[dM��ɜ���e�0���|��m�C]�y��0�ZI`��@*��?�?��z�(� Q$洫!x���v Z�����U����s��wcDj%}Zg1�c����o��J_�zQ����j�&c.��eh��8-Z-��W�
�,t�ݘ�������D_L�m����&z{X�����{"nƗ
�u��lz\BKqP����r?Yc�o4�{zg�W��þ�v��Z�,���;%[n؄�u�I&��󀠗�m_���oΘ���Sb-2���ڷ�(�`HԐ���̴A��1�nP�9���B�.k�+\ˌ�O}���a8<����h4JQ)FAxCBث�fѐZ_]=4Z�S_�SPhU2��@u�4,�������-�_�

/YQ�1pѿS3N.g�cfR�ܹ׈��� �AF%$Pm����:���lF���uZ��̫�Yyrg+3v�����>����zF���y܅9B�;t~�S3
��7��.Rn��)�L̙d�z��Ε=��F����û$���7�
�N
��A� ��ZD��]_'V�������^|` U���Y�|��[��Ԡ)Z�G�i2
�[�K6�K;��<'��"��o�kX��SԘ�g Hb�"��A���^p�;#��]¿��JMd��A���r���~�}�&B��S�O&�	gY;~6u�{���a�G��К���QmJ^����L6g7�77< b�9�\ߢ��ḹ
)�Z	���+0�U֓<�d���3���S��۞,-<۞\�TQ�C�?���75��=~C�Rz�h"�K��՜�{��ܹ��)�����(��{U���{r��OG�J/��:�uM�#_	������3jR)8����k�y-?�vT���֘e3=e��H�3��%�8LN����m��gZ��"�4�6�����-�0�gf����2W|Z!ّ2mn��Nd��s��2�/S�1�N�{�a�(�t�TP��j�^������J�-n?�ց��M�o�fnZ�Z��		QkdQ��eNF�N���1� ޯg�&ɺz\EB51]P�I����X�e�8e��:�����37��o�z��'+Ml#�ƒ7�J���N���n�A�ܥ~��}F����ʄ��F�%͎jz߃GY�'9NŁ^���\��ʂV�Z�أ��(x�٧�I{�����1�����g�����V��R�טY���"I*�^g5�/�@3�l�ra[4�e�G�@By'ێJx�W�[ༀ
�W�@rq�R|��4�����c�{������p��@�op�Ύa�����F�[���[�U|�?��K������%��Y�TI[����Q�5·�t[��A��ib�{�sw��C�A�e�j\�h&d�a�o����%GHЧ�#�f��֥QE��b�#0O�<Q8��/(��]�$�3��A��4� �sU=�ɦ��&�=U^�M}7�jB�̭����ε����WC:Y&�w�7MR8�<��>2��c���f�V��A�P���s��D;f�[V�C5���%+Ni�ë�F�3�����V�NG/�15mH�CMĥ]��К�ה7�����1��<*�T�N�0���\�P��Zq�b�����K� �g�8��Ϯ���f��v*�@�ygK���A%;����\ �Ƕ�GCk��c���!E���	�K���`�'U���6݀�p�5/c�6�F���j��^�:��{�c5��Z�w�@�����֯&aRI��@)W�SJ\I㧱D�]����8(&u�?�<z�����N��TRqm��ť�����j�<� �6t
�q�/�~5"F���.��,z���n+�˟Ts�9���
�64���E!ѿ��y��˗>��dGjc��7oc� ��D��a�zq��:�&b��V�`�4�����@�1����2�q��#<��\�տ��!�F�$��z/�ҭ�6�$<�B���c��������(�(�d"1��#�q���Wb3�llEE ޏ�|��j0��ԍ>���AUG�Gn���z�?���Vi!�2>3�?�
OE�&-�Qm�n0<P� ��X9�*�PQ�gGU(`��E-�P�#3;�5�ƴ�\�c�����Iz�ny��\��3^���)H�5��@3v��yi�h�i�������