��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k�EsQ{�M��6��f��g3� �8`pb�-����~/�]2��?�2�)ļqM�F�H��/W�%�� �숉��Y����5��Q�ͨւg�vU�v	���Nc�:�AV��]�dur����$���3c�&����k����'M
 �����sT+�!N��N�2A/@1`ۨPQa"��eG�����儕��"���ے�r �8s0u��}� ��:O���eUb�� �wb(�~Q����Й�ѡ��:D1!����G�z�i�!X�ނ�o��%i �Χ�9��X��SE]�F���V�mjyYw�$���'��q�bI��	�ɚ?΢��A�e�K�6eQ��[/�/�H
���~2�Ө�f���w���XZ}FfU��&�A� s�E��t�VG�"*��
���4�x�=+y\V�x���r���cա������1d �{�5~k�c�P+�a�!�}�W�ܳ@C�F�hy���K��s�{t�Um܂q̺X bjÀQ)� ��m_,g�g�C���s+G1f$��&La!?��O�YL;�����]��m��W h�2�HB��6J��BJ�H�?�8V��W��^����$�Wd�:��]���ނ����Ͽ7}���e���!h�TP�D��][Q@s��fjX*��9�o�ea�ޣ�r��z�*�$��� ���F�"����B��y��m�m��o��,m^�?.�!Ɵh^:��	F^��=�9�8yc4��@�s��)Tэiʤ\�-8=#F��A�5{��G��x��J��5��(tf��hޅ���-%��ᇐ�/Lr�QE>�J�~-Ǿ��/z�������(ݍ9���㗵[������G��8G^��K�a�8w*�	B<@��6�B�OʰoI��i0�Z���q,W��F�0�Q�C7�Yx7�!1��0��=�,O:�K�l��J�l�QM�I��-do�pF����0	����b���oN���r������+������Sf�
l����6�5�jaT����nE!?���.B�n���7�N����V�� �W~��C��Iju�@w�J��ֽ�4]?؛��ЙlJ!����NZf��=�?|�����E�Y���f���4ǓW~��Ep��W�Ӧ��SHh���7������K\eKw{_I>�/�t	_P�N��O? ��I��y������Ì>� ]����V����&TP���!m����ms�`Og1i��X��T�3��7���m����*^r�L'W�o���`�V����ԚTdL�@3�|H�99��d 2���c��<�g�C�A������������?�M�o�x�u]ʦGv�R�,lm��'�'��(c�Y.4u��й8'M�{�"���7X-�"IHj���lN�o~�C����Og��U�D�������D w7vZ�c�,�7cv*�e����D�`Fuu�y���˹�Gq^k�P���3��A�����g� �@p��;�I:gc@7����g����%��rʏ�m2�+��y��,В:=36b���5BL�҅7�S2a�5x!��������	�e7JJ��^�LY��Ρ��*y~�ۈ@�h�=]㭛u9��a��D�sЃ�Q2�PA�t*�`ۂS�H
 �؊L��٘z���Hж����oGf2En��Z���-RZ��y9�[��p*�L�7��$�s�J��\+q��J�7�!�e�~�]{kJ�Tf����*�0%
���g���Ք~�`�Oꘒ�.���r�ם�]��6]���9b�Κc��R��m='�%�`���%=m�K��ˎQC6v��ٌ�A�4�qۢhZ��~8#cvq�cA�V�02�ڦκ�e1]����e��_���L7}�k�x����Ӗ�5�Zm���ʅ�Vj���8��o���W��r�5���r��F�z)(2;�W,��5�Ǫ ��H@�v��Fk�Zn�P�izn{;ѐ�[[�J녃o9�@�?�vw'��"寍��Nf"|KP��� N�b�h�����A�,�,�j�2�Nv�XV	�{�s����i3�$�r�>��d�;�?����A��~�t[���	,�m��(�'�/]J���t��<��Ԩ'��F@�C���*��ʻ�3� P��n{
��ax��`↎�����ᚹ]W#���
2��бC��`�Cx��Ϯ_�_�hY�¤b#��PK]�D읲fD��"��&��˨q!B��L������{��%X��LC#-;l�����G��O�?%QB�_�TQ��d�i?R1�?��b�R3���	!�K��w BQëc�8��~�$�G,�cl�����\r����eL��3QX�����}128���}v>K�m5`�@D�hiG+5�[;vF�V/R�������C/�Ĳ��9����!5�5�0��q�m4%��i�D�9��Q�1>�vP�}�Hi��v��/��ْJ��=G:y�ڹ��;��<�ʺM����KcW)(JS0:�uD�-��ei޽�EDZ��Чؗ�9�x�=5�)��.Ӣ���u���I��S@c��Y{۵j(�F������#0Smf�����O��%R�B�"��/KB +��8��rx��x��-����ޯ^Ag@Bd)Au�C3�n��IRt�HPM�LR�lT�K�ȵ��R�ɻ�DAZ�W %�	G�1Gks.�����杢����ە���3)��S&��S糪D��_��CЇ�c���+�K�3מ�)�&
�^e����&$e��`��%(��T�'@��w	e�GT0;��+���y@Y��r�6n�ݦB$�]?����X	VgX/����N=gM��/q=�h��O���>b�%X��4��3�䳗��l]ъ�o�sά�ǣ��_L�� ��;�n��,�Q��o9����5��t���2�kU���x�/��r��hkJ6��P����Zd����ӡ-]T�u��\\Ҭ$�V���"�,*{I��n�5���;��rE\cIԐ�m͹��㎓�C�d 8��}�Ǎv���OB�i���r@=Lj��3�H�-Y��`�P}[	�q��az^���x˂+c�*k�	�쯜Ǒ�Q�3>�� ,����:T��j	�S�|}�'�I�%��ȧ��,��N�׵ Ӯ�� ��o�����*^,�ч�ǖ�Zq�0ݧ�1F��C�^2�
�{6��E_��A��P�X�$)T����K�����g�|7�O�oc��4�� ����Ci��/��|�x��݂[&+�X(0^
�G�%oJh�V���r��d�/ �P��Z��2���+_��XΒʹ&^�������Ъ\���Q�{<{:����l�b��5�2�������;bvS�x!4�o���β^���6wY�;����;nV�K�`����E���Ov_{?MEz�������P���u�u���Т����*��}Wa9��&jz�ȟU��)DB3j�!~�ň4E������̒~s,���Y~w�t����B���h�G�k�p�����u��a����u:&bTm�k��(���Oe\%u�H�0�Ϫ~�	2v�n|j(����KWS���M�#�m[�����q���XB����s����*5O�Q�IP� �O!�4H���04[��h���O,����=���xC�5�#�� ��0<���dW-�
����;5��o��ʼ?��f�����̴���W�A	*�u����I��K��O�y�M���$��#�_�h��'����'-
e3x��6��Y�ы�$�j$���["����|�|b#6�� ��kY?zn��p�ǄP����mʰ�x���β{;2��UKÁH���*7`rm�tx¦'��d&���{����&c��'�7�\w���2�3�s`�/��xKU�7���X�N��%�/-��4�Uk���Sq�^�E4Ѓ�"�,� ��r�d�@�b�������w�q��(�؏h��Jh,�`��!=��e��7�E�k�/�b)�T�0�o��\A�wJs��g�+{�ViB
��Ż��Ё�p� X�Ž��5�#���֖F_p���O%�(QI>���
��rn�{�,؇��&��H���fy��ol�_�-�bxFQf� -��g����i��G3Q�0��|1�s��4N`a1<��M|WG���t��MF:$��j� ���N7���7S/�����	+��=t��	p�f���(���mE.�3���$����6ڃ̭{H)�۵C����G�}�N"��!X�r.��s��K��f[\���4�>Vi#i�I4�����<����L'֦�u�<V��F�Mt�=�I߫lϥ[]מz�#��*��k�|phIY��W�H��}\c��Ғ2㺎�ރ߁��=�����fwdUhA��̌�@�O,�}����C[�?��
:���2&F�Jl�nG9�,��3�s�1ײ'RC�z0�'�t	/�L����;s��2�M�?�2(w�
#т-m���Z���ov	7=��eEw-�y�J�N%�z���KL�E['X���R�����Gf�+�2F}��%��Ex�sK�C�+���-�i~f�>Z��
��Z��n]es/I����C��7��Ԋv�S�"J.c���^���?|'�V� bb�q!���#�{��Il��/�2�&����x�˯dM�l���q����:U�C�$�kՇ�Ȉ��[z��4�ii��l�j�6�r�;�MI��k�;J�95޻�g��q����&���*�ᗯS0��d�$v���#����iɥ�FKz"]`8����آ�>���'X5�Uj%Y1�v�3���+Ҳ��Ѝ+���Yv׆B�4�K#$G\>,|��?+q���9�D"�`�V"_ә]�<�+�\�,Y�[89�����[,�Q����6yâ/����"��j�/��^��GdX�<|/q��ޛ�"n��vPq��,C~���.�21Ќm-�nʵr1J��fGZͪ��%�m�al��c��
f�w\��Ed8	�����4�SY�u�K��B���e�Z���.)�?�[���g��>����e4}g |�<�2��T^�� <g��q�P��QH��ɕ[��ݭ�a��<�OLOj4W�bB.��v;遴#[��4�F6��=�	��L_��D�SO�+��\=C���%�?2T� ���5����~^�j2��Om q��� �O��������0bI��2�>�j�(*G8�S�����^kO'�"w:��&١d�,w�&����լd)<R�kYS�Z2���G��E��+K�� ������Uf*�����[�}~��%�u�J�|�L�4=R����"���.�����Aę��3�o+��1��&���;��d���F}e�L?#&+���C�����1���f��y�QsW�;�}�ғ���|����W�/Qm*��C=I����̄=��%k6{U��E���I�WMY�4BT������fU��� �y,$��}��ߩ8�u�֠֐pH�����W�2 -�яr�!�"��]˟������cy]��A!����j�&.�:>P
�"����&8��)&��y;c�:�V�'B�C��x��\u�`��yzQf�kn�Ñ�_$Ħ�K�a]�VN�Io�c~^��'�K��G ��3K��.�n��xb�Q��>�RǱXP		��a���QcCGi~����S�\{Lh��\�-;�|T�u�#�Ĩ�p�z��!��@�u,�L����;��fH�����U���^���H hP.�t:�tQ���A����}���g����6���<Z�D ����*����t,���[Ql|�!~l���:���h�&�V"_��J��x�i�ݑ(���K���Zf�ugs��T0�;�5aqJ�_��=���b� �G8�X|�6��}�?����0O//5�Pwxbf�|�)dn�8�1�/xXm*!3A�iNY�a]G^�aA�� ��ȼ�_]mCul�
�݋�/�����/
����@I�#p���	��d&T��N��-zb�}�ԾLo�I�z,�}�Za�I��q�;	�-ͭS��j7�� ��#gm�ky��ϹB�Yx�p#[#*�w��O.����ËcW;Xv�����{"�f�~�[��0CW��b�i�����8��z�1T�}��?�t�ȫ�z^?��.�������h��&�S�j�rs殌����uwN]?4rq�_9�6�7�ۢ+V�f�!a_�?Qh�uK�ҁ���D���ҝ����!�|�zb'�f�e�s:N���&���&)TI F�臅{	Z����`��;xG"g�o~�$������]���u-�?il���X	���d��Pao�n����8K
D������j�n��4�chM��F��-?`'���W/�����g����q��<d�.K�-~ n]��?��`��t��T�xy�Li��i��9%tU�G�Dh��� �c�S�f2�D�o�k�,��hK�hՙ2��{ �Q�vص��F�La�d�P_2��}��X�3 *��޿p;�g
gd�ֈ C�w��3?T�wc3��.��rVS*�p��pg�J�+��C:>\�i�g�n� .}G�6T�;�vT�7�]?����_��.*� �Ԣ�|&25RN�O.���C��|U���83�&���,X���w���C���Y-U�6Ix���@��=�UOu}sp�6*�J;ŉ���uک�3e���/�n<�0M��|�s5a� |�@K�-2�A� ����G@�����������u�Jh���*v���-%���&����q��'��~~�/��jS��i.Y���z�Md�[�_���冴f D��I����Z,EQ������ ��}]Oy��R9JD�����yuQ�=�&7]F��:=AJ��2Nދb!B� ",�>�{�h;ѝ����F�S�-y��wI�&�T5v8��8M}w�8%����AZ�C��/��Ďs|a���N��㟾JfO����`K�I���kls��2��n0�+ML�I�4v�'��5Ҷ��~VV�:x�-^�A·�q��)ٿ��$��8+(�'^�$� ���@z��L�Z�?�V.�[{��S|�I��|�fC��)o��\�p�^�]d&�pI$�v�k�j���|u�̝l��ǇK+��Y���:L� '��aJ<�W���[�7����+�dG�m�
9}bBHZ5y�1�v��-n�SjKV��9}%񔙟$~@`�IAS� ��
k�yMy�s��ƃ����KS��mQ}9���=��)������X��[I�E����V�B��!��hFt�t�>�iddI����L;4�b뻒��V�+-Qqw�I��_�Y.7��ַ��Mq�c:����m�	e�3���!Zk���r���2PF����!��dѭk Ey]/hCݪ=;)bә���X��рڀ_����g�k1e�K)Nf'�=w͔yHa,�s��$�'w��A.Y����+�2#� ?�JH�Xr��2�lnzń�Ck䳌� ^�	��Dʽ@�'��_ ����X-�4y����翐ȵ�u*�Z�����)� J��y����DiB�,~�I���Rsx�^܈ �%�$]�.{������":hd�Y$CG^V�'PtK���i��F{�)zև��]Նٍ�3
��W}]O��Y��~1��k�V��4�T���gm�b��WQ��>�a_{��D�³�v�Z�+���l�9#��r��Ɇ9q�A�s"F�pi+��� )lP��q�Ljv~�	�K�Ig���rIPXG����&��j��gY�� �f`�<䀤�3䁳Cc�֟����`=��	����L�X[(�!N����^����8�1����B�]d��Sx|�]��|��=����&ϕ�<̫��Kq���V�:)1Ry`(�c����`i�ø�%�Q����ya)�9�
G�30�IT2���� �uv�B/D�!a�&/.iZQ�lscoH�g2�Q��v�c��K��,]��?eԈ��Դ�~n�Rh@0b �}�Ks��$͏����r6P�4`7�W�i~je�z�C��r���B@���DZ<u�G��G �� �൏i'>"h'���u�W7Y"ѯ�4ˉ6d�����v+���j��G�͸ҘC4�VL+���L����>���0�w�$v�jo,����1@��S'�Q�
�(��h.ͯ�5Q9e@��y�dB�Rܾy`�(�k5�n��~��,���C;35Q��r����#�_��.J���W�:�)��yf4����p�J�!I��(Ka��ɲK�)��:R��q�r��B�?�SC/7|pa����cY2���B�޽����8 ���G�"Z��$�!'D�O
%������6z=�I�W�C��oz�Իa`UR[��3��M@9�S����9����q�&��tq��S�F�0DXLұ%o���7RKaѻSJ���A"]�f�H;K���(�Q�~���D�0 w�K��Qʼ����Hv�)����R*�<���X��1���l����@A��ɐ�!�iׂi��qe,��!��o��7��I�׺s��Lʵ5�@.*-�6Q�`k�'�͊�