��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI���!qp�6ht����B;dv
�[�܈
�/���t�!HO;���;��.$?�'�-#ܨ��q�X `*Ƈ'�e,��Sg�Bno~����1���V�0HA�=/�c�����)7!/2�����&��������N��Қ	Z�G�i؈�7ХP��^��S�T���4a��I����Zp^�B���,��1�W�؂���K�U��=k{�LcF���)��Idᦿ�_�Jy�����d��iN"����#�,^F"��.P�P�����9���})��ւ}�?�T��;_O�@0�|&���7cgKD��PD��댜2�.��%`:N���n�@�8�ݘ55{�K�l��߆,��`QJ���ɘV��kF�B��+]�4E�`�8�`�-��a$�$$�.~T������n`-*k���_�il�
�J��j�E�@��z5�o�v��W��D\?_��mdk� @�ĸ!�'�M*w���	��w�%+K��*��Ճ����^����1b����l�z�e����J�ڶ)M��U���J[e�#c֟T�`О�H�LP�ָ�q�뤶K�е>�=_ߴ`*}�8ٓE�#y���(l�C9#\p��3��*p��3�<k�I����k����/μGq���z�*ݺrM�m�r޵!L{]*�>���S{dE#/b���Auǐ�j�%Nǿ[ӤSdҟ��x%�J6������^�������ɜ���c-��*+NY�䡍�T��By�
�OcNY�(/
Io��~�d��Pe�$�"殖+����❰��<��]6�������ƢuI1u~��Z�����>X`S%�|B�q��Ni(Ug�^����Af�E}�}d��~
%��e�ɢ4ٟ�"+8�f�LfCz���}�XH���T��6��#sV�0�J���G:�����S�����8�5d�ɒ��P(�\��g�?u:S�nEv��M�O�z\5@H��,���xs1��G� %� ��m�Y��*:ax��a[K�w=�'{�p,y�ֆ��o�"�1A\F�.�]��G�L񙦯T#:M�=˪) �����&�l��f�����|0}�δ���I�qMJ�@_�M#d6�/��SQˎb���$E�(k4����#��[1YT'>�vl[�p��>9*mY{/�[���r�������͑��6�v�ez�
�?���˜w@���OnX�	̟ۆ25�L��k-�3�?o8� ��MX�� X��s<F���]��)h�����Cs�ZP��ΩEP�']�X�:���4�Z�_�g\�5�0���@ڲv��#�lX����z��H#��d�4���&Gl�c�?����v#�6R�Q.Z�ȼ�e+N�FS���`�%�12=P���8A_�qC�U"�(e����/94�gRI�&-���>�����=C�Y�bޮ����p��%]�\�Y�?{�-�R���ܤ�_�x�o1�f�>��	,��k�~����*;�0�e�P5�ᜉ�j����>��� ��������V�D֬����a��;�~�PU��y�n�JZ�W`腅��hA~08S(Y2Q��t�V��:��$�|� �J���9	������B~ f�v�X��Uf3����������!5��a ��̩<�T��>�J��!�o�*��{%����iެBW��k��ɍ��OB�w�?P�U���pSO���c��ܹ)�'�������!�7���'o"%�)������=�3K���K�P��\h��T�'�`C?gu�����a��j���es	oh[�E���������i8��%�mm��
=P�v��zTf�;�Eh�'�岗�>������.Tȱ����v�N���%��Aa	�^5����PD�c����O��j��Z�L��;�wz18�H	. �#�<��~C~3��%+�V�`��(��|��v��B큍��I�e?�W��/�d"Uҥ�F���V�4�xc5�?�_}���}���H��-l�9��S�!
@e��GS��V��"ş�i�?�S6-��H����}��{����ꤊ��*�TM%���n'F�"O4��|�*�M?���&����̐��t?�av�%φ32�QF9� �ҒB��Y��3��y̳���>��>�]�Jcx���WAo����ΐ�h���'�����5��F�@��t�����A�q��ޡ*{3	T�:�DJ�2�,� �P�@E-=����P�=���6�@FT1�ҥ.�����b�@��BN�����#�z,g��`oY�D0b�ןp�����J"�a��V��k�><E�	��SS�广�E�yuce�WhQ�C��U2#��Qi��ɸ�lgyPC����Z���f��_�o:Č +j�M]�ИRfT(�E�*)Qs���Y왭�F��"���y}�