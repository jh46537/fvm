��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c��btdQl�E��*���7��ܽ֋L�a��u-��z7���i���n�̍8�*���[~����P�q���\ʍ��c��j2�"��\���`�.�.3cYO���Tl�H���	�2�n/�e4� �v�-�M��������	���As������gi�-��9����	�{�pٓ.�]�[�m���HV��������|]����,��4���yz�N�E:�N-�a�m���\�'z�uO)�v���J:��~O��u��$����N����v:��T�Q�Ϧ�+�-.P<hL����G�"Ƃ�t_���N��ǈ�r�('f�Y��nF`���,��D����J�T�u�oP\���Ц�^VtglR^!��P|��.}Nk��� �;y�	Ew�-Z_�BE6"ЖS!������25�t0=�SLZRx���u�H?��3�bMR�/��f۷�&55W�ݳ*�rȭ_�Ek�|Q���g�0����4ˤf�NR���1�����r�KO��+㷡�y���D�=I�Y%�fp���^����w���K�0���:�wi�M�f�a�f?�/�M����Pa�&��#��/>�	!����H��V�X�we�t���G�,j��F�m���D�o�l�)P��i��iWOM�g�i�5��R����r��*=t_��l,K�ي��ټUV�}�o��cĒ#e&9�U��P>�������nB��2�Gp�*���\u_��T���)����R���;�¸�߽9�oǯ�:$/�[R�O6����i5���F2Wk���ZZ��RF���YR�8�uѥ�������N�}�R���A;�+������T�S��	�Yt2 v'�M-�Y�T���X��D�#[��g���%y���W ;S�k-�Y��ۻ�F�TB�b^�l�<{�9 �H/�P������Ub�Sʅ�`�mN�t	Q�'���<��΅݊t��77��2�niۚ������X���;�R�z�VH��#��tB뙙����~rD6�,�(�D7Q76yXY��m��tox�Vִ��2oǕ������s����`SڴP�L�G�z��[~}�4.����Ϝ��-��a.aK�`M�9��^��&�j�R.����ఆ�c��6jϣ_�I3c��c�LJ��\0U�������a��)<�������\c4��ߊ/*)}՛�#?І"��b��z�X��o��)�7\����%pA�H��-�=���Bi!f�� 䝫�xU���K�!W2��91L���Yz�Xp���@p�Y$x�@��!��d����vIi!�\fN>�o>��ջ ��-�������g:sY�o �Ϧ;�~�C㷾OeX���Q��"b�k�l��T�@�%C� ���Шl�a}41ָ�jP�\!�59�6����C���)Q
���zVbpbs�Ϳ��h�m��%�d��*�9�l��R�	�c��d��n��u)��̢���"[��ߋN���Joʟ��K��&�s?�ju�Ţ��"r�=k�n˶�k�Fj�\��Q^�T�|�_�#�ϧꉰ���dD��5}��}fIp�T�.�� fH��`��h)ރZUBw�Ό��2��z�ÏMhiPWW����r������/�V2��H��ه�����&0 ��\I���we��ّ�����:�SA���<!iN�f��f��R/�K���d��3O�|`��W,욚�R�ܼ^nJ"����j8M���D�Q��ɀ�8�d>K�b����F��R��_C�z&�pe�ߡJ���b���+�Xf���i�����F#S q�������?��}�
'����8^z���K.8U��tK�Wy� �ݴ>LZk�M�s1O�¥Ǜ��;�]�����w)�OXm�]7���s�V�Mr�XU�>�w^@��n�Qc�Rކ��3�!�{��^	�������I����W��d�3���Q��n�!u��Z�Z�-$��-���4D�`@wb�{�]��y�����<S�O�I�ʾ�(���|��"�d�}{������$X��gÉ�$��������~���:?���з��s���?{NU���bʡ��}��f)����1I��0Q����<�Jt1R���h����/���&ſ ��?�����5�e���G���@@F\�yR�qWg$^�
�Zs}Р%�b�vS"�U+ a�����K;<���o�|����s(x�'��t?dl��K���³�j�]-E���߂9��d����ߜ��1JfR�Ex	K�v��J`6����0�p�/H�	Ű~���PJ�c�`���� ���go�>W�B3��WDw����@� 1�-)�,�9>A/�~�,k~��0ۦ=��(��U����6'."CKq})�ڶ��b���B��/������f������<�|E���gb}���mwB����"�S���|&���Æ�q�ߡ���Lv�����c��8h�Ia:P_��%��Y�!�������R@�� .U��&��'�e��G��M4]�qE[�x�'�O5���	��D2r�O����3J��#��%�{��w��f=F��IaI�K-r@�����e�&`zo{��;��Γ�D�����Q>�Kpm���Od>SY��۫��iS	���X�]�ZY�R�5$�Z��;�?��kϽ1S_�H�shb�/} ��1y����O2$.���(-�Z͕�w�Ol DWq4�
h�ט֯ޛ�-��r��r~y���X��h���*�F槖3Og�,�	n{�U�Ks���AR�n6�k�L��X�9R��Gҽ_�����g�yۯgi�EY2k	}ۏ��ż7�+&�4%�Ӭ���g�.'-=��r��q��5���K�����e��������߶�5�*O��WH�������p�	f�VC�Cr������\"�Uί��g����V��~#���S��|�����!�����6J4O]�Tj�g��6\sΩq9���V���g�\m	Cd��C׍œڛ�gfw�'�FI��i��	k2��<:���y���-L���iґ�2�a��%�7H���`����������B�8y6���*��Rc}�&*!VԦ`�fI�4��jF5�"�=��;�`u���K���w��-c�u������f5���Es6��G<$�0B���їAP� {�nV|{�v)����R\�p���ٞ�1ƙ�G�xم���0��~6��:��R�Z�&���4�W�D�h�\2v�i��u�@���֊-Æ~ �T�,�����k�	~𣍭]��̨�} ��,4�-��=�r��Ϟy�Z��T�{l{���Mx�cGύ���Mŝ_/ -�	�
���3I	=�Cd�J�Իg�C����t$ʚ}���7��@�kx.&�xsm�WK�ː��|I��q)��	���s"Y��Er����:k�b�nG�
�<o�R���7��[�J9I�H���y��.3�]4�-�h2�m��ѿz��kSj�O���QI��pl��Yd�y�	���'	|���i@r��}(q:4��n�bkGuYW)_�4��d^��hLo�k�Lɳ�0�An.B��+���CF{�/_�{��Q�3�,wW��k�R�똯����
�~J#�Ի�l�jy=dZ��X45V��lxo�16F'��*�s���1��mxʛ]9kT�M�"b���/C��hRP>�EQ�IR�t�(ڎfp�)�R��^�#/����Zg��� ��!��Yp|�?)�2���M�7����,SY����^�L��������9�(�}�}	���+M�[P���2��z�1�SZ�.�U���� �`� �rLHE;�d��d��.���:>B�9j`_x�k�������\Pe#�,�QH�\�(8�q� ��I"��J���� �3C�fް L�󛂄�,�?㣾�J3�h1�<@;��|�*od	e��t�c�P̞齾�]�_�C"�0��u�ؿ���̛#�;��c�n�S�6HGgaӑ�:�Mnw������Wj��_�.��f�l�M� �Enw����)cmR��
��Z#W��4X!�'̋2�h^˫變=�����Jژ8�u	U���c�ʈ�	�\��+��T�3 ٹ����#�F�	�LeG7v&ks���1'����k&�Ǭ�����s<}- 1��W̸�� "G��ET֪qv�$ HLA"N���I�0s�5~�?��E����bh\u��9xy� Z#��`���yx�P����Ž�6�tdYŬ�|�F�E?�v�()D�I�ێDs�8xU
Q,�Z��KQ��ty��G	�,h�G�L���%W��Dw����H�Y��V���H�-�%�Rx��mC��N��2���\�ӧI�q���s<��7��(]6�LA�T|���e�K@ϲ����/�}k��L�R��e�揄�B��~��Z0zwp)�:�$��������ߙ���޸�W�%�O\ѥ��2�by0 �_."%�LK&���Kj`��3�Y�v�&D7�iG>��&����_Y������#Gii���Iѓr�Jl�4���U�/Lm��:�����v�"�����۽!��Ye! a��a���ß�"�� �gsV 6�]���^9�x�I����o_T�>��X�P�
��d^�i�lg���C��"�3���j9Cp�Bo�t�w��n�=���k� XDz��d*?�K�K�H�r�/i_��*�0�!R��V0R^T{��	)p�d����Rֶ��7 )��2J�$-����G�-�ޟ?�m)���v�Z�u��s�tzn�%ߨ��_��x*�C&i4`F~Al|=1���*�v������HtH�qK�"WPR�c���YP�s�I��u�R �b�&Նy��hԊՄ:��`ԡ�]�ӰvB����ةH-0�V�q���"���k���i>Ly��������5�>�<s+%��$�ɩב��x�xS��&ZU�}2��,cֶ�˾^��� z�ZD��E�Ռ�s��g��=B����!BTp6��n&(�!��gt��%+����H+)\mu�:����(�k=�S�UZ����4����S�w����2�Q<���'s0�R�G���H��u�@l^w4,