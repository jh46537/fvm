��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O��!N;�?'ǝ�{9�1�\��,�L�B�8��V�R?��[6F+�+�4"p���n�d�#�$؍p�����.�{¯q��ěW�F^��A�S*��|��Ea)��sz�$��O�+�d(�W�n{�|��C�:� O��U荈PjZ�h�'#��}�Z7��-?D����͈#�26���1�o%3}V�9M5@�����s���F��	+�5�������S�/	��;;�~��g��JRyyҩ�M�'������Q����4�1_A�<�����E�s������?�I8��6U�3[����[we'C	�De��m�!L�����;ܜ0��V�~Ջ�r|��˛a�1X�=��
�M<3��(&�<�<���U�p�b��)��+1��+�����=�	�"Eβ�,�������pR�Ry�+f߮2j�۞o

�,>��������wX��2�:D�J ��� ��<���h�S[��h��-(��(�s0�9��5�[t��s�Lm�����S����f�fQ
���3��?�$7I��Vٚq*�T���8�!yxɕ"��f���&���4Y�v����^�re��F��������]���g��D���?��EH���2SM�>ZT�Ӷ����k��ֻ,��9p��3��XoS���,������vtD�S�Z0#���:0��8��Bk��{����7��e�ecQ�6~�|��/��8������y�dgO��4Y���S�`�_�� �8|C����6 �N�.���]�S=W�h��5_ @�WC8��#����d���.'4����'5���@FjL�D6)$2Ctc�,?������	5��f �))�\<~	�*o���>_v�N���ZU��9�`�ly��.l(]2ȴG�
vꑩ�/���E}n����'�ZG��b�U� ���-fɦH����eÁ����&�"w
0R<�{����-.H�b���r��.�6=�{���5�3�?,ۇ��;ր������$�6%j�r�D���|�ֿ�w�3蔀�b�pM�-1�3�vȨ~/��X=�H̹j��.�V��������}_�����4���ѿY6�_0
H����Q�9�֯uFE6>���P��9Ԭo�zD+���s��1��E50=�+�����sG�(��SB���?�a�o�C���q��W��
8.����G���͆lb�٩��2������'/~���~E_�I���p�'k:�M�������ƃ�S�z�S
��ƺ#v��k��؀t�Nf�IO��7ɷv��HuIHt��Dr}���,p2�S?�x8pJ����d�����;d����J*-B���H#���
NNK���s�"<�"�PA �C�OUd	:��p�,?�;���p@99qNb���QO�ηxLꪩ8�`j��T�#9��8#;�3�d���iW�5P�IÈO	L��H��=ؼ�{@i
� ��W���h���������]�Jz���=���M�}敐�0G�ֲ�"Q�t�Sy�gYL@Y��%�����{QKI(�����%�S=����;4��A��0w,g�f�7���:?�S����}�������"d�]��0Ae;�R�~�{{JF����Ӣ�Y��`��z�,�+���Ҡ�~ �cd/�����&��a��"�뙖� ۇs��\��C&AՈ@��Ϻ�Z�y�Y_���{y[L�Z7ceH��*4�\�Pux9���WTw��f"W�H�E�XoX������lO�\�d~]~�v1�����l�#�ź���mJ��(c�f�����ۓ���,G�J���l����f&^;l��փ~�<�a�X�Yrb�~�F�	�.�{V��S���b���B��?����k(ok��(72�"�FhhuKf���Խ�Y��i9�$����7�9Y����ߎ:��k�(\y5�����*e ����1��w��wz�	x���ל,�#��&�Ǫn�+˥���>s�(P��p"����8dǟH�|9���6�XC4k��W����y�b�s��Î(Y�r�ͧpJ��"ц�.�Z!���U3L��d�O��o� ,
�'��T�1�,�!�a���?�
=ғeՕx���x4�c֫܄�I���%Ta��Wz.��64��\����yy1��U�4al0F��է�4���c?I�w�P9����	�L��������c{���P�Ƿ���@�%��C\�� ��ōt�H/�4H�����6��i1=G��0��KVl�"�q��@/ה��^��_�O��"�f/�l���_�����~���j��i�����ς��ݱG�� l��fG�km����,�Г�HO���$�S<�ZE�&�ny3��_RF����0��`�:.��ʕ;���B�F�i�өvGH����z��:�
�1��
n�]�Y�HӍ/A �� PR��y��s%WI��^�g˹1�E�yhԖ�SKf���!�K+T=d�-.�"1���5�&�ͯ��@���!�C:�C��)��2��ȿ9����fD����ɩQ�u�敂Z�o0-U*O�j͔�����L^'U�b��x�o��I8MM���� �|O"��m�v{M�k�λ1E�X���S/��V�]��ǋk�|����^��m
7/���'�|�_�k�)O��a�i��H����Ċ�#�2/q���o��a���S�ֈ�w󻗑���I�bOJ�z�U`L��Fĝ��d;�0���'�	��+�f�Ջw�-�z���&��}
�2���5�k0o9��d���&���Y�>�?�&���]��(���f�����b���NM�\t�\x���O�*�ALmx�?_������u��}SP����~m��?Z�ă�A�$|�%��6ǝ��q;�wr.D�in>�.�ِ��=�D1�