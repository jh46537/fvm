��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���Ox���0��?T�}�D�yBl98�锛�l	`�ġ	d}�:��PƸ����~��R��o�K�jV�,R����vy���3����O���Z�����g�̼A��v�{�7
��5�¾����B�C����������r}�:ش)qqa���·����BW�4����"V�CL�zhXo�e��6kT]xl(���%lT'�W���'�N�V#�L�`�`�Xy�6$���:��9I��ì=P��uS�I�w��������F��<��s��y�i�u�����ml�G")�O�4����}�,r��𯴢}�鑪 _@�y�Tkt}��8!�JŜ�>9��C �gl���-����{���Z�*� 9�[�B���c�M�͠�+�G�Yy"TGz_'l��2/;��	^F�/	b2�ܕ�Z���./k7iǶ�>��R nS�}O�i|�y���I�J��ohD/g���\��'o�_Xn�K���{~�	�������B1�-K�?�m��w>���:b�Ri�yČ��N�������ל�J�)�h��ͣT|!�C�4�xl�C�Y�Z��,OϱJ��R���e)=9�e��R���p8��7�*}:�M=Z�9��(T���3rBt�{Ndpz�N�whaR/��_p�V���G-�/�M�1�����W��ԫAv��H�N��_��0�磊���~����C�ޜu�s7IX݀1������ ?@%F8~}uF"~^{N���h:A�P>|h��X]�{��2�2����>v���H�.WPr�CWv����p��#�|�/f4��Ҙ揍�8�O(h�8��'>^�p�H*��Dثz�Dc��V~L�+zTU�w���LU�?��+ ���ud�A�t,�!�A��B���ung���a��laF����	��h�&f�ษ5�爔��5�,��|�Q!�6��,�Y�$��?T^j�|���FU��L���\?�9�8��Wr��� 쾵-�*J�b�P�pcMd��p,�E�[�c�
�'�r��7�O�-D���T_;��1��_K��|R!(GŜY�u��%ڴ��?2����{`.}��a!�PsL�Q���.�z�G*�O�;�r����s��[j�
�6�`��tv<b�3�Ha��p\R�}�
���j� �������a���]�ʔ�%���U�p�=�)@e�pz����Kv�U�qG�O1(ʑ4W�vץ~y���;��������L|�P�̫z&���)KϏ�.?y����\|�D(�I�a7��S�W�<���Ԫ_���g��D�446�cTQW�$������엝�̤�.'?����K��\ʃlX8�����*?[T�� �ܕO�T74U��g�7�i�sI���kǂə�|!�@��9z��*�l4DI����.��0!�!�����fc���cߵdܹmlX��z6]���J�[vBmb�V����G��,_.�Ɉ�̜�'�ƊwD[LHM7h�lӖ�|T�X_�קxt�����B��n���:�	kdu����S@�M������	� C??����S��ZN�Y���,|p�Cw�G0k	�U��4�Zv-1i����Wv�$|�#߄�?��۰��S�8�B�9;T�4��&��B_'�}V˯/�0�Am�4�d�<���i���X�*��'.�< A6����sBo�8Yg���Zػ�jǼ�=�G]������W� �ƿfѕ��Mr��io��D�����(�����g?"?y���M���jI�I�+E�m!Dc&94����د�r)]�3k�c�ǒ�nh��\�7��	�Y�Ɖ"W��ys���ߥdf��gN%�8�Dxw{�����*K7�L���k�_7������o5��u���Iq��i�����_7�?xku+)���Nd�o��?<HɕYf������ͼ�\��e���;���q��Y5��#�1�Rt��r�#%?1�V�|>@?�HEф��?O��I�|�����4�cQU"��8�������Υs�9��u����z�>��W�Rv�[�0�o. _�Ө��[�2�#�=�^
L3�@T�]EPͰW���4��x�FK���Y������Q�wp/����y��<�'�Dkْ�f�K4�����fպ���TJ��֋�3t���:)�L;�{��R}�hZ#"�����Z܍;��`�7;��CH����&`���7E�iwn뿩Y����R���q��!Kʑ]�s����`y�h�Q��ew!��\�'���&�_	��DX\��hEB>���3[}ۧ�iM������'꠮5��>w���� �N�X)F6>a4�����}7����5�0��g33mыUY�Q��%��R���I�b� ﯩV�wV؅�Րt�8�g>�=l�]�6}{{�ְg���f&���"i�1��H-���H���`N|�H/�������ak�6w��YH�f�ή��M<��.�i
͛{�T�X��nEV�����Fj!�q�Ry����'m������%�ϸ�*�i�k��_Vόwrn�� ���;F���q�P���DdM���OD>��2�f��88oy��GR}Dہ���9�NA�t����������|�^�v��B"3���?G୾��1ԧ$1�����i�<\�q��JYޡ�-?�Hbnh݀Q>n	��P�8�|KƠ���df���L�]��7�-핂x�+{0�D�-��TA3��gp�Sӫ��	籬����y�=�8�
_l�}1:n��2J����5,��Wl*V�C��e�G>�}f��Gm�����oE}�؛�M`e'�ҙs��;��2��[��)w#G�����=,��S]��!4�Dm7��it�w6��Еp���4U������"�6��F�ʻ�x��{b�T��.��bj֡�R��W�9�z�Yy@#�����	k����� #��?���1��0�'�e�?io<�U�.Bߍ
�a�ß�CB2� (_Z)��l9X]=�����Uru����D3�ց�V���8�"}m,��ɟ���Ȫ�b�̠��}����}���F�2t3�#��v���Z��]�(���F,��1$ #AO���	8,��Q��D��Wq�?�a�	���;�h������x��1���m7H�x�#i�C�nW��������v�ޢ�;�����&;X䧛+Gb`��z��U�3��戮��КE��"�������}�@��= ����.�;���;%��}܅A1x�(�:���-m�g��
>c��ٔu#��
�� ����5vfBn��Br����_��<m�#�(�l����_��
%�{+o^ٚ�1�u��E�����nE��t��F�h�]��
�t�0*�z4?��Ld2��koW�2:.����6�: �$��yF}����H�Z�w`6/�\^�Q�Y��%�qx�h:�^I�t.�D�Q��*�U����CV�S�L\:�c��C�:�,�y!��-Z�{�7�8�?,c�^�c���|�]���:�D�7b�h�T����K�z��
�0z��c��a`��i���2x��x�����>�Vuqb�����!��<���z�^������D�D�_��rJ#܈,A�/�����V[k�H��ݍ�Bj1�Dʶ�;j�cK�{�8-�`�kE+
�N��Ȕ�T}��EmA3�j���Y%^���q�x�����/1�t	�sJ�߁�>� �������R���є?e���T��O�\=�Q�ٷFd�cZS��
��!��Le +�y�3��A:ϠPF]q��$}މئ\�!���F�il�߽v�d]ُm�O�{֊UM�������~w͐Ĩ�4����ƞ'�#v#܉;�>֭�JL��A.�9�}�/Z��
��#��7��5����%�Ϧ� ��R��q�]�M����+����c<%暐���8�М��
��w�!�q��'Q�wVn�'��$4i��OgZ~��iM�=Ƹ���a�O:iۛ��f��]��縼���/v�GI��K����_�5{��=�֤V�8N��Tǭܐ�E���3]����O��u��J��e)����K{ws[�h��.�K��c"����ǪBdR��V��@����}n�}	�{Ͷ����pQ,B����+x8�o�b>L<����x���焖8w<b�~(�_��J���@it���a(ָ&����83# ���"�\.`?��ϗl��/�_���M��ו������|�mԾ�n'�b~: uEsq�bt�j!��J�E���4I�ڢ�U6�f������&\]�<k̷�A����H<&��jY�gYsu���q�ޅ�e�>��FDAɶ���8�Vj�ǆ�����7�c1���\.A�G8�B\��0W^ʟ�5�<)'�0y�Ҍ/�9is{qF�ێ|�
]W~	�p�:C�aR <k�4�Əb��4�8�m����e��WS3�TZq��{V�6�4�L�૿n-�?�6m]���rEzW_�Bre��¤(�b�"ZZ������@�"��/�/����ڞ.w�s-52���0��
��K�;aMB�}��������oN~34s����)0�nQ)��$�i\9E�6֙T�g�,��L�OQ#rE�l��.� �Z}��\���*�_��E���k_�La*��1��]�e��R��?/��P�NU����'ޏ�Q���>%6��q�.'���'�*(��@1���"b���j.��`�!�h���!M�}&��`b¨ui�6VR��R�҅����.=L�4�O
E�,����	�����L����Հ�����v�� ���wt"�zA��[|���D�F��JbiFY����0�^���S�o�¥�Żqդi1���WO#'%Q/mG��Hx�M?O_�N��A�������.I�_�/���~��ɚ��M}�D�E����.lG�jS�#7�K�ٽO�����V�Ϡ2F�f��/��Cr[�q	w��L�Q|L.���"��9&�)1��� �~&��AnNh۳���ɻ���`A��k���'�89
�{����	��KN�٣���v.��Z��3����t�k�$�\��Q�:�I�+��s�sb_�/�K�����N��1)��� W ��տ!M�Vυ$��:$u�ߌ�)�4!�/�O	%;.F{A��+T���s��L*Gf�7"�1�p�S�/���T�6w���[_�#|8��m��	�+��0�E= F+D�5ʬ�����~ f=�8`l�/S��Ai8�p�d\ro�����9Qa��?���tb�߲�3n�.�8�-c��<�ݓ�b�GhE	2a�u����]��?�MsT��Q���5�ǀ��tCqE���Iz_�.5�Bx����bxG�2��;5n�	v���]����W��S��u+�&#
{&Rm�۝wW2�5�����):.��AO������P�����el���aE
�z@A�0�P�����!(f�ML{}C�V���m��(bںc3F�w�30hJA����'��ǵw��A��v�\K�z)�k��/w�>R���)zi�$��%�X&3��}��)�>�O�h���V�U��0N�dn��VdIA�D����L��ES�B��BNq��m��io��/��`0[~.����#�a�����`�0;�� f�V�:Ry��3��š���wA�:I����~�	��B[W(ٶ~eq |�<7��4[JZ\E��s
A�7ɐȋ;Np�ӛ3��'hu�	�	
��.����*¡;�v��y���q�I��f���8�M�-Z�f)��Ӟ:ک�=f�Oo����%Z���Ц��X�Dt Ui�h5���Y2m��y�ph�����v2����4$�|}o>����H��Q�u����|!,�n�w{�ݩ��� w�&�
�a����L�h��˩�,�B_��d8s.{�_���3Ԙb�P�/�m{ߠ����*k�`xB���[�'�5I'��#��QE��pPZ�B��t�f���Ei�d��aaV�M`W��~�H !j�ti'�^��������k<F@�����sos��jў��u��{���Y �=�u5���Kj��b�!U@������;�Vw��M! ��mȼ�lN���*��%[j���6� 5�t5���j@fùJ���� ��r��^�Q�]l������xfګ"��۲JYg3G��76L�d/�g�BrG��V�C����&	�>�O��̉���|H��c����k�;��ۇ&&K5�@���_�>�F��G�_�d�Ъ%ji귢���U������l6�O\�Da��5����1If4
�j�+)>l��oi�"�=h�"�������?_L&�U��hZU���7���F�}�Y��_r4୥a%�]r�Fk�y�|_��]og�m�H?fh7���e(,n5&�����N A�Q$�bTڙR�*b8]po:��.�>Ʉ��߂qٛ����:8�_����+�NMH��i@�)�y��R���<���3-S�7#j-S�{%ԅ�,G׿Qom!Wf��=KkSI�%t<��~:�׃:�݄��� ��C<��ݜA0�/+��C۬�
i�Ń4��Ȉr�5p���]�s5�$�j]�����]�x� ��y�׻�K;�&��Qw���3}{��0�\%�Pk�vnz�KG�R���G���W�kM�y�`��������eH�ݚ�� �a���lj�%m
�\<1��%y�E}�+G��Ms�x���,bʁ)��L���M���0�fs�\`������ڠ�̑��N�VP��ΙI�8��9�d�F�~��`�Sƾ�6�� �����p���.⍰ȲԐ�_=�k�L4�aN�1�]`!/T-��EJ�O#H?B��Q"r�Y���L�K�(}������ձ����y]�^%�R$"3GL.R;���ۙ�q
�����_�Ѵ��m]��P��E>|��>#8:������j�BȦԵWlK���]\���6|�TZ?#����a͑Y�����2Iy1���`1k智Р���w$�����r��<䃙��=M��}'����ضb����g�OEV�v:����z�VxGh��	ȺRp��nh���Ԅ��*����tA ��8YyK�3/�Ǜ�����;����$V� ?L�XѤ=
3��PߟR�w
�8��'{ sK2�d����Dx?��C�2�LQ�/R�����%��0/5�Z��'��]t�������3h�� �Xِ	�ۜ��%\��]/��yG���	����Q��g������Xl��a%�Ҩ˯�P%13]���5�p�jY���qضt��ĵ����m��^��!nȒ��@g֪�|	ވ	�+�o�o����)����D.���� �(u�����r ��#���/#��'�*�sL'ι�-�t�1פR��gO�ނ�=�������BX�B����^(M'G������)	M�T���22��*��͉p�l�HE��`�c�:�Z��Ѥ����y��H\����&TLS^<qT�rg�������>a�O����'��|�X��%yy_���¦��8+��Uyw� 5*�/6N���$/j��֣@��vd"�kg�F�o��k�� ���|H�����m��V��bi��
��XB@�y!� ��C����VO��U�Z���z�Tf�w%K���=v�����X���\ZO�ߨ�vJ�eN�T<�?��c�O�8¼=�-�|)r��8��7]Rk5���1�ON ��oS�n
%�V\��Y����(���� W32�}�HNE��7��	�="�c�k��ʄ�p�3�{�}P0�r�	���
��e�a�#�ܑ��ᢜ�t�Fv*��ʦl�*,s��~݌ݿ�ԁ~4R��`9wH�=��n���E�O������k�I�5���i���cG|���b&}J��a�}�{�9s�~%�E$��7@(�\�7��u���B�k�>�����6LWΰ-�o��d(��"�z��ـ�]�'��������J���&�2V��S�q�٩H��5��ph&�}s���곌Ick�fU�z�޽�-��Fu6� �@���b}ʴÈ�ʪ������&��v�[��E0����Z�����H��XK�/q�tVW:Qe�@�h�Mnb�����)�ޜy��G2P��&/~�@ؒ��~�6Ɣ� ��oD���;��.�������!�b��~I12��>���k�S�A)܆����1@5��K��-4&M����a�S�MW�8<��̧h�3#̶J�	�N���(��]��4�3Y|�<s�@zP�zS�#�0:�a�x�gM6�d�E<,w��.[6@�K���iȌ��>�-)mpÃ�b������U��IZ��P��塧8(�f�,�L;B"�����^p<�zn=�f��z�Vt�� `�p�G�6�U�"������������E�F�E���d�i3p���\�Tr]X���]��A��1�'1��-O����b�১�Y�ף�.tQ6"j���K�;�H	<*E�j�Ø�����24�lī�PYސO��R��3q�Wy�Υ����q�:ȽX�bP�٩/��%0���vaI	�=�#Нpx ���}�2��x�J�72�5���%���V�b^��=�~,�a^��S��W�X��H80��UX����>��&��7[Z;N'N����4��^��<���	m��}��w	(w^~B��i�\N"���T�h��¨fx�8-�ˌ���Qk�pp�aE�)������C���p�����w�y�7�~3�Qu�MS�>�[	z��d��"F��t�-0�8'����%��?��Sf���$ ��^/y��`Kg��SYO�Zѐ��5z����V��-XO�HnQ�r��Fo�$y�-��lr����_Ŕ��3�(�v�4�	�~[}�ȣz�'R��Ķ&�R�_w��^߾���J2r&��L%�Sz���|��l[����GN4J��ڇ���*�
K�^
�DU��lXj�����m�d�w��!��uz!��X��e��ȗⱂ��d�C�;7*�"X�"�N�Ï�Nm�� ~�ru3������8����f���5��c���|��M��ؓ��;�P�T�S5�4�y�cW!��>�7�~����q*}�����)��X�kb��\�Ц��9.z��,�]���s��G��L�8{�\ڂ�U�6�C��mO��\ɜ1�i=����/�"�cv��D����z�h�a�.�����sI�6��֖�x���˛�ڋ��QIl�%x<���3n�r�3AE8Ksk�,��[=�W@P���[��'�&u��'�M����+^8A����)$��j�j>8wF�W�6��L0��C`Nj�Ϸt��"�j�%[�(=T%����wds8�}QSJ.I��]C��%�2��˗h�X]�9����M+��J�hr���F͡6�谾�5Z9��Rb:Ir�?R��'+q�\������rʐ�·J��� ,��ʊ>`ӳX)�'�\� �n��F�%�����#;�a����	6��L����!-�07��1��Y�>��Ru��NzOf
�m)�dW~b�	ǎ�1l${��!Pp��VbS���+ۯ�F����?�'�eƪ���u���r�0��
��Z��͝��y�pe�]�Q��ʔ���A���>B��s�d�3����P�&|-7����O�މ�=s���6߭���	jM�6d�C��X�z��c`��ļ1����r��f�Q�l�Sr!\�x]����L�B%�;X3al�|m��D}�ƥ{Tø�nh�P?!���S�K3��e>��u��?rP�2��]o`$�[a����s��-�rtB��u�촨\���ʺQt�i�Y1 �I��D4e�������|V��#�GI_UnK�!}��(M�.68�1�����˟Lmg�y��Ft	A�Y�d��aG�q�6ȧ�7�$��Sώ2�.L=!d��c̀0�����b֫8/�Ly-o5����mA�s]_��8R2�U�,���a� �0.����6���3z�Hu�%�믆ޥ�d���RW@����n��FI��NA�wL�a����Z$�TB�JѢ�P�q j]3��5�K�1v�<�-����d�	
 �y9Eb�6�x k��MN���c%�\'a�]Lc�!���.��a��-�E�y���l�ўG�t�C����Q6'u_�:�j���W�{Ə*+��Ϩ�Bo4g��Q~�4��&;^1G!b[��itJ��*����w��i�6���36��<[U���gG��32��_���n��������$nݼ(�F�e�1�$.�q�GLƸ�����O;��Q\
r�ǈ���R��,��l"����Q0��U�J�a���&�Z_@�.�]=��&�=�:
�������q�]vl��F�Y�5����3j�f��??�/g�PH���\���i��lˮ�����!<�&�u�KgX����������\۴r�]R�Ʊ���O�&q����"�Њ̘�R`ȁF�[yTn.O�K��Xϫkrޛ�?�Q�T
+B���u�-�&J�[W�u��G��	ø��Н�v�����A�$��������|
�>w��ԥw�� [Z�O�LF��t������z����ҫèD�3�Ń�(�3�^�x��w�2  ��F���O+�	�Wb�H�R�Z���<G� Jw�AW�����炐�S-�b��a�&�n���O��{�&��:	}��9Gk �:���5�����kI���O��D�6n��tw�{��;�H��<�Dai1�OZ"��Ԯ�"�a��n���Ѣe'�o|��e�B0�X�>�e������P��_VM� �p�-��I�<_�1�5T>�қ��0���3����O��{^	�& �R�F����$^#��-%�Z��
��]9�N�ŎOv`G�����ϴcC2��x�g�k7��3�{-it�H�:�0e(�y��?!�E��%�?��G:���.�4�J��g�$Đ��LJe��8M��a]��nO�1��#D���Ea+�ɂ��r}����>��}(�67IEڠu����p�["�w�pB����҃K&��(w�}��jk S�4#d��S���@S�ɺ؎� ���.�d��͒�v:U����lW��s^o�kX]=�RB&����6����%����^\��<A�+)��y�{�y��2�;R6�wBR�r,y��n�p�wT�C5�߮��L�S(�Ǜ�B�'1ܽ���nǠ,�������n	�R{nކ�X����;����1��y\�S�`��>R�VPQV��r*��1GUT������uԥ�7Ȫ(���.��5z�Nn]=}F�o�2���P]{�ü�gBu��hjEY�S�89����<�����ihc��%ї��hETq�.��@�H.��FZ���d�G��O�z~a9�A��O�>���_���.��l��a�0:���[\��u��q�>��'���*���9L�x���h+��k�Ȯ���Bz旈��pP�ahݥq�-K�^�#TY<A�)�@�-hu�@Y�RZ�뉧c��j��2��S畝E��ϱ�O��KUo���6�Î�YA�P>��t�_�4�i��"	뼗K�0!E,Ʀ��CTO�@��U����j���]��x�0i�S�4z�Z��kl:�nu%�]L֠�F~��H����T��^�%���@>�xuk�����	�~�=ǘ�D���j������h����x$�����ʹ�-"q51�%n��)��2�'���^� ?ڰK�=� 1!����Br�V�
b)�����8��C��d#��	������-�՛���Ê�/#ۃ�զ��"6i@��؛�YV4�=&�@�VQ��������[��7�����n��Sbo�m {��`_]��^T�	�H*�����#(3�B,��ym	��	�Qx&jz
�.0x5����ITmt�^o`�' 7�Pz�k�:���C��j�H�)M��{�P�(2�I��DvOs�9�&̣���pHD������:�]P��rC��TB#���������k��U��xJ��[IX*!gOӸ�/	 ���dJ���f�{N �$a��}3tr�Թ�e~}���e��=�p*�_"ik��4�{���W������`��5�H�h~,�2@v]V ���X�U��e��i�?��A�_���M^��~� �6DaE2�����.Ǉ�wb��2
\k�ר�=�P�A�Ե�}������J2ΰ�ȯ5K��ʭ\�R��v��m@��:�׽|HE���`���>\���o�F�o���
�nާ��G[�Zw� _~����a�I�|x\&^���%��fP2�y�b�[ƍ����8(��R�"5f��S$ڎ/���M��Ks��Rn�{+��eg<�|���΍���|V�w���=�?����%.L�K<��B�B_�a����J�l���j~���I[a�7R	�@]����5�G�����ϧV�i7΄��� �0ɠ\�1��uHw��d��wV��~�ȧ��l���r�^K�s�ǃh��Gq�WIf֕�]�w>�x�!��O+)�IP�� �TPH��+��=�ժ�#��NT�ˉk;ű�l�S���N�W���U���<D�R��
lEP���8��N��3�����>u*���aQp��@o�idv�$���,.�ԣ��8Lnߑt���"m�Z��qU��K-_�R��5�,��x��&Y<��Te��E��3���Fm%��xY~��G���Ĩ[�I�\!�T B�O�p�}wT�1��9��;G�A�g;k��#���~I�8c����P�����Ā4��%!�u�d�2j�"b�Hv�rh]�0f����I�)g��Y5�POVni�*.��=�7����7���V򱢪5
$���ԕ,WK(��~'t��ᑯ��(#_�����C�kI��>�������� *Ut/p��pvi�H~v�5��D5��9���gS2�q�]X�P���A�\�[A���]>�9�����%M,��+�������5I3�����Cl�(|`�~�e3��R$�	��>y����׍U���,l��ֽ  t�l˨j��ٓht��1JMj>��$bIl������-l�6�����W��l!�#ϐ�$����ξ��D�
p��:W��������sq���M�L
6���} x�}Ǭ7�IB���x ��i^�����j_C���-�U�/ǌr�U�%W[��:>E!t7�)�@���(�֎��}����]p4Z�*.`:�o<O��4���'	�'Ƒ�����$�r/�Wc=l�s��Pq[8ȱ3�G`Z:��
I�Θ����Q��Bd�{���f3?�f�o)���m�	�S��LeF:Ԥ��+�N�ݞ`���~���w;����t���F� ��դ�)d���F��1�pG����p��������^�+8���_�jц�_GwG�-zhk:
h��R�+�@�a	��Y��81"W� ��aoP��/h�=O��=���6,*X��֥N�k�vƪJ��v
 23#�3�*�d�]�d% "�����S���L�5:a�k��B&#���"LHQn���b[L�s�F����Wы�oB&�����#��oj9Z�M��W���Q9z2�h2����j�kD}~����1p�Tw�D�˕`�kJUqk�|}Z�u�1���}fL"�?L�j��bIY36�����-p/�Q:�T%w�9Y�ow�kY/��vW����9�j!���K��%S��W�*W�K:1B�n����s�Mis�Ԡ��jKL*����gwΠ��Z��TV��e���ɻ'��:���>��}"���(�1�K`_!����{I���u�T��ҤC����Ԥ�%,a�=ˑ��迭t�꺓yZ<�UOMĪ7�s~�f��t�����r�|p�@.aF� áY�OSt�i��e�:�u3��W��a�F�A#�R�.���̗�	`�+Lc�V�G����#u��
��k��}X�:0�:)��o0[� ���ʥ��L��Y�b �ٌcW��eu��vE�y	\~8A���2pp2F.�R~a��G�j����Ⱥ�]c��ON�Ω�@����y������ި�>{<[�^q]�j=۪r��Y��l^)(�qGSk`�k��H��#�v:4�v��1R[]�)�۰�����&M(U��Y��:��|0L]RvW���q��ƉsՏ9{a�ye�~��8co��;	<�ś��>+�䝒14$?��6ĭ��"�W-.ŗ�5;7��' ���2%��u/K�.L@�I@
�=Z�r@_Cɼ͂.�G�w�j4a"Tw+���L�h4�]�]�=4�-� ��èH�:��\��5
,pL��T�c�$\� ����k����i��|,lM����	�ɸ�]�2��$Cgl2��OA���'��t��3{���69�G�[�|�����[8C���G:	����g���<.R��nD_t� d�麉>`"t4_6F�6���R�t~�A��������"��<w�q�^ۮVU�&�i��l�d���#���Jp��M5��Y�e	�`����-�R,X�d)�3�M��?�z�!2�~���k;4�����O=�� 2(�A�>��w�ť�',���q�Ą?@]sF	�-��	"�6��s3տ{t��d��0oB�����?��y4.���_�q��~�z��^���s����NM�R�]�J��:�������ĸcS�I(��gpq)����x��O���v=N�����
(���5@���M(�.r��		�p��i`�<��2�Z@ Jޕs9͎�i�����X���C�T�`#�d�,�M�'��K#Y���}#\=8��2}���H���WAJ�\5�R%�~�UHφ2s����Jn����}FQd8y���TU��n�ڟ�a���1d>aߏ'� ���8����`N«�ӽ�L�\;�%Q����9|Y��� ��ƕU�kE�E	��P5��ө���x��úA4B��Vl�ޘ�0�(�	�yi�v�H�v Nz	�#aFYۿ>r���6}T��z��?Vd?yĎ}k�&��gȐ���W�*���)�#��+�����"X�I^I�����_��ˌ���"�+:�� 0v�
��ww������5�U�f�>��,(}4�� Q��7��lY@�������.��ɚn��js� V��s���b�i��<�1 �`\���P�CܰH�|4hYy<��(!���ID�V#�6��p��<2�ie���(.��x��u�,)�k��5A�1YA��6]�]�`��0ό;{n-5��(�s�m�3i���5T�*İ݊� ������%{�qj,����GH\,�s��8dS�q>�~N�[�u��)x}�����^}���Yx���Z��wm��O�fϻy�?9qc��4�Rk���A>��f�D����!���~���yiǉ��Q:��K�8�uյ��bY��IQ���ۋ ���j�U�K�s �>u�m�#��X�(�K��P��_)�9*dF�S���j)�(1�W����o6�P0�� �R�Uo�:�(�I���ֲ?���
ŏ+/�r���?�n�ad�/���*�s涄�q��r�OB�g6|+�G����G���8TW�2�p�Y��A�{tt����o��Gk�f��&v{ϕ@�T���;5������t�l�iO�����,痖582�� {�T�?�U��LQ��l�K�߾�[T�`�$�����zb�u�hk2�0�ߙ����i.�������hQӡ���ZZ�lδ\I��K��Lvxx���f���
>Sd_�Xq�E�?1�w{�-<!.|��C�]�T3}؈��8֨n�g�h�V�U�ܺ*@���d^s:�ᜟ��y�o��nj������d07zo,�������R����K+B�.|����ֳS}���IԅT�g��L-�����g? 9���cdN��4�->��h?��tA1�h���R�����'�5�� b�ЁG�ܤt�A�v1�`�Q���W>�_[�6;WN9ы�_h���;�?h�:�� ����_�d��}TmjT�lz��Ѵu�T��A�4񒑳k<�C
�]f�&��!���Vp�bC2aiO�R�{;�*ث6��V2�Sy[s��/����<t��X4����<���� U�N�sMC��3�:E��H�x5C��!(fַMv��������5�Z������d"��Ｇ�KѤ�` ��eҝ�7b�I�t�QPz�v�X��'����/�T���V�A�K��}�pt>ϫ
���C�Q��b�1G�J�(ύ��(:�AlC�*��sdʑA����{�I\#�BRf �]1�Y3F|�u�b��P�!�]�9I�)�������y. /�}%M��~}x� �{�3���M&8�����.��vq�d�)��_@��������[QSWw�"�!U�gx4u���޿��'����!H��5 m߾��*��Z�RvV��hK��uj�!y�ד	m�`A��"��GK&�ŵ�&S
}��0@c�,�bzz�ZI�:�t0@k�rѯyA��H�A�鼋���wY�3ָM<"d�L��Ňz0F\&ǀ��Yg��P���<��Mñ��=E@pE���Q��k7�AԻ�M�:��f{�����mFJ_�|��߲�[Hw�YJ�z�D'���N��I�*�1��L��1���F�Psz�Iud�R �p��L���a.(��Fh���&¶�A��$��dp�jΠ�L�:��W�Qx�A���ı|�T+\<��n?�����7f�/�%@M�������Eu/
W#��Ob܃��M��<������N*��sD���o�dP��?�ǹ4��d��W)L���׎���V��<�`k�������.������j�!p��zy]+��q
����6�.�LI��{*X�����)ׂ�r!��v>�#wV&�wh�����=.�Op�rZ��9c{�m�=�7N�Y����_Gw�:�2������B����Q^;}��!��2�yfJA��@s[a	�t,��/�p��/Hcv�_��Y]�f�J�}x�\i�ڜ��*F��u#�#s�	D�0������F� *�Ə�\��|�я�=�-Z�d�@�0�+|��<Z��<�Ԯ_�@���K~��BJ-�h�{xG����$��筤K���8����W�
s
��i<�����bb��	�}7� � ~�������Ʈ���ݹD�˴vÃ=��g�ѐ�7T��7O���V�s�B^��3�����3�	��5��k�`��㠿���m�ܙ�>�;<K��u!��� �"��M��Җ�v�[VO]���Q�*����X�W=N6j�i��Ϊ�8vA�K�i5�t@k���7Ӎ�����f��֤fҁ=�(�Ѱ�)5��$[�Z�<�d��j��x��z��*6<2�:��h��+���Z� t��Ķw��d�N��x�-�� �	^�^s���*q��7S�اS:����Z��GP�L�I�{J����{��o�>�NX�]��e��1��|��n��vl�!�wR}�rc�P8Ϝ���ShC�@���h{u�ՙs�n=�{�	�h�xzy�S�A�q�H�X/Fˤ���&EA#���bs.G�0��K��T��ě����G�5�W_6���ƾk����P4�Z�0�ߌ��s!��HS��v��Kb����2¡�IxuWUn<^�"�&�Ii)����>(u��������Mgz��,fG[��>�'$�ک=������_e��V�|� ����)氪gky�nV�[�{r��-�,v��ٳ�^[�ơt�),"��[�Z�Y�9�-������_�߃�ܾOa+�Z@[����]N��hQ5�^��5K 6�&�s%��J�R�6�ǽ�3WrC�֢9��������L���{n&��ȵ��qp�1J��d���?�oK܁���V3䚸�)�z��?��3�\�.����K�r��3A��QV��&����%d���6��V���1ߐR}3�wYpE҇u���i4YS��YV�&B4M��=D����~��՗�u�;ύ�����f#+S�m]l32���$c�%��[r_PI�0�P���]4�">#����¦"��Yá)�x."�)i;U�'�+��aߡ��GV�7h��p�u�S��'�5��)n��L.����%0W�)-x�TY[��3ڗ��`�~gA��ܠ�U����|���X&
 ��l-��f8 B_��Z�p ��g익� �)�)�k�L7�Wg6�g@ùӷ��g�3�-������[�q�F�l�s�����e��S���z0Yf)�丬D�#�����W�4���t~��Qa���)M@Ux�]a1�r�<M�㺛<e�q�3�6�i8ක�'�p��ꑦ��C���(�&���ߔEM���/���Һ�m&�t��^d�9���jqi
3o�7�%$�?ۤ�v��b����m掬����Hap�Y��r�A�e%�P�!z�c�����H��9t+��j;�,�,��TCW�:�ɕllq=�J�0/e��+ً@��^��>�������:��]ă^�zڿ�uB1��͎��W����\�f��<�����j��v�5<H�Ӟ�|S^�~��*8K��N�۲ج֚l�5KĪ@!�u$�5��~47j���J]�g�{��U7D�X��]�2.�di��GKq����U߭��®
˷�IV2�k6q�R�½�:���J���M�����Lh��O]'��;_�F��t���|ĕ_�������u�Лs�6Rv���ϭ���[Z0��|��-Rz��u`�>xW�%"�v?�x^2j�o%(*# ���-������zW�D�0��9l��m�M;�t���Rv)�^�]���]����&Lq+���$:�(8�.��>��ohﷸ�Ţ���ȓ�v���x�G�T�FC[<���1K@�¨�X�IT����*��Ǡ+PX3�88�9OBzs�<f�\#�u*p&� �;mU|��J v�,4�&y.���hqLG#ΟFf�Q�\C�̛v�QZ\�|%Fy��q=�Mov"Q�a����9���6�&X ����`�����?�6R���4�۝?~ɪ���xJ��}0o�A��1���k\ӯ5~�N���Kw7"��`��ín�bqk�
<X~��WwJ4C�X`g{�ؤ����Y�w�1���k�jK�jr�{Hg��<���ů�n����[�3-��+w�6oYzX��N����2;/����� ��R���N�.h#�]'��#���5@Dz̟�J츢IM������?�o/�w�IH� N�=DQ����ؕ��j;��n�/o���oZ4��lHb�����nP��`��M�sC�u�!�0�V`�:�۰v ��k��Z�)�+,2�T)CI�?��B%����Zu�.���)�s���ʀ%~�s��9V6�T����D���G�}�v�;�W����
��q��;���y��~eā�{�'�!^~5�q�/)aA#߅�`�+;�����$���bf,�Ɉ���Z��f�*��74��W�E]��iXގ��T����YoY����$�8f&ή*�߾�6ek�g_�"0�q���Uۇ��b���&+4���C�!R�m���~�fnG�t��s<�_P,�t�Y%'�C���'z��۝N��V�j�Xq�f��[CTp;r��N��&� #�-zz.F��(׌�i N�w�#(7��I%������0��/�Ywv;o���̯i�3B�_�i���U���1���y~��c<�	S?��	cp9x
r��a�NEDV���@�8�:��J���b��hq��!��b�˱7W�;���*ɖ�{
l��*�� D�H7���ú$V5h	�ks��E�I2��
�m�j_S����<4\4#L�$������97�'%�Ծ���!F��7!j,��^���|zǹ�������.��T��3%hX2%��X������uI�x > /�'�bkHuTu��2�ړ�,lb�	_A9��b���!�o�n�P��G s;���HZ���u�L���2�e[/��`��};3�=��z��]W�V��AB���D�Ύ��<�L����i��s�xgY�S
�J�zy$��u_Q��mK���!���l���-J�zT6�hVZI��:䋯+��������B�X���T/�I)��ɦ�[��M�vhȁ�A�D\�j�sD����)�����|*bXI��\m�b+e�@X>/Wga��y4+��LW^�
��.v�q:��B�y��ub�4>�Ծ�gd;��@�L�{�
�r�X 	����oa-S�m�m]�JL���7�ɱy��kK>Z�{�-�K�+��Q��T>�a҃�����Q�����P�,36�j�o�xK�q��-Y��iՂ�`��gZ�5���X�����|3�vK�u�4�~�2̠��"2ԩ��{��+��f($b`W��6q*!td��U���ֲ��~��`�I����6�랈�I�o[E
�E�m̀�^������{j��	��<��ZT���V�u��N�TN�-tiрZ�X����.���`�;=ye1mʽw<h}H�6Yh](���`[���;&�YP�1���萶� �S�'�_�n!X�l��!��O`��;�3�f��%@	\�Pt���}�V�zG��='���`݇־��W�����zB3}r;���d}����Ki�:
�,W��@��ax�+�h��Ԏ�Y$S�|F"��W��)Z1z�D���s>�t�(����#�������ΰ����l��<;�3W�����L��^�IFZ�m�M}B�a��To͡HD��U!V���Dx!��mP�v"�m�E.�����H9�V�,݌�p��#և��2�G��x�v?!!wN��g+҈�o1��WAT�@�t�)��\�G�<G�>Z�ӓ���?�m��ǎ{��bj�$	��c��[x�n&��E+z���F����z�r)���̭��q{�@(y\_��v;vʨA\4��E�#r��"���y�;�C�ǂa�ze�O�~e��gad]��m'��L�i�mO�S��h?��tDp��	Z�(?ޤ��3�g߫f�2�d������?��[�"����D�M)��nr�枕I_|�����>�7�:��_��Z5Nk�i��� 5Y|L��r��-�{���Ӧ��]S$������O�;Fpu*ĺEm�رs�lx�b��+�����6cR��$5�,�{��a�)�jt�<�K�B�c�=��<ТA��`���cp,c״� W����84�
C	y�^Q�9�ٷ��_��b�/i�0,�^gl��oN6+Q�Ӗ��U[_e<�'����Z"��d��܂�:�����P�7j�lV/\��P5^L���­V�*E��,���,� ��d���V
��.u%!CӋS�r*��Z���z�LcW�J���,�r�w��ǯc��4W,�W�,x豬���>ӐȲ��1@�/�^�� T�ޭd�F�7H�@5yܽ
����:��h�>�S�1�H	\��
F&��N���o�@Dz�\r'u������I�"����N�]EP���DῈ��j�G�k�=��};�����M.�1�V���C���Ě@H��#�D���@wM2��ٚ�(��R��hzO�m��τ�ew�%z�2E,��5��O�Z����{,]�I�O�ģ1���T��f|�c���a�կ���[��HN��~�H�gӊ��<c�3_�� ڠ��M������)jg� o�M�j*���BC�	�"�9��e�f?����X�jln��P�lB� ���C*�3�\z�`~7�y%�F�"�.·�Ht������\��[����L~�ʐ���~��P����n�ɢͬٍK^[��&	Qb�:&�O�k�XOu_��? whg�Ѷ��T��5�+������W����~�6��P��9 �B�3>�Ѥ��k	�����jL��$��T���;���,�9���������?F�ϰ�,&�E��ڀq&c�q���6�)��;ڋ��-�