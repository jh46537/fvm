// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Fl9v+xekOChYXa8+6HZCJcMGLe6+T61dNWdnOSTbPiFTh9ds9PHVw2Mz3FTnB6P+
3L/7FpXE37XMBHJjPXXinklwkvxU0OX1zH5gZflWvJXbMv0DQRe64O7W23kJjWU3
bVNEimGxhBO7w3VGyKVUJufsxkS+aZtmmr1ZpnlHD2E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 28976)
3RDPFhp/PGnvzFbgUFv1BZ14Fq+sh9mAu7QaeOWNUJ/wBm+S0aKQpK2QpQFI2aL+
5zar856ZRRpg9WHmR99wHDEBNAtazQcaC3kPmIWx3C+ndLGocA/gIxoyrOHm1S22
GCQlEVHNyl6l8lQIklyHRxPjhZ/QeZcL4BfC5dsvqnziPJgZ2XTWphBugsPS/aor
572Dw9c+EB3XLkQoxP9camg/xOKVGZ8ghioYYTI9eva98bNEPfMZH7xOp/FrMdzz
y9+x/1J7yL8BjkegWWRYeSfxETLtm2lyK1AyIc7GvDFxQscJLASj5E45YaVuJtMj
JH502AD8u6wqJz8uTuQgPU1QqgVWf8BHjhheX27THlYsODl0Z2/si3PpxZE1xhsP
d6E1qYVu07cK8xpvmeG3WzvwVUS7IcZkl+dwDZ+xfZsiuu09oeuXW6PCJTcnneGx
EXZmItsKr1HG6sH/YqXYMBVjOde2SXqPdaiAdswenwG1xtfZ5WfQsR9oMjIsgHth
xiPChqNsBhWyB0Xy3MUJ/YMzbLHq1y6PnFWbqf6bIEyjlUajW5S9nG0IHsVh/Ifm
74a7fruuVxDZ2n/BpZLzwKv696zyhaLywO1y8FDA0d7Jej+jqxwRMws9KlKYb3QF
gUe2jXNKsMz7C4ZaB5aF+yg96pbp3c+LfZNe053vlG+9bSaMi6oQwx4q6p7uU8LB
oncZ3T8c4V0LTmqBFeDR6JcGuiRVNfMKC9I9v0Brb2y0wm/sazMXWGkNtPyeu9Ya
bhgT/cUlHodMoxRJrgsBvBelhagkyym+lBfiSb5d10aMa/z5Bxkn0imNsV1iVzgZ
3GHbTCz3y696Df40LAddYyd3FICw0EXPe0XCnluTlTjcdtuN2KdC+WDUjC2yr4D8
r48j9U0knX5CG0IC9Tc2lA8fyMa5zrQDPzRKEGYTCnJwZXMOL4hvw7U2QFnPWjTJ
IDPYxWcg8PQxTVHzxIJqAgCfwIKb6oc5/WlfFqPvvhSbt78SK+yUx++VODDI0ox5
wQKMimDFyLanl1ocZlOGJqPee8vTRBWEFD6VjNZJjK3OD3i5dUsjlXFL+v4Nw4WX
uc8KqrHQ9huZXu8+w+74DRl+1aYv4K7c7LSnm5t51MLNR9gPaHfSps5KvcdH86ro
KPwdgUvpaiyAGus0Xfr6uFnOc4Ak82e+Dq1aB90rNcUm9lK64K+lbOsKSZ9rP1Nt
Ma4qsJeS4lJw5BFZYMpwqVP+Okxp0mVD8PhvFUx7NLzRr4AGeDG+9pAdwz4Bfq9e
hrETZeR0RNddlVubHPlMBYdeYE0WMReQPt9E71KZKL6vgSkAUOpyGvRXwSYE4ofl
YA1lKoyAcYbdgnaqhLIR3/BxP2eSXs1efH9WGaEgRM7RYqyO1QyvN9wjE8fCdmW9
iFHypR3JycjSeLzn3ZNzBY5R2Rh8llBKvIbSjkz9skUA/cN2iUrAgtl5vLRKTqAA
r7sCzfWnD1ljccd3Cr/HH/Z/CC4QLK9HaRr969DnIlR3/SPE16FqMNNwM+X7woYB
XkekZV/JIDKHa1vFfLQOJenDK+Q+MmamaIeQ0tUZmGtiRUWSEhEX4vP+clIVrlNV
0jogKvBjlCzwZfoW5nWY49qggiqYxs/PptT79PwPxLOdPSLiVe8d6aSyS9qCBcjp
z/73+A5GO/U6NFxh/HAYLpnBOlzzhgjt7CeT6bbXrFmVt7bNGn3WGD6cJYjv89jA
qDyj8xzA3Fmum9oxH6KoKbU4mdFqLV49iu8X5cDiZY18kPiP5+gf0c4pykGKUQq0
VV/dl9kXR+780grpbcLPfkpMvnP/O9xqJ9BLA1dleTrT6zKkC1BTlWfHuWxDT3fn
9BBRRA1J6MdOpCP+qk0o0CMaVVBtjCaXV+yPtN3IxDKeNatVmnneuehhuZ92hGe0
AQkXlhflgTfLOw4ZL2OhuDE8DD/FkRci0OzGrayVVrnf7HCsFZ5Q2Pgj5G8X0US4
qLsHgY7YR9gVu7bRciIHcjlLZUfwdxppgX1AOG/67psFMklmw/z4BCF+l5sS4jnI
Bq34IP5hY2EZJxen0W+a/ymU32RV2/8IqRSMBCvgVPeJ/pXTG8Zf1ZyRPdOGAwZ+
7tqg0QkR+bNFZ7Lq3FuTDc5IYHCX6wEpUmUIOqOQYS8LwQLwsGBVGc6qT5YrQlEp
kCQuQjhhZ64GC+PL/oD9o75WBdjOiKxZIahcqTm3KE0JPWtXhmkS6oh/xY6SWeYi
ZXpuVbgwVrxbHts5HloQgGMdlyXMQb/uu2lhS0KwNtixZC/zM9HMUtl/Xex1cfMo
GCzWBOkBpDRU6TyZTZ5fnazNaaPSnxF8fAFWv+Tv8ueiojiW45YZvzlg6k7HbeZu
TRIiv+r4P4m2NV7tr0piczYV2nvgDA+eg4IgmLvPMxVg/FR33ZwfbCI2b+bx/8YT
B1U/KXgLQ8RFLIMUOZjwq8Fo0dX4a1Ne+b3Y/cN6hCDWNizWv0CbHI6m+35HJoIc
gGbBxQ8B5CsKgoxKc+whUfwB4TLGmgOYBA7811ZCRHZy+bp3UAWcRiKYkqF/Xl1O
kXFFY5gDGljrhdYeL+hqmeAGcfWCVUnvjjBFBL6CayIh94tvRZY1usTH/zSWI/5z
8cxPB9bDpFCFuTJYkC2Sj0kANKx5ePiIaidgwPKI9wkY+uL+JtVVZfcNcTZjBnnI
pHKdc5h2JJXEzVH4G8u4wD8v8lToFJOa14XUP7XpNnKSD3bS3QHLQ1DE+YyJqiUt
GMPtSrdjWnu2UBYJpSTat/P1592JMJxvKdvG7w6YvuSD8ZEefLLiW1wwHB7vG9+Q
lw06H6ui4wSTbQL/RDSRTwdhaCF5y6Qv5utdRhroPgHdMuPM8w7ALF5Y9vYow3R3
U8UHZ+sBWu8AyuZWnjIvbqwxwGFxNrlAXHd/R1X7j4s9l/bfFkynU3qAQ/HF6p5F
bfkzrELRfg/BK7+qPPpYeqTeTzVsSX/joFDRHvenOGu8jU+UFNslbYl7v9pmTysX
270sniPfZnDSofs52v3FhaNXRUajbqBIJCdnxlYS4FBdZWC+zaN9zyyplUHS8JB3
Y0dmO2vfdq92v6Bd8y/lADUUOu2OMdCv7ghArGKDKvNSe06a7cVmRI8WwiFSbEvF
euezRIsCV2a9D/IsV/jes7fdRJVuFXSu4egZyNrsDr9ypDqiTF6mHaP1eVtBGOQR
6Ytat6UnQ3svZkoXt897bEf57AvDYG+GCuj/54wtfzQ+9gZAfCwRJVUuLvEvtQg2
lSyGTo9m906FjX82fO1kjZMnNb7jlESIvtfuPZcuJvRX+nFRH9tHXvQ1W2wp1Rrh
9Zwc5y/5udoNYSL5CJ4iz3/b8yleNmi5Pl2n4FiPFSN3/1xWsH6WEGx8JOWWmAv3
geZK1VIMeJHv3dDZu2M26/q73p+zfBi4EVQa12dcFYNEtA+0xiQnS8HCJwoUoQD6
M+ZRPuA4v0nihBo2ql2MXaRu8DuGuZFNo1r3bLFHaDjnSglYE+g8lOPxZfi2Scar
FtFWz8bVd84CqL9SEvMxuZdcK3N/SEV0lWpnOUX3OQOUNsQ+3pzHDAQnCKDwH7j3
2ECwfYcKhd5Az3wiGyrsl1YJ4XY7bjiTJ5uETZ940TgIwb/nPXa1/FpC4XJg7Nz0
+rikK45jUGsxBoRu7Bi56N/SR9Zg5CyEqg+4brbV9GNrNFpAhg8AhxcJ1cCCA7yr
g27JvlaDTdWaQq7idMulSasQtTRAqc+uKmEtxITi/GzAfVZ1bjAS2AyLi5W23fO3
3V9wyOxuV11HPC8HDvvK/L4CIr3Q6EssFvW3ce7gmek24yT7BQgtFSkyCGuxrQmX
r7C/eMWdddwiHNRTOfwQiQgFbY5lMEdtYcIMkKLXJH9KgfRGIoYy84XxqSQtYSMp
pXlKtEhmw6nwp7gHzoPohO/kQWw4CbzTco+YMjvO+V6jmvZy+vNNm0lWRYinCeSk
N+cjUp4q+cjkkw7vVDvD1cxzd81EEuSIV6/zYRgYaGYYwUqEtEpORD/P+B7G6SLU
A6UQDWmJ7KLTowy+J8amIR4j41H03HLSWJGhStpNDfLawZVbkVclo4bTzOsrI5wc
x2xXqqT3Uf42J6Fy8vbTeS5F6g6cns0LaxWfoywX5wOHPZ071OgmKHvASh0q9YTy
pdhvpNXlCU79Kw0eEROlICqCLaJJaNYU4B8DDlUx9YufIfPlokV4sRUAm3g5DTZy
/gFXll4qlieQQB5nr+S6lKwaaAy4Qp/qJpPaO4w+Kpfn63H5iD+hkri9d37XyUQT
7fsRNl7fynDZcNiGj4+79Pvh4pUlSk/uZtNnPVZsjHnJEm3rw+QzN7ucSDc339zk
Q6piCQLY+S6NhakrvcDRiwlvtx4Ybvvs2VBUUfMdFPfNhca0KpCQHalavkf8MEAU
1qkUbKseimch2LHAMlljfvLZmUGh1KFpwMtSYL0VtpPoboQOX/h9Rry8iV6FjwM8
ViQO1I5CNZhXDB03zxU5SXPdtA0Z3MsShZnKAhxQGx9Nn6KCLsmKELqFFcuR1Fw+
iL9Re0xdZiv0HN2Rf6xrF9fcGVO8PS+JuvOukFOxSJkjnZyKgMZzUdu05vWJRPQI
upJ2x1RfYXcTmiM9PvGuUpvc7kqwa8AkXzw0DJ26nwyNOBPY+Qhba/lWFrwi9r54
+tER5eIn6uC8xjL6+6Ecuq/a0O3zaqQqru1FPJoau9+MUQWWbTc5I8X0yzr747r1
zpZr7OqEjOlJ08nPuD4dD/bGNt5T0QtQdkjDLqA6rpd+jNa+UFHn5Wd/7JCMTGly
Yp6+8yGfIJZVnvVyY+aALIyU5Mx3GwKArUEUe5tb/0+QZA9COdtbDSF1cnPzMnXa
IneMoTrDNB5iA55aew3uC0BOWWvTnbjTiN46Vu3louc5q5lvyr9Uuy/M29Gg9HJr
OZP6+j42w1ICI34yRLJm7NQtkaa1RLa/64B4OleBCETwBgQCDccBtmFVJAfAiXJo
0i4/oLho/sqUpI9z+ZKdELx6ZAUAKsRnTLYY0YBb3dMNsdIAH+QZBmslAeymwuka
tDslfSSaSZbTTf9XDlUx919RYat19dlZMzfsYH5QQUxL17V8RffUp7YNMXEB6xEE
ANBO3SWyLUmnewL1mIiN6Kb/WylhDCOay7FU7nav6JK6LVN1vycruedJvc22aN0j
yTwf5lZWjYIKOVtEAGExvon4BJzFCy17IzstIklKe4+32ANrw7HEXtoHJ/FjrsSI
Ur4O+fjd8J/NxJqhHiEbFAgIvdaLiB0SfJFhf/lTEn87xZOTzWlfJnbzuo+Ap3+m
VpY0Y4DIu+33F1VMzA+MiNxJ+Z4PaJGnahnzJm0EC8dVvuxpz5aDelfifZGhnq+d
2zz8qMzLDyA6H+Q7GYrBp9D2EAaF9DPa4LYTax7T+oQJnoaxw67/N+daBzgUXHIk
W1pWTUxGI4wz+WAj7ZaWtRuc2ZWaceQRbqFffT1VsUKd/O6Id/UCnfMZdfFyuH4/
HHmpmkhW7LcC+QbXvk6HKoBrbK+rPEV99vaSpOX8jmP1V4If07aZHCqZD8TubGrd
zLCfJQinkarnuEhY+qkLycowNCnB3mvGZFzfHWYJyWaZqgy/6tJOE/1C7sOiO6hv
51TV67TQEbtUVy9qY8zOhE2shTgX/S2UbeIEcvtkbgLZiMu/DD70gANQu9XzhctN
FKb7XjdC8SrTihwAPzEt6EpOMbsF+Yyf+XjQXDC7BvfZH8kN+VMByNQYqwNmGCDe
s6+Rudq7DsC9X0Tvf21GshgWbEyo0RBmrUVe2GNSd05wP1zintgrHg7g1WuPcJOd
JD4xF9/FvhMm9hSFwYQAmIkpdKKonabolh/wfZqT//AGDUY2VLw3vg/GVpGuyi9e
BhtDiQc7TwIqdcVsn5VDlSCKRxQ1+YuLIJezTkz1OhNzLlr4b6Q7woeLGSVa+tqH
9a0ykdxgTNC2cy05LLcBl9Wwd3W2Iu/GEy/9Gq1lBZhYQHZy4+/Wlm5g7j4UYCZ+
uF44+K07j+fX6fIgzpwmRQ+pT/FeVBERg9xnF57ESlhuZA8B38gJCLTvt+FiXdrC
bQOCQt4oY76PPB+KOUgd+/GQTlYRm9J5U6aLvuu0qa9BnOIsHQZzzdn3yLFVDwWO
13cZmhwIXfOCQMztjeP8YMvyGNq1po68pkjNiA6e/VbQemIti0ShBNVGvh9cImLD
D/b0J/JyVVooKuKAMmoybOu9Xfu8doqUnv1aReu1O6YsagP/iTzLqJU7FyZAUt1a
tSjNB6NHe3Y7EfB8HdxUvv0ZoIwiOQffwnVVKWmxjhKi+gpyf8/IyRtwfRdpvk6b
ogAW6f5klr89spyqlloRc23Tm53fZDXticAQ0NZ2IJsJBMRqQe2Re2zWXzW9fgnh
fNS6t9PQlLRTWdYm+qFWP9ZSs/+5UBtSxp1BWTSAy+n5QN+MC4hOz1vremjuBXZZ
E067l9SFSUhNEehCaFX59Eqs80TcNoL9wQD/uzCgGgpilOcZQ1Kh4hjnyH3LzQfU
TyidB8GEYxN8yo84zMGZaH7b54hj25gf05n1oGvj9zdwr653ehuDVmKUpSMDQC39
ZAkLcIlCyjiRIMxXBEnG+Iz+FAaVM+3UX53BRRK0truIgjAj2r41YaJSJQFt3Nmc
he+zopaN47vM1hmTBtnlkK3Js/lNQUeGSWF3VlpDres5T2sRD/dag0BvLyrp5irX
vLdurBVXsaJ0skIzRrGioDKFpCyV0LWt9mDcID/yYt32L524ShIyWsK+hRFVpKi7
bQdy5IJkQOF8L2pnUwvh3YeHunLkdS13BgVElD/JkrITlMzSIr0lKSiumG7MpeAW
C2b8OgfNvqaXCoqNVHV8z2/UB06VMWSPDpVUyh68z2mMvBTCpXCnnN0fL1CsWRAV
Lk26/sLWsXXF0fUupyEEp0tNxFtsR7aLsf/izgYg5TA/MZgMoOicpQ5KhJC+VG/4
MxXbzJktQ0vjTaNWDQ+lNHpnM4kFrjMEiBBR1p5LxTQP22Mgi1QMl5C4ftgqY6iS
KIILa7ZM42OfDtzwlOyEU1fq60p3NlhgWH0rl9f1jzxxgoDiyavUi2HHfL24OEaV
0cPo00rDLDH+TWZOLP2vLZSroiIPN6Cbq1XWPvU+U9Os3SC++3ALnFHL2sC2Zmsg
PCUSWsLX+wGRQdbpZOif+G987r97oS1G1FCPGSaW7StvoX4Ws4ubjUzgfYK3UJzc
gUKk2tyBznKMYYzUSchLYeR6FsWT7eZVMG4QOO9wsNi56AMxa2PyYvleQ7xGUxVq
7er0bNg8qeaSLm+QdXrapS+qSshMUW71CRXZfrS7W1BOzENW7iFp6MuYfAQZDHrb
2hUWvbDnexDh8yHiB+Khhc//JFD1Td8RgOPYGx17Ayc+YgjJdO9mIwghBkD/LfQU
hNqyDfwBntgDQzZtQ9QpihuV76Ipr24Jk/fAsfaI0/guPszai4Q5z9Rc9CSJbeUF
No+b62qRPLAlrtXdTMCdlLT80BHn0HZ0cypRXm7pev5iqtjvaAxuO/ynoTncMSAV
ygOfVXhe0lJCUGWCwrEYwy82fOZCWsaZI7koViG/9u3otfX4aVh0/hnRy8TW2uRo
xvfeczQMKZkZ2NXDfalih2YZnPiWuNd+eYZFgO2ofUzFRPOaOFj4lF8HfKeiZF6E
2utqKdo0XoZtX1+ClU2IIHaPIE63mTK79g+2kzvQn55tN0gv0tfAHb+2IgxbN0Fw
CdflpVvHkRGERycqCPYo4GkkgkNNhRrrhAdRsbknUbHtr+5g34E6GIWxEQLgDjqS
tgSbzJn7Erx7twATUWdm+lwpKrfsP5K0Zxcgnlhh6tx5tFdXlgx6RgneZNqY8zRA
O6HYog4NWC9CY7b14Awx9rUfDVfpfKZThCJeUAsqoezbSBeQSDDtM7QzEHbynFHG
FeUYla+D0XhgJAWFT3m1dr4+Nn34RdlaZe0/NVUf8/iHr7zvyMcBQ95LKMLCCiQM
a4kkgkroE+7t1XlnxO0YUsL1w0Y4SIFVRi1lWE9Wn4qY2FXoFlUaogsuqEEc0/+1
xWp1TidbcI7SoaqNn8osKUm9Fv+zPvdczr/eT5BBMLia7m4Ibf/PIY83WG+lTAMy
RA4SSRWhKS9EA+ILLkX3VfXabq016my3XGgk6tnaWNEgdNEtdGlth9H9e2yrImX7
XZJY/ZWlFfA/Ihx3/jko3m0j/PLx9tqAZpLPVXgbQKuF82vRtE2fp5IBqfTH6uWj
SSNWPPS2hcvdSN9zpNU5MzBJ9+e7RgJXDWNexjd8vuOLlMXrdYYolJu+QpSSQxzI
roS3m+vCRFqrBIJxAKbhMwCN2oFh7m7lSenO6YzuV0gkgFa2SSeSQrchwqXM3F0Q
+voFwmJsYME9tGWDMJO+Qi/B6u+rozfb3bJ2PRhAlgSyixWbFKu/ULz8E9dOyLse
Ngl3+7RVBfYken2No/EJ8Wc/ETPZetW8Yw5Zur6U0xxQYT7VD8DtetqXRLJ/5+pn
mXOXcXD64jIaqYKCNhNoU0vc63IVNgwP05OmbvM2C9NHewXal3CjBCdq2T5RgdKF
5QDqTDcor3CAsVdQlciI6lySsZt986FoC6K9icNwafnHjRhvHepx1BtqNYO5jdO5
x+FohrQwG8elYxnDs6iJuug5s6hRtjvcaWogJCcHN4cVZp8Mvak4d0H3C1my+zmU
P26x7C8vV939LRod9RlwAFqSoKuqXiESSm+P0e47jg5iNKgHrxsPlgu4gQsMGAuw
xi4PkLbjmoBtfbna96Bjy2XipSfX78i2Ko13XGN4Ur4Lnwfs6d0qp1KLhuXV5WFN
tpXQ88v2ZW1WSNjdkpSVejSdAjOyZux2pt1xzRIOFicQcqMu6fkWr0mdcltJIq2n
ShIFbSDlKh73Q7JBgDeJW1Uf2l9nRpDT/wBfVGMpuSrXpXA6kJVYLmIyRWDH+imB
MHzze11toDHXjnQyipVbfWE2tyjFOhSbqKflzLPbHvY7i/8n13KEmbQ8Dt9nWYiL
v6uIwz7QWXYIhsv/A+J1Mx0dMivUQqcOoHW3530K3O4kuR7Ojo5CpvHlz2UGkSiR
CLCH3s0SZllhkeG9fJd+/XHSq2L2ZqkyCNpeaPfydm1n27q+O7kkYF2h6gwoA6XO
Sa4GmU6SgPU01EBDBbl0WeNEql3unKOt4mbi2EJO+udA047XnpjOHqDsX0AV6yeW
91RYuBLD5w/ZsY9eMlYKw5UDsakKldJ6k4fSorcAc2j4lMSPi1rnLhY+ZH6qFl9x
yyLo1bjXTxZedi8B3+ihN3n3CdcW5voYjm1EUWdvSudXPajja5d1w5tbmylTKW7u
WGgu2WVfIw/A8U7OQldQ4SW1qahLK1munc6NPddg65Ai6X4OenbPdFkm1qy9clh8
5aHIlHaJCVJjZsCCxkrK3EupBQ6ce5k19BNrJCgbK90+WhbFO0J12ZbCQopCLbOi
onIfh75BFOL2TfJnadL5UN1ba04BcNNK3S8jqlYzv4qjaOC9DGelMNlflYt2H/6m
isDooTe9qSeUrc2SceIb5FPMrnzLyNaLXxuc5oQn/OFEI3pLMMY5r8x5lbHLQ/ys
LvFmc6BdZpE4jT2Au2ACef2MDx3l1MTn7uS2lyXFO7CNkReo71SnsnaJGX22OrWl
LqLddMPGM0ucrs9vSbJtUSaYMmQJsNbLua49egznBOonswg3m6g/5YFqnwTQnb6A
PM28OjFAbIoOmpOMRi6oCQLLS6Gc8V1iR7R0F994YMxdE9QDsyCWPAnJBd3OPr+C
l5+Mgx5BljdD+3YNWKRar4qzH/bHqo64H7FGYowkVI7vghEhdkM8YrqRLW0NRb26
Fm/w9szdKVQWkfsO/zfksYyk8wF7x6M1rkZ+uIdnISNERfbahdoxeCwl3VUDc2sq
6AIIq5IVvWwBJQrBiIKINTy0jMm0CFmqdJr0bd9FxP6lBjekfOBhYx3ToR2S+4Vk
vbRh8qJQYLJ2FWgznQlw3CB1oIDPDKXR1lw9zKEQCx068hhYuCxlrDFFhUeoVMDy
+iVf9WlO59wdcO7KmRrmcuuHF8UxHeqgdO3hl7e7RTBuuExG755Mof6qxPGtOFPG
AbVOjHTSg6B3HDV2SsrvmUH/kWMyQtXpCKN7iJo/U9QmYhMPUHsL8SOMsDvHkemC
nkFTYEQ7K9v27iOqvcSm7UaqD7nnrtLNahIyDJTvDHVASYjb8Km3D0hWX86FEwap
dxPzfC93Y7Qx0p7vhKK5IVCCQd8JQDZ0YiaNZ0B3mvpa592FZqO/l6C+5rjnezfm
tRp+yk46C73BRc9ihFLwdkm9/7ntkJMGqAGrWjea7nkAd5KiJdnbP7fT4hT0uWvY
xyQZPqDZJLrCtInuOHCedQHJU1znQHcYCgKZ2zGXaCUGec/Mq4/F1R/uY6suqGvm
P/xRwGKDpGOF6WgeWRSHTbXr86DXtB3lsvC26qd099ocBSyoj/fxSft97kd7L+Jc
eWxDvO+na8WkZHqDsZhrILL7h34olb1lEUCRmze5wf5sRGlql103ReUps1pgYYA1
NRiML8vpITp3s/mdd/v7UN379a1lU4jlDeNM0PWZCrgeoI32OdFV5uxOdSSaFlh9
ZZDDxPbgDuTtuoRiDJdzmMLQrEimvV7I1aXG2S3mpAf87NhkOFXGhN1EU7T7mbd2
ciD2uUQNDR1bGp72doIDcpHESeLDchKFoSY3DX014AIy8CHA60/Xb0nf00kqfMjP
ROmCKiE3LNCFn16YY7+jc596NRwTiOfIypbTHCyN7nffwJ5qHtNwN/6edtCU/PRv
5cNqR1DMFErY/QfG5FFX4Pt8RBmIRjo9J507jTq/2D85wHupnwcRrpCQo25RXJuO
FK/ALMC9q09DHbNwtHQMy0ZuXEEWS0TY/NSrkRDlmikjK/6uw0r3FyRIx/Z+rDPX
kclba5rcuB+n0wdCg1Yan6awiQODcKRoimq+so9wdpmYFzUMP9sTCiROT46Pxlie
yg9wAoS89iIMm+9Z92uaZji/T/TIQKVERKYQy7SHDJ4b809p/EnHxsCXJqRf0RUW
9Cq2ab8iK7TBDYB/boCQ/ubo6YUE2zK4j5ahnrhrQFlZqPIvG1/1ZLgDWtv1aj7u
1BeVaOOgne07pNDchpBlBhk5ozLoJITh+7AX7AKI/5jFuhe4f6W93R3muLnl6Xvr
djE4/5enQCslilkmbvsoe4dXA+92fZwVd1csRfkr4fOrdYhpZqFcb2aYWy98kBpT
0Q9FG+9AW2/66QN2YRDx4oM+ppFvMv1ymdSGpzJSBkXYf0dRrhVmWoUXkUZM2TC7
pELnALYurolyt0Rmnz3qC0S/lY2/ZHNA/kmJPp6f/UxBK9WXgk9Rj97ANu/VLstC
azEeYTCrJtKr+RMBQJBaVASev1IXIoxDEQHgpVCBlHFz4JYo1fGL+KKfcZcGHOJZ
NN6J1jrVT8l+Yxe568ITtDbGsqYSVlf3epl+MoY+XQiRRNYUmCVQ0T9EAnMZXXdx
BFkg3x3Zp5mf9IluPrG17OOVqz4Mjs1Hvhf2WUe8NaANSBFKXwfd7RIsNX/9CYbf
dS5cGl4C3exMbZ550CXW+A6HEXnCw8QicCA2qxfXJ9/0hltatUYn3sEcY1VQpYnT
xatexHuA45DfvvZ1Y5plFSlgwBZXE0sZQEd1If4+oWiVX7oUZhH/lLKYw35yq8Iv
TxjNi83ErjmH24U928Py5lzQVSuJUTV3oIFZVXjiGcF7CoQVBf/i6oQ1NLOeGsO0
bssXJw8/DDLXLm472mXDocDyCktFQ8f5FLcpD188lPyrv6Sv2/U5k73PlthwwqJq
M1HSVC8eTliz3jHrSU+s3iWaI19UMHAWoLKz83RE4NQ0804lKcuflUct28q0wXS5
W6i1fuBqmRQCH3oc5U0ClnyOjB3IuUw2gKpzcInIsdjaMx+o/J1j/scyrzy1macH
+D0DiHEez6FJsq+ucWk0S4RWqaDa5S4yIJ4y88G1fxV47FjCmmoe9CpOan5F7VYX
Hogw1pcJPahXPDEfRhYKjeUypSns7kz3hq1teh85YmO+JF9Wnh3Pb6YT5HAimQMi
WqF+++VoCL+322N5kY4e95K3wFIM8ucIGGG5l2ZuMi7FMAmx8bywXygpKl81Xr8R
MBsC1lq+940pVxb5iIiTc6IHnJnQgEgveYRMtDZdcbhKBhS2xImqzmlKpfza01jZ
7ZqOftyP/RZZkpxQBmAe5c5yIbdqi5Mml2YjOuMZyQFooocqdDR/HnKiTGrQ7OXH
NlZbdHyEBQNUI1f7C0u0Daa1VaEouO1erjUeryC8Q1b9irnDIVZnvzsuwCAENRbB
WUQmv3OolPSD8duqZUYUvIGObfcfdwHIVqA+GiC6YKMxYZ3zEf8R15Zt94IoPqMG
noqmgmDyIW/KlavZxWnLD9+yeHhHtE7w//fVeB7+5VVLPiTgHk/XMOBvxfMSh4KF
ovwve9tssXOOqum+DmsVDdtlkmTyZTPWfG/5DUf6FBo+xKQvghjag+2EO39YbVC0
SoUWKXnE3H1Bni78IWpHAxh5WSr3V2+ti3+a9QeaDxnlawg2yYlEMkT7BplVQp/O
Zr78K5PKciQChyDVXGj0lgX0AwphYV+WExLDf/QQ+YkPvrE/DdnWPZABVRQQIzg9
JLM5YpUVtFj/B/I6ooQEMWGKVdrTbLAMqM8JojtlaroeuMqv60ABme5J4vjhbm+F
NKGmRteBkXruxv7d9n2H7dPEP0CktowvsR3X+M0eubXJ6kB+Ncy57kstG94HaDsO
41zSgVMLytAC3Wl2zkoP2evJnBOEbWpHV3nwAChWG1nJuecOSQ2B6or1pgQYn1Xa
0m94RXg/+gXaYc3fXVnJQE60FPglfZV5qhQL1B97PuLxjk8nkVLJSm/lC0Cv0/UA
zDDscouKerQQ99kKK4MEH05FZfVcKIWfaTlG0+gfUC5Rjz0fI3PR1A9+fdjb8y2t
2QX6JAhObRSTWuGmobsovqcOAkiYkpD0b3HTY7yR6+6rKlO3IFnJZ7qERNTgygeT
TVa+Wky/Hzhg+Vn700YvRpMCAmNceghM3Lr4NvrhrYICDGc0AUcu99+QmDTzmLoI
0KDwrAyKTWsNiV7K6BQcLh0lyOakiSyR2rQVO4KEofy6CgSuSYks0OhLtpAt696Z
vgBvOr1lbs/LG+Kuu55/GysZZy8MQq2D3zGs5iMxGirkaYdqTXEDFGBgRVoRj4u9
Y2S3GT9BFvhuVZ49AlGN3WemLRmpgZmAUrWX7z7cmVXBfQ+ICfWjrE4gkME86V0V
uRiGmRDAblAB7lBZWdgPo25KiKz9dkUx/pUfxDFFlwGdeqMFcCzjzzy20i0TQVSr
GPRM+qiWaYcpm8O1s1ACKSCDiyCEUf9omkUFK2qelWboq8vhJqop2ejc4vx6uSyz
m8A4pMvP1RMBv+ADPLlBlNFsTdrkEYaBBtOzFH2+T68KrYmSZyGTTAJPIPLLSuAG
Oy+/rdJ4b6I9Zb/jhZjHAO6we4saRNwsHtmiXp2+kq2rmeGFI0UclvMMe8RUMQS5
zqIOafu0MnpbMX1QZBMptfqRz/j7xZJLeH/OGK/l0VkO7UJkZHHtNbZ7+McX8iWZ
voq5BddKnosf3lIeAL/OKRojpBDGJEZEGIa1F2ii9uQmAEgfR9saWiEG38TaHA2s
WFC2VIVQso3eu3fKhDqoVgj7A+10cRA8tzL2wpJuyfN6bF62cSrvcj9xilGCLAKt
WO9Yx14EuSDbJunVU8RhMg57MDufrJBC8via9pC/93VEveU4YI6UGn9kwff2rTcO
R4gDde1L7awp83YscY1CUaonq02CGZD1w+/kJQMflDUf2YtWhSJYSkxHr3iyJQ6U
6h5/Fih7cFbBSHydS2w8GDVKcZm2DVy1qGN/zoczKP8U4U7Bw9yAetdxeWcHO1HH
7aHZKpOwN62xbppUX9rUN8TYuMa+d9aS07CbBHjQjWalEZviVfi22dhD/jlqPVrq
ouyFZX613fAKMjRHOa2KiPIB+KmLDulluUmdQclp30ZJLFRfgUE+Svza77/PR4lC
P0Drq/SirY+ILyijIcpbDjNw13iv5KEJi/h2m1+c8FXrLNwOiuD0hxj5x1mMWmdg
hC58WCGwaN8wTSAAg/BpVWXgiWBaxsO/IGbpNeYEJ0MItsvajegAXTlRjsEXqIRy
FZ5OtivC3Jfvi6lajwqjSI/BbfR1JMyLv49m0h9BmtoeqWMIBSMaYk43fB8M6Cbb
W4OdS5NE1i6cv/RBCE40e5WJb0BmooXj06SeUA7CTPaQ6qY3XX9mjO9SIijM2PK/
ue/ol66CNcPj7uG1hWHGUmp5iiNPPPMbdnSGR1hi6H6QrY7HQApvwZJZZ8V7ewOL
pMkeSRu/z5EnCmG2X9Ho2ifQ7Y410JYQAmmm1RZyJrblIWMtgfXuo0mZe4oTonbF
l7T6jVYsEEiUKTQNeLZun4cVil109Jgzemteiec9DqqTQ2Utk3Ai1Wkh0qe6ZQzt
73BJKeo71P0W3E0A1tRV7Qk5DXfpFUoUBFfLddFAR+p4mG7pCi70X7UR/RO4B8lV
IcKcYoeXCy3tYEsbNBbLML3CtX1+jPoiTRyEhigKVhoRJbraDoI6EmZe0hSdPl1R
Vzo7mp+vFiP+Zbn90rvhcl489E9JlOYciCuC6Lb5zUrikutS8S7vjpQNnQuSVgNC
r1zDt6Bpc6Zh4IfopWR7hbwEhFpQZnJSe3IynfJtt8pqT0RsYpkoN8CQ/g2hmeEj
IFviGVV5LOaC/LDVxHrT87oGwF2AqeRZc818WuFx9Bnzaeyl/WOhdKb/NfRJFqAm
H9IsE5waOIIaF2CVKt6ELX0Mmk3QzJmP/KNaO4oddz36aMvmpIA9TV2TlZbSZCfq
8FbqU5S4WVSR3sxsOz+0GaYGvgTfzsK3IBtOaPvgyW5dq2PMMYUrYYjY4uOWqqRP
GJglBkQfq1VLRrC9itIKSC/8Z3Pr3M5JoaVIzOqG7GeNZLLPaNaZ6AT7U6z8QcGL
5Zjw5YWrEXWZ33BbB5xD7eONkB1rV1SDl245xqoRTcU0pTNvIXeshG5ukhwgFQvC
W3DndQGr4lCuzdqjfENJY0miA0P1dH08WDWAVrlrjYx1S3xjN6Iz2V7F+hl3mFkZ
k4GB8AxzqYuecFjSaIXLvltQAvzpr8k+3d47hqXu67nx/xSvQ6vzXGE14oLGpYQd
Gr+c+6V1B4Z7XtNCGZKXfIBfpNnWiISVuMou2379jOOHO4mmA6rW70Ti5G/XBOHS
alxiuFtm4v2J0BxqsJ60WXytMtf0FD9bYML9PbbfCan4hWilhmMqRnCXS8UC+a12
ehT4YttyKBv5lAzGvZ07Ucs8cV9l2G/BvOpaHmaqhBXUgKUIOn+uV44SoXjvH61a
TKl3NDI18kN0BSbzNSEbmn00lJJjdx1hksuNuI3kNEWhQBiaxoMOtJdzOMKr5F2l
Ysq1D4HsjQeeoqu5jVn7rBhSP1PaP+TGDPpzBoNrb0zD6L1p6bTZK6mYVBQsTuRM
mFL5zbe7xaAG+qZYWstTQQyXwoFRP3N51SWzHd4+jV1pVRzIQeZEp8OXaYpYkAwd
FdcvRqoRDn48dTh4Rx0PefTW2uQntShTrt839pVMMqpXkdCXIh2THElW6VvXDhPd
GMmS1otozmiltk1e046iPE/LXsjycqDSfVlsMzqzm6ed9c7eMe07Zu6fQm5og6fp
YMZ99kUMlcCBtguUlFMiYJCppUr0toAFGwCIRLi21ugOumMv5UfvMdGPL65N1j/G
VtqhF8OF9efrRqc68ibXbUjriVZgPCPeV7+uV9ctyGNJT2iI5Xjifq1Zg8u0zxpB
68jLeubyoKUnPoqOu9VB16/fdotmYsT/HiZGnalmm2QALHygg4GB4fC1Y1EWYQhl
g3lGfPCXVTc+Rr4+V4hvxjXHTa24oEPxWxv9t+R9aoGZwzumfyIPQ29Yw0kxJg08
xpg+mhzfHzkchIAJJU/AGxLBVUzZQixcrOnG3yIL5eD1eRcS6YwG9PaElV7U9Rxy
LWaAgEcZPpISOcaVEH9msj1JO4w7TqfNOPfstTQ5w3LLlmKkFm8sYd8Ue+lVweRD
j5y2nPeE5+Z1HjWQukLXovp1clelV6l68epQ7oWcckgK+arcxvSsVPqoP4/HCNvr
LOXZho51eDONbrqpV/Mc9AIzpXQwGdgNC/zvLiH2qsaVzx+XFmGOI2tE5X+veHJc
JM/eVMZUZB2fd+GHaPEu8lj1yNEgaKDAdwzkhAJIi82P5RhWSEBGggaqflxQZfeC
XsfQgspJqekR7ixc4aNPTkpz+HHyVnOMCUhN+tuhv/HkmCgpvweLSLieCAdIGYfY
cWJGZHWcg8lMC5nFjX3aeu6EkoeOJt0ejB7gJkjQo+VjbmKk3YAqJDmnhtuy3IIP
N6T3CcCcp5svPJ7a4MqktAGOPf72neotl0kcvIxawu9tL3c2kWKnVu/1S73/IJT7
sCXywjDM4tticnF/TrF0uj+9UXRT2tRKSXXA2nxQhezR0YlaV9XyWcO0h6ZnHToc
oOQxGv04Om0ZJ45zNhJVqwk04xGfOLKdtwG6hqpzH3g2bxQ8PD8jvZyGzEl6w5r0
12VYVEnFIIiefTlZHAWwYtIcEn+EObZj8ZAXELtwRtZwXV0CI9OMZKKejfUWeUCV
/w7ddo9mDlnIq3EXA9sjs9FFPYMpoDeFxyddBZd40shP4yR94KKtuG/STUpHoTYB
+dseTSuxbVZ5Z6/xjkiQJ2M42Hs5dNktpJsWoP/RqFzIoFeatLIEidjDZ4drANCg
/lAzLrZSjWdjF+eP85AnYiRYk6nPbJMv2gEFNno1jz1j1woowttsQTOtVKjreRS0
M1oTeJZHD/5AZWP0+3upTj1m0v+Sa/h1SliWM73PVUv0jJKZ4aU0tMxDoGY0heqM
JIrH2p8BcgO1VIQ1tGE6BwILQc1qSTN7H/1SaUPF7//NXlK7jktm35jZ2QPDc32d
l5kU5+/WfUQekhEYLJJm9lmp8XL5vCH1BE5gLIzKGZKUHM6dZGVTGofexkRE9gyh
LOBCmY6nQ/6Iai2s8q7Gd9yd84ZJiDOJqqtp9Q9cy+YCEgdSCtwu3vineghfeLfX
41iaqBkZQOeWNwgPYVRnLFo+WhcbyeG+QgTwWqoYvBvGC51iSELn9j0X46im4Mbn
nFROUrhj9jdUXsGUhFTXtTKjpKcn3mM8xD3rpvfSWs9hcNGLvohpOkQem2/bkNBg
4ZcqseGVrEwhkhiEEN+mM7qQO7xSJGEO3yO7oTDmwGGhbDuxCcCE5Xm5Y4T3okZ3
aqfiF1H28H/v1bmMpuyfvrmx5YsFWrE7pr3DqIGTCYRJw4OEmHRq96f/u75QHzUv
y+aheo+I6UQk2QqtBAfBdchUPEAkn+XfLpVEu8baUwvZNs0EuzHOBRkMQ8JFkERm
WzgF5v4KxDRUdNEhXtsPYyh/HZMaUeb925Vh1YOs4UtjxuvnSTrNFh14+hKnjAF8
kjvvlN6YJefd2ky82sWLTdgwtyLt2vNhQhIu1Z6BzQCg+Gl8jcbf1e1nuTwggo0L
Abe+g9/LZhn3t+7hUA4P60H+LrHBWjUh4zmb82evBAsJYq4rwyeXdfLW1LqRcGxG
/Wc67EcO7Zain6LVLn/2IHhx6f/OKRdXZNskCbfsnCvliv+YmaOW8cRCHT4qC4sQ
w9LICApP+AwPdaq3Pdw4hf/MFWftuSbILOR7cilhyqk8zHZ36wUqvNHVNjfWJttv
jmKcRs912fb0RXl+XASloVfrxkEmlwbQ+JeteUqlFtCo+I3Ay9V4XSOXHiW+rjZw
Il1zKTw5ZH9cUfvURH7U+1L7SeNgUqZ31H0yDHR8Iv7bSkPa2Bmp8bjtJ4vNr6np
uw6G+SDvUV0GFB8mQg3AyAfsS6rNUalA+zJBr7dSApFCqSDqRmZgwGjnavPaOnfV
Oqe2yVUVLslSVjDmttMe4Qt+KiNHxdIZmLGiwBcNFQWc1RCNVOw8g5y6BRBrVxtw
B8cnyn59NWZLN5Q3JbCK4M+Y/Aoq0RDWnhY8Bii26L3Aj0bTMZdCXT7Z2oMtm4Aj
WEd8nbX8CH+gqGcZT8viCxj1FYDkrR8EypR4QPqlvBnC66eddV4G+oXrMiv/dVIC
a+FrcjDrJedRd4tcSz72c4UPytW/0X3rQeqabFjAuUVSW8VQSoJH32YDPe+KA6ES
as1YnGs6za8M6IcIrRZ8lpMJrSfdrimgMJcLpznj/+mZ8O7Ztu6lNFTivBHRsYJG
SX8eN8tPppbTydScmJW6FKzUnsaBCkrPFkr/bJ4nNZk9JYJ8XMx8sRYypQiH0pnG
Y13FJmXEsqv3jz4/58YuzK3a5rmkT58SnX4Rv41x3FfuO9o+DpWvDk0cp5An4XQi
cX5FvtBwXJn8l0zBBRFiKaAJ3w7fa/pqmjZN4E1/HvHAwXnT3ezFboiPoXNxZOP0
E3hECAlvND34CyQxWW5M+YOKyYEPB0daqE0QeXrhgPi8OHof/gCX6OEOXnJgIzA9
YE/j/dxsRGy0lHEF5NwZyBHvSD6Wl5xv/ituEMaGtcTZ0CVHIrdS71fArMA+Vtte
cMCMt17P9MwjOoISW3hK7fV2l+vsZP3SF8nuS/VBO0H02BEP4wYx2dOKQHgvw48r
lGvTCCCQ1RBmgpBvrq/O1C38e4oceMsfwSiWBjVSNZjNIRWzVwqy0eFDHNcEZ+Gj
+yLcC+Wo1dCJFPqXI4kuNWp4FExf1oO2HdPUcO9k/QryniUC84qdG+FAjTTWfika
GlOgfSfwo8d5pKcKgWlCST+KGke6Ma3bM3nfsF7W4BaH/NolUL+n7ul8CM8eS/rp
ZfhxLf1YDhKnSyuKt5EgYGSmSCgJHRGRiljBLElS6blKcJRwWbJ2fFQQtrxE8E46
6lHfCNaLyKp2rlO/Dv5z6QPCfQj1Nsjia8d6KlHfe9ho4cV3Wk4M9TMJtyEF3nyI
13KRBvOFMn+n5TzDqyzENXF8lszeoVdE3XwiNnPfKaehRd+JaD6D+DoDIculTmWG
twNidGzbDjqQpde6Z517ZMF5Ob4vNerlrzgYkeJBbUOp2DnvAAtGguhtqnxFLNYr
gILD24bIlkAUz9ff0bFAx7TmmmlTM3qkWj7rMyLNMd8x24WwoqSYX4N5yLgx/BkE
vX6aNIjNNcH83iXTTlzl+IC8hNvlIjk9WVqMzQYAZ9hHw93ycVRsU37QLIm168po
fA/JvfwMIsdkPqDvTkf+EzYAl8IURx7ovyAJ1YcYZzkmV6xt+YDr96J7IEGXPpeh
+UFvf120m+HS5pETGhwgJr9FXqebtuEjmj8op56knrziok1sQz09GMyouiCxhHLp
mUb9QfeFll90sHAiEfrSHtmKZdQgIlmHlZ/nPOXYCnNjZelTE0vwaz38x/LHqsEO
LprrOkrkMzOk1OwSHdtaV8iyCApyZjFV8qdzhNC9eWCgi9be+m8IXRCjnCcRQ+tX
HVTCWsQQTxmmbBHapz1cBjUWJ2+CCh7MZLuXWckNDamCfMEdWvuK53f5CdYUmPqn
mm8pdPuKRBYijilSI7e4qeG+rX33WeNRWuPsrcxKVd9RMthj5TtA1GAwukP+FFRQ
5Arp7AC38s5Nm+9IyNWWaIEfMZIDGVjJyLncaBK7vT73k4CQDE9GiR9XCkbPe06w
EXq8rHnPCnpb3R6jNBuXQBQIgbvh/LmtIdM9Mw4RA9ni6Xknh1hkKHnYvErnZoRf
E/swDlzJyKQkoLpYWeGvKmAwrEzV3mL46nEYM4iN4UfxljAfkxnurFA9o/Ao+ioG
csYWskzxZHnD7MGimK9uZrRYouZT/BoZl8FoeVXx1+mYnfbTOpA6ugbRCS5Gfydj
0ygtzviJMBGYl8RZjx26662ik2cZp/Z2a9XOPrhBlfHwQx1xkW4NI8Rtg628fqpg
mjsmMTo3PGDqZEMmypJqgeOK0imr1ZzcH0Vrwnm/u7xXLGz+BVzeCcwTsm3AnxjG
qeRZGkxIneMpI1f60J4FD2wmfpSCsTDV5nYiFq/VGUXQD7L+PtOGiDKNszNQQIY6
tbQP05FR3AfZ0DhWAF4sWBJ/fzY9z+1/USeIsLvVHppI27ezu0j/98JQ9q2Zh3LN
MkLDXmSBVSk5DHZepVPLz2UsH+BOov1MvCjkkdXkPOTcShtXy6g8oIqj3S+5+NX7
rrbZOrQdqTQ0o9j8XL1MwWx4drzcDaoleqmqjBeRkKdDBmxQQxirPomgrHDw/dp3
1TLIrXHXqiWbEOGOGPJVZLX2oEgN4idiv3ZY4qlKKODtuVE46ZhyhU+atshuKd/A
XxcicXZHbqA5obIMmZAIGiT0JRwX2yfTyVUkEdymQVSIBNTPLs59O+t95eZPQNh3
SXKlz+jKwxnj3PhHJC/r6DyL61l3S9Elo8/odqt6cKCBYhN3u5h81k0hRv9ocKjU
JRDXYH1u15RgOLrbX9GPxYc8BjJl8BdJmj2XRVoOU/qQf5cKf9cqKvlUz/OP6Lsh
29oJ7npXPADrsbL7bgni/jLTDb1DnAu78Q9ntoC5q42IMvNCWrSnb7iHVIc0Snc3
etHEFaJUjEKXAmoklrVNEsBV0BCpQB/pmLKA7bz/sjnH4Mwy16beFe9xyfxgBVld
zQJd/KSdWZtNZf3KdcTKp+dxMDBYrHfAarl3zRsSUaYwvTohI5CxzUDi9k/528Yg
kLNoEWBBQcAq41oRMMiL+CX8wUnUe7TJKQdEuWd3WA5J79HBKWrTwsDmyXYpjffT
QZeLyFQUK5fofso/UkaeyfPEj6gejN7W7IOBt0GF7bzKfYVRdHIqkiPtxuZU9Xoc
z4K2/7PQis9MOCNc59mvKyfODBIQP9nyGoG4QjZkUDK+p/8I2PNf8pqrgqYMGzY9
jtLU1MASv4U4abb1dNqfQdRNHAv/F9igUJATPzLM9u0xKdqyO+Qy7ZnftglpSGEO
7wywtRwcz86Fc1uQ7ZY5p2fagudEo1LT87g76Nh9MOqUHeF6icBu7sff6pvzjDn0
iwtEHVKwnRAK9St5l/hnk9eI2wVDsekzHvpCmMFAX2+e848Q3x3hzKRZGgpu4D1Y
GuOsutBPAJTt5fwl+GIzF40018A31pOCuSPS9gq0Nm0LSC5hjK0JyzNYqyNFnKK+
MBxFKYeY5Eg3FJwqd+1xYs+6PXHEDzJt8IqFvUAo6IelG2N8xulpKeV/T1gDIK8T
qzN0SJl54nJXPVC2CEpYH5frzN842E9wNmEJsXTVm/MaeO4shswIlCa8LyAfr2Cx
VFLhd79eKaX31pNcIvMirCFzpJl/fCJnc21nMd6EQ14x69LsWcEZQyKRZM/gccr2
H5ni2NDbsuHYfjmh7itPDKcV4ZOVg+1WkjeAWeZLI1vSsiU1pDMegjljibpa6Op6
0vlIdQS8J/JmLEzuwQdPiixmrwgtp/eoD4St0KBMyZE1Iq9HdG7q16zbiByLnk8V
VMVHAkuRYU/oAeLdM4k6Fet+GkMlZ6TtJhLmjoWHJPE5+bjNOFyvCqYPpTuvGuaR
GKiYyIo0m260GKwWb74SiY+/36zWhWAb2dVN5zS4o05l18PufCK1iuuUfzQdwwo2
UR8eEQ7OLiihW7XZq4hA6Xra18ZcJt6MxP4QGHoWgqi2af/v5v7WSgAgEk6OO9ui
BwJrpWisVeb4FoZN7TY80gkRMipZ3hrXuAPhfZ9yHmyeSbFgxAa58UNpfGqg6+ap
FtPJmOxxsJr+HznT1TsXd/rN+FpKDquiGlSjNmxp+FpJ/58XOskNhGppOGtp67iE
XPg1gLj1DtMs4HOKrVP2QUkfVM7rO2BZ7Q8slR1Tff8+qoxgA74JprxCb9nLEJVG
Rfod0y+Wc2+jnWYTBcSz31AIwbwJGDVvL8E9RSdHstN3g5t8BZh4X/Qx5C1GoG1o
grcL9y8S9Pl7b9/5Xl3m11lly/MYwZ8MWkqijtfbgULFaAKUMkfsV3w61VQGQdB5
PzuHQMSOBYtKajvxpshoDPvUBDSy7JdD8uV6Ljy86hfBDx+X/Bskb3xNP6+L1bDx
KV3xvLs/pvxp+T/RnchkcJ802l23Z3QTqfGJ4CZpmKlSAPU3EeKfuKs/+coXQ1R2
f+f6mgM/xa9YSloZAoLdV/zTlGMLJUcPNZZGGfR9qCKd0hS5nZT7TTI71t6BAfUJ
6IqSLFdg3am/Gaj4VHIn2aumonISAy8OJNDzHmeOtwM/+jX0SPPTQTPr8bE09h8e
SyZe15Q/yU5YB/n9lV8oOuqgQ6Y1w0oL88MLESsCR0K4TdxdsEqfwCg1++HLcq5a
FddwE2Z8UBZrgyp1yXzTxR3/2x4TWA1wmzlzvIRx5AhpcOS0LkSLiVCZxo5aQ/Cb
TNKOqbcnhNLpYRZXaGEQRpX4cW1S6HsTQbrQPJ1B645sQvfZlS9Lhjf1nd6LwWoh
B+RefVrFs4KpHdjjKhBAYMdQwlvbF7GfMhsNj6m/NEQ4x6tPotpfqDzo61vq97Rb
caKhebpwuJzjbOK7Zf4auaJ6jD7mhxn5VCzx5CfCwlp+ZYDe0AAVWZpgLNHCbYzV
+v8do5BtPafr6ILw60I8eC8pdid+xh1h+w8JMD+/9cEY7OpGAzIsuBe07YHdDvAp
sMKHyrinUuBonCwBp7rtr72V7VB87SgXxJGFQ4N/cLFfHKvF5hz+bFIwWgFAxKFc
e/4HaOD/s1Vc4Fb8vhzPlG7Jh5XO2HCHWF6YxuPGFSX0xdsnGkveQfSbuaxnpmZh
nyG0w5/hTzlApYhKEir0W2duD2pAGwnHf1kyPOU4vq/io9OKycKyPe6y0JRQ5TMf
HTDm7j7Db7Q1UKYAJIlv4V2YfrXRTP4NKdHFpS7TEe0tJ8EUCOdtSYYxYUDGxgfo
a1fK4Y3Bj0q0J/UtJzaALKY3PcH8wSgfrsVhMihFr8Ru/JvjTHbqGXr3CGFXD6t3
Y9t3UANpUeIIOuDQXjPVpVSE3YsOijUXFgWUq1Vq1dm6XcB4mGEyaPjBf6mkzVGH
iVaitITM6SQqc+PfOZI9JZ90ifPL5RZD3BufmZpSZYvkqW7NNTWudfG6x3AUwy3I
nnVWt3EMyVsU98pXgOPryAn1Ksx0HN5IJKN8QohFB+6N+aH2vKfin7RCheQdkFuZ
i9P9M3N3ucKY0AofvYtDOBMhTn3CJX9EbL3GR9FX+Y9JWkN1BxoPdhXXOjpwBM6q
SB+JmMyRSNBCumtUjElafNnKlzZzngAozkUzVjz2fR4mZXEOTpU2KzwUbyk07JAb
wZ2APgOOW4//aVyGoyle0XU4zoz7a/8nYaEDgRE32yk9g8H1tXjKa6cnIlpb51fq
wizB41pRajNUXs78SB3Xnekt6rzSC+3OWOfKD/CbNxaaVPteDF7KnZSPGrDaV8rB
1xfMDx5a+WmWzivzX7kplbCJEUVEIp6qg2qNNKdUsiP20wYfzgro/UsUeU4nKznb
1xV/LlwBOa5DoxGLzOmcEa1CwNoGvVQ2yGtjMcth6K/dtHbUXdn4UBQhAKEOHev/
WM5Wa5MkUClzXfg2NhShh0/7uu4p/jF0QGHavQSK7YNLyRqDfK8yzBejiBqJ7UAT
Ci2gZ6UIlgXSwOd3lwzHxqvibY7XmcfXt3kg4mqudrLvl8Q3BCCnJ9A56CgnGrPH
0bk36+GCEyl4AV7vGfq8wz3FT2sw5TsS/0fMN/Bbji2zWL16rkDJFsjIy/ep+s/b
q4FHxdU0BMciw7Gm0Dt/iSoR3lbpd6CdgnA4lAzxy81uboRXbeBbVhkqFMH3pxV8
tYZvbZAepjlOdgV+teWquCLulS6WRqGLzLMFLZ9ObKZmfPOFgztINLpudkBoziwx
pCdpnAbQ+5Bhut//P/phovmk5d2RPneEpR1k9tirWum85rF7iSqOGn0Kt5El9452
W62S4huaMl6SHoES7bmz5ncAxdiFGON9h1WgRgaZ/0UQbyJZvgKLzdq0LPSEGNkI
Xk3R0ZWLJmXFm+w4EekH+OCsNrebemG5QkJFZAR88v3qXVzkcDC9wAEMvt0o16i7
mRsKO4M1kEE/2OQVa6b0uSNbyRcvdoajNunGKutuhqMf6j/ILAAVeeED9zIgnqAk
fDnSEl9FgSv81NSy7I/fNVxqNmb405ssMvAwXTMmtX5kPrOqnvhCj/q+XTSShXEO
Ch2K7GihKUzWeFPEupQDViJTr/dsDlJHe7XaYzNzaHCtjXkGbS0TlkOJO1sx001C
bAsAWgHVpfpkQvY8V7agWpp4hW7Xb50Xa9bXtV0CKBMUrz3WXrxDqYzcfPc+Nc0N
5073d8obEAM2X4twpnv++O0vJF855gG5IDun8/chd9IOG+hsRUU3Ovfer/piKRaN
Uhe0Au+Vlla5IcC8A9+3OFO2CSbbq8yxhZBob+1H+lfHycLAC0q8N8AIj/hcOr9w
xcctoxENv+A0JqzMGGYTS/7qQyF2SXp6wOKaF37TT96MY7y8uWXeVWJ72DcfyFYn
dBS20IljTnv+I1QXnjiQqcy/ynSs2elCzz/TOYp0JMLEBvps46ZNvzZo1ht3WvvR
W8TWfth9tfjVZwbK27uVFjrF8ShwT+3JLWOy5AdoIjCo8o/lwyAhp9DFrGsNl/Si
yV9g+Iapd6b8nyAUWgj0ZFYb8VJKoc6FhZI0PUGFd+RaY2pIiSNK3J2MG5BWP8V/
LTWXrNioKZ9bnQJ8LgA887wm1LORG2nM2ouU8D2mEYe4BI5qi6AHU6V+LCUXNbGk
B57U63dJ7lIZo6f3kNkzRPEnac38pVaRghDZ0qveL6BjsnOXD0oEi/GQC8dt5DlM
OCmfwS/8hCQKx+wpEkj8FrABP082kqze/bPu/RTK7ojiOhnONM1OS4PZqEVCq2UF
LYRN5fe3VhW5xluW4Xjh/A9fuPmCfUk4cIyAUQn7ILxdo6hGKT0/aPmNZE1Q0YYy
brou4NcUvGogORqgKNi0JMpNbZ4eGxK+xZNbF3bbRp314l9xBROoZn6Hq8FGm3IT
QSvBxQLm+CJL24kKW0N8Uep54cT3xukofoZ7BcZ1bj4qM9LbnETH/tHVp4LjkFto
3QIBGKrcEdrR1TptSxBV3CTmdMHwW2b1NY1oC0VI/UIAtGmNzPpdLrZ60Ev0ymoH
u+mmOczi+oXDVEt9CwR9P6q3TKpwDgaR0uVV7zjpaUyYE0pnroWr1knI+r4lM/XF
5UD+lPT8yhCVnHz8muk261GdpPQKW360xfkhOlGtiaeb6c/TqydJk1p032g73k6A
XYnJjtLs+CDCCz72XCkFF3Cy6oO+ZhCRaZGDcL8I+G8fxQVS+oopHV9nby81uByy
qUkL7JOnt9hHae/1jrO89n4/lvgyp0UwqGm/1fB3okWODTq15LaJSu3tZLogHk0k
G3AF7eTjENPxrCCblabUUmqmsTKCS9jeGOC0QxPGOcd/QG0wqydVYwYoKbl7z2As
QovRg9RxHrj1Dg8CP1TZutvnjUGrZluBCiQop5kW3AYdz8eGMq0LF9WT+qFRFdqf
X8SLdaWrvNp4xBeTxD8gBLDFkKmcL1DFY4OmxfFJVBJ8aJ/ApCuraHXdFKhATO0z
3XMzZSifkmw1MQYLziutKWUI0STzmnOd5AmFNdo3twuS/XzrrYiuSa/ocfd6SdJZ
O27HAjFKxeRxBvGt0GQ8W+WOOdQeJGwX/DUZnkQMCJf0B9HC4QISf2kQbbAZRHb/
0/tAaBAR4RtWOhsD81OTRqTwvO9uaWEBFSjqOrOE6WtIpWuasL7uBlFH1RiuwX6I
Z0G3C4iqjfomvMMpKePW7SZc7GTAGdCzitNLRwhq5Raa5pqBza09/r4H04KLrlLj
xrX1WXO9uU7PMpYC6L9A6iF4kPUgxqZAVv5Bo+NWzfXQKy2PsTozh5D+ie72BIRB
PlIyEgEQQAZkyex2fkebjk8S0vgPijtsZyOP/6yF61UqE30JRA53LZwQPR+NnQ/3
sgPn2amKJ8BRyqGeXSZPrDIpXGFB9dm/czf1MrTtsXYxPWzknmkyV6zmxk774lQq
AqRnqHz24MOQ+m8Pkt4w5m+9qVSny/gcMTTQgIo+UyxNcp84YQUWsqVwA2ka1UrU
gZvoAUixxuu5yljjJk5sujIMVyXx/DC1ijl6yPh3o2K+BvFGF0IZ23MnXi2xdxhN
hzi9gHs8ACu28BTObLo2LeKcI/HpZ5XH04wia1LPk6xG9xW/F5xMXA1pheRIzjYG
zsHB72MbW/+KyGF3m3wmezVYntDkriKnEDS4BLMttrMcNFj7Aa81yD42/c1F7wMZ
fNIx6Pn8dPJ7lMMAHiS+SDMwyNlWmQn7CeGEZtoCm9U6KWdDlP9SD1RQ3ZbI9lsL
spkzaFmHcCNGlRmQ9xhyr2zXXFSB0xIeKjhWk2tVvedUCqxSeWTY9w4biPsjXziS
aOLoy9p2gQTgDShwD3dt7wfEfVAfG2miVw0c5av2+c5TprImRthdEM7yTvL2MQam
wMSwg+0D6vywYNxDNmGUseaVbo8LGTKXXr4vrxbDZLfQTmZq9NmV4JJgrFGQNR3C
c+gQ8lZ3+CKDM1pz3NCP2f1rA3jYfFJGLsm78flkGCeqorw4bFXoB/VfQZyeYuLJ
n1F0IE+1qaqtJCcAIlPgv3zIMUbZ+/+6UC3UfmrGfhiDJ/ZDy8TltGe4NFZgW6is
+eJD5g/JyzkY2Uif7ck1wIN7phT1BMSId0YhAWXz+KMjWi2n1I1/fG5jFZcnH46f
TxjCtS+hoAVQYDRi3uqNQh41rqA5CSOXoBj61DvZOQw2e8vnoL4w3FpTGr9Da4b5
i3r3xBPXPwyGjJSJCf7bDJLTyiC2S870BgdWafwMvSLTrgV2rPEag45fInqDrnkH
OJ0B9AUiXwYV2KK3cQmSb0ESCl1I+BaxkD/Hlb6JMXV6S9WWDdbZD8NI8zSQy9Yr
7R2ptXn1K5IBq4287yDl/kES0vLWF+hWBUBjHgDX02kY8qjYDxcFbGvYE7kuDR5A
dvqmhFrNQcGPFVZWW+KpHAb1QQfO6uEtwpo7CuswYyLHfMsytODAla2GJEJpuMR8
wspXqd6UxMzH/Low5BE/zGZxdV4bfVMZhCpWvHY1y+e1eSEzzkDu+fOCK8xqGmwN
YW8SB2ySS6enEqTbT4+mpU8718rc84aEelyI0WtXtNszOL+PQV/QvOlypr7j6qC8
Km1/csXBcJKXOm4keW/Fkk9NklxAYOVGz38DWSJ0HhMpbeJB6546I42vCnEOvTQD
Zm/K5oR88JKKFpufj1DcRH5JzbZYrSSTgZ3zwrUjOriFgdR6FOkNgX1n71BYHQyE
4/fO8HFx4jVmC413+/jnYhEO9OoJMuxx9p/Kk0xRswoD7hVtfoW9oRv12NhrAapa
SoXK/rDAg22oPoM4wcTQVkSHVSEOFhh6+3L6lYJaRYlfNU6Kb3Fu7IgkwIBDopSH
TCzUs4EBUWx70M3cIBktZjrCaxPwsaAaZC6awKwZujimQUUWWAi1vISO1NwOP3Jj
Uim6HRrYPqsN/PC1xDl/sZWcb4EJnQ6Q50nRjvVwhb0+aV6KJSWuFyNbQJpmjsjS
K+93boULmkmBP2d5W+evDyNOSNhpw+vCsIXlKlLQwqA5g4FckzbCnUEuAKGI2zEA
sqmG0oVQpviD7rjZhKDrq+dBzUY2mBZ18Ou1NQQPww+kRheq28169KdQaZXheZ6d
LT3Zf0nuHprPIS6Fklbl3jITgct5LPhxlPvTwB9LD2Ss+M2CQQdLIe2wrRCmvpOC
2Hq3CGv8QO7jln50YItTlr5OSDX0J3e2FOA7pbRed4sIXWSwgeGd8StuICi29AHP
Q3Bn+aRW8GQxZZAepbqmelsHvIceNW5sRbn+bkFJwI6vOWDIXfCQN8igEfvo/mbF
HcIOnjnOmo6uOea4nViVCtTf368zxqhsBC+VT8ICfHCFYaX0JhXUnThBnt/83+lr
ewpNWMnFXecjtdJy46VM9cUiGOqxf0KOv/1WJRUhH2tyWg+0FavHShjjInEjLHi4
FaqS0vs6nhy3E10eWCHfUtrzz0SRVk4V05q+0bys8294rxr6nOFVimM3jNbixdKj
F2W37fuJjw9VrtwiaQAEJya5EZRsoyRJdu4+DVzC5kSwkWl+K8IwLKo2302LrwUk
vscG7xb0AVP08Rp49ZIyO1hXqxcT6PrbXC/k9Encnej+gz2bZ1xc30W53djfaYzl
nGYH/CrEl7hAGNWD8z0A0VS+fSHVVtJIEi6PsCm4Yk1YIBopiJhc+budNiTv3505
BnVxKWXurollhUIt0r2M4bQreA9VYGSErUijMHMjSw0Nced8pkBWHcN2jI9tLUBQ
cO4UcEJ1WQMUuVOIfhNuVsGjzpVYoFbLdG1lv+2M8+q1d+DwP+6jZb4enT0yczg0
A9NEk+9wB44n/kw9RQfTbcIk74GNXlofRndvf2O2S/lb1s8w3WBd4M4UuiUCoz1F
oeo7JQZF5jviMwgvEofflHV9efWkYA30aUyKhl/LwMZgY5INzWjJwe3PjsRg9hid
RXADDFCqpV4kvD4sJhPBzb3xCiQZwco0RksJjyfRlpse0TW2/k7W1/qVSODNEttN
XNmnAEb7QdXsozQlflQstTEtZXAcBIR201iZSaKunNyP1TxSE4vMKXqM41PxLTVM
a9cKv0r+UvKeTc/Sq9ThbrPfcAcnAoIJM+bw/F6wX/+LLQDnK+IBgZDHZRWTKADJ
klNOCRazRAisw33mhZt50NqoN6zA1B6A3KRafTKC2QbHmQDcE5NaHUNdJLAovEv3
MyUcQwu6qlR80NTcwJbcGVBBot6JNAsHEZFhMEik7esG0XKaoPmUSpSxfPoceHw2
tOXkMbZyDn33XGa4Gt5bvecl3vwL9ZDR1d3cY/m7i1KlQeNBjX5D5hhj1+ojB5aS
YlfE0ojOoABTh8wW3VD8vmCv+z/TFlmj4HVuaBhZXdmZ7RmoXC3C7rZF5+4Qv04+
lUrdLsaDHsZNGo+KVpcd+ooUyklN13W5CJQYaulMCpnq2opTXQAMLCVKrCX6Ccjd
Z1aP0hvDEoaiMBHSP94RZhKnX0alaFWjVW2MPejpaQPJ6sxQJ8IXzXB92VoFEiIB
zlzEjCHc+EJeNIU2lsO8u1KymGuWm7vO6Ik/2oyLNIe+1SahDRtl/KZ7XiUo6xCI
95shyIzRNRO/h9uJH76Q1PKusLjJ/tUzL6TFCHXp3cTyi2EUdFa830LPX2TrOGBq
1V48FCUiIee79m+rkfA6qAbF5+u8o58TeNNaYxvONfMl6yd1FtPqVQ28bJQBXg+n
tKZi5xx7w3QNj62IoOpbA6y9N0hgT6BstZ9akEGn1z7vKO3CSlYjfqH6G2I+RaM0
GnA76rcPAZPKbVmCt2WkDkNfpy9bw/MccIza5KJeh0qS3AjYc0iWuFndrOsQ9nGA
2vVsL0kQX9GWVFwMIhO1dSgiimb1SuAjgh2MfRRX+rbJd3P5RGMS1PPlWswfs2Nt
tXjYKeexs+Q6C1a79UDJ0yodGxkIMTfV0ADwgxCM1Wqx2VzwafFagYnfrUq92w9t
fPpju3Y+Iz+qCj2FC5nt+zuSZ/SSO1Vqp+1GoVdGdXBcuPc2edWwKyQdk0jmtbnF
GhBu3Z04VTmb8i+s4E1Q6jnOHefI+V/grsclCMggWPxZuxbDRtZPyH2hWNF7Ss4F
jnqGI0VzYYJxPOlUeQfcnuJb7QCqf5m+rVPxQobIKTdaUl9gnkpSCWEmmNrxWX5X
ZYld3f6rzlpMxlsmYGuqDSQXSM9n5BbD2vWbK3LZkIl2Od0/u/DphQnUtywxuXaO
qA1ZE9eiZhEI/vzYOBm2TeQDF7maMwKIuyM6Lga8Lv3cZwzKoY9jECvnxKy53UEe
p4dsN/UZb+IGUQxY6B249Jan3uNBjjyd+MLw5y04wQD6vFukeqbhZzh88OjnJQvU
dcuiBw7sPxkV4YqXjewwpeZHGa2jjcgpygxRg3GMW6zE8FebcWM520wX/IcCohe/
bNvcl/lvRCbSybYBTT+sURQtsFWeOHB0UOB3i43kKNkApxcT79Zv1txXLYnXswL7
OLTFSgVog/YObszIkZtz5wT9MZytxvoVsU10aPrSqUI8ET6S1SYPbxOfXWwNdlrE
lMcNsJ6ObKQmvTGGmNR0jLEa8uTvuEUUpoO9aotPXBdWmUsweFvbuO7Yp6isBrTR
x4rzulaTfEWc2/PDgID/zUY+MYcW6NdEh10rVVlha9pgC58vDZnxVFNJT+lQYzxN
8qxPj6vD7sdKP7nZtwfOZx80m5U8rmk1gFbMOWhp0KBffXx6xX9xUibzcAvxc5mR
6en87vWNvqi6t2asgilg8QLQeZvtk1h8dAdcSoiqWUmkPrGzEETV/u0puQWAGkYF
0/WsyxYOD+aUhOj2fNXcMiMeB+7F/OhRdcPYnFRNVzOn0v1+7T5IjGJyhl1nlUAy
Nmk98IiFxpwvSdxO/61chgUe0yjUkP0x+72ThKtVIcQUwXL7opvcfOJvtHqWencO
iloB82F9nUDhlmywghvPNjukNIGFySbTTzXr2Pdb+DTX+XmhWyCftUW4HgbKUrpb
AzgDwtk0M0/hLUb399L0I6bOtmfC4VExBSdMsHfyFuQOCDS1vwWAKLJluh0AuLvC
qBy9EWHC/jsOpAj29TvbnqZNxAR5CnASgfyrCIHy5e4wqd+EcfxRWayLR1Y4Cizw
6SNMV6BD/S9DDdWJCE70G8t9sRif7KqC7YeOkk3dxbjmlaijnLBa8CxPIhU12VTc
Q69IPRVbi7BdQeIf3PCcQTDe7V60sjCWrjIEWXCO5RpPlixGFmQarws7YM1GCQrv
4NyoCXnawrSaTdsvlpU+lqUGA49bFDN0ASD5cmB8D4QVGofqFpRWD/ErJErjJQVP
MAUd/lWdh6zVlShP1KM6kKpV1hxoht9hxWk5Q1gLV1D5i4ImWCGtBWQBMVTdN88l
rDekLWeULLZQ1dAk7HaEsuYtMnvjZqKjaitK1UpuMnktItIqhZCt5w6/HW3TjOU/
eMitHq1Df1eQF9CgduFrQFlXtLib/Jy5VHMer3h21vA7F1QWnEC7/4QdSjXyaADN
fOpBZMM/chPwTIPVwdlHSDoEo0+76+UnuLWipJhsMDsl9ZWRUnbS7smWUGxC78Hx
pAZs1UrlU1SOedBXraIayTwM8vMsFuq+Px5jdZDkETlgQANQ94R4XiB1Y+M8oo/+
bDUAGXTrCifQ2SW16h0dTeCAwtpSdu5+zePtRLw4XjLPOKi9vlSGfDujlCWAI6KX
1k5fko+Ha17rjlmTZ7xJFK5Pl2AxoRgBWlBYjl85cMkcPbezS/6YZo1KGDZTUs3e
8XihkhBa7yydmQ0YNTwdCGtVT00F6XgkeGpQfialJy7WTxBpK4nvAKxnjhVnoEBf
L0HE61MBKVfNQG9wo0/+q6Lmv4tjyLljcXozysNFxea3SdbEJuAdKt4q0uEta8VG
gJjycym7gRF/zgV6YiKcUO+3OvdltJobSevDreA17XqtTZfDAB8EiqPp8MtGwtvf
a8EzQQgklG7AfmpB6FmUL9bjeDeiBaBf6MgiZv5tKoQu6FU4QOP5sd6bAzJXylGs
ZEoNtNKfh3XPkXKUvY3wv81EjyVE9U8XgPFnjAOwEECUZbf9D8mIJ74BXi1zlTJO
+gxJEsIr6hM5SKAmh4+SSJ5uqSCMNiAnylF4wdPu/YkBTUGJTpMsF4J17CfW87t3
g9J2z/14NEPAH5ZNtwbDK7gVRJ/cjXBAomQTQlZbs6b9pAfm67vbv3Yn1tIe8Xuz
tL4qVAq0PqWNxvTC82syPwcChMOlm/3R9SE9EY9C0sXd0IJ89JDaSMGq0I0XaWIs
BhW6WJ7s1uwv6InjX7bAo9b20mBcWAlG/hgrkmEgZz26ol8GeSkLVVUEn2R/eKzQ
E2pa9gariy1Jllcn6k+9l+3kE68yykGs2GQCVJiFlasvemX8re4HkpBNTdC5lo0K
2bX1GDs0xM+jeRYJfUXLS1ngEYiDz535P/WQyytRImnpAGSvc2nRO4wUD+s1pKnT
8RI5UsJQwp3+AZG1HkQlL0v02GXs+q1pzpDciJ7OfYtMPo2MIp6WwsNEd625G65J
QzhwQsfSejj0MlnObgEp9NTqGsE6hIe3RzXIP677wpHFcRqHh5lH7zA6cOdpfGUx
PAXvic2a9C6HoTEMbn4bEGZ0r1CxYQ+NWYgd0OFiuXw2iiK4Jj9JlveJMgdEIElp
zCX7ZdRb/oi8kxojocWXpnROjVRiY7YQ1r8vLP9oSB2bvIFj6jnCYCcX3nAV+6dJ
OTqY0soRUV+EwFPXafumzWMjBcOL2ly9gLjFl3Ord33K/+E7SjUE2CYbAIPMzkXK
i5ydYjAv3acGwU87IFsVFwKHtgKqUfP6w5X1tCBd3TfHfkrvh4A7AsC2HPjcAklw
xvQbzjDQIjaA1z/5Bf3hw8Mu0XUJnVcf/R302i+E0RFeDnAYF8FUmaUAuvWhEN4Y
I0ovJvrShXeQh4UwzD0zAZ7ynYMDNSBpcfQRZeuoQKWyLlHHlPVn7WtN75NYoLhp
lYlTWxNIzAoLh6hCx/3Y33s24jvAQ0GOz42dMI05/1F767oheJ9r+QpuyGOazlAf
PgmpFWQtv1QquNJds0AEuKpJ1uAp7CUZV47ZDScAsGqeYhTO6BnEBQHTJ+Pbt+7S
ENPyNchbqHbLYJswzt8d0WBK1xmlCwtZMPpFkMlkTJ+eiTu47OmemC7VZ0AqfyPQ
MkyIApQiQxjw+cYQS+PzVkGcyVxQzACTOVH02a3Zl1mmuxNk95bsBHxJ6KGpWxMJ
U7UW3OVTqq/8O5YIg5lKHEbcXN1aQsVl0WaH+L8DdY2lRrNixi1FSdToKNi8fMc2
JqnFm71v0T7oDUDODqzClHLLXRlQaj8grui8mvC0KFvNY222H5rlePkowWbp5qeY
tkdKxE0aQAC8CwSKACemnRLNIhw5rqRAWulzqgCqLDsx7h49J1/Pepzt1JVz7Qqu
Vd6TcN8lMMMBqybTTPN9gZb8uIGnoVJzYDbwBdmNRwLjiK4Aq2Pgh8n9UEEOI8Ms
YOu9Yp64/p3I/vE2Y6R3isVJUjB2kQZUiUvBdvCcqAfHAL+7aGq+EfTCyh+8tImZ
DXWRTG5uYlqgv5/1DCHKXHwBFBHqXVcoTei7uSZB21Tf1m80ioxApkEn6iBbOt5y
/vsyg1kJxSwiKk/vrit5u7QQt6YRqsXKdvSghX7tqjD07X2KNGgm/t6tL5EBnwTz
AeUZ1pkOJ2hJPjrvUtF1XPBwr1VD+wemMVHNleX0cVSqoLAguKDoQAzTzF1c94Rh
69h5IB0F8h6MM7yLFobF5K+EHpB9jm2eVRneLBmWc9usL+LmQe6AzaFcNHGUsY2v
ddiHA1BtsryDIZBKnKIMFHS3qmHuxbPBXacq8wQFRXTI649zCBOQkGl274NK4x0r
JF5RGiQ2Mq1y4tTn/iNJ684WSaozQtPr7zGbiPT8laOFIakexELvadjMsaFnN/LI
nelXBpOcGlapaIWQDuVdDQbpQguYF9deHAffqz5c7Sp9k/wFyqmvH2b19Wg7ij62
7hI7MZW88wgFxsAJK6qrZ5ccbFwPBoVTzbuvsFbP7W90XzIlx3vt1++w3u5dcCfp
sG5b+W8BrNn9XzlCQTVlTUyq3KxrxmunTPnsRZXLnc4UQauD9XYrh0cAZdpCMp0I
JGvjbcJhnI7b36Yx1QUxWfU7v6Yv4o4Hf+1Q39JYgDNzG73i47anrdbmfRTF7cfQ
kP1okZUXYaq3347kUYTXyGam1kBqq1l/sUumyl/FoZjfjNLIIt2sJ/1oJLypjwE3
XliDX5xrcFh0SBeHLBPDJmsu0Qu6lfN2n7+i470uBGgqqSxmunju6YyGV52Xc8E+
X7GKtludqQtuhHcClUFGPgvptYQhsI4N/S2iHyA3vtDsYqqgMMTGOXmQJl1FMI/Y
X8dmaTB0qA5OCB5VoZdmI6lzegBxZFD65ViRFSKl8xlub+vSkkV7HOOqOHpy3tnV
qzO19vZde2asckUYbsxFNF41hBwQC4EaEu9DL/B5bWVNBgTjSoR9GQeUTPOj0V6o
dY1xB4dYyJCQYWZyMaOteHxhhxQtV1l5/FqWNMNeAv7cNoZYM0zW1CPzeHFuH3oc
wgRwZBDMtad41M3+MTCD2PPUmV0aGhn/sT6PglTPqxr+MWQpLQsJmyqSuZrtLAUx
TgfqokwE21bIc9hCLleOHMv/lISc8YiD0XP0NU23rldjCxurlnwlWesQuywhRf1y
toLe8RaoQ8TpJ+islbHXG21/MFlKXK1qXEul4yudHF24USQ2ZeHGvc91qVMSa1Jy
gptzl7QnGkP6noamRndBTvmlxF3YC/21Uq9piBhKwIUh6Ox+515w26+QEDd4flab
sXEEpf0pL4w8sZNcJU3s1lXwzRyKttxCvug7QOJpA9lS98SFJqrIGW9s4sj2mng/
S4ku8hndZmdWcWnLFHhGBkzVwqmxFAZzf2eRVaO77pC8nd7WUz2U6CA8P4WiR9U2
mOmx2iVHxSaOjXr9IdALM01zTHtfCpc305j09JIuwpFuc9+DiSSAx9EvDFhgtxub
QBDfFsj2HOiR2tEjbQ9Xa+ZDXsM+Jy2NRz7EW/4MbeOYhBq3WEKaKhAN+ICWgBec
VXgTiFr7H3ac8pGjnrjU6LH+6GM8Mi5XLSiraUY9wUOGDyBVq5HaikQjV6mW0bMp
FyV2XAvn4H9SoQTHhJMcF46o8Zl8YIQ0cLR4hA3elf0cS847XBDiR34J0Q/5n5Qb
FS4gdbq97F+nWf4Tm53mehCuECnsIFrkdANbi6vBlkXoBdubZU6xTDHknmY7u0Pz
zMH1pkS3av+0wiqf1Huph7Pusmv2oIDRBJSxfah2GxQmlJXoI3yV+GBcfjUjXIbZ
RvMhXmJ9kbJ6Hi725JMTNUcAg6S13Hxkn6dVcl24zhHqa6RunPGAZmpdfhNznrsF
G2J5rg7on6vmdXggmgzjJcpNv1i7LAeh1XQzt2+iTv305HGlDuqeDBErXj3dIfuV
oP/UPM9CZpKYB2dxixWItTartiw+dEZXkKwnnyaTg1HzCdcQi4HXviOSbkd9X99Y
B1Fys242TcMCqXcD78DV2lHOyVqZT3Lv7S6P02MU/jHqBE0RzRaL8sfyzASdEJFo
aNjWoTN9vQmk3eGbs0Zm7J/tyox0g1UTGTwcqpTUUq5yAhh5v8/HRckxPcsKgUHi
MrdqqvvCq5tO7RC4nwPHOnsCi6NvnVLlZmR8q4Xw71+I6xJLKKuOeTjNShhFQl6Q
RuDVUmd8I6MYU+AddZeFL1SNQyCz1e3hT0T0BVqrltGesprn3XdsKsKi+xRlNiII
O4XgopKyv1QOcLAAIvKngWJUTdtABTTbbAL+A5CgrT+Bhzw7nIKBuigSJHWz/DxY
slRI/61bGjEgHQtQh+kJkyIrtzizuRzoYu6p9bUFnW9vD6Gngws2AptVPtUHkx/E
2I/k4M96V7X2hT/TT4eMLl9XdMM64A1RWwPZ3tJ+LINRanYhnVlcqpO6iOIazs/X
8lDTvE/IodSZXCZgnORsuh9BC9FtncrWAgsxiINE7TAgUYWY+zwwOgccNJi5t5Iz
T/cTAl6rVhuxdKffjMEeBZSEQ3ghlgSYMUTgkbck4VBRAXYazgxjtYL9OyiI5Qgv
/lt7dof84LxO1OLkP3FaYAoSI6/CtWa5sTAGEkUlueSKpvhMRZLDebokuVYvi46B
5pZZ60RyAdG4rdnR80c8uQDNgErMs9udM2CNxDYQN05oQ6ypaYMjjfSt/Z/ds7lx
GribgEvwTk3J9V3Afy8VfxjJgBHPR7NFqHKXaPRifR39r694YqqhfIdSusMpY1a2
F+jBTmNqc2Nnj47XXztd/p6gq+x2BmNw1L/RTVhKzP0pdzcww4EIu9zf45W/MlFt
Q1lknwl0fEeIZCRkXfiwGAAaIIA5l2plVHdF/Wj2aeoguJO/MNuecxliU08wyMmE
+0CWF2Uog9b2DB/hrz3xK6oEAOqY1TANj90uuaPa7DoShA5CCeiC8GRBRF7NF6hK
mCQ/x0aZ4SlF+jHMX6J0+NYcWe+lcoVX5PfD8X/Lt2RZOz99SqqadLJbNxG7rYH0
81tZbEyV0jzoU8KrFXW5n4671GwZRfKcM0ckOft3SOW+0kVDRhx2M0KOVdzJU2rt
A3MFc9Uz4AaeCPyKtDIS88wRfRx+ajklN3rOrAYCBOM83GIbKZWPQrEsCcocCNIU
TsphIWtBQIcsVh7wIN50TlHUyrcEYzcsUCTvpJaZ6cElEoItiD9F+knLsAKtWRNm
6yzMf6lSVJYdSEnkWvIOmE0jxn+qBMUjzsQfs3lPoBtIOLxPplFANyssdk+0hyox
dC3XcpRgIb0kuJeuYD778GyWPmaeoLW5UHbFLQ50zLTQsloxO2qjsAc1TSfmWxBA
fo4XgLQlUxZJ9nyWhqR2bbPh88shmL1ZjjxkUt5vLjn2fTPZd2JaaIq5nctZuAvr
oX59GHxVOqraYRRRS5J1azOgGMFxmQT7lFSlaqU2q7koavmxqvrZtXvzS8BNsCiD
+JNMG0HhJL+IyzH3CxZOS+cqpzXjK2CAllTg6xvJfuE75TGB6Fhrki8Wpp9rTuaG
PLvBoZa+9RzI4m3hHWEhO/U4pbABpWxW0WH3Eub/qx2HCJ4BurwSmN/fYAcMSDwe
tDBCAICeB4AjegJUkP8XooiigRNmmREsHvtlMccUPtJ3YzQJMpTHB7+DDiDGf4Eb
j7Fj/qVORRI3JTPv2nqsYP1sis0qBUp7g3tdW0HFMpGMBa5yesj14r2ugfNkkjes
C650imK/ZpepvEejAVGmDVqxyjsu8b5bDmJ/U8UWt70yc6SH2prX+bMfVnRywwqo
hIpl+Q0JI/XskzUtigrlulV4lbGglNT3Qf8Y0qcnuvSm6vEy+tcoyyylaLDNAmmr
SjtbACKdB8wqnUEkumWrcMRupdhAiqlv/XGE5AKGegxF5re6HoSMWKHXtOaWcy1K
Z1He+RR4HMzAtt0BxaixoQTz7qQbmKShMTd8bD5bSpjlkIxYOySo+Gl0X8h9LzzB
6N90DDoeSNAENZ032lV3boFszgVCDciplN554Y4XwadE4aQ7DXnMN/Ik3lrf6Who
LOsJ5DAPaW0pEdAB2QPuruYkztXGmg+9du72dVnvColgJQ1lyD5AOtHNRxNVfPiH
X6f3oFGB2Zvc5CXjTvl4rDyQzgMaliSL2binfMb9VFMxlXWvOMonY8d4duNwX1e0
ukocOV7nWPQu2oSDju68ueFk7TuKW+rIeGYRYmYQV0b+nb6qLHeP1hzb5L1/l6lS
03Js6DLGd1w0+Rc5yMKfIYOP0j8XQ4vuPkgHewZAN8Bahxo69WEkQTOyy6hYbM8L
g/xMT8DwcVaxn9ZIqhOvnXafymrpMs7+QocaWdkmlqAj4jYIUB+YLCiSbU3P3gd/
mlosYxuhLLC3/1ConxiuNOj10uEWTcz14zAiZaJ8F1XRLck3bOYurqrV7maBMJOu
1MCLcffQ3zdY2R4Lzko8jzRarM51n8aB50ZUacwNKOcJC3GJXSiQPK2sIw6xRLVv
2CeJ7A1TCgIeZNr2DJ/Kf9QnHiCkn/z6fYRqUxZqmGqq03BR2ciPcghewvbSITKI
30vKBvLcZhIHUVZNcltRkE1qG7xdcUVWO4e+0N9dFqgdfTxk9EfqyrG/r6Nb3KJ1
gqIheDcUV/IyYteaX0Pbd/RdInrV+u1QdqaPe+6brqNcuRwRYKeIMfv1JDa4dysn
kj5McwPKZk2znWqj6wiKcZB+aTmvnaKqWdn++f7i0/SVtQvzTdxm3tlcCMjENGe9
IK6zZasUpmoLZs2HF4zXeKLKHr0q+RljB785obOAzguvrcBNbdN8O/lGmCApS0X8
tRSiN0ZsS5MYI9/9qbAl+IEo9IHUlBJKM9sVahkpa5FXAdL3YdZp7XL7IxVjRhxI
pi2PObDx8jzS/OopkJFUiu5N8m1MhOfKhH6TZioEObZFuFtY7BmX5kcSZHK4o/dH
47+I3QYwRgGlWVqyK2bdlPtX1LxBFn2M/CWt5Y/VaMfnyGjrlH53u16DDBNm+UTp
3glngoLCu9vNPk7SIrDXe3zs3U0aUbhTxg/OBpp/AYBOkdngGpR3p266Nt0/mZar
FEbvY07SrhMm5YH5G0+zbBfHbRuE8BuHpUQ6ZJwEk6wRuUhH1fJz6gcO63iBjq0N
bwgGZA0bLwzmreLDCxrjvRCybrQI71MiLTvh/fixbAbUoFQVPMAk6t6l+7KbV6Of
2cbg6aWmfxWfVgnK3YkZ9rhuSRCwo33kRxNWh5xi8AGGak7oGg932mKK4gVOHlhU
RA7FQnXVlvgnjRrjAjdi0Tzg59FjxsCHq11npsoTL/h1mOILEVr8eBiMQ/8zV1p2
0TwKuci/PWiZY2+4/s0cYZGp7Fzndgch73mQsxHCWOFbo3/lHfSYni+LgoUynANN
8Bt5OAYZIOTtz/yM2sPzRpkm3uAa2F0Chjx8mgK4omjzsb9aSvIySyjf4rUB90Ka
inV1KVpcT5LPxVUkQgZJLchx5ue2kyg7rwa2OyNo2+g=
`pragma protect end_protected
