��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���Ox���0��?T�}�D�yBl98�锛�l	`�ġ	d}�:��PƸ����~��R��o�K�jV�,R����vy���3����O���Z�����g�̼A��v�{�7
��5�¾����B�C����������r}�:ش)qqa���·����BW�4����"V�CL�zhXo�e��6kT]xl(���%lT'�W���'�N�V#�L�`�`�Xy�6$���:��9I��ì=P��uS�I�w��������F��<��s��y�i�u�����ml�G")�O�4����}�,r��𯴢}�鑪 _@�y�Tkt}��8!�JŜ�>9��C �gl���-����{���Z�*� 9�[�B���c�M�͠�+�G�Yy"TGz_'l��2/;��	^F�/	b2�ܕ�Z���./k7iǶ�>��R nS�}O�i|�y��ည��s��KA�O-@��`u�p�1���F��-^���Π٥�w��\'�YL (g
���s�@�9ڬ�!m�L!]�\���� h�u�#<���=�f��ww3
Q�f�%� Q��S���t����fZ�����c��ʡ���әO�qʉwyGP�#��S��"=�n����ƾ"�����-��ߍ�2�AG����[ uݕ0"���e�L�qȀ���9�����g��ʷ����s"Yz��'�`�%�=dr�`6Ϫ*���6���co��W�V�2g_�f�X��m����B���(%"�q2�}ԟ��Y2��cפ�@��K)�`�.���U������b��)�3����wo��?=њƵ�S����?R۱S\'y�*�Y�i����t��7-���=�J:y9��9�8���H<؁h����!������1dEs\�n�!�_Mo�w�Ɲ��}]<¥�wL�Vcn�M���0�
&��?wY�rg�{����0��_��II�L?��KjR;��m%u��Y�Ŏ�-W��
�Y7*�ZU�Z�x>���ds�!w.��G��A	�hJ��ӟw�h������������/��Y��Qz�r{�G�W��m�ޛ�1��O�,I|�����Q�~��=�+ݥ�aQ���|�P��Z`��YYq͙ʠ�E�m"�sH�y�7�U��*(�آ	��5���nrߠ���a��^VS�xG�)~Q4o�М�	���	�ĶP�Z�g�q������{���tz�;T{��U�X�ы��-�1-'Gܶ![~%#Q�h����M�|�" ��K�P�ũ�7�\��إ��eg�l7|��df"?9?.�ĥY��L��zR���hGvsi)Bd�1
��v^���m68+�&�E�A��7�:t1E�3��F���mF�/�=En�9A�c-�#��]/��_Q�֞��A����_�?��Hܧ�l���*��᝾�d`�\"Q�.SG���ö��R\�5S)��m�	F��Jn`ܺj�w�L�����>U|��~3�O��TJ�M��x�:j�&�� v�t�Ǝ�Psϡ�+����D��Hq
���>7�[<r�@�ke�����s'P��Y��:�aki�����5a��x��"����n�ˈ���(_h�d�E����-�|i�K�BG��z;��������뺔��Ё���qĝ��'!�R���+���ў�v:�R�+WM�M?9��
��!Bs���a�k���%B;Ced��v����Tr�U��a�̿����hb��l���~���S���dXFYPԚv����J�>߉��Q,�Q���M۹�E��ug�G����̄}4�k� ��`�t�x�c���H>r��Uh��/��e��,i�'�J�|���/��p��c�֑$Dh��>dC�k�pѰ�Ã�Ԩ�!LА8��o�h�{8�d7��3��|@2�E_o�C������6}���Va�MO�]:5M��}&���+ne���X%��PQ���.3�u�TU��}.T�c���{7��;��v!f�˴���0]ЬD\+�J6}��yʖSgq3)�+I]�x?�K���kj���� 1��4�����3�{�'��vj��\��w�č�_�+^��~!ӊJ��z�P"��xr��K<{��p�0�1ܐ�������C?�u"���q�%��ȅ��E������[��4|E�q��?\ˤ��~	�x(_����-?��~t��^u�{�\�F)��L��љ���0 `7��5i����<�]*-�L� t�b��Vp�ۧimy�e���[J;�k�˪AӈxL�w�����I����R:w�S�R��c�5x!��%�������z��Wl�W
�ܱ� �D9��}�_u"~�T���-Gr|?!�P&�Ӱ�jR�7�� ��W�]���T����ڙ{R7��~cŗ�8c��n��ytfse�Cڋ�P�,=��g-X��^N�y������wC6�P�B���F;,�a���GQ_|��i-�N�Nic��=<9�&_M�� �~��M)�nPXMU_	�zM����`\z�3��O����+���옩pO���C��G�����T՘�a�9�_���ͺˈX�#�PR�FUԓ��N������O���;H�{��o�-��t�P�`�d ֢���'�M�����*LU��#gϖ
WNB�Z/�]��_�µ$�x����/����D�$��'����j!�u���R�� ��K��1ɴ��	c��m�����Q
�`�Rx����FXiյ��Q�v�g0/ztܻ�u���pq�
[�������Q6�T����&0O1�5L��7T֠	�1��Ȯ���FK�5��r��'�\2�e�0dCXa� �^g���^ѓ��G���2Gho_NSG5���A;cOi�̚B�G�����`73��M�,l#02��fЄ'S׎kN�D����o��5��Ϡ�ȩqo\eiT}T���~��t�0�
�?'� 6>n��1�F��k
J���jl$��~Bu/��ޮLX]D�>�u�Y"J0~���OV�F�*pI�oA�b�c�ǉ�+ �Ƽ�Z��2��$:�YEKz$=�R�=��2�ʦ4{���]DDA�~��ׄ�Q�	
�x�"���Lv�v�s����� %^%�WN�*�z��bt诚4��Җg/�y��4�|�s��9s�{)1wrD�]s9T�-K<�k[1�xO��Zn�٭���C^K}��gر�!Ӽ��0W���)�9'�Kz�j�R�<�O�k)�?
��p.-���t�q�
eJ�g��2���Y��tvH�r.�)�����R�&}Mz��_Ƚ�؛���;�5.D�T�#L�Dt�"�ur��jE*���z5��I'I�3����PR˿��rZ��mkM�oVW/��u�B�J�������=
��Q�Y|����43�j�hG1M*	)K���4�l"���Ve��6�."v�û��1ۻJ}]U��z8R���n�R8b�y�n�p��XEY���:^@f^��@B��p	_6����	H�������̿1fK
�ˬ����s��l@	���5�'J�u��/e^ �h��x{a��?_�H��S�iL�e����)�l[^�R~
p�򹡁�e��魃�tJ��L)���;4a�[�]�*��,�5	/�L+������L��I��ZS;�ndtf}��J]S�o�H%�>�i"�	��(J3��k�g�;	܅Vi���Q�����YW_��=���&��B��������Ȏ`���N^�p��?��|sޙ��Û�_�����6Y�aH�wt^���X��-�ؤK���v[�\zU@�����t�o����v����i��a􊛂N,��M	���_�c���&\��lj�PI�3h����01��I?��W��fB�:�Xbҟ��Sc )�M�Aߵ�<��UY'���W ��D"�6�]��_�U��=CǙ{���w����E�G~+L�IV����5�Z��f����E����Ui姲�ӽs�m9T�r|l�`~[������x�S������(�ى���v�y�N���)M�/7*�����8�B6�:;�Rr�R�����@ˬ)�j٠����KzW�π.��u���?����ÖR�1���Sǐ�+@����~\���>[����
R��_�tB��m 	ߪnR_�y��2�i�u��F��i<:]wM�Rb;w�&���Mo�|�htk�)�KmA��&V��P̴A��ai�L*s`(_��_A�v�u�o�qe��i$�� ���H�x"��#@�.� ������V��^v���� ђ�쌌q�ӭ�LS�1���>��
_���׀�	[{�_[�|��ٓK�CO>픝S�{f���^�"��k�v�vp���� ��駓�2K�0>Z�6;M'��[���˝�KX�K5_7j=	�T�DRP�?"�G� |�qn6�� RQ[��з5�k�i��nF=iL�������6#�Y�oS�A��ڠ���o�N�!!�a��fk��P�U%yp'~��-�"ܶ�i��N�ȯ;OQ��#�ћޝǸ�մ\UR~(���6C�WHU�il�� &+���C��I#E�C�u�`A�������a�NF�B.���\sl�k_���rF���7`��Ч0��t��}�a��]��Ү{�8����Ft��=�ɺNY��z���F�j��֢���`��ƍZ��1��cx����
*�Ls�
�&���f�Ϧk�O.�6�"��]��iq�u�Wj�}�E�`���Z0Jg�!{���)1�;�����3k���uZS���?�����/q	�K����~v�_X9��fG�y�Dn��ӟs} ���>R|Z)�+f��(Z����� ^p��^!�U���U��Z��9�K<�<���t�ؽ|�e�Բ9/���)w&E 6l�=�T��P��|����h�4���(e�D����OJ�t���.���'��߉�7c4��a#��� �>p��>=rW,�ާ/��wJ0����b&MТo��Q�'�Q༥���)q%"G�{;9N�$���xGCG7�"R8@<*8�C+l�nN�=���W��@䇡:��p��%2%Ҁ���!�0
/ض���`ؖ��+F�m.��ps

Q(�2�o�l�:�����4���	�4��i`��S��İ��Ɠ�w���vc9�G��SΉ\g����0ɖ�,�/��&ܿ	�[��ލ����6���C4���S�)R��#�K@Bv�8͵V@�/�����:�������<O��0����]5���m����q���d��6����8Y�r�<�����+pw%��Qu��2�'�E�i]�-����1K�ҿy3G�D~Qʉ��o!e�AXP4��P�zUQ�!Q��Z�F,v���g�{�2I�:Z#͘a���,ڿ������E�W��o�e�,��]��3C%�B��j����&�4�^��J(Ym27[���@�?��C��b+�z?��L��e��`�D-j�b�]��_G+v@��C����\qQ:3"�?�~���-@�['-uA�;�����O��v�b)|�a]�p�MGf�� D����w����fA�!�*:�Fw#@!Jk�ѬPX��Y!N'V��b	�]�w@}�'����^sɶ.��2�L�.�Ѹ)�`�|�VOph�>��/���W�b���:��k����9�V/��Z�ž�^���95T_̇y`�@W�F�ޱ��1Ȏ��f�|��˸$%F����Κ&�����
"̠4�"q����x�HJ�2Rs�MMYR��N������U�v}*����bk���3t��C�T�Q�,M��3�w1y�R�#7Ag�'z�H�����Q�[���!��� w��8�XxI�u��[�fO��<�>*�<�7����ױs��c���|���z���eg�^�g��x�]sc�oj�&�	����L���p��P�h��`��4 &��&2�஽R���va�s�S�zv���u����ɜ�B�Q��K!�\���]�Fk"��wn'M��p�P�6�m����`��B$j�F�賹a�%��Ib��VQT܄5o��DE�b3���K?�;Eu)?�ݺۺu/ztyʐ�����Y܎��#^�(�>x��c9�%s����J��	wYK'����� h��"���b�%�-{?�me��I��2�g�D�qp��@ey��]ef��M0�D����������Sx��K��b����DGH����˓�F���R�0d�v���fMKyF���'��2� ���/T$�Ɗ枥���p�K�R�S
��oYjּߵS�%sW�_���!`⤋�%��7ڀ��+^�M�r5+\Xz@����\�$�CkĎ�0���zelSl�0]�w^5�Ź؁w���P2/�J����@��f,Jy�� ����7A!�::�x��ҹU�J���L�l�4�q	b�^}t��2�`�Q��Ea�����`��\�_�h��(�)���U�Rlwz�����1�Vs��ލ��WTs��b���B���ˆ����G�,^tJ���F���_Oz� f�	�HA�J��?�(..���m��)��J^E�����H��%��E0&�b�.^�['�;%O}��D�?�B]9�[��22�)u?����@SZ������όԭ)�W�|�=�L��HdhWyJ3L�$"WUᒹCT ����[?���U��ٿ�b4B�#z��dw~����v����NC찹� ��W1�I:s����|��O��X'o���ā}ԳLE�>�-��!�߅�#;��G�W��b-OU^�f%�g��'r��G |V!�be�� P� 5.�U�b�>�oU�:e�١��`�RZ|����.�L�?H���0P��Κ_��=�QF# �D��j�%@���0�^+ ��!&njހi�H__<�
�7��	-�`���	�q=�b1��1!�n���ze���a�+.K�z�bp�-	��v�W+�R��n�z7����h�Dތ:46���s>��S�;#�ĺ�[��2G{/���~;���.��E�v�/����xS*-�[��/�� y����6�I�����[�0�o���Ր��8���5%rZJC kI���j�	>�x�,�<�$�6BQ�*a?��҆$����KX�����24�H]DNd����9v�ksWV�6-|��I!��]J��*~`��Yn���P��th���F�;������Dm�?0�^&A�4���v��LRHW<�`�gy�`���"&��_T�A�pq�mR	wuo�D{��~����^�a��Z~{g�zO� Vc�V�@���"�7�����9������s�Jyoͳ�5n�ٰ�����8��G�\��Ȯ؞��a)����������l�4��~х|�P�o��!
�2b�� 2��H.g���%�Aت��$�� o:�F���O�$*��HLD������9�((�o;��'X>c�~B&���+)���IEz��0���0��G[ SI�n7"t���A[���Y' ܬ���A�!I���[��K1����a`���A�H*} ���#$dBdU��Q�Nװ!�V��n{�i���n�̖E���a��Ohᣒ�3��i"'u��s�[9Y���4g�{�H@|N.�v���=�$��[��^eaQ|h��*��X�QW)��Q�����P��-�|���p��^qq{X-��k�t��L��(�I�`�l������8, %�����
W:k�+��,H;�j�v�X��->��qH�=����Y��C�`B,M���N���jC�t�v��$���{]��.� j�igJ�q^�Ll�#����t�y�/�T^]��@}gF������3�7�٩�ėJ�9��X\3W�
�UK y��ف�W��}�T�5���s�d=�LPׅ�2�%$k~]2�׻Y�/a�Ld$��7㳽0���{#}������y��H)�>Wnzh{�j�}���;=FL��2�Fa"��?]�G��ԧ�8�Ov,�0Sj�BeaZ��[1
�;��a~�}u4F�jG>~�S;9\8�&6�i\!��+�O)���'��P�?��*I�W���7N�,,���a�R�X�ҳ�Kd�/ʍv�>�GQ=�'�B�6 �_�d{��mJan�����t�I�C�p(�"�g��ԗA[�[~y��mz�מ�P������H0�5���N��ێ� �������$?zg7��Ӈ�3���H;�m���CU��A~}Y�E�"6k��R�
�=�����$q�I�����hQ������iI_�I����ό�@�b��N���-*�4��7��@�`��\���d�M��n�T=������Ƥ�q&Mo��̡FXˇ��B��<Af�ۭ�L��0}"�6����ct+v�ݲC�t؀@bu�q~��9䢦ex]P�T]�cZ��0G��jc�9�8��x\\+�Ei�(�wZ��V%gz��wz�֞*��e����2�'�� �҄����g�'s��9bo �+.�NK;�@.D_�,���i�ކ�ɣ7��������/�����'��c�to�5.��!�����{tO��F��Ÿ��)A�I�!�覰��Lv�x1�i��<�|-����X�P�o�`i"W����nVH@�t������w�������B�$z��ێإq�:���2� ( L��Q#���Y�Z�'��=���1�iµ��0)�Ձ�4΍@�q���{�֨���u������7ʺ5zm�Mo=�"�<�1Z(���ͽ5;�F�++�H��(��	�-������۟=�ƔQ0�~���$j޲�CퟅG9E����Յ��7��nڕ�^��ۯ�i�"UW&�����bk��:�S�/�l��~{֪+N/�-,�Q�h��{dn�V^*(�Vf���1Z�gj��`���μ�q�)
2��$b�eND�'��c��X�Z[��Č��>^��h�kZ�R�l�&B@�n�D��/'����C
���#��Z!�cSv�!��NbQz��wdF��-��IY�5X�a��嵹���k�cz+O>)����d���B�4����4��Tt�V��^?ts��#f�bf�8�U���$1�'����P1�Gv��L=��I��Cs�sT;�3`��J,z7�j�j�b���3L� ��UГ�.Om	����ExG7��v�x��[ܔS:���ߒ���6�Y�o+�c��\���  N*��Eع-p$��O�!�7H�a�P��q�w����va��cG�H���MU��l5��kֆv�].�>�H���cM���s��+�%�q  �	�ܑb�zb�nA\�7���@@� �_�e�jO�G�)�'9L�:��Pue�V#OE+���\ ��/L�FX&�.��w��$��V��a��n�#tE�K3|�7>"~�A�;4TM� W�	S�!���f�� yxf|]�]��s� ��YoX��`�)����k�I��׷�YtHB��Įҵ���J�H����>s�}N#R�/f���nՖ��F)��	3�5��aU�`�=�N�yk�����q֦�����޾�j�mbUd��M% H����!/����1����1R�xRċs� z�I��a�W���F���+����	v��y�;��rwrY�79�K��P
|�3�*��j�y�X�-�
iC�h =����T-ք��{�Ĉ�~��R3n��s3�k���s����j�<��i�r�\����,Q�:��T1V1멤�c��:ӀlQ`H��'�!��u�0!s�[�h'*����'A��M��;!�ٕ���8T���A@�Ig��9 �"���d��粌�*�tO�QE�HPu�>Iv���QJ���W{y<
=�x�b�JG$�r�_<�z�9�){��G�D+��,j�E: �H���O��@��y
se�Uj�$�6E��QBE���1�B�4� �G��p��S�ҁN��c>��h�s�D�v[M(;L�z�Ͱ���|9%�En&��7z��>��U�'��N�g
O�`�������I���=�hg/g����5�\U�>'")e�	\?�R��)��l��4�N�]	�s7R�i�
�Wm�I@��E����9�?V�F���7IX���h; \���L���r�jA.j2�J���-+	�j�yo���K��D�o�C��jkR���E�gŷ��1IV�@���@���~�ч�{[�A��sb�Kx+�/�.�ЂdO
?ɞ�eh�8�����Jü���Z,a�/?G��������w` s��`������)I�������
�@�c�*A� K��M���9��GY�&�y��?CS�Ӈ����V �)�c����a�R��a���CG�ߨ�ǿ��X����"�B�Ï%�]���|�P�n�YXx��f@?�s�o� �ɤ-!&>u���D&r�����rv}:N�/��t	Iڃ޽8���`g�xy�X��U��g�_�E鏹z�drF5�E���| �"�M���l��/����)	����D�Dc[y�4j��K�X�-�-R��l�1�G��0�V��*Tf��lR6u��tQ����?:��,������c�Ŝ>����}sV I�+R�<6	�~���Fz��L��I.1�kn���^�;�]I�g�^Ւ�������������4i
xW�t�o����߂l����k�a��+�5]���<�t${��g:�dw[�U�Ċ~�z#����{�CgY]��'��6��"k-����`��(2�r���EIJ�9K�:�\H�6s�����u�[�;74�r��Tn�GG�(al�������e�%�[�11Eb�)��엃yrB���KJ�z�6�0�W��y<�4�����a(to��(��9�E&�������������(T?�g��D��:��0-PF�e�S:D!��)�v2��HŤGkH��1U2����s�}ZpW�h�$,��Kv7��0��%d�Z���Gd�"a�jQ��o�-���
6ŪǮqu��S����E��`'��9s��+��kb�Ä�l`�f���Ӣ�|�3��#B�1z`۲�dhMn�"�N�7#"���4��75���FW�~��RP�븝��e[{^Pf�t�ᳪ�~ͩ��e�I���m�R/8��i?�I��H��own�b�ש��-ݑ�����YFʝ~��d�g���#q$e���`{  	)at.1ؑɿj����o�t(�I�R��c!|���Y����v"�ZxQ���X����Եդ���;{��*��]�Cd��P*"�\r�D&0-@�I�)m:�a����ZiM��ۡ�E����Q�";(ݢ��I�c�v��e���os��i𡜳h�
��৙��t��3ȹEș�W��1"(�Z6�����	��/B�2;`�|��;��-V��#�����:�͚��pL.��+�F�^O�_�aQ�͋h��/F�5�K��gإ�/����N��4���k>su.J
jwaP��cL\ K���#�D��FA�"<�D�Ϝ���Bp���3�.�4z��#��}ه.b;L n9�y$�s-kp߾�N&���"��~0YuN��(�>�308zm\-����^hc�e��e�ഺ�N�6�ӂ���uj׀���q��Xڙꦱ?��XBEO-�}�)�_[�̃A8x�֦�����'³�	��_�}����c�w���8q]�7p\����'
����w��A�_n`��_w�p>�9=�n�.�[������yOD(���GV�;�dڎ�[}8�S�Tp�[��_��Û#�h�+6�s����
�w��� �
b=�Z���I�n���%�l!�o����1YP ����(W�)ndq�!�������˟�S�t��a�Wa���<����ȴ"I�#*%�+ḍǐ=����MNO� @���6���M�T���Iaw��i��?㞲���xx�$r$�_������r�֒M(�����V`�@�H�OY�ù��������Zr��1Xf�BK��g���G�$�jI�q ��������$ı�L8�jug�i@=���6���V,+c�ue��L����n=1I��K'�nl+��v���