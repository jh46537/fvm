// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:33:00 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OLicKfLTwuUeOibcuJSYHDc2rp/oykYM1621TWyhRNm5ssFS1gTx8o6cNRX5n3XW
5Dpgt+0Q0BYSchbyRyuhqyO+ZQzLWtPJi1xs1bH94B+MEKa8DbE3Tbu/R1LPHlIa
cBGnZ7XdHRBIqlKTQGZC876qexBSnl4qGc2y2MAL9gY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2656)
vgpnbO3g45Kqthqjf88K5pl/69JjpqZIx/Qo6TuqXUb3IVXp0i4GGCtSXTcWpkxk
+MVYQzcG0YBbLLY84m5RdflTItZ084HIKUSqXIFx/G444DTowLtLgMYwl99/6Pqy
y/BubbScyZZqQuXOBE9q9VcbgIalJOXPEj2spM7ARJVkHvF/KbY+4EqZ+REa+aL4
idtlSiicLptl1sCwD88t7tBpDSrj/GiJSOH0zDXxTQEmkQNTwl39ohH6skbX89T1
QWBLCrPoCzVxg4gOT+VN+Mu/GB/N+paEcJuGQLm1xuxk3OjPGjywxlOOvV5I/JA0
FQOSqDubXWZxRwUSBNEq0aQ1A9KCzKikNOInwO3RqSR35eLOotuBNi1nRbmCMVrs
exIOjDGotXYR79JknGGjKAo132ZE2Qj+Wams22qB/G+tTcVd8w+pL17rM0kdbiRf
XP2DA6ZB96WsMvQ1Z95te3lhTaCGEf9FO5MBCmeI1ERnbyMqogXXNkguX9oYrx8L
5eXmvd+8A/v9R4QQurlzySMXGxfH4kB9mURmksWiJzhXZ4q0hsSd8mBdlne98N2f
IdTD+twmLw67e3Zq0y/nM+UCS4Dw7/35oI4Ib0kvYyGuKEbs/Y8uPJeVPkHy5Z2O
93atMYqx1RH5wOG5G23huDS4aqk2YASN9QV7sP+bnvmxBCb0uEqrHjY6+qg/csRh
xblILk7K38V1q5XX9+1OrwwZX8Vm2ep0NubMkV7DpANvibXchE4bUjra21reUsx+
r4kABAU/ZlhZLMfEeK+oU29F7v8JHYBRHTuRQW0uljo5n1jE9Jk7ZDQVcFfgu5PU
C5D8fKuf1kpcXBSTm76eQBZ4foFw5MIjZkiCPpzcp/y2rXwU3+ZhPkJpCmNptKO5
2EvL2bbZePo0kjAF/DFfD0G0YEKH02ltbu5Z6M1EtAzcJdCb9MoDJLOe+26fI9uF
FicjfJQvdakNgFTQQg5jNfnMhtGYW7ENo19vg122NOvjYnIvVJCcNWdNb7UQw5Hy
p0IMLC7Ur+nCp9jBOpfzEm0XBEAqqYt6O3QJcW2w4mXwpQcBE3DYnu1nAj76QrAz
YEIcXTQjowIx6XZAmG3aVVoX8mdUS6oQ7h8qYt+oHuaxZo/2emNTyTbvEOG4H/OU
lnag+JzkQIgZPg2RUCqYS8jPU2qiwHPpiw86auaE3bsMc4tySlnn1ggpKqMW8ADQ
1pf7XsAOm4KzY1fCs6aH+xY0IXYEjnbuEvsp+/cSxzPQgL4apf34Kj7ZgvNa37p4
SaRKBp1g2NLJ+8z5L3zHBMuEcLdrKFAFyLsOgpW0y4pCMTgJVOAsYq4q1YipaxGn
xiW2hy0cXDlAsuT0Oz+6GGlbHjNNDfm3Dzs3cLV6mXNr1vrLQ8dvnloQBHoc4Zob
S0khxGCaY+QP3DshccxVsWfRgQOgS158NplKG7X/w2mdQpbWSLfPx/RdN1DX1FDN
CgcA5/mRQgijdXvO9cjk7FrxeQqnstA46S7HUQp2gQiYLrwsTz32T2hxJB8JHMLQ
ePkqrVvOVf08szDu08M+Z1nnOQrIup7NdTh17SnWyk3GWqqiPaceWP3WUxYISLY6
MT/9wQgwnygULX7ymTh83aDAGqqX6PofXypngD2ZzWpOpWiPHeplKTAwAkm8Yuw9
2cF/N9GmZZ1WRBYnFS21AR8fmG5RO91lnbi7Du/CVYh/Gsr3RGmDHsn/ZBNehK7G
/nxurcJujMVMRk6wEhhiMrPAvNADLggFvIYBxwv4UKKZ+cNPqexcfDUWeNmF9zFX
Y0Ow5/wtQmO67pPiLHYnSLwvQQkXvfhVf+BOvyyolZ/t5H3NtH5z9EY8+cBo8l3k
7ETwN5a5k3S9eqSB/ebrDUg5eONyLr583e5L4NVQql1toXWT2ylJH+1zOQoP+oR4
VyVnQwgIB3/u2W6ale/LO9i3kdVnUXk3knjUrb1CoSONsYLG1VMV9lIoEpNwnfLJ
S6q/BcowZOZjj1DfUPuydzJ7XHeN/nfZv8SffhYSIb/Q3x9FlNXkWYjIfvqsNqVp
fTdxZdGWFYkpWDfCUmcQwUGSetMtowjlBvh79nRV11yIKvX9UzFMPEJcx8IHxlyq
WHS/3IkxCWWTwQrRyTH3gSWzOmGLvjnjvoQxzbaZZSZ+UtMuwfqzANsCfD3vWg8v
EAS2kJPXHWdTy0sO2JA4FyWYjc7j2Yco2xXyq6S61NZ68vXgvRdB0JEFWJXmeDSv
IsLqScq66WofEmJfMj9uaKHNEAW3aaaNN9dZ7d5ptdrocpXKw4PZjLKK9RPP7i8q
WsodP1A0mhDCCR9vXZS5NPcsZPYqkihTcUwG23NDVEKitius1OFA/A2BXLOxIpGf
CkmtIPkqOMbKNR4/VDZ4QoaIUSv9W2KJuu10QQgp3mgTnbF8HJXihVjGptM0wt5+
NUJ52dePeRaCLAPbK0FRTXV2oaOE5aOxEjYdV3uJcsfkipJuMlb0JEzj0ajDiZFo
T605CCTBdzv9UB5AIcvJekvte5fl5ZtvlvqqOMkazRp7TwvBo/taxrorxHlFeioQ
o1ssZReR9cZeP3sCf79IVRJpWLdMqKs+QqzjBhZ3pVd8jDZcBr82J9YzGF2n2n0X
DAHMHiiEXlafUoUrusCVMCGjsKeltlLO9ieN8p1TXXxCxA4352V+N5JWX2iGzv6J
A5RVjQ2/pokjJeaLW7JuNA4NBwbbOu2wEghL1tQ/QHFizBT/qBdtY0fL6xm4Cmst
9vTp4ZIP2ZR9raOH6F3ef5JHL102RgOFQRyqk0LUksdjS/yPMgrhuHY5sGrzsOoD
KmuvoPHlo4jaS9opKc87kbAGGWKLe96IxZXqKoB3ZP831SRLeVnQkEzG0kjARlXU
DomIAmjL9s9SZvUi6pLgL4qBNSpOE987GV9W/h7OxhHwAaRuDG+5auln/Z/Qcx9v
o0/ljxahobmlwUSr8vCeLpbmPNeX5yydHW7TmRmnM9krQrLVFXUCpeGsuqu5z0Yj
8CJyDK6zj1D7bzJVB6wcpdlOX7gjZ+/LECDg4E4Ji/8KRXIBRtkoZ0isWdGxrVqj
oGaBy3cymhgAVy706XeQli1qFFxR0+cpgkCCzFBjR/LDkzBccczRVuwkl4LBov9Z
EoOjdLV237TVgaVYvEnE7kqBOIU/RMifdtDaOvgSIvW1lBc2UuRzqnsjiMWMZ+PJ
Nd4j1Vgsic7oR8FqWP8upng9kNJmjOx7SlbnZ9hxx4Ok3kK5vKpliwnrJD3hd946
Ls2kRDjzciEr2qfJRUqv4/vsZs5An39GV30OrmsL7MvVJ4ucv2EswEFkjcJyBh32
orZw/SAL/FG5FHrYgj6m/er4HS6P47ij8v3rQAItJu58UfQQRUYC6QyCO6a391x4
O9GtAIHrY+pa3TrkHM4vNpE0PG/TztXNXX+JwIecEnGc8g7QcA+GDVWA97mxDHy5
lwib3kdLVh0H2NvI3UmWAxFGQDp5bAWIn9xrsIJGHO2pz0loGiOg8sFgTHS11D8P
aqmLlxkG74UY9xv4EL4vUg==
`pragma protect end_protected
