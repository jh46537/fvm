��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzG&jI�#�aW������r�2"ݽ'=}WῶO��n	`f���UW-�}W�8Vg<V�j�F�HC�,�x�G�n�����q�)� 8������l5޸߮�sh\�N$m��Xkf(����^��f���/1��CS���@������%�l �Ģ����oV�-�	L���E�y�խ#溂Yyą0q���%�M�e<�u�{� �%��ݳ�bʑc����ig��y�(^G�#�lʎ/���Y�/�D�^>�%������LD"��舕�@��&���hs3��ٿ���@k� �Ei5'|� �a��2��i~��X��f��O�M)�{mY����(�����q4��/��#o����-�O���'��Ϫu�H�T�������ENj[�`+l�SԗHbo�P�s4uC��Q���M��T_�O�� *��9��� �[{������:�j]����Uu��"w���Rb�l��6�w�i��Pfpo�?+�:����C��Ӕ�H�Ϥo�]N��ka��P���_����ޟ,�Aǿ�'��L�{�?/AJo@��v�2bɵ!��������@�O�O�X�A=N���g���s`C�ɮ7�h�?d5,��S�l�3�,����m�ɨ��d���Vy���s�8��F���;�-�D�[�z��u�(�@�*���l�&_�n��y>;�=���0��k#��5��$nH+�7�+`��t�bDu��̟O�>M��S�V�������F�/Dd/q{�Px���pM���ꩊ��؄Cq��[p �B���Mti�?�r��F,�
��?ī�ɕV�E��&������2Z��CYf D���n�Y�yj��������j�͍rF��`�Ƃ���h�~��������q�;�(pQ��,������c~*�*�����7�]<�g'�ߐp��9��::��)��՗�P�R���z�!QmTB;G��$�^-�9y�{��`�6��w�
!���F�����M�B;���EP��B+�M&�R*���A�#�JC0W�w�8�cui�egt4�*�����|-,5�ᯝ]���Â?���� �9U��R)�˖�|z?���{����ӄ`��LæT�K�q�c�c����ϊb/�hP�����E���q{��c�
b9y�M�����e�ĀICT6��3���>oĿMiZ��?0<{7�%;h��[� �/L7ʆK�<J3<I��\��'~���=|w�J,�D���Ǹ\D�+��JP�����������6�١WP��8������Ry 0/�'���:���.�dP�&���X�d�����0
Ŝ��j}%�p(�Q
��ƨ�����	��SQ����)�biO~]���P��!�Mw��]-��\��dD��M{
�~��t)~\�S�����u�sk=�>�"��,9f�G�����نLA�����(�u���t����r�E�'d���C���P�=%����/��L���=�6����v�� ��.Jb��o˙�&KN-�$�2�X߷���h�<�c(w��"«���D͎����I��P��ۚ��fI��H��;�fCw�؛��8��f�0,4}*��:F�����Xr"���[����3�4m���|*P����@N���+�Yݙ�tz��$9�q�� o�;eB��.L�;�uU�ef��{���pF��?��ܠ�������*�U����6D��}h6K&H����_�-�u�E��B�䋚.y<
Ѷ-%��m���D�[��e�I<Z�~C�ӆT��n��܄A�8��c����?� �p���_z��v�qVs572�A��8\�����i�"��vF0q� ?���(a�G�v8���_A�{�A���0A�M��sՎr\4��K���C��)7i6D��Y�[W�j����ɒ��Hf��|s&?�G�X3mP?ȏ�V��Q�ܑȷr��J��=HP�bb/����.]}L'�l��+�n�ޝ��E���vw�{�����Ben�]V/S#7��)k[�(��(ؕ����w�b����1lm?P���������Cմd�P��Tu������h�~.�,^��E�l����,V��:��u�<���-��=��Lt�Ԙ5�aGD[$�CvH�דڗ����&ep�V�2:�Q�Ւo�3ߎ�!b�X���;��6|�t�6p���w�z���/��FM.g�jMf���bf�M�����|�=�yN�\��n�6B@����M�*�8�D`& @���l�wW�0�{���o�~�X�+���-l���x>'Nr] ��+��ZV�O7��V+�������tΥf�1!0 ��sz��Dm�)�c�QG�mp�N�J~�X��č|��g��[�JUw�딟.XJ�c�5��*#�)��klh���	Tx �����C�8A7�� �/m[��p�lB�Y1�}J��6���	��,�����>"B�%rᮾRS]�$6��⍰�Ӻ�����_*9c��	�߷����)�A��ҩ�k$k#���5��O��ƫ�@fm��ȳweţoE ��\�F>.wG2�^H�ĝmR!"��ߋ��]�$��N#�-7�X�o��*�#�X�g��Ա-�9�E�3�]���E�����aAd�b��ݶ9��԰�xM�́5Е�ӏd��^yQ2���_(Ig�t����:��̇��vݸj�AjF��ϛ<P����VQr��k�܀��I�O�.*r&>�=���=��md���u4K�ț�:k�}r	cO�D���hڇ=>��NF���O�PX�U�MEC�f߀C��3�efVmM��ݦ����A�.,uK�S�œ+�G��˝.:��Np�n��)lBVA���Xe8w[��m��x}������
��J�^Y�p�-�
	���4��uh`�d��t�N��R	��ݗH����ݳ�)Yw2�KC����*�E��'�J�����A�!��f��Rcu�m|��'"=��m�"
�x��5@Up�^�-���vX��ӕ�#0�,к�m�f렌�N~�B�g���Pٌ��G��H���HЮ�A�c$r>�@��+�~�?v�"��gz�8zg��t�5Ԯ��7% �]��H5�݃�1!QI�5h�3�q[�}>#9��%���7�Pl����K������CC ��5�]YÐ��\.��;"�qk��uM)E�A	eqP��ݯA�6q�g`��#d�H���xs��,]��`_���z���/Ѱ�F��8���.���:וOƟ���|�Z�Sh��L�����A�\s����0$U#z��E���rl����m�a���p���Ձ@����|S�����".y��HP����{E���<*iM�'�H���cx�!d���>��N� ���i�x�9*��<��nY"3=&h����LnUk���	RG���ò��{(�LR
5U9'0�����]��T�^qĴd��Z���Y�~C��8QPI�Vo�8���Qw��@��.�~������-��z�%t���PP}����\r9JRܰ��#p��B.~������� ��0�u.�8$�v���4��>M�OB��+��OlCkn �H��xG�̳ӟ���ǳ��Q�rZ�k���:Я!'t$k������_��:c�F�Bg�E�A���д�Yox�<�S�Sbbns%^�!G��7��O{M���<�X.�ѶK����mF����[�pO9�QGk���D��o	I�|X�s�[?������b���$�@v���-캢���,x�JIYz����ZA"�%YK-�;g4�{}Z��)��ѵ?U]�8}�v��O\?h�q��z�E'�HD
���({�Q���-�	�'f4�|)7��aݵ���x�2����a�L��Ϗ�y�Pϊ@�Ë���cZ9�z�W���έL�hI����;8�Y{����qc��`!|Z��Ұ�,e.�L��ΛZ�i��.:�(�L�)(�C��
��Ύ@�>�^~�kt�Ny���b:�p����~��
kIB�Xc��tT��J����M��
��E녡�2Q����~���r��~���J U�-e��+���4cY\��](Bl�����3�܅�.��P���pT�-'Ɉ^wgY�4}_̎�胔㜏~�4�}��_�gd�s�M�I���c�#^��]���-)t�D�9��$�7��?��b���9`7=Bw^d����>��W"�W�1�����(Na�^P�2w�^�򵡝;�L�fM��.��(�68Y�+�H�S~V\�*� ǉ�/��]pkQ�;���DqYe�����%�v�J"�zjR�6���?j��t����v�E�$�+�H)��U�7 ��\tb�Z�Q;ü�h�p��D+� ޯ�hM��Ge#�����>�������s��@$�ߊR�q�j�[☍%h�}9Qo!�+D۠V���\��ݎ��PQ��ƲĽ���/�(�a�F�8@:XP24 ���.�ۑv\�	s�Q�)b��d
.yX랒(S�ݎ�����FL��E>FzHCo��1��<�}���sy�����u�f9��s��Y��}�-�/���5��Z	�qP�^s�_ ��b�(����D�*r	24w<���{y�Zgw؄���qC������SXn��w{3���5|�O&�|g%6�rJ�ML�c������fee2*��¢��7��җ�y(ϟY\O�p���vץ�W7LO��1�W�������K�����ǈT�ՇM��Ñ�ŏIhF��D�m�����#�� �`v[~3�al�b��yg�2\J{�:�]:�5�ͽ+�,*Q�%K��c�s\��9�O`����JCR�X�HC��j�)lSg�칬it��{���1��%0%�/9�e2o���>��?��,�6�H2��7i�3D;ǘbF�����۹`��]]oF����t Q�v�ȿ�V�0?�����T�	} ���>�����^Ŷ��c��d�֕��7���*,�WՐM������nv����+���،��k&~rn��IP���8U�W�*HVM�c~C�C5o
�+�&�G�
%I��T�7A�-�R&�{,McZ&����#�݀�	��^W���߯�(����-Y��C|��0@8�!�-�j~�F�F�*VC�x>��r0,-N�6��d%��^�
~Xx�yF^
e(�Ğ�g�Xe��-�D�}Ѫ8��..��q4Hy([���<�������o��o��
J�G�Y67�K�jR���nX������1%`�6�v�r�3�g�Bsi6�܏�6��O�3~������V�%�pf�6(Ck)f�|2�s��7�����չ=}���s*ڤ\i�eP]�}�M���7�8��yY�^wMi��V8�B$0Ƞ|=i��9_n�g=N��!h�_)�DƱ8��3R�Ss�ƴՒ�T�Dp\h����7@���	�`㌹�2�u�w*�A���p���[,�1�x��,xk{��kA�`��\O<��d��'�AC���#����a��8�_�L��G�'%�U+�	�8�������l�C,�t��z%Ɖ/r�b���f@������N����}Jh!�R���hm��=���Գ�#'�,9�n:�Fi�'��ϻG/��@4!��k��[O���P��"��CH�T�W@�n����`S�,�C�Yz�Dcߐŝ��1-J�y-���7ϯ����}n<jZmR
����	&�a��澕��GG��j��� ��r�3_*�u�<.-�O���L#u�N���*�G�6�.L�$X����8�2�>D�)���ɚ��L_�H=t:ϥÎ�q4݅�JY'��Ж��\�8%�1�f�:@Za�� Sn�3AKD���r1Y��Ũ�xy���&��o>&��
�
t��j�@���A��6_��O�����ݲ=�H�0����+�s�o�+����.����2G;�a��
¡�N�;�SCh�o�g������#t��2����eњ�Z��J�ĥ��%.t��4�j'�)��`��Yj�0N͸h�E%&��� r8p��e�Eba����µ���%%2�U�p�nqqs�\��TSi<"
���W���9�hH򯪑Z�LL,1z�׸�E����]�� C�X\��P8�c4��X�Hbb��Q�'V��31���D�V���B`CE/�ض9C6���QC�޴";��Ю:�=��Q�h?��g�Ov�>����#��-��ne0j���L�+7O]�?O���N���aY�{����03n���|���E�C{xz-������,�y����&���`P�itӵ�W�$��]��4��Q�(�7���n�Bb�8�Fo�;N=A��G�:���p��KnxPX�gg}��I�Z�_J�.���:��M����Scoڴ{_G�t��� YCo�XS� �}���_�H��N/�6ϫ�}�����3N��t�(-]O�b0��N!�
Ij��A�S��3W�,*ǔG��ZW�m�n��q;�7�C�ɩB�@πx#�����4!����-d�4!�V�R����t,�	0זc*��f�xb+�/�'_H���fap95qnD���ܙ=W�:��
H����~��Ɇ��6�TG��<J�hN����Ο���U��kȋ c5�7��sۭ�{��"�}=;��.L>\<��vX�j����b�mg���knCd����#�$�z�?0ל�a<��w�x(O�h>���J4�Y}k�ؠ����_;5X���M�fPß���͂=���-�6UJ� ��'�SB������>������;D�B�ԁ��\�$��{k��R�@r�rA��N�����\=�{��h��jè	�kM������Ѧu[H2�ӆ9��}��Y��f�{�#0�-ӟ�X��L'e�>1)\/����b_NeaG�B��#�T�wpm0W?�,}�L�!ܰp ]�`2Â�i)ߎ��r)�O�SaC�D�6]��٬�M���)�G���D��v�+���)�A�7�l�Y�kW�.$|��L�V˒9�z���'{��[�شǬI����,%��2�e�&K�P�0nGq���%�f�NSh��&#6?[����I���L��G�\�̩u��	�<���;䤞0I��=��Z
�9�vJd����M�[?�a��x����f���`�JƳ��7۹y���R{tF� �t��� c�e�ޯi��AG�<��L�� ���{M��P"��2�D� �IP��q)'#�*Y��eao�^f!ɛ�i����VX���=O����W����	�۟�7-��ǿ+ ĖI)3�ȡl��K���J��z��"~)����8�,��u�Dy{4�wr~�M�<!����y�ӷ1BG�V+=����Np�L�rg9���e���+n�K��ACB�@ l�%�n�Q/����.�:��i��3:0u����h�Qx��(���Odg�|8�^�ӻ;����ή�UJj&O��p�1�� ��]��GQo#N��C�e�a��N���L�-n`B����s+�"I���)����嗖���W��̻z'<��eEU�u�?�����O�8]���|c�kc���/R`�:ԥW�����J�A'��y�\�r�a�TO��C����Ըv��۲Ϲ@׃ uj�����ܸ�[y�yҍRB�q2lU��K��D�,��i�f�[���RG����v����Hw�����>V�`S��6'1���ߧ�z ���2��/t+��ˉ�	\����P����W*YA4���r�Lh�����f�J/Yo�>~o�ᬺv>{�C�|$ԓ�hk(
}J*� p�}������H�%~1Ѿ�:��f���BgI�Ģ����xl\�x� ����G�r~h�>�B�z��%s��(�C���
	&��<��8a�ϧp��W����=��=���+JWɓ�p�+%СVed���BQ0�L�KY5��-��DX�JQ�P��~X���<@�Y~MXG;緡�9p�,�b��L�k�9��,�K:PE�Kv�3���A�G6�I��K�Ĵ�:���Rͩ^�;��,W+x