��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����p�0�F���)�ã~d�:����f=�n����l�@>O�Њ�۸"�#~����f����S��UT���������בJ���\/��2����r�X����`Ir�K_�x6YV����(�/�~�k�q}����;)���3~�=�FgBBKO.��}�@��z���̥x�6;���X<�����~2�M�2��$)�sFaa��4����9Q@���e:TWrt���z6c)�<�~q\M6�'����/ q	-��# � � ?!3�m���{�D@� �+P>�e�<>��]zF0�P}��N�в\� �Jy�Ǚ�j�qAw�IX�Q�2�6�o7�O�7w<S��H���y7
W��w�Ӯ�T��Qg�"D��^�U�L��u~I=�5U�$��n5p�V����B�E"i��z�MPBo�,{�օ9����Ka��s\�^�d�h{ѻ&o��ÐY��~	F�C������.O�8'��Z�Z��z��|PkT�� �O�Jr7n�p��J}����3����&�L�{[]�B���Qn��%jZ:�,\)���Б����X��%�|c� �^���UO�h�"��L��:���Q�\�9�hK�[�3�Xw���쪍���9�F���nFXT���F����ܮOBi��}~3P�F��*�z�[Y3,m�f9�DQ�����#��Jn�	��c�H}6j�� ˧Q�f���ٛC����^fh|���1�]�
'Ϲ�p��@��f!'|�� �
e4�T��.Jm��믭E����F��! l�^M�~lx6-����0��Z���9�;�E�c��qH[[d+�)��I5Ђ4��.~��+Y@+w"�=�9c

�X�2D)|��#Ӥ^EnI�_s/�
0�I����2�w��N��x�\��HK����e�g�l�Jjn%8��g �(A`�j��6�������Bu�郲	6G�Y�jɑ~jNp��0\^���'\����&�����b9�5p�~�N��i���V�a7@��9T�`�8������o��_�f��GB)�<��V����0���Ix�����G�}��*������W���Nc�)<��4v����;pLC���w~�v����	$2�ױ]���\[�`���"�V�#T�˔D��f��3Y��h� '��37c��x�$3�?��y��x�F
� �^�sfj�]gyp�t�V��lT �7�ef7��0} �&��V`W~�7e�o'$�
x��s�@���>EQ�ε!�s��rm�-Fs�]�w@	�o���YS=PR6:��32�A��l^$�OI�F�T-���U����������T.�O��C���%m�{o�c_��������kӂ��řZ�h�/��D����ҒT�Ff�U�W��\�3�_�s�����+�𲮏f�����4��<^�0���.���[�����F��Z���.��exG�M{�j�;�hm=��f�-W�2�&RR���k�w�CQ=���#%솇;��<C�h9��l�����z��>BY
X(6�p"�
7������q�հ���۠�G
^M�\0�T؉1���E;^m�2ua���L�cP�8W�h!9O@uhB�I6λ��� ^��~Fa@�ZR���H4�Wr���`����NB���w�k>��N �1��{��4VqwU/!��}��/����H��?/�$7QkG�ib8�b��ͽ�Xfk��nw���=���%�~d8���ժ��š���l�w�˦� $6ئtJ�Cl�K��T����܎K�M����p�li)��6��7G�*Z�uZ�H��_|����)�xQaN� ��Y�F����$�[c�2ԈJ�RJ���N<� ,
��$��*�M8[�#��u5��b�����H� ^�I�3Vࢨ*�w�.B��E���	��ئ��o!mY�Љ�bZ1����",o��&;��.N���r��&{{N;�J��@ջ]�5�U�󦓮c�����:��R�
K�������u�V��u�R��bB����\S a���X�8u i0%���^en%������Lwst;�*�&L[�y��羀Q�i���H�IƘ :O:w~�P����.��I��1js~������k�� �&�8\R���%���8rǆ�8�S&��!�yȵvo��s4cx�vi�8�W�6;� >�T�!>��������5_�e5i+f�����a���~��������y��x�ï<�n��GZ��K��!��`��3p4���o��ܴ���<��`5�z*��.W���pH��s��3��uu\�D�j�:�P.{g�bL4�ag��I�O�-%� �0Z�Ê��Ę����8O7��k�1�-"�V�H�x��{$��g��o��s��.��r�ޏ¾�9�ɷe��[���s$m�ͨ*<c��ؙp��Ơ\��g�ޣ�t8Pg�4�]|f&� b��杲��zr-GA���ݜ��-̲�r�9R�
���U6���<]�$�)�D~Nv�9}��)�Ck�v�Z�o�ߑ����K�w8|��%?(�PT �mdV�p,��wƉȕjQC"A���T��9[}JN�
�ۛ7mGd7��8b�~���{�  �w����7��{�S�.R�~2,6)c
���ʐ�XZ��j�jU� �>�!����=�0r���$qs[ʔ��V�,�]E�H�	|�>H!��|p���4��א�ᡍ¶����ޖ%|��<��0ۭ�F�-��nY�(�R�k�d�Y�yT�N�rу������;�;�L9w��o�nU�n��ߝxYe��G���j!��?��X�5�Ffn�S���]�a�ؑ#	���%pČ���T=���S��m(�$Bc�u{�c!�� +�,�P�&=�>މP�s�8[ ���į�R�����a��@bz���,k
+�1�K��y����"��S ��v	�Y%��Y<��O�����&��Xel�lҿ���r��.R6��S�aG�N>��4<�.��4`�H�*�����xO��7Y����Fc2l�d���gm.^!����҉�l��U��ᛘƾ{�;	"��h�O*A�ϥ4�	��9����z����!=�9��\� .~;���zE������9`���M�_���P��糝t���/������~7R�r����3���"��i����b`��f_���4��=g�dCF�k�le����FP�@X/�}�"8=�D4H�?T�>�'(g+ feڲ�`�j�V��*^aa�X��찰�K�!��\��H�v4v�1���5��+L_'{���dR��Y���r�U�������ӈ���o�.��)�e�l/f�@ J�3.����rOW����@�̜�}��D�{�ڝ��ŧ�A,Nd4�gİ/x(����2�p�Q��'��A�&4�v���{��vީd�;2!vE��ϝ���w~̭�&�Y�]aN_����iw��.�AHT`	���m][k;{4X/G�.� ��2�`���1"ȰA�\[�~|��>7^f��0	d��$�I+E�UQ3���U�иU�H1���V6��JK�oqj�nL.��@3����u2���!N���~�(je����ۣ�.?���ϼ����j�̦�;��pk��~�m��g��Loy_�� �Ipg�_�0kug�����sN^ е*�Ķ� jG��?�F-�&}{��$�x�4j��:Z�4��?}�8�l8�D�I���)	"{��t�@d�U3�FRX�
guF�J���7dwۉ\�Z!��"�F��٩�N��z���q�޽������Zw ��7�t� :�H�7�J�`�����۩\<5�H��ά�������� ѷcN7�~8~*� SF�Y��c��-(-�L1,�.q�����@q'>"�<�N�w`Һ���6'M�Ĭ�o�8fi�B��&%��O�y�9@��u����^`�d=�gmJ_�W��Ύ~z
����,��(_�ch��=����+�Өڪ����E�X����'I�4���Q._*�4�L-!Ro�����H3ny}z��	�$z�6 �CF��u�Hod5"F��2a�i��T��k��s��{�p���綉������$ q;����[���|�<�`�멢��i*o�<ݭ�z�����p�L-w�sD�sk�|�Up�sU��<C33��1�a��4�RH�U��ϊ��_�%���RM #�Z��B
�'����[��v4�����MEQ�j+6��62���/�]h4����l��c��~���O'��,XK�F0l��dM d،���0��Xq�;���>i�e�������ΰ�xǫ��{˿	��Մ��.N�sc;j��[ЊF���q }��\���S�Aҋ}�H.��0o�$���⯯���I���n�ZG��F�E��YEaԐ��}��"*]w�&zo��A>���%�H���f��} �?V8q4�>�qA*>M��;1".�$�E����UH�I�Ae6$�wY) 4�����ؤS�wyO�P��-��,~�*�'�:�a���V�5,G�a��޿��y�
7����i����O^�7Jn��h���)�N���Y��Á���q�ք���k؁��5�XYg� ܕ�d�#��1X!Da���Շ�<�d���,Aj\�Q�g2P� ���E�܅�i��7�/�����������&��g ���'�|��td�.��lK;a^����l�ڷ{��uH�����U8�5I�������&<���d��޸��myq���oA�c�4����l��'�h��u�зԟg��c���F%kf�d"q5�.6"�t����y���<�s�¡�>�o�3�k����֍Oa�.�U�@��k���w�` ���ʲj ����4���:�騾�ଧ���-Po��>�,�_���wĳ��听��l�b5{Ysl���k'v��ʟO�oo�6ܟU����oȾ�h��S�/�ʻ#�3Z}Wvx���F����;�{�����O���l���J�Q���7��J-���H���+�=Ĉ"�h���$O��º--�rav	�?s�#��&O���|�7�QGF����%DV���t�]��څ|���X0��
����/*��2����O�#�
 ���C����V]!a���Ps�V;��DZ뒗�hS ?O���4I���Jͳ���Q%]�~,k�f���fC�G�/�ӺC��g� �J[h��3��Ѧ�R�NKgκa{�ZR������*��a�Uu�|�P,:��T�K���a��:&9�=+@l��Ri5���QtU\�wO-�ړ��I}�mK>~	�e�t��[���`u�,W8��C���"����� _� ᧂR�`��q:.�Kb
���P,k���!i���ܤ�o�>#�*J�i`i4��Kۚ��� �fhOB�Jw��L�J��L���E>e��Uj�y��F�:0B��ץ�ۃܞ��$r�L���{���Cw)����MUfZi�k�ӯֱ���$�z�oQ���V������q��m��]���H����� �B:��+���\�;�
�U0+��ڛI�Y��)�½��ID�:���@w��<r�7��
;	�[���������}���ez�HQ���P:�Ԏ�0��ɲ�-Ǻ/��6��5p���H���OD�(�ɌJ��6���,�a�N �4�����)��^_�P'���YX9�SJَ�m�����q�|�@{<��Q�)�������&b�S��9�q�����r��2�"z�~	�18y��@-��?�+�Y���Rn�͏�ܜ����k_��a�련y�{���U/84*5�� 3��_��,�0B*$��v�r�K��Hz�?�I���nA��	;Z���E֗�]�9_-�ԈJ�A@�62�S�޹�_�g��4�
��H�)�j�<w��7N�gI���r�fsh� MĎ�ݷ)T\F������~�9^����#A=S?7;�W�-,mr��mNY�`���-�yn�Z�����`����D���ƣ�R�^�6_YZ�Qy�w��"�b��7`���D�i���?{ã���~�N5i����;���7�qF&�F�9N/@j�TK��;)�u��L�א�R�f�Di#P��uQэK?0gI�\fM�<3�@����)꾴�;K��<��T,�
�aǅ��ڗ�hD��!|�xuqT�����DE�Mt����f7��;�&dx�l��u�$��ca���B�y�m(���^�-�r�/j��q�@�^�r�.���������έjM�`,P=ܢmzH�V�?�;P�o��ou~lW�֌la1�v�~��F�3�W`�!���f7n<������(��?��ƥ��M��W(�N��Fw+�M#�-�Z&X	��z+�vӞ���	�8����[�:�U��Y�Td�xUJ �Rl��|4Z\����H��y���.|����spa0O���!�<p�!y�Znm�3�!���bn�~�;���R�����5�[��\��B�?�*�<��`�.(�$Ą&�|˶Ͳ�`��i@1�[�!p�}+�;�s�-�J����u��US3�g%jc�h��%i��
*.�^�s��k2(�-�Z���_��"m����D`�cB�P[�6
&�l�׹I�Tl��'&����;����E)�Q ?h�Лg�Nl[0
H��:� �%���6(�N��;.�Q��Rp���k���V�Oἕ]�F.�x5t(G̪���������ֺ=����^}P/?r8��I$N�����Ն�5}^:BNR�Q��f�V�[��B|:�XJ�[�s�Iot���cM{>��;�8>~�m�����H�z:]D�hR���^�����IU��g�H4 �ښ�u	�>Z6����E�'i�73PeĐ	�P�9�J��|RN[J����=Cɜ37ޙ�8���P���B��

y
H��"��mܶ���� ����h�?�wR�v>��Y�=@�բ���^9�w�	�6m�Z)xF�V��ct���/�n� ��Qt9,����Q�ay��k�{����7g���GL��x���䑗�2T����GP�uY|�\P��c^?�K�>6���5��_�*�Djv	
��=d��bSnkXͯ�u�{��&���H�+m��0�>/ǜ�F{��4c�8 �}h#�U������MѴ�W��~gy�9>K3&����E�PG�6�ɡK: �Q�㡘(~��e�;uA>��ʜL�O��նR��E)���oa���M��dj��Xw��9y0C�&xS]O/�����f" t4���]?o,w�V�<n����h�LA���rf�;�'���N��`v���5��Iq
�0��s�6G�1	�p�	���ȧ#��f�XFÇ������z�Á�)g^�x�^5+z{������ũ;��-�r�v+�N�-yU���O��_m1��2ć��@�B�����X��=q�T��̦��-��t ��J���x�q�4b�v-j��~[R�QM
��U7���.A}tZ��*]p���?kNM��|^�2�� W6?����9ֱn2��]F�OB'P������5��� �Y��*�lB�.���<���%M4xں����j�7x޼ce0�)Sh��<���Q�\]����\8�!�3��k&b��E���C���{ڭϩ��D�W7V�"<�k�n�D�=��	_O���0]ɣ!b����}9-��p��n�ĬIDx&_=c�JڳsFl���a{��,���OYȅ����
R�,"�=<����Ξ�M�g��_a�T���,�0]X3��8�E��<0�Ie�+,������ڕ7���B�@P���9�K�\3h�o4�����|��K�U���>^W��t����z�\�BB�u9����Ud��Ѽr�r��� | �M��cT{���f�WR{$T*�3\��$[;�)�&,Y:�G,>	E�.��3#9��ޝ'+�v<\�I�lGi���0�����C��K��א� 1�D�>�Y�|�����D�0�yy�Ke����F+�	wN`	r]DL`TT|�:�(I?*2�6�u	��ӧ���ӊ���?�i�����^���H��K$��Mߍ��	��D$7ğ�ZS@�W�]��Q+�P�p���BBk�}pM�D�E�ehR���b���3A�Pdƺ�a5���A��7�)�O��ckAdG����f�
�:#���ד4�d
 �;B-N�5wu-6z�R����L�\LJ��G7F.���h�go7hV��>W X8��	N�Q���`8��&����Vôŗ�� op�yr{@K[Nݘ	��5�t��'��r�q���СqU����|�!��㦻+���n�u�;5��Π�`��E����T�~O�}A������'w��#�0�zK^�[۵�i����Iyq�y|6�y4�u�5�����si=�m+�%!P���v�/=`y���_�h����·���q��j��L��/�)�g�_�IE%43Z�Djڻ�jSuC+J S��"���{��E9����c{+.s��b����_G$��m�i��� i~2\]W�-��1��4j�bK�)I���Yx�+ψAީń�6]�Ath�g�fx^ȴ���4�d�����z-J�־��){Y�^�>�v}��fG�T�K=��^(�jQhM����eʶ���|<�K=)4���@�ar�8��)��\&�/��e y^"|�U��ڀ�Vm"��՘��4�!z-�}��Tf�摧��5�����N56}�i����m_�DD�DL>}T܍�����Bm�aj6�C$�N����}�%��&�7~e�i��<�=�#Q�^(��o��_%_��
�<����L2H {)]�	��ҶW�f�y�<ʯ��P�i�����n����i���>w��+�⭖�I�/\��DڣP�h|`vj� ��j�۞��B�w���T�d�n�`�m^���t��	x�7�"�ވ|�*��:*�Sf�F�ݰO!��?\|�ԁ� �L}i�g�N9��R��� �}xc°��z��]�J��d/�;Df�d-�3�����
0ht*6J8��U��<�nf�ɧZ��H��O�$.�%��x��D�&�S�s��[U�񲗅")\��=���{�2�!�,f�n1K�r*c(���K7����B��YS�2i+4p� ���kL2\f7�;�ezSs�_�y��q������RJ�� "�{1O�
Ś�c8�K'����."
|h�}_0�"%�fL�˸��īw���TFc�
I�K��C��>P�ro1	6%���Z��hna��/��c��i���s$���9Cɳ[pHI�v�_���uV�">!Qm7��>0�@�R�W5͚}�����u#X��%�^�E,�9d�h�Ԃ���;ػ�󂙆�2y=���NB�S*�n"�D!/R��E�f�K���2���)�¶[)�t������*�@h�Pd�*��al0;�Ƈ�<]���R�S�]����V���_@�^��Ri@��Fɞ��%o����/�\��=9�E��3�8�}v�("h?�w���N3�Y&c'��,ܯ�/����M��6���i6�pŃ���.�/hz��K�`4'#����U�Iҋ�*���e��x�]�𭋘c���M��%�	�"D�-'d,'b�uE�P+�b�sIt.�6��bu`�X(D����(�:���~����� ��G�Cz5W��	�2��펚o7��I&����7:�ƴհ(&�$�ǈ�ъt�
<=�ۛ�҅Ŝ/R9��}B�cR�-���o8c>��<�H���m��fӒ3��yv�W�׈ڨd��کR����{/����$깘%�$c��¼���,������j��N �el@8A�H�����O���M�8����j"�
���V�L2n�^��K�H�h�/뎀p�!��,UaX�a�e'�Xo���U�<�w��n'(v|8��4
Rb�P21���wu]k��h�~R`�\�Y��y�0�3"w�Ta"�f�=.��Up#��<Ĭ�n'�;�0�	V�͍���2p8�k�����[��N
lo	8��|�`k�k�^d/ jj�u�$)�No�ǘ1~��u���
�~��S�A���E����M�;1�'A����`��0H(�4Ү; �	�������%_�A��̪E�»�����QƽM���`C#���P3�jd8|�b��7��z�]�E�_��o���0m�I��s�T_��*��	3;6��?#��J|ИB�ꄖ�)9��b�"�>�(���D�?��˶����r��5O��=2��-��jO�@����"�5��?K���d���C�{z�K�.�i!@���a,@�,��Tw��{�����E:�[�}�(�̫�֝	���a
�*�j����&W7(9�dy���������4�iX����v1^&�8��k:�fg�޳��"�s��C{�y���/�y��V��?��,�(7�zz�z�|Z��Y�iR�^�c��TH�#*�����Id%��A�{,�N	���R�@��o1��rE�=��WXy��Tl�]o)q�0��)��c�26�B��։{���MlxoPA*6�܋�؜y`���;"�$�P���A���j�@u�ԣ�m�zCI���!���",��̛m�z|� ���Ǫ����ðrQ�iH�Ż�?�Ewё�%�M�EɅ�C�6ȕ�1��
f�&&��[XSlL߉����8;�MR9-��ln7����`8d�|�	4��*�'�1η�:0f[BOv�y^S����
I�K��6v �'�#)T z��G��+�[�O��E Q([����U����xI��	�d�>�ų�X9�g���o�0���X)LE�a��$�b�;*�l�Q#@&l��@4׵�%)���б��{a�g].gv�4��TU��z����/�ي��{�%��³����[�3��ӓ��ED�;&�2g����{�10x��2�|n���N��= l���W2 �e���w?'	���
V[3uƅ|�u{ο��� >eP�q�v0�c�7�JD�(��ΧG�s;��	x T>0fv���e���%�@�c'*�+�c���Y�۪6IC+|�UU���S�m=ӳy���`�>!-k�\w��+Q>�[n�@��9��~���i|6{v��]��	���-��%��b�^m'w���/m��)��9v�+�@�-Fd�[lT�����r��&��*� �����et^9D~��k{�!?����G��1��B��hF