��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&&l3[�ɀ��t��*�Q]	�5��D޳,�+��YXQ�i&C�K')�-��Ev�\�Xg;����H�	1�,%�E��pM�ţ�n4;{0}�X��l1�
�#�]�m��u�;�9�p�cL�B�!pV���>z�L[�u"� �.��*oѨn0`,U@Qπ��@�u�W�)>H�U
n}҄%�;Be�2��o���y)���[��iVLtre�N�8��n�;����3�GC� ����<���kȟf�¬�[Ml��`�K�eૣ��R�QTU�!�	һ0����=�ג`�=��Ç��Q�![��>����[x�Iq��$GD'ݡ�n\�L��F��AQ��ֳ��g��uh�����'�k0�_,[:�b�M���C-I� M�R�>�W7��?_x�h��H�w�'�����&ʪ�k��A��0�	��f@j++��ȶ͗@�L!��4B��]Y*L��l���	��]�1Gӈ��o�6U!z���Y��N��p��=����Հ��l$N�QAr|2���%��=��� s��-bW�%�󲢡��a�L�$�����M��uf��?D��Q��s��_��E ��(D��LwN`��Nӕ&7��&Z&�'�ܨ�$� �Y�)�G22�&D�x�Y���_�gÜv'�9YN��F�e}[�H��P�Q�i��jP��%��;~CL��}q�2'm%$��߅�q��ٷ$W!*>(C�:.����wE��p��$/]'�딛!6�4(]I� �2���?���J�!��4�PˏՂ&WV8v�)`Y�G�xHd[V��5p>ƶ�~����^��<j�w[��0�)~M-}4z����
������P!l�@(�����}���M�e�4V���̼�����+>''|�呠�kۼ9�Q��A:ε�LU�S� �3�TD�{A`�tl�����n(X.#�A��,��ñ�-�	"�~76Y"G@�R�����utH
��Y�Ě		������ԗ�d�'���ftE��R0�_{{����vm��-�l��-��7/ǿ�z��M?�=�7L�~�6���&��k��_
aw���)kQ�@׃:y�Q�`yKH5�]���n\�|~��F����C�@�yJ?kg,g��BYi�Z�����X�R,�W���@�����Y�D���C�@bO5�du�4�6	yG@ܛ��h>�T�P�=���'W��6>�A�(~�
`//8>&�?ؚ,;��$Z��C|�͏rVJ:�'[7Ѱ��;����	Ȑ@�X�2�+��5h�	d�[���dbD$�L](����[��k�c���?�j	��L8�V��C�W���
x5��Q�����WYߐ$�I1���d�(EjǬ{='t��۫�;�����=s7"�������o�s�8�.7��m��v3�oo|cŢ\H+lcK���I-��b�@I���\F�
��,b�WIj38�48INt�U�5���g�"|<�\�L�*���e���iC�k��z_�9K>��R4G����:r�n���U�OPߗ����������A�Į�%��G�	�I��۞�)��[���gX��qh)&�A��ﺻ�]���tE�`]�}K������B�]byo�l�.+rjr�Cť��@��_�s��f9S9#QM'2	6�N���b�i���WW�2�	j��_s[�����#UO���Q�X��bN} �?|�f���(��U�Z6߇{l/�t���6;�gfъ ;� �
��'�J��G��Td-=��zQ������G�r��4B#^p�7I�Z�{���^f;3XB�I�����S�,Y�>w*6���cg����јV|u���.1H���ܓ'���Z5�{e�F�����,]1��k
�A"�YԌ0\B,�����i�8�g��΄o����S`� ���Bۙ�D���z!aUk�c�V6�f�HI]bp�=>�#���  �XeGG!X W��Ϩ�$�':���?�?DG�N\I2R��7���7������*zu˱m��M��^�i������<�8/ݟ��6�P�W�/�ٴ��Y7F,�ڃʔt� �s�zb[?��ݻ�0�u���,	z��@L�G�x�צ�����̓�Ni�R�j�ŦL.��{�CG��g!{e"���l� ����]Q��
]�MX�>����s��L1P��*� 2.p��Z�-8�u��T�<���n�(ǝlZ��t搏�����j���8�	�zk(j���T��#������jn�o	���N����8�[����2���hT��^wz��h<����޶�#d�&�a�� ��ם��c��}V퍛:�����T�(�(x��`!�r��� ����}@Y���F��<JM<|�{b�Bs�*w����G+EOz��>��_��N�ԌP���z�+�j=(�� ��lvG���%i?O/r����f����	H���TKۤ X����g�,٬��m��)��7���3ve���4�p`���#|�K4Z�n=GOQ�X��mS}Ar_����f��Nǒ�#j]�K#�ݴEbp5V����O�&(gaG�Dͯ�t��cO�r��U���`�ȍ��k~�I��KEI]�DߪB�/ƅ��p�*c�`'�y8��c7�����.	��MUt'�J�?��{�9�`�rz.���w�q�
p�R���Js^K�eN�gL*�	iOP�DB���6SV���EI��Ķy�m��%tn}'G�N�����kAcd��6b ɩ����J���*�Áv:Ћ��?5��9�	���2I�Ph�QS�'� "t�6V��D.����������Xq@>Z��?�K���{C��:|�"aA�D�B��!��p!z>�&��m�������<RLD=l2�R��&n@K���?��Rힳ�J��!�� G�-�:̩-����9��iEDK3�j����������]�d����U�5Ｊ������a��	F���\�/+��^�XtZ�����u2�����yK`�]�	��"7^�+Lu��~�;��3f&��z���}�V�(�/�����SЏ���� ��X�iH�d�w�0�1>`Mh:���SaGlzx����<p�����߫�3�Ӎ�R����&$����ރgU���i�T�f;7�:v/����3*:ʎ>����� �%ށ��֢�C-�2F�ku���5��{�u��@��+�4��D�14�f�dԕ��-^�`�h�I0D)�f�3���Dy���� 4�ƎпԷ��mâz1��^��}R:H-8����NT7���Gu<'�d��9���Q��F�M��Fj��U�JQ�k�
�.��ȬsEj��[��)�Wq���܏w�q_�6��I�D�B� ����\Ӭ��D1�_�~�����8���4֟o+��(��PG���Ɇ�T�87�	��N#*v��NFs����ʫ�r�@q�"��>�﷉�%䮖�5�I�F�O��M~ke����a@`t���.^�%�<k4g���6Z���n7�����p�&�}���N6���ќ�;Q����'ǻ�s�Lu�1�4yD9�y���_�g���=�����R���M�&*L�Q;��WVn K���}bj�%@�������zB�o��x������Qs�C�~��X:��t;�x�#��z2O�#V����;������cD���S����&t#���Cl�,�k����K̿z[3,��h�Wλ�:�����%&���҆�@�l�Ĵ]�7�	�!Vݷ}�f�'����c������^Ir��inwoC*�y��>$��s�;���Q,Gd�+�Q1�1u���3.,w ?�6*	�+k�WG8�>��8�3&�-,�̲w~'L
��I"�X���td���re����Q{�Z�Q�W�~��� ���>�����Z�OP���=�((@���ʻ���֏�)����o")�M�0M�,i�F�Δ=�ۼ��!��B�&}v�j�-jH<e;�o���܇o,��A|�6e�!������^o��A���My��{u��L��%�Hv!N7R�s��0,���"8�/O�X.?ʊk��]H>��K����z�8ԧ�=�k�>���G6�m�p��xj�W�Bg"�nh/�����͚jπ����α�A-��8]_1�wՓ�]��ܼ�]<���d쮋�� ��7��Up���)i�.*�N�ϵ���)�b@3u[�E��E|Fs]\�|m�V�����+�#���M/	�Y	8��8O��OlYJ&�ᴿ�.E�Z2>�p_��q��[�`��Yğ��&(4�����>(�*5��/8�$�,?�韓F� k��L�:3n7r'��N��Z�"��V�pٛ|���Bd녈$�(J�f�%��'��^|��SM�-Jw�ے�2��/���{���L���͚�2�bZ�w���X>4'�W����pV��"��>�hO����2�~果W�� �|`W#92��Z8��&�F�H�3C������QZ�9�'�tK�� (Hn6����Y>uځ�;"׹Z����:��j�ބ��k�̽q(+�l�)���ͱ�r�+ ��G���^k�U���C)�b���V��ƮA���c��A>���}I�H���\���tw�QVle��۸�W��U]���9ȇ�n	�SטE���]&���X�Kdb�AiDv�f��ᝉ�ݥ�
�:;�f0p���>Nq�.�×�τ���ޱ2e]�	9E��&)\0�H����J���H��"�߂�[tZ��8�i3��F��pIl�2eJeJ��E����j��
(��B;'��z?����m�r�
�b�7!� s�r8�i���k��_fz<�#�]NE8� 7�+�`�������S���r�v�s)�Ii[=�X�[��S��ܹV"�n����C���^�j���mƄ:C0�w�P۸Q�+y:�rmSO�8>�H��'��H�'������/��mw|��ͨ��� ��ڰts�k���~\]l0�V�T%��N�2e�mB˨���f,/��b�+���*�����@^p�_�H��_�F0��v��y�ф���|^G�΃5^���0�(z8O#�:q�<�E�c	h~O0NZ�/��I�Pl�\��q�< ,��Dl�f|m`jX�5��&��b?4�+|m�d8*����p��	�:��b�t�ӟ&�-�!����4���靏�ȼ��;�s���;دθ�s����:Ԕ-q�@#�|7T|Qs�Lo�M�� u����u���(Y�Is���Ђ�=~�+ق	i�v��ݬÙz:gb�I�P4�VkvG^�N���>i�c-5��5�vP I��:�+f���!I�Ln ��"���\�j���2w7;F����3�<�6�����t!� p��n﨟"�������+�Ѳ��5*(F�3g��f�iB[5Ii~��Γ�[�eb��җ=K	�g��M������(�Q1v�Qb�~(�X�1`��ꦰ7{�/�͊�DlF�Ki�9��QR��k89���}ë��=Q9R��P���,�j`���(��4�q�Gd^CJ�S�F��P�ș(p��YiʜP�Ԕ�u#�;�� ��f��L@`�����%�)�ٶ��+�;#k��H~�M�oUd~�� k��mX|��3R;3KcM�5���0F$F�<�1�{�%k2�+JU5�1�����b�ŬM�6~B.�_fۋ�?cF8}��N�.+"ܭ���ϋW�9��Y`N�M��{{+㨓�B�x2�^D�pn���Yxw군�S{�(}�����k�
��p�'/m�Ѩt=$�����}�i�Q(f�%ç!��f���'����y
�r���� ��v�,��N��c�����J5zx�:�~�Gg�^�.Ș��k�|C�#&�!��spt�L��F!ݎMh��/�@@����7r�rBM��6��wzN)�6;a�S~����?��p����=/�>)�2�(�d�Ɯ�Tw�J��_���(�m�Um�(=�.`䋲�!���6r�,��m�DRH�wM��{z��5&5��zӺ�<n��s�K�e;�x�[�tr\S�OW�S�Ry��K���?,��L�=�Cq��yiݐ��,�����HUVЌ��k'|l"�2!���r�}���d�^h*�|UX\��� 1�q8��OL�xBH�nM��\[?�p6�ޖ��U¯7<	�Y��:g5>��[[�!�$_��gO��z������o��W��Q��G����Yko��Q2e�y)�'k����7�"2���F�G��:4�����	�Ӫ��K:KY�LvX�
{�9��V��G��A��l�X�;w�w�缞�0ܷ�
ˮ©߀L��E�D�����T��@_b�|)y�)��#R��aA'6�T��$k豘dp��4�%�FE,�q>��	����D������ W��\DR�@�p�����mRi{L�N?I��AނI2�In�ϼ�;�kZ�w���SX�
��0m�s�%��[���:�?[@<(|�@?���^�F1Bmѽ�a����>>�2���=����O��jr^�Y��,��U0��'`xH��,Q��a�0`>�PG�M�ߵ�"ΉHWih�;�	��hYu�,�CF���C0��}�ڌ�wZx�o:�eɾj�)�6x,Z�5I�Ќ>%�ZZE���F��C�#�m�ڮ���yîy�@s� �h�P���,�[^oBq�	&����&�ڹx=�Y�ₜ'ƀ ��k��y�Ỗ���O���$Q� �j��h��Z��n�r~{o�
���?�Wu��#�ސ ��o�29��}J���9�
�	'�,�l����-��N�{@�A#�j�1ӕ�8 �M�O��;��y��7�.L�|}V�>��-�-9a�\X�m$��i���4P����Z�$��lE���L>�=�R�P$ۭ��j��VT{�C���t���6�1wo,(����0{�0��֭Q�b�p����k�F��i�B���pm�?~���Y�3tt��g�f��l�Ͻ_�龾��ʜ�8�{����4�ؓ]�$��.N�7��_�%�:+_���Q��	��K���Fծ?�$.�a�������~���[i�h��x�ܷ�j]���[[���ο�=�;D���!T> ��8F����ԉ4"a�M'�a���Ӛ���y���|.>�Vټ�$������L�h�y�V��+�fx���"��<��������l�.�ȅ������2��+t�5o%�c�'DN:./Л.yW�0���W�%Fԁu���
���iP�P��M�ȳS�)�\�P��җk��R��[��7�I�7��ݞ$<]@�s4va�2�򀹱��MA�ONĥ��Y�ͼ�H��Te%kV��It~G����Y���;6����C�YUx*��:�i�<�Iq%8�nSg��!�ܢ|x�|)�4ǁw�w�%$4ɒ��0E��װS�h�C -�^���`@>PW���q���ɦ�k�d(x,l����i�^$8;�Ӏ���V�s.:7m�0w��#��[�A�������Jɨ�2�]�+|� -�@!