��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�Y�f�ʴ��d�m���8P&B�� ��
�˿F!����i�xL���G)35�У0�Y6ɓL7ɶ�4[�Z��K!�Rʶ�������*�r��ug��51���ƅdӾǇg!PU�Ձ�j�$�6/�s�����a�8B`F$��cWw��St�\nq 	1�	",pd��]��!i���k=Sq��+�rƅ2!6�!e&{��֍ܮ�� ��k���R�II��� �~s~�d�dOQM.�F+�������1!��E�Y��"�(cJ���~��`�6G�11Ed^�7����Vo�T��h��ܣܠ��*�_q��m���o�r�ah��$_Yp��F����++���ǋ��`���u�&T�k��U 5T�����u��H����Q�����0��fH��Gr�NY�Ic� ��>]�x�G�Ro}��w�H�\�r��K ��-�S�Y��7�ن���b 'yYI.��!;8w�yph�v�j]���v`(9"H�+�L��3PʐO)��s+���;h�� a�~�[��Բ�f:,�Uw�+1ÆpZ�I7/\?�r�9�P�O%���J�V���������
`��'��k�������L=|�=͔���`��
+�]���/>6T3��������5A?B ���tF�񞈲�G�9V�O~lH��?�,������3�|{`�1�;��54M�F���ץ�(���߂�	�B���Ԅ�B:��9��#R*���F�;/&��դ$ٍ�,�V��ۊ������6M�1R}��Q��'�rdy����y5����UN����?T[T}��4��e;���*�1�5�p�s���m�򩋆W���*�
Yhh?mⷬ��G�u
q��x4�o�¼�A�g_�=*�����b�@A�WT#�`X&L-��y�(���ͽ�ȘL�`?��2k{2նY0���hU�	/�����(�����j�Qv�ω�)���ԕǧ)���
J=3�}��H�#�NN�/�HmD��C"/��>�Q儭�F�J��?�^�kSibQ��o�(�9�'��r�����G�R�j����z{upMV��cO��|[���x�!��I�_{ �1"�����4`@��s�7"���F����u��jUA���"�~�QM���gD�[j���£Ztn�?�}b����1_��d�1"H��4�L�l�<���~:S|�­�x0��3f3�������o{�]X}o�u��3����e�Pɳ�78Q5
>�8Ը�ZVMG
VgN��gt-�~������X�cH� ������<�4]#�E��a�^�V�:҈���g�= �k�(9�a4�x5p���)O/�CgYs+g�y��j��C3N3Ϋ��ʬ�0��،��Z��{`����R����i�=�	��8AL�P��(.�F�zknR��r�5#��j��WVLR��V� �"@��/�-G�nF��#iؐGJ��o��E�B�O;H�>�� ��Ռ0���2?��\�d
d�[`�C[�M�^r��h��%Z��2�?7,�Ȁ�(�!���@����T�bꝦ�?���h#� ���v-V
Խ1_���<�� N�uZ&��N_S�#t��NL`���>�������.�7�Q�4a3�_ěLD
'O��E=����yD%�ΰS��{�zc@��y��l���.�gt�WK���/���3O�l��y��ؐ�ܖ�-��C5��vtc�kg�\(P�������
9�S�B��\��ڒ	?��T�,�$���mGDGjԘVj�8K{j-�j  5�a�?Fr$\���眯lb-�NOڭ�=�y��B�Y���(B.���!�&�q9s�v������_$i��*:�c<ȗ�Ƙ��to��p�c�I�:R�Z�X
'�
�w{�z���@Ʈ]�F�2
����
�_��Q�'L'L����'ʦ �ް�9\�yY�(����P��T�Z��ށH�.v��BW���A�Aj7�E��o"�O%�����a}�ǼOd�_�jdy������t$}�K3o�;;8A0+�;8��5�[s��t3���Kp�/����Sb�X�:�<�6{�kֻ��y�S⥠ۻ}�� �}p�"M�m�@�� ,�s�����UuX���<�5@�d`G�+}�]�s�	�*4�O��q�*)UD3���B�� ��M������XX�æM���/*[��	'�2���?4V�.q5���+4�8�e�ȸ�r�[@��A񨹓����g\��u��OL�,�����0ɞ���b�����q٠u�9P�$�����2�9z��?#�:8΁Yəۥq�}���剕�'����|T�㕋�Ҫ)&G�HQ@._���J���n�1 ��FZ�=�z�>#A������T��:�M���PJ^YM6N}���ٴ �/}%�q�PȖ�P��ջ��odyfT$~�����z��(.� �/a�L�|c����<���:�� �[;��I���#@Pm�$��$�H�W��RM��X��#GZ%�=��k���z�#��1ӈ�f��x�q�_ʓ{>B���C�M�ub�ua	<�트`ER�n�>) �m�}���EY�(��pvmjs#�<�>կ�J+�[�J�e�WgT�x��ҝ��`6x�D^��;�s�)nP wr?g:!����pA�������������A>M$��2�f�,m.�əb�������W��]7H���0_ђB.�k/n�ً�Is�������z!��|�#|/��i
��/sx��$Kt�C���(a�����vy�Vѯ:tsx��x��C9G�EՑ��!�s��L�t��3�#(B$3��C�5����92��2�d#�+�U��h��	|�d$��q7�t�"1[���#b@� ��Ha�U7<n�[R*�#=oY�Q�����n��v-%� ]�E���^���1Vu-���FhaylD��X�-͔t����;�9]lZג3�-��A�`��&Y �q�N�Ǐ�L�D��^�C\?�6�/鲕Qq5E��;]sef��s)�^�,JWA�Y�~ �2h�h��W���$F���g�������Ɩ�ǊD�������Qk��6��cO��)��V�
�Zd��>F��� � =+˒7�߾�6��u:!�p�1���Gj(6^�ˊ�V�?�oA	wmn&\-٭S� G�T��["8�\��TcM�i�}:!68�� H�zfq��
i�P�v�Z �?KE����>�:u��el�`*?k��P]��t�[�z�b������ӣNpG�۝�.|:���H��{�r��=�k�|�ԟ>����k���=�p�y�͑���E՜R��m���"����,��:�#�F��|����6�p�9%i����L_A#������]�9`uK���9{&t(q�<�!�
��oLR�5��$�!���t�!�+�~ZԦ�H�k�6���ص�&��+C��"Ym���d�J�n��<Ō��l�w�����ĺ���@��r���q�9����J�	��:��W�n���bq*~S�jc;�v�-����oiǤ�5
�so	�ֻؘ���V��{Vmb�e{>P�Gh�r���Azj jN����R9�+�tʍ���d�Xp)�KMI��5|k�1��T(��Q來eE���p�&D���E�
���@�RZ�(����(�F�<�勅����[9x/�������r�b����,w^K���\+K�JL7�w�7m�4�a��k�8|���f��}q�P�+[X�`B�r�d&7]߼���3f�̨B!���p�~~�`�C_��}�����Z�b�E�-r���Z��eԂ6��X���k��r2�>}Bt�S��l�Ե>Z������ɬ6�R[����UǼ�+J��-�"��|�����}���p�뻢��@�8h����r�Rl��#V?���Q>5��C����>]�-�V����D �y�'dQ��a�2m����L�����i͛m֙�jے�W;���Ew��$�5�'uY��3N�bB#�܃���᲻Z���!깐���V|�d?�r�,���*�fɭ�^��A4�5��}2�;�E1��N��+�{���@.OVӠ��`�m��.3s���MJ�ҽz��U��R�ǈ���v �$��S-z���#.Zv�u�|A@=�:6���o+�.�8ĝ>���^I�՞�C� �t6�]�O�|�b���4{3ai���m����|�l<iZfH�F���{�"r�x=WƱ"�^~�-�%��K����&=�NS6nk}�
齆�Z��D��\����LS}�@&e�� `�����qXniHׯ��<?Q3���뵐6���x D��+