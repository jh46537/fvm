// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:34 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fRLKroGb/mLOe+PoVksMBlBEwV1c82fkpbkk0jrJWKlrBxRFbVTh082mnPVdcGKo
nOKLAhWwA7/Qjo7+dyeIW8APokCrWFHlj8iGJdxp7ISrugcBGnvQF5d0pSSfyvDc
c5vUkPj5vK5LHAQeE/+ZkmaPi8n2OfaIe0HgtsgHwt4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5568)
kpMIepCabBJqylZ+9gKmvhGO+fzn2KcO51aeB4Kpm4fiTfADZqfA2X/KQ24LPWMe
9r7bmWLSP+E600ZDJO290ivO5361NT8p0gUU3QU+TQg64iVt0oAiLZNeShu8R2G4
bPk78vDYulPNz0hdKZR5P5P2D68i/fZ0JLCwXY+mTiJykeIkx/8bVH6YN9QdjkNT
h4jd4UnKGC1kIfychGlVjhSrmwqQHtiTvpiQvPLkfms3al0xqb005/Lzu6okvpKb
w1YXjrXng1NucY1fJJ5bLqvIJQ/YUr2h9idm8Zqlc3uAMtSO3I947pUmCpSSYJFG
KBibxiZIsgwVxt6/QP6cnsR6R7SJAAsMAOQy+/m9HLoy4Nq3OY8OdkqF6GPwUK6Q
zhQ0+wjZ+oTJ0wREG0gti/H77dR+/6B4TJqy13zoiAsOSJcLhBmxxyVsq2PDU5Vu
T2tGZqtWSxODHeYickuDIv+rn8v444QLcKZ8yAeh8We3G3gRlM6773JCdlltLdpj
dBMjvzTNQIAko7WUTgQox67OwlpUwc4l4Abu10lgnKM5e7DBW5vWVhowQ30RpNgX
WVBNWzTbAYxz4oR772aa5IdL1Q4bD/ekkpnibm4XoAnq8Svpzej5cIoY7y6eOFLh
Fz+CzBQ2RINN/X8I3kH7dYmgmjbhpKx4Clvn+Fiv4Zn+jMjKpBkBOX4UymMfq5s7
15jKT37LBOzG4tUA/pVTC1yp5tyLctuDdZsR+C+BHyWTYQZD6n6HUpZK8zzY3OUI
VWG8fEE2K/PqSKXpy8QoyG0A/lHZPmAQF68YBEut5H3acrew9NawABgX7Z+Wu4WQ
dhd4HX92VIFeUpGjFZIbF0lC0K6cdWqhUwLUV7ZEpnleMZ/Pa6E71M7aW53dYq/G
mvAML39jwZKe3m3Yrv6xIUKCpvZ5ufDvDR/M2H9WJwNXtArOh6us9vFAchSnqEDv
U2YWzDw5XOvHOZOl3j4zhwcl8CTCMOyoS9GTBOzxsWLhchlo7987eWvj1rDM6pQ2
xLsnl2Uy7WE75bLXE+eAwKli9gVF5+kA88d/tmALatYUZL6apnImQJClTkHACKMy
efw4WnjtgdzpJDhTC9iV0KtTkz1aKiAZMUaRz4KqSI8elBJYa5ol4cyZdRa1CnYk
yeRQEUV52CvXcJG7M5jIMFKJHoQHKFWAsfcqVNRIALGaaPmEvncVug7KIAy1/NMF
2xQxTfvCX0yzD5a0Rt8KajTq4fGb4atQ6OcOmcZNwlWlWtwea4S3slWOayVi62x8
dmcQjGgWNbsWfdbr5gzwTmXI+P8N4s1Gt9LS+WBIehR8hSzjyyqqv+s1SYoJ9DvP
yjjrjYAB+gR13cGkaj5EVpYVQmNwwrHefguuXlC5IUDC5D/kjK3PE/LM6LNtdqMX
Vb09Ma4NieA392AAvM8riSO7XxpRd5ERPibme/ZsNbdAdCCuHAZemT6grdyaJuRI
DvUYiz1hOEoPbbr4s2ZtuJNSaeKlPiOjL43sDaTzG7CiKeq73hmnex1BXUQZGQ79
znwAPqZ3o9Wb11vEptVSI89chV5fd4myZXKnKVubkgftHh8rLLDAp1+1y5wKfg80
NfX2EFp/pKQffFvWUd/GpMscVHs5WO5ASRKBv9+M+4OxADOKSgHuZRiV0cYEaaR3
S2lcLUqrLIoAhizrOFCKujFC6zyw6O6aVm54/KYrckrhnrsXnIgYGHRc6LWCv8xU
phmhlGEVCyXkfxij7V1CWPsk1qqKD0sO6J12OYkmn6Vx60RtFOJrV5iR7ujnFxLI
vTyCZs/mHrMQeJmtcqUS3xydgeAJyQnd6n8lus4gg3kduK0nMjm7qla5JILwlqQa
M2h1QjnviZeQkc3hmpy9lha4hD7kcGGLxCzam9LiqtL7k7iHA8Eq+WPLCduMhrWL
aJeIBcCN+A9s3irIqsuoKDBk51kojncj3Fa8kVEQlg+0NWzsgwIi3tZtfFiIvzu1
o5Wnm6JoYF8bFic3oifWqESMObc0XYmZWSJtZ6Wm0B0uasMP/crlG/vgMuJsl1oF
JeILxjMJqAWjDELJQZieEfr94aOHMZyMOLA0qj2weUcQHeySWY3DWtWTnMjw9I0Y
21YmdO5pALfytkyjkdtZ41P0XJntLktipB/BiT1wT+xK9s4iTgHlMjsDCbra0mUA
4+UNesbyzVtusKHt2UUP3uehES3PsqeGPrOTtvwLx2sNgtmyXLUobDI830qedfrZ
ze1YpAreY7Ge2UAgfzDVvKTpfeXDSslydDxmWMKtse5VWL0MZZgdCB/G04FRKqXm
aFRCxsEyFNFfknGJmBhFqflBknqKSef4yZmNoS7GfWr9jPzqlwcXR/+IrD5P8IfC
gTzEWlpw/rP9NNd9AAV8g7lwSfrUEshLIUzE4d+I9+pB94C1XzVeHtGoaOm1GQNr
iKlAebmlMJU4XzCiLFtz+AuyrScsyrGT4SO7RurqlFljIv9vTuJyOjgC8czg5tWf
4z+/xOp0E4O0ChriqCKAM/stGW7GvowifDH/KF87iwbDTsKsfQhD9c2ljBevf6oE
jdafrYwG9LKkpw+OMdMTALHvnuMTnAJA41Qp5ptJ5KzkjDRt+4+LkLk9UC0/TmFC
VEy0B0x15XWhNCCRKCBrj3hM+FbVvVs89hAyiSIXiYizl5Nz+N6owBnAb+ci0NQ0
FxNGnYyWJGXI5g0HU5soWKP3v/vg18aks2fV8C0JbZOzvaGzupTEFKETQGFapRYO
SotlFxzmbbG35ca09ft+tJc1JPhcKi5kKh431ldH0CD48mlsHQQBR9jHZrJrue7Y
f4OIsHGfsvualiNRUzh+J28JMr5FNE1xrKqyqRRrW7yszPhjJQMvq2mK8STaLczb
fwavsDnFthsNH6dHn/8frsV/VB2aeTtKZ710s4BYAr3ZD1lh2rkWkdc9rxHCZK4p
lCA24TL+VKHq66GSDFi3F6JbHmbBMpjXndHbQUtdZdxxOmSvnOlXM/LeyJOdmcfj
K2x84rMCq0seP8OyyMD8yfVbQdfz/a1epASUaq2hiOvHDpUq6JYXKGhUDuf5arNy
6rVKa+pziX1uldrFNpXe9WT+EoDV7VU79XZaWajUKoxoYi5K2LznrE5fVziDhSnd
MdtxEI6SAW3PE+/07AQb1TDSARUNRMCLUEoLJeZXGSY4FBtEvTWBVNhwlrjBBhyU
tvxxGe3lNxa1y48zeuLz9pRQ7zZu15BWCaH9OVpF37TyHU4ep++EGm9bJvoXXd6u
TnjuN/1I5oQhnCSTe9M7Y0vtG2v66mCr9c4Kz2oRzAphceXoC7i/cIpx1tdcw7Yz
TiKZW0vFhEwBWk4p/xzD3xHD9kVCbl5/dlC9NOEma2zBcZj+qP8rV+OSfiFCi94K
/WWRbDHzJT6/01o2d401fYmNDrmw8Y9VapSXHwJZ1WsVKKr9hOG3bYe0MAzd4vyo
t91Uv3Km2jvP4jMfgV37We+nPRQcV/AhBcEhQIe67gXEVZ1QqdRIrw3v8suoKKR9
/3XUHH3a7aMU8wo96eIiXFU4zTW3AhwNNJ7PD5g4ZXSCEjYy/DQOXZBrjhNC8VeO
s9UzgN9IPW+VX5Ec+c4fJokB7lBzX0cfoiAX9uZRvgeBVqwSpXPmJDkv9g9GpYbM
oVpNBmq45Dn+Ik2ZU/3cxhZSRqkdQ7GiF+9fC1VKO59AO6odwEML6aKKQR/1Cxd8
/sRwa4DDAByqlpatj3JdMsrSWByzEUW8NJoAQkwcIfPBQBoBn9Vu7YX+Slv/Ctjv
5E9hY46UgPRrXMIZAvwP5anAq3x4yJfQAtyx64Yswv01dKG88Y7S5hozhWmHx66M
e1sY0zDhw1gJRYgZXTIKFDAbaF+iFtVO4q4FeJmd+XbEiqOSYDFS+vwejneYoAIU
SdsbGqALQ2pDh4QNhHW8C8YrVGwrokW1RBemwIUmf6VBVNz8E0QOldxTA6Yn1d8E
MA0YqTH52qznqZmQcCxbsoz4nzOGicK5/iQliS/57CBuuAQ/3JAJMMqrn9ZEwHrp
4hRjMVK/22TzMBBfc1+e3bhBQ96gezfqxED5WhQBVn8oqBo1mtNQwO7LvYAEWtIl
5xrVIiMBLKvWDP1oL1YkBSouVK4Meusj8Z50jcrb7Ayr1TLdZRDDjR2OzVoEQ5Vr
LqSxWX67Yh4ULGec0SuhNGHOUrRH8kBizSHvVqDb58wi3cNjs60jOA7PwReFqWeB
kwOvh37MQf5pfDMzNtRFUx8Ax7ACgW5tYAd2UJeMdwaljbRYsfbfKi/ByU1savLA
7Dh7WQZTjSzh1Sfx2bjqbPoi87M3rhpWCJWVahQ9pTRqzUskSTl0W9HiNP016r3b
EG1nZht2HvRY6PXniiiej9TwyAdxe+K+sEzovK+3DtwTZUQVPrrEEL3VAULcNicc
/31OKi0NJ8moMjBS9kXIdY64506DM+pkvCnpKxIUwtS/+u5Xx4LGgrMJ1eCHYdWw
0ZUa3Ekikpmnj5Y4plxk9hR9tQkkE2p5rWPJDvLrW4lxrFCdVv7eK1Xr53bXipUq
m9mcBDKuP+GYrNp5+5OpsjjF3wzAyISOqyb5HJorIakPEYFHOs9uxZ9PgTo0Z1Rm
cHwqLnmug1Vc+5qwtFjr/oBKr/ljYjHK6KiaG6zV14Y06B9fW3Op5ijMFSoLor3v
yVEVIkBXrA7eh0w7r2oRMb0lGMBoFx6Ly5X71qf7+cuJKLrUIFSzAp02X30UcRAZ
7fdiLYR2rq4eO/23nmp3oUWnr0Tz1NIGG975Oc+W+1Ifl1z+EM7bznv5BVKruKtD
wAVaeXYkU2EJCRtJfV9Oh0MCUGD5aZnJN6Habj6rI+Zw08mYfjNdX33wolLIs1lX
lcQsDXOU3NlYvm2z6g2fJc6y4WHHfXXu85Vv7Xodxakl/yoeXp11Nr3M3WEh9TPl
61VASDm5U9ZqPX+GBKrMn1CweuCFEqrYQZ+/WVmllV1FeC7ERhktAwMlFpmKHRwg
KYSVQjCd/cnHZzvmb9pWjBehYpoooteFMYHPBKVssqQta8SpAs/oAb2P1J0507YA
xKSojrKsmIcK0OYUlN28fl6ZkKwP6f485bTqlcTTlMSH1HP1HeJNosbDs2lI84sp
W2mKFnjwC8HGhUBBW26qNiUGjlS38PfAv49Fq5nh79aKFHMicMHIu1haI6HGFwK5
1piQ/McCSqukjOc+wxExKe126DFY2UVYCkn2FsxAjdyNQ5qs5BsTKcGY5hFjZDVk
eSdwipXYsFAh7EZjFZq0zF4su9/KrgvTZI+i5uqM9DXvYJBc7cf7u+lmhyQEB//J
i0cvZTwA4X6WgaDI0fU3HPkGX1sfD3kBkMRR4FiCTjZb8cwMbtFsLAi/+Tnx6aiL
JHW9auvkxNry2iWzT65JNXMSHEcs+98OCxdBAakNSEFGvPVz4/suoEdeBvv1TBvP
b/9zmNhWJJBSEutnhE/p/wRtu4s081j3nFtqwFNQ/LX2ZWUUB6Ty4qmEzV+gpdcb
FY6uk2cFd6CoNeqkoW6mA1y+QISbwYZh2PlM3LVq9Dbx6XoAKO94oAGf09m3BubT
/zWnufqCoqfxi2RtI05dny8lOrhdBQ5/AKmaHtrvtiIWGKef8RG9agEEvSOQIsUg
5/pxCQb0pVQMBejw8mpa0Gb4ZCmip8f7CRT2dULpGIL3SKH/SyXEfT5XEJtrzlOJ
6MAcfGVL0tiJfQxNfUdAxUZzWZqgcjIDW1/XCKz9nAkLcPP5faQpLmQDirSm34BO
lHUb2RVT+tRVt7+lGG0BKn67+Y5irpoScwJemI6Iz0NR7azq5iO46N9HYViZK8/0
JHfq+TiNYK7qqtJlfTsrnQrvFIRCdFLNRp/FEsHaej4lNksYmWhjbhV4RQm1jUh2
b+fkS164vso9HGuqUKHwDQStL+OygHQRXppescPhsYeacbYsSs4lKOucQUUxAfHA
dx4V3tcg7Wrw9fc1QP8/abEJDXDTklmvp4B/ZuGYvI5al9JSEf8dQsBGR5L6/fEC
ZAKJ6LuRGtxZL3Xc8K5Fui+2hoO8a2Te78rYypClah5JgL8GcZSCpj62JjgAaSXj
VakPUavQU7L0gdBXiIrVR44TISzejcyhYLLomSiIiNd96G6cba4UHZttz88OJG4k
3Tnuk3l2G8+VTlNbv01XCNRFY7zyS8zZJq0ujAWd0+6kX7d5MYELhQbUdxs4j3uO
WX8BYLrFCBZXGRVZ5CIFe4jkmeM0i9pb4+1dFhWLmx0vEZAzHM8i1xkiF8c1rQ4m
8BOenyoIf2+BaHbTZWPn9TuKhldnfi2c/JKD70sWLsVMKBKMDRE8wPTDSBspq+zj
LlhIpnU0KpTccOz5Cz9LGgGgEDp1rWPUYsfcGtTTcNWFcFaTI9e60B38zJyq56/G
m+4Sf65JPFKNZNGT1D256YPcM8PcJpjIioUJFurZT9v9KA+m7nVdSrlaCCXEuGJH
c0dI8xa+a42/ZNspIqBfCHgyAgWGG/RSQD+N9SlHnJ6ZfG5BUwT2KjwHsWXX9lFb
ggG5rfC/lf0n9FeNyt3QSJHGsPS6ohU0xN/bNwtp+6j3nEDARNdJXz93q7BMw7kG
BW6crwj1KHkhWTNelWqCNYcF2fhjCYU64ZxegDsb5arvjuLtQ7EuTGQyEhpLRq1a
cGsPCTcptMcTSl2DM/fTvOMi2P+9iZPCn/tJsXFRv03dpnmUM/BxEM3cH00kfQ1c
CSAfU1rqEITQcIOeZUUX+3+LWWANeEF5xzydaeo8AIVevQBsTYBTZUVQ2uInpTrL
llAxG7CTBtLFMzQDpME/0qDxwvDZwBD0JX3lfm+9WYp40YCpES6m08nPgAk2XnLI
C6UwKMlmJRwHcJ5j0WAQRPrzpxyHYiUYdjw0BxxyQ7P0PUrVVC+WEhUTPXZCiHGo
kd3W5CJMjJMoAPk4Y7AIi7o4ECxC6EbPQFcGivkdSEbP0jR632SKSAVZSwteR5zt
T/nGSry3/+/TloS59qf8wxQ4gyREZxXTNBoxJjzBacSQZgdJRroFklKbS756fbf3
8Wu6BdbTlLExd7EkWFfcnpxTouBNA816LuFx6ti8OTQyEP3QgROXz15cFzsyvPQM
u/1Vb35lrIjkYbtlmRhe975udMVqwlaJNKTwV9vbNNS1+yCKsjHKL74LcGZImSyG
o6UJ8Enqps/meysNhhlDa5nb7mJUp0ObKwtv3NZagEqPlQPf6kccJhpO62ZvMnIf
NASd2tufRGstqWfQgyJX9HFc+5wu7J6iCU3RGzQyKf1TQmql8XIYyklDmCRMIYsS
FQYXHu1yRRBWKVGR4K7dcdPVtWYSPL9pJyOvQMvq86TDn9dIiEBq4oZ7AxP6862w
Q26kLx/2iRMNZOOQSZQG2ht06dZbIw1nlQ8/eUG7bmg9iiNbAyhoQYfmkzJ7NHj5
`pragma protect end_protected
