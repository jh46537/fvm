// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.1
// ALTERA_TIMESTAMP:Thu Oct 24 15:37:46 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iTeud6t8DF8XQ4nc5LIIikgZyf7Dm3aWiA3c+2vdEKovs1/Yma0YdsD3vR2STNjE
RaPq+yhobXSsGLYnz2/+sO6XCoXSnLcGKEG8O8vNLYuDtYE1ZPxhx/ACTMnnNnfY
uCCHnVAb+JPD/X99GTXYiRuQIPJi2E4iiiB1RSsEUxs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8592)
5UvQjhQNu2J+UD5yWx2cHlwgF6Lu5qPKAGXISGZ8elcHd2swbq+jJt528nQjPD8Z
BPzqmehT49iVvjvvGx0CzoyasiMXbLgtPWh9a7hlKwwozdKWD2KRhq4bSmBfQkxO
t2IsSKvHXjch7toIpwDJeVby8WIRqHY0NMeSClo7bcjvIhykMuEuZW7A25BXKkYU
EnVbdQhKxUBo2Zu1ZNYLtxNQqcxWEV/SjMmkTIC5ZHsqxX/p345wNUrs/sXkGKqF
WlP8uqmkcmMa+XglLHqjpjwsj/tlXIEeu7yN3xAe6gDgIeGJ9xZrmUedf0+HzbUB
g17ONFdvzfTwBAanxFAgxsi/OlpLvchUMnVvtV9jcClmuzc2hIvth7KlNeNUQZMz
lquL0yx6LjuZJgtl+3UVLnvkXSKzRup5qfC6X9vVe/wgeFB6d5XPDJOwHjzMZ6S/
7Wl9zhw73u4QkJlr09Gwo8DqaPlIUvOrJRSLd0Y6Ofy7uRggN3LFMf4kZuXloWwv
kZg0+xij73UQz7eE89UnlsYANY0uPlvUq323QEPaoIxFUIxxlXogNTCVVqfNNMvl
1RwI2xHCmrEgpec3kummBph5u8sOfxoa6QOrjdDfrO/00gmP8/gHlewsjiRYeyLK
c6OiURGOmBdCB0IH1uyxBejg2O++1To0oQV042GMAsxMbGlp7FEy0HiANnVIaN+y
QNN2HhwA//mxdjTBov+NsuDuWTQkZz59XSyNyfcgUzOtDAyUnKO1T103v5jVYde+
ViWGGWreuBC2wkcFOTRM8CzBWDFKFr4kJIHqG+ho3hZJ4m3DUipzsBQXHMtY2jiz
dHHkSRFQd92LADl6iUI0UvQ8aJlGa1jWkl19asYFlsEDmOtIWmAMS+7Zur1VDaUW
7O3QYpX3FpNKwSaAE3TB+XkncvhG6+CnqzULBHtK1XwYaW5maDfPx5ba14Ukzk4W
9+togyD8cKqjkBiy3K7FzAOSYc8gS6rnB7zdhgEb4auPfpwAA1XEfgfWnVAgq+/j
adqPvPh6FSCywKmmULX1dUDRY9szQ8medjneaeNFJdp0UogGykYGOZxMKuuPtc9S
uP8078RynS3uH+kkniyyreW301I+Z0McWaAC2FOwjwf4DpDPYSS42XalRt8+i1cY
3NA/FQnIEL84koNkVmt1gIx00dcgKpJFxcx28njioywrQ3o2d4GCdGmiMu53Vvte
ma8bRb6UAskJj5F1VLJ5jnfzbDlYAx7Rb0IoHmap5iNWBKCUE4PJXMgIKEmPISOe
gByarlapM1gxJ/qV8l4nCnQT43rX8wxlXpu5ehHvWDNkGrVPZB1E09wur9Wnk/AP
LTWUoZLK3p5J2V9AXNo0Vmc1Nsgv7xgqMM1w7Mj6ERzVY3UEIEcofH7SVkqPumg8
WTdfA0BJqbunXPQChDLEM5xfpkw7QC2jRvJIc0yWQcKm0C8zhDxuFUoO30HuLvHr
LIgvXMXscF4e6M5alV+5rjOuzHOUfuHLznn+SL+ZD/gxiHyKpb+TGLIPdHwQ1dwX
Nk0y6Sf5UWnCkZZaIrX3ILzFdr49wwVMv3uSPqUb8wba5KtOz42yL1+NJVQ5yq/v
uvVyaZZ3zRvy6irqE9d11JvIA4p0FxPrNSpnVoK3YL1iNTl2Y+UcC8+b8IF6g76y
FlvumFoIPPBmthFDLfETgLJi1gRNVB19179HVnbi7FeOE1KrMFgR9IDBjPGLyXAG
tktuQbmFv0e4uU6sYP6MORIreT1UuDDt7tHKb9OxCMfIDw60ABcdnVY2T0dbxRgj
VB6LSd6a12EKjK5Pejhq3J3vnM5BXRkKKpz3Cyow/Iw7b1Iy8VwAId+K7GMtehlz
Y62gXDL7T2ehS3VABU/l9T7q8wIx9DgTHb2ZHkxTdJNhfpYiD7AmaF8kgzWkBGQ/
fcjAoMfoQHgmSTWnXB7dlMvmPV3eU/TrdGHoNHo+kfDP9PfGqd5jElwkE8izPLxg
CISNxtZ0CFO18exKmAs50uza3phGXDBuXqSpKod4iyq6WjvNCC24byh7CNQdtlUR
tR9RPbD8t+PwASbWP4sK/KosiAvvQSPs7sTgSBFuZyaS2zcdDTBlcZTqMTB64o/S
1W30m8QqAYOF5sGlPANtlFy638msNl4fZ1YW/nprg7OPkxC93/AQVcu0/r/kcMmv
CeEcNY7q+DCQTZpAzhXcXjPnU866AzLXf+LVtf3LpdGr58bEQkNyAU5mWIf3QN0/
Nh2iDH8W+v6cP5TyweQ9mbY9x9nURM2FtOSTtTG2kP9at9yat4QSl8dQdXanr1+Z
FACWELpbif3FsvbdcEGTIM/k8P0tL2E839okpfWMk6VctZN3rsrIn/2ObHqrdp60
jN0TOpvKWdYeLwGG4q3NiFJxekiLJP3ap4XROaWkmyixs+qGSftW0zJRh1OOWXFc
4FpVWsHTqHvk9EXgCLGGc/nrkmLHyKfm4Dh2YE9UuBwKH2GU+t5CkCeaHeEzU7m5
N9ED+dHMyTaN6Wwt8CWIwvYnDybbEwi1ff89+62REoit4CaaaD3imaaniMaclTJV
VGx6tVHhE14mQwNqpVvvdLbRqRPiQGTCgNPJ1iVwZaaAJnrtyRhWIfEyHQbAISvn
IQKXxJXeI+LIbd4L6vtjcQzxUoouucgFz5NutslX/kKZKKiWZ1jIZHaKFIMoykRK
j9UiDX5Iz0yhTjtds5cQBSGReSkZI6L82svaNJEVcDUYwHAKDCaN2LpE7Mh5xguN
7NCGFUyWKcNkOmL3HFQLpXjHgtzkGCEGyl0ECf0JB0kjcCD739qJoIeHijusNfpo
0bQQ/Edg967yW8zhC81T1OgOS1DhNvCwd9UnpAcDJeZDmHBRWnXEGTre//Pzmz6Q
YVKvoWzy7ngnMag+A9HEY1S5zJ8ZB1YqHpnK8urNfqUxZ7oial10JYIvm9Wyg0HO
X6g11ZuEzJduBUwEuBpO8zKrpxPCExEibuhrrdtqELTFN3dj4j6ayxX0XLifx50Y
K0/yy5q5XxF1bSdMK6jLN5aQOAeTl0wOAiy28aMMMDDBUGCEdrDeCDY81bS0yHc0
BjQn8z3RA57eG2SQ2aO8d5tAzgJ9v8Yl2G8ykAgK8TFBI/u6l/eeU4efCYOpkv11
6PFtXF+kgj69MGCN1EOB8OaZftA/RMz+vGyYiCe4w/9BYcRqv1AnVsndLw5A5Lyb
O2SH+y4cVLCG36UkYgAUmWYg42MnxJEN906fy+V6o8riyS8nRICHZupd5epgG/tS
/aw8B16p7ibtAkA0J9kMEVFGpi4RZzi7wQfVkfwL4/CamtZDhm/WiJ5zoy47zCt6
OC2W2lcgtjazbFvzcpvkPSMdU/9xGucVzfZpfaJt/t4FoQ8O/wZPWSiJGd+BUBdu
pjrXTvVZlD7fd/rYm/ALZ+3Wp+k05tw68o49cxO2Yvjl7hx/JISAUnAPHI/IBWPM
mX2bkX8o5FcSpvB+ON3pkVDhQuWLoAbtEi+63vJlmeHFmy21UYvuMZ7+VSn5fzDJ
cphSz9e9rfqNCAtcoo+ZfcGmB6XvoDyUnt10eseHnK8t6BXQIzc7DKmRlmzfcaC9
gjzQcW+bTB0zeDJpMs9QhCgsn7HXnsaeBowfuHU6/6WDsb2zbIv2Wt9rTYKgydxu
TB+wusTztSVJwq2E6oTUN1Up6NHVjQWEaCNmGMYoa7869Xk/IvzPIpUnElsk8Bgh
QLJSjjnO1r0a8KgbLrWkEjHIF/nlxenMuI3bMC5qE9Py90ow44KykdZ/+ih+Pq3w
a9R/uvYM+Qw/ygsXX5xznR15xFARXNQTr3FHxJWsw1gm1aqAaOiPd2c+Y1EP9kDC
T4LMfVIspzuIcrwhJKRWYRcj8bOkmGWVOJiXIGSdgiJdzr48p26KVUfsnGj/OKf+
2nFbGH+0jhvBoj+r6Omo+8ABUOxR57JOWUQ+4uQPnhOJnEOI0oc4vbLt2j41xUWC
pgVLcae6Zw7ZQSfQs3+FH/ze7QzvyaVO33L8w0hgKBhmRcffv8ZiGIAs/iEdh7Sl
W6J4tdRUSPbJ43gikrjRQWPViO7Lph8/Hl4WQ+4Dtt5KJWvHk3ejZOzAK80740SL
4t5C/1Yg/LGmN0gQHrCwce9Yc3IItHwhbdTuWUdaLFZ+DbJA+dQymbv1b5/uPyPt
a0sQBjXxc4DatU5JfOIcL1H5Z6kQiG1ibzxuSo0kmHPmxoaurkN2KjC7/3rhgsva
tzUxXKwot+hmfiMlwxP3HNuB62tizdmXPdn5SICgxEB/F9tQcD3VSvutqcMxerEA
YXv8qC4g8y80pNTp45YVKWRFhFJlJsjnwkHBiMYf9nIV6GpHrlsQ7q2pviO5JtwX
AWkGUbQEPFhBdnOgPPQOvj1Ap6hqM/WMjNNgQYR28nfmI3PfkCIRYP/m09BnoGQU
lCzoFjdhaHN3cTQfeiUCNQqzWzi/IYyT6+sKonsVb4d0sXxFiz8YJfh2W48UKN86
aVqKqzBANkGXDQ1LN7/KRqBSY+gEZBZGElhYyPwFhq3VPCjboJpbEQ/FAreyQicI
Ub7YXLydkomDv2TCEKifqKKXxkLglnQNkYsiMUejKFsn0i+KpaZ1RkDoIqu53TCC
GSPBmEhHzK+KYI/9eVwW/2PxsBFED3UBu4isDXqDanU77EG8CqmodJoCmKfneuno
ek2O9GmZY++UNiKSp24Pj+16rDh+S/fVWaujR0Qh5VvBxHr+F0uUMsM/Y9/JlJHc
F7EFYdBbZDvXTaATPOkBncUvIoiJigiNNWzgL2XE1s8C1WLpjVbA27lE9T5qoL6P
2pTpwhMawjBn3FEZlqOPQYy+Q6iilEVhHC7caHEx8cagllndd8jftc6oEFkBVXy6
kYLfA5w2TwU7orxeWnOln1RX0YkMfSqbhJ5v9QOCHDAdOTUq0GmgrY3M/DfMoBXi
3parlxxMqd42RenqEnRQWxe4ED5rLDEJJvTfFjPHuSud10XNBxbLnQgbFUuEmOZ4
7NvEOm+U42RH7BYXr6Jjo3KR0kEW39Q6nohfRbEqm12bv7VFRJGMhJOxBXJ43iP8
I7A5Xg+h1xKe5VbqJQR/EPoqF78t0oYPFr+doGbcq8j0ypIlLuy+XpHXx7hXKWXw
hluseKXhUS4/rO8k1kZ6VBAfl0rItefdbm5/5x5//43RNOvPPQXKbFbDk8s6MMW2
sgtZbUEHlqnvZ/73cXwNTu1nBPE6C/qzKtfXdeLjUxyjRC7x2QIUi6m6kkCrkL+q
b+wtC3nmgFs7rWLXL09STijeJZIeUzQOkDgUWlVyr50hX2Ocpv2hMuYh5lqgqzpe
RHLtkpqT+aUSpX90HP6+Pd6tgSpdIg7xbjl886qvxZ+Wg8IR/O+6DlHL7qZRu4FM
M2F64DhA2udT4aYe4H8eiJeIvdPKHm3k/Qoab4DIdtqZAWyYX/pQcZfVAOvi3hHS
HM78YZurEz8ENXALQyZufOi6Fub+hPyatVv4tsDVAmOIaQBj1AtRv9C02hVvaoAN
dBEo6cyEIVtMuF5iU7KJXwD3/yEvOQuuF+jq2sQSJEt/BgtWB9ygFG6NiVJR+LgB
gJJckeSfir6o29fAep1+qQ2XLMVQ/SNVB5drFt12GldUimToOKIJsxu0fuNB2O8a
xSmt4skZxc9mD1UP0Z4ne3Vlo1qXvhHEby9+yS07YTeWgRCANMskOMt8mq6WR2y4
HFlUqViBJMRUnqka7faoPX6H2YkxUbCG/rXdpHFFlK3BjokbhcV0JvTYPNpMVzC+
GrfybcAfov4jtwpMcep3ykvn4jaKKyZkrtZJe9wij+WYPjs2WgcSa6kd3JNQ2nO7
TsTbO0cmM4NbfKEWrxMPL0mXgMoo8RNgSmS2XaNWG/XGFbSDCeweMNg0r3w81Adz
zJafUQjHfwPTfe7BDm3FFcTwaxX8Am/AQK8g/1Qg6XLW8vlgoAzUnSVEVwsDk5eF
kR15iez370k89rHdlv+mrkJlbHpdkUtzI1jWCJes7GkTbWr2JHWTIGk12mw4iwQD
VSq+8vzMtg+3YgLVFaIFeAIuYf5pmBhfNa+/vtz8agIGie7pydt3qE4SjLBkfalI
vpjRmg4EQ/i95BqaYb88MH44oMkfvtq8F+9aONXRd4n1vOTMCPgQygfQAa0iSLru
Pnq45XA4P5ZJBlVtC/KkWryXkaDRyfxrfKueJaHluSedGbjwQWauu60t0q6EmyWa
J4ScURRirrbTMa8FIJhXRXugslxwsL4qSVedynEr4oCs0TeL7q1FxHIWmSnKcMoc
rFmz1W6MPL+m79KiBOUKiY/LH1lXe5QtCnqGWY4lYBuz9cfc83/k+eI9xiLmkRud
nKVFkemds3tDDY4KsMEp4vfLs5wi2NMV3OE0WingS9VVAXnd+3ek1mhk/7C5CYa7
xfG7aNOc1/uvdHoFRQm9WMZDMIEAwK2YtKHBlJIpl8yaIAQRZscc41FMFJG9Qhgi
aWlY+It7cRwz6j6MEVGNS1q0FxekxY6QWSEb+RPDGjPAoTtRzk2FmhVJPyRBts6v
quRBMJr3G+kcSKW8055zCP9OptyqbXQqnfvRpcDium1gua4nWGEwQgknuJG2T3Wy
TxwWunT/ZHB1J34wLXxZlVaDvV4Z2gpLC6fesFaJm2wEge/5YeWSCUJHDVZ1HuW5
o+5D4F/aI5vo/Ia/Be6gjEn4M/pzHp+B36VfolJXTpuh9xZ0smBVdgrXSubb5s7s
t2qdbMMRZoMoZlFRzDnthsoMXb1TuvkAUH1x5rbINmqlJ9XBLS+JHhl7epoTVBw/
eC7nBgDsQfK+D8F8Z7oB9ex7ke6uoNYhUkFgjtd2exu9IYRkks8xg5fSDMuJQpOn
8kusmYmu5tH9ralNh90jvNECwEjX9ihz3rrlkVrGxLKeXdsAlpIqPpqzklLIKZ4n
vqT5T2tP+vLExLYjFsv/MfZQQgep+K4bNwoWwwyDlkPdC/iAsvnMtXc6iG/mvT/c
x7PzuZHibEPZ1MEkP0w2aFuTBK7CtL+oUiX73LC9GdJr/JPJKzKRlNAyH/QgV4nf
qywK7eGBvGWs0Hpnq/nLaeQvjQKUjrtM74lskLd4fA3AdmJzPZU+qBPDyWp35FN1
RbQzifrgxOntVo+CCe//UXkD1MW6YMOH0Ow7iMYFdRJWYzHt3H0nEdUXGpFUQ+xm
sAxbmBQ767Wgbl1QS4A0TXh+BX0cYI4GbbgUkqJuKXtVxFo5a01IvE+KyEiPBmVY
UnaDjzIQWWKfbEPTYDOTZHoaX6dojia2ub6xf7TWNUSzhsfUPgZkHJUIEPeOaS79
0Juwker+hpA52Gl7KofVS5GFgyOXtpUWbk9iQoy1r0oRkQKWU5769JsIYTt2N73H
sdKi2rLFGHaFvuQCJA16LLkLyo/FgqGFTaecLQ3Y2eZwwaFB5rVYV7Cmrnjm/F2n
3ZKgBhqHtoNahxXu5xPOBpWtAo+Ug8qcNKtT5L4NRANAX2oEOxMwEvquREvkxDNi
iEwzApnlDFiIaVus8MopvFIeOYNsR+BfNB1t+eW/fa9F+axMfrCsoFXuW0hqPVTT
HC29YkKk5x9If4MJfDT4kIat8w/bvVcqBP/175wSqezdQivpzsnTuot5nSk0O/Yq
YzVDW9875ibqCiUwWCKSir7akP9SYg9LsTozY14M4xtK5cP+CGUkMHFb7ynn+0dk
bEDIvMwW0bOJsrAbfFjAQzM79LCt41/CO+DX5ijwTp++9z530srS/5LdkNlSXpxY
xYArrb4CebSc327kC4QqSoPnbb/J4EYxE2QnNpnzL3M8Jp10lIMA1/0D2vYVhLWp
UIkpPc02UR8aGiHhdYS/um7vZdzwm5CzqHvxCI290FCVqaSNuk7B3FqqWxxKRsuj
Q9cRB+ktLcYJUWrya7dvPgTCYJjal4+TLpGK9Nb3z6qtRUWrZRbQHJmcUfDjwFAF
os8V5AECEWAdV1Jb2I6WNFlHd7wToDuMWS9MNoxL+kIZw/aITCNkYUy6SOmJNn6m
bH6s6AvEzCGkX91JaTowbD0tDEsiVrgYVcf+zl7VmdS5chP/Hzi5jmQhwEez6oEm
9nZ366juqOEQS5lbPQxgsCPUIkDHUky0lPE9G2PwE4JlcApc2//gksgzAnvwGfpk
hfhtNO5B237EIdlp8AeYFtNKLghr4hFTCV/fZuF0k+YmdAZj64t7ybsrE7FIg1us
Cu9xYIkzFZP1zymslII5MHXQ51Ak9UKcpj8LD/0IMX6DSPksIk3AAhCFxmVGS+Z3
x0l0q7a6zLGnMeJYEGOfLbw9Nkj5YYs7xoonYzvBIkRnn3BY3n/HtXNU4Cjh+iKI
shcmRLPtfTaPi2Jg2Sh6jFHL+IeGJJYiwxs5r2OXAlBauvtwpEJZTKFEKZYH1Enu
Wn+UCvIVCiTZhOk+s2PkES6RrL9ivoKh6oljw/de6NxqClS2KvUZXP5Z4HehtDS7
Qs3aUfK2t2KV+V5SZ9IrO7YQdRaIdisj5anQ4u8hzkeFh4TTQpmQBtgOa7E8TFw3
JIzKqPb3nzKPNhcxKBhxVOHgLcbZd7e6w/JBfm76JvETB2WflIxHiEGFvM90avoj
limo/MHwiDyvZ1eti5fXAC1aET2dUHIyPA77HzSsDLInX3ValnsCSMXMldXuMHSX
RxqNjpVBTW1kHtStQbXRYg6yoNCwkwIXFX+vJ08+i9b25nRD16loDMCzq4Vh/1Z6
CqCy1ibcZS1bw0LtC3ic/AKL0npLNzfD6LAL4MMUxFdcY8OzZU7PTzyJnWrHjUou
AA77lltB3CSu3NMd6leqlEBMFqqmMbXIRGJkQ0oqgXlG57nt0euUUWF/vyJl+JaK
yIdY2NMkSpgNw3MSKhSbrJxd0eqkpeTzoyzA49+6RTN4LY38W1B8uIj4ahAnskL6
/KLgomNnvcs1RAtPKNl1RYzdpSjFjLHj6fhuBAw53NmIBCTPItJGG/OIIA5a3Y08
7EYQeVcHZQS+PiTriFqiAdiHJZ+x0HvrjowHIwqd94kwApF4hpMmRPkyqpZ5W1VS
BmAc4CkNCtOS0xFlksbFKj2FdMO0Zn4SIsCTX6pKN1+sEsA7M0RIuDo8d2Qr7HvB
8FGstv1WsvDUu9/dE53IHYoo09GUPj6UqDEKDBL9xev1Qu6PonC0cXoTgfRyYP0A
B2s0AFTzjADgHDFQUmeSWW3KcGCT7m8dlyTC/I7r3TJoYSiUPO+91hWgC6nHdXMP
f24hUKzMn5GEqnsbAhMnhaqJj+ZRGg27rFn22aShJZAeBqYxw0of5Q4wzD2YBqge
JjCgVKO+ssJZW5w1yh5Y69vmvTvrVgHEsNOZWuDcggJFR9hKpjtsJS+43TxghyAy
eLAyuSYqMFZ7+86gEyTBqjZ8XKmJjXu273haOGt0OaR/ynEUaCWOLlXut1dMZd9D
DcVURxB0wpzJ2hFVN7RNpxjujFcijhMgjgl5Fumc8JmcL/V2bYRUcjGkrQostOww
WJUdOAPBJZGeucrGeZruc53+BRdTuRGiYNxOulOxD0wFotz2zDBsGNCdmatm4Occ
9y+0i7MDDAJNmbe76isttsQxu9UMlMkxdIrB8F+AJYWnNzHtcZz9bBwj1M6KEkU+
XNsxiCjVPiW5Sf17TKrnuPJlquWOPHnwVrWvfSk/mfJUJbKWmqhRmd6P5csG5HvX
kzx3cLM8Iuu8mWAKJW2px0J4pact++mD1zuJKGwrfEu+rYuNO+UWSc+dyVPl9JPO
WRSCifhswiRBnwiQaVWYFmjPBu8hv9wxYsA2JFMEYHzqynWltcm3h2XADAqoHxU5
VQAciKuN09LOZKCueaG13A1aCmtXk23IO8s/7uq9YM4TVVTRDKa06eDnnixyq7z7
ajaGhaymTRQZghubzz3MLxT8elEHdE6dllJ903WQMHru8HsofpTSAGMtah21jf1r
6mB24Tx9l4IH+5Nmf2F+Yre4F6AmU4qP+HhOD/nBZ1HOEwErNCzUO4tkmASmjNxm
wyRLtZ76JbOFeRVcdjvDlv/cnr2mTvdIyNQBB04w2VKOG9lG5HEAelwAYB+8lMQm
dwfdnrlFJs9TKnn61XvhaLBXGfECfE/qSOi7qraq3RIOHz36EXDjpD92O6R/fshj
VJNKmbQIxZr78kJLP/HrLpjxoaZ1d6uOi+GqKzi16a+/Qd/jEN42ytlWef31sZPs
hYfVElCD0+ZHFcHpf1sLOljQw2U2hb5j5ABOVpdCPWb5Fp/uHeEy4UqwA7eLpmDg
k+sb1UMA6qx/sVqpoMDL+9tNXe0SzXGZtlXtfH9+vCou3vDTs2Pia49LydiEmDju
/rDbAFyLFcwsoNuq+vqFkZLyfi2wBAVlAAf/ou/7WXNM68tkvazORRH/wmv+ZS9Q
6V5sgJ518rkrzsybZyt7PXcWV0OJuXrFvdS3hwNoD0W1AV7h/wV4Evq9vtu4mvFm
8gEi34aalKwzlsJNeIppBVdkHY0x1w4H5iipWwbLH4obo15e2AXxtcL7IP2AdUEb
fsXbbO3ZRq17kEfkc4wjXTGcFQsnkXn1IdQFLY+TigbhDRSFCbe4A46J64v68kts
rZdLRVaNZaVPdzAA2IyYAS4wGWiDlv48U9fY6kTyLqAV18WpWAAwDk2WzB70FYMo
yGTkHz4KsaXBeofjlsnK9dX0xl7QbFWeZdVQwW8e+8t/ozhA4vjAHYTAQxIA0is6
e9Yx2Yw1tuv6efaYHdZkNv4LCDOMOuU0JvrIatcATkLSQq0/Xv7ozZgACveK6VNW
8Na57XC/DcNbitUery/5U/YFuGBy5tPXNmcD4UOzmKW6Zv2tIvpodmXYAfeYea0i
mNSjAXMZuQFsZTuLsuk7dtdf9AHh4N3HKL2Vu5QJxD3JAF4Bq0bxQgSPSjz4vaL6
XS4QwlEGd2KLcd2AaJQemgC9VA7l8NnRqysAioA7sqTGc10BoxAZyoFYfnMcP6tJ
XTG7UEzel3APx72v8W8UCfES71X0qbv/YK+P4BPIykmoVin1t0THD66AhB6ZLTpD
b8Y7WbgBc7feejaZ6z7uxag/VC+ahVkow2P+J/cTJvQ7LB1/oYzp6PFF0/iFRDiA
plxXrfQ46S5Oz9n1sl/FjyAWFrm/xi7kRsdz4+q1PvOPZ1walgDSp5OpsGyh8O2O
nniZUfJleaz7EuWRcNn3WUMD4cQElWNT4PaDr6N0AoFksiOv1zEZr2+94kiwk0Bx
RE+6rp4DPy0Ea/3RBI1wggzWBK/i6pU/nW9Uq/jLXxDlmSBuoOAZmckbdu1yJ6ZT
LwZGJiGhoaKVA7xLtCEuHbO68BXqj7BghapnMEcZk5W4gtE5P0z5MUFBIVAU7Tx0
HjFFFg7EDcEObwK6ooXCCklrfhN8VEMG2hNEwvMS7IavqgNS2w/sm83HtUbuRLh4
JzQJcCCP7zfwYW+GTc9M2y0IcJvbg2RTcFpkgx674HE2jFOl46ZGD2DRQZoH6ei0
`pragma protect end_protected
