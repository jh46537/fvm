��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�^��h�����mb��feE���0�8GI\�VE�|E�T	dݹ._lR<���<ߵ]�uj�x i�/���r��Eg�佗`Ҿsb!`�ĤF���u�#@���}�;(Ԡ7K�#Yo|B�&N�	n �*�3RR�gz��eO�a3(��Rmʬ���e��v��3Yt,�k_�#G�:�'��b��gd9x�,�T��ƶn��o$���~�|���y���'�t(�PXD�5x�w��-���X�5���'v�\<��rm�~�wHM�\*j>g��?$��D����vǹ���)'����*x8�!n�����B[P>���,�S׌1��Z��(gh��Ws[�a�do� 6Qup�CRړ�+���?<w�B�*�ۍL�X�y؛LxH���tT_���/�Tj0��!�0a�rngMX����J�R��$�axi�žw���ۡ16���]DǷO.Ϛ�����D[���ϛqˏ�SԅX_��z�M��j�;}T�Ё��B���aA�r^�i�o�g^.��(}�����]$R��!���^R+jg�˥��Y�.��}��p0��wo�~G�ˡ���L�uK�i��r�MkB�WR�=\��#=��L-Bw7a��ĥeZM*�v=�N��[?L��v��#�?�H�y󻥤�V'�,���̿C�P��[ ڳ��WV��H4ڳ6�eM�\�TSVC���E/Es.��H�1E��$L�Y̓��%d{�~���E'*��l5�P��� 
[qd��Yx��B��T��W�{?p���H��h����	�	0I(8���s�a'�ۿ�,�y�BDh�БFT��������D���D�B|�gب����ũ���r�u�'-( Ϥ�?�r����w*��sf}�lZ�`�2����4Fo�-Um�C����������KL�p���G6��%�I,�C��,V��7��
-+L(�v�1Z�A$Ԭ���Ƶ�ԁ����#�1�V(��lڡ�B�w��8ja}Hڢ�<Yu���_r�wA�9K�M����/�w1%����n�#o�w�(vŽ_i�,��] ��SsUQY�MG,��hN�f���q�[}�?�R������|��/�t�X���$�sC�� ��>�fH���`��i}"hѧT�;�9��O:#���u)s7���^��i]������-ok-O��X���1Q��C�,21��D�KӒ�e���9,��2��$���YxV��C]����}���I��%�3x�~k��}�Џ�53R�=��J탱c�����uΔ?�����{�Irg��p���͔2�Ǎr�U2q>�A�"u��j�P-�Y���b��c�BU�=iV�R!�IⅦ޷;�K�qf��\2{�Q�ȅ�y�sI�;��{d˼�Iu�{�e��n�\���[�/G&O��k����F�!�ˁI��w�}7��[����: �b�= �S`;_�Vr�Vs8/�L_�K �]������X>�'Z� xDձ��������Ň\.�J��Yf)j-(��uJ3�z�2f�[.���&|�,nT��e�#��%]��?t������"e�n����E�XmCbO���IC�()���>�oy+`LM5}Z���&�U[ܬF��Zc�Z�\Of���[Ń���l�����EK���~ѧ �RЊ��9P&�o+�l[ޑ����	(����X�&qd�C�C�s�k�!�3{$be�7?��3���u�Rt_	��6������UD�0t�HP�����i0��s�=S���H%0��F9E��_y���J�	m�tK����2���a�hw'���R2�zTJ����QԨ��㰒m8��v�+��RW����-`']k���U������<��T�:������y�6B�[k�;7|~�|�NxcXy�k�^�����E&���r�f����$-L߇~��+9]#U��>�T�?�������!���! +� �e޴���n�]�2��T%�1�Q9xè��o>�u��]�F�\3��8��"���+���ص��B��z���6R!�?pŋ�3y��e���S6jڰ~��J�Urul\!PO%�n!cm���� 2a-�)}>O�0������d�[#�k� 7�Rg����)��_[^��R@�������{ߔ��Hڿ��WT�^tr�_������^)�0}O W��B������)��׼IK�J���F��|�!cEzq��o��рB�˃�⡈��dջ��J`�]���p/�����3�H��$��n�����w��i��~���MG��T���ETTM���]���o��]���\Ϲ` ?{?�ܳ�(!�0坐y�d�OҶ��b�B�жj
/�������]��ս�s3�sw�$�,[�!s�Wo��f��j�!�7��%6��i|hǦ)55LU�j�eB�L�9�5)�]�����m�C|��x��m^ *7P�=}	n���QyS�ՎiM.�n�- 7V��#�M�
�������;�r�,K���}�p�j�_1=$��� �E�K/_"�Ǐgjd%xX�&��'Jś2�z���X�r�>��l|G�;� -7�C��;�0s�����~�C���ʻA�E�!��q�"A��Z>[�P7啨��0K���f���A��p��ǈ��P1����k��u�sj�B@�@��z�����1�kJ�wgtE&E7�]�Ą�-O��ht��@�M"b �T>�W��)�qYV��ȱ]��~m鿱Q�?9KF:���s��>�ޕ��]��DWX�*�cw�%(�Bw��Y`���-,c�!�j(�����F8,	���cu����h[���.(�J}Yz2T��>FU�Gא�^��u¯���+�X�dw0�.�K����W4�'�\�q��i ��'��#G����|sf�Y��m�p����&��\?:���) P��5S�p��p���D��S���dpɱ ���t�U�+�/��u'�R	ٶ3�K� �����k����0�r�ʿgd�V�jqT�0j����vvy	���
}�

��<��l��>��"G�$� �w�����8��؎I�Kh[��� X�JP�c���⢎D7 ���F��V�?�ۏa,0h��:�v�� �ƅ8�K
  &��w{W�I�̘]sp�'����^�x�i��^0���n	���='�;}�S�z�}�3���lj��.(?E4��*���5��
�u9]��l��Ӯ ��Jx�!�;I��Z�.��}��;t��ŉ����YM�܁@�축%�$s���St|�*{i�I��!�ɬ���%���s\x�Г�3��Z�*���)-��O��Gh����B�5W��l�}������)�~Y��ԡy��Ѓ�r���'������%��ԕlV`Ը|�5�o��1����m��G��O5��1Ԇ��������Q��#�`�dR��OS ����|�s�$����/S%�T��Q	
�\�ǈz:�n~�=͗��x��wZ ��Ɏ�K��B#m0y{{�A��j89�G��z�$w;��pA��Ka_&o��O<m�|84��mi��B�/u�QC�]�ّl��B0 ��ϧz�yC!з�-�/ ;�b2J(O�=����yX�Y����d�uX`W��5���Nב�e�\芀	c!�tN1/0�cQ�핢�O����Ҏa�(UW/�J=���*ӈA1��N=�0������E�Rr�I������W�~K�1B7n"}�����D#Z�G�/Eˈ�쑭R�u|E���N��X�.:g��(��%��I�FP���~�n�,J����K�������3	u�q�z�JD%�=�S�>�X��M���4ԗ
�Q x�q��y��/+���gxH�^yqE�)u{D��m.��)�R�#�k}GY����}�͊ݹWoS�I��vK�z��2+ˬ�v�3��(�����L��CZ��v���x�����u��#��()D�my�`.AY�&�Ԯ�X����<tx$�K�Xw�����^�a�>�l㵱/(��4G�����C��J���q�F�3���c�T�w
D c��ud��V�-�ѻbT�F)C�Ϧۑ�ßg|2��&��ǂ��������̌�ڔ�1@��)=��t!�>W,���;Fe��F��v<�ř&���ٞ0��ŮԴqЪ��g-$WdF�˺����9��PVҵ�������2p��v�Y�7P
�R+��xk���P�$ފ���B;�\]"�J����,/��|�j��B>�s����c�{�����"T:���Į�������Ȥ�~W�W^�D�\�^�s��,���4b2��.��6x���To�ƭ���I���I�a5�k"dB����bxG(��fi�U�|2��v��� }!�vP���9�^���Hxuh�w�-�������+���"��*䛻�g�}8R�L���S���B�F�E���
�2Y�����A��x�a���������Mx:�M�?�j�KDJ�a�XL�X,[�A�Z��!c�I��y��oP�q�  ��6� x���J2�ZPd,���9�
�es}+�~�@��x��*.�X���y|�jB���z�͒:���?0��ʣ T�F8GS�(��q~��^Za��x@�����_��y�3Y[8���0�L�� q��'�XlL��7#���B�|�Y�^��HZ�!s��Z}&�Z����2!���i��M���-7e|�.�f#�e�VϷ� ���4�{LN���K�#��;�ٷp�e��7b ��ѳ}f�4,����V�gO�?�U.xT9�p�)��?��K����0Dv.��n�2��^��׺>B��u���l�J�P��k��s�u�:V�,����L�����쪺ڿG[�Ζ�hA �2f���/��f�������N�:R>�1�>XIؿ{�r����7���0�4}����8�m���f�lUFO�X��J����u�/��jŏZ`h
~�!���DLj�yxP��(q�[z��h�
�X��0��[F��O3YzL
�I@J~��_`����A�Lҷ�X�{�=Lz��U*��u�Ka��z��] `a�4e�/?8�������#�ؑ�٧t��<�V��%����|mx��3�d4k�y*��1ƭOZ��*7��O����&A�'5˖��'�eJf4�����:).Z��.l7������'�����B�0����!��QA!s1�Qn�?e�����i�ъo9��O�}`BM1�R�)�^$��E�R����{pN)�	xu/]EO��	|n^�'&��"�1t�m.��*�*2A
V��p���\$D�-'�J̗b�z=���*��C�0r^*2�Q�i��4:���=���i8rݺ||�=����>�P���QE�J��
��#2�RI�y��xE���.y��E�)Sc�[��i"��l�?����c'�?�����uU���M�@��N��N��o̢P������U�T g�xQԗ�,6	��{��&Aw<�����fV�c����QM���h��w���yA�*>	OXJ�Oq�}'����$A��&b&�=F�#��1EQ��JF��p�%U����I��F����y+i����Vx�J(���'>GD(�^�\Uq
�Ϭ?�sj�z �N�%
:	m'��{d7��
�|dS��]����qp�ѣ2�����F5�&�{U!2ZrU~���
�eH�E�EѸ�� Rm�`+jwӋ�b��E���EC��G��F��򁯪s�鋺�w	t��Ϝ)�~�W�����"��g����v�QT*9�%N�iIW�5�u�WE��b��q�������ITyzf!����o�@uR��y���z��������*ܰ[ZχGU�?����4m��'��m@�����?2����O""w��vC�ND�$�cl=i�ݱQ�ӪX3kc���N�k���}��npN���Y�e8��O�G������kG���%�pL��3�B���_�LS_�4E�t闽U��d�}��Aa��t���Bh�z��(T�Ω_�XҤ*�G���st����A��&��������f6�.T[d�����'�u"4<�Q���ɝ5�$t*Y_��:��M`�\;�0 ��u'o]!+E,\���}�Q��Z��(<�3{��q�+ɹ��lK�q��e�.ɬUE���,��q�:��ȕ�D���"~��{+�j����"�`��:�X�3&�<|0���{W�;�i*�3�jv�����SP:���h�����<v�����e-r�H|�q�Yn�ʔ��2`��x&�e�1����m_������m!a�Q��{�	iw��~[� f��ǋ���ӟ�N���ִ��@����bQ��N:���z������g+c3 ��0ЈWR"/���,>y:X[uX�{�Gu~GO א�����u�u����B"@��c|�0c���|�-�é�V���c�[�!=ɔD��/�-ң"b�����K�>>h���Hy��\�����lGQ4�^+���~X�#J8E�g��9��@6n\_���V��nt��]]_E��L�+:�$P4 �t @4lZ�2Lq��$�pلf��8p�K��ãc$����v�5�5�isᢇ.7�oՍ�M=f�GVymJ�(��Gw�B�>Q�=M�8(?�QB��V�.�qa��*yZY���Wʾ��+�B8�ρ�j,����/V����Vz:T[�����q%
�Q��A&Ԑ�mK�ގDGU�e���?܈��yV�b:a�.�j���B��bStH,4Q33���Vv~R��O��[��1`�"�Ec) �r�H�Q��?\8�`�U(l����&�&b��p��/I�s����$�;�UGj��3A���!�7��>*�LM�o6^�['4=�D����1zЌ��`|���� �Fu}�8!�8`����r8����X�R��hؠ0y�P�i���l����J6G��x�&ܴ���$�Al�.^T�~M����$`-�eNJ� l}��R�|_�����m�&��_b�����$x�j	���<��W>i�'��!��E��՟�����S������e�I���W��z�AR�pp�.j{iᭇډQ�4V���i��M 9�hnB�����
h�S�p��PI�hS恽���508	�*9(;��{?Y��2W��7"q>�:�7�����rruu[ c���j������xC $��d@~!?�ćhL�v^�T�_q��9Ŗ��v�)?.�Ї31��4?|Y��$G�3���DBO 1�jB�P��?�cg	T'��\g�>�`
�c�w�Ԧ��b�,�j��&g8��h��wC@a��wۉ�[�uLg�%�ůx+G�A(��e���kD�e�߫&	��#����Fa��=�Z��}yx<���߰�M���4>2|ch��&`�*+ve ��|�ݠ��>�>�����T��p��v����vf%�o�7��Hs�pDw�ܣ.��&2L�����b�L�;o�ewK7w}ը��x��3Ɩ"$m@m�j�������N	P�R�\��dZk����Ҿ�@��oÅ�*��&O�EROAٱI�����\��'ơׅ'D ��OcT��{����^��綩@�P�"=��S�r-�q����H�0u�'��c��6��d��3�� �����'!�c���;X��YrU*u���)0�ժ|rlʦ��G�vk�Ny�H����7Sz�!܁$���5��{�G��xwBu�b�-��Ap��e�L��.m�aÑ����Pr�}��(�U� ����qCe돵f�o꪿�o��s�&bL08�1c˓8�T�1��M�\왩�����M��7:㘁@�&��&�J̞Z�}9��dr.dО��)OD�{�u���Y���9�Ĭ�]='�ó?�z��ʟm}�-��!Y:4�>m���q���9�yP�.��L�	�on���p8&��h�� �`���%K����A���ͅ GO��2��πA�3�"W���-cE�u�G>��ܰ~o0�M.[& 5���8���)\��a�W�3K��"���fT�xF߁힘�Z5��!3)����4쌵�Xm-b��l�=�6�+��F��4�^���%�o��3���.�(Rq��3{*W|�m�@̵"�4�XSePB9��~R�v��"����j�&2�=*��8E!LLkw�h�B-��^��ׇl`W)�YE�щ(�j�I����� @<>ߣR?��s:�ԛ�}�$Z��h��@��>�0eR�X�B�ۚ�Pg�Lxs4gSC�%W�>��Ã��Ȧ�g�HZJv-0��T�^)E^�vZ�39te8�gz�5�@��*�m�op��=�П�=����Բ-�j':����(9��-�m���]�sN�8I����<�O0H5���7�!mq�`��,��-6�}�nU��� Q���$���30mA����ǲz��_��� �<ɂ1�3�8�8%��
���\7�R��C������m~���2�byk3ᆇH�X��E�&	n��P��'^1�lF�T�3�=���ὖ��YGXC�|z�m��	[�$�e��w\S����	hҎ-��i�M����d�Ҩ;���Q`�X\l������h�s�`(���{mN�?�b�6��i����\��v�\���,2խc�J�p��g���HdH���}��t͒7����}��2�+-���Cq�����P�&�v��fjl��ߤ��F��_r�M� ��bG��* hX������Ņ��"��V�R~]�r�NZwv�q�av�`��g?{KHHk�c+�^I�s'�����w!F�X�&FK-w۾߽^]f�lM� Ÿb���xgW��2����¬��g1�|Xe�9�q���h��nUa��{ʮ�A�$�Yp�>��f�o"O!�s&����� �f�,7�	\�̡.u�ƒ�>��Z����;���U�d�<�Q|�X�W�)'(�H�YP�� p�.G�l���ɉ���o�&�h�[�J�X�n���<���8�T��ܭ��KA�XNӘ'�=��h��5Y��t[�{B��:�V��8~���)dz@�6��}#�S��4�]P�&�UA1u����6�N=�PW�8����U���m{_OP�j��ci>�4P��8g�1�sɺiT������,�9|�4���Ncf��ִ��Old�s����y|��x��?���&�����ц���2b��M��+Y:}�����ǁ�]����oF�I�F�	�d����W ֹ�����q�M-�)�A!���R�w�}9?F(v��LT���Z׊r5�C�a��G�-�!�)z��
<���"����a�h`ս��-�aN�|���1�8dس�w�L�5����������@}���@v�&������+G*xӋ���~;�u]@L��5�6��*�u�	�[��>�_x+)IV�Eب*��u��r�Lg5�@GQ��v%i���r`���M`x����0� � S����5!ݟy��^wp�=Ź�ܙ���&�$�4}~ "傭}�.=����y��'FFy�����uK	��a����	;,��~�i=2I�SWv^�"Zֱ$�*��Y����>�^�`lYS�`3�&�urc�"���1�b�!�\�n��@9~%�ɦ tJ��&��a��8��D"V���~�/���qj��ӟ��Q ���
,ǐ��N���%������\�ɭq&XB#�j{E�@�Ƚ�I��%sn�]�]���y�Bd ^3�6��X���z�sb�^�-(��@���)��jt)��bfp�:�1�Z	0oV�j߹饘6��r���������A�_?~�<_����c�p�*�
��g�(}�k@�/~q��V0�^�I��ŨV�.���,�^јb�Z���~�®�O�[[�GU�o]�q��4�i"��w�����q�.ڭ�Y)x���|��Ԭb�;��� r�5o��ސG间��:�x�H�D~Gq
Yc3҈d��W#mߣ��<�d�e\�Zf��֕
9k�K`��b����#`��]�X��њf�D��M�rlrOB	�B_�_
�
Qf��<@��ig���լ��,���}��h
E���� �9�] �K��{2��t����/%�W�][+ 9*��K$~'sE�t��>}�D����Uޏ���� Mc��8E��O���#@?��B|�X�_�m/X�/��8�"F�΋�\�:PA
b�4���2���Q@�r�r��m`�ܻ��Y��S.���	I�w�w�kh�N$��>w!ь:���

Sp�
�!��iSϜ�����-��ɮ��m���/v��Q���剘f(y��Q��<��R4�0 Q
�ޘ�D9�����M����/پ��X�見2�.��f�I����A��= Y���P$�_�pț��,�̃�a���"69�'��q�,D^�5���<�Ү�q��gܔʦ�Y���r[���ApCS�����!����F���}R�5���z��eB|�����Y
]dP���2�sе���zP�/"�=o�vb�U�ŷ#D�	���vz��S&��@��Ȗ�a�+�#t�3��H�bf�qc&B<�k����SaF��Q��b�!���'";��ۣ?u-��u3����b�@ %9H�k����J�a��r��7���bsO�l��W;W��{�� Ԣc|�w��b�F�L����d��뢛�z��<Б��#)2��o��c�FA�Ŗ+oD��,�WN�j�i"}d���{�klM�7E��11�U@D#e��#;��(��H�q=i�d� o!Q�L��ة:���IH
�����l{۹�5Bh���om]��� 5z�%�����n��Z����#�����On�	��pt���p��O�r�Lh�����Wf�,��t��F�z��Clz�N ƹ}|L!�[���v&T�'�{�Y8���T.�qyY�DL�bJ]xN��7���ݾ��3e,�́����g��ۡy����ks��#��ˎ���eG9W���_sfX�f�� �z�����|v�S��2^U���j�����?H��*.J�jԨ{D��x����6�+�9���c=�/�hvŒ����N�I��	�|�\ �^-Y��:��W���k��D�_��`�ǯ�ҿ�oU](�A�U��S���C�mkN~�1�ƞ�y��1�]�~k�,�5q�l,�`L�r�����FD����u��Ψ�a'�I�D����r�G!����F@��q�H�B�ЦA��K=�'�8yc��..�7�<���<Jtߓ�(Z�҆��[I��d���_z�뎁䍕�3�R%2<6���OXw�r�JY�r<���l�ޣ
��HK�9�Y*a4��藌N�pw~i�q0����kO�����)^�=$�w�l��z�X����%{N��EΝ��M��^(�*�4$�a�D�	�He�*O�7<������Զ萻�� ��bjyJ�U��6B�������ҁ��s���O���f�&����C�!}����:�e����'_Iu*��Cr1za��̊�\��Xj9�p�(�^ӡ�o�tT��q�:� R�N"���uD��,j.����}���2��Ny��.���<4��#��'�1�,՗��pRf��8���K@����̹g�.���eo'��|��I��qRo���ՁP�P�ZX��uR�6���J�%�bd0�<��ε���iA�HU ��u��S��B��'nj�_��Fr�[C���oi��4��� ��/�!* CZ�wn12��M������	��Fߗ�\�h=��V/ؕ�Rg1��Y��[QA���g&g�q�`es~Xm�Q�+1�f�3S�P����N"l��s��t=9 ��Jۛ�(�8I\H�))I3�B������Y-���.;�Q�q��~%�[������3U[F��u�`'��z��\���0C�E�p�F��|g��{�����wu��5�(#,�Ĉ����*��OY�ɤӭ�t<���]�S���~B�1�1*������K��eO�z�i#)Xҭݢ���p~pJ��=��T�q��O����X82��L��߄��ӫ5:�HV��jzІ�P���j�hoBp�obV6��b�W��yyV=U!�阍m$|��ӝG���K���ߟ�\��?.���D�~ȵ׾���tj�ͱ'�_qgy��Z|$\wWV��������T����+?��w��0劬�Y����o�M�8�wLhXQ"�|�_�����>/D��>�ohk���*0⍧�^�.�ĺN���)���Oq\L�.����#�du���l��Mó�q��tYRnR�XSȲ��(�V���ȁt�h�Z*�����F{1�9˹���'?vhP��T�Q��B�C�,�l�&j* �풱�M0W������e�v:l+��q��/�9qM����!o5�����U~c>���l��C�ADx��V�u�[8�L����+`��SؗN�GY�����1�H�0��**�s�ok�JM4T-ɫ'o�%�� �
��K����:z�K}�՛̤s��K�����	7m|�#gk)=��Z�оg"d�.��N�0ԧl�z�-Q�Vid6i��r�r�N�����y[���p5!(v¾�X2S+l�.y\`(��T���^����pӍ�ԉ��<%���z7���x�.�kD�A$Fo1�k��G (Ы복ʚb��-��_N�X��-c�O���{T����ʋ/�I%����$����v�b�fd,+O��\bݶ�$Z���+���aٹK�'�ks�k[ʃN�g��}��(��̈BjdQ�3gH�N�]<�c���yC	u�Iձ� _�@M19��oW&���N!1�iJ�q傎F�S[�=FO����kn��jp�C�(t�(�L��H���+7�%~1j��@WS��� e��>�y���9�!p��Uv���m�������C��t5�B������dwRIᙖ�KM����A!,�W���"%_�ls�K��������XH�h'���ڊ�{J�۱��~�wb�Z�
�s��t�G$y��z�B=�Z
F*�)������J��h	1���ԏ�����׽Bt�`��dE�Wt	�Ҕ�0�%��,���K���j�%�D��z� �+��L���gq~����D ��e�zR˟���G�}�l��0U��(״J�0�B A�?b���'�[?��$������vq�����(�ZF�+v�8|�2��j�㘌�0���l�X$]��3/�^�ߏam��s���2�����[`K�U�0�xQ�!��/F^�����z�����&�T&�gP��a$<~�ei�YX�����M�@'��F��vf�1_�G���=������{>M��C��*.5�sv�=��~&��O�O_4�f��F"�2䰏s5��5�`�Y�ZR��=���K�,9ڟ�B=���J�I�CM�L�6YQ��N +o�8NV�*N�a'6zQPU�3n�W�3�v� V,���ί'�����y��"�1���v?XE����+�H�@�7����o�5Ց1
�!�n�m���u�N}���.��>������.G��t��&C��,�(=�9ڀ�z�B��ܭ��{rp�#�.��[�����o��>v�y�Ԣ?�n��Ś��H+S�;��H�6z��)��0���-��=@�A��g���0il*0	M�NH-�#ۆs�]*Hd���߯>�(5����l!"��Oë��Ly�pe��X�e{����K�GkU�Z�t:�+���Cg�:'���`A�]�<5����6ޅʊ�5Π��yԟ���._>�+�*�YQ.c�Rl��,�Iz׉��Ԁ�m�S��LHC�>��ïh�h���O��tdl�>���)^�*>>�C�Y�`Ih8�N�;��U�!��-cOtF�C�c���<As�)mqo�<w���cu�Q�Ͱ|�l>��'��ȋg�Ҹ����C��1�a[M���+ Oj���%>�'�D �u���.d���a�b�ED:��+�����uqӌl�x2c��)u%X��J،w�nl��{��rv��lGu���h���Z(]~� =�3�e\9�vm���f�H �N��E�1�+����Ӗ%_���'�`d�2��R��ԎS<�˄f�,�����T̉��q��8����8�&��;M��wgѪ/��=)+,�-=�N���l�"#�������@�}�`��"��@�>�%�g���B�8`4�[~�"�R��h�̳�5%�Yc��L�1�-����q�PP[�&��ێ+
�w��9=�`Rf�܎Wk���e���Q���-�s��-�bdf��.{:��c}K�M�7`��O��@ߖ���A[�qN��>",f�BE˽��U��r��`ާx�C����G(���4"<ǈ��CC���z��Y�R��x�+##XfUD�|s4�]�D�/h��3t�M�H�K�y�"AqNEB;.
�4Ύ-R+3���9g1c�^[{�pʶb�N�(��-L�x��Q��b�=��"5� ��ġ��^��}���C���jΟ:Z5�2ˤ�LM%E��'��%_�P��!�+h�.Z�8*����N1��
w������#Z�h��9��ƃbʽ39B��~�:�H�� T�}&<���+��)z
�מE`	���u2q|��=��b�"Z�ʩt��ҨY����Al8X"2mRQD�c���ұ.j�Hr� ��ɮ$Ŵ��Bz�Ѐk�٩�;	0�d�5�V|pQ�<ԢX�db��o���{/��|����>~P@:��x7�]��j}�g]#'4��0�3+���3m	i_^J�T��_���CN���n�A?VZ=� �S����R��tG|��]��@1���{�"��z=������W��,�!)����&���:.�P��������-u��:�s�G�@�#�.������OB��@�Tf9�gm���?ʈ46��?�U��4I.od�6�up R�rVQ��]|-X�|ط�< �A$͌����F�T�d�M`�&�)����*�Q/��F2��x�o�o��Z:i��v�n��Z�S����]a&���� ����^Jd!6rX�8� 1
�j2Qc�P�3�QN�t�.Ŏ`��5R[\�z=�t|2J!����6b:��ٮk�Be�=�+63K������Ĝ���	5����D<�<:wp5tE��0r yT9=�^��y����@��|��6���ʷ�ޥFk��b.� ����r]��H),�d8�.��"��֜�`�z�o�jF�6jP�V��ZV������-������!_�l�1�sF\��k���l�<��5)�6�f��A�q��Y��Id����ud��\Oi�{���􂺡de��%Α�vn���S����7C��2%�i��p��,�!�{������d8��wB�}��d<; 8����<��fA�,{d%��3�-	TA-��zck�/N��"_�%#��T��j.\���@�!ͧc�K�G>�H-,�F�Dn�^������-��Rn%���wk iۯT�v������ �/�A7�f�*�ϔ�p�&��\��1ږIy������P�$�o��3�!]���x8�/}]�2ǻm(
;d%�Tg)例C�E	Z�/+��U��e��x�4qBA)fH0Y%�o�Ԃ���mX��I��b�qϴ�۹3v�{x.@��T&�+�x��B0�r�=�H�q��7����:�@�� &��^>d�KN3u80K5w{Ii�h�����)3��ʆbd��ng�=��\�|Wvc;�|����|�����U���yܞ;V�~���NW/*�K~r~a���*�Ɩ���ȓV��p��~��r�rܝ�F8M���z��X��?��qJ ?8`��a8"i,۶ Q	*��D���]i�j�|��{��>�RjG�i�����`+��~�iy��y��/�#�3��;C�`-	�^ӯ� W�BW-$K۴���b�VT�^�-�6�y�W�Ԭ����"sqX����>A�pL��r�N�?���۴�"�V���j_{g�;̂��RËW���Xa�j�~2�_ӛ�v�@�z��y{�����j�ݡ5���~
�mC܅�ik��7����@�$�Po��|pT��Z(Ν��8�%q����1��zX�M|CXE�eau����;Ka�ɼ �l�Ґ<b8P�3�oe�+\ݦ-����q><��c�S�f��fӾ�4�l�@A�=[��z��x�u�adB��ں�e�\��m6��7_�mfص�3��b7�>y>�ݘ��+���N�-�hg��.�W��� *�Aj��f��F��k�K�"9&ɬ����l��0o�_��,������p��X�Źtk���Jaq���؏h�D9���9�%`�6�dr-i��}���5s�C�����u��t��O\b^�����3Z"E{fk�X�j��H!F0���U�v֤5U��k~;�|��l6(J2=�z��<�-��be*��8� #��&d@`/��I�vm��g�%�;렯U�-���,M�7����Zy�xi��)QS]'O��g�4�ɭ��xX%�j�&�\!�}���>E�d����볶�D����}7��.�&���*g����RG��ME��:�]�����GMtm�;%��ҩ��-�`[��J�o%��0@j�Al�"�<$f
��n͢4�q��e��D0.E�C�_Ĭ�&�h����(p��ZNSۀ�\���*
v�bӠ^��c�W#��x���gFW�f��j�[X��a�8���`���:�}2[����+~57E���Υ�x�]m����^^.1�^��o��N���Y�ѱZLwc8aI|�x͉H &l��\� ��d{������6�%��H[8�6R���I���Y�@J�p��> �5���$���I�
&p�[���0~��3�g��@ӄ&�6��I<4&����͸�ؐQ�i���D��ofMQ���'v���Fc��O
]y�
ժK�A8��B_�%��rG������W��;����!�}|�������&*�SX$�_�����b�"n9m�^�$;$~�~�I{7)��9Z���y���gn��f�>���X���4��NRJS��wu��6\K�<<r�RT�P^aY؟ �<�A� H(���و5Z��R����Du�W{�.g��Ǉ�ki�쟼�w�3�Ow�����<$�Cf�Ҋq��6� �g)6f�&E y_Ya�O��t�Ax���=ѧ(�6���Y�2'FzM.p�+D�
�v|F� ,>9`sTD��&�����l�#<�����K}��M.����:ܗ�fp�.�Q�l[��,s�MP��LY��88�5η)r��[9h�Ɛ9=a:�<�"�I-+-<|�YRP�F33,�̴����� r��@?�w��,o�К2�@%���U!D�B	%�d�ܹ[�Ĭ1����4�\u�e.�����AOAw�#��-S���.]����(h1���bK���ߩI&ꤛ���۫.#h�	�m�8WO���lͅF̛�o'�/i����v��lq�v�v���9���I!B�1�����ew�O���f�E�	�K����1���X��^���u2�g/�ȕ1�>^u
X綑��Z�²���(��4�%=�C�8�0P� ����i�9���Ȱ =��^�#sؒ�
Ą�?T�)QxS��+��h���������P����6��s����<�+�U�
êt������ٱj;S���zV;P����?�8��|�3��H��@Gf���m�����
�=���CM�-��Ȕ�+�#vZ#"�+,��<����N��fd�ol���%��7)Q� ��^(I��!��Y�].3 Z��pΙ^��M��Z���&��}a�v�R=Z֕X�Ӛc���l�8h
��L��O�\��K�xּ���σ.�Ҵ�����QtX��Ft[^�o[բk��!j�ŧWr�\}�c���Z�a�x�?�ATHsYL��QT�=��9��2cj�y!9�#{k��A(�:��8
��K��B�����K�0�w���'�r�U!
(�����y�������A2 �-�㰦>�MV�6"͋��:p}�aWi�#2���.� �V���	xN�rj��������
턺X�t�#P0�V��E9wT��Sc#�1j�=��-�4��U�.m�;~w��:ۂܢ��Аށ��f�`g�bJ��A�;�]����U�Y�b��q'�Q"����`v���Y�m]��؎���;���V�8�NtUJ=��W'��� ��N�p�&]�KBig~�j�_1�خ��#��?�l��jg򸽱%���(����vy��>!���+�!:�'�U���	S�y�M����ȑ�v���b���l2i>���+��"�m!��*���8��2x_rЖ�ug�M�#�(�<v}�41P��Ä�h��>ɭ�H��k!z��?����9
�`JȆ%��z��@)�gT�)눽Z
}vg�Zs���t�ybCM�;��w��ۉ��ς���`<�-+S�PV���MU�M�fa��9�)W&6�T��ήM~���0�p�mvV���C���N@����A��)*��Sd�^W�M Hӿ-M@��F��l�x��p�:O�l���p�6�,\ڡm��g����x�Oj����4p
���
�N��c���sE(#4��%P���12������ ���F�}�O?
L1�H�NAg�1����l��{-'����/*�������M��&}A��g�����H��t��υ��P�}R~ܒs����Z`��r��Z�ku��K�=�b1�M�/cV��f��j����j�����UХL�l�u
���:���K^�A�>�I@j��(�ͪ$Q[�̚��5#Uz��H���˦��	��k���!����?��
�T��w�uM�t$H_��)
%z�ݲ�x�LY1�h��Ψ=+ʽ�I&� c'}Qo�J)I��.��D�u�짩#wm�q��-�I��U�R���H����.~������
�U�2�X��8��2©�O��-�����H	�[O�����#0�+_���R�ܩ�����6
-$�%mX6�.��9l��ܜTm�m�{G��2��ל��Ӫ�K�e�E�@����9��b�>�_L�����$ �i��1\����]�'qf�~�÷=�&�k�4�5�MIiƤijy��d��R�#�0ﳎ4q/�t����oʬZ�+��8;���}I@�n�qhx�i�W��'t��^f�PM��Mr[��kYt!�:z�U�"/�,*�ˤL[�������"&A:��+g�<��>�3�9���������-��c�6��N0,xş�k�y�чEl|�YJ���\�������@� �M���D?x�F{\�G
}���i?f��s�5{�������'A7�}*�ȋ�H��ݾ?��]�(��Ր�����S��œHy�w�"y�ӈ�}�@hp���������j",�r�陂�Э;��)�ʆ��J10��;�e��lT)��A|�V���x(����E���o!b8��دMJV� ��������i��-�`v?����16��Hv8 B��v636�j�P��/�VPB�-7+$�YΤ�{я�_'���Lm/i�]��P�K����]�c�T/�ƽ6�5�*�C��aC��sI�;ϮN��/��޹Vl�#��A���y�K�^��+w##/�гD7{fǏ��_C��:��!b��m����zn]=��6 c��F��04j����S�I>z�DޒO9��4�T���Ƅ1'g�{����<�؎6ҷmF�'�#a9�B䓚MD�����<��]���?����*8YI�����8%�L�^�m+�GJ;�1�-H[b�������K�﯁Z��.e#N�t�A}���#�r��n�UK���?>������YBLɬh�Qy����" �ܴ�.��<v��o��HX���t.�m"��һ�.K��p)��K:���32����pq��߈sF��0��b�<��S2�6�X* |x��Q�|���.��4Q��>��%�$�r�Ca��KdA�����p��m�֯ʠ����Ѯ��7 ��
6�:�����PN����Ƕ|���m-W�{��}=Ċd=�>LH��)�*�<p2��`�QW`����IV8vD�����Ǖ]�e5mp���>A���:2�3x�.�=�Z�S�]׌s���SϛW�����D��Ī�ߝ�"��Ps�ڛ�*�ԉ P�]�}�v�J?;9QȄ1���ozȹh�Ye;��j����&2�CaB�(��)�(D�M[^�I��-jCy�v$�Z��JY�L�6��@}�F�Fa��}�ex�:Ic/�@Ś��m��(O�M��z��/�X�&$S�!������+�Lx"��fc�_���ِ�:��6����S��\V�t;I��� Dt�?�ȃRgnꝍ�nzi�x.����TrB�9���r��k�ss(�h�}d& �����.�_�)�n���=!��^�c�;�-g��Q{^�l�Ё7@Q�8�n�V��!��p>V��B$JId��)�yE��Ќ�<mix�5'a�𕪫��P���etW��x4�oA��r��)��" +��j�>oiI��ғ�.�7N��Z�?�D�J�M�y#�8�R�B'�c�f`�ߞg���ߵ�B�c�aK�t�YK?�������p��3_ſ{�iA���6�� ���ݥ��l����O��O�M΄����l� W��zP4Y������J�0�@˔̭��<���B�>J��H+�P�VlI38hѩw����3 ���r�`��*�'z��#��v�@R���I)Dxy$jp{�&^H1	��������(�D��I�����+���.z�.Nz�X�
��#�;fܪ�6�p�qg�-Ϙkn~��i�њW���� �o�'Ӈ�YoO��A�+'|��o}��{Zh�`f���M,�ŝI�V����z��f������=M�,CX�sX�2�S]���V�ۡ��"�A&���K�#�d5��w�f�gE��v��RtIjn&P�W�N�"��%�`��e|m�s�r�q{���I{'������S���[Tvj�"uk�W�ӈ��;�q�F�	̔|c��@q���?�[@7]i������ha�}Ǚ�,r2=5������cH5v{���C����9cQܨ(l"��+P����&;���9�B2�.%�Sj�CZ�"c������%����.�~TWp�R�5����6��Y��T�#����K�������iQ�T�"�V�q}���*s�[N��]G���eUGb��'�(��y2��M@�������Ě�f֓�q�GG�\?h]*�ep�eh¸�X�2L����C�^�|��7k��������Du?�A<n�aمz<���Dv<�2^�;�J�b-"�dZr�r��H��ֆ|Nr��
*҂ɜ�
�0��h�¯�8}>"B�HzPE<AEb��C"�{��e�jN�~pwR(�m��0��A�.�/4�U�Eb���vc�j�>�4�ء̄��䦻���`��6"����7�$�?򜚮o[������dI�A��G��R�T��o��Y�eQn;o�ރ�_�����R�m��! ��{�#�W�G�{q�XކP��Q��3�]_��n�Yɯ^!\��K���(�-�CI0-�R��-��E53~ZW/E�	+g}����Ekh��������8�V�-ۗz�w�X���U�d��>}�I�?C����õ�פ��'x�a���9v-�~/^�DEd�v�`S@�'��6]w;�Z�l���-��<;.�z|�����.�,;�ˮ���@��d�k��3،�A�Ya���$?��\8ڱ#��(�5����g��#T��^}�$t1���X��oD.���Ф�C�B���Ѯ��Rfa^���/�^l9HZ���m��U�oR�k*�P`HQ���Jf���WA���o:�x�eZ�k��Y�Lt���a���� �+�m],R���E�� ���I�+�(��Q�O��<:K���˺�h�V�֬���d��M=��I�9��g"�	��l<m����$��ϩ(B�B���e���(hk��(�?8���Gl/��K�aZ&�Qas�68�ߐ�혹Cv��Ư$��C��M���8g�o�Haũ��t�|1W�Z�B��u�*�ۉ&�KҒ7g��J�o�T
��'m<M�۪'�X�'��p���$���s`	E#٬�d�^�,E�!��Eq�UN�i��Ɯƫ�J�e��T;Y�1d-��6Ƞ[�ƕڰ��K�\�6'��}¢e�ך���b�Z쵴�xO�S㴰�nEnd!�Ukqٳ�ve�Qvg�T�lr;2n���v_WԔ0�w���R��⊉�%����*��;���e��H�$�u��[F����P�V4���Sn� ����_�!2�O�?�{?�];��v���)�R�H����7�c jq��kv^�DeaL9��I�2��tf���8��v���ۉ�#�����������MߨI�]�i��W�����;��4����^��j���5L^
���p���_!��u�}V�����b����=�o��CpM,X��*i�>|eTm�/��N���n4��Jʁ4=?��_:�*h�sAlyl��~[��Q���`{�2���@9+��U���6����R,��L# #1��NE%�Է0�w���T�K��R�!xbzB�@kC�(�!R!��?3�4x�S"*�f�A�������$1?�+!#*r(�~��t�ڽy:>��g���A�"�[�7Gp��t�U�[��1���o�:=���L]� �ϯ$N�����#Ygƪ�R-)�'Qh欌ՍcD��wKo9���M�fu�9j^�KI�Mb.��dh-��p;����U61��u5��L;��{A�̽>�`I�l'��f[�Y�J;R�h��J�h�S�R@*J?s���:�Ȃb�7��j�Y�{��Ͼϕս6�a��By����טt$Ǡ@�	�1Q�a�C<d�����!��q(P ��#��tY�Dh�&����Vv��T���&�hl��Plx�ӦX���9��ﴒ$Π��@W���H)̟��-z��;C����5@�П��h0�lL�"��R7���yl�j��@��B�Q��=69N{�t�oaL?�CB���7�1����n��%��t�6` ��w8[	���UZFîG)H\��xY���������9
�w��L�XM�8���va��B���Ch&޿����J�P�1�HI㱦�E� <��+�����]
��qUkߺt�XE��[Ԓ��X�����>�V�W�gv��zd�8����fH�/�T4k�	� =ia��:���b�i�14ٰ6�/��S���ܩ��z�h$����a��G>���v�*FSe5�>*Kj�O��a,��>��V0�S]�X��1l�^�Ј� .:�N�"[�K����� ��2���ոێdQ�25���7�8������T�<<V( 5߷�a����I�qy���0?�w�t�*�T�q!M-$ieP��̺�<���sS/q֖Ĝ7��>����G����y���.�k�I�ž�l��h��i�G��
I-?�x`���I��A�}j)��Ό\6�Հ�`A:ϖ�
\c��)��d��p�v�So`�Re�Q�Ga�Vy��$8E�W\�����%2�DJ�8"u��C*����h^S������<-��[�6��y�Ғy�UeR��ڳ��Y(��rk��K���X���o��ʅ�6aA�R'vT�YsXM��&���Q�����՘�h�%�Fl��l�F��r�}�7�}8Z�|�|b"���Z�O;�17���5ߏG��T2猓!��Q%?Migm0����P_��@Π��"�w!Y�l7��#Wz�U�ʓ�[�)ź�H�1��%�E��6k�Dy�SwL��� ot��5Q&f��82��m���P*&}�͍q���o�2�^��_��EI[6��%��~�M?���t�jp�N'�J��ߍ
�2A�?��2��G0g6�($c����V��:��zWapoXV3��{�`*�N��	�#����^��>F��V�6]�5RH�ˇQ��ഐ̳�#���<����k���V1&��T�l9��=@�l?K�f�Pl�(���V#�LU�q����y�����Z��Т����=�
��3L������&�4t��O9�Z��еz=��K�d@�y����[0�L� c�DJ�]£JH��t��o���巭�Ԝ7߰���I�:%�svk�@���[�Nyga��d�̥�l�&��K]_�ּ�sC��=��V.��`ߣI���3+��N_�K,<q; ֜��*����3��_�7B�*�l��Ժ>߅pm��}&n������
�A��dn�^G�C��b�jF{rݎ����C�9#�۲�V\}�}�aa�����7�!�����
9�f<��T�����)_m�}N�hrY�*@O3gV�����z)a�  ���S�N��k,x��s���m��gGN��9�5U&���M��\H��}aa��Ĵ=ը	�y4%cw-�gZM`^_Z��xRp��[�
2s'�!W

�n7P
��V�2|�&���Yp7
5�磼�������Ĩd���t͓Sb����1�!����2�t��\��I�=�)$Nظ&Y�85;�n1e�vӚN�}	�w!��0_�:��1�$�7���G�n��?n����D`YB)�b����Ჸ�*H��3`!e���ƙ�|��責�2��3�����x\�_Rk�5�틮B0�=���5Kr�V@�؞'�}>�R�~Bp��4
��C��� T��j�%�e�g�����RӗW����V4�m��M��KwB��,�5����9�������i>>�$��ڬ7����1�5v�ʮ������2�G���ޓ4r��~$9��S6�Ͷפ�f�{\m�J���)��8v��T���l��ߑe"l��Q�r�~�)e�4�~��	�~JLo�K������\B�/�;Ag�֮^Íu��+K��#ht��:3���2�zl��lWc_�C?b�. �����\{mC>��4�E1~ziQ�6���M��݃|-�*��}I0���6��Ͽ_�U�L�&  W�u���wh�-���O��t��<D� �2��^��ؾ�K�r�K���@- ]�ڎ� ʅ-׾)]���||���ivI+��B���K�@��i��h�`/2	O�d���D�U�:��G�,L��{�"�\��r2��}F���L���ߤ AL+���m�eTD���FX0KE�C�I��w�?��ʴWv@�_�-�f�cǃC.��I?MK6���x�l6n��#A@�)3ٻf���5N�k!6g! ��/���<��LݦN�)���Ȱc��D�>ٓ`�/5�8܅�~�ف�Z�P��N@�����|���hwH�Y��^�ɲ����/�R�`2G%=�~Y�7�F��Q�L�%��������q�0�S���27z	��p(G ;�<mT�q�m�8a~.�L�����FJ�#�˗������ F�(=n$�����_��ٵ����r@IE��,�J��.��Ĕ9���ؘ���R�Ц.�rꌕg�$�KG�6�G�w>d�G[�_�q9$�i*�Q�Sx�dʜ�`��YMi����o_��?��*�^��\;㛳'���C�MR�E�uo�l���M8�؝�௾ݘ&\~�>f�J��8����Me���ڹ�^�%��C���:���j�,����?M����4��k�,$k`w�J2�:(/�:�`�A��A�>�)(�
$��Y��N,7S~��r2��Baњ�pY�k+���b�\4?=�P���J��u�C�jZ]l��C(��
N�u�ߢ��
B�$�v���^Px0� �����y `����(V+��y�2H9��M��2���6���eD�9C�k8{O���/��������u����*\�׃Ҍ=߄�G�ܔ �m��EI�q8O3� ?�7�T[ź��8,+<լvq�r4F>n0a�l5���'6�w�p��&j�х�#̼�����r�1���{�͸?���b�o¬�#�j]��E$?���7Pp�z����?�C�s/������|5�'`{F�i�;ڬ���H/����hl�؉N��2e�Ni�zGU5ľ���ۓ�6��"��0=4�����-�,�pj���zo�l%0�A/_�N�57�Q��MԸ��ɓ���1:��A;m���1�P��33]� �����n��4�����'��@zO���	q����۫S3�X6M���̽�eb��{�E��mX*�;��]l��IH��'S��	� K��D��ՠd�	 �������&c08Fb��G0�.ev�3ߧd��0��h�Q ^!���ӅT"k	:N�V�[�H`��5���8���bɀy���[O��qn��p橇��P�w�]Pj�n�����������O����K���Bڡ���N�[��q�f�~+��QP,7ӄ�M�!Y�5��ζ��$]���~����X�$�~7�j������ħ���jvD9�=E���M��D�z�T*�ο@x`y���x����DZJ<��D�\��B�E6��U����]��î4rA��2�x��+�3��p�H&%�x�U��|m��BS�&XX ��bC���cQ��Kb��o�EZ�L��w�w�:����,Mmk�='GwZG?�����8N���T�\����ds�~~�C�{F����2t�Cto8Ah��1�� R�O�5�3b.�5�j,�2��N�%�����d߀f���,���D��+*I���~�����9e��7X�ɸ���Uy��`�#a��ف�i����u��5�^������1�P��19�<6"�8����_����I�e�7�)A���
"��Y1zt��j{��G�|�/hl�쳶/{	�ԝ���,l�d��Ӕ�yQK���c�JTe:!LV4Q��N _���TNX��I�Fx�����1���!yr�ux\�����7{Q�5�)[��I�1�h��R�J�$�j���h(���88���6<���z�Ö-.I��IR,�d5L���K>'y��tGCxP��P�h�&��[���x��;ȰqP_� '���;����m��0��^���/`y�j��EU#��(S��HI�]���u��Z�K�>�U}���8�ސX�Uh6	|�+|��K�� ŐZ�z�����T/������L��3����ki�X,��+uu4X���'���Y�0��2��7�ߞ輀����v�b��ϰ��+���(�C�%�?##�;��*Y���l��"f��߃�����ů��<�x޼4�����s6(Y ݄�a"�UQ鶕?9��=|��lڗdi�@������|[�`d&���O�j�Q;DT��_V KUΑ�D���wyi]p�dGe7�S���:�g��R��:E��+;�y�����������/(���I�jh�F(<��3C�>6��O=L9���Wq����0�L����4�Z3�����W�� )l��1����>i�3�d�JS��JB۰r�7Jd�r+��-�S��f`��Â4��GPS=�Su��0�a� ����v<% E$L��o�r"�0秌�ǝ��w�M�����v�+\A�����.�+q�]��[ۋ_H���<8&�%?�VT�T��K�!)�|�Q�/���uԓ���;��XMy�~�^��1&�h~4-�$^&��X���{���IE8:��6���]�綤��ֶ�����>[�>�}�~�ƙ�+o<��4�ɿUp_���톎����S��N��N�h���鉶�:v�9W�E�1��~|���c��xV����?Z����+�Hf�J#�D����JU����T��gZ���;ؗ�2tq@�H���OR�5F"���ExX+UV|s�����d֓�&�Z��٪�����(-t����Jl0I��kTp+aa�
� V����]�1|:���r�z��� ��B�A<6�w�����Zx0���)t1-��)�n$6	��n�vժ�$o������y]8�~I�dL�6�_�X�k��L,����x�zYT�y<%Q��~c¢׳�7c�t*آP�x��
�C�A�e�j� ����3��\�L^�K{ۆcc����a��,��R8�����ێ�����i[�>�p�܈Ĳ[` �>Z��c^����'6-n��AH�Vls�>��i��&�4;�˕��T�
�W�C�뎃��^�����Qnv�;ɗ�4����B�
�z״� �?�d��\�!��O���JQDw��c���\tM�c)��F���Y��*P/J��lA���Z�� ��wC������Z���3�݌(Y�?��!Q��M�?��2������{��u�ݼ��R=�ɷŗ���=)�u��iz������fm0�?`a���;��9Pr�I˹.bat�;'���_kw �ֿ1D�sHzY5-�����Ѯ�"+����'�P������Ʉ^��nϣn
+�o�*W���o���������5�v�"��`�E���9F"ʮ�SH�t��%Hv�c��D�VH:���-��R���m%C���a'�y�1~��̐��u�Ӫ���?�ѿX/��� b؅7����!�~���$��,�zң%z�l*��*�6"h��<}֌����/3'JW��(�}Q���V�٧��<��-�'�����g1��q0�	?t5�#��\c���=��i>2Q�h��i����ڨ�+���%K�s�<��:�ޏ�����~�?f��6��TF�aYӇ����?��sQ׺V��)?+��Ũ�6#�����p�.�dr -�;�&��+�o���,�*\�!�4o�[|P7\�8||�nm���)[N�<���"�b���_�ɹ̙{��;�ڣJ����V�u>��D���ŀp���w���LD�#
r�H�F�jyõ������ �68$݃Mo��zNO��~>=�б���N���+�6ҜD��A@�����.!�������j� w�薜꽯�X"�	�z���NI��-Q�Z �yr���Ɓ����x�Eu���-� :q�=�$��S��痎TY��x�vZ{�-]�p���d�kmL	2�5���(2+����SSn��J��:���� ��*����$�)���_f}�!s�B�M(�@�4��8��?$!�[�?"/v�kj"S쿵�
��-�am�Z�]!<ʞ��W	�_��*�T�;�G!_�א�/@a\?,,������Q�=ag��1�T���}in%�`-����U��'	uVIp���QW����đP�#*�+�9���� ��d{�~	-���@3��oP*���_?�:8�������8��0�+�fZ����[��_�8��O�_��?���t����?��&�x|4y×Sb�u�"/䣫�B�Cc��ʛ����b�s��ϊ}�����2�*��i�̟�5ې�V3?�-?!��!��U�����e��y�̊�ȉ��!ݏ���DhU)��]�߽�3᧳y�x �7�r�|�Lt޽�6��o���R�#�+�3�%���L&���MК���(�9����إ����X�Vi��$ RE~�}p�q4mǗ�9�&�j��%K������Is�VoO�Q���'��݌�A�ڏP��qW����,����.u�Sl�%�-�"W�[%�}^}��#�q�'x'�	�q����͚O���U`<�wk&�v� צ4������8��n��wsub�����=�`Ls��{�2~ZRU) �	��_T�/�}�'$����N����IHi�&��b^�
H�H�2�Y�@����8�*Q�W�m ��j{Ɔˡ;�R�8�[XT�R+DyLj������7��?.��K%��G@u%���D��k���{=�n���(����S62�[˚)|_@}3�o �9V�ʂ.�G�E�r>��Yw,}P�N�p���gdCZ���=�<>�T������F�Z�nj�=G��n��m�(�j���L�\D*Qad	�.�D]���Z-�����I�fS �$���D��}^ �����}�`mf���!��D���;��g�Ϛy�������-�[��Z�+.������o�t�)&���wU}.tN��<;E�=[f)V߀8=�`@�['�G��1p�S���.�F����K��{�9��s��W���^iCC'�S�{͊�9b�Kx3�r�H���D������1Q���\u��.�E�Dq��K'�ͺv��z�XVЏ��Ax+B���>lE�E�r^��_�����;c��Z�.1�*�wE��%5��wA��>z�~����!F�QVR��d��T�	 [߶��J2�K�wձdn���nu��|>�k66�h�t�p1��n�%Y�U|^�C߼�`%�/��GS�*&;M�)aKP٠e!�݀q�����)n�l���[�G��mQ+�(Ѡ{�9�Z��<:�r5�X��ѩ��������Ҕ������j��c '���:�t��w��r�,���F�fmU�Ғ�%�"�\(0?ݐ�҂�߇�$f8�95�E6�/KC!S�<�`䍫��@*p1I�G����?(W�3_=�#2�Pz��8
8Ȋv�E�	#˼���-ZU9��ˢ �U���=����,A���lS̗�0ٔE�Q�	D�'^��3���)R��C�t�W0�����=t!{�ր�ar~p'��:`t�G_b5 Qe� �|�xF�d@UٻzjN�y���W����¬|g�����/��z0��y��qs��6��;�)��(^*P�������r݁�`�ZG�+����Ap�2%�#�w_�KVUR8.�5W�*��gQtc�a--����C�o�Uo���D�6]# �"�'6�+[�O״̝\V�E�w�����K�!@�<:5b|*{�@F��D~F�[X��8�(.�������#t�4_X�$" ��xK�����W>m���*u���ok��k���T���=PS�eRWv4�W�t�;�*-�,�B?L�a�1�h���;w�c��B��������W<�6�k��P�M�TZ#oӖ�6K��B�����͜s���>��օH�T�����w��h��7�0�ׅ�T�523DK�&lW���0�p"S������L���o+ۣ}b0�dL=@횱�m�QJG�����@�c�W��d����7��/J��9��um�fBk��w_H8-��N�O꛿��o��L$i%��ԦR�B<��f>{]C��~�-���6�F_�>���V��z��q%�D�I3�5R�0�"O��o��?,ş��m7(��sf�n��C��7�������@Gh�$������p�����^�Q���ɣ�x��4𸿵F!���
i{e*jC� �Ys��� �ڏ�aRڽ!��M�aY���|�i���d�,�}��l�a�b� '��-�,���>*G!(�QD�� �0���� ��������zխ��
4���2	`�@of�x0��o��V�O� �	1>*��T?�������:iU7VZX3�7K�+v�'��������NH<�{�Ol�a�/��Y�.��lzP&Ǉ�3��p�&}R}�A��W��6��=��0�Sr5��mvzxa ,h0 }i'���{�r����U��އе���K�'�7:j�q�a3�z�;=!vɼ��l3Tf�/۱TScG���=9��i@��tn�>�����zs�9�5x��s���#��e����� &�M��:BBb��w?R���<��v<p��u
a���+Z�-��C������L�i�/h�N�V�^+�~ٹt���;�k�D����X����Ni�hx��	����Hm{� ��m��oD:�E/�3�ˮ>���?&XH�rM���O���
���X�i�q�cC�V�]w@��"�&\��?���i�Y��8@�����п�#wՖUkjc:"X5BJ�):���4ߎH#p��6��Ȇ�M�i�	�w#�H�dA�sA&���rP|Fe��,�r�v�c����M�E�� x����p��UɎ	>���rs'Rw�*I��' D���<�A�<պ�c��}�U i�����X��ꟍ�^?��!3GtZ&G�.���^�L�ق!I&]去�HQ2/�ќ�~m�b?4���Ճ�M�i��n���)��&Lc�\*}�A:�C���k�ܓ�{�c�O"}�KU\�P�J���l�(�V�88�BHn��:+2Jh\�)�(>f�r �7�B�;<dG�n���ʖr���2v��,r*�B�iT
���FrA6F%Q�Lr�1�H>|����.�����Un�1=:_�Փ����μ0=�*�ȣ��\���\d�&�)�����w�G����@Ŋ�Q�xd��<�&�@���Kl�<RaÌ�$
 �'?����Ӗz�I�~�"\C����C��Wܕ�Z���@������7�,0,����.�Dt0��9K�}�dJ8u-5P����7��U�ǭ�a�,���=L{��=� ز\.�=k���˞����5[b�]��!��kO��<7�.0�=bB_����)U���}������D��Tՙ�Q�O��5U*�����k	k��	4�1&�ʔ��_o��h酋�m������{vA�#6����(��!�?WA�},�VR�������7��'�*@/]�w��וb�ױ�ܪs�H�K���8�e�%)���)�pr�v۬�K ���Ǔ.��k#��]A7�5��@X[����1�D�;5�3��|��`0�	�VJS��i�oYk��8���@e �$�k��)ƧʡP�M=�|/�����G	Hu� ���>�!��]��/�r��WoB\����DQ	vQ����p��@�N(�w��p��^�Fq?v�M����"3v�4IIP*��l�{G�FO���t@�_��9�t��x���<�?l���ϣ����]5s��������(!�d��-F�/	N�B�[�P��~&�O���|-7��f���ę��Ҵ��Db2���7�w�)�QvE�ͦN��R^�� ��|ٸc�䉿p�륆��*�������{a��Y� ߣ�-���Wՠ��j
�Ix��{�]��6�̚-���9 ����\E'�IK:���]m���]QOM������]�u|��'��g�o�j��'���Z-�E�9��@?B���ur)���1Z2}���
MU�!/!��In;�ў�A��:�?㞰�i�Q��g���.p훥�o-�*$�� ?Uρ(Ÿ|�)F�ډc�2dN��Q�\#<ad�����f`ah����	����Y�s21Jݾ���Ao3�t;�Ev ��Ý"����/�(�A�w%����	�""%�
4�����D��
I"�7۽3�z�V>_�� ��`�k���؝�z����0S�и�溆��/����Ji�<'�r��k�}�:ݝ�>3�~l���^�?�GU�g���`���^p��Uh�h��\Ğ}66	�s�0���Z��
���������O��O1�T��z�B�0:��Ö$w��l}]��2���&����U�Q���3������jby'_}ո��B��\�ͧ��p�2H�(t�X����v��f�JE������j �8L�^��<�&Zs�ߗa��Lu~]�-���<1�W0����7�Dh�ɵ�{EK�\�@��2֕�����р�7.�rfyF�m����U���7�-�_|�҅z�S,��WvW��&�l��E����6���9H� �5^���w����^$)�U��_�
�B(5��m҈�D�ڜNń��w�@V�v4U���D�17i�gvB��#Ǵ�h�bpOŁ��*��U��T�P�@u?m�\�pm�o��7$|=���M �U�����E'?@�_ ϛr1�t3�SD���(T��ݝܝZ���O%#y�=��nX�G�c��Z�3��T�A���ƞ�I�Dc=R_��x�.�� �C�"Et֠�>0O��Tѱ�`��"x�"�Ħ �Bd }E�˩���!�c�o��S�z^����U�6�D}�|���".���h�`v��������>u����kp�����i��Yj��B$6�X���A2U}%��6��9�tsڥz�V;CTL>�Ic���")�S�	'^�K�!r�~��T����D�����9��B(	�J.X����y����{#b�QH������Z�:$��ɥ�.��ˈ�8�'��l�̟ͨ��,N��"В��U��M���������S(���Rvx�GRs��l5"R���m _��T��'��3&�8���/����þi^�6o��ǚmM�C���V��U��j��8/w���۴'QKۥ����B�)�ٔH2�\kf����Y��D�(��@ף	-�O��"3yE��d�����9�۠�E�i�+g1�)�M�����52�l�o����U�S�jK�T�%��Ț�g��Vo�Lpm�$6]�uX�+̚ݵ��0P��ݷSի�{>^�+�A�=`��s5sz��y�^F�������$�%�Yf�7����_Ȏ�+��?�����
�>�,�	��Cٗ�����o��W�^�_i%/mO�ڙ/�6r"�?�̹�;��:M�g�_*�6�(�[�7*�%�)+�+?�%����%"/�~�z박I�L�pc�g��D'.��]�E���@Q�S���R�}�G|^�!�?��*E���0tM�Լ�$�}��:�/JE�{B��I��[x�Q�Z6��I��������B�ۨ�K�4'����S}�`��x� (���2�'�î1qf��?�'����i]���FzB�j�?�۴�+p��~� �	���{4UeЁe
Wb|��GC^uQgP0���Z%��ɇo5$��񘻼�g�+�p]�E��ѣ�i�0