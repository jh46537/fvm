��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�Nf����>qXQ�J�y����
5{�D���??���s/�I�ń���!��a�pCP�����9:ٕ���$�>��S]^s�u���pW�Sۢ�Z�l|�۴*p�&qx��\X�	���&���ιQ�_5�Px̯[�e���ibU����կ3�D=�rO��TO8S�,�����**�'l|/){oEŵl��C�5�(P�֊�1R	Lo��,J��"���/-3Y)Dɭ/�'ah�����Q�^@75���
K�1���r��-�W�vU�o5*!����'��;cQH
����"�4�b�dD'n���� �M�ǳ�J�����X¸W�}w�Gk��"��6or6�����g��(- J��O��8=h��=��5�p��E�E�5v�����Y�TCn���C5�1o���ً��pl��>o�)��c;+�!?��M<�AI��Q��Y;�H��E��:�)�pj�1}��H�~�*�z���
��_�Q�|����F�F���.��2�K�M��pp��2x��l
Q����:"!�Z�C��-�6���ۘq� zgUU��校���/��Q�	rf�[���G����X���w���7Q��FFfF#�$�A��s'�J-��G�ĸ�c�#2��$AS���"���/��n���n�a<*�����j�x�+Nx�q���/e���c�E+z(���N��8V-"���>6���g]��GfV/(��x2%:}��a�7.許]pm�>_�x3i�5Ei����%�����";��K��~�R��U�M�اi�0Tm����!7 c�K��ח��� ?��[��l��֩�mIh��Fs����s>K#�|c������cw�"�m[��)(T���T��ܠa?D_r0W>7<.Y�4�g����С9�^v��~��h.@�v K��
?{�}Ħ;�P��C�D=v�+S��9�[��Lr�#o�8�c�
䴂)���߅�z;�ء�/K��m��5(ۥ�Y��(���W#ۙ�>���{���n���3���h�h~��J�4yr��a?;Y(�+�j?T#��w��u�{�����]g�Q��}�2�8g
.Va��&�>�p�wj\XN�gD�]l�_�,�뇖�%H���B���l��T��'�"Z*�??n�	�^C�"��w���V�֒�"��*���bXJ8�3��'�f���ú�Q!%~���|�wȺ+W�l<�
%C�$��)���j�޿���R��5��^�����Y���p�8$�7��u4��D���I���V��)=�8�KD��>£��<����ޑ������1�v�X�w�5R�-���v&��	tU�����*�]���feM�u���O�Xӗ��G 6�Q�J��:DZ%�F�\�Q:d�P��k>L�v? �a�?vrF���|���!lyz	�>X.Ř#�A.�E<d4�h_Y�w�m�����}ϟnߘ�˘�!~�lW��s���4���`A!J{q��Ry�~b�ṟ��6\S��-����+�TQe��C��Ž�x��0�N%)�,0�215��KoF@��^��t���嘪�|Q�W^����m�Hx|���epLi��Ksx��);ɩ�X[i�g2	5����%ϣ`����Ŝ;�ZB\4��͞�[P�Y�������y苨A�
*r�]�8������>����"&�3ڮF�� ���g0?+u���S� 񯉜�
4s��< zQ��P��������$c���Q�7m�UPSWXU�gt�,��d���#�7�{�7J�HǢ��G����A '{��w�c�#1Q"�tfڐ��A%��|��C4� %�^�	>�#iF��>�V��"A�,}�u�]����Q:�.[Z�0��K�^��e@Ɔ�lO$�����wF!񼧃�z�*j��:�A'9x�iMjw��s��ǺȺjQ���ҏ�P�u|��U����>�؄�ꠢ� h>?Z��__b����w���8eF ed��/�fZ|/E���,�L��Tʃ�h�*�@DҊ㢏h�%(��&h�|{�ƎU��a�>�����?�����y����S/qe+��ⶉv�*���x�����EP栽�1\A�4�>Y���ժ�߇-�ǈ�He��<���\��k,pU�$�#<7���A������x%s%�r�A�+��C쩱1���ӆze�Sx5\�_�;"���Y����|�o���+p�b�k�� ���FA�r�\�v��Hc42��
r��8����kCx�XV?�㤷��f��d�k�ޚ ���-2����k<lV����1�]��Fe/�b,}.�c�"āNP��>�jF�>h���JJ�T�GWh��Y!��m*)���	�Mp�9�O<*��FY��_���DG#��9�j�?}&��kZRI��U�
�����.�����s�	�q`ޞ���,�&�C�)q�P�9��MԶ�Z�/Y��l1ow�M4W���h�����^����T���l\��N��jb�^����"	�*���ꎍ�I�.Y���ZNF�4��b���ٓ���i�]ju	=A��>_wS���PCO��%�����j�p��yÔ�w`M�]���XX�6�s�Rj�ϖ��!�l�2sI���;���$��I�ױ�jqC�\B��o�v3������ȶU_o����࿤Hu���{(��3y�_r�ߔ��(-`A��_L�5<I�z<����}/���;\_@���{��;�0!�~��47񓥷���8�	=��O�D��c.�-�i�g��NǛV��*\�޴VV�)({�p���ү���@�n�|��Cr�p5��j��OU i��7P�ds����_��s��!V=��w*ѲI>�]��x�EK@j�_�f�����X�d¼�au�ث�幟L���0�r��k�t@�������x�@��?�(��r����	���
90߂?�o(bfN,�;�D:���ѿ��3@� ���<+�֤�v�1�XS�T�i��-���"������ϮШz���"�����f�< -���Ӕq:�Ou�U����H1��@-Q���@�+|�QR^ȆF'�E���-LHT����J�^��J0�Zmx���1��_5�ix��Yp-��Yܡ���۷�,���R_ap�{OQ��ߚ����e���gS�#����<ɋ��}�'Q��t�z~R)ԋ@�������r����8����������E]p�|���0�qkN� �X�
����Z��r=�W�IA�&:���6eAi�2AE~}�Y�J�\��~{����Qϣ_��An��