��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S�VJ���ɾ GK�rA�!��}�x�E}ݨk�fի�u�(���L K߲w�.L}x1F2�#5H�:�'))�6_��\j�S��W��w�.㆔�[NQ�6��iM�@��9��eh��L�@�Fb�%FZ�"e��R���W��@�s3a�����膂Y�:�D���!G��j	�E����}��Ui����kh稯ka�"������e�^��6�ɠ�Ij��-���jW}e�@,��=��\�`�Ǩ��:>_2�)����������t*�� *��%/��X_0�2�KwS9�ڪaԟ�	�踷Q����Z�@Z|�歊�)���ܰ�K���"F�"�;�ŰS�d&>�،4j�o�9���xD��h[JH)���m�tS����\�ɑ� �n�{ƒ;PM�����>"s��R��m(ɠԉؔ�W��6���ߜ=�5�%�_��+*�o/�Wv/�nW�S������50�u#�����=�O�3b�w��Z,L+F=5�'�?y{��yN�2���D2�m� �p)*�CW��F�7�Ye�ȼW�xs	p���-0Gnނ���Q��	��q՜o
����D+�g��!!|VeG*�s�1� y��!��FXV/ao�
Z�#o �xE5�_�=��جƒ�K����#������\?xi`i(d����#���&S����$��a%�o5�H��}\�����?�ՒI�W��+|Vz/:�2�T�K���f?�k��A9���d�̺}���6���K�����T�ʫ�n?�塲������*}�Y�9�{��S���c�{ҩ����H���qn����qh��W�"�&sL'4Z����B��,8��w��BFd�8M�Y�b�oe�Wl� }�$�ՇD�O����r,���1�υ�\\v��<Ɗ��h�L]@�'�Z{�e5��w~��t�qJsP�X�q)��"ˀ�-׍����������@�(� ��bx������O�3�Ӓ[O[	�Q�����c���x������_��˸)��+��hNۚ�-�4�G�[��T ����r�͸���6�GY����G��E<Cn'C@>^=0�DFj_�hEň�
����6Yv��ݚ�n��r�'U�d/"�OS����<�N[�-��������O�oH�Xd�K�qF����mʞ淛�vKBDݽ��F*m��W0��iH*�SM�-s��a�fո�5/?�ز�yw����Ʊ�^3�T�%��ޮ�~�N'kK�u��M;�&8&������0a��B��{B�t����@ֺ?n~`š݀۱�
���
��ާ���2o��E1��*?�X ��1֐��g�0� Z�(ӖrA6��r|�5���"M��� �zrU�Y����A��-���Ӂ�Q����Z/*rl8g���1tFC�c���$	�����K�?������5w�"����xG��i�&�k}�k�*|}Ӣ�#K̉|u�_&�o@&.�
�\��w���ߌ��L�S[ {��3J��2���F�م��%���}~t�:���]�;�q.~��j�+i��L�_|D�s���Qa�!�_l����=->݅�����()�L��̾��94�ċ�2C4�N%�*J��&�+N�,'/0�^,a��]S����;�A�H�Ȍ�6ua�=����F��%T\�4���K�I�2Ӡ��R�D�-nt^4�P��y���ڹ,]�j� <;�f�I���\JY�Y�����Hu���RK�C��p�2k�a�M�Ǭ�uR c�H��(1����" >��[:�
�⬿�(���r<3Ku��K���{�/�6���w �z��݆�����-�u� R��o1O�[~�����?�b��)�9��L�	l�vh�/��?�g]be�*N���)N�W�ZK��x�)`�*R����6@ID`����vFګ7��*�^�ck��/�عx��Q�
>�]I}�b�&D%YD�E=�-������m�c"+�d�'i�,R[��a�p�O�2	6��c���~CÈd�BRAڬk���t]VKĕ[�ρ~o��������1��>�t����c��x�X,�F �h��������ő�s�֓ 
N/�m�y�VC�����B�������e��ѱ�nBx�P˿����H)�������p��W�Ϳw��"���4�Z���?��m���
Z�a�&5�=���Ԩw9�����j�����5mM�׻-�z��EN�C{>�@/�Gd�:%xə:�9,���̀C6t� K�Iγ�.�����d�LX]9B8T�R�����l�^��V�ӆ�i��4��g�s?AtH;?�Lw-U�yg���ủ��k�0� �"����<���o�dƗ�pBg��#��r�a(��ho���V,�b3�u@2dk��'<�t���GcV0�]��,��-��挙��*��^���Q��Xomj(j���C4�]J�}$��b91qb��@t�+L��4JB��5D	��x��3�1sZ>Vب0���� ��w�?5\hea�������F5lCҥ��v�֓m~����/-*��k�D{�hi�Ђ�������Z�{t�1r5�\z��Vb�Ki��~�Z����?�� �,�ֲ��l���}f��ɑ!�`��j�bpǖ�8�e�ޚOK�պ>S�E�Ni.�G���
wy�w� �Y����՜E�'��gQ<�w/r;Ł쩒�Ǵ^����U����Ƨpy�6���5�kD^�m��f����"I�S�D��H��y c'�����an��(��E��0�!ȱ���Ԥ#vR�K��y��	ϙ@���2J࠙��*g��A�\R* �8^�el�G�w�_��_n��C�h��dx�H9���٤{�~7|$t�fH��Od'��08q��P�v G�Z,���R���Ȁ�A6��&�y�p�t]��0���|�af@BE�� _^oڜ�)DJH��c����0�t��u|�F�OG��<����o�>Z�<,�^r�݇�4%��Ѧ�x��*�`QUߕg��>#g�Fʟ�J E���N�I���J�p�L�W��I�Y�$��6���	������t���X�B�-��X�e2"��<�����[3�=�}�RG��!�W�܈4���l�C�"����$�Y �;3��ͭ����Ҭ�
�;�?�[�{�᧔����w�@�]܌4$
���3����輻Ta P%2P ��C�N��pg!�"Cy<Ԅ}겡6>��k��7�0���X���ෛ&��q����]�2��'3�3�k���iuw׋@�q>2]lMT��p����s&�d�IIJ߇���k�[�0W�b��h��(b�`]�JI?*
c��^��$Zz��LI��t�@�`����2�KƔ�ȕL�.Ȑ�����%X�TQ�\U��U�假"���T�s�?���;��h(ZU^385��J����4���Rw��%��GxV�'�)WK6��T~�"iS�A�0c�̚ώM��<[��Eϕ����y�(дּ�Zl�"��ܹV}0�>\�ɽ���g��> g�O������Qh�;�xѸr�ȿ�h�B$��Eҵ�r5�w	�$*�W\�Ф=��`ؚyF��s8 �4��6
䮽�a˙w>��]*r��@,-� O,��S��Z��f�� R��IC���O���d�sU���x�ҧykz�m|���X���8���Z���6��2gB�a��gֳI��X�"��B�L��Įd0/��V�?փ�r�U��'^�"����?�����_�Bm��š@�wymx@�i/�"<`|����+���b�,0��;���fz���|�}U0}��KҜc��iz���l j�t�v�$�n�!��D��s�����::��&/[�rJ��x�xֻ<M$f5[�'��:�������l[P�E��
m yB�17�Ѻ���B�w������jӜE���7�	���Z2iIO�aƓS���	�\���x8��b�JR�WJ��4Dd�P�b�����)^�on�����Sj�3[�n�ז�]z�I��� �x�Ci�h�b��)�ܛi�s1|{'���p�SAE�1�P z��!�F��4A�ެ���Ȧ��2�T�w5̘�S�N�Vցs��� ֌>�\�k�m��E��P�T7=����X�#R0��7MSW����=a9�I9�QcnHh OB��9��}Z�� $XL�VU�f:�Xv¡(��In�N]��CC�/�SK')�(�%�������I���
�l�Ǩu����oH�cA�m����!�c鐏�1f>�>t��Q��g��A�K�JN�FM��q�k��S`��'(��ݪ�(foC�2�\ё䋚��*��/�bGr�'3b
T���D�����q���&��&��T�YP��v��0��'')%��P�d����G3����������c`(�����gi.j+�>�y��Z��Q�*(���
�������l����ߐ��`,�&�zz<��'\��W����	�Ԯ7Z���wє�V��W��Ӷ,�u4�ͮ���3��X�e� ������yp����lν�;����O���$�ޱ���� �:-���eg ~x�����3��lY���.ΌlܬA�
��.��1R�"�B��y^�6��c�Ak�!O��X""pqz�ʋ�9��9a	u?�]��4�Q4i�9j-!��C1��M���}��~�0s �Ír$N� ��%u�ӈ��U 1P�������2B.�&My�H�����w]T��J��9uZ=�@�2�:�o�<�77*`�H/>��d/P�1z}��pp3�g���1%�6a^�=K�W)�M�?��BK�-���|*��̍C�%3���Md�L�j������U�;�
d��O�,�3���=�{S��X�4��	-#����JȀ��pkk���!�)��K��~����+�o���B�G�C|xg�O�����GK>�Q��7	Y��O,�kMwv��)f�O'X���{���Γyoc��S�֕Ok�=o�Ⲻ|G2}L4LȁVBKŀ���%����D50w	H��_ݹ���߫���ǝ�єă��'4���+%��D��5g8G�����e�J�E�gp4�h�Ж�����)�3��
8>��-��b]D��Y=��wh�qm�§��ƭ��s�-�.�,���V�w�Wױ��2��Pk{�Ŀ����{�D1�E��r�I,;a}V���
�L@(���!�z�V�v��� J�U��ِ۰��Ns�aa�0+����4謿����$}��r�h(~mkQ���v��B�C��b�!����{��S��K!*%����F*\wT���Sl��F���!,��z��:�U�6@�"���)jFK$%���������V�ͅP�{C"���r��hjk�0s��V��u l�������_���Л�� ���WoN=Ê+������Y��I���GP��eb���P�O+������3��Pͮ6O{=!I z��`G������W'�h�WmEw6������'I�#�4Ҫ��y�R�wԯ�ύ?Q ����7��V<�2���ro%���{�Ba���]!PDkj	f).��}�K:Q�g4^��>J#���L�Iy3==i��fj$彛yl��F�?$?�����7T���1fC���:��5�A�ٲ�EO :/�%�u;��y��K�es9U�^�x�)Z>9B̺�1��s�*���0�1��c���C��`]jI4lW�"���Z)āc�s�~]�IOy�Y0�}�5��W&/٧"�X)\-�l���� v ~
RU�bݲ]$ym�p|"}�H\�X��Ƃ���]��x�ogG�R~��5- $	L��
=ptw�>�#�<�	���v�y?m���/_`��!~,͋%�"]sk�GH��
?{�B�hO`�1E�ʁ���S�Q�tQ͞�\���(���z���Y ���ȧ'l|瘰8�cLUp�k��	�f��������f}�#@q��z>~N��sɞ1ޯ�T���Vj���YaOPk����p�w�Y@�����8t!8�"�;�1�'��`�W�����hP׫��<��+a���[�Sw�=W��\�U���N�j����⃿7^X;IT��ȓ"�"���#C7J1�:�Ac˖����[�m��ԭ�gcǳ����4�`[��� p�i��\��B�F^��~��p�S�?�(�,G"�OGcm2%X�Ւǃ��;<[�0�Ts[�w�5�ٔ�܋��Z���:�`!��r���$�>��ڤIL,�7��L\1t��qe��eQz*;H��#Ld��'u�Cy���?qQ ��v_�A�e;C@$Y��r*6I�R��v�/��p�!KD�v��b�ɥ�'���]0�/N�����zH�'͏�T� �)�;���~ ���,KeNa3�-쥫�Y����)�Az��C��N����i)Mí��m䤫�4���AH�hh�"�{Wt�p+�'&���,h����	.h4[�,"�A�k�8d�H������h+[�#�h���n$�h	��6��2��_S�	:�DT!��*J	�r@��aX!P*�����8���\�?��-�۳a��x��	*a���k�KP���S��b��(5�,B@�����1�'Q��������|:�H�_qO�+�rn}t�(����R�qt�Z�8FdF��jOq`�N��܇����r�P�v�(���cHj|��<6m{L�ޟ0B�-�4��J�9.��jY���E��'p7�x�&O��(��ka�an
��{=����$M��j��:f	��PDH.��[�ը`�/>�`D�Yn�y��l�n��k����N�4(��״!��֡zCb���,Z���8[���B�W��k���)�Y�_�����7`g�ݧ�9�TM���}yۡ��X�K��R"=@��QB$ �v�k -w��O*����m����-#פ�]z��m�E��oDخٶG�ndٸhqZ���'�L�/5v�,�h�>	����F�8�fn|�(�mi�oc�e�	z����?�!2K�2����R���m�ժ"�~8�I���s�C<���п�u	�'�QU��|��Nx���쿌f�3����\��m��w��jo�@#�U����(�?K�Gki@�'8$ �(���M&�:���Gb"�Z�"�.9���+b�B����l�ʭ�_MY�ˋ詰6�e��$I80