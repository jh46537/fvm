��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��x#PcJk�� � ��Z�q��Ւ�K�$ꈵ�(���&m�%r LFy���JCLsOBl֏�[��״3��,z͙��ƫ��6�gJ��-)I���h��_���;�*���댗�P=YoVs�6.��4��s�F�Z��DG�Nq|J]�2�&~n[c@�y�d�of�|=xC�ŉ���	�t\�q'ԇ�1�4�s^e�版��˰K��r�f��!}v飵r�x�9C�3w �tʐ!�,�!��pN����� ,
�@��K�w����q2�!)0|����ė�'��-7�p��=3酞�J�t�d�����7�x���,���V��Iѧ�`�%@Bl�C�[�o!4_3�pT�DhnC��4�@��ef�-�����g���>l��:����@���Ip��J}o�e��m|Te*���G8{!�m���
�J������U�uVv	o��X{����Pwʴ}Nܮ+�}-h|��Q˗��������>����s>c��T�n>��t�S5��R)JBn���z���i�>l<k�����]��Q&���4�	��BW�q3ʨa��I�GM-�Bbrsm�?��"��ov�a����u��0meY@@�mp��
���Jt \��Go��ټ�mYN�/
6�T;K��"e���i�q5d��+�Z�y���o� ��=>�f�M䲸�n���ę�%apaA�J��]ךc_�
�x��689��c�F�l@$��7�`j˓��1>�X2�#��߬�ּ�ce�x`�l�c�<�
8g>������1���\ˇ`�3)O;BBw�M��Rh%�*�?�u�13��/E�/e8���Ur{,����U��fr��WU���
FԊ�����UQߟK�\���m7'�P�H*Rֺ_��߸�#Z5M:�f6ȴ,sb�A>"��Mzw4j�vdX�V=�E�D�����v���p`�I.3�u���.�^	]���=�6fޟ;3���[F�k�����]�������und��=~~W-E�@�E�-_\1L��t
���HW2���/�j��|��>�6�_���:`�&'�䪐��W-����4�o����E����������Ž�+�|!*��C��}�&�VP�FZѯ�ƃO�P�����@������7�pA���A0JP@�
ǈ�(����s6�3��?�Ԭ���y���$ɴ�<����6BL4%�Y	�h@�Wz�]�y��D���G��-��E�໷�x!}�o]���/Eh-�(+V���������%`BJ��=�S�RT�X|"ȝ��s��)g�ϰ�h-�#�\�5C�]d�%t���0k�	��.nGoZՠ�v�&J��MT�y�N�m�IC�M~9�
>��Y���J�i��&�aX�u�'ү������(��h�6�H�0�n��V��:�q�I�m߅�4=��1���{�
�Z*���X�|��4^�bw&1Ci� �SKj SV�E3�iT�Ї��m�!0��6���r�X.�;�����9B:'>\�CIC�Ys%wx�UG敒�$)� @jU���diQ�)�G^�A/����q������B���"烣�y4�"fz�e�+�Z���3���ؽ0�Ɇ�d��{��߶�	����#�nQ����nOP�8��a��[W6�;����^�0���� }5$g�M��k_N�P�eU�g�F\��d�}��l_}���~��⍇�ڎ�5�ՇH�k�����KaB�o�{��+�{�1���1���мgTĳ���9=�y'��K���WC�V���
;�roo�N���Tl����kE	�����6R��r
+e{,*HJ	����%oי��M�����B-X�s��o;��Yjm�S��`I�������a�L������z*��R�J�!�%b���k�%��2��>ϼ_�"�F�vu29�G}kׁ=J_��i�%a.���6eԌ�<IvR���yd+�|o��Z`�q���	KijZm��P���8�ޘ5�A8;R�|l^��&�>�e;�'��/��SoD��������_k�f(%M��a��!Պ�����)��T��,E��p��3ӛ���U�f.�"�"!�ʉZ�@�@�6X��G�3��иMH�����O�G��*� ����h��PhPWrU��+xu�����X��Z�EXTZ�R�t�C]C1uH��IM��@R�����)��lH��	 ���=������먃tl��;o��c?kk���"g|�<�!�v�7{�u_�v�(8"��t��-��xﴻ�9�I�&/="�U���ՊCBs3���M�z��1��h�aׯ؝^�<BZ_+>%0���r��Si�^���̑'w/�$P�
)�2b��@q����!3��	�	��p�}�jų`VOR�G���M����lT�\�,y��U�Q��`5^p>�w[�����j#��=\x�7��8`�e�.�F t�D�+�;�h-T\S��/���Q�ε�kn�����1�ʮ�ӟ�*�u(�Ӡ{&� NJ�����]����v��Sl���l����	�M&4�\ʐ�&0||0���O��$��jV�V�9����0yaBM�P��R�l0O)�YT�Ti�2R��ڵ�|�$j0��V��Ie��ݎ�2pm�+{E�V�V��G��çy9�2f�%��'^�$ZlAy���#2��=�Z�<��TI�^x2vix']�����T��ֲ�3T��ە�p�& ��i�
@x�[\�2|̠��:ő�h�����*F���df�Wȶ"0∷#��Piܢ�L�J�m�j�0���\ɻ�%� a�)�r���Qh|ϰJd�q�^;�M��1����Tz2���rj)�m$'Pʍ��I��n�/�a��a<���8�q���V`����s����ߓ� ����mè���3Pl���?�*��Vn�"x0P~��`��#�Sx�|*H��2a��_6��0T��!+���Ų79���S��:��)�W��#��F�W8����mK�L�h�e�ķ&mB#],�ř���F�:��΍���SI��s�#��'���V��p'Z�P;�H�n�=K����Xl��R�9�X��r\x7��n��^j��������Q�z(�4�GB��F��� �91�j���������l��Lqju��)g�ӿ�ƭ�=k;�
} >���D8�U�&�[vft�Ra����Z������
��ޘ}��*K�꽍�Ľ�萹�������it����i0G�a����-тOk����� .�����!.5��g �F+zl�f�nʬ6l�vS�6M�b�rp��	�v>����B#'���'.#�0��Mcc������rD��8Px?�TB�˯$\c�� ^+W�>g��;��
8��6f�N��R��Ĭ�!�`�'�듼 ���r`��#g�(W-~k���@7r�f��^	.�,�rK��g�����x��lJ v��m�4e"�>H��*E�w_11�9<�)�@���#5N|���Aΐ���I*y��e	-�K9�_ڤ�"�[W��h�Z��� 3p�H�n�x��������f�C����B.�G�/���9Lo]�cwk�M0j6SUt������益M��eo���/Oۦ;I.�XZ��Y\����g�>��C �����טJ��鉰#����:�X�鷙z(�.�z�_��mB簫l��0*�7j���_���f$L�t3D$�d~�������g�� ��c|e)�����B�=@���1~�Zw�������E=��:�����š���W�N���b:HPk�#�/�j�ȼ���_��?��Xd�V	F��ݒ:���a�K����ӹ.�VK�V"~���NR�w&7$�f5D�I02 ��l@�gU��JF�ȱ��)�Dg�9`�3x"����T��q�*����=��&�?c��E [�+��Ch�Fd����pg��M�l"U 0T��z�
-��3����2]�S�k��y��_�wX��(��F^���sT�3�@�r�ps%$�^��!��	ߔX]J���#"��P���R�\��|\�X�7�P_��\�Β��@�M_,�"�.����4� ��)�P�^?��.�x�i��i�ZAܩh�υ�J�p�:�������T B�C湡�,�Q���˾�� �SD�re�_C���kr�����ZD�LW����%�i��Bx�E�Ipd}�H��ѡr�\���KE,�����Qu�w��PFzːiC��Ղ�(%r�jP�-�����;m�1Nx�S<G (|-� �R��ܼ"%K�ȕ��4�c�	n�2x|!ە���n�R��B���pT������mGUwi
B��XX�,~V�O�LO�^�YK � T���tP�vM�UWI<* �ٿ�܌��m6ր蝧Mz�� 
����h�ȩ���q��v~�$hݔj��u���ݘ��|����U����{�B���4.�rT��]XL��8�����Pn�3j�,]/�+~�$\ɣbZ� ����i|��P�#"�13]�{�Ɨ�Ŋ8uRW<~{Ƨ�J���ڸ!:rU�i�'Λ���u��N+`犸'D%�)#=4X��`�{Lp+����A�7��f#��ٯ�E�k�7D�����R�����K�_@�Z�|��\O�J\�^������[�'y�������INx҅�V�$Qo�h�hox��㬄:T}�-�CEwm��3�{{wk]}�3=: SJ��҇ӝp0+쉹f�N ;���Z����
;�l�@T{����em�_%�@�,�A�]?��BCIq�r�tt4II���B�#}�O&���릱�����|ym,g�|%����ξ��mh�S���w��,!.�EMf)����K�^�����X�@��,c5�f���i}���
�a�+]�e�JaqS"EN��8��t<�������*WeԻ�]��Њh���ٮW���zh.�.Z��Y�I����B����(��A1ѲY;��tl>^�[�E��r�1`*nC#�g��ї�|i�I�է��&�\� H�!8�-�G�Q.U�i	z�� cw�K��>���z�ƥ�������[�����V��X�$�Q8�\SA�Q�lն�Wn�+�3����OxՉY��ͮ�u��>B���S��@K��ِJ�P�T�N!��ԛ�U٩�}nԊO!�g;�[��l�zZ�h��}��Ԇ��6��kf(ĢO��4��6��U7������w\����ޗ��賋w�J�k�O����9���g�}����.kZ~;eH4TP�j6�#�4��U3C� �Ɨ%5{�b���y{DC��;�Gy	��
��*�e���V��X��so�Yۣk���ӳ-��]��:Z�8C�G0�D �pQ$��ڴӻ���y �<V�Ñ�Z6=������>"�8����Ro��ˍt%L��J�5}D���8U�R���,(0Ys�����h���o<_�aE<x�?�/z���m�jɴhr��S�;�:%��O�
a�A9��&����E��,P�3e����F[�fJU��QW𳚛���3zp�à�����DT��7�����Z��Ǹ	�&'i�O8�[3�����1�8k�ܶ���j\�H�����x3�1���^���~Y�����(��;�jQ)��&�?��{7�T�3�?쬽��a� +T`��	,�睙c	�Bd�aq��H&^�z���{a${N[�`��(�>'���Ny��n1wB��<�lͅz��F��\��P�W��D?�g,cR��JƂR���Q`녺�e [S��I���a�]��}k>��Vh-QŒ�͑�@���/�-�a��@�4<XԔ8�i�����t��d�Cb�.�r{��n� �#�i��/���#����;�R���6ŭ@ZQ�є���>o�ۍ�9�e��ʥ��9)��%MƘ�F2��F7n����D�V�����+�~ެF	 ���u#��Fj12C���kԟ�WQG?B������课��:����&F~q�D%7] b�@�o8�z��?;f��"|�g�R=_fگ��nڠ	�7����w�󤅛"r���r`�J�	�]�)	<mѳ�2C���a�޶�9ʠjX�+��G#���'�Ӫ���Hn���`�N���
P� :�O�9k�
�iO����U��E�
�*R�4CeЂr����C/���b�>%���R�)�d��
�d����xD�27��Ҽ��WM��$�a3B(Zr�p��)"|��(,��� V����psi�#����J\�ʛ8G1�ۊ�5�!���#@�;|b�9'��"�ᅱ�	D2+�wG��Ǜ�ڼ���)�)�!8� �p��6H�E{j�A��CB���A�Z=0wX�O߈��8� �V�!���\����t	
/,�A<��v�]XӅ`���m�Y%��9l���FӘ2��U�u�T*R#D��#ʲJe��o���*l���N�"�7��#?�|`���b�L��o������r�wC�۠ޗxB�E��_�ӵ{�l�^h�]ۺ�}dKڥ0<~L��t����l�A�k�*h�s�**r��=O�)��r8���h�<��C�+l���ۣC��	|�r�N�S[��<�&~�,lбek5���
��5��s~$�A0�ؑ��K	��I9T�8�=�ֶa]$K���^?d��.{sRxBRQl��>�s1X��:��ɲaҭo3����g���������˙'M��>+��L�%Wn�kZ${�i�t���Bf �AytiYy��Q��G�2�����eGm�G..K*�A2̸Id�S��)7��t��ūq�Ly����'R.oR��a�v��r+�K�T^^ە.2�!���0���N���Ԓd��qN�r�h��H�M5X[��P1��C ���W,t�ŔއŠ�Q��=�ixaE�!���`�4��{L��W��~�H�����U2�Znw�͂�njG̸&��9��I<;�{��}� 0+�C�����y�I�tZ������h�r8)}0f���Xvh� ,��9ܝ��oVljI*�(�;�����<��a��{�K��J��eq>	Y�b�H�X3y�7��`�\|@	\�ci�p9��$_�����B�h��;�+���K*!�bq]�h��n'9��lna~�2o˙���$jo����Ѫ����Uzǌ���;_ [�d�����u���ϜӪ�݈c�-CV�uL�Ahp��>f����n��F�Z�S�5�,oFR���-.*k&�J��>vI�͘�@�у�vr�8�$� 0N+���2l���J�A{��ma`�g �=pr<)�Җy����@�̖���0SA]R�x@�&��"��^ ��s��w�겧QʌsJU�RWol`C���S*ioͤb Y���S����(,	�;Hv�� �3kCͯ�!��Z��K�=m�U>���(���� ���ew*�4�I�Y�vo�*W�o���|��wEm&���S�fد���eQ��/��5R�S�
\��s�m��nnR������<b���]������>ymTؼ���n<��zKI=<~��h�=.�<�y���/ؠ�w�m����G�9|���5�'Inu*F�t�_�����`�=��ޅ<��z-g'��|��Ml"��l��P�>d�q-�dg��f��y���
1 �9��ʓ�,��R������]�u�I�L ��ǎ�goXrI��	v͑ԥ�R-L7/)',�w��Uw�w��_`(�1H{֌�i���tr�:��<966#�߲ vPv
O2���uuӫ|�лja���i�5�b��|]T#�8?���O��9�c�[t3��
�7g�>W��q�:T��*�Sx�4��R��dV���5�Hv�)<�(G����&��]B��Wx5S9�KP�5S	�c�5�1�{�AZ�DH�\�@���X\ãH�چ�뢙�f�k�� XD�r�a����.v��Fi���x.�ɉ�d|�����T���2,(�rє�Ҏ!Y�������n$D��:p}�d��V�����J�H҄�C�!�!��&��ǖn���]-�_��Qb��J'��
�)͖��؍@`�M�w��ԍU����R�DG�������<���V&��ϓ��T"sq
�~�@��E�\���m涾`D�b@�i��ʊ#�u����p4;�����*#p4�����Ѐ��� �(���qT߁�yzu�M�w�|/8����1�y�tG:��4�$3�n�
�X3�Ƥ9��^��/y�C���Р��$^����=:�B7)�j�f��_T�W�G�Ñ_�^����}�A���3���׀���+��Я3g�L�!�=��uǾ|\�'�1�g��1tR�Z�P�8i� ��a���B����X��"��5��?��~m�#��C�8K��(
`��:e%��cF��8��� �'��d.~߂:�g��-��~d͒X�����n1�hp�D����d^�d�cV����K����p����.L�3%Ɔ�s���6��7��1�����/�����|�sؔ���A�}�O3��cN��Y '���qb�$C4��z�	��&gU�_�mUܼ�=�?���l���`�o��tNaf���u]�����.��ޅ�:n���L��9���5K��z�x���O����g>�?�)64���!�Kqr�j�'U�G��"5�%?��&��Y��6t�G�#	ػ�'�B����_��"��lpD�"�u
qg[�z�I��.�<���8�$��dc�8r]PU+��Pc⻃-��_�� ��AHځ��R�h�]�$�莠��}����8W�0R6n�K�3�M�]��XXvפ�a>R�@���C�V�'��kŋ�p &j��y��߁�o��c'����������c?-�d~#�(y'iͦJMa{���&ٴ*�j���zs0��lxm�ܲ�#Tj�K�xd���Ԛ'�V�_ü��փ���^XD����4�m����zW�Xp
ͧj�;��)�����f7l����]�
��6�mS�iG���E�H��FH.�CTTn�c�w�~rʠ����Gq*>�?�62���c�/D�� Kz��)���L1�$���#��G(�>�gZ�xV��B����5���T�^ʉz(�}�J�id-F�&,lУc�.,�!���WHݛJ��1��G��fp����s`�`��`K4����Y �"Zo?<�dDK�o�mKV����F�i�n��gsJ��<�*f2���SD$����E�n�1��
h�&�g�^יdR�[��U�AU�M�,���C+u���:���f���+l�j������^��tW|,����� � ��!����c��籚yU`�ˍ�'_����NO��]LW�Iwjr��c�g4���+9�\�Y�cՕ�U+��qb����>)��t�.<d��pch�bO�ZΘ���iF��H~�	,��w�9���иz%��!{xI^�BET������Jqp�i2`y���]�M���E��U}j��z���c���&n����� ro��_mL±���HLϤ�4���m䈠NO�2k����.gs����B-m�(�T��0��FDwH�6�q)��������2����ЩhxE)?|�`|jɈ|'���/٪v4^1�B.�p�2�P>M�h�-/K���6.g�K<��ρ�g�K<��e����x��9����5���`QSvF�2�r�?���0�͒���� �2�'%�E���/�X�"`G_�P��][�c����J�/o�����yD�+^��NrH�hZ]1�ùSM�A��^g��� ����\Ć��\�!�Q��$�R⒡
G��wnp�D����7b�'�;��s�T�"�i��u4<8�|��틝�D�m�vh@g�*�Np�o\�ѐh��X���0w�m��e�Zk;�Z�qUQ�0��b��Φ}�v�9=���y͆cF�	M�rR�����<�n24��K2gFn�	��B�>� R�q(���g�����{�T�.z�+�aB�@�d#C�]��ܽ����Y�y⹮�[�r��F0��|
�P��O����g|ln`�y�N�IC&ײ�@@ό�Y\��U�j�~��%8�T�xs{ ^�m�e���|+9�G��M��rN�����,�0|�lﮫ��{*��+:����8"�_[~`<�L@�niJZ5⇌+�6��C��������i�d���ח�Oe(�_�س���,�v��@�o(����ϗ�2	�~�)A�� ������>#{*�?j�FrV��D�G�����oh�����:�P{�5��}a�CwW1R6���W�)T���㱍�Zc�^K�ޅY�*�I�m�@��H:�� �T�K��{O:�ч��k�B�B'����%`�I�F���Jx��NΪ<�3O񤺃-��u���*ꆚ	�00�P o�A
[���)3B�|�Ӆ�^��Z�"n�a<�~ZY�lNĭ-��P��,��n�Ӑ���7ҧ�����&�]���Y@C���Fc�������X��y�N�`'���r�xX:��4�@q�:��9r��&nunڔ�?2i�?�FqdޫA�k�r*���I��-���Ƕ�m,��$�^@p����+�ԇ |�]�hU�e�E%�L�lݟ4�4��4���LHv���&-�v�8TB��a]������0IN	�ss�G������3�`U�cQ�"/�%>y��w�T��*�85���nx�Zz �e���W`�@�Uܤ௩o��UW�o\s
G�Ř=`
*GK�7vl��1��3���rPu� o� ?ਬ�hY����١8���2��\���1���p��4��v��?��Eژ>V�2k�}	b���ƩI����~Rk�~A�ʛ�7v_����a����B�K���ҵ�_�Te���[+C:�^�UC{tx�,?S�%�➽%L�yBU��𚚏<}�zS���,�V"�V�c�*,��D�w��<��鈝4�\|���.�ܾW(���%�6ݍ�h��8v�ޯ#����c|)Mu �m��%ZC�`��=1����*�V�n���������ndßb>*�&ˍjξ���W�:9Ź��f�Q�Su�8�vN�����x�7s�	^s+�kat��/���dmC��%�_:n��%�C/�9�*�Ri]%�w^��<h������А.���K
P�� �O����"q<2�0V?Ԝ6&U-�� � $L���џE��c Z��S�M�7�EA	��}�˜��4�T�?+G����u$ ���`�z��B�Z�@����3�3����8�S�D�ǳ��X��-�J�"5p�F����W�A�{o{q<�%������hl5�Q֘-%p��]N��F+2�{���I:�JhkU�0�`�:h�YM6�+��qS���W ���xI����D#�}O Ŋx�f�!Ź���
"�k�Qp]|E!��tI�I��K=(��I�����JZv�v�s���ٺ��ëx�_"��w
�������m��Z��;�3=�&���+�;ٰ�l�<�h9m����tiO��r
�yG޲��D�Mܶ� ����L�~��@$T*𤍕h:�+"�2D�U��.�0�-^n����5xi5dN0��0�,j���aY�����,w�e�qR�%Xc��CK��
�,�6�����WΪ�����%*�?��ke%f�������iMy.�
ђ��h��u�?���7�'���uͼ[�ε��A=G���*��!��2У�D�ǉ,�K ����(c3X�MH�f��g�}q����d�<�UR��K��qP��vU0z.b�0�+U#2,�;+����6�!��y�����r�}r y �[�`�<���qgsi�3T%�G+=��x�q�^�c5��x�`i��/=:gr�5%!�Ru�E�<0��Y	�1-Ӫ& .�4�O޹�iӞ>� q��9J�|�	�W^�"�%�͜&FB��������Q^Jv�b���~M��|?=���τ�Q���	�d�4[[�iĊm��&=�ӱ�h��G
j�Lo��4x&@$�+r�м�
�r�LU�u�z���NZ3����j	=�Twa��&��k`m�!���.U����*X�� �۷�X��sS�ډSi��)9�[i��x�	�vO�Jt�b��ޞ�e�����!+�j|��%��'t�^�#DR��O�=�I����R�o��n67�S�����W�]�A�������H�6p	��C_cE`�Z��,�����5V.�.�>��T�:��"��W"���/��$�G �;������D-+��;�`E��$/�vo�P��"��@*,��8�iI~Zb&��cl�'9o)�.y�.�އ:���Əx�ޡыn��I8�Y�-�,��4ۏ?7R$a�b*�m�e
H`R��]5ԟ���28�����[-����4Y���3fw�0�j��W���L�o�J����{
��~�+|!���X�4�����1���Ĉ��Uzl�᷆	�?�fJU,k���_a�E6��	%'�X1���:Alq`��ҥ���R�kY�/���M8"_�,W�ɴk��� ����[v�_aX�I@y^à;�|���Y\��I�#�ws5�ҕ�W������O�����!�x>bw��h���:lƭ$T]�J���N�v"O����Ȱ���fKW�*ڍƂ�lHԷ��P��6�/�{?cz�NGtM���`7O6�Ncw%M�J/����?����Ĩ���E_W<�"���t�`�5�u�BA�ϭj������ n|�2�
��N�,5pW�6��D�6�c_�Ts�\z>k�b�5g�ͱ�(��@�&�[���D|�3��3���x����9�*��*dv w��4�f7 #�w�mSB�Eȯ`�3�Qp$��)���i�8�Ka����SX[�d {H�Ҥ�!0�	q��h���^4���l�=9��Z��tOrOxɧG���t��,VԱV9�ߎ����Ш������8'��X��X�-QR����|� ��Oj�F �ǂP����w������b�#�����+L��`�t$m�Y����5�ZF��.����:�p�W;>:�xn(�ڸMC�T��&k��czQO��A���Q�*""4Bb�-��ʍ�zPU�b1��~R�P���7k�^o��C��_�Yl�����:�����[��z�V��P��ocg�MK���Y�e,�{}�j9��7B�����q�HN�7>�x�	$���P�j��� �//̽Gãh�?�ݥt��y��Ζ�ݴ�\��zF/��u�^�j%I����s��f%������V65R�<���>�ܢ��z�� ���Q�p�(��P�D�Iy��M��[}3�h��֠y�����M"ޡ��P>�%�05r��^��P礐�w�K��Y�����A~���8�}$�z�d��_�
^��ږ�!��) �]�V8�V8WGm�������˱�y�s;�0�ǧ���&^�y$@�mJ����OlQ+͵�y�1�3��؁w�݇��e�v�C�[+����۟f�p����C�GHM��9k��? u�BEv����dh����@0\<�L�a�S'YSDk��|�S FG�T&}D���"+�},����҈a'���L���Mxw-r��Bq����!�>߸n՘��;�`>U�;�2Ö`{o��1I��K�"�����z��q�Q,���e#8�ҾG��!��(�k�*�B�U2��+p�AF^P��9��r�����͠���I��3� ǆV��iRq�x� �k_3�X�!k����d����<��[J	'� $:K�O�����/��H����p��%�+�1�M�"��zQ�W��� Cs�0р?"]tX�w0��>"���4�x��D=�'Q����ʹd��J��ʈ��)to���vD�y�:Y��t~l����<�D�6�\��U�5�R	��^�����բAG���ۡΨdT��y�O���VT�D8�cb��	���)x�0AF�k��;��B�W�	�])f������W�v���S�śBl��B/X���.�*�OfK'A�A4�$����h��j��g5�|����t��[�ˆ��q"�R���z��b�l����/�!2ء�w�"�L�g���xʉn+�(���t|��CO�n�˂����lh�͜65���a��e�{[T-����y�u��{>h=_"�����PD@�o�>���=d�J��*8/�����}���G��ڼ�"�H/b��Ʀ��h���4tyK�͢&|�ՖhR��0�Z�v�!Z{Z���婘� �^��+��[՜%�wA2���MQ^v�M.aK$M[��<�#��e�	��y��z�ሎ����P4;���֒�m[�Ļ[�.,!���?w��`�!Zȯ}���P�	�E.�ű��|Nᧁ����E����:,jϜ��AƄ�b�v��q�]���?A�hn�$4�;�sD$ܹ�7**�z�{�wW�vD,����(Wm`H�>�*�Ȭ����w�H� �A���%8i�E���7ݻ5����
F���ٓBKXK����ȗ���Yu�����)��@`^Y���9%��m7L^[t�maי{��D�>R6#KYo�	arfN%�\�G|?g��E��,�����Ӑ�A��[-���ۈ�X�6���I����)�/�����#���4vtk��*On5C��w^��A?��Bp��s���V����|�75O4�OA4:�ðƴ���I��'yuA���/��̖����."��c�Ó'�v�M��MVݪ��bb ��~�;P��-��J0��\������>���M��[�Z�z��n|�=/�b�J�aCF�L����VXPa[�Si�!S�G�AN����t��^��.�4x�o,>�_����L*��A�s^���r�װ-�h�H�K�#�He���,�<.i#5��#�%�o�ₛ���ޕ����?���va�[��	�=*�ˍU-7�ώd2��9G;�6Pw �; 2��iE��NM�K�H��H~�/����dP������m�I�yט��W,'�l�M�O��W�QmPw��-���X!�|Y��<F9��E�w �$�o�p�GC��4�G
�K�+�uZr�� 1_�;�OS�q-�x��֗�&�$�Ϻ��1�=A���gA�F	�0ˉ����#[J���^�Ӗ㶽��[	6�P����ݡ������$��rQޯk���wNTD���q5����p�����9/J�L��nk��V.9T�i:�L`�����ǳM֣8����O]~�E�4S��.��� ��!�M �����S��8��klg���5����?_*��5�t��n#N�{wAΖ�fV\����Gv���^;�`~��_�bɩ�DdO8㪻��
��@���4M��=�*͏���  ��LY����7��4�`��E���r�*��0�^�M�࿁_b2�c�d麫���:ek����xԩ^��7=�J�:z����걻��1�G�=�?��̴�v��Oq����%��Zq�bE�̃�l,γ�b���+)f[�����Q�����*WHW�F���Ą;n ����L�e��&���𴿉���y1O��ׄ\�,#�}��ڋ�kh:�\M7~>)?p����c��ST���%t��d�i�J��F��p:w�\dbb?����F�<dZ�}���Hf�/�l�k9H��y�ۂ5*?#�+�6����O걫	���4�Te��)�,@�C.1�3:�h�,�2EdsJOXP��I�a�������<`�4!Y�ZN���]�Mp&���gLIL�N~�r�C �C�$^��a0Q��u�Ws)��j4#�qd㆞%�/�lfG�N�'����p���鷭���(��@O��93�� u�ֵ�i)�z3#��C�ͩ�k6��qBV��y�N PDE��_6�܃�ipP���d�47��3�f�O���]4�'�6N��Z�˟p��?+.���|ՐKG�3�"*�M��������1Fvt���j� pɉL�!v5c�BCV�>զ�ɤ�D&;G��Y����D�V����jș|����5��!�\��Æ�����&#g1�9�Ns�%m��-6�}��0�d#i�!��_�` �v�Ҳ�r�g*]>�N!_�a3�ʫG���~H����8��]
�V�N��(�SI{��u�6�3������󇮆�����C?5g���;i� 3�yS�3r+�^���W\��V2m�\=(;