��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(|����	t!����YXRe�������U݈�NׂI��h� cw����X�`��\���� �o�H�RLҹ�%��!��*�}�\���&�!Ԃ�0�K�~�B&�p'�=y�wV<'���PH�y\�^'��Y�����������D�x� :
�$�<�W�%�������=\IX�xTSa�n���3�q���$��H�k�X�������(V(U��L���ٲެQCE�v�6�m�C��7�䬷iW�E_߬Z¸�f��G=��E;��Qc�dg�clE{��#�c�T��DV3[�=� ���w�	��,���̏��i�׷�^�v�/��t�rM#�5{S��pͤZ�66&-�º�E8��GhE��Z ^����V�x�)I(���y�y�*����J]@�r�������n+~]��k�b|6� Ӑٿ*)L�4��cx�/������e"ѝ�1
@���#g�G���`�]Ϙ@�JZ`$��᫯b�Q"5���E˝�_E�����l��o�^�ٵe�h=��\��Y��e!%Ɏ�A�<Loӓ�ZGR�%�$:�Y7_�HB.Ɣ."��X+��z���d�'Cř+\@� $�M��gƍ��D���$��-�*Z������F�{n :����Od0����
�F��@!����<R��5�U��;�7F%m����<w���C�j���򾻐�{}�D�	�'(зKz(�5���1˝��p�g��~w�Λ�a��Ik�m|���;��`H�2ބ�����qP�|���hC|nFj�]'���e�s1�4���{�s9�0*�Au\��}�Ky/��u��L��2��Z6�d���������`ZP�c�$WG��$a�����,բe����o���.���rF�,���*\�U̦ŲL���(�d��Iid����V�nL�p#� ���v�/�:Go�g<�"�y�U��I��W!u��O�ܭSQ��!"�
��øt#���ږ�F���U�C���S��d���>N��v���iv��8�3Cr�@��v�ȩ9/��kJW:�	k�j�f��蠍�En�dq�o���Xb�1�JՊ�0ꍶG�� �Ū��{{����km���li�Ƿ΍,K(|4�cNWF��#�)�7�����\�àm����m��
p� ��;؞'��ii�z�Zy�EM��2t��F@�|1��b�?)3�i��5��De�&i�{��un�9�`�7��$Mګ5!���MP�����G�Ɂf�p-
ވ�X�~�$*ϊ���{�\*x��ș[�5���h�1>�r5��*�R�M���Sk �0)��d<����B�v���Wz f7�1�	�=T�U{E�܂.�����d���13l��}.>�Z�������P�ߟ��*���r��|D"^�+�ۄ�۱����tZ+n.�a�]�2Z*���K�ՒB9����C�2$��$WE�]a�z��Mb��,���j��!�|��չ��z���?ԥ8T ��#��������
�w9,�X����'βz4_*�S�*8v���e?kΝX%;�/`iU�޳�g��	�`ܴX�T���Z�:�jjZ��k���"��%}�����(�d��!!g�%����F�^�v��o4��z�t=	�����:�H�w,��(37���+/����}'�y��pu�m��X�����ʄ �d0�ܮ;���Q�D9�-��خ0�y���6�Q�x�8J@�#gM@�b�{��łzm�H2��؆�,�XD��j��B[ �^�rY�N٥pa��J�$Ee���Q��Yy���Ke�U(��~�'�<|�:�ά�~(Qq�^�3�B}E��Aw�ΰ����I|��˻�0�xp��8�zg�a;�{R�yIw�*L���*MCW�] O:���(?1����� h���2�<%���@΃t?��AQ1f�ۆ�`UyE (H\P�����M;���u6XPV�lNV`��2GY�4�=���hWO�g���O(�I�3�l��%��� ����m��P���ե����f�Jm�><��IS14�7�H�
-���Yn
���7���c!���-Q��
!�Vl's�Q�$��J�W_�M�!���ܾb���|q<�[�Ч\�>e�G�����-���+F���`j�|�Il���6���əUA	V�ߋ8N\����F~����|y�2'k�jbO�����EςM)W 0HϺ$#����S�<��7�EYY�3�Od�ܚ�H+���GڤW�ʙ�>�h�nm,n� ����+7T�K�&�U�,�w��`4t`pA���D�����yϦ���q�^ʋ��%�NL�+��~��d/�����>���aFy+�	�8kFddi?�C��*S����V�;�L1�Ԑb�MV�R��$�k��e_������^�q!�%l�{�Qt�5�$��u��$�M^���j��,�4%����~�n��Va�{��?����a{omZd�`�uj�r�x��laO�C���q��(e�w������*,���D�!����K�
m�;KV����
�_�v~WD͓�q��a�e��̧�G��Z	5�+����
"��oJ�!l�\+�0C�xt��4d����P"��rz,�9]}ͮ��ڲ�"!��^>���.▂��?���2�9w�+���hό��M�T��nw�-�m����1ed5*�h&>�Uew�h��J�j�(~n�����|qF�H7���Aq����[<��2P}qd$ۘ!_b]V�Ͻ���ث���?���,݊+'�		;�[V��j����c�Q���-�vOݬ솫 �-M<�pѨ�9 ��p���� 0Ho��yd=4�x/S��"��w�o�u�����.|�J�xvŪ�B=��%���e�����&���;~��ub�+ظ��؏�e/�/g�&���A���EC�ߩ��������3��_G[��q� �*xe{^�̤�(�v���vۈ��lE����p)�$�1��R1S��ǧeí?�y`��e�d��k9{��ۜErӈV\��YD�;9!��=�,	��� ʷ�T�Q�fU��4�x�!hK���-�#�u����i��*j'&�7Je�s�_�����֡X]�E���fQ�XHVp�"����(A���F��ߠ����sv����_+]P�{` 	������~���� ?ǭ�V��E�j��IbF:��xBmKE��Դu sJ��=Gl��b�-	����H*f[��;N"
?y)�
�-�շ�����q(��=��h�c{�JU�ڂ�0ʔ#�*������1	op�g?��ɓ��v��kfcp����l3�BG~́3p~v�5A쾩i�S<a��45F~��qQ�N$�`�ˌ	k�9����	�蠡6��cUf�hGWl���F��5��'5!���.F�J���+�h����^�wr
ޞ��AG��&������Z_����z�k,�D׬ȣׁ��E��k'�#���}�o0�)���SɉC��,��4pw��Y)���?!��+k���&H0'ӣ��tZa�X߭|5C�13� v���x�*'- ɸh��Ww�W��@��>p0"DX��@�r��WX*&M�����N�묰��-����D2����!�C�Kʣ�ƾ C`�۪�2K|��Fϊ-A�D��RA;����!q�"�M�QHXb�p\��Y�1�����"�昸7�xvhͨ�%Y#���6�񀊓<�q��:fp~h��M�2@l�;�Cnb���BMR�Φ�����#�5���,��p"i�1��!�n@� �ȗ�M90���{�)l��f��ǆ,��f>_̍s���ãs�@*o�>�˭� d��䉄�����Fu�E���^���?�.E���?�� "�`���q���"]��#rRU�������3͈CVfTV+���T]�0��=�1����Vt��\E�,�湼��7��ߨr�̻��w�\���m��8ʜ���(z���3��L�m���:Ҕ�m�Ͳ��^f�npCI���]"4
�����	?E����_���w����ߓ�����-�~U&�|a�h�Ԯ��F�?6稠�Y�"%�pQ? ͅ����Ad�-�s̥�9Ԋ�x���t������ж.A�X��kI����dT�H���06b�k�������f��<N�7����r����x�6-��}�&?����^r:#�S����8���$Vʁ;�.�9�b d�9.�r���@�&�}y�%��@�ܩ�i�/LS"Q:hhz;U��/;;��7�_fZ��M��ɖ�P�qdA׶(��W	x����5��tOe���ǲ@�bLC�`�y����	�_,�P��t
̈́�@[O����U'�0��G=�b�%LT\�
���m���/E�"��_c%� M�,}ok��/ō`��l�)�Ey�K��0�u�Qȧ�\ʝD�������Dd08�
��<���B*˂�==R��$������L�+ɛ��<'�qhAJ��t�!��;�a5B6���x��phWz��rZ`���	����:x�m��5M*j�J�Zl���;��{�"j[���:��6EL�#���q��F-�S��ڶ���4�g�r]�(��7�iRW	��@�z	+��d����P��GfeM,ꀻ��`A.�����4(�����RK̓�eG��9W�[OΖ�c�����0~NZ�ȫ\O���l��@���FhI�;PN%�-T�$^��h�3lyS?�!	������HU�ՕM�8�sH�����K��R��Į��`�0 �J�S�}�'�!���η�+]�fA$	6�O��쟩�4�J�?;��-�:n��n�ˤz-�*q�
	��QNr�ō��������f��m�l0�JG�Ǣ�� ����J�BZq)�w���R�BG?1H��G���Y�q���K#ţ�1 ���*9��kVc>��;�'�/��azles�dDg�ŉ���b[��9�#�,J�O��(����uz[0ܗ˾�L/���th`�ogxE�X��R;	9B�p<�-�*4T���˗S�>"��@���;Q�K��m�p�X��3��Y��]�^bY��V�{�vu�u8���F��B�_��*�x�n^y���������Bh���2�#�0��W�~�I��9_�"Z9-d��|t!S�ϲ\+�(�s��Fd�Ԃ��4�V�R��Q��)�	�M(o�0�i:o�+��Kx���2��g_*:G�9�\E�\��sz��%�D;�oaSgP���(!��T*_?�a�-��a������@ƇV'��G\�$��ǎ����U��jo�DJD����	P�ۘcK�8$��G��a�����l�36��ҜvgP�%yZ@�r�6�C�^��Oc�q��q��?Z�;�0/�?��O;��E%6�g�9�ܘF�z*�N��~���߼��3#�V����7�X��Ƣk3wߵ��s�:'���`�	 2��.��/\K=s�;��.DN���̧��H ��BX�Bj^}I v�X���yҼ���a��ƿ��t����,VSSVG�d��������#��P،�l�F]���!cO\}m�b�Υ�.[)H��"�6F�ӷ�"�Ux-�[��+8�^�KJ��A!�Zmk/���^S�BM��3M h����e�	W����9�G�X���ʭ.���xN�i��������=6��c���yX@25�]��l�����晥g'$����?�F�󵄗�U|��쩠/bFX:�[�9�EE�\+��=�O_T����8*��v̪ҺG�-+�X���c�։Q�3���A���[�<�}Sp�r۶$j$�C�ܯ5�(ۃ�������e(�:³�%�2���}�дK�1J�y�+�m�}��}��݆��au�[��B>'��H��Jƺ n"=��GsѬ��[�L�ğ��j���)��d�EI�$�g�4��I�ba&�4Λ�"E[rD��4.��?�q1�H�Hl��ɍA>YVB�FԬ��@5����HP���ѓ=4U�4��@� [���Bpf��`�a����R֍�籜���n?�U_�t��6VS#����:L����j��CH+06��LCK�a�'�?��&:z1Qbp!U	��j����^Î*�����
�F���D>M��8]�xH��g.�Zg�Ȓ˨���ъf�=u���*�j�s�������<�X#���rr��*:9�]�q(�0A3ytm)1�W~j�)J���r�Vf�09��^*׎�e�a�'��u�'q�ղ���A��5��S	2���#B�̤$�<d��ĄguC�ʈy���.���0k�f`�5�����fV��c<'�6a�����4PӒ;8�� $;��圐�x�O˸���
�
�\��]a\p�w��=�
w���Q����FA�'�BK�3�����*�Ag鄚��J��8�3�$�e-~������ec������i��9�yX���ٸ�;RY����$�P+ƥS3C)pD&dB$���5��;1���� ��2�����l�;�����7m�!�?�a������