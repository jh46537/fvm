��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""½�c��ノ�!]&P{re|ڀ1�(=CK�{Y��C+S�� 8I*�oһ�s\�2"�^`!Y�XeR)���g���]�)!r&���:oK�چ��,"n� �R��T+���5j0z���u��T�ո]�Oh>mF�pa��� )�Ճu�n���`�-��~�k2��$� 'T�&US_;gn���k
C��}�N�����c�CG��=��e%���D;��)4�H�  t֘^4#�[I�fW�m��S�R �ne�/T^��+D����4���m���r�ر�b�W��N�Z�2��s
WM����'؞:�|>�Wp��fr��;p�@�		�� �y[�N|>�X_��AI ��	��wW���1y��/Yx����I�O:u�~��ݕy�g��[ɷ��,���Z7�UK���z�`�Iʬ�PR��=w�3|2ݒ,O���T b��f��CF�� {���,��	�����ʘc�)a���PYn�5`DyI�U!v{ZA C�w�b��n}#�/��Y����<=k_Y�EH�"T}g���������v��A{���C��NX	� o����:U����w�Y���x�'��~@Ls�o>�ffZ��Q.|��珄��؎3�}�p�%4B�$����͸��HR��V��p��\$i~꜊�\�%���H� '�a.��h��	Ť)]7�T;-و쵖_}|`CYǭ�q>a'{_��$�(t[�>��pN�9D���a����qP瘌�K}:~��S	��[�� �����{(�c�<b0�k��95�m]Op��Y7헔}u�0�o�-nB~i�ez�����>�ˏw�.��FI�H+{D�B���A�G�;���ԼD-��G��HƭM���v�t�n���+�ep���%Y������Aa�����u&h�R���W���D?+J:tȿ_�5ݑ�{��pT�Z(e(-����\�˄7���-F
�NH����2i�,-Q#>�����L8����@X7 D�a���K7`��aL�����`�V�<O���C"B�v���E��н�"J:ۘC�I�,���ε*����p��0G��:%W̨ɼ�&� C]
��T�KN����'��HD��͉؄�8.Mp��
c#��"Um�e\yj˳�@|��y�У"���+yd�.1I���v��G���|��釯-�Q��P�jk�#��$����J��B�\����GH�v�:�G�k<iy�e��18��\1�K��ٝ�A�fJ9MsE����,�)��9ZD�U���yLp��i`��*�̠.�b^���Q�h�r�\ND�yjL�a�N�N���Y�L���K�@!��.xP^.�J�T�ۀ�?Rs���W(x���ao2���`�/���D��N�S
}P�֑��q���|4�����(-*�8� ܎O%f����� ����sZ�om�-iB�\\�)ı��9��J�K5��,�MG�I6u��i8c%H�'����5-� �<OY>E�\m�Q<�?�N�6�8l��$�)����W��=aSKmd;�^�"�IHM9��[�VFlz�h*��ȗ�:��u������B�΍�)����������`��Ujv���*	V=�������j�������6T1�S�a�?sC��سoMz9Y��Lk75��q�>�{MqK�9�-dv1oN�%%�
��D��h�j�D֮�Z��u�Ck'���Ϧ��AC�M�AKCqȼ�����Kn�~+����8���垠OB��V����Z]�����El�_�]ߤ�X�ƺ0�D~�j#�}c!�˴��7����K��0�R�:��_��(��� �������%�;�)�X�k�DI9��=6�"���
@ H�O�5��k*y9�6����[�qß`�n���(��w�a[�/H�`{:e��%�Vk<5%kB�m�nn�˗`���ˆ|����\p����ݿ�k��@g�՟��C�h�|��p/-,6d����\^�����M)(��r�j2!~ )
�%�;{?q�e��!�*7���"���;Z%���Z��n�����wJ{+�G<X�Փj�ap��e�+0O�Kz_=썎
�y��f@YV}w)�B	��^y��[4�<�>-�1m��)���c��S�:��g�Br
 ����Jss�ֻ�;8�R7�	(���F���x$ #�,T�@�	�g5?�E����}��w=�we@ΒQm�OV-
�͖핔f��"��t0�0����apy��,�ka���&T�����2&���:d��4b^#1	�����t��M���FEc�x�}�ĉRe)��]_���IuU٢�ƚ�cFU�ǐR�W{D{�r�Rk�YJ�J�Z�K.X@xN'��zU�o�U'�(g�� �� ��/�l,� nbP�4nҿ�� �%�8%��"�T��
V���֎-���;1I��(|���Tޗ�) �OF�!b����ub��ɥNY3E�;�x��_��˝���M0�Îx�T�~pp� &v�C�:�o�G��G`��[w�k�Ĳ��;v�f�I�X� �x7Wv��:�;_��o	�2��ʃʳEɲ���MBQt�4�1�}�De|����>�Vn� ���?rDk�-1�r�m�䱼h<r����ɂ�c��gp/��i»�e���:��'Y��Є.@�+��(�HxV�rq�k��
�8hg��`�:f!��0�մ����תB=����aDV��B*	 ��������۱� ���n�ܹ�o��{�N���#�e�A�gY�9�F 〻��8=(�>8də�=b����Sɴ����v��XWL=T��lF"���������tG]^��jy��.;#c0%��*BG�=�3x��L ��d��ntV!XՖ��!lu��1$����N�ۣG:���-�Bg�˽"��#u�W�F�j�8E�	�W�IJ��O�Jw�o涄���I5��+��"�oͽ�ey=ƳXh�fAװť�A�jv�������;�E*ɱ��D�C<Cpo��/=�@����i*�z��|�H�d��,�H��kQ��
����i�8j�T_!5β�n�QM,6ĸ��`�s�I�7��i�hsx	�/_��o�c�L^BO� t%��&�#�OC�b���rs"P��ըP�q��°t�y�].I����8ֵd1��h	��C����]������.e0���EL���B���q�Gk���P�M6���ţ�Ex<��G���ѫ'�K��ƙ��EA$zcO�4	��K*��Fej����"��̨��ÞS$O��O9�[t�wE��e�]2cT�"�eI�1�.��Q.��FO��?����8r3�L�p��C�Q��`%��8�|�m��DXϧ���a�B]@5R�73�l�U�{�K�.`vk�����*�1� H����pyy�n��ٜHVFM������K�'a�~O����S@B^'�x�0R���"�B-�)���(�`#5�E�3HqPoV��(����Kf�~X�J?\_2�)���暋ѾxʮtKi��k�o<g����&B�ͦ:�ً�}i�яǇԜQ�̚ic5%�8xEC!��l��ʷp���yR!+�����a`B�<�_�W#���f�S���xa�^�ΥU�S�0�T�p�ᕖxr��;h�+E��}(�-��c��]Ap�8]�)�ۤ�%��d���B�E������S�6l�/��G�n��+�敫a��gE?Y����]�l#��z7��:q=d��du
F�.�2(/Z�e��s�+���.��q����'?��n8I��TdL����!�xL��V덡W���S��+81���j�"��T�"��x�h�?^��o��_yb��}q͛1���2��d��{fiä����r�@�� �2wT �6BB���)�΢$�nδ,e�͜���=_�q�>�`v�_Ʌ3Mu\�j���ў�b�2E�,�U-y
�ѫ�.��������6�B��ʰ"y��L�"��|��?�;̅j*k=�>]&���YVA3�oD��C�#�����~�x�{��BPwfƸ�ɺ:XR��0� ҷ*f���AjiP��"j�����Yp�N�
\��|�Tbؼ�
JC���F�Z�`C�^�
fh}+>�r�P	�!�4�7�����G<h���)���WW?�LD$zj�� \E���6j�G���瑟e,p������.�W���<���	���0�u��8�n�-�U��k�@�E�%����({֪f�E�0��|��p�U��d������u�����`9W�TkN�DUC���b��r;��lI��:�c�ѻ���R@07�0D�& C�5���O1\wL]�#��X#����ܻeY�ʹx���<]��8K�?�!����*��^i��r��E�g'�&��Pಐ�$A�$N�CX[se].��r� �w*���$�1�� ������y�oː�>�&|.��r��Ⱥ��nRR�fŽІ�.�."�	�	@����V�T52N,��n���CX�Ú�*�HA�TC/Hm��XPZEEa�/}|u��j��,�M$��	K���VTuU�T��PX{��oq7N^k��  ��E ��m����	�C1�׏�0���W]p7�²}�Э����e,��L�,P�v��$���
T�eK���@���i����m��%XR��Yu=�G�e�{y���)�7 ��ʠ}��ԋ�ޮ�R�$;�r�p�D�d�0\��%ਣ��4F�Ė���Rg���6������Г�Tݳ1g�)��0ng�D�[����$�#��xYl�s!�9�S\��p&f�)܅�-Y���xM��s`Zg���Z�+�D�	'��iv8/�OD��ck�"���Լ�N�
���X9H��A8E !�.*(�����ռ�tړ� �P'SWɂ��p!��E���y{ch�'�s/1�虥�|_�Ĥg۪A����+N �Vh�ꠗ��� ���~t��u��ޙ��#�s^��ZE8L}~ �f�ʸ5Gj*� �D�ֽD[@<U���
8��F-���g�_rύ�ϕ��K�c<O�j�(m�j뿬"��8�%�I���F	�ɱ?����E
C����N�|�+,�~s��o�����m2�1S��u�r|!��l)ݫ����q@���0"�gh��Ӡ{ٕ�?�����]�k"(��bW���VD:�2{g�;�K�e��ڛ|�����Q�*�$��F�M��3$�_"؄�:���t�,}�G�}��8@L�ȽE�e�=���9�!�0��Q�O��'�-V�G��-:O S����+�%��c�g��?i	����q��5�%2�{����*>'r'4��4*SPH�=^?iXV|��\qaIj]��4�h�s�"A�и(U��M����H!��t�{�~c���,�bď�.��z85��G�G<p\Q�����(Ԑ��{��( ����M��+�z�|�&��ȭd�00���?�F�^�V�.�ҹ&�(���e~G0ˇ�:�ʲAi�+�י�N2�k@ѱ�����+�|�l����%!�p�\����+]>_�]i�6�7a����"�Y���Ϟ�葩q��%��zڡ���q�ODM�̼��?l��52��g>T��փ�������.����3N��Z��3(�s���og�A�����]p��n��;k8^����c��]�"+%��)1�]������6�|��,]�{SV�I����T�f���t�V�ղ�e���L-�>���w���}��#p�����Z$��!��9��&Up����9��T�Y�Ⱥ�"�-!�{Z�����������w�z�\)����# �ސ�e��2�{ٞe�u�#"ǀ�a�		�6��F:0�nA[Y?�$d#�P<���1��x�C���w��#,�z�2���dQ
�ܺ�@,�
O�2n�
�4zT��j%�����S��ᯡ�$�����Bn���<�
V�ԋi���R ���;s�s9ɎL�;U�^�sٷ����zbT��5?��x�q2�F�,<���;7��&��P���*�����o�Zm��8��H���2(��ų�\=B�%˲�ڗ�XU�i��OJ(*p_Fh�*<9e���c��V�b�������o���Ƚ�����CD��Ѝ�gM��E��bu�z�����3 m��2m�b���j��c�����l��a��H��1M�%����`��ڜ0��~$�%���~��h�"�y��R��ps�N�N�U���D���\3�c
q&�{D
u�4�J�xu�mV+���zD�|�d� ����lm	���o�9
+w)A dy�l)n��F!7���J���jYdm'_����a��0��c�4abN���%������nW����d�s�[R4m�Q���bҋ�'��yJr۳4�ť"q$�Ϲ��T�3�
Y���Lq�ZU�MT$��U/���)7�P#ʥ��ѹ��࿭8 P_��l��.^m��~�?|���� ����qJ�s�4}����G��HmI�R�n�߰���p����v�@�,�������R'>R�lZ�:%�ig���x����5�l䨊����5�`�)���e��vs�2�W�zc�}7�b��Q��+�f!�H�7z�̟��Ʊ��XkI��f����R� �'���Y�������@Fm���Q�>":.?ͳ�zN���>V%C�����i8wu)��dn��;���n�U�1�!k9��[���hqKIf��!건�����W��1�1O�=�UM"o��cn��{�*{�����O�L	�5�$#�pF?,rhe���'��� �H\M9gɡ^����z��b��J���,PX��9�}^N�#��^ ���۷���MwZs������9�C���K���°!� �Z_7��� P�ЯO��pI]�����{�Cu��8�q��(<���/�-J����bk�@�5�N&�Y�J$2#���kڽk)=v�s�Q�����8Az3���M?�Q1_����%Su�'��E���j&��	�v��p,ڡ����Fl���G��-��A��@�j��@���n�:���?���O�<=O?��x����z����?�_͎*�K�Y�I9MH]��_̉��v����B�-�
����Y{���w�'@7�֟�D&u�{�f�[N��a~T� ��>�%�c�����q���rmo ���Y�k���X����-Lp��(D��#ߌ�3FS�ʆWD�˟f?�oz��5����G�$1ghQ�3��i6%Sx(y�^����8�Ջ]6T��c��=���e4��5|8�����/ƍ�N�)�%KK�+?�U��7f����~��}����g�t9��@���(%ve.g!?�8�"��ji�B���t�}O�0@�����	�3k
��ƣ���*J�W�T����x��#~���=�q�k�&��=j�i��hF��D ���#����Q�����k��h�����X�StdsՃ���d�E(��f
��d�23��K�h;`�K��j+c���٦߼k�*W�+�(Pu��A�X���{�Sd& ��lI#��ˤbg���!�'D��}��BK�`{;!0�W$��(�?���x��ˊ��l�_P���b��g���ޠ\����\}Q�N�N�R@h鿁��$P{�l{�����C�n6��@���lw�@N��x�Tuw�TC��F xy�:]�X������n���:��.Ni(�ȁ]�E,�l�4���H��q̗����c��Ǵ��w�W\��6R���A��h?-�������I���Nd����B䏑#[�ă'�ڽ@qL�A��A�<	Ɖ�5�R�8׻�-����b�.��3�Z"M���y�v1��_e>o{7kIy�oؚQa��D��������3j�������d	eR`�K�BZ��s>+��b���'��(n��jyOQQP+lY��3MB	 �y�A����}j�T�鞱|�	���q��@A����T������fB����t۞1W� �c�*���#� SA�ȬH�1�8�#[X�LK�P�� X�)x�+�v�z��/V�!�%�H.�8�!}O�k~��B���}M����>M��کF��_�8GL�H�4�e����*�NQ���4�7.������������^Nq~���|<t8(�����L`b�%�nGb��Z�m]	�om��1�����������\�Jh��8�e���4.v*g"��v��/�c:%<��p�߈��%�߃�����8���C5�P�vÏ�юJ^_L�9W��BQR���N�'��M�8��']��L�zx��Цol3k��OI����:�Z�E��Z�fpE����c�([l#?f4l�>�U�fG/�e|MqY؝�㳲z��I-�>LmTG4o�Q���3�1���x�-f���ER�3W��������"�R�>sl��m�����������y��=K�)���Ż0�VA�k^�Ov�m��ݚ��Ѧ����L�ڸ�v��[�-��2&���W�l���nOM!F�����L�i�H��^�7���y;�����"�N�	K£E���g�ퟌ� �O�	�J�6���f���ì�^���6����9���Գ��A��(��_vò�-��\�+,�ډ�،��Q�i������@��+5�f�$�8�m^7W�'��SNAW��n�=�!|]a[i��I��L2 �^�:i�� =�}�y�����Y^�������C��խ8�}o_<}!����yVyI'_�H$�*b��r#^��6�_�]�?/��sݚ�&����ZSQ�I�1w�e�Ղ���`vO�m{!O�G�*����H��Hْʹű#�p����h�#�e�3�s���yN�G*�����>L�X]v�cS�y�Ϸ�� :-٠��ט��ݕ��u�G�ي�^Ȃ+N��&��b`�j���`�(y+>-��K�UU��	0ð��6���:�Q�G��9�>q���ƳX�J�����&-2��3T��ɆoF�'v�J+����V��|�$�4řj+s�?�A�� �g4�>Ί��c����&�a7�dvi���?)ڜ?���	^a���}ay
2/�r:H\��Q������b+3��E �3�$�r�O��o،ovz�@1�r�)�k'V.��{"y����C����bL3����ުso=ńtc��F%gGP�aWo*�.�WEx�_�=�E������g��p➞lOG�[2yVv7���}�z�(Mj�퓯0�:�$��`�O	c)�]h9��/�*�U�n�N-��J4i�v{)��J],��B)�&QC~���xz�p�TG����$,*(>xd6�J�_ 3�V�z��v������<��D��ǥ��Kń��W��6��,�(��:M��,u8ԥ�j�gC�>�GKwV� ��G��fC茼��4�1pd?i$:`/`�O?V�Y4��l�Cl��M<|��"��2�8�R� �����u�y��R�'"�_	����sV:o�����Ⱦ5��?�^�.��6Z�tesX!�t4tT��Y� ��~�^�ՙ���vغɖ��9 o1���;�_��� ���N���M�w$����o��9�5)�L�\Fq���0 �H�#��¬f`4|zz;:W+P��v�H?*�Ğ���>5�����I��Gn����^�k��8�JXSo��A]��\s�^PM���}��