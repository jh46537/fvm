��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_���+�#�����u�a�� �E	,a�$�����DH�"|>/NN����8nz�b��ޣ��j2(!'rUz�c_�Z���!4N�ǚ���}(]�19��������ڽ������+��'״1'�Ozd�T�P�,Ҽ�ٓÓ[&6=��kI�w���c����'>@�Eż���٨�Ӽ$S�J�#�w��#���H�~
,e� RI��%�(E�/zx(�iYJM�u�`ۙ�YAmN1���,d~��g>�����CR��R�i:%�1R{�R+f�ָ[�B���}�>��Lr�,dm���q;��N�&�d��Q�'3�ʜ�%�� �^�=���Q	�gy��Ik���b��E�I-NOvޟ��\ēm�8Ze{t�U�쵠We����3�J�7:�ͧ�J�±���{��*\�H��<{:�٠�5�T����7��3�b�&��w��J�x��}⫹�E<o���6IE�ފ6�6$jq9��n|�"�f����6���F)�S%~ca���TP�JV�6���.�uW��e�<�%|5��մ���]�<��]��[��;F?�9�{����.�	(���{VOĮ��d�-�·
����~,7�}ܢޅ3��:>����.���C0�'[:�t�C���M����-���7�w�-��G fn����3p��;8��9G^.�����$��x�C./n�Pn�fXL����d�H�N��D@���2`�� j��
���/,���H"����l��Й'�>G�P_X��ɹ�Mng���+UW�����vр ��Oh������������_�<�2L��H[�C��GB����Y'�@������v��|w�cYpgU��]�w{pJY��V�VT��~�`�0m�(kSB��R+nI,�n���h����El� �V9�v
�,T����+~F@�T��W�x�q5�T��t8:7���hc2T���6�;%������ª_���t����Ļ1��
9�b�ˠ�U3��j�i4���v�bDNB��2	�ғi��eV) ���$��g�y:��H��s��D����*�:���iߴ�:u+*�h�Y�uz��2bbb}��o~-R8�a�EU�ώ^��ݲ�xcϞ�OܼY��v����q�~�j.�lM��t��0�����8c�7�4�Ǘ?�Z�5�F��9� cb�]��*��dy,�o�О�c7Q_��h57m�b�ꬒvul�2R�-̊a�p�8%�^�抈�q���=�[�~;%W�!vOɖ�M��@}ل�oY"��a���	��)��,����^�2�:fiym���ɺԘ�\���A�"ʲP5��� ����O�LQ":��,W<LB�)����|M���'(�U�	�-�:v�0�unjKו)�ۊI��)sk�	џ�p�-T� 0s��%4��!��M�r�֌��w�[��	?}��@�|�g
!c �J_,�������To���n�޶M22).�l�[�~l��O��w_ҡ��6�h,f��~�uI�I�N����
e39x�"��0?�V���*=�*���ɔI�-/��ߊ8P�u� ����9��|�C���si�4x>����qE��T��h�2)%�ZK+�j���s:E���\n@p�}p=2����Tb��S!h�?�����4�m�%��ܭ��NG��ʽ�Ną��qrs�z0��{N^�)y���(%q4U���B-�h@�Ys��ɗ(�K�d����w4K��8(׼�����/15�}3� �01�V����&W�����w������d5�*�TNTW�Bn1�2Ǣ�p{�e�A�
���ٚԓ��\?����~�Q��j),��1z;o���T7���0+o6M��P�JL�_�� �Wx�ě'l:�r ��A{���9& ��t�!YΚY?C� �/���!�6�R�7�p��v��X��UB*�#�`kɂ�t*��Q��S5!�(A�E���q?�r��=Œ��K�mz}�g']]��l�oRM�&Q��|/8V2ĝ��_-�����~/0�8��>�7�f�x�z�� �%ai�̫����X�W�1��������!�{>�_T�����f�h���69��t�E�O�����S�D����6۔�>s�.X<. S�E��O��B�6p��8l$|��,vK&Z|t�dQX���:r�k����V`���9�˖�~���,o/�����.)�>�g$�k�V;�?��ɘ�ۍ8<��=��k�Yl�$�q"���H`�-��ﵦx�kX������;��}�������dK�.B�#����=E�ji��-\X�l]�1�e�)1���9;�K6�9װ�F\��|ƧXXC��')GT�=�7�j����f@���P|eb��1�~o)���@�ױ4�Ϫ�K���W��������j�X:����;����a��\�%��w��yz�sI�><E"��wF�@�^��*s�ߓ�Wذ�,�G�҄�^�U<��k��n��8n���-���?�z���F3`l���gR+��r�c�A3+hB�au���{-������L!Uj�吣�|[#��f���L/�(��Y��}G����V/�y��*������&F�]�A ����j�@0��+�"��I�N�x.���>=��ق^�g��CA��X�ʔ���I��n#wɢ-��Ȁ�@���f�갬E���izqt��ew��s��3��\S��c,@�| ��2o�Ex@u���%H|��˦?&V��{LU�������C+�Xp��.�b����6�Q"��7'�yWѽ1�s���O�f�!��5�v�=�~�v�Z��ռή�/�Ә�i��W
+AU΅���9\��j��9�$�Bl�rᎸ�/��}D=~���m�����N��q=�~p\ �wd�ܿ]�0Kܦ������x{�qz챺&��^g}�)���8+�'n�[Όl�N\���?��$�l0ZG����O�����g?vbN��A`�B`0~I
`_�Kb5�۲��J����e�����܂�D�b4�ut����v�Q��?��5[ʺ�5���;�V )��3[dd��:55�o��t(�Ē!
h11�q�Z��5�}rU�X*�BO{��2�������0��2Ά����)�d0� ��x?��kU; ��5̤͒�Z�8۶�?���%i7�KJ�b`�K&�|J�@ϥ���M^�懫����5���6̪TZ��WpH-�[Qr�A�_z
���'�;HP���S�f�Um�>�eg����p�96�k�]�#�n���-��+<q��HcT�t27�.g}���ƈ27��u빸O��H87xZl�O�������0}��~!㝩���0�,_	��1�*b��g���`d���w�*��� �J��6'�<���|J�nRlr�R���_T�߾m�sT�J� ��4�6�y��>�����×f�S��ۣ�xKM�|�0���?���o��
2?6�=�4!*�6n�v%�ʄN��59�C�]?K��"�-���uwL�DP��< ù��(&�U', l�[J�j��d�"Y��m؏{�S��!y	���]�ukn��u#>�Ky����d��9��w?$�F�b��<�<a�_ �E;�b;s�D��.��e�9պ[B����m�H���"V�c9�����}I�|?t6~h��b��b�%��MaO���
�>x�V��@%�)OK��!(��^R�.�����XP�J0�O<�sa�#��=����3��dY�gT7��?��z�u1���6�}\�^x�wY;�:�<�1�;���|e�.e�:������A�$䂞����
z+����D�	.���}�嬰�u�����Sc��*az\�NQ.*�G��2�[�y�iQl` ;Ĥ�#���!�Ĺa��	A޷�5S����xU�N�3��Ic��+拊�f�_�����h�V�;��q������/,>��3mT	4��������O���d�VO\��؈��.V+Ѣ�KN_�T_8��n"�����Yv��ed��	��������e��Y�o�^�G�r��:��k!�[��hR��r��#��R;���j\qe��9��r��
M�)�R.�L:��k�O�>uϖ���?^8�Zj�({�i		�����~G5���0�ʞ��ѱYB3���/�h���9E�:�)>ֳH^��\F�/ȡU���1,��/%%�����)�m\T⧌��t����W�XՍ;���۟勵s�ݒ��7�E���	h��t�� ��sI�0t�~�6Y�^+��d��an�p ��nߚ������}��m����YS��#6&:�Q_WO_W��}M�}�lb�.E*�����_�+~���<Z���d1R�#�<�������o������I#�aV$� Z��R߆\�Ѩr���(y��j���/�����<tK8�\a..����� Q^���
��N󛙩���@�[�ߛ��!oD)K���@����X*��g,�`3ӯjQc�b����E�m��=`Ǉ�3gB�6�y���k�2�~�\��J5�1�����'x����ʹB��e��Ӈ	���ŰZ�5 ï��ru
����8�� �l���F����sL��K{)tS�@����A�j���U�������5��%��-Hc�l��$�>���v�&��^��#�S����P�e�!�ʔ!e�6�.�US3{�������e���J�L}Qϸ|u/�f��s.�y��5�O���V%>������g�#ڷ���i~�=����g�~����(�qi�\����?4Hk�Gf��ɾ\��<"��^�
�ӭ�0.%���*������ڤ�ܐt���T+g�����x�M�H;zVB�\�Msk+�_���3�1~���~���=�����A���W=�=QV|z�V����ο+P�ĞO�,{.\�W;G����.(���r���8E����O�GkK�����s���)ʝ��*Bz���s5�v���sĞ�g#��
G�Z�2z}]D[�%Z[��h�H��Ԥ���	�H4��J�`�/i�KVι�{bN�j3��8`8r�K��P���󥡺��Y8�I��GƸ%�P���X�iF]�B��Z��6+D���m2n�pe��6�>;D�@�
fm�r>D|"����Pc}�Md�.P""WK�Yh�J���5W��8�,�g��rV?�쉡�2p?"�3􂉭ԁ��"�� ��iK_��8�P&�%��'۬����� �?n]� �V[R/jPֽ[�@ң9^{�-@����cui���R��h0��M�
�$���P�j*����֒��P�����R�n��#��k߮M#F���!��M��� Ȑt�-N��l�	9���&���O���/���ד�4
f^��6�1����_��!��HpÒb
��O�)�|k�V�ĸ��[�,�ó࢞��گ\��8��$����l+`d�VF�&n�[L�M�lb��i�+v�c������+K򫨞mw%Z�ҝ�J���f�&�i�V����[e�X��LV5��+� �H����ii��k/���D��ߵ$�� T�`�:�x�ʴ05Z����b4�t�W�dFiNKk�M��p��x��0���?�ٔ�"3�	��emP@�D���=�5���5uTq�h��V%�D�Δ���b��#+���w�uW���л�0�6Y> �{�er�|t.��>�J�x�ڛ�k#������F�IE�Z`c�]0���1&v�U;�̧a��0K@�T�B�9�¼���h��3�[��1�