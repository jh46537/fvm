��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�×M��������`�X⯰�]<h��� U���o`7� �$'8��o��F�H���G������R��qd۶,L�X�u�����(���B��9 ;s��*�=��ߞ�A#�D�p��&�f�}�u��/�/��	��e��,��n��I�8YƱ��� ���t�
9G‹��Q����.9D|�+�3��q*����kL[�o�|y��//�}dL��O0�H�O1m�9�zo0�����A��D�!��BB��6�s��t<�"�/SN�	F��������
`��}{W3�á�c�?\l�����"Kz��L��|��=�Ӛ$O��g"$_�ƿ�
m<%9�	���Y�ja�H52�J��> ���M�Ќ��q�æТ�g@
U�" }�i�����у9|�h;p_C�$|"�v�zݮ�z����-+/�ڰ�����א�@���E$��.�<����_lA�d�X�Fa_evLh!�.����D��Z}^f���0=�Mr��2��Zw3�Y̿�_���٫�������ΔW���[H%W<pm��ZI�� ��yz�N�k����}u�CżZ��j�c}�"�湱F��X�S�Ǟ�Z����ת�Vi7�T�� �Wռ�H�:G�"�qs�Dz���忐3j�𓣼R�5X%��'�Op�qC	K,d�1���7PR[7�&�A�bA�{���z����&X���3$��$�6� ���r�ZQAz�3��t��J�ݍd���g[Ӆ1��9�3f��|�����)(������и[���/^�֟F�/^~&EsZ]�О�='"7�Jf	O���evc������Ŵ�9�%:*1�n[�!˿�Fll��|}�큷�I��[d|r!rBӿ���&�zH#�C]�=S>]���G\�F�H(�%���dzQ�[Q���#�|�_ئ��h�G���i�dȋ�*�˥%܃"ݿ��J��1��s�Sj����>�o�B7�d���'?��m�Y��z���	��R��>�τ]��'7�<�f�s���f�d�ɢ��br��/��\2�Kſ,����C���3	��.#"�M�^	PFgb�3�A���amQf�,�^ξ�;B���+!�뜇V�4t�y�E֕j�ݠ����2c�7x���.�g���uFt��\6�Fbr�WC<�a���1��8Y�(!���XظDR���JQ�6���=:�t%~�7�&��%��oh�L���	�CN;K�O�P7kN���e��G�
�[���Q?JV��D�Va&�!��'W:��I�Ș��Ȋ6�Ms��Tm�>*����,�ḑ����&���0O�+�#����.�S��3	:��3��~0���dC�mo�Ov�p�5Y��k�		�Y$��f������Ւ�O6�f������Y�`�����[D��>z_u@�ػ&[u�R�I�.u��ݖ?��KyCT.��鏄	djuD�����p�*#h��Ǚ:��ۑ�ԑ�źުI:�Q\�.��:k��)�Fe��;�O���`��2<�����1���� �=����"s����Թ�@��/ϭ��H�C.���"/�C��+D����iDS�zm��7Y��:�����<��!w�
�T0=V!��ӹ�-���ʒ3�2��[�C����TrZ��ɵ��ud����|�704bt����K���;��n�b��T���K�T��!�btM���3���xs/��)V�"䰢��)��2��ޏ��x��	ǿ��3��2϶�����@%�.��Or����>�;����|hʪh@ޒ{����O�+ՄS.,��<���˦�f��~TEL��\Z��x`��(઒) �M��jT�<����w^uQ�g�%/����ܣ�n����g��ŧg�TYKT�<�y2c� ��?8%�$�E��5�B3�c�Y S����s�Kf���[1��{���<��c[�o�����j@X3^$����O�㈁(����r�~�����=l�Gӭ�ˠ��YSI�JG#��Y�B`�ɒ�$/mx��''���?H�v_8���6����e<ģj�l�\"u�'�	-��忥Q���l�㕋���"_�%�����cۉ��H9t;Ar�8*��\QHB���j`z�l��X#F�v���KN��Z����<d�����,݄��]�&0y_���i|��#f~�95����O?yW0��t��;�b[��/>U�܆�Ay`l�\J,��1�KI$!����e״l��E�]�;��Т�s�|w�+A{�i��y8VY[��2_�pkɌ/�5�D�d���b��NV��Y�\JFϏ��B_�H˫�W7��>��H�s���tԛ9'/�g�OO�����ک�0LF@c�[�Ae��huv~{�.y@�����!�`��P5,IM _��q��`�i?s����V�xC�Ģ�k���Y׌m����)/n����	�����+���k��O��g�}"x拤�Ͻ�*�0lMZ��*ԍBs�B����(]���cT8�W{P��e��V�9H�(��$��o\����v����A���DR�ֶ;��c�"sI1&P�b�f��2v�ۨƿ�&��AK�b�D(`H�d,�Cq��u����Ko�h3"xT�1�9���}10<��`�$Onn����41e��<�9!��R�6*����a���hؒ�?��SZ)� c�����լC��V DƖ�ﴀ�����#�w����,,��٤4��X�M7\��Z(<S?FBV�� ���(u�1?3�����<���	�3/<ȧs^�K�x4������A���B9�_2�����sUb����h��7'	ӂ���PQY�m���׾Z��L��|Ў`�~a�|q�@��+9�@Mx��	��3������.��g�k�"rݮ����-hVO`�fL�l���3�K�v����������(����JF��<.$-.�;�D�{V���!�*�w��V"f���x���wB�/���q�%V��/��)�6���@d����Wi�/!�|�(�ϴl��.>[�6oVk��kFdDg��$�f Z!��wI����f��b$��84z��?dEӡ�\��2	��1��W��:�S�\��4Dh=xK�t[�p�#�H
�K��@|a���Q�J��r�ϻ=����EDz�̢�i�J� ل���O�����$��.$�C�o|��؁$�̀�E�]l�q���<_�Ԃ XVh�$� �/Y��TB6;�V_̯�����W X�z��ύ��-����<=����&qFJ�u���.pR�T���ߕ/	�ܓ���W�ș�2�|ی_�0
�
U�FC���]�eƖ�.b"=���לrsܘ2�%9wIXБq�d^�*|�c�Q��1;0��-x���ZG�//��7\���������0���/b�߮��ZҊR�YJk�A�?'z3�4��P�A?b>l(�?����Ũ��t<d���YB("qG2�E��!��S��`���w+9�f�:L���(�I����˄��&x�5_Ħ�'UP��|=L�(o�3$�hu��CIX5v�q_f+���̰�K+��u�ObZ��L��|�b�gA�l��č����?�[U1�Y����6*Pz�P�S�ݶ�@� ǝ4����z�7���t�R�W���z�P=��L-�p0�` ;��~� � ��)��|�D�7=�tD6�1��"ʸA�i<�&X��'�A�3��]f?z+�Tr�h^GNl�=nW_���ո=(����]�vvGZђ	ˇ׊��*A��P;ֵ�v���V*�&�_�⌶[2����i������mW �]Ņf�;t{��1��U�S��%:E����3j�7��GE�B{lAi����//����.'��c1P=�qn�W̃\���l4
��1͂������� [�7����DY8O��[=-��:Ѝ�eѲ��+�oB��,��夷����{����HM폱|0�cd� ��f�<�7'�@'�p�ϯQ����x���,��7�Kw��T�Z݀������:2y�J�-��t:sb{���s(��������ib�=Q2đp�'9��2>�R|��i����Ô�<0�`[���&��ztJ�C�`�����_��m[��@Hp���?>�	�9a�:W���$��|&�E�8(��]?��2�I\�)� �A�C�:�nA�i����7�>!�&�m�G׸`R�(�X�T��y4����x����.(��t\DG�E ^�V�5d����u��
fB/g"���U���BO�b�T!6V�j�ֲ��	e��ܭ��s6~e҃K���w�/x"h�����^�4u����uxȎH'�#��z���"8�X��9��=�$�Ƌ����ñG��{�2o-��Fliny��9�V�[s���ށ�s�A���V���{zCHu������E�d5!�Cdy��A@t�c�����Ik��$�*a�)����֒��ߣ8���k���R���i���޹��,̖=�D�"�/������yAn~���b�,T�V������a������e�<��f�(e�Ɍ,��èp�
Μc��_�Z}p�\jC�����A�H�����A���܎�?3F.^'�M��*�!i �l4|��[��Àl�H^���m�i�r�h{�^$D�g`��J��A���^kԲ�Up�R߫}���!��Cj���>��*�I�m�\�'gѥ2��.����X�=�����t(w�j�f��n����� ��k��l�(�js���bu���
Z�B��.��H������NJ������,öԐ4�v��o ߌۀò>�crS=T�9����8�!��
S��0O�h����贍��t��Ĩ�� uἢ9l�{��bJE����ֿ�?�#�L4H�!� ��g��6�_�[��.MI��ρ�}��1��˔����>�QX���(���>�#3S���2�
����(��Cܑ���v��8��"Z`ݙ��2ʭ�ow�[N̛��l��(�>gD�@\����[\�\�2�m���&�JG�<e�S<��1�YM�~q��ˈ�K��:G�,�:o�6���ڗ����,S�����KB>m���qq�=bL2q��k����e�z`�XϢ�Q��g$�Hݎ36�H��\���u���4�/g�$wxzR��q�ˑ�޵��$���hQ�*3{�����?s)T��\��\@��G�f6�,4S��� /�Gj��%�T@׶ � Va5W�]β�C���M@24���)�h���:��tښm�w��ce%G����l�w�\5���`Q7.xgCU~'xz�-*�◸&{�.;T���1;J���ʺ^ B6��e�ɉ�����cF�g�u�l1ܓ(N�U�����5�a04� ���+F�j��9x�ʭy����"/���C��ө˓�ȱ�. Q�7uy��q��ľe�ʏ�4��}/�şT�Zt�%����SD\j~�J�K��[d6�z� �����X[���ØbS|������&&��s�)�5����7���r���O���Һ�l��)w>��P̑�?�=IC��K�q��j�N�0��O5q���j�uҍ�+�����e�+�J&���T;�Q6�Q����\���D}�*	E#�'פY�}���"�г��ݏ�V���%�I���7�o�L
�8>������M�4F$:Dr��B�3��z2�,wk����������Y�^�f���(�0��[���n����4�ɁC�/nI��ⓛn3=�${�e��:��ȳL���>#B�����Yי�W?�NΏ�T%�>�U�:�V��y�M����NHY6��oe��*5�t+<]��t����K�?�P��<�9�;kˬb��4T'2J�����f�C����(��"�Ih:����ަU�m-1�@�Q5��wP�J�֝_<��f�q������ŌA�dq=^Nq��\��a��,>��gC���,v�W^��y6@���Q׶�bn�:;���89�f�����U��Q{��y��M�z�т���������*�a�+�7/b��������с�R��v5	�ڻ�k�@�S�I]U�7pu($�2�F���y�(���˦
�'}�ｰ1�aֶ�EY܌Q��&M����t��U���<�p&�$^��?��y��ؙ50�$��8���"֛�=�LQV�H�"���e���+������F�@uM�%���T���>
;ļ�m��
�Bn���Mc2�ﴵ���i�%;@	���ZU�B��>��DM��i~y�L&���"�/�>Z�{.��J�=;l<cK���HskZ�����~���,w2?�W�J�g��䘱�BA-�0����+�HP�O��2�Yb��� [�¨|"�5���2P���S2���;�C��89Zv �h�[���Q���O��s;Y�w�ͭ�A��4�*��(��f�3&C�6�<��3B�~�b��	�`�BKy�_�r�(�z���8Q��su7���S���rE�.�3)�S8��� �����<�Y%�;r:��9uK����lkq�|$B��c ��!i9NHS7N9��q�@�����3Y�I��[h���k�k7����c�C3�6,����!dAOxH V�����b{�>��K���g�ri��7�D�ڲ��������C¢�_;/��i�_֖Xqj!��=|;gy�[*Y��W���
m?m�v��W��	+8��
ـ!���sc��P�3G��J��I^I99,-�@	����tg䏏H�M�X�<՞y��)��ɀ�9�F���>�O��b*��jW;ƭ���eѼ\�cj�u��c�-Of�`���񱈷�i�d��Y�����S�uO����iV	(x�p7E�p����|�e�"ER�������i2js`�.��Q6O@�UVڣ<D?mr������̠F�9�.�X����-]���1�=ȍ��G!��J��Ɖ� (U�����t���D�IOۅ�c�e/�}��R�&"֊(K<�8v-}������aH�+�O��ۙ�GuO}R[�p���Z
��B�J$W�U������u&��-d����O�`�[�,��������i\&0v%e�ϼ�
	��`��=͕�)2��G��b�_5	�|��W0�J�mz&��3Z`젌������P`�v��%��C���4�����T�s�)r�+pմ�����+�Ur��Y0<��\k�μ��,��<���Dq�Sb���_F��Ͼ��p��Q��l#�I֬��&PH6��c@�>dv���h�<W�ѝ��b]����oܑ���/X�)��A�h�gf��CMUs[��np�-���KW�gw�z��	0��{�
���D�h�_�@�zxֻH* ��ʅ�^/{㋃�e�3܉�����W��w�	{�A���6h�Oj��uN�yÛ�S��������[�[�2�{�� �i�;�%�(pw+�+fO,N����;/ت4�W,_O��� ��\���D�U���G	�#��� |��O�:�^Q�\�W��*vB��w�h)9�秴{����p��֢+��0s��{7O��G��t�c�G_<���E�^d��H�|��?�ˮ��2w���x$�8� ��&���^U�����:�G�ޤ�LB�_�?X���0 !�BB|L[b��H+���..?��e�G�����A{�"V�8]f��)p�T:CN&5-Zœ�Ӷ���r�=����XO��Uu#E�tW)�>�?
�N�W`�2�$j����#�^%���RvO7�i.Jz^��N� ��)���/r�9A�
��ج R��2��F�֖i�@�!�/Y�wkB̉6{��@�oB.㗼Y���0�2�d�ͨӣ?�� 5�+�Q����
�l��7��������<��  Vl�qBE:��jJp��D�Ngw9�<w1�=�#���1:�2S��� ԅ=@.}�w�Q���B�άؕ�x�6�f�)�����F�6��P3\bz��j�9���(��Y��YA�y	�T�A����G�����>z��Qlg^�2�Q���	X3�1�!0���T���X�ʌ�Z�.�}X�B߂��e0���	QLtRru1�,�&��P���O끫t�N��/4�'�.�ω�5�����29�tO�#.��P���j���W3SR�y��*.��'�^�{'��^Em��d�t�����x^�E��/T�T�ۀ�f�$��AWiWݹ�؈VW�Z|�x+M�{�L�J����mk���-�jl��>6�y+��;��v�E%��>��W���~��)A0�Ct6�ה�&���!,��Nq�;�z`�c82ƕ�-L��	6$��&P�F/���t��֨tUې��[�����c=%�y{�R�Vh��?�}߰;�u(-�� C{�25�H?z��2l0���t7�J=(a��B;nBC�	��J��+�}��*f��n�Q���'Na���NC'J��,}i�QB|?��Bfk��p�c+äY�s�~Z��{]��`�o���E�|>�} H��F�D�G��F�Ь����Z�^��4�^WE��>�Ίe�a���u��ԡ�9Km�~��7�q�{	h;ŝl��n"Jw�G^է,�,�����V�L�p����1-<�C��ߓ��J���\��M>{��Ҡ�L]�M�Iu���'U2+���-&������%���Q,�iD5��_u9t���@1��7��r8��TNl5�g6HXh��m���R��f�##�x�t7�hb's�S ��1
��$g'\ ��J�a�uɌӂ:�Y�m��T�f��#���S.%��'$��aDa����0�,�q�寛1�Eg�H�3�2&鱗�Oe7j���Z�[=4����18��8m�~?2�[��0� �N�e�rLT�/�z5�Ȉ}�խo�:���NYI� �:����:�wc�[үi*=~~�#ɂi���2�%�X�^�q�D)�������QLZy5�k ����3y\p�/?qI�-��1�KhҕC-�FD{Ql؇#�W�v�]��Tio�#1aߚ�yg27p�?
NZ� ����������	�D�UӦ�E�	~q�ABZ�u�N�P?�P��K�,w�?�׫�2K��Wt׺�U����������zL4��)#����"�L掩P�?���+��	K����[eB+\�l:���D���I�DɓfV��=k���g��X����!��^b�(� C�w�ݑL3���1�t��A��c*�����@\�� ����p��5��Q�i����
?8Ǭ��k8�!�qy���(���ĒF(�ʮ)�����*�������ъ9�ƹ�G�J ����(|$&�v��"�	镟b�^2&�tdED}�����O���XK�_8m���]�ooфW4�Q�g���h����]v�B|&�SҎ�ˌ�ܮ���XA�Ή��c`h����^=��.��ҪW��=w
��=fN�M��Ttt&�4H�W�Y��.m��ÓSϠ\�~;\$�E�2��Z��s`90�31��m2t �4�Z�<�I,MŘY$]=Ӥ�H�A���p���}�N���*} @Z;X���E$mt��2~��PwJ�2�1�q�EC�ak>���a��Q-�vM���%��aT�[�Tگs�n���6.ޚ��.�yH�M�EI
�JV���M�� Ml�њL$���Sr�"�l�@�<��U���=�aR���Č悉OBk��.\ޚڬ9r��M�E�Z��y2�N���KF�3��U��Xö�>�E^M��z"��̹b��P�p� nqg;)�����Q�\�#��0k�f��� (Ű��ܖb�(�(�&Y�P�~9��=���7��~ 2Vh��p�})�Gν)v�e9U�m���a����&f�mJ��<v��������l.Zwr,�0�,c�֢Z��1�������ط�t� �TY�W�-J��~��@C���N3�`��/���w��K�^���̬��};<ˠ>��w7�dmR6@ǅs��t'�͑ ��
���G[9�;��%}����f�.����6�)�p�H�:w"2���Nָ��B�x
#��q�u�k�)��iͷonl��B��	����m��1��8�Ry�L��o�{qI|9���,�Qzhvm��s�~�Ck��K6i��hl}$�8t{�r��ou�,M�{՜��a�ZC'�aq-�ҨNf��U
{�֜�����%g���4�m_fث�_m���K�SW�-l�$7�:�����x/4���,4:�kb�
P�i���Q�d�#>�{Ju(��*j�|w�U��c�pd������p�Np�'(��ɭƹ� yJj#ö}]x]��r톙�ָ�JHu�XG&�c>p���'�,E�޳fEh��`'P��P���Ic��i����ԒS��cw�J��$��j�ZO.�2�/i��I�MDԨ�#��8���Y]�X�7ʈ|��u*�L�� ;��#Y�����V<X$�����VY���aN�"JѷE/7>���Y�/�ӫo)�{�X�������e�����O�S�	�2PBf� �����P�Ds���O�CA赫�<t}F{vV�?z�p�ϒq��,Y��%ChWȰ����P���f�(���!%���+��B�`CZ_���֚L�y<-����V�$���Kpa�m�Sf��v_$[j�Z�3���	���o�&��Єϙ��r �pw���h�'*؜���:�����7"���m��,���o�<u�7W��d�A��˥��8�1�J�l��v���Ϭ������P2m��G�v�-��m���?zg�ZFvJ�g�d��@���5dƞ��3�D2PB��e$�FhPp\�}��K{�!�;r�B�"����M��+���w��|oI���6#�^��CR�<Yz8S�^����ٖ�Z?h�_����*p2���L!��Kw�?G��q�1�8��8S8��)7Z�
�t����=zQz:,�˩d�>�[�	1���X����W�����2d��(�Lh<J�x%�tg����cf�u��䠋.��@pX�'��]:u���qkL�(ր��Eq9�=p��U-�5�t��H0?�]�������G���|�!���1?�����$�?T}�m��Ѫ�D�i��{b(iP����sR�a��>�v$���g��~���ޮG5{��w���j|24b��_���lr��噶���O!vU=������v�ۘ*��;8�s�_&|+�,������F9����8���'����-��"uKB�7�����oH�[-�����Z/�=�K�xPJ$����
o�ڿ�z��Q�(�[��(�m�o��$v��f�1��:6�`
��6�tس|���#uɠ;l)��o�[W�=v9��L%�MaRK��ڏ2�� >ks���q�^W�����W�)� �m��!d`��S���E#�I�M��fi��ϧ��W�����xVX�ہ]�2�>��P�ͅ���=�/�����h2��kO���c
��M��.��ֻ/����%��@�A@%���o���`a���6"��)���=zC�hdb�
7+h�c��ݸ-E!�\1�\��֞	���d�M��� aF�9�ơ
*���b�&J���2�:�aK�s�h��L�򊨌
�'�rb�T
����5��>�m�1��y�f��7p�i� m��2���/�`	2T� ��T��'i���A@|�p��y�j�$�d�@����=�`/���U�Y��dC�3ߚ)����? �:v[*�Oh�x���\���+�kZ)P�x�����^tBh��W������3J����v\-T�q��M/<$ �spv��峣_[e_CB@�Z�h�7�2�mI�@w�ŗ�x�:��v�"�'���8���x�c��k�Ϸ%4ˎ~�q�BsN�����qb�2�� R��Z�R�ʁ���W����BiG