��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm����질�95J{۠���D<_��`�vM���yI��eϝ�9�b�(Eĥ�����6��0��Grh��<�h���'&wOû!�>�k�N@'��".LJ�Ҍ�J�,;�K<��X����6�.B� ̒�|�&�P �#E��zk����e�m��}��4°�Yۼ�7�X	x�::��]�$��(8�e��-�V�ܝ]R�2������Ca�e���*l��v̈́AtO�;��;�#Qp�h0�v�)�l������
/��o�m���KM���.���B� >�-k�S
(��%1ve���LNP�I�AU��&!���Y��C�� y���^9Z;|�V�m�D�.�jU��*	?AK�kwA��<S��5)?x�l'h\���5���]iVR�KF�?��P��(d�����l�ܹ-q�Bf�!/\*`<��@(5�8���"�M�Ic\@^T����:��λKuஎܹe��z�����5��]�޴ &]�_�_>Ie^d�����
&G�.^�0Ӷ��Z��g*,����F�T:�+�9�G�skEI{�������v�{y���7h���ɧM#�U{s�agF��L�i!�
�ҽ��ن� :5�ݫ,���V��r\{IV�5$`_�19t2<ګύ�L�����3�v9��SS:%�`�긽W�f�:�ٝT�8e�8 �K�nh@m*�LV�hs4:�6;	gaVg͞���.�]��I�,���~�����%��@:�)��h��E�<MƅB7�����0q�O �����p�kZХKd<>����~颲)�_ޯ�YC��h{I���-�  �	�L�oa�Am`����lYc]S���s���'kX�������#���z�RJ�����uՄμ��&�/��t���>NKw���}��g��=&yޢ�<�J�'g�I5��1h�u/�@�;��7;��<���yB���+��Uѩ|�<�\|=_�}���<qS'�-�-xA��Mz�$�N6�}��u�����0C�m'�g�s��Ճ&紞�y��L���.KGٝ6\Ɓ�?w
zT%��?�3"�T��XG|� z7�7��O��ꋃ2;���)�E�;ҋ�[
��J�w�����?��i$�0=~���ڭ΃����⿭9PSdm�_/fZ{�PRVCs܄����Í<��\S)��PK�)��2d?����/� ���U�K���s�l!�!g�d��2�y���}[�.VmnG�E�`�V�P6f�1R�E��	=����r�PES��FZ2����[��^
8��c
�8Q��'H���̿�7RQ\�jJ�|s=i�EC`��So��pg/�n����Ni�����qW��h-�2b��.���p+F6�B���ܠ͌8{N.-��q�T	v\�RrK���ڇJ����?k���3`�40FC���
|/"HB��b��Wм�O��H�{ p�x�n���V��޲-<�?�&�g7��(B:É�6��H�4���ݜ��=C���y���,@�{z6�������Ǣ�
rq�d6VT�ݪ�$K�w���F���e�s�Ə���w�Z�x�{'��i{>F�n�t�#�x�5\�`�e2o�HJ!_5v'PRj5fi���x�?�;Z����D��a�J��;��;��1h����oA����6���Ӿ
~�ک,��̵؃Yu���=(��4M6��^!nՐ������x��<�;�&5����(��m\����a��$v3s��"6VW�3�Z���Xq��&	=�Ǭh�J�y�\s�3g����r�)������a.r���>��M�UzG���"�S�^ �X�r_��!X���`��:�q��_f�:�}�p�i���2t1{u���/�7!2�W�	�#�SD�.������Q�_���d5Z�3�+�甕>�h�;�_�~9�������99�Z��I�u$fA_=�����" �4��T/h\��YR�i����}dk-q0�atK�XBM��3��O�S�|;��#�fC�����O����B��3xt�i��2,x����L���8X&�bK[>���T��*JVʮ�R@���
I�%������c� ���IG�"�q��9�r��@s:.��]ޒ��5�>�bNv�i	�僣~��QvF��X�9���Y�^�9l8�rk?1q���2��c|dH��H�\���Ϡj`�~Tar"-7YC�=��Ia��[r��)�:<��0��=;׾�[>�::��/&�M���{�~H�����;�h�E���,������.W�d���˄{�[�k3,�Y!��h���Y(���G��.�f4*c��[���{�B�y���I�@�n�k��m��3*��c2�:��]}TF�}�\�k�ڃ�����H��PZa��P��b��־l�z�\`]�����?|���Pg7�3a�XܛY��һ��P��@��XoW�AC Ë�y� /��h��$�����܊�MW�u� w-p�`+�r���KJ>�pyD�'IA>����1�`���i��&nIq���b��vRv�K�gZɞB���A݈�����w[�E '�	uKy),3���ͯ���.x�)����u ��P�;U+���g�Z�w~�lrw5(j�2F���Ū������`�N��׼�$��e�J	|�Z�\��`�c
�{#���p��لV�*,K�U�����O�j`�(�ٝ�[8�v-�Z9/���e����4B�ͨ��Co�W�+j��H!m���Ɲ�����8��c"�K����f�X�o�A����7�&�x�+�Me;.��Vl�;�0���8�@ �ʐ��8I�6]}Ƈ���i��3��A��x��3�l�w�p��,ə�9H�CƌHf�?�k?-`�������l噧:����;,7��!!�2��ga]f��`?��K����`GfAݞ���P=O�t��f�o�܉�HPj��(�9�U���`��%�4���;^v�qՉ0X0�>I����e�S�JS@�kQܲ�lB�G�������珢i̋���%��RV���5�9��P�4W�7��tR2���xOPB��r��F�����E�t2�6��Z�P#���"=�\�pLT�:�D��o��Xr�L�҇k��IۖR�W�QUd.���-鶡ǞQ
�G�E��*S�����z����KUC�͸��/��cGxƣd��{-����C�����q�:=����x�V���T�'Q$z��b�@} =/��R�65y�}�k���M�겂�_je��Sl����~�2[�$����˔T�(XW;�69�����쒀V���#�׳�غ�:�ܵ����@��?3��'򧠟[^��#����b�d��y�_R�B�j����r�\��u-�zyq0
��a���h}�*.����/�>X��w\.Kg�i����nEw?J�Һ@���4�4gm2`��o�l�l�% =���}�iK�
Fw�S21mRV�Z�t���ԃ��|��<�:� N��#��fO�Yb��b�s�w�i�%��za���Inn#�Mc�)b
u���� �TEL�ØL���a3�	۱����W1��ܺ�g�l��Jw+��cQ���KEG0@ߵ#��#�=�*�ઉ����|�c#!W�0z��� \#\��r�὎)�qjU�r�>(�2Vp
S��'�.]��&�,7�����A8�TyB���D�<�TT��)�pJ�-wӻh�d���3�ZH8�����Fٕ���x[��mET�~g���[MΗ��(����{%|��N�!/����ޝ2���a��j[�+H��/^G[�d;v�B���+\���d(F��	�w��!̧�P`w;�9��V��(�T���CV����'����S	C�
�}˃���z�JhU���Oq�q�%D��Jy�=t��%ZLa��łVS�d���'7����9ޞP�<��C����\��W<��z��u���z�]��&��~�����0c/�B�A���=22$!��!�c�caHh�ɂwU���'�J�}���<Vꭉ|qL���	����:/�{���D<�s�K��n`�H-p�h'o��o�0r�xs��B�����u
$����=��Cuz�,�2�=���/$���=�U/v�.�P�}W��è��G
[��E#�_E��g��}
=��n��x��jtQ�d_�"�z(~ws´����ؚ]�ʖ���3��pI�D`�F��4U	!�����T��6)o^������[=�]_��ݢо�8�Ya8��EE#l5�1j���ŀ���g�M�p����������h�X������02�5�R �.S�Pey��>~���p���%{��~ ��S������me����[�0�_^��ʷ�![���#4o.���#�&򆛞<��� g/)���ٻ�BV��EB5�{�:�δ@W��^UF��JΒ��>}o�n��g�����Z�Ӝ���:3��fvP	l�g��ˆ����9�^��E�oLݰ��2�5�����M�_ۅ]P�4P�W�T3�n@�f�^�&ʟc�28���4�,��&ÿ*��#n�QS���$�6�ݸ4������`}��)��{j�+�M@f_?�5��?Z�~�$)�P[L��қ�t�r����%��"�dF\qI{���,��K,)�������=(��aL�:Fa��Iq�&R Ϥp���ѱW�r˩]�ج������<-����J�޼:�2��!yb��K&���G ټ"ew�bt�]�Ыj<�f#27_�Ib%Fq��3l�1c!;`@�sяj�l����-��zWf4���7{ԬГ�J����I+��k�N�I!	�]lMs}BI��R�Y���p)� c�Y �K�I�r�w]����:8tܔ���F�,#f;!%^�##q=��H<��~�[���'.�8ut6�P����b5�d�F1�^���[/KÎ�C��B����[F��_ͨ�\�<����A>v0t�Y׸s�
`�ѝC��@BK��#������8_�^�������`�bŒ#E��٘Z*��lx#�ȑ=�S���<)�}b�;	�\�ɔ�B�~���ƙ(_�Uh�G��߾~�T�b��7�,Ƙ�^��W���v���"nPRÓ�K�d~tl���J��h�uH��6+������*���زJo�+��:mY
��0��P�������A%'�$0�6G�1A�J�T���;�"��{��t�K$,@�k*�ڏ/iLZ�\^)�}���H���gO��n����[�ƀ���"\ ��h� �ϸ��	�v�a]�)��:u�K�����t��(!���0iA\��2o��l���	M���B�ˮ���P��fQ@/���Y3�B�CVI�n.(�9^�v+��mcZz��h�����!t�G�n~�!����:��4����0/�j,M�����!�n�2}},iA.Xq��1Xs7AH��*c���X���M��u��T��rE�}fHj���d�ʘ4Q�x!�<�{�p|��������"���_�1<"@&�����AO���)�c���Nڐ�د
�ۖ��L�I��*�{�{��/�y��s����v�LS��3�"��p=P�(�n�����w����?�ֱ���As��\K
~�Pj�G��q�9�l�Wb)��#o<�%�<��9����$@/@��6��M� ���M8=�Y�^D��r�I`vF�.���wv�4 �3еLg��+s�b��Q�z8��P��y<g�U5�7����R��J7u�v�,�=)���x���?���5��F���3|�l+�5ȺK�U����kz�
���aD�C�����o����� L|z��v��ߐ^����9�&������u5���`'G�n�&��7�6�xQ�Z{��\��.��}�T	��q7l7��h�I?�ͬ�$���h�;]��CQ�����D�=�,)�3����Ǘ�N[�ר���f����7zW%V�ebn^��5��7� x;���KQ�ϩ	���/J#�/'5"��tQ��ߴy��R�\�i�E���H����yǢ�xk8ej�KSq�m�����T� �K,�]0Z�A��X�+��-�#=��� �Y�c�D�R�$�a0��K"vuδDo�����g�z�U,L�	\�{��xO(�K�A�ZQ�~u_�&��L6�:�/c�����iJ4��'�މ|�F>K����&QР)4����t�٪���:t8���`��V�ޚ}���*E�]�H��-�����w�����X�Z�8���a��N�v%�֝;G�<�'��C�>>��G2��̶��y �R.��0�e������f�[����P�z���G7��>�0�y��A��c�*�1�_ɼ��HA/���.Iu��f��\���UX9��v��z��<�ʈ�)I��,���)�ӀP	�5U+o:*!�2����(m�4{�i�2οؒb�#]��ɂ\�.�J� �C�迈��F�'��0Ե{�s�&��|77{��7(��g���JQ^*�]Z o��/��)���S҂ScӺ�8�l�\��HM�t��a�""i"Z��p�%��4`V�B�6f.��E9�֕Z��2Z	�@0���a�Sc����x	�
�L�أ�5����74�e���a��}),n�l��e�WS�#Qs�b]r�*�9d{=ܬ�ѱЬLK��l<����u��|J�]]a���Q)�eU�7��Ƽ ���A��_��v0 _�8bq��lF*�6K�(-4�+����|���Atz^4a�W7-���λv��{4W�TW!pԾ��=6������v�Ԙ�g��2�M��eY}�^��}��6�{d�a�fhӬ��MJE�1^ⱺ|�KIc�J������Je5��/<2)�[�V�����O�PVt�����?�Þ���v� 8N���=����ؽ��94���ܦ#T��.�8��P���߶}�d�9W�������2,�D
e7�X)s �ו9'�&ı/
���}�w��VSU�46��ᮧ�~S�E9�=0~cvD�;4�S�9��m|��L0R�����!�z��w?�SW����N�A�6ް����]ɭ=�e޷�߁���l���r����<�G��-�ͳ�-�7���3��c���P6��KH�A)��KjQ�'1�:��P���ӥ��z�Kt�
˅[��4���d�����"��=8y�.NWup�l�'�������g*
��t�	ȿ�42����n[5�z��N�t[#�	G��5 �֫E4{����f��5�(.8;��u���h���'�((�K�'zq�zw�g�X�y�d�DgzU��u4"���^0P�[0��F��OEәY:���#���ȐH�<���rrVUuǾx�<�Z�0�#w�c���*^C�iH-��t�/�Q7~�0$˙a��/�t[&3�����0��8Q�1�2r)��M�.:'��:�U�f��ޙ�4�K��A����TZ&�Eb����E�	d3E����6��u/~��`p�p����#��4�t�Tm��t�l���6b �=�z��}���A�Z�V�9�D�eV��@r�Q�W5�D4�
�}�����q�N�M-��r2Dw�����6]*����Ov .��P�b��?�b*מ뿷?�f���οc��aX_��@�-���f��>.A���M��ĵH��<�oU����64���Gz�tO�0J���g����mQ ��;ԍs�.m���w~#A��n���V��*)XI��7����k�&f��x���l�g	��v�vzƴ�� I���W>ʗ�<B�t��ι�>