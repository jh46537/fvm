��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�
�
QT<W)|Z@�l@Rꦯ;A�C� ��.��W�m�"_��ͮk�N�]y	n]�N/-]��%F֠�n�Wt��{C��Z^���UtV��*��k�������!�kBM��\���w_0� ��;E��0yЭ���Z�Z�<k�n�iۂ��3��.!�=��l�j�'�>���情�z��w�"�)�*��}%�$\�#����
N$'+R0�����-�ĂJr�rZ�*Y'C)/F��"��Ɍ�o�\��xү��ޥ��k��e���$����?���_z�⋷�r^��n��e���4)�7��O%�?�ՐS|�~��o�;��:�!�}�i���.{;w����/p�?DVd3��ؗg_���h�%ؔ5���=B��_�|���w� O�3q�r��I:�b��p(�Dc�t.����9�/�]�*�)g	4x'�ۻ	N?qI��*�nY���;J6����݉<R���/#ݜ@��_3��7jr΢�!~�@s`\6�rGEQ���ý������y{�B���V�6� W��;VK�2􇵰�'�	��-4m���x	E���i�̲͔M&w�D���,L�t?�҆�6`�dBi�j����XV�qc�u9lũ���9�H��x~$'�W�I��L�̉�/���;�7�ݡ�:խ��D� ��{��scS`�"K���&<@)}rc�_̜��x>B J0���=��:a�@Cl����&�z�Ug�/´�V+p��W���l"�]�>�;
K%	�]o�n8�b��}�E��*�� UEQ�}gv(�A��7in����� ��W�%u�y[d7b%���ޡDM}�����!g&�������Q��>Yj�y�p��l�b�x�7*y' g��#��c)�� �Hf�=J�~�fU��5�_NMuC>�ͼ����w'r°�,pe�ƥ�Dd/+t�-1����0��Ά���[cPɷ�1�HX<i}w�X^
�4��"��G�Z(�Up��K@��O*G�s�
�F/x�V�Ct��u}y�Է�A�OE��N�dK^m��D�m.j�����}��\`YP��g��Is9�wy`SaD29�h�9dϩz���D�eCiI��le�0��C����w�ז��Ȳ�0c�h����o��%��sbpK`lS�*� �v���sXܼ8��l|�,�"��NN��qHʜZ��i�Vl_ê�^y��O���}Z�������Ou�����%��c��	�}0���֩�N��7B��W�R���kl#�!�weC�Z�Zò�&�?o�P�>U����y�Uxt*�!�����j�൝%(C�no�5�ho���BU�/gg�9t1[������i�7�O���x̃�|ܒ���Dұ:LJ�35���!��Y���a��0�]%f A8�?�g�Q4�S/��)�B��"(9������W����Q�V`��.��*B�ߖ ����2PL���Q�@��'�:(�%C��e�&��9{����W��g3�]@��j��b��M����Z���VX5Z��t�d���|�;t�-�ʖ3��Z6 Q^3��!�c��r������
�F@���[�5����A{7�;D��m�@n�AO�9H�I5�9R����\<l&R?�c^ȭ�հY����{�7�ǒũ��z�x�ޣx)2���*���Ժ��ꌉ}�Ӫ�c�wl�-�������?��O8r���I�b��.��.�����p���|0J�����"�0���}���pW�{��E��������؆m�?��j�3)n�>[�]÷c�_[���	��2��e��Q�
���K���!�?��nF�alE� p�[���h���o��k��]l�m�����p6�JB���"�_B��f޵S�_n�����?*P�»T�̞�8���}�v��t��6��'.�$]����ڢ����?,@�Û@k���Y�(-� ��L�T�v�oQ0uf��@�A.d��{�������o��i�V���N�|/d<�!����N�C�+ƃL��E�޺!����{\㩟8"w.w ��5�)���^��m��)���dU�:bS��]�|?�'�ٛJ�C�ovnS#�֗h C���tx����&�[�;�W�oz	��3�(�ʥ`cw(�#{x�c�c�x�m %R\�zT�`�ܷ`/)�/�(� |eR<��j�ť�{T�4�I\�b��^oYO�d��w�S�Q�I��9K��O5��o����,��oF{uQ�p�w�b��|>�F�4I?��FGۿ����uS����O���*G�<�`�=��|��P�6����6h]�<`y@�_�dMV��bw������IYa��g�
�Ц�!�@�$�8`��ĸ�l�LY��&U���L��M�M?
ťmQdND�4^��DqR^��j�.8X�v�h�F�V<=�����"�\kF|E�1��x](�����6 �*J���|m	��.�M���垩?C`�N��8խ�j�1��w�|+ >꩙Y�ބH�y���8�D$+B��j�+FwM�c�k�ȯ��s�Hy�}���ْ/�r��}/�7�`4�<)��ri F[�и�7~���Y�����~m�)Q��I-�ǎ�Ν4#��s�+m�չ��QB����{m�`��_Ԗ���-���]�37"쿨����|�鞠%�Ξ�PG�M�C�l�)���1���e:�/���y�/���+ i�eg1�x��g���Uc6Z��v tu����L*ibhu�!��:ؤ�_DK���	k}e��ݥ����kf����ч�ltĴm�p6�F5�{�	m�R�3��R�5�V	����]��lDd���{@�R��*�3�����9}V���/aD�~���a�G����� ͦ}����R�P�Qsz��]��?��B���ZC�X�R�ܣ�	N�$A��9f��:�`TPBb�KevG�Gנ�B�/�:pГD����!:��KQ��h���Y��&�������,CYZ:ˣ�gt�"~)�Az���%1��~g)��K~�Ka8�oR����+1�y�W(Y	Dl�+�G���^��|+g�1�#�	nzԉ�m)t'x�Q*�PM�͒Hh�@lX$�p��+}Bs7�6
�zόы��꾔��}?:�u�BK�����!m m�f���(�n�`���u��f�b�|/��[cs.;�[͂��ؗf	=���`(�Y��A�+CZ��bO9���Iʟ��CQ��]@uV>~t��g��)��]�0�W�Ͽ%+���,Vch���t�.s.@�ԃ'dwe�\oN�PF��1�{m��\6�m�q����k�$�e2�Q�O\��a p֎��$9�����QD�F��.�Hf��S�9�8��[uy�S�{74����UDϵ�R���-9[D�f'�;g~��?��
��Q��$�>��Λq�`#��d��S�.���-�8�_ʷRo{�:���(���8DH�l��)!����2g.���d.d�hʦ�-iF�c����aS�>��v���d-�|K{�tD��C� ����'&o��u�������N�;��	���Dw�,�q�A?{R}�{gzM<6�s��)�FY`�� ��gu��Vxю�EҵT��Uo|:��)��=c��F9����_��+�J���WQ"b)֝�0�r��i@�V���WÇ>w�U�7��b��]蟌�HHj��&�:�1z���y��-��e���L�,b=g��q�P㢋c[�D���|�8�X�tG_o�t3&���/Ѷ���{��y��*;�̶��䍋*R�<Þ��d��yO��Ap����H�Q�*�/����s��xgRu#)���c}b^9��;�G����v4���\3�ϖ����a׫f��:���&L~k]����V`�<d�z�wK��N�p3�a?�ߘ4�/�H:�҇~� �s
�f�mA�3''��cʪMkvη0��@���[�0�A%j�"�ʒ�\�X��	��T�S7-H.R�?sF�S�7(��m��Wsd�wǹ
#��F����d=B�[�=��,h���[����b���t�݅q�p��6#�r��6��%���Z�|~��L���f��5�h�f�L���	��[+��z/br�)���s�~<��ȏ�^5�v�� t���ZxC�V?q�����3���"2��Z6�K����c6��4�퐈��G�ș�,Q�� ���V�����Ƣ������z�Y�"����H��ZJ�%���w�,���\�;�y|�
���sAS�5�1�y �8��	���#��#*K]��rza�3�|g�l�I�1�~%yfO�Z��6 �3v�Z��^��Җs>���I�T?�e�����d����æ>���?ӱ��2�r卼&cMn*N=��u�H>���Q���)k��T��������ǥ��L��J|�񟾱,�ܜ�O�V�.��Y4Tʊ�[/!���w|�#4�Ϊ'��p��
�k� M�|�x�,�v����f��%��$���-�������������R��M�k��B�(w2x��鏣+W/\@�R��P��βUAШ���g���1I�dmύM��Du�nC��OI#h��ԩ�H�oI�w.J���e���V�4-��Bd�&uP��U1���m"�����.4F-���Z�ͪ!��KZ��� (���#Y$7���`3a�v�W5X��8^�vD��#��vC�bT�m��c}c�/g�O�W3��G*XӼӁh+��]�e��DR>@�s����d�x�|�W-��M�!#)w�J��-d
JtG�\�&ڿs�Q&�MUp���*^�c�u=�S�1*�cgv���M�kСgT�VmR=���<o!�oX[C�z�5��=�8�	�J��f��Q��v9�ct��ӌw��7�]�(@�c��I(�m5�>X@�`���L�6�'3:qų�9�������)A��I���Wt����(*
�0d~�G9���As�N^���%��Q��l�Z������b#H��N�m3��?�
蟞_�X�e���ź���.ݻR�cU4��	-�k )�8�z��RTv�V�$�@֧=�޻��䀈�`[-��p��K��U�����%ש�i�rf���=qV�ӌ���9�5���eV��ԧ��Xp1�~���˩�D��$$M�R��  ���0�0:��A��dn{�o��ν�Th�kE���>�	���nB��z�'��n��R�穘����[��36L`��\���r�'%+�#�Ӗ�4P�e)"��Y� ��'l���[�.���-���ϫ�,����<�K��t��K�aֻx8Um5a�O��/`���?������hSU���w��Y�P�τs(��4"
���0oF��r &3��X&0�
F0��,9���S�l������p�c����e�����0Q��f� z*�6 ޫ�i
P�Ag��^���у���׏o��L�#�b��w��*��V;pz!t�cn�E�a��U)��R='�����[�N�����#$����#bI�w}����Qy
�
	X�U����,VZ���q��'��w'@��Ga�9��χ~g�����=u�X+��Uy}h�Y��U܁'ɳ�/AO�`�1�
u�팣\³:8~�~�fh�R@R�0�k���J��V1<țlF��q2�J�~,Z-)�2�U��C���ßgԳX,�9<����2�}��] ��оx�s<�!ך��֑�����QoF��޲A�%�� k���k\�vo�o>�[	0g�F�n����wd�ͽ~R��Z׭ �?r;������'��i0P>��
�i�ep�ۂ����ȑa�AZ��*�5z��gd��8�2�Q�B������T�tr:��Y#񛨭e�,f�M�˻�G�"����m������9����W�q�!��Y
�Z��/Y�Xv�@�H�����.g	Qg�4(:�=�s��H���k|�(r��a�xFt[{�dOj�E�1<�����/w�+�����B"�$E�AnhHk;y*1w���]b�_�	d��J��_Yr2\-O��@i��4z�N���`qթ��y��FT�W�*�5����EQ�B���>���H����y����/K����(%�(9�xђ�؁��<O8	���B]wֵ�8\]���ВP�%&���?�� R�a�a������6����]���X����g�ire�p{�ũ�8�ë&�`^�~ -����Y���W �8���?�4����[���P�CX��>Z�8m�b'�Y'��4KD	�ty"�Jz�/v�"72��h%�*/eݍ��FV�-k�]kP>��/h����/�fGr��߷0m�����=/���+	k�>/no4%�	B�ϡ��	�d�H7	g�a��,��bV�7���Ul�*����D��(e9s�Z�]@�	�e~(�� �Xgl�))m�Hf	��b�ט�*D-.ȻV��_ܲ��${��j�@��� ���eU͗}��
��t^��"�Pr_k����u�����k��R���W�u%,�ܴ?���"D���c7�Zq�2q�4(�bB\_b��L�j%�{'h�T��9��J����O�����]'��:��T[��>j�z�o��r�JR����/"��K��Ŏ��;s+Ff�@7C�[+�9v�s��W�x6��#�dp��y`���枿̫��=#����.����U6RÇ��@/9m&�d��W�K?���[e�Ip�M��x�:
�G���2��)����ڌ_S�Z����;G;X����<ڏ��.��R�LRAa\�At�8�|O(]��蒷d���o�fo��O��[��/��'U��3:��O<Kt��O�JB[7�8�9"�\\���B��_�|o�M�E�c ��B44���@�畫��&�r�����Sϐ85��o����ǥ`�򃱵�9$����g>��ތ4=uνQ��_li�Q�� w���pI�@�~0�/1��(B8R��ڮ�^�tI���z�S゜}���j���'ks[��?�"A�|s�K���'�ނ /B��<�y/�[��m  Z���B��(B���<�;ki�;��Q��E��ǫ�0� �7MZf 
~<��`���D\e���!Ǳ�d*c��9��9����e��gy`u	���J�����3. �/��_+�y)�Hm-R~���o��zm�d��� c�b{�d�rZ������!|�fz�D�k��c�#B�iADN��r���cq�H	� v^8C$�����}.�#&e���lڠ:@LU˒%��X�%s�"��K���^��.A�S0Ss��������I��v���;�l[��ٕ��h�^��{UAi�͆rMւ�k�Zκ�v��ۛv�������xj|��<<��*��7ʄ�X�v�۳�;�������ӧ%u(D�/2���t�0X�Rݲ���_������&�HNb�T$�w!��~�m���~X��+����e�.�E�=���}��5�`�*\�I��di�g���p�Z�s�5z�j��X�����{�'�S�7J��&�� ��[R�("�+�e���.]����r���`%��_��IHg�54Z�p��K|��b��iDc��u�%P���_��-|�B���@�6ܘ�U�d��qTy�)����K%�����n�q�A���+�}��ڍj�����-��)�eA�9g�0䇛�.֍��[�ְLb���fe=��&�Rrh�u�q�hV*�HXu>����5]���Cɡ�Vђ��B�] ur慽<������0M���ֽ���9Z�Brh\���x��q��NW <Y��M�%\X�v��qEk�dH�S�f���|�뉖�O��T�B�x��^��Ve|��X_�;S����;�lML��`Q;5fZ��ɩ��^�?�9��Y ٵ���=�eL�Br�ږ�����A���I��I���'���!7� ���0�)�f� 0�c?��Ý�fF��� ��A��o�Qp��~L¶}v����(Ǹ���J�����C�5�U�+�9��\8�l&�%�ʉ��נ����I-�y�G��n>����'+ ��R:���6�\�����L�sɲDZ_��C��V��P����ڡ=����f��b@Uv���)wB_���o\f4��/׾����<��Ig:��A��(��s����%�����?+��,�;0_�P7�&�#�Ђ��X��|�+�,�vj�d�C�xd�}�Аa�%�Y�^2OТҋ�:C� 9u�3b�<�,*����:W����W�4���1�e�oO^�ye�=:l���)��'gE.��8m��U��l�ap&TZB[�q��_F��}�d3��Vfcg�op���6�dr�~��0[����v�_5\�S#`��:�P�~%�mh�#�Y�A24�BN�N�>VJ6�ۦ��%����	�2�P;y��1{���8ٿ����ie<?��a���MU���!�MLw\�-�p������]�� �O�&o,r#�� lq���LT�8i�w��@���#ݐ�-� G�4&scr4 W}���޴.>#�����F�0���\В����4�E�G'Ϻg�3�BD�W���U�!dp pMC
l4�����ѝ-�Ǥ��� M���6�t�g	��_�z,��	M�|]H��u ��{:����((���l�b\�+�d���F�{���&Y�]�����eQ{� ��֜��` ��;ߡ������3�Q� ��9� \��pK <o�'O���`m����-���L��h��*�+�����&�вn^6>�����W�ew�`u��&YeˑK�G%A�J�]���>�e)�������&��/v�A��Z�[	��fc'&�:�	�V���*�J6�:Jsuf�F�84C�*R�WD��Qe#�l��%f�*H����J��vX�D����y{3��/���0x�"590u���(���TZ��|��sW���=�_4(/����N��c�^��D��<�W�,��+8*�@F>�{�u >��r���tKhO�.�X�zRo�	P�|F���C-�{��������)���O1���ĘPCq�M� p8z�����뢇�	H���[P.g�/�1�'������ל��t���c�9�[�5��31�_i��W�j�Z^���Y���&�����O�,]�Vo!"p�"Sl��\YoK����;9���n���"�D���p�̴]����Ҵx��'�nd��˄��3�&�?��B#*�:�³;��F/IS��źo��Ew���]Y��2�!Q)�PW�삩��h��lc/L�d�u��f�P�Ҩ&�t��Ґ��'��V������Y����\i��B&ǩAĚ�F�S/iͧ�gS`�
��kP+�q^o�q���q������4s��v��n��#����%��H���Q���k��oV�=�ԅ-�� о�+�Kt5~�]����	W-��Ӵ����,Ve0�6Ũx���Rҿ�������=!�˃�(c���A��M�}���'@�t�П�Z84v'O���H˶T��r#���No��.�?���V�Z�L�6;8��r���b
D�{��HA�����'���I(:��\T��;�h�\�o#����Vz]�P�k˹�uO�ץ��kqw0�	���A�)[�s|�]|v�I��DX"7,�蒨qYf*��9����L`R��Cg1��m7w|���E7�%^�1k�7^�-�����h���c�W�79���ߡ����&<bRM6�ot�s�U�E���Ô��)z���JR,A=��î�b���w��!�iw
�aFA��Ȝ��B��Ӵ�'�<^:-��A�J�*��X�v��3i�ۂ`�t��<���4������ڳi\��)�11!�ٰhv�)f.Ӣ�d$�a^I?���Fǻ����v���A|�N2Ι���6U��C���l��r��kc�	�-7�}(\%h����J��e����io���$5y�Yi��{����=��=أ@�=n��sv��y2l�'��1p�Q��g8$�x��DDP|���ӾY�N��3u��p;�����Iy�_�����<)+B��8� �Mr��KG	zN ��>w���v==�Qi��*�� ���Л ��߱6�����YM�)���߅��[e��=�x�H�F4ÛU|Lͥy�h�>�6ܸ�"L�O�Lo?�ln>}�8��&����8��Ǡ�_W�T�l̐u�!M�Ђ��KK�lO�ݣ����_���;!�@��aT�ew�Y�Oå_s�;!]����`�ڶ~5G��)V6O�g}Z�<ҹ�h�5�$&�{�q�4���?67B-/����Qӿ#>�hjk o�ìs���>��r1���݀cv(����_=U�eFG+��J|��=�pu-.2m��V�eN�D�9����x����0�O�T#���4�]�B�Fښ֘�F<`��h
#�#~r'*x�/t�n�&�o��H��fG4	^�yʽ�Ǚł�}~ꙇJ�WC����i1U}��k#2��� +�x
�yU3(�6�4�����(?rP��ZE�0�({_Z�u����|%��ۮܹ}ձ�������}Q�z�������Qd�P��`��`���{��[g�kmni���V�罗)��Мԫ�n$�~����a�+�nn��3�6�Hf���������⑏l��-ZһCi�*�{��Cދa��J�f�t@��R�F�jye?����p�ή8oigg�V��_(pӧ��F�WE������|BD���ڲ�&ž���\	�SVz6���}Z�̼���\y|�����D�V�����0��`��J֤�h�%-+����wC�m+�� ����#%�^M�h��M�$ˈ����@))λ���������U^{h�*��i�>'�w;
�{��(�WP���y��Q���D��Fި�p\.a�w^h���� \IɌ�(Յ�7�#g:BV�=�p
��OXbV;��ލ9Ru��!��8z���	��e_`��5�m6�a-��O�_-s!=��܍f=�?	�A���T(-D��h���
(����$g僾 q���r����fR�KYDg��.�UNs�����w f�Q�T���{_���aј���ȡ�&�����/k���pXR�s��jɕ��Ң9�*:��88����8��U��r