��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C��_�+��+��^���vZ�r�Ln�Ք2���x��)���|�#�1pv��0�7��
=�
�{�J��@ ߕ���Y�b@�����?0 �1�>���*�1(�v��}�c���Z�^L���n�
Ɣ|K��~g߂��Eacz�����Pz���놗T������u�7�s�9m��G���Pi���cN|/$��&Q��/�]Za�l�����\�K`m	ez�",1*��e�6����) �G�DC^�H�0�b���g]�����a�`�Ͽ�.ܚv �Xo?H�6
8I;�8����J�;�%�	����
3۴�����"(j��^y�χ�Kz]���"��3E3"&_�\ �:���i��1���Ω4��W�]q[�p��~F#�t�����We��x���8C�F[^F�`X���m��vg~t��m��zq��aK95 �uu�æf�w�~����kt%�K�ϵ�+�qJ�g'ߢ$(��TyLb#k��#~EC�OH,_�e���8������ e�W-/�/���Z=�s�orw�H��G��WXEi���Ǣ(§5`%�6~�2������5���W
�z�t�N![��H�hi�G�'���GYu������/�̚�M�h��PE�DF�mc�/�\���0N��Tj��̨a�Ž�`��������RQȣH���.G�6��)��0ȱR�C���/u��J��~�+�̪D�r�+5��@�Y��!�_��"����q�J��Ig��xK�����.�^��ƽ��0� �I�6Ɨ�:��Y-͆ �Qķ���!3&�����ռ�
����kݳ �~	ҥ�=�xͲ��]���eb<��s��RW���!�\��h�<S�!�R�1~5H�����T9��K�R\�!#, �P ����ڪ�q)DO�=���%�:^�'��i��Mӊ�	��
���Ҟ����r��B�0���eY{sy�C���r��tҒ�T�<b�+���%Jэ' <!����������p��"}�R6�^���;��!�o���-,�;��WE��oH��`mLV�,}��6����g��Խ34�4���������O0MI��_��y;^*�j�B�� �@Bn�$�� �~��(С�Q4q� ��!��dϱ�B:hI��*
Bjk(P�\��2o�@�^���~6�vA��sx���PR�Yձ'��̫�FNmE�h)hc�4���r��v��#6{�:j�[�J�W}&=7���O1���.�.΂�(�oRy��!��T��eԗ�LV�~V� (����q�q��]��B���֖��d�]����L��xZr�I��Gm�M.)H�*/�z��o
%1��T����EJ�T�����Xz%O0�rv6��;�[���.mV�)%I0�V���Blz���R��c=~��M�S����?݃�� hk�(�}w��y���h��,���X���N���u�[t�����FR��F\�=c�S�����l���s�j�sr�sX:ߕ��<xD��+S,rf�b�i�� Ij>.�y�)��a�)�[��I'�kT�r,c�+d��5 ���xۋ�\o��U�>��g�� �F:�6P�*u��z�v���]��J�x���>_���,ʄ��ǠiM���i��ͭ�s�z����nǒ��bYK���E�