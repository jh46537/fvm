��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9��Z ���ný��M�k�����[I$l�^!T��8���c<��Q�<dNO1f4���&X�#J��Vn�5�]�ȩ�B���7���!3�):������b'���0�Ξm4t�����{)S�>�K,����Di�0߁�JL�Q�bxLӂ���b˱�x��3?\�cA����Xĥ��k�����k�?i7�ϖn-��|op�`���;��������HJ6a��-�<���r�'�r�fڒ����RĂ���9t�_;.J��<�"��+���"��۠�2N���e�r��L��zg�?V�X+p��e��[����dԌ�/��e�_���d�j�͒�d˄*	m�������u�!��lgLs�D�)�N����b;�Æ�n��]r��:��FV��萸F�p��SD����"�s�{oxeHm� �
�x(�Ŭ�;�3�5Z��|x�R�#�ɲ.ز�V5�ΚY���HβU0r%=AY��*�2]n�͂H����ⶪ+�Ȗ�s��Y�ܕt22�e���;>l"+�=�/rÞg�eB������7Y?�Ǩ��rؖ����!/�t�t�v�i���.ʊ���l�[h\�vuQ��������+����T��T#���0A��	��H>�i������+6���	��NgۘO#llua� A�5��R��Ɵ�}�Q�0�I��{�@� �����1vuqf=��=߁3�`u�"�o�ee�N�A)]���$��TG��K�9`����Ϋ�.�8谸@V?n�:)�b4��a	�/�3��鲋@���r躽Y�،��-��Z� B���iS8�4�VM�A�R��,֖W0M1��!m�#K�"4��W�2�����N�ݯ�==�K7ۚط��w�@� u��U�`:�<t���m���VWR�C����&_q� ��*7*�nQ/P>�Ձ�w����>�
��������zш��b�Π�B7TF�Ec丮y�ɏ�kCT��K�C:���o�8����VQ+�����q�e�b-��]�r,u��󑈶�n#�z>E& �U��� Ƞ�)n�Љ#�am� ���_�}�!q�����Xޤ��34yK�Hf�Y=�REwa*,���K��7�dL�ɨ7�e�r~��lq�@'���տH��ۣi��!\Lد0� QU<G�2���/�f�4Â<Ǽ�C��P����tO���s���8�D��gPc
�_>~���Գ'CRˆ����o�	]F��K��ۓ�ک+���9�K�J�������S�b���h)]�����k����p�>K�1J���%�QX����{�J��X��l�`>G��#�DFs,��'ug(�K�^�,��.� @�HR!6��Ch�����s��(*t�������8�H����Ok-��R)S�Y;s�����@���8���'�P7��n��K�˨��M�Kj������EЩ*��c!	�ay��S������s)o癲M��n�xM�B{��i�<"pq7T1A�H�!?�g�2n��ԈF�&���hua��&�'��D���[�&O��`�X�����)9E4obmH͔�O���Ô��{�� B�M}:dO~0_%}�X��Hі1�	�������ai&�V���2 ���]�~�E��?�N�l��S�5��D�N�d��jn�Db�H��'�vwڇ"3i�:4�@�Z����1���y�<nu�~�˘EtO�J-k7r�i��[Ke;�m���n���-*K�ZF���
P��P��;Ws�TbL��<e�%A�"-2Z�|��FF�����B�!�w���)�!Рօu��E!-�0��P*1�Ŗ��\m����Z��u���4�~RƼ^���7uU�R�޲u��g�����`ɗ��m�'r[���y���Ԣ6"s�`�.��������SЄ	���8�Pta��� ��M|��l�qLxp(r���1�]�a�����\��=R�!�Ú�lq���k�!�4��V�D\����ѿ�+J��([��t����},�c<L�%�;�a�=��T��F�C�'���z�j��˿���Fe+�Sǒ��4`���h��c��l�%qk��o�Q<w��9�o�⌊�=����C=���֡��]�V��T�H�Nù�/Z��/G�.O��������Ȍ+����2��j���%�qܢkWd��T�xx�7�Cw]'8��7k�h���}K<�<��r6�Լ��"H�`����L�ڒ^��F|�	5Uw$H�\nCߏO����-S��Gg<#}���x�[�Lk;!c��=��Z��`:�U�y�Di�Ά�X�$V�X�ꢫ�k񺬉&���-��O��-8�� Fz8�7� ����4y�{�q���	�Y�ތ�j��sl�w��%S�*Jv����Ƈ�H�d�dIu����8�'�U<"\�`��d��ELC��mt�yzW&�mT��Q~�I��ꐤNm@�п�	$�x�s�R󯰪g�|�?�u����4��S�I��*=�\f�- c�ݹ,C��׺����[���gS�T�rkH�3�}]��5�D�Q��^ �V�%���H�tj��&��y��	����������ޔr���Ȁf���	���j�:��y1Ǳ���@U�HI�Y���e��9-W]���%D\b�?�-��[�gs��a>;#+h'�7���������*�4 IrZk��)!��TU�~\F����ҿx%��ś,�0a�)�g"��%��z?��~}&�\i�ga��c�;E]�Ҍ�͆HR�N2ρ�k�P��C��y���~��=j4KT�W@��212<��L����2�$������,�b��dڡ��� i�/fHݮ�a"���-W[o韀�w�~��$K�'�� ٍ
�yb��k�(ꄇ{�~�-�D�E�(F�< �B�>��)��7�tA�X=���ը��M�z�E�lm��~�գ"iQZCd'tMa�2m�j��ȍ[��yϙV!Ѹ�}��^���������&x<Bt!�D�<N���XE>��ًGѿ�e�����Y�n=-�4P�e�W�����F���F���ъ\�r�S���7���t�u��s���M[���		a�|b�G;�6%���o{�,:�D��4��n���(��j�������x`72S��/|)H��OC��f>�{������;	��k��EU��ˮ��p�
}�n�R8�e�����y":S��ڡT�!��+��d3l���=j#�7N�/�q#Q�χ]7@;�"P8~D�S��Yݩ����#��D���B>d ��mF�u�A�F>Ӯ��۰�E�:ZyK>�Nο�����
~���Da��k��|�}Nv�wƼ�V����"^ �A���F�\:�EsY88}��4�8خkU߼��ѝY��sJ�6}�KNp��F�����D�$Eo�3��wLz뼚��;�	��$��RkU^�����Wh�9�F�� H�����M��ϣ[���Rq��h]g]$��@��z�#�)$?7Y}�P',�<�ZY#C��qqK�^�?}��́C����B��,�'�{��S�4�K�@�Km8���8��O~dv�W��k�&�	�ex@O�ݩ�龬�1�\¼�] "D8��,���ؚyz^`���c�����>J6dSߊ_��z��Ơ9��1�|�.��o��J����7?C@�H|�KM{��`��8���;.��"����U�]!.�?0�ߥu�Z�[叢}���~�O��؊���%�_͚zk��uN������y�r,��p�F}� �r�XJ��UK=d�3�T�?��l졾";���sF�>Ɔ�jz��&�R `h�t.�a$����b�]�h�~�a��H�d�}��0�m؆ ���?�c,�m�G��(��ä)���N��@�vD2Z��c�M��z��=��=�1_��zoE�G�.���6�f���nʊh�Wt��[ij��V�O�wV;�+��I��޼M�nb�^��Ifpˢ���<T]So���T[;�]�J2���g*O�j���tͯ���T���Nm��+�4�8��h�����P���0}���滄�Һ�g#�AڀsR;����������Tv�$g#_}H��:>s|�� 7���
�	N��.��ķ�v�������
F���g6Bp�p����s�<3eVp=�z~�"�{<�,�oH�J������ɷ3�S�����U�{��9�֚��Qǈ�;o��￁9x�ct�H��z_Ƿ�R��9@�N�wp�c�c2��`6�ml��~�3+�j��Z���:x� ��U����h��p9od� ����ˣQ�{(��E�Ȉ�P�R4��5ΧvD���wA����ǧ���ˈY��B^����@_����	��2#��r�9(��i���'&�E(u3QN�<v�Z<nIZ��T� s�|��Bfbl��0|��/!����z/, s<�����*/��D�ա��WK�o��/�Z ~lk0ԫ�bz�2���e��)	���F��!!0c��88�S����(yg⟢ފ)Frm���G:������*�Ӓ��Q�x�/�Ƹ�r�Q&�iM�cduw4�(��D���;�����9Kf��[4o���0�����]�X>`�{}[H2�-ð���7͖H�#�Hq���ZA~��ќ�|��E�p�xw�Bx3ё��$A�_���4�|;�v�Y�+�'�[��^����q��.ݹP�1l9���5yʳjeh�Vl��gfMW�4�[a�Q�l@�*0���..�(�l��"�Ε[Pb��:�5h���y)��� Ib�w�������J��f��ϫ�az��§Y=���j�@c�$3��tj-���T��-�:v�qY��