��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��x�_H�Ew�8�v���+�Mv����pR9N߭k&�u��dE�8t���g0� �x}�3p�_f��#�`qU6����H�Z�F�(�5�ҫ��	���c�^�W����a&3���L^��F��1��&sŃ�H��cS�w\�gS�S�]�ƅ'iIH5�WYȆZv����j|:�<�q����_Xl-�z�{�syq��:q��)1��f����P�dMee���u����l��ƨ~T��`��b��k�4��}�#���5�/M�^�r��#/�}����sK�^�����>������8N��(z����)7̵:������F���;X�.#F\_� 2k9���X��TI��y�>0F�'xOZ���{�O6O�Q͓�_��B��������^���+58%f�a�,��}��
�)�H�8�2�p�0y_�eL�Z��8vD���I��ĺaLn}�sM6����ئt�= ��YI�l�%�@�&5	&0���ց��O��`!vv�69������T<�3FĄ|~Z�a{��~f�M������T�G8�"��bK�/[09���O=߫����\�H����7�:���GǶ7�9k̂n�c�9 ��/H^9!��i�
�}4�v)^=0����Ҋajr�Ka����J|��.D����:|�_�׵��+��J	J��!�h��0+��'��#E��Q*�gt�36�Rzz<����գ����g�����-�G?��)?��K�D	2�7*������ص���h69*̷���,�dF�g���զ�����X�iu��\�O#%s�Kn�"#ж����n��x����L��ec��uC�G�He��r[��1�S���=T ���1��n�Ou#F��m�Y�/�F/<|/�!��Tqڽ��7��b]�Ef�L����2
_�?'&�!O��N��<�^���XB
h�|�����P1a�&�l��A�	�[�ԚW�S�f�x�8�Iɱ���_�t���@���H��|8�K�U��2rԈL�Ԃ��%�C�/x��m����?�����!���+��v�UL!�.�Ivn!V�E���g2X�x�-��������h�]�I&����Xހ�3����7�L��Ci����K��t�3�e*_?���7MP�'=`��-��,�0���J"�}��e�"0�f���>����#Z��z=�wG���]J_�����1�<}����Veh�B(�����^��C��}�l�,�q�yE3�h ��5E�>���E��ld��4����V�`H>���V������Ey�'�f��H�� ��=���gLh	K�c6d�f"e��I�
�E�0�h�����:�{;�H�r
�ɍ>�f��Bc�p�9��S@\�'J�K <O�(`��V^+�'tS4Y$������/b9�x�4|԰�HK��]ZJ89�e���P�4�X�B�N�����T�s~�l�]��}���ڐ��n��N�[�nqB�G����>2�r�n�wi6?ZD��㣇�T+��W�:}H�7�p�4�h�^��@�Տ�YLd�YU6�r`RS��6�ek��z=�7� X��۫s�Zw��Lצ��N����*{N�>��<�	b%0����&m��~�D\2'x	����c�<��1�}�%�o3p0b�������ϟ�!�N'��&(\��+�H4�m#@V��4ws��w�r�K�@V,�!(Fy%�Û:�ɩ�)�;�s�߳}0�<�Q��s�C�8s��'/i;qs��u�7S�����!�n���Z$݊w�u)*��REI�?�)6U���B9Y/dΟ#��U�Z�y�@�>P�X�3}�N��-���q˅�;��HO�"ᴸg��w��R	�K����$dm�Kz��j�&�E-V�����-7"�N&��M�RXh[��HV�r1���}� �F��rlp ��>�x��<�3���Hn���Gg�B�Cd��~]�N~�� ���@K�;����gq	�ѻ��R\g�uUP��9m�����Z8n?�M@��>��a�sɥ&Ѕj?�'O��P�{�����A��jb��겱b6�"+ �Sd�WJc)��.v�Dv
S8-Y�S$�+�?�bԬ#7�~M(j|������7<ʱ���ҡt�����U��T�y��M.�������Шz��$��X~��ܠ�, ^˄E+�1��wp:@tw�l���{��&�׀&��/��rd�p�������R�_�)j��J��B��l�G�����#��L���l�TcB��J��q2��]�;�F`]��G���W��`��5��|�VG9q�+,�}c[�t�OƜͩձ�e�y�@� \�~޿U0��>�W�ߙJt�à":�l�
4� :����x�I�y?�>��ݑ��Dp���0 ?|�LwjO���e�0qieT��oV��Y���R�bP�K3�o]���ꔐ�}�<��"j�?�Zo!G��,����0j}���E}Dd�6b61�������{�ӛ4,\i�E�h:�ٙ���ِ�7����2 �� x�+��2���(tt��,`�%���ū�8y�n�d7
HW��$�UR`����A��8���Seܻ����5�!G^�ƞM]z��r�f��X ��غ$4���x5_z�A9�����)�ᦛ�����az�<1/��y���C_�>Z~C7��
��i���o���K�� �r�Uw�p�������#\H3��{yx|%�y�H�_�	���>��Z_�+�&�=/" Z�6`��>�E�xC5�H���,G#��
#\5���+�m�c��i7?��Od����{�/w+)���if���ѮJMx"���Q0gq��?��ٌ]�:�_gpiM)z��E�8E���V�Ƭ����'0?@�~��B2".�IP���լ���0���`&N�{m�j>�����ſ��\��J|}�ݲ{T�$)���%�A4b�h ���D�^^���ۓ��� ��Laa7�M���uv��"��	��hV�Q��I�f�&p��klS��B��߿�#4��#� 1k=�i��茄��>A�'��n���<^9��+XYTg�$ڟ�S��o����9M~	��E���mWLI��Te���{�p�J���Y�h������k��I���ؙ*]��OT�h��jNU��j� ��N� os��W׮��XÌ>��{ϔ����㞕,���'_D͵��?.�cz��s+̃b����p�]��b�]ۅ�[[x��j��f�Q��?�� ��Q��K}4��mm`��B���<�\��sa:)0�4QV2bh��t���A��2���D]wL�K�D�l�n�	>(q��,yǆZ)l;�g���N$�#�MG����i;'��Y��R��ܺG�ڧ��7X���	��(DA��6�N��h�&�
��o��-��M��6����hf��z�Y}j8�y���?c�?��a���ƺ�Ne��E�����[�ܞ85�\w�H&���aƴA���2!A����Z B=�ar;�*���H�.��Ѝ� �'G}�"M�A���O|^�� �9��^V�.)�&��D]����6����'��?|��l��[�/�!O��iת��5~������ǌ�t�95n� ��V���?�:����
B!\@Q�P�[��_Z5`ڎ3on�X�\$����5{�o��Q�H
�SGB|!�pD�c�	
�k�3��M�T0̶ mLIU����ܓ���uΚ��9d��cJ��m���+�����+��=V]n�BM�-��N�Z��V�,��� b#��r��r�쩝����N�w�i���Q )jܠ��%�.�s}��h���� �rk��s��{�xB1���xUpz�Eez3~,����G��7��8D+���R�6g�K8r�u'g���X�)�2�/�Ǳ°d�s~ԙ :ְ0bqN�Wmk-Z�p�{���-�Ds�fi�mj��r�7��M�i4��uM��Mʠa��Gb�(=/�}��CX�SS� *��}��JUv��.�H��IJ����%��@���F¸������}r/���"�r�:=u�@�4cԔ���g�]?S�.>V�u�>ގ��ґ��
p�		��x��Bl'������V�T1�s2j�Kr��FL�g2������R��[�@S�+{/7�*��G-�r��.�k��#v�+�ֆ��
����	��Z���+Nq,���Vm9��F�lv��Qv*��pO����6�4����]�e��Z�FPˍ���e��G��Z� =nQ�i������,e�T�n�2���O+,��\=T���آ�HT������%�s������g:�޸@I�$�h/V!ۀ�/��Q�O�1��G7Z^Mh7��i�/��
>��`-+[�L���Ҟ�/j~�����i��R�o�W�Z�`}�,�3�\�/F=�X��~�t���BLY�z��]F'�T���#Q*��4�k4�6f7s���\�w�@>p���5�'�	��&Ä�&�ɗ<�{:�;v��)l+C ��kŧd��6�_S@X�T�R�[~����Te3�	�
��9�}� ~�5@�)���+��"�?XE?�Y%���9�yz���LS%�<��9�T�>]D��lP3}s4+�*��O�:�f���ݠ& O�68��|/��pϭZ��fB��b�?e�l</}��8��7��6�B�"$�`�ʎWf;��|/�/򜂷���vr^�[�_��߆!�_�p%v�Ա@�8�C��X����e�^�\J��g�p��|��9��K�0�Om��+����D�C�U\�Τ���:�}9�t��!���S��-�e�x.G�[�-??Z=��t�b��E uh<�-!S���x���#���GP����2CH2���	
O�t�L�;K�P� �ӌ����W�u�04S�f
��&�O4E��Nb*�sOX�m/#!�&}��E�01C."g�鵖q~�@܊������D��K��ɴ���E��b�Y�����6Ae(���V��ߺ���F
���k���z��U��#koIgP����$:GG��%�<��Hj��\;)���/,�.z��z&���ZK��+ͱ�}S<JL�1M���ǋ�X���"�7�-cυ:����l�3��6���Ivd�����!�݊t���Ί�u�gA�k� D��*8R����x���bw�}{�Ք)�~^>�.]��V'���_Ǹ5�&��6(%��wđ��fkD`"춾:��Dt�����(���ьMV4-~9k{촓̼;QŜ�4yly��]p�9%��D�8��M��|�,�c�bf��'�}}��70AV8*y���X	B��
�f�����|z;�^`.�3�u����#������A�|�t�̽�cK��ݗҸr�4<R��R?0NϾp�R%�^��q��T��Eñvh��Mn1���=�W?l6,��<#S*s��~�?�7����!,���,��q����wY��
Z7"h�ZᐥJ�J%� �6�M*G�����y���mVT�'�&!P�˧qo��Z}���5	T�}�� �RϑP�9����(�~y1��G�C[�H�>v��RK�.��)�p��o�:��SO���>LWd�,.l�e�R�#36�	w/.b�G�9.j�>��͠&�Y�(�����R˜�XuR�z�W�l1-"�^�׬-�m$1�F���6|ڮ�K
��ת��I�+�g	��8�k��R�Sy���֗��*@P�/�>2Z���}}j���S����	�����̍w%��>.�W�V��h�E�%��O6J3*i�&C���٣*�HN�n�sF�F��D���V����o��؈K�5��qi�F�� bD��^�G��O�O��i���)@K��rM�D�VXW4t۳���r��<'k}HwB�ҹTC�a�������v��0����3��Nl^�B��J+�W��چw�i�Ik��״�@dMx����]�ȖS�4��՚��E[���M����eo�df��c�<���n�Ǟ�8�d���Y���lQ$�Y��V!а�|c}�����w(��x��U��)�e-�}�n
dݘ�(|/�6*���WCٖ0�oE��/�|�"���1F1��T��-�����tn�g۞�d�,��e�H��N�G��������	��x��g���~�e>��53AZ{!����}k}�gZ([�5|Q����Hw��O��t1'�g���X� ���H�-NM��|�	�k:/D�����9�6����^�f� Ԅ��p&�]�x�$nC�^�C��Sht��p�_!MGzs�\|�����&�M��͊[7�#FQNk���r/�݃:��1Q���XM����Q��$4ДL'񫨴������#|��d����Be/����x:+�t�±q���₎16*�Z����L��~�O���>]�UIP�B��?}�De~L#r.c��'�Z�5�����]��T��O�eV�CK�ή�
�G_����/��b�[� "=3�-��p��m� ���1֑s�۸h8A�7�@t�MB�=:����S�3�)�!+)V��~������p)ꚉ��ʕ�"hw%����Z$N�e���닮�7�glOT3���0�����u/��B\m3�z���Q���b��W��U\t��]J�X�+WH��v�kV40q�tT?X�����������p)8��Ղ#$V��N=)c�����g�]�00��h���1���j7�A��;@�9QW
4v3NQ�r+��,�w1[_��y�n��C���~y�����ƊW�o�}��u��.i��#�{Z;'n����cn�(	A���-Lɪ�)0���CFǬ�;������3v^3�F<��a�H�f3����)�]���]�I��0A���*r4�J�� P*Q�gE�	_^QO��6��)���t8��k�<��a]�E=~��iG3U�-�#71���O��
	���T�Zg��p�fY~bۂ�A�� g]w���p�0�'�+�<C_��s]<X4UP����L5�֜�@�5�,
h��?�����Z�����=��p�?n|�	g|�6쐻�~A�V�'l��V6Վ�k�َ���C�����,m�,��$�cb���}'Y0]R�!Z����A�����p�5�Gx"�K��Rem��)�IX����`�q9q���r��\�hh����t����6sM`�Cz��Y�\P��M�_+�q���'K���7�n�I0kڣ'�KB]���ZS�4��ŷr[X�p�j"_P)�~�/RS P���YPɘ����o��d pK��,T�M��1����*�d/]ѼL9�)�����q�dol��2��X���_�����ҭ�V-ت�_}a���L�{�Aƣ��nt��6�L