��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�c���G�J�,=N�{�P.�*�@�&��^[��Ԇ�Ă�#�a��� u!��;*ջ�2��n��:#7��l��8����k�D��"3rd+���]��*�a���7�a�W�Ce�L������ ��5u���#��)�g���=!5�g]4�y��t�/�Y��Kw"������u�J�M&
Rܾ�a=�;�D�.[9>��_2�j)���&��%O���b�R#([��%x�E��8[���i��xh Z�ulN�"m*��5ߡ��!���ʛ(k���=���&�}�n	�i��8�=�(=��>چ�����[��/��#�qĪ�7�������m�훓((IF�YZy�r�z}G,mJ��&���\�}ֲ�n��i���*u#R�c� �zP�Lr�U��]o���� J���Y�\�J��_ա叫�#�/��1��":0jO]�T�F~���?r�c$,����Ti�o^��f���eq�d��U[/���s������h~ߌ�o'�%v�j9���sY����2D� -�'%��Sn��x���}{<
��i���y�+N�i��.�w)B����&�`�ܜ�ۮdA��@���԰g�TF[ņ�Z�W�y��t�3�����jC��� �Ջ����4��S�/s�w�,��b��u�ƶ�>��ґtչ�J���F%��j���`���C�3	��@A�#��|���H�E̚n�s�ワ3.���lrӂ�|Q~�]��]�\!��F0�݁ʃ���Z5�;.Aw�� q���p� V�N#���m�R��6���~���R�t���[�0R�Z�aK&.�>����?f����!?��$:a'�/)�P�~w�@��z�G�g	9a�8�F�!Y����U6�<��#������ş�Y��Gٍ2-F0��eJ���XݓJ�a��dgT������� ��1�!z,�g�
�"��2��1�|�kOEV�TZ��e&S[��n�S��� �d@\�E�3����&w̜E����+^A�9,�)��������.T�^5N��8j��{:/����
�d^��U��N{�{��ҩ��I��Rǀ$Ɯ!�M�b!��~��
��Wy?�g�����[��)���lj]�.f�Q�������(AD"�d�*D5��v��rv��+����B���v��թ��� ��)���9�åCC�!��JfU�%�.1�`����nNf3�Ʉi�=���kH�� ���U��%`
e�R�} v�~Ǐ6��dq��wΤt���.υ���֣���gIM�B�r���I��|��]��0̾F����4r���>�������LS�.��@��NY\��`�Ц��(,%ao�!wU���<X_(��u�S%=-���
%`�����CٷɅ�H�`��ef�"UB�ˠh��4?{�>��zm�t���}Ik7j�y��xBA��J} �	/	p@�"��n����ơ�Jf�ހóA�BE̮��GV�H6��R��h�
#A���x����O�Q����7�@ro
80��Xn�%��x�X}t*Z5��W�<F��������Y��n�'`]��:�%���:`���Q�}u�� O��r��0�������[��l����j@D��3{�U��IÐz����jfj�g_�S�pN� ��`���U��_M�/u�e�E�,��@��"���G�__(�2���w
����>��-���⥴LѤT=�N�C�]�'�پ��TV+>T���"y�Zw�����f�7Z߲�@_��ThD�>��(��F��ءz^���B��IH���ڔ��ORH��r�c%\�K(��8��3�f���M<��m�i�� �����1$����&�5�
�!���Mx����՟�c�w����"�}�q�Y��q��R�譢e���">���a� Cb6���l���{	�/M����
;S��C'3|ko@e0����x�3F5	�{FRq+�Ҕn1��X�@�ښ�Ǎ����C#�Z=�9��	��宺@s�B����%��<(��Z+\�9Πc�(|����{�Bj��p�~�p&�^�C^�\o�L�P
/a��(cC3���Q�Έ�Z�/(K������TF��"�}��\q*d�(�V���?�\[�-�J��s����3��"yFx-�V@����BN�M�S����@:��֮�����d~%��͕��f��}m�Y���#-�ʤG)ߑj�</��FT��A\���Ƿ���_�GM�Z3���q�gp��x^��/�>`��%t��§z~����eit����>}�s�P�T�Ha�fq��p`=f�MJv]��(�i�8���S#�,�0����ow��j�H�g$B�D�'�."xA8�'i��&����t�dJ2�y����%yF��LJ"����K=�7�r|.fC��J�AkU���Pr�<6�"�;�7�\����̞��a��i�N`�x���A��G����f82�;+;�{\E�ba;~)"�bj��X|�KE;��h��m>��B����P�����.��)��8��s����N��+��N��3m�FTZc����4�a�[�GKx	�~h/@&�<�6�=�	�����~��D/jf*t�(bVqW-� ,��1��j!����hE�S�u����$���m��K?��!jJ4�_8��.|d�fZ���d솤�mV�Y̙��/֮�W:��՚A܌�wڎ����5��F	9��ΐ��'���\ts�9 m_�|�nE Z�g��9���7%��k��	�k�LW�_�������;��&Υ�\�ɴ=RS����ԒQ�P,|Qג!K��n��a�T�yn�������@/�/
��ПD���A�8�>�_،jԘ���Y;rnЖU���͡�]��ƶ���Sµ����d�ˑ�<	�f!�QPp��(���y��b������sQ��B�#/һ�~اe�0F�5Q�6?ϧ-���}�O���� �|:�{��.j=�,��Y�N�f��F��~4~������밬��,���eu���LG8�.�b�2���%���+�4�V��_?\Q�K���������Ʉ?��k�ă�[�<�⥂�k�?qӗ_h�?ήޥ���&Eb���-9��z���G?�p!�g|���}�u
OrC��x�����!�O�»���745����0�������-D������e���0�C:!��j¥䥊���2���ib��7qj�t����������s � �PLD�������fN/��.�����h�!g�vI�!P}ٻH1�t�q�6���z�\R�G��#h<�+j>�Nie��V���z��#��,^}%�W�O�C�� �e���B���	=��^1R�ӈ�^����z��J�`����Z)��sZJƴh�Y�Fgm �^g��$��$ﰅ�lK�\��,2�G���5"$��5G��<ŋ��3���u/�Ð.�����x��Q��AJ:���g="]L�ǅ���v����{�\�6��/	�Q|^�He�g��� M�M�h�w^[ʌNoQ�|�M��q�;�.������=��0��{����z50uf݃��2a^H1�_�`���Ζ��/8�v{S��K/']�.�������',�36݌(}��8� G�We6IeIH@�S���J����h�e��L8�]��/x�=��l�
�Mɗ;I }�/���N���ݵ�l
4���A�Z�L����ެb�]��uK}C��Tv ��.��%<i����Y�P�*U���;�i�M�fKy,84O{E��{����c��u��ﷻoy��B��#��P�.ٜ�*~���^�� :�w�+|�@��_�ѡ�"H����7��o��O�P�l���w��sIfh�X��7bZ̯�oȘ�D6y������N�P[y'))`����h)15�tڳ�����g=#[R�s{�e�z�k4�cM�i ��)�� dQq����}?i]��.��U���C)1v�w?r��)�j�X���7��:'.Ȕ�[��d��
�l-I�N��hK��<�8Rlcm0E?h�1bj0$���z?M�P��Lt˾��^���u<�S<�Q"�9� K�R�� �Ҩ2��
�WFN�S�	��bap����|Y���C�/0y�L��~/�G%x���5��K츀+�^�s6�;x!���kB�����mFv4�@���!/ŮUo`���~@��f<.G��b�a~��>�ۈ�ɏ
  U�[�՜��n"�Y��s����4�[H([�
��umH�d�Ld��Cc{�4�cC�'���4$��Ȩ��y��+�L���yt��R�!M���V�za�j�֡��p5��Btt$�]���G!t�g6c�&'�0�8x�����؊�_�bz޻+��i�Hr�XO���]Wx'\X��Hu3��/{<��������~}���+�М�����H-�)M7��[��2���:������Wr��+ PEA=QFy9s\3�u���z�wG_�zU���B�0��|�	_ܛ��Me<V���"��c�)u�S��Ą����C7��Ew#+��'d�)�Li��N�(�6隈*ĥ_rc�ڭ/'�A��^=y݈�x���'I���e[�j'B �)��$H���Q�D^�"յ��Ь�:q$��3�����A�Ա��P�ߋ�U���O����"�~�|�NX�������� ��=y��7��z��	�!���Z�B�C���]gЌ�}7�7[�-芤%rU`���aw��>�r�Z� ^�|�3��w�c��,M|����o3R��W V2G����U��j���L��\
�c�R;���|�P�g�j��Q���DXdV�_�cp<������l���(���������Чt�i���%�'��N��j�T�5�@�i�Xل;�e:��ET�<�h��E�ʡa�T�WZf@$�q.�H�LѬ3�d;f����t���<o� �������s��J�Q�ß�Y��e�������T<���b����',��3�5K�ޑ�}���C��
�0�����J�F �^��Võ|'�^���6��͐��|��B�UXcϳ�XؑK+�ms��x&@$^Շ􌬓W6>`QzX ]=��,�yl͂��lΫK(�:�e3^,'��QO`飼�]�Z[���j�����l�����пLpuғ�x
�(�!g��o���ӂ�K��`7��M���6l��TS��C�m�Ϣ�?����6�Ԣ�tf�u~m[�:�w��J�J���مP���$�j������7��������5%�e�� �����z���u��/.*�3��؆��=F���z�N�7�4�|J!�G���n 6x�&>�p��U�<��xX\N������*#���c�����݄���|��z�����O�1~��R� ���A���,w�dP��6�Xj�D��O�X�őӧ�(��A�Ps�,`�
E�ɧ.�Q[�`c�}�WO�M��:�Y_�~�~��#�O:�\�`�ƕ9'��ZqF�T&��6eJX)B�K��k��.r�lD�1l�i����}���F�/����gr��=u�i�p����t��2?��K��~L��z��k�{ى���i�+�����&�	�F0�D���z�����hƁ��S�ࣁQeZ�'o����χ|K����7֜�,6��1Ϙ�y:�f"��M�s�YYk8�sc�/|��I��=�KK�~yM�,]��v���F�O�Ξ��TZp,�&UC�I��8T�К#���b=���ge2Y��F��)�fK��B��h��Ԁ���k�>%C��4f��� GH$�a�!�2W��� ��yDQ�Ob�I�c���J2*�C@�5�[�\�}�I��A��BĢlg��2�|�:<W�[�nQS�g6C�0����8Qu������vl�W����	x��/��l�+b�FK�)E0K�nzn�ο��{)�X��bV_�|o�Gy�[ש*�X;|����!F{[����ǹ��
� 3�y�ƭ�<��'c�h�\>�\��QBD7��{�֗�;��HR��U�6�xi��o�h�37���U�B
c��C��} ��^�|�����V.�[�q��= �[
Q�P_?k��8���]�N���3�X�[e0�^/�e�j�3��<d�"�Nz�������}Z9,Մ�����m~�B��eN�*��ZM%N3J�$��^��a"��K�Bkh �����0���1l@� � �j�)S���h���l���RE΍�ܤ	��>�	p�7@��0���3�ov�!C����3l�t��0ߦK�
�=>������0�3��:���|:*����t�{�g����V�w@��`\�A�>��V��96��?��ć���D�2��z����������*��O#��1W��o�