��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħB`Lr�@�>�	C�k*b���f^��g�{u�$�u�崼�q{�//�������x6�Es�_�~�n�=02Y�{}���ٱ�,�i����b���)�Ag;��m���	W�=H@D������P��>�X�����	�GsFMsiķ�7���~�rS%m�?�$R�,��VŷG$���ި�Dx���O��9%�q���kn`�3H[�e8`$Od=��Rԝ�)R�mxt�0��hOL.�\3,���*����=�� i=��sr����@��ag����1�[�����fg��(ڼ\�ًU��ȏ�����e�������Q�%��&��Y:
�8��|����L3����;͝T�l��1ԿkW�ߴ�|t&��D"XI��Z��Q����7u�r@㻹:�%�ň��+����>p��ӘBx�b���D*�/�KW�0��(�{�6��.z��hrf�3=W���N�3�q/M�H*�z�b|)�ml���e�����-f�����N�0�W�/�<b��*���T���p/L���l6�19�u�3��{�t���4��.6���ݲ�q�SK��&�b��[�R;�	'֙�pe��}�ʚ�X49���ڨ�oG���V�b0V�SB �M]S�m�o��i����5wy�|E����9bр-LQ�����g6T����*ȌA�x�
�ޜ.����!'� ��e�B��uG~�\>N�)��KN���V���ͱ�H����m�9t���в)	�ڠR�.)�]���R�����w���-��x͑\+A�3��vI+�G�, �	?�������8
Țt~8P�� <(a�����A��f>�.��d���@���)sy ��D�gd��v#�\ȭ��e���	`(�ai�B�T�)����6��.�i�ɥYA�A*M�j|�`> �0�5�v�=�y�xRJ�rW.�G7��z�xM��4��9$כ��Y��"��� ��S�@N��X�j�r���F�)�C��5���riՄ�<�@�C�7;K6@�M�l:�h��i"�Q��G��G?{L=���Q�w����4��{��C�/gi6��MK3���:�"ċ{��Dj������L��G@�ߪ�����~g�SA��f�V�O��}�� �T9g!�}������@�s�,���Us��z�v�8��D�|�z�a��,�:�wp��E`Nu��H�V��>1ぴޤ �K0w��ł�ܓ$B.���m�$�V�yR��8]]ƋBx� � � $M%��͆�0��˓����x���/ȗ��mH,���yG���PEt`�%x�jL�Poe�syiN7�>�~%�az���4Ӻ������z�����Ixn���'��3���p_�v����C\��Y�{�&T��Sګ�.{W���8���,��
�_�2�����if�,�N!o�o
_7Ba�q����iY��g)�ul"�/�" �^�yZ�=7�bJL�3��A��_}3���#�ֻ�Q���S����en�2KR�U�敃enk���1v�O^O��k|�qV��@�;��_R��=K��7�?C����Yo�Y��Tɥ�fJ�MB�A.��H܏ �Lw��D��|B��H��@ ��~c0���������@�7�k�����]9H���z���a%�M3�9��π�])�v�(�*hG��,��fo����Qid��<�i����0��((/�g<����*����0=X6�L|�M+%s� �� |�L���Hz� 5�_P��M��0X�T��at��#:����Hͯv���U�,}a����r�0 >[��OI�o8�b_<D�Y{k���F������PE�d�,(�G͂���j�!K�~	C��kY�%��7p��c&�៭�c|����6i.N��B�Hb��j�ы�C*�����z���!��VyM��?2-�A�PF�3��vY�\� �<���S�l_�����P�V�C�CL�w��oNR^��rPYgAʹi��\�4;~H��#�f�}�1��
�.h^�C�Vq�i;��g��t��������o���iE�ǌl���
�1֏.�$��cX�͇�6��U�yERF�B��/��?�;�	5yE�ÑDRJA1��s2�5۾LC66[��-�n7�i�p���-��������L�Aófb��܇kW7L#Re {��%�:������e����]���	���w=$z�Xʥ��J��	\&���c�\.4�G��*�|9��`�hM������2����vj��Ӫ�k���Ŵ�JG�	�绝5�U��8Z:�Lp�}ރ6}��xZ�г۞��{>5�c�����p}5zYQۻ���+SHs�+�!�
��*	]��=M?A=X�������&�5�?V}�BM�(�T���i��m���:w��y��U���d��6�m�=���+�VE0B!2 xM�Tj�/�G�xd�[�Br�;G���z�a��zHjR�e����r��r��{ȓ(�<�CVf�Kq�ޔ��O4�b���K�����������b0\�8G?]��i�@�@��E�^؅��_������j�e�V�0BF��Ӕ�<o_p}�+	ˎ�PCg��=u�|YR�8Ǭ~a=��̵��M=��t$���<G�{S��k�J5+�\��ߋM�^R�~m33к��Cc���Xw����N�upS�<_n.��|A�콯�T9ڡ1�O0s"���7�Љ+aP�ݡ��T��V�J &�pr,��y��E̓A�w����7���A��)ZU����	�<�&L��Ƴ��q�SF<,����� p��2/�;r�*�^8E���y�Y��ݒ��Ra.%�7ꦽ����h�^�o�4�p��G�֒�x���gf�a�G�&E��\������eJ��	��Qɀr��9AM{g�0kHvд;����'-(E����{<�?��`�w�S�3w�mc����k��r�n�ԁ�%L�i&s;f�A�ɲP���F���5�;R�'AN���I�Y$'���^T��lv�ظ� (�J_{l����2kS�9���Ʌyiª�w�hU�RC ���&�*m �uЖ �c�,Z���e�.n�W�,߯�Ay�� ":m�ZpA���3��YQ?�����}��ꃷ���.�3?�K]t#��4I�๵�^iO�1㢕:]'kN<�h}���u*����u�+#U��ui;�q����aD��Yk��w��D �?��܌��̡�?��_�*�"�=(s�.c�Gd+V�2��d͌f40V��Qz�` ���Qh�)o�3
�':�-�dR�% c��ğ�Y�.Z��)�P!N��	�k��:�9�'��tP���ߡ�{����m�L<����L9!ј~�4ԋ�h�s�ʬNc��Y��<h�w_ן޿CH���4�K䘡�̍��;<M�&T��=�{iP���BÜ�EQN�{|:@�!,������o�ܕ�N~ ��h���6�����B�RN(�
E����Pd�V(8O��E*���L��J�һ�:��	Ts�i&�GXiyo�XU�*$=std	Yu{�]�6�(L>*��D�MTZ�;�'=k.1"�qr#Z2�u�����رwS�0�a�ׁ�>!���_���Yt�����s0P�oF�Y'1�=��Yf���Ϟw�����^��T���~�ẋ�P��V~@��ӥ�B�$y4 /���FFr\����-��R�����f'QY��gU�<�ۙ*9dr[^R��V5��FDɿZl���h�o��@^�-�e����6�*�{�O�e[���RIw.i�$d�+Y�����ͺ�o�(�}'�$ނj~� �T2so�4��kh��kBdsQ�������H�]Y��6���Mq��.���g��dJ����b�T�!�]*٤��O:t{Gc�_'��C�|�<��B	�8����0������7a\K���u^e���s�r߽<l)��&> 3E!����wM}apW�4���㩶�_��[�	�d(��SLd�B�ŤS�iQP��2�#������ާ��UA�99��������2ʯ_ ��1�1? �T�ޗ�� �/�W��/+7�Z3̱Ó �Xa�������[�\�ٗy���YR��`� 旑2	ɷ?RD���t�!����+�l]�v$��A/!���Oɷ��@�i?���I���T�:OU�[N�w��{������[����ˁ�����B�y��H����`����u�������s+Z@���ȩ�-����*^���l�e����7#�;#�
��R4PY�oO�:o��_el�om�b�
�H�ˑ1p�z�p����<@y����c�+���04"���9�� ���E<�bdPʏ8M~Ʒ�rX�y����&���'�?�%-��e�Gln@RS�>�A�$��8kuڧ�oB)��_��ѡM��h�ݴ.NE�'���5=rY^Z���k�8GdOv6p��Ö@�A|���>a��l���:,���?���v�8lp��X_�c1R��N[,]��y�/{[��"��� wtߍ�~�/��`��5��F��A�|/�N3��}��'J"�A<���Xa���$�(4���~�|��{{�]�yy<�]H�2�M��;��+a���'��E{�qc�g��(mf��/�(��x[��$mm-��u=��+%l�#9�
m�ل;�k�,�8��i�a���LƬ/!J�L
�CZC(R��
㰰�A{g�c�$#�d�"q�x��OTa�z� ���a�㹫B�gPX*{hp��Q���L��O��[�X����:M��s�۾��0��XJ΅��
�1����586�?�-U18`��}:2K7�M��G���oE�q_C�`BQ��� 9bO�!BŬU!j7�`���(�9�[�n�pi�K��l��pf��/nb�C1+l��{�Y�	5إ��G��Rc�n$�y��xů%d�.��H)c�yMj\Pħ6���/���EG08�@y��-k��z�m��Q>@<��x�c���A+�ө6����j�^g���a+=������H���E��;|r�=�(;^��.������r�C��Ri]Э+����Q�\�U.יRKA%5��.C%`.���>ȳ/-�c�-��aMǃR�qs�]Ӟ���>�Y�c1�w��Z7w��i�lL-����B9������;Ca�ƿ�m/�q��3|�2�X/�2酖r5�������j�� V�'��z#8�"4z��no_��=*_6_R�!7T��h�FGƉ}��TR� �yR��,���-�O�������"���1lB���:�J!,�����n����B~��LS+�N�ﶯrb���/LG�����!����x0vn/ݝL��0�nz����Hu%Ϋ@y�<���ui�f�9}V��0���Q�`�Y�"�����ׄȅJ�:B{9aèсg�)�|��`3 ��d����k�9OC�l��$��\5o��S]�z��e�=6(,9��L?Ɩ�{�Õ%3IG�D�|\!Tƙi��oqG�� ��2��J�g��EX�Nݏc3�+�\�ߐ&(4�8�x|�M�%OP��$��^h��N�ti���Tj�{�^�#�VQ`+�>LbWL�`^X��� ��+QW�p�����ƙX2ʵ�#q�Z7}�,�N�sKis�}L�=�I0]���6�8��˹u���9R�m�mՂ��;_�l[Ir7�wXൌ�c� G9y�%�G����fL�@/�y[?L`If�z�!P�s0۫V��4CJ˱�7��+����dj�>d4N�]��`��gjMߟ>�b��6���%E����R��aR��9`�����������]�j��޺�>ۥ�O�_��� � Ue��cyn�R�`�{��q �h���-��礝/�%����$�L����� c��=��J������Jv������� �'k�� 5G�F���*S"�잃�u������4��8��*H��B�`��9�$��S���@se�����~,5&��2�54�]�M9b������R�%��"Ӡ�	��d�C�r�i�8+k��.�r1	��,NP٠$�gەz~�M5B�m���A�f�K�g5���{��JQ�ڻ�V#���Ȫ�:� f�ÁT5;���녑u��6Ϫ�2K��&F�l542A�B �6� ̚^��~~W0��KJŧ��8P�����rπYD_�~W��U�8us�S4�^"�	� Y���}m�@��������ު�D(�9�\$�L�cs W�VY��Zp,H�������*��H<y&'r2���f)�V8d��~��K,9��!�g����-T�	F�^���;�1��^�f>�u<��X��y�4����Os�+Cm^\%&���q�Jd����FK���1���|�(�\�% �ZS�4V��D#���*&کɎ6(��ct0�,�X�{x�Y)l��^`~�mΨ��[@�z|��\ U���߯�m%�z�������E/L&^����s���o��G��N�(� �.htֲ=ECPdX!�����!o��C6ch������P��|[�6�z�K�q�� <��~���%R����|��r欣.��K�بgF�<���M�Z̼�%��
;a&XU(LO���Q���Q�$Cx�}_F��:�<KD�as�:�FM��&v\��b���f�tu�f�#@���d�=�O�t�B�"���,�
�9��"�����#�\j|/7�X��]:���¢; ����D.�/l���ʨz�>�$�N�j�_*M�8��|!Vt�~���ﶫ�J�Dpˢo��v�^$ע��0�j�&��涯uY�k�ʐzj��Td�/C���N��K�	U�V��5_�դ��?�[�@1j�1>�o�
g+rU�K������.�	��7_���K˗g�%{��ft�+q�8ρf\&�3K��k��G��V,$U/wnk���A<j�-���W<p.J�j��'��dL�MW�L]�;|���*M�_��'�6����Ѿ��)�ڿPMc�v���e)���G��E=�N���YP��}�;�jQaK�s)��Gf���ILoܜ�G�}�-�SYM��ƣMwz����� #���_�Ћ��,׾ɺ��QJ!xb�k:�LϧJox��n8���T Ү'��^h��5�Re�*��t-{Q�f���<��k��E퉖pztg-ʲ���+�����5���X��`�[�P�H,O�%�+�&pHwBGK��DJ>������!�5����9߸��F���R�����|5Vz�Y-×d�7��7f��a�����~���A�����٧	
�~��@�
��,��*���i��*����죀��`�����
�$��;��m��PX��\��nL���ZZ(K~5t&�d���v�W*�d�>��M�y�O���n��O�RS�L�2�r����m���s3$�\�i&���Ǥ���A��\����*�_�sL!T���vq�;V��@�K[U�t�W���1�-6,��i�勀��}X��QYE;�Y����X �\k��Jt��:w!�*PT�@._��06���=����C$�
E�����e�Π���="p��r�k��_u��,�4��g�L����Y5��]��>f
J���1+~>�����S*�q���Y�i�VU@9_ �23��g~w�@fG�9cZLˬ�+��;�H��)�;�27��E��)���?��b�|~3Iy��1��2k���V�_�ʷ���+GL̜�� �� B�{G��p�Co۲�{Ae��GT-V�k⦯�b��o}��q:F�i���/k�Sdc����{�N�r��b��R�!�ܯЯܛ�f�ز]>Bo�V�3f�F�ȣ�|���v�j `�s#�&���y�;��զ�Iٟa�1պ�)��q�y�]��_Fe:���e}U�~T�_���]����1^KP~�p�r�'�Ֆ�CfC�6�����x7�U�.��q"�1�L�����.)��VB�����b���S��Fx�Q���+��cY�^�+�Nq&�;WL��������G_#��I�7���
�j:~`ӀJ<o��M/��LeY�a�h�MR��k���i�_q����[7Ĭ�d�ED#�9Lp����vD�_z�b�,!'�͛ÒK�nl�����`�,�-����>3٪�M�1����P4�1��YU�@��s�A��XT���������Ң��̵Tȱ�[S�U��سȯW:~J\����\$�pP����ƶՀ�pxʽ"�<lUDQ)�w�ͪ_&�0�º,�!h������"1?ὔ)��Z�����`��t�k�F�J	C���ܜT>�`I!�cN�W��h(�p(����0"M�l��:�����E�
����f9[<�����F����h�Ҫ�@�ͽPH��R��0��9Q8%?�?,��"���2Cͱ��3�Q*�P�ĵP�fL�d���t��b���W�+��-R�{Z�yIH�;�p�N!*�����M<�]C�;�	i�_�^�=n�0K)n�b���wSj�����_�C�6!�
�dH��\�k�L�	 ��y`a]O�D�9��mF��~�%�\{��A�B�ss����'����Ӭ�*����?X���bg��htvv��J��"��E^�{Z��j>�+��=�ڍi�S�WG��ƻ�.X�0%-gS9���	��h}E�?"n��]o�h�ݮ̮���3��7����+ST�H�Z覇�z�P���@��W=#X|Ca_�&3����[�b��]�Kũ�yP���#��A?��|������[P%2l��������W���\�	T�*�8e�����������+�\1l	02�s�m����ȣ�Uf,��P�osW��r�c{�J�C$s����鉼���<~�x�\9S��'�x�k7��#�����?�?E���YI�D�c����=%$���8�;mn^O>�0�/��Κ")��Pnx�:!(Vo�䔖�S[w[��"B�v���+�Y܄��R��e��5r��	܉���������I�����@��j���:��t*���)�Iه����## #]]��'L�Ũ�j�_�Ǧ�&�6�1m���ě���?�:D&������N����!A���A�#�BE
���"��=6����F�%�v�i�fe.��#��B��-��`����Q���^�<rW���E����I����P]L��
3���&-�'3��V����8}��/5�n�`
�xˈF�0n8��P�����F��oP0<t���ө��I86ŝ=�����tj@q���M}��biq��L��?��.���Nr�N����)I<�M�+]�3F޷cz�M 4�+�8��K�s-4)Z���6b,��#��v P!���-��4���Ny��{�����gR�\7�q�v�فU�����"�8�񸡔1F�će��D(j�a��ad�x\�4��H7	�2��S�p��F�L��ߔw� / �#2���Um�	g��QɊ)�*�iy���E�(*�UY���`����ZME��Y�������c�.5s������B1K ȇl]�>s�J��oV�����;Z�_�͠�lC\oFX�L8;s
Z��O�M��q����3~! �����ʁZ\|.(�6��D�O���g*�s��S�%�����1�^y��_�,�sw��2���_?