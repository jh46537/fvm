��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,����۝�gW�Z7��?$J��w=%g�?`ԝ��# et�L��#�e�LGtр̎����-�0��EA)���y�Ff��J��/��K��>&~��Oe�s����b�C��H�+ɛ�y�reVE�+)��J4�tG�o��\3QL�9m�<R %��z�9��K���~����ZR�8H�0�
lr�m·[�ZE�rU�'j�B�4��m�e[���n��q�[�RT:�u�`�7�>7��<���d4�\fD����}����C�����TdXw�J�9h��U���:"���XI�T�=�y�fB��9�����|{�W����mTto�����)F�)��������5Ҵ�hOꇄ����qۙ�e{��p�?�ɰ;O�Ħ&JV��>ο������ɏ,{��\�&��R�S�GC|����ĳB��sإd+Y�<Z%�����r
��$�R�k晷�i零%?d�+�_'l���.t\.�z��4���x鶞T�� 20�/E�fqǽ�[��&f�����S<s*���7���=|h�snM��T��7����v�f�?��sej�7�k+�<ry�?&�e�܅S�I)E�[�̴�G�͌��7P�֨F��;��c4�![-�7Ms����z�Q�|��������B�
x�i��K�T�RtyOmI��2O�p?L��$�I��\k��#�G :�o��'	lb�f�S�GiI7��b���?�`�-~�Tx]R�~Ps�gt�e�����r�\V���hJM4�a��C��΄Ї�N�[�%n^y��K�Sx��R��\9�qc뒓��F�Kf��;�8h�#��z�q��I�C�l�z��MT������ �<�X���@�!6TT=���f����!)���O�A�|_e�w�ՠn��'=��{y.����jҪ�$�\|�Snz:S_
��-�� ���2�wb`38D��OB��Jn#����p�4�³Fm��3�ƥ��_��:C��9�W�_xj�� ;t
�9:d's���}�n�z^�O[Ͽ1�T����(����|/� Z�0��\��'���*n��OѧsOdT%0]�d�G�Hc8���g�flZ��cv�i��h��s�7�\\A��6T�7a�%*A��P-��C�C�t��)����7a��o6�m���E�x�~���dz��$/��sn��یe@;�L�h�}��i-�DJj2���fx5������S��z7F�X�h�3yj��6@3M��roiD�aV`GO��H�|v.қ�g���W�ۼ�g`>-�	��O��T�:��~\�܋8B �=�:Ƀ�E�N8��BԏNr3��4�o���OvA�x2(�++h�.���}�13ep1-����t�=1��/<���@�-XY�K<~�X��$����|�1�K�����(��=�U�y,"6�l_�gq �h21Ż5<>pp��b�ʾK�&Z2~#V]���'t/��fa�De&v�a8_��r	.4�oЭ�duc?����؟!4!��5��O�x�T�>]�{�g�|cJ �@70�헩C�-���߅�S���n�9����s���;���Q3���{V7�P��f�F	e&�F��3�"km׈�O���Y6�}�(����:�|lш}B���?�m��*�Ŀ>A����7���� @3�a���\�J�?-�+����D.07�� h��y@���������}�ܲ�	3��D��=��Tu����PC���?H�h�m�C��>ѡ��e���x<=<w^�q���@Ϣ4Y��s1E(*�7���*>�$A?\�a��������_�y�v��6�*bS����d0ޭ�1�A2!e�f�W)��/Ep'��ù*��j�����������/Xz�1z��|����O�!b����x�!Y���l��:��Y��r$��-�8i�{lI"v0	�;�e)�\U2c��]���t��c���1�&�0A�7
��[lOҺ'IӠ��`3�8�Kڙ1�&��z�f_;I�%��6�H����c�k���s)�V�pF2h���h8�G�8��q��
[�(L;R�luP�c$���D��B��L5�[���a�n3���ȕ�bU��H��+�s��<TgH