��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z�
�xpQ�	g�>�)5�Ը��Rd:
��01���9��6��1�s�hU|2z>�WpF�T4��.��=������/�����KwGl�anhJŮK9`�œOF��-&������9�u��pe�JdV^'p��@P�b�����P�{� �a�����Q�l�#�"�,XB�ރ�_�W$�jç����?��O�vO����	��҈m����z�ݗ2'�{l&vHG>h-�J��a�N�aA�'�[��H�b(���ꊡ�ۆԃ3��Y�E㗋.���OL���H��=@a���;���F��b�	T��7?��XU��_;�?~
 ]W��
 D'�:����}D>qP����� �Vނ˿lm��z#�s��$ϛ.�c
_ Cϸ�B{��ִ�2���g�{�L}�g��+��2�/h�*ݞ�J��] �/O�2
Ԑ�L�i�zE5���)T2�hX�ա��0x4E/ю䌫�'�f��� OO���2̼Ž����R��J�kև�"���=���.���>��+ �z»j�z��l�3idց^IUy����u�[��s'
���o����)�$� qˈo���ۻsژ�x���G�Ky�ڶM&�aQ���(*dq{k�����@D@nM���(-:q��L"7Z"RK&-
J��z��_�v���,8u"��@5V/exGe�VՖ"kw�r�S,N���԰��P����.����Ȼ�$ �"�D�S��U1�j��hy�������GA�ǉ�Y���r�����c��5��OC�A��{�a		��u��n��v˳�N]<�Z��"�hw��x ~��E�k�2��EG��ȝ�*���H5�k3"�7?�{.����Axi�X���D�x�Kv���g��n��4X1���~����ߤ�>P_%2�*���ݲ{O��'FQ�d�p��5�[��С�s�f���ڽ���e��.�,�U鼽|���<~@nE����!O�7��:�1�6N1S��z�ȺWz�/Y|���;�VF����SJKB�]�-`����t�p��v�%X��	IyM�ȩn��đD�H׽��]�����f�1���Y�θX�ᰞe�A���j[��#uE��QIF��+#�Kc-�_߄`���}P$��?j�tD(���q�v�0X�p��-��r!�h1�g �#���d�����S{[���ͭs\��4���X?H��I�x}��nۄXkܭ:��+��-�)7�,�X̳r���%�A	L8�������z�h��g�2|�e�Gu� ���u������ g��j<ck�C���`y�cw�h7�/X�ᲅ5N?��6���7�p�E��l�7�Jo���\�n�<���1���W������Z@Uy�Jͮ5��U�)] �%��#�- ��Icv��Z�#���Ʃ�R�K-�>!F�P��<�����.hgH; �_O7�tU�UX#ĹA��#�|��&k����Q�����ϴ7��n�^�;����|!>o�/t�q:C���~	��g �0|�Ѭ�}��q�^��q�LO�@�@qWt�'���<G�0c���Ty=���b����Zݲ�8խ�i�U]ug�}���P�Cn���<���"�=��M�18�;cDY����>�c��vVս����*�79�1�[��l���8�&2�K �6���qK��8��W�s���,b(�M=%�BL+�~&۟8u��`T����;�e_��o��FZ��sG�3�Y�|'j5���(n��w�,t��ҧ��si���QԪwKI���	:nr� G� �̨�څm�}4o6��어��w�q�!
��ɼD�0��jMZȷ�~��+r��D�)��Ǽ�$��ү�٩E�������S*ej��I�G�=w�zW�]@����ɇђڵI�no��y)����$4W���z�ݔ�xA�93�T!���S$Ŏ,	ңKÿ���"��B�5k�l�|��b��_�ʰ=�@6	aG�@�k|R�����BM>�]X�\�3��bG�hlڟK�^.n�P^8B���cJ�����ۨ~��U�D��h�uU���+���ǼuH�%;<q$�Jfp�/�3&0ܙ���PR�~�ˀļ.�2��1��� ��:
A�cW�H� h!D�m�e���q��o��*Qգl�Q��6܇��1�!.`�L�B�W�AE&�	AF��Y�*L�41�.�=��v��4�qw����o�aO7�71�8t҄�:�sm���Ѳ�3����c�tt�y��R��)�\!^�/� �,��]u�%�H,y�YCƑ�A�-?��]�-� ��w.qD�t$�Zs�i�>�\�2ݧ,��΂���q��u��>��t{ۋ���_�O��Z� Q6��o$�iP6H'˗�9��7C��a�X��n�0F���
%�læm趣}�����B���_
�0}3��Ｗǳ�:آc"`����r�f��V�kYa�t�2��3s�6W���{E;����\�f�t]���ٻ������kS"�>3-nӭ�w9I�
Q�t�,9��~$��\�y�3R����b:���3�-�<ɾ�Q�_���X?Q��T�3���hTdl"������|1Yp�
Bַs�����ka�FEA��)H��6
��ZBn�2~l�x!���-�\/PɆa��&��r� �K��UueKȂ�2fY�����)�����$�h�z��\c�Z�?~Ł�O�������\:w&�J�P{ ���n��}�K��P^���4M���!ۮ������B�n�H$�5k�?����?x��X�cU�wLd��%��B�js�d�F��3ۀ�ԇ(R�����$4���d��L2�}Y! s�G�F���ݓߝ��;=��2C�Ӎbr���S���^8.�*}�>.��O�)�!��v�'Nݵ��9ۗ�;�	�TJd�-��'}�N����1�8h�U�>q��<w�����|��g�x}Z�(���Z{71
Z;�h6�ys�I��k�0�>z=B^{>��l��=~2�! �w��~D{0۩�9��������N�w�A�	R�Z�p ە�7�k�o��zb�灗� ��������^���z�-��C���W�xF���t�I!o�ʽ1�}nΝQ1=_��o{��rS̗s���y�ݻEimivm��:=-�/���(LѪ:s}�������Ƽ�-���v���8ֳ�.:Z����f3ꝱ�o��,i��M!N&�6ny�*��n���YFp�%Ť���98@�Xv�
(߶�c��Q��Vk;�j�꛼tSޑ�[�W��9(wU���_;Z}q��Xwu7\�Q��*	f{����3"i���C��f�R���<*���-�.*���=�BE+�]&v&6���:�'�ܗa*��2^xV����A��';d���l1j"�xn�����`�F�;Z"��'�~��d �|玩��g��k��ʑȤx��;h}(��VfF �:R��|�g�E	���g�`0���޷�Sn�ϡ��g��c7b����*�9d�;��M���]�*�b c����h���Kn�9\k-+��� ���=�_'K�]34���o���Z7sW�G4A9@� ��2��\_���={����f��sP�Mn?reə2�m�:7��b�׆x����x��B(Z�&�H����z����w.S�.���`��lS���ۓ��|�����69�Yxd&@�f��}rc B��d���J�q 3�
IGy4��,�m���M��[��j��¥�S�~e�"p�ŧ��?n]�l��s�]�u���#N�1�d?eܷ���c�0$:4�0k����oE:?/��p"^�բ��+Q)a$�w�s�P��"#I���nw
���NR(�=�˱z�:�P��7����`
[Nh�p��?f��&a��e�ͧI��\�������Ӥ|Qkؼ����Y�o\p\6�C�8�S"�m�K�'�����oO�"��9�g.�����#�&B�k��N�q��D�̞][�˓]=@WL׏�a��R��g0r�H> ���C�W{ZP,�2�P=��R0�I^j�oF���x���)�!f��"�P�H��[��})�.Y��5��j���e$	x�,�͖�����x5��K��G�^2����.F��b���r�.G܆��L}e��k]<qq~Ǎ�}��_���6=.mAC~r��xw��Sy@�s�:�h�^9~�s-��7����jݤ8��U))���i�8��-�[�����0_x�a!7�ڔ����ᯌJ=�*�`I�}�/V+�՟�&/Gq伱��3]��cL*9�.�̘CӢ݌��^���D�J���y=�����~���y[p�����-�! �B]�B� {8(o��e���d����<��Ձ��}Q@�`d�K,��H���F �������e�2�r�(�
�+(.V��8��f��T)� ��J~K�k�8L>G3���jb~h'��=�G��L��}ߛ���X�U��#�bݽ,���}y�鞼*W���{!	,bz��I��k�FU��y1l�Q!�;z��k֬�) �ˋ�i�~����w�h��[�x��7�s]G�6C?��+�.�痚���cs~���,Z;�ͼR���a�����cl�ĭ�o�l�$���4$%CLOqh��b��V�G�1����t���ӫ%���D����Ři��.�X���D}��z1T�fu�}8&���&��KEa�#��2�wMs�E�0�A�$