��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�������s�h�qQ Ҵ�pp%�bs�!F1���|W��ٍi�\��չˇ���7Ge�+��9�*m@Mm��A��/f��XT��݌��GP�s��Ɔ4)c��f6�}jwS�����r��j����Īf�t�8J�gmdD����I��h9EWC0^����T�
�we�g 7H�����2�^/����t��PY��Ivs�b�q@>y�%K�~���*0p�w������
��w��{R�8u-C���_f(ZG��|���/zg��P�sIY+�e���<8%���⌚��8gn*rp,����_{���W���J��fM����D�~ۂx�Q|�hCުŶ�_����[�����������=�՞����6�����o��B�#A�����4��5s�32.�^�`�!c菂Q�h�;�wטvm���Jy�#�d�d��_ǫ&؁�	_�%[��1QݢB�&��sთ/A��4�,;�w�����C��k�e4ƫ�z|��<�I~�/�����e��4$�	��j�u�ar\_����U'��vB=���*������V�L)�ߛ�~��~���W�x{*#��g_��;�����f
�6�{`y����O2ιl_��,v��[�G�c����1c
��:��^][F�Z��[��Z�6X@���<
���Ωl���M�5 ��"N���m�|���5#�!MM�^���=NL}w�M�܆�ݞԬcݗ���0.�+y�{$b�5Y�$��8IY�d=���Sgf]8'e�h�^mG��8�n��b)8��R��;,g���oA埘Z�씽8]h� ]��b��o�vS��O�����2c+�1ſ����?���)b�]��	O 6����0�P�oH�O?25��vc�<�;�Ck2#�(i@Y�-���%A8k���̏t���u�'k����đp �)��?��q�v����]@�O�?�"	�#=b�pI���O�N��K�L�_٧�}���֋J�2-bGe&��Zh�P
���o�G�x��Jm4��4O�8�US:T턤� Ĺ���h�,F&̥��:���ܐ���� Mg�a���{�P�K(((�;`e�([��)�3S
�z{~}�F�\���|(����o�t�������76~$��F#$|s��3΁c�υUj)�{Do�HZQ{�x^�c�-�\�d��dy����ۥva��.��VtȦ(ʋG�E!�m@�R���%�y�^n���ό��;�"\�5_v�`�ݒu�g���V ���<W�����IϢz���P��R�B
U�9�B<�������
�O�R`�f��OǬ��Γ��I�9�ߺ`�Jt��������lef�Ϊk�𔘖���*��uG�N��ou��4��ѭ�-��t���J�.)��N��Ϻ)���[O�ϻ�XjJ�2Y@���i�N���!�ՁVW~�خ���5��,T<0yۭ�\g��^�`��1���A�}����.�S���@��7^�Ckʚ��{�����QZ�EfW����D[�$y"��˂JJ������B��vF+�Y�VYQx+5Q�0����-��}-:�!�J�Dj(�GN.���y ���A�+��r�뜔�$�SZ���o|Y	��̆*��\zt{�&^��[����z�9�C^_4���լ�f��.����3���H�B�$�ϡi��j�|?�������/W����IX��i�gzz��HEZ�l,8���q̶� ;�n|�(A�}��Z���FC[�w�������[�Q9��RP�>�q�i	��YO>̡�=9A����r�&ֽS�@�l�����b^Q�'x� �޾C���޼��a(7�(s�<���͠�L51���h�%����o�� �z=T�K�Ğ�oJ>�a���5�Z��(d-h��-%�=�>\K/]dٔ?b���I���N����_��%� 7سv���Pp���n+D�
�Ly�����H�w�GP"�Xc�6ۊ�48j����i��zQ�w�wk���3���Q�c�e�
U���f���	�6�_�Mu �=��I�/ !a��˯�"�exC�tw!D�
�	{%����I�s�e�w�^2ɳ���w��Do��.C'����X˓+w��z$�'����[�1P3k���މ�v�D�.�,7g���Vz��{9n�� � #�����U�� ������E��\�F�A��Vq��X|���!b�]����� ��(�t�Q�G)��U���*����D�ڦX$�=]п�!��]^C��v|su��a^��8����ɉ�"Rv��b�QP|2�R��_���٪�Y�?�ķ��a�B0�� &)j��s��Q�r`66:�m�?/@��[O��R'�k�g�)]n>Vfa����Y)��wp=�L���nO���6�"����>�I�=lt8'��)��7�7^+\tD��ϭ �G����Rf_��X�e��8j��S�&�i�����%�Wז�a9A�E|뛴������_T�'�HHr��d���n��"_4'u�N� �Jجnbʓ��PN�<���MI�/���i'�\�_�Re;E�:��_Џ��'�-��E�h+�`|˅x���-_�᥽d���?,�/�*S����x�� 6�)����VŹՎ��A3��y��+�1	���^��N���D|��aߋ朣�����?���9)�N"�eav]T8B�O �屮��uP��W�Ф����!ch���\��e�@�g8��l��8��4\��)��B#SA%����rW5�ܡ]{�� G	P�mM�aõ�E\TH,xݿ=�!ԃY�N��pa���V&A���<�����OuL�x�޿�Y8�i�0K�!债�p8w_�u���8e������.�)��*@3�[�3>�sԓ�4�s��q����@\I�Y��ߩY:����W���	7C�%���.�꿓����ٮgٳ�ɯΖ��Z1�׫.�
�^g��9��.��#��l�p�1:F�I,�Lcdg�%��[U���=�G �V�i뢇�1IYL��C�l�٭����mP�Q)�S'�A��<��ݦ�����]Dn4~�kEgyZ�b���=���*\�A?&��n[̾=*v���;h��.�CޠC�M�IѦL��k �1{3���� ���C{�l)Tf���1��;�ƾ���t�q�oVm��ت�A����%e��M��u�c��%�_�cbs�[���:@�Ԁ��S�#��<�;�a�ʝ!m��2��ԅ#���{�w����& ~X�ƾJ9{mCg"�4�߀�R�䶝v�7��05k�W��{����P�M��D��k �
��ڐ�c�ٿ^4"�]�# �oS��k)Rd�@y�R���d���f�H���Ӣߓ��٫��u��eb��̼x[>�,O\*�_��Vj�2�_��K�]L���n,�x�(FV(�6O믅:�Q'������W��ק��U��2Y��M�E9d{�>�0Ӆo���� �9�x���&�k��Qr`��]�-
��
$s@L.��=9�N;��P��{�@��F�f�k��<yì�L��c����{����g�VT؆���!�u��� ��e����69^�oE�Q-��;7������h��I��l�iPR\w����=��+ȱ�&�9���2s�wyꀒ�
� �ř[z,>Z��r�Q;ċz���f4�����M�
�Tʓ���G1Q�\�2�S��B?����:|��L�S���oeH�)���~t�i�t�hI�x�÷�y�[�3
�B����U �3$I�"V�"8��Q+�UL@q���M鿔�r��l��OT��[�|��M���a��Y�����2�Il��wj�K)e�I�:�`�#�3��o�ܓ|S֥��F�ޗ�'�**�(�z�cu7�`\}�t��x(��2��J|ȵ"�.�=V�O/���nu���D��d.A��&ֽ���t����b��C{��d�d��Ε�=�o��=F��U����Av}����$�Q/j�t*%���\!oc���򄡎���Q%cZI�5����dH�����B�ƚ�P�Q@�G�/��J���)kFL�ON/��ِj0�Z�#Y��c�b��:�fӐ�RF�U���eNj��M��ڝA.>�&�v�\�`-���vH���jH�#D�B��ޗ��b���e8�JK"O�ʛ=�����.���L�}d4a�)����i�x���{lD�r&x����t�+8�e�z g-�6c=w�q��`FǢf�mf�.p��:6�O�H4����x���k��}�������r�j��m�`H,}1��Oű�&q���	�P�ӆ�؅9��sbP�}xRXH�2m�^�|�����(��a�˩ݯCW�����q� �����n��@�`ݏ�PH��ʺY6C^�fM�p����6�%��6wz���2M0��:��5�)�VȾ=�L�;N��J''uS��8���B&��7��UTOt�0�����ǯY6�!F[k^Q��!����↉�$��F����u���,�
� ��{�xdA?/(14,Z}��*�/0���fC�@�u��e��w8�i~n��/�6v).�]rnHn��*�sGMZR��_�Ӕ�7ם�qY���#V�������ꀿª�k �6��&�6��K ���Y���o YD�z�������F�"��)��z4W���W�>�T=��FxfT�j<�d��y{|���Sb2�b��#����\�=�HɎ�զ��_������(n�Eむ��
(<5e�*_ݫ���,"7�ak���di�TsX�Џ�DAށ�.�A��� ӏR'��_�����d�3~"-P`Ŗ��Xޢ`&J��{>~�_b ����H,�qB�T��x]oR_y�pg����I��B�r�!���h����հz��C�#�R�L��-f�v���s���DKȤe��T�a������������_l��:�2(��Xf���
�J�^KىG{{_c�N0�^���'��FAA�9F�.K&t�Ҷ��������	�l~3��>P����x�����d�z��)��Trrv-�t"���,Ec��w���m��ެ���R�����s�>P�R8��S��W*B,.�]����UA���9��Ek��+G�-����mfș������`Q�k�S�%e^n>��(�1}���B�F�2-��ƾx	�a�����u,��A|�7o��f8��o�>���Oٗ��Ǩ�1e�??�Hw"n<�E�b��f�\˄`6�=�t��UBH��̫K�aB��͡iU{�2 0�i/pE���H�;m4O�����C�	?���e������� ��ϡ�}�}v��zS�#@X��A���k���u��[���S��Cx��\��&�б��`�UN`��,j�_@��Auv���,�V�aG�)�ӹ�Ɲ������O�)�׌��K�L�v� 8���T7�� �c����\frv(y �Y�au���$�X��	MH�gV(�zN�CY��5I:wDc��EeBϹ��}�=�0+.�/�f�m�{���Tc����W���`��ʄ�ҭ0�VpO�8J����X�O�.kr�G�b�����h��;�W�����|��P:�o��h��r��Z��N�U
z��M��Z_-Ojkȃ�	+��^Ѯ絠� +���y��_�)~�]!��Lii�$����H�ʝ�'�B�zHJ(}l������p2�^ex�>a�H�a9���]���
���f.��8��6�BlJ��.P��֭���f!�2�w���zS�������t96�֡s�~����6�&�Y,�.	)כ�qÑҬnxs��9��<��kS��H�M	�x��"�x	-��y��d�Ӭc�����O�E�$��OEq�c`��_4�w�l��^���مR�XKܷ�v'K�X-㮂����^J&9\����W�A�N�C���?��3]��9Fq<�$3I�Rj$�y[��;�>=}�����+e�.�%��Nv�gʌ�r,��AG�2�w�v}���4'l6�p�Tu��1�����6sZ�^�kλ�X���5������+��nٞ�����J*&&���`oj.�<tc?�T�6�ov,"�7t�q�G����wr�rhz8L��Q��yݭ�m�e=�~�V��]�Grh�Ȯ�S+t�N�߅��goj�	����+���.笫[��s�M	4�.�/�o8��C���)]�u�;K��<P�}F�&����#�.�'��&��<�k�|A�l/J��9��G�g�:e.��yb�Kb�2J^�ѡʏ�r����U��g�vY�;�٪��|P�0\�?v���£��GȢ��G�a�g�
�m�b�[�$�G�����>^c��I�u5���)�� !ҰB���]�7=xY	a��~1��[���l�� �E��������Ұ�E�$��?�x���G��q.�,I��2�� ���m�J+�& ����h�ЌXC�>�t@};R���¬���[�����:z)9v2c^XF���*:�K�Ui+f8��Y��7�=�W��0�`f��"��&�Hm�n��u2CZ�n�f8�����:�$t��3'ڠ��*��޾2�~��|<��<z9	��o|���s'�T;F/��՝v=bՏ=�Y��&�Q��޶r.x�	��G�д�KD�>(y�f꽛["Z=�j�1tv�H32o7�`����|7�łdyD��$$Y�êk�ь�8�
e2��bcn�>A/�î��"��t$W�Lw�$�Z������[��O��b쩝BK���a>of�u�b�K���g�'��Q&N��<�jrB}��s�`j�g"�xTI�26�X�$�<�z����u1���l�-��-$�������%&��<�����|��=1��2_
���|�ֶ�6b�C�6�F��_��O��O�C�\�u4��
w0�J�c���(M���v�׋
��L�:��ĩ�r����$�ؠ9(�V�[,dp&�ς�t�T��1�'G�اF�JQ�wo�ɟ�IڽQCW���e
�v���P;No�@�ser7C�;��tͣa��g�\M��]ДX�C�v������2\��x��R�"�R����X����,��Yy�(��|��z�Ͷ�����D��}X�C#%���,�&�Kwf�_S5���:����D�F6DZF�
��J4���- P����1�^[k�h���H��uC�s��8X]$Z��3��x��+��+[PS3�����op{�(.kI>��~
�?�x�d�vE�lZ�\��'���b�؁��V�8���/[]��rDI��s���%1�`Gǳ�$���,d�g_�iuti�>�΂A�<��ğ��YD6 ����|ip�|ag�m��6��43�s��X0'ŅA����I����;�ƻ���Ԥl�H:�'��_�֤l��ceM�*;��yqݒ����/&1� Xv�S(�����=s���wWv������	�/�3�[dj�!�n �N�7�]̚��ˤ�p�[Rw��6�E�ju}m%�y]n Hz��m#����&�JԌ�6� LG4������nY$�O�쟼pe$/3�J/�Qq�ڴ�8��� T-����p%�I�sK2cu�U3᧻snv1q
l��1�Q�/HR��򫍞�.Y�^�Z��j7
�x���;�{[���k!�rQ��~��S#l��-���ŷDZskEE��s7�x8nY��H��������q;��O��^��wx�����8�p/IL
���ƼC Qi� L��蔂��G}J� �]�P:~��H���|�3�%��k��_+F��rޭ�9�K�b�S�I�87f?����\]G���)�B؞d����u�����mo�.{�m������Dg��f����>��+v�(��0�Wrv��r�&U�ւ�4�C
������/���h���R�F�(eh��Y1Z���{#/�pO�LX�)��������˘Af`���/�R �յ�vn��T�ۚo�ݳ�%6~h+���}�,�g܈`��iC���B�M�dh�ȫ�VH3�\��ꜫ�p��:����;���mΫh���|�`�v׶���E�B�V6D��9�?��������HU�v��h�ۉ�%!��ux�6�Sy�P(�
�?�V� ��B;6~��M���`���ԇ~jv�q����2V��яlM�fI�S��`��?yk�����(�^̺)%`	�h�ȴ��g}�����~8r�"U4�;
]��o䌓�&���A2�L��֫*E��p	�nk���$�郡�������U����`�^�,�J��N�e hC�;�w)&��͏��{&b6����'z/�PJ�F�
�=�~!;'��jU�93P��T��U?���'�`���;�S^VF�6�8�U�VJ}.�7����w��)J��'5\���R3A����qO���SD��(B���|�b��Ǆo�zl�%-��lɗc����fle"Z�����������faGS��1C(j8��'�F:�A�G�v�*7l�spxY)��ĵ�ג�WCk������m��|qȄ򓛟��N,�^��½dϏ�B��A��MH�t�ȯ$���I�=��r�5�Ԅ{�ea<)}ذ:E.4��icRTV�^P�j��Uq�:�h�|̫j@R��@Ǹ�����^�ѐ�jo�]� z�����ck�=���cT!�E��1�F��pǜѼ%��+.D��8UZ*� �B��:ݚ��l��iSW;��عx�����	��'%�m=R��m`#��o>��P|-זּ�I;��Y�W�	�)��'�s����á3����e�8.Ǯ������E�byJ�Q�]-�[�� u�>Sb��%�z��r�훑��=�{	�I���aE�ͼ��!M���\�K�!~����r��䄜_�gT'P��%��|��J�h������g�E6�~����Z���8�F>��E�#��bqlR���$u��hi��M��]���CK�P���R@��L�~5���Ku�#[���cVؖ3�n��q)�[דF����=>j��������Gwb6P��d����Ll�7\�g��4�~��a;O˓��m��2P��S���X�[�v�&iZ ��V��mj��:h���EP���2�;ފ�n��.'S����W[��l�心��D�%��YE��f�V'�q4���T,��ְ��%#թxF�B�wp�1D��� 1��L�c�6�>��/���T��`�%u�U6�P�p�I����|�o0QP��X"���]	����H�JV�ِ*������U����y�P�͗j_#�edy����"��G*��&qC���8�G�+���O��T��(����8�]p����l���9W=';�T�ä�g�c�n�Qg��U^�nbN�5f�F��U��L99������j��	]tF=vb�W�~8��$o��'� �WH���VҏC�́����H׍��1�����B�+]
��L�����an�6XJW�ɾ:�m�f���v��\J�0�t�orm�Zgpʄ��멣�_r۞?p?NkX
|��,�{̹+�Ӫŉ�Zũ;��߲J�7=��v�~6��
8�Cp����\�'���:߁�N+�.<��m����_Z��\�l+�g�I�Lfʮ��.3�T���L�6��.���?{�w`=]��c#Zf81�O��C���~��w�f3Vb7��C���d�v3�8T��th���R,��*}�������$�
�@��n<�(�Z<��#����F�F���	����%��O�hX�U��*�M��lF8����U��|[S?; �q�|5�����|��)12C�$���'9����>*���V1�;c�.��e'��M�"��v}1��h��R��9�8I�n��0�º�:�����O.�bq{��kG��u��\x�Dk��ɓ���d*SD��6ϒ{X)-�p9}ʮ�z~�>��:���_E����_��1�e�J,Ų@�� ��V�H��wn�P����������n�Gi�4� /+�?�9#��7�=�K�v�H���g� ����p�\�gN������z:�h�uqU����!��8n�4��<�{��v�b`Nm�&����ee���F�K��~I��.�&��w��%�*E��:��P�y�x�A�"ʷ|��
�4sZ�H�.Y��s�!��B�{�E�m#�ݬ�����˶{�:%F����o.�R�w�իE����;���E�*O�]z[��I�XW�����De�9L�bqC�ɫT�U�Y��P�nݲ,Q�c��"���ι�,~��7+R_J����)E5����|z$g��=N̿���Z���z�0���`���>]u��^#�R^�ÁԪWl#h��z���:���SzkJ�ňȃ�--x5G��������2�����WQ�V	Ek6)�<�f�_�ZS[�"O,�bD���ؑ�]�;ê�w'�:b��v֚���.�C��%� A^��<~�Cm��T`
��,:�gsDD9�+���au�ʎ,e��7�G_8��X)aNJ��/�DPB�M ��ȷ,���P[Q��P��w-�O=6�
�t
ϓ�n�yZ>Y3�Ws��62�[O{OC��j�s�-�"�GH���K%�����:�,����K��P*\�˞-�?	������f�����z��-X.QY��S���+�bm�,~,��K���T���y�J<�
�{�C�P�+Y@�S�0�8oV�;���� ���<X��?
W^�zu��f�T�42yg�K�e��CA�nt�#�5��m�U>��'4I��#'�"���N�=�����x���)H�p���F�,+����X���/']�N7zn�م"f�ğb�ct���J���Aԟ.��6�v�╇I/I�>���jF.o�#���_1/��-a*�Vx�H,
��T�����dɒQ��Q�S�B"[i3� ��E�]��-�!����e�u����n"sx���'o��G�������	^L��ɴ����U`�A�f)^k�D���w��~����V%jtN��E7�Bޤ�����"����񨊾]4K�"/0.}?�ԣ��C�?3	�t�"��vI �7�)KL!�Z4@YP�K�ǎ��H-��	�\�jGx��CO�s�+#�՟^���xR���IjN����  �{�+��]H������Q��/z&װ��q�p���=z�����p/��h����-+�@	������K0�(�|�&O�%3���39�?�;��V�D�Zꗲcu�k��$�6�U�mٞ�j!Lr�Q�@EU��c�����hg�LM��nXn���8P��W_y3@�gn�7�le�QARX���Y|"V;�i�ԁ�n��w2�ݵ��w^y���7F�T���t�Ur�P ��"�cΒ��>����I"}��>	��$��ϕ�u�@��g˞�b���f4�����x��T�t �D�.3J>#�����I�ٳ9M�����<$	�C�]!d�%����VR)'�ޮ�M��J�"���9|��+��F�>��<�����;0 *#�&��R ��x��}m�59|��A�cP�X�-�.x U���#�q��aƀ�6�ʤ[�p4kD�4ڴߐ���f�DM�Z0��f!43��S�s%���t����EP�I��T-�������5�^�s�܈�
_���O�yH�����b�p��\�S*�����q�6C�C@s]�����e;p���I�1ƸR�9��w�a^�9+ﱎ��b閌�ko��J*ވ�	������`����_&j��^^�L�Z����˓j] �?�����b�'�H��r<��������Y�2B}HT�,�q��Re�aU���Rxo�Z�@#
�u�z�	\gt�,� � ~�'*��o.C/�y�8ܳ9��% t�x�,����Of�
��"�UjV<
�ו�ia��7�&����h'��]s;�ǲ=��[g,g
#�y��qU��m\�WDrK�=%a��t^�6�������w;��v��F�:����_�I5q�bg��s��=:y�>"p�1sDF���+a�R���5"�	��;�g@e�6���ss9�N��ȓZ�y�.amt�/��@aǬ��t۲��1��W"Rd��&wh�m��4+��g�-^��ECi�̳��ڕ[f��}���c.z�Ôo����K��d=b_�����	�V�H��� �`H�/m�ۉ{|��fu�����5��Z�f3Zj�<nI[Oir�l��oo�6\ ;�KPud7����#Ѷ�0:���к�<x��)�;}݄CY=���K�h�z���3��F[�?ʉ���|;�u"���zlH��q
�m��KdH�/���.�\E�N��3v3�$*�3���fŎ&mO1OO�'���F�3��=Dhs�

�V�2��R:03�����+]�Ҧ������sf���E���Q\�q�7����2���R�����֟S{x���d��UpoiG���(Z��?����O���5���A{)3��}��4���0�'f����������c*�ɛ(U���o �XHρ/��}�X%�Z	�7(��$�<�@��~a^A�Ou��,�ƒ\��B�P2\���J���o�ú��7q��J-D�k!���>}�Ժ!4��j�h��ݝT��꤀ɵ�G<��w��2¸�}������_��Y�&�|Q;���e�~�Ø�	N�Q>u�W�X���+�W���}uPM�;6*��bIٖL���<�� 3�d�q/Ω?{g17F�do��u�<�W�""Z0k��`�OB����'e#0�L�<���s-*]@Q3zm�K>|&`�a����%��]�^��������E�x�!y�����k@���+�'�8k�jq��l�R���e|�f�>�P�$O)A�Z�'ɮQ�ب�T^HӪ~"������=��|U��h���E~S���l<����T���G�{��3Ƴ���Z�H=OU����:nN�F�sa[���T�B���w��Κj�"��%���&�}6v=�3w��?��9Q��8oS/��%�ǘ�_#[nF&�Gb�R5�^�F��*އ�T�K�%�H�����9u �Eu��d�[���e^����'�Ѐ=���zg9_	w�jC{f�����ҟzW��7��B`h���
���G����THVj"���w���)3�OZq#�8�[I�;�8��[�7˔�֬��q�#��e�-"ui}0��VH�5l��O� ��{x�јS�c��YrH��#.��)s����G5����e�ۍ<��Z{��Һ���g��M^�BD`�ήجW;���:~���f�ye�o�o����1)db�-qT�Lś��L9���4Ű���#�2c7qqۆ/KO:�0�?���ɖ�0�>��!���S�����V��k�ˎ̛��_k����F	��"$�8�[5[�h��ŢbzR��9����k7���e�*��V�[&BK\:V�(ۈ�q6#J� ��u��Ý!}H�H�t���Ҽk.2ev�J�/ry��������R�M�<��>Р��#.��-Ją�%D��(�0����]�R�q����sC��d���[������<K8�w������$�{+ꗰ��T�)ǈc��7�.w�E�K��~W�؀�p�����q���"N81,>�u@fw�څYYDTd�{�ą&�������E�E{�x���T`3k���K��|�������@R�{F�@�8�IM|n}@����-�+�;G���S�0[7��J"�9s���oL�m�K���^�D�PĮ&!��>]�\�<�n�X煯/�_I�nc�Ad�"x�:%({���y��Ly�7!��(���]�_k�q�ݪv����G'����,0T<�w�&�E��I�S�}�Ei�˘���.�ȼ�Pg"���I@�A��ޕ�An��t#A����.�+5��ʠ�E�,�&I�4�[��V���ʹ�[*u�\��#���q��" \7����Tހ�%��+T[/8�Ogf � ��/���]+*s/�\���%X�T�y;���;AX���`�I�cg���|���t�B��0`�o:ǃ��t�s<?��f.ͮB��g_�A������)>�P:PD�V7�N��ju��AE��5����ߔ�jG,�C�����Z��������J�o�P7<O� &��q7.�8��/�}
��qӏ�(}TuJP�IUZ�6�`v������Jj�6g�����)o�cE�b��̝����!m>>�ܱjF���Un�]Ӝi%� z�=�{ț�����v�A��K�goJ�u�悡�+��%ջ�tK�%�^]�ͩe�M�e@�J�c�T�3�[�5��ŀ��8�Lt�l��).�R�����"�(^��h���>��1�,%L��ͨ�]�}�vq�z��Q�J��糎�8���P�C��IO�g�����J'T�!~�!#^�
�8����J XR����Jr���x�P��ڂ�d�"O�{��4�zDS��t�~X�D�����,�4��;���k��o�:0�}�b�l�g��њ#y��xС��W7�a0�f8�����u�5�������#�v!<������� �9Q��(	�,8��R:����4�/�a6�Z�qR�*��{�3s�E+o6��-6��VV�J/>��oڠ�䲹���nddJq?
A$J�%��&�IQ�*�Deb0�E��'8	f�خD�J������S#�(|�u����ު+,Y����#���Hkm��0���������d�=�J�AH��ZPK?J%�,���đ3ȹ��n"o���[jŚ�sG_�\*YU��IDuLR8
�uFϭ�h>�t-�&7 hDuk�ܷ8
<+��ϼU�y\:�PvYh]~"��#Q�	��Z<���iJ�j��&���x~ݘB��w�5#}�����W3�=`F\��0�o��)����|g���D��y�J\�
��3Q�A$���a�+@f�2���D۰٥����J�ޑ䡲$�P����5�>I�[q� �1W�ˉ��tl��3��ƪ�}�t��� b�4��"ل�X��/�D�������bWk]�qD_4�9eEE�\�+�q��XY�InT�Y%w���׏%b��h�MM �
�0q�5�J��-�5e�ɰ�)��N��#"���UfLT+y�?F-�l��~�B��b��U3���q��'�0�y�u;���y��z.��z1�f���O�#��Q���\-���V��#X�o٠o�>����_�:ۉU���������f��������|�]�,.l��֬d�X�:yF<P �G��8 y[�!�"N/m��s���i>�N�2b�y���(��u��i4�ц>�T�2l���$�V9cpUm|���J&]ѽ���{��5���LyA�A^�r50���B`\߯J�߻�+lS�؁X�G�\�.?��(e��ZɄ�������U;���6�z��j�sd���`ؕ����y��ԌM|+����GZ��M��*	�q�dHB��.@Gڷ^<����$��ٳy��r���S�|�J3y�D�S���j�R��Cd|����r�hNgw�*<5q^��S[�䰾Gޞɒ\/6j]�vh� s7$�����p�zA4]I����U�ف{�B�������7Zy�r'2���!�f/?2�#�6s���OFi���i�K�tm���.3��u�
�1�b���1��S�]�e�n�}yK]�@$��;�c�����nē��X>!�y㯪s��B��I��q�/z��$��L!K��)"LG �(��9.:ZL����^N.�5����A,��3�m����V����b{�����o��CN�z]�3	�����C�x�����o�ݫW��UKֽSL�vh��Jm$�!�ߊ���ٖ���]t�Zٯ��룈C��z��JQ��:���#Op�3��� �%* 8 �F>�C��ѹl��V��F���z��S�{ReF~e;qg�ѩ���+~9fN�7�c;jԺ������a�2'��w��boQ�}�U�}�hU��2B��(�[iɧ������&��U\Zp@_yZ<7�e� �z!��vc�z�Y��Q(�I6Y�~�+�?|�2��S����'��f={!ݻ�G�`^	>�6�UqR
2��7��hꘄ��9�ձ�
��z�����P�cT���ٴZ���g���o`����a;����*&�o�G$={��]�[�J͊]R����w���b0�5W
�f�^�!g&d/E��&Zm���.��Nj�H ��@lB1���{�S���&	f�����v��O�K^@|�Vc�a�D�7��5ҥ�H7��5)���_���i:ί/�_3�ʯo��O
��4�'�T
Y�2�xF��~�^�?����,�6�[s��+}�
�m,�N��N��X�F�
[�����5��TFN+�R0/�Ul�&�N��s���83ۣ@��K0>&u�5�,�s���)U	�@��r��I��Jg��KDP�\-0�S�u��#.��֊*��*v��f��Πɼ�ʕ[�֐�wьA/_/w��Xqc�G�φ���<�t�{e��}m¶��_a����u6�1��c�x��̤�0Ok(���|��͎;�����;����\��`��"A��Vhxc�~��?�S�;*�R�(��O�gP}�Ͽs�ܗК1(�|�����l��2�	��5���ϜBU��������3�.�pf0N���.J~���զ7;�����wV�#���)�[��)�aw�=������nU�;�s$L��F���Ȣօ � y_�3�2�%'9w��ʧ���-��\}�/@;D��}%�A�,B�=�:)X���jC��9�:}��1���7�c�S�M�s$��`��8C8D���*!Pu�̈�©��ĭi��F��V�Y���aS��k�~��PY�<.I~I[�IY�,�M�5nu�\��qr�ᩱ�Ƿ��f��\�kx�^ �fMd�x��_]��B=k��T�ш�ʲ~������7r[��4X���J�_K�%�޴��'8�8�F�WCW�1�;�����C��a��C0��@���|��t�����Mj���)��~��Bî�E��n�l�̜D[&��2���ݡ�����"�d[eJ >a���nfL��
K�P�+f���*��V��CF8]⏑�>�<ؘ���z񰴜'y~e�.!�y�7��ᙼp3��*���{�(�*�vzu$�@j	i+�@�����Xe
y'=,�öe��,d8>����L�uH�-���_gS��|��S;�t�������y���z�х`]�]ĝ(�h8�Z�:�$�0����]�D)_4N�9�.�D����ӺL� ��
����������ZE�t0/KA���Y���*l���?��Fe�m����M"��g�(Z��B�R(�'y��d�&A��������jɜ��|�YDB�RdTQ}���f�#��5:Le�\��' �~�H��F�p�o�F	](	
�*���s�I��� �!M�W�A+���# �O�)��*�)���)�wn�>�e�)C5���%�[
�Z���Θ���^,��a>r�;�r��U��Nzް�[���	�vPxwT�\�υ����?�G���
�|�{85�ᾘe�)
�w��c��k�C�(5�	�~�K���7���{7��y�{�핣#ہ\�M�1\]ju������NS�b��&�XD^/#��9�!6X��m����La[� 8��y�Ь\{sS�Q���`��q65��\��O�'�^�;�k�0�_�����>��m��B���.R��.�8�\���z��꘬7P| �P�!U�Bi@��k�yH^.p����K�;
P�C�=���"ͺ���f������Q?��'7�3uw��+�[��R�P$N��3%�Tn��5��͓����ݶT�+;�~��MPu�,�wC�:x���*s#���i�,�5V�Gl:G�Qc��ߌ4��R�%��W.��?ᯬ�j����7&�s�M�W��A���􆎠��9(���\bg�t�%	�Dv�ڴGĨ��$��rC��4��#�k�wp;~��j��;��022�b��MH�\i�/�%S^��|�b
$O�>=�x`a@��꼈��l�Ŧf����Z/>���OshH2�
��_'t�(���5�+�˩Ab[T���n R�2�'����%s�l����8W��a&�.�Z�z�M�pE��\k�w�x�K�>~��&W\�.�2R,.��}���I;�6�@i�%������lɎY�5��iMvug�����?p�=_j�=�2�n@�K�V���MJ���jU��a�Ju�*ٙǆ!"�(<���|�o ��D�D������8
(��*����J�J���� @g��S-���Z�=G��a5���U���6�F`�K�+�����>֙k0����xvj´�Vd�db��+�rdhc���=��"��cOC^�rt���t��a���t%s����xm�?U�cP����-��h���}���p�z��J�q���:5�㈟��Xו���39�v�L��������*�;����m�!��D�G*EoѤ;-�j�(�bVʠ^V�i}g�kO �}��s��uab��؀`���^4�:��+w!�=�1����
��0�A���4d��M�$��eU��C�������Y�4�p�� XI�Ψ8���f�E��|8���Ty㲿��e�P�&�{���U�߫���oB��,��ȼ�*�ꯃ�"䫢�߫>����� �k�	�����@zA+9��,? �5�墸���`�Mo%(sG=�6T�BȰ��.��9w�yI���uij�-�cZ��;�L�-ݽK|�(Q�����b.;6]��T�X�P�}� `��u� ����٥L����<p��g��v���.�(������5:
:őQ|�.V/��x͎�T�o3t=ʈp�Ǿ��
�o'�ё�F��H|�����X�qe��Y+�f,�C+#J���+|!����F�LE/#,L2��<�q�o��im���&�VXG�o�uM��1	�05�*$T��� g�UO�:nˢF�$����6�-9��*�}<�s�+�ײ�0�,������:�}?A[�˵3׻s`|yj�:�$X��hQm.�!ր�X6m��F��Ԛ��a $vS�F�V2CƬm\j��1��<�`0���O3��� ;T2'/��������d/�s�����UX� �2����H�63���8;�G�1����Þ:�Z�Fh��`��ݑ@���>�]xǐnwG-3��F��$֡]ZVsmZb�1@�������+ڬ?���h�����ĸ@�E<nL�����8F�����7��nz�_?E
�h;~�����C���
{P��vn����f>�d���K��0���K�5������	�ĥe��	���=WET��@��uEUN��'��p���*�+����'>_��K"&�00P�K�mA7�p�e�TiԤ������2��hEﵘ���3�:�&��k`�:����	)��4U�b�ֶ���<��ggڕ�"&����Ј�� $�^g$�:?Dm#In��t�'�0[9�<FK���E>$t	�E����%��5���zvYTZ���"�1��-F6%��Sv���b~�3?�9��N����NCSG�%4dO��	|���3��VS�a�bE�Jޟrɋ���.f����9Cl��������{�Z�G����L(��ʼ�oˋ��=�%w��uf��g�/INh���*w��;���<��ϩ�ۇ7�t���9w\?937��k��׏�7�bl��� "���
f)�"����E��(������E,�\I"�Q4�����5~��I�q�ݐ��p����J���HjG����;��LZa*X��;��5E�����f�������㹫��$���c��.X�tr���?�� GN��v]h�r� -��8�/�nxˎ+w�u#J��.�PhF�{�c։�N�Z��`3A�6�/�xC�Ea�1M��8@�d�P]
�a1vq෴�TE1�sJ
eǼ��/�a������1���)2���_�$"�	H
<9�d%�[�;y�����WV��I�7mG�7|S���7d��K8����ԉ�I�m�.<{VdZ.���>$�E�������hC�z��^ޟ��)��6���L.�5r(_�D�#R�gd;:s�˝��`&�Z~RJ���v��Ѓ���1�������s[��_�s���S�s�꯲�zr�KY`Cqo;<>��z�X���0��a��IM��X�`PLD��P�O�|H���]��#�|��6<����d�	���X�O٪���䌾3*84h|T��v�<L�V֠��v7��L�(�@C0*� }:ㄺ�٥��x����EN�&���@�X���������wDZg�[^J׃\�}<#gbZ/���r|OF��l���g�BS�����-~����M	(�¹���_�PQP2>�m��a����-އ����A�!	��� �#l��c��9�_Nx�Bk�k���趦t�����M����L�jI����G�n޳��hR����	C�j����yz��]�n0g�U8��;1��h�|§�rŸ�l ����Md[	�.�����iK��i7%=K[���0xA�D!B~R�����0�6"�����2��/��3c`�f�O�ظ��̗�� �[5��� �)�������8�t����+�.	��AM�"�^�"�[-��!���~Z�}f�i!��nB�����^�W��Y�_<v¯�������� |�xk��} C;�$,�B9�A;�%�=]�\��<^q`���l�ͽ���![�Ą<_m�N��#fZ�wcOlY�r�{\.��
�Ϳ�	:T~�Z��<{�h�.)��HGP��Ek�C�/]8��\����+����¥X�d�v��v���|A�S|i��|,�+�],�1�Y+P�,����3�z���&2�g ����f{��4n*i�5�ho�=���Y�`~�I^oY�ĢA\��)�YK�Պ�!6v;�\pL�%�m�t̍�>ނ�9=V�6���3�L�؛��䞘U<Q�x,��	Q��d98��TJ�9�V�ֳ�Y�8
%d���	fČJ����JS�v[����kw}�st� e�'�	������w�24�8\*꩑���oV��?{S�jΟ���.��i��Y�;�R!CWй�tF����>�U$* �(e�������|��#���bgOf�	^N�C���kz���t�%�����m0y����_��b��;Z?�م2��{��d�c%��Y��d�vG�U��p@@d%GZ�D��-�g���ɷ�I�V�'k���Y����և�+��}����v��/z�P�����d��\|��l,�Zkmj�]����������p¶Uj�� -]v� C�7�;��!�
�`��^kT13z�c���E��|��٥s�A3�d����Ը̡6*�G
��^��DF��ԆDР�K��m�n��W1��C��˸���=��h�a��e�^��aP�&!�ު*7�t�[lV#�Q�� �?T�����R&��K�mw��ΰ;[��]���j�p���Q����
�\ה�1�mg_x�s��hj�b��2U�26y>���R�d����B��	W��I.�bqK�#�?�bpeѪ��c7b���7l��
�-����T�\h>!���W�P��=��#&G��.���z%�X���18�������˶�ڌ�3Z+�+v~U�!��6����`ʾ� D�D�%x�T�߽ [��B�v4�[���ӗ�=�ng;���h��	�֢�헛�F��ac�x��R"JRyy���T9T,[���&�z�/�W�0���w'����\'�ʜ����u��h��""��Ò��H�7L��e���3����Ac����,5b����94�p t#����@&Qk턆�|�O����8�i�����]���E\�fh#���}�EȔ[�xAOB�$��Vlә��P�2\#>bڠ���Z�[���&�����I���P]J\�\J�Q/�Gy�"R��l��w�����ۤ=Ms;�E�'sV�6�
31H����:���a���+i���*-&K�6�lS߲��a��R���D�v�n��!�6a[>R���q8d��7����ҍ�.��2��>
`���h�w3"�@f:�d)?�\~_w��Ejdy��~���L�͚�ؔ#)b�d)�o6���RB0#�(�Ym��0���Z�;�WOs����R,��y��\fM����Z׀��˿F�;��T���5"����{9��o,���V�Y��:F[X\�+��֯�Ae�̼��ؼ�^���-��g^���wa_�%Գ:���G�3(2i�! �Wjt��ӑh�Y������?x�G����k�]-�lz�����>rk�:�(}`#C� $Y~r�1�v�T%
�l9�+���i�Q�PwS��ū/��/�o�ڬ��֐�����O�?��h�p��Ǯ>�n��5��O_j�?���A���8H�գoi�|�uäw)�@e�)���r@���� u�'�Ƽ�(V|~�㊼ԄB��;Ѳ�z� G�{���:%w@��Mθv�p��+j�ݛt���d�̹�7�A�f$dR*�]��;F:�f+ 1�y/.Tb�P7�.��95�i��o6ԅ_֮�D��sh��Y,O�xW�n5Y3�C)��!�>h�Xc�Os�_hd���E��X=�hBͽ[��d�8�!���ه��ܶ-�f;b=�
	������y'�}8	��|.���>�y�����VDBSq�_DwmL»o���: ����)rW��uդ n��;���3��+�Z� �a��x�Sa���vku��s�V"#kB��p���V>�V�D�����3��R�c^}�O��-꺊��q_�`����b)/#@�yZvC�W4���~XY�y�������>\���[3v>� ���	�-���U�x�J��7#���(LrQ��Կi ]���2	"�ٚ��a��"\�d�����Y3q ��:���>��o@��V��	Ͽ�j�& G6���1��bRk��o�lG�J�{n�4a,�퓷
5~����iAS��1'�L5E��r�a^�i[�rp��|��U��kDyr��9ʾ�$�_��_D.[p�~�J�́?oe^:�L~Vf����(�����
�N��Ba��.�U��X�0;�ͺ��YT���ӿ"�r�����Gr#���y�(Ҙi�4Wsu��Ǌ{ V�s�;�QPRvw�:;Ŷ�-"�#>	R���eZ��O����d
�; k�D� ��D�N�,h̦QȭD�����5�I�#�3�|�=|Y~#9qM��,�T����D齗���x�l�>�d����^"��D��q��Ħ�(�6>|�
���jk�)K�Ө���y���#oZ��P�c���ƾ�3я�D=�f�_���NX�=�W�������#wq���K~|��?��m�C'6��8x��XJEF�ъ�~����\���o}tOݗ��.���W����\Y#!�-|�FഅhG�TU�I�h/��f�j
C�ĩ�r�{���M��=׺�W��~Q�zl��������@f��ЂS&�gx ivTa���6"����X;l�x�dW[l��8��wO6Зa|�7��9I"�M��t{����g���k\��Rd�S̓�H���p�¬���r���.v�Bl3x��;��k|S$��Y7?-�i֘=̍"�y調3��C_���c��dC�|Z���Vsޑ!�r��� �ζ�Ehܳ��
����� B��S�Iq7�S��u�!��\q���g͚m�D��0�k���i�'pQ�rŰ�[�p�#��^:F�=�lC�G��� ����U<���rN��c���'�Ҭ���A�����Kk���	p�D�пQ����k��h~�EVS�,��#�5���2��ԑ�l��{�#Q���입�<�Q���l
c���`�9�9��$Al/� @l^�_�.��aVY�W�	�������8��k���1�� 	}݀�{��,�W��)�^W���y>®�)��������5�eUg��:��oMm�u�{��b���e��Ȼ���+��.B�S���,B���H�o�&FܲDB�F��ͦ@I�Aރvl�괽<������j��0�|��� z�z1��bzw�թtf�ciX+G�	��]�T��Kڌ�Q��L��F���|�U*�n�3 G�s=.V����י-m���!�k�=8 �s��?����Z�$�}��⺒{]��Tm�6E���&
���T�ӒP�u���o�-��q �\@���7Jkr��L�3��6�`������D$�ϰ��c��}@���#�/��b�;�8r��F,E���gcѫ���LV'��Rj�'�����A%q�N�Q���W��{�גh��4�b.p�j�Ų+�dU��O��:z��"\5�E��-�=l���u�G3�,� 9�B�
�u����g;��}'k� -&�l�hn�h��1f,zg��&�iN|�A����B_"�-���x�Q�
� T�-�G7:KW�*�GLqz����:J���@�_~�t�r�R.�{=�b8
{5p���9./
�c�����P���S����<L)��Jw/���D����{�� Z�i�c_"H_{�*ݻ��T����t~wٵ�ϋt����n]����?�J�V�=�ڇ+�;EK��ǚ���4�Z��=�m��Dq1������:'�cxT��ä�����i|quA�Y�O�~Q�<��u�� ;b&�}mf�o����#���.g(e�}���U�o�Y�s�;�
�ť����<�����J���p7;.STӑ4%�G�2�wGdV�ol����4�R�v��B�1x�L-Z//	zv�d%������L�8�1��؞���[�s�Ht=[eI�����8�)�u���]n�����Xx���̸�}����=��x��_,ΰ�4�<�h6C�	��Qͨ�j����ٽ�aM�l�(#�c��[���ݞ��B��T�L�������p0@1d�Z[�9'; jZX��ሚ��B�wʂw�E�1$�����F_���ݱ���M�1��I�@�'��~�"~C�/��%��P��F�}: Ԯ_�_|鑪b�w�ӿ�u|(�WTuU��5�0K��ԲhG���� jhD�~'ZNtl \ ��z\�������;  %
m��s��B5T0�$��)��q�������Q�-qg	�@���� e�#<C,'�+m6N�黅�`�i�(��X��m�aٝ3�F,M�Ms��|���O;:5����Q�q��Q�;CQds�+n��o]��ȧ���e鹩v��wj蝒�>S�JGJ������;��)��B+s��e^���$����9�����"M�'[��]����q
q��^�}�-�a�����H�+ң
O� ������s
��;L�"v��v��Dhƣ�����I"U�)����;K�Ӟ��~����L��x�I�쫦N7|�"�;���l(��jM�?l������*�S���ZE�	O��D����V8�l�ÌQ��%�}j:#�AqM~R�q����d�Q��Α=.�n�Av;��#A��L܌���ÇKb�N��0�Z� Db�=pk��a{�}
��5O	�+��f�̎���R�?%`�K�tK���.'c�S�NEK��(�����M_�IG��[��K����2����uf�׻�!�,2��A�(�IY�Q��|0��X�u���	`�H|lg]�L��*W|F��6/��F�E�!���AS�+��i�H�بς����y�ыj!�>��`��!G��j�����6�0�,����;����%��0�ϫ�_�=�@����a���eɨ���,!�N���"l��%�
=>�����*ؐ�<\Y	������d)���'U�
kR�n|b7��.��l����t�Z�r�fKZF�BG�b��.�5�:y.0����!�W=Š�Bɵ�ߺd�¸6�۵~#�g��ɻ�V���ܭ{�Al��1�
ik�}�=�A[�g'�5���i�	�}��t�Ώ*�Pj�U�=hq�@
��ުF�xڒ�����0ce솢�'^���=|�vȝ�w��w��^��q)�h~ ���.V�J�f��L�:7�w�.�K�#USM���=����qFG���9ЧH����K�0��v�֋r �B��z^V���ddp��͡�M���󓔛UBB�J:�/�1u�KR�N�7s�8�+��d2�d� ��QZp�w؃ԙ�#�U�N��ǰ�tN��w@�Q������&q�;7��ڸ'g7 +�8{��t���E�	Km��L�q���dp)A��)2^��Zv����e���P~1������Cu�Q��~�g��?˲q�=�L���Q�C<�tS2�R�P���}Ф���`6�4_�`�震��F!���X6ɞ���s@�����;�̓��k�Q��k2�O��t!��kmMY�˿qF��d�*��^m@�����Ψ�(S#R�$�ş2�3�H��V"��iuoc�j���x��;�e=��+r��F�ʩ�[��Т3Pfm�o1����ֽ8��!A(�!y����7b��b2��&��D�x��,���������<�|����0� �ZY/7��xE�IA560����p_�FB��QIy	�ir:��ҢX�"#A�Й�����l�y d�㒫q��t�����ʲ����#륱棕����Ve<�����'Y�$A��	@�6��,�D�i��0�=�ЍD�^�@k��f�����(���]س�?�Y���+��L-�}�se>$����h�)&��׶f?��gE�R���df�֥m�I�R�3��`{m.I*c����(^)u�S,�|+����[��h	m^Z�~�N�@�s�m�02�e�>�!DjoK1M��j�A��@������`��IR�[���k0�G@���ə6�l���o�bQ��$�8��b�"�n��?���wp��W���!b��Q2��`��������"@B�/ §��0�Ѵ��M��E����Ma�o��iҏ+DS��`�Ka�Jv�پ�ܸj@��s5x!0꫔�L���U)���|	ŀh,�Y�Pφj�BMMT>J����}�������w��������1��5�;5�h`�LŐ�Zzg�Xf1�URU�j��Vu�im������$cNú.��+Z;V�:Kqj��r�ei.�%v���9�|����y �H�,DOm�^�rb��K[̰}�Q��IgE�,����{%s�k>�59B�9�����_y(|n�՗��36b�Zn��;ʹ镋�����|�%�ZF8���xT�8�N\����̾i3Fp=G������n<?p�I����p�����o��x,*��)�����p(<cp�M�x#YYrGD�r��kd�_/�"��j� �0CEZ�$%�iCZ$gj�h��{Uv����b,E��k,�+eJQ�χ
t�-+�g�$8M:0y�@�Y��K	�(/�rP
�� q�Q;����9���qۊ#��EP/�N��J�3:ݨ��dS ��¾�V�o����Y���Y�#�]���-ϓ���E#by�'t=.v!�J��j��.�Q��R!_u7�(�!j�X��7G�^��)�`��[
�H�b�S�f��o]S:�\�.�RWK��1Q�1�@�pH^V|{��0S�ـ�
�;M��O�i��T{��I���di$��~IT�l�PhM[&Pb>=r#*��PD4O��Cd���R���cj"Zh
H�60��[������5j|������6�c�O�@}2�b�����^)O�rB�le$�E�#�;'�����	$1�c��ɧ�h�״:� I�,cy�t̕�jђ؛��s��P���,�=��0��[�q��7��]�^q�C&�������B��������v�l�\�X�t��_%�܄(I��L�|�lM���?��h�3uG������V��P�+]o�>��r"��|ʻ*i��a��k�GM��P��M����	�� y!��l#0~V+- ��vJi~����:E���6��a���n4d�4���3���?�� (�����3�.�_k�7��*�nǣx�O����sz�zY�����Vʸ0�����ul�_��"�	�sZM�FȚ����Mƿ&�kG��o�8�G���"W�e�<���ۥ;��_�	��~`�a/~��'���$vY���
��} R:'��r����M֤��H@U�G"[F��.�Q��c=J���&vf4��h����<��t���m�,���,������t1�c�ܕ*�+r3y4ChZH�|�\�����Э��؁�-N�G&^�'n�;��ވ��2&��W�l�xrqr���@!������p�&�Uj�z��P);�|��F��kg3�d<L�"OgX���&��y	�}�m�W񮾩�k3���[���]�����������6�o2�GP��(��S��X��ا�L�����;+U�%W�ƨ�HnT���x$#�~Nj�՛�|"f���v�E�����FP���^��Cx+`V+�1�?Э%@��S��$<�����j:~�Of��A�`.m��JV�!��Ԇ����sp��+�,����o�.Y,��ʹ�0�i�M��\�]4��)�؆�F��ZDY�!Dם�W"�2��y�xcs7�;�쭶���R7���f�`�Gh�D|����s�[2B{=2���8a�z�=3�Cn�~���PS�D)w/�����3Z�B *{�p6/Aշ�A8��w�N��%��� 0��=���l]]h���-�P6)N�D��,��w>V���?��\|3��#�v�ŋPg}�ee�}1ҽ�&�F'/'8�/��;����'�{ك��!��I���&����p��a�&g�ݤ��7$������ۄ'̽/�e����{�8���Bo��id�K���8���e&�����"`M��:�*�Y����e�V@�#WX��w�|z�T�vy��8u�~e��H���wa(W�J�h$NVafGg���	��W��v ���I{���p��)f�Hdc�~�uV8I�600�e+���榌6@���u��*]�j� ��<��D�Q��OXfd��7�6_�I��p��p��V@үkT7��d��,���,���[q.~��= ��ed:[�a<#�Qd ��� MMI �[=��L����ps�r��,��,�k�JO�@�4�]��#brH��b����?1���W3��@{���@����:���PV.p�O��׽���$3l.��Q�ˉ؋�0�	L2��eu$�Ԏ	�=�G����KJ{	�m�}�^��ԥ�0L��-�a���%�4�ݜ5	Έ�kZ��e�0U�}|����nW|�ǡp��� ��{�s�/��w:��^�����w���Wgc�H����b1�Y=�D޲P�>���%Ok_wdg-�U��&ߧp���C@u�������ͼ���-,Z��ZͲ�{~g[7w�^o8 jxB����"�:S������;���aMy�:j���S��֑
0$�Z~���1���0���2��M��MO��h�S�D�9��P��Лh�@��e�jˀ)�N)L��z���d�<�Wjr��"{ݯ�,$݅e1b���f��>�|��K�լ� %F+��Z�S�����7�i�a[	��r���AsMc�Ms�_#��EՅ�e �XY��x�iK�����}�-�5�H�j������7�*b~��<ϯ]���<��$��tIz@�x�r�̜���a;�W���s�/� 5��:^�xҹ�Y	�óq}���g�c����&'���w��.���ét�A���p����\�(�Δ�߿-mGƾ���ʩ�i��]^����tU[M1̺��*�ZP��xM���Ӧ+�d8��M�G,��L��h��K�d�,:7��r��A3�ʹ3AtōR��8ǆ$Q��-L�N��~�t�Tŀ�ʞ��a�����+�����a�ҷMo�ݨ]��b�8�u,Ɯ 0��<���/<���K�5��JB�5 �X�	gs� X�����UV.ZN|�Z�4�x��x/��G�V=I���3Ϩ�'������<�S~�1�u��2r����!�)g"�U��S���Qt�����_ �[����
	/mP�ŀ���ǝ>��i1�s���.�[�lw���s�1,�=v��j��|g�l�B��/ګQ���m�AC^~,�o���O��w`R;pC5�ox:=��W���}�!M�Q]�^<���D�21���d9�k[�o:(Q�%���Cn�Z���E5$�F�؈j�IXAaZ�'�+{���_I�Hqq��Ti�{ $R�;�V��#S�x ��۴j㎺^�ʭ�J�K�ξk�j��h�JT��CI��HP���b���"�ꫩp+�˹*�V?=ګ�\m�w�u��,'�q,��*�� dxA���hL��K�b�`=�<Ft_���
�|[F�<�n��D,X�0L�Ó�AS�E�nĽ�~�P����+{6�wL7edw��[�O����8�ϓ�gzLX�@��`�<JC��,סz��$��5��9��2$kz�je-�]� Igdz�BF�J��:�Dᔘ�Q�*I4
Px4o��#�jj�qC��y�s�љ�M��L�OZؑ[�@�dڏ���[����HI��I0?�`4�G���| J���4�,aV�4�R�?�ei3�s��A1f��ʢ�����i2B����}|�X�r�#� ��.�Э�G��xo@���A���᎕@a�3"ʶ��V�7�N�ސ��O8}I�Ǯ&g=��]�*G��Q(�t�E(��U���U���G]l+�,����@"�<��V_����3�9t��q�ݜ(�mY�`ׯ��q��8��q�'�t�rAL<����B8������6�ӣ�RԑO&���+bK1WkD4�u<:7O��Dq�Q��؁�n��\��a5�6��V~ �m�Z�e�D3+����.���r4Ǎ�5s<������/������I��b�%������,�J'Zv��2��̀!H-����M��ǩ.JD�@F��R����/�K��\M9l��oJ�s���@@���o;!S��!V�:�=����7Eg���4E�$IiL=��ц�S�Px�VQ�5���hV$�����&�{�0�������b���糦�'�"}�ڿ��Fq5�L�硦�����4�p	���∿n�H���l��V(���:����S%N5���C]e���wX���XZq�_��?hx�<��G�����:����lj��7��Z��ۃrZ�b/r�����4ڸ��.s�1C��w�D9�`:��$;�S/��T�QX�qP.���I���DT�f�m�6hU6y�0V0�>H>�d͸���+����u���ЇL��%���� ��i��>%j�[��@ l�m�r��
$	wy9h9�iE5u����G�PrZ���
����mT�wLT�C	���:��(��#��`���f6�����n��hD�X�v��)c�ǻ����V�r9}Xl�~E��uR���.0�T�v�wu3�r]�
-�>(863	��4�+��<�6j�F����@;����w��'�'�jRF��g1)n�fԛW�P�sŵidn2����9K�k~V-dd�1��0�	���Sj�/���?�g�@�ҽ�ωH�䉅� u����3L[h촯xtؙ��pB��C�#/�}+`�G�dI�xm��\qzo�8�1I�Fr/��2����;����i1�wc H!Z\����$�"S$���.D��MF�s��'���.R�[�14�3�2���vC�����m}O(�YO2� .�M��Y�J5���b��B���� "<x�3�~*����#m�;�-G+U��W�� ���&A�����=58�t�S-�F�0�����W�R�GM8������}C�0d�&���W[W����xz������d�9p/75Rɬ	зg�j%`�Dm0�(u�t@�;¼������Nx������l2�٢F���C�\��JhP�ζ�&*�fד�n����a�[|�-��R�Z-Yh7��ͥF]κ�v�oP��s~����=:]�Ӏ�
��,P��$��'�_���Œ��rcX�zS�|�i~f�r���|1YE��t
Q8��mӴ�� �E��!4�&ʫd�ob>��@:ǧ���=�㳁i_v���_���[��!�[=��#�26rI���.K�҉���*���WT�[��=.A��AA�u�?�#�>TB�e� �����<���$