��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъQ`/�P7L�*v!�x|k�܄Cs=ŵ�4n��mJ�W��Ű�9�Y����1�����Q��� ���5���/ 帏��}(���.CȖ{�)����l	C�����qt�ݯ����ȟnWf-֊��˾�X~��q�Ҋ���Y� >e�1�ɝ�	<��E*u_�@�ى��|���
`�>�ur
�(�>��{����k����1'�Ox8P���,z��{dO�l˃�Q��������v��8�Wx�+]l$���7�!i�>�on0��h#^���`��n�!�G k�q FVw�|L�~`�(L�
�P~c��l�����G���b�xr9�e�*�@��
[�����U0h�vmi��~5Gߧ�5�"�U���e
�;��3���FF�dY���Y�GbB����!�)	��b����N�a4��ɷ�m<#� �����D�Ϯrv+�@����o�]*B��N�ǘ�S5����8K�[�f���@�r�� �5S�̇�&��`1Ҵw\@�L#�؍���(槈������A���IZ���]vg�U�~�q֧>#�u��?_��i��3�TGc�j��"ؙF�T	M�Z���ԎE�-m��m���.��e��*�<�ПJ������j�`�[hgI$�:*���T�1ߗ�r/�O9��Zf��z��t;��V2}t���u��FwxZe	"�h��.'�]�aI��n�F��J6�͡,}�Ya"��N�_��!t����R�#Sc�v/&��[R����_����v���7���sTQM�R��Kq/0WCa;�FmEjG����q��L��B=b��٨�NHK�x�{#�L�<#�Y�r�w�{ڱLٯ������TX.Be�r�}6�aÄ6�	^��o�`� &>��|�k@h�0"��%�aM��I? m�����C]�KV:�^R�ޥ�s��c�"9�;�܅����R�f��~�w��^ꀥFό�V&��
\^���:�<��8W8�k'�
�<���<\������@��D�VԘ* �7�Ƨ��
V�'q���$Z��51v��	76J��E��[����.�s߮�Y������'H��3�mr�NY$�I�geݱ�&�iƭ�Kt�� ��U'�we�6�K�|���*i2����2	�^�p��������Bu����s�S��HG\�;ٵD����h����hC�!�>β�{�L�(�-5�o�/k�n��H���Ap���"�%K^��s@E���R�.���u�B,xlZ|���&�)FnwU��`��nW����n�b:�M��l@e���N���9��c��Bc�M�_�e�^�ԏ��m�&�t��N���y �﫷R�њ��r��7��5��:� �w���%W������KJ?-8�B���:׭�K=9�HӋ�/|}�r��Q�\y{:���7��dYZ1T���O�J�H�鳑���Gp���+#kA7�	� e�����`P8඄1�����p;��^�dKe�{�B����Km�����yc�K�H�Bݔ�
��-�"�O�ѫ 3jQ*S7,�u�4�04�9���i[�бr�t��$ {B�Rj�>�s	I��{�c�;*��-Iq�SPJz���;�O*�;p��$n�^"��\v\(���
`��{昇��L#�<~�zj�#7NӪ��/u��/��2��V�7Y��m�;�UX�Rއⶮ8��sj�������J��G�10o��ϋ=lR{�
����$.|�b�$2޶�	T1�FP����<��^���0	q�lEZ�b t/df��J�:0����'�rZx~���pmyo�l>{8�I�F����P�{c��
�ݔ��n�p�ov��+>�r�%B��(j����J���$��:�и��#$$��>:�غ]%��aR� \����
~�ߡ<.��$7f�u�=+@��@t	D�L%�����1��#B�?�� ?���CA+��U����!T_��k�/!�5X+�cC��ED�t��� ��S�U�:x���5�f�k[�Ol�����uu����7��F=��.���|���w�9��6�J����Qǯ�x�QG��9�R�a�����ԹdNj���cO�IC�	�d���A�*>��ϛm��H��VO�Y�8'�b:U�ޙ�>0�r���(;%�#�@x���~��}wE�R����������+=��F\zK��z�a0DU�W��6ڊ9e(�&�揣��[5���;^�d�Q���["�@�E�B��X��2������m���a�c����.��vZ��i�W�Q*�@���Tܺ8{V��n���٫�����T����{��Z!ә���C��/�0I>�wng'��M��#b�Q��f� ���e�.��+k��:�_�è�)%>˕1��g�\��Rg�ݮ�5�֖,CY,R��9�3�	.��e�~P1)ʾ�O�A2G�5�����Z�2�&�@����N�K�Jn�o�^WC,��o��7偸�������R����zTՑ��Ć�f"�1�����MG�M\����8����=ke��c$� ���0=��� s�d��*��-���Y��'��q�屷���(2Yz�J�Cz�Dq����@�j�͛�?n�j���U�p?9�d�FUo1�|��L$�^����A0�tZ�i�}żbBA�j��C���9(���fΧaϴ�e�p���S�C�ڟq�������}"��߾�߈��)���cq����/l8g��o���L$4s9���t}�r>���[�S��ֵ4ff8A@���[9"����Z�����"ҜtQ��X�Y�ݑ!�{^Pj%J��u�f�r�eǁja�'(1j�ϩ��(�y�P?���C�<XK����ce�GzK�4�%;MK>`�9�N.�E�D�����l�B� y9������C�����0_�3��'A���\�J��l�Q�z׌��jo�F ���W/�͗}h��N|���@��Fl��͆�I�&�����D�$���\mSh���B\JH��d)&�����d��$�m�"�\k��:_�T4�8ztM��Q霰�_��ov�m�pn�='��K��0�*�9��)JRdx�>c-�y�}?rB'�bK�5� �Z��/Q���C�%�濝΢�Ίݬ������.��7A��e�k�0�W�L�ՠFy�g���1a����'
׺��+P�z��_=+)~�'̳��M#��G[k�9���7f�~3H��M)���V�W�S��&�טt��»<jf|��nC\e+���`�mɕO����?�.J]��y�.yؐ�S���?�������R.'��C�-I����[[��Q�obد������)+�d���i��\a��*(Z�ʝV�0N�/"���e�
eُJ7�T��~��r0��:`����g��J�`z�HO�q�ޏ�K\��1�9�NE^�~Aa�]�y;�F���Tq�6H<����M3�'�~�)�R��3�fq�y$�)����uՋ�ʋa�� V�9P�N�!�@ /��e�/5D��g������S̈6ܷ��r��;���m:�!Ex�qݎ�_���T�4�Y�h�y0j8�v�
b�tY1v��m�5�	��0�?��s���,.�Һ��'\�=�k#���C�L����%���oi�8�.���fm}��C���2M-����mdI��P���Ip��T�lte���Bg¨��^��3`cj���/L�in��S��ku��Ƥ����d�73��Zb#� ae��3�2od臶�s29߸vڣ���-�CG��o�N���߱�y�ѻ�o�d�03P6a��Q��� u�X������OE�ݐ���X�S`�p�@����꧋�ez�(x�R-�h�(l�x��4��W�N7:�O�γ��(��r��Ϝ����M��_d��գS�FͿ-�4�w���)
l�n:]���	�vckwB��4v��d����n��*�/ZX�]������M#�P�he��y�t�ݪ~�;0��b}�4_��`T.�YlIˎ�$T�h�#U��]����v���t����m��-��by'h+1۷��6�p�h�h)T�3�wڥԧc���5�R��Z��Kձ�8t��s���̞6!���JY�xXK��{��ű�N��'�/�*@^Le�|;�E��&\���f����Y�3#ڔ�=$��/%�OA���"\��s5��5�#��V��!�ȥC����5\?|7��t��(���p�E��O,[��&[Ҙa�of�v��.�T���框ۼ��p>:�pr�P�"85�ژ���f ׮sE���T?m�R��ڿ���e�i�]�'X�:��CL�l�B��)PC0�V�I��em/3	��8�ۼ��UN�Y���~CQz�ܭ؏�Ȑ.u`;�f����Ձ"�|�ŗc���6�=ZS�Hy)��Z7�ɶQ�R��zŃK�XKH\69PO�`��_���`�ږ����:&6��3_�xJѰ�8��� ��h��1���p��H�⑨��G4Kߙ�F�0��xɦ���_���c툷Ud}�qJ]V}R$�H\���fM��K���k2:���p>��_t������4&+Ç����&5y�<�L�*��J(�п�O��T�@逧��md��5�Rn�t��1=�~�L[Fº��WU	����u����\�IU�\R�Q$+���p����M�;Za`?�)�inU8�2.QP���{��(�����Y�|m�o�@���q�8X���C���@�|F+h��G1�V��q)o�Ie 6��{�LV���ԽMD:�0�S�S�2�e�%Vq2�	pzl�y)�c�8n!~ӿ��m��v�?�X�U4�q�n���e)�$8n�WG)n��>�r�c,�4l�6Flm��`������\��|j,���t��(���Y��@�E34,Chs;H����N�0�]�!C�O�%�lS�3PK��d�1��Kek��ZN�*t�z\�TJ
��u��_z-�!�
{>2�M�4�mׂ��p؉�/&w��Lh�3� �� ��3��1���-ō8�S�����*�J��:�H����fԋ���o=a�S�湩��:l��y�޴���Z����l"��a�K�MQ�b.]r�2�Y�J����QrmŉuX����xA�]��z�c��Sa�H��ޑƱt��������$3��9��MΗ��Mf"-��Bo��^�c!������.v	_�1���� e ��}�'ƻ5��s�&,��TdB-��1�:1X�����]Tr�ҧ��4���a��I2�/��nK��3\�I���� [�{�(��Ѧ#�9�xԵt�F��`��D�����/Z�KΊµ���S A6<xoԥ�厯v��VB����<�x�4 K��|q���l0��"�qd�4Fm�͝��@]��)(����6Li��_ByM3��J�7�!�@�_��c�0m���/��c����y�[��\CH)��(QSE����Ը�.�
$ æ�x(S�-:TRC���#Z
� �� p�դ�R8���P!h�^p����K�킢,
�T�3��.c���B�"�?S��:�b�@D/`�&N�l�~p4�%'86�jSY��w���!�Cj�������5�ĈNvX�D�;��	�A�66n=T�Y:}z==��f,�h��<��P���R��\a�ʀ�������,�0ūW�9�7��{g����Q�����%g�0�)]0 �0��~c�]���g��D�ۍ��p�ץ����LHe�0B&_�`�pZ"�`�WC��[{{�"ݱc���?aF�"��T?��L/u:�mD���Ύ��o��!F2� ���ܼ�}���4���N�-~c"ID)|�WZg~x��盒��%�vɩ޵+���4)>]����_J�&0 ��W�V5�R���Ʀa)&�W�2 �]�X�Q���&�T�{�̃�['�K�HÙ6�����\�4��x���8�� ���'('�z�'HT����/_�I�΄ϝ4��+��ڀ
�ii�eWL8��e>�4�P�hYn���e�K�ղ�r(��h�e�9��Q]<+գ$���=vz)MQ�*2y�d�c��л��֟�-���&U#t�.3�����C�Gm�H[������g!��\�EM���P4����稍шRnDW8W�`I.��u�=~-��c����~D�l��y��S`O�J�8��%������q厔i��
|s�����gʒz�*�٪�������&0 7���&xC�7�f�	� 2�1xkK��LXX�-n�*��YNm�B��Vټsӏ��غC�SC�u����X����Hc5Z�AF4�|��L��Q'�پc��j>���q�'"Oj���~2�	��k��nS��~�l���4N�����c�M϶oJ�.�9�jW�z �/�HQJ	1i
�Ko�Ӆ��X�By-+$����AR��S�fǨ��u�Ұ��^M}��_�r�p���~A�7v��'��f�@�O ��͔��)U��r9��]�ŀ��w��Z�+��S�X(;!s�6�9t�'M1#򸎜������S���=�X��N{�T+G�G�˱�ǒN!�o��l�ng�����>�k�ZSߖ+����@�]!�T0 ���6��<��iP�������y���b��-��#��$�B�n�ܪ.9��'d��)b=�ԗ�Wj�k+,��u��C��ذ�%)ۨ%EN[q�Yw���ʶ��2h|>����nW��2��5L$��cu��?��Ґ�����3�F�r/M3GJ˙�a�އ����$ ?�y;LQ��H�7�ǝm�B�\�:����b�j�Q;u�h�B�Y'M���ɦ$T�ՙ�VzK�K~�_V~���d�{Zū��;��vB6��
��r%^����T�m���N_��h�a�B]�u�*N*L����H =G�H�R�7˗#&�AC���8Ŧ�����/9Ks�+��6��� ��9!ͥ�'.I����^�7���YC��/�	����v�ʔe�A���Q���_7��3h�����n���?�^ކE�̯�-���Ƒ��Y��Ӵ�����8sV9�z�/6dy9�P�t{��x �(CF:��S~/�o |�U.u���}��Ңt���.g�z��&��O�n��a���J��X�7"ɳ��tʼ�9�3�]�^l���@/��@�`j$T��3n�`��0��֡g�1oQN�.�Ib�[Їl�&6kD��F?k���8���7sp+�'q4w�Oל^��x��SΩo�q��}هp������n6��&U�Zd�	=���:�K�`O�-�!�&�\�$����U����{����~�+>�DL7gT�vJ��]7�G�N�����x��I��P���Rq4Rꆾ?0&��{}�����}q�R�-_s�T ��A�g����~�e��������H�4`�:�TJ�\��{�}�Fxls�^\���Pj��|r��5T �\�v��4��z��H�+s���ʊ��"!�c{��ư�����.C�].��̅���p4�G���]�����ЈI��f:A�4����0���j�'��U�]���D���&�0�����@Q�G4ǃ�^1��L���j}��`��$��U����O��ϡ��"��[��l� �1�Zü@X89������>�kC=��`8��z�?�>������=K�M3� �;��Ϸ~i��X�e���çV{���}��˷�3� (�H)�E�1)p/�}H$�\$���E:����Y8�jRy�b)�a��cDA�=@�Na��)/��t:��ܧ"��
�<��Xд��f0���Y�A��s&��)�h�VP_^?��S�%���%5V�
`�O���X+�������F�. a+������`�����X
�ׯ<&��b�i�9�/�0�O,ŭ��Z����)<Bw�y�W�7�.L�XZM�*"�1�=A��L�h�|AJK���̛ut�9���繭^��,�2,U��t#;U�f#D���;Oa㪒��*��V�[���@��ςG���4��G��*P��D�{���Bp���u�$2l���M��]�]۳�`��e� �7�w��C7�'T�.o��-�N�f'��
������YaI����.5N)�x9�.��~h�^�7s��NB�����ר��:>K�!�����%�x�wg��7��X�ȧ9&�*я 犽��e����y�5���//,��~GS�� ���M�l d?h�"�S�B��x,)��Ad�h�Z���B�Q���0x��n4U�Aܒ9q�𵧌S��Q�s/�)�.��_� k�$�~��$�{F���7�Ec���NNIE��qm�H�����<1��I��L�n �7L�ݺ*�>���8'�O���k@�hʠ�^W�����2���8���˨ ;����R�`5�PN�q����S�y�j�p�Ic��sw�h��b�%;�N�8��!@B�/�^�l�W
�]ٔi��g�������neg�����&B��w���ޒ�Ƭ�Y嬺����������q�$�z��bXq�K���k�Bon�p!b�l4�\�I�`�9Y���.o=��z�>�2g�V�=Y��>�s�z�ֹ|���������܉��C8p:	��oE�2���^i��z}�����l�>#�ݔ��J�Mv�ZX���q��2����$�0G�ϡ�%����kh�UF�#�ٰ��טSƷ}�8�];�R���h!���d��e��J�.Sp�gX�m�2�GdS82o����}lRv{�qp2��)<��rC�!�X��b)풝�Up�����p�<[dH�Zh>	k%āO����G2���b�eW8�
���ľ��J\{u>[���{�7�a�<3:.F��� z2m+F��o��[})(w$!L�v-&���үӃ���I�#�h����{D�CʙwuX�	�}�r���쏽C6��itBxS̰X�,x�U.^۽���|�
Q�����2-`�0ŝ��aٝk��3J�o,.�����8��1���j{��RH��`��B�Wm0ӪQ�ǲ�kw�����iU�ԙ��]5�cF3rh+A����
Y,��UÛ�;�f����ϧ+vU$g�"N��3^DM���d�/�@��5�ystY���+�l�[78oR�\�V�Xp�k ��>�����q��I֒�Og��'�h�<3&`��ْL�������-�л�)f!�Y.�Q�Fg���F�F���~����"�T^?������v���_Od�%ɢ���=�6�RB��r�SQ���O��P9�n�r�W�wVw`)�z[�R�e��8Z����y_ �V�cg��cc�w����#�1k���'ŌY����z�n,�{@��vq|~N�k�%��@m�� x�1��S)��������|�*.���qN{��ʙ�2kT24�F�{�vC�I)�vF���m�p�]���A��ri��6×km"Bߍ�����!���qS�5i4���;x�ķ_�\+3JĆ�L�����p��)Vz��`S�o�J|�FF�yh��/I�f�^�hq@ٻF���'���띊�)"�A9'���Ѓ�*q`ݟ3�;;�� �h�l���!�`�8�2�)�lXx�_��qB���ZVz�cXq��L�Vٲ|��W��5�N�� ���u��/���E����Ņ�p������R<��Σ'�[��D����aj�_�6\�~�S���Zi�C5�C|/�.��됼�U7�x$�cƹ㊔]�E/�j��=S�MɏtEY<6*'��ЕB�XI״)��:�.(Z��H�����M��[��^����6hK����\�Ŀ���;��k����<i���w�\����aqRC��������a����v�)�H��W=ÿO;�v_:�7_s+鐑�/0���7<qΌa���DA�0�w�{�$�c�T��*����ed�j�3��cz�Kq�����*�V~�߾�,��n��+��=�T�3R6�i,n������vꩫ�
�a���8�����υ����j)����j#���4��L���n{�߄F=���$L���"@�y>l������|Z��_��p�ذY�������r��v-nncm��8ʲ{�s΢D��nQ�OFy̒P�����,�7"�6'K\�^LX2�5ļ������=��:��楤��1u4xi��.��ad;xŤux:�.@�w]�U���O���wYLhy��;�O1�9?7�N�9�;���~z�H�F��j����|�;ܺ�dڴ}���j5�tGz�c%t��v��a;�]�7�I�xih ���&D����h�qOi�����qr�?5��x�oȅ��¤cD����F�_^P��[��'W�? �:�Gd������.ͣ�\N��(�Y/���^�^)4��������܍����`^J�2k���Ņc�\�P�kUc��Z������� �s�t[%�F�񨆆���y����^�8ne��w-��|c������i��
y.���y��6A7�o��{�|b(w�x�P��5��Gvj�ር����S��*��qⳂ�]r��A��%��kl�½�r�|���Ķq_-gB(�l<g����A���8ke�/Q��F=H�q?g�
^m�ŋ�x�_&Ưy6�)���#<m/^��'wtCR�6�x���:����2`�e�n8׎����i�_�-�
��
+�ל��w#��e1�|�+L���Ԣ	ű���I3LT:�Y��Rxqp���������V����oi��������eE֖w��ޏ���e�Z��@��F+hr����K*�*g�]����~j�S�K϶�4+�"�Q�����[�q��#�����o��2�kP�5S���U
DUP�y�d�����g��`���J-V�~*�{�Z�+6Y顝(�Y/f�wc�A� ��Ҿn��q�:�w*�j�[�y�p:d=Ʉ�Q��!���Ȣ�ߍ��5�	�d���G���
y||(u�ȝ]��
K��.zj�:b������Vf�"RU1OX�O�^ �W�2\Ò܅�W�;1�z|pV�ﴼ��ywgQ�\�/�z�ݲ�4�4�
��)d�Fɾ�co�S����zT��:;h���S�YTm%FH�إ#�`�J� �)�����R�����vM_���z$%��y7Ub�^��rԥ҆�����>:Ƅ	��)�4	�h���	���
R�&���Ԫg�8�u/z��A��m����6P����u����OjQCJxr6�O}�G�9ٟ�S��N���B=A�ߔ<^��Րsp�K�I$����{P���2a��Q��6 �!���j��妃Y:ʍ�v����ͺG$���2�E �L"?����: _�F����O@�{���v�S���N͝n.�;��Q�L"�Ŭ@��X��[����q餹e���xBM�"$��{���`��Z6�@��ӥ��>x��o�"�7_43&M��3���)R->(X���s�Ơ�l�1����:
1y2T�z����5��<̛�V�ws7�u��ѿ��%�,�uޢBx�y�+ѷE����اJf�`!D��M�Zl�J���6��X�Ԓ�'��~bqp�.���2|E��%u�W��������&�v� ��Y��kH�[�҇�Z8\�iJ�zK�eν��:�B'�|�`��#i��d3hz�Tv���~HL}�{'< �r��PL��	�/�l'im{/ �рO
X�/�u� &�7�k�Aqu�`A$��R�9W�r`�D�Q���}�g�X�L�E��=�q��SP�jCC�$��G+,8���3���Q��0w�s�y ���9�W*��J�Y1��̷�!ٜG������Ѥu��U�T��/�6ƍ��A0�]h�JX�N\>o�[��M�M�*`�b �{�����M�ph���M�47P�}�z��_���<9�22Z��D�Ҡ�=�܈l�6��wI�(�<#� 7\��1���������ka�.�!���-6��$��F-U��T�k8/���)��+_]>�R�=�vR~Q���K&ॱ���m�Ho�z������&�*9b��aZC��|C��
[q�b�S��1G��zmN�WR�X���p��-0XQ��0�N�ݦm�_.p� 6,��DB�X�\)�V8�a/Db����C?l[���&����k���'�(��B���NB������(�j��1�#ɣ��:�f��6�1��@�(������`K���_��N��|f�zIf�+D��Nj:F!Şl�ɮrF�C7����̷FAs�X�2�d��f�ښ3�#�6!`�8SܻV~la�|.-����k`m��|�қ�P���y+ĵ<���Xf��nο�+���
���P�!A�9������g��ǐ������%��jx��d��ZG\'Ż�R��z�^W�5��X����r��dQ��Kw�ٓ���_�y�ww,t�ؠ�^���9��{:]z���.w+H�rч;�_���=���˔�ʣ�����;��)�ɣ����+bDnkNV �t��6���s
e4�v#%���7����9�ꦊ ��B���lj�������P�:�Hb܋�-��%�UJ��KY�8�'��r~ܥ �L)�_&8����jM��T-$/��᧛k��ۗ�Q�h���Τ��s�^_�L<G
wP�������p�t��t&)_�w����TXw1˳���~gC�hO�>.��<�p4�!'65��K[���β�9�V]�rgp�=s'���S���YT,������4a��"���9W�֎�9���0mR�y��_ϳ����4��ui�p�]���g��h�%U�i���ѡ�-������:�'*Z��J	�����eu��e7��N\��T)ξW�̅�N����XE+����O0f��f�D�� ���+�\.L�O���V��|58�yTP�C� �8�]��"���fz���'�t�U�o���M^=D0�3c����Ԛ���=63t�l���������"*���j��m��;������I�Kdt��$X�F����|�v��ڲ#��d��9�t_2�K�׵��'�|�.�c,YB��{D]�U33��%f�Q�Fô����w:Fv���a�J(Z�YP���3����Qͮ�,U��|��R�Һ!�T1���P%��ر�I���,�GL-s�νC%�n=��*�j
kc��;��@���k�z��W&�������o�McD�"|��X�dn��M<���?ѧM���'�y���PQ˾[�I@�D��j���	��������V��Ô	��0�b����!߳���q��R6 �~��!X�Q(݅䙾�N�_'Fˍ�֛���w�4'~��7IpNT&+Rz��D���25�`���Jv��pҔH�0|[�5`Ji�J�]9��X��+{4���0�\�+�z��/��vH8��	A���?��F�,���n��T|��Gez��Υ슌�|��]���[N*�����E��6�q��h�cW��:\`it����s�,��t4h�P�� އ��f9ԧB�c1���xد2ŷ�1��_bd�/���e_?%���޹�Œ4����'�q���$zG#�ƥ/��H%����@'W��"�<��P?��N�U�UZ�'��i��
�!C��3?�Ɨj���
�8f-(I��m���3P1�(�2�[t�ł��O�b��-d?V8�Q�Z3]�������;��A�Bݬbq]���];���B��2�@(�����Y!Xv�*�^�$�z+Q̓����e��V������ �O����ӯ��1Qǳ�ܛ�ܳ�n��1e��	��Q�[�gI��ݢI�gq}C�y�_�l@\��I�z�Oa��75VH1~u�[њԸ�Y��6'��P����Y��dl����{��$ �J*�ў�59�ox�ӕ��7:6�x���.�Fq���q�-Q�!S�Y�#O7�XA��)cj�ƼK� ���'_�j6& pʆ�����4����xR����7�A�7�Q�G�ߔ藮��\w��09�E��!������6긁����'pTN���!Ƹ��.� � v�V'�#,vY��e4�^���5��ZZ���6ǳv�Rk�Ay���/�c���e�IIH�7Ӡ�G]to7y���<1PCA��2��R���{�J(M��6Ez?EHh"���G ��!����&�l,�'̇��R��p#H~�$������6]�o��gK�~�%t`^O��WY�C*�=&~�@*��e~pO��=��26����/��rwCY%�����S2��@1>������lH�c������,�ŰH��<Mx,2�=3�1�Ge���Е<	v���k��21��IdxRŢz)�a���7�X;�`�V�����)}�I���� ��p��Y8���"6 bO�A�W��E�-θ��Ә�h$#��-�/b�����;@j�G����g�l�{���1�ٶ�֪��PlO���s��`���Ֆ>t�W*'c'�"���HFȹv�?1Bޝ�c�"���������%�@��ч'�n�<�YV��>;sm���c�n��_t��r��_8_����bv˺�]�˗k�^�R;�,hJf�K!���-�r���^�n�4�wAӿ�.n�l!�ks�@V&���]���-��P����p�X���,e"9M!z������B���G���z�1�.}q�����aUp]����0�p��0r�`���; ����~�|����f'�ӽ�Ց:$�U�ý>Ú��O5�Ζ4�b����%��i��<eR��`-N�a�pAK�~ښpUaa���������&�<�;�Bx0Y�<��f�C��o�<!�mi��&�&�^�s�vĘ��o�zC����Fn[U��	啣���W��'�ӭK[�bs2R��2yi�&8*��^x�]㋡�ےUD0ꈣP�	��R�Ɉ�ZwO2�Gaȅ:�1��h�����<n��J,�<mi�,��D��y��k�Z��8,�C��	nާ-�dM�]L��x���B�UV�%��]��ǯ�P�F�
�ͤo0��m���m��Z^ʄ�5ʮ]�;�Z��X���"��2Iq퇌�Y�9Δ���w��ٛ�wYX��XoH��O�z�uB�<M�*Q����MD`��+ z�i���[[Ib�ُ�2I T�V�k����F�`��xE���S.�����c�yru��ƣMg��&HWw�=��t� l�](P���P���I��(o!3����S���_��̔!Iޫ�D�:��I,;'zf=�02��N���0��i�Gw�1m�3k�+�Z�����|+��:Sn��ٻp��*�����$n�J��`�b�ܓ#dq�H�Ҧ�C��`]�!Ʋk���{%y�L���63����I�2�O+k�hr�vAou�ȳ��jv�G�o��[8�m��OrW5ƣ;l�rf)VPJtx���7��Y�V�RL%�K}-�΂ ���	@��Q5]X�&XI���j�����	L�/T��� Nm����S��c����A������9�3�H�����
��/���s��t���V7����ز�f��>�|~N	d0r*�[l�T�C��BKґ�&�4��퐃�~X���]�0����?/���3I;np�<#%�*�$�%$E�)���@0�#S�w�+D)U�q�@����~r�j-s%�p�2���ɷ�S��y�ޢ��%VƶfV�wA�E\9F8�_�)�Z�Ƥ�E��ȑ���A�R��o�OKj-�k����M�?�\M
	�ȏRر��<���ao��*���쎏�2�=	)�e�!�����q��T��}�?=ۓg���A�Nv����ޔ�"�r�S�4s1ǾC��ԋOY���μ�F�7� EF��%���8O14G<�Hn¶G;��Iؐ�$�������S��3��{��i8�D�25�g	��b�B�~V~q���Y�C�X�����+�3H�g��>��F���<.�U>o<��"���D��M��(AN��9E�^���l]�SA��2�_g5F�o�#�A�vE�t�;�O������<d,aܛ����$E�S���8T�v��/�_F�I���J;�嶩P��\�p��t��@��I�Q�������H�c�e�ճ��h:<)0$��d��	���U׆>��F	�������'�SNW��L�L�HEQ����'Y���y��s�2�PM^7xs\����N\o���JE��$��
_=ŷ��Ԁ�l���eX�X�ߐ�eNj2�O�6������-Jvc��rO��<̆b��zj%���M���U�x0Ƙ�c��r`+Ю.Tj�+&S�VU�^��>*�T�k	�T[����+��A�梆�=����j99d]�ox3���yx�(rGK���'#�:�"�u|G<�ች�ƒ���V^�KVZ�o����L��H�p�ol��ć�XQ||Nt��@ͅ�����;��H]iQCU�^yG��u���e��`B@��|�ƥT��/+"bVZ�w"��%~oE��A���W1��2���RP����OMJ���lR�J���8���xY��?t�/�+�0������p?f*�
��QcS��:J���z�O��{?�at���,3�;�^�*6N�ήq���H�b�Y���(�+�$Ky�X�LW3�~�i�E�\b2��_��V���"?�q���O&�|H���B/H�!�۟��`󱡥nt~�>0�#�|�/�p5[� �<oJ'����[�:�PD�T>$us���D�F�����;yb|��RT����!z���$�O"Ӂ��u��[��]�En7�Ov�1�E�JF(�
����9X� ��3!����<h%�ݫ�&�D�	�'����B�Cɸv
�X�?��Fd�u��{�@�Z���Z4a�z�.?s cPv|���}k1w����X�A �3����.��ur�mL��@ ����8�� Y��N8{��^ӑOPe�k_򀶲9碇=�ƾg��f��0/�C|.�]Bj\��Sg���Y�/�g��o()oX<�	Vv��%����/�W��#��.t�XŐ [�;�T!]��"�u���&�*O���~�b~2})���ͳ��[@w����و�jNM$	X��_�iJp%Hϕ{�����SztQF�S��z8�D+h��"ⶹ͂B��pe�`tK��D|gq�,kM�<} �Һ�Ӱ�	��Z��:�	i59hEy�;�31�$������,��k��M�ۉ84/�ȡ�,�b!����Ak���O���詧��5�bp1����D�|G�9�X� '��5x�� V�w�ϊ���ȈҜ�b/�
��w���h'U$Ӏji^�#>� ����g��>v������0�u�H�р�;<���@6�U��x����|3w75�-��^�BFÝ��`�6\�U�m�|К���דC,��<^���\ 9���1��s�!�{L-�vy��A"��f�0iܡ����M��܁��f��R�)��v��J�Ժ�7ɭВ�v���������pG��1��<�Es ��Zb�sY�
���a�:G�E�ꆳ3~`�/W�.��t�e/2�Zbn�*%o�  ]�w�A��S<+]��+x$�Y�_���n�Ƞw���xu����92��R�`̸K������t�^q��e�����/TcrnԪ#�Id{�_�?��H�����DIcr:iyq��yMˬ�|�َ����D �"��B^�v���Nb����h�Xޢ�ϒ�N z/n�Æc	�T�<�]�is~{"�1��O����MJu��#w�B�#��1߰�k��:�2�\��͇�w B��c#�,��)s(�]����Fg2�֞UQ
��_��T�}��wt���mH�c�3N(�-�|�%�ğ�a�D�w����o�}l�M g�5v���ٰ�Pj�E[w�bf��M���Mރŏ@���������1�Pdo�����v�n�RΟ�4�ft���w.� ���H�!Q�mZ��E����޽ꚰ9�a�7d���J�	�E1h����I,o�����w�2�sH�#�6�8����<��$FwZ%ɏ"�I���~N��L��< h����Vi.�vSٗ����ʞj�}�g4�/�c7^fo����<���y�'���N�����E�r~��"	� 2FKp]�vw«����>��v�r����o�l��`H�m8O0�q�c�7NZ�,m'�$:>k^��i-|fҎ�&�|S�p
Aw���cR͍#����~_�&�ME���5�M\�R���/�m]��`	�d�3y�ta�h��B�g��85����#�}r��B=�Z��6�C���%��@1�ٰ�4|+~&a���V���Ǭ��\�l��rbL�|�����k�J4�*���&���7�D{r�'m�5J�և�����nFWt��#	����X|�Ψ[@�H� ����LL�p߰/���B��$������8e٦�x�'�#q۽���n���y���ϓ�T��S�,�[�A�ҏ>�Uy���)!��sq���X����ʠY)a8<Tg��O�m�Ӈ6u��	J���S�2\5A_��\Y<v 6U]�W��:p����T�#�M�5:^Bq�y8pE%�/sR�;��$��_о1O;ј�
�,-o�:��G�9�k>��6C1�u \q�g�h�����U�6���8�g"��c�m�6��Jm��~_�`�F���F�٘�O�n��{�@�f��I��@Zb�Y_��򁩾�q{m����@�K��<Zػ�D٪�W��?�yqܫ76P'KމB߀�GR�i@vbrI׏��x	ܲ�td��jx��qٜ���{y�n��#9�Z����;��Ga�p	T�����2�N�M�a�Q��6~EO%pN�@f����-���VQ*0�X��ȗZ�[\�/�T�_�4�����I��v��q>7y��q=B�U5�4^�b�U��O��*�#�8�,[��>g�YN[������0O7K��r6�kV����m�+���31��1���Xˤ��M�+ʅ��*"�A���V���݌�2�B��K����y�����w�C�uWZ��&��Ő� ���6�ލ��޺���ه�����31CrvO�Ҹo�ݴ�1�1Ä3�����sЖ�����j(��
\�l|vpb4���w~�/��)1�sCx������e�]Z�a��+�|j�'������I���/+K^���{h;�&��2F�ޘU�M�}_1{�"Q���w)�\�сx���_�̴�Aݬ0�ٓ�����	m�K��rNPFM�*І<��>�oy�p/lW/ �%a�o$���LB<\��E�������g��s��7�S4�N�5F.� FDj�!��v@B���<��]V�tCԅ�~�B3^�Qp���ʾC�	�]�xk�H��E;>�v
�o����D�"�s�"�ڵ3 '�j�Ii��V�2.T�PU�z�@F�9�5`���I�s��"���?��<c��
�'k��C~�A�P�����JBʦ���Y�x���9���3������z�,������V���TBm/[��{����xqW�8�p}�R�BR�D�F�L�~��;}c�͊��0��DW��t{�p:_�tx9���H�n�Je[d�����Ck���� �`O�R��������X�N�|�&S�j8~O#W���n����z,�85>���.��;�x�j�˃9�B�y5O��4�t�l�s�>���?]NnA����G�z&F���}1��J"�z�U(����EYY�(I�k�(;��RqA�q��>��Q{a��V���������6#� ĥl+gU���&TO7�w���
lM�?xҔ9܊`��*��bK&��%�m 9c����m��g�C �!<!��鬕n>�l�8�s��V���C�v�s�p0�
*���G��G��;�#UOӍ��,V���bggϙ���0li��ג�|�L>g7�Wb�*XSp߽aڽ;�����B+u�n�����t �0!K��bAJ�UT��>v��� �;�kt�q}8�/�A��Â�� ��}P�ռ�$ f���À6�fK��f�9�QR�E+���1�k�i�
��F_�����JL�.F�����;�?�M��yv��FZ��B��2���qĝOFJ۷W�8z^m���[ RYa�xp�u(?]I��[�ܖ���}W�~��W\��1l�.�'J;_h��p=���eF�D6*��y=���2����(,�8�Mx�c��ԍ"t�\�?��u�	m�I쀡_�w�d.b"P��6���x	[9��rL}z����1�!;[��@�sUI�Y;L��	�dT��S�?ޘ�)��kQ����}%ET���~T�]����`�fQ! ��9� ��W���w�l!F��XO��%�1�GW��E�ZT�w��y�]G�t�يW�hLkU��P�2� xŸ)�����g�3��v��xW��m�U՘�	��]hix�gڍ���Ll�����W��-�O9|���}�ݥ�ۜt�U�|K*@�d�#B1���1���#X���]"&CI]�65�n��z3�zaȣ�$�����8�gd"�L�D��H@���h��"(
���gA��θ!���f�v��#7�F|k�?���I[�����v���,���Z���a�D���<@�"V}6�4��,Wɔt���r�X�57�2n��� ɨ)�����c�����|��ac^��deh˚a� �-�;�  +�K���R�������y�k���^^�<ϥ[�f{ֹ�꘿1���)��FW@|��Sv9VD�?PI�4�3�7o8��}x��C^/��,�\{���Jqc���E�εܝ����;�:ڍR�a�m�P�&����e{/�]q�Qdh�6w:!���Y�M��X�6vq��E2�}ɣ�˾F)�U_-
�1��b��9 ���(X�4��p�[;u�(S!y^B���Z��	��GC�&�o���ȇ*�IX�����:e.}"�Y�����t����[���y�[�=�M2$���3k�����qV'�x��q��ʦ<�M�
	�]E��w�B�60*	�l�q�7{Vp%��� X�hyyD��A�B3��'E ڲ�� >! ������*q���	��lc��Y�@�V�C��Re7U8!S�t�������C�݋t�S�H!�5W�`�8[�[k�|�t��͆���t����0�7E�:�;��Nf�����Y�"���v.�!�eN��Q�ՊאY�`�Ք=�7�iӭ��Mo~�����v9�]�A	L�2�g�<}r��L�(��U*��#uq��3ވ��"��u��)D�$���A�{+���8�Jgܰ=<��+��]ԥ�0��<�v��:馏в<�1Yi�XǼ�&q|Xr�MS�6������Q�]�->R":q�f�zI���
^�撱F�پ�M�+�i�@ۦ�R���lĚ�����)��(>�J�+1����IBv�)��x?7��őHW��
}c̘�g&>-�� s���Iz�Z�� H����*��0�$��gWiA룿><��!T=2��������;��In���N��� �z6V�j~�F�g@������?»�|��_P���\, �'�_�q{�<L3Isօ�k��PO��j���2�.�&Xfd9��4��.�x8��K��j��(�F�o�Ң���,���$4�т(��)�e���e8=������΍��*�Ly�o��8!�J�F\1`4��1���%�7�?\~�>!P]�fI��YN��|����@t�i�Kz/����j���q\��L�¸�#&�9���G���q�v?�ر^�o���I�9��	v�;�X�wҘk��91�y�c<g{����V�:�7�I�3a��(04�`�9-�Ѷ̻��P]�����W�g�V&�WQOx�	�u�~���nF�Aw+Fwi�W�B $o�5o�T4�K���v3W��Y��/�����S��6���h�����ܐ0͐���I��a�uxs%���"�o1�_�u�{�|�,��ki�<�{�e���a49��Bg�]�|�$<��"Y}u�x�� ��K����g���#n5��G�eס���YX� s�Wz��W��FQ|$��,]u7��#�;s�L�^'��ڔ�����<b�S��N ��+���Ts\���L`����	����j'O
	��x~@Z�z��)��1D4�B�Ȕt���IW_��5�{��f�ԁ�w2<"a����f.=<�O9�Qb�<�Ȓ�19�-)�M�>���7���kG�Y���~�<%<9hȞuD>bAM{wt��FM���������}]x6E����P�G�]�cq�X�%I`����E��H! ��*|�����Q���)�n�Ɯ^�D��hN�.�庁.�Ab����\�J�A
�����QyT�sh~Q�g������d�@'[Ю�U\���\�A|xT�VVi�'�����%�`�{;�?�T4��mj���N�)u��l�q�"d��Gз���� p��:R�@��s�?��]�K��a����H�{�c_�:��/?7��.�K
���j���I!%Pe�J�_�I����h�O`\�ی}~��So��TMt���=:��jN@ݙ�-�Z�w�cʬCo��đ?�\w?�8ך��P{[��,4|�5C�/ȓӋM�l���0��s��Z�������;e5�eBz�3JX;���<�~�:"]�.9�=��'tC]n.H�?�N[����m�`��qУ��M��!�߭ ��Y�!1g{��p��[)0L���d����C�UM�)F�$0�L��� JlNں��^Â���r4x��6ۮ�8ԭ�/����Һ�Z�5�dO>���џ���٭#�g[�}m꣔�{m�ٵP���C�5����c�O@��u\�`A�=��`��
 LZy'%��h�_�|���ͽ�r�+���L�L�dA����Tm���,>��)4�+u�A���]���h-C�f�O���n5�tO�Gd��A}�$ӣF�E�A�gݑ�()���LT�|,ߚ{#WFs�څ��߀��I�vIOޏ��.~���ߊ0*2)�p%f��b���:�~6��l�>~��7T�4C�mO�&�X����o��}´����٩�]�כH,�k��O+j�pu�[G�h��+�/���P��%&�K�W�/ү2��kp�/9$�������K}Q�ሩ���F�٣���1�:K$V&�+����D�Bĕ#�fb��H}��0�����'=�/}�*ܩo>r;.]�ƺ�՗e���N��*`�K:ԟ���|'>���1�+g�-�����0b�>��lj(��FɺCt��&���c跊 ����tY����d�PP�������r����x�"w��v2���0ĶI�j�%sȹP��m���J2�҈�H��|`�}OHk1�.�ok�����.�.��~Ln�C�p�[J��O�>gS�o%�w�*[�����닖���:�!�ՁdJ�N�e@����G{���"��fo�8�^����F=	�IϢ ]�Q�p�#xw P=�HO�4��v�bB���<2d����+�iV�����[}i&x��$vކZ5��Z��4�����V,{��K�|��+P�d��E<Kd*�#�X1�����ȓ��ʵ��u�)��Ms���R~�%�XTP$jG����}0�+�AF��wXeVN�X�u��g�N�|���'W��3��us���&.f���.D{ 8c���M_���xu��^�nh�1�&��-(���2��RH�`��r��?�V!�t�C�8�4,�Xsѻ,���d����.<�i��*�X/�I�5�͵���`�mi�q	ʴģ.� `X��J�ٿ��4f�:v<0�3͍*$^��U��/r��(+F���"�Nf^�tXs���*|[gG�A���7�/u�� ������m�eY��{�0it(1N����T����y/�	#]k#P#7��2�w�[�ӗ�VhȆᴋJ/�����m��X&:�,J!�5�߬��kj�j���Ͽ->[��}2����!H(�.aJ�j�)�mN�
<�g^ΰQ�Y�?I���o�̨��3�
i\���%�P�!)E������?�M����.&#�1"���3�� 2�1��*�I�A��S?*�3{",�ή���bє�����0��#�x��D�^��<��� xqB���>S���)��T��5T$��n�<�(R�"�`��*��*e�kh,�])G�Bz��*�}�CB(�*���!��{�@)�J��_�M&>2n(Qd|�?"i���	�w֝�"L����wH����>�捨�� ~XV���'��eX�_ynt���9��#����O;�W�K�Wҟ�π����5����7��HlhP��Kx��g.P�]�V8`�YCi}"�����nc�r%�LI��Z���>U�g�]}�
 �4�ڃ�s�M]����r��3@�&��1ZV��:D�tF�6�n���xȃ���~�J�n"��ǧq��;���'+�of�>�P7lT���;�`�퉎��k,S[ʼ�Y�Q1�g��R�j��,iyh�wF��oL��Qž��,4bXQ�D�*�-ĖDT���������{���ن @�z���4Q{�$4z��A����=[��!"ET�~�.�ּ /�x
��D[p{�4Dq!g�q^+d�X�P�F:����6g�mX�1���F�� �OU���H������&r�UW�Ndm�%{c��:�	F���Y\�#�[��!٫ݥ�}R*��>����D�wL���@zn�:.г�
�y�jJX�_.�g$0y�F��׸z�g�����nB�c�t���,XA�\�{gN �~��gn_)+�Cy㵏@Q�G��L������g�@��Q�n�?�KS��<xϾLJ��GY��'O	ؑb�*N�9z��C=}*�A������ݎ]���	���j����f&nm�?qn��:�"����
8>X]%Av//�:�˄�l!Z�I�c����ˮޯ�wݨ��+�[!sF�ו�ˢ�o�sQ����=�b��hJ����0�(�ǻ\b��6�m�ʦ����iSc㣵�0��S�(y�"����Q�e��w�2T����'s0�[��m�n��f����Z���K�fU{L�T!rJ4>�f��dB����m�\��ɇ�Zb"H��0�A6�N��g1v#ko��&e�n�&�`��`�it���v��r?�����G��tsSk,���o�MՖ�n������vh�Z�i�۾"2�ʹ7�s��:u&08��e�U�*v��Q�s�^�!Ix6/��è�2QN��j�
Y3��C���i-U�8�h$qM��:u�x7���:�r�I�rc�4��D�ض��'�VJ%n�a�����]�k3�`�:�a�8�f�/��"ݛ^:4��
Z��8����f:�:���Q1٤��������=�وP5�;�:��]����"�|p�L5�ë�,��T�� �v[6�&�|8X���"Zxl�ގk����}i"M�̺��� �m�X�Z���t��K*�T�ǁ~ꂰF%�8D��=ua����iq�lT�su���Tveꚨ��x��E���g�#���
��qNgyjn���m��I�UmF��WM�{C������؟w;�� ��)&�6�6vi��^���HB�~{Ww)��+G�6ɺ:Ւ(E����{��z�8�E���J{���H#Κ\6�?��i$fp���.U�L?c6ҟ@�6r�A��8Ǿ	�"�?��x��^���T�1��Hy���JAs%F��s�а��f��*�|����T����pgg���Tru2�μ������� ����+1&��{ܖ�*�ȄA;Ǵ	8��KP���H�k�y��� ģa�|�nK��n&�;��G��N7�Q_�~����ḥ�o_V�A Z�9�^�^��H�k}�{�K���-'�̕53O#՚��r�nׯM�|��?9��ϹG�~䣍:08?,=��D;o�DF�����^���~�<h���J&���㙊MH�qצ�)bg�bTԄ���]6�d<��k7*��L=؃�>��� GVcO0����BU	|a�F��kBD^|��Ar���{���[���a�U������.�#ʔ3N�0���Ы7�N;�ih���[��܂Q�$_��7��؅w�t��=BJ�����P�Y^V<p�)ót���p&Ϧ�]�^iW��q��C,�3����:��f����Q��0� �y P��a�E8U��sf�����N鋙P�^OL�#�9N��A%�Me�)}�i8eW2>�Uku�.yX���=u��*(W�*�/��4��U��Lˆ����y���!�E��~����XT����-���G�\`*�ي�Z�V�vӑ��͖��xB,͐Sk5�J�.\������f�l�>�Έ��J-��y���M��9ܖ}�ٙ���޾�PY��Y��E-R�m���'����mҍQ_K�f�8���7$[�,��N�i8B���v���3+�&���`�Qج���E����3	tu��7����]��v,��[H��4�ᶙ�ږ��!�}�Q�?����@ڄ��)�l5o�S��Fyc.-�w���H�nu�|?
�T�l�t���x�hs�s�U�� ޭ' 
�� �JkQ"���
�+��O����b9O��|X�dNΜ,8�f��wI���%�x�5Б}�W���3h��9�hoD����Q�����8���n ��p=S˟gۼ���L���"6��y��ZS��!w�Ő ���̟6��E�J���k
�Jq�֨	�6x��֨'�ct���axo�T-�i���TXH%�������B��I��->���QA�J5T�V��`���	4�;��h{jv��՛��.����A�#�叄>M���>����(|�v���qc\u�h�K����f�G�/pg��ku0��e�4��'�)0o��1YV�ÿ����XG��w5�����v�i�s	��;���=�f�M��v���$��p����!�vuT)c���MgN��r�� �}�o[ Fj�����
��4��K�}>7g��1�o�B�Ě��~�g�P=^[��$g�<��7;(prg�V ~r�rjt�����G�B�CT�^(����� ��rp]�@>'�\^���J���#xԭ�C_u�H_�����{�Q_ڄ����D$��W�<����w
bf5<;�!���U��q^Z<>:5�@8f����:#�>�y>ǗNP1@r���jJs[��&=�e�����u�BmM�)���N"��G�N��.����axf㠙����AX�:x�����	��r7�$��#s���!/ί�r�-�S�7�ύifW5�5zÌ����Z�R@c�%s<Y6��Ѿ�z,���,���������ku¯�<yؘe���2d�˚��P����@���l�`����kǔ�X�\{�Փ	���J�?=��o�$�)b�K�A
���9���S�#d:�b�`I�Ǜ,�ȅ��iHo����YT�{9J��l�Z�!�P��Q4 �/��S�C��������J^�����W��L9s���Q�p���f;�@op�U�''#�]g����Kw+���۫��nX����������9@]���<�#����Vx���ȼ�hVb�gm�'򡈍f[���ҍ_3{4?EyZ�O��chw6�jI�G�h6Jo��P21��>�"�^�9j����cN���0ْZ��IL�W�	���f��r��隸��"�!jsI�,m^��u����p�3���h���)NJ�|�1�o<�e�	${1���IK�s�V��2��+mGC/����j\uƜ_dk�Z��ܱdҝ��Z���*5ƅؚ��J؉B�/�/��w��\�<{^6-�A��iV��џ�8���B�c�M�'�jM��iH�v8�f�p����.�UF��D��--K������UZP�u/�Y}Z�I)��2�f���<�3n�P��ł_5�q�H������0:�R��$�H 1�����.I��0��H��	sX��#�$4�ĺD֤dk�7���5Z}`����N`!��;�P�����^b�����YْZ Ȕ�ϕI��8"�5Q����p�Ժ���� ��q�P="z���㢙"�\oC.xj�O��y�PB�ȱ�sl������(Ze���p�pڜ�o�!e�tt� 8IźR�3�,�jB,f���=�2��[G��W�����Go_`s>X��zXN�:^u�x��R4���9)�p@�2EІ��I�b�w����]�<��4�瀝��A��LX8/�z�R5=5�l[\&tc�w���"���p/�b�QM��t�4�?��C����%9�:�mXs��D�V!$�����+P����W�)Y��~>Q�b�/_s��CB�(iU�c�EI+��_��rOY��:�r��o��{/_zk�d����a��C;���&��e�U?��G����'^��� ~��i�[�(PU��8�����'�G�s���w�p�2H�8L���yS����W�q�,�O�G�i�;,t��n���1,�BTѡ���癩����7�����S'g�����]�'	i�u�+LH�Uӷ����H��Cڎ�ʍO��We�WTܯ�Ƹ@_������|��6zI��Ipz!5y�#��^�^^�*@=x����v]�YlX�K�^��e��u�ڳ�"F�%W>A�[���r��{0e����ɤS\�t��eB����4A�p�j��5� ��,�ٚ�d��#�m����+�j��"+rd|U[h��>J;��Q$Pj�3�%��$ߣ� ��Y��һ8o�^�tD�.�D���Ab��h]/�`�p2�F��ќ:%��ׇtnu;�Yj��x��BB����p�d�$�e�,y��˭��f�0����Xɂ�l�Bv^l@�Uh ��}�Ď� ��k%����7Q�uBCZ5BX��C�8��a��]Tڃ^o����@E �2�Z�r�S�s�~;�'�jS�,~"��Ғ�XT����OW�o�·6�z!33�`��ga��7��ֳ��ܲ���Qp��}�8}*y�`K-Th��uY��z�����z����A��d}M��4<����܆��k_���b�.m^�W,W�A��|�5L�e4�t�F\� �bH�8���__��KEd�����B��M�%�ͫ6�22s*����Tϱ�x�Z� E���v�/��Ye��3�>*Z�;�Q�뀱�3~�o�� �͚浳���Փ�YJj��7�|�4Qݕ�*� !��$��j.+��/�V�<we�l"�������b��:�փ��5�H��.l�����L@OS� }�2����΁s��LR,�̚>����@���C�������Xʭ����� ����R���h�X��ڃt��ҡ�C����2��c ��]ǃu�ѡ�\�C%{j7�-w[��T��x9�u2]�}��I)���IW�a�&5��`%���~H�/�������t�8�=�v��@��'����'�R�wM�O���j`���RB����*��ȡ"cs<XU��>�L,6� �8����nX���i.��e]a�Vp܂�|$�y��y���8�f��޿�O�3��W�P:'�z�.V�g�W���+�W�_�+�gr�V�x�[$F"9�یr{>1X���X�R�zą4=\ ��a�y��X�vFv#	�^&$R��-�D�-�����[�o���ű��� �9���苖F�m*���O�7�~��9E�l2�lm��t>��������ކ����^�y�!2Vo�~�$3��]!nG���ڤ�2�� ��#��3y����,���T���C[���.�m!&�H}gQ�;�V~���l�}�(L-
PPGO�$
T�K�E��D��F�� ٨	-=;QO��a><kq��:_Dp$�T[�;۰\WV�)e�$<��/�!2�m:[����y(��Ï���S| �DX����(W*+_�WH~�/&K���6(��~�Sz���)��V?&^��1# v�[���]�����A-C!������n�^4s���$���"캯`tX{Â�KD�f���Ӫ��S�}�^|.Z6"|���������ɦ�z�>�0���7{y2�E?yoT��3��E�Ⱥ���9	�$fZ�_���b�cm���٠<�0�|�t����7���c�0_f�r�p��n�MX��ǾHb�Y9u�9@�K�np�	�S|ξ5�����md��;���8)��z�%��Oa�Q�<_�E��T���$�}���%��3��y-^�����pWBi/��v>x����n��5��>i4���_�ZUQ�oZK���q:C|���;�-�D𞻘����k��"�Yt#�@��;,�ܰN��e�Xh��䣙��=����H��_)P��t�y;���轖���._��Y��XZ���ʷ]]~�;�}8*�bؤ\,��~4U֎�H�'J�ޯn���C̞l~._�[�B��ݍk�v��]�3�U�b����\��3�{�s,Z����0u��?��PAf��F�Y�*��p��#�"�<`�hU��׬\���������M�&"������~���3Gݞ��yW&*i4�׊4��-�մ)ER�qp���U���%<~%W^c=.,8�rCF�*��E�.�����J�P����*-82s��UY�]lr=��=�?��ߓ*l���C li5=�Ryr|,�Q턋t��I��A!����������M��Q�!��V`�k�@$S���(m �T�c�e)���Y��? ��ҩTP����7qY&�j>�B��t\O�0�+r�/���D�)`S���4N¶於���hx�v���ˠ�X�6�I7��Le���jj���K���E!|C�T�C��N�:�O�j�r@�֥�h����7Ґ�wi>fУ�x�x��b�#b��FLǙ�����Dt��<�F:�w��ࣽi�?i����kz�a
̔K��+�'���4��(�{G!\CF��Sm�����F��J=맮���M6�����zo>�e�+�=2����<����SPP�:�G�ՔNnz=Cr�_
�;��K�s��/�e99@u�qR��,BGD�(KW�_�C&Ld��� ])M�������5ɺ�!���.��-Ά�&ʆW�P�����֎�]��1mlK;����
�A�lk�� @[d�me�����qn���y�aɭ�*51!�T��~$yd?��RG[6�nti����G+� ·޷�ٞn����yn9�,x�E�����g�����ccX�͑.q�h�v(njd��������K���^�νJ���E���K+�&�	 %���:��ܜ��& �/�=Uk�V~%?J���OV2�z%v}��&�����c���&ֈ����)T"�Ӵ,rZ�L����RҲ/������j�Ykk�A}�1ٮ��� [;x�K�/@ǣ�cnt�[�Z�<��0�)E��#�G E#wdO��!��)<��E�)$��G�6B�BJm��\+��G�<~����w��l8=�TD�,�u6r�֢$B� TT�Y�|\�Y��Az�I��j�<����������F(�SWb�d��������J���B�����~�[�0  �Oc-Nq	�S����q��EX�m�c&#���bB5K�\7.���?���Q;��c�1%�:bl�E�ln�+C��0A`���'
�A�|�P9q�[��#�9��M�L��['��7�DC���3�8p��K��C��ς.D�Z��C��;N��X3�p��8�df_AE
 �܆���:mAg��{�p��Hk��:�jZ�����b��У�&t
v�>����*�_xlG����������ڱ8rVi�̰��
e"5�.�&+O���Z��󱜅�r��""�[h� !��t�S�W���b(�Cō �4�#�9̝@q8&O��
�m�K����tj���W4�bέi�/��d��I�F���|cd���d�^A�\q��ۨ���.��÷�k�;~T�#�,~�RO�
w/�C衉Ne��?���*���8;�`��j����k�����$�-��(sbOb�'�]�B�ѥ&�	�S�X�w?�I��4�M�����X,���մK���:�������T-��O+�6�)2��G����(TJ%�#~��O��[�;>�}a/�>������.iɜ-�"�9�V��[��z"�G8:�Q��v��-pR�4\2I����3w�F���7�a��%Џ�u~�q�����v[ 	�y��������.h�e��.e�����Fľ��'Ҋ<�N70��Orh�qsc�:�����2��M��	�@jµ*�͗���*S^bq(?�CA��]}���l��lj�8��
r0�c���.��Kh+�1e����ӜTT�q��=�������V��_����3=>�QF�S�E��Mu��16�dq�`���pXl0=�j�:�/ �hѵ %Y�M�߱Trs��|���#�}�ԺP��̜����o���9a}8�t2�rNaM����^�S C5�VԕbG(T�LY!g.��*���>�JP��Yq��^�S/�h�A+ �AL���m��O#F�H�Z3�Y�t�{+�u�v뛀��/+�|i;��|�jkO�h�"h����p*gȮ�n�
����>�9y���U�d+�b�c�w&���+uwU����HW�e��?T�K�|�9��Ţ����TfW�\���)�<�)Px�V��'�z����P�-����q^����X/����"��?��t�#�������_�v�A�/,������'��f��ٗ�/"�WZ�B��'Y}���^I��������@LDt&ډV�u�p��$Y_he��Ầ�Equ�Be�QP{%|��S�D	�r�]ja�ժcu��lqy�?'e��;gڗ��=!x��!���  ���X�nh�����R�$��y�_YCg����F�q��kR_�^	'�ܳE�e��=������g�]���/�]f$���U���﹣CM�.��Xd�T��)ul��yb��kp���0v?K{<���1��YJ˲���0��8d��{�cn�8�_$���U��e�0�����z�2���ݠ����/;	'�i��ɞl>����$pGك��dd�QI��L��hz��W�,Y����X��E�#�����7���ɥ~�0�=�z�Q�c\��FA~/+G�(���,���=hQTޅ��.��H��k�^A��1 ��j� ����hr��s^��eཇ�����o�%���ȥ�߷G�F<��x�*���Z&0a�)H�DJ��s57I�t�d������#�l�w&5��н���0~�Q^��g~�������5a!y��uR���v+{d���m;֪be��B�y�U���&}�Sյа����ro@6���u{w�U��
��H��.
�t�.�QH�^����;��Q7�;5���d�N	�1��	�@��K�r8��覃�,�<��&z���Ѝ�>�!O�I*z��'{}�+���ڌ̿e�`Ͻ}���x����HP�Z�K�l-���4a���1
O�/41��P{��9=8w=�qQJT)M{�b8~����ʂ� Q�f9_ab���:�0��;���8��du����x��.�{�u:���>vl�7�p��c�O	��I{�`��֫���㾁��:q�kY�]�)K|��V�ݭ=}��I�0�=�oi�D�@�@�T�O�L���ʏ��F�j�̺�tXT+����
��5�(�� �ljŠ�4�0AL�=�6��)咞"H广/:���۬�dfdf%�k�����r��ە�6�y�?kL���Um��T2���Om���QO�NU���%���G�O�a����H	��jw�/z�0�E�e�.��3�y.a�+@'Q�_�d�� `f�d�CO!x�D�1(5��>������g�-%�`rF��{�9�n�11q�S��#�p��h�ry�|���:>�\�<-��۝y�QkQ0"O ��ϊ"{T0珲��j	�.Ä��v���bAЬ�_9����k�͏���׍�:RF�7yk��@��܌��A]qL��y[�M�#�O_�� ��S].l!� Ҡ��_����e-0�!h�-�ϟ�y�?�P��_M0	=I�N1�o]��|_CD2�\r����Q�B��{�K�EJ�~��|�(�O�s�-�-���r(�da�֕[E��$s�b#O���4Ѭѥ�#��CW%gldp��՝�>���[����|d��RA�1�UO_�2�"@�}��}b��;�#N�>v�9�Y�Z���i��O����V4t��e��[�	�G��y0�a����=s�2��~Ȅ�Wg�b%S��������59��	a�[R��;�!T�g�����H�� �qn�����D�E��:^��lo����;�Ҏ��m�tNjj�u5��bQ�q+��v��R��}�^
����_�72S��������S�t���0]������R��솎m���y��q{�C�NZ���뜿8��Ǿ��+��W�ۣG���U�B��t�4�*�ڃ�϶+<+�by	�_�RUoU���x�7�qv-�Ħ��e>)r��ס�S��rմ����A�Y'x�N;�-�Sh�v���H��T ��ʩB*��q���?0EF���і�<}.��uR������4b��>�!o�xa���bĒ(�E��C��<`*_�U�ԝ�묹��ۋ�f�eN��@��7o���[{�L(���D����k��Hz�7;�y`�A���^ŏ53`M��\���*�F�##1���og*E�d�[<t�>/���;(A����f����`�����'%�y��R���L��Uw��K���aL��g�2��R�̎���8�Zw7+�fű��$S���s7Q�B��\��e��JE��T�S�K��C�ۖv�1���� ��p)��V�9�7���ft���j�����;C�κ�.�܌�P�	(R{yXw�/��y���9�&��-��xu
�R����1*!G|Pt��'���7�Wzc�Ee,��NvҘ��ݳ���a������1���'��՜�^c�����a�;�ݥL|����yJ�r�U*��<�X&�%��{���K�2�54`� 2^�O1$�P�.7��FU!^�(X�Y��2$XH��Е������4�
��r��V/����*�.�"
�R�lVkƊ���b���0�`�0|�cʀ����i��,"���o�ٍ9���$��<�#kgn"���x7ho�D��h�7q���_�2���;���5A;��F�c�W����/�.�?�@�l������ ��&��M�"��y��u��K5�wq*�PRh�����[�q�{n��|%���]��qˣ�<���K���4��&��2P`��ݼ@O�'O����} �Я�JI(#�G��v�<ߞ��W����-���N�[~z������mJ<��������z��Q�3Ќ��ը3� �Z��d)*mXw0oorp�7�~GXחxDpJ��i��[?7u����Yz��HO�A0vS�p[X)�2�E��,Ñlj7-���1�٠2\�B;�f���&�l�]������O�J@���u�u�sd��)"����[���D�i����$bV�6��s�<���:$��n ,��$�??�����l�b�-+~���	��6�ج)��jЙ�>L��j�X|pA`��'��!w��N	Q��=~���^R����;h�.�V�|��>�"�Tͼ�5��s�Ì6
���^�űE�ORʠ'��(\�~�M��@�Rr�2���OCx�57�r��Z �d;���b�Mqe� G��D��
�"��5��H_䜅���?��.��2�Ūa����6{�Կ��� ���d�Y��)���!=MT*�
��<B#jH��n��T$�X�֩",ȻFR�?�+'�f� ����2�Z�Hh������8b�]�+s��mGR�]�kgl0�H��p�.ǽr�V�A	�̛eՇ��~_���6�ga]��d7��|qb˓ �F��OE3l#3:�5�)�~�A!:�͚H�������-�����>��h�3�B�+@X�]��������*1<�&[�S�`�8^�ʛ_�#�����_�:�b7^C�)����f՟���\a�֟* �[����!��H����4�;J�"���D	��ղI�Urt���h�P��O�it�!�۠$\�>U=��8q9�Uy�xvwƹG��?���^H2\ߊʨE"��k�Wb�N^N'f9.W����i�lo�CA�`OK˂�=ȻO���k�ߢ2\���鹀\ b��>�d|��h��&n��,���:��n�L��k.j�ǌ�< �����y���foҠ*}�[�,
�|LN�\�����t (<���������G�>�L�m_C�9GO�J/��Wwꉭ^( ��	�e\��G�7ib�Uҷ*�H�B@2c����ͥ�x;
�k:.E� �X���2�x
X6�
��s��'�Pey)�v���iHiJ^��>�v�|�Sv��6�ă�<(5���ߖ:7�*Gv���o�B�$R�j��(zm���c�R¢��DL��2��ַ�r��!�y^��( ?��,/LaԚO�W�~���}oԞ��߶�CQ��]t�����f�?��_FP� �/�܀�j�y��O�D	�
�zZ�x�g�8��1�{Q-/:����3�l|W��]���^�
c0��՞��x������#�7zMȦLzM�T�EBf�Q�J=9����.����v��0g�"��eq���8�6�?�l�w�P������m�]5<3�Sf�_ۏ��	��������+Ks67�L�aK��5�咺�ҡ��g��&�5�PE� ��y�Q�Ildj��k����9���{�tRL^)�r����^��a,f7�O}(��l�����!F��*��<"7�O>��<��g�n�}�,|K����;���nx�1���h�]�;[&:�T.n0I���]J^������Q3��%L��J�?�o�r�����{3���kS�p�Jҫ�H�Y����C{ߟ���k<��gfr9�=A��oQx��TӃ�0�p���^� ��?�r/
!V�j�w��	դ��@:�"+�3�/Q_��1r$хG��ؕ��ڄ���1m���9����	x��f��0��g�#��&�k莄,.�wn��8�m�NwSB!�(a�F��yҡ���`�hZ*�!(pk>��9���|�Y?���&���5������qz�T��f�M\p*�
�^�bL�R-	�+�P������ar�d��'��/�aq
f�i�)��I�l-<v��"�@�.FH@�2��[Ƌ�,̌x�?��:����yF���p �C
��
��B4���\�3����ʆ�z����#��6��h?c��g��־�N����r��L楯����R鳀�(r՜���pd�K�6]nN��N�
��n����$��"#a` �ҷ�Ag}u}��]����c���]2l����)Hwne�
Ǐ	a�.I�|I�&q�Pmˢ(�Kfs;���z۳�D�\��Zѷ2۝�t�x�����t�c������ �,~�?����x��W�V�%�3��GD�bDj(n�˙7�S�aW��Ù���
5�S� ����6�sJEjxd�lp��=B�J�_��}�TI<Љ���Y��*�Ꚓ��`�����;�ʬ����{h�dʐ<Rr����h��Mi��L�}-u!��Z4��ޕX��/sy6��$�%=v{,�f��t���#5�U�@J�|�4��=;��
eB��i��V����d/��Wm!a+���m�� ����g�m�e��i��(;�x�i�Q#S��PFb2��ei��'~b�'�w!�V�Hq��X�
��0�ټ�<6IOqo�� T�&��٢no�,"}La+:��,��o~������U�_p�+�}�K��=��t\��:�gE�B)������f#t�)*��,�Rv[�un�4��ۥ�gw��S/q��A�hЂd?7{��#���(�I-	%�1��@�6���I]��N��)'������o��=5��.(1,}BY�3b�$�Q��vd^��!�>[�
����������a�G�_x7�
�BGc��O��0�{w؀Ue>�c� E�,��4����hba멈��l`ϱ`���6HLӋ�d��Y��y�\�m��
 ^t�yg���ZP�^���F]F!�ȠE����v��:V�u4FI����[;���l���;	��q��8�1�Hڱ�6M�N��Dy�r����)c��Ɨ=��ꌅc�Ozwyr7&�f T�i|�_�m�Gg]��>�����n���lE�&�H�u��ɲ�ƌm�ǡL��dpw�p.��5�{0��=
����QCK�nڒڶ�,���)��"$U�XK&������5�����u��@]7���cZ�U���5�LY��ͼ"��^2�6ˇs*���eX_�o-&o�W��C9�ڝv;6�
�0��m F!v�����[�́�6�1���0L�+=jO�)"ֈ�]��-���	�<�n�"/�J�_�ٿ׋�˅;��ڼj�r��]%
ža>��*"��o��+��$[\9�?�5?r��($=�����K2���_ar~�ID����h�<b�nJs���g�6�t�0�½�E�e���U?&fx(�aBE��#��zH�gz���R�O�����m(ڨ����PyWk3[���z�ٚ�y�nO�j��OsG��]m�������W���4��zxî
5��l�xD�oN�}�N�����Dt_��k�2���;:���p%'�˧@�F�K����# �N�;�i��3.&�N�K�0
���}�7(���A$��]���YЍ��KHޏ*ݵ����:{3'���o-�;�g5��1���78)|շ�]��f�(!+�F������\��7O\Ux�s��A&��W��r�i�1_��P��I<H��߼�uh7��w�ӡ���خ!��)}��I �6єh�"����J�P������\�����@yN�WG�����yi��-+L���<"�F��E���G�g}{�+�[�R��b�l��<�)��+����ɰ� F�LSCr�%l��֭;**�;����8��P�Pğ4�I�6��WVPO�AG?�_��л� �waK�5���6��Ⱦ:MB��d�(ò�}�ᳮ&ن�@�/2������RL���3���Z���r34�F��U�F�K@ՄKQ��k����h�n:t����/�>E�J���K����Go'��m!
��w٫�����ơbh��z�zUX��?.~�����xM�'���S����hJPq��\i�Z�@v]�|NY=�ʞ��1��j����q���^�&Z��TsU��;ۈ�(���"��˪�O�4&Fk���<{ڭ���=�	�AEա�Ҳ�p�f���ЬУ\s|�F;��ÄI�&Ћ__�%��ю{L��� S�OO&H��	��TUa�GM�n��r7�!�rF��������ɏ�r��&¸S.�3@:xX��J4��T/:�O7�(>�u����ɖּ8L謹���cՕ�j�7�Q:�W9+b?φ5�[T��).T]��r�  k��[�K t��^�y���Z��Vl8�c��Q-���+�V��B�¹�Q���ϕF�i)�6�m��y�,(c$���5��/��Ud p\��K�|�t��[�!`}��2RgRxa����ˆ��?S4N9r����X�����bMC>�$ěH�+�/:^����S�H:�lOWk����(īX�ߥư��Z-�LL�#����cn�p=��`��
��:�tH��Nm���8��p��{��Z>����I\�k׌���IC��ElF���7�dڹâ�O�d�f��k�?��N��ZP0�����'�3��ɣ��.�x���%���H��O����^2o�_��c
v�O6ξ��9�z�5��E�%2G�i+�1h�V���	���Ǎ�<��*Z����C\�L��ny��&�*6b���L?[� �$ �K~Sk�SX�e�w:VW���ET�fWPi�ni�n�; h� -1#U|ʹ2�ʦk֐3D+�p���Z���p���,��;H�1Jt���� ���ǀ�8vGkP�	H��q�F�BlQסm�}v�#1S�	��y+�c����et����v�럃�D0þ+��<�wf�M�M`Ei<��L���.�ь�Yz�Й`��~��E�Eh�h�G��n�������6D�9D�/�V��qTB��)�H-��]
����[�u��H�n���v���r����d�ʰ����9�L��RK7�P�cV(��OL֧,0�,��BQ�RC�7=���W�h�n�� ���Ό���Կ+��mF���Fq�K���m���L��i�fo��Q3k���6�uSx�i쬘P�pb�YW^��Y�F.�N6E�a����C�5���������=3�U~�������8"O6(*�g�p�uQc�+�����h�>+� Q�C;�V�"�G�e�s��&�%4D�/{��͵�ZT�(Q
��E�5�:�R	j�4�;�3J��HfW�9�~�x��\~G4~�S�!܁�y�jZs�PW�	��x��F����r�[z�dGB8O�xȊLg��T�'Y_��*v��dކ��
��� xխ_�����1lJ4�	�c3 [/�,=��:.��nM�ױ�^�5f�wMb
�M5��� )�����}�5t��_��:$MuKK-�$V򪥝 �L}��5��R~/�Y�K �iKz������f�bb٥�j�E%
p�t)� �T��1PD�(��r��"