��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��t��t�!����֝{�ӓ�[q�Ѡ�Bʌ4�Pq�{�@I!�wz,}r�����:!N�� ���hZ9I���a���ֵ���U��㍽�����ޤFk��ic_Ow'�����
�J|wn?[.���� xd�=mq%�P�3��B%B*b�^�� k� l�n�a��o�����$.v�ϡ�O���CV�<�
����=�)u�t|�
i|
O��E3����baisѯ^#
�	2�c	0E85@��Zl����hO��a5�)�ʪuI�x��S��\	�mfL4H���a驞,���!~�u Uh��b(���x�&� �
	�����8ɢ���!0�+��BJ�(0W�J�e��g� &y�""�%��٬�0�B�����_��&@	����a���?�m����S�������s/�_��p��m�l�Z��/�	i.(H��R�C��%�E[h.]�A<��N%� �/��\8Y��|�һ[F���6E�Tj�
�G����t�w�I��
b�k?f���"aޯ���^	�A��'G�g���xNh��fk3TCq;ɠ^�gp�X"�����Ԙ�����j�Ԣ'�������0�N�ʩ��\�P����j?�9��e׶H�0�c'�HwS�֍�n&wpxu���,�j�|�m��}��~AT<EfIc���M�1 i�Z�tZG7���5�{H5b	����΄�DO�����8~��C�ѝ� ~Ģ7�ފGם�8afiҟD���~�������TbY��Z�A~��n���>_]lO*��Q)�N-�^Q�g��ܬw��5^JW���"R]�]u��Rވ�pk�P�;< ���n�T�j�1��f\7�-���<$�~嚙�w�>����|<�7�-wj��*��yeC@c�2���I�)џ��U 0 �����Y{�U֗u���n�N\�h7�����U+'P+����r����*����&��Њ\����)
n�)��x�qmL�l��J�,oL~ ��c�%%�{��,�=�كO�clg����U�?n4���z2k/��|㗁���=-`�H�c2�YI2�ȌB(uXμ���/�z��Pq�� ��C��Z�ߥ� �VN|`�`X%��&�����[,�T5ݺ�%E���)"�N��3C$\��}��jRq�RN[`rW��C��-P���-�a>U�~�S�J�Q<.E�9�������ev�`,	'-k��o��CZpFmK!��aJ�w�?Ů��ʛ[ \^-��]Đ�����kBl�o$�$��<;g�M$��S�Snk�_���>V��pf��c<	��!��%�C�����Vl��W���u��ѧ��'TW}�#�d!&���H�ݭc
��uf�b���"P���5�R�Ln/�\���C���P����E�i�g��x�Z�#*Û\�!��)�
�_c��&�^� 5�6���2��g���U������Y���~#�v{��"�8�7���4�������S�|��*	Q�(;/U1��G#M�'�lT�6~m[�\K.��'JB~��a�1M����ߒ�cU�o�cN`-ih�x���n�������{��y-�Qe���h�h �.��P��Vk�\�֝8�}���P`�x�U0���>O��ݥ��9��K�D����Q��|}��O3�)� :l�6���-��Ù׬i����+iV����������|�M@�)-�On5ѧ��g?���W[�bw�Z �N�@��@����y��/��ED��r*M����@��: �+!�j*��:������AC�u\
�g��'2��&���v_���;���-��%��%��p8�-��uW������c��P�����G�Z�]�Es6���_�,\��K�p�� �Ӈ(1�\P�ߏ�"^\�|�y��U ���k�O��q���w�	����ؽq�p'�!�s@v;�����{e�]�\ƀ��Y�b�PkF�l�/q/)���%^�l�
I[�{(梢�_���<g8�	�	v����"���;��?�cUپ�ʌs'��ۃZ���h|o�+!4����[����t�C�x)�)z:�=�sߗuL���oi� E����t,���Zjuŋ�d�{�T ���S��7������ʐ
B����������u�,*�~~�����.�z)����ɺ�(�!� 6_�$�ա���B��q��}�2�����o
bv�l��<� ��b{6��=��I�FK�{������ϙ[����KP�������$�ўR�F���@<�c<x�]�3����B'T�_t���#��gF�;�9�pOo���i!ǘ�tPb�|��a"�/Zb+V�?�ɳuǠ@%��#�AW��)�oV�  JKXo�?l���Hw@7O˒Q]We5��\Mĭ���ɪ}�o�j��V�BL��/�x���2�`y�C�+'�� #��O'���Wk�4}�5	�4S?$(֥�Hm��H}P$ ����2���������"������$BJ���R�y:�Eȿ'PVʹ�(��P���W1� ���a�DT&��N�Ҹ�_'��i��ZS`���}���m1)�9��7�GY�p�����r?�r�����~۫�w���Q�d�I�0=|��B%myLy��	�(�tZ�vL`C��:�Ό����&J�/"Mp7W!�<�x����Jm.f�k��ˍVJ]iHDm&��g��}Y�ʛ�I% ����u�� �� �O��<��#Vf��6T�v��)S��e;����{D3\�oJ��8S�?��<����h*Wb��T���Ȁ9m�'ͳL������c$a;�t��7���^�WD���V۽����!i]��_�	ӥ���'�Ѽy��I�8Ia6-&"6��-��X��7�+���֏��2��f�M� $5Σ��t���?�ns��l�2I��5���U� 3S�U�r�܎V 9��k��3����3�Y�|0���V�C��)H_�.3��IR]؇�T��x���;��[1:E:�P�焢����f8��Fޕ�û��Ä0�|l�a��~��R�f���-����yJ� m��=|� ���7,H(cj2�8;̭�L��MV	���h�� jB?��î�/>Կڪ��h��������'��~�o�{��"�$>v�8L���7W����(u��b��F�%TX�msw0C=�C��1=+6l��V�/3��Ύ,𮆿���@=���!	�d��īj$��ʂ6�ӈ�Z�}q`&�u%�Ųg8vWg4!v�ٱ�Q��֪�b���yr!UV�������T���QY�![����ro]$d[]r+
�Ą���+ݲ��5i���%q,�^���բR�"�d��k{�*_E�jWJ�+vG���j1<�{�
�����F �<�.�b�<*H_Sl�����{A�Y%�[0Q��+L�}�7*��z�źg�-oM�,p ʇ�X��ˤ$N�D�!�hu84��߭T�qV5�oͪ�u���m����'lv*��v�Fl�~�x�t�q�d�o��I��{'aҽ_]P����c:2�C��r�(�Q��3��TG�ΰ�k�� @(��2!+�$U�~|5��B dWVKܧMt�u��p'<��vdxR���p'�A꣟��p=���y��t��m�	Ͽ�޲��!��o����<%��2��q�?��tO��q�n��G��̕%kǂj)]6�ڞU�\��+ٻ�}��+cx�I�����p��H�M{�����BRx����g�2e�p"O$`�p#62�̣h-��Xy������ڀ�H��_uT�k<�ܞ�ښ9-b��b; �ke��x������p��Ԉw |��=��1Z%�����>�r.�u
�d�
fFbj��.7����qh=Z�g}�Rm�r>]�">n�!$s~���r�ySz��F!���i��9ͨ.�R��O��#�FO3l�Nv�3	p?o��)�k��y����މ��ɼnѼiB%��^Q��M�ޞ�M�3���	���iq����� �4ъbD�O��h�'#}�}:]���am%�Mv�U��B��}�X����~;8>#���3:_'��m;���!��׸T����O�..9F��>��/r�'MkXP��gR\߫���W�M`܍Xm�?�Q'Ξ���Z���xw�/.�R�����V���Ac蚿/a�S�琉0A���\j�<�� ��A��}1/X�CC�@ݥm�H$�dӆm@:9P��3gA�*��A��ǙtN�
��$�֡��8�y♞͟E������In�:3GnVo ��3�4�����K�&��Γ[��?s~�]d0C���Q��<�����^ė�����r���>���٣&�%��HFs6�d�Pc�5zX���M+��^+ӑ6��3�%Ėn�V`�'�"�(��Q�H�f���Iq4�fn�O��v�=l34�Y�qR�Y��Fݎ�)�/��I�ͱQ.A��vҮ��q7�S`p���:��ƂݸF�:ކA�i_Ts�3���|�8�����U
��E��ڇ��g�x�`Կ�d@�آ#
�x�??����;����ֲ�h�q$a �7v�s`�k���V��ȍ�v�'d�����'n���WɁ*�� �7向H/��&əp[T�����@R=T�f���(�Թ�s\P��̤#���a��䋭��k����V�:8�Л���q�>E|PSt�@sc2P5�E�쯄+���6�n���5A������}#�/Hh����R���gp�����BS��3�< ��O��+!�~���ߌ��W�xk����U���ސ�����v��6�cJ�BQi�zDO#�[8N���+׏�8���y�6�=���}k(eR�gT�C�.�	�)7���L�
Y��ݷ���$�0�gY�i�v��yѕD{���F�2N��ү֟iB)w���٤�#ӏ಻���qF�|㡬��^��I�� �b��=7�=�2�g.�T(�9<��Uh�syA��x-�<�`�ł��yL��hx��?�zƛ�c�^�\PD~���Сk�#-���qhR��%iWv�:>W<vn�V4�ϖ�l'U�|1�7��]��wQ	9j��<����\0WMVC����S��MK2@y�����bAO��	n����#S�v<������ ړ���h䏅�N->��?�Pܡ	����+y5�˃A�&$q��-P�3,o�tӒMIV���]�uO/Q��T�q��=�L��&�f��N�֥R�C�g�RХP��J�>�B��'x����g�[��a�l키�
ơ����EG�F֤�(���X�J�s���Qj��s�E\x��>�!>�肰 {��d4J��Y�e���ɷ�Q����b�H4�Zi@^\�"��l�M�W+wG"Z�9��p��W�B�w�s��
�����3��Z��]��;#US�ė^��k��ކj�V�]g��ю��0~�|�'x��v��GP+3i�v�-�A��?*����[^���X�/�dӣ'0i=�L���0�~���Y*��^2�dQI`��.N(� a�=����wdm6�q��^ovDI�V�VZ�=�p]2�ë�G]M�,���	ߨQWm�V��s�`��AA�����Ԣ�X�Bt�a4��������G0����K.����uoa�q��"��~���)%{�c��}9���/�����p���yF6r���ҧ-"�I���9�;�w,С�����c�g{΅WpL?|]�__V����HꙬE;�b�]c��g ��M~K�C�MA�z��HqI������TT c�K�Z�F�))��7�F����o�Pfπ�S��џ��R�'�x1��5���ȗ39XҾ݈��+e��՞���F0���6N5����Us�Sz�ۥѶ�[��S�ҽr��Գ��0�hB�3���d��F܊tdX�RE�ITx(l����!������4d,�DE��������ɱp.ccf��fV	A�N�K$��3LX�V|�>�7{ (PV*�nM���)��͘�y�X;�Վ��|EIA��2ˍ���W���M3�T����%�d2V�i��D[욋O�!a�k�o�?�[�+4	*�t�OD�ʫj�4QJw�.�Xm�+�W�<kn-mIt�����x���H_�!�t�(�F���@Bt����=�ʰR����
hg�x	�;s���ō{������+�4�D���� z.��Ͻp�M��V�7 [HK��>>�K\d�t�b4�&�-Ak�Z��"���^B���'���[@kǓ�q�l3A���o�!m'1�:��h�W���E��n*�IC��������7su����9�7@�7����,�O�v�s��f2O���"�;4׳��q8
7&`��Ž�D��M�3�/��]��^X'�<E�4��(|��@
����=���<�-Em���+�MCY@����u����/�@Nj��NB��÷��"uZRVʮ��r�xZ�y���-�T��?��]�b��')��bz�J��k|{r4�N\H���5=��u��0�2(�6�y�7�=��M6�F�c8یpX��-n7��:'����IͅށZc�VG��0�ٽ$���T<4e���$��9n�����K�p[Ⱦ���a5V���Ǚ#N4w$i�qB���T��$��I��fP�4��}[}���F%��#GL�/����T��� ��d��-��N�����- n��뚓kΐ� s��- =R<*���/t]�I��;���׌~��@�'��`̴�����.�����=�j�J���d����_����&�{�v�/�=��e9�E�\a�m��iԺ�D������p�%�g���U�w�L%uZ,��^ڹ*x���D�O;�k{�ea�!$p��ڼH�^%��:�)}�����<���^P�c�8�,Uw���NÇ�?�)�����)k/$�ş�S�)�6���dO��a��f�{�Ɩ�؛���Wo��qO���eق��?Z;-��n����j�-���� U�o�P�<,EV�U*~^�m����`�]^����
h���& ���^�$˞�Xxʺ�U:�g����={xE*_}+�4Є��1�?Vy�0�P;	��� +���6��׾7"�^�/[	ёgA@<k�9^��V[SC�E���ˍjiXf9=��aE��z�8{��MxjMb^	^(a�t|� ���R����f�u+װ(+�9ߜW�M�B�2z��Uǚ 'E�����N ��ô����R�t���;��p�~����H`.�j��A]��3�47(��أBO>Fy��x��VA%C�a{"}����0�ğ͝UM	���[d�����r~��F�)Ī�Eh�+�����}��L[��֘��+��-�[���n�Mskm��bcO�A���z-�h�� �e��e��_���3�����r�~ͨ�f�4��S�1�ӻ?Y��e���D`�$j�7;����!~:DA%���8�?���q�g{���o
��֤P,�}�,�s,H��%�jF%ϒbW%��/kt��xO�;TXƮ�l�w����7Hj����9����{�cvӌ� �4�{ Z$0�\E(cy��Q����x ى�l<T�_��J5!e�e2��rGW2B�a���/U���C3=�ĩ�6�\��|�C@c�Z���� {�P-d�VḰH�'��b��jOi�H�qyq&����֘W.�t�����C��s ��z��0���|��ְ�jK�+�X+<��4�w��'�6���IPI�g����Ί���5�c�v�.Wf<o���y��z���O����N���� ��ڢ�3t���U��w�L���X�F��P5I��-��>&�H��PE��x�?�lQ��QH5t��%�����x�ɼ�B�q��3�vo{��7��*����lh�p�'��{-Je�����P�w��yt�P�A��濲T(�n'
�x=,9|�rn�`X�A��ڛ!�(4���k&�eڔ��N��}�Y|�.�9�$�4�Q֔)a�<��0����s��}(h���7��z�x���X��C���w؀�� ��cmÙ�)�E�rt���?�\����jOGo]�u����u4�>���;���i����"N�ٗ2=$7�`��M��\�7J� �5�9UFl$�LـS�;P^�m.�n�JD���{���
�,*C�#������/u���Xl����_K����V	D~�u=�M�@萣B՜�����MXy\s:�9�_X�遹�B3�Qߗ�����A�,�GݤV���Q�ռ'P�S�QW��GX�4��;'����zx�C4O4�\�g|�I��}��Aؒ��{�)����8N)컊���#�G����v����R���
������i�n�{D���;�!�h���58*�#Ҩ3��-�BzB3�[���:�cG4�;�{g���na~�K��RSQj��tn�g�`S�����ؽ�x�^P�DTU�=�Vދ3[-m��(�6G�j�C����?�wZŒ��6�Ω����{�H<;8�#���.��X�Ӽ$; G�Q�y\����ƺQ�`ZI���T7RWan��X��ɍ.��!p/T卑�&�#@�W�)fצ�K��T�a�vgl�f�hr��#Er�β�#�]�mZ;(P��^#�����aPB1��n�?�^YsF����zUM�_�>-@��
�O}O�?7�⏗��Q`7U&���	�p�l�Tn,/X�����Hc'��ko�
�h�<�#TI"�����it�g��["2���ܚ=���L��s=��xxg�\�r*�����`֝N�f1,�<��Z�7>��e����9�b�4�]�>�0J��&N�ڤ����C40_���I]^B�� �됒D�!�e=���3H�R=�`b-\�g~L��l�>O���UN_ n�@&����B����h���+�5[�cR��1]c�F�m�D<�+!>/��c-dJ�[40��=ʤdE�խbB.�Pn��>�氚PO��"]5[��L����Q�:�Y��v�B��6;�'밢#����Zаl����H����w@�2����u�5�H��Jc�~!��M�(w ��B�����ڶ��b���0E;K*��	��W��O�'[Ott���!i_��c�Ty�����DQ�B�
����Qo��wxb��ۥR��ן��p��N�(�o?�5�(wK��2� �-��_����wۣ���A<��[���8b��{�k�Wt��c��Yjrl�k�k���/<�<���l���[��׵��F�aR��Y����ʑԾ���3��|�WH�?��q4�YQ���uJ<s���k(+K��I<� � �J��˜~T����Ss���ֿi�[���"M^*T+��CR0 U+�ϰ��
v�?�3H���P٭��w��٢�N�8�u�����g�$
iZ���׽ʄ�����p�u��z�J�����KwO�Z��b��κu#M��*�WL��N���|-�~)\Zt LJ�K^-8���lн���H�xr~�&v^�V���;|�Y�q2�v~I9������E��?f�[��]Haг`�&�륚I��e��>(�N��hL�rff��RW���	-��[���4iKջJ_�ߴ�VC3L[�}����mzh�7U�YHCd��~�"�l��(Ҁc�r�m��ke�o0��eUt��`m�E�g�������@Z�S�
]lv���%���t���}��NkW���7?Է��F�y���h�@r�����0ξ���$�*�RuKM1m�����j���8��wPy-A��9��_g":o!�n�����w�Z�[ʽ��3U� ��
�
d͝����/tw��3!��J�LV�݃L쿤^������7����8|^\e����� ����׬��-,b7-b���"3\��?U�%@��R��gD>��ua"z�RM=��@������?���}�:���Ym��4�;U�J��q�}!K�E���&��U4WI�_�&���Yj�
t-=�uϟ#Dg��3�k��O���z�$&�δ��d���b�Z�K��eHԋ`W�p��fs�~5�����͗� �'NOA���3u���)Y������� ���,V%�%(#����vҩ{t�����B}��Wbn�uAU⧃Ǚ�I��,���b�Y&u��?_kio��.2����b��Ѷĝ���u��V��P+�����"�&�I+wZ=����<0;��:�KaK���?R�3�B�����+��	�#���r>q�`�0/�3/{�u��WB�����8B����D�&߹\57>�4.����L�[��r��C�V��1��??\�T���
�~Rb��;d%G�_�(ʎ��t�=�# 2�K��k j��ޚ�H�5�C6��8�<�u3��P1o�x��h��$X�(�!DF&,�`G0{<{X
��P5�f_�wØm]Qa�L��'�T��%s`�3��Ø��I��9���X_��Cъ.�h�Gz_ݨ� K���dRc����(����xI�����8�tU>Y�Dż��VX+ђ����0
��4�1\̧[�;{Q/�a}}P��$
�����/�S��;��G#P0���-�������^�,3T ,�l�nh<��b��o���P���_^< K��B��X��.vٟOy�~��w�R�H듻W�,~�_ȂM���U��
�.�w*`�c�[�3C"��<\�O����%���i�����׌o4dh�q��r��d�sPǑ���WlS^#I��)~���%��J�Q�bՁ\U��QQ��qN*/"�04�ܙ	Cͨk�-B�(Ǝ>hn)
�\H8-P�қUX;�[3�~��p�Ҏ��`��B��'����q����a���Y�����'P��+��͘fiǵ��tt�f�Őmr�K��&�tA:�\	����r�(;��`��-���;�}���:�(
@0�d��9��[��w��Q���Ȯ��*���_�?���^���w/<���S���f�!&�p�U��$���mI�����)oq+��p;U�򳘭�pX���F�Y�n��!�'�ЦQ.!��l�j7�H�� PH��\���\E�Aw��]0l�Y���Ie�;ɳҫ��&&c�f �\։�d㔋b���Y:��[A
J�s��
�g]eV�������G�Qy���[�i�EM�y��1s��Z7�l��#b������}�U��qB ����Ɨ�t�|�)i4��UѴo����t������B M���ތc|o�fˍ	Z�Z��Y���ަ�Yꅻg�����{;l�'�Tj�`��� �]Tj?�=a�BΜ�':�`.�*��;HLz�> �>U��}.����E!uP�������H�텳�� �A��)ng/�뢆7�6�a�2�a���;�4�J�Ȏ�¤�[��C����N!PC߬D���ڏ���IF��Ӛ
��ٌ ĭ��L��>��g�"���88`ޖ�<C��.�df(�
%�@d*���n�b�!�