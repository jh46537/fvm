��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�&=�N���,^]9�O� �R�d��/=���H�/�~6R��2q["�2�*�\'`�y��To���N����"}Ԩ�-Y����Z�Y&%cA�'k���C�>�=].x�>~�ONU�4�,PI�ѓ���~ѕ�Z���rZ�DG3���}�+�}��{���޺H\�H�Ɣ6�2)�y?���'�n�A@��8�<�y:X������]h4�G�9
�����Ƽo���.ά�-x����m��ϛ耖c�Q#�/��O��{�7��(��n��WzT%")Lq&���L��?�{�A�/��|��l�Vm?ޘC7f�U��~VƊ���f����߃�GS��,y�<��yɹY(	��~��h%[�䙗d���_�����:�ر9ӎ�kGȘ����׮"�gun��)���g�͹#��k��Q���2��������S4�%H��F%T�MJ�=q
U��p��?2a�M���X�&y�[Qy=�\n�D�9�L0U���Ᏽ��1���"�r���sX�gO��Ϩ��~R��Q���L��h��.��֧.���>=�I�r�d/�-3Q��dY7�9{�����@���0�=F�?Gx�~��@�p@U}	��g�3K�N��.M ��n��E	�.��WY4�=�.-��isw�	/ۢSI��h ~���gi�b�,�<�b����!#f*���I�}۟8��7%.=��f�~��Nw�$PС8>4L�����x,V]�+�|��b��vn�S,��x��"�V�����M�&����d��cc�L��+!6ȜvM�A2�vz�:Rsx�:���i��Ի����M߽�)�5Z��T5����Z�+�f��5]�7%����X-��Mqc�٧�� �����Ώv_$ =lUg�0�|F��b���^�#J1-cتc�#�ܼ^����8i��¦O����{U��;G+��󫮙_�*k�	�H7͵�&�� ]���Y�<?����f��+�ŝ�HTLq#�{�WJ���u��hp�Jٽ�7��U*�L��߃�|R�#.n��K��G�Kg��	>��x��_&���n���;��6b^��pS?Z�=�h�jv�'ʱ�FB�`6�>I��+ӥ���p�)
�C�r�Gl�����?��nk�9�_8gS�)��A����T{���6i0[ mK�r3�Y���}�S�y)��i��lv��+�y��*�0_Q�!�>R���T�!Y�R�2�N�~�6�xZr�6=_a$�7jIug4@�]�J߻�CpmB��]�y��'�H3f>���׆�]����*h%��s��Q��x�+��YO��@>k��к�v-W���e��Y�ǂdH#����7���J��� �2�h�ݟ����ھMB�4������hF�j��呟U�l�S?��gw�&�)⋜j�;�FJ.g̟��.{^'%rf�� ¯���X3�z�	B/+el*"���
(1i��Wj���/K������=��1�vw|-yME��.��zI%ȟ�q,hUpY�/�c���& ����|ī�T�̬xa���e:w������L����#4�3��F}��vR&�m�A�Uc)���o)�	Y�m7@�pO�usʹs��2(���εF�0�r��zp�S�
C��Ϸ���ڌ��?�Y ��>�WǓ�.3]����h( H��gp����<4Ȧ���.��m�y�%�v�rKaY �S����s���Ä�^���F��N|6�^��,?Q�����^���z�&�q��+�l��Þ��D�a���ggo���7�>��f��_��3�d���Œ��( b��L��1|��%ڪ�-HZ�M�6�����"���x���B(ϋ&��K��=��2�uo�V�@�P�C�d��T�(M>�٤�#���cD%+}���A/�����������̎�����n���@����L��m��#f�h�PeM�Cy�:-5�k5c�M�� 
-B��'�
����z�$W���Û3�+~�l���)�Y�����Y���W�vJ�O}d6�o&dX�-���>�R�@ug�I'�_��fv��b��E��Y[7��u�;�|٩zRT�zc�è%��.K���wק�R9EC<���+���rRv��6�֯�h)*�Boh:u�:3�ӳT�q����I�M�՗
���K��{ek.��0�Ʋ���K�M���R����i7��+/�D��H�5#q���,�RB��5��VW��]��e��r�n�]�VjȤQ��t"mRf�@K���P���� *�1R���^1�d���:]Qi�Cz�Ǡ�����(���)5��ѣ*z�R��aN�v���4��*�P3 )H�c~]�=��ND2�+G�Bm�U�ܾ�t�[n��~D���{䎅*O}�B�(@�H�oWL��"y�p�[��)=��Q>��l�r��f���s_O� tE�_OX��Bxݸb�����T ~'�Q��з�	čY���>��I��;��G����l���������w��XN��^�%���J����Lp ��+�MЦGa�]߮�޲X?��N��%���E�ƞ�ud	�8� �b���|��S�i6ʃߡ4}p����TI�a��:��X�N֚C*�'���u�*���^Sz4��*M�i�Ȼ����}�x!%���'Ҧ�L����DJS��q/��=D��^���G���(���*q��6�D�~;H
�#��rK�W	Dlo��ߋPjO��(A���%:/�K_\f�U�(��&*������mG*�m��}Cޘ�@Ƥ�`�1<s�B�AY�;������'�J;0�4��Z�}�<�n�$�[~`7���V���������5��V�:���#�&�h>L{t��?J0p�Z�%[�uyK0�Ӫ�g��ѩ�c
Ð��K�����4k3I(���؂>�mJ|����-!�*A�W{���R�N���L����m�O]0?ɽ,�wk�|9��}d>�U��1>�ʪ1Z��F;;X��I?���ċ�����) mϕU̪������K���W� q{�t�x�P(9�O�-�k��
$ר=�׎O�E%#�u������u[5�l� �j�q�(���*oȏk?�S*7¾>3���
�H�o>2X}�> '��;;�X	�
<!v�eVf��9D���]�:o�`]_�2�$�l�4�����Ӆ�
t���Њ�&�r�b���ˡӥz��u���j���ۗ�B���?���S�Ow���e⩰N���v�U٭0�^O���Z�3� �*I���.�n����e�Tc,��y(�˔$2ӪI�܈�=���߬� Ļ�u���PU��9wC��f�t���۶�U�=Y�y��Yo`]��V������0�a�X0�O}���Q�;D?|��m��{,6�x��	����W����e��p�e�T�4��{MH)]�_�'���uA�i�d49�\3��[��h֩3���0<Ȱ-���`!��,N2l���<,���{�0�ugش��N��S��=��0����(?�"�a@���B� ޼�6�����c����ۍB������#A����!r�E�)��G_�qo���Z�a�9H��F���{�g�0hCټ��ꥭ@��t�V�+gi�b�U.��ʚ��ք�V�	��Hh�n�sn�����Ae��D-&Z��7�@+A��VfS�K�4lT�K-9`�x�3��0�����g�Tį�g�8��n��f>6�|A�8�lk7��>X�5�r��4�+�v��b���;�[�U�D�G�ǒ�0hzA��'�������5�(�Ht��<_*̫��0h~Y�����ԿY���壠`��I_x��K�d�8=m��f��.���zւ����炩Ff;џ3�Z����k��m�S�n��]�;c��yݟG;� �k���S�{S��[z#�c.� x�7]eN]:�x��:`/�H�[�lr`��z�v��;�>_�i�
�-k�ל|+ȴJ��u�Y_\`S����+�x���	��i��/�3w�Ӓ����g��DK1���� 2iyph��� F�f�)q�=�O�|�H�V�[����?����s��d$�����+e��+ŚO���"aL�6�?�)��劽<x�̆w��IgB��c��7�/����z��E��ԍ�B��i>�U�*��æ���=�����%�#a�J4��t���F������/���3$G�kNS<��t����@��,F�?_��_�M[ҭ�ɱ7��F0d�^,����W��7^�2�N[bhX6�I�A�.*��c1�>~�O�\��:�=鍀�l��N��@p*��U�:6�L]LlP �
�-%��0��$�ZzW��`�ړ[��B���Ǚ5�R�p�Fr�#��U�����.�:��"����[f�� ���Kx}�+��>�f��uρ�
,�� �ɫPӂ��m�F�k�OD'&w	��K��P�k&�5�M�����X�T��!���<�v�G���:R�zAHH�9'��a�l�3��X�7�2�=D:�)6f9 �tge= lk�BZ�k~�/���I�y�^��Ч�@6�Qs?*VY������.6)&�I��ȕ)	��Y7TZZ�Gd��3�����eM�jUD1B�o1}�t��� q���}�!d-�����g�*m��~���)�kwt&��$���=/S{������xװ1%�	��w�ؗ�oY=���%-2�C(eJ���JvX��إ$K��@�&�\����H����d���6�Ld	���*kI�Ƭ�������ǽi(��剛bx��RQ�u<6Ԓ���
��2;Os�V�K}H������/	S�������v����X1��P�$	w��v�t�e�)�L仗l��?��u|�:W&.�Q�ŨX�tj��n_/�)�a�L�:z�B����'
@�!D�����q��Q�=��������#�',�,������k���Nƒ�=�Ҟ�vK=��@r���*$���9@Zp�}��f��rЋtú�7�z� �N.ĕ����P$0���w�[p+C���#:&PEdp�,=�ꓼƘ#�T>Kj��jD�d3&�88�	��Pk^{�coX��[n�hyu��#��M��\�y/W+x����[�9��b����S�=�8ýtS�`K��o�#�O�K��xû��!`��";h�uʽ�w�z|��h���9;U��y*�P�|��~�a�Ϯ��ԣ���}��*���T�x̆�KM�d5QA��CM�o�ӪU�	��;�&%�xZ%�q��$U��
����TpF�o!g��-�)I'^�I/Y���QY�E�O��\99{���y�'�/p�A�'1��h�8y)D�z�n܂���2&��z�7�#�{s/���噟�2	Ǎ��I:{���ݴ�����o�,��q�9���p"=O*P���dg�����=&�IR� qz�- R��s���8�i��ܿ����-_��m�]�|K��(�(�n�!u����9�Q!F�=/��=Y-7/��c�̍IDC_�W��O\��f�"��	���oQ�؋j*q�����_�����%z��#0|����
I�$=�%e\����+is�2��
���M���*Yt�?0�#}���l���nَ�Z���1��H4���w�H���/2$��
��� �N�	� q< wB�M(�5gE��>sP��K/�f�ÜYJ��o�R��@޼ӎ�,޼'�n���/v�8͚�ǳ�(����oX�h�UfhJS�������@q��	�^�Bn�ﳡ�b�i��V���/�C��b'���Fl���8# y����������ZZ!A`��ӡpݮ�ˋ[|:!K#G����h�~藭�(l}�R�=�5���4�Gj���"ڑ���.Ֆ�u+��q<�}��P֐-��	�[��hG{�I<�A��ߺGX&uA�����p�c5����"��9T8ʔ��-����ѻe���\Sprs"��1�`ň��敜��dݕ���(Ӌ���M3���Y�>��~����N��o�*��oXõ�'�V�E�CK1�A�/�/�Ѫ�;�_$T�И���{��l#8��p+K��4
��ҧ�өl�·�}+�YQ�J�՘v�F߿J���Qh�#9s	*��?��+�BD��Y��b��W�6"a�/cq�1 �$1�jY�U�8����ƨ��"�%���_�X�}�PНxNF��I������h�X��n�g��,�GJ�a
C��"gF�d}>�5kXp��Z=��EGg���h���}D����A�X�o���tR�?�H�����t����j{�;��Vߒڎ5=u���_�J�%�^H���H�š��_`�v{zg�N��H�a����{�
�)�@�5����%+��uMD�i��aV&���?�������h�7f�FA���2�h�ϳ���.��˷�x��x',l��DN��*4J�S2�ѫ+v6�R8r*�w-��X;�t�BR�d��8w�v���K��!;L2��2�jGp�}��=�"QO#��z�rC!�mI��%9��)�B�C���5�Ċ���*%w�꟏��U��%�g�ǆ��b��q�e�>�.��t���O�܁�G�b2�񪥕�SV�=�#ʖ���1 �8�>S�e��ٯ��1�����ċ���:]%NI���:Y���!�ř}-��4đ\�+�#&}�n�������z��Ĥ����6�ɻV��7h��B�^�2^~L�Bd{ʟN�V��'p�X7�T<[L�`'[uε�;6�nA�4I[�f�}��|�����*����q��ƣ�x�g���	��~h'�ʚ0�l��� ��Z�_���!5�>�=Ul�L�$�V@<oX�r�t0qqK�%��n�4�P�P�6hrۻ�Ʌ*Й���g4�%<"���EƉ�i�x��c�ϓm�g=4�w��XJ���V8��b���1�m�챘.f�|�I'QG��qx,�H�q��]��A�,�>��dd��_˽���/@;`����b"(d߹�-X��i#�U�^�ΐ�$E�t ㄾH�~j���X��>���25�+	�6�}�Ae�����?�+�.�k�3Zb��\�
���'�w�l�vX^I�s9��75+ͩ��r0��0h�)�g,bU�y��y�-���8`��a��#��Z��H�m}i,�tLi�Xj�b9̧c����g=,龓sb��#�(�����j��?����B�@�,�����)�Wh���X7��xqUTjK3(��zL{�UF��޾B�Ղ��tk��_	?�ffQ	=�5�}!�3���� ��-B�M����$2�L3g`��na���t���p�)���8r������Zƙ� 9��I�P�`4���]�X\��L���8'G��Ħ'��Ң�F�z��Cr�DUXf+=ڷv�+z��a���dh��͹���ރ��x�_Q���?�8* �����!d�#����h�AҶ"e!^0�='�I�k�K+ڴ��"����	ٝQ8Yt~>�2�p~ ���g���U��2-^1������J�hŷN�+��|s�w��r�v�)�b���) �����Ҡ���F�"	��^:J1����9-0լ��D���9t��^���{�i9+��?������V�~�L\���9��n�m4&��� ��腍����>M������Bg�JN��ӻ����1���s��l����'1� ��/��&%-�m����* ~puB^k@�oˊ�+�ȇn)�����-�C$*�79;����젫Q���QY��
)+H������
�dD�Σ5��!�� �@���ϲI����U�h�����]�k}0�oS��&� '�
:	�J�̟\i��R}0���fB�w��k��qc����R.��=N�m�Jpd�\�Q�݇�Ye�!�h^6H.���7��U���
�A{=�H,��*1�^�٫>>}#��K��;u�m��Ņx<g�m�ov`ٝwj�}��6�/�D�-@�+�|�S������3_�iT"��#��Y-���D�������oD�`[�r�J�J�N�n4���Xr����G�#�b��O��5��r9S��c�`�n��m,X�&���ڊBOy��@-�"�w!&�K=m��j}1�	,P����_aőX$��.;��#�d����ή�z���&@���tlE�Eh�\J��Eݓ����T���0��a���N��XM�J�ϒ��X�4���r8� �ɪ��ؚ������b�|�����.�rIy�;�Y�]�i��M������*��*ٍ�	P,'YYM|�K8���@���{e�Ǡ 	��wGR�zn�K�Py�E�Hq)^���_J�����/4)�!L!�W�i�g�.���]�m���?|�pk Ȍ�e�#%B�P}m�[��jq���a��p�����h��8�xd���g�[C.�X�mCvr%ẩ/T��p7?U%���6h�.��ܰ�<��u1r)7S�J���F�6�HgSMד�2.��b�Y����J���7�Aމ���v˖�,���T9�����(�xnzU����t��.�E�Ψ֒�	17V�� 	R�����jڂ�3��hp �s`��z⊑5U�Iv��Jd1��`�ׇ�6�Y@�IY˭�n>�vG��z��k�%�'@��N���F�w;x�XO����s�g1�p�>w|,��(}��37����0�E��d���Ĝ�3�ۃXW�ɜ������.$��[���O��s���-R0�r	����Q�䅺R4�`�1e�.��K��LV①�o��^z�l?֦xh���t����x��G�w`�E�)��9ht�T��`��E.��ВI�4�X�bB�Ƨ�c�"Yl7S=�펙+�J������������m;:�j�d��I�����|z�/��������f����_�K�U/��R����(�\>��)\��Y���Aaܨ5�d���L3���/f1s�Z~ѺFz=�wW��pS�a6P�ir��{��|�)l ���<.����kT
Z�2�\����1oU�5
)o����t s�Sţ]{ғU�/�od\K�]H!�!�a���2�͕B��#��#>�Q��=:��9B�O �ͧ�����uڄӏף&������˗�v�A��zq����aw�,�Q5Rk*�qv�,@���=�hQF䷽Fwߝ��S���'�V�6A��~)������+ga�(��0��Vs�3�{B���Vu���+B���h��������E"�܄�ڧ�$���J���c&ճ�Cq� �P3�T��D쪊�NA�ob��	�Lv!�#��fk󒖴�WH���j<�0�o�?`^�'K�ڡͲ-Ay��E0DR{���c?��?�5����C��\�P�jT�!ٟk��q�9��S2��Yl���#�]�����#���uG5�j�e� �oen�{��	@�xW⺔�:?�Y3�X�����	�x�4��JW�y��`�j��&���0�VH���K7�o1_�Y�T} ,���[�h�Ϣ��u7�P�s���W߶8��\������*�O�U5�X"a���xdt����6wߦ�`KH~׸{����E���Z�W��p�fǲxr�Z��Z0?sC+�C����7
n����`_���8��o�6�l? ��n�T��N/�J
��.>����� x�|[���Q�J�[�P�Q��B�V4pw�m'n�տԛ��Rr%P���^bQ�2-3r��&_��H�~s|�;�P2���l�j���n
iXm����&�7���.��P��e�^�E�v�(흧xYT	�s��S�ēe�uX{dZr}o�p5r��?!�ľ�� ���g�UWQo�Q�0���4���4�>�Х[�kͼm#�1%�N+B�ڸa�SK��رy����Aaक�րǲxyI�h7����E��tclh>j`��(��zP8M������3v�cgH�Sf����^��)O�GF�:�u��H�����H-��.��l{Ϋ�|8�$����L�i�vl?�!��6e���k��f����8���>p�ċ����Y����w����X�(��	t��	??{|�r��^ж�2ʵ���<��@�b�s4kו�Fh�[��Z=o�S�x�t3�W>�V_����[���*C�WC���/���8z�8e�55����'�w]Y�.¹�������i�RL��C|�
R
 y��"R�ڿA�@�Si�Z�uE�������/���Y�?z&4��vѻ�5`�k��P�1�{Jh*�T�Q��p�f]�C����[�d�74��#�A1O/2��M�'�1�C`��r�J�.��Xl.��X�~t�6r1ᔺ�����G � ��A�:�P��u���ru�����,4���o�f���᜴b;7)��<���h�Z�ӍDڱ9(M�$�Gqo��*����	��`	i�.w^�x�J	���2������̖�Y��G���������rNQ�9���T��-�*�MCU7�H�2�A]䌧Ǚ�;�H����Ĥ5�?wE��"�Cgڈ��/� �:�H�M	FX^�
�o��xz�lmXuD�}�}:Ʒ�{� `���1>�����?}~Y�����:�71٠S��`� ���4�O`X蠿�����3�;z���0~R��&��ͣ�G���8g���! (�zpT�) ��囉��t1�3�҈���tPX?ȼ��@� �?}@ُ��� G�%㠴���&�W@�n'O�Z͟@����!�M�$F]�P_���n�tKg���&V�^kz��f�״��-����.�wn�3���&��?W��W^?a�%vj�S�H��G�Rʱ�>���#���HN�@�Q���(�C��"�"�ռ�~��`;�K�	v,�����\����=� ��	<�c�_X�K��?�Y&���¾"(�'�C�r�uK����?:� ��<�^K=�ͨ+�)۲�;�J�b$�߶}�ix��mFZR��I�8������0�5�bX�*���1V�s\��U��;B`m!�)WL�u�1���?a����)�*bͨ�M!|6��5�*� %�/��}@��i�.����@A��1�H�M�6�L����Cpr��~�z
����{�[��l�KAK&�C�����RC��+&���a��5�K ?��*��H=�����ȁT��ZB
�.XW�Ш�
V���H\r�XU}T��n�v𜑔%�-��$l���ޏ:iOj��m��.},���}������Q۸��T>T_��,�{�$��'��ª�=���"�n�*��K��3��A,�'|k�ox��&:��0E-
�����[��io�YK���E�gB���4H��cH��V�����V��u���5�VA���Y�1���ldK-[��~z���M:���[�Ύ�Q��yc@�A�XgR4�P��ͺ�%��7��X�-L�X��%�HC]n0�Z���+��ߺ4~���چ�D>��oG&j-%�:]`��-y�	Ҙ������m�f�̳e�1e�S�� %�^�xȗD�`�O�oք��XK�!"!8���\�л� ��L��m�N" �䗸+qF#� �R����jB���]��l�޹z���S�"��(~aV��g��[	Y�=�&�z��^ڢ���V�a�1ceUv���v����w2�P[���j�15�,��p�Н)�s�/i�H"¹䑷�%"C���u�@��
1#���4��R��k�N-�R���榷��Lx�4���A���!"�6^a6�Ri�3��,�=������[,0��Tm5��%�q0�{��U�ء�=E�}���H��A��e@� �����@LD�2��x�4��������ϕ;�L>�nl@���J,�W��"�	�������h^�VLs�����O��ֺ�j�f�~�0��߄�����X3R��M�\��Ѥ��f1�	ZU@�:QE+�6w�3���_)\K*�Ԇ�_9�R;�`�ȑ�KeKD@��[hMI5f�`:���BDB��W�e$��]�m�ؾK�Zmk�U����Ik�T$4����==|����sƯ�J��hler_ φ���C����O��"9��J�q�����tw"	CL���E΍,i�Z����'�F5��n����R���/d`<ih�#����3§��NVؕO_��`��l���{8�h;q���#�Cn�M����Ƨ|{��GS�c�����V��Ӛ���aiW	k(i�� ���(y�,�Z�@��+5v�驲��sg��vE�D��<
B�ӭ���9�*�\lG��za.ouc����`8��mZ��0� ���ic��}�=���u�YQ