��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}���
�,=����ڳ���7�kF��oݫޘ�$�?k�
�MJ��Q ���q؄=�|����!N��і��v��RD��"e�/m7�mY����p ��֑L�3�׌FaӦ��,ߝ�>��a+�=q�{	�T�|3K�:�*�{�����`�SKE�U%k���a��!^��*���H��9�g�g��ᷰ9:�����j�FƤ�lB�9�c�E8�o�ݴ�'%���7�ܴu-$r2G����o^����3Y��G��Ff���n�m�
%�y��ȩ8���{�r���ط~�U/�r` �$?A�@Y������e��=�Pߑ�
f��zB�$��SL�������������e�2ճ梬�� ��\�4tT����??n��nʸ׻I"b�ŕ} �I�
��8�M�_aX3��;�@�yuDx\��o�a���T�[6+v�a�d�R�P�K���\��sEP���ҳ��_�H
oݸ���=�=�+I��q[b6h�5ݚy�f>�T�BN߬��$�m�t�t��f8X�J;k�)wq44��BTG�(���]�П�o�T/���%+$5xDZDoT?P�!Zy�7:q��h�����̊d��3,S��h5�:��jtt�gw�x�����%A�Vs�o?�TO۴�rd��U�D����7[������3�K����i��y�aj~�ښ�թ�*,�C�"�s�'�T��~��.3�+�V�ϑ�}G˕���#~��N*>f�~/��(�%Ev v���e���%l��8�h7�4����HllঃS�u��C,*�bOV����O��������Z/�'f�n=g�]iU
�G�|��?�4������W_*[��ũ�N�����(�)�f�̶ăy���'&>M���H�O 5HQ'�������v �T+�r@$^��?!�����0|	/��*J���(so\'�)��`�L�!|	B�&G�0ò�����~I�5C4�O��E�ik�?����]!3�	y��4[9�6MAآ���Y��CAr�����-���p��D�3�A��B���	���bS�;�s��b����̔',<*�GG��&�#.aO;�Y�O���?���x4O=���#��n�\z|$K�^�Cz�.��\����!������+e�*3�wy��������A2l)
����
�7]s��KR�EI����B���x2TS��vՙL�#'uK��C�g���sm�L�<h-�:���k����F]�{!���7"*6}J�,�t��?>m���m��d�b�-���+��>�H��7�_�O�I� 8��jVUrn�h�LM�|�iN6�to����|�v����gL�ED|��{����3�:��Z����m����!̶?*���qDb����՛H��++';Bڕ���q�9�5�NBN����mZ�����z�X����Q�� 83;�iT3�]�ж�wp��y���KB��1��Ʌ�ڤ����8P�N��VN�y+Bsd憁	VIb���Ӟ�E_�dx��9���K��9>�񮚶��N$]�8�IGM+ED�л=3�"�G� �ݎlG�����K3���qR,U� �gL�L�����]l�|���t�J���v���
�D��l&�IJ����\.�rR��K��T�i���4Ĳ�F��K7��B�u�҃��xO���^5���ڬ*���?��o�o�lka+!bI%�!��3v�p���YK��Xi�X~�	�?I���LM�±��X���z��1�	:�kuO�ړ�����(2�=�<�����1N�f�w~����F�"�[�*�Z̑H�B��|A�js7�Y�����o���U!*���ݨ�\ ��N���������Ai�> �MedɁ�e{����4�a��u�E�S�("X@��H�����Y-"���Y��W%���:�f@��X<H�;�/�Y�И��g�����]Ӷ��,���ME%ў#6�b�V�˾j����S,r�c1�+�� 	9&ӟ�	:UA><^�z���O%�;hIM	������Eb<�k..�x��L���̸��q:�X*���f��[ YS>"� ���
�z��e6�[���x���1ד�zAd^�o��ʭ�g�9��D��$\	�h���iY�E2��t䮾�T��e(���[/����Cm?�CٚR�����ʸU�CGK2vWޏ�)>�'�K��tq��N���h�6�,�4�A\�m<��� eM�Y�W�yB��msE�Z:	�S �Z:}�Q��ſ����D or�[��V���b��W��<�xt [�w���m+p���s��X2�/m�x�ۍkT��C�e���5)�yO��Km-o�q���p�������
ۋ�����B
a-v�d��<&2S`y��(�����6Ol��5���}���g7������T�K��S�m��V|&ﴇ-n�X[�0xd�,��H���fȏ$���~N���^�y�Jg�ϮU	*���Y�p����.��S�;cB�-��݁Z�1���c�y��X�ƪ�^&谗��c�;n�b���p^$�=�H�5�,7�d	a�OI	���"���H�qdkD:d�]���rwY�����(7�j)"���<Ҧd��P[uFpk���F�<�%3�^�S�
����
�ar�6#
�5�|����Q���f'9�m�Z�!��w�ŒK�T�BU!��yW>�C�|��OC(s�z�I$LOuU�"�k��_�v0q�E��5Pr�����\ӊ�r�o���(R>BBY��b:�qg�!Y$�\�G�{K�q��;F�����x��������w�R���忖��œ��Y\4BS4fũ�4��� ����4��z� ��H��N�/���o���h/�.�ɮ�D���M_=1k�Ea���mo�CL���1�O�kf�H�V����Y)�q�S�f�n7�%��v�5{��܃&�W��� �aHe�G�Z4-oCU)o֚��փ���$'�rd�tA� �H�Z��U�HX���L���O��C4+24�ޙ2s9�M;�*)�����<dy6@����\y2�-˰�������Q��6��;��#E�sQ�i����������v����&�R���@�Gg$AK�hĊ��M��̣K4��\�.�RW�����ȸ]%K�(���.`u3(q ���4g«�h	����ƟuX�����Џ#�2�Z���&;�7dB�>m�D&��3�F�rrU�f�}AV&�Z���U�\����*�R�����
�y��tr�}��*��i �gO�43I��SZ�:�����Ug#��R�2k��A�eg��O��u_�E�e)굮yC6��Y|V�b�&G�ֽ�'�N�~f3��L��VU�)t�Ԅ��5����۷��H��z�Ki���[='�d@�ۻ�E`K7�:x�ѱB��X�xi߅m��"��.c�-�ӧz�
�D�{��Ó>+:d�5cG�> rꗒ�p��*��Fޙ1l����G�?��S~��j%֭��0���GJ깖$�����g��E��C��$���6\��0h=¤�����*��en�[�%5���&z@eo�]�ڕ��9��7n�-:U&��"i^��>y����?X2	�$M�dHUn@�ؗ��@�����&�hg,zg"�K�}~�_.!L^�0̏��5�#׋:�W&�5.��
�p�_L�w����:Y?�?��/n���A(k����!���w�4C�͙Ou�asO*�ޔ��`���p�w�V0!��k㈒e�־��R��%��
����&r�a�+��y����^��ar��54N�/�����;
�ˠX�m�Mm_p�7Z혂�f�P_b��מ����d�E[�9.C�t�Qz8�팻�<����E;Skm����{�Z��r��Vb�gm�e�`�2v��ۋNL�k�$�C'��߉z�n�M v����J��%�	1��*�V��բcf��X��4�-��:҄��hD�# �����	!�b0��)vb�/��S�#�`p?��B��L�� ��[��"i.���%�U��o�0��v|>=�5�wVa�kMC�@=�L�Vn���Hb��
��.$r�{��&/ls�߬O�`�
�9�ȵ�hv��ґ���YnN?f��_��b[�[y����[�D:@abګe��(�;Ԯ2��`O~�&��L<(�t�y߈���MZ� g��(�� )�cϞ�t���˺�M�t�x-�U��d,��Q8/~\F�M$�$ް������Ջ������xf���0S&5�v��DO��Z���Ҁ�y�o}�S���2��MS(���~���lb�>ek	�d.օS[��
��	G[j��$���nT��=pp1(���ǭ�J� L�';�C�(_^@"P�?��q�cv�!�7d�6"�F�f
ǘ���Y�,��P/�V�w%���c)�vu{_������#6�"þL)R� L�*i�z�c ޞй��&��ou{�>+W�Sgoi�>�����yU!�$!���}:Os�q++>"Y ���z �k��(��.f�/�����q�!�PUi^imX�c���,]_ؿ!��z���Q	^��"�/Z�G��CK� �MI�O�X4$P����ex�n�1�M�q�nBc���:ѐ�ם,��)�YPpG�P_o)Ȕ�^��6۷	��K��<�O�6.�}�w$��H�W�@m���ic�X�<���0��ұ���_�zu2N�\3(N��loq���j:B����"�R�ي:�A����IA��N�@Qǌ�S��`�:��ƴJB�7�<2�Mv[��-B�8W�+�a�C��ly����q���j �r��(
����ͣ�ucy�*P�E����)��]D��&p�\-U���>-�[IWw9\�������ΌpG�6U�F?}�i�_�/�L�YYx<�8�����_��t@��hS���@��T~n�o󼆷m���b�s��G�^Wh�X��NN�c
��9�=�KG�1PT�Ȯ�|�:l��q���BL��E�!%!}C$s��b�맚��Ca:�C*���"��F�Y��M�3���S�^rȀ+5�����dB�u̼z����{,�ZktJ�B�	J;n���|��s��>�i��tй���˛1z�����/�,�#�I�����=�"�ci|��N�T�CF6��1K���"�,�<�Ɂl>&7�j�=�������<��Y ���ى�� ;�m�7��i������T'������Cmg�%Im=jC9��-m�?�4��K9��!�8k�Y�����j0�G��b�I	EZg��;d'�`vI9���|�t-��+6?��V�vI�H���!*�0w�P+�b�	�eߕ,fn��'��[{�ڛ���� ھ`<�G닚�:)-"��w70�Vvf�����BB��DmP3[�Yg�I�l��K���G���W��	�!+����˭.%��-2��1��oR��z�H��QO]΄V��A�j~l�r�U
q�GT�*����j-!F�l�@
����(o$V@��!��H�뤪0J3�x,�%t���'��HF��b���x��:�!��y$L��(�	rg)a7Lj�4�����]���p�[��/��;������U��_x"�0�[����Y7s�x<9��B�,�
Z`	��d�Q>�)Z���Ș�H{EG���|�������B��Dá��7o�E��g�?j�w������֌V⏋[��G�j��]�e�D��T���]i�Mmz�h,���O��]%�e�%�P�g�9�Oc�+3�9���&Y{b�Gt?��s��v�Z��D^WK��!f]&?���胫${v�.t��F�hL]�CF����uC�[���z�
}`@�4���lc��1�H�Sƴi��'	� ��)l&��Qb���dl�7L���3g�s)g���D��w��[�d9O��C�C�бD��X�V
��	�v����-��k�A�U|�ܠ�T�t���<��Ѿ��[X-}�2!nrǻ�6�8�"3����V���}�R��3��LΗ%`bo6��K��W���P��H���#���fbX��i�\Bd�z}I����V�O���5���e*W�B�AX���.����֧v�1�^��Jq�V�v��j�}��Y_nO�X4�'pڲZxG������y.���<"m��� ����y��'�x}�28-	C}\Ɉ���c�� �� \�cS��q���6�BD�ߞ$:��f\�[1=^t����&�!D��2���/�s���(H�Ͽ�C$<����8/1�,Z��u����aƖ��*���+�1.߲��`�iY��,���O�2�.�٣�V���`�a��п�4˹;��~����=��O���]���1����E\
	7o��:�4 �̄������n�2}r:�R�O��>�k;��/�m_Ti��p����2��B��~�΃I/(�ACI�:j��:�.������un^��)\U��%;��A�U�gE����\A:�	P�������j�3T�|0G,�؛qR�����/��q���P��H(P�sP>�0�Bּ��I٘G#qɒ��YW�i��g�JL�q�.ս���Ga�� �o.3���|�����t�a3�a��h�o
Nf��$�9��rq��ws��&�R(l�\Nc*D��Y����Ď%w�٣�+�h+`��i�2���p�ǔ �s�	�H��?�}��b)�XA��,�$|�%OQ\Rl7�V��Ư�6���_z��/B�h��)�r������v��Y�e�j\�[^7�E#����:.�J����	=�[��G�s4rү�/�\nP��s��Z@KL��ˍ9H�W��U Ҡ]���J�H���f�g���v�W�`��q�����V.��3��[����I6�@���:��nP!�heٺb������A �o�"X�2�ep���8t$�m���� ��EGv��g ��x�h���>�y��&ݴ3���fu���{��޺���_F�ͧ撑�bc��I�?B��=9� �M��\)�:Rų��;:�u��:m��u"��n� ��<�^{% 2-@4=- ��a��\Ǩ�x!��d[�	w�mkV)`��t0 ���o�j+����>����U|��M���i	��i���f��o����2��$k��*�-%tx�r�`�$��\Gҫ�-]к{�XR�޻�=(�=���;�/*I�m���QfXDƋ	��Cʢ�����HӓEZNv�,�>����o�Pvv���w��*��x�:�?O7Kg��2���s� ���������/�uP6�;�6��kF��b-���m��I,n@Ua���jPǙ���=�ŁM�W�Cdmd~X-�ÿ�i^G���&�ڥ����\�'\��%�i��g�pv��7lE ���+~��dbe�c��XZ�bN��Hu���.��sd�z�l���8�!�MR^;��dHq�fY��O����UTO���,#��E��Z���t�WpgY�&�nuKaB���28ƖF�/��o�f�߇��&���U~���w��qmEQ%����s���Ԛ��E4�we�ې2d"� Zu���n�LN�iB�x�R�����<�bi�'%�`�,tUA��#�2,?�4�H� �\�3lVh ]O�CI�z�7�&38N�&Z�2}Ht'��s&��j�w@�NԤ�K6�����J�y���L؎�].jPs!V�۵G�~g㊖�ؿ��Q����DFqR������g� ��[���(얛�D�1wu觴��OQ�e>wjxM��
L榻D)���^�̶m�o�9z�"��o�nV����Y1��
� 1+�/�p~��{�G*�,U�<�����o��n$�AP�WE*y�G�\�j������iyG������ڈ�G�"���x� ZP��&��Ej��DM��.>��#+ -E+����<D^Ռ*�p��z�ы�ߏ�y&�w+�2/��`�x�Ӹ���	.u���q�&N�R�?I�x�s啃��>�����@/���+9F�������p�Pq'��`XX���w�N��'5�γY��n\�L(����7�����:��%�W�l�ʧ�|�7F��\�\Bl�54~�^f�q
l��l�����6�_3�-�0Oō09�MO�˟^�;7����WC�d��C�s���h�+�8<K�F"�^�� ��q��H������a�$��*����{��\܃�VS��iŅ�������[LB�5׀/�3��yƥ�(g��ų�ͣ;Ļ�m>��q��#����m;UW�m��$}�p}��O��I.x���9I ۼ˒J��	�y�#:�>���YS���h	NA���O� 
���5�ُ�Ƙ��HDޒ������ɫ�x�Nq�p �!O6�2��M@��T�s��tUV{�dw����y���N5��~7�ks�a�&�k�,͑%���lL��[�R
ՇO�����ْ��=Yo��pW,��Gt��~�,�V�5��f_]��~�*e[��fz�*~���f��RI{�Di}4���>M��1" LC�FLx�>@yϡ\�_�n�I���<P�@7���_�`���?o�V�|��0 &�(�U��4�j'%�)��e�n�͝���I#X	��뾱c*]C�1b�k�N399�/�Â��Z�5i{E����s`��1�^~��Uhf���O���iQ=��Q�`��%Y�Da���'��*H��Q�S��r<�-a �z�`89_v[!���#��ēgTηk������:�%"9n(���MY���C�P&�yh�,ѻ,���/Wc�ku����E��~tF�c�'��?�(OVyC��9�9{���<��7)�����č+�f<5'���iJ��j�a��Σޑ����hSj�#�{u}��C�>��i�b��Wʖ|�л!��y7U����Lu���a���gM�Hɴ�HD�������Haf ի�?Op�0��\P8���
n���t.;*00�ƜaR�&��="�q�O�U��8���с�����q�Oń0���"���5(r_�=�B#lKf�=�#i3�U���Le���FG�?�6�����p5����^۹q/��H#�V6�g
�wi]3�ۭ��IG)@�Z)��K��g�&Xjݩ�˂���E��oB��Ar�E/�"^��
�T���dQ�f��,��k����u|��`�3���_J 7���j��tX❁}/i�NZ�VRah��N����o����	'���@v6�@���U��1M��u�)�����YC�W�S�zz�oO��̨��lb�UN����%����(G:u��9��O8wv��(+��㴱&b��ӂ�o�����Ҙ�~�����xex��(��4'a^�l
$�Kjg���pA_Ҍ���ɥ<k1�DcS�$�~Y��8���F-��$��jI�[����s�Dٗp�4� оS0ĸ��T�u0o������XW��Z?t�-sU�E����$܌CFN�]����Ϩ�c�>Vw�(����%�͋�ʨ�����U��忡,+O�'�0t��-tc��Qc��?
z�ւO�[�n�w�|����-l��%)�����A��D��3F٘a����$�����A$�qZ�>k/���	��wP��+ ,�8r�u���7�$'c�*��Ewq�ӥ!�ǔ5z��C���8�~�Ϥr|�!o���1E����hm����]���Q�$k�D�W�r%�?�XU�|vI)c}��+3��b��^�Z)�ix��dwy�H��O��f#����#�h��)�����!I1���X2���i��p��0��]_�:���!;���ȡT�\p3�eK_E��Ģ2��w���xU�J'��{:��F` ����V�M=��y�>�G1K8K��UJ���l�O7s��٤�k:��ߤ���������:��?�Yd*]���=Fi]����/_@�E��ղ���B3*D��r��v��d+�]��ѯ���:G��;�*yڕ=�Uc���Ú�1���s�.�b%��O��֋�X��FF�IĖ�P�Gzn.��d;�� ���8�ls������5β�w�I����rc��,0���`�o�p6�+i���+F� �͒�y~�@-�ϊǅ)?�.n�p:2�z҉j���Ӱ<��6/�'�@�HƠ?���#hO
��Lu�����D��=���v�d�j�52\�Zױ3�髐ϕ��]8�k��q7�1Y��j����o�k��8�s��O�J|�C�u�M
-��q*�v�7�B�'��8�i�d�L�]j��5N斾��CT�r)H�.E��µź��qBwTHځ�h ���?��)�%���v�m;l_xmTG ���RB%_��y�=��Q	���o+ȳ�����o�/���u�xɌ����r��i )7��ՠ
�.P�4g ��Ü���w�ȉ�*����s�����^Ӈ��)6<]�|����Ɠ�hu�J]�WI�_��ADp�����w��#��b�#�7�q���l�hS}D��^�(�����i��U�mQ�=K��蔝~ϯ�g���#�#\�t�AݟO�A��[5s�^��F�3o^ִR]i�h"x����	�'��Y(��,̖F�I.8�ڜ�-�-G�-���]lfaE.A1B�M��^��0��2;�騌�%:�aYn^hCE�q��_2Xz���5t��E?�^
�	����+���;�x-�;�����4  {�d.eC�G�=D&Xh(��#��:.4���%6:��\��F��#��ts%Smj*:s�f�ϟ0i�z�
5��ō惒G{�a����X����i�M[�������z��O�w��`fH�r�R�~eu��E?9���8�־=,�*�Y�����X�����6�q��9��2O��,Ka��n����� ��0e�?�F�$%ջ�Mr�8��=��.���!��
�6��Ϟ$YR��F|���UԻ�yx�aM���������=v�Ua� x|�J�3w����E��&��'�l���bb�fU n�<�B���L��d�i�iu��C��1����Q�7�R*y ��l}�×z��Q�jQ5�LP�:�lp��A�������#�r�L�h�2^C:���u'�c<���C���J�G�d�s��y��F%���*v����8���O$_�y!���Fj�y�\��e�:�b��Q�B6�Qk��ۇ��,��A;{{X������^~m_��QQ�����'�_M�H��y��a�5�a�Yu֞
^��A�!���[y!�z����	��6H��`Sk%棈�h�x�� ���� �Sf��M�6��"�↲�®l� x��~e9��s�R{Ó}C��#m@bp�.�H�g��g�	�=��$��m,kn�ז�}�
�(�o����B�����"
��W�u�f��Q�
k�Z1|~%D�h�%��;�/LP�P3l�Jo�:	��'W]�=9��|�%�}Q�G�(*��H#CG�7P�^�O�?�HJ;�3�^PCY42y!�>���u�d㭡���H�b~�^-�i���*8��%OiXXb����n�	u6v������?�Ew�����~%�������y|fXp����R1���}s��?1�Qf���"J�塙E�����>�R5��ֺ�o��`~D��"�.Ɔ'�2Au\�(�f������`��k�Ĩ�*�s��;&�X2��Q��2��uQ�DR;��qc�V��:V�L����PO����N���ɾ9�5��g�������-���D��>*��{�C�K݊�Q��>�G�rh({w\�o�ޜ�'M�]��ݰ����ag�'����>ϲ4��S��?�3k���Q�[>I���x\��.����8��h�>,�U��Y m�[~����i���#_��̼�^"����'�][x,�R��Eh}"�b�{U:@����ک�nUBQ�,:�dS�ǻ4��{dU�J���2"
܃?���XV�E\=���m�p�ҫO�Mmz��&�S�����c�h~��*�"�P+��w\l{@�m ��d_�_Ȁ���KI�}�����X���1��w���*1�d��(F1�W!��Gr�1>�j$X��w�2q��#�0`و�=�k����M����Bہވ/"��l��*	Jb;�F�V����0e.��3j uX[���{u�̓2k
1Q�?hn�@���a�\v�6"cqG����]I��I���'y�ɯ�'E)64�U(,��[�{�x2e<�VC闫���󌛆Rʇ��sL���J���||RI�j9�����'�����R�eyg>�Q�I �<�-�N�B��n�jqF���		���y'1�-�\�N�Q�1p
�Oy1:�1An��(����)���������p����G!�9��!\�l�	E��ց����h�A�7�~k��y�R �#tb���<�&�Km��9l�Zi�Q��f��y%���怰3�+��Y-�S9U�o"䦉����O�؂B���Y�d�H�L,e$ͫ+�_B��_V!B$R���Ȧ�8�G�=�b��3���$ �P���n�3�`F��r�h9cC	�j��Aj�z��+�w�� oRo�fyYw������E��Y���ǳ#�rw0g׋�bsI��Ia��j��+,���T[�(?�ۻ��-�cP<�\"?��߻��8��y�s��џ�~w ��7I��G�]7�wۤť!�]
ok���+j.ah!Q����?C+�����,�2=KO�L�S���@6q�쏊��i�uQ���f�P^��:�7L&̓H�S�MkQ�W�:Eƿ
�N��.��_��~��s��P�'��(�Ε��w�0x	�R�ߪ��9/�sQ���$�i��0�}E�yw��<�'��L�G�i5][���K��&U���6sF����޵���D�4*��NR�^�S�+�*�"ŁI�����[���@���HK�����{Ps����9{�^��9"� ��Wږ�ѕ20,�0�$�q�:�<|��"(:X����O�$v�m~jUݔr s�������H�4�'���g� K�����;L���6�q��$�
?��M�0-�X���zD����k����J�S�/��xb�:=���e����.WE���"B+������Z`���d �rYk�E[��6x=e�%��ZZ����mPB(��/R��� �dL�
LrM��� c8���E�
�]0�2L^���tF�R��8=u�EQ4o�� &�DT+j��Fkm=��<���ϡ�֊X.�-�xrY�1W]�2�\�t��1�Pd�Hh��%�e�gnxX���*�����@��U�uM��M�
��[Xp�"C��m���XPS3H�3Ǆ�a�,�%)1�E��u=�y63]C�B���U�Hy�M���1�u`!G�a$c���2������i���h��y��TѹafQ�at�]g���� �h��f�-`��<�F.��*����&O��P/���c��M*\�|�c� uWu��3Da��:J,ߚS�`��� �*�k��2��IJ;	%4�J��0U�w���\���[��~"IU�Z��� �����Lu���ٓ��O.F��ُ���J�BX>>�g�x_d�g#!*(�i�m�7)�{�ҟ�UK�ţ��{�lL���+�*�O��eO� q��a\#�Q���s��X9L<Rͻ��(K�IA?����v@�+�p�Y���4�@�ia��h�i�{��NY@k1H�7�6�3��z��5��'��1�GϬ����wҟ��P�0�ڙ����&u���q1B��D�i���_�A�;]Y�(=_o�=����n��Tbߗv&�r���+E�z��]$�qE��9�����qy�hJ�B�^�z����Ǭ$�]2Kݐ���@ǉ�$b@�R/����Y�Ƒ���ɀw%��ixL�ۨ�ꫯ4��1�"�oM�W��	�B�:НDK��5@�ԁk�9��A��b�{r2�,�<^�ߎ���Q'{ҿ"r(��BB��R���͆2᧬�|lD��L��M�ܘ���ysm�M���*��t;��m�6W]e�1��a�C_k�k�BK�ʅ�ш���>K����V����Ab�c�-���>�ߡ��¹�%�k�

����by�x�~��T%���R*�n17���!�|��_�U&R=5��G��A�*�_���H��VF'� �C��~��Q�g��t"j
I�5�Wg��
��7�:�F�v��)�	©g���H�"�)�V�چ{���/�ht��{;��-$ޚw�	yѳN�q��& 8'�8�Q����}��Ī�F )�U�;�ߨ�`_����C�>��r|�>�S�uE�N��A/G�ż ��~ּ���ΰ�L֙]M���zM��S"lkM*���ƴ�=.�?�a~�T12�i��Pm%q��ґp�b�.G�U��&�6?y��Oǫ��w XM���op�H*�־�R���X���f�V��P!�<�d�(�����ku����7ui�n�^�ǆ�*Na��RG��ze��5c��@����A<=��@��_*-_���[�=H�M{�~��j���q��]��N��'ɺbQ�����f�dفal���h	xb���r�]�C������0��6 =����,9��_;��7Ԁ�Gq�����T\f�<��q�y�`[SK�؅�{5���6��Rь�4Jk���P��
����Kq�C�߮��A]�=6o�K�K�9���F��������<6NbjM�i�~�����|�ج�g��Ȥu}a�JJ�Q򐘐3�]��&�J��sEo��v�*rd�v�Y�o����
��>��lq��h�ɦYR�آ�½Y"B%i�}o'q�J)Cܞ��u�h�a��IQ�����HIitV�`ν�$�g��c ��B<m8��������!gW��>5��1XЁ]��\���Q��Wh!�з���'�n�-Q**��BCT�VoNŵKV�'�;�s@�Y@r�߃���td4����	)�O�´��[���NA#L�(�R��Mҗ��_D��F��-��/ؓ�0iX�]`��=9����/mA�~m ��+���JMr]h�5���)��y�NY� �k|ݗ����QZ}�--���]�`�6P�W�ӽ�
㟥��~r�Q������OT�)ڮ
�4Rt��B��!�d�l�a�n����R��rQ>�$���o��{����z�4�BK�r�I\uׁb�e���\A"X�2�&)B6|�Z�̿����D����W�f����]��}�m���U��f�h�� ���
���P�*�i���(`R�n�ط�ď�7�W�z]�u\)�;�z�3$�d�����ä�6�:�K(R�-��$@Q-�����=p�y$���ҧEٻ$mKͥB�����!Os���OY�-4�3�i*T,b�jP��(�����s��qv,�3t>T��#��� "�!�z��p�x��z�*#�%������ �-�6{�iK�M�����U��ԁ@tS��'�w������,��|i<��F�6��lm�d:`^�����0c@Ē����5Am�n��r4�'�S�Ps����\)ʋ�+4g@�y�Ǌ�?�ת����m���3�,����r�]��p�ژ�Eֺ_���Bk��^�jK���n�L���WI�Qr�@p׀���b-Ek��_�jdz����so�׼��]��~pF�"h�'���O	8���z�73`�PR�md���b�˝IV�.e'Q���=Sz��vL�@���L�.��\�GԱ5ej7,��R|\a�{�Q�T�#���o����{�Ź��8�#�B�A"�9��$��k
ɣ��=s'����s���ϰ�{�/�%�T6���W�R�ر&M��=x�+%�J�A�������Ϋ�N+�\�:��4VK�A�������B���|�9��CB�%�u�M^�f���m�|<���'+G H{�T��M����AS��PѺ�{C���s�Z��a�\��"_{�}����P����dC���טxΗ��_�[�3����0:w�D7)@C	O�g�ga��"p���AB�M�>��_�%��jJ��-6R���A���g�W��j�%��p���" ����d5��1���I�$/x��u��Z���r£�� �)�r�m_����&!����6�-�V���Qxc���V��D<��� Ճ�^�5XF��MT�g�Y���Z��RM�%��.��%�y�8=7��6���q	8��R�Zc�:��a��U��?��Mg�g���.�T3���NY/0�c�'�G�
8+�;���9W? �~��"��+o��f�F�;�
�9�����M� G�i{x��|s�����o;�]d=�1(b�_�6�W$0h�D�W�_2
����D��A���S��Oit��<���QkJ�S����A�� ����qpY��2E���k3��	�z��P�|�TG�f1�_�/Զ��������u��~��'�t%���>�E��Z%�l*֧�8���d��䴩֡U�
Sz_G��U��,X�ŝ3>�ހ��Э��D7+l8���Ox�\g;�5�f�-U�`���ɇ��oL��׹��A��=�0�ɒ,T0~?���u�X��z��i�˥T�B�h�B�,��v��*ؤi E �k��)k4'�x����?L������A:�n���o�ӊ�&M2�1�؎���)pzd5��=9�����y�A:Y�b'��L(�oc]�&�(�l��>�o�>	{�%u#?��H�]%d!r��u�.3uh>5O5���)0��q�k�yミ/�yu�b�fv����<Х5J�1 U�	W��wR[m�>��u���0z[A���wd����c(��O�p-%u�_t��q%4�� �6�Uٿ�W��ld~���Y�rx��+t�J��g����N���ܖW�[���袹��G�d�w��3�;�R�	vMJ��_���M����ϫѓ	U-�+r�-���dɬ���	��2:�+~��pH�(�u}w-���u΃i�z���9B�~�}����f!&�x:��?���o����5�`�|�2JG�5X��U���������'ZE�y��Np�\c����D߱�/ ֤�{w'����o�cXRh�����x.~R�G�
7y7E�Ԩ�wxh�DtrVѝDx��X���e d������kڅG0�Ey�J�I;A$�r���<����蓻*-��P!�^%�_]�,���Ua�O��#Rػ0h�DY*��y��O����}A ��2uX8ϐh7�s7�Ͱ�L�)��J�UP�ީ\Ǣ���7��)�G�U=]�H7�jke��	�ͱ��©�Kl�#����k�j1q������l���X$\��7]���ý17�Ӣ�G;]���-��|�m��țu�<�-��y���cO%GΦ�_�)��I�8԰���q�J�ǧWl����Xo-+�]L����@nZ��LT���L|�W����XS�9K�� ��?�!����ȋ��L`]�����:tI�Z�����Ǌ��pT����ߡ4�x㝲��#������y�^��3�O�q���� ��/����C#���a�S�������=6��M����v.�*���#1�����Oo���5�����h��:�!�;`K�m����Hڒ�5���4:5e� ڵ=Mj�]��D\�4�z�䏬��BhPvtr�fʹ|����p���;q`+ƪ�)|l�67,���?a����v�)##��/��L�t�&�w�W.�_&��oZ<G5w��t\��S7Ch�V�&�al��0z��ʑ�I���]��P�T�/��lVm�DԱ�nⰠX�b��6t;�7D�@7|>p��}�'bœ�\�
5�pG�#,2Z�[��+]!�,Q�Qu��sP�;W���S=~Sِd척���'k&(���&��0M@���ر7���H�7�_YB�Gů$���Cq��^�B�m�O�o�GExV�5� (�߈=<b!;�k&��ᑂ=�;3sqP3��L�h�ưb,nHUU� ),u��C.�+~����PWհ7j�ʹ!�T��"�hY�$
��'Y�1���q��f�yÐ}�}�g؜Z������S~�ポ��<k`�$�; T�{i2��id��	����K1W�2��B��V�jVsD��*BR-��bb�L�GM��&$���$�zKdr��B���eה�j�x�����(��i{P{ҲUBx��O�ɒ��E �v�FT:Ƅ�֜�K��-�Z"Pt�s�����]6%I!��ٚ����<�(&�o�8;m��lz��JA��{wqt]��A�ay�Q(%L��PS/�ּ�_����d����Li����3g߭��~&m�a*�ࠏ2���}����y=�ua
<2�����w�D�Q����O�+^�)�12�U�%���L2M��iɦw���s$�rΛ+^�ꄼ��*7����͵f?������{�,Ө:�y�ը���F���x{�\8Wu�Jr� �p1TBJqD�S�W�Du��FQ������y��_���m��9�R� A���F s^ǋnD����:ZIckEϰ�W`!{�9ih��n�F�7 �"�i ��e咄L)ט�6�<W<�6�,����>O�.Ȳ�ZB����V�|GH�Ծ�ڄ�_ݲwzt�*�Zf;ح���T+o� �}䘔���#$����\�w����8�o�EA�����<w�����	A��Kx�VK4�)�����f#��酜!��OM�R�Q4���NlĨ K�mk�z�~�� �݊X��M<θx��]���vA�O\�xnN
���^���]E�֋�J&T�٨��!�Sqs~�R��Q��1�(Qab�bU�4�R�����b'�}�r���3.)1�'�zڴ3��}�� �P��7��`Ҧ��jC���pE� �#!(����5�;)����I�9w��e���]/ҳ�}�,���������"�J�<����� 5T3g���V"}���si�Jv�1�D.�&{�RI�c��7��FS_�/p|&H\¨a2�f�kv��Om+B~MjփД\�6�q%��$��I�OgB��MV��Ka���ipX2N.�����T������Pc���{a�ƪ)"�u�F�,Y�!Ic�}d�&w!��7Rz�Ah)'rll/��+B�ě�0�����NOE+�*1;?�?��p]A.|�J%��8��|���5=A��G��*����E��x[�V��!�mj��{���-*�G�4�"*@N�v��d0[2'N�(K�@&kp���Z�#�E_�������w��T�f6o���qMڳ|����`s�s����]&�{���y��bث=S�\ O^�]���l	9�Sg~�Z�P�i�My�"����1�c>��(��[�2N^kTM=_�����~����e6q���)�cW���f�Ð�b�:�*ᕐ���	?Ym�xÁ6A�v6��T�7��� @N}����@{u_�o`��g@��(uʝ���f��)��[ ����kgR1���$�̽|�5���bv�?%��{P���(__}�_��Q���y$o���+t�V	L��㕖�8�!�1�
�x<<����B43E#��^��j��1t������H��ʁ5p�>Z����e�Ή;��fQb�ځ�;s��0��>
���k���܄��ټ����@[j9�ۙ�\?�An�d%�m��3�4=�J�n�/�=�`�v=�D��.(�AM��v�H�]Åɟ-7yP�L<`����X[��TE;btd���;CZO|=�C�e�,A~򖾓M#Z<�U�I�ʤ;�w��~NY�7&z�������'����I�*���m�>�nF�M�}�X.����C���
��b��?�m��~��uX�V^xZ��� n���2�s���1���dí{��!�w$[��>J��ڕ� ��?��onMX���%��1�9ma�̎U>��T��Жl�l��-QuT�����<]v"�%�Bqߧ�^�~)m�:���}�Vw��>�Hpz1r����u1o�n��K���
������1��|0.�½�R����� �Ef7�@UHrpf���zZ��0�rr�z=Zw���x41Y�v�$Ƣ��oq���^���<u�h��B}h�m��%��%hB�:�E)�D���$���*������`T&���X�<�����s~�'ӬP2�ה�D�p�j{.�t$؂��?L�Il@L��'L[�k ~����#T�M� ���\ J�a;>^�?�[2�#�w�pv6�4�k�ĳ(Ǐ']~�yk�|�膔�k�r���?"��X������V:��ҲQ���{.'�s�����]F�����������t&�[���2j+�gDT��po���h�������j�>߸cV[
`-'Ds9�-"�L��V�]�N�����Ln��?�Ǹ���A�鄽Vލ���ԧ�F����d����j�׬��G挜�rp:�yݮb�v�U���̧��i#8_��u"K �#u���xg�~X\%R"=G0k�:p�,yE�!�L�Lݴ���)��Z^����`��=����z	ڗ��V�-���DI��S�zj,/f���(�O����LH�s�a�>�u����|�1�m�����W�_��M��5�����J�S}۪@��@d|K���!	�q����� 
�D�@8�/�K�b��c��R>�� #����?T݉�HR���������؍=5�3`�rQHli�D��'�}��-��e�������s#0R �Χx@PKZ#Ɠ�#�1���,�7��7�lM��i�(٭��i�C��Y�*���B#<�e�(~�7�1�9'�=���1_�"Q���˄c�sa�o�ę��y�6R���ee4[ Ԝ�RY����������%R0<�f�Y6�$<��I�ɭ$�y_�d׋Ƒk���0���>s~|�"�}	T.q�A���w:��������\ �Sp~e���aG����:���s��f��j8��P�������>h�v�����d��-$5ae�/��@-}��G0FcA|�M�4�$h���#
�ۑ�<�C�~��FI�ߠ�>�9�P�61�i��%5�c�/�Q� ����E���K������ۉNBiZ��D���@`�����W�e�i�?É7}��U��uFx Q���"�F��,	��\Z�⻢��c�}�eG�<?�r��H��'E�$^��� ��Y`9����q���a��5�{�8�Pz�ڝ)9���F�@�X�?'���_�։��ե�s����4'؇T=�{z)���=�_�{������(�+\W�1֨Ʃ[��Oſ.�9��atI4L,��)^h�Vkr&��$x
�7�d�`�k����X�Z�g�߅���O�RbO����Keڧ���=9P���	s�a[M���%΂b0������/a����kC�2�4 s��g���~Z� w ��I�7Қ�����(7u�2H���95R=�2N�1��K���ˬ"���h~o� ����)�%j�����DO
i �Ka:��������s�E.��b�����AF�-/6C h��N>i�꼊��nZ�[��m"���Jτd^�aѺ�Fy��ڍxuټny���@6_�c��-*J������&o\��/�.Ą«�u9����.�"�g��p�D֕��Vi�|����pW��a�z�B]z�Cm�ο}���<�o��<��ɔo���:�z�4Z�Pϓ����(�	\ϲ�:[<�}v�?-��M1aU:?��sa��8r�!��� ��p�(��i�1I���,�&B��vY���ԝ�)Q��6�1v�����ξ���Ě���!�ܮ�	$h���#�և׮��DZYhXΙp�*���*�]���8eb���aR�1�޴"�P)`�S <kXj�Ƿ�^T�E B+�:�0Ե?����/�� �c_:J�yp��V���31����rm�'�����m�r�s�p�dl�"�3w�Y���o����(��]Yz
��i��tF���A�dQ
���\�6{�:/͗[���d�q��_��/+U걀X�jX��6A2R9+Q�����d�4*@��1��`DՇ�V�u��4V)��
�݉��5����R�G[$JsӠs�Ӣ��,$�����BG�8�%=�fmlbxM�$��wbN��.D�SH�cN@�UZ�������IRB��aЌ�U����ֿ�#��p$�d?2#ja5b����H�{WM��#s���z(���D�9�aNJ3}C�;$�mzr�"K:B��g~�%@F�dOv�/����E?�T���a$��&�	?Pg�X�����@?\��dᅕ�1��,7@pk����*���k0��_��e�4s�MTg���^�o2����W�G�����O��� �/�o�R"��n\��ɓND#���i�2]r#��'�q���i1���C��?���*��D�	��>ٽ���c��'9o�8�Zz�
�V��y�{�8�7(��.L�QK�_�՝Rn D��4F.�y�g�$����.*�?(�����i����|L��]�3�k<;��C�Wk��\I-����_m�<[��O�-�s5c��q��|#��n��/��7�U�ƴ?Z#g���<%�)>F{  �����N��n�,��}/�m2�n5���&�H��s!<�
�������٤;��?��5j�zJ[��M������Fk����@��!^v���hNS�Dh&\�dW��c�Õ�4$�)�+I���?�	�M����eF���ף�՜[��]�Ȝ{'��V����������c�'��V�O6�6ͻC�',��4�bƁ�3�{��+����}�bT����⪀=*�������3s� �wBu�_�N�@9 ׽'"^�,q�Xc�c��+��c�h,#���x�@h6E�:PWȰ ;9nҗps����� �ë��lh)����_��=����Crz��7�0}��@��-2vP x�p��X�^S���@!��I,��R]8�����2ǷIv�[Cq��?(CZ�������� =�ZI��$�(�\�S�+q��_��f|���D�c�PwA�Fw�$SP��kD/x�s�-H|C(�o��B�e	+�2���x�c
���d(������I
}�/��OƂ9��-Qc�`�;-[1����p��s��<�A��� ��s%��:�}��.�c�[ф��R:�=�1�Y�?��e�
��ՆFA]b~���[�b)l9���?��ؘc�`�a� ���$N���2�m��G�'�G��h�,��MXP���,>��X��_<�5%�S�k�p7�U����J��,/��QҪ,�����m$.hցo(�DdXE` ��y��8�a?9�L��>r�[� ��<�E�����y]�4�c?0*!�~b��`�i�G�X��g�X����'�C~ g��0Kk���W�=���XZ�ͭ�}�W��I��ˑ���k�a�J�=���D׹��
M��f:�:����o�1x0-���5�^���N�#gA�0 I�η �&�΃����$�lq^xA����Cv7�|���PC�hM|��q�ێ:N�,j�t�ca
��fr���ǤO�
�0	O����F����Ztfx�E�`t>����W_��z��N��cŬ^�RWx̠���m q�&U �!s/�v����x9�sT�s猠,2���z��*[���wn!+��]�/P/$P������n���4O`�~00��>O�4/{J�I�,���5X$�n(�c�启l*ڧA���i�ծ[SBq%��b��:8����;Vy�eam XZ'E�.7���-Gy���-k��gg�
g`f;����~{����ͻ��Z������Wট���tyaO���rXm4�W�
;R�Y���y,�D�D`�֨n���!M��������J����Y�P03�-H胡�=\�N�g��L{�
`�R6�S���K�/ש��;�]�A+J{&��.���Lǥ�nv/�I���1��p�QX�^[�0lp����H�Z�)�E�6w��#�	,]^ .`���u'P�� �(wā�7�W�{a�&��t� z�VkC���C�ϔ�L���ى���v������x����2s.�S� �+�r��t{��c�dCfYQ�	�Ѽ�1�-�s~���+�3�	�pZ�>&�t�{�v)h����Șe�"���.&�K~��~ y6�N�����1t������0L��u,7���͙��6W.��vS���<��40�������:�z>%v@1�����C���)��6����qkG��CItX�e��?���|�,�	"�aҷ�O�|R��������pc���F�����|���@�����gc���b���� �B��Y�`{��j�yS�Q��5�����#�cBg��A�0^5#�Q��d�� T���=�8C��M�������3��Ӎ����.�sՎd� ����3*�>.]D�ÿ� �odjw�Kb"ETo�r f���gt��,��(�$�GhiP���Ȟ�}:�͔:�H!��5p�N��&D�%.;`a�8�@������7�Z���L�	0�ꓶ�n�¹
?̰^N�&��Q���G�$$���� ���8%�^%
������������1y���/�A�NOXq^X.&�7+��"r޽>�cS�~�rq��~�8���zJ�4�@���lD����u�aa��~-���qʔÙϾ���a�#�0Vqў���X�?|��P�lc�w�!����<������l���U���5�� "
�`j�c+Ӧ+(VP3�1�?\do�D	t��^vLC���/&_O��]BY�V\��`�-6�H�J����\E]J��ߺ��|'�c�(��(T�C�"}[��Ts���;���&��E��A�.F��|�Z�?�d)bLmLD!s�o���I6�2�f�ۘ�@:@B�m;�C�9��\N0�N� t�70��o�a��'Rܶ���~��͘��vK��_\4�ǧ"��zX7 �C쏂��?G�殼����2�JL�LINz���N0��fW����G>B3r�2��ك���)qO�i�bꊯ�;���@�$�逰c�=� �ۤ�'���Ld�u���j���]�q�?����l�Ra����X�)d��։_1W4J{��A��u�:wc�Y����+#���|�:杝�y4�D�T~dN�2ӭ �������^�V��0"�k�n���|V��-:U����IҘ��)I��j]Ĕb^Y���G��W/�t�WHd(��1ܥuӾ%�M�r��,�R|Ջ(�a-� o�W��z)v>�e�3�eɒ���ˏw��h~jш�L� �V����;�'����x
,������.z�^mR�1��ٔ���)&4z����i�� �?�yy\�F,L�B}��8�I��[~����\��8��"�B�s�2����ʦ��2H�\���w�HL���t��<,�ڋ�CW�{�������F����\�5,�ގ�+�v�)B�!esyq�����i�s���#�Y���e�iuS��e�3�D�=�\Y�,h��kT���W�uRb"~T+�i՞d��ւ�z����	V�Ӈ�����۫$7IMX>-[u���T��h�
B��Ų��s�`pe� <	���AqNV�w3��r�j���a�3�d�m9&��������.�"e�]��<�#���z�Ƭb����#Dy�1𡟚fe8FR+�ġ z�ЍY�;���/RQG鎤i�F��4]��7|�.�P2Vs��oǷ?hҦ^�[+�:(
R�%C�UV��*����7��r%�\����$���J��Wf� ��^��� ���^o�`EKGw��Q����Y�D�V�xp����ө��(����T�Q'U]���O�.�a5���|���O��b��s�6�1���z_>�[�x��
*~y$q�.���ݫ���9i�\�"�e}��d])|C�}p%H't�$�/�HUD��%�>��	m4������U�0�3-}�^�a}�?:4���*~�9��j/>X������c����bc`#sU_��X��	bN���s/0Nfx�_��&��@�>�5�{���T���8�}��`i �_�C����s�2�ɬ8�
��x���'�s�)bU_?�Vn:��0���NZwֺ=�3�6k��:�%�9Fł^.y-�D��I�)���B#���#o �Erq�WSr�kfҜ���U�[Qbz�>�De��&��D�hqh�f*�H�k�	���]���
��q��\����8��so#��ژY.c@7�U��� :��k��Q^j��F{�R�Ӊ�hP�k�U#��;�n�@���%DJ6y���(�و�1k�ކ�i��q7��B}��g7,�}��M�@�8K&��������IL�>hBK���$��Y�c|A�{���
���WŲGU��%ө7�$e���*�}�z?3V����lb���9k ��'h�bu�W���<`gTWV|�h
�Km8��q���BP� l3��:�� )yZ��"��p|p �I-�H�a����~7�hxHg�>X�ĜUV�E��{���1@8����Vƾ���X���
ˣcq*���:m���������S��e~#�퀶�3s]A ���o�_�����k��;yǒ�����c��N����ǻCg��q
��FLo�^|�!�2�-X���w"<�h����^������'T��ȁ��,�^�n�b�W	���@�Q�������`��>��,���?%������g]���7QeH�I�N���Rz��
�}����MhI5Z� �f�̣�a��Zc$��4���0N��q�Y�OM�����%֤J��e*�Gi�@`���*YA~�,�a�Vb����ї�BN{�ҵ��u8��2쮇3��H��	�w�H��b�)��aݿ4��uWR5��~v5�`-H�Ey�U��}���p�
YH�nI��^ϟ�����L�6���us�)������4��p�Y��a��n@��8�v��-ǂJ�l׎��|��<�.�Ī�R���V�˘�h�?,�kh)'�^4�hL�_�UQf�O}8�)�~3��#%�24�@��h���%�4X�t0��+��|�O�Ʃ��T���L��:XX��p�	w��a ��>ޜ:�01/��S#�Sr�1طc�2�'-�{U�Q��61f`C�{B�����KA�rB����H`V|~�@���DD�$Ԡ�E�q��KP�A3x��E��^��,yR������9e���0�<r��=��c����w/���Ջ�@�3@}f��̈VV�[�i�"��~�S������w~ly���t��m푭�ij;+�ŷ�n��sd��tV�1e��l(�qb���M{�\a̳��3�͈o�àR	��.ƌ�י90�� �2�������`�H*��N��P��#�DU|.i�|k8�2d�4�i�Q��������Z���ʱK��D���cȶ�'��K�[*��U�F�3�|\���2o��a�����2r@��`�4�0�TE��݄L�2V�����%�����Ջ�]M��,j��8
n=Sd.�2q_�?3�Tw���|�w����*0��v`c�H'g������u!�#�|�jG&�=��	#��n�M�e"�($���H���<�SK63=�"���ظ��ǸNF���xI��8����pa��_\��)j�|���\����@R_P┨ӗڍJ (�ϟ�y�qJ�D�T�We��v�aJN-�_��_n��=&��[3DW?���28���bW�����]�fC�M�ηt�R��4�����Ԟ_r1�nھW�2�����+�`�XE����?��l�/�T�z62�%�6/e/�1[���%j�Cq}��{��c����K�Xu�aX��U"l�����A����'1s��}n ��W���P���b�c�=�_đ���r��
UK��5i}�c�uA����J0�i1��H628�[��K^Ww~����;ā��a���#@�!��w��{�����n��`��_q	z����{�$�1q�,x�vN/����ۅ�(�k���B�����TF-���j���1��'��:1�������R�N_Խ����Q�XF�icWd��!�*I��>x�^��d�o���^q�2)��+��.�W�l�f�ݹZA��:ӥ�|� �����I��˧،�y�(uw�\H�q{Dᕺ����ӳ8�M)�~x�j��Â���B�7�"s���X�[����K[�����e�/�`v�_,+�����A5A��(HN��g�T���e=����Ь�}'e�7�����V�1��#i#��-�.�[�k��?�x,��"R�t���P�<����,�BlD�y �F�l�4�؅%>I@Ik�8pM,��d@ω� ��g��8�1�̀�Lه!�&h�>��ʜQ1�3���~��|+�wUlX����Z��"T�z�@����i�$�-��u*�Ȥ�v���x�߅ʔk�Q��dnani�Ƈ���2�#M>~,��~��hp����=���q���S\��ϔ�7�.?Ւ�I+��n�g{h�#�m������O���S}�Bd#�oF��z�iٚ^�Y&�N̆��8�zI�L����$q��M�U�T��=���ȑ��� %�r�	�s�jx4�U��^����w�>ֱ�Cp#�kk�6��j�gMbr�l�%�&�\�z"?"�Rj��Lɑ6ޫ|�JW�.��QD$s�~<P�I:	��،Y�����v�B������Op���ڛ^�.����p�����;��녾�:y�_�ۜ
,�3ˡ��;(џ����#~����M������'�~rp}ƫ�3O`>�8��_mN����.�K[����<�~��)��h'v#2�nq��h������a#�C��bx�_�
x���u�