��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z��6��5��g��P��^�d��54�k�I�d6\ N�RF�N��>��;d�R}dG;��A���x%BI��HL���p}1_�dc��hV�HHA�y�c{�9��1��Oy�Q��A���1��&��1E��W�X�[�
F�Ɛ�- :�X�QՋW \�ؔ����)1T�zuê��k�똌ʇ%����ۭaϔ���KU�Q�mԦ�+�*��Y/�5�H�^���8���z�J�^�6/�m�+M�&��f+�>�T�<�ۚz�*pI�ܢ�vq�%5c�7���:պg,N|�{�B{qF�@�EI�m�t@�}!Q���,���<�t�����}*�r�s%��M�u�V�3��Y�N̘ҋqY�aqF	�Y<�LN��[`:�A�
%��X]��6ꓻ�5R������&��7��QY�=Y�l��K���� �o)f���m��XKn�f6�i٧���L;���o�U�ũv9�r�{�ȫ�I�gN�й�Q�Sz�2��HyçV��5�L��Yw`�$��/[]��N�&�*��2���̰��"�d���A�! �����Sk���i��I�Ԇ���0���h�I���4C;���m���W"���ԯ���9)�˫3'=T�	�S,��u�3l ���^Z�I��D)��@REe��<�zs\rGЀ?�%&OHx�����%�1v�����'�D��(+�;1�Ї����|$9��~A%�o��r���9 �\Ξ�r��3�+w�����Q�vfV��I+�/��o��u�'FU;>�.4�I�T����,0�:g����C���������X�QΫ�÷mq	/^����b��y���^A/���af�l:���|.�d���ɴ��r	���͙���E� ��ܵ�x@���
T��^�\�Oߺ� ���Z*�H���`L G�&)k]��iI��(��@w���4�-����`c@oX�~v`��7ۻ�[kz��Ӫ�jÇ\�::��Om*��[�&��D�lt�ڢG���R�cL�l19�EC��x�&��XU0� -j&Ԝ�t�1��L��b��Q��Ž�oaMIO.!�[�,W=d�nLS^u;p��b�^jW2�<��6�Y⊶+:sLc"�I�Hi�0*��n�uR\pI4�i��A�8�!�uD#>���w�ρ6�Z�~KWQ�]�oL���ջK��b�#e��ɻ�f/�
	�¼
;n�6p��ϖ��4tڨd�nO����̂���[=���]�Sʰك���@���� q;��ߜ=�3�^�J�z���Ϥv��f�$i��V�*(�x��ш��#�@N��
�~����r�|�0�ɴ�Y�?
n�8jW&S~yd�z���&�ε��t�*���I�"YO�3
&@��e��Nnp�8b /�Z��Ocg�m�'�6d����UL -
���ɶ.ǤiD��s��k�:��i�O���r�S��K��yJ�� �����S�T���;���G���G:���:�=Ŀ���F��S��)��0'c�����rK�JlȽZM�6��i.�O|�S{��I�꨸&��?�
j"_`P�^��؃/ѬPS�:Ƥ
�'oܹ��	��J�L>w��G��E~�ͬ-��9��\Kq,���Măw��q{I����:J��Pƕ�n��220?�U�A3^��~{%�-��"��L��}h\7�.�����˺����]�k�|��;��.��J��y�F�{޷.] ����<�;AYk6�,��:���7	�ܤ2Iλ��hm<�<��.q� �%���F��3 .Y0�v�y��Cx�{��w?;��B=����A�Q3��2�b5?�TP�$�[	�ژ�9F�5���`ߋ�c�[�����G�6�F$�(�B4�f�7҆4�ɏWBދ+�[�njԛ�����ߔ0�W��ѯ�6�;�!�#Յ�|2n@5aA?�#��B��8:1;]��
v&�WVD�p~�dj���̵�Z~G�V���%��`��}�[1 ++I���9:.SG�P%��:ؾ�x���Ӫ�m���T��;��iO�Vy�J�b^�ۅ��f'���*ne��(D�[���*ƕy��������h�>�|�u�v�!��n�&��;��i�;�WQri쒭Rz�ttN�k�%0vk��l׻;r�ނM�}kƽ1�� ��2��ctv��j�������s��/� ��+�S�?#�k'�p����")Z����C\�cG��֎����Dlh�s߫\���E~^�����;!�E�ȇ��9�҂v%�)]�Ʒ�_��D�lR$dLle�0���vD���nr������C��k���"@�gg��}ފ�8!�v�)��X쳳������֑!Ҋr1�Q���}#�JT�Tn7��}��]�E�;�� �7ch�@�z��a�I���rc��{��W�Ge?ڥ�uf��Ӆ��Z��RN�I�&����6�+�P	��7$FJ�����_e��������������$T���0x�a,>�3d�3(�v�<�!�7Y�H��7d��AH�7��o���ڮ�f��o�k�n�����b��'j�c��N�v3S��a�fW\^��Wy(eGI�|�=�~36[���#+m�sHC�L�x�L]��f�L-��A}�w��u����y�"'����
�p���z���_�}~h��I��WE�Ζ����\�0�[�C�hKz�����U��*p�����p	���j��<�u���5Gte�t�4�خ�}J}�(�Q�yZ7P��>T���q�L~�ŧ�!͵�:"U��=��)����d�}p���$^��1��u�[�\�c�G�,�OQׄ}�_w�R�'���Ҝ\��9���WR?�3�V��K��|����C�]�$���$�ܴ��#@�@��X>h%h̤�x Nb^�ō��I���y�#�h׋�1���5��w���n��B6�j#4�旱�-�<����Ќ��8��~���\�/b�1��Ż}3��:N"�j�{�ZK~ـ�m���A���h��7
βE��^�	����c飜m��Dr�S���$:�c8O��e��������[v��w6�82�H+����q��J<��k1�5Hu_���^����':ǫ�4���QqSe����Q}`N��TI�z`��/"�,���Y���s���7r�x�>ą��`dڃÑp��\��أ���Ҥ����a2L���fxY�%�x�.ѣ?��E��<d}�f��,��T���a�������eIh�����%�wb��k��o���� ��mP2/�!	���<L�4��8Y[���F�A}ߪ��Q����]�;�;_��`|����u�$���]���G���<SPT��I��o��'8F�W�F0�C������ej~�� �6���WO�pm'7�ZF�%���GP����*��8'}�����ޯ���u�����y%m���g7;���Ϩle�ގ����	v��7����|��hR���I��W�~�KX�e��
)EJ_�YA�^��rq<=�n�9�H]���P��h�Mo���X0�BOK�q�Lr�δA8{�L�@�£t���[��K聇t�������W@�>kS�!b�]�$��΋�N;OR��5�+
�?�Z
C�u�K0�x��I>�ƭ(����޻��|2�^��UQ^�"v�q�b��^��m��> ����,��L���z��d��A7��	9S��=�3��j�\���@��)fx�~�\��]��E�����i��X�)'�|����X�$�<:��S)kv�;�[�� ;��^Ď� �Y���`N�L�2�:F��\������E@�1��a�na��jB��"�9&q���`��xE�7��r�L'
��H 8�����B��:Z[x�@�'��A�5�	p����?8ؑ2`�nDgM<-|E/b6p+�I�����9����ԙ*������{㱞�W��20F�Ҽ��k�qS���^y���'�ϸ� m��Z�"� E��&����S�����ꀗ3�(f���y䰴���\�L�bGe����D�̸
��R{fx�'Zj��`r�{d>��/�xI[{�m͡�Y`tJ�4���c.BS��Р����%�|c#���4�#�_t�km^*�r���J{�~~�R3�H��y� =,�w �)�Xwc�u8 �8�9�b�x�Evw�Ǟ�$T��6�7�΋�o)2Q�6��C<�^�S"�I����h%����*��H8�|��+!N���V�a�T97��z�IZԳzX��+t��r[�<n�!�`;8�3�8cQ4�6�R�#����b���4�&<�zB������2g�<O`�aL_����Z	�23k�R^w���F��4A+�E7L �idT��ڬ�67�u����`��%�:�KDhH�[3�KU	q�9 ��� }�;���|��p#ʎ9��ʖ�p*_pK��SBiS�]YnIl�Z�|�E�5�B	�k�o�	��bĻQ

�ʬiD7���g�(X�_��klFUݯ0�#q���_,�����[�9��;d���P�O����C�{[��'b��q��Q�ֶcV�Ñ�h��)�j��Z�_:%�l��ML�B$��ԴD�V6c���;mN�*����F�v��l����A9�����A�7�9�2��Ha�u頻���8Z�zb)<�������9d�{���PU3A	�htF��f�U���"���I45�����eH��fk)R�Z��~b3���R�=mj��n\�Pd]H�4�}R�	>����ǌ;,�#>U��L���YCIi1�]�{jm@c�rX}������%�@<aM)c\6�[Q�;�V`i�JMN�J��e�z�� � 'O��-�I\�l�R�hq�4l)�s/�-h�,K�'G��r��_��}Q>�E��[>�@O��2BǕ�l�)�j-����<��H|FR�.�.x�S��JQ};u\�����;��C��uEEl^�(�q)�V۷�2Z�{YBj̭3���1��gY	wm�/�f��� w����c�sP��4i�.͆�N�ȫ�{�"X��눥#2͓��)��-� �=@��zo�-�%��
�U�+���Y#�<�Im��z^����NS'/���|���w}��=2��rѡ�`�X<�g�����p0���Q��5H���'T7�!�In��k���y�l�z�"y�i
5�Yl�Z�]��: =��Zug�s]���5r�"�SL����e݂�d�j��7�0|�ZZG�kx·���L��P����ɐ� �Հ6�1�W�j-�ӲhE�.�����Z�T���g=��pR���tѬ��ds�$�\�=x��Lq\��6�R���
�w&� �(��x	1%�ŗT40�Ҥk�-��Kï��^sHD�%�iK�͑<�v���̿��ox����H�|���{���c7>xo��u���So��AQ�ȅ.��v�#�<����,�z�wp�!:��\d��%a"�}�{a��Ӧ_�ע�F��eBp��<�)�����&�u֕�v���၁'/?��+��r�~s�2ӿ$O���?����ֆ�h!�Fc'n��.��L��e�/g(/�h ������|6/$O���O�K vn*�.��Q�� '�Mx6�w�c�o�F���sd�R�"3�[���͎�ԭyE�BR�i�6u�{�7"*����k�)�i�k~5j��BDj��U�Zp �
_h��`�f�ϛ?5a��UA�,-����f�����"ݠ%���Q��_�k]�]����X��o]>���mŨ��)���gz㰬bAX��4m8�����׏+<N�������ZQ�>����2�g��[݂'�y���:���?O%q��Kv��K���6)����}���ꬹ�&��L���_x얫�ڻ�?su�ɂ�����
!�KJ8!*&y���.�t���9����ƺV=��'�r">q��kiu��[V4e����3������8y|g(��ej,�F,��(.��1��u��y�����Q�H�r��X͊�u�CM�Aяѧ++8��+x��B�$V+J6���/.;�?+��&y�ꕸ��h& �6qX\�����d�S0�(���K��V��p�j�5�e+y^��f/ԡ������R%N�7$s�߈.輪�P��n���ه������G;����i�*XRjI�H��"���;wa�?=̹P��i�kI.p�B|뵗�oE�Uetf{���G��{��͊~!���.�k��O9\k�%�g�k"��}sV�ש��(����b� ��؈z�����K���'�:�;�,�U�\OC�P�̈́�a	�%�Y�i��V��O�e�;���^��_{�p�qJ�b�&+�o$�wȓ����pPQ2�e�����п�jS�FZ����F��ş @|r,���ֻ;et����/7UP��/� Λ��y>��0�@5M�#,�ϳϝ����o�%�ԭ�=����^�ál�Ȉ�q��2�:zXJ�����{ǻ������e�/��@��)
W
�M ��lWD�<��b��L�6��Z����]�b�m��w(�g^fՖ�g���oqׯ�8���`���>�Q%cZD.����<���8˦Y���z�	���'�Zo���7hI�<9O� ?�ƴgH���uy]��d7�S?`�������n�Zb�C�9��v������d��I�6a�V̋vK�=B�-����컞��4����;�&�	�����
&�z>��v_w��Vl5i+w�!+h5f�]���n��~�3P�q���-tm3�Hu/F����
o�i�je�{ �0���K�n>%i���U�!m�+/��9H�t����y=_j���������#�z� Z{�+2�O�=�f}[U�}�b�y�	�S�S����˧e��.'��!+*e�5��MK��� ǒ�n�e9Y��e��	KX8��;]�̫�|��&Q;J�2�����(Jp�.Ο�*�i��h��G�x��O�V�^Lr���z���RU�ǘʝe%?�8��e=dR��Ŋul"LIL:�3+H���G���Y� ���PX/�$bOͷ�l���Jq-(3Dr6�S�2���)'ѵ�-7.[�5�-S#U[�"�[�`_��7�WgdQ�Ib6n�TtD�#�'G(��