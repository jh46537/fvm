��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&}�d>l�ImV��*�"��C��@�Π<��Q&���4ZP����[����F�Hr�#�f�v��ݠ%6=s�`�{`ȹFCe;C��jЄ�1�'>:&WZo�E���W�0�_{�����+%��KgOhG���x�j�$�rր��<�P~�eg3�':xZF���D���̔"&�U�m�:���]������B�'q����Q�����D!<��FN��t�MZُ�
����4cQ@�#ؽDT�i�7LZ����3
�:�/.-Ð� ����<bԱ�͜���%7}ssV�?t��G$fC�$���LZw[q%���~Qm�h"�A�g��*	��6a�'�	ӶiN����2H#���f����6��<�"U9�i_emn$��/~�$�2KK [���pzk
�r&d�!�+��d�K�q+��U1�u���8+Wqp�)����Y�~,�rH��D��]�ql&EV+���1�y����g�%�Ǆ�D%Ά�B�d̲>os���$����}��އ���ME ��L