// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:35 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rL3f848zXoYdLAQUh8hg2PdqQrLmT3zrGni0zAoreAI2SvPkm4yZ6S1bqJvB2JxT
sgMc/Q1x1oQr5+6dZRxFdMvf2a/omf6BfRkb500rUptLBwtlDa625i07oMu3ayQG
OceGOL/BlNRmwEdkIi9gbgQRE2g2j8OJwSZLq/53W8U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30336)
/WSaaNJerViZNAtxy2AHGXDNpClnNba5UpvXGcj3Hstd3DtpQvS/6vDhfcnOdHls
CCclG/NqGK6hVWgGDCgodT4YtQSfP3BGjGvMFzSxA1VeQoeQIagfBHA9Z1xBLfAV
34mt1ffiqcPKQwOWAi1v9kyg3mQTbv2y3AFvmmQ91dTAbEA5t0r1dgZxYy+oum5z
csNFUUI1mVblbAcr08oK/mluS+EMwDbcW7dCy2WG7TcNGTrUpYDPg08/VwtybuLJ
eRvYndgZsSIwZRCgpXl3zxOcDR+84nSe1P4DjrB0AoN2QRosFu3Mw3+nfoCOhnQ2
ra/7F8Wc8C4ZOCsFVuh63IrSN+Nxt3IMPZhHXcUYs4ewsQX/c2Vpso2W6jvuwL31
Btym0YIik6ysemz2rzORRik9ZH8nQGzjMxFg5jNco0RPlDdPccqzNHLsn5Lhxa1X
OqJ6DJrNWz8UXMe4T9rMCi7t2Fh2iQE2iq6guzZ48rPJfso3MDctZZLocOqiYWOp
JJoC0YYSJqvY4afI80P8LXi47PuOAxk7+CR/nWXtaIBhsrKcJYG/tvTR30pqTXas
ZH5FOQZ+7Rz3Lzc8I9RLI7xDtFHPi3/c2KEDh4S/B1m+YywdpI5pPoB05BGSY4QZ
FdxfB9sjahff2gKr4F2EmwAUPPEN5iVKsp3t4bq3eQWvDRZFZJFwVyb/57Sg1LZC
q3OMHHndrn+ACad5kvxX9w/1XGe+Pasm7kmBZSxT6UJ8A14Ws4Xbt91srvqcpgu+
Kr6vnA5Mp74QQzCaUpMyMY9gXwPlfoaU+jYClPjZIAlX3jiIoS9qQxXyJ1zFBBQM
xc7ABD0ULhsVyeTsIGemPAjzJTWpMuRSeOtmKwCrd37N02am4AIzksz+XAfKp1Cs
YIq59857S/4wNIOpuPMstvVxM46u32s/vL2m6o2JFcSRkQcmzDgL9nQ2BbL563jn
kn0sQfHnraeVGcgk8kLMyMsuiWxaoBJnQ+vlfm0InFOpjrHW67PM5tC4BJDdF3zl
kP5Cc6nj+6kMqJPZwya6/wzcvUnWeZ1czDk8g9bmHZK1Btpce7UM6t9473qkTFo+
czkU4xHCVALfBuBN/7OPpAm62GdChGQO6ZMO+7hdJEmR7AmzxFe0gIOt0LnN+Fo5
H7YHyhCkUqAHBVIveMxdKh5p2zSeLbNPAIBgrD7R0ww4RSpfBRVa6F94wN1l/zSE
OQnnL4FQCgjbPmPuUQ1zK17dQhL5CNd+bhDNGJnsWKBAXWojGwTSn8U+iQxZ30sQ
HdftC0N1R4J4dzJhElTK0rfNhGXTqGJg4IlEgs9HiqxjzZFvV4oJDXQp+SfSFo3D
Dv1D2VB7I/tVpeMhIO7iCvYuFbmKeQ1iObQT5+x8U0FO0pO6G1jy4gS0Bfd8C5Ms
qlbtXKEpuTQPbochCTBqCuOEHTKXhrCnmX9ROK5CNrogyHW/1AyBAjUh6eSBaYOB
WeQCHP0DdS4kJ/vWVcXW3aPdunMcfXUAgjn1Ff8svE5PYVNkGntpvmi8mP1OKno2
15P5Qza38GXpcRF/e0wXC+p314N9+il/stdn0x5EcABCRMC25Dn/69QddiKyspFc
zaP+a3HIOoU+8DrQam9u2V8pXGuaXVNp/AbfcX2Golcn7mJndXT1Zjle98MmOHY9
qVDWH+unMyTwBOnu1f3pAJ+iOmmLUJ8DLLraQbcXzyLMlACHrbtSX4GdnxDdohfC
oUWX9NVHpF9LhGs4MsQDIYAyiw9vSgtfWoCLJfKV0xTbGLKJrCZtbA1LUiuJ15Cm
kMN+DAKZ4n4eN5gasI3zAJlYoYfkSGGgNh3raWCA032AfrInlIvp6xZImTEqqwsS
VpSRnSZ0RbDrSrCGMr4Uyl5+Q1SYYE3A/KCdcNSuvh6depdAvHwKPZCS9YM999Aa
dp46BYw5WsTWkEfCUVHSAdCmnAvdWLJukPUu6Adm9QkIMsZGgwp/5C47zktPVoyK
AZyIRxkE9IqBNZrOtZnE8tARsro98tKBthGQGN3LsB6sCm/m80xlq2FTk2gT/MH7
G44fIC/cYCSQmUWfU7FtyrsYdT3Ig9U8IrGxU1CTg/dv7PIIQeSum8qVJZ2gNC4S
QfZdbLtpeBc1NRdsLs5eSHvLSzrx4QJS2fV4UINKAKoRgH+RfBLpxi0jpRlngYPN
RQLEcyuenfTDi7zIL51luS8vGKuq/eQz2VRIonMBFFVJYEMSgRmWSAmSkXulfKw3
wZ03N7Z47SzL3rlF6nFRYLGERyed55D3ZnpUmblCUmCft7Oedua+LtJjlnFYLNut
BR1GfcihH/A7g9jsoop/mFT7Tm3ZZuAmAzYkAJ56YIHegDXGwvA+XJRogCRrVSXQ
UgQTfxI4knK6hOvJEASfMxm5FHLbaiQGpzKsWMONxUbrrVlG8m904zVfn+nnmQAT
RGhugEg8Oym+Zio1OWVzvoEEidC3wG3AXnM84DVMTHU6oGawnCpuI1aV/V1XN2Nw
Jc1pFxLntNOqnwK9R2uxepyulTONadJ1HfFBGoJEDjQYVEN08MzAX8PdNxuw5x00
TJIx+oK5fLODha+dp1rWnhcEI0UEsezrS+3k1vQ9G8qBeqIo3GEtFBx7Mcxy0Fho
t5ypqbqA8uVAjt3Sbl/Eei2fA4GMeUQ9rkLTpIQt17+oQf7qjXtUJ9PwARTqVV3X
Qa5rezn28QhW3k/8cKNWzWX84oJ9qM0eS2r+yKaRZAgTQ8XzX3PMT/LhVOdHJWx3
pui6Z4fdqCsJDqyF0dkEomTyfAk1mUwiUuEG0xfYtajF7HO5ngrvAzr5r38dGn/i
nmYFeDoCtzrJltWk1QMZTuVwW0+lNaPdh5ET+lmZKv2fwED8z0pzt235KTUuMBSl
gWsM5b03q2tJoPI2Vva69/ZqaVI5uO7O8Y0puBkAHmnJbwkyb/yACyFgRNfMCHxu
h3esdGqeamqVKlwBRQQVJTj7ubyQ5USzcmObRWoDOF+R/rPBEwEY6NYUg5gFcOKP
mJSeOJd5dlJCJbvEPRb9iVRrKUHnnk8Eyx9sLlZ/kplvJo2Sf/D1ijF59UcN6Y9d
ALjAz8EQvTu9uxNYsKJEpcb+sTSZnx7eXCdZvg+GVCnViFBmjXeSpqA9QVgumuwD
snW1S4HsktkLD5wuVwhwQ4Jan884QHIPH/aK72G7022NO12jAuMOPYKrofQgMA/U
EY/JCDdSSpc9tWZ06coB5Zy96TzFV00qfFFTugrv7A0A9jwKAG1hZMv5IjdnjFmP
NiMIk3NG5f1H95ixt/flCg3qOX3xfVFtpbuzRDG2cVLSwIgex9j/raSIvKwDoANd
Nmy87HhpdoxAkXm3FsC4LNvdyZuXE/2vV0hKeE21s28MFIu+p/6HICQVejelJMd5
D5vL4uBxUVEF51qY+XFqQTiMUBow5fH86GFeMLS+3enMcu5fnlQa0F0jGbNR3/AW
YhShrANb+j6pZW6zDJ1nyekYNVtBmqE2Yh9v2HXSDQEak9sWJSGmYQwiWBD/DWox
hKwchKWCnZgpptTT0Bn5kOhPK1z5wQvsZNRvGgHx17wuKg3CCJrJQ55ZBaPxiXTB
IzOuFwO/ojqQXskRRNfIW8X25+jC0QSEmJ67/KluR3AVf9zqYlVZmF+ybqU6DfBs
42KFopICKK0JEaBt0X2PgZrz6adqhp/FUKHowQDJJ8yotbFS2tmBgx4mMq4A9D+R
dR5y1SAKp1zjrBFGY9yuDPNufYHaOv4m5juz+QtL7zK/HFEN7Hih+v588zr6aQDn
ItfOtn80ZyNt0jp6MaZyHmEm+wE+lFFNo2FjPXJ7iTVVvY2aHz3YOG2+xheRIY+6
9jNv/s8sRMbwO7YnAJeTUjwZk/3NQgomWTb4UAqcoIBMJnKyvnGpjB+lYXZTVFVE
gNA+Og9Rzov173qY/d9kKEpMOB2KPvbv+m9JkWAvwM4cm//lTXf4I1jbCUASAqwT
ewuGClgHbB/p5fztOxyMljt9bHF52yLDE3N9Vs/jHvO5WpjkQxwMdK1cNhak5Drz
HMs8zgSFQAhaxZMLXDdOI+hGAESJbtDPXwab+AYHCy2VSl0aqEIDsYq462xtrwR5
ghXz0tcurCs5ewm6raHUUVbCU7JSQ5ipElwcs8+AZmRFIT64UUdijF5kedIkbfib
qjZDe7scV3MPxuL/8hqz35RdotR7PcfF5ao92oLf97oW/APmLKg1Sxy0yE8dBMxA
GedEyAqmL0Nw/G6MjcuzWdoEqLXTeJ8bNWtcL26rtIRYhaNuqmKhou8yjbIN+bqw
zXUPynKFwW1tczyLViYU7YHAbr3YA5mJChvN+BVh3wQdUetvyU2g8BrqPR68Jdcj
xPucliHbL3P7mpx4jK+46+04QdUOHZ7TNuRvsQ5n27xJDe3RspdvXTJ+kOAEzkhE
FwRKfn/sdiFewEp9NGcco1W+oiaTcYGbZFF66iwxlDjsPy+qgtOXM6YeayUA+cTJ
M8Kzra3SdGqFAFOaUnnqwhKqxXLYJdFQR9D5pF5cS7NPfUbAHgbPjf27RS56THmK
zJ//qYyhpKmexMITTZ7m/rhZqC9OmiVXPFSl3gmatT3lO6ehKj66E8vVL1zMYPRe
ngtVLeESc0b57n4VrzOdNSOJQSC+3Kgj3pRJ9EQxUNL3pHZtZl+i86gjf2tY2AiJ
usNcBk748pRHa+pSlhBUw58Sc83AXWdC2Dxx4XZCO7CZras5XiBV6ejUe15qseho
jPpRSlDCl9Gc+YdNnTpVPH0PzNFwIS0q3MlYoftZrNOY3UWGJnnk3ZgBppdbJ072
0vq4B0bJG+tKau2EvLwj5dpxCP1QW39IN6qIaLm9fp3TZ4CotWOlmfmu3Qrv7qsM
gNgHRHjTUFD/ncpCd4VXEcf+1vzxyll+Xdqo21Eby0XbuQWXMrhRkQF+FO9LETJO
WriFYHcfxxoDFefYMtjlwLihIiNEOqr9hJYOEWJKqjg9GDS+VqltEE4q7K/1+SKb
1ZYLvYVrUAIOzRoSd64qtfXJeeFB1uJl61+2k5WJfxHJd5EWhRrgKj9fqNdYUBy0
nGaPHRDut7BeDzsyP7BNsJzyibFptaRQa2IfNjzdyENFFna+GTxy7D9FgReqK/j1
VfgET/EUCjaLWtgZW7s/5LLOkN3WH8wNQkySatopU02hq333DRTOYyzuhU0wVNUB
UW65BZSDNt3nKhsxTuHPBHnl96lC8Kd7a9qF2yJIkz1uOkydEuvPlN3uipUwMaCp
rmeavpmBs530bgCBl5GjnvbVqazMz2wA3ymJTKBXi05Mi/Sfj071AiGxD0vdubTv
okNJG7UKWD9jcuqDKi6XlbvI8JsUzZEqZ4fKtqutgs10ywPMFgUL8ZsdwYuwhEqN
xyjmb07TFeK3pVBnozP0YCO3VzxO+mh3pV2P7nsf+IRmCPJCkCUmUuIthPJnk+wl
E7hqFbXZjyQFasWfImlLULu2pO898s66JysFYQQ18VuVB+0I7EoZXMizMZAD6Hc0
ux7ixtmTgP1dWueZOD42lkd/txPLSkxm5GHVTA9riqfjHnmwnD1RTISlcOie/UKC
UBrsvYYznYlEaLQFZ53YoUpX6V7i7ysxNRT4vdYdTdEPjMhPPkmLOlhsC9z35LJl
p/EIp0nad7K6Ezlny8TFiEZp4qWZIeJQp8Ia1oaMQ2qL1T1MUlZ8JHCBfELbcrg9
kpauCiW6UwompZlIQUH9Zj1pE5oZwxD96Nc+3U8ClqIB9TJWMOQiMtVrxxt6KDyj
g4WP/35teG3H1fPfjDsxdkZtBWPYPP7ZOxSGzGNt5qJJStJ98QN5TTzEZy1SIiGP
HUhYeBmNupgWONZt4+jzETHQtAyVdzeOhzNqtYopnKy09iapuqNv7dMGZ0QR/OlZ
MYhFsJ0kWI18A1RZbMeNRd7Og9XtT43fX9xuVrw47nleNPq/XlIotYRYvp4Xz4Gr
wxmaEg60m+PvRPlxE16LAIJDZOshHcS8LJfqUmhXfhotfR9WFuE9dBlylnnY9d+w
pR571ah9BZQx0ZE+lhVl5ci2twGeLSN0tMHfc8/hhf6WlYeXUmOEs/lDo1TMJeoL
8XYAtftxq4s9DTexn1VR+WqDDtG2pds2/Y68fMwQS6qrzQxCmx9Qwf6DpCV0r0Cv
UEmW22BYPgKiD0QyM/4DIYTvrZi8uggSmnzMe3gTbenzfwJiLFyWnG52rq4e7au4
CGPNkICBb0vrPaqk/54qUXKz1djKMGAYjZ+drK2hncKXSAD0rGtDqWkKPGSjBVo7
WwEeEB0oSBy262V4zkDuuExvQbWVdFamqKoJeeFmn/Ri45exFCoxyFMF5MDEwy9i
fnoqqzNna9cufI3S0MjBjtOJwOQpfdHHGkC5oMzDpLGDt0bAwz4dzW87wn7oaitU
C3LqMnj4MKEQBLiLZbERENMo7UJ8Y6OZVs2WbHIKUsnTg/bYvaqG82sGU5oHAlcF
vS9kbBVX96g24oFBRmIuw0PYSYyMi7HpNsEaPjz2loemOI7iWRfrh3ROJsIHMrvm
e4q9YuNc11tbjRhgUNggjP1GJjW/KwQk5ywJ0J1kIZuS1i7CrfFTdWcTc5pXw5P5
ViW+JSKopbuBP3943q7KxmwrIyri/DPeioiVcYgg16yJ3cMrubXqSEOygVdLKaZO
0CDA+GrLA5FCq3cxV2p4pmSYwEpbVgdnbHpKlcN3TcDH8Tj9vk3QSY1HIG9rQDLZ
vak5FJjj37diekVXQ2MdkgtfBYoECKaA7a3PsE34Ysic70uJARoVCo8zmbcKJ29y
Wk5HIeEGrupJhtznpC8fECv4q3OfW+dXVqFNT6hr6Yft077jwTd/hCfGNTrANBD9
Vtx1DyauiVB5z+hNSvPw78TimFt2KX1jWO61jfV5GEQ/CZzRp0Fwd/Z0Q5Eub5tJ
l35TIdGJQuim8iiqvQJY+WJSqmyl+EeXMrgnPT24Q0U6Ro+phjGMULwkYAgqY6/Q
x1l5ydrVYpn0SOp1c5aSYDk0znWr1VV1lLzdennAlvGkW4pHSpTMvgColNcV9Mys
27u9QpTByQR2agiUpd8q05TjqcbkEvHTLSe1oqGrHt1Mrzp9ujoTUrrq76gNVvpQ
+bC/Ebz0w2Md4T3DNHnVbKD66D4rnr+ko60XekIDvpVrHok1Ho7Efpq7ftEaQe1N
K3eFvH9v+vYpPp9SJVkLCITdHiX0xTO8+aj80T9JWwNXV6DcknkrmyXyROs6suSn
CN9Ws1nksjuM+fiQQhHQ5SCjkH+VZmPQ8p+gqpkCoGWc38MphqVJkYbQIXps0994
K+5xiO2Pe4dx4i+HgImRkMsrSCap9S/Dy/9DuSsSYx9RuQEJoXfPnKxIAkoIEKf/
0278SaH98kd4We54QoqAj1cXt5kEMkJOWdBvU1geGKTBGI2Op/f+FBDfXmUPS9Qt
mQQ4+5vkWYw3RsDK169KRUJ+MOPT9kwv1vxEJimPMrIoju1nwgK/YZvezUstI+3l
39V8sd3TP8G5z+qrm9kx6QmIl3WVNPLTDzPb5GUGBzRIuOjg5ceMUBiuz4zF6wL9
ZGTVnqiLivNOHEwicHQ0tbHvIye5zoZcItpGkhX897CKniqC3RYuGyIup42lOO43
7kh6lhouMz1vU+9BfEs7kYXGY2uL3V6HHWnIjN9suvtG3rut82eBE+QfAycJrPgN
lmPq608C+EJb7anI+TTJqy+2bWyoL/SsXnHZCiS4lbvp+YfRCMNRYNM/+1GAUBbm
SHjhcY5YydCuan5mzJdXjTI1k9x9Sx94viE625Tam5NRHBe5U17ng85Nh5cNxcaE
Wr6TE75QPH4B/+0iPdYueTySSN8r8RXNA4gnZdEJf3kdSzVmYwdycsQKrVl/jpqu
Xc5t4INvBG/ex2jjaSYvaASu1bXMOGb5Ah9KOznK4iWhUcam0GPbsyP8oGlJy7CW
Lmy+gDk7SG7FMN88Vx/cuzi7JRoijU1VkJeu55oOhLu3gxwXKhdRanvt8wSvchr5
ki2jdGqCeB2OACCyM/v3dWPj4U3sDA9dn5LGpfIbtfURuBWjhPYVTFMbvxp80h9Z
NHp1Y9r1BPFiV+o+hExO3hfwowcw5uxjqCjgVB78dx5GUFSFa/39qODH9HEKQHEc
M45wEfg/B7t3Ag5F9eAuPHKiEWrTpVi9lzTGTLmARXYRhCpwTw6nkTl/hB8lg+7x
FJa+UE+GGWRTkE+KukdtvhoQtb1njeaY0Rg7ziEaFdrqFYM5Ac3hCfJP/SNTr0KG
jr7Putz/YFx+X1LK2CUIUGxIdXHbTPRTCp47SACpmw44EzCIaWsp/ZHOZIgyVKP/
kvjytFI2bBxJ8t846rHYGwWAkFDdQ6vrUHJbx5glICOb3LVa02KA/tWTXQazGjyD
BG6xmcxz+hdu0tyY30NXmb5/8WAy3T0iOu7J2q98r9P1+7S+JhePkDv2KW+R1tmI
Tarppbgjy55Z75g5jwiuSdb3x5b6Bmm/6oSCmKP/6tUDv/yYdLdDV6GVY2oI8Upt
SplGDhUCx+XMN4oF5e/8X+hRJ3nLiBXu0e3TIWcLgKSVHchM/LROqRsoTu0ihZLA
Y559/SpYoNorNc5ERkxlxk4H8WLBX15XdzRyFWip+/mSY0DRS3VeSYAJrGdiWsmE
jofc6PQ8+4N7FpLJe7lqRdWU94euF4QSdA0ubPA34uz0Vk3YrqaTMXKavhd1uyOq
ORIUL48Rp89rlSr9j+gmaWXrxFy10/osztcKUxPu4e8fukgPKbKF3gANcuvhXt4L
lOA66DS8nvqMAeZ4+KhM06f9y5pwm/aPA9/sv+PErV6lJuHpay1d2I2KX0SgAynF
x4z22yRdAhIy2GfAc3sx+VNHaQBCDe7J6fPcRHgsfwy6TW1J+zKfyjVXOzEOsmFu
3Ob/X58YO3fp8P9TFzkJ9rg/rESQoVyfeMkgtlvLm6KBRKNeWvVyuNtto3wMiTiC
bbyjaYqR3BI9HNNeqcWqsnYc9bFbqI1Eh4HZJi7cj/JzJcOr1uqAuqQnCkgeBsQM
1VtGiT6Ywx8eECy61sZ5D2xcpkBuzQbbCdqktIGd8tNQgVkg4d71euIUVxg/2wq/
qjFmYBx3p/I+4HI4GEpuL+sgePyApTGp3X0a9fz34dbjOlus66x/ACZtfQji2RfF
JcD3sXQ9BMUiCZnWsZdgZzfsavVWyx11PVe1Cy4lF3tHN8UiDFsgNR8dXMZutMLe
xmdIgTESCmG3hGKtHMCDT9xp6uEIyIrBLZKSdoDVUa0XTWwoAy9L0iokxmzY1k4t
5t0Uxy2M7+uaJHvrYwKJcY/aFdM3xVQJjHAm00V6D75FLlhgKF6bMlgytXYQPQUe
/QDiiw2gO52uO05QkVNioXP67nTFETMZavT+s/oGzbhUNn/li5kKQ6JJqG9xD6/4
U8VgpfCaOCfMl8dOcuubeNIy5bp+0+WRl+9/hGbBtZMmxwL8Ilx9kneVo9tS5NxD
igZmvwQzqwjmlVUsmRRlir9B22nC355Xz4ovef1gGkWQAx/Ami23vQGF/b2VT55J
rwLm7b5hw6zMTiWi5C6r0hB1XqqqFj6ykFledHy+xbYPRWqqqX9XIonFsssW2mN3
5KnooEZK8jcRmbHQ7TP8RRShzddaLYabHtvWE/830TTHKbhaKBgcTo2EE24Dsmiv
MDZ1OviiS0U91cq7cFA4sxJyDP8a0vyADTS0kSomBdGJv1loQyDQDsIJlKsbpRFi
4Vcd7dvildFZbEp6785IVDyn4ijxAZE/F2/F7Tli1wWMA1/0pJ3wWfI7pbP2k8l7
oee+u4cx+sf7WMZGqeESMXX+ylqtXIbfgqJLV1VGThQpFvJH9gs+JSjei/Lz7sR9
O63x7sl1yoV27TUBkIrhQHZIFNg32OjpAuTbaBQbWRoXXOR9cvsGR+jZHhKpoN5A
18M+71oG0xqYNVacZ1QsO+FWzgGIgBao6UcmS3kb7faHCVhvLgOlv8e97CkKt9ZZ
nBnhySxLgQp318oOs8Kt41C5svZ5tsxo2MZqVSSTNWxqPLi1DfklFkdU3xPpWoWB
GIBvG07JxNOl+sTt23L4V6vujza0FS1UDVgAeRgnO0eR3woVbO2bvIZ4jpx3AQGA
YsaVYsbtc4SZvU3pATFk2oHe3C/xUYh0nm666Sh4FhkMUAt8Av3i0G0Q0R9zSzyU
pEHpIEbbddeesDFgWkn4Fyf//+sILMFSz1DbGvFyzcrlCd+uXWY6iuPmL8fwiBvb
B2wi4SS4HPzItPVlcwSLPrkD6FUkPywjH5L75RZjN5BqB6+VuiDWe9igRQtLpsOs
8gAE5IrYisYAkFkAcw8RdDH8IHQstMTvK6PFxgJ2YnIHAAO7GolnI2UfETTW8bsO
bNVT14DmbH2iecssTKRQbFc3LgCUC71E9Vc9tECShAnPkztZX/vgvdRWvR7j2J6m
NRdhGG8m9NX68VeEqOIpGSLFdPQ86Dnembno88Ot9N4SW1PDgmircazv8DxqE2zF
f+bWhQPlApIcn27maEdx4zfZ2arJNKByzBqRk5bm2nfyCqYBWq5su3tdZJ7Hug+A
XpKfZTlJ9p0wqzq+TfYm5wzD0x/5uOW5uyrLCwG/zzBNQwhtfhugBrFVQN5Fiip8
cVnIjpdqsh1Oo6+zCoTwX8QmrB/nuQIsRDuvmOdMVFji0Ow8xBt9RHKJJImueIoI
++vAw66fQaeSt3MJk4mSIqUCW1tX1VPgQl9tAaW5Zlm5rtDh5PB8hG/HCCzhas7A
niqESy20C+5A4b1/4Tjte3Expz18xVoDDud9VrkT5xrC6hoLfOuJr/bC0f8IvLkc
ZLlGX4TFfrQAjyHESTFCWtzz/2G3Z/qYt7SBis6HVIOI4gQdEqJEk27j2ItnkLTk
ic/EuOK1VmTj+KdLuyQg1bGpzHw73A4Arde9Plw3K5E3vs4qMf7lEh+a6HME3VWt
kEihO+la1xAW6Qvqs74Bv7W3nrMCLHuvVYMrplPPfZgnXUQzsL2cXsqrthheHR7P
0OTmgSUViC5nvU9fY+Dl1wmNc0PldHTnDbrbSEF9WaDJueDBi2niHChXYPphfUJz
OA+cUk+7Ds5tjnrmfwhlQ7vPDJFqV4e9LPNOeryjaLzTYmyTt8yK5uSGE627Te80
fkn6alyk8SD6KoDUI/Jg+x3EIp3LHA7rRiwMvWVijklS4i/IGThzAOHhR7tNpeK3
oZr2lW4BnQbuo0/D7s8W2zDbuivy0yUTLMb+BV6xH0dxQMRVTqDdQXSaJDnzxDSj
2XQQmU7uQ2LqAo9LDXdIgCEOIyShO7u1WzEec/njaysiwZnHKbzhyUwmCCZsb9IS
pZKhibY4Npo8CAHdL3P3gp/94DIei3+NxVDL5DUbWikaZ5vBqub1rhy1LeRBB0SO
tiyxh429JQnR4YMfsmtoTLpJ7jFmmdJadbKF0UHkplVT6YodSj4EjmoMT25mJHsT
3bEnUDN117TCDbjqWbDTBz2QffTVxO+y42KUacqw5WZYCXpwHczzC/8m+x/lMnzm
8Ipc1IN/CVW6AQf70QTwEn53B2CP29WDV/Zc6YCciHB7kKMLsQktbts7k5ahiYRF
2pQHDvFNhc+HUZeD/vP+V6AWip6rx2sh5afevpRTFcXaNXbZxfoGCBWrWhMtxft0
pMhQj22G5pLwH6nnJ6goVwBikj1gS5L+9BOj7OHkfQKhyHsUoXqwOaSxAXZtYc40
bsxuPJZYCwtYm6ni7Us4BefVCq0pnPGZYp9X+d3aw1of2FFw8FO1fy3B1qpHcLwH
3vaeQorqsznmjOlrprGklmUO+Ih79Azmei8S78hQIt37b9L/cdaYHfWO+stN37Uv
DS6fS69/2jfaIYElIcFcSeZh1wIV55K/zvwyUayJq15KelS6CajpwdobV7N75LU5
cwqs9KNJQkqkvsbcMhaBIkkVabnRdMZBMBHo8b3ebFps8nOHE9Nsx4N0TAD9ju/W
/2j63K9mnMyoB2Ix6F5yBUKZ6jbfuamfiLYxe3J5PAO8pAAR0lyrso/NVin1/mtc
vPt/Iq8DiD+BS3SnS59sYTYLYX1k+55s2TLzECuTl0bgBNLaFqMezG8z/mxsiYYh
stWOyeBdtULsOfeVQsJlMbQnIucQpeEGMeas5mTmDS1fMu0Z8v6j13uMZ+Ichoa4
0wNsR27yb53ZDmrxWisDxmu8nl9WOh5vLGXnnvm8pjfEMVCa2AMAzrVRRmg3nFNc
b2VtqeCN3VsbYYfHFfYf87UAVc/gFev9drxNbeXf+6Xz8+yqwdcrTocf2wuIjbQF
1RhOjMl108OTi+qGHX/l4ub6aJznJrbMDIf2wOcLlhCQFctdvvzS87RZ8+a0Sdsm
I8RJyHiv1RFwsUnIvneFQaj7jVnvuQrB+4Slnyjgu/w9h4VwpVIZ5HgwtsjRfghu
iGdeWbLAC85xW2vMSo9wo9xU+TZdOIqC9GNI1VkG3EXXtLFwQnovcXEw8vlQ/q5Y
AyLCobbzcmEsvJKTDvXAJTEwScNcMy4WESUP2TCM+CMmAwiu1Ox0uHcX1rdpMk2a
k5oN0dCQ1bPtUGdwqvHhzW+PhlLVC1gItNq2lEqbfxkdmP1C/3lotyow5r4Rtq/f
8qjTgm41JuT+2yNYuY/EiE44qmveVcNNXi9W6TbceGE1Qh9e5+y8wm9U5EGFhllN
XDoRaPVZwR/7ne3IYWvm8C4TeWDPReA8S7uQypguh6W3jGJvJCkmBG6dGUSqmZa9
CQDAptG/ocPdmQlKPuqwhxy+1abWJRh9NIIiG1/A+0H+pjCRnuFoz17VkfQRbOSX
lf4YkWcEXx12A1mcO5TYJ9EzO11HcwUoVqP5jyFwKqh0G6FdeNgXaKmoT5UPGaYx
Y3UygB055/MYJBWSIEiYiH4nY8Rqb3j+3TV0FttD7yaNP6CB0eCi7OsMp0prRzdP
VtiGDUPVxzGfEuHml0qPfBm5uZJ6c1iNX7bj2APPmRC/YwsF1ybBHoqRSR04Uk03
BcVkgSD2HmlOYNCUXYyZzdr5FB1l7PAwFunS6dY0XRFXItba+Xh9zmqgIy9Qh5KL
J4aNdc8zMjcc7/ly21blN2aPwJ3BSpXqzhlsLgTr3UJu/GU7bBiCl5Gx8HDki4gN
wsQGCFgp8osD7b0+MxnJPLCuIxdet5nlk0ubmw7Kh5I2QDQAYBa30J53KnfjpavJ
twaa0xhPT7kCdPrF1yL5fQAs/g09r3MOyood0FpTZmQmS/Od6XoVlVE4vLoXx3t/
AIVnTJ08gj+FcZn54if7iuIPutx/yZlZP0xPZeevdxhtMQOAVshObPv4XLl8NR1K
uCkgBn5bkvu/BrXF5wUsWN5bi8nthbQ4YFy/zgKRW+tkCzZmVnU6HClBnhGwoV8I
/tijAB0AaD/V7mJZlh3Ep992PciVExTqtYZgmINCw5Hsw1b77dn7b/ESOdj1BIMQ
hQjatQJbzWjZMh3/1d4fqLMUA2qb38GBM+V9kmOM08h8l6ZmSDNRurOzMTv+Pg1/
N+/bJTYZthE3h3pR8q9xoz/GanPlrYSKac8Ac7Kry1aZlOUZDrPykuL2EnI7pb/M
MEIB2NV+39fBY9LTz1x2EAuOLK9jyCrSQZowhO1X7hmHQFgpvTGkz8GMLJQlEmfj
IPXI+UeNBLqLNbkZNtjxGWXcD1s+hnDp7BUM9gmyYYNtA+CHu4OTONRMxwVOzQ1x
ntTZfVnfzciaoioyXy6fwU/Z1qHoF+eDxacjphQJdLrSDxW5Mv+QGMGIc4bsaS3R
s8XeRLvWvRen7A1mkoyaHtL+qB+zSbIMUUVHFPNQp/wnja6aKSGxtcM/1jFG9yhK
ghprX/emFy0Q6/s9xpaCbka7XTKB7kKWn8htr1pGzVBhV93zz6BBpqYGps1DKqne
3X4pwlhlmGp5gI7jdN53+kL45y6CWWEk+308Ibm59zys4/nbbviGVjq+otach++G
PAKOsl08wJwU2mbXs/qLmfezx5195ls34bmz4cQniRyi3Z4c1oc1V9nZcaTP6jGy
gWS5gzfWnjvjMRcdapHykD+57dsBZf/4dbAHQNm2GA4/o6U/L9K8jBu3wU15cRGL
wvdxEfV9nSYlN+gLgHyIqh2GjAExMi5y5CEXCczXfqyoJiwd7AQGrcZwAMiM9Owo
H3xKHhnuKbrc80NdXbZg+8dWKpJdKTpYDUuIi/VO2pB9rPQRWmV/FbRZI5MSSjLG
5L1lRqyXWPQAeaNsciuqa9WknQyHu/s+uXMHn7RFf83vBxBgl+qSn+TNBmMWhb1D
ynYMZVLs0c+AFNk9S8A20i+gwNF1trud0Ktc0P1How/ZILqXjlGA3w4XD7slZNR8
9tNH8Z9LKQ1hEgrbAd4hB573t+YHyUchwSfoR7r5yShHO2/piCUtnqlYgtm8Hcsq
bMN5NavyJq6CxaPMFLu+yV50BoX9bojjeABW3HsZ3IIrsHLIrjLEaz1K4+y0HzKe
kygjuGD1aSQDbZu5toxRNsGdbTh+Lo1SD2HippB5Ch85piqbNFIIdl6Q6bO11/H6
6NAjSJE5NhZSyR2hImaH6K8aHrN56NzQq/FRv/ZM3AcbYiZP8BvIp7+tVJjvkPIc
T/rKCR/LQECr6WB7UDIgvN7MFVeAifRgSqG5f17J4jUNyVR7dXix8rpb/symXpIS
BZcn0I9DQlirG6jqwfYXvYmy4oKpH+07uc6ClRRANStcSxlwzsqKGMs3nGY1XNNV
BQHm1qsCz6jd77TzR3V4oTNt/vJ9Z6whvVbk3670RoYN/kHbV/KoLQMrq/IdVt41
bmzhZ2chcr79D0jmpewhNbNF3/Cquf5ZAwjHwtqCUrzMoO963ClhyK7mkE1lXp3S
f4L8KKvebb02XfXawfW5Tqcb8LQL1jpZeyVw2bGun8/zdZE/CZmjjo4KDLVM4N+I
msEmJMALukPPcP38cBT/pcxqTrW9jyo4630Lh2GH1dzuZIc9m6n9u2rlAJX4Ye6c
Yo7fT7D2WRuCeyIUf8L7f0R5kpw9DAjDPgjDhmkEWEVFdI6K98BpfdBe9EM6TGyN
J32S6Vs9N+r5Qi/kgkI3RLc55LXcyDXgAfzB1orwZxveOW4lqpFV4evVwmBpVR4H
ZQFzGhSHZxXBRwMtjYo4h27tpdZv0vKSUCc83xynkFL6rUh0dyHTJNtn7oYuY5vO
bsdaT72iSUiYjkJC3D6GxiLGolDNpUZUaH3qZ5UZbrgpgxPV9XZNl5Zs3oFL7y2M
Sz4prLaEZtJv6tXyiCrXUN6cgGTglXS3zTUvs6v4S2cYsG++xQwn45dAGLzVhwQ/
O88DDqmJxOzHe0XKSl/DSNFC8WYesEv3+rO167Kjg7Em/I46KHDCXycEN2ce5Tuy
0Z6w8LTF7lnKEbgajy7DNr2QcpUXn5A6LO+cL5l/crOvpOdRbh8Zc4AGXeIKSsgh
EDhyEmfFlRkLomABAqud0AKd133lggU44D8/22uVyFwj3gs0JrLTBtxB3TNxL1R6
NHzhPU5GVVL07ElFPB5Ge0N/H3IVMYbc0XS/J1qCtRIHtVrrLYqSyV1SwqK7vdmI
E7B8FGpkGna84godr3AOzdvrYchJeZq8c1juu4t1z12n/WTWXQzq7n0hBGq0ckf4
xP1qH03I93vAJ7YEyFA+I5DmplMxIa3HRS9qKFqrgyxAJV+DR8jiNlXCAELnxxdU
+q3C+w/iYq38Q6UwrOic7O3dteb2T5Db1oftzi/YRAOh3F4NNRjGiJMkb9q9aw6V
058B7ecA8aRbx/4dCuuoqf4K2DSdE7GPXyKwG+PxLO41SBe47zURfdAjKkuTAK6U
y0+PpIPP1u529sM3uqxznOsC0AHMybYKgpsfTk0CvJ1xfz1GspN1mMfzfdqIMF5A
+9/LlSG2DQCutCmjq2fUlyKcnr/xTTJBXZ1LiFsffuDdYG0AOtloeAFDmC/RfdN3
wRwoWn9vhMItPZQRJg9Lxo20Xtf+bus5NoZQapUIsYQhIIsEsmLIqsqWqmIzf6AD
i/LnHEO9ylHLNHxNVPe4npfAVCEZkMtNL5pIxnkVByunm5kUhTdPwFCkegVLU5xT
xtuILII67vlxHd4GeglvBCAZD68VYN3JfU+HUOJApT5xjwXbcMDN6rCimcb2LGtW
bogyPfbvR8phKkdrAmEcOgCxxE2q1Kp1kGeZvdRQj6U/styQPOUN6w+yFB6dEpRA
HIMaLm8g+u2tZuIYL/KhEwu7lnXN64NDCeOObBNwkoadkOjeXuBlQrBHQwlqdqLt
nznFnJnaGs3pmJZBMHh6V2jhljbQ/RItZlbAv/4yvG98QYwcsrKF/EikgEeLbuan
NHkERR+hwqHV9vj7iOhXDrDoaUxA7o2UWpMzxR2r5qCKPlbXrTdkshEniNxJBm0R
kkJi4sHnMm30t3TKl00E2jTxF9OVSGAeB0iq2NS8Z0wpWpTuaNrNXR2C8fwG/J4Z
YRlBZeQFVOIxBHeDZ4yOY56SmiwEjU+nTyle+Z4qjwmUuOX3Vp0v2UWSVa87/Hwo
JLdII1mnI9iKNZY9W3wuh7NPQODRA3nFyMvFpYq2jz0Md6MyF1F8OCxl418pqvwP
ifHMLGuM6pxgtZVHwpmJe+g/FJzCe3jZEHIq/eyvXgSlygU6GKA09t9ixwYw2DGw
JNeoqFP8+ZWbi8Ijtqe+vMe2uImriSP4ic0ycE5/W+6eWZOyQh/qnRS6fk++rvZ7
KkjQYtJ3w69jsa7OuX94Ep0WVUG+N3eZIaIYwmp1Uq+jzjoxIyCiMiyMIM/1BFGe
fGmf1XXJWRki7xDGiCINThTgS1Fzg9A9waU1nqaEbSGaoUzrvQ86Jx1N1/yVAQJO
mCIpuJEUyTmpYyRhwfDL2WjqnAv6c7zVgh+e8d95X0x8Zs5T7aPE/TxECd+J/xLK
Zwf2DHY+Auym9m10R4//ZPxqHMbudwDW0QLSZam8FwF/jdv53ZPnHT7nMgFOxuV1
0/o5Jybn15ReegMaEGIG/UCA8WLkNMzgWmvDkU8RosMtymwFodhm50uy9GeIlBPW
MzYnU2cHcvRScfqr/x4fTzSM6LkOFChptYkncT3Mgnj9kIi+q19LP6ikmAgyKep4
iV0dYLMrO20/2wSHHrppHoqGqAGfUnTHFOaNnLqyCObpHKc8KgsT6mGFWsAic9Ip
6gVXbtu3LE7OC9fJ1WHfJV+yEy0k8NgZ6CgUbwmGpqtSedIB0nMIYUKJ7EfhVj1+
dltlwn4FkIq687uOhSxY+PQR9Nt9bzN4cnKiYpjTBoLHO+JSmSpbROuZ0r17qg7P
zoGKRTbCVTJyxTJTCmrHfywxqS36eoEk6Ia+SmwnmzeILQoMER8d/0b9xoq+d/3g
ssnBF/BQbZwijrHwFWni4m4KJ4lUkr75FMT8DIFD9MszlznOUJ4IRboS4z01seHC
3KyUPEt+3F8gZeAMv6zPdFxoq2J6/hvdw6mOXn2Vd3BIwqV1DmmCXHPXJsTov/Bb
CAdX30EyWm70LROOCluo/ozNjLICj4fnto77ffRaYEUE3L/tFmM6S9HBCQ01ZDvi
HzcrPGnQA38rDWHWRDCaz5u3dGVt5oX0bQVf05N+m0XvPmohvNUTJMqfXEvEOlW9
bV7X3iQINwdAnkK6oD7ZmGKh7i/iEiJLio/Y3n1Tr6c4k4GPXIQNWAjuqaOBk1Z4
NyrKtYmworoybMHB5ywoII2aJMxr2P2hGjZA/DadfUeGeQVlT7gOh0essJvGCJfa
rn/vXNE2Xf+w8+wL3BzbZtBjVDnj9gLcLg7uiKUf6PUHFAfmpDwRvMKMJyB3tfdj
Vh2oQ/zqo/zdv2gkTO+DomS99q7Zvdc7fTP5Laaqyx/FFNEKoQNV0PnPX7AwFEnF
uxteJ+wFIZ5LGYPrQCNMTG0NTyZ2VJ6n+hXMNqqsYEAmXsszbvKyIwc/QBHRch1J
2EOgcH4d5ePVjG+DUVMZIZlC1EQhS6ba4VirNVbh6+JTkwmmOwFbomkIctV7yvxc
ACDoAASA2lMzaEAVr6E2VvSCbSIwrzSuy2AVTSj6m7AtmIxnryL4wGnXry3h+1Qv
FQ+Yx9O/XVzQcey50uSz33/DNMKRwD05CCwDcZHJ4LkteXgHaS8GnWkYYUKWFdGp
vMw+Y2mZLD+hvUlFoWMpzXcimjML/xMraUO+SalOL0YVtwYPdBeiIQRYwiaClwoq
GCrHhvKoPcuDPjTVBNTIZJ1m9Ae6qIH9VudE00vF4qGMRWEhW1UxDn1bDnRomtZn
1RtFzGLeNuYnTxa8lH2V9f0qEmf7zq1LbwDVwu8whuvTSsqCp61+Zzm6WfhMJvoP
kVYkP5gLGIsvCxTxJVTzB9LAG5Wnh1WVq7EsVmVlm+Iz8ZvHJFLoZOdQhJAp68SC
IriWF4CIT8osx1G7fv+yGvGtduFYNcm7cAqshw3FMQvmDSz7CqmY76c4O9fBum0C
2jquDWs6yooWFMHYJIhriO5C4hfZS234N9sypvrnqTqnwfGk46mOVBmF7UhasWjg
2ci61xdRaMCK3+iyBqQs3d3aNZOIcBXObvgF1eLfohGTzb8LUVBZE46IZ3Ba9UnJ
Rph8YltNZ6RWXbQDw+QpaPqKRQHJKirVaqSVT+GpxuO42pvz0PiGU7i3aVWkIqDC
q65xCAvq7/gOAt0AqtrDEPawtH6aqihfuo/RannrfTUkPiCF+mBuvnkfkhRUBA3i
5z0xio3eq21HXA5NCELdss5HiismrwMe2210MO/GOHE9lIC3zr5mq2ufI52Nm1G+
XcEQrK/SdU+7zh6BV2IFXEnnDcGJgfXGOzOhr+vyudhDNE4df4tX+Xz/xxbf77eX
AZrjemV7VH8H/3k6Eu2NKovDrNIYzu/lLtQI/HRsEvP9VY1BsA6eRI73+Qs1Mipx
47RmZkeTe7MPz0CwALwoyrYT1O0xEXMK6QxC0H5TjdlivpXvF4qDxgwJeuxNE6lf
JHWGmwdkZ+HeyNItkXeB0qaTsygJN9EXhbdweHUx6bcUcsiuZKmUkcxpbDpF2SCm
70A+IRZ7KDFaou1eH41FP4LS2901fJhdTvmm2EdNVYymQDVDVpWU/lC0/ywjQ5Wm
N50am7OV7XMtpV/uGqEVukSnInaTvcObWw7nemigsO4+Ew4UW0gsF5D9GB/Z5WO4
vVA2IXMiyoCk+5r30W7QWL0Pg0wSqfHxrYekbGTcA2VJpWOl40F5UUH7SOPNr2V6
nktl0K+A1u8dI9QvKOXOPLV6q4zh2Qp5jM7l/0rHei8AHtlsowtV6l5jO6TV6Ogz
nEpAYFRW0Dla48QgST26uQ9hi/f3iCzVeq4aDZ8aJFxpoMDLck7jeL6R9sv75WHe
3gwqVzPuv2IgbvOV/gtzqhvVHt34spxwEHXEZBG1DsFfEE481ucgfry6sJizx18G
PTiYqL9C7ozGtaGxJEb6L9uU8MSxzf+z3P5KQmyaPz2qjx4rWkd5NEDBL/h9//tn
1AsZvsO8FVOZTS87y8BT7EVltaT90TUDeCAdbC9osxaT6avaJcRcuE5ZbfUaKqmZ
gYHk/HpGN+UOKoESltuHpxeXgDU2nf9c7hN1hgHPAcWCS2LJYQ9RA763SlN0fm2/
4hXI5b1iP0DhBCO9dLOJtCKYdfGlofEBSSuX/si36VExasyJbwi9cF7PrFxAAepB
m0NCmn5SWqcOIpopQC16tics7bjlqqoFmrZKWTp+Gfn21kXPUKKgFDQ4pXGwbauI
cbv/a02VgawmYm79j6Gv8CkqdlPXt8fTJBQhfJsjaBnkqkuN7oIprAU2e/AjpZwp
lL09jSbxfci0T79cr7k6KB1d4S+uqQjJN3djEnMjd/ojJ0o8evOcJ1EPp8od6Xij
u8FoKqm1TvNwe2A2OpB1NQX0aNZU+BNOleNolYJ2/nduufJZ6JYMBu5gmBZBCz5g
mM5QeLSUYteBpGwAbpBcgYzC50znHcmxvQIwKWJTeIu8Jd7RhTaN3FZh3kns+7ii
uuaZ2/3ONYLCdOGxwP6Fq6r9I9Urt0WK8RC+P1xLQ2I+vufUhYq5wDn96kaZ281T
zCvV0M1jHgOBQ1S/aJBGDpUGQxigjK21hdlTqevOyrjms+oNSVLCFNUtP6cGcaoW
GAK5RbirlCYLgmhKiu4flirec915kqo39f8pqCVovPxyYNAaQEaw+84rV/nQ5BGI
RjFHBzZReMrmvIATJpbXOXbXdtbi+Z2vW6gKXNSjm+s7WBGq1Wg06WLP1eR26uMT
jhC87NqDBWg+9vTugsz1NGMIBCcP7t2aRPZ/aw9b7R2ezgX3/SlUP03QmDcmuVUj
Jg0+SYIN36MdbUm/ry+VkxXC3IjnSwddM0r05tXAJOixsrMtERuD3fEJSkllmF0C
7s0bxRsVPR1oNOXp7e7q5W5w/JFDQeKv/KKg1Ioj69jySZKcsfJMDcKUpDHcfvEe
T26S89IAMBAbFYa2eqQJPwgvX2S5lZvj8qGq94jZNwv0BmcXZGeC3z597dK96k8N
jovPFoErQCLeKIirBx/ET2ITUqmryX2kJAyFhfjui3AYYePV5LzLNTdP/f+GlDgv
y0TQ1Oy3SJN0RzTXh5VdakUpdwC5LxrtfUEekEpzqyRUAgzJcXxEuEKSYnkdSjG/
Ktd0Yiwm2QNlGhYuXZ+J85xqad3iNXFami8EmEcutuDMwPUIKG67xLJTI9DFX3Zj
qeNEePitgH5H821GRneGRmHM7ngERxHVurmvwN6fTgZOcEiswAOA6Wr07uvZxgg9
b5wKIMlDgIGu58IcFXgB7lS65inw75QXqkmwPbRgVeXmUlTG/x/q5GcqjvR1ZxnI
zFCG6PPVdtHoYUv2FtyRLmRGtcn3ijiTng4eXQNtrnpnbs+oifGZqJmVe0OIwfCo
jzPJ/FAa/fGGjow22szowt4aIU0jOBAezuYooedbOGUGJC+a+MsQducO5nHJf13E
xGuk8EkAI5fLMTdbLwm+EhsBGSnwpnsx4ZwRUac+WWVXpe7ZTYbLuZZi4l0xF+nI
nKjjyjcbIRZm6Wk2K8Eek/5XqlBfXrj0ZRc+VhbO7cWswrXdguSnxRkap7/vALk8
6IXN4YRdjukKyQMkMNPJbH3hCglTVgAhSxEaT0wE8QOwh53Anugy4rk0tTwsu9dl
e/e1eZiiMrX+YGZSpleEappGmEBvmci87aivrTWvyC5Bwl7BQFw9F2Zl4HwShyWX
jLQFIgVa2PR+tJKebD77CVJIgyL8uJWAmm6VHABqezVVQHHOe/S5wbm96aCxphkl
iWh5k+vFHtEMwFG5ulDUN7S81EUyGwExvqTAebtXyQrX1rBnCjZUZ3NBtGDTUh+N
5xx3oEmJYxtjSuLWq3J/GhE5OZgJk8BlUwgz+ey1bStGOquAUNreyZROOmvuOexE
YkEzGhZc4a8y3OjAzuP4QrwH8bipFYKQ4gcvCCpVi8oTtrkXga4l8HVA3H3zR6vR
ABmoNQZQ+ZvDeXTIJqebm20gGLaQXe+QZjJy6gXeClkBGOLy/QNaZ00j3ntbAX2O
Q3W47WCl8ykKOSaP81ojak+NyIs+RpWaYtBgQlpsMdgbIykAXqazm8q89R5TOta3
cDQRMNnrslmJb7YaT5l8e6qUZwy07/g2+1xO9QctP0icA6g028ozW2y94p58nvFP
G7c5p+uSDcXxkfloDlZF5yFmpU4Jmq2LHRm/DYrI645ex6o+jlCLeiRYBMwYPec9
34X42UKHOLeE7Z6NGWu+YvzOF5rmeqhFuQZKUVrEV+Qc2zXz5z7F4aRcX9wLGkX/
sPASQOkl/jSlOI/BDfHGJuRN6kj73DaWU7JxQroQ//ZGEc2oXiYufklip5Cu2bvg
ZJksTybl+w2oUMF034weWV/i9RpT5xH5HcSFQOH5NRvfj91edJkeaMkni6yOfc/v
K7tgIR0ZpYA8BTNZrkApCxcUrcHV+EzODEJcRiA7IFKxBvEtMZfimvkOKKBhP3R0
ncIJr3NoGYt4XSMe9wl9bQ2+5RnGIpDuOofbdTWXDIYte9GjUt7p4+FY4FdD2gaE
kOa9lb/GiGk0Xn3O6dqEsGwLP/1V4npczEbrkqDqURo7vAQQPYGzAYv0AMdwPNe0
HvS77OZqpBNz6swAEVPBw4wQMKmvsz0srFj/QmztQYa9fcnkofxAkWjUtQslkcpQ
87XohXklcyyjBxJcDsZbSnD8ANm+sYoeVgNjD4DHKMI51mq/Bu+8mf+PoEQjd4nV
FVznQF0DN9Dj3wImiEt8G9lkyQK8Oh7RO3VxO5GNcwzy25Z1YalxOw39mobaU3Sv
5HXCK09LDp75za5+zbscsHkxo4iomOJoCKJMtO/Ti+u45YpdzfqLtLuo9BYeI1Gq
09bgFnkUeimNi7Nm/9V0SjUegW+SZAyQ95VSGm+21FWq8cMnfLnnjN86iqpAB8EG
YjAfC0RtAoOReKA5cVJxr4xNf+NyjGvz6okSBx6ozSkDLx8+Agt3Qo3wSIb0yJ88
bZMC9VMtUn0PL/QfHugG215Q+CWTzPOCfC+KgIev8K+Iz+SZuCLNHrOxBstKMAlQ
vODz2u/M2NPrSOgwzfDqKZjnl98fSFwYHO0BiDsPJ/snJYX3ihPiV/jpkmdyQqnT
K3PAXZWwSwLinxvVZAZNdaeTWn42cVnG4ZJ0hh1+zBeGakpgBaZCyBO+Bf2HDxkJ
wmaP33QV27ZAAMBgEi5qbLSk131A7Y0gQSr12yIriKgsS1+2oJkVRGZhlYYH1je1
80N7/e0my1FoY0dnm+PjIg8zDNUYrX8n944qY0KakhtHT0qxMvfNNpDXM4MyfqCs
DqAgZ24fKR8UJbmOwErMI8S62JU8tBS2H8j3462lpCO1slfQI+SMl6azh9jdM/qa
3/jGjOBnLx113sVsL32Thsi5UGPzQstsfJdMy03Ih/DtFCnplTU9f3y/NR4X7U3X
bpbmghPkV63Fa/Ymvge3cnArO47PdJt6e7uIfbXxQo5Jp1/mmLAJUW5or1iSEJfo
ymQrlTeRpNYOq2f9RC2JJu58nWE7GB9llhTADXwRPBLIPdmzqtFw4S6+ygjg2GdQ
AWPDXtYdPQVSBIilyfoHyVeb7RMG+g0lXymHDt7ldyN4ZkBmt5y1ujwvwIWtFR/u
scCHdywwj4giPeduR4naTcfX0POtOlX0urIFJ3jGhMjmnprEHvPjwPcMm1jHghKu
HR8L07LlDoAW3ysGpvb26ehEl9LLL6OyDFJuM2Yp2eyWiY1mm7Z9sheTFNyXLjnj
FrbCXbXYzMurBMOKy2cggoaEEeScJiqsj23qasIBqsewOUCh5nAP3+M/5EkX0KKo
vodnWUJrXMG2cUd2LZHeljeSSEItIIMlK+VmU7sCo2bA7Mi7GGcUbKUsVZXvOoZ8
6czEu19AQJ9+poVxRTEIaXDel18ytqYVLgZShtmO+07xIN+gE1vGAKsaMb49rD6Y
udMKOvzM+HCjsfK1W4Ptxa+jlUoVGYHWqfoFEuoLuGz2gAV4RkUesM07WUlPmw9I
xquRS8DXnZMnKtCnb/JtASxuRZIJDyU3DCoOy0V5sTFZWNaHlVel/gVnPAE84T26
SGVsRRE96VFssWtefiihqsD3BXd2uxiPVoEoMWLCraWG1Y49Rqx/U0kr4/BE4Yhk
dX6ZhfNjt4O7pk4oMsdeoKhVKzDLRflDEx8rcH1Yv5uai7cLV0oX9q3AT9CFu5vm
9kAHkny9PaeQd3iqLkiH4GTNaVCsSp2ADjDeHFMWykTxL60NpyPNf6LxE7Uzt7Mv
Kx3ee/C9QPhwY3zUE94uMLog8E0CwhMc3cmuNjbW5Vbmx9sucEGttnJnESvKbkTd
ESvLe+BEey8Gq7Cv1ZZaFTU+M2RXgi7QeZWqfc9JJc0uc6Go6TZBHKpVBf7InkOV
kNOYcBscwFLgwcmFW/pmo9PAEyQdbqlLI6tJroEHKf2FhdCo+EMDyLQJJqTH6j1k
4cC+7eiBNz+wWx0lHFwuY/Ee1BnQef6+I4kJNyuqmrq/ZcnTzrhzu++iSUdoUZR3
zCdElNTX2MdEo0rilBzknrYnQXKwz2d13eqNBrt3EU949gsWxVqQMc1AR0VOq8/M
uLVoPmeO8qBqzAJOoHYJB7p7mu8suQqix+vAlGdZiU2hbCu3WECQ9tnjBybZWMjg
X4Hv0lWBKhPXhNtRQCnc5x3DltUf2zhS/+PBWdTIHieewDR4/jYZBrnJKbJ9zmNC
52IxEpzqKzWPOKJ6ickt/Zb3Eu9fWSaMhbYrfqUuC82wEy0KfhR1+F709xS7bIYa
lmniUmPjnJspnu7xfeBRiycjULrRsObBPsPK+8kvlDI5FAXVOkCSAZdCOPodTUK6
dXZJj/Jz+ac4FEl4L0RGa6IePGwK1T2ZAarNWW5KFUdqJpF9SIg3B+BCUik2fE3r
VuGIf5eD8O1jOGln9dIN3lfrPe81UveiP00ElkG6Nz9tS+wE7Du9GCTi7SRDCNRj
gt1s5GkaWM2mSN8ObxbnnPU/dDBvKPUhyyv5I99FqhsctZUSsl028R+FI3C/tWYE
+ssG8dGH2Xvfi5akyTUcCzaIDXmZdGFsa3phq1CvyRPjq/mteceQsdo5s7/8zEWi
yEZ0SF6JjglbDxV7MtOS56oxnvSi3ai0HAWNFW2SXWcPcNAUXxJJf3GHAJ51ML3W
gcjK6RGXaceM4tqyzcQPpA4HYlev9JvUBZBotoCLanC+fqd9HyUO3QSXVhZfJdP1
v7vxQ+0CMKMrw4sQl/qqlYGTGslqUB5N4cr9B4xgjek43bc5g9Tz+istt5V7d2+6
iGdsxJc7Q77DevSRgcn4Hbsyww6IExSgUTcdCD7i2iU6wgRUj2k1W6oIfW2Y7Im9
l5vRzQ/BLazVE00ecvFMzUieyxgnGtSHvjXkvSs3OSo0hQzui1FvLz4QILG11e2+
KtGD4r1t2xtjwXv23tYwKfDCopifcXE6kFasncWURFWZoEdf6/YWjaoF2+Ng0BXc
roV+PrVW81Q27nTi+2OhP27MHvrBOvD5yrGvcLf7Cow3mz/ufmLQf4o8at2N2NVv
YXTJ7NQ6buMyhdGVtUYRJ5A1GrUXRqpv9PZdTSPXrUkIrEIQxL2FgU0IH5va7T0X
WQhTpo4S6Urc74JotYZTOqNLGGTqGLMTbC60TMx7eVfL+C52elXLSaS3N34JtIbC
s7m7B2KS/Ta2tBdaAb5WPCnMc7IX/VFZbWh2iK1CgcZDK8rB9AmWEFxLFHqy9VkD
sQkEwuy6rMx/mrR2TklkYsQqFOrWqyS9z3duf33rG9O+f+T1ysqqHqEiv0Xe7VfY
TKV+FkECNik4mMa5mQ6I1H83gBffiS7+eyPHvWvJjs/hvc5Ym4g5PiCynQzAnZ2y
n8vhwFzJfLWHEMVwbhd+67TG9RAGoPzVSUOwbbS+j99NXYF4ie7cNg46M0/EexUt
JXAO8kGUJ8hjwxN0ZoXp0AzNqJcRgA+GcFIqcW5c/xXIlcJkasHLzX/Cki96ozh/
40AcA+4N7E+Op+5VlFSzn3gxBDqoyn0HoeBAU05HKwoDiC+l3bSsez64fMhic0x2
zyh8Aiu9CnGKUaOIL7ByDVLwDCFgpILYkt64qDS8qX45VS15VCTQBCr6F9m5/CuQ
Qhk29Xvs2zU4iJMff0MPDdiJSdkh7IAxC4dXuo5NEwYOH+DUyjeVWqIs6O8JNHS/
GQwt7ykM1hbN6NIUtR+o9tlge5YouPT2wEn/yzC4oiL0pnzx5sVUPEHjZEeEw0sA
n6NUpPlT6zubmc6w/OWFmf4SenIA4ojMXIMZhHiqH7yZzUMOAggTY5tkz53RQhAL
U8iAB+ovmoh3c4hh94QQa4F3gPP0Ut8gAldgOqMM7LhG5UJuoi42i5oisxNt3ER2
IhAZeOp5bxeVQA9l2hKQWLTqDOmTzBx2/cz0oyPxm+Aha8N1ZyBkNlS74Ag/oyTe
i9L4jpCQ9Q2oEXIGZxpD3+Y8AMdOs+E+BAQn8Vp7oSIFiomYrnrZdZ+3ZLS0D3WX
GNIi+ImEB1kz4NRuHLlMjkhI67L0koXsw/cepyZ0z5u/XPA6XwPtciD2XzRrHvOl
a7XUBW0l6TxPwwI6VTLxqqHRP5xoYS+d9qTDPq5MPJL/nq11ExekeqbfzKGVa1lE
Rh5zZXhRMLNEg5ebhYs4pTdFCmR+x/kXLV0R4YDp2SN9InSpzRt8mLh97yGSSLdB
yK9DOFNE9SYkAXCOo4ngd3lGES0raxaQpbi9jCDSpHKjyjveKCuIvZFaD2S8yspx
mmqgHwbZajX0O/SM5Bp+93tRtq8HKZpq8KQ4/Q4E9YCbwSA42Z92hRDrGru9A/ih
/77Zd80nC1im6VF7aCbSalV8kzLaAf2VzxjIGP19RO/8lvBGroZnk9KUOvhPsp6m
EkepirYHdOt9DaN+AXf9NATTt0bD8JWdIggD0tFaNXmfQ9vQomeJOpAhdd3mCcrK
K8+v0h+Huv9rMpRHHJX+Wy2UFedTncc8+rsOeUg7s6LSoPVM3Tj5BBkWgXirtS6S
Z1QMqFlNShdGyXpdsy/LET6PuuTEb1W94CAT9V6t8jbKAfszuK8eCpzIXKHr9ai9
UPoNAngED0YGBYaPPDPLVvl0ULpIBR59jPlT/kRrf4C10PrqBDZNEU1w0s5pF0xo
KmWADLk9WB8npX4j2CZcOlk9edBsB1IFaYwZdfQdb+4SHPBQHxe8IEVag8s0Kqw+
ODc7lXl/6QNzqnsdT8Cf8fep3irMhKpzBGadHhViFF9UTu//HiJkK8dUX4PKh4Y2
rWz4bBAMtk1a9dqbDQn2x1aG3aqWA9VDgqdH7HFc/zcwXCs52bj4L4ptYE2KFiiQ
K8/ja9xersc7b/BXVtF6XS7hwjFRfo1uuOyatsVmctc4JQF0qDkiA8RuOx6gIXig
TlPcmxgzdGTBCDINFgdKJOfdCryApCNarp7CbyoUw2xYX8rb9C235H9Jjz1buxlS
qEcn+chRVgzIoMLYslw1/lXub8QdRLgiEduq74FjVDLKsbcPbpY3VH1qRrXISdFC
M8SZrsyAHTB+FiczNHwpiQIzsGpYNM/HMB2KOBxfyKBoufh6m20hl9UgpeOdjiO4
erJO0RECOheZjP6TwHMdMr7TmcfF87jVg9Tc4zTyg4Stzb4pTKQ68SWAGdgHPxTC
53hGhw/GD9skzKIn+G0/VH0WxjZYp4iQHzdz4Zlrp6Gvfy3NK93bETNZ4QqcFBdO
6WFQnKpOkQjR3rJa/n1KQJHVTVNZVzlwUUNFL/4XGmycywaW4K4jO1KSCj/YQ/4V
Be8mAVAxXNp5K8bntX8NlN3zKfpxukWUwagzhBtWxLL3/f1r4ohiL1wPPQ0q31Mz
Ri11Q/+7R9zRqUBlcITWlwKAp9gvcotWF7pzms+YVNN5vjaVJWehAhwlBP1K7LWl
CJeJmDKMMq+8v3I7S8PiziYSvCn5BAfDOp0Xd3GEt1xleVsi4iMCw8+bTdP/qGzo
vaitILt4ne8zOpZetGQP/8QSIBnRjNhz/hR95+8RlaTNXVnBs0MLjW6lX8f1VpJo
yUB5YiVLXKRIdafy5Mb1ikTGIyuH+jeGiWpg1a8WMIxm24lUTF86nxlGeGmxpUwA
U/U3iqny3WClgH+svZsx56Ywmd2td5LhL9Odp28rtO+92NEE1fMW69tHQDFkev+P
iuXmsE+QRZFI8ZvdqK1h7XIzTsrYuymQQKTHOdcZ0OJsAOoPIk5mYt5Pmg9Td8cX
W8paxuykTIoDTc14aDSpZmlMse40HC0Kg9Oe/sMIRhklAWVwf/o724AydR1wENB9
YrPYnT/aIcsDMO6fW7RH8MLdPqQ5DRsIg0wFEwADQDPcjbZFJu7WQZ/1aKBQP6Sd
xWHAR6A31r8Xeb/QJEI0/GpC4QKFtr5q/I1+gO69s50Kq5vJIRDsOmakrkOXZ4fc
gLgmjnnWiyBXOfLo5wsuWFkKDlApvdQEZ+M927vt/NjC6NoyfKw/BWg0yHANfVFI
cHpSc16xIFE4VjBtipiIR1eoJxKmrX0ZBAPFUIPUFsj+lq/sjx90sU2XqAWvEcho
/NYeTx04wvA/NYKF2Uz2dcZ0jNpgZ88s69+d6KNf3C9NOQGpRe6F/Tned3/Jj0Gv
ZF4icfi3dJtVThnVPOztuwjn3BtQMO20LSUf15dBENRppWRlEKqyZR+E8PUQMdyt
aSmKz5aLHdFwjkV0ZWdVVQv/5JG8/mcrtIAF+Dq632cTS9jLXeRxNCVIS3elkv38
wVs/wWj3I5Ukd+o/pHiolUp7y1znencNU0gsyNKc8IW64zmppj+oq4KBHQuTAp0L
KqTpibS+/B0gUXS9Hlfdh7pfUJpnLvN/4quJd1WmaivKYR/W/Vx1B4W4i2SZA+SQ
ULsM3/Ql8TmwN7nVFprLZJivxiFK/co58DJ4uDqqS/cgUS84YxH/qznVMLIPVx4f
JkQgfGt02fL8LPRgaEeLDG1vPiQAJePtKsSUXjAG9zPYsSIw/1/8MjYHlvdH4gK8
d4DYtBabIggYX8wATeYEbIWJySlPE4wUZobWagwVFIkUEwYm7j4O1N9zAA5B0B1i
WJ43XFMaKrSmOdMQjn6aj9bjZwIVh8ORkh0yeP6WKgOnejYxjkblmFaBXmfFYWs6
1FPqkRcJ2qK393xQqNFBxq7PYeZ7MmamHAryGAditnqFKsPitgURHUyy8IuXlJD0
3mFaoSsNF97hMgofxI9CpHF1MWKzn1jmZu+JfMlplAbdYMCMva80W+JKp0ZucbFE
SBq572Rip+2jYrdvJdmKwQfgzOkSzEyuAWmubGuRebzTv9lb+hIlrLOAJcIuKoWg
OTdlzCmjvCSZfFfuiBb0R9nliDIpkYCfGePZsN/RHV+02jBts+xFUhv+xN+oNE/o
GJAVipKAKKM3loIcWSmCpXdJSl7KLnqfE6Ge9nEJseQRSPNXZgWni4rcb9FED1Ph
SoQOusJaxBZ9ZgiYmgeSOGWpig4aJm7TAyxVJkQgM9tYtqFRGSHO0jpuLvYKNDmP
DpSXWlcg3jQYYQdki1G91oYorGFFJgcxalyWcRlLfdeSrvbRl21sRTV8UL947PaY
LI+de1NtN24HhHK+mD9RJdy6VCQZqrKYNZseD5PkdKTq2NdfzuSS85HZuCSuL5Xv
TA2qP92rbM5AN/3au8gDIF02xwP9u1Q5DwdQrW7Vj+zmkBPJEWJmwaKJJeT87RFP
Tm2xyDuiE0MROSrJ+RtDfKiJJZIjAvuzdEEqLhDgXh8C2AttC0vJIMeMxoiQTsT+
Pe54xxqieUg2Odah14goOqmSilZxb8Y1Za4+/WMXoRqNbk+yZQ13uvmSYoX4sJJd
wITNWBxuOkbPi+PvmMFXQC7iV0bgW6E2xy+r2OaQufHrCRcYdmwesFtc86EZVvW3
Twbwjo4U7D/H6Vjlyl6tYBYJ50/zxy0g+T76y3on1skSnDPT6zQ7wp9sE/R/1bhP
LJSpk73TPjL+CF7jGIQMmEKCaFlv9VRZnzj0WCIb2TzZtOXqFzbp2r9bmFtCOp6e
6ISRG3hMZKKlZu88l2NhkrG4e5R12IJ34ZhEkhwCKPoo8MbIDOE/tVxDzvPuUzz4
YrWqGAHxJOM+ZeilkpvrBcKScq0hMoobeQ2nWYPX9ATLLQmEyjtWGp7zFdhC8dwZ
Q49naFPNuFW92yj9R7esrhzfG0xFJIfSYRuq+nvYEdLmwLXX4I3Z0mSaT/ftCMUn
3jF+Jx9iWk8dTmLR5tyH7mcbUE34nftC46WQRVGcf9cjJ+D+xYpFnHA/7tAn5GgI
1cLoy4Dlo6mlNLRi6iuWNBdqwdasSZMRsxLCp5esBQp41QGopov3hkNq6pHz5G8V
Xv57vhwVn5Ky0THXGrwV/jnflib52C4dD2GTf2DZFoqOq52jDv1MtehBkhepEyml
bayjHCX2vx0E284XE1HnkoRb+OgMgB2bbXS0RW7qwW1NSOVWIkcNhp0pB2CumKHt
4lN35vrRH13zbPAABItNKPFeGZsNrx5Ce33hFg1pc0kUwERYe2SSi2g0pF3P/SNV
URDfAqjX681oMk1AfnHkRYRVFFsPuGMWzRu8XH+2/ARZMtI4bPHcTq22vlhR0Qt7
ebKouJPS5kxu/ZElhdKzrX9B42JwGZawSuebc7IqPi2hr/S1Ev3CQZ22flUPSNKl
U46tUJ5piTAmUOn47t9Evv5YgS4CXhN0+z4UlC5NwVWih/gfIwv/KWb8DT/b13qb
r8b9QUQhxhRAH2kC1Btyd7mRyn8WkUCVwKS6SrfE8JKk7HRgtoInvnxa+B7O7Jpz
D14+lm1Xp22VzWFQXXPnPiBYXu++KPdjxVuFqfz1T4evQvjve/uR/JS/TkOz8XTN
JvnFpeGhy+25Jle4xErxyDYDu7HG7B5CzPG6iBgYfFK1ZcSNducEuXRP91m7qytn
FOO91z91IkxRPpYV7TdgRcjhB2a8ZDUhgffzNHGH/mftxG+L0MqmcqcqqtRWJVQC
SU1ljoTtG83W42YOYgrqRGzr2Sxd/oXxqLytp/DhZsa1MSud5/DBbWuAQEFxk0qT
VVCqnicU7n6fHz9vcX215MDCPUNVMVdzBfmZ6s75o8xXSlZHJ9w11JcqmXxnTjW0
91kPdw4m1jZdfP2XtvrxV6PhfTzzZ3/RuoPGwMZnA3aJSjM/1zX5uMtnqbof/c1a
dx9B9fUNJCl/MRPmfG8B66L+VQ1R/1Clo2+Z5ZmhID4HrHtpXnpyGfr7b7eD8IP/
vHQsQ+6LcXIgt6qZuTlRfFXg0lK0h+DVs94rVk/VXD+JqBeAgzQtHdt93ktSddbp
laNljDAqBinpBSEaq7pQ7qR74W0D5f0yqBTZrud7BaHHVr4RQuoe8pHIFNN4J+/i
LaGuFenDTiyploQU2e4w0mqt1oxttnSPB03fuuKdO6DTss76A4Q3DJ0eMzeF0T/V
HrtNNn92Y2q+DXomIL15Aoe/FuvaTGoAA9y5GX708csGodEdn2JYlu5lZU699DtX
WxbYbdvuU0KZRy1DdFrHj8Hq2c2Ea2k6UkM+Jl65PIWVcncV7DEVqm2D++ADxFvc
ZchWf7ke09ez3Zi4M1DKMUugz9o9UTEPjpB/K3Xrca75rB1EbJsmk9moSvpONkwB
r0PSEpDtz5N64cu4/F9pZEmCNqHWiD/dJBk5uHTr7hIlNS3xoBqw5QDiTTmONmLZ
1a/pvNa7/WHhevIK3K5vAr7wVOgLyr0qbhlfQIMVjliBRKnRXw4BAvQB2YlYzMVo
yxe2A/fDzS4j9e6bffxXPfJaZOO0lV4xo/Hg0Uz85efB88H4lxT4e53helKBu4C/
IA6QtGLTbOchqnckDDPsfPLoMjNgkIYsyNmS3vvLvRjhxJ+NOgXCdisRNUYD7XCC
j9ULDzJoWjPbWmqtHSXEyzpUAgp4k2Orq34dw91YRkLIz33tv8z1+x9MEB+yx1DQ
GCggtEg26MV/BPQWhffI+UkKtRSwRBQj7WDdDbVHHiyVeRsPpyhAE0ESYa7OVDI5
bBeb12tEWoktsAvN4soFlhcWD/XPWIjEAnz0+0AdnYzG3QDzY+xcJnpd/AAH/n0r
l98xo2AmLHPqtnAtzVPD3noxAapn3FIUFADIJqYyeUzfIdJHvk8PzUixhCcIjp1C
TXWfSMmoFuBWcC77N6YTwPbJ51JTCv4xOtC5wTu4InRp2cWO55kV3+DkErirfFUj
Shy6Tb0wl3nqUsCDmysP/DdcsXFaGKExeEeLlAZ/9O1OeGHm2MRAktmVFwCbtdqk
DbCOygPMtyCYTaZ62Ky92/P9zoDcdeBq/PlSe75rB6AXPuJPXWycDX2LbYZbw0mq
xE+TBjM+IAxTwCcxcDkBGLPrN2eh3q3XiCm+UNOZUsNqQP8+hooVNN9hppst6rm3
nS54jsnnU4BwfPvrQ454Y052zGss/RU3yjZcb0s2rjlfZZ0VfL72YTzlVcjrIKq+
inpm8qB1HRH30UZBiyMcCkF1Fs3IF/0WvMQ3SlRHF2b0GW5cYGC3axqoH9/6XWn5
3R2CI64WkciePgt1VptCNEAM++uIZPr/EBsx085YrwptCAqG5pLChE8KdBXGcnDl
7yd+/81H08ZXKEf7HolXX6ZW4hCPOK8ipSVMPxhYHEuMWOcc8tbjw71Y6jpHrtVB
U68No6I5qTX+nW+gerVsCqSQBCehkb7m0Rc8ZS26cvgqG2DMlRrjFkIIOKWv7d6R
aW3z4IAkTRenzG/952eMEVPlAHiNg1cM5hePK0y120qtmoPWp8Z12JpsYgxp0kd0
rtgHmsJT6Vv+QQSMLWhDw1ve/jp3gHrLBoXXXZfVcffiizMGqLG+8tdx21DVN2E4
68Xt2xjpAp9Uzp26kAx3Fz7EVhXE+6xNsofIMkzU57VvbXAHtF9Zg/y81GghZS/e
1D5PKjum4sf7kom7hJasZUTvvCS3xHVDeZHJpqr7P97oSmoj7hZtHbH3ls413pLI
cOG0ZI/GskgjvF8wusECA042oo6qNOUsMVki63VSVF42fV8DHtvyiVy1xCVhl0mU
v+i8Ea1L6BUhW6IFCzgGcIedV89Mid1MoWXXUBJbEwrzVO8RvtBjEtupC41V/M9+
KYExwHXnagOfBvA93pBtdfZx1YSJrKXNbMjKFF2p25GgGXWmdchx7Rh3RUzKPQvH
tNzQ0yPupTsW6k+r4IEBPExYvSobWNiyegjuwZN4xsfLcorJlkYNw8N0xFZShDoh
RKv1k7UlJFIlg63v8RU6kO2hHVgtJcfx4tyZ+MXk+9hz+yf2e9evbabth7cWrTHf
aZmbIJ0BvJ71Ny3SRlRTngGD1V6bMmFKrBCyv9HTmLvg0Nz3QlbtugX8k57fG8C/
mXobyH3uMnx23FP9KkGEkC2T/AIpWi8o0mJQ1Q/fKsN+CXqbFo2JtZUoFDA0b7LH
lQp95X7cw2Z2MK+9dYFOYCKRyfwFnbfhNAZApUUC9zO4ScWRO/O2aGGn25nvJzsP
Ak22Gb15dsRP7OdqVOJI9VNcQG+VcZVHWRw4T5w+fnSp2GJl33rIH5DtbjXYzWkh
1AA7cgr47FAa/ccQb1ISDpFnOdocdu0O6hkNPw8VXE5kUoDN6vEP4JOSTv78VesB
UB3hYu4ox3XNZ/hYLqJ1U4cBtveTBgy8yf1MW4a2yQFIki/zXcrxQ8cNvbzbp+Bs
UnMQbMHWH3vIEs8aaY6gSLaB0mU2PFPCFTYCCCmaLH85Es47XmwYc5dm1c7X9G0G
VRWv1O4HWGSUvSI+m5RPN8uhbspsvTh+EOigQrtvgEaGy7YVde+fuxJ/9nXuBX4C
t5N3ptLbcDHYbAnoHBzJ/YHFVGA/CDuoCxu15VGPBQQ4esHXs14xxYThZGfNzV84
0hsTRzew4cjy0v+cGa7lNfUyXhYmSbkSbEuXlYQnw858UV88tU1Nd0BGy/ZeEXi/
Ls0xVkn18FtzXbL06Co38PZ3LNgO8h+ck8dyUCMdhOu/TU4Ed/GiuNe59DXqrKel
lO+1T6XnfrnyLdxUEgZpKfb4Zq0CYdooSN6c84pUNX0Xi1TVojLS2c/vNlovWEIh
Ybrvh+60ij+BeLpQZu9rs3cmvF6wHRmb0UVVsVDpAUaM48ZCiYGm8LeuH6Z+vaIc
8wKbeqGJUJM+MGCz6Z9eZ1jAHzUo+Gd3EIMRE9i6tvo+TgGfcNvvMVs20KlAQ33v
gVuKci0NHi/krJtSaHd9IqAqvPE0RoIN3oNRiL1ZZAn/j6FjcFRIOBKJS6S7GuP/
EdvmW0LICn3w900+3nys0CRKaPoQ6qi35htyqXIqRv94ymWSRGVxT90noljakSIl
bZFRlGLK88m6NzPj79t6gqGrF/Pxpr2kl2XOs1feHG5dCY61OeM6xS49LXwx5G+V
26LEUYxjgfYs1iaFt6zT5t9Ef6mEjG6F8gpW6low+10vm8QjX4asqJm8g73/AOwr
gZuktIoUfn63wH6+hDWK/2GP76+Dpo1GjXIG+1PdQj7Celu0CF9wj9BlN0NywhSB
TxuBxMDb/OE3BUUByYB6JU2pdKMBKlY8O0Ih+kzkHq/FPCcKWsRL6UWkt69iMYcP
8+R7gg/BbGVcSptv0fy37qvqDzhgj0W8V0ITWNY0z/tIm0HsNBnOrKmhibjB5+NJ
kKnHQbpjt+lwUQlP7wZOM/eC0VWM1qKqTSn/j21rMGUK6+DL20PLx29RmGxabc7E
7Mf61bFQM/EE+nAESwEYX0EWIkRFzNpk4HnsX4sklPhCA5kF8nyMIWxLlm0ige7T
U4XzJfm8ocjhQIuuhYTtcnJPIGioZxxOYqbOV0+HDEcs5BnrqIscAlYKbMSdAxXQ
8o8B/J2f64OeTxO1h3y5DSRDg1WmEeNNJ4tIDTVioFAnVlKylVLQs0taZvjNg0Ng
6jje8PkYN3lSwiz2L4xZklYIWAyI0XoTQPEJAxX+pMHA6rl09MvfI9nEfikZElgB
SWLUy8MGB9/0YuSDlTAOTLmwMIYifohi7A6LawIq1LNiOG79Vupy9Tb8vnOozIRC
OcoCg22kxf5StH4IhYmq6FimmvYLpV1lrf66VRPjULlq4YvIRbYT+f2QNXgrh30D
t/RFHnUdfQayFBpRflAzJ/q0JpLbtUc4WzO51lvLaQiLkGj+3wOUY2baYGEFSKLp
tg8HCSRqWJh4mOkemGlH/etlNJVodgiKM52EwLFSOX7+CwkqT8ilEzWbjSmG/GlB
giluA4m5rfuQrRPZPr0LLTUniCSSxPa1r55y1SlkPFtB5VlB4O8gSXc6N2GCGVtu
1k3oohrLHMUvejCgfbkjcHI/v94+lAkgSiy3HGAI+3uDMAOlKVUR9P6Blk0RIx3O
n58fTJKlCc3NMxCUdQTVQ/1dRpAPyyGl/YWtTop3m9fb0ZAvFPrBNYtb/KAgDbRw
ZKxSLtx/1DtagKY/+lQhkW8mVpUX/BxKlB7Tg5yTIMttY/AXiNzQ470GRYb3OF/j
+KEqpydJK4W9DOoUPNdJDmlBTpDSrIc0Hr5Fqahb6U/7pP2L2qhdaaxGrmgZFDCJ
ydjm2oYHJzodOOQ2zCArySVQZ3luv8M7AQxFkkeohXmD40ATBIdsKJpJ3Cmwd9Af
4EHf85gGNgFDrlNd+zbne3p6n5NTg7NwrHpU3h7PtOOoX11EYYg7bLwCPeIN4+1q
cGCPPcWSFwxtCnufPfFDywWSv4sx/sBuq9zhIixtnTOnsL2iVjJgccqAVAwdqHzY
hWeZHLyMDrlrFyTC5PXlZ4ErqNOlowKAz4rG/9UXdkFWku/ZCp8ljGFD8kpUh2CH
Qei5UQnNovT8LVQR5/9z884v/e0fMAEdc2ZlL0ciN7rharzxMcURTZqunsDfEQ7y
mKdCDnJFnhMFBmq5gHOEdI8A8D64knmx6wd2ul96JsYrXVFjAFBN3Gf9UaVF8Ste
GdD0Pzq2qKrCixEJrmVwiipfe4XdVCiG8xfBUuyBtlkZt7iMvipIvHn06022pa/u
CMupNvE/1jL9q1COpDJ0tLUoQPaLvod2h34D9kZWsIjiTmYNKZzVlNb/wfqIp5im
YbssId9gyGFWKc/PPfOacqPhc5/UDlxgvBuZ7bFdBBUPPY1OmK+vN2oxWn0mY4Cl
6+ZYJW3hUBaMU9CH16w4E7gSthHKbjrqpeqiUx98MTfyba8j68H6pjoAkE32k0Zr
iVZ8pbeN/4vtbRT8oVlitXXfx0mcuX2BVZbpJGWf03vPBU+xN1N6jYoG3Gj3GJRo
yFUL22L8diTqRSwzqYhs82bIFGYFvcSbIoujXmorP4sabDaHBu9b7cyLuuEcE2/x
U1HoByjRQgg94WcC+8oLAHpkbprVf4WYgZ9WOASSYz1aKR5EXmRwiHAeRZZoHEgv
/P7OnwDH0MUnoT1hdBviEctYncQCj5jvaWOad+zzTRyrNaeIxqTTFaae9oQJEzWR
bf2F3Sqd4tyvp83GTe99w3X+qoOv7lUMafM0LmlE2SCU9+HfQvP0HdeGKpZ8GXt3
AzplJMz/1V+u6GLdgRoPCsxedQBIaTkuZEmyGxx+SttJqTGBsjmtam6x7JswhAFW
OR1NP7H68lAOTJWeLDEtPcncJnw1msCt1S694Glgsc2dDxEFvkVyX3GaX0FmSQnY
FZPMAN0oZ3Yh2czj0ue3Eapul/DZw/diIFhuKeT6mivajVfy2RJLeBj42vd/GuUv
mhfPmpqFsQBudKjcFCoW1Bg6a1w4bYPSWp8ICQdSYhKswys3Uy18RWaDWW+Etpip
retQb0/cbgotRpbuzsFAF+xo7DXh64aMzfY9QL/ATb7jxaORcrgV/kW9u2UOkfWO
23OsMzA2sbKS0CJBtf0vhF3BzBJWdM//wKEI9eXTccWdsFJF2r3tehlRGNEMrcWd
JxaXY4DA5ugaHc9wgNaEkupDWP68TbtYkLDI0EKBTHNnAfQ0Gas61yiJF8NGV+df
hjzrzVD2w9uhVT5dP3EqatxjSC+abx10qzQbBUcsErlC2XBaUCusvGBqQ1RZeDNI
kjvsz/bzbeVKu9YqC2Wzj4OshLuHLddx4ym2i5I3XD2qIu+QNjQ3OCq1chcUZIXy
4lZwLheWlmh0b8LCSOPBCdCdaOlg/iCua+r52RMV9bOqan+H9M3LOz2nvUiDbvMd
3rUQSJ+8l+Xz2hJKLQ82wjMgGMZe0pBQ/jS2n50GWT71rm3RI4WBUISmjUQCKWBM
y28rjqII7ejHu353bQX0ADEQ116yf4xFkJMzq0PGFrnL5ddCTPY1YdYEPqkkg7Lk
4GSPizmfzY3b8zTa3OQN3lx+t3uvXB2kD5rk1faiY7WnAVER5O64QMROZt1jZ0cr
gIXfdfMlfFWrwJ/tMsKNfQI7fSLKGcFNMm1v6fiuTu0a9wRUDdqjGUW7pzkf9BdD
1wGSE7LYnooLNDGQuk5JOUkIlr3kc/dnIJ0322dZR5UTlV4wqM3XBadhWzffGpBW
Yce05C/TsN4rAdZqMevKKEuHcRLamKTU7O0EFUyNu+tXDCDkoOUV2N/yC4basGg8
BkKcQgtr2fEVisNC0JBb4QFytOWhJhaGpYACC+SxEjQtX3LcZpXtk8J6nOs9eHEI
ivmgIBtOxdUtLnDNdLcPwlRrgG6mRBjFLa3VVf+UdZvUvDn64CnSPVxPhDHBMMvJ
WDZM2LZFc5jTayi4EWLPeN5rMbYfi35ObMlIYRJi+0E/uiR5FM7Ui7NhV+ttU/kD
D8bbt1PKDFnV11+dd1XGumTe9PeI7Y5SkhVZZFg06rU5NkYn892t4j2XUU76EX0L
GY19U5bqpliuPRlQeHAq8PG/TGWdYMGEOiHWWorU3bstq+ymhQcOyOYhIhsU4HLN
13YEaWcbxRxlaDJ2i58OgZHNiqHVSV+96kwh3lcHDfZAOw68FLxGESLbmasbXq06
E0UjFdM0ped+BPYXsg1nP6wpxGhCFX3IBfAHEoppX3AqXEPMk6uLCrgA/AQB8DsY
H5UgWQaxDlvDR8/6wcJhdWEEJ83/4S2Fp9nMqitoiQZkQxeL/f8ktUJOUVXWJ4bm
wbso7bDzzEM3/sPwB91jaQfgKGeamPw1X6pfoQkLPPhtIDq8HbB45zPF5ZM4noQA
l8+c3066NKihRZGZ3Ti2kxa9PGIRh1sSEdQhsx+6dAv1oq51e4mXZRVjq+7b7Dqf
00vvxILaPgRqFgbSD8BzDe++ljJBq8Uy6iF6gEz6/B/D5zObaQteV+4fG4bztJGV
RAcsVVzAqAiBprIHxETAyr2gaZyRcH0bYRHOQo+rUVIWLIUb3zy8HGw3CrM4r+rR
V09LO62wUF7eSi5fHE/6NfrFD7G9j/IA5Tw53Y9d2IZcuA6Jj1yXeAFfAIw/1ClR
opVO1pqoODAN+jD5p/b/03/9fXEKfYGvYo2iF9tlWGAK3Udd+K43qQak0AV7fWHr
jWI7oV9tL2fDeVSoptBYdnBO/RK53SDXiKTfcUEzyNj/zC/k5isEarr77Vuw1xNk
HHtu6nQlnJGoSJmY5I/Ru9GdhJGSdbX8TbghbEkh5r9Z2/iJoHaoNg3W3EgzTE9d
4Jm2C9B7AM7EQYA48DlxIdvuEZX6IpqnXpO5/DMboPMBKE0Vzd1tbSQwwHBKlSxe
ebdVW+s6+4tzf9H9FdW+BLbq9WKp+xDnzOlenwqEBe+X2b/jgXseh6TAFazFGgaX
Pvps7TAM0b9Hu9YjY+xxeoFsXE5+IFUP6Xv9uAqMujjZdXLOl8BTVWAohlcYVGJk
9z2MnYlBc7i9PaBg5z4IUB/7tql9cTbRpAvR7Od/cRae46HMeT2UWqdDos/OLM8K
PN85+O8bD+InTAcWjel550evzsa8vyVlUP3/91oj19UhHnEgXFF9rlHdOZPGZJHX
rCcgDKewsJ/H8jnbjLbBs77IeKavi2sf7WWeSO16jto0zV01+ohejrd5UvrBGxoh
x/gG/SJPVibpJlHaOxEIwW3NlqZZHYuQWI/8Y3h6yJIHaSG/osrKNpn28vSQkrWG
RDKuA3Fk610dbub3ARQ27r8nqCr4ELbX//a9Y60KWP7YxX5E7HOOQTaY1On4IdW9
yRlXgAN069qIxAlY2FG6bfPnedKUbZfdOP3Q0E5DivfT55DLZKYH4AlgRvRZgbbl
SWmD+qbKEyGBBK8nHWIfefZmOJ4OVi7bHog1IIQdV2NwdDRJh/yOH0l7zexlN5MD
p7VW4tB3jSAXhg8yZUoAZmKCtGfaGpQmDmj/KnVfMBPf63Ngf81qrl9AT6ferqFu
7WD7CCph0sxkzarJbYg9PWJlUcB/0ck0i3Ws7FhEsWQm68ujTkKBQvQ27DA9RxYZ
kpeBUy5858Gt/EQxDj2xNaIBlD/pjX99yilwmTcV7YPcixiM/wirt4FPyjBL9AsM
oxon+QynyhrHJsa3zQhygYKcwaZRwJWWZyrR/HdMDFcZAIEFyDKBJSuKY74IIbP5
tcgHq/nlaTuQODViRUJoNL8qM8/YT+ucFh3QTWxFDuNPAPQvQXcQBU55jP7yk8lf
lMuT7q/bbphQpMdi8YnNW0zCFilxp9WqX91F3TLETvhquBEJ1YhVJZpZGPhJ9ip4
LQPZICRtqoHLlx8glowr6LAs8QKapIvtzHSEuGG4ln8fpQWPksCAIcmN+U+xmfau
GNuDbkaEYhFT8xjpOuyNfsCjvUahTWjVFr5u15LnDpemrfDseAXFZLegLdezBv5L
40QLZkb7c9K2zGukHf4mlo2fh3Vcwq3fxVmmwvvFDCUgY92nuCTTMEo+4xKFHIQW
sCr/yMN5SPB4IJ5MHJDAWtZSjo3kLrBUENTrjBMLFSqPkUqg+H4tPYNDdujU6IhL
nTkwDHGvVHfvAHqNzQCDoojHNgqA0UZAsVvcbYfwqD4rTYyMsnhLjQuhsTrOFGCL
WYnJ3Q6yw73MH8ga6yAssgtUmsxGDPGOD77BZhRTlHXfYnLA/wHCPepjIsrajTJJ
/TrtN39+ZXQbM8O3V+L5RcvSNyRb9qHE23T2qDvIzBTvT2QWgbbFKD9YcXecY+DH
2hLHVBWSYVsgBDWt+x/WzNAjDgGSbBnpNqz/cEmhsi8s9cihwvBERRFu8rHqz7Bv
HAhl/JDXhkz4lfsoHW3oIrP8PBIrx8bFfO5jkchOLeCpPEtJ5gjUBmoQam26fhsQ
nxL7FKJN97lukjv88MCmsu8AlYMxlaMOZYB9Vj7+rEPeZOd5M1XEfGd1+CmgbSkn
CpqlxQw3eknMU+eOnPpWcK9Z/CFK6ik86mmNnu1LXA10qsTUA6BKHx2KgOcnEkf8
tQAr7aOy84pRt9PA2AjrceEEPN+ti0O0Ra7VcesscEqHl9XsdtNUnbSljt2i3SW5
RHM026buyZQp/z6cPdvjRRJZLOyzmUC27DB7gcxzniVNkLrrn7MPbN8b9NQWhF4r
u1MNNsGB88YVlAgt0N6gUnzv/ZpOU0lAQVxuWBRg0xvm7RDfiD5D4g+9FnlUYJXf
3YZgSrnpWqcXIvV4w7G3G3fHKWFznulcr2bP4+dhYQMQqjmlavcP8RX1TI1A5aIx
/QiPAxEAVYRMgLh7kKqIRzgv10FlSvbBRVnk12aMiUkbDXfXwJPangHMo5pV0vcQ
MfRg0E7VMfk+aGx7ggNn715stTJW0qeWCMwMnR5AshnpVpHtHIRwF6dNwA/p3TRn
H0f0lnIVF5l4AjTYQwdNMqeBbAazO2BzzCd5oClqGto+i88dhUoZ75yB0SUWfYpd
2g1bNYAsxZRczclkiKGlh/UXCOagWTilWNbsKNQnrFJkF+utgSl5bb3ecptTqiUY
P1snse1xQZlIYCzpfpa17pruDFV2y8gwWd6chbJmdSZr0emvnEVbiCq2c6wYCzRg
APjHh2fQzBxrD7+OnoEMWUkVoTI4ZF6tRKTFqb5Y+ETUd0lqHM381eo8kalHfigC
zBbXyLDRwjFG2zXcHS8IvjEM7xcEY+/+49EWnHs52FZv31JdHnfDJn+VAs1SObFZ
`pragma protect end_protected
