// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0
// ALTERA_TIMESTAMP:Thu Apr  4 08:27:56 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NYAa6Q/puWSvrbMmqfpcnR+65I1vN8sKNU4tzkNkr10A54hag07GbZyYFvXKX/Ft
pse4FSwDf9srqEBxVsJGjV/MEm+gG7tRHFfb73HNGwTxOwFEe4ZnPfsjDYYC6pDZ
bM91bmJOGRpt82u+X4xxX+vFuy/o0qJ66ZgVF7lSvGU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30176)
Z6YRgBejRw2N90/DE9ppgYPPa+8e0bWeb72fWF9LwolEYvK0zo3qa5lnL0wWW8Mj
ziwt/o390s+bMZKbNv8JQFxkzWwRKC5rjnTJh6rNXyGNf3Cti0KOAsirwWCgQYYw
pMn/aIXh+eeMsAchO1swwpUhtl8YMjy+JEjDR0677pFl6TurUn09uDyFRIn8JpTV
wy3ondBtTLoc4N3YG9/4ZYQGPZyGyhXm3wchtW4119WOQA7sBZr9v/kEHYAFjVSI
Gjs/K2OhYUL0jDh/fYfvfFiR+qOqM2t/J5RRpBmgg8pQ8rjWcyk90+AEwhZu/pif
gBoU3j+ii2R0Xih0KVfFBvvnLJSjCXN54RrCz6yznyVApW0t6Gyq0TNA9y1LKTsP
Cv9EfLBPWjCl/RKrsCHupLzYk8ieSmEoIbprN5/WLO4NfJqdojf941rK0LY6MX3a
fr21qFjqWqp+V1sO5UpO50xCRX1j2/GilJrK9E1XhbNOm6lsohCT//oz60DHAofz
hJuOJK+AsD3osRBHo5DloqUZq1737b2+JRAlP344DqHCtOwYD6CP1rPkT5cgNngk
camfPAlqjKcWsFr+pymbD9tjYiFUFlNj6w7+JGN8qlcp7j/UR+eYW973GfxN8Ro0
i0/VjeJmuJX8QAsWbX9i3Go1zdQmCGuoeJKJgO1JnHmL/tS9JTOqq152BnKvjCu2
wxjNJyEq5GZE1Sxw8xxOJ7tVnllB+7kBCvQGe44xTngMy3BVdOISoJq4k7XHFpAr
R8D4v1Qm+B1KX/RWdGDVS88bdu7PQnP35EtasrpqEKubjjqFNNTSsq70SL2YZNCh
reN83+hP8Qp0+dTarQb3wWPVAAnM705+vMm529bUAPSx7L6baqlbSMc+dREEpte4
5hok6u5a3/3bm12qQb88XQBitE4GD85VoxthiCmc3oGOD8rBdEwd7kP6fKehocro
seK13hPEW8qI2ffly5c74fSAfgX/jSeAbWB/uaYMNhnQxdx8GfXaOC1jC4I62lg8
yNroWq6jO7vlD1O5++um6Ih70qCzZC0PbKQmJt7z4SC360aZxDhkCj0Ur4YUS2W6
yddoM1F8uyRa23Hk818cM81ll51VcjcfPnVZXW2xyk5eBpoGHS0+2Byh2pP3Yvq+
kBBoLi6PODo+y64SZKLVo9GztnmXa7dHUQ7ewaynCo9wSXwFcf0xuGnLmQkjp3U4
g3K99Md5FgNyWQ2qpfG3gITUpce7Y3Pg5vLI+6NbZryHGn9sAZ5BadkhzytmfDc/
iBbR9zHzSggJY6OS9OJsre18FYNLClZ1anzttKYgs1bxuj/yMDzw4H41NtWa/3be
7FsYH5bF4gQqMR/0ZSGEY+fJziUHqKhmGVCvJ7O7JPtzFQDkGrAO9zSORrVpK+Vl
y7lRCM+jkAHnb8Awi00x2cTO3kjLCLRD4eLm7MijUNh170F9U85hWq2/Ejj7t4i5
fyT7UGZF1NikIKrZT0JA7LZMi+pjrCQxdGWjht2xfk936fCFkLC1waE2NKpYR+cK
b9TaUM8pt/DbDXpSgtyX+NjGLboEyg9AnSXMQBZDR83rlp6ggpt7EssEKbr8+mXD
wTJc9vqn3+C3g9mVEm5kmPvtVx9o3DqcSmT+dXKHmF1lwwnp5VwTQv9wKOoE/0MV
F8LSO3DVfIy212d5l2eUcUi9EClO9XpM4IHI7V6g5jdvSKqErPEcW7IstB0L18xa
4q7Ew3CQTUAlTxbaCpKlw+XzgSc8BKz1gohR3CtXSKncmEJ6WPTPTkK+TJhpZhJO
NW2I8kH3YPgdYb6zXKdtVo1TZvnhZVK1UoEXqCqX3ydpVMo7BbcmCMnuQssR6dVl
OxThsUHFZbak6yZLymiiiVELD9ygqrrBcLw679L0jnQw98Wz6mtJsIB7VwT69pXN
HIqodtbWljVOkg7jT9i9TpKBeyUo9prRej5JcA//wKvkuqMs5SaSjH6aNWBgvKLm
8OCm8tfpE032/xxbC13ls+r1P4CpUHYA+Te6YHhPuseg4vFAThWTnzRkzEKuBqid
TLU1q1JF7FIs/5fJUSbgogegRX4F1bq+OFPBoe4UiYYL3MpXau7vdeayjVjsVFa+
96Bovb8NHXzdauwaw/UXgZbVGqDGR21lej8Ge0vFTFTk3U3DWeOV85eprxtL6UDV
825PXUTGOElxk2Va1B78NkCkJNZv2GPjjBaaXdwtcrf44bLZUkCS0M63oWC8HVT6
RPzWN9OZntp4dHxpK2MDi4gmiuouyQ+HZuYtXHqmL2+V7KZUIE2PsOnR40giVfDg
pYji6Cl+HdMlUCrli83EUdgXdSMGdMcXco3/thg0Yk+njLzhJMBxnoqC/jYfAj74
SRkaV76tCaEsrrB1Po7JfgW14x7YuJZQpPfQIaKE9R4PAVr/Ns+Nxjdt8reSMZ60
aXgFggPmbPGy9BofCi/zCEhlBcp3pvtj0NmWU8T2E6fGt6odtl6f3qFFSIcGn8lH
4iBOCg8GohUjtxFMUv2W5Hg43GR7ibyoRui4AaGqqceoqMuUV9ztBisIwdcj3tri
4SgRQdcYjesRCzo09k0tP+AcYiGOJS3uADw2aeAAdW9JxONY9DbiMXFE8EPnzdAN
r0ItjLBrWRqsjYH0ZSDg83qlhKDApryN4owbj2eTqDv2in6jBsae6QVjL/CtPsnc
TFyMHothsYQGK1xh3hoWY05VXEmUzUwiKDbCcFgz1d0jD7qeANg4PxMlPdFf1QpE
Otxb9PtUcw68MCO5ighZ1CbRHTbKctMAnf6KbChriaIODm9YDbWTRI+JdxgAhWeX
bXK54efIt7T+HDaXSRtX2GESajqSXU77FcXcWFEG4jUuHV/eE6Zw+G1rb1PNrmM5
TIT1KVyTpH8PsIkL4rdfgYLEV6dN6ovPriBq+nmz48u/XFFh8hOy2EFazN9Wu3UZ
Tu416yz7POZtfRVzaLTOMwRtzJLfhrNgN68o1NqT+qY0sEyJwFc/d94jhiZwU/Hk
DXNCeD9QnM/Pu8rkXkpEz+4WysEnBMDlaU3dApqnszp4rMtXYjxnFMLcFPfByRtX
rBJT04BJtRrhwb0Qg6subsByKumacHu3857hJ1LhNXIFnZUeCr6vbz/LJjv7yD1I
Q53T1H4RwMUU+6rFFVkcRbsqG+zxpU5oDhIpA86sBSK1vHmsbSNzWieUJQNkmrhU
V4APUBwHMZ40KkxyxegImPECIaRWxBqGXGns7lgk1AlTrDx9CgJvuwY2YdpudFsV
ttlNsgN/3X0H11+iQacBmpKAvc0k2hfe5c+HCzJJEATDe1zaehcBX3G5JmU4FV+W
xsky1Rd3FWBhA8fnHFe/oeOfvdMoT35UlneMbwpQqyIOuLl07OS1HvW24ap2VGIx
tHA4t4G3cSoqC9BorgRKAVSisCnUEjN5ccZSovDZv5f1XdSe2MBKSsKMhbBX/5ba
7syGzUeiprpneE3BvZMdxBp6V1KbbWLRtHfgDm6eb44/w0vGXki2/ZjS5MFP6Dan
1SHPJC2ysIkbGZgeC3L1bbhEaMV5cXSj7nvklW/lYk5FOsIgYGqVgh69oFFmZ4MJ
SdhJWEKCleE0bbSUOFcVdMhtXwd4XZQGiTRiUtIcJu5/F1Mt8XM+zsrv4f433C2w
zyKC8XLlOT+RDIYZBOQsPGVXtvCKjrCLr3+GCzeg3lRmYQ43qGlfRqcutRfB6enB
aRcEUAUOtkdsAUjbWA/gDpi+2jEjiQ33p6+SmYWrGYBLCg0XrFJI7CYHZRx8b8sx
ovBk2pM8zD+Kh4Wg6gAxINkJnDu/6+8R6utynA1O7kPk/FTqQsAUTwBkTeLsfHVJ
LuzImyALp9N/8wN9aYhT6AqBjrlbpIQMFMKwKoRwaRvezv+4BoOQkNNh0fCHlhfq
OrXOJlcXxbyBY69TsBuK9Iv+0WVdF18gUzL64weIR71pvGARZb6ydAAeaqveRVXI
1Z0P+/E2hXS2xjDIq1ohrfPExuyuGdeA0GmmDOe4emn9FAnacg6ul2MmOyUIHK8f
v9TqEAjQEI4WxpzDprosGGLG6gWq/pc004nem4rNvJXHFUTxx7yn16TJxNplqZTF
ocP9V47hhywDM+31zSaOGz6dniMCIoWh8V7ScXhfVTeNkyBcrCl9EiPzRRCHiyz3
8Ff16NDA8YPuUnVJOZIobvCN5fcKFgU2TvjmE8eT6mHNOtVZxu+PKHerCL4tKBMI
e+9QM0Nt6utunIolQ2dcr9mc2Zb7tH34ZmRyDVu++z1yiAV5GrxVAulW/Aoe4GFv
8fl93VRHbpCyktxuWtrSka2GR3ghSzN9yf3iLOwRXjS1DZbZRGtu/3uN/OEpVJ45
99UL27ohn2uAsdmu9rygPj/uso+ywpAu5zv2QLBjgu72J5P1y54rA0j9E7xxJCrv
x8lb6sjaKtuMPdmYkG+IXJ7l6nxDW1xEkS4u9FwOoAcgxbd4N6zOBfM3XhWoRfd5
xefOa1K5lLiELodJ5AFHXkG7Qi4e+OiMi5DqVG50ygdlm3iaLIePhXy7gsgRttdk
e67eTWCFBiWsWgj2zoTy/TwW4cjL4H+8ahMN1CglldAeVFT4FwtpdsQNxtvDgZQA
0/RwPMg4PLK2IU1sY6Cb+fkcf9EXpk02J/uMank5vvENv0zGx8OlScozxF24UGoV
DyWIKXgHiipZT6gvG4C3OCeoQUdE5pi8D6Gs9sP6xOl+B1Nk0MuJV1ED2J76SUrU
Lzrue8T97VmkGbdqUUn+/WfE5Zk1pNO6mMB1N25TZGbhehhQiaubMUqJ/WNzFYoM
oa5rLDeVkmXDWURemL6MxooLCuRpGHOmxUBD8goshKBbO+8q1AMNyN0ND7NqKs64
e6gSuFBqKoqks/3q2oC4GuUt1AAXqG/31GqX7LhuuJ5oai5Zbe/Bg8wP2vS86mr+
L+RJp0cBm88BN/ApZOud9unWTzZzQBjfDfV14tUd2pVJ/oiqnaGQPh1O2ucitriO
t/vq1hkSZWYgilrtEw9eUzPWtbN+E8ZHmf5xrDD4UQQY8TtYQwNE054FeIJHgPpU
orn5dUH60iRxupGUHQfxAM8a9dRe7ThYU4DkxqW9VDkFxakfS+qCM+Al1HZpaVwA
9ZHCdRjQUl0Q0KhebXjMfpbvi5MTpKjZmHRhjlURvittfo59Na6EQS766zgvfuPv
amoZGTYUVfOKoKcoJqyopBWUCRDqVhShSj06GZ+2+av6lKOXThRC1ezTk6h8Nn5G
S9NsrpUJUWQtWBKP9YvdAeF87+7VjAvPvMsN+9QbVFKn8KFvnl1IiOtIJFAwBHr9
OWkKnd5higY/Iuo/jQOsPGdxKig19RPtQIE2ZpxoPKPrCKMPoDJJGMcGwJ1+u7k0
Kbw6NnZhj6GJPndPU+Z8gv+um6s3iX2DO26CH6WsoNnmwXyMtOtQ9iVFC54m+3bz
7pIYK8sJXY6EvUDONreu9RgPlfXn2D0APreegcXJtmhxzN8ifXrgBfsIg317+PW4
E+O6XCq0SBE9k9dOTX2ZJ3zycnGzcM9l0KnAd7rgJmO0V3arhw3Lx/VaWEneWCwm
WX8qQajSvLmSNNhlpItMCtWw916QrCPjR8pLl6x6Ssw+uqDDEZEjwvvf/n9gDlkj
lMILoFYSz9v/6toZuQ8bfxFrVEoTxWajNIlio88JY2VJh64QD8ma6I+ycN1v7bJZ
b0ASqFE8dRSNgguRhKGY1NkuGDdmYsrc4/ymaiG4e7LW5hMdUY3YSrfsB2q/9/ry
tQFwJWBajduXrJSWsXRxuVUZUw2pcaB6iLKVTZAKpx1SWH3+160z30A5Pz4XRtTD
eyRQ/swIjs7fn6WZR63xdwA8syxiDP1MuOuSD1zMtbR3dMx6nJb64L32t0unp4ty
416DTavrqPIFKZZMED9Cmq9tXPo3TnQ7a8Qga1bBe/sqB0oc90MV+IHPGQvCeM5L
1adc0eFU3UX6f+kV0nPEIrqzq4v0Om6ET7FLDUjg3T2gOvEtWwwwml3c9akt222R
iT1scbP5kk3aKlL7WIw5r78zipo1xNqJK4b+E1fp5ZLisDQw2wUmKyLUKtz8ryWj
tFPhHT6Abc9tbXWHeYBITjB2TdYDhngIrv3EqNHWerYWm2sxcflWZ5yVVBbvb04c
pUk7FiX22HeOQZtKT3derrk10vGb++TJok5qvyn1kkM5Ly6hgGo+kZK4cPTuLvVl
IWOu+eL9nuR4bMgACExlJ4ziIF7ZI9a1EjKEyIRo9ZA1e9fxo6r03+fW3kf4vN0C
mciKI3D52l8M7+ainTdnKkBIPbSa7i4QeVA4NgJqxxka3ONXP3p00K8ano61TrR5
dXqSrgEWdedmtdjzxIPT0k+ZYn/imF8noFV3yeQXV0p+tUnFFUZ7bfgGd0PUwQ4K
ecHyGpbl3PzZ/IEyu4AkFxVnKymBdtwqtOjR54ax6c/bIZwyQf0X6nDZ8Ga7fJX6
7RY47NBWzJHwGmF3/hFj5wIGr+/Mr8QL+Z8Ku3iUIlaE7lq3oOim5NnLEycMc5lD
9g8ay2C27yJPg7Jr5HudIpl4+DZPutJ7jIrHmfJymH/pdB/lpqcz8RRVak0gaLgc
RKiVoqY28GnxTiARX6G72nkwnBYxBVxAkx1awj4r8elthWomKFGkQy6FBgGwlrlg
KejirMQEN73YxiPIRFnV7U7+aP0DDCX+RM/m3PrPuXJKKzKEhC1SSnoqbpoa9Ynx
Utu8lv0WRchHGltm23Fui2mSyhPSsxAVWHta+3CF6ZoV2DtvRAIsZ7jHNDfCIfNQ
lum5bbO1BCGRuYZmMA+25SrjazfeLo3oLwdiwj1MH4cYv51eKA4fYSWXinU7kKbU
3p964pcuKAQFdVMw7nN7HC1uSy4G6NifN9hkDHeQIq/S5bVvgtM+jINxtz4dhZ7S
0chAPI7iry/lF3TDcn2pQepJRz1H78Kv2x1NiMvRJpOLZCgMHmM0EVRvdkVbUe88
e32TnvajB8QdzLVi8284ZzE4j/kuNsVTPdLe5adAaDcrFc6/WeLZPp7Vr+m2RQAG
QoPe5XAZJGKgFVuv8DAu3kdHrCXugaKyqlF4B5N9x8PbrRV2FToZYVSGOhIGO6RF
sz6p+LNISCdjOZkN71staaUDg9Qm2Q6L9kUt2uuZQjxv7scC0iXcwDnYuhvSiy3v
hBOmB1JupTtW5LIMiEwpWxN64WRnvemSRSxhCoizPwzvQapB8MuV3HpllvxDLNWa
t0xE/oGqZsUGRP28wUREBRzpGk+RP6s2afAu9qVMu5wYYFGjV7oTXTCCmJ3iFYaC
W8Slky60up/IFEgQo7YLb07nZF+4ObKG7olB4/5+rCoYW8sfvX4BgUVMddKfQUFt
WAU8x4n0C4kdqxyQiTDBRvnwgzycrvVQTTXgtJ1eEQthucD+Q+zeinsZDKJ6Yx06
iU6nkjiSLqcZeG0JXa0CnGT00OGQy4DHTHZ1Gri5kn2YIef9ycih+hWmdo22qgDk
Os/rQVwUgCBLJdaO1XF5nsgPt8H2BjOV3onXStAE964Abkgdv5bvKRmoPocw3geJ
RvBEO0Cw3UtoTYzmOzWnBnBC2Wlls1kUZz5SG3xhM37XoSzhvBaOIbIwhEj1eYz0
H6JbkmuSi8FigXi/47hxOdpXSI8GUnmWvbm9Nqi+mXGCsHmHZMorqSgJRrsQL/Ta
WV/3rrDZd5os09r23dAijZlYWRAzTHKS3lgwzHxPMwBWbcF4X8wLR30xzaMq2vUL
hFjyd8xoQlAJNH3FRfMN5YkHkSnUTZhKJWZ+o9lQzSxxVTUqbC77us9GD5G75IEu
M3ygNCKcdT154rUv2swc6S420pGAbhoJu6Eu0kqq/RNv5Lg3GVSXApse/HkC0KK2
7L6nakbN6vObEeyCeo7uXVRfGuSh7+oijK0lqzigQuFBawUdxluJwdLgB4suE2QQ
xkDjcsJhPjumWP48R9+4fjrZmkNwKgP3ecEIwqpnZHn6zB0CMIdL3jvj6w4qw3fF
4uuSds1DU4LeUWK70bMF3cVTyCbECA2X3IhO/XHpXgdti28abMwTBx1SNXvlFXjH
JmMB6hAsUyIm2fwtcycmFjMFf9ZskkpA61rM4Qos0+dM8owNzUAejIFfE2jLTNoQ
lk7GZzeQCzWUkBSY2149DOz1SeuHZuibJ37rpogAUVgP60NyjkJUYnz4o3afgGQp
3rtNnS+DIYqVc+Hp9qAreLtL4Fa6ZwQuTyuIyPffQDJvmdaPdMJ+g28aBXPrWndO
NG3r0ZhVdiNZnFeWLqVLlh9Gyx017PY6/fzwoIHQIjThftfpZ+bcbAPJEPC5bfw9
aKpn2WPlRjw2SbyexmCQB3dzUkuC6OWBJ+zAWg03rqiiZwVA4Fu2y653gNtp4Qud
yl93s419F/NNL4KMnzIbExWiOgkciwcLLZCm/KBct/vQs45YQ0hwVNrZgmvPUjpD
kdYvCWtV4R/SdEo25avndO3h5421iun4wMJQCev3d3aWC5TayLkuRfpdT/1pNEt3
qE7cynliGQIRRTPe++kQEYvWSuXkdiNL7kbEgIuOq/NZXXdwAoXPn4ThZ8/92d6B
PPkgenrte5djdTn/EljHJi94Md97ykC7cGQ75wshXcFsO7ZsUFpGm+ZhiQSCT/P4
qjsZs6nQaQ8b0CRDhXSOVn0arF/xqhDPxmMXgl6h304GxK5o5gsxYiEJ/vESReyT
eOOAEYFUsnqAIxOmBKNH9mqLa8b1b8hb6NbyrCL53x87yIaX+F2ybJyfYIAPJpOz
ggiYUj7K26YCESGMppIJ5WOorMnX6TTOw4gQv1Z6W42r/nMMbOcyjzkTv9R8EHuW
e3uyMgpfE8FeBkiNPG5bOOFSZ7TG8ohRdnFNu63vMQVeUsH+TYLf6f0etdOdQXzK
UAfoPs+86OrR0ZoCg7rnejDdFhktSFnhJzKQwLN8i42FyxcvCb3Fsb9fu3MfmVdF
VDqTH+jhiRspJDOoJKC54lls0Z46x7uHzmnVlcdaeNoVfN8N3E2XpxyHmCwwTV4t
cadngZD6LREXdV4zkmVZ8NRDbO939sTCcabKK6pDf7njDG3gTj5YIgpRDxh+KFK9
428YKR8NuXiX4PZmDP9AV8QA7RzgTv2Gg4nfj/AxekeB/zRuwKZLFbl9DnAUNzqP
GTlU30Vx9pbShNROIMluEYZ/lYJIK8rYOhiHnLhX/eL0Z6SMGVv9MpzE6eBuN72D
86D4BSMqSIlUOCsDm4x+KPWuas9A1N/t5RONyVrVzOoCJc/0+hxyHS/axQJgj5TB
YIb7r7mWKvn2I/XlBYv02wfT/Ko+VXUN1LPigtXuWvqAAAkmF7h0JlS+TgLBtHgu
C6TfkICi16FNtooNEYDQ0dfJj3R8AUp06SpkGvoiUiihR8bGJYl2tCE7tMTPeVsn
udJQrvYXA3xtmXhg8fjSB+aFgiqdms8WkpPqp/HpXb4Jk/haoSqxKAoAch+UKLI2
H2Na4Namo3P9zxa3TSYDw34Rxc4nnU3n5oyx86a6oZG8umAxEtuYMdIFO/i4k3b3
DcsSOtcCHHLgtkSaL3tIbYKOp5OHRqpDDAMcoxRn/84zBiGwhu4Gcs9lWwkhlicX
e+NdUz8f9w+bx8VNUhhM3fJLCgmRdkuM3HNJQGfCarlMjNDPGUB9bQVoZjn6WEIm
IzL2ydCvVJWUfENguPWG2HlC1BT5QD7fCyU+pIuuEIBQKPEghmkgmqdGQ7iaEDpV
M0PV1sKwIo2I5a8GotL+WAhiO4L05Ola3rqDmWCTktVNWm2tvHdHZ99sCxBl7rxT
ulws2WnJLAKREY1Y8sPWS3QoV2ASebO2ojszYZcy85ekxrKiDE+A8goy7qXYbFqq
wpIm3RUjVVurMtnvvV/VZhcDjYgMyiDepkVUfuHETlke7kHlGN1N1TLliWr+VhUi
woX6/9jLZzJVmCM7xfgY9xxyJk4Qlula08u9BwjZPj41z+tx/Hhi7/ezVMcW0rAf
bE/s0u25bX9qcICteV7vLmisbR+tj+SMyk4TLAi5O7lquunF0hz6YeYhyY7BXrvI
zN5rq3PMi19qUrecVlnimTpklHVPA35QHsMiCxzU7tmL/Dqq89IO+7wuNmuD+3fT
zXObEnWGYsQ4biXuGPDeYdInEvH6eiShdFqg/kBGmhCdfNfdayYB6zhDPAcRossV
2ZDMJmFZhdQCgZ2jObWP6AYzhbujR31ulUue3GStiFyJQDZxKUeoS9+dklNLioqo
EMNN8L2ndIHEf2BEr9OhwoMFw7LVZWX9X2nrpdkS16HjIVkfH15Bc4nsRZg6J7nk
PuLb/3a3RNihkTsHvWcqssFEmBfGZLZTLFtIR/UNV9E9tBBab9ekGtTvDMZitC3c
qZRcEF4TIdvrLF3Bd8w/LYDt5Wqr5xXydgnq3vZ32ZBGZ2DUmyeLvpUmxAJZB1OB
JB4ejPhbp7PKCCdNc/0rAr+LwFmHrMoqBXbAGmSTC3f6uHIqzjCB/PMljHgsoE+M
IZFl8vIMSebp9FoBjC1sivZQ2D+kPOdXkas/WAdwwTFsREkCcy8D5p9yiFwdLkyn
5V2vOWLyk3TAWI904d9Ywob1ZWLfoY3/K3DkmqC90qPlw6YssWzD7iCrTifOODft
oivGKeKPwJMmNWTqVc94APxj5L5p5tfKDZawo+heo//xPWubH1XzN0Tu9P/FFCGE
Cee7x8ImFlkmpTbMq3r9NHSKA9wcGntZkkCWB95/33QOhn2sehkDj6+YCjs1ZrhB
nw2hIPAEzEjP7hC6iB+2TnoCqrUsqvQJiw39z65ucZs4Umfa2GZWHBUcsv5PRMF3
qRYaTKCziJzhVDYFIr7jaDyyk035JaSmCk8Jv2undjofm6/2V7DTv3k5mdE3bJv1
WQB95Z9U63MSESABB88pBgtdDpHCBXWjqkmPna1lGT4oWpQseLtHz2gZF0i6APTB
GuR87iORcnBKzHMlDJZi/yhKDYBLV6tfhrlwQ1ghfc4emNRWMmyLw46IHTJo9iaH
hUFkgi+1i58kbNp7yg7H8PUGVS9N5QLTiuesqSEe3G2S/LdSbSXCbhWMyGZZxmhg
al7MoxZ3nZU/X+yn2MOFvWMORkvtlaQ1x0LDH2w5LJlvHt2CGdjk85Yl6n5E0GdN
EYskORUGAVcCbAjtMZ3hd2GxgHRX/VcL9jgyUJHGzTf2lKQiSBtkFAdRN+FRHsTn
vm2e4RmlCIY8PlKiNGJsQB0slF/5II/tCwx7V6krkDG8f57Vo2ScvKgs9k0OkYTE
9kclaqzMKRIdLaVTlvFD5L/FuSYbzCKSBkj9xmBbBi+nUUM9hy4IWBTw3bG/aJ4o
34sTe1pLUh6R14BNQJaZuWm91QcN8tbRwEOHwn21RXTQwYBs6pslDWI+qOGoQLWe
pA+bW/xm1p2KEUd6G9uWAoshl0MnxVBSsk0oLx5AJCkYCG40pGfcXpU0kHryh6aQ
jpmZjIFdfbDV1kgDUF7G05PsfPTB7rMBRWib/B8a5+LLOEKWCe/BTglCh1mfukSn
4uVw2YL4gpbRT60VzVsFJISc4PUdF9sSK42vmKJiShrw4XoyDwLGrtFAo45uM7Gk
N4Q3xKPwIX6EDmzbYG+CILvkTCZ1JEsnRzrM09IYw2+xkUfyEib1O30UC2MfdviZ
RU6FPOkuuaZuFPE87Cyutgtdk/ugKmRKUbaOExQVFeDTYUSftuj0Vv9jPieNuRnd
VgDB34TOhxZOiPUxexa9Qo3uptkwyKFJUdJDM9uykP8RVIY5D0GbLVH9vfLdPK9b
P1NJ0lXBOIm23opvDuGwqQ1OQKnFBwHhLTr5Ac8H7i6rlKnpdk/ArzAm5oO23wm1
sKEKELXaDJ+UaLADrYFmxgCZSXgJfcW8lV6h8SmAZg5Loin/1ARCAKY7/dLGdIRz
4BfVYLX3xNUo8hwzRT/7pt5rOMGidYQgl+M8C7kYzARSWxIaBBC9ccVyrR46YQ4t
6zxwiYzhmtULXqwxRQYJFFJerMQP84Z9oa/klC4QxYyoZsN749siKFxYuybYMhjr
LpFjsKyPVrLVUpxPZcl+5hFtWApYOJpLbLod/nOJT5IcX5xDZl9XifyCtzG5Gg/z
9Vl6/qmhJB0KROzUobD+ELNnzxj/gWjPlbT5xEbvWKUfbcJIWteD0+RE6yPaqDbz
DURy8Ch168lhCrUDUXrML/MaijgZg4IP8TCQvCVlg8dgfuuuUSzjpm0cdn70l6Mj
Z8+qCRvQr+hYy3w10H8s4M2rZvkhrrxFlJktPCKgYqTjzV+rJP6ij/jQW8I1eWlu
3DFxHjC8ce7Mi/y4zpZMhp37l6gNTc7GY6A8NY0RNNKbFfxyxe8sojv8mSaxpVg6
edY89vFi1YpYJh9FvxrO8W6COTLyudkASAQTK4A9XsEz2kbTB8ypRbIlruN9jK6c
GgCubpeljE1rr8z4Y6380d56XOST9ePiAPMIW6jDQyPQD6O+i69hBUxtoHu51LuA
1OYHz6aFxlVVKO5x1PJn8FZXcQYv0QGIGCpwUpYdW8Iv3ux651Zu9raNnzUh8e2I
KL/XKOnxFWg3i9JnC2UJrb3GrGPTsgGGRYIrrKJlpQ7uj0sBiWyDuTnIStdlLTo7
RFol2X8f8iSGKZ8jPbEo+ZF7pLG59Ha6jIHRO5AmwrxAmnHCn20yf5btYgXqlo1K
7Ly4AfnF0VqjRkgR1ymp3qDZ6ZgGcg2jDkpdjXQ4FGAlNGmmas/+svm/gv5NDdu+
buWvGCzRp2GTsEI01rEbWW+k6/VMWFI3xvz1OaZw8j6+NGoejAYRmt55qOOFkgWq
aUhwyjmTJr20CYdAT46RJ44ySvcVKSbFVwZDmHkvjGPK/ZDMWpklp2+ng03IHYSO
KTrALmxSmdr4GbUOxvleRiHWwC41WNfCgCwrysfNoDwNqnqJ41r8gXD8SS0ddvBn
fcEWNkN5y1ZOYOBVC17K+Xc/imSRKtdQvtn911cf1xLEnlyztM96xaom39E25KVt
efbaE1Xko0/UUMwYMoJoUROTCQboZayXiSWkMp3vYZIRAB9niI8cGe6z/EUET5AX
usjJ2EdzvgvElxEI4LNTyhcroVpYThLnpXfvYZUaBjnKWHwk0D+m+SBOVNDFRgo/
7Dwnh9o/XeDk5OgzUivfFZQ9dV1G54EPX7eugAfzs29HfD38+a1cFXh1bjNH2ypB
8+l7f0fyOSP/dQzoKOhkygGyFB6om1hJ95L7vC3AuEx39C9PJZ/D4MBkXeStD3id
pLHhuCs6lOBWamTcnj9kE8XOSM08aAUbQi3tJy2xHESCc1enCzKCjp2SlWNZpvFZ
t8bBEeR1tlVnurKh5BjmdDyGcB0on0DUyjnsR0bJTLhKNSaZxFAy0p2aWvobz3n2
9qfKe1sRLQ5UqYw0xkMpYUqBSuifULO32+DI3NaBFADpusgRkmonjOqNNJgCPO0C
L9WURGBzyzh9yWQX2Z2OsxofiQ7t51N9WSdhmPQK/ERpXOLYJ/ooOFMv66jOPVeX
Jj+Zk6Ff2Ny1l8DOIvxlWaKnfdP2/y128fmixaXuyocLdCS2WS72vnYXZs/rAzsB
5+hJdp7Wn9QyuI9JXsvg0Ywq36oj7K6U4iF+NBgmMKq1mOOLdjHScTFQLyN7fZ+A
LxISVuAeqdA8dN1VTa2P4TX1BpKTRfbpGwLQhob4jBU1Mnh/3uqpWdc9cKCYA/+u
1oDnZ+3iDIwUOc+EDaCke22ieFJ9vewkMf1q7HJPRMzwBzN6kc4Fu9mRhsruzqwl
xW1jFVC2vFSQz35wgCh67py/0nEc1246WOjATeipncQ21mAmu9naqsduEBmrZcQ6
MvI+xrHuF1T1NWO/nVAJuEmeIMyldxuIbfU9CErzuV7hsz1O9Ah4q1M/wngmSSK/
ZTSKiQqLjefWyPmO0jeFtyo6SBQHjQIBOFI3aXkVK5FHojkIH2lzFC4n095muqF2
bHIdE56vMXixZP5v3Z6gb5p9Rx8KPBZ9o/dkix7hanAy02Kjh8CIle5qewbfnzF/
EMB8Sv9V3pPWZAIMJ1Mhdnqolv0K/cgCt3hAR8jVoGL4Zig+n4HODcC4mkPeb7HY
l37equIWQT2ZhZDnxHuuiXCP0dOfkDmOr3ogP5bjidSHv8fDtzl93HblTCe6j8Xh
1FF91IH0Y5Zke4Kl6/nbdVSjKKEd2rx9YNClF3jhQvWEvOOL0rbfV+NzlzEAwoyk
c169dhE0B2gW95Ik0lIxStKpM7J1icCJ4ZG6RDpcXfOdt0oBmfJ9pV9FarJo17ty
++d8vF3vfhNQiNVQPRE2jSMGzGoGAE0/MjFspwmCEYyBC6mcWUWwwi4JZ0fW2+p8
KGVV+otWgste6YTW7V0+ahaPlwwA6FVdzoaZAPIujKTtUHdsHSbwAHBXlyxf/GJY
+1rS2qWPE9gNdteCpzmVJhO0jkh7LOysJaaaOQQzGaGxp0JkRILLqoohyyGorpVO
JCLf0vby538Igq1O/LyJ0pcfslDjLD93BD9zOlrXhbzb95yOW7FsNN0JKnIXyc9b
qOu7hs/jjgvDiHvcXS8lf0HkLek1xMDAytQMN6vfBVGhjzIG3Hx/JQxORQKY/Fgf
d492RrA5Vjbli5lPdL0L78hgm8Rcn6WHvZiet8wPFQg94L1t4Q9KijEYNxV2d/g+
OiRnCalCcWvKmJZ6EbSzHb0H26tyyYZ0MEqJEjTlw/yOD0h0M2V+2DeGjWkcVB6L
faR0o3a/sQGD1gVYUbY8FFbGPCGb4cu3QRJttwESVKMcwBv8syav6PD653RwHBNl
HRWA8Ewzx+b2+FuqeEhUY3a9qzuxldT2w3m6kJ+ho+LWVwdV+ADLSXcjlMFwgTIn
H8Ua+YvjH7XKuFaJK/B4TYZ3bHkpaHosJfIzOlu/rhNxkPUkbPTdzpgtCknbHsv0
1w+QUsp0QQHFaqYUqHjDKJRdn+LFahA+Qkdvqutc21H9b7FQA4DwEc2JpSNpho8l
UNTjU+5n4warGWBu8iVTR7dcQN4imN7ReWf2O8RqlM5r0IRsV5tRaHzURjMIpsqW
kJ1OGn/MJ4twR1bKjgiPgL4rmsleMqH04U0X+PSUj5et76KgfVnMFVJ026Ehx6lU
Z25nqCHbJVbSiXyPCo9v9jwzvkz7l9fKAdpFKRkYw8HrtRs60p7v5Y3sgXmUc4n7
4yEfYP5CBsmx4ZXVRmCCbHdYmM5InzaQ7yhBDNmY3ye0LatRQwfjrkNejty2i2A3
fvGODOfb2XNsLOhj2dnQ2wAwIxYAT6MUS1LuFRH7njEXLEJNt7wHdIv1smTvqYk4
2fRebktvR0K84mRolfbmf09fC4dL62iuNyYcP4L5ShS9nEgL4Fje8INY94B+Wm8M
P1Zp0qNT19U21iKJDKsnLccnhzYTZbPu83kT0e6gY8KCUJqlfWgOCapvat71inIV
eVlKFO/uZejjG/+KYycRAg0Ox5kQAspT9X50mPJkjub8lQ05FLZzNC2KmuB8wtjl
NnSzpqQaURxAfJQ16pb/eqr3HcX6MGqQuem9EIS25Kj+VGEewYszMZENUNVhIOxO
ffCK9NOKAoIJxJSMH+qFW2JlM/GJ2m5lNPueWb8RGA/V9Xe6ZL0ILxjUmlGXhNZw
HHqBCOcBszgJBI8zJBKqoUk08tm6UD5I+sai90gF+q61yUpGlrfVqhKW/bO5p3U/
uux2vC4W+h05gYz8Fi4awKXPQg/rz0kMHzdX1IlQwuvWjnT6363bej7v2SuPLXB1
Bv3qxnE3uHa/YogX3dHqMNvAZ+aL1PlVMwB1j1TdL1ARViD1O9OAQMXHpaM/njET
vRc46QEFqzfQ4DcQq23d8ZuaF3cVkQhMa7+JczQmITlrRZiZy7LKRtZUIhGr++FY
Qelw3Uo0Vc88lZzQukXeHEHIcGVl8A9EFi/w9x7n4bGIkwPgvfRR54l2Rv9lDb0J
xga0YgsJwbo0tk4PqWEoEfbvpOk7l4RPOvvpTfRWMlIaTVSVNLg1evLVMEskJuRu
B+QIceKOzRUSYjwf+vXnt8eOy23gAndnm86ceg6V40dv8jXhSrA4ClqwpDx0bm15
eP3+bxPK99DF6LSlIplq9oQujnjPa6LO4O6uXT6MZ4aW8W/nP9X6KoqT+l0k+Tot
yFN4hy5neLPTfUH/54Fn2Ob9sWJfAZZ9WzOZkINcLJEpLkiqEOW87Z30AsyW6zUd
qWN2QuurcgFl1kI/Zqe38bK1MlApF5uDNdnIUzHQCWyb4+GW6QHCfkqkFfVkRu+b
lEKzZpH9N0oN3HITHSYUa02pkZCJJiNNAoSmGo4V1cIXfpxNYwpCw3D5eDdmBqhm
/o4LlaPk1O92Eb339tKqedHHE1GY1K1uVxaM5JonpvxndK+WShQ2uPc0fmgc0ad2
mCGwF0/qFZhD581PpS8uIxF5GpA6F1VpQbQ/lJ5iJ2Rpce14EKUfGY2vtuO324ZW
3BSzo6EsVHFMSqrDKD9PSMkeHvaV1tZdDz6SRfFRmQeJaSrYgmzvWVOdlpbrR8LO
Mp1QjVvuzsHqHV1n63ZaPWVO5rqvHgT1VbkYjYyod7xipVl1/gAFQ+gcfNG309Fs
v5bzKhg67prVa/oK1ZSn3ZhhfPyl+oVN5ro1/J4kwHvlOeqj21qElLQ6HzBc6JgK
9VNo5zdL2QaaTEpAMdNmAk54vM5x30/nI3MT02UlRqCDG+Tk4czzv3VhCfGwnikc
a0JPS03jP/55Tb36q3qv7y7RKqrHYO1wltzNUNpZuOtn2+3ugC/vSkqGo69FiiuH
A3p8f0j85oaNS7sBlmiD5FDJjA6plyST6Dhqbbvg5iTHX2b+s6a0xmZaiPxGwzmg
NgRFsLITamgc2Y4gXdAp8fx08v8x7cG59kmLQwsIs/HZvVaTuZs+nQI7lKjk6BQi
bzN7Uu7GA4/sAgB94CjjqZNCRccdWHf4qfh5nYVHmIvBN58/zpbqHbNDLN92b2NR
07prWXejOpAaGuLMky4JVk/Yf6I9lJpL86apQsrIEYM7wgYYiHh1XNSEVz6YJPQP
zLOQ93yPAM7eHiJyB4SP10Ix+Nc8aYVOLhaNY7+IpWr4Fc1LeSDSrEwE6RQZzJoL
c6CvxD3IPXYSWst2iXOekjaHSa9KMXEHHWaYeSLYh89K15JuMYPn034V4xSnCsQ7
2WmgdvZGBJe6WgQ9xEVyENFBUyHlCp2HFso8KF2Zj6Gk2zLyjTylT5LLP9MFwnpF
9HK8igLJdF7vAaGTvgTzg4x9+SDldamZElICNq6TlnpUya2Mol1M77g8zt7p8C4a
s5A9nk7qag0q+7IoFjbrNNTCStWoQcuyDdImaFAJRBl90kSxTiALpcwPhnexNm6G
LJCGXCoDuRficcd3k5FmvxFRCAXxdTJlyIJfzkU2jyVj6cS/QgbaNtvtrMYzk6bi
BHr1fslJ2dhIuwRd6/G5bcr105OW09ljzpdp5ekaD8EswYkQ42Fe2vjecLRgZ0FA
XBmTwvsIkTywL00CnXVoSmrSzShmGHz+L0Ln3Cn2m7uMcanU5/OVLKWiyS4LRkfG
cPmZmWFK7qB2IVJxQKaMRs8d3qk3k8hPLWKusLIYfQRCy3O3uW7bga8UOsatkG8C
uA/Z0I+4sNkoeV9kUU7RkKa7ei6eIe09JTg1I1WcSPEhY/TNYHVxM+JArv7IPeqZ
7oqS6jsJC90SH2Bs6KYDFV+Fbs+hL9bNRpZVf9sfl0blQFyYEmSN3HcMeOqDUAUN
GSMfOuWTNtY4sKu0LAwVkyTBPiYDfmqNEbmUUOFCaJKTDt4yY83AgVf+TdeJkgp8
8m2VnIaJWbOwsr+QQjzOxrMooHfJQtwgOHGdPUG0zwL1x0kZs53dPk8yca/DPezK
siwzW9fenbTtCNYpIJy4tYw+bg9Uzc4Ycc/I78ZvgYq6I1wpNJc+ecsgQlOBY1YI
6o/9lxeXqJLISiNbAvXT4UH1jJkDhzpn7txyj1zLTs/9A7urHBUH6F0B7alBPtbs
jv5VQKqVoWzBVKZA/yvNMso4xM6+3F0Fcnk5vEjgjMUTZ2wXKwq4AIHOdbG5BZWc
leirIKxZx67iB2ITFF7nT28f0BMj84eCD0JwBGGl4zf+s2qD573BjAwtRAI/yV6W
8JZpyC1jYwDj+hPoCAOW2ILMxjvB6LCLOyf+4hzBhRkVwPhIrMX0+xOsxI5zAg4c
AuI8PMRIcIpE8FvXBpoF8Jd9q3IQO2XIYdvr0657cU4iQri9i9qSv1zokG7XqJ/p
/LIKi0S86cBuEh1lHQcpEW3iCj9Wh1JfSDJQtQmvhoUczvjyFyk3YngUeDUBJKSE
k+IlsEgYlhCbzV2SstyvMQUZmSoS5SNBXL9SD78774rIy8k+th8JO4BscbAG/sBK
3jlNzdDIHdM9BfgsE7JT0LFBXpG9nL/WTIPk+vi9ymgl/GLh/Yky6sYS9BwEiZ4c
HjPn2VIUSN5moEzeds6+yhLPkekrtAcQ+C34azsmdRdNmRKD0OYgPr28LZ6Qwp/W
Mr1VWUVfMLOGj2GV+wq69fKsOHBB55dAjd5DEh+90cYKIJSu2gmTuGFvzyenUYHP
ZRsnH4MFp10jAnOYDYxnk1kTKGethW7SIPu9UkU07trb1asI4E9RYP7kR6Dzu0TO
vCWQ+YXPg4A+S+1iKd79N2c/EiZfSdBdqggR7opRj10qc/cnQbT2bFZiu2gpVA/Z
omTL9P3rcSOoO35EMA1BtwDWDSAhs0m9Y/MHD86zLToC1vkINAgp61X3nz2Q/svT
djvw8au65Mt484KuwRgeYB7wSC7d6ppYPJhvcpoyIvAuBDfgMZKOTXZjh8wpfIU3
56vKxdYQsbwVTjZdvRums4vaIJws4nfVDxQmOCqn2qXg0wXWTFfHkINYOLqnnkCl
MsuCIwsjd0/+ZTHiHwDse7c2Qfb6IAO4rGIAWibRZ3ShEa4QZhcYuVzC15vXKLUy
xdDpFFMLKuKRpeKxk1aBFzY0fz6sMFMYIs2AGRPSHNr4GMdOr8ASJclSDJ8OXjVB
wAZdQIOz3cYSFCx1vEi2jvyCB7h8JWcllB6pFAkqpsl3Qikl1krZj34cTBDEPwBw
a1eMw7WlQaQXPbKA1iVfwrh+a18VQJecck27Wjp/FZXHJyAjVn4gbAu3vCARE+E+
gv7jnD2ma12Hl3FAMDQeG8ySclm4Ef2QWMIFGFFt9q6GF+2/p6T7VzjoZzKfLSVk
O1cO4l1aSv9bykZIyhV81W/1o2MxrtQLaiivXXXFjPeD4qDbObhLXAPYTTTLQNn2
q+xBHKMiL5QxscqvG377vUmBhytKXXwtv/FPrdSsRcEWRq2uZ/Qvlqvvqo+pQEwo
YKScRFWililCVfm0+nIxV42CV9nvqaycYnYKOUyN1YFb7183yQK6KoIUcUpAWW1s
3O6xE6Wa+2YsjI6cEtXcBZklK5ZONVAwdmKfjiXF45hq4Tor7KMveww3AnCzQsgx
y6E34v4p87wzgan4+ro/gUh7DgaTWnrFASsj3AiuXptdqOsXLPuOoOLzZy3zOwGE
1+w3uc0bQMeOGGwIgzh74LHLTVXlBCS5CLXdnyt9+Srw58jeUpvBgkuAGYgcdVaw
TAW0TwcIta6f3EoyuZa5WhCpyqEkIkIilpTKhK6YGyLgMvOz2mmbx8Rqml94mRN2
fQSjJFnAWDrgdL7sZMh7FD93TpH2glbf2l7Y5LiAubs8pvuTxAwrNXuDZ4ZtXWJA
foBXh1dgIzxi1TatAvz5W29lxQc9oxZjSOBDK8mEP32GIR7O35IgwZztNHp+6oCh
649s9I1rjIzt1b/AkLkrmGkEZGVlZYOjiij7TEOSMQFYPcyf1M/KxW+6w6V5pknf
kN0BSxJ/dkyf3pQci9cLYcFJvhuDIJoHjNZFoif+BXFzcdXWZKLDJpCBIWWye/y3
vztX1n6/9kOccnX/o5kbOEADF0fQKsZcq4lmpBzSS/4EnyrUBjI3QmW7JqfZVcCy
LFnluiosL9pPWWrJp92eXylOZLZF4iK3c1if7rAHkuR1mFHmbuCHk+428Cf1TMVa
UHpcPpp7x5t+w+Ha/T1w7jjqu/nXU3F7dBOANrBlBobrsA6LQPZHv2LWY+daW7fz
DVbIShKsKnwMXYWbMrJPy8BIoAp04DFjD2d+pRlP+W+aauRI/kMypwcoTlgtRvVh
37R7c3DoCLpjza0u3cQfn2JjWqoN8hOIh1RhOlQ7N6Cez9fG+ulsFG8vSJojKtGD
oHhv0vNUgFKEe1NOVQQ8i497kBHJzrv4ReexJcmYJje4hwTkYVA2aWfLDEtgijEU
nB9l+SrVq0yEqtVdfOI1pHDqBWE5UO0E/q9RzytEPpMlZ+GwCKUzARXlI4igkNnD
1kOwgJXBcK7ojM6V3UT6bpelZNKNCXT+v6U1/luYlk340f9wkSIVvwZJ5sCLCFUq
oeIc7y4Djs6K25BmZoGUGV5mK1coXfy+0Cs2PxZLXCTzXd9HEdIMNX+SLtlS/3At
75IRYYUL54bbyOMW3GO70WeMaCQJeAzKvs0IHpirfEDZjYbuyx4pQw+Aal49vKSZ
HByBuI80L6sxfn5EYQVz1il9hhj2+jmN8aG4msrUtCWZW+NBNxmUkueCcWxgm9FV
4TBff4UY2sdHF5cFt/lOLq+so05/f8tBliyr/HhPeVX83QDr9tA/Y/AiUQUaGtAX
dSPeU/yxMVBMgl3AZtYH8OGbXOQS4zhbPiUFpIdtVp1r8bQFGU8LIizb1V4iInGv
i6Y1/18q96ieeBV2x5SpH0He/v590xttBxZFi/9G3p5oPE//w9DVUuTxQ+RiWqKU
/hHlsix0ylM0mY1wFfGchNqKo14x0vWWNCZvLfV3q8inTwnDRrP9jtU9RhqoLVC7
D6g5U6NlkHiLenCBz/K97jygoVa8n9kbdYW4s2XjNp2DUnkhXXz01jz7u3GVXOmS
0/aQ79wVzrUEdGJCOC0cfVw7nIH3EuG/uy9d1Fy0t30wcNOw66nBABYq+CBzYCW6
9fh6pOuGl5EtYmg5mqVvaLRgBteonquFelUt/p+tD/be8BogMObGi7GtJl9JFa9T
nOt0rp7nSrFJICO0hKKcMSex4sB3L3iCr7Dn58E1X3MZML6AbLvhM1bmQJ1WvYQo
qoaaRq4Xa+rgvWEH9tj26yKfR1DiHLyfa3wC83plQM/JzUdjS+qratvtCvPKC9EJ
NeXQBTuKWJmdOxpiHiqQn4lJzcgsSDiSTSpPOSG3/IaMdCSXMfQTy5DAyVLimyhR
rs9kh7/WiI2H9A6nhtSPKRMuLNzkZLI6l6JgIhV/yvXZuvv9w5s/wu7+liqwHpwH
9ZMg/MrOpMow18g4ZBe4rjkjFRareS4lYGD6dpMqF/hloF9lraovZ4UNGHOYMJps
2slNPyH0Ri8DvPehelpWkIwAJ7dYbe/Zbf3HLmyBhzcLc5+ryv/YKd+QQ9SuxQWe
M4GEMhgVBSWYMHat/TRl/l7SOVEDaACFiz1tLRAUUXcPfCcdwJKbAmLzWJ7WJtJ2
JZiP+s7MBg5/vW9IOoaSE5J1dIOijo/OphceiluhADQ5c1pdaoNqgLUk4mVoiFFp
IRYrTFt5+WGINFMb5AJ/aZ1n0ZcEVkqgXGT9vmcjhDTAwQl+o9XQWvGiX1Xkuba5
v9m4YaDG5Cs6eQG8NnKMZAv28dWtVQV/9Jbyn52zNRXo0aPKaDECJOKFs684EQ9+
FEHeKaIrTkAXnmiNHYpBAfXLKPHVjJw+46PmUbm1mV2srAhsZGADw5CHbAfBEVNN
xcDA854uUbOcRYFktoKKH0TR4qh7Bb4XEECEaTqr/pC17ntkXKKGHeSuqVREKW4G
c13ojLZNEuZCPW7+ba8bBSmXfoPgQZ+4JEjj6FousBZo3A86owJf/j5/fq+hOgL/
surNtFKxmYro7teyJkxQOsMyVbF/wtm93YfTULma1TwbokE+MhwiS4YCwQewEELd
QeVb3mqRh8ShLHkv+/VhRB5MoruDWCDcZ83Vb+u6NbqJ6FNSYK8DtN7aSnvdGu7H
MbDX84/OvJ18P30nHWsQnewN66xSu92AID7hnQAYWZGzRZPO0m6gFZ/e8RYXPijx
qVXb8RNAIH1bQ0IvJ4t9xns/dYLLI9K2G7oHjLeZbLvIxiazDMUHQ9qM+HXpQPBN
uLW/rex1wKRK6xO13fb65GVPuNCIrnMXKXrtpIz3j/KGoudg1czwG6Y+JEvnIhrA
SCFKeReJFqqVkXlhOCta/lcNEConhtR3lQDaRiKtwJxEc2jOapq8NE+gxN7RYql5
gklAvgMLGkGPb0wp5F6cePseGxX7nVsF4DVptbKr5p+FSsHxWtu4hsVaJtCPsk8b
8H7kqNDQTEREMxSoKGGPyBG5IKAOpxO6JDHpbzZaJbnpf124ZxKmyMatZWTtCBac
ZCxXJHFABRYmA/sQHB+dG9wZ7xJCEWHUjX7ntR6daK+UiNPlM0ppo+hOWybhU8jI
WbPhotHn7ruROKEKvfUhtK6kqhg0e8wJbqHJMVEF1XPY9bHEks8JJO6haX3emLHq
T0fvb0ttZHaY+TJvO7ouszGajsuOUWNQetVGPuNm7kuO/sh4BD5ifhNnO54p3vwB
j/+t7GhHzOgklKpt44WoyD0jVuz+F/H9/dQa6aSnkGNpGm9KezCzsFXJQQ6yeAU9
bnZVSVbIO5PMjULMSHJzblze3h2SSYurCNHDoKBFCuZOuAvojBvkSv7i+uRbMNVz
vEwrbJ7dRf3nC5EgwLXISFEiUlJN+NmqsiikIypdmhv7cU0i2UDivT8//p2fj/hH
t2rP6omiVHASVo7MF/mBeOV8O2xIHiLxQoWMRLl/IgEdng/irQS/g5WtsE5ffnFD
vEU6fM3+4HrmVNzdtuEp9H85u0g7AVrjy2vNezZws8r8Cn5fdFJMmjLXsRe2BlLC
MTXlpm/lTqPjUOVYMHx2zUmDm4efS5K9M5+7ukOhnRksCgsuREXND8xhs4vsd2xp
c2UYYk0i6VBGMr64iHrKWOv/LIOdKXFtpVccUUfril1btidj8dimQW927Pzj46d9
baI71BNtHg6V28nFr9qys76xL9Z0nfafCM4g6v2nw6x5nU9e0DPp1B5tHxGf5LkK
CMAYQVv+GDmrHjz5aHCQoL8wts0EUsKD7UhJhAIvU0CAKKD4Makb26pJO/ZFKzNV
GBYTuQeb/syvMmuvJ+CNtXy5Hqyn45f4d2b5xnAoXvFnALxiqRBdXBX4ux9olqkR
9lI+Sa/0blNZXgtZ0kW1/jTIFuvW/gXQCBgPeP3CQNI2EJYYRaWGDtaZ/GLBB9ju
a/LPqapU+D6n0n9z84QXaqTfhvcOnG50CoGAuRMqYZTjuMjlPUzwYJT1RwpI9uHO
bvCR2NrK0uQslRvwmXcYYwnyqtwdPsYAfZYV2+NHhm3YCGJi5uWJAJBkctgWYQfz
GQL1Z2ZHkoP0QI7dtCXoCrFeHBiSGy8kc+NY13LiuuZNyD8AuHSrS7ysIjC445ww
Xg5xsb8FquM7jr7kWhNRP3Jf2DIn3wpIa9CB24poy/1Av+Tu57m8OqDTcu1jGY4R
rv8lpuMcWdG10CReJuYR+ImAkMpKwfCkNvcrFoU83d/JTYJUbgmm36Tfx/0Zy5OG
uIYSJwLbF55oXndYgBj6/1eokLh+IqxLsYVqnFcp+mmP7l37EjwC5QMTIT5TVGiP
0vzt9RT4OxXr+S5o00OWg6FzRkb3R4LK7m0jloehEg1RkZE9LdOr1sNYgMoufnal
PTCe+khCW16nxz0HN7vC54Qm4NZ6P2t9+CWfAuZiZxIxNuM0dSSkLNCYxLjTxAU3
TQsRQdnDTpr2vfcb6prXMlGhE1qXdXstTULFAaiMGzOSveCegWu8n3146drT/Y3i
RPsy21hfMolMtBmtVYzwd46LnPNvdM4WqeXr28ChpEPpPhe5292cN2BwpKOYO4um
xB+bo/uBbC7mGyp+wY+zdTYV4bDBhV7K48T/3Q1w4JlGkOmNcfXlgOgrTgO82YEk
v+7jRBuvgruowGcCVquGnOfpbYk15o9KIqwIPf6DZbKdrVYjSbWZ2NmpaVycGINE
FHf7d5Oy0IiFSTECe/lwinWvJRj0xv1QCqEmNGEzzoHJCMa2Y431a4WkW7WFRQ9i
gHBQ71Fi/3uQwUkcsjxpXUrcbXdIo09KqciRAvnvBRM4wuAX4RlKr7LurLkrgHxV
joh4w3HOdvLgxHHqUkqIQxlJ6oC5NZCnKVW49Lbh06Vn3PCs0DbKOU1eyGkaeXsu
E/i1luarJhfsUpiaJHEj4QxgZmE7KEa/NT0qsQCc7Q8KD2JK4jlUWxA2FIoY/0JZ
v9gRkJFqjcOzbji6pwEGg0ZC8aDtjcaGuVEIhNRJ7sPXMEff9DuftXKuW3sLOgGY
TtZdGINpyqzb/3gBXa+ub+kLksZCLnwFYp7+m3DY1iK7h2oAwztQ6Fd5tMgKfGMc
8ig/GB1pDvHwRT4OCv4JoL1krkfmPpB6K+ScfYU1TT8PJeAc+C/Q3L6CEHiLb5D+
8YwpGAaUxDa166aAGYw4iLahNubwHbAsvtDh6dItp4MocmiH45ZqDlakC5XngAsY
ZQL8fC6qAtfiVosfoicuoG6dafDnCKE533jJzOHBIwHVB59PT9g6zvuWkldjN+r3
hqvYGiFkWLsfBGb07bQrLeFwliFx2cYh1hcQpi+AEpowCJL2X/PEzxgBjKLDhGrj
qeLva/qp22BF87D5RDuWo9ijuOnO5WxvBtz00B4Ip/FVkN8tuEoSXqj4j8sNxrPh
damykriYLp9DCn8KqBgVeX9DDXICFChzysyh/vIEh6ysTv7Z4NFZ5c+M0GgvNQJ3
U09sg4Cgz4zIGVUL6VspzntGENeRoQqHadlmVtTWKpjw1grPVJEpIFf1znFVyVT2
hwGiG5WEKvg+7iOcXCoQ4EfL+suFJU6JNeDU5vXsJgGRcPwZ7nUNxAYW8xquqPjM
RiX/DzSMe6FYqmYJE8owiwlA1/cELuFGFPpe8Xj5Y33DuAWC/CoNQhyAWC/uRiar
lB7HO8wP+9YRwckIgatBBdnanFocoq1geeH7XUT5zaCXsa9ha79LUvCy7tnxn6zt
Sz3GZKb/oDPIyakPDV9rVfHyeHaFi9BVsEt2wlOUK7Kwpv97eAU/aqKDvakJ6e0/
Mbb9ZsG5kNRBzSvIzcLiinD6mDU2zwsYzs+kdbk37Wciwe9UqbMQwfpAuo7bUfam
iHFu4euud+Muyir1+k9/3fmyIb+Ew4Re46+BFYdpDB5pBR7+DVqY+ntWUgsXyHes
jvy9jP+lmrql4rHUqoeKQXnrVb3+yFSijBcuqFb6DAW6LUTTNvFlYCqqQsx49TDv
o4EXn2pdpf9zg/vPy2E1KPEALn7w9aUYPfgilCC+VxkQngnzuTferOp5xXEKK72y
pDHOLobc2ynXe1GfFlr5H94XArYfbvMNhRHz8LWkAGA3IADWDRAxn8xaNSi+q+tG
VZ75H+F7TJxf9zUsIVBS9tul+I8PmAm/zkVtkC/frsxXlC/tXmdecieJpm5D6UhD
H2UMDrfflG52lRxCYgQ1tbFXR9dSuL927GWvNCFqNwY2BiqeGorizRL4vTPTXUZf
GbfXQGDhPiPtQlw0P9byDuoz6MJz37rGmbLC9/baFZDB4h3TiZ9CR3b0eSXSPu2f
CyqvnnHJoY2iAyOkm70K40iT6pb7tIsnrm7UeNim6bnK4qd/H4HN26LPhtaBHiQI
dPFmt7KqRDOlFCwUGdboZfzicRZ3mLiAqv+as8pbjvojxMSd8SQ3dDWUzYKrV4Ff
btuw6kavTlMGD7Cz6+bzQmIv/OwgbYyaWxfvlqXpehap2wKkxbPBVNtphwcEao/E
29lLfnQOCxGEYVc5DC+b4sHudjn64hMEWVAYxfUJfl3/0gKRyIJyDuopWl4VK0mN
sBGcN4wPJ0KdvkCWP4NqGHlQygarRKhzsWLX7ryxtuWwYQKhT0pFTsuhbppyN8R7
nBuWFaD5YQtt4QhNOyhhryoZUhpC61VESbXLqx4Ynvua6jTN3D65ZMgaesoEJov3
/erKKdfr5U+v+7NqCwmWEAsYJxv/esnTDFzeQqHNZAFji7Q6ZLYFBBAVrL5be2fs
YFdYXGofe7W+LrF+4liCUWXaFGn372mwLzqV9duh3P2/31IfqmsBsRDJUgExddh8
dyzURUSt4phGZuEaFw9tVlGd3wUUBdXKcx0rGpaCbSGhztPcKTIxdtlTiXJXaQFD
UhtV46ZQ9i3UJW/7b1tR4R8ZcQXpxwIcZai88K3mdMmKiEehDfrD31cj+2nNZCoT
BhNIESDvkRvJQ31db9fbvhCZ9s2cLpRUhBNUffVKknZ7Cv2WO8AQZNfImvIhS+O+
btkOSMN0XdnOF8uOx0YBptF34RbNZjDngPxSjY0phuCpPVxGuGk9GUF91mtHZzfM
Kls8gqEu8SItcwFTyAuvHr2ccZ9vXBxs5LjrVfO+f2Awz3CcFj+5T2uZuh3qf1Xl
zrjkedZRMIEw7p0B730utjM7nchjYfTy0DlQy01QMaE7S1fNupPLk6EHc2og47Yt
xBox+tg4x6S8g8o3Jz37e07zfBUjTeMPP3MOiSxYLBY1beGYJnQgOUgOgFwvZuCN
GQ1NNp8VSw/6sBPF7znG55TDOYeTntSVycgXnEy4h1/0EatyqlK6FBoUgB5Fysy/
0qYY3+1WI2wdzl0V6T+6ez/LsZYEZJO3zAi6UxKloKIh+SNf3U3mGRCK0rfLSR/m
105O3DZwvJg3hS0KKNwpGX7Ua+IT/GBW6vEtbPqJcp8hdasXEmmfg9b9N7n85v4d
8NiBqtEU7+HmGQdUJraM9NPxUyUC02rFUH0OpHc+Zm6Fm5kgS2VloCMhBi7GGS0c
yOoV/pL7orPbSMOSNKdlE/zJ69RL92qA5FXVl9BGtbtTh702BM+d4rGfFrtKRIdy
ZLOv5/n299KDqy6cdi+7pK2fspebLRzJ/Dn9RRjef5Gn5YnUCJil9lajw4AkoFhS
0IOLbADlztUpOGZm+RtVkXSWeA26+EF+JCpLY6VBhOBoLYKSEj7GfjdfsNQOjipd
lDKJmqnFQ/Zm8gOiJCnv7/n7y0gXUD/EYEa9x08TUGgPtf/bFEKNVWQgNPqcZc5x
u/tg7B4GwOEVYlVfO6kCUCPV/uModAG+Yq1l6SKvKRwlcFia6fzNju6X48lUQvbO
od2Y6ZbmnHYe7qZPbNk0EGMctrbW5WSihNF1pYqtQgRviXlt0v/iM+GBJ9qSE9WI
9XToSwnOeizZz8iQj5cL1IIzRcrwCqRu9QR1wFzPpp/VK4ROlOs3WN/V+GjBEvhW
9S98x4fEWajh6xAF6+SpysTvDOjgPDIuMmMN1Pd7Y5graA2L/BYXLJMkhBliFtVy
zCSV0u2zN1YXPPe0dN7ZGpnudzRl1za8PLBAJHb5rDznEaHQblH+Mn05GjYufDMw
BsytfAwLuUakUxB7G19aV8lB28MqBM5IB86N/XTW+PmvziRvvDKKHd0OFHSpMNtK
74kHvdWBKcPi66DjbHEXestePFpSpNKAzvhi7ZeWL4XMvaauUhJEqH5//ilWP8A4
NJpThP0w2D547FQSOMh05K9vCl9MTn46b5X0tsBf8V0OKTJKqGtooEVygy3qsMd4
s+svPB3mhyPcoZ0OI3w5iV6PM8zuKqmHYq0fyDAVSOaC302tdxWsEUu8IKJAK9yJ
27hXgkBedxQsn6HqmNX66ZahoHXhpU6/aKpt7YNpYUkjSl3vq6gx7pez+HQ0Npec
XSO+UzSLQn0RS0pps1dp+LtD5YaWb3Fgrgo8TfAbxhco2+QjLBpQUoP2Hk9td9fd
5tcbpUMx8Gk9iuG7dlf2q74YDdNPB+Df3WKPTktOjbIp1VCt9GsQsmushv81enr5
MIVzZxTlC5o+p171ANZoL6rR5CsrTxi1XVXx0uVLOfHWNZEjHK2accEqM2n48t1h
Ozvnhx3A8qH36MTHUc8RFr8VOJdt5ETS0wF2LZLWgYmUfh0XQf9YEEiLWLUSBiNJ
W3EZE7QEVCTB9inb4U0YrW/mmus9HskD5sTmmLs7FbEyoy7vy5eIZV3oRL0QVHAa
6qI3rq7Bj7e/+eEz5wcHy+pl4XIbHXYWzgpvi7jbUIPXAX9tzbr1z9WVKKdcKuS9
AqaIIT5omGJnZElT8hAyfKbPugINBGjj/n1qO/kLrK35yKKiik/CJnGpqAfxOcO1
90kVFTKA+qdlrvSZ8akD/cWv0LXqhzwrrnzlcj9kRKWoa0btADcoxqGdm2RSU4kG
/v423KKQUJTGfCCQ7DXpyTGtMijbWqUFxk0uPJjpF+l96EM83QeqQ+VA3j5HvLxO
HwpEMpd16PWdwFDoHZQ6FeFhAcRWf1U+DU5R2nC9lAIvR6LF0isLUaBnluF7p1op
jk8joLR33kM+xjzGP9IIjnueFBm3VaK43qYPYz3Lxt/4imk3JOkGvyXkLWhH3qYD
ww/AtdDSZNGD8cBD67tQA3KHjZIE2oGS8jxlO2CAdjRvgFFk55Yb5kFYQU1PupoN
Ggoj8xdWZM3Sqqsqtbzl+34gwzCZWEy0SXqUnG+wWaRfJhXi7UemSLVvDF4Vww8f
QJ6XI2eKrnjjk4Bjaog4a8xWo20uahm/43eBlSzAvFnXjHWzNv9v5kwk++qsLp83
uLwqld1efwHSUlPhnpLFwZ1P6r6b2hscZs/LWFLpqF/hDuly22yIIodo81/G3cwx
d0AcvVhvoBYymWC6MEXfD8g2OUFDFwr4hwpVeSpEIj0gOPRzJFWLyX3nliOqZ4Od
yrqMQmOOfXKY+GS22X5t/G9IyfdBqAd9D1sWTRVaXAimslSpSY2bfuQOMZb1gCti
sUjMdbzh0QWWahc57vWjQ0GCSq44IGZY9R55pw17Nb7O/IUSb1etJAJqjlNraSb8
8/pjhi2E7kbL9rkQM5tXU/kfs1g/8iwP/ktJtSUzBKlT4TdLqwpzNeO0SFRUbyR2
q5gbOr1ipKXNcE5bqKwDx6w+TCdmvFg8LZOmjeQMOTM/6GgqjP9zk8Bvj/Phs15x
1kcyL9DaQOJKPPoRc/c7sEVi7Bn9SI5q7oTmky+B4DXtCIBpexIJnPSOHZAp0SUc
GsC1e4fgtlpCyfQ5zCoDcnzPhxctoGhJMoOwjhMIhxw0g7NyriWps/gZ3kqHryWi
JbyTEBW/H23hxTcxKpcrtDR0l9LzrNoFA5v72YVtb8PncRRQgaRfEcCIMpS0kIre
XbnL11q8LozwAt5GBQMXu9IkaOREIwLeQH/oOlfOUpd8zR3Q8BqxGMtszZxwG6mq
JDVGz0ntXUEFaIYbuEJTOoPi+XoMIwH8oOwgy9AJWnwH6U6Tc2kpimGFt4kX3fOF
NuGor+6KY8ML34BF05fUPMHwZROy3HbowtDmqn3rd0dVbo1jYqRo6jelOKXNlTkY
GBoB6znceRpeqM+8IRnnpgAwgBBSCvDS3Zlbw680tlTl+y7piDjpCb5USgdxwO1H
XtshcxTK5e9WVxD3AZMmqFS9/E7P3uTvi4XF+y1kbgiZ0Q1qheyK1fAz+YhiMm9H
bRJbr0n/co5rIszylYsL3WMFZLsyAjpOo7DXkz62cp4YDRTYSLPzERR+VdbXKTFe
amGgZhnJ+Sru/ek7zO+vYl+kvAn1c6ibkZqzKilBBvr5JskXw3nz5gThC9saOELr
bT7c9NvZtFek3vfXLqrN3MSNa2mO6brv044S+QYvP5/w3YFBCBYlLPXK3CYcp+Mt
ORoDHzo0EjnHP61/ikg3W9uVQIwxXM1PMoRaT/3U1x1uMrcSST4H2QR6P9T+jeHw
e15TyrSmNayRwepuxRGggkMB/RiZwoc5Ew35PYBb95JXTSI+Ctj0GDHXn2l76hDE
wxNg9gPq2NHytCyuqqvjETItXIaZsDIXGRyY1MTRVhPbC1ZIEcqNuO5XZDtTfHJh
0VWBbaNvMm5Bmskn6hcHylsP+BfDbfW+MZmC7LzUqdVQZnhGs15Iwokn7ZR18wSw
FD6l96oWbFL0zfxQNsMBxSxNnbueqUcfHqyYJmY9USVgPMOgSz89nJHwxU/T7hSI
qktl0AEhc3Kh4e/sQhQkoJtI+261MyPoekzKNrgJ+gJgyULRMs+lu37Yy++7EoXy
0FMrHh/VFDKD4GDZBzM9OPcrfgFQ4BbPrxTkrS+ok4dDm6y6+QX/TJdpWDtlI0um
4IdXvOTTbjXgpDYbQPAWTXWWAdJvCEn90Ld8DNPHpMvs5Po7f2+eQCsdnm/6dk9o
SIqOQsmHnmNXsqPaBUPI1nggodidXQBq1ue+5Rah0CjBcdofLbwgV5RcL7tg4vEO
iAnM7uHhUnEUnYY2hWpF8FKKIkG4Zwfju7YLTpz8WqQBLj+kJkzZPlMuX1YmBhdc
k6pH+NpUe0Hg6txhNsLtNIasz/3TxjCiTQdjLVJuy2wDKnt3yX9pY3QNF/qoMHeP
fT0leTVffzmVJCB80+q3V64nqJw3AdGp5imT6gEzZVXBlQrOwXCFWKd6t/ejtYFs
X6a4fZ13Y3P0GHhPRkWjNXQ9pLYgPtIFsojKUw3w7jD3G92ceeTXunen446WUUrQ
HO7LGHDkci7M8jkBWHPAgv6/NH51zeIjbfk4dMxZgZ+FSBc2e1b9jecWT0Ybw1yM
udhXdLGeT5WyLlEanekemOhplyI0vDbHydaH5lqIDSO9zZfVjbw0yksRmNONqeOg
SSxWV450QDnC3Zb2Rs+aZ0dW7EcL2iLec6JAtdnfEoAh9g3+WTxukFzJ/qFbHihh
RkPc8QRz2KwScKL42sHjtPYGO9OpeUJ0v+6Qm/3En2T0C2rRmx8LvKEj1Zk8hOXU
hvgLbCE4JXX8PGKZHLJ9xttzrM3H0apTKn15r5Tpbsk+oV22TV+tS2pCmnIJRhDo
cH/OfknOxwopnW4wf1Fm8GefJLyAmkBS8+fywPg5MXDBrVva4xFF2VEOAQmejcBq
g+QhZ/ZElsyk3gBbYp07ROJQQZrldFSYICwMhxCg++RyxY9VXEIqnmiTAo1VYf9W
unIfvkbq658uQ4+31z6dS/lIIjnl1Ne0CFEB+IBslNvDPwt3OKvp6frMWKJbZvBe
zDx8WAzz4jsymQKaT7cYTdM/0xeQ6HbY0KQsOIoxw1L0H6EbnylepeAa3cUkVhid
+dw5HH8j5qyUd51qWlxKWmoHEv6dyvmQ2aCWSRNcXHkbypOoLoc+wb9QSu5gbE6k
mfvJA8drIO7yTxB4lFOQiGlGD4MmJdr4UE/vNlVQJcmFaXK229bXZg081mY4n9Py
0Bdl2307/Ctnf2/0ihQ6au42yKQHgpAnpFt212/lRaSzeh6RkxP6LJxz5an6GNbv
O32zXm+bEY4Jkf9g1xrC/UdImZ+Qc2vK5reyaxCzg4BHku6/txOw0HB9Jr5oimA5
lcRfqs8Bda6gEsbiMzHAvnLWtJwKGtEd/48XshdneIxjwLtvyQeRcZdRv8Vr0pCR
YYJjZ4yP7+mg5PXrvGqb9uYi8qNhWDnBRYc6IHyZQ7lZn8kMHpqrP9tV+JhXCz6u
K7efxKUebXLfAYDa79IYLRq8Mh+131uA/gdOp2UuX9ZAYTBvwX2F0bN7xghBWV6c
e0iRGEFbClZuubWXdmuSzb6UzIfX0bGt+fUeJFfpuBQkub3x7sQDKqxrE8U+uEbk
MPoxrtEgyTcyJuQqCuJzEU+bR+x05aPVRJYg+iRnhrcooiVyPA8Ca1ak/iDaBLRJ
ZaKu2uD8Rs7GBx/FKgrOPSd7Q0f3FME8/cSOqa22+2D9SEhU5ZVvyzL7lhLS2Hb+
v8NptPtcMNuG1OaMKRHiB2L52ib1kTnhrpW7Sshf2UelTAj5nVXB1/xVCbTtVR8J
pem2QRhLPwXBYsFfzdU3PoOZMhzQKgtKwbGGRvGSkkl7EjGUWVhr3SFKMSuBup9I
WSiAxx0ufj7GtkeZ0WyvzoO39rf0ttRjDSlZRgTlx9e81is9sz1g5ZSEKp5UB91D
y4Te+AQkExYwOrQgP83W1RzB75rkkmkj8INsJBIe+w6ZyoGBoDKSqkUxhPVm35AR
2j8XOvJTcPCg6ffSZXZ+PY/nqns3GJ5N1dwppbqHk+PnSWAt74nlOK14gLPLHkzJ
xKc/pXxiIWv/vXwldnNLY5rE40iGjmol/DWRXBUSC8FXMO7VzAWtGj5NrQQSYkcJ
iwUKXIS3rrdr1P1ephVfto4Lo41tktRo2Dbuhm7cbwHLCA1q2VM18S4yg+KDJVe2
emnQxgZ6ET+vQXBoLn/Aim5d9HzOWsjX1/Kh3b9BuhbVsMpIERUTlqBFGfeSVL4w
oLshg4b5b/K9CLmca+IjzA3hzKBQALQugYaC3T0hCvZN+iRMCUNMH+oYzhokIc7h
Hr0u9XqNNBDBDL6sFVPeQ2a0c+kf1FO/nSVt3/R3anbiiLqjKOEuuTpCNJ34Qp9r
5phkywc/yQR1pr+zOvZHI+xtPkivv7jceCaeHL27Wp/t5Fq5BDVkPDJH5mu/WCPF
jx7lZG64YEX+rIYjMrcq/2eBSNruPT8viptsD1jNxbnGetPqB6YiUxlHsLMdq2ft
AB5gTawfADD7EhiT7lXS7tsPK11gFX6/XG7Sfh3GNKIcjR6RQkCv0CSL6zq0gBde
8TB14Gip1IsSKY3tnOg67Yn4dwcCYcpvwvdFLli4bNao3mo0AQl/x6HMXlFE9B3M
Xigks0LVQQPB7e3l/6jjTtOek+DjK+KC+kMMxeSoEUD2TF35pPgcLcU5LCSRSz1v
j47pVU2jDYx/HyzlA6r3ti0OHxeEZBjXrLnRoZaUfjaLuoLEE4Cij0uWfCxKvYVb
jPNjGG+ia/ZhGgkEjhXqBDD7GpPR6CeJfOcEj0B5uCJCRnrEakHOvgdrOCDe9tT7
dSxAdn827s19r5jYtMuyHKHgR+p5fJQa454qzbUd2UmGfzkkCoSNt2qVCKiiAjRk
xZjOaTe0nEMSrt/vtjPBlh9sOgLCkAefOUIGa+dEBwuHXhkjy/ao1scVCrrJTVLn
4v9R4QlAUgXxiJi8tDyuZLc8Nk5Tvm6O+jMRBNY2MiVS6Red9J8I5y2We92szanz
FJZvuq9/Pb32aO6YGiPLqg053scgl9HZXC00o1dP4ILuXUJBFp8Wfr+17Q0M9Uys
etBqH4L6JktvZLgEQb7ExvjP17dq3iATzfPAoLBWj60RKgVbjmJjjXzzSSEv5u6M
TMe8obToiSm/bfYEdt0vf5sPuyzUeC2Ha9l/1aY9jfn73Z0cbQJeb3DiNGpiD5Bf
PcPybpxZFamE5o9p+6kzmZ4bMnk1rnnTZXfCKAPYl75U+7kSsKCcIqLlhhaBEE1w
oE5zfGThByHbjR9+MbNgHLtwCQmLg+nOtAP++FMNpd+vvjLC1r14cBIvILm25mk2
EVAGX3MtpJRX3BzKNwX/cocGMmo98hl1Nv8YTNCi90i7ECoZFfNReDB0/3J/d0Sl
hNR+BBBMyss8crkMCpZv6Hsft9i+7oFpmSUriOgIXakRFiU3G9syBI9jKMqjh67L
X3MfAVwvYFdZQzm5QSpEL+gueL90mojoSlZn6c/8bOJOWZfQct0Nk2+thmkP72Gm
tkMm6YQEBRJ97wQtFVpoQYtJFWTmTJ9kUw4On6Iuu+YqEaBcAMFd0vZ0MQP6MANc
YbHbZaT2nXmpV0v4+ZAi0iZGX6uQ6wA6EmcSYxPXCO3+MqCUSaBXlsIaakVGHMy4
DfbEzvfefzAghe7FU+o4PI9iu7qFMbIyws33Crosgfxm+Fm5E3UbSot5z6C+8DhJ
+9hhG1KNVcIfoINBELVQth6IBkUJRtr/k4UmiWTZXeKbJwLxswK7o51jK/RmRNFc
9ubZBcxj6qv4J/uzOyznyq9iiTIdt6/nxDcTQT5q4Q34fOM7FjdwcBIf172CJgWB
PWuUveSd6ttiTyXEAX2F1hugxZf7vOtvooAnMp40LZyrMLpdJGVD3YLqIMgWN4O4
sB5Y4P+tvkXTZpOZZ+Y2GTBwX0VDIemxeFY+5G+bi1BqrgjPZutqSSiKE91tZ4u6
L2JPO8n6SFrW7RQwRIn/qjWmGjVxun9THwcNPkvZjpsk/Isjf39DKSMmeY8++wje
XC3GXW9eKWWtmN4iB0oVmIyz8zyEJmsYUqejWUK2JD0Psi+9qJHMLW5O9k6SY8ro
lZOHJvjJ6eQPLqbl2pWqX1/hrg8HMYFkhmSFyuRFPbKulAtgAzdgs+5nulGeI5br
rWm86xTBKapwh02LruAMe2tX42LtBiHIbsLmtEf/TrzIgrWaHmijpstvM/MA9TJl
pyHxmC6dmiJE14vnhoz4sNJjcsD2Zae3/C0TEpxd2COHHU8om3jh9rHaGWDlawdb
kbw98Uh+9UTzAvSLiOoC2Mr2ClGqs8lwu19hnZWMSR/mDxv3xVIxKYFA1cOB+MFs
tFlp+PCUhGjfHfHFhXAfaKYDBqRtVG6PKM2viKtP76Zss786HZpFfg2MzYY2i/rA
5jUgrfjkk5cDAw1kcTVXlI5Et9MTUlyCnwSEyj/aNYuhu0fdTkOuRVsrLnZmhNNW
fEXjjAlx6HdxEHnd8tFTsVXC0USTSLtTgg0bWa9S3FB/MDcbV+MUB76v18ILLK0G
kZHuGD1u4YncRShkmCtp1E5jULHuXqRz+OUmTITH+9XHsz4QLt9VexK2NaUFSV1J
8Tg7DsYcVmG1KZIUn/4yv0FyhNuYEJLliiWtDjyuMQ2buQhZmP5So2OyhAkba62A
q58oyhLEIKtpKrEbra8LLU7FvcFg6QVJE1EJXlLKeqpUkaYWimqPKzO54nkKKaZ/
RF6bKp1F/B1BM9wNj8SrISy0rOKFu1/pzxP+TC6QJ++YJ7eZ+smjis9MOvt+knz6
aDLcIGELcjuYHS6QLxTLgWSgeokD+T7qXfGErPx6enSUZ5D+JbWEAuMAghUIBCTE
d/yUshigQSAh9CspDGZJY/vK70OWnYXtmCEe8OWTBRAXxR5+3M1JgoFsS1Xx37Jf
qAQ0LptTaINQqUthy+kBIdXUSJDL+sNkiLH+weLKfo5BQxfe2X7mcwENpTqAlz/S
+P+GL6f83afsVRdCIjKyKx/ah4Q9r0c0aXVIzTcMGowbb40xMbc4Osh5nN8mN+Bq
JUJokcSKxxyEbNMUY6OZEqmwZUiDKQxyKEHzKZmEGdz0fjynWDkdvBPeRawvwMT/
kAyxXzAkdA8li60cqVgkKT3d3lSKcgArNRVRvyI/noAVask+ZCbCoBLs3JelifZY
D8TnqP27jDRD07c2wlFrqQ993AL9oNK3oN94+CCSDKcz3UMwV86FfrVWWNaaF3h2
q27+qvGeyu/E3KBJNfxLyXelk8ThYbzLx2ANchsIqs7XebpSZmttD6LNGu4Btie3
bFwjSEgt32vs6K0rK2iWzkc4MI2iC4vWhuxInDdXtUM97JcW5wnCVKRffJDdpmFL
3BPJ0R0o6IrtKPjiFn+l+KdoUOuHodGogw3C7/xcqQTW3jV+TU3xsdqJdNxM923w
fr2QAUFoDv8zDv1KyQbOGh82uc9UkfbxgJ+i3LKGA/U+xCCVHUS3ZImw+xLLDemG
xjjFb93bu352BqTjoIj5eMYuMj/l3Ap2Nml+nqzqstl5iwBNk4i5k9beuV2S1QbX
BUKLaHZTMOFobeKntg6wPqQvgWLx9ic/Vq8T5CqdOJ0i7VNPq11JF41FEZhFCbh2
YkbXCF9G8AfItBkVeswOtfHeHyXYGLr4XoZhRzt3EzU5hfidljB3VDmYbXCgluzK
BqiNwu5Y/WKiYV4iZLlnk62YJd/NFcObf9p4CI8tMBIUCAJxRDiCyzQmDL7u0jxQ
LxN573KR1n0vrRKVLtgqxJ+Me29y81fpdueV3TMmS+w9sLSfmgR8ZGhME1uUFNCU
66WhED7CMFm0uCE6ERWDiZ2Fl3Y/u43XdcN/2SkGbw9JqB43YWC4K6ly1ioBwCHf
4iwNbdPgq0asiTiPTYG0i2Fib3Q+S0dPIDJOG+SyRpiIxHm8cK13LhvtKDm86epO
PQAZCgxIsYRZ2F+XwQPNiCGhuE5XTc7QUMSsnbZL50jbaRqnFIzhHLFZrYUWzyMB
ewkpfVyoFyUiPH3l+qgyzZNLJfONWcFN7pS3GXcYG7SyoHzisNBzRFQI5bnFPE8T
7bkGgVYIX9ERX47KDkZuX1zknSmvGGHSsOck/3arK/+IGUrAuQkUFN6LP2ESxdFS
reyFcHWQShPTzFA/sQ2Uja6KA+mHOWzTmx04eRBOLrJfx7lG5QFsjJ6Hhb7HOGcj
HkntmJtKWSowMHPFWwP8Bvzo6WWfDfZe8HPW6YWK6TpBrPYohX+xXGoJek+rSloS
COHbepS/wbI8xjcRtM7qai/26bKa1wUK9nNvd1/VcHOVelYcw4URhI0kJhEUF8gQ
+PCDoEgDrOxgw2wqxO8ddz/hyFwRbctJu4t/sXret9gZJG2g9KF1rwySb4DYE9bI
A0PWQSUwixewdpAUFtvKJRe5ZBpbjO5ph0KwvClSlcYoYvgpmL5KQQofk4P9SGT+
FlR3zngHaDXm6OhZ+nONwjXwpS5+lJpuvzdy9Vj2UVte/5ZlP0qQISC7rCkxGcdR
2vUgyfSJvWJnVHQMgu2CVmVcj/bc9jk5KMTf2ZkPmaHuNyz/XS0r6T9Ezcez0GV2
fr879vem1Q7EtCNvyrxCAs1ornQxc4aaIT0q3NByhDyebVF9gPWoJMlLDrle1EAa
H2MXrKlRydpmTrU8b/umrZS2plKasJ6KRaXtlQ98jnvpLwwGClPMrzCb1EajOXjS
xZSesSuW2D+qZ8Li9zit6sS9sJ9diMahV1AAscAyWt7Z8Jk0O/E/qX5+BPEgzAaJ
92MtG7z0znauuBhQBYxbdsEt1lf/4XMC4G9tVeC6CDHHQWPP2XwxxwlAPHY3NEN4
I+Z5VdVWhXs6ICh4Tfucju4tQCfKxfrOlxw5VGjMmEGT51j2DTuzKTsRt2l/dA50
AjVs8K4mKytvGktqiwl8Zv//v1CTT5ILbBA/LbABjkf9lJ8F/q9eO7vqKyX59Iuu
VHjIWu6y8K4KHQlwStC1y573WXO7Dqx3JmcELQJ4rluRU2a3wGCxefiS3BbDJ54d
WbiGRgFF0WA3cWYC+MDu7GJ2qjsmZS4+a2MaLBmvfpcLOHus5QUJwapUKjesjb7O
NwzDWseF7fF0xUB0tw8EDuCJd1MXP+/GbgaH/P6r5qVG/guesqMHIKc1zC26o5Lf
Y95Me1d7Sa3JFmnW/gf2eIYDBJ2fDOo8XO9szpmX7wZFKy1vUOUpOHoTA5Wr935n
8kuHWEsfVJiy4fZT0PnQGIP0CnPbjW3z9jnOS958SwllM61AMR7dH+ZGo4KmVKOp
N1mnTu/0GYQ2Ydcy6P2IaWb/85pep4r8N4CYAh27eTivQfd7PYnR5m0XIJyqSJkT
w0QHxfD4pst0+n9r1w3hKbNYl/GI99l7j52YjeP7LMWDtHm50uVuYXV/bV/LR99N
rKSjuvrvXOp30VVVEDj7peW0WYedxFSOMoPz7wYu1ghfO9iSalWi88Z3JWXsA6n3
CyZuV1jTuyYiTo0hf/Qc++bm6xvlb9O2jqVEo68pqCpbZ3zgXLgJu1PgSnv3SM6g
zcQ+pMJvrs7S2wzt8KVglru2dhmNmahI8mmQRdtONsauyPYbm6Oq5/+L57DCJLWL
8MSi1WSb+ZjCYLUr1OqT+6UazrUMtswS598cLC/p2m6mlAoR228WpirDaUMhtWux
DeQpIoQjT3gOihelLUAdV9gnRcywwpVWHwIXqUK+NP+iloxr5q3Cck9I4urWuAjJ
47OS7R1GFSR8uvseNjp+nxvrokCv7JU23e4DKBzdjzkt0k/qHhor2P8hH/w8MZye
hFf00f1t8fQMDJxZhzCMWtt7/Dd8mOspncuv85JAcbQeCKTR8zUaOq/ZbXP7MrAd
B6S6Z3aV2eYUPJPD99JopUVnmNMN5Gpq0eGsK1EUgOq/HwQf7pr+liIs+E6bkdIU
Qk4qDfgRGQfQQcqqYOiEE25FMqXnK0hmygZq0LLD6hbNfT/ISI8XD5gnPtUxfyk5
tLmoSg5sHhyJjQZrNYn5hZ59Tq6+n67449UpQpUM4g2ZkZCZ0H0+EotkDfkCF5Bo
cK3CLZNiI/bN8hNZJeIB96lGtUAWIQVJm+06DBdUQFYFwD3oZ2Bu0nGhrOA7YuHd
R6+6sHjuqBD9BOeJGfvPDL1WAuhgrt0tBZ7l0XamreAquyxIT65CjmKdYKtG0QzW
bpNTCk+6CJg5uMHhZuYWxQO1+qwpdltXZgQmOS/DExuv0Wl9yRetOcoBn3clY4N+
4EpkBvTRhuZ5VGcsOdPAt8UALabyrrSyFl3oAwGfhmSyPbJGHw/XpkRXSBtMlZ5u
ru5Xx4F/7mpBt+PfnS9KY/sEhiSB5qqbmfXBc/DGfxxL2E82HEfpDaRni//GOYZn
zm44Au5u0HOF5pOtTao10zQil546JSOIqA4SN1Jfmk2vMDPt9MFhzycgL40j7Jdj
jkc99iN/8Ji/o7HHGmgSKq7vY7Dkqt28yAVDbdp+/xoCV3yzw5uwzfkvQdBRf0iP
p/Mirg2gFJALqkalotP8fHgC7IWuIpjPqPcoP3Wpx0VVMi7vZ3HeXN41l4ooTXps
1es7YM72hVTwLtY0Hfw8NrykW54KFvgmWjXKqIbSDtKfTUJxvIjW3l7rkzcqW0rp
Jmu0f5Ev1Jl1GJQA/OtP6F6U/onxllOGO1zjMioroEi+fyv5fRibjyH9Eej+8D5T
7yl8wZ/9DRjczG4DRabyp3N4F/T7I3/BnaFhOHRzkowslod61+gdzrG9J5gIWLdT
lTbVWwraUEuJRqQ6FDX0C1VTnOXQT3wzuGeV6BTDqG2bJ4+9P6G0o777/vCEjra9
Q0exouSqflUKAZ60dtQ6gU/+2hBgFOOE4YBQPznAV4YqysS7F92FMvuVXGL8IMA3
5sHoEhblZ9RDU/2a7Ez+pdwGXtZMeHeOWma3F105mfmgIIC6kgQpt3syKuM3Mcw2
K2U9GCa0fsrJlUuhfd9l9VeM7HCdfI5nmw7XBDrWXB8C0Hj/QTS33QlU/Dwowrtc
8bNJg3TyfvCX2qHn/R6qXN+z7+3wjF176+iWPRI7jwRLm49ex4mClMz0Ezjv+rsn
SBwQyQvRz3aK0FO5qhdGpi5pWfiGA9v/AlBorL0MSlLmrVySkaaTasxjtrNIpvl2
ale52MS8k05frZ0Q6k6ETpc8oSRLdehUuBklLCJUj8vDgaMV4RCEKmiM22ZrO86E
I/X7HnkSfB8HZhJRxaDt8M0FQJyN9Io2yxaIKMoF7ByZan1pEz9oR8u6iBuM8Fo+
jr/uRdOBlf7BLnTIYA5CyOHIMu+SrYBBWTX1jhyxx6C+csKSTqWlP5Zs5DOv3qHq
RInOxpTefENZ6BQLOc9j3pwe0jdaTsvIJcepQUkNmQTL/NSNcNIzROTN590sSQUD
ITA34cYVOKwMbrpUU+3Rsl2PrcR7dtpxX3AsvyZgytDF6KsOF3ZmkDgjqMReSWm/
eLI9NKEu83d587pI4882NzwN3HD+G0jSjCVwDSNHoKL80/145RpV9AUPt3X4V7xZ
t5hVJkYTi3FHwgJJW+oEV5o2qTMtPAvtOe6QByrZr7GT/txntW7VR6UbwAE0pt9l
mNWZjYGChuleuI1MdZ6Wtxesane0ZwDbukWbonqsDCFYZJPK0sx70amrd/jMH0fN
2ybC+doRophJGRqN8qoZ893YuDI2YXFfAqA5+jfTuChR4RBAte+fFgp5SvF+Hd9J
sjo5RPHpka+ff61hINhBLt22kbZAaoNuvjrxZX1onhctiAqQ+ufLHV70BD84aeR9
0eYQt0vFBOkyZr4Z6M2EjHC7EDme6+umWWsqeyyMfAjWKgatabyhRGMnsHyrg4PX
ijgl8HeCP4hju9xExpsPJaaOtZg9q4sSNcdoFwXgopcj8xAa7nZxroXB0kyIL/c5
4KDGxaD1hqQcdeXDUeWWJQGbdksypg67kk2EG9j4mCxO2TdX7rqfmQMwkeJsQwOk
bMVliNSv2Sqc2PzQgzu4hZ9dFxu5pdsjZA0SXj/5Pg1N6zJ607Q2fMXvEgeUrnC+
HMlkH981zTjh9o58v0YckTgQSrox3hxZEsSN1+r0AMTBgxeD+yKYOb2rHJgzT31p
9LVyZ5V0fW5ZE80LxxGMKSK0H9pl0EcWTPrCy4VffU4=
`pragma protect end_protected
