��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħ5,��kF��#��o`�Ylw�ve�ѹ{�S��@Лw��\&@_��9�S��]��}4��<������?����N���M�S?��g�Ǣ�8��l)�����E�t9���ً���&�z72��!?�T|O�Ƚ�����MQz*�޶��E<�p6�w���d*^K���pْ=����j�<�1�
<j��~���V�c����N�����:	������J�������0K��ri��y�	p����zze�ґ�.۝Dt:��.���"f�������m?1c�?f����2Y_!��;t��:����
B����������+|b�)��`Q5-��4�k��{�9�k�)�]��)Q�>��ΜӰ��H�+F��4R
���#n]�H��w"�^�|�53�D�;�����
�Ҋ�(*J����Hk��$~̓K���I���XX@�R`9�U��~�%�8�yK|��/�Rj"����f���m2~�����T�s���p�ɐ��QQ��R�]��Y��6���M�ڈ�}骕xm��S���, Y[�-+M��Ƌ�H�TS�nT��TҜ���ˎו+t��!ߢ���XCr���U�0��HY�Ϳ��r��@��)c���Y�Amm����!(�&'��uc0�NF^�`O;-9�7u��(�4ɭ�9��3�+��!`<R�G 0��z���d�ƦA��~��rZs,��1�3�[�,<��瘬R�2�W�C�/�?����sE��O�ɐ}���X�������X8�I�l��Q S`�b`�
�p�1ѽ�}H����T��B�&��V�oUF1$qN28�b�#�yfH|hq��P�{r�YZ8������8��E����#1*���@�%a��Z�g���"��ESǘ4E�競��P�'l��&�R_��Q� 7�Ĩ����.���m��'*�7F��8w���F�k�ݽ���Ո�7��;Uw�-�TD.;�5�k��D���2�m��O
q��Z�FZK�=aD��k�1m�����+X�Μ��9�B��y���S���>a,�{"܋�&x�D�R���� Z�n�]F�?�\�&�c�qܶXH����:Q���
���`� ؔLI���N&��do����=��	����?�� �l5#��b6>�C5�����I�rVx�h���
R�.F�1fk4��/s�4d6kq蚟���+��A�@�0���h$.p	����of�C�XV#T�a	��h2%�K�ʔ��'H���w�G�&䬼T�aiZW�lJ��k�[�茈,^?�a2�gW�I؅��Ԉ���Z�34�*��{��}��9�I���,`;>�yP�R_yY��hiȲllH3�:��ΫVs\&K�p�J����`�Z��m����;���:����+��3��j��>��W·�ۧxH��+D{Bw[���I�����������$a"W.a��~?s �:'�m�D�T/�1?5��m���rt�Ԉ�\|�7��" ��`�˲�k>HU��!M�P�_ʾ$�&H�eK3Uڝ��	zl�a�v	�����Il��#Hk��X����{���:d\�z㒆@�����4��Rc菠�3��q]��k�p^�f���:Kzޒt?X�Z?0��Y�����$俭Kz�}Q��{