��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb&�L�S��O�|X��0aIo�Og�X��H�/�?CE%�A�^�3�+�75�|_�Q�r�<�<xE��.i�!$��ݷ��5/x�b�������&F��+��
�{�Zb��1��Q�sS�1X�ӣ�u
���r��&,}r� �D]ʓ��|��IT&�E�-C�t���+ʞޛ)�Bk.�Cr$cQ�%O��,�ey���FqZ�8�+-qG���8)e�>0�o�I p�����s�Ϥ.�S���8e ��l��너U��������˗3���}C�Ӓ+�% ~���-���4�j$fV��
� 7���pi��3�_��eJA��

%ֳ3��}�;M$�X4�*sB/���-�A�*� ���@;*���Oj�0e�f��lvLX�s����ܕ��G� .�&�q�$d�#��O9����ʟ��ԉ\d9u9�O�ψ����O����Z��3ʬ#��DO�X�9�!e���ق��
��n"]4���XJb	�R��O#j)����L3��A�+x���2��L�y�ZQ�"��y�u��:�έq��㒬i>� d�`&`i�-`�p����~�I���_R.�xD�#G�8�����j̲ ������6���ߘm�k��x�oT�E���C��q]��ᓠ��#�J��s
PE5.Ϧ_J7��f��13+l�$� *:d��h!�޽�j] �S^���9i�^R�?NW��t�)�)9�[&��^ �~i�l ���9�|�����O���ZR���»��2{:g�#=�lgD,�|��X��ѿO����:�ڈ���p�� �#0�e����\��'�6]ar���+��@�Z�.��.�V��������Bv��`L������]�n}�4�p+���Os�O�d;`C�֪���aN����v����{Ĺ���ڇ=�R�M�z��Ɇ!��W�*�C��o�P�q~&�b�f2[�)����]�P�%�ƻ/Wg!yb�a�N�.��~lX6!ԼjO����N/�U���`�bQ��\���2�9���N�[f���#%. _�0�C�����
n�ǣ�B��C �(�V;5�k��I~��������O�L���������NZ��%�T]0���Ks*�������h%��J����B�^O�u��;�Gm��A��<���0\:���ۿˇ=�.|�]�g�#�ej���#��c�N�9�sI6���`q���p��PK��T����U@j�D��P ���X���@%I��E�nAS��U�&�3��6��� t�� T�����ب�8$�2�q6qI�ln��3�rD���\ =.2�Q��{<�U�B=@i���&n��so�����y:��J�^ǒg�:w�D�mdX�An���§�k�1�D��A0���=�-� B��.\{��f�T�V4��-��|_�M�+�Fj��ݏ�M]�+��5MD�m-to~;�T�|G�F@>��@�e4�{g�xN�&�%�\���2#"~щ��x��
!���o�"|��|�t5*�fn�2<ZT84����Ty扜�zt�~W�T�>���9��}R�}1��w�E�%��*ǈm�^3�_��x�cP��o;�I;Z��8c��o��c(���.���6%KO������yx.]�Y���7�h5�|5�@hd�<*�1���e�
��R Y�;re"����%g�@i�dL�y�]q���:�]]�
b�U7�Z�������Gx�W!dq0�
�h��&[��,
����P��$ �d~������6k;/���+�V�p�	[�Pڎ��g�j�2��{��}��:boo����
���B�(��mI�qn&|(����s�Uh�
��r�!�q�=MD���$0��N� Ir��+W�Q���9��4s=0j���w��xB(W��1��,�`�=��ɛ�T�6:2�A�@�${��L�;���]� +����"J�L͢@s�H�����r�T�T�ѡ�#oP����̈́���[�}�N��֓7u�!lȡL��M��w����Æ�q2�fA�p�MdK.?��s��;��,q;�{����p���b��nJ��$";�x2��������?�G����mz��(�a:�����E�5��m���E��r(Yr���t�=��#	�@�4+�Qj�y!��ء���Z�|����"-mHR��bQ�I����{�_�', h@W���|�K��6��ϊ����w��.�-����"/�����c.��s=�@�n�%j�?�(t�::�"�,�E��')'21@\��u�����:���Ѝ�M�H:T���+�Z��<<5�~k�Bň E��0q��.�f��u��݉"����m��c!8�Sm�w��˺�G������.
�CO��PQ�)y�CW�)HF%a}����E�U�wW�L��ċt���hw?�7j�I��]�l�.���������
9����!����Ʉ�t���ȴfi��2��:
p�K/����/�pN���/���1�������.d��?��<�j��=-�Ɲb��M�2,A(�����0��4�ژL�Zm�PK���Э ����p*�	��̞.d#3���!З!R��$����Ƹ@�t �!ՠP�a�r5Z��NH���-������`�u��ԵZ������8���c�%���e�O��0s4XM�ݙ��ˈ�}��?����-k��X�c��۟Q�z|�����>�X>��U�@��Z�`w��P2�����f�N
��񁸑E
�-���g������|��Ro�m�.���퇚�Y�lr�|~yIu[.�͔.?��),O_r�F�+�����jc�x�r�Wg�!����ǡ�	+_;�RvA)z�[ѭ |�Ɠ�چ�_!�l|�4��vw9�#o�����Fu�h_�Y	yJ���lN�5�MaUb��M�.���]�v@�G"� �6Xf|�EHK8'M�l�?�Y��`����Pe�yφ�����a�|
� A�>��*��L�0�1��L�aV��d̆EJf�Q���e:��wޏ�<�1���1g7��������'R %L��>b$��`N�	�q�xk![Kb	z��@��ʑ<:���'�l�&6���Z��6[hPU�"�ļ�YF9�N6W�!������@V�3'3[2Ml)f��Ig����o�H�5�~���v��,����u��D�����R�>����)�K�RIر$��#<4�G*��A�1�i��5����.�($ ��X������u҈X���0��@�����p�ц6���o�H���%��ܿGTS�y^2��m��6��ĵ�����S���b�~�x�������K(}
�:]!�������C�<�gp5��%,� O<8K����ο=�y8ZB�V~�$P����ڛ��I���x?5Up��Ӿ�5����s|J��9j�B��SB�:撞 #E���\��bA�89���Ff>g��%���)�"v��	�I%Ґ�U�h.]���˸N��ƚ�oFM�	+�_���o�T�4���Ͼ�j�+�����/�4�{��׬��c��kb��{ڌ�z�o޼	�,eK�{����
�-�l�����#��(�E*��.R[���Ua �)�b�S��*.*(=�4/1��Ğ�W��b�e��YĴ�O�c�ӹ�K�$��ݵ,ZX���s	�-��w�@����S��f :;��ўX&e&�!)�vlKĨh�[5◐,��K+��Ƌ������=�*��Բ�ğ���xUC�*$	pM�n��bx�Y���$���I,����]�B����F�w�U�jÊ�)ސ�L��Bt�� ��7Vl�H��d8�[����d��")�х�}�hu�a�.��iC%Qߕ��]Lrč��F�����7���ڗ��l���9����GQ騐��xjRy9�����i�*ۧ)(�/`MU�ϥ�������k��]�i��=e�������&��=ٝ���w8��5���+o�	�� ����@!$� #�7�mVP��8$R�%�-H<�3;��AGy�<�m�8�W]���&�R���ͳX�?�Q��#���ev�����by�/��[����V$����~wԮ��4�7Z�<���]�Y���M^�dg]J�x�G�~P�ͬ�f�t���D�S��u�e�H�����0�R��+ َ�\:�|���煟i��2-�sM��A�8�f�~����ҕ# tm�����R�*��rګ,E�����������ERoLi�ϧ/�ݞ=Vg�xh�P�6c7��c�<WI�,&;�������9�����(�S�-��*JI/b��3���'��X�,�U ��#��E�� �S�GH��A�d�&�����09��*�|,q��b܂sw��ա��0R;h��.M鵧�so�X�a�CQ�'V(�o�a}u�hu���5�<Y���A�)�@�?����8v�ź���y�4*�k�D�6�������� +���W.�B���o=���\��&1��1�p#bo�/ς�:�z!��I�"#)�`�xL���2x�N4J(����pL8:.lm�f����&,0/���V�6`�Hq~#���AA>*�Uv�v'buyX���n�5�@�?��&�
m� �4�Kj��@Eb-����`N�-���MZ?r�lN�|�� "L��K̕'�*ľy|�ah�b��uT��Q���oWh�'��RzA����0"�4e�@�v}�EZ��ץ�(�r�<7w[E~ڪ�����D;�Xj8Ћ��Ҩ?F^�w2��tH��tAw�8�#�И�#�����W��USWƩ$��t:/���/ZI��F;�$.UY��������Aq����� g���F*�S��>DΔ�ŵ�)#n�o@�U�'�b�,D�a:�w��P��;�u��m� �3/�ȺL�j��Z���p��ͷHV�����P�^̻��Wl!$ݒ�R�tsI�B�ѽ��N�����������U?�"�j6�Ύ�tA@��+��xt+��{3Q��Ѩ�����S;����;E1.y,���@�D��s�i�[eRSk���Αbwh�5�*U5ҫ|��D-Zn:�.�KZtX�mz�NQ�!�Vz+�a��[4ԇGP%��Z��&P��Le4�kS��o$g1|����R�-��^��F{�Oz�{G��W|�t���.�ե�\����`,7w������T�o�� ��ᓿ4NaTcB�R9��n	�C�Y7�Jܕ���ܔ�m���w��������.�V���.��=�����E�FQ�5��=���k��HX�'��̧��s��{�j2�����&:�~�㜓�'K�ƴ`AqEH��'r.�.����icG~�dẲ>r�q���/v�o��*��k���nxr�3I	G�D��x:bbr.<I������VA�S������� ���&M�g'/*�@�y��ԏP����д��D��?�~�a,�n�d8�-h�~��V�+�9I�2m�\U	8S�V���d��Q�?�=]"�f���o�����t來�e�&O��/��w,wy��b)!;i7:&y��Yѿu�:�a�D�����Z��[p�]٣����E��$�3@۔�R�p����K�#ze�����<}��uu�Ք��_����β"�vd�2���:�t
�e;h� ��d|r *s��� 3B���e��m�e�5B0js��
*��ؔ�A� �2qk%��$L&�3aHO 	����l��b�A̾����M���^�5��Slg6��c�,>{�,��(��W���.���6�U�ڨ��B5,k`�j��c����(Jf����P4!Ƚ��ctlpM-F���%�75��cx#�覾.���b�W�V���#'���v_�_D��(V�����T��r]�@�22�QZ#�Ѧޒ���9I*��W ?������W����Ag�a|��bQ�X2��G��m=�:�[���9���&?�\SL+��*J��0>�%�}�VA�F�W;\q��x�J�&�1ׯ�..�fڪ���'C_B-�^܋�<F;)�(�W|�M���F
@$H���ob����lS�H�ڭoY<��8��r��r�������Iꇪ;`��	�\}��Q�Zpcr'/&�v����~���&o��O"�Ia�Sx�^g��-�.��4IԜ���O�D��1 N�cQ�$?F�����ƪYE����89��ʶ��>��,�����,#�U��h���JkJ��y3���=+1�$�f�T�c�N�!�R0R�<V�n�x_g�v�	E��$�ʿ/4�Ԣ½���+fv+�A�9�H���J
����?��$N�g�"�/B�u�@T����i*�	�W�X�l�e��s/؊g{�C�i�t���&�dz�}ӽ\�C⧧8���dYwϭ�٨�/V�E��Ŀ��h�� ���z����Fq%<���2W�2Q�S"��1��3�?mߵ�̋m��:��(3,�Mh�e�,U�ůr������-���DC�dX�>�����zp�/
mR�����=�y��Y�'�/�c��zf�r�;�Y҆�Ah�P����܆��i^RK?��5t�	pR�z��W�N�P����V����SY�"��LQj�s��Yv�[��i6�[����Q��\��!-;�L%������s��woxwy!$qƛ�@*�;��`X���9��3������zĵ�r���ӫ�u��ɂ�U#P�� �o�+�e!z���".h4~	H��E[�+�5ґ]ƞ{�_������� ꘉ��e �;��̌pB$g�ߧU��O3�h󱐞�|���\�]��h�c'��s7���'t�2����nH��|�Ѿ�"�`Lz%�t3l!�w5]�/�����1k\MڌwT��Ƿ�����N\,����<��7�����f�� ����(V*���4Y�8�	ˏ�ls��%����&�I�n�o�����
�Hՙ�Ѱ�tUlm���g�n�|io��T����j=�ħ�]��� �D��"lK�Oi���#��A�`���g�&>l �sN�O�k��X�oS���$ٟ;�k,��%ʀ��f1m�G%A�y>�:�q�B�fFz!��
"������5t:�$�_7��:`� �8�d+�7�|)�|$�FR���W��Z��V-AZ��M>|_�*SX;M� �~[�c\9x��޾3q��=��,�d*�Bpd6^P��p�𠈔P��@��_���a�"�w�)\� �4R��P��l�*q�h%b�nP�������n�mU�,��s�|%{��x�2��i/�+e�V�w�>���������ʺ��������b�z���b3��N�������-4d��'�s[��m��C�.C�q�~�_�ާ@�"4꥖�� ����LT�UW~i:��I��ꚠ>R��~d��ۜt�N�(�P䍖�N\9�dkǮ�|6���e�z�"f+��g�Xc�8�[�s,j^%7�m�#�p���9|�i$9��-J�&ظdpo\���d�w`�؋٫+E1��M�?�%	����׸Y��:�g��C�z`G7�;�w潗S7iw��.,���\ݝߋj��v�@���H��&�Eo�O�E��W�+�t\�8�ԉk��2�r+_���t�-3ď����/�KݼQZ�G`��rJ��!������4��4شX�R9!�$�GP" �w���ۭ��h>���9�G����S�t����"ݧ�Y��Am�E>�j}�Z;����$��9Њ6�׺:J.��&��9�+x`�Dyk��IC��	i�%6�o����6+;H�c�ժT ��U�w�LZF*G��V���0b'r�vpc��|�o�L� N|�U����l��װӓq(K�3}��V���Q���c��i�X-�1Z��5O�\����_{�l��>7��/��I�cկ��PRK����0X���=����.ݤV�5�;�yo��^;��L0�	Gq��-3����OJ�>�0*}���ȣdI��f �)���Chd���@8�vD{8���.���V�s�
�����A��5q�������f ��hC?�(R�A��o����t���u���t�;�DU���B�{9���k���%�NeYc��#�C�8��$����
v3"0�v�>W�W:��]rb&�C���J5ȓ�klt��\�E�Cl�v{� ��s��H
	�����z�^�|�"M�I������l���v���R=����ʬc�B���B�(�,�@�ȏ�8H80�s!P<�����}���?Ն}�k\O8!t��Б�P�Y�[��pu历��lW�m'�6�oB�,�u.��/�1Z2m�N�>�aL[��-[�
��}y�M_�N�[�Ծ���3& 7aY�22�/��/X��Z���=�������K�(7�j+ $u�/I�Uq�C!�.W%ߊƑ�t�Xӣ�|���&#K��	e��S�����oEN6Ϡ��� OR�M��/j
����0K��|O4)�w\��Q�~�i>�@�=(Z���0��|KlHv%�]8�u7q �g�j��|Rԫ�Ⰳ�1���mͅ���t�ՏUǲ}�	�7�^���ipt�3R�xG�ޝ7��r��,�T{D���m��c�-2I]������^b��8P��U.��M�dD�C�]��'Q���5�.�(��n��oc����C�Uر�=���3;��*e�K^�0p ����j (:u��6V_���ԡ�OE�(�����]e�O�|����������W�S�y�
�x�E���2:>D�
%a�:N��c���|�����s�Z�4�#��A���� ^�����W����D������ �N?Y;����c_J)�E��N�h<8=D4 ��"�i�E�Mi����-��!�k���csD�N͉.H�&��;I����}���ݨ��lx�+�'���L����7#�S�6b���q�.�1/�-�}'�O�7;��|(�B���B�Y��Ò� �\8�}�ќa?�ӕ(����U�w&����sxG�K����Yq�?q���Z��9�ʈ7�*���y��P�|w}��x��h�=�z��-Y>7��L�^ ~��;l�Z���h� p��B+-�����(�p/33��/��Yn��B��~F7���0����� 10���Nwfc�pu�lw�� ㍟$�7�6�x���������M%v�[����߀�NY����<���KU(7�T��!M;.pqvp�=�8��x�1���l�g���������ֱ�@b@z�)��s��k:6����\s��3b��2v��N4i���_۞�QрT'��%><xO·|g`�FL�<��[AH��3�N6�Q�nCiv�"�z��da?%�����T��x��[_��B}y9Wg�a�s�_I(�9�PS#�J�o�\a�(dd�v^=��(���OɄ���/�S[��\^��U�D?��4O�$gdTh7�<ϞZ%�'�A�$S�=w)�IQ?���C�
T�	�6U#s8���uZ�I�o�X�z��y�$�m��6��PWH��ݟ23��ٰ���f"1��|c����]a^*�A,����t7-�$W�1�͚â�W3v;�a��\�T<��_�g�Y۷V�&l�=K��^�#����Zި]�"6���Y�?��Ȱl�J/ʷZ��z��k��";�t�$(�N(�L'uZL��4+0�T�m��W�'WB6�T�:��:d��вLl�p5(
�
'��Qwt�h�^T%j���;t��w3��6`[B�d�a�a-���'^6��d�|N���D�-v<����٬^Mmx�S@�͉~�W����GSc8R�5#>yF���pe����s`T�s�׻��5N	���w��aUD[��wO�($�ݎ?9��9�{W�m�+��) ܨ�<���֡=��Zg{��Ղ:7�O�rty;��؏�wY�4����5���>��p+c"]n�d�Dp*��eڰ�Nq��k�N5�))� f
pF�^	�L�?�W'�H�]�疁JC%�9��֢4P�B*Q�Ww��ջG��p��k�Xɂ�&���3]l��e��kt2K�۟h�4Sv�i#�\x����2J�92��PF!��Se(B|-l͏e��
#�8�%�ϐ�v�u�O̋С�4��n�.�`���ۙ�/{4#_����@�C��c6ܤ�{[3��ҹ����M|k
�BAj8R�ߜ�qV@]�/o;3�s�;}�U)�� �0H�_՚%#*)�܈�����š�+P��.�`�BޓS7p[��F���?�,�<��`�Ǿ��A�a���U���S��*��"t�>�a�|�z��Q��D� �}ň�`���dKeh�e��W�UV3�8�9����1����Zmڟ���̊$�[�\6ѣv��Ga�sa,���ZM���>�l�j6�NV^�4�����P(�5v��4%Vu�h�Yh���atQ�eū�S�_�n�%�ew��h�G������@���+���w�^D�,O��Ow0�d�	j`�)���o�Cq�����$e���th�3ſ ��C,j�B�����C�y��C�r.��?����t���Ass�6	�V�X���fۜ�^�3�c���YB�i.ȉ,{<Z�&���)Å�+y���|�jG�&l'����9�OlRۨ^߅zI���ս���H�ܢ�Q�k� ��������\}��.��'��R�����������"_q��/��p"���w�Ϭ �p�*�f7��Y B��_U��̲�PEhȢF�k�MRվ�S��rF؂w�n����7O��؜��aȭ��<���ͯ�1�1*��IT0�j9jGd�Er�n�����BU`}Ɵ%���ޅ�J�laP���ofA� �����s�,�i#�"�2�oa��hi��cs]�f,�ܕk8�C#fXX�o�F��;��
����<�=K�B۰��Mem��<��a�ct�r��t�������� ,�oGL�v>���د_�4�\;�J�����*���d�tܚC]tR��*8wd�jZ���/X*3���KRI
�]�#��$�$+�AG�R�#��\gqf�F}>
��T��y�9�,VU����G߶���g�C��m�Q�w���^��k�E�xD{���p&��m���|x�E0ԃC���zvW��{�ѳ<�X��a�w-�P�h��Y��f�4.H'��,�p���ņ�D�rĝ��<@0l���՝��C����O�2@
���Y
G~=B�P��4nŒ��(eK~���&4��V�'Cl׻N��t�O�4����Pw�"<�4k!����x�&�����{l!�&{@݆�]��R�(�1�mR��0d�~נNv챜���&]�j�A�Ql��f3�=���t�<�fCj�X������(HQVt�q'r����V[txV\�&���6��nV+�������)�[�d	*Eo�5>@1T�3݈�A�[���64O��@��f��2F���,L�x�@L�>p
��\���˗�w,���׺rc%���x��t���4���C^ո^v�0qq:��8��t��ν�g�f�7�K���Ď�����&��1"FXd������w
ud�!̚ٯM��ܭ�����)<�ˉ�m\����/�&W@2
q��	�a�?�-\K������4��Y�O���N�W��z����"�-��k�t6��G��)��To�ֲd��-V�qdl��AQ��a�i{�J��!��ᥝY�℃A�q����]}w�3p��@����3��}�T�#v6pv��Ʀ��\��)�Z ,�~4w����i���ͅ+�6�\yAa��T{L���GR.���Y�6�M�������˴�+�o|�Iy���+�����m��^�F��z�q��5LYY�]���X{>&��n��?���@^�T��E	 �,k��Q�k���2W�9����u����<�� Y�_�Ͼ��xs����4:�.�L�h>��7[�L| ^�Uy�N7"��E_�~1����~3��gyUu��~-t�|hn���3;t��&7d��Vv��͞@{o��վ'2���C�J9@̳��ȣ-�_�a
�I�����ÃO�������M��Ţ��m[_�
���.����;Ǌ6a)ey��%�+�b�Y0�)�dj�=�;���Q)MVU0��'lm��> ):zR���l�]Vk��T�b	�:�5DCEF�Տ6�nlmPv���,�GB�����k�ezE�>~����k�D��1����TÚ�K�?	��E��0�#��vD�%	׮zqh�*���ZN�_�}B�
�u@��W��'7��fu@^\˥��/�q f���
�4;�ɸ��A�sw@��D��#�#0,}y����_�~�S,�W��4���QT�{��y�ڹ�巽�gs!�lq�JX�ǔ_���#$��
'�m0+�e��Q��3��y�7�� 
�f/��ѳ(������l��2��. ���'��"�o�����Ϫ��!���d
T���ڳ#�k��^�$�k]�~��Q7�k|�Tӱ������5 H5��wx+�f�I�Qc��ɝ�HͰWO�#�����JQ.�K���ZB�8d���_���$?��_�jE�t��'V�Ieݨ罔.��7u�6� ��T��9'D9ѽK��Xw:DFG��Z[��q�*,�O��Yn2a�o1	l�&qPZXY�7}�\UY�C��2�����<p���F�Zib4�gJ��u�}G�ݿ�F��l��{|�k�����d�f�7o�P��p���vi �j���z��u�o���d%k��M�J�9ݥ��ck�����/]�k1{�> l����k;���{b��,�be#û��8���C�I:>�XI��OU�0�[�M����Ѡ�+�\�9 q)�
o'`�^�z�����a�Wf=��]]ǕFL�ܦ_�&�8f���9�^B�v�!Q肹����Jr���Y�<��Z����ͳ��4�8K���:G�4��L2;����O��]�
��{��W�٫e����2Xoq�W�M�X�&
K*A��O�1"H�?�!�E�Ja�@�HV��}^eNy�p�Q���<���mTˤ$����=�b@Ef�`i1rx8c����$��]�
�] [�ոKhԕ]��=�C�P^Y��[څ�]7~��{V