��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0�����
����'a���en�,�=y��~{��i�#�sS�Z�àx�WW�Bg������𓇴r�b�ex�Wv�c���V[�4+9o]��\�S�������_���]U��J��]2c���L��<e�@�&���jX�3r|~�SrOa�{NR^����y�R�ΏD�|����m�'�m@�q��S��Ƣ,(�jݎ�4��>X���w�j2�)M��&�wU�=�a�;�k����K���b���ʎ�\������E�\��,D�`�������A\]��J�o�A�����^�.�c�mC5�h�9����N�
�.�C�!�V ˘�٬.#�]�	ޔ.�⏩� j4pTMt��U�uW#�����3��ɐAw����/5���C�اDt�����e���#�h�e�W��QyG	��,ct��{6k-���w�Y&=pK]kS�g7�̝WJ� �
�Y�X�K���L �n��ӡoQU�Iy���r���o2k�aYDx���v~WX������+��xe|F\u�R��0?ked�1G���U��'i��Q8{���=X��c�H����Մ�t>�"��ĵP�f�J�#a���:09�n��n����Z0�6�U�.h����V����	��7�4�N龗}	k���!�8���;W�̙Bnz��I��{��?R�Sߧ�	����dx�^�_����!4��dŤr�ߕ�v[���c90��0��������l�����T�7!�F�<�q΃�-&0m\�9�w�H����?m�6��:�WM��\�qK�\L���l������9�&���E��<��ͥa�/��=^���Z���`4�ǵ,���~�tfXL�W$���nL����ցLE��$���k*���(*��_��ˈ���zb�-4Ǡw,m���;}y(R�ü���~m5eG��(nX1���ן�*	WB�,��r�?
����	qv}tȲ��9��[h�5q�`��_��#KбnO�봘��5��'=%�bތ!:hL-��~l�a������a�(�����HR��D���Oɬ�%$>-������+S���)V�z��5��$�w�T��l ��S��R?ӯ�}T_5F{��ͱeҾ�Ȕltvբo{"�}�W$�L���c3%�pbp���Q/gyJw$��!�N�ˡ��Vs���˄�7��Y�C!�RX3�iRr��n]���wu��2	�y�r�(�%��l�1G�
��1F��ʝ�k*gZ�Zw4�|J���΍c��k`�Ք��ehr��5���\���㥲g"¢b�X;w/6"@����@H�l�chvF���#Bg��=�,	����ɇ5o�:�X��GB���*,uo��u�oe�xF��NVWg�f!���q��>�����t�>�k��i�-e�p�c�mr��3tQB��i���}�_�࿔k�v�O��maI�q��FL������3�ys{4�l�݉�����k�3�6ď��S���4ǣ��$�TdC./z�%���Z��JP�-&!�g�U#��W���( <�,��5��Q¨@FՍ�t��'�X|�iQ��m��/���}�G�����(49�!cV��$}E���֑"�����
�"�I�K\�hʯ���`A�ր���DUzY	N�OL=�J���j�.�����A�g��^���2
9�[�U�O��E�H�/g�'�pa���L$A<�!��@�	}ֱ��	7P#{�/�,2�p�w:���e��ܿ>���Hg2�F_bw�:�T:C�=���9Ђj��{=!k�A��H�Ӳr h�Zݻ��"��a��V�l�4%g����b�`O? B_���l;�,�@��w7)!��c�?�����ɰ>b��[ݦ�H�h�R�P7���Iȑg���pN"���I�l�<E��)Ŏ'f+{[G}L�M>�ݢQ�����A	�Wdm	�O�&B��f��>f=hx��9RM��Z}� ��$5V'	�Nц۝I%�+c�aw�J�\4h�4�)q�)z��
�Iv �ƥ�������űW��s���*�Oxge,�W��H:(�1<`�']#[@�%�N�~�Ay�k$Ǳ�X��Ճ�	�ѧ�v�><�B�4����ٺ��ʂ4g^T�R�����`>:QqB��	����Wv́�p�ε�������薩�$�C������6�bq�Hzч\ �4�|H{c��Ő����,ג�l�9����[�+)M�諧L4������8J��M�'~���A�'���0�6�v���m׉�;rI�噰A�2/�emQL��~/I~��ݡ�q,�����)��n����HΎo;[�8MV�A�y��w�@��5��kA�#Zt;�֝��R��p������Y��(�^ u	�WF^_	� ���V�"��i���	B$�N2��x���b�n��iLo�l�I����J,r���/%hp��C<]Nn���6�Ξ�^sT=��an^����#2$�e���@�����T�D�|#6�Mt�0�y��JB����xn�\�f�W����@d\�� ��qz��������������g%̎q|c|�'|�RL���-���YI��gb�c�h׊��9`�U/V��K�k��8�tݮ�?�
�@<eڵڮ�_�[W�(����P&��`?i�Y��"�h:mX��������m�"��3~��8�3읱��F.���lr�-�쇼���
"������U�x�Y�5�-�<g�L3�$�  �͖���nԊ���a:�/�ό�o�?Or�o+t�>NU�"_�c)s���c%iF���%��+Ƃ��sv�ο�b�����tn��]&��{��i���2է����������B�� RҚ`��/��r�Z8�X��5�o��3'6�Ȫ��Y4��&N�?U�jq�>���d��6�ȍϠU�=?����,�S�a�怫Μ��t<�K9���.![E���"���L��yej�N��t�d�e���L`n��yiCY?�Nɯ��g��e� �k�Ȏ�+y留9�*+I��i�~�n��@J�%2���bU'�xJ]�o/����I�v�nHR)���RW�?7�K�6��|���{'��Ŕ6�X|Qi��J\,@i'�6>+re5�����J�9�}��9SRab�|�_�Y8�� �h��=�u��F�ѹ0�O-5o�9�)la�5f��`�5c��e���s�7���q3��+��~���i	�	
�J�Dh0�����1|o-v�RK�iϨ,vU�+^5�?ƶ�t���m�|�(���d���X�j�
9�J�jMο�8�c~S��Z��yQD������q�,���"���g������|�926���Zt����F������(�^b\?��� ^X$l>��f�U��6�$^���0ͭ��o� ���>�ˈ�e�&�ޏT1p�{�a	���4�I���F`������p��D��`�'�.MI���5'�����w��Ӣ����L���/�� |V/������c�<rA���~��>���4Ѥ�ۺ�bnd��9���=W6��D���8��~f��$��d=�W/}e��y�Kׄ_ZU@��i�=�z�Ѩ���CX��=��O-����z^`���"R�6�b�4�)���Yhr�|���>~M<��
r>M��e��ӟ	�V/��g	0p�� �ߒ7Z���\*�wv��4�AI�!�G<`Ҿ�}4���g0�q�5,I��C��DfZ�B>rڴ�H*�$q�*�=w�{f~3���!@:*�jG�k>8<j�͗�ی+���0���Z�l��js��]O��rpp/کx�>��OQ�m���qB���4�B�K��>O��m�"s�]�^C7<�wl�Xqu;y���~{�s�¬7��r�������	�ѳ c�O�h|;�om�'��ï��VH{j�z��z�j�ņv?�o0i�}�ʍ��y��'��8Ɠ��T,2��]��U�w�����w��E��1�B-��8|�P@�x��wB0�ɐ)m���J@3-	��V��S_���1l�&	��H�Z�B�%�,B4}fY�$���C݄�Y�D͕��zL�YrE&���%��ڷ�k�����,#��M �žF�A@Z���'���4&5�-��}����N[SV��ŠXd����������͇5���yJ�\$��+�`�#3P��+�|��M��Ö1XPHу29"�߀�<0�$=0����2� �nW�&r(~�?;�u]1�%;2��|��ψC\�� l}I��m!i$�� �+�b� ����p�H��*O�/Ūg�޹��6*�4�؄o������S���q��޿T��ܳ����T���k0J�|Gq��8_xy�e����B���o0x�� �:���/W`j��*�r�Q�{�"o�AF����z��0�Y�
&�7�T�