��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�kw4o�e�UU���׮\m5N�5����(y(�~9a�U�K��<�w����GO�O��U��@\���{�p������}!�)g�-�H7-d���D��������(n�k8Z�Ř�-��������{�Kݐ5��������Kr]�:�"��z��Y������|#_G�ڊa�d���r��BK��x�K:_��o�l�L��i��a/l�0�������9��lc��Eץ{���SBZ�)�4o`�ֶj���qψxh�	!�h��v�D&�)/����څ��2��5/˔�h['㑣$�;�=���v�ʴ�I��B1r�K��?��~8U����ߩI ��S�+d,C}��z9��2�(Ǡ����W�W:������~�����yZ��>#��]�84
�wdk[3�i�V:H�خ"c��a�����	��`�'�����=��gv�EIk�r������@Sg�
m<�w�?�Ie�%,@�n ���<Ǵ���#�g����� E(� ���us�V��QلՐ�%��[����iFE0Z�@L�2:p]��e�����nGSy�Cgd�~��/�Gd��//��k���<��9DN� �5��t.Z�z'�����5���8+�����DG�ѐ�w@�/�P���_�-��v趦/Qʿ�t�Ϣin`~�����C����D_�#-��������䤙��B�;_*V�O��ln<C�s�8�J=�c(���?gs\pw�Q"��<����6=�!�^�p��������8kZ��N)iS�"���L*'M��z�t��[yOF�Э����b!If�����[�@SR(�q�3�[�;��i�� ���.���3�}��k��߆�P��cQ�˧��p�U��bs�%��L�FV���u1G��<ƲDO����	����ُW�����n�V,��`6�[��."l����a'���	�ƩR�Q��UzЂ��b/l@4x�L?�(�+��Ї���ǓuO.uʗ���q ��{�0���I�n����+���i̛�
��![���0i�	:�m�
��$����������b�G�(�@\�p\1��0�ԍ�f%;�Ď�7t�U�@]P�4�9J�^E�n��E�-]�L5^�ݦH(�5⁠+w���Ǣ���x�#ߠTc��:�N����%y��|�0�ɮ}�DQ���ͳ�����D��)ĲH'{"�p����qshI���7f$l�q_�Bm�.v�o�ӫ��z�~�����v��1��>6T��	���z�ͩ
r<N#f��S��MQߑ�`�"^%ܣK<�3N���a�u�g*��E�j�W�$	>�	�H���*q�ϙGNDN'!�p����R��.���EA��Ɔ���!�n�A�(���#�8?������W�����/>�Q��cD!������:�J�Q�J���u~e෕z�&���;�����5�A2��P_ڛ��,��"���=�>�!e��=n;7��{w�:�G�Ŋg3�ǗAs���w��7ņ��=�"���XLj}���Y&N?q|	M�j��OnmC�ܨ+6��IO��laC�;%F�=�B�Y!�q�UmY���-���Y`�u�knl��P-A�!������.�x.���ERW1{3�f�S1�
����Fj֭�")���8��n�{��a�e~U�C �O�Z${|>u�9mZ���^��]�~�����\�m{�@kX(��J?��g9	/�k ���.�9���b����=��a�b��v/L��>|���;M�e�m	<0�h7c,p}�	d,�X����i��:�D�
��qIr��:����#���
&����=�џ��!J�e1����Z�X"�2̈��<��q$�_� ��6X¬�w�UV�U��ȭ����h���=�W��
�  ��]�L�kC���όQ�l��[�y �HY^GZ�L�|9��[5e�<��9p�:��<�K�n��/�p6
���A)��`'�j-ƻ����%�]o�����׈�tv\�_X�QXjs��@��A,�e�1�8c'��	>���#|h���n�*0V�f@c�T���[�6PGJ W���M3���f�6.M���P�@5�X%mu������Ұ�%��������mR�HGx؁	�6Uӎ��Hg㓍�*	���}�Eⶹ,)��`	G��� j��6�弚˥2�۞*�y�QO�����xK;�д="|&�6�i�r3�3�T�<L��o�;�ӻ��m:h�բ1�ɇy��R���n�ehc�d�]Jc���YB[>
�ʡ
���",�B�;��m�³�W��2Sg�'��L�V��5�M��h�Ԃ�@��IZ��Dn+ν��Gݠp�8v�3���cJ�g� W{��@F�M����@�0Wj�^^����������UbH9�Α�l�qƈ�fh�\)�1�w�5�'R�q�Sa��ڹ����8�N�}Wq��J>�yZD9uD��a��`���C�`/q��J������d?��CP/�q�ͪ��>IY�`�:
�ӻ�� jE~�����Z<Y	x���p���Q�י��b`h��F���=Fe�YSF�����ӵa�1Zv��7zR*d8NL�����}��d�mG�'���Y)�ǥs6b���_Z}>䠜�T7Ż���&BNk�Le�~�r��`}�X�"���;BC1Tר"Ge��un��h���t�{��rtx��X�JGҙ�ƞc��4��I���W<@�q�AO��
���k>k�ȼ�9��9��k���\,���vk�g�5�c���GһK��ꁶ�A��p��щ�5E�.��q�l�2U��g����]�,w���~��)�)$�i�Б��� 8�8Gl7p�Kײ͢�|�'�X�r
�[G;����� x���n�|--��)�#ї4��	����8�FT%u��qC���L�^�:�`0l�>��x�#���� �z��>W������#Μ��c �>�|��s6��Kt�[/����\ �t�|��g)ġZ?���|��E�-�"�Y��mQ��L��MqR�5}�1%,U�ԫ;����(�@�6���i�_s��?�����:��Fd��B�bu������A,�,O��h#{ۊƱ�zr�ti�������sʗ��J�N��S0=�����N�O��m9��!��=��v��?���i��{v߁�ݽ���;N4����CR�_�-h9�uU���`�u�B޲S���4���Y~p\������W�Iq�J*V�WM�}BU�TM&���ǲ��S���}t�d]�u��O#��ؕ�ۓ�h�����㺒п�o���=�y�P|�ё��+>ʷ/�7��wL����"a~�	:��A�}��L��<���{d��,	� �,��F�֨M8YS�}\�G����R� ��UqR���������^R�ֳ�#�r|1��	˹�r�pR
��TY�A ��i[*��xSn`��!�-�����	
b7�{D����l���ع���T)�m��U�<P���uA�N�I�łQnӣd=�^�[�D#㎃���8�o�a?�uW�~��&�ڌ�L��B�hDH{n*-�[��B�ŋ�9 ]oF�S�~��j�u dU�d��m7�?dE䏎�o���kz���A�Ԗ��Tt;�Y(�Q��q��ɷ����GL���!��+q���W
)�w��]�i��i�b]��F� �l#Anln�cz�]V}��#xxI��{���
�/�*p�X(
w��N5�3�N��0�/$��n,�!]/�K��ͬ��ٙAt%W�-lK���k(�+& �~�@��f%��!$����/z!MQ����ܬ�׳At]�+�$)O����p�mϠ��D��0��5����g����m�X�A/_A	$��M֞�<u���k�i�2�!QP���qTJ=��k(i��pבz�Q[e�H���x�*V��n�yS?�E����Y�I\��ޒ�yfh�DK[��P�/߬=�\˨���>�lDc ٿ�<�}�rֿ�bra����W��B�!Q����V^kZr�.�iru6��*d�H�N[�RAPJ��j>	�K�5o�?<�ǎ[T��/�B�v֏�>��Tn���+�w+܂��t��P���I~/�:l�b|q�[&�(۳fȭ��}��R�'a<!1���wx�C������3�����'1o����iL3i�$jA��.ȳ12�P-K_�m��q�{$��"
�d���1� �p�|!��i��`��(�~4ѿ=Ix�j�`O=��7�� �ou'K�s���:l���w["/Y\#�GNh�b9A���J�9��w2������^��(V�/z�
X�<��1�{��=�@��ě@���(J�d]��6�p;&��YA����K�l�F������L1�ΏC���{�J7,��jߡ�`a��"Ae}
m_YP�ak����+�(�ӫ�R@(09�&�a8�@5R��f�� �#���O����(Z^f≮��ͫ!�U��s$d�ز���De2�0�l@Hg�����*���5Cyrz~?�ql_��߹^�t�O��b>t	T+��$��T�_�HK0��P�ҸᲳ�댰IJ�2erƟ�����F}�8�M��D�
���Y�,Q�U�gp�ri�9	G��h뼒:n1»��ǅa�c��6��r��Z���Z4�l,�i��n�eK����ǝ
�NY�O�`��'��_�_�C~����vFch�BIx��������Ե��	U<e���4P�i5�_�B%)'�Gt ��%S���q �J|��ѵ?���[��|J{�fXI�ii�E�ؑ���:�����K-�?kI`�C�<}�g��&�D��Wxiq����WHG`�긎QHe��2��W%1� �J����7�pS{�&�wf�){lC�&EJ�V��tX�����9�b��ypld-����j�B��+fD�ۚ������,�B`����x�5G��4� <����#H�� B����Q�gb��H��b�%���y�0�T�p��_�ŝ�P_��W�ŧ�&Ď�>w(�Ed�ѥh)�y	��^�V��ذ]�k�{�	8�t���R�ʉ\�B�F�lq{�*��;˿9���W�=�}3�7���c��1�q�8�SĽM��2{wt/��]@�'�U��+��3s���?���+��e+*�N�ߔmMR�3��^1��
E�c�Tq n��'�e�H�B�ɧ77l}O�:�4� �B[ �ٺb�\��6��B�� n����X��S�4h��M�qh�?k3O��6�Ҍ�6q֤t����BUۨ�ЍT�����P��4r�)C�d�,5��-J���s�r�f��� 3�g��$��|�<	���&���r,f
pIȇ��\,�������D�� Iw����WȌ������[bˋ��t
k_�_S^zn�g֊OPr��O�䚨�Qs9.pRԟ%��x��h$mq��1r� ��1]�AB�"�B��t�f��@�*V��XPz�*��^#�M�U�I��uL��py�����;W�DdEu\��b���lA����`.����yIE*nÈ�P�K�1(T6`��E&�i���.��r�@/
ZsK���d��U��ҭe���D����eG.k��|�x�_^,��6ָ���'<�x��}#4?�w.C��WfܮY��7T#.͉���F·ǞO��9?أ���jj 
�TT�&�ұ���hc��e=b�W�u��hZl忧·!�(� ߿��Z�垂� (<�/ޖ�M��G[��R԰�Rw���H�9�-���r���Ԩ0b�ټf�f»=w����榡�R�`딽d���8�n�&4�̗�K*t�qU�'ؙ��܆�Z_غ��.�f��D{�*W���=�+� gi�=��h�_��j�p�l�k71P������{8��oC��TvD�b �Cr��6]J1A,H�i�i�>�q��>����G�e�x[�3-�*B��������:L���o�(�~������E��j���!����%Q�� H��=�PD�t&�g=�u�6)�UwD��Q/��R���˗�ؖD�=ֹ���k]�.<X_���|�D�)�C?��xS���n�E�2��Ew�%��~L�J��b:<��Y.ϗk$PǜY��D��FscC������/��~�Y�X8Pw����U�j�ˮ���p�Y��&�<�	�f�	��~�ns�˪���
�ꡣJ�܎�א��L�J��y�3e�3$I����ߍ P��۲�gGU3w���$#$e�a��J+9d����F"����uS'5T��K��v�H�w�^?g��eq�f����d�Z��S�S�5�]����̱a �k��	�[��	�V7�ZuL�U��q�g�"��g�@��Ȗ�#�l���3j��hRTU���r�7��W��e����Ҋ]���Z)�G���ϳ��Z�p���T ���8�	W���ỻ��5�j�_U�jeJȶ}��3�`���U�4�w��Y
lwN�?��}	�1,���rcL���7�-�W	٬{�r�riႚnp4M�iTj�-%���L����� �/FIP�r�|����������u�+�qw&m:ꖸ{��9�E-�sХ��e�����>s����&Hl�\0��H�w�d�x鏅N#z����d�l�}�J�_G���-�� kA�NLEy
_�~���Ű�^8#"��\���P_b����xn�+x����!��_���1'��V�.�~�v�M&�d�/�!�k�&E>�fc�6Qԋ�WqdhK67�8�f�u�0�98�%�e�W8`dFXfnւ�{{~��0�aO��><+TP��,@	0����o(��^4�w�%|���ׄ��Ö�@K��]U�}��f	o��ԃB�^�P�Z~!�P���	9:n�H�i�1�W��UPQ�8!��z����m8álm{-\U�"Ar�L/<�zks����QW��F��9G-U��ւ����*$��8�oF�����V]���U�\G�]�nؘ�T�$���c{=��������>��9�088o�$&�����B�]OBݳ��	��y����|`��$�$��G�`>K