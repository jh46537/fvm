��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S�VJ���ɾ GK�rA�!��}�x�E}ݨk�fի�u�(���L K߲w�.L}x1F2�#5H�:�'))�6_��\j�S��W��w�.㆔�[NQ�6��iM�@��9��eh��L�@�Fb�%FZ�"e��R���W��@�s3a�����膂Y�:�D���!G��j	�E����}��Ui����kh稯ka�"������e�^��6�ɠ�Ij��-���jW}e�@,��=��\�`�Ǩ��:>_2�)����������t*�� *��%/��X_0�2�KwS9�ڪaԟ�	�踷Q����Z�@Z|�歊�)���ܰ�K���"F�"�;�ŰS�d&>�،4j�o�9���xD��h[JH)���m�tS����\�ɑ� �n�{ƒ;PM�����>"s��R��m(ɠԉؔ�W��6���ߜ=�5�%�_��+*�o/�Wv/�nW�S������50�u#�����=�O�3b�w��Z,L+F=5�'�?y{��yN�2���D2�m� �p)*�CW��F�7�Ye�ȼW�xs	p���-0Gnނ���Q��	��q՜o
����D+�g��!!|VeG*�s�1� y��!��FXV/ao�
Z�#o �xE5�_�=��جƒ�K����#������\?xi`i(d����#���&S����$��a%�o5�H��}\�����?�ՒI�W��+|Vz/:�2�T�K���f?�k��A9���d�̺}���6���K�����T�ʫ�n?�塲������*}�Y�9�{��S���c�{ҩ����H���qn����qh��W�"�&sL'4Z����B��,8��w��BFd�8M�Y�b�oe�Wl� }�$�ՇD�O����r,���1�υ�\\v��<Ɗ��h�L]@�'�Z{�e5��w~��t�qJsP�X�q)��"ˀ�-׍����������@�(� ��bx������O�3�Ӓ[O[	�Q�����c���x������_��˸)��+��hNۚ�-�4�G�[��T ����r�͸���6�GY����G��E<Cn'C@>^=0�DFj_�hEň�
����6Yv��ݚ�n��r�'U�d/"�OS����<�N[�-��������O�oH�Xd�K�qF����mʞ淛�vKBDݽ��F*m��W0��iH*�SM�-s��a�fո�5/?�ز�yw����Ʊ�^3�T�%��ޮ�~�N'kK�u��M;�&8&������0a��B��{B�t����@ֺ?n~`š݀۱�
���
��ާ���2o��E1��*?�X ��1֐��g�0� Z�(ӖrA6��r|�5���"M��� �zrU�Y����A��-���Ӂ�Q����Z/*rl8g���1tFC�c���$	�����K�?������5w�"����xG��i�&�k}�k�*|}Ӣ�#K̉|u�_&�o@&.�
�\��w���ߌ��L�S[ {��3J��2���F�م��%���}~t�:���]�;�q.~��j�+i��L�_|D�s���Qa�!�_l����=->݅�����()�L��̾��94�ċ�2C4�N%�*J��&�+N�,'/0�^,a��]S����;�A�H�Ȍ�6ua�=����F��%T\�4���K�I�2Ӡ��R�D�-nt^4�P��y���ڹ,]�j� <;�f�I���\JY�Y�����Hu���RK�C��p�2k�a�M�Ǭ�uR c�H��(1����" >��[:�
�⬿�(���r<3Ku��K���{�/�6���w �z��݆�����-�u� R��o1O�[~�����?�b��)�9��L�	l�vh�/��?�g]be�*N���)N�W�ZK��x�)`�*R����6@ID`����vFګ7��*�^�ck��/�عx��Q�
>�]I}�b�&D%YD�E=�-������m�c"+�d�'i�,R[��a�p�O�2	6��c���~CÈd�BRAڬk���t]VKĕ[�ρ~o��������1��>�t����c��x�X,�F �h��������ő�s�֓ 
N/�m�y�VC�����B�������e��ѱ�nBx�P˿����H)�������p��W�Ϳw��"���4�Z���?��m���
Z�a�&5�=���Ԩw9�����j�����5mM�׻-�z��EN�C{>�@/�Gd�:%xə:�9,���̀C6t� K�Iγ�.�����d�LX]9B8T�R�����l�^��V�ӆ�i��4��g�s?AtH;?�Lw-U�yg���ủ��k�0� �"����<���o�dƗ�pBg��#��r�a(��ho���V,�b3�u@2dk��'<�t���GcV0�]��,��-�p�Sp�t����b(��]�n�zd�N�v{���G��Ԩ���̤�ۋ5i,�Bf�7������.{Or� �f[�}aq�OP����8tj��I�(��P���Ⱦl�^�h>��A��2�?Ef���!��Y	�\���<Ş�>��z�4�E+x���,�J6V;1�z���0�?�^��w�r^4Z�d��"�]/ywN��V�)����v�4_u^��?����0��� ~n���/��<7ak���x�e=��v(��2a-Ep����A}��,��h�Ӻ�Mu�h;8U���f��N�z��̡3��5���/i��)m1G�W�`XB�)ʥQ��(Z��O(�.U|�Jk�;+���׶��������
�pu�$��G|%5��v��V�#T����%��/�CA=0�XD>�� mieC;���tm§{BT�(ٰ1W�j$�%s�^IѼ����/UG-vmgYy�o��lOYh�J̢�ٵ����ڀ:��#�~Y��u$.������{��J��FY|��\9�"1��<U%��]��|F|�}�#<���s)�ѧd��r�)��Zt�6�⦐T��q�?����o���H���MO<�
� x�:��f��X�sp��%r��s���}4@��H��H�Ha�s���,-_Xi�ڭ�Q�Vc(	pG�(��5�<5kD����������4S�L��B
�w���54`�x�k2�����/fc�§)��[n��^}"���)Pe�K�z�'��73����Or�&hr�;����Xb�S�v�U���.��(15���D�r�L��a���t1k�[o��U�K2<������?�o�n@[w���ۖ>�t�dӫ�6A�덮.�-,UƩHu�C�Ϥ+���`�T���T wU��<�[<�Sm��W��w{�'�m����vk�$�v �1���ڨS�|Gd���m����}�]�ġ�)ƺ��NB�h��M&�1w*���<
�������h�(\���t���j���߻r�n<F�����y�fZ����=�؛����B��«�a�_3Ȝ߹��z�>��
�����<�\�B;�k����w�'5˵S�-V1��j('�y�Dz��Ɯ����Z��LȄ�q��h�4ޢO���Lc��UA���"�
/W�!�$Z٦i"NNcۡ 0���>")S��niֵ�wE��p�����7E���]iKT�2��+�������2);���p�M�(�1�-�ǯ�2R�kzے�޵��7���
�Nëj.ج��d&��8�}�28�|���R2`��O���g�� qi� �k��ß��<�����9��|���A0�j�'��&{�F�J��S�.k5�]����wvH�}�p�$<�V�SZl�ȥ�P�[Q1��H�
�R(kW�|��	j[h�I�d�87KGCy��`zahkY*�(�����v�GN�Aα!5Ys�m�=�(���X�V�d�Ğc�B8�8����w�\�|Z��[k�~�&K7��9<5�Y����Qd�V� ���7���ϰ��5Wݤ��k	�y^���4ûj}2��b
��)�|"��o0�&E��pF&��_f���'��Èő�'v@M�I�?�R�������_O�	�t	���<]��!5�[:ur0CϪ�������Iud$���fVo)�A�é�l#A�z�ʠQjk�.J�3�@�Y��2�龜�8a��2����~�I��{p	ؼ+Ss�Í�bq$%��ﲗ���K�K6����a��g�x��3�p�6"��C��2��tb� ���tI��%���"��Zq�rF�"��HӺ�	��{;��Gh&O=s���m5����f�>��N��sl�c�4ҘkyH���9��u"Ƙ~yeR#�D\��;���62�󿅌���)_تt�ӯ����O�lC�).��v�ETc���'*�����<'BLx�0}خ.�5�j���3�>wI\@�F X�yWf/���ܿ�s�-�����p�m~��J�R2���9�Q���_�ٟړ|r�Ğ��~����H�l�L[��\wec��RG�i�JN�do~��/�mr��j�"�R'xD��T������$�K��c�YW_��
�E���O�/�dG����і'��iЩ������9���:����Z��K� �?��v����6�e_�BY�r%2�f���$\�!��z9k����H망� NE]�\>o�0�J��ƀ.0�ޗ��~����0[y�{�epzC�eQ)�H�M�5���dG�X��7>���U���j���V>ˁ��v̙�$uZ���"�h0�B{���k-�~:�)��P�usF���b�(+<	��n�Y/�o�#���J1�
!���>|����DY1&�:���ƹ�.�6tWa^\��c2�?ӂ�C�������aVR݁RP*c�g9j�2+�a�W�՘R��B��n[_���;��-8�ʺz�y�y��\o�ғu(c3�8-�,��������[!��|Q㭿�bgo��3��R�#R���B��U�-��Ǉȩ^�z��(�E�*Ѭ�acr=�E�H��s�Qo�"逸L�7�ᑻ����G�HW)�C�;wY
}������%z��M<C���K ��Tv��\ y��&��)�?�):�r���x(�PX�_�O�o(z�Oq"8�d2�����Zp���Y���{�Y�_��.R��ǒ�����e��Pn�.�<�`3+'	���΁S�l�J�,�-c�s���i�mlɄ��?�g?�̠Y>��rA������G���L�o�" �7��_.J���R��@�!I/��E]���q\�R���F���ލk*��P���"�^1\����Y���BI�2NR��(�A�ۆ���4,qN*�~G긄<'����^su��n�б����))�W������#�71�&�^A~tí�z
+��{����ϓaqHnyhkҭ�?N��{�L��Yпm��h���5\��ߎ���L�Du텩�[���٠g��Z*3+X��`M�X4���(F����`b�6|�H���O5���'�ǅϙ'qh2j
tt��
�J�?T�<�\������؀v$9���Lܸ(�DrRd��QnQ,��>AqG���6�Js��T�������ˮW#���.�:��Xrx]�I���*4��o���z���$����SCG1����M�X��������@\�=�T�rGî�?���OY�e��ݱXl�~wA��oؤe�QֈJ��c�l͜����qUn�@�ݳ�餀ˌ��ίuz+�z;��|�K{���Uz��R�Ť�Y�L�W��߅��N�B�g��Yss�8�ˢlhᦨ1�3�8����Gtw�L��ʖ�}���:G��P��V[���ʲ�ջ�+���~}n;��^�K3% mKlmO���(�j$x�L�Q,��_��%q���\�w;����0*N��ˏn�Fb�CN���d��}��8�\0�:�充.]\p��$��~H�T���K���?ښ���;�.L���b�@pq����I��BG�\˯Y��Ƶ�?4�&�)����$����agc��Z�̓T�7Et\"HBa�I0O,p��.M����r;%c~[��~n�i'���K����T���K��V��7�ф�3��OAC1���I��i��?��_��쉉���O��ψ6}���H~�-�/Z���}�̨�{��>�#?�3Y2�Z�0��W�j����Xڣ�R,��=ї�?|�_������y�Lo�p!Ut�
G�E��%	u���\�Sc��k}2�1,��e)�u�U����,���?� ���%�.��L�Vu��S+r/��V��vPo��U��y�[<a��4����ZJ捲��]<|�4~��3쒇)eHiX���I �> �p�w�r!"�y�f2rv���8�qh}b�����6����K.�U�	��^$)�Yb-/fc���p#��j�f����t���oa���w��̳�Y ����C�(�2���x�a���K�coJ$������#��9�����O���7�+�=�Am6I�	�H�E(�$�q<��+٧1[*��.v�^>>.����G�6!�c��R��Eo9��r��)���5<��y�+�a�<���q�;c�H�����r��]Т��B
_�-�lj>��5U�����b�vXubjӣ���1f�ܖ�c�*�=M�j
�]ܽ��E�����.KR�`w1~�,
�u�+�C��Б�X�����)�f��c��#�+:I9=�4��e�s#����aIN�"7���R�n��t=j�f��N0��;~K`�l&�n/mF1t�ߗ��fD'��a	m��#�������J�b���p/��5&�2�Bm����h5��-|8
�ׄ������17- )qĂڝ�����N����bB�´�0f-�`a{����]�G
h�Ym�Cw�҃O8�z�po�ifi�>���=t��bJC�F�����o�eԒ��r���BSH K�wn7���`Δ�fztf����J*݃�.�bAp����\��V��#ra����@��/�E���#`�'꫗sw����͓*���꿎`N�����|j���m��΄AFM�s�x�4=τH��Z{5�f�^�ɶ6��y���??����r��j�q��� 1�?x%��5����Fxz���j9F���Z߻�#F~I�f9�[ 嗬������Ǻ5'aw���m9*��[8�.��В�*][*ڍ�
��