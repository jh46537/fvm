��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�a�[W;���(���=����n�|`&��'jJ)]E�:���}�M��ȹ�ۏ̙n�#^�u�y �g�D^��I�Xww��#�hq�㿕V�#�m��(?�H	*ҝ	=:�xݎ̇~��$�f~��?޺���T&#�s)ឱY�!:�{X�B���YD�}@���������N�ٌTt���yE��k*m"��z�z)�&Aj;��Y���=�āK�NXf^E�ȩY�ת[w�z�i��8[G-m���3.l��z�[M�V�3�_���e?������ԝwWB?p�A���%�֓�-��҂��nb"�Y[�a�-/E�tX��S�p2PO�����)#��T����!da.���3-��[#kU�2a�4��p=�5��bmX��mʪ�Up����\<#O
�^A�^>8@۝yʑ7��u4�7�[E�����2��0���NƁv~H��O�D8$.��k���"��1�8/pN�}��c2�K\^��R���Ѐʾ�:Z˽��z����R�E�]�V�@B@!z�Dt���D{0:�'a��.Ʒ|Y�e?�c��Ѧ**ܻ�RK������f�*����:{���5�u�W��f�[���(;�L��%��-Y�j,L��]7Ƭ�.�RC���a�^��C6�(�B"
z��� �P�w<'(2�P�x��2<;�5�}Z$����\��y�AQ�P��[���gtA���@��� �A�ۥ�)����w"��D��<�@�ye��G�N�����r�s^�sBt.�#.�_�v6��]Ĝӡ���SV��:~A�P�\�%�ǭ� ��S�K��z9�N.���\/*�H��W�H��1�%���C��!�4�b�d��LMn��Q�@�wU6'�T)��bWˇV���㠪Ӕ��b���DQ>����p���u QE�kӖ=OBLA^%�|�K{��� MAO����>D3�au?���y���
u��+�p��\���N
����NS�d����� �ѽ��1�Qy+sbK�F=D���F�#��v��i��p)��jt�l���zѕY� ��\�u��8Q�iͅD���q]�J�;�Њ��d�5����h{�U��?�j>C��^m����;׾�w�i�EUL����1i�	�������4辔�c�y��v��$rV�1�s ����3���㪂��ͽ2��;%��'���!æ
D��L�'����aa��a�������?� �B�JR*�n�i�?�G�	�u�^�\ �+<��/��oc��h�7�Ə=� ΢qeAO�A-`�,1��X4�K=��%/�K8�p�h���0���1�bC���Sa�����{ n��=)�2��A$�<���/ T���2��A�G��Dx�� W]7�t�:�N4!���.�D�#ADp�ྺ�,d�aT N`��~4h���M�'jkpY���`���Ɵ�>�����}U�`�F�;K��E��:	�6}��@�Z�b�Y�D"?�����I��ǒ��za���6�F��%`H�U�+F��k8�!nrL�k�I��HI��7���jz6��ͼ���Ϳ(2�qɸ�/���+CZ&M�$h����b�y�A���#Ń|H5~������=􄷀�� o)<O�p����m�����p����6"V󆀾ܩ����>	ˇs����#Ҿ�5��:r}Z@�z�f�_�=tI�ܧ}���f^@�Y���P�a��F��N�Ş#3/�<�:'�Rc��dͿ}a-���&W
�RAqS�_7��i����g�h�g�c�xk���"���kGfe����%��!�6e�\���i|zb܄���i�\�%�9�SI���2b3ZUMp�}���"A��������i}�J1e��ć#�����dC��r���S��I��5*-+rL��\Ŗ=���k�u�:"#wO�WO �/5?�>�����piE�}�vUNp�}ޔ*��	�
%��X��i2��8V��sy���pt��j�;C�~� ��+.� }�yʚ�Qx_5b�6o��X-�M���a6�/H���6�׶�ǃ�V'��1�5�ZQ���aצ��m�jgGݲ\�����������8�D�3}[:8�|��"��H ��-ME��b�b06h��8#KHEs��q>���i��h�~§pe� ؚk�1Ր
�'ȫ>��
�mz ��.]���%e�b�OX�u��'�Fd�w�f�̛�yR(E�T)�;x�����F[�|?�6��6`@e�c��
:&�#L�e1��	���R����BGr��� 5M#��Cg�Ǵ@��o6���}Xxx/c���{��0�`B8�yUv��M�@Cb����u@�o�݉���V�u��Z��^�}�W��l��n��A�)��څ
�[^@]�Ch�lES�G����֒7?Z&]i�JN���oW����n
�L�ӥ�?+�I l��x�Sџ��4�I�p�2��¹��-��:A@M�I=\�ϣ��&�ap��ǌ�"��-� ���m��y��=�����ঞH��[Y.r�"���Bd8�т�+�]�P ��@�A��x]\qV#lH�8NЂ��������i��W$����ɥ�ڨ�6�q~}z�m��@�Ji��8�i����%C��/6�����Q�u�p7�1#ڹ�����B\����.G!V8\�Ӫ��<��㪗�~+�y���ϛ�OO����hR�I���}H��.뭐�	|�V�=k����e����Q��pX��c�����l�	L��sC�c�j��m��hBTh<��(a9���0��3�F����zd���:�(�cu�� $��i�?�,G���p�al�L�[&,ϜU`O� ,��� �[^C
�n�a1E��q�W��kco���J�������H`�Rf:�W[�����G����a�=,�6�V�����:�N�;��+ҁ$W�?�`d����"=��d��HC̉U��F͙X�B��K�wn&�{"
4�j_�*��1K���U���g�T�ݦ&G�ʢu��C���;<��FF�G���b��J.�l��ME��LY�T���b(�����:�<�G'd�F�<���0�b��6�}�r�Z�5��>x��\㿇�cC[c����Aĸ��X��-6�F{R���m��G�'ʆ���A��9�������;?��-����s〛5���&�4r�L��Kִk:���̋�9�6�hP� �_r &����=�]�?;�*ڼ.�u�f:u��i���rI�d;`*�y}�v1��C�M����0h�F�o���E �� �Pp?{5+���)@�\TثH1���e��E�p_N��pQx|Y�J�ݯ�з��2۲��M�|x"w�߄���w�dz��0)"Z@��C�V1��ms4�`�|��e>�1�m� �L.\q�͸���On��ߋSr(:JJ5���>��~��/�U2���g�⌋�j�yV�Z�U��������b�[�b\�f7�p6�ۂ
��%]���ˊ�(�(ϮE�n,�I�s���P��<�1:�`Hb�\��{�,sr��:�����	)z����P���C,�o[��щgO�]V�&A��'�k�� �y��v~�I4�w����w�ďq�qs�%�u���UF�O3��g�9����5B�B��O_\�S�W��ZB��A��l���G؍���f�O��ꧩ�q�ۢ���W�ʘyG@W�Z^�&8%o���ښ������F0xQ�-��Zo�����b��H�79�5Y���N+h]�O���K��z��/t����D�=w��������B��8���8��5B�£�+mI��
E����m�!57�5������R"��1CCv�Wtw���oi�Z�7O�R/�T�]�����Q��dK:�Y}��H��bѺ9�@�~����r& ����A��.�����,jO�+2M��08���;*�_�J����8���#�A<m$=C�d�3/A{I}w�b�C�߾�'#8]b��-QbB`�h"Uhd�H+�沧'�h���{�L�	�J�ee��-d�x6�=`?����M�.����4ï�E��?��E��_�EM\�J�/��� ��5P��J��H�;����"�y1o�C��ѥJ+��2Z��`IY(�Fg1�����4��ª�z1��3r!����E��BN����Q���"�]?5�	�{Ea.�}g�(���W����\N_��
k��ה�G���^�Uu���KE���W�.p֋�jjͥ��#y�=��=y_Zr��)0(�Ŕq.�~p5!n�>��{�5���MʊW�����B��եu��3
�W��u'%��K�0�k��ϒؗEbUl�����.�x� Kb�vzE->	@\_�<mH=��j(���R|!^�G����rC2���[n��}������Z%��慆�A&p��D�pbP�f���*�WɄ�M;a�O��}��h�U㹨GjA%z}<W�t$G$)�e�C֊�H��w�f��Rw�X�g�eSti�a�썘=�ai���f�ɣ7I�y���V1���L-e�Q��ӵ��1S�b��&T��۲!x0�E{�s���<�x��pev'O/������IK&�p��Ց�41�5�v[�t��S����8�3��ߪ�GeF�u�=m���g�~��z�|pD(��G����&kʒ�U��]�]|���yq*��{|/�ʉ@L�`گM\���^1���k��C�H�k�Ǹ�چE}�*����&�<�9�y_Y^Id?�d�H�kݵ�q!���8(J���5f�a�R��˝��;|����3*�G��D��3��&=�C�"ϵm\eZg��ț%����A�'8��e���f=�ڸ�^i�����;�TQ��y����H�L�-x�,$%-Jl��J�a��Z0v{ /�Ym�W�~���Y���A���ε�Ao�7>�Az&���;˚��s���0�Ox׌:t=|�D<X-��:�I�;�_�.b��>s8Q���r,6��m��x+`_!�U���-���)�8���dӻ��L>�I��,R����#�5.��!�5g��KV���цL>�?�,�@gX$��8U��b�%�wg[v�����5�#;-��'׿��J�1[$��9�s��f�zO8r&ŕ�;/�/j�𘸵Xh�!�F�`�����BG4���z
�=����	�����]��gaK�sjE�^`�q-�U{�>�8�[	�v�)�i�Tg�Xκ�x:�"�e��������6�.r1B��.�r��Y�ɽ��j������$��i��Ղ:��d�*����-�3�N�Vs�<�l�C|QĨ����p�<��� �mz�p����	�?��1ڙ�������R�r_f�F0���E���O��V�'��q1@��$e�n���g�`�4��ޠ�4wV|O������ ��S�)q��Z�UL��,��7R�dR��@�d���u�PWu���L���o	�:;+�Fy��4�_�:��$�tzt$���G��3�)���[�����Af/�ם�a��6���Q����w��_�.nm[Vz�k�x^�������U�@�:_{4��*>t��ߚ
z5WD��5 ��!�$���4)R\����]9M.*�}b��Z^�Ε�%� Kf'��S>y�����\l���̀��w/�x��M�ӣY#30�,Giv(d'qLc��ny�Ц�_A�������N���5E�`{�w�q�P(�<W��	*���-���I�A�H��=ōV{9I`��ʍ[n������< �k�7;�v��Q=2�PheH���c�13 ̧59Z�P��{��=���	�������`��<}�MҦ[#Uu{����!u��v�"����ۡ~��{f���t �ZL[Nj���-��A���,[�5���_<4Np�U����~�e|���EB�������>}��W���1���X?N�a��ōsfF���VPt��mޛ��*C"у{��ɍ��;��E�(_�"I�UdY<�E������/���Y˲P�.�oʿ�O�zK�^��VffL�LϷ��8��\���ʕX0��@��f��6��e��QQL�c*�!����#��s�{��b/��5������3�X�c��O�T�.����F�I&lu�!�/�^]/Ŝ����j,����ثl���ûA����NI}oF�ƌ��>�@�,���@3bn�'�xf�*���+(ޙm5�y�G\��6�� (�˦JY!H.^U&b�K���r�L*�$�0֫ �'�=����u�W�A�ȵa�(b��z�)ߓ�b[q�z�C��,�q�����ʰ�X�vg��s�C0��ܸ�S�~K���«���1�����&�[��.�> '�1��C�ǩ��r�#��}�p-'��ȴ�?اVq�Ub���T$	�d��iZy� �B9L�H�����J�a j1�ɋhA7p��:Z���"�D��Z|��I��>��9�+r4w��wM>�Z2�7_e�LS���'�G���[E�O�i萕z�N�>��Aq;�a�i.dJֺ���ؔM�]i�X��J�t��n�2v	CN<�����C������#3J����ҹ�D�df��ɤ��Q��üh�4o��5���2�ꉳ�P�3��70s�)ep'����G	�G��\B �r�5��9$F#�`/�	�J��(��4oP�����}�2���˓�l�$�=��P�Jה@4��flԿ��P��*�.W�"��Z\>�_�f����z9��﬷����k��i��D�Hv�C�՗�O�!l(���-��q,⢦�}�^�mkX���l��8KW4|;Ɍ`s@�w�Y��*Jhg�kBN3�43X��sd�{
����"��)��-�c"���z/��Gݱ�ָ�����w���i5�Q���T�3�}�Ks�S��]t��y���A�7��U">�J����&Zn\�:e]	����4����>�xF-��M�}\�=��W�������1�q����)���(c	M��m_�R�r 8�3/���j.{`г+\J��B���&:P�k�"﹓�����f�]�\�+�����.�ա ��=<��_-�p�s_�:����ة8u�eS�R7o *NO>����p��F]7����4J4#h���X��9G���%t_�u����.�2[*�@�t7��\)���ٖ�4+kY�w�)XG�t�~�j7�I�I�H��y�tz��3<��Ha�<��"O��S���ۛE`�9�)�/.$sT�laC�-q��C��
S$���!�d
���{C�̇�r$~�,��k��!�ך�	*�:�L�&�q�k?���T��"�dW�b<+Q}�yJhr�e;�o2�aUMO�(��^�,�|�	��� �Ja-%�O!�K��b�����$�Ͽ��w�X*$��	��`	�N�_m`�y#���lF�|&�ff�Iu�<O�^}�V�P{w�4�r�z�:�X��P��͹Cidw����`��A>�<���e����+eT3{��s����fM�|�?ѿ��7� Ў"�y�߮?{����ʜ��Ћ�Q��
��{^��Nyr�����΅R����$�k���7#��&]��aB&��٫�k�rxG�J�D�l>=�2��Af���L�掋��������$m�g�\��>b�mc;�F��;�{���>s��J�l�u�\�^@�X�1��HO@��~.�b���i )����|�Q�L�����"(��gk���`��x"�y_�9G�^m��t�B���ChqtM�R�Ę�\~)��qV�?��꯼`�? <yV�/U6�Imqƴ0����_�av�0T���̿*/��|�<�e���(��i�*ZH�ʶ�ݴO���m���J�g8IH�>eX�#�B�|i4����b����n2j���dؚ�:��C�_��9�����%\G�i^�3�(wI~��_D�0&�Q�g��7f�'ɬ��)	ճy[z:}�ę�� ��H��X��6�9�)��t��Ie��ա%gmJ"' $c��4�J$V�K{��׭�x|�#P(���3C�]�3�|q��|���+��|�]>m�8�G��	�C"�^�v&.D�`�V|ٜx�Y+�B^Wo�f;P�x��\���nư��d|T��W��y�n�D��ݹj<�M�'�S������h�	Q�셾P9!�3�l����J����mqJP���:=�?���!�G,��R�g#*$sP�$��z�#t�����~��=�4�NU*��v=�,@��n��i��~a�������>�زikn�k�^%�t� ���� �p[<l��6v���j>��ٹ�h>��R$<��'ms�	���"��˂Ԧ+����m�ءf�MN�1�ՠ���o�3��AIFkbfXoD��00K�G(��lɊ��zK`\��	���p�}]~)i3(�������ħ�~�P�Y�d�ޙ�Ke"�
u0@��RY#r����sP$�m�+ ��l�r����}�3��Ų��K��܃1S�L�i�;A�Ļ��,�/��_^P���e�k�W���W�N��ڹ�=�q�QŦcL�8��/堈���"���o%a��p��&1!~)[��6�%_� �������0�G����S��8���:�T��9O���Wc��b2��8ᚐ+(3*�;cVMޯc��뒋�Ϳ�� 숛e����?@ٛjW��*0#�Y�:OS�A�΋LPB��cq'r������Z
H�8ut>�v�F���8���k9"۳�F�D�w�X��S��DJ�CZ�g�[L����Cx�(2R��1�������Z�z��� e�}���>�H��.��ϫΨY�"Nf$�LF�U#rU	w�O�Nb��Վ�u���J�fe����Q����8���ݣEW2ܷ���eɫȉ�T��"{��hʚ�$r��*<���B�{��]�VCH�%p�u
������/^mC�t�+���D�3�|�5�x���_��n m��6��<傷�n��t���?��_���]]Gr� ���u	G���������c�ۮ�'#Ȇ��X|��s�TP�G�p0Z�ThTR�7lP���غ�er�:��ѿ�C'0:�����O��׳$��o�䩗4r�A�|U�<^��������I��Y@�q�����W�˺%^�G�p�S�]���6A�PwE�E.�h���1VJ��$����PsҮ,B#���N6��jY�}�˧ʻ_��<ӿ������=_5#����OĞ�4�([Ov�c}�3*���Dʲ�9�DJ*��?TM1&�j*ӻ<���_8��
V��kF�P���bw��F��6"�T���!թ��56���.� ���
�ݐɅ?��(/[�3�Z��5�D3d���st>%������X���}��A���Jpg���G�[��� Xy�1����@Uh&�n�>Pz���` %�T�CL�5���m�^���]��!�������޿u@���ݕ����Ү���J�(l�ٞ��ng��	��UT���x�]����G����p-O8��,��F��"3K�?�ͷ�'���HM��� )��޵"L���տ�]a�(A�-a�M��!F��鸡]�UQ�<���YHiǔ�����w��`��yk5��r|�%�bJK��K���^�N�<Z������5N� S}[�����x�-"~�9���K�J�Ћua!����c���}��0�>i �ƀ����!�p�y�S'Ct�W�˯��Z�)��B/���o�0�*W�w�5+K��x�Ȥ�}s}���-�a��W��L8B2`w�1\��c����|��0�8iT���ޘ�X'z� ס3�'� �e��.��d�0=�U4#�(#zZm���Rh�r�2�Y��D���ݑi�K��3��a��E�-�[�QuXA@���m�&;��$��F�C�)���k�ܓڠ�B���7��ǔ��#���*��qo3l�b�ڻ��$�=y�Ĩ�?�������M_���3I��hI���D%J�p���<K�Éq���Rsqu��>o���]�:O��RV�t0�����C�K<�F�ADr����N��P��l�2�^��$\_�?ӷ���Rr������������:�P<��=�=k8w/�Ң�m�Y%|To�^U�P�@Z�_�����#�[:Y��Y�K>3�Ik�X`�E�n��ժ��Ir),r|�Ł�0�}&�)�*L���&k��,�{�eou�����!X�/Lf2�C�8&Kl��〉�Ě����^��\�`.Q8�ਁ 1$�UC�/��m'���c[9�w�$�z]O��%1�\�f��S���&f3&[u�:",S������LkF�zA��YO�p�
C�G���yt){��ȵ�w1���#gz@*1�M\�]x5	a��r�R=�����^AqI��*��lQ�݄H�j�4�.�>9������b��ʠw6쇟����:bY$o�T�oM"`���=W	ݘK��F�A��5E�
�[�"���f�3?P��r]�t��e8�sBg��pt�v\߂�Vz�4��B��􀥊s���h�p�^�yƼH�A�-P�iK�w�L��x��/O���82�QxCZ�3�/��c���㊔��b��1'�F~��	oЯ�J�j�	���G
�{1��kp�P�|r�~OJέ�bm�p�[m�XѴ���?�vA�1ބ��H��zw?���C�����C���POYO���Zk�� {�-����m?*��]���7ε�(^ԭ�I�����c�-�q��ZP7ѡ�@3~�Gy�^��_+�૑w�+/��a��W,��>6Yoe�=���k�"t�d='�.�/��o+����/��h�K���Sxxu�O���*Ey�?��A���ډv|i���Q�m��@we�Xq����m�Cr����$��������C����ٲ�9�D�K�,(���\S�+W)�N�����K���=F	-3���8�zy�u�P�W;DIXvS-,��Rjmk�*,!����4�,
��i�I�[�$)	Z>~?��h�6� �u W&�$�_���J�
Ӛ:p�Co��,yk2����"ń7�xu���M�'.���W(�9�}�͛'�Ԋ�N�8�n^5%ݻ�a�<���v�$:l�IE���-��D�p6�9��i�)Ua�)l@����Vz]%K�������X3�e�d�?96w���{��� ��e	����A�� �E�$m,RY�o�B�5��G�ֆ��g1ow���0LW�G�¥��ٟl�퓸8�;T�oi|�j��QA�*��}�8��	e�H��\5lӤ��Ѿ ��R����T���#�Vt�M�<����b�F>w�&s�A������ٳ	=�D&j��-������,�����Y�˱8�Q��UŁ�6=�~p�r�h�ͱh-�<���| ����>���U�?Z���tC6'�.�|'{p��<�x��Whm��|@������~������=�܄�1.ܡ?�Y�l�q��~<(]69uF^�|Rm߈��"l��DG=�V�m�f�C��=���/V�@O��#�s�f�E)���.�A�t��J�J���Z��>�nd)yY��΄�mA)8���0�����{��-g���D"�*^�5��M㬎����,�(�L����v�J��P�Q�k �dH�}��uEΘdFўs9{b.�Cµh���s����A����O�Ƒ��|)I���G~^gm�0�����@P�</���	�;���w��Cl���Ph��kU�3��ʏN�eӫ�K�G�GG�Q�b��)�?�{���q�sm3o~*7����2JҢ����O��I]ꢢ���*,">C{ ��F���و&ъ�]s9u��4�V��=.Ჷ'~~�������ͻY(��죠��s��W:e�[ό����Ҩ�VB׼u�C�2�N��L���T�B))���=v:�d��c��X��Kc0����&��՗�J)9����:҃0 ��~K4a�//U�C҃^�e�[M	N&���S�,������s*�1����u��%����t�P�:��C]���[?27�K:F�N��E3B����q���V�z�+&O@YD���Rj� *��Y�> �4�m���y�j�h䰭��g�Bxv�tf��y�.���cѼ�f5�ZQv���D�JZ�\Dڠ�D�ק�/���u����!:E2Bgym���n$�9f.=Agxj�)Zk��FJ;S,+�M�����B��d{��:նSW��Uʚ�Xᙍͮ�M��"~ R�6����_��Y�"=Y�WGF>��J

��hE��@H;�Nt��[.�a�"_!,؛V>S1Ot'֖@��Z���1v��O��U/hO��a7�ǬC�@x��	���JS��֊L�u�.�:�'�����4~ L������͝�@.���/�/a�j����A��ן�l�s�V
>{k�BlrII�x#�X�x���
�@U���O��r[0w0�z9�8��HhC]�Krtf��~Bѯe�0��a.,3���Mަ�����E�Ă'd뙙-c ɗ��o��M�Y(�^]Al�׋fZ�C�͟hH�߰����Q���� kI�Ä��(p��� �. �ɨ0��rp�V�k`�Q1�տ�*��f5%�t�Ы�t��w�_r�es���C��ݭ
�u�37W}�0�C���}�xl/
�t	�61Y��my~Dt��hF�ن���F߿�_�[":Ź�!��F�\�����v��!; N��g�^�0�6,`Gr���'B������-��*l.�Ώ�@j$�g�tڪ*	>m�f|n�?�'k�u���G;es�y�*��:P��eBa�F
˞�"N�{�W���*��Ⱐ�Ok	j�g���GZM/�vJ��#�Bȿ��(�:@�q��e&p�NB�Ǧ��y5����1i�p)�Cvh�Ƴ;t�q��CI���II]�TH�M؞F����s�Ge~G|ٿ���P�G㵖�q�pX��($}�=��4��8�Q���I3ƙ�}�iDG���	��""F�V"6���d�EW��n���s�� 0<�﷟
O���(��n��V��{1��X�Ǯ�?�F��59T,��Ob�s��O/��X��=��X�X��w��l�_%
�~�]J��f���ԅ�����5]$�}*=��qR�
樜����C�'��ŉfN�Clg#P�&�6�t�7��0_�{Fm��g�a\�*Ui\ӔGB��G�HԄPNT��Ĺٸ�A�=�Q�`,�vճTr��\d��)\����Ν�e�����ٰʖc�\��{�s��E���ˮ����TrUh�A`�d+ˀ Z�w�H$�k�"�X����x2 F+�I�KJ�Ҫ�[y�c`L9����h��6��;�ٖ�����+%P~Q�OZ�c�_߶��Á���t��<%Sd�fJK�ҠF=n�+H�*�d�T{n�_�����ƃ/&��A��.f�V��Z��	��|�� ����Fjs���iF(���	�rU���}���h����XU�����dA�@=�T ;��Z.X��HMHP�<�>��p/�Pr4�?<}����Z��z�S���R����`����5�������V�p�����0�%�h�)��I0+�b�t=L�(�Y(N���ELn���т���k�`���r)�;k�<�./��#�)��# �nH�5�H�*�m���]*	��4��b�v�p,Q�����ǔJ�-JxY�(e���EFp���o3p��=��w����#}	�9�\��;������2\�9S*0GsA�*J��FȌ��;
��U[To��[u"��Z�wJ��ш�l~Z�g�� !�&��)���E���<Up$n3R
�N���ϖ�%<= w~a��jA?���3S-ЮuESʽc��?w�v xƀe��q���SDǌl�@�k�gYfTJ�<A�,�v��K2�B�^����R#�G	�Ao�l�v2��ce=��K!�k�8�>5��s$0}1��ᩗ�-��.\�=�"&��$Gu��L<R5S`�{u�烃g�˯ΈK��w����}��E�?k^���(�hۍSZ�<��?��&{9�Q��:�4�]���	4����8%����o6�bH4�ǽ������=D�?*�y޻9���*���@m���)W=��я�4�2oC���et���r�$ގz�ʾa���Z0��obt,i晝I%B�+�9w��j��In��	����������W��(]�g�E~�*"0�a^�P��I'~"�r����81e_I`+��Kg4׫��#y�U'q�O�yT ����>o�QѴã��\CQ�[�-<H���;:./1��W��(gh |�^�x�"�1C��[2�q{�:"Ab)��(�= [i��2�&�
I���h��'-��,0a�E3u�����ڊX�eH+�5�hVI��}���Q�Hg+�vLJ�������eC���jF�l|s�f.Z�e=��E67R����U��5�&N�g���1Rk%��Y���C�?��~�����F���v�"�X�[
a�ț��,1W=�f�S�aRU;ttj�<�h"��bg%y������������me�dr���?xd�V��{��9�i�ݕ�X�6ID&��������W�<:n�;B@�v3ˬƎ�3�X��㝌2�Wt"Aliշ^���!��ʽ����Xr�1C��2
�W�:?�$����kq�zG}�[��׳��S��]�����U��[`�y�n�<�,=���"Rw���{�L0���C�J`R�2���#����]HPT�i�X5�?C?a#1�&a���+C_���_OWKB�.NM?*�����%��XNz��J��^��L�;�����Tp�����;��՘a�N@E�������,�l%�mJ�������dm�:��o��X�C�^�[L�g]��	v�K�&e�/�6�����:G�Ń�D<�H_�Kܶ��� ��%O�2d��껎 ��:�4 a󘆴d-��"R�HkXH�6�@��������7�=���M7�����i]ޮe�o�te�ސ�<�jw���
&�"�y�5V"�++��?�T�౬κj@��v4"�b;��7ˤ�+g�z]lz�50:�e2ꠑ���T��[ �N���žQu�|,ֶ�����`70�9d���&d�;.5�W��-.�v{�vLt�zj� �P�;G���A�j���U��Jew���3�0�y�QM�PUO����%��p�2��/���蟮�Y��Iי�YJ<��U�洓��z�v��i��!mߔq���*!��u���Ed�N@������o^�}:\���0�joy�d{J�.(�O�~�l�i��T�y{+U�=-��|�$��u�� �N!�����_�(�������A{�ˉe��y��(s�hq���e�&#�^/�a�����T�0XF���)�t&���)[���C\�/U���qy6��4�-�T�a�4��0���vh�P�Љ0���O!S� ��V�%âxϫ���]�=�x���	MAٶN�=���g�7B�.a�m�gs8��E<'N�D兢+M�淾��Y��5Nd��FF��~!�տJ*��AS�3�ͪ?�����S�aC'_ݙ�(K�q�WӾ)�9��-��2��gK���ﲃ���f�N���Zͅ	R����*f�v0Ö\��$)B��{f��`��1e��
;[{�Y����g7�����c��8I6(H"���r�:�؇����y|����榶�j�f�o#"3�ت���������X��)o(��m��0��W.��ďϡ�f��Kd{=;.�2��bO��	gc��GS�+%7Ҭ�s{�u�q�0��]���a�nZ���O�Z�ȹ�ѯ
z@{�J}�����3�j�l�gb�rC<i��;�!��B��	D������R��$ 
EڞNf�]1�j=���x����Dl$x���XI��������?�e6i���"���w����3�о�x@@N�I� �|:o
�t�t���/�� ��E)2�h%������~l5��9�!2��Y'������7R��!�l�R<�j�O>a8�+�RW���Mשq��&�=t=���۰�;�ӯ@�\���]S<_�^7X	ʱ�[�.�R��B���+N�����gEfԱ:Ez��.(��P�r��Q�x�}f���Źq�'��0;h�� ���=ո�*��v�����bR��������̧�qh�ն��64ܼ�O��/e\"�%����o�5;��%fO��0	Mt1���aY[SW�m��x�~S[��L���sJf�D�^���n�L���mk:�y�J1����5&lժ�(�Z��|��f�n�o.O�"ܚ�um둸��`���F�g�y����ꆾ)4�J�jɪ3yU-�n�o��� �C����!4KI6�=Pdv��_1�&�>&�?ם���K�W*/*��{�G�#�X���&"X*@�R	#��9yr��q6��r]]/J6l#��(�ީ�<�X��hv�>��u��p'���6G��X��3�
�	�T���� �E�#X�͎�C|�0\m�S����'��_Mb���r�OL�H�nK�b�n`B֯M�e1 � zP�$̥�������#���v�̽���
����Fv�\\!r!~x�CV��ǩ�Ϸ�9����H�g_���9�pC��Ļ�K�?��Ge���f�P��ZS�*���C��?Y>\M����X��X����@z�˩g���=����v*�]M���@.�A�C��茀��F`=l���jr쒒d�cn�'9cԣ��$�9p��Y-��ӓ�M�-�>a�@G�����m�a�s��CR���f&|����/ɣ��.��'�� [ݠ�ۑ�/��l���4��C�����[!w7I/s��e��	����÷�ԓ�� ;�/iLn�D,@%�]�4o�І�11��r[[3l����̵Z=14���R ��BU��hZ�4?�u��h�'ת�A �ٳ��:N��/�j\�(C;n�^��KΛ���yO-�x��_u+��B�QZb�)~���k0y��?H�'<E�Pd��-�{;:��a�5F5Zį�3J����MBw�32ZZ<v���ĽXbQ��_�Ae�ixJ��8څ'f2-�+�)Js�k#x��l*	�.�cD��F��ݞ I��Wx6j+3���*�ǅ?{��CiSe�٠p.�q�nߴQS�%8�*��i�9[��j$FR8�ð�[]>IK�wu>]�'�d��&a��,�}0!2�d~9����)i���B��<5�~��+�~E� ����f�U�'m��]�^2�:�ݡt��>% �X����=�|���~�#O��v���پ[�Q���'�F�tp7�	|g'��3��S�a��_��6�><���e���AP�/�. ���TJT����
�^.*5}������P���M�Ѵ�atI�ԟ�\҃���5���Jh�xU��S7�$��xD���R�+j�4�I���dRE޸[� A24�d:M-rzq>�v�q��N2�*����bR7�������֦�������z���G`�������ϽJ�4�������n�/���b}X�Yg����('�M�B<_�'r�v�r��W���A�B%&rO���̧���A�K�2g?78?̼@��� �f��,[|��O
u=K{BwD�s�+��>e���.���$8�XfC)�O*�_��M���|P�esڬRv<�d1�P�tzl+}�-�h��9��0�K��"�`�S�#�� ����̧��KS��̫�8|`�v�6��\R�l���b�^�]����H�C,�+��!vVs�d��%/�~-Ь]�S�۽�{ofXф�"��G��rR�~Y��j�����_{���C�/�I:(nX󼄲��%�c��ߔ�}U �;\\���W¸א������	l��L�q��?
C�����":������Q`\�Ť�JA���@ֈ��2!�Ā���{�-4��q�u�vɎl�e��[����̀�h+��ح,ʋ�a��;̰�E��������u
>3a8Q¦y
3�a�o��;��M��aDa�p]F��l�0��(hi�~�2�)5>&jV�s�"���Rk�s��V�܄\{���q���1�4	�-H�]����1K�鸡�[���֥I����@K??.v�H�H�mV��z���֤'nfU��s��t�S�h'{!�V&����1VM�9�a�z�T�q���0�f[�����ѽ��	S\Uc�id�nD<J���~�7ǘkz�H�= ,���7D%*Ro��רּ�6e��s� p��R
tz!+/	W��L2��j�5���3��)% E��f��q����