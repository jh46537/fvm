��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^S��A}�N��G�޺��Mj�;c��� ���^�4�p����#v(�z�7�b��=��ŝ�C�G������Z��I�����!:�{��[Dx��a��2s��푳B�`�~���W�������C�&� ��u`_�+���!���G�t�c͟�3�J�WoQ��(��A?�E�B5bX�"F�y}�c���#���4m"	6�9�T>���6��4Ume��H�����6c�􏂶]�<�=���*�~�*���%���8����C-�d�^W�BW�}>E�w�3.c��$�<���u��j�h�r��1	6�C��ӖV��">r��, �ڑ�vv��I3�EHG�q�R�;K�������,�D
\���~�@ΆR���
��S	��e2Oյ\�D��봮%�N	��N��r�b����n������P���
�������W�ǜ�Z��D���
Z�b@o^��R� �-��OI$�Mؾ>��χd��U7r�cו�w����'��P�~�p�@#�u)<�\�p{�����q�J���$��"��T|ʽ�^�s]��z�ν�Ǆ����^oé��ʃ3ï{�0�JIݻ?�
e6��n*�)��Ohio�Nk��a�-!ƕ[�X|�. GZa&��d6���G����@7��p�~P�S�~nne��<�f��7q$���,&{���j�T����j���^�V�u�SԦ�9_�� t:4���4�sÍ�L�G�1��\���s��F�ɸL�}�<���u�8���@@;�Y��6<(p�'�7�iN��B}�e27����3�P򔒜��q|@� �{�x	�X7�w]" �0�̽W�����
(2���.��H��I���J$_Mǁ>&�����IZ�T���3���I�R����j�0'�o�F���L���C�w�/�����4p��I[�Xݍ8����n3����g>kKuy�w�a��/k��ܠ��!'�ݯ�+��������?U`�9�D��]kt��g#��}�q\+�j�,�J�{u�Z�Hנ���S�	�;`�-7�Q��$Ὃ@؍�WZ��BM���W!�+��d.]b��gBѩ�;�Ru�(~�B�O�&�5-�]	�V�
 ��B�UyT��I���E�i[w�6����C�k�mB�u���~7�V�Z@-W��wP���fq�pn�%� �b�@�k�4�o"��z}g/��j��b8L�f��%15٬Dh N���[\A�D� �UR�u�K�V@6�R������AʷV���"Җ��'FfŃc�5Ĵ��=66�5�P��p$٤N����qMJdNb]NqM�/���_�[��&1kd��d~5�`0�K��{���o����5�ԫ1�K�	e���WT47����x�=ݭ���I�ɥ�+�Cg�C<���}��T�N�w��,�vQcl�>z}`ό>��1ȱǌV+INSA��LŚ��:��f�$���w���!�+Z����:��ns¼�9��x�Я��U~& �{��r`stg��=t���L���|w������O�o��W�̈�#aa[��_'o�X���c���Ư�3u���/��M��^�|��;puv�Qs��j��%�vbH��,�Xv����53�$��[���Y˙��=IL�Q���h�����Ȟop�Q�d|f��ܵ��p�l2��cX�u�>\�T8�O��Q��l�51qU��82���=�������Xk���f.����_�:�85�I�2������Jsc�͘A�z�\@�A`��!X_�U{*����X)�9�33��ա�I�I�'����*���M~��	v9`B"����@oTT�Eo���	br����UZ�����Zu8*�b��]��%�<���;�کB�h�Cx�Q��o`	�\�q�ń�އ% ��F��Vl%�
�v�lbvj�] �eU���Y���0ϣu�Yq\~��ϛ��C�7O�l�-�bg�Q�x8�S�&q8PuS�Z`B��vG��KKwl�IO��&�&Ճ��
_�"���:C�XV^�d"!�"�u޳��$������_(�u�#	�{�� /f,�q�[V-Z+��œS��0�P����^/:{�-�'�7����;�e���Dl�=3/���^����=Z[}^�	z���I���@9ĵc��g8���[V�@[q��G�6��)[��!EBD>^���=/���R��CbQ�F���9��ÏP�xd�W���^Z����ߝ�T���<|��_:�iQC�%>�&#�M�J����2}���]�6ğ����d����"#v=��ߔ�XB�'+���)"q�6�|�Dr$��_D'����B��x|�5m֘�1=v��cm&�?�ǲH+�Z�}� ��ɵϱb�*H�U�g���JǍ?\��]�����C�/n�ꌎ�7Z����ו�5�H�� *��?�R���0k]��'���)�6�g���@R%����*���W��p����*���8������+�PR^C���j�9�����1 aO����Dd���L��DX�=SDM��E�VˀD�H#'�̞ɲ`�i}7�����=f%�Q�P����������b���rl��� jA�A�Q!熯�:�(�\ �AA�����Ƚɪh�\��{>�)� �a0a�f�@�/�e��H
�G׊3�{��2����pw0Iܫ�΃����r�b�1X�@���$�"Ya�5�)a���R�B�"�S@ƽ�O�P]�b7�����e�g��([���A�H�*w`U z���4*�*��8�%�Yd�,�Z�R,�*�����Am&�f���rd2|�9�bz� ���|u���jl�L]��Q�ݹ%�CN^�k%:�+�Z�.����O�V����]�ęl`[e�ʭ2���¯Z�M*��/�]�u��i�d���i�*�O���">d�N@�j-�l4s�M��U��Gu�k��gcu�ǱS��@���ӟX��1��0g<q�?ӯ�����6���ǅqg��+a-5�l�j3��@�z���ca+��΁}����� �Ueܳ9��O��Y[��V�ߡ�My�I(������O*�/�^�W��>�����3Z�%��rF$�%V��ԡ���$�%��y�I���zŉ_����=+����'� ɟH7�����͘���ʧj�l����OZqPo^*db��+ѳ�_�Pb�uf�A���#v*��)�]�u�I����4��Qʽc�fn<~H�^��� hQg:Xz�)���汧&��}�j8�|��2���ϣv�v�0<�B���p��0;}V�IE$ǡ X{:�Nc�Hs�H9'>"�Y���0 ~oc�����La�BX�'&X�q��@2���X�TThs��]�f�M���G]x�̏ `cإ�өw�e=e����ɚ����� ����ҿ�d��DG>㿨�	:���<��Ny���	�1Akw���nVBr��x�r�D��e���T��lm��b�sm�_��t��_F1����v!����˥�4.������d0���G
=#q�j�BR�����>?`pp�	t�{�D�??+�����lm��R�pv��r��MV�'7��%�tװǫ����^eg^�p��3� j%z���}y�����X�oԗ�vax�+JؾЯlt�A~Z�.�y����v1z���'���	e�x�ܥn�hڀ��@��Kt�*F�y��9t/Q4ϴ��w�x9�FS9��˱�֋r�[O>]�\-�no�܈^��z��g���0�ҡYa��:��5�"Q�Rk~�Ur��b2��Ɠ�n_V�d�/C��Ym7�2%��f$U����qrf���m�o�l�y*x!V��P�Q�*Ƣ0贽Dp�&�4i�]`���ge?H�<�*����5�������Ɩ��\hZ������SNY!����  � ��a(!�n����4�_>H�� m+�]�S���(�YJ��$`��5 ��Ԅֶ�h�ާ��R9�b�2]������JT�̒O��<C-���B�a�8�|��K
&�7g�
7������lJ{=�����"��hw紩 �]�^�Ȣ 
^� �j^�eaq�|�:{��gR�Ϣ�y
� Q~@�_�x6��tл��@��Z���t�:�.Qe$4]D�d���t���fy��³�b��@g��������:�� ��ޝ�
"���4��_�"���nX��|Y>ܭY��R.��{гy���T�A���=�α� ��_6h�X�_��l%^��d!��-{�����Y��QB��{f=m�6 �����c�����N���۞I�e�s%���>�r��+��:pYϨަ�>E�Mxэ@�� �4��	l��S$�C���s�;Y|´0P�s-����H�|������LiA�s٠;Sw��!���n�R�5�?Xi��X�rW�ܜ�f8����JR58K�S�N�K�MIt4�|=Q�R}����}��C��y̤qU�m�K������b�X�6�͝cE���
�i�)������Z��]y��T��yo����,t�7^�]����]؉���K�QRt4��؋�a�)��E`�^s�o�;���gŏVh��v8��u�.�;dv\���I���U���m�D�PQHP���h3��ns5�O�dD����\�e��"�и&�/-!2�=;���F�uD�����U�-S�Itg-�P��4�VN��q�5F�է�� (
����b��,��6��5����K��T��w��ŴΛ�y��j�E{�Q�.J�@�dNQ���ݎZ2�+e45Vn�l��d|+�-�N1�H�]lP��=�_�y�DNY&j�)�H�K�$r��0c��Z<Q��{��$'�B@V�t0�h7=�i�-���*f���B���7JE$ 0(s��y$�R�?XcJ�s'`4����g�,ӫ�伞�g���J*gG�܃�	6�,��-i��Zm���롪
��SY�ބ%2Y7!��f�&ɂ��ҿZ�s���o���PT}�K��Ch0����j��C�QΆƅ�fM�I�&d
��;�3uq������Y���o��pq�P��ͬ3�x�4E4VJ��&�_��L�c�m�����1�6Њ����Q&�x�u�՛���H�:�C�'�j�@�l�X�E�-'�lӋ�X�^���?�5�<���R<7:�x ��_H
��ߠ%Vc�)�\a.�� ��鼱s�p����~���[S��?�R� �����5��c��q�	uԍ�q W���F���T���!���͑�J{���E��[�yH%w�UF2���M:��Ӣ؇@�:EI������r��	a��铈��]�Ax�䉕.�A��%���פ��1��Zp��\����p.'�qF�.e�RVw��`�C(��Klu�*6�K�z0�����#���J�X�����.�}����"p�X|s%��품�U8
+�>¬{�N�$Ձ�^U*d�u~��"+L#Bj���Q�y��J�#��j���t�f$#�#������G��	h�Sf0>����Zv�����F�=���n���!By2�䙅�=��0�m��\nA�fŤw@��s�mp�������ҙ�M(�d��L�(�'/�e$b
��jʶ��{Xȵ�SE%Ԅ����tC���b&U>�����������M:b��A��K�3�9�@*򷽛�u�eȋ#����1��y
����8�`���������H�<|3�]!�;���>�y$�J��є��cX/���j����,��^B��C�V�!J��<�(]�g
�l@�Qh8y�'�I�%�O��g";9����}'�v�h<}/Œ���)�ӳ�
��Ŗ:4��6εf�Y��,�`9Wd�	�����\G���	J�M�FAޣ�w���� ���py��Ŋ���]�e����v���S�P��K�s��a�:~�$��dJ�}�$��(���j^�8_Q�nm�:�H��Kd�zX"�X��7M&#���C�k��R,��s���(ozMOZ�ŊK6N|����v�/r"����ًf�)A�������/����ͦ[B �u�dYYL����QlH