��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0��؄i���^�{���b�e��_�@�*��Ht�'��p�z`��A�s\ꗪ���}�SAu7 ����G)ž�,zJ��S��H'燵��� �K�����I�ze#wH��1���nF^.݊4T�+�J�ֲ�i�V�, ��B�������&�)���� �$��E��i{��Hܦ���ٔsrgAM�c���=
�i�����<�ix�8/Ƅ���rWo
6m��h����b
�wx�^~�t7��>�52Z�QI��NmuG��@�!�C'�h\�e�C�Z)9��
�v��YP�椻ޓΫ���	����NloeJT�C`�",	��~���m�l<���y����c/X��S�h�'�f�rv	Q�爳���w�k��*���C����H ��5 ��$�۹�����ۻ���O��SF#l�KI� r�(,���T�,�o�Xn��]��?���Ĩo��ٳ`�u� 楯#r̎����H�z����2�)��TT��aJ]�<�� s�:����
�8�.�[�;� �0�w�ޭ��f�Fx�����4�F�Q�T ��b� ��43���`�\Ҿ߯#]}���(WaU���,�$���@_��w`z��yq�c�
��Ȍ<v��^�i�;�+��:��Tӂ�Q8
���`1�喍�ܿ��ޟ�u��wm��3�f�k�x�y�PT�����t/���fC3&4>凌0Ւ��2Ь��i��u�.6�k��D���\�pWV�P������A���-���#��7�%���A���7�U�ɥ\\�m�:��D:�6v��Q���^���KJT,��ͭ��`��v:��}^¦k5�Ci0!!��=5�okQ���|`�������!�a$?_���#��a��u�)7�w�hs�W��*��]��j
H� ���M��[�Z}9̄(Ð.����@����%#�V�b�����d(��F?{���p������㨈e	�����F��*j��Ь�`�nә98���4ӓ�[��'uU2��χ7�A��Z��-'���'D��O_��o��)2Z�·�#c��;5q���������2?, ��Q֮_����M'v���gd�r���|�FR�+�U���y���c}��;�3"��y����~9�/;k$��!�,����� ��l����Q��Ms���ޕɴ+ۆݫ\Hhy�%���RJN���y%�:�ܙ.�]M\����mL��:P��6�x���!�G#q�O���?Ք)[�J��Y��ܮ��QϮ@㟛�g���A��*|}OVRc(=����dHjo.�>��0/���ÿ���/�e�(풙T/��إujt&^��]<4D,�##�/R�m�Y����&}�ł���'�ύ��k5R���د��܋�V��@Dmi���܍��vJ���Pa�1c�%�o�n�RmRw�X��`yuU8�R������S��
����{l-;��
��-���854 ����io2���?±nt��O�kK�d�Sxm^��9>/�8���Rd���C��c����88�0�ZǷ������O���v�y�OZI��������T:��/!|�CE�/�Bȧ���YkW�=��H��٬��X��<�T@��u�sz�q�>VǞ�����A?e����g�2��j���/��-���{:t}	X*�+�<\�kB���v8<���)#p��`>GW����7���&<[��4�8'UI��o�x�RI���/d]�i�
�y���z+�I܁}T�f���/Y1ʲ?$��[;NwHc#?:�}g�鐚J���Y���j�Ӓ����u#��uYb �=2uM��n�^�=����%�������>H���8�����D��KU9�Șٓa�n�1�c�(�x�V��2A���H
h:�;�g�QҤ�eka��������\�+ˍ�Z!ͥD|,'�s-���57+b�`U(bu��	'@^]u�jx>���0��Rw��\b�A%^e���_�1���Rه���ZЩg_�\�ɯ����QB���tL���L�� 1�[� ��[!v8���}�2��R�-����\���]7B�w�O�}�h0D�/�ZU�A�K|���2�a�F��8'�ׂ�Z�G�Mp�J�1��$Z+��aei �&	S������ABQ�ffy3������� ������,	��J�"%e��JV���M!��-�q��eI���0���?$εl�uX����`�X0����\i��+��Y�p�9-Ba���Z�=�#�<-��7�]�F�J���M� m��ȇ�[��or6��{3�I@=�zw�'��>ϢV��'.^�T�0��}�IpI�,���$J4R;wQ�,U��?����D��c��{��1����O�UV�mˣ��m2�,��2�n�Fq�a��i�w[�pw�\Q':$�J��*�Ow]���s���V���e	�ڎ�]�q�vZ���:x�<&�8����*+:?:;O�ȻZ��S��,M���QZ� �<;���=8M�8�
G�W^[F(�垝�&Dd�Q.՜Z��Gl���O�)q���i��#�+�� ��C���e*k�<���M?�-HۗW�~��y��� .6"�y�]"Ǟ&��^l�X�2��
��h�2S�j�-jp��&z�IUb=�A�5ˀ=[�_mo��Jn�;S�d�u�5��ej�7�֒� ��c�aE�����|�z�[`V�<!��-5��ds� ��N�GN��E�d��#"���7��Ԉ��ޮ�������p�FD]ب���%��*D}�ߗ��܊���?������ �><�p�6�_�i�'ѷ�w͒��{?4;�m/�qS�Z��*��=!S9�����t
�y�5a�����A}!!'������gR+4l����13�Yy���Yh" 6��ڂϿ\��<�NӪ�^�Me�M��']�To����I�vT��q�8Ƞ�+j+����ÿv�J�S�l������L�02 �Rb�Fʵ �7�t�>�A�Oޥۋ���xW�h�z�R5A?cRP���}�2�u ���7X_��;��b�yGF ���'ŨSj�Κ%�N��1�^���eаr����o->>��q��cR/X�>��2�7γ���0zإq������)B<d@�����t̓�����uA��z��wBE����2�E���E���E�Ϩ�#�����K�ܙX��Ц�:�9_���E���N�k��P��<�o��%���?��Hy.��ɝ<�4R�I�0��-<�n�.�0�la�x�\Gi"S!Xy�/ �����;�:��"�E��0��d��n�}�/�o���!@B!��aJ�P��̒/}���ck�