��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzk��f�-�ך?׌�1� ��n����4��z�����%}=�k�g�+'4h'~k�W%�x��<�,:0%Z*~�%T��8����LJy�oW��V��q�lj�eG=�s�#ø��A��3�C�t.�K�Y#nHX�Dֲ�q���i��>Vb��ฝUY�
-u��d̯ẓ���S���CbF2.A4҈[B��)uYz̎�z�
k����ǡ���N�����z��#����m$��7�RҲ[�\�*��͂��]��4P�������8"��Ҝ4;���y��dW?��ښ��E	�k}�GAO��%�1*�y�~T���x��w���3��epm������(�^(�R������B��(߀l����P�1uPD2��	F.B:;'���-s���F����� �X?\�1!V�Y ��Q���D��0uN>b�;2�C'���:����X�����
֦7f�19'��ɎEt�w�����������Y�����~\^B��m�E���cTɞ�����+��Q�[��fsE��v�� �ʑ)yHJU'�>c:l:��B4�&��"���	��uߧ$:^B�xc�?��<2��/���vp"�b2d(��E�F��Cnp��1{�w���}�u����۾�r#��� !���q��l�/G� d�+,{t;�J�X�v.��MX�5�R�B#�;��
�q�[��/M�}8��Cb��9@�T$���F�|�X��&h��!���b�e��z����5[̬�R��Kd�l�w�۾����8��X�����<�g�E'/ێgxX�KI�n3����⺁����]��5��[�K�f������P�0
���lEJ���轀�:��-�
�?�P�C�16��q���+d�`�!K����݂�ޘ�(m��Fi�븴���i�Q�����oFV(�,�qZT~o <�9�׹`J�u�?&��(�_��[ь\�)J�z����j
8`�k=��xN�˴1{y�qaAP	]c�t�E���p��K8���9V;H/�O~ ،�w������@y�^��o+Q@`������ƃA0�|�� ��L���"Qw z��{3�H��{�w��cd[��H��/�l987z4j҄�Y�c7�kb��p&�� �j~��h�x4J��F�����V⚭��ϣ5�Ƿ�&���T��B��LJ��]]${ښ��~ć��D�<��6=ˌ���v"����Iq��*ϕ����2M�nK�$AWm�Ar�U��q8��j�n���:/����%H��e�@a�CPM:�|��P&�����h�9d	^��� ��q����9+������'&��x�.*7��?+�`^��hv�X����ى�#!!��(ӄ96�jp���
�rWnX�1��Z)�8��b;:�oN�?�~��f�����W�ߜH���Sq�+�u�V�,.\/�a5��	9�:5�|2��&ok��`�:߼l�&�	� <�;]ϳ�ZG2�^a�H��U��B��/��� �:߮6s��j�wr��;7Rzp`ar"��4�b�a�8>艪a&��Â)�����R��I}�^t���x8�T��e��)2y9=?(�纀@���֮�h`)u������ҝ�r�	ӄCOٰ�����8{e%����*l�>n�ilvՓ����Կ�+��5�h��d�T�y6#�>s������׀�@���U\4�~�Y�t���O3Q��i]|����$��nm��_4i��՛Ȱޣ�?`�C�9ޖ~��(8�h2���e�\rj��O�qz*�Y�g����K;���E���{Kb@s{A�̀k`���:��l2�1���_� �F�O����Y
:v�����n���/����e�5�Ib�m
��3۫�>��(��Y^�/!,�ǖҲ��X[%p[Y|-�i3Z�or6}׫�_�Σ�Z��sA+��p�I6��� ��ԇ��J��-��5"W�������*�5��e'A&�Ee�(4]�glUV@�F��������LH��T�4X��L��^�9�j�������	dU�E��0o�?�ڃI�2/��]��8pyN�k1Csgu(����!�据�Ӊ�Fp�� l՚���-8]�#��^����}��U��ƕŶ	x���-UU&C�l
�`�K�c�Q����7��r�X��N��U��Db����%\w`����� I+@X$�W��J��,Q2kI�u�M*`���^�9@rw�5�,��3�R���څ�ڋ3g�>3�̵����0_�[����Ih�������~��`=XR���&&u����3����p�T�hR[�
����F#�,E��C�`�j��9SP�72���9y��<'О���3��K�V��mp>Z����dw~u5�h����������Q�S�y+��W��	���}��-��1h��쿾�H8ב��_}�(�5�p�I8p��~xm����	��[�{~�튻�p���'L���l�{�v�u�D�.M~��В�p�*p_�/���f���=��럘��D����8\�g���Y,��Aj����B�˦�	��an�k��^XVsGh�]?u�<r�����K]�Xw[q�2�ٗl��lO�H$w�������_O��H�z�M�?B���'�i�ye���}o/����M1 .�u�x��[e3w�r��4�ې��2@ k�C<�/�\���1�\�aF��i~Χ�Ʒ�I�8E���6��3*�6���g�P~��E�R��c�k��|��@�������2M�Ij���".:�5�ܟ����T��WI����\%�a񨾥�>A��)K{ъ^�c���3�S`��S^l6g�⍧��-7*��<�*.��׷ol�۹�#�,�wA�	?��|�n��x�0l�A�Z����K�_��KAu�7�p��A�����Z�(�Ï�����H�l���)/��DQ��Ǹ���R���y�/{�!�Eh��sZzT�����Q��b���?�U8�݂���XK�aR�1!0B�P��HX�Qs偯���:���g���Dh�	�``��QD��~�3Tz�qF��ZT7Uy����"�'�0>�ݾM�x��F3�R���SԴ��|-inA`�p�H˾�a��ӻ�����$a�I<Ð"�y+ut��Oz�
^ў���yIV���	��cp�:�H���IMns���ߘ�^QJ���݁�Gc���b#	�J������0��|ɻU>R׀4]���nȞ1'{r��8�1U!�wn`~�Qi�QG��~�l�4H3rp�uo�Rқ�����~%�g����`���	����C�X�7�!�0��-�:Y�ʽ��jMS�B��ݖ.�����`�n�����d@4g�N@����V�6vsR�� "I9�$n���#0�4���3x����+���yG�^yXyAz4u#9�!1Dͷ�׵k��n������($�a�!����G9�y�v^�Z��sX���GNL� ��d�-�д�"L*܇��&�7��+�Z���NXWa��b	�q�'�p��Dw��"�nxa�v�t=w��_V‣�>ƣ�B)��F6C�9�T�V6��u����Vk�ok�)ϞJ��A� �Cy��W>��p�Y�cK��!h����[7��t��~k��傧;m�,Z��f/;�s�.2��j%j�F6#�.z�2ɬ�B�MP���.�71O��K�h�qa ���$�ʷ%�}/�CF��׾��qP��ٲ��ȱP�U/�8�� �ѡb����A���W	BQ/��-l�"���/l��}/W�RV��k3��,>�)E���L�6�d@T�ȧ�ʄ��8߲�PЄRsd"feI,������jtg�(��j˪�9����3ӡ	q�HH�O,f�bf�C�_�TWo�J�܉]�/�&kS�T�J&�T�H}{1�����I"��<��mb��ߌ{�@qq2Mh?yDҁl�~��[�E�XX�>_��$��rL炙o�Ф)�P��H�JJR]�m8��E�͕K��l�'d����&|t3��}�6?���%�Jx	LbR�yQ���O�������[�m	3����3v[�_� Ng����J޿�|_s�K:�/�k���\G�"�L*:����b��q��=5s-��m�d5��p�(�F6"�(��0�b�����e�ʶ�]�.�U���A���7��S�_��A*�L��oڒ�Xw=��d���ӳ�1M�̈��&�q���$�� є5,mе����;䲯ё&|��{���I�z?��g�
0_/�0�N�U8��ᩔ���Oݦn2῎XXHl"V��:�.0`�p�;�Ǳ
T�Ɠw�U���E�0Z�N3Jvͳ��#/|b��X�<���,̲Y��W�G��i�n[����(?}��-c��ix���Mz��^0��"%F*�i���i�	b$U�u3���My4t�����?Q��a�ג��-�C����0�s-�4X��E��O g��'�ۈ�.c�h`[)�Pu��s6���?���1ހ.�$-�ٿ9�#^���:��Y�d�r�q0���x�c6�[�ٚ�E�O5�v�4+ޜ�*�'�n�h��Bu��]l�l����o'�4`M���f�t�&>����e���,�۬c���fJZ�#QnӢQZ�s���������A?����n�û@� ���zY��|�*�ꇇʧ��+�ԯ��?��*���F]�RM~tm0{�&��������uɂC��?�K:SҵMD�|"�nK�9���.#֎�:��`�ڼg�Qd��.��(nVPg#�E����E祻 ��$�	lG�ۻ<�.�[V82oE]�R�4�t'��6������%�����ā�c�q\R3(���١B��Z�j����psԈ���|˲�`��<��x�֚ޠ�==b�2���F�Cr��k�65gi��!���!���)�Aw�#.;���Am}�H��^�~�L�ݏ�Z���W[խ���������4�+���։��X����x��=��$��kD�ø��O�H~�-����E���/�V�͙�}3D4�sx��|ݾ�����A�^W2jDT'AH.������noB�>ѝ�!�rM�-K(QH߂t*I�� ��}0����P1a��Hy�>��$D\���7�s�)ݻi��,�wƅ�a��ژ�!��Z�zGP->�
+?5>���CEö\N�0�C=GcZ����\:��'�K��?��x��#������{7L�L���S�M��$�k*
�>��]B7���d
"���fʊ�����DR5PZ�x�[|�SJ��x�C|(�,M[��d������h�:Ec����9)���>e)��[,j�wV�Š�V�c�_���H^?���6�F;�������h��D�<;�����r�a'#�@�&g�(BR��!g���w��N�o�����`���{�A�#��a9V�4�������V�B��þ�OM@�L�	�r�]br[}%�<���>;���LX�o,u	��Ej�T��6b��'�PA����Sь�ir������1��Qa�K����׎�C��X�5{�n��ТW���s�"�\���=���WB1ǆ 5���W�Y0��Ŭ�Fpl�{|�<��	� �ɘ��O�R��;=��"��=5q�Q�7��x)(�`ɩ�}�w0M�}�����/��N�P�Z^���i�I	���Q��z��u/p`�p��E@eLI1*Y��h������?�e�������GϷ���+X���.��Û�?Gi-7��v{����Px1IN"��d���'���I�0���7D)�D�^AMqaY�m-��9���6��"�n�gA����b|9�U��G���SE��P�p_Z�n������<g/�Ä��-�h�����6�����#H��B�����U��F�9�Q��{j�i�̼y}|�Ք�VY�I}��ɒ3�,�*��8��vB�,���4�,�|xAN����%\a�s��MX垺k]X[lOqx�|
�!KU0_�E*UT�@l��f�t�$��j
������j��6��YD���`��C�WԳ���$�%j#Ѽ�G�?�_�Kg��"��P��R��uڞ�nӥ&%�Խ���G��%Dб'Hd��n�g8Ͻ���s\��Dɜ���W���oI�8G/-��?�D\|btL��Se-]���
�OH|�_������V0�(�G���\ҙN6Ɔ����4,!��'�n��8|.���խk7*sv�"�"�,�\T�Sf�i�E���PV
�H�o�2�e^RxȦm_M�Rv"����)հ�3�]���'Y%����<�nL{�X�J �MF�B�����(3�TϨ�JbF����6Z 1[g�G4q;��xG�2�[��LyA(['ӎ`�+������@k��ԹD� �LR��V�Z\���� 0g�]j:�:7?�0t6��퉸�E���&�B6g��FͰ'�*Ѱ�ӷ��=X��94	�K渥;��0I�
�)<�L��88����~��g~m=��&�[���Hfh ��a�Rq�j����x�Ե�	}Y(�R��dq��^�+=�x9�8_�%s�M򯝪�@n����Z�
ې��fWk?���\�����-Q��J�º9"��8���x;���k,_�o��^bQ8��E�ُ�_!"���i�C𹺃�5� �-��PZf�s�1fUt�^��<��m/�1���?��F�m�xb1�)85��۫�Hǋl�IL\�f𺳴�5|\�:���X�H"�o�-�x7�Z����ԣ�����͛��1�e�%���M*$ߊnRc�dy/���#�� Y��Hً�o��LY���ӑ�p'���a�شFW$��K�=35c^�߿�\9�����Jc�N�־W��װ���M|���ApP(�<�T�0�(R3F��
��B����>��1�4���ԇĬ=��q&�7��Q�iP����9n����u�Yl�/1U��A�kU��a��eq��Z��=JX����Uo�͋ܝ�_�1s6i�{�bg+;j�����:j�L������](%�/�c�ÝP��Xu��O�uQ���)WB��&�{wrM��(z̄�+��v�~�-Y�c��$�e��#*x�$�0��m�s��:�ڍ/0D@�v���̆�P%�Ȅ����
�͊��E9cZ��6�rta͞`$�.��=�4�?Q�V�q����s����O(��|k�d����YC����3a�֨��=y��*B�*�7q��^�l~���R��תp�#Rf���iM��s��(i\�`0p���A���h���gD�ei;.?���v����J���O�y��W�˖V��i���<�5�����$���ęq������%k�}ը�j^������a�U!��=��\`���P���v���K"����a��g���Q�S(�X{����#��SpE�҄7�s.�箾S��uAԴ?��4�[?��'-@�[Sjьs�T6	�_	�3�i`�|ʪ����J�p���b\^Wd���&����B߃�2�0�Q�J�{��򪭄�M
�ab��ʣxe.s`�0�F�D��I:7L��=n�^��(�{t��=TJ�T�,�h���B���Y�����g9�}1$�P�g�_�����_1xú7��~ޮ�$-HL�Yo
3G��Ix�o#����뿋VC�fo��JY�%�w�R*h1��t<�ì9��,�Q齣���8��{ʭ(�3먎�YZ�A봊�V�U�6^7~�: x\�*<<z����YR`�kÄ�W����Ɂ�?�b˖��"K���]��0���W9k���;��.���_�tPIA���a}���s�0��ly����)�.I0V��5r[�5�P)<�� n��^���(QA���V��+�v�E�줦��q~q^py^������df��]���b���&	��>��� 9��){S�R�gA�y��(�h;�@{R�E�u�t	H[I�%�?�LN�m)�;��̌���;����������UU%kS�U�*����C
���@�F4,X����XCzK@c5&d�#���1C���U��.hR���2~nA�}���s���Պ!E���zK�>�^
���'��b$RLT#�N�P���j�6��J{�1a��0�.U̀�M	 ���]�%��GQs��{�"����N���q��f�V�N�+�wGS��NG�H�Sя�4I&'W+.7U�H�Bs�/:��M��v_��[P�����1�
�v���D�3����onE�l�^����1����A�3\rZ�4�s�������+�Fg@O�J��4���y0�F ��V�U�Y���8omV��v���\��79��S�G�y�9�gD� �ւ2Z���u�B܄d �F�1'ps�[�3w�E���u�Qm�T^F�8�J6�}��y�%x�5�`��'��o��ゥ��ء/|��	��_J�=�V��F�c.LX�@��8��5�\��]�J4�?�[u4��S,�2 "�Ja����k���
MB@�f�H���^�����P	���:V��q����Bv���e3l�