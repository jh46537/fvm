��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbж��ъ�]���ts�c�I�B[��>U����ܝ�N��Rɬb΂�b�`��VfR��w��clf�e�����7(�ɲ[����k�Eƹ�-����bl䎟D�ɡ�Nu��F�V]12���ʾ<�(l����۳���#���d��P(�F�nq�ￌgRhc��s��/^}s;�{�v5�����m���ؙ<8��LB�=�������n�*΁Eճo0"~�_rl]�cB],�@�I�p:y�IkI��̋���ӗж�f�)���'�gAL�e������v;�����B�WuܐO���-x�<�?��`�j�]~/^w�(��c䩯��<�R[�h|��S��L��ߴU*�
1~����ÆF����8�)"dO&�$5Q��Ϯ�)
���Ж�OE\������D�$Zn�l�S�+����/����g�!C��`^�� �#�� �J���H� ��nDU�-��5�e�w�x�})�<M��p��\��35��+��4��*L�{���>Կ�V9���].�^��"����!�8��6��ҏ����g�=�&<�4�Oő�*�~��"�M�wM�iPNQ���1S��'_���0 ��ͱ��$��N�~O4{ɖ�[_�v��H���_z�B�S�f����>_�?~��^KUb��nu瞈:��%lӌ�c�5�s�X��b��7���Z'�i'����8�n�,mE�'�T���?�읍{��eq�/'m�Ԃ�n��X��S|A]��3������cHExY��AM���_�d�z�"~��6g��|�}٩|�Z��;v�W�	s)t�8w������������UD�ow�v(�~Q��=A'lT�-"4�GLG9�/�h�q�%&:v[H���ȇ#�۱ۇ`��9���K�Q:k�	������"�~�V�L�sT�Y�9/r?�#D�y ]��A
G
Һ���������g�i�>f���5|�����X��/���T0PT�#�(�C��D��$|C ���
V����E$�|b��>���`��lQ�V�+d�<��%o�&x!Q'F���������}���Eٕ�r��o���wG�/�����%��Ts�}�d$��<&��W�-o�B���	�3i����q�w͟�u�� ��ǎ�"�CտFa��QU�
�ȭ$8옴WSM���%Fdr����K�ޭH�ȟ�|#<Ĉ\�G>��el^b�(K`�;�Cbmӓ)�LV����5-���k�̬p�DU���Ѣ�#: �'�m���冇7�@�n/A���qn��+�;z$(�̼~4�kq�q���Q妼>&]sW�V���?貇�x�Ƃ��|q�p%g���+����AL�
���Iz�w��1vC-^I���$F��Z_ʐ8�_��k�U��K���?�ө�N�8�̝դ����[	�4Cǂ��*B��S\&4WU��q/Λ��2ƥ�3�!4q�[�6m�,��T�D* ��tm9S�o(`���z	8�f��E��HE۾�~�E�U��$�o���ϩW�U��
��~�u�hpR{���2��F����U��"e��Syo���f��-�`ȂU��po�` _�N��_���{H��t��B��*��˰�d���?I��K Jf�(
�}�D>fU���p$���W#A"��b9�O�����Lk��~��k�����ѿl��]ǘc��~�rR���fU��&�^y����w�u5��&@$��[OF+�u��of1JVn��'6�qb��h\W9��0Y.u�m�i:A��m^�mF�_��5__��Fԇ�Ā�?��k-֞؄)�" }�Vn��x����7���p|{w+�%�D:%�B�c�4bC��d{=������H\��W�)��c��$�'`#�q�C�f��3$���fy�I��}�;�/(\c�@ �5~lLcH��$1r*ם槟�3ֈ7��B�Fr]�ૡ��������(&�(��4���x������S�^��ڲG�,+�I��� J]�e�l�ݴ<c���&�)<,��\uN�;�?-�4Ja��n���i+Sg���^�>�+�--�=~ipE-�
�^~:�%2�W��_���!u�5 Z��,W�'�er��I`iw�o���{�qt�/�T�5�5@�:,����T�=ڊY��?�!�L?�hN���������"���S�*J��^�p���-��������hF�3�����̛�o �#u�Zˇ��v|&F�6��ł�2��`��I��3�ܬ=�e�>>��=�n.iT@U�@����,��E�qE��"\��.�gU8]��!|�\$�FD���`�A�p��~��s�����mS�w��!�gD�=���Y-rP��WT�5w� %���y�a�紑n��?����B\�Hh�?8j<9.y�6O�@���o3~7�AI?%���ށ���,'���Y�^�ݲ}�t��,KcW�"��-3g��L�2Łd���q�-�}\��%��R!�/�uv��?����Z���4ԕ?�����)!$3���?m��:�1cա|�g� a�jcaVc��-Q���A��,t���t�n�ji��p��\�T۶j�V��g���T��0��';��t�v�Em����T�Z�5C�� 'vq�^+�cJ���"�c���
4��^�����w�]�!�f�q�g�b�D�B�Jo�'��F�v�A�6w��#x:�̮GV~�LZ��Z $�r3K�h��(fLy��<L�}����Hq���ǒ����PVhL}-o������_9b2��r�,�.G
��m��{}|�ح�i�B�`_��6��2���տ��9c߅HƷ�j��
j���ڈ�&y��୨h��5tGu+���V%S�a��"HKQ9����G��.����h����D8�:�_%��1��WE���p\�0��O��
�����|��uno�a���맇�[i/9�Kb�dY'��]ꠐ�ڲ�nd�.[�I&v��;I,�x���hC�&k�2�:�w����.�-˿Y�$n3�g�砗��	�T���b�5�.}g�c���N�X���k����?A�<9��cFW_8�b�R�ԯ��1�N�C��~��QbkD 1����am�x�7B��g��*M�<;R�/��G���T�-�ukuG�\�(�AQ|q5�����W�x�=��C�E�!�z�����<Q��[���2-�ռ�.�3�W��H��H(��M��NB��;�nG�rGr-��ޱ��X�>�T
׍;�!��ZMy�'��"�%o#憎7\~{���V$Ĺ��d��/�~D���e��(jɋeJv�G�D�7�3��"q�ڌʋe��A�{��H>��༤Yl�����a�\@P��4����o�l��e�
ue�N�!L����x{��|�K��|�'+��?L�9�[>��q�8h�i��o��Cޘ�_�gi=���|
<<�8ѿviب񊢒.�8.�r����@��t�H��E�J����>�q��4�d��c��#�n�B�;P;�\��j;�1�-�4K�։�l���5�!)�y����[.�/�:���G��c����a�l�H1�rja�au���k����q��oC�N�{�0�%&�(4��A2Ȅ\��[��R�/��1�fr�[�2Ώ����\g�~W���+�f�f����ٴ��z��������y�X�>����w�Xw���_��Ji>yŧ�����v�#�閾Ro��:ʱ8S�M�w Izl7Ay����xI"�X��x����X�t��&f쓎���%2���h�p�q�J�'�����0"&�b���2�>'����g8���=���`�@���=�� �V�ȸ�����o��I1ɿp�'m֦�/���X�/9&N�1r�9��yQI��&�~_�ѣ������s��4dB^�<��C���ݮ������:���������m��<���Wz���?
97	D�E�� dB�JYRsO�?0�"�{MK�߿�3�X��8������^T����n��Dԓ��42�`�W��R����Ƀ��B%�p�7��3�� �З���G u�\���`1���8*Ϡ�7I n�,4t�K��,؞_9�3�F�Ϟ�4�]ֻ�Х��-��¦!`(�I�se��Ju�8��Fp��o�K
��%� Ҍ��yXs��0�����.��vc���b�2�2���O�^�j�46����v7�~�+��Vu�2恬�>\"�� ➐
b���7䁆��6�uH���,#ћ�Y�7���������6���ً�*�:F��7��Jo8�+7df5{5G�
��m����otK�����O:���z&�v�vo��S��H�9U�HS�em�4YupP%�3�t��s)�<s�`N#� 7�S�&-y�����2G#�2?f����8`��.����۲�š��u�-�����ɱ��X�ձ�.z%3'�t��x�=\{3y)QЪ�:�O�P�'\��$���_�F*Qk��Ips� Ὲ0�dxI �x'��W�D*�*?��	���tC���2��l1���[��}l�d �������3�`�+�d���q��;>��JE���Ys�{}N�W
R��%&��O�ҏ�9<k�o/gq�f�d�c�e�������ơ7�˼Ėl�#zT�,o��0�����|� &z��l"�d�G����.��9�|O�>b)Q6VH�	i�O7�q�j��i>���E�|h^�����d�v^D.w�(�kh?_#/¡����;Wz:�qs���<���q�8��^>�g�.�o!y_
��
蜓�h5��+38h{�y[{qA���WҫR�r�\	C@�Tp`me�ߘ�h}�ް�������]6��]?&t	�������&d���)�@�x�$b���ْ/*�[�?��3�C,/aè3�1}ގ����lt�fܥZ	�[ٰ����Z�];��:P6��=��W� �H�R�yt��5�kz��6���evǳ2�hvി��锚I��`_��J`0Y���c.&��zc���cc������#��%>��Fd���hǒ��c��0v����Ő��J��8`�j�z��廬��=�֝�9l�s�r�x��x3C�IBi���Rb�I,w�#W���"TުI�X��5�oR̊�x��&��|uщP����u��<��y�4�$m�,�-eḅ@/D�9`L<X��D=ybZ�L�c7giH��I�����l����N}ZI��&@)��FQ�6�W]��P1���J��#��R��q��(�HOC����g�����RWoVȾ~I\��>mӞԯ:�:^����VLggE����d�+{