��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb5�	���uYC�т��z�4��Q&�2�hv 3�����,�.hR��{��+�;вT2]�	�T���D����]s�Wn��y4��{�hY��v���ɒ�s��2XD_IlI�j�5 /QR��C�Nv���Й���8	!+}�t�-�4w�
O�su��S���.��g�l��-���9X��D>fG�	�*C�rF�Y�j��A���
�V��s�Q�>�ʨ��+��<:�6�a�g�p�ɬOB� �K*$�hw��ᥣ�7���xn�=.��/�u�8� �7�~x���h��4��~A��+&��,��,���)�0l���P�2pl��}��˥���^�hk��}��N]Yr��"�\=F�ܤhο�YZa�� s����w��ߏ�I�j�4�0|O�:V\ЄsHd=3vm�׀6A��S;Rg��҅Vm���8�}�㣢늕G0���D,�|)d��sYW
�]a!a��lUs�JX��k��5�>�C}����P=�HW�w*��{)�ʈ�V *>�B�\���
Y�ZH�?Zڽ�`T�e~d���1��e_�M��4P����)t���K�E��{�ȹ��r��tı6�����;��m���;��_+�w��l�-���~w$M�H|��|q� ~�b)�Z�4��{o�+mw���*k/�sR��+*���3�V��{�\�)k-7��Z3`FC��ݢ��q��z�	���hZ���VG!iv^��nڗ�5s�I:����*����Е�j���é���Nh�����LY����k�rrΆ
)�xA�\� &@6]=�B��cY��y3���i�ü�,{�R������q�:6�K_bXI|*�	���F��7���%uJ,3[`���k閄Ϡ� �O��$�J4'��N���l��63�LN6�ƗqH(G�
h���xl@����aHԛ���;�N�y��5�Y��e��>{Mү��*s��;%�ٿ�6�.�b����yVf	�kw��8/K��Q)Lv�Obg�Xz{9�X~]�#�$KW|D�C���?G��� ��Q��x���&E5pe���w}eFT�>4�K�]�./$�$�j��E�@�]pq��p �;o������=����˻]����{-�f��'������J�p��%���=���2t�	蚑�8��f���*��~�	|fj�ơw_��s���I����R���B�
�VTs�����fE�.��URC����Y�o�ڛ�b#�t�9�xx�ہA���Z����O�N�?|b�]\\6�q�Va��*/2��J��2�[m|~�c<���a�{b"e%��;S��ǆ��S�f
4ʆ� ����7�+�F�e��wx���;�����A���_2�m�N`qX���������[�ss@<�H���nA7.rlԱr��v������S�T�{�4^��1��1���)oj�[�j����$1q����i1��)��rb����O���B3��I�p�3������*�w�pb���t1��)g~&�bQ\.5���6�H#	����әhfϜ"�]=��D�%�����@(#�6mO�e �Ap�
��0v#	��6js�ON�T%>=������!�8sFaň�4Q_�m�r��tQ�U�����A
��"7�R٪*��3s���j�N��Զ{����	���'p#x��Y�d�F�oq�F��n��)��=�~cJ'	�4���N��L%CRqǵ'��W�|�T�s�TP���6Tg��@8p���zҩ��QA4EuA��2^����f��85�C��X�����+��l�@��bA0�/��п=ݯo�A�Q��1#G�[����*�ȲȴE|f�v��t���g=_�H��N��Ȫ���F��pTY̽u4V��Q ��U2��BDv4|G�o2C��D���R"��Q��OБ��łE^J7�he;��p���u�ͷ��|iB�2�b�6�!���d�'����!4V����;,R���D��H����Q����Nw#]t��)��%�r/��;l]I6>�%I�����lȶ:lʮ�@�ᾍ�c��hD�}�1?M8���f~ ��RXI������E�_�p�����Wb�N�kݿx�x2��H���辬ڷ�ntcWq��1"K3u�̷':�CݩxMܵ)�_R�/	(���:q��81d�C�`���9gcY-�h�i\H�e
	�0����}8��gVc�^ <����j<ES�k��Y^TӤBlo7�W~�PA]�$����SVW�ѐ�X�$��D'J4�ԧ=z��͎)�ر���z�NJ�y�����Ӻf�^�Ŗ��g����o�!�k��}²����X�$�E��H��0׸xhL�Gi����:
Z�3���r�|.���8�	�G�7E���˥pBF�U��e���h���h�}�#�r�|��@Z�����p´�ʭEM|���LDb�r`d��&�.��E�
�5yr]*�P���v���hR�aً��4,j�J��5���b�������bAh$�i��M�K���n�� ��>�ߦ����L�O-P�*�9��<��Lw�vv����{��(7.~_����������-{����3h���p{'�|l��b˽̒D*����騘*Dy����.�U��{w�,ce���:�x[�7���ZdZ�֤�fh��.W`�YR�������Vή���w����\�b� ��9���:���Q�����t��������8:HZ����������&~��Dd����H�b�C�2�s5�8%�K���E�!e\��}�_!W�,��}�~TV�:w����b�&������W��FBv���.��p�>����cw�!qU��Z�MG�d-"��b����Vr������[�K:��މ����	1qދ�0��W�`u=���������4CJ���7�c�jG��EXS��3j���ֶ]M=�A��;�J݅��%���R�^����<4"�G����NVV�|்�V�-�Y�Sv�HIo%�cl���&#�i���T�rn'������H�im�ee㹧_(}kPu�b+�9H�^�Ji����\�����uR%�P�h_:��bO*w����x��P^c��~����T�(������Z����@A#�r�׺x�)8����6���(iPEP0��HQ����0\��Р�_=��c_@�$uP�uޚ��މW�.�3�<I��C�*�%}�j��b��d ��;I�)����Zc���كw���ׁ�W�8^�1�F��֤K{>����tJg�^�F8�/�e|w������� ;
��e��쟁��P�����.��Y�F�+�j,��*P�����A��3�!4�k:O�~qȆ1@�:�ꁲ\:QZ�U�0w��Q�o��z�P�R�����gb�p5�G�A��E�c��*������ag�Xi~�\<ri����G�_j>0��z�f-�Y�,�kHE��|�� �QA;�2�O�N�@���݊����&��뵆b,H��h��x�Vi�U�`�z�� �}���
Y!��
��k��'�E�p�?Іӱ��-蜋��J���e�<���&/L2n	]�EJ[)Q>�����q������O4+I���[·Kk�\@ژjf{>LpH��R�SC���ۅ���l���������:VN������QgP��v�"�)����ٽ i4�	��em­ž��򩕜d}�-�1_yO��G�B�UC��ֻHs�K��B��X��O��ic��7��a>�z`I|aȧP�`�jBcHua����d�N�lz��ݞk��L��|��i��d8���+�h��5�ZF�d���<�RǦ�N�@�A�׽#�1���vƥ�;�t���<�yCja��ۯJ��I�i����9��y������B=�����y���K��i}�yO��c��b��_�
-���j���'����βV�@���1"�f� ��/Z�����F�X�F�����o�%;;���in�;�|<��������N��XTJ^���徤�]�/԰ɢ�mg4M Ü�A��O-\�7$zɕ{A�t7[j^�5�x�����K0{������9/� ��[Æ��,�u�{w//'�*�?��M�`A�*B��'Kq��؆?5��_e@��]��U�!�|�Q-��4�@�!r�܉6�z?����Ȱ0gk#�V�S5I�W�B�]�7U4�zl�i��!)Ӓ�Ɋ���ޣb�F�oKt�k�sб�B�5�Q��o}P"t fa�3^���c�))�t���J�|��������Z)�.:D��x��z=�Yj�LH�14��}/��|�6�4YS"��3Ҿc�b*�z�����,��'n��d�}�N��:�L���B���n�P�[)*��������= �ٰ�b�����\P,��yW�@���M�qtM
(��-汮L ���y=���!
���50Y^�]�B�}Otz�i�L�& N��("̗��7������YJ	�ǻ7�N	W�'�$5]?�m�'ӣ���0�����oy{[�cq�b%�k�d/!O�q�E.ir�.kwB �(�(� ��G�)�T�g�f;�F^�2Z���bs�إ��o110*��:��V���wX��5w�G����k����$�Ch�-Ѯ�1�����F�vT���q�͢����ǿ�^P<sO��U���������˲���"#�oV0��Ɇ�A+P�+2�+B�$�O)�ȳ��֑��
�5 �Ɉ� 2 &�ɐ�c���G��W���>?�}�}S���z+���x�p*�oRVq��l��uTL�x�p�Ĳ��UJ��;�zk.|��]]P-Mp��̇J�1�����HE���!lB��~�)k܃Lȑ"cg��.�l�H�D�� v����[�q������ X�1��=[,7�}9����J��[����$�q�K�ή�}�(�TO��^���<�F���W��6=$�Ih���C�3�2���@�hA ���o�.��o��}�X�s�IT����'���J��Sɷ���s�P�]h�EH�ԉ����H�r/��M�Ua�Ȗ$i����jS
�%�Gk�Լ�{��Ĉ�,�9����,�UC2KÂc3e����O�<��.�`��@z9h�|�ga_�Ѣ��4�,��f�����	�pp�0�>�C�U�Я��WPNP@?i��T��]���Ĕ�;5�胟Ih�����������ˍ[Ut{�׾@��Xp��8�U��kȃ#�YA�'�hb�e8pZ����vYF׿��yer�-���E9��:���Iމ�{�$�`}Z���ܓZ-�V$@�V�
7�F��C�L��[v�`�@v�>k&��k:G	2�!��F#]��E�>�J���R��x�%����G8[l�Ӵ	��l�l�F���ܪy�������}��� #/5�� ��A�,����w����)��<�7��US��� k�,���-�k�z�a��'���@��g��ˁZ�n�ڹ����G��WCӲ[fO�,����㛳�ܕ�ش/ZI4U��y���wOہų=�8h��)�wAӎ]1P�HMr�0����ޞ�0��r�E������͘P��U��\��]&��z�cb�ɥMiD� +��::��T�	u�6�@��+YM1��?c�Af ��L0bj&!y�?!g��� �Wwq1a5�?M���:��S[1�/�Q�f�!���  aE�V�̟Rl�\֚*/�6ާ4�I�j�B�U���dL��<x����I�������f�f�=�e ���h��FG
���9�9u���z[�n���s�t��X���#�}u�g���zW0���98v�/��/�Ź�?]U�.�f����d���8�a}�U��8#_l#e=����C��Y	�Μ]�p� �-��YB<�\]:�Ds,���·W�hS`��9����F��`���@eߘ	�-s��	3�(�L�k|,��;&��ǂ�af��a�pR�0 �-���2
ɤ����SOZz�}���PB�@��l}ri���U�*|N(Pk�Jf�˿xhBb92K��YHM�`���K0��.9�تM�:���v@O2�e;�+b��IS�4��i��5���1QY��v���D��%7j<�gB�������ZY� k8ܦ �>����p�;0d87�@__�R\c@����D]��\�����������U��'Wږ����Vp���aT봌]ۻJ��W�y\IJ-�_��,�w�u~�5�)�E ����ܭJ��R�˧�ђ��UY�n��"����;W*� ���/��1�+3��<N?�`�rԮ�z���#f���be���^�!,M�4(�O��cV�@΃3ڊK-�R�*��s��������w�ӏD"�>��9�(!���D���2qQVҨ
�40�x���\�P2�f��Z��ϳ�$�C��2��r����sie���[s3D'^�Ӈk�2�j�.��Z��O�A+h������[|ui���2/�̶+��CGU��2V��(d���t����8�$�	DG�9̌�D��/f�:�o��+'�IJ��>�6���e�4����`5�O�<���� }�ɔ_�1W���Uگ��GV��>G��y7��=2����d,:�x%֓��?��2�����'�"�_ �ɕl%WC�x��!�̺��G�AK-��IjxJ5���/3��/����8�1|��ӵ�f�W*�H�j��m����5�Uc������HܜiJ]���1��y�')|�6���a�7q���E�Y�0gJ\m��k6B�b��d���u��0�)n&��ӳ���c-�>�y��0�|֯?�M�~�y��PP�l<��E����2/�]�q'������.�{���.g�P�
|���� �͗ �u�(y�40|���<�_�����ZU{�Pcr�c�b�]B��m_��Z�ٱW=pQv��A79�����_~�ig��\����>1�q@�w<4���3x\HG���Ő�U�'�d��I; �'���l*^�'�y�a���E�L"�|���󷐣z�N�$��Q��pmV���n�'���P���,C�� �D?`���2z/֚vZ�<u<z�e��oe$CZ�(S�q�a\pL#s&���^0��:ж�ㆁ� ����܍׍�]�i3?DĿ����g�8�4��	z\���,�RU�.]�~l^��V�Elݬ��rͲǙE������Ǌ���\�W��p�װ2J0�^�H\�����A�vNrh�$��t�4$(^!�]�*��P�K3ݔ�K����鄀�~��ھ_��Z���O��q��\
zػt}�җyK\��
	�7��nz�'	Jn�5�{t�0v;�'�k|;�0G�����-<�1h�u�f[	�coj�d�����%�F����b������
T2�u���^au��y�:�I����]�0�#0ݑ�l]�A���� 
뒓v��p[���6;HsΑ�n��)2�)��2�rMzh,>��� ��<�,y_���Β�0hp�Vg���&�?��9�T�cZ֐��Wp/�~[���(����58/���_����Yb}�ͦm��^k���A�i���_����� ���h �:�#�{=�t�w���CA8����
�Y����)��A�5Y�u�p,��u'��+O��3X�J���es��qi�*�������U̖�n���Լ�X�LX%�4+^U$~^�Z� m��q_j�C>�x�1j!����/ϴ�ު�n:�A��)	�Ʒ��O_ӓ��f��EZf����J¨;�d�)�mKio�e�5`�Buf�+%H.���a����9�B)cU�w��j�lr{�JI����^�E������FS�<��Vv��o�����+�C�Qᰐ\)�a�����b�O�i3[!;Ja�C7�j�ڪp�X�T*�l�1�n�DJ�8
I�0(o���Z��n����	r� $��#�	����<���4��|U������olW��iB���ܠ���T�5p�R��*�hV��P�!\���d��-�����OZ��d=3C�N1��;I���-��$�d4��n���
�f'�*��>��ߋ3�C�;H���A^�����[�)��(�T7着�ۜ���Z�7��ϸ�� .2��"-���"qУ���!�jS>c-w�x)�g*��\dd��6�`�w���N�Ԛ~�H��}-܅��R�9���6������m�R��R��֫XS����H[��ǯj �YS�~���
՜�Q���k�v��gݱ3�Ԣb��h�x~Wv��)�i�ʙ��@����c¦|>�\j���e�4��K1]Ia�v��7�{t���K:�V�D����T?z����&~��ڢ���QMv��j��+��
RQ	o��#����C�Q"��r���H�Q������.�E^z�w�ԏP��<$O9��*(�<��	�-�Jީo6���Jw[~�=�ٺLw�O�Cx�f�Ef�\y"�?sdE� է�7��-,ag}��(�b�VѮ�L�ܦ�p���[K�`�ᎭC&�wM�ˁ������$��F�仾��RA��`���x�WR]�BB��q����߳��£^ۧ�0#��t�@��cn�X�N7Z�I�?����}
F떝�ѭ J�iT��8�YXR����m�
)�;�c��K��=����n�x6x�	*F������9��+�NQ�4���
2���Y~vo�=��*���%�5��R�=E�P"�5�嗱@��.X�9��D�E���D�Lک[D��2�MJ��GI��ד�P�=W��i9U����$�҃�8	�����a}�����!̩k���f+(���F�y/���=�F��s@�~��΂�<�g<�Ӱ<�"��`܍���*��N�������k1m�H�x^�
�.)����'�J��1 8�42�uߵ�ˌ1�9��ܺ�~��D��?���T�T���N�P��4ѱ[Z$�D6I�	��	�5�d�����1��ҭE�f�٩.g`OVD�q�:flCL��!f^��&���!6����s�ОGjl�������Խ��?�����
&H5k���)O���HI��e�	q�Y6+*ɸc���e�1�*U&��"WZ��k�;�����*�|�I��mC��2�&&�R8��Xl�b��JZ:�+f��h���5'GV�^��@3ŀ�}T�TL[53T��T������^����2�����r�m�$>fHm�M��<zWTh O�b�B����*m�g�-�U��U�����I�/OUj�
Bڦ�ib����Y �T�?��#g�!�Ywp�z��5?��q��S*·��K���f���\*_�eL�}G���-�h�:=�S�oކf�OK�:?'��)�1�\��vCn��*ӲCv_�,N�~��Jd.���e���+���3D!y��
0@�T+B��>4ǛM "�)�&&>�y�6�Bh�7���~�:>a�p�c9��P`U�iXF�F_��ڦ�Z�Ǻ����Qf�Bqp�X����1����3�4Ƙq�9h�eu]7Lt�k�P��������U*q/�]�҄,�c<y ��H�k���̌�i�'�Hh�����F���B&����H�jS�렋��]?G���z����^��8ex�:��=�m�h��h]�Wȍ�&�e��2+�K�G�.��(�]��?�-�^%�i��a,��2�X���|�ĕ�1r`�"�~��kU[��&.${�<$�6G_r֦n��у����1��c9ݲ�Еi���H�ܼ�����]�=�~�,-��-��)%��=��?x_�0bc�;�"�.ß���;���g"V72:S0e��ץ^6Ӈ��<�R_�}��!$rFU�l�o&��f���цc���7XNO�)S	߱㻂M\T�=M��f�C�!wJ�x6��a�F(A����5�����Ky9���ːv;.5�u���+�A�#�P���J e��>��ߎ��/�A�w1����l��B�$I���H+\Sl�>�CX>�7~>�(�P#����zr��%�6^�����:
o�З��V}m��j*��!I���~���¨:�2�[Z�σ8Z��"E#�겸b��¡�Ȃ�73p1��J�l��<<oC^��ĔE34X�n�yr�|e������V��U�|2�tF}�5�,3=y�BI�CmSCySi�d	}:	5��ө����[�y�:�4��/�J����ri]7�<��*���av{�ս߷�)�\Zs��=��펥0���j���je�/8oc�>����a&/鑾��<�mY]��X҃�7G�-Ϫ�V�1$ϔ�Z��V=B�fu\S5�ƽ���H���3��H�I4�ѡ����Y/�y ls���lW�]c�{�C���Q���-���מ�k�o�Y��`m�T��"��u7�x=�X����g;�v{Ef)�n	%EZc2�3��=��4�_��N�C�]�+޹��HR��#`4��O�;��a�:&�`d��~X�Xl����|TY���4��Y%8�
8�Q�5�y�����[N�i�+XC�sZ:H�(��A(  �*"�k��\,�f`U]�\�p����^��U�?8�3������d�_5�ȶR���⺴�h��I�9*J�n�p�.�*W�T�0Q��m��Ȟ�m"���0*�*;@ͯ�m0����*�����R�՘���� �Z�rb�����첯Hp�A���w����M�uT��3#�~F˫s��Ve�n�m=YB�Ԙ:���Ё6=�\-���t³w=hL͠v��w��o�P�q��,~�!w�ښ,[Է/+`�F���:�@��5O�Nd�ܐB�Q����&g �q�5i��LX�\��'yc��Nz���vݠ�9Sg��Ԟ�!o����~D��нb���=v"�_o�b�e� ��
���T<�'�0�'��L�A�&M+ �1�`�-�̃�ѨzJ)G Z1Nx\������P��+��#U�Sno#���pq�06%�[�E�[���Z��{���~B�I��V�����쐇�l�-{�gts�P�L~�L$�6{�keQ�F�my�Nh��}���宩�@�$=T����
����*J{�[��8��gس�U���_W6����	�rMc���cA͔(�ʵL�;�Ӏ��ymԛ|<4`vH]�0���)���J�+k�Tp��j,��
��O�lO$� 5V��Ow�1�K�#"�X�iԋ 
�J�O����?P��Y�RW ���}D�� �gF��z��9l�66��e�~rE5���b��G^h\�r��z A�����C=o$��hR�O�QR�6Y�l皦	\�p� ;QΓ�{��뢤��_rQe��P�).EeB[6h�#�
ŝ�	�7&?3A^9��zN�+ް<A�������?V����w���vU�X^MC_�<��gI����T�7߮#(;�s�ېwS�k��ܔ�
L�z��^/yxX�l39��(���vP��]3�N5,2������ON��h�SN3L0g���ތ��R�ӣ�@)��$2x�g}�pr0�V'Q�#EjƲ.0����3����}����g-|`n����?[F� M�:_'L �������']!$:�C���y܏��?P�l9�m���G��1�"/��?�LU�%��Få���*N��� GK�O%��1��1�����v�C'�4�����x�)��@�7l����c~���N�<�Z��)�$M&���q�������¡*�&9�I���
IH��<�J	]ϊV�!����������Ґ���8`5r�Ʀ�

~`B�E�h��!A�aGm�.�Bή����QEB�%�-9iw\.q����Cp��ez���x꟢�^_\�o������u����m\]�D�Ne�|,0Q���g���q�%ion�'��=����ѫ CA����mN����&�)c�0<��ȝ8}ԣ.3Q�R���pR����8%�9��[�{(�����I�E� g�-��I�{La�̓�Dπ����j�V����s�ϲ���6��o�u��<pgKLw�bm�]�{4�#�Y��߽���ZY�����E��͖�:U�;E!�(Йiͻ�8a�"p?���<�������U���@U����k�ت�h�#��]����
���Xu���a#G�K��/т���f6���c1��W$JۖFAu��m��9���+�<�>��9�� �mw����:^Z�y������}���{i]�ўR������c[�L>Q�1��jo�g������2��W���#̪����������6ӏڂpSb%���n���0����~$X�1J&朕�4J�6F����+�o�^�4L /�=c�6�۟?(��v�f[�=�º���u;Xf��t���S!t�uɣŇ�����$��p�h:s�Ċ��Y��ĉ�|�-�#����ܻ�'7�<pb��Iʛ�}(��I�F�ř�����vl�_��4�18.��vY���-��ː���э	͕�.�ʾՎ� r�
Μp�CG�=A]��7n�-�+�{��Nm'�8_���furD����&�"^���_ˊ�M��s1��;��5�����`�J'�'�8,��j�@Õ�<�O}�??l�ow�����O��F�H�����H�d%]�.�O��8��<x��iV�����Z�h*����(�^�|6��?X�ѫ���ߙ�*�u�61��ܴR/�ތ�����)��?�e�)BQ,��+����w��>R
 Ff�&����'��d��&�U��D���JhW��p!*2�N+��2�Jg'�Pz��u	.N�3R��AuQ~Y�CyǏ��
��>��hG�+�ʀ��H�Y���}N�ԜB���c�1J�|��.���]q�v� �x���Ff��&/57���r��<�MCPZ�	x�M�tZ+˯6��p�e'��`��-Zk�_��d(�10�v�G�5ʃ���ֆ��[�;l������@�(k��fA�2��E��,��đ����n�D�Ͳ�O���}�W*��-l�ĝ������,)�E4��}>(ϲ��*�U�R�xSZIJ\oK�7�8�6l���&)�T�fK}?����� ��hB��tw:���ϫ����?,�N����pZ[�b��Ψ���
w��0F�p+LW��1؍�hT�˿�C�������/�H�7sp���{m�H���]��rf��;pRw�olv������;�T���$�G-x���v�<j�Jڎ@���R����q���Dy��	�cXtK��]��`<������ٗ��2emr3cք�~t��UOp�<���W��|���'�"�Ƅ�Q>��e:!L��s·�qO��e��J���T,�Q��gփD����A+@�sg��h�F������т�����H\���f�j��c�f�u�0��:1����'P�URD�smJVWlF�Ὸm:ILȳY2��d�2?�A����k�_�(/`��1՚p&7E���� ��&�xcm�w[��F��v��)F�w��V��mԽ6ÕJl�Fd$U'�(3܅:csu|V���0v0�'�'c�S�V`A`�$�;l��yЪ�1�x�����](���/��Q��p�LXm"7pϝ��-�;A��hnD�p݅0p{%+��Ȼ��x(�O]���1���y�!�#��]�af�I�)ɅqC*����6I1u��F������Ҁ�q�KB����?��]�%,Ҡw�-���e֮��-,o
`K�Z�.D��S���,�ko`�C$>;��7��h�]�c��sšY����Ms��e�m��۹�qz)��_Ξ;]B��
$U��\V#��yߓA��G,�x��F�(����X)�|��Ȍ�x2'��`�A��'��y�(���10�<(~y��D��[��/�t�%`��P�h��s({DGfߘ�<g���	�l�L�4,��/!�Ŧ�*k�N`���a�9δ*%��O�V`D��m ����~dШ�@��"6�ERަ#�S�f�R&�����&w1mԈXY�l�}b����su/1�Ͻ�*�{F�Z�-� Ie�6�Ĺ
�i}`;���I�7�2�Ĝ-l���0�-2�?�6خ)V�dMϢ8�A�h�A�7gSJc����h��[��6Ԕ%^zv�����i�a�{�+������t�,����ml���(0�8~�ݸ�1�.=a'��FA�PM��~`ɸ�@�O�|-7B����|W����^��e ���"�{JAr"ؒ o�y��r0Ua#�:Lxq�o۠�06kErc�a�n�c1둰`Uy2�y}�p��5a��r�g�ECv��럘p7k�1�`�A\�9.�`i����
(z���8�a�Ve�k�-�#I �W�Y(˒��+Ob�Uϋ:�K��*5�Č��K�K��\�<e�uDW�M1��m����	�:�Y@��M�sʨ��&)�m��sڟ�i�	�NH�T�������QR*6��v���S.�U'����JՋ�������胛<��Ig�[3�.�|�B� ĸ�xsf��;��Ml�i���f�:�r=0��k\���4B\'U�"���R��.n�7��9�H��xV��Y��8�y��#���Q��!2�LV2�=*1�j�o^f��ӤqM��s��F��(���p�?u�{����C�Q��a�4�<·����k�#9����P�Z����O�V��3@J�S���~�c �����d� Kȟ���h�օ�[Nb�r�J-*Ҽ����[��!b_�j�/�SZ���0
��fj��=o�Ң�nkNo�P�0&���MR��ߺ��W�H���Ws��a����$�w�ļh�1�`̬dDj��հ�2�h쀮��N�W��E�fx�gb:|~�����g��VP��XvQ�uW�Jf�]o��Z��7fP�J�N�)yQ��l��;�T�ű*U*U�&Sf�e:�YU.�mA�����HJ���	5�._lտa�m�.��E��i���dN�boY�@YDf�\[C�
CA�ܱ�t��<�>�Ջ=�7�|���.Q�����}�/��C�Wl�`��Ǯ����2X)α7��c��]�����\Y�2IWH�=��.��1?z��������0���%y=)a�EF����(��%��K��@�%�G���H&x����3�I�;	�zh~�m��þ[N��H`6�fs�E��XP��叫���^s��G�i|_�_܍U��.���"e`~Q���F<H.�.S�o�y"U�\agc����ɒ�= �zl��D�*�	����䁕���\AN++��D�PY�>s}i)in?v	���q�!�Ns��gP�Z$;��C
o"�
}�Fk�/	��d�ݧ���W<Q%�������8xY�c���2R�S���t��U���pl�q�$�'h숍X;���
'���T)�N�9WP����6'F�8�!A�iM>�����*��5{�o�ߦ4W͒�3����/u��TJ�-<>�S�Ӷ�]'n��O��=u���Lh)#�U@�~X���N?[�r�0%�,c;���-�m�Ц_� !W_*ED�v����z�:ab�����U������dv`�
7��$x�f���Ȫ{�O9Q�ڟy��z睭f��rӛcq�`Ii��T�E�>�cw�)4��7�toDeXH��&!1$��l�Q
A�u�Hx��C�U�2�c6}h���a\/�S�?�tAKd�ᲁ�u�����p�66�!�.$A�@*�G����t���x�(�T���e�Ѥ�X�PyKIP��D)���o�׃��m�%[��gm�+⠽��vM���Q"������`�X/
 &wG����-\�܂�rҧ�g�p�.���l��D/��q��,�G���ֲ6���Ί��V���LB�.�V[#�,Z��H�N
��� �y�\���>�L���tv3��V�h����C!yW��>��R�ޭT.U�C-�˞�Ny�CU�~��(*�I��Kt=�uJ�ʙK���7���e�&;K��b��D���a�ί ��įĤ�Z2M����[Ca_������o��;0��pa��j��_�=�:�Mj�lgC���`
u��l���+�5 Z��N�|�xF�/�8	\��D��ѹ�\�J� b��m\?�Y�q�:�1�&�1�2BV����L .�o��/����@C7 z|<m�/� �b��1�p�2a���A�J/�����!c⿼���eQoL�ｱ�0(�w�s�4v���ZV8����#��`�e��(�N�*ŏ�aZ҅k�(��r�=�l�n~P=Gi���il�Kwd��p\��]�>�_ؖ)R���r	$L����8��2��#�(�@�����_�j��yA�B��Q�������F�d��d+2&MIH1�|䋤#���ty �&���m�+�}�)p|�L��j���9G���:cw"����f_�͐E�M��A�,1�nϳ�����_~�u�,�бnN�r��w`���!7EYU��ù�Ďm�>����ܠ]qM�F�rV�,y/�ln���m��*< �C�8ϒ��I�snb���U�l]Qw�8+���iwn��?��9�g����ص�Ú����Ѫ
���25xgL~�?��zB���2�)@L-��ώ{9�p>Td^|�a�oF���<B<!s�1�CSC�P���˲RF�����5���	���j?��ݣ3�����]7y�fzIa�!Z��03�S�Z[�~�����3�����𔍴&�<X�9ڂ�TI;E��3Τ3�R`^���Wv��e"��b.�;��Y��zUM=y	)|�������c���TSPx�m0o���`�#�o�����,#E��8�tcU����#]r&�����N�H�X����)ʜ���3v�d\��xS�����r�B9܍��3��h��{��%ג�t��r�."����p�����.%�Fv�LOGU���y��*}����Hay@��0L[O~좍e
F��ᢗ>�tT6%C����Hь��>\
�%M�3�xy������"p )����\6��8r��w>��ϻ�(O�
Hs�
ιH�]�*���2��1���hA���|������p�]�"_D+e�܊$�7��Fa1����k>	�N~�ʷe��-;�D92�#:��kl��"z��e죶(�AmL"����=���:��{��Q�L�q�E���$��Z�Tod��4��pIE�Di�*H=lq ��e҉ㆋٷ�����;�����0�䕤���7����U�d9 �ӽታ��'�b8�������V�c�N��-����k�b�a�ԝ#�d~�j�OR�<��4Ӵ��u�b
x⾎�OD�FF���8�mɓqq	�$����yl.��,p��Z��� S��g��
=2�s�mv ����]�<ڞI4��r�W���n���Y����d�,ns�n��� ͽ�S#`�9佄��!p):�҅��c@m�XsK=FӞh@4e_@,��$�{�ٱ��BBRŰ9%��W�)����m4F���aq��fIp*�����	��3-��.��z:��\i=iB"r�>O����.�ٗ܂<�:�m��.�ލ�y����N�QF�6�����'����y�-���gB��%��v���2ٔ^Kk�Pk~BY��;.Cl&��z���9΃��hT���)�Il�3 �s��p�1�I���G�[k�L�*�Gi�����U,�O�Al��ö_�^�,tA΄*T����R��F�Wd�c��r��ֆj�l�C�9�j;|+R�`ӟ�3�Y�k3c��wB;6��!�	�;3���Z#��A?ӫ��h˴�q��ZMbc��ȴ.�����L�Gm�c�E)��2���埫*h��H�HeO%:��Տ�I�olG8�a�����-=8��˸�s�u����i�
�#�7ܤvT�F�˷Z����_���� J�L�+����`�N�Ok�d���$�vI�8��:��Q�~����z���m��n'�FE��5p���A4����C�aK飑�QVr�"/3���"Q��,�Q�\m�o��Ԃ��d�.f҆��+�_���� ��ۊ! ��I�ݲIX���O�S���P+r]O_U�xE�6���:<Ԕ�6`��9���;��ܩ Ib뭹�+���eLUZI{'�)M�Ί  ��e�]�ܗ~6��X$ݻ �Տ�vT%�(:M���)G��he]��=
J�;���N�T�:�qV��\rl��{�,Vn�: ��\�̟�W!�������௫{�+,�Aa��U��z�0}��l�&��Gy
���-u�|d0��_�ص�&������vK���E�4j$8L��wek*�i*���y ��b5���N%�;L�{�p��R���5���u�2j��5x7V�|���r�b�0��KdV}bc�J�K���5Y�VԄ?���v��kP�{� ������"*� J���kF) %����L飨�J��}uVF��F�Y:��M\ӷK���Fhqa~��b0����Y"|�n�<q�"�I��HA~Z���t��uHqS@�z=����(���OP�)�v���O�77����SveH�y��8�qU�w��������\�c`���D��!։X�.�=ȦA[��d���"s@)���)�u�"��	7ns�� ����ԦI���?c�
P/v)��w�j��D���l�r�c^|�n!���S	������X��K��WCt��u䅁�紿b��[γ�����=1�c"o�|�R�q�BK"�~n�4F㌢@�>�a�Q0;�Go�5�D��.?vȸ�k֑,�ۧ� �~����-)eMڤǅ�u�u���h�[�&B�{'�x >/��le�O�NW����aV���G)w���5\���io]��Y`o���pO��'�eSL�ڣ�J�����Q�χ�6���4���̱�U���q����Q�]Z�@��X����u�{�~d�1�6��R��Â��u�u2�!��q��'��`�I`P��%�y9��j��� O�����W�j�BƵA,��q:�K�C;�"/I�	���P���k_�v�6Į{�Y�R �`��@}0�R��1zL�KU��oG!惐򄣾e� h���b=�䊽���0ASd��\���1�܉��	�O��� �'+���~��B��=��9�:��`FV
��퀯:����<���!H.�i�2�T�`���5Ӎr�n�u��=��$~��e����;g6�ro&s�t
O��i������_�e� ����"�J�,�����B�ԑ�?	���}��t��+gw�|@�xâDpZ.�?�}�leF��5t<7��"Ӊ�O (j7v'k�x�C�ٽ8�����#��G>p��߈��I����6���|Ba7��^�A�BW"�v>�Y�P��17�MYk�L3�5JQ3߆�Y��w�2�ي��a���f����"=�b�F
��e�U-۲p-O����C� V։|�5�*�k�	�TTy�c���5��i�B�[ ZlU橣�!i�?�1��Q9L~P�u��Q; &ob��м��/h-�s��gB��QO����s���_ [읝�����	f�aD�YL��F5{�V��ʝ��������L�(��w��7G�S�GN�A��z����c�M�!��n	�*S�J�0�d(��~vbl�eu�v5�-����v�1��|����&���}ӝ%�ų��9��	Q�������bT�l��ьd��.N^y����-�SɾdF�%ˮ$��۠72"bꂹ��"�N}����X�� q����wa~�4t���mu!��:�M�&?�`��]�cmQ��|3��l�Q�q�m4&��L���E"]�&������E�	1�_��,'�M���)��Z���!<ߥN��E��V�]I�ϳA���63�2�[�k����w�m�ʪ����bOS���	� �^�Mv����2N�'k�\{#O�=�?�oC�I�H��Z/@}"��GW�@8�f�y��'Q�c��g���2���A�g����	��#Ql�2:�;�V���}8�T�Ki^Y����O`�
���Eb>��4���V��7��F�Eh���=�N���j��G�fP ��J
U��4��=K�EP���dmp�٩�d�����km�w�c��;��Ӳ\������L�T�U��x�h�Q�'����^Yʿ9O1s�t���b�(sn��a"=��#��f�E�І|'	�FR++�C����:��g^�L1�_�]5.jmߣ�O�Tu�e����\��(���*}g:���'J���������q�z�U�i���%߃o��˝}�5S��\JV�τ''.-�2�q@�ж�|g1��*7��N�2s��9L�#;M6ݨQ�m�A�ۥ8hɏ/L8k@nl���F��~�Y��`j�:I��6NJUT��W��$q��c�3��`}�|"ToB�LT0R�2���������c� ����㋯�w
Ƽ������*�ڐ�]ߓ�x�4�ځ���u hOg����,��1�������Cak�^���씥�v�����*���4S}%̈��<K -3)w����趽�|ޡ�Y��F���D}cm� �f��`�^�(.WQ"���bD�	��_F
)�i?�^Q�
��2]�v��O��;�X���[]{&�簉�ݵ0�1�w�!���Lu�o}"��~��Brs��i��A�5�2�2A��u��6�-ł�v�������ɳ����b�����	�	�c8�TM���'��.�ݫV��,�_����]8X�_-U���z��_!���CsVB�JԸ)_-�GT�.��Pc��+~��U��}�J�������#�KS�9Yz@�D�,.��Ӿ��r�/��0�^!�=�/˥��h��T��S���+�zM�kl3�?���U�!	S�SŁF���� 8������},��b�SL��MN"�/��$����"���r��[�=з�m�<��uA%�F`<�\-m�*%Fӎ�td�:=%���)5�hq��\2Y����>VQW�s�4�����_m��`0f9{j�����b�k'M�L�3�|]���&�������%�F��q�#�R7ǅ�p[�kEU�{sn�
�T<��ۧ��hq@B�sEu2Q��&��R(����q�QtKy�Z��� fͮ�����J�{�=U�9p"�aO?!��*	�qq��cB"S1y�{d�5،�KBT���6֐rSk�Y�����-d�p�'K�8�������R�J϶N�Z����/q�|cE�O��g�ΰ���V��1֡}�;��=ip���#</]>�.�m�N.�8���^��^G�?Z�rn&b�*��n��k��}��X�`n}Ua�+���B�������tX���PL^�/��V�L&��n�[��*Jk3�b��0.�Iy����@�&8�H/��4�Z!�Y�0TiA���]2j�*!���l`b������C��6�n!Cݑ}̞�V�I�ּ/D7�s�v��EEs3�\G폩ahňt���X���Zb+��!�-���H���k�\O9�TϸS�Tmh�Ϯ ���}��F���dhn(Ŕ�h`(����p�s�����@E����f��A��C��}/�x|�P+��mD*�ma�(����@L�I�Tf�wi[���3��3���)�Ê�������`��6[њ�B�9H8 �	���֞���Bߪ��vb�S�� � O✎�ē����؊32"Xie� �-���"ǩnZ����W�I[,���j�������wJo�4���5z����ѷ�� ��p^&-��[�C��c��lS�Œ��{e�`����9t@ʵGYV闿oř�7_��p�j6����W�,z�E����R�Tg�	�d�48hݙ�m��3/�f����+<������\�4������ҡ���S�q��=���u�E�i�'�n�ԇ U�pжׯ��4�n
�}��8"hz���P}i�r�Y�6̬���;M��|d����磌�*zըY8���[Ɓ{慼rMSy'gL�*�54���dlnȿt�:�*>,piv������d�d��V[K�E�<[�{�Aq��0 ��²�A�)�à 9�8�Ƃw�Z�f�iJ5X�E�y9�j�Cŋ�V���`s�D��Yt_n�t�;qS_��Mu�2f����Պ�L��)g��^�f\�F�Z��t�!���5�^��N[V����Oe%e���$�����VB�~5�hF���J!�����}����d��]�ߴ	�>�]���D쒪ʠ,�TbWQ��
�������z���v%��T��s���_��!���I&�����2�I���D�Αro8�
�$��1a?6ܻ�Z�q�VN�\)�?�ِ��q���J����2q�������`�'R��q��nM���7�ޘ�p�k�������);s�#�J�qa���R ������Nܺ, ��A��Q��$,�2\�e�����}z�oBi�J�:{��~_c����� ���Zjz}U�
��1�a�r�wdr��� �#�ţl\5�[憎���1�]o �� ~�c�NY�U����o����ȉ+��q�@��s�ߦj���6�#�� &PS���ԩ�3�ď���?~?Oz,a���ho����*.�m`OP��i��������ֱ��u��܁Ď+JNN%��r��]k���iK5�Z�c�� ��*Jzt"�W�+]� �����6$��4}��B&_&���棕�NNdMY�i�h���g&)`|9��F���:��ٷ7bӪ�qS�$؈��+���-�]�G����=�79<a��|��!@;$C�&LjЖ��=�}��Uv�g��D�Y�i:��������y����J
;��U�юv
�:�H'��q�H4�\x��A�ۆ�џ_|�K��B���4=�Ep���h.T�A�]_�]���b��������#k�-����,,)x��h_
����{���G�)��Ǧ�hI�	4|S=p�J��澰�w�L�����x��|w�[2oS<͠��xs�#�B�ݻ�or�h�Y�~�%�Ճ�̓8s����19��O���Qd�qR�z�����zl�zkN����g�!��k>C�$���cFU�H�C`4�S�F ��Q�Q�nyI樂��Z!j��i*�E3o�R>��@�T�,����h��l==�G%Y6L�nf�����^��iy3ώZ���$=�w��=�fj�	�b�fq13���_�1�<M��E�u���z�;�P�C��k%o��GI7�
EWf��ru�\�(6Ty�,�K��?�B�C5=R`�sB�K���3ɺ����J;�ɣfwQTH-1�/?����N^B�����:u��z���D�����?#]�s����L��fѾl��0��uk�	�0�f�'u>n�z?�:mc�?;��w$�^��@n+ߗ|L�M9�+?��� ����o��]��>j�=�� �uM��kH�j�4��	ʫr�MF�IrI!T���=�Ƚـ��:��>��5��Ž\X�5r���o,��:s��1����ӵ�+e�%�����}w����ɤvXl�26h��s�ZH�5��/+�<'p�d� }[�x�pE�}��s{�ذ�qMo
�Q���3<B)d��qx�s�<r��穳;RJ����,�Z�a��Ҥ7��s�{dAaFf�ʟx���ϝD�G�GY�w�w��\�-�JY��5џ�ڭ\���(���a>j���.�M(�,A�[�Z��Vz@����1	�����T��+���˓��Nu'�n�9�Xͮ�!�4e��y�;��/a�?vX1�h��j{�jun7#e,��5�u��KM��p*��mC2Q1Q|�:�����A\�:�?D�jgx���
�0��������Sa��Lo-�����+텧�\�v���:�|��k��ia�d�Z$�5�T�k�%)�J8h��=͏͇��^3D|�T%���B˗�e��!��sEF����.��t!��N܀:項�k�Q;A� ������t��g"E����s���fq��7@y%�G��g0����E�Ut"�$�>Sv9��B�<0���'3���.�O1#����^���xP��&P (�$fmZl*Eջt#	�H���]ʹ�G�}VAտ4H����Z��_�^<������f���6aÖ<kޑo��rUË�JS��^'����T����$�]�#h�g�E\8��M9�Dӻ�yf-�&�̷�(��F��Qc���:�*�� �-�K.�U�yVq%J�Et��b�:K�6���u��*x@���ޅ[���\P@wj�-�4�ƶ ����,o���T�{��$��Ѯ^A!�#�(^?|�U�p�.RA�v
n���F�Zd��4=:c��zw#rg�θ���®IBp�O�@'��Ξ�~DP�ߢT�d��t/B4���t���A�����P�i��Ð>0J�b�����=�%;Y�C��Dh����|��F����˜�ٸ����]ƝuAk5K��.��M����B��9V��҃�f�����9c{v̚㋯<���嫏V�K�[:��[ߗ�~��������:kH�����Ԃ�
��D��p�����q�S����p�p�pwK�`�I|����x1� ѮJ��<�g� Ҷsd�'��Ɋp���t,P��r>Ǫ>��2��M?��q�v�е�E^�w���k��`��m�A[��6`pJLO1�\�)�\Th��xN2#6\�}\�W�'�b��C�Z�8?Ƌj
jso3�\��U2�#l�hr����8��Y�_5N���w^&����0*��U�m��n�Ia�CG�����~��F�3��G��Oc^z�P�?>�<Z|���17+��ib ��~<$�aH�	����k}6����A�-#���9��Uzc=PhC7g�5������6E�,KK��8&�>��P� ��alXъeL�_�:S��/����W_'E|�I����܅�=��ȾC������}�b��iA�B��Hؕ��^P�Q���G���zTh�)t�1r�4�Ĵ ~�ֿ�;����&�P�Z�uc�������X��}��5,�AR���v��F�x�=�Z�I ���k��nO�S1�!���A�g��� Ζ>�����tu���
;�	luK���䆨TRش�z��406�M���a�'�9T(��X/�k��H3DP� /��i�ay�f���c~��\��
��^������b�L'rwڏ�0����8��fJ~��2Fh�$���G�>�Ӈb���}֔�!OC�Bg�c��� z�uY�<��)y� ��ǘ���qmW�2F�r�~�U���9��q��7Xx.Fm2�1�ȋ�s/}�@t���0�Ͼ�K�P�R��@9���+:��z���d�ٵ!���>��
Ѡ�s�#g�.�@�,�_�������8�x?��x&s�o��sV���"!W�O+= ��^3���ӄ���Jl�ސ��5��$I>%7aܔ���))e<�H��F��݋�b�@r�W�f�J�9��m����]3�ځ�ЈL�eX5]w����R� �螴}2)���9s<D�>��W'c�1��J��C��荁�9k)Hw�d_������z�V������L��od�$"��h���ɉ��E*ɟ�[%G��u��W���w��G����m��\k�'��������u���"��@���s�8�,�ϕ���)��q��HV���i�]jLe�O0�?���2�Vʦ�����j�e����T%nn�y,����e���>��Gr4.��&l���@nbjY���(qF\�H��^�g�*3�G�0�C鐁*5`�w�mI3�ze�ӵ$\���|�J�V4O<�%"J6i��h �#���R�y�Ru�Z�7n���\"�C=���R�fT�$�gᖦ�f{���,����j�QB>������:�w
���JT��e#=vHs�7oؾ*H�ME��#k=r�Lv����hQz��%ʈ�-���P�Ѽ?��Wp}��5k��c��Q��bn�}�oә�NxU5���hg�Y�?x8ok�)�"̨}�"eM?�E&���ED5��ֺD�uQE�}},Q7oR`c�n��X�6c?�������	��WNe}�r�Gk�&��AT8w�4��Q���P��q "h�q�"l�'��G�X+��
^�+��F�$���,I�j���NVfH��P�T�S����h�0(��SqT�	<6�_�7xd2�J�rƿ@D��V�����g��|�n��˘��~��R�c�GDnP��O0!^��A�NhK��;�������C�j��A���
�X�����5b�+�@2߇"���$; 0�Kǜ���=|e�����>����ȚT-�jD�g�ׇ���Aw��Bڧ�g��A���|�/pu��Y�]I��)܀T 4�*'Õe]3B��@�K͊��0�7�g� ��N�v��x�ڡ����{ظ�쏷P�6_ZM�{2~��xB��)�O�-�y�7ɨ˛����C��|�3�ts�Z�3�9�%qc_:<"���p�ML!/��X#�xܖ1��ea�7Jd��D��(�
��}��9 uQEݾ s�(չ

K�����@BG]��<_Z?��R��(�B8��|*J庈C�N�z|ӥa�pv��u2=�!p/ia^���W�s��& ��T%?;�Ϗig�m�Y��K��e�PVj䶹2 f��S?s��R)d��=�Ԭ�4�i��#$���Fʾ�e�x���c���iE�$+���[�����0�uK
L+�k�׮섚�����7G�is�D#��j�*�\�ׯ����
��nf�0��=y^��-rOw"
"���=I�I�
��h&}G�<*�!gψV�J�Dʙ�C!����4�a�eԚⁱ��/��><3H�vI�ˏ����t���9 M��=����
�;�qc�L����ŃM�t�)�.b�T�BB�2�E!W����=��$D�V#C�WX�3��A��q�9��&��pF��P��	P��|a�
ZqI�.Y�0��2/n���L�0b�q��x����o�׮�bs��L��Sn,X��\��S�D�q�0b��4^��I]��m���2eM}��;�p�if��ts�Q��'��1�H��q$�'�`�ų���%�j�(�r��2C���&K��Ld�'��_٬��݊��~u�֫�1i�)G�O����vɗ�������ӁQEw?�+f��f�sX�*�w�?�&�CZ�QA��������i���n�F��@U�hf���x�F���x��L�.V*��_�n��	�z�K����9�L�H�u�OO�cW�q�3���Ԯ���#d��]\%1�y7֍D*ϗ�G�N�oaX���N|�cX��F�I/�Kl�ŏx��������!�f$rC}�����+9)��b�_ tfB`��R��.����DD�fQ���R(B�CaӴ�2A��9jy�O�o��|�L�r�m��u\�B��RO�6��ZN��<_�U�Ar� VXy���;z�cg71��!T�`Q˽�L8�'9%�)��QفN6q�g��s��+�䰙����| :���s�}�_�q��ݞ�ŕZ����^T����8�T�ۿ��er�@=�|)(�-�P�}%g�� ��b@c&I�y�B�(���wR�����҉�Q[��´�>?G�slS`�s�ݯ����>��9�g�]xJ+ؠҞ�	���䜭�Q`4&���#��i�o����gu�� ���?Œ=�"?O&��|0M��/���9v(i�4�jD�f����$�z�yEPr�n�;����*KpF��5��b���U>;Q�����L�,�W��x'���z���˘1��Ϊ]�������]P�/��!�-�K�t����e؍ʏ�}�<z�5ilJ��r;�Lb'~E^�k�⟨&����&�3�E~F�3ik���;�����&p���c'=l��$��x=H��'����KB�7�~�#�cI���!k#�� ��Z����4�"�Qk�&z�d<ӍV?�u��t�Aix�i
�US��~#�"��V���xIbqȡb@50�+H.��}��xM�Ǉ1��"{�+�L��VKb�P!�p�3ڛ.�i�]XK5�,�&ڗ�y�P�����n�ÅNFr�������x|<vv"q9�ݹC��/l�V%�4y1��s�i�i�x
u[`�4K;`/�D��(Z�F�l�ѧܕ��4�r�In�uX��~��	4 )E�K�wd�k��C5�\A�yјN|�Z��>~� ���1g(�$q���V��rT*�e|��6�OR����+��b�Lt�.�7��^_M�Z|�OP��:�t�4��^��e^f��rw��GMB��G���x���d�����ľe'd��n��-�,�d�
GؒQH27$��@G�O�;�� ��L)�8�tӇ(�	�{�Z�/6�U�\U�۔�� f����̠EN.2ד���d٠kK���X�B�PɃ��G�b���dr��QȆ<�f���؜� �1~v~eW����{F�tY��\���#i ���\#.�LHD��H���ȫ�y����6�����U�Վp"��N%Ϻ�@ܗ��J8l�>���F��D�nJ {����F��*��>�ҏP�xȒ ������{W���
gQN���I��.�3����x��	��F�EG �ǽ�$UK�l�)�%K��
A�I D�/^�R����δ�)�G�\;k+���;-��R"P����o��#�Pb���dn!�,�W�2yt�wyc��5d)W� t�5�"'��e_���{U@ٺ�e0*��	��k!�f�+��9����g���3�_��&��^�)����,�������F_,`�2L \�ē:����g:"�����2o�I�n��y.����ʯ��� D>��F��c2���y�����h��#�N�,k��t�q����]c�Z��b�
'�ڒ�3l�n,��Z²É0��1���~�&��oI:�-�[b
�x��Đ����d�]Д���m�'�M`�	$RU֢Rg��lkW���!2�Cܚ������]��>�m+sy&��.���c"����2��+$$|/r�����?��*�hY-��7t���,�T�|`�M��rRT�����-���mDV]Ii�;�܆�˳aU#UVR$ɼ����ϸ ��`��Q���։�/9�{]���s�~��ƌgBs4�wӸ�[>�x{�vdiN5��đ�q�:'�yB�[P�/I.2���f�V6�R���k� Ds��?�Th��!<����~�������N9�,7ۀ��-�f-~��P��C��0��K��}|��_&�E橊���*P_���!R~��<�iЪk���6_�o��_u�	��4�OW��|���-�,����5_�Ρ�~0S�J�YZ�%ST` ����w��Y�- g��K觛���ӕ&�ȿ	��KZz{���u���� 6�K\v0R��%��� X<���4�e'���v��/� �J�'�����N���=��P|0߯�AL_.oh�����&[&�0^Z�-T����}d�[�7�U�`����SP$$ۋ�횃��"��µ��;4e�[KD]��Ǜ9���s9�Ivh~�����ѠTsy�r]�V��&J�y�Ƥ�u���1�z
�|�G}nl�>��b�-�ے��?��V��:;{��>�~���9ޭ�q���ܨ���5v�Ϟ#���w���'7e�ˀ�ɘq�
0Ǡ�|���b�g(��X�l�N��5#������Ӝ�}J�+��J�(�/�
�X~���7B�lnֿyF9���t-���3�d�h�������z�C7D]t;{-�z��~�)wI�gac�I�/��P��U�=�H�|$�j.Ff�] �����}&l��q8�U�L5�c�z��8� ��>�$���p�R��^2��R`F�f.���Z�C�R����L�-���c����β�Uv^�t�%z4�����m)�-Q�-�s���C���B��0��*s$k>dԹ�A�
�Y�� 

�􎫧� �x�1yc�$�.��c�N��:�Ϙ.'�$x��@��(�+h��Bڽ?*?��]��$�f�#�n�7;5��8�e`H��ՔdM>���㵆�CD�ԁ��~%���ɸA��9�+���OkC¥%bY�a�׃<k�C^ \�a�騽�@�iP�؀��9\vl>���C.�㡸<�),�W���R��m�O���4D���S�h-$+������~�d�������1ɢ�����:p"�ˊ���_1(-�0�w4̅iW�oT$,�8a�~$V�e��ŋT`��17���dճ�.<�:��w\��"]h��_�Ă�Q�lm16��C�u���T�c�}�{�v� ����I/�5�L�K׌jVBY���]*52��o;t��'O��d�A�1�1�W�qfX9/�ͦ��@���Z,�ɪ/���?4�^�2w)t�p�,7�� 6Lh#�t�z�g�V%iS���;���"�Cݠ\�¬ݶ?�"���e��U�#%�B�WHao����dp\��%1�IJs�	���$*�u��>&Օp�;�6b�>��܋=g�?�8N������mZ�����:d 2q0l*$H�-1�������twb��h�J��3�N�i�����ܡ2Y�]��۽�N��0pq���H���W����!�e���W?uT������tUH����֋o<#��̐N8��8�[��<��Ms��ș��;Q�rknB�,�K�@#h�_`�����Uha��l�Zx]W���3�#�qp�)�t��u�=eQC�%}�uT��Fk�y�&��=��j���a��^��d�j/��.��'���lr�����E )s.ǜ!Z�p-�<����X ˿����0��h�0�7�g�hG��%\�X5W�n���ţ��:S�ݦ��lv�3c��	������B�np+�C��虿��A,��5b�mI+�����(Q�^�h���\��83!�y)�o�OGj���ώ�YpP�f��7�t�����tf�񨟣��7ۻ���g��`-w͊� CsN��T���������y�* }F�]M�a�Ei����ySvڊTD;�>3ߠMv���<��3�hy�ca�aj&�K�.�࠺i&.p4D�������j�`����d]beSә�1�2��J�j�����	�c�����L�i��F% @��w�����^���c%#9e8H�]?�>}Οũ���!��cDm�M�p�g73�v��|��N>ֈzo$D��[�2��/v�C�j#��ȓ|�)�6ˮ`Y��;8�x�<���Z��k�:���»K!��b$����n�Br{P�I��Ѵ�ݸ�5L{s�*�?O2|D����9q&��b��^���9䏋E�/㰎�ͻP�z46��}1�Kf.%L��6ۼ���<N/���>�c�I���8X4�:��%jb�DX#W�_�-�#L�"/ W�l�,�fJ��t�=HAm!@���kѽ]�M(�*v�ݍ��@���\]����>�����J�����uV�,���դLO��{�Vg�q	kqp��[9ae�PV|Ѳ�㷑~�J��/J� O	�rM�p[��5�,��A����������k��i�mg����klc��|�wezt����C2{y"`
{/=�lP.�0�h�2+>�Ͷ�N�^���?!�j�>��{�3_l��$��Qufh��x��S�o���A��vy����';��ͽ5�+�Ȏ�f���CD,ՠ����o-�����LS��\�,��\�������f�r�at������J��3m������H�	9�*Λ�"ON��x�?!I?��-�O�����F�/���2f�$��1Ҕv����+Qq6�9m���	��Ct��>1s|TE����+�������%�wAO{I�b��wx�K����CA'�2#���,;���t����%q���!��E���&u�~R$���C���7�na����` (Y�I�]fT���wڳ���}8@�������=te���H���H���(N���[����+B�_�nؐ|���2{3%��*�����]���
y�tμU��}�XL�ƠzH��pIX��
�!��[@���ş�6r�i�9]s��]G�,��o�����`UI�����^[�?`�|���%U�N�
&���E�YEd����qA?A�)P="DQ�-���/'��}�Z`�L�l=���R��O��U�g��U}[�P�J4c�h���:)�į�D��4/������?�Gن�̢��a=)��,w2����fFs�y���L�{yW�@�d��Pp~.E\��f�=s��g����'J��*�~b�ׯS*��r�/�q����g쬥N�Cޞ�\��O����8I��v�2���D�މ<���1x�g�����;��|8�pb������t\w�9��q�,-_����3w���"-���uH���0V$j@�Vz���m�OpQ�}���;MP��.��c#'-���!%ut�Q~$�;�jo���X+�����˨��z�Ղ���JP�iQ0S���'ZE�$�݁����v�h[���h���14��?"$B�؝]<�_6�����QU�-i۽;u~O�Q�R��c�,Ϩ�n�����a{H����͒�X�:ܠ|�3*�j�HrNt�n��B�L"��c��aY��$M���lx����/���"���i7�|�7�wz����Q�o�]����>��*bH@$�V��_��wX8�aN�7{���!��	��%��D.�C�����i�U�2�} $m�!�@*�/e�#����e�u|� R�oVI��.��]��'��wyA(<'H�s������?)�>�?R�BQo�_�1�1_I߃�ご���"A�׃C����G�ː-R���O[�4t�,cA��sB��u���ZjPo�SfƮO9��ǚ`蕜)��Qg��+�g1�ښ�0��(�h��_��!S���.$�u�_d���{�+�J,�g���<A��NJ�۬l������?�RB0��D�g��"5��w�%���	�3�UH���i��!v^I�7h���$�� ��4s0q�6
֏7�+�Hz�l�j|���"x����)�{�]QH�|hA2���aQ�w��8��,s5�.��ϐ;\6:��v��I%@�� }s�HpP5�A���-�]���z��jH�?��`����Ɠ��>Q7�d�\۬90�-�[�7�����N���c�T��ۧ	�L���o��YǺZ �C(���}�H��;VB�.�T�R��2eHFďY��:GKJ�G>�ر�	�ht:CC]���)D2�����,�.t )��<x�~hg�P[s��{����4�S����R�$��B:��uu�/���ٱ)�V~��:�iI������eu3T��lrX��3s�q]a�uT3j�ө�ʂ��SԺU� �/E�̈�]��t��ɞ���Y����h���%ܳ�S��*P�'�h������y~�265 �Ny��r
�.W̝�5���{�Sm*�_=��#C�� Ix)�!��a�|�z�����D�9���|y��d�]�h(qT�;\�R��n5�):LܬA��/�,-��؄��!�|Z��w�J��$Y��|GSZ��5_:�RVKmMp+a,�{o�I8dw�ncӦ�"$�: �;'�8�D�>�p�ܐzt��R�3��j*vŘ�,R��(	D����"�֔���vu��/�ǪCW$mj��Ƭ�MƄ�6�3edx�R�;?���?���s��|�[��VC]�1E3O�R�Ui�L�k�m�n����͒������G$��7zt;@����-��%�]�D�ҙ���l�y#��Ӎ$d�z8�V-CV��z��0a���& ��ƃ�@Oʷf��%6n#��	���g��T�*L�kh6�`؝�P�����䚅���lc��%�ϮNϕ�����z�
=�f{*��`��Q(�U��:��צL���m�R�{Ă}*(9�hwV+������7J�cyP�� ��}�A��rJn�u�7LO�B���a��դh�8��������VX�@��Ě1��:�[�C�H�ܶͅ&_����b ���(������̺�<}�N�N����W57ɛw��ņ�u�}g��Q�mh�뚥E�^�eLÁ*�*���ն*j2�qt��+taXc|�dN���8!�y�HŊ�V3��&���
rx���[�?h!_�d��{&�ۦ���7��h�ޑ���tI"�uʊ�-��SɎ�� ��"�zo�A�GOWۑr4q`�O��]o�'j��SɎH����m�^2�9��'� ��k��?�� �����Ύ����k<�{pQe������x�4����h-��|�%�x����bH����ֈ�ybhI�?$zH�A�_�^���N�~���.���6���f�?o:�����/}/�;��G���./��з�fÕ �*8�W'���<@\�o��}73Mn�nx:ck������	�ޟ�%�äc�"�i���G X��'���gT�ن�	���$;��kC�v�7Y�pZ����\j�T�`���J��������a<��ҟ�2)XN�ئ��C�t�?�3�}��h�p���@(6D1@��v�b�區f�ѼE��6Cn@$6��;i��(s�S�{5�D)̐� ��
����+3"g LK���1��t뺎�տ��*���J��5�tZ�xO�cq�_�*�4�'8�
��;!
��4s7+���bո��-j����垹8Q��6��|�l��3&�J�w���7 �@-�$��9����b��&��Mm����A:���AzX��FBeS�����/ #�kio���:�Jdm͞?�6Mt����Wn�3Ό��t�FօkI�5A��1������D�շ�[��8��3r�>�H�9>����#�����Kk(O�����$� �5
p��yo���&|���\�\'_�;��@-` |}�uA�p�K���*��F�*D��{��*wVd]�s�}�'yBZ #���6_J5G������,�E?
R��Q�C!y��%F��y~ �Gf�O�"(~�ٟ���,�֍�zL��DF�����YMr[:�����4���H����f�[�\�#��d,�q�K���Gĸ�]eS���gX˲�z̾R��&@{��7�?�};ʧ���'�g;�����\(9^¸�hw���	��z>v���Ur P�ۭ��j����=�qC��L���&S��J���| RNhq��d#����\���ĐqM���yl#P��|�"����n�+O�F�L�js�~���9��0ܾ/���gT����F�v���6C�e⛛N�(�dk.O�mB�,����S4�a"�P���L?��v/��q��r^C�gaB̯����r{�%{���T�5j�[>`]�|ץ�b��
Rށ�֜-�6�0A�������4I��j� eiվX�m���F����DRT_�	��~d���g�rW�-��br����HWP��Pz�8d:4 �ᾊ(� �����Ko��i\���vؽ䩏Ȟ���{��æ��!�$�T����k��?J%1��G$o��z��iX�yn{��]������:3����pY�5�F��܄��RL�Z�<�N���i����p�+3���7�3�'�%J7�4~0A�i.\�Rbqi�ؙNE�����[�B+&}�!{��沶oX�g��/��
3D̞���'�a�qA`Q)z����ƺ���SS� ��{���9�Fnw�dE�Ⱦt� 4��{��5�TZ��Dyc�N��0�?�'���9�D[��D���R7+��-��k/lg|�nU'|���ݟ���`�;r89��nL@�9�~j�؂��l�%��D�{	vn���W $6�t<r���#Y�By�>�D�l��;��s����*����pTu��5̞�l�\�qq�V�l�s?X���Ub��z�p��<b���sE1��V�ȿ�TB��=��e,Fϝ>��R��I%�`lɞ����$�ut��)
t���DA�:��Z�ւ���^��7\���NvԽ�-y�9�,=dUƩrO�����1��`B\���/�)2�t����\@�7" l��Ε���;�f3��H� 8�_�Tug��D�V)�����,��ڪ�VV�$�n�����ȘN!�v���=|؆W�Y��3�S�L5O�TXwh-��G�dw±\��Y�FG
b�S�ROyZ�:�9G/���n��� A�K�X����������ѡ��m�J��:�sV
����G}[�L?�KRɳ�m���)�,�Eݠز��K|���X������2�**;2UAS�O$�܄tW�^pq�t�h��#�F]��:!E��@��y�)q�4��m H(�+#zQ1� /���[���}�?��N.{�U7U{���*��3���)k����ދ
���7�\~k!
��rg����Bl"��ƃ��ȥ�卵�q:�Ɩ`
�J_��}����c}���),O�gŰ���&i9)xmI��AV���)QR��W~�Rt#��-
�F���Hj���/��}�\u̥DL�x�#����#s6�/dU���w�r,4BQ���+gK���G-B�|gT�MPYEz$�H� �%���*n��ڰ�0�A��)��9F;˿�����H]3,&n�>�W[7\�����F�JI��� ���A�������m�*o�7}F�+l�����T������KSpw�{ΤAP�Zcd����BJ:C�S8��?Vς��p������+�	9�g�=��dkl'5Uh G��Hw�q�F��GS����
V�қ*�ѭ��^	'���iJ"�S͗�}��0��R��+��=��$�_���Ɗ���l��\���.VXN-�(�B���P�O�~��c��;(�wN;"������a]V���?�Ш�p���wۦ5��:c tC9SXp�['Y
�3K�^��m�fƓ=�*�_"�5l�=? =Zh�g��g]�zw氚����l2M���0�K���\��Z,���!��qؤA��4P��0%8'v�$�J�y�4�C��PS��i<��b�T��1,ԭʏjiAs3���x�PKJ(�X��m�e��D���j��LP�|��PT��9�]��K�%��(gp~������f顐<�Ѥ�K�?�l2����O���B����]4�j���ލ����p߹Oqz{מ"V~��ވ��2*�=c<�3\����<@�J
���6�����<^G���y�Z�KZ�1�6g��|����?�NW�s_g� O�ߊ��o�	�wՏ�&��#H:EkԠ�Fؽ��*�ԅ��E��I!o���#�7㹾�A�����tܟ�P ���+�ܻ��TD���F�\};h�ߢ�4�يn��
e����%~��C}�����O2�b���%D��9��9i�N�4��,.XmX���> �U*��<�h�u��.����Z����%�>�������x�
0�������=�^�`�h�Ѽ1Y]"��Jp��/Z�1H*<Rp"�������;���EiY(dO�؝g����/ �_0��v=,���f�"���rbVY{��[���	�=Z3,Jn1$�֔��N��BjI����S�?Z	m�λ��6 H5{!���8;���
Ϡ=Қc��mk�V-D�t�a��(����R?2L��{H��u�2�3똨0���8��|�_u����Kk��;D� ����L2a��&�26���{�H/MT�k���G�"P��Ҫ[��!5��(#w��1�r�,k�ϟ�IK�cm�(}3��h{����m%����N����stm�!`�|n.���^X�u��R��7�)���+\��F�*�JF�~|�����// �ꁂ{�����q*3,�X�@���׃ �2Ԣ%
��r:��n��i�����3���vHj<��ȹ��*�0!���k�E���ay�~Y��Cpqw8�hZ����k���qv�0f2j�A3i�˔�^��Tg&���#Nq�nYJ8���V�FPC/d���i؄B�	</�=b�A6��a�*�1E�m� =k'<�)Cas�Y�����
�lѪ�k����A���[X�]2��gP@3�5��������@��{rpW6K�魭/�lQD��<Dc��):\'/�:{�&�!�~��g@D�$��p�#.�A�x��IXL\=��������6�����9����e!�$.�~U�F�z/�9��/)���]		l�(��a�Z7@�{.�̎�b��FP���m�I����lG\b�� ��h�g'�z Z��1�������ϻ�9�����D��ˇb9d�J�b�D��jc)B�G찤RKW����XO�<�p	Z����#0q�{6!�ã�*�8R�U��S�=���/�()��S��/L.�@��;�+��+�N񘜶N�<�%|���B��L��"�g�܁�gf	�7�K�FAY-��_gJ�|��ͦ� ;��g3Tn��v,8�<%���*r��W�O'5��aw��&��<�B����J�F�5�=ܴ��G~�èڿ#7�Q"����(2�YJ�D�R�k�N>pB+W�f�Ĭ+ڪ�J?sN��u�*߫�`�t�J�#A���Ynr�zG)���+�v3�1�|��%�{/`Mľ<h�~i0�(	��@��]�>����sSK�-�R��T�E�!�\�V'�����a�1܂��:9���Z�b9�`����f�QX���mEhY�*x����o�b�d���h�ugN򛮯ow'�y��(����
�7+j$pQЩ�d􌮒%�u����3����a�_�a��]�0����`�9����T����~$��f�� �*y��uҹP�2���R�WOѸɟ���4zɞ.��38�8�u4����*^r��z�^�����F�9�l?�m�����>�"�[%3�h��x�a{�eE+O:8H:a�4ޣ9�/!Ue�����|i���<���&�&�E�.�Eܠ�v<D&qu�mg�Z'~.i����J�k*���lߥ�ɭA����٤���5G�?ֲ��_��Q�}!%�
�����ou�?�ۄ����5FiY6"Ήe�����n�>��I���r�&�+چ�5��p��T�C��<��d�u�8���(�H����(4�5-Ĳ�FGe���<"�-��H��VA�|Ì���>��a���u`��#5 ��܃&U�1�HH��R6%�MzL!H�)<j-��}�I��h����1	a<Qhe���rM��F���=�bD:�*	7�����<�@���J�"�q�����B�tC�yp`r���G�5C��?���4���O��׈WD�N��Dk�J;RP�r+��@&鉊> `���f����G@���T�>e�7A��	&&����sb�9�HX�����6W��N�"a��`A���^��oe�c�Ɣ�-�}�{H�X�v�EN�N��ʹ���O+˝/��؇����^2�;5�؛
^}7́�˾���/�W��:rq\�΁7����W�@���K�S��_"�A���D8�|�gKȕ�h��2Ǌڠ���,��<��z�H��uW��K������P�6��w!'`����m�c��kӔ3q�
��t�}-~�m{������Z�@��h:�Ӥ.h�,d>s���P<$��	B�T>�ɒP!T�o�Rl\���V�}�� ڍn���s�8��[0Ҍ�ңز�*D!񫳸�-��=+����Trf�?�����`z��b�����H����%�ݷ���_�q�qں~ņ��$�;!�۾�������|�+�ə $YZ��m˝.b�2����9.;"Diɭ5P��nDF2�0s��RњHל&�P�t{W�4`����7e��K
i
�&�@�v�p1ٳ��Я�����	J�$��"�,���r7�]��[�8�\ӛ���+��J����.㭧˚����([�+�X�ӱ��ߊ�v���[6��y+�\��ё�mmN�����z�z�)����M�����d�xPǍ���2���T�.f����L��i���|�9�@0�H�k���.����M
zpW�����>T�;=8�$B8�N�Un��Fc	���y����LϠ/�Y&�� �s��`�Y��w�X�|�w�R5������@ɺ:�M����i4Ȯ�`k$NF��q|��e���6*#�F|�u���ktȃK�:��r���$_Ml�o�%������ܹ�Q��T^:̍�7~\�l�X�����Y�h�7|D��)�B�9�p�"/�z�����]�K�|��Q��ޜm 0�:��'�O:��WI������z�?���
��X��!���U�o��,�sPO��},�=�N�훠썝�4�}��b�s�4+��p��=o�!CUio��O:�����q�}�XꧭHC2����7���]��cpH��U�8E/��xɳ�2?2{��=HK�E�0H�/�� Q�eI��J�!�:}}<��H��vI���m�C� ߐ������'!�����EM���dԌ�� ���h���n�b��R�X��������M�]�Y�0�f���*�2�N����|��h֛��K
�k�[�P���c:�3I�K��"*�ߜ���p�������;�^Q
�6�W��bְ�6���U�T���S������$��ߣ:�#�J��6f�d� .�2S-��{:c}cZ�L֗��)ͷ�jghڕD�ղ~��_�xZpzz�m��6d�%�|�^�`d����N��&�xD_�!�[r��7�̸!��y:��!��.�#g�;�~'�]/UB���]��w�+5#��IĹ��~޴l:��`��Al��d@�>�Q����؟���G�e �Hb&�!\z�t��X��}��F���I�>6m�!��[o�)E.ƹ�Jke����|���BǷ��:J%��u(��+��fH�t(��s�'{�HE-�|\�����4f3n�V~?�kć3�S����S�olT����&��3�i�3�K�0'Q��TP����g�j�wH}^	��%�T�Xj��B��Sn[�aEA{F�f���d����N�^�ŊQ��3Ĉ;T�l$I�x�?�d����@�۝^*��Z+����[�%�`��� y�����Mß���\��,���R'��Xcu3�&�6!٦j9�d����3q��L�?H��a����'cI�$h ��G����6|��T����~��85ob����[��OkS �r��h�*�F��襇Ռ m�Z����s]@��S��LĿ�&N�� 3	c踂s��_M�����C y&R��U������^��SJ�J< M�0F��Y0L���c��l�p(�:�c�O6-��	��a�r���]�˱���2�\o�?>፺h�Jg���ڇ�cu�&r��O�R)رR(���Q��K�C
_f�W"��kY�f�5j��J�s����QiS$rࠠ�i�}r#T|�fT�d@���S��N��{κN��u�D%ZЄm�s�ю���Q�Z����X��O�L��V�i��̞�[J Ο E�g���G���&;�Xߔ8�6ݕ�8�6T�B<)ư���W�`�J��*鶒4�g�K(��\�����ŀR�����Zk�U��z3��Ѿu�4���"jK�\�h�'̓4	��ۺQ�qL(��g�6:ز�K��.Ϲ��Bg����.X[M���Q%@TV����-&�9� �F����x�૪
���Ȟ�.}������S�(s��sht��kO �sXį�0�t�Z�Ӗ�V[�8$F� �1$��ʓ�;\���·Si�p��i;!�T�9جU?�8]��E�4���2�]Ă������>}�-K���W$}%g]s���g��@���^�݌�t����NO�㒬4���
����b��M\�CMGn��'k��y� "�<bD��ʌñ��O(�{��=��c�OY�,5Q`G��7���szB�S�����^��P��Wo���>Vz(�����#˟�<��n�mx��0�F��.�ۡ!a隖n�������~1��YV��U�;c��GL��8��s��K"��W���\��y�X�y�'��1~i��'/Xz�J�U�R:�k��o�_@����1�Iik�iϺ�q
��}S��l59_�|�c�i����P�L�%@d��M*��n�Z�f.^J/Vu��V<4�j�l@�B�>ki)zF#�vP.sd�-E
��+��S/�W��������2DH���\^P�K����J�Xr���C�#�����/��f�r���ڵ���gm^6��.~��d�XyUJ��_����û�m��7^<�������_�����r\}	ISC������%^��{���-�9�FX �w���4��D�z_�� ���$<J%��6,y=��4EoT�dqsV͔Xj��"|���t}4���̗���;5T_}�+Br��r���6���Ⱦ/�㔎�u�#X2'�)�U�-��${:D��'��>c���|F�ǩ0�Ս؆i�i���W��yb�S���FƼ����;o����tݣ�(�g��Wa����8���I���&�z6�@6���_L�`.��j���s��:���i_�}\���tU4���t�5c�eG��':x���!Ҏ�A(�3��W9���/EO����R&��7 ����㖉����J=��y:ɖ�PLr��\�5Ƴv�6V���J�󐝮7&��r��@n *Uz+i�ZPs���C1�ã���&����ڵ���"�
>�c��9ji���kn1K�F����7�N�"Ds�Ґ3Ze�1�@�C����������U�sL���r��"7�}��f��Ig�'���\SH�Kh�d�f��!>����p��-�!�R�{�iE/o(�d��Ǻ6A��"�T�430g��t�X�
Q�b�`yƊ����.�֔�+q�^�Ta����MZ�L����FB�0G?�7�_�c�����V�y�L�s>t�3��[��ܭ�J~,�X�F�+s,j���ïv{'��Ζ��F{-��\�N�G̓�C�Kj�3�H\�%}�Oa`�.z@1��
��γtƴ9�yĂ+��R�Z��G�/)/I�.�c�x1�L��)��9�lQU�u�p�z.�2܇�yCdtű�k�\����[�?}����U�g+!=�f�[�Lh�G�rf]�+-��rfT��M���PuP�{�8$ �K2���8�����Ɯ�is��q�Ȇ anX�j�Us�����d��gx9b��ݯx��X4kR�c[����U�u�W���q*yc�Ӓ�sn��E�'�­����ed@��U�>wV�hכ�$���`�'�`�y��G��w�g2F�\H�@1�~�团�5 �Eɩ��b����V�Z8��E��j��"��\f��;?��dz�f���;�ԉ5��,VC�w��a=�EH��%FgM����]+����[��F>�:I���!�-䊕w�Adc�
��f/��=O��8���c���Q��\�����K��L"}��	�������Ac��.���L�R����E�ȔI�uE/�5�0���RO����>�=��g�@Z�SE�Q�uɑ�`3;U>�Ѿ9[��?�Qoh?��]��e�"�y�w�pJFJD��R���d�,%�x���X���J�= �yҵ4bL�LJ] I��0x���*��� f�oQ t��0� 5�v�����2CPf{���r1��b�D;�*��.<�jG��0�'�-���]R��!$��D;�Fｨ3�I����-�迉��ڒ_s˪�P!oI�^B�L�-���{lT� ����h㉜|�C\�CJ*%���q"�޵lh�!���;�1�b4!��#F��L�*ʃ:�A\�Nz$i��~�\cϹ?�L�.�{� ��Ӑ9��!��M�q�aEfp��P�z?���N�5���⃦����޷j<�x�@�Y���v�������D���O��ﺷF�/������`(���}������F�f^g�%��`ܮ���ȯ?1�3�5o˟PN�����'� o��������x`�t	����B1MD�v���!�0R��:evq5�t{�FX9 ְ`��(�.�&|�_����;sy��ɹ���rI��XU�v4�O�b6�n����ʓ�(JM}m�z#�Nm�	�v�*���o�	o_M	�(�əo���rD; �>�G��j�zuBa�V�%�kl�o��1g���?�a�t����:lȸw����ԏ��e��Tܒ�����`�0qX�k�c���C�˽|*�[crbG�P~l>�щ���q�VG��`*_/���@O�˹����u�ډ6O�ے���{�R�?�"�@�
}6�C�0p�_���f��gG�2��I ����V���H;�L����br�T A�(( _��jl�����)S'�0q,�w�>y�[���e(��쑜k�H�����[��K}����n��s�
E�P����\�'MOHDvI���ze�'�ϝ9�t�e[�E'�g`�(�-?�8�æ�ڲ!���E>fӓ�k��x�/r�i�}:�'h��_�sZ[�bAQ/~�j(F�Bz{an��>��-aL����6X����q��#���'��I{�a�"#5b�n�W06Ǐ>�l|���M.�@xF0��SP�M����D�z<�_E����FEb�ڙ
,X~g�����@p�����d>
�A:#��E�{�����S�'����i�"�~�)�K�	��Rx�������Ǿ}e����!Tp_���w�n�bA���E?���]��g=/�� � ��2h��������z��I1^�l��gw�j-#"Fj��@iV�e���Nj����_�W�'����2���X'����2R�ky1d��÷XP"��jW����'")ǂG�IIj��KX�ѡ[I�R�|r��TS'"���`~/H1��j)T��*y��H�C��oޘTf;�HlC���R�`bl�C�yZϹ�\�2C��,S�<�^�6���SW� �ezC-���f�ޗR�o_$�1b������߸n�O;�yBW�Ԥ a� y�q�<̏������Ϙ����'���	RH�mp��T�a׻#��~�#���A�:M%�E�(*�h�i5Z��l�2��55N�}���'�,���c��hU8t�۩�Km8L����e6㾃f"���P7�Zu�-Hx��x?�Ŀze&���c���+0�	���5�q�V�G%{ϴEM�Y��֌����[��&5��iaf˛Ҹ���k�KRC�	�&�2�MKS��� ^S�ضF��K�zN�X>�����&�i��߲B�R�����L�����*ם�B��\�	��X\�ke��=�>���p��9�F'{�]����ф�L�J�=@�s��[�*�W��[U�n�����A;,�UI Mj`.��������^���I�Nb\�s{G�/ϾnQ���^B�&-�Ml�vk�����`�Dv2,��o�'�Tx�$�p��4o��2��盆N�,�A~F�K�j�ؽ�T|j���H5M��%6�	��J&�"~�m��(�����������A|�@MRI������\I����c�5�	�ɠ�ũ��\2�C��Zx�pS�2���|ƾ�5 ��54��>�ΠG�`�����2�(�y9iҞ\��x)q��D�
�}�܏�-��BS�V����Ԡ�M�ߐQ�4��A�����˓���������4�����]�i�k�<����z������J�jU���r^2ل2Ac����c*x#���ń�=3��G�H�s����GNE�$��ʽ��g�r����m��5n�X��2_K�����z���m����%b8Ti�t�	�7�Sj� +���<TE�a���2����?�n]�,wL|�>X�9f����3j ���w�)���)=���_߈�4b��EE��Q2��G(��mbu:xe�-V���q���
�I�	����ҍ�#�Վ[�u1L�s��!(�bw#5���4GK��EƊ�M��W�fw���J}Mt o6��Y0 mZ�Sm�
����t*��g¶=������Y�c>�bS^�1��wU����^^]:P������p�R�"�?��{���ͧ�aj#���k�kSeI,3���Gκ�B�.׉�8Q�z�������B�<|��:��UV�>F�������2���0b]!���d�	�4�F�Gm�=K2<�{�
��!E[�MQ2"\�ב2`�NM�fL�l�/�d�(c#Rn�˔F��HD��)U>�I?aV�o���,�ǐ�5���M�p��[�%Pr��>�C�& ��;����o�h�r�i���p�7ˁcT:��+���!�@%��VXo ��:��sR���� ضW.z���� �f�w��j������s۸\L )>�@���;�@�m��6�(˾��h����\R�z�F6��L�x%��cC�ډ���0)X�P�3,=i#��.�5�}�͵o@�C&ۡ7Eu	�x����9?� ��F{�e�Pw�+<K�>��Ak�XJ�gl6���퇨(Np9�˻x5r���
��|4����+��u�����Kt:�q�\�����5Ĩ�9��+�E��*G[��TuE�b[��Z�h�a�,�<�o�I�Ι���>Μ�*��,�b��������s���i+$�8��X`a���a�����uv5}/RփPŪ���SH�1c��f�0��N�����LD$ɤ��4�|�%���g�܌_�y�Qx䭾Ү{�̪n�s��7|�c G7��(X���stˁ=�<RL��L�vD1ȿB =/P�(����������
������#�t���J���y�߱Sc�Y��Ղ�J	�1�_��'�bK�ˎ���M�����#�&�@�"y3pX��</S�
r�����W#�8�2�����PKUR�nv����}!*�ۚ*l�g06Ҩ�d�A� e N�ʆ����m����4��y��n����@x�
z��hFq��++��3{s��=���1=,�?�X�I��t0��,�G�����K�?�⿽��v`B��c�#z#ڪj3�Vqv��Οnb�|@�@09e����u�>��T�i��S;n��OMF
�v�W3�A$(���jX,t5z��̐�^wQ�j�Ysrаիt�" =YK��P�w��:���HY����'0K�S9��A�|�/��a<�2���.�$8"b�j컋>E	�:�R��k��9�ƨU��O���`\���
��4�+MCQ�u�S7(������(;�1_i��No3"^5�N$EP�����g�X�h&m�%22���t3����������>,�ū�2EH2a�>hT~q�VDsLv:���������#��/(����q�Z�A$��H����gҊ�v�zUH1����À�:(�tn�]���p��p�D��Xi��r�t����V�ň_]zĠ��;GQ�!u"���.t������߳!��t�"��T8�w�҃�`�JXWw��n렻��8��GQc��Rq�םq@z���S�!/v\.O꼙s#�vN��<�lzLkq�yWuP\~��%�pG�Ƈgdz���\�?�rH������e���k�-Y�����Ҵ3&�5�V�Y]�֓M咮(��a�j�;|���J����I�r�ϼ`^v��&�%��%3�|'�=*�?��a�!��l�$�~�������?�D�R�H]q�@�3�/�ڀ��R�<��YPϩ����������Ow8�N�������K�.�l1�S��WIkl�x�6v+��^M�SC3,o�Ϸ�:E����yd��7h�?�v�{��m����`���f���)�(�j�I�C��9��+��50��l]���Ea��wKyX��h�$బ^ǆ|pf�+2G��6b��N�b��h*��׏��r!�NǮ��1%/��9I�3v|��i12�Wb�������q�k��E�7��m ^���R��Vқ��i�HR�V�W�"����e�R�����R�72�2@6�y�)�Ffd��(���$�:�G[�Ʌ]�;�X����>	���:Kˊ����qH����02�VD&>��S��Ќ6k��K���7�<� ���O�x�\0�t}���(S�A��Ad��[�irI?��%����%R´�M2���5�@N[����֙3ӝ�� �y�ں��Y��,Q�U��V�� 9�� �l,tP���ka�|�Jd�l��Z轸?����ư��E�K�q,t���o`w+8��+�[�ڕe��>Y�"��1.y��A���GNP�_?�j��Bg�><ؗ���~3��0U�]��*��� �b��W���SP�nE�~��L	ӕEy)�;�33�a��P.'z�ȱF�qn<Ϲ<;H}tlt�{�ߟ3]�>���uU�k0Ym+`�@J�Ī�L%��u�P���≙UdD���{c`�f��U憅:[.:�BS��j(1B�S��\���A�u1�����ui�.D0��s͋�!de=,$%;����G��!�C��66��9r�<�:��S~�%o����pdRx���@7��P>C��zq-�j������FѷY��p`%b��߉Ρ����TmϠ�1}�^�E�F������ݍb+J6-�>���<Qy�.�g)���<������k�|Ȝ�w������6$��t�<�qH��w<��������V�$�g⷟��t��{��G��}���b,��;��t��^����~�2pִ�S�)�ѪV����+�lΈ�B5T+Gxu�˱��+>��-k+�h�*���r(��ӟ�-�!�F<l�t�<����Ǹ G:V��H~���b`�;�G��ɬ}�8�<��m�#�;�P��7������p����ޅn��o˒���A����XV&�ފ1��_є��9���'
�Elh��iQ���Ų��2�;����^�fOf��ζ9З��;.�L�*�bZ�v7�a����l�Є��?X$c�[�4���L���Z��*4�$��ݻ��o,���N/�:W�o�2����|b��9s���ت�g��]��R��f3y� 0���|�χ��'�@� [�Ư�W���J��[���h �vpc`�����Zpm�~�V��uc�ȭ��$uz� �!�n�P���L~��
�7�W���{;�ҕ^��{�|��K��fmG	���w�&���"�����S�c�'�Lx͡*֡z,�{D3�gÚ�8&x~�''���o�`��O�.=�h�"��Y�f�W���U�.���%Đw�!6DE�O��̝�z��)\5�-�fs�#8�C�xh��f�����F����&�@1V�仆9 ���?�uF�-�����:f~=�U�&=4M��@Iva8	�&a1���H'�Qd%
�ʯ�8�η%+;�jt�d*�����G�����R�#'���*�^.�\Br�c�7�q�)���h�B񤊱�1t������=f���tô���Yr1���(�T���2_s�ѳ&'�`�&.{� ��c�a����4O��8q������xwU�"ڎ�MP� ˚�|%�zX⎄�k�����/��i5�������	�Y��L�/�J�w�m|�n=y�aR�Sv�7�鴝�rkp�"Ԩc���#���7zbM��w�؁�2� R����M���b擄ni,�^?�>�yNG� Gs������U��Zܺ�*�������,�Ǚ�
ۀ�T�`��_S Vx�$� �T���iI��]x�!����Պ�O�2�̣�أ��,[,�G����p^{,�����es ��8�@�q�Mu�h��kϺ,����!������t!�ߵ<��ev�u��O����Г�2	7,���y�ۚ���6�V��a�:Ǹ@u��r���~Q/�/����b��4X\]E���-�[C_B~kE�/M?3�p&���C��p�M�TDe\���d�LT�p&�^�4�)=~���){���w����.z�������	_���sbEt�<^�R�/0!b{��Q,C�*��+�ȳ]���$�$�K�C�I�mK�ߙlQ���z{,���/��9���C����$y�*|J�yG��dV���� 5��V�s'�Ӟ�I��|}>��Tclx��EτU�W\��Q�zd�G,ʫ�-�3�wK���]$�0���)G����3_0F~SQ%[έ�����퓇!�k�'�Տ�Ke����9hB~#<d��;�EP
g���/� �L���E%���u'�(b?��<Eh�u�N� ��_z�:2��&}�B����� �舼/,��w�4N�-�>�S���h��xGBS� �SCo�%�F����:���#�(��(� E�O^�6�r��Z���&Q�;&|�0�3Xy%���r������ˋ]o��џ�z;G�����G3ҙ���4a�1�M�`��2���d�F4�'҅�]���p��`������ �X���)ʈ�	�J��'�����֤/.(y�h9���9]��&���`el	U�Y{K���ǪBY��D��[;�|`�D�A�`� ��~��<�\����%%H-l6-�@P�ؾyf/Ǡ���:�X>�E�2��(��j*��~���^��ѷ����㴀�k�2�"V�5ў��jl0�a�����ke#9�0ij�zN�V�s�3>�U�3W];FE�9�'��p�˽b�{9.��06v0�VT��h�9z	�$J�F�9r<�W�Ʊ�fQ���W���۔`CȖ��-���)���ڏ�q�{�ƻn��I���~@ִ�a!x���6�c#�:���f�ԽE�k�(3Y��΅�G/kb��n��R��5��%�ϔ�ܱ�&f�.�!CCe��_.�l�D�*�bU<�[�-����z��wxՠe�w��$K�������׫h����5�:P�(��w�#����w0��^��/,�캝��I�Á�5�$��`BZr螟����im�qG�2����
 �ҫ<����ap{�U�#��s��Ae_�`��%�6���C�����`�
�P;�L؛.4�"�7�]B=�GĮl��V����y�7�/}K��$�nx~�X���p��(�������p~8+���,�}e�׸��٭F`��Vbg��\�I������1�³�~G�jJ������'�ng�����X�#xҭ��n+��)����̜2H|~�*b^���BPU�$駻)nI�����w�}ņWr,g��˼��
��bї��}E�-�k���c��K��� ��=f�DJ��;h>�r��F�9D�+�K��s乤Y��"l-�/Vy4����+_�ʀV�b���[w�h���@7�C�w,W��a�$V1��/	xe|Ɠ^w�$,H�~����J*es��	,q�~Yc�����K��mT8{��.u^�P΋/��>Y�~��M]�K[gE�����F:YJ}i33\)'4e,|tnG�^��S�t�w#1�ht�>�d̹�ADHVu����\X�ĂbM�wq;�|7�~uc �_�jF�f�P�ܫ
*o�̲�)�Li=R���_*pՁUp�tb0`��mm�=5 ���bvy	�F�T��
��~n��[�E$
%��2�.�(7�a�`�͜�JZ��t�u��p!�}�_J�f(�n^�eHC���bm��N�_'r����Fˈsx;�C"x8Ic߆,��L���������`�No�nw��Sg�L���u�&\�>j�O�_(��1L�0���I�
l٢���)<F�@6emw��S���e���=T%:6�-�3j��vh"���BV�	�U�o;� ���	=�#.�m�7喚Q���q���UA��94M���W@�(�\,(��clv���Qn?=�yr+�
0Fg�;�XB���ۣ��u�f��)m9�Z
^<�����Il���jE�Fxi�1�8�$#F�/�0&���]�
���#��8��A0�Ѣ'_�ëE�5�F���>��f:c"I]���z|��,��v٧��&-��f �{x3�}��1��^��p�"���w���g��H�FРL˯D�3_�b��o�{���|���z�������k���[!��q��L�;OL�WY��
]6�tB�a��}'t� �������/�)���/8'�9+�`@��@�d�-�/>۵>����C0EEx�zfI�Q����l��S&1�����k�R����>Y[�1r�^���� b��Ҥ@`�K����>��)��><�l�gRk�!C*�\��t��vT&��0��L�h�{�4�!?���X���_�}�S^��ܰE3���Lo����苃	�עZ3M}H��?aj?��k��^ӻq\���t]�vz�����P���!3M{��h�bg��^�L��>�\K5�������E�CsI�LyI0MP���\N*�/yڹ+Ɔ�g�E�;��>1:�M5��s��F�7_DM��R=�*]8�Io�_Y��3�I|���T�8B �SBJi�C(�;ڹC�*`ٽ@*q+I.��hY��I���]7c<t�Ԟ���d:�˳e�~]]�7���%��G���(�)�q���9iQty'�z���> �+�%�S���щ7�����\l ~��J���[�=s2(s��l-�଴�a��e�[H���Z�k5D� ��D\9V���^&����� �#Nཆ ���40���$3Y��$�5�z[w�U�ͶWpd$�S�J%��܅��Bj����E�ƫ���;��*E�* �a�Iy�C!�����ѼY�Td:Xp�[��}�ˑ:jکF�\\'��֭<��%U�VfgӧP0�	�ׯڼ�{��X��[���RO餃�UJDp�&�^ �q���J ڮ�ߖo�f�j@˪i��=}���8���{{)
��� N����2	��|��-YK~�B֝v�H(�&i���Q��vvT��(���`�_p��E�}�m&���l���G�$��'����Z�_tcϋ���
"�~�����r	/Of�n<v�C��˭zJ�ת�E1�	�(�Ы}vfa�Ǹ����A���?���B�x���~�?�tW��c�y��3��ǖ�3��N��<܀�N���=#���s��hVv�62$v�6���V��=�D�$?�|�t{�f<�)�]��k����X�vov\{��T�E�,��::�Y.�LSn;�L4��CF��[n�~��z�|��},Q����w���(��Y��_�-�	�����?�ʙ�(x	o��bU�v� ���Y��i��]�D�A���5�@��oNn�n+΢�l�明�1�D���t��8E˄��::��T�;�:��V��!R�N�DW@�yx&ɣ��ft���6���+��gd����8a�З>o���Ƞ�b�w�
�pU$Բ�b�_P�| ���ō[-�{��q��xn�A���Y�e`�0�1w��e�.�Gκ���u�(� �u�s,[re-:Ms�s��W��fn�Y����}V�jWA��_�%ll�='{�~c�������͂�Z�,��Q�U"�up�S	j+�90�嘪�@3�8�� �P4�Ꮃ�P� ��+���9׷����/�t�F��'��~��,��Qŝ&k%�y �Z($�6n/�.�
%=O���ո�u�4�d4h�N^K����������Ɣy�c,f�5p�'���~�tW����>ھ8b�T���l���'|�¿,1�M�D	�s�U=�Ǌ��.5X�b�b��Y��t%�D=2'^��崓*	sp���j"r ��3�@��$d Ɗ-g���rW��l�f�e�:��b�b�P�Qn#�N�ܷ���ASY�����=�*B!�"��0��p�7�C��Z<�]�E�����"��f�C#8+��W%溂�G5x+?�C�b��b��f��/6]��*�\*G,�] Cg��}��3I�袻k��^�(�ޒ�-pR�ì��)y�@L��';��4u_��wn�MR6r��M��t�=>Ş3#�NA���1!oS�kg�;gA$����@.���j{6g��.�2|��\ܢ��0ރ���c^�)Zf�ӴGf��u��P=N�ߗ���wς{ˇ�,{qʩ�=WLP�\+ӈ��'O� 5Cw�W�F.d��8]�)m�H�~7�x�E��X�p�Z�m+�*)�9�A?ܮԉ���Y���GOg����-ް;�l�%N���w�M��iA*!�h�\��p��`x��K�f�hrL.�63���ڲ�ZsR�88������n��Ċ�)v�%u�I��N@�
�,[H���z�WB(S,�zU(��&���
���zG$B�����0	w����N��\Hg��y�N�'�YI1����g��p6)�7�Pf�/˟3��k�g�
�܆=���S�tO㩃�*���A���	W��@�'-�i��e�`�U�
�0A��y�U�FC.Y5��$6� 7Z��nB#����~��Vo�Scc	��ڟ����2.{�B����u`�W48O�^������&����Y�jb&R80qU��\Z2{�Y�����l" G�#LA�PV������A;���JB�)��  �����p^����IrkeQ��F�M�����2���Y�2�;rR/�ؗdО�]�LC���+$��)!�g �N ʾ�IiZNI��$�p=���By˴���ER�-��M:\�3CdNe��V#����]9Aaa�L��1v��'�l��8��l��Ǌ���u��?i+mⳁ�(�)�\B����׸�ʧ������	�JYV:���s�W�|�c�0N�5��>��F����"�?9�������q�秐�!1��0^q�ɭ�k��>��xnp�}� �SqC.�CW�hɴ��{y���Ia�[�)m�f�8�V5A���g'���荲���!�1@�Y�G����m)w|�AtB¾B�R�c��~i�8������T��Z���=]^���8P�
:65ـ�}s|�V�΃�䧮��B����,xd�������#ү%�#��y������?��Y)�j@��������sl�3ܮ�w����G$��G�"=�8B�#��7��m	��-��)�['�I�mB�o��UWiH�X	;� J�^����`S���$��%����!��5b����b�eB�]d<*ʤϒ|[:��ݢ���)���K��5-i�%��&\�аB
��<[h�"kpCc���<&��a��dh�Wr���6L��r.Z�CyU7����5����VԹ��CBL8�z��� ��-4�o�������㖰�'�C����~�ٞ-D!_ �O~�a�ܟ�>���c%�sk���g��{g��!C�&ϑ��#\�[�A����1A_D�[3�6H��D"�c�jŸEs�:�{�Nn�V�����9�j1�?�[�`�ą5�>+�q`{ԙ�/"SSV��i[�K�u}.I�O����4!4&}!|�3X3e��[���s�zSe>֖�����A��ũ�V��4�VaW"�AoS��'r:Ze�F0�_˵�<�/�i�_���x�4w���� �X�3D��?W����g���hj7<F����>5
�<5T�i܀��6ת��NZ@W�ʅ��>\��}V����0Ŭ0[�P����M�\��řu=��i�*/W�!�&>��۸�y)6�X�V�O�	���#��(+���*ډ|XGߠ>��p������Ӟ�:�Qݣ}"�`cJ��o������d��/�f������ݘ4�h,ex����{K�����qR��v�2}��$əE��b���ʮ�&�(g8���A�g�����.T!��� ��w�ض.'���7�MI,�+����F	>e�V`#���n}D��&(qG�.2��m��,�w�;�=�~>dGS�i��q�l��[���2sT�S�+�}ч@��b.){͌e�  8���4�ު]Qя>dc����%R�0G��q�����;;t��(CfL�z^��l�h������f{�G�+�-�@��X�F���c�1b�Y$���F��L�N��!h|�A밞�q�N~v�*���tz����+?�"�V��9������Wun:��٭�Z�Skp��Q���~��]��i������:�s����D�=����w��+��bSè��։����������*НJF]��PCR���qb��d��lA-.-ƌ���ό�k?�,,��d��k2�:�S�߹`Sk�|j�i�5�W�q� ��2�����Px6M�M��%QZ˯�ߨ8d�����u��ã�f�ꀘEM�$��9)7ӥo�5c�#� qr������m0y��yZF��r�i�*9S�����j|bAi���Q�6qe����u�nW9gG������,�Ay�W>����i`���Vi�y�Ӌ�¥vR��a:�')�ǩ�>q����>;zb�N��Do��|�y��E�:c.�Z2��D���Vז!��`q�i'͛Py��L�r4��ڞ����Ieu3��N�W�O@��t��58�ܬ��O��Q��m���
9�6����[�xT���O`D�|�~��V�2P���Zӟ{�{�ջ�Ġ?�10���5{K�w�jB��&<q���{���ej��AO��J��sG��;�[�����mS�ˈy�u"�����,}�º��<2��y�͎�b4�=����n�y;�ޠ�U8�&z�{��x^R�O���q��~c���{ �<�����q5��8�e��R�+��L�+=J�^z(��9��}������b6+�8iF���ԃ�H�%P=;.�.�c>6�_k8�ԫ��P��v�g��%}rS�MS�[�X�3�i��M,���C�����l�w�U�� \Xf�0T?��?�k;�G�Vqi��.��f���N���qK:S�+�Yx+��^'e� �[���0�>-�v�5V8�G�sa�����w)ST��>~t*E��dA�3j��D�u��D��6V$I��p��f�^�`������������4��8xN��AĆ���4�P���U��4#v����3��J�E�� ���}[bU?��������Id�����EWMD�%e�Dj�Y�`�XZ3e�:�7�}o\uT��M�s2�p��t��C^9ǖ�������Ruop�8����_:�\����KP�'8���
Z.Ŧ��\#��*R͌����tB%�?�Ņ	X)�x]�d`��5PK`�!S�\��F�l�G�\�1��y��ZF�y-���<�=c{��"��V��ӽH	�����M}��L���4�Q��@��É�ZФ�&T�cc�w�A��#���V3�v�+(v]o'�P��~�fU;���SbDSO�T���.�U���|�$OO/I���i"rY=�� IU�����]#�'�l���+�e�3�4���v�{�lo�Ѓŀ����!�v(,�)7R>���6��\}�~L�I2��d9e��@�=�YnF4N��ڇ0�;�ARE�WE})���iA��O�����b@�nLȿ��Ak�u�}���{֜���Z$"�<���i�x~�g��q�(��������rx5�����n|;$5��M��IW*��A^�25���i�g ��%|6��\H�g�z���#�0	3s�����
S��!�������QjB�ۇ���8���h�Vs���5��K���"u1|5ނ��2H��-�H�F�&�x���T�r�*���� ��ی)�)u'�o���[�� <f������Y$��CER��h5!�����]���䄃�p��̐ic�Ua�Cf��jڹ��F�?�,��g$"Ad��	��:��.��ڲ*.�ӕD-Y�@Qڗ����Upa������v/ʭ�".>j���ʘIs8��3Q��*d���.��IŸ��X�k��$N,s�;��#������)��jR�",�-��nBe�X2����J���) nޑ���f���W��۱K\'{��Ѥ6����'
�H+Ylh.�Z�Զ	�"�T�X|�[�lk�����!	�L$N2�ؖ�O
.��_-c���G'ܷ��M���B�u+��q�s#�H�+zøj���Q���Աc�������p�}tO^�]�DQ�0�2a6�w��>Y9٩U�d�����)/���_��ݦDU[�<�O�04���J�q%�IM+�π�)�Η-�����6���s����O%��邢�υ��Xê��-y�Z[�MVܚ���n���Ė8Et,�Q�p���=�M-#�t֍���?�[�0���lseU$�3��9N��
k�r�EQ���N���î���W��KJ����i�dQ�bv�X�����4��߱����h$��d�/-i�h4Ok���_��x";���i��q���8��y�����*�X�S��3��qf����� �����)wt�3ʵn=~ٱ/��Ƅ��5oQ��:e�7��.�	�|�*��n稕�S��m$D�LNGzC��Ν�D>0Ӫ�y54�n�:
b��KN�\m@��C�Q�����+`ң���\+�0
�y4ݎ\���%�sFy�f�c����d�9MWn+&��1����)w�v�$X���8c���X�HMVwO���5v
�a�'wj�2ۖ�w�I0�s�<�}	�������Y�\#Ȇ"W��W���w�b��ka� ��M5��徆�6�S�<]�cn7��9wi��ި1��r>��ɛ� �)+D�Tm�3�o����5�hb�$�p�����y�S�A8|��A�:t��Z>�s�aM�~��������n��;x?��)�!3+"ap�3(�IIc����4���'����([�h���ֳ�ҬiV��͂&���`��]��t#MSQ�j47��!T;���~�M���Sco�\�v���<�Kݞ�D��ɓ8�b2�cՑ�b��Ǜ^��(��3�	$p^�ai7�9� '�;{�����-�#\Z2����3�D�R p�J�e9��#���S
v]J���n
C���E�dN�3�&�=vDɤ&Y8�~�1&k�u�നص'�a��sh~��m\z�_���\�J��?���4*1�p��5���n�>�gu�m~��0P���t��:�
���	����(i�6�L8DC��E�]���w����V`2�f8�T�ˢ�����[��T6n�5��4�7���F�6� V�6�s����I���/�����6����V��*�
�9%86H��u�r����u�+l�c����0&0�]�o��ͬܬ�mP���o��%���� `4��1Ȳ�Gm�G&_��7E2���>���9"��ty���Dˣ`"c�YH1�����{�f<����Z�M�<�ᗻ��E�%�����-x�QJ]��u80w��4dlt�P�C��W��I]��׍����䟑Vjo��� �m�.����l�n8s#?k����T�����t�t�� �������4	�B,�7���7�Z��<��	��	�w�Ϩ�hWe��6ۈ�1F[ǖe� ۾׷ʋ���N\pch;s�R��t�.�$�
�� =��~�L� ��*�
}UO�Ӣry��X��VI��o���7��!�F�MX��>�?�,�E|�n@��>��W����3���LX�9��m�}���,ܶ��w����C{2,��۶���*ndRb���[`�I����<u�[u_�.�����n<"���'3���X�G�wnٰ��l��c�H�I:�~:������*�_�����=o�`ק��r��� @>�[=�ň,�%�Z����@r�_i5����q����xf�?-����j��I��݊K��4���X/-���d���t�#��j�k���e%�W@E��r�vA�P����� ��#_9�jA�5���9&�װ��\'6����2b=�����]�. x�0:�Y& .��R�����~)�{T:��b
�r8�u ���!x��mQ�چ�y��"��\��Y[�$];��'C��}R���Ǻr=���������y���0&�Np��}��Ы�������>��=�@^S��|~(o
<£~��n�p��ۻ"���p�N1��PN�EW��1��8��G���)~�_������QW��?B5� ��T.�"�3qAN������x_V�h��2���QL����8��}d�'��sJ�X��Jk7�.�QU[�f�֞b^�����B\D�.r����INp�U;��T��>r<�!�-d�dm��[_�T<�$o���(��jИ�2�����R���P�?��ӥ�6{�J��x�6��8;?�| ��/K��+�vyH�<dg���ۄ�E���f�A/���6�x������q|���Na�T��b�rHZ]j1r��Z�X���b��HE`*�����Y�h:��mC�&�[�l�=��	i����F�VM����N�x�����(;��w�#��UzT��1�W�X����^+'����3��E9�{q��Ҙ��9���D5�����6�^�Ө�=tqާ����RV�,���R�n0�Y�Ӕf�!r�*�w�8�\JȫlP�\j��+k֜���Jg� `�^n�;:A��R�g���۷��H�)�V�T��W��@!�W�i�$U��U* ��{y�|0�6�\�O=cyg@�����錰%aCC@����7!�M? @z��-�P� ��$"�S(Vs;¬��N�J^�����v�p��%V:����8����b��"E�"Lt�ڇ�Bb�z��Y{�a;BR;�/��g���=&,0��N_�w��f$a����	'$а��/��	�S�\jL�3 �#�ab�����Kw���Bm����×t�:���`���#�{�����6u��=�����(����j=�~Ubq�C��2����Wב.l��7�|h��k��U��$�Ϲ�V�����
�C�����+�"�7:<����-I
�Oo{B�<��^cɹ(��֢�`��<�;�D�<;׹���pV�������p��T�K烻��"*��rd��	���h�Uޤ�3Shݿ����ex��c��}�o�����u8��������:EnWm�\7~�>��e��RuR99��W��;�J0БD���e�NV�}����!�>%T�ϵ�����ݪNG�_��ܜͮ����X�ϵJ�*�$0��G���5�)��e��:0U�	/n��B��WS"ͭ�9�19-#��:�0�߆�&G'	��6a�e��,2i���p��A��A+f|�0#ʨ��V��B��F�S��-�Ė�DB|�ϯj�I�=��se�L���F�$���œB�������MY0��G�/�,N�H�&�uQD��s�B���wI�m�su�����ݰ1I�P���Q�bC:�Qg	�G�
?���I��?,�w�I�3�#�ck���iT�ұ�G@\=��IWaT��uA��+jxN�9�*E(G�]������G���$�ma�ޢ�9�����6j2��Ca�i���j��1v$��Κ�HH{�+Y��˛��n��t�;~��7�pΑ�ՁO/9�[V��7
��?N���DAsi�Qu�J��ݣVT�ϓ�*���bx,�}��k�4^5�9^�I�ui�c����i��ɋ��a 
�`o��4?���7��T�t5n�c�76!��kn]r��m։|�_�j��=�a����@�ēb��Gj�N�
�x���t'vE�$��p�[����-5�|���Z��8L�)RjK�G��ög���x6Sg�w�o���9p���3^{�[ES��/�v�EK�?H�Za��0Su��y��BG���`ߠ�#k�1: �T�t}׶�Ǫ�^�P���6��N���A�"��B�fTJC��� ���V���vM�<b�"�~�][�����*?��۔��� �^E9����a�^V��&0T��R���4�=ƥ��l��g�4g���
�g�ʁ����b?�j����(�������E]�Q���I�IЩGu���<����(e�>9��G�Fi�� Z�W;y���ra�����E��p"=�TRn@y9���'��rT��_�T��]���0tbg�O��T����}q^�k?A>����b���9�H�L��3�g�:�}_�@��/e�W�"��<c�磖�ru��Bl�H_���
���>�*�ڴ�
:�����ˑ0�m��U���E{��n��,RY^\��?f�T�����إnz}��Ļ�~��u�KT֯SU;����.E�,y�(!�ϯ�G�?!�su|��|��a���ٶ�&%£I�C���,xpZa��Iy-lP$����|Yܫ=i�y��|�+^�z���R����Q~�H��e��+`���<��p�ڈD$yO����xe����H��*NH[��ğVh�u?��:_���/Dľ�j�fV)��h��<]�n�U���Blыx��.*��?�nv
4��M��M+����m+f�X}��p��Hq:�m6���oS�w�=!]x���V\����m:��4�p�z�!�B�#������bN
��3l�g����E�����J�gg3���׃�)Ɖl�����=���]?�c�7c1����!qa�ɀ-[��٧��$ϸ�1o�"M�ZGsNa4�Y����+Tj�W
Su~p�7�$��9H�D$�X.�E�����j���Y1ǫ��|��2|j@�#$/��HOͰ�ϦR��fg��W��ı�j,ϖYT��E���w�J�0:���z�XWANb�����]t���3���|�ڻ��s��G	�;���g�O�hp�tt���4G�����h�eG�Jq(�Zś@ZX�Q��32�[�b�:������`*{�<�ۻ��Y���X+]Zg�<x�4�kX���j����R�.w�Ŗ��S�5f�ҶM ;�6?�ٺ�A{�a-�8�;a�w���y8y�`C:�-ݶZ��ԁ���ZKC�HL�E^v�I���?���egu��h�u�*�D/�����i�K}�f�7�_�|s$��Z�Z�%^&��c)T�_ �U��	M�x�$cI=�F�3!�u`�Yt�ωX��aC7	_�nQ	ME���1=�(s
6��F��#6;Q��c�p�bi�F�!}LT���6������>�ض���%�$:����b6:�O�AN�%�p`ޠ�-�=�JvD�.�c�*S��e��nLW��8��ARy
$�~�`�tZ'T��lbeGGS=)���'�M�֮d����,����Y^�����a\��Ȗ
�8˨���jZ-���<C�f��Oɢ`Ɩ.b��F��̧�_�R�Z�|�ش��ڃ�r�)�.+��آ.���exk��0�}�?�[�a��t�������wQȕZڦ��?o�I���:{)��9�Φ]�8#�d���l�6.> 9Ws�`������>�.�?�^���˨®m�O���3<ߋ=E*����Ԃ2,,�H�վ>z�n}�����9%�K�W*�j��Ի��`N�&���(��_c����`�ʬ����_O\B�Ͽ���X��Ӽ�����#�X0/8RJ����D̢��Ă`�X�C^�Q�W�p6"��K?I��"-���ɘ�G�<ˀs7���������+���C�]'��+j����굵���[����P0�D�V L�e��h ���T(��׫�2��C?;��h��L��z�cg<�|��]����0������U�5�w2��!iM�6��/��ɉy*K�^�T���L�o�J��ٗk��%�B��M�"#o;X���ջ��W[� �Dvzq��W��f�Bz��_��4�䀎}�?p�0��B@
�(�>��-��s�0_���s�M��<l���u���B�|h%���ĨTV�z��?]ȁ-��м������u�]$�<��H|%��~&腔�ި�j���������*`.x��7��F�MSb�f@��F��$Yx�\�e���pǬ���7��F9�/���u��Ś[9��
�u�a�����3��J֏�57hJD�R~Ы<ely�^%��$.���p\�ڀ�Ӆ��/�����B(���f�h��.&M��˼mS#�S����r�k�_��]d%��C2��r�g
�"!���7����k��=��@�9�d�vM3>�q�.5�\8����O�ƺu�o�����-
�4TC��NT�(P��P�
PcI܊l��Is�Qy�
��9p6���cf�W�Bx�ibh#_��6�:��ܳ��ہ�b꟡&A�~|+�W�Xg/��Q|B:��Jf�گ�윊 �Ļ�f�*ʑ�]� �k���$qѹ߱��D?C�XY��L�&^{/s.e�=V8"�s�����6��ڼ�V$>�xw՜+��GW�1Ҝ�3i��U9�޳��bᡟy������\�����岵��� �T�Q����܈>�J/�ZVV`~�w�V�[�Z���"�� ������]3����B^�%��Ht愈�.�Y�`ܦ,�9R?�{Ue����%�x;���[�$�K�����E*z��tO� ��Y�Rl�E��6oj>Ѽ"6�F�S��-auw�/��৖�*?�O�ȯd��N�&�Ѹ���6���/�	��Gj�i�|z3:ҔK��M^v�f�pKf�4l]�H�ׅ�O���א+�V+��~Ѩ���=���I���,�d�y59G����L^��ǽ��xp�;�O�)����{ڵ[�qQ��g� �dyT	���w��/�/B�{4v��-����i&J��ߎ���#����{����*)��k?Ϩ2^�	B`�'��\�?�^"�Cu�%����4��M��'N}��,F�qo�de� �Q��k�h����"��f}�*ņ>�
q���2o�����>�Zps&K�ݐj�3-J��밯�����W����'�g�;u9硪�%��tL� /玡��"�zڿ��[��r��[����A1=����Q�����c��n�M>"��8���aY)q`�=�����5U�'�2�Ӏ��FdZ��o������*Bb��}^m%(���fB�%\B�g:
���;����TBT���1Y�]� ��m
�A��(ާ�J�[�ߕa#Jj�e���\`��r�GA�LM�
rci��<��p�i:����G|&+!�o�s ��kVh���c�-��3Bh%��[K�`2�}:+�h�ٝ�K��vD�$ȊW#�ԞW���M �?�U�z>�v������	�e;�a�g�8V�02`;���f�tt�J�����T��rX ��]�Do4<��/��}��j�QhR7���^��Ԁ�e��W> 'ׇK��F)�>�Z?���ʡ�}�
k�1?�N�7�T�\}�'�6a�o��b��Db�ݮ����c�V�X&*����r�#H]�����Y�k�pX�6\���\d��hg�w��
�M�Q٨v��p���&C�Mu�Ԟŝ��m�/rҊ���O|��`�pC����]����Q���R���/T}2�f�>RaY�����Fo ���"%ђ澔QgnVvu��_D�ǹ%?<�3Sb�J's��zIja�I�L��C�b���z�b��m�����~���`���m�G��{<�������sYqs�q���-r�r�"��6�
�+e-oz�Kl�q��s�Ƅ(o¹G��z��\�yu����0�fS�D��Zv 	&�@�	_�G���3qE2>�%��a�W��z��@��5c>,�*پ'���x:���uD^��r4	�h�/��PpK�W������W���K�%.��)���HK��sh�o��؉c\�FC�����d���x���
�'���7s�{���w�dhS�$mV[�\o򴵹��ׁ�j�?\�'x�G���wF�+�����?��<D�L��~u\E! #��m��U`��T�:�$���x?#�'���SN]�m��N�뎛�*k�w��Ч*��ց��J`Q	��r)�r��e��+DSȵ|m��'�c�!�5U$�"�]��J#��l#pl�e����Z�mn���jK�'tZM���f{d����g�35.�e��h����D�n'W����Cܝ�"J�r�@��Mw���;�
=���NΔ��_�e��	�㝨:�;����9� ��|��vB�q>��d�2������i�PǙ���u�hkz�א�OL��t+���cT���Pj�(:E���SI��t�����U%T�R	�F�o�I?mY\�`W�]���I\n��ƌ�X��[�ꝑ�V���z�������3˭����?���wNX��ѣ���G;?(�rɊ���O��>���k"��(��u�Wf�e��)8z��/��ʤe��`��ĉ����Lǒ����6q���"��'2�2%�+���O_�+�"˛sdb��X�LZ^�fLg=O-�&���3����d�B����*��X�?�<�f!AO�%�r�զ�]����\Ȇ/^[m��͔R�k$m�<�Cv7a!N)s�\��Y��<f����)��iG��g���n�y1�t±6&��Gc��u���\��,ȷ�v�k�į\���9. (��[Z
+.I>^�r�U��G4��e��ˎ�0�iгq��-eS5䇻Ľ��&���}�4#
ze�8pj�\�k��Db;2�o�]��xԘK~?�F��7�R3������s�4�1F�0��B��}a�YF},JR�ϊ��@�Àڍ:;�,ğ�t2N[y�/Y0������[o�&�2q�d�k#�+�K��qe�LZKG���Õ�R�:�#)�D���j���3гؿ��p��@��Ȑ��}B�����H���_��V�B#y7�~��c�6�ځJ{Y�-{���3(�z-%�
g��,^Q�o�+�g��H�֝J��(�	�R
g��{��m�h5^���V��cR�����Wss>��MBi�"		��-C�e�˔ʼK��kȩCnV}�B�~�jC��+
�yu�F����p䒝_;���X�Dc'� <.�K.A����k�^�:a���w�!��w����� ���2�z�z[�������G��~��Q�|�Zf4��/r�Ïȅ�)�Ĭ#�qI㞦c��ד�y�	�W�P��^$����~A w�ǿ))��	��P�6v��@�G M�"͘���(Z����O�b��U��qڙ�V�{�H�(�f�_F�to��N�|�c�ٰۣN�J ?�n��)4NW�Z�:��{V��
nu�����EDJN������=��3x�X|m�T]�g�4��2,�)O���c�V���f�Q� ��?�rP�6�r�[�=M���F n߾VԠk��"�
`䶲M��?�k4bCI�񫤓j;Y.k��:�g�kH�����]vk�!��\~�u��Z�C��c��E�C��+��G��z\��Z(tJ�Cڏ	ok�k��!E!���C�_X�~7�����;�)Y���&ϟ-A�v49&c�^�d�|��}/����U�j�I�|��inAW��Hމ1���A0J��G����K��j�������p��ҿ�n{�>�+l�K4y<�q�}�J� i�e�N3wħ8c���Vm=�o�-9�L�{¯������Y;֔��@�9t����P 3WP�&.^QZ\XV-P�,���[�aW�fv�����Ǯ�b�0}����/=���|�`��#������ ��؂6}��?��4�?S��t;7}�2A^7L۾<�`rKFάS�Ve��j5���S؞��|�~��Ni΁�a3dR=bA��r��Ĺӕ��ם�+�Cо�(���
�M�KgB�',@�Z����#�G�(���Úh��k� ��`�[�
�����,���*f��N�=�`��D�5
C91�bd|=KQ�A�.���NS�啹X��g�2�5R�@ު*����9H��%���Y��@Pne�8�_�q�i�=�<�=؂���~D>�J���p�a� 1�_��(�����2 38Kr�� 祈p�N�s"*�g*����4�p�~��Y�x�Z
IU����;�S�	������Eȕ�>U�� �Oz�o��oop�]^�\�l�Dm�3��΀�-H怩��w��Y����_���G;�%���28��8J�2���Ƣ�S1jȭ`)ΰ6�ma��a��Q.�,�	��m��]B���,��[�/Ц�NPc�υ�_��eʆt��g7�pc���S�7���ߜ�=��%�}{�X��-"�v)<�/��X�2h�u�G�V!خf̈7��#�a�ի�&Oh�^�*zmJ����]�p��_���_�a�)��J��bVN��&�NϒZ��B�v|�f�S$C/z�����w�̧{��Oꀺ=�\�11h��
��������[�o�/��I�Cp�F������ov|��k5O_<r��-���|	�1k�v���*�Y�	J�&E[��kQD!@��~j���8H�זF(�� ��O��=�R�ie�	�Me�x��lA��y&����j�b=�v��d�>����X�jQB}�[�zx��S�\L���������EE���i
��ʛ��^�Ş���i?ʤ}���b���2����W
��$��@r�ғ^Q ��[L��~+�6��e\d��	k�oEC�L�N�2Sq��uԀrm@0d�H�` gU9���),'$��x?��X����� �2(������Wn� ǋbmDr�������K��H�m\י=`Y4`6`��.�S��1`�sװ<6��^�O7��_Q����q�ZS�A��յ��\��A�M4_s�q:琑�T� !��de�]���(���'j��U�R�N�xO�p����ҧ�� �����_Z��m%���V@�{ۥT��!��r.&�>���:��$�������:y�.lw�'�P��r��֔�g�˭~�WнB�>��:�?����Jp���:f��V�2��Rh�>��1����l��&(r-��w1��4���@6�S.�p�bd�"�^�l'�esa��L��Lsb+�ޫ��W�?��ReQ'����1�7���=�L��U�R�M!]Mz"�����UCQ���hAp�܉K��!&\�Ƅ��^2A꟏i���C|��06lf�j�Am��eC#�rʝϮd	+=��"^������ɜ�Du$�)~^��΋�� ���r�jY�l�[ �~���f>v�&u����4a�jiomւMأX�(w�Y�w�����+&"�MM���^��
������95m��H�<��Y��uj������?TQ�v~������ �҅GqT�)=D<��|pgճP����l�S��Vyu�{�tܻS>xĚFiQ���D�����0�����*�[��;q	�*�#�����E\ݼ]Yz�C��,p��L ��P��Th����(��@F2+����O����۴�q��&�5�L�s>���CH��Ĺ[�y)/wNR��(�W��q� 1��Z��mЇ`{�p^ ������A��+:�YH�E�A�� 3���^���b33j�Eƕ�n���PFb�U�nl�$�Z�;��w�p�9�$@��?���g���/��.a�<�ʖ݃A �&��yKErC��Ȳd��~�%h��;�J:h�z�^*���� ��(�. 7�U���K����v�xt�A��ݺ7R�I��n���NxE�)�=�e�w?t9<Y�9y��)EvW�5ธ������������l�`"���еFv� jy��v�|�O�;��6�#���1�TE���H�7�}ą̶]7G8R��ל���K��ʵ��v��$�(�BαѰ,��xev�*qj^ �Y�wAo�Ih~�*�Fn���9F�#:um<�_�_�i�j6�z[�"	��k��W��}���g�=��t�q��pa���*��M��dƙ���� W����[>��t�s�Ę)�)�����k�0f�W�;Uv�l3DZ	1J{��Ǵ�2u��=�.(�:X�`� B�SEޭ7���&��ߣ��z#^��P�2�iψ�~Ė&�v!4�\ʲ�._�S�s��rn�S�hY��C?�>��q��vc�s�p/���؈��~[�S+�l��\��65��7;{vP�̀�R�i 3�$���"i-�'^-!�#�6�(��~�>#{O ٗX��b�"䛌n�&0<fꫵ?�.���8��WC|���1)�h�������5����)ԏ�+^A������5���]-"^�ʙ�Q|���:9Hg���Au��E��*!���2ԟ�a��tYXis�d���0	z�-?a5O�劮Ƭِ�*i�D� �!P��m�p0�^��s�,bQb�K����o�&��$C8[��ƺ�?2A"\��R��/�A1������@s�}s�g�����+�uҡ!��h�B��8`H�6N�	��8�Ai��Y#�R��F�m'�G�HW�^���<�wdA�g��ƥ=(�ֺ�N��o�؃�q�&	�	8��:,�&��o�<�t$��j@z��d���k�;v��R����H�᩻�>�,�����5���_�QGz�n�s�1��+�M?_N�7e#�nƄ<'��L���Qdd�$e���`sc��Ar
�W�
Dy�1���+�K�{�� �END*�ڊ�뮊w|(�l���fB��.
lca�2 
1�}����y�����!���"섏�D茰�'ps.Y"���"4X�ԖG���W�e�"�}�r��.9����s0S*�/eG�A�#���Sqsm��D9ړ5Zux*�N2��N}qA`�>O;wˢ�.�20��39�z�zU�Wo��r�3�n[c��8�	Z��R��!]@�	�4`���Q4(��#Y��I88۵�J KcM�Z������˭Q�C�Uj%�n������I H���`U9�xr�t��,q�{����� g��1�Ɠ��&_PBe��f]�l�����]���[B����)Sp���	���u���ec�'ۧ�N�t�Ѭ�k�9��)Q+`�[��o�Е.a< ����۪s�2+ԸC8����fI.>�/V�
����]�}Ja���Rp�{����M��Y��P���,���x_�!��Ǔ$t�
&��1�^oI�!�{�hMB����u�CL�0�L�~�(�55�D���X�;C���ϐ��Mo��y�`����B(팥fh���M���I�^N�[�nt�<�����)N
�b�;l�D�)���&?%�[����]����p�
PU&�+�%�4ԗ���׸Z�� ���2<n�`;gj��?�΄���v�̏���5)x��`PA�[agG,,}dm���U�ɨB�cP�Ak��*��W>�X�TQh�%h/�L�O38PԎ,���tv��u�*ܐ��,��_Y�k�!����j����W���❲����e�fo��|4/�6A��qp�!hk�4�P�0k3��1�-���Z��S�M9g9&�(�!�f���Ykv�E�e�NG?j�j44Bk��Qyg���d/<�:�#�L�&�{:B�C�E�=Ԏb��֛���v����P�������Z��t��|�]����x�Gp��d��ӌe��6zT���ج���8L=�%[P�yju��v�>nM��-p�>X��+������굴��kv��>�t�W��?W�p�A�-��<����[}��S���ל)��ʄi��9��/0�O�!T:�(d{��2����:ٵ��i����?�;�/�A%�v �J�����Q�ʉӿT�$&#b�"��r��L�H�z&�x��`��n3>�--d]�f����.����������3�)����8�^m �����~��?��5��]��f��}������,s���D��=k���["�D����my�^��K���U���[���B��u�"� a.)QyrY����.�F�p2~�(��I��(�fq~���oX5w�S���1V�oHD�l�F�����lVp��AP�P���\� hu5s��Հ��p�VUԷ�6��D��ԓE��\J�d�A2�^*�T%���|�9�_�;i|Ư�I�Q���e;d�ʢ��Nڦx�?o�9�~��SZ�p7�l �05ֵ�U8\��a��s�Hh����h�c��P������6Z�{�ɝ-��H�:,9� �<R�� ���nm�3�Qc� ���˥:e�eJ
��\͡:����ˮ�%�(SRa"�Fw��rU�p����dwT�f�$��Ű��m	�}���sϕ�e��&�_���"vlYn����wm��x�|I���&�!یR��0�yv8S�o���]�_]Ouw�n��۽,;��)��y[�wS3�RAn�Ff���9{�뾫l�	2q�YY
�-��@b��n�Gx[8�$y��W~�>����\�G`rJ�>�p��X��x��N�^[�"�Q����΀d,�Q��L�(���vf��7P��H�n�'[�+���^�X��j�q�8!Rj5�\٬�72�,�}P0@+~����Q��*��Êl�M�J3MQ��-e5x�Ӈ�� ���̾�>��M[�ZL�F�[>�����û�H�Sx_��r�@�M�C�D�m��X�*Qwйr��(�I�L@'Lp
���*�aL�R��U��ˊ%P���jLï���ao��%�� �QE\�TM(�dD��af(�ՎL��V(2��	-�z�������:�ՊT�t��&���g,[3���R�2�6N��ղ"�f���-�-{=U��Z�AT& ��q�Y0R�E�9�8�2��3.͢��o	 ⴬��-�Œ�X���_>gDbH��i]=b>J(//�c�a�ڍ)>���{�2P�"�I*Z�9�3}��]��'�B4��6��MX{����&�����vx�"9�۲�]U&�~��N
�14Fe$�ݡ,����D�ҀK���ٟ�%=��N�2��qLz�Xp��1]��%<��i4p{f +;#$|������BO(����H:��a�\��%]*���z�4d�)����K��e��>��ܴ��:�_�7��l�1s�Mg��	�Ru/�k}1�з.�	lLF���̧K��F;��%${s�!���>ӂ�qP����^�fO����MbZ����F�3@km{O0a�|���h����\�ZN��������7��W�urȅ����������T���]��Ѐ7��������e����1	���%���+�ӏ�C����V���	Ŗ��'l	�a�Z���_�2���I���U�>Sv��J@�Ys�i�t�w`׮+�������cP�`�3��i��Y%���WE��V�����j�ܬmI�7��|X������Y6(`���;�j� +/�8��ʡ�d@��T��ݨ�d|��L�Љ�d�v��يc��!��!����T�1XB}�ؚ��׉Y��N����v>6�ji����w����yb#NӚ�����VNG7y��2�B��#�thiB�˱�,NU1�T�j�����"J�ar�x���We����}��������L���"��A,M�7�^��}�\:�Xl}ћ���!����)��-�De6kw�x��Q�/ ��j�����RL��8u�S���N���2�i9�d��Ɇ��UO�z�&���I�!�=�<L�y�<������(_[ꃵ�%S��B6ү�=�y�%���=g�<9f���uSD���x�̗�i��?�soµ���=���3�t��<V�QF�	I�ڤ�T8R�<E�1{>q�G�\�E���S�p��,�g$�aU�"�{G��p))Rn��Gz�6μ���6���s���<�4bQP"�K�%/��$`����{��ı)��V\UV�$�My�8��}�󯕔F�2�	�G\���*7��>7ב[s�#����tDG ��X�mm)A�c�,g���'�9E2��"�O�K�!,�)���g��፛T�URG���B�k쵬{i�>��������e��@�A�P��T"�)��q�btOY( p����E7/UY6��R��!��iv:��@O��-=7\���tgV�0���>�)�[��T*h{9�T9K�r����D���UXd),���[��x��]g<$��	���Y�K��	�]�~�Һ�P�P$�U��:!b�MyC�uF�?��<(9�m+]$������t	æ�X8�Pv�,��ض}�ΐX)�)Qr�oQf���[-��@
�Pu��CS���-⚮P\��ó�/�QT���������.?�o����Sg�j��W�Fq!˗��f��H�g�=���TH�.�����Ӫn�q��p���y�� ��FFFn*,�V�7'j����к�`�(��#�'�8wLv¹��.��k��cdu+�����_�l����#D�� ����o�"�d��*�1I�k о2G���0�=�0��
���!���V�����Ɗ�g�x<��!*I�9�#l8���k�e��YSQ�yt]����uo�h��\��'&�L���B%F�J��v
]�~�V�1mAMm�ͻ�\��~H��s�#?�*��v�<,��+���j�>7�t_7�S�����t�Xj� ��㭼^��Ӯ�����?���yZ��v��]�A��0r�z��v��(X�JU.�0�a̓�n��sXH*�Th���I3���0#�U����>9S�U��GE��_!�)�0<�ڟ�Ն���Fn-��:��8w�%�s�j͸�+^a�{��-tp�6�ͩ4a�G�p=�U���U�p�c�G�r�i]��ex�Ȧ����d��U��2<G�lY*�P�1���ayQ���q��,Uy�k����$���ѷ������Z1�z:K6��>Tzwd �P���=3�OS��P�o�2���j/#L*�����&z��j{��.�蘓��,�dm�H�l:R�1��H�&0�~�-�1[UB�1�
��[](0i�*����B���O!ڻ*�HoM�j�k�t��,RБ.q���S2�E�.C80�:A�����#3] n�dI��Ye�hvң���*���'�Ld�����+�tUUכ߅F�:�q�_
Ltμd�+���`އ�eM����@�Q��ۃ7Y����([/�kTZs�F���S
��rp�ʫ4]|�U�ə<�k�%Ů' �j+p�7�EG^Fym=�!1�����a�kn-���j��J��:��E���M��f�XTv�����5���ͩ*G�$r�<Ӱ�L+�>�_l,���ܲR��g\��4-|�VN��py���~�/��R`��H5�_ݞ��+�b�W�v�M�K�&Jv^qڢ#��]3���d2��"F��L_�/aݙ�kV��u�ZB������V����]�a��d��w���X�d2��ri5��:���Eg��I҅o;ӧ��Ω�v�%^��G(�P)ҹ_����y	*�x��F��I�+�۠7�d��i��ّ4暁TG<�����Ћ�/�Ū%V�z��9{J����&Z6��gq{���\+�VD(��=[�|\3��IPZ�tg�=����}�,��n	�9k�.��j2�rg��C�����M�X�l��c�Ʌx2Z�!�%V���6��1+�ƫRx�h3Ĩ�Dx*ɾ�r�fh��qn��Jx��pM�*ǝ�n�6��8󒊛Պ�����q����,��V�7��aR���Q�RN]�AB}�5���}�B(Ӻ�l�&���|c��!��hss�=�Z�d�Y���o��X n��V�p�T"�vn(����"�����>L�k��ǳ�h����u�"�Zu�c���<�`�,M��B:��2^�v��d����n���y(��LRXp�������@.��a���������$73��"�{*�P1H9�؇K~�D�1�<e�Lz��g[l`+5�M�Z�- i���t��/���9���օ �K��j� ��(R{�N�W�x����Vt������Z5�z�Z~5��ŉ��='��ٖu����5P������7N�ՅI^ɗyӳ�)H��5���Q����J�`�k-�+,,����p�1�8�'x�}ϻy��r>q�=°��ad���,Ę
5����2�!���zձ��j鉂{L���X�ϻ��6J���l���7�PwۤX�+4�.�����&Q���,�0��5�ա9D��D/KM�6y.���&h��R���[��ma�C�|�1���3��`�7f�K��VY���&�e�d�]��-!�96�]�h�"<�}�*��� FZo�l�
�)$��Jh����2�?x:�!Ei-�F�-�nDc�(�,["��i:{bK�3��A�2#�3EvU e��(���<�"����qbˌ�\�FuH� �1�`6��e�y�AT+xkۑM�W��I���mS�xJIW¦zk��k�k	������?��X&:9�3/���k�-k��bAZU��S�.u��_*��'�ۣ������-f�L���H�=�2w̞���	��S�EmH�x�����q�'�t� ���&K)BG��� �J��oI�E�~`�����@O���_�"��:�J?
��r8�7�]��G���O�HiW7�~�\{�v;͹j9��[�����X=܆�B��7�/�Ī3fl�Ԃ��\	��d�
��th�*���+2�z��y�빉�Ja,3,\:����D,�-�	ɡv���l�/�8�Ċ��b�E<��r�0�*'��#��t�+�t�s~��CB
id�o�:�`��kk-9Y�S�c��$�l�0q9<��$�V.佃�!���<��~�����59`����v�ty���w��f�)�����p��j0[/G�q�P��8}��ir7��g:��*�����F�\.�N���B��a�hD	�Jax���l��E������К�t����˕IO��ةz8�q=�[P0�2�P4>�;҄�\)&�����b�''�y��+B�#Mqy��Y��ߞ+��	������I����;	m��>�#Uwd�ƫ|Ζ;�D2@��8��L����8��#H*�ָx��0��.T�i�����)�B�<�܏�>h�K�l��Tl�����1`����^��T~yc*W�?�Nc�%�B~�C`�ɀr҆�e�ST�q>A�Y�{�����$8��,���^1Ԙ��O4x[x�2���̿��#���i��V;�0�Hb�x�Kj�z�r�A8g~|'�ax��/�k?�ӛW��wƌϺ���h���F�+�������3�\>
q-E_a`��uh��a���*
G��RL΄�&�߃��n���X!$�m��t� ΢����6������f�Y`N~�^��>� ��]c9j+�Ƭd��w���O���B��M�@��P�!��D�]�@&�=p�H^�UE�#��U��@��=�*�-p�)2�����6t$$ć��`^�����æg�%i#ܹ�&ќ�0Ho�r�V��[�r�&~���]wg;��2m�7��O����p����3����K��_��
���E�x���~�x<��� �/5��%��l����݈z��`1��(�`S����>[�� �N`+_�(����̼��jZ(W>w���Ԧ�/���y1�IV��w�K6��:m�ި���'���8v w��X2:�[�,�?�Y�m7�\ބ�ߞ,0n_F�.�Զ�^Jh���X�o���� �6�gC}�O�ً	C�RJ�8j��,*���ГTg�?���󛑙W |�j���	�_��{�c�i�%lގd�b�.���'Ŏ���8o�*|�1H�QA������/�����k�T}�Z����B8>�]q�
R�O5��~�=MW"g�&Imr�qƕ:�6/�\��e�2����?���W�G�>�/&_��5tYd�a��v�\Q�G���%-�V~i%D�������EM��4�����<ʒ{gV� ���T�0n���G�O��C���(T�Q�±ǜ�2o^��	V���5ɫ�Vn�����t-�̀G���0h�<n̒Q�ɐP!��?*?�̭c�6�/�9��\���R�����[��B�$�)�@]��Z��s��T(�A�PG'np����X��|T��"r8ka$�{}O�R�gi��F�8�YU�b[!}�1Ec�]����?\G�������84o�]`�`������<����7�Ǫ�r�r.�<��ٯ�=��*��`�{���bs�R�%�s�a\h�R�=��w���R*r*�L8� R��n�zʔ���c�A����XXhZ^F�5�,u\�b�QM�%kѢr���C����A*w%R}���[8@k3BK�$<P�PPp	�\�7U�rh<�Q�J��>��V���H*{���ja����K���љ�f,�蒇fR�^��<�l�7��Z8}��k)\պWNIT�S]� ���6�	��p̮)� �1���ts����I�7����,�o�ʠ�6��kfd\,$K՝dW�����*��WNc��3&k[�Q�-o�������Q�$ l׽�M}�ccz�ER^�N�!�\�� '-feq�>Y ~��ְTf�=�նĻ�5��W��0ž�'v0vc���TlF�]뭋�x}h�0uU,�����0�L�����;7v�x��B`%�e䆹'+��8T�$�~���H�@�,[M�0+i����ʇ�#B,��YA^��xm1��g�����UHZ�Ƶ�bT�x�.coZm<�ȗ���%w�澍���	�CG�
�)�v9�J�*e���~��"�	�@�Њ�򲆩�X�;V�^�=  ���Sbi�����[/�%\����ں4Y:[&����"{��V��N1+��;ea/�M������</���$��)�5����7�o�v�hX�'����7m-�s�~]���C��IHRM�xJ�`�1����̱rG�F���>nD��I�a]�m��O��X��U�G��غ+*���7�L���@T�N�q�.�eF`�N�)��,�K*ɴ�?	B27 Ӥ�X^����s�իO�/�w���\�.��؎�c�J�Y�г�:{0`Gzz�)�-��3ǘ�\R(E�-����2nDMs��6u����q�yπ�(�`'���u���񎂫A�]�"�k��d�r�h�)�ǎs����2�=��=׍�/h�J${��x��T���N����������j	V9I̗�����_��]���p�=������_���hKz7�Pfx��`�g�;Z0>����>ّ�������qx�w_պ� @{d$��jo=|�#C��I�`�pjg�� 6�Oz�8�)�H�β��y���v�X\j0��Ť�@� �1$�F�<BK��K��͆C@ ?��ӽv9��@��*����h>��ZVPt2�[X,�k����h�/��Ck�G���.�q&��}��"n;�_'���{k�j@��V-�C-�5�f+�KdA7��EtCۇ��Z�%�f�+_���Y��L"H��['-f��	30Bc�Ņr�J�����Q��W�k��_𼙝��*��o#�LZ���$Ȁ�Ui	O�2��Y�ɭ}+�,���P�!T���9#�y������hd��}1o��>Y�[��&�]�O���y������	Ĩ������""	-o?�U���s���Mk��,����đU:�­ �u:Ҏ׋m̽~mbSc00��U�X�Q��v_rx���>�2@��R��ON� �|�g��ݜG�D#�\��e��!z��&���W��!G�XӋ���C4|&����������6��n�bS�\ͽ�z�A�Zo~��t`m-_���fmδ�v���~6��Q39�����F݂��<U8�:ܢ��2S��~�&��c6�;*�\�CA^.�n.�~��(��S�K�-�6�.s}f�606 I��d�j���Q�P1+���A�EO]/-�-�q��v�n��J�y�2��l���@����� �vá�iƸf\��1��.���
Q��!ZU�$�����v����sl�BV �������#}��5M}�w���ϭm�=�c����T�����E���J�%�]��=A8����M�WY-�&T	G�B�`��v����Ts��X>B9�Lyڏ5h~���'R/��I�/Q�y;#�C+r��ç��-)ێ�y~��-� N��am�Ӑ���)���|B���Z�,J��d�6VՂ�i}�;0~��(z(���9�,���u��������Ŀ=� �H�[��,����W�7�E/Ҫ�|+Ea���g������������������nE�s�`��(~���<
v��ن.]���D#`�Q�Iʐ�ѡ��C�;��t��٪u��������O�W�J`Gڝ5��������k����+�gal�`�v�;0����Мµ)P�{E֭�q��_�KT�um&�_��\Akdm��9�~-o=�T� r��.�5Ȇ�,X����O�p+���bϩ~�Bg��l���d�B@�Xq������[��\��=ݔU7钰R���}��v��XX�?H���Ea`�|��o������WN��G
�$�v�7�9#����3G&8��P탇��*�Ӱ�gr�����D�f�u.?0��J>I���T3)��]��H�C J����}�nst<�l�fL�S٥]ed�n2�a�����Kw�=DGT�/l�c�VyBP<�Bm����Kd�Y��~`�]�h�u��^ƺ��fz�H�I��1�G�_C%F�%�߯��6�g�&Ar#.��J�O�Gk��k����~��wa
���� +7�7���.K��ʀ���G��V�a���b��i�7���38��K�%~Z���lsY_8}���ߍ�e��p�1��a5��zf:�@��v��p�n:�Z6�'��a1��D�t���2��j���5N���\~a�.�B���Yr��p*����_�LsNxS�z��y�Sjj��DԊ���!�����w_��� ��i@���9yp)�-{�&���!��p����0�^^�2�D�$v0���IU���Z�c�ץ��b
y�_��>$%r�C���¢@�� �7�D���#�;����Y��e3�-J�G6�z,��/ߒ�7�.��f�*d�/��hl�ݭJr�R��Bq�Vf�A�IWU��J>�����q�l�y��7�6�����q2�;�kDH�R�q^��dĩ�s�0+Y�X`k񲛮o��K\���+��א��k!�9�s�5m-*Ȱ����\5^��)@K?%�ة��n7�t��/rL��r�Com��	Bf<�/�f�C���A���� !�a#nW��P��Qz6y��Fz�1���YRC���޻|�}�����$��d[ssHષc�>+i'i�K#p���%�"&r $H��5I3Hp����՟����U	> �X K�����G�y�E|���hS+�#m�� �?Z^�0��N�&�b]<�^�@64��W~�8�i(a[ޔȘ`�R
���+������n�$���	���S'��'8Cꖔ�ɘ������ʹLd���7�r�;���@�H^�K�#[��.��c<�h[	��?���͓�W%��/�c]�1�1�9M�g�Ϸ|��
a�FsGu�w0� �k)ϝ�1�
r|�������{Gχ��'V��vw ��I��[6�-��1��\ջ<v�SPC�Ֆ82N�kc�V���/\�h�ٰd��>�F�F~�G��ǒ��; ����T3U.Z���C�,PΦ�Ew�װ<�Ү�XY��l�{)ߚ�H��嫘��[�P6�����K$�j��nCt�q�U¸��0��jF�a�I�BP8D��^�Y",�x�+V-�7(S��{���#�в�2Nڇ�;����f��˅�q�j�⃬���6�5��.�KQ�`�c���(�oo[&��� ��a����1�j�᚜�b�\Z[,w �.BÇ&���
rh+f謫��7�?��@�1凇�9�K$�kIǶ�u+/v�ٝ����\���z�W��4�"��;�����چ�4npDh���尀k��Z�0��'; 	S)�7s�l��ϔu9I!\���z��=H�V\<z���=��4
ZL{1c�`��fo�M��ĆuЩ��1�����@�x�N��b O�c;\�d�4f��F�;S_d%W���
�Aw�kM�\\���lWYugTv@,�3q�_QQyB}?Ĺ�E�(t����g��]�(�9n8��	sO�ѥ�����Q��3�ll��H�r��8�x�ђ��z-��������p�u������7x�Ӣ��X@�����	z�@c�'�����s.7,��a;ΘL*�nZO�*CEi�!��1[�-ȔW�G� �����c�?����Uxo��_p]��<o���h2]����d��V���~�����?.�"���B�Ι���H�9-����@<�9g�dCjصv8�Fۑ���)���-Y' �U�u���YJ,�Jwn4�W���h�m����;���+f3��� O���^Å�|q/�T'o�={R��@�����$ZUql~������@���[A�aZ�V\�d�B��$$�D���1��D�eV�S���wy�����װ�:���[]�9�g�IjN���+��� �2}�Cq��NvXG+.:��^��Ҡ+A�A��$#k�Fq@�	oRc��,�����y����h�ד2�F\Ƭח�����E-�Ľ;���$!i����Ԭ��d�VO��(@����#��9��׆۲]�uq2ޑIk`������a��x7�N]� ��~W��Cb:&o�<W�3%S�VI��}s@v�'S�r)�9|�ݐU��؈��L�K��W���"k����a7�����%����A*�r�5�	��9�O�-�9>$Qe�ϒ���U�S������@R�����;�����w�K��k*D�������r~����*�G�x���zC2I�3����J��_2Vw�Ckʋ�?�Za�Iz_��?�r��%�~G^	�x���1�hUڕ��^RGm��7���=�6н�Z���vu�u%Х��Lbn{zJ�]w�AK]P8h��A��e��> �idv� 1�R1���ٮ����։¶K��n{_����\�
j��}p<�1jLVE䥆����A|L�Q0� �C
��M�=�X��DgM�u��"b�$�ed��tܐ��v� ��H��>�Fj��}h�8��i���s��iy|6'+��{&-���
��G�D����*��T3�PsgO.�MU�*�Ia�l��m��\ߑN�0��I����}T!4A?���@0�W�J.IFwv�c�-X��I�O}o�ѿZ�')�1�PeI�IU���h}%��+)([��ͱ_:�c��vrRM����ʣty���P9�VA�PE�Ó�X�)�j6���8�H ��UvF�?
>���Ta.�Eݨ�'���Հ�+���dċ�1ס���� @x��ƺ����yeTO�g���=�%8e�Th�3ʠ]/_�
ۖ�-b�f��/�� ��]e
T���Gc�~���8�l��/���#��� ����q4����W�T���+-�v9�%�� 5F�cXFA��=���l��#�����V}T6Z��M���x����?Oǒ;�f�����a���BA�8�̠���C�<����Pr�-���m'��[3@�?l�@PF51so1�f��|oB�����M�G�O�r�;��do��T�~����	��,���(BՂ�������`}u�G��Tv�p}���{��P�q����SE�X/�+VGwp����̊�
��N�CBҏCtd���%\z ۏ��V������T��l���,�.B/�p�}n7K��v��^=Ku�(�R��&�H����u'�ė癇���g(��$5�bhPGΏ@�zL�ԫy�'/I�&X!�1a��2*-%ZR�Z�11�ȯ��6<�|ǲQ�� ;+[��q&��z�d��,��o��������ڱ����>�
$悸�#��0G�-w����+�ߕ��!:���2��R��6.b�Cz5�X�xi!E�x��D��iӌM��&� �������ey�+<����g�L�N��{�^��Q$��cP��Q�K�r����ϱ~s�~���μ˝����6�߉��`xs�7k�\aѕz��[����Y��$�ͷf�&��5e�u7B�E'�|��φ5cD�揞Eb("��d��w:408������>�v��r����쫄��uם��3�V;��ȇ�mi��@����k�B �C�T����������bNb]JK��`�MqL�.C��.4�H��3�e���x(����pќJK��
/�����P6��ڤ378�U�btN�?Hgn6`�nOe��P��+�sAHzm��P黯��c�9�몭!�\!}u��n��t�����R�lR ����D)�6f���'ܹ��%7%����!�P�pGQ2����$�j��/o����\o̚��C\��	,���5��b�����Y��"�pC�5Upbx�o��n�V/."^�c~ö���S-����I��5M͜�ճEL=ف�ə\y/���h���S y~��*6G��(���٠��H�9�_V�{XN�C�QF���en5���r�<7B�V��>�N�+�ī�������2iL�}�1�)�2���
A�J��,�1�
÷0{�MM$Ҿ�/�Z�n@�?�c��yT����/d/L�l��[M�˲-U��bK�z
2�L���N���{>��? !Hq&1&B�l��Z��'L���츲�N̶�\��Jq_�����ҟ\@ߖ[BZv����gC� �3;�,�;��դl/�%zoB;�ຜGj{���k�-g஁&p�Wߥt\��}4Y-�Bn_���Cch�v_�,���1�?���1Jl�b�op�	�&�`�Kp�����=�#3Ui�]\��t����a^�;�ޣ\D� � ��U���.�l[�Ks����b{�չ�Z�Z��*+ͺ�}$:��Jn��n�%ʽl����N�;^Z�'p,�e�ӝ���9@�s���~���i�^^*�#۵�@=�,�G�����~��#��1�4�iH�&�vb٫��_�ˏg�5}�<�hC�~��Փ�*���Rn|r�` B�b8_(;^"Y��J�{�Mz�d^U���~�_�n��8.��Ј�l�C��a���w��MGp� yAC�/�4�gVA�����Aj������۵d��L����6"u��B�|����?'7�j��J������1Ma�?����@�U�$L���JcKr�Z��YH��ֳ?��=�kn=s/I�u�[��Y�^P� �䦝�T�[��'H�#��g������7p����p�N�CK멨�ő�7��
��.��|%�l;���9lg򼥱��N�
v�tGmo����eSҢ�m+�|�j@��:�.A`q����#�~�ڨR�~��SiS{�v�����n�#�u��~��ݦrE�+Vt���%��c��sa)��̪�����h����$"Uo�в�AX��^@ы��ZM�_��������}Gv�p.��>пj�R�D��f�U��,`��T�ޜX��ewj�����- �Vޭ=�5S��%w�V��LH��w�_O�������R�?������1�>���]����-�������Mi_;/�U�4/mO�7��������t���[]K���%���z�W��+�A�^�G��:��3#��f�q[��=O����Rd��Z�m�ttT$���SD9���8%�C�t�A�R�WǴ�;VLQ��\��Ŕ�d*C�P6�X�s3���CtАe]נ
eFA�QT�}Ā�̒�����E5&�L�RdB�8������`�:퉜t}{�.�_LU5,�-�Qo'W���~��NVlV~�q�W��tԸ]��T:�C���:hf�,��e��kub��A}~9ry�/"Z�.���L���.J�bS@��w���[�PB5�g�e43�`�9�IF�A����ɛ���a�+%#��ˑ��3����[0�S#5���m���k��n}me��:��e�g���o�NVK�,0Z#�%E�D�����8�6��./%���;����!q4�G�,褝vk\ǔ&ʥ��c�$���1��&��I��Z��R�o��w�)�xʲr�.2Jٓ��%G�3��¤�E���;{�^�O�)���ǼJ�i6kR��O1�<j�[U���b���W$�27���:�p߂-��z �t�H����3���+OI�@0D�m)�#ұ�y��pެ^Eݛ�5��-�S6O ���k�w N<}�[�ܤ��('�i�h`{�W7m�&�Q]�����Bu(�mnqP�]�߽�A�����c<���\m�ΜbY
�����wh�v�^e�|/9�D�gٶno��a�}�	{OO��vr��З�}�f/�·y&���2p>X�Na?��!�ua)�u0=eV��S�����L�fi�p��.Ui��5f��yq�q}� �qiX��dC����r�?ʵ:,bq7�y��~�����G�[~�@d�d~�&&�K�/ ��9��M�#|p�ھ�nQ����O��#r�J���d�杅>��x��#_��R)
�����o��B l���)*��O$�d�
��-�C`
υ3���X֟��h�.����J��X7K<��(�"�M�7������҃e�uV���'��$F�q���!�l�fWrܔ��N=h�'�VXP��e�WϘ1n�\:`)���u��uӃ�lD���zn��ړ4�xK��y���GK�0bv@n�Gt
�)��$9?�[��j��ʫ����S�h�>B��.��Κ����V��S�	�_������lK=�ڔ$�;ƙMz\K�'�9�u�u���[i�G�4��AD.?T��Jg	�<��t����w�C<����H�t��G�K-Z�3Tp�Dϋ-������<��wxK��= ���0`�{|-=	%hg ����U^�n�iNG�誒MVq-w�,ЩJ�@x��?1�l� wJ�	u/N�(b��Y��֝��RgO�\^�HrG�@�SF��ç�[
PO�Df��TMM���n���&�E��	�"�gԂ�UnfIڡM�*cp6��^���Cj�G#��>2���c?�[x֞�|&��o����#l!��H˽����_-�aY4�Y������4���t�3��.��)oIp��x��(��+x��_�F�튱i0 v�o�ʫ�b=�
�6��_�����ڶ����%�];�)�K|5�O��C'�.d
ߜ�Wi�fP��^2)��ؐ�
�����k(8��ޤJ�`��0��ћ��[�";���{��3owje��� f=���̙�]�Iޙ)��)�F��{�&�����X��"��f$�0��EJP[It����u��r���~���1+_��).)���_����"w;����b���H��gH��t�����+H��׌ҽ)C�/pa"g"�WU�.�+�:��9(q�D sa�/��2�)�{I฻��W��g�Qn=�${��� ��?! ��kXY)�"Ѣ���DM+��]"S�t]��H�7����ak�H�Hq3�&(���J�J~T�:�6��b`#�G�U���d��LM�$$��[?��H�хٟ�Dh�2�(�7�J�39�Dp�ײX�T�q&$�0����t��@������wJ$E��?L�W�x����˴7����+��ǵ�O̸s�������3��뻣�\8�c��K�__rn^���|�j2��;�_m ��.�b#KF�K�u�B�O��Ao���yw,} �z�>�����������g5��Ir:��P89�&���x5�v�|�`�%wM	n&	��2� g؅�L����Fج�D���OL;�`׾�H�c�^z$Mz��Bp��zq�/��N�F��bꞭ*����` ��ў���g��-JV��8�mVԨHC��jo#�5V4�۝h�1�lQ�J�F����[t�Ij��wi�&�,o�]��a�4�ajCM���ꀿݎf�E�^���c���(���`���{�@�D�B�F�J�pFp�tw���[��5t�������G���}�!}j�I�MH���k�Ƒ�N�u�FR��(C�5�.# Bc���*kR��
2��Rࡻ4��dI�)A"q:PE��S{�ܰףz~�P�M#�����q�i8,,|14��<���S>%H�V�A?��0�!
]#�~���E[�aջ|Rj�Ô��/p��2p�x���� ��2.۳�o����|� �v���ٿ`�9��ǜuql
����;6K}Xu���g$���<�FO�F���Q���s5��O:f�?��s֧�G"���^^RL�1��$"�VȚ��z�w����0�i���t)��p��Φ��H�Ay+]m;��r�&���G'ؓ~Ր��0�r�v�t���������#�����;�gO娎|���G2bX����,߯)�����{<g�_�Oc�7�x���l�?�|읦�3<o��{��m;=[�ѭP���"]���?qr����J�y��Z�Lk�l@T`�p\%����6I@�3�z@tL�܉W�F��y㑆e)yINl�*��Ub�,V:�!�.���׮Iz�3(��ce��2�7ș����c~}��Ӆ��A?��S���^%{$�A0�|���	�I�|)���+�!�B�,���n����� ZB��ދ�Y�c�I����V~J�eT>A.�Q���]9ְ�6Y�&��!�����o��t�BO.Ȗ��/����X t�ۢ�f,���qћ�b���o�w�`])s���n�rI�����!�`��~S�q��~����dE�qq%E�I�M�Ff:����C���:�̟z�&��E�3Ȗ$����ٹ���]�w���'^���<Sd�O	��C��XS9��^.��!ҖT�p�8�(��&�@�X|1��}��v"������Z�p�H�P�I�I�G�z��O#��Ο1n��{* �9��]@P�% ݙ���l�9�H�	#����@�s�")=�!K��D4�uA0�f斑���qU2?8f��]���0QZ��2y��(�Ln�ſ��<I<�xGdպo0:!їO�Mf/�f?3 �?T[$�����D�'e�k�wI���ncL��NG3G4r����J]��4\
�Q��;�"�v\�d'��¾
�$��@	�u�&:��b=�Y[�Y�NcgJ�/*�!��%��h0KIl�?tV��C�y�(LL�~낂'�:p���}2g)�_�3���M�½��\}k<8�V�H�1s����E|A����e��u2�j�	�_��J�A��y�v���z�	~���_��h��?G&�<��}I�+Yiߠߙy;�$?s�m�9��剉Q��w�L���{�+y��9�K{V`U�Ώ߄����m����,��F5�6�-�µ|�����R��V�ϧ�����~�OXQ��1�@F��Ұ�Y�N_? ��������p��^��#�.�7�~q!�7��OF�Ř�y�}O�H5DeD,�-(�Zv�F|՟!���c�>������͗Iv��u2���Y�F*^�MbN}k��h��V��Ѵ\^Ge�����]J"=wd�=�V�s\�XD�E#W*58�P���a��S�����8� @���]؅�𘺖]Nt��V�+
^	L�FJ�%z3����`����ϟ�$m���we�H��3D�4�<l.yKf�&?3�b,/	��Aj0����P���6~��o~��3�H?�<�%!vc��aE�P-RE�/&�T�.W��e� 9mOp9 ����#�
���@�jg�,,���1���\zgSj�~��__^�x�y������&�P�WO���<��>1�)O���	�Z�rG�y�?/	���(hE-�g��p��ѵ,i�F��mQ�L�	c �u���9kD�Ik���zƃE���0�N�'V�0�V �}��TL;�ӗd�Z��`W� �	PԂ� >AM��MY@�|m}u���6��B����^d���Ip�вL�fx��4O>hrI�1Rk\��NN�A~�ķ^��|Cݥ��Xq&.Ϸ� \.���
�y |`�5���<��+Ч��}s���"�)����U4U���e�lDO�}D2�胾V�
Ü�c�iS!/����ƌ$�E��8d��.��$���3�ߠ��PoO6k`M#�n_|SrS������۠" i��uJ'�a_�i3Ը��+��k�m��w|Y�SSC��?���~9�c[�"PT�|wC��tiv�8��\��'�Y����G����K�00��}��8��C��Fl���6��w ��m�_�>����u)�����~�Iw����!�y�XE1�
� �Ì�p|B(+@ȕ�wk�v���G���.���3=��]����.=��.x>yC��3�WW�U�E8����yX��3Z��p�5����0������NS�z�������H��:������Z���r�tb�R_���W��DQc��	�g���0'�ix����zS�oH3���Nb�l��Խ�5��ޜ9�����\t�Ҁ �$���C���셠U�ϠS	)���=��ڎ~;�`���?D!�ͅ��'7 ����ŏE�ʄ�Ϧ	�e�s8�P��
�_��L*��À��\�`o��WF�����D�᥃�4�n`!IZ�;0�Z^���	��bzb�m�U˄	��0�#���4��'�gk��T�ȃ�d���;��r�zŽ�h|�LL���� ��<
9RZ"M"ǭv=<7�&oF��d��Wx��k�tԶ�;�Y$�@�~�h�;����_>3�e�L��OA&��<�Yl��Hz@���o��!*>�Չՙmb&=��$EJ��=1m�]�����4�H���-�����DW����U`K��t�<���
����Χ#��yXZQЭ���N�#IPL�͉�Qa��>j ���!ӅY��͵G���E��D2AExP��$�B��B�o[��w��]!���5�`U�ӱ���/���w#N�1�>��.(.�(vApſ����Ϝ���k�Jj�\�=�^�:P�N��C��su���YͲ��xE-�]A5�ofy�� $�$^�+��&�_P*�5,��&GG[n�	6s�r:)�����a���k�B��h��9&-���̘���$bVl��Y��Bz'`�u�"�kO���tC���".�S�__r_�f%2\!��:�sXD�p,� ��i��NJ�r��c����=��*909���X�#8G�]�/��qh������ZC	�B!7�����]Ble���`���Vb("(0a����"�k��<�(-p�Vӈ"s\R:���7��J�҄tu[�)�j��	F��vQ��^۬���wY�4,l[��� Y+ik�ȴ!���kk]���2��$sW�����B������Ui�c��}X&��a�(z���}����C��JV ��Э��4��\Z1)[J��ԏ{���UkS'�-��e�~>��2Cw`F�.g��5�s�1�X�[|��QC� �`w��c(�K���>�I8��Ϛ�si��2˽���{�[��:H�
�t��Mg'�`p���N�~�}Us�a�������Ǣ^D��	n�D�r���{#�KR��e�_tU��%��(�<N��=��y ���`��ͼ�܋�A��ѭ�B��\"����Ow�iT��GR�A~%���S�@�*E�M�:A�L�!qW�u2�-��:�:t�� ���``��PИ�뿈
1��C,4
�Z���S��!g=�'�R"݆�2p�@�O��1ۈxA*^ʹpg�v -��r��	1~u�t��hb�Cש�03g�3�V'��Nr��<6��*���¾����FƙP�W٢/�h-���a�7%�􆉕�N��u�֊!sg?$e���g,�����y�T͠��#B7y��o��P�y��/��7ڶ��.K�����4�X�)� @���$w�T������vѹ���#Ka��h���.=���^DR��~��E�[[�����`���N���J	o+��T�L�,�|�-`��̀���`:S)�����ֻ ����\�����	d�����r~���16�"��9�sT2������퇪 }ؗ(5�ƌOt�D3U3n���ӿ�G������2��?b30C�,q��RP�Χ�0����g(�'3b���UG"$0yW~^��cA������*�ٌ���u�¨��Փ���2��(Z��R{�?�q9�_���v��z#;�z�I�����؈F�c�~�A�"z�>�W���31��f�i\�������Z���A�_����3U�H�Z	���Q��6J��
%c�'u��G>��LM�Ԍ�MUM��Ҵ��3��	�+8V�u����9c���^��a�����߽�
��U�Q��ʟ���=��{UJ7�WJ�4Ζ���8��6G��$�9�t��
#�Cl��'�c����<˕��-�5��3#]qm��
����c@��#��r`l'�^�fXU�|���L7e���!�kz��������4[�t����^���kb����Jt�5���B��r��Oz��.�v)ȏ�7ϧq����??{�J?�¹�H�� �2d��U�'���V����U霣~�F��3&v~Ψ���8��@�3=W��5'��Sq�2�7�����5�튠�o(+�
r%4!���j���n�&�c:�;@2��Ċ[?���1���8�#U.=x�F�sF�J�=ui��6�4H�;X�����:d���0�nm���W��wx`���sv-��������&(��v�OB/��˙�=Wa!��d8���@3H1	��!�p��UL?��>���{��?�!�:���_G%j��2��$<��v� ��R9�����E�I��:A�W�9vM�Z��&�r=	�]��Ш��w6G�Pe⦩��/7C>?�}�����E������!:����n��,
���#)���Yb�n��pna����2���JIL�ڋ@��Bi.2�Ƣט&�&�:;6�����&*$��d��G� �+���m<�]{33F����T�'�֫hk�o�
{���+��b��~̈́=��b�8�q�Fvʕqy���u�-���d�Q�d�˙z��9�����7w��zWSͻ�]e0}!4k���4���z�o] �2�Y�1ɍ�be����ʓJ�v�7����7G�lx���hT�.�|.LU\��0g$Ğ��v���2��p�1:р��{~/bɵ�@�����XE�Ur�'�..���9���J��|}�����U����9�A0�:��n������ڿ"`�dŒ��3-;i-���.n��G�x�/<A0��*�UkR\rg:Q��$w�Co�94�D�*��enD��Ƅ<���:�<L@�L�x��s���E�E����T-��B|Fk� �QN?��U	�{��na������Ƚ�E��@_��9_�2�ƙ�ē��p��1�����h�=�?D�Ɂ��[�A��,ʅ!����)Ey٬ĝ�5�1�G�u�
HXc.8B����1�i���z�k��,� |��� ���K�8�޺��u*�~����_l�"����m�m�,ǧ3C�Vh��\-U��;+fr�.���7�>o-xU��O5%��C�讜b��rU�ˠ��N�ZM��`6=R����8��k����Z �.zA :edrh�6��#��.�xHQI˭�ϗ�@rIh�Z��8mh�I����7^�/�˜�}	��ۋ����������;��Ԑ���/!����F��{&mHϕ1�R��a�a�?m���J�+���"����r�0�Ql�-���P�7�8�i�Y˹։�:���{���kJ�Q$f�LO�I�L��n�%�o�����V�c��޽?��j/ 5��Y��_�m�8�\Y�!�D���8P����3�+`���n��{&��ԑQ�Y�R���Z���2���z���,4��� ����"�}��O�@gn�690���$;ä*�Z��sZ+H�`�Ҿ_��Cv���?E�qr���w|���s8݂K�d��x �����	���T��+����{�k,�3c{B�����*�IVf޾���t,^ݖ50}�è{e��|����LMTǽvV����Sb�C.�X�w�vz�����.�v���7�n�%��d��5��
�r��d��dl��٣�;M7���teH���,�I{�
ͷ)��c�����G�������GV�"��r^�c��Pg���~�|�S� >�d�	;\2Do�"������T���Q&����1�6ר��{�=�	�wm��5t�ݸ���V���H�� ��|�Nm�QF��q	��%*��\�M�����y�{��Mh���$��e.S�)t��K�,�婮}\�R��o︖E���5GƘ!d�x1�?�z�6$�
6�}R�8���j����g�	��bv@�.QE �P+t��%�j�'auJ�+�v1s�[Ԡ�;�E����8�2a@֣C��n8څ��7�����5�;忠��A�����߻�KzJ�}��he$�Z�����DQ[H"��(X�#_x7���+�����B��,h[���>�VI��>��� �OuOާ����5υ`^!�_���;P�d�{K�t3���w�4���W�#�~���ki
>��y�;e�K��Zg�2����C*�������f��w��!� *rWQNn@��	֨@P5T��e/tV�L�)(M�TMc;�	�� '����!J'�I�~�W�?߾�|9�'ۻ�	�9�J�yK�֦^����pTgJ.��5	ȼ
/�ȼi��޾�a�]��,�K;�y�]�|�X��c�@$?U'�KV@7ې�HcV_ÿZ�
��}�hm~w�q�W�M��<�]�j��5E0k-�*�4P��Bn�\K��Vn.���'�϶�\�,��Mbeo�?�Z�.���ޛj�$���(V9��g�2�>�SҐ�[�$��-�!�^y��5�JׇpR����N��r�|g��[��,?5Ƒ�����$�map ����S>�p-90��ђ�O6�'�x���ɥ!�'����{����B��[�Nlh�}'�I'��t�.a�?E]�hD�AK�6�������@�P�0ǩ/����8�lN`�EpJ��u�pR�L��"�EI� �F曉}J�P�lo�T���o`�&��%�j��0ת?;µ¨A�G�����QޠB�H�G�h	�Q�o�N���~J���嘏���|Ů]��y��8Bc_����S,8���0�b�Q�B\��	#�X��z'y��}b�e�r��l�y���h�O�[̸������4{!�M��HG1�|ѹb�]�Rk��{��!�P��O��vtzy峍<R��W��	��Od��]ҵ
������TP&�m�FNpn��8�5����{a���)��1|Y�-�o���v��p���)~�%͕U�bi��r��^�G�L�F,v!!�J���5�J��I��l�G�A��FBj��$9�G?�� ��Xϖ8���gU��i�A���Q��Q��5�"���m��y,��@�!ϱh�H��.o5�8Q�;���*~�/��Vt=�+��'�"_����vC��[�nu��?��1\1�[��G�{�wx��m�e���� ^���^�f�� � t�������T�(��.��l,�����Δ���d3S�衂ޅ�(�${����Zo�z+2k����
8uF�}��3�������}찄�J)Ϥ�6{Q�_���E�b��B�Һ2J=��Za���Vt�H��\v�K(H$�ɇ�6�<�
ᾷ� �,#��&�����@xM��84W���?�~��X�MS^�@a��b���Cy	pϯY󠌁@ł�,1��/e$��{^�1�=
=�f�|���A��J�#QQL�`H��n���T��G⒣��mO�ey3��1r�3֘�1*�q��	������\��xƏ(�w��1�/#�	�U]/���Y>�k�$���F�T�d"�ּ�����;5��H2R@w$�2�ݢ���A�����ݥ�_���dd�%ͯT|��猉�u뢑Q���P�W��}i�)}�y����g�H�i�.��N6�Poo~K���\*�?8îS�l*����\6��
}�*%�5��:�I�#M��抪�:���_�n�%DC�����]�W�e#٭gx���y��"�|X{�룇�1䙯����ƝE��({�Ĵ�8p��\�j���d��x\��`<�S�Ƹ�O��#��o(�w�
j.%B�w��·��h�%��wɒ����}�xt��8����2#�����ҿ��}\4�e�3a�x	���X�I $'��q%0��@c$��~:Q�@�D��āy��}�*v���Q9����v�4�ky%�`b8�����Q����M����E���
�Ƒ'J-匫S�\��l'��	$�t_�05���v�kLv�>7�X[0=5�͊���R��hc�)k����W������Ϙd�n0��gv��g��U�"ZLC[U�Ǎ�I+�ywS��{�l��0�U��diE�L|t�,/7/�4k��Va2eH�}�����1�i��F�A?Lwbb:���pPͼIO��R��� uT��
2�⼶8���:��=�����"��y71M�� �)>U+ �P�|0Q,x��ϩ�̮Q��>/�ds�"1��0z;<��p͚+մ�}�y$N�� إ�D�����c��]�#�I3�#~%%���l��P%���
���f:+��S� ���H�~a��H��7��$��L_�͂ue�������y&g�>О�Ƴ54=Pu��xVuk��[��02�IPFr�¦���n2���},;o3Yҷ��ؿ;<�
��/*�쑣�}=
�l�+Z�G���D2�߰:;�'�ˬ��am�����26�ª��F�~y�����m1�����23�۔mz�	q��8�Pv��~�ci�X[�铏 �W	U�#		7��U�����p�u�0�H�?���J�n��򭤗C gD7�:h*�$(�0�1�IrЍL
�0w��0J>�+�ؽ/
b����B�� qb!G�1u�-|��%֟9O�jm��]EI���i��x/Ro�g���c�;�����Z��!("�z�;ߖ2 ��Q;g<�o6��z�G�A%A�e	F�]�k"��j>|�a�Z������U�qP"�n�;�Я�p�=䣛��%�	�W�<rvW����2�®��F�~ݱ\*���b˨`�}��Q������_��=��W�K�m�ј)�A�j��HbBݵ`���I�4����&�*c���F$ˍ>��sSHR�EI�ɤ Ź��������:���=��ֵŵ8�~�Z��FUB,���c�CF�H!�?��zo�W�)� \����|!�K����	��+�Q��<	f
���OQS�˫�����F�ϛ��n��oeB�"I���i�K��J͸[rD%@<�0ϼ��o��f�d�2�!ABce�t�R���!2���E1�d��;&����3������I䴗�u�Q�i��h��H��Y&�7�\�4��r#�k6X;� ���ĭ\_��F_}X����EsL�z� �Ţ:/mF?m���,]�ޖ�����2���U�e��;�a��SHr�����B��.|O�f��=�?����A��/$EG!�2C� ����@�+C��9�5�v�+KY�^}Tt�̎���ƅ��}��ܷq�ך ��J<���@�G�����4�6y�P���=��c�\%_���^bD�l�,�p����,8-�{5���[22g�4��W)�����=���N k$�hI��˺���G\��j��2+�"����J��E�~�:�!@�&�ֻ�@q�#%ߒ�Z��QYS?6|k^^�Pag� B����>�f��6b�T�q[�A��d��hw�}ZHf9��/(L�-ִ����֬��B5����e���o��w����7�)��.aT9�gCQV�P*��1p�_/t��:&��� ��F3��0_C�1;����,>MY���K���N�>�Q7�G���lQ>�n�d�WQa}���@�ݐ�w���"0я5"e^0ۖbɨ��D�ٸ`�?WӰ�X�&�u͛#(Lz(�������}J��5��i.��-�,�4�ؿ���U`1�GV��D>�����M�Q8�.�L�i������p�%���"Hӂ̈d�F���%�q.\X�B��;�E˜��Ew�����8ܓ�H=�jqq5n2"���y�Uz�4�_��������t�n;<����P�e�a�_H���xVʠ(�u�΁�X؀ܛτ���
e+�e,��袊A���.B}�/-�{ݭOi禎���]�'N2)S!]�u޺���v��;Dj���k7	T���-u)�q�ۂ�C.KKL��)�&j+w��H���M&,���y�ݦb�DO�Mm�؍���&�= �Vp
�� ��y�і�'����hIy@"��a���+�&�t[���V�K瑽�F؜�N�<��CX&N�J񵨉�LD� y��R��p��>����3��1<E%)��Q~����������HF�:�,��&�Q�O����騕-bj���w5��H�׿����n�В��s4���RcK�b���s����=#Q}+Q˻y@t��:)��	�z�=�:��}�#�њ�K$1��s�kj�U��p��kB�?5�p��'|�#8V���l���7צU3''�?h��ҊD~!���'R�A�e4]#���z�,�X�9���!�c����Ww�^��-�f�����Jb�rS_�C���Aݙo��X �����Z�b����yֹ�%��Q�ƭ)�'w�%�2�(������퐛q�X_�Pt��'H6�4
��s��{PvF�*�>��#EA鱓���%���[���Y��UΐJ�J(�^F�׫����(�9"�.�{(�'*����x�,e?^ �g���l"
�mp"����Y�v[�S�v��PW��W|���r9�Ze.���y|��J�¹�!�H�G���)�*��_�Տ��:<�/UpR ��e9S@(py������(yt[Mb���o�o���-�q$� _�Gu�w"?���a2���Ѥ�a�Į���?��XP-��lĉ2���M�-���w�ߞXh��d����Y�!���6���~���p��c��7�*b� $�8/��;@S���P)��Ű���H="��t��e7��؀__�^Z򲘸@�6�Gܒ7}ޡ״-.J� 1ULJu�	td��Cx���Q7�i��O$������R�c��ӝ8A�<�uV}�	�P����H�A�e� �]�s��vJ9x� �@�`�4	�ׁ�Hr���~�[a@ #\Oȹ�"c4xvs���Zˌ�"�/Wo⬿>�M�`��d����?���QF��2 `�å40tm�he�<	�j?IҲ����8�����/��z�����u�w�G%�(x� f��8���iꮇz�F� <���ք-�W�1���$�q+��O�����ʄ�]5p6n�>1s~�X�^�8`���~�xL��H�@g%�k~�CN�#^$�N�?A���)��_�_#��� /T���dޝ|�X�U�GO7�w���6��^W�\�6��!��<r�=#w�a�
5��k[;]�� El�bj|��e�e�Fʛ�x�ũl�L��jd���҉�������
C>>d����?\ՊΕ�[�y�o�X�!:��Msޱ�J�NHlI9�
2��Fat^�A�y]GFF��X1te�wX����f����/s�jy��7�<��Z�ǜ}dW ���;�Y)�ϖo��������h��2�X��e��Oq9#у��y�oέSe�}��a>�DZٵ-bp�&Jn�C��\6�H��BIe�.����v�l����i�6���:��f��CX;��X��g��\ϓ�_�$f�n�&˻T5`_)�k2<�l	�j1������xe��(�e���7Y�
������b��)W�QɶzZ-�Ih+p���Z�	�B��y��3ZJ��Y��U������B���V0GZ�(������R��V8��lʨF��n�0Q�bڞ�h)����owʍH�\�Ѯ<2+��yC\>D��X"�����uk�����8�8��H���
wl@?$6� ��ӛۥm�^���H���i��(3%f�d�=l�F|�	R��Q-w�斳8t�eܫ94��`k�ڸQ�t*$b��w��(��u;F�TX�`�::�x��KF�����8�,��g�����B��1����ԬxR�I���kP��3�@l��*`���3W�'�:��cK <��) �'����!�c��-l=.q�kÚ�����Y3z�aD,Vv�E�vى�_�#�oi���+��)'��C�T]�O����Bț��5�sj,���Il�iE6KQ�&G(@ߜ���锴�* e�w�<v�zq�^�f���F��'X�0��M�'��J2h��\S��H}?�ZP�A�h��j�kٶ�xŌt�P.�f
]
�v�PhGP�<����@��[�nY��{�h���� hh֞e�e�;>C$Wϐ)��Ol�*� B7�{T��Y���s���U��<;t�>�Q��}�2K�a�����*�((�<3��s�'�7�a�y�lGIl���LYFx��כҽ�)���k�-#&˻m+�����a�Yh�%j��F�BODҥ�Q���2�u&����S�@$���-a�}�f�M�@*c͟8�_�B<�Yw���a���)S��wŌ{1�[�]r��t��'jW"��Ï�O��Ʀ(C�zVb��{m�n�_��ɟ�L72�F���7��cI��X��[o��s�V�{�0�!��xy�Z��|.vu��=x���*�xF�mvM=4�H O�q#9�墇5�&��u���u�_&XG��~S׿/������&Uk�~f��	����P�:V�q)	��2�e���{�ǰ�D�nC`������b��2{b����RE+�k�
��۷ �{���.��E�O�����D�W�*��f���n������,���U��`�!]W(�LH�%Z�����}s+��4�[5�32�7�w�.l6+�P��{�.°��}�zo�W�rJ�]:U��%����|�G�y/�U�3̹�MP�
���}?ݳJjaIu�Z��iס,��nQ��9�_��@P��;i�ւ�/�h@����O-�~��j���g�@B�/�kf&���2'G��E��5��e3�|�8=��IWc��m�-x]��8j��F\��{'���W-�{]�/%�_}h��y�1��] 2;��W@�xȹ����!?I�+�[N��X�}Iw���7�|4��D����8_���j�G��
m8 U����D}�y��
E ���G?�J�=.�P�6W1�0�ܰEa��٘K�ңҷ���PkH(��� ���_#���3�^�ۊO,��(2���u{ rO��3!H<�%NDPUz*��yc���<�E�P�!���X5��A��CM\���Θ�����W�{N3�����Ǭ,���Lk*���@������Z��X�}RKu��9'�?���gco���bʲ	"������6=C���B�Dfe��	"���8��j`��Y�������c_�ص$���������`$�E��
x�����<R��a�������|z��j��"���,f
7�_m<�S7~r��𝑻�9M�(�)y��\�Ԧĸ����R�bl�&sƷ��u�~k̚Q���S��P�� 7����2�J:�>�.���2x�,hr_%�W��1}��2�m��`�[�+�u��1p��uѢ��l�U�DE���.������}���D-��w�:���0�>����p(1�S�$jr�sų�h�Iq�T�L�>�-�QW�)cّ#���n΃��Ǆ���e�[��'aPo ��-P��y���LK����`Z���0Ş�ؽ���eH��H��M���oB�JUƛ��VV���1Z�4�soW����;�0d��wzh2XA�!<�`�>]F����- �t�1�w#��U��\����(�ʢ��I7�8~ޢ6��,�e$����u
���Zb�o�|����膁�,k'�5x�
��si��A�?H�p&���I�����@ݮ���`c|�{vjcgr��L�G��)�@��p����������|�J�5��ғ�c2�j���YQ�T��;L�ۨ��#��U~�;�S�U�O�M�k�U��b�E2�7����!7��3�ѩ(NY���\�3A��+��3v�v�.�i���㬂$Q�E_�T#' �d�D՘���O�x0��V0��09=>������`��bz�*]�����*���Og�����>b10vH�v�e��Id����4�*�w�
Ә~�M/{2�wh�m}Ze8�y�W82^٘K����ƍ~�IͽF�1�grz\v{�Ψ�'�sd�P�
���	n�;sr/�E˛�X�MH�~�&$�	>"��o��Čx��78^�l�E�+bq:��������T��(��ἴ���$"�iWʜ"�n�֥�B	�_KĒaΎT�}��˓����J��r�DRiF\;��o�����j�����m1�=ď@Y�䎒��xV\,��b���Y|�*�L����VmX��T��� �����y?H�5�P�7Pw����c`��K2Ɖe�'��1�� �0��i���e��.�k$��,gN:����$���ٱ�O-_
�����46ڵ��b�e*�g���?;#4g�凰�]�Ib��!��_�~�,&��V����2�X���!3]SF��{��l{mI�:$���")\U,���An��u��/�R0�d��������j�^tc#v�(�� ag4���&X��q�q�=!���q쯚� �L�o��w0-Q	;�k��\��6C��2�V^PoH�ɰ]�B�s���kjc@>�˥�Ҭ8����a�Cʃ��>s����=4}��T����,�8u�G�sO�e��
(oF+'(��\��i����U��T<}`����7��O���LG�����+��/r�Ny!o��Vf�|�aD# ��*���a Ҿ�1�L��z#Z����v�e�����̐�8��GO@ŗ�#���+L�dE�Rו�L����X�� �q`\0@�5#��8�UHr�(_�mB"q]B���R+Ԍ2A�;��6�DN4P`�:�[�W~���תI���o{�ϡ��x^� �:�U�T4Ǽ񚴔d�_��z��a�Œ�n�1�UTv�ދ��F� ���>c��\�Н�aNR��D��m� �5�w�op��ֆخZ��.qh����t� o;2ݻy?��a)���kY� ��|T���<�߈1���ty�������	����O�B����%��h
���[dՓjTl[�)g��c���7!����|CUs�}�H΃���%^tX������:o���"SGZ�!�)>����^�r��L����uv~�M\Ο'7/���,.��E�j��кaI8{�h�Y+�*��i[���5_��\�S��M$-�KB�V{�Ըf�5�f,/���� �"�����z|1��3O���aRة`��ۂ�D�K��Ze|.:�i2���~�w�x�1�ݛ,Z������,-l���.*׍Sd��Շ�Qh��;��+Xf�Ϫn��5-��m�8{����u��?$�6�x���i
�I��o�/��e^ܳ�!��3Z!�����
�0�܁���Vi�P�EЇ8yγy�0�UP_@�9v�R�T�(��5cW��\����D��+	9�߼��S�-�=a����qљ�-���hA�z5�7w#�[�^�֔���@�_/���n�N��Z�:���澿�N��Ǉu��*_}J�̚��m��f�m4�~�Ӭ9V��ls�$W�=���4s�ͅ��w��l��	S�~ؼ@����h7�i?��5�����W<81�ii��s�.*�pO�	�G��?�̻����
 /R�5�3�,����ת�<4��͊�;G{���[�멶���r�+�0G��H��{�/����_�DW���
D��hZ�_i*5�yD_�of��K���Һ��ʖ֡���������4��O�ט14��
fg���zrH�< ���Ne)�u��H�kO��Ϋ�l7S�@�7��y����WX�٩҂�>�r��}��S"����{5�@����{���*0V��yF��P���5��6��[�8��Ϟ�����xM�����W"	)��l�e�_z-�i��>�$�����E�� E���.O��<H�|6*rʚ19X=�ƑL�V���'f��kh���ma���_^��o6N4�A������?L��7}6V%+���ֆ�[�3�
��������pot4'���>bu��RF�&`�������>��\�zG�,�׏�_q+�|B�Mѹd�5�`�6v3G�[�$^�_q�#���t�WK+�#XL/ڇ��rH�;�~l�B����h�ұM��[R�x�NI�K�/�f�\���8�� ����t�/��Ɓؐ����������|C*��r�D��0�d]M�����)I�X,�Ֆڴ��}G6��(�U����l�qyn�F<�ت"+��>�J����3)��y�I��Z��P�~�M�Kp�o��`~��D?�:5t�!��vZ3{����ܳrr�9�����:��F�u�����I�}�L~�b��~llVl=�<���Ӣj��*��KX�HD���P��	�5?�).%d�"�CM�
U|�����X�&��	��F3�p�O�I�Gjv��5o�͌ZHD�e��R:�	�e��Q-z-52	��C�H_`�4���~�M�����O��e?կ�H��BZO���Lyꌄ��(~&�V�Ĵl�����=�sF��3Z`����ݴ/��5�J��8l �������7l|�%R�v���6S�D�0���������Ѵrg�s�r $/A���P��W`'RZ��P½m��drѵR�=9�4l��_�|0�7��|eHF�V�^� �ġC�ب���"��6H%(�h�L/�������������'��G�SD��pwl�fǤ@%F|�D�l��!�I߱ӵ��H}�M�t=
����Ե�ED��,��=��X��v`U�'��7�
����g˧jd��\��^Ǔ��;Qy4����9Dl{�-�B��$��\ג��%lr.V?>���H��~��"$*�du8%�H�����o��a� �{l�u�k���w%��4f�+�Tx.͐��,쾿�.��-�@Ȑ���GS�Rq	Q}"T$�|�)�͗M��!��� �Iϫ8mh���E� ھ�~���܄Pՙ�ڭ�*��������U��$dl�s�S����N�x�7��(a�|�@N��f�v�����?��pK���(l�sJA����	�:38�XRP$lǭ4w7���٫�/�#7�;�C���ϟ�{��qu��b�IO�H�{d��a����M	�Q���6� 17�3��B�r e,N¢�_�*� $+E�0'+�j�	��d*��sڻ�7�p�����ΟQ[[�L{��t(^��1�S���B���j�꘧0Y��TZJ��L��1�kV��9[�.�Qr���S8w��ןV=끝8�L:��KBo����G�H�3�cl#����bfաN|(�ۛ�L��L�ם��fX�am�O}B�� �^�+�&P�ġ����a��R�Q��q3V�.�a�f`���%��%�l�ܦ"�Z��`8�\�l���G�@�Z�ee�PH��V	���!��j�A\�m��N��v�Eڼ�0�j9�-)%��4�	׊�BVڽ��7� �Í�[�V�4�'��`>q�I��e<����#�/.�-0c�v-FF�Xݷ�9	���.t���ϹRx�yg��]]��䶁n�7�g����s���:��O���㉕T]in��B0k�*���f=���1:ĺ�J�X:��yIx��c]�LT�р^%2��d��+�n1�ڟfN�F��s���;�c��mo�Ϭ�,\�D��.�+���Ȇ��/mCzF~���T˞���9UJ�A���W  ��Q��E���r��ݤ1�.��n����}�<^�.�ԑ�_K�#�jVRݮ��t�a ��8f1&���@ZY]!�,�N��a����܄Q{��ŋn6��B��6H?���A��!m�zx�+栣Jc�o=��'�؟��2ŅX'C�a�gzP�ֻ%��n`j�<ΰ�VwS�x%P�k�d�5?io9����G���w��]yZ<qi7�K�a�Y���zx��E�ⷍ�=v�h�B�s�oҋ 󺐂���m@c����i!��ń^S=�:F��fl�����y���P(DJI	Hpiί�C��<�^ݙ��,z�PO��K����
ee��Rk�����x�����s֬��32�*�un�	�S�Yri_:�'vV\ɦ+z���p�8q��e/��'���b	f���C��\q�P�p�����Y��jAp��J+�q�Ğ��0����K��1�1�Z�E��m-FI'CU7�'߱��=���ɖ'V)�C��nv�\ׯ��s�>H�ް��$ɰ�pڐ&$�I|ݡ�{w�Ț
�P�V��LwAz���K�J���}��կ����6��#y�����q�]y��d}��@�S�cD��C�W���*�0D'p9ڞ�\�dÓ��D��'7�
Kd磙�X����(��m�`��r���n/O8�T�P�&q�[s"4R#ʽLk<t*ߒZ\�3^��D�b:�<,9�&3�PH:�g������9��ΰ����ˑ�P���H������t~�e�������x�I�����H��X��È�-�EIA|�����ꝵ�?ݕ5�Ae���I�9��:�5vL�A�x	]g?�Q3.�
��o?�V[�CC�ZQ��U�V�rj�3D1�`yu=���@�E�s7���Fܚ��\G ���_'���ir"#~�E]�@ğ��b��*�7�Yی����5�o�2Q�V5o���m�b$��>r.�/H�z���u4�=�5[Q���>$��r��o��}!�7������i�-F)M�����9�u�����<��f��8����cᦫDZ����Gy�X�љ�������ҽ�k@�R�Cr�qQ�P�.�qʕ}<�gdַ��!�l��A>ՙ�-&@���Z�wE�Q�m���j{�����.��Ϝ���0���(���>�I%�tA�Z'T2j��BhG����������EK�G<�CP���q6��
�s��-�u�@*)��O�g�j�>���;����We4�J�dR�^�~?�����z��F�.�$ñ��{n�j���*���S�3�#C��0�}��c�q9�#y�\K\�J�ѰٜC�hYmԓJ���/@�djJ8?���H��R��4��_f��޺fw+�|��*xX�/^���b�/O�������e(2gߜo�މ�b��E�|��*.�&�Ɩv�uB����^��*�žr}?#���?�벱���E���qӅ����@u�%Vx��d8B~}���7��{�
�B��f��8�a8��l�%zĆ(��f�x��V�HpK;�;��ϱ��<���G[[�����2�7�:&e>)����s�n�2�.$�Q�JsB�@��`�mj�9��8�h|����:��Cb=v2-c���\J��)$j$�*���u�5�,��t�ڂ쟯p�?n�gs���h��� 8��n��GV�T�W�F�XY¬ϟPc�� /J;Ύ5�uN���L��(6;XRLeo;�V���Ϣ��d�V�3��5�e}59D���_�*����@�n3)ǭp�Z%�z�D"0?n���K�˓o��Q�p#	����� f�	��Ր\�j�k�����3� S<���L
�+��g3�'��֟�s^-W��?4rp�0�x$xk��q^��G��7X �M'�AJ%����Ǳ�(�a"�W���
�ڄW���Ã-HB�n�(4Z�u.��T[:��*i��~:E.콦���*��ث=ڦv#DlO�iX�����6dKx�޿�cP��Q�2�4d�S�F�@�+$���c��`��/�@�,N� #e`">U�S�y�ZU��=��D����iҸ���-��JC ���z�KiYJ����p����7)fD�����:��:���d<�&] �ߜ�:&p��#�p`l3X��O����{�MX�����pރ�|��]�,���3G������S�*$�Nf�KD��&�"��i�6r�;Z-N|z��]�⮉V��������c�v960�Ŧj�A�'Y0|�� mY�L� ���¸E@A����t�[N3eQū�Q� c��B#��͋'�&9�b5��H��-�F���4��k:: ��4�S-�7 �i�⃂�ގ�Q�
�嵫A�m<�lת��!����I�h��r?�o���f��	P!�@�n�W&��n:5n�ݐ�G~P�z.����w��>����XevȦ:0�]���AF��.��M�,�^�����uyW��ٓ h�k������[q�����2�Қ:�o��/zM)������"�pgk	�J_�V��~��I���}��f=<����qȹr��J��-o�C#��C{����kI.�u��X�.I0��p���¥"sv�O&+�����	MƤa��#�0�>��nT��B*���HS\���춅�ه�xu���J�����!3\���h���6C��V�.U�J'vi�a���,:����G�D����p���?i����W��`��|4ܨI�>�*�>O&�#�D4�]��~���W� 	��WK@�7��Ú��d�#K��㔸4��*��<MM�3��c\z�ereC8�n���D�1�<ab��	=,槅)��`Sg3~v���4*�b
h�NR����s���0�{��1Eʵ|
���s��[f�ŭt�$N�J]���F�%��/�S�0,UN�\��v��)�~�������l	�mZ��յ���q��`�	HfCW�te^e�z�;N0ܿT�L�r��2_���&3Z�/�LX�̆.`�kh>���{�F�1����m���H��JM_����V�\�$N�gβwp|�8< ��-�
��H����:������Ķ�rQ�&����1�Ow�!���H�����߷�$D��}�
�b?w�#�9J�[ xG[��#�W�g`�[~�{���mɪ�]htջ#�������� �ė�1rHW窀� K#:��	�g�	��pG�kDI�Χ�z#�e���a}^dă�E|D��QU��nR���"7k��68w�<����	����˖w��&@!�A*C�;���E�|}f7L�J��Qn�����4���A=�#&�+а��D�+�=>D��B�|L�0q/8eǦ�΄���$��!�|�'F�v��3yHq��]w�s�x�.�o�4��`���4�>(����/%�3��i1����?���QU�[%>��).}>��K�B��|�k���0EA�s�թ�qs���?�0PS>fw6t������bf,������[ǧ6������ʕK�-��cD
��?#(>/$��!,���LӦ��=�j�~z,B˕��Tvh���Ό����g��2�h{3���x����v�Q[��춻?�oTL<�"�@q���R�}���R-�v�����F�P[3b��i�2�-��������Π�MۣO$�y���PDy�?�+rd*~ ��#�(}�Ĺ�e���֫$z�ε?���04��~����KBz�K��dkH6��Z��P�j#>�]f2�rp�os���=HN����WH��STY�"ڤ�?��a��c��̌Ea�t:F�i�WT�[U�UÓ(�'��袐�~,�JBr����ˀz�wU�ҧ钳;&�T!��1Ḓ
�&�A�?G�?9��P0�h�U;nx�%�x��Ko٠�.�8������ړ����b|uV��
+zZ��Gˋy;
IS�U�ʔlP��ԭ%UO�sC�~��leIS;��`J\�.Y)�:��$��ϔ�T��-��x�B�����u��m>��dE��\����`W)B:F->�i"e<W�,YX'��4t�?��!.?/D�Jz��"�����`Y��A��8J�SE��1�|Fw�1菣��׍T�ׯ�1��9U3��"���-N3]�9�uv�kiet=��O*+����=�E�d6{
���m��:;������a��2�̜� 竩���r������y�6�T�1Oj^�Zg��q�o|�9��� ��N�ڛ�7�ɞڂ,i�ɴ��"�+�%�!�w��2�re� Zx2���������k 4�Pߓ�|��Q���F��Ȳ�RL51��8�fa�Xa�etS+�gW���#�g	�^i������D��Ö5t�*]�d�@����ݻh.N���ԝ/��H8�j�ym	R��>D-�B6�ԡP=�@��T�u*�TĲ�жK]-'���
IZ�d�OЋ�!����w���t뵔g'z}�"5�w��$%e����i�k.z�_�~ng��a5r�F�JԒ�h��Յ���	�uSG��=p�����꫕�f؏�JDb9�h~�$~�|�qH/�º�O�Q|Άl]/��V�i�[0������͵� �W#�Γx�LP����㙜Y�5�	�u��eN�qw��)�+��i$��Pȧp�]0����nk���y�������3	�	5�>�Y�V�R*�F%��:��78j�Kw�S]7[���EED�q۫,35�9�nDO��!�1,��9��K��{��j�;[e,O�͜�G��mh��f[��:�ѕJՋb�F�pf����y�iD�aWUߵ0�RзgZ��(�,:_'�9-e�&��[E�h��'�̑8yσr���$l���7�����s�}u��YNF�E�#5�:�>��I��4*�|m_4q�Z~��[����7�^�0�Q��t�'��3O~xV
��z��AA���}ou����e�%�u�b4�SaK��d�����pT�7V%?d�|�7d��r���@;nY��o�-�R�S�&�����D%�!*SeH����{z@�Օ�P$?|OދC4p��#��.`�J��蔟�)&w����^*V�G�W���!-�~��̚:�Ac�+����C��ɏ���r��&��5k��;6���o��RhT�0�\�	��LE���zlcz�SY���:�W�����_�D����#l�nq�=���������CW� ��mޙ�T~��P���FF�Ͻ��'E�>~Om���hLC��:������C��i���"F^���)��Kd�&Pm����`h��"6�F��3d���|]

�Fr�Nz��d�.cw�tI��>f��'�6����k�W:�u�m�fO�䢐����_�_�g��]h��t��u�P.!.ԬZ��x�s	I?�QT��4�� �w�2]�c��qP{޸k�>�����Ƶ�:�@8�4���ٿ�6JE�J���AF_��k�̤�K��Ծ�EmJ�� M躄#�BІN�rfd�D�4r�1�>*�c����(��9m�ry�����K��b����\i��7pd5LG1ȍ=RQk��[��.�3>�x�QC�C%�0&o� _�T������}0�o��~���Z�`�����=Z,���A;�&M��4b ����'��k��z3-��c��ps�Jl��4�3�2�_�dEb3M�	�/;B�68`�пr*V�[�.M���@i�gz���j>~]�v�b1K��d��KM�>"c��Rc�q�SQ1N�H"(��ײt=���PT�֡|���"�8ev��{��D'7ռ\�g[������H[�m��Q'Z��.6A��J��QS�	�����-���n�N�W��@"���d�,1(b�-�L"Kϗ�[s:N��0�_����j��IʄZ�2�8�����M��# ��[����G'.��f~�`G6޺A��J��|�ڄ�J�����Y_���`�۵�$&g�C�\hb~��xz�.��3��;J��*��X�qj)r�<�>Ml���`�g�=���+�~����1-ֳ��q|��(.���������ble\B�h�2��ĺ�\Mw��jҒn%��N�.+\�C2K*�(�ߙ��b�֥� >]��b����Y���]d��w횎ন�ZM�j5���J�b?X�\����ò	yd��Fh�)㵚5���4�*�5-�d����v=y�|��ٔ�m��r�n!M�1���.�v�B��V*�i�'��c�t��h�-j��o!���
/�-%����9��Z�j�=ʾ%��P������L�)�����A*w�b9�ϧs�K@�CL��+A��x[�S4�.Ғ�c��"Ӧwo&����Bdv�+���X�����LWW6�F��Uv��m>0�|,��\��:�$A�oK���Q�o�+�h6�{?�)ڤ���h��zA�h:��*K�4� �#F���R���FvGK\U�K\����!ӯ�H�?�M̜V3$l��r7oеoJ�2fN=�*�����Q�iA�3�r�Zap�H��
C��K֦�BM���-���TQ�ʜ���&�:�$�{�!�9�%�mMr��-��m�ʒ��%����!L]�E0�x���e!d��F��4�?i�s�\�T]��->�Q�5>Nv�0��dW;����)�D��O"^҄ѥO�@��6i��g�&�n�D��qq�8�;i���J�.)��q�n�e��J�eڑ���p��{����;�r�Dom2&��]QƳ$]�����=:*��Pk>t4���?Y����!�2&Ι���[��$Z�������ρPC�ج(K�Z �/&}
��_�pJ���`t��A���b�X����I�������Z��g�R���$�O>�tU}N�mL��i�yG�����`Ȕ:c�Ë���E�z�0Y�[X���%	W��n�%�mb0��1IRd�У��2�e��	�����;��f$F��@��Kj�-[!���N�P��k�\,A/�bl3�ǛW_�R�,�ڌ���֛ao����V�D,&I������-�(�@��|E� z�,��R�_�.�Yo�K(s��y���?����gK�P.��"OX%��Ʋ:�U��o$�me�'mh��� ~���K��jl����-������r��P>����ʰ
^��l�^��h�d�����Ȝ���g����4${W�2�D�y�����E�H?��|n�aCsL���WY�	��=����oD��˚쥫bd^D	,֦�Ux�Q ��h���^FJs$\���F5Xh3F����=:�}��[W�z�����������.�s�F,�xÙ��ޗ�	~^���#_����n�U�$�E}Y۠+���"EQ�1�ra���� �1A��z�C=�э��֏#�`������(Kᒵ,ԉ89��E����] `*�2�}���7>1������/�]�_��%���S���g�a���e�sm\�$?��v^�O�9��d��>��5�If�PW��R�/3F ����@m��0��fH�k�UG��d��E�M߼2� `�����h�f�Z��:Z���bN)� v�أ'��DY8�%e���^O����J�@B���Io����������Os����K���XH��jx~iGٕ�?ʑW�������ډ�Rb��P�m��/_ϗ��;4���(`C?~���	J{	��z�nꮍ�a�Z�~����*�\����&�z;j�8Y�+fep�|_����{@���>'�F�� 0�D�{2�Y˫)P����)K�:4ׯ���x*�����@�C� ed���J�d��8�~j�^P��K�NW�� >T�/h=&ei{�R$�M�������;|g^e���6������ pT�؈�p�M��2������prl�d������`�2&;�#)���GCn<�F
ܨ�J�O�{��nî1x�K�=��UT���O��ֻ��(7��?zF$2P��O�v=�\?��x�q���hq�P��kp��#���v��E�?[�*�_~�4~s`#H��h[c4x���B~��,w-8{Y��x-ҩ�)�&�+�>󄱵����0lPU{���Àx��Z�
�!��]?&�3��j�Y��.#�����O�*\�~z2ґT}i�xnE�������%������B�A��0�>CC�6������"ָ2[������C��&K-��nWu���;$���ȟ���;j�}��2���oϳ+��N���7�v�v�E����YeY�~r�9����T��,�h�P�xF���9��e2�P<�͊������'/��i�0�
�ҭ���)��D�s��y�֩ �
�Or�����|6i8���)��K�i�{wX[$�|1�y��� 
첫���j�_�zP+�^u��ߎWʐH��h�q�Ȕ�^w���"��mp٠e�s��I�(Hy�n`��yb`���b �X�5O� f�j��t~���^JbX!Vf�/�O��6`���*=�R.��h��Bs?C�*`_1�b�s�P�+9ԟu<��;��c 8s���!ԯ�tx+�d�;�@!�H(��%^)��SZ��Ģs�@jx����1z����S����P$��0x���B֪��\Aq���F�4��4�ǜ�7}�����.�rJ[��.�(NU��$6��W3�S<q>8����{<a��+�w}���AO��S�]U�����O��6�b�l�b�1l(6��s�Ƞg+�sγ~q�3�?^�{�,�����/�K�U`i�YJ��R�,��Fs#�m�4�[s�k]��1;Ґ�5XF�=ͩTэ��������@�����-9���6��Y���е{�-oq�*I�q@e��T3^�5�$S��d���V����JO��7T�!*
wT�l�G#H���q�.�����.�T�87������痒�L$��)�ގҸp��3C�����8��CXJ-,P�]ĀoR�T��ˮ��K|�N�;�Tm^���W� �-�/P'e(Z�X뫈�I��� ���DQn�{��m�$�kN������|.���58�2r��zLa��Q��e����T�*���4�;�H��J+1�=5��u�k�K*lvaq��2���' =�M;����,�"�S���^��VHt�"��J�C"��VQ)�n��x-|��3�Zr�_R� id�JEb�L��s�p6��c`� �?M|(>�8X@��G�#��>B}CMpD���a���At���R]PB��0nϬ2�P����,mH*���o'�/;�\E*颒@�p�<B��h�2�I�v��S�ڶ��>��C��5�HHL�p���aGG�n~~�/�倄��H��|+���}'�Ԟ$�3��D�wQ��2���g���`Mi�ƃ
���":i8ny���Q\�V���h�CH"�Q�9�۳/��^�8e+{^��=���3{���K
y���^ڜi:{oG�5�%s*����fW@�c��ݙ���t��O�y��'���.�B�b2��k3lg�w!�7N����e6��4���7[mx-�_*l,����|��8�V|��Pu�2�o�\'C�UJ�5+a{��J�:Ŭ]�:
C�x+�DXzE�l�Lݬoh�U�w67-��Ƥ�qp�L�].x�͇
�Sp�c�o�s�ë�P!�M��s2��n�X��L���Bvڅ=��$��/,�X�!��)2����6��(�%��r�Z��'�Ķ�jqVK�A�J����O�z-�7*�`u�4�L@�o:��^�8�SGJ��P�7�O�F���t�A��t�R^hP?v��{tbX��)�÷$s��G$SR��}( �'^�Qh0Pk�^��ʙ��gUF��N~���rw�֋ad3�d"�~g T�0M��繃�3ƪ������1,���44yY��?�\p(��>���yBd�pO�(c�K""Z��}��5�F:��LN��%s���+gh��B
�
�X������9����Ac�?�KYQI8����)k�3����i��Q��#��:��^j1U����8pW�t���ҫ2%�z�����E�im׈3s�S�RF[�:�)�����j=#�h�E1X�\��͋����ǡ��O"�%SBS��יഺ�-���g���ǌ����/"�) TZ��2��^����ޙ�����i�=]��[�L?x���E`�'d�>��7�k��r����=5t���S���1��jL��!��4B�Q^hoo芵O�};;F���!�cu�#���\ݵޢ/Y��c�(Z) ��6��5 �eK�'��r��Ao~1%G�z����M����AJ�G��:D׎�B���t�tZZ1gJ v�P�����O��|�A�Hp�M9.i�T��,���62ޓ3����X�{��(����"��+	|��q��'��~�e0�R̸�,��z ���u�%�$�k�)�9�04v��п��|w~'�]���q	���cL��v�z��m�&;uH6=vnZ�{j�z�uΤ��u>`�o��+����iplf*�� 埋�Y^ �Kfz��K2��^K�F�Ls\�3�<��	_��z�4j����M1"6P�f��(`R*�a%�NQ9��&j�zR��=��^CZ;.���������؊�0#��H{R9���PR9�އ��n���c��O�Dt��i����(�G�f�ձ#@pu��=�b"\7�{���+�4l �1�vk�Xى��[�oM/ގ~e���h�q��0RvD>�pУ� ˧�%?�R8��-����G��}*���!>���3�8�����@`0�`E<LRfx�'I	�s�p.q,�Ѩ~�W����[��v�=��+��_ 3��[�	��A�($�iԪ����w)35��@���xG,��uHmzm�j7؀T�ZR�S��ǡ�[��N�{P%��fE������"�v�w� ����E/�%���ո}�R?9t�u�x��k����S$"Z�R�?��˧Z�g1,i����������4��oͰ���Hm�s��5Ct�>A�j"���O�8f�� ��z���,��m!�RP��^�]��#�
�fK���\���B�,�x1����}����WI�T[W�*.�����/-#�kT*	���ߊsTQ��=��0 [d~3&9�%�N.3���i������#�Մ�[�}Xܰ�<~> �}o�W�f�zX�	@��lB{3r�&_Z��Ko����!��H�/�Ai�8%:��U��^ƯX�;6��ڬ��E g�U'F��U�����d��p��9�Z�}�o����DN��m��j@�v�A��c������W)e)��Dw�+�UW�1m;�#UI�c�'���D�Z5ʵ'���T���G`��I��Xڄ�}��|�v���2!,A��%K�B�5H����kV��>Q	 �L�biynaJ��e�o!ʍ���-��DJ��%�����])XTp�e{���h|���{4_��4�+��àQ3���f���
t���7C$f�#48=L}и�ѓ^w�z��*)��lj�A+q�H/�I}�3&�~�И�Ż���[��`���C)a��+�&un�����y�=�&�����K�S�+�V��ԻG����X���q�k��n����9I#}�q&8)��zT�/_�gae]���vN��5!`��ߓ郤B��S�JQ�L/ַ̙^�\���S5���'e(�n�����y直�[~V-"��⾰��i&c;��_��$�K�ҠS�=�N��J�G{9����?���'!?��.nL��cE��X��ǡ�9H!9K8��^��H.y�����IF9O�v:�qo�䗍X�p�G�1 e/�=�=�i�j�W�y ��5�˓O��&d��|��f]w�*��P��?�Fs}P�?����ح�,��/���6�#[��)�w�,&��"�0t#f�2�2=a�;���BIY[?��u
�)��~i�&���hh:���g~qZ�C��[���D�WP�V�8=�ą�Ҫ҅z�%��R���RbyV�0�m��:���O:y�U��.
qu�6Nً)��	��[g^���`��*�"�l�>8��K�!��)�>�[����Q�.�s�#�u����f'���$B�[�ڵ�W��4I���޳�����w���.�r=�@��^���'����ȭP�4��J������7���s�N�
���Yg���pF��\��:�~M�j!�B�1)Z�<0��ٛ��gNUX|��� ��-�MO�fb&3�L��eIZ���ZO�t"w�<vz@ŕ`��X=�cIy������\�+���Q�\Gk\'	ǲ%����xOZ���dDy}��~~��M|:-�ʤ.˿aH[�1Ea'����|1�;B����)�7�sE�Bo2G_�ס�*��.Pث�������>]_��Ŕ��!<,�� L�VI�-W�3E��u���$��-�6�<�_8�7Y���ع��"�m���Gu�C�v�5�
�1@�Щk�+��7�U�6d	}G���Z�^'c�2���.������^޼Vt��v������7[N9���T��ē1�T��!��m���ܠ�Q�߅pj]�R��D�i�ǯ�����3�����S��,����ӼD��D0e=#�va����:�c�c�f�Y�N��ˠ7t�1�ӮMHz�D����4EA�q�?cU����X�}e�yiH/��q�q�e1Ju �P�+7����U� �ZL~�RۍU�I�J�Ӛu����a@a�B4�x�h9آZ��/�!0����x=���{x�xmRޮ�jN�-a��j�=�:[��w�7Do��k��7���MjC�g�?_���s�S�3����F<b�r �+ٷ�	+3є����vhj��K�7;Ov�y�o�k&wo0%��cݤ��ɼP+������o�����P= g���]��v?�,�d��6ۧ8����$4Da}��؄��2�=O�2+O����6����.Z�|�cr� q�i+�o�)�ɹJ�A��7/�i2�/V
|��_���PƩ8���lGϔ.����g��9��$g-�B �d��3��Ҫ�pM���qq�Yk�c��s��6�ScTi���d��U�^}h_k�l����^Q�;|X8���V�[�ӡu�L��%˼��xۚ��$W��2�qhrz!�@�t�eԱ���>?�թ�
�N�]��&�-�Ӱp�堘&���+���_?ê�_
�q�@LU����f��ꂋu��:+u-�gwN��aA�0����S	kd�[��wYiΰ?&ӗZ�j�ւ1��S���J[n�.S�%\�6�#��b�U�F��b� t"�џ�Q�	f����'¦E�� dW�qz�Pp��W%
y�3��j\
"�����j"�Ġ�~��n������,#�eS~U��<�`z�:��zWBA�!��A<a���[���D1ȋH��R�h��� ������4�T5�|�d4�Zg�	l��Oh�Fx�*�Q��F�
u���9����O.S��>!�����uҬ}�TfY��~�2
�F�+���~1OPϝ���+��;���3]�~�<w�=�xK�UcL�k51�jb��$���+Q�+m�A��Xhƾ]�~��EݓU�l˂�*�(�μ�V!h�^6n��M} {�h>�>p0\a#�kIoT��u"2p�{�kDl��S�ku� 3�G�`�˫�4��ǎe��ڛ���u��1��i�>����h��g��΄ �˼�����DMʊu����E��m�S��р�� �J��o�^N�}�>�+����a���",�O�����ʯZPu9���-��l&sQ`r=�w�X���$�LV����m����.���?�16�j:dV$$���
Z���gρ*�����S?�&��`(����\�Fn��ҳV-jW�/i#�%j���fȢSO��b��9�l$� �om�����淣��Lwb�����x�H�L�9��b�nN��˨D��w.���&LM:|�����Z��2
��C{���=��g0����k�>�$I�N���M�����(���3�t�u�M���:���^A[�G`�tG7��H�w/�W� a%�v���e��m:�M�${�'�>���҄k3����2s�\�F��co��h^�
fS��C̼Hk��8V��H���j}{]���y��{�,�OX��-��	���h��T��6[�BН�ӧ�c��6[}�ikT���,%���tx�������<�"�?�z���%Q�/L��a{�v�J2��W#d��3yO���z�/j�tf9۪;�.���ɢǓrq�^{qB��uNA�OTo7�#������7��$�k,乑Mfɧ���,�j�:��Y)9���c��x����LH��;���@�3����;�Gk[�n����2��4�|�A	��z�+�9�gɔ��tj�`�-�6A��dQ��u�b��l�C�h�B�m���F@5��I�o�wv�A֥�bB�6��v����JJoj������8�O��Z�����$�B�<ȭ%U��'� 7T,��Z����%�'% �0lM�n����;�֬�?�|quO:HM��'P0;�g�⫭������X��_�Epg�\�$�6�Ac~,ܺᶒF'����x��)�\Ig�	�T!��:ˣ�a����k�evt8K>�yu�����b*�
H߸�8�Fy����h?J/��D'/Pd�w ��� c��_�`� ��X�yK�,%2o/��Ư6�\�j��nRPU'K�t��TuD�I�'�����0�ݫ]������;C���1��-֝��^���Vw)	��Ѧ�:�Q#��VW>/~����㵤'�b�p��`Z�J�d����P�O�T�缅��Md�ȳ���TR�\�y��;��s�����c?O�m^:�&;u�7b���P�:���O�F�i���KMmp����e@�$��^x��s���V&�Տ_�^�Ck(�����˗8'O�ܨ�����DZ^�j���mԡ���%.>}�7�Ƙ�>���T�����Љ�����҅St�����ޢZ�.�@�����wc�i��}��Α���CQ�Ȫ�#r��e�HY���ؼ=���N�R�R��5Q�)'����c�� *��y'��:�Kl��ϕo�c�A��S�Ok����^EKDۦy��k���~.7ixmV�m�-��dk�{���+h���:|i��|�9a�{a��cV�Q�E�aAbז}:��0�LM����ڊty�K�4�
2�M�	����u���B��l.���.U��;�j��3�>i��@�6:�.S�O��E0:n�i���{1�:Ii��.����by4��~�D��{@����͉ñ��v<r����hPh~/�=�g;I��:����+j�G@ Y�� ����y��\�A׀vF�C�gLˀ�V��í&|�-)�Ol2^����`,D�T��dPnj�Ӑ'�݌E ��l�T���*���M 89���fK��4g��֑l3ŧe�����(�j	���O	�t)��1����������L���h��-�|]��_��.�h"H5tP�`���8���4Z%Yb���i]�Ь��Й<����b0��Si�����n���S����NG�:���"A}(���M��H8��҂۠�~��M`����|����E���H��������������,#��@xyN������0���^������7�0����t����OJ�I�imN1�.;͖���yʡ��� ����
��~ ���FK��('�ӻMM3�11���z���k��H���]D����8H��j\鏵{�>������BK�= ���1zOm��Es����/�m��K�NW���m$��4ȳ�Uq��l�l��Z�?�>*�G����"8#5�	#����Ž��}��wV2Ӣ�4[�XD1��h�D�ˡ�?�a��@�VGRE���0�4A�D�����ϝ)�[~����u6?Ά@��?S+� ֡��<��Q�|,C;(II'@*�@!�=�ea��{�ٕ�n)h�y�;�&����`Z�8n���A�X��z3V�@�=��*��J��"\�5V�@����3j����]ߏY��̰T����cX)Mx�LLdn�H��5���<��(_���ZԱR��'f��(�N��+#�Y�!��R�
K�?�r��,8η���#^���\jL?�����
�a��z6�����?�*Ok�����8���~��d^���v`��H}q�A��[�BӼ��ML�T ����u���ޥ% ��_#����"�6��[Z�m���,,�ĊqHD�D�N��r�P�L�ns��/��R���k��3�����R:/3j`�<�M�<��C�iu��=OTK�/aFż��ĺ��)�F�ࣂhI��ځp	9���L�Ѧ��̥/����Sl��a(>�I���5:��������0����w��	���� �S?�JrG�8�~���ƞhZ�^�U��h�p]H��1�]먪	���v����#��{�m �V�a$���f�l��{N���7�ـ��-)���������x�r���Ɯ>v������aظ�/g�>�i�O[���6���QD-9���(�>�v�G<X�߮��Ee�Ǎ��� �֦G���,"E�I�����8�-J�݉��k�{�"��@��7ϹB�ꑶD<
5/��B��M.���.ǵ"<��}�f��.E���ȕ��;��2!r'K�nޒ7ɌO^M4@0I	��eƉ���(��29G���}p��l�o�WF1��6c��a��o2X*~[�jW�3G�#^OHQ�^gQ�uv����
ѓ8��U]y�'i�Y1e��o�#�!0����~���$x�Г2)��\�79G���sb�dV�WՉGQN4�7��G@ַA�kXh�ꏢԜ���l@k�T�q����X9Ne��;Cg����B�s_������Eܠ��Nk���G�p��A(�5��X�=����=�&���_I�nW�?��O�2�Wt��O��)YN�P���^��.o����K��/�/�aN���n��1d/U��M�X��L�:�1�z�`o�{Վ���C��R��he�u㖠���$O���V6c��O���Dbt�������f�-F�ɂ��^�F88�ֳ�gO)����wl������gԥHS�$��|��Č��~a�2=����� �������]������'\�xm!*2�$�`�����D�U�I�{���9BH�wd��J�I$�H)Մdu���|�#�w��x�k�}�g�T	������1��T.�/[:Тș^�I�4�$	~@����m1��{M�j9BH�0�j��X�5�^Z��w�VS�_�;<�W�)5e'����{.�KIT}C9<fw���3�����Oy)^<'�J̮a20+q���y����դ�d�z��@���{�Y�oɆ�&r1��/�F�Q�M��V�=# �_�mč�z���؂+sR�otM���Ǜ�}D��M�!�G�櫹n�ڃZ�!�h���8Y��#�ڠ�ן��%�mq��kr=w��,�7����n�<�*��b�C">�6y�� yU��ԻR6��!=tܼiiR�~3�~rc�|C���>z�U6���U�i�����-���� �� R��݀�h��J2ېm����JFE@9�q��f���T;7JD�]gE�%��s�)����d;T��Ȩˡuhn���]�o���LK�e���I���u����!�N�Ɖ��0���]�ZZ(T�>�d/��`��j��G@g�#v�:o������U���`��N�v	/c~ ��g ��_��i�!Q�V�h��A3@� ��_)��n����N��K.���Jÿ��m�x�/�e�&��l�XXk���2׮�5O� ��M1p�����̗����ڛ�݋O$�K�F7�_X�Iوj��s�-�o�G��3_�f���ū;L�b=D;?�N�N�~�N��0q�. �P�����R�%����`��]�"��z�W��ZX챣5��)�+���W���^@�^F�+�x�!K���X��Ukof����ѷ�`m]�#S'1���C%�G����l9I&v�)�z{�oh-ٕ�+�����S?����Hj$� �d_g���P�v(��ӕ����B����PW��aJ�cۼM��q��I�k^ �x�xZP\"�h���Na
Y�@w7�G>�4�4k�ob,4M��$�;+�2$]�`��b9�WD���H�LAG:ɻ����m������@�PG�keL��O�!{�c�����_K������q�o˞��!���qb����~Z[{KCϘĈ�<+\
��2
��5�P$l�6|*dG�4���2�}
�'~!ޢ|z�۶*���8!W<+�N۴Q�g	m��<�WEP��'�5�ߌ��C� Ú�Ѵ� D�hNE��b���p��п%m����@$i�t�0�����]b.P��Ճ��!^��P7qp�#���n��%�Y��u��4Rj�s��s�f��Tq��s�Kr���@��ZH�E���x²ԨB'XF�L����o�li9G0�sW��f�6��_#��p޻�����Z,�q+L?i���������Q� �RK���ӻb��N�o^3�
�D�ĨB\���0[K�Ǟ~3�.~����)�/hrR�Ͷ"ј��.?�������k�֑*Yw�x�5;cޑ������	��P ^�s��$"
����D�����i�۬�.���y[��yТ�48E9�M��-7Ų�4���˷Zُ�aڻa�A��4�1�|-BٻNG;|C����2��%9��fѻݧ`���[8}Cf�5X�dezx߻�}n��)��aĦ�xH����3NOو�@����m�/=%2HL �I���`�O��	��k�A.KC"�u��D+?,2��DC����~T��t(k�_w����*z��x\GQ��&|��`2�-�dY�AJ^{�j lӋq!�G����-r
�j�Q�\i^��r"U1��:Q!�������,�2��tw�+pERSH~��S=�UMY/����1�w�D6�����p�:�I���>\��:+nm�3�^@ �b����6L<�0�����K��e�	/�|�tc���xێK!�.V�@ʍ4�kj�mē�L��='+6�+�tM����8C[��#/?ʒ���!~�1#>��1�,[�<웼Qx�Dy�Ĺ��t�@[��\��LS*s��i�+��a�!����A��w�*b��a�sx�b?�j�!���- <凑;|��@���U�c�#!�յ������Q�<���b��l1�b��ҥ��jX��n#��aA���a���PC,W�TW�l���཰��ƹ���������K��l���[E����P����k�����Z}�*Ƨ�<�t>���cA������rT 7W�-�-�T��l��sG,m��"�K�F�q��?��'�h�Qx�A!��f�;�b1�r#D��^5���U7h��(P��Jgہ��O��-?�WvSKIz6�.�<��6��Ǩ4�%�'4E�d{��n�JF/-�&-�G?��#Qy��A�C�dɯ�H��hP5`D�����]�TGZ�&�XP��V�Z�a�4���PM��x'�i�)�N<V}�(�XB'҂X��=K��r�O����b���LQ
����s�q3��z��n�3�&c��t�K�X���V5	���=��n�ǥX��au�l��pH��rtZ��C!���l�7�� �V<[���N1d�扤)��&toh}����z'�`h�UdtSH�Gz���ؕ����}�"��q��#	*�5Y��N>ݘSs2?.�܂�0,��J�hE�9u�GG���xj�*��x5@�gn4Ө��1Zb;G�'&��CE\Q�2NJ��Z���G�'��V~=��&o����{��`r�gG�ʬ�C4�.�+1c:�����ڣ8C�H�⦞(�̠�=��=K���y$]�}0��#�_5�*>���;3,پa�����-��<�[��0�)��p��� ��և&�����z6ػ�%*�����c&^O��X)[�Q4�]\Ri��}?���n�Mm�$UB�I��%���g�7��b�&%U�+��s�9�).�˼]��yMT���޿dg�v)�����cP5�>PX*��K���A���M+V};�"V&��W��X$!{�Mi�|�q�b��9l�I6��vpK2�{��qM��G�����@d�A���)nXpN����w_�a�^���<^�J��yb��%�l�I擌�e�xY�A~A�|���N�)�<%Կ�L ��
���.�a-ņ}H�`o���D }�,�3��Kӝ��5I�F�i�֑A�;�ە��Vxn4�Z{�Fi�O�Q�.���|B==�!&q-,J����d���!�kM�0߈3zP�<m�(�q�6#�/�{���j��^(\��iy�;���2���a�1�eR�!.<�|��յ��q�(qؒ����x�I
L#�Vl)��x��#$��X4��'�iB^8RG�},�卢}F¯luº+ju��e�ԋQ�9p8n�XI���W�"���nD,��~��#n�}����y 򧝤_��~�
�*Q�M���|��jc�����"�'=>1M%���X	*���LG��ʁ��I���jz�Ƀ��Z��}J�ˁ�$/=�ǢUGC��Q�B�� ��mļj2�7�:ݏ��=�g�7��/.��fpj�HNO���7]�a:1�Ȇ��N�4�*r(D�>v��|U.^��u��a1�����¹�)7����z�\���U���˧jDY�rH�z���e�M�S{³���.�С���e�)ք�1�1\�Q�I�:�&�r�j,Z�����u�O�5�e:�|ݿ�s^��$톋�k��3ʺIC;�� g����?�z�t�PTܘ�!�OJ������T}���+}����X���J��ES3�f+BS�moE4�]���㓚#� O޷�B��0���o��'�`!2m��՟�hI��l�\#�B�:���iB����teq<:�kʋ_��b%�j��{�Z�i��{��dE]�m�P2�^��k��_�K�<D�B�+����c:Z)]��|�ݮ��4�	���Â�M'Z���7�c�pz��m�idiY�%d�'�L
f*J�LX�.s[v,�:M�e���{v؞x���٣p_lz�]ۖӷ�v椳�`���
t��y/3J��!�5�0�m�'6�>�3�f������L������Һ�Y��!����:'o�6�+]�5��-�~�y�b����Syx����������i^ܹ�nc�ٙ�<d��>%B@7��:|�#xxM�!�
�Q��N�%ʈ_5�M��,�~���_��N�����0��q��/k�;:Y��Kw�w�kdprT`���љ}���d/l�\�\"���Q���h�n)�j��n�rI�K��C5 �����P&x��P	�u�竢�~�����/�!��d�Ur�Ek.H ԡ��-�'UO���v�� 	���L~"o�����wj)�1f�����9���۸���vO�{�^Lum�<��ؚ����s�p�L�5��U_���$'�>f��}	��H1�Z���##�\���� 
F�n� �A��� �A��
Ȇ1|�k�/pʆ�8@���2·h�붧 ���.�g��"U��za��¶�m6
�V����FEK�<ﶺ��D��Ouɼr/�L�3�X��x|�Xؼ!�+����W^4�/��k�>̈��fP����+8�p��i��W˔q #O-K%��#.{Oj�e���d���4gxj�q�N_`-:p\�
��ҷ[∮���]5I�ެ�Ѿq`�{5����2�d��Kd��0NGx��_ә0�5�'? �h�r����0�pm�{L�O��e'xĈ�?����f=D랽0�y��l� �uP'��fJ�r�rJc(�!�<Ft�A�r��e-�y�
{{�x�P����>2pEwT�ϫ(���Q`��ʲ�l���A����@�zM��m�qEad��߻�h�1�R��X�>��i]��iw���:fht�e��\��������nm�^*%�b���e��C�(rj4?� hoB+�jרh14F�t�Y�QQ4Q˗��i���-͓�g��-��)���v�a��[�Ot`BC/����P{C偷�Swﶨ��k���Zg�����SM�4Qϝ�v�o1w	���@�1M�i��n��k@���l&<U�ʣ�,r��>p�ez���ي�14�0�ì����p/�Y}�]F�2����|��g_���}����C �Y` ��ӘX����[L��ԍ��r�_���.�#mM*��6��QZ�ΑN�N�ǭp��%�z�G	���\v�,Wu
�7����	�h�'ϯKcvea��r�;!�3n��S�{�m`��e�'��v���*D��]!FAU�b��&��U�ݰo�:�����h�X�Q��`�׃J�q�����8�-�ᙽ�_�"�hxRdЭ�E���|7
��4yIyŤ��/Rɿ�R�����D��4�K9(�+U=�ᓴ�	2+N!)�ף�ܫ`*�e"�_��Q��&��!�h�����C�pt2m����9*N�A���T��[t���g�(L��d]�����ό��h|a�9�P���;`e����$F:��~D����&�l=Ԩ>�gf�I��5	��� (�[y�6+C�x�m��T��]�Uc��/��۾>6)��X7x���;��b�qF	��ن�^(�ϛ/U���r��C8hRN��|���Q}�_�~�:��S�:��K��i����kmr4g4"1 �{�� ����|i��3鐴�Dvf���U��k�
͆y:�w+�7���i~�b#��
��3��Z8A��}�=��A~��A���mw
M�'v��$z
������z}�:o�W����TY���t�k�ӕ���l��aE�&_�(^�|Nbbt�t��)$�7�ԏ��۲� �m��<�0� G�İ�̷�ӷO����T��z�����}Q~��62{(�E��R�v���t�ݐ�� ��Vn��Z&���&�Y��OX���,E����I��vA��K��:�x�/��Oz>Em�#��Lt������h'sEb��5^a���@B���c�DQ�m��	�W�>�ָ	�Q�Bx͞=��؄���G,�b���MT�̷(w����b��Z�7����Sܼ��vr$Ř��.ψ��"e��l�z�	u��IԺ P���hL�9���IB�UE�A^��6��E��p�� �ՖpJY�y(m� s�8G{KU���bY�S��`	�h���E�B��{Ê��������a�҉-*�%�0=���1�����ڒ��HU��)�\k�F�R]�8�ƣ�֨܍B��c��V���טD��zl�dю��%^b�|����Casj(C�����2��o��t�L*W���GQx�~��Z{YUSn�%�Z�kP�n�  m�t0��	TA"��8L��z(4�}����f1s?)���x�{�Өkq�����+/�QeD,�b�>OQ��dԫM������4��s��i,���KzI��m1^�HU%E�`5��]�L��9��(x��ZC����q�k܋���F���h���F�����Y:mR�\y��W��w2}�G�'��L��أU�hdv��^x�jQ1��J/��Y:���c|��F��=�r��3D���}Y�
�2�)���'�G&�q�8ڦ.��(
�͑]���.�H��0:8y�~T�>��4z7�D��(��h����Z���7�U���])!�:>L��ZIH�H~ab��^x���Ł�d���bvr���@w�O�w�u��H�i�w�.oxuI�V��&�&�=oZ$�C�?�7�Ič�G�օLߣqG�fN`lw��ؿ�?gE+�mo�퀏P6Ҥ�=���ؤ4�s
Xw�q�������UZ���Y�-���~���Kƕ5F�3?\�y�a��f.�
�I;X��Rl���%��I��ѮB��:�[��>{:V4�12��r�vf�T^a����H�W爸�F���q��(7�[+����)0�*󢯔���ê�S��_��+�`:�)���(K��$L���t��^�	�)�N��B6;b�.ȴP_1VM*Pp��tF�!]KO2�x� 0H؝!���?�<���ڋB�1���/	��%��&[�����`��M�l�Ԏ�[�١�ۦ<�˦�2��s;0��/�|��t'놡J�@�"�l`)�:�Hp��g���ж5�w` ���%��AAJ��m&
�ᧉ�$�e���E.��7!׀��^�H��6�Y|�5*�z1�e){��n��������<�%������!�V�p����>x��{���p���R�O+�b��{p�7�m���w0n�o��a�;�d茼i%�ظH��;%k6`�#CX�zВ1Y��@��v	Pڧ_�_g=v	bV"㾕���Ȭ���ʠ�!�S�+���1��J7��QMjA�����sc�q�७��.7`j�>p�R�r$':�AjW�\^������Gg��_����E���_A����.�RV�ɞXq�~>�SJ�4t���I�����J��U<ʙ��?�	J�QJEʮ	�VyOk,��àņ�4�x�)��t���t%0LE�y6�@&�;�x�}3�b���<Z��(�V�ˈ")i����r��g-�,�K%u���ա"9���t4� ��&��ʫ����nX����pM��: ]��pm}���@���>JGgl|���	M�ޥ8�z��>����۬�l�=��w�GiS��v��
�閛U�#�`�Kb]��xhJײ�s~KNzT�{���)x7���&.>A��\Բ8(�e`4ڑ�{�k�9\��n,[���{�O0�+X!�yӾ��^�l�ۗ�����A�9ޭ�����o�k� G(6u#Q���V�p%|�=�����WW���������khe�^.�sx F�fT?p��!���s+��ڽ3x����o�{�`���͹B�_�ܚb�=�c�����?��+w7��G����Ma��G�LM�MӴ�� )1/㦰��Y����	L��������~���j����ɔPY&���XA["�; =�;)E���i���e����0�L���)�!�������Y��PM?<�&�j*��!��j
B> [�z�	�Oc
 R�rG��a	jM��4R*R>m'h+�_��~����&s%mt�����O�@c���%&��HВr�����95�����0 ��8suCok?�09���d��m�0��b|ST������ټ��j��'P���W�E�fg��ұ^ D�	F��f3|�LxA\��S��
�w�� hF���0���Wa��q7b����%�k[���e�ʔ9c�멹E�w*�����qRˇ�Yk�S����Ϋ�(�u_�cx�g����V"���l�1Fox��h�L0*SWJg����ؕ��Hv���ﲏ�s�e�S
��WJ�����T���#�J�G��F#�L��9R��i���%GC|D*�u�.�&�H��MF���J��X�{gO/Qǻ�R6�`2�;m��#�����CN�
�+)��F�]G�� �$�f�	���c���b&�%�9^f�&�0�����Ҫ�Q��W�;$�Z�f[aڂ�f�b� @'�]�9&�P]FJ'PW�N="�}�ܯ��g��{�k=�p묵����1<������qN9�M�ّb}Җ2�:W����Qv�n����Q�&V�"r-�`��B��Z.�l��
@��+�I]�r�D�vp���-�ƕw�%͆9Ǵ���
���S^����^Ī����p�ȿ�Эʑ�-	F%�|m��|	,+e�<%F�L�ec�na�mC�r!$��b�nF�d���z�Cw[ZI�-|?�3F��K��Xa�A��}͑#���^�f�p��N5w=R��^�v9�q�"4�[�Z����$���ࡿ���#�_-����p�(:t4�t�n�)��I�v)oؙ�皈k�҄%��dE���P�r�RX=Zǣv�:*ѣf�`-a���F�7�#l4��L�a�[w#ES��G����	�1�0���n�Ǿ�[�;>�EG�J��}2�	�����)F)K�-&Ej*��+�n��!� ���K�S��v�|����)LdGg@�ݿ?vN	��6��F�E`ˊ
�db�M_�U��>�}@�뛏M#�p8m��������b7oU!������s�H	��w�A΍@�`&]Y/�p꠿�D:y��bl�Զ�8qS�
8�P�j1�Q��u4���~>�{���B���-�ي��#���q,on�H�r�ǹ�7��#�~��tCS�ƣ���#�>�������)z��ӂ�7�m���bZ/T������%˄!P&	��0ߦ �,�� �Rg�x�WE�*Pă?J\5:��\Ȭ�g�k��/�L�����@mYf��_+�מZ$�R���n϶� �~�mT8E�����L�P�vk׿��[��Ơ{en .<@��_�a+�b���a��}��:j�[�+|4� ڒ�m�ERf�P�����.��aX����h�;3<E�C|��[#z��pl�݈���I�d��QK�@��z��δ��XO�]"�J�Z�qu�+��D�����F��]����/�*~�xF;�
�`F�����s���}n���>���]���7q�I�L[(O����a��{Mj
�Q����/���9e��M24�H��y�᥍i'�R.��*r�9���;����l�����ڑ�������V�b:D4@y���(B����>Y�Ɠ]#�95+{K��!�Q�i$_�����7�ca<�+��P�a�c4������-���`�Q�*���b�:3T�q��l�Aq�_׀i���Ac�|��7��K�����`��K`�����f�l��N&���P�ۯK�ݑ6������ �������Z@~����q�0}3���z�h3��m�� ��l,�%�&	i�OQ�#�G֌�{	]�\M��E�ǩ�r!?jL��p֗��}M%����^P����4Wӛ�j� #!�Ғ�f�R�k�;K����cyv��ח��(]����P�_�U��$0f�L.� .��C,�%?����@����G<�K��vS^q+�eh��jV��R7����,-F�� �+�ak��h�$HK駰KIY&4�K¾/�^��>Z����%���ʺc��u��m�m��d(@L�������d��v��N�.�U�MT���S�}'9	�z_���3�ŀ��u��LK@�i�I�F��!�찃▵���2V��[�nw�2V������5���ڣk���'�R�D6|���K[��l#gu�tOK����!7�;V2��Knub�(_�چ���`��Rgfr#Ӹ��s�~�S���\�F�$�s0��=��؞���`)3� z���'�`�+��k���j��:�u��)��lH����Y�e�5dնQ�L0<eKŭ�|�2�CL������ue6X.����|�ej�{F���CUkB�b�,�t��m��� �}jg�>}
�����K�c�p籎�!-��h�nLW�N���D֡o���荰���%�}~߆a��k��F=��a��&.+�B���u�@��t�B�W��J����:}gn�n.��ˬA�	U��d�-�;X2v�h[0M���G�y��A:�����;�%�k��������ћ�#O�_ƞ暕a�qXtF���P|�n��A��9jv]�����AaU�ud$��-�q;`&���s�Th�Lĥg?�}�w8��̽L82�|��a�:;��X/��h�z�����Mf�����e�D='�~��ڵ��x�Ei��sF����,̄�����ORZ	-xiy�b���l+�af'�o��q8���Vh��Y.�]�|�11������#G��SA�%�T�;���k�,|P�8B��A ��Y����LQf�W�� �!�M��=��+��Qs6����q� ��hk���ƶ�H���CW�]���X�{��i��:��Y������w�� �x��;�1l�С�.��%j7��흻�:��?����k�x��)��u8D�1/n{
�0���Z��*��MOl��7ћ�iv��E�
;�R@�|F�H�j3t"�2��}�Ad�����`��f�L�������".��@���z��p�+�E��@��o��y4�O���@�l�&�Z-����� mŐX�K*p��OY.��� ��4A�Q�IkȀuc����p��R$f:22�1W���z���>�|t�YC�����!Mۍ>�ޮa��V]�48�7���f�������,����u��J��F{��n�Q�gx���j���1�=�\��p�U'yV�	�Z���,��w_؁X�4a�:�]a,�Fcm	03��G����̕�~� ��8�޼�Gd�X�nx��00��3��d�23.��(�L���{o�Vk��M���a�F���dʯ��2���%�4���OZc+J+��Z�=u{k3�B.j�Ӛ����U��l����3��A���Dg=�!�}��8!�1B�F��ś�
6�����=CQ�I�s�A
A�1Խk��v�h�ǒ&�"��؈w�
�* ����s�\���_����ʱQ��@��VT��ʕQ�z��R/�0�!�xu��R1�����(IN�K�M��+&�&��?c#AQ�W�S3��]-F䙀�?���Jp�l`��̌�����O�拖���%4�h�0x�"��ٖ�P+'u��*.�I���K��|n�p;�����Rh���H�<0[%����&��`V���U>�J�O������+<�:?��� �'�C`�Gb��v^�,-�p������c;�z@����VI�Jw�D�SQ�p+|�^P�C����o����X��r�_�Mt �>x���jIBK��҆�ҡ���3�2�F��=���o4���+i(kX�6h���-��j#S]G]���U�ת�H8,��4;3���uJ�����������7����B+F�_vX'ԍ���-�~l��~�X��6wm��$d��j��N�2I�І��w�H�5P�u�d;9j�bhA���jIa	 �3.	������$�������o�|�=�R |D�c����ԈŖX��-~j��a��)�_���չ9%]��9/���Y�+V =��^[�H]���3� ,���8ꇮv:�h��%#��f�#��n]���>|:vC�5b�\3�ȳظ�e���.�B鴐iT��zU&줘�O��Q�D�E���["s�T�N��S܂�4�,�"ۙ(7)�f�m�7����� ���h�Q�����Ψ���OVQhXZA��}�j�
��`|�$#ž;�m�).�ޙ�.9�zw̢e�c0k����0�ŇJ��pI>�դ�!�!����9�5Qz+����''���+m�^u%��D��A��~g����5w���H�X��/�6f*��c��ܱ����q���A��?�w0��
Y�3s�Z�(�ξ�-�|���x�q^0���G6 Bt�C�~&Z8�}��Rx�s�h���[��KJ���v�2�5Ӱ
qɛ�fM]4*���rvs�X&��M���C-~;�|��?��\�5����,�'�0�(N�k�j[8�:h ݼo�)
�(��<�->�.G��;���Q�)�`U�����B��;ZBo��f�!��B��)
P(�{ALI�㊱�plE����[J顔S�aO>k�Q�3'�N2��O5�Rդϲư�/J-g�<X>��f�G2����������UY�����6^�t��{�=�>DO�]\�����1��fZ���;��5��K��y���pwKn8��:)Es�)�)lZ�������(��8�sN�l;O�!4#��s%F]�H��mLD�'ׁ����f��`�B��nk#�!�Z��U�E"���t�V{�y����9
H���QB3vX�|��6����p��3���L�)���n�E>	p�R#4����G[gb�F�p"�GCZ��kx�U�$
6�!w�_�H���6{���x�='���Vj�nV�̯�(8�J����1N<ܗu�h@;�d}��ë�~[��֐�!ro��t9����ڒv�GM�6����99���ܐ�;���d
ꣴ�۟Kl�X�h��I8��Be��`��K��I@j�|���}
��Y��T0N�N�?��ܝ�6�~V.Y���u[S�)���Z�&/�r��d�&gך8�wf� "�)9���_���ݣj����疞��m\o�u�r=/�2��zr��/���<ԩ^sőev%��,wz@e�DY��L[����eb���&�{B,��Qd!��"�E��Ԯ�k������
p�G����^�9�m�Ln�4���iiX�h���Y9ڧm��1:<��|�"/��9H�]1�A�Djz�fc�$Y�UJqQ��S����M��;��5���Nm�8�d�+eDP�UCO��K&-��d)�A}!m��`�[�WrVg����hOGm?��wϊV�v�Ę��|���ѤQl�h3JS����ū,�'tȪ��n�R�%��3y�C��F	�uܓ[ 1�>eҀ���P|�����g>��]
�/�2�5��c���o��{F���l��������F[�� ��bSbf�
N
�Rʥ
�����aȡI�'jkW��qLC�+EA./�|IۃU)%~��`��_�|p�n���*��������	��V%@ �P�8�Y��+��>�w�&���!�5�Ε��ʷ��$���5?�(A�;�K�9k���:��9���):}r�Pƿwl�i�:�6�h� �Vd�8C,U�\�Ή&V%xQ�d:D眳�˘��81��{!Q�Y@Si����؇���bH�5�BxFf���:!�_Eж��ϒ��%G[z��$R?;�T5*ܚA�K9t@�	b�q$ce������q�g��*"�����<��h���<m��O�_pP��0��ؼ�h0� s5�B��og���S���,1�8fт�X٥EC��	��P��st:0�d��$w��TP��.Ae�PG�#5��O8�THK7ۑ:*?" usG[+<���I�﯒҅�=�t1}�HyW#Ē�Нo��[v���k���r��k��/��,,����2��N�*�l0Z�]�&�<�������"�%��lCJo[����찁Mz�Ѻ���t[�z�Qs�n�D�
D,�,=�Q�mS( y�u@у�W#}��T��~)# +`�˒q���`�`�/QI�SV�@m5g8��}^� �U�����F�L4�*k�a����.��z��\�U=��&�6���$�^o>�|�����w��T���N�����K�a�!��<�؎m��2S�c����+%ˈ�9Kqͮ������n��`�ZT�$��p)Xʝ�d��o3�UHoX���p�Y.�/�kՌ���^�Ezy�6�ۊ��^�Su��iX ��`���9��כg��맨�`�d�'.ƷY.\��]4"[}1�#����R�ݒ:�� '�`�#"�U�8֭�tQ���g���v`���|w�QNw�����>�o"H3u���u�0"����g���^[˱mC�	��*,F��mhdL1�l�ĺ��"�˛��m�-J0)W�H���
�!
�,R�Ky������!I����3κ�.:�åB�L���g(^��v�u��E��/�����[G�𜍹����HX*��~Bfu�b����d2W�/)�xrW�|�4�.ɓ� 	ͧ��&I���9�1�dD���,��X�Z�,6r^)�_�\"�I$�4��X�����q��c��y����ƾP��E4F�%��v�2�HZR`��n��$���"�߬�߮�=�;I��{=$��Su
�ez8j�6jS�FƵ!s�k-�zKp���~l�~�Е���{�:��� RZW��Zk�3/����j*A��`���_Y����{�ʩ��A���\���¯'��<>x��1��u����ءb�Ve&���G讹��r��jo���t���
;�EB������c����du2���Ғ�:ۀX���!�g���m.����q��{�(I�&����������
E��g�>���Ѩ���Ejr��Oe���~.��U��h���%D��[	�?
3����͑����(���L%k�����P�7�yV������ MjG�,��O��6��ڟI�����b? l"���(�ݜ�C�%�V�R����
�L�9,^�	)e帉�5UGܯ�X� ,/�B�No���#����qϻ�]I!+s�\�TGʠ������f��VW�%�,<ݢ ���,}(w�(�I����#�>�+SO��l����|X5S3��{�K�l�J�L����F�<�h&�q�ծ?���h$v�]����ҡ7�^+�)��l����8��<TC@dP��dDԟP�ѐ�q�������`�O�(�`�/�k�r�%JvV�*�gvLt�>��4�gi�x�rgdk���;�W�����2��n�ps�h��j���wv��>�i����zn��,���~�[����/��E���FM�Ĵ���"Y'`�Ӥ���KGF�� 9y�Ȋ�{�^G.��`S�y��&��`���6�2��s��O���SI�-��{Xf�>y����f�������َY?l=i�����_ciTGQ�[�`�Ix_��99]1ϡkK�7 I� �b���z�tۛ,ɺ�<�-��~}Nލ,`Q�`���gE�:���V�? S[��Bz&�kj��^�8��d]�^R,����EY!v���͇1NCن���nS*�ǜ��\x���N+�5��ىͺ3x6o5zW+��=�,f�*Sڡf�L��:�YO�e�����5���&[5Ǉ�|הn}����_��?{���@hL�=�in�&+�4+��������0ac'��#�W�`��{b��-cIl����β8�ߨ�:%��y��^n㙧��=�!�:_��250'G�4�~��{�2�*��o���_��V�x|�1E�
�Vq�a3=�q]��}�hs��u�?���~.ﮑj��� /:D!ʑ|�A����E���v��{�O���D��A��KΓ�!��f���V�z��'�<�L�v�����\f��_�k��I��?���۾=������O�,�"Ls���:	�Nl�Ȑ�a�����E��[|ػDi{P~細���?�������tl4	[0V7WLN�Q�2xk�ZO5�v���Ӑ�3�8;�'��ׄx�s9�c�S�7���d~`��<��i���>���Mtz)>��D�>�֢M���X;�%YL�õ��
�
�y.AR�蛻���n�U4
���,cГ!1r����Y<��Hؠ/���&�^�*T��(9Ť���i٦]�3��.�b��v�p��A�
<�t^j�[�!��QU�r�uq˔-Z���5�>��� 2�I���f4��Q�޹��w���Ȗ�(�ED+�
!�'=���C(˻��B^�OhL�*n:���dE$��<������ �R��1_#��Ǹ�Yw�0$䦱�J��l���kK�Z�|V��h|����B[}�$��Ep{W|���EA
�$Ƙ15)(޵�����b�? ��]��K�mwM��/�����eO��MX�Y��A=��~u�o%�:P`8�%b�'�&�./�0�i6S�z�
+�Ҽ��tO��-K��O���x`?�0�u2�wT-�����䭆�}P� nT��K[8�
�@ȱ&�V;�q����)��>�m�P3�&�b����1�C�pa��z#/h�4���X����#W��e�ڙ9oq�쌷��G��/��[B��M.�o���n��3���ƐrO��Z�8E�x�.�����|�q�����gc�~f��������z�u�Z��_*�Z]���lAM���93�^���V{&��Ob�'t�0f�WY��F�	T��otc�:��E#�&w鯣��s�4Ty�a�*�����1/���{�ukV�X����f�޴&��(�W���_�	�����d�kZ����ח��ߌ �(���w�沵�x���"�p���K��\�(��;(u��3�+�P+����N�s.�Ɗ��g�+�`̏��}{˃3�m;��ୖR��֨D�3&��$K�c;`;��̷!ٰ�L<�oB�O�=y}�:���K�&b[���;�0�S܅w}ש�/$��/DL�!6�'L�7^�?�(M����_�����F�4����횚e�=�_"W>����,�'�9���C�~J-\����)~��ߵ~�b\�v˅����uYL�a_-��Fߜ����%�����솿���Sx�ކ��f�Fȗ<��R�1e`���"���:��3�@�ӹ�����n�͚[��R*@7;���T������j��A���r�h-�2F��ӯe�M�X���b߃I�f��9R?i�U�~!��QĔr��=��d��y*��=f&E� ӬKu6|'O"��g,\��ww>��q|o�2��n�zʃ�M^��%�x�;2K�w\�� T�R�շ弚�G\������^8']��2��a2��>����y\�i|������C�Ë��Ĉ�U2W�Κ-�*YHI�Y �(�h�آq�Z��qw�#��{�ܻ��ṡ��ԋv��R���5��������]@�� N�6.C۷).t��� 9Fl�ȫ=�>v�� wi]�4��	2��U�̈́h�J�0&�f>�L\�����w.x)¥���k� 	}.�1��[��!7�_�I0S�u<�k�a�\O��ȚYY���RQ��ʱ�v����Z�/���.���,�g�Չߩ����E����ߩ��|����r0w�Ӡ��%���}�<����t	��כ1T]U���S)��-�� p�òd�F*0�b"c5�ߞ�$��
�%$���a�Z̰�l���\0Xzp�.U&���w��
c�h���Db��漏��j��#n�ЬI�*��-��[��¯�9�H��Oq�o�W� B��_<�ʵ�����FU�I,--"�x�/-�{�ۜxn
����3M�:��ۧ.^���zE�x6����l��mj�&�U����$)(ܫ��9B�ъ��ܲ5�� �J��tW�SY2.5I���7@A�͟;:m�w[�돰�,��_�b�1�8~v]��T^u�p�_���-�t�{�I�?�;ߒ�LmA�hI%k�	U�E�09q�1˄e�D�5�ŕ������A�pi�fi���]���ш?w�3��#og�NmsE�a
m���S�T�fl1�0�J����~�M�L5���j���!5�3Z̾�L~�v*�!	����Ȃ{�9��͊ � MĪ�o'1�%^��$����CW����\,�V� �KEX��r {o�� ������`*1��:�3͇{R��o@�0����Q�7��.'���r�bd�?��C��9Cw[��]Mz�gȎ)��Y�PE�6���_��Ɯ]�~K�O��Z�c��E�}�0ه�o)tJ�}�j%H/�
	#D��s��T�d�����Or�j���C(�]*`��,)����J��| ɔG����u�ٱ�d�7f���1�����
�[ �����׭[@��/��oK�5Qrb�AXr�p�y�dv\m���ҧ��Ti�����~Z	~*�7���(>�W����hz�}B�	�4�t݉��\mSZ�R��XF��w���S��w�����[ L��\��d
@s����K�d!�+�����{V�/��f�ޒU�21Y/��+��q��cq��E�8(@ �'�$���������R�L&�oR�0�|_��5��ӪY� +��1=}D{~Os?niՔ�j?̥Y�]�Q&�RE[fU�۪���t�艗z���*�2l<�A}E�o�]��53A�Q���j����eW{Y��G��n�"pB�3� TG]A�����~(��Cİ!�"\=������6����س�(������[�Ȩ�5�x���F���hPGuH�d��:ɟ����%6���RDG������O��K�.�GPNN�l����׷k�>�����O*Ѝ)��P$��ss��*$
t`�2d�@�wi�#^e"�UC��+�0�jc����T�h'���Axf�)Dt!��{�eYc-�o��A�&�[Ȣ<'yS	�������n�#!����&�í�ˬ�-����	�]���IM���z��޻���$��_lO)��涵����6����\9`?4���/)+�_�.���~������~<�Acڷ�?����܇~f��4[�߇M���&�o�����-�7��E���4Ò-��S o1B1F����e�R4�q�N�"�Žxq0�d'!nD)l�|ρ�8.g�m���H9j%�Y����#KZ7?��.�A"J?b{#N��r���	HTa(
_~,�s��;����QI�n�?֦�+���P��r&SzJ�vѱ�v���ˆ;�]gy6��Pdg����8Wɿ9=W[��C��-�1a����f�8U��]��(hN)��8���u���ԟ{-��7�o�(���>�mvj
��X�Z��$�cx��z��m���n�0&��6�݃�R�����Օ,�ے��Nl��6�j��g�*�W���m�C�c�d�drD���Cڧ���i����h���^Y@1\K:��d�j'G��A�"�͎zO���S�E멪�\׿������Cw�&��4�Zܕ[6i)�1	���dHu�U�� B�aZx�<�=���L�b���Z ����&4����SU�=m}�d',�A�+:tܠi	��v$"��ե8K�p66�j��{)�]K�D��M�DN~,����׸
D��wN
<���}�H��њ@���<;^�_�m�Bh#��v�R��):M@u��Zp�g��|�^�Fw�P�`=���2I�����ܗ����<E����P��#�	��3ӌL�+/{ 3^�S?o�+f*n�Lh�XkO�Q4��� p̀�{A�I�2z�� �x�~#m��w�<�J
����H�k
Ӿ��B�	bf�7H�>qm��B"pE$5��^zI�2��-���{.`�ݶ*C-12���; ��g��)I��y:��	>}�- 7ʎ��W8�D�����6$��B��N&]<�U���:om13a�2��;BW�_=%�A�����n�t%Gn�vTF�`�7����~���8)�r��W I�n�����gH�"Z�2� Y��ۧ�3�~���.���ݭ��Ѹ�rh˚��E�r#��C�w�Q�4`���V�"�Ϥ�en�Қ�(��a4���p�g[9[ŪfH��G�%&e������@���ɒx��HreΗ��&������돏�4y��.P��2�7ײ7lI�qWw��FnUu7Mj�繻������;��o��������䂘U)w#����`��/^��T�T=��9�8��B��`@�{zg[��!rw)u�3�m���'�<��/ߟ1����8��A�e�D���'R�aK�.��&ȓg���d�c������=:h����P�>:};Z<����3��nu�q�S�e�f��������w��g�H�-:N�8����X[|�!�cl|�y∱.eX5�F�i0����btQ{P׃y����tQ:�Y�	�N��{u�W�:�b����>S�C��D��'�L�5x�q�Y�W�w,!����������>e9�Q������׹�]�*ݛI���l��:�V^@����V٧����)���о����2��3��Ƨ��R$مi}����~�����Q���"5�x���4=b������k,��@;�O����i&���n������Їb�(c�\ơ�o���-�4x�o@�Z��d���aok��&dI���0>Zs5�~E��"�~3�0"N"~T�@%->����,{~P�n��H�Q�����/���^.޴u������&�R��LN�U���^{����:�vV�py
xכ�
k��w���	X�^S������� � �Ѐ�G}�A�md8"樠n�.��-�>�Ε���t�fȳe �:�uE���N����(������wg�Zym��7S������jx�b�W�����)r�RxU�Y_��LC�4ڭѲ��.��}p*�є�y��AJ�5D��^ӺZ��KPa��!����B�H�o+KԤ���Y�K�[�Z�mK���8����W���(��L��0?h��Ʌ���������4Շ�E%�2\7��*�M��&n<[c�jg���}H�;��㳷L>�>dR�֥����	��hi4k�N]Ka�\1�!9I�ur��u��m��H}K�n��F��X�	\�e=�[����J҉�?CD~G�oC�C\�m�W��9ϫ��}P�h���̆��"���"d�9���J#��'��;�(��S����^J�Y��!�O�^g>IX��gd�WSC�½�7�Q�<��*��P�F�P)�~� #��$#����vq~-ծ��%��i7vv��ܜ��'��!�e���j����u�a �/��9R&i�@�ٓjp��?��p0ԅN2)y����L�(-��鸫Q@uq3��7 �rA��V����,C�X����K$���$���)�߸��Ri����0��$z�(^��h��RHWՅU
���󍦶��h�R���.�}@Ʒ��1�[�U�M�$�ty^����8#���,�����E�@s
��O��[s�����%2��{燎�YSҫ�o��%K~�=��ߙ�'�h��a��݊Y]�r�T�ӝ���E,�:��O���a�M�R�9h��k4�Mowʴ�jTc6�?��Bf�Z�/�w���.�wd�a�E��ʸn����D��(ȸ�FKx�ܻ��.���P���1��7�VRf�T�1tC��qY��t�{��`��#�*l=����~����}u/9�>�e�'��#Ѷ�ar�ηG$��?���)�P���ku�^b'��l�����E$��ܫ���?�rI�|1���As�э�q����d���X��ѥzp�ӽ`��,Egtզ.�]��+������6�x� c�F̣�$Vt�es��m�4и�4܈>�:Q�;8��yf@ی��愚"Q�z�������n�C��݃��H��j�{����ۗt�������V�^� ��R"$*�A�&(�CF}4�_�H���f�C��3�ţ-jL�	��ՠ�ď����G���{ �0INO3�y�^NJu�9���][?�o�H���G\eK=
�1�0 ����:��t��b�j��~�)I�=Z��r�=!�-���x�Z��k�\L5���\�ܺv��7����v�^���t~�aؕ��n}�f/�� ��t����qx�=��!G�[�f�y�cW�lEb���G�X8�r��G��k���K�wg�ֿ6�O敭�zd�� _�q��7�T"�Sx�b��Pb�Yq��9�G���ޢ�  ;��v;��
������M"&*���J��)vH���B���J������S\ ����&��Pm�M�W�����w���|�4L>�KP���6 b[b�����b�Ҽ�tȏ/RҴʮ�2
�ù0��Ӟ�A&�Ũ���/.�� /�zQ :�m���$d_M
PfX]@2��K��k�T�7��R'�D�qF'�`�}�l<�5++ÿg�!���� ׻֪n�[����)��^qK!��Y�)rVjwK,8h!����F����-��X��B���^C�̃M�L��HG75��~�,�غ
|�����H�+p�R�c΅/�v�!j��k����5/�崶�D�_�l̟P�+���w[^�de�T�G�{o`���3�~'m���𺸈.��fΨ�ۘ�#���;AyK�D~��u�,��E�S�2y�k� MR�K{Ѯ����]��'䟍v���&���|"x�z�р���h�ft4����%�t�b�^�?bn�Mb����db�eM��
��<9�T���%�+W�xo��10�/]����'��ns��1��ꗶsn|*⯣*�m�B���c�N��GcC+^�������?�ɐ��g�Y�ʱ����iR�!r�{VhZ9�`��������ѵK"(��?1����-�E��R �f�o��j���ӘO�'f��m�gK�kZCϊ�V�]l�3 �h��ջo1ڝAl�I5���0XN�NYn&M�:a^�`[P�r���0ʐ=�C&���q�I-М+�S]Hv�y'X������H���Gӝ9��u��Ps�+�~�+�����?�G�/9V�	��kI��l��B�OĸhjI[�/{&�������O�˷��ρi���iIU0z��`�g���i�[5Um���!�+V#$����eV����m���kV�#>�ױ3�a��I����Cc�"�H�P.���O'�Fg��H��v[�,�>���������6��0�M����`��g��/��2^k�g����7��-z�6h�^�I1���0��@74�01��o-�3��o+P
��'W��Ҭj�&*�ͱѸ[ ؆� z̷��f�g5��2��i��v:(ez|V���d�����M��d��j�uCy���@w�z+����d���kw1�����q��8��AI��͜%�ĭ[�������KؑL��'k/:T@V2����GF	�3
�ˣt�'��)������f;B�f��ޞf\�9�׾a������l՟Z��wk5IG����oANCk��'�Y��"cɵ�ocʶ���u8�g8V۽+')�v�O�(d7+ރ�qxF��,f���T^aT��h�pR-KH������`��jd�-�1���D#��\,�qTز�!QK9P.#���S~w.M�T:6>�O��Ҷ�;^�(�ӗd9��n=���a���/�!�i�x=�*s����%�I?��|����mJ�-��M�>��
? ,��[�g�ᯔ��p"�ݚ�nђ�?�"���	�� �B�8sc���%�����0�����	4�ɇ����;�oR��
f�tȿj�L��ٚ���Ē����z^C��d.��w/w :17��j� �d"!��Y�wo�l2G5�r�ɇ$�x1�R��C���\�������4RBD��`�'%ԑӄ�_��b�g���<�����0�(�t�m�@�B�B�����@+��R����e:��9ɬ�����>���]�5�
�1C>.NO?.�"XFk[�]�ϕ��o�����q,O�Ы���7)Oz�1ɬ�G9j֚�٦�4_����O�D��b�D�l��pJ��h���ziodQ��Rw�J��K�5�S��3R��I4#
_��D�����K�3�)���|ɠi��N��K������j�n;��ʊ����	��-,�1@˔�z���$E/�R���f��!� ܴ��;{m�	jLA���lE�*4�*�4�2d 7"������4��,�1���F:�[K��-�q��q%���֎�����ou��!2h�X�a�@6X�DE��H+�j;����'	P�|�����ʩס���;L��fD&���?k������Qy��U� Ca�}(%yU7ؾ��kl ��� g�<�u���9�h\
�;��K�π���.��ط?w��V[-$���?֑�7Ù_�^�����+$��,2�lʻ��#�F���(��������a��U��To'�[���5���F�����B�W=�C��f�C��?����CpG�Z����N>D�Mc��M�҄�T��2�H�ч���a��P�7�L�Y/��G��'G4��\uk�5�!Pn�Uf��0۟)ĭ�Qv�ؐ�lx^��ڢ�W$2�	��n�/ȑ�԰�����Gf�:	�n�!�4�;1�rp��E���:'p���.��F�qYi1A�|�8-�D�k_��G��F��j�g.x�o+���d7?�R���w�y7�sd	�Q�P"~��j^|�����&K�C�7��V^��2Dv�2 /j�n�U=�Y/����yV�)�uo0��{3E��ai�N#�i5��*�lEit,�Lʔ���<C�&)���5c�ۖ�I�����sZ˧�pJ�
b\h�����%X�����˘rѫg�D�a�E,�}�H��"��+�d[b�5(�@�~�Z���2�5k��%aaMI�{���C��g���K]����Bg=,�8}�@�n��^o�G��m�84���g�_��䫴T��#8n)ff���.��I`���[:��@�%}flʖ��hN~�{P?ue'�o�E��2������l���㇠d�:�����o���������ѰP�ۼc卙�\�y�B	�,����g��:�J�c5�Zs6��%�Z\Q48tn�seiT�e0�׍\���t"�59���Q�V0k/{`�Ql&�%�pfG`������� '�H\n�j��Y�[���>Z��R���J$�r5{hά�N����|�� Kw��2��ƳĜ�*:d~�c��?p�s
YA��;�J%��\�\���Tb���]|4i���I�5��Fb忚�feӠ/�Au�\��p�K2k˝��qj.�*�O��-L@I�<�I�Tqw;4?T��������:�h6�Dޅ�;9�D�Q�>���c� �M�Ak�Twu�6a2^b��UM3P��d���赁��*�o}�l�&��θ �ea���Ǒ��LOp_������=�Е_e�I�FI�Sr��<�y%��o+*;4��D�8{�j��}?�`	F<̧t��q����0�G���d>͕����Z����n@}��u��.6��
�+��8{+3������J7��@�����
0c/�a�����l3�T5�DEX���tz���z�85)�x���pW��I�*��ɻ�0�廙��|C� ����Jvg�����nj�i�eA�Z#�S�
��DQCJ���bc���+�=��B@�躇�.�F��^̸o���Б?���Ca�,`���iz�@k0�����f�0����l����wiC��>�쿓s�'����?�SS��j�@� �"�J�%Q��I��ã=�2Óm�L�K
�&l�wc�ˡ_aL��Zԃj�.p��f[�l��dm<�z4�C�Û��,9W��q�i��/[k�#�o1����������Al�s
��j}�S���F�Gൽ�oȞ����h�m��(r���+7��<(/NՉ��)V~i
�=���\������/C<mg�̻	&#=�FB�,p=Joc93�ӯW�yAG�h�/��\$i����Gr���/�I�L~O�b�.��mTi��;���V�\K��FA9�&:8��楬���q�F�u�c[V3�*7�%L�hM��*� +5�j0��<O�F���=iX��;��+�+]�A9-'���|yk�>!�:��Φv�ԝ�q���F2����cT���'߼��J�t��fY
�������d���#�\��?�/d���z�k��i�n������ s1�_�'���(14R�����Ц�nk���>s
A	�MH*Roc:�P�6l6%?y��Rh(qA'�0����7U�pb�7-N��e`��7)�&dkdc�*���8}�k��J�G�Ī�]:*+�M�$m�;�ĦpK��8a�ޱ;�6���=phf�
�S�=H��5:���:�%l~�� 9,kZ杀���TN<��Dm��:� *��u������Z��Z{Mq<��e;�<Ȋ�/RV����X����{����A�����ǭsֺѪ�d_5����=��oY�=ag�*�}_�6����4@ �'_
m
����>��G ^��$�#|q���;;�f�_�����ħ!X�.sa�f�7�0���ȍ��W�D�xna���Ջ*y�ᏄƵ���`�<�m��'� .���Z�S
a6{�ct��1�S7��C���g:�_ϫ�H�M�W
��,b�\�>a�2q@��c�]�_hSH��� !z�Ԃ��Ia#��L��/jl�!��G�yrmu�I����ix9������<2w���}{�^����=���C�z�./�gO�^qm�c��G]�o����P�AS���í���81�\��p���E(�Y�>�,��Pd/S>`�P�S<��Ic��H}���@RQ��i�"[��ax�=	[���;:+��ʜs`�*e!��o�+�x0�x��e�w��o'�NH)�e�}������:�D$�x�������g5���KX.�Pxy�Kf�O;�O~��!�CvĜX��M�6C��!%\N�"#�KrS=X��z�Ee��}\O1�a���o��}���R���ujǧ�`(�N;+d��)T�#�a!dbQ��dv��&Q'Z
����)*\
L��l��
�%��j�;���oۜ�+�`�`��8
b'��?�������ޝ�gކ*�/�;����s���]}�By��ɞHQ�x��[f
��e�,k$ gP���B����܀�OKĤLһtIn�Dhpl�P��Z�oCjb��
�(������+��K,a�Z	�dv��s��;����7n����;l���C���qi-���2��S�~E� �b����/9K��	2+])V[�A�	pl�����H%j�x�Р�XD���"�i!D1��1�"�xT_p���ֲ?'�s���"}�(#m��?Z.�z��7�%�n5�c֞l�!v�x��s�����w-s^%�sor��#��l�}�}ew�� ���֞�[���ZO��N�F��f�9� Li;�'P'���<���!�]�g{���p��^����U�o���*R�V`�_���&�ƅ;W��زw��ts7��Y���C�x���y��o����W����)o�w��g$�`P���k�	�)yG�������ܬ-%-b�?&�m,��D1�^�V7���	q�gYcxi�@�uE	ѱ`�Q����)!$:PfM+A��F��sD�=��3������N_okVI�{D|b5 =&�/�^d<����c��6��~�0��~���B��@�A��������9�|䴣1��9�x�:CR8H����\-X�Y: 0�,��6�ڒ��A����=���^8���t�����SN�ǿ��"��$	�*�5�2Eí�pUv�Yx�'��Q�9wzb����.��s5�����ΌS���3N�N�Z��� D)�-4���,��/54ƞE��N÷(�=]o��_A���a�^���*�.1~ɨxIhHV{�ڬ�s����<*F��:$�%s�i-�x�v���cL��{��w[���jHB�zF���nQa.~�i�����i ѓiMp;Тٵ��+;J�O�mp1�����D4$]�6����K�}˹�7�珿oq��[��X�r�\i�۴
�A��<Y��fil;��a��������+^�ԁ8�$W.�7CF�|i�z����}���n>B���6�65Ǿ�Y���7��f�6#�ۮR��0�V�T�u�Xz)��^^N��Ȱ+�3[=O��F��i���]i־26Ҵq�:m�L�&C�E��I�������>EG��$�3�D�^Y�D5ֳs����x ���.9���	4��9�Qt�މ|�(u#ND���l�	�~t�����Eh$δȡ`k/�j�m,v҃wkrވ{ˤ�����5�#�N�dU+w\"�����aO�^�����b"��6�D���cs����fڛ��3<�v�/��/x���h�3#���٫�����I��|�J<��~����d��v>�N!�x4f������<Q��O������3����}������{5s�ٙRi�`��}�`�r|W?R�>�̑i��)�TZٞ��
m&�@b��Es0|�e;|����&u�U�/��3�;�h��WS鄋�Sb}��'���پ�t�����!<����`&���hC�]a�G��	|T�K2ڏ�u�]��s�����<N�
2"P�5��KY�s)#�� \�=W�<��/�eE����,	/C��ûbĐ+����H�*��2����a�Pח��D,��Tg���C�3z���]�M�$WkY>��8=�<���������6"h�K�P�#���h�=_	�c=A�v<�o�?�Rˣ�r�\J١S�C�2N�|�9l\�)��X�������5Vd +�@�F��ԁ�m�Z�p/-��&��$L����j ��Ӹn`C��	Ե���8@��`��Ui�����L��e��	�@�R�����&�m5��?h 3-+��)v���J�]<�4���T�����:s=�t��<��iȠ|�ƅ���0��L&���T���Fp�������4D3ؽ�3�<9a�~"1���w��Rv0�f͟�A�2k���f�O��\�f�K�1�*��y�ԉe��ڃ��2�����܇x���τ��;��>�-���$�����+�/���_��'�ZΓ�����V�N��2U�<�X�u�U���2�)E��eR~��JR�c<��lf�ݯs���g����3��m�{o��<Z��K�/X�)+�38&:W�ڍCɬ�iq❷ѮNfz��jJ������rYG�c����D�Sz��<f^5�J����;F���L�-ĥ��B���� �⯎��˥�R�NZ��Y�oN��d<#٧�B6�אAa����[�\M��2�o��si�������"0�/ű�g��k]Oj���@�?�Er��CT�,��u]\Y�y ��]�=Qp@��ݼE��r9}��;��F@"S&�����a^��W�eyK�R
(�4���F�ϵ�I��uf5�hJ�3��_Gq�N��a՛tc>��]ϵҸkj~N;��j�-FiG��:����q-�m�a��F�;Т|�����NS֢[�5����Mw�騻19Ȩ��֢WY�r�O���:oTlP!3@~�ͱ�4��F g50�/�FY��Cd�S��(MX��>F"�[k;>̓Jt�t�Yc{Y\>C��]��e���(�����|�q����&�Y�0<|܅� �D�w��sT4	�~6���X|�p�������S'�P,�c�������s7$��d=J�x��C{���m��	��ƹ�JLHY �9Y�A(��oI̿��~�۸q��Q��J楢b^Op�ݥ@G�^^e��9����g����Ќ����q�0����$�c�"iT2$!�Fg,ɓv��kr$�\a��A���m�v�v��V����l%�n*Z���n3���5P�vΊ�Z��}"�1�ނ��T5���I��}>�����w���x�%�{��9-���O�SM"��һ�co��c`$�	�}q�M����3���~ڧi��+��������p�.Y�鿯h�!��1�1
|��x��c~ꫀ4F�^{U�`S���������6߷y��z�:�.s<�踇\k�W�N�V$��x%8��@���_�%acs9!oMs<���1�� �xV!s�oF�yߗ�z�C���,��dEnl9���f��n��vT:�Y����p~�+�K'������98�T�s����H����G���9���,I�1U���W��Bܗ+��g�WS�_}ӄ�#��#�k�z_���#>K	�գ���Z�	t�1JR���L�_fj>�[�cP+�뤥F��1z�c�Ճ2�i<�!("vQV G}8�:�a��@t^���լwCŞZ$G��N'��/ջi͵�O�]�N��6���>��.���p�>��!F�t�ȣ(�_a��U&�e��t0B�n���V��e�x��.�Q�[q��-��8�#�Gj)�|����׵��{H��:\��V��cz_�oB��݆�\����ča�0OA��>�@.:UGtf¶��|R6�'�ޜnKlmm�5M!bnH;�������gso�?v��m�M�h�x��Ш����6�<���n�?^e���L�+����C����[�d�'�6AGN,V��RUL�*���>L2�F�^U]�JPD�C��%5��Ħ��u,��u���%_��t#gVHJ���F.��p���J�����Vt�v|�r�Q�?IgΟeD�umS$����M/�E�A�ⷋIY�24DQ��$sl�h�j���,�V09��*����nDE�!xĹ�{Oz�$���E��#F�h�`�� P!ؘ����Ս�&�Ȟ%�j�m����㦕,ar�P��'�"��8q��p)k�=܋<VU��KޅD�.t/!��牂��OiOR+4]l�@�>�$V��g�|/�'�g"�����;�����
fQ��q3����rF�]�	ֶ����PwO�$��gؘkD;��O��h���D�{��̤k5Y8(np�����?�������y���Z���[���$�\6��A���{2��m]�Q�W�|�'�V��7H�<�}p\��n�ޔ��ɽ�8'HlU�}CWK�*�5���Hl$N�j�΢��� ��o9��uϽX'S	E�3��ū$���Q�^(�:��"/?�qE�!���hK22���m�Tn�;�E���Pq���A����J	����8�ر�$��w�������:�9*���4'�n�E���CF��؀���!�킽4��b�c�~dz'ۯ�L;�2P��5i	|�k)�g���t!�(�`s �8�4)����f��w�jg� ��r�bHrjHҎ����@���
^3���I��(v��:>��;v��rr+�����q2�_�{����4���:h_�z+����|��X썴	 y�nRI��zoXy�P��s��^'dwFkSP�A<�g�f��r�B��e]�ǌ�������������f���0P��v��
�����Y��X�e|k���t0*���Ǣ��F
J$;.����������'��lQ�K��ւln�_21ټ��k	�1���Z���x�`�l%.86��.Co��Q�iw����;'�`��1���%�~����q,���[��-L�VK�,l�V���q��A\7��c.�w*�6y�OM�{[K����d�>G]=\A��"�؞a��j�^�d��b́��Z{�5o��Vv�zu��U�G3�V�>�Ɗ�:B���7��=z7@*���<����5gq�t�2b�?Ic8ƿ������۳�_�>(�/L �u��z8~?��A����E�4ٰ��,Gi���3���2����o���KZ��Zz#�v*N|�������%_U�W���'��/J5���5ź�$�΂]�('��<�dw���u����3�gp�#� �JH)�{l
m�'T�,Z�P�2����y� ΊھO�K��
y���7�}�D�s�E��L�1c16���W�(��D!���k��M�HB���K�]���f�R;��D�X�0��{*T��Yӭ�-)2M����-����+�$�s��%~
u�UD���.�fRF\���ZF���������_�vS����𫻝O$�,�B�=��W����/5���`�����Pqo�\|�nJ�3e@G5�5k �o� 갸�u�e��*�ٞ�fS��!ȣEK������X�P@���PRA9������j��=��}@�F�A��K���~�0<����v*����U�ğ�JO��^�8z]������%��AjӶ�ͥ
�޿8)1�2P�t��� ����A�
���da��~��D��Y����u]a;IyϘ�T���x�k~�qG{A��I~�����H��G���Q٘�p$�����L�s��"�zc���$��O�৞ٹ�D�m��=�n2�0o8=�:��m~�:�fhl�v`Q�PU����մ���瑛������S�yg�ő�ժ��D�8#x��u`�����z[���ə����^��e�G�R���-��/�BC�ҁ�M*�5*���̏��{)�ٮ\� t���1uAZ���	�t2$��B,�Bf&0Q�;���R�����7ʲ>�P��w
;��Cy�0O|ز$�3Hf�[��L����`��{?��pW�X�~��\����f��ގ -|I���;S�w$�54{���bP��`�'Ѯn�ڃc�q����y����I��|`,U��{ľ`6��4��r������|p�"ΌҜq���r��53ߞ��8,��e����:���x�B\��a�'��pI��S* ,�pO�+8��.(�
�")�8��.Cm���ĭ[r���=�=!{.��i^���C��|I�˺@=��3�I1�X�){���A�m�=9�9γ���e+�i����m�'�&���)�H���A��(��{��]'S�-
})Q�xp5ۙ�`aeC+sv�� 7�s�IX���r�@�|gl �t�
/I�}}�w��[�׆>�y�>�t�Ɵn��([_��h�{g��<�-�m�A�v�GB�4$^2�r_c��u�a�� _��O��MN�i_ 2'��1Z�x���:��w֗͜;w����!vv�~��;��?ũ����}��K��?a��+�d��	�J�=��q�Ԅ�<X���r���:#�ǃ-���*^A*S�'ȇ"x���f�S���
���cʹY1��e���Qo����w�Y���èb�?��=-`�dy�@ߩ�W�dB����Uס϶�T�)�8n�?��#$#�v��@.��3}�Z��Ⴣ�6�}_�EcO�)�����e����ϯ��@��~z�=���.Ic+�n�Yc��s��A��4��'�~l\�� 5������8IH?��Q:o��-��+%����iU��a�]�5+�φ�*��m�
<��J٬�ǈ���g7!�:��b�lp�G[��5�E�BN����p��:q�Kz��I��r_��ڭ�l�
-����^����m��HM�r\5	��:n����HR*U�Ɗ���N�u�r��Yjv��R�&h��ǟ�.���w@�(X0�;y���}���O��Ѱ�i,�e�s��jRY�����H���bh2Ǖ�ow&ZN�{��X�a�]�e��|ѹ�T���W��-�{66dR�Ks����S��%���<+\��:��Q�pElDn�|3��W������� ��	ߦ�}!��p�u4M�>g�4��8��ʵ0W��e�p�q"��\���,/��Ɛ���e��J[E{x�)��x;C���r?�^����w���'a����ߺ#��0���ވ|䠢p�]��e�r�ӿI�ǻ H����Xs/
��x˗cdc�Vݱ_M��W;� �m����4!E��@#�~
�'^v�)1�J^�+��:�N���c�å�\<[>{U� #�N�G=����ؤ�tk��wpW(r��T�J�����N����!:H�TmEw�K���$�v�`;V�;���M��A�8����X+)?�H����UJ�Mn-��t�ApJ�x�E�n�Z�ܾ�1m����Gq�NHxN.�Ձi��x�d�OQ���:s�ܞ�0��[��qo5A�����x%�pF7�ﱪN��L)$��}�6>2��K��V����5*�F��+�BV(�e�S6�V�\K_�: �3��l�s��}�$�kb��F���mJ=w0I��e��z�dRrәz*E��lq��h�rK�
�s֘�3j���I��4"�TN�#�\9$�.�gΣg׸V�9�B=8��)������9�wv��B��TR7S5t�_#�s��Q���z��g]_l�.P�}��մ�-�z5^u�H;�5�Tu�ݚ+q���7��'�E�m0�]�
۱
���QY
���:�uyc�xFp�!���Y�^c��6V�ZE���b�`�1ԪG�M���D�ml�oĴ/��O��K���aH|�f@K�y/Yſi(Sd�t�[��0LN��ȡ|	�^��.S�eY�=�� ��c,��v��|����)-��|'#�{��%W��E��e�虅�jOW��2AJ�Ai� t�{�@J��
=�GA��G�N@��袰]2��==@�5߹���P�DǐG�.�%iNE�@\�4��$�%
܋e���4D]�����W�E>�J�3Ńf��F�IY	W���<e��]��o����cȲ��]�������O-yO?9 ��<ggO]��ҁj��f\`��AЄrj��i@k���*�Lj���iH%�"���$��ǎ���;��d��)�(���VFl䐜�4��m/�uCet�E}Vp苽~��)�k=��T�r�S�<kz�c����Qr ���t��U=�t���Wk���[KM�ƈm�r�d���`���7<=�4h�I�ׅ�a�̒d��M��cJ�<Z���Ͽ�Q7��e[C�&h%�����'v
��֞fÆ����h�b'2��#%��l�Ⱦ�	��V���c������	M���Уp�b��C3���5���q/Mj�-�%�<�b�~�߀�\QE�8��e̻��FEt���4�/F�&o��ӗk��ȟc��
�i�΃$to w�i,�vh�f3��@��ۄ�n|��2�F���Â���򓇳��?��Śp0i��
.��&��c³L��.�@�� �(x
̇S5	�� H�%RG-W�o�[NPu�5׻�	nE�ʍ�$z�������=�گ�p'.hZ�R+�Q]�S�<�����| A׫�8���k:5���G�Q�Ѭ&r+2/ⅬK��¿�ց�x��u"���a�@No��д���c�J�+��O���l�؃�۲}jh1�,��X��sG<��LZޡ���Pź���6G�j�OM4�*�'�o�4.+�S��ɢʤ�p�_�6���X�eC%�\Y�/L�@�)�9��^,���uѝ��VWY�: ÿ(�[zoV�-�a�RI��T?��l��>��۾�sj4LqB�ן�:�r�E�'��{�Gu*��E��z��8	�*���8߾#�/j�U��јB�Ms�a���V�GPΔN%�q=����򿮵�h�g���#T�y�&d�7�a"���%��[V��"]�
��5ƙ�!mt���4���$�lˇ�+�"~���g��P�C�K�X��Р�x�΍D��\CB1��T2������2x�ݾb?���k�.�ˤ�{Z���DA�i��=�]AI��w>�k�������5���չg� ��կ��{��]��L��]�:�h��!���lj&��:v4f;Ddqe�5�5����]Y��l�|\?* ��W��pߴA�E_�E}�)�3�4��?�/l������U���*���ܴ�O,��z�O1�>�L��I�$@�����p.�?�_����܎�\��]�T+��]�/\t��a�c��/��؇NKM�
�����D7c�+��?��U�Mtr��b}H�u*��;復�M��n����77��۠ ��}j�h1H�#�8���@x�W�oKj�Gx�3�O� "��ߊ�'��F�鴺e�S-�"�)�5QY]���#A0�{��pP��(QL�Zֺ��Á�~�Ư�[&�'�g%�r ��Cv��4�c�9g��>�B�.Jz�yTr�A�ZK:f�~�!��/G�/ ��� ���g�<h�b�S�!���y\�GM^}؛����p�Ol}dJ�(�S!�\�Oy������k�!]��Y{��ީ�[�	��OĨ��0�f1n��ǒ�jn�p7j֕S�`����u�=�}چ���W~��EaЄm^�I��AH�Z��uC1L��G�A!��]���i�w<(�W��j�x?����Ta�`����;CG�#���R4��@�)��Md��fD�Y�� x�{5mr��\����;��4&"i�+q���[X�x������y���yS8�a(�"���w3)H��*r��y��j������U6y��$G:I���0ei�`�e�ο�~xѐ�p�	�.�D:#XP�Yz�?w����Jo�'ki�����-�5UI,FY��p�<[���{Y����(����
dʚ'�&>��q�pb�ʿ�
US^j����Da��L�MJ襰R���Q�|���w�qk��Ѣ�{}����:�,��̟��a �l�8z@4"�n�֐M��a|��آU�g�*Y�����n�l��gu��<{lx��¨gOj�ZX��S����c&D�� �5�>z��t�w�������ef&�f�?��Nr�iv&n|,]���eIY�[��dd@��`ݒw8���bw�S����"yH�^��(������jc�+x�)Pk֟���zq9�sn�[�> v9�WLV��������Œ�,ʵ���ޱ��,SN�ȩ��dH��v�b�|1
M��F 8ږ���\�T�����*��,悜Ä�eS����)?^�^ι�M����?!�S�M�T̏��"LS��ZA(+��&6�|��vK?B���[������gߋS����'�9Gk�}���1�Q�l�'@�:��z%��5<p�M���#�2�6�Df��c�PO�4��g�}�X��:Е�B �G�z���oe�~���j��4��Tw\��:��t��6D��Og�l�=0���eܻy���P�����E¹]"��7�Ԃ'-������$�Q�?�W�о�d�`M�=|��B1�Z���k���RG�J���r�1����l�)�<��^�"VM��F54I~�����
G��8	L^M7,�@(1���Nq�~X0�����j��x��D�zۻV�0Eb��g5q5��K0����:�!vyI�3e�U��N����&�ιP�4�A!c	O����1��d�*H/x4O�{=|���� +�,�Ei�i�J��33*��4��Kٸ�r�x���I&'���m�?<�&�{�T:����2����n.���4|����_\=kQ��!��3$�@�*ș'S��Y8�;�S!�Ed1*�1�����OL�[?�$Z�f��u�#�w<0 (SOGS��{+�]���]D�aƵ}�d��H[݁Wj4��7X6uc�U�g���	c�֮��*5jKi��h�S?�iUĮw0��QJ}m�%L�?��W~	ʭ��-sb�׫� f�%d4�:�1���O��>Z��q�-t�1vN���l/k�>;�_Tו�xc���oo�F���D��ؿ�����sK��t�t�$��� �KU��'Ex�诰"Y�����)>��h%�[��}ed�z����kE�n�t��*�Оęw ���V���/�/�<�QN���=L�[NˏH��n�?Ièۻ�?wR^�($�Ɍc]ʰ��@����x��䶱TR�8"�r����5�IR�՘>���`�j���q�oj v���֡�Yp&�I���{5�[�=�eƃ���<$�Zr��CO��?��I��e(���	~�8�O��Ԩ��籏D����7{�U���z�4��+���I�6����t����0���-�fnl�?���X���V�W�)̦~�)��%[HW�ۊ��O"�iD{5�̮݄[����s�z�
%�F�B,=x�y��,�F�Ȅ���"5ƁE�EV�
t%����R���{�eB���q��6���_�h�ˉ�|�sHh�����N�R�Nzsƙ���yM��j'&���q����D>�m��G?���p������D�E|x�:Bc���5��!	ud M(q�@�˲�9+�A���3Y��� P�L�b���!ɅT��֚ꓽ�#�:��1D��}
Ǫ��	.퓇�%S�ſ��bd�6RO`Q��b<[~�TD�1���x�������Y��Vn�k'�<H��Pn�|�O����<7�(���DLs<̈�53/]��*C�������^��ǌwG���7^s
Two=G�f�?��O�ܭ�9@��C�O�G�,��K�u�S��bS'��+o�{���:/��u�8�n;bB��[�L��3��u�d'l���k�T�>	���l�t[2,IY;Պ���]GGm�p���D=R�y�^-�8@L�. �6u��!%�(�&'�r�m�i?x��b(*x\M�W V���^�v�;ipS��=˧hb.=ޙ����p�.7nBD��o(��a�A[��&i�8�� .[=��C,Y�4�.�,��������qMB��I�b��+�T.[���$�0'a�1_դ��r�86q`mZ�L4@ft�d[b^�������n��k�B�i� �ٕKc����n�"���pJ�s�@e7ǀ���=#�/6_�r���܌����[4�&�/z�/�w�PMP����,�ɡ��z��g1��P��bO���h���g �y�B�����kP7�Ɂ�����aұ�8�]������������ވ�0�L4�^�G#|%��U��k*��8�ҵ ��!=��F�l���ɶ
r�g�f�jIϥ
�30xZ3Pp��&��@�K*9���x $�Ж.���I"�>��R�l��x�Zw�=�j�A"�����XgLi�C��JC��%kgG�+_�1�a�ղD�5wĪyQ��:i�𞞑�@WO8 ��_���5��ʥ�٢�Ҳ�M]��'�ޓP*Go�PD������Z�r+cgbѐ^�	bһ��"�!��7�)���0����>�b��Q�%�y	�ub&��!��mz�h���/qQN�wu��3eW$<K-`Ye��km�%vV��PFf&���o�����G�C>c�xBp�Lwr����^��9Z����=KG���,����@�2����PTt-|b��TT����S �H�ݑ�tw/���w�#t�H��M?L'�ĿO��i	�y��I��wE!�4nz�Z�}����*��S�@�_�x��ßNF��o6�~n��3ȘXj����j�ϳ��i'���*)�kw�P���%�2�R�!y>"��gm�5${�K��sIUݿh�w��9i?a
ʷ���ճAIM�8��*���[G�vā;��4΋]�QdrzZe�5εk(��]G���&i+�~GW��O5DI�n�e6:+86.�@P�.�F޿6A^�o�Y�0Q���&��K��pCS��cf���L8k���D��3҈�~f�p�/��'U�Ū�X�e��̯2.���ۋz,1�:�k�5Z�3����X��&����ڥ�M��x�}�,e}$����i�M�5t�1kk��m�j"���e�i���`j�5�c��J<F�X<��b��#��%�j0
F��uW�isڤH`�
8�(�*$o����!�2'�o��ꯝ`�!y���1�+R:�
��:���1�{���d[��c����p(��al�k�[>|y��?V�	*�z�y��Y�s�W�e򷱞m��*��t>($�����'������]s�dXF��`�]���vGp	:n���yg�dӁ�ZE��b�ZF�#}�;���W�^q
�F��%�)ݖ��m�W�j����h�ip�L�asg�)XuY���J�Z������v+��L�N�wq9�Cq0���`��#|�s�3Kgڽ�7����f�I�WY+�	����~�L�Y�W�N֩=wGL�2뎛��m�n{�ʵa32o
�>�U)V�Q
b��,_�T�5�\�����2�S�i�@�Ӥ���u�:��`�=K��Q�+�SB��m��z��E��򤓎��G;y���J�}/L�c�fn���Gˏ���'����С�w�����B]���m�Y���W��8������'<hZ�� w�
^F�`���K2M�}_��_*�l���U�j4@�-f�z�2w��,Ǌ-�������K��?�����h ���� �A�*Z6qc"�7��S�..���g~"�:��9�b�8���V@3n�i�y�d~��&�m��8~���<�S��G_��Z���S-4N{�s���jx�NxV�Nj#E�>dh�@�]!B��<#b�iG]�ǁ���g:ܻ�|έ��H6v1>2�J����>�K�>)���(���%.`������(
�H�_ct���6�v8��3p�t��*�ɕ�~++i�i�lճ�/�X�o���#D(o�8)�'4͵�>���vN�r��`�@����q;ӌ���-�VһR��r��3��i&P���56hÂ]���V��
葏����E��QT����wH�R�H;#}~Ld$�N���������~Ƶf������.��,�'�^���1F�f�Ұ:`���zP/���B�:�b�3��SCu�)�p��+u�`o�U�N1��w\>z��5���A�����?�́��砼�U�Y��M����|�	���*�E5����Tߡ�%�4�!S(PE��!N_���z����r��g�� �E�)���u�+��:��ی>l�.a�]�����+.�`˒�ER��P�8�	��R����Ʊi7d���Y'��Oy��1Ay�H�����q����D�t����>"*�!����@QD�1���B�v�W�ܝ6{V�=�AfNf��0'wM�]{f-�����`�h�����~��Rj?��\3�5�Z�i���r%zW�r�İs��v)�̦��5���'%<gwi�$���G�����e��,[�� ?��`j���@���=f��s#�JjGa��U�� }�a�<�j�A 53�v��-]�j w�OAJ����@��u:����zdT@�#�S��[X��Y��F C5^�/2	�f*��s���O$T������q��C�P����G��i��}�A�\ۦ=��̹֥�@G� n.�6D^����w�CJCb�+@�i7~8��V���pP�t�̇���
^�$��,�o�s��^�SXc9����
�:�����8[�����}����U ����W��˺�/���8n�gx	��a���������Q�E�o�|8�%��`<��?�b3�38�s�s��՗�
�(��Y�y��!yM���Vj!�8�mZڲ���	�&C>�n<'��bߝ6<idn㞴/tr�ȆL�
.��B�����J7�5���X D#�V����~T���&��_>���2W��@K0�o��N+�� ��G`�c�*\��L��]�t�	�������"1��hr�k���h��z�}�qϺx.M��1(<��@�a�Q�-W0���kC��Q��!h>����FH����\g41�"[,ϴ�'&6��D[�����T&ڎ�U޳b2"��Xt{�9��!Q�6YD��l?��ezV����a���o�|��	Q]ǟɷ��q�p�H{�o�n[<�u6��@�LͿ��y-7gaO�M��9����DD�׹����rt2�*��z���65��Z[�1W�x�C ��hIS@���kM�����U F��,Y��vX+ԢT>�]`�xN�N�� �ef��(H���b8��o��+�Z������̡��� �o$1�jS~�.�R���M�N��ޮ�!�(Zt����"����$��q|K�
�	���	��Y䆩fr�w���H�d�����8NB!�p�!�ge�U�/��l�S�ǿu6�����gIZ �h��MM	���+��#��h(�f��v������VR��O���&�M��}0S�nc%i� �mM^U+@��_����-a'�GE�M�n�s��ᙕQ˫���l36�GR��'����*���[7�r�"�:���f���_�T�x��i��3#�-�T��o�[S^�hIJt��C'�LZ-�}|�_�K���~Gu�6�!=����?\��<c�F���qry�����Ʀ�����&̧��z�����O���$�^4T6�*��z�<{��-`�)xV�NQ�7hP/�uc'É4`����c
|�Jin�l9O�|���;�g�͌�:Y��~�u��ӕ���-�@3�j�f>?���1&?F�cklh~��.g�&:1�+��~�z`�۸]v�b��d���`p� ��N�¯�S���X�K�l�SܭW�YF�]][I@1��{ͼ�7_q"��IKV���	��)��*�mr6t=F�uV~2�M���[+�B.�%�+��1��L�m�����t��_��'Ӡ���b<�z�:�[nB�~������o���!���4����Ն\c�7�߯�S\���@MJ5�XT�O&�%'hvo�:��h�Q:<�W��$e3���]9n���������`�IS�*veblTB�K��_>|z��֯ީ�]���!�[��A0����s�o��)�s�qGqH� @��f�7A���L��i�y�L���k�dkL��Afp,��
&$�
�|L�0�2�
2����\'�$U�lk�5�Pr�F���Zs�ep�ǹbs����ԛ�����,�V��7��i� �)��϶ȸ��g6�:�����\� ���dfrKI;���������i��o���e�C)�3��h�_WΥE��!������u����0�����)�T�_����ig��Vm���憘R��m������T�nZ���^i2�����Oe�%����@�a#7t�}���(aZ�V	��6�'�3�~�y_��j=�����T��wa�TQā��8A>�w|/�q��֕���^�����-�vd-�2m5�&+�j��S���R�0�Gru4=�+��{�,�pb*�aȪi3���e�"(ŋP�Q=��F��+�]�@�(��G\�EǼ��c~���[v���%�vf,�b�q���%,��S������g��������W�Ǐ>���lY�\�N}��f�`dVf�L�&'��3z�lak�/��ξŽ�x���ҤP����ĕH�T�-��#��"!*��V��o`��Q����9���Qk�V�*�<�{7���|�PMZ����F�6I�o��\j��Y���fh�1�$��"O^dWIV���썂1;se%�PP�;n�o>�j��
��偉x#��5�0+}��$��9&�o3�x���ȴ�B*��w��`����~�ҋH/�KSu�[)�����c(<���1���Z���N_���)z�)�{m�j!X�(oi�Χl���bA,`Ũ7����� qJ��o�GS��n���'��I,
����D��ޛ?9#�\<��P�y��."s2�'���L��b�Ǻ��&#��������w��t�l�Pےwu��ՄAu1�� ����2@�.<Ry��;K����v�[V�{ڒ�;A��	?c�Aŉ�q�ؕ
n�ʛeE<�.�~r�x?(��vɡ�Za��B��7�ZQ:�H3�o�߻d��׳H*gq�ڦ��ދ�����ҦL��ӖS�1k�ۿAZ���X�	qt�ho�;B��	�M"0�]=9:8��>�]�Y��Sn=�4?F��z�__��ַN�^g�d��N��Y�I��{�g�[�� ?4�	�E�
�J9[�?X�Uݿ��
��(�$��з�}���i��ҒA���㠶\��R
����1�mQQ��]]�8C��V�&W��g㈺�c��Ǩ+}���] �*	m�z?����,Y/�b4˝��7�m��� �m:>_��f���&ݘ��d�E���-�@w.u\�U���,�)V<.c��yk�-�Wa�󊅄?�L,��]�WS���4NO~▜�W�c����̣V��"'������KY*I��Q�g\;��(/�J������}�,v��<��u�� h�Һ��{���`�ސ9���W|GM�L��֥b��>�5����^΅X�M�1�9�H�#�-��+1������6 vbeNk]"S��oD�p\�Q��n�^J���ݼGw�󆱔�-C�9@~��΋O�'`k�b�Y��tX�Te ���l���= �7
u��������6K��D�&lԄ�������ՈM���S�JZɸϵ��`_���]Z�7�J/1�cLJU�2r.D�k\�\f�1*&�,z����VƤU����s��{�.�c�Hq��-�|��(�f�!�dO*Rs��~�|��b<j��^���Cak�s	t�b�P���c�(���v�|�JRe��,�,��m����P���T�-�8���l��"�;�W�iQ��s�[�N�Z��`S2�(ν6=Мf�o���gԵ��X��j�����\ �~D�C3�8�G+��*J�q9����n��0�?��/���,T�6�A-u2�w��:Q�q%�8�!*_Q�$� v0R�oR�[x�O��?��-#���}�^z�M���?tbcd��1��Y�C�>mv2�i�6��Ǿ���"u�lA�]u�G����A�{^	(�Hm�$�������G���y:�0�W�1f�Y68�B@e#�#�`6+�M�g�z�GBΐ	n �����u�Ey�bڊ��H�~.=(iSh3���vήb���U�����TU$�=ra��)k�+3�vKѕ��\���N#	g@�rX�o��~�S�L��1�mΏ�����Z�y���A�H��F��ϡW���-&ŔCf�e>Mw�Xɑ&�(��]���&pvӱFȨ��f�Ji�[�j�C�F�t�H�D*<q��"g-�u��ߗX�zj�>��*��(Rڹ����`t��zF@�HegS���?)���yi��<�P?����"+T�	�΢�B{�����Nn��7���:@ ��qFN���f��h�u�Ʊ�	L��ͤ��q��l�x�����AFt��0?�N\���;#I�p0A��`c�������"����e3�=�_M$+�-�2Qm̠Y~-��F&��(0,<����4�p�HxN?�)��{�T�v����=�_H�i,��3��0t�[�Ʋ�-�Zbv/S�-i욎�3�>S4���xpk�\Y���W�����Ԧ�2�5߅��ׯ���w`�z��|x�f4:
�266R���;5�I��4S,+ǃ�w��
�t��SY���p�y_#��sY�����S|��}�E�p1��-�'�ؒ-�$ �j�A*���!G��_+���R
&a�/��8@���V��$ə;�V�8Fjg$I�.�>G����`0:u�bX~Ԭ�襰 w�b��D������벿��2�Q��� W ��>��$p��gog����E�=Ϊ�c<M�ն�.�(�p��R�P�������G�Go�}ӵK� �+�\.:�2/�qD�����c���0cz�s��^�ǝ������i�vxF���nA�i��I�ό�n󫶷����+��a��OuY�6�������/�Vy���ndbV�����,0'����
9	�8i �c}�R��l�ϙ[�
�~P�BB��2HUzk|&�Ԋ ���_7i��ō��:�!f��~�~��K���`@��N�(����w�AB83���E������������N삻LQ�w&�'�X�h��@'���@��*���B�{���b�If�ǋtV�3�_B�� �����:��������X��T�0�pb".l�N��q7�wO���c����˽;T9��� P������=Nf� 7R.of�\C���2�~�k���V/�v��4���N�e���k�5㥊b[�cZ������=T�{���q����<M4�������k��Ȇԟ�d��iY��Q�(�D}�
�V�h|���чiD�՝&���eJ�2 ��5��M!�R�0���w�l�m���q#,XX�@::��%=�~�B̂a85�ɹ����ag�'7��*֛j)#�����o�$]\>���=��D��VL������E�;������ �h3�(�w0V!|�a��u�6"�S'�[Wnj^R���s�֚��EН�q�ͯ�Z�.o��T4SH���'�vmZ&EQV�ɷ��#sy�~�����V�߆��Fܠq��Ш��E~�,!�Z<�,Ds�S���oz?��QA#[>�������5DX��O"�Ї��s�Gkg�PRA�^��3ot��G��Oh������㰲e�`*韹�Rb�b�0�V�~m����h5�wZ4(��"����U�p������b�4B�˼&��TQ��g�}���o��]e�*+kr!K����n��NY�`��µ��^�rM�`�+�!�cJ�8އ6P���Y�0.��^|�
�G4�3`�SZ�h�$l�8�<�� �<^	�$���y���q�dȟ��Vb���@4$6]���Tv�����h������p����f1d`�B��r��ьZ��{꜕A���%�$$��Z��<����I��9��[�QW�~P�O������x��b�W�{�O��t���(#�quol��%1�-�] nM�ʩ���34�%� ˪ϗ9���0?B��bȵM�~ѡ�u��r
�Xo3�������e�*X��|;�xW�}��	Y���Ay�HS���<���.:G�>�O��F{�^5��;7͜��6PX����6f�V+�bU�l0���ć�K�c�Z�t���b�]�u��]�m�p7�$5����oWP>ὁ�eF�=��w���o��C筙���q��(��m�K�R�Бt��"� �p�a:�{��7�<_z������a��mr�Nп�5������Q�V4m�o+�i�u6h��/|��.w�/�B����2�ZB����j�:h$n�����X:�E�F�$z�A���%��ؔ^[�
�X��c�x�$/jj O d����)���Τed��R�MU<���,���Ak���1-b�*XD=<��j1J�G�K�"S��0�J��b�V�̕@y�_�ۅ�tJ��l��T֬�c�#�n��Qk?=���j���[,v��\X�^jPa��6X<�s#����(�Hlb�}�*S}���XK���'�V����1�DX� ���ۅ�w���[��9%��;`�+�ğ�a�(lll�>�W���P�1yx��� s��Ǒ�A�p{R�����sn�
OU��+1�����*�6�؃4����Zi|�)Uĥ'���^/�ꞕ��z��rb	�V�ғ+��5�*��Zyuw����#��A�x�"wf���y/XH��������,s��*,� �OFP�2hp8e�v��������9�}y�X��o!f����OuV*�\�A���Z�҅�(����듞0�����i��(bH����(l�o�x�*z�nz�"Vr��|�f;����+��`WB��ȃ=�V`ˎ���zt��Iu���#��d��Cjw���pQ���� ����+{!,p�	���ۗ,a��]{�����V�+g�*Pf� t�;�`��J���niSg��{J���u��\��W�H�hU�Aк�/u�
�yt��x�B�/�bYk��8b���:"}D�N���m̝�P�����>��V�
�;x�LnhZV	c��C�X�I:$��h
�zi,����`��q�2���ђ����K%�z�b��B�����vO��Y����2�/����'�!B����mua�w��5>� �wsNa��Z��U��P��"��y�2O��U��r&mg�)��t��T�]_��L�(���HՎTƿ�E�����_�ԡ"^K~�9s4PTO|��*q�ԀQ^t�Pa>����>����x�YW�z#��zz���Z�^��L�ٲL��v3z���n���0m6Ub�r�S����B��t<ͨ��`�@����$ee��";��H-��mk�����o�Vr`@�E6ñ���(|l�2[h[�:"�P�V��{N�IX��ɠ��4G�=ԎA6��EV�y��K�DU��l���b#[�SW�t�=��������b�f3���,��`�0�"�l$�KI2��܇����y�m��>�8E68}�D
������P��uP�{�`�A������\co�+��S��(|�r�� �oU�l!��_
�4�Zm�`3��������V	���7s45��C�L)z��	J�����Oȫ���|�����K�JK[<i�x�La[_L�d^�XB�~M�/��E��`�"�25O�֬���Au*plN�5		�tB�.���1Gi��T�Ȱٚ7�I願�H"��Q�3](.}��|s\#p��g�2W4jOszIH,����se:}"zT��^�Fv���@%:�-jBFs!W������*
�3��J����o ��7 ��OT�����=ns��E� ����z�r�>#L�c�nH�l��z��cY�����rC'�+c����#$��~x��YL�y�I<Ғ�w��� ׅ�]�a����^/_0Cޥ���=�d�l�R�i F� IT�8E����Zg�h4���i����¼0ҡgqz-PK(�J��t�fedp�#e���p�
�����2�8�6�_����&�3/�>�`�q9��l�Z_���8|��K7��z +d�R�%H �8i�掗��;9y�$�M�?WPj�/��	~��V�,e��| 2��� �	���3�q�]��C�Y�T�F\���(?��M���P�>;��[��@	����SS6�ޞ�V�y{��K�1�(����� �yV$�А෡.����pY�-�n����j0y�x�`m��}`ww2A�	L^�0IS�������k��V<��Kc���6�]e�'��l`�J��=��2� ӌt�_�]���&���h?��d�D�%H�<\�R_.�*�QA���z(@�%�`�}�&ᒯ����C>(/�
��{E�~S��Z}һ+\�X�ڕ�8`AĴ�Y��(+�.��� {NԪ�X�$ּ,?��Kdh�� ~�����a���A)��c|�Ą�
V��Z��I4@�ӷ��Wnn5g��g�XT�UN1Й}"2$���$�(��#���!;�˅;g#c�sz�VB]�ف��g��jJͳ�P *���BX�ɉ&Uq���TU�D��C��Ԡ;��N~3����K�g-RF���s�	�e�r�l}js�9�T�H|�d@�{�ͳw%Ǡ�1�$P����Ģ�������_��4bO�3<��O���i�>X�����H�G}M���򛻿��j����M%��R�έI
D 5Й**���Z�����&7�3	��n},{3�K�\����P�zWf� =yr�3����1[�I����|ð<{s��`�(g���J~���r��Wi�Mx�'~�j�$ϫ\�F�����WJ�}�S���n��F//Q�#N���!F}-V�%Q�����}�6��	��=���XU;r�� �+���6���9�x�q�@���Y�H#�Q�l�D����to���Oޞk��n?. |��Mti�#�J�ŋiX <� �}t�s�%H�|����W�é��_4'�:D0�#Ֆ����f�I%��Adp���If=B����E�&����s4^�]�D�YQb�y�~脒_՘�) �TM���'1���#���)�s'�ڞNW��`���y�*{g+F���C���(�?8M�����|X�����i�#�.t�GT�� g�)�՜�2\^�g�w���rW�J��?:T�7)��w��i�:��[�.3)�.�xȳ���7��vH۽��v2TIXg- ��N�pO��B�J�OΏ�(�� �+�*�q�rd�����7�Uω�ʥ��>Wf �{^Eh)=�À1����B|Ĥ����{h��sgU�7:^V���R��ɏ�r�N{>��'�(�609+� ���؀���O�:�\e7�\��l���m�<X�"%�IWҲg���qT�ҝ;P����̌c� gU���l���U4\�((�VaT,b�(λ�+?���ј�sf��[,V��z4�����ELp���Q�0^�I��
�3e����?Kf<�s�R�6�h�,�mA��9��!Ul�*��ҙ�y)")ʲ���'͝�XȫuF��v��r���m|�i�Q�4�b��ߌ����Wu��,�
��gx�d� ��j��r�6�3[��:���L�F(PB�
��t�,���P}?�\&�p�y�oLa��;�VzD�/�n���9�,�x�Q�؁�1^Y$b�do�(��w�O���ꈷ'�ⷑ|j _�)�7�D�+��,G����¾��,t0����
}�b�0�l��c/s�l��ثY-��0���p_3t�\��Ӌ5�莙�a)(Q�l�����/\ό��~r8'�D�4�K���(��
�̹t�e�ٗ�ku#�����g�|1�ޘgB����'�q�%z�(S�d]�ˇ�!�W����:�ݮ�E��+_�� UL`p���*��~�_�}8��.��H(i�+p^�
1��Xr9^Zz�<���rc6z꣼$#���]�Y�v�2R��2:s"?�.h���Qx�Ԣ۞��X�E�Fx�v]2�vN|���Qfr��8�:��V��|'�2�E�U�9�ZT�S8����gt�����r�����goZzQ�k�\0k?�q�����m��KT~��oA�M��ĿH*����)�(�Ep �F�$ԛ�{&O�e����f\{�&3���P��p�$���ռ����Z��l�aT��a� L�8D���!������S&����(�w���\;	a�ڝ Dt��9dMU�㕢)M�ҫ�����!�Z�T�&|zH�U��k{��Z��^����g���]�k��O������S@����l��H�跃��B�:	�5S�;A,#RA�$W�dPM�8C)�����o��ʰ'\o.��rB�	�4{n}A�|܄t
S)x��Fk`�I�@��V nȣӚ`oʹ<C��̏aCq�A�jZ0&Ńl�ڪ����IM#��=&�.8��|�eܲ����5�;�\Q���'[bYߚO�5��k��bB�9эu���}����4��׉��Ll�^??��4%6�1Y �1=΍ f=!�Ae��s��0���� �X�=m����S�}������A�y1��d/7��*ҭ�+�Z�w�>�&�T�ge>{�%���.Z����\��������	F�,%�V�C�`Űfąr�R�t`�G�!N%�L)-+�Q�d�Z�Ԙ�i*g���O���V�,�Cf�`{���A�5yE;%���Ly:������tAo P`ę�Ib)%��c�Y,�M�W/��C8e�2�%<Ba98h���4�f'JE�тxͺ�ŨϾ�A�zp�_7�p�<��y��e�a�:�p���g(���u|l����]	�|I���8f�n�����?�W�t?�d��l�ԣfp�+����8�Q�W�ע����a�2�̬�����~���tB���Ke�g�6�,c����x��B�������������3���=h�R�_�;ט�[�r���!��"��Q��_��/p�����3o�.`R$B�~����f��{����=�i:�k����T��E>��j�����0`W}mx4�!�z���b?���Y	3�'Aj����8}6�z��-�ތ�}қ�T�}k;��*0d�S�]#hy��,�.﯀԰��@~E�4,k���2�I:x�-��jg?���xǅ��C	��z�]?���u�z<}c�[��md6�(Ta�ޞ��M�����[?����6�ZM�J}'�2��1a��.?�j�o��;��� .�����ֹ6[ZL���,���i:B��u��T�lPZ3a�6�\J�l`�Jgu��]�@�n������`�S��^�i.ه�4Vc���j��ļ]�`�#��[m�&Ee8�UB'1��HC�#�'N��5ұ�n���y3$�e	6B��[CHG�:h1/��������ʾ�a;[���j{�<�������	/�kE@ԶB�%%�a�"�t�c^�B���Mo6����PP1����O�5�z~S@��<{"<�e#��HC�Ps���?��y��?��u�o�b?J�O�Q�E�M0`;y������!�|��h?>@h�iТ�]	z���wַ][z�?B7��.�r��=��G>�w��!j'��XE��� y<s�F�ue��^��n���`�̞2#��&\���Wl����9Eq~1,�%[ɍ	��n���i�#����޾g=&*%P�~�-�
�`�8uBȳ,���O����*����D�7�a�i.������W�񥨇v��"?�]}��Gv�<���wzgr|�u�d,�^Տ�ǧ���l�^:߈/b���=c[�vb��U���/L	e��d%���������*���g��SQI�ʎ����^��˫�:$� s�A���Z�b�b������y�(�7��vM%�O�Wϱ�����Q��&y�p8'�r�u\HK��������D���%�'ix*(2`#�=cOu�eܲ������
ui�#i��,\�4)��b�n���\������C�/�6Ձ�L�+Y�9���~s*�'�cԹ�]�o=���7�>�i��I���i 8\��է���Me-��@b�$�ߓx6����i�<�P1=z{ TQ8�I�ￄ�*�a-H��Ϻ�)iX��N��αu��N�,9��Yu��ҋe����!�v���鴹M9�����K(e.��lA�wr����i�>�^��~j�8�޶���g����V�]�E�9N����q�r^�L���O���;w/�ؒ��W�
�[�Q�����ۓ�GfI����x���e�zQ�2u�M0V�F��H8~N�F�R�ZX1qM�Z*��#�6g�۵�hdo Q�+rzX>c�rQU�tC\e��u��1���\݋#}Tُ���\�o7�ﵲ�d�:Oْ�pEYwlejI9/�)k��2��O���l��[�����N���*Ϩ���gB��3B��ó�[6��ǲ�6��i��C��:`\.�f󅆈�3] x&x�ᯠ>��^��3���%S�j�F�2�fV��{���)���.J�{!��'�6yx,���A�>~����r��p��Xh�d�mB���u�qlz��&9XYh�[;1������|�c��(�_�aR�V�����'�����Vi��jc�'}��A����1���3���2, 9iNT�d�d�[�-|�$�	L��ԍ�;��� ������w$s��rД��1�~� ՛�Y-��W?�G�<੾W��;`���m�~����?��L�o�o�f�^h��N��MT`Ӫ�Ʌ��;9V�H��.�|T�Hd�
Kz�x]k�|i̙O�kʥ��؆��\�����1!���"��!��b�'|k4�p�^$�5�Ou�H��^��ꔴ������@��^��ŃW��*X����67��P
�$L�
�^����,n@����܌�������ҍo$��ፀ��۹-%pȯ��y���s��r�^Y4��ͮ���6L[�jM�B5�|K���,O� ��;ME5����R��29\���j/W�Pa�~}���PIt]�g_	�r��K��.Ԏ�X���y�l�5��c1��p�
�l�������b���@�u��{F?mL��	�����3,�]���B9�dw+����z^V�H����r�Hpe��-���U���|b��K�e��`�Ws�f��U��SQ�w��+d���:���ό�6��`v��s^$ny��&u	D�f-T�Es���#����-SV��߮�ȯ���U�8Ϋ�i�;�g'�s����ie^M� ��Eھ&��������qXW�
ǵ�l4��*(�L)�|l8n�/#������"��=O�T�)�w�Sݒ��o� *J.��B��h�7�˫g���81��UM@��g���3ǘB�ҝ,�$_�NO���.Ǖ���8s�����K�ҭ��m������z�8D5>C��/		&ڷ�4'���r:��/.�Ŀ�$Tn���F:�ϔ��� ���"*dZW����r��$bN^H���a�x�f�l�{�U�\��pfr����Wbc�1��1�b�!��<����B\Y�Z�9���^��IE��e�'���V)ܚ�ag�@���䵅�}�Fw��FX�S�P����3�I���8>�Y`�UI=�}�SR3�>��o�x>mB�%nO���
˱�έ�Z(&���g�5��f�-�EtS�!�5��u��S��;��S����
h+���dr�Mo�j���+�_��h�5��mÎX w�o��Zh�� �`�笲7�py���p����9_g��:{y���	f�Xn��L{��a7M�X�{Y	?
,�T�{���6k���Q�����+��hG����"�v�^^	���8��Hb���� ��?X�A�u#��{K���P�G,��y�3��k뾠p"Sd�H����_c%�K���+cn!�� �8
��G�U)c��N
�"��&�c�V<�O?�(ʹw���˺QI�p�D�k%8�e�gR��s}d�<�QQLA��I�˷���ǝm4C����0���9=af�߅�Qf����b+�V2�ۈf�)�"1���G(��Fe�1���͑j �gw�%�x	9��)M~9N��[>E�=��+#3�d�M��}q@�R}�� ��pf�Ȉέ��c({b�@��[��"k�E�^⬊��IW����]�a��)�@֋��L���$����1�	�u� �(�=�U�&ERe����5�^��O�sR���C߭d(���e��7�5��$�n�«J��]�V��D�����I{1���kdQ��_���引6�̞�<�W����
{I�k�[�'�rgu�}��ét�����pwx���'%~�NQ)o�H�BUc?`����]m}�V��;JF��fإt{�d���P����j�,��8s��<�a��WI_8ʋ�W���fn'M���!`�2Vy�T�/sK]�� i_�6�~��$�ǃ�g�� {��|�I��i�0v֭��<�W�+�j+_��X6L�#7\��oćVl�����I�x�+��Mˢg������U�"{*��\:WL�6BX�qc%�MҼSp��~��20�U��$r���$�����!��2�Z���s{��цy���q����/�J���s5,�pf�4o"��(����/�"��閽9�\��tֻ7�
�9��m�,O�*���#������ЕDؕ	 �Q�?=ˁT%\�)I9�(���U����M-��w����+��F~.͈��[��1{�CI�I�.l$4�K�@g$���%������yO�D�U�
�	T���k���f&���>��������\����cjL�P��oq���
N���B_�����9g̊J�0��Lp_
�u�dPe��� �C����
>��9����G��.���I��"(c�WF����}}��{W:q��þT�5:��w�U3YD�ʙ��B�Ee-����C�I?8�p��#�p�q�N�Һ������IZ�G��Ui�z�5&���_n����\�PY��O+��*�/+1��-���G��<^:�f�X���(	Îp"JH�g������]Sp�N�=�R��4�]���V�����x��k!�t��=�*�v���5'EY�s�a��^���1E�Y��4�S ��0�e�1ʓ�T�7��Rg��'���$}���hw�o@�����t�H��{#�㊫5� v��W��ݿiU�hL(k[P��2�{&>;���2��vǆ� �;ۺyS�Z�{z9�"*?�F�V������#�5��a���X�3h���7����,N���6���t��u��o�?;�����c�Gk8g�~�4���/���X�%��͹7ex�b!��S�e���BUE�,�?�W�B�@�Zypu��5'����`_3(QTӸi$hO@�.��d�g���(�<����rE�\%��b�ΌW�!*M��KmP�E�Avppl	�:�h�;T��1)���>�[g���l���6��!:���}ɼj���ar��u6	�6�,�Y��x���?F�,�2��u��2�ö��jbvy8�|X�l�C!���ڏ°��j�ܫ[��X�����tmj���@��O�|����mdF<8����`	�p����՘�꫐@�@ӗ��[֭a�.���
M�L����\�q���H���.�0~��5^ڰr(��ȝ\�$�ᙚĮ�^F��:��7;�1DL�7������[��}�������7.!�YB�-`��RZ����;T}��c۞k%���[1(7�!�`R&t��m8���ؙ�>�:����*���r7�Ƹ;D�I�>�q8�d#�e�'+�n-�w�Z�0[��; �������_2O�Q�]"��N�1��^U�{[W�S^�1T��A1b�aT�חR߻l^љ��N�21�� C�v^����ޭcKz�4r�ެ��a2��x$bU�������y3��H�N7��� ��3�Y��\M|S�8�)I��+�w��D����|o8<�O���c�r]!����8�	pL�1���3�+�x9��4� 2�P�����3�z�;kv�n��.f/mD��wc��dZTn�i��[״����.6�gގ�0���X�r�yk_'���3$��I�y7LCU(���+	|Ȗ�QZ�dg�;׻�
��+��P�=7qB{�) ����M�����aN����rUH$
�j��d*7�R0W9��%gg�V4P�*,��(���H٭D���p3CUX<��O��w ��Be�M�[[�Q`� bqRg�_cL`��<�:�j���Q�E~�ÜQ/
�C�`a�\�$h[���ca6RƗ��З��cZZ56{��7���i�陷�
I�0��r�G+����e���%�<T�]�3$a�k��_���'|�8/��c�H�^�o\�ѫ6J�����A3Gu�ɱ����u0�O�r�ќL�$������{̭�������Oa���������˰�h���#$MrB�U��(����'>$��í��pM_����4��c��U����;07�Q ��/ǽ�/�Ng�DH7��!xt�q�U�ڤ��Y�>��[f�e#�(�J�%����!���z�9x㰌@7��V{?�;U� j0����c�H�����Ƣ_�,ckS*�D�� ��mR'��H�ǘr��d���)2h��G@߫�Hʫ�����p�ku�[x����� E���D*w�te�,��>�X[.SoWtYu����j��wL<�\��}���}<Z�0�kd�5֒���J%�~���k��.H�.a�{̃���JD[��T�F�9��N�o�H�M�����O=�ѷnI����Bx2Ɂ���%��i�M:����v4�A�A8��=�u���e��R�����a�[��n��0����Q�2������x&>��"F;��k�@ �[F�yN�/��|s��\i����^�m��`�}[r�V�M^]�ou��%�_o��% �OC������ w��%���\5(��r��h�`�Y.^,�c�DU�ט��F���,#^��������¨J��T���󴡐Z��ca�F�������6�H[�j�B�����+}>�Q�,B�L�_WÉ�'���?�7�i��p�b�
kV��<�����17dɨ�hA�*�e�p�;(��0�[TɭK{'S���8}#��|Ȃ3bV��C���t��'���Ѯ[��7 ���7��;m�-P�}��7��4\XJW��f��K�K.��k)E�&+��o���bH#��҈p������ũx1�i4�VA��or���B�<�PB.��9>�
����!�rV!���	��fs�2���=�.�d5s���)��|������R�"Z�[c��3�z��7�=�tJ��t��8;C��U��Fb:-���	zN�����v:A��kkۅ�Ç��'plI!}�vR�J /Z���>���c���h03?fz�������_��u+o<$ٱ��whd���2;�v��7zv������B��ܣg��
�P~����� ͭ�\�F ����`��$m�v���A�%!�-��ͼo��PYK7���&)��ʹ��]��f"�
�������@/��^D��I~",��'Ǫ�Lf���IP:(�?���zR�kZ�W�X�7dp��]����|�8�Y
�&PŽ�tTi/P�(X�
���y��%�UG*Ϩ4��OhZz�g�N���&F�b�.����@67(9x<�}�`�>��+6�^�ݵ�" �?���{��s:���Cj˔@��ી�)����)�Q%�qi������d�۠�C#�0.Ԟz�Zӆ6�d�792��4����M�=��&R���X P�����?�.������ѓ����_���?��֤�N�7�,a��|��+<��_���p�����D����,��. �+��Kc\uH��F�i��;�7\�t���7�)ϵ�W�wt]�dӣ�Q���ż�c\�Wi3tG����������[���s�&�M�$��X�%}.��.���ləRK
4����+����3U\�bh��h��%���H���3��T�y_&���rm]�E0�aU����z��<�d`�^ҝ�����"/^"�'�o2����|�l=h����}-�l����4M��r��9��^~�2`NϬ�k[o�O�i���n�d��ac�6���K0�E�O�|DC��Qe�A�Z�.��ȶ�74�ʞ���(��ҳ��=��F��[�:$�s��M_�1b��J�Jc�m���:i�USr��J���o�$Z)���i�����6�C�4i�5rc��{�n�Eg��KGF>�dTsO}�/ �\������u�Ϋ]�w�T��4F'(0�d�|(NIM�J����G�C�t�+Z^�L�</~�L5���H��þ������4����,��1+-�`a��q�nUG}�qM�8���ed���X��
#���-���hb�T �5;�)�¥76�+��R�v�n��w���_��ou�x<������`4�-� 4I/h��Dx�V�TR�0�Z?�Z�(��"u�b7_Doh%�CY�<��4��i�Z��H�9n�]�����`&j�ykGܝǅ�a)A�/������&�����3@7��{��~�Ŗ�ϖ9YԀ��n�-�9��"�*��k�)���k��jO��?Q��� �
+PФ��W �Qn!���h�o��A��|`Tt�f�ި�?'�ȉ���0\N��m�)�o<vLAb�^�L���]r�/l�̷X�d"�φ*�(9׵c2�<]�׹�����+��E�c/�<�����df���Y�mU��T�0h�X�;d/�gr��A �JD)���5J �(�?ٯ�e��Q�ن��.�rK�0g(y��}�����aop�Gtye��Z��ݖ@H�Ҡ��g�#P�^G?��-v��y}w4��Y�/�S�����,a��Ȣ�s)��Ԍ������]��F�m%Z%�SF`�a+�Nr+��ky�����IQ�+��T�Џпh�U�>�r��×��ם)�9d��5����<���I361!8Dg��0�P��|�l2C3S������Je��k&�ތ��i��9ԡ��-�QhB�g��� �?�D]�KT� �O�$�����q�C�;���>��z��Y��K1\���(����wq:�����"r]�:��w�����\�,�[DW×Fm��N��̏N�����������5D�U��E4M�EeR�V3-��'��5�@v������a*����;�ڟ�~���4�ق�$��z6�(B�-�w�_���A����r�Ņ3H�Gm�z���ݐ��N�=�\l{�:�#������,����� j}v��mݣ�&��4�������IJn�Oğ���E��c�(�f�ɷ����ԁ' �ey�^��HbϦD��BC�l��w7��ѡc����L|�cr0�⎹y�>慩���4j?�Y���,��;l�ߋt?3x���
��՜�w��]`�{q8�r�4�����8����.�/!�'L�/�h�8P����H�7cH�:~�}���`�������JY.�'�� ���P���s'|3;qe�9�0�7M��4��|^c�s�j/�t�U['b�!&�V��fG��L諛`T�d+aL�0`�����ˑ�-)��2�G�o.w=��$H�ν=P��a<_I8'���7�ת��6mx���h`+��ҏ�5��͛�@�"��;p8}����b���af�+F�tO%����w���3C��o����:cU4# ���@Y��=���I�[l�L�=۽��g� ��T�65|e��)���@ �/%������rxf� (���{s��E���j*���c��`v�]���x?W��9^ޛ��1u��e���(ZW�y�N�B����$:���ȵ#���d\���I�jn�tx7l�.��j �iڊy�K���Ræ�]i#�j��L0t�$ºSQT�dj���_�_���l�%?��]�s"����JwRW�U�u�
�1-GΪ(t�\�8#���ӦL;��z�Ԥ�.��e>�z-s>'�E�pY*���N���������й���n�4S�\�+��O,��wk!���Uw=���ΐ�	V���\cΉ?��D�E��K�1����|��^e��ċ~�$(<���p�W����(�>g�[A��)q���ӿ+ĩs����=�4����}޼��4�$�.���+���Ai�5��� ��{ʟ�I4�9�<�u�~���g ZN������V7>��Z#�B�W�;fX� ;��ׂ��u$s ���l|@toT��פQHҏQ�t>*�+.�0B.C�y��-�b_Z�wc���s�b=jڣlE����mp���u������� �3�R��_��J3��Nm>�S�.�g��.����8��~�6�蠘(�>p������Rb��<S�^�7%�(/S�����X�_9%��9�K8;}�f�ւ��j�#wG�G0�>���^����3J?Tɶ��`�Q�g�0����D�t���2����ۯ����vn7V���4�4��#���K&�(igZ�SɊ-
g~	mik�fu�K�i�{��{궓@��yz��
�����F)=�9�j�&��d-��-mY��#)�)�m���*;I[Y*R��ȯy]*(.^�"O��W^L��K�j�Tv�
]��M9��yu1{��Tg��W���
!������=��B^�y3�(�'F{X+�����O@���&���Pf��"�C�%]E��*�%�-�t�����P��='luݻ���io Ʉ�8������!ƿD�Ҕ��/�=��3=\���k�~=DR+�-}����/'�����!���X���Q��UR���{'b���YO7�ZpϷ�J�b���/�6)u�nk��҄�"��#�CU&�H-�+�I�(-)��M��`����y�'ہt�B@i?��j�~�f�m�gt��>�p��q��[u����JɄht�J�v&��d@_��ߡ���3�5��Ƚ���n|���
6�|AAf2`�u3r����4	.;�,�@�d��/� �	�3��zQW�=_aI�J�����u�B��;��^���45�A����N�N;_��FUx4M?��z�
QM]���l| �]�T7� �BV "z�S��uQ!�F�D��U�G�=�]����B�E�g ���'�т�	�zL�Bfxr�B0 ����V���� ��~�|(��E��7ĝ����,��2b��!��[��@�V���̐���!�?�k��-Ҹ�W��yٙ��ˤ�Y�fBܯ�>W���}
���;���+}�.���d���4ź��ͷDܿ����~�Sq�[�1B����;�r�c�IEm�hP�|'�n>!'d�u���Sd"�s�_Z�� W�-�)E��{Vi�=3�xJ���{����	.��p���B�_�F��]�Qޥ�!��K��ȝ��+GH �NR3k����đw��Y������/O��]���r׺�YI�0II,m8��?���d*�������J܃�Ѽᵣ�)���j.ǟR?����5} ��–UZg�0k�_�G��N+��Bw��|�@P̨5��Ҕ�����:�\���b�6"V3��sh1�D�dϭ�kqth���	߽5��~}2`�u
J��#S�k%2*0Y������\H�ӢMHw���F�܉c�j��A�x1��P!�
�I��`�f��]���%�/1[T������w[*z�?{ڼ����'Ӹ�obKA����Y���D>g|2�c��'!i֕��A8^��!��	Zx&ى̒��8�ʾ���[�$)s%/C���\�6��@R�>cCQ�t/U��jEә]lK*|_R�=׀�
L<d� �5p,R��r��jv����o��t���	(�J�"��� x��57��T�~���O<�^Je������++W���Qɸ+!�����=|�x4.I��a-��� �|cĦ�� ��9��ߛ�--;�C��,��<1���
�C��m�DW�lb�r�u~*6kK͐/�'�1 ��|������^og>�5u>lа~��Â��a�W9Ma�������2+m�ȱ	R8��BO$oH���]�+����^�݋ª��܅�q�ρ�~�O��=T�]A_�F[ƛ�6�n�~��gR.�@�j[N�#��ѹƤ�L�a��eƸ�"d�-/��p6�h1�Ф+O�n�o�>�Dk�!i��<\���O,��r}M�zK�I��*��:L;V�1@�L�a_3�җ<x|�8֜Q���Ն�3g�?����1ol���5>�9R*`y�>��N��z1���/��;j.ò����%�����b	��w7��L�N�
���'�۞U\{���l�Ծ�cβx��;�MB�*�r�Y �SL��e��Z���� ���� ���A�@3��&�
������B_�J�|��<���×���8�9H�����6Lx�V��G��Z�2A	3���A�{ȟ��3[R~"'�eP��Q��:���]L��[Tq��	TS"��x��ҕexԟ�qZ��=K��knMy��j0옅(�c��=P%32P,l�h����9� v��	}e��y|��*�Ȱ#'�C@֕%�/�é�t����/��E\pO���S0w"k��#�%��f�b���Qt?k�^2�n��jgu�~��uބ��� �Au<�O�Vw�aj�9\�d���ܛm\N'3�=%Y���A5�e�N�r�����B��LuÒP;B�\ m��\l����(�I�Z@E��n�s��mY���1Z鷲$j�Q��H
�Èj��j�\<k���K�(���UEW�Z߶<6@$��r��E|!wc?fhT�t-|xc�Y`Nh�]�w3`5�9��@�l�=�|)���ѽ�S��R�׽�Rp��=	he���Kr�ʼz��R~���B�`�&4\z���}��%ehZm� �V�Ybu�\D)!ur��`.�d����b�t�m�,���p�^�BE߄�V+x2ڴ�#ӛ�E�򵚚f��a_r����с�j�}6o�.+��j�R��%ߘ^�������Xrwn���C��#*0���^�����4d6<����.,,���.�4�Y�B��d��1В�<�]��(y���p��	��$�D�:�t�2x���3:>Y���w"X���K��;q�ǟ>1�q��H�ʉD@��$U�±�;��3�I��)�p�L����r�j���J�~��8�l�9iH�%E�"#�%P�)p�z?��1��S^0 ��~,�-�.���5���;�m#8�
h��N�z��S8�W��Hp��0}`>
��;^6�P!M�����"�C��|M'ҳ�	?^(��y�� 1���.4jS���C�[��d��9mg,2	t!��^)����}��u]�U�<ӫP�X̃� eԉ��;tLk�:7,pLQ�ͧ"M\�O�1����ϣ���q��7Ș�u-���J�(�e��{�%:0�[�<�E�eUkc�r5��i�]����s���.�/�v8['E����I�Nj"�/����I��+��"����F&�»e1�J�(�{0�x�Chtny IJ1���#B�)������mU@�#2���^�2o,s9���>?���� 
��n��^A}��.�)q;��wsT,`f��,�݇�e���*Ӵ��FJ�ݧ #��Yt���2"<
vs��}�
�^��0�@��Dq�4	dQ�١Sj:�����M��)J����쇈�a G�b��tL
m@�.Σ�Q�����	��'f`���6���+7C�yOl���^:,�.�g*a��	�xO@�q�u����3_kQ��Lz��^<�c��oP}?�ەU�+�5�D�L:��[��:?NZd6%�J3eE�2�i(��芔���b��c�H��.�ٗ��Z
'*�SI)��
�`78.G��K��e��X^�Io�dH~=Xb�mL�5QM�l�|��-@IW0%�0H,ؓ�`� �����~X�*�`[F�b�C'�O�UEN�I
Rz������v,�W��r��qN�`p�|��@䆓���|����Rw=o������ɠ�������􍜯ۗg��XDF�>�`�O�ܮ0Щ�X�7���ʒ�}��X}���^u� �vՉC�4�Y5h�𨊁�	aG�� ��7_]~�l��jxS�vH~i���{���E}���-q�<q�l�N�F�
�"�
;�!M��3>N�CH&ɐ�X�b�D�Ǧ��6e��5~��Fy�]%�K�w�*T�v6�Xd]�z��4LXv�e�D%��E���X�ǐ��­�