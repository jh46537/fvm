��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>���;0���[��q�N/[85��1d�nޭ�!oX!�ذ��p�ޥ�4��^H��*��i�f�m����l��&�<�]\�8e�44���k�t�CЇ�+Y����^���($�?�`�\!��?>���l3�d%�	�]�_�J��^���׿G����y4����bI���Ѣ �4�L�:�,nmE��HHDJٰ��B��A/Y��́\MD{�+��<�Fb˖,�r�I �����$^�tL v�z�ڥ(������k4zV�%Vd\�l�̽��b6��C<�������2�	��ډ#�X���sYag�v	M�¥�.���9��䴘
0����m�}d������W�R�S<�V�j4I0ҙ�fd���K�]�іn��$]��z����}�7�O`��r\]1E%! ��)�)ua�(x�= :��i�(�1 �`Y�4ZK�W�ŵ����l� �����t}gp>�a�xp�Na��q~wms���w��W���YI�z四��x9Mcp7WY�bR�r%̺�*ΦW����R���������|���{���(����_��\p�N��&�#1Vx1�z��iqK]Bؒ$�Yj�=�d��	�3,��ZʁR�����>�^��$�!J-<��1�m������� $��(��~�n��<�m�Y�B��#1�PJ�.�D0 oF��NR։g5$/�6�$>Of���Q'A}HD�RY�3tVƍ[��J��l�@
�Tg�|2�Vu1�!�Ȃ��L�r*z���#�����,�gp&#�Y%F:����y��s~��)Z���*�#nnG+=�*�Qc6�0��E�E.n����ݴ4g̖�c�B��X�	�������w�\�����G,������::fq�q(������}����e�Ƌ�<.S|It��2^rŗΏ�3� ��S�7��oO����P�����pk�;��.�n��U���ԢO�B��-2-+k�X�=ly�d���0�Q٪a��\֗f�1~b�O$B�å�����f��{�I袶ķGCw&�}4�и� rxv��|u��iqo�Y�ꑢ�62�?j��e���YpY�R�4C2���q��e7�+Y���w�Q$��4	�S�D�hΓ(X]��^��O`P���c�
a�(�P�#.4T���n����E�#��h��ǃ0&���K�,B����P��C��/&��(A/�#�\� r���+$��c�~Ѡ�Kgv��(Q��􄧒��9��>���O@tKV=ΉD(X�C&�6}7��N�p��]�z���ɻB����A:�rVa*�}�>	}$�����\=p�D�(-����h�H� 5�w�����dW�k�=�J�l���@F�:Y�\x0gy���+z���6���	E��;��ܝ{s�D�|
0���F�����w���#'+8���U���~�=��K��4X�Ь�w�
h-��V�zy��\n-}<��Gh�QWU�1
�*�{&�{Z?Q��J4*;�^���jFG!-��k-��-�j�
��o���i!E���q�R�[>�e�Q�����p {y�gըt�CC�_?���6F�n��k�є�ͼ�0D+��ͷ��Pf)��l�+4ɪ�6���4Jw��XN*�X�g3DFE!������CL�3�0��0��鸉�`a'��^��b���L[��z�һ"Γ�u�=A��#PU��|��o�Gճ^^�lM��":=�v8�c6 R�P���I%��0�?�h�y�ӗh5I�3|(�U�#z�;��=�1�Q���]��� ��i����0��p%� ɷLx�"%l�H���l�<�s76�'Yg8��9�Z�řv��`�(�(�p�d�0�>N
Ʊv9)�3C���>p�i���IJ~C���t�+��icq�S׋qmX��ڇ�Eױ�.�K}�oî���d �V4kŃY��Aؐ��+��W����ڱO��.Pq��k�߻0�_�'�/�5~���h���)���7}�ɻ1��=%5�h�Go,|͖0ot�S-X:6&hӯAԾ������(�S�
��棳�X��ڢ�Cux�868�^Kj���-W8d2�b��g�.k�,z��>�̤7�8��Ԉ���߯1�37�9��A�x�q���Ex�-"-�#U���n��I��j?�|�ᓘ�(T� ���Y��w+U-�0�����w��f�����oW���Bss�>QP]�!������l���ĕ��K���z~4�)�������638c��{���V[��i�ñb,���=���Ƣ2�m��>B~��O6�Ç>x��^�ǂ;�g���u�����yh��>��Ɉ������\\���]R��_K�Z8�ƭ<(���8�s�;d��bE�w�&��"��X��,�xJ�d��8A����JE�Fÿ_��^����Ɨu�u�G`
w�p��rDn�Ν��S��dߠ0W���9����|	_Ő�;��Q9E^"������ـ^�a�ٙܣa�$��T��e��һj��B�I���,:&W��^�Y�DM�D��G{7�W2\����|�����k�x���\��~~�y��f��� �;���:�b�LQ�oQ�\�;�d��_�������픤T������n�b,�|���4���!�J~CxVPn�-1�Js�%�GxEcAiCxfj���mP M�ET�q��M�[����68��-dhi�i��K� ��c�V,k�
�Ƕ�Yt*_l�G�Ɨ�-�x�ofa�Hں�����s̸+s��˦��t���*4��i���s?^�5F�<Sn��$}�ݍ&Đ�(B!#������5��핔Z�f�#[e*�s"�����#�t�XO�韹s��J�T���s�(9-���OZ�J�*��f9nR�t����3���d���m%V[q)2I�K-s-4~l�4�7z��rTO�u��Q)�e��:WMm,�Ź(��6iGx������n��݆U1v��&l�Ǜ��\�2��\�h�g��+�a�nW�{U4yId(��AF٢�s��kck��X�x�B�O?sO���ŏ��N��J����vC`"�d:�6��%��� <�-���
ȎMN/����)Cezp�e�8�H���u�b#�dz�>+/�rp����j�s��jTg95�yJ�����\�)0�������Gm>G*J(dDo���Ks�K�A��3O���]F�2���t �ĵ��x}C��h,�z�.���W�<Us�#~b�7?+��:���mƉ�ˏ���J��gD+n]�\B�:c�3��Զ�!��$Ǟ�������
t���R�n���k�_�+��8ݾ������=�Ŕ��L��/��}����b$�|�*X`q���L����z�����Ӥ�g�`����� �6ewz$4R`#H�����7��R�x�?�F9畝�|(�g�P��T��v�-
���Bi	� ���a�*2���=��d��<}�����L��m�^�fT �y��mE�"@&���G�>	��w8��w��`���XY�l�sY�s���>-�Y!�0�;��:,�!�D輨\k����k=�\o�~�25����܈=ٝl�"�}��|@í;1��PGo�Q�>�sf~���Jj��Q�w�&<K��֗6R��"k�1!�1b��!g��3N��q�3�����D�E�8�/���i�D���Y�`Ў}+q��:2hG@��U�h4�93��{8�ܾc#�ٱ�/�n.u�F���.�}��q?��2Uݻ,xd���3��sxe��7P�$$��
�C�-u�l�:"�+�d�y����=/ �	���5�����A��Dg�[�6�')�3�1�4��^���k�L t;����p�h�Obݹ�Y-�U(�E�?ily`�e +�ް�Z�ɠ�P9dxQ>ە�}'e�`$Ove�cjŇ9ʮuUȢ�M��yӅ1�[��5P@ܖ���0�����lx{x?�+������._���>rJr5�:���Е�v��/��]AT�� ���e�t,�#�^H6��/��^�r,�j���^s�^�z����/\N�]q���}��6�	��X�t���֢	�s�e&��k�>N'�u/v�I�DTl��l����7e���=W�B���(*��o�ީy�ֲ�[��m%I{G�x�c�4�mӼi��\��Nj�Kf���O��F�	c��	�
�y�\ݼg�m>(�8>٣ZCaH��[���H��'(��jcP�)�-�L�@o�K#����Xtu�߉�!�����~Lgٙ��(�}z����ǏpG��5����gyР�Q���I��&e����	Y",�E1�#����[�W��B�N.�	�d�-�`N�R�;�:���+@�@-j	0R|�0.��Y��H�a؟иڿ".m�����X��U�	ۄ'\#�(y��l=�}�E噦[���@�4�0"�+����ߖ�K��8�b#g�@�c�0Opj�����4xn*hZ�Cy]~X��J��+������/�d�{f��k�%u�����jN���E���C�u�����!�>|@N�S1�������Ͷ�"��ݳ6��tN%�Rʅ�l��e�aB�����l�\g�j��������CKI#��XJ�o}(z5i+��F&�y��y�Oa�6T#�:�É.+G��QȊ� ))
f~����#��Sj �.�x��u[i�������}�ї�'��9������"�$�^�`Q��� th���>'[b9��8�v�!m&v��u���LdD`����B����h
���ŉ�)�<����o�䚎�i�kzk0ϣ�S�R��ߣ�14�JJM<\���#�*���]G�)���;'�,ӊ�>����J�#�p�M�wM9�y�����P���92�=#FN�*��p�A=ĭ:ц+�-�S�,<D�%���̀��E��H���<. U����qX����=�JK�l-�����ؠP�����&,ns��#�9�_�F�~,jN�s��I<H-t���\P���`�dl<O}�؛���t��r�X�/��0���D}�-�v���`�g5����!��S��5��v�a�ܷ�M�c��0[���?Rc�ȓ�h�*��)e�-��FK/�J�`�.}ztȑ�٢�;��q���i~%&�Ox~4��h���$4xm��ߦ�6T��+f�1�v�D��A�b�־�K� 0��8")>A�>�t��y�?�#CZ.����nxٕ�>zM(Б��6�A�[?�̋|�i����V�"Z�=4�e���w�^q�ޅ��th+|<�U��e�E�l�f��ȦHz$�����K��.�Y�}D%;vg��ߘ,k���M�'�Y�5��?6�Z��a�x�_i��a�<�?���д�x\�pݪ7tt牀�=?�v���Z�%ƤGg�Q�8�8Fq����!ҙ��%2ށ<ԏ$?Y3� ���Ӂ�ؚ��e�ay���y'�,ĐK7WR���Xf��`��H���_�Ū����$�(�ާpr*h[3�sJ�SIe-�Nk���l��W3aMȺb4�l�$j�VD$�?�Q�-���z6�S^n�YI$����J��`�u	��)���$Bn����q�4��&��}31g�О�<�4���-z�&��1�0�_ng����q�7s�}�9���ˣ&c�Ut�q��o��l-�p�e��l� ����깣�.Ϲ
@j�W�e��C�q��@䫜L\~�E)dq��[�$�X)d�џ1�}K �J�������gˤ�3U.�	�p|�,���Sb�k�ߑ�D���lO�S�p��@CN�a}�d�6�I�/}�3�A7��d94Z���Ѳ�����H�����,>������B^u��	���3=]B�E?1 y�yW��D����e�<�2�D@��;L�;���s��R�r�q8BR�[tb�o��Y�