��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�؆���o��9_��ʵ�Fꙣ>��IG�C�����TD��=��v��ޜ�YU�~EZ_�i��ݯ����yϋ�?'�Kъ�n�tOZ��kzA2���M8촕v�IA���}OK��퟇���\�>�����º�P�>o�QSO���!��3��0O�s�se*�}��ɩY@�js a.�۹�W@`#��ܜB���$���U�(�c`����T�[�]����ש�̊�xx�~W�u��?9���z!��`h<��O�X���׺R���ؼ�JE�>.��g�q���K����Šks�b��Rp�e�S�f�m��XEU�Nh����0��<d�R]L�t���ּu, �-E(L5�x�6�0Y�,�r���pl�Z�:��l\)$����>`Ig�yIbB��\l��));��9���_����o�_ܻk��-��8H ^����nF�P������[���TM��d�Z��� ��;1C�d2�g���5Q왊?���m�X� |�D.
n����#����@g.�7������XZj���^2�J�H2�q�Nĝ΋�RW��9�������1��g<����Ya���@���j���h��gh�m���<��X&�&�z�Sj�?֨;q���+��q�&?
R������f�0p�w-�)���ci7��F,�O,hA>�Q�֒�*�G������	�|Qjւ�𗈎�?�[�3��(�չ��W��3����\��<����=���eŪy�v��3���N/ԄK�#��R���K��2Yણv�}u�T@���<m��	��~���\B�Rٰy�5d��W��>�*qm۱֔�A=��k��?ZmL���z����ɰB��N<N,�ۜ5ş �-�6�g&UE�SP����a9��K��k*e���P�:��<��-f�))ˇ�R��� �A%/Y
��.�xa��n��$Xn�Q�[�U��o�4֚+j&�@Mq� ]�����c�ȣlS�g���\���3Pjv�e�y�$�U�9���iN����Ӟ�uH(�ƅ�?v4���@����wn\�88��G���P@��,����G62v�������ۼ��$���B��_]�OI�&�I��#,@`��q��~����[uoY��c��Z��S�D�&]�ȸ< p]�3A<���.*���?������2Ҩ�$��:�� lO��s^TG�@�*#~���N�-��4&S�?��L�_�λ�b���aӚ����:��*�f�_��'y*S�s����|�!�7�0%��R{��5A4.Φ�ya�=d���`;&'� ����������{�T޲ak�����^
�y�8�?������'KVr�� ��7�|��9��$�P�GAhg O�=��P��7���`M1]+uh�����K<�B�p�9Y������/1GF��x��	��s"��	.bA څ�?5�ǚ]�Q���7��2�:H�l,h���0��i�J�!��L�,؏���_�4(	�
C&ѽ��A"a0ϪPhxʜ�>�߱Gu�"̰&$����rpCް�m���K����C�E�rk�zZ���>>�����ADU�U���Bp��u�h����x d<m�>|z����ll̓h��(� ����� w��d���A �Fj�;;]��|�~�)�Y{g��*X�
oI�$V�\O��٤#�x��oZ���0��%�2�|Ti T�k��c!V޻O�S�F��B珜E<cZ�6�)5Ϋ�����a�7�3Af힛�Ϝ/Q�騶{��EGz�����+6�:�uJ��Ǭ���|���[�.f����!�>��q�G�QwJ?0G.k��˨�	�X:�ޝI�tl��D���_���j�����_T��`ø�^%",ڦAr��X��X����)�R�P����p:�V�\3Ty�O���ng�q-�JfF�U�����/jm��_�=bDS:]D"(|nbZ|[�9�5��Q>��~	E��`�f��ɣ�g����z���i�99����QZ:,]*�Y��*��Ѩ����}:g?�+�|8���g���@�ʍX)�����������	�� Zy N���b>�&���e������F��`S��nc�tq�Z
�:�*ND~>V�
W�%㛀�'Z�Q�CP�%2���2
�Ha�M���?�� �̄�Z
�QMv����!~���\��И��r��|�v��/�$8��e�]�_V"U���/���e��{x���b�����Ļd�x��W�Ħ�&�����B��p��Z2C��,L���߷��)V�W�]��y��9Fɹ_F�����5�2t}3��x,�?�Ne1����/���*itK:b}6%�Nǎ?
���~8&j D�0Q�A��ʷ�4��u��cl�P2���I��@�n�{z�0���rN=�jM�%'CĴ���Zy�p�Sw��cjhK��!��ڊK�����$���[D��� �/q�I��8�w����j��8eLM.f�S�5��Yc�]��l̃~h�K��ӕ"�w��5Z�s�4*�&�t�/����ߗ#b���0� *[�_��Ш�rso�v�-��V7�gƎ�)�	�@�Ra�}sN��tO	���в~���ך��t��|�n����D���e/H�6��)��l��]�K�O���ۮ��PӟQ�Bp�,�r`�w3��YXBrq�77 ��E�>� 1H���Ґ'���a�qRӥ��Q� pX������.���=��Ch��F�m�:[��XD��U�N�-&9�m�;�Z(���@]4Ʌ�5ͷ��<U�w�-���Ӊ:2:�a��l��Y$�����]���Mj�U�X�1�[M��h����a`���al��]�C@K��H� ꇷ����� �C�}��Ȉ���*)U��ncjwI"��Qx%Rs^�}싟đ\4&����N_�gr�IvK}z�� 4���έ�F���HW��(��E$�^�O�:.� �-���j�e�y���+^��K�� e���Rd��D@�VLdc/2F0���N~�vuQO���T��1�#�J򘲿��3�R�^��ɽ.9	6�q�yη�	���Ŭ�3p6`p�6�ACV�0����1mM�+�'by�kJ�-y)��D��@��b�\��;�~���@�QNp����� ,���Is `�}	Z���N���tuP��_�������3T�7�fa^C�Y0�c>U�s��,��OuW����diC3���6���)`h������5�s�%��9UP�_����PѲ��!ft��Ba��q)|�h�������k�k��׋�l�sF��d�!���eH������M�M�[C���a[5��T,�ᕰ^5�Sv���-2.p�/ "�v�Ч���خ]r������&�c�/צ��.yJ������j�7��e�X��힛:�~�8�7�b�&4#z'�9�EF�ثsM���؞��P{�r s#��81����<���Ћ�E�*k}����7�m���TZr�����ʿwJ��i��~��3��.>��۔�`X��>��0j5�������� ��_Ŗi��%�$�ʱ-��+���#�#x����#�������kUwǘ����iB��P������9����Z�N������p��]5K�	-��W��dOt8[$.�V3�������g���aUn�6XD'��̳Ŕ�a��1
��k�L9@�hCFS?�!�a���9}�9`i�\�d��-��J0�fr��&l���H��ă�miǌa1jFpX�
A�F��q0��-��i�hb��(Z>=ʾq�x���S����FsMI�:rK7��U	��)������9���5`�ӄX:��CrX�����V�`r|]�L��T�>�"r����Nwv�by����xoP񲥙�B.����>���zA����w��/ﾞR�RkC]}��Ea9,���y``N!0Z|pV}U��6�m	�T�m���]�����. �)M���z3`} �|�� �:�%$���6V�u1z4&�R;0j
V�7���RK��Dfs��S���	���@��u�n�=� L��:�y�^������g�am+��2NI�h� �ȱ��UF��N܍�+V�&���AI[)�;q���8xHn$��#X��Mi�T��&���W���"�"B�6�f���+@nCO0�|-��Mѡ#!P7F��ݧ�7��ɜ�-@X!�"DI�;A�Ss����?���ݺ����e+�g���H_���z���V��Z$�-��&<d�����

�V��C�S>5�HH؅I�t��Q��Oբ�)�$��&���.�p:���݄ߔ����'J(_LV��Cs�����r�C:!�߃	�څ�����v
M$�V����J(�%$YQ���v(��WJ)�V��S�;y�p�(�1�����O��8�<������u���и$B�$Y��r�980V�Dpᩊb3���B�_���R؃�J�-�ߑs�����4?��|�`��6W��XX��E�)�aȧc������Q@���yu�i.{}۲�����!���ӏ�l�w����������	�8qJ���
��7��u�1����4<F�l5TES�VNQ9~}-x�[y�+!�C��:���m�K|�<��&�%���&4J����fV���E�(C(q���y �X�A��k�e�MY����������|�D�f�Y�ͧTl��zU	x����Jw�XU�䃦��,\d��2��f����s��� �)��u��b鲠��[6(Y��L�m�j-�����|�_c1�ie��ƽ��9���OX�G�/>�Du�H�YO�rAZIRI����M��z/x�\+�JnT+���*m1�~����BL��$p$��( ���62\"_a톦:s�kەVD��K���O;]u�*�2K�����#���n�n��;���:��"�$�d�{������
����+t���5(/_ɠ�f����=z��<!D�}Gk~��忁h�/�Ms{"ULߢի$7N������>5_�7H�+�L��#��%"sH�lu��.uF8��G��y�Y�2�`P�/����+��o_\�����S� �g�.d�<|�ik<��#(����M�̡Ϩ̘��/Ϸxf�aix���	y��,�D���oB���&��R�4�s�"{�;'#J,��>L.��X�S�}��x���	�y���9C�_��ʣ��4�J���@�Cu���^\���@�Hi����n�5��n� ���$G�|[�"��6��k� :(��ߗ�!���θ�i��c���'��jsŻ�����R0h�
��2��J2��7x�Ϥ5�oB])�,�����'f�E7^��^�h2�i��ɛ�茯��ýE8�3�g���_��ʩ�ǎ��-�a�:^��!\#�/v5ae����A�&,��wq5����W �"6eux�Jx���9 ���[���n��?53�@K�m���p���wzM&��8w�ܵ(�'��^��O�K��<g�[����_��-���}�`j�Q��#J}���3�5B �n��Lz����6�mA��lA��j�J�h|u�CR�(�]�����0�L5�uodF�x%��^��
g