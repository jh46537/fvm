��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8��A��t��
�]W˱�ӆo �I{�C3槏��ff7 8��6���7�Y)`6�-�7,!�=�f�&Q��"�qiK���ﳑ�ɃnT:��J����""ӜJT��Ʌj����uo��]B1��IJ�P+p���Ү�r���~$̬�͇��!��||�XG�@,U���56=�t�we[�Ax��mԧ3C�d�u!�R�9У�X�c�m<>$y��l]�
�tf�?�� ^��fdT<�n���r��s�?��Z*�����)��Y����:�v���c��0�`X���}m�z0\)	�/O��Q�J�rV�SK���&�v�!n!	�!��z|�M�%.�.�\��R���Y�q��CN�`"$�T���9�w{��˙�������m�![�Xxug�i/�~����ʠ���t�s<<��3�54s<���\0ΗT����a��	�ֿp'�����v�Fd ^��g���w<�-��}`������ �	پ1�F	���l���4=Lf}����ɺ&x�,h��hZ	P�9s�r�'@m���d.�%Z���t\%��6����T�C�i���yU,�:FJE �n�-#U�+�IS98��x�
����5tgޢ��VL��`>A�	$��;,����ԓ�|��<�!p��Wp�3�EW�a@�J�uJ�����L���<v?����n	S;�MՁ�z�x�Nf���X�=�X�Mlq��+=~����N��ϖ �>�u���3�����q��&�_��Omh�E`�I*��sd#��3K�T�2K��h|a,	��},VE���;���������/k�� 0��@���E�����G`�-5~�9��"��)z��6����Ȉ��ڡ��|��A�#K�H�)���%έm�8�Ӓk��#��\6�[9�W�cLt�e�LF��q�L��
y)2�F�9F��n���'�24u�`�~a�ߗȽ�*�p�+��ө���T��*���|��+]�K�xXo�f(��l��L��I%�D~b�h)��E��7}����T�dL�c.��A~��҂>��4�Y�չW���<%q���Y�2Q�`����ЎX��Ic�f�"m���PA<mV=���<�}b1ϥ�:� VJ'�z�ɮ��]�'�<�����X\���ơ+� ���L@�l}c1�]��#�~2�9ƻt�;����4�=(0�տ�؀�ܙ��8 xy;�����0�Y��q�om��#0���q�Js�pUkGp�U��0�[��S�g jN}�ӶK�������=h#|
�M�s��%���Dtq����b���es��b��J���ѿ�'II�sro����1����{�����S�k����b֛�u�"N�������̎2�9��'���B~�I8��^�>� zt��AH�!��A+=���8c��͢����@~�{ ���%��� F�!,:�z��,�-�0Up�8�����Pk�Y	A��\yv�O�xd������ퟘ�� ��`d��Տ�k���ݻ�aI.���S��"����t�`n�xa���)<�!���} �^*h��J���B�3�<<�`Џwv]��E:�����9�*)���&��������L�_V�����ń+����7�lbz�n��"�`z���qX����4%��y�2���!V3��aH���8U)�$4m�Sß���\�X��5������	��5�IFԙ���A�e�ڸ3FB��IJ. �`�ܙ�~�B�&��Mo���p�ǀ�,���&s�ʵ���w�y�Y����D�Ii��L.��X+�>z@>y)��$�µ�&N��Z�5�����J���M����x�=�Y��w�)b��8.qQ/���DP��ۿ�Nz&�	�%m����}?$*E��)Wqt�{G���.2��m#T�-�7��X�IطK��lM'����^�+nqݸ�PO���.P}#b6K^�&�88Μ�����&�V8ΡP�h[h:Js��^KZ�Y�A�2�BD�n�`�_�T���W���2��v1�,_���7�9��Dk�W��fN��%��&l>g�����նo��'�i���F�Z��p�$4U�s�L#��Ntv/_h��58��ke��?��Q�'G�k(ږ�7�Y^yĆ<|Bb{����!�a?>A�5'�z�n�ny�ā�qӣ�n7`΍L`���\Rs6�����:�SnL棍N�cd6k4�n�cz�PAP��n���&P�zRXO����0�_0L_b�����G�L�h-��.�����#��k���vP
�$��fN<��č\تaN�ʥg�^i;�I�J+M��=��#��]�~|
�d��q"uHL�����<�-Tq��9
�,���2�>�s}��ԭUE��l�?V�Vv`��]�]�z��8�����̂xوX`��,2ƽ�E�+�G3wڀ-�n�hZ~�,��j�s>�����ƙ�ה�C�� ��[]l�_���3�v�w�:�M�W���&��6��z�.�jm���faY����t���f�K�cl�t�W���^�{9��X�����e�t���2����s�$��M�^}y��Ɇ�yM�Ԙw���+9|'G��݃e:؉�1�0�%kL��9#D�]@��v�kV:J&�YT��ۇ!���� ,q M�F��=������@���ܟ�E�fU����n�>(� ~�O��$�vvH��k��Y��_W3c��WwO���Р*E�pj��!��EZ���<����(}u�T�)ݛ*�~\؋x�O1ax�M3߀l������1M�m/�6��>.���?}���2H7���x e!���hs+�od�/U� ������~��Q��M��s����Xy��a+=�vw�^��Қ�@�� ����J3 �):x�c,Et4��G��M��
����{T;����=�E��/<&6&"
��Q�$�~&��0'���f���-�姒y9e�+��h9ؤ�a��a�u�
�v�W����:-?%ÿ��I�.G'�nè��L>wt=̔���c����jw#d{��&t��j�����tM�}�{��3��0'�9���dh����e���ġP��.Rﲹ��j,jiD�ܙR��]pϸ=p턏�$;�u���-T�8seW��^Y}�|�4j���X�;�uF��ʡ7Ҟ�)s��\8����k�i��#�?7�5��A�7����"��0o��$��Cheup�I�ؚ#� ����0��)z�d�%�����B^T_���u�˘��T��}0���y��F��>`�v�67���&R�'���S}S�C>ڟJM^Ճ�5v8 ����G���3{�G�$D���;��Ș�%�~Nrl��{#3c�9�c����P�㐤uމ�Y�����^c7���T�Q�M0�������=�f#�W l����A5
L}�t�QF�d�u*qwd���!I>������2��q�d��x;6Y�==��֒�	/fj*�����ͧ c���Hu��%М��f���kƑg�K�fMQ�-�4Q��������@��us�]�~�R��h��´�VD�n�c{���ח03��V�Rr�f3�	
a�:���]�o#�.�����4?�t�Z��Rp� hW;}��%���{�:��,�����e���0�!���u�X���������z���	�)J�$�+ȓ����4uzor�('���K	|��)73e�Ƭ���i�j5��,��e�׺z��d��@��y��)ט3v�Lkc4`夽�gjT�������/Gm}�sO�M*^�m��yo��Y.WQ��}��% �R7̥��#V�d�l�KE��E0*,�@��F��U��*��O�H��4�=AJ��!s[dU��ۜ)��C��߼��������\���P�2� $-��pg��V:�f7�BCS� D9n^�c�6�J�X�J�ISd�a*�w������I��KR��a�1��ݏCCozr�c�0'HHҧ�bI��|�h�8n{�V����@���]yR�\w�Ⱦw7z�5�b���w��/
W�oI��{Y���aW���Ov.�� �0��B�32�.��aʝ��E�|BE�i]����u�6�̓������i������ۚ�ߡ,��k��#�ː����Y���h� ��%��<r��{8穓�4�%[��'^�G^$�Kק{�X��w��wa�E� ^#�W�QK�H��1����Gk��!��n���,)�YS2�ސ%�}z[SQ��h���T��o�i�ȥ'�U5�$b-�6B�p���.GK�����B����5=�{)r�D}F�����c�GQ���S�ۼ�3*h0��I�~:-��*�����{��q2j\r�LO��3_�A��}��F�f���,]Yd=�����a��[�`��ɗ�U5R(����A=��F��n��(�6-T����i)�ވ�޶(�a� 4�?m��36��Ex~��`I$Z��SF>��j���g�0m;���(��T��0Ck����ݕ��Ӿ!A��fM˲�7F,�%�n���0�g�.����jG�Jb!�Fu0}R��ܕ��Y�KC	�����V����=����i`�SkX�]dg3�?�Q�<?�]�NT�N6����U���A�z}�\��"w��xu@l��}��;��� }��ǽiPu>��E����������o(U���Y��p� �1&׶l��.�%vAp����7����kW�@4���n���)a[��Ϥ����`�z�_5�F �S����_����>Z��XV*i`Z�Ekg�3BoC�=�ޝPcS���1%�*nZ��6�����e!�|�3x�1�7�v����48~�N���w�
/24oM\v3Zz�i�1G�S`#����&d8��0�I�U�/]tt�ja��1/�_�⣇�l��( ���۞��_2��Җ�<J�2��K;�����h������d���yԪ�
�0:�N�`��2�XTS��>��������o��jKъ���Kr �ql��jD>�d��s���:����_w��a��֎��/	�{��i����#	#�N�E��Z$ӈ7[�K_�Ɵ�[��=�a�4c��G�O,ػsR�pi�큒�҄W�Ko���$	Ć_!�f�<ÈTY���e	���yE���	�ѭ��k�"��Ͷ���HKZ�݁��J|c	�nT"��I5��#/��"i5M$$4��l�匁�%ʅ.�*4lk;u�D����X��=��V��Ǉ��5>�B�X�)<�L= n5���I��e֑B�!+B�xq6-H�>^e��z�G:��W)0x��_I�e�;�9U�Q�Qh[�ȫ����*�Mؿ/�4M ��%d�X_ tS��?�Ѧ�әH�a���e6Yn�Foo�9�)�#=�S�A�wXnV�e�z�_b"��I�Ԭf��6����g����@�\��w'�e�XzE��2 j��G�
E����D�����͍pX䋔���F^�i�qC���0�j��@��ߧ�8�)�&����S^TR0 �NȌZl�UG�iD�'��\���N��OR�5��4�[RO	|/�O,�Ɠ���6��
c�]a.*2o���^6��z��&8�A�s�C;I�o~��"�I��o�������}}4�Х��ן) �Y�B���m_�D�-XvB�B�����e�"��������XDT�p����Ҿ����V����'N����*����,�x.^T9��Z-?<\\���iwV�Qprc���_"w��N2W�h�K�佽⃿�>�)��UB�*���h�[���x*�j9uXSfԫ黹�%+yuN�6����f���,�ѻ��ވK�`A�=�|#}�xO@KJ0m;�1|я����[ߙū����w	*��E�|7�x��l��4\�;��� Jgk��̫�S�R��N_jV���H�]���۫ȋCm�r�Y	����4�N�ܨ���[N�������xn%zM���@��u��!��hj�o�Ҳ� �^k�_n�f���2~���/�[�]	1��q�ܾ"��HC�IgG!k5��N��`/��^�;rfz ��� K��Ō51?�z�
�!C�E��FѲ$�_7A�L,2*��:���9�w{������
.��W����k�@�C��q�R,�u�m@d����n�L ������^�����s^]��m�(O�~�V)x?:��5�,#�%6� c�֘T�X��#br9�����5^��P���Ab�p�Q솥vk��.J�(p���Y7ˏ�I��ͯq�9���ם�����*�6@D���|���11Ȁ̉y2 �ce��O&[7�K袨�>+��`��Q��BTMi�DZֿx��UL����Y~N:K�F�
�(��m 
��ʼ�Q8����ğ�fu��i,?��c�v��+wQ�b����RT�~-��v㇭���de�5h r�qu��~�g\t��LN��߉Ap�H��b���n��ڈ�x\�h@�Δ'P)�����-����Y:�1U�r5%�`�~��l6��*<���4f���7���ɸ#ڰ]7R�a���X���0�_�� !�GI���/Zp� ��潘�%l>���Y�0����h�g����n!��9tS�����_�{��9���1����?��n4>|>6r�HA3��A2�i!:Z����k �~|7Q�Ox���BƉ�Z��nAGoN��J�����GԞ�*2N�03���_a����ڔ��T:�lo�A�g;|T�/p�������\����$,���5+9�����z�$�k��ۭ����}%z��I�N�Z���F��Ń�r��[�Y��e�^a�5GL�����5�t��p �
�f�aΥ־��8S�=a�m]��r�\�{�K��~�`��Lf��1t�� �~�fOW��uz�?�zi�4�
r��!�-e�e�)?��d[)'ԑZnL/��X\��4�35�,g�����	��+v�68Y�嫀a>-��p�%��������i���'ۦ�1��^0F�E�{x�-]��:Z�zj|�f��]�Ai89������'�"һ<�ɦ���|@�Yf�{b@t�v�1͵��l�����k���lY���*��P�r]�u}ž��A�M �"5pݖ����鯱d7�֨Vi/��*Zߛ��{"t2T��y��v� E�����G(>�V؍���
���C�W�kl -pL1�
���Z�F���D�軋�xl���Q�.����i)U`��B���=��0=1���<�_����RWsp;����3��|-)�2�O;�0�e$/�x���-����:��{��J���M�������)	���ݡ892���AJ­��B�q�����e/��ď�ga�R��Khql<զ�gq#�\�y�Z��}l�E�?�C���JNh����ˎ� ����[S=ߥci#NI���0U�����uЖ�sU#6�Bj>���P>T��:�%m�G΋�-����WS�]^e3"�*2\���4�.� �1*��H�$�{Ѣ���U2�?�3��@F�/ϫ���r��¿�&C�~H9ڧ8���E~�"J%缇XU�V��-[��N=QS d�^uQÃ��	(K%ww����T��Ay��z[�lH_�m�?�R�д�G�3�N0�֞moU��{ �w��lc㣕�Ai[^����F��HR��f��H� �S&�y^�R�����'ܿv�,}3� Jh��p�Z�r`��<<�f{`��}�ꈱ�;?�#���A�k5G���ō�/N�Y�S��p���d��*K��[[Z�1��zO���
����w�H[���̓����Y�Fa���?	�.�F�m��k���WI��t����(wk*"�2�� {���kߧ�&Q[�b�ab��˒VM�:��h;�T]`ѕ%��|�<�l�1�c�M�#���h會�۠�B`����y�����m��@6��:�K�OqѬ�a�*u=W��<�̓��1}����Xv5Gq�4?r'^���״9x��:G�2:�d����0!�A#o��^o�n}���"8r�@s�]2$s��$GP��@u�*��M{(�M��N�x_kU�<U͡����$3Y%l��mx�#\��B�����n(㳻}�.�l5���}u����fd���m,���M��io�b�N=�kq:������~�'5��`�� 帧�칍�M\���_?X���uYjf����b�d JM�7�*��T�!G�������@Q�J������q`����W��������Ę��I�t�<��]^�U�흥� X�c���,"�W�'�uV�Y�)0�+���B۝#]� D�|�2Z�(RH0_!Z8��������3���0�SO��K8���P�J�P{���q&V���;���� ��!�2���R��"��o���RF?����I�^77�^�u2C�-bҹ+��i�_h��:�CR�;(���:ѹ���Xd�'7�/]Ҝ�����#��`��O�s>����B���W�0��E���[����Ρ��&�����a�ɢ�8���ؘ|<Yx�Y�	�HPͭ+��Zj�uo�`��!�%�+����Q��f�٪�85Ì.���ϰ �����[F&\&�*��H~�8�Q(�|ޜT[�7��7)K�����EqcT��QDg^���8V��J�V<Q\@jl�/Ѩ�$K^l�p����([إAW����d��?0K�+�)}�C$Ӷw������Q�o�����7��RR�'7M)�+ȕ�lg�?֫X�w}�?�b�
�C�WD�$��5"����V?bc�ss���h��rl����d�l�?@I�S/������`Ow�B���2�NK��Ѹۨq��I9�׉��BX�4���rI�������u��YP�Ϊb�_�m��<ƣ�O*J��ꋣM���D��d�e�����%��M�DM��zQs?E�t�+�ָ}9a'���NE��A2��eH���9 ��> ,=�X��(�el4�{ ��k��vj�F�7�ڨ\QQ�qL�b�N��S�D���IKMԶ[t[Fi֧~��_�\l^Ř�`.iZ��o�$qp�X{~j�0����i����h�QU�+�>>���~��ܫ�����������i ��+|9k�V'���a�c$dQ������)�_��-��cv7��ASW�d�lJ�D�go�z��3�u��/�c�5���K��u0�PN\�������k���sT���r��j�Q/;!N@����^]B7�G�%���cL��y�}�V�K��M�D�֝����v��T֜T������������y�{�=&����y�a>�F,"��&�@<.e�f��\�!E �;;��u�߁0�Ȑ��Q@�i�^�@��O�o��4�/�h��̎�� �)�����R������(��l�aV|^���e~��4Y���@a�[��k8x.���9���}:��|X栣fͩ�U=�?z��*X�G�W'��cR�
ً5���CQ`��=
�G�zͩ��_�qw#<���`�sh!,գt�L��؂WQv����|@N&�:J�s�H����@A ����ñ�M?��;;Ay:y��f>l�glV|��""������ތ����� �Gұf��&�aJb+��Z����B=�Gf���b7�3n���)��hdmwP��� ��P���䷩!B G�g}�4��&�P�����k���J��_\{<�w�1z�t�3��$���:�b�Ub%��a�Ô�]Պ/����b/�O�)�^3�Ȱ��L����"dz��i+>*�䧝R&�£�?NWr�:7@hQ0�Yu� ��D8#t��9�I�{bE	��,M����((r��!'�2����ʊ���&�s6�Yi��B������$f�q𻣆Ȟ�m��P>p~���<�6eh]������"�S�G�f���su:�^4酋�6��z�k���J��U����Fٶ�)LT�BT�_G�!�o"��=@t!�
�p0��)����=�6�l>ܮ=I*���1���"8�4/�t@^Z�T�!'ϲ�)-���}9xm��Qrtj��>�d>#&m��,��Y���	��m�'S�f��y�-�	�śp����?;]����_*���t���3�m?}m�(8���i��vU�&�~��)\��"���5"�@�T.�nn�w����<I��<�'rSt�T�י~0�%����6L�����"ꆕ�('trL�����VJ+��歅����'���� �I�D�lG����a	T���s�����iS��� �d�l�>�0�Y�/^+���E�&3�Re���p��Gvq�kn���}�pl��o��ޞ��TF�R�#�I��jTķ!�+��Ia6a��b0q5�nJ�#sa�f�����?F"6�t��%�@��s�0��A�
���cϴH���B���&�"(�y-?H����P�j���� JEk��
����-��k囧��� `ܻ�* ��r�M��l�*�F�l�(T��Y@�v�~dQ���#��R�Up�;x�$Ξ
\��Y@����]��k�ճԽ
�$F�'�M4d��j� �o�������61�+��J�YfLC�&�!�C�����#;�p{����/���g��"Y\:����}�zD���C��������ס��刻�qw�ͯ\ѯ)$p�`���4���/���=ʹ�u0H.\���!��b�<L	��\����X�M��r'~�)�3��pbW�}1����l���M*t��|kg�)��SH�9[\ڋL�uS��Å)����s�tx��*�X��6�)��]�.�fiC�K k����L��	ƛ[�G��{�bˬ��<%k���z�T�;5�Y3M~m�����ط{?�<���/x5���a�E�� ��>+ߐ=�wa�F��ME���Yr��?��?��}�1[�t ��bX
�!�3�(�C!Wxx8���k�1~a��˘}�t�B������? ��ԻI��a���8}��/ ��]2ce��r��#KQ��t��[��)͎�!:����y[�6̩�:�,W�r�p�owC!�O�-g�,�HF����'F��)3���i��P6��!��@\
'Yyna�]=!��)Ѿ�@�=�Q��,ji�o8��cx7�΍5��ǘ���'��RҞm95B�'�{�0n�@ ��p���Зɤm�e�7����$�I���	�i�X��ۼ9e��X@�����L�*�և7WSO@�P�thD"�Qq��$m� �-	�@�$� n޺�7:�vQ� �m�[7z��vARa��4�@�C�_?�őq;���Ow�ZQ��]!�Q�٤����Q������J	Rz)}���AJc�È�|�k��x'�=��ܩ$O	��G4%�Mw�#?#��|��1r�Am�]=A�Z?Q��.�l�Z}V�[0��Զ=}nv)�T���v.V�lM�!x���D���c�`�lQ�wrdb�ښ�I@&�L+gr��s/X���[�d�p�΢���TKE�t�x�@��.�m���o!#��f5�������ԫZ��#��G�[��>����^h� 7D~tn���H47w�F�	���3�'f����{��b�>���ރO���UGD0X7tߘ����>�����9f��z�^�̒$��@A"W\�pU��T��N(ө��s"�d[�t �R,�:�nd�!���(�Y}FUq=����\���h���Xv�0e�P�Y�g#�;/\�W'I%��6���
�@;��[O|1�+�jp�q#���tx�{�V���f��܀֪�cS�� ���&h����s��T�Z���D��&&��|A�B�\ZʣᎪ��5MEϳ��������	%5y_Ჲ����R�"���K��sH(�&�0�t��[>��w~���hmdC�M3h\�|�����
njwJ X��>��J`_���� �$�X�^��̞3�*�t�h;I��9�O=���9u��p�ޝ_w
P�_B:�r���o&|���u���2���6���g�1�Ĭ?5]���6t�+K{�ɵ�$8$V^t�t��������i>�|k�M6��l�GǹZ;���"�������v�x3kb7'�2��i�]�X��k��`�QUF;��঺�0��k�cE��갷>��N��Sj�Cx��t*�]R��4��/�V��=�M*ì9V�eL�B}k�1ۨz�$?�SV�����S��F�&]!�0�) �}<��Tz�c$1H��z��P�
COm*cY���AKF�ьx�PQ�,��2	��Q�?0)t�s�z�ō;w�8��$�y+�"y *���"�ˮ*1\xj>Y_�z,�h���O� _2��y~�0�B����o�%ɧ�Z���j��K>���F�h��h���+D[L+_��LL_��֣����k�U�`е��F������{ϡ�x]0M��hu��̳�8	�=�T39[��5o��O����p�~���7�g�'�k��аʬ�\���n��$��艽C�ψv������eTe�;�C��1726]#A�����c��z��[�{f~��`��='B�%!-н���7�{3Li���^�����_�h>���YZƞ)k�WF��Dpv�p�0��/�ɒQ�� A!1KL��L3�����=��P���$='&.�85ֽv>��N�]Jb���/+ Zze7Ҙ���wպ�"�F�9R���GBj�FY��V�oص&��1��z��ܧ��(�:�${-�heـ�V�,�w!�*:"xG�&����N��A�v8v��s� s8�#�� -��\����R�N��i�{�>�1
�7�Vx�P_��CNkhӃ�� 5z�*�?�4���N���/��֟�l��r��|�RZ��&b��e��Z Gz�p�A[�2Mv�>����T�'̸�ª�6_�^�%�����#��u����^���-���x�(���K\��Z5��em�ͻ�=*�x�a��vr�N|�t	��S.a�nyc)�J��bv���AnG�����s7�؉��q��^+�����f`+��p��?!s+��>�-ikm�h��O��MP�}���>r���p�K�~l�}'���:�_�_�tk @\����#_?��`Ŵ ����'ԩ�R�@��������&VoK�d<�KE_�yФ�٘����,�n�T��yc������}O��c����AC*�����.4s�M��?�K��m�}�_�Wʖ�)�b���u��ز5ѫj����Xı��!b$��+�U�"�,���Ad��K/�M�ޣ3����BIsO� ɺ��5?1I��Vl�d�n�8�3V�n�,m���+Ѣ�)�Z���8���y��a��k�i\s%}b؄�\�)����+[�Ë�E�/k�J�(�z��%K��{`�M=�F'l(� ���p��E�����<=�Z�I��{W�|L��]#|Nj�I�R~7�	��ɵ�%�(S����%/�����ڸ��|�i�`\CX^p��0�出�"����y��J��''ڳY	Ձ��Jy�/�ב(��,$��/��9�=�`+>�P�3�O������+���
�#̽QS묊TqO��n~��R�N��J�6>�e��%�r!�8�R�����K�9��d�ӫ��r�t%g�G�' �hX�o�|D3�X�BMT�KQ]2��wa�柟��e�vy�K��*���Ǯ����d�af*�b@qL�Hɡ
2�V�#�<K��1E�C���$�svD��
|�"�zm���lVy�4�����qY�g̑"���e.����-��E9�^��D�T��@�S�Ŧ��n<���c�dVbA����\n�i�/��%c�����-HY�1m ��h����c� ���в14{�De�3�y4��С��c��������,6|1ؙL���xbZR����A�Lφ���%��g����fh{�l�����6]??bz����B<��f���L�������~(M�C1 u,{8KH���^đ2T���^K+ڸ1���%o�H���MjuE?7��l���f���gi�)��"a�� �dx�;њj*k�G��5|��mq���|�Zp���+�C���gQ����-�*`�b2��5����K1o���Kؾ�\���Ux�Z���^d�VT#˵`��|L����mcXGjB9B���yY8�15k���FBH9�M��� ��jRg�#]�%c��7