��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���D�w
��p��������Yx�;a��>��H"���z�'��!� ��������	z�D��>ܱp�H�����7�8@�e,*�y�wP��6@���e<B,�����p#����W}/d�q��+VV9�,;%�gǥ��g��j|�}M6�$�������Qg����h�%`u�H�'�Y��8�8�?�yU[ �Y�a��r�1�Ѱ��|2�.�z�<d]uc���V�Z����<��z��亳�I��j�]�x9�f�4�w���8U��r-��b�x�ȥ	w�a��DY�c��:���ir:�g��S7�pP��Ƒ���w����� ��x�i]�cΟBy��$�>��T�s�`}z��I���C�`Iĥ +}����%ώ�F[@��ͬ�lv�D������g�ҋ,9�����P�/�55%q�s�T���MƄ_�<@H��-���t���x{��>��p�6�CA��|���h������\��5p�Tp�D�y�V�G�RP8������J��V�f�� 0�z�c`��9���|%Q
Q��J�#󊡅�Z�tKr~��S�0��h���v��˼+�A}�#�� �)������.�Y���0��\��9ɫA�W�g;�n�H�O��o��:�!m�B��4��b�Υ�Y�C~��qF�O&e�"p�m�.�6?4��JC�9Lђ���qt�p�V�����	F%�:r`��a�ߌ��q�x-yF�M�.�5N*#��8���'$ܐ��7&�e���!D%2��R���X��@U���>HQ�WYn��"�1G��Ҁ2�%F���(rx�!tx#�g���
���������S��{ I�oAR��.zA�*��FQ/��8;�%G�J������ �i�;�p�����X����M��!.o�1�K^q>��S#q-z�Ϗy>5�Zr,a!;�������d�7���eK8�������T��ݣH2:n0m��jy*�a!���A�=����M0p�_MN�ZH-؄p->���'JhBr{�iYhXv$�S�7s�,�+{�q�3A}�`�i�|ωo��'�2���F�cڊ���=����ְp�M�����1�ޱ�5���z�Qˀ9t��9<"���lą��;z�_��]Aݷ���F@��o6�G��5'm�A_��k7�̕Ɔ�U`��(�b��CC,[�"����/{�_�Nf��G:,^��Dr��:ڢ��?=e:ɜq]�����`$��ÄFy����4*9&���E��8�H��,��?��د��/�<U��BY�5`.���,��ɍ~�+�Y���t��x���NϜĺ�1�[�xw�Co�jQ2�7�V�e=�(�C�$K��x�I}�mL��k��3����R�0r^l	Y�D%�cQ��Q����4J�؁b���]�W)�7�7N�l)t��"4,������.��<t���EF1�`,S���zk[�q9��pOP��r�!<Drrr��cFG=�-�8&!�\ۖ��^���%��|����??�`)<��C�%	��їB���V�`�n��p:��=�y�%;��u[5�������FR�\I���X���uri�N���i�O��:57�}��F�}%�_nM�������um"��:����,�k �U.G�~���*�`��f�᝛.447���i(
�R�o^g0����DpQ����I9?�b����Wa��}y�(D�abۻ�I.��bwH/��,[ (LVm-8C��X������,���-������>���OO�!�`�/k��z���A�vÙ0�����ZF�ό�y�0���}#�.:�h
���n�%R�ط������G2~㾽�~�L��O=;aNE�/��t�r��ҕ�.�@Ȯ�ɞ����s�M@Σ =�9_��wȟ�T:�1�v���sc��c���zb��'y7�g֔���U&B��oĳ~&]��cr�%�ǌ��-E$�ES*m���Ⱦ����j5+�AحZ��wu�+e}R���zp�Dچm�'+o*^����#!����wTq�������4�@U�եrp�L��dg��H�nI�GW\�`�Z�=ʦ�:[nb���00�	��m�^Zi��{&�Gl�����&�e$�pbZ��}�v�P�U�i�ſ��q�w��K������������L�"L��Y�;f����34�P�ViZ�p�T.�U-��h���i�&����T�e���B�eZ��Lkȅ���L��.�o����rw�`�&_S/G�?7�
?`lkp.���0���&8T�7�_C��L�ǢPD���Jq���p�x>F���K��	�j ��0��ݍe�1/�f5}��� '�g�"
����������ݺBG�`Ȃ|ZQ�Q��DZ0/uI7��Aek��|-ܶZ��Q�2n���_w�; ��"�SF^U��,�͒S�;i�ʟ���-!����	�_��%�sd�\oU����J�����r�g�*">�J���j�ݹ�����-���識�-����)��
��鳇T��wOa�_��?3#򔡊��kW�'�~���(���Ʀ��!���%#r��,3���{���c�H9��_�
���!�zql�.
��[��Y`c����������\̐���>Q%2�s&<{Vy+b"I]���8WyĭBoe�����h�܏�d�%�� ��Tq�������Ea��'h&�t���J�� ׊�O�%�6����[�e�DPf����l5�?օ�{!FĻ���A�Ǹ?�E�=��|�wo��M:P!d{6s�OlR�\�_n��ܻ�~H�O� ��9���0�V�Ʀ0��브y?�Wh} �gm�j���9x�P�?��HA����.�{줊���S��w�8�3�Q\W@́����:���8vNʶP�(��dG��ݿNR�;��ѐ\�E�����w:�����s"���Q�*��v0�=��ro��ʅ�_�(y2�ofN�Ѥ+�z�U���~�'*:��il��r�v"�Z�9������vR��� �Sz��$Uf���g�hGbF��/c�1"�$�� ģ�c#��&�C ����W��%�����ϱ���I���AE���#�p����V��Id�X�ȤLE5q�v�K����;7_���"�˱2��Hc~4���=iK3X'�H�O�b '��KV��8�tE�Cx�*�%e5E�� S��>�;#�Q��nVt� ��FV�!��d&�c��'��H<��D�{X!�y`�������az���C���}¥����BC��m�t-���V�S�]6�盡���5�?�P�:]T*E	��=��ϡ�r��(��w�l��f��e�Ŧ���J�Ig�p@�m��cgw��	���4W��;���|E�D��}W����M�DW�T'I�.�W�]d���/�a P/��3����kЏ��#A�nB��?�(=,!c�����?n��.�Ư�!q�0�4M�~>/ē%�։i�og��F�)qY���D�դ�'+ �v~�%��R��Ca��
��j�&����J8���ŷ�a�a2wT�=����X��@^��^�-���?�@��x��S:�>����~ݗ�<T�]ڸ~aü>��gzzA�Ξ���ϔ�a��D����Op��m׀�} I��I�t�Ǿ;�H��) 2,2	f�,�Cl�"���5[>�>~۔roP^�Q��`�}�ar1����S=ۑѥ���!̢� �'�q.=���MX�B�/�k�wK��36��N&3��S�������Y�����F���in�pNC�w@j`�� [��x��(�
OVh Z=1Y��[���7@�,SԻ5��FXc��"�%N�E�l9��E? ���g/'_�`LR83��1p>��ֆ¶����D�/�>A����Ώt*�/{�Ҝ�=�m�6rO�#�����y��c��2T�q\ku���k�g��+wu���W�9�/��̍��h2dSs'��8�)���}����*�:gj�M��P1���is�/E�I�{#A3~�,[4}
!-�%F���b��1�I�h�8U->"Wq5�����Z&�~��h��Ћ�y�L����\��������Cۑ�®f����W~��B�V���Q�a6�&Up=-5[�SP��Nx�Z_^&�[�k���9��k��L�e��Qm��b_r=}O��)@y޾ζh8����UOg'�枪�0�e� �HM��f$/!z����сs�C�f�T#�����W�q��^�'uf�J!J&��^�[&mpȉ3C����Eht!b|�z�[5U���Z��+��լk�[�|5+��d��rgb���٩s:&����5{��L���r<!*Rʵ7t1��{BᆛΌA��*Ͼe��B�7O�/F�ɘ��3��i���J�lU�G�L:�U����{�m�6�&Q$;����;�J���G�����m��9O^��C�gQ�[����I�E�����cH�� {��ɕ�#��٧�M�zy��zuv44%�����F�y/�5��4\pQ�bs�s�F�����/mGt!��=�7,�?	B��; ������V+�7��$���������C�/�O���^��̎�L��!��&f��d�X8\���6�t
O+�{�D������Az�< Fv⌒�Nl1���՜����v�8�o�[��О��2�I_�/C�n�>�o�C�\��*��b>�Q)�UB䧠�T���:�BY��DF���@ J=%}�0u�UÏx�H�aF~@z�TcU��f.'��55�lMw����H��0�b��l�32��jpW��w���K�w�X��EBi�u�^j7��Ba�Lۣ@�d٪��ܘ��[��n��\��j[���O��u��^v����Ꝛ!]��V:��<\�Ct������u��kx�� @�&v���#ZF����B�<���y�[��������񾡳�'P��<�>l�#u�Ң�|Q.�&��Y���l;a�Dp?W0�\��U���ݹCc�' �;��hz`T���ߙr���|�wăȍG�L����wi����H\���Z��]N�|_BCG���֯gCz�d��Z4�t��Tj�B�"��v[�yI�ȓȖt��2Fwv�!ET�nE��T��
f��%���˦#��Ʋ�U���V(�q���a����f�#�9\�J��֝H�'�m���/ۑ���m~�%��ۢ�߀4��A��CO��f�E�$cʰ������$3�	(��&����x���]�H��.&q��AdE{e*ۍ�&�oJ��/e�n������5�O��O��S7�4�P]�%`������h��p�9�Zz 7�*{�J��I���q���J�RE9����)zO��pM�=z������Fz�V��[F�:�z � R���Bxg��z�3k}���U&�#�m91�kVȎn�nW�p�Y�>��
/�esc?���.�<y����Q�Ԛ�k?����N����3��\�U��Y���@6ǪK����(V
#̗��b���:�VR����Ԗ�>3�O M��7�%��C���$��Y���Z�Z&���&` ����c-Ã���_���T#	��x�V�z.<t�S��=�#�D�r\;E+xv�F����0)���YK������C�%O�\[�pCp��k�!q�@O���ʨ�H1��'�o�Z�|;X)�,'1X
?J����H�2 ����{ſ��VBV���@�Mwv�'���6�y�i?s��ف���R}����P�P�$=N�7��G�8��Z�
�`G'��]�^�!��;L�D�鐶�D��9��2j��.�v�C�0�k�mj���,
��[{��oȾ��T����)��\)wj�0 �'����YJ��l�� ���u�R�7�ZxD�`�Y�-��)��d��&�#���nd���= ��P�Zr�P�Y���I����W)8�Q�)� |�'�7�%uH��������i!�W���#����q��k�C�T���\�*�.4V��p��55���H���-���q�lK�G�B���x�,���?20; #	P��a|��"���1�F�?�y<~r>ڎSZK3j��Iy�q�g�ǲҨ�v�{������Đˉ:m�=��Z�.�����gn���1�3���0 dBS�uSĪ b�Q��&�y
1A��X��-k@\2��"� n �yu�=�fH�h��������������a�Q6�~�	x�g�b1��Cǟ�Tn!y{<��C���q�h9��B�s�j	[�#ԝTx/l]��VU��	*�{ѵ�'S�b��`��&�z��uy�Hj�p��39����\'���b�����R"������c���-�
�o�w�9�c�"����p�apC�	��\$��s�b6P��z�\�U��ql�k^fP���SCá�?�������Z��'���t鋑������Py�4��"t=��	v62��i����UY���c�%Ҵ�P�ۉ~�˳Q�[��Zx	mT�����cOGo ��P@��`j����R�0o�Ǘ�#�7񰜩W�D<H���v१ز�S�J�����r���.����o�*�A�"1��J')��8��ۅ��cLjC1��QO0�1�o��U��=?<:Gi5)y+B_�k�/̇���"�0!�����AkzA����"pZ9Ę�\>���)�ѹ_O��y#�����
HAx�>}�no�<���ar����%�w��9��@]C��>��������э{�\���5W�Z���c��ըǘԑO��o^��+(ϧ�)ߜ����K��e����$��!ȜP��FU&��FV5`�+��_��T���u7����A' tn���#
��ye����X�9�F��Ƣެz��R��k��H`~�鼽�\9j_���#��'z���5�_��5j�X�9�VB�{�}�.��P��=��}� ����͊���
8�"gU3+!`���A����ʛ4q��)�Z{�x
&�>V;M,.�VM�%��r�Ύ!�ߩ��.	O�R�3���a�$'�Zc��#z}�n{*�]�2�1"��ĆE0i6�e�����
�Kpf�X
�e�����V�T�3�4�H���oq_��~}�T�����iS�C2��w,�]�b]3��<q7����#��o�?x����Ě��F�E�[*c����a�V-P�췳/��EG�~�R����A"?�ߨ#|&���G?�H߆��%��,2�"�u��_(���5�%e��l~�c�=���!�D�����R�+�+��\.�Zbn3a��%ႡB'Ȇ���\�����l|������F?�Y "]�F�;մ�8�(��b�*&�X���Nte/�`��\[^ خ��?��E���,mxNH���$�vj�mR+"{-���n�*O����#u��Š�P�rUB����f��[P6��-}>&*d��1�=�>,�0���aZ��a��}|<�r�d�Z���AQi���t�+�t��g[8�|�J�Ǝ����\Ҋ�����_� ��%�<,7��l�=�8���F"�@4�^ܠ�L�(�(�?ZeSR�Ό���7������dӭ墰��E��)��*v��@���6B���a�!>L�N�:��q��	0�L:��-4*펗���0��)��BKz��CМ�����E)���U��
����O� ��G��b��sp��J!$	���$Ux�[nn�7p��z��	�pm�Eh��ԑ늋
d�k[���z������C>u�S�WW87/�$6T�ۧ�U0usL���2�I��M������?o���N�+O��ۇ��;!/���$o�� �V�G��;�V�!��Qi���5�E�(|�`H��9�B�
����qu{x���.��Ԉ��4���/n'�և���<, ێL����I4�c�����N�]F�ݹf��̈��˹���Cm��/�f,f�^,U�ԧ��빔_,7��]"�0���j����+�%�Wd`H��W�$��TF1�׬���c��`ˣ�8�����.ޫ��[Y��v�,�4�=���{���s��ֲ�Z�j,'�Xn��{�ʙ���yG̬��o�h�����d��+��|x�8�=�9��ڵP�Z���ʀhּ��',��M
�Ŵ��ZU��\��L' M�P�czo�P^�����j(0��y�ZEQ�jW�@��V
`��k�i�jyN\�����F̹%f���b��@|�QB�W޾�V��}bpN8�-`7mWIc(47�Q���ɓT��P�W!|-�K�~�jAr������؟����
-x��+������ӈ���gʶVI�r�0�pBШ�8��Pߘ����Wݖ�Q����)��[�����O%cr��)@�{��@�io�ྯ� l�0��ژ��m���
�ORz�xW���4�F(g�2$�G����:��۰�Vܼsj�.�(H����7��޳�����ϝ��^��F�M���	
ĸ��C0FF�f����`ZĨsR_*���<8.����*Q��� ���6�ڊR� �Y�B��dR�p���5ɝKb~�� ��l��qR�it%� 1�I�*���6��4+�����b
���ȧ0��X�i��;�v]����y\
1�Ns�py�b;�}�,����)����W^%��޸�9,ېeԝx*=^�p�BD�H�\�ޥ��9PP_�;_J����dϴ]r�O?�X������V��|[K�W�{��;�>�Q����!���o��'�ۢ�
"����_�v}q�#Ei~�B+A�e������g�C��Χ'������	��%�D���`�kO�R�-�=UghI�m�A�3�	v�^�y�E�`�ϛf3~%�(�����w5�lڪ�'1����$��f��sF8�fY�H1�mJi�0f�y��ɳ�.;��|S���;GQ ���N��E1?��7&z��!�@���AW7��ؕס]ƨ�i������ys��O���9��kB7�c�Z���C������7����H�=�����R�<2���@b����Z�v��m7b��i�f�������E��]k/_�p�D��$c*XS޴!Sb"K���3&�336��y��8�X��-�U�I5�r�l

2׭�s���4T�x�#�0��Z�;Z5�����Na_�Wۏ�͹Nޣ6M���캒ֱ���c������oe{G �+��w��)���&��A��,ف�Oe�������T�6��	p��Pϝ�J=H5uY�2��qq�-ޤm�c��'��b�w�2���`_����O�������0�I}X[ĵ��[$��P;U���#��<U�yd�)4P��8@#�[�U3c��`a6Wɋ:��␖���L��Ƶ�d��1�/��C�$�t���@����;���l3��C�Ѭ9�h�������R?a�x3���V֝>�EYU�A���X�(9��ܥn�]�f�C��;�d�+��n)���j�`��%��q��˭J��TH{�KpCp�I��o�s�w�=�,�Q��՝�Hv�㛤v�z~K��XЊ:Ǩ����kx5��k���t�_r���Ej��Č34�\E������Zo�@���n��P�x,3���f�[��1��K٠������J��8*]�^�B��a�c�O����S��ޒ$Y�v0��Y��_��i��Q�l��NN�4˱�	�_!��t{�G� �N$D,w ��,��L�A0�h���A�U|%h>��R%�e<�������8��`x���O����T���Q\}ɔ�|ȪL�ʐ%v���V5��**�X=�ÝP����ʀ���P��>�D/��̷�Z�����#c�jI��d�1?�n]·8��/����^*�||��\�w�^|X���4hp~�|�ߴH�#�\}z�3MA΀�m� ޶���g�(��Dp�t&�箸�.8���_H��gv(�<�m�#��gعQ:��jN޴წ<����fV����Q�>1���'��$�\:�[�V�~l���o����>@�.������V?a;��qE��osaj���� �H%q���e��\4��F7�:uAoMa��W�T<�j-&���C���_9�I��0bc4��lٲQ���6���e}�t뼳?p�7�8H�rv
I�}��H�����=�����'�k��W�����[��6�e?+!�̃���yQC�4[�
��A]Ѯ�Ĩ�K��R`v	c{�^�� ���Z����h�tA_�U�R^���-�2P�߹to	��	��B�p���`�&�[�e�k��7P^��h�������Q���i�Ұ(Dģ�}���>D\ݔT3g�|ky�c�"����oY4��	ڥĐ\}�מ4���~ �ZV������)ӫ�w_UO��X����95Q���r��ΫI\v�����
M8���i��>�z������]v-<e;l-��C�Ȱ�������֚2�����tQ��Qe���ȏp��?-�>'&�u�r�z�~$��U5Rh�X��'���O�(t�o2w��	*= �e;3�ɺƄ�N����H����3~i��ܛO�΀TC�lgG�뻭4@�8���_�7���w\�+��0}��-g옄 �]��k}����3J�ZfÌp�-uW��LjVf���"U�f���{Ta�Ws;�E5JLTaO�2 ���*��0�����a�רv���@�r[�*0�
�旹B�,�({`�U�Ϡ^>�ȫ��j)a�hX����]�ӐU�*���
dU�, ���w�F�(��MB�%.Y-w�����·K��w"�v��:��\����#KC�_ ��pXD��,D�XB+͋7_"�B7a�cR[���=�Ȅ�g�@ϙ<o�)��S�]�]Yy!������B���\�Xf���~�N��1�~����6<Y�uu�X��_A�1y-e��h�����2�}�[��~�Ii]4�x��C�����@5�p	?����l�z�0�i�Xl�#�-��yx�

�}�3�{�'_�X7a=��NM$���O�;�n�J��(:ډ�jٰٚ](v�s����qF��"i��L�� ��h0��Ӈ����?�eܜB���
�-���}%��u���o���-*��+x��u2��T�	�2���Ee��{�
������7��\zM����7ͬ<��k��`C0�vbm)j�5�3�w��' Ш�_�(�N�ma�L��{\�.���m�Sՠ��UD�U3%���Y���*Wt�4Ɉ��#�l�,���#E:)�D��n)g|�#��O�,��3a'�dɠ������x�i5��v�J�*0��(��kC!V�������}ѐ�Z��!)��Ȓs�j4Ss�>���"���hH�dD*\x/�l>�.3�dsھ������.C��l݅�J�)�Z�?{��K���4����<�?u����)й�]���L��N�B�|G�Э�xi�@��?y��� (�Q��D|�흆�c���A.��.;�_�/J�30;��/'�p`���;	b��[���H~�_u�I�ӟ���dg��w���#�$�;�r����4�"�7�-��2�NuŹ2��W��z�<0�I'�',�O�i?��!�~��^M ��|B�I���Q���9����
�&�Fd�V����d�
��j7��`����6��Baz�%/E"a�1�V|w����H��k|�D�pU��p>^kr��e�T��H�J�<�+S��Zh�_��p��|�^	�ڻG>w���-E�M'�}5�#��Ë@��[mb�#�И�vȔ���\�w?�-��ug\Ӡ��<�=ST�o�b�nP4�(����}����n��Q�#�t �͟J&W؂�����*M_�������:���)51�Teg���Ϻ�QL�B�[�p�N|��s1��d�Lr�&]}�{������ѫ���Da��n׃��d���~e�rS3��6QN ޻���<�\�Th�l����gy��K�2��}��Ɉ?I]�1����-Y�}b<?߃���&�0	���N��hz$��Î�r�b����'���r���E\�H��������( 4��9!��ʄ�K���<݁����\Zj��.Si�:*C�6춁��,:��rM!	�-�K��cI-볨y%�!�N��ϛ�����d$�?�8C�!߇�Mu&C0���f�F#�ha�9k=�2C������
�.�����~��V~W_,F�Q���T<����0�tj-W�s�`R�M�q���Zv���mz��ޖ�<D��J���#c˨CRI���!�1�83�=��D�$�vn�u-�C����A���M`P��Bn ��!�Ee�#��ĭ=�H��^ו�5��M}�J�:�H��d�W�V�>����ñf`�������Z�Xpi���c HK_���r��W��t�e�X���w��7/I󨉣�]Tñ=����X�O�J�̧��n���Ϫ�]���pI�T����E�����K���t�U�t�(��|�hc�>)��vS:���bߺ�_]H]�9{:Þ<���i�A�Je��2K�85M�ż���bUp�%�0��$�Ǎ��>���yo�&�1\5
 �;�|��+Jf��`�Il�;�C]��lgVJT8��e/�X-�o�����~��o�����{x1�j��c��3�p��ZuE^c�A=؟�" Jg��&��G���9A��u����}U�#��n]]1���v^��BB<�c>���*J��C	#��ۈ,A��n� 5��ᦐX�hD�p4��W;�&c��J�j���Z��C*|���+�`�Bݯ��bi�A�~�+s�Bʠ@h��A�U��Ee��1ɉ�3���T��#����E�� ҿ�A��)x��pa/�nLij ˜�a�V|�ORq.v	)�bc��.rijɾ�f��� ���ģM�g�,m�n%1*����|9�qZMqΘh�W�r?�"ҳg5�����jX*�?�g%�����yJ�� �$4�Uq��P���sF��/ʆ��8O3g䄸b7�C���쳠��M~_��%�uDb�9�O���_��k~�4�a{�I�7����������UM�|��2,}����� �F�f�xj����=Bs�e4*�Bmz�x*�$����f(%��>(���������æt�i��R��	99���b�������c����8���Nλ�T��{�XX�� #�Q�.�F��a&K0̘Q1����O4Z�+th4�7��5Ȉ��N�F�b��[�7o��o�|�, 7Wܹ �Yb���A9�7O>;�Nx|�f�=�@	��$�є����y���� ��y1S`ji�0}��$�H���-��- ���$���,�L������h�E�e9�ñ�!Un
��M����E(�G,��ܩ��6A�Z9��z���.nww����}b�2`�s�<��	:������if�c)�d�^�ǽ�Dz�T?7p�Hv*V:�[
ͫ�����n��#5O��yf�w�"�]�X��7A~a����*�}�m��n2ŭ4�^B�R��K�k�#�u15(���S(��߄�mo�] Qny���{�
��O�37�O��|����.��weٵ-Y�ht��f���ʌsҏ:XkwE��0�Wu���V���,_E�J�HbTDт������7��ح�>�(��J�d�&"�+�'�P�N:֦P?k,��TV���$/�q���_�������:��x��Č���l��C��[1A����s�.�� <�wUFo�+��c��Aa�ԀG�A��jt��`y��M��Q�����t���OG=c�z�q���7r|]�A0�j�Ae�ރ,���(�8U��Q� /]�h��F�|�
-���ﮋh��!�v��c����=��md#�`�ž���~�ت��I-�aޔe�[a��$��)񚪙�TUK7�X�.( �����c���Վ$�^.����x``��`CγS!Z�(p��s�LB����Z�wɈB��ρ��1���to��7�b/��$�-���t�㵿�7_�.�p���F�7o�䖼\خx��C�ȵ����G� �7(����Jy�D؆fC���J�9��ϓ�mH����@���>i��T�m{H+,
C|A,/05Zm�CG�s��{c0!+HmM�1HN*gO�k�x�9�bO�w8N�Q}<u�!���~j� 
�J�*�H���p���KG�(�� G(pz�q3\ �u�=`��3�L|.?�Y<���}���y|�9��������Pm�� bweX���?��ݱb�%2���#�DQ�����·��-v��f��q�	q�����4{���P�xv�)W��O�G[|q�}^��4��c�_�0G�	�����^�O�<L���-��<3y1f� f�㐨�����=@
Ѓ� B%t�F��W&a�y���Lӗ7���eZ4#���rn�q�H�iF�X��2�F��3��7�8��Ȁ�;֟X���o`��������exX����9��.E4����t�w��a��^���oo �:c/#���Zy��;�/7��;2;�'y�l�2�2�����.E�ǪkTC�`����Ⱦ�ˢ����]�1v���&E�Wu{w��!��%L���/�~��I�Q˂L���/����A�EslZcD�w��A�����9��Jh7�1]�������� ��A7�����Y���3;��ģ�:oZ?��aȡ �j�.�)��nLPp&���/5&��])��Ò�sW�՚��x��R�EWf=�>��K*R���q��᦭'θ��`�w�\�d�%+�xfq��.���lYS��isAW��c�������r�"�l��弤��dϸw�w�� A�P��x�O:�cR�
ᧁ}���`����5�-9�}<"욆��K2k�&b�ńZW�V�0F
n�T�3�R���N�gHxpi]�l�~e��g��%�Im�[�F��"WŤSW|fX��K���3�{6¹���-qd������#EBc+��S��\]Qӿ;�;v=�1g��-y����~In8U@�V	tp���l��.�e�O�yۤC:�p�/`=ޙ&���\�����T���� jqu��W�Ď�f��9�h����w�j �L�^�� �!(��<�y{&E�k��y��Q�(���i��T�{iDw1:�zsH����5PvG��L��Ђ8x�Aج��JJa��:�"�`������N{Z�b��xdfu5(�����ڞ�+����I�l��A���>�����U���1����)��G���:�^)&�4�n|�S�;b���`j�դg�3-�֭�7�k��IWJ����"�6M�&�+f�����R0eH@��;��Ty�9C�[^s@4Ͳ����q+���q��E
��Ôc�{�����5���ׄ��H�a�>��f�hq�>��Q�<����(��a�����5[����ϘU��:��Y�7�U!�c*aهn.���*Ȭ�N����c^��hx"в�9~z��'�Y�>=�q��"��bK��ٟ�0� ��+�\�ʄm`&�êT�W�&Ϸơ�9�f�B�8��j���
�^r9A�4ކͬp�zp���;�T�?d�+Yu�u�$�ϰ������Mx�{��>~��$���ryC�o+ՠ.d"R.*��6�f3��A�7G�!3�����|�%��L`�g��(���	�`
�V�;J�rL��y���tg��VA��\��\�M%���d����r�K���ht����Mx���A�a���!�Q;pvr��34h�ҭ�P)�Ҹ�rH��F=���;��﹯Z^oyJ��Ʈ����ʭ2�ԟ�e��Ƒ��8�� l����K>=#нP=TM75��K,N4�
�8<�T��U��:K u�Ƀ�|𱡨�u���S-;�����|�Ԧ|�t7A�[="êp�	f<͓���Ի��%X��o|-�/q�]�c��8HSn�I���U�/)y����Fu9�n$"�+}P-���P6c����يO�s`�p����=Ӫ�4�q��}!n7>�"_*�
C����>�X�b�)^;z���յ�,UB�Em`�_l���(Cti�D�ʽ?�]�E�E7�7K��-R��|��-\f8�|����� ?E�;(�>���p�d/ض~W1�ǡ��c6)����>kZ�7+��RJ^L㇬���cɞP�U>�ؒ8��1��*�OC�����
[�4%?��-�;$��dC�p� �[���ŵ��Z��cA�Z�^���~l��G[�w�Ѝ�4~ ǰ�/՞��!`���Oa6Q1��E`RW"@SL������Cd����!V�v��ۙ�t�<�isV�8�낛A�1�H�?�ǖ�.�[�'����Ns�Mu�$�����ؤ��Z�{��[hy�b���p[�u�D/��� ��Hb�W�o�����>G�e��R�ӂ�+���P"�IWz��Iv�z`M)7���{��9�
�w���_L���6	�D�SƼ:/��N���6�	�^Ξ`� ����j�:������#�R&���Z̒�	n�I��� oH-MA,k�~c��{��fZ֪��1�oפr��w aOEӥ� ��Z$� �&�C�S��u��7{t^ȼ�\�����y����-�Fץ{g1Â2���.Ij7\�虘*XM���:��_��ިx1{Lp�p}� +`�]��wis��^V����DUJ����Nf���H�lT�K�7ΑIK�� L�R���/Kn��g�0ð�+�<��p�oN+a!����AT�TNRn�#1Q�]d��|_�c3����U9�Fj@�JS�E��b@�����c��!�d�ͨ-!�޲\[�ۊ<˽8��ͤ�Gp��:�s�`R��3[�ӆ�'*����KL���7��^�zB��s�Fx�W	�!<���S�伜	ꬖ��BR�l��a\Z�d�R��x�㮟��p>7��G��ܢǦ$Wg�|�`)�?�c!���;���t��v��^f=���!k�����Z\W:y���;���P��8"fV�>�F���O;��K�-���ܕj���f���l����-[�?�E��R�O7����z�.� �`���o���nq�E���`1�4~�5N�*�N}j�ݽ	�14���+�F���48B�X�BH�˵{r� ���(X�ਯ)�݅�&[i�?-�� ���YW�#����
�`!����w�#X�����/9�Z��`��gۅ��V�@Q��W��e�Ǩ�M�"�xP�t�D!��\�E���c�����5����T����	�Ś�O����F3��CA#t7��I�r��0 �����iuc�tJ�Ȃ�&z/�5v	e�n�62�w�"B�����
,��(]`����_�ï�c���?��AT�#����(�F���?��>P~&4�7k�bT��j��8WX��&����?��0]�Bu}|���{]�s��=�4���jA̢��V �F[.�2P�Zg]�Xv�i�R�����|M��$���d�YA=���{��ÿ���^��'�k��D��W���Zf�-�pb͜�c��d:|W�;6c��Dա�Ts}H��r+w	'!_5H;�.l��lu�g_> xd�������:a��l�/��M[,�5�%kP� -l)�g�ߚ��R�X�쒿ee��]��2��R�W����}97���\�3��74
�3j��������& SL�N�"_���)�|��ț�0|�������X~{0�]�]H���M�:�*�L��)��_N��2��:�i����X}H��)u&�{���CK^�آ�D��`��t����d}s�n�@�e�{�k+0_��ɝ��T���\���	�Z� L5�?1"$��4�7���yf���G�]7�:㌦M�����n��2��p��7 QE�E�@��}��w�џKr�wU#"Vs�S�?LYyX�����v�o��Ǣ��@e�m����ÙAH�� �5-�
���� (���X4?������l� �aT �:�p����j���uwx���#��b�ҌmJ��6���4��(@c<� �Xk�W��Ǟ.]Y�ԣ��b~�?Y��ؚ?0���nC:;J|�]6m��g,�S���nFA���S��_�'b�Zѣ�ŉ�sMy�%+���L`Y4��0oXlH���$��qy�d�*�2lbC����Ą�GYZ"k�,�&�ѮQ���Uz=,�l��9����><%J��:1[bR��{
/��]:#[��!s{mм-o��Z)a1��̈��x� ���WM�G�B�q�@���M��>��P��S$�N$�Z]��HJ����6M�
�UV֑���"e����ք����Vo,l�F�a���z�vڎܸ~,��0�ǽVM6�3)z�e�l�yt*T�;|�ߟ�Z�M��!I��o�����樾�k�{�)��R���e@�ӛ�c|(��"���TV�s=�� `&�ڡ��֫'y�..I��1�I`�{��Tx3�U��v��9]UFX�Q�v��8vD�����}UL�9�ˌ�v�jFG���M9&���-Xh�΋X~�奒k�I	(y�V�ׯʃ����Oƥ���{Jt�5�k:B�fW{�Ģ8=}�!#|�W7%r�Ļb���@��j	�����&�BnB�>NS.P?��VV^!��:��þ�H}�rrv�\*�.Z�Bl�|qO�C�&�p� �|��_@X��el¶��vt��7�RA�Wb�,
_�
>
�\��ᡊ��n�ظ�?/5^S��:�+�.X�
��������|�Ѩ�9����!O����uM���AX��~�
�Y'����r��S^�0�Xsa��H$n�����X5!:XU��_����C�@�S,�I��`k�M>e��$��u�˔»�vUx�|�沯����kK���1C�sȡU��髖aŋċ��A���w��,��]s:Q"���*������ɰ���ѤsZ��N�;�q��X�����H��M�~�0Pg��էwd�⻪>e~�bx/!
�q\�3)��V�#y��� �(�8����H|�N6�㉛MRA�xx�|_�g7��GS��oF����2#��g���d�a�{�[��уR��7���;���6$�ԓ�'>cʼ�{�4�ktg�S9+�d�SIH��\��mt�����PI�R�1����-y���Z>��54o�^gr�(�\�b'Wh�S��jģ�(C��q#�+����2o뻡R���3�;a�¬�V_��F��pgl(���U�g[^���6��|LH�0j<L���޲�����wٸ+��Mj������bX��+ʢS!�D�!��#��+��Z�P�?�0��{�I��
�耲G�f���_8�_�_���`���Y3o*���rA����%��y�4�����`�h���{�i1�5|���AZ�c��
\\��%���콅�E���&�h.�A���>�P)�9�˰��`TT={+����Ov���j���pЗd\vj��NU�xC�D�I����_B���;:dm��"=�����.��7��6�y���}�zpJg�r0�l0&�FGc���WZÚo~���C(zx������?�(�F�aH��IB�K��~�H��b�)��D:"T����=Lo�ATMG�(H�D7�/`d�qI�V��Ds�6�X�~>7����׍��),�R��2� y
�IR�ɜYl���R�65QG� ]�~Tě[|6�Z�9�F^�I��l���vߪ��}E{O���Z�.'W{�>�μE�킩�I߅�����	����:6����[jR�o��������?���-~������e˼)�����,�vk��9��w�ؠ����q@��`q{"ف/�_�\ ,��G|��Kh�]�Y;!�z�f�DO0�|z���9�E�#�X��M$o�j[A��@۸IAx����$<"���=d�������WԐs-��N{�G�{,�����?�����ɩ�	w�9�g�������b��$*����[ѽ��d �W����b�_6U�x���M���ޤEf��v�1�kGQ��i]��������6UN�yr�N�i����������e��� ��޵��r�Tn׎ם�/=U��|EО\Y\��!z���3��Z��v�Ұp_�O��(���]���a�^F�ޭ��@���Zb4�vJ�{-�Z�G�P]]�D���K�7�\�C��5L��h!(WQJ���]�O�5ߠ�m`��i R	�����y�
����
S�E%���	Ʋ���9c��ϸ-R=z�/=I�GlcK��W�!"~Xr��E���h֋���U��m�|��Lp��$�5/<�s��ͬ��Z
d��7,��K�uo�L�П��aS,�F*V�h`&�4�]3#��̀�/U��i[�\�ׂnd!hf�:�&��I��a@��a۰��k�r���ᆣy9�[z��Gw���8>��+O	/�h1���	w��w��9�y��َ0�c���#���w�SԜ�s��aE�H�{t������A�Ђ�&:��kf3^�c��_�5�Ճ/��m����9a"��\Q\5�3���'�J+�N��C;�+�l�u�y�D�Ϗ�|F�ǰ�(;oP��T�I	{5������)�c'�ơ٦�J�����@E~�0ǹ�{a��U�,���&{3-[��[	�f�7���R��)��Ι�o�h��f��6�m�l�뀰v��\4[��~'���`:���p�9�g�ã�R55�+w�"ۃXe�e�����A ����C'1�w�F�h�3�X4P�UЎs	p��9o�m�%J06�Nc����*?T^���[N�(��|=]��_Iv{?!����K���c�=e6��V�� ���N��Lr2#fz<���͟FgH�����Wh3���kn�ObT���Pc�<��1�#+Mrg�T��-"�(�
�C��;��ԣ��A���@0�^׻<���EȾL�����2���=�Kj�-��S��K�49`+l-sQ{hcx�|C���k�m-;�r��G,N�uC	�5��x�"$n�ϑ"�Qظ-�A3Ф,>�g`c&Te	�Wh��)O�&�3h]�hnz҈��͞)��Xq@�����Q��D����<���oI�9	�$�CG�Ȓ��H�y���$�j�7� ~�F���_uI�b�"���\c"�����.�<~��UI��I��{`M��cB"�5x*�U���wm�ܞ�&��ʫ�q�rW��>�����ޘ�1�R�n�)-�h��U���f�xy�p�?B�����z��b�ze��,cq7�e��/J�E@�E�Ӆ��(�ѕ���:�nЏ$�����:(��@�N��#?�?�9�4��ӂ��j)	�*u/�ҿK�)�����d��.���U��OM����� |�x�KP���@ �7Ĩ�_*�sp|�-��3���S��3� z`Čj9�H��LHFk>�7u����b,��0�˕�|FU=�O�!���5k\�µߓ0��Lj�b��S��Զ��5�%����z�'��!xԃ;�x}���j$56P����Y��a F�sq,�����ޜǙAcܹCD�|�*P��d�!�� ���l #c>"N��lL���q0�kh� �:$E�&v4�2��ՙ��	C�(���%>��]��4�BQ�X�/q;���m�խ%h$�=�ĝߦ���,9r~C&[��Ԋ`���;�,���a?�ǞG�$QI/s�`�Z�[
��)P'���W����H��?4͂�k��;y��@,I	ۣ|8 3m/+�:ë.Xy�z�hY���Opl�{�ZS��FTG.`T������1��!�-�1ƿr׎h��B�v��4!�a�>	6Z6�b��];t��e���.����{�ʶ�8<x3�����;�H�R�-�nyC=�������K}(����M�me8�D<�7X3�D�zEٜ�\l۩U6�4�"�\��kA���=F���f��K�(�YlR�']h�Y���d����ݺ>/!�B̀�;\���ӈ��5�Di�H$J�������c?vl��F�(����`��U#n�Ӛ�Mu-���U)V]z(�ZE���bP*o�< �쟭ظ`��+f��Q��8#|�F��<t�}���d#��c�>��$�!E��1��z�iW���ů�x��؆���h��I�+�n���C�%�15G�����,������G.NzJ��2*+�����k��;9r��E~?E|EE�jW41P�s�Ӆ�Z�T��%"�,��r����2팖8y�'x�f��+���[)�g���(��n��;"��1���4"Lu�6�?�6`�[�E&\�HH+��>�X��0F�A�T)q���$�/�,�qb���|��?����v����ͬ'�.n�n��eXYj"w�X��_F���]b����]9�� l���Y<�0�<㏾�@���Y!~�:Yڈ���T�/�R}����zz�S���J�Q�'����!���x���yr,z<�+�6H�1`ڮk�Q�2��<�#�rN���@�E�]uÒ�;.x�I��/��t'�Z)*Vu�Q�����nU�QMx�xƀM}��iV�~'��� �T��Ksqv9��2Y�/����ޭ��_� 7Ԁ�|��&���ũn�Iǫ"�j����F4���uE�OC\_��Y����Y M���>q;AS�=jڻ��O{pR�ce]�׎��Q�tO�"MÂwǑt���qzK�'�8h6p�~�q��߂��8��x�S�vߔg��X���$�S�&&Ē�q/��l�PE��#F�O��c�� y0�3|������_^j�� @������O�H񳪞�I���Ε���hbi�ғ��.h]��,�f�z�@|Qt�F����Ų���w: }���%>�cK�6������~H����� �ܒ��"k��%�w����2�#����?=V���ln8��U>�t#�a�{�[iL�9�هx���+�h�R'���6�xzhhG�@��Ê��O8c��E@޼yN��Ǳ��`���x	j�����%�A��Ľ��YeOp�67Z����kim��p~Ugͼ��']���-lј�D4�]�-�F���3��P���~=��>`:�FzJ�e���dc��Ǚ6���� C�mS `l��[#����	KR��_i�X�I=�GK0��D$��a�-͛���6����W�]y��?Н �B�>*�&�~�X������f�֪�v� DxY5@��ǆT����r��F�lA���n'�����i� <�e;s��
�(2d#��]Zc��k-�!5��j�GO5�w.|}n�:.���'Y��� [�VDW�y��K��]�';��2Jp��}�Ԛ�.uHN@�WkΆ݌v�h``ZJD.��V��@Zd�"�?�@~Ā�~��fn9�I��/�՘|�����`bR���m������8��a�<S�3[?/0���l]i��H�w�E;������?��k`�;�����g����ר)��D���z��!��xK���'�e���]�K"-	t]�;��3�-iD<�x.��n��J֎�YIM;��7�0��c�T�,�����N�/)R��>���U��R�r���l?h�5C���F�C�Om���N��W�B��M�W_��_=�`�U���B*�I�/��T9!�9���sL�b��ֿF�������S+ۛ�nq����?���J��6�`:Ӡ�\$2G$�'�o�|��З�ΰ�R�T-��R=��q�d�j�D�[sI0��`�&����.3���\�/�h_�X�%8P�P��y�µ�_�W��/�
��S��L���9d�	��.�L��Yjs�$�~�0���G�ú��L�],ևd��ў*��K�DZ	�2��Gs���b�W����O��iz����e)�v��H
*�$��A�pڌ����)&�#����lwx0>��X �M�9��hf�����t��e�)�K�tW���G[(��O͂>@���8t }�5D��m����n���&$�=z���cn3���	P�� 㴧����r��<�S[Z�.l���`��W���#�G#D@T�uҾ�0$c��H����l>�N�uk�y�D�ɲZU@�/��U���1L�l���_���-�"J�
	��[u(Bmړǉ9厹3��7��S�a�@$�q�ur <Q��-�	D ��r0�s�t�v�=�a� �6���/�l!����D�V_�g5W;DR�$���XF~O<�:~�'��9������TzBV
ϱ���(䈭�H����C�5RЭ���&�ȿ���t@�=&#��nw�w��Zx9��P-�:�~�Ζt����)>[��*q���W��b/ꋉ�Xx�@fEs�w�Tl�r�v0���tn��j]�L��H���"�|��2y1wP�*�.V_�MO��1R�a00h%%2"g�bd�M�7'	��#�0�XH ��L���G���y��Q�ycjL'�J+2Q�S{�44206d��l,���\�)m��7n�Kg��q�n0#�	�3����:��޴�9�v�� �q���um}:�u���B�~wc�3ÿ�$##�@��aqYu*��e��< 4W`���`fʍYw��Y�RVm*5�����u���!�us�gZ����qԥ��=m[�K�=����L��,�W�����f�tx��-��Tvk��M7��pU�+M�*��u���"��j k7�d]@�����g�""��|�s�H'�\@�
�(Uu�pg��d�"g�%� ���2��3�%�AĔo8�.d 1�q�c���� 9������g��g�Hz��q�Q�)�X�����q.j��l$t��C%ۂ� ;u�D �1��jRr��Oe�|5�p"��\�o��u: ���.auN!����J,9�)�G.��kݽ�US�M����K��y$>�q`Dfg�P�
�.���?���N0�T��';&�`��{����l�D��h׻�0Ě�Jw;(3�2}��eЌU;���0{)��@��a?`�ɶt�p~���#��Z�����k"Xo�9�s}�Smط͒���t��ʁl�������߼���%�Y�*�jq��}y1⧜�)B�Z~'�rh�՜������4fe׵T;��D<Y㎺ �3�]"�>�0�WǾ�3L�������ޠ_��҃|�.��q>����Ր�B(�޺}Dx�*�V�m�&��܌By\q�ړ|@��Vj�&��M��S�7��=�����ZSU�V����k|o1�H!�7�N�T�۞��*���婨�$H��("��a���C�s�`@����/��G������x�EV|�}U��-�9�[8ߦ�>�t���qx�^�].O�r�W�}+_�,����S��9Y�>��&0��s�^R<@k}t��(�G�<R_d�7�����F3��7�ƫ1Yz�\�I��˸��h+oN�4D�oƃ��� Z�F�%L�8X�x��$�p4�y6(�B��i�et�:��]���q�MV�xjJ"���cц��S)2�����V��G��a�p`UfZ�9�����91 �@_���4�9�i�/PE��"j*�kf�{;�0݅��Q�R���jB��f*�LGM�����$%Z�|<��Fl����S�{}@�u�(���5�V���co� �P�i��S#;�N�׫G���Xl��ЧI(�}ʠ�i��̚F5����Y������t�.�Qd���
�saݔ�Upb�� C�3}s��,٠T�V��e�jNll9��&�ϓ�ƴ5���)q/���҇��o��B��zُ���x���d�10��n�-(��<�6x�3�-�d �?�����:��r�'�Q��B:6��
�l+�6��&.�'Z��l�xd��ze$ӽ���x�7�E	F�̷��o�s|}R?�-2��B�������3��55�OZ�MH����	o�}��B�]"�:���K_��y�g��Y>	]��2|�5��.Y9.8�IB���]�<k�(�Ά��(E��{���e����&�v��
,� d1dˈ{~z��'��Xw�}	kՓz�ΐ��F�/l�8� �Ml��Z����@��X1���xHy�$m,����ҫ6P5��#(�1��	\7�#�����#ӑ�������.fm)EM��{X�<�=sXM�-��/�M�0�h�t��N��Ȣ�߱S��8����l��F�������T�F���ݐĵք�w)N��DK�"���S��x����T��7+�x�L��;���Ќ�I��_2ޒ%4+�����q5�h�$�c�X����N���oW��f��}=��ݓ�+f����S�D�#�h�#�Au�����a
����'9��ʄ�-��X�IK�>��GI��D�"=��Fo��i�����(/H�:�5�dV�'w��І�d��9�B��1�.��E~p���`׈�25���V6��hC�o�J�	ً��Y ]cWց�{C�����B��bK!"sہ�i��I\�����ُR�Ef�4�M�ݿ5��X�.q�+���3�VbR]�!u:#l�3�!��V�H�6��뒣㴼��룗�0��.�m�?6cPK��??
x��머�v���q �-�gS�)�chq�/E�
�,��-N^�#�x�Êޕj�ݕ��ۣ�. ���{&������y^�u�Ia���AǷ�
b�T��N���-�%.g������P�`����_{npoV΃��h�n_]d,u�7�ǽ�D�p�tE;�@[��!�@�m'�K�7�e5���n=�Š�ޑ�<|��нO̰+���"����I��g�zR�1<Г��&����h�e����~�ʂ(?����1ǃ�? >� Ć)����GG���j�R�B����(�?[�CE��n+�L��wO^0̞Sb����Jѯ�L>_��fc晰�	]kz[���(�`x<FK�`MLQ�{���7�f=�=4~"k�n��w-�����FSV��nYo8��n��Z����m�,�N�V��;9�GVVnG%�����.V^����_boOzzeT<�&Du��=ʠ�g�@��L�)��,D&ϔJ�N��釱�������Y��q�	��/�W���d]Ok��~Ú(�مw%%��A@�������W�u�[Go�V�cܖL�D'6���7����9�'�c�r ��j��G��9�`���ө��A돪�P�	�Xrnu���6E�Hp'�3��^�?�M����d�m&6���!*!��A�t6TՐ>=��<ܳ�!*p4f�D���ł��.��â�\��L�'�.���&Sl�i�H&(Ŝ�b }�(�����ݸ�~\��R��\�M����{g��.���Ao?,�С.���bo6��������d߸�� ���S�"
4EJ��ȉ�����}��_p����A퉭�Om�k��'E��/!V3"j���_bS���@vǚ{�7lM��^���kRϴH�Ȼ�V�A�*LI�����<R�А^�I)1��VP����3��)E7H"f��R�9�?���Gބ�u����M����B��S,��}X^X7OR\���n�\f΁���rkm���g(Qz׼�0� ѳF
p�E/���%��~g�	T�h�y���w%_�Uoy`�G�fT��s���o���pX��Y9����p�F向-K�G���"�2zCͬ��|0���q�u��)����`�(�. ��c�ۣ���^_L�z'V�����6��)	�Rʴ�����#�R�y�ġL�x�s�މ������� �t�\.�+w�WI���dN��Q|2�@��<��AfVjHvPȃ����1t.P�|e\(��Q�C'ؒ����lyH���S����5��d�q]a&����X�%#�8��&�w&�H��ǘ�$��x�;W�����aԸ6�#Hj�;�0|4!JP37~+E֦LdI6T�|t]f#于%�������Ɛ*�Q���ؑ�p�CW�C�M�b��}\t���V�lC��Ccf�B&��
<ޯ������>��i���̟}VD �L�x��4�z��"���,^�^^��Q2�����Ʋk3�F'�u��aX&y]���mDk�������������Ȧ'<|u��_{}E�j��]�=z�I�%�XYOZ�tN�_�>��q�5#N���=׍�t��5�u���E4Y�� O�p��dH��&��"� ����T�m�W�>�49���Tӊ0�2��H�t�ơ9ùW��8.�E�^Z\9��Y�tr�I�~q*�[X\����"b>�fn/���fFdF�jŋ0W�9����z$����Y^�"9�n*g+��2�#9`D����3WN�'��j��ZG�ιxC����X�?'�x���F�'%��Z'��C�弯W��%+��f~��� [��E����b��hi��tfHd��������f<gՕ�	]cz�Ow�׍'t�ڌhj�R<��/�]�w���6�Y���nB�67�\�GP�鸠Aиώ+�V���M�$�2�়'��O��H���Kԫ��CCh�u��@�o�6��"0� ���V+�둢a~�S-c��r#��^?��rN@����u��~�Ű�8�hM��@o���"xl�������%�������o�ήWÁgCN���k|���r$)枡��o漸k�q�L��N��#�RuRA�S:s�^�}Q�	0+"���B��#{�;�oD�= ��W���A���յ�r_
��ꉕ���K@M�vd����/�[����V��nA׀'�{�4��ח�	vԊV�e��nM������ I���f/>J�:�{�u%�8�f�T=��:�r����O��8�k�&E�wk��'��F���>����XzX�L2����j����]�4��ǎ�O�����kp�Zѱ�Q�&'��:���Y#5���t�>{4`$;�ף��pժz�}[N��!��e����i�