��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI���!qp�6ht����B;dv
�[�܈
�/���t�!HO;���;��.$?�'�-#ܨ��q�X `*Ƈ'�e,��Sg�Bno~����1���V�0HA�=/�c�����)7!/2�����&��������N��Қ	Z�G�i؈�7ХP��^��S�T���4a��I����Zp^�B���,��1�W�؂���K�U��=k{�LcF���)��Idᦿ�_�Jy�����d��iN"����#�,^F"��.P�P�����9���})��ւ}�?�T��;_O�@0�|&���7cgKD��PD��댜2�.��%`:N���n�@�8�ݘ55{�K�l��߆,��`QJ���ɘV��kF�B��+]�4E�`�8�`�-��a$�$$�.~T������n`-*k���_�il�
�J��j�E�@���tΰ�k�`D�޸`|�͋��s]b��l�Y�<{KZ���G��R{��J�R�{��&����X9��ec#0��(EVЯ2�6�W���X�4����a�?x��F��a�Rq&���U~�R/�HWT� ����~�\�i���C�b$by�K�(OR/�R&UNﵦ���V�g��$;��� �	Z�1p���.�M�{�=[B��4K�	�2�*C� �:g�8�(V�Θ���?�`Ȳ !�IYS��b9�޳u��$U�Ά�X 5np���\3NO�J')��Y|b�d&���΄eFăܡ�KU�J�*�K���$� ��L퓏��q�P�����#�LT2-�����u���Wn#%��~�ҝ��K4��Aa90�].�(k�����
���J찆���r��`�"|��
�l��¶�I�M���qi&�1EmL�>;{a+�toU��G$G����|�B���7@�7�73���<G60\ش,Wӟ��ƨ ���g��!F��b�Te\1B`so��[��1�ؤ�Nz0������ٱ��mՁ�Y}o S�x;�>x��]{ښJM��#(��*�R�����=<Ci��C���)D.��'Gur��X�&�1�?͟#+�V�	�C���Gͨ�	��bA���*�܂<=�$o"���ΟV�����*(�&|�J�.̅��(�j;��[�ěg�c$S V�^o[�g:>��s?\aK�o6I��O�$����ƣ�N���0���x���L�v�+IzT�}}v�$pƢ��H4���VײZ�pR�M�i�]`!4JϬ9/!&��,e���T����c��4��[�(�q���K ��)	��BZõwzF����k��0x*�Y�-J`�B:�$ZBX-8Y�@m�
�6��ޱ*.��٭�I߆�/�&�m@��U~Qc������`O�y��=>���PїkD��}@p�D���1h]{� L�������&ť
�eh�V�}���>![(+�s�WV�O�:CY�,�D
��0��>@�x�?�ɞk�
�|�S�W�-�J(�e`N���f^�v�j���'����d����H��Y�Os���m6h�(����<�*Ջ/T��K"�<j�L�I�қ��sB.���I/E���D*����?�^����X�V�K����Pz�;%��Fn����WѣtX�[n����\<D[Cr�١%��,�M��}$�4e�n�f�v�Q0�{S�NFd#�4������\�1ިV�K!������U��|�k�¬��p��"��Y�5�QJ^�>�:����*�)x�U<0WƿA������,�M���l��c�W��L�(�ϵ��� ��N>K�a��Q4I0�_})& ����Eh��%��Mo�����Xy�!r9�U��l�p��%��6�j�o���d5�mR��̭�On�$���W�t���9䂛l���E�26]�^@���A_8�	�Ի��~���4�]I1�2�~{Ŀ�M�`�[v���v龹���i{�������%p��ڵ�CS��iէM�)���^���BV�4��X.��S��C+WE��bJfizs�A�E��?���#�
��J�gN�y��Ȣ@gWI.���~mp�zqşIVqXV�/�$f�f���٭���[�v��ޯ��Dx7V9+��`�J�>R�Oi�[
C�Q�����ә\$��u.! (@H}�� N}��L����?�J���o'O��nP�m�7�e����)Ef� �LV
��J�mw"�p*hG�\S�׫�'$�E���{�+x��CHzS�2_V��L	'�AT5����8���4�&Z�q���	��\0��Ay������YJ�qB�x�Y-�;���,�������q�!�z�d�j�Z\F��ɀ鐐}�3ߣ�s��ŏ"xE��uSY�?�5��<�U�2���s[�+�T.�z���ȑ����y�)aC'�زS
6�ŵ��cn`g���5�9�&Y-�|P�z�}�v�).9*(sO���U7����*Pw