��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbѪU�g��L��Q܃3ZN/2^䀞\D'��ro6�~E�S�c���Ct�.	�"÷g�ì���@7��Ii#N�GA�Fk���!�G�S��ߊ��v��0��� �B`�p���>����(�|/a�01e����ޗ���?+��#pF���Kr�j����>fj�lѪ�w<|��rX%-�O��}9go�$�|~��q��9�;�Z�to׏�OFG���,N��<��	S��aMSU�Ig��!��7��9_�ww˾���[��]��:�5��2��]�XP�btrqe��/M'�L��-���׸�&ҲY�d@E��9��ٳow�E&�O�*M��",܇M�0A���*�;j�+��w<�ɛ�Wߖ�<��]` y+����*��鉼@"7��l�D��ˬg`C�:�W,����+�!�����e�����,ڳ|��XL4��	l�&�|������Cͼ�#���ʞ�H��eȰ1Cƹ���^�d6�)��}��V�"���=O-dL�1�mU�I�6�$�N4ӵI�R��*.~��`;�j�Ȯ��,��j�3�P�3
k��L�[T\3
��;u�~�L ��?�o��ia��$|!�z�+�@CO%�&i9�(�k~�IX���WF�%OHi$�-�N� ;~j�浄� ԥ��9��%�K4�]*�
)}l�ڎ�6�pasO��~SΉ�UD���@T���\���+��%�ϩ�ڣ���O���L^�˘�ZU���z{�F�Z�n����	�#O�!ɵ)� c/��>��j�]jf,k=5^��$��������f�b����{��>�	�L΀ƚ;_��h�Q7tOv�"�E^���|����Q5i�I�I�@�b�����J��p����1��֖����Е�t?���&�F)}�x)L�W��|�t���g��[���]��ö����])���y]j��'z����N��	Ȗ�b�R�� 9C�����D��l0<�xt�!�lL��g��;�q
��5wW�������s�JC�hj��~�w�⹻Ez�s��.��a�Uw]HP {:�����ȿL��#D�4�xMRU%G,�K����7�'��bA12l�Ӳ0/��J�{jN�˭�9�0�5����,Q�:�[�X����D�	�[�xh��>4��Cu2�3O�h�|�2P{00��|#�v\���0�
,V�}^K��%��.5>���v\��L��b���L����Ţ��n$=�}����2�#��I������#d�!vM��E'xƩ�Q�k��T�M4n�*��۹6��#��t�0ҟ��X;6S������u�g����>��\��6k�z`�4K4�b���V�#�Q�2��7!��<�s���:\�P��