��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7*/�Ⱦ�oP*��bo�O�EoNR4(k�����S5Ɣ?J��K缀+�I&&G���Q�����zK}b��9���+�C�YX�e����?���_�	������x?-NL�CLMa0�dTɒ��0{�i���W�o��p{�?__��I>�t�/��z�RO)��q�qȧ$����i�(N��^�\W� u(�=@=ͺ��*"%S<E�E��r�YY�HPb
�^����S��E�P��62�xk6���xL�\R�
��WS�N߀1����k�{x�d��.�nZ=�Fj^!^�k
����̻<���i=g�\mɁ���UXB��*�yo(D��t�n�5����>s��w���~Y�̍H�P�^��B�S��2�v�Kw4Ő��6��T{��V�Rlx� :��v�����A��몟^"��鯱�?�]���:��m/jt�]p�?�z{���ϩ��]TtȲ& 0rJ��\����Ǎ1��ܻA�幝 �-���wV�E�j�C�I"���q���ߠ�;��c�����M�~N](��0.����]���l��V�?,�K<v�Q���4NÏe.��w���(S���/�X&��7��?r�2�������^ļ����3q��;r���4�t�: ܗ���0���a(e�O���O9g���2�_��<q6�x���#�y��еyEv�I/a�����̢%
�WDb��D�J�c��i���p;� ��L�k
�e�-����+jq�tQr�Uw	)���ǁ]�H�o	j3)����5��
_�R��/*�/��V5�x�4@��-�!�@B����G-��]E2�Fбr\�\�6�����3�Z�y��{�H��6k�-���h"W}�Z�l����P�y�?u5M?�����nKH��ǶpQy�9S���]���S��79�~�s�x�c��%����:�;�`��&m���2|IF��Ig��'.����F��7���,>��>�O^���)F��n�<۱��Ѳ�h*k�Y���R�t��ᘵ�)�q��1��	*h��$
Jً�ez���e@Ÿ�^�{�DWR�Wk`�K]9���2
�c�{���8�d�� ��Eь6 ���� 跦�o�癲T�ԍL�|��ɅT�^=�E(<�h�����琱��[� �q3����cM�C��1� ���)vs��W�7�'�r�����s�U�џ�3 9I�K�l��2�!e� uߍ�߃v0�U�sŒ{;��7nw0�T/77q��������ת�XTy7�g;��	K�1+f{��%�.�$%h��O���d�;KkՒm'���re�2>�;�ҡK�2m��3\�M���-��d�+Q45N�<��eVǣQ�PFU^SąH"�f 2��4V]�;��?�=��_�Aj�q������qLμ�`g�V��o�DPh�7b���#�CZ �ޘ��s�f"\&��V�Nh��ԔV�s�Ž�K���V�9�@Q���� V�H,���|���l�!������3#�&��.��{r�y����Vud�%s���&7�����_o�J#?�o��	��-\�K�Ѵ�!)�Z���j����jϝ@a&�^h�I}�-�b��wY����Io\�Xa۬��i��`�u��y���2�Y�@�9�ȆB,"V8/={�ҋ�6��'�s�B4�� �������757�]�G�R7�7�`��oi����j�y6ƀ Y��sQ��x��������ᇏ�׵;֙���1ě(~�閁���CW�E��y�(�!62����dԯU�;��"F��}�UbpT�ݠ���(1�ȭ%{���G�C��>���6Xp?�2���{c�����3Ul]��v,?���1ܪ>TE9�Q��p%�E��p�V3�p��[OU��{A�����J�kp?ù�2z��
lE`�R�W�����lgC;`ɦ�7O`�ǹ��fu����|�'�?؟<����٤|{�=�N���sA��Y}GO�Z�%y�_I9o!p��rB��"|��a �d�S���ʠ*
�e�-� n�p޻���W�	�>��UC�O
��u+�/g���r�y���!&��Q�Q'��&�*}�"cq�m�I�Uw>ԳB��g��h���b��ؕJ:W�� E�`G�@�����^������|0��H$[+���������{@���6��e��	v�6�.	� qC��A����J"��eK��>�P8���h�_hB@���z�U�:Ҭߖ��qR���^�J�F��z�kx<�^������92�k(挠�6O��A��H��w�.�VgI��;�]����N��ba�_8;%h�5�3���t�3.x����.:�7��*ؠY�*2�]x3I�qNݳ ��~������b��Yp��S�wl�I�cEגN��>,��⩡=mi"����Jk(a��#�Y�!>u4���I�V�qE����U;��e1r����OM���� ��\�Ⰹ�2�;��ծ7�F%9o!���4r�r xH�
���Q�E�x\��R�P�nfz�́<��Xs%���
��'c�*���W��o�qJ�߻6 ���U\>���f�ێcv�!E�����&��!Q��mI��f :F�]�zKW�s����h�e��@i����<b,�?�g)rT�7 ��jCנȨ��
	$
!�I�꺑Ⴑ��=nv>��W��V������ �s�f'�4)o���Ca �oC�)[�
Һ5CWS�b�y��֮I�} �u�d���V��확��v�A���F���F����`"��w�
�{$��窤�_b~uD�9�7V���Y��BO-{v�7�uF���o�FM�U�ήjV{�M��6[|�g5��� ���+�T�'��^gc��/�LO7�,�6����ř$M�	�
�8	�������t�������{��<F�F��Z;u��4�_�����A�`:��a��m��B�Rߏ��+B�LB=�ػ��( ��E�"S�W�C�h.�<��{�ǜSV6��i,n0�IZ�?����]Y�b���|:�ozu}�&^$CP��_"jڂ�#�.���P��VQ����2q%Y.J׈�`�g�ʇ�.l��i�=�:Ŭ�_��
���Ts�\ި��T���̥z���m-'�i���'�F�/�w�~O�����=�h�r2�QՌ�\���i���O'6��E`��.�/��c�\;�U�՘}C���e������Jf),�b;X���M��I�`��y�cNٌ��ۿ���چ-g,���/7�/���+�[M$ô� �L����{*�i����n��k���r��jSCWO�L'{�����'�_ۋ}���ڊ�|!ӿ�S�H��Lj�шy�%�"A���-=��~����OL�\��͉ޙ\���Ġ�J�:r��l�Ӌ߄|)���F�Z���Ud�J�����#�8�,���%����l�����K(Ml|�X""�/P���JH�C��{9bY���B�
8������*��g�C؊ӟ@&�x
�]��՝fg�)����`�S����!��?�m���yV	vۥ�%�T~�L��иT�h#����}"�ۧ�^C������]@�,J��S�
{�j�f����U�Q&����|[�<z�^X7�1�lOӞ�{�%~��B�{��p>gm񢴿�ol���k� t pi��t��o'�d��hl�Mʯ)�8�7��6r�_�/w���G5RY�Y�p���e!�Q����B�������7^^�����h>"z��1<����<55��j"�}�b�� �i��c������������B,�':��ܱs�g�x��~������1%�!�<x)ſ��c�^�V��Ѣo�����䱵nc�G�t�&AZw� N�@
��AA�K�����oLYXj+q�d@��"d<X��*zp7t�˕>Qi�٪3'D�7ɝ=1L 0������wvIU�-��^	`X<��tE�EU��Ys��|(� �lz.&��$�P�Xe��k�CߊMc������j���Ro�D���W�.�HQ��,C��3a�r�� v��;��͵���rV�>�����
�mSń����9�{���:��E./f� ��6�/�(���I\.�*`Hw� �,Ha����q�$ryZ]\��~��:۬��=%2����m��O�3.BB���b��u�B��X��u;QT4�):p�aPIk�۱܊��sj���Q d���1�em�2G����|:�XC��؅��t�ԩGV�5v(�� fU@ߌ&3�c֭d����٠u�p�Q����l�k�WwD�"��7�)�V��@+��N8�FfX�E	�a{���7f�o�WL�+�-����_����n�R�;�����6@�ؓ}R�N��`�w�X<��{�1�Ĥ��v�9|�G��B����Bte�W�ŏ+��^, ��+$'�};m��-9c>�C�.�r���5ġ��`</`�Ƨ���H�w/�ɷ���<,ԇc��&TN|��EN�:�8?�q��Ûg�CZD��=��tL�h�F`��S���{��rW!��
�l �M���kޤ�<���H�Ϻ�V������Ҙ�������\.�xX�3�a!���F	3��	&��\zn�� ����}�vop;P�A�!=W3*lG�#,�擊3R�����6{Dj���|
��n���yg4���W���_U5�`�(P�_�+�]�������sn:f������s�Ԣ񩌹uZ$��[f3�Nt�ޟ���0� u3�u5H��Mo(g:y5��
��g�Tc��z: ��{�?R����y��1I�6���ٵ0¡���������O+�,VI�	���.��[��S���,����ٹ�}Cw81�~"6��?b�gsS��V��ꮽ�|פ�����5��Uq��H+��9�&�<\l�o�n�k�ܵ���䓶>�y\1���������v�ˏ1�&�J����%Nw�'-���(�:jʍ�Ap+�5�K�)�0,;�]J%��UE*�,�3��iX[ഹ�_U�.�
�n�/fI�4��V(���=O؇hh����Õ[��F�Snu��?u,�uIes��C� ��mY$�U��DÊ��&��ƪ�(I�L�r4��V$�M!�x�Y�Z�8B񜐁?�K��8F�r��hV�cd���;��o_��G����8W����G-��8r��~���W`�1�ⲽ��j�O�{ g�ʀP��N�m*Yiwu_�`#:���)��k>�a��b9��飃�Q65�1Xj�Bۚ_g.'�����_���.[�Ak�VG�^:�,^0�P[L�B�{�53�?^�	�a|�O\Gئ�3Sz,{QX�L�nXD���zww�Ͼ`~�Ӈ�s��/cA��+�U�WEޯض~���[w71�6�`�C,J�$��D�x-�j�1Si6j��B��c��*�l]J��&�o��us$�[M��Q�`7��A3��cȖҊ,��E|�&�v��`��T4��ziȔ^L���ǈ�E�D�vo!���tX!�_���ˋe.1t۲����B�s��M�a���n�����7}�S��%ڲ��G��r`r5���<�Sk�:j�܏��/��WY����i��I$���.$�4�� ���E��%�J�ǃy�h����m����b�hѺXk�5���ֿ����B}��h56k
�~����?�@8!��l�&��e�E���S�a����eR�[�����f�U��;_�<n�'9V&�k.Z�Z���:��)JE�~s�:`l]ۿp�?�A�G����G���+�K��a
7��;@�J�E���JP
,��7c�����ZI�Z�P:��+�íQŸMm?���$���`���ݰ���z %�B�Q��9�Z]���!�{}�}�ա�k:us�<�����.�qQ�E��e��F̨2��|�u '�:�~����JH����u���ūZ���O���>��X!�U=�aı/��g��t4����3��O���m�D"{3��f�	�t��.�a���8��î���M�CA*|j���摅�6Wp�J�r��j���Eh��rvQ�����w_j�R垔���g炠, o�.L�J������Y���ϡ˰����3�$��T�ɾ*́�끞_Hz�y֡����!�@m�jJfzX�#V�Hd!���UX�?��\���aT�j�����V��1�m����?�,��U�]��7�Y�|���Z�s̭��-�_����G�_�s�;��Q;���C�� i<�hm��)~YI��V3�fD�'n1���plN�{�i�a3꓉�Sо���b��\���*�.`�T���f�#�9��l��o%B�4�4¬1��V�P~��n4x�
���X쓐�$�x�WT�w�}Og��HgW7�hOp��]�h:�L3�J�;�<�h�qh��=�sҙ�}�5@�ό�{i�?�f�*�}�[L(
��J���"ynڈ]�>�y�R�[��D���N?�0G�AJ�|�b��K�6����/PL��m��#G
�d����s�ꕗ����n����;�ٯ3
4}��^67��6��$۟�0��'3r�_&�$y����8픤>�㹷9�uz#�٦��	��;h1?�5�'x�]�K������gę/�Х���_ɋ�����~S�I :d:�Pg?��2�5f�r��O'M��)�Q���P=
�f|��vG��Q'>� �ψ.i�#s2j�@[��I�&sZBg���M=�ub��ڏ~���}�)I���=�⏂>�d��/�%�F�꫁I^1C�I�O�k��:C�h��lT�Zfj�zR��L�ρG�19����n~�%���}���'��k>a#����������_1�IJ��u��C��V�_d��(@�����XN�x[������ɢ������*ދE؍C�B�X7l<<+z��t�u��T;�+RH��%&�
�^J�[7Y�a.QY͑����oK0��=����0Ӹ��&Q�|9�⺰�b�97G_����:"��v|3:���3���kG|L0������������q%���Ǫ'�N	�c1��1P��.��0-
ڕ۷��z|��,l2�V��]��
����>��E/q���(�ڨu2��=�N�	���w��9m���&�:,�ST���f̃1]����K�
��\�󃇊�z���ho!����:-���fv�*��VI�h�����<6� ���?����vD�쿩���K!suq�n�}�Swu���]��yx���	�4툲ؑi>l`()=�����}�V�2�1� YՋ*2�p�x�X�+Tq��������B��)f�%L}k�wL����]{J����g%Y�g)f��Nfp�`������#��-JY���X9j� "���%<��{����_-`��ϫ�i���#~�.eP�c�����-�lb ���o��q�/:�]d�(#3�o7� Ze:Hd���qB}3�(�siB%l��_47T��KL����{��!�O�m�� ~[������=�o�zXIw��=F�B1pлqZ��Om���'1��<ڤdb�T<�V�Q�X�}ܬ� ���}]�-�a�G����BD��L�W��G�H����>><��F�Lf4�I���>���v=�����Ü���{r�H�呎�z���FkV�C�W A�|d����!n<���|�/��`�֮'1:�-�{��i�x�t- 8s�%���ڿ���2�M�gL�=��p�d���H�\��d��7�yJ�3g�&�:S�x
���%CCf5k�I�ⷳ�N����M@37�I�Ւ�y������[��t:��sG-b��ɬߓ+��6�~�l1w�7�y
�Ŗ��� �߅�%�k�uq{����t�`��I��ukU��[�
�w���e}柅��M}�X4o��!从�1����,l�*�<ݠ��@���B�<��3���]x5�^8���9�ПfW4b����(�k�ʮ���TM%q�3@��;\�#�L��s�:�^�`�hc�6�uj���A�4��)�~��j*q�h�w��@�������"Ɖ,	���0��[g����<��7��o��k��1\�z��t��`[ ��q(5�џ�dI��T�a�ȭ�8d�r^����e,���e��7�`t�Jn�5�|Z��/��<2I*^�� ���Q3pBҊ*�绁�s� '���k��D�a$�b���u=ǽe��K �i9�P���d����9F���Ԩ��:�rS|s �U)�ce�I�h���g�>̓PH`F�����>R�3�	}�0~:���XB+V�h)�YLA]�֝�QUD.�t�d�_�H�<�y���V)A���"q�:<�]�Or�.�f�nWXt5Ӊ�1���!<7������� �V1qԔ�n�]�g�}t���ّN���`|��|��t��g-��P�g�@�|M���x	Z.E���0G�3��NkZk����(�7��H|�*�o��L �@hᥪ>&#�vo/h'V���X~�{yá0�r�ɿc�>��
��h��3(���䖉��?c�f�������OI��č�cت��-�_�"��x���!�AR	��_��o��!�N�_�2>�V[�*�֫�pr����::�9��f��6w3�������2R6�^�~LeQ���}g3Ѕ ,6�;�7�L\؆�H�.WZ�?�"���rϖ��6���ZZd��d�u�>@�����p�8 ��3�p��0ku���v������WW��ޞ�hݒu�[��O�����6���}P~�<��.��ã¼]���F	\���6��mc��O���|��W���e��0Y��d' a8ʀ}W'�zql�=a6�k�v���+������1���6\���}˾s����p�c�I_�f�>7��s�ȿ�0tP��M��,5��u�5�@�sG��BEأ懲���Hr�Hr`�|o���;����㆙PZ[g�9	�1N��_2'�y�T<�Ni�d?�Q7��Eoi����i�H��c�l��CIP������`!պ$���B��n�F�/v8�֑��x1���Ӹ��ĳ;��)QIU�i��sۮ���W�9
R�e<��j�������z�v.E[pD���q�G-x���O��{oӋ�_��������!��|Nu��"�Lw>�j����Z��d��)�]V�Tn�2 �J�m� {[&�oвKg�������V�Cp�r��9��Bx��,B@^��e���<2*�]�U�=�-[�_���2�J��4Y&�O�9Ѭ�w�:�g`ʧ{�`0i����ؓ�B�L:ж}�<�����,�qN����HK�z��Hp�3~#� H�+ه�׀9��پMw�E	T����zؘ����8�2Y���W���Y�?\�����>4�J��X�()Z�V&��g䌗	�[�V�4�$�C�mW�������>il��a�q���Ȅ�/���%�A=E���j����~L��+�J�edʉ��W�'��v�a�z;�Dl����z[�pC��i�a8����M�[RdY���PD��i��NWh8��]�hC�P��o��94���q꿁�Z��OZ�ԯ�&/@����N��ܐX	m�����h�q��+�q���x#����l��rJ�؋rgu�\��
-���lJn[�+DJ�w��s*��|�#�'.>_�K�a����"r���Tw��WNg6�tܜ��JO/�'܌k=�Ɗ��unf��k�+�����h*X��j:N�C��y�n�b�TG�H�Civ�%���-o⟮�W���L^�ث�C�[�u���/�3ٷ�Ѧ�-*���R'%�X��Ͱ������Z���m
o��_�ý=������ál�G��}�ީ	����d��ӑ��A=��?��:�ؐnt\��U }ށ�PO�C�o}�&���n���1���x$K_(2߰84�E:����r z��>�ԁ�Փ�J������%�w��P2`��`�A:���Q�6��VŒ���� \��Oa��n3����=�4�mtcf��zKT�A4�����|�!��qa�׀������Ei�nПq��v�feHr�|	�cO3���qt�f�dQ*�%�����2����H��H���O~�,���Q�i���cu���h*�N�%���
Z !FLj�bW1��E@�)� 8�d=��Wd�g��Z#s����0�K��{ۺ*ڦI�ڈ;0Bp��,h�����#�2V7�JK��L��v�
U����GO�[��v��x�?����76^A2�TpC�edd�L�֚�l�1<�LY�<�K�Rܿnh��9��*v��HM���& ޱ>��l�~����-�z����!�E3��hI�/N�4��CC�+5���b'��v�� �%)���ӹ��=GK�����Ԯ
?+?�C�����#��7vtm��D�u:��"3����"�?c�IH�7�n�o��� R%�3�l��	�~� v��sP��jq�8E��Ee�"�|�/�	.�Z�Yگ���>��f����	a��6}��pt��1O�@�L�2�	��G��oA�o�t��V�{� �:M����(���-Hhҽ�o.a����+LA�k.�/�VbЋՔ�%Vе,����<Z	�f�`p{�V�̫j�Ⱥ����Lc�+�W\