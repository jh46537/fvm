��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�9��.=���`s�r�<���s�0!��k�k*e�x�6�#���:d����U�����Y��0�ہ�	މ�eQ����F��C��>XH�Y��0�tiw�FS�0���n�)�	r�e@y:�Vi�)V��$4�ܝȡ�>�Qyކ�8�i���G�����m�ܘ7��Q�7��F	޽#M�9��>ÔHy ׀�N�e�����K�B}��j��(�?/���a��YW࢓���ڊ�%J#Z��,+���������������蹱{X5m��:/��#���`����;��L6s��a ������͊�(�Gϑ���0��f8����i?��t�-4Y>S���I����8%�aR5���.�|H�.�������7����Tk��x�DXǋ���t{T����-d������a{�\5�f\u��Ŀ:�$����j߻C�U*�b��+�c�y��!b�/ݽ�@��c��-�`M�bD�����gm����>��c�wB���P����ϦR㴹n��;Z� ��K��)�
Z;���}2m^^�m\�o�)�Q�-g����[����χ:��Pg8�ǋ�B�(�'_"�?~��q�=)��j�H�3p��W��\�<���H���h,�4Z��d� �	Po�׬�u+Ѷ/&�y^\�|\��+H��f���'�m��N��_�B#ʋ��$Hђ�%���8���hWG1țy#l�sjا�1r����;t;�#�!�1��o�ݑcc�
}3n�y��Ĭi�~����'��S&6�r�����E|�m_u��RLS�qd��a�,��AW�:1�M@�νE��&�֎>�6���eZ��"���ߛ׊;Nqw��-�jV�@/� �槷ŧYF��=�ه���@=0�ک�t@�5�,��L�( � �#�I��I­�M:��^�������J��c��n�4��?6��ٽ/���3�-�9?��	s{�$�a辒���&��/��Y���C��f�obqc�\I���T�Z�$�	H��E*�#qPP�e�r��Z�e}I!!	�Sf_P�I۫���!1Ր3�j�Է�) r�^
����9Z���2&%!�����e�j�/��s�"S��Z�vĨ��g�<��N�)�M,ʊ����Z�"�Rjx���Υ#�,a\5�̝,�G�,�MA���o�#Wk>]w�I�'SI;U��ڎ�z�V斵<�/m�c+?�^$`���hB�.=/����{�(��,S	[r�7灓���f�:5
{����a��,�J`�B�W�·@��Gˈ��N����A6'o�Z�W�I.WU�ц3������P��!�z��R��%�:n%x�s�Dɷ�"wƓ#4s����NaA��#А��)�2����rťo|�
���&�����{%��G/n���V`T�Bϼ �a啂Ja�*b�*��~�"y��U%�b�|^�'/���Xо��� �\x�DX��3Y����N�4�B�1�Y�.U��8p�5G,8���6�g�TU��o����e�CF�^��'6rG�{1�C~������������]��A��5ɥb����ΰ\�:�[��*���O��+2<�{���'��~���#���Yi������H��f�*�H����n�:�ïV@Ix�y'd�g�gv;,����w`S�m�;o���N��=K�hW� �8�Xc��<�@& ��㓏�M���^�El��_ċ	8�ܯQ+�6�nf�b���]
�yg.Z���\�Y��U���'��SqW�	�x%3�ea���BC��l��/K+~c���b�b���.^Y�������*eR�\x�n��u�������� "'R�4+���`�<Ù<�w������[	�KK>�7������8�'���h�=� ��=���%�J�~z���+Ｖ��h�#ќ��h� i�g�Ҵq�4�C]�@[�p�\u㈛{��W���+���B�H��H>nT	���[nȻ��BJr�o.P�q�� ���8��_���%^�˷f����P���)^s/��q��|*$% B�OOX���7�dR�ѱ��hT��{���'X�*$���/����-���
����1wʿ��cՀ5u�x8�Q��q�UA�S2�3��J���v��M�,>Bi	(�7�>�}x�:U��U��'�	{��U��3����~���X�Tw�h��xo8��א�-�^/`\m�;]�+��r�)���'�!]j�>�p5Ǳ3|�簯ʽ����OW���1���G��-������j�ƃ��(�<Ҿ�h~��Ӗm�yv"I
��� 9�}E���^���;0HEPq*�)�����Ϲ`�`��������S�/'�Hݼ(`Q��W�!K�o2H7BSV�=�{q�(��Sz����GV;������D^���5_xE��5i�H��;[��菻�Y�1;�[�H��]�X���\H����t��ڣ*����Q�����ެ <;G��f���)����(�h⛓��R@�h,�An��!�,Xt���;0���6��ץI?|ђ+��#�}��6G�[�u���eZ3����'�����;��P!��k��E+1�:�9�m�:�
���QYf�M�5O��$�&�L��A�(H��vK�5ݣ!el��A<(E�W`���G�^����̧/�4f��h�"��������͊H�6�ĺ'��*�&`�C)�*��bB�ugu@�r7+dV3��6HoR���̌�}��#%o�U�E[��/���0K��t�%k0���ⵅ{���Va =�J/�;	�_�w����4��c����/�	�ד�Ha+˰n�=��=C�f�������z�����ʏ7�q�k���f��^Tm_5�-4���������5���5&��|��:�s0XS#�7�ɀ|�[pE:�T���)����3�/DP���X�|����հg}�6������[UY���^e�;ߚ��;������b�Ѕ.�¡��e�C�{!7w�FՑ��K�b^�O*Px�o~^��J5�)���r�0�]/T���-[�����{���䗰�n�������!@�;��-��_�UB�ba���q��̆�ѣG�R]�����;r�]�hcD��@�w5o��7)�[4n�SqJ��y;�q�e��v��A��Q�Rp��v�Ó /X�c������V�bw�Q\��MvYt+�Ne�
逯;7Z���:{a[��T�ۄV���F���g��;{���U���=���PY
呮2���f'���I�ygv'�k�Cq��guu@�"f�~l$�M�t��b�y��W�����}��7'
I.]\�_�m��4�@�h��BC�W�
�3
���at KO-7d��'��~ʫ�(��s���Z����I����EY��}� I�1ry����>&�Q����_���0k~���%����bG��#d��c!:29�)�4�>�Qيoֿ#��������.���?���{�"cQiE�(q����P��I�:T��D��3@6������ї�X�gBo�FĶ�߈6�$���I>���@�B��v{rM�s���C�G�L�� ��m��v�)�m�����e�ϯ.n���6�<1L�1�1���Wz��}.G��{&�)�a�h�Nud>\͕Y��S��>�3��m.Hȧ�q�1�����oQ�N*4���6��lb�m-��3�x�:
PA��={PL�v��֙���WY�{�&X?7x�u��d�hj�u�<At�����A��lU�9kJi��/1�7�K��|�X${�Wײ�|��ҍ��$�P�_�~K(\R�(.S<�������1�i?�̎�O��~l�X�/�Z��uʋ:
��B�?1�-U�"���:)��e�۟=V��^�/(|�t&)9����K��W�\���^hT�͂�2��EUA<y3�~5-�.�߫�]=�A]F�z�BD���9I^���Rt�% �_�!�f�j��z$�F�Sq5|F�f?�<��y
)�����۞�ЈB��;�9�"�_������<U=���LY���"�Z�a�8~{�f�P������XA�=��Тz�'-w/�zCSEg^e�"X!����JC�z"�>+��"-.U3�S�@��_|{>�n�&*���oil�z.M�mD�H�&� ]���lP?����tN�yj�����q�dK�<�:�7&�"�)�%�Pn����-d����^�r,"�O
3(\4�T��	�'�)�=|SPlB�/@_$�p�c9������^q�xcݠ�jO�f6d{�}�zM�`�����u��?`Z3��ע���O��1��]q���������_�;��D�Ic5�fN���&w�s�mj� 0��aM��ks����PҎ7�=�4��^��k�V���y���%bC|U�Ju�
w&2���O�s�H�R��%\�	��J~>��3�.k{X�H7�PP�M!E�ڞ_N"w��΢�j^PFޑ�0�$�ҌzVK���K�C�����m14���t�ˁ�����?�?�t T�����8����Zq鶢���d#��*����w}Qo�r�ɓtFŚ:�xsT""|�Z+���*S\��K�X��;Xv��юo��w�QS����6$].��X