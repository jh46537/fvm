��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>����rhhm���%�ñ��\X}"y�GM8�,�eP��:h�Z�{|��L�~�t ,������DN�F�	�:j-��u*�zn���{�h^���C��zlC�Wg1MH����{[�rx&R�+0,@Q:/��ц�?yU��g_b��1���C��M����훅�[�>F�?X�	��ϟ�]w&A���E t��/y[�x�b���튟Y}
�]�w3cGTe�����F;;�A���|-�¤��^�{�w\e�+����"-�v�E�`iӆH��n1��Z���Z"9߸���֦�}Q^�t%��$w��=6�e�C�?'G;n�F� O�9�Y�,Q���X^��"�p�񔺖�3ЄQ���W*�'0J��kq���>|6d$j���V�+�{��Yf[�( ���_��qd�pY�o�4�8h� 
��ɴ884�|�?�!�8��љ��*t� &˷�TX�sx�����|��tTv �x_ +�)|Fd�a`En�gEos�x�anZ�9zyf\�kX�fdBυKJ�(��*��ib����4���ř5ؗ��W-�P�t׆Ͳ��$���6�HJ7�xz�����cӶjQ4���S�Z�~D��}���jƘ��R/����މsB�K;@�]3�j�u�T��8��`�+mkY�4��B"�+�	Z�L��;"v�����9s�4��1>���da�����au�uۮ�����B�ai��J0�J��2V��#�p���)m�O�3#�A�B��0jBAgn	���ƣ�����ݵ�����.Z"x<p���-J����1#�;e��C�����4B8m9h��,�9� ��BjU�����np�-�i6��-��J8�����&�Tꃦz)�,v�l��t��2^ ;��^�lho�����99lH7���I�d�8��? �n�� 5կ�	Ր���J.'w@"d��}E�J�Ώh�HL�w�J��0r��a,�%���0��w\�Ť��X�c��=H?,���טgw��J,S�&��3����{�(�{�*�~Y��/�l��^�\�݋�a�"Ʊ�s�~�Ј����څ�n�wj��t�P�cs���8�+����BW7�17�����A�L���u�E�H���/ٶ^&���pK�)h�O�/���F��;����h՞$M��Bʧ�Wt��^�{�zy�%������i�$U�y��}�x_��T|�Ep�G�[]򚕧�-ВN�@󞞟W�i��I�����������:$ �g ��9X�UTo��4�/,h}�kR������k��	��"+��X;D��I�9��r�o+�z���sA�Z��@R�����͋�.���QP"2��sO���q�J��+԰6ʵpO��r�vr�$��������&D������X��"8˦$���ѿw� �rEO�2� |�e�d�6���#ؖ�g�;q���_K{��Ū��A�3�h�n��
'�tJ�R��x�.�L��}Jh�2����1���S�(��S�i�k?j��~�5����Ŀ�ۛ�t����Ù��d�����*�zT>V�gN����g�TGሬoM�����4c*Ҩ�V�����^Rӕ�"�k�}H S�R�2yͷ��G3z��@�b˿u����oN��@>�ں��ӽa ����/��
b�ǣ�\�,] x"���)��֊v'v-�T͕\h�S��5}xǧ�S5��R/x�h��,Y���Al]�ۜ��'h+�TQ����w����{�$ "qD�n�vh����g���,Oa�}'��Gq��|�\6�|ƍ��ѥ}��<^˸��c	�-X���7��� �e;����]�ĳp?r���"X��K8�>1�;[�8��V�6S$��b�6����Ɯ��H�|��`/T�G�X�s	|'��iy�@�I��c�	�T��b����M��s��/���8�x�ݙ:qK���]�&�����^��2���{�ˠ��.�Hsfe��G1o��V9�\1V2v)�|�u��Ujǡ����b�. >���凊(��w�����P$p�r�/��1�2��f[Q_�gʕ��)���/�P�I]��
��\'y�X!>�C���@q��λ�r�ϾC*z��a�_�W�����Bm�z;2{��x0Xg��v@��g"5؁�c���SP�J��#a���|��^?;&�jj-�oX�l�� "�/���c���Uk�/�v�#�t�!N������(�'�8Qnӿ��wV@)߸z�(�9Vl�����s�������oܙ��3�j`�t�����j� �Ӯ��)��[B�Wk�UWY@}�dƵ���'p"����nL�a[�DJ�������-��O<�� �gx�6 R��G4��������|����>�'=V�s�j C�ԚH^���rt$$�]i9q��)��q��!ƛ��PX�������PO���=*��sE<�$��! Dk]��zw=`i(��!��`f��0�Z��g-��2�Q�sz'T�>nQ>�ś�H珤3����V�*Oα G 
K�n+�ii�'�4aJnڪ�x�E1@;?�?`��-iBdȆ��z�9�m�#}���܄�Ai���įW�H#��f�C�)�U��uo5N�k�TW"#�d��X��q��F��f²W�J9�����T(A� !:\[��{��]1��J��K�x1�m6�#z{d��0/�mfaȅŸ���Ҹs�w)W� Qe6�n1��Ɨ���xNUXMm+zґ'Đ
pdSG��j%$�Q!�֧eG�<��K��v�^�&�61=�j뽂C�S	U�ݷ���t�-�N����Ϙ$�g�<��ğ�Bf�4z��B���`cV)ݥj&g��0sx{�*F[�?��u��!}��}��HZ��ٓǊp*Oh����I8O������х��e�Ҿ�HPX��2μ]$`��H�#A�n�q#�	 ͚�>�)���hu�C�_��ꂦ��������~��7AW�G7+}{I�h҅�2�����`i��f�j�%�{4Mѯ�ҡn3��	6�b��^�v�qm����"�ۓ�	u��&��Ж$~	���OΤ^�:o�
:���[�ΐ<�=�`Қ�O�Ow�YI����(���1�H�6�SD@}fZ���Sy(���|cp���κ�O����,N��;!N[���;�����I/��ޱ�4��-�r3�c2�%;�]g
�kw�k6��!�+���RA��k��i5����_� !��S��09��y�(�!.�&0I�\n7`T���p��=�=��ǻ(8��n6j[�0�$S��]�;=��.�%#v�o[cH�0����$sC��5Q!{�v��E~��|�Lj���y;���9+PI6�����m�f8X,�Ds�[�m�v��-�V"C���m�9p���䝌��ިu�;��������5I<�*�<�d��@��c6}��}����tU�4��7:θ:̎(f��#&���uD<�F)%�~�`����!,a`�V�;l��r�ka>�r��!�}q"�4��{Z�Vp���c I
^��7��S�bG�0�@��G$��O�Y8��O}M�	�7�VEћ�q�}���oˀ��v�]������	o�ŇJM���<;\굷���qzx1a%��i95���n�H�C��bo��	��I��eG�h҃�@r��7�<,�8�D����	�֣��U�r
�%���ܳb���������{�NF,CY�a��%Q��G�hٳQ��������9�����%���vӬ��B�L���!t�4�������|�D<�e7½!l��^^׶0"���}�z���.�ٳ����t,��.�ʃ�&�Z�D�O;���S�<���X�7�_��vD�_�t.��'sE�\�$WC�� 1�S
̔N�����ǯ�&(Tx2��E�d��`�-w��(N������q"���g� /4�M�>�r�H6B��%�8��"��AzǱ�L�-ų0w�zy��K����О��'����Z0ݗI�}_n�zu�Μ���9�6
_�}��qx*�0[��i�B�3����Դ�<#�)�Q�#oc��0��.�}� ���r��1�)�k��m\�����~��E!{8RZ�98q�,���6�W���b�(��ۊg��>��줡�K��	����PCi�)�Y0u]@kԬ������|+sں=��QV�icZS*�6:�o��<A^�J�7�ǿB��d�!L�:�����O�FȚ
�ºtʱx��E qD)�`g8����ܓ��'��cT��i%���
Z�l+�i"s�2�S��7��%V�ECC�av�+�ӯ:���y2<zi�B�]�
��d���~�hY���������L�eg)��6�ؤ���G��Ь��"~2������0LNb_�5��3�;�T�w&�{/=�T�g���o&(&~+󗅐?-���û&^�:�[4�R���q�,���o(Tj��B�띇�iZ�4P+��Z:	?QrSV�u[3�k�i��)�|����}0mU�[����%|rs|����uE��������|k�\I��ι�թR?}Ho�~�.�ƿ��x)�鏳��@�-\�2Z!�]�{��%��!0��;g���8S�|跸�)�NF�r"�<�o�l5������?��*O����
�V���R���^b�rT����6��d�>3X�q�ܝ���7X88��>@��f���0%H��v�?�);�����/�h�m�^7�:�U����E9B7O�+N�0�jT�ʒ�*�E�I�]Ax#`�VI#�rt����VE)4��4�G������N�˘�"K|6�ü>�O|*�p� u�n� ɟ�
�Ȇ�88��QT����kY]�.dY�="Ův����6���l��i�.:��5p4;L~�y���S�t o0�y�:�#��i(?��i�ef���gP	�a,3
Ls/��E�1��I�����^���;R���Zb�6_�Ʊh������RX�KF�%j��#���	Q�0̑�m���4�+�I݅S9�8�$����|ĉz��?�u����Mr6�=�+b�\�[�Gr5=���i���POE�Y�~2e��d�w{0d�֢��V��6�k�t�DD^�AL\h��Gɋ_�|c��%x�
�Ȏ����):�͏1�M�P73rv<�|���o��ԋsE=��k	5E2޽Q�!Q������?�3�.�g��>�zɾѐf�<L
P�;š���ͦ	���9���H�1�V]n8Χ����Wi��T�m W\9��� �I0~�������Œ?T�?�e�]�H'�r��d��!0��=����O�}��_5w<ʚ ��"XdR�P���iA�QYid��׬a(��w���~:�]8rb�J��L�WQ3�^�V/q�Ag�:M3=R<-p ��[��m�$/�m��`Û)������������o#��Z`��G-���� ��$�"��D��:�]�y/_�!��_���_L]�	0������T�Pbs������j�~�yl��V�tP�ߦ��wj`ޒ��|���%bz�ax�������(`�M�v�e^x����ˍց$�a��~7����*�q.c���l�͝�0���n�{%6����t���)@&����GiG��OH1�~��E��Y���E�L*��[�%�q�	F *C�@�����̲E�`�4����,�M�ΊTopA;
B�$���P�x�b��գ�z�kc�XR��(�S�X��%�h6�i��h�vl��/Z%_�@I�B�L��+��(R�/��ci����y��VT W�q�!��l)�z&O��������V�);�aT����\��J�T� <A�!^R�L|TGăx����Q �l��۶ l��7_���M�Tǰ:EĎ�vh%L�1E�8K/IPS®����Ӝ�h(�"��1��FĔ�����9�§�"����e��#C��i [�u0�\��Fc��a�]�8`V`�ғI�~F�����_�2������HZ�J7g��h'] ¥Q��k=2d\t��>��,�ֆ��xX��ͦ����������a�{�nN.ّ�<'Rg���%�?�l�4��C]�,�NW�k�F�S}����H������iKx������xe^-�7������&��b�oU����������cP��:(����K��P�YU�#|<~����gk"�Cd���YQX@��<�r��
ƹvv���2�W4����g�����D�*���4�\򻼽�E�Ж���e��V��0Hy�����C
)�@ޓ}QCC+-�1`X�dA�����_S�e�,�-9�I�k�屙4I6	�o��0�2H�*o]@��ׅ&������9���G��[��|_I-��"˝8���o�E��Y���t�%��2�X�]5������-C+�A��p��+K�;Ly
l��Z-J���ٜ b��[ �-�@��%h��|��y,�6�n�R$kS	r���K�v�m��'���(q
B#Ms�'�E�������ԂVt�F{{p�F��8l�K�� ��7|{��r�z۷�h	&oJ_s����^���.;cb"$)��qp����n���3�cB������c%G%���rhj�3�w���&�R`�y�� gP���ʚX�	��EcM�w�w>���C��WDPY�*�w�/Fu��ᔶX^�º���e���!'�W��{<�{���p�I$+�)��9�EL�뤛6=`2�(�hK�i���<������>����$_�`�k��]ˇ��gkV-^x/HA�z�g
�
�`A���Ɯ*��z�L�r�Oa��PN]E�2�x�uq���h�oM+���o�+4���";�gVw!�oKIGi��Z�`M@@N�R�μ:�����W�o�{�m�݅$��]�_"��B�壳�U�O�v�@HX��;.r���D�$ػ��؋�vÐM��zT�0&�f���F'/��o=z2^�r)�� �kM���X���Vem�ſ�_:��c�����Z|h��n�DIC�k�v	g���s]�C^�?Ν�*���:��~-hg1C�Q��n��ܙ�w汥�'v�x���l�dO�'�8&g^պz�e�0D��F�ʐ��9@���۳��rnuEAB#Rb���� �TW	��X��ߘ�w	�������!�Miǡ�a�\UvV1k�xx��>Jx==#��h`\��s� mf�
d���F��ͭHp�'JS�G;x~����H��\4}���p&S4��-Ԩ���D�t��+	���~�7���!MWjG�2�q�S��Rr�OmDa��`	ő��"aH��Z)<�2QfmǂW�uӗAL?�r�`�;!8Fi���
cm��/ܦ�
�+M�!�ZIѠ�W��[sjnf�3ϯ�G��\��p�_��� 
sv�hmr� F�x��PҬ��e�f6����^��[���S?o4� �D/���W�l�(�=�@����!�\��'~9س��7�p�Ь����'� P��U}烽%�j���RKX���MD���v����:�M���p(������Õ�UV�l���a/����\�$)� ?2/���
���%��c�-�ҋ�^.�֊ٺ�P_h�ϟ��zj}'�
g���m����A<eE�_g��*H��Ko����Bu��BHgv	�B�٘��2$����|I�"���o�(���g���&���J�fk�A��>~��W�UUV쩇�u��&����)�>��>����<l*Sj9˷��sٺ�|��{����oOM��&	зyV��Ki�IX�q� �u������f�r���Nj����k2�چ[�R?#���*#�q��l!��<j�������AꞆ�Ŝ|��ꅵQY�"H�"��ۯ�����UDT�V��oe�mn)2�/ڂ�P$0{�bf�5퀢ME<D�fN.S��g��z��� ?O�+��P�*4���Րf����B5t\9�]I���u��5f���7��BĠX�
��d[�\#W8��o\10�ޠ�#k�1hD+<�qx�#I���8}g��c�m�"�a'˴#8@'�ok�1J�g���L(7��wK�M���V񒻳\�vL��A�Hh����!���$�GJ ����&��UY� .�=j��2����w0ک^7@��D�߁&p�C�"�r��k�f���'��O�Xi ����74��Z�xW4ګ��E�k���9v�c{�`%!��'6�E6$o�Bj�t���mg�;���o�]i�<f�L܊�TT�(d*��]�`�:�ꛦz��;�D\t����Ӵv��Nv1�n�kT��8k�F��3W.$��s�=D2_������~o��p1�h&�8g�k��j
��ÆEISd��	�M�$@��#�d��$�5u.��j�V`f�GS�Q���N���"�W�tw���cN]�S���/ʆdp#g&�*;�`��U���=�@�Va��jޱ��a�o���kqu�6b��um������ԞR�������R�����R�#GlҖk��~�������"�y�}~��ɇ�	���}��;�/Bc��y���^Qz��Ր� M�{G���/�џ[��0�ң��-EH��ݎ=��q��H�췜D�(�8�W�/�U��\ʗ��7.���c�j�*%�a��g�C�KGT�K���t�E�t����]7�[ݜ�����߉hpN]��R�a)��J*0x�7�0aV��1���/�A��^`L�]yk�Iz̆<3�Ĳr���l'��>s�Ĕ�=�&=�&k
>ى�J�"â�h����'�0$���m��N�1���F:D���Lx8��^ �\��۔EA�gF����u�T��sb{|Tay5ʘl�h�9)�n�)�5���a��$� �2Jl# V���H�^�G�܃k��i�2���`� *�*�K0!m��^�GB���T�J~��W:�0�4o_��e^���'�Aߤ���-�RD�K7g4��L�~�Z��+.�����:�cU���l�,՞�[5�`cq��8�d7L�/������~�A��������:������Ov�U�;4G�, �I%��*�V��8sb��#�W!���K�Ubcؐ,��v�Z�6���.N�.�����y�dx�r}^�l�E�U|j��>��
n}�tyQ��."��ؐ��C*���]G�;�M"%�C�>14��S��Lp���0[��Kv+Л�Ɖk�?r<M��ӭy�nf<�*�ҷ���q�'��%,��,���>���z�5>-�K�/����r��eh��+}1k�ƴ�&pn�g���g.e�JJK����`���L;L��KKmk�����C��%�9�NTUN�������'�˦�9�ǈʝH 2�Ư�Z����q�ކE�e��#2%�+.Qс(AH�
D��;r�RG�j��T����X��^�}���} ����{�z�h�,��'\�(���~��mg��������� g���p!̙�K`��Ru�~ʞL��2#UO� �uo�r��I檝f��
Ս�o�%':��p �<����,�k�Y�zǻ� ���,�޸���.g-֦����Tf��j���
�|N1��{��Ad5o�;��	4�4<�$�U�"�x��t��ꎵKq�P�pg� V��ę��o�v���Ϋq�`pM@��Dޅ�J L坜�Ap74�L���>��K)k���v#͆�Ic���۳�`�|��P_7>#�mo���_�,ȲL������I�SJ'�eۄ��\59�\{UL��;��}�O���DX�:����a�K�}d��>�����d�U�vb�YZ�{[S�/�		��_} &&Ƽ�U�^�$ke�d^�D^����[��X
b |����{f�������t�aR�c\hc���9V���ʏ&�J�_�0_M:��Ȣ@�e��px�����#�����Jal�k��EēK���R�(f���d���J�&1@����{����*EBL�QA���|Tq]ܘ�xe�o�����C��Pw#�g�lΆߺ�o�IR<um��[�>#u�,�%�Z���Z�g�� ɠ�>�^+�+臿��h���YA�������ܲ����De�%�og����\��ϘYÚ>�`">̛ZI��v��L{�i�����9�]q8뼅�`�j��Z���Q�����Mgt:R��!{��r�:���t6ξ�ʧ\��	䢅�'b��@:>WL�r��n��(�:h�Hx��Qf�����-C����)�e�M�G�EnQ��[R�]՗���D�gL��	`9�-�r�i#��&��ׂel�e�p7Si�oְ�l]��.���S�8Q>��� �sj*��|��CD��fI��R��F�*wu�C�������F>7����K�j��%D���ڱq��:�3g';  2��;�Ï�td���ޑ�
��%n�bA�03�B�("�x��6��c����#�������hM��ɬ����+�S�E�.H*A�2O�v�;ER
oi�fE7��ςq �e=���'6y�#�Fkg�Z�qS�!@�6��}�Q3�ۻ�l��&<9�q����<1�
r��Z>T�Fagn1��^����0�+������-b6Oꌓmi� ?�M�&��o��<��x��n���j����>��,C�{C��7���?A����K<s0�O�z��|��~Q��
ʇ~��ѺBw�Zy�=� ���:�0Sa�Enutϼ�ŵ�A�k\�:�`,r��s�KD	��-<�6T�I�&�*!�"��eJB2�.���)�^z�u_[���?.4����d��N�,3��N	נƠʎ�}�ǃ���܊P�Ia~��Z���NϺ�ө���b �̸�/^܇8s���$�e�� B�*\2�V�|�[��ǧ7�a���ߠ�I�6��&2�	��)$+��"�`@Gt�a ����3P�w�'��]��"���+?`��a�@����EY��*sy]����݁����Z��b6���w��7� �W�<'p�6mH���^�p�|W��$%�￝��!~�4��K�Ѫ����b��=�[���mP�Ȱ6�^�qCߍ�Oa[R�r���*(o���.��WP�n����I�����{�.��~:��|dR0�s�_�)��iC��1�/�ޞg�m��Lۉ������)��-O�%���$�(��]��NK|8��{_{�dO�ķ�+B���.n0���gyrh |��5 ���Rq��I�ݦ����c��n��f�.8�g=���ˑ�Ds�"c̉�q�ֿAT��+_��q��Z;P u�+��=��`����,<����q��f���Q^�"=�Ú)�}�na��?d���K�Cs"Ɲ6�>S�~����W��˗��8�8��}�(xmB6����(X-J'�=����PUE�1� ��Q�z-�� ��Z3(��4�{aN�J$�Q0���}�cH`�C*aW�_��i��VPH5+Ӎ?�߾��T�QՍx+\�T!u�x��̺�R�>T��H�V�-�÷{�EZ2��"�WJ�
��W�G�{��MB�	Z�x���v�U�W�h��!7���6�gG�Yg�[xMz�����������<��&k������(��?I��屈��T�;�Ӌ/���x�c�Q- �j���)9s��
�'�c.�a.��UXP*H�]I=Z����У[ NW|�$#�'L�G�p�΅w������À��ɸg�s���u,Q��ʦ�p(�?��
��&����L�� ��,�C]�T�ϤC4��?m�?%ǡ��+�����AZd�ԉu��*�
F�؄�g��ܼ� �����.%�|"�]=��@������^Ky]܍l��R��z�E	�"��L�43�2O
E����4Z`N�$,������T::�����!�P��}d]�� ���Z�P_
�>m.���pU<Va(�oJ�x�.�EDU�W���2��H���HhU N�Újj��sX����B��q�3��.�-��O'0�3��D:p�搓˒(#�]x�wX�w�o�h�3f�۾��_4nZ0<��B�寣�k���Rj"���%d �\�[y�^o<=�T���ͳ.�#���$�s�Jp���)]RlH$�~��_(��T=�J�H[8�Mm5Dj�ŰbV�2H��٘�@lQ����l&F�n݂�u���7UJ�	-�µw~�K�~%������oajL Be��c��;גJqw4�e@֠]��8 k���!o�?����C��B��:>��1J�9G��Â���Z�?��S͙ʹv��O ���u
% �qsz��v��_x�>�n~�"Y�h��7�&��.��0��O��~-0�BXY#9��]��\��Ә׃N�S��X�c�P�[~M���O��va��V��d�(&)�]���;��2�5Oa��q�jx(�Oz�QX���T��0���h�ub{8o�&tCWq��Ӫ�
���n5�QP�f�sൈ��N���E���Vn��/�+�i��>/>���Eә����K_k��15��	��4.�H�v�
[A=�b#Y�<f)4f�Q5��@���K�-h;[*�SD���WDg),��f�>+X,�\㪽�O�ǇcG�Kn�R�O���C��d6b�����@���j�9�����&dT����9�1f�������6��d��y����^XU�FA�G�i�Y�P��],��`B}�Q��a�?���K�3���2�E�޵Z��� ����j&h����eڝ����j]c^�wd}%��{���z+�F�c,�M>����k\�G.�x��E:�7�ekw���k�ݲA��{�dumY$���|ҥ]9S��`�:�oh��9���s��z>L�*z���l�*+]8ق`G9~3��*��^A�oj����g�W�\����w0�N?��W���<P5���M?�B\����Ko�6��M�q�?��V�+�858�1t�
NΏ`�?�g���ֺ�_S27l�Ɉ����1׾�aD�~$�����`��GR��5M�:=N���u��\� a�[���+��x�(5��}F�������J��οPc��x)3��Ȉ��@22iW��+տ���Ei�����zw��Q(L����T�V�2��ZZ��^ʸ�ȣ��8��b�B1��p̌�K��6ӫ�6#�.]3�O�"�8��@-LH��Ή �m3���e��`�"l�����Z:��e�Zw�"[�#e@�#�v'���X3Z�Ө8�x���P&�Vq�,Q��{10��`�]�R�YΤ �`H�>f ��̳���|}}t#r҂e����G���Z�W��J�.>qs^a�}�]��
��?K.�ᑚ�;D��b�&*��z��dMMK##~�y�	Ѷ^���0��$7U�"�F���g��ʽ�p�g���?���h�P�$w�r��/�����T2$ҙ,�Ȅ��m�(s�1�Pw�%��8[���=f��� ��K��/z2��]�%� vHⶽ2���M��>'cZq�۳�|���s�އ��"CQ18��Ò_���F�&r�̅vw�"��.��@��:�Cѻ���wsG5F��c��Z�Η��GbwtZ�˄*$�'�cb�Zlư¾ǩ���h�rY0��X��+��R���+ٔ?�q�Q�"^s����'�F��߄/w�"?�ޘ7�E��#�'�2�i�gY�|���.!�-q�cu�=0[�3<����%�ڛ��*�E�TɈ��P����Jb���=KU)_�ʺ�O�d��.	ċY5 ��*�,L�z%��BiN�te�qg���\4ds�.WH"9v�-.����Q��̏�� �p�e��<Օ�YJ�D��u�	��//��Nk��5��2l�c2���Cy�9;��p��+��NV\�~��sL�M���3bG�������mz¸Bo�r����NC�>#H��5��E��w�3��a<X���}X>��D��Ɖ�00�Ǽ���$���)�~�(/`R���=@*U�������#�xaN�:�ɞ���gG'Q���T��|�PS':U���m���j4lJb��]}M:�H�  \E�TkRAm ��$�H�Z-�����r�F
bQ�B<��;�!�� 9ȝ�o�¿]ח�!^q�"��(�?	3k�gP���_�,��f��+ؽu�)&����x{�:;����U�hL��o+�`��C.�޸��Ȏ�cRr�����F�+���l����P$p��1���FD�;���ӟ��4�P�8���3ՉT{�{Ȃ�v�1~n��oB�'���sŰ���1��;	��w�*�Oӎ�:�Jr�`D[_�%�����	�P�'D}��d��*y��'�<Y��FlyT�*�`s�σ��%�]�m��r- ih�j"H�6fg��R��A�-� �8���_^'̠�,�TS��kB�D�1e�� �u.ru���4����PY�U�G�~�5�d�)���8�\�|���M�Y����E�*@��؇7l���yL��>��N:ӈ��5x�=t`�����.�j��,��ᒼ�K4�xက[�vnܹ��͚%����V$*��Mt��tz�����
�J�YĻ��v'�������6́=�k���|���+�����V�L���Q��D�֎l-�Բ��84�M��%{y��Md6��K��q��Sm|��띌؎�o��F�T��ϵ�]���5�dB"��gX��_Q���f�.x�0m�E,�;��>�>�kq��ʝ�,����+K�Ȋ;���h�e��-��@a�iu\5p�
�"X�'���V�⢊g`}��]2j}��J�����Jџ�t�,d%7�ޯ���-�x�Xd�+߆�"@"��Ee�IuD�Ro���4wL�1�L�6q���c`�~܁�̦}��ǵW�9�$���L��j@~�B�l|��a5~���#g��!���ƒS���l�兀&�	hs,�|���guK
<��p'�'�n�Vk�������~�T`���&4��	9m�.!�L��"3��!���[
<���l

�B���~��ب��� ����:���ޟ��><�-��-�	���kf����*H�� �B�%�+�y����@���}�T ��
Lzv��7��e�#[��ԐO��j��m��tc��8T�Ιe)�z"�)m�>�a�ZQ�`��+�Fy�Prf
ȵ�[��I?+��e�qc:K�#�k��-mi6���#�	1[qve{�G�\�㓐]'A�eYCʐ�=��%�E��_���EeL>��58�ۧ>"|.N�6Dk�_GC���X��/��� � ��F�(Z�{0�
	p�t �K~sO��><F��)]3I7Ĵ�-WHOv᧚{�ݷ����O�,a�0ǰ]��}֝�B`M��1p2���{Ͱ L��,!�Uv�pz8_9{�>D&��Ͼ���?�����d�dU饴gF�cNYP�^���8��^�R� kN���YA�5�ڸ)^+��Y�V�� 9�T}R��î��=��S5K:��S�H����RB[�>އhSRwHNI�(G��A�Wθ�̋ÞO��
N�3MW�J<z�~�(\=�-&��2�A�R�U��x���`Sa��N'�*�J�e�^�z��6���G��T/t�N���G;4�jHǴ[@�U���R�ҥ�|ݕ�(��w�I�i��jT�0cY\��6��_E����R���s�Ѵ�G�b!�CM%�y��:�I�(����߫�����+Q�8Z
Z�(o4��a]�J�n|���p����e�Q���
hQ&������[�7P{�4�̤��ˑd �tY,�=�5*������n"V�sd�	��<���ip�]F ��OA��xP�s�}y�N�X�t�C�B����>�z�殗�Dc����#ڊ�#�3��s+�.#;��9 `���(5�^��o�s�� ���w Y�=������jF���Ζ�f6Ӛq��1H��Puf�����A����r��^*��ރ�����9��Q{�6��8k����:�LU��K<�1�Z�jZ/[�4@�C/�IYKҒ�C�c�$5��C��3�X� �=<�	��)v�_��{�>��O��{A��v�A�Q3����o�����V�j�}
�%�XtvXƫVe��!�x��:r�Fp�b�W��EH��x�'Ԇ����ִ�t�Ĉ���#�Rl���@����Ee�	�i7�=�� � �Ceb|#~0z"�Y�:��mu�>�t�W%�3�Xv�ӰU�K��
>i�E_���Pڱ��=s�z���`�;O!w����+�$��1��W���['�%Ə��6�'-?c]c��t�%�2�A��C����!�>����ԫy��7P�]��E�I7�3C�+�r��1P���+��CB)�ʡƋ-EaSr��^�JӋ�1]r���0|PC�aH�������e�n�*��*o8t�|! O�Z�U��㭁�R1�kB�����>��]F�}.8���m���Oc��+�v ��e�?Ll����Rz�]>�]���?�����Q[�;�Q|"~UP�B��_���E�`B���n�6=�?ޛ�q����O�_��H�)|��]1��:a=1�v��)��b��F��C����d�W�b���"7���2���lo�Jm������7\�kլ�	e��Ǔz�ٹ��Ko2��8;�ͯ����Q\��GS g�NB�����"%	�g��S]��aD�����+�#�,a�*L$2��z��seE8�#0��)mಬ�?�'}�H0��M2��;Y
��%����b��T'ז#~����7FV��
�= ��^~<�[T���9�g��B�(�}�����_}dK��� n�2Q�[q�)�,��4Ԋ��a�8��Z;���:�@���KӴE�!o��LHKI�XV���tO}.>�c���.i�~a�M�|�>&��R���ef*���{OF�2��o�Y��1�=�,��*��_�An%ALT@����xnw6e9h����s�D��;j��=��!��\��P�B?e��lv�L�b���w����nOSL2���{#鋱��A �vc[�pz�e�Pđ^
�X�U�-�8;�Gp�G���XNk�5G�p�Vڜ�\�8�{�%����q	k�B�����ɓ��ks�|�<����}�mt���HK���t���`����c����}�(�	l�^��-��V!o�3�/������U��;o��Uq+F#��z#��96Y�_���8��~7_-���	(�p�flv�$_�ӵ9���HZ�s��>RYQ��Z.+��s��\W�x��yzW���Q0Z��8]d��{����2�.�u�-��.>�w�`*�a��6�p�S0�n���3=�2�Թ��_M� m���SY��z�N��:�b��Z�}�iꅣWXFF�P�]�6��7���+ �"/B����V�����x�^J �Iϸ�<������iS���i�T��.�I�����ӂ���M�'�Ukh'��żڱ:_�(�@���b���s�V֭�֊���j@D7��!ڎԩ�l�{�����>Uٞ���wT���D�f�b��!��"�i}���$}G.�΃uA9�4�fR�旾�=�Y�~��c�%|��$���XE2+��&�������j[���V<3mÊl�o2�Mqz�Ѹ�:���|���+�㧗�R�둍^�!x"�����x����N���}�f����/dT�w}���^m>����)���<�:�b���֗�yl�ꂠ��T����&�N	��M��2X9��rs�~���A7�c}aoѡ�y�����;�e�UǾ�n�1�
�7JN�]����D��XA�V��iJ
��[Nz���T-�UNP���C<X��Wƴlתyi���L�_f�����|���^K����`HM��%�)���Z�7!{�F�BLc2S�3<�} )�Ϻ���ǆo�.K����S����a!���/?���_I��c�v�KS�is?��Ұ��g����a��c�F��<~���9�g�n�&#P�!�t�A"<+7��WX���4R��J���|�=t��B�}.(�4���^{�%���a#�>�
]�î�/~� �y4�B't_��d���O��N�j��0����|qV�}[7�f՗\pC�w��s�r�[���IK`=�� |��Zϯ��5EϜ��y�t��s񊧔<
V"޵��6Vl�)yD�������*T��\-��s2 ��7�1)����:���2<e
0f`(t*K�I�㽭�m��l/䀊5j�t��z�l��wc�q�������A$���\�t�[�b��ؙ��=�����]�����` l�n]�,|e���ׇ��E�M��'�2K�üli-��+wh0'@+ڬ�@�HBŔ��y�@�w'�;�X(+^d)9G�S��$ٻ8n8��R��w���1#ʽ�$����C�!a�5�s�	�����d�<,[��i�_�T$M�{���h8�$O����ځ�]<8^���:T��p�+8���x"���;��[k(�~UYg�x���'Gu^uv�o�Q�t����	
�m�Oz���:eTB́��j�Jm�ڪ�bO����{,��F�J�7���d����2�����=#>�]��sA��g��s���C[1�N�a�]�%�	��!%�l?�j⾷�m�ł�W�ܾ�����Oo�*i0�k�0�ɂ�$�N�Bx�&��%���/�c�3��Z��銾�FW�-�F��=�V'uu:x��,���y�^��Q���8��"��Jx�Eq̶�m��Ա���6[�U�K��Ca�@1w�}��k�M*/Qz�2G���\7G��!��R���p�����J������	y�XR�heH{�/4J��&�����L�p�S�˵��
�<I=O�OQX�^Bv?�(G7k�|�[�[����� �ODW��W�7��>�*�ޖ��ˠ�ŲoSa�}(��p��|g
j\�|LF�e�B#�?�h�Y��w��/\�f�<�G��S�hlЭ��.-�����}P��|���{�*�F��?i8�+��t{�yt���:��<�
4�5�9Q �����>���l�I@,S�2�,�wٷN�A���K�D3��A��(5�ͼ#Ǫ.�F����Ȑ��rX[�/�/��>֛51�LZ�RlV���&:�����ՔM�n����	���2�1��\/�c��c�a?��됃���d0���9_���	�J��FU���&�!z��b%�v,F;�G�IT��K4��4,@���f,&��4'����[���- ���<�U�iz�i뽉�1���<;k�g��	o���~�x��mi��Y�[n����\Gr�l2��^�w>$e���2��[}�D�����'��m���Q&���?��&ZnOD�e�
�@H������ɶ�Vq݋���W��;E��AH+z���2������]֚b��f+&�i��M��+�J���1K�1?�{�A5L,7����F�r0��
M��=�Q��jWU�Trkb������&Yz�9��Z[u��,��YG�b��m�lo�x���1�uQn��@��v� ����k)堿�!��@؈�)gV��,ab)���ȁ�l�uC?�J�x�Q�|�*'X�l	�!u�)i0[�~�y�<�M:��у�!oW��^��pbK�	|�巂�!\������`u������,����YS�Dh���pZ0�}��o�&� ��o�P��a ݺ�D3D��	ks焖:�ٛE��¨	7��u��ؓy<["�y8���=����`!�w�:y�̽o4���1��fLc�=��f��V��u�Я�r~�{����߲�{�����-�:�$o�A̡��M��:�AN4ʍ�ӂ�"�D�x�W�p*�ъ� �O�p=�,{�M/�;)G'0��ֽ�s;��>N�X�~f�F)�CJ�7m"�?-y��[��l8��$�E�i�ىA�~\��bN)��|�m_C�ZO�'lV����0��cD�+��}ؕ92Ѧ���%F��9��n�7Dh%SBf�6�B�0�]�Z�.3oY����B+�n��쒕0�G�ر��ʞ��J�q߼�Q\DZ�g�U�٭n��Hx:��S90�� `����K[w=�˴bt]��Yy���uɉ��� �<�7^�Ǭ �9!a�"�J��s_-�{�Z�<�j����|�Sj0�����]Ԛ������k��2��G{j���ij�&�@�En���7}=����}%k���b"�M5	ˁ���'����n"t*�28���}$�����â�%\:��N>/\�rUF�I�����	���S��XY�	��َ>Г����*Wp�c���ݰv�B�F<Ҥ�b��Ң��E X�Xe�{�O�\Q���i�0.����>�{U� �gGb��7r����~J]{�h�Y_�Q�s7� �����R�����9�Nƞ�'��)�����,�wٙ<ג�X����w*�	�1�8�Pk�{Fn����p����w{Dc��>R�M���[Y���f;��AGT�� �u�HY���o?\Ć���ϥn�6f�4���;۱*�LJƩg�Ճ�b�_��G%�\�3ʸ�Ơ��71�g�ƾ��!��vM�u�vu3i��5�3w9���v��ۥ�/ �����k�,���E|�(�{�Tc��$�}�>�2U�z�&��2�ۄYw��7������h
zl��#����s�U���	��GOhG%�l�Ь"d����~I$r���
��=W�%4|�W9�9V�_���tt�+�����@�N�H�R��~[���vͯm3����n@g��J��E�C���������p����Nm솸vX�?�t����͘�)\����3L�h�:�_󽊍�y��j����CQ�JaĎ��}Gx[t�m��q��C�œ�k/���^�����OeqUHaė�N'����1�I��jÁq�_��mx�֖ٔ+��5�_���?�i���&��V��9�.���>7�e�׹W+���o��W��#���E�-W�+وG:8{���.�@�o�Q��0t&H�~�#�AU!R}Q�tƂ*_�ϱ�2=f�S�d�_��2��%� ��)��if��<a�T��8~D\O�D�Ò�Vd%�e���r������-%ȉ��R�!P.�%Fk���I����Myi%jy��J ���x0��ȕ1��P�'�/ፐ��7���� �pz�����ѧP�˕t*<G_Zѕ�~`N#�%ϋ^�"�5�Ɨ��S���Ua���D\|�*��əX�G���.c�M�k�sS_/z2��G�-Y9E�E�l>[J�����ϛ�V��f7�'f|�"^�3U��|�ސun��a�c&�΋z�J"��-�s3����H���Kz>@��"����*�,��,�"�o���p��h�i�dO\�s�f$,/���a�|���9��M ��"H��q~���DS�\�J�n2ޑh�$��'!�x�p��d�*d�Zd�̸u�g6!)K��~�W�ġgf?�Ns~�������ޞ߫~
�c����{+s�`R�;�,�����y?�%�3o�����B(��_Yg�SK�e���'�����wMl˖¼�q���A#�N8s4��;�8vO|E�G�2!�;�d��_Y��ɮ��>��[N��&3��Ȓ'y�z��ƒb����0���WI���yJ���?���I�dCǴN05=��1�j^�7�)�͇-�ح8_����8�ܒ���w�W���L�l��p�`�&<�E�O�ª ��
�$+NTOh���w�B��n��?�0�`2#i���p7�����C�)�TA!VA�l��m������6Ĝ�)��ֆH�	�s�������UzwY�Gg��mP1��D��0���HM��x\��l���=�f׎��~�{��M�1�(<MfF�+��c��* ��1A�cV?�|���82<{0��3��҇���UG���92%�	@a��Z;J����l��� ��j��yw���D����ki��SmP!A���mZ)�ĭ#4Q㴙m�,��V'��� y�Î�q��>w!�E����ۉ@�ք���gW�*���ʘ��	�O62��E�`P���va��y�x4���d���<.s�LJ���fᆅ�(y�#:x)}�cyp�����xJ�̤֑ 6=;�����wI)F��CP��0$3<��Ben��z	AGK5d��D����.c1��sj	�䣴�ā�h�DEl�n�a^`�#DG���h4pD���(�#(��Vz�{��fjU)�����UO��O&�7���d�YT�yì���U@�*��ĸcj�U!E�J�QEci�����U\ W�����gD�ce'�5��W)}k�)��nǘ_3�H$��꒩�AĖl��w$��\��@	����A�gx�<�������%|C�B��I3���u��N�2��B�m�!�;z��*������]I'�f8���&�b�X�X�+`:Ј�"O�}�ok�a�ݵׄ��������w�Ѡj��rƆ.o�M�#oC5?�+�x6$��(V�U9���b��p�>���FX)��Q�b)�$;�X�Ʉ83�j�I-�p��G]t����E�F�cF�C�ߔb�Q�O�L �(��.��P�ݵf}�Ί��űj��Jk/\����nHhLL�SnE���x���|���F�;������v��D����e%��Q��J��.�lܪ��+���J�{�FL�x| j�I4���8D@c~�B�g��qH��,Ky�E^a�l��|�D�� ���.{�m,.fB�nh9��"iH�����y	ޅ'	Q�t��-ֿaA�[�m��Z	Zܠ,Y�C\�%��|9����.���Q���#'�f��n���g��T�L*������Q8���`��=jN������p��'n�B��\�ۖ�8
�3Nu������T(C-�B�섞rq�?!ѐJg>���4
( ]>��J ��7��fr�f�k&�mǡ���[�'���H6Ssk�8�1����Nhx�1WJ�B@#��f�� [��o�j����^l��r������D�u�Xql]Ɂq���~#9�$�rU
�iԴ�����]�7�"@��lRZA�
�N��Sr�|�����+2i�9��<�7Y>h�C?ڑ���4�%�t`�E�9G���N��.sJ�u]���'��S�!�1����U���Pe(���q��������&��'�?*.�}����م��C�+�gFRѳ���Ѡ@��[v2��P|��
<�/�: 3؋G��Y��&�I�RlD�`�5�<Ah��������6Z-��@��f�*Pא&ҙ�������80)� �m"�nh�H��b5"Cj���0�n��x9����g�r��Z/�x`�����������H1q���h��4wR��S�,|`�
�r.���V�O���0�P�ǈ9�V*1��گM�uQ,_w�hǓ=���Q4���|F�����P
D���p���M�+��`~����t�`Z�^nn������0���r�]i�J-`ܰ~���>Q�d<P���U;Hp׹�l9� ���^��/V��Z�|
٘x����t���c�Z�6���8ǅ�K7}�ceEe*�6�~�ܾ�ܼ1t�����_���&Ѵ�cPDO�aV��<r~�W�ၭ��c�&�܄������ �$N]z��reM e�Zc��-�}�ѫ̃.+x�`訢���}�'qV�x?]n!y3���?�18���)�Da����)�|�T*�c�=��[��Bx�t]�S�a�&GT��m��̭x6���P��ؼЪ���xB����B��$�:8v �3/P�5
�e�����
�%y�y���c��Sf�J[+�3f�TD^!mjػ�;��o��,�Iw !&s�nd�;�a1�[F�ۦq,	��&R�Cç�;�-?-��s��^��=�Y2��˂�C�fh�;�x!Vx��9���F�����):��� -6�7��Wz[�q7�a�B������>�U�����|�[�4����
�u��;�m��d��P�il⨯S섾�Ԫƹ��a'?�٨=b�OО�A����ͧ��MSJg�/�l�T���ȡ��b���F{��+�O���;�q@�j�&��Z�8��ʯ�+ɲh�~��{O@.G���|�홌-e�'�c.��O�ҳ�%��:����,gDT��谩�h�o�q���o�ݫ(YörW�>
)�0r���D@��Ȕ�Gz��yǓ�-Ѵ
C#��W;��yo��n9'Ayp�.{��'BGg�QI�xѤ��㧋��50���Qr�:��@��OWֳV���uk�<�|��PJl<I�����q\ÚG��WU�]���1��ml����Ҳ �"�wRh>ڢ;@�MA���p R��۬x_7L�<�`�'��	M,��ц��R#	�(��1�6=�)�dO�e̟��N��҃\r��L�Ѳ#~�w�۔ (s�	����&�,���	1���y�t�9T��Z2�ae<�v'����ګltO0�OVk[qBt�)�ʏT7�Ca�vc|��/\0v��# �hl�]�kK��=��VM�>I�8��/�r\�g��Sŧ�Ff����ez���CL#o�`�״��}�񸤪��iW�|�΅b~�+#'옢Q���y�F���s��G�5��0��,l<Y���l�mPg�rl�%"�G /����Ű*��H��6�|�8�ט"5�`��UB������'8�;�4Պ�ǫ�.�ޯ&	��u	�Z�)OV��&Q������`��;���?XJ��1�ˢ�*	J��C�M��*�iÇ��8��A�(<K�;Ol�ZlS��T��vk��Ii�ֈ�<&�ۛi�W�ʽIa��o���`�xn/�^�X�ΔZ�*�$�����h9�&q^TV=�po����7�;#s���G�������0M�Ů����5+����j�,|�ʕ��w|YI�,����ۚp��]��������� {��-�G<)0�t5�0-J��u��u�?
�����ק5�S�A`A`c�f�D�T�h��6��>����(� K�ICw$vn�2��BK�����@��_<p�M({�n���+�*}w	jh����d�T2���fss�p�Qq������Β�y9�6�Q�3�|�����XKtL�6�?[9�6J�P��S.g�3'�H#S8�>ן��^�Ϸ�ڄL'��!����X�i�C�"����5.�_~*Tkw�E����6�v��x��`i��C\1
`6��\�{65n�'�,�-�	�������Y,�S�LTȩ�1p�MO�2� ��AS�R����m�U�g�W�8w�H-ɼ�y�Y�t��d$u덫�tA�g��l�����c֭6����0�uGd��`ˌ�A� 3�՝�`_hs��U�r*��{��©�~�	�@�)C���d.5�� :�"`�M����!>���M��+�q�ՇBj� j���ēU����&�� ���w�&KvA���!�.��q�%�p�!�!1����-#�&��^W*珟Zma!?��,0>.�!��%��|IϨ����V�J}�x����/8����^����v�C"�$�+��:X���K��F��/�f�/�z��Ђ��"��j�D�j��U	P�S�	�^}�\&f��`�z`����>l�ۣ�[�}Gm�$�c�X�<8�����ږ�3�7���_#���ʏF�M����*��$>/��"���&��4e���g�j����|p����Pc�$+��wNWvi���e>2A)3�Tܨ�b��a��nճ�a��#���J���:�8���/e�� 6_�Bd��N�n!�zn��2"�:�<��zh�H��4+"���6���a?��Pt�]�E=�R[{��u�Zт&�Y�KX1�RQ�T���Z�9��-�}�)�R�\�po�rJ<`���=��av�}���o.1*����1o�=ְY��hA[p��{0�ևT �l�^fz���Xm�5�7@:{3@A�b�M�y�O�V���m��Z��W���f�~����ʜr�`d��5�qE;�j���V��o�E�c?M���mM������������[!-��+,m�U.;D�lc^@zO�t�2�$e�O�6"nF�����G����b& ����.mh��{�2�����ҧ7����S�_�T�����^^*����"�`�\����c��d��z�#����+�X�lJ!����&�D,�����xȭ��CN��&�B���'�;Մ�E��\����r�����. ��sY���X�3Mq�����Wu���s���=��n�O���^ncx������h-{<�����ʾ8�����5�A��֭l%�]�q�"�W�^A!>۔'!jZ�wm[o,���6$�K.���g�k�B��sP)��&RD)�Kdu�jM�h�q�<�;>Sb�$`+
*di����R��Ʋ����g�#+����c7AG��a�ş�e��ڳ<��
3�Q�?;���,M��A{��Q)KX��V�۷�ô'�n+l���6�Sp�r E�uT�e�T���� s��AQ'a�o�k"�v�E<�@t���f,�L�h�ɽ��^���@�DSb�V�G�K��U	wGr�_s �h��x^�Z���Tgh����B�^R:��@�ywY�u
�B�q�>br�������:�CӤ�7om�,��oㆸ��� ��hX�*��*��S��ǳ\�l�@�_!�3���mb$�WؓB������X ��:�1=��YD��G��w֚wֳ��U	���>UJ7��HgT��>�
zɅ�lCܫ]�k����lx����+\�UQ�3-�˽^9����f�<��ԩ�ˈ�[>M
 j�r�^���~��2� ��J�P�Q�"����bx�&�myh�A��
E�����R$��;�t��~�́_6k��R�-���d���\�<Vj:<l�)t�xS����/׍n,�7��P[O�<��d;25�fv�ID� �j�)C}]��&�ָ��R`�G@sIn�x
�FY�d�'9 'Tu�6�Y��cH�4|T�s0��Q<�Q����LOV;ܱ�H2k���.��jS�)F`�>��N�3��Yς݂n� �b���,���N�!;r����҉fzé�Y�PY.3m;{��	�Ou��O-T���j[W"�^ �"CR��x��H��H��SЗ��@jwvL��Djο��������˝-?�w��1VC�h�P�k���5���&[�R�m����xOPG�*�v���|��pR���T;i�_6�!�tn4�sjϫ�C�M���Y t�٤ͷ�!�/�?��X����Zet���� o:����EX�ص&+)�1�g�:Aƞ�>N��;.��]���k�� P�PFg�E�Ν�Y���{�p��x��v"���i.�޳_��=�,�����	��Y���3��fV����|AX�0�W�ƶ�4#���N�"��0�0TV��� K2��=C�0�bj�+6�H�FԘ��а�{���BPQK�V�Ӳ$�ʹ������4��S}���'.TĹ�'o�����ݩ���	�qy�4�p�2Q�Z�Uѷ�(7�P���ճ�{�l�Qg��Q����G��3�8��$��ʣ��$��[����Z�-iN���~����mm�)X�����eG�����7|