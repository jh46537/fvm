��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw�a�[W;���(���=�+V0�[&���`�F�}S���5気�uM�W1�����j�@�b��Z�"<��/uMZ�ɒ[�AuQ%TJw���b}��O���R���6~$�����!��S��-�M��A�K)�~�'���s�^z4�!ݖb�+X�YKù,��)ۀ�Um쯠m��X�����.�{�Wy�/d�7��#�l������{	���&�����	%�HϷ��bW���0��Ϭ��� ���s-��Yh��ہ!��8���B|(gՈ��ʅ�>�������*.���F"z��F8�ot�p�5P����?�Mw}Wm��4v�� �<[o�虷��u���sWؼ�G�Ƶ�YEw�솶b-a};�7�՝����:U7��A�(��2K���hD$���N9�G�E@�;N��,T�X�T_�:"I:��g�Aܵ6��)���H�Lzcz*��ZVn �^w�����V&c�i�1�g~�k��>X����&�]D����O���g.�҆ī�"����z�;��`�X��
�������
��1��C.��r��`�7��J��2�6Us?Ň���Kj?�F�C�_�_U�D`��\0x�������w�%>��V!S�,d��ӊ`���|�V��2E|OW�+��G]���@���_s�뮫rf(Ti/�[ZK�]zY��]S�	\k����U�f;1<O@�2x1+����cfz�%�.�(��������q�w�L��W��:3|C�/�������%� �����|�3���Ԍ�����d�!�
4�ڼ�����.���1�8�,�99l��t����0"�=0}�V8���^�ξ�=��qe �y��՝Yucp���Ē���J� �^�0�l�lTrU+�/��"��)Ư�!0���|�YZ�֓�X�#��1q�.�}�o}��ԅ5Z�:��"�4z�抍�U���[��5��~P}�f�`3~Ytڷ��s~${S�ܠ~�}͸�B�t�po���h�b��Q�5aI&W	)j���77ە �qh�´���Rf�N��{��V}�OR��Q�#}��5.|�[ʮ3�5�o2�WG�+C]�ˁ,~F鬦'����ܲ�dR��,U'Na���P�$� I���C��ƌ�&p�~�c�[.���F��!v���}+�JZu6s5F=�W��0�Kβ���^�(�c-s��S�i!�w�,�����;�s�4en��eE4aa�#������mC�?hF�i�j=�c�.d6��2��)qҍu��	5
�d�As�JˁG�C��o���6o�-�)q����o��%SY����JCf�V}�	ߋ][�2�qa��ү�ps7�S�c��G��gة���������k���cʴ��!E~«���'ެ���dy#�u��\�{��I'�gg�ű�n��[���4a�AU��a_��b�Ƒ�p����,6U���wx2W3�����k+��os��+=���Ϯ�p�os](}�o��=�r�Q�Sez��
�2��+�Q�1 J��,#bTKIᰉ*�R��2L�	��)��7��Ї�b:Q��w0�mEYC�J��z_�B��@9UG�벓�'��%덌Y_�{���F����V&�~����yf/��OW�O#�G�L��9�#�1�}_B�r�߉>9��-���L���d���6`O�����ہ�M0���H#�q��?�Q.��!�҉��9���.�T�1r� T���eޟ _��\k��'���L�0	m��O>Zs�2Q�뤛ToGjG;�p#����������~2��&+E����r':X��q�W;((�
Y��1��\/Md�o�UIOX��'J�ܱ��ܗ��4���P�#8������};i��p3��� ��W����t��%A쩢���0��D�I��D.!��Q�#�k��:8����*<�aD��=2�	�#�Шb�ir��b�(������V��@e7Աɧf�گ��!�����tg�L�ss_p2a�%!���fc��^X������Ig�'Hx(�@��PY�J?lhO�U�Y�)�c\�-[}d��!��y���VMg"��W�Â%9��Z�F�xa���2������j��L6��}����l8�����1��˪g/��\>�X�~;�f�[�#܄��J�����F���w�~^�����Y,o�ɽ7�ꋊ2��c�ls��׷�]g6��4��V�������|�ǖmB��"uN�ȸ��E����q��L���F��(�-Vi�l�N�\)~��k�-є�{�QF��u��x���ǐ�L�ץ�N1)�} �	~��T/	��X�����ߩ�'�u�F!��"s4�-8�8�ME��-�0�P�]�q�k8�F��~]k�5p�F�#ڕy�l�dX)фѝ�c䚓�>�:��j���y��~ U.�8q��WUFO�t���3%�6�c-)Y�p�~��w�c ���[S=hH��hmq���4�smnp���=p�d&�p���sn��L�+�aW��|l#�8d���#h��� ���ctI�7�2�8L��q������>~BZa�6��T_�p��~�#}�yI�<�nfw�!��-I�	b��mJ���v����3Q{�b��AŠ�*˥�fWƅ-�9�Sb��n}�i�9��T�lX�b�'�L��6({��.H�������'K��'Y�k!f�l=���9�sy�]2�"�\���L�Z��(������,?�ϠQG�����3��W��A�.�V��-�&�=����e�O�~�i�T�ڭ�O�rj7U�g7�v"�c�*d�:������FX��~�m۬�)�xs�����;f1�@�!��$�X;�_Xl�||=UE�kQW�f&�yo|9���E�I�)�NsM9�BD8,���*P։��O��Z���S��e�8SO�;�Zl�|��Pzj�d��w��8����iH�9�T1��H�%|�<a����D,^d���U�`�?��>+��l�l�;
���= �Ny!:���e-s�*��-��E�u)���s���죰H�� B�D���I�6�QS�,W�"7!�>�[G��j�n4��j�P���.#��&2B�j��|��{t��%�����b����x�p{{���ܤW֨�^q��r�w��D#B`�Bt0�4��m��#ρ�]��z6�t9�/X"�/A��d[�-(+��o���E��g$�5b'�)�~ֻ�'o��3 ZJ6!��Q)�Z�#�-@��YyP��y*�7��_�F�Y82̓�>7A"�1����I��.R(,/��8CT�Q����k�[���w��c�gQ�� ��j�� ����G/T�0(8���?�ٷa(�rlb�S��g�h�&�����V(�y����3���CYj�r���I�Cӡ����h,���4%���M����'��G��X'UU�$҅�Qy2sK!0���?�A�|=��&[�`�X{�p�E�}������Q����u����K�u�m���،x�nU�H�b�%�����|�Hg���U�N��5CT���v'z�f�1!WkPze	*-A�%���n*�� �q��`Hy]!Y0��$��jҺB����MWo�%��-�r���s4O�����?y�-��P��;K��b:(7|暮�ɧ5)�=��gPH]���ØT�M�qۛE����"����&����!E,H���&j���������rt-�mmh���h8�e�h���0�
��DL஗k�i~,����u�CET��/��(��w{�ѓ?���74K��=���j���-��Z<{X�}a`����EI�� �m}�������bFEw����`�.O�U��q�_φ�[�:�p VAK�xe���<6��կ�%u�S]��I�k�@o��� � w����[���
'� y�M��]��=��:;�VR?��~p东��quX�2��G��QCaZ^���R�%���^���p�Ȉ 3CgA���o��]Q�^�i�X���~c���UKz��)�#��zB��rA��]RK2 �I��(��Y\
�<;=}f�j>0&�eI��b��a���e�Uh8kr�>��O�Zm�}�/IM��S4�v���On��	6vU���*mV��pn�!�d�y�h:�^�� <�f����Hz�ą�5�l������4]I�t��/�3G��͠UN�F�)�.�8W�y�� ��,�ޒc(o�\U���U��y�)ۚt�X�b$���,>��츐Y��Ñ>�q���bF�/���Y�y�>��)XNEt�Ĝ�rv��y�r28��H��H��E##;�B��$����X�"�3/nā� 6��E�ŀ�> ]ẻ���3�K����pzZ����?3�Ţ������@�������E��Dޓ鸎dI	!%�Rjx�����u</1O���gv
��奢��ޭ�X]��Ld�B1�-T��-