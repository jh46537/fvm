��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��W"���e�EN�gz#)�)��a"���Ⓞ,B�$t�{����c�,�-��� k�4�	��[%��B�?���4��\�@e-��� ���u����'᣸߬Hӣmy� q�`L�S�L��-|�,���Ξ�<j�����̨O��f��U�,ﭵ�h���voҭOu���[�)n�g*k�<l��p�l�O
����1�e"��MT����t���*��<�i�Awd�;����ECF�ZC8��&屹_|��vlj�k�G3�*�萜�(:L
�>3���v�L&��p4pt9y�%o:b��A�f�����
@hQ6yP$�Q�f���{��R�e�5!�d᭟��7+UZ,���!��I�= ȑ���C˥rό�I�iy���3�V~/�N�6!�74@-q�^6�& �shn�'J|�#"����,�[����	�ε�Q]�ł�[���	8�m�}0��Gi�=mc�W�N�#��%���"���z��0��2C�Q�L���f�.���,`	�߻�ke�P����zhD���P� ��v��Gͪ��t!e�ι�`�w�Gܐ�bPƓl� HU5Β|��A���׋vdgyeˏ@����s7=���3�#�~5�[ߗGI�H�c}���of���l ,���f�sDfI��x�}�sӕ��j��0a�FјZ|��ִj�L觘�Oއ�q��̈́�N�y��)e%i�s2�qNSȷH
pu�!C@��R�8�7�7@n�1����������#Z�9���8@V��nF?�>s;`�3�&�3�T���춦w��h�Sł�mØk� ��T�s�W��~�.�X��L/'l���h�+@�G�W{ŏ�a_I��đ=f�;��&[��֞@��(er��Źɮ��ʰ!~}�	�41�2��g_R���&ki~+g_��$qxQ�>� �7__Ɍ�B׋�+1��-�=�����L]�E�$�r臨�(��.����=�`"+���m�pi�{H�$��0z3�+$ܔh�\��@Ȍ'S޿2krѻ'+�`��M���>l/��������/H�v'�o�����8�~>%ⳍrp5~��̯�;HQ�Z�@����)c�7�j>���h�G%`%�7���щ�+��1̢�����P <�"mOCW+�UJ�ʓ�K��&��m�6����2	�����D��]���hr/Z�B���FBgy�p�%��z��S��S�]�.�A�V҆�2��1��ވ���1�����1 &�g�2�T�~��n$�������96Od.��\)�(-FX���2V�U��7�_m8)�%=�]�{G���N�p���@И���{�l���M�a#!&}���ޔ}S,=��oN��4��\2h>"������;�>Z��w�B�S�;:g@��E�5��2���⃏�����e��̞rTS�l�A}aB�� �mO�o�G�_�Se�{�Mu��|��4�Ά􏰘�����R�>�3apf��/�ݦw+���"ȣ+� ���?+8Iũl'<`L�Ql+�T�F��A��^=��J��������$���Ԏ|�U��xF���Se� �_�5J��㸚a�4�}&�zߔ�b��i'Cz< �_\����t�C6�'���щ�9̇L8F�{>�$[�j������Ȳ��:z��&��{�= �.4/��t%�̙�2*��*�߅./��nD*�U' ����p
�H��މD7�,�~�}�8���ũ� ��nV�to;'��� �����~4
ϐ�,&!E�������^s�U���}�N�aD�@���D��oR��0�N����-6����=~����n��?��(~>z�9�[����0ڃ;7�^�[�|�]}ҁR�,���J��� �r4�wL�l�]Wn�cM������n����]-����u�d�m��䏎��$[U����a,b�Ẁ7_Jw�%v�X�d�!wB�+8��#|�0�-!������̀V#/'A�����W+2��%pß��� �!�&*c��v�Nls����сz&i���޸ ���:[&��M��Gn���Ӛ1�&�*S��ڦ�M�|{�Ԣ��� v�p.=��̖����Z|���r�@N��7� G���<��/��%�B5�L���~��m��o�#%:��g7W,@�!d�t��)>��p�	Dz��b����s���Fl�މ����4�nO�笄�=����Q ?��BI��|3�άp�dc���g)�t���m- Ѐ�?�׀����y~�=��^K9�/����T�3�uj()�hU�3I���s�pS2�g�&c�B��*a�GJ�4^4�c�!�~��fa�k�R�O/���0�9*��q9�[X��R�7c7Mz��-�b	�u�H���g3��S��-�Q����d>��|Q=�;��ع���&9Hw���赐�Jz�����@b|E.H+��T���*T���1���AO_�Xdc�JEg�����h���Ϭ�)�(<��R�f{��Q���:`�l֊y�Pt�-���ɜ��u�$����$C�"p��2��3ŰXG[�e��!���?L�3�"���y�+D#�b��[�G��[-���g���ẓ�tdk՞߄��e�r�t��4�|Bbi;��hG��CsD?��k��#���_�Ӌm�C�i��Ch;����w2�,G)m�dnb��[�u��OQ߯�~��)sF<ث%�ۡn݀���uH�=��?��D�s�� �Z�m��Ew��FS���E���\���!߈v;g��$�%X�$�[��z�P%w��G���tζ׈S����xl/�h-Ϳ��u��#<$�a��Jܱ�{gq�� �h3��5��d�k¬[B%4�+^�{��3!'k�FC�
z�©�>�S�6�uY�8x�f�8杪��n&��I���(IS|���������b�������(���>��B��v��p��ä{|�NP��YIP��pU,i��j+�;ɷU�_g7�L��Dm��L���䳮�&8��5�S�H��aG�U%��Ⱥ�*���� Flas����(��^�U�Hl�9�1sʌߊ�!���Z���p �)��L���4�� �I �{�{��k�Jl��U��B�W���IT�"�\7�H{%nѩ��j���7Kq� ^[�Ȏq��Ghw͒`�JD�����j�d�k�l�G�,~�*�L��ːYk�(H��i�>��j�vR�J��z2�\q��Hٯ]��jj��0CsVmJ�o��0#kb�Ht�EnWDk�_Ir�22]9��e���b�u-/���|T泋���B~@���d����<�.�A� �;2�р&���Y�L����I�'�d�_R��Ve���(��צh!!��c��:u}\���
��3>R���-��� !�m}��]*
E?��2m���]�9��#�DZ�6[�jc�ޜ�A\���	�����+�����S�E��6��g>v�����?R;�>Ng](=����K�oH�2sw�[����,_���I���҄���hR�ӟ)<�&���?"���w��#4���
����8P�ȇ����9��IJl�d���QN/:A.C�S`%t=��Tf�h#�4��ZF��xE�TN#ߍI ��K��q/ʗ\�g~���G/�)��OE�V^�Y�v��Ӗ���Ef�i��>�L������*%��T����g%��i�/^Z�U�.n�hXAP�a��<:����2�o�-{s#����Ӯ�>nOx$�L%nwL,���+��r�*��S8(nw�� ���<� �Il��,Y&[�����`���{@{M�Q�V"!v\S���3�7��"Aމ�}���O���n]P'Yh+�vu����5N��!s1�5]�Fy{a��Щ/g���v �c΄��,tk��w��f��p��/���&&vKf� ����kzg��^C��2!�(�fq<��骏Ѱ-H���^�<���O%�$��RՃI,��U�'Y��i��-3 E�Q:�< IT)�n�v�u����LcG�u0�{O�A��Ĳ�5�`�X�˗����兛\�'ʹ��pkH`^ZK>�4Ҏ�_��K{����A��/9Ab���fQJ��cc�X��0_hX%��(�^�'x~�`9���Q��W���+]����aD�,y^d�~��{$���!��$[Y�����4;�3</��,��k>q1��ٮ`�É��,i�-A�}�B��a��y��7��}��(�4˛����~N�x�t�y^�'��Xc6��a����?��F���MddK УD�E�1�����7]S@�}��^�dz|σe�5��d#\�$����M�
����Pi������w���)�t���"?ݺ�d�#�b�=�*!�!���[�$��D���EEϛ#>��j�P�����m+���ț3���_
��{�X�.`h�{f�q��v�*�YZ�l#����̒��L����Q�^��A��s��łؼP������μ��<��:
��P��W%�:�r������u���'-�j��R�f�2g�����*|�A~��O
H�`Ul�7B�'����d�t/��a)�+�5۰�E���qgm]���R�/@iS<�����(߼s������@]}W`4�����*�F���r|k3\K�(։ٿ�����U��<a��j�(J��}�C*��=«����od��<}3�X�λ�s�E�>;��5�<�)����Ī��.��(�/ڑ�=�v��"�P�_�ʌ]׈�G]�~��Ϟ%���Gb�͸�Ȯ���l�u}><��D��6���/�G���n'[Lc
4 ��L�����@����L/rF�X4)漲��%��.rv��8���?́<0��#��XZ<��x'��C���Cf ؞���q��:�`\A�)���L��GNa��^�=�W#,����$�xֿ		�bM��@�;t1p��^=�=�(ժ�����=��9�����@�X��Q(�O$<��V6eW��$�7Q���}C+X���^���B�Ь�uA"ꍜow�
��]���U��� �%�;�
�R���D7	n���"�V>Ξn{G\���hEv\����I�]�1]J���}��m��%3�pc�v�ȡO��i��>���ݷ�D'��@�w�U�.��'�3�4�n-��[3��J-~d�iR�2����ݺi;�b�&���q��D���D�7s����8��P.��=z�����׿@�WՁ�(4e�2f֫i��1!�2[�����o�����f"C�SM�5Nv[�L{�)�HI�އN��k��N#)���%M��%�~A7!?�R��^/�jx���D��l!�w�m0
�L�uå+;L��S�� MWR��|;S@�j�}�� 7 ��q�LY������odg�
�}xN��2qy�|6�vȌhh!�ջ�j�y�3��s��5��lW>r�)`E�J�Bc"�vh���,Y�/Aq��
Mܓ�_7 '�������쇤8$)r7�y��2��up{C�=�K�3P���s骲�c�92��q�
�O�1"J|q�^jg]���@~u9#�Z�U�q/ܫ�VYzB۳1-�������`"M���=�]�6�b'�0�m�KK����u���ά�RɰM�KG��[`�Ҕ,�#��{r5�6�;% ���n)�w�Ċ�V���?�_���N�⒦$2G�#�y�rh�y�J���������A�+�f=t�u��G
��Q�����9���W�jk7%���ĸ�@�yV�c����w�Џ�V�l�KyB�!��@���d��5�q��F�Vt\D���44?���	*�t}�:��w+�����Pz`����2�mR�c�3"!��<\'��'ggPF���)���Z�=��L]h��4D�8�DNeO�p�ٟ&j-��?�?
�6md������$<�/m���˃n��y�!����,uo
vW�?��(޿�������Bf}����jMID~�+�8�����ÑS�{@�3��6��f-������lVE_�z*�g�4/~�Y�Tpn�鑺��]pO����m�[�.^V�����Ak���_����������ڰ����۵�G��f��;�9-��Mgo� �3��-� 	�<T.��Ir�A��h���</,�)XТ� U8�:�5�c��G,B�J;��B��(�Vho���l+aJ�}��{��c��v�Y��c�A�>�h"�)�5�	��! {�h?���wSn�g��5$�A}>�T�ǌ/����6�;��0 �[�M��;�$�������xH��E�y.f��SG��u��e����3��_����?��{�F.�VF��W��Rk��9 ;G={p���7�O01��m��P,�F�7Њ���5[02�a�C' V݁(�q&�"l��Ay��B9��ߎ�~�/so������^��1�/�.!}>��hn��kQ	��]�����6�s�6�X" ��1/��+v�����>��%��{��ΐĜ�KzY������sԊQ�0z������9a�=�[���]ic�PcZ6�����A%�<��P~W-����T�^��_,�{�EnĽ֖H{�V��Ol)-fXA���80��͘�e�\/a�%�ԍ޵M�9��iW����@�h"��Fx�伾�@�8�yFo�a�c������.���%�Z�2��`]-T�Q��3����r �{����&;���G����'�h��K�VM�*��Q��˒M���/�g#F�=��j�K�Y:�(z7Ų`���涣>T;z=��!"�����֜�I�� Sy4Hl[]k�(�����rS�\���Xz�mY���pls�-)h�gŚ����(4B��ocw*��}�v�s�t�'DbW����-�{�.8��9p(� �-���o���Q��q���8��.�( PQ�ܳ0�/5���/���<I�� a����Y�����}�ն�"���e�%���!�5��Q�wʬ`���$�?����?h�W!�]��嬨�N^��)B��rr;���U�Onx��t%?����Τ�G9����E��^6�t�<��|����g�H���G��$��������]w�W�W��H���*�`�kAZ�׬&��'%c��="�C�S����N�r9;�S?�4�����f��3���Ӝ4�P��v�!��=;�Z_5Ε�YL������w  xbj7���2e�,�ȐěȖq��ʏY���H����_|"�q���4���;�7�}~v�\!���3ڃ͐-�ff�&�RZ�.�yd���>����ptEX5#��UM�tzi��&���<l��Q�E��D������B�������c�6`� ���?��қ-Gb��:�^���}�˻t.*�Ǔ�,� M��҃���WUr��L��a�x��U-�5ܤ&�֘�8t�`�3��Θ{L+�>'C���g"��Z��l�q*f�1��R�SW&j]]b׻��~0h�#94w�*(��d�@�`+���C)����/ش*�Ҽ;��F�;#)l�d/u�}��&I?1�p�i�K-�ԫ$�o���x�_�`E.���Gċ?ވ��GO�]wܜnZ��I��Y���5���B�";v�3��uO���F
�ɒ�B�Yr�f�ƈb��˦��l&)������d�e�ޡx���ɝ��"�<Q@,�p�ԇa���x�Ĝ$�f�AKau�o.4d�t��6b�6�x�88���F���� ށ�˞h�,PzX {#5����,��z\�����E����W��A��D���GW�A�����{���ᮄ�' 0:(AB�n'zS_$���
����F�qOz��?o5�s��5���d��l�Y|��K_����xs��S7�Y''h�*��13�F��W4t���s�w���g7�v��A��h.�7��ov������TFZE�,J���y�`�o�O�d�꯾ �ы����=�n��.��������������px>$�!��>�B��[aތ������s	>�0�(��΁A�t>Edr���ہ�7q��>�����+��&����.L:��&j�7E��CZ\ոIz�L��
�"?���w�����v�p���5���>��	��<ȡQBi�j;�HF[��c�7�4N�.��%6�ѶXK��{��q"Oq�5�V\D��ck[ ���_d�� i�9�䕢�&9��.;Zc����[lmKٛʄAV\s�����j	-�#pLY�J�d{�I)�R_��3��y]F�E���|W:=�؆4Y�G�[����H��`L�oY)�O@��D0�iv�P�_JeV��_������@b!� ��/&I����Fh�4G�?cS�4*mˉ��Ͻ���)w�<U�1��d\gW1�#kO�����#v�a��[�+�u��k(e@�M����axP�$�~ ���R�>������.�n'qE��g�����s��{̡�U��wҬ��³e�D���0���p��d�p�
r
׼;��X#�T��2Kn 5ig��Qo���^�C�=�L���N�m���jy3�����Nn��]��Pk�A�i���Y���k*HYɣ��ߕ�Ⱦ��Xo�:�O��U�o$*!�[y%b9M?E~��H��`=�u&�O��`��֍Hƛ,�q ]Ɛۼ�tжA�ڣ8wQ\�w�+��^:�)���Fx.]b�'E���RnCfe��2���������!��| m�&�Ǡ2�v������/7�|��50�
�p?�����|�(�BE$��!��%���1Fq��u���0�݀ �,�4\�Ә��7
.�B�wu7R�.M*���^���^��f��j��W���Z�������)|��'�UX�hh�0~X�d� B�V�R{p�޻,�����4�xP�@E�[!|�D��ˊ���[�����}!�PrQ�ޏ�h��ʦl����*�;�k�;������kU�6����P�^Q)�T�<ҍzօt�O!�Y2�]7x�t7/���O�[�E��W�ۙp����<R��H�{�!?Eeo�9��{�eVC��ƹ�s���|�5?�Z��(Ǿ?�̋��y�y)=��ݢ�*L1EqN]2V�"��=|��[K(`�;2�_:9J�*��Q�^�0�b�u�敷�&;����q��#�u�ܙH���'�@�V��J�����1�Y���{��/�y��S�#�0R�nwI6	�����`	rO&s���[���}k-��|�tm�DY�- ?�y}��j�y�VG(���RM��őx�[pa���������S����=�����i<.����S���U>IV���z�
�4wO��\����ئ��������!��R��p�F��0��}��a��y������b�(��M�0������轂�#�z���*��>�^�@J�D�o�u|< �2����$�������g �� Ú `S�k����8��b�*�7���d~7!13�N��ɟ+<���3t��,�ۓ���%�}1�$�0���9�80�6A�v�<����dU���yӈ�s3^pX�G��������EBn�ԡE���3�o6d��5��ʢVtP��ó���͸[�ͭ2��3��A�2薿̧�
�/�=�m�K�!���?���S��ˌ���50&x�A���<��QC���{g�����A����������ߊ��ыb�Ek�[\r�G��G7���f�|ʮ�6o	tw���Գ��8d�Y/�B�������X�������hQ����P��s0�lS���<��Æ#��~�����Z�ў���rza|H�݀@\��")HP����9$��<S8 3/J�O�In�Nxh�B�-D�4���>13��q^��8��>���j�KH ��[�∄���M����_L�H{"^�*��YQHl.�@�&5h͛nH���J��I��(�*!��Q�F���'��<6�YJ]$�f���Q���%^S�� ��a�����Ѻ''�U�ǋV���j�;MGg�l4ȉ�LY��ɲ6
��?���V->��e��&bz"��T5�3}z�#=�[9<l��5��)α�6���?IW;a���) �*���n[co�'�n���w-)��d���V�j�7��.T?i�.]����خ�lYy�l�E��m=U��ul��DT��Z���Tz��R���c'蜞��h��-��7Ѿ��C��6��ސ�g��]6���nS�y��Z��������K����<IC C.Og�D�̼[������y(�92�l<Z"��I&g���e� R��1QI���<}�@���{@e��M59�q�+��g�M��Si�g��=ƅz�
l�-���Ͳ�nV�T.�P�	�n�E�{�ʵ�y;;T�i	�4����)���}͌=Y�T�K �tw��sN�1�^����1��6�*�k���O���?�V\<����Q��㿼��Q���}�8�E�hO��G������ϖg�k��U!^ZN&������x����[��� �MΗ�GN�:��o,�L0�o
�] {\�x�8*����UAH�J��8�[����U��ծ]i�G}%�(1L������ʊV�NvK�P�U���|��c/�Ŷ3���^����7̰�0��#:��L��Ɛj�ഇƈANu�R����>�����(����J���"�d��$C��&M��7P�}�x��f�s�?ߨ�'���7̺i�MxZ2�ee+i��6@<
��rr ��w����,K��=��]���ɰ�W�y2fP����:"��&&�ƫ;^�	\�ӘXn��tg�!�d_���݋g�I�@��$R.~V!	�9�����z����Гj�",	���`��"�{��9�n��vc\���9������������ԏ)������o�3�����#>B��(Wu]�hY6�Y{�����j��,�ƽC�ѩ�i3�YI��`���,�^P��UJU�U�	�[�6W
"�3�r�쨖���+�\n]ccȫ�ޫ�{������*��דjҀc��|N��hsoϙ�<�*Z������ϗ��-�CN�Ղ7G���9'�uQ�ǃ�稓B����6���������-%�?����k5S#�k�{x.&�2'Nr����qB�4�����V%�V:�������G��?�IN��3����m-~<�I�[����۾�,�ѠMŦ?��=� ��щ�|���xǼ��Z�xEJL�Bop�YKz�nL{'#Πr ��ٽ{�!�~Ӆ����e�ͥ���U����Ƀƹ@��46�g4ja�`��継1uGU'�O-�7����)K"�,<���I����g�oE�|Ҽ�7/ov��N��J:�������O�@����]�k~q6����T%�q wV�L�P��vaE�V�����Q8���Ｄ�k�RN#�bcS)����� �D��	{*8����P�����-�T��:a�ed]x��Jg�]�J�� #�MKݮ]�j�X��)Y����;�s��������b�৪�[��>L�#��1���A[%�׀�^.=��!�XoLeS� 6��Q8Ψ�>	���E�3Fm�t���I�B� `�h��|p�q�Y
��h�eȑ�Ў���~������6h�B�E�f��?,�rV[�/p�P��+��[��ayd5�9��j8�w���q��i�eo�O6ҍ9xo�*��j�u�;V�����(#�z������7��b_�f�������&JC�ɊrG	 J��,�m^x��֯�$�5J\.�VUQ�W��q��3�c�X4=�S��x��6��~�u%�g��/���ل�b�_����)9į����a��D:k~)9�\^�ՏB"���S��c�p��C���| �_A�8o%���)�v���Gr!��؇�@�Z�>qz�S��U�n$z+F%�!ֽ��:n�c^�=k?f��6��XnS��@�r�i,�1k��Z�7�B�i�+�s_/��?1&53��0RM{�U8��[s���W&�)�3~i��>�e�j�~)��V�fݒ��d��������t.��j6UW�W�� M�1@�{�����=���a/̼�%��6/C|�
�^���DV9`oT9&/L�G�4�N
���Sڧg 3Έ\3{j̀����K���܂Ғ��hh�+O�U�?����Xkk�o�m!���?��6N��z����������?e��ۡ�uK�ļ��E�W��������n~�w��N��"]#�����d������B��aQOk�������1n��U���X4��d���ө��?F��^��0�s�AX�x�݊���w��p��"������xR�W��-�0�[Nd�
X��w4�i��ۿ)�/���ߐ�)�Y��)k������l�KD��_e{��#oUd/���%I�a��(�[P�]���d�F5M�z�ց�t^�����Z@�E
��8��j�3��G�����J;iq+X�4�O����gO�k���S;v��䔈6/o�w�����%�~�R��^h����H2���<1�+=4�>���!�}�B<�A��1涨8հJ�$�(�ML���� C�&�,7`zqNǬ-t��q^����J���^5���r�0Puj��@���߳.�وC#<X�+�����&DsH9z5)ԢBP��B	�������z7�.�-F�2#)I��V��M4�jrX�D�E!~GpD�n|`m�9L5����tr߿O���B���f�n��x��Ϯ��õG���O��J+� �XD��P�f0���U!�Kh�V6���NaP�A�Di�'g��;�0��P�羒%����1���LN?m^le��z��k�6[mM� ��>���N^eYs��ߏK�*�٫�S�b�{iO�s���=`Dy4d�ed�0��w�b����ı���Vi�͟|O��_�߂w��X�<	��U���/y�EՊX��TZ�r�a����(�2�9��$���׽br���P��m�ԟ�뷆ira�R�.�/�^\�N�7��y#�n2;�`qC�֒9�P�OcC#Hb���Ŝ���Q����x��)~�&2n��}�^{�$����i���]���n9%[��um�6�|B�3��ܻ(�b܌��R�=��d���I��Ⱦ1�_�����KN���su��f����-&7�wʋ@��@��d��)Hg�(�{f�p`��
S�]��ܭ�i=�Zߑ���]anA��6+[��7�D۳��L��}��Q�,w�����n���0��8M���G�C/@��yh?	^�},������u0�����,��VQ��M����V�@�O�����g�\G��"�K]t��.���r+�E�3��tPU	i5^��&���`���q�8��Ŏ
�c����I0��߷ݛ�4`���������. 7TQ��4b��G6�.+_�@�,l}'X�O��mM`��r�����hv��Rd<�����b�(����y4I�IL���#2/Z�}U�)K��ϳ�0 �p4�Ow�iW�k�v������Dq��J����ir�]ZhՆ�w��")N@Z�Hw�����b2Ҝ+�-&h-�M��i��5bZ�Mmv"�5Owc����a~4MMu5.���8=��<��M��O"��E�L�.%�%y�I�SF^�l�D�rp�%��X�n=��o�U3���RM�?0��o7�A��]�����Z�M���*���H��:E�$�x��]�A5%L۰le����ϪxJf���(�/�A�5�x�H7&f�ʲ�"A�} ���ȋ>��-���2+kjU�h�U8�:e��.p<l�i��*qҤ0}�m��^�re? ?��]�
�4�%�epӳ�(s�(�}���i�x닜�!qG ��m��WB��=WD�z�� �c��(�ES�V�=1?( F�=�`m_� D`H�{{j����?ƪ�7�^�L�,l)`�0�8QT�Y���	7�R��\s�(����Zf�bv���M#	ྈ[�:���4 d�	���$��`��;4�טi��:V��BӖ�s �G��s>S�ܒ���[V�n���]�%G��g6�(���H��B�H�e�CE�'t|�V�o2k��T����7�ya+/1�S`�>Y���ء�VA�g��aD#h����P�:z&�&�Ƴ/�}�[)0D
�\����Us�w;�lq����z����6hѶ���g�s�,Ə�Vz�Aj�0�ҿ;zyt�$�W��;�D��1V����[�y�����F�g��e7��25���%S!�u�5�j��8�;�S˹gS6/y�_��x��c������Ë�34�a.���c���ĺUJ��=dՓ��b�!������
������4%�$�^�"1�]�����-NnRuFk�L����L��Mdπ�؅�){i���f�Jcʪ�jl� 3�1�zF�F&W�e�_���=ӫ;���u/{�����������3�	a�%X�3"D��JY���/�BH���F�mu6����1fQD�.�'`�	#x"��o���-Y��n�v2Zv��\�H�����u�W�
aЭ��4q�J�ԧ�+�N+�aܜZ�ŵQ��:G\���yė���h
�p�ʝ�1�%s)�����(�;���(zFC��H�=�e�ˣ���!�4rx|	���;%�@`�
���V�m{�9���f��\<Me��0��#����Tĭ]���PZN8x��U�C�`��G&��������8f�T�IP�rUP��{��R:� ;t-�X)&�w�j��mt���/CX�xv���W;V���[���կ�"������JL�6�%��Iu4��|�R������a�� � �»��h�	*���_|J9Lt&���g�NX�]T�p��dV��h�J��7đt��M�.<+Ͷ<���@j�"� 8XH	`� �*�PK�wq�)�@DN����_��`���ZӐBNR�<�Uu	�)�S�(��Q>m~�N��l���ڈ7��6Z�+���&+��tN��`�=b+�m��|ayć�$kB���o�VşF�C��j�?�V���5+}�լl���+���/���4#
��qZ�\�`皫�a���v�Nb�����*�>���Ģn�:kĄ~y��|�[�$=�[rm��c��nI��8 J!G<)M�P][E�~���Ob�c�tHt���k����"�\��Yu��jw��o٬ܦv ���{�7�]O��c)�Tv���7��W�g�#�TQ{�U{���&�'�4�9B3!Wr�2/a�*�(�=�AFg:�+Dw���� �|G*�����j���X�s-�<�S����S�.ЊNRD�R�H��xY�m-�����ɒ��z�2y�KE��( �'�
�ĕA���*�c��{�-筎�|*��x|&�7�K�#��͈���Uˑ6� 	j惓�V��I�V;V��4�bݿ�=�����$[c�p<�	�6�tesBيc��Es2����g�fc�W�Ƒ^�^)����l��������41���Wʻ�JIx�~�����Ev���i��L�nʵ��57�\�!��q�����-�Z�̹��v|�v�}�F��m���4�zJRb3p�f!�pE� �z�7㓈wBFq���#Sg<���P�.!���d�J� ����>�g���0r�j`�BZS���� �4�_A�}yB6z�\M���E +:`;$���QJ�/��릮��'����ՙ�����AЙG��Qي������^�M��9�Q��;_Nd���b��"$�i1Ë-)I�QV.W�l�  gE�=d+���ٕ±
U���2DM@�3ߧ*B��~kf�:)�\�H��m'����ǁ�4Y}M��]Yk����B���βȴLB�9�.�$��홸�P���SAO��g5$3�+����6q�e����������*:�Pa�&�=��=��M'��	x�o��Bi�r��|�<�ـoQ($�6�1�V/��]��"f'%1ŜUPpr%JG�T�;��Hr��(��S���i�K��^�f��	0Ñ��H������j����j���[��4$�������![^yzx%��}?����!d�<��Y-�~�lU4�!����&�m��a�~`��P�~F�K%�l���YZ'.�� ,7}�\����Dp��zdn���ب�*�t�V�_�ٮ�[�����%��>Z-�H�Z���jf����ܿ`}�U�2� ҏ ǹa�n�A�F=Hv9���H~h��BÜ��5�/�FJdN�V�([f=��)��hXf�$����h���\��)۪���t���wh�`�O+��j�z��1�na ���J�luC�ɕ'��[eG�ᔠ�}jc��Մ"�'�{�g��uLZ�\�&���d�hI��R��T�gCi�,�)�a��"�8�s���֓�e`G��	wcD�u
�z���cSȻȈ+z���&����
��gpT*S��S�&�⣅�\��T�AG��+����K�h��/��kz�"�~,�Q�=�Ng��I��g�o3xøj;l�� �
��*r ���Cp���U��?�&�7�4�L�&�=r*���@�B�<x��������D��K�h�@%&�
uto=A�W��P�xĉ�<����et������K���L���ly��Ƿ��
r��iI%�a]S��O�r�f��:!F&�Oi���e!F���7�1�;�XP?	ﰵp7q�����vE�Ǝ�]Эj�yDZ�Z�y�!J���������m�x��㝤�ɩ�;�8r`�DʫÈ���j�ޙD�X��f�����z��̗����m�����Q�x&.�5x��M=\ԃ������@^�Q� �ZY&�� �
�|zm_��L��v�0�\��;��J��PlɋQdړWGb�f;zQ��A
�o?˓��d{X�:t��y	�U#Jي��ӑ�)}Pb A�3��dL�myC��z��^UZ
��������Wǧ���Am�*�j@Xc�*�7AiU}�=�ǳ�E��P�����8:��ʪ��7�� Q�WI��J�I�����X��7�(W�Q������~�� �t<{}u��5�:.Mn�
5o"�+3��]���nC��?�Zh�Y!I�ۣ��X�"�\�Y�Q�?�\b�
;�[���Ĉ"�x�'21e��%�V֩�]
� � �b<�n�k�������c�����$u�C��1į�������ښ�W;n}�s�i�*�L��\s^|�����j�g�0���T�
�����{��,x��#�/ks5���3�31S�̾�����ė��b�����i��r�ݴ�12��w)
�-�׼��A_�օ�,bk���]�'~IrMjP�kb=h���,�l��޾���))�������@&�媊�Gl(cv�s�����S]8 9ɲ����(�p;kaa�u�l��K�r`H��p0��F�R�ʢ�+;WD"�+|X*��Ĕ(d�qjP�$��[o�cQ 	:-��lY~�B����S��7xL9-6���	�S����U��:�\��Є9`j֡w51��z�\'���_=v?�V@/�5��jYuz��3��@.�am.J��
3������Sa������������ƚ�@���3��M�ƌ�B�W��+��h�$�nJw����*�e�oO�"K�f�1�}�v�L�E�����Q-�y���}a���IS��
���P���R�!!�/yyX7H		|�����Z3��#���HUr^p�,�:�]mz܆��^%�mJȿ�8h- ������� WNJOJ_���Bx��?����a��&�>����o�!y5�1�X��~�Ec��M����ze�8��3�0y4D����h!�8�A�Qg�p\��7�Й�J��]Ŷ{�m6��+��{��?��%s=���.J��yzl d9���B�]�}��a�I�}q�:k���d[̀N���[���.�e;ܭF$ǵ��Q����sp�y��ʑA�T�6�h���=���7mМ�^m �]�������>g��CP-����-���;���̳$�����ZO�xK�g�\�s�[�E3s�#�P��#���F�,�W��l,å��r�����b��0/ȃ�Z�}����mH�I�)����>��*��Q��G���S��9h��˵�_#�%^��X�Wו��sK�M�-��{��jYR�+q(Q��jF����S�Z�H�����.�h�n	�++�^:<�����t�֭u	�W�  �a�O$h*���Th&Mɞ1�8��*I�(V��^�b�|L]O��}`m\���5�a��>�&�[d�y'ZY��:�X�K��7X��U�Ǿ�M�A�E��J���e��u0�LGOӥܔ����u�}-Y��� �� ��fɥ�%e4W1���2d4���0�Y��~�.U��_�':�x5Y*9_�K��-iu
�?}*E�ّU�kLh8℧⚻I|ɨ�Ы��G����/Yr�]-��1��kL3LJ�lx[G_��_>dd�l%~E�ه�ںsv(<�胝K�+fkl��ڀ/���l�Dlu�^2�Tg�6��_p��0(���R�}N�)�򉢪�u�_j��ð$l8{��~q��|s�b
�.�B�^`�[@�8���������JM�t��ka�9�aܬ�B7`M0��-ӈ�)�J�٠��d2��*�#���݇�^�]�ߖ�[U�L�