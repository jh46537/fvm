��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�
�
QT<W���
I2�0w1�	��4�ж$�
^QG5U�I�N��/�e�]�XK೽V!��&�{,����ANA�t?,��t@��ٶӜ
o��!9#�;�T�[�q�N�KsW�fUÐ��6vA+�Wq<�ݴ�K��n��<<\{5��ͮeY�;��zp��?	�p���G��c("'�T��<��+��Z( ��,#����h)��-K�� ��2�?Y��'�f��^3ٔ�R��N\�o0�(&����<B���ˎ�?(|������0F��2�r
�{�^�vRK �1X��j���>�EdS�{�	����x�����%���mV9�,��Mc!6��&�e��mF|for��`bq��A�vHG(.��#p�	u�Y���!��a�zVa�5�*��<a�c{�8�aj:PH�l���)r`����+z����U�\?V����/to�k�mZ���0��z t��+
�SN<�b�i*�B�CDa�S��!��}��2/�$o'�Z��s��^�4��_6�`<ARC����\�����{�H+lٗ�g�$jc�js�����[ʹ�v��� TT�8���8a�fj�L`�AO%��~��P�=�쫡��c� N4� o�:�G��Иz����X�����Z��!�s����6U�_j�����8�6nH%�a����:
oF�#���~��� �ȐkXAmx��7)̾�Wmש�zlELg���M�>/��6m�kъ�E����'-L& ��;�U�%��w����d\m��#���\0Kuoס���O4z$PfU���#�a$-P���hPaKq�w6xdu�.��l�~�U����Ǐ�=#~$	Ͱ�+Z��&�S�L���')ťc����7K�Nӭ�  zZ-�^��/�K��7�O���Te�;��Qy��v��ʡY�m���8c =�BuR�v�lk��/xz��:�Xt����Nm�/�'�[�l��Z���^�Ʃ�����3�.s������dt�2XN�qA���W��V�2�2��½vT�(��ZR��ߢ��-d��R��>���{��TIxx-{���jDMh�&��1�K��qg�b�|fs�`-��~}d��J��u��Y��SJ�0+�Pf��o/�o>^����,D1(�����=]��&t�5.�*b1@t�
�%�7�q�����G$�~��#���9l"X� Kw��:�B��yR�i�`�PE�*'c9>܏��>)��ŗGy�S7���aqgi4!�<0��q�}��JI���q����e�ى�[��[僚0����u��7#!�P�|��4bv��Y�8~�+ͨr?��j]��}j�f9�MN�	�f�2u�����N�e�u�&���>3��*�_�D��9�@Z!}�My��l"�)���?%�� �4����Q&X�m�@-=.��xl$�vW�Ԅa7��gE/[�%�S����W���148ba�z�Z�]�%���p	%�Wۮ���C���\-���.fZv�NKW�!c�	S��� ��d)%	:Gf�0���߿c.�[��s�~����Ħ�].e+7��	-� F��KH�5?�c���]M���و-9!p@v�Z�+�c�/��_�<M���4Qk�nJ}8id�u��.��r�G7��/��2����O�h�T~J��Fşb
�28/��+�2�@M��C���Y���_��q��v���|�֧��E��ƽ؏L,㷐�K�5��%��z�F���R`�d	U�N�K�Lx����lH�����~12O�3��I��a�V�?eB���a���D~P��~A>8Ɲ��^"�^��(}��6�X&���r�������{Z:���Y�N�k"ѸK�)��s�<�_
�_�vty��*��YjO`��z���<���KU��L���CK4L8ۼ�3��ǹ�?b@��13�~_YC(Y5z���(Ħ4�5���T���ܬ���C$p6fR�p��g, *�O�Y�O=U�HPp��QV����&)������g�����	1G��u��hi�>O	���
�_2��G�b?�g���j��n8�·�N{�v;?d*��\������S(8C�:J�ί&?Ż��<��Zử�̚/��*���d��[���� d��������̺_5�$�u&*���-b`)�n{<W��྆u&|]$�QcJ���*��B�����j"Z��2�6?}3(w���6���s���=��0;Wl5��M:�֣��|#�[e٣�
�-98L�� 8�8��yt�i.�G���:8ٟk��4E�}�0/"�T�^�<��J���A}�L´�� {� ۲����-\^*�oO|��&AR��:> ��i6Ͽi5c�?R �1?BY%8~ۗ�V�d|�:U�eZ'���t���~͌�����b�<�5�����{��׵�V�r_܌�X�Kb���yT�Iu�v�Y�[�&I�n��(�/��6Ctb֫�
�b�&`_{��ef���o�_��Q�Z5E�-�#��/-dr�㢙�����N)$ɒ�NB�Y�����ͮ�[C�]12�:��w�;Y�"��/X����b�	CF��y�9�6>��F�o�����9+-��p������(� �y�|<�{�3���A�LȰ�\��
�Fڊ�,¥+�Q[c��L�/�8�+k����y lB����*0~3#;9�QO2F��-u�]����U���]* ����
TJ��.�XR�l����[rZ�� J�� %eg�f���1|��z��nOC/��o'7PZ�0,��:$u涸/��x�9k�V���Y�e6�v����N��
~�Ӵ��N�\�Z�H壘�ϔ�צ˿#�,��K j�+e/T��+d77}sȢnvy����Z���.(�fck��FTe�8���%ZaN�O�n���\ޙ[۰ A�v�u� 9yA��W��Z$� [�A�4���~�5�������Q6���78%������h�˞�n!��
j���'<T!�:��Yq��E`�p��]�������/��[ds(�p?�hs���k���g�'��n����焵�C-=�}ڠ݃�7��{ҧS�yB��=�g��5���WhiV|�����׻�-]5�"V��О_,K~����;� �h����y"+�p��|��Y�������1��WU�S�ıՏȧ},Y0� ���a�*��y-����W!&zWnG��$�Z�6,�Z���ϒ$j�[�i��I~�Z�P�ڶĢ:f��"pd]�lǿ���hLJՙf��)r<�~�ğ�� �ν|Zf~�z���J@�I�2�E&ź��.ww.����̱�ԭv!����B 2_ua��� (Zb�]�ye�h4�,��8��HkU����Ml_1�#M���>�8��i�N��L��|]*�^��h^��Z��Rk��"�|�8/��J�Jdv�[/)���W$��8%%�����Q�+�ǈ��z���l[�d2z���}����� �(D�����-נ~�t���c����eSo����$�L��_�7��L�u����!^��Y��L�r!��R_jU���)��ZO���|q�k����(���%�~ :M�;��p�/�s  �0�M���hi[���)U�TW����}��X=J�
���,n=y�.O�ث-�I��2}��$�,��特����� a�H��z���p�xZH��UU�X̵����	dڨX)�
˳�x��b֊4�QU�:ᭂ��PjˑN^
n�E)5��[V�il�i�9�IĮ�zd��$�+>r��El��"��l,\�_5�]����g2Ǌ���z�$����,�Z@����+[�V[#� ��w������x�����BǗ!�'��T$_.cIQf�Rg��U���k�y�>�jX�B����A�^�,�{ښJ�|J��ԅ\6���ɕ���^m/�|�O>UY��6k������-5�]������\*^��-,�^6�?C8�̦�+ZpP���ļ*�1�J��2�/�p�~�[h�
SzQ&�Jw�&1�(�V��#lW������X��ǘ���pwϦ�S@�D�d_��dB�z<G���t��{ŰX���`�El�q����T�<{�Q�i1�i��^���؁������s�GF5�^,�(S�wWP"���B��9޻����t���#��7t�,�3Z�>N*����<j뗾��\�������w��)#*�̐0��U\1�[����r���&��[�q��稾�f�C���#-�L��wem��^u�����G�qJ~�_D��� rMh��d]�َ��|���Ö.�6z����н�>BB�B���3R@1�ZL��mdVD/���<��T8
���d�ŋ��\��jv;����t�~6�����V�~e-�'��wG/r�~���B��K�P(�\���S"�u8�U�S�nz~�I�qF!��O���������xĕ�E��=P�Bʷc�7 N�����g䕍�=C�d���N����DD��ZG{��~�^��3�b�P�ƁB.�?ܞ�&��
��5�����!��#���㡨m9�} p�Å�P�w�����@�g���NA��R3��ǀ������ -Np�8��rj<MM�+��n�,^�_��Ugj�"���/g�H_�ͬ+�և�g��+�q�m���]�|��2�^7�S���8�>JPVU��&#:Xa�F�c �� �f�C�\�k�`��E�&� W`7p2d��o�v�j�/�plj���,8*[��x>�2�#��v�v�E:��{�x���]�b��@>���߾�2�����SŽ:5޸j�h�D1��7ZCzEXs�� ^iBq��W����K�ݳ�!����<������B�0���[.�t�T�h+1���	�]���.�t�#���v�~��M}A
d1�$��e wjk5����O��nx_+��v�l�[���8a�����ʋ��%�1�9�<gu\�|U�r9*b�q��jާr�km�9�Z�6�{�xɁ�#�������t� �LD�S��Ki3UCdj��5��6<%R2���2��H\��aKx�n&@�ְG9v�Z�����0V=�y��yW�e���q�Z��$� �Y� 
^�U�2��Ez@���j�MT�:i����������AE�Q�g�Ugu�V�aE�0�\��-�T9�3f��nli*�}A�%!���ѧ��n��hK��G-��x�3�.��;Z�?w���X�>��/���n&�Ɉ%*�v�YUm�2q~f #�?����~�S��Z�6�����y��k~�b���ҋ��i�ǎ�SI��g��}�!��#�n�� �ʪXv�����bZٌ���y�.�v�>�Ǵ�˒����c��LjK��.?�K0n˅l���l��k�������Z*h�k�ѓ�����6��G%����S f}�8���!"�u�((EQ�4��~>z�G]4�pD�˄�)v�TM�~��(F+ϟM�����'�`��G)i�� 9��+T������	j=�z(2���t�P���/�@{�WF��e3�2��b"y{2�{�&�V3o9(urP͏��!����U#�2����K,�z���9Nµ�h����w�$g�ĥb�h��J�����|�y`���KC�ٹ�1F�ߊ��~
��g����P7K������P�*xi��J㔗x���z��L?4#wlyzI��e�������l�i�>�[�����0qC�+t�=�QG���G7�P"+���q��T�߇�ܕ�K�t֟���$�_!�>ӸQY] =��ܪ�y�D�(���<<�3���W���P��|	f��f�O�&�n����EhA1��M�	w\�X'f��6�R�DkG�i�NA�s27D�%+g��GMdu�g��j?�����d���H�������׏�'�M�c-]fM&����k|���=�bb��p�|�Ys������yd�b:�lS�D���W���
�;��>��i�99	0DFPʝ/=�)�j5|3(�5; �m�7" �X��љ��V{K[g�$�������|X<ń�a��Y2o��s71Ͽ�>��s1T�ؑ!\��Z����7f�ų�7ʪp/��2����U��{����R��m�������b�	X����lac�[�N��z����\o��b�g�O?��9;�[�,�(���Kޘ)�Kӥ՗�����>� |�1��3�����T�MC�jP��F�tO���
-��J���nh������i�@eZ{���E�x/���U��>�,�f�KJI�Zg�b���,g��Y�g1�%3�`%�ϕ�Bޝ�g���D&R��x��E���Ѽ�Дޓ�}��ʖ����<��#�^���4����K��@�6��Ǿu�jԇ�N�2�u�*��
n{\���������b|}�xʴ̃���ו|`n�9z?<�_J�7����b\�p��"WD�������s%�:)��G7"z��7 ʟ$����&�l����j �0&�y��o�9��F����@��Ѓ"U�c��$g�;����=@��:�ɮ��X��X R�̎N=�?wZ����}^�w)׈�s�U���>
U��m 6�����^=��1�֦�X�a���vv1�F$��O�� �ȥ�]��X�W�h7�ՠdyK��fc|m�mo%�d;�"�-ʲW������j��r�VS�&o�)���I4����v�j0o�{�T�[g��H�Z�W����qp�rQ�^.Ӻ�Eg4;�$�>�ȣf
��t>5-�ok�����r�4K�N�<+���|O�_Գd��o��B��$k�[�{���==��֔�	^U������0"/�{C��L�	��UcLk�z�����ד꼇� ap���/1ڌG�ys������Rg��(g�b]���2f�-��;���R��)���"�@etld�{�[	�Ktz�f��7�/�T?�����e��e�c��4���6�8u�R�h{$Q/�lY�zdO�X�!G�A&���3߀X�|C��f�bn�����´H�Z��v�ߎi��$��#��.i;�7$���ٰ���k1�M.�FKǖ_��lup�;���y4 ��8:�0�[���O+�����Ds��}��8:(�3hM��f?����_�y�B1�dxђ�k2눯6����Z�B2��Hf�+�/%:n���8�j9�~o�Qz9������I#?���Z8��%'/� ��� �߹c���<�X�Ċ.RrƤ�D�xS�=�rW����.���$�A�b����Qͧ��3�,h����[KiQ"[�^*�Z�k8��%vk�N&�)Wҭ��`�rJς�.������r���Ss"�&={��s�SE2xH,f�[Y8��B���3�|.�?��A�.H�Ņ�q�ס�49|����}.��xc��������gqNwb�f�eۉI��z-&w��`�l�RT��3��L7t���MZ�r��o�'�S��`���:�n��c�4LU�.nzH8���Zc��w�q�x�|����ܷ̒�v+X���V �a��q_~�DX�Q�ZF�M�(���]b�bH��Ds}�ڴI.80� l�u"��&{A0E���-c[���R4�p�G� 5����RͲ� ����e"m��d�]���y��1<:�&������E*'ޔ CS?n*�Q�D�Q&�j;��% !ʂ��	aJF��R����T�ȍ#`�⇒��Í�N�e�n���x��̓�fF�*˞LH�����vt�$џ�2Nt�dP��1��x���nL�����s����@4��T+fX�C�X�b�2=����̲?�2C�U���P�� �g7��������˧�a:#�Ձ����$#����ڐسek2�S���/Q�m�=� !�$,}�a �TE�Q�ew���v��#o��ەg��V�z��,��Ϲ�Qhn}5�����^"~Z`5���!�4�� ���������>6h�QR�b6�׬�`�� ��0ގ?Ԫn3�}�腐���$5�'�n��ջEV"zj��R��F
�h%_Oy��*I0�1�%\��V !�����J��l�^�wHV5�b6m�y�ƒ����s�G�M6n��mB�gĞ���	�����s^����u~�7��i�
���VT���~C>��;8�ąpY�P#�Ʒ��7�����'��@����R:��"�Tl�õol�9�j|�%��{�w�Z"޲?UrMՆ"�">u5�_#so�J��P��;�B��	z���/%�KT=Y��;TN�&+iL�OEeP�9=;!Ű��ث%$��_�U��������7���s�aal,b�t��3I�a^�ᗅ3�����:js3�h�Y{S���9C=���=���_��~Zm��a�����D��\��?!v!ϼ\�<����ɼƗm"��Sp�������L'����L���IH5Z�t��}����'���!p{$�p��?�����˗������/oF��m%ֺ��A� +~H_��>��Mo��+��,�c�(���Y�ה���QFO�_O����G�%�G��͸��#�#�H ���-*� ���|�?�IV�!�y��#�s��}}�*rI�g+&�w;�c��NU�UO� ��ſ(�ʸh�?nE�B��� ��g�=�9��[��IEyO���s\r�#�A�g�`�כ��&8Y$���<h����I=<K��N|�a������AP3��h�2�e����r`�qN�{�ʩ
�o_L�2^v6?�^�T)S�B����� �L�(q�K^j��\3Ux��� �/KJ�w���*
S?�GX���\�d�u%F��j����u���!0��:�����N�WR��;'�fҜ2�Q�ݜ 4�7{�<��:�T��y���K�Ew=^���q�k���� 兏)a���j��3ތptok�d���RjK��IO/G��3�ud����iNf���R=�4�^gE{ J�QA`jn����l5*��$UvW�\�
�?�ܵ��dw������!�4D��c����3�p�Ϡ�����a��1L����Ó./w�5ɗ�c��
���_�w�.$r���ע�M��o���d�H��$���'�-l7}��d[��&{�A �X���A��G��H��، ����2t~T�Mś��B��`����'`��F�"i(�a/Okc��ĉ�sn�uY����9�}��N��p����R���X���C0�m�� �!ɱ�$����t��0ן<�z�c��
g�}B����X#�a%2V��@EO△��(��H���<�U)U��ќ�h��-���؅l|��K���mv�� @	>��״�:�]`�@�J�=u�Uڄ揳>.��A"�f}�����k䑵n�H����X����U���� ���=��S�E ��4�5��3��>S�7��Ha�Lb����-��%�g*j��>�2~DR',JV��EdP�-#�d|[{���0ȩtI`Ic���e0/��ڸ(�a�߷�e�L+?�0�9��I��y��C����c����)�'�n�S"�����/��|&�/q͚�y��yMh����oM�0�-;Np'���h��jX�|���^-XܟC�����k>��1PkG����=o^6%D��6���}��{S�Z��9n��ܹ��C��<R�t�(��)(��?�Tɻ���x���y����so�*�L���or��4�Z�p.����3�w����h��H��(q:uot����ܢ�S	=�U4;��qYvD��?=�2��
>@�G����x`�>�#��S��{��ۍ��LESf?�S
�Ȇ����G��pd���U���}1(�����tCw�{�o¢|`��P+�>��wޫRф�7�D�(K���Mm�oR�����Yץ�<�$��bC�K�}|0Ll���_�#C���$ϤaJA{�v���� f��MX��I�� �^;Ց�T��>}u#g��,����0�/A����瀑�ޤ�܌EZ4��;�
L^5�����Q*2]�-I��~�D�b�sSa��PW�s KN�%YZ�Ng�M0�A�����o���o7b$�O�R|5�K�iX���w�*΅sr���2>��gz�Z�Me��݆�ȿK�F������� Y7:�b��w��P_�0!K�w�7�$`�g �B&����p��Y��|�׼��_�>;�[R�)*ד�ق� ��[p%�9t�Ff�Bv\�����pƠX�_OR�~G���k��e	w�/R(�J�%�T5*y�����
i}G�p����Z���Fշ�y;����{tT���yR:S�ǔ+=Vȕ����7�� ��{oT�]V�����!� '�s\���n�®2:|�3�@�0*\�m\�	#q�0���i��"}(B��p91����Ţbd�T-�x�=��.�y��R[{Q��]��~ٌ��y&Gk���Q�ŧ�	����@�oׄ�ru���2�.Y�QN�`�G��6X͉�EC�A�_�8q��ݲ��,��g)n\��#�l2�??���ۻ=�~ͥ�{	4�E�J��j���r7E���Y�t��~cs}�'N���'����j}
�e�8`�^"�x���"R��}DdW��#��<*�.'��jw�W,$�S�h���d��G��5�lkL;>x�/V�l�<Mx�Z6�|ܳ���y��G$	~�0�	���ә_���'�N�%е��
��U�򝽾�na����׍�Q����\W��P����o�D�A!Ƀ7��6��i�I�[!��!�G̚�����e*��Sn�k�2Ѓ�I@������w�����*voo�a�ֺ�~����X�i2����U�@�Ӆa�R-M
�+OJ����-� �L_*E\j�G�{�ܒ����2(�	#u���_��>α�֛�g�����g%���'[�A�(�c	��dR+�����]�T����|���5��?P����_��Ƅ��u>��
�:	-�.`��z����Fʦ��˛\5$}��I{Ai����3h�R�s w\���lB(�����ڨ��rǒ��A����"��rA��!�0< �D��y�Yl�b��w�,n�qλZ�M�CY��l�+;i<�[8�P��-�P(n��/�Ed���8^�7��"��(�e=Ş�嚠�+� ��k����:Ea�}d��EL�6�[�ZJ'EMH�+{��;��j�<W����E��{#hVպ6#h����y8�Se����l�B�i!i.���wl�9h��_a��n��Ho_L{o���=����谸�l��T@�V���t�UmUڿn�Q�j�����oJ=c6rO� ���¨s����$�����ϡu)?$C�6pDT�n�]�`�U�F�AɅ|@]��:��Y�}�5\����XU�X��.��{�M���"����/����0�}�V9�6�B-�6&S5��
�A8K���>o��1D�������I�3HN��@t")��'Xݽu�g�/�s:�b5��ϑ�<�3������_�����#k�#~�zw΋s	�ҽ��.j��z64(�~�n"0RL�&12���pKL&�Zv��U��.5�U1�\��"�y�DsQ~��X�=A�W����1f�[;(��lr�xV���_����pK���z�o��t\X]z�W�2]6I[���G͉��Q���nd�0&�K�}��8�˒�V�.�N=�qU�@}�W�Ul��I`��OI��.�����s������*�!����1v��ϲd�6�dE���'jV��Fwk����ޑ�*��*��.)�ae!L���c��&_�{ю�~{=��_2�_J��+��P�Ћ7+¿��}�O�_�8^Z�hQ@]���#'G�Ga�n[j��0��_҉DD_��c$����п��p��G��rXo���^U�p���9�0���Ew�sj�U�.TXc�rpI{�2��]Oٞ���<Q�j.���:*�6Ȕ��5��$(Ćcmɋ�J���:���Ng�v��-4�HD�U�r�4��ي6j_w �~�Mr��e�ٮ߬��3����e�{G<8�$���4D��:`!����w�b�W�&�wa�_m�Q |d�[@m3���&L-I�M��J:oo��6c�lGԙ���xq�����K+~���>��c�E>��M�{:�Z�7���@�UM?J�BQm�-"�p)��ˌ��[eBl�z݂��Cr�k�,��ݣ>�9��;���Оx-�����r�4>���#'��dX<hey=^"E�7��<5}�:�k�"�i�t0C���@D#K��&�n�QB���E��p���
ߕ,�Q�6Zm��	�"��{�q��gF dr����4�W�l��if|B�?fĆ�����0�Vh�����]jA�d�W���B��ݳ��.>�$��gc�tSÀ�b�[xicb�E�f	uF�ɹ\��E
���(�-�YY�^�f'X���\���[�"��ɲ���N������a@0tc�Ag�K8ˍP���ݨ�-K�l^af���X��J&��D��UL;��-�=���j�KG����C�c�F��VԓhL����i�:�?��
%y�����,Rg
�]?�v��q4��@���y�.W%�Y�(��ik�:��?�]Y|;�<�@� a�Ao�T�Í���^� �S:һ�٢���)Ԅ����'1~��8Ċª_��k��Z�Ul�ב���*V��Z�vA+x$_K��N��?_��j����ߝ}�2�e��$wl޽�}�#������ǟ3��Nl{d�� 4�գ�G ��^��rw�ۡY�~����:W��bQmxO��N=��w�3���8� �'�u�ᰮ6��8
ܑ����OJ��o���s��`Ļ��+4�N����$Z�C��P�ϵyB��٬5u�C�G�Ľ����J8�\����4�-� -�m�l%G�|��Q;�_�������|��ܹx���{A秦���[,M�2LO����OU�B�4"�cdX]t��P�*g�H���i��K�-��7p�V$NbT��Q">�JnG^�N����lq�u�	�=���k���9��rJΔ�6;��cSnL�l4���{�u��MX`O�U�lWǼ���{F�2)�/b'�i<���r|���;/(�:�A��ι��+���/��Ye�����K�f��tN�G�8��8ĳ��(nC��K�8����_l�b`�����Yb����)8`�Ѯ�Cş�c,} `����	cb��J����6,<�B�F���k���b����ĳ���ď���_Ćk��2ye���L9�uڌ��B9�XD������؟��sm��X�'��U2m��N�e�Lg@3	��:s�GqT�����9G:B�q��uw�.�L�Gd�����X��#���a�?a^��z�����CN�yK[�R�D(J^�ӧ��k�,�C�d~"d�o��l䨅b�;�����j}�4z]���.�&w��Q�
�����D�,�r����2W���ʉ1�9.��`��a��<���0Nۦ�@��;�\[�Q�U<ҁ/_��YS;���֢m��`+F���Ζ�0�g����V�F�Gʦ1M��CK��h��FK��I;"�m؇�����s������4�#�)���b�� �2iB	��*y.!#�G G�B��7�X���)
c����������H��CE��_1��	��N-X�%R�?�Bu�:9��c�Rx��OI eE�Z��U��7d���z�O�I�j�g�``RȎ�;�� ]�������oC#o�}�'�e�UA�}�/�*1��n�ߔ���}e�(����5��O>{A�¨�6�$���rބM�{S��#Q�I>k=�wE=)����C�	�(�.�`�d�ρ*�[���
�֦ck��V��8/޷�0�5$[������7�.U"N�|$牵k����W�d`�۠[6�DO���o�V�����\8�u�������u�vB4!��g}�B��ą���pdk��żI��������*P�`�a�T+w($ܑ�*V{����E�ei%T��r#5����	=��nO�m[M�h��C>����	�*�4����E>�g�얢���M��j�	���.���A`q+�yU����j�U�������H/��}� ��.�Q�5<�86H3c�����^�T��#���D���~���W���8�d�,/����Y�͚�I�|�'��60T��-�Q)�&_�ډ|f��Z��s{ ��p|�鳌�M�#&�ł��l;����W�-b�H�2M+�*q�7��UW��ԑ��5W+C'���+wfŁ�o-}6&�v�2�X�"T��ب���k$^-���|��4���P2�s�1?7n�*��[����>�2��Rc0KU��
�(M��#�` J��rͅQ��\x!�����p�.��.�� C�<�4q��L�pY��t튛r��񓾣�߆4�)/�XL`�E�	�ѻZ�F{�B�U����W�I#�~�GΎ���F� [������Y�D@�0�;WG�~�(=�i_��rQ������{�)��=�_v�8�Ô�MA�	�@�BX�T�*=Y�Ӕ�p!��J�� 3py�'��ǻ3��題�u=N�����Sl���|*"���o{`�`]��;{o������7^�F�M	Kcq��R���8��8; ������kf7�ńk՟	ҋZ�������m�C�g2�밶p�_��#�q��vL�]4r[u���
��!]ȹN��d|U�uj�mUk��+��i���YXpW��l�&rVX�~�R����e�)�׷��d6p�ݴɋq.or��m����B�7��o��g�+OO�r7���v8�G��7ܽ����o�7'TqF��� `B����r�=A�Xٮ��ǖ��s��"oz������YFD�-2��%����$�MM�!�#1��g�/���M���A�]F�#d�7��H���˭v#3�i,�H�n<y�z-�¶�c�ʛ���*�b*W���i��,DC|�}��5���iJ����<�A��G�E\��=���[������9����=���$u�G�h��a�� !��ʗptL2N�F�6P�x �۵hFv�b�k���kL�g�Ahy\�W��-��0����Y:�.P��y/e\�%��=���rO�H�^����E!�M�{)cjdH�j2R����6g��z�d	�������$���i���kV��֘l�!�J/K�O��5��� j`J��0��EV\��e�_J�]<.���D���ʯ�����}��	D���x��#�!'��*g?���2"�Ҹ:�x;D�hx���
��^4/|�k��<��f��Z��4}�����+������HFQ�cR��7���ՔhsD�F���(p���5
?9�씤��q���k�8�Wƃ<EƣR�=�;,���^�,|���.2^*�Ӵ��<8E��q�[��JO�"Y+􅾼QȰ��i 1���'�07B��B�L�>3��/�0'ӎC���r� G��h�O�.O������ki!ATo�"�4�i�K��y��:=c�j����N(����V��8�IC������N1,�E�6/�>�u���K�%0��#t��"s���t���]HJ�~�Z�3�)��V�� ���R�93Z�c����M��]�8��������J�j�e���y|���G�}����-)�V6� ����'�۠���H�_��w������QU���x�5.�&�������������g���=؜;Ϗ���5�]߮����N���e�}����	s�h�Xf*�U�����gۉE	���HV�;#���`�d��L��+A#�Â����^G�%�,A녒5�m�O7�� ���D0���t�{����(Ny���J���޶�L�E*���%�Hg-�%+r^m�n)�g�̟�-G%�6p"���`l�k�!D�T��o�`>K:�WԨ��#���A.����������8S2��ٺd]�dn�=�G���R���=DN|���&P���Q2zF|�4���2d�F���ue��:&��M;4l��=^`�r�9;�+]���R�^�d|T���d~$��ĥT"�6��]P��P�WAN�Oѹ�����H�z؝ÁKD0�عhg���p�%`�e}q��n�i��]�gJ����MGckt�q�@�vZO㇦���X0/
�9�6酨25�'_���@�?�k�D:Xs����c��\{�S�p�����="�59y	���H&�@w��6�k��jW[cׅU������\&�1W�Ր���A�$�ϑ�0�ƹ!�i��@�	��H<-C�kpV;H��.���
P�ߺ�K�d���b�j���q~ =|��۬$+#�O6?T�����	�}�ꡣ��6�����? �ױ�nNz.�G�sL/��� �_�E�?��^�����f�t�}T2��p��Ώ-G.O�s(����ˢSr���31+ .��R+�g�_k�|���E̗\	<��K�쪷��N�q�z!�wYJs����/��۲`���~�цo�G�wjy�:���#�.�|8B5������^���D�"A������_�I��K-e�b�+��u5���
e�ʰ�L���>�O���Mfd��Y�2m�hE����14�O�"���|��?�1�c|���2R��t�K�u��� �jh���+]��ݚD��BF�Y��<�@F"��:Ą�U0]�Tmuu4D�m*���lѫ�)��J�!�:�~�b����)��V=�9���k������V�����	���ԫ�Om���-��-��H;��B�V���O;<+?<.�<Ő�p���k����yj�c��Ō�W��B���}j�	�*@<G�y��I!ˬ$�u�'j9\����..-?�{�������������C-o���f`_�ٮ�7���V�7{��R�oJJR4���:���]��J���y��ǫH�_�$p������c�[�A>n�{��p������wԴ�-_��/`�"���\f6�d�?�Yr	z ���k#e�B8��P���\�#���"xCQ*c�JM��b����A3{x:*O�3��/� 1b�k����	&�IK�˝���|]W��PP=$�ql(������\'�d����3�n���uG�H;[:� �~��{�ȣȊ�D^O�����C�e�2|݊i���b�B�`�����Z��I_�܊��:�����u$�e��Q��dƠAa�z�"�.��v?�i?W�q;*'�z>��<Ūn�Kt��<���E�e�E8���O���쁂�Gb������Xd��U��x�/њ��>�?sv]����.�\(���&p�':�̭M�ׇ��xʿj��[|#G��ޝJݛG�A^�nu���4�ꚉR }"e���[��;:���{��F+Ԏ�9B��k�ly�2�_��튓�ۑv��>���%׸�C�v�������u�Oʿ+x�l�`@�2]��l��å|vP@��N"�ɿ�-1����r�'`�.�T�8�����5N5gR���F;=��i��Bޫ�CD��9����������=B�Rt���L����{e�X'��i��Go�{��n�6qE
��\��`�|0{q�N�\�2K,�� ���5�_�ɩ�1��!3��k�"3�%���4!�%�B�0���SL����$	�=T��-T?��H�l��O%*e�xnF�8��)�H���	a�����v;g�9��Dx���F��1�D,��֛�5�"��A��&N���4�����M��$�7��8�i A�ǙLM�+�Fvȵ���8�;�y��A�2���O��4j��ti�:�L]����2�|z��DN�|2R�˃ߥ#�e^e?ʸ��8݊�4C�8�eZ�1�r�T���U?<S��b7F)sClKA�a���Ȗ���q�P�S�g'?�:��8�i�нp�L�t��Ǿ$#�XSפU.1�fY{ڪ�����ݟI�L�Z#C�s�`P����K��MHf�M��-�S���A��}���!�����K�5�bd�t�Eq�,p9�wn?ʲYf���^�VY�H������~�~��!����sB�K�&QW҈���H���y���*_�ݟ�}$�듓H+/i(ŷJn߿���ļM��<� �Z��j�S���w����g*��z1y��-yu��@��*�g�S�=G|���@r��{W/������}+��/��h���=6��Y��~a�-�
� �(��ۙ�/���Ie��(M�f����/���8���w>c����rFo5��$�_+�2���6>Iί��.���N�n��)����ٔH?��-��z�V��y:�0�4�Xn����	��ivc1�'hL��y��:�Xy�ϸ��|��uzO����nzrE������(��jg�!�K���YC>��v��[a�*�4@L+b���G"�[ 5g�r�5��mUZ��3[҆��S��#�BMU������}��J�y�Y���L�9��>Hؐ�:k��U��z��X�P'"������,9��	JAc��9�hvHĥ���
4��%ؼ�7'������4!��J�j� �����edQ#a���Q�	@�a�?TL��5��F��6���r#�u�)�xc[1�&����z�dV)m6ɴKIK��ӯ̤�G�r���_�9�s6?
Fo\�,�>-���j�D�������YO�⌊mc�r�b�s�Ʊ���{n�y�g+O�P�4 ������f�"8[�{��E�7�YVv9�5(}wγl�N5���e	{���/����<,�<������MR�4R���t��1K�c#�ΰH�ʐ3�Zr=x`X	���d!{ze�4{�˧���X�������OM�L��\fÁE���"��3O�D�P�׆=�֯����h����h�>��n���kJڃ~�`���Y�1h�۬�T]��|��$���w~�
>�DMX9ܹ����Z�ˏ�q�}cI�����y�״�;���rJiJ`,�y�Rx�h\�>�'�z�vn)�韆 ���'J�װ���@A�$���c������n�Iim�B�����£@m#�E��Mr������|�����+��������!�iv��4�����7&~���h� �&��k�ty�Q�_N����)���'\g3��[�rz��h97f]Ry ��m:e�
��KM~�O�fш��!ަ���^٨�$����,�eSneʕD�T$���L�&5�Ț�?b,���ο�Ց�D|��W��>��ȿ��]LEƜ�ث~$#�=ŀY4�FW-k�Ä�+�W�2�E����js៓��}qJ���u��4gj�A]�ʳ�頖,������/�Q?��l[��0��\{I�*�[�V�Vm{Z%z�!�-���;W��`۪¡y@�]:7�p���~i����j3��q�ܳyO�$��2�4�"�%U�kԪ�uɣ�zm�����j�I��Pa)J�7~ad曇��*b����)�4VF��R����A���|�@��feF;؋,�