��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb9$(>RK��N��.��q�tS�LfN��7��y�����U��lz��5�G�Tȅ��&�=���a��W���9n�l29@�Ǯ��|Ŀ�t��4�`�j�MSJ ���`�->FۻƜ���T�	lU���ςrXE�H�tp7���̚����v&l��<3�~��D�6�/��crb��^�^�9DX��.-�\K�b̷?��I���Y�֗��TH]2�{�Ӟ.�ž�ZM�`-K��
&�&��Fex���qJ!g_V^��n"(ɺ.r�2��|T:�e�d���Hzr��p��Fl�|�6M��
��A��r��Hz�=��D[Tn�#�OKD�0bV�8�X�a��ﵥ��Hl��D�����Xh
����+I[O�_��3ڤ�u�>LΌ
O(��%48�<�W�=���p|�5+ڇB�I�õ��{������UҨM���Yi%���{l���d��kfV�v]8�ѱ♸����9�ˤ��Bg��Z����΀�/1�c����
���ҡ�#\J�L۾	|�CQ"�p$���8�B�i3L�,nTHu��E�L�s9w�+��)�n�WA�{�yU�O�Pq���S�8���cz�.!�91��� �����4,�9/�*}����=�H.��n诛����[��J"�8zO>Ŝ
��Ѭ|4x9 </&���w�13Ew�������t�Yp�F	�Lp����慡�ՊT�')9�i�#�i����|X�hѿ�m��^�XI-
��F&B���(���Ķ�w�l�Je�D m�N�T��v�^�j1<�i����D<��'k`��r��9V� ���_rT.%lʖn�u��LǱ��N��=��3zKӁlk�B2��ÐTWw�,3�Slҽ��`�t�ǯ��!��k�����R���4�[�wM����b�������	��4�vhd'�%����R��{�Q��w;��R�����aU�G��%�x�~s�c�v[�gWDEHH���xQ�aC�{�IL�$�=��.l54�h��E�p���@��o+M��YR���!g7Q���>�P�3�(�G24��H�2�Ѫ�KK1�#!�^Ÿ�۞��/�z6c�^���Y���blu�m��ٸ�)�G����g�ua��EFIV�̡�U�6������x����ז���>�i�тw.�XI��S�:_��T\wE�s�7U���x�Bٰǟ�0F�vU~q`���9cWr�W�m/e(��X�[��Q������D�*RoL% ҄U�L��a��My,�9*s _�س�(7B�����)Q���^�(��̅�S6��T˽Q�pvcC)���e����:( ��XB���5��u��8+A�d�y>c�-z��e8	�+v�� ��%�V��B���g7� ��m��Q�Ms�D�bt�} F��(Ry��Xo����y��P&���!�6{�����l
�V��/'�u�P�cw�I���o�������D�,�?�=��Д�B�^$O4�O�.z�����Vo(�m�8Ǎ�Β�O�Bp
�ڽ�38���Y�XX�s���6���̅�7$1�e e�����;xo8Z��;h{*�,[,�q��L:T�ԏ��Oή�P>�G�D2�sR4��~�?6J�)uI%N��}�(d<�ʇ�i���JRRu	
Ĺ��j������o���UE5�%�1�}�4u�	���)�ߝOI�G�#�2#�	��꫽����[������d͜-�icGJ��g�ŷ5�U�\�</������7��B�q�KM�8u)5xAP�r�Dۓ����t�Y&���ׄ���pe4	���J]e�i'd�ܲ{����O������|�I�@%��U�Pӫ9]�/�Q,�r�W�~*h���h�@���5u���"TM5͝Xk�n6���H��~�ҥ:�{�z<S�B�q�Lk?A���V.�bj��*�+�3���q8���~��Ҹ���\��;��B�0ޱ�dpZ���f[\���=A���f�������ڭ���	�p@���"'�V�MI����r�p;��־�Ww����ȿ��ѐ��'���~x�m���\�8�@9��ʓ�C�[����F>%gG�9cT��*y��#�9��I��� '%��X�.�����Q��os �ȱ���>?ɐ(
�s�E�:N@ɛ�,lf� 6��n*���N>�G�>|⃵�����m��,����"�=���ǉ�b��Eˉ�hj����I#	�^�UKFw�T�z�8o����N�P�3�5v�
�c}�����%w?KC�1s|�Jt3��,��F��^% Jކ���[�oKȭr��ՠbʻ����TW!G���Y1�Vk�B��#�����Q�#~%$��> DB����q�A�J��ʶ�y+Ȓ����,&̝ٷ�rա)�v@��CQ��9���UT�G_�s��G$�g�W$oP��m�������@����i\��w� ֱe����G��{`����A��<(��h.�L�v�}:$�O�
��r������apw���lĵs[d0�.ve���a�@7�M:+�(���������4r�#���݃y��+x�/�ߩ���k{���n������_^��qtA:
����-)�
B>R��naח�_��)�gS|g�pê�i��Lee��mo	�x�ֱ#�_;ڛU�9����cyo-ŗ��a��fC����d >?�l>���`�T�'���nG�<,���K�M�{�\��'̩q71�YkS.�.u�.A�ڰ�M%C����`bzە�c�+�Y���h3
�30ə��[�d�ژ@�lƘ"��FwYb'[r����*��zU������sg����Vǀ�_�X��v ��B�P�i�Y��[�1è?T�;���(�%M <�᩷�!U�hb}�l. U�N�>� �G�,ɦ�;�|>�[�_b�v:�p��# ^]�&�qZ�k�OϿ�@�����C��{�Vc��0#s�w�mTG
���	�M𖫘?j=��ޙ��m�p��+3�c��|k��z�h�q�M���C͘^�z���X_��HCt�A�ֵ&�iAK6��473Gpj.!�2Ip�\��p�ݖM�Xp��b������ɜ`��P1�J!����3*a��ߋ*���
��6u��{X��4�Aa)2s�F(,��)i%�9���95��6k{-͇���i�%&��Uw��7��
c��XPE��/��ؕ8�M�:����en{ot���D@r@!��P�c4]��@I���#ߕ�F����4D��H+�1=���ҹ�Ѫ��˶f��Hv�I��n�O�9���/2q[��j��]�]��yU�8��H��`	�V�ý�o�O`�c��{��_˧p��m9�j���e~5L���A���aYj�禎�ap|I�?+{j4��7Kp�\	$��SkjۮDз��0�4�q�|���.@[f�Q����n�d <k��xR�z�<%�P�����O�O�2�яJ��Qm�vn���H��	&����o��D�`����*�d+�_�� �z��^���s�d�wGn�!+;Ki����,���)�::;�IH�l&�g�Im�89��������f�"�'o���n&߇TFұ��ݩ�tD��~q��s���=-}��ި���ةcl8���#�<n9K"Bہ�n��_5&vT�+���ڐ�R�メ����|�p�o��������j�cx(豱5��,n��l5�b����z�����gEf	����33yX��CW^�۠۾�EDA�?��8�}�6�-������Z`����������&�G�o��^�DzA�m�)��<�/�9`�M�sj���@؃|��X۫҈pxk2O���a�ɉ�V)�L�eH7�#��]�߁y���Eh_�?��q�MA��s�����z8v{x��bUu�m��yF݃�K��_X>�ȷ��	}��iX�,0;�(�a��CZ���>�|P#q.!�e��Z�d,qa˰䭽�V�!c2D��I�l�g�V�VD7ű8ץ�X|F����."�P�[Hy�����2E�{�$�r����ժ*l �f�O&,��6�#�%]ض���CDd��s�fo�%�' J�BVxN�r	��d��d���Փ-�K�q]z�N����xQb�_N�2 p�j�#��U����Ksw;���b�`W�Yˬx�$S��