// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:31 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BVWp8u/fcpS2+wzld6wKJaHyaePYWsWdJtxw+mtMt/inmDHm8doT8R0cp2VRJ5Vm
8iDA1LIC0I3VpP0IO/Liefh+GNv39lVlpbFE4EwB9e1RF64pxwkflJwU+FtFHGOw
TemkaybqOlzWAmq5dzxs1cEiQM3Fyi2S0yRX1ZhAJ8E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10608)
GZmQ96oZHT+xg7psX7kvgowSgV+gyK1ettZY6imMjX6/nQ1G84nd4hmHHPEBdVng
YLg1ypXzADvS4Vv1aqhburXCzrMmurdr3TT+fLsf0FQo0TecOxmgPnyeETN102ua
KRlQa8xAamKqcc06liAUInd/kotgF4uRoVEl8SUgDhBxEt+h5AU8j7x8NyRJ+MIu
yDfOGacye0xRu4XXiulANxMkbrxN+Eiun3AgEDIhNUFCHeR4H80wQ0W1/1GJy6gc
QVNjGORAuxNvZ11ruUXNmYYdbf3ADJvr0RCYWFRwx2WR5fMUhO6qqrnMz8bhksKo
oLRYutDYDU5E9H4it6b7YQbFbBE/yqGxIStAMbGF4zYujRsxCfNcchWveBiCh2Yg
cK+WGaYXLuNApdozawJGGZk0+BTJ7Qr9A23t+UzzneusC8KB6zhBgYIRAGIcaGvZ
SXdhXxa1ncnJfyTspAk/csJzzoT0gdBVCavjERc7WZcVvS//YdnsHoqW13OXPahf
9mN7f2QKi19cCgTLArdERp8nZTbRP4VZ5nY9HQ768dvcONXuTR6PBlF2LpsmHnWs
I0BmO3/8G1e7udA86Y94cZOwBuU7NZq4o9ByO4Orflc4WLqWvCMtYmFUDikN+Eo+
m0gfzRbz06Sd0mKQV4cIwes6dg5hAOVD0VchnwxFqnf2oJ5hW1z4xkrfcOo6ij2X
9+5lLZWRXIEDCC8rAAlgZLWAphQbeBUP2Ro+BuHVnlDee91weryn9H60e5QgYp7D
xjpPT8Mq+/1p+Pb0vYtLQcElEwITAqs8I+R613nCh4GZlR2X7F5rIJN34sK/lJD4
5OXXPBoBRpEfYEm2rX/csmtaODv/TYZWNv9kpStjE7RMed2pl8qYEqHl+l3vvHqb
ZbOIUc9f2XUQsDS3SQruIWfFUluEhyhwKNtvco5BbvWMKXG5e3602UW5DFl2wsdY
xFfUF98KZKpoHCdoWtY48f6P2OSrP/zOlF5sntTpyQmFrK+ddcwRmpg3BpVTEEtY
i6keBILM2k+q3Z1Uo86IOoyT4n59aLbx/yMqD9Yhj2nv32yC92vaGAAI7Xlh03hZ
A2r5z3XBioKSyRRVnDLNuRMbsHvfdn130wEgonOUYlkcsJcAuVbsGwDyfBMuhO3p
5GkECRN+maeMi+IXT5zWJKJi0yHxOA2u1V0u3wcXFXoMWBuq+QpexSM6XLWEUVOo
5/nQyHZK+lUGN6tyVICG391Bt6+5GeMSLEXEKscckjk+/P5ZiJvdbWzyy4YnQwIK
ikwKR2DxUwiGhoG4VwlSpPugMpngyobmXCb4Yhn0fr5QQD+3a1BSE7HTOt0uaOrP
AgRTvtw/lTvwGl93TuEX9XU6PBPcqwLCRgHga6kVFhU0YQAv1kCgVWCvaV38WVsq
WkLkxat3QibY2AXOZiduylWPF5za4btCfhxTD8izLf6R/utKmC+dxoqefztOPfV8
mP7FJ/FjsEiL2xK+aKtEoiFq4rL0Ly9R0zZTJv7frYxXSKnKJXF10/WdniP+O3Ys
M1k3phEo1bZrgbYNWBjlS2apJcwtDR2K2Ai8aLftT2a2SHuP6cr6Jcukps+EOd0N
3Mvzzt2zV80JFaz5tzQAx+WJp7SUopg9z/S/ohtAFH/NHwU19sIB810yuug9Rg4B
hheH76oFZdgV86qCXQZ43iPtLAQ1kBR+HXOUoxG+2pBmMlDEzmm6MHCJQVimmdh+
fy7updjoVa4FVfa47Dxnb172Vph546p7+q9niannLEyQX461Qx+Djg/OhNIXikYI
DxENLA+tThzxxU/gGBImK0sEmI41EWEMKouXZEghBOS2ApL7jl1nlRLRqWozo2TY
qlOk5+QuDN2eMZP9PsqGg5LnUSzrDM+prlG3sgAuAtk92Dz4K0HjjeDga08GcizX
4iMWyHoQm6JQYO313173+9USMyYJbeGuJAzMD3zqqGKgBs3vJzjLVtqXQ6EwWnFr
KTkgvlUYLmuujRgMaxIQx2NPEEzzAfvbRiZmTfqm0xhuAvS11FSR3q2ho8w1+KNb
Q2ZM2v6+V3BqdUlXMroEZkDNSOq9PcvfwkA7nP6EPZm48M2lkYVsLLqL/mgRCheW
Dp7Mo9MuY/CBZ9hqTJQaGtBPyzJaQku+qy514kRH07d1TaaT3HcYuHr7MwQc1xtA
0Lpln9NTOmiLfy2TnJ4DgGxotcc/G2uOQ5oz+2auZBBQVn/ch8TKYoItgYqdoU67
QOgAYLMEGVsFhsvu8f0BE0G9KpJ27IEz7p7l91LaApesE+QgM07cx4+yZe2q0VUr
LCjsfMgytAqV8T9+MiR0YMFXYHdqzR+BBPei+IvE5Ywx0gHwjbxreTCykzPxVB32
ZYwy5aFpCRCtLCdO9OUCS1dmY2czEwkLBUZsXF/AT/SfTSB2/StFrglsu36/GIPx
AEZh8Kxncc7x0XLnCet4YnWG9aQ/1wQ9cdm+WKixTRFpkvuQ6KdpqDXN9dMc2PC2
wlTXzxl72UlEoAyUU5X8l4HErITCPDJnUCh3vcyoq74S0lR5HNiH0b3Feeg8OiDi
tANXOAnjPkndSyKCAvBQGR1HEj6FhvNXxpSeK4RJbnWFYafrsu5anQ3wNtg2WjYW
dpogsczv6Dbti3LIvx9d7bOE0bC4uZfSZKwx6P0zZMxoHqWUkjx5rikSAbNzakyJ
jngQu6Z5YAW4FkKTjAXMDpCX/ND49c3bZdfxxguJdsDoW58/v9eRA5EJeHJUQMrM
YRNLxtPSAyMz6Xq1s+DeGiOdfj3UKf6azaTuuGd3pMaYlq2IMdI3JPJb42M/BgVf
FOtHc0Gh4ZNrmU+Paw1QdtZGjsIEoFm6O69slN51UltMa5IoxYyyPmtSuVHNcru4
v4d9IVqBxK73lTI1zSULPJCnBfX3tW7WQEGwsBF0mkqiAgFwH8T0MyztqYeb5ZYE
dJ87KP9s7WWka80JkKi71xtURtwKGnWdiNTD6A2KB8GHftj7r/JNWUVYpsvltPfU
6N42JVVP+ajrILT+Uuk+ZBdeLcjnehKDXYxsny36ObChbbjSWKKEx4XS1d4UJeeV
kjbIGTp9eVqxRzXwH6mbdXOoBsvgMXkdJkoK7MMuStmRBRTWWEx3ivOx3voA/z6E
u7wTGRV2TtuTId+c5Pg8ag7F5k+SC+yxuOT4RegJ3zCKwV0usA2D9Cz38kZ+CeFG
C6YtaD+cVFomXl13YaPwCnAdMt/DDkcWRvKgabzIw6AsOAyXvVeOWbAWE6NAiOfW
BvKtmuybBTKXfMrjgIeqAFJP6YYvt/AUtCOSB85gvrph5nXuTCq4fRBguO37CRK+
Z94BCvuA5yivStWBDMY8mFVMTU5ZkoaExQtli7w6SZwK/xd7jzBb7VYBrOTofIPB
B72otjoYyvRinfwfoVcJvA3RoSQYhsubkY2/hI6ksCnUxRTCaQ3kl14SP96Z+VqS
64ikHw30VAfik2QjJVBxVmpBAd2toRyla9s4krTWVbVsXpcG6jx9aJyAxjx+O03I
yZKNVyVn5/Nx0q22J0r+wICBai6W2gYhPCHp2sKXGFhrBxtHbKOyhoLfQXY64Fnn
MZF0Ys8hdzMVn1WV73SX5j1+FLWt1cV29az/1I0sXIU1d5qxs7rawKl/j6PV4gl2
dynrjmk9gPwKEdpg8D8ZXDz3gX7DoJRQrSl7xTBkmbXijH3+x3q6hRC0H/lHUrj/
JSJdGwWkI4G1PVh1+wZlaKif8IgGGRxxsP8FMJgKyCyeYJyw36kthOVQeZ1LlvP1
1SPF1XNSo8QlBRwxnBvLNv+IDWOjFimmP4923XLe/vCqJr9Z0jj8CnmQ0utlkwdu
cIEiaq9c+U79UgUTZNOz1UDtYnCSDg9CJ3ediMqtIgZd+V/VLljpPUTiI//Tumbf
KNcs495hALeY5gS6hksbbRxILGFHCgZBrRpcadkV89sgxdCIHI6AqaK+nyQggQm+
3O+js4/VtDD1zgQu2TZBVXlZRF2t9OCQCHQaXjaUoQbD7OO0gjDLzkZ4fBdjw/Dr
mXTZJu1iWJrFe8Ja6COcVGUpToJ2PyoPAyffgToNpp6xLXckuMzidnEAfmXhqY5a
+opeWMy+mbvrh4hnaceIpyqGyWLExty6/mAB2yrr9K9qQZwIgdTqRudKpA5uU522
P8k6h+U/2lUNr/iBlL5PFacOYNcBvt6vpX1tX919YyAiVwPuD/x32qA/3LihJK8m
nqyf9NC6iZJjj5kbZYQQN+HQA/f/p5cxSEwveye3Snd/kuL8bd8/zK2GHFfTq/w6
f3p3MZT/a/4/WRpkTKjfOtk2xKahCVZBxc+Dx0wODYe/ivbUtgs/C5pPbFyxwDtf
fgKyopVLY3DxHjgDhJaUsAEwZyAC3z4YOCPS6uUR+AB2F9nXb9a8AJi1E25NKnwF
QjmBbP148640R8TNd+uyLjrgsgBDB7uhRnTZxn2CSiaCO/Bmofjxi42CEar6/5Db
Cd4pbXeJ9Sq0ewiNMlwfo6i9jhNh2AvZg2bFJOB4wLAeQE08YzKLlvbaq/jDcsKV
MKI7ME/uBe2+gRWBqFoy7Gnr294cnnnPuKOHcUbg0Lb4xisPNAWsOpRWZkTU9/S7
QIOUmTXln+YCfgWJ+zN8lI5+3Knr3rcAYrebfEECvZN+4a7D1nPwxHV+X+KUPLcP
VKWtu3drbG2m3ZPQvuXv8hA8SnslYbmO+tCrTUJQK/SOSi8x5LyBeks4jInBseXx
Ghtm79ntTrN2yT6TBRBMomut/3t/Tg5JcvRHiPu+MqELGPX0HNQOTenQ0k4FmttM
0Go4EnHasGGujgt2aHefFH0soMoWAlmt4XGy/94eKtehoSeWBWr+k6hHuoe87a0B
62a3VaSCkPD9xd87r3KLKrGFo9Se+9YQpj7Fj/qcb+yxMzW9zehnyPE4Bo7+0KuN
REpSMLTF9sVggvHA5C7R+PTyz1ysu6Wf5puV8+HSusDI6SO9n6tA+nr/6GULBADD
MGA8xzpzoCMqd7OIe7T0KEXDtqCG5UU1E2VD2nKwKba9dJIM5e1xiHOdcsr5ejy7
dGfhvJQ4yz/6WNsv1sPLWbC8NmJ484zt3Fd+hhLj8dcSvduTU2JqkZ7h+mWTJhso
tJrzWIe0mkqUHNDEi5vFPz6tRFA75GQUmbYWnmsX+qCkVbwyNuZQ8grBWnHelK1z
NfyUbr9KJ9WCggsKsR/pVvalTUJwo2tCu/kCnfps9CqkZuCJn2DPvCNuusM2nf5Y
JbPMPJjIcnhTplbWdz/TszG8jzIbVt2Oe587VCJ+qnZJLhucodevpaTEQahtPGe1
e9p0yFWq4LvC2CzACO6CczyU8v69FoL3CPvs14SmKcZPEYPDjnXtp+n1ojk5ev8z
PUggjjS1brqg9v2tMwLk6otswXOtAntpdrdnSx4g4TnjkLerGFpDiR3DG5Yqn/V/
TyZOOISDQhBTeTuGEqlOVyTDhjL9XvOjgZX70p5jFQmYaa9yTcPYdwufwYK1P9D8
VwaSBuqaaZv3qjX68VMXcrIfJzhn4U52JR7c7giXZl/sAIJHUNIWSwBI/xFcbYss
1RVw4Xf6DBkcv3hzs5YdrKjilQ5afO2Rn2bjpdWOK9kESDT/QkE28dGqUGgirtSo
z2HUyyyndqgg1kYiOrLJQVyo/YV01/Qg2kerbpKscQ9GvnkMztLC8NzSCYAFtFR5
FEYt44qd7OgMH9fxfpmt2SHzbvBS3MqEbOJJS0gOJob8+EpaAeBXMfMS6ShvEGE1
5gC8nknDFMA0+rMfGPkSxEwjPfxL20ebHYkHc0NHcgwy+EHZ6UI9kjyLAsOtiDrm
q3Vbn1uaBJll74CYOU+FKGKCmGnYKYNcpEpVS0TBPvvQ0FgxQxnQtZ9AMtOwKTiY
p3Z1hZlcDLvwMqhb8hm7qz/mTd/h/nxtOtmyQFK8833q91UlhEbY0cq0Its1+T2H
Lv2da5RsXrhv5iEhBOwBUMuO3N/+n5MwwCubn4avLY5DyYqCe2idPJBZw7OHLoAD
urcrKy+HOE9UbJVdSeSAN0m3gVGxzrFdhY/GUZ2uRlyf+bjRmI4e7Zb80qhC7gTM
Cdzg28F6XO7bMcxnuhMPspc1MVEAn9f5AWuHF0aX/CYMXgmXDpje2K03ocsZLh7q
s0GV1/BWYKeUU9cBGUoHglKT5z8sb7CZ7Vvi25mcd8EXApVlnGLuHWO4feQQmxlJ
7qBCAJLYHrcIAUjO49Ty8FiT6QCUvU3VlwRxEJJldXrWuWR4AvgNtq6TV6xhGwyI
WwBirVj5upgd/6VcJ9InBecFOsGqRYkyAopNv1JdzjdwoO/C9PDtWkmnLz4BIrQq
ML9XXglrHj8Fftesr27cZ+w/Ku2oVnLNx2aN1toexr1/2nlco5y4p5RaacMcWGsS
z7qkEIuXGNl0C4Aa5u3WNZSPF69WolzCSwFQbbb8RfGzNYA1tv68esZ5ngwwIQxD
5RO6PcwBiaUXgmgr22+5effsIIEhEv5pdNOy67twds7GgZWeVACgXUfHzIA8/XH6
HvxtS2sbg8oXKTRCpyzGUvEKxffjzNPY1ib/dlfNDL+WZzatX2mjXi9XnpUybbhd
ShgyKyzHMzjaL3ERO0lkhjrcWqpW2oCHcvdj3lD6pgDnwIwXN05JJECozR7eemkd
SYByFHFa+G2o4pRVAMZzpPQJy3x6mh5c5mSpY4W/fVRz55G/U2O+14SnfKMdnIyB
gjIpbz0qJy22qgcwefq/nTe2QDUUx+KPmyfVvTHGMPG1VDVZMa3/36mADK/rtxFW
NSfC8Sz8mB78u3D5fpwpFo48P/YpZ95f3kHY1QvNd73EoU/9JplvISQ4s+AWGcSv
1xUXgfQwxdpZqPPJ0P9H+kK/aew9tcKiAXASWJb2AzRO3TQVn5rxiixgwpIlhar+
l1KK0DlGFpXqcuX6ah4wgGtgG48d8RrNVU8gUCt8VsrdLVtaXN20+mC3gouCdmvt
EFnutKZQnlWBosM0GGD2sSUzdLr6HndPpP1sTDxgtkPhwY+wVB9ewRTqoxVavI1D
+Bnv5Cqi4heDPKf5g3ZJT/PC6MXVxL/QlFpnnzygupuvW+Mb3FhuCuHbw9+5MKRp
IeeCrJ38AvFnlscDDELdIVwtudPTyCuqLg0Ie+CIjH0YGfsi7lLbeNwu6oW5PL2H
5iYYf+7pYV46E45R/vRvZuePkurvDXIf/g4Cfz4CzzJJ97XjJdKRDpj4IzXyrQx+
HGvk05Gduiij676V/xzb/ngq8hnoSNCczbvzaNj21EzroMmj1mbSFOeBg23a4n0C
S3yC3FtBBnKzGI8OX3YgRnpLGO7Oq5IKyVWpGgfjXWyQhDjaeLovAc9cKYfaPozb
psRl6JYp1WdoJbdSzgAtVFgmXTWQzCh7bQzFL/PFE0UhGrQxcP3N1qnKo993hV5j
AuhUvR7UraSnGSKvi1yADLusoloKU+ziSG112Lh5qWqs6O8pqYwzPvBLEg5hIf5p
cvL1ozxCeOw2tHlAn5YE7c4+tUfRiAxKlZyfpskpKNYZajXgk6sK/Myu3XnSSMm0
SQoYlnxNXhnDNHajQBztxw9z20rdoxNmh+x0gPokdvXzNykFOHFtZ+nl39oevftJ
6jlF5t9KyFbIUlQ5yw0H4HYHz09Qu0rTep4eIqtMHD5oRlFHqqsHivN6jNrGjs0v
2gq18GMATjCPVtFYQsK2SELxZ1gVdnLpn4qmkIKxjrVwr25AVlx1yTWC0MT2+J9M
ppAVgiQDfynzvS/AzGvfS6KtCIK0wwIPy1jsczIAnBdVwXcJquTf/qxfVeJhQATb
N6lXVwlAXJTFZtRQbxwAaJvY8NoXucYjoArC4pb1iUflDL02tG3ZJVqEn34jsGAW
O45ug5VOUfPIXde40IKLLDp96OENRS4Mloc4hPQBTdWqEHqJiICrX5DMIGq6ee33
OMGaAos3DLibfFWn8WuokOSbfE4BDi+N+Y6WVgoGR3t5Mz5AQy1E5h3kGxNgerIQ
0wPX1F4C57R2nQHP558iHjYdtW9WdCGgRxmqtYtNRUF2eWHbDLIIJ/YGPmhG2iBO
VbgrGH15RfBXPUo6/nW1r9/T3l/92mgZmNAC9KtYJc4WnJdW32f6bAD0yl1yxXuO
P2robuibLWp9x8MQQdJVwUtu/dFycanM8vPo29h9v3D33MVtBGi6RdbikvytKGIg
C4KFKQ5wciLV1nMu7/2D87TiTpfLj1lPokelzxFZMsiFZ50nV660J88S2Iu9wV9U
OLK52XJZV26z38i4YQc8zgYYNz5535tSo/sUP1jXlxhQ0nUVmV5eBig6i7RT1Jfy
JY8IpZ5shnwlOEdKvqppH5rtU2VFmMlAqp/LXfDj/lUdAuvyyWNE8SjKnv+cwVn7
2qtTxuCchHn8DCVuV354WG5iWXliP1oBaoShj+7dGm/k3taaTYRlDGjk7Lrxt54b
3Qha7ddLVOfLmcWfVGaULTEPyU6osw8wP3+KrYsbisglL6G4u43MMqEySepSID6u
yuhbtap2o4Y3lOejsjXl6mGt0C1doCcMQAnrKlw5Z0RL2pUbvGsAqxHFhKIp3cuO
SxiCkEbJeaOaK3MpetN0P8GEIKScttsZGq3Vyg5GH+1B/95MQ3cpdPBMwwwzT+Pd
rrCIuTS5IJdUOcmDxSKfJ2jSjeDFQ5/JN/Qk91bciDSg8Y06gpyc1MA3WX2n4rvl
VjdYTR635SKi3wP/IHkZB4I4SI7uLepiaJ0Uma/jNJGSRk0Jve8megmQxHUfw8eF
6wzazM1uyGW8G6G3weJ2xvwv/ucLo1bWARgFmCChE5y/mqu/lXFdr/pMCFsxAFei
/Z3kpSVjunuwdJCGyn4bmxEqBz5Z38MA55GGlJOodB2C/QLIQBb/hkljApEafuHs
gJcAbnu4ovnVrkM/Qy9naovmrjZfvbKOmAuvWCER+27GHDr8opov24d9LfTb22d/
fdZ177fzlciLIhekjN6xHVUes6ceyJvRPkSvhkW+OHj6OzNRykTS3cIr+NnX9bxv
2Yh6ulY0669iKwllUvOwI27BTfQZTn9JrFLuA7X2gn/UVG2TN+Jbum6xwTOHyCqq
qu05VXurkrT4YZ5ZSL46J3TiRv424C/JUcAXjBV10dMf+Cb+3lH1NsWAXNoQczlK
gVYK0I07SbswIJ3xLxA/T56mlbimRA9F0bLcf8yAP55FeuYTFhhKxUIJVda7TkRo
QAl1m4YO7fDwv3jwrtUIw+fpXQ/cP+cT8afl981MGxfuGQlMygjyoY6+k16ZnN05
P4pAOYsIe2N1MsqOP9Bwyp77DORwijnYDdVLwSVb6+Vt/6U4wzbXwHQeBcwF3WWh
Of1imP0cXQZvUy228Xi/ONqjSKSqIs51diWhXec0Hnj5FW1k5vKyAH8kNTNPxS9f
KAm6eOaZs2+UK0T+O4Sd2QhlWfc8kJ6AJsdNUxUnoXcPRZGSufkxAyavHXY9lfT3
/KJAw1TdxGOn0ch1Lm7H3wI5Oa9b4z5nC4a6MTRj3K43QscMTGmje2PJaNWeEiDw
nbj/OdS/aCuDqHBhQfYtrSs6hoe+OM3P6G5IkCt2cMYO0UjMyIDkuPghR4P9Ha9D
HBInscuukDYKhnezQXQtLf7PFoz8d10XW1CE7fWbuaLMkqhdNw10iXERqlhPP240
Bqre3vqXXZgeU4WVrLLnY2c2K6Z/78eMFsZM808D5jVZ5bPy58PcOXEhTegivotn
BkZLdcm3Z5YMiO6w9ucHY/tgD7UX7LHK0F3R2RYnOh2hI4qsSLJvBOdz9xQm47RC
NRnYDTRk0HOWfqucKK5EB4lYP0L3xgxBhFpDeGEeX7cTTFVm1T2Fmck8pGOnqiJ7
g6tJmMXR3RBKMsItHczoRQ+vetP1MB1x4O8lbbs2qSWrVJnOauyzeUdEs/eN2Npi
ljLGrYKo5pj0Mgt3rLuJvdtBxKVWrt3+B7AB/9BsXxlcVR7KOYS/g8zD0F1/5AED
YvDUZ2BqUackTPyiGrYHnrOv1/g2Ufl3y37xbVcEtBdMdgCATGQQfM469TXKD3vQ
rL8Yp/JdskZF3Ft6mLQXzB+LDAEl5kpySUMlBMxTtNAjESw9UwDF3OuPgRt0TrNP
xKjmJ9x4Wbt8Gj4MU1kNyKRLX3+NJO4P58F1q5+ESBmlvgLy65Le49f7btJoSNzW
3TRNsaniiu6oxU5Ur7SPtt86+szNae8no9aWxY0KN7ppTNbzZvGkns3y39Vr4Qy3
nh34hnVzV0SSvCyPX4QajemrFCz/HEjreOvShaAILCt4zxnW/twJnTda8em0OGNp
2YR2j+sKcJCI6gnYLhvMgXOpdCSdEgnTgF7/4RKb4naSJD+daoHZab0YS4/W99Wd
sKMKkCPgP8cty2a5s52Hefx2DpeTae9hgGcFm7PywKzy41i1CxBnnsqD8h4UQvX3
wbjbLYh0HxS+OCNgN9uygfpvLO4bpqo2G9dfvSwsIKYjPe/ZojPVe9xS2TA5cItO
J8YJ4efqsqQcl+Vn1Yt3jthOllebfdypGR/buUGszh6pf35mZgAzS43yutil9yZX
ObBzCFdmsBYOlRhWUWeZiaDduGkHcZOrpZjjsbxBhLTuw6vrHca6LvHp2/BNNyzD
rq2VH6uzFzP52AXyJs4yj9fm4hvWrSbJv4svE7MJtmry7Hi+h/ow8Ut2dYDFPswR
IHItS4SN7BZ7moq0Lwp4rpaJiUMl0CS4Lk+G0MWuWXiXb1UXskpkLilQk8iHJw3G
GisjD6zoHPcXfkPHMn1xufD9xIvgFG7FBDJuvh6KQLpW7atjnjoKbgGkUO1OmmP6
pGyIZrX3lm/KfZ4LLL39FzZYi5dMKUsOHdZFVHOwtCn+E1qv5kLus+900OIyp3Ge
hx4Uvjv7CSaZW0SZ+lIqaxHwOBG6E6YI+rAvMgYVFVDvj+M9KCNycmeQSwqJgGBB
wlZmQTU5Yyrohq5RtFRSnZECM+RK+ewqb0f6qsK6Kb7Gbfxi6FUyC4xz86Oy3v+0
YPWYbDJ3EbyND40dLV08pm2rQbR+dhNN3/F969MNKaiNAPmyn0S/X2fbh/hqkN4y
S04f0cr1kUsVBxaWMsVrOBynwUHBuAaCLoLaUA2GGcbcHDXOPXVpTua4BgEZPhOv
kku/is86HIdyRtshcxO7cmng+MxgMuARgj02CJ6dK2yAPqB69GIcnITQ33zGD+4M
pzwoSp7qcL/oPSZgaddFX3E2XQwufyeMVwRjdeuSRrd5+5T9O9j3iPAbqzUXoE96
Wj+YaJGXota5JBbQRSri4C8XphMEybpZYRIRZjJ2qXv9KQXcIvof60BUB9Cmkkpb
Qiznu0jnBue/okPNBGEe8l1lKWcOz4GBDbsu6D6p/SeN5ouwO1cioJy77rJRxPXW
ubn1w5MWZnpRu/y8HffMN3KHhtrvPdvDWcqVvapvAsZSdWOLsvzwxQ+5h82Ok+9g
dqs+JSIju5OuuGQHH69RvC64ftaG/W4t4sN9BS4N/myhm117VbxH8UKM46WNEe4+
bKVKXVMV9Nl66aiYaB69EumZRWS7AetmLhH7WwxP7PgqqksKaOJPIVoTE/5kzzVc
7atHRy8SZfvTU6xWg4/Fh9iQg+h1pxjcTUKz09izw6ZP3RMeb10ql8hpH3iIpgav
0Bfz758iiRfP11k81HIit/sxw2cuKTjHguaHK0iBn8McCvH/W/dPA1IA6aytaeEQ
jWKUTmHFoMnh9z2aNDdXH3PVEAAw9d2qlgO9eoyHbVQwwui7bIXTzCMnhiEbiRfq
wpPFqJgSLua94lgBuS/ZpVaKDSeFIPDurG/qb7nXlF67hr0Zr6z2qV7uEar2sxco
4UDfLSfKacbzsNuvWt5frgEbWz96eM6U0wkzmfjpk/ylrBv39IiKHQ7+1lv+IyIl
bvewvspuTwjrzr46Qy+HeTb+bPpM2U8zF5kJkjfawIT+1nDctgzZIJeve6LmREIc
oLd7kZX1LL833xdbVwK8hCq6W4cbHU3yxFNhdy2BLurUp8pR15yg27yhgnaD69vQ
6v1yT/r6yXdhG4h+8Csrp5eV1psKYF2hoCB4Lw54nN+la1UQ82tAhEc2br8lNj+s
mPVIC23NwIHyabLLkzPUWAVrbW1clbc19P1iVYVuGcZIOr4OfulnU9fvDUYM4zMM
7xuTyo2FFB59LpzxQr7lMaJ97niWzhce6Yuaq3LvicyWGQqC6IWS6fI/hex7dVmt
L9O5JE+NuuJufuyqJyUHUqKYjoYg4tnYH08Qi4cVZJdGzGu+Dpo633ytUfBFrMGF
PTdjZWP5waootnMLhh9UKh6AZT6HnLQ30fA1FhXeX2SbXjv0ZGQ1oitFQ8l2MH1x
T6KrsklMT8/qy/pr79n7Qw29oZzjhBgxuSMoWnr8xptpEMaSh/8X1s6/Ls8oj37Q
cfvnxJjLCgrJI94B5JaB1qiuOSFH2wwCJjeayWvomUxCd505EywexPuZpweA5nd0
AOjfAfX37eRgMx/4aCzAF5GodRLC5HmzBhNLhlRCRdrHFR4nfIyjGrhPP3mYs3Lw
ve6PRnuFw/8HK7hcvNWvHQmkwi+eHBoUxG0+ZbkE9wb7h9NRQuh+pML5abuEnQ5Q
47alU57o9XaOINayxUsZUwJyX2E5sVTBqN/3PZGcu+KsV4nrlqb/rcoXRFbugx+P
s4GtabBqsuPn7rcLUsfDjyRCZHBzUNF8bzUImLRmKBnAfeeDQgsfyYxkvpl/7Ntp
OFymCChOnqUS2XDHhL0M35QBVNDWABQXTPotBIvtOt08xZB+1hS710ltT0gp7VgR
s7j0uIjl1D5saZmZi7Y6ZNOsnO0TU+wjhdfQaOQfwhHUt+DKXqvgmVG2pwwgY054
PFEzNCoTpAqKCXzHLmCKR8WR9nUMkizc+/qexWSYQOhHp1ysGTgBZiZlAEJDhV3w
K9ETAGnxD51NjrKtJa0e+xYPH9W+0JzF4dYmcAfa1Wqqf0Ct2snhlAOI2cRhK2s3
fD1Fe2PxHT/5LGhkgZsWLDga5O7df2DOZAzhUgOo857ZgiO19xt51YoXeGukBU0o
YnFvpVacval4kGWNw0C1ZY20hblMQkQnsw1NZ5v5ioQ6k+2qefTl/UwhDkN7Y1cY
NyHMm1Nf5CUbbUw/S1QIe+TH3fxDKTnDq7rxy6LMiBrzprzktYWlHCU6XRMrOQ70
QgOJtxG/10LLUmny9snZC/9butW394YQSjWFaJier5c2zYWQ8Idvfy7q17Hgtegm
Ofq/NyVGHeu0IUYwQ21T0XD/qPk6+RqZVsrcxurz18TorCUina1J0L2x3wZiL6fK
O7Ns6fE96S/yzeT506a4P1Kv2AySx2rXCP7o/DPZukTaY1+a41+Ke5jho+IE7+92
jvdkZJz+n2s4/L+NoODpcUyS33wnBKUTnWCXpIq2ZrgGkSXW/nILPykvIYJDiSlY
Lj/RpWMZUY80AejfU1Xv3zQ8IL2Tl+4LRcse2FTx1CHHCz/uKoOiNVjJk8SOj9Ye
aRYnuh0oaj6NpFhJzbm188s9WqQfkSy0dEv9QdqhaHj9VY44WvUfcFb4Q9zC1y8C
SAdOJyrkiwaZ9h0O3SZxrgXwbGpZ5U/IuigY9VnqR4yU7CSP//INcm7OTC2RCi7S
QXkfhf1oagZheWmYVgINVX1/vfNEx7CRga8xxE4Upx2oNy8EohvzO2jKjFaPExKY
jhwG2r+o6drXUNkCOVdj7XVA8dBaUJNnglYPLk9CXmpcV7lpuoKDHY7Ps6e+pEuu
Rz7FoD77mpH86wg9NtnC4vbOqqrIc0wLi8SEpeYSwTAKW5zKqp55UdVVKmkSMusc
wASu4cUVlVB0SVG9MqvmEqqO7nR4aiDz/BEqxAiMqKgmES4IO05ECp9B30bZMs73
l9gPl0wSx7Io2zT/I70YzFCENRp0uVy03+jlLglMXvhSYkVeghjuUljKDhyR+fZ/
+EaKeHK9GDdewG+n/yxh3MoDC8tFEJFYTORTjaTrS/IpcwAqlWhDpyuR4lzllQ8r
hTIg+8rlu+QJ+xz7lO/I/0e57Y0hKju+S99o3RFVvA2FyAPwKftnicrYUxsziVr3
jMpCdn2tRIODSPwPLQa4g0gPHfS7u8TGgOBXwAhpe4q0ily0Eo6qlEANxEAcPYQb
`pragma protect end_protected
