��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����:��=3�J�r	=�� M@Q �:���!+��?kC6U�T/���&��	�bK����V��D�Db������V��yfʀIG�D�Cs㠆�.�`OI"��\��L'1dA_���%��:��c���'P���G��4BS�_VW�#�6����ZT�v�O�! Q1�fX�<o��3���x4��̢�!i}���IZ���C} ���ӣ��L�l�,��Z���#)GO2��ׁ0 ���_y��7�����m��n��tGo$�=x:�U���������3�YX�"}�ۋF1�0� �-3��{^Yt_-����W1�>_��M�-�����������&9�^�?�ʄ�BϦ�s�V�gW��ĉ�Y@B��9`wg������t�I���Y�<���A�T�L�Z5p�C3Y���D��N<�;�n6��y��S�s�ok�G�n���Ҕ����b�騂�
r�ҢҞ���ɜ&�uT]�<*��,]
�о1�N��.f�j�
\�Av���9�mͰ��o���-�z�Υ�d
�?�0iST�L�`o�<�7���o��Ӟ�)�r!���'�P5O�^Vt��3���Md��4'89�^$!7�HT��簩&G؎���\����gP9�	�R�{8U�-�z#�(��m
a���Q�]칥ȯ�"H��6f�uw��� �Y����)�����фJU;Σ�loS�G����C������@wEX����\C�����)�M[m�������r=)4tL�B@K�o&7��n{��� � �#����	�[5�ʏ1�>���3�7���h�3��p��V��N�vHo��?$kvjq� �]�a�A'�s/G�h����`�3�v�.2��1�F;[v�ز�1Wb��,�~l�sZ��H��%)� ����8OpX%���<./��ᢞ���C7w|�tE9�� ��8�__����[����%!��M-2Ƣ��Ka'0y�K;Z�[Ck��m���(���q#���.���۱/����YNhl� �t����m4�]4#P��_�}���b�xS�Ur�>?Pߊ?�%Fz���6�lkE4�BnX&qt�� >�28|�7M-�����e����	�|��ؔâ�VЇ����\�`�Ă��U��Y�)���]Um?�kU��Wދ�u���J�-����J>�����O��TI���{������j���F�Q���I,�>�يe�&{ި���r9{�vNZ�S��\��])R�:��z�6d�&=�հ�FGَ|wR���bl�ċƶn{�.k��^����F³2	�o��� ʑ<�u��bX�Ɯ�ٰ��a�L�*yD�[�ds�݅2L��6�χ�|���p�""ޅOR�'R]@k�>���k�?h�L�*,�>1&� �kͶ��9W��|J5�L%�C6��������Gܣ4���Z��a�p�#b���� �|�"�!`��ܼcyqh��qW�0\پ9������}>
���4�t���"�R�-;�k7�05v��p8YD���}�'�ԝ����c�k�
�v[J�����~�0۟J"�Q�ő��O�^Lw��� ��OQ�eN�>ΐ�F,T�T�`��E6�4�p�j�e"1j\�K��@�)�����@�����+Dj{��"�P�/>�^L������뚔a�D��W�E��{�*{��� Hyԅ�m~m��D��r�V�c�9K�$��5��O�P��͡��b��O���N�S���-����n��/�(�^LZΎ����ְ�J4ʕC����JXo[�U&�}Z�� ���6�����ćY
-]9�e��p^�9>�KEw>�	,�Ov���l�a�Z��V���6�f�1P�����vJq�D��ԣ2�>"Dl������*�4~ʵ�_Ed�^T��->�t���qg���F�dmis���c�F���=���R3�Q���e�\N:z��y��EYDc�M�y��.
�Y<d��]R��9���S����	/�;�DB�!��g�28" �k,EY}�.YT]�"!��TJ,B��Z/�YievI�(6>"��>�\۔T�W������9����{�O.yڿ?7 G$N���az8W��e���+�Q���VB�C��3�M~��1����(�[6me�,j(z��q�〦�}m�[�ν�@S�P>8�͜�ِ�Ut�S	�Y��(�?�59��N�%Fehsm�r�d����8�(��Z����y��[�	���p�Q	�����9N�Ƴ��#�}PT8���~�l^y��Mw�b���G�vfN�P
m�mf�<rI�}��C��52aZZĝV��(����3m����3]�C����������*�ע�⅟X��8kL����ZCg#*��jة��r1��*=ّ �A?_ψ+N~Rp�;�0���%B�_g5�Ȝ�I��
*�4"!�1$l>0h=zU�D��e+6ֻ��F.�y�Jr�ίv�cs4�	?�����e����t�r�U������V1:=����X�ɂ��!Ѩm�Xm��eҭ��1�n�doϖ(�<��%�de�E	LV�*��3X�_��(�A�pu*ĆX�g(��]���w"�fh�8j���l�Xr�����XҔ�(M)�[P�z�x����]e=�/M�g�G�-��R�{���Vق�W{j50�O$	�4�B~�[�
�t	S�V4��U���T��H��v�T]��h]$�ζ��� ���Sn����W��~&�F���wm��Fi3�ȋ��\3�����ZjOn=�"H�7�c鲦iR�g��ö��r��C���Z�c1�� �Fs�e����ѵ���O(�Wn p��V
뚆Ycv��W�/hs�Q�$�
��ִq����W���Ə��g�I�m��'��a��l^�L�4V1�M�Y��k�k��,R�I�M�����W ��0 ��u��<�*��t����&����������VP�F9r �3��D��z��+��bW*���I�P8 ��wWZ��۝�y(��a�*Aϓ���j��[3�Q�^�b�	Y��N/���l�#w�cHt���X�݇�2����?w�k�;l.�U}>��a=�H���O�'Y]������]�jS�Rch)�9�Y��ҊO��R�2=���4�n�C;�z���#��d�=����?���a<n��J�Z�H��b�|Շag��[$V�����w��-Ѓ�����h��m�R�CHj8s@�qx[��|k�(�
�F���Xc_�R`��F�}>S����i�����!b�<C0ʷ5��QN������^/�h/�˺fo�"S�Q2�y���R#+�Z
���g���'�5��q�skA� a�l{���&Q<Y�%���<�4�,��K��"! ��QR�s�<��q�^��B�-9�al'�z^f9
:<|}�����/����R�!�-Y **AjwW*XdW�)���DC��4�?��������ω�����7=�s^���=�tO��F9�[�����S��&�X��{�l�����x�.K�]��1���HPhr�ގ����VN�X�o�V$�"Kn�ϯC�\�L��I@��a�?�"�c#��D8�M���H ���F�=��;~Uw�"�8g���wr{�c+wS"��Re�l2��{d��߇+:��`��O�� �~C����TĮ�@#S��cb�;2��ЅȢZ�e�\b�w5��"���Ԗ���1JK^�]�ܖ�:�2�. qX�"���W������;�l�BC5Tٱs�w��A�6Z�y�:�D��AD���ܘ�c�����XjtB�'��ݰ&�xI��T���<<^݈�AN�.�"�kr>�����	�o'A�)��U�j�1��`���|���U�h3���G����̒	�3v��&�y�Ԣ��po��[�G{�HW�1S�
\���\3h?ɻ���\�l�o|����D@<�E�ʑ+�J�]�|ڞɣ#����Լ��vH�\e���a������/؁�$��-��{��m�`8x̉?�t���s���;����������x����ڈ��uW��g��;R01K}���څ����jE�ToO܃�Z�?J�0!����ݦet"g�BJLP����6���	���R[֯��ݳd�{&=8����i�`|[��-N<܍>�Rc�i��cإל'�#Z��7g��3��O���ͺB5�u�B�#>�?W��e����$���*�d�D�)��x�r�+�s������I���d���}������U�����1Dj�HV)�ȡ@N�>B���!��?Ćɂ��%��m"o3>�_t�%+<�l�Q�z�5|�F"P�Z	j�Ū`4��X���;�3�A��@+�)���f�I�C�;Sɾgr}���ͪg��4��>�u�DB�n�v�,#�]oN��"��ןy0'@؅7��V#���v{��z=���m�Y��^��J�q�]����|�n�=���Qj�?젃n�@�c���"w<�u�n,�#n�hˉ� Z�S��o����3�d��d{��H�ĳ�8�p�C��>�Z�Y�mh�.s(=�3�l�����/o9��߬��"J�#�M�	Ԍ�A)�v�C��`T�m��������y���~ʽ�4��y��U��)(#��X%ݮ/���0�K��������H�1�����DQ��c��?? +�����'����)q�(�7�R'{E���j���
m2����Z���l-�[��y�:�BˁyA˷5Xx:BE��!{x��Ɂ���t\O�o#��!F.l���2 Xv~�(��=�(W�1�p���K��=t��� ͝Vε��4�Mp�,��Y�ш��b'�:B_���L�rU�y�.w���O�u�˄U9�n~Z���UF�[�2#<(Lz٘շ	Z��J� ꛼;�3�rB���|y
��M����Y�r@+�Ĥ����>Y�}��KX�!�	c���l������d(��Ʒ���5ҋ���Qk
��̽
�.�"ٴ��}�OH-t���B�W�LҬ���Ƅ�da�O��ݛ��nM�ˈD0Kj���KR����T���������	5 ��I���\_q�:��UQ�!xϳ��~�t��zBp|.�c��H��t(_�����/�.�k����Q��!1$`�s�e��v��J(�qy�X�=�+��o,~�
>æU���"�r���������fj�ތ��+��D+ÙS��oWOT���ۊ���
�>p@	1�o��������!x�xi��9hXa�[PGE����~4g���}*�W�G��j@�[\1����b�����-��#u�a�h�z�� �_q����e|����,�InE��HX�"�)M��Wy�����KV�pI���fH�+��W�(�������~��c�A�WV�ͬԪ�����$�nQ=�Yc��;��ど�����"��9�LK.�����KF`�����\7V�UX������l��	���y�?[J��q�|�v�Q}�%�sa��b�yQ�f��7Q��CC^,H�k��X���7��ޗ�D�� y[v�Sd� Q/�!�)@��w��(�@׺۔G��;�*����
�����`�F�������#��s� � ���r!�| A�@;����Ie����`<k�H�	ȅ�ˑ��{T9|B$�țO�!g���T��A�����B�/͖�خ�eI�:���b��2��L.�jD�� қ��2�waK|S���U�I��7�F�E���>�6� v�!�����G�e��؊吢�d"Asn��@�+']��[��9ZU���0�N�l{4X(<��XR�2���J�>4R��y=wa݁HP裟ƍ��G�E�Oᢜ��4��t��+7z�����e1�ľ:l9����w�5�ZV���Qu�*�p6b��%�=K�����Q>MB]�>a��+��j�V5�ؽ�4M��g^�R��me�}�;��*�p������`M�:��""���GJ3n�A�|�K
c1�G��<��ۋ�v��Dq]rDD3��a�>f�S*Y�ڀ�a$2�}k��=��*�ᴃ'S�q����Tԅ�,qaM'�Ս���t�a/v���9�X/�Q��52��M-�Nzz���VЊ�;��k?������3�y�	�c��v��DBX��v|�=��	C����N��J|�]'�_e>z�F���
O��HC |���ע��LC1� ��yA�[��V�����9Je8�O���|E5�k���=�xY��trP?>�;�$�Oc�9P����p�L�_L7����P�^�8�I��w㽸��K4������ P�N0ՂJ8�O(g��捿+3�z6������]�N���z���x2k@߿���h���d���:퐫�9r��1�̿������rT�b}�X7O6��SPh���F��}�Qm�!@×|��>��x=ò)9�6)-cUϺ��A�x ���:�,��+D�jAaZ���ۻk�s���yV�߾X}uA9R���Nk�ǞL������<s_U�"k��q�z㞱�L�4&E��i]�}�wK���C��N��9T���r�w��h"��}6c>6|.�1*�|�r ��MlO�f�:|EJdPe"�r��r��+cJ��H��k�˦�Q���0����@�(���^C(��S�X�h�����U������"���?��*@���M�ŖH`���/�B�>��x�K�@ S���?u����\ߞ��"���@�T׶�/TV_�7�O��H�����τ�-G��- Y���H@�*�b���bp���~��wK��ޗMf��}xY�C���y�'NI ���?(!�O"�vϽ�z��ܟ����[��ޠ7Ѥn&!��0�R���P�C99��C������a���na;�&�V�x�Qb��<���##��՟2����~#���<;�m�c��]�M�U�Ik���A�c����kt��#]#c�;$Y>,k�g&��Em_9�$@�D4�F�C�����S�Y�i��Z�S$O�'6��n^_byj��C��X5H��;ƝZ/�� -}u7^�N������z¶AF�W���r&3UKG��w���c�=90-��Y��WMO��|o�Y
�[p'X?.*ƾ�lH��}��Ӧ�cΒ�*�]�_C�C�=z gu��e��%���� ^��?�k:�>��������/�L����4�	�%�s?��$M���*���d)��⦠ ����q��;�1��6�����*�j:YHl,n��V�\7u	dX;\�9oz�o����5�G�|ľ�r���ʤ�ӓ|6kZ��޼`��BM�u���%D(a䖱����4�OKkU¥���6O�4���cFH6��K8 y��bF�[K�&�G�b^\`�=����i�<,�QνSwA��*�i�@��D1�c�����	�s��ui�=Ǽ���n
� �=��!3��?nNs�p����K�c����Д�L�d35�t=�H��d�����D&'��RoR���d�>��yU*��N���2��P�'}9�oB_���Q�=鷽V��R�4Ж!�7�y�������~̕v��kq����S!��e
����y5츋 �QY��~6`ҟol^l���f� (�Ɓ~G��.I�Q�M52b��?������n����i����Кe.�>�������P04�l n��|g��I��]ih���fz�U~aK|Q�MQ��n��(��%}+țN�ؿ�|�a����PHaU����sg��A�7�.ygI�>U���������{��:�,*�G{�iH�S�����ë���D��hdz���
.(-"Ą
�!��N���(���{����3�|��*����&c�m扑i�z����PM��C=ȍf�X��BZ��i�|�"�X`�gA��XK�ͲZ��b�&L����K/)��u�V�6�*SR��Gi��f���y��������EL�V=�� ��]t?�.����[���A(�dɴ�b�z��5���/�r����'{��s<�#Q~�c��kJ�]�b�ք�דƅ��B��V?#�Z��h��/ze�\Y�����gQ���)@�&���M6P�����`�`}���-�L�,���N=^��K�+ۖ �KR�5���u�g4��d-���=`�����D;xv��zW� ��V�|�H��30g��'z�8�/���	�o����U�w������|��i���J��\��)6>)�Q��NS3#�5t�y��N�Q��*;C�>MT�d�<�{4qlnU}]�um��Vz����5�&]�L;
�fw*5V�j�~	���wτ�eL��Z`�[�ڧ";�.�i�� s��U�����!.�ZJL���_�Z��qh�C���23��QmXڵE�&�^y<RN���"������M�y ��k�8��+�Ux;�	A���L�zf�������T�������JBN���Y
WRz�1'fy2z�Z3M�O� 0��j����i!M��s�j�����Y�_��qVPʈլ��1J?�h��_*n���3p=r7n�u15^u�8�)[�g��np��Q�^��f��3�!���\cg�؞5��D��2dI���+�AϮ�0�����n\��'3X+���7�b����|�bj���+�⭣K0XMoϳV��"~����Vv��9�)�"�E=,�q�h�rT۾pr���<����[�6�/�$QL)�G��.�K��m<�`����^1��8�s�i/��A�9X�dN�=�(iyPI����R`Q�0r6�<�J����F9t��82�Lz�a��Q��=El-"�jIə���z���=>�2:�
�gsu��ˠ�c!d�����M�a�X)8Q��3���Ƽ #��u�T4E&S@}��-��a�gIӵ �(�M'.�� #��D�Go-zڢx�2�ȳϴ�w�cq��%�� (�>���6�wQ�>�����TD�Oc9<���]=*�:'9-N_�@��ח�9��[1��;��3��P��B�y;��hPɞX���O�C����l�]��-�8��9�Pw'Bh�e�FZ�`�y$I��]G�"�s:�1���p�����D,�d�t�fi�0b� ?�e�:�����l=S�<3bF����uoyUw�S�}/�}�|N�t�֬�|��k���Q*�o0��%�."�]N�~��\t�N��}�N��Č�T�'K�O�tr�`��v�s���7�ǡ<�u�W	�b�F�k��X��D��E_�ʝW���ȑ�{D�Jx\R�
Qk��A��ۅ��4Iq���(#Q6���a��^ɬ�����߹����HG�&[�v�M欮j�jop��bc❤3.,��r�S��	���`M��-�b
����3L��h�GyȻ�ݲw�0ۣ��DN�BR*�$��"E_�P�)���Ӑ���;� C�mX�ސ���'p���N����ݠh��ϫFda�3b$k���Q��M� �x��ID�V�r��*奃[�1���u=i�_�I�;�3#|�/PZ��E�*���H�rM���Z�@\3�Zn��3����;0j�Ւ����s8���j��X��f5=���T�Pªk�g}(=z����@h�C�o�5<N�H�Y�u~��[��p�8.��`t����6��z�ѯf��6LD�i�k�v�\ځ�ܻ�駑�69<�w,T�z�EuL�������>��gv7w��)�;�Z������D#KQ��ŉ&mLh��}ٰF��KБґ�?�iW�.h�3��i}��E|e �m��J��W�����)�0�̂G���56����@q����	�����J�Z�#�_](o�[T<B~
�(;z�Co�\���Jr;%�����Eg�Pp�ks�ҋI�(�U�W�11}&i
M���o��Q��0v����P-�L���g ��\��������PF�K#e��ܬI�"z��)z	�4JiY%ء8��� B���EK����Ԕ��]>+d�rU�C�<��¢��ڀG,
h����^��{;~z� �{�I�q�"s���)�%�� �Q	)���_=���]Z��	m����Ã����/+��=4~�V�����2�cOXkv>ސ����l�F�:��H���jY/u��T-kbz
��w��]OYr�T԰hyǧe�#l.E�+�Zݶ��|tK�j�d��I���ʗ���؋|�C����"���mQC�����3���,e)���m�e��H���ё�k����9Ej���!:D�;�[I�|�v\�ص��5*��� �ʲw�ѽ��[-� ��_h�t�IK�|��v�Q��W����7���!�(�[mT�2�7{�o��>��v{0��)e��![����IG�s�^YGCtL�(����/|��n��+��1"l�"bvG��x�O�ȩ�@�Ͱ��)��SZ�e��i���sﬁ�m����+8�{Ȫ�E)�;���Mڍ�5s�'|�"6���h�� �����,��vs�ߕ_'� ��OS�ޅ2@]��1�s՛�h�7 ���G���Z��1M&$Rl�P��t��{�Q�O�Z��["�|�7�������)e��Z@���w�25���ّ��t����Uv�!ώs?��8t*G�3ӊx�x$Ps붏VTzȾd ��+�us��?_>*�ŭ��N��W�wZ%�ATqp�#HԀ�G�G��
",zƺh>��FIx���f,�p4��R�1���'��B����C����პ��i��@���'�F2��'�e�v0N���"��65��є.�PX��}a'��%�T �Dpx[)F����{d���y�����*�|� 
�1c�� �Ҭ.�ӣ-c����O��I��$Ϗ:���e�z�֙wKy��a��lU�j��I��Xj�I`%��v�^F�>엺�k8A��.���f3:+z����d-�r��VL�� ?:O��V��I��`t�p=��_s�Y���㝸,2��U _��:��P�]a�A��yϔ��.ĕ��G�u��qPD�c5C'h�3kq��A)��I*	R�`�]���v�d�8S� �S2��潓�^P b�Hc  \�?o�S�Ҝ����p����xN+�<�v�w�$�C\Y���L�RF�1�Lj����	mZ{��.�K��Yo�*HG�o�4TIT���Q?�_�Z�p�C��RH��*�N��my�Zn%Z��޲��LHS��w�~�Hډ	qLѼ'(O��qݐ�,101I�n��^b6��(��d}��y�A�8���[��}#s��J�$򭖓|��y�����	�%�ż4����u�s{Rh��X��:��p>f�T��eXim�\'id�^�X�,R��M�`P��4-q��h�$�h���$�5�W\���m'>|,�K!8,W.@��e����žX�K��\R=��p0��x�gO�Z�U����Ot���ُ�a������e�`�7�' �E�x�Q��N�)h��c�huB�fh�?������%�V��K��u�B�5���I<���o�^�}�
j��~����A��x� =�K8�P��Y.�i������b��nR/&����w���d��Ĥ���/��%��̳�M����N\J� p�}��(���������C@N&=��iz�Lj���b��!	���D�t���$l���d ,�dAUXO0;Ӯ:9`(���T