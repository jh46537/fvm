��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����,��f9t���3>��Ձ�A�7M ��uj��M�0��{�ơ�Wa=Kg��!洭D�2�&�6����2�����X܋��x� ����G1���w�S��3�C�1�9��1+CH�<3�vwN��F�T�\#[�'I���ҒO*K��V�6�k%���D��Sn�&$Y�au��Q�/���OO .�XS}���9��k,[=0�hj��V���w��:g�!,;�(���1��+�\�dn�!��S��Q�j��:"[s��em8�'��v|h17���Kz.�0�!/
��3c��V��=y@��
9��O��ܔ4��U�ϒy/�1t���iy�N��/�L���\�q��oԭ�����jX-��ϸ8(��9��1��y<�c�N�"ǲ4�%0H|K�:���	�e��{U[�S����a~U�
BU��dk�	C��k�7Rʟ�F,�;�c��H�.)��@?���\B�Պ�'�;%�'p���	VL� �w�$jTpɑC!Z��3���r�I�D*w,��Q*.e�&����Ћ�o�%��e�Л^Ӛ�/�P��"ц&m*�8��~ł�s��U�ε]u�/e���>�"�$J5�q��c%��Y�nil��Q)����� ڸ$��3\6�k�(��66l]��W��n�B8���Uw����"(�	����9!P�
��w_[-������g!V9js��a��&6�z�"z�R��_��Ŀ��E����>v����wm�g��J����V��G��/��R;s�O#,"�M>�tOa���xm����=��K=�7���>���[/�}�yV�?Y��ן�Ohx6�4���/�y���%�O =���(nfJݘ9v=�����ہ6L�;�(73����G4�˼VȆ�b_�~�B'
�ۇ������o�Q��!��enu
�J��3�D�iM�s�����1� ,��s� $��3��y�ZdVK���	��e��<� /�2r��l/��<�P�!��!V��$�$j\���l�� �ޘ\���B�.�^����:f$���9�����jYq&����-o�*�h�::zPY-�߀
�QS湋Uk�V�}]�����ĺ�$�yU��k�����5J;�g��nѧ@��Ս/7kL���T �ey>��/s�5ퟞػT���#S�Uc)A�Rmc�e������d	��,�}���u	8Ju3�7;F�ڑ��'r��$-�˹iT�����>�h�m�����w#�&@�\�Q��<Ѥ�u�Ba�R���D�@��\��� ff?ܢ�K�s]�]��&&)�V(w������O����7� ��@��� O�8��ۂ�F�e;�퇕�0����j���r�9�|8^wA�-9��&T�X��]9�(��T�}�#`"�@#�}�^T'Nٙ�����
�U�^vA�~�ܢ$ǩ�9�)~��0�����^$��"��dm%�W��ژ�98x����R�l+�)�Y��%$`�(,aB���O���34�)��|��]4�@g�;k�~�Ǫc�o�' ��Ū��"e�oՠ�?�L6��E���[30Le+�P��ulR9C�ȱ��bI==%��xE�ET�31"
�wQI�TN<����Dp���;�a�o�Y&Xœ���B	�#���T�9��3=�AL���1u_��|���6ʞÎ}H~�E�w��EzO��`������"�z'�o� ��D��>��x�?|��/v�$/��� ���l��a1"� @��9�{���t@��ix��0�)��SB{����z�)��R||u|7��#� ż}�
b��=��I{ ȶ�.y*nq�P�%�?���k�K����r;��2���zBnuF|�թ��kG
ƨ|o��7�nn�S����nRa+�|a�Z�A�����0�}`;|`���3?�PzB`�1u5���׉���a=�Z
��=������=��|��el���(9�;ZGz1���� � �2�U��gQ
�-Cs2׀~�uܐ�l�@�����&/&��0.5,ad����N�����c����A߾LI3�-��D	��暝�ů��5�|PŜ yZ.l���x+�b�@�~�/ȭA��Ȗ����kp��n�.�����<���8�^@��ـ�?���74�C�t�	��U�0�LyN@`���I�g������FTVS
�@[���b0Y��uN����F٭�*u�f�H�%�s�|�<�Sw���jc��t��Q$"��J[�j�˺2��������C�\{�2��D��>T�D0�c��R�Ò��ת���2QAS����0r�K��- ����V��!a��?\�2D�闣R։��nQ-�y[�3����&P$��b�{�Ə��I[.�P̖fhpM�@���(�����"����-v�C�i�y%zNap'ʓ62@��"!��5Ă�1c�Ϊl�9m���(�� M�>�ϧ����y�[�cw�X�0u��Mm�j�1VO�y��Ԟr�r��Wb٤`����m�ԭH�A���4�O�ֽf�C�ۢ \�F��-�:j�9�5���e��f�Hr1�o���>��'��R&�u[�=�{q�~��ܻ�)t�&4����T^��ѣ���~ ��EJ�f%jw��N}��탹o�{���!�u����Y|r XL)t�4�5C���q��mt�P��3�w�
<�w��3T���=���6���)Z��#v0�zL+����_���)L���N���`罤`��,�^�sDU�C�+��@x�&��� �O�b�qT:�4�q��ƣ�d0[� ��Ϗ|/�?�䕿6��~N�����
�;�2��A&F�f�O/�_1�6�0�j���)�ޘ�I�,OZ`s�RE9Y�?���7_��o�a�e��j��5NS��k�8Qo�t�U��'��_�5r�%���I�GF]���8��e��U���[(NzjzQ`B�c��ifr����@`����81s�y���q*|߬s�N\`X�IA|��el^���!TK�9�[��x~���Q'��^�}���Px?�؟�f�-d�f�'�_L,/����B��W��P���D��nҤ��2[)��DFD7s
8*"�:�z@5���:ݔ>��w>�������\N���4o���B-�*�������t�x��@4C^x���HB����n%�-X��b�ٖzae���7�c&QsPb���(XҊ�n�/`�*�W<��yb�CJ~�qv�W44x�HH�x����MB�b�*コ��n-L�Y��<]-7��&J���7�:d(xPUT�d=&c�tqX�w�:ݏ�Ku^l�����/��.�֮�JG���Q���/�h��F����լ"�ŭ*w��E:������E��X_>�l�IԞ�U�9�WW�U�	����4�w�<���J�v��������s�@"��}�2a�T�����:���6S�q`������4��
@�@��A�%��f1d}�氡nWJ�Q0V�%Zf��]	{W���Qi�L����Q.���DE鸐Tar�I.˩).
7�Q ����H�~!$�)�� ~Ȉ�
��ऌ�Ԍ���uQ�<��+�����hG����LE `���&Wa�_#;80�y�E�R��@@@ʺ�[���'�09��UO'���n�����8g���"���K��=$[��Kc���i��h�}�@?4��Oѻ��g�z�voE�{�����IEK �E��q�p����%ڬ$g�_���,7ёq4o�U�I�ܒ�EX{��$��v��#ڱ�\��e�]�X�elT��u��cw]x<�-�F�l?�l���6Z���'S���a?�!����|�F��?uf��|��:���vB�A�'���>����Gn�� �E����u�B���t
Ǩ29^����9��1Vג��G��ŵ��"�_&�F�åt�Mf�e�`�KL&��0�H'H0���5�Y:s?X�AP�������R'��1��B�ڤ[|�ƥ��F?�ob�"���;37�4����oN&�%��I�N�����(Nt���Ȝ��F3�L�����¿o�tTc�y���ڶU�"0��i٪�@y�����X.�Ԡ��X��pk���ۗEFP���X��5R������^*�"2���&�Q�@J���1�}��6IN�E�%U�f��s�����E7I����yH4������@�g87�5��TĽ7$�-e���vi�]�G����ŏa������dM��
�2��7����)B�;U��M-�˹B��N��ӿ�gx�8XHD9��ECO�+��Vz�/R��R��J��[�s�j��f�#����Zƴ��b�1h�Θ���#/�E'$��@���N��O���0��Gg.��t��e�\�'�#��=3���	��"��=|l�B���~�:�g�2�HZpbZ<��1�g&$�V(P��g.�B�H��B��l-�
NQ������L*/��A���I��T�m܎Y��?��<׏����o6���?�R�J���qf����{���#��I�;,'�@bWN���X���,2�̀[)��[�*�i��׵���m��=�\��%���sFnf��e=��ad"�������0jD{ɨ���o�e"�����#fS6�߰1ƛ�v(��-�
�����C;(�(z�E+MaB�I��H����)f��_��܉�3ji�OA�����/|$��@�>����YBl\)9�M��q�
� �,;{@Nj~���Vb��UDO�(�\�o���X���j+���eB��N���)�M�,��c���T`%�j��E��[ݬ���\qFn-�'��7�;��g�Y[I�gB�~I�M�>hO ��$��]��(�󾠳3K�t0f|���[�T��l��}��Iް�A��%�(�?��8s��Sy`pF�e�s�*��;_s�=��$��˕KYmp�p�F���Z���_�3M6--x�n��7��G
<�}���Cc=Pu��֨� �f,����dm5�o@!�&���J^�<_��N&���)�M� "z�[�v��E h���_�1^���[��Cm#��2���Ԝ�
�1FB&/�XZT�КH�Q�+^�>�0Ϲ�6�EXѿccx��L��q����8�O�����XE��Y���èꭂ��(�t7��\�E�o-��>|���K�''�\j�?N2�
����I��������B�e�-��}����ܝR&��.e6���Q�W�3�L�sJ��''�9BO�q�AI0d}Ә�N\��*�^D�����;�>%��&yć�ݽm+��*C��9�
��﬎�n���T����^�j�L3r��X̪ ����<��J2�CȐ����u��Lz,X]3+x���%��BD����2�|WC��[d���#s�bq	\F��68;%3,tQ�|�����oT��E�Gm�����n/�;���/﷈F�snX���k_ vЕw�1^�Lo?AL��B@QL�4^��ӆ�r*�!b�|��Z\ƒ.����ܪUr$����C(i��%��		�m�c	�޳W���z��Ӵg�ڬ�n��m��V��f�01 �'1�G5����6�$���ROJ^�K�?ruJ����z�� *�t����fcV�$Jh�,�t��3#	A� �u3n]�(��D���KFY��[�o�S"����ZІ�g�#����!=|'/���\�~j[փ'��ƦY�`��Z��Re�H�r�����3L�̇��iS}�se4�I�&�8�HE�?/����b�U0��g�:|Ƴ��x8�wv~�����	��O��л�6�� ��Ǖi��6>i���sт$���Pa`G���`=�@(f��Lv�lH�u���L���ߛ��Pu��hZ'���";�R2>���Ƽ��8������v��br+���/�$m�(�����Z�w�U-�OL`��1�\ذ��=ʦ �����ş�1X��L�������w����{i��%tj����Z=XM7z��ONL�s����ґAƻ'��)�T|s܎_���ũ9ʗ�����b�F��t�����	:���K��	���$���ݢ���h��i�Ay�����)+~����,��E��l��
o��!K�w�(]c���wjP����kDBP�MǙ`�%N�--��M?P��4W��SB}Es5�Y?��mĚcE�u{���@|%g�9�_I�?E�߽�b7�rg�5�v���Ja��;�y膹�R���������Z�J�h�Z�8V�5�l1+�I����Lf���׭bm���
�)+�/ˠ��?���ދZ��4>��$��}�iq���ǐ��D��O��	$���v�=�FT(8�'-��(�B^�o�I���fZ�!�{�D���'����ZS�����X]����8���+&X]��J�@}�:d.jB����M�p�*<(�����Y�I/�
+���N���k���:��J0�KCOU�~3�R(�v�����@�hӎ�4��u�2�����%G����MQ4J&m��X�.uqqD-�6cY����r�ա�M|Q-N�F�az9<G��Z���wS�U�տ+��olN�Aw��Kz8U.�DxkC8�ú��J�)G!0���Fp��n�(E9�S'��7�*����p�SH�'�� �[�:[�1�?�]�f�D��1�L�Y�Df%nw���[��H��1!�e�p$��V���y����l��9���婌������`�A�v��+���2s�Cj��/�>�n6�*(2*J�3���<@{9M���������vͽ���|�����'�`e�dZ�mR�<�����nS�O� LAH���bu�䔳L�5��X�1O��*�y��Et���:T}��U�rjh�7۞`�[���̲�E:k�k�[Y�|��W�mHV���@�Us�Y���|,ܣY͕����nk�ȓ4���K��
���>�&�t����R��S��'ߡB2�D;0e��m<��3lC3V�U�j;�Ʊ���P��ɥ�s�D�զΥ��`��~���)�އΏ�Q��
ؗ��2N����ϟ�߂��$	1[0�4�ޘ�o�6&����,b@�!xU�+x6���?$��|�!��u�V=؈PA��^�������o:����n����3u"��'�In�?�Z��wVU�cF��蠗���]�=I,���#��u"k39I y�M�t�m��R$�bcvk˒�sK�htISE=�T&�o�~&z�l�i�Mo�J����a��N�)���a��Y뷟�RdG��L���L{�����R3�h������i�e7e:�S�:5���]�B���b��k����b�R�?p)�Qpu~Ɖ��n���1����Y�4"�K۬S��ـl��3"%Б*ȻpOfJ��B͌�N0��GiO�������;׵8����Qo�0��a��/
E�d����IΫaX�_ut���x��@�[�%/^⫁����[�L��Y�&j�4�6�t�����*f������[��໩"���P�|���7��Չ�7H��I���aJ|� ���.�|���O�ՙU0�*�ɿ�H�^�S�Ԁ2���ڳ�049m�	wࢁ�����-��%=q��h��B��"O��������?��D�5�:�U��cN���N��
�:�x�&������.UnUB:�ĻO�l������rO���~3X8�~1�aa�&[�_	�6�b��l��+ݠJjP,��}O�\hN��l�ecj�'Ï[H�]�wH�
�q�6 W�T�YT;"	i��s�V�$\4�|����+���f���#W-p#J�P��Qۼ��%[��3(1��\�/��M�ʑ)�~�G7���ސM�'���3���*�"摞�J�W�]�L�^��FW��c��GY��'�y5B�R��Y������j��蠻�E������>��.�{q����m\otŜq~����U<]�!�2�vf����oӑ�6+`6��X�%�n�|Ỳ��F�����2mC�n��@r��L?L��/���30Ym�L���;�y�� !a����a�a;/%���KЧ^��}����޳C���^vD�2�}�)��1�����ճ��'Z��!�ĘgbYW�ώ��L3�էj8�Ѡ���'I���MM��h��[��n G�oF�7��n���R�)��J�����f��[������ryZ�������s�޴M���5�Ou`�U�La������2�O��6�C�f�ؕe,}��U���K3-�?�$riqE3��%[�<����r�7)��N�}�A�Eڀ�w�[�������ZPoV�@�0��	�_j��FG������鍅���t�ٱ� <r�W�n�:ar�<�����{�X� �	�_��)/�0�L��Ke`���d���|�r�"�_e�!�\�jX�T���le�׌r@�S��w^�WND�&�kR)�m9"����2��?�0�71E�J�c��{_��׎�i�ɠ�����%�C� v���8d�!V��g��1��b���T����ƨ�R���7�U���A�2��'�錴��д3�������d���i�[�}�x{�]�BA�a ǟ#��Ɓ劃
���fD��L {@Ҏ���Td�$�ޯ���I�����>����F0w�Z�џ��g�ZS�����*��/+È�j��x>�'��FPpn�س���( �$������G��4i���j޻Zd�SO��RĬn/T^Cm���~~�'}n�9�pAن���Zw��[��R��5��"��F�FG��/�vд��N�'q�p�R�;ݬz���ޠ�\�
/�~�[�Q\�ͥ�$��^���܌~�oҝw'更4J�˻3��~��Yxd��������[Lw&�àV09�g\��U!�� ��iV��F&��.���!:v.)���Eʋ��>�>��Mj�l�%UM����U��,��@g*3;�}��sBv5���v�@���V	]H�GxP�Ԕ��V*�^�]�{!�-�����=`���knBhi`Ϝ H��t�3b�z`�\�̂OH�W�ǟqM�y�xxP9�_]��)�;;��@�]{4%��K�_�����jE��2��	�z�ZA�/�]y��u_�~R,��#+ȝl��%y��U g�X�b�*A��w�eV˓�Lr���U#9�(g����?d ^�g/̶�hpyX���O<����
Y�Ln��&Z�k6�70G�Ŕ���@v���SXېgY��ө��
��\������){����C	OVW8�N'phԲ�-���>�q��
"hȹ{7���Zd>v1�\��N�˯j߯0[<D�4L*R1��z��3�����	Tw��Y���U�z*�,[�U����9	�\Һ&;�7�@�'�(���}e1x-��P���̭���ʧ�����Fs�rE o����������k�M�V������q!]��Oʁ�䏱��1��/�)ٓ",���c
��ᨒ&�u�+����sP�Ĭ���m�n�� $H���� �]�*̋&ʒ�~����C�U���]�k�^�P;��h��qG��)9����~�+�t*�� g��n�����������;r����omkeP�W"m����[F���I�5�Vj��𪨡�� ���î�U/�U"���Z�oLe���5��'�aپ�lk[��5!T�UF5Qj�.�Z�<���'U�ɂKV��-��vW���.��b�d}^������^���_=���T!�@o��|��4b�V����k��k�7N�CU#"���L.`������i�J�$E~�,��5&�_i0��h�����#u������ �	'X��cr�V$���\ /�0f���쭝4[ ���J��ۓHC������5^CI���CR�j�͠~���Ty~��MRk-�ʼJ�8"}���B�a�[�a��x��"�ۡH�Л=<�J�S��ˎg>N���ګ��.�_����1A��f��l�us�\	�o��ngb�!.ɩ�Mk�l�7q�cp�z��k�gII��m�h�V[���9gM��.�)!X��ѓE����a��� }�b4ɓ9��ǐvِ�.��W~� ����IK5�wY"����,Њ�\�>y���S
�J��V��H��ljt�e z6؛p��3� �(H6�k��j�03UP����2)�:}�#�[SؗTϛhe�J۔e؊����_� D��2�&1�n�P5�B~��2QݞYj(�x��ژ�M$m`�r��z.4��皅�ZE��_�B)$�Z:�lt�%j��䑢� P���>��N�Dte���Yռ-�w�%��v˾/F���̕�Its�˂#V���z#�����V$����gM�w��EOi)�/i�v@ǿ�wǗ��������
��*��-������;ji=u|%�"����%���l)��@� ��y�e� F\�����=NXg�
V��)"��HH+ԩփ�r[&��h*_�Ū��/�eDa�p�GQ��3��z|*>�4�$�&O׷�zũ�s{���Q7pn�X}u�1>��:���7Y��9ɩ�i8p �І�"G�l��/d@Űz2��`�8��¯'p|ߎ���e� �����X�\U>p� �C�(w5�Hq�i���jb좃[<�B��k���7�sP�0�[�~M��F�t���y���\d�P�g���D���BK�jI(]�>�.���)�=j/���tu�E�Ch+F,Je��ku���c�T� w���2&d��,�5�<�^��\;��O���������W?���5���>���:B�&����P�k>�T-�c��,���>�O�:7Z���/�Sl��6b�/����mU��p�w�  -P;|���X���<J��1
zra%	`�)�K��nT�������n�����:)���m^�y��P�*!㲕�rZ�d�����i���6�Q�Ah>��YY)�W���0���j���OW2��vvS	xx�c�E���MH 4�>����X.�$����KK[}Dq�R�D�����lk�q��{;[����]��-h��0�C�X�R&s�r��=�p;����gV��[y�ʪ�we��΍�i$�>u��eLX?���a栶p�8iV4x��>ק��G8=�Ĳ ��������n�,�/3����k��gI��Lӗ��3�6����Kc��U��E��_j(E��A�Lմ� �n����@�e>�9�*���}w��n����,���O�5�Ԩ�?�7���CԲ$�f�����48����]j��W8'1^�-�Ʈ+Y�>��{p�G�56�hp�$nm8��T|}5�m�����'�����_P/�3g���w�9d^����.�aS�2� ���g��+sb/�.�XÁ�u���`+�fp�7Lceگ�T��	���	�l{Qu�F�',f����a�����<�E� 1pLh�p���(�'D�)����ݵ�L�U	'�ؐ^�w�Lב��k �ǹw�O\`�����g�����o�0��,�c5%��?M��]g�^СV�����q^�y��7�x���x>&$��n�kV�Dȴ��צ�u����f<�
y�6��s]�j����-̾�=��M�ݳd�|�&t���H�x�q#l�����NY�D6�[��:(W�"��gY�~>��o��娮��9c��E�C��X�m��|�P��h\���Ȍ���%]Z?7�F�bz()%�� �G��jTs�����(�e�W=!ό�\Z�0A�[Y6��ReηR�#�4�Ng�7�P�7��H�f7�T냰Q�f��a�a���������q�Sh�}�H<m������h�71(�K3���k����9�w�K�[���b{��?w)����j�}��7�, C�^6p!�IJ�M�x�{�r.���p�SV�%x�D�X\�������i�j�����	y=H^�!���b���'�xǹ/7U]mX��=Щ�?���hD)����_��'-悃�w1U�
I`�$������jQh4����'4k�a��]�Y|a�y�+�6L)q�M)H�<�jC���$���ն��}�sN�O�S몝t�9�Gh�&�C�@�̝jaI�X9<�}I�l��ꇎ�7�;��y�f����0������J��GAH!ܮ/��eЌ��H��TH_��7-�f!���W���r�(�Y��ev���,ͧ���+�[!�	�$�󥃝�n2���63��\��m���10�7��[Ӓ�,����(f0�/��
�h���}T�{H��S5�-y~�PD���{c8D��V�w��S@�廍�]w��6j��h7G�/��
3�Zk���j�6.�Ξ��ͧL(%�e/1g�#��3�o~MH�{�l|ft��
�;-1ƽ�aE�7ںVh	�@�lh����ʖ�Z�l�#ڶc%�����\�߼1M|~Ѵ|!hL.n�	�:�?rq2]��g�$������I7� ���ɓd�EsM��c�,�˼3U����[����Y˥�e,#|P^|��N�M�F|�׈q��9���o�� �����Se
o�ؤ%���E��m����]-��"TM��[������4
m�u�A�j�3����3�\[����x�C�&2S8�h��m����ި�5P�����-X�����B�on4��b�E(V��Ϛ�%ޙ.��Y�����A�h�����gOt�<I��_nz���x�A�^=��H<�یZ쯂��w�L$�z��hyB�fBO�������ʴ�*ߝ��[!m�J$�*_9��=��1`�y�(o1�s.J��H��o���'%�}B��0|�Gw����8�6e�%�$�����ײQ9��Q�q!�P\t+sUg���E4\��S�h]'���+`���[����B�.)  QR7 ���fC�&Y��5��X�F�tL���"�_V�Φ(Zy�OJ���})ud`z��l�y0�	EpT1��J�7��� ���D2��B��N�`�ٮ%^7 �m�AG͗}W���jJ���V��̘W�I��O��O���	TiQu_;�x�����)��T��A��E'���Z�B)o�r��_C�W+��`��Dx�����u^<�����<�v�M��S����p�w��ܹE�ҋ�)�R�=�������O��qdv,�!4Pٽۘ)�S�#�M>����� �M�&�t9E3���y��u�&F3��E�}���h�?�=<�a"�wL�&1Iݪ�(/�C�����4�/
�6����;���^�N�PU�%E7�Z���S�V}�&d�����3�������&��i��M���t�ȵ�T�X&W)|�A\��gq�6l��˷�"����}�-�Hj߮�.�B��"����1̌-s�S�#��!a	R�zh���H���׶ O�Ff�s{c�\Khph5��F1�w!u�E�`k��.�c�奦j�MA���xz������&��Ȇ?��b�3�7R".��1�� \��|fɛe��zH�%e&JV�x������������;�~�Ѕ]g����F
�pS�����/���x[�ݶ�W�����y�����1��Z)hR�b�3��Ԣ撝hE�m�=������Յ
ma"3?���=չ�G�}�1r��L3i��ٱS���H��&3	Dɂ=%�!��>dK󞑫R������9CT�iOB� �P*T���zn���{��>6�J��#h���}{������-ځO�9���p�ط(�-�<�\%W���}��ŧ�t�5P����[�ㅋ4=ٵ ��;2�B<���W���#[�b��R�p�����}4��i��o0�<j�$W��Ľ�券�6�l���u+>X�}̙�4 F2d�9�� �5qf�iU��..��
��@!�pG�pC���֟���ݰR�K��A��~��R����;�����
�'L�r��,����BG��.Y�
�|PE:��.@tC�R�+�<)0f�'��"��0���D!4��j�Hv^� W�ܵ�-#�]P�j���Dn������|A����`���줍0�����`ʠ0@�֎c��\Qqt��9%!�^��J쑄`�A �K�x�,��rE�~�)�ߠ�<�����1¨�H�V��f�p]P�� w>�q����؇�2��* ���,��9��x��٘i�^�f�������۾y���:{�c|R��8 d�@�W�|��.�%���]DL��
�"^���a���w�;Q&>�}o�*�[!n�N~�a��n���|\�Ѻ����y?ӋO��/U�[��� !��@��"/?%E�9��m�m޴���P��/�Wˢ�T�l�Q=JٹДE
b��J!�� Udi�X�6,fI졊�^�oz(�$��.K�ΞǱ{�3[�;�
PM�Ȑ$>~k��Gl-M�w	��j�����4hXy�K�[���K��3)�z�S�J�?�R��/r[�K��(�kxk[8�ḡGLVO��Q�Z 	2���e���N���eb������&|�����M��'�c��?N̺�A�����K��Ty�[
/�3���C �|3Nj<h��M�~�+���/5f �ޏ��8���ٗÜ6f��9�����7�O�0�ch�!7��W`��V�&�}[���ڑ2�<�pcЬ^g���AZƕ����yݦ��	��s��l
S�%�,��G�v ���C�R�50�=d�x����J�D&��L?A]�lATil��{��6��J����ϸ�	����\��oB~=����enMV�a+�n�t͓Vⁱ�sMN���a{�!��}�,�kK��a�mғj�ܬg�Q���I��N�f��5<���A�Q�B�x���Kkek�����Q��0�۵}�T ��ћN"4vee�� ޾C��O�.��T�U��#"a�0��a��z�h�c��66K@Ɖ�Lw�@�\�D☷O¾���R2�o��>+&u,�W["�'w�70u�jQ��>�-�ֵ^u�@J6��%Päf���KUzp���'�]�\qe�F�T�a�v~��YT��e��`��"�3�����m���3f2R ��j~,�{Q��N�?8�l$+�Ip6?���P=ߟ$9�W�#��</=�.�!�h�*����u��	���oJ�����x����L�NnO��|�|wݤ�T����f�r���f<ucIa�£5�������m�Dc��CE��[�(]Ʈ�5�`.��T�g�/�R���t}L�����Φ"jѕ�:���z���J{��bA%ylЮ�)�"4�W~\��DuI��cXc�RQ�2*o�S)�Ҧ�,��O��1U�H���`�	�I�+��Z>�ת�[��h��[��c�G1��؁,[����"����ƍ�,9���g��GQ�[J�9�քzC��+[�a�V���tӮS���}ʾ��1$o��ɖ,6��ezy���	R��V&}�
_�����7mo?9�*Y��pz��5����trw����d�}(e��a]�g���`��+Q�F�����;�,bB�/��/�cQ}G�IYX��h3;c::/���t�^��Z>ODyo{��H$���.�N���1���Lم�&�@��п�"+��K�+������A�{�H��DԀ������K_{h��|���Ka]'vE�@k9V�	x��b�Vm ���Խ��bP�[_z��g��>�[i���� _y'n��e�莺m���[/��C
���N>�i�dg4�ծ͊`��u�U޺L����3��d�$(����Xė[Ѧ��^/J��u{�g.�
�S�a�q����i����B�����W���������!l���z�]�-6˹���2mó����&��իps�+����2';����Z�i|��}	v/c�l�N	�k:����.2R�O�e�w���L��ݎ'%�>]b���(yLχ�	�ִ3��T1b
t�I�Y߬����W�z�v�����w[��ffm�捆�c�aH!2z�KI��X�jO�C�6�T�_�Y]2�}	y*}��������H�����iH�V��6����O _،C�Z:���	���Y]䆁������
	Hn{z�i0�F+�,f %�yvaт�vA�N~y��a�������TvQ7�n{]�������jǟ���+�% D�ci�Mh�ec��Z=��	����E�#��� Yr�P��������G��@�֔r��z�n� "� [u�9�<D�#�x�(���G��u�m|vb�ޥ��7�h6���:OC�����P���
x�߭^R��,8yQ�w�N4���sc��\T2��/���j�Kz�cu�Y@ֲ��qK��s������˰��ٓǾ�K�@�Jߝ����.�J-U��~Մ+�;q�A�Y⃛а�?9�55�a��9�O+AE�\�b��-�C�
ն�5����F���KW�6ϵ-%�/�CٝZ@��Lf����ϙ���]��}�0��Uy��9+�eK|*�Y�c`�8C&��sEM ^CZ~`����k+�O!�>Ո;�85m�h0F��'���*7#x�&�^�f��}�U�}u�/+~Eͭf��K��|��� ��gV�����)�}"d�5��-�?]����8�����R{��.0#��a��z$q�G�%���i�銱L�$�����xã���r��i��	�X *#��2p��(I���ܫ2+-�C�:a�r�!7t)y�E����B*�p22�	����'6[��-�M�~���KO31�i܈C����D�
~�:�"�n�&vB�|����J_����Y���9����"7;��dR��}7�2�R!|����Q��>��a��YF��N��Ţ�4�#O9oX":8L�\�ʱM�$;JJp.4 �����2e$�y�
��&�m���_��Yvr�Z�)G�K��rT� �,�wQl(w�gj��A3��@�m�\��#��M,A�|�zcNMN��w���u��o7ŗ-O&��Wܖ�
�!�nH~��>�X���Ⱦ�H��"���\����MG��3䨗��w��Q�*w0]�B�!��j��mͶ������oDd(+�Odq��}ĸ`J��CM/Y[����Pi��W6�d�5D��W01�+F�9<��=6؁\�^�l�̝��ym� ���"pA��\p����q@���`�#ȃE�l�~m8��+�i���h	Sn��edF�������H�/�G�S�v�̓C>�fN+���'<,A;�p�dk`EeR�'��g��J`�;J4Ų_=?%�Z����d6]���k�@<�c��)�ށ�{؎6�0�c�CJ����͓��O�%�J��~M��V<�`��Jb.:����Cz��Z���*ָ�}t@��Y�~���#�מ	�@'C��Օ��1�e)��u�Yfs��҈����T�&4�
.��R��VwA����8�-�sbc��;��ppt_��������U��@�m�n�Q��lگ�DLd���^���3����E�����nu�~~��j'D������)˧�1�@�ņ�o6&q�ほ(��"��ͧ�'57n���%�y�$}�[�A4C��/�}�@6�dMX_M��.�_���rP���׶;�Tw�aT"
��D{���/,�Q�<�y���ؤ4!��8��Ҫ
�ȘX�j�.��K�a]��l��{M��/�U���U��M���g���N��k��qe=����P��O<�w�ߤS6���{��x���MI��=��Q�5�𽰋mM�y�ڞ��$��6�)9,��{15��z����Se�C����p+Ph�HZNq�g����WihI?��f��l8*@?�=¶�AĝS��u�����W��g~@��)��=��iE�@G��/w�>�48)V�#e�sDnV���7���F��eVL�P�[�hR��<)��3�(�{@����c�Zd�J遉�$�zd_�{c������0�P���5C=-�dD���kD�ŲZ|��`�_wOE�u6��a�g�j�]:~���j���L��h�f*:b�.=	SX�K�k߳����H'����Z�8j�Y��Np�A�X��˲x����Ƴ��F���E���H���1<t?w
�-fh�6��i?�~x�*bj�Iӽ�o(�ϖ��5���Ҳ"C�{ZeW^WMS�0I�W�~��[դD���GE@������E븲6&*2~��PyX��D�`=�N��UT4P`F���O͡Z�}^֪I�����s5�N�����.�����Z�I[ܮ���qPࢁ��kw]��_�j'0��~�T:JF����lq�qR�뿑C�7��J]�P��Or�|8�V?~ ��S����=��Pҟ�����t/�NE�������O�I���}�d&��togs�0|\{r�=*�U{O�k5�=9��C�6׷�ir�$�'�:�����-���{?��b~Í����R�%P@֕�m3@檢$[���Oͱ)���d,����RlP��(���O��}�Ru�כ������G�P�r�Φ�f��XT�;ibb��:�����M?/Q拉w�ɪ�w �ED��?���A=ES�_=F]4-˭8,�}U�|9����a~�﮾K�ӯm_e��7WȀ�WP�Sn�@섚��!{hsX��E��8ӯT/�հ�R?�[	Vd�ʝ�pV���X�(��	Eq�g�i���a��jk��*�N�4��@)�~�����R��S��S��Z��y����Xc¿n�*�����-�׏,�f�ㆵ�O�cG���~NGp�}2�vCl���??%JįY.���m�2���4 ��P�xف6n���k���Bh�y�7�UR�����!B���"t�Ղw��+�g�W��Y�٬\C�a޶+#L:H�'LJ�A��eKWλ��oaT4�7}�z(��U��x��u��d%�F�e~I^z0�9�4�<�(�������p誩�����.�׷�����KsNF�92�4�4o&�A�,�B��^$T�*Qqo/J���9���5hȟ�� 8A���Q�*����d�E�_5��Gm��Q	dS�Y��������Ob�1��������#n�����7�����"-�e�l��vf`篗�wt|�?��!���4$\�+o�ma�-K� ���2/�Π���c��L�u���/��%�J����fi�egړ�����3mO1�w�����Bry*>N��X��(v�*/O���L�3��w᲏�5J!���Ap�ux}4Jn�{�N�7�Vd���9ﻇ|��&���
�+�A�	O�煠��PG=p�:�<_�v����>�����ɫW�*A讼��׭@xzX}����e>�2:��uM��; �h�o�I�B�?�!:wL��,F���L%�T�0�K��bY�Dc�Yl,�U�Ђ�äP??-ȐɃ&���E��O`�v��Έ��i\8y�=��]K'*G��I&����jz�"�lvv-G��_բ���b��������6��h/D6�tB6U(��W9Y��[LP�>�0AT@���}��L�n�u��96�]���آɓ��]P�ie�87'99�{�Go������H�D��7����?�۹����j�qP������D�fGqh�C����+l��9�=����e$��_C� �G�Y�:C�4�=-������������z�C�7��9[�zz�F�<4ׄf�Q[7lk�k���A��(��&	��
<G�����7n��E�bi@����SXN�S�� Ҋ/,�zT�wW�@dP�L�ٽ���HمO}}Dk�W7Y���Z��8f�8���v[ET�'���fM*JQ����:��Ĝ04���
{����B�)�%�b��F	�<�0ڰ�����$t]��OA�����-9E��S�ϊ�nP%�mj9���D`���[U�Oj&�y|gh?��v�Ą۹`)��!f���h.B���D �cD��q�hM�T��(m�\y2�w
�f7aF�BO��ͅ�˶�h{䌭�0.4C_4Պ�����'˘���w�CsH�r~B|����~�8r&]��/���v��N�KٿNK�����(�͸��q��aX~?��;����Ŕ]>� "i�16b>�ۏ-5x?�y���lVI�a<��ۊ�iE7;i�����>8��^U~W��pEF-CڈHڷh��!��Y�l�D�Zp�Vq�#�����o̙K�����uۮn����θ��Ä~�g\��K1,��� A������;�*��d~�:\���Ɖ�I}
mNf����?`��#�#��o��U�v����gy�|�ѧ=y9��Cn�w�J~�� g��1�R�����2 �;�Z���k��N�>�9�	8S�b�sy\�х�vV�d�ڙ3��b��ݣ����T5���,�z��F�I��� g�	�ʜ?3���I,�{އ�=@A���H՚���hd �LL��8�{��x�0R������Z�嗙�O���Q���[1���#A��IYyh���{����Sc�._5������/.M�� �ĸdȎ{�^ڗߟs��x�_��
(앧C@�rN&�3�x�{_ ��{��]����u��&7D��V "� ���lCN�M��?6�������R�櫒@�y��:WFE"� }b�F���^�^���%rDb��1!�ۈ=�kC���zV}���� �SZ��2��,6h�"�u���@m��)2(.�owk���n4�!�8H]ђ\���{�����>IS��Ȑ��Tn�3�&�Oy�5��8�����jj\�{�1���=6a����U�e�,�t�^�~s��S����@
�!����O�^t�5�9[���p[��b\��i����]��.z��H�}��4���M\�o���P
���T��.]�:�Zܦڑ�:�^��#��_�{q����B���Z��lIZE����:�1�k��.��>�>k��S��1�qeN�i�S����;=R<2�sp`[r�Ga��ْ���2�j�÷V�6~�)Q���/ǜ�zi���6�Ԝ�_끇����"�b=��b{�ڑ����O^�[���n����2C��=+?h��L.&����<i��݋��Gh�a�j w��aЍS�#�$΂s�����{�H�l�,��s&L鸨�Zk�]�����8��xY@�s�?�����L��I`1�8Zpkh�f�W�m�9}{s5�M\��!���p�Q/V���/KEf5�޲�b�&%�g��t�����)5�t��·���'�𘇗j5������ ��F̤�"\�#�C��'��C���L���D��Ҫ���h��
� �	�ܑQ�p��YzQئ��d:�q�Fb�?xA��ܖǘ���_�6�-��޷SC>�����5N�mx���tJ��E	��>��s�tl	�]�p��(�B��9�o�x����t�7��	�i�'Ǝ�O���\��|�I��F����Ad�.�?�5`T���IW� Z>Wf,���^�����[�v�iTI�B��/�#3'>�z^�~w'��U%,)D0�C��$CSĿş��a��V6`�2,����dXO5H���d��2��(�u�e�r��qZ�+�FT�y7�;1�Y���#4�&�"?�k��l(+v��zE�;��-��=�q�х�w� ���:e7\�5a�T,-�h�$~�훳�Ѝ�=���|�*�ĝ?d�uV�غ�6F��]��	��i苬��[�;���m3���ͨbiO�U�j�@׆L�����=��}�i���Ym��	�����IYbp_�����.8eԄv�$˂ە�\�No.�s�bp��x�)��cem�(lVAF�m��}N��H��Mf�q��f���#�Gx��[�?^����Nxwf�W�#�����}�䔠�w.;gJ]*�@b��DZ�$9�7k�D�o�f┞l��t����� �3�Y�$�1��D}����o/eޝǺ�	�_}t""��	:��1�����]�N�c��~SOjMڄ�zdӁ��i�fy8�~3�*w,��/P������St?�{"TH�-�u��w���T8-���N�(�DA��h�Ob�+��[E%��AZ��C���;~�uZ>�=dx�غt�hܽ�J�;a��7E� B��X_�C�>'gY����o�l����~�`+��<��2ƳlK�*�<���Υ>YpƄ;�R�ثj��'B��*�C�d�/B;����ݞͣ;���c�B�X$��$CB�MP�����0�/�2��b��S�z�-���SJ�O��L��u��Zs�νM�
c�,{�"��b��q�S���RJ5��9�wE_��� �@u٠y�ݿ��<����}��4cuz[��ȪGW�S���۽ �c�<�X�q�]h�{j���硞'oh|;�ù�0D��I'rs؟��xH����V����i�����Եܒ=��S�-���z:|�,T]�T�����+u:9��,�BAP�0�[��b	�{<�B���K�*���e���'�e��E����u�&���w,V`�}I�+������+�T6f�ѣJ�?d~E	h-L]�-�E ��*��m
d��V��Gbabm�4�+hF��fR�׌<!Ecu�wWSF?I�9��ʱ�iU�%���%ؚ�,���r����`����Y�vYyʷ��5�G�������߭vX+=�W��<(G,�P�.���*5u��(���/,�5[���D��\�%4�,������^�竝���Q�Uux��>�1�z\���Y�C�t���?f0��3}�X�Q��?�nO�gIa�5����$�Q�5c�e=��R�.��ܩ�I�N]���U_�@���RST�*<����l	x�����ǻ�f�t2�� Y�Kl2)ܓY����چ8У����?�S\I֤5�e���0�:y&��dF։H���2��	�r�@F�a�$W��>1Њ;�7��k����Ȃ <�ا�Q+�_2ݍ$��o���3�8.f����.��$nnzAFrw�}����ʕ9��`u��U��-�8�}��d����WuqR'9*��6Ȃ;o��$n[UQ%�29��AXL\ ��[��U1�d�Ha���~��H�6]���fD�z�A	�����k�l11F�@?LV�+w�V�K�^��ց��{IN�U4�&z�'N&�=��
�5l�̲hz^:���fuq���oҾў�\D��w+�����{2�%�:&�?Xw�	ԹN<X~�L�#��nb�<���vݎ�����,���k(�N��~W�:	6k�<ѯ�7���V!�� �_uH�%�<YR?��>H(�n~��O=��j�O�y����s9+ ����B��i�)ů����+fG�Xj��ǹ��B�n�o[y?�M}R}�⯗�7�%�?Z����^�-L0��>��Epy�G�\�?�]'�Y,3�щ������l�ŏ����\=�s��F]��U��*�"���.�a���]��ޜ�ޖ�������)�����;A(���Ļ�`ە�<]o�1jg�yb��
��l��:-`�I��@",��*<umG��b$�籭��n0.��Y�QA^����;Ne2­�T�j'�sؘiܜ@_ w�[[�k>���ȃLb�6��r,���U����bvp�8+Ni#G�ѻ�А�YL�`kFf���n�� ��ִ��������~�B���������GA�F�P�;�o�|�+��
��=���m]nxq(QL(©����80���!�����|�=�J�z�WZ�7	
6�!j�$b_5f�0��#��q����;��	@)��&k�;A(e}�\9�ٴp��=�HZ�"�D���Rzx`�ns ���:��="}��������48��(���"��������=-k�m����$�i$'X�)����!� j���P���(�����FrQ��ʔ6����H�E��S�Q��!��$?�{������R+�;�TkU�F�M ����nvR�*1�A�����r�I�w����L�)���_�c�_QK�F�S�o:��%���7jA���2�L�*��9���A&�H�"G��Y����W"�0���{a��Zl9�ҦY��5k~ĭk8*�� ���';u�sTd���� K��c��x�����N��oUv\�Db�s�Dz�}�cE�)#aAb{�]��v��B�D�WM�X�+�Ls>ߴn��v��ǧ�R�>���iH&�e�a;b;D�M��Ql���j�JG8�ЛՄζ����a��㯼p<ꊼ�(ق{�WhW\��'��3��3��bnۉ��f�:�8�:Ç���J��n�b���),�h��Sx�sAd�~N�""�7dQ�̥2�>�n�g�2�"Y�`�.V��fч��i�t$�߽�eׅO|=]"��a-ql4�.��i=~��-_�^��'	�%��7]��A��c�V=��o%���p��{�J�I�;��A0x�X/eV�����rsX�rÑ����z�l���?�΃���bN��gQS�~;��bͲ��e���u/�f�g�E��&p��_�3k\�b����& �D9�Wj�Kܱ���]t����:r����ڗP�,e�В+lMڧz�b�K"�e��ɋ�� b.h��.���s}��O�f���Jy���Jϐ��˘_�����sF��Me�$b6D}����9c��N᳒��	���5Q'�;�f��U,qR)�@�,�︥��<�P\NE �s@�;�Ɵ��M��ou���,��#�O��v�jDV�_���7���y�2��C����y��!���Kz�L�a�@���*��d
�vXMb=��8#��^)�1B���5�	��U�Rl�@��bLӖr"��X���Ś�d���}~9�֔ű	v���
�%t��E]�ů����e!̔�I�.4�	{��`s$�ȶI&��B�T?����@7/����e�P�\�}U��;-ثpP����0�Tnݑs�ꈓc����3�+ÉT���3R�0�U���K�$����X��'w�P2���e
m#��Iv��ϏT�̈����)i���w�d�O���t@<3��C튡�-PF*09� z�.��`���"k]켔����!ȼ�a{��
e�oRԓ���2�֩Us��è�d)����h�fAe�Ō��p�j�m=0.�>�����������l����t"��JgU^�D+xpp6��栠흆���_7C��-�\~E�A��B]�^`��.���<��?���@��� �v�;���3� 4l��-pH���l�������[������U��,�PA���{�ǩF@�cK��4p�t�W���S\S�!�!Q|�-D�C�I�@���t�^A����ev�
��K���TR&0��tB��U�3�> ��ާ���3�V?���E� ���o(iГ���4 �ċ;�?dn(g1�/��j���O
��=|�9�g��G@��羒O�D�
uR��u�~Ϸ
o5(ˁ�d��q�d|ڇi�k��a��]dE+ώ�B�E?��B�\{A:�H��C�%>���`��qD���ɨ���w���P�p3fMZ��x9۪�T�ج�O�UKi:у�ҭ��9��ٴ���̶8�9��&|��Kر�8�k��U����1���\��ܻ�Ӏh�zP����H�1�2�Y��nm�u|p:&Ǚ%G��x737��z���b�.��(?n��<��S?���
��@x�I���[�~�9K^��h샛���n�ZUPc��_��EU\jo�������&,�#D��KُF�GB������ru�����\^�۝���J-F��i�Q�l2���+�vs�7��ʔ�)�Z���{@��W����n��5�J�m^>�(�w:=E�e�+^8#�`��+R���S"pu�[��l{��6�����Fa�1�.�jQʘ�`d�}���Ґ�B��`^��c�a�ᭁ:*�r��D�7�	�������%V�L �w����k*���j�C_�|R	<��7Z���0��%y�<���`%�s�9��]�	�g$Q�9��^f����.�1�e�X�r���22�G����I���J�)O���qt�E�\/�V�MM=�V2k�i6woUa�*
���%
)�9,OT2�$w2yE!*��G����AX6�J�f�K6V��u�2L@>B�{�Ovw
na��QJ�y�8���&%���)v�{JЈ����*��:6B�-�*�.������B�
��1]?���M�k^���_�z�ރkև<��Ҫ��_�Q�*���F����C�hz�wE��[RL/�c?;�l[U����
�{�3o�VKVw+P�]��[	HZ7��h�e�q�x�W�x}6P�
UˉՇ�S�a
�{��~����D����9��۟�ꈘ~�$j�>��U:��w���D������*�~�tܐ�z臄�'=�"j���p|J]7i�Y����00���J�З�2�;�]R9зԍ�3���4 �:��g�}G��?�c��`��])5,��|T��Ĳ��t���iTuߨN3x��e��Ȗ�K��n=]uؒ haU �0�"�m��
P������^5��E��u��F�I@n�ƫ}M)Y�� w����vս{�xP$��q7x�D�o�����q'������)~ p����'�[�tiڼ637��� ����x�o����*Ь�N�����4��0W�I�l������i��j��T�*A�x��Pp*��jG܉,�<�a~V="7e�6�~b$ �s
��_��닁�]�܆������e�v&���/�t9S]����w��K�lӐ��i��o���4.ɢA�N����,4ɥ�­I�g!{���G��w9�L�㽥D�җ���a��g��`���gk�dܪ�`��U�{�VD�y)�ܰo`CN��*b+�7c��}��"w��3
�p�V&����u��h�����
����T�&���F�T������h���臄���CvW��<�|���|Dd�A��G�
�E�c��R��a���RT��%�C��{�ɾ27u��z�`)9I̮0�g��5J��e0kɍE���~o$}��
�`�6��q��6�"(v'u��<�	�����8=�#Y�7�sH��ʙ��������-Cl s�m �i��A���b��t}ϼMǃ�sbAo�3��˭��(�/�ܞ1�r"8�qas5v�2�-��^���쪎��"��s,���P�"p�Z�"ꨑ~��KN�ם@w1��h]P�3�_���4�D���c��~(~�3���L��m����5jy�F\�W���|��(��lx$��K�/��=}�4>1O����AZ)�i�2��-��+}Ͱ}dt�m\&$�~�+��Ⱥ#��QR���oa�%�p��ʇ'��X,�B#٬�dyGְg,P�J*~p��y������Zq��lZ�����O;���^b�+��ƪ��'/CY����M��P�(y��o����*xe�Y�W��I�BgnG�5�,�f�U��B�hq<dGM# �^A�Q��AU�	?�V����	f��
�B޳��a=xgZ����)zR|8 �}\	�ka�y"Z�?֋������ ��;&|�G|B($���0����*�,N�ӄ���p�wC���?
U}�t��c��8�f��">*U��MB�=�|��k�����ǰ߅Ɏ�R8l�=�s�M]��)%����{��n0��y�K���Ӂ�Eq�#���g�q�,g�]lb�F�;�0)BZ�o�ʕ����4z��r����@�z�Vhf��6�+U�+n�#�8��V�[�-Ē��9��q޽�]"���$ug���O�q"�6e>�H,��0�ݼ������P'e�Ȝ��Đ>*�)t����^"y�=��nAbK��0cO�����gZ� 0�<�ichS�m��矓I�<�ӁE	<`8�����|����Y�L���Z`��\�l?�}Q���]F�Fx���Ց7+��1��6��*�����Y,�������q�&�	��$��*7Լ��`-�;Ez���$����@��Z�IY����2�5���M��G]�L6e�F�-z�V^�oi���������#r.M�;���y �_d�4q#��FK8��6:+äI�����U�af��o\p:��ke8�� ΄Vt2`PW����+mz��Le����l����5#8�?�X�9+R�7>XWT�$:�N$Qs�w�y~��5p&^�%>��o7����Gu? ��n��|+�8����1����2=��0X̤@'�U�R��ٝ�	��X���iO�U?�a���bQR�Q��V6V��ttH��A�.��������i�D�}�NWl��k5���wض1�ջLn`��g����E%��-6m�Bv62��Z��=n+�P_p�~IsOV�D
�b�Bq�܃���L�l��m����ǽ��fw���21��9���R�QACd�SuX�'C7�0�f3�
>:��h`5f
�mh���qFɴ���8��[MZ�g��%��M��Ԕ4M��О-��l�l�m�J�_�XT	�̖%����%��KP9#.) ��T�t;Z0 FK�<	�7@EW��%~�;�хh*n���Aucκ�ep�Mܺ��C�!f��VI�t����t�����9@3��?��m���(�C7q�w�y��@$�"w�U��ˋ�n��S���G��5�F����-��ۘ�6J��[�}ރ���n�z�L���,�9+r�������޾j��	X>�m���e�����-*4��ә-.�]kI����ۂb�b1g����1�J���)4���,Qӥ��ɑ u.��8wj`.�9J�"������ly��8G�A�� �K+�X[R-�&�'��L��^컻�@e�$B�-m�V+a�u�Pd��m Wl��j�g~<w<AG�Br�g�z(��/�~#�V5U<�5�è�ؼ*ۊ�M����"v��UKخ(���"Oj �F�/K��T���F��%�M�e;�W����1?v.+;��	�%P�|�8��4k������Z&���d�3%�ˬ���/������ͼ�_*�k3��l�ֱ2�g��&X9e}\�ap��h�|6�w�Qh.ˏwqW�S.��V������t�n����?6S�~�ω}_6�̀,KY:�����`����o/����蛢I?���5��?�Vꃱ�E�e��^x�o�[I7�3A����`�J'J=suRB%Z�u��Jg\�EwC�Zޟmǆ��&�ɱ����Q�����7�} 	�el׈�7잉m�i�Β<����m�L2��XE�c�#8���'nX�|��?�7�H�뷯�)	<D�����J۵� 
���]$�%�P򛵯j�B&՗� �aMwf#G${U+�A�˷�B���JUug9�F�ͺ'wD��`[���P����C����É���
��à��REP墱�cCu���]���~M�v镳�	�a�f�s�(��:9��i�M�� ǊJxR0Ê�W)kg&�9�f��r�*�?sn� �R��6*E�=�v?--na���CYUC�uY�c5X�ly�>3��������|�����dc\6_o��L�����mPv tCHc�{s�]ґ�S�ӆ`ѥ7 �8砦����Jr{CgZ�w�7���FH��N	o[�4\O�������ф���q�ͿT����,��c�C���,"R~Ĳw����'��$,��C|y7�9�`�ca�>B���Z.F�3)e���Z��O*��j
�صi�Nǰ�a����^�Y�K�D"��U�i��[j��8����J��n6�Gf4*=�����4l�>W�}��.A�ę����R6��x���X,��ƑɴB
5�?\���;�� ��-��C��V]���T�e��I��b�A��jn���6[�0�����`O"]�3_9?����Gҭ��Ã���{�=U�lIYd��+F��ҰM֝�:(�R�7Y�����tRXf>{��ʧїcI%5�xu7p�VbJ���9�r��7Vv(��Ƨ��O����\��<���䵟�8�O�H6��H�:ߠ��r���2�߱�̓ȝ�T3���_�z%����KS�c
\��I���GkBMg-\�.���I�[o;\�ÜÕ�w=��JBI��׃��8t�BH���8�2����v)�_���1�����o!U��{ZS���>�+^R����6���3��_Oks�[S% �1��C����ք�;��d�A�wե�~T<WvQC������1ǒ��Kt��V'��F)����{�5�PL'��x��<�w/�d`�t�˗i�k=��|a͝�Mͪ����?y���ӑ�֪�>���"�����R،H'�		t����Kb�9�_�4��D����gG���
�A|�ߙw�l=�%��2���ƃ�[���r/��U
��������/%��:~ަ7in�zh��/�>N���L옐�k�����Q��4t���_���Ӝ�5��,7$�nΕ:FT8J��)?c��f�M�DI֭n�VC�f��A������0�d���3�nxc�'OΈ��#���N������Z��-���	'/����{m'P��W]:v�q��	�������)ٙw��$釕]���!A`O���#�0|ÖM���^�/D�w�.ש* FL�m�i�Q�m����h���6��� #Q]�~��E?���1�ɜ��&烕�0dݶ`�Yw�=�F#��<��)Շ�}�_��Ir�9�D�!�Øi�����[�pi��f���(�%����D��x�CR���\�Z��m?�d�c�8נ��i�@��Y�<AE"���pJ��L�`1Efܔ<�qG��30���8Ǆ��J&�a@N��L�q#O'Sa^�-S�Z'ܹG��ͯ <xZp�8�Rφ "�F�HϢ���B�/�F��^ b��0N}->�f��l�>�C'u�"ZX�?�۰	�����5O,��(��"k��3�gI-�i�ݹ��u��6�.���C�k9��0��8}�ߙ��I��|i/�~S�&D���N��0���\��h"5��7��I//c����ó6t�#)|8�C��D�j ��d�m"f���}��o�tO>c�z��ԭi��\��T���(��˒��kc8��m�,S���QZ��%��l7a7͝O������Gj�%�諦�BI�Z�酣�j�:���H�Ɠ�������d�aհ�rzTٞ��2w��%�~���Ge���x�RR����c:+T$ �5[�������B2!�;�0���ϰ,��Gn��a���ׇ�)���2��\�����Qܹ�{E�f��i�8����u�"Bp�H����+}\��~�,���&�sW^w�IúII�r1f=�(�2��� �]?��9�TY1��%���n�V�����I�v� ����3tH#0�	έ���QP	��6�u�N�nʖB|��z<�W�]k�KZ.~)�Ӱo�!t� p5�7�����>��p�/w���.]R1��]����_\�-�)��lk���緧�E"����LxE��Q��z�>�'�������Io[X�-���]�k����?�pm96�_^�2�z��+u��EU���8���-�e����+Zc�ƷC6�W<�b�v���ӄx���+O�h�3�T��~�3��2�A���8����7t:cA;�)��1�م\�@�D̯m�؜�]��r���d#��t�ڨ�֟��n� Vz��=�4@�����)%6���W/Ipx�K$�զtj≀O�<7]=7#�g�do�:�T3���a_��b����[ޓa9"x啃���8���m_J�g90��ʂFl� ���G��-�{-n�1+uO�g"�S��FL5����@���)��|hU}9!�7K�����P3ު#F�>4[���۬5vn߷&�����G�T��!���@%��ބ6K�ᘶᱲ@�b�b���չ
�w�O�X/I�{}��3�ݲ�3�3XU�J-4F��\�R�}�q}>�3�fi¢���������,��@%�xσ�͞U#C[4_5����2��N{�%b� �iM�]u:m)Ố�T0��ߕh)�MA:�SK��Z�4�g���S[?��s����p�1A|3�����,��n*�~��΢f\�y����,���t�ux4`�jQ�ʐ&�|����a��O��v��&��Ʀde_��&i�R��!#�l�\�&�.E���$.	{����`4�� �C�E .z�. ���/ߕ��
�'��zG?;pa�I��m�d�ԸM⒋U#����Q���!���B%}<�/�9ys��>��?+�*"��)�$��{��S୹k3��`�V��Ի��ˏB](2��ἴ�].��`�nr��{ ~�z��(]�>���`u3!�|�UkI}\P��k��f�!�k�ϲ��u��3���8�#�u|� -Uo�d����9��Xf��L�*��-D���{��=*�eʰ�OOך���W�ט���;˙:1�4,�C�N҄�+�^E��sFߎV�o{��ӕg�8&�l�-�=^��<j�_���P�<<�YP����5일2e���Ūf�'%mC|s��Fv"��?!SY/����)��������tJZV��C7�f �������U���9�V]�#�ؼ޾.��T��5�=-���zy�b�Zy�;����|��Ƨ�Qd�ҫ%[;i�����[R+�y��@cR!M�1�6�E5����J�om��#��BS���V��,�|s��[���F��iM��h5����1���ru��yK�Q��w\ǟ������1!D��IL'iw!V��>˳��ö<�.�H+�V_��q�6^����s�G$��[fӈ�F7��8ц� �|6;����;%sW#�h�$;�[sz��!��='�ʨ�;Ǝ���>�#h��z�I�r���i4[��Z��h�=GW1���a�� ��1���G!Q^��b��#r�
Q쟑&���`�'* ���V:��~Qc���J���W��'(����d���up6ؖN��˕�.S�{#��U9}��_�D���%E0*��B�}D�h�=��Dp�q�@�z�+�_؂���ו*���J��:�$�;���V%̏ۍJ�e��w.����vm44�f_��q�y�K���y1p��.;ɠ<id�,H��!-��a8Ac���������]�;�{��P
��l���8%��3��Z-�Tש�"�w�Ók��G���>t�ӡ;��&�bw����b
����q�a�i�η�F.}uEqɊ�W�T$P��&�{��Os[����m�x���t�p��%�
�P6�Zp��X/��x�%�(;1�eAC6��_¸����
B�H��a�DH�@�n����n���Ur��2��kd]��mG۪��2�Bu�mnB*Pc�<�(���n�CW���L�'%yQ6�i����4<�d�j�K��ʉM�&b��6���!S���j�.hR&�g�I�z �rRjqQ�4-Oa�����J�,t����ֲ~"��Q?v��"u��\p{h$�Q��*t��>r0�����y�O͂���U����Nz�BZ&�R�8zRBK���Rn�c�<A�3�ë���ҡc�6X����,ϱ���`cx��?��;+VE������D��W�ǜ���	?�8��j��i�O��]�a!cl4���/���ߦ�]%�����_X<n��N�	oj-�n_�ԕD�b�w�:ߝ`��{(�v?<��2��ǦE�~����yf�s�c�gv�h0J4n���1�$� ��g0$t	�A(���q%���j�qV/�a=���'�4Dj��F:��	��"�6��Mhi�P��'6w+J+�Hw���g�u"!Y�'���n^�i �2,T��>泽�H��s��6ҷu�����^���Н�V���ڏ&Ь;�H�15�J�4D��2�V�pϙ"�0?1�2mU�eJG��r��T���l��6��_���@��c�JU�S������\<4=�^?>�g�O���_jf��d�f�x@]ų��A��%�%;�ێ_wZYd3�4���{���#S��NKN���a�Х��W��P��|������s��]p9?��8�/��Ɲ���O�̛�M�U�<�=j�JfDj��1ϕ-i �s�A�. � �2�{	W�����)�g��z(���,�*6<�Z��cJ�Y�V'-Y�!���n<��͎۟�j�$� ����� �k˽��.�	�e\Y���F���d#�v���=��HIAU��vZ�Ԉ'%
sIM�8�fLSE�M}�sxtՄC��)��F���u���>��ns�9�$h+�l�0�@yn0��oG���Ee���U�ڹ5S��1�1j7��� y��c�<w~x>y�3�_~�C�gހ��c�����βK"L

Pj^5|�u%}S�jݽ�Λ���Jd��y�ft0$��c�"Fns*1J
 ��l��	�=����-����4&�oz�Cj?_�ӵ���M�0��@����E�]X�5/M�U5��b�A�憯�����RC?�j͍�L���9�
��8s�����#m�\;�����G_���?%�3��X�1�TY~+���,n�ř}[�N���i$E�{�J:3O�V}���|6"�]S��-�����rf��[i�c�)�}��Y�iR�->}�"��+&�h�p��x�J,d-_�ܴB3@]V̮@�iN���	>�d]�=����KA��"Ty�&�K��h��1ų<!�!GF�%y���2wԸ�����M�B�^n ��!67�������m[�n�R��H�����L;d:M�Cy��ee�[�%�X+�mh��u@�im �u�ҫ�o��or�uR��p(�X��n/�����%�Q���N�����>���i��M���3O�"����Hl��7Z�l[v��Z��l���*�FZb��ٓ�S�h7[.�;�.��C@����G���D,3�?�Z*���=��4��L��ESǛf �I1��הt�']*�a�w�j����3��%xdވ����˶>�����<wuZ���=��j��i뙖���F1���	�=���d��;g��-%n*�/����5��Oߺe7�҅�`�
����J���u����.�b��ԛa�5����$1�	&C��V�B�2�q_S̿����僯�)��h}"j�B��|cp65'�O_)GK]��K����8oAz����?�Z{���Ț�'Ii�_~˪��eU]�/�X)�2�����t�r������1�2&�=Ʀ���Z�_q_rh��{i���W��n����'Q幱B��0�&;ܷ��5v����w�b���n3\g�~��^�MG��3�u$�(��B^��Vx�\Q�z9����v�%���9�cb��
�J���i}�!�l�e�������%�6����֫�l���d���c!HA��Z��!v��j��m/�~�уc��|�E����I'Tj����U��{W�Ҟ&�6������b�dB\��.�l��h�|�wE�!\��ED)4�G�z|�	�7�I����{�w���R��.���%9{��mxX/�J�	r"k@U�h�
��Υ�#�0"�M����<U* �K墪-$�\+�or4Y����зx{���O�B��lJ�b?B��so�5$���{Z&�Q���y��5'X�M����g������Q�b�<���O�4v<=�ĭ$�l����Nc�I:����J�#�g��|��.5'@�?��do�R}�K0��S$�a��oFZ"ݬ��/-����	�2�otS�)��@�`�*�X�dp�]Wm����ӊg�D�!�U@�����cF��%�
�46+������W���m�����M�hs��R��:�n�o|{I|�����4D�Z���op-�q]7�͒$�ct�<�c��s3q1�{��u�+���T��
��r qD^�kl��|��%)T�T�m�yiwE$�L�2��S����3��u��cR3;�����|�>�(N2�lR���k�_�t��d�ؾ�����]M��1�i�[m뚘!!�e��*���v����@���ph��X���w������y((�C��et�"��qR����Xw]l^��ª7� 3m�[^[��r�)`}��g�Z�����ؗF�т���[>�a��=N��^�+pMт�Q�3�e*LY��Hc��2�F0�$UfN�R� (,t���c�>Z����F������
��魄�JuU9H�`��; Ӊ�A���U��sS������Pȅ�=3��~AR�����З$Kmt�Y��휽%��sAQ*[B�8}>��D��;��q��M�	{*���N��9��>'�l�ȸڮ�O^�5�����m~0RĈxM���X���}��c�ZTb�A�[�������';Da�����%��U�$n���pO���'T���3Mz�¡��W߃ R�ɿ�2R!
�T��6�U=��9��C����R�O��p�Zn��c��;�&<= ]�|Q����=�؍