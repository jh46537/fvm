��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb�����jA����'J��V-�@m��Yx�W����A�.�ƋB8/dq�4z
��»Ø�;����/�?;H�G�ai���'3-D=R��@���\�&�A����w���.�yI6����˗�UF��%�T��巎����몢����®\&Չ5W=KA��ޅ,bF�?N�~�o{�K��\�̪@Қ7�h���%��ԐEktU@"�BSیv�z�#���d'Q���GޕF9���9����Ե�@��t�u����򯜈[�i��y?h��{+���<s�h�!���.F�%f��ڋZ�ie�:0Sgp��av��pxь����ɝ�ihIeH�G��ꮇ �j�yC+���T����i3Dؒ�0��~�R-�����Oqlo^�����ʳRo�3,���;���?Z�R���j5�Ԭ7�k���*�	�{A�sz�P����:fc(����=?@�n�F*�6��{�L8��P%��_��Q�*��N��ay���#�D�Ďχy#�m0���韪U���r�L�+�7a捦�N]�Rr����@�ǗC�"���������a1 �D��
��v'�E:�8�N��ApQ����#�8[2�������EL����1� e��6B���|��|�x���������h�F?z�% w^no@�����v)y�LS\���Ɏ�k���U}W��)���,(d鄺�2�_��fU-=0E�H��Z�`�����+Yۊ��S�O^#���4|#�nd�Bu�8�p�F����dsEԢl�:��: ��W5����|zZL>���G�8��ݟۤ*"pk��6v�!�3F���g�b����s{�	��W��w���M�!�U�I��;uN��ހ��ޏ�ן�\OSr�j%,�uP����`,C�>L��!J�7�w��(	W)a=*˭aQ��!�`��ܣ,���|��riJ�T�4�]�q���ڟ�{{���j#�l��`;4��7����ײ5%X/Ȼ;����G�&�	`o��M��4m����*���;��o`�k6��'ק�|>~z����e���|�ޕ��MR U���}�?�,�1�m��g6��bnW��� �3�j��r^M�`�I�J���tbjiF'���B�_v��v�y?i�#�xjH��<>�qd�ZT"�=k
�u0�1q��PbА����͡L��ph9U4@Q0R�>�z8:c)|v
���`9azXJ=����Ef`I$�����p%|��\�Ea�:zU��͝"$���&�+۲-����^�wM��n��|�*�uN� �D���^�j����p��\H'O6�����S�s�J��C��G�<"Cy\�fjӢi?�`\�}�pq�(�Gڙ��F��m��I��L�w�^�g�&pF�{�E�e��/�O��;/C��uת&��]T��! yNK"=�l��dk�O�뻱|4��!��$K�F�!ʍԵ��H^�b2�<������g�t^Kc\�~��H�04�G �~����lDxV���΋���+C�m*�UL�)Q��*O�I����o��I�1��O+�;?p�r����~Q7y�X�.��� �>�{�{_�o���;1ъ��q^d��m,Xe����F��taS�9�;T�8����">>�j�;ڮX\�A�]ND�� ������lyހ�	�yVmw��<��D:�$�C�}�cv���^S�<�A}2��w񚺧�˧�qu�����CV�(N�4̋�h�VYω4�b����t���{��Y�jE�V�K����G��`��w��i�<K�C�W�8�t��X������+
���M�e�n�l��p.���Y�O�ca@9F	5�i��O��@�}�] �~�SHZwkY��eUeS���#~	@$��� ���5��-�7��"���2�p�
��Nt^�U�mσ��f$%P�)�,pWQIQu��?7�Co���xފ���O̹��|y�J)@ɋ¾,��iQ��\W���4{��!����C��VV�"�&�~l��s�:��3ж�< ,����>wF4Q�55_x����H���}�ƭ�>�w�؞��e���D}�?�~�	��!5�9�Ǹ�v��OwAg�d)C�8��g~��׽�x �{=����R��&�<��;�HcG�.r�-}���7�#��D� ��,����A♗}lH0l�����w*�\��-o}{�(��-�#[���d�I�5%�B�r6�u0`Za��\�x=	�\��?,�@�Gt�!��aŪ�on��/�p �ҳLAe����V�$τ�$�9�	\v���M�zJ�h�q��]�W�$�v�h��qu)f<갠5Ӏ$�Ӊ��|@�^%���#��{Л0�Y������ȴwk���0.p$�LW�C=Ն�ɠ>A��7�-umUOwmW4�fcp-��p	�c��A�ީ{��`��<����Jqx�����$;����0x��,,q!,!^'���^y�]�=DԐ��SʻӍ�J����/�����ޙvL&�S.g[6(~�pa��AY �⿷��k�ph&9J,^��
'�l��ț?J��;wd�~��a�Pu��9 0�A�S��!F����.*L�g��-{��U]��RM��{���͵�+U�3.Rf���s��)6E�YY��q�����78n�L�j!�n� g#j�ࢯ��t.	�j���8��W"8B��͋��G�*�D��j3�{F�������c ���2�%��ėa&Z�Fn�%�.��C@�����B��m�v+��Tү
�ypfrK3���S)e�|����EFXT��O�G�I��O��jӌd��;!��q%��aiX6+2t=�A�OI�}twՀ����ӑ���}Źyٷ��!K�}/�e�Σ�W�_ֻ�}_�3x�M��p��L]u�������~UtlC���E�|ϥ9R>v������r-9,|�i�=,�@�Ɵ;E�1go���/#G��#嘯9OI��҉�>4Z���[���W%���������~Ү����)nX	�c�$��x��+��w�]e�tм
�@�꾸)|��N3R���F3�������x�E�����?c٭=�$>)ߑ	�s���̐�����R�LGk^|�;��#DG�Y�"��[�0�ha]|�N�a�*HU<,��@��� >9��<���
�E�Y|>���91�#������G���ͷ�F�!�nF�ϨN�\	�B[G	1{ߖ�u�&�2-�� *�1�YE9��з�=�x�#�w��BC��t<  �*ρ bY#�&���w���F��s�}��.h]%,N�lWe�A�&>���ı�ڎ-��#e,��:C����bam�>�P��a:]����bqoF�Yݴ%%��CH�@�m�/HR�E�R�o)��|�3���oD	�ET:�HM3�,�,6l|r�FEBDp�zAߌ�*�n��	�F.�aR��M��l��h��pڤ��}�
�@�c�)F�#���=�@�{H$��o!����D�<�����)u�@3�@� L�w$p���Q��0y_�F)�5!��Ӿ�οݏp�:8$�u�]�2�_����Ǿ�����ڔ�T2��
M�A����:�}�hg���iL�] �6
I��i;g���� h^i�JL�G}^�w��Y�K�7�`Ŧ��%�l�������z��|�=ʰN�,����-�3xT%ЭL��<���w��$"��	��|�U�4f{E*���G�$ޞ>I�8�P�6����� ����!xyѣ�g�3�б]��=��'HF���#��>1j^�6��ȱ�9HU����ٮ�������6=����T�0r�ݘׇS_<-ܛ��Y�����~de���l5Tb��>I��b7;�k�M�
[e���c�uԻH��X�&{��k2JPMm��m72b ��zJyXC(�qJ��߆O�.�#��.DIx��VV���C"��LD�h<W�zSP%���7Vx&y�b�8�'۬��ˣ�9㿂"��PǘM����_vI/ ۭ��������mSԌ�ׂ\�n|�X���^�g�m�B����o3-��O-�����v��i��r�>{�ǅ�[�Q���JH���FB�r�,����b��ۣ��7�!�h)��ϛ�|����tI8z
�(�\�o�"�x>�Yӊ��eC�(��Ϛ�\~T^?e�u�D�A̅<�h���U$���/:B(Ϫ��nQ<a�j�`N/

_8p�����2���\#2�(w��Y�M�cp��~&��0-�;B��B=����cR�[Z�p�S�?�"����&r2�a�W�
�q��:B݂�4椁wno
�9%����/TK��`4O��]@�;����F-uI:��������%�(m����&�n�Y�+j�9���Rh�߽%����4k���O={k)��ό+���3�_��(q;�"u<'5�*v[�I���
Z҅'ukC`��..�e|'���~\J^�Âv�qL|��Yty�,�Xe��$��u|���K���b�ehdJ�L̀���<��k��:���O�u轮a�~$���'��4T�~�u_���qZ��6JM4ZX�X{1�_�F�z�Ol���4���@�Nt��C�|^K3���CU�0P<O�l��^|��2ei����R_�*��d��n�h���f �z�T[�OW3�:K�����ث}�I)1e�ut��������/0�������p�')��ׯ,?�?�����ͫUGq�׏����0Q2z@O�t�F���gvE��*��0Ʃ���hl��k,�X���h�Z)+)�4�5'ł��G9�>޶	h��W���_�VT�j����I�!�!�� �(�ECӐ�_��d�!x�5���=J��5�o�c����,�A�\y��i[�����j����8=f[x�'7%M����Κ?��n���t�
�B��E��b�r# 6BA�TY$Ӳ�L��k�悅Q6hzbTye����?�[���~�
���ž$�:��?�Y�cil��':�Q���ُe�,U�[�/�
��rZYy��|s�w{f�ǅM�
�����PD��a�K����of�d]�ޭy�֦��|p�a۹�X�W�Y���߾��C��&�N\��<&���δ��&����:�9��;����mOѤ�W�z͗��7��B�Z��R�D��4ɐ֯��y����^n��]��<�`��un[�L-~?�&����h��
Ojnk	��^��@�