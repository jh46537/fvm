��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽���^(2�� +]�ݻ;;�w��>vO��@e�@?_ï�9d�|IF1|��}L�k�|�Z�Qy��I)UP��"=O���T�D&[ݥXa3 .�X/��� ��DF��!��X��2=`6�l�gQuƄh�Q;��j���h�u���!����sF�|��j(�xs=���W���	����+��E�ʹ(�ir��0�D#u|z��%��m���a�gO�I}���n�+NK�S�x²y�ρ�����5Wo�	].��B�����b����R���I�F�����f)N��U�N���[W��S9z𘥵�#B���T�z.�$��=HzJ�&MuӚ5l����CN������\��G�AK�8�yH�~
�B��������5��ͯ�h|X%o�p�uw X�´)��>2@��0�]Ӗ���<?~�#B/�;)ݒ'�E'-���  (ؐyIC��7��	��f�7���`���r��E)��,�R�C�cg�P���|��S?�6�B��k�o�~��	mb����S��Aq�8�GK�
��~�*$�K}�Q,~οg�����p���E�����ʵ��Z�oy.��)D���i�ԳN�s��a�=��o^��p�3�q�,R5"fTQMܹ�Q���G�j��輴�:��[�[��{Q�ڼ�»��7y�?�M��`Nj�Ei+��[�x���?Z��˔4�e��{�GX.��X�i^�^QK����>"��b+�.w�������Q�7�)�m������b�n�r�ﵭ��$C|��ꯍ{?�hV}G�i�����a8{i@������G�L�8���$���ʬ�,3��2iu���j�I2=q���K�IRcX�e0T.����c!�1��;�L�.]1�J��O�(���@C��"�=���ۻ�Uv��(J��]F$�h�[�S�+����lzEK`m該f��l>�j�uJ��0�l#�O��f����w����Kz��0A�Y�c��7�e��w���˚)r���fꙺn�i�������c��O�$&�4yz]��*�ȉ݁�RC�K��1��A���%�˻� xMD)z�/b�'qw��0rg_�a1�B��#];�M������u]�ʭQ��h�fs�P�g��M`9�������**�
)��4�=o4M%���ј.B�_~�c�Q�[q�>���U�-��a�.��n�>��J�u�6������,�~qX��v1Du�'�ٗG���DtF�(d*���R�O��!�yb�z6�|�j��JH��M1���lV`z�;����Ы�exM����cCb���Kp�l1m��vGxf�ھل!݀�£�:D_��
�� �`�"��EL���3A�Nr�g����<6�N-rL�u����ƭ;mm��I�ǻ�
�bc&l��8^�H"��L��	�Ĕ?��O�?2�8U ��kրų�Ւ��+:*���[�w��Z?�u�Vs�~��`����{�*~��2��iP<�l�[�蝐�g��m��1�~*�u0LI�٦ѳN�l�������z�<��y�Z�;8����(6%} #�a�薁Kyu��5�2�l�����'�gE�۷��W��3����y�i0����3k���;{FO��)9 $WQ#�HP��0����oRX��B��Ė�퇕�9�-���D3!���.f40��Q#^�+戮6<W9�� ��'@V�q�p���
'�z��ί�m

�Ӏ#:���·���q8s�M�I�<�q�z�/���� ��&J��F��y=d�G��#��0D٢����M�.���(�C\$�0��p%�`?{O[Uoڣ�<�_aa7�W_`��#3��]ӗ<��TȘ�DƮ��V�r۳Z�y>vI��C��-�tE���0T�?y���������|FO�.����aC{,�\@����ó�O:�=��5ˋ�N�.��t�>y��ê�]�T246���~p�E���5��k�-�]�=OȊ^�f�� ����o��&B+��S��#�(�.�e+���ƴqg��6C��2D��.y�]��2W��i�f�E�����!sݪh��Y�o�^ir!����f�E/�J��D	
���������"+e
�nnx�K@T�R����sLL]�<x��7�@��e�4�6����|�Brk=�V��t�����,��&;ǻ����.z�(�bO�+a�R;I��'ѡ��;�-!�_�zi�?��~p��7"�G�d���U�uU09uZ�J#��p��T�k�h-(�`,����G?���L�B ��h��X:����G!���*ҁ3}Z���v�V �GG�9^�X��K~�+�U��B���yLevӷ�_0b��R����$a|`^��{��'�A��������ЗL�&�
No,���Mђ�3 ���S��HR� ��f؆_#��΍��|��7K��.R�v*��Q��_�QQ�� ���։O����!71�8>:`3��ޔv�Q��6/�x��MC{�JUw?�f^U>�K�V����"��OA����p��|��&�g��n���0�g���u�t�o�.::HL���Ŋ����9h�ۆQ7��|t.�Ђ\�