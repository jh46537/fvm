��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�
��)����\VH7�d��:q��Z��
�'��Rl3(N�~`$�u�V����I��t���Y'��W"���<s ϓ�T�F?���-�ܚX==@c8�j	qPH�	��\�`���Y�ÿд�9a*�Z�Y+up��Nɕ�f�����4�e�͊Qm���A�|�v�H�v�Յ���J��P��M�븓Dp6���8Y��<Bfo3��$'���rVn�}��
]�FMu�� RF�9��d��\`?��	لZ�i+���1��Pz��;�����f�76F����,�8\�TUMupé;�f���/ƈ�~:�YB�"���h�W�s�s!z�(V�r���#l1�˲��IT� �v����ǿ6�%�D�����̊��� u���A�t�,Z��d���7� B��7�t�xQ1�|�n���?8�[9ۘ��?�� ���f�ʅ���ڹ.hf���T�8Ĥ�����lH��R/�M��ߛNսK���bL�1�2/"C��w��o��J��(�02�
-fZ��h����/�^���*�������DuB`J~�����d��������8"�3����2���.�O���:ϝ�nP�?6��k�y���Fq]�egh|�@�'���yH�P��k�ob!�*+��y'M�K�D�8��jl�i�7����}��Ӥ�c�C�?�:R(\"��7�S�E"��GE�u�ߺ���>;�=�~�74������Ifq���Z��il�G���'o%�gd,�����X�XU���/
��OpuyT���qd`�f���4t"�05�8�.����Y^��L�h7�L�� E���VQ�.�Ar9L�[�d�qAUZ3���c< ��K�S}����[L�7��Y@�r�5���{x����O����ag��Dx�"?��;��s����wg��'�p��-�"������Ɲh#���
�_G@��R �6���{9�?�����S��۠����c {���]3���	�s� a��.YZ D֓��GOCy��ͮ��0�o�Z����9��u�~�#�f�|��HK�UD�v	��&Z+ZU�j�A��U�>\E�c)g���&�9�0<Ox$�0i0���✦��LLhR�r�V��q��Н�,r���g�UD
���{���}!�L$V��������z�����J���2_���� Ô�_�T�|��l���V0W$�9N��q��>�.�� �Q"��m~�?;��˄��>�H��~��a��*S�����\����'��Kb�pu�zH��3��Y���w�~ʀ�n����}됳/⾏Z`�j���s!��/�n�	�J����
R堀��ҏӰs�ѵ��fẀ �}K}�n>Iͬ9	n�]��D�qԞ�6�^�t@Y�M�*��5�W�%���)۵o)��e7r�w��kU����U�"��B<�u���3�o�XåP���"�L���{F#u?��X�}�S�^cn�d �PC��! W��(�C�E���0hF�9W=V��8d��!�Qu��p�##���*ֻ<���kW��P��~0�^��P�7���Ҫ��M��I�Ԫ��֞��pl�P�����r�2k�iI������UjC�-7���)-�+��̶���mQ[�/��b���n�-��l�p"��r�L�8H��5*M��ɖ��!r��_����'� 96�dM�n4K-.�!H�w��ǟsy�zc'd{���� �7��,��y�vn߱��-�{����� _b�H�����lS��,�됶&�a�uٳ��sUD�Rm莀��a�6=iPҍ����ڋa�uwD�u�~&�)��Ƶ[	�0X��f5�c�q}�I�|�n��2%�{�"�~����,V���f�(�^�{;�^{���Z�u�ce,v,Jva"�}9���n=&H`蕋o~h?͔%�P�&�射��v�w=�������~Rm����Հi4J���6q�$�H��,�� Re���,*:�Y���*�A��"�l.Z��3SE�J�ߣ��iO��n����j�5��ƹ��kml�S)���pS���mꋢsS����Cwxxʥ�]���Hw��~.	�/� �]R����al����ue�Bbci��	j�EȨ#<�M��ލİ~K۔�2��)�by��ڸ�9��2m=�UléCSz��:@��}�&��E��L����$��3��'G��?Tk��+2�J �֯�,����}�(֙�%+~�ฎ�x��m�s=FSN�Z��Z%�mV��!N��
o�J�$�?���>ܕ �Ps%ԽJ�q���̕ TS����Կ�FK��f�i�����C��U��v #�T��Dx1߼�A��vd8�Za�K,��zKcI:����6<�����y��B�(}sd����4�y5�U�篅'��2+X�Zkb�
��j�� �R���dK<[�Y2
��>����=�1*^��ft��\�����h��Y���?B&�U$PWl44yZβ|����O����C�]0b��Zcz��-�ڥV��#��F�@��b�X��P0�_A��b�F�U}���@�?'�9���^��eV�.�y�r�?d�N["������P����4˥�韞��u���3B7h/
(�&*@{�y<5�Pd>V�ۖN�I������p'��kfX(R��P^�ϵ�?p�����z��=.q����uHm3��z�Fyu�r��ZNP˛
q�٣����&5�~����*7��"a������?��#��"�Y�pz�mg��$��Y�3���-Y�����mW��En/c͇5c�n�:���n��.O�Ң��Ђ��8:�L��0�^�<-�?��Yw�܈��"3X���hbEO��A2mav��S��l���kb�%�E*� h��Q��=K���*�D�8d��+SXk�GKf��&hܔ�����>fiӋ�u*i͘�nh1}�����G���rz�L�_;!�xZ����س�s0;|L���гΈ1�Fx\qg;�y�o�����O�e��~YF�`�׽�<����.5��~q$vFr�ܳ`����Kl��w�:w�WnzK�
���"#N�j{�͇�����k�'�%KT�2��!Ot���I�Ů[A�О10�� �R���/�p�ht�2�ԓ���U(�Y��B��+�Lc�% ��L[�9��� J���SFA:4`agK�]�Ѵ��tq��G�3�^�v�
�����9� {02�x���t.�"!:g��2�O��θ�)�ª.�p��g�r-����'�jn@g�T���vlJ ���������	!�I��-�W���ݠ�%��9�~&��C��%��?�#��u8�)�� 7����Mn��C"�Tp���
����B|�_���:8K=Y��S2�NM�Ow2�+3hN�4�v|�������
���h\�5�Ÿ��2�e�SO�%
5r<�T^��u��}��,�^��0o[/��_�}�X/�P4�݄C���j!C�g���Ɉ���V�S�^ f�	��⥣�C����7��b&�j���7�J�H������B.��?����cҪ���yך��
��%)]Jo��ջ6�4Z�� �q�C*Po��fY�Ĉ�^�e�0�#���A0���8��h�<,"N���A�{�x�1x\��ĩA�����k=wI�Z�����YNx�﯑/Đ������8�ޝ'b�򮮼6�d_c� ��N0�5j�F�j04<�����wzt)�"_z0IH�0n�։|��C��T����`C`r�n&)���`�&~˼��yޑ��z�"���S�U�@�!��(�\t���l�=�8bu��T�����Y?�,*^r���m���T��4���SM�PS@�"H/F������?Xj��E:?�1�Y�sg�z�ƵJ�u�9Cƃ�Cahw�'%��2*��ɯն���]�f�r�\��;������y,K����T��1?A���b��sa����P����D ����� ��������"��%S�u�row��	���{��A	�-�WM�}#��ۑ��5�`��,�y�W�%�:�.*Aã^��|v{U���%0����k2��f?,؟�Fp�f'�5lc����[�����`�߮���CE%�.M�,15����P+����j*�ף��Ӻn�0��.pC
�p���mw��� .'�"ˣ��+z4���h�a��� �|��(���k96M����Ȏ������g}��p~N5c��=�� ��r'ֿ���nQN�ͳA���K��r�R��ś�)I�b�:X��ΐ�yPe�~g�j�s��]6�^��rJ�9�HŹ�}#s8P�JҀ�I���Z{�ɤ��B�? Y�hB^�'s�1�Q�-yC� �s�G�nϩ�t�����{�g:����t�Q�~8����[`ӫ4�tw�n�v�����&�s��:g%���i��|;k��(X��f�� ���k��a��M�\q�d��m�sA�hqU�z�r�:�6�����l M5{��G��'�^'bzb�%��,UST�֗r��~�GZTi��M�Ck6��sU�,��.�<|�d��L��3�4�8pH�9��<n�|�$i�A���S?g7xR���Lf��bₛFO����	n l�&�Ɨ�����=0��լ�[B�_"�Tذ�������h.xk��%C��c��>�4*�H�]P���9Z�@�o�u��ҷ��xyڞ]��^`��X�[����wu����e*�I��@8x:�V�X���Gz��iP��+�9N���(����;���"�rj�B�?��췝-Fj��)�B/�i��c���N�6��4�D`���^g��J�o�\�=��NM�`����bI�CR`M��\��q!t��%s/�B�`����Ԟ��K�������ى���I%������;b���C�>Qg�yR�ǣ��o���	��Q����ʡH�7o(���}��(��օ�K#yCO2iǖ"���	��գ,ﶮ�j����b������S�Y�n����Wou����D�
7&L���%!��v#��^S��n��2�DǢ4��W*��Fq���!�L���vn�.�Ɵ���e:ѣ
6��EEԡ��!Kc,al�Z� 5堰�cH�DR6b߾�lb�Z�gv���7�ct�"� �i�PvEʆ�\�|~ �z��ڠ�Љ�l��;V�_}.H^�/�Y/33YO�[Ҩ��.V& O*�'X_�lD�
��u*Y���?h(�ϓ���<!1
�SID��p��3F�^f�G= 1�='	���є"6��W�,�|~W����*��f�"VM��fVb*XǮ���TL������2��\�1�ǰz�V���Xo|Yם^�/�ǂe�+S�z���ߞxbz�b{�db�N�Zg��b���a��`�u/qhuS�M0#�E��vV`�����?�Ѯ V����:
�.��2z���j�U�K{����!_κ�{P\�:Dy[�$��G�-�D�)�d�*x{(��:\�N�9�?(��i��h7&Z�_����f@~	��]�QB����0��p��٥�Z�W���T܂�,Ƅ�Su�����J>"}+

�xfT�گ�ـ���5��$�Zח��Y��y�p$UíH�^�wO���?�jw|;	����ڣ<Rӑ����o�l�)�}4k��~�L�e�a��:��衵ZCi��-��i�`���XTm�0'��M��]M!�V���V������'<|���������3;�0��W�,\��&�oyu_�JhMN�t��3�v䖺�����;q��6���x�$'�b�8'5����`֠���-�I��90~��-T��9�/�P�����������n� ����#�uf�^j��艥���VTJ����d�]9�t>�MU�������U�xnL���(M�듳������0?	<0H�<�Q��\@��[��SE2�(�t8a���~X�c/��cX}7���XNE�[�W�:SLF