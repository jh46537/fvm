��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�c����W�3��1��1���s�9�	ܝ)Ѯ�k=�nW���M��K��M0�%\[��r�ʕd�
P��;{I�z�K�y;���9���զ� ?1Թ��Յ��̜)���/0.o�m���Ɉ�;׃�"	С߯]b*�{�E�hc'�`��S�y���{��Sc+�eƲ���곦=,j�������?�ys��N�ߚ^E3 �W�`���<z�,0���:�&���&�v��CƏS,��˷� I�q�C�
@�n�PB��l�<��QJ��
)���Ry�)=��X�&?��O�6�rJ��XG�����S�����i�R;ĵ�1����<��`Ň�"#���?c��(1���J"�/U���vWcc�5�a	~w+���hW٫��\�1�/Sk\�Bw[d�e<�Z~`�㙇�A��;��G�� ��#���a#�X>�O��ܡ�Q�Dm%Қ�ak��05�L�*�{^�1���5�K��D2�ޡ��Pbn�4�0G�k�����l�0�=�����Km��=T��y��[�� ���i�I�^�v����S����!5"��*L�\�6�%��7���P5s� �u�c٪"ӻ'���?b�������Ic�w��܋O5��rKΈ�G��n�fS��\��~8/GQR�4Dbz`Ex[�	��`W�b���)���\�/��e��aBۗ�lԽ�#y}0C�+�}>Ҍ�Tr<��K�,T�~����D�g��Ҹ��]�@E}'�fuX"�2�1D�1�h�%�	��F>��*o�]�����fd���
vv��V&=�j��H�A�^�<Hf���!�����0�N�<�r����".N)���di��4tB(`��P���#��Z2>x�Ś+�S��eR�D�9'�8r�hmq�0gj�&�v��Fh�2���k^�6�i��QRsgH�	��m����)ָs}�j�2wt�AF�MW����k�m�4R����㍠��	�,rʢ�ή)�;�g�mNd����=���bM�ҿleϿ�G��U�l�Z{e���M���PY���*����>�@p��=-:.�$&Du�sብ�Dԍ��d�:O4����t��<O�V�ע���*�)�rmͩ��A*� 1��Ѩ&�Tn&�EHP?{�Hcj9V%,�C>Y��ޔ����8o_�bj��ù�pQ�8�?��P�U�r4�~*o�N۟ۦ��j��Hg'�N����WKb��	@ތ�/IX�v\��
H/�Q ���xl�t��w��Y&y���c�mKE.-\K	�~�rt�N���k� F�/��yN��kn��]h5a��O�*�3���_i)��k�p�P���z�eW��l��l�3�'�v���o(�T�s�����=(���(�=���}6��'O��Bl��U�K�F���V��0
'4��A;�*�x.֙��K˺`ʯ��Z�����p� �'?h�4j�[�t���q��a8}�I�|m����[��QM,���o�e���ò�E'��<~Va�Z?_oP�rP(D	΃�bS�=d����9%�"]��4*��c�ғ�q��ˀE������wE���P2����ҕ|UC����!�e��N�d������ !nјj�l ]W�{B+C'��x���h���Egp�ن]@��C<�����������Vʜ�_wFUA�d�"mG��鈏��ږ�Շ����
�j7zr����V
H]�d���(�ex��?��FkȲ*ߔ(����\����=:rߖe���Xb:m��ɡ;�@g���莒��F��8��G�Ӎ�޷s(��\=.2���q
��t�F?a9�%��_�PwJwLi͸|�y	wZ>���9:E��4����6����?��O?�M�k�Y���όV�'-Dk����U���{>�D+t� ���,��o�F�S��K�n��e)�_wƜ�"������Ւn���Ҏ0t���&7Q��� <�A�cx=	%��)�"~�ud���h~�豹WK��O�q Vԁb%�7+�4�O��ZU$�5[,
��u@ޞt��e�� ����,Rhb�_��ﱩ_*Fj��Ǿ^�p�y�u!��T�Ѳx��2×�7�Q Y�b�' �JC���X
3�?�{b��VIr,�K�\��T�� ѱ�G�59��1䝃Ol4�����ː.�,��E�/ԫ��;���jA���2�T��93$�GOǺ�W㰜���rw�-_�>61)e�rT�D��]�*X"���o����i�	�����tk A�TB5c�pS��D��`��v�\8�]����H�-��TN�H� G�T�@���*���^��2m&�f�=`��w5EG��ds�T�{%�>�	SG���'�̀�
*���x�G%�^Z�QN�Q�����ZI��AS�y��n�� ��:�'&�G�C�m�Nz^��|��h��N ?�^0M*B���Ё��Q�!8e�0y �K�ȪP�k��N�Tw�it{+b�3|����uR�ykوW0a��54hZ9��@h�O���Ur�^R�����u����7��a#<:E�6un�8qa�"P��T�`2#ً�:���E>�������tn7����{ꎄ ^v�["�]��T���0��;)�ɼW0У[�Ry���.�����eL�P}�2����ʪ��Rʘ%&�͙�㝚&V_ݏ;�d�Mm9Ǹ���v,E6��:�q���!d���Y���R�����wg+g�ٯ9zD�k���6Jd�.����>�� ��cy�D���չwv�2�l��YB��.�Z���qJ��;:T�&c�HGr<��RH�L�oPqP>��&+�&��#���=��ò����[bPC!�:c���c��	Q����܀�Mm�ZͲ!�A���z\�<c���b���Y���.oUrSԭ�� ���-pʝo�
�@]s�h|n%Őt�xd�l��ܿ=Qv�N-�rT��n�Ya�"�T�F]0^�エ~��>�:�T/Ĥ5��?���j���$4U�����H�l�*����ݠh�|��?:���h�th��R
1DRE���'m?�[I�"��ѣ�"�+�=j�?��X��ԛ��{��A��n��_Nևn�ķ�hi�4�����[��-��߇��mȞ���(i�(�;/��>�����������(�O}T����>9�~lT�$�o�|��7z��ePި�%�՚Ɓ��}�qgWԤu�b�2!��;�iX�q�K%��(F��1OY\>[�(Z%�������}Dr ���E+�'Ho��h�9w��6��گ�	���/���+���Y������*���Z����rV�J�ķJ4����V��e1�ط��۪��/��`��=2�<����"C�j G�ς�������^��;�=9q��p�"�cfwA@����d�2����A��9����_���a���+9a�^3�VI3,5����2fN�����k�����1�Z4�^�c�j�@�+*9�>���O�^)Q�L����MH�\���^������ .��3�1{#�����K��*��5�G����~O� ��4幵��
�$ �n�)�|��Ã�B/����8�͵�]�9j&��t�[�8S�h$ŒF3�h�̳�$�'T����� ��9o�X>149��͖n+� �4�_"�-ƛ�qp�d׉��m�bf����uag��\+���Vb��M�s_]�A�3�������!^������c-��{�����$����W��m��9�}耤9o��}��fsdg�7�Q$X� �Y o>��Y����B���K�#�ޏ�,8[�YV�C�J�W	C�4��_�.=��(�&�۫�j$�*���/M�B1D�*Ծ�3j���t�]�����8χ��o /��>	5(�`E��R�����R�ڜ�OV�2� �Q��)�]��<��oSO�wr�_-;)�CsC��R�ϵ\��Y��u1J\���B2vX@�h��5�?^�Ѹ1�yv%An�XU�ou[{tW�u�5tc%E��z��O^qm"pX�%������/e��~2A?�P�%n7����P&��
yب�R�q;/�\Mז�0�xZ�`�Б��h�a���a�IB]"��s5��.Y��L��.rBӭ)����Εjk��B�6|�Jw�J�x���P�8��8q�К�e�|)b�Vzm<�'Q@��E	�= D��o�J8�=�`�5�3g^jq�d;������aS�-��u�@�E��~�z@�����t�T�
/솏O�d�
��2�%Ƕ�c�4.=�h���&�mv�����y��S֪�+��Mat��ߟ����@�D )�?zw�k�@�z�Y�I��	b ��7�gn��HAN�[�th��4Á$Q��E!Ed`��^�j���9�p0���8�MfK��Ϡ`��E|�֪�^�G]y^�N��K���]�2l߶�N��O�6���^��wV�J1ʌɺ^���S�]~�Z� ���ώ�~����7hz�r��	�%J���Qm�#7�q JB9��h�� O^z�U�����9�*U���5 H)�L������A�
Z�j�hC02���G\z$�U"�k�u�U�;��C�`�t֝_�$�  lwb#��׈�i"<��%!�"�����R@�����2��.iY�X����ͱxl�.�K����.�ɛP��A6�΢z<��<�'jK'7m\k֖a�"���U
�2��!���˧]Ƽ'��K�L��X{���\+i�9�`I�����GI�����d���8��#_�?*�m�y	����j�H�!��W��l+��vb������U�)}��:�h�Ůi.�N_gD��Y��VXz���M��C������rv7�6��X� ��D����%
'X!���'?�(��8ʴ��/Z����G3(�L5	4i�����WM�|�j��c��Am�?�C����YC�.GQx��������ȕPEK�^��4��|~oΛnx�� �#=�CZ\�ʾ���a8I�<�Sժ�ë�E�q��6E��
�n/ݤ]��J ���|opj��|�V@(��7�|�6��H(��_�t����6��2�)�e��i��PzAQ��Q��&��3Y��#��.���K���L��(³�Q	h�y�7���J��w����Ʊ�B`Ht����=X��0y��)�����,�;4xWhr�¤0-�ZC�.�UGX�A����r��A�Kk�&�M²���;�J��U�h���� �
�[�s���e���˟Է�Q���!��۠11&�Xc����L��1�zm��o��'pP�t�sa�*N���81��Yk!9��7\����U�YU��%��R)BI���/U�Z�2	�\B��flq,��G�.�P���5[��	`ՌbӸ����1FNjmg:���"�X%��n