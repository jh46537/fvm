��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��x ƴ �A­,��z�FŕV~��֪������a����4��]�/�7߽�ʈvr���#�����X�`C�.�eQ��M��w9O�@�� �kP8ۋ�ǰ�]_g6����9s���ikz=�`2�c�F�O�@	��Ϟ�Eo;Q����*����7��}l���I�	�Q~�N�ڵ�V⯷@��z"3/�.l\�������-$�����_-���1�oR��uZ�v��ܲ�/��zT�#�\m�ͣ��%�~Q@"�9!~"����~� 54�_���黼2y��2J�`'ԧ�h��i� �M�4��N'�g^0+vnu�����vk�M�;b��\H8�Y�Q����<z܇������ o}e�mA㟗��� T,�Ȁ�3ZM1L�"kvס8u,�2Ձ��H�������/���yqP(��[�) �UcF���4�ǟ��d��P4��4���a:'S��E�5����^P�Qi����)��Af4#�R$�O��~T��%JMN������_���ԡ����̖�?9��`���A��
���Da�9���G|��;m�`
������ҿ��*�P��0�JT�T�HL�clN߇:R�4!Bfj<B�n�D$A���}��% ��F �zY[�B��������wL\�B��h��PTE|0PU_!}c�����5����9�w_���b�f��bn����U���Â�,��RȂ��m�3��QY)["RB�^P>��*����ܑ��(��#�2N���i2o���P�_�ơ	K[���4�d���+�6,K	�DA��p��-��ou�W:~�o����
5��	����o��8ȩ�`C�8K������#����R�٤�� �����K��ѓ��`��b����@����
6.6�U#F\��|���Q���)��N#�}�I��x�U7�����uʑń)�{��{�B��j>�xv��f��\���SO�SX�����E:�@!T�ʐi1���M���������_N:��z�U��d}�:?D�C�\��5�L[v_��y�M����V�"�[%,d�{��C�>��l�J���2 �V��rz�ؒ#��ե;��<��<M�,��|g����~\$^��[���}�"�_4e��Ä� �Q���d��C��<��6:P���њ�(B=�[*����0c��P�T���.`	��n*�5/��e�����r�T���� �M02�T��$��k�$`Ο�l9aa���fG�_�ʳ�	�.N�N����P7_Ht4��y �'4dK�(��~��Y�QqG������Z w�8)�
'[����Ǧ��_4�Fxx�J[�<�Է���x҈s
/|����O����:Xe�5�67L�PJIk���dV-d�J��&Jv*{���- ���M��G���3\�o!<_^ �LT���z�{aab,#��$��v5����㈅sU�:�����S�|ۍ�f���L�OM�R'�~JL�����������q�%�>���A�0� Că-�=w[N�3��-jn�%ˋ��Hv�K5��@�����l�VuM{���@�͠�	��Uu0���$.Q��le�-!ol	3L6�e�D���?��;�TRNv{!\��Jȶ5;kp��m���Y�O���M�CV�&`�]��xhO��Eᓩ��j���� �NI��^y��	�����3�����F�LR���"�>ɀp����#� �d�~P�?��L��u#���~nNI�=F���u5�� ����j��q@���!��):�-�L�P-L�Yj@k���4	G��`ov�C�Z��TDe
NK���fx�z��̛��wBt-^����Wu�ǒ4�F	X-\0������/vY����7�\WG��?}n�2TFj�7`��w���\4j�by>�ڙ�˛9L�eu}O�,¤���"Q�-q(�}���%:�/�>�����h���3.�#�4iJ� It�;ݯ�64��˛i�����:��,���݈rr��d��l�E�hխ�6���-�]�O���ٟ6�򀵵��^,�爏|Fc� ��	��7�1�ߤ\�4����ț���ֺC�D�]�t���R��Q"��TX�%��7O�m� �Ϭɷ3���ת�7uZa�&�3����j|�4�l�H�KY���y3llz��<�>���{�;�����+D�/�NPC=��3( ���<zzV���CuNQ���������@�
*�}���֊�i<�����lR����Q�.�؊�����Y��R[jA��&���Ƞs�h I�C���VRk�����ӈĄ��3��q����v f'�d����N�0Gӄe��T�:0@�%�y.�b��+s�v�o��W�}ڹ���<'����[m��]Y�E�`Ι�K(�u,���5�ӽm�Ą��.�Yi  Z|q{���UՍ������fL�(R[��"�`ӛB���6�O��̛K�s鵎RD����@4*k΃��XX  �o��z{��]�#>~6'F�V/��h�4��֔�(�vC��ٳ\�B~���#�F>X�ez�R���UNE����o Y<-�G@�O�^�\γ�3�� h�F�~�	���Y�iD���}�+�M��"qM�#"e�7?N�蛾�ia���Bv�.c�|6�U�I�:�i�wp՞b�r�5��������;��)!%�6+$�|�`��%%,(� `)��z�� �!��1]>�x��~ ���-1��$�T��«�u�-ƙ�΀�5�S�r�Ka��W&Ј�.ڧ�j�Nd�+�cE����7x���=�ٰ+92�]ZH=ʊLu�+Npuz�I��ߝ�Xj�x�G3؆�5��=
Pg���/?~3�nWŹ~e�G$%F��_�QA����#���c�kO�ʹ�����/��k��䖠�{���/Wӫg���H�r�ߨ�4��9��f&TA�[��I���H�bTz8� �,Hަ�ꚭ
E�$���$�ć{�Z�c��kTĄ�j$�&�d=K�޷��Z �����[$��_����(��{箴0�A<*i��-ƋRqMri R�ʀ��ϐEc1��,c��!l�{��#�s�+VQ%�]a�M�$� ^2* ���=)=x�w5k6�l�X}��(�ƇV�F����?=�B*�%�7��h�oj�������x��V��=?���e
a�M_��9���A�I�z(I��O��׿�~��,�*)�#��嚦�}Z]���H�e/�V�G��9:�Rm ��F�M�y�$u4�O��c��a5x����,� /`I��]Jy�����R�Q�=�RdTS�M9P1 �F&�Ǎ��Q��6�����ME�0�X��m�In�*yw�o�y���o	2d��za.K������_��|�i�Is0�I�zm�c�`T$Ex��*�
��Y�1�<9�;� &��v��m��I���D���"�ۗ�j�$o�u�-��8�ʏ��qh����AZ�F �a�H5~L��*Ћ�˛&���G��qQ���C����Y\�n*c�=)hh�I�j�S����Nh�|M��W˩�/�"υ��^1��P�g��q)���+w߻:sܐU/�D�t�)��Gs��b���|o��f
�S)%r��O�-	���g�0LY�a\��y߄���N�ń��\��=x!�b��i4�~�ó���#Oz���ж	j[�����W0��*�I2�����u2+4����'}�)�Z�f��L�(�t�a�H�����f�G�� �C�~�Z�O�-[��I�(��Ę�Ǣhb���K7�k����Ϙ.R��v�;J"��6�P�O��&�[�8�x9`�f�7�o�á���[�+ts�BC�i������ⱸ��q]HÃ�.�v���?��sۊ�v��v,*�1�L��
'w�q�
���� �2��H����,Rg�+y�k��[�fp�v����A?�wu�"m��~�)(�0�J�tZ{�s����,PԚ��-66[|���)�UK�78�ٟ�Vq���_O��Ey������~1�6���l�7�P	G՞�;Y�8������|j0�wo'�4У���݄Rv�MU��|d�q�0�^��<[�MS��7`�F�s]�7x&�χ��XƘ؁��ܵ�R˦�#��	������\9��"�c|eS�C�.�/RŤ{�c*a���tB]8��ϕZ,֘����K�E�:�1S�ɍ�D%�;��]��x!��!:��?��UZ*�a
�Yh%�2�>�x�� ���|q7�npߤXX��P�݉a�W�����I{ԅ̞^x�4YR�fă;v���a	&+��N*};�v
_~��z9lJ����qs��gG�|óK�;T���2c~� V:ߒ2����QO�T*=��A��a�#��LN�Z�Qn}
�k�lEo��������%��jԡ�����dh���FF����Z���.� 8���H�U�I�(]���c�)6��e��yT�9�J*��vH�K��m'Q����wb��}�8��9�:�q�Xu�:E*��06���m7P�}ڒk���:k�<W������}<j9��˪�2H����n���^F�6C��������G���-vsHXGZH&�^��r$�ȹ�9%��R�Y>j�N`�֯���t/�T���!���D���t�k�;�SP�++�6�,�Z�K8�n��ŘJ�a��Y�2�d�(�s
_�P3�'�ۻ��e;�9E�\:!>Pg��_���%K��Jn���(bU��;�Hx�K:oj()���mK��H%!2 �3I(��~�Bz����o�aѐ:��G�w\�LQ)nPd�`M��J|7��I5����8|���_�4m���*��Y�"�#6	�PT�.����б��/8�0�p�a��Yve�ǃ�<�(| ђ���j���ҡ"�(͋	ʢ	f����UO}s4�`_{�%�d�	,�"��6��vP�7p�.:h �w�Qc�_*�(;�b~����d���`�14�s��\%�Q"���B�`�y��
%4n0�W��n�n��kjϟA�����wf�=Cb�7�#�g�K�l���o���F?m&��J�M�|�<���ǿDL�!��CB�q���>��<��A�yl��S+ Fo�V8�Ih�u^᧴��U&��~3�>7����b�A����B{�{u�O4��:DU��k��&��?h���CR�<�+�0��AB�k�_+����:`���=�.Q ��4��lk ry!�f�T��$�߲�c}#s��	��k���&��}Piv���f�V���w�F�1|�����δ�&@ƷV�B����,�>_�cb��>d����D��o���%yxB�>8�)?�����C�.�<���d��J��t��u�}�n�H���#�h�U�I�,,H�;����Ո��ߜb�;I�J]>!p5+�z�
[�YwRZaMR��&^Ԅ�F�������Ϸ����-� �S��5Y���8��3�+H[h2�hN�2{?�}_�Zmi%NF�J�T\GR;�f����ع幬r*�e��]��t�3�OM�:�̈���$�:��Waר��֢�p%����e��+\��D�mfO��樖>�����I��-Ё��-�+�2Z��`�u�3J3������k�:*el���ˋȇB���l<����V�5�m�~��&v"�z	٠G�/*;M�u�)M�oxLF��k
fy��
o�/{jJp�qX׮M؅w,7.]�,��[��+
xI�	���i�]NRhs��K����e�n@�3�zn&x�N���"��ur�w�[�K�i��	`�H��b1x\3Y
P�͌��.{��XZ(�����n�J���W���8�F���2x��	�2C��EW"B���k
N�K��s�Q�=����<p��u#HV����(�.��2���Xcر��8��>:������Ё��lE_,$6��G�ow�-R5�Νj���ƓD�j%S]�?�=�/�a7�w����-��U'q� �U�͘�1a���}x'��~	j�R���i9D����r|\��-N`�m$<��;��%N"��gcyK�އ��s�?�J���}�\�]
� ����d	~�G��B�Hl��SکDdSS�����)�����c�-��		5��H���S�^vp�/��nw�^�?�;�d�t�߀���c#��vf_,�㑡�w�R��pVJ~����Z���^?CN'z%��ǁ+A�#�I�#"�����66���Y�t�ж⮀�l�d�[�[�x�j{�ϝ�_����үЋj�I(����fx�=�� �����E-�\��c�Υ�֟��H��u�l�^~���r���U��,��_(�B����X�w�/mø�`�dJ��^�!e�S6$<Zd�3`/���:"g�O�(X&/��"�8��gB���������%h`��k>�1
���A�s������*j�1�t@ߢ֩���JRnz�*�d>4o�!B[���+�������s�v�Æ3E��j'E*��O�Y����hk����Q-�3a
91�Ʋ�ò�'��w�	���Phw���tWb{�hh\?a��>]��r�1���Y�e�<[A���I�i*�f�<�H�zoj����,���5uWF<���n�=��q4@EJ��%.Ԝ�%w�^�1&g��!���%P/4�Q=��.�DY!d�(�����y�(-����ݩ&��i���9�hі��f�n"���x_��������J͈+&/4��'��|�R�� AY�|��^a����� {�q�$���=̩�����g@r)ӽ�e�{����xIؐx�������|����;��C�]�+�aOkv��%�Bz��˥�W	�~[C���N*��j=�������48�p��%Ʌf���ߗ����Yvۢ�����������"�2'j���,0_�w�����h�-��/��.��{x����Hd&S�� ��P@����ӿ{�ˁ�LvK�B��[�N7�b�l��%��l�Բ�f��~{K�}���.`��.JƉ��O�=a��|	���p��w��R���5jZ��Z�S)[����b�ZA���_���ȕCU���e��vZ�l���ހW�E1���Ӯ1'r����R��ev{R�\�R������^{�J���@�ŗ�L�%�V�֚ ܚ�\!�=��ߤ{)o�<\��C���Z�%a�dS�ɡ�N
װu)F�d����(1-u�������	W�-P˗��������
6�P�*z���_�]��)�!	��bE���1.C��NTk:u=C��qT�/v����=D6�J����uI� �~� dm��f��}����7p�9w�Έ{��	@�X��9�`�xrN�@��}�+�e#X����@2�O��A������q}����YŴ��~���|9|tN�6_��l�z�}*-��E��Y�C`Q�4�:� ���A`x��0����<c��$�JW�Θ�J��XO�E����LG+'��\����d��]����B���$�����<aءR1��D@�(3��)��J�lP����o�\>{�fE#I��$��{�^��n�.��4�4x{�&����Qʝ���#�|}B��'l|����8/P���EA����ƕ��e�|����Юt�֞�o���&9�~�[m�;�&~�(����1�e�@yy,x�Ш�_wi��kZ�UlX�����/�HQ��P+�W<�GAw�u���- a�At�Z��R8�>V]�x�c}��?[C��N���B�H#����tc��6Τ��ګ,5���Jp�����El��X��>(�2�����
���K\!�ۣ�p9̀���+>p��r��ڭ��`�fD��3_��f���7��yy�v��ō�!���ޡ�1K\ݷ_��\ZvӀ�4�ե�*�������{ފ�ð�U�߮���Rә�G�S1�Sࡧ]ذ�飌�Q�o6Y�7��<po&��
3���μ+���9jU��Ԟ��D�,Ƥ�tk�GH����I�)��f5
lu [z��f�|T91�=��:Wy��)�]���K���|5���64�~�Vb�\5p\e����b�{%��"��vd=P;|zI^�=S������ܑ�1
��渤]��2�Yr0����0�8�Ard!�4AR\���I���qIy���ǰy�������{�o��1�r]x�����fK�*{��3/��P����B�zz�p���/�Kg�8��-=�M	��=�z/��M�$��2KXދ6����<KAS����k\����b��h�b�wpe�^�� W\�����C��E������7j*H���٬�V���j�f��]1�[�j�A��J�B�W��v�8�υ\��!��6�|�b�(	�\fD���1��N��oaM�c�옚��_��E\�'J�O��ꗅ�e��>f�8�:�x�.���İ��^�b�o[��5���g�W�i���^	��9��6FX���|���S�
���P���s7;_%��%��X��.�;#�m"�I���!�FN�U���ʋ���'k�J��܀PRG�V��6��yLd�.�E�{��1�h6>���ʁ��J����}�uyS������t6��zWS=���z�+�G.D;wK%�%��ׂ��#&�0��se:DV��d��S״�Z�)Z��2�;�K��8��} dL���(�Y��[/��V0�>{r�u�D�/�u�Q�N��n������C��|g��.;`����P�����c�+)��^�ܿa'�a!�g��5�눀'����~ٺeޱ�����<}�Bjt����(��Փ�]��|r_e�6X�9"x���R�n�T�D��v
��a+�#i��]0��\�[�����!�0�a?��7��Q׉V̡��Pn���fJ��OO����IXp��>i�������("X�#%I�*O�F����c�i��
��C�nID��D�B�&t�2��������f^�|e���і�+2�j)����4~�`��;t��@���</��}+_/�Ԉ��rv�9���nבQ�w�%����A����hj�����f�����_`��.	M��u_F!�k��)\��^.s�����z"��\��%\Ɇ�F����/%�8�o�6�-�`�!7(�x|tsx=2(/#���K@�`���,����v�Dɋ�����V/�鐛���eԱ���O
I��`��@�V`\W�&����<,�(C�o^}�W����Q������k��ժ��K�z:��n�p9d@��)�h>"!�%m�+�xv�cr��|�K�U7�:H_�/7'�O5����I�'Ka�������V&\Ai���w����t��4_�`Qk��u�H+'PP�Y�yƞ�m�����'�̇孥�F��9QՂ�v�����1�E�%���"�a"l���-������&��&;F��'!���w��P��l}8V��`p���>މ��
�J���;e��r���g<��Q����o><0�ᖟF�}/J�";���FK��e-<"v��ʍL*Q`t�ܞ����;�c;�,q�eh� ��,���y�^\|�E�K����Y,��p9�0�� 4� ��M	�+P�1�_Eѽ��?��?��A��<!�8T���o�g�>a�I-��צ�6�/'�mt�8E%4��L����s�2�1��������E{��e�y�[m�b8L�i�P�zm��"����8i#�Z�Z�P����DC�T�P�sdt���ی-����p��Dr��ɶ3͑mg~#6Ŭ�øF�PI��g�u�X6|�B��`�7�F��4��ɼ�`��?-
o�Ya�RI��:݅?C�
��&F-Sߺ�ia߸�ð�׆)�� H��%���y��7�] 3�(�N1++��R����;�	��} �E�{���䅑ܱ���������)\2I2���3(�
���� ݐ��M�*�&�����x��avϬW7�]�<��s��U�\Jx������B4����S� �Ӷ�g���Ղ���V�t��Wqh������D@�}%���ʼ ]L����C|qQ�Zw��y��ф����{�Qv�U���-3O\Gg��J��E���qq���Y��ҝ��II`�(��p��� {O��X�&����8���"ۛZ.D�V��IE� ���
&����&-s��d�R9�C�
�K�&���h�5�y"�>���/;��϶_�n�
��3��\e�(�g���G��B��z�[�!L�8�~t�Y%�""�#L�3^���2�?���U#����XHDm��Nu��&���՛��a��َ�`U��X�'Lx��ء��!-mR4A~�%^;���}M���&��A�]�f9$�RN��!M ?Nv��#;j6���Y�A��{u����@��g������q�;(?jn�!��
-�q��]�+F��/�#G���볽��5�v�}�>U�jg���"����9�%n�a������O@���Nm�E�Y�ꌠ�c�eD���OZ���H�"��3���͍V������M?1�QY���]'C�!y4}rs� �st|(Ir��"*�y�3b�'���D�����VR�,;����k0��N�|�:�����蜗n��r�03�>o�'��7�e�˞	�$�q���N��ߜjSn��0G��� �z��5 e��wE� ����1X@�w��Qrہ�'�'ꙫL�XO8%'��#��'�]'0V*�L�u�#�UB͚�����}�,�]  �J���Y�'��t�q:p�?�z�9.]:���dO��l��c[s&W�BӀ�i���Y,����v� ��ЊZ��'��YI�xx�
���(g�>�B7�BJ�o2m����`�0��:�~��ۀ�ɠ��:��ۘs��d�34���ڸ�����N�͉8�P.��E�����e��X�[c>�Y��L��ּ�o,�s3��@�kI#D7��I��{҉��L.E/	%�Td2���"�����?T�C���+�������&���pr���=��O�Pk�Z�ں�2��m�A%����]$���ɸ��+����*`u�FSrb���#�ݘ�\�F{�$�ݺ��������n�j��&l:��|�j��!����RDN���H��1��IIx�p�C�����^T뇐�Լ@rS{?��ڈJ��e����O��'�(np������7z{����� ���MqB��FlR���CTF��K%.z��O6mJ��;'�fE��n&N��m3+N1�q�
Y���$&
��
1K��%�Ln&!kK��k^/��[~TA4'�$r�[�]��D�� |IY�ʱ�b,��6�R\���c:�/�t�8�[L��7��:�2���7ŕ~�y�؎�J�F+�R���ܧ���@ɖ;!��������T�2�s)��r*�ӡ�h-�<�4H
4"���cS�+nS��h>�טsy-�^*ٍ$��XH�}�t��n�'Ùc�I}�xOd��h���Z�v��$�����\�u*��8�8kW�g�����Ӡ_5qG
_weXki�a�:˅�bC��C0�᏾��݋A#����?��!J#�r�n(紛ԚN�Fn���׺��4�rzC3l)[��:g�,_b������'Y�m]BЅT�M�����R�����U[+2�{E�ZX/�O�su�<�я��wBs���ۀ\S����J�Hn�ڹ!WG�4$O/L_��P;�+�+�,i�� ��y���/'�~��T��=������9���"=�(˵��e��
B��R�%��ѳH�!Qn�k���Q��\W�Ѳt��U!p�s���3XNO �dĲ���E-�1ʸ8�K�FV���1TPŨ��Stغ�-:@O��|32f���q�+��9�*GU��"�T�x�d��q�9X���f(y�7:����b9A�p�,m���E�5��_7 a��6ү��:s��`��e�R����T����}��������HY�#>#u�]ϑh��_��9�N�@���:���a6IYնb�P"d���W$��LY+R���
�`i��Q���>�Rs)��Mu��o�s��H��pQD5���@k�S�A���<%�*����S#J畕(�nl�K�j��Y}�����xh��(J��.1�tFEP��N�9��)�p��P�����qQ���H���˫���Z���N��p��?�)������a���لWP�V!���S�SXa��J�,=�?e>a�֑�o$Z)H1�%�=?�W2�QY�R�ޫu��i��{����W��9�������mϘ�g���?d��6U������
5���3�"����Xek<���	2����W`��=�؇��<o����@�Vˮ��*_��M���H�$��Q�~>�;�w�r\DĻd���5l��ߩ��v��/ݕ�f����2(UoYF�`K"h�j�c�ɫ"�;p �/A���L����1q�g�Qo�j�V)��n�=�7��Kj���X��������77���������D���+C]��B�>&542|O%��/!1�">zi�Ya{��ǌ�~��-|$��v_�'l����stQS�4e�j���a�|J$�dr�N�$��}ua*�?���r\�V(�)LА�45�?*ȿH�;���tf�k&X�u���![�K^;�`f���T��HF:�RY���*����'Ћ��f�
��D,�B!��$�������|�8�[��\�K/s�h8��^��Y���G��ѻ,>ZT�]�L���[ˤ�w?k�k�� ��һ��(y��H�2��՗s��e��U&
����C\�S7}V�T�l���u����s%N�z��|fG>�Ѭڥƞb;��t���g�lH��j=�ѢP-�"� Lc70�Y��n猅l��Ot�V\ϲs��16ͽD�v��q��
N���޼sWAn����g�w42�,u�βi@���b��b�� =��W����&����=�nAtSO����I��p@N_>pȻ
�Q���ꥩ:Z�4T��N�3ك,7p�#(�%O.�ټ_�0��4\Aq� kʛ���s-H���<P��!D�OF�w��P�t'�F���_ф�C�0��k� �M6���9���1 :U�7�p���_�ֆv,W�Ǐg��Xz��3SP|;�,��bXQ[Մg����%�1��.�b�/���¬�I�'s��E�#&��c��퍚�n�%�#ԽI����0j�����@\W��t��P�n��&�������R��V�`4��	��GTP\�|��G�mV|!�vpc)�@)8#Yy蘣�R���&�9LY4�nv=S�D�n�5y������Z��Ե^�o���4�ݍqު���q��•
���E��Q��$�mI�]G�{���BL��_�V��4s�>wT��o�����Ou�4�@[��t�Of�[\� �k���oQN	*H��|$��QG�R��d��<烪�Ĕ<�'�Ǆ��'h�@0S͈�6?M�|?��J3�fh<��
Jq��0�����K�E�j��\�щ�°�P�K�#�nC�Oms{ޝ�tjԸjb�_�t��,wr��0��i�	x����7_�b�~��Ku!�*<pE�B=p�*!��l��nT�9�NqJ�w�s`܌�bq��@�o9}��f<a��P�Ӄ�(o��h~�3�F�FsI�T��o4 ��qP_J��v_c��I�eN��JUT�Bc�{�D��V�[��J"��(u�=�L��K<�����O��~\��4��_�C����M	B�����Fo���XG�kPV,=��X�]r�����My�il�0�}�S�q*�f;��{��|n�K������G.�[�^2��\)ed�����DÚWL�,��|�x�8�I���J�
��i["#�ڋ?�rְ�/��v(���XQ������7�"25O2���^ q�e���
��~����0��{�u��1壶f�2���r�c���p�<�&����M�ѱ�<V���2�z��gv_��Y���/LD�;�ŝΌ��h?IU:j]q߉v6�ﵺj�L[D��LM�2\�D*g²�9Kn��-%0	~���~�9x+��Z��ò�j�,pcG�Y<��؂�UM��[�5���n���d��T���k��Z>������4��|M
����8��H_��óF���)_. +*O����°��A�4�WU�שCifjv�cB*�,�0PR[̹�-p;t�*����A�̀U�v�q�I�\��)~5�� ����aB��Ԏ�ٻ�fǾ9�͢����8�GI`	I#�(�σd�!�M��6�7#�[�RQ�;��q|JΪ��U�ـ�G��ƌ'w�ҋ��C�	�w�ͣ�*+�֚7��1�P�=I��W�Ę�k��]��\͋1���m�U��V;����;�2���ݻ�X����c�/x���$�[ϱ%��u.���/.���/->sݠ·9X9�TϪ�
�kua��=o�.�K�_�ss89�c����>��&"D�8�۞��Vd@���λl��Q��ns��!�O�#o�$�v�7��x�y�{���_��.��[�k=�!�kE�f���K��c��G�rq�U53pf��哣d\�s�d�"g��\��@yX1��u�V�07i�Y2���I���-n/N�Jˆ`Ɯf����(�M�%�<�H�H��JI���ɜt��>-��6��P��Lp�Y�WڐI�[�g���Z����`��+�����i�xPOc�=��pg�&���֪���� rX��!%Nx+�,^d,�����0$��1����M�	�}��^�?�u�N���2=p͂�t]œ��dOLKp�RO�V9�!�"}q���t"��Ū�54k�:�$��9�Ŋf�e�*%��}���$4��3=��w
9�.yfo�U9��4.�
m�Yѱ�?��?x�6��D=j.���d+P^)�@d����p�y.F�L�wUˉ�'`d�svG�m��5?��Y�2Ae���Z�[������ȫ�S&�{B��$A��v��d�n���2J�|�������ś�ѳ�,�#���p_QW��l�6�|������F����^��5�@ƛ���BN> ���D� ŒS�(Ѝ��%@�����P�`� %]���q�"����+�X*�\!w�mvum�o��di���33�ݣ
�Y1"�7����U^:r����>�]��t�[1��n�i�u.LF;�`�|8�����i����u�!�D�`��Q����%����`X*]H6iNk�II[�����fSW�~B��� ��~��T�a��v�vU�����ƪn�0�]�B�PYy����0ԋ_'S���!r��2v}}*?��w���1C~r]A�/���yV����/gM��ԍ}���ZK��nî���:~�4�c���:G�����mu�s��UwH�om���`1x��Ѹ���#��y@#Bj.!1�����j��.��=մc*Wg��#~�.{XӵH`���Fha�XA�rK}ADU�s��QPW�'%N(�ԼPǚ����bM�J {��k�r��d(�j&��ů��u�j�ֹ�c@U��2��3
=̍�0�����W3�����n.b���s�B����^��l��\�p�ՀE��ь�h�P�"��>3�Z_��N(�r�+Ї��"39w�2#�۩v�j�zwN�K��-C#�c��n�>�4�Q�}�
@�h�8�Oj�1�ĹM��L���i��/6��ʫMm���0y���|�=��� ������	��.� l��3�@7�7��r)ú�=n����(E������U��'�+�蚃� �y�t���y��<��Qu36�V�?_1I�¸���6p��I�P���na��To빫K��%B�wγ_\���ߞ�n>y���p}��97Q�8��NV��G�(�[����A6�^�����2xa�Ϙn�E{j�"?}G7KL�X�`Pi��5�D� 9����} u`����VP�7Vq����}�-)6�r:���{����6y�X�vdyl
��.	������J��z�O$�1 2�ifj�n�����dqХ��b��K���b�{�FO��|����@���B��f\h�;~W9q%�f���U?/_�l�L����a>����s�W���?"ʍ�Y��0(��4`�VGB�H���̸������0��ڸ���N�Q�q�H��CYG�g5'�z��f�M],�����v|[��W�J���bd�w���"Q�5��}jFIfkD��u.v��
R�*B2ji�cZ�8q�C�Tj��M�H[ڴ�h��˶*�k���L2�ei�aPL���7Y;~W�݅4�������d��	�֖;��
����l���� �V�f`{��'�e�.-��]���G.`�J�X�:��Zב�y�-������+�?�+�,�xG��a��\�CEi/���JԴ�J�[o��$m6�o0n#��Q6�-�8܃��-F�N�\�a��M�V@岳n�F�o�9`!֪�O�;_ ��^���d[��	���^���t$Y�L(~���g� ��>�'�刮�dE�P�8|�L���ʗYP�������gRm8�������h[h�2mM`t��}�R0���R؍��]ݴ��ޠL�^A,ox�bCs�k)��u�B��4����e+��=�j1N��)�BT�!�F�)oMo߱��s%�a1��Dz�$�L�V}�Ad<:���?�=D6���0ﭏ�<����H���q��9�PeOt9�Ä����Zzt�q�D�e�]0��y̘�AC���6��[o�Y�w�qeꓸ~Kw�,��d��b�I��C���Jn��q�J������G�q�'�0F��Ô��z-vsH��.�(�g.�������c��v>��������O���dM׆��A���T&�s�M�܉�^�͑'
����Y��	~!܄�J�@��S�Ed���mF͚��4�g�����d������V��v;,��Q;X��I��8�#�<�Z�o@̕R�,Y������}�+��|�S�'��M�Y��c�f��F<�:�u^���W&�~��:"�3�a��u������3�=��D���񁪏~#�RnC�6bQڡ�y��Va�5�+�_��!q�~P����uP�!�S������8OyR�Q}Uۭ����0Z	|���Ci4�s����w<�g�q�_�)�C�*Ԝ�i"D�~d�|=k�%�Ph�����H'7���[{�� {/��O��`dG"H���D�=�c ZP	�Է�Ĉ��Lz��6�|��J=�P�%E��w��W���g�3�h��18L�����4���U�s3;o�ۊ���z7]��mUE����3c#�X��z��UkfZ}�@ʆ�\�_(��f�r�ۡ�ry��/�D&��Ѭ���#�E���I�\b�9O��|�C�n��dz��]����pGDjH�X>��0
�s�sa6��c��˙q�R�
�(�b�W�KA�a�z]x�b��u>�����3��S(w5Q�X)��{�$(��ea����)�Թ�.	W|y�ҿ��V�"H��O%�lOfI�w$�Z�pW�j�6��~�I��d���:�+���~�R�w�@]{�&�t�p�x�W &�wkFX�ݛ�"����7��Ʋ�b�9/v��U��J�	�xBqcM�h��"�(v%K|�.l����+��$4h��c>���" ���:c;｝���kt�I��.r��|.�f-���)Z?(��֊��u�~����!�_��م��iJ���{���l���6?|B�Ս�1x���)b��JWh�����y��/n+>��.}6��B���6}�}^q�Fcd$�5+�N���2�Q`�z{�2�E{���)@���q�LbYsw�4�o��Z�@�{���m��J�����f�|��=�a�{)B����e���qPf[[�C/��pJ�j?AdScMCM��C$�$�x71��][a;��EK�L��BI���|Fu���[;�iL��&�k����Z�H*�!«��:��h�X!9�*��r��c�"����%J�jw)�ʰ��N5�ֻ�(q�y��*�}6778��R�̼��q�"�m1�%���9��v�TQ��LaW���Y-]�����u>\r
r��� �T�k�z�N�5�������P�����
�ؼ���0�*�4v�^�{!�Qݡ@��1u��UЇ�4�`�E��� He0b���[A�2�i�	�$�l�:���rGM1�u��1Kp��'�1ك<� 0@?]��燄%���!��z�+ρ��)�-����P�w�=#s���b����5ŕ�z>����9)ǘ�`��[�dGDN���� sg΃'-���}Ht�/��狸�[%�N�|+�{�Τ� ��oh#ѾM߁�~~7qފy����s[��2q^�/���S� ��ɴ� g����J P�B�sa˱�!��4u�3R#�k�Q@��jRKǠ �h,��i�%�.C܀>]���-�"��8�Ԯ�:�*��6jN�\�e�����-=/ه T���fXHg0~�Zu��ۼ���-�2|EµT�Rug,��ϘD@W��'#xCHqqG��Ϯ=��3�Ȑ�3��bJ�XH�+p�U�4��Ï��z�}��9���b_�<_u�^V�S��Q���g}�����-����"�4�NΥ��,��ΐ���1�<�)���/��oUZ��hF����W
S�rD]�p�j�q��:�3�b�۱7�� P��x�Z���򼉈M�;�i�A|�w�a��ɔ�x~u���O��煆��M�'#}�0�S�5�������G��#��|1���8�LY�~�+ظ����N�7F�c��J���|U��Вd��p�$�u�, ��,�٭���F�U���>{��8�(�?6���� ��P'9�@�ĭ��6-"��U�{�o��HW�[��j2��~�C���1�=@����������]�uMb����O�j�}��\T@	��+��R+k]����Ge���(�l�ǣ��˟�������]�-�-;��mTEY�vM/�M(B�b�/Mb#�h�����]����f�?����]�m]��q-�
�L�L˳@� h�xYĬ��� �e�>�
�@�ѫ�Df��e$8쟢�GP(w���xô:v��g�����'�{�P�/ ��[U!9��@K�xش�9�6M��j��Ů���t{NQe�f:W)JaN�s�ch��4y����Ѩ4I�)�s)��MfR
X?�tt%�@��rH��x��Vo;�/k�W�m�`��N�jV��Y#�}�����(u"F��`��DT��H5�.Y8#բ;e��h�9�U֥U�bӹ���pّFd&�Q�g�G�@�Y `fE���֪�C	��f�����"h��j�;�y�U���s���Iut{�|�D�i�Q�5�M��L6�G�}�
�*:EB�Q�Y6+Jw��)k�\wB�R�2�M��X�"[���IQol�m���M�UN	�	D~�H눙�\^�e6Tζ�@�h���8�̧�R	��8^���5���Z>��}����Z����l�mg�e����h�ٽt�,�7H�ף��&��9�����q���]��KUc���\j��s�_'N��c����:�7pQL>[NPF�������SԐ��@\_&%��x�d��>r������+.c������$�{��G;�E�J��v+�$r���x��������nk�#Tc�D`��~�d�^�[ܟ$�6�@�]�|��P�9�_H��K}����t��,��C�.�2x�|@�S��8tQf���_�a���� ��7S1�a��y�{�qy^uP��%پ���F�Ҙ%�n��E&o,�W�Ek�|�|Eh6qJ�8���$�j!x��9\����|�UV��/��;�0.���i��-R�&?⟆��m2��'t�Wm��z�%V�$��|$˯��S��@zǥ�A X�e*�qW?3K�1�Tp���ɀ����(��QK�26�L����z�b!���3�D*�+%fj���B���WA����5~{zm��qC��.UW�F*	G�;1ٌ�i��enǼ�-T/�r�v��dy�9Rh���	p���-�63�����yHa��c�"WwVT�Z�RL�7�^
���a�6��`�.����Nu��k��}�)��V����%����l�6���1$;<<ӭ�B2��k`c����%��  Ic]��f%�I��=a���؃�1?b�E��nC�w�ť�Y�kC@�t�G#�sl�#���!$��*O(�Y�+���E��%�n��j�[��$IA�
����c�Ø���=�8�wkۺZ	��5��V�أ�"UQ!o���/��Y�
��i�F,V�D̎UD���"��XU��qBX�*�L'��$2�΁��� ��+�S��OHw%���y�dg�Ee�OE	�y��:���v���~�X]z*��i�&`h��b��E�˅�C���%0���[?����*��!��s(�j����jv�+�I��%Xm�K����ތ[�V:3���8�� 	���2i������ 0�7����t��Qb�x�2�dK���=Xs�����$��Þ����
�\X��8l����]�H_t�{;{ RhCy�����'+J�EBN�B{cݞL!�}�c��j��>
l��a��yng�O����␀H��=����g#��X�|a?��A�KU��
�m��0�ڒO�PﵾbJ�n��/���c�q�������l$����z�]�����,k�Fקw����G�Ǭ$�FM���"6W�QM>^EK(w�O&�ՙ��9j���9�鮬:	��5`��c���9O��[�!�������@1����,L�ҡ�S����{�PΪ
���DxL�m&ӫ��7��0�@ A
K��{���f͒So!�ݱ1ti�Ծ�J����-A#�츑���jx�c��]�r���ѱ8��y��Z��z�4�M� �3cQV�/J@W�-�NI~3jW���a����%Cs@T���f�sq�����p��x��P�D�o�[?���C	D�����#��v��9�A��̫Z%��v.�>6��. ��o�G��w�$@V�
�8(m�jk��h d��Y��1���Cr��T((-�N�^zN��1F��L�ph�g		$}�[��m2�(ă����ᴠ��H��K�V�8�y�9|���q���Ύ7%�<�7FV^!�IV �.�LXA�g�)ds��DJ%9=���$�	�`��aOx��T��\D��Q�]7P���	��ICVM��$Q�Uk�`p��W������]�!B�����y��H�����05���)菏��ud��L��xʔ�����?�o�ȧ�������M�n���?�d��ڰ�auH�s�y#�F<�$&����o��?���WC��d�����a,�N"�N�'��Z&�N:F�F֯�1�Z&�4i+��!��o�ژ�����,�[�s�0���I-m��zY��x������Ig�O$_o�#}n�[�y8St;t��#q0|�_��7�\$��.97������g(�3��y��$j��q�5��F�D,�_)��u���q�*�'i���8hs�{�������0.s�j)�~��2�`��*��vwe���~Fb2�����L���?��0��]����·	��P�n���#�|&�h�d�/�q���z�8o�ӁTa��)jFA�?Q���V7�|o���#O�v���"����㭮���9�Ux��B��!�I��?��
�&T�j1�$�?T�g��N)o�t�⍕C1g(w_]��O��j��Ѻ}U��$��rv�+�J��MWU�n��~��ڻ��}�IȞ9ny�"���<�`�gfD�YQ9Q>��FT�*�`V����nL�w�Of9�9�}$�X�jDo�DW������@k��T�������d��?�`�T[ϳ��5dV/���T�l\
6WD��z�S��>�����se<�Pt���1J����<zy\P#6L��|���?CW"*[N5f$�Zr�dt\�>�p� ]��X�����VO.#�X�K����Z�c$s{����0�{�7tL])�#@c���@�>
sm������k�o<�F�g�a$��f�\���_i�tP=���T6~d�^SH38�=�&0��o�i��O��fC�f���9Ի��P�&![�bIBV�]���)����zYE�Gډ���-��<`:4K��r͟1ܙ��^�/���v>�����Â�WS���&�K@=�K��}.��[��QB��ye6$����?h�P]{�*@�}gV��%w����1m��->�[��[(�ϵ�J�+�%�N3D�����vS 8�*��,�@>�Y��
�E����?����` ���OV�mT���g��B���w;u��e��gj_c�>��:̇����n�oŲ�ţ�nI�8jR���0vq�t�~r�_��H��R���o�"u��s׌&�/əF6�|��i��"E�a�Cg��kn^i��i"1}�������������*>�؀B�t��`wM��8K�ړ�gP�;�6�޷V/�����8�3<�; �|���ֳ���g�뎳,���ض���,4_�0\�wBRi9���)�b'Lf�Wur���U��:�R�w���D��-�J��Y��L���y,�ߌ����8
؉].8�U���x������&�t�)����䍡ё3Y� ���W��&c�2�ȡ��V���^�]�þ�U�2򼯔mE:Eze��'eX�Sn@~,�}�Cp��� Ş )�fw h9�*���dϸ<�M��j��oO�NG�"��okjB��O]J�2#�gjFB��ޞP��J���%�<?���3��Ƿ�""P�5�ZC�r�Ii�Jh�tP桝z�� �����>�-}�C��M�t���eK]i�z����/��gY���T9�ڈ��;�;�ej�s,f����_X�~�C;N�vL��
�.F8VY,�w{����U�r���;�KqAu[Zc0%ԩij��N�K�.TO�XR��%���e0�7�.~�:cy�`O���G��lGu�2��:�n������ѫ�26sw��r���
��<uz�i4[���D�����7�1���x���5c4W��#i��]��+�l�ul�����{�e��+jЍ�6�O���=��W���Y۰��|��=�e�(\4��2\p`�PX8��LG��-݇�=m)wiB�˄2���3^�R�#�b�0 �f [�|��v��w�am��&}R�}@��g��8D'��_�X�����4eL��j K6Ԅ��]�a-8��ýt��-?��ףm�yZM��O3ay��]�g���"�\�8K�E��\��=W�V:>M*������t�n�<bb�R���f�Eq@�X��\�,��x�����g����27-��J��x&�������g�P"`���Q�'[�����p�jJf��v��av�lAxwÑ�Ǿ�Y0La׆�痜�_��p#���P�À�e@�iw=r7���B�Ȅ���q��եc�P���E���S��_j�ŵc\���e��e;.[�$���(R [���x��X�B¸�6=>�>���%�7���c-m�,VRe8��PO�����2'Ӊ�����=\$���vxT�V@���}�v���"-\Ln����E?�v�[���S��	*�%3����5���/F〔��(uxK��(^9:2=Da����-�w�S�J�C�{*����.j��Ic�ɥ�9�(I�&�գH�x��4�˄���^{}��(�uki�3nO��9����,y+q8��;Ʋ�,"��עKvŃ@��w�[��F�$��'f��+%E�q��(hf2�Q\�Ba�{�����E%!��M(���\�G7<�!�	��\5�s���ubU.�����0e�D� ��X��@��ʮ�n�eW�=�z�?O��K�y�;9�	�4��x�U-Eb��#� ��N�F��v�!A�F�Q�b׮�`��I���3�rX���R��|�.��IȐ�p��?��Y�{�͌d�`��O�C>��W���ϡBpX�����d�5�e����
���$����<�$�;�Ji@��)��c>C��v�Q�Tp��� 9n�yPz� ��ɮ0 n.Z�b���"�N�T^aaS{?�kXė�C�F,S�l�}��z+GQ��qLѯYt��
P��6�M���:%�۾E��4rq�ԅ_����M�����g �Վp��������K�ii�9�7�%��u��+��կ#�@j�e�!U�`�Qu��-��uB%��<�7�w�=���̝���*���Fq�-�	j,���~�Z�~/�'6��ؠ��{�ݗ��FOC Ezŗ)B��m~e�<br�ޡb�:�vJ�֋9�ʘ���w;�8�}r���Y�]������yB��_�`N�Y8��0��~��@ ����_���֯9i���q܆aY&z�:��B>�Wx^�������]�1b�[�0�6xlA{vq�6�G����Bs����1����B�豧v�\���3"�\%f=�QU���q]r�	��63�����^t�����C�a2	�-�o̠^��������,P��uO�fDfG���LJ;��?`�0��v�:��2K�vitFs(X��jYѩcwa���u�x����\��`Q�|��@;BT��_K6�A����M�DF�^Ū�N�g��q#b��zė�'�K�����y'��V
=2�-��y��K/:�ZC[�'{��G����U&F��9i�8v����D=rE�v�t$����j%�rb:%%t��y2��
Q�N`5�t�pCr!��;��Ϩ�Q��WH2/rW����h�7v���8 !��e=�ͯ-ƭ������hG�MC��2Ëp�7 lO�%,�>�r��xQ�
���6��~Ҁvk�d���8�%f�|{���!�ͩ��[r0U-�n݉w�\z��+A�,V.t9Eا����O$��{�IB|��N�a#%�Z ��N�܄��JpD0ڕ�͕A~Y�M��2Q?��	�'��.�O^<����i�7N��U�yNq�7���oΖb�o�}(�nP>����<��gA�zɻL�e�d`a�'��1d���F�>M�	Bғξ[��^TWȺ�8���i��(&^�4 <�ꃮ���-���7�\�6FW��큕��A����y? �.a' �j',��p�;�"�<�ܐ0�\պ��B|!�C��b�Zݤ!ڃ���7�|¾x�2�N�K㻨03��X���XWz�A�8�5ܙ�5�@{�������i������е�!X��ݻ�������4S����\����ۓ�N?R(3�����(��t���7~� �2����I
�-R��g0�B�9�)���.��s9�.v�]�I�R�o���	@�� �����|D��Ik�A{��V�R�S���d�?b�s�DI��~�J̱I�}W/g�t�r +9}�i���������X�<�B��̊�Z�b�߳8�����´��r#�����ꄕ�]�w�Vv��đWQ�tB9��:��1}���l���.�ț(G�Z�V�|����`!L��P�_��_*Tmo�#�c8l���vL*ִ�zv����
,|�$���M�7��ð#Y��`���BZ��v���a�h��̐6�0(�,��7/�Da=Z��^�$,�����3�>�Dw���=Fn�
!ߍ�jZ�|P���\�=����l��dE�ω ս`.1o�?��C"K9��i�J%K �2��Òc�lT����[�(��IL�2�%;�V��NRFBwk^�cCe%.��zѻkWu�_�����4�)_聀x~����^Xk�l�n�y��V�EW���q�1���e_�����7(q��yg�-M'h�O�+�[��;�W��Z���3͈��k�Mv$��	'm��I�
%|�Hp= t���3t��}�EdC�*.ȷ���������j+��X�x�P�=�.9����De�zj�0Y(��&W<ȵ��k�����!�d3�:.�!W�[� �Hc����z3y˲S`��dڰX�ڡ�"�{C�kuǿ�v�YD|o+��c�� g�l�o#�s9��I�-O���ܾ��� �~�F$��h�;+�����;���^�:�0�4st��6��,L�(����W��6t68F�LX�6��<���������D�2�! �R�-ek�D��,Y�\���pV��QuJ���y0o�����D���o�k6�%y����\���*�D����Ng\�����H���xB�m(+�~��'�&�ՆS��O>���?%@L����]*�[у����M�ً�s��A�����Ni�6y�ޑ���P��Ǥ�{�9@�x�X��_�s &h1}tT���"��h�SG��Z9Qi��4�H2*e���g�x�I�T�B#V�?!��eN�T�d-]"��0�'V
��� ����i�4p1k�a��w�f�?Z������x]�n���8ϴ���,^awq�ܡS���=�F�����g�ZG�Nc4Sv�E�����kS�^�7� �F(T/�d�L�~�M����d\B�r� y��%��Z�v%A������t A�9EZNIlm=�b�R��T�����v:��ʛ�$٫�i�l���0��T;zr��Z���O�⾫�s�z5 ����9CB�^��v>���#B̀�b�!��k���}��̒n⦱��iޱ+������6�q&���mu��1_kV�[��f�R��@D�/����w\�2i��_��TV�O@�#P\<#�����L<k̜�B��]򹳌#��MA��~�ʨ�$�Ad��]8ʹ�H���=���N�4�.��K<rbc��m�k_��?�@���r��4��4�k�ɤ{�oC�Z�<iq�]/3��-�Դ�$����ܯ��MR�.#�i�b����A��a�+�y�C����r���EL
�}�G: |�W8?�Y�G�n��Ӈ�<oo�#d�5[�lD��8>����.+���|H�5�|��� PQM5��*F�tI���������98a�E4�D�C�DJ-�pt(�@�vul�"�)I(�y?|K)qbJ֍�������칤D̛<�S�/g#g/��v�E���$tDin�k��7OA�mZ�}{�@9 ���]{ݤ�D�SQd��@��7�IsQV�}��l�!���˿jL9�^6�!�=���8+F�)BVD��"V���<#z7����m�0�Ä��F W�����FD�tjv�}4�nWͯ�Ft¨�N?�[�*��z�`�1�@V�"�pb�s�+jV\���2���"�W�,�pp����(��C����@Ewє�τƳo	�Mc��) J�g�O�QW�*�l�����dWI}-�)�>�:��G��yM� Dy��nt��0w5�Bֺ��Q�Vr�͊�rj��DU�?d�-�4����]ʣC���*�X�XJ2e�_#8Gxdg0���n�\T#.j�[�Jފc�8{�@H�n
�#�S	=�Ԏ������'!}��K����O�����}���x9�����!�D��~v��0Q�	Mw��D-�%l8f��֭^��	��.D0J�Ж�A�CS�%���Յ4�J�*���ȴ}�]�k���;�w���w�]��as� ɪӖ������:��5���n����G�:�������L�d�;���l�1��@�nC�?V�츾����h.bp�e �JE�{��h�Xp�7��.�S'(���ݜ1X:�C=�ܑ�Զ��{���
��o�JKe	�d����p�����l���?���e���1\oEi����OW��[���_:�[V��L(��$f��?Х�fV�e{��o>Xݣ&� 1#5�st��G5F*M��x�ӭ�����c�H�U{��Bj`��"t�4����sLK���s2���(�Y��TP�d#^z��T��(��-���+�:;>2L.a9gլYz�������e�Р���)��Ӹ�4ɇ.�7>k���ZUv�xJ�&oYU- �
�L�/�P����&:ο��6m��v�d�i1��V;�p��� �>2BA�9c�,z{�D}Fqi�
���xڟ~zYuJ�>�������v/�,�N�G%M鑮�lJ��1�?�_r���ƎN���~�ZHH�n��/����Ȕ�x:� <'ĸ�������,hQ��D��D��[|yR�ׇ r��	ES@���KOF�P�d��YFZs���c�9t����r������Q�|������B�^�?��5M[��-�?"ʩ�pB���qVk�vQnR���'� T���-���=���_������[��.0�-Y�r!}}O���xP�P�+/�f!ǥ���R�#C۞�~V�U"R�٩Æ�
�weo���o�� �^�:U��A޲�L�E 2�R���mñ�>ht�9v�z�<��'����<�����3�7���OVƶ�(7�jG�idt��n��3
��i��+��SM�&�Ҹ��cw�7�=�����}�...U���F�;���Y%K���J�:R�F�*~�n��z<naK(i&H!<i��5���h�f��ew�� �$
P4/r�(*��@Q�pE��Օ���2�yx.K�]MV{��oW(�oQ�Yc#A�~���"��^C��.����>"��l�S�!� Q#���G�2aɴ�ON�s:"���@g��O ��H�3~x�~�f����ز��/���Ti��E���f�b�OR]D��#)���_�6=0���sKM�N��^��hI	K���?�g� � e>��~�h��Z����][S�q��hQ����P(rm��h���!<d%v�_O4�؝P��a(��W.�{� l�  �W�\�|��D{i��M*df���!�O��8��@�(Z>, I�)E�gY0ofN���o�H��.��z�c�
����h�(rPJ�2���/���E��o/�
4R�c��%�c�z��A݈�#S10����v{B~�]����x�d��t��ī~q`��&����Ts���sb�1u��_�'�b��x�[�,L�G���V��un���P���X�3�T��vE���~�;��E��R�ķŎ����y��pA��)��%j����K�C�B�|b�>/��=�+��s��x	˛��ٮ5�L0z��8i)�5��y�*�gε9�>�n&����M�>�qP~(�@��S8�
� �N�e��7�,��u��y����2t�.��l!
9�@��4��b_�p�����$ͳ�������s��bS'e\��R՞��!JJ���1ر��z+�*�o�(�e�,^3sG.�� ��lP�u�*S!A!�d����ԇ
�9-�P�e�N`����ι`f{}�"#9>ň/��tvW�i�
�1i�����S	|n���~!�C�����'!�ةQl�S`���C��w�q��A�1l����A��3�Z0��r�r$��;�����L��2{!�V�M�u"�v�1p|�ϳ4�!{vN��E� ���Խ�3n��JlD~Lt�j�r0sS��� 5F��2�ĂG�q�~�ۯ���u	�	��,<3t�T)��lw�i�����,=!��Da-;$��#*��C�=�V�J�]��(s���v�����H�^0;��a�m"���"*�3�4�ă;�L����2�"l���0�.�_�`�I;�V2���E'�d\)��,�k�Z����dڸN�� ���"qJ(�!G9y��uw��cɏO
�A�^�o�)�ʴ�|�i��sS�']k�|[�&m�`��/�Cbk��!sH�f��[	'T�T���դ+����S"��%�UCw�>(����0��/��6�7��)8�k��Z����l����t��n���m��"��ټ���\kJ�#�!س�f�3�;�^m�E� 8���:�4@)������/�.������(�����j��`i����j���Sy2,8���),����a���to8,�#+zz�k>Ic9��Y؉;��t`kݓI�-��^���G�����}� ��-�@W��mm���.`L��1͍v������2��f���X�Op�U�E:��2����<nW�����^�L�f�[p6��A��m��f��r�He����c���`cZ0�`�ڟ�ҶU�B[/#vc������r�?&m�PPU�S+vg���÷���t��|F�8Ǽ��DJ"�1������c���i�٠=U��L�3"��r��YI.t_��W��s���Xe�O�*L�.UZ8����28d��`Ǡ��&/���Y��Q�g��Cӝ�;fXF�.����ݜ��E��@Siz)9��
6&eX�Py��|��<�x�Pɣ,�k��YW$�ꋽG�(ͭm���PO�(uN�]����sF 	dx(46P�K6��:	a�;�� �Y��ZI�&��yn�5²��F������o΄�.�$_�܍-��죊���i��:]��%d��� ���Y7��1��~p	gb?�S�!���T�M�mWg�x6$Fh~���j��F���o�
T%���B]i-.bA��/�������b5^��?�6[��
�����"q2�W���.��i��/��9�hD[�4��̃��JB���I0ǽ���4�÷�E2;{Y���������K<.�hq�tB>W�[r������X��{:�u&��ǜ�|�_o�ʦI�6�~�ggzsjy��f)D�7�v���8|�I�`�U�?:?!�3zt���m�0�g!��>g���
v��}�m�{I�!�f-{�v_:��s4��(v'J�u2rMr@5}����wHi�7{�,����֤HH����&F��!���(c����j��WZp��%��i!_�x�.|{5�9j�E߈3J#?�^牝�g�����1 �T�*�I�
��>f.��Y
���YC@nw�z�E5��rF�+��C1���m��m �X�c��/It�h�pB-LO�z�^���ι죆���}㝯� 0�;h8}�f���`��}$)�~������D���Z�GV�<6{�>���S�0k�.�� .TWbs$�mW��`\GH����j�Jj��[���z������s)�d&J
�-_߂��x�yp%�kKB�l+�Z��`���8S�+ڻ_ɒ�~ٴ�^��l���o��k)1t$I�븜S������P���(���<M�+��l����B����ۃf~���6�n�-�N�\�4�P�{e1%_jI���р���)������p�=B~5e�N/֒�����i��YG�i�.oa��0��2��F	�[/J*� J~��Ҩ�X�9b�j���zg�oOĀ�Tyyv��5u�#u�0��D>B2���{)��vZ���q*�1p�n�I�Y�aLf�n���mzmж�=ܵ�(\حgi���g(���Ff���Ϣ�0�ۓ����e���jf`�{����Ru׽8��ڥJe�E`G\U�	�<OW�O4���Ddʡ� <�����`i���-$��pg��]�Q�io�r9�~*J��7 �.#؏Qv��7O���+�w�B���M6�b�=Y7���x�����6�f}�I]�NB�!�荿A:onҙ�Q��Z��оx{'��Z��%Ҋ�2���b-&�3Q'�ق��@~"��E��
^�1���蝆F�S��gaL�ȫ,0�l�����Dv]ě]���[={u^o�^�)�G����&��u_�^��� އ��G��~yX�p� �{G� �S�&��m���tz�l�����s��Hl7�Z9��*Q��Xb�C�w�9�)Q����M�W��g���?2	�R@���d!)�7 +���vA�ƣ�4���˅*��5n�J�{.�O����eSCy3b��y��6$t�aO���倳z��<	�"��W4���ݕ����a3[��6�>:T���*��1�L��h�V-*~�$3��#�H�1G���F�H`�u�.��L�A�Ŭ}�F�uO4�J�u�[(�i��dӌ�����sȁ�G���8э*�8�7��ù���AK�\�?�=+Z��B�z�QJ@�*>���Ԣ�T�v��,�2c��}J�5�/�U��^ٓ��@j_��RN8!ɱM��V����kq!͖��DE^�H� ��UϪ����ӹ��X�Jf�� 7)�hčZe�2����g�o0���Z�@�}3�E 	k��a�
���I��߈$�R,|�sШ*��?x����Xv(³��$�-��SD�Ao8��%��@��T�����پeg׺����ǲ�o8�)e����	�얆���?Xi�H�	� �=��xĜ�w�;�zZ6�$?�P��2y�)!
�#zA>;�uk9O�ӛ�-褌ʲ��<�+͑�XLF�=q��k��lmoXơ�@�?᝙W�Tg�95�m/��;xd�y���F:^�Ui�#eU��xs�r�t�T��m�i��Z��4�0�Į�i���H|��Ñ��s�ke7ޣ$n�h?da�c��R��*=��� ���NI&�L@����SH�PH�,�[X�y,_�W_����Y�
*<�S�xvl��O硒WQI@��4X�-��RIkJ5Ex�,��:1�В�%���{9>����t�|�=�I�迤#w��vb������xuXx�r5�m��&��"�o�Ԯa׌ ��1q�CW��Vz�7��I����9
Q���c��g@.
R�2�g��`ԶV$�YYHT�t���ٰ��?�����=�lCr��S�o�,G;��dx�r��BY���lG�8Bjn8���N<�G���Xe��sՕl�<�j%x�&)�{�)�pqvm��V��g��6�����E���WE��,Ec�ЎhY���:�#���~�@G�|}�~�hES����x[��:�'�Ep�$����TV%=C�j��[�[Yl4Ee;����x>�/�seG`��8m��C/s�_E�w}C�o�C��On���p�}�M&&��>��kՄA�A'�S��|���떬�\7[�<�`��Q((*���k4%�N3�Cz�D�±^��\��y�q��9�(�t��3lǖћ�t�6��Y.�n®��j:�?�wY����|�A�Z�H,��jO��Z�T%�݃�b�l��2�,P�C?ðSΧ��;2�bKKB����t�ۂ��,��9N�S��H��\�u-�08�t#aD�;\0�3AH+o��|OC�
x��o�Oq]�o��L"#>\�x
pط��J&ԉ��G�J���ۧ>�P�zTƵ�D�7y���W*��1�j_6.k�4��a`x�`��ߨ��oD!xR\O�0������n!���}�K�u�H$�Y�Kjʲ���,���1xɰ�P��L/ѫ8����S$����*���/�kh)�v(����������e$��Pѐeo�^�N1�u���O<�z~LE�Cq5W!��9���)�en�ƛF�=����,C��CP�*�X!��� !L�׏�&w��4].��,>�r6p3=���m�e����eH�%K�0k-"��V�����M"���Q�K-��r�>����C2�5������]LM�wd:�*�9�G|���YfAi��/ї$T9��֘�EV�ôI_���R�/�m\!�vUr�	��/h�&m�������1(���b���Q_dewhD��c���H/�5j���̧����E�!�{����Q�f\X�HY �ų=�U��6;����bi�Sũ�LL�W-���U��f��Y/��ߊd7�6���.
Y����J}��z��ɸ��X���p[+��u��Ec�#��������FVB�{�wn�0��)���@X(0=_�+�ܤ�O;�~�+���%��a�ИSq��t9&�y��M�ʬeU�FB#�b���u��*~i_2&wIL�&� �V��|�Wt�w��`��R��[}n+�Z��9���T~��z���;�H�P{.���@K��&�-���p��v��y�p�ms�K��	t����Ƥ[p�ظD�yS��ޤp�b�S�ܰ�U��h;d�BdL���wJE���!��&сf���m�a ��ĉIG�@N�o�bCt��ؤi��u&��=��]8r�j�/F��b��ҐEϑn�g��$��v��fv��1!	���C=t����d$�]�4�k�!�j��؉r��ݡ(O"��]=���Ŋ0D�*$ڗ@=�r�+��Coh��Q�+��+������4�X�����z@��R��7���n
ջu@��<�M��U_����^($�)�7W3oD�%�hè�ݣ?y>�7�6La�>��ukx5���@���"��\��H)�T�_I������LΖ�������f�ݠI0G��&�5b���Qgb��L�r���F����"ը�Yֺ��2^蘋`zU�G^�3L��K��}�����Olf-�*D�[����־�'�=u���o;���9E�L�b�G���G<?v?(�N`�ь�N�)�����-�}R�,N�5dǯ@�p����Y�<�07z��~!k7��VT��P��AN���d�7���g���D�,~~�@<�Y��8޲Y}�&�{�r��ʨ��?���4��lz�ʮ^�$J��L������<��efB���"9=�qp� ��ﶻ�an#���iBt?z���BȤ·o��,��)f|���|��d5�A�����{��KD-�75,י�,1/�4(�}���˴R�֯�G,����O|��8����v��=-@��9���o���N6����y�d̳3PA��1��!ju86H?��q�����㟐{���U�@i���Ӆ(Z�D��u�
35��?}�nֶ*^]+<��g��8�Lr�x�;tZU�D�]v*c��	we��<�A���Z�',�����ɔ P��#v�h`R*��Lc���XΥ�5��m�d6'���c����X��P��𘇙�q>�_][�b�!��4Y�����t���P(F�q.A	�7a�PΡ��Cˡ����6b�X�!��r(g������ *�w ��v��_5�>}r?���@Z�%<�Zh�W$`�U@�Ͽ_��I���8��2r�Z0�Ϧ.�V���|JGi�>0I�N�f�.8ȚYPLL�����n�_2�2��� ��<�[�K���� �jp�9���� J;�b�{����@ˠ[6�Tu%lӛ`c�\Ns�Vр김Om�S��!A��؀��N����
�=����Z�h���MA�3�n�$f\���!��0�ޕ��EH�ꘓpV��I����zw�$!�KE�lx=m2��e}<����Ȝ2l�QP�n~��#A�۠�ǹH`��ŭZ�K��(O�W�%��zT�W�b�`^ѧ�Ƥ��@=`��ԗ�&�dQhhv��C���?�/0���ҷtL�s�j�3�X�47?�^�u �X܂6S���v�c�������#,�¸�K�h ���#��?��?�V#��MF�u���jh�*k���xK�T���5�5���#�l�)@���Ѓ�&{V���rH�&��~�v�jF'�ٳ��S
Q�MmG�/�71�#"E��Ge���t�r_��v�,J+	|!II%y�T񏭨I���A�+���8�o;  e�	��-�=H!˫sO�����ŎLt`�ۑ,
()�j��!�uR�mxp�0�vJ8qi%�֘Ӷ&Qc�2u-
��R�u�N},xqS�� �_s�7Ü�e���Z:�R0t�ZԬ� �)��#��z*��2ȉ�Sm.�ֆ��/I��v����%�t~:.w�?g�"��ď͖���I2z��ft�O.5��GMc�����E�|�h����;�(�2-\j ������o�_З�E骫^M�s�QE;m�����²�6w|
�Cz�j��3w`qj�_�)��2�Ŷ���"t���G�1x,����@KT7y�j�Q�Չ����3P~�^'C��!B�$�O<������2=��k����͋od�O�ށ�̊QI�&%��O1�Q)�n��5��J�jU�7�1xC4B+ 68�"z���(�I��=�B�Mo&��۾��)$aO�Em/	�r���=wVx';�Q�,ڞǊ)���1=�&^�! �9���f���Ee�8/5A��l؟��J��ɵ�]W���JJC?��*�dU�,�'���~1��[�q��J� ����&⭟V��A�-����VS����tQ	J?��e��`�v�E�
�K��Nc�T��*?��r&�[t�&�8������˦1ggF�"{ɫ��y�BԎ4�ϔŴI����?�z����_.�]����#���0�
(�m�HMuZ�Kw*��Պ�9���?��� �Y����G4e'��n��;
�JQݧ45��!(�$��;-0�A�k�'"��*v,5�Y�_`���³{/p���HH�:�oɡ�WB=|?�Y+�Z��1�7h�V5LBS~��,�%��7�����I���%?v�1Cj�����O�.�K���y�-�	�y"	�x�Q���.���]YX��<#�zzJ�v��O4��?+f�z��m�����OY7%��`3�%�9ˑC�����z�w����Y�\�6��W L9Yo���G��<~���+ϸqpf�:
s88���{���=y%�/�J��tƚ���yF��&��Iy���COM�!	�o��Or��	BB|�C��=����bɒ�G�~�r���qҐ���<O}S�
@l�V����%QF��Jx�eI:;�";S��mw�Ҷ0�bUȣ��(����i�i�XA|����m�.j�|���+eA���
��������ާ�}�PW C�ѐa��KUO�
E��)@�;ѝ�+M	+.�p��B�:�m��xC0��-�����{�Չ�'eK�(Fv��g���5�xR�����;�v��`횵���}�2
��7}?�u�{�&�̉s����
ż���1���_,�Y U>k�r��_��������_.����^���#�q�+un���qKr���3���Z���S,���3�1�n������_b*��|黇d{��!����$Grz��'�/�n1lo}Xm�3�bʵ��54��n,����;kx�fd�� 9X�W��e��;=�M�È٭+ܐ���(��fvs ����P�Y�R̖n��@�̅�]VF�-���Lto9��=�*<�⫿gQ��=WYB8�_p�tp�1�{W�L�Y�)"�=�x��f�31�O K����LUт�����%��~��!^�����M�-��t�A�v/�Ș�ͦ���,���[��i5�;�kyOh��PN@������Ė��_|8uY|�ҩF!�n��ȶd�s�.��M���K怼E�bJ=�Oc�ʫ���j���o��Ў�:�I JnX�;L;�vLݣ�Q�8G3�=ڿ'�:�]�!��|�W����.�ź��5�
>��u�8��=��B��>�Z<��w���v�-��F��YC_H��F���н@F>�IH��0Y��˩=�b�!=�$ ��[��BH4���T? ��v)��v�I�����/��� $;ܰ�p-���s%�"4,Vu�j��yBm	B��s6����O��\��:x=�+@�!e^�i�h�~a*K2�����R%�-��W�b�Uma�u�g!��A��N��Ӥ(jDA��_]����\����8=áq�NT�®"����.�o)%rc�,�޸�һН�5X{�A��0����э�B���1��"e�cl�����(�ن��q��������(8\��Z���M|�N\�|����|cv �\�_�CR���*�����j�jc ��[S�L�Jm�}������9��Cg��e֪�<>4D�܇�%u=�<(���9��6W~�B�������̶��D�[5�V��E��,d�;�cs�)#Dm5����L���E4�P>�vA\0�[�\���5i	�p@MT�maQ��Sdĩ>PNT��t�=�uAHg�=ݓ0�E�5��^�-)��=�K��G��m�4W��Ĕ<w�8[>B��U���UƐt�u���؅���M�.{�q�^I*(�ӖQ����7ߣ����l�X�ؗ�(3��Cs��0+dp'��>Z*vKOYxO����:�V"<�!��V�E����\°�i��E���/F���ߨVF�����8ɧ\I��tSmm�.�aU#����Tl�!v�޴T��ȴ��`A���z��֝�u:�d�Ǳ{L��O��<���8���P,^L������^�Zs�����'�>;��7��F�*�Lo�i��fu��z\�����5���p�0�~)�2yus]5�T���ͻ��r�HƱQ;ʹ��_���I&�Ê40#L���(����a�F(��X��'ڕH������R霛���� ��#���!=�.�$O�w��n�[��My��禠�T�����C]Х9���G��n 0�~��g̕�$�P�S�o��Oo(��q2jG�Be���}��%2���Y�{����z� ?��h�5��;��l���)�;�Ԙ�Ƙ����Rkjp�Qԅ���J�Ӫ{4#��}���S��*�#�|�<{
�y)�-��l�34��''=a=�X�ݱ�8��5�#	�o���$�$e�S��¢2�I�^�)���P �;Q�ԤkP�'�'mY�T�Ӂ���\e�v�}Q�mX��=Q������s�H��O�Pr�1	�>��dY��uE��i�,�CP��2�S��'zT��e鵹�9oϡO@��8a-4��k��ġ��	�9�!���k�3N��Q��#��ZG��ژ0D��@$���f�}�Vj�<�*4�d+�&��3�r`�J�2����s��#���0���� ��]�)_����UH�]�p�F�5p"�чH�V��T�?x���q-��\|?K!D��G��CD�Pm�9����MD�inԹl��H�I���$T�!P<J�gS�{'��`�'dL�❲lW����m�CK4ؕ	�&}M�
��b=��N��C�L�{��q=�e(d4�V.������t�A��i}ʭ��|O��h�4�A����Y�~�{�=5����	�w�=��$����u@�U��P�O*
N��z�)���z7+j����8BǛ?u�'�N�m��G�0��7a�M�j{��S�F�R��5�e&��¡�a�_��u��!��O�A�ob�F��}�{�J]��������g��{�%j�u���ZD�����
�*��\�3K-�ux*�f����<I#�6���Ԣ�ih���{Ɋw���Z�?E�`8��e\s ����nF����?��q��hp��;�	�r~M�5uE�ּ��<`��������JlU�3�u&h��G����s"X���4�%�50`N�tsK����oSW��]o積S�����<��Z��T{1Q&�J���sֽw�á�i����T�@���N���U5��5JW�İ�+�m7mp���W�3*�2������z�"̄Hb�^�F��
rSuU��lR���8�&��&I��>Abx��G����
3��^D6�I)��ۼE���n����1�J}w��
�N�!�wM�-gm�zx\��S7X~�Ir������)F��!��m��Uߙ	�ȋ����nt��~�������=��4��h��� ����T_aC�(�ʆ�����k|� Ea�Hk��V�����e�7���h%��nb�v�@�kێ�Ϙ�Lhd��ک��;�.	�)˘9�62�Ǐ�	�M�KԂ�O�%�+�U��RE\�Ϛ;����U,IFQ���Q.A�����!��F���SM��L�B��ʨ�#fărX��Ƕ2���2��%V����k#�f�o����d���`T&T��8���7��g}�=J�b��DC;rfdM�;��'x�F�*W�Ȉ󭢑kL`���������U�X�>�e�p�"�b�����U�/�Jۋ�v��o�z<-��$��'��� 6�G����t�U�u��/Y��i��� ��j �^�u�z��C:O�;�(�W:O{�Y+�3#:���"Sz� �h�m�@q>� ��˕�hw�ˉ)(���z�[�b�[�?���4���v� ��oe~��J�T���Z��+[xWJ�9q��_�[v��V�U��H3�����ľ�T��^�2ۢ0wȎ��E+H�l��u��,�²����V�]3��6`o� M@��0=br���e��ɯ�Ǐ���\���t����C��k����C�����,������īF����;�J/x@�_	����4�{>���E&��
�����E��@��5��4f���:	��/�NfKc����Q�js�c�@q.�]����lgu������a����RIuU����vI�ugd%�� �]_7���s��jS�(����7�(�ĉ�����zu4>	L	QJ��ͽQ��\r��
3f�okR⊢�;Нg���� �F����N��B�L1׼i���zQ� ?�C������#~�k��k��Z�~��������*��Ȏ�xS��3��/Xaq%��'	)�C��`�X� ��]H������V�� �9	̑�a�����
��Ǭ>��ۣ1��>h/4���ʭ�ֱ-��rC*$��8G��n�O"�\��l'5b9��FO����w����Oّ����
ݸ�A��*L+�`��p�o< ����K��%�,4�������mcԆ���UHm�rw�g�F���=yn��ճ ����@H�s�*P]z��<�/��OXVy��G��~���w�6��a�Hq����ΎY<f#m���8�A������#��J��� :E��D���K��ս�]nՕ�{$z���rrc�c�AOƿ���+>�-�*Ue���`�-8ҡN�v��=�C����Mq�*Ц.��!���IQ�'$�s�J/:�(��.I�����<�"!i!=u��Q�c[�i��Bx�*��ƶ��� r��l�)���X�?����;����c?gF����c&���cv0b�Q��xΰEFB�M2�"�>PC���6�Q!<�;��R�7U�~���o�#A���,��hEZ/0����C�C��}9Zh��1�]���H���;��a�rƓa��8���/k.e<��xᘂ,��gB���z������`.���՛h%����'ŒH"�-���J�.))��t
&5��sW�?���_�IaZ7�'ߛ�8�MYX��u����Ty��-vf�t��,��U�Y��Np2�_�=��e��}���k��a�zn`��$V�!Z�8p��9f&��-��L�dr���D(���~����V�=��>��}�X,�e���^�E֢�����;�WA?��=ӟ�Z.�d�UBnj���P�T��0Xm��'x�b�7�B��� Y'Jf`_�7~��,�n;�sb���	��A�s���0�v�x���f��zvj��OZ�4������{7���q����=��n�`|n�mD�΅�H���u��봷�+�,&�kk�usŤX������~x>���e#t��3
A��&����@��J_�q�9����hL�����7�F"�Ug�+��I�*���毄��54D��ї&��6@M�ɓ����z�C��Ó����F|Rq��ph�(4^R��Ѩ�!^v���2���
+�����l@n{���H&rrYpK�
�K�[�Ab��}}"�������3�V��?z����i3X���Ӳ�l��S|���.�7M8�j�ٳ}��+��Z��Y�|	0d��2A�3sn�p/⡾]~��MN#�/O9��u���&D�w8�W��je�!��z��-G��V��K4E������Y�]��N�I�x�{1�MW�Tős�� �(�:�"B~����}��+m����[�}m�㝒��J���շ�0t.�aI~��.�2���l/q�~�>Nܚk� 7y��n =�T���e�T���[�H�|!�͙��jb�NҊ��=�+�����
4~����N�W ��E��ihl�+y� �`�͝2��	�~_��+�z�⍼	5��}����x�]'G����Rf�Fqo�ϰ�D*�/z�Hv@�şk�P+"�A��.�>*k9����F��˯"ᶫ�J�7m���۹�ߵh�K�;��ɸ���,���F���̽<9G�)J�q�2�y]�|��]Ddv�G�9�kG�H�#{��K��{��U�ڶQc�R�j�l��g!��
0�2[�.����fըG=^����Q�^i�������j'|z�"��
bF��/a�[̞2B=�H�c�8���~d��[����Fn�9���VZ�����7��>	��u_�"<��oѦ0��Μ#�"����P�Y���l�7��' ��_�H���aY��6�`�p�L{��'�ﺞ��Lo���y���uWu�)3q8�r�g˙��jWf�!)}�6`��?��T�۲M�HaM()�g����G1����.����Ů��_8���� �*\C¬8|����x��b��>�Rk2C'���T��><hfL�t�ğ���ڕ.�z�\�Q���K��EG��fV�T�
g�_��M� ��x���ǗZZ����COL�?��*�c����H��%xF�ޗ���3��+)���<�()�tg�Xql��q�6�`l8�&r�R��7�[��X;q��)w���+�u�$��V����3���''�Y�
�46�9�)���\T� [U/�Ux->�'ϖfN�b}s�mG�D<X؈�o$$}���;N��z�:��u�u�eX;yv8�U������f�/UW l�����M��'H,uX���mؐ���*�w��1��@�Y����Z�3)�{�ҿ%f�P]��qA��"�����B���xa�{���QH��3� ��_�?2��tO	��>8=��]�u��l\�B�?e�q��;�tߜ���;ݗ�\���}��~|�%_�C�N� ���a�'��[��a��+�x��7�J(�#����5����2� �8�=�6) C���'y���P���b2���b�M���&~�Z���۪�3(�4�)�׻MH��9W r�{Ad�3�T�l��NT^a�(hc*���P9��
���݌<��
���?�a�4QD���J�`$G�&���\�%����f`F�ޑ%e�v�P�30��uwn2�
#��3p0t��,V�3,����%�'��� B�p���ד[31A�H�����s̜�#tnv�nv��Gt�$/l��%e��Q�g��%��1�6 3Op~����VKAz��Nv�rc����
Zݱs��X:��b>�ex�;��6qo�)N(�(@�M�:�q���%���M��;'��*�^2J�����N��l�E�*_�-���e½i	�>��Έ��`�������ǍN��O�hv��J��t6������9+�a!р����%�i���|���/�87[s<��FT�� G�R����>�T���7W��|u�T;k���Lg��۱|B>����/6�:[<�aAi�aʩI1�:/E�`��-4��[I[�5Aa�M��C�@��ͳB��M��<0D[��c��ζ�����C�%�KdLA~jN���2��J��顔7S� �|���!O�l��K-���l0g`܇��r^2��a(3�y-`&���%���[�R�Kb����0)5 �� ��I������ �X��*n�����՞jշIcQ�N��>%o�.ΕAy4D��(A�|�0���L���{��D{��<�S&=�H,	����ϰ������]�z�,q��s��R�+��(�Ǝn5���mO��)�O5x�i29:L���(J�Φ�6����Gn�N&m��T"�����jQ ���-D��:������騆�"<�	&p�1k(jf�©L��48j�gXk�����
K�QC���$�"����]#r��S"���&�B���;p�,��6	�9⣅�l�"X�du�xL��X��na}�w����	J��iV���|���M~���Uz͂�܀=[{ øs⒐�8��8B�I%/�ƱѐSz�1�;���Ԧ1��sI�S�P���И�go�R%͋x��*7�����&|d8F�:��Z=��U���@�ɰ�cE��M���l�դ1�R6?)�\ %r�w6 fkL���a��֫��ⵋ0�	�M�>�S-g;��&0��8Jg~}.c٪Ww]���z����\D��[�2A���?�݄���W����X+I}�x[1֑��G �s@p6��������<F.�.h�&o�S8qhfB;�}���e�5^�9�$S)1���u8�k@# $V���^������d���`��5����Y�
��E��AكC�5�̗��V���XXO�Ux!��k�*�7��Y�	��\��a��۵>�| 򄨼���+m_�%i���JY@�P��z8�f��/��e��YqL�˴����Mk�1�;�s7��i&��6�9{u��Dt�4���[�	�>�cC7����|��|��`ڋ��	R���A�3�6+;%C>�?�ݐ�1��)���tgT�i�B_�C��v)M;R�M�� Q�s=x�E%�q0����/ﺩ���p��R  Z\=0�)�<���v`��U��b����ϛ'�S��,IxC�e�v�ؒTPW�g07��D�{ψE��nKD�n�|��� 9BX��)s�K8�Z�۵i�#3�QR�I.ɨ�?��Z�}Ф���CεB0T���Ӑyq d%~�]���=�Tw �un>����o���
�Mk#xM2'y����k��ܭh1�C�Y�����	�ͺw�V}�w��"6i,����_���z��%H�R�L�"\�v����w����$�����{�Q���;����jԚ�Y���ƥ��k�4Q��+e�#���)�%��1� D���<�\F~�����l����b���$�#��%���*�:�� w����ol�rh� ��fy[��`:�,t�F�{�%y)v�Ԡ�c�a��Z��";E�����Ji�%m��L��5��o������GAY�}5��;@xu�E��m'�I��Ii^�n���i,r(\�@>�e�Qa���M�@��f�,�*��$i�cQ
���'��<~�I��K6y:gTlm͊L"�m��8=���:�mDT�/�Փ�E�wH����s!�(��ia�6'����z}_���v��3��2��3�8F|��Wp���s��{��9����Ԑዬ�p'�l-�(�x���W0C,Ãj}��"���c��	��ȗx�N�X�o����>7���]c����h�7I��Q~!R�I���왂�;.e��/8�cW��;`әŹ����NI��«���M��ϛ���_�c˪.��g��r�|�r1�B�[���ܠf�O�G`�N��w��nn@��S6�U�͏��@iln|�6Q'�=xb�\.��h�L8K��r�%x�y�҂
R�?�&����)�tB,�5*���>흢�^�pq���Ki	�����a4��>ʆ�f͕Um�l_�0g�Ju�m�%��1�Q�5��*���;X���ϯ(�Z _&J�\�����	�(s�{0(��!���e}'�ߠL�n�1�I���U�x	(�8�h���L��3:8�B��bb
'�Xq�������,ݓN>�"�a�H��:W�Ǫ��$Ŷ[�@KUZ3B8I�B;3u�؄
_{C[� [P��od@[�r�sY��!E�J$�]v�p�C-���(
��M�"�:�j�HS���o�� �7CI�,*�P�o5����M����%	Z[������tu|%E$�u��c�/*h��`���N��"4N����AG�J�E�ɚ�VJ#�-q�j�"c~��IvU
Ľ%�[?�R�'EWՕR,�0B5�G5�S�pG����s���n�e�OQV[Ե�a~="ޛJ�A����b���f�E����A�u>v$K�1����P���i�?r�9�����O���?�o�\vΈ���YU����� ����Pa�[w_?Gb�uQ� 9H&������0�j¶0�Nr:����b�z��:A������cTMB`�����~�E�y���Fd9U�`����i"2���X�r�?��w��lȪ��)�b���@'b�Ua�hYF��[��XoY���Jߏ�׮SC�CKM�!X�j���]W�������s����Tؿa}�{g����ft�����A�!��g#�6K���� ������'��Ӌ��8��u�q�o����v�H�^�tp+��")ٶ�'@�'�40/����^G/:|��!��Ww��ܑ�/��2�q�stok ��8;����Sn�]@ٵ~\Z��N�R���}[W�6�>����.�_�#YfV��7!�w2��EP�:oS��
B����XI\#܏��$r����ߚf�3�^���y�0Fj�1��X7�B����F�GЄ<-�>�G�=�K��aB�K��-ݽ�[,Pй�m�Jq�35����Id:�N%J���"��[�.5	x���׷r�q�����g�鍕��p1�Rj����M+�(���DF����]ā~��7���n�G��"~��ֵG�0�Ѳ���+��%�v��y�,G�5�p;c4��c)kKw iU!�Ԑ�\��N؅���ӸI���D���z�Bĭ�#4/=��A��G7��s�`��K�yC#��Ev�x(���>��࠵�ܮծ��C�\(�3����F�ȝ3���^��{al���f�hdv�xD��	r9����������[O �LqpNP�G���.�CN���YEŵ���N�C��2AhQ�f����*57��hóH�R��x���:�t���Ofp}_.�r��;9�{[苁Ӛpÿ�	x���>�V�x�!��*�K�TN��|j>rap�_F�/y��)���):Ň�ڂ1;i�S4�����0���MDH�qw��Q�q����~F?���*��ݒ���y�(������V�]|�S8���.
�=���I"%�j�af�x�C%���u�|H��i����W�vA���wח�?��wK0��*dt_��y�9�V����4"�6V�"�hb6)$��u��@�᥆�NB��o9��챔"vie�l�P� ��GvOj���B������:�zl�:�,W��{ߡ.^��y>�/���
�&h��?O�K~���҄��)�Lʖ�T|�X`,v\��h(�=��	���6��2�ݏ$���"$�������'mgk����M�����]2�B�������۱i�'ˤi>��0��bVTMdm|\tt,x��o４wBu~b��$z=gq���
���#���=�3�t嫱B�L6���orRRv"f��$K|�F�4�^gU�����;&�&kk������ӱ����A�/X2��s�T$����rY�5��U��䫎�h�>	#w�盯6~v����P�']�!)��������'�����bػ��J�'��3K�'�Y��k��v;-�~��P�LG�����sg�^Ĺ4ۥw]��Or��ְ]����4=cz	1,M^D��)�0.#��Fb��� U� ���/�pP�V����>�ps�<��!4!��\�><�8���ˋ��N�Z5�v$�=:�c��[,�{�9^/׹h�sj��Hִ�k�K�ɉ���,�dyqM�!�'��h�L�j}����-�G�k���:�E�ZGN���Ǹ�4�>���
&�,�9�֒$�*�9 �{ūv�;ö�J6�J.�v~8��ɓ�Ӣ��_�q��TnP&4��~�$�E�G�&7d���Ӹ��us�2��I�7�Z7�'�h��֐��vF,�)L��������-b�n�H�6���Y�o��^JT��p���g�
%�m��v�\��r���k�grR[0}J6�#�nFꮖYxX��Q�-^�|� ��B���́1=�}��s+��
C�a�*B��7��癋V+Qt-ʆ"KnU	���}�@�X���c�In���a��w�bB�7�n�~Ȥ4���o��n(\KF�v�rkJ�����g�;,��<��%��*�-Q�@Xև[�G��dLB9�s�"Т��]{G��8"�o���� ���,t?�RU�t:F�D⃣c�c����S���[�����Vf&�����m�$c�O,mw�i"��X��Y[�$�7��ggZ��M}���回���o�g�?�L{A��ք�<]�8l~D�¤~Ɲ[������Ta��E	,����x�R��L36���6d����M���B��V�O��) (�o�7����/P��=�a���ݹ�lݔB�k��^yP9�DL�J������sA�ȌN`/%#A��k,�"�ߜ�ʢ�̼+�����:��mF�X�<�F���:���1�BUJ��[�Z��H��}��U�gW7T����<�u����8��ߐ��ns΁�A�h���5V���,���Q�-�(�N��)~���J���px�X*ߴ~ D;�HT���Y,%�Cַk���=2C���7(yp�<��V� �Ĥ�I�.NMIj��*���&1,�Dq#�
���_�ͤh`zH���p�d���δEO�'����tú	�:��G{n��6=�����X��(�ޣN���&��kK)0󿧽f*_h�*cuST�=��"��1mr�^3�Z׶6����_���%���H��ૂe���^��U+�ȤƷ�̅�Ӡ�-���.�,��@�Q�� >����f��x+��,��Ne=T�#E�rV'�f��u._o�y|O�8�B�̛�F.�U�h�.R��j���+e�NO�0@��6$�.5�KW�On�G�ij�Xq(�����p���7���.|a�#�A�<�9��=���ZdP{��{jW�V/9��������9�~�i�Zxcb�d�TV�Y`+�n0qB�zd��w�K ���O�Kp����}7z~��-� ��.��[�ԃ������Y���EQ#햙q��>xBA;����1�1�s ڒk�3=N[t5�b^��Z����2̅����[���r�VL��h�+��@�|�z�Z�Ӭ2��?�;j
���Tq��A�e�;.�f�}V�?qB��Y�2l߽s5s���VpX�t�/�&��|	7���
���R��
N���SNz���V�mb�D�Bm�Ɓ�Q��f�yk�r��s(���ҹ����\�S(�8�@SS�'��W�f�P��!�}{��n�}�?��z��|�O��S�(n$i��]��5قԔ5F�8՘9�<F|^v	;��x�\�o�ꀳi��De��׉8�����HL̡3M9��p8���w�@n(�i)H$����"Gg���T=L��6f^�������~�a���S��X7��2���Q���(.�y0�u�n�D���j��_�R&/Q0@O5�񹻖`9�t@��>�%��BHj�DP�����%��S���	>��t�YO �r];,�|<�	���Ogd?\j 	)���&�,�4N���_g�5��;�Ak�φf��
q3�����F��g^&cq�ޖ�gK��,��V���f�MON�z���E�5O��x��	n����|�f������:�3�R�MA��nN�=��|3�R�̺�P)5��7� �g��ׁ��z\��$��)��X�G�ƅ3�LY��F�oq�'E��Y_��8�.�/Z��B���N��>$oO��Mo��>҆zh� =s�-�Fz��	�2\����Q����lr5�]5�a,��6w�y��KL�ZCZh�~���鄏��T_�/;l��\\+-	�Sju�N�x�yJ��S��ƎR�1?9��A�$�d���1����X=TFשּׂ��ԃ� �㤍�j0M�J���I��@p��L<�q$էoH\��Gp7!����5I��m_�ѱ3�;�_�eJ�y7�i���ٗ}.��Ŝ΃8�f
�}���_"y��m^�$�3S���)��	���
ۗa�0��u�c�P_9,�\@��P���?�� ~���tK
I����b�-T�?�.p���Խ��^�1�+8�I0QY>wl��m���7-Ϳ-� j���Q�l�<_��D  �}�J��d����i�/@g�h���{�P�wUuK�@����,����*g�������	¨����Ȥ��U!�o-ʅ2i_���/����6�d&���1�p^����e���ۃ~��Wx���i�&�UTE-�T��.Ϊ�^��Rhxm��Ë�g��	=XÕ�R�<��� L����)G��m݂���9���s�bD�*�G;O��.��3�m_>��*aTX�qdD�^�{'�m�P*w�������"]`����>�+�^e���
���:x�d�x�;��M��xg���D�Y=i��5�]BĂ�DX�%�;3�6NF�z����lU�P���BE|\��P�U�;�d[I�	y/7]�q�%�8�;�V;�
}��b4S	n�uH��ģ��雩��ˎ�@�$��W�i�K�<��U�v��HR8�U�2�PW/

���e%]!XL����-�+_���	O���Zߥ���u�)�����b�x<��r�L����KO���n��ё|��I�ڊ��ԋ��G?���� ���_՞�!3��]xx����?.d#��Ss��]$�ke]�����eH3�n��<��$��7/�n�2�9{$����"�[X�h]�iUҌ����j�աd<֑f��e�=z�Q�c�76��ԦCX��B)�J��b͠���iJp{_���8�6AFp����o��m��������<��2G~��ֲ�/h�+<�X,���ș4�ꄆ����Ol�j�ւ9�`H\�F����ɤ��rt���݂dw��_{Ӹ�˂*�b_��<�~|�,���)�пre��n���|�%�����H/I���[nO�=b�q{)��w���GHA5��j�C����C����z|b�0.B'f��݂BNc��{=�e\ɏ����։?غ��|��/��2O����ɼ=��h�1�]JЊf ��H��Jux	Ú���:��f���x&Q��9��2af��FJ�p?!yq�Pe�7N�]��� ~R��!H�=hl�m��n.���*[���-���)j�ρ�=�?B�:?��|�p/Λ�	^���Z79'�x�[���z&�'U�Y���d�0a ����\�.��2&J'�fe)袺n��j��b�h:K�d7�:�y�W4�	�U[0��>��Q4����������"�'�TT_n6�!Ά��1PRj�1�r��^Ā$��5�j���5]7`8�8�*��7��4$X��D��Y�@�[G�7%8�d�70;A�*�$�,;c�\{�xg3�:	��Js5��םOg� EĴ�r��M�R�e�>�魤�nb'+#6�HU�i��c���n�}�g탺[d ~$�Eww��~���P7dկ���&�'���rm��% Gě�>x-�3�\�����d�O�ul�0\/�B1K�����Wm�(-q3�M��U��Hc4s��bj�pLZ�~�F��WR>�%��H&�7E�� E�2N�����T�q/艓���hTM��)~pm��F�c r�?�lk��4,��5����\��ٰ�\�hj�~+V2�0�(rҒ~�	� ��.xɝlK�&�&?��"Xb/��#tf\噎�9��4!��X���׊Cc (�J�9�b`xE�D��q��y|ĉ
�C�
1�X¦h�L��?��f���=�/%(����n�0*��m9n°�Ncb�o�]8*�)�tE.� �!�j�u8_Q]y}���t��k�X���3�����3���n��9��e"�)��1�3։���M!�Z�B�����a���V����)yf�SǀUTU��{�Uy��F�����\���۬)ُB�yæ�(�\R��\o��"��;�̳�\_<~�-sbk�{*F����G9I�o�Ϩ�e|�e�p� 	��6��QS+f'ẓ'v@�d"�#��6�U�e��+�3�D�VC�G�kqX���F�/'�d�؊e�}��4�j�z#}@}�I$4�;��&#��Ł��' |G�Td>�S�p�$�e��+�ǼQ�G�۷DE�厤[Y��$�S�tT��#�2&y'�b�}YDK��'A��&g*�-:Ϛ|n�zzI���;,�`
qn��pPm��؊ܘ�ޖk��k)�-�|����(�����c=Q��X�CQ�� ��Q�rU>\��w��b���J�V�l�� �	��§����?���Մ(Ki��*��݁B��4��0L^�z�'X'<sC+�9��j�&�d�4��V����d+u	��x2ԼZ��[��XR?�0�@��2��8��U7����\ z���b���?u���|�� �x���o4�8�t�Y�j�:-ב8c�{��eߒ�ı���GA!�}�b�����_ʚ1��t7�M]oU��߉�uǨC��q���Lϸv.�DNQ�~�G����(��A���́�MAt��|fVw~:_K��iu�FJ�wu7	Y�K���2- >�7q�J(2��Ƞt���y%dsʭ����iF��]�Nq����k�ۢΌU5b{w�L�a����8���%�q�#����s��j�$'t��x7u�<5m7�O��d�8�j�1e�g-���qp����n,��δ��n%� �IyX8�u�P�|)ZT�iu�p+��Kz���jZ�k8=xu�=����%�~�N=�C��F���>�2�>J̛ی�!��vr#�𝨔��7Iu���.nʿ�0v�)�����T��U��Ri<>ʖ7�8�p�=�_�֮��v�5�U�p�o��z���j��l�C�H#&Y#3��
q~8����3�2��S�"�$m�|�ʠ�&ߘf�:�>t�lcg	�@�L����&+0��{�̼*z��$}�D��"?�})2ۈ�|uP5R�{uQ���a,�?�$A��O���<rE�t�&'t��ȿ=c�Qdu)/$u��`;�{ZU��N��ЪD��M��>����Q
�tj{]-�&�%r�?rW��;��kȘhK����Z ȃ`��ED�?q���w���5K�(�{������0�c\�K]��M�'x�;�9�/);�&93:=��A�~�ܒ �?���<�DǦ�W��}i�C�"���Ha���&v����M�NiBeA�hX��W�a�i�m�Mg
��uLG	�x���qz͹��"���B��P�����N�J"ߤOy7�I'�&R����Z�1��Ҵ����Q�R��mf�U�C o5-�=�{��Զi���
#�H�7>+(Y��hμ6(�)�"�J�b{�p#�n[4SPP����v�P��o���u��S�o@M�+K��V �@U�òB����fX�	iV�)��n�'F��N��A�s��$�\8�1Ȯ�a 9�Xޯ#,%�cZ˭��n��ݣ5�u"��æ��~�?�3M/Da�(�� �.:)l�Ȁ�u��3l.f�a>K��@�.bu~�s�ɋ0�.}�i�P�k��d�-�GW�G²�O�er>5�Z�6�h�1k�C-*�g
�\D�� .0�[����Qzq��-��'h fq���B�Դ�:5̉d���Q�� p�!7ѿ[,4N��N�>�1����n�:������Um�~VF�)ێ� T]�}g��NK����Q(_3�z<ߺL�LO�VT�6��	�N��%ߟ��E�`�ST������7ͤ�=b��v��9�؞a�H+D��툓ک���)���^.}6�lΣ����&`z%aV�Y�7�E�4��[FM�<6��f�2�1?'� `s�W��lO�r���@,=�Nt�B���;n�������,K�|c���^�v��uR��u��޲��gll�h�N��N�]3�іN6��r�:�t>�aQ��M�M�Q����F�3�K9Fr�~v���(��[������2�P|�Μ��v?X����a��̗��U3AO�N@�QExL��Y�x3��G�7?x�"`�	#`N��J����H�B�m�$�Z���q%Q�� �+��� �x�l��Nb\RU��&
�f̿�s�-�}뷉1�[8�	g{�+q|	�V�D�u����?".kI߅8�����x��{6Ax�]{�sٵVO��^7F"��#��Wra�u>>���*�2X��|���L����Sru��X���A$�w��$�Y�|2��<����CH�!���l)�Ҽ�I�yH���,��0w�KMI�{��+�#D��zj���?PLZ���5�����CWt�C�����m�DF	�����2hk�G;���{2�J2C۲4��l��J�Y?�����������l
�]~���җ���&&���2�ZL��Q~�+��<�}��ɶkGc:7�vm"_zvhv���+��/���]�A��W5GO�]���O}���dHQ��#��l�[�e:�8K"@�	GQG��Ŷ�����x4�3��Q^2- ���L:6Ib�m�hs>b���O���a
�cʑ"�DE,X_�'q�.�gSZyƌk(�r�t���0��u �m��!%�4��kt�8La����
�4·~@��[
�ઽ�w�$��|�q�CttᬂhS'���Lu������
�qt�`�%�b���f�Ul�)�r�p�\6o���+�I0�,"�₈�D�J~#���͌�&� A��� �#V��8>�U�;s���$�l -�PS+�\|�����$�]�*��P���j9�{~1�W�Z���妌<ET�2�p�������l �*��t�����բ�9~��ő�_� ��W�?A�M� ��\��ը���;�c�W��t+8�Sb�+6c�*A{�.�����l8'>
هA���R�66�%O�w��'�^�DĎNpLy�6�9�N��S[����i|R�gb�"ѥ,U�a�?j��3l�4p��A���,_��-n�Z�/X~� !܏�)ȿ�B҄��}�fֺOq+[-���a����s�َѥ��cf^��]8'>G�i����m^\�W��l��p��1�Plnv!�R%�8�b���XF��p���+��a����l�&4E!�X�)YLS� �yB��I����1�����]��7�}1H�N$6;y|�)��+
ƚM�s�a6sb&��rh����o�F��4��v��N��U��$K�uP�(׵���zی�� !��Ȥ`^�2��o*�!�����3���w�g��v�E��R�m�Q���UO^3]����ٶ�:��km~*GqS����ʢ���Ǧ��A�,�3�w6Ю�QW�;y@�$h��8�[@rԁ��sL�-�$z�|���qw%��$]�w�9�*���wI�R��D��#��[+m�FZ�<���O�&�em�r/X� ����7��ȟ�(�JI~t�������ʈٮi��T���#��BY�ZS�������{F��6�g��Pi�}�h{�������k��ؾX�}MV���T��� �`��֏��|zG�yx\�Ol�$��L<����G�y�{#?�����^jK��V�-!0s��iQQ,�� ����k���m9���a'U�ma����F=z������#M��K� 1�PA��1p�Y]��ϕ�$��o��.��V���J�9�yoa�kZ���
���;B(yd�8Ļ�\�xB-�d+}e��Ci����n�w�����߶˽���!�;"�@�td	�6o��)��/���R���+�am��f�~�)�6/���+k]�1
��͌�7n*� E�U�.�Ӣa�J�}��!�Y��_�w�១�SŚ{��5t��cx��$u��D����'�=�ﶎ���:�z��ܰ-~4\�����s��Q���_�YLi�a!���jC%t�rzlK�ZS�F���mK���뿘i
x9,w<=;�)58��iMq?[�KY���Q\ǼN�ļ%�Ԅ�S	�Wz�<�k��{*
�<�E��`J�[�O|���Y��o>�/>m1��n���c^}w,{L�RYez�B��f�ip-ؿ=0�!���m�MJ�� 8�&���d�"4��vGŁ.X���^���&��~V�$�E�nw
�)FP��7��֟wK��@Kb���Tz5ً���5ߌ��������7�Z�kj&H�os<��ʮqs	�Qj�n��q�	��sh�d�S����-r�b�$lT	�'"��ң_䱍jiExw|$d���FS�B\LȎ͢�՗���W�A7��,#�8笏�(b�JcnN�^�e��P��%���[]!G�B��P�Ug�7�v�B1�����X�����K@�m��x'��wʡ�Q�������ƌL�$m����z� �	�K����퓕��_��m��s63O�szܑB� } ��┭���*�u���k��6�ԃ�$�>�6@�h��b�[�14�y����O?#��û1/z�D&	���>��(���D����g5��f�mR�k-+R����o���mN�5�N��zar��Ŗ~���<���U�����\ٵ𫱜]��gv��������%�|.k��5-�H�'Q�O����/t~mrf�[U�q�Yr�T#��x��K��oe��"��û��%@�����	7~WKU��6��/��)�̡��vi�0"�u�N�}�B�
�?)�u���W"��fq��.�_ڼd�;����}�)�i31�f��%A�&�h6Qw2�37u)�Lfx�j�V�-��'���a���)3���s3eGμF�5:�M���H��	�)(ߡ�6_��ÓY-��Y��R��ô�Z�_�;�W��xyj>ə`� 4W���wc:Sc�*U� �u��%z���g��g�e��'=�/���X�oZ��_�f����h�A�C�T���d�{XU8����8��G����I**rB�>�Þ\1�uU�\�l��`��#�(1�Ǒg��`H�a��O�%Zx�&a-��r�Hy{��y�q���si`v��ڸ�Ы�c)��OZG��ƹ�������p��o&
u��DӇ����k�8�w�S�܏��mCN����� �y�o�	 �U`�:��q~����e��w�P��+ψ>BwU���uoq!�sLPA�+悩���XK��� <��r��R�($�ت1�WV���6Nf�(���Z1�f�жd4��뾽T�M�)��L��o/.oT�~ƒNf��X��ޟW?��S�sƀN��|>8%���[Ĝu�����%9��\?Z/�1��C/������M�=2 $��ϩ��iq��K.���r�9�]s"�n
����n���ɚ�õWu)돢� T��m���)���� ��XO>~"��6��'�?ݓ#����o��&f��}A-�	:-����+֯�9|<��|<���$E�쁸���4 �sd/��?�A7�S���b�8��Z-o��G�.���g��5r���V��f*y�㎵B+��L������~DԳbq����-Ǎ�H@�}iҝ�Rh�\t�l��H�8�rCKD��{��@�(���IX�
8��Ç�̽��x8T�W����+��Q�ۣt��U�v*>�.IEH�J����Nv�>�µ�y��XMd?�@��á�jx?{����s�������
w]���o��m߱��˶}��:l-1�7ޫjUKK�S|��u�.��\�E�d�RJ{�5M~��������z���ɞ��3�C�M�Vmd��uշ�T �
�J�\�9!���X����Dk��D'7S

9k��1�y[�Qe������4(�D�O�ʝ�4J0��m���;��f�3�g��2�����oh�P`��x~�era�@<?�F,�՟Xi3��m�Yه��e�yU���T�+WMa0%���/�S��L�_j?��k1�3�h�G�\8S����	1`�=}��Ő}�(�v�13�x�5��KwT�Nq��x�Sq��pq�0z��E�Q՘ꙿ2/U�;�;�t�N����?o1�Ή>U=:�[��[������|m.����s:�0T�n��	e��y��V\%4)�"� �>���Zskᘗ����eF��I:oa��uw��}kb�M�1�(�Dh���u��o�A��:{85���@J!e�=<-���5�-�W
�{
{��p��� &$��%3ʹ�S�t��3��Kטv�M�^I4q)��.�_,���_�&��؈*�0`Ӡt,R)6q0���I��|���0�6�Oі!!wc�Z��u�H�l� ��^%j�����+)�Č ~F�Y'�Ck�u���,�B'1����q��:Z�|��ꠣ��6��I�iLEcQ�3^Tɘ�j
�Dou��(Wu�1��ƥS��V�o ��2Pߘ�f��w �� �(ކ�{����`3�xJPt�`��|t~!�wbB�����AfTbT�X����?݃��(�X@�VԸ�������g��lE��2 �2���u�+����8�c�����8Yvh�AF��x��>p�N�}��"Ԑ����Uy��2�{ Q�$�pO�T�Fy2���ʭ+�j�6���ˊ\ˑ�ǥ���披z������W����~��]�=�DZ�{n��I#DnP��/<�:�4�A�.J���,]>-UDH4)K)_m�e\�+�5\��m�ǃ(q>�p&���h��xg���
�y�����P� YHt�@ыx����9D��+8Z"@FCN�rI�\e���r"ǿ �N˓#�J�x�d��6>��J�C�ǐ7��*Z�y2Բ�q/[ ��RҬxn��l��.I|ݵ��o�3��	@O]V@h�;�������L�r�V�;c�?4̚A!W� ���ND$X1UP �;���A1p��A{�x�p2�W.�5�R�l$w���֠�Uwb�;?�{�U�2pħ�N,Av�SC��D[�o��S�G���� �$�LD}��_���/0�U�"�� gdYs��'c��O�; ]V?�\�+�������&*�(E#���ۻ#�v�R7�k��i=;;2�/�̘�jQ%-��%��y~�m��ӗzc%"��|b�"��"r&��G.�8U�-�ub��JM�V���|u���l�9������������SEA�����J���_�=�<,+"��J��״� ��QC_$<#������Ŀ��9���xtX���ܕ�.���h[!i���*ّ�b5d�����Þ$ۚ��EpWZ�~Cu��PZAdM�M�g[#�<�8G�	b?����6��_"������a4��l�\�).4��WE���"�������C0ei���-�׹T�����im`5��L���hȌ\},�O��y����A�n͜?g-����^#X�ۋ�{Iт���~^�hk>�H�����X-+�]"�RH��b;疿(��E	ŉ�#���6�^V+�}@�v#%[�;��3X�4�o����x������i�<C�����ϝT��f�>�F�J�L�jx��	}�S�6�6�^�O���R)L�x����yg ��l_�H����y�_�,#)�^C~�)[N���aʩѶ����T��\�V����kHZ�߯8����͊�;t	�մ���Ǩ���6ԣ�AW���&ɀ��ZRƸ�)���	�Y���ej�ZrgĪ\u�$��i�Uֈ��q~��1v�����zZ��/�Vt�}�aUpf�k2���	��](���ئ�~.}���e��CR�؀���f�9�g��U��c���������	<���/=�y�`�������TU9�z�Ͽ �dT��T溧�c�@S~ǜ}-�u�4b��Đ�A�kK��*v���M0�lLѭ�@�C����y���ĚH�8[h��8��|͍@�Lf7��Z����$�MZ(��ls��h�q�}�=�ߌ�0>Q�8zı�K�v��{{�`�/�e�-m���zN��^����'�p�L�NDyN��ި�t�te�����VZ�~�i	����Mc�߳���2O�yz��7{�p�&�3��V~�l� ą�S]/c��0�*{e�ؽ쫎V��`?:�L�f�v�=ɿU��o_�h�D,�9�X�A�a�Pvt��7KV/�ΰ��^�	�t$���g��Id��[{P�]HNq�V�s�Ç��H�?�7�<���	wTꭀ�H�7S�F̖l��:��� ��ё$S�9�c��A�ħғL�H����'������d�ţ& �TX*���Q����0+�R�i<#��3�9�t�	���Y�g�F�xPT\�"S���b��~*Ep>6M��	J\|K�N��<��,�>���'�Xl֣(���LZ���{)�~�=+�vQ��Ɋ%l��Ԓ��c�����>�]\zW���\Z��hϓ
7���hDE�i���z��O�iTD�"oTˑ���n��:є[pв{<I-0��'�R:8��T��%��UƦ���5���2�A��(���
�-��qOP���31�!��9�BP�	��M6mb,���܆9�#�Jp���a��*v�Y7���mo�mI���$&����|�T[��e�Ë\���b5yatV'�1+DY�G%UD�ɸB�J��%���ΓE}���Q(�M�?+����/`U 3�ŢR�$�-�\��ɡ��C,Q���>�h�8Y���rR
ι�+�~Lˑ��1�E��ك5���'�I��,�:�̭n�����<���Ŋ��h��Q��%�J�&iM�Vp��'�a��#Si��Ll�����ji	�>�UN/��(ܙ�1�;Z�I�0}�?K��L�Ū��g��ؓ�B�\��Z��M��W)9S `L�|�؇ٺ7U��qEE �k
l,���2�{�0��*�MM�񐬐H��,aV��^�7J`ɴDɟO�'�($�� >�Ws���(�1츂^)���?jB��@�Qau��k0�6:�~Z
~�ah��^��c?���Ҋ�����:]�{u�7����54Ը�+��f�j�@Ҿ���)>c���d%\��� �	3��p���9���"�2?Mu"��.'8��"���H;�<ԏi�*���_W�Fx��fj�k�� 6���Һ ����K2|b�K��Ɉ!w�\�}z�?��T���~0��ǌ�Ι�/\�>�}�$O> ��3}���:��߾/�N�b[�	��$����x���(��X_DY��|�/�^ba*e������)�C�7ۥ�|D6�2"|�v`d��O)D�TB������K�w�{SW���������5���A�upF=��{>�0��da�+�h-��J�=�~L��!��θ72��k�i��;u!�2���~�GӉo��_KA����>^"��m�M[�K���Gwx�����̝Κf��~��������Iڨ�v���G㗨���d���R�
�LݴJ/A����#<ug��)��	l����{���M�����)���q\�r�,+����zSe��K� Z�رd��>6h%VW+y��߃����
�%'F��𖫙{�]���>xyX�t�?�J?t��@�,h1:��ԯ:P�f���t���c���L�տzgq$�	N���#��%�Scͭ�'Ŏ[���¹C�bF,	�.$��a����1�d��Յ��w�p�&%	���ަ�Lf�Y}�yi���v���]ui��#���|Y����}%p�ٯ��}k���Ș0K� �Ky�B�x������>ZG@�l%	�*�����D�j�G�}�l�Ѫ�,���"�b����D��R(_A8iu���3��΋�TI�J�׍��?6�5�`V`��<}�-��Ti+�:n,�0���ZUT���y����ۗ4��%�=��>Jt��,�(�XV���C��5�#a\��b�r�1;C���U��	aU!���an���nj��[P���b�dq�5���1��|�� H7G w�p0�F�x�I�)�tF_�O���B"� �Eا�f���ȳ6 �M*�\��º�I�l��;����P��?ඛ0s�:@J��.�B;��|S�L?tb�3�']<]��i:��S������B�́Lũb�Dy?D�}<BZ���iX(5~�v��F���o&��k`J6�=��O�4�P�@́%�.��ߤ1���ɇ<�{&U�D^ҋ��h���_�-���b����=�nA�Щ���Z׽��Wi:����TͶg�/�
�1�)��e�g�
�Q0�����Y4TI�D�o�2S�_����3�9F��Rܿ�k�#g���2�E��ټ���M�X%*��5�;�t�9��VvU��]�� �DA�v��ZK�A��t�-��:�`��)p�P�R>�C~'ʹ�.���{
����ȺlE˴�t2K�1Oa����D��� b(+��dB��0]p�_�9/��b\�+p��V�4t.�=��觛��v7H�lq�,��Glng�FA�ë�E���|�0v|�rA:��3A!��ŵ��v��DJ^�PJ'�3�Uk{�K�g�#��l�]���Ȁ�ntmX
��g��F }�6�Mv��� �.\mc�U|��<&�?8�����
�a�[���1;1rڎ 8QXa�ߧ-����{N7�j�a�ճ�Y뗔@����1�	��z2u�r�ç:6i�uo�@�pu���4AfS��LG��z_?`���!Ϯ�FRAf#j�a����ޢ-)�cr�M��ٿ�~H�l�e��P�c�0l�0[�fmQ�������biJ6~�k��b�m�B�,�?=]�.��q��gw�7cA��GG��xH���9_��lD�Ǜ�#� ���4�-�pQ��w'�"R�߽���f��(��8pe?yh��c��oXm��3B��V�p ��.9ڒ�?���&p�l�^&�Q�'����p�y ?��0�_�q�+�Vi��|�2�.��9�Q_@-̂�[�����`� ���� 3�?�<�H����\ҹ�B�P��>v�qf��BV�~M�:�^�fȝ�A��:�&����9�%���R����5Qgv>�o�[��u�Hs#*���%��A���y�������~�=�w�����<g�����P��b�}-���J�N%����}��\�q�HPx��&��'/4�P�~ >�W+�Z���:�m�4E��
�L��*i��%{��U�^��O�/��I��!�,�ug��8n2�b��P~#
�΄����i�bL�u�������B
S/���%5F3[@�o^��O�Ưi�ڥ��d0'O�T"�FDZ\��c2����\f1��gkn0��{�0�a~��q#"���g��@��.`���p��+��P&�$h7�rD[�Q�N@�l�[�(U ���e��Յa�����l�	,�V�[.�EV�?����X>�B��񫂇����7����~:�L���qEҬA�C���Ri4Y���*Ĭք�L(1�������Zǝt{.JŶ�t5)?P����I�g����U}�^^��V��yά�L�GCu*����[R� �����+�������|f��H'�{���2��>�����X�6��v�zjf�%%���Z1�w7wӂ_EI����[aƋQ~K�0Ц�bm�|l77�6��H�����&o2k��F,��?i��)��%.�ʎj��v�Nf��>�����+a�f�(`_�ﱃΐ���Ǎ�-����������c�H�9�{��슡L�|��3]u��Y{�I�(�_�`��ak����Oŉ��^:$�YZ��8����
�'�'-�{�ĠtkD�H�C��C{�FL�1���S.u3��
8�� 𰷥�� �,5"l_�ٽN�ϐ/�ڽ��e���*P���P���/�6ie�xxͶL��LnE�[�/F�c����
��'#�ڛt��J��eܙ��fY-�Pw���.z���k���X���.�l�>���#s�lۙ�5m�e��}mT�q�ŉ�kV�FkҰ*�ĸ2v<r����/�Ɛf�8H1����&O'�t�6�6�1Q,K%4����5���K[z�KO�l��Ć�٦5�-_�,:Ֆ�Az�1ANn�kqKvp��WY\�3{�.w����p?>z.,�Xh}��2�Ma�*;�t��$�|Ѻ;������Lէ���)CP��kL�Wg�]qa'{�J��,���̺���a��&�"������%��X>��e��q�Gc�s�~�D:��\���:�w<�?9f7�1�d�KV�h��v�N�p�P�BONo���?��π4C�h=5F����{ז1|��k��9��{�f��~�[R�!�Z.c�ip�1K����3�Ԃ����r�	3��԰Ģ�\+V�	n~F~�3�a�Y��B=F��}����V=DO�����.D̰;'��UO	 ���d���>�4��6����V����.��TɒU���_F�OnR�b�
��/��JR�b���(�Yt���(#F�nh��+��5*˪�msy��N��6"պ���zG�
-�O�ҫ�����@4�@=��YxfK5��ܚ~��ܱ	�y�O@�c~��A<�{�FN_'M�b�Y &���(Dv&�&�5�e�J���RRsI��>O<�ٖ��|���Xq5,�P�p<�k���&}�"2��MC�y��ȇ�]��m�ܘȷg �<�|daBk#E=Нr��(v�|5�K^z�g���(���������h�0�՘W�Rx��:�����>���� c�m0��x��fPj^�ĉ�崵`p�b�K�fN:�-�&�M�V�[(
�,�R�Y�U6up�	�EU��h��wGA� W'^F�>����Y,�4@�ߔҦ���\X�ѐ��['�ϔ��mN�E1�o��1����N�])����ךY�[s�,��-�����~z�����Kq�6��(~Ɯ�C��g�g]�ӌ�c�;�OM���?9�r
׫�@�y��u�XEp���>�[R��T7��s�uΘ�L�@�AR�1kmU���~�A�=d7�)y�A��]sjƖ�|��`��K��FH�h}������9vZx��<�頩�,D�ňŴ`��R{���+��z(�e�L�~R:97���$����	*�$�����0�{{{D}a}9s*�;����|M���=]^5�)�����@�Ì�k.�@�N1�BP��F���^��/!��J-��>��{)1`E, ��ȐnLiVq�I�A��0V�K�h(�IV<�.G*�����.FC��i�,/�+e��-߾gy��������5R���K�-��-���_�!��ۚȷ4�|.�1E;�>�E�;␄��-c��㵝�u��)Y�|��Q���6�߳!�[�Ӧ����̂O8R�	/�*��s�\�Z�����1)�����^_�M9��q��M��k���I��k�CH1�z�E�c�p9IJؕ��;�{>gd,�� ]��aP�}C�Ds�n����^��t1�$t�YY1�J�e��ݼ�����Uا߇=B! ʷ#��v��u.�h��(��:Yy ^J������}/���a��'�1�pHwv��<{����8$(�eQZ|䭛X���'�K573�G�*꟤�`���ɾB�w,C��NPR��bL��0�d~��S��Y6�y!�oa������%�������f�����sVY2��
ɰXw�@2Ki���MNJ؉��l��t�X�*@�P5TTz��uyA$�[9Kz�[����'�J!�k�F50��Y��DL��ǗˢJ�YB{MR�j,yQ�icU\�W��I��W�t�N��"<DP3
Ň��ewRv�� �� ��p��-���%r�3=1������{Yc��Y�)��C�N�i� `uH9j,AL�~��F銋���ކ�fϷO�%�p���`�ϊt�Q�ъ���\'Qj��r-���/���"�`}s2(^�Z��R��.�X��:I�8(������3��0F&��A�V$� y���9$�P}s�-O�ж�5ʄ��Hэ�������V;���	_�0��.B�UZ��b������E�h -J �Ka�ȍ�i�nΫ�xM��^x�o�:�6~t}�q7���*T:��z+���|���V8�VV�gY%4v�_7���r0��o+�v�A�b�H{n6Z�*'��!�=�[��ێ�3�@z�zocF�K���
;9?=y�q��
:p���I~6���E�#%ݳR:l���9��i;R<w<�@���i쫍�����K�@�4qt�`Ȍ���\�ׇ&�t� ��[��rs�W:'�KQoz��g�I�H�ySҐO�l<���Vh�������V���8>��R�-��]@�z���C�h)�v�}�^Z�!�AX1�=s��R�[Ref�p=���=�jdX����q�TUO~Ѧ���_C��H1T��"ҳ3��?�Pz����>�O���m�bM��y:�s�,�gC�u�9VU��	��pU��K�w��.K���_I葁��}奡:�ei��TX��Gש2���Q���4R�~�«�[�?��W@he%tJ���V��3^S����Γ���k��"��8t�$�ӫ�A}�sYM?\4i�';�$WZ!͍�*�?�#"�{9�Fs��X��F���ܙS� ��د��&�˂2� �R�ϞS���Z.~iy���"��O<"ǻ��7�+��s�
�����d���w�v<	���;��z/\�n(g��e,4�ʢ���b�Z���g5�ʑH�PRc}P aG�(}��$"�y�U�u��e�h�`О�N�h��������G.���%�9�Pb�"\�%$���ÈV��T���� v�q&�Sl �>�Ʈ��w.�����iod�I}y[D�2vt����Ȑ|��crь�m�?<D�`�<�Iف�c���-��=M
�~��*��x����:[�]�O�s$�w� Р)(�Cr��z���ܟ`T}Ȉi�߳���A��e�=S�X���SV9�^�?VO���(i��C�r{ɟ	u����O<�Bɐ u;�����	&#�<h����&��( �	 ���sJ˗}� q<�����N�w�n�c�����3dϓP�jԧ�V������
d��9���^���x,R«B��mk7�$�&�EAX�����M.� �;>P�iN�S�yg��Z˟c�ӵ-}V��	RF���{��*���q�ܮ����8��YGc�Eu�-��qn��%0Zs�;��wػ(Q��]���-C$j�*<]��ӷ�,�j?�>
�܆:��0a=WZ��y�7;�/�g��P}g��'.AZ��k	�����Cҥ��&}gy����	�������dI��7�P}����.�UU�����::(�@u��K4�K�PA_ߦ�6I�CBW��fjb�Z����a�'!����?��L�%(���$c��p+D��
��N���)�rΎC�D���+��z��[m�:	I�d�n���Iȹ�~K�ޖ�if��M�I���9����.EP	z��_��C�[�n�bTf���u���ح�d~��Bp���31���>.�&�7m�0C�e��i�jYy�eȾ?�p<z|mڞy�(�B��la��0:���P;� 3I���sZ&��/�:\�ܘؼ�}�m�&���� �a�{�		�l�w9��\N���տT�^��+
���,w��jp�ƾ�dp� ,���s��<�ߎ?� �h�FV4dQ"u���&�٫� \C����C��R��~稝dm�R���V�d��3wT����U���霾sq��C�C�+2��'�5��P�BF �!,��Ci�f��$/������Q.ڡ
�
�qe��	sE�)��V�iAׄ5M��ˌ2)EC�w[�;��e͵T�!�Z73��i̵��I������T7�ј>�����;�[C�$�7SL��
HT&C�}u�Ҏ�H5ΙaZ�B���,/<��dŴZ�Rv惮�R<%���l�B�̩l����IZ��0Gº���3ɵ�5����������5���()65@�f^}PEBL��ϺM~� �)X�:�;{��^�nrp�)����Ӯ�B�Gyɚ�!�n�Fi>�VsV ��P�������W�0x;"'�E��k����<-�{Y������6�-��$����6������!O��d��A�A�
��;p9�<���� �i��������O�Ǳ]��&�v����9_7�:�%�)S���pT�^o])zu��ɑ�ߧ	�M9�L'�kW$i��u[�}J�����6X�~�1mK,J#p2tUr� $�Y<��47yp��|��u=�0���+v��̻����Y���#��c�11��oL��Df�+�CFE'�ҢrAե짔�XZ�p�HZݱ�˸�8�o�x+B7Q���3N>�V��K@�2�;���ޕӝݫqT��I�W'��'���US =÷⤾62�5b��a_1H�d偛���:�b�	��s�U����RT���Lb]�Ds8�>�76jg8�o9D��D����/��͏��׭��P�^�0�KVjG��P��qef,���Xr1�}躩�d�����%`�o���:�ӯ�s��쳬rPsZ$�2�,��c�h��>������E�~�k-���M�q��R��mx)�9;��e�c���<17�3Gr��.�>��F�c�w2x�@�V�����;�'$��j�&��a��\L�@!E�QJb}E�r32���Uz��1��������8��27� ��GW�=�&����DZKm��%z���Ա��c �v?	i�$�3���9p-4��*�w�C!<(R6�UQ��������i0WT1ψ�{�B�����0��(pOʦ����a��brQi�x�������m�>��οh�͑��T;���O����ZƏ��̋�=���@Y�to��ۜ��3�H���63�.�<�l{2��f��N}�~|����n�O?��A\�Ȗ܀f��ҳL�|Ԁ�M㝵������5$KʥB7�?��
t��r)W�����XΦ�����T�٦0�l�����c5B5%���u�rˇ�)v�@u㵸:9Vۅ���IZqb+��_��4�t�y����>Bh�������)�F!������/����p	�����ş]�سa�@���������]>%�!�q���.�H֤fp$-�~�J�@}�(K�e�8	Nw�'��'��.�'X��d�y����=�6�!��zbY�g�-��ѝ�f������>v�y��}�&���$�)Ul�!��Ab\C7�kkV`כü�O!;p��cz7�=��I��H����nY��VZ���&>�����@ ϧ��Y��B2s�w|=]:����ӡP���;��E�{ʛ�1���I���8Y�K+����X^��k�j�S����T�o�w8>H�v��H��5�9����x}y�$=����E5�|z� 8�+y���M�q���6�\n%az���yc�mH��b��)'�+��f��x�|��xl���S(�2�7�0��xa����P]�
uZp����$��NQ�}��Q�ʺ�\�а�
�9 �({1�)�����4{�_M>�U�ܖ�}]F'���S`x��-��C�fE߾�9>�H�+�j���3#�����AR�����x"���z����[̺�[��#̔qhHkTP�K��0r��y�=hX�bPβ�uR��> ��(hc��>���̖��(� =�]��U,gBb΀���H�C� ��a|�� !ijX���w����_rC��50&R�)5���a�#�w����b�y����&鱏��wԚ1�DcjQ/������BaTv�,����r�X�� ����� ?�^�lf�_II�'Ҏ�p�����G�Iu�r����͚~��6;�8�U�=��0�P��]C�_݌��f%u�m�Vg�bE�@]��"e�	�Z[b���������Q4�8���� �� �y�1�w���^�k�Y�I	��4$1M�Kc��Cv�;R.�1��6�uP&�j�!�ؿb��MG�{"����
�<��p|+FP�`�y?���O��9j��FKv���ћ6�cN��7:=5��2��H͝��L��D�!��vS��A�rq�i�Ã�#�Qm�2JZ� ]��-�N�~��AVā��B�߈�e�#饀W��E�zz�O�ȵ-���Ֆ���@!_�٦���^������e}A�ut���\�,���M�&G	t��H�Y��A��F�F"��A���Q@�tM��o��3a���V�������9tQ��}r�	F�)?���kA���c;�I}G�#��#�A�w�u?�<���?B�x5�6mgB�*4*U�f	'y'Gj�'ZXs��\H�Ii&$?�!���J��V����y��٥�S����{. t��i��C�F
+��A�j�P�����?FՕ��<$�!=�/���B����O�b�[��]5q5O(��G�N=޴����ht}�q�Kx�q�
x{����uRΉ�w�����ê�ޖ(<`���������1�ER3&�iV�dt@�l�Eo�s�B;rix��|4� z��Ai.�t�$ܩ�D���Z����tJ�/�g��
Q��X<tD�=����v��6����=Bd�<S��-ݍ�҈�]�7޹���͇@W�c��*_��|ãN�D�H����Ev��A���8@"#lN����wN�4ދa�f���ʂ_�-��+�f��Tz����a.�`�<��&Zb<���l�J���}b��>u�n��Yӭ�9��:�1*�y�D$�b�Է��c���"�TW�,!�G���z�i��!���=���Ce�p֧��EΧ�����s�����0d=��<�����:\'泇<%y��xK�Ш2���q�q�IZ�7��$C�@Z��ҎG�G��3�~5��8�\N{�:�N�I޶m=��I������&��(|�B[|�_���a��S��6[W��`!
ejnP��^I�Ҁo���d��k4�U�|�xdM�p�"4���
0 ��EQ�N��+���g����Oy(`UB�K�6SPd�tb��*��uE��yt`;�^-?���q�7��Շ��&������FA����h����ȶ$�ƶ/�'�*�F��K�ʍ�E�>��UPRjT� K�-C�����VH}�+�n��,
[-^�v��bd��W}�g"D=-;p�.[+�SFX|K��w���{)�ݬ7�� Aa�~ӎ�^��;
锐ƪ7�5r����z��d~D�DoD�а��eDX�fr/@3st�
CD��U� ��*�6���mq|L�mRI�Q��oQT^��)� �A��#���&�(�<$?�Q�$��C���h�~C2�u!MTLy��8n�$��J�hfs0>�Z�Y w8����B���
��;���.U��L��׮�#��C�j�c>�q%���ñu!���2G�������1�l�O�	3L˖��\J�$+誺�l#1!���^�x_9���Ӣ����K�]���R"^<&-�9õ��V�T2����Y*�Fԟ��U
���0�{R��%��m-�<vR�-��[I�i�є�1�Bٛ��-vnK;^wR����8�g����6�}�����j�CO���Wj�;d�FU��n����6�ى�1{B��U�[�ͧ�<3�QX���m*?x=q��+	n�ɔ@�*�����E�n�T�p�z�b-�&3���]����|޼�6�{���D>�b�m-�N+��	�y��P@(��ZP��b3!�V�i�6
K�Nݒ����
�X���4�5�Hyn^}թy�P�.��pyJ�ǰ�7�̻��N�FU.c+0�ˊ;�Q��
&li|�VU�'��&嫺GK.U8�9�O��8�{��+�
)�ې��q�y� k6�
��J|��(jq��EA~����ћ�	��դ��ۏ~��밦�d�78�%����Enb�(�����a�yN �����x�����T�1��<�򃄴2#�����pF�w��}@OC㔪�+��ۙ�_�ET�����]S���N*]��n] �p��]EH�l��.W1���ŋ�_?zG��A��{�s����]X��&#!�3S�qv���3AH��9|�p�����5;��bf|���ƞ)(w�J�i{��@�r-���c�x���uU��R��z��B8�y|٣�v�l�� m����7��;q�	@ S��*m�u�����Ӽ�����>�U�v�ߕ��L�2k�e}*֙e��?���AfA�aZ�۱g�V�Q4��`zh2e_���f���-{c$b+���A�?R�{�9l`�s�����k��?�^ ��+�+�`�0�����5�	 ~�v>���њ����o����E�2ՍFa���(E�^�����˱���%��zCő���9�!kbF�S[��VP����y ���K�!���o�;������c�`ϓ��sj�GO���
��N�b�r}�`�k���!� �b�Z,j}�d��������:�+`�h@mi$EƝUa�Xa������'F��ֶ��F���Q�i��~ؓJ�9:�m�:�0�?�1�tT�q� �ͫ5f����T��+]�hJSkO'�s����C����g�a�Z����=w`�|�쟂����Z��^�~ů��������Cx{�6���G�X���;����j�G�!����T��κ1D�+zil�唜=Z�4��'lV�dʒ�H��s��ޮ���thmd:���tO
q:� ��� ���x�Sv�^t�8L�S�x�X�T�Ӿ{��b��'K̙SO��$�a.�H�J�����v�oxl!)-cT�mzX��9xnq]���H6�	�H���wLm<	)T\E�"l�g�t�RYP��n[z�]+�P��ń����f��>�R���b�n�/��89����|����yz�*N>�{���m�b�Z�����ϑ�����C�?���ӧ�&iN~��yG��N��J����tZ��]e&�	�|&�mm�ǑƘT���#�K�#�7"�R�4`���6od����R��i�I��/��u0�oV%����	�G�F��	�Ů�׮�
���Ǐ��00aa�XIЛi*h ��v0*�II��~���_K���	T��
]��[M�e�ȷ�xSG3ac�pn@�Y&y���5>�f`����B�������h{���G��ొ�M�AH�̧��颱T�^7$����gXˤ�Q esg�)� s&d�bwBJ&ww�-�11_�ϴ���Bζ���@)�!�ˬ�G�_};˷s(�fN?O0Y�
>�׷���h!t4H#li��AçO�S�;ߤ��1��^�4�ٌ�ցV�Oz�Lݡ��R��a�er40��������%�`�"d:,�"C,n_x���������N��n4pK����� "V��w
��	��3"��z=����ף���v�w�wa�ȴ�E�(������N����ஶ��' ;-����hlQV�י/QT�4�/òH ��@n�8R%���u�ᆁ�j;�ӿ�P�|���7b@��cD�lMq�OX�I�eJ�����vM4�~	��f"N��4��w��~7��$.W��D!#�H���]��JѓF^�r�7;8��A����P���_�r���#��RJ���ׂ�J R�˥6����,#�	t^;_����u"�	�BU/�p�.86̗|.��!O8O��H4��5�y�ڣ����_ڢ��dzl���*�)��4��N�AQdHҬ�y�-`��4Gu\,{\�:w44,��nY8�A���
�bQ;'�_�8ҽ{	�T��w�h��؊�{i�M�v ��Ws ʚs��G�	�Ǘ$�k����xhU6��O�[��f�RtpEb0��`<ҿ���T;概�cI���ǃ�YP�+5E���c+��ta�X��'�^Y��8�Z��71�������C[2V��G)ř�ε�[����d�xõ혛p���mR���eX3���F�D�c�d{*�-�Y=�^`STͤ��CW�_���R<j˘+E�:zd�I�!�A��a·�z0U�RA�Yzn ��diy��l�O����Y��~ל/��7�ƶdP���}�#o\=cauf��j����k(����PY�6�\���Ìr�����A���˿~���N���}�48�@����k 
�@�|ϛ+��Z�zv-�RA��������:�%8�`����>=2/���5��-�k$c�0�����&p�fG`�َV5�Kݽ��	Z밌�h{x7��9�d:��Ҧ�2E�o�e� x�i�!�bp����!�!:
^���gy���	�!��N�h��B	�M3z� IT�0�`(�(~��pV�Ps@Rʘ��l�3[�*i$�Uo�������Qe�|�Y� ?���"#,U󿋚 ��\�{a�7�O��H[O���6�P�Wk�o�\�#꺹6���XQ���x0������l,i�n^G������R%:	��1�#������W_̌�)3f�Ĭ��,�*���mɋ�ݷ����>\���� .���g���Gu�>e����x	�;b�d�4Ei�m=����рz/����ږ�,����I-�U&p'�3����*
�����Ȏ�S�e�VU��T�I�/8�ǖЭv��N����������q��5��<zE(��ܹ,�ck^���/�Ov�i��3�u���U��	U�R�A6��n�r�A<�a)�hC��^\��L�=�|h��i���*��s�,��
��q?_�M���E�S�ӘL��`z�<��a��C�<��-���zV�x0Ǵ0��TGC��^}�Qx�[ic>Fd�&�����C�Z#�EǥC|�J���Dda��R���Ν
���z� `����c���Jѵ"Y@e%wr2��hTY�Ժ�5��Eb�c����$��%d#J���j�y���;���4a��ጢ�oķ������bT���?�^�?I�O� V�sI���F����dR����òw���.�}��X��	�}�/�G�^ܖ:����x&�- h��c��?��[=~��N�!@S� VN&C�1 �"�8�d�"�l/�dбV�WT'xq������-7�DX�/q���Fц��ԕ���v}͵���|j_�#Az{����W�FXY�/}���fH�s�D<��γ}��藊WY!=NOWy�K����X�K�z�Q'�.q\:J�J�}J{�ZJ�2���wOfX�2$��ѯH��M�sXSQ�y�'�0B�=��P6����L�K7+W��ܟ��U�(��*#�v"�(��l��P��`%��I}%Ȓ��<�~�x�\��5�_~Ss6�:���]xHV���v�;_�I�e��f�f'���>�l�v�3��ܨ��o�ג�W�ac��a6��Z]M�P��qR>h�׮/u�Q��P���ꙍ@�7��srAM�������u�q�N)��r�C�ėWV�?l���­���UT��<p���5�B���$�Vo� ��9�I�A��Hݲ钍!�=������$i���Y�hCd���ȿ胆�K��t����*�Y}�\�#���D�J�|��M��֗C�1�bt(�u����I�0�A��Ris���=����+�L�?r�fp�慫`��/�~\�GB?�k��V)�ۓE' ts+�e��Ct�#HV﯉���p�}�Rԡ��Ο/��r}��A�ڟ�v���r�F�m�=m{'$���o� (��m5�$=�V:���c�4��is,E�ruq�����؋ﬞ�B�4�$�	��V������^竈�W�[ے5T� �9q��_qƋ��z]��FN�I?oZ'�"{�RC6V/�돈�
x�V����]�5L�Y�'�3���/���������@V��e=�g�: ֡�� �g���ݙ�n.u|�
=4��#`|�D��-�[7aK��R�,-�))�jձ˨P�_�^�営��&� ����A�?2��ǀ�����<+&A�]��+�>
�K`[�I�4�+,�΍���e�b?-�1I�2m�fd�%w�$r��ɤrZ�Nƀ�YsO�V���3cΉ�	�S�K��E�`wT~��sV��a$�?5H���n�ϯe_��+�|
mڳ�m܄J��ۣl�4�&�3f���|���.G��͑U��������|����/�[�lº[�< �n�\��~�s)`��n#S�?/�A�L��9����C��;ꑂ�fe��O>e"���R�Lo�+&�?�і DZ_W��$�Ӭ�k$6�pͥ�{�+D+�w���
�V�u��6v �/-&jpz��;_6+������|W��-���Y��I�"��x�j��dB���D'����l<�g��A'�J������������������J~�ğ@ �k9.���.���|	Č��sb��� �vz�o4�FNAZ7�\�8���$���lD�F�iW�6��P�K�&'�jib�#�,+AO|��K���D����58J��ـ7��L�������P���~���O��aw��	��@�(��'j�ZOO2�v�r�Q�!�}*���'�؈��J�ʝ-�[q��t�Hx��6U�w�~�f��TWN,�<��L_�����
z��Vځ�%F�]����.A�4ٵ����\���ִ%�E}��2��e�a��Ār��_�Uo`��֗�ꦑޗUow������k��+�I�,O��������u�S�z�ڀ�R�AU��ݜ1B���ALl����F��I-6d�Ñ�B�$�u4�<�'6�i;�Ԓyeӊ����$�jlaJ��;ۣ5�{�>N�{Jun�[_�d@ �&��_��8�����$�74���"N��X��& ��~C���Ȏ:�I�������~
)h�(����\��,9�k��� �S	-Jd �X�z���-f$�E?��,+��3��}�v��]��)Є��!EQ`&ɡ��hx�΃hI�ӷ�QV�]�`+�5h�B�j���ǏW�Qf�=�����3�lZc�LG�!a9���(B'ɍm |e��z��R�ǁ��0Ϻ�|���f�N٫�7��,Z�)R��j|nÌ!�lB��Y��q���P��RJ��M�Oz�ȭ����[s�F�kӐ*�{��=I��mt�<�ǹ��;5������=�9�M�һ��ջ�!8��<
=]J<�|7"����'7ǥlD)��~��f8ƛ����gk"��՝��e�v+!#�������i{�c,�8�n���g�}�����":����E�K���e����5�w�oX�|�+�˦<��@Ja*W-�K?�0�� Vu*���jwa�M�f��@BtMO�4��
(%����h�����)�J���|���{�*��!rj�X�Gk�G�:}T�|�-�<\]�q�_-�;彫_?�J�o"f�@����`ձ-uQc̵/gL��B��l[���$~o߫qZ	T�*���v�{F'�v�9y'2[�|uS��W�؋��?�Ld���P��5_pM��[4!���m>�׏6�$��N��C�8����56n�$����b�<��J�&:0��s����:W4��B�v����!p��m�˪�t�'�U0�M�yظJ)R�CV�(����):l�{T�nv��^U�Ř��h2�t��� ��j%��x�@�?�$b-k������ra�V}"Y�(C�p�z�����]�I2��ݱ�d��8<�@v��)|�ey�Gt���O��E�UW��p@[j�+�D�7��R?u)PK^മ{��b��^�j������tN�ң�����@SJ�+�=[����ύse�|�����h��B��*�x���nS�k�+H�;�-m:9{CC~�u�-;���i_Gњ{g�s"i�\�'��D{����cC�悁crwTE��'z�~,�"�MM�;H���NX���}��o{Fk���O\^�Ox���*��a^��Z��3������������&�
�]W���&D���R��('ddǼl��^����3[�
���v��FPt�����U�;K���a�h��`Wz\qX8�a�d*����7�x��[5b�E��3	���l)l(0jnr2v.ukT�)��⇐4k��1cќ��2��<І	t�,�R�UBf"��Ҩ�~h�(��e�����11��J�[G�
Q�m(t���p!�Z��qQ^8 �c|��f����j�M���������)����ΰ�Qm Λ�֩*�u�Rdk<�H�Hl"Ų�\H�<������u(�T��� �B�x�����ql�p�xQKd���H�숭V&����O�1��ۿN��2#�d=�(��@��x"�H�?�����4b�g��X�(l�+�������%Շv�}��J�xt�4=^�3����q��ɢ��x�	�	-�dc�nm��k�@x"���@<h�T�ތ w���*7w�Z�g}��v�a-l���ܙ���x���օ�3qJeC���nJ 䭽
rwn0�\TŎ�Kv���+���C��$O�F����2s��rD2�C����C��⸏;��{�3J���)�3��A`}w�i�Î�:fC�M�e~GVz��a���BiAel�%��NM�h�P����$������Q����m��1z�D�����)�����>�+p��R��!���d��sw���B8l�3ӱy�p�Z��yۋ�X ���=N*�X�8uVr�LZ�M329�N!�6Ù0?���~-_�pHJM4V�?Bn��Z��
���T�BƝ���^%�wx�o���:,T�=�E@a���r�[��bE'�x�X���L�tQ���~�F}�P.��v8���?�.9�;Z]�kUݞ�OQ(�QQ���*)��	yfyĈ����J��2s��RԼ�������jꗧY��O�zi���"�����'�w�� ���;��\��0�L���		:_��\Iߠℹ���Փ�+4#u[(���#j����p(�ϮcY}�7��e�om��"%},�Q^ˌ��:�\"[�	�䥂a E>�W�{ᴕ�
���z�{�C"#杙�p��[V_��ģ�Z�!��{ߕ��}�3�Jя�kڅ!�o)��P����h��Pw�
נ��̓\�LZ�u�T�>�\�KDG+ݔJA���S�:�������P��	Bo�JN�%`���8.r]4 ���%s&.?{9�a�D7��+�!���EH(�K�y&hi��"7U��{�*eDQA���WJ>��R��c�����"��>�}��'Rɒ��b*���}�CB��!�6�V|lE��C�����h���U��.�ׂ�%����+�]mL��T�m�/�"^1(�lq�0��.�i�W\��#�����9�L0�/�|Of�4ꅲa�MB_��9�1N��;vo�j��+��V��9�!d�pHU}Qkh0��^�{��z�ZT�� <�1.еmX-!<DT�).tæx2���pω���+tu�ͨ^-��N檶�`�Df��zRtR"�޼O�t��B�%!�~��Qzz~tD�<�8���� ������E�*�e�y�R���r�a��r����,���
�6��s�^W�l���FCک'i&p��{�����&�U���$�|c�}|b�2b�
؎.�l��D��7�乥x^
�D�<j���҃&0��>���V35�MxV8���lk�Y����ԇj��bUr�$&ʔ���tW�[�A���CՍ����ƅ�;z���4;몆��O�4���PR�"��ok�uu6��#�mZt��+fi�ۜ|���J`�ӈ;Yؙ�릯K�Tn-,���+���(]���5�]if^	w* �W��
M�˚Z��|���*��W;�k�s�܂�*3d��Y����v�����Q������\<�Ch����E��� �L��wL��㽂�S8���9'�k��#��-P�[C��K�G�7�E;Ei
�Ske`{ƨx��$�H��@��Ɵ��O��f������U������*FTyO��N����u�� g
Q���+���F�D],=���3�*�!18�l�5���Y[���`���h��-Uv�Z�ݗ)h�G� �̅oмŒ}�`��KdH�T���7S������\x�*�����I���W�/�W[��!!񽄮H%̗��/0MA�Y}��|��j%�� 9N�C	�a��^Yޟ�~�y��}���6��^���U0��<�?$�i8��s�� ? ;.iVXXM�^0 X���L��C�1�S1	G'�uѨ��E�f��.�Sf�?�{fϳD%��Y���Q$�S5�$<-�;����m'��4O'�#{�=|��
J��Lh�uJK�i��d����\��*�g��;��|h�G<I��`S�L*�4�8�7�:�h�3n�L������!Y)"��h��|��!8�xŀ�ߙ�|��#��Κ�q>s���_� K�/S����R�]}lm'�1;},~��h�=�2& ���1txڜ^�UB'ܠy��d�!r?��\9�#�W��^�lm �!��r�HqMO�5�N��-8� ���!1��F�E,t�����o[4�W��S��Ēպ(�����5�3s.����P�����{�i��ʷԬ{l��>�S=���E������d�����n�~�a�C��E*mYPi����!���ޒv'Ȩ����]����]{�Bk�L�#����v�C��y���ҳm�l?�\Y=��[>�����!�y��a��OjQ��iA�����Q�NY�g��u+ˆ��TA���/]��]R��\�6�#�7�h�R�<��^���:�Y1���/��N,�j �����j�ӎ�� cd�r_��?Y��V�$�Pt�z�:� �G�����Ď�,{
e 䒋��v���O��	�.!���%��gN����$����.,��pa�d}�{/L�}��n䯒Û���)mO��}�����@dJ�ۃ5���-!x�?��,S2�9_ǘ��nQ���e�U�,MF��A0��9��CD�I��^�]�9����<9U5~����4�Qϭ�#[���Z�T"��OY��{�M��q��)+/��:�9g�Gqr��u���n�p_w�������r�x�G�ʧE9u�?�0~!ɿ0�*3��#}���/��ϔ�&kJBT�������#�ZbC���v��	k��7hZ(�2���T�[�
��/g�PG�ಋ�@hLo���O����j���	/���'f酏�v�Ŏ�QTc�z�{x-��uu��q�����`�, �[��[�7S���Z?�3Ly��qatD�B�,�/+"�<L��Xe�F�M������~����.�<�x۬$Β�F���#��1����)�Y�;{��GN�v|�%����Fv��(�:a\&�F�㲓��ZjŻr�:P������x!��4�sYKx����B�mB�
Uyy�KR'������}�Q��*xy`.a�������ڛs8�e��Un�e����(-P�?�F�z��F+{�Β*����X�}���D��GZ��0�R��k��X�bD�wwag��@ݔT^]o�UI������g���,��w^���Z7���.ǡ�U�?5��^>�9�F�3r(�~*K�OWa�����A��z�I�7��)���|ղg|��Jy�XH^��NSe{Z�-�6�Y�T�X�s����t�H;�Tߑ-�FEJx�8f@�*����>�DM@ޥ��*��iN�)��+�)~�F)���$O��r��6�$���=0�>���;e-d��O�^|I,��I6Z�1�z�uo��	0�aP<��<�N��|��ۿET�E"�nA�X6/e.�.JLq��2SyՁNz��L�7��U�<dxqa��-,�%@x_�c#2� ��)��[W��,1�r&9�Ŋ�gV�<��vCb��=vo��[�@~6��7���R�?����y+����<|R�+���ɯi6�>Ҋ���0��61�|dh�܇�qY��������{��x�UJ���&g �K�����oy����~c��!�*��p`�@.wN�wH~vB�����"���<u�O�=v3̸��} �糾sIY�Zi+X%ꓝ����ĉ�S�����#Z}ZsV�Ѳ�߅Z�=�	)�!2�7���l<�*�s�(@��HE�5��Zf#4�W-��?�v�J�a���$�p_����b�,L�Ӏ��FS���=��?uG���&ڻ&F�`x����w��1ֺ�R��^C7qލ���8�_,����7��j�v9OT�&8@�1�~�}��M~<s�mV�H���}��֏!��
���S����ϐ;�8.��6�����2 u�n��ǔp�K�\.D�$�o�Z�iZ&���&	Q�vt��b*-�����m�O�����\�F�L���#N=1�@#�
�~1�ױ�}��sZ����(֨�ھ��裹��F����~niJ��6�WP�Om=b� \�ڟ���c�~��AmJLKWǼ���z'9he�%<Y�EL�u���9�:�mʺC�k��.o�Ύ�^}�)�4ݯ��Ϧ3j��x�US�/��� �� �q��y��=�{��n�����(���Y��4�ʚۼ�K�0Iu��%pK<I{�'��)�/�8�[��ݮ���A� ���P��4���E�0F�B����Nb��[QFCH%� P�<7ʔ.�q�i<�zsx]�4N�w�_o���7�{�W)���䲦@J�&\<��6�p������+�#&����zYk�O(�)#t�}����IGeYkmr����&b!�~w���(�a�
-W����m�X��|��K+�@Ө�D�xS0����Й��V����\'è���u�kՏU4��@���A��R��3ۓ��CF�\�_�KC���Ï���k���U'F2,6�B����m^�a�tT���5(�(CAlu��D=#���P�"�C5@TQ�f:�`�U.}H�P�y���9�1aP����h���6���[��>��m��6�;9@�m���!3��w�D?6]?��ÕX�mHn�	��|��M����{�݀�+v�!�59�Mh&UI?I��M����@��@ø�՜�N�h7j�٭ �������k�/��?#(��'�?�t+访��|g������L�������M��4�M�~��0�{Y|j�2����heD��D/jʗ@cv���5H_�����-�u�����:�/��5ѽ���ὑT:����j*b��J;���B�dytӒ䯘��8��&udr߄���&l#im��QI��iٛ`��B���V�f�\󑠿�$%�~��
�;c�������6U�N�v��o�4.��Ih�;���I��	}�:�"�_�}�Ǜ�2z�|miJ'�^�Z���R�dgj@AH;aub<��;e��U�v6�^���	e�i�tJ֏�V'}�jc^Lx��Z��㔍'PVRrB���Q.��x�-�/Uԕؠښ��s#O�P��F�=Oi�7P�������W�k�5�F��!�W.p݄fp��L���J���ca7��hƑ��T�6���k��2��nO�pr"Uzz�����i�br���]z��~,Z��ܑ6�op!�&H���3�!46&���
e<���+��?Ft��o�F(�7ZU���L�p(���
���@��ws���B��c�dC�`����k����5ho�����ہ�p�#@ت����s�/�׵�G}*m��R#$?Y𩆁�^���r�T��x9.QܧC�t�*c(�j����T�� ������7�w��h kGJ��u;m�
�[�
��;=�זU��Ǳ�6鉮U�f1�G7�C#�3�#�� 4W�e.u�t?6��q� $�V�eo8�g4n޿�l�����c]>J���gfRa	��:!BX��jO���m�-�dg	f�x8�'Ϩ�GZ�7W����<���5l5�z߅�}LN�p���P�T=�%V��IJ܌d��B&��~v< ��?HX�֎$��xb��.�>�GRu���fl�5.��������GIVB%�#@�J׍4��<u���Oí,���N9��������eT	��O{D噒ɭow�Ʌ��nzfǰ��?t{W/�4�Z����`��D3~��6Ws�ir������)���Z�׼�����Y�\�xIL/��"����Uo�f�P�����h��3�As��0��n�1xܼk���M\ha�k�s��b�>Pꢚ��=6-�>��CgZ^�!D�R����k�$Š� �j=�2��/�>FR8	)j�������?���@�I��f�J�eb�ɐ��b�R���[0��V�������7C�R�;u|&0��@[K�p:��m� �{^b=:����g�]?�̮����P�Q�;n��ձ�N�-�>����������ZsR���÷���z��\P�x�U=X�\�|؟��Uy�����c��S��� ���OM����u�*e����z��d�@$+��ٷ�I�q�"$���U��
�*�vehI�z,f�%gH���Vs�.nr�����3�#Sޫ0w4���I?I{W�d�q���=̶m3� ���L�j&���m��	κ��S��8}^�<�I�1�"X�+0��p��GSu�(N�����~	��gb��n�q1��|c{,�? �4I3��[t����h�dp' �Q���fv8�O^B�v���v{���yn'�)J�ݟ�-?���.
���o�H�
�������SmCԳNd!N,^�'��prLӞ�E�}<�ː�w\�~7���z��V�my�����:<������0�	}D�|5��O]1Gn)�߷�[*��1ȏ��i�zJ���� ï�Ζq���5H��gIU}��$�X�#�0�f�����;h29ik����IiQ��r$2�p��y3>︤�U��v��z�Vkd"�v���ӯ))-�c`C���xә�O���7φ�j�%6|����3�b|���5�����d���?�l�FO�5�����^�<_��/�}v:�|Dy��z��^o;D<�� W��G
�@b����P�u��
g����-��ͪ�������N<`'�ഥ_XNG�${b�Ǉ�E����s4�Eei@�qP��t̺H�FZ�7w�������b�C�9����+�.h�n�� c�*�@aK�
/[�"�������ǭ��
��Q-p4��.���f䝈�6ī�J�" i��Vk8#�9|�U���̮U2�.§������	d&�.̢�'���K=�����z�L��O@��'格q�tŢ6%�s�{({�c=]�T!_/���.�k�@g�-pmmU�tC��њkG=��e<$�ż%����D�A5���.���u���t<�T��̛c#�WD�Y���L&��f	ޜ����+�� XI�k4!���s��1�Cd L�=��Q.�p�S�O���5`�dYb_f-�ͺ�Lx�㣅*��N*HV�.�}]��M�_h��̽Ӥ��J��h��Cr�q6�_�}`����mIO�����I�O�;�P3�5J�E��~�~���m��k&���z���	q�8�Bl�����3�k]���ǴŚX0Bsh���1��H�o��9�d��XOxݓ�5J��5<�8��U�[�f�ǟ�@���5(|�;�` �BrF<�v����M��q9SJ'h��!�2V�Ps|'����s:'HQ>�U{��>�O+0]y���{w�E��$>I��՜9����\��^�x\�h��'�eH��s1t�ꂭ��#щ=w`nj*3�.'9+�8j?-�4�NL�a��y�9��٩�6���6���A�8���EE<F�
nhNw��^n���Pe��Ľ�Q}��!��`�K�\�"��� ����A� �y�|�Z���<�\M�IQ�)�.`�!�Ȧ�(N-/�1�7����h�-�X��+%A������
��g�ӱ�9q����EZ&��t+�#�q�LW-�w�F��]���-���tx�WX���ֿ�!$޵<"v�us�mN}>8c�S����)�E����2�h2@��΁��ttLiЭ�	H�a�$��aZMMT��V����� ��D�D��
�iK�qCƧ�Q���]��kA�����p�9��o����A�4�H?S'#)�J�q�����	�(���¼�S�%�
���$��E���RI�T���5��s��Y��APTBkt]�z���d�BS�"�$�(}Tղ"��Pf�uֶ�ꫥ��=/9�k(WE�d�ٰ��"�UB�L:���.�{������r��SO�9�!\&dx��
�}Uaܢ���y#��YL~��Hp����ߴ%������/�5��-4�#X����?°!��z7�͏#d����۳H���Ų6�k	/&�q�!� ��4��#��IG�5�u\��m���g������Gׂ��2O�5:GY�&y����ne���-m�N���R���F�B02���ί|�!Ǭ�bJ�M
ޑ�k|���g���jw��W���:R<�Na��H͓�-E~(y��Q�Q�&F>w�+b�՗���Q�j�ov�[��.�N��i�#����N+2(��<��	��/�I�KL��^��(�w�sld�WlH��NgV�T������e��inl�¦�Dl�p.��n#�i]��|f=u{O�}"��Ag�k0��Y�yPd{������/&3-���bC�9�P��!�Ҽ���1ࢺ]�V�����=��o��#�� �� ��=<U��>�;SɨY	|�
Ɛ�P������&�|���)�в�LcF�i���i���χ��@���#�k�z8D��Om��K4^aFW������	��͉ȵLX������I��*���®ܢR���Tp���fIXǨ>�	{���3�icP�^K��*0��t��(�R[���.�Z��~zGݜ��%1�͒���Z��aO�̜Q�^�h�-q*~L�#l�����U��v�_�o$��[����l�.� �^�d�U�PH)���Q{��kI���a�SgTu����5ؗ�>�/�7�(M�&����9��P�Ķ?<s�;�ݭ�9!�oP���H����9n��Q���O�u�*�Pɩ:(�^[��Ҵ ��-��A���X\FUT|.�H�
���Fs�&%i����� ��Q�������2�ʣ�i�]F.ߺ[Ϲ��J7����J�n�
g��Μ%=^���{<��	�Pi�D}j^*�o�K>~s��jc���'ͻ�����/�F�^%���.ɂ A�z[��$'~�M������R��Q����(]�&n�{!��'&X��[��P�WE<	$�L��Mh��L��8�}�`��A���;-��<��[m�G��|��P���~^��r�-���O��͋~R���&��$0�w�L55�Ӑ K�]��ڽ�|z��|>i��s�=l�D��ɢ���߂���%����kh�4~�����%��
L�P��,�q���9��ԊS����77�+��g`?��F ����R�9Y����(�B�z��!�!��p��h���t����ԙ�k�{����[
Y�V}5z�:��l��oo&x�!��8�A$�VR�e9��n ��6����S�������f%,����C	x����n��n��z^���ɂ���"�V[6H�������iQ�1��xn�%T	'T�!;�g��0v{َ6FQ�=�d�&���>���/Hzvx�i-������(��:ID���z�Vg�������0J���X(�+%m�\�DU3A�2ח�^+m�����,���.��:>,П�.=�!$����C��6� �ȇ�ʩ��1�C�x[D&ʱ�;��;�\TI�UZњ0����6>���-t ��x�.l��A��$��N/#�f~[��e<_����gj���� u-e Y���>(�`�:ocV���Om�i=�y'E�o��Ɋp��G�s@���j�i�������,֪8��e*�xk�jM���~���>��g��g��W�����˔}[ ��捸agf	�,$�c����X<���1n�u�l'���6��ꎪ���Ny�8�3�D��ED�R򿩁������H�NO��i�`�:��:����L��7����[��C�Z)v���@Gœ��L���-��c?�ŋ	�9O�đ{@����]:�+v��/���2x���Ifm�Ff<)o��-��_��J�S}@+5�Ң͊������ʓ�@�lX����tX�Ch�?����X�n�3)���n鈗JA�y���w4����u{ENkݨd_(��z�R�l�h"%;��]��F.<d�����FX�6�]ca�!�~���z�۔���1g�,�PS����fs�6�m����]�ػwqe�w�i<B ����Z`�0�&@JU&��&^�R��Ue�<~	�7!��g
w�ި٨?�9� ��
F}1�e�|qaG� �$H�2�¹���d���N�
��CRL<�j�a&����H�@П�"��P��>$1�, �z	@;m2H:2��4��)8PLQ>� �z�7�����j�x�|1
��˯G
L�%���.��C���Ase���|��/�yrt�;X#��2�ʊ�P�̌���ԊҖZG`\M���e���kb�_�^�~���d���6v�B�7��k��dA�R�8A�ˌv��<�)`4��9��:��imI��ű�`�*��"7��-Z]����D��:�s-h��$2<ٝV��u>�ID�j���Msv�"A�+]��;�Ƴ�3פп�z��c˴��T�hzT��~�"��(���v>��Į6�5��{f:5q�o$1w��*v���|`׏x��vs3YOZ�f�r�`���C V��˝; .�1�(ӟ�4�(�.�Y@`wJ ���R����cG�!n8��*8����\�|���8���u�$�Xw�PU"��q����B��ӤA^׶�C{kbRL�]����Q�W����b�Ɩq�H�tc�������('��W��:�Cy�4�p^V@�0x����ƙK%�ř���_:���}�c\7�{7�����]V��p��p7�1�/|�!��:����K�U�|䪗��������I��ΈY�N$!F� G�X����)(�GF4a=>���2��<��"��ht�A��}Kŏ6��k>F�/i���_�"�7���)6���Z�K������
Kx=xt�_E�E��.h�%�q����%UAhv�i��#�z��$r�s�v9���lk���1�G��/5X�5��W7P����3:�x�9�hص��w�ɒ�Y��nq0�.QB����@=.�n����a�~����k�C�v������j]�,���DCI2P�=gQ�}R���"z��|>�������i����3=������Y�0��������6s��O���㯌`�]5�T5��@��I.���r��o_l+�H�~��_�Ԣ��-��u?AD�N�3ͨ�(��d���8
�ή
���)���/��"��X�V^��b\Z]�K�܀c��ǯ��j�g;�s�9,C�6f�3� W��ʤ�J�r��B������6�-����\�"��AH#J�=�&��F�ʰ璦X�g�J���|���f��vI-�L�)ʞ�����lZ�¦��И�=8�:/��4�����c��K�/)���b��gP Nv�������ՃoR���OM�j��n��`�ex��˸L��L�5�������C"�q�JA>�S�o��R	�~)�#���`5w��� ���Z�o�&I��{]�~J;�A2�7�o��{�)�q�3�Hو��1��w8�ݟ�ǛщW���/��s��C�7N�U�����N�}Q�OLӯSy
~��"���gG~޲Y�q|�Y\�6�\�	��qO����6� #�%t��0��.�F�~Y���Ӭ�?�8J s�h�"Pv�U�pΒC��\i���u_�[�mbj�՜)��9���.� �gk�W�����y�^�{�wq��9���(�-��A�,§県H����~,�J��ƇX�g�U�B��Ls�1*8:��į�G��U�J�->�/͵�#�A���K;�KxG�� �nf�KY�\?���Oh��nW���͡?�t�c=������L��?�	u�c�]]�+g����(������K�����o�A��^�gM~-S�x{80����@��9?T�BT�"�����hL�l>Kd̗����,�0�������ζ / �@�vT�;�7��-b~`@� �>,��[��/��b.�d*`��C���c�1V���X!�<�ݒ��}�� ��V9�@�w�w�Y���'O������B��񵫚}�5N������\�F�c����Ւ��[s�����v�����ݠ85������)&��8b���'$>Z�H5�P�ã͘���T��3�!zp�"yu�k1p�z��4o��k��"�����DJD��	]&F�gZ�>���)�����խ����Ս4 �.�m>.D�&�����F[�G�ą3��яj���1��\c�-��f��"G��:��$A�x�����0���}����(Ð�A]y3.�'��.[`�~�����1p�C�f���
7�����b��Q��#K��_1�sb���^�Dסh��"�	�s���S���1ga<��8z���$]��zj�7�Ѝq��%�ͻ�E���e��@��~֮������ �UT[�
�O���Z���JN��<�2pe�4c:l�hX[E�t|�	O_A�Oɺ��3.3��c�$I�L�+Z�j��������y2�N% nJ�w�Ng �t�!�����S0�JW�J�7����z�� ��c�2Q��]���:�I�T�CB�s�B��G�j;T�삣���*KUNw���K���^�Nz�Iщ�Vx�$� 0j<3�/�lN�Y-�a*�ȸG�b�DN�}{)��"������)��g4�-R�[��ٜ�wZx�o~�ү��|2ZE��i�S2a�E�2)G��)�m3�\XK�%Uz묑���:�\C(���������g�@�W�502�&��̻��9Q�L����[2�{OS�kl��� ���j���ԏ ����&�K�c�rX����@g�Z���@����~�H��=�k�U�)~뤈��dK*#Ç����m�Ԅ�VV�8ū�MJ���g�d�%�0�(B*��a�s�}R�C=C����­fo���bi8b����Vŧ,�y����A���Y8%?�BB�]�O���I5�t���Y��~�E6�l���	����F��i`��_V%��WG�5�	0\�!�Vku2Z��Zjo
����[��Y�2���O�E{+��s��}zc����>�-瓹��L��(���!�"FV�ivaI[� �kA�_�\*٘!���v���iI��(��L�C�A�>1�`��Q0n���#�2j���@l Ɖ�.�T>�3]/�VY�D�r�P�(A��M_�Q�]��rH�<�-k�?�=���L��g�*
��&�
%R���#��77wp{�܉
�N�w��?\�q)����5�Vf�Qy�'7��W�O��rÂ�ԕd��z|��E�K�D�!�hĳY@����Z�8�Wի��@���Qʘ���e��I/w��4�����|�����M���O�d����e&���ОU�pB&���	+�Lr�E�����=V���\芠G�[\�mO��#q�S�����ߥM��t�"�`�'��D��"�+�	"�\	P���,�b������K�&z��c�X� M�a{*���ه�=��ޢ��Uc`��t �r����J�o%$
�icZ ;?��#'-�7��=k_�s�@&����v��1~Ȣ)��b[m: l�؞Z�Fm��^lR������LI���5&�gZ|�LӴ���s]n���킭�gڄ���HŲ�y��RxJ�*`�^������¤a������$A_.���SYy�Sip�V������ة�u��VSin<s��c����ځߋ����������[6΄���@[O]�!η��:':��g��Hi��d��lΠvF�F�^���yU3c��#������q��ܟ��f��x_)�2*�½蹖L�LI��Z�UH�o�;�J>2�[�D�8�����$3ux�6v�|���������s=��"u�n)�B��G醻����ׄ�����5s
h�����ů��1���YX�@���5�S��bt��n�nK)�����q�[du�UH�SqM h��Aw �������!Yl�����
�l^EltL�\G��:&�M �s[�sd祋���6��S�8�+��F/�o�$�����+
���C<�w50��� �� ���No���7�5R�Cŕ�U��d)2�;�±싽Q}e��Up>����>/�	[ �J�ut�����֑/��X%���4�+?3LKv���Ԧ$� x�pw����1������g�HW�b��FO�6��%�|�:[N�ܗs?���Z<YTb�Sd�f6�­Y4B��ŅEy������f�v�j�߽��w�)���;2K~���Z�,M�����t���D�zKґ�.kP�t7竍diV�!I�̷�>+�\�g����o*��-��E%�V�)�d�g�x�ݏx�S齵��F�(�Ň�%B-�e.���Ra	�Ҭ�}����0�wO\���_�z9��Я.�R��7�(�� ���&Z`jwfgɼ��mL�� ����خ4J K�����-U��9�4��(�qx��W)����[�O]s��閱�_ ��h`�0������H�&������&�\��Vhj�� �#u��{-ϡ@�m��U�6�;-�V%_9�~OtZ��6����vG�/�D����i������F�n�G2���0?�����ÝK�a���'�o-�����H$3{{пK:>�4���,[k��W���<b��ɟc�;�J��^[z����7.]b��p��� Dư���1>K��c�*Qh��U�V��A���c��Y��R;�������O'v=74��i�٤��񬒗��,^���=��'V^U��cS?z���,��3�`�:�6�U�Lm���܄�,�5|x2�~��Wq[gټu�؇-g஗c��M�i��ԓ��i�`e����q<檻߽�˂��z��$ktQN��{��o�2e������<���	�̎�guT�ά���^����1I{���eˣNC?OoQ���8��X��	��/�rv غۢ+��<56!�g���LD=�L�Cn�W�.Qä������ 2!c"�=<��znٌt~$���?8�Dt%P����4.IlJ��l�Yߍ?�~9�6��Bޫ����l~� Z�qؚ�-;1��ۯ�SI�#5��H�[�7�C�1_R#����P��U
�O��� �D �kĒ�^� ��M��iV�m�O*��w�,3\���	��Z�u:�L z���{���ĵ�����	τ#06]�yn �tY`*���}
s�9y��{�d���g/	|�w�[^YL
s7��2Im�C���	HG
�+ �͈�d�y��� �H!�>�[�'Q��A@�@�t:%�=�Xhd�2D���8�>kYҀdZE*�a�1�r��0 �L�r���5�c�U�(��_�=��TC�;�F����bu�+�����r�frm�vJP2�q0|���X�[����B��^��J��(�����ߜ(��뿚�K\���ӷ�s3{�_u��b�[T��^}�#@	���/���as���u������}DL��H��$6�
�[3"�h#� v� �,1$c!��}�#�9IHC�͘�{l4�����.r�=H�(+��]\pb_t.��l���X�����D4���T�"��#�n�x8��u����ōg��	�\�J��Ʊ�J��`$@q'��1�����*�h)¯n��}�A�dఞg����ԞCg�����kO��t�P]%7lf�8(���x�j6l�#i�%xٸ.�ے���[^��x����J�~I"����}S̚����'�����9�NYv�k��8鈱Mr�ͤ+�B���|�H��a�cڇ8Cf����k�̊!�H���>����[�1�}UuNW'�`��K��ďh0���P�A*��z�I�X�z\u�FP���@x��"��A����U�5.m�
M8Wv�C���!����v�f�@�y���Ҝ�+QL�.��p��z��Ebq��3B�j)��y2�͢��1S
��A�!����R���ل׉�Vw�mƜ
�$�r!�r/8h��E4��^�?c��.,S�rW���W���s��w�(���tǩ��z߼_�EK	$B��Q|�>���u�1�Ok��7%��7SE�GG'��a�r�Q�Kd(�솧k���AQ$����3�?��֒Ar5���!���3qn�q#�w镄��A큓FOj�ް'�r_K6�8��xĈ���V5+�ΊxB�N����u�X՟� �-UsgjE��������>B�֚��q���c~�0�֓���J��T[J-ÕL���%M�^�������{�'�Y�"��ms���=:*�[#rV]NC�/�*q��ʵPy��h�E��Uh܎�D"ǩ������N�L�C@��~��␕'�w�Sɵ�%�3靂ː@9�U��cmg c����@$��J;�Q"�� d���&P��SA��z��#��J�=�������.��8��[j?{Wu����#��I[�ہ����2rl)��<�����<��C�Sm <��+�C��
�2�(DV�3�o�r(T�O�2�[�7 �c��b&o��ġ�U����S��zvK������D�P��i(e��1�����wB별"�J���a��=���36T��X�,E\_�JkY �ùr���B��e�������:���T+����\��àO��Q��"���d���̸�h��I$L6#��E){q��U���Yڎ�AuÕKe��(�z'f@&[�~��WkȖ�� ��J��-9αz��Ìu��lϔ�q����ؼQ�e�Q���$�u8�d���a��:�:����)�Pu/�Q�X��lH��n8��ݬ�5m�(*�~~5Zl`�|��ב_`�-Hg���_oWɞ\�`��^ѻ۔��9�y^�߿�A��J�L���Y�TV�CR��c�H|�V�6}�K�x;,|���F
q�6䡔������mk{E�p��/��b]WaqUL��,�OD^>6(�9v4&���[_o��QOY�(��w�qD�����!���tT�ä��y�gqY<���&��o H�u�j:�Z�o�?K;t�#����ëP�g��x��_\}1���ǁ����kR2�F��S_ȧ��O �5Jn:Y���<�������
%zC�t��>���d"��.�Rw�G��hY��򟽻L�v��IWԾ,���T��w�׹�lh�:ei�C`���Yf�VJ��J�͗�Hwg"N��  	ky�9�~����\����P9˘j���R�#���l��p\p�Pu��-�~���B47��H�\;설x�Hc��Ym��mc�[��K�ۻ�7�K\��	tc�VV���+�v��8_p��B.É�$h�8=[b��뉇�-
�]9n�[.e�P�I�c����4�]T�W���TS!��V�,z�G��@g�N蠰�uh�j 1?�����N�^<:�-?E-Λ=�@?�;�zW���T��얈� q`o�܌m�(�3��/�5u���4��]J�F���:4��90p�2�տ�>A��`�<�Ԫ��?&+�fei�=�[����_~��w���n'����M�x�I�h��OHyUx��:�G�.�B��iw�����O��xnݱ0	e��5t�=��i�X����w�KU�S���.���~{ɣo���H�7T���hJ���d.�/���<҂��lI:[��񋶫��ew��mw�nz�g��hBp���*��$�8k#�?1�3K����5�T�j2I�ڳFT��Ӏ����^3������І����C�օwH�A� ������x�Z%c��-b�������@��#�|�LB#���ǹZ�WD�SY�Z&y#L��t��H�o��pU�`5�X���(ߨ�Ű��y�������`&�PH����d�(s֠�`4���yٟ�
G���))T��6u��I��:L,��V��C������ٮ"}�B�)��I?�?����Z�R[M4�:�����s��#w�˖/��ߺ��P���u	l6&�Uã���u�ͱu&e�Уr�J|4K��ॾS������~�`�Nk�ߑo�2S<b*,"��DJD�4��0�æ�6���u���K<��	e�)~��~��/]ZQv�o�:��r��Cmm=�X�.�,A���Nl�m�ꊒ����ǩJ��G�9%�?�T+���g��Aֹ;�2A�X�Vj�]�IE4�� �j�]9%~�3�(���@$����������N3a���W�_r[^-D�7@��8�i���;ߔ���j���w]�5��-���R4���l�]{�B� ���$� �}V�v^����׈���E�n�X�ܾ���)P�zLk�Ah�ģa�M�L��/��
��~]�<�����~�֮Kt�Z���ܽ@�z���h�CMi���n���ἡ����v��+�@)�^�}�βfs�J@�;���ڀi��4���v%+s,����7�,��V�������J�pϷ8�([jq:KĬ߽HVw)�Ɏ�J��V
����oW�+`q�,�z����˾��}�%g*Q�9�	�%ވD��"�Vs�5e����/�����K'_�
��{�F2�G-l��a�eM��&rp�,�R���c~��e�0�45o�e���E,�#0-��eK���hd5�rRUe5Q'�h~����PM�$�-�}��ɫ@h〾��h$*0��ٶʈ:�Ve����e����s�bۋ�0&\afR��t��7���-ݮ���M�ۈ���6d�ڿ�e��@eNda�4@�D����2��%(8t���gw��j���	,� ��hC��.?MHG������B=#���R�AW�L�܃= 2ux� �f�!��r�����
�/$r�o�	0�����WN��v���4�#�W�몵J�=h?<�h2���Ր�[��r �߄]�� ;N��(�CBDN�������~����}���т��(1��\1@���e�-�*�d1ݯ]~��_ͦ ��Pӄ�I���W�h�!����w �]�٠�ʮ��'��g0�">X���܏N�~�mP��d,��Gz��C������X�����sVѵW-�qB���F�� 4��Vd�	�z��nv]�Rb�l���Ϡ
�ɋ�Հ��E�o"j���{=�Q�B��JU�
%�Q#�@���fc�����ҹ�����H���L�$ď�ϣ`\���ܧܵ���lCj�I��"m����=� �ܸ�<� $�?骪�.�PU��r����Ȯǉfk_Ȁ��cMtBȕ�@	u?��-¼�M�lj4�c^MX�F��b��T�S�B(�����-+�������o:��=��T�o�M�Z�P.1�v��ޞN`��}9f!K��r�b��n7�׿�ӧ�=O�woD��ī������x"f�0�� ���]GՒ�[��8�ɖ.`0�I�5�F��D�N�nt��%j�����Cx��?S*B�I�].�s���7����*)��|�,'1�_�b�Ï����_�M�F�w�HI�/��&̼6Z50m@)�ߢ��(�*�ա��ѳ<>�p�v��CU&[�)H+a �u^ ���]��L�����1h����
A}eB@�.�7���/��+9�-�6Vs�$��R ���e�HoWy��\���$��h����y5X���Pv	�L�7JsE�Ui;��YۉA��ٝ5�@Gv/�_�V?��|!!��V3*k�T�r9�S�H9N�D�K�,��6�X�1zRmm|�A�(�����l1��r1E�9I��{Ƨab߳���Ju2�Hd?�(����a+q��4�S�2�>y<���ނj�xQ��D���:E�/�-��*;�8��Q}Ak{^��av�m���.�+~�(\�Ler��q/���5k�0`����sB��7�k��߻�=R̐�^ H������ݮ
-)�țr?$���8dҨ��6�f��4	���dGPn.V:[0��C?��%�m���i�(c?����b���	]Mt�����VL�ْ�s���֛���Np���T�뚙�2��c� �{a@�t#�F�R��X=�
��4I�؈e���hu򮟹�L0��X��%RlN������5J�S��nD��*N� �KVO���䒂����
A�/ѧ{���k����6�Z��;�W��D��>#g��Y�N�FLzlJX���v�ik_ö����3���t&��3��,�z�x����Xw���s^Ξ�J�Pz=C�����r��ENG�m��s�~��p��S���V�D1��s	�$�D��R�Z}8��7��!>/]f�|�jK�ؠk������Z?'
�A�;]���>厁\N{n��L����z�Ζ�F�Q)S$B�; њh߼��D`�P�L>~�-N�K����
�ϼҽ���p�����gy"���/�0���pְ����UY�?�]0��) �gš��Ykڡ6;#�̌���$����;m��#̚P�X<ۥ�l����X*��W�h�-�ᶜ�w Đ|�W�_�?�:�F�8��*�,�z��y�ͣj:��-�P�,�{� С���yU���%��J��1���R�t��Bc�hE7�u\\;����t ��H��L�kγ�J8���I�m�E¸����a�D�UP��.��~墿
d5��p� �S��iY�g	�~W�P���r:���yݬ?wa����^��('�\v@���B�D^`	:r�	.	�pE�-��s�LE�U�=�Oиe�D�3�^��E�H������Z�,Y��V���	�-Y�_��� h�n�(qA��]��Q�R[V4�-Τ>��ݐ���� #&�v�+.P9&�r�*"0�Y�m5�")��ǎ��O>� ���4�5r�Lbøv�#��!s��UA!�#|$s��x�M��q6��n�-���BQ?NF�Ņ�4"�	[/Z��x.�R	[�y�vַ�۸
=�Z��������V�/��*r �`Va8N��G|�V�C`-Dpv�st��V�Z�T�[M���8Jq��л}�\̼ђ#5aW���"H!��s���`��g�Eh=n
����G��;�9@�%��*��z�u��2Yh�v=KF
ѷ{F����'2�F������/W|\N6�zVbT�nb�!sx{Y��cT?��]��L��m����ܤ�S7�����}�����-�h��������u ��;O���w��t0� 2*�J�����%��M�e#@�?�DK���<|�+<�F��wPA���2����n7vM��0��4�C:��x�[�յ.���E�����#x�4��`.�}��m�g�%i=��b�!8�
׽E\��ku������z���γ ��3خ�6F�y/���e��F^9���rSتY�)CM*N4q����8�O�/�N�����5��֡�v��3�2D����%H�#����Z���.�xqo���Q��3��c�'o��v��*&�#��KU�&^�_��%V�q��Oۉ�N�U����UxΗ�[��t����(6�b���SAt�ކ�2+���Ӽ	_+�����L+��5�u�	�G���C:����C�l��3/b�Ɖ�YqR��R`��DN��LsnO/�	�؝qO��r�(r�Z��7���-�D���ٱ����bt�}��lM�tNpƵbm� ��'*빰���RTl�Rs��?3�P�^ޣ�I�y�y�*�nM�Z�c$~�°mi$
3N� �8��K�H�����aZ����͵��?=�2y�L6��ų�C���_y��5�\\P�1O]fh9\��K�]L�&�<R������%�>l,V�rc&r��mj�H��ʺ�s�	��x�g۔�(�?�l:>�e  ^U/���IY�Z"��`�����!��>�/~��d lSXaJEp���)�8	(�7}��l��D�v��+����j�6zXN�	(��'5'��R�k�7�%�*(K�Qbs�0�'/�̞"�Q&WӔ�r�Ұ$%e����sM)�!��a��H(�LE�CǇS.��Qo�����P���t�޹v�IƗh���v���t]"0x�Z(b������J�NI�%�W���i�C�I6 ���ϕ�,z��Yܲ)�{GC�՚�l��R���,.��{?�[�#���o-��?�Z�vF f	X~�W��:Qm���q6`?���8�E9������L��1��.�﵈?�P� t�؀wk0�^�K�bH��;�Zq5|�#A����]) CϪ�'��	�b����|5=:�_>D�8"=�%8�ݒ����[�p)�5r���I�4�shBV��Iͱ��C��1ѕ��,D�W8�v�8-<e�A���ޭ �����-�͟r��-��qш�f��\/�a��>/M��o�Cő)8k��C����m�3k���������Ѕ� 4c<���"$N`�c�'�EI�d�f��s X'���#�`�@�kPX�>�:�)Cʾ�n�oH)�T�W���'�����������4Q�o���zD��z���D��+����9�ӻ��	��T�@?+���|�S���8��n�y�?L��a��yv���"��M>�7����j�gx+��L���;�[�T�R;UX�_�ރ�D������~�{��OJ�+�{[����a��Z�O'6��0��yKɞ�iz����=�@Oi/�f�����p�]0��:ԟ.���+�n���rϥ���ݖmy݄�!GkZ���q#מc���Ŭ4#���h��p�����v_������$9o��u9�ce*X +q�Hb����R|�P��{ѩ����F�yJqm\NQ�"�k�n.+ڽX�q3}��k�\ ^H���񰋷,�����f��c����``ގj$�\%�v�U]�x��}VK�� �˼'Q���@K�����^W�`���\󽯍kT�<��uC�O������G�	ޡ������?��7���2���e��(����-r�w5J?ӪTj!й#'����t�TK�������S�����.�ޮo8^telC�2�MO
��p����{���e|�{������� ��>�3���K��#�P�*��������
?9�������������̕=�P�uMlY�o�1�5������%��nXǱ\Ω8 <��4�`/��ϻlv�5��a�c�Ӝ�~�.��nfV/	��@^t���-��S���4���F��/�p�I�GhgwI$��W�`d�	&^����f4rbT�z��m��\ʄ�K�b+��+\����N�%�QX;�kݒ n�x�`�lHb�g����]s��ϔ�ٓ�:�8���]E�keƍޛ��K��`ȗ����׊@ޕ����]��)WDT�\j�p��-���n6�(*���=O�w+����̔���(@�̄��?�f�E��� >���X:�pTuF�AT�C��o�d ���\��k�ܧ�z9cPl+�Q� ���dTk(�T��r����fs*�l)�gd��WH|ܒ!��o䖶D�s�.��&˙��u+�����?�[���������7	9��Ѻ�'�G�*;����)��M��*�!�d�� �[���8�`t���\!E���9�J�au�����rF�D18 ���ybz�ѴW���^ŗ��z[Ke�,�료 
���]e�$s8o2O?q��F&�j���� xJΉ�[��^�W�����>���4bP�Cn����<�u?�/����b�xJ�tm�9�K�'�ID�[����pd�Y|x�#�������]��B~���RG�o�f����h���a����:�����Q�8�-d��|}R�!Գe�� ��)b}�T��������%b��̵�� m�u�V���{.ߟa�A�*$�́�.�ָ��Ҭ+JR����JY�w��ܡC�� ���Ã����x^��ٖ%g�X�&S.]zrXE�C�'F�'<���ק<p�P$O�IYp�	ʸ���{l��ӈ���Ӣ��#��r�e�8���{@����'w?z��ųM�MB�߲s��`�m��P�Ut�6�ר����ض�8�J ͷ�ӊy���ﶷ^��)�!+�U\Rꗑ&�m�D��8>��^��"�CP���ŀ_��@ ��P�|�7~�����Dj��'�i�<iM�������w��K��O<q�z���#��%M�=���[��#�C�U��b��r� e�[�E�%��#$Z��������d�`AN�A��k�",�3�d|f"Í���-DzC-�T��<H,�>D�|�����c�}�� �����&N��y���t�읤T �_�p���_!�[��̯��j��w���e��ыl��u�˷3Rq�
=�1K�F��D��]#����l���g�X6��3�T[���ž
/z���-���q������#�����7����a�O����>(�?�/��x�
Wh�bjKɲ��?]VU_B�%A����iv�r;5���p^:����1����~�-�K<�A1��Y����˱#
���B���d�2�"�N�ģ���i�O��ER̗��Eҿ�#���xX�f��p<��A�=ِ!5��==���f��Jߪ�3���sO���ELg��F�񩦷���)Gz}�A�և�%<����ھ�n��j��}�0[�.�ʁ��z=!�O�`ڵDl&�8�#���yF̠pXV�Y	��h����5)�NG��;�}�e��O�&�b�}�p��&�sT�RdWNg��*��,X�����Ĳ�z���ä�Z��}-%@M����	�����P���|���9�rc�E�`aMq�/���R�h<�-��2�9�gN<�4*�('m�s�<��#Sb��\a�u
�[ua��1�V��9-�	��+���;�vb�~ԉ!��x�����:J�z��#.6
�B7�-�Cb>i*:D���B@Y�z $'�2����! E������WXdAJ�N4�ZI�k��{�I�5 ��/���J֘U�>��4�Iyts�( O��t����~�#�I��X{��� X�5��N��u)_Z��/0���陋�U�@I�V��mB$`��ږ����;���E7�.d8� ��ETn���݆�� �����b�礼�KQ߬ƫC�li���n��J��D�${G����D�Q^�)f(!�;c������'��#�!d9�ٱfI%��Y����8)����78
��P��
Qx�oŒ d~�;�{0�b|]��֏���@��me�)D�ɥ���'c��)|y����`��?�k��E�}�&[�p��?�^���jZQ�
�N2J~J���OgA�s%ئ" -��*$����d�9ä[�A�Gj�@פ*�6R���`����w��2��=��
n���R+NǄ��� ���9 ��ʹ?�'���Ր�_�l,:�1���Վ����
LP�wa�q�.��A�#`���6o�S��G�5h���D�@G ���7��0�B�Ϳ�p^�G�E�i��.@�����J�ų;H�{υ�.E�t�A@v������4�l���5�s�j���P�k���틟w���v��}���邵{�\>��  �G���gpU�.���q=��INC�5���KE�K�Xv�-�k@�#a7EVN�N.f�5��+�A��a�\�	�Ӊ�$>DI�τ/Hy��j;j@e�~g�D��]\CGc�Vށ8�!Ē���gQO�?����E.L�\�(��퉕��9�3�M�q��'N^k��t��?b����-�JfI�h0}��d�����:�P���E���>�ک\���O��"s��>���>�J:y�!��>[4�6�����1�����f��@���t��Zz�Z$BE�O(���-�+N���X��PC�e�},$���M���x?�u�
Xct�a:^o6�l�hb9e)�P�M� ����}�^����ݷX�����܍��R@�6:�8��'�'Zo�lg���p�/_���H��b�&��1���_à��Gρ�tG$!p�� |o�y�_ �3 ���1�pFE�NP�����V��^�$����5�u���0I��Ej�N%W����0���#�ƣ�����m���h]�d��pdkA�f��.c͸6'B�H�&@.ڏw�3�_����d|����BVJ�3����Y[X�Mn����ҺF�d��9ou�h���&Hl��*���� y(ĺ��XN8�-�s�J�w�w��:�p����&�eg11���3��;r�H���X��|"9���Y��lL�)��H�ٽ�^�-Ӊ���ށ���*�EĿ
I�����#gΥ����d3��v{�XZ&���Bt�r�J������hoX���	���6)������~c�}��ؒ����ʩy��I8.�;���M�'�Y-�޻�KV��E��f �Gi�\g[SE�7�Mt�eb(c|��{ 득��"T1�N�u4X�M���ÆX-���>��J����4��y��6��͠�/Bׄ����� ���E�!�2�dKJW����6��M>,/�2x��9�'�O\�0�k�����Ҿp1Q�Y����ل��P��|�qW۬�Tf�M�?)|7X��zU�Ѥu������-�M�gh���
�d��$[�e�M�:D��b�q��,�cW�C�Q��j�n���m�ڲ�C��%�De]��.�*%��qZߚ�(.��?�qW����kZ�):UŘU$W��Ӓ	-t^��b�ᅎu��^A�lTR��;-�nmi�doRŁ[D��\�<aǏ���<�����ƨ
>���Q|zi$����A��y�|�q����"����0 ����
j����y�.���:�J�ͪ�)��n:�ʹYU[:��ؚ�J�w+�G���s��{�7)fH��wA[�1o���'�v���ghFu"�����X<��.x^B�%������"�s`n�'��bBd>��c+H��N�qB�NS����V���|Y����?v��.���}��Y�d8MsS�[E�-�L��&6Ε&@�ו�SC��̒�~6���3���ƫGCޕ���I�(_N�ƌJ��d�E�y��ۤ�ט�G���ϲS؄�C���mx��w?jߎQE�8�	�$o)f�g�E����|�{ei܇X����~8p
�Gl`�Q��}��NU��aVb���dAp�e(��\��C/o}4��}���JeYJI�υ�c��[�|���_�[y�\ǣj�����KA Z�pluT�n$����L��	�MC����O�i\dڋL"�M#o�s=��$�(�b6�X���v��_�Ώ��7��Y����wT'����L��1ˈ��E=L�rGRp����
�$�����1l��LqjD9{aF
A{��8�$ ˮI��#0��:w��i�����I�{(>�S��F}���K�G���y[v9��˽Y��7��VF\~����X��2�;K.V�I@���LK�|M���&0iy��k�o��<ytO���\x��
�<��`iİ�e�-���޵��a�����0>M��l�Ns$>�F�qw�I�2U�-��^?��F��1U��G��@nf����9#��RL�:�(a�^Vésx�F�� E�ь�֩��J}��f-��|��U��� 4R�)=!H9@��!�+2�����(�&����Zp@e���JT|�����$�풜�m՛��ѕ������%kj�b��_G�I�&��쀼�	'��������<K)3��Q��GY�(��g�4�_���@���\��x�"�@�b�PmȌ���P���M<���n?-����:��py�r$c5�\3�Xm�bIo��q'��By�a�4B�5��0Pܜ�r��'��p$4mCZ��
ܝ�Oc3�{s�y';tV��Q��ޛ�t.�}��PT�M���a
:8�;�we#��I�^%F���$�]>�"&�#��U �Zb�Wʢ�
�&z���ޱ�=��4�z��k$�B}��:W,��+AH�(z��~�27�3Q��H4��*�I�"ʃW%�"ч� >
��-y����RUxHF��ކ����K>y�2
`��f�+Q�ϧM]"�^IQ6�۔��'λ�t륚K3�Y��Լ �)�i��j�PS�G�ɏʠh��n�m+�ʫ�A��_�{�?�^�
I_,�`��Y������(���
P�����C��=��h���uҪ�f���%(�*3G�﫶�n���AP�����I���)��<#S�;&ǒ����S����a���ͣ)b	�2sՋ^�XKM�+q��I���c�SĖ���%��Cc^Q�+N�a#f˦�-s�:ey����/ez��0]�Q��V"Lpӑ��J#C�F��(?mQ��srvR�W��7om��<ք��0�	���}�]�f4+aq1�rxV�<���3�!}W���K�k5̦ؔ�K"�nA\X7�(K�2T��FB/��z���X;�2WP��z��h�֡͘K��5`Q��_�g�ģ=�ߠ�\r��L׽���n?�w�0QL�<Wu����ӛ��XM{fp�~��DY�%��