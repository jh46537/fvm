��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&�T��%�h�B�?f���H9��?U�7��%��5]�:u�j:WZRto��{�3}�(�JO���A�����ǘ������a0���^���B���R�%՞���SP��]$7xk"k�&H�(�. FC��`��ƶ},O��$���}�'���mX���K��Z JrmтH��w�|���v��N@:5���  i$�˪�Q�Iq�����r�?�E?�Q�P���9�IN�F����:���3�ِ�`	�L;�� S�W;�I�M�������^�[9V},�o2	�Y|���\��{[|x�}緛��-���`|0�66*�VGgu`eJ]����z8dN�9ۦZ΍-�(�}N�^�GVG �z��%X�H��jԵ����<)ojV��Ή�m����� �9/���R��g�mR���yP���|'V=?�� �I�hP+R�)�56�n�`�Q/i���l�����C�}M@m��0�XVDF|��9�̅�5�]��Rd=�S씬�!�H�"4�'Zᶾ��� .,��O��c�$��Վp�����r3Z緖� ����^�k���ׂs��X�䒊U�0
�K��4�E�-ղȝ�:ݻz9S����/�����7�����&�V:�Ck�_|]�jq�f�ե�����a8 ۋ&���>@�r
��r���Ϻ���q�~�M��݈|9�K�a����ȇt�A������_�{�0R�s��<��O�q6�v2=���7��~Ä&���$}CUk�*��P�O�XX�J�d�֙�����kA���Mr� ��RrݜgVǖl䦔�ꢙ���ef^�a�W����j����!��ȢwA5GwD2P�����HA��0��[!n$4���4���I"��2��D�
y�'gښ���5Y+w�e���;�|'J�dh��T����K�b,�\�MC�r0�=�{e�qh�I�A�l�z���9H�v۳66��)`?&�sT��܈��A�O�98d��+�T�BCg#�瀯n>lo�&S3��]+7c���43�!�Nuͽ\���­_G/��Hn봠����; ���ӻ67��5��P������$����5���;�\��OR�eW��pv(��>�w��%9"�V����m��~པ\�.�`��I�Ҍz}�i����������:�:9��W�Ȕb��͖�p�����8ݛ{&�}q�U������"�+�%�9��?ۃ��aR̴mV�><+@T��D�����FP�`(�y]����Mv������.���K1&�#ګ�lX��h�&u�^|85�\��_M�:yV��B�dCǥ�Sny�/���e���{�Fw��T)ɜ��RjgЪ�D��ɦ��
�Ůa{��7�p�h�5E|�S��@�9<O�l��z��y��m��$6�}�o��b�h'�Ody��u���t��9���������R$��1]��ڑ9���������u������1_�q��ɀ�J䞍P��u�:Ψ��3H}�����p�����⁔�|E�&���|��e���T�;T�}FHA+�����?<�#�D�O�u��]����*Pe'@3`XE�yg<k���8ݕ�'{��c�B3b�"�~��*XK���P�[��~����/� F����"���_s���K����l����F�Ec�4->Z>�k�R����l����;��GUa�(�5r{�v9�Y�*p�sT��{�𹷃hM�����Vk���,y���F<�:�o��8�+�R����8�BHT�z�)�G�E2�����%��Kp��-'�pu1.j\6�,e�ޏ�qT
���h���ԣXI�58,m��*W��
��${��Jl���y�Zsܩ�Q�'���(�OŸsڀ����=ݚ5c�ѫ��@���h���p�˧>4KN~ڝ?͞����,���iɞ�W:�j؃g]/���ʇJY�~�Q���s.u9n��/I~��/RF�X,��_��,���D������T��!(N���$?�~C�e޵�d+F�t�Y����}u�cEn���2�Ċ�}�b�X���Hf���^�w3N���8���p����?����`�(�����B`|[x��[��vE3T�+^b?�LE���u��p����? ���х��(���د����ӯ��#�0��A��!���>N�l�R����Ź�J�!_�)O��{�t��jOJ��ê���)$��xx��۳��*��~ړߦ�B؂ � Q�P7=lSY�V5���IE���@1�)#r;���&���儸�L 9#4��9w����Ժ���/�j �p�]��R����sGf~=�)�X�0M�]^آք y���D��'�Xtu.|v��;a��_k'��x���9�iv37���}:ӿ����Y?���C_p��s�8�if�
K<�#�/z��Hz>��m�Ӷ���']�  W���]:6n���Bt�H0���N��fm���	O6R�%���Ӓ�6|х�D�����ی�E�#V�����6���T[^Вm.-S��NHJ��Y�j��n��j?���dY'U�R�d.�I��_��	�@���(�3:fGzG#ܩ%���}� C����|㸼UKxpY��U�NQ�����<$J�����rcl�8b���j����������WX�`"��u���Ng��B*Ii(�1c�ō�AU0/�.H��2��"V7�qn�����h�V��*�����R��K�$˰�/�4G��TN%DKa#��U0�&��/�!yԮ� ���X�d���/�2o�g4fF*"B9'F��@��>�͘�,~K9|���F%��JY�����sp�a'��Kj�*��3�Wa�����(GQf�	��Ƹ��'�j�6~���L���q̋νES{��30|�Y������t�Ȁ�w��	�V��6�/���!~�2k�8x��{)��l��ݝfm�W=Z� �:t��2�l)�.�^��e^�w��3�.4�J�����v�Ѳ��a���󉝸�����������)�F�x�u��jx62>;	��Q��칺����۠:��Nf�Q2��)	#��t��0Sy��?~�킸�����D��c�i�T��ws��,D0���F���x\�ʜW�
���ԙg�z1��/��$kV����@� �k���	��A�T��� ����6;r��G��[��
���C�X���TyC�x�����3�jM'��_�b_0�KʀS�����C6��C8��w�$' 3��]PF^����ZKd4�}5k{~I1aۦ��;O����+���X�ea��n�3�_:$�H��� ���D���c�IԖ�E@�~\��OA��,%�����!�n�Jk�>�j�Ϫ���I�;#�)j�U.��E�0��Y���!-��lW\��E��#�A�Ix���7�_SŀL�x������?��Z�R��]h)��ۓ!��'g��/�{����I�P�߰?��Z���R���1d����Ӫc/�W�RSF@��Po��	-�`�qA�.&�;t��4N����+O&R�yCx�b>TQ���S�:_��e�o���r���+�W��Z�{F��%q�?�&s'tP{?{��@&�]�je7m��%"����*Ie~�tU�Q��\%���~-�qz)��E��.�]����_�fַ9Q`���]9�c�clg��	��Q��q� ��%i�dF҆�ۮBv��n��V�=��W��A���/���r=k�0��L3m�A{p2�f1�i��W��|af���m��%��[v�uA�7�.6�(�#�<]a0S�d���8#�L���M7�&k��H=ȣa�l���2��s0�����<��o����'����bR���aCG���~z�W{�flTO`آ��r5��;~>�q�[��	f 8��.���(S*U����1U걛#|y��G�;����7�ʩL/�z������C��E���ˇ���I�o&�qTd(��d�'9M_�jNTI_*���<]Ң�t��7'�J���/tv%UC�O��?��v?��9mp��cN���Ss��Z,\4"��J�/�3E��]����
(w'��� ə}"Ս�W>�)���z�������D����)�wC��t=	��4��YL�Ǽ�I�@��aq�HQ���$�)(�:�ѽ�N#�E��n�@i�Q��>{D����9�q|��p���Y��,�h��M�y�\{Dk�Q�В��O6HJv��2z�D��;|���(kV��B�r�#~�fv� ��mb��D�u��qrb4������U���W.q
.�jԆ/��B��<W�*���+5���N�.�d�r+`KCQ�c�k3����,՚�n%8����g�Im֟��̹f�'Lm��3�i��|���a���^�D �q��
���;����1]E�:+ׄJ5��V��y׬��[۟���3�jW��l �K���<B��]���M����P�xHd7�ʸϻxg�i��Fl�=����ր�}ar\��Av�����襹M�H�(9�'��g�74Ƙ !��^���]�9U<d3�5AT�������^�֕��c(��T�u8����(�sjOl�Dn
n#�8<�����TO�9�,�^��l�����a��r�a�ÿrW-;� *�D�I� ��i�&�1q*k��"d�F�s�P������C�(Esd�G!���� �����Qh`\��N��J������������oL�ߩIB<t��IY��j��W���.^1p�/�$��})�0nwe���u���`A�yYӫ�x�Pܜ���.�/��g���-7�\<�j��R7�1��+&�o#E�iRǝ�2X2�)�nޣ�8"��@�Q����[����,���b��Z�����#x��&�ҮE� b�p�
���h���x�q�����8�2-�w�Pu3˚�7����-U��S��J��[��U�����/\�� �~�+��S`c�0m_�LY��'`|��V��B�����̓/f$�{��$��5�kCۛ	Q��B���q���Q�Q�������U6V��y+,3���y�yi���Mz�L��e!��ܚ�5�M�ŒE��OL.Q꿓$#~�*%������u��������|L�
�O����Q�:J��KYC[a�!N�D��6�u��i��[ȹ�� ?�"�hl�0W-�d�ԑ���yЦr㤜[r�&��14�<q�I44�KbW�{Q2V�&���!yT8�%�g�eK���U��4� �>���}��0�_XB�H���11�!���c���hK�?E �"�.�sL~�!�Ъ;�s��5�ȫ�;D}&g�kD[�LeS�����.���)V�mγYH�a{�_�^6��y��mB�r	Q�7lN�����jPj�YWg��@�!����X�:�@g�uMFѽ�k	5����4��|V��_��Q�;`
�
�l\�݁�R_�I�yQ|�߀�4��R}�f>��*�t�>lM��}�qc�]ze��b�$��o�r���G���߽�K2�)M�2��
��#�Σ�ˀA��=�-�tϗ�e)��w�!�޵}�P�օ��0U�X몜I�i8��7������}C��`I���a�!(�f��cN�['e���m�s]�y��$ϡ�6uW.Ntn)+���p�l��~=���'�"�tC�T{��j_w���6�2�f:A5�
���9��;��4�5-�f�E]׻8V�N��f�ץ��d2��jv�c5�s^R1a�W��2DfX��Y�\�W��}�g��^Ѹ���1�yu�$�$����~A���6�>��sy�XܳAB���u>sƠ�_9s�R�G�z?�;�Q���i��rZ���|!�6�g�Tx����O7P�Ch|-c��&?i�x�-Ocʒm�eۑs�=Ka��>LP�<�;1*��~D2���ǽH].�Cq�h硈y�1 ���T�
�w�$u�n���)�	��%�@��:Ն�(�l$�dCFE�s�N���V$@p�2ɇ��kl��.�fh�Uv#��u�m�z�����U�H��D×Ҷ� �7a^�aFL�%8�N���	W�	��J��.c(�.Sͽ%�x��Zp=�����)m���G[��?�N$���E��fN���g��X�oJ��w�m�u�@㹰�Z	�喐�9B���0��"�xg��+�j$�ڕԪ���K�u��{
����Y"7ul<v���H��ʖs� �}7'�2�[*T��_0�fV�Χ�(�l��E�fY��M&�K˖��Bw���Q$8ͮ���!ɟ�h�[6i�p5@���I7t��ğ0 k��p6�bN�:��l_,��D�_y0��O��
ڦq����T~`��A�HXv�����ܐc��M;t0�(7�U9��a�`�[�	d���1^��돧���a���Pz`P����  I��1b(;D�;3�0��rO�!��@��j�8�jd�^�g��h�my�9�[��~uVx��O;|D���_��M7���vY�U_!�D�}�����-�����̝�y�+�"	Ɇ�Ǯ��g�	�<�i�sl %��"9`u�Ͽ�T�Z��q )�����Y.�I�����6����z<M:D�[C]�y�ݳܲ�߰��DM,?615��������T�3)�C	���2`i��E|P�'KN�&8u���,��|6%tmo3�d��4���1u��l�x0-ey�b7�����,����0o���Z=qdNm�^V��KN$H0��d@�?�Ķ��Y=.�M��Z˩
6�/�3�Ðm~ �j��mT� �6��e��N��h�RYZ\7u�wT&��5�g<[I�9�=��і�Q�a?����}�́س �ғXH����1�$@Yx��ӆ^c��W��kM�a�C�'��\�ğI��(��X{;��G��0Y+DU"���և�sQ���Y��d�Ave���)���i
9o�)�B�y�h��;�!��0	��w�aBȻ�Ń\��+/�p���j�N�3=�@�x�U^-�n�ˌ�hC��Fq�e�DHFE٣o��W6	��B�W�M��X��,���O떽�5�jX?���T�k{,Y�[H��+8��G�f1%�7�2�~��B6�m�c�˦�;6̼AhE��a@�ɜ��RTL�;�`7fzr5����{H'�����12H����	iBiz���V%�b7�5��o��l�/�r��1��
�PBx���x�I��e��a�>V�o8M3�Ч`+�gͩ䚦ڇ8��˂#�& Dabc|Ry*\L���H���v�g�a�Y�E����rK��.Ձ����F"e�I�Aʡd�S����_���������8t�pԞ;k:/3�Y�T#�r�u��qIm��.3��2���r��O��}sѲ��R#��ˌʚ�
�������a��2�-��C�	q�:�C��J�~��M�g|�=( ~3��p����i>�&�(��{�:�Ƕa� ��;D
7�iKAiz���g�`<@�rw�o'��	�x�C57�݇q�����>��kn08���<~���F�/��[e����J��0�D�s-:c�t���"-�����q��;���>G�8�ѿ���"s[G ]��H�Lo\�e������y�Q�}��(�G@o�D;8p�x���z��nl�&X��XD�ToN��W_%��W��`S7ƨu<����*���#~۳��QFҿwt�c�Za�0�e�
��H�
��1�=jFAy��A�_����_��~8Ve�!�5�3�j&����t$G��ֈ�Z����v3b�Pŋƅ�=<�`~�L�>'$VB\@S�,��
pG+ʯ�WNw����!����e�43��n��Te�C7�F�E$���C�����tH�)3�hM��r�׳�wT&����K$wu�G�/�v5 �CrU�@�?ܙH�O<��)Vi���b!3��ܕ��6��|�<FKI��:*j�T�gj����J��:⟤O�:��r�]S=v<��	���8������tl��q�6�{pԹ�)��r��9�;�#�13�
���y�>ژ���;����ݼ�B�����GJ�k�8�Zw]8?���s��?�n8���M���Y��gւ���4ű"D�h�Y���=�}�~.�8���-~\%8�3U�KQS�)A���0:I�\ua�0�;�PN���POp�7ʜ��=���9Q������-��u��F �z��c�@ k�2�m%uN�ox�������+�����˭�l	΂�-s7���i���
��9*���	v�?�e�к��Y�iW�-�9���G�l�V���<�:cL��j�i9m4H��)5)w��U���WH1Z��wP3&��F�ʌ���ي�e
V� `_ ��0ڔgu�2w�Hq��]�%B��F>l�z^L�8mϢ�� �B����X����]>c��$��p��ǀ����f�-$�[��9�T߀\��/��WUX�E�wO�� 8�+�X/�$�;��E�1�3�E� =��Aȿ�G�MI�	���������]�෎��"b�V'B��r�S6�J���K���?(��F�u��Ì|E	�o��
���P:g�Q�y?����p4�;J��3T���%�ڵQH:0�Z1��]ZS��X\w,�|��͞�B]��ӻ�$��+�����%�|�R�/�Q6���{)υ���)�� e5��p��@��ou�7�X��ڮ��	���o�2U���v9ו�q%���ū(cH����J�-�
 8Zd��Y�3����#��H��"���ݾ0�?(+<�襧兆m;�J���C)M[��W�B��Z��������a2ێAAbM�@=�cU�'��+�#+���Ʈ�(����qCYH::$��a[`������ϲt���wj�S�-jc̵�Ψ��
�z���nDݍ���*^��,�{����T�w^N��>���0��u	׬�9h��-P�<�m�p;��ur_|Ǵ��.O�vv��J��8�|�х�zͮm*/��ΑsX��*fhr�9�pCh�	-D!��ۄ`�:@�sQ	���M�֎f�ɋ_{#7!�E � a�Pq�p��u��I�x?�D���qw�u1����jP$$���+��4v��h�n�Œ)�y
7Yx�~���3�s�=�=%�X�R(U��\R�7uTXM{a������Q�B{����E5���v(H��8��+���1`NԸ��TQtC���WI���w��T��'�
���/%ſ�]�p*���4"#$)G:�h��6�5$/$�h���t$�9je՟��(�����u�����FQ�X���_#<=��!�C��G�P�(\h'��Z�gF������-O>׼�� a/�;
@n�ֹ0�va�`Ơhy;(��y6�c�T���\���몸�K怊S@Z�'k9�;���#���[p�7���K�R�����������F��GןzWg��NC��A����K{�V�1���72w�6���RQ�!y�]jWX�rǦ� 7ݏJ��= %Q˗f���PO�0��7`+����4U�f��N�H{�ֿm�Oe|�K��%B�Ӆ��\X�2��g���J�}�t�6�I�AQ���[�w��3��P��K<�L�1�'�dʙ�1�_ǽͭ5��pJ?�90&���D[ v�	�P�(H
�Y�� Z��h�:��)��L.6sv�{[�϶+I���X��I����<k�V�<6B:"�Q����;�z�v�N�@��w��פ��M�iC}�+_U��L�As�l��4�qhS6,u�G�Q9#���v`�ǰJ|��OWSE��#��yH8 �u��#��FI�(׉p��eO��E���$�Xu�2Q���D��z1�1n�X#�a�=�%����"��܃�#�w�V��bE��"xR�/PO�
�+��$%�Y6�(t��b���P/�&T�j@un9�))4��"��M���q�z~���Z�8�_���ȁ	�\����y X%Y�a/p��J��j��!�܄h$z�]�c@����>�3�d���8������S��"T�H�c}�^՚{P?3����eq�D��jV�򩶆�ۏ%kC���	�8���)t����&�b(Z�hg���F9�O���0΍n���@ݍH�)����f��xe
�mrZ�N��z�Ray |����]��sR�>�Ku��H�%�� ��^u�lݺ�&��-�)�Br����A|K�Z��k/((��ٰ܊�\Q�~{�t��E�tQ�D��ycth?J�i��u���[4�;��N��bt;[���Կ\���q8Xp�e���d�/���������@,GkĹ�[}�qw0ɏ��*nr9�p��t��v��~G
�$���I6�v6I��$Ӣ�p��LH���O�f)��T�ǈb�B�,���.ɾ��(erXp�>r��S˭6C&:_��੡MV��:�������v���olT��7���������u�X�d�&GO��d�|;�,{��]����(Q����Ky?�Q�+�O�wOҨ�x�˸sI��-���� � v٢G<�@�#"
�(1IC�O��䦰}��a(�E[+b��� $�(��"�_�R
�!��E����c�c�L_i����nd-���&�@��
(@5�pU�| h��(De�6-7+2���ڽc�p��:Gaǈ0a���9��4�}���Pz�7���~���mӨY(э!YL�=�]�+6^u]y�a�hߟ�,���9-�8�q�㱧;el*����"��<=o?��ˀ��ʼ���AdW$�t�V9�sؑN�}�,y���s��X��#i#<<�������ڻ�An�w�az�y���Z6<���I�>���Y�L?�,4�"$m�_#	j��f��hi���JG]�r����E��+�T`@p�������@"���`m/ؿ�-�l�܁��*[�j�<��F�?+\�|�!ytK#��.BN8*�9x�3��y0�,(&
"�3�[�6��