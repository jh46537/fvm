��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVbs����e����`#ql`NK��fC;�!�����J!X�v�����@��F�������秺nC���>U>p�o��m񍏥�'���n��Ԯ�'��؎��l� 
��0���u@T�|�J$�Ab���[�)�Bƹ��'��T����z���&��˄B��W�Z'�(����S) }���$����?�Pd򶗶�
\��#���Ӹ�2q���ҁͧ�x0@��#g��T��x�����0�AӍ�.� �m�CSN!e
�Xm��l! rљɌ*�@��W$�a���(e�:j�(gk�r�:��)��o��x�&o�{�I�6`�3�`��]O�ux�a�)�sLC�U�>;z�)�0|G��r=a����3R,������U�B��+��	>^<�Υ��t�gV�'�'$��=�G���H�V�����Z�lfCp�;�J�����x ~�w��l�2�՛����{��H��C8c��o��v��ԑwdꤝ�r&�.?��E.>���PE������BZ H���_9��z� ����z="X>[0�u��c4�Z{�Ï2�q��&8��p�PZG��nQ�I�gxi����Z��Jv#�%������P;Oono��oV��!�!���[3~�/�jo�v=��ٿp��f��>�Kni�a8��7!�dlʠ+����{��x����uf
�A�����<.��qk*�j4���AmǑ�����gi�2&#�?V*B:^�a2�-���.�(p��XC�:.����B�Pa�(ʚ������i�dV)q��ǃ�a������̃�ɋ������܁F&��a�� �-E���Y�&�@9U����{� �����L�`8P��A!���F��(�)3���Z���:����e<��L�ӓ)EsU�� "�dq�Ɖ��nW��6�8K>�6��5�a��PD�-���}y0FT^�qZϡ��3<6/9h��{�M��7�7�)�?�T)dL���?.�m�x�zW��oj1��hZ���;��aY��#L�$��"��m��C炷��2�k��1�{�E��n��7IV~_=��9����<��<��������'�֮�T�)I�)8ɷ�{�po�$շA�fK���(�p���߯���=S"���X���5������kNv#0q|�C=�h���[W�␌���ܯÃUg�:���f͗�Smu���U����/���/M�ч�l�ҁ��K1Yq�LD��k'�^3��8�!�����Q<���� ��O�>qz�CV��݂�át�Z��?΢o3�����EwJ�?��n�HF�*��av}ʩ�	�l�ڇ#���V�m�W��Nx�5����ɭaUNdl�)H� x�w>��)JL�|gu�Ad�����y8�/z���#1���ߍ5m��sx��;[�	U��o��\P�	��lV�O󾨔���L.D^1��km�������>"�:v�p���~��G�
:nF(�I+� &��p�1\��[��I����8h�u�	
6�+:�Cj� K2��_6�Ę�ًg��TblEhA"4(}>)C+V%+�*�mj���A��z��@1���R������,WSv���N��c���n�B�{,!�]��r��_��aL�x':2>E��\�0>ʩ��ή�2���ċ���ᰑ+��`���9>�����|���wQ��Q��Z�F'��к�Y�>�
�����A��h��⊔�#��HydT~̃�����=���BC&	M�w������`7��0����$"���<,��Y�`���(���}?����gN��X��;�l��2?s���*G<��FCP=$\������Ɣ�W.��c��	�A���$y|���nz]@���8��?7h�}--��A�	����EF���fr��#���=#M��0wC����[v�Z�:� ��I�yO�F	����ؔ�4Φ�	(7^���ܷ���� �^v��NR�F�P&?�^U����t�'M��䅵�N�)�qL�:��@5܆Ӂǧ!ͪ�� ��R��E�詉zJ_����lc`�D����5�����i�Y���U(�[,����p�̪�i�r���Ci�f����zd��YgW�ʊ��F�)�5��LӾO�_ ��BO��<&�
ʖǫ��/�5�Emy%Ҩyڟ��|�h�g/ӇL�L�OF~�O���iI��Z��9;�C#eb�/�PbE�k�L��A��j�uH�X� �-��ݷf9|��.G������RD�7aOe��x����\B!�a.�<�?��(a�D�Ŕ��G�#`Fpp<������;t=���՜�}��{߃q�/�s�%�������8&���x&���)_+�#S��
�^e@��z�Eh���_ZC����u�1�n)� ,G1Kv$��9��Kj���c��V1�޵�\I�k���C������aބ�(�y��tyr��b�� �d-�?��J�)8+?�w��3�k1e����� ��R�vr�=e�^�%ū�\<���^$ō@����m�
ݽ�_��[�֕�[�:��>q钝`Z����X�u��� �S������`�^l�^�p�����lgD�\�В���䈖?'���(j�ֳy��D�z�9)��:��+���R�-����AB_n��پ��8�z>����DB]�
`��C�uC<D�
�EAtX��T�,_� Ɉ�h����?H�>`��>�Q'����K(R�z�g쉞{x�'	5tLE��?�Iy.�F���Wq���A�7ϡ,�Lt-{6ź�E�׳&_GVs=�JORPPN�Q���_�x����\���Q>���d�ڶ>�}Ɵ.�ط��$��%���R�Å�Q��4>�b�Z��$��W�&��<M���r��ֺP`�O"��;N�õz�nx+�V�A#5e|�1dRI�Tq��{�x+�������h��!u�l,�f�j�ȡP)�GV {�Bw8S\��̟���9�mb��YI����b��_k�'h'Q���-��Ҍ�BYgG��I�����l���\��͹�V�n����A8��B|7C�{�sp���:5}����ZKԈ�\?t�}k�NV��,p_�� ��]`w��R۴���l�o��3�Zi�w>#��'≪�*���o��FV_�3�D���1���j}�?�D�V�wO�U��M�1��y�O¿Ժ[f)���bS6~yF�����v�������>�F�ٕH�B��op�䙗�{����؟����n�M	�'f���N<D7j}!M ���Ko���j���B�k�l�����*���K9�)�ٴ��8�CNT��a�ъ�1��J�Ǌ�@(X8�x�Ӵ	�H�?��X�#,�r,���S����'Jc%>(�̂3����i�Sa~)?T:N���N�@�M��{�����~�bD �A0D!�G_�*�${j�o��νCZ?�Q�J��	o�O���B�+�w%�v�1d���$+��Ȱ�l���"h��{���n�_Hܡ%>���g��i9'���tw-�q���^���1Q�ަ�����\^s�Ȃ�tM!�3���Gޑ��<�/8�O�������i��G�_�=o,�\�o�������=t�)�6� ��.u�-��mÊ���Iφ:���9�ݭ׬6��]=��/F;&�0Z�%{�ӗ���ُ���_��) ~�d��k(�C$2��ߞA:�J��9#��SK<x��c햐	gog!��)'P;&��6.����d)k��M��E��XId����a�e9M"�Dy�L�n�%��i���"��{p@~��L���p�;LC�O�cO��_S���2����@��:�8p ב��MR���Ufq]�0�ɱ}�6){�A3��������s=ɓs��+���b��w��L�ӅIS�� N��XnLES����6�ଵ|�/��У+$���xw� �E<�#��ǽx�������Cç����Ó�+��ʀ_����NX��8��J$CT���k@��L���@��_J(��%y�����S��fT��	�Gj��GY%[4�_�K�gRakҏ�.��߹�<n�p\��>m��c��j�Ȫ}��`�����3�B_
�����<�x7BV�6�~J��ЋTLj�l�:�z��3#��\����CU����r�Q���/�:��/ �t`��z�f�J�	���Í�Ya�4J����nU�nA��qa/	f�ޏ`�~@�W!��\E�1�e.��������.=շCe��������d5c�q~��� �H
���ݴI@7��oj�?
S�6t�@@R333���'��ϥ��B��o�_e$����`�R�s*s@��k�g�@<��o5͌u�e�Ok�8�Ic�~�GaTQ&
���L����O�����G�J����6���/b�T+	Ai���� )�>�<r
�2#�e���M�>�gF?�@�SW���1��
7���=��"Ӓ�wE�X�f��o�C���ƴì�^ n\r�8s~����`y�X�A@S����:��uu��u'D�P�� p[�7�w?e�	G��n����s��*n]h��w1v��3��k���!I�sP�L^�,˵��������NZ4��^�wZ��ޒj���2&1OZ�)��'O��>K���[cb��eh�E}�-�m�j�pqpb=�hCg-� m,έ�,v/�B��)��V��Y�ɼKj����ӽq�׌@�XrT��%'�����J�w�K7EJ#���]J��
�l�j� �/�7{'Q�^���vǿ(�I���W�0�1�"��G��KDh���՚��{�l�� 3r���3Fr�U.�+����bƲ�	����R�9n)�ă��}�6x5R�0J`�g�!byh�h ��MMn��a~�� -F���O�k�i���X��L�Ɏ��Б^s�J9\R���@R��_��%�<�ɪ���k��x�Ѧ���G�6���L2�:���V�7;��'Ѧ��VZ�h�19ū��5)�kl�e�
� goN��V%<���V��9��`)��\c ��|O�4����E(gB�Pq��\�+���?���-��jU��}��/�V(vQ�<4[��.7I���M�؍�Ō�Q�����(c�j�����5�HQQJB<��b���	��g3MV��=כ �F��Hc9_>����H�f^i^|�װ��_ǳ~v}!jY�`�F�S�H|����T���!4��Z��U^��)!%��!U-�!��%P�6|p9��0���L�>e�M:5- ���A�d���lGD�ǪF2#�v&�����^�3}Fh�J����6T%;n�����6e�0�@�Ȓ2��(�>ܝ<�������á�`K}"Ը���m>PQ����*�{��	��ƕ�{��u��GC�����ٮ?����s{k*/�pP�;" �
�Biy<u�0��*Z����E���z)�Zj}�ܚ����ZѤ��nc�w�u�:��l;{��h{*+b�c>��W����pl��.�6����d�ʄlg̰1��B>W�4q1�P��,�*�bp����ٓ��T��Kw���B ��i�-�΃�DD�"*�r�+k{�y��k�va
n_�n)ή9��}��|�c,�+����a����p�׋UI.�ט1����3���a�@ft'^��j�%t�Fi��-�^[	���S#������
�f ~�Fbjlv���o�t��;���,Q%�v�C5��us�F0QY�1)����|�j C!��ɴ��������H��N���rd@]L�Lk�l/M��V�Q.����֘�Ŀ�ᢵ2~_�h	��KJH�;�vNt�(�T�� ��#����k[A�d���5����x������SK��84 ��NS��r�J'�Gs��p�QeJ�Ӫ���m*�7ca��]/D.;�z�kYϔ�1��V�*���e��b����gn��������Q��0�y��qƢ+��y�}Bȫ����Di85����:��5��+C�x��j��j��������-is�����Y �F8�w�\⒭��ڸ�iP x�ͮp�*W���W�PW��f�y�C��h�r�-�b����)�`:$o%Q��Q���G��ɋq�n���G�����c�D�l��8��{e��߻���A�\h��F\zG ^<l��Z�E+��x�!�Q5--x����c�0�)�$�k��]�	�Y7Y�r����V𕾿�q��Y��U��YO	\�C��L��4s	X�I��E����'vaC�j���T�������C�ޱ{n����!d���z�nl\
Y���2|l@�����rt>R5=P���5qi�� P	�HHf߽���OQ4M���?,���X����ZB�sT~�A��ƃ�������-*���Cg�s}t��vO�WWI%�ktO?�W���>�`Y\��s�	�
J��B��%f�%Ki֙�:!��C�R]"��2�x���M)#�[�
Z���v�b�NA28���h6�+���kPR�p�/��?n4�^��H� /!�ߡ�3�曩����z��#��5���P���a(�Fۿ��e��sQ0��kN�쒑r@���7HǸ��D<��N�L�n$���4>e/������� ���t�z���߭Su���<Pr�cX�~���ǫ�H��I��OR�iA�B21��ĊotV�g�o���eau+�)j=�sgw)�L�Lω[!N���.%�XnE��3�#Z�}:�;܋H+t�é�(�#j?$�܏[Ȑ],���ξ��$�������؎5��3��nq�S\R��<�����P���Q�n�(��6�t�ݚ���0<��N�r%��i�N��h���vp���}�쎤ԡF�O*Tc�s8u����j�4�4ck�f��#�e��S���*D�i��D��\).�l� �f�ݡP 3(l���P$eP]�O��d�^��P~+�%kn�A�@�������L�dF�h�S$ˇ�;\�r�dj���+P� �M�E�w�ZI$*�A��V<��-��%(tJns�F�����g%n�5�f�E/~+U������ܺ�"ў��fkB� ��/+��(!�a���-�#h��ٺ��x[��{3%iN	o���HC0���?��#�-`Qѯ[��/d�+�#4,ٌ��4z���쬧K�Pt�j^yD@��ddWcVV�6ಐN��i��Zz��f����;
e�ZN��E)N�S�P}�6�+f!��*b� 7>�����Q�x|ό5*���u1��E�]AA@�U�m n�+���	�a�e+,����� &��t���k���t�h�.���SS P�=v�z�DA=�@K�	K����9ξ�`�q��&(sPrI���0�	I�s����A�Q�T�hҋ���շZ�@��*�V=��|A�*5��"�;�Nx�&�ش8S�����
0�/o6�;6୦.���1^�{�JmIb0팘�G4C�??�E��ݐ+�f�e�Ue�Fϝ����Ib�aN���'[W!��OD�e ��6��=*�l�-h���`����lo��HC���ak[�%���%)�@ �B��%����i���H���1�,q�Ӓy'>�'�hW�Of���j�ap��7���p��W�;�[+�榵oX'd�����g�"8���o#��ѱ4�����}����HVd��9#�����=�hh�[:.��Q>���5�fC�eL�³�4`��b�4,� �(k���]�S�Z�37��fZ��� ��z�Y^�D��U���g-Àϗ�]�>�K�����2}���G�	���Z��|�;���N-F���2~w�@�8R_[�/�g��e����t��j�2\�����,j��|�q�9S�Sઘ̞���M�5#  h?I�H����s�߂�֌��>�|�᛹�۸(Ny]5:G��z���g�w�l�RP�I�8�<�PA19M��°^Z�@���2�	~��Gw��Mj�>���Q#�I?\z�����Zu�A�+}[A�［+ţ[���8ˍ0��qZA޹0g��2	�͍t7x4s�������B���g�𦧘�Ѽ�
v�l����5_�������Ϣ��B~`ⶌ�5���N$����nJm����ؙ��(3��s��y�4�3����T��i�|��	T ]}��r� ҏ�� �A�g�@^����U�W���饇�2B��QW�l������gR�5����_w�D�������徢�) ���ЌҎ����[[Ş����YV<I�Q�fk��ݲg��~^�(��9�d$�39S�fm�!���N�N��3��PXEj�t��O�e�u͘o�y���w�V�E���֧�t��LX�μq�Jڦ*]�ϳ	�Vh4�+�DG��Aiz5J�ٸ���~ہBI&��Q�4`��������C8櫶x'�һ� ����@��V�I��'�����DÂQ��W�)��m�EZF[�#3���F.+�<*�	���(���� ��w+���i�K�.6��%Gu����H��Qn��ħ>����}��T�J��jQj
8������D<K��ۣʺ@\2���~�R+z��U����g4��!�\�7L<1Ʃ�l�6��,���c}u� �?�m��bJV�(�3�Cܣmr���N�~��郿�� X�b����.�<9����@r
�2�S�(�!6��&i��x\�w��>o[����G����	!%�Ȱ��{V_G�v	�����梕��ZM���fޕ���OНuL>f w_��5.���fY@(�y��	5�|%��L� �\c4
)b|�斑��z����3��qd�%30B'��W�Y�B�Sޅ�G�_-�4L�=��������1����C�XW5��X{&�
�7�K؁����<2�k�ǃ7p =m��m����is�A��x�����	��7n\�$�rMũY���DHS~�˦��[\�2
���Y�ی�@70I�Y*6�m��<�^"�iO��@#��q�Muwp� q�p��҅��HBxr?s���R)N�!���Ǝ����	���$!a~D(� ~0N���W#K���!�yW&��0nq����=�1��X�hQ/�i�&�
Xe�#�'���u��L�,j��<����ݏc6��n
A
`�%������_�u+p�OaS^6��F�40 `ʵ$[���c�x������4(�d�
�˹G�a�u~�T�;x�ư��B�H")M;F�a�D͘L�> 7V��e����~6�n�^�z[qһ�Aj(ˣ�z�PF����Cs~g�ދ}|�Ҙ5�V�0�Q�ch��c8*�z�	��.�rԜ4�[AUf�O��s!��u�:3s�Ƕ��Iܐ̢�s^f��"�ЙqXD��ۺ�,1�7�6��I-��_�BK��+��"���z�æ��6-�qw�9F/�06�Wͳ
M�̭tVg;@�e��Fb�A�t�><���>���#ŝ�R��킑�C�L_h"�d���-�;<wy��)�	,C�ooI"DЗ��<���Ӽ�qԶ�A߀��'SՒ�^�:�,�"��<g*��A�Ė�.�?�νm\>��J���!� �ر	��̻��v��"w���zv�\B��xkvo�Lb=~��+^}��F��+vd=(><��a��G5���x/&��G�����=�<샴rᄄv1�����6o��2�݊�ْ�Ԁ�G����"�<ި��wM�4oE%$e�DU;�d\�^�!1�|d�.��,Ģ�k��v +m�/��L--ؑ񬯳��g�=;X	{+	�Xj�=����n�.�6/�C��	�EIHs#��>Y�daӔ<f=��;\���!^��@�,c{�r�7�RÞ;�WZ�
 �ßg9U#?����5�ď���e�����#>[38�5���	.�T�9�_������kC�{���<jyz�e����s���u�`�n%�O��!���?ف�3[�����|ѕ2�_e��k��E��Q�L���(�o�7L�AN�O?�]8Ǉ<���OukJ����7��M��?,��ꌹ)��� � ���GO��s��_{.�W������c���R�Ψ-�K��������-8�fm�a���"���������E���
���w�?@^"Sy:�q?$���di,jz�@����}�c�����տ`H�Hi{�F��<��o�G�H��v����-_{��I����u2���N$;�Z��m��W N�� �������|�z�������ZZ	��mn�����3J���S���4���C��	m��V�~.%*����0Y)�刻��6�n#��!Ũ_W�Z�[{bL���1��r��!���\�W}��nLB�*�	ϡ7�pM��eHF�p�.����9,�*�fp��T5H��&(�x~�腷�H�8��>E
��pJ�w�8����K� ����ޛ