// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:27 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XFXsHTDwbHLgfClXGe0nmJ50Mf8QBWSSd1umy+K3svjMarGc9xH5uvFqDlJ17bSg
FxSQNWQQD10hTTugMFW09avF3YKEn4Du37Jrk+gGDcfVJ+VHouKnKmdGeZsKiVMu
048GzFxF/fP6vuzXJ6SNCeN+xJDG8uJdJEbNkJGpUNg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5232)
5gsj3mtXDINSQEUGHXS6I43aLAdCYqKLw1wQShDB+ZcGdV7POX4vU25dHoxAFTeU
JCmy12jmfXrPrDNedKrA2cPIIxkmTOk5oqphxVfyDvI3lWM6oO34s5NxJsoqivWm
BqdgwX5GskdIzAXgwJfDubZwwF4V6mt0SFG8KlhT7d2U9xkNxSUm2i6cKn/VmaiF
YylTD9kKqn2AbrfbI+BGMjWXxF0fW5TTEzZda29xSZ20/xiLx9ijnSfa7/SEfc2f
SgQMJBOX5ZTqbqsVWsAg5X/Ant7OgmelmAMm642Z+R9kPaiHOTSgjum4GTiMlorf
dLyspE80cgTl55s1a5Xn8iTWkEQZyJRhWCKpLRNhZgiiksZMajjDn9upjIlA2GNF
21wxVGn5aqXMSiio5DSvWjqooGfQcIhW3oUQoUghKXPDbiWtnwTFDw2SdhiwKxJf
mJZtgMRjvI1Iy0igBSaw8Qcmfjx+Q93LolfDRoF/qKVWM/fNnuT+OG5XqJQsWAO4
Zq6+e7qZD8efjkN+EZCOwzhM2jRUbBBOp6tycDEA2Jm7agg969LyeHWBUXwGzBqc
en7UoJrowNwo1rG/DTSmxaskgtPDWLLMkU70aEARX5rCNGpuFabk2gZtk4ExhB0C
OdXLM7yfrmuA26KOehu7HaLkHAwYLX4dblOU5yfsliprRD/tkFH96I3N/4U45WVV
rDpmqbmEREAk0X3lYWb3LMeOYwkQFhUJ0eRLkOuNCgWprD1BkQXxEOH8pecKEqtP
uaQFAqpjtj3LQ8CPJOFUwphXBOP79V1aQgKE4EjhY2eoR5ZRxyD7uObH6Hq7N2Cw
nUunvX3cKz5v+a+zv06/2TbTzFPRIJ9zRJkwm0xq5J+4f2O3JgAn8uZG9RbZnq6N
BhWdaJhfl+jqnZnlh3fvR6nvrt0b1y2K73muONOI2/Ify8vfBqNFGCrYnr1shHM2
Zkx0bTaHDUi3OHjz6lqWPJlAXXLlEd/D1CHDp+wE5TeZ3ze75a21HA2l10wj171d
IMdhR0nctKc/OJT9BpghbqfM+xkUGzsh+pHX0h1k09gGMYK1QF8EgDUml5h6yQMe
NqqtXNyVokIv6JsP0hattSx7IHB6UoU6sa3729o1qO5xTNsnl1Cv02zIs4sPymSQ
TOQf7RQGdngrKAs9M1uTUGIk2frNWVQ0mpvvnoXVaeSiccA9PSpEkAjrBYP3rSz+
q2qdr58UPjWW3wdQJbzf88CTv28BJpG1NAhacn1mM8e4JOcD4gikzpGvtYUigbUd
OtKm8/cOtfUmmhYciN9uFuTTD4jZ9jmInsP3HZk+NvHwgTwUp3EwE93JHgxqyvhz
wtVvPU3T4+JZleqewrSxPOyErHYl55GQkV1NA+4NRfGcErEkX2FAGel1Y7/wVxyb
UQg9b7j1vsnwqeHYf4sTHWO+blfLo6wFWcmEe3ZH2S++tLxqVJN+Dt6DPDLPWbNf
SVKGwB4Lzod2ZXxUp93m/okA0TY2wCn611aLD0Y3PlH/Qqdsni+e6LyxPGs/ETKJ
bytL49nfPNmlcJHDjAK99Dh6OrbwS5tElE3xPZ7+4WpiBsYgtmX/abgu8ZpxibUx
5YmP7bknFLIvkpj3QAV7TATl9IVnU3d+t3NzwX8Qc4FnRM+mW9FEjZ9s0H3oP/9O
VlhvnSSR9Fy814N6XPFMJNrJd1WTugN8hUhQr7ugFxlPwp4Qbfnxhms1MlkkV/Qr
qt1i596hfAc4uQaRIWD+qMP35Rkn9ANP0RUnjuYwgK8INAufq31CgAqUtYHXflMf
W5BfHShCLduJgeSCE7aLsHZD9SUsl9kgVb1aHGQ/knJXpjBk3BGPSxFmXOU2sPGA
SE7sU5KzRuOTPA/wLirQ2LQCsB0SVkZF80fH1tVg7O28B92Fq2njx3BrFCSCFVeo
atj7aFHFM3IH9NWyW2zzG5LulhPa88MFlW//W+0UAAbllCaY+rGGe26YANvPbZHk
z5dvFRZB4EKUGkZp1MuhKSt5v/X09KgSCB4ohS+qlL9OHJoGB4eq92ywRb9N6AL2
/BmdNIKXcmduqR9QV6S+/b73IpPnMjtz5Us5MCSQGpYDBTqBk/l7sJfzqGn871V7
9xFck1302gUOdMh98s30BHyMb7OjkYlo2KjvSGki4/02WwYCoMGUb3Jo9XtGWOJp
G83RdlHFz6PLaPSE+RLa4iP20Xzz4xBhFShxWQ2Pw2hPtyt/Ypw+nzGI8qHdF8a/
uKh1s6kRw43/zxl/FNSf2W3M3y0wyPDTrAGLD0h81vi42Wapds7g1OzWEtT8H+c8
7pdH+afzt5OsjejilvWkS03arjyNRDNwooWk/z61JeP9L52EesyInBbPUB3nFxr9
12Y/Wt+kDXYFOzGvVL0o4/1V/x1/4RI0eqtTHMpSrQSu8hRsE9DzX2vJ3rsfT3iu
WgLEesO5GFebpBBTPQQ25vhaNEtidT3a3F5K38RWffJ2bfG01r4657bbgJ2qon3Z
YPHv6fjjwZoIBDnN5ZH4rXaiRqc17aqDHAaz+4GZ30zrqYM5XcaQsYnmw8wq07jb
sFWVt3h9Nrl9AnoQDjRr4u/u/o8OyTqdnZvztHgkwhOJOmDm4dc7EeY4kLbVsaqu
CoNrVbtnk8QF9g7Tfj3cRVDmMfjDrJcKTin9I8xtOJok6YzCuW4lwwTmy1NX1c1C
qhVeaW2vPv3io8cc5JMc44KDTqeCNSrwYPzQbb16MOC3anoc/Mu6hPppa9fuCY0d
wHXlWhcITMl2+3+Von98PQqLuP/HTUuPh01h75v5sAo+TrBZyVRvNQeqIOWuQMoj
AKtIwvkWszpxW/91IlO3JY35G75Lu+jz0tln6IDDL/1MeJ+uBkC3Vm3AsBIWjwM9
tJHS7yujrh7+mXU4ezfwYmjKf7KNp2DueovKrbswPBa9DZPPYdb7RkgF6gQVqc0v
iVt8cbDi1OKb3cHAiZrVPPi67tbmrwZ0QDMrzw2S8IEK2AqtsU9bwtoxix9VjDwC
wNWWzKU6LgkU0E/xF+EDZe2mz1ECqRKzhx/7JTRecYyltd3JHbhHYoJrMOiVBINb
TmcuRIZnceTFVu6BotzesBJ0NovuKKPvDl0fuPGNwqtd908BklvfYj2otlF2VTmc
OfM2W0woebP4nDFxy4ULuaLZUzznxVx5AvcixhagcBOcMhn5EsQA7b+yyAkoe965
I225UIBLEIa+UH5lebuswUxUPkYAefxHX8M5huPPVPtZPub7neMqx510W/6jsMfO
BBFPvFlnMffAK/OGvNq5skF6CVPSi1Y3d4dQlvSOCMlRE7FABUAbQu1hoCSfavUg
wn6CBZqmvIkc7uavgkut2OHmj4d3XN5a3ifbyP2qqigcna8PfavyOmeXVcZKQJ1I
26oyzohK9VC+sn7Lev/q8WM25SYNjfmd+PSlcLj1ne3BfD3gKI4+7zzAG+pDRk/P
UoDqc+S3VY5Ap/1XQaIa+UznIWjUCV/fhtzHIVM7FTMUv5Y1DWMDZJ1Hl8TKojAV
di36g8Ae+eZZ4dP7r+1OK9gok9VQ5CuaqKH7RoVJ1cjXX25ik2fwARK9Zwia7V83
P8rczdEAC4DCLfGWPmuySoBqiYGa/aNym5mmve1zjW6SzgbX5Fb5VdmXLFxjD8hr
LdBFEO5Jea7cXkE0YH/RK5UC4xtTFptF6SA7cJPt9zPsuC2qmD2xPCQGIyrQooFw
MlnOV71gNVHqsikVZGOPha1FBgFjpY9NmjVi8nrkYk2PzCVMk/HyB6NEwWB6nLFf
xlmamSgbJohXgv+Xu4WJnZZZDqjho+CkE7yfJpXtasFt8hrvT7QRbIp3NXmCOahz
9oL1NwdmKsA+SXSR/ErA4WxtksL3j7eItUkLFNI8s7A9e6hgAdWELMtXtr6xgz+n
rzWaXz9VPh1BQmax2oo2bBO5j2eg8wbIv0lOR48N8bRTMG4lZCnNxP9500D20H0K
j01/nsjethTm3+U+y7uhu6GO2HdHUTekE4AkFiw+9uXIvO2dJQnpksHe6lcckZ++
ujpbFwL9qJbXwequQC4WCoftKY4DBKaFBzN8wPexKx9iYRJk9fWLluOudsqwUpEz
EUHK8KJquYhoQLZB849BqgjMUxAO/z8epqV4Q1053Fu9RvDGyGih9x8d5LNw8zsR
AIUGYEsD5KfhCoflPuhHff0PdiJAi34EU4b1eBgerPueAYrpHl/Xgx9sWvMg8771
96XefD9P6ObgMsRDbEUwxv2GUBZkXgCa58LFPbADt56n7txTtcDnzqEiZJFRZM6m
ofjqEiuaA2eIML4n1tzuYQzff9s5QloqXErKYSfdnZ8MQ5d057sHwxH4Gs2CvUQt
4QkY32ZCUr5X7RsRsc+GOw/yOPxUTylTkRWbjGRKz+AQ5N8UXmsWNkqPjFza99pg
C8XsoCDncZTpiQ2IM2gtpm8PPSlR6BmUIlffLdX32jq60KkA76AMxM/Kc9SNjAu4
VBYjNv8eiXkD5eSA7WhohgyLgRtF7nbT1W4UFmITq0x+dtXXGzXLLUZ8iXvj8O8Q
injm5Wh9KsriTRDTMuqZKCWRTYG5o/DvBcpE1VWowokftsrZcchz/4ugmXC9ThHT
k4omU4km1MWA30nj3tqVqkGpftxU2J1+LNoyuapUdk4avhKEVexQhihHAeKAL47R
goaxmVc5WPW8i0/QPthhfHoZibQknQhVKX6lGhfx2J8WF8dfC3wwbYGQw449zlL+
NCD1HQpU4bE7zU9QV6l2YyFogEYsbHnyWaFQEguYgN3iXdm4WCUyjfhtCSYnjTjg
zczVsHodg3TZEd7CDrFZEtC4bRPuXoYyvXGqoQmtljE4d0tz2b++rgkFmCvoeDN0
g+cqXZzKRFwbPDlSYQlLuA+ZkiAhICjx5l5QSob+z4CRZ9IMkPghXOZHw3Ap+mS7
rbS2ak8VtDKEptPoZHGLGdwr8JJEOq4s1eyJ7YsND655eO22EsyafGnTs3eVKP+x
p5xEv6KEVMOlF/oBWxa0Co6QVZks70lGnyrL3alMp4fJHMUJ0XfK9/rwSe7Jlvpv
cd70xEvwXyL6/da3JYGEgGT6S9qAU8PNq3fAhyIiMZuueC77qHiNxXKMldcPfUnZ
4T2D9GsJ7xTk3oxVbpH/8VZNKGRBogRwFczJnqlcE2bZLy8oPtMlsj2l6QjIZBdM
Wk/Z7pS/ValeWsVwTQmLoXCZupMcMz9GCbN73IoLf0du5ji+iFFJa4C2rfG+8VYv
I0ebHUTbmbZVyb19xwmymZz72ZGJM+8JIeHjTZM2yLy3uu9By0+V9cuuK5eHdnK1
QLyt8ZxY8zt90tYWMFIBjbEdotxBPl+uote+iUUWLPl7rr9a0fPCuK1k+k2c+3ot
ENoRqYzYseQH3xBcEo7D/jEWdX0MDet+o0RHE8q2pNyw2wpJCn0CimIgbWqA4BCp
wuL4ShbIoMBklFnjrdAWQHNT6TcN3eugD/wzu8NhK26QPg4RzxJ7h6wTCQQxekf7
zRFKvRHmmfqYHgGpMtwG+i60kdT1MQtKYnZ3q9q9o9AGoo4yBJ1JBo4Nc+RILkuK
CvWHt6aGt/IC+7c+Wzo65/+9zqpBzHqSfp1UZZsAxlxy38EnLtFJV9M5+OVUU8K+
Pi6ItPRLQHWJTCIRVG/XK5l1ZZKm87p4RimfrqnVqmza15ReywPMVUociTBbth3S
eg7hdp1Acd7fHKGkeNV2fA7SGwp3uzUkWyQaPg/hQx8RDIx6y4+3kdk3YjtMq5Y3
UpLUZ1k2O4631RbpY2cmg/L8AoQN9U7ZpWYZXpMDKtEi3jDIe+Aua9+zDkNspPzO
261oNBOdCOLDNGBaH024Qbt6A3kZWouB8+LmfwEm3eHUb8HnQXeccdNYFFAa2KF7
JkaY1uv1PcPAolzyT1mmAzrT86ZBSO0WAmPbSdToxdMA2mGO8OaMqWM4HdK8PjCE
ct8zb94Atgartzf+zzuI8noDrAK1n2RnTew7zcMWqr/LTjUYnSZS3zE1NuXwQH2X
Subp4NdyDLORwpK3jgDUR8ezB4kejUiS3I7AdftnUTRG5ASCaNbE558UTSrm4/ad
t2+br2fUwyaR1k5pvsp+GQrM7vPG4Bh1EOeKfSyobgP3bP0QGqIIveuEtM4k09YK
lzc1kd9+CVyAtnJ0UChhT7IxBfWwo6I4j0CY0Fuwqm2JclH9mCHcjdr7iKweqm1X
6N7KWYq9QUv/7mXMMrkQt3/n4j20D52lKp8KdKZxoSXv62+KrwNJo1mkP0grNUGO
i9U9Dv4zgmb0dqPFAajMAR9OzoYBMeneebC3s9o6cYECusfj7fAoluJ4UT9wNK/t
gZUG2SZTCj88vFBW/jwNPPWTlDUM69lb+rvRPrtjCw6DOJzO+K25QEWlrL46hwFT
xltiaMUPy2mkOMy8ZNwmeNYjnemspZ3IhnIWQ9qY/p8GC1vB7zcv7AQ4y8QtIrEC
ccpHy+IxkVjP9fNO3SzIWb68Q/sBLtXiev88rF2C+D27XnTBieQ8BM6ctIdDvCRT
7lHQ6WCyrML9+HDTNsKt5EXdY5Z7ZkLFd6ZzMmP9gRjZdfnieMt1e18h0WQdp0NB
2cNbt+mALjNL6WJ72dYUjRtai/MUj7ew6pfpujPfVRtaHvts/I0cVZLCSrFg5GvH
BQfFShpfg+/tLEPMWDuuzfHKxnHgSKBL+oDayYdCq8aUQoEvIPemaVltZM7YON4U
8ittRx/2D8FMAbGfMK7BijL3qZkRpPtpOlLE9CtZ6RkA4V2qTU3XURFJm30Ugscr
Eb9ZulY3gBrOnVDro4lH2wCP8KPG7pIz66KwuN1RndFkfsOH0JZ6r9OjPsMx5ymG
1zIOUqUuVmj3FuEFvSiMBHUM7jtAiP7PhuMyi8r3hDzc+utekFLDGHQq4EOgkqDX
scSCqNFjh6HN2cZOFHuFdit/h9UJySq3U4vbxJ0QQxvVzPP2Ti/8vHH51sm8c1qv
`pragma protect end_protected
