��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@�ԍ! �AoH���;yE\�U�S�r*A�*�脼	�f>ߏ{�Q`�q�8fu�(���
�Dl�#_աظ<W���KPYra�^�藴ٽ5�Sc՚�Jhbkp?c��L�QQ\}�w�@wS�eB2��v��P:�c���w�o��f��L]�Cl*��Y2X��R�l������fY�*|M�	3�r_�N�t}�"?I9Y�ϯ��d�Q헧���H}�Ce�U4M^  ��
�@��xhuМ�T��UY�M'B���J������������T��~����R׉b�x��w@�/���N@ㆍ����\p���	Z.s���ڡ�v�DOB}H�`r������ b���%E�uzR�%D��z���_#�{.�������j�X��.�d��Ԩ�a�	-�8�V�ǈ��p������V� ]�W����+h�f��� �� ��K�p��q����$�{���ɼ*�"�\��	�!O��:u!oub�R�³�R�Y/t����xL��Kt,�sR���[�Ig��؊C A#9(Km#�&u�����u��b��b(���دY�I-��8��/M�W�v�%bϧ+���8�{0�G�.��]e ��|u'V��-��U	���8�T;�>q����X=�,WaS���3/2h���_6��$|�&�aF����V�{��-���.��n��L{��8��LaP�P-S�!�B<�� e�R&�������Ƒ����%Đ)�A�"�ےbo���k��m��d��n�*Q��v)�Jy�~�L��.e����j�<��+�'��kҽpr�˚SR�}$��4��5������<�㸸"��i@=�*j������P��[�&��-�俿0��j�<k���rT�MB��$k؜��r=�m��mbC����s���<�B_\���r�]+�2�*���y����;�ϊ��-���t�n��h��?\0@�4�k}�͵�M�� f�oΥN�T[O�I�J��
q	H�i���5(�4��_%��������/����O~o�y�e���Ƅ�yU�XK)���读��JWh�&�_����xI.tNP�,�c��3A��'���\�%v�;ʖ��,��ZV��G��2�uP_�aB�,���bTO\�����-<r�� ���#��a��q�龱�2���,�{����6��1D�͎B;���k�ߎm��˙4'&"=���9ٴq�r����2�U�( ��h�TM� 0�������]���!gNO��\�0;˛�ȥ{nܴ�	{�LЯ�}�Y���X�w��f�V�>���L�+����Q2����sIse��瀋� �ԡ_���Oi���cV���:�i��5: ��O��R�Ab9⛿�M�D��S�q|�	6�3w�h �v����bǬ/X/|~r�w��ɓ��-� 
}1*��C����m�����[h�q�	�g�m;7���Q��XP������E#��Yڔ+���<H�N��IHJ�a����/�"m��x��?�Ri�&�@?��*ӵ4㗝�=^$b�ҿA}}y%������RFS%���B���g�&zx�	ݡ���1���t�l��,�~�$�S�U#��`��?q��-����N��:;�^W�Z���RN4	�a"�{kY>�Qd:�p��1�L�=qw�'�*K�Roتx��v���j݊�U<Uv��͉N*1����n=7W����\�&v�v�`uiց�b�G��:�8�T��2������X�}|�,'Ñq�u�[�ﬢr����^[�0��Pࡱ��`�*�=HE'�		9x��@m���Q�( �A_XJ�8��Cv-�a|�و���Vi����_����C�`q���_R��Z����	,���s_۩�Zs�~!^_�`�A��۴#x���WL:F�(R%���#�kvh����j��0����暟�Ֆ��c.��o�/N��N��E��3��1>G|.�� ��b��b�S_��9��41}�ҷS�AHk��oGI���ŮVdC(��Im�G���*�)���sN�~@|���/��W/�F>5��Sv�b�&�Y�`�>������.���h$\r��Q�]h��Cх�Xh�"�C�7�R���;����u�$���	ց_8Q:p�E�s�>�1�̂�6}��24��ً�7 �) �He}����Z$����E�*�8fSn~i�v��9�i�[��|�"ȷ��8�x�����\_Ҿ0�����uxwo���'�N���� �t֣�B���W�]6}-��Ў3��t�Yg;j)�.��J�H{-�����G,<b>~W��Nu��J%�˒Y&�Y����^85X��V�~��j�����ֱKIޓ�"@�QG��u��y��TĿ�9��:o�*��Wx{B�8��Bs䭂)�[�u���#8�U���9��+�E7��P��ES�����ԯ��ro�H�_�^J�o��4;E�X���_�<��T����UR��x}A�U��I����G�/\bm�l��hf��xGTݎ��W��"#��������
��$�w��2=e��7�H�p2n��-5�E� ��h��ոO�PS{&:?@G����� ��%�f[�)���躢�2��I�4'�؋����3L-V�ciT�̏��� .���<[X�ۀ0Z.I���e�_ox�D�ܹ�{��}D�%o��9<���tN-�n%
I�