��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|�p�v���?��y>����d:��}$d	 �!x�;<�c��"��4j� �xNd���^g�+b�s�lws�{�F���tBKѿ���Xd�k�9�CU0���������k�g�5o�S�G�e�wc��E����T�	�]e�S/k��ޥs��M?���8u�J��t|)M@��䯻�/��#4�OdM���8�XF�D	䎖�=NGR�8���ӗ�u�Y�7��M�{e�{
�R6�T��zw벃�?��0��3*����.�b���9}P�ssa�p����_���� '.��ބ�4`Q��]qUC�Y�/I';"�{�O~W���U��)�����-�fG5C��)��b�/�	!�	���~욤�K1�2bbEĤ��`EL봇"�ҳzlN�W㟫�n��{��E�&T,կڸ�� e��6���Y��N�Q�q�u���5!�����@6��H0������Ռ)ݓ��i/9P!y�x��:U��x"_��yY����b]��NшҬ����cw�ZV���K���q2��V�T�myV��~�>�	N�5���V��LZ'�E�1�}R��TS�+6�mU�t�^z���j�?�F�#�I\�h��_�ہ�٨ ���̗��+3��p��X�P��n� ��p�,8�W�Pt����Gr*\�qz�72K�ݴ��Z�Z�|Yq���sJo�����?s���7�՗��IǴ��]�>�j��IZ�6�&Ρ�{-�r:�!��b��X� ǩIG���uL}�s�	���R�(o��~%�&�h����Y����MK���[��Ь>Qn���/��W-�k���+�kA-%wih�d`>��$]C�O��r?���W(tZ%%ϼ�dRpIa��tB�kp��Ci6z7{`�G ��.�[�������Xpd����q�������/�ȃ;� ��R!�O��K8ج_����7f~�r(w�*u����9Z.k�I(r#9.���1G��_��610�� p�G���ǭ�C	C��J��L�	0`ƨ��N�`j�.��Sc������Fa���ߚiم�K���9+:S��L�0�9�p��x�VG������N�*�5[���مQ0��:��1��|�e�s�b�Q��j���S���X��|�R��q9�l?�+� �2ϛ��e��f9��u]�O	�$�0H�\f�5ցOY`�4�������i�I�okO �>rC�g���r&�{�s����$�A_V�3�oA�_R��]�x����.�Dg�QbF]f�]MC�A�J�z#��q��44�y�ͺ^�SwzK\Ԯ�b��.����|�WE��������'Xm� v+���3]�L��t�v���>i]�F�)���IаD��|!��Zv=@DH�J�}�t�Sl���HQۏ��6~�K�29�x7(�pL=>�����u���y��O?��u���
���XI�����e�����Z|��<��@N�B���dK�s���Y|�0�����H���-���6S����+v>3g?��a�u�8�1k���t՝�5� �8ؾ�T�n�T2�DjD�^扷>,,��?���m�B�fP٤�h�驲o%Hۉ��_-� +S~_�j����m�Rr(@6µž����ƹ]/���Q��)��e2�q���Q}@(sZ��\@6:�̤* m�����Y����U+����0u��QP����x[�����W�^A�OR��O��r�qG����6��s�`�@�qZ�3�����ah�RoѺ�@]��>��H��|���>+O-Y�!����(�������J�ڄ��+�#3�I�@S�)i��j��*��XG�T�emr��
�[��h)�y#A����
��#	I��H�-KU�p��M)���yN�=R�Є�P�W���T�ݹf�j�/���Fذh7�r�����`�v4���C�C��*�Nq���=ZAS
چ�0��ȿ��&�d��r��&��k�8E4���k��������l�0A�u�}&}m��I'c#&:r��vm� 9���9T:��]��}3v��x.�ի���秱�-[9�C�{�(�(^ZQ��n���G�^	���6��3:���d{OIF�;-|ȷ�?�/����д�����e�K��ߡ��^ݬ�)��i�5%?ڞ�j���� 1�N���O��k�GS�Y���\�
U�^k����>/����y��[8�@C��w��=�����e��4hW�qu�^\MU����Y5!�VK
�
bl2s5N�%[w�[l��� |w']/�x���M~a���W���o����7�f�%�8p��ދ�t����H+'7=�>�uM��r>a\����[\�=4��2ޜ�´��fV�'kz���J��:���p�F�k��{�鵐��ͤw����K��p���jE�C�U�9v���	��j`f�������QTD�;�@���>�-���>�rv��83��\gX���@��)�o��gnL�Zbf
#�`,�ײ�76uu�|2��6���iRK�֐7��5�!g,���>4�!��7b�+U̴xD��FX�x��������$Z�N�l!������+7fv'�_?%J�ڴ��k�X��"�b���VJ�1��*�I������i�>9Hw�s�B�P6эE0jdSF�� o���ה�~�����h��R3J?���e��b�\����]�GE��X Gkw�)s �͑�@><�Y��B�SX�����;��q|M��4ѕRf!)���2�ƿ`��0ِaE�X��qE��I���2l��,*��?H�!i
��;��]�sf X��)1�تp����[(a	�}�X���8>d $�4�s�\�/�-�x {?������]���c��H���ЅReh>&<v�h�W�H��x�I.\	�)ؾ���:�1��^�U�ߢ��I8���Xe���+�n ����Ӣ!6�v��%a�ۑ��'�F?-J&ٴ	�{h`w�wF������C�F��ּ�Y�a��9�[���ur�<�&�,�P���@HP�X��y��,Ҝ#!+y�+4�Kl��L�D/>o!��$~	�Q���J�
��2��k��U���ݻ���}~�kd��^�3�����*���j6mߓ0m<k]���^'.�/$�+�ǜ��]?��nh)G�)�	�׼�X���zsI�������Q/#����K��~���]].]C����T-Dp�1r%bPqCH��N��3������J ����Ռc���+���e)�ly��\�s�ĝ��8#w�׈�9��d����;��)`�j��L��z �0���#�O���W���!��d�/�~̎�i��x��t���(��Ҙ*�T�Qhytz�pJ	r������r�\W�)����aT�Q�ƎQ��[(�0[�yW�<'vk��8{Y\Qל�lcp�������6T[-A���i(7�F72ќW��~�������T.a��ۏ.�/
�nv�sb�ݍM�U+�7�̄�m+թ~�B�H=_G�u�g�7�U�	��~�9V�Sv;��fEѭ�"�R��O|�@Us��%�귩�om ���� �'5���e+�$_�2��{�v��n������.�D4�O~<�������4�9NW E��*�0�N't�WԺ*aV�<%?����H:�����Vz����ʛ>�������P��'�3��*�m�3���WfL*���E�[����w�l~ ۉ�Ȇ����d�bjT���F��Gʅ��)����JmT/t�57��9��.��F��
��ܳ�Wg��+��\2R�6�/���ȉ#0>�q��O���v��
K�y����,Os1�����M��r ���������ϛ]5�|�}�_c�Ya;��S��seR�!���f���.}H��� ��({ ��b{���mF23�+��Ȟ���Jѧ[�z�5��犵�Ts��h¥u�~EX�9�-�����H�q�!�c�Vf�ŭ���t�bﰯ��������pݙ�$�����w��J��C�J�����@1|9�O������U*x�����R���2�2��!�F��~��Q��w%<%]���Jg\S$r����3�]9�ng|%㽹����j�~�Ux��H�v\5%S��^5�c��np� �����4n�3��zۼ6�Dp�~x8��m�B��>��K�}��Ma�\s��f�;P�����D@�C�L+�Wߑ�2YM���;�D�]~��@}'��F��`:�x���I��.^���F�	D>*�:�G:�>������Ib��u�|��Z�= �����+B�hp�$��K�}�3ۚ���P�h"���!򝝮�O`9�f��5���!6]p祉Wq�������`�2q�r��@�Æ�Z��?q��ϬCl�@�綟���Н�&�h	ݝB�LGo.�&��[�7���/v8fa�'�����3�����p�Ae�����:��:cO<�f��ד��VXi�U��I�x��,�4z.-G{�&c��ٓ����n�8�x�g��gͰ��}��1�EjF[�ӱEU[�7��*t�P�̘��!��V���!�aN暔엷�?�.3���U���E-���2��V�x��V��62׵�ǔka����#�V��΄�|#�l������k���d
����{�}�X�G�-��q�Ƞj:&�W+��~�P�2-R6��Np�>�L[�S��)�Of�қ�n'��/��ꩀV�4<�0��+��z�e+���TB1O+f��Wd���_O�:Z[hF4��>Ll{��<�~���&��z��ك1]W��E����~T�xeE4�w^\���D���ݸ);X�!,����7D�\=W����I��� ~����|+���ْs�yW��l8���a�@N�ߜ�q6L7���ԇRa�K*F�}t4�c2�>������:6�,�l��A�gq�7ok�[ڽ�=�b&��<�!��D2���O6�@'?e�C@�����tt��0&�,����CQL
��L���!����9��v���m�
�`�d絔�C��ήH��Ei0� ��K`�.n�F�1�nO����Anix�����,S���1�����w\D��ҫO�t.d&¶Z~ㇷ�T�J����,@�vJ�7bekE����xO��k���\��&����/U�a��\rMc����͓\1�>B#gU��`k��ww��k�N��Q'�
�ͦ�=̷Zv� iX|[>+.���!��^l�ό���b�T�EEsr[g�߮�1��������v.���]������AC��f�J��$�?�LokB@��獩X<r��^��nd�[b��������_���#�aR솷���qPV|/�`@Rp�|\��=�����&7�Hk����bpV�yB\�(�d�<�F�_oN��_�̀�l�>L�p�s��k��5�Y张�{O�+�ܲ��_�G^A`�i�3�\/�C�ǈ��o��V:���1A�U�Er�ג�,�}<m��M�z�j]/����p�E{���?r�C^g�w!!Z�g
D�x��IE��u�,��-0颜��S̏�390|�}"L`^?J3]�8+��NA|!|R9��q��鎝�?����N�3rC��|r6�z	[�؍=�����ެ鰶��ma�fƯ���_9^J��浦\-�Q#S՗&o�j�����'�nP�7Y)��Ը�<���9Q@
���k���W�6 Ű��(�޵�� ���� �2����t_4)�Tz����5w�2X<d�S��\>3�`�#���~��}Hi%���~(V�H�B�*�ΰ�F-���"���$k)zjL�������T��_F�Bq�S�"5��
v�f6A�sU��g�BVދQ�1�t/���⠠�UR0㳫��ož*�c��Rq�cCw�(��%�NA�F��#����Jh�U����@`�'��Nc�E?h�8���\�K��:5�"�v�u/��2F�.D��T-��&��S��Jk>]ڍ��ם~�5	qr*���Ζ(��|ڒzW��#?Q���u�O�)��ox�犮�i�����'�E�k3�����mY9.8²��'��`��a����#��m):ᙲ�Q�$�U�c2@�ViƐu��r�t�0��/�k#�Yv�R�@M�V�Y��o������R`v��Y�n�?2q���*���Cr�G�������K����m��$D�xC��x}Z� a��k%�>�֥��l|K俘EB����Hb?�V��/��N�7%�b0<s� �;-�77�ؑ~��TY��`�"H�L
!��A�}��l����(�֘��^�/���6� ��{�/~�+�h�H�^+��\���iǇ�H��:�IK\�J�SV�,l��q�i-���>Ja�=�X���T;���=�ȝ���bɷ�@ �R"�ɷ�w���\��ݲ\>�m���#��p����IV��:�2���I�����[���C�_m4 D5c5]aD��aow/�d���t7��@�VJ�	,��l�Z����8�����> �؜zj�dnQמE!Y�D_�J�iR�� _���}`z����X�bPJ(rI���`���D�t�7�@+~K��jq��y�7'3�s��л���t��q�^�g���d���v��k�����S�����Vh�ov�,å��`�Z7�$�#���+÷;å��s[�D߄�n���+5꧔sW���6
�!,�� CpZ��h�H�S"B��E/)(&�{���9��ώjO��?������6�eF0�>I����ЛS���f4�Y�U82vE'z��Kq���&�Wa��aKI!?�@��b �����eO�����	+(�i���������<�3<NS�L�Q�X���~ɯq�p�sZ����������/Mb�{��J�%�]rMD��ގ���=T:�B�	��HT^	ؽ7���.ݳ�k݀i���	�	���uM��#hFPpfGfE��BC����'�K��]L�;ٍ��Y�V��g�)�T��3U٫��M���6�ϟޕ�\dy�D�.��uP��X1,)�3�z 0q�a:�I��MN� ¼�L"^��6:lHe˞a�]����|h�,#�V��PPj?���)w���bNؚ��'W���r����F�i/h�����r�]&ώ4\�`>���>M^ia�����}c�v�DBB�Y��+��@�]l����Wp���;�5|��\��j ���r���(˿���]����VYYi\���>�/��\T&3��1Hgt#z�z�Ͻњ��Jc�A@^��T�@<�i��؃�(?v��r�$x�0pcXjt&��L�؂��,3W�=����b܂�@����.&��i��.����f�fy����10,Q-Y����
��S�	���L�"��5��U��np�A�C>s��oI!�f���h��K�6�ʝ����j2R0��k�t���R���p�qɿ}w�N��)#�]]�	��3SK ^!��f�,yZ�y�(r�|sX���[���l�_bF���6?e�*�'v��K
$�r�2�#�՟%���h]��Yq�����v��M
9�@��z���1�{�XgqB�0\��V���Hj,p�\d)�,��|
�����hg��/dx�dxX�)����L�������J��@˟G�A5�w��)��97D��(�GU	i:r�Vo@����k�)�R�>�Ow�}�?�&M��YH�87Y�
fsY��-kĮ3�x ԶY{
��u"9�$YaY{��gk�b��Q������&�6Q��'-g�礧�ZBz��m�u�h�oD�w����Θ�����n8��6(ܡ��c�lJ���a�j����i�	;��!b�؝z�!�R����2D0�r._@�nZ��V&'{���@d����Ȕ6����Ɲ�iZϺ�t��e�^� ��ϪŇ����NK�Zٓ�5�)���8��`%;%{���0oB�\�|l��������D#_���2�}^�ev���A�w�!���No��f��d8�?��Y�;��o�;��<�r�9��1�3��riΩ�=`viˣV���E��	�㩆�)��0�;O�/��Z�0�#1�����-Nd�?V/��_���
�T���������w\��+��V�]�s�Z^��r��w�OX� ;L/1_#�`���!펚5���l38�|5�
_���|	�>U����"�X���/�����<)"���|����Sh��&/ًo�}�ËY=e����������g���T����������Vx�q�2.��A���06~O�/������t�`�Zȹ�z�(>�#:a�A�/ں�� ;/��Y����[�5g>)�\�$(6������?%~��j��U@`q 4d8�d0�ڿ�m1.\KBc���ri�/�KI_��t�P9��l��"��^�>�i����wЗ��g}҉����Z�3�v~\(n�ު�qDd�8v�e��ʣ;�#�����"9�����.	���WG&@M?^6��J���Y�b��`�wS�5�����[���d##a���ԕS��ȑ|=E�5���ᾖQ)6�A�X�K����)u��lZ�d��T�T�1Q\��.gW�����W|���&�0%h e�?6U�lO^��2z^�>��U���4�DO�į���)��c�� [���5��|2�sß�4-W�͞����YWY�Dj�2K7]|��ja����"���HZ5UM��i���`�!��*Rr���Wիl����l�����h�p�J��z�^wy�
�!CZ��#&�fR��41�����4�f��."{��*(,�]�'��Ӯ 5��#�l������I�)s�qq���]OPC����o���2���R)F��UD.o�؀���q�-�&��'�_��*��}	��,���.��cN�z0bc��7��zx��9����k���o��C-<�|�q��F�jή�4ѕ� w���ٚ}6�������ZD��Ը����O_���6�5Ʉ{ ����?���fe�{�G�*t%�1:�&M�V���9��0�"��e�$��ZQ�G�C�R��;�N�?_��(n�����)�O��>�3FTd�Y��%��}�:�
��B��q5)�s@
�= ��GҴW>���a�i����l^M󳰁����vgڢ^���p�a��
�?�E�dD0�hw4��}8�! r����"0)���<����c��@|���qL�{�2�3D��z��:;�"JM�P�s�q�v���1e����g��ƻA��+�e�B$�z/�ߧ��.v��YKaY�U�蟵���.hH �W}oh���k�Ƨ{�J����ǣ�?����NM1�@����P�+H7�=�m5���wݞ{��$�(�_�.�>�$�\����m�N2*܅�(:�Jxk��6���;�7�O4E�NUxM`}='���q@8`������>�:��)�����Q�K
�1�,��ܪ�]?��\�ޟv/bl	G�B�� 4��,d�H;q�!-L��e0�ӕ�k$���8K���u��ps+��>�d��Uٚ��6(�b8�\޳��ZcEZ�b���F�0ỻ��obM�9������~�����[pq
P���� o_���V4о�{5���s&.�%�5�����(�e.l�%ڷ������/��c�赜+�� H��g
^�G-��4p5@1Q����1��m;K��$͡���H~���߿�a�}�z��boUv�h�<r^A���,��͝z���T��G�Y^?�Ah/�{����ˬ2"U��E�ǥ#E��(�>�1N*��3@Ƞ;59 �e�*h�,�P*�m�ª��{�A�'���ȱ٫_"��}�'&��!�R5�4p���׫�].S�k�2N�IL���+_BA�	�x���[i7�Rk�^��C����2��Gy:�aʷ��nd�h�{�g���RAu�G�#����ڣ��,�)\�I��i�� ��H���1YZ�F_�w$Jhآ�tٛ�����0?���vI|�n煕��*Ο�+9!�H�e
���e���,��R���@��]DVd��>?�|p���Pӓ���l6�l�6�E�~	�p��|�H⼡�����C�BjM��Fl��n�-��g��{��� O�
�C��o%da��|����/g6��K�nek7ZlC��-v��?�n��je�����5�K�<ډ ={�昨�Tm�h<bs��� 16��Q�u���2sC8�����1�Wp]�J.����A�٤�/�E�T�fe$w� L�?���� -嶊᫣�ȃd+��I|W�<}�IQ��2�Z؛p��z��޽T8�pB�AU��L��Ǌ�|m��qb��r��r��ߐo`�������z��l�ؓ�����{���q��[�����F�}64�.ڲG�������I�[&�?C,��1�h�an���h�M��b���2\}%B/�ً"5���u	�p{M��)� Ѵ�gwl�I�c)�������b6��܃G���큭f�~�¤�cG�k��뉔��ǅ�ޙ�%_����%`�x� �2��z��f��2t-g���=�������2��n(��A']ֹ�q�a���{��]2�)`�s*Up1H�޾��+S������7:.����t�p(>�����`�0�˸U�rq쒽������ӛϫE�sّI���Bd�pЛO �$� &��ϐs�'�}�ɒ�:+�G'�s$AnG���8��+��L�B��e=��=�'�nGA�r�T�貤� r�;ϸ%��s΢�8���=������U�Pb�8���b����b���\_����d���Rm]"!�d��%���UEA����#���e2��yCg��M�r�U�>�p�C��Y��p3�#��)�3�fO7!�������F�l����֛7M'�8�Cflr ]x�zf�Pj��J�oT��f�i���5��ƞ�|���zy)YP�<CNs^�BH|��l� �6g��B
ժǻ�y����u�.Ou����h=�<�g������zg8�v�E)iϷ����-hc�!�XQ�	��M+��_>�`��.|2�LNclR��6iKڼ?�X�_ܽ�
ҵi�v��W��6�(�Y��/u�5'�񍅑���5AU�Y�ȹ"�J���*L-���_]g`��'c~��8����󒸐��*�Q���ڄ���|�@�r�˥Hݖ�I���T�U�)�m��ʔ���dɓ+��,�Qa�$'���3�� ���%Q�|c�kq��4n6� ڟb���/�b|��p=iX�B&�+�1��2����5�\�8�����g!�������E�%$�=���Y�-JsY&��j�wI��񷒇��xA$b\�=w%�)�L����6����\&՜]ѡ�΂l���!�k����V�fM����Co*��S�֖kU�	�A4�3�R���cv1f�̸]yK��4��q ĔpG)FE^��3���)-��E�	��P]�;l�a�c�x����I
r��N+�'����ũgI�	�@2�q<B��[������HWĖ$2!���;N�j���Rg����f6�e�z(�`�j��y�c��ά]���\^oߟ�&f��t �Z�B�7y���NK��b���[ĹKs;�&+���Y��q��?�Y2��^�N�7�;gʦ��%��3��a�"8c�l_��o�¿�
���.���� z/}�����(�1�M��q(z2d��F&�A�0}e���y�DF��s�`�RL\���uc�D  �s��
��6[�(�����*�PH��p�8�+_p��Fؤ�����m���'6��7�%KQ�����N���H�eYpZ͏'�d4�FȞ�<J��]�g�·:��6�<ʀ6dEĎ�0��6e�d�M��F��	�7�A�͹Wa��D%-ٸr��`B�o�O}�~��C�L/�C=�	���cԞ���Omr��p�!�ѕ��8�2�����7��������n����������� ��s����;ޣRh��I�dMS3�g���XB�L:: ����Rk�{�?��.9>� қ�d���'�� ���#�����@�j{f#�`�z���߲T��^1G�~����"aI���}(��v9�Y�Qo���_��@؂� �kdL�N��,��D�U8!F�[�  ��@�dU�#˞9g�-���ܝ���'8ٝ
s�X͟y�p�֬�2u�y�I�
?�L�nJ&��¾e�it\����D[N�q�ͮ��o�c���D��2�@�%,T$˨�W6>�+��BxR>�l�;?�۟��6�����y�NA��Z�jv����`��s[��\�?�"jL&i��~� ���eX�� _�Hy�/w��1���y�$3��<���e�5r8)v�<f�w��2��vEG)Xm���4u�v��)۟!��]��ش�R��;GyR�[�@��w0��Z������/�ɃWza���Ҙ�EBrz�r5����.��z����҅��<��$��<�$��T8 �y{ &�jR�\j�RFXD��ZJMA�(�Cbp��/�24̄pu\�ɷ}(o����^qV�h��Nu?S���OFS �.x:a[e��>����~a�6X3%�j���i^�����,Fq�]�+k�9�'"p�K��I�;�k�R�ۜ��4���k�C�6e���P�q x����%m�1�oD�$���0[����f_��F!E�@tν>����%��7���6���W��0/�J
L�WY&5��=����y�PiW�#�C���U\�����!�$٭�g\�R3��~�rJ���V�5B·���C�Xvt�vj5��$�̈́��hW���g�k�-|�ҫY]�*j��PuPE��ю���\��z���~�u������F����'�zMK��{hBNw.~�����_����x8^>�"u��,��D�G�W,�~m�ɺ���1Ǡ��۩ʦ��2WB3we�P����p�nΔA�3e�K�����9��T� �����"(�Xi��a>�<�}��m�*���h�a�5�x�{�28ю�V+X'�����m�p���)���c�!�~�\a(��mU|ľ(��35D�B�h/F�/%�A�ZioQ�)�,T�]ſ�B2�Ϛ+��Z� �	iŞ�����^�2o�uX���?*Fƍhg�;<��b�wA�JE���z}�l���C�~3p_7	>�;������_J΅�V���|�:Gi�7�0��kپ��q��e�4*���p�nD���2�lL��֭��h]D�4��;�WS�@B�T�&����r�������}L`�n��vB$n%��W�[m�T*���;�Of%`v!D�ʖ���\u��.�e0���^��D����ba,��䚌��le�:}g�O�RH���\ƾy���x���W���5�<����+�e��C��n!e4�5���H��fx�sU�	`�8�aĎ�e�8�V�>��'�\+����/20�3��;��l�ش�)'��(Ǉ$5�[��}�5|#���y�[J�~��Ԛ+5�1�'tRd�1��������i�px�'jd����c#��O��c�o���3�x�Y���9E���	�����9Vš�i
����ke�5K�mb��m��>di�SQ��՛%������b㰧��f�z���!5ew���$^[���3`�$>Ks��b�q,s̰���f+�½_����~4�������6+QySD����v�s�!!�pT�漢�ǬJ���"�B+r-�����t���D�X|�t�z>�&�wcj �PRE��9��f��T�k"EҾ���>г�}}0u?+��Ƒ2D^H��|Gp�	BB\0Vr5P�U�h��+�WT��_�'V37�b-����XJ�a91��y�"X
�4�Ĉ(%	�R�A���T����ِ�0%�jʵ���9�9��VMǐ,��w���<�J�2�� ��Fl_�uc���x����c�{��`%3,+me�1��h��T���[ls-�����l�h�d�ܤ�.����|͎8O'��+H����������lS	��&5�Q
Ĵ�b.���>�XI�G[+��Xō���ݒA����{�y���'�m*jMvp���?���ɢ���:��f�е�I�},xT���5ߌP*l [<��X5[���rȣAS!S�b��>��B�[�bd@-�s0��n�8����]�|G�hfZy���0��taf�/1����0\�,�{g�AH�r��j�uЭ�v�g�M�����xB�P�ͅ�A�V�$�
�o`���%*B����nP>�-@]���1��+��9]��Uf-0�bx������ ��*��&WAC��(���FWT(��p�;�$2��*�䐐� ��?�e����a�~W�ڞ�~s��y�ш�|��ʡXy��c�E��(VB�C�4�!C�ft��8�IF������I��R��)ȯ��P52�{f©zm��r��n���n,� v]��HӲV���>�ʰ�}=;�(�n9�z������՘�k��=ы��Z��#�ǁ_V}��2z�Tj,��r��1����of��X� �����)�<���7��SY1�ڍ��^.^�Q�at?ώ6������R2�lF��C�H�-�&S��(�C��kс�RKp���4�d�C6�����q��0�g�>A�s;�����muE�i{R�����b��ɧ\�[�C跴���8�i������v���D�f�)��f�aE.M��Ď�8�K�ؽ�:g�d�Ĳ�7`���9A�[� ��B��ser�Q/䔫=YG�5zrʞ���gI� �yr;]?�^8"�=6��֏^`yw�N��D��NO\*Go�f��i0��ʂ���E�<eM!��k���)4��i�9և�0��ؿfq���}�vj��Ý�
�Ծ�������=ZY���� �gZ���q��pj��&�/�Hk�6MY�V!���
�Yv���Y���{��rk7d�ć��� sX�@eJ?o�7�DH`��Wx)��1�8�Iʠ`M��^Nb!��ZR7:��mn\v(��5�l��E��)([2"p��,1wj����?")�5pT�2�r��o�A��BV��É�� d�Ҫ�ص�t��7���f���f)��}WV`��,^�5�a����`e�g��W�1��aM"�C:���x���`U�k��� oPgǳ�d6�+3E.(����q�]^�FH��i�_*Oh�ԫ��*Q�b`1���Ղmo�Ǝl��RY����u[��3��Ɩ��83��3[IK� ��G$$\�4�X��-}�T�B���θ�' 
���<Y�˺�����_L�C�Pz�o�q+s>������~���D���̠a1I�
Pn�:�u���Yc�^��=�b�3�F&ʿ�ӳ��_�0X},��
�xA�+�~�<�JN�󾾘Ġ"AͅG��x�E�	�w� � mr���c��|`-�$��2�45���� �&����a��]��HJ�剴��~e�� b�=ٵߚߵ˖��땑�����Y+�&Ռ� EP+{vl6ب4\[Κ��_<p��X]ˏ��v�����P��Ƙ�_RoIx|���� B!��t`ܒCL��e?`oFҬ���#>�sCQ-�ظ�FL�t�i���Γs݃�G$�ڍa}V��*�'H4��e��e�d���hOU���@7��m.P%N_Hch�A3���[�_d,�mHʂ̶��3�.޷�g�F������a�Γ:/[�(��=�z�\S�T4q�,f�x�N/v�C�����'��І�4���ohG��I��Vφ2o�Π,䂦�rlIT#���p?�'�^[K��.5k>��)M󽊇#��a@Z��IT*��jo�C��w������"��2��:G��+p�h�W�Pe,���ȏ�Hvy�ɇy�U�BY�z�+	MRYIL#d��{��{�ߥ����ax����
M�A���=L
�~��@RR��v5�zP0��c�eǔcj�5-E\�����yɬ�Ӫ ���m7�<'ؠ>���*��po �o�w��>P7�3A.�^Wo� ����S�cB]����K��2�����]$�@�k�wR���9�y����/%��W���#�1� {��Xwj$H��⿖U��i�/����
��6t�A�gi)�_�o�֠�+�M'�zT�4a�ב�"�,{�Av��!{�G���{7�2�>ӳ�_K=�zU.c
��7��s-�ʢ���E��.�d������&d'�h���=.k��I�n� ��d@&�ш?�l�͟8���5+��|T޵H�N��7�θj�9A����(��j�r"a��7���:5�3�Q����3:�.�قAZ�b�:����#��h��-�K�W��;��/������l��T���"U�p=}�P��[�h_J�<\t�fy��*䁴�cٮ+�����5/&b�cE�6lU�[�+_W��#��ꃤ�T����E7��)��f�i(<��%x��.�sF6*^@� ���㳰��b�G �eg�����^���m�a�z�\[���`��Q4�Q��U���={�O<��[��&
?��|Ǖ��7�^��B��׺p������kO��;ɵ:��j�4��c���jFn��6�4�b�xW%��Z��8>E���,;4����iZ�vR-ÇnQ�4�3Ӻ��]�'enl�&ї�ǽ{2�-�AF�2i;X���TM�k
�r+K��s���Pf�H@�C����JsX�'����� m~����%$���uͲ�fճO�^�4⪿j�>�/�#}������~N�~�����F��D9���V��6�Uj����EY@A�@ d�$�|���K�K���$�2�AN3V���(TQrӵm�
R��k�k� ���9F�%���-	9�L2�
�޽rhQ9{h����� 6�x�(%ޱ�ї#���>iA�+yh�Y�7ҿ�>nO�y)@j�v��Ш�S�A.X��#X��s�~O,�y�B`��.c�5�Q�2�@���L�:���SΊ����b����/�
}1k��U���ק�����PJ,�ç5�;��	"���;�2g��s��g��!�Y�G ��q�@!l���=T"r�`���|�(���U+��Q��Q4rUv�E�Ц���F�K�0�j;��MU�Ad�Xe�v'��ǭ`��>�T���F]��:%����؜JwaC�˃����`���BG�X��WJ�>��:���x	��hr����Z-��B%��Re�,�~y��y#��_�glTW��2t�|qc-���<�Cݣ�2���Bsn�F5Coy�a���Y�&V<�s��4�caF��1臚�G�Xl.b�HW���ooN�`9?[qԺ)yt�VM�:,��8��v	O��$��F"�M��\1xC�����ܒ�6Cs��viJ��DDJ����'-}��9?��	�(d��D�\����B@XsS"��g	�o#-�X~��m��+ږ�0dԅ\**:"�3�id�����قy81��j U��j:�Sn��Gox��.A�g/ŭ�_I��~O,8q����)���JSj^^<	��,�4��0͛n�j  ��,��^E7��ez����u���b+ �A������,>L�A�5�Z#�"8jizI;U(b�sq|�H{ڞ�؝�>�<����QZ��>={	e^��/���o�"O)ˢF��<�'{3�[�A%�8��"ʽ�Id����@7G`'�^^E������ p|�O��l^�G+�RE�[K>s��m=��Dý����L��)��<��IFZ&{�8A~�I��1�yEs\1&l	<s�	��x>B�y%&��z���_2��8�g3�(�w���<�ݘ� {ʯ�T�H:V ��'P;�*NV}r���dq?���zȺ�p���y�
�����3쵐�"N!�u�i!� �2
����g�;����̦��p�A�����H�>g2���'t0���
i 5��Ĩ��;.^���y�o"y��qئ�<ǃ[3���~ѧ�ZFx�_���*�P�/�[�T�5�S\7�P�&�����Kֶ$PP�k3���Z�f�l��:W�Ʃ\��+�"�K6e5�Uk�s��7 Q�����?�`:c>�ƫӮ��!|_�*"|ւ(9�a��ԇl��ߵ��^�$
������Q 2ZA��|
W�2�w���oT�O�����������<��4�����w�G� �j���e�x�Hi��f�7�"`�~x��Nw�$�&��_�n���K�qY\��vN�e6�������T��h	�!|�+'�����Om���g��?�]ֿ�]��5�?�^��}��E碡)���;%_@�׍ ��Z:���]{ˠ,Mڈ������ň��`�
�BK~�+`�Xֹ?�.f�^|����A���z�QC��z��q>I [n���4�]0w����j�z�b�V�������`��cT�B�7J��E���[���j]�~���H�V�����u↡����B� �vŴ�w�=����
2���d�l���3i��}�A�
�w*
ڲ�}�N	���o�Y�684� ��y 9o�[�rBL��L�yI�0���/A��%;����(B42�6F״Ps��F �P ���D����G��	ܲd��3�(�u�ۯV��I�p��Q"�U�k��k������x�ח�w?�>K�Vi��OYGW���S�+a���x4���4���|�!:Ȍu"�PF���J�r,�I�3�P0�I^��%���ʣ۲����1NZ��7�=}�>õE�pw"��g������UO,����!�D�a�oNVȢ��F)�V~M��	�ʜXŠh�ڮ��.ֲ�^�V��SkH�,?��씼g�l	�vmq��		*�z9��F��？VN�bW�h����1 �k����Gi��s�2Q��w�թ,9�)N�K�9d�078,�.VS�/��]j��1���ʰ�`*��^=�㝙����e��Faɩ�Cbv��b�'fh�눒"��F4�J�>u�spY�������5#b}�߹�d�E
�'�2(��cހ��vM�Z=��J$ܙ�W�3+g�����ZF��6��v0��Ý����/���ZT�6�/GR���g+�<�.P�lKU�w�|v^̬|n\��5�`3h/���+C�y�Ņ���DSr��w���5�kO�+���w}Y�Pa��êޖ9�~[�f�F�U�X�#�E;�A�[�co��[��ZDmA�P%���F����B�����G2ҟ�I���M�B��������%c&b=�%��I�:��~)�S�{�u	O�6-%4��P��p����مo�1~�ё� ,�Sۍ�����a���>\���%[������M��.�8�~# s٧��~��V�ͯ8����iJ,D���=�E,�A5F���α∪/~�aY��
��?������Y*���P&�2Պ�>b�,>u3����^N��U~��d�ѴC��9�gBg���V��6�bS�DH�V�+h��X������fc���1Y�_D���P�x\[��L�SV�5�ׅ��y�l���=�Ҥ�N3EK�ux�!ހ���>g��s`�̵�yjټ�u0�J{��b"�9��k��p:aq�$��i5!�<J����8��!-*Ci]eW��r����tI�Ӈ(J½۸����S�V|�`����s6�Ԑ����;��C���%=������:@-v�۪)����&V-}'�/ZL[�x�R�2a���0E/��}�
.3=a0�Q�[n���%��I����pI���	>�Sk�U���I6�FK�8P�
J|&͌ez�?%�wF�̡L,�i�29lg��3f�)z�:���f�V*�%;��T�ycSyS�1A�P���GG�3�ᐕ8��W�Y������R�Ǖq�Ne�O�'>�,/Fϩ���œy_��ѓ�Qx�����oVȖTlPx�AX�3�=�{�a7a�\ '��o�!���[���M@x9�R�q[w��D�����9�ܴ�|�( PJ�!��)؎evn�;��V Q�ooů�0�-"���x?X\Z L�a�;���vG� \j��C�Q��>v	('E�z�)��w"l݅���e*\�q��hD&A�7�Xr��k������)��$3��R����(>�֞�f��)w/C��ry�yj�Y}0x���j;���\_ה��yu�������xE���>�����Q���]Y���bE�?��l�f��w~�4{}�k��Z�N{L您�<U"�jZ%�l���{K�0
��1�L߃lzx�/N^=Y�\�-LQ��)�u�	яr:m��8ũ��������=EwX�b��zi�d���)	ES*x)y^�[K4�y}ϖ�ɝs�� f�W�"^�d��/�O�� ?����G��
KjQ�v_kr���B�Ҳ���CR�J����2�zVٌ���Q��|[�G6���g��"M�w¨���ٚ���OR$�Wp��\λ�ӆq��D���*笊LIqɸUL1p�-�8�jn�7R����En�k��[N�c^?��t�|C�h�Wr��yMϲ�_�:�`�s�e�	-�k�?�҂&	���7ʮ�����~�P��|��w�-��o��k�W�4��s�=��p5��'�F�1VQ!�0��V�b��8'JƗɗ�����(�m{!;u�����E�Hh��r�[����R�7��涸]�Fc�zO����	ۛ�����d/�7hE
$kWn�/�(��@�f��r�O9�d� ��\ʋ|��f��
T����������)����f4�Fa���:��\B�)m�߲Eb�:���6��
��$�nL��H�cgY.�u�������R�����.����D�tV	�@����Axq�[�0�+�W��牍
:��FϽ�(�%gD����	���}��R�C��C�񾿲O�H�����7��=���B� fl(�/��E9��{�al�S�,�8�R<>v�ə]�"� ��CD��x���b[{�c�z����)l��'2�e�!8(�œ�![������^-�ԧǤ���G����Q�Jۯ���b�m� �׋d�%�x��4TbP�auaͽx'm�:���KjѠ4��ɼ;�qu���(�r�kP;t����P��L�<��)^��gK������"���tcv�J�[_�����p�1��C���+������0����{n���u���t�5��>���|���.���8��;�k%0Úu(�}��f�Juo�Zi��%���Nl�#�-�ދ���,h���|�9+c/�<�kف��(Z��>���k���-Z�n�����5�YO�1��J�U�ָ8�iV5y�`�y&C��%��I��.�!q��:��o<�~�,��c9~��K�k�I� p��kt3�4e~��)Yϓ�'��!��a���.�V�l	��m} �(��&�� N9�Ndb��})�͇y�q�]�꣧2=Gv��G���gd>+~j�"0��i��p,�Bۚ1;�]�e�o3y/Aa"F�T0$����ڳ�<I<�傁�j�%x�U��h���Q𠆳ؕX=�M�i��7 녎�5����b<�^�_�� TȽ3���Dq��SX� ��xe}��G�š=S0�|-�(�dg��)G?E�F�i�R5����m��_�e~��;��f�4��vIhJc��hz+�Z��7�Z�q�_P��5e�^����{��A a'�B�� �ޣ~�$�:=��ԌB��?VSc�i$0�@��}m�`��8����&<{�:BY�]� g0���_���^��>����3��B���4�� /��w����R{ҷ�D�I`d D�\�1���7'Gt���OJ���g� w�ԋ܅ܗ� :��;�~�S�p|�dQ���W�2�I]f2[3Kb-�� ҚS �Τ��o�����"l�/F�N�5�\��}�i�c��L+��[�NGJ3��Ih��DAd
#;��+�E��X����߅mtIHڐȮ ��UFR����)�F34��1y��ߊf�G�L��x�L����P�W��N����ZPb��2m�$�y�kT@9�[E
kC_����/��w��0z!���E�P�L�T9�٫�1����?gÈ��I�<�� �e�=�+��8%�����M`�t�#iP�K����{&��Yk�P���v��_�r�,++��/a*�0�r��
����
�;W��k�=�h%��������L��d����,�*Ƹ`�7�fmz ����"�U�4<kmv�3h#�4�s8��'��&
�����D�"�\�`mIK:v����� o�P�̝���)��Ś% ���-��`�6����Ti1�K*�f���-�� Z*��������Dt���h�泲7*}5����x�!����'*�4~� �=j��)����G��ߧ�n�a�.�x^�qwbS��j� tU� c�o��Iܦ$��j�C��.�݀tY�n�����*�E��wL���8�y�}�)(�p�7E���9�L�����ԵB��\o�K@j�|D*�e���f����E�R�#�aK�� 4-�� �fC�<U��c�<+	~�[�lZ��������4��JU��Vz�bh�sN�&�D��P�'��U�D�Yq:�6����J��g(�;�3�%�˥�b��F	';lTR
�<9(��70Y�����r������!u���9e�o�
ե�
kچi3��H��[��7.&��)k��<����r��x.U�R���g1v:�)�*g���Q���]����հ�tɾ��x�SWP�0��y�	EN�3u�$����\��_��MD�"ϹO��:CЎ���!�X f�h����\�X⿿+��A���@�]�3���ߜO��]eƀ��*ISEm�0��U8�:o�
����m��V!pGV")��[�,k�_W�0��P�V�Oe��0�&6�}U=y�pR���hQ>ns�nB�U_Wa���<��9�T�)q�˸��S��s��:���$k<�eY�o��Q@$�U��M���=����=,�c�H@�ӥ��oo��z�)��B�ݪm����Әc�]ȑg�[I
/�맋$�}LQm;x$� ��BA������vE��1l�S�ЧP�p'�Ϩd>�[��s���e��9����"Ɵ����U9)U�L ./�������/Gϟ��z'!�¼x�=)t�ˊo^҃���[z�h�E�qY�9�]R�E4J6֊�h����a|�6wDa/�"p����;��d�0*��M+��S�Ӧ��cdH�% s�4�(�rP����4ye��:=�����]N?U��U���Pӛ>n#u\�ymz�咶IMC�4J�!n�6t�X��:%>d��H;�`@k�m&(؁���+!��8�����2�'i�z�љ%
v��hD�Øؽ�5/�e�/���e��-�~-�fU��~�s�H!�C(��&�ķ���:��2yuge!}E�s��d��0�	C,]3�288W�
x�M�y�sD��D�C�m��ʛiꈹ���hU\ȓ2�N͕s�ԉN�j���Y��H����V'+tG@���?+3���W�N��/I�ZR���kG�"���e���0�R��-4D�"��u�jB����v\n��[�m���o7U<}��o�4��m[H�1[�k"��J,C9��J�����߇q���0a0L= �ri�ũ��>YQ���rh�ƙo+���������m`�K�~�*������mÎ�%�Ǣ�����,�F��bn�B����g�cH˦.fJ��Y��U�w�l���ڲ�A��WN����&p�C`3�W����?�{�)(eGo{�i�Y����K�2c�6t�D%1�~X,�ل
��F�ŋ���ќ��Q�"95��K��3u� p��dd4y�"�3�=���?� b�p=��ܭ�����5�6��v.P��k���:�*2�YAtv!�@�4��ާ����X��c��O`�=qg��7ˮ��=s �ؖ�+&�N�?�R�{�D�#�AbGw/��rmKYf��'��$���T���V��2co�D��e��p)]݊���9�-��Y�~d��:�s���q�D#��m���;��f}sn�9���!e���75?��qq���9���#�ȅP����w`�I,'\���gzO�Ch���ݮC��Z��)��c2,�%�(oT4��9�0�~�K�c�Jq��H�zY�\���S��P*s�ـ�U�k�z�.V@������b���B�3h
w	�����E@ߺx�	$���Y�x��aM�w'u��}�pU�c��D�<%��:-����v�v�!�E[)����r(4�+M��#��������u�<���a� JE��O��N�QR/��yI����k��do�p�KO+�@w���w�\��嘜[��%F�G�zCRǶ��Z}L�1�����sym
Sm��0A����lE�6��}7(�9�S�L�?�M�r����|h-��x�����T�_� �'�	m�Ƿ����ߘ��	s�ش�AA�w��YH���x�1yWAB��N�#��AW�R6)�%��Z����DOUH~��7� �qjS	A�_�;X���˔)n:��**��Ft=Xw��ls�@0��4 n�e�-��X���A����6��ˠ�z��vӝȉ���.�w�Q�n_=��[@�:����Q��8[d9Ǌj,oLݯ)Zp�<sJ�_G��Qb<�����2`'
xr���{E%(�V�V(A#�/�r���/���<�]����nz+��Q�Kɡ�Ԗ
�Y3����ŷZ���(2�Nt�	�m��Sf]����i�[d��b��="Ǝ�&�D�|1���.'dh�Z[�/�	A��[k��=u�H��!O��Q��z�.�texW�ڧ��h����p����A�v�L���E]��j_s��3���nN`����d�-0�ƪ=��a�m�ήl��j�"k�Z�B*F7�� �ߟ���������ܖ��L�sIJ���e�9���Z�޴E�*d$���ȓ�DΣ��P����,~^D�ޚ��GG3#�LO�zo�:LRck8x�$Mǋvu�y[��4{EGBus��eч�Lt���Yv꠰������h�[��#�#&ȁ��w�^�V�K���g���Ʈ�Ώ@�;�Q-M���[۪'_��nD}�.�x�8:^�J���F�e��� �Y6����S9�:%�S<��K%��*^��\�ս���T�tG�����B� =��d?]H�?m���29���զiS���t
��c�5�{�N��:��N�Im��j��g~þ҆Д��-�jD-�X� �=���z��N��S`���(C5eᵚ|#b��М�Ԝ���%���N��hbo��	HE
�<�s^�����t�+BWt�,ݯ��v,��U�E-���y���|�"4%������F�g*-	�-���s����f?YSx�?�Tw��jA��Zq���<��-�la�Q�hƇ�m2N��84�_�p,~^gu-R�<Gv|�0�?-��
�N%�*l<�¨��ş�n�6}e9�K�m	+g��%H��"�a�oc�?C��)�����0��k�I[��;�XY�8c�������6h�vڮ�An�߰��� q�6baV
nb������9��~���%�����Q��޶�0��I���_������7NX]BA���Rh#�ip����f��y*Y#�N�L�e��i�c4wu�3�p��ۅ�AI
�[�N%��� �{S�%F�i�_����z����vǟu�Oô#�FK�N�q���y[���ֲ�!�^4.�:QGV��(_z8��"��ݚ��f]��aCd΢�(m��˟���eG%o���ZsVt�9����UD�?C�Э�N��B|�w=Rk�}@�7O����<�t̹V5 %Fq�����q�˙0ؽe��KE�B�G��b��"fPt��d�c� �!l�*/s����7�e�˾~����G�.�5?M��\���=Eѫm�f!򵅷�!|=�1����o������#��3��΀H�?��R� �|��o5��L�rP���ⵓ�����T�����z�&CxH�ej�I��}��B�bv�.b�LRP^�� 	�aܴb;�mŕ�ݹl.� ő���e1�OS��1�.��`l,�<�"�?S�8�\��6~-�q�nط��cq�/7M<����FH$�e�1��G�E$z.�"]�Zˈþ���ƾ��`��8m\=��x���4.
m슑]7�,��Q�e�-��ؔ��H�mB�����I��&?숯�ȸ���^�vU���g?��T�9ꩿ���n\:���Y��U����NJ*�t$�#�wܱ�sƈ"�)>�
�A���4K�O��h��ϓ�2Wx�3
hZ�br0�L�#�޿5ppo��� ��Z���F�n�ЖH@5���% �!�C���s)-K��z1��Z]����KD���=�a�'o=�r�_�AXŧ����	٘"#�c�j�����=���Y����ؖ�
���0/N'̂�K���2e�&0ĥ�$�r6S��d�KZ@�O�G���1��6�?�X9ѱ��t�TL����`aJy@g��Y�?�H3��I#u2eu1�F��v����:����k����=�����=�.!��6���A�o7Ç\�LH�f���SB�D�3<�&m$�9�����Wu�,-4Y["a�d��Ɖ��z��z�Z)��:������D� 	%!V��G]R�=����z�P^Al��ў�}�{=��e�-��]���J�Z�ʹd?�gc�]h�T���u�P�_Ŧ�Z���V!�8�m�"��Q���N�Ʉ�9�-�A�V�Z���<B`�H�ya���m>d���+�3̾�x����ͭ�����kBr�Xض�p٠��m�νQ�L��A\�����K�������3��J��ㅷ�Lz�����-��K�ː�@��wZLa����f$�����	������>��\��{
w|mv��<�ܛ�'���hqґ�s�@O���,h{������-�h��>�����X>Dk�m����r����c���"~lU������ۭ�V،��j��d�\�\����%�{�gڛ�o�@��Y42�[����Y�(���=�mC�	��<1�Q�e{��!��_�C}4��i�q�g�\4~��D����	"G:J��k΋q����4z#f�WOm5m[7Q�&�o�5�O6L�B�]X�#��DH_�B,��)B8�\l�f]%��M�.l[',�U�b���Ѩ+s3���у$��ts�+�ʰF���F���煯�ϷeM��<�����[+(a4CT�e{a��sv��3���d�&�`~&����CB�#�;B�B:(�����G5v�F�le���'WˆeZ� g������Uv�������Ш�QA��%=�u��ſ☦���s����z`����RU�l ��Kqb⡠���IT�����[=�%�����`_���t;$ת���G�u�,E�����\T} ���,�Yq�}�w54\�w��{���82)r��F��9�y���v�Nv���FD��+⌲U�#���ǿ	��Q0lf�8��
*�χs(t����D9�)��+�x�W/�?�������Ԯ��<��fN��ñf�|�
�]za�Tj�qUE����2�����5��ώ��'	�E�\�y�I[�t��%MV~��&魋�-_h#9R��a�H���!q�����<��,)��֚�J)��y�������zW���N/��K��	�o	���#|����gw�2N��ma�m+���h�:|����~��b���F�;��,r����	�3�RǮ;��ljnT�rm
~�v�:�dz�\kCfh/E�D�'�����O�r1兂�. �(��HuA��/�В�2ҖIH���e��]��2;gq�&�H@d%��v��7G��Gv�1)��$�R���0���m_t~�a4N�h��{�����=P�=Kf�1]�T�f�-���
� T8%_m}kͧXn C�Wcv�
|&z�Pp��1�m�$����o���v������R�~L(+���U�J�oc�?x#���"�o ʾ
=� �9?�!	��LҽAD��ͣp��O	:z$:ëE&�m����>����e��ç�8�0?������!XO�,Q{��K`i]2��L_���0Mⲳ��Vb<����1\��!\Q��GG��b�?�S^�(���#��o�R��� ������ﯦ�a���B�2U�ǐ���ͅ U�k.:e� ,?�fB:s��T�\�e� �áҊ�\��U}K��.tЈ�R�'�~Eέ~#�Y������u I��Д�F43�`��+�٧kk��=6U
�`�(P�m~?1�ev^����Q�3X`��߄���.���ￗOQg��޴��T����T�*�!�\须-�HF"�%���6>�!�ɯ(�}HjX͕|��G �2��b���;�՝g*Aʾ�h�/czK+Y}�<�fJp�lLj�{��?~�N�=l�y�;S���#�9�&!�
:B1�+K51�lb�a�O�k@�O�э�V��Α߁��"M〺��i�HW�(�+z�A��bϒ�w�<f�CB��Ľz��Y��6ւ�kQ�܇3lN9Ԣ	^���7!~眀
���h*��~�8�vi�Os�E�3�c���������1�G�
�����hJ�K��ݸj@@�hH�0K�R:��(�r�n��:r�+&�w B �W�
���Y�ɯ���49�-�q���>�5l��D��5v�o�f��T2�L�ޣ�VZ���R@�S�!�rC��:'�GK�*�0м�.�����s:�Fg�m�bMm���3W�9�u3u�O�kU�b�;)V�H@*C����7W_Dk�XK"�����I1'���\���y���/,�����h��r~�׬���y������_,�5�W;� ��4Z"�`�U�Չ�$���1�:�=5���P�<g���粞6�|j��Y����tf�A��r��\�@�� ��.q�L��t�2Uc@���EAnC	!�[ߪEv$ޠ�)���ղ����p��%�#���:Wq�͔�q틹@�����q�`0'#蝿����89[7�&���ҥ
�ere+R���n�:v����Yg�T>vf�g���^m,r �Q��҄��$�u�>@�,�ՄE%�elf�f���`���Zu��x���Q�+��J̽�U,!�|�<�%�?�h�n����P��pʏq�4���h���5B�!�)�8�,�y�d�ro���4��;,��asN2��~Ja/n�:6 �?�y]��&T�7��O�̰g:�N������׎�ϒ�~��sҠi�%Y-���+������n��hPې��l�������urR��/w:q	J�#�f��$�|����Y�])�h;��{:��bu��{��~tM���f2�Rf�v_����rUQ�n����R��y��tq�w��Eq^+��)2��Z�&��)��1�+˿�ʠw�mVVS�a�Vfd֠8�y{����ĉy��/�c��0uU19(�_U�Ӏ�&�Qh�?�����]���;J���H@ӑ9���n�d0�D@�\}mU-�cǸ��3��4�� �(����M�'V�;���Ȳ������?���
�Hp�蘑sP(,���aɎ��2T]��2V�ݬ1G���k(����^�tl��ݦ�g��E4�T3�R���A�\�����n�_T@o�^�S��w��3�����1�e�aV@QB��)~}�h�W�+��"G
�����h�xƟ�0����,�^SQex��5�Z�Z]�SR��Lu|c�{{�%�̤�.{��܌��>�b6�,�f�tL����M���ʜr�F�Q;E�w��o��t]RV�@����4�X�05K;@�F��?�j���y�����۱b�|�2�$ӿ��MĄ>�	v5�w�KV\ZN����O����� Y�Xρ� E����`"���kx%�t��Lm1�f/�N�[9�n��iXx������T�ۣ��h���TG������-\^f`�b�\��<J��g�h�eȮJ�X�O��,�=V�M����o&Z��T�e����>s�bL|^��Z��W��ΐH��-|.�LI�����Y���/�W���ch�~��,�*�\��y�3�G�:kF2B�,,y�BxÖ���Q�kqKE%�r���d���U��K��N�
)҈�����뻿�����đx°�x���T'�[q�����5.j�!�x��T���hR�\�B��=��p�~�@�S�I�0��C�Rl�v��G2�٢����k��!��boǵ����"��:2y7Qi�ɁX[�.����3#�^7�ih�($ls�&)�2�L�k(XVE��Bu�b �K[n��Ĝ̍���ď|~�9��Z�R.�K�H���X��ܶ��M�mzgI��7%E��2�0m������c���w5�B���$K9-�͌Ҁ�؛x�2�6�)A��y�p�A,4��"���V�ޘ'��F���5"�����k��.���Ni����h �{���k�O��k4�=>]��� B?7�
�Հ�`��n6�IVd�
��w���UmӤz�c-e↦�B�����&�6��b/fO��>g���}tDri�� ���U\�&���k�F j#/���'0����6@�^�.�er,T2%q}�1�Gk�n�hS��5�C���	��2�<��=Z�="}n��vr;��9��d���R�K�����u�5k=
��ܧG�vD���0q�1P�k�&ć�9�VX�Wé�O,�4�Κ����i�2��3�"��Dҵ�6ip!v�ΖZ.��s1�7�_k���(zW0}ML'��K~D��Yfh;#1�q")��R\��jԬ�o�b����Zيu��]-�%^r���!6�>��_q�����9�r�'�z����\�n�c�:���<p^f�G�u@�d��TI�=Ź��zyk�-���դ7Mf�������F��Zs��՛���5�r��Րڞ�n�}��3�pVg~j�6��<