��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ又tY�����C�f:OY��(><Y`s}�^@f �v���z�S��IE��f��!��U&bU��zi�I$�E�B�Y:mw�Ak@�JNi��C�t�&ND�3���&��srd((�fEI�6������d��7q��
���a�J���k���o����Y"~cL7|+uC6�&��/DGQ���P��f+�		���M�X;2<�`^8)_Z������3��,G�z��z����;�t�S=M#vE��U";����`&h�{$�N�+t���]�I����
I�E� �λ�}5����$В�������ʀ��v�k��7|쮆�w�ձ��{C���H�xM?ǽ�'ħp�v�OG�� ,���ymc����#��בsb]b>�ZFQ��Z�A����&*ݵB�ǠE)tu�
��R�z1���in�&~�Z"�7�1�+ӡ{ L5��f�1�!K�7�!I�����e:'�A��\g�X� g@l.�+����$���C��O@���9A|���B�ݶ��.���N��P���n�)��eV��L��Z����������C*��ʥ�V�w��Q��E@{��ŕ�k��NYW�H��0!�D9r��w��`��_�}�-`A&0��������o� -��gs�w�+k��ʽ1�W�w� 4�P��_H)ᵈ��p�����vb��t�v蒖�,?�j�'�s��U�Ɇȿ��&K	�8���E �C��.9�������U�����4vO��\C(u�d=�Z6��t�`z��]��>�b��������it�����G F4&����"Ҝ&���ٓZ��i_XKȣ�W\��/I%ª}q�<��!�/K��6��5׊֫@�o�G9�/`[�N�a�����B���R��BA5}#s�NMAr�_����O��W�,��y�`8����������l7*9M�Y��G�x?.{�y�E� �`ѯSR�fv��8��-Pfi�K@L��id��� �z�!�v���ͻ��vh�[������O`����6�8Q~�">���q�6�OS�J����R�l0�O��S�a��#�ϵ�dqX�؜'��S͒�l'8�9�/;(��e�@3?*�./���4�Ҏ)-�6Ip�VI��f�U@���;�.�^�<���>dLu��v�;��L����9qeg�G1KRT�f��SA�p#S�aI���S.F;��9��
��#[���E����Q�y0���@��:�E�T�/:����Y�DDrMs�e�XӅ�l%49����[����]�F��ެ�����O��ں?t?�J>�s��(�C�O}xzf��OQ��lKT��+�9I˽�m����$�U5�7��Cf9iR���Q�"�Hp�#��Rm{S��t��/h�7?�>���	�L7����E"&�Έ����
+�(�+̳����m&���9���SAĹ0W�������ﮁ�� �;��ꘀ��dc��T=�SU��,�-�h:s��Y��e!�'䎩`^`�B*�N�xj0�p_�<�� .�a9��kK��G]�!��cf����Ɲ�x�[em� E([��P�\sR����<t{�V�*�h��X2�E]�����G��U?w��kŖۅC΁��N�hs�G�ˋ�_�F�}��e�����e��wz��c��(�1kyS��O��<0���r��dn���C��MI�e���]s�-��jA���k9���ɤ�-����?�e�C����Y��}B'1A�m��y��>��W�<��9oarY&n�z�W�l��eY��%��:��,�G���I`t8W*z��&3�j��������"�ۍ>c���^X+/ ����6(x���Z�9#���L��{�<Z�-;1�����V�4r�CYq4`B����G�Ȍ�p��ɻ�z�|p���3��ev�dq��寅c[؜n��d��ROԺ�V�uo����%����P!�UQY��4��E=`b(j"�\���ZPR�: ���͒�MDY100�<7޸�v�