��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~3��Z�������# ��d|��̪�����PAZ:�;� ��Փ�?�}�F�ԙm�-r)��]���m�V[��zA�?�p�,O�?����5���dk�������'�]��i!������&5E��PN=����x��ҤLh��c9�`���u�˄x�]�-SZI{�i�]y�I���򾃺�㎛0���PN@k����D|d�F�Ύ��k�p�.���'o��'g{B�n�n!H���qʢ�n榕�*�wYOgs���0-���0�X�:����*%3�x%i�KU�W�,��3�=G�-5�&��N��= �޶R<�#*3E�"�~�7��.��ʧ�P����f#8���͠���VDĊ%*�C�8�$�x*X��TŠ~�!q�a��ũP��{L�.<��b���Ai��@;#�����7�4�y6W�[�,��%Tso�9`P�������������AW)�|�|��%��1�}�,��Jw�s��wX��P�ӄ\J�H��:�^�uNPM�_mZ�(�	5��Aq��de�l�{���O#��n$��w�Ty�fS�wa]|�|�y
��	��g��iE0d��Ok��i�@�}4n\���<���߬���&��h��s`��-C�n��#���sӬ��U$�����L��4��䙓�]�3Y���^�^��s��C:x��=�q��(��`ٖ��2�hP��v����c�����/�F(��t�јi��v�SR��n�6�0ڃ~W�C�X��_���4�#c��0Q�I\���j��G�6h�����[��}U;6<��#���l��/�,Ew�N{y�cXv�����!�?f�|`��ɛ��w�6S�a}JeG���4�
��r��C���!���Φ�t>!��t��z5B�do�so�A�ŻrZ~�t��Q�6l/��/|�ɹ]�Y�Ú!aMw��a)DC	�d����@]"Fֽ��v�&oc���������7�';Q�ĺͻ%�x�����C9�Y�X��V{����_��pJ�Ē��U�����^���2e���E�#Iш9�e���A�W�F,�o�	�$����Kܰ��()�R�j^�)T9\�q��r�jēmD��B��s���Q�6i�wd�#��iňL�J�t�g�;ӛE�� .�
���CNTa�O�IA��G
�r�ZH[F� ���J���Md񪭄��#���0h���I@��
����UM��zH\S��H�P�L�5�Gؒ:au�|R����zW0��i�٢#��[��U��Nn�nU���9����6`�ܵ�*և�L���_-(K��C�s��e�j�����>Өi�����9��[�V���rp���g�o����UP��Uj��RA8�����7T��(��d��L}�/
��C3�u�NԹ �|���H�p�|�X��.�!W�e�¡5���ñv�-�� 1��R1�-j��\�a$HS*�k?��Z��SX
���νKW
��ڊָ�}O��[���.Q��w_�9x�,V���<��P#Uލ�b}-�`K�c�>�!�.i��~�/��A��t+~����h@v��{M$i��$Dm���+M�Ɇ&��hT��n��z�	������a��1�CBG��%3� ���W�n��l�˔�.�ݢ�G��LO9�`>#Sc;�=�_���S��u�&׏���	j�T�^�y����~rV2=҃�j��T�����y�	p�>RE����� �\s���BWW�LG�Y�m7���5�f��V���C���x���k���y)��m�S���}����N\\�6s|L���J����U��ק������;�)W��N�׎,T9JOc��� �PBl��q��]��+�aFG/�����g��M��������s@�ϴ�҇�ap��؎0���//�3��*i%�7]�(}�o��d]��rF��2�W�[�c��<�tv�Θ6tK`)��D�������ħ��ȑQ��C�~�ܥ0(7�t����F���)� p��>\��\�L�%�!�x���&�Y���JbV��(�3��v\.v��L�ه�TP}Š���3z(FF☁�H:��vk��jU���i1�E�[���5��!�h� ���!��l+ǾK
ج�خ�� SBA{����c8�&�u��T��]�fM;��W�� @�0��P33����~�ڌ|4s�i��G9�p�?�����]Nh��~7����C����G�4d]ͅx����G��=��?N�l2 Ħue��Gy�l�O~i�iF�H/[�I���)>��/�,�~�h�ʊ�ϭS��-T��%�3�Њ�TW'�&��J�Ҩ�8�9~�=�w��.G�Δߋ���*��N�_FG>z��.h��\Z�N�j8�B�S���Y����P��!�L�-�Xr�'����/�l^!��3ô�~2��TX]�)�	�0.	~, ����e��F���8I�Ǵ���e�g��j��M!pZ�lZ��[�<���ڎ
mҞ`-!�����RnPŅ��c��{k�|��!ͦSo*���9rNM���IZ���X?Cp���������:����Q����y`گ�m�)�5U|@�.�(@͑N���H8�
��y�P1��ߒm ���13��z�up�Թƕ9���a��)��G��Z&��\놐�S��9�|uXL�$*̀�ўWN��c�м��)��Nu �j`袧^�����p�B����7�� ��� ^�o���y�'��a~�����ĥ��lE-0�C�td�!�'���lEC$.����?��Y������9�����z���_<B�-^��d|�A��_��U�/�����X[���ݺ��l]�jA�N�� �(��KIcO������d�KC��B,Y��1�H��Ŝ)�5�d��Ij�g�-^hm���}��Ӛ^&���X���u����<��"&���I���>�NI��uS��'�G��uɡ&����~�'ez'��dQL������5N�.j��c-����'T]��V���&PZ�1a嶺FD����8�SX�T�h����[:^����f1�(}S�Ħ�_��8�h�$Gxpix��ޑ(�ǲ���Ʌ�FE /4 8�q#u���]�4Ϧ��Y?~��.�]I�*�0c���|�NX�p�	 ���%�89yݭ(���ɹ#K'��϶8��D��?�j�ۭzj{(�9�%	O5m�^�e�*+,M0%}���̗��ϕ�kY+s�5�z̭lxԚ�k�FT���l�}�o����0����Y��2J����$*L�\Fנ^��)��ؼ@gGC@�{Q��{uZ�_FdMo��<�I�b��9�X%��
g��R���G3������-����}�b
6)�։$91�S��=g�W�FO(�H����
c3�.)O��q�XACZML�H( ���I��R���*>��A�
�5��]��N�^'$�$����q�sts�?�@4�)1H3O��iHO��������4��l]���W.q���[����%���cs�:��5.9N� \O���+cv���5�aAKj��$��4��<���$E
>wƹ�T��җDT;���i��� ��z�l��|A�ތ��m,��w���Ѝ�S3�m�&��}�/�i��I3Q��m�ޔa�D���~ z�HM�m�f���E���S��a��Ws�tٸ�Z�>�Z�Fs]�����'�����0A{�7�����>����%�\Y���<�q'c}B�叄��:��K�7jr�Rc�<�4��VJ���Tٰ�X�-�T�&q��fQ�5����sE��z�u���^�P~�"G(:IG�n_MD���fn��ʊ�����)|y^^5+�E}���򤄒�9&�rd�2g�Ԡ�O�>G
�	��DWL��Me���8\�����jؾl*Lě�z�t���ǡkCg�}�b�W*����=-G�ƜLPT��g6Z�Y0�_.�\:�@���Ә��4<��6���N��B�Vњ>�"__���<��G��vk����GyHm�{��}�l�=1���1-���0�Ђ�9}E�d&��M�a����G9�gޘ���f�fQ͊~�1v�N/����֪�f^L���U�! �)IA��ب�q��[��Ů|��h�ܶ��E�J\
��"� 0_�i��(C{�e�[�Sp��#�9M�B��}3"�_Ă�{Zdj1F>3q#N�V����-��[gw4T���a�<|Y{{�Д�S��*X��PX��f����#�{��8�V@:������8��I�v~�S�9#��qy�+���,���r���"�����zM�֫�i$��	P��U�t0sG��E��F�o?�QӘZqm��X�/J�C���)턶$OX�5�
��'QoJ�Oq-��=��J9tܺ$&���(6�X�1��Fٿh�fG1�������:��?��"�,a�8w1�'M)��Eo�[)�l�IǿeL��r!ݐ��Ya'3�����W{rLrAHd�����)�֗��u� si�]!�>٠�st�O�[j�>k�2�<��ӊXL�q�t�^� t YU%��)�~G?�UE����z'1i�M���&<�_����� �Yt���]L�o��%��C��d�3[�
��*��g��.O����`$��=>��D96	1�|*�O��Ŏ%1��?1��B�4�������A�@�H Ԧ{z��(�� �mn[-��ڦc�xt�z�D{ؾݡV���E�-`}I�{m=�KQ��a�=*��S�'#�z�A�[�P>�8��@I} 9������)�(�Kuv�g!�6���x����������:�P�ɉOV{�A��)�Lb�@����M!��Zv�.[�zol�q�"���p��_�/����d{.W��E;�'����on�.�PI��㧦���v����^P^��H"��+���H�s?5���W��Wq:=��T}�f4�#V�؃�U�߭W�U2�\VkIK���mmZlj#xةB������s��܂��]�|��7��T���׵����XX���{��X�v���|�2�O8E���ar�扻<�X�uJ@[�? :2>�V
��VF����#�#f��n��?0��Fr��k��/V��{&�Pv�����1�J��r�.X<�F�؎���}�ɨ0N��*f_� /B�(��Q��L�o����씏�ќ���sg��x&4��3<-~��ڰ���3�wU���mA�d���ڂ����G����Hґ
�~�ߎ[�&Hct�FD�V�w.����~�̟n}=��S?m�����g��ͤs�9c��Ag����j�XX���1���(Y
���D��$��tT�f���^(O~-��%K�#R�2�4?�' ��M	�PT����f<i��>�t;�J���ϐ���$�CK���4�F�D\C�]�Vc�g�U���[�Z*�����������V���:�د��)����-�C��芥���Zb
(��Wt�#?�!��cG�?��5��h�b�/�v$ �99��;x�>���V<�';Ei��Ȯ޸v��&�V�EQ=�WN���5��tAҊ�+($T�D�ne�p=:���S�^��F���H���-�o;�u���ZL&�r�������l.e<,�;(_�<w��+�=�[��_�	"�O�φ�0lIG��:H�|���=UkHs�����I���=97ͤw��ɾ=���Av�b���;;>��'e	'�y0đ���3'h��
���m���=1?5�l�8�D�]o9лJZ\��}D9N���	pm�4��1���=��(�e��������H� > �-��Eu崰oC�@4��ÇF!��AW��n??!ɀ��'��ہ���+�S��
A���I�.�>��q����@5�\r�/�h��)�JN�.8Ω|Pg3���8�X����0F'�K�Eg8�̜�	�L�t���ax�G�X�%����<2��+2�Ҫ���0��% /�>m@̉M��*���.���҆~�!��_��rl��V�Dç�Ŗ�ů����D㘪�ӑ3������tو���`rA[�N�a��CE_1=�_s�Ş���栝��J�'B���sN"��ݖ"��5��5r�F�Y��q-���HJ��.gB��r�KU���f�~� L��i��0��Г��/|m��x����}�1<�@�.�i�:Xu��u`����#�!6�B�N�2�����S�w��7?IT�w�j7�#�.�����iu|���R+�M��r��\5f�p��eU�$J�����*3�]W/ŝ�;�_kY�`��������]�S�[m�N����X"��*���EA�o�y`�����19ߗ��1��YR+���3�0�� K/9�QzO<�\�b!aJ�u���s`_�DvhR��㘖�A"y�y�2� P	�L[�%^0J���7L#�}��T��!ҩz��U�]YԲa��2�&��3
\{��ր��ȯ����")�M��o�E���p���K�AC��C a�}�T*�*<IѽE�HbN/Rv���o�|�kc,�u�<���|����2����/�U��:23���e_'+6��1kw&�d����;d.+ꗵ`�M�T�?�^w���	�O`�ګ|�<�QAG�s|��2ʾQ��݇vB�6}�A��ε�x����!�/m�G���oj����b����5�sW�3w��&�Q���/��q[��"zK�tG��"M����NCF��n�{h�V�CA}v{�<܊���,�� (��Zxt3@/��U�o��� %Կ�K� ���d��PG�����DG��k��3f��t�j��_�u�R�+V����1�Ї��J��E�]

l��rB�i"�Ĩ�B�������u����){��b�[�D
y��.�8e �.�r�P〧!��ޤK��<�!�7� 褊��:�<�]�>-�@m�n��9�#��0�p�����,Yao- �A�y��uGD>x�jR��0���cߝrS�0�F�N���d+ĨCE	&�u~2}��J�ͻ������  "]5Si�j��2Q|Ǧ��o_�f
�;��?�=�!1�@��R�\E��N;r�̋\r�O���#wE��jz��
�ա�C��N�t��֖G�d��z�1^s�h�]��cْնd�Fg�p�g�x�g��Q���ac�u;B���U�)���|�*jwZ�����ǌ�B��R�6l�b�h�gsiCMY�[�-�N�r#��f �d�ܰu�q´ߛ ���I���t@=3�p�j?ݵ��X�mi�P�V����4dڷ&�2��"��/��r_>&s{��d�乙�< �d�~Ϩn}5S���2��t�t�D}m���
X���<i<��n/���^����Y�/���4_�DF����b�T�^<w�����:�yyբ�<欗��f�7[3���X���]��A�7ȥ��!�5���ׯǟ�gj���5��n6Ʈ��;d��{q�e�#k\�(��26�fHr�(I��f�t?Fl��0�kV�	=.!Fz��kh�E���)j�k��?�������#8q���o75W��:�ω��,��\']'à��T���Z�j��/ŝÑwEs��u�g�����t�L`��y>�m����h;e]Էk������b�����T\��VE���ABkMe ��+�Ю��mg��xc&$F�6�ʎo�o3(�B�)��Zq�S}�7�l �>[�@�WlH/4��#s\��p�����T�*k��� |}�J\)��M��I�P��;B���E-}<�d�;8Gw�<���gY��3 �3K��A�.�2�9�v�c%�]�k�a�ˎ��#f�H\��j����`
tr鐕k��X��ml�z�q�`�񇰛���1��g�I�B�d���[
0�Z@�;��:*�waH��ŝ�T�66Oaj9�[e��6 ?Lq�
�u 0��c;x~e$�\���
y�)�R����ƞ�z�"U�C��5���?4v�m='��b�`���wZ��Ȕ�������V̚�8�|8��4�j6�Q��Dwk�&����bO���,wI1�d�5%wn�k�~�:Û0�/�^�t*P���8��r>;�Z�����}qI��L�G�-N8�,V�G���N �)�)RM�DI��풋o�w"'WS硡��?�"x�\����:m��~M����3IvY���e��#	�T�7	�c�u�QOT�|Ԩ�lϝ����l��$���ƽ�F�=�q��`I�_@�T��$�����f+����),��o�L�����/�"�x��_�*��<�:,�������eY�9S녜պ��s�G7j)�ESY��0[zh~��4%x޼�j!��~���?%YZ_6���ʨ\L:E8�d�#V�����+u�Ϭ��8//�*5�e�
b��<��J�E~Y�/)�������6�ǔ�E���Sb����o/�p(R%�e���.q�t�s�_����8Q-zu̛�J�Q�,d��xAO�P�r��w�a�)�M�H˭�C��������'�&w��'�+b!c:{4��m���I��_;�ne�r#��~��'�S�4����Ǿޡ�b��p�nl]���!#|�SPmЯ{i�  �8�J��ې�O��z�W�P��Qr@sHv��o�z���H�@�p腫�;���V���6�&�`i�N{��!߀��QcJ>r�>,
��_���-?;�v��w�Wk�Eң`��$�"�~[�$���]���J��o��3�u��qǩ�۬�}&��2k�z��c��~mצ��o���ꇳy��+�q��N�Lϭ�Gsw	ky�X����:��͢U�*RB��Y�U�J����G8uUS���ji��~pp[�y�Yt�El3��m��#}��~�#J�8�����o�b<������d^T�c��=�ȼ���C	���l����R��L}��,�4ҋ�����Xh�;�K���r� 5+�7S�YHKyx���ӅR����W��x�c�g �K�h#�Z� @��D:�G��hW���s:��T�释�ʚ���Ԯ�$�{�
ق"��T��z