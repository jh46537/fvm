��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����x�7��� ��{���[�l�
=NQ֤�G�,�*]%�|'!al�p!/�J U��Z]H]��ՊeB|Ɣ�u� |�ׁt�၏-_��n�ȩV��(B�]8�:���ee��"�Z�p�A٧[t�fD;�� �@d�+uu�&rf��H�}�߽��O�����"3���<u�5պb����������1��Ƞ����V�3|�Gi4J�VEw��Q¥��:����\j�$h����=��ʾ�,\�o�`9�\��ܲ�,��^{,&ӻ��&S��pcD*@�r"�q\�� ��'��~^e"5Q�J��e��U��[gJg��[{K��VF4�@������}���s��ոƪه��xb��st����Ʌ�1w4�vLL8L����Ϟh}"���.��?��m��r�2�xج)A���VA�{�n�1d���sKoR�_��Բ�Eg=h��@�+ig����f��=+K���t��;QFZ��^����J��+~�|�5r'�E��C�h�|���;�fvrxV2ш��xPN&l�~�8[��ŕ�a���E%z`"{Cb�޲*bb�_9P����l���y��&�AX�`e�8,LRp����hQ5���JIE�hݶ�B����մj��O�}O}۬Fr��9�f=�|����w��Ձ���yI�Ҕo'4�� ��%^d�굆����	�@�Y�t��``������{��~����I�;L����ȡ)�P};\�혏) <��2�:���;R����Pu	c�Z�� ^���2����%+�Dc�`7e����hߍǯ���y��׿��fOȖ��s���6>պ��ِ�ӣ�V��'M]n��(+ݱ��I�]H��:sǍ1~�ƣ�i�y��v���8H�p�Ry�7��R<��:)<q&��A�!7<`��2��F�4_2���qLH�E�U(E���t%5sDq�O/�W� ^�����y�@�N����lnF�9��+�
~6��O�%o���� ��@�`-j�x� X��FH�r�fWXgӏ�GUB�sK�ONw/��HĔ�ԥ�h�ϯ�P���3���J��?�Dd!���ۈ���7����ax\�q΂�Fݴ���z4s�3d5����5�rESY��;WdK
��&(�,L�J�˞W�S �h�. �YW"�=`�z%n��r �ֺ "����L� e~ QPlwXur�iX+�}�e�a��������ح�iG��^s�%O8S��t�2���a���)���Y�ֈr}���*F�;"F��L�@�����xK��Po�k*��_�GEC�QO>[�SJHƿ��`)��LJ���p�l�5�u���y�d"D4]���)�5)���
Y<�cg/�ri�\Z�;�j�A�r��'��+�8��A
���A�Fאd������Jj���9��O�ˀک�Z�FߝL��+�R�Ƹ�r9���V�^8w]���K�A�G0�=�F�j���Ŵ���dE|s�"�рS�{k|�ޛ+��䞮b�S�H}X��ӻ-�q�6F���;� bA�2�8V�:хse�CץPGn6r�s�2	!o"���d��'r��j����D��5�~��زg�+-�j��4��������b΂�w�q����2c��{c��&���1GD��z�#�1���%Օ�e�#�&X�Cvz=!�ij
Mheѩ}�:q��Fᖡ'҄K�V9�X�O���N�{V	:.:�$Sd�2�3�i�z�ʴ�,�o8�5),�1��B\���RC�v�I�>QmeL���<]�'�w�5q�*�d���F}�YN<Ӧ`!lxiNL�d�v�Ew/��^ć��Or��7[8F��e+�ր(���{�4��?*��}~X�a�B��G'�W���7�\�X��!�9h������� W��\��o5,�A9�9�CiM�ԙ�|����L6 ,bg9�p�z�nd����H��`1y�`������Zw{F$�n����'�?ڻ�_�`�|�ۇ�Y�p���4�b�4uU�a�lˉx���'lXu�R3���u�-م�sᶩ���v��<�2�'���  �zسƢ���4e \�t�\���lAc|����ħ�0��:De)<�aCʶ4�%WnO]Y�;���k"Lt��C'�E���\�׷h�L�p��9��ѐ���J�����#� ���w�4�ϔ �&~���{o�b
�oa��$1���t�D`�hӠ��!o����������)�2�q���2o*�V���Q2�:Pш9ox�P��ć�L��`�o/r��z/0v�pPMY�,z5bk���B��f�&=�r0��s�Å��W��-]
��S/O)l5J�o*C����ȒAFC�7�Yq�h������ֆó�/g�T��� D��J{���VN���}x9H�: +c�Q�~�y?c$�t�L�lh4Rt��r�\�x�5j�:G���M�S�1�ي�{�F�4�'>�εq7Џ�,P��kU֮�
8�Q&EӜk�����-�=�0)��EN��y���V+|T���G���2c�$m�w���%�Q�@��JW>W��E	�Kͤ�3�Z������E�0H>Z�#6ݫ�z��2P��On���Г�u�
t�XY�\�wg�ųJe#��3�o�>��{�b���"ƈQ�m�@��T�)������'m��ˁs�w�&B}��#����a��S3��+}p�y?k��h3��e�TQ���Y���d��?����2�(���,~*Y��wC.��}~ _�׫	��C�W6���g����g����i%�c����폹�=ڒK�N��/��$vI�th�sn`��
4�Ȝ�4BY"�^�U������ ��xj"���T�~�N
"e]��R��i{�~�-�j}_�	9�<�� �ah{��eή]��]��/�f�DN~nX>1wf����K��r(hV_qB]�����~��Kvo�[g��p�@�%��čW�1ʵ%5f�p,�[KM{	�����.�lŔ�}il�jl��JM��JG{�kf�'���E�g^���]����{�w\�97b�Gw��sޏ7�A����Af1������3N_�8�x.�z�s��?�����U�Q'":��JW���":|�J'���y�%�Kn��7����@���[|�q�.8�o>
zR��聫�M^Iz5��ʤB����3r�� �����e�c���x�|$��n��3��au1E��lך²]r(�_!�m�1y<(�Ȯe�<Z~z>%A�(�mw�`
�RA^��rے:�8T���=aP�Fm �ЮTނ��fKˉc~Js18~pМ�{�c�=w�¤c��6#�L�T��y]�v�RT;��07�!o$�OdB����d��ݳ�mK��r��L������5�:�#3�#m�c`�?g>Y�����K���H��m��t���U��c&�ZX�5as�����r(���@
���bF曓!o� 
��\Y��ij#� H�p��Pwu�/
�NN�<�R(= {e�Ȇ9�6m�5z�`!�t��ų�5�����h�iQ���6��m�B��<���i��%���xq*.�"1�Ze�%�ӫy�N�=��1dw�B0�٣URm&�E� �Vn�z����Q�j������u�F�����[�s���mo�W
�8p�����Ѣ�\-�����,�O�J��N:0p~|������O�_�t	���$�_����;l�9��Ӵ���?��e��4�6���_[W���ј�3��=�7���Ѭ�j��6k��~���@A~�ً�>�V!��Ph�5@�;�Dh*/�ϝ��{�q.���;O�^�#������G�R2����U5Uo���H��@����ex��e�x����,"8R�:J�%4���
����40a�ˢ���Ry��({�X�� c�ru�OC��9��wc�,�?��3X��O����q���]�K������wQ��l��_�L��@�F�e�5 q�~�|X�1�&���լ�
�{y^ n{�W��1FNف���� 	y����ػOF���\�"HrfA���������Q�!�I8�O.d}��H�ht�#'2\�hza����i��u��y�sMz��Z�8�u���D���66�#�V�{�8�]	1��M�FT3.��S��6�w�OcԘ	K/�蚮���{���9�Mz�r�#��B�?�>	�H��\�ifRJL�#�)5�=�3 "i!����K�x�<;�z*����X�.���&�*�˫�R��&G�I�z�^�Zk���MPHP�4��ݩ�#f�]ē�Fq�����!cnTz~ze�C��n��x���Vd��ι���-����9>_'������n���\�I�%��c}����Ԑ�^8~��T̆����w�?�:�t�0�E�?�xo��d�B�����H��i�E���v6��z��4�2&���\���R����Z5Fl�L�.�	�/w�t'?Q�Z�S}i.��g�	�]	��%�4{˖�p��w2������ۻ���VP�����ο�ڂop�$�Ҿ���JP��Kx��Y���[;�9�a�NȒ~�&k�}�lT�R��ӿ��p��'X��b�����)Cdy��	�^LQD�S��!�]ݶ�!X}�z�������
]��c�d�eo����K�Uѫ�+��?��$2�
���U%�󐝡�b�˯dm,UO�K\��mi `'J���{�a'uw$�3���E�C{��/��R�OƓg�B#� Pr}T��$�J���wLNA,�'q���"��s8��XTq��4._H<h���E�z�^az��L���9�̄NQt��o�����^rN#K��
������E~�~�?/�D������"�/ۚR7��d� �3ZFOg�w�i�MH����J1M�$���]���ĵ�,M��-��lD/dV f�le~��	f:}��=e���<]uȁ�H�ث"H������n��N>=$x�I�? {��^}$�$T��aٍ��gn0�cM�����[�E��' �Y��=!R?�a��j�DZ&��X�/�XH�.�>�\��XR�V�}FpUe���Մ���웻s��y�R��P�
�(S����a0(_s꾁��QD�
�L(�¨��G~Vef�}���,������ɹ��tQf��0��!b�ꮛ�{p=s%R�AKAO�xf��TE�*i�w .�/����z���o�y�!����8�K~��������#��1����-,�x޶L��uPú"�l�?ΤB!�a�.�t��/ǘ�B����5<D{�)�&�}���V�@��~����D�!|D,��[��0�T���ݯ����Ɗں��"�߽�ޜ|]Xݝ�Q����T��J���.7�>�[]�����M%�|��QG��k4=�������5�O���xoWd_�?x&���k���0��(�L��o��i��\��Z�Vu���3�@@��L���O�
�<�!�<��/��a2	@@b���Ӎ
���$�i���T��\��&P�2�P����;e�ʚ�	�J��;\6�o��p���lw̽��g+W��Q��� �v3��cr�p��J)m���sA�̽�N<w����o��@^�wnN˶y��Ǯ���U�a� v���-�O,��a2ۋf����t���j����=��|<�/DZ}V�J����hlш��Ր���]B��x�U^A�a-�9w�K��eا�o�`Uǿ��"��; ��ud������b��jO�g�;E
Jԓ��!�>�N�����V+��2VA���M֟�)Ye�����>ֆ�$�5T�A�Q�+:�e8���G����5j�4��.}V����g�W<�ey�ch%D��'S�I�!����7�V�R��
\�!�B\�?���5�0VC�Ay���@P�2�����rS�b��!�-�ip~l�(�(1/����Iy.��7تwg��+i���c��a藒�a�I�.u͗��%��@:;B'Mv����ˏW��0�b�W��5f���	E�G�Xe�dN��A~��hpE�������5.t�H�N�г`5ꥀ��\�`���5�����0ߌR!��.nd�cY��U����U�:Jd��o@<[��DB��W��>�OЯzx�tC f0J��tt'Rb��C%̐P?��"p�����~� �\t�&�rƳg���A�����u����=h�[&�ֆ�ja`i��xg��]�+RX���q�ܭ�N)@��؂�f|21��5�V�eAQ��Ch,���E��/Z��T� 	"��f��$r 	v�ѭp,����j��_[���'�NɵZ�MK�lC�^]�JhjѦ�W�a\��5�l��Hў��+��x���vJ�A�0j.^�_3�Y;�.�!���X艛g"v;������W�u��
G9�v\������Z���B)��1L�滺�8/N��vZ�5rhy�kN����O�#(+�q�1/���l]�z�\�