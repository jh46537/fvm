��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S�VJ���ɾ GK�rA�!��}�x�E}ݨk�fի�u�(���L K߲w�.L}x1F2�#5H�:�'))�6_��\j�S��W��w�.㆔�[NQ�6��iM�@��9��eh��L�@�Fb�%FZ�"e��R���W��@�s3a�����膂Y�:�D���!G��j	�E����}��Ui����kh稯ka�"������e�^��6�ɠ�Ij��-���jW}e�@,��=��\�`�Ǩ��:>_2�)����������t*�� *��%/��X_0�2�KwS9�ڪaԟ�	�踷Q����Z�@Z|�歊�)���ܰ�K���"F�"�;�ŰS�d&>�،4j�o�9���xD��h[JH)���m�tS����\�ɑ� �n�{ƒ;PM�����>"s��R��m(ɠԉؔ�W��6���ߜ=�5�%�_��+*�o/�Wv/�nW�S������50�u#�����=�O�3b�w��Z,L+F=5�'�?y{��yN�2���D2�m� �p)*�CW��F�7�Ye�ȼW�xs	p���-0Gnނ���Q��	��q՜o
����D+�g��!!|VeG*�s�1� y��!��FXV/ao�
Z�#o �xE5�_�=��جƒ�K����#������\?xi`i(d����#���&S����$��a%�o5�H��}\�����?�ՒI�W��+|Vz/:�2�T�K���f?�k��A9���d�̺}���6���K�����T�ʫ�n?�塲������*}�Y�9�{��S���c�{ҩ����H���qn����qh��W�"�&sL'4Z����B��,8��w��BFd�8M�Y�b�oe�Wl� }�$�ՇD�O����r,���1�υ�\\v��<Ɗ��h�L]@�'�Z{�e5��w~��t�qJsP�X�q)��"ˀ�-׍����������@�(� ��bx������O�3�Ӓ[O[	�Q�����c���x������_��˸)��+��hNۚ�-�4�G�[��T ����r�͸���6�GY����G��E<Cn'C@>^=0�DFj_�hEň�
����6Yv��ݚ�n��r�'U�d/"�OS����<�N[�-��������O�oH�Xd�K�qF����mʞ淛�vKBDݽ��F*m��W0��iH*�SM�-s��a�fո�5/?�ز�yw����Ʊ�^3�T�%��ޮ�~�N'kK�u��M;�&8&������0a��B��{B�t����@ֺ?n~`š݀۱�
���
��ާ���2o��E1��*?�X ��1֐��g�0� Z�(ӖrA6��r|�5���"M��� �zrU�Y����A��-���Ӂ�Q����Z/*rl8g���1tFC�c���$	�����K�?������5w�"����xG��i�&�k}�k�*|}Ӣ�#K̉|u�_&�o@&.�
�\��w���ߌ��L�S[ {��3J��2���F�م��%���}~t�:���]�;�q.~��j�+i��L�_|D�s���Qa�!�_l����=->݅�����()�L��̾��94�ċ�2C4�N%�*J��&�+N�,'/0�^,a��]S����;�A�H�Ȍ�6ua�=����F��%T\�4���K�I�2Ӡ��R�D�-nt^4�P��y���ڹ,]�j� <;�f�I���\JY�Y�����Hu���RK�C��p�2k�a�M�Ǭ�uR c�H��(1����" >��[:�
�⬿�(���r<3Ku��K���{�/�6���w �z��݆�����-�u� R��o1O�[~�����?�b��)�9��L�	l�vh�/��?�g]be�*N���)N�W�ZK��x�)`�*R����6@ID`����vFګ7��*�^�ck��/�عx��Q�
>�]I}�b�&D%YD�E=�-������m�c"+�d�'i�,R[��a�p�O�2	6��c���~CÈd�BRAڬk���t]VKĕ[�ρ~o��������1��>�t����c��x�X,�F �h��������ő�s�֓ 
N/�m�y�VC�����B�������e��ѱ�nBx�P˿����H)�������p��W�Ϳw��"���4�Z���?��m���
Z�a�&5�=���Ԩw9�����j�����5mM�׻-�z��EN�C{>�@/�Gd�:%xə:�9,���̀C6t� K�Iγ�.�����d�LX]9B8T�R�����l�^��V�ӆ�i��4��g�s?AtH;?�Lw-U�yg���ủ��k�0� �"����<���o�dƗ�pBg��#��r�a(��ho���V,�b3�u@2dk��'<�t���GcV0�]��,��-�=�Pػ?��j%�V��� B��$�H���(=8���f�;GT�FM��ʨ}I�-�PaV��x�I�)�c}ǐ��_�.qc�"~���+`�)��
�5y��*Ω'P?�O�����^+�����/t���F��u��G�B�3���b��O�!�*=k��:�Q:A�2�{��ԝ�Dc��J5A}��&�w�$,H"h�"m�cNUs�t� =�u���6����qOE�UƑz}P�pD�WF~J�L&̕��(3�vU~�
nQI� `��fsA�
s�����W��\�7;�p`a������8?�K���(���Ӡ�E��0�XP��!ZpЕ1E���
2J����Kٳ(a�oC0��A�<vi�pLԒ�0��,�B��&@c�ЦTˀ������S��0�Ʋ��k��2\#���*ۧ����}.�Jj"H,y��9N�on���JQ��ɉ����i�D�`�މ��N"��	��5b�A��.?G�q���J5�:[1 \E��r)��v~쨨�����l�F()�K�_�R�=�s�aM?(������J���5X�5맿;s�k��?I����)\C�u`XMA8��TC�X�Ҝ�nioٲ�ڒ�. 7w+g��^�,�����c6?�a�0��]�R�ϝ�ў�a~K&��4���ͯ#�0�i�{S��f�}	�D���^0tr���oE��
W{����15Xt�DB��xe�g���kJ��Q�N\�4n��몦��	k$�41/^<�!1YdKƍ��б�+5�{ ������C�\GO|b!{}��BN�N;$΂��_$�Z�� 򂕪kH��.��R����ըu���L���g���4e!f&d3�Et�-�����8!�յ!��d-7D6sac�~]�?A
g���)\��I�쵍3us'4��ڀ�����
s����~��X�Tฦ�H��:����Κs3Gr��/`��ʞv��=�V�p沅֛e]@��^�f�:Y�6���-�cQ
0wG��p -#�(n^I�QI��N�e�^#
��{�ڳ�?X	��f%Y����t.��P��ޖ�\�yQ?�@�0U�[G"o�Κ�����)%}e-�y93�8."��|�)fQ�<�ݬ[HF�ak�Go��!���D���g�3�� �RѾ"��r�s_-|H���	����)�`r��(Y�vI:^M�����j�Ҭ`)E��W�5�m#y��V�_a�`�ݓ�F;nn�-{�����U@=Т�)glG��Gp�e��f����Ł,T��D���'��|��*���hlk�#$+Ζq/IS~R9��v�0�Z��&n�߮��7�!���EE��JҪ^���Z,zd�B����
�;5�,D��0�/uk�6�T�0&K���0�P�v�>	I!V��L�b@۟����M4Y�+�P��w|���_��IUW���"���"��/��=ߤ�� �"������r�1�7����\L�����k��Sקj�K�� x�'}����k�'�k"��$�n ��ct��$����	р�u<Uj�OZ���~�Vr1K�� 2t�J�(��*��D�p�'�#{i���dU��4ѓ:Ԅ�$���j�
>�}���;+/.Px�2���3�Dv��!� ��-���'���͌���� S����ꛮ��@ K8j���{|�*i�)�q=�<��γ#��Q1�.�εXEI%��<f�"��2����Ǟc�" �A�UF�4z�����#	S�ʝ��k%خ���c���m�O^q�j� K��{45��f|��矪.���M��9��p��t���J������0c��$�\�dq���u,�W~�+n�m�ӕ(�װ��P�D/�U�M_�ja���w�<&�?sѓ�����_WkgZZ�s
Q��g��T�p�{��ړ>tL�"TFct((�1j���P0�W����!g�� єϞ�ׇ���`jv���w�}>7��+.fP���~J$��p�aWǡ���E����*K�$�����f1�WrB/Fn��a��Ѹ䓴�pMkyAzS�˨c�$m�6�^VP�D>	 �(�L�0�y��&,!���^�.����* �K���MU�x��	]SW�]o�����ã������zP��*f;kgHx2�������п6~� �j8?
q�VIE];W1߀��R��H��U5x����������S��F�>i%	����Ћ��� �> �>e~ӚfH&���v���a���{��U:�2,�QPfY����_�m��h/���F%�c�3h�/����� ��Hz�I���_���i���d�M*��`H����D�wу�T��sq�v�YwWnm+e�}�A�?((�mZ�v݂HYVi}ܹ��,$�U�mU��h��I�&��t!�ڒL�eE���a7&�nƄ��{�w����(填�!� �0�Q��ǔ��{ʃ�xol�������Q�_<���C��,��:�(|.��,h���n�P(�!V�:-����bs�!}�%=�p�[��B�:��A}�̰gL������Q:>�L5lR|`��0�OR�[:����#n�Ŗ�@�m�1�p�X���6x�Y��&��Pj���k'r[��be�fi� �R���������`<��Z�w��^s�ݾ&��K*��_p�#I����,���1{��fO�<8��5�׬v�
�[c�u;�N��B��\��w��Ot�E�O�"x&(�$m��iY�/�T�Ԁ��+����q�	��G�y5?_S� ���{1L
�sKￏ�o��*r\��7�L������|� W��\�Jy3~��G��$Q�l� �^_Ҵ���yI6	�X�`���sŊ�uϼJ�c�h���"��n���3�{�w ��:J[T���w?�|Hrf1�k�G�)X0/�s�󻉺X	�A�	v�&�!$n0P�g�_�o����Rz\���H��k)� ��)�o&B��7Ԗ�nUQ�.�Ȁ�h�L�v���\|?�n%�p��`��o�@$�mK^
�v���I�o@����1��	�������|z���iS*�ݾ{1;i��/eO�Y�bsm�s��I%6`�3w�v#<:ҡ�4����ѧ�L����u9 B�-�T��W�0��y��K���԰?s���z�n�!��躲 V]�;E��n�v�	,�pc0�7Y�)��<�0gs���՛�dˍ��뎁��3��}�/+�6��R�'�y6���?+��q�k��h�����@'J����CV��H��;�Z��h��L�Q�gE�7��57Fx�!� b�z9��� �bg�w^����
m`�Ƕ|��/��S,_{���}�o��%w��)m6��=��z���Cm�V�pm��q��|o�U��}�A��W �jˮ-#�r����]	�:��<��;��Z*��yw��	��%sȚ�$��l:�{�<)����]Ѱ��u ��wy��E5*]�����F@�.ۤ���`�|f�ɒb�:HOM5jW���/�]A����OK׹\�E�^�Rl����?�,/���_/	���.n�'�I$d��p��%��i!���t4]q�5mtm!����>붇g=P�^j6�'e�׽��{�:^6��w��mY��a��^��p��6& n։$�Bu�)^�6x&�
EWω���,DI��9e�4�EQ����{��JW��������F\KG�>#/�2Tb��Q��rο��,j���oFq�B4�1��mf�*�uS/��Ӭ̀O�H~����[Si��~�������D�C�7!���0Za"ڐ�Bصs'��� ��X����x;��``����Q$C��ӯ�ۆ�<���P!�0��h�|�?ȗ�D���8���؉��Ф�/0!�8�+��_g0�R
�Na��Od�/�%���̣X�ȱ� y��p-tZ�v=	ׂ���J�a3����-��;��fU~y?2� A� Z�bh�c\��/�*�z�k�C�u6���u�c���⛧�R-/����#�Ul�[��bG^ihP��}q�|-b�|Ȓi5���=
m�a$nH�qj��},�]�y��ַ��XI�c�� �͉Z��ב1М���$�Ѥ��v�֍(�h��PҼwt}��UKDF��A9S��7��1��m.�g��ЩWƯ��$��]}]D�TA�K�"��=#J����0S-�,���N��׆�S�G��'���?�Z |��P. fX����CXn,D���y?c�zgu7b�6������|�]aި�|b�+���qo������?���G+n�����=��~ٛ0U��L�769p`�9�>{b(��c�壞�Bq��پH�<v0��r��W���M[I���|W^�Y>R�J#	�n&c"1zb%��:l7j{iJ;�S�D�3!�ީ�u���AZ���hiZHS��lf�C|%�o�$� ��~�G���4��Ձ^��{<������J#׼���2Z�s��Զ+���n�|��:(�cxJ��z�D�,��Mվ�E���cG	�Qx߹�~nΑO�!�skFͬ�y�ٖ?��������hc�x�v�l"A%�]z����D��ɬ��|M
�8w���,�˱8��>u��N�O� ��,"��d-$���t�L}O笔����Q��-]6�\h%����8�Go|ŷ$��KH�f�:'3"7��ݯ�R���.dI/I����,`W�NYVw�8 ����a�x��86��A��欌Do�6~�>bι���yCI���;�{�B%eʯP�C	szO�t�L�mlB�"��/�+e