��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&i�uˤw���Q5��xzJ; !p�-�ߵt�Q�וi��L��:L�p����6L��9�x|z8��� �-�� G���ݶ��/�W���ek������pc��l~kS�N3�;f��ԏu�벗��%L�L,��+���ڭx{'���W�S�.��U6��N:�'}k�AN�70A�^.{�f�·���=\Ђ��6����~۠����;8���7�ݠ�{j��	t~����r&��h�! ����i�
5BƵ`�>c?.hq�6w!~�Z���.)������G�������7�3�0�v7P�f��{���ȴ�z�ԧ��!Y=!F��������`�}cO\U3?���r���.�c�M�5r�赂�ɨ`e����g`���TdŬB�3��.U��qō裵vN�1�_C�nQ���D��$�( ��
='EyP��a�����]>�©7d�^���=K����\zq�仞{i�.��cG��h�^�D��pil3Ko�6����z*���\!띙7!#�!bJ��~�5_���ګ�w��U��G^/`�"�߾L?�X:��j�CDQk�H'ً#	�)�������#�Շsx�=~�r����
�9{���7�9����.l-{��q$?+�tw�F8vJ>r�`H|V�'�՟���V�QL\���T�H�D�P�J���)��=�.��r�X�^k��冁<��r?�F�2o�AW���RsZS������u]0��y����d�+�����5���I�j��n��P����(��!	�]�Z�����)8��{�t���a�G�c�]d��aYI��x_�F;�D��z�X��D`,��-2#XoՈ6����6q��֥=��[W����qp}[�j��+��O2�-H�'�0z; �S)�#�,7����k�&g�B�a��x��u�]��Efw=��A���>1�-��� �u��\�$g��2�5���%�{���lUB]�$���c<��=9Έ����kĲC0x��^h������������p�5h� #���N��d�L2��!��I'�_�@�7z�rD�0��`퍗)ծlx̀'/s�T~�7��P�^.g�����	��V�p�{x_��E��ٻ�?9v��yh�W�D�Q�QS���5������ry@���H�';P���)�h7�|���"WT���4G2�2�K��3��՟+�rF �iҰ�	Bj͋�m�S��1ٳ�6�X���1}|>�N�2C�h�����
�^�Epj]Os(eb�++@�e�6�>��+����΄�c�ez�
N�ނW��o��̡�@^R.y��{!��W&_���q�߫�u� ���z����@���� (U����f�)U��=�8m

Tl_2�a��l�]��/�ܪ�1b�րu�k��S5��t��n�+����6K�$�����֛�΄��vL"f+�8�KQ2f���w����\��X�w���s?yd��>^�߷z��1-z��d�y�gV|s�X�����F0�w)�>�Y�b�Ǘ�e��$ڂ_e�>�|3��E��ә�s��M��L���1��Ru夗�����?ڼE�J�/,5�[�����,����)�B?�U؋������=I��@x)��=��YJ�2�iI��k3vt��pi_��؅_g�]�x���s�]_]<2V<D2|�RDB����bt�Xς���j�k�Om#�a�O�*2LLN������\(f�H�`*��Z���k��Ia�W�/~�?!˩+��M�nzw2୹Z�Os�B�}aEzf�������|��Mb�l���G�x��5h9�ҞN�������O����i�=�>�E�T7�z���X�A��|��y�?h��������0�87ҏ��E��@���]sX<Y��|������ZʊO�]�铘Vų�]�ʮӕ$�:+���t\%�V顿r4~ �VUUb�ᔨ-�uoL"l��0ŋG��K�F�;O]ޮ��K�Nn3ڇz��7f�tXx���7J��m��(�KfN���;���:)�MG��:r�� .��gi�{:^��}��i�R��#����Ϧ�