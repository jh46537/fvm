��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&k�㩓���5�In��D���-Nx�J�G��0�Gb��_t_+�`t�ɢV�>2��y�|��0�E8/�P�5��~��@�egzG&jI�#�a-&�2J�@+�������P����ۿ:���δ��������lK�����D�;�ߜ�lS#�[�g����.�}O�)�  ��h��TVIE�ʇ�n��ES����uG�[�(��Zq>��⨨լ��`Tb1�l>����_#�S��5��D�����9ӚN����P��p� Q��s�]�6��G�k-\Ν=��#Lo�F�a
<E٫O䤤u��yh��&R*�:�G�_���@R$�m�E������ٞL���3w��d��jMWJ��ZP�ә�ʣ���'�D�x��O��2���W]������&5ңr4�-��|���,�e��Q^3��[T4�3���"�]��mUk���O �uLM'�ڬ���m�q#|��)U��WllK"_XG��ԅ��@��;�H�nQ��fym�g��v��K� �[Z�w����-�-h�x���>>�fV0i���2��.�#���F�� -bT��E3N2˸�Gk8�4��c��T�Y<!\�x�FxѰt�H�RIr��SI�0t�}����F�$�	���|a*T��~�/�rO�&q`�������z�K��r�&K��� di����:-T��v�EiT�����pD!�K�4��t���A�Z�In��'�\�u酀YD3�,~�C���,	��� �����!�wM{���bp���5
:�Q��ν�Vc-�����ʋ�[>�#�=/T�Z=��BVTh'9j��V�
��R�֠��(`{��W�d�P��.y��<\�����J�O�`]H��Kj��c�����66D�OI�<ٞ( E���0�������*Wz���fi��6�3߽����*����>ZV�&"��X���^jP_´��悦��ؽUc��M�։k�H$������'�;T/���F1�M,m��XC�k�/�J� 1������-mv^}F.�n�j�qq�̕���[���\��	�%
g!���s�+������e�	0��n����>
�Y�0�&F!ˈ].#��~W),��n��Ox�CDW捠���C�E�ؗ���9�(;��ˤ0E��x<VZ�R{{�p�p�J:�'׈sؘ*4�w�[Y�.���ϒ|���H�2�����n���W��z�s-�!�(��̏g�_������ �,��AF���#�_������
H�c�OL$qfw�2�޸m��W�o����d��0X0 ~BR�;P�"��=�����'�L�'r-mc���%3n!I���J�=i>#�2�k�Se���m�� ~����p�a���g��j{�(����qQ4�q�f�"���f��ɯ�ą�{~��m�?��l:���_*�a�aoY�\@h��p�A���*)�&��pc�{3�sa�^m2�����z��A���CG�X�X���@?Y�{�l8��6>�����d7��c���Sk#�����r�O��D�<�Ǖ�����N(�[�2 �A������&�����?u�1�I��9�О�y�T����fc��^7��:���
���_Io��:�x״ET�J�f�p~�׽&=}�r�yoڐ�9��Ìrx����c'M5vT��#������pC���u]��J�9*,�)���ʨ��q��S�R�r�Ʃu���EXk���G�1��5���Wvs���L�>���C��6h|�Ʃ���rC�N�p��"c�1Rj��9/0��e<p�Z��򬥶B���
�V����Y�\�L- ��{m��".V�<��G�,=t��C~ws-�C�2��� m*�j)u�o`��{�Vj�&x��[��.��FFnl9��� g��D�#l`t�����}[{�*�����[���,(�$�'_���[cgߵ�p�7�8cО&NpaF�=�[�`^����p��(_� (	�`e��by��p�znw���Qᡥ��o��?���uƔk��a&��$n�O��p�̂mv1����#���\#�p��|=�L��VBesn�J:.ȥ����� �hq�}���r)P�s]-�1���x�ߒ���j��0mH�a�� �?�߽�����x�JB��vi�JZغF��h �6�0�8�d�Lz�ѥW�h�Ȏ2Q���l9IM�YMqz6���8뵺w\d$쾑O�s� F�z��;��"��־o����#v[�6���Z�����V�b\��D��^Y��:�ĤU�0�k��)#��[�E96�n����',Y����z�Zt����0e�8i���'h����`>��{߸��_)�gf��$a/-�#*91�������;���$�,���X�=NKv@ܫ��ap�ˢ9���sءAF F8V30|�e`
�/�%M�?_]��c:^H@�`I.�U����Ђ�mE��c��vWȝc���&�� z�n Ɠ���ʒWZ����rL����b�.�d��<&��+^K��f��*�m� C,ߗ�B�F��J?U��&�*Ñ��I�����~���_�˼^Q�
qa�A��鬻*6�CR�*��Q�P�q/(���`�SdtpF>d�<29j�G�R&=Kk����}xJa��6�=@ĸ0�D���������<`Z�/��Az ���D<�ĥ��
����~�t�;P��c����Uæ�K�|�8g�C4�gs%��Q��̤��A�(\-�� Q֝7'rˠ�R@XC��MS������au��3�3�@��j�VSZ8�ў��L��@jf�@��(��C�o��rX���UaZ]�/6$�\��9T�V�\�"�8	8~^���B�ӣD�k�� �A�d�|�UMȟr���t��D�Ƚ������M��8��#+�Э#V9���V] �;cm��UnI[�@5�~�r.�q6ǃ#g0*/V�8H �o��MAr��6|����n����g����BD��*&/F��Sg&=�5e������of��XpN�vk]�1:�'���4���ۯbͪPƧ�Ra�0���u�~�Ȫo�XGf�����t�Y�(X9���Dw��W4[��۱�W���a�kU�M�񔍜]iD�ܵ|Lmf�hiu-�x�]F�n;�[��#�b5��^Ce��Ե!?E?Q��iY�A�i���X�q�utń�A?���*��Pm�Kj��т؏Ø�dJ>o׮)��`���_����2�nx*E���k���_���.�������}��h�(�aCk��e��h���K�Y����E�����\��u��[�g�6&_E���X�F!Yz�h���,*nզ�5���b�� P���/�!>l���[Ԗ�j�A&��h@� �@)C%O&h�iΝ�$e�{&�kU���ն�a�G1v��v��H�D�%g�"�n*�;�Q5�$��X{�<���=9��<�MQ�p0S]���
������+�`�&B����M�5I���h���{��$	v?ba�a��ʶ]�zq�5lй�X�rg�)+U��":��#��%!	���4ݒ�(�O��qoq��Mmaj"��������8�|U�t�C�t���6 �a������%3�(���x�9���I����}:����)�%S�%`��?[�m͸mTg�l&��?�(���gO��ne�,'�J}.��!���H�T���}������x�$��j��K!P=�m^�>�QQQ=܂��\Bc���zw�4��g�k�I��@��b�}1dC�R���h����4K��iD�3H�p��q��{�ɑ��2M�?��;̲���'(��v}����6u�B2�^;e.�Zp`�Ŗ��k<�\+��a1���X�M�Z�ބ;ļ
i�iw�'@�[#xƺHPn:���'+��"��޷Ω�$v̕�<�j��\S���ޯ�B7���6�OB����E",�)�>�k�dβd����.���\��t�׽�-&n4ݔ%[�&jn�#p'�O�}�	k��ګ��V�5��o����'�
�B0��2�b�͝17�3x�l�~	��Vgcn[�~����ґ��~� Љ�wfQM����!�%��a�`��?��l� ��"��>�~�Շ��$SEѫ�mf}�#��M���$�L�T���â�����&Ev�37~Z�;��ɨ���W�J_��y��d �Ox��I�~#V=��c/!x�0�3����,c�y�o� x��F[���e��_j�Ja���A���|T\͌�F4��osH����Y��s�h��.��Q�Q�ݑ�����<�b�@�&B���)xTZ# o�su4G��T=��H�i�2�e������O��} ������hD��'p���%�t=Bjڎ2�}K6!���5�*�l��8�-��<�~IZ:3Ws i�	O�9���ቇ�q��QNbȧ��fA���o�Hv�I�;q(g���0r�L�[�i�j�>=f>�Etn�'��-�P�$��=[W.��h�K=�퇀�3�������7�v���{� kQP�TPrL@qؠ(�S��A_vm`y���˟�� ֽ��ur��Eؗx�J��l��U�ɖT���͞�Y��v��̸���L�!�t�!s�,���Y|'���dB��� �
vC�h
���g��w�z��K qN,�f�?�J%=��͹�=b�(y���Q�6']��O��b|��s8�^;0���{ʗ��T@kT����k����x��5b(�o�P
&��I�R <�`5YhUj8Btd/?:�ۇ�v�]F�z�&*��J���S�F���-N�[q"G9u���	�h�y,�e��