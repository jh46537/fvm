��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&.�[ʽ��@xg[����W�%;ʉ$�ړ�(C�H����Z\��=@t�����T�YČڜ�Τ]R��7������n���f���"�N�	Q�m�� h�~��\}}�2�x���ge6�D��{u������gp�o?I�O|��<���J�+�T�\i#���q󴰅I�V��̗
��E���-��Մ��ൣ��_����Rg
9�g�I��g��.R���Z�B�FC��4^O.1�p�/QH�|�SXm��'�7��¨"�=xuG��KPHh��j�fܨ�u9�#�M0���C����t����_�w*�)~N�A܍R<^�J��#��`�`j�ݘ
x��}�n	-���:��?�h��P\�&�^�y�A����̀���S|o���Q}��v�-,����&L�a��|c
10��>(��9��s4l(������+�1if�Ta��ڹs���v/��~�zQ���͝<Pk�ec����2�(}�؅��1ү*�4H���y�)����] ���-R���ޞJ}���7;�!��qh��B�B����su��v��������!DM���V(Du�"���f�u��ִ�rt�*����s�Y��A����G�$�e��.�6֝PRIsס��G�z��K��D(yH���I�ߧ9���n��N�3���2��玡�=�"*��5��l��<Y�&�0�̧��`����|�K	㭪������vic��+�NN���.RBq�l`��2��"�Z	:���z��/���2"�/�41�+��;���[�j�7%�'����~fI�RCo{��x��s�ڻ�����1���Bt#߬�ߩ�Fp}1�C�����L`/�k� tNW'��X���Q���;'L[�������˨_�.)jڃ��]�^�Աy���lt̸-t>ñῄ�wo�\���=@��;D"�<]����{��R��[ C���A����.Ȫy?p_���U���Ů>�M}Ṛ��G�����z��0rg����p�9��Ϫs��.: ��}#�R�>W �'z�J�ᱲ������w�9[�I��~R;�8��{�o��MF�pa��t�r��Q�Nc�R�^�Mx�O�^��u&�\��]!\�[����?C��c� ��v�g2h��̂{�:�������e���~�4q�o�[�!�|�jZ��w*7���x��h�9�X��.��r�Xq�l"�� $WժOSp: S��B;�V7#\�n=����9I5DLNY��:�,ߍ�<�ԓ�쫿=�o�K�Ѝ(�0V2WA�ֻp
�qae&��*�v*���Z-JXSW[\Nuh�a �z�Mc���h��;�E�tb/Ǔ���ӸKkHW�,T���8R��Juw�0�5��G���
����2N�A�6�>����=.�0���Mn�L=�����9��.O� ~���
XtW)�1�e�S���f��eA��C	�EO&��)�A{�o�2�fQЀj�y��km����+��)5����)�rZ\E�M���E���-�8R� �ˋ�d��=����9�XXјIP����V�o*�˫�4���fP�����l��*�H��:B�\ �G �N�ɲ4�8�����j�dH�r��pw�f�0ej"{Z��@��vqZ���й�E���E����۷��I:���Gb栯��bgr,:�M�j�8�ҕ�n�ZՖ5�ɭ��8P"�պ��M"m���k��f�z�L<JA�jV<i���xu34����T�/WY��#Lc�����x�ƚ���gv���� �y�*�sW竘�[B�W�	��}�ex�_k^� 7u갴 ��/�����0�X���"�?	�F��2 ��D��J���O���]��F]6n���+*��nZ:��H*��~���Y��yG�`Y����[�r|��*��\v"���]�b�� �����.hnB5����'���RXU^� �0iT+v�H����Jn6~��l���RÊ�}�.}����4�O�k�f���Wg)��rY�Bﲕ��6X���s8cʊ��zz��c&��WP�h���5�~�G��p�^�1#G"_E��� ��f�D��3�́��g	�v�6���S梭m������΄	�G���1v7$�W�����y���(
#��?�w��&А	��s�LSRΫ��U�D�[Q��hlɿ�ue���r�8��Ă�U�c!s��m_�]S ���,��v�	�!��P����X�H�_������1�\�H����\���es��z�s7����0��p�
/��1���؇/E���Eϖ$��B�5p��֖�$�J��%"CK��M���-��)'��WI�!��ڥGܹ�k����3��v�Ҳ	�-�ӯ�ڱ�̉�`͢=�MI���|_	�|i5�� �_;S5���0r�8<�(��:��'9%���2���h����M>��Ǿ�7瑥�y��#�W�vɝ,49��{Vv4�It���Z�Ob��3��%iZ����&�2#�G�!��T[E�w]r�V�e��k����3�2�&V`k�t�((``&�r���CិP�V<d��M}ҹ�rEǫ@���=�g