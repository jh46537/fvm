��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&����H�� %�]̪'�;��U�;���,w� ��U-�
�u>��.�Xu����}��1���]$'��b�S���'5��-K:�T��0R>q�i+���֩��݋� m�2�`�B{�'��mi(��[i��,��� �J������w��4����V �z�Pf� 
ͬ�	~z��2}|s�&�٧q7}���߻�o��nŁ��`'?&hT��B#* !➝<@�YF�F-�^i��F^%+�3�t�w $yL8p�W��yU�t�}!��L�/��J��M�Va2�
������SD~�����ز,�
�֯��Hآ]ք�>1ܐ흜c�n�Gi���Y�����Qp|�����t��S"&�5��x'�h�<��DS���ᵁXW�B�3���E�'&�Cr?\�4FA1���lJu�F���ʸ\�y��>����\.��b}snf�9�)>�������!Q��x�ߢ�]��Od�
��`_z���3 ���<gX���iRؑi0��~Ќ�f���6��"ߧ�k4h����R�q�7��z��[<��������VI��׻ޏx$�(��qXuq�(1��.���<��(XޮWld"�k`Y0L9��%�G-lY��c�#�r�wǐ�����=�+IK�`�9��t�i��\���q�7>d:�>����w�z��H��)�l�xC�yߡI�.�v��8%t��9��e%L�e ��:ťGC��Z� ���^�9�?���v6��%M$�������sYq/��9�!��/4X�)/3���y��w��Ԩ9�g�w�G�u�A�\���v�A����Ŏ9�k���@a�yG�\�w)�-��7
g5�ZO'���Ԇ	�>q+]Ӱ �!�����d/u�U�>DA���jI�K
iQ~�I�ў�҉����)".5+�]�񳆩3����*�S�(��>6x��	
��"����3��<D�~-�S�÷d���4Q����J׭��@�-��ȓ�K�� ���Y�n^��.6�Z�����Y��%��7�H9��Dv�Im��S\v�-���u�S`��K�` {�>�@+W��Q$�2��o�|�E+`��
��"���t�\�I�0�hܨ��;뎲�,�E+%r���sQG��	}ȶ ��ፌ�}Cd�ds�m�� C��E�[l_���K����mE��c��-�6Ae_�����]ƙ����Do��8��ԭ1	���[>_􌴖F�DW�W~I#�a^��k�fS�I�s!��j��f=Z�w�:����j�a>B'c�h����P%��Aqi�PrK)Q�V��ٵ�i7]�s��^TC#�yM�g,�%kڅHе6��&E��1�����`�|�H'u�O��2l��D?{�B��T?fx0Ҽ���"ʢ2
�G�_�ġ����Ŝm2��]{}����b��M8�Ɨ�K7��ob(�tҎ/7|����ZR��tX��n1��t#b�\n$O\UL�Q=��
�����|���`_��s����E�X�˦V_n��%'j"���cv�\��PQ���>B"`I��N�tp���ƙV+�:�cNX����x!l=�:j����=��Ҳ�5HN ����	��?�4	q�1h�
t.k׽0����H���.��O桎��wg��Ը�r���c�(^�$o+���ī.G2\���Rsľ�[MF�HR- �yveE�6 v<S��V�ϋV�yP;xBU�O�͖Z�d�o��O�HG�С��ecO��)�>0B�dU
�~B�|��I�r�;s�&�|�\�Zvh��"�ğ�%$#f^�J�Wd��o����P�4�`C���Ë��xZ^�Rd�g��s<�㣚b�,u豵�#�,O!�￉j_ٟ+���*A�/�ť_�,5���*���$p"�&]k�3_�����'����r��tӴYy���\���D 2DӦ=i��Ԇ�mV�qv��*�@�U�b�XP3H��-�Eb��9yR"\3�=2��T���S; gvld��=�B}m�"����f�Oڻٹ����u��,��y.gsKo�!��' I/1�,��k��k��L��<�Hϴ������g��f���?������D�SJ|�����X�����(�w�l?����P��z(iq��F��V����u�Q�	J?=B\�聱ft($����r�C0`}���ȳDu]���D+	��ދ<m����؉Ч�Lv,�ZH-��m�ָ����*���%p�7�'��Ό��ֵ�&H����T�JH��C~5[-R�(��,XX�Q�+���%w���։�3�M��grQ`.���2e��Z�3�G��x����\�$����m4BC�$�UmM�.V�Z�/B\� �L6h#@��$��X�'��<�@�baN��5�S�q���oa�� ַ�� ���R��H�1b���}�%V��?~pV�� ��Uū.5@��Է�lF���z}�i��3N�+�W/s�ί9I��t��,RNwmn;��k�#��q�i�KM�Q8��@tGy�h�%��_�(�I��~吸���
�휁rE���2�q�5g9�i�OOl����ڥÜ>˖!��;��ol�ߜyg��/n����Ʊ�q��_���f��q�Gv���]��؉m�s��h� N�;]L��9��6���_YiJ��%w�+2���ħ�㚳3U,�$�����ީ�N�'���'���� ��0�{1����]�u��7ܳ<�]��d�*�)��z���ݟ?�r�C��`!�Yun��%�F�Щ��<Id�~*#�U]�=�����p�i�ط�*���^s�M�=eB7��۠	�^�ԉ0Jڿo��>rK���b�0Cl8"�Qθ	a�ȏ죦�z]�@1lÃQj�ܻ��f��O4��C��13�ob4�!f���͙�}�'�=�,����z��FT`t��:c�B�Z�A2f4�J�
`�Σ1I?FK3+�������w�-c�Tr��Kq����v�H�Dɵi�mbE��%�� ���{~�^�^~?o��q}^MEm�=V�q�!.̛}f�KqwU\� �@:�D���"��R�P0oD�0̬b9o휴V�n�3�-Cl�Hm5a=�Ʃ����L�J0��/C�F��/�+��ڬCQ�c)6o.��슨`��Ā.�ё7P�#ee�Q�#-�([�+B%B��<�Sj ��>���:���:,0��Ү� g�Q?�P0(iUP`�E
���|�b���m�D�9H~zcb�^�/��>�H�f�z���\�DI n��e�����?Ӷ���p�G,3`ǻ�Y;FN��;��_�"0�?��8���%��?|���R�դvV~�|s�}{����C������P�貇~D����疋�1"���Y[.D5
'^�F�J���WBg��<nv�&mMiM���} ���ڪjR(I�����>��]����o�j:���/�ЮOU 	�����I�1]v��Jv���t���	YV�Pծ�mig�I�]�ѯ���o ��bTF�%�QUF;��V�= ���]q[|��TR�W?�2��--$0&4=�����'f���R���� �[��r��@V�#����=����h@Sf���~,���ӛ v��A��M�n�X��[&����.c��O����
�����tN�t����HUFY�q�{�C�� ;9�����&B��ի��\Q3���YS�q��⾆��1�m3��Ef�F�w�
�h����&�NE8Isl�a?pq�Ǣ\�ְr'm�>�a�ET��x��XH�w��J�{e}�q��!g�A&��]H�7�V�#4��(�u��Wu'�ΚJ����_�ˇ!����	h��i�ƸJ[z�?�q薢�U1���׎M�D�2��p�����W�p]e�j^���7�.PV/A���}7�X]^��w�4���@�wV�NC�<���dҤ2�ۛ��>G��+D�Ԙ(���W������Ժ��]M.�1�	�����7�*��1�
����<��~���bw�{�Ot^�d�+�B:�7��x!P��a?q
��,��P4lU�-�sZ`O��Vb���m�Vȟ��|���$|���=p�����T�-�=r=s���"+���~2�K���0�D�q���2"(��J�Z��e�79�<��M��<2=�%o�Sڳ��כ���H�5��������É�����n�f����)bF�����sۭ�c�����c"�����&a�_B��5�p�}x�Lf}��V}������i��S�G	ʽB�b���9�0����K�*R�8���6C���=�S�g2%�7��E�Sw��I7��ݎ,O��Z���s���¶O �y�-�>��r�~�����\�k���#�s�����޿�O�6Kz�J�����������5�ic�S�kn ���,2��5��Oψl¦�>&뉀"m���O��A���c���:�s%�����-�6)���4����O�:��,i�@��VA�ٵ�U��{;��E*;�q�pa���A��O���/�+�	�+����P�{q�[�1dF����ϨUzI�8�Χ6K)���g�Q,(����J�����f�3fw����=��:`WU���������җ���S%J>�$]yc��K]��CK���4B����I���-r�$N�b����9p�lV b^|^��ȗwo���8R��&�X�MG�������KczB�}���t�� #fC/�?+p{_q�ew�8�h�4��C����h�t��et%�d�b��>8>Pr<�������s�`�9UUă�{�(c�wS��A��k0��Z���PE�ߡ�:�T-a'uHťn�_n�dd�o�#9���̯R�����,�O l+�M*V_�V���"�r��U�d���B��!������1�����JR�ADx��Lܥ�@��H�n �̾U�^~�`����9~>���c`D~F���9�B֕d+��'�Ӝd��>��qn��N��}�cв���[T,�|� �����Ԙ#K�nuê]>�˞\�ys%�p�)�n����� }�G����m�V��5��p;�H�_ˌ�m�����,o}�S �����HS���FzJP}!���mf1�4�w�7g�@�I��\�1������}%-�r�89�&(�Nb3�<�2�t��X�7��u���2J:��\߀�`��,@_�/v��ҥF0#M?�p�[j�啽4ȩHOZ�H���v� �V߃ GX�� ^��;%�|�TC0s:��!8	ⷖiS�ữu�7�Jg��Γ�^c�J�A�� �2U�@(z�]�Y�D87$�A$68������#����b���M6���A�h�0P�q� �s:»�l8����:p�� 4
����D�^�
GN�#�b::��� ;X�2/�^���sTǗ���8�T~���&T8}����Ϳ�QVZ��=�t���z����I��M׊����RMG(���fj�qWe��C����� �YٍM��[и6N�J�o]���Y���}:R�`�H��-�dz�*sb��h�t���]������h��D�pN�i4"u3�5H�¤_��d�	5�����Ē�/�['�Pb��<`�=Ĺfy�-�}�b��O�=�A��6îh�<�ao��4�*���ţO�4���Q=$3�S��'��K��xBS	���"B�\�3zvu}�3CA�����Փ�h��_�s�z��S�"��SU�u��p��<?����%,��m���٫/�E�.�$T�	~T7y���jc��R��(4z఍�����q�Z��/�w�|Q̛�J�E> _�b�Bޚ��Lj�Z%o_����㰾j1�U%s�i�Ԃ�ռPן��\�v�b���T��UY�Ӽ��!w����<���ν,$��}&���HO�j1�Ǚt��B1b�l'�t��KW+ǩ�R�Ӟ�K�c�E�V�q����M-$����L���mOZ9��cµ��y�:R�[
I.����%
@���B�^c؜�W�+j��v��Z�t��ꎤ���Һ�ݙ�!�N�L�� /�wU�˵���m�~��]��hT��������l�9��/	g���̳�+(��_�p�d�Q�h>�VZ��p� 8�C ����2[J/޽��e��E�U����&�@b}g�0�kѤ�����'�9|S
�K_���BOsb�{�K�ML�����x6���es
<��)A�/�=������	.!���L8#�l
k�3���bYw�I�u����Z�Q����Q`Q#p��D��F�#�pl����n�?�h>�̋Ñ�X��y�J�#�n!�V4�d?����X�Y\�]��HzWTMEq5�](���8^r�{aH���R��ڛ"�K�t�P���_�u�4s3=��\��nj��#K�6x������˚[�/�7K;�R��4�q�Y��C�o3h��t7�K=��g�eet��	������u,��Jo0�)h hן����5�:SrD�<��T���@��=	^�ܻ����� Ԅ��V&�NjYE��e<<�P xg�I������mw���b�;��S"�d$���1���}jooo./sz�"� `�&���:\;��Z2nS�[.���p]LH�uN˛��
��H��)#����Qo���r^�]9RP�]�l�g���c�/��M
H&s��	�p����j|��-�{*��#�Qc�B{q���,b���2r�LxP~/�@��@���Q��u��E#���>�_t��F��RZ�*��?��T�Q�<��~�f��� �	ݢ������TQDi�OJ��nV"U���y�����	��H��J�	�'7�e��W��
�^�:~u�R�\�C�󲄧
�l��W�
FY�Gg,��\R>��N՞L�~Y�G�L���1��������f�L���jՊK�
�|l�y;-��!�?ò���N�V��n'���t�?H�$�L�-s�$:�#�G|.��h��@,����b����P/�9�gs�b^_|�M��:r�]���p��FG[�`讍��,�߆fɊ�2:�jv�����a�	e?L� x�i���-�t5���~V{!�<8�?��L��0��Y0w��
�w�X�,����NH�i�0.lU��=(
)����Ь5��;��Y�n����p����� ���^UK�,
�5u�S�H����&*;�{eֹ#o��'e�3d��	�!W ��pXc0	�i3���(Y_gb\
�՝�gp��q����������RS��IL�:p�YI�E����PHl@N�/lj ��'�)�񐔑���� I&��H�s��t&��9vQ��Z� vin_���M�.�k�`�����mn�m�^���|#��1�	�:�Ĥ���ԡ%����o<�1C���!e0���}z��[Sj&ŌdU{6�{�XC��s i���rٱXQH�7w9�7�L�>C�Ξ b���c���N�]����Y��R��Cu�&S��]�B��V�1�Ɍ�:���8�e)��9��>Բ��_g�gꛀ�O���9!�2��/ �~���L.��Fz�k��[S�Ѓτ����y={�6��,@��+�T�t�uOatF6������������9�� ��A����oIާ��2J��k��ҕj��LN���=�ޗߜ�^zr0�H��m���%�l��]�u�i���?��~.�yj���>�ه�H�8��{UM=����|W�(op��]�0�����k�;٥��á"�x�i,��.Nv&{}��	#aj�
`���,����Io���E����F�mR�$���my��\��r��kl[�Or�]D4��9�h�]���hy�y�Y�������x�=K&k�ϯ�c�}+��@���ƽ�c٤ b�O�N�����Ɗ�w��=�X�z�qC�*��x���럹	�38�怘.�Af�"0>�tJ�����������xL'�Z�F۰�m�f��ִ$���[;2�RO|h�!�����`Ǡ�����%���