��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�j�� R�3��8��ji	jXo�֢�VM���Y��JK~��vm��J\�k�*���兮М4�<�op���r|r����C����:շ��ծ|[�W���O:I!cm�]W&
kx��v��#��ށaf��*�;�\����d9�D��XE�����(�b;oν��o��g��Jޘ?��SL��F�d�u��7�j`÷0e2ŗ��J�$H�pWҩ�7,�ګ�ٲ"P	�c��\I�\���qT6���L@��()��WPÏ�p��F�jF԰��"�Q`�[�^���@�f��P�X����К��	G��H~@�F�L��E�i؅�x�V���ӛ�iF[A5�������ǚ,?�T�i���K0Y̍��:��_���r��2}�qM]{u.|`#��N�xD����e���E1����~~�n}� �Tj5
e;�����=7�"hU\8��P�<�`�Eܙn��ݵ#���1�]�Պ������O��ʾ���]�M);�jI��h�:d�1�d���"��5���C��:�X��b�7C�k�jXA��R�J��|o�E�͘q4j;�� ��JXh_*<�����*U\]P��F�+5!ܧ�m
� q�C��-�DYRR�Yh�;�zJ&�x��DÇ�M5ͮ'՜c���Wϲf5�w�S_+�l��c� ڻԀ!�[�(�h���D���r ��R �ퟗ1�7!�=��ض�qk}Gupx�f~�&R+��1j�Fz�w���0��9����H�v.��QRpVb���M���Z����53v/�&M�,4����R�_��΀�@x�Ť6{��cH�9=��;u.m��e)ʤ�绥��ҝ�-Ql�K���R�>ÍMe4�������#js�*���(p��@Ґ=NC챎��`���֏f²�0+x�Z�{�m2�L%[�c#�J�[)g�)th�g�/m�5iw8I		��l��]���ع��{���J���o;@�A�w��%��E)\S�)	������^GQ.�h���-O2yN�q؎
�g������qO�R!!h#D��f+�� ��O;����?F�&%!^9!c9�����5�1ܣ�ٛ�3��=7�Ji�3�lN��Fb��WdB1e�����1�{�{�3��xg[+#�@B�&�ܑ ���wYph>͘�d�,�=s����a�Q���K�����;��a�"D�u h�2$pff���-���0j:���l�^,� �*�mNt6S��vn�"iV�����eV�$q�8r���na7�(�VnK���f�t��� =�q��e�i������"��5��t����6�������Y��F'm��+`�j�PJ�5�	�{�5V"�k`;�碯��li��JL~qd��f�Hl&AO�ۅ��WF���FO�8��Utg~��n�t�������h��$J��h���kL�������N7-Qi��I�5ub/���3�����#<�����W0n?\��o��L#R6�_����Iv��\��ѯ��)K����;����^�k�Li�A�m޶�<��1�aט8G#GN���C�<i��ڌ�n_ ^c6������	4`�aP]�qI�0�"�@��Y�x����V¦���I֑U�1$~[��=�w� !��:s*���zj�?�N�"�]'��0�P�&���Q6��@È�a�#��Wb9�.��:���a�2��?��N����dd��φu������؋�W+�<D̋R+C��X�B��L4|F�k4��51�[$�=��C�5�	�導q�+�G`�'K���`�:�7O9$�Ͳ7R�����<���RrZ�����f��?(pn̉�S5�
�{m�#5A_i��_������l����l���aN�𜉥��4�R�l���I1b�!� )U�d>
]?�ZQ-�~S#���TN���ե�����Z1-}�Ķ�f�4a
�'�<�Z�f�,�y,z��/���Ơݩ� �~�-U�/=�/(߰��@��a�7(�z���q��`<��rc��H���Z���/n~�;B�St�v����x.�ls��6��ڮ��Y�D�Zfp�Й��⪖�;��_�H�Y�++H�:)&T�����Rz.�nEM�;�~h�=;����I{�'H�����z28�P��|xC��]x�a.�2��kЍ��:����yQ�Hm�>[��v�C�c�b��REl�<-s�s厵\�����e�5��Շ̌��G���e��)q1(i��e�/����յ��j��(��%��Z?zMN^ѵ*��T�E>�=M�� Y� �xё������B{[�ɠ�x ������[$A�1G���,��t������+�i��i������x��e��%�՜�EMT.E� �BP������k��+,,�ɸ�4y�9>��DbKY�V�}�[���kC�(^�R�Z�S�;5�G�B�H�T�EXI�,��6hF"���x�:��  w��24��&��		�%�_��ڰ�eP
��givM�d&r�K��R˻� �I�#οY�8���g�=Y�y��E��ļE =˫�rG�p����˘F�c}3I�|@`_�-��w��&S�U�<`��gm��`�����^30�r�g��>x`�7�������w_3 �i-{�ʰ�����cJ��=,��5�"�[��->�?�N��|�KM'ó(�laӎ:Og.^�e���ݷ&��8����'��7�����trT��cw{W���0�?��8����ʙ)'q>���f���p4�nbuz�GWG�C	o[��q�V�uO�q�Dd�Po�����0��QDy�2`c�E�)m��xy�Cc-��&
l?��K�2��q@�Q�}��r?m�)Ԧ?��_�x챾=�����İ|�(���+��,V5��ȝ�v�	�H7 B��N]�v�N����%��;��C��+��/逾O��������N)Y�����D�K�
o�����P�O��������
䧜�� rnx�Pd�S�6��>�-�����s�f�	���G��z2m���Db�n��yɆİ�0w���jc��CsQr�rIS��0�)G4N��L���^��>s���y��^��!�4�a����T��Ck�;����7[�B\o�0S/����lM4W�)�gK��s�]�;�U>�����A���{��2�zU�7e
m���)�G@�ͯ�yŞ��Q��A��"TG��as�����K���RI�YU�tֹ�Ϧj��W��W���:Y5UW�x��q��T��R�6�[0�1D3��r�q��Fd�ҏ�̀L�t�
q��T,��@��Ǩ�����B��Fp��y�C���
3n�܃[����c(ԅ~�  �r�4d[����Mê�9)�;1Y�sgW.�jH�<K�ᆸ2���=�e�Qo"Q巄
�|V�eZ�2g�G��pN�ܼ��P��KĠo@�R�{~�ܛ��4��Wp?<j�K��S>���$�
TX^���߷���`