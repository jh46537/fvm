��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&HI�Alta!E`���Lm6i�^Sn\�c��I>~��~e���We�ُ�⍵� ����k%�Nna��<�kv�x�=s6/�Rp��_6��h��A�g�6��O社3�XS�ݻ��;͈7L�-��^n`�q|ڹ*Y��%�h}�B6���#���'��s��\���n�y=��!0@%h-�tt�p\B���"yҒ�:��h�]�
��J�;9+$Z]4D&���~k�ڡ�z��a�jGӶک������M���)��h)yo큙l-�|���PE1��:�ozc��HH97h5�ǁ��ipj݈&�B�:rZ����0 Ț��U�?��ف�Q�j����+�J;�����ytK��G9P�F��t����st���oJ@47;2��'"|y��`��w�`r�+`4}�
"�f��(HT�VO`o�.����ٟ�h�d�U�@et1'�B�{h;4B�#�~�Q�g�@��5�r0���� 6�:$���mQ�$��z��˙Y���A�.�t�M��몟W	��>��y>m�L�M+e��*�g?��u��6�+��\�y�I���.�Ʋ��]�x|�=|���0�"��Q�c�8X�3�t�Z�@���P������gkf B���qWyw8�͇��rwcf&aH�+�@���lĆ��������?����m�C��i����V]��9dSqJ���Ͷt��	E4�bh3�u��h�[w]���X)�S�ζ�(--���N�E��R�:�ߋD�}_�+����5:	$7y�in��E���7��1�_�i���'<5�K�Vf7�p�w�{&Y�M{Ƥ�O�(�aY��t�v����B�36V!R:�/����W����Z�/���Xn�7'��`��|,l]���ݻ��2Z��2��Z�e]��j璦����y=���j%��l7b��:@.�k����GI�����'?���_�C�SX�v��W:"��7�iA�<o�����aܤ�B���?ye��A���xK��I����v�� g.I�:��[^�Ns:`����k��;y�} �J�c�L}q?}:a�v���pOݗ��C "��	#�J�Ȏ������_ ҟ}J]��gS�� 1����K�f�5���ڎ�+%�H��c��V��f�I�2Ia*,id�
�`�>�J�G.^�Ve�b��:��/y�H.������0�7_JX�D�o�-��ځ�Em&��ȟ$���`��jj~�4Ik��D�ʕ7_��A#݌�#Vl�r�Vj�'�`�\F�k|�ЇJΛ��F��(
���<&�4������������^�i�����#�n,�/�	����t4��m���S� ��x��ۮ�������"-�#i/�:�Z�� jk�:2����� 5$�??��4~b�d*���Y��v�7g��3�<�=�z$���#q�'��]G�Y�_Akk�p���U/�u&�Kk��$����%)Y�C�t����
i���Q-1_���l�/}�aS4!�����l+B�}Y�J&� UH��y/�hAr��C. ����7I8����3=n�	�w�J���f�*,�����{��D T�@�CEA9L�(>א�ڀey7}ș(�[���)i�Wi����Z݌�x� ���.Y6UЂ��-�7b�_�d�J�.�O�� 3Ð�Vu�E��o��^ci�&���6l��ݰڑo���B������>����-e�^K��*P��J�r&bY�N�[�0V�&i�Lᝯ��C��� S�j��̏j�lb��t�P#f���/)���E%A�?�gh�����H9�z�O��t��Wm]�7����N���G\/C�^�cd<���5UA��zF��Ll� y7�D�0�n5\��ꯦ��N��ҡ�dY:2��K������O�H}����x��G���x�H��9Ѩ>wl7~����3�6�~s-����0!�;H���k��j� 2�L��4譀cŅ�ا���v���ɍ��t���MY���y����v��w}��Y�Kkʑ�9')b�l9]�Y5�m�ږ,���J��2��糱9'O��n̮
��{�]����E��!J�jY��9���pA�+O��mj�>M3�j�A�q���o��T�'4o����F[=�����¬JX����$��3ų�9�����-�U��܏?���-&���r������.�QC�
t�V�=�֮5�Q��k �l�t^�:�+o�or�0�+�5>�L��۩������\�:qX�)����� � ����EE[N5Y�qˮ#�)0ta�af��s��1b}ܴs�[avP�6��	���v�ݼ�ҩԴߠ��{<��l�"���#��D~�kj�U.A�!u'f�� �$|�u��.p��E���<=���9�+̨�{7̾L�*6$k^�
�J)�55��c���4ۆ�����p]g�Qt7݋K�̐$�I��T�W�����~�a�g3�!�Nq���.Lu�o��#��P�n&q���GRaI��(w��q�����,��$$��`7��ݪн��+#R�G���MXE;�b�&9�T�����_�"�MC�l(��P��<�O���[P )�D�[[l��t'$�1;ca%��442����GiR�"����I�?@Ń�j^������n�hb{�ъ�W��n𩀏\���`����E���>����N��K�lC���;")���^�dgsr�"Sb�+�i�i\��Q�}C:��ǜo��"�P��7�X����x]�ӥ��:x�#��i;3�O����u}U+�P����m�b��"I��CGH�v��`"�qS��N���h�X��Mq���S���
�F�uЉ��H'7QR�N��7ۑ{2������$j܃M��~���D-�u�M%��$`�E� �)}J/�4��ly�!*k<�������b~�SV=l���Ch\�:�YUgK����m�14|�]Ptj�D�
�LG"+��O�(��t3��i�ef_ڻl�Q��(kU2�W`�a��Г7�q���7$x�
Qdw㞇vnPO��VrC��ɳ��V�׮��moH��o��v�;�e'B�?xºg?��T��"�(D��D�}�.P��@W4�/I	*#�����6��|{���9sY�GvU�i��qc�G�4��A���E��4�辍�s���y{{��c\H�+��`���A�c��-�]��S�Mem�!}�^N�y&���s�9�_R)
JJ0