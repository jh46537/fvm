��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ�P�H���
��l���Y�󛳅���.�X��}�X�����e�O={�9�����Q6~s[V�%^
>��a���t�f{�Z�u�Z���	v��3t�mW�=O��H��si���X���W��=��&��K)��kG��I�1�)�
��Ls��_BX���~ SV��X�$���6��P��Y�ۮ�[m;���yjl4�k<����g�_Ԟ��(%�D��0B��z`Ąu}�$	}��(_]~;ϸ2��K[n�����#|b;>���V?O�W�z�95+�y:Ac�EA��ƭ��7\E�q+�?dA�z��72E����n�:��YU;�[�YY):kC�Iۉ2������:�Y(���3ֵ6�!�|�5c�Mo�,�5�IFLjZ͛��hvfCp�����G����Jh¢vw4˔l��h�C4�|�>e�Ҫ��s\Bĩ�x���p4?(B���1޷�����w��sG;�V��y���P[��T��uE�: �|�ȉ%w����Y�~�+� �N�L�)��`�ۏe�GM�4l��"�UD�j���9^B#��k$A�����/ȭ���Vp��,��¤:�>��gG~��>.��~E�:?��u#L������,��ن���_��RTrxCp���u��^~�������SaG˂6wųf�d"�A�BgӰ��@�,�P�w!��Q���:��fP���o���=X��o�"�B���p���C��%Fz����v����Y�:������e�/�!��S˽����r�B������W9�N��
I�y�$6o��!��=,����x"-����d��ˠB_1j���\�@(jY�=4:3��'��/:�k{de���ӱ��.�|�2n���Hx���]|��3����ņ��=4��X���&�ᗈ��E�W���r�d��^n�h`��S ���=tp"ǅ����}=S@�S��� �\2�k�W��`H\���W&�#q�´_VFi)���}�����	�	�,r2��1r�ﶄ\+��MĻ��C�����%o��oH���?#�*v1"ELB�\���[�Q&�S���>3>�p52���/�`�T@KDż%,��L���>~~�2�Lw[����ATY�U��Z3! ��J�;�E���s��O�Z�,��|$�.o#\�L���h�2�>�5�0�BPO��|�t�Z�_(�J �}��o0qW�κ�1r�1��������-w�o� ��XP�*�{J�	I6G� "��c����@�}��6��L�|��#�0�{�|S;�(�k�FiB��i�st��ʉ{q٥~J�*�٪ݠ�^M�|H�����WLrޭX���
yu�(������IP2��!_d�2�M^��Jn,�0����q[��Of��4<[�sH����3,vnwl��&ǩ��P�����o�Bͷ��֧��b���4ݴ8Ant�-g&�`4+�>8�krd�����R�Y���86�3J���}"N=��(	����-4U%�����b�4w�p��ds��٦~����km�|�Ô{�5R�+���h��?��á�h8�X.7h��x��q�v��%[��&l�Sp�G�LO������\˗�@/e��:����LKxSX�k���+.T��9��IT$�#~M�`����vJ1����ռ��jRUG�jż�>�CG@N�dxFw/�}�䮁r�^�%&�CE5��5��R�C8�d]ڥ\�W�ç�-�q�ڪ*��KWvT-y4�CtǬ~�-ⱅ���ٸ�l������$���w�w��d4蒝Ȇ,ƳC6�$��9yhs��>��be�p��{��03�؇Ȫ-��C9VL���(\(�<�U�Q����(-����'u|��B�F-�FC46��$~X-�}Fd�p�zZ,��O���,�F�u0>�ށ�Eg�w��V*�[�3cr�G��?��VCgG�H��]#�4�3�}]�b'�r���m�!��΢%0�)/D��(f�9�Y�5rA`�P���t���o�����,K*�^�K��!0?�s�p��D�[0L�o*rtd���ݤ��m,���فt��A\gJo�\�Sad_'>'�~��MD�Sa)�0�뙗�u`7���u���h	����մ�<n�� y�%�ϗ�B�����Ɓ��x}d`���k�tk�a����R5(F�{ k�Bo�^�۰Bԁ
\�&=����l(�<�I�]�]�uSC��r�릇q҆�����E�r���͘�$�$Y��q�O	��T�%���J�D�AU���z�2��13�X�K8%F>�
d�})���;�NT��6�WJ�1��s��>M�Uĩ�~���oX#��s��j�c�t�M��+]RF4���|RN0)ǽ/�em���'��M��9��f�m���<��`�B��3�f16D74�#��s�o��%�q���]kd�(�ݡ\�����9������C��!~U�F��XsHM�E�m8%�n�얛�����Vg�l��Y#�qݱn{���D�yp�,��n�v|�@���-*�yi���	r�,r���߂Z��&f���RZ�0pO���
��y?���d2L������v��%�V���I�絉�
\��=M�vm49�r�$dؚ_�8�{/8����c=U�E�?� \��PS��~A�����Bd�9+����xj�si�?��C�����_��h͞Uo��֑�>0TD/�ʒ��/,��'�P�!�����hpfa�p���h��T!6���SJ
�؝V�ۻ�'�}�y��d�#5"WvD�F�*����Mt��'���>�Z��욘�p ��#�4�04D�{��_A53u�B��}`��~�A����؎C��Q����r?X����5�p�?QV�֝�l�>��A,%��v��Z^ؚ��-�{pKT�@�]�xmF����.��`Ҿ_F=�s�D��/+*QR?���D���}$��s�(#�2N�F�����B7�q�UdN��N
�P�w
�>w��ŀY4�����GVfxܴVK2��,�n�D���brNM:5�c�?��4�<��6PV�vT�ǡP%�Q#I�O��h$Pۚ]
�H?+�{+�'�����/JLQ3hz*�vyG^����ҕ�lh�z���;��Z��m6�c]�Ad#PM���f��+�&��O�0��ux�Eڂ����L���r�9�/�����:)����z�2�&f{MՆba"�f��P��%��>4�5�Oi�32��R�Ș���(��62�� K�t!�����\	d��QB�?$�Έ,��#�<_t�r�!��;�	�{����Y�Y�tۉ�|�>H[<c�S{
W�ɤ/����7Hğ�֖dNu�Km(�n>�����iht>���ň�����X؅6T�BΤ���..���������8-~Xs�1|�YX݂�b�^2D�S��7�U8oj%�����%a���	2['�s��q�^��lv��5�vG'��T�2������e��\J~"�I��H?��"<���P��D�i�NZ�Z��6���r{.��b�~�������ծ���E��8&�1�)c4�A'K�h���]:{JGC�p,¶M�PA@�U<"K���kL�,�+9���U��.*>�����)B�+F!�1��_���0�'�ַ	�*S�ɋ4_'=Z�	��@���b{��'\xV@��h����Y@��-�={m�E�5(1�p�T�C���6/���&��w�F���~�VfIn}X- �~;�2v��`P!�hŮ9TQƋo�_|�3h�%�+�/R�-�Y���H�c��WTe��YT����*rMߌ���~�8`��x���bf����t~)єX+-=���E:�0F/��m�\C͂%|]<����P�܌I�gm�r}k�cX�D��+��4�}�A�)tu���`nq��kN��F*�