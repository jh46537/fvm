��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�w�\պ}���'d��qx�Ba=��1�@t�lo�ܦY`f9��GU��O����5y�k�wy5� e%�iHF�K~3��Z�������# ��d|��̪�����PAZ:�;� ��Փ�?�}�F�ԙm�-r)��]���m�V[��zA�?�p�,O�?����5���dk�������'�]��i!������&4s�����	�O�^Ȉ�i�pz���j��;¬q��"�޺A��+NT���2o4ƙb��fZJ1k$$.�,��C��{r�cD؎ (�>A�xq�Ou�"f�X��ٮ6e-��0Z ��*V�7u1��y�*��w ���Y�92�<���?NS�	U��؆��p��l�VW��O�"֎��CVt05���?*v��*bi�����2d8����/,�`�0(fb?�v��I@%�S��%�Ǎ�^�ݽ+7��Lǐ:�Y�oTq��iǼEOf�x|V�n}?k����ede�7��&*)>RecF�Ƥ��p�0F3�j'o�0;;�6sWN��rR�a�d�l�����^�|��\th��v�ݓpi�F��ql:�~hq��ur���(f��T�[y�/o�
�����3U d,Ryb����z���L�@����-{�	5����HÑC��Q�`>�3�2���I^M���0V�0� @�s�=���e���'��ª��k�8��k�c"���{�L�����n�9m5/D7�N��!��G���D�5֚�M[��
&�BC���	�s���D�a��bϢ�b��.(��!�%����cI��Gx4�C���	);��Zs��k��'Zwʧ�+�
=�� �u�������A]��;lRW嬋��`��K�t�x����=S]"�m��]B��sD*ΟB�ͮ:�,)������t�&�-9�o9jj�y]�kR@Ǚ�	|�!��6R���To���	�l`�v5������.�e���-�]#���.�l�h���-�MM"n��	CpՀ>ֹ��UT�E��pb��<X讖�$p��T�ճ�c�g\: v�Z#<���O�����o%B�F?���ړ�-0�:ޯ�wh�։x#WP�ŦjiH^08��K#S�|6W�]g� ��8}��d��brH��y���4���pz:��;��p,M�AI,��! 3���r��|�<��ОP��BT���#��<�����Vx�.Xr��M����k]�� i*u����E�� 9��ߤ�<jq�w82�DuA���d\�����J�:[U�Lq'~Snbꤛ�Ⱦ(�G��~�� �xv�E?�s���鰐�@��
����3����4+�p�x�2�.g~�r��H+z/�Ew]T��R!���B#i����%���Z�3��|�1���&x�0ο�6�_��_��,��h!H�&Y[wp�޶$䴡�s��0�o]5�I�$��+�Q䴊A/����JLq�N�@N���V�xw=���Cٜq�_}�����>ϡ|�5Y[���� �U|�(���IMwg\7g���o�ǘ7wO4?��֓���M/2�ۭϝ��V��R�^��疐Ȫ��3�ޥ�x���:��v�Gt7gn_�*^�T�,c������Ǵ�����[R� ����¶����t5��f��4Ǧv���8�MZ���E������B�)S�
7`]"kA�����<Ԑ�9N`��(-Њ�b׃8�E���審t�~e�4�{���h�b9$���i�Q�p��nJ04����_>^�ϖ�4����![�5�D|>�8&�	>���k4�'�1� 3�%��ms��& �}8(���r��V����c� ��>kAQT���a&N���_��@��Bg1��Hs�<�B��ߴ��eL�` +{\qD�%�1B�t�вb)�6̍Gۇ�;��՟��Rp��%��Zx��7qG`�'*MH�~�	��,zgS���TU��E��$�]{�Hr�YgːW�e��o�m�"��e���[E ��1I���>��>�+���훒B�h�Ż&!?�f<�}��Z#�K���,-�;R��Y���2��_t�|5�`����1qk������:�՚p6i��*�B�5Bnio���K-&hL��/���j`6��h	�18�:��9;/G�+��� ����$����2�d������O�Z�u�+�!F���ћ$�%ג4A{q��з]%7 ���&0�:��e�E%%^̏�mj�JOO���B|mIFV=�V�/9���D�?��dP��7
��@A �S���
�7�ͼ�x����[�L;�0ﺝ�ꉱ
f�{�O!7�#���'�IÛa�5��Z��fWBL"��*E��X�4���uzXh�ij�n$"P$Z��X~��z���l�v��"�l�kd|���Ȭ��&�A��>�p�9��&�g{�׻�2e��M�-�3���}{�/ET�zGO4s���;�~Q~�;�pz�PH4t7�����5L����.��������S�K�l�Vr�,�F]�<O^6����y��@��f�F���uo�'���i��:ƪZ�46h�Evy٥kW)�x�̮B��$��}*J �E��OD5}b�㉥������lU���X2���&7uk��q�Em��?�����C��i�#/˜O"X���afJ��0�d������(1�B�^��$�@_���I��a��Z�R��h.0��/E�o-i3F���/l�x5�5g�%�g�1'�Bd�)�_Z�v=9�zg�����ۋE �V1A�ϐ����Q� �O�v�Na�4�e�C���j��Q,�g�6<���M��*zJ��)F�Ȱ'x�69_�N\ݤ;�Y�d��=#���z%����x՘�\��Yh��N�F��
?ն�����8�����ז�hd�3O���&��j7n��R����n@�$ԗ↧-c���I|_�,��2	��Ԓi`�`2؎F/�M�"������&r��U?@��\W�6���X�cӊ���ƅ�R(���B�z��Ӵ�v3��������|���*~Ѝ��y���;���ֲ���y��W.��x�0�w��cz[b*�������W�].ut憡�F~��l��{އ9��i�j��B*�@�8��ԯM��K��k.��┯l �9.���� U������-�(������K�$�fxe��z�����% ';Y�؆�	ݒ��R���JT��d¿�4L�#t�1:3ug��l�/�V�n|2��X��o���^��Ⱁ���䃿�>�����W�2�О���\�.$��@	�����m��+h��m���m��o�G��o���q΍�OE�?6f�@*)�C�����D2�܅�̨�'�"���+]*k�����1:�mUe��sK��$1�
�/���9�x�Q�o����sĀ/�}�,��C�!>�f]�S�F����#�!��=E!�k�2_\�Ǟ?(E� c2+�p�[��qZ)M�݆�l=��ku�\�=/"i4ny���	բYL����2���W��ܝU����,��G�J@��*���Id@F{COL��A.b�Wc��T�Ӄw>�L�/Zzш�(��T��YFģ����Xw����oF�qc��"�������ڀ诸vWG��%���@}���9h`����βG��x�U�ц�M���L}C&�Er2��ѻn������S�+�H|wnti��n{4t=�
\q�= ���r���U��>��UAΤd푱6��̻��H1"Kǿ9�	�7���? �s��E����I�������'1"t�1��d:[[�aC��ѣ���g�\8��7�h�,�Z�����{���[��]��C�1F �#X�`i!�H�k��y����iY��#��=7�1Y�}�˅fy�6�I�
ß��(/ݔOLeN��߅����_qK��<����Ð����O!b8�8f�^_�e���l,��*�v$Uޯx�u�'�v_�3�/k�CF��o|��oT�*���S	�e vYh��Zc���>=���="�3N7�T�eǀ�>�1���@(�hԁ��������j�I%����W��Z���ؿ�����W��A�5�<��>aVb"i-3y�`ON�,��Uqk0��A��!M�u�WL�O�>�>��Rښjȱ���z�@}ʥ�i Q�#�g2d���A�UA�i�������+3ݑs�n`�.ܞN0�:�EŷM"�?��g"(⤹N_4Ǌ�\�� NTW��tf$Y�8�b�ʫi~��cn���v���䑈��T3�+�q�:"S���T����F����:(~h��ִgʟ��&/-�q�Z�S����U�z�� ݐH�Q�����Ϳi�{?W-���n�PWw��������=��H-�uԾ�؂ݘ�]���:�*����r��krQ���>��XٳH���1�Ё��$@	��(��?�dcm�)�Yܮ��OY�1�&A�9�}�5i���_?5��0�b�e ��V��-�o����4��`|z�r�;T��U��n�R�e*��q�C��
1e�Snw�ņ�m�� Q����z�?��Ԙ�%A�����|�0��8�ƍ�va~~�S	&�����r	��>����,5o���	X�@2�!�Q�k9��p;���"�]�3�@�ݖa��I���F%�uS�	�μ��D�2�cU��J�T���m���ٲ&^���B�8m��X��RLO(K3���7? ��Z�ov ;���,����E[9�����.��`� ���JunI1c��	Q
�-l��uJ���D'���
$Ǖ���u����zPnX~"�_�X��J�-溝�LͩJ�̞K3���$��s_���3�p�A�(��3�"��Xy`��W��L�r"f(.7�WI���+���
��}8v��J��=?rt����f$MimI�%5;(WE�,�ԌM&8�;(�|v�%1� ��u�J���㶫9�~�-�#U{X�y˞��d���,�hHڰW�v�HN��3��xM��w	�.������'��P��S��g%������@'��z�LOX��j��\�gxw��\9(�:)�^8�3:�:NMF�9m�jv�4����52%��6Mk�D��0�;[�i~cgOaǤ�I�u�⧨�%��Sq�����D���"��3��ߣ�#�JDi���m\�n�̴�Pp�6Ұ\�/��J���Q��r$$� ��&�.}!�H8{g����
�?v�|�e{:��CBc0���S\�c��f�qG��uHgG�n�p���sa�($��<�)��>n�o�9��&��&�L��o�2v/I��ī+^yCW���_ף%���K�9���p�f�<�r�_�4 �xKu���a��m��
�8-ʐ��Tԉ-\�:9�IJ�D]�%�'ٙl��+�o��9���#\ ��tr��=dk�r)!r@M�*p��i�>�����h��M��`K7LѰC���QY�	X�?�����}�>�c4}`Sg�	���?PML׵�GK>�q�S; 
��q_<]�n�%���1���=z�t
�6 �+u!LK��	�r{F�B}�SJ����w8z�������W�2��L�gTTTNmBc�����B�[�V�9I3^���[b,Z}��J����NC�C���J"[�<x�<)f�5R(�mw��� Tr�����	��l�Kp��ep��B*ɣ.���0���p2ƙ�Pw1��葢Lg�&J zMdF�E��s�� γ���<�VF�����"����F�C�4�a2k($V��R=�ߢ�HjI����/�KC-��L��)##[�y��a����	9zi�4ȓB�����b	&3�$8T~�7#��B�0��L�&��I*�2�O#�f��~��bj�(wYE7�}`��-��������Hjq����[Z[�gQJA��{nr\1 T�.!�iZoHVR�1�O����w9��!՜��q��5U��4�~�q4�fc��%�� ��)on0)9.�XD0�7����7������4����~�$�@ Kx��e�Ë����[��+}U�_��y�!���.~q+��f<ؚe�}�	��;bʝ���tt���9,�����*�:c�FU��Rz*`�)��DW���jk�Zz��S�O�E5��UjY��h�����%#oؕ�C�_���6*9xǒ��^hP��y�@ע,6煫=���;xt��\{)OE��~+Q긔����K�қR ]:r��[s��\zG��_�<�W?���-�Tâp��)<S��~�������$h������o�i�u�v-\`p�	�d���m���G�3��.����B*��3F�b�S��[���E�Ȭ->�ʎ]x�,ZP�UQ�X����a&����A�,I��`.�Y_�BH1΃�����z_,� �=8O+�"F�� �#�H��:3��t�x��ί�A�i!��	�Id��"���s����2�+�вO-��U9npLkf�/қZ���Q�v^[��� �S��
�N�m��"8�k�!���
s����E��X�E&x-����N�j��h�[Ms����}o+�y�C�P��k]�H4�����������f�NX�A�� a�\Q���.��FK�z�����惒�I��Z�&���Ij�z��,�Ƒo	��?x�mQ��MW�wŜG�C��l��Z�1՚F�rI��v}�>&T�դ����x�S��1�Q�q{IXhdl�׀�Y�1�~ݙ�,�@�S%�#��9��*�������b�f���^� ձj��=5<���)��N��{�o%,r4w��U�[����D�
 ���{��YB��T�}��ԁ��f�3��jlqv�&���Ō�-�"ph]YP�(���,
�����7����]�4&a�~Pa�zqƙ[a�J-Jm� D�w����R\���J�ߔ,$V_������V�'H��䪴�������������D@�#Y��%�yU�g��z���ݦ�+�5�Lƈ�8�9�|��3��'x~�B^����}�.6��)(�bOs��d��������S��K��	�q����+��n��Q�#����$ ����4�<)��nq����㖝��և&|��շ�CH@���PEF׋�*�������%1�f幈j#�p[$�p��Ђ=��ޫh�@>��(�o���E&���#����M�0�d)��M2��a�v@"������Z�âq��M�:�u�t��QE,���)�F�<KH�/[����y{Po���g��)��0�����/���$�xԉZ~�����a#�?��-Mfe����A���Yo�����UWF�G���>ś���	�v�K	-��Y03K��T/I�?$�U���ǈ���� 9U��f�dۉ�9�1O�X@������i ���HI罒���:��/(�f�xk-�b܈L	~��w�fX�5�}-ٺ$�oƒ��}&B���,�2�<���"[��_VDU�qܗ�o��ӋCՃ^�J�Ӕ���	ڹt!\GM��h�^�4P�\�*�y�{��O2�ς�WN�7o�|���G��|�(��Y�o_�b�g��0b��;Ը5����c�K��z����-����{������QH�Ӹ�����@qG�L4��܃�0��/��h�e�K���
#?f`b[�J�	�M�c�1�"�z!D��J�`�����f3�-����ԭ�	�����Ç��gkF�;	x�h0#f�43O�s��7f-v���ض�W�K��i~ۑb䝳*S��n��!yw
r���UN��h��8�|�ӧٜ���Z<����tp���i|�����zN䏂���q�p��і;�Oh�D�%o?��B�j ә��r�O�|��볷������93^��XU�r*�?/ ��2����_�A�.��;8�M�v�+]��i�8�S��l�����F��m�r�3����!m8��{e�H���7����׉�w�ő��&�f�G�Ճ	�(�z?B�>���)׼�f�����V�"����S	(���w�1��ًԪ>M�)������$g��W���_��^$`�LR���b��d
��I�P&��(�/���u�H����!P�9�I��5�;C�^6��� ���SU��w0�1ͺ�S?:� /�굲�����7ּ����a�A�ҋ]�b�B�$U�PY�M|�n��5��<g���e2�wD�#�h�g��f�fB#��V�.k<�a��}����E�J5�Rd ��lI ��Vh]!
���K�fY��S���#S)�֝0��`l#��8�w���1c8�����ZX�8g�l�����?]�T�F�2���]�l���nuv��-Q5������r�DXT���߿u���U4��NJkB�]��q�c�2ĺ��S\�L�R��EF��G��R���y�TM8n�-Z��v��$�q��t
�D[�R���t��D�`nFa��Py-��8�%�j�Ɵn�!D�*�+��x��2Bj[ɱ�j�KFA��8���Ĉ%r�@֭�!�q�3 <!
ڸ�rO������`h�J�)K��Bc�3���j�C�o?G ��=�,�����c����߀�)��lE��/n�:��*i�䅱"������u�@�K�	E3�@�Zo�:N���q�|�H��laU��MA�%�V'��2���My���_z4ڱ���By�Ŗ)�"��bĤ꫚��|���d�{K�����L`�3�:*Ns�<7UȞk(�1C��������VK��Θz�g���n��oi8�Y��m��0����<O̙mM���E@�x����]�FLM�3gT5hj/�Y#���Q�/��$pZ`7���`���08�M�Sl���o���$`�w��Е1\�7V�S3���<B��R��a�O7�"�ND���S�[.��G�ʻ"`Y�I�ċ�oMen�s0�<"��6@��fq��C��`k ����CE0r�,6�Q�־��Q0Z���l�ǖ)=�h�@�=�&���Z�i�JQ�އL��"�7v��c�`��LX�����D�1�0'�P�2;���6���w�f9�A�ir�z��zMo ����΀T��V~|��7#��+>h�&�=��ГV�~�Q��QŁ�Ƞ6�5d���'���f�ۏ�C�Rr(:|v��4�A�{�sQC�'��uce n�R� ����KYF��@�K�;����5�j|P�+��و'	\�J� �վ&s����#,�ρ�jM!8,���������0���h�6(��g��'��n�����9�~{�$��
�mr܂�&�]����f+�l~b�#Sh�ǈ�����w���f���r��z n6��o�%���f=;��-sL��P٢�{/�$h����aՑ2�G߻ל��T��v�Q4^X��j���!�U�3�����(��~�����;n��X��dxS'��C�Z{��A2�0AV�p��I�8|j6�>Ҟ�nL�f�[\�E���!�û_YҊ�dG�l���Sc��C&lGYܜjo������(�H�(�{��S!33�Ż����P��2�Ed�,yaR�����=2��Ψ8�2�����(�=�'����|�z�J���Q�����)���ɿ�,n~�Ym���ڷ��"X�}}�,D�:�m1*"���_��<.)�p�x5"�AU&��ܖ�V+����Uo�0}�w3M	�M�m�s=��⣝ç�Ò-���|{u<��W�F�h�?�@�﴾�#w#�y!/�Ñ��x�*�)�r�(��@H�o���ו������g	f��BNܯ�����|u��RG������"/p��:+�{(� 5ГP;(I�m�q���"$x���N ��}Lw�ǲ��c��o(RC;5"IY�*�!w�$_G0&*'�T�G*�u�*�#o��/W�f񎨩�����ּᘙ+њ���$ O��(%��ܔ�VS3��_L�u�{C�R[u8�>#$Q�1|�
�?����;�c n�1�Ȃ�14�ݱ,Rw�ng�h��]�A�(����\e?�#�3�7�2��Z�!@�����e����Y�"yCyV�$�{��^��\����[#'�� �g�_.����:M�X����
W���X�+�2L���@�[��ʵ{���^nwp��7�)%Q����8���K�l�+�$�~E���Z����x�cW^��ڂo�ʧ5"h�����G[�P�������h���%v�^�� ��t��z"*_Pvz�jn�K�݌�&O%���}�B��Af6��YƉ�w�F�P�+��p=�:Z9��r��R��!��<#���0[oc2�fnX�Ѧ�>2H��iZ5M�-���B��?�U,e^ ��b�>H����ڹņFL䋏o�;߳ ��tl�ݟ�ܡY�@Ir�����H�#�I��$t�p���h�ix,�Q"g��q����p�r�#XL�y�.oc���JaY@Q�J�`d��dv{�Y�`e�_f�oP�r�n����lK�g,��rp/������*��ϳ�3�S7���p�A"�z� 7rμƖH�P�@t�ȣ%�@pV���|d��w81Ц8./i5�zuK�;$ �5��,�&�4�NH�I���<�Z\�L��B��!� t�q/bථ]z�~�7=��IR�"�VA�\p�\B�qv3��cqvוu�I��=^��o�:򏖅|�B3��.u
�u&t��k�h.�Az2&�Ʒm�0C�6�-x5
���8$q�)51 �_�~��wi�o�6c>�(#�?�|���P�r��*ߟ��� ��"2��/:}w
�P��r?�����M�%�u9���v�{��g���6�]č3�u�����Y��hn�g��I&e��m�b�]e����{P� ��(��b��g�.����jObl)����89G��łҕ���7t��1�h�?{���u#�d��|ٮ%P(����sǳ3Q�D?�/�S�6�0���\sQ�SzA�z>�� ���A�69��g��}yw����草�F]�8������eg��t�8�(� �Н-`:^ȉ��kz���Moc�D�h��P&�+���QR$�&%z�J}��9
�q�d���߭nW�e<��^7���?�ќ�����іV�4"�&�F)�t���i؋�26儝Skzϕ���vZɀ5�W�Y�}B���tYU_2\ �	��S�G�\���Yж���ݷ���)p�#ʹ�$C=I�d��\4��@�z�4�����?�P4��tLY#���A|�|t��㔮����l�8wG�N���r��O�ԟ�|!d�����qVx]gԉd��