��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]�7�%��	+=vJ�c���H��|��	>�6����"!���>����|dI�3uh���{���DiPθ֟��A}h��¦OR��ү���x���ݯ��cK�Q��;��t���冭,]��_�aI�m����+)���R!�湧���w� "���a�$�C�����lZ��j]����5�A͎�0p�읢b���S��T`XI�s����;��bk��@���B�X���3�o��kf�Zc�L˺��G�ʅ�` �a���[��~�H#���#9Ux��k��[�m�"h�%^ta�T:!�
��ІN��.��A�d�b�S��qEN}b��T��W��E�"���������f�a3�4�U�\(�/���� g=�.���)��CIo�v���Q�?�j���Z�t}�ҋ�p����:�MO��Ԡ���,���z�y����A��m,�C�P�?�q5����L�r���,*��l�;����3!/KRU��P;c����H�H�OS�j�G`����5��P���4{�rKa�!���+̱�\���S��pc���F��݄g+h~��)��r�����@n�dS�U.���+��Zv9z�<�[�'Ŏ�k�$�%�%Q[<G+�2���M�b�l�B�>��n�y6�#�(���Bg����׷�ǟ��m	�9Y_�v�#�+N���'Ƒup;��<Pǡ2�iЋ�����6�c�\�O�[�<�� D�[�:R�Ǣ�'XK�S������̯}���m�%��E}��h�xޣQ�E�w�̥?���'-Zׁ�XkNh�"cу�m�����Q22O����)^^��<����<�
Fɐ�){�g��)9Ɋ3�d���'�R���9j��V�y��ҿ�7,m�Y,`{7|�;M���%�1��LY��P�<�������@�������R-N+��D�qIJg���!�,,��a������D���+A�x��F'*}��&��pU�F����g�ILիU(�H���S�w�KD�bn	��}�}��t������W@�Qd��I�h>�c� ���z�צ/�/"��R���^ŉL��fݙ�_w���w���S{�G�~7���r!��Q;L��ZP��`��1H��S�Q,{xx	����Ή�WO����R7�k�U����QD�1�Ό�3��jM,U#��`�g�e���)`(�C���P��?F����/�`B��Oa�e!»���Vy��~mD	�ܿ�|\��5ga]>E%���"��خE"-yyAĪUW�95D�C;�X�����m(�^i��;�t ��#�����k�5�Ey��u�����N�*�熕�/�VAdW��T4v�.�<3R�}��bO���1w���?Ɩ��T�L)ĩl��?D?�ҹ�W&�u��G!���'(�{ 4c���E���%���.4�(JSm�3e�^:yT`|x/��B�>��,�t�Jq�%�qr��A���/4�HRN��Ί��w:p��'�˷34��>,'2��q�B�'�ri�v��B>�k����2(Ahb�I��Z
9�-��I|:$�a�^�^RB������������i3���k�����Ԓ��B1��X�}�%Z����'z�_�x64mhOm~(�� '��U�B3��H��.�6��K]v�(��`ჸ�<D������Ö \��j.o�ShL�v5��SԲ��z�өY߫�%��?�'�����"��@�_���B��
�k�7�S�b#5�	�9��K��b�3��j�BM0� ��@��b"u*C���o�˸�V��v�$���,ް6b�?Ph��lL��5�V��am�!7��!A{؂�ߢ3�"=4�Ct��B�b՜H�+O�X s�ڼ�R�O�Ū��������2�p��>�N�hqQ���hy�ro���(�i��[�p-�ݥ�d�ri�x,T)�!�-�C���$����|��P�I���m\�`R�`r� �]��7���4�N����Ձ�ݱQ�A�������?���=ׯ 4#�&����,�;wM�n5��D��t~���y���Y�)w���zځ�
/��<ǔ��g�[c�)�d?	�#/ "Tq��Fd�U۹��P�������>)��` cװm�=zf4[y��aɝK�.� v��i�_b�l=L��DVG'����� �k��:Yƺd���|5��AZ_�)�f{<ܒ'���YO7$C��l �������:�/��i#K2�J�p'8�>��FM�tp ������k�o�o�?��ؐw��dA;x�ᩫ�Xppw����/�-P��BB��|0�γ���N)��4)��ϴ�6XIT��G��&��5$��!/��8#�=+��Z3��
�L�Vk���^r�p�C$���F�nw{e��Mkif�jL��ǋ�+�l�m���wz�G���>�8�j��" ���N(,��
�������A2��'�3B�����%+�
z�l)٧f�X�ֵM�c^���e�����9�
uc�=�������`�#�u�M��-�!L�&b۲+#{?-d��n.�b� ��̓� S0�"�H�����,���B��3;�g��;u�M�S���&�IY ���!�{�}S,FT��~�M��-��RI��a-�$�o���)Rb���ыǝ��n~�r���@&]���W�O'׾b���Tg�B0�����-d������,}�N-zn�/�Li9���Bȗy�6Ń���������l~E��%��B���MPL���sgx��]��c�瑲9E�El�L#�~�W��|��>���q��Y�R���ܬ�H����].�>_�&U��xz���W숟!?]����6� Ĩ�9, �1o�\�#�`9��a�u��X�4�	�0\��M�/��c��J�x���/:���>���a�u({�E�6�f��}��&0�ٶ�_Q+���1���%\�4sk����y%l����	ؒ?_�C^�o��{9�$rl����ԯ�x� �)��d��׳���#��`sO�ׁ�==v��� d�Ic��՚\�ӭ�	��W�p�Wh7;1(�B�od.>s�ak���2+���l��@Hl���������W��jz�}�0P~�*��=�.X�:����2�
�c�t8Z�Ê��v{J�I��X9終�L+�H߇ .rCIב�2�YzH�ґ ࿇�x�$���W�X��GH6�]�+T��$���8�Z
�����=���*	P�P�2!c�k0U�U�4С��FQ�-��%s�������]w xV��Mf}�@@�]�,`
�DG�U�=��^g�?�q�$D$�g��Z���F�z��t��i�s?���OY���������]�X�"��3��AR��#��y���՗��WO�o�%N�w2%c5��ͭ�����Kf�b(e�ܱ��Q�H=|�PY�߼\@.!�&��4�I��l[��X�\�D׵"��$P�V"�mp��uT�z�AvC�sT:�ۡJ�b����FSHP� �̮��ؓ,.h��I [~c�8��������U�Z��(�V�ױ�N(u9W��DKqӲ"��6��$d�;�VV��a�~[�^Ԡ؋Lh��#�����1���Ҝ�>�)l)3	��C�̋\�c�������N�f���܃N�Xn��T� O 	A^�p����N�q1�,�r��pBiɦ�R.��D�xC|KR��/S�w{�5ܓ^�%
 ��u��GM�99�ۨ|l�"UU����a^!.`U.�v�
Bؾ���F*�al�+��$�^�5�cLh
~��V�'~X��sRUa�-٣ݬ�h#�,mMED�i���%��:twʲ��]�WQ��f��C�� �"�H���~
�d��9��M�k�\eȲ ����6�	���A�y�=�] Ξ=�i"��=�����]M�"0:�k$���!�,�C$��$	)����e�ކ�%�iT�d�6�ϟ��z����۴�$��E���tNt��v��i?R��ޡ����x~m�Q�Om��$QĠ�C�'ZN�|����T3�|00O83RGcL�}���,���H&8Â^��'�)���~�<jyy�/���zP�s�����B<+�����@t�(ʷ��65�F ����ҷ��Hĩ�U�+}9*�N��Nj`X��,������&��f��Y���U!I5� � yvx_�*���}W�������TЮ!��m�1;^�B9"�ٷ]\�6�Yp���:~�I��\���E���o�ƈ�b�2�=!�;��5E���c��ͲY���A���-D	��>���WQ��M�ny��9?Gz!}���UE�	�"���@�b�����p��7t8hp ����z�Ĝ� �T��k�Bn�M.��K!qg�Ǳ<¹1c'����]�߽ǎ,��}��t�B���!�;H�(�@�,�֞:��)C�Ed�u[��`q����K}Ǎ��FJp����Kh5+���B�=��٦�G`{�a���c�4{�M���GQF���>z��묐8�Ws.(�hpX�����6+���=;_��"�΁��v�;��Y�m�r�5(T-���J"��C
�pj�x9*����m�����޳�kIR�5�~4&@]�ӰN�1��U@h�����Q>ʧ:�zq���	\�4�Ҭ���{t���<�'�39-��
�t_"�"�����������e�3���R�i������E�-Wu��5(�Rn�S�����j�&�lW�fě��`W�H��m�}���1!2�ey2�PC��ú�X9'"M�U!�f#�8��`J��`��&z�������lw�ԋE��E#���s3.f���(�,}0�����2���l�ao�թQ��չ�e{��ZL�U	n�
tQ5��>�Q%��ʷ������L�Y_�E�$���[�]]�Q����Z�׏��dt�H�'���)楂�6@`���9��b��h���Z꫌Ӱ]^X���!�t��=�(��,�����#�u�f�k ���X��τA��\�)a�`Mp.��7#�RVOS��P a���;^r:���:,Bא����T���.��!��f�>�U��D��,�%�JW�m�B?�g�[R����;�>�/�+$i���cE40},Pg��-����S@�wS��$�ּUdHbr����?B��#�x\�8�_-i��X?c*t��o��
E��E�t�m�e����cE��)3XOJO�I=��H|ȯ�����F� 6�~�&��G~�wA��R�x�?�"T��V"�
 %�gS5اF=M(fn��\����� ���X��3���d!�߆�_��ʘ�7neu�G�e��z'6���B��+�����rJ\W�y�g����w+
E��f�G�k�9Ѱ�B�~�� ��~�Å�w������J��.�];�]AL��F�����S��	�����	IWz�X�����A�/1�9������je��VY�WdBO��s�5�8U�#Qnh���*|�Ҥ�2_�9��,dW]���L��n��h��R�
�v�0م>�Ō����3o���w��txE	�EBR
���ZX��[ħ*w�mPP?x��G���2��
Ts��O�V���7pM�ً�g7�TR�����"?뺝�d/Ф�� vɈ�����5O	��;&��h�~d:�x"DL;�h⭲$V9j�pש��0;�g�5pq�νM���!Ӝ��0DM�/Z�?�����t��p��#��1�/w��ܿ�n7�`J��U��F4��=K��W;�Q��"�����B�2-�zC�,36t3�+�Ioo�c�������Ba]�s�.5|�(��ȜN���M�:a�dR<c�$E\��Ձ��