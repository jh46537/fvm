��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&l�d\�vW�muk9%��˧�*0D�	0K�#��uЀR��S񟼶D�NaLK��ܔ��I�g�
���S!ی�ہT�������a@|��z�M�=����D�F3�g�;&"��rN���p�����Xݭ��8�~�0����i��;ݏ+��ↂ0�?�ceR
k�&��;T/�h��HKIw�|��&3.��Ů��p�!Q���i(�+��gX]����\G��/"�TDV
x; ��*���1$���'�os�G́�C2�:>�r��]�#A��]F�~?:6�,Ӱ������4;Y-�����|��U]�Ԝ���6&F,O���*Tkt�Zzڠ6]�ޢ5m�IS��Z䝤����VX��@)���t�I��Ml�k�{F^��-���2#��q릍@�BF(S��:�����jm�â.]"�	�i�,��Z��GU�՗��5�P�N���Lh�����	"���>�֞=]Kd����;�'��D�Yj���I��Kv���R�]���}
�jD�Kh-��W��M�� 	����eD��p���.��8�O���lD�Wa2]8)�b�;p![��5E���I6�����>FN�,5��y��zo�����f�_p)���P�Ey������0~$��^F<)أl�Ϥ��uvLi�9���~)��:��2�ӾG×)c�PB�7A���n]ue�q!L{��:�e��:!^���~���m��R.J�N��m�u�}�&�+τ�J6�����w���O~؀���.`R��BϷ|���}�����jx�n��筜�w�^�O"eT�� *}�j{J
T=9�H�i<��&I�T&Oũ)C���l�ׇ���blg{��әUaˢ���1��w���.���6�o�"�
�i�q.����r'X���b�"n1š	̿0c&!�H�k5~�vrOK�i�������m==;ƅYä�mZ�����ZB�:q-bF�]]jYi%�ꁰV-<]�x�(�GW�#�gѣ��)��c���d����ە(ai4��G>����jI��$g�ߣݒ���7R����ˑ͜x��5���.CU�Ǵ���n��$;1u߳��33�R+�@�S� ����(��[$��P�p�!t6]���')l�����؋�����w�����*��8�~`���F��b"��/� �N�����܋�+h��a�Ü��^;����|�קY�U���ҞT��T2ƫf��`�����y����89K6��H5�P��m�-�cw�=9�E�<��G�υ�ףC�)� �)���xo��bܙ��C��x�(o��j��/�y� ��h��!�EŁ�?�:��L2����K��<�.�n;f���5�`2=�I�@��ﬢlSYFy���} ��`0��k�7���`4AP��o��D����lt������˴�t�+sh }"}݁�]�����a_@�w����/��[�T�(0�Ӟ�ǁ�N��w~���9�	Z��Jt�V��@�b�W0Ifz�	�
L��2Y 7\�)�ú�ɲ�����ޞ!�s̮��;&��o�'Hى������z���)3j`f7pB�E5.Z3���"�r*z������{R0�f�vA�ې��Y��k1_�We�(t5濱�n\wQ�j���N��R�y��r��m:".+a��4��˻uI�#L3�3�L���@��џ���9�Z��ޕw�"P`g��ȹC�[2��n�� ��}o� �K��*��t8�\�������7*�[�9kn��&S/�4��M��1o*�@�{?�l���9�kY����I6/�S2|�����-Es��yr���Hf->��U��Trl��U0���O�F���7�t;]���y�G�ݓ�1��a��ϖ�9�]D>��ǥ��}ӀW��J���܄���<6m��"�A��?�mM^F`G�\}n���8;6է]�4Tz��UҨ7� x�k���
�pao^Kf�%P�>s�)�><�� ݏ�Ġ�+�M"��P~��g?�)x��OD�#�M�\�$������������+A�g�G���Rm����2 ��5��5/]��d���sY�;3����V���"����Q����b�J�h;L@���{T=J�7BFI,��]Y�uY9�~h�ЄP�3�A��l]v
r�83������pX����8�5��\���O"7�b�����?���������}����<�%��^~`g|��\,>Y�*j��y�����3�%!��}��ϚgK� ��ڞ���!��O�`���5�o��&�p@IQ�y�d@¡���ke���Q��A��u��n���{}�^���_�T���'y�,-�/b����Y�������`b��PP����V�^bW����P�nԦkF�����\�*���0�!TAL�����E�i��+,Ȇ�k�p��	��8vF¥�����7��J��H���y�b�S>�x}궊+vb�@'c�f]S'B���"�I4�=���cG���8�bE��^��(�~�3\�%��1����"Ab��,I�Ǖ+D"$+Y׀�f��֨����9�C-��nb��5d�|P���Q��� �������4���\���tƢЏ��-d2�GFE �$�^P�.4B��qB����3ށQ��(0���ɟ�{y~P̓��������ǈ���lQ�ؿ�C%�������qG��Z�<+��h]�<B�㑪�˦O*`����G\�W�xOF��1��AN�W��}��E�PY��-���Z�T��O�O�ixr-Ӓ�+��h[�C�c5ɐ��l��@�Y��Wβ�7�*�1*�F|k� �d_*n�ߜx���o��Q���c�ډ�Djw'R�:��D9�4 �伬�ϴ��U!sV���V��"|���E$x�L��`]����y0�Vc�����[���z$����eȦ�8���^q����d����wF�bK'd���L�dTt�z��G���5���H��ج3>ZR%Yg�Me�$ӷ+7u��@�][�n�H��ݑ����Hs]�{��l���e�5O l���.�OoW�_���&<S�G�潪�����?E�S�c3�����0����:[t(�R {��� �Y�Џ��V�	��B��B�ւ�[#�A��K̓0����%v�����5�z@�#��
���l��	�^=�v�����C����(N��& �j-:�}c�b�2>oa�i���֝�ϊo�6���'��k|�sPA�!|�~����-�F���PQwn4�'�@�5(�V��aw�����з�7B.c��d޺'30�&>̫7\�gl�I��s1:!/7ɊDܴrx��������h�l8�"��_�"�\�6~q\ Z�#K�1&�OG���_�*c����#Uo�ѻ���aJ~�Ѣ�l��J]*���բ���(���3��H��O����1J7��o}ZR�g�Y���jP.�G�d�$�5QY@I�s3;�y��MS�<>:�ä�ܑ���T�5*/0Ms���ͅ�YG7�`� ���g}�_�M@�6@\�$�T�	���r~��2;�"�X�}�1��u�]Z9�Ը���p�p�vRBI������� mM8��~��k�]�>�(�l'�C�ר�#���S�ޡ@���`��5�r�Z�̌"3lD��d9�ŝ�{G 鷫9������>�~�X5WJ�Dd���ձxrb
��	n%j��<���+��ޭ�6�-��Z�<S�<��s��+�,9���$�k����9ok�7[��+�j0(c�f�t����j//~ĵJ1j��>����U��V[�y� � ae��M�K]�
�w�S�{M��E?����w`n����m&k�I���e=5�*X��m�@C:��f�զ�Șt��:�� v�$�V�Aw��n���Ҟk9׾Ð�b�c[����!z�X͏�t,��K'�M��Χ��~~{�)v�A�L� k�� ��U�Q�QK��0��-G!�=�/������e���#uu�$ݟt#��+H=���9R��:��=��)���9*�-3����[@���&��2lC,I�ge�N�V��hx���W�)���ҧ�P3,�d�9��Pt '�&���ZS]v|O%�ZՕ��� 8�:��Mv}WQF\<��k������@R�)�FA����oW�E��k��>:�c}X(��a>�Mk����B�����eN�t��d&�dx��P-���T��Qr�6��Ag3~dJ������Ine�K�G�����`bC�"�oV�R�7	�$?j��YЦ�Q��U���Q-�<�{j �G���d!�&��%�5�+�"Q�L:^>�W��\�$�F������Рh�!r��� A�,O텨����1��:�S�w������4��n�>�B8v��x<�&�
P��ǘ�)���$������k<g��3I�l.\�@r��B�����.O�T�yJ�
����c;��T�Jr#U!�.�ԅ !�&]U�<wc�"��$a�,<�J�� ��8��WIP�z���K��1]�xY�g�|;�J�íJ�O+5 .�����MF�����W�|_s�Gr��T�|��=����gZ#���BG��TfK=�����`��z�sb �7n�/����%}��K���~77��6p��/���*U�9�)�$0��� �~#tzj��`�6]���;>�z�.��NP"�O(؛���2P��l���Ei�<i3���$5�R��;6~�z��j_����!��w\ݩ�0�Z�&s���.�LJ�����z�Jj�{:���>�A�;5��ˋh�,�9��2XNt%I.��Ic�s�h(�� � ���{�g~[#�)}�`'D��P��������(��络�5��p,+����>/���牶�F
8W3.�H�d�~j��.ECDj��[=�Vt��؛?�f#$�%��,�A�`�b8Y���Z�#9v;�J��sp�\�K�|rP��d��⇚~�,t��p�j�/7��U,?�#���5a��`)���%�&�r��Qj%��D�k����xPe/���Ф�m/����w �p݁*��!�"�̤���2e�z��BI~v��T^J�R+w��������RLo�R�l$]h�)��iOr�)��H��KὀgF����T�
�:R^�4b����$�@!��|Ĺ���,��Ǡ	�)�UgYf/�*�`�*zD����&@VZ�Ӵ��o'�2w�c�����0�O�����(y��J�U�GM���rG��m�_�A ��If��	W�D(L~�L8�5h��*"*S¤�g�c����{����|�=A�)/|'I�e~%�C�)j<� 1m'��.@�lR��ᒯ�o�o�h�wj)��8��)�TIJ�4H��t�bHq��Y*����'Y/�G���A���)mzzFO�m@��缌�f��HK��be��rH��dv��Mɵ�FA��ߑ�> �ȷ�C�(����i]��s�,��=�ܻ&���ט�QЩk��4�~/�o3Р�$�ゑ,
�ow�@�⁧�K,:u@�6S���U��퀃�+W`��8����E?�'~Di��[�Nΐ#y]�0,B�%����)�b�jXc'�P�:�ȩ2���դ���]��/1�z����������Se��j�����\�>v��c��&��Vm�䞽���ԓ���)�7�(�_��n�"�;���������\��>�@�������/��oG����E���	�
�$Bȁ�d�n�_͓�#�$�z�S�w��f��Xǎ�����#�t�O��L@eu&^����:�lQ� ���r,<�"�V���~��1ҽu;��eƖ�x�D{h55�E�V����dȢ�n|8�D���p�A����9��s����m(>�r/@>������ɬ�^�ˬ�*(��J)MC����s^Yt����I���YJ�B�(��Ɠ�m�w�8�eJ������VV����ʸD-� ����/n2���V�>�R��shaf����8�24=�);�oz4�T�0�r�a����]�v��D��
1�E�U@Q�c���k�z!�� Cuf��nNga"!�3�ɝ�*�ֺ@L՘$v_�zƙ��׵S}����@�<gG[�^����(��EǰLQ?r���B]A=�����EI@���ѭ�p��w�L��Z�e����@���v���kk��$3��	au�c�H/h$���p�Tì
k�	�$��1e����M��#�o�b��F�3;D�R�җY�^���X�#cLϓ���LÑ�@;ZQP!���<Y{��jS͕�P�`��s�AT�`vO=ܥ[�"&4�8��S��	�fOp_�\զ�x�K)��'�4H�G�} \�,���QF1�� ���(#[-,�C������g�.�ס(�7��kŶ��$#��,��Q@���WZ���WTR�h`_�����>�eO��ǵ�k'b��&�;'G�)�~�c�F��+؂���t�- iG*�h���p��������(�I��ϟ�W����G\LS���a��i�[ܫ'�D�8jP�B�$)����׀~p��|�g��-�o��gc�n��	59����K�����Ѻ�"NK'X��]Fy���$.�>���j�6�BM@�{"-�ZU�AF�W��)�X�����fL�f����&���
JVt�aB�hf�b�K1��oK$�+��q�a$�}����/����agR��{s�bu���¥P��}�C�Ugp�����ר�� a�:$��F�n=ЎD�Tr�PEA��^<�0L���Ʉ�X1��R8S������� �x^�u�@�G0xϦ��؊o�\��W���m^j"�,2���t蝳��-j��_4����d�V��,��Ƣ�KIK$ԕ����دy3�@Ƒ�����>;�*5I�oo����u6O/��$ ���P!���6+��8w��vǵ6�"�a9���4�C;���`^:���������`T��3y]!��>U8�]�?�ˌ7VSw".�o�<0��i���D��=�R"�V|�q'/>w`{1�%g������9zu���Zpdh�=iڗ�m���yD4��6���;�b+{�&حWpxiU�Qa����e��؅��=]д�v ��eN��\8��S_�߻�	�뻄#�$�(趓���lʹ.F֔�]ߢ�������/��Qч�i�6����<I'����o�-U&k��P�������|�&۲| ���I@�&��7%?�Q���T"����7��V�M�D0
��Mծ��O���w+�,mk��wZ�[�8f�?���嫋�c�_��%�� �ا���G�>��]x�q1vRx5���A�E�����_p`b��
kcՊ�j���6-z�س���%�D����%���c�Y�,�W��?U���i*�,4	�-r���d��j�lc^�j)�l-�����+Ч��2�檪�u���\��`�s#d.�ɻC�X,���5��D��3ZQfM:|��V]���ܹV���Z+؉�#@~�z�'�Գ*@�SSMOǤ�D�]�6�ղ�ܙ(�����I;'A!����Kvt�Z~�W3ԅ�*ĭ������D)��k�Ǡ�ߤ�V��| ͪ*�J����3�ѹ�w爓/��\R������q�Z[P�}�o3�!�;�6؞Z�]�a�?�Ce�kBa_)�w��C�$G�����^�
�kp�2�I1���j�[\po
��ϛ�8�8ezlb�Ҿe��#m��B!�Urc�X�I���%F���L�e�(�;�3-��4Z<����^�� ��Y��d}���I|���ΕV��6K�X�U>2h2wDWL��Y�����ޞƎ^ t��-�����6��V^K��ǙH�\�QZ�_��z/0D��Iu#�����6�#Z��Q�����9�sZ�
dÄHP)�����C�F��#�@��a��ZN<��o��~��Gnk��з�%��Qs2�W<Z�F���w-M��*))��_,��r'���x��&?⽞ZG�h�Q���|�J���s&�,�/�R}�	9<�wݰ.��;�{Vv#v�������������T��>���U��x�=9��F�豊��5W���
ǹ�u$���c<=���H��L�D�jw`Th?�I�T��ݭ<�� M|��v[F��T�� T�7�Ę#���:�~p+Vi�O�%��O�/J���4P�aIk�Vtۤ����议���O�?e���&�Eڵ!4�%w,i����`1ز<��3:�0����� z��B���o�!GzK�WαUG��yp$��cAp��|�6>�xQ�_�u��A= �S�=�PZ>��*q�3�z��q��f�M�����[�M�صNS,�+f&�1?�ý�����uo0���z�ז�I�N�#�%z��S#z����B-㊈�rc���_�Lg�9�w���>��"!m��Q���x�؝�t!�s�*NI��WI��Q��^Ĵ����B�?�8F�e_�C�{Bz�EK��d� f][�&m�)3����Hk�۔���:��X�[�����"�A\�|���m,�RR�?�Pt1�8԰āk>�dA�Um�38��t3�������Wůx����v7C��b~"�-3�`�SM߾VZm~=��� 	��bI�������4J�bSt���L%�S��� ��� 5xw�o:�����;S�?[e�DYq&=���1~�[����I�R�c:B6�b��
#�q=��/ޫcj��f�$�ui�'m�P<Ɩ� �����V9�?��I�*8K'
Lӆ���D��U��x��MJN
N ���%Oh��o�'5�-O��~B�o�;b�T2P�Xm@Tу��hW��kr�X^h�&2�Ij���fD���LR$�����������D�JzdS}�2�*�
��bDe6����+�SMP}I��W��M+�8�&[�F��o,r�4�jm={�K������gD`�1d�Z�A��>݇R�,��Ȭ�Ț�o~�7M�I�2*@�F�9^�����7.s��O"��c�6����X�Lb�Oն�Ƨ@7C�
0^V����l�p�w�E�:$��A3����o���N�yl�5H�!F��D�v��j?��5�yZ�"D�������q��a��˨u2Ǉ�t�� � �t	��R@X�[��\���ܶ�ɢZ+#��u(uw��Ҍ5��:E��� f�yYM�`Om{r����\��<�ԌI�w�TK|ED����6�<sAxea�5�E8�,��{ɿ�ź�"�����:��ns�0z:C�Q�y�0���M���*� �9]�2���6�=^�0'G�[���DH�kp.Ӧ�+�8��6��@���g݊Í��[x�/~ �����O)�x��ʹK�e?f��\!jt�����sH�Lr�H734�-���6l��rLߜ0����D��^�,� i璍�����Q����]�m�RRC�2e�~ѷۢ/����@w��:=�<����ӊ��h�ū��D��a<57�,�z�U�5���l��&��HW+x���I�� ��n�s�Ň��� �5́B��̜��ig,�z��>~/�:T'���raJ
��`��`�M�U��s��L(���
��C
bPG L����*������ɂFә����C��0��]�B5�{�y�(g��P>��u:U+W���H�[Ǝ��.aI�,4�U�e��xZE�{�6g��OrD�9�ه	��h
�G�]�2]3I�b��z�3��~qx��J�HE�;9���˰ϡ��I��(7�K�s���(Mb�ͷw�ӈ2��Ū�U�Y���х�����3�,�w�[z���#��w��צ�,��a�Aqpj�_q��3��]��V){ui���"Hp�����1
��x�P��4�����=�����N���!�*���A^M'�T�Ɖ�H!5�zJ��N���W�Ձ���n=R���`-ǎR?^�D��k��T��K����:=�|iH�kͨ3��EU�G:]�6�j�����0�5���0��鳢4 P���6�P*��9��5tV�뻑��'n��
,8X��&���D�$d�+�I�ݙ�"_<��>������_��&�Bt���Ҥ8;�~C7' ���M�/'<�Bvk�: Q�ǫ�}d}�p-Oi`��vMf��+��r9���}i�e͔��t��)��-�QB��7��8'��a��A�˯jK��?LS�2�����&FycM���{eQ�x�P���c�t'���F�D�x���Q�O=`�Qs���+�.3�&��S2��΄��
�i�˯�[1K�nN�n qN}@z�ʠ�����0��:���(|���G�
x�ZG��Fc�Q[��j��ɣ��0�Ko��A�6	�����1�րD���R{�"ni�s�kp���t]s�$��!JBc:�?%��2Y���O=M��+yYҷ3o2��և��S�:��fy���v�L�|f�o��'�H���K8�V��{Б5ʩ$"�P��8}6�q�,r������lȭ�!�N!&ZG90ͱT��yN6+ܩj�pq*'Zz��X'?)��ꋿ�ԯ��Q��I����zN+��g��5�1FU����mb�jH�>�a���x=+�?�X��Ȗ�ǥ*��7��@�l���jj�
�����0��H�ٹ�_����1����'�0�������!B]M�Yd[���	�A|��jiDbD����VI�Rטu� ��(�x]j�h��ŉ���{*S~%�X�"�Dn�q+(Pi��'F���X�@��Hh��������l-�0�u"
)H���5��d��sG�0�a��D�wO�I���	�s<cJG!V|�C�Kb���v�N�&�̢��-��?̌C-�??7$l���gke1�!�&@���`���e-k��1�}�ޏ}��`i�1m�C�%zL���,X�#�{=2�O9���:���z�Eه�<o�b_�?��݊~�������e���'���)8�<N-_@��sz�x@�MB�}!��g�I(��h��9�����;��-u�qh�N���s+��x�H�X*��pr�>�Oԩ�QQ���E���<��
�=�^��A,�3�D���w�x�u^�pշ�8Ұl��~�Ҧq04o�ꭋGG�7ǺO�r��N�enm5��$����D|U�7�FBi���@ۊ��)���@���i+��X�]4��`�R�3��C���p.���'����4Fs+��w5���ۖ��C+l��`��]�3ِ��^���'ԛߠqL#��Gn�xA�F�5�_� G�|���s���K�9�&L�F���!�����nES4�P��6�Q���87f��*��5��kh쩛W�M���-@|2���y�ǹ��oH�B��u�qLE�S}  ��5��Ze��^�DpG�^�Ȅ"�m4�:,�v"�~�?h=��:([A���7��QD�G�1&�N��֪�5p�����܌�P�� р�~E�~tC��{�+�z?��M����a�[C(�(�� E�����'�������#�F��m�c��o���i��=]�Nw(Ủ*|���@���"ͺK7���D"ѐ�E���TL��Cԇ�o��g��^����}�5��X鱘�	�8��j_[p�??ڷ�^�.���P
0g6�;����*�f��^�Dq�U:ľ����?tA)8����@��p
w��]�M�%�*<x��	�[z�>��!��n,ݯ�A�<��^v���|j� ��Y��o����lN�6	3G�HLV��%~.xuZ��5ho����8��ba��D�����uBش
+l�����]�� �G�I?r��|J��L~�]�_���vHHLLjKg��T$w�k�AfXFB�y	qB%Q�O1�S-����7gP�\�B,y�@n4B���̀E���j�Lh� ӌh뭺l�I��F�?�����x?�o�sQ?�~Ҽ%�Mq�� �(Vnu�K{�����2�s�Yz����V��Z&�:�Pk���mڳkE}ӓ��5�V�y�T��Z�5�5���ǃ$�.f�\;�Y��[S�1h݊��w�*��		�}��x&a�kxC��x����Xߴ2���t�=�rdiVgɫ�Y�&HU6�6�"v��\��߳��)����P�w��b3 /2����u�2|��,��=!1�?�����0sk����b1*����0�޻�����@ ���� �g�>�T:������R�������%����#Š�gEדL��ĳK���v/pO�J�ƺ�Y`b#U�7��,ۜ�bI��b�Ap8��5w,�=�BGr��)Y���(�0&�Dyr��8��tT2��ظ��S?����G�nn�qf���UJ��6^�z0�b��AX��w��.~SB��{P��A0a�%�~GƐ85�(��Б~�ЇpD��=�d��,��gtJ'�Þk-7明�r��J6:��:c$�9��C��]/��k�ѱy���9�K��2��(����?����S&���6a�cRC��M��ݚ��o38�d ������"��'�޸M�?�x�-����jc����3�Hꈍ��?A�D)&�����W�W�|���L��9V`�s�+�a�?)�Nd����UJ`A&���w����v&b^ r����ٲIc��#�-8��_%��������@����gŝ9q�e^�t:��Ê��AK˨\��ߠ_2d�{�n78P�?H@��&�Hٵ��Ĩ��_`ߎ��"a^I�Zbgt�J@���f؝P_����j�FLZAM�]t�5/�yR-l6F5��y@l5d�[!�6G	(F�K�ĥ��G��2L!О�J�'s`g�b���hV��P�	@X�"�e{}}^Gu��d?(�!=<La��z����<� ��k�y^!c���}R�l���'��㢸EBg���ۆ����_�xXJ���)��]�v��)僁է�������(�5�n��0�c%���dd$
_D���8B�խ}�7�u���v���f�Ԫ���4�/������|���~�-8�"������ϝǩ�
�+��9�JĥD�!J<��)ﱳ��H�))��o���<\�kkz
ؿX�a�
�~��o�CF���L�ߵ���B��]WM�Q	�ZYPu�%w�%�x����O�)��;��*�FҞ:;�ye�T/���qt���Rya��G��$���+��P7k�� �_��T ��G�3�=D��{��]SyN�3���C��W��?MW+p�<�]tK�T]\N71�R��F�I�ktwaα�*o����dM�Ap#�ܞ��p����˳,����Z�.F}<8��:d�$�y��0�����js.�L�G����Q�q��`!�	��������������̛.�z!�3�R�8`���ڷO�j*�у��e��*�����[uX�?���;X��6��g�`gF�O���|����Ǜ1�v �`��.����g�_Sm�]�DS���>B� ��ܩ;�)�5פ����#~�� ��tx��Mh�E��� �^��t�Mu��!r������59tZ��sD��U�sS�09׮�����T��ǐii�M�ߘ�����ք័�(���a)��c�-%����r@��H#�7��2��\��Ăx^$d�r�������0^x�b$G� ��H�-�Ŋ?�co{ >_����c�q;>h)�n>��Ep�*-It�C1xDc~Y9x�_Y��x=��h��0[I�һ���\��Y���2����d�t�Y��!����0ĨP�60�1o���
�D�H�+>'�PF�M}��&���CE�~Y1��
ؠ�hʩ��s��x�/�D�7���Zª��������L����ח�E+�c�큦�2�0z�*3XB�������8�DV��R�M��PO�l�D^a���Aj���躒G)7�`�]�B���Ҙ��"]��O$"�,�R�vsz��
h�f����.��A�
>UȐ�є���?�r0�AG��eu�-V��Ū*Y�8M%��a�r�U�	�^��C<>y�iQ/�\���5�A+j�����H��V��D� t��pFa5��m��lG4{�Xd�n��	�8�����;�<��,4��.����kz�5͑�{��H���!ц�����!<]�o�r�1%qs�;G�����zv�1�5�ǎ����+=�_��-�}���*���1��/	3V�R��a͜�+�@tT3�AC	���˘����*$jv�� ۜ0��E陔��)�W��xo�j��V(�|�W�&N�R!B�o �?S ���y��M{e?�b��6��*����_U��M���T��\"�,�9@���8�^�
'7�,�L�����L�yU$7�"/~��sS)%J���S ���~k�0��k�"xRC��̫�gj{2��fF����$�7�Z��3`��(�0g%Q;n�0�6S]R�V?�Ol�E��\yUV�6A[ͨt-���)�T{ �-�W���B��0�#Kdw�#G��Й�<z������a+s��Ҙ���	�V���ܭ��2��p��^n���R�k;E�^ҟ�O�W���%Y���.+�VV�f��.K�v᝘��g[V*c�4��(�������a�
@����" �<�8|��<V��%��@���nG�����n�z��o����n,'u��b�֓���n)F���?�g��2���>��}�k���X\��̑�>�,H�n��^k��
���&����3�x���y�<�MJn(�<�c��uJ� �G��OH&/�h� .Oi��h=<�90��1	N�K{�+�و�B���o�ͫj����V��)�'<v �K�	�Nk���cZ�@�D�R�Q���a�J�� x�D��Zk�U �dE��|���_:,�H��G�4���,V�t�3�%�혚�4��,y~�ֳ@�$ˎ�chh	��c)b����`��
3u�I�|��"P�ԯ�&)�v����Xw���Ug;R^���?��&���bl�wQ��\ѯ�l9�������ބ���ed�ە�$>�2w ��L+4��*�%�v����l���H����Fe0����&�kU�L'%�=2+�(���s����>�����RP��7���nW�g��P����O[#�����pS��v��D�f~�\�Trrd᳦A��%~UҤ<Ր�
���j����SFTQ���[��8Yъ	p+��g���w����"����Xo�5�k�&�s�1��I�A�/jtL�i+�R�Q:'cSi �R�.�:L| �jS��<���b���X�W4&X{#�>kH�x8��
�v��2���:�i I}����(���l!����� L� ��/�Q�0�,f��&�U�Q8O�BG2���+�I���A���IԬb3�`��&���e�V��B����]�r��Z����e9�=��U�
�>�q�	
b�F3z�e���a��U0&8T�Zf����'C�P1ؿ���M(c�u¨)(8�9�7�$g�a-���M!�#��cv­��W��jR�S*�5�4`�j/��f�*Jk���:s��XPAoʉ;Mz��� �NRVM�J}�*4N3���w�iI��ƉV�GYr��㝸�
� :Ao��*ef��2��>���c֩qY��Y�i�KI�BT۸��;�Cyn Uu!���@l�W��X/��Ɩl�YEg;)1V�4���R�UW� p�X�r��&�>�C� 3�dl�) �:a����h'?��c����M�{����N��H()B��rx��'�mT�{�?%m�}v��uō�q�Tl���f(.�Z����Co�Z���p�a*�T�����;�CQ���[;�>=BW��5N���4G��������\����'_�\/mE}� J��f��/��1�^��:�E�!^��I��\��lIb�[T�髕m�t�;�خéܱ�ΰA�v��_����/����p���NG��uw�-�Z��L�o+�U�`���7��Ya�Zx�zJ"R�F�]�����.�̘�x_�%K:�Oÿ��yd56�C�k��D����zx��`��[c�=�G6v�jY呗�-�~�i��ր�EH�r�|�=Mg�O��P�Q�r3Ev�8c��砅ۯ1�P�h��Į�oҗ"���=�7�L���;��4E	��w\�<�ũ�6�f4y�
u�����r����[����!P�=��ٝ�S�!p��pu\��fl(���1O���M�
�-��������5h�B`"Ϭv�obZ�J)�pA�1!v��7J,�V�1�~�:0��� ����dTb�[�� Ъ8.*ҵ]�j0�,�������!!^nU"�p�}��b�]ӫhd[,�M�(_�kWH�жXk+�o��(�N͜�K�:,�.��Ug9��������A��,���㹷C�BF��Y����0��c_��ca'2$�_���u�f��!}B<L'���䑋h8S���'�� ���ہ�C�����ou�{��a��6��[ri������i�Sm���B :�d��0��5�)#o0���MZ^�s����n��6����;0ͿOL��t�AF�mAI�4�f�D����|����@W���Ǖ坵����BQtyte��y߅�i�-;K�&iz#K'�����%����t	�(��w2`4��	߶��{�1�!&As*/�b���V���+g�\�f��B�P�n�\���p���LWE��3=�ǽ�s�D�}��>�S��^l��T���*��c&n<rǛ�K�f+������w�CRn$���E��p���U���O���/v�7�»PL	��x��<ϗ�PFo�+vG�z�V����h��Yp*B�����W�V)������}d�(i�!Cyt���jĆsy�G���o ��L�p
t�|N/���]�?i'�m�:�B���W���F`����m�,�9���\����DQ:iJ�f\�D�niޕ3C�j������)R@p��^6��Rk�7�]��tY���k�J8jR�Y>$|d1���9�fh���o�SXs���C2r�N����~
죲�<�b����{+�� �
�������hf�9���/���a٨I��_�ʰ��V�����5K�]�s��Xw��P���]_��&qs=.�|߿����[������c`��<���!v����K�SC�3��ZB���葃��"�c+ys�\.���i��������8G�:!+"ӽʰh�!�O�YS���%$ԇ��@R�^���0��+���*+͢�A_����K��b�IB ^��"��`T$�eS�/_r 4��r�9�Ymާ���Mw�4I:~� �S,:`�ȷ@�E�f�k�"Z��P��9�H�n��:Y�i*�Y��X{Զm�D�t���`HmvH��Z�P���jP�q6ª�Ѫ�d�CU��$L�`f�Ku�цtCooiZ)/e��X�s5c5�t�s�uB|3W
��񁇷p��7>�������qN�wFM:B�uB���~9ܟ��`�+�$G�G?(��j�����T<���Q��~�2�3�bI>�@��0T���[��l��@&�wz2]�@�x�h=3��W��F^q���Β|��jL���R�l�1���8�7Ec�}�:11��e����(d$/��f7b�+J����>	�YFy&������U�rW�3�9���*���T��﹈n��r��X�'Z�]W$"��E'1�����t$�\�D�.���!�yֺ'�{t��GЋ^S����S�e����9����X&B������\K}�}h�,�$�2���&�@4�������g�r�Xx�ϋ�aJ���);�s�_z��S)��|�����bDkk�%;�,{��H3�_��Ѻ��u3��leV�?'�y|�$䌽�O=
L�B�p��ސ�'�Yړ\K:�7fe���F��XS�>�����6I�N�fɏ���v���:��RЅ�r���v/,3��EWT~��n�
���Fx�]�4�"e>�+�z4~y��U{���O*I�
�m��1���3��P&�{m���]�G���=��0���b@�d��҆�@3-�<�Ѣ��Ԡ�\x���/��;u]�#ft��Ӈ��1�H�jN�ɦ�2ZiK���1��	3�/��v�C
ri�cM$rn�PG�T�zم���<�Ζ0$X��^�Nk�����F��)��h_Ѱ��^�d	�����u'(z��Ώv����t'i�5N�1��@�����~���,�]�,'|��t�]s��HfS�`W��G�%���,ӂ�Z ؽ��\���$� ԯL���>�+jD�z$����#u����B�b�~cޕ�j���#�/��xjA�4�90��A��Q�@mO�1�󜿚���/��lM�V��Qd�h���[rd8e�M�+�b�-�7��k�W��;.��`$E@��:�V�׆2�÷�Z3��IX�&m>�S�*�g1��S�ԟ��:�2m*��>�;�Y���V�w�ge��k?O��?�wde>�?)�z�1���D�]E��O�?�`b9LV��p
&�����Tr����^h=d'�C	�o��3r���B6�f��K�H�!n�M�7���z��A`P>&��Z��e;��ܓ���v4��(�4 ��6�5� ����"S�,��t#y���G8��X4�cˮ����Z{]��U�V��ӄ�k�5Xs�{�t��f�Ӕz<�gpy���S�pB�մo��z�b�����	�t�Ξ�P����:Jמ0?V�<T,��څ���RPL��~5�_@�&SVY�h��I�e��=���"A��!L�ӌ��߱��-�d?�$�7U���m��zp����-FR��Z�Zs�����ҘR	Pæ����kco���UZ�n���|��=)��J�����\a7s6�[��,��\/^9i�����}�Չ����\�V���'=Be�q1� 2����-`�P�j��h-d�ԁ� ��E�z�n�?���4Ӎ|�7k��������*i�J�� ٭{��ҫ��o.h�(w�����S��4s�Е�àq(�=(X�Gى����gr
����'x�_1�����/b������  ��G3��z1b�P;h���w���eX�m�y���Lɱ��������7!�;;9�"'s��G�O.�����&�x���/æ���1�����ϯ��}l�o�qP�):&�1���љC%�;?�x��`���X��8V���[�8���h\燛*��~�Y������K�	��99�]�9ϭ�ة���xc6� 8���Q��]ǈ<u˾�����[>�����ٶ�s<ZM��TM;�5��d��b�d0k��
q��iU���x����<u\];Ү��I0~��{a��tvhvbq��,R���fo������E�����z4��ѫ��&E�2����2Wvm���"�@����zEAÍZ��n���9}u�T=0E�Eg�9��ܕ$�:��,�%��J[��*��)֐lҥI'3H��w=6�h.�
ߓ�\�i�Ǡ�VP%͚X�����@~�Fs/���M���5*gb.mݮ�#���^�*��֊ښ�YJlx(���Y�(��1ï��Ju���)z�|�����O���pZgp�a7Ϣ��H�H���W4U8������7�_1 K�km�a�+8����ɂh&��3��j������������c	�$�Q̊ڟ��&L�E\�	�=Y�e�-C�j1�	:ӷ=�󲨀#56o�	��Y~;QD"
��Mؒߋ��^�Б��&���$ȹ������a!�5Y�tP��D{��0{��u]H����s��$>����̻ViK9���QH}�N���2H�kL����(�3�7+*0� i	�D�-�j�1� �Q/�cf����Lq��y�꟠v�ǂ@7sZ,�s>���K˳ ��7Ybtl��@.�hT�H��[�<�
��� nb;ȟkl�70t}^��q�V�F��a�gi�XN��-�����Î�r�|�=�� �m������'��E�J���9$B'���z�Ӵ�%T�<�[���%��X�m����9"���F�'n�o�%���4�K��v���Gӻk�vxAߗG�d�����((�(ݸ���):�m!�N�c:ʡ�՗r�Y"Z��jg�-��]���<j�t~��ht���q�F�߈r�8Cr�%v�R��9����4��RJ\D�d��KT��7߻��k�eX��(��PÐI���M����H;�7x�%����7���tѫ"7g�T߻W�$�գ�R�2��G'8��k@ �,�!=`J1H�5��Z(���^	�6N�6��j��5��L�,�
���[�N�����y<V&5�^������)���QK�]ϑ(:o����`6(y���}{Q�3��D���lߩ�_�;i !�
&;�P{�ہv��A�˯?�i�!m�W#���P����j�,"kê��)L�G��6����vdP�������=a*�_����	8���8̋-�"�t�䫄v3ҩn�ז�t�O/�b�n��1&H$[�g��۲���**���v��x�����k�[K@�C�(9jU�Y��(���K��i�
�|�e�=�A�T��Wm�>��?��ntcѵ����G��ؿ"NZ��T��T�t��]��)�%����I,�)�&ۗ ��太Y���g�q]�ް�I�+��${�2��M�*8��3��J�7��������.��d(�eM�Pm�-�ų�j&{�$?6QH��\Ԑ2m��_�/���֑���mk�i�C����P=�ў9��5`cM8:��u��3�&� ��d	<=]A�B��ȟ�S�Y�<0���}G<�.^���])�h(�Y<8N�PmEо/=|V[�V5��W�X�e���m�G_���d�=���e,k�[<�3P�ȗʼ���r4�����f��j�Y�i�����uڱ1Y~���Cz����ܜ��|[�U��/uK�7��N�.v����,o"�T!|ʍ�/u
�I[9�S���zeN�t0C���'�Z;%4��G��1��9	oG�m�^`Vp���Jk_q�AwLt� �Lo������--�9��2�T#�:NS��M%}��[b��������"m�3
_�śK_'���:�\�f��,�An�#*��F|���~�m0��"�ۈ�.M�6��R��e�i���?�z`����Z<O���Di̖8`����Hfnn#�)@��� 7*vX�9��.�}��5^��|�n���g)t����3��I�D���C��Ks3½UgXt��' �1K ̭�+�9 >cBCg��f�3�G�{7u�u��S���ڌ,:?YGٰ�En�Ƿ�sk;Qw�)�O,���]�C����p"r�Y��r\�|2��xbZ�7���1ͬ'���$�u�0�f�+ ��
Nk/������1��&�����f���p��n�c�b�|�6Ԏ���S�����{2��k��F��r�k�:���@E[ ����}��l����T��3TdhV��j���w���>�9�n�Y���d�k	ᯀ:k`Bv�ܭ�c�2zx��a�������ۨ3��n�+r;�N�(���Y������]DVhm����@3��(�8���f��m-C�Om6yĮ��4X�6���G�r �A\�\��N��J0�Y�.���9��]��r%�}kW�
{��q�݌�Y�`&z�֧��ǭ���/����a`	W��C�;Ki�T���|No��.�!H��QH	W-`EHa�q�Kb2>���P{�H�۩��A.�п�?ln��N��͗Fޣ���D�|�ޔD �" �0X�-��_��}�ߌ"=`{��S��� B�#�(��8�'A5�ή ڝ���_��G�2�5� ��Fu�Zo�:�� d�W�ꨮ]*}����;
���.i��7`�S�S���Sƭ�K��<�+(�;zPV��6}o���yLGذK�c�qb�V���i ���١m!W/s+gi��ߙ�s`��
���m�����;c98��;�Tl�<O��A�5�:d�=d@��|P�q27"j9\��o���a����e	��l"�]H�۔�sȳ��/cx���0�����G���1Ai{��&��rV�H�R���uo;�np����pQ���T/yI8��*��}�!����.^�q~��;ؕ�l�'��D<��I�a󐀄�B���+c������O���0m6���8�s�G|���Sd�&�}�C_R:���L+
�9�/���ri���HO�����5v_rRg�=�ۊ��lO�r>bp�VQ�<Jx/P�g�y��%��.-#�He���%	�b����e��817�{܀���q��Vi{?�3H�Xw��mLX���s��F��y�T�Ҵ}}aC��r�����KL^p\���� �."�g�[oy�#�) �J���n�mZ���p��U�;��!�n91�=�q�#��Tl�{�NضC�ӊ�Qm��b����Y�� �~�-N?,��V'�}���A�ǀ�p���W� `��ص�+�'�xWj�i���".��.��3����<�ru �	,�8��qeS��H��B˖�g��Zj�2g�⿉�5��� ����G!m��De�|�2W�2��u��9	���+�M��&ͦ��hnH;�0�5&��;��d��j���Ћu�=���ͼwF58��?f�e�|l�a�vV�� �X�v8���+{մtƾ
��cu�_"�b��T@����+���ܶ��&�s*:7���}1f�,Ϧ�WD+��ƾ����_B�Vߔ�Y;�z�RR�ԚV���9Ctߕț�^v�o,���:þ'Z��/�$*O��j�L9*&N�d֭����~�;�	��5�5������n	*��UZ\XD�[�������f܁VD��n��5q�ma�~F��o��coWe���k�\�3Q68��'�%�" ��Y7�.�9�4��⭻��C�2��雿hjUH~��.���9�ܠ#�ߴѾ���
Y�TБrB~�
��%� >��Pu&5�'��BンAf\D�dÜ�����ỼM��º?'�%��K���/!�7\�q�>W�i7��k���g�cK���\���U!�է���]7<�����s�]84�I�uRlN���
�5*/�����Ѐ̰�a�w����\Ą�ׅn��)5:�����jɩ�Sy�xP�%/��@&1�l7���l�<?�.w���b��9�cgF;Yz�S@ ��p����&���<PRf��g�u����1U�$����5:����5�ZnV��'� Z���}�zd၅���m����Z�5~��o79��$%���j��uRӝl|;�UOj��6�h��p�<�w���$d��hZ�N��������{Q*�e�h�9�q$���?�<�����|���, c��b�a�����lv�@�ӂ=���Y�l�AP/�H'�݃-��_4[F֞�N������?*��E9gg��~����_�6G�X�5��">���e�E �n���vlnc�{��LJW�QO�9��~�	?z�]�����!�Qf�ig�h�.��]���~
4��P
��a�Y�?��,�|�鐔??k���뗊�3�;�����Z�����M�=#���9�v7���
q%
PY��܁�ޅ�C���̔Q��+��uc"���B h`ק�R��\B~�vA�x�  �8X�W�M�p�����9�O���g�Ӂb���!b׷�[�@4v�Oő�w�|Q���5���`���Fz:�E+���/���X��|eQ�D#�?����vEX�	s��΁ZA?D���	��Z�%$��+�iO
�[���ip_I:|2�-?���U�!�:��i�X�!7{e�I����4ﱳZp<���\+��e6K>,�* ���Mn��#��ZV�?��G��ݠ�l`L$�C��"�~����� ����1!�G����pt���8������^Oq����L�F��§:��*���MΝ�YjS�i7������F��w6�@"��6���_�����(���J���F������7���6呛*�X�B���]�h�֖��Vv>F
�in��ݿb�+2XO�	iii�B�+��v��㑐�f�(�Ϛ���3'K{�ȑKɑYj�ϣNî8��C���q^bv4رE��i�����X�Sʹ-$�Z�Z����&��Y����sFA��ڻ��.Qf�5	�	�Q�;	ː�s�%�k�~y��WP7V��_�	F��u����LW6�E��X�A�@��{Y����I.�<-RM�����U'	����;�,=���c�K�㑙@c]�1m!i�L����O�Y��sE� )T#"�Dņ
��8yit	c��_�k!J�nT&E�Ρڇ9+:���O��Aq[�i�w�CBf8�S�daI¥����e� Q~XG5d�<!R}I_򋂵n����-#\��aR�Kn���]��Tc��:_�K�EO�R#r�$��H����\�-C�u�����7c!
�h8MV�P�:";��XZ�Q{��ȺXg�O:��$a�7)^ƚ]�Y��0F�'�\��Ί+����'�f�/��g��|�l��
�k.ZQ��O����\�)�M�S�ӣ��M��;�T�i�"�]�N���J�P�]H����j@	��A �c��]�v�φ��y��ґUr�1���O��)��fb�&e^�6�6����`���ȴ���������������L��gr�Po�?���d�G�����m4���u�\~�ie�-P6����J@]S����։y�KW��j�k�":�1���h:��=�� ���x�d��(��U��=��Q[�ɏTXP#!�i��{?{�3�'^���\`������Ub�#O�V�z���?�y�"��h=&�Y`ק�چ��cء��l's��i�������]#�׹{�о�hc?$�(�������,�PF�l���P��c���k���������3���9Աi��tQ�ÿʔ_�g�[� ����r[�A��� p�T�2Q�pk[�
h"?��pp\��)��DM��7'��`��}M���8��s�%sR��_�V|!}Me:�`�v��å��5�V�E�׺�eC�^wu^����¥kPB��#���>�L����H���K�K��9%P�'⚎��x��_���w�x�W���� �=y;+��U]�4 �^�q���&k�T��Hv�'wFEH���. ��� s?`Hy�r�R���z��^ �S��v���Z�nywsW� l���P�$L���7W,�(�pM����4�0�3VZ�6X����Ӵ���e�K��4M=Nv�G���jGF$~K���^�p���~�EqFLev:uW�\�����a�a`��l_��i�P���o�d �u<E��*볆+u��
k]T��]�5BI��!�t�Йc���톯�����rg��ԭ��0�����04!'�U����	1넂�d4��������=)��b���؈��1�B�z�|X2�����w7�}x��y=⮘u>�6�O�2떏�������mx��/����ˉ}Ŧ���M~�\R����eXp0�9]	���0����@�(t%�֖�C�c%&1�LW��޹>�k�{��UOE��Z�By(�������Z���.f㍘R�eY�ԩh/�}e4q|�=3�:���K~��7?��sT�/��Y�*#J�Wu~y`���h����A;���u�D� J��n�nT�368z�u�z����_�
s)����L��$}0�o�H� ٧���$Xtj�����;�	O��� �j��%o�A8��P���}?v��G��*��<IR��#/�=we���D��c4��{�1s*�H2[�?��%�,{Sc���0O� ��������Z�Y�{�Kd�T81�7*�O�t��V/�:y����F|j���j 6��&��͔����QJ=S��K���P�zG��y'qO�k�[�����1�����G��+d�O����1�P�9��홈�<l���5h�����EL	R��$!��L�T�F���XG�f-�
@�cV�ۉ������v��5�dHּ�6�_ll�o�! �][?�V�Ra��éX���R�$��Afs�p@J�W}���h<0!��WӦ�������������
���(����Qc��8&p�(��Q��1�Y�|VS�33��;c��c0yHNS_+����/�%�/}1�PYߝI��Y���F�]B�W.�}7B��`��W��v�M�s�����w����_q$���,���NF����W���Us^@2:<Sս�aٟhP=���~�<���*Ȉ�=������+�3�ۆ����r�x��#��ᢁ`��3�iH���H�N����w.�g�*UA�������X��D��G������Z(��k�0QZ�Ξ�������A#l���S�s�IM}	�rn�UR�=Co��'��=��S)�a-���oN|(�zm�*����K�J]`�h��w��n� ���G�6���=+�	<�Y�l�56�=9b�@5�bR�S��O�&;C��<�o����S�#���iRe�[����JpIp!t>�p45~�� �L\C�����~�Rɜ������|uy�"d̈́���3�<
�+��L'�%�6-�{?\�jh|�;M´���E���s= �����4#?\���L��?K�^b�C;oh�����Te�Z�vP��;�8 �׿�0C�N��Z�i����.)�= O�	�d ���$2�j�4[� �Z�����ܲ�2���&Q����Ȱ� �pK(�@�b���[Ws��\2U?��[3.��=y�'�S_���%�>Kg�_a4�a�JY�:㏂tܼIǴ�@�^��Q���V�5��-tōV�d���*�>iG\��K�mi|m6clq6Ycv� &��`�7T?d�Tԩ����'�k/� �ia
�ۗăڹ���9}���+��k	�O(���t���=x�L�)4�'�bx�u����c�����{�Zs���m�}=y��zٟ�̈́�B
\h�9��{�O�$�)TV�g��������.kcח��~^��@v�YR� sPjױfi�cV��S�S܎����I��J�t=o-�(}�˺�(/��U�{ș�,�TΞ�DKx�&d��InBh�}�@��9�r�["��w�0mA�1��Ya��CTe;�;d*�����"}٠��f
��[�	N�J=-@�C�d�����C��f��C>H���x�<��6���Vbo;�h��JT�
���"�ICc1�[lT#ޥ?
#�U7��X�
/pL����Z���S��s"z�^��;#/��s^�$x�^������wdz���E:v���;U�*��="w���!��n,٢!1!�i�08ox�DZ"~s�#�Bv�I�AWO=��S����neV����=O��]�
�:F�{�˫ ��}H*;�Ib^/���/A����EX�uZ5��y���+)�,�k���l8�eW���F?���5l���n�M*�Df�!q�:3)�%�x�0��t�bw :G�[�\-�;�yń�I����rr5�<��@��[EإxuXi8�&��EN��'ebƑhuf��1`��h��=�G�8t��(|��^4��Y:"�o6����$5�����l�Riga������<NC�%J���fu���"1��/μ&6�a�pp�P���-x+\�>�+{l�^�M�u߳/Fo?E��x������@�cӆ%e��U�UL�v�-K�il�����OZ�y���J)��9��\�~
b���T�۩t.������D<C8 �D^��g���#�/dV�!��V�[�l��_iّ�%T��ZպrZ�iC�2v)O��
.U(��x���#�9i������/�x4�[1
�ݳtk�5A[�u|3��|�b�Ǭom���j��������q�6��
��ML�߼�6�q�N�1״C�T�&����A�|A��"1�c�$�- �{������m?a��k�>מ��jQ~*����g�#��c���ypH�Q����Zg>�KD]�0�?���g��x肈�D�l���5�O�����C�����y!��1�l��ȿ����P�U(�P%����j��%ze@#�a �Ɉ���ޑ�[ ��F_*�^�;K��v؄P��=��5<g�$��I����U�;yM��������9�T��A⇠B���R!�>�E�0��  |�Hx�q-��t�~��c��Ĕ^c>a�/��]獐�T �X����W�v�r���o�n�wi��GH}R�DjA��ي�[2���w�n�  ��6Hͱ�;Ƕ$�dE���``�����ͩ�����E���	�&|�������N�ǡ!�¾��z�����^+���ɍ?�b�!�b�G�SXi/&����ʪ�$8-�����gY0��j	H/`��@9%�s%�����H��H�U.���r�@�� �=K�/_��@��2n|{�T��ݏ����R��7eGSn?��;}*����q�OA��&��������b�,��;TRQ׋+��0G�1B�S�
�"�r�$�բK�Oz$q�'@g5������H"�i;��7�v$lKxhDze�H��܊'�T�<X7�'m�O��5�{�VQ,T�.���l����L���-�z���+! G�w�򜳐N�����Ǵe�P���ry�����{���vqh���9)���&��2��xQE�^�fl�#�mb8�X���±)(��%/V�k��sDEZ�ߣ@��C9F"e��h^[�J�P���p�Y���bX�Ct	�8c�N �o�Ħ�����G�YE�k�m�陏�wXl.��z��6�� ܔ�U���r����Yи\h/�q�)a̵h"?�#vv	�tō��9�S�E�x�����gz��,�s���0P��ё��yK�򅗹�������P�J���Ze��td�aH�����1ߎ6����g��6җ�.���:놄4�(G�8�"uMIbe�39����4 ,��얤c�K�>���7��w�$S�dfζ/�W�K_Z(E��:2t�b_e�%�iAF�ƈ[`T.ዶ4)�����	������T܅�+ԟ�<���ٞ5e8�F0%T�ڛ�ܝV�{����*���e?�099��c4��T@z�Ο9�@>Ĕ���'R��k�?����ۡ��B���k%�W��OHH�n�������"�t�<i�/�\/D1��"P�XSC#ױ1a-�"�_���!�8X�#;r�&cK���P7��e|����}�\�!��*z=�տy����x���FE�i)X''��"Ӟc���h���t�o;5��{Eٱ�J4��,i��IO�]�F~��g��[�,(}�w�>G�+�H����YM�|�J����|c����b�g�U����x��i/Љ�\����mM�\Ǘ��ڜ�=�M�_�QcWk�2u�����g�����E�E	i{��9��7��\+��y�h����v��4;+K��g������/�3�r�����,"�W��0I w�Rﵡ�E�؜�"�	���m�0r'�q �\f�Ӣ�b5E���=�����	9�EoX�B��5o'I�ї\Ԇ��}ut��^R������JU���D%�A�1��<��f";x�8���F,?i���}�݅�\C���>Θ��K�!�>�CC?.gw|z]�A�(P�����1�lS���JF�JI�a�Qm�����UC�Յ�'S�����P���~���V?�n����ה��>'�s�b��d�:?,����� �y�g�t�z�B�T��X��s_0��eI�nUns��W�,#����^t�	H��+���P� z�s>%�D��#�z.���ϲ�}��D��O/�!����a��O����ُ�|�6*�dǘ?�`S{B�a�"������S������?���.x*fpHlV��-"��q�ɱ	o�?O<'���^_�L�>�����������Љ��3J}�M��t<�1/ڴv�������c0���E2vLv���3{1��X��|���0�;#~�
	��Z8���ho�#t�����1�����i�s�C�mY�lK�����2f�6���zm��"��/.�.Ǆ�t��+�f���'(���LR+��0��s	K�lF���O�kZ�������Pܮ�Qy��#�gt���T�k��U��c~R��i�R$K��(&?��DOZ����"@`{�jP�f��t�����sE0T��~�=�QEOu��#��w��#����`��x���RQΜ�?z�:6�rJFS�D������A/Imd�;�@��یG��$����r�%^ܠXι��ٜَR�w��NƻGsӲ̋�~�E�zƯwHs�}�t�K��\����.����5|-�I�";U��sK��F�@�#�qb��,gg�6��uIw����rO�.$$j4����`㎳�BV��*a�wbk�2?�'L�&���Tb��X޵sf6��v�]!x�y�y���" U�E�����{�kP���P(Z���g���|�O�ʧ.�nZ_����X�&:#�q���o\�fO����=�5 ��A(�)��s�|3+��a���JӋ�S����>�U��	�c��f�^��W�bSg�T"��e�o	q��)�B#�?�F��CRX����Nկ�V0�SJ>�A���MH���ݽ��v�!ts���:�FR\),�mY��}DǴ���^�
vN�S�A#��'��ľ�-��z8����p�b�]��[0b|�q�P@7^��Nn�:���a{�L+���Ԉ���z�.I�����tl�*�b�n)�(�5�f O4~o-"�OI��K�k�p�wb�\��f[��赏
�)B�������]w�ތ�h1�����s53�Ǔ��IL?L��A�y�q����b8!`�Y�f<kZq�w���mfԕ�ٴ-ǱGN��� L�g3m�$9@G_o�l�0��3!�dʌ���(�99�ΈɍPj�~�Nm�m�T�&�8�A������'E��U�v�Z �VhU�(ٷ�:��X�8͙�����1�֬��<�)a-�������_>���z^T��ͭu��V(���|u�݌��&#���q��L�f?�#y�
���G~V�9eW�V�QC������W�0�|"��(�)��rW9e����,����Q����Y�C~_	%��塬�,&��p�7���j�������J2��c 	�OP~l�+#��t'�z��<��ݫ颽7�7+$�g�1�Umk;1����^=`�ݛ�m������h�8��&Y^[��@��:�]i�bz-� l���2e���c���?��@�^/2"���V� ��ko��t�n��b��<r�kwL)�k��K�)_m�p�Z�(4�i�5m�e��.sx