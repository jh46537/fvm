��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��U���S��1�$g�O�ȣi����|�璐�Z+�cc�n�-Z���"�����KB�]wdX��yԒ������!��Ǚ�]��6�rӌ"=	�I�{�܉o݄*U���Fm1���LEO48D�,>;vL�a�?�݌�uA�
��w���.\�f��H�.&��B$.��b����Ҽ���K�转��-%�N2����$1���=p�"��w�5�e!�f�b���<�X�� ̾^4�GX^w�*���RL`��{Ș���z���|`����=Q�c2	���D���S����6�E޳Hn�l|s���Q[x�MUH'}�G���ô�\�M�\��,&�U.��3�'��"����z.LՉ��ǵ�h#�"��Ԝ��KDSY��X^v���k���'[Ȇ_��	v�z�F�� Y6���qC6_��yϐ��bKj��s�!��m�fS�� 7�I�7�8���IF�HJA�o�����jz쪁��#<�o3i��$L>6.1F�#�	z�z��&ẟ\�a�5G0]�W�� W����F����y�E+crqH U(�t�i+����?���;�p��� R.�	C�
E��O���F��� ��c�� ���_��z�	!��t�xW_��L��e�A84��w>�=�-ݒ��v\�<�0����!~Z�O�i��$6�/Y�t�b�j!vr�  ~�m�z�=���H�̔����0��� �9��g�2�4+P�E���9 kHTZ�o�;�1�X��"��S���lO���	����Y��4��?�ٟ�ĉ
�2h-�:�&�jr
��@�1/r/����j������
�\L1��zqF����ǄX�2	{�2�V&��O��Mls���O�R�w�@����56��$�%S`Y�YA ��_�	��(=�u7���}���
�,=����F���ޱ��xL��z�Z>��<4�@{1�W�Jj�"l��ƻxW��!2gI_��.r9�z�I�w ��W��=wʒ� !ћ0��{�տWq����s�O�eQ��B���`�f���?�:Q�i���ǉ������U2A�� ؒ_�Q��ʽ��^�uݕ�}���9� �D#��C�j:��z�~��f4-�= 8&=:�u�W3�T��}�>Y� ���*M�6C�躓l�Mkk3 ������f�j���QPj���ĕ��B��kͳ� T���z��-1O�v�W��'�J�m����\�D)�T)Y��̶]�_`L
@�d��Ǳ�ֈ��7��l���^�@�s�[,3��VA�}�*��՞{�x���QR�U�#v�e�;\_kSUb�%2g�$�<aS!��3��M�ኙ���يi�˷��g��R({�����!�7;���d��NI�t�B�-a��Ѣ�[�\��b��#PIqē(z��Y��sΩa�y�|���uɺ-�y�c5.��-����[RH��J�yXqلi�Ŋ}�L3��E���$�W���P��ii_���?�x��>����h����=ϯ�r��~�~oF���v�z�h_}�|R�_����g&�H�s�z�՝��в��(������e1B�p��	�5m���>��!|ⶁs�<3������!�X�UJЭݳ}L���v��� �]�y8��70`��*,�w�O�4�)§��'���1⽩a9�)5�nR$Ȧ���J0�	e+u�l���*g:�27��E�����/�\5$��	b�e%�wA(9��h$2�	�P��<Nx�8����i�������̹���V�Z^]329O{�J
7A��s�p3 ���Af���H�[m3n���/z������~��W8�}ϝֲ��<a �{��~�W��(.�P2k?�o���IWQ�.^bi��d���o�6@'�]I�Q�[ ^��K��>5ۋX��(����B��
6B�� �<p��&���4���.�P�V�$�ә1I�y�z����=E�/�bg�y�,�FK�+̗ߋ���;c����D+�k(M�-���UKϷ�
q (6{�Ng������_�w�#A{�ax�d��F&s�F�[�`�j���H��EЋ��2�7A*��b*���.��gC'�%O�TCA�(����R͇qj�BƆ�/O}Z ��os�5���s�0��������-�Y��6�������2he;�p*��WɺĴ�r[������<�2��D��?�q�� �R�@ǝW2�m	}f� #qa��C�yB�ZL�y�\��P��*�&d�j������X�&}h&�?/y��:�M�G�i[Ax�d>`�`LVE�[\T�eD���(��D������1@�E�k]C�r'Q���N�k��e���wȓ�e�&7G��=ؚ_���}&>�.ǥ!�6_)�c"']xB5R	�8�9���[[�٘OH0eHx���p�֧4J����UʍC��e���/K{;=�Ҕ\-�Uҿ�9\����H�q��&�P��E�3�@H�^��O3R"��(��;�tT�Ѓ!~�����n�E��]���+iG�ϵ� H%Fd"ەe�I��3�d��%O�MH�!a"�
�~<����̧<3�K�F�4lXٻ�����&e5�H�X"���a�8WpF#��W�o}�S�A{���A9j�9W\	L�0+rp��㺶V�fd���Ф�\h��A`�4�~=����:�𾴋e!��sB깺H��D�(A�Ǆ%�{
:N��M
���lS���	�:�W����(cmn�R�e6�pbۊ�_%yX��$��/@��G�'�2���8/k�Kf4���iZ��=ؤ׭����[���)�Si���B� �x�����c�����)Vs�ΐ�U`kq��_��/r=4����i�ESMu5t|�Ξ��d��6N�����l(��/�י�c�p�V�TR �E�s#�k�n��h� �:��|�&L��Y�g��/�N��KUA��Q8�n)�P��Z�%lh�[������YVU�mp�^�Żk�W���kcB��h����V�"=�|�ݬ����;dM;k3����=0�cG	�W��Ѩ��7�zY���t�ī��fz��|�k�k?g�c^>O[>�N7]4�חҳ�����7"��2�����8ЈD��N�r�����˶�d���8��T��]��h&�C�'PN�v��iA�j�/����$t����b\�P�����+��M��.�2ѶD������@�R쾪��*&��Z�([j} 
����k�s�5a[�����o��Tc��@���_?�+�ɶ�%�(���#YڃG����{|ף��4��5sމ'�o�U�s��Ӂp��FE�4�n���zN�_�L->�����Dc�\�\r�e!�$��-�e��ĸ.�7��#`8-q��s��(
w��q���)��k��X�]ѝ)F����݅��ѓ�K�CR�1?��_+�@L�����6�����Qk)�*N��KE��z��}\��Q����P���DA푼��
��R�J�s����bG5��K*���~�̳������X��Ã��8�m�b�1��V�҂�=�'�$SL#�L��"vT��f�ד��e�Ex,��6�=Q#F���FUu9l�����3�TDR L�<:L*�&�G!�R��p�}�3ِ��Ԋ���.5��p�������>Bw�C�"��ה+ʲ���� ��NDb��Jc�=�[���i�5eޝ�F�K%_jh���Wִ>hI;dυv�:)�N��Hf��<�,w
�����#:�gk�y'�p��Y�~���og��$�{�����s�_<uy�LO;�܏�� �;�0�>�9*��:���Yqk�Ca��anW����*,0���;^�/;�O��w��_�+��`�V��z�E���_I��,6�[g�\�9�h-��6�����=_�b(�D�E��?�*A5 3դX1hL虌��a�����%ÿ,g�a|9V��a��r�"X��CW/z������x��i�~DOS6s�0Id]������ F��L$���l���h�&�#��h�|#�mK
�81Ԧ�.:ۛ�G�������;Z�M����l\Q��2	m�y�A�X� ���H*.ǌZ#����9������K$'�K��N�S��bZ����j��Z��S�j8�Mq�b���p�Jѷק��Bs!K����ۊ12;4�M�s;T}�!a�h�^S	�u�Sj�@b�-�I��͢]����n���E5]F��%XY���V���f-�q���@[9Q�tc��/y*ڽ�Am[ f�8$ϙu�YB��}0�N3�dl��F����Ҕ��7U>��ό���
!{n�^B#�4��Q��:! ��� ���d�>?����?�ݺ��u�C�u`��U��6�����a=_4��7�OU��*�@��x�E��(���.Y��6/�a �����g������z��O�e�j�:�Q-�H,QO+��6*Rf��vq�$�$���k������T1��/��'MT�;԰�@Y��z{]d��d���� x���(ä� +U�ڐN(�g�P�A��YA^9�|��q��m�Y��e$k�u�!Lm����h�i���)�6NC#��P���!wb�u.<1���7��������'C](���W�a��@R�e ���	GQ��c	�<v�03'W��^�$�g�2��i���������ǂ#�Ǳ���fn�l֊�**�k�/j�8�~�I�Ď�TF&�y, �~N__d�p�*��SG�C���k�'p�җ�N.^�TQ�\���>���,�����T�
�W���I����g{!M�Kjx��m�RQ��O��jEE�j�Q��;l�����0{`�N��P*�<�$El��t���+K�4)�:P�z�b�j=�^Pos���S
�����-�Ȼ����\O�|�O���sl0��w���+Գ��;a�ӽ�������E�M��)���D��l���ʻi��)SC�����wdר`��&��q�d �8^`�S3�6P�^p���KD�C�׏�c%!����t*�;]���Q"ա��Kw.1{�C���a�;L9J�e�A";^�(�*��s�-�q��H�8_L =���f�_=f�����C8�$�ÁY�,�_H���g~C�7��ڱ@g��֢�G��/PN+=N6��go"���=GL�f����@z~ޜ��9 �>�i��Ćla���}urs��OYq!Ag)�F:��N��4~�J�h3L'�1���e?6����n8��4\�ЬS�h��zĤߛ���,:���H�-���41��E݇�4�%����^���O�+�"�<����(�|^�K�/4���Rw����M+~�Z7k��FS�S/�,�B��eJ_��~����S�I�v�+�Ƿ��Ϩ�����H�9�H��.�f��Zvc��d4�w�əNc��T���řU�Y��hr@��x�\��!{� �F_
�{��)�{V���32O��2��F��|_6sYc�+��r��\-M�-gxO�����"L�_@&�|�6Mߝְ��bz�S\Y���Ү��w8��E	�a�E�������"\�ν���R���
�&%�f�Mp$�:CG?-Y,>~�M" �X���j���Q��0�T��p�ւ��P:a��s��eP�Tt����A?�eϵ�F�Fʫ���4Y�I�|Z���:V�������\���T��ձ�sl	b�����n���j�~���V���;��wR�����K�Ҷ���&�*!�齲�.J�0&Jr�7g�v����S�tO����il*׏�@g$`j�@�>ps���_Ř����V�����V�Bı�&�>�����*D�L��"� 	�;�>T���:n÷���/��U=�@����](� '����k�-���?�~O�x��7�6hD,��'h:��pU�|�8�J��s,iȱ%{�g
�Ҿ@�%��eB:��-��Da�~�L�I�I�	)�[*�#)�J�m,��>�'R(&-��,��Kbm�w�Z~��0��?�J�`S3j]j��L��¥@֘����gU!lI|�� ������i_`�Oq��I�Vd�C���6w����B/@kD�G��Z�W�_- :�����D��r��Q�9�c,�6��^����n8����@~X�����:��=��[Sn�E^~&�
Z�$5˭�1��M��*��(1g5�����4U�ֹ9���@/^��������Z2�(��`�Da$G�������~��?f�j
dXX��Xػ��;�	L����W"���,�e_t�K���mE���Fg�����v���I�P#�hO?��c�d�:ٺj��o�}n�<�3Mv�?�qs�5=��n4�g1�t7��D�Q[s��-P������A^���Th<�7���9WZB������iؕ�o^S���X���n�i��#H���	�]�(by(� ��A�l���x)6����!��)-PJՄ/��b��b?�td�xc[�%��c��^��A]��-�^�5�p�9�������.��k5W�W��!k��ͮW�=��Ȕ�}�|�Y�A5� .K�l[�5����jq����(�TI��!��8���~*n
G5q7qY9r��K�&�`0�ت�C�z��"�d\�"0�[���R��̲u+���# ���G��ﶯ���"�M}� `{�l������2�'u�@U���ۮ�{x��9�4TAA*����L���9䋰9�Y�(��&Pq��9P6�#l{)���^�p�l63c>�oa���r7ݖm$����W8����=(l2f�阡�a-����~�Vn�l�yت�J&�u�`��!��b 8�� �EM��I)P������!�g������N%�[��~�D�B�-�ȬnLWCHns^�\�@S�ϒ9'�Yd�!gO^4!f ��f�Q�������qN5LOQ�sNJ���Iv�Z�;K�;����G���&㪽
۬��N�o��+�!��t�U���X�1f&��������"	���|������f}�!�E2z�;"�2�A֟Q�I��J!��rAz&���)�(���q�uZ�+�!�C=�J,�굼r�6ue%�Kc�k�m5����kGP[B� 5A]���~��IO 9Y�2�J1bJ}�T5����UEj�x�'0c�z=I���\hR�.��%� &v��+4m��a��	����I�Ya�vH���]��Z��@+�&5=f#��L)�r۷�L�(Fy(�wK{��5M�Rʃ܄3ߙm$^/��N�^t��yh5��чK�������2�9�zR�:�L�l�/�=�:L�&}ܯč��봀c�W�و���'Q�Gt��)�oQ1�n��b�a�]���9�{/�RE���I�l��S�t���xF���@�I�ߺH���HB�T�p����Y�z�4��������xY%�HY���R��A��ui��d��/����C.�(����s	����e�h)FS�s��b�ʎEk' 9@�i|���%6TyG�rTlO�IK���C�� �:kSb:�G:���_@`.H�D�s��إ�#۴�����E��c\��Rj�|�5^ⳝ��ǒ��EH�l���ރ#��54h`
�{O=�ŅV����A�}HмX��R
Ek�������v���� ���eB�&����N���%�L�����0��H�`��gY����:�)c3"'�d+lX~�"<��ז�&��pE��<St�n�\G�s(9 q0>~�
�j�u8�*V��B\m����;��^��қ=-l���W#ơ����Q��[�����}Lz�΄C�~z�Ӹu~�a[%�{`�˸���֎X��'�M,�ֿ�,F�
�ŋ��������F�e uqƈ�I0^��������X��G��r� �*)�D��NѤ���DD�Y3�x�4�j�d��H��!`�Ķt�F8���]�I|Ug��~SL�/��#%�䡱,�ɸ�'��3���H5,���60�J��-D�+�ƽ�\��	����/�e!�����ߡ�J;h���������D=�!�W�o	�ȕ�Z.��.��G��;��� �Z����o�K&R�ì��y[Z��=�f>-	��՚j�XH�u���G�H�H��j	�P���Ģ�ߢ�����_�d�stS�����(�ihp3��+��V����WAX������h]�����G���IB�����|����ғ�U`�VA��Jz������،�G'ހ!������EA~wPђ~�<����r�D�����^mW��\(�W�L��tt_@����uG&ɚ@��v��%��� �����<<a+���?�����Ӫ��#��]�*�.iT{�S�n�s�A��,��B�l,v��d7R�A��`h�9��wc�ma,�יiK��O����ԥ�b���b:�j�6M�32sQ��Oc۸�d]ǿ4����"Q�͒��3d-_�ƻ>�"����ć�`tЏ/�c����]��%��g�ʭZ��v��b�7ʰ�.�;�qʸ������z�5��TΓ��j}�D�5�ƂH��Q�3E����P�$�ӆ�G���T�x�I���c �d�>�ý�l4Mѹ�XQgP���ZAV^��M?o��Rs��/[��od�g\qp�o=��\tN`G��K| �r�S���CZvi	F"�Ebu4c��_�����"bm,�6h|�aPB]@l��gCB�s����fh^zp��&���<�Q�\����Eo��&7�M��+�q��sSi������v����1�k���8ў���+���f|딃E�y�d/���� 4"ܚ�7]�ou,~�'��sPT���{�ds��J_? �R�k��<��-(FfQ�����dI�Z��B���7.gf����C���M����b-����#v��>�A����FMna=Jf��5]f��<|= �݇�d#�&z�ǃ��/c���?��	m̧߳?�U,� � �no����|O1��'��\|������U��F�amJ<p�<$�8��.��x�-m6�\e� N�p�r�7���b���U �4$�}�"���W�'��|��P1K���uU5Sޚ?��Z#����UQ�?�1���� e�� HO*`��Q�#ΰ<"Ii��/���G�-�p)&��1�$w��b���߽�ȵ���*��ï6�2�$��X1�����L�\�˷��\�"v��}R��L�a��S�m ��i\e�o7�2d��#� ��ـ6���ĒMEez]��_ِ=�"��3��9�,�I�ݐ��PzjVn!Q*獀654p�6�zqO���h���n*���GXk��
�8��.�î{7��D�/�	��i�3M�?l��x綄�K�=h�K;���|��Rh0f�5R�n��(Z�3ѧ5{��F�ٱ�g`[�)��m'n
Syz���w�kV����U�!�p�'����m߶�.7��G QB^AD=�Jeal�9����^�h��n���t��	�,$����at�9�U�3x-�`��"vY�L��T� ��߉�3��ۢ�2���=��d^���zT��{����3�z�{K��	�)��蛜�Igˠ�Q�G�cZ��V�CɃ�4ع�����S�I������:z��~>Y�QU|$��.0O��*@�Y9)�=��p7u���v���兌���(D�1���m3��7�@�	�k��J��4L�� 6mp���M�J�YȤ���J�V���l��ʴ�DɀP>^���5�!oBJ�s���~���r��7�+����9{����D��-�s=�1�����D@�q@a&�n��ؕ��fC��A쫗���=�Dپk�D����&O�K�~�<�	ZVDvrT�_�w��:��({%����U|���O�gr��A��q@2-���ԁ�͑��e�t��D�NՊ��"�J�O,CC�v�
�!�%+R���R���Y�J�}�| 9馘i�d�Ë���2����r��MB!��mHA�z�� �`s�MT��'�4���R]'/���}�m�~<�C��K���w,]"����1�!��:���n��h5䎦3��V��[���P�Ԣ"p�����Hc�9м)-[�EC���k૗�J\4�q��l͂{�+��{9>�*�e3,a��`e���E�>p�ZĈ�#�T������Ic`��V�B2�(�
��h���R"r�����QT�W�5��l`�^�9W/P�h��9��@��|I��Hɀa��ߐ�Z�	-�Z����K�5�"�:rUE��Y��GY�$���7�yW�y�9�m�R����|r`Q�8�l��m����^����$7���i
_K^y�:/ۋ�thDϧ<�Z��=�"O�M�UE�K�:�2��B��#j1a:s��+q������j��NA�~�;H�쳏Ko�c�����Y�f���MŬzI�rR�5Z!wJ����Yfʖ�y�v��`��JYWl���~�DE
Ɋ˙�gx���j���6�VٵW,A;����ձ�48c�L�פu8����,15�G�MF�PRQ��Ph.M,�#�%��m�aW�O���\�)'��\��S�U�$�B���W�9��I���k�r�K��ւ$X+9�Ӳ�I��)z�ǹ��P�"G"�V̵.15�>�h;n�l���F�+5iK��O�ˀ4[j��j��I��IN�Lq�R�<a�}$j�o�4��S�U�V���Z_��]���l���p��f< ӷM�|��WZ�D��zV��eo��x@ɩ����h��a&��Nw�����H�"�uې�9�;8_�*�蝱��6<��liឮ)1ꕭe̓el�O~h��Y�<��ˉ�"7E8���gI�L��,���%�_�6O1��pAٮ�>I���?�)�ʼ(��*���{|^a�'\�`�o&�j=���AW�B��mruWW�Z�d��^\��$�7�JO@����f��L�
���c�����`�e:��YQ}G,|J�P{9z�'^��K��
c�&�,K�X���=Ǒ�x��8I��_P�������N7�`	�/�D���&~�˨�L���P3�YkDA'��~6���@Z�q;بj���wF�ɩecm*��ǭ�3-nP|9�$�/ᐞo����D�K�!���%K�#�Utq�=�u��j�	����j��dYWP�,u�;_��.:�?�%Y�G�����i`��G���oe [��{Q�B�O�5�G�!q1�?�Vy���)������B��Ա_E����7#C�"II-����G�}���j��#�y<��J2((�����6/j�ޓ�ы������E�$v��'��?�7����0:�����엲6���������
����M_���#��� �H��8�x�_�1Q�������IOh��@�[�V�-�/�uSh�������
1����d��/�9[��(�[�c��i�9�\>��v�ٽ�.%�TBV&�_��
[�L8s�:�e:��ՋJ@+�kE&щ%:�U�� ��@��hA)�k�G;-I���b��=%����dZ�T&6�﷾��m^~h ��>~�I�r�m�2��}�c�C�Zi,65�fѭh����5����2-P���F^���@����g��KcYUG�f��7\���wݑ��A�� 	�J@bi6���+���^��Y�n�����aH��=ۿ��"�P�4%������q^Rt�OO=����o�	$��:ҕO�8�@աd��~���Æ����������,�!�K����r�l��3^����ͧ�ObU���B&�q���p^�h�#@�	�s�[��p�_͎v����?�B�{f^�v���������oW@�a�ǂ�=Hy�àz�^�%��]~Wo����մȶ�#W�uw
�ץL��P�\�b�:1�����D\�A��k&������]*h����%�c��Ѧ���C��`��A��D���u���m�ƁX@Pu��\2�X�����O��y���ׂ�_���>QK*9�u�T�Y&�oY{�%b6ti�ҙD�!�0j��ҍKZ�HuN�X��A�C�A�^���� �2po1 �(�N�O��co���h��|��]���0n�t���7&���߸{DJC�M�fv֒� ߫NF����ce\���"eI׋HթY����o��Еʷ����\ ��5�#�'y�A��b�CxI��&M�3��;��|h�<�����X�laKF�� &�f/�*�}�Qo��[��ĩ�"�5�No��ʑ:�)Jj�qk�����Q��,�̀4d�bܤ�c8M׌yB]�%F7���oiA���O��N���xf@�O��T�7c�Rf�)Gs"6���K�ф��.~DKФ���.ġG��o6���t#k�
��=��]A�PoQ�T�c��='oa���w�Fg���B�K��B�ɡ�ў}��x�%��a[4�M�`9�Qs�6S�$��z�Ji�����(.��oאP_��o.*�g���U�c �C�����۲��7�Xბ
9OA�6��p�It�5.�o�5:�|4̑�ݚ�9e �N�_4�\?_��?1��~�L�8��g!Ĭ+�P̹jyE\D���Pjh6���w&OOfbNg'�Ω.CXZ�Q���@_%�lZ�\h�5�<�d%��1{��o�VI�j��� �]�
N���=]���b:HT�a�4'Ue��*=P�2cؚ��pa.�����}��9����m��U����Z����� �a	��bM@�˥���읉��o#`1ۢ�o�9-B�Ma J.�d�N+P�*r�gEI��j�������ք�+����Ŵ���#v�T���4q�C�<�?kr��w����U��[�z������Ѳ�0��O���r���w��τ������8r��#�b�
��[J��ލy�UI��]T��Y=���'��gUQkyv�k��6�RV�Rca��E�b��g7����Z���2Dr]:�h���$�ïQ`��F=��#��#ڰ��q<��M����-�;�7)�=��xER��3�D��hj����m���Uڿ��y��%G���5�u�]䟠�ˎT����`��%D_�B�_�c�`'�c]��.,8Q=��2a
~��Gu"���n^�׼��&aS>���l_Ujӈ����p�\�����U�q�A��dI�la��u�"�.0D}� ����P�Q,��<u���}ʦj u�Jl�m�;㥳�ҁV�,L�֪�2Ԯ�������B��8(׍:�|�b�1�T��i�/f���IAڈ�V�;i�b���l���b��g}a���e��]�=&�g��@��Q��T�IƶK���u9{��k��1\=�K0����ܹ��Ć.U�6�T�QBv�����W�P-�C?�G��^ ���1-w������4�lkf�'E����5��ɖ.�Fv��ڈ����ɛ�d�t����"U�Us��m*�]�h�`��(���Ր@���|5񽊎J���V��t󜸟��`ם��-_��_���T��7Y���Fqǋ�.��K۟{!�2H�;�^���3��U��+��m�#	��숡��on��gN]����g�]�C�(2��D(��=�p��X������w�["W^��Ͷº��C�;�S�ik"�9��q�t�3��=9�:`͠p���.z���L�De\�.z���`������8�>�\�\�ɠt.;�@ ���Z:�>��p�����Bz�#�=�U��iau"`Q��������j�԰�H�H%X�?�ĸ��VC��I����,��6,1�CO[�`-�~=$6͊:�� �2� WRs�&��u����]iݥ��Ə��)��<� (u�)�]&��㪿y��X�t0�j�x���'�Bo��ςG�1WsP	s�i�'.�6�o��JP�L����;���=���N�������]��^UB3�obl�9��t��!EPc�yQ�����2�^q.֪���$�t)nwrD�%�2$w"A2���#��T2��K�-{oܚ��DD�(�y��DGO��.^��]�h�� 3�}���1 ��5��G:�Ο�n��u�!�����M�'���D�a�l}�q��mH]��G�xo��"Lk�}tJO6�~:2����'S�u��$Ul��TBg�K}�o�k��ޗ�cσe���g(��el�Q۪�
O�,�����w�bv�~J���G���R�M�� ��@�<�ߛD���B���9G��aR:���|<��>}�ۿ5��֓O!�T�h���i�hpH��޼�xQ�-��Ō#l�W�?�R?X��1
��K�}�d�u_�1���� �(�;	��\�f6���,�x��-��r*�!�#v
dV��em��Yk�䫜t��f#q,��)0��Ý���p�`RQ��\�IŖ�C�:�0�a����V�X
�cYK�=�n�%>�
̯
��njY!l\�o�4D(/��"�z?�P�0��X�% ��uj�i	��oBs��(&끩
�<��h���D4�7�C_��c5�"t��R�x�{�g��r�C`Sz*�|�������}��l�d�)((&�p?�铀�0E�>"��� ����ުN��p5���VpHhT(>����q$��kc����|%�������R :�D��"��N�*������J
��e�+��x���$9`�L3ys�����<w� Y<�k
C7Ü(=���y70��\@�{m�����f��:�T��5% �R���a�4�8��Nߨ�w��Òg��=.���6����h:vua��ԁZ��xiv2"��J\RNsc
|y����R�
&��Ґ�0��p�Mw^I��L�������u5#����o� ���lʟdl�V�|(���`�����J\3>��T������w����n����az?�_FC��c���έS튡��P�u{�cI�QU�؟����U5��;�m�tBT���Q��+�m��1�$��ּݳ�Ǳ[���>U�����1r��?%p6�ˣZ]R���te L1R���F�j����]z�x5���;��2��Kc$� +��g�,���:�JlZ�4hi��Q�03w0
Y6
z����_H�TT�����~IP�A ��J��f�Q�4�1[UX�8}*��m�@M�)VY�a�B�ͶQ�r�e�6۶�@�9�cs0ߔ��N�s�� ��������1�uC��tEʐl����������7�Gn���%d�	0̬aҪ����G��>8}^�e��c�%9s��dq��W� Q�U��U��%y�uE��b��A��<"�l]q{��e���Ǿg�����;��8|��w�S�0�\@Hy��_ /:BS�����{�74�-4 A�Q[���T9�J���F\��s7Op����X0:��A��Acw;0<ڏoeL��Ҝ�H̶��bh=.v>e���q��VH�,C
n��L�B�]X�Խ��23�(k�y��`F�գ�g1�ێ�,l���˹�|���Yjj�{;�ۈd�G̰�.@��t�����e�o7�{�2Ƌ���an�y���@��=�Ws~���`��)u�*]�Ŀ<{I�#}����/���mU� �<?3&:}I���K͌0R�Z�%��[�op4�U^(:KxEY�Ԁ�-ܭ������r���z���3ϵ���T;�d1-b�B���gb��\�26L�;�������� ���_k��rܫ'VN����^_�����8m��nu���I$ ��sV��C�����u��JȂ?��� �yn+#����Tf���f��Y���������b��z'i2��a������@̘�	1��s;�'�O�S���bd2�m��	��?F�<��q���}+��]�����lF�h��v�.��P�E'���/~��k�tGh��9�fP)�:шi�Q�#�94S&kn�g[F
�+ǳ�0��t��35�X|ˋ�h7cɫ�4:�+ǨS�817IV��x��9jK�h�3h(W��"��T,[msE�b	t96:�.>��}����z�=�PP��.��։���v�bU%ō�8e;�w%�9�9��B3M��	6m��`wfә���k�~I�P;���hdN1��-D�S�GH�l'^�Z�<C���N�W��ɒb���J9'N�l���H�����5F�A�Đ�e#��;����M`�"1���e�@��D��cw�z��$׉w��(;��q�@k����`�9�.�V��,��/s������j�����"��L��`xw�%Ar޵ys��Ҟ��
>�:��qJ�8P����t��s.�k�~: �z��Ѫ��O|�m^�r��jb��-Ȅj�١�Ε�X�" C.� ʢ\��4I3��/ה`����|oq�`�] �խ}bQ�q�Q"��v��s�8F���|zx)E���d��C��4�ٿ:m�X.��;���f�i��g!4t�t? �	�`��NG��hc2���.��M���2c����uM�-(�l��΁�r�{�X�1�k��ϳ�q�'/x����(q�)�\F��d�N�I�\��cP8>�S�@���܌��]��)`��f#�U�[�'j���R��S�K'����а4�$�_p1>e�Ϻ�t��ߺP��x/X9E%��]�g�;l��|?$�05�pP����"#��vox0J�0i����;L�T���0�@�J�m�6�]w����%�ƽ\1�K��2P<�j�.�-��y :���U��dn5�j�����XF{e�Q�h�x�y�ws�C�C�F�Dxy2�����,�QۅLf_ ʼ����eG��"ۗ�C~�O@X���:$���G�a�M��+�Cʃ��`�1ڡ�K�������c�
SHj�����`� ��g�$lJu��x6��["A��#	9�c�s�w/�ʈ�'t�)�Ǥ̦?�9KH�*:���<������;e�
b
�c>��S�Z�>�꜎p�u��ΐ`�DETY�r+P�ҹ�M������BN����WG�l�S|�z��g8H�����������;)����r��˼��E�)��=^<s��� �A��Ul�@u&�*���f(��;�������ߧ��Lh-��\�e ��+�
�����8m�	���m���nW��.i���(�eü��\}���Ȋ�W��^+�׳σR�)�o��c�	��j9eU�����I����%����3.�����=��Wb���0@f"�ϩ�KZֺ�p+?2��3���* !N�����
F6�`c��0"��1剣K@X��9�M���˾]h��mB�C��^���$�	�9=i����F��ʢ�����c���� �.6�|M��*J���</I� ��8��z�T�T�7���q6� {A�no�N����Pj��+�-��R�j�ԕ����1�����%z���u�o>,���v�/Ekr?�Ĳ�NN�Û�n�y^����0!� ��[��@U�C\#/�Fp�\�5:����-<���(p��h��ݴ��k��\d���ě�ߩST?7�)N�(��;�	�'j��0Q��t/}
|q����|�@L�����[�r骴���ιK[$`�k�)�L��K�BHx������"��{��;�i�g5��A��W��/��Jw��+x�c�=��b|�D�o�'��\B��qi��q|z��Zse��T]H�Z�S�DB���Z��H��.;9�xYp�I�:�g�s� �F�;ᕜ�᏾P{�eNj6�%�#R�S����$L,>���d��R��\]@GTÄB��:�3���-��,Api,�Y=���O�I��U1|�ŹYB?�|��䖄���g�am2O�@T���&E�����d=�=2à���m��Ynr�BJt�;�ˌ�;%0�Ҹ���u�q�U9�/Ԓh�ޡ���)r'PR�"v �)#���5�9i��0�j���=�{���n����Ow6�m��gQ��ɂ�-aO�)��ag��w��P0�����D���@��g6Uɬ�r�"�� ������ �fx�|;�U��������:���gT�E��Ó��d�H��p�K�/���W�-��D���S��U�oo��lr�f�t��YU���;���z��rv^7�۫&n�����~��i�߭np� ����ޗ8�Y�\˯2���	P#�ik��D��ҽFo�%�}@Sy�N���~��%)�!ږ����O����*� �Sw���!�~Y�*�Ґ݆$M��3�9LnJ�^v�4��?�P��Eo֋8[�D.�rf��w"�ʘ��d٨r���J�TT���������z��*( �>b0K_>��X_̺ᒔ�л��ܑI�}�)�FY����ok��3�Rٰ�zEb�U����C4m���Rԡ*��H��9i?��kO�ےŀ����fV��݅�"�2�f��-�#�E�u���$k���\~C� �����zoTp&����_��,r���|����`�,T2WU�p�T@%�"]`#+$>1A��Pʚ�(L�T����p��rjƭ��Sֈ�by�uʭ��D��8`�FCe1�`�?H��d�GI�X��L��p+��׾9t��2tw��vm��S�E"m�����p#�>d����i��i��*ׄխ��jWZq҅J��-d#jz���#^Ç��q�D�D��#$�D��1����Ʊv�fEy'��(�g���a�z�)������<2�gW�gT"�
���s������*!��5�
���p3 ,����!/������}H*}@�t�޺C`���f�@�N�V��&��z��*�/�9�<��1}P��;��Z��kԬ��cY`̈́&��>^�cG�� ��L��<���(d߀ZU��џ��f��%�z�Q���*�8��:Y�_���H�K��
,�죢aEʝl��)�Mj4��?۪�:�1���f�RB0���21崵?����������pq՚�)�V{��9�q��
��w��b]��p�}/��M^yP�mQ(��U�X� 3�5��dI�LtV:{�]�\_��)��c�b��3f�e�Vq��h樓{-U����Q�Z��J�^_hW�z�ŭ�J�Μ��#�}�X��&������À����5��ϫ>Nn�\A8ɏ�"�j���a���s�k3��Qw������>��R$�"X��
����I�7Ktn�L��3ʄNSm�텔kNd~-�!�T��b�9����_ؾڟ�9J��5�8����*u�oB���=��)j�}�y
NF�{����3L-1U��Smp�d��
��6)��.
��vPG� �J$A��5�Ps@�u���*�h�e�5���dW2��>/${'�K���gq���dTV����l5��ԭ��P�n��U5u��ƭB�5J���V|j�|�sN.�����;����Z���=b�uc0�ߤ>W��f��ɳ=6C#�x�dh�蟜#�"B���(�$���iR�	�M�Ī��?˝��%������WҦf�-:v��Q�ّΉ��m�7y�,u��P|�ܨݕ,Tmx,T�(q����l��/&ɠ�����pW+��U��BQ��(�Ryt�����Kb�]�Ǖ6�cF�L=������72���g���>)��l�m���^�̊
Y'�F��	6P�a�\9�ڂ�)��`7�M��cu�{؂3�pM���3�\����@U��y,wo�+Vww����`�#`�>�Q�4+����N��˥�J䤇��;vS�ўLr���1AqG���	7�MΚ��J�p�d���, O���x���Y�x�|���w2)o@;�m�6[�5t����������?���N�w�vϯCFc�r_��o<���fpD��f�3�d
����ܲ����m�x�qbz/�8�%�濝�N�˱��K�EH���oeC����Q�+�O&��(��L�m{�	�����6�A��.0}/�r�`#�c��<����x�}�L_0��d+���^/���P���;�>��E����H���X6�6����K�˼=s,o��B����kd	g_�[��^��d���'�Kp�4c :�E��ie$mz*b���6�6~��w?q��7nY������h�E�\a�QtV"��
�p��cX{
��j1���v�`�ٍ��稺�B�Ex�ȳ�>����t�	��y��&|�����f��]�y�jԘ��u��,�g��L<MV�����=S`i��s����n2�|�G���d������@��}��0N
��=�&J�|���j��ip�p�b�ʅ&�����=�H��	Y�ѿ� JI�F�b��-��UQ��T[oLM�A����V�Fj
���-w�� ńy�i=ߞ3�$N8�V���~(l�[_"Aޢ�1�|�&�p)�)��9q�ҭ����AU�C�ڵ�	c�S!��į������A��s��JK��R%�X��W�vnJm��gR��P���r��s5PD"���Q	��6��rn/E+LA��(�7���u�S����;��ع�DY�򼘘����E��OC����+�Q�:%�9���O�O��JBl������=%x��k���~�;�d����#/�@���g\����IK.���.aR_��}�1���tlX�b��+�T:y8�9�����VDC��^�yF���_6��$�Z�\H���6�L��Y���K�_>�:΍#�_T��\��#�_��� ED�W��ef���X���:
��HB��7�냺h���Z�m
4�(SP�*��F,DM.g���ݗpY� �Pu@�:i;�B���gEiEUɛwG�1ਹ�kٷ�f�}gX�"tg�KP9�i�&�h[�ְ]x�m�7�	�%Z]�Q�N��	ъ�IY����/�X��+F�m�N��YkA��;������� ��@]r�"{+O��ۣ6��7�(�{ �=E��虍�T��p��}�/�ڦ��]i!*���l�ɸC��jt��D�s�����A��#�t,�����ɍ�!
�cĥDu1�x�g�r�&�|C;��˰aw,Z�	�˾g��yM��5n#m�m�ɲ:�\���� me���oO�>��E���	@=�ulB��U�P3�zĀ�1a��뇪I荦�A�k�%�)&O? �
��[���jKҹ��\g�����[W��/�y�l�t��?D�Q;v8��\�B7�L�/nLb`�Y�6(<?Iba�эj�fJ�gz=�+z�B����R�߹ǠF������/��y��|@���Y�m��~~j_z'�j��5G�g���]�k�� �4�.|J>�#�N")Qw��x�W�R�}��TM�c�P�H��̗`�T=S'gK��B�S{���P���9��2W�l�j�&�I�D��+G���u�V��6�:�i���V�tg"�K�{Sk��� U�A�/bڶ`SR�6��#ym[s�,��F�ؓ��bk.�������a>�S�̓�9��Wz @�u*Ux����o�[��7���,fPEd�c��=)����j�ÄcE)�y&�;[��C��7�y������	�3ǁ�.Zt���Y��D~h�y?�3�!�Ag�Q�ы1 �eD�RP�r��9����B'~����X+��u�푠<��^�",~IN�bL��
K�v�G� =�O�����$�Щu*�R~)H���4h��+ɕ�|����HG�{��p���hd�jqȷ={hS��,�a7�=^��"S����d��;]�w���n;O@8Ȼ;�s-Cn�x����:��&K�(�Y �l ��	�>LR󱹔���KF�;����\�rR.��K��{��"E�?Þ��9�L��[${7�g��t�߆�8N�XQ�Y��}���=L#R�j�u��-�(yh�c��gh�K���^�e����U͙�va���y���@�����$z��du%b�\��*�4��rAmC�a1�F5������giK�:?_���ߔ'� &<u���Ui��V�;g,I:B��eӃK\�$�۝��{��kdbo!ߺ���>=�ZKo���>�)yBO˻�a�2�2e����]b
vgEw�-WC�H�q�Lnђ�Y((�)mv�MӘ{u���Xh��']+��8qՆ�I%ذ�і!�:�ұ�D[��o�n�	x^�kŚ]�8'�=�տ]K O_Ad��΋K�+�x>�����:V��žI�6�;x��^�{N�1��6��/�U���^;��a+��.�/��Q0d����X���n@%`��.~��J��uc˯�5�����6ht;�!b6qk���Q��M���f�a������/5w\U�EM_;]M�b+?�O+���.�է'��'Wwv���`���<�}�"־���ꑮw >�6�T������zŉˎ8��i�i�3�~�oq��8
�������R�v�ž�ؖ��e�R����g<�yb�|7�j ��qC�y��]biQ5	��z�9j��l?�f$�û�Wu#ܷ2��:t�pj0���A����0o�� u���(#�*��������NX�������H$�O��gD~�m(�{cU��H K�ơ���Üs-8�:F�����޷~��"P��-�~f�y.5�br�IUo�2c���ADz��D|��/k(��6y����V��{mrǃ`R�ؙ�pJv]�&@��4��Zk�ul��j��>%F���He����0���� \T�l2^c�(�6�̚�s�L�/�D�N��2��T��
h9��/2��k*�h�j<�sDbRW���6��h"�zɛJ�H���o:�HU>��q��A1��#ҷ��������۰瀜�prmf���������n�M�7�VZ;��q��T���ϡ�$dx������0�g�S֙
���~g�zȠ��RA�:"�i�5��\}�e.[x6k3~6��=Q@���A��&�l���v_�o�#r�f+ݟ2�<x�
���0��=�&��??��8�kQ��]<�D��m{�*����};�ߎ;R7�Pw��x�+��=2��漗WXq�ٿ_Ϫ�FeNz��T�3�).����0��{Gf����{1���$���J���	x蚣N��\�m��΅h7�76`��7Q�he�F� �;a�P����LYW��� ����S��M�-���n���z"'�ȝ�X�1{|�k��)$VW�N�Iϭ���wY�Y$ �{�ƛ����h#'��t,;{`�6�(����c��ryQl�5]��?
�� �N�5a�zC�r�Q���8'+ؚ�B̺Jx���2چ�~"&��5�/�j�]��M�h��5�{7l��tQE:�?%��|"�t��B�bt�t$A�vʳ ԪHk�+��[D�+�P�Z��g!�>�M	+I{��N(%Y`򃗉-��C�� |P�@���F�"�	U`/s��躘�E=>�����#�(U�p9rE���.�O/}�m���srk��x��0�]�I
5&qmd�B��������%�|Bonjp��r|� )�a;��>m�MC+(O��D�x��Uj_�L5��>�핥r)�1M�M�5��9������77�V%���d>j�!Sx>�@Cþ��ɑ�1Zx�M6�꒡���C�|G�9X����`B"��͵^�u�瞇�#Twp0�-S2���ז-��I���4�r{�3�=hx��j�L����+��YLCA/�;�[�U�QL�wI��!nա?��Ð\A�{�ӏ=�꺍7��a7�th����dQO#�<��HQ���1�_D�}^��+�)�5/Ү�i�k,�[޴e�y���̚��C�Ev��ʒ��dS����ۖ��U�\6e�"�R�8(�R:s�j���8�_����H[��n�f���Tr���	Ś_	�7����_!�n@���JW�A�VN�!!�8J���Bt<��>��S8:\����¾��z���B�_9?.�x�֛bxԴƈ]��iO�� ���P~���y��r������*v�~��?\�ږ������[q�K�r0bW�rQ���"��nc����)~�<6�'����a��|�걦$�db4H���g=X��;i��J̯06Dp<�az����m$89+E�p0Zkn��.��|HgV`/�������w��ek�T��}�i�c�쭞���<� Àz����%|{�؄��3W�'�ܺ�� ��XR�yo�Yt
��^#_3�}�}ƴKt�o۲h�c�H�
�D��.��4�2�O�z�Fvw���[�sf|]�zL������GH�O�-�,�h����Y���R���QG7�͵����Z��q��ޓbN#�v�΀�1]|3��Q��x�4�RS�WʪPC�0���B�{3e�/�#T5W:��5�����ZX�Mm5X ���YD��$�BfRc��A�.F聠D�0���+�E��23 P&jJ��ó�ԟ���R_hR�w�R�>/q<k=��(�F�2�̽uI? �0eò����غuS>��ץL����\%�N��R/]��;��"(���Fː*��1�*o����2ya����.�����+H�RUP;��]���L�G��gBW� _�5��Q��5}@�i����=�-獎���}f�2�ȜA8j�ZK��i��q�-`Y�IcJ�{3C��� /
�gJy=���ћb)�Е��a\X��$֨^�lf�S̡ߺ,�G�"�+�^M�3�V���H7k݃'(��|Ɗ�j�B��}���ė���Ŕ�ii�B�@��B��T���w� x� >����a"�k�lv�U�h��M��4��P�[H.��I�X�Z���[��Uɟ���4�EW۞6�7�
~`��')�5敯�$��1}��)#u�"�F��շ��/(��-\T`0iG�y!�h����0����p�_�������:+žC(9��]U�&l����9b-��j��c\t C���E%[�������&���D��e�uC��T}�{�:��#����]�;X�KUΌ����쀉�lB���j^��6ݱ^*�i���G](��4�Z��1c��E�`7�4���L�{1�d��,�6�~�e�{_�+

�w֔8A=w����I��m ��O��?D��2�_}{������ZP��>Ts'����2��o�GY�2������I�xS����c�����	�����8���/��̮D�p�=p�b`���X]V�~e���8��[��6e2�!�Or�����gF��yq����01H��ض�z�g�h����+e��"L.灶)�ʵ{�6�� ��D�n�f��d.&�A�[�=��5�LKf��t�]�o��R�7\���jAa�L��A	��%A->�VL��e�3���3�ϧgC2� �W9ς'5�!^8Y:3,��sP��A�pŒ!=��P:h`4���U㣥���.\,}��5jۼ��ܳ.��!��n�]���Q��18I\�Qz;&��Q�0k�%��&/�D��{�g�$� G�g2�sH*�����Hg
�d�|��g�G_"?�d�
�%bv�����tI���煅� ��	v-�V�L�0��� Q�o���6j�E{{٢�0SV�ѵ��Ym�L�#D?��]��ԫzB4���s����GE.��(���^��Pr���f ڼ����{!b��F5dM�ȌߌAqB�كIy��>	)´R<�kv��+�:�7�ƾ��,��R���4�툈�>c��@:G�&��!a�7�_m�69���n�~��_�p�^��#�zY�Ҡ�*H��m�1j�I��U�X�+��`�l'M1�tJ�c^l�
��݋��y���k+�e����ʩ`}�ʜ�*��b��q�T��T��6!�!)u���<u��cU}�~�:�,h�E����M7�3hS��kg��M�S�%0��-�֞�����$J����i�i5�8�W��golD`\��euBm��F�X?��F�-B�r��r�FK)��_�����ˍE��m	�ƣ���)Wqc�����S��O�	��X�x��^]�ͫ(��U!Cbp^�A�Q
K�1�(-�/��[�=jȖC T���e�e���ǾsǾ���َ�00���&���>j.
�;ݯ8)��{�F�>i���:"�mr�褶D���9�r�6n�x�X�BZє�S����-?��a��(Ny|�\���Wc1_��g����R�s��ԧ�I�=�����J���t�%�����X�_qp�+�Q+Z�:?�/���0�X��*V=��FǏ������^3��8��5�'�g�I+�����S	��ր���Jd�L�E/(' ��!�7V�? K0m�7�f���pGz� ��6Iǳ��`7齶t8~�MٕQ`�{8�c֒!��X��LOPc����Μ��;ޕ�,|�d����������r�<�
L�������(���P�{K7�T*b'4&M:� A���. =e{��Ѫ��S�z�^�D4(��2��N�־���>ɐx;P�2.$�HFTW����������!~��|���S.���x���OT��
'QM�b;`��gd����к1h?�6�Ks�U��{/A��m���sDrj�a��B�<0�熊�-�v�h�(�z��=:�_���|k�YV��p��O]�A��63����FI�I)�-��~)HTY�$�����5����Q+��1IN�� �l��G�c\�tgŋ�@��,Ӯ�][�r����H�(���8!ĸ�O�厓e>�z�;TO���m`A����ͷ�ܫ�|7λq1]�
��f�� z�a;�a���[�+U�tL���/�-�k��P����l�D�;@�k�n�Xx*��F���A�~Iݠ�B��8�%�֩�@��|Z�)�a���O�@��u�,�E2���dP������\d�P��_p.=(��"j�B�/��υ��?E*D	rs��a�&F[���?hIS��A��ך���J(l���F9�#v� M���w��=����ֳRJ��K��+��u��w�t���A�H��N�
{>�ĝK��E&Vt㉲t�L�VWҾ�^k����r��ɨ����g���ޣ)��7h����Ĝӭϼ�S�9��A �*�~^�z�b��A���gD@��LQW3=A�?�?wl<�Yr0�B�s=
��ww��A�F.����F	�nm٭�*�����L�H(3���	���q�K��?W��̛EZ,��o��r��|��2-`E�p���u��Eʾ)A�Ą5�Vs�mn��킟�۝��1���>
ϐ��v�j����C��
���Ь�Vs����f����av�����>�pޛ>�dtS[��胣D���lp�r��x�qi�8�����o��o-��R�Kؼ;,Vit�L�)���s\<)X�;H �YAo5�\�Q�H	˸�/��<��W7�б'�i*�މ�.���>� ص�|���y;�-��1�S,(v����T�-��7?�痩�-�5`i�������Qd��!dIYP\�<�G3!��7���ז���K��&������@�����G���S�i�T�tn�m��9�!*�Cl����	6��abyj=�hŊ��z;Bq���sYp"Cj;��8�*A�=o�����x9�A;�f�|܋^1p�X9
�/ߪ	d��P�2H���3/�?��#�\w���D����Cy��RY�z���qG��	�R@�*�"�B��Ծ�I�j"�����`�4T��e�X����B{?"��۵�*���i�q{�-r�)��~}�zG���b�+�2����IAs�t��=���R�b'�����AԬq�Ln�|���ō�$�P+��kQ�K$�������i���ֳ����=NV�ئ<ǂI��{"Ï��h���m��oˋ�6^�f\�Ι��W/ϡ��=�8
�@ �:Sr.���$���z�5}tM�Ve" ��B��*�	���.��J���OV�u+��$.�z���	H �E���&T�ePG�&!�1)0�%@��R�Q
�Ս	�=+Dl�73���tx�J	�=���hn�����(�ۙC|�n�g���i!��}�+bV���7�~KpaU���#�Ĭ���}`��� ��=�Х�d"µ7�<e�4��� �<;�i�=؂�,�5�\[U��� ��Z�4VP���8�H��S����e��vL*}��]�k���U���+Zy�c�S!w�23"��{�����[aa�e+3Ԫ�q�&��+ �o���n?4'�A���6Hz�)z�L�y�=%HǉZ<�^؈e�O�5Y�%��l��w�����| �4Pt�d!��)�yN��Vj0�ߛ�-����KU��1���g�0�N'5�u�ŠZ����ɋR�z�n&�θ���}�hb�P,��4R��m���
o�i�ckAI�O�`n��z�~�������?�&._9�}G�)��U6���1;x��α:6-�EY)ٌ��
b����qV����Xmj!�������@Ăy�0��<������]֎�tHP��\3:��L�A�����Q�Ռ1�,�=|?D�f�]Q�����z�Р��]�H��1�̢�{�$+���6����~�>r`Y�_l�N),��9�l��%BH<|�|�ĵ6$��f��?���pd�ְ~�(�T�f蚭A�3��_U����S�Z=qၶ�>���s���~��
�g��H�ZfN�c�2�^7$.xV��:S탑&�nJ�tyX�c�� �ylE=��8�YBA��g��]�A�'|���ʨA�"?@��W\Ḕ��q��f-��߮@=>9m�������`6�\2#^� v=��1<��dw�����T�jB)\���6g�p�.D��Ɗ��̊F���
*���ʻ{w�te�گW���T�q냙��
����}��+����U%�п*��`;�:�������ɠ�4G�1�x���O^�p�BK��K��3rJ��U��=}M������~�|��k�m�~Ѐ��u�ҹ,"x9�����Xd���i9��趻=��JZ�T�L�b�3Q>pQ,�@muL�Y�l5��&��X�z5�m�7� C+F7�{��!���;�ü�PLR15�BT�&�#͸�^��p>�����BN'���e����L�/��~�''���A�P�n�C�
�l��g���������:����*<��\�.R)2C��t����9�����@�����$����x�'�V�8��qQgDbθa��w�q��Inf~�u)wPy��ԩ{�{���(��&��à�KO�5� R.��I�j:�P�%k.8ah�0��D�Y�s���N���G���|(����|ͪ�wf�\#꟦p�O�.SIM��2P�6��}�fθ	,����2�y!,�>�� �����(!~���'[@v"fJ���Z�XףЪ��ҥT�N��STh�Q䂁�v-��֌�e�E�
�?S�6w5�y�$�@��6��iZ�_[�q h�n2s�\��p*���޻`���n����	�Q_�V�1���G���\*l<Z֔���}iM���Y�;�y���."a�%uッ"b����@E˟��-ڲ��ܱ�C��=f������rkbՀ�))/VKe�	����K��$Ì ΋�)"w���$r��N'H&J,!`�>6�v�w��?=: l;ڢ�{_)�y�3� ��Oa��1G���L� ��<m�a��\��Pa�VZv� k<�jdap�|U�	�n*��EO$+�Vr阘�Vt���F4p2I�\5\� �;��[}9c�$#�}ޥu�P�}�ϫ�\�����c$*�<��{��Ȓ����&#�+z�J����j�ע�z����zjX�՛�,8lT� �b5(����)�tg�'o9A_bv�.p��,�椑k�.P�6?5��Pg
��l��0��l���M�:�	���+����f�k&Uڠ�a���o(-�P�g0��;����ktO�H�l@A.k��.xG��^��c�m�?B�����{VN��f�O� �@�
VT��ʵV����wR���g<�Y-Ϥ��~�/;��i� ����^�ܣ�l������%��:��m�=���I����U�1�y� Μ ����G?�s��=��s�D<�X'�wUj�x�c��������0�Ƹ�`. ee����G`:[8�P1@�s�df��_j�ӷgcƝύ�����r(���?����$�p~����{�R�G�N7it d��> s�/"����l\�jEBZ����ZR�'�\�F?�d&t�F[�M�y�|c��;�A��y����.|��3fcz�0�D���@0�B�p�������,E���X�w���IʈLp~�g|�wt�E�P��J�qv1=�;����tSnd�#��J�r����96,��t!8�̲MJ�W���	��jܟ�Q�j���W�46�n�q3Ћ�vl����u�Xn<�Pٽ��%��ӱ���8�����jN���X+.���I�Ys��p����-�����(ǳ�<���?�~�M����Eh��'4 *Sc�[C3�LR��ڴ�;^��+JF����}vc�P�t�t=�+*JAi�7G�X�{X�h�~	�O[0��wo�6R��Ԁ5�����ӫI���R���T;����s]����?h���\ '�M`
��o��Z�FW����ER'��\�1�Y���e�-��qH���y�%�����Tpl%�S"m��oe���J�����rɅ��$����-�:X�?8�p(�U�Vu��߱aBA��s��"<
����,�cT��[��y��}V�E��@1 �~�̓l��R:����&��p	zٻO��4�!H���������=�ݓ�5֜m�v�I4f$�\�e�8C޾zz��$��ɹA����Dd�\zs_��΁�+�R.b�w;��9�H�hIr>��� �LG��ԗOSx��YF�����}CnA����Z��:�V�\���+�Ϩ6�r���z�����J݃݁J� D�Bq���rY}��X��ջy�E���x}�8.^L5�9�ضrm��)h 2����+ϟ�IbS��um��*�!���Qa� �k��,_�0vB�N��9!8ܔ�#